* NGSPICE file created from diff_pair_sample_1411.ext - technology: sky130A

.subckt diff_pair_sample_1411 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VP.t0 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X1 VDD2.t9 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X2 VTAIL.t16 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X3 VDD2.t8 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X4 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=0 ps=0 w=11.55 l=3.39
X5 VTAIL.t19 VN.t2 VDD2.t7 B.t23 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=0 ps=0 w=11.55 l=3.39
X7 VDD1.t1 VP.t2 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X8 VTAIL.t18 VN.t3 VDD2.t6 B.t22 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X9 VTAIL.t0 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X10 VDD1.t0 VP.t3 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=4.5045 ps=23.88 w=11.55 l=3.39
X11 VDD1.t7 VP.t4 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X12 VDD2.t4 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X13 VDD2.t3 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=4.5045 ps=23.88 w=11.55 l=3.39
X14 VDD1.t6 VP.t5 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=4.5045 ps=23.88 w=11.55 l=3.39
X15 VDD1.t9 VP.t6 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X16 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=0 ps=0 w=11.55 l=3.39
X17 VTAIL.t4 VN.t7 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X18 VTAIL.t10 VP.t7 VDD1.t8 B.t23 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5045 pd=23.88 as=0 ps=0 w=11.55 l=3.39
X20 VDD1.t3 VP.t8 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X21 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
X22 VDD2.t0 VN.t9 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=4.5045 ps=23.88 w=11.55 l=3.39
X23 VTAIL.t8 VP.t9 VDD1.t2 B.t22 sky130_fd_pr__nfet_01v8 ad=1.90575 pd=11.88 as=1.90575 ps=11.88 w=11.55 l=3.39
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n21 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n57 VP.n20 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n19 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n18 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n115 VP.n114 161.3
R23 VP.n113 VP.n1 161.3
R24 VP.n112 VP.n111 161.3
R25 VP.n110 VP.n2 161.3
R26 VP.n109 VP.n108 161.3
R27 VP.n107 VP.n3 161.3
R28 VP.n106 VP.n105 161.3
R29 VP.n104 VP.n4 161.3
R30 VP.n103 VP.n102 161.3
R31 VP.n100 VP.n5 161.3
R32 VP.n99 VP.n98 161.3
R33 VP.n97 VP.n6 161.3
R34 VP.n96 VP.n95 161.3
R35 VP.n94 VP.n7 161.3
R36 VP.n93 VP.n92 161.3
R37 VP.n91 VP.n90 161.3
R38 VP.n89 VP.n9 161.3
R39 VP.n88 VP.n87 161.3
R40 VP.n86 VP.n10 161.3
R41 VP.n85 VP.n84 161.3
R42 VP.n83 VP.n11 161.3
R43 VP.n82 VP.n81 161.3
R44 VP.n80 VP.n79 161.3
R45 VP.n78 VP.n13 161.3
R46 VP.n77 VP.n76 161.3
R47 VP.n75 VP.n14 161.3
R48 VP.n74 VP.n73 161.3
R49 VP.n72 VP.n15 161.3
R50 VP.n71 VP.n70 161.3
R51 VP.n69 VP.n16 161.3
R52 VP.n30 VP.t4 115.392
R53 VP.n67 VP.t2 82.1111
R54 VP.n12 VP.t9 82.1111
R55 VP.n8 VP.t8 82.1111
R56 VP.n101 VP.t7 82.1111
R57 VP.n0 VP.t5 82.1111
R58 VP.n17 VP.t3 82.1111
R59 VP.n51 VP.t0 82.1111
R60 VP.n25 VP.t6 82.1111
R61 VP.n29 VP.t1 82.1111
R62 VP.n68 VP.n67 80.7699
R63 VP.n116 VP.n0 80.7699
R64 VP.n66 VP.n17 80.7699
R65 VP.n68 VP.n66 57.1205
R66 VP.n73 VP.n14 56.5193
R67 VP.n108 VP.n2 56.5193
R68 VP.n58 VP.n19 56.5193
R69 VP.n30 VP.n29 51.5827
R70 VP.n84 VP.n10 51.1773
R71 VP.n99 VP.n6 51.1773
R72 VP.n49 VP.n23 51.1773
R73 VP.n34 VP.n27 51.1773
R74 VP.n88 VP.n10 29.8095
R75 VP.n95 VP.n6 29.8095
R76 VP.n45 VP.n23 29.8095
R77 VP.n38 VP.n27 29.8095
R78 VP.n71 VP.n16 24.4675
R79 VP.n72 VP.n71 24.4675
R80 VP.n73 VP.n72 24.4675
R81 VP.n77 VP.n14 24.4675
R82 VP.n78 VP.n77 24.4675
R83 VP.n79 VP.n78 24.4675
R84 VP.n83 VP.n82 24.4675
R85 VP.n84 VP.n83 24.4675
R86 VP.n89 VP.n88 24.4675
R87 VP.n90 VP.n89 24.4675
R88 VP.n94 VP.n93 24.4675
R89 VP.n95 VP.n94 24.4675
R90 VP.n100 VP.n99 24.4675
R91 VP.n102 VP.n100 24.4675
R92 VP.n106 VP.n4 24.4675
R93 VP.n107 VP.n106 24.4675
R94 VP.n108 VP.n107 24.4675
R95 VP.n112 VP.n2 24.4675
R96 VP.n113 VP.n112 24.4675
R97 VP.n114 VP.n113 24.4675
R98 VP.n62 VP.n19 24.4675
R99 VP.n63 VP.n62 24.4675
R100 VP.n64 VP.n63 24.4675
R101 VP.n50 VP.n49 24.4675
R102 VP.n52 VP.n50 24.4675
R103 VP.n56 VP.n21 24.4675
R104 VP.n57 VP.n56 24.4675
R105 VP.n58 VP.n57 24.4675
R106 VP.n39 VP.n38 24.4675
R107 VP.n40 VP.n39 24.4675
R108 VP.n44 VP.n43 24.4675
R109 VP.n45 VP.n44 24.4675
R110 VP.n33 VP.n32 24.4675
R111 VP.n34 VP.n33 24.4675
R112 VP.n82 VP.n12 22.9995
R113 VP.n102 VP.n101 22.9995
R114 VP.n52 VP.n51 22.9995
R115 VP.n32 VP.n29 22.9995
R116 VP.n90 VP.n8 12.234
R117 VP.n93 VP.n8 12.234
R118 VP.n40 VP.n25 12.234
R119 VP.n43 VP.n25 12.234
R120 VP.n67 VP.n16 9.29796
R121 VP.n114 VP.n0 9.29796
R122 VP.n64 VP.n17 9.29796
R123 VP.n31 VP.n30 3.17991
R124 VP.n79 VP.n12 1.46852
R125 VP.n101 VP.n4 1.46852
R126 VP.n51 VP.n21 1.46852
R127 VP.n66 VP.n65 0.354971
R128 VP.n69 VP.n68 0.354971
R129 VP.n116 VP.n115 0.354971
R130 VP VP.n116 0.26696
R131 VP.n31 VP.n28 0.189894
R132 VP.n35 VP.n28 0.189894
R133 VP.n36 VP.n35 0.189894
R134 VP.n37 VP.n36 0.189894
R135 VP.n37 VP.n26 0.189894
R136 VP.n41 VP.n26 0.189894
R137 VP.n42 VP.n41 0.189894
R138 VP.n42 VP.n24 0.189894
R139 VP.n46 VP.n24 0.189894
R140 VP.n47 VP.n46 0.189894
R141 VP.n48 VP.n47 0.189894
R142 VP.n48 VP.n22 0.189894
R143 VP.n53 VP.n22 0.189894
R144 VP.n54 VP.n53 0.189894
R145 VP.n55 VP.n54 0.189894
R146 VP.n55 VP.n20 0.189894
R147 VP.n59 VP.n20 0.189894
R148 VP.n60 VP.n59 0.189894
R149 VP.n61 VP.n60 0.189894
R150 VP.n61 VP.n18 0.189894
R151 VP.n65 VP.n18 0.189894
R152 VP.n70 VP.n69 0.189894
R153 VP.n70 VP.n15 0.189894
R154 VP.n74 VP.n15 0.189894
R155 VP.n75 VP.n74 0.189894
R156 VP.n76 VP.n75 0.189894
R157 VP.n76 VP.n13 0.189894
R158 VP.n80 VP.n13 0.189894
R159 VP.n81 VP.n80 0.189894
R160 VP.n81 VP.n11 0.189894
R161 VP.n85 VP.n11 0.189894
R162 VP.n86 VP.n85 0.189894
R163 VP.n87 VP.n86 0.189894
R164 VP.n87 VP.n9 0.189894
R165 VP.n91 VP.n9 0.189894
R166 VP.n92 VP.n91 0.189894
R167 VP.n92 VP.n7 0.189894
R168 VP.n96 VP.n7 0.189894
R169 VP.n97 VP.n96 0.189894
R170 VP.n98 VP.n97 0.189894
R171 VP.n98 VP.n5 0.189894
R172 VP.n103 VP.n5 0.189894
R173 VP.n104 VP.n103 0.189894
R174 VP.n105 VP.n104 0.189894
R175 VP.n105 VP.n3 0.189894
R176 VP.n109 VP.n3 0.189894
R177 VP.n110 VP.n109 0.189894
R178 VP.n111 VP.n110 0.189894
R179 VP.n111 VP.n1 0.189894
R180 VP.n115 VP.n1 0.189894
R181 VDD1.n56 VDD1.n0 289.615
R182 VDD1.n119 VDD1.n63 289.615
R183 VDD1.n57 VDD1.n56 185
R184 VDD1.n55 VDD1.n54 185
R185 VDD1.n4 VDD1.n3 185
R186 VDD1.n49 VDD1.n48 185
R187 VDD1.n47 VDD1.n46 185
R188 VDD1.n8 VDD1.n7 185
R189 VDD1.n12 VDD1.n10 185
R190 VDD1.n41 VDD1.n40 185
R191 VDD1.n39 VDD1.n38 185
R192 VDD1.n14 VDD1.n13 185
R193 VDD1.n33 VDD1.n32 185
R194 VDD1.n31 VDD1.n30 185
R195 VDD1.n18 VDD1.n17 185
R196 VDD1.n25 VDD1.n24 185
R197 VDD1.n23 VDD1.n22 185
R198 VDD1.n84 VDD1.n83 185
R199 VDD1.n86 VDD1.n85 185
R200 VDD1.n79 VDD1.n78 185
R201 VDD1.n92 VDD1.n91 185
R202 VDD1.n94 VDD1.n93 185
R203 VDD1.n75 VDD1.n74 185
R204 VDD1.n101 VDD1.n100 185
R205 VDD1.n102 VDD1.n73 185
R206 VDD1.n104 VDD1.n103 185
R207 VDD1.n71 VDD1.n70 185
R208 VDD1.n110 VDD1.n109 185
R209 VDD1.n112 VDD1.n111 185
R210 VDD1.n67 VDD1.n66 185
R211 VDD1.n118 VDD1.n117 185
R212 VDD1.n120 VDD1.n119 185
R213 VDD1.n21 VDD1.t7 149.524
R214 VDD1.n82 VDD1.t1 149.524
R215 VDD1.n56 VDD1.n55 104.615
R216 VDD1.n55 VDD1.n3 104.615
R217 VDD1.n48 VDD1.n3 104.615
R218 VDD1.n48 VDD1.n47 104.615
R219 VDD1.n47 VDD1.n7 104.615
R220 VDD1.n12 VDD1.n7 104.615
R221 VDD1.n40 VDD1.n12 104.615
R222 VDD1.n40 VDD1.n39 104.615
R223 VDD1.n39 VDD1.n13 104.615
R224 VDD1.n32 VDD1.n13 104.615
R225 VDD1.n32 VDD1.n31 104.615
R226 VDD1.n31 VDD1.n17 104.615
R227 VDD1.n24 VDD1.n17 104.615
R228 VDD1.n24 VDD1.n23 104.615
R229 VDD1.n85 VDD1.n84 104.615
R230 VDD1.n85 VDD1.n78 104.615
R231 VDD1.n92 VDD1.n78 104.615
R232 VDD1.n93 VDD1.n92 104.615
R233 VDD1.n93 VDD1.n74 104.615
R234 VDD1.n101 VDD1.n74 104.615
R235 VDD1.n102 VDD1.n101 104.615
R236 VDD1.n103 VDD1.n102 104.615
R237 VDD1.n103 VDD1.n70 104.615
R238 VDD1.n110 VDD1.n70 104.615
R239 VDD1.n111 VDD1.n110 104.615
R240 VDD1.n111 VDD1.n66 104.615
R241 VDD1.n118 VDD1.n66 104.615
R242 VDD1.n119 VDD1.n118 104.615
R243 VDD1.n127 VDD1.n126 67.3487
R244 VDD1.n62 VDD1.n61 64.999
R245 VDD1.n129 VDD1.n128 64.9988
R246 VDD1.n125 VDD1.n124 64.9988
R247 VDD1.n62 VDD1.n60 54.9801
R248 VDD1.n125 VDD1.n123 54.9801
R249 VDD1.n23 VDD1.t7 52.3082
R250 VDD1.n84 VDD1.t1 52.3082
R251 VDD1.n129 VDD1.n127 51.0914
R252 VDD1.n10 VDD1.n8 13.1884
R253 VDD1.n104 VDD1.n71 13.1884
R254 VDD1.n46 VDD1.n45 12.8005
R255 VDD1.n42 VDD1.n41 12.8005
R256 VDD1.n105 VDD1.n73 12.8005
R257 VDD1.n109 VDD1.n108 12.8005
R258 VDD1.n49 VDD1.n6 12.0247
R259 VDD1.n38 VDD1.n11 12.0247
R260 VDD1.n100 VDD1.n99 12.0247
R261 VDD1.n112 VDD1.n69 12.0247
R262 VDD1.n50 VDD1.n4 11.249
R263 VDD1.n37 VDD1.n14 11.249
R264 VDD1.n98 VDD1.n75 11.249
R265 VDD1.n113 VDD1.n67 11.249
R266 VDD1.n54 VDD1.n53 10.4732
R267 VDD1.n34 VDD1.n33 10.4732
R268 VDD1.n95 VDD1.n94 10.4732
R269 VDD1.n117 VDD1.n116 10.4732
R270 VDD1.n22 VDD1.n21 10.2747
R271 VDD1.n83 VDD1.n82 10.2747
R272 VDD1.n57 VDD1.n2 9.69747
R273 VDD1.n30 VDD1.n16 9.69747
R274 VDD1.n91 VDD1.n77 9.69747
R275 VDD1.n120 VDD1.n65 9.69747
R276 VDD1.n60 VDD1.n59 9.45567
R277 VDD1.n123 VDD1.n122 9.45567
R278 VDD1.n20 VDD1.n19 9.3005
R279 VDD1.n27 VDD1.n26 9.3005
R280 VDD1.n29 VDD1.n28 9.3005
R281 VDD1.n16 VDD1.n15 9.3005
R282 VDD1.n35 VDD1.n34 9.3005
R283 VDD1.n37 VDD1.n36 9.3005
R284 VDD1.n11 VDD1.n9 9.3005
R285 VDD1.n43 VDD1.n42 9.3005
R286 VDD1.n59 VDD1.n58 9.3005
R287 VDD1.n2 VDD1.n1 9.3005
R288 VDD1.n53 VDD1.n52 9.3005
R289 VDD1.n51 VDD1.n50 9.3005
R290 VDD1.n6 VDD1.n5 9.3005
R291 VDD1.n45 VDD1.n44 9.3005
R292 VDD1.n122 VDD1.n121 9.3005
R293 VDD1.n65 VDD1.n64 9.3005
R294 VDD1.n116 VDD1.n115 9.3005
R295 VDD1.n114 VDD1.n113 9.3005
R296 VDD1.n69 VDD1.n68 9.3005
R297 VDD1.n108 VDD1.n107 9.3005
R298 VDD1.n81 VDD1.n80 9.3005
R299 VDD1.n88 VDD1.n87 9.3005
R300 VDD1.n90 VDD1.n89 9.3005
R301 VDD1.n77 VDD1.n76 9.3005
R302 VDD1.n96 VDD1.n95 9.3005
R303 VDD1.n98 VDD1.n97 9.3005
R304 VDD1.n99 VDD1.n72 9.3005
R305 VDD1.n106 VDD1.n105 9.3005
R306 VDD1.n58 VDD1.n0 8.92171
R307 VDD1.n29 VDD1.n18 8.92171
R308 VDD1.n90 VDD1.n79 8.92171
R309 VDD1.n121 VDD1.n63 8.92171
R310 VDD1.n26 VDD1.n25 8.14595
R311 VDD1.n87 VDD1.n86 8.14595
R312 VDD1.n22 VDD1.n20 7.3702
R313 VDD1.n83 VDD1.n81 7.3702
R314 VDD1.n25 VDD1.n20 5.81868
R315 VDD1.n86 VDD1.n81 5.81868
R316 VDD1.n60 VDD1.n0 5.04292
R317 VDD1.n26 VDD1.n18 5.04292
R318 VDD1.n87 VDD1.n79 5.04292
R319 VDD1.n123 VDD1.n63 5.04292
R320 VDD1.n58 VDD1.n57 4.26717
R321 VDD1.n30 VDD1.n29 4.26717
R322 VDD1.n91 VDD1.n90 4.26717
R323 VDD1.n121 VDD1.n120 4.26717
R324 VDD1.n54 VDD1.n2 3.49141
R325 VDD1.n33 VDD1.n16 3.49141
R326 VDD1.n94 VDD1.n77 3.49141
R327 VDD1.n117 VDD1.n65 3.49141
R328 VDD1.n21 VDD1.n19 2.84303
R329 VDD1.n82 VDD1.n80 2.84303
R330 VDD1.n53 VDD1.n4 2.71565
R331 VDD1.n34 VDD1.n14 2.71565
R332 VDD1.n95 VDD1.n75 2.71565
R333 VDD1.n116 VDD1.n67 2.71565
R334 VDD1 VDD1.n129 2.34748
R335 VDD1.n50 VDD1.n49 1.93989
R336 VDD1.n38 VDD1.n37 1.93989
R337 VDD1.n100 VDD1.n98 1.93989
R338 VDD1.n113 VDD1.n112 1.93989
R339 VDD1.n128 VDD1.t5 1.71479
R340 VDD1.n128 VDD1.t0 1.71479
R341 VDD1.n61 VDD1.t4 1.71479
R342 VDD1.n61 VDD1.t9 1.71479
R343 VDD1.n126 VDD1.t8 1.71479
R344 VDD1.n126 VDD1.t6 1.71479
R345 VDD1.n124 VDD1.t2 1.71479
R346 VDD1.n124 VDD1.t3 1.71479
R347 VDD1.n46 VDD1.n6 1.16414
R348 VDD1.n41 VDD1.n11 1.16414
R349 VDD1.n99 VDD1.n73 1.16414
R350 VDD1.n109 VDD1.n69 1.16414
R351 VDD1 VDD1.n62 0.860414
R352 VDD1.n127 VDD1.n125 0.746878
R353 VDD1.n45 VDD1.n8 0.388379
R354 VDD1.n42 VDD1.n10 0.388379
R355 VDD1.n105 VDD1.n104 0.388379
R356 VDD1.n108 VDD1.n71 0.388379
R357 VDD1.n59 VDD1.n1 0.155672
R358 VDD1.n52 VDD1.n1 0.155672
R359 VDD1.n52 VDD1.n51 0.155672
R360 VDD1.n51 VDD1.n5 0.155672
R361 VDD1.n44 VDD1.n5 0.155672
R362 VDD1.n44 VDD1.n43 0.155672
R363 VDD1.n43 VDD1.n9 0.155672
R364 VDD1.n36 VDD1.n9 0.155672
R365 VDD1.n36 VDD1.n35 0.155672
R366 VDD1.n35 VDD1.n15 0.155672
R367 VDD1.n28 VDD1.n15 0.155672
R368 VDD1.n28 VDD1.n27 0.155672
R369 VDD1.n27 VDD1.n19 0.155672
R370 VDD1.n88 VDD1.n80 0.155672
R371 VDD1.n89 VDD1.n88 0.155672
R372 VDD1.n89 VDD1.n76 0.155672
R373 VDD1.n96 VDD1.n76 0.155672
R374 VDD1.n97 VDD1.n96 0.155672
R375 VDD1.n97 VDD1.n72 0.155672
R376 VDD1.n106 VDD1.n72 0.155672
R377 VDD1.n107 VDD1.n106 0.155672
R378 VDD1.n107 VDD1.n68 0.155672
R379 VDD1.n114 VDD1.n68 0.155672
R380 VDD1.n115 VDD1.n114 0.155672
R381 VDD1.n115 VDD1.n64 0.155672
R382 VDD1.n122 VDD1.n64 0.155672
R383 VTAIL.n256 VTAIL.n200 289.615
R384 VTAIL.n58 VTAIL.n2 289.615
R385 VTAIL.n194 VTAIL.n138 289.615
R386 VTAIL.n128 VTAIL.n72 289.615
R387 VTAIL.n221 VTAIL.n220 185
R388 VTAIL.n223 VTAIL.n222 185
R389 VTAIL.n216 VTAIL.n215 185
R390 VTAIL.n229 VTAIL.n228 185
R391 VTAIL.n231 VTAIL.n230 185
R392 VTAIL.n212 VTAIL.n211 185
R393 VTAIL.n238 VTAIL.n237 185
R394 VTAIL.n239 VTAIL.n210 185
R395 VTAIL.n241 VTAIL.n240 185
R396 VTAIL.n208 VTAIL.n207 185
R397 VTAIL.n247 VTAIL.n246 185
R398 VTAIL.n249 VTAIL.n248 185
R399 VTAIL.n204 VTAIL.n203 185
R400 VTAIL.n255 VTAIL.n254 185
R401 VTAIL.n257 VTAIL.n256 185
R402 VTAIL.n23 VTAIL.n22 185
R403 VTAIL.n25 VTAIL.n24 185
R404 VTAIL.n18 VTAIL.n17 185
R405 VTAIL.n31 VTAIL.n30 185
R406 VTAIL.n33 VTAIL.n32 185
R407 VTAIL.n14 VTAIL.n13 185
R408 VTAIL.n40 VTAIL.n39 185
R409 VTAIL.n41 VTAIL.n12 185
R410 VTAIL.n43 VTAIL.n42 185
R411 VTAIL.n10 VTAIL.n9 185
R412 VTAIL.n49 VTAIL.n48 185
R413 VTAIL.n51 VTAIL.n50 185
R414 VTAIL.n6 VTAIL.n5 185
R415 VTAIL.n57 VTAIL.n56 185
R416 VTAIL.n59 VTAIL.n58 185
R417 VTAIL.n195 VTAIL.n194 185
R418 VTAIL.n193 VTAIL.n192 185
R419 VTAIL.n142 VTAIL.n141 185
R420 VTAIL.n187 VTAIL.n186 185
R421 VTAIL.n185 VTAIL.n184 185
R422 VTAIL.n146 VTAIL.n145 185
R423 VTAIL.n150 VTAIL.n148 185
R424 VTAIL.n179 VTAIL.n178 185
R425 VTAIL.n177 VTAIL.n176 185
R426 VTAIL.n152 VTAIL.n151 185
R427 VTAIL.n171 VTAIL.n170 185
R428 VTAIL.n169 VTAIL.n168 185
R429 VTAIL.n156 VTAIL.n155 185
R430 VTAIL.n163 VTAIL.n162 185
R431 VTAIL.n161 VTAIL.n160 185
R432 VTAIL.n129 VTAIL.n128 185
R433 VTAIL.n127 VTAIL.n126 185
R434 VTAIL.n76 VTAIL.n75 185
R435 VTAIL.n121 VTAIL.n120 185
R436 VTAIL.n119 VTAIL.n118 185
R437 VTAIL.n80 VTAIL.n79 185
R438 VTAIL.n84 VTAIL.n82 185
R439 VTAIL.n113 VTAIL.n112 185
R440 VTAIL.n111 VTAIL.n110 185
R441 VTAIL.n86 VTAIL.n85 185
R442 VTAIL.n105 VTAIL.n104 185
R443 VTAIL.n103 VTAIL.n102 185
R444 VTAIL.n90 VTAIL.n89 185
R445 VTAIL.n97 VTAIL.n96 185
R446 VTAIL.n95 VTAIL.n94 185
R447 VTAIL.n219 VTAIL.t3 149.524
R448 VTAIL.n21 VTAIL.t12 149.524
R449 VTAIL.n159 VTAIL.t14 149.524
R450 VTAIL.n93 VTAIL.t5 149.524
R451 VTAIL.n222 VTAIL.n221 104.615
R452 VTAIL.n222 VTAIL.n215 104.615
R453 VTAIL.n229 VTAIL.n215 104.615
R454 VTAIL.n230 VTAIL.n229 104.615
R455 VTAIL.n230 VTAIL.n211 104.615
R456 VTAIL.n238 VTAIL.n211 104.615
R457 VTAIL.n239 VTAIL.n238 104.615
R458 VTAIL.n240 VTAIL.n239 104.615
R459 VTAIL.n240 VTAIL.n207 104.615
R460 VTAIL.n247 VTAIL.n207 104.615
R461 VTAIL.n248 VTAIL.n247 104.615
R462 VTAIL.n248 VTAIL.n203 104.615
R463 VTAIL.n255 VTAIL.n203 104.615
R464 VTAIL.n256 VTAIL.n255 104.615
R465 VTAIL.n24 VTAIL.n23 104.615
R466 VTAIL.n24 VTAIL.n17 104.615
R467 VTAIL.n31 VTAIL.n17 104.615
R468 VTAIL.n32 VTAIL.n31 104.615
R469 VTAIL.n32 VTAIL.n13 104.615
R470 VTAIL.n40 VTAIL.n13 104.615
R471 VTAIL.n41 VTAIL.n40 104.615
R472 VTAIL.n42 VTAIL.n41 104.615
R473 VTAIL.n42 VTAIL.n9 104.615
R474 VTAIL.n49 VTAIL.n9 104.615
R475 VTAIL.n50 VTAIL.n49 104.615
R476 VTAIL.n50 VTAIL.n5 104.615
R477 VTAIL.n57 VTAIL.n5 104.615
R478 VTAIL.n58 VTAIL.n57 104.615
R479 VTAIL.n194 VTAIL.n193 104.615
R480 VTAIL.n193 VTAIL.n141 104.615
R481 VTAIL.n186 VTAIL.n141 104.615
R482 VTAIL.n186 VTAIL.n185 104.615
R483 VTAIL.n185 VTAIL.n145 104.615
R484 VTAIL.n150 VTAIL.n145 104.615
R485 VTAIL.n178 VTAIL.n150 104.615
R486 VTAIL.n178 VTAIL.n177 104.615
R487 VTAIL.n177 VTAIL.n151 104.615
R488 VTAIL.n170 VTAIL.n151 104.615
R489 VTAIL.n170 VTAIL.n169 104.615
R490 VTAIL.n169 VTAIL.n155 104.615
R491 VTAIL.n162 VTAIL.n155 104.615
R492 VTAIL.n162 VTAIL.n161 104.615
R493 VTAIL.n128 VTAIL.n127 104.615
R494 VTAIL.n127 VTAIL.n75 104.615
R495 VTAIL.n120 VTAIL.n75 104.615
R496 VTAIL.n120 VTAIL.n119 104.615
R497 VTAIL.n119 VTAIL.n79 104.615
R498 VTAIL.n84 VTAIL.n79 104.615
R499 VTAIL.n112 VTAIL.n84 104.615
R500 VTAIL.n112 VTAIL.n111 104.615
R501 VTAIL.n111 VTAIL.n85 104.615
R502 VTAIL.n104 VTAIL.n85 104.615
R503 VTAIL.n104 VTAIL.n103 104.615
R504 VTAIL.n103 VTAIL.n89 104.615
R505 VTAIL.n96 VTAIL.n89 104.615
R506 VTAIL.n96 VTAIL.n95 104.615
R507 VTAIL.n221 VTAIL.t3 52.3082
R508 VTAIL.n23 VTAIL.t12 52.3082
R509 VTAIL.n161 VTAIL.t14 52.3082
R510 VTAIL.n95 VTAIL.t5 52.3082
R511 VTAIL.n137 VTAIL.n136 48.3202
R512 VTAIL.n135 VTAIL.n134 48.3202
R513 VTAIL.n71 VTAIL.n70 48.3202
R514 VTAIL.n69 VTAIL.n68 48.3202
R515 VTAIL.n263 VTAIL.n262 48.32
R516 VTAIL.n1 VTAIL.n0 48.32
R517 VTAIL.n65 VTAIL.n64 48.32
R518 VTAIL.n67 VTAIL.n66 48.32
R519 VTAIL.n261 VTAIL.n260 35.0944
R520 VTAIL.n63 VTAIL.n62 35.0944
R521 VTAIL.n199 VTAIL.n198 35.0944
R522 VTAIL.n133 VTAIL.n132 35.0944
R523 VTAIL.n69 VTAIL.n67 28.7376
R524 VTAIL.n261 VTAIL.n199 25.5307
R525 VTAIL.n241 VTAIL.n208 13.1884
R526 VTAIL.n43 VTAIL.n10 13.1884
R527 VTAIL.n148 VTAIL.n146 13.1884
R528 VTAIL.n82 VTAIL.n80 13.1884
R529 VTAIL.n242 VTAIL.n210 12.8005
R530 VTAIL.n246 VTAIL.n245 12.8005
R531 VTAIL.n44 VTAIL.n12 12.8005
R532 VTAIL.n48 VTAIL.n47 12.8005
R533 VTAIL.n184 VTAIL.n183 12.8005
R534 VTAIL.n180 VTAIL.n179 12.8005
R535 VTAIL.n118 VTAIL.n117 12.8005
R536 VTAIL.n114 VTAIL.n113 12.8005
R537 VTAIL.n237 VTAIL.n236 12.0247
R538 VTAIL.n249 VTAIL.n206 12.0247
R539 VTAIL.n39 VTAIL.n38 12.0247
R540 VTAIL.n51 VTAIL.n8 12.0247
R541 VTAIL.n187 VTAIL.n144 12.0247
R542 VTAIL.n176 VTAIL.n149 12.0247
R543 VTAIL.n121 VTAIL.n78 12.0247
R544 VTAIL.n110 VTAIL.n83 12.0247
R545 VTAIL.n235 VTAIL.n212 11.249
R546 VTAIL.n250 VTAIL.n204 11.249
R547 VTAIL.n37 VTAIL.n14 11.249
R548 VTAIL.n52 VTAIL.n6 11.249
R549 VTAIL.n188 VTAIL.n142 11.249
R550 VTAIL.n175 VTAIL.n152 11.249
R551 VTAIL.n122 VTAIL.n76 11.249
R552 VTAIL.n109 VTAIL.n86 11.249
R553 VTAIL.n232 VTAIL.n231 10.4732
R554 VTAIL.n254 VTAIL.n253 10.4732
R555 VTAIL.n34 VTAIL.n33 10.4732
R556 VTAIL.n56 VTAIL.n55 10.4732
R557 VTAIL.n192 VTAIL.n191 10.4732
R558 VTAIL.n172 VTAIL.n171 10.4732
R559 VTAIL.n126 VTAIL.n125 10.4732
R560 VTAIL.n106 VTAIL.n105 10.4732
R561 VTAIL.n220 VTAIL.n219 10.2747
R562 VTAIL.n22 VTAIL.n21 10.2747
R563 VTAIL.n160 VTAIL.n159 10.2747
R564 VTAIL.n94 VTAIL.n93 10.2747
R565 VTAIL.n228 VTAIL.n214 9.69747
R566 VTAIL.n257 VTAIL.n202 9.69747
R567 VTAIL.n30 VTAIL.n16 9.69747
R568 VTAIL.n59 VTAIL.n4 9.69747
R569 VTAIL.n195 VTAIL.n140 9.69747
R570 VTAIL.n168 VTAIL.n154 9.69747
R571 VTAIL.n129 VTAIL.n74 9.69747
R572 VTAIL.n102 VTAIL.n88 9.69747
R573 VTAIL.n260 VTAIL.n259 9.45567
R574 VTAIL.n62 VTAIL.n61 9.45567
R575 VTAIL.n198 VTAIL.n197 9.45567
R576 VTAIL.n132 VTAIL.n131 9.45567
R577 VTAIL.n259 VTAIL.n258 9.3005
R578 VTAIL.n202 VTAIL.n201 9.3005
R579 VTAIL.n253 VTAIL.n252 9.3005
R580 VTAIL.n251 VTAIL.n250 9.3005
R581 VTAIL.n206 VTAIL.n205 9.3005
R582 VTAIL.n245 VTAIL.n244 9.3005
R583 VTAIL.n218 VTAIL.n217 9.3005
R584 VTAIL.n225 VTAIL.n224 9.3005
R585 VTAIL.n227 VTAIL.n226 9.3005
R586 VTAIL.n214 VTAIL.n213 9.3005
R587 VTAIL.n233 VTAIL.n232 9.3005
R588 VTAIL.n235 VTAIL.n234 9.3005
R589 VTAIL.n236 VTAIL.n209 9.3005
R590 VTAIL.n243 VTAIL.n242 9.3005
R591 VTAIL.n61 VTAIL.n60 9.3005
R592 VTAIL.n4 VTAIL.n3 9.3005
R593 VTAIL.n55 VTAIL.n54 9.3005
R594 VTAIL.n53 VTAIL.n52 9.3005
R595 VTAIL.n8 VTAIL.n7 9.3005
R596 VTAIL.n47 VTAIL.n46 9.3005
R597 VTAIL.n20 VTAIL.n19 9.3005
R598 VTAIL.n27 VTAIL.n26 9.3005
R599 VTAIL.n29 VTAIL.n28 9.3005
R600 VTAIL.n16 VTAIL.n15 9.3005
R601 VTAIL.n35 VTAIL.n34 9.3005
R602 VTAIL.n37 VTAIL.n36 9.3005
R603 VTAIL.n38 VTAIL.n11 9.3005
R604 VTAIL.n45 VTAIL.n44 9.3005
R605 VTAIL.n158 VTAIL.n157 9.3005
R606 VTAIL.n165 VTAIL.n164 9.3005
R607 VTAIL.n167 VTAIL.n166 9.3005
R608 VTAIL.n154 VTAIL.n153 9.3005
R609 VTAIL.n173 VTAIL.n172 9.3005
R610 VTAIL.n175 VTAIL.n174 9.3005
R611 VTAIL.n149 VTAIL.n147 9.3005
R612 VTAIL.n181 VTAIL.n180 9.3005
R613 VTAIL.n197 VTAIL.n196 9.3005
R614 VTAIL.n140 VTAIL.n139 9.3005
R615 VTAIL.n191 VTAIL.n190 9.3005
R616 VTAIL.n189 VTAIL.n188 9.3005
R617 VTAIL.n144 VTAIL.n143 9.3005
R618 VTAIL.n183 VTAIL.n182 9.3005
R619 VTAIL.n92 VTAIL.n91 9.3005
R620 VTAIL.n99 VTAIL.n98 9.3005
R621 VTAIL.n101 VTAIL.n100 9.3005
R622 VTAIL.n88 VTAIL.n87 9.3005
R623 VTAIL.n107 VTAIL.n106 9.3005
R624 VTAIL.n109 VTAIL.n108 9.3005
R625 VTAIL.n83 VTAIL.n81 9.3005
R626 VTAIL.n115 VTAIL.n114 9.3005
R627 VTAIL.n131 VTAIL.n130 9.3005
R628 VTAIL.n74 VTAIL.n73 9.3005
R629 VTAIL.n125 VTAIL.n124 9.3005
R630 VTAIL.n123 VTAIL.n122 9.3005
R631 VTAIL.n78 VTAIL.n77 9.3005
R632 VTAIL.n117 VTAIL.n116 9.3005
R633 VTAIL.n227 VTAIL.n216 8.92171
R634 VTAIL.n258 VTAIL.n200 8.92171
R635 VTAIL.n29 VTAIL.n18 8.92171
R636 VTAIL.n60 VTAIL.n2 8.92171
R637 VTAIL.n196 VTAIL.n138 8.92171
R638 VTAIL.n167 VTAIL.n156 8.92171
R639 VTAIL.n130 VTAIL.n72 8.92171
R640 VTAIL.n101 VTAIL.n90 8.92171
R641 VTAIL.n224 VTAIL.n223 8.14595
R642 VTAIL.n26 VTAIL.n25 8.14595
R643 VTAIL.n164 VTAIL.n163 8.14595
R644 VTAIL.n98 VTAIL.n97 8.14595
R645 VTAIL.n220 VTAIL.n218 7.3702
R646 VTAIL.n22 VTAIL.n20 7.3702
R647 VTAIL.n160 VTAIL.n158 7.3702
R648 VTAIL.n94 VTAIL.n92 7.3702
R649 VTAIL.n223 VTAIL.n218 5.81868
R650 VTAIL.n25 VTAIL.n20 5.81868
R651 VTAIL.n163 VTAIL.n158 5.81868
R652 VTAIL.n97 VTAIL.n92 5.81868
R653 VTAIL.n224 VTAIL.n216 5.04292
R654 VTAIL.n260 VTAIL.n200 5.04292
R655 VTAIL.n26 VTAIL.n18 5.04292
R656 VTAIL.n62 VTAIL.n2 5.04292
R657 VTAIL.n198 VTAIL.n138 5.04292
R658 VTAIL.n164 VTAIL.n156 5.04292
R659 VTAIL.n132 VTAIL.n72 5.04292
R660 VTAIL.n98 VTAIL.n90 5.04292
R661 VTAIL.n228 VTAIL.n227 4.26717
R662 VTAIL.n258 VTAIL.n257 4.26717
R663 VTAIL.n30 VTAIL.n29 4.26717
R664 VTAIL.n60 VTAIL.n59 4.26717
R665 VTAIL.n196 VTAIL.n195 4.26717
R666 VTAIL.n168 VTAIL.n167 4.26717
R667 VTAIL.n130 VTAIL.n129 4.26717
R668 VTAIL.n102 VTAIL.n101 4.26717
R669 VTAIL.n231 VTAIL.n214 3.49141
R670 VTAIL.n254 VTAIL.n202 3.49141
R671 VTAIL.n33 VTAIL.n16 3.49141
R672 VTAIL.n56 VTAIL.n4 3.49141
R673 VTAIL.n192 VTAIL.n140 3.49141
R674 VTAIL.n171 VTAIL.n154 3.49141
R675 VTAIL.n126 VTAIL.n74 3.49141
R676 VTAIL.n105 VTAIL.n88 3.49141
R677 VTAIL.n71 VTAIL.n69 3.2074
R678 VTAIL.n133 VTAIL.n71 3.2074
R679 VTAIL.n137 VTAIL.n135 3.2074
R680 VTAIL.n199 VTAIL.n137 3.2074
R681 VTAIL.n67 VTAIL.n65 3.2074
R682 VTAIL.n65 VTAIL.n63 3.2074
R683 VTAIL.n263 VTAIL.n261 3.2074
R684 VTAIL.n219 VTAIL.n217 2.84303
R685 VTAIL.n21 VTAIL.n19 2.84303
R686 VTAIL.n159 VTAIL.n157 2.84303
R687 VTAIL.n93 VTAIL.n91 2.84303
R688 VTAIL.n232 VTAIL.n212 2.71565
R689 VTAIL.n253 VTAIL.n204 2.71565
R690 VTAIL.n34 VTAIL.n14 2.71565
R691 VTAIL.n55 VTAIL.n6 2.71565
R692 VTAIL.n191 VTAIL.n142 2.71565
R693 VTAIL.n172 VTAIL.n152 2.71565
R694 VTAIL.n125 VTAIL.n76 2.71565
R695 VTAIL.n106 VTAIL.n86 2.71565
R696 VTAIL VTAIL.n1 2.46386
R697 VTAIL.n135 VTAIL.n133 2.07378
R698 VTAIL.n63 VTAIL.n1 2.07378
R699 VTAIL.n237 VTAIL.n235 1.93989
R700 VTAIL.n250 VTAIL.n249 1.93989
R701 VTAIL.n39 VTAIL.n37 1.93989
R702 VTAIL.n52 VTAIL.n51 1.93989
R703 VTAIL.n188 VTAIL.n187 1.93989
R704 VTAIL.n176 VTAIL.n175 1.93989
R705 VTAIL.n122 VTAIL.n121 1.93989
R706 VTAIL.n110 VTAIL.n109 1.93989
R707 VTAIL.n262 VTAIL.t1 1.71479
R708 VTAIL.n262 VTAIL.t4 1.71479
R709 VTAIL.n0 VTAIL.t2 1.71479
R710 VTAIL.n0 VTAIL.t0 1.71479
R711 VTAIL.n64 VTAIL.t9 1.71479
R712 VTAIL.n64 VTAIL.t10 1.71479
R713 VTAIL.n66 VTAIL.t15 1.71479
R714 VTAIL.n66 VTAIL.t8 1.71479
R715 VTAIL.n136 VTAIL.t11 1.71479
R716 VTAIL.n136 VTAIL.t17 1.71479
R717 VTAIL.n134 VTAIL.t13 1.71479
R718 VTAIL.n134 VTAIL.t16 1.71479
R719 VTAIL.n70 VTAIL.t7 1.71479
R720 VTAIL.n70 VTAIL.t19 1.71479
R721 VTAIL.n68 VTAIL.t6 1.71479
R722 VTAIL.n68 VTAIL.t18 1.71479
R723 VTAIL.n236 VTAIL.n210 1.16414
R724 VTAIL.n246 VTAIL.n206 1.16414
R725 VTAIL.n38 VTAIL.n12 1.16414
R726 VTAIL.n48 VTAIL.n8 1.16414
R727 VTAIL.n184 VTAIL.n144 1.16414
R728 VTAIL.n179 VTAIL.n149 1.16414
R729 VTAIL.n118 VTAIL.n78 1.16414
R730 VTAIL.n113 VTAIL.n83 1.16414
R731 VTAIL VTAIL.n263 0.744035
R732 VTAIL.n242 VTAIL.n241 0.388379
R733 VTAIL.n245 VTAIL.n208 0.388379
R734 VTAIL.n44 VTAIL.n43 0.388379
R735 VTAIL.n47 VTAIL.n10 0.388379
R736 VTAIL.n183 VTAIL.n146 0.388379
R737 VTAIL.n180 VTAIL.n148 0.388379
R738 VTAIL.n117 VTAIL.n80 0.388379
R739 VTAIL.n114 VTAIL.n82 0.388379
R740 VTAIL.n225 VTAIL.n217 0.155672
R741 VTAIL.n226 VTAIL.n225 0.155672
R742 VTAIL.n226 VTAIL.n213 0.155672
R743 VTAIL.n233 VTAIL.n213 0.155672
R744 VTAIL.n234 VTAIL.n233 0.155672
R745 VTAIL.n234 VTAIL.n209 0.155672
R746 VTAIL.n243 VTAIL.n209 0.155672
R747 VTAIL.n244 VTAIL.n243 0.155672
R748 VTAIL.n244 VTAIL.n205 0.155672
R749 VTAIL.n251 VTAIL.n205 0.155672
R750 VTAIL.n252 VTAIL.n251 0.155672
R751 VTAIL.n252 VTAIL.n201 0.155672
R752 VTAIL.n259 VTAIL.n201 0.155672
R753 VTAIL.n27 VTAIL.n19 0.155672
R754 VTAIL.n28 VTAIL.n27 0.155672
R755 VTAIL.n28 VTAIL.n15 0.155672
R756 VTAIL.n35 VTAIL.n15 0.155672
R757 VTAIL.n36 VTAIL.n35 0.155672
R758 VTAIL.n36 VTAIL.n11 0.155672
R759 VTAIL.n45 VTAIL.n11 0.155672
R760 VTAIL.n46 VTAIL.n45 0.155672
R761 VTAIL.n46 VTAIL.n7 0.155672
R762 VTAIL.n53 VTAIL.n7 0.155672
R763 VTAIL.n54 VTAIL.n53 0.155672
R764 VTAIL.n54 VTAIL.n3 0.155672
R765 VTAIL.n61 VTAIL.n3 0.155672
R766 VTAIL.n197 VTAIL.n139 0.155672
R767 VTAIL.n190 VTAIL.n139 0.155672
R768 VTAIL.n190 VTAIL.n189 0.155672
R769 VTAIL.n189 VTAIL.n143 0.155672
R770 VTAIL.n182 VTAIL.n143 0.155672
R771 VTAIL.n182 VTAIL.n181 0.155672
R772 VTAIL.n181 VTAIL.n147 0.155672
R773 VTAIL.n174 VTAIL.n147 0.155672
R774 VTAIL.n174 VTAIL.n173 0.155672
R775 VTAIL.n173 VTAIL.n153 0.155672
R776 VTAIL.n166 VTAIL.n153 0.155672
R777 VTAIL.n166 VTAIL.n165 0.155672
R778 VTAIL.n165 VTAIL.n157 0.155672
R779 VTAIL.n131 VTAIL.n73 0.155672
R780 VTAIL.n124 VTAIL.n73 0.155672
R781 VTAIL.n124 VTAIL.n123 0.155672
R782 VTAIL.n123 VTAIL.n77 0.155672
R783 VTAIL.n116 VTAIL.n77 0.155672
R784 VTAIL.n116 VTAIL.n115 0.155672
R785 VTAIL.n115 VTAIL.n81 0.155672
R786 VTAIL.n108 VTAIL.n81 0.155672
R787 VTAIL.n108 VTAIL.n107 0.155672
R788 VTAIL.n107 VTAIL.n87 0.155672
R789 VTAIL.n100 VTAIL.n87 0.155672
R790 VTAIL.n100 VTAIL.n99 0.155672
R791 VTAIL.n99 VTAIL.n91 0.155672
R792 B.n1050 B.n1049 585
R793 B.n361 B.n178 585
R794 B.n360 B.n359 585
R795 B.n358 B.n357 585
R796 B.n356 B.n355 585
R797 B.n354 B.n353 585
R798 B.n352 B.n351 585
R799 B.n350 B.n349 585
R800 B.n348 B.n347 585
R801 B.n346 B.n345 585
R802 B.n344 B.n343 585
R803 B.n342 B.n341 585
R804 B.n340 B.n339 585
R805 B.n338 B.n337 585
R806 B.n336 B.n335 585
R807 B.n334 B.n333 585
R808 B.n332 B.n331 585
R809 B.n330 B.n329 585
R810 B.n328 B.n327 585
R811 B.n326 B.n325 585
R812 B.n324 B.n323 585
R813 B.n322 B.n321 585
R814 B.n320 B.n319 585
R815 B.n318 B.n317 585
R816 B.n316 B.n315 585
R817 B.n314 B.n313 585
R818 B.n312 B.n311 585
R819 B.n310 B.n309 585
R820 B.n308 B.n307 585
R821 B.n306 B.n305 585
R822 B.n304 B.n303 585
R823 B.n302 B.n301 585
R824 B.n300 B.n299 585
R825 B.n298 B.n297 585
R826 B.n296 B.n295 585
R827 B.n294 B.n293 585
R828 B.n292 B.n291 585
R829 B.n290 B.n289 585
R830 B.n288 B.n287 585
R831 B.n286 B.n285 585
R832 B.n284 B.n283 585
R833 B.n282 B.n281 585
R834 B.n280 B.n279 585
R835 B.n278 B.n277 585
R836 B.n276 B.n275 585
R837 B.n274 B.n273 585
R838 B.n272 B.n271 585
R839 B.n270 B.n269 585
R840 B.n268 B.n267 585
R841 B.n266 B.n265 585
R842 B.n264 B.n263 585
R843 B.n262 B.n261 585
R844 B.n260 B.n259 585
R845 B.n258 B.n257 585
R846 B.n256 B.n255 585
R847 B.n254 B.n253 585
R848 B.n252 B.n251 585
R849 B.n250 B.n249 585
R850 B.n248 B.n247 585
R851 B.n246 B.n245 585
R852 B.n244 B.n243 585
R853 B.n242 B.n241 585
R854 B.n240 B.n239 585
R855 B.n238 B.n237 585
R856 B.n236 B.n235 585
R857 B.n234 B.n233 585
R858 B.n232 B.n231 585
R859 B.n230 B.n229 585
R860 B.n228 B.n227 585
R861 B.n226 B.n225 585
R862 B.n224 B.n223 585
R863 B.n222 B.n221 585
R864 B.n220 B.n219 585
R865 B.n218 B.n217 585
R866 B.n216 B.n215 585
R867 B.n214 B.n213 585
R868 B.n212 B.n211 585
R869 B.n210 B.n209 585
R870 B.n208 B.n207 585
R871 B.n206 B.n205 585
R872 B.n204 B.n203 585
R873 B.n202 B.n201 585
R874 B.n200 B.n199 585
R875 B.n198 B.n197 585
R876 B.n196 B.n195 585
R877 B.n194 B.n193 585
R878 B.n192 B.n191 585
R879 B.n190 B.n189 585
R880 B.n188 B.n187 585
R881 B.n186 B.n185 585
R882 B.n1048 B.n133 585
R883 B.n1053 B.n133 585
R884 B.n1047 B.n132 585
R885 B.n1054 B.n132 585
R886 B.n1046 B.n1045 585
R887 B.n1045 B.n128 585
R888 B.n1044 B.n127 585
R889 B.n1060 B.n127 585
R890 B.n1043 B.n126 585
R891 B.n1061 B.n126 585
R892 B.n1042 B.n125 585
R893 B.n1062 B.n125 585
R894 B.n1041 B.n1040 585
R895 B.n1040 B.n121 585
R896 B.n1039 B.n120 585
R897 B.n1068 B.n120 585
R898 B.n1038 B.n119 585
R899 B.n1069 B.n119 585
R900 B.n1037 B.n118 585
R901 B.n1070 B.n118 585
R902 B.n1036 B.n1035 585
R903 B.n1035 B.n114 585
R904 B.n1034 B.n113 585
R905 B.n1076 B.n113 585
R906 B.n1033 B.n112 585
R907 B.n1077 B.n112 585
R908 B.n1032 B.n111 585
R909 B.n1078 B.n111 585
R910 B.n1031 B.n1030 585
R911 B.n1030 B.n107 585
R912 B.n1029 B.n106 585
R913 B.n1084 B.n106 585
R914 B.n1028 B.n105 585
R915 B.n1085 B.n105 585
R916 B.n1027 B.n104 585
R917 B.n1086 B.n104 585
R918 B.n1026 B.n1025 585
R919 B.n1025 B.n100 585
R920 B.n1024 B.n99 585
R921 B.n1092 B.n99 585
R922 B.n1023 B.n98 585
R923 B.n1093 B.n98 585
R924 B.n1022 B.n97 585
R925 B.n1094 B.n97 585
R926 B.n1021 B.n1020 585
R927 B.n1020 B.n96 585
R928 B.n1019 B.n92 585
R929 B.n1100 B.n92 585
R930 B.n1018 B.n91 585
R931 B.n1101 B.n91 585
R932 B.n1017 B.n90 585
R933 B.n1102 B.n90 585
R934 B.n1016 B.n1015 585
R935 B.n1015 B.n86 585
R936 B.n1014 B.n85 585
R937 B.n1108 B.n85 585
R938 B.n1013 B.n84 585
R939 B.n1109 B.n84 585
R940 B.n1012 B.n83 585
R941 B.n1110 B.n83 585
R942 B.n1011 B.n1010 585
R943 B.n1010 B.n79 585
R944 B.n1009 B.n78 585
R945 B.n1116 B.n78 585
R946 B.n1008 B.n77 585
R947 B.n1117 B.n77 585
R948 B.n1007 B.n76 585
R949 B.n1118 B.n76 585
R950 B.n1006 B.n1005 585
R951 B.n1005 B.n72 585
R952 B.n1004 B.n71 585
R953 B.n1124 B.n71 585
R954 B.n1003 B.n70 585
R955 B.n1125 B.n70 585
R956 B.n1002 B.n69 585
R957 B.n1126 B.n69 585
R958 B.n1001 B.n1000 585
R959 B.n1000 B.n65 585
R960 B.n999 B.n64 585
R961 B.n1132 B.n64 585
R962 B.n998 B.n63 585
R963 B.n1133 B.n63 585
R964 B.n997 B.n62 585
R965 B.n1134 B.n62 585
R966 B.n996 B.n995 585
R967 B.n995 B.n58 585
R968 B.n994 B.n57 585
R969 B.n1140 B.n57 585
R970 B.n993 B.n56 585
R971 B.n1141 B.n56 585
R972 B.n992 B.n55 585
R973 B.n1142 B.n55 585
R974 B.n991 B.n990 585
R975 B.n990 B.n51 585
R976 B.n989 B.n50 585
R977 B.n1148 B.n50 585
R978 B.n988 B.n49 585
R979 B.n1149 B.n49 585
R980 B.n987 B.n48 585
R981 B.n1150 B.n48 585
R982 B.n986 B.n985 585
R983 B.n985 B.n44 585
R984 B.n984 B.n43 585
R985 B.n1156 B.n43 585
R986 B.n983 B.n42 585
R987 B.n1157 B.n42 585
R988 B.n982 B.n41 585
R989 B.n1158 B.n41 585
R990 B.n981 B.n980 585
R991 B.n980 B.n37 585
R992 B.n979 B.n36 585
R993 B.n1164 B.n36 585
R994 B.n978 B.n35 585
R995 B.n1165 B.n35 585
R996 B.n977 B.n34 585
R997 B.n1166 B.n34 585
R998 B.n976 B.n975 585
R999 B.n975 B.n30 585
R1000 B.n974 B.n29 585
R1001 B.n1172 B.n29 585
R1002 B.n973 B.n28 585
R1003 B.n1173 B.n28 585
R1004 B.n972 B.n27 585
R1005 B.n1174 B.n27 585
R1006 B.n971 B.n970 585
R1007 B.n970 B.n23 585
R1008 B.n969 B.n22 585
R1009 B.n1180 B.n22 585
R1010 B.n968 B.n21 585
R1011 B.n1181 B.n21 585
R1012 B.n967 B.n20 585
R1013 B.n1182 B.n20 585
R1014 B.n966 B.n965 585
R1015 B.n965 B.n19 585
R1016 B.n964 B.n15 585
R1017 B.n1188 B.n15 585
R1018 B.n963 B.n14 585
R1019 B.n1189 B.n14 585
R1020 B.n962 B.n13 585
R1021 B.n1190 B.n13 585
R1022 B.n961 B.n960 585
R1023 B.n960 B.n12 585
R1024 B.n959 B.n958 585
R1025 B.n959 B.n8 585
R1026 B.n957 B.n7 585
R1027 B.n1197 B.n7 585
R1028 B.n956 B.n6 585
R1029 B.n1198 B.n6 585
R1030 B.n955 B.n5 585
R1031 B.n1199 B.n5 585
R1032 B.n954 B.n953 585
R1033 B.n953 B.n4 585
R1034 B.n952 B.n362 585
R1035 B.n952 B.n951 585
R1036 B.n942 B.n363 585
R1037 B.n364 B.n363 585
R1038 B.n944 B.n943 585
R1039 B.n945 B.n944 585
R1040 B.n941 B.n369 585
R1041 B.n369 B.n368 585
R1042 B.n940 B.n939 585
R1043 B.n939 B.n938 585
R1044 B.n371 B.n370 585
R1045 B.n931 B.n371 585
R1046 B.n930 B.n929 585
R1047 B.n932 B.n930 585
R1048 B.n928 B.n376 585
R1049 B.n376 B.n375 585
R1050 B.n927 B.n926 585
R1051 B.n926 B.n925 585
R1052 B.n378 B.n377 585
R1053 B.n379 B.n378 585
R1054 B.n918 B.n917 585
R1055 B.n919 B.n918 585
R1056 B.n916 B.n384 585
R1057 B.n384 B.n383 585
R1058 B.n915 B.n914 585
R1059 B.n914 B.n913 585
R1060 B.n386 B.n385 585
R1061 B.n387 B.n386 585
R1062 B.n906 B.n905 585
R1063 B.n907 B.n906 585
R1064 B.n904 B.n392 585
R1065 B.n392 B.n391 585
R1066 B.n903 B.n902 585
R1067 B.n902 B.n901 585
R1068 B.n394 B.n393 585
R1069 B.n395 B.n394 585
R1070 B.n894 B.n893 585
R1071 B.n895 B.n894 585
R1072 B.n892 B.n400 585
R1073 B.n400 B.n399 585
R1074 B.n891 B.n890 585
R1075 B.n890 B.n889 585
R1076 B.n402 B.n401 585
R1077 B.n403 B.n402 585
R1078 B.n882 B.n881 585
R1079 B.n883 B.n882 585
R1080 B.n880 B.n408 585
R1081 B.n408 B.n407 585
R1082 B.n879 B.n878 585
R1083 B.n878 B.n877 585
R1084 B.n410 B.n409 585
R1085 B.n411 B.n410 585
R1086 B.n870 B.n869 585
R1087 B.n871 B.n870 585
R1088 B.n868 B.n415 585
R1089 B.n419 B.n415 585
R1090 B.n867 B.n866 585
R1091 B.n866 B.n865 585
R1092 B.n417 B.n416 585
R1093 B.n418 B.n417 585
R1094 B.n858 B.n857 585
R1095 B.n859 B.n858 585
R1096 B.n856 B.n424 585
R1097 B.n424 B.n423 585
R1098 B.n855 B.n854 585
R1099 B.n854 B.n853 585
R1100 B.n426 B.n425 585
R1101 B.n427 B.n426 585
R1102 B.n846 B.n845 585
R1103 B.n847 B.n846 585
R1104 B.n844 B.n432 585
R1105 B.n432 B.n431 585
R1106 B.n843 B.n842 585
R1107 B.n842 B.n841 585
R1108 B.n434 B.n433 585
R1109 B.n435 B.n434 585
R1110 B.n834 B.n833 585
R1111 B.n835 B.n834 585
R1112 B.n832 B.n440 585
R1113 B.n440 B.n439 585
R1114 B.n831 B.n830 585
R1115 B.n830 B.n829 585
R1116 B.n442 B.n441 585
R1117 B.n443 B.n442 585
R1118 B.n822 B.n821 585
R1119 B.n823 B.n822 585
R1120 B.n820 B.n448 585
R1121 B.n448 B.n447 585
R1122 B.n819 B.n818 585
R1123 B.n818 B.n817 585
R1124 B.n450 B.n449 585
R1125 B.n451 B.n450 585
R1126 B.n810 B.n809 585
R1127 B.n811 B.n810 585
R1128 B.n808 B.n456 585
R1129 B.n456 B.n455 585
R1130 B.n807 B.n806 585
R1131 B.n806 B.n805 585
R1132 B.n458 B.n457 585
R1133 B.n798 B.n458 585
R1134 B.n797 B.n796 585
R1135 B.n799 B.n797 585
R1136 B.n795 B.n463 585
R1137 B.n463 B.n462 585
R1138 B.n794 B.n793 585
R1139 B.n793 B.n792 585
R1140 B.n465 B.n464 585
R1141 B.n466 B.n465 585
R1142 B.n785 B.n784 585
R1143 B.n786 B.n785 585
R1144 B.n783 B.n471 585
R1145 B.n471 B.n470 585
R1146 B.n782 B.n781 585
R1147 B.n781 B.n780 585
R1148 B.n473 B.n472 585
R1149 B.n474 B.n473 585
R1150 B.n773 B.n772 585
R1151 B.n774 B.n773 585
R1152 B.n771 B.n479 585
R1153 B.n479 B.n478 585
R1154 B.n770 B.n769 585
R1155 B.n769 B.n768 585
R1156 B.n481 B.n480 585
R1157 B.n482 B.n481 585
R1158 B.n761 B.n760 585
R1159 B.n762 B.n761 585
R1160 B.n759 B.n486 585
R1161 B.n490 B.n486 585
R1162 B.n758 B.n757 585
R1163 B.n757 B.n756 585
R1164 B.n488 B.n487 585
R1165 B.n489 B.n488 585
R1166 B.n749 B.n748 585
R1167 B.n750 B.n749 585
R1168 B.n747 B.n495 585
R1169 B.n495 B.n494 585
R1170 B.n746 B.n745 585
R1171 B.n745 B.n744 585
R1172 B.n497 B.n496 585
R1173 B.n498 B.n497 585
R1174 B.n737 B.n736 585
R1175 B.n738 B.n737 585
R1176 B.n735 B.n503 585
R1177 B.n503 B.n502 585
R1178 B.n730 B.n729 585
R1179 B.n728 B.n550 585
R1180 B.n727 B.n549 585
R1181 B.n732 B.n549 585
R1182 B.n726 B.n725 585
R1183 B.n724 B.n723 585
R1184 B.n722 B.n721 585
R1185 B.n720 B.n719 585
R1186 B.n718 B.n717 585
R1187 B.n716 B.n715 585
R1188 B.n714 B.n713 585
R1189 B.n712 B.n711 585
R1190 B.n710 B.n709 585
R1191 B.n708 B.n707 585
R1192 B.n706 B.n705 585
R1193 B.n704 B.n703 585
R1194 B.n702 B.n701 585
R1195 B.n700 B.n699 585
R1196 B.n698 B.n697 585
R1197 B.n696 B.n695 585
R1198 B.n694 B.n693 585
R1199 B.n692 B.n691 585
R1200 B.n690 B.n689 585
R1201 B.n688 B.n687 585
R1202 B.n686 B.n685 585
R1203 B.n684 B.n683 585
R1204 B.n682 B.n681 585
R1205 B.n680 B.n679 585
R1206 B.n678 B.n677 585
R1207 B.n676 B.n675 585
R1208 B.n674 B.n673 585
R1209 B.n672 B.n671 585
R1210 B.n670 B.n669 585
R1211 B.n668 B.n667 585
R1212 B.n666 B.n665 585
R1213 B.n664 B.n663 585
R1214 B.n662 B.n661 585
R1215 B.n660 B.n659 585
R1216 B.n658 B.n657 585
R1217 B.n656 B.n655 585
R1218 B.n654 B.n653 585
R1219 B.n651 B.n650 585
R1220 B.n649 B.n648 585
R1221 B.n647 B.n646 585
R1222 B.n645 B.n644 585
R1223 B.n643 B.n642 585
R1224 B.n641 B.n640 585
R1225 B.n639 B.n638 585
R1226 B.n637 B.n636 585
R1227 B.n635 B.n634 585
R1228 B.n633 B.n632 585
R1229 B.n630 B.n629 585
R1230 B.n628 B.n627 585
R1231 B.n626 B.n625 585
R1232 B.n624 B.n623 585
R1233 B.n622 B.n621 585
R1234 B.n620 B.n619 585
R1235 B.n618 B.n617 585
R1236 B.n616 B.n615 585
R1237 B.n614 B.n613 585
R1238 B.n612 B.n611 585
R1239 B.n610 B.n609 585
R1240 B.n608 B.n607 585
R1241 B.n606 B.n605 585
R1242 B.n604 B.n603 585
R1243 B.n602 B.n601 585
R1244 B.n600 B.n599 585
R1245 B.n598 B.n597 585
R1246 B.n596 B.n595 585
R1247 B.n594 B.n593 585
R1248 B.n592 B.n591 585
R1249 B.n590 B.n589 585
R1250 B.n588 B.n587 585
R1251 B.n586 B.n585 585
R1252 B.n584 B.n583 585
R1253 B.n582 B.n581 585
R1254 B.n580 B.n579 585
R1255 B.n578 B.n577 585
R1256 B.n576 B.n575 585
R1257 B.n574 B.n573 585
R1258 B.n572 B.n571 585
R1259 B.n570 B.n569 585
R1260 B.n568 B.n567 585
R1261 B.n566 B.n565 585
R1262 B.n564 B.n563 585
R1263 B.n562 B.n561 585
R1264 B.n560 B.n559 585
R1265 B.n558 B.n557 585
R1266 B.n556 B.n555 585
R1267 B.n505 B.n504 585
R1268 B.n734 B.n733 585
R1269 B.n733 B.n732 585
R1270 B.n501 B.n500 585
R1271 B.n502 B.n501 585
R1272 B.n740 B.n739 585
R1273 B.n739 B.n738 585
R1274 B.n741 B.n499 585
R1275 B.n499 B.n498 585
R1276 B.n743 B.n742 585
R1277 B.n744 B.n743 585
R1278 B.n493 B.n492 585
R1279 B.n494 B.n493 585
R1280 B.n752 B.n751 585
R1281 B.n751 B.n750 585
R1282 B.n753 B.n491 585
R1283 B.n491 B.n489 585
R1284 B.n755 B.n754 585
R1285 B.n756 B.n755 585
R1286 B.n485 B.n484 585
R1287 B.n490 B.n485 585
R1288 B.n764 B.n763 585
R1289 B.n763 B.n762 585
R1290 B.n765 B.n483 585
R1291 B.n483 B.n482 585
R1292 B.n767 B.n766 585
R1293 B.n768 B.n767 585
R1294 B.n477 B.n476 585
R1295 B.n478 B.n477 585
R1296 B.n776 B.n775 585
R1297 B.n775 B.n774 585
R1298 B.n777 B.n475 585
R1299 B.n475 B.n474 585
R1300 B.n779 B.n778 585
R1301 B.n780 B.n779 585
R1302 B.n469 B.n468 585
R1303 B.n470 B.n469 585
R1304 B.n788 B.n787 585
R1305 B.n787 B.n786 585
R1306 B.n789 B.n467 585
R1307 B.n467 B.n466 585
R1308 B.n791 B.n790 585
R1309 B.n792 B.n791 585
R1310 B.n461 B.n460 585
R1311 B.n462 B.n461 585
R1312 B.n801 B.n800 585
R1313 B.n800 B.n799 585
R1314 B.n802 B.n459 585
R1315 B.n798 B.n459 585
R1316 B.n804 B.n803 585
R1317 B.n805 B.n804 585
R1318 B.n454 B.n453 585
R1319 B.n455 B.n454 585
R1320 B.n813 B.n812 585
R1321 B.n812 B.n811 585
R1322 B.n814 B.n452 585
R1323 B.n452 B.n451 585
R1324 B.n816 B.n815 585
R1325 B.n817 B.n816 585
R1326 B.n446 B.n445 585
R1327 B.n447 B.n446 585
R1328 B.n825 B.n824 585
R1329 B.n824 B.n823 585
R1330 B.n826 B.n444 585
R1331 B.n444 B.n443 585
R1332 B.n828 B.n827 585
R1333 B.n829 B.n828 585
R1334 B.n438 B.n437 585
R1335 B.n439 B.n438 585
R1336 B.n837 B.n836 585
R1337 B.n836 B.n835 585
R1338 B.n838 B.n436 585
R1339 B.n436 B.n435 585
R1340 B.n840 B.n839 585
R1341 B.n841 B.n840 585
R1342 B.n430 B.n429 585
R1343 B.n431 B.n430 585
R1344 B.n849 B.n848 585
R1345 B.n848 B.n847 585
R1346 B.n850 B.n428 585
R1347 B.n428 B.n427 585
R1348 B.n852 B.n851 585
R1349 B.n853 B.n852 585
R1350 B.n422 B.n421 585
R1351 B.n423 B.n422 585
R1352 B.n861 B.n860 585
R1353 B.n860 B.n859 585
R1354 B.n862 B.n420 585
R1355 B.n420 B.n418 585
R1356 B.n864 B.n863 585
R1357 B.n865 B.n864 585
R1358 B.n414 B.n413 585
R1359 B.n419 B.n414 585
R1360 B.n873 B.n872 585
R1361 B.n872 B.n871 585
R1362 B.n874 B.n412 585
R1363 B.n412 B.n411 585
R1364 B.n876 B.n875 585
R1365 B.n877 B.n876 585
R1366 B.n406 B.n405 585
R1367 B.n407 B.n406 585
R1368 B.n885 B.n884 585
R1369 B.n884 B.n883 585
R1370 B.n886 B.n404 585
R1371 B.n404 B.n403 585
R1372 B.n888 B.n887 585
R1373 B.n889 B.n888 585
R1374 B.n398 B.n397 585
R1375 B.n399 B.n398 585
R1376 B.n897 B.n896 585
R1377 B.n896 B.n895 585
R1378 B.n898 B.n396 585
R1379 B.n396 B.n395 585
R1380 B.n900 B.n899 585
R1381 B.n901 B.n900 585
R1382 B.n390 B.n389 585
R1383 B.n391 B.n390 585
R1384 B.n909 B.n908 585
R1385 B.n908 B.n907 585
R1386 B.n910 B.n388 585
R1387 B.n388 B.n387 585
R1388 B.n912 B.n911 585
R1389 B.n913 B.n912 585
R1390 B.n382 B.n381 585
R1391 B.n383 B.n382 585
R1392 B.n921 B.n920 585
R1393 B.n920 B.n919 585
R1394 B.n922 B.n380 585
R1395 B.n380 B.n379 585
R1396 B.n924 B.n923 585
R1397 B.n925 B.n924 585
R1398 B.n374 B.n373 585
R1399 B.n375 B.n374 585
R1400 B.n934 B.n933 585
R1401 B.n933 B.n932 585
R1402 B.n935 B.n372 585
R1403 B.n931 B.n372 585
R1404 B.n937 B.n936 585
R1405 B.n938 B.n937 585
R1406 B.n367 B.n366 585
R1407 B.n368 B.n367 585
R1408 B.n947 B.n946 585
R1409 B.n946 B.n945 585
R1410 B.n948 B.n365 585
R1411 B.n365 B.n364 585
R1412 B.n950 B.n949 585
R1413 B.n951 B.n950 585
R1414 B.n3 B.n0 585
R1415 B.n4 B.n3 585
R1416 B.n1196 B.n1 585
R1417 B.n1197 B.n1196 585
R1418 B.n1195 B.n1194 585
R1419 B.n1195 B.n8 585
R1420 B.n1193 B.n9 585
R1421 B.n12 B.n9 585
R1422 B.n1192 B.n1191 585
R1423 B.n1191 B.n1190 585
R1424 B.n11 B.n10 585
R1425 B.n1189 B.n11 585
R1426 B.n1187 B.n1186 585
R1427 B.n1188 B.n1187 585
R1428 B.n1185 B.n16 585
R1429 B.n19 B.n16 585
R1430 B.n1184 B.n1183 585
R1431 B.n1183 B.n1182 585
R1432 B.n18 B.n17 585
R1433 B.n1181 B.n18 585
R1434 B.n1179 B.n1178 585
R1435 B.n1180 B.n1179 585
R1436 B.n1177 B.n24 585
R1437 B.n24 B.n23 585
R1438 B.n1176 B.n1175 585
R1439 B.n1175 B.n1174 585
R1440 B.n26 B.n25 585
R1441 B.n1173 B.n26 585
R1442 B.n1171 B.n1170 585
R1443 B.n1172 B.n1171 585
R1444 B.n1169 B.n31 585
R1445 B.n31 B.n30 585
R1446 B.n1168 B.n1167 585
R1447 B.n1167 B.n1166 585
R1448 B.n33 B.n32 585
R1449 B.n1165 B.n33 585
R1450 B.n1163 B.n1162 585
R1451 B.n1164 B.n1163 585
R1452 B.n1161 B.n38 585
R1453 B.n38 B.n37 585
R1454 B.n1160 B.n1159 585
R1455 B.n1159 B.n1158 585
R1456 B.n40 B.n39 585
R1457 B.n1157 B.n40 585
R1458 B.n1155 B.n1154 585
R1459 B.n1156 B.n1155 585
R1460 B.n1153 B.n45 585
R1461 B.n45 B.n44 585
R1462 B.n1152 B.n1151 585
R1463 B.n1151 B.n1150 585
R1464 B.n47 B.n46 585
R1465 B.n1149 B.n47 585
R1466 B.n1147 B.n1146 585
R1467 B.n1148 B.n1147 585
R1468 B.n1145 B.n52 585
R1469 B.n52 B.n51 585
R1470 B.n1144 B.n1143 585
R1471 B.n1143 B.n1142 585
R1472 B.n54 B.n53 585
R1473 B.n1141 B.n54 585
R1474 B.n1139 B.n1138 585
R1475 B.n1140 B.n1139 585
R1476 B.n1137 B.n59 585
R1477 B.n59 B.n58 585
R1478 B.n1136 B.n1135 585
R1479 B.n1135 B.n1134 585
R1480 B.n61 B.n60 585
R1481 B.n1133 B.n61 585
R1482 B.n1131 B.n1130 585
R1483 B.n1132 B.n1131 585
R1484 B.n1129 B.n66 585
R1485 B.n66 B.n65 585
R1486 B.n1128 B.n1127 585
R1487 B.n1127 B.n1126 585
R1488 B.n68 B.n67 585
R1489 B.n1125 B.n68 585
R1490 B.n1123 B.n1122 585
R1491 B.n1124 B.n1123 585
R1492 B.n1121 B.n73 585
R1493 B.n73 B.n72 585
R1494 B.n1120 B.n1119 585
R1495 B.n1119 B.n1118 585
R1496 B.n75 B.n74 585
R1497 B.n1117 B.n75 585
R1498 B.n1115 B.n1114 585
R1499 B.n1116 B.n1115 585
R1500 B.n1113 B.n80 585
R1501 B.n80 B.n79 585
R1502 B.n1112 B.n1111 585
R1503 B.n1111 B.n1110 585
R1504 B.n82 B.n81 585
R1505 B.n1109 B.n82 585
R1506 B.n1107 B.n1106 585
R1507 B.n1108 B.n1107 585
R1508 B.n1105 B.n87 585
R1509 B.n87 B.n86 585
R1510 B.n1104 B.n1103 585
R1511 B.n1103 B.n1102 585
R1512 B.n89 B.n88 585
R1513 B.n1101 B.n89 585
R1514 B.n1099 B.n1098 585
R1515 B.n1100 B.n1099 585
R1516 B.n1097 B.n93 585
R1517 B.n96 B.n93 585
R1518 B.n1096 B.n1095 585
R1519 B.n1095 B.n1094 585
R1520 B.n95 B.n94 585
R1521 B.n1093 B.n95 585
R1522 B.n1091 B.n1090 585
R1523 B.n1092 B.n1091 585
R1524 B.n1089 B.n101 585
R1525 B.n101 B.n100 585
R1526 B.n1088 B.n1087 585
R1527 B.n1087 B.n1086 585
R1528 B.n103 B.n102 585
R1529 B.n1085 B.n103 585
R1530 B.n1083 B.n1082 585
R1531 B.n1084 B.n1083 585
R1532 B.n1081 B.n108 585
R1533 B.n108 B.n107 585
R1534 B.n1080 B.n1079 585
R1535 B.n1079 B.n1078 585
R1536 B.n110 B.n109 585
R1537 B.n1077 B.n110 585
R1538 B.n1075 B.n1074 585
R1539 B.n1076 B.n1075 585
R1540 B.n1073 B.n115 585
R1541 B.n115 B.n114 585
R1542 B.n1072 B.n1071 585
R1543 B.n1071 B.n1070 585
R1544 B.n117 B.n116 585
R1545 B.n1069 B.n117 585
R1546 B.n1067 B.n1066 585
R1547 B.n1068 B.n1067 585
R1548 B.n1065 B.n122 585
R1549 B.n122 B.n121 585
R1550 B.n1064 B.n1063 585
R1551 B.n1063 B.n1062 585
R1552 B.n124 B.n123 585
R1553 B.n1061 B.n124 585
R1554 B.n1059 B.n1058 585
R1555 B.n1060 B.n1059 585
R1556 B.n1057 B.n129 585
R1557 B.n129 B.n128 585
R1558 B.n1056 B.n1055 585
R1559 B.n1055 B.n1054 585
R1560 B.n131 B.n130 585
R1561 B.n1053 B.n131 585
R1562 B.n1200 B.n1199 585
R1563 B.n1198 B.n2 585
R1564 B.n185 B.n131 554.963
R1565 B.n1050 B.n133 554.963
R1566 B.n733 B.n503 554.963
R1567 B.n730 B.n501 554.963
R1568 B.n179 B.t17 346.901
R1569 B.n553 B.t21 346.901
R1570 B.n182 B.t14 346.901
R1571 B.n551 B.t11 346.901
R1572 B.n182 B.t12 291.103
R1573 B.n179 B.t16 291.103
R1574 B.n553 B.t19 291.103
R1575 B.n551 B.t8 291.103
R1576 B.n180 B.t18 274.757
R1577 B.n554 B.t20 274.757
R1578 B.n183 B.t15 274.757
R1579 B.n552 B.t10 274.757
R1580 B.n1052 B.n1051 256.663
R1581 B.n1052 B.n177 256.663
R1582 B.n1052 B.n176 256.663
R1583 B.n1052 B.n175 256.663
R1584 B.n1052 B.n174 256.663
R1585 B.n1052 B.n173 256.663
R1586 B.n1052 B.n172 256.663
R1587 B.n1052 B.n171 256.663
R1588 B.n1052 B.n170 256.663
R1589 B.n1052 B.n169 256.663
R1590 B.n1052 B.n168 256.663
R1591 B.n1052 B.n167 256.663
R1592 B.n1052 B.n166 256.663
R1593 B.n1052 B.n165 256.663
R1594 B.n1052 B.n164 256.663
R1595 B.n1052 B.n163 256.663
R1596 B.n1052 B.n162 256.663
R1597 B.n1052 B.n161 256.663
R1598 B.n1052 B.n160 256.663
R1599 B.n1052 B.n159 256.663
R1600 B.n1052 B.n158 256.663
R1601 B.n1052 B.n157 256.663
R1602 B.n1052 B.n156 256.663
R1603 B.n1052 B.n155 256.663
R1604 B.n1052 B.n154 256.663
R1605 B.n1052 B.n153 256.663
R1606 B.n1052 B.n152 256.663
R1607 B.n1052 B.n151 256.663
R1608 B.n1052 B.n150 256.663
R1609 B.n1052 B.n149 256.663
R1610 B.n1052 B.n148 256.663
R1611 B.n1052 B.n147 256.663
R1612 B.n1052 B.n146 256.663
R1613 B.n1052 B.n145 256.663
R1614 B.n1052 B.n144 256.663
R1615 B.n1052 B.n143 256.663
R1616 B.n1052 B.n142 256.663
R1617 B.n1052 B.n141 256.663
R1618 B.n1052 B.n140 256.663
R1619 B.n1052 B.n139 256.663
R1620 B.n1052 B.n138 256.663
R1621 B.n1052 B.n137 256.663
R1622 B.n1052 B.n136 256.663
R1623 B.n1052 B.n135 256.663
R1624 B.n1052 B.n134 256.663
R1625 B.n732 B.n731 256.663
R1626 B.n732 B.n506 256.663
R1627 B.n732 B.n507 256.663
R1628 B.n732 B.n508 256.663
R1629 B.n732 B.n509 256.663
R1630 B.n732 B.n510 256.663
R1631 B.n732 B.n511 256.663
R1632 B.n732 B.n512 256.663
R1633 B.n732 B.n513 256.663
R1634 B.n732 B.n514 256.663
R1635 B.n732 B.n515 256.663
R1636 B.n732 B.n516 256.663
R1637 B.n732 B.n517 256.663
R1638 B.n732 B.n518 256.663
R1639 B.n732 B.n519 256.663
R1640 B.n732 B.n520 256.663
R1641 B.n732 B.n521 256.663
R1642 B.n732 B.n522 256.663
R1643 B.n732 B.n523 256.663
R1644 B.n732 B.n524 256.663
R1645 B.n732 B.n525 256.663
R1646 B.n732 B.n526 256.663
R1647 B.n732 B.n527 256.663
R1648 B.n732 B.n528 256.663
R1649 B.n732 B.n529 256.663
R1650 B.n732 B.n530 256.663
R1651 B.n732 B.n531 256.663
R1652 B.n732 B.n532 256.663
R1653 B.n732 B.n533 256.663
R1654 B.n732 B.n534 256.663
R1655 B.n732 B.n535 256.663
R1656 B.n732 B.n536 256.663
R1657 B.n732 B.n537 256.663
R1658 B.n732 B.n538 256.663
R1659 B.n732 B.n539 256.663
R1660 B.n732 B.n540 256.663
R1661 B.n732 B.n541 256.663
R1662 B.n732 B.n542 256.663
R1663 B.n732 B.n543 256.663
R1664 B.n732 B.n544 256.663
R1665 B.n732 B.n545 256.663
R1666 B.n732 B.n546 256.663
R1667 B.n732 B.n547 256.663
R1668 B.n732 B.n548 256.663
R1669 B.n1202 B.n1201 256.663
R1670 B.n189 B.n188 163.367
R1671 B.n193 B.n192 163.367
R1672 B.n197 B.n196 163.367
R1673 B.n201 B.n200 163.367
R1674 B.n205 B.n204 163.367
R1675 B.n209 B.n208 163.367
R1676 B.n213 B.n212 163.367
R1677 B.n217 B.n216 163.367
R1678 B.n221 B.n220 163.367
R1679 B.n225 B.n224 163.367
R1680 B.n229 B.n228 163.367
R1681 B.n233 B.n232 163.367
R1682 B.n237 B.n236 163.367
R1683 B.n241 B.n240 163.367
R1684 B.n245 B.n244 163.367
R1685 B.n249 B.n248 163.367
R1686 B.n253 B.n252 163.367
R1687 B.n257 B.n256 163.367
R1688 B.n261 B.n260 163.367
R1689 B.n265 B.n264 163.367
R1690 B.n269 B.n268 163.367
R1691 B.n273 B.n272 163.367
R1692 B.n277 B.n276 163.367
R1693 B.n281 B.n280 163.367
R1694 B.n285 B.n284 163.367
R1695 B.n289 B.n288 163.367
R1696 B.n293 B.n292 163.367
R1697 B.n297 B.n296 163.367
R1698 B.n301 B.n300 163.367
R1699 B.n305 B.n304 163.367
R1700 B.n309 B.n308 163.367
R1701 B.n313 B.n312 163.367
R1702 B.n317 B.n316 163.367
R1703 B.n321 B.n320 163.367
R1704 B.n325 B.n324 163.367
R1705 B.n329 B.n328 163.367
R1706 B.n333 B.n332 163.367
R1707 B.n337 B.n336 163.367
R1708 B.n341 B.n340 163.367
R1709 B.n345 B.n344 163.367
R1710 B.n349 B.n348 163.367
R1711 B.n353 B.n352 163.367
R1712 B.n357 B.n356 163.367
R1713 B.n359 B.n178 163.367
R1714 B.n737 B.n503 163.367
R1715 B.n737 B.n497 163.367
R1716 B.n745 B.n497 163.367
R1717 B.n745 B.n495 163.367
R1718 B.n749 B.n495 163.367
R1719 B.n749 B.n488 163.367
R1720 B.n757 B.n488 163.367
R1721 B.n757 B.n486 163.367
R1722 B.n761 B.n486 163.367
R1723 B.n761 B.n481 163.367
R1724 B.n769 B.n481 163.367
R1725 B.n769 B.n479 163.367
R1726 B.n773 B.n479 163.367
R1727 B.n773 B.n473 163.367
R1728 B.n781 B.n473 163.367
R1729 B.n781 B.n471 163.367
R1730 B.n785 B.n471 163.367
R1731 B.n785 B.n465 163.367
R1732 B.n793 B.n465 163.367
R1733 B.n793 B.n463 163.367
R1734 B.n797 B.n463 163.367
R1735 B.n797 B.n458 163.367
R1736 B.n806 B.n458 163.367
R1737 B.n806 B.n456 163.367
R1738 B.n810 B.n456 163.367
R1739 B.n810 B.n450 163.367
R1740 B.n818 B.n450 163.367
R1741 B.n818 B.n448 163.367
R1742 B.n822 B.n448 163.367
R1743 B.n822 B.n442 163.367
R1744 B.n830 B.n442 163.367
R1745 B.n830 B.n440 163.367
R1746 B.n834 B.n440 163.367
R1747 B.n834 B.n434 163.367
R1748 B.n842 B.n434 163.367
R1749 B.n842 B.n432 163.367
R1750 B.n846 B.n432 163.367
R1751 B.n846 B.n426 163.367
R1752 B.n854 B.n426 163.367
R1753 B.n854 B.n424 163.367
R1754 B.n858 B.n424 163.367
R1755 B.n858 B.n417 163.367
R1756 B.n866 B.n417 163.367
R1757 B.n866 B.n415 163.367
R1758 B.n870 B.n415 163.367
R1759 B.n870 B.n410 163.367
R1760 B.n878 B.n410 163.367
R1761 B.n878 B.n408 163.367
R1762 B.n882 B.n408 163.367
R1763 B.n882 B.n402 163.367
R1764 B.n890 B.n402 163.367
R1765 B.n890 B.n400 163.367
R1766 B.n894 B.n400 163.367
R1767 B.n894 B.n394 163.367
R1768 B.n902 B.n394 163.367
R1769 B.n902 B.n392 163.367
R1770 B.n906 B.n392 163.367
R1771 B.n906 B.n386 163.367
R1772 B.n914 B.n386 163.367
R1773 B.n914 B.n384 163.367
R1774 B.n918 B.n384 163.367
R1775 B.n918 B.n378 163.367
R1776 B.n926 B.n378 163.367
R1777 B.n926 B.n376 163.367
R1778 B.n930 B.n376 163.367
R1779 B.n930 B.n371 163.367
R1780 B.n939 B.n371 163.367
R1781 B.n939 B.n369 163.367
R1782 B.n944 B.n369 163.367
R1783 B.n944 B.n363 163.367
R1784 B.n952 B.n363 163.367
R1785 B.n953 B.n952 163.367
R1786 B.n953 B.n5 163.367
R1787 B.n6 B.n5 163.367
R1788 B.n7 B.n6 163.367
R1789 B.n959 B.n7 163.367
R1790 B.n960 B.n959 163.367
R1791 B.n960 B.n13 163.367
R1792 B.n14 B.n13 163.367
R1793 B.n15 B.n14 163.367
R1794 B.n965 B.n15 163.367
R1795 B.n965 B.n20 163.367
R1796 B.n21 B.n20 163.367
R1797 B.n22 B.n21 163.367
R1798 B.n970 B.n22 163.367
R1799 B.n970 B.n27 163.367
R1800 B.n28 B.n27 163.367
R1801 B.n29 B.n28 163.367
R1802 B.n975 B.n29 163.367
R1803 B.n975 B.n34 163.367
R1804 B.n35 B.n34 163.367
R1805 B.n36 B.n35 163.367
R1806 B.n980 B.n36 163.367
R1807 B.n980 B.n41 163.367
R1808 B.n42 B.n41 163.367
R1809 B.n43 B.n42 163.367
R1810 B.n985 B.n43 163.367
R1811 B.n985 B.n48 163.367
R1812 B.n49 B.n48 163.367
R1813 B.n50 B.n49 163.367
R1814 B.n990 B.n50 163.367
R1815 B.n990 B.n55 163.367
R1816 B.n56 B.n55 163.367
R1817 B.n57 B.n56 163.367
R1818 B.n995 B.n57 163.367
R1819 B.n995 B.n62 163.367
R1820 B.n63 B.n62 163.367
R1821 B.n64 B.n63 163.367
R1822 B.n1000 B.n64 163.367
R1823 B.n1000 B.n69 163.367
R1824 B.n70 B.n69 163.367
R1825 B.n71 B.n70 163.367
R1826 B.n1005 B.n71 163.367
R1827 B.n1005 B.n76 163.367
R1828 B.n77 B.n76 163.367
R1829 B.n78 B.n77 163.367
R1830 B.n1010 B.n78 163.367
R1831 B.n1010 B.n83 163.367
R1832 B.n84 B.n83 163.367
R1833 B.n85 B.n84 163.367
R1834 B.n1015 B.n85 163.367
R1835 B.n1015 B.n90 163.367
R1836 B.n91 B.n90 163.367
R1837 B.n92 B.n91 163.367
R1838 B.n1020 B.n92 163.367
R1839 B.n1020 B.n97 163.367
R1840 B.n98 B.n97 163.367
R1841 B.n99 B.n98 163.367
R1842 B.n1025 B.n99 163.367
R1843 B.n1025 B.n104 163.367
R1844 B.n105 B.n104 163.367
R1845 B.n106 B.n105 163.367
R1846 B.n1030 B.n106 163.367
R1847 B.n1030 B.n111 163.367
R1848 B.n112 B.n111 163.367
R1849 B.n113 B.n112 163.367
R1850 B.n1035 B.n113 163.367
R1851 B.n1035 B.n118 163.367
R1852 B.n119 B.n118 163.367
R1853 B.n120 B.n119 163.367
R1854 B.n1040 B.n120 163.367
R1855 B.n1040 B.n125 163.367
R1856 B.n126 B.n125 163.367
R1857 B.n127 B.n126 163.367
R1858 B.n1045 B.n127 163.367
R1859 B.n1045 B.n132 163.367
R1860 B.n133 B.n132 163.367
R1861 B.n550 B.n549 163.367
R1862 B.n725 B.n549 163.367
R1863 B.n723 B.n722 163.367
R1864 B.n719 B.n718 163.367
R1865 B.n715 B.n714 163.367
R1866 B.n711 B.n710 163.367
R1867 B.n707 B.n706 163.367
R1868 B.n703 B.n702 163.367
R1869 B.n699 B.n698 163.367
R1870 B.n695 B.n694 163.367
R1871 B.n691 B.n690 163.367
R1872 B.n687 B.n686 163.367
R1873 B.n683 B.n682 163.367
R1874 B.n679 B.n678 163.367
R1875 B.n675 B.n674 163.367
R1876 B.n671 B.n670 163.367
R1877 B.n667 B.n666 163.367
R1878 B.n663 B.n662 163.367
R1879 B.n659 B.n658 163.367
R1880 B.n655 B.n654 163.367
R1881 B.n650 B.n649 163.367
R1882 B.n646 B.n645 163.367
R1883 B.n642 B.n641 163.367
R1884 B.n638 B.n637 163.367
R1885 B.n634 B.n633 163.367
R1886 B.n629 B.n628 163.367
R1887 B.n625 B.n624 163.367
R1888 B.n621 B.n620 163.367
R1889 B.n617 B.n616 163.367
R1890 B.n613 B.n612 163.367
R1891 B.n609 B.n608 163.367
R1892 B.n605 B.n604 163.367
R1893 B.n601 B.n600 163.367
R1894 B.n597 B.n596 163.367
R1895 B.n593 B.n592 163.367
R1896 B.n589 B.n588 163.367
R1897 B.n585 B.n584 163.367
R1898 B.n581 B.n580 163.367
R1899 B.n577 B.n576 163.367
R1900 B.n573 B.n572 163.367
R1901 B.n569 B.n568 163.367
R1902 B.n565 B.n564 163.367
R1903 B.n561 B.n560 163.367
R1904 B.n557 B.n556 163.367
R1905 B.n733 B.n505 163.367
R1906 B.n739 B.n501 163.367
R1907 B.n739 B.n499 163.367
R1908 B.n743 B.n499 163.367
R1909 B.n743 B.n493 163.367
R1910 B.n751 B.n493 163.367
R1911 B.n751 B.n491 163.367
R1912 B.n755 B.n491 163.367
R1913 B.n755 B.n485 163.367
R1914 B.n763 B.n485 163.367
R1915 B.n763 B.n483 163.367
R1916 B.n767 B.n483 163.367
R1917 B.n767 B.n477 163.367
R1918 B.n775 B.n477 163.367
R1919 B.n775 B.n475 163.367
R1920 B.n779 B.n475 163.367
R1921 B.n779 B.n469 163.367
R1922 B.n787 B.n469 163.367
R1923 B.n787 B.n467 163.367
R1924 B.n791 B.n467 163.367
R1925 B.n791 B.n461 163.367
R1926 B.n800 B.n461 163.367
R1927 B.n800 B.n459 163.367
R1928 B.n804 B.n459 163.367
R1929 B.n804 B.n454 163.367
R1930 B.n812 B.n454 163.367
R1931 B.n812 B.n452 163.367
R1932 B.n816 B.n452 163.367
R1933 B.n816 B.n446 163.367
R1934 B.n824 B.n446 163.367
R1935 B.n824 B.n444 163.367
R1936 B.n828 B.n444 163.367
R1937 B.n828 B.n438 163.367
R1938 B.n836 B.n438 163.367
R1939 B.n836 B.n436 163.367
R1940 B.n840 B.n436 163.367
R1941 B.n840 B.n430 163.367
R1942 B.n848 B.n430 163.367
R1943 B.n848 B.n428 163.367
R1944 B.n852 B.n428 163.367
R1945 B.n852 B.n422 163.367
R1946 B.n860 B.n422 163.367
R1947 B.n860 B.n420 163.367
R1948 B.n864 B.n420 163.367
R1949 B.n864 B.n414 163.367
R1950 B.n872 B.n414 163.367
R1951 B.n872 B.n412 163.367
R1952 B.n876 B.n412 163.367
R1953 B.n876 B.n406 163.367
R1954 B.n884 B.n406 163.367
R1955 B.n884 B.n404 163.367
R1956 B.n888 B.n404 163.367
R1957 B.n888 B.n398 163.367
R1958 B.n896 B.n398 163.367
R1959 B.n896 B.n396 163.367
R1960 B.n900 B.n396 163.367
R1961 B.n900 B.n390 163.367
R1962 B.n908 B.n390 163.367
R1963 B.n908 B.n388 163.367
R1964 B.n912 B.n388 163.367
R1965 B.n912 B.n382 163.367
R1966 B.n920 B.n382 163.367
R1967 B.n920 B.n380 163.367
R1968 B.n924 B.n380 163.367
R1969 B.n924 B.n374 163.367
R1970 B.n933 B.n374 163.367
R1971 B.n933 B.n372 163.367
R1972 B.n937 B.n372 163.367
R1973 B.n937 B.n367 163.367
R1974 B.n946 B.n367 163.367
R1975 B.n946 B.n365 163.367
R1976 B.n950 B.n365 163.367
R1977 B.n950 B.n3 163.367
R1978 B.n1200 B.n3 163.367
R1979 B.n1196 B.n2 163.367
R1980 B.n1196 B.n1195 163.367
R1981 B.n1195 B.n9 163.367
R1982 B.n1191 B.n9 163.367
R1983 B.n1191 B.n11 163.367
R1984 B.n1187 B.n11 163.367
R1985 B.n1187 B.n16 163.367
R1986 B.n1183 B.n16 163.367
R1987 B.n1183 B.n18 163.367
R1988 B.n1179 B.n18 163.367
R1989 B.n1179 B.n24 163.367
R1990 B.n1175 B.n24 163.367
R1991 B.n1175 B.n26 163.367
R1992 B.n1171 B.n26 163.367
R1993 B.n1171 B.n31 163.367
R1994 B.n1167 B.n31 163.367
R1995 B.n1167 B.n33 163.367
R1996 B.n1163 B.n33 163.367
R1997 B.n1163 B.n38 163.367
R1998 B.n1159 B.n38 163.367
R1999 B.n1159 B.n40 163.367
R2000 B.n1155 B.n40 163.367
R2001 B.n1155 B.n45 163.367
R2002 B.n1151 B.n45 163.367
R2003 B.n1151 B.n47 163.367
R2004 B.n1147 B.n47 163.367
R2005 B.n1147 B.n52 163.367
R2006 B.n1143 B.n52 163.367
R2007 B.n1143 B.n54 163.367
R2008 B.n1139 B.n54 163.367
R2009 B.n1139 B.n59 163.367
R2010 B.n1135 B.n59 163.367
R2011 B.n1135 B.n61 163.367
R2012 B.n1131 B.n61 163.367
R2013 B.n1131 B.n66 163.367
R2014 B.n1127 B.n66 163.367
R2015 B.n1127 B.n68 163.367
R2016 B.n1123 B.n68 163.367
R2017 B.n1123 B.n73 163.367
R2018 B.n1119 B.n73 163.367
R2019 B.n1119 B.n75 163.367
R2020 B.n1115 B.n75 163.367
R2021 B.n1115 B.n80 163.367
R2022 B.n1111 B.n80 163.367
R2023 B.n1111 B.n82 163.367
R2024 B.n1107 B.n82 163.367
R2025 B.n1107 B.n87 163.367
R2026 B.n1103 B.n87 163.367
R2027 B.n1103 B.n89 163.367
R2028 B.n1099 B.n89 163.367
R2029 B.n1099 B.n93 163.367
R2030 B.n1095 B.n93 163.367
R2031 B.n1095 B.n95 163.367
R2032 B.n1091 B.n95 163.367
R2033 B.n1091 B.n101 163.367
R2034 B.n1087 B.n101 163.367
R2035 B.n1087 B.n103 163.367
R2036 B.n1083 B.n103 163.367
R2037 B.n1083 B.n108 163.367
R2038 B.n1079 B.n108 163.367
R2039 B.n1079 B.n110 163.367
R2040 B.n1075 B.n110 163.367
R2041 B.n1075 B.n115 163.367
R2042 B.n1071 B.n115 163.367
R2043 B.n1071 B.n117 163.367
R2044 B.n1067 B.n117 163.367
R2045 B.n1067 B.n122 163.367
R2046 B.n1063 B.n122 163.367
R2047 B.n1063 B.n124 163.367
R2048 B.n1059 B.n124 163.367
R2049 B.n1059 B.n129 163.367
R2050 B.n1055 B.n129 163.367
R2051 B.n1055 B.n131 163.367
R2052 B.n732 B.n502 92.1847
R2053 B.n1053 B.n1052 92.1847
R2054 B.n183 B.n182 72.146
R2055 B.n180 B.n179 72.146
R2056 B.n554 B.n553 72.146
R2057 B.n552 B.n551 72.146
R2058 B.n185 B.n134 71.676
R2059 B.n189 B.n135 71.676
R2060 B.n193 B.n136 71.676
R2061 B.n197 B.n137 71.676
R2062 B.n201 B.n138 71.676
R2063 B.n205 B.n139 71.676
R2064 B.n209 B.n140 71.676
R2065 B.n213 B.n141 71.676
R2066 B.n217 B.n142 71.676
R2067 B.n221 B.n143 71.676
R2068 B.n225 B.n144 71.676
R2069 B.n229 B.n145 71.676
R2070 B.n233 B.n146 71.676
R2071 B.n237 B.n147 71.676
R2072 B.n241 B.n148 71.676
R2073 B.n245 B.n149 71.676
R2074 B.n249 B.n150 71.676
R2075 B.n253 B.n151 71.676
R2076 B.n257 B.n152 71.676
R2077 B.n261 B.n153 71.676
R2078 B.n265 B.n154 71.676
R2079 B.n269 B.n155 71.676
R2080 B.n273 B.n156 71.676
R2081 B.n277 B.n157 71.676
R2082 B.n281 B.n158 71.676
R2083 B.n285 B.n159 71.676
R2084 B.n289 B.n160 71.676
R2085 B.n293 B.n161 71.676
R2086 B.n297 B.n162 71.676
R2087 B.n301 B.n163 71.676
R2088 B.n305 B.n164 71.676
R2089 B.n309 B.n165 71.676
R2090 B.n313 B.n166 71.676
R2091 B.n317 B.n167 71.676
R2092 B.n321 B.n168 71.676
R2093 B.n325 B.n169 71.676
R2094 B.n329 B.n170 71.676
R2095 B.n333 B.n171 71.676
R2096 B.n337 B.n172 71.676
R2097 B.n341 B.n173 71.676
R2098 B.n345 B.n174 71.676
R2099 B.n349 B.n175 71.676
R2100 B.n353 B.n176 71.676
R2101 B.n357 B.n177 71.676
R2102 B.n1051 B.n178 71.676
R2103 B.n1051 B.n1050 71.676
R2104 B.n359 B.n177 71.676
R2105 B.n356 B.n176 71.676
R2106 B.n352 B.n175 71.676
R2107 B.n348 B.n174 71.676
R2108 B.n344 B.n173 71.676
R2109 B.n340 B.n172 71.676
R2110 B.n336 B.n171 71.676
R2111 B.n332 B.n170 71.676
R2112 B.n328 B.n169 71.676
R2113 B.n324 B.n168 71.676
R2114 B.n320 B.n167 71.676
R2115 B.n316 B.n166 71.676
R2116 B.n312 B.n165 71.676
R2117 B.n308 B.n164 71.676
R2118 B.n304 B.n163 71.676
R2119 B.n300 B.n162 71.676
R2120 B.n296 B.n161 71.676
R2121 B.n292 B.n160 71.676
R2122 B.n288 B.n159 71.676
R2123 B.n284 B.n158 71.676
R2124 B.n280 B.n157 71.676
R2125 B.n276 B.n156 71.676
R2126 B.n272 B.n155 71.676
R2127 B.n268 B.n154 71.676
R2128 B.n264 B.n153 71.676
R2129 B.n260 B.n152 71.676
R2130 B.n256 B.n151 71.676
R2131 B.n252 B.n150 71.676
R2132 B.n248 B.n149 71.676
R2133 B.n244 B.n148 71.676
R2134 B.n240 B.n147 71.676
R2135 B.n236 B.n146 71.676
R2136 B.n232 B.n145 71.676
R2137 B.n228 B.n144 71.676
R2138 B.n224 B.n143 71.676
R2139 B.n220 B.n142 71.676
R2140 B.n216 B.n141 71.676
R2141 B.n212 B.n140 71.676
R2142 B.n208 B.n139 71.676
R2143 B.n204 B.n138 71.676
R2144 B.n200 B.n137 71.676
R2145 B.n196 B.n136 71.676
R2146 B.n192 B.n135 71.676
R2147 B.n188 B.n134 71.676
R2148 B.n731 B.n730 71.676
R2149 B.n725 B.n506 71.676
R2150 B.n722 B.n507 71.676
R2151 B.n718 B.n508 71.676
R2152 B.n714 B.n509 71.676
R2153 B.n710 B.n510 71.676
R2154 B.n706 B.n511 71.676
R2155 B.n702 B.n512 71.676
R2156 B.n698 B.n513 71.676
R2157 B.n694 B.n514 71.676
R2158 B.n690 B.n515 71.676
R2159 B.n686 B.n516 71.676
R2160 B.n682 B.n517 71.676
R2161 B.n678 B.n518 71.676
R2162 B.n674 B.n519 71.676
R2163 B.n670 B.n520 71.676
R2164 B.n666 B.n521 71.676
R2165 B.n662 B.n522 71.676
R2166 B.n658 B.n523 71.676
R2167 B.n654 B.n524 71.676
R2168 B.n649 B.n525 71.676
R2169 B.n645 B.n526 71.676
R2170 B.n641 B.n527 71.676
R2171 B.n637 B.n528 71.676
R2172 B.n633 B.n529 71.676
R2173 B.n628 B.n530 71.676
R2174 B.n624 B.n531 71.676
R2175 B.n620 B.n532 71.676
R2176 B.n616 B.n533 71.676
R2177 B.n612 B.n534 71.676
R2178 B.n608 B.n535 71.676
R2179 B.n604 B.n536 71.676
R2180 B.n600 B.n537 71.676
R2181 B.n596 B.n538 71.676
R2182 B.n592 B.n539 71.676
R2183 B.n588 B.n540 71.676
R2184 B.n584 B.n541 71.676
R2185 B.n580 B.n542 71.676
R2186 B.n576 B.n543 71.676
R2187 B.n572 B.n544 71.676
R2188 B.n568 B.n545 71.676
R2189 B.n564 B.n546 71.676
R2190 B.n560 B.n547 71.676
R2191 B.n556 B.n548 71.676
R2192 B.n731 B.n550 71.676
R2193 B.n723 B.n506 71.676
R2194 B.n719 B.n507 71.676
R2195 B.n715 B.n508 71.676
R2196 B.n711 B.n509 71.676
R2197 B.n707 B.n510 71.676
R2198 B.n703 B.n511 71.676
R2199 B.n699 B.n512 71.676
R2200 B.n695 B.n513 71.676
R2201 B.n691 B.n514 71.676
R2202 B.n687 B.n515 71.676
R2203 B.n683 B.n516 71.676
R2204 B.n679 B.n517 71.676
R2205 B.n675 B.n518 71.676
R2206 B.n671 B.n519 71.676
R2207 B.n667 B.n520 71.676
R2208 B.n663 B.n521 71.676
R2209 B.n659 B.n522 71.676
R2210 B.n655 B.n523 71.676
R2211 B.n650 B.n524 71.676
R2212 B.n646 B.n525 71.676
R2213 B.n642 B.n526 71.676
R2214 B.n638 B.n527 71.676
R2215 B.n634 B.n528 71.676
R2216 B.n629 B.n529 71.676
R2217 B.n625 B.n530 71.676
R2218 B.n621 B.n531 71.676
R2219 B.n617 B.n532 71.676
R2220 B.n613 B.n533 71.676
R2221 B.n609 B.n534 71.676
R2222 B.n605 B.n535 71.676
R2223 B.n601 B.n536 71.676
R2224 B.n597 B.n537 71.676
R2225 B.n593 B.n538 71.676
R2226 B.n589 B.n539 71.676
R2227 B.n585 B.n540 71.676
R2228 B.n581 B.n541 71.676
R2229 B.n577 B.n542 71.676
R2230 B.n573 B.n543 71.676
R2231 B.n569 B.n544 71.676
R2232 B.n565 B.n545 71.676
R2233 B.n561 B.n546 71.676
R2234 B.n557 B.n547 71.676
R2235 B.n548 B.n505 71.676
R2236 B.n1201 B.n1200 71.676
R2237 B.n1201 B.n2 71.676
R2238 B.n184 B.n183 59.5399
R2239 B.n181 B.n180 59.5399
R2240 B.n631 B.n554 59.5399
R2241 B.n652 B.n552 59.5399
R2242 B.n738 B.n502 44.4582
R2243 B.n738 B.n498 44.4582
R2244 B.n744 B.n498 44.4582
R2245 B.n744 B.n494 44.4582
R2246 B.n750 B.n494 44.4582
R2247 B.n750 B.n489 44.4582
R2248 B.n756 B.n489 44.4582
R2249 B.n756 B.n490 44.4582
R2250 B.n762 B.n482 44.4582
R2251 B.n768 B.n482 44.4582
R2252 B.n768 B.n478 44.4582
R2253 B.n774 B.n478 44.4582
R2254 B.n774 B.n474 44.4582
R2255 B.n780 B.n474 44.4582
R2256 B.n780 B.n470 44.4582
R2257 B.n786 B.n470 44.4582
R2258 B.n786 B.n466 44.4582
R2259 B.n792 B.n466 44.4582
R2260 B.n792 B.n462 44.4582
R2261 B.n799 B.n462 44.4582
R2262 B.n799 B.n798 44.4582
R2263 B.n805 B.n455 44.4582
R2264 B.n811 B.n455 44.4582
R2265 B.n811 B.n451 44.4582
R2266 B.n817 B.n451 44.4582
R2267 B.n817 B.n447 44.4582
R2268 B.n823 B.n447 44.4582
R2269 B.n823 B.n443 44.4582
R2270 B.n829 B.n443 44.4582
R2271 B.n829 B.n439 44.4582
R2272 B.n835 B.n439 44.4582
R2273 B.n841 B.n435 44.4582
R2274 B.n841 B.n431 44.4582
R2275 B.n847 B.n431 44.4582
R2276 B.n847 B.n427 44.4582
R2277 B.n853 B.n427 44.4582
R2278 B.n853 B.n423 44.4582
R2279 B.n859 B.n423 44.4582
R2280 B.n859 B.n418 44.4582
R2281 B.n865 B.n418 44.4582
R2282 B.n865 B.n419 44.4582
R2283 B.n871 B.n411 44.4582
R2284 B.n877 B.n411 44.4582
R2285 B.n877 B.n407 44.4582
R2286 B.n883 B.n407 44.4582
R2287 B.n883 B.n403 44.4582
R2288 B.n889 B.n403 44.4582
R2289 B.n889 B.n399 44.4582
R2290 B.n895 B.n399 44.4582
R2291 B.n895 B.n395 44.4582
R2292 B.n901 B.n395 44.4582
R2293 B.n907 B.n391 44.4582
R2294 B.n907 B.n387 44.4582
R2295 B.n913 B.n387 44.4582
R2296 B.n913 B.n383 44.4582
R2297 B.n919 B.n383 44.4582
R2298 B.n919 B.n379 44.4582
R2299 B.n925 B.n379 44.4582
R2300 B.n925 B.n375 44.4582
R2301 B.n932 B.n375 44.4582
R2302 B.n932 B.n931 44.4582
R2303 B.n938 B.n368 44.4582
R2304 B.n945 B.n368 44.4582
R2305 B.n945 B.n364 44.4582
R2306 B.n951 B.n364 44.4582
R2307 B.n951 B.n4 44.4582
R2308 B.n1199 B.n4 44.4582
R2309 B.n1199 B.n1198 44.4582
R2310 B.n1198 B.n1197 44.4582
R2311 B.n1197 B.n8 44.4582
R2312 B.n12 B.n8 44.4582
R2313 B.n1190 B.n12 44.4582
R2314 B.n1190 B.n1189 44.4582
R2315 B.n1189 B.n1188 44.4582
R2316 B.n1182 B.n19 44.4582
R2317 B.n1182 B.n1181 44.4582
R2318 B.n1181 B.n1180 44.4582
R2319 B.n1180 B.n23 44.4582
R2320 B.n1174 B.n23 44.4582
R2321 B.n1174 B.n1173 44.4582
R2322 B.n1173 B.n1172 44.4582
R2323 B.n1172 B.n30 44.4582
R2324 B.n1166 B.n30 44.4582
R2325 B.n1166 B.n1165 44.4582
R2326 B.n1164 B.n37 44.4582
R2327 B.n1158 B.n37 44.4582
R2328 B.n1158 B.n1157 44.4582
R2329 B.n1157 B.n1156 44.4582
R2330 B.n1156 B.n44 44.4582
R2331 B.n1150 B.n44 44.4582
R2332 B.n1150 B.n1149 44.4582
R2333 B.n1149 B.n1148 44.4582
R2334 B.n1148 B.n51 44.4582
R2335 B.n1142 B.n51 44.4582
R2336 B.n1141 B.n1140 44.4582
R2337 B.n1140 B.n58 44.4582
R2338 B.n1134 B.n58 44.4582
R2339 B.n1134 B.n1133 44.4582
R2340 B.n1133 B.n1132 44.4582
R2341 B.n1132 B.n65 44.4582
R2342 B.n1126 B.n65 44.4582
R2343 B.n1126 B.n1125 44.4582
R2344 B.n1125 B.n1124 44.4582
R2345 B.n1124 B.n72 44.4582
R2346 B.n1118 B.n1117 44.4582
R2347 B.n1117 B.n1116 44.4582
R2348 B.n1116 B.n79 44.4582
R2349 B.n1110 B.n79 44.4582
R2350 B.n1110 B.n1109 44.4582
R2351 B.n1109 B.n1108 44.4582
R2352 B.n1108 B.n86 44.4582
R2353 B.n1102 B.n86 44.4582
R2354 B.n1102 B.n1101 44.4582
R2355 B.n1101 B.n1100 44.4582
R2356 B.n1094 B.n96 44.4582
R2357 B.n1094 B.n1093 44.4582
R2358 B.n1093 B.n1092 44.4582
R2359 B.n1092 B.n100 44.4582
R2360 B.n1086 B.n100 44.4582
R2361 B.n1086 B.n1085 44.4582
R2362 B.n1085 B.n1084 44.4582
R2363 B.n1084 B.n107 44.4582
R2364 B.n1078 B.n107 44.4582
R2365 B.n1078 B.n1077 44.4582
R2366 B.n1077 B.n1076 44.4582
R2367 B.n1076 B.n114 44.4582
R2368 B.n1070 B.n114 44.4582
R2369 B.n1069 B.n1068 44.4582
R2370 B.n1068 B.n121 44.4582
R2371 B.n1062 B.n121 44.4582
R2372 B.n1062 B.n1061 44.4582
R2373 B.n1061 B.n1060 44.4582
R2374 B.n1060 B.n128 44.4582
R2375 B.n1054 B.n128 44.4582
R2376 B.n1054 B.n1053 44.4582
R2377 B.n1049 B.n1048 36.059
R2378 B.n729 B.n500 36.059
R2379 B.n735 B.n734 36.059
R2380 B.n186 B.n130 36.059
R2381 B.n798 B.t6 29.421
R2382 B.n96 B.t3 29.421
R2383 B.n835 B.t22 26.8058
R2384 B.n1118 B.t4 26.8058
R2385 B.n938 B.t5 25.4983
R2386 B.n1188 B.t2 25.4983
R2387 B.n419 B.t7 24.1907
R2388 B.t1 B.n1141 24.1907
R2389 B.n490 B.t9 22.8831
R2390 B.t23 B.n391 22.8831
R2391 B.n1165 B.t0 22.8831
R2392 B.t13 B.n1069 22.8831
R2393 B.n762 B.t9 21.5755
R2394 B.n901 B.t23 21.5755
R2395 B.t0 B.n1164 21.5755
R2396 B.n1070 B.t13 21.5755
R2397 B.n871 B.t7 20.268
R2398 B.n1142 B.t1 20.268
R2399 B.n931 B.t5 18.9604
R2400 B.n19 B.t2 18.9604
R2401 B B.n1202 18.0485
R2402 B.t22 B.n435 17.6528
R2403 B.t4 B.n72 17.6528
R2404 B.n805 B.t6 15.0376
R2405 B.n1100 B.t3 15.0376
R2406 B.n740 B.n500 10.6151
R2407 B.n741 B.n740 10.6151
R2408 B.n742 B.n741 10.6151
R2409 B.n742 B.n492 10.6151
R2410 B.n752 B.n492 10.6151
R2411 B.n753 B.n752 10.6151
R2412 B.n754 B.n753 10.6151
R2413 B.n754 B.n484 10.6151
R2414 B.n764 B.n484 10.6151
R2415 B.n765 B.n764 10.6151
R2416 B.n766 B.n765 10.6151
R2417 B.n766 B.n476 10.6151
R2418 B.n776 B.n476 10.6151
R2419 B.n777 B.n776 10.6151
R2420 B.n778 B.n777 10.6151
R2421 B.n778 B.n468 10.6151
R2422 B.n788 B.n468 10.6151
R2423 B.n789 B.n788 10.6151
R2424 B.n790 B.n789 10.6151
R2425 B.n790 B.n460 10.6151
R2426 B.n801 B.n460 10.6151
R2427 B.n802 B.n801 10.6151
R2428 B.n803 B.n802 10.6151
R2429 B.n803 B.n453 10.6151
R2430 B.n813 B.n453 10.6151
R2431 B.n814 B.n813 10.6151
R2432 B.n815 B.n814 10.6151
R2433 B.n815 B.n445 10.6151
R2434 B.n825 B.n445 10.6151
R2435 B.n826 B.n825 10.6151
R2436 B.n827 B.n826 10.6151
R2437 B.n827 B.n437 10.6151
R2438 B.n837 B.n437 10.6151
R2439 B.n838 B.n837 10.6151
R2440 B.n839 B.n838 10.6151
R2441 B.n839 B.n429 10.6151
R2442 B.n849 B.n429 10.6151
R2443 B.n850 B.n849 10.6151
R2444 B.n851 B.n850 10.6151
R2445 B.n851 B.n421 10.6151
R2446 B.n861 B.n421 10.6151
R2447 B.n862 B.n861 10.6151
R2448 B.n863 B.n862 10.6151
R2449 B.n863 B.n413 10.6151
R2450 B.n873 B.n413 10.6151
R2451 B.n874 B.n873 10.6151
R2452 B.n875 B.n874 10.6151
R2453 B.n875 B.n405 10.6151
R2454 B.n885 B.n405 10.6151
R2455 B.n886 B.n885 10.6151
R2456 B.n887 B.n886 10.6151
R2457 B.n887 B.n397 10.6151
R2458 B.n897 B.n397 10.6151
R2459 B.n898 B.n897 10.6151
R2460 B.n899 B.n898 10.6151
R2461 B.n899 B.n389 10.6151
R2462 B.n909 B.n389 10.6151
R2463 B.n910 B.n909 10.6151
R2464 B.n911 B.n910 10.6151
R2465 B.n911 B.n381 10.6151
R2466 B.n921 B.n381 10.6151
R2467 B.n922 B.n921 10.6151
R2468 B.n923 B.n922 10.6151
R2469 B.n923 B.n373 10.6151
R2470 B.n934 B.n373 10.6151
R2471 B.n935 B.n934 10.6151
R2472 B.n936 B.n935 10.6151
R2473 B.n936 B.n366 10.6151
R2474 B.n947 B.n366 10.6151
R2475 B.n948 B.n947 10.6151
R2476 B.n949 B.n948 10.6151
R2477 B.n949 B.n0 10.6151
R2478 B.n729 B.n728 10.6151
R2479 B.n728 B.n727 10.6151
R2480 B.n727 B.n726 10.6151
R2481 B.n726 B.n724 10.6151
R2482 B.n724 B.n721 10.6151
R2483 B.n721 B.n720 10.6151
R2484 B.n720 B.n717 10.6151
R2485 B.n717 B.n716 10.6151
R2486 B.n716 B.n713 10.6151
R2487 B.n713 B.n712 10.6151
R2488 B.n712 B.n709 10.6151
R2489 B.n709 B.n708 10.6151
R2490 B.n708 B.n705 10.6151
R2491 B.n705 B.n704 10.6151
R2492 B.n704 B.n701 10.6151
R2493 B.n701 B.n700 10.6151
R2494 B.n700 B.n697 10.6151
R2495 B.n697 B.n696 10.6151
R2496 B.n696 B.n693 10.6151
R2497 B.n693 B.n692 10.6151
R2498 B.n692 B.n689 10.6151
R2499 B.n689 B.n688 10.6151
R2500 B.n688 B.n685 10.6151
R2501 B.n685 B.n684 10.6151
R2502 B.n684 B.n681 10.6151
R2503 B.n681 B.n680 10.6151
R2504 B.n680 B.n677 10.6151
R2505 B.n677 B.n676 10.6151
R2506 B.n676 B.n673 10.6151
R2507 B.n673 B.n672 10.6151
R2508 B.n672 B.n669 10.6151
R2509 B.n669 B.n668 10.6151
R2510 B.n668 B.n665 10.6151
R2511 B.n665 B.n664 10.6151
R2512 B.n664 B.n661 10.6151
R2513 B.n661 B.n660 10.6151
R2514 B.n660 B.n657 10.6151
R2515 B.n657 B.n656 10.6151
R2516 B.n656 B.n653 10.6151
R2517 B.n651 B.n648 10.6151
R2518 B.n648 B.n647 10.6151
R2519 B.n647 B.n644 10.6151
R2520 B.n644 B.n643 10.6151
R2521 B.n643 B.n640 10.6151
R2522 B.n640 B.n639 10.6151
R2523 B.n639 B.n636 10.6151
R2524 B.n636 B.n635 10.6151
R2525 B.n635 B.n632 10.6151
R2526 B.n630 B.n627 10.6151
R2527 B.n627 B.n626 10.6151
R2528 B.n626 B.n623 10.6151
R2529 B.n623 B.n622 10.6151
R2530 B.n622 B.n619 10.6151
R2531 B.n619 B.n618 10.6151
R2532 B.n618 B.n615 10.6151
R2533 B.n615 B.n614 10.6151
R2534 B.n614 B.n611 10.6151
R2535 B.n611 B.n610 10.6151
R2536 B.n610 B.n607 10.6151
R2537 B.n607 B.n606 10.6151
R2538 B.n606 B.n603 10.6151
R2539 B.n603 B.n602 10.6151
R2540 B.n602 B.n599 10.6151
R2541 B.n599 B.n598 10.6151
R2542 B.n598 B.n595 10.6151
R2543 B.n595 B.n594 10.6151
R2544 B.n594 B.n591 10.6151
R2545 B.n591 B.n590 10.6151
R2546 B.n590 B.n587 10.6151
R2547 B.n587 B.n586 10.6151
R2548 B.n586 B.n583 10.6151
R2549 B.n583 B.n582 10.6151
R2550 B.n582 B.n579 10.6151
R2551 B.n579 B.n578 10.6151
R2552 B.n578 B.n575 10.6151
R2553 B.n575 B.n574 10.6151
R2554 B.n574 B.n571 10.6151
R2555 B.n571 B.n570 10.6151
R2556 B.n570 B.n567 10.6151
R2557 B.n567 B.n566 10.6151
R2558 B.n566 B.n563 10.6151
R2559 B.n563 B.n562 10.6151
R2560 B.n562 B.n559 10.6151
R2561 B.n559 B.n558 10.6151
R2562 B.n558 B.n555 10.6151
R2563 B.n555 B.n504 10.6151
R2564 B.n734 B.n504 10.6151
R2565 B.n736 B.n735 10.6151
R2566 B.n736 B.n496 10.6151
R2567 B.n746 B.n496 10.6151
R2568 B.n747 B.n746 10.6151
R2569 B.n748 B.n747 10.6151
R2570 B.n748 B.n487 10.6151
R2571 B.n758 B.n487 10.6151
R2572 B.n759 B.n758 10.6151
R2573 B.n760 B.n759 10.6151
R2574 B.n760 B.n480 10.6151
R2575 B.n770 B.n480 10.6151
R2576 B.n771 B.n770 10.6151
R2577 B.n772 B.n771 10.6151
R2578 B.n772 B.n472 10.6151
R2579 B.n782 B.n472 10.6151
R2580 B.n783 B.n782 10.6151
R2581 B.n784 B.n783 10.6151
R2582 B.n784 B.n464 10.6151
R2583 B.n794 B.n464 10.6151
R2584 B.n795 B.n794 10.6151
R2585 B.n796 B.n795 10.6151
R2586 B.n796 B.n457 10.6151
R2587 B.n807 B.n457 10.6151
R2588 B.n808 B.n807 10.6151
R2589 B.n809 B.n808 10.6151
R2590 B.n809 B.n449 10.6151
R2591 B.n819 B.n449 10.6151
R2592 B.n820 B.n819 10.6151
R2593 B.n821 B.n820 10.6151
R2594 B.n821 B.n441 10.6151
R2595 B.n831 B.n441 10.6151
R2596 B.n832 B.n831 10.6151
R2597 B.n833 B.n832 10.6151
R2598 B.n833 B.n433 10.6151
R2599 B.n843 B.n433 10.6151
R2600 B.n844 B.n843 10.6151
R2601 B.n845 B.n844 10.6151
R2602 B.n845 B.n425 10.6151
R2603 B.n855 B.n425 10.6151
R2604 B.n856 B.n855 10.6151
R2605 B.n857 B.n856 10.6151
R2606 B.n857 B.n416 10.6151
R2607 B.n867 B.n416 10.6151
R2608 B.n868 B.n867 10.6151
R2609 B.n869 B.n868 10.6151
R2610 B.n869 B.n409 10.6151
R2611 B.n879 B.n409 10.6151
R2612 B.n880 B.n879 10.6151
R2613 B.n881 B.n880 10.6151
R2614 B.n881 B.n401 10.6151
R2615 B.n891 B.n401 10.6151
R2616 B.n892 B.n891 10.6151
R2617 B.n893 B.n892 10.6151
R2618 B.n893 B.n393 10.6151
R2619 B.n903 B.n393 10.6151
R2620 B.n904 B.n903 10.6151
R2621 B.n905 B.n904 10.6151
R2622 B.n905 B.n385 10.6151
R2623 B.n915 B.n385 10.6151
R2624 B.n916 B.n915 10.6151
R2625 B.n917 B.n916 10.6151
R2626 B.n917 B.n377 10.6151
R2627 B.n927 B.n377 10.6151
R2628 B.n928 B.n927 10.6151
R2629 B.n929 B.n928 10.6151
R2630 B.n929 B.n370 10.6151
R2631 B.n940 B.n370 10.6151
R2632 B.n941 B.n940 10.6151
R2633 B.n943 B.n941 10.6151
R2634 B.n943 B.n942 10.6151
R2635 B.n942 B.n362 10.6151
R2636 B.n954 B.n362 10.6151
R2637 B.n955 B.n954 10.6151
R2638 B.n956 B.n955 10.6151
R2639 B.n957 B.n956 10.6151
R2640 B.n958 B.n957 10.6151
R2641 B.n961 B.n958 10.6151
R2642 B.n962 B.n961 10.6151
R2643 B.n963 B.n962 10.6151
R2644 B.n964 B.n963 10.6151
R2645 B.n966 B.n964 10.6151
R2646 B.n967 B.n966 10.6151
R2647 B.n968 B.n967 10.6151
R2648 B.n969 B.n968 10.6151
R2649 B.n971 B.n969 10.6151
R2650 B.n972 B.n971 10.6151
R2651 B.n973 B.n972 10.6151
R2652 B.n974 B.n973 10.6151
R2653 B.n976 B.n974 10.6151
R2654 B.n977 B.n976 10.6151
R2655 B.n978 B.n977 10.6151
R2656 B.n979 B.n978 10.6151
R2657 B.n981 B.n979 10.6151
R2658 B.n982 B.n981 10.6151
R2659 B.n983 B.n982 10.6151
R2660 B.n984 B.n983 10.6151
R2661 B.n986 B.n984 10.6151
R2662 B.n987 B.n986 10.6151
R2663 B.n988 B.n987 10.6151
R2664 B.n989 B.n988 10.6151
R2665 B.n991 B.n989 10.6151
R2666 B.n992 B.n991 10.6151
R2667 B.n993 B.n992 10.6151
R2668 B.n994 B.n993 10.6151
R2669 B.n996 B.n994 10.6151
R2670 B.n997 B.n996 10.6151
R2671 B.n998 B.n997 10.6151
R2672 B.n999 B.n998 10.6151
R2673 B.n1001 B.n999 10.6151
R2674 B.n1002 B.n1001 10.6151
R2675 B.n1003 B.n1002 10.6151
R2676 B.n1004 B.n1003 10.6151
R2677 B.n1006 B.n1004 10.6151
R2678 B.n1007 B.n1006 10.6151
R2679 B.n1008 B.n1007 10.6151
R2680 B.n1009 B.n1008 10.6151
R2681 B.n1011 B.n1009 10.6151
R2682 B.n1012 B.n1011 10.6151
R2683 B.n1013 B.n1012 10.6151
R2684 B.n1014 B.n1013 10.6151
R2685 B.n1016 B.n1014 10.6151
R2686 B.n1017 B.n1016 10.6151
R2687 B.n1018 B.n1017 10.6151
R2688 B.n1019 B.n1018 10.6151
R2689 B.n1021 B.n1019 10.6151
R2690 B.n1022 B.n1021 10.6151
R2691 B.n1023 B.n1022 10.6151
R2692 B.n1024 B.n1023 10.6151
R2693 B.n1026 B.n1024 10.6151
R2694 B.n1027 B.n1026 10.6151
R2695 B.n1028 B.n1027 10.6151
R2696 B.n1029 B.n1028 10.6151
R2697 B.n1031 B.n1029 10.6151
R2698 B.n1032 B.n1031 10.6151
R2699 B.n1033 B.n1032 10.6151
R2700 B.n1034 B.n1033 10.6151
R2701 B.n1036 B.n1034 10.6151
R2702 B.n1037 B.n1036 10.6151
R2703 B.n1038 B.n1037 10.6151
R2704 B.n1039 B.n1038 10.6151
R2705 B.n1041 B.n1039 10.6151
R2706 B.n1042 B.n1041 10.6151
R2707 B.n1043 B.n1042 10.6151
R2708 B.n1044 B.n1043 10.6151
R2709 B.n1046 B.n1044 10.6151
R2710 B.n1047 B.n1046 10.6151
R2711 B.n1048 B.n1047 10.6151
R2712 B.n1194 B.n1 10.6151
R2713 B.n1194 B.n1193 10.6151
R2714 B.n1193 B.n1192 10.6151
R2715 B.n1192 B.n10 10.6151
R2716 B.n1186 B.n10 10.6151
R2717 B.n1186 B.n1185 10.6151
R2718 B.n1185 B.n1184 10.6151
R2719 B.n1184 B.n17 10.6151
R2720 B.n1178 B.n17 10.6151
R2721 B.n1178 B.n1177 10.6151
R2722 B.n1177 B.n1176 10.6151
R2723 B.n1176 B.n25 10.6151
R2724 B.n1170 B.n25 10.6151
R2725 B.n1170 B.n1169 10.6151
R2726 B.n1169 B.n1168 10.6151
R2727 B.n1168 B.n32 10.6151
R2728 B.n1162 B.n32 10.6151
R2729 B.n1162 B.n1161 10.6151
R2730 B.n1161 B.n1160 10.6151
R2731 B.n1160 B.n39 10.6151
R2732 B.n1154 B.n39 10.6151
R2733 B.n1154 B.n1153 10.6151
R2734 B.n1153 B.n1152 10.6151
R2735 B.n1152 B.n46 10.6151
R2736 B.n1146 B.n46 10.6151
R2737 B.n1146 B.n1145 10.6151
R2738 B.n1145 B.n1144 10.6151
R2739 B.n1144 B.n53 10.6151
R2740 B.n1138 B.n53 10.6151
R2741 B.n1138 B.n1137 10.6151
R2742 B.n1137 B.n1136 10.6151
R2743 B.n1136 B.n60 10.6151
R2744 B.n1130 B.n60 10.6151
R2745 B.n1130 B.n1129 10.6151
R2746 B.n1129 B.n1128 10.6151
R2747 B.n1128 B.n67 10.6151
R2748 B.n1122 B.n67 10.6151
R2749 B.n1122 B.n1121 10.6151
R2750 B.n1121 B.n1120 10.6151
R2751 B.n1120 B.n74 10.6151
R2752 B.n1114 B.n74 10.6151
R2753 B.n1114 B.n1113 10.6151
R2754 B.n1113 B.n1112 10.6151
R2755 B.n1112 B.n81 10.6151
R2756 B.n1106 B.n81 10.6151
R2757 B.n1106 B.n1105 10.6151
R2758 B.n1105 B.n1104 10.6151
R2759 B.n1104 B.n88 10.6151
R2760 B.n1098 B.n88 10.6151
R2761 B.n1098 B.n1097 10.6151
R2762 B.n1097 B.n1096 10.6151
R2763 B.n1096 B.n94 10.6151
R2764 B.n1090 B.n94 10.6151
R2765 B.n1090 B.n1089 10.6151
R2766 B.n1089 B.n1088 10.6151
R2767 B.n1088 B.n102 10.6151
R2768 B.n1082 B.n102 10.6151
R2769 B.n1082 B.n1081 10.6151
R2770 B.n1081 B.n1080 10.6151
R2771 B.n1080 B.n109 10.6151
R2772 B.n1074 B.n109 10.6151
R2773 B.n1074 B.n1073 10.6151
R2774 B.n1073 B.n1072 10.6151
R2775 B.n1072 B.n116 10.6151
R2776 B.n1066 B.n116 10.6151
R2777 B.n1066 B.n1065 10.6151
R2778 B.n1065 B.n1064 10.6151
R2779 B.n1064 B.n123 10.6151
R2780 B.n1058 B.n123 10.6151
R2781 B.n1058 B.n1057 10.6151
R2782 B.n1057 B.n1056 10.6151
R2783 B.n1056 B.n130 10.6151
R2784 B.n187 B.n186 10.6151
R2785 B.n190 B.n187 10.6151
R2786 B.n191 B.n190 10.6151
R2787 B.n194 B.n191 10.6151
R2788 B.n195 B.n194 10.6151
R2789 B.n198 B.n195 10.6151
R2790 B.n199 B.n198 10.6151
R2791 B.n202 B.n199 10.6151
R2792 B.n203 B.n202 10.6151
R2793 B.n206 B.n203 10.6151
R2794 B.n207 B.n206 10.6151
R2795 B.n210 B.n207 10.6151
R2796 B.n211 B.n210 10.6151
R2797 B.n214 B.n211 10.6151
R2798 B.n215 B.n214 10.6151
R2799 B.n218 B.n215 10.6151
R2800 B.n219 B.n218 10.6151
R2801 B.n222 B.n219 10.6151
R2802 B.n223 B.n222 10.6151
R2803 B.n226 B.n223 10.6151
R2804 B.n227 B.n226 10.6151
R2805 B.n230 B.n227 10.6151
R2806 B.n231 B.n230 10.6151
R2807 B.n234 B.n231 10.6151
R2808 B.n235 B.n234 10.6151
R2809 B.n238 B.n235 10.6151
R2810 B.n239 B.n238 10.6151
R2811 B.n242 B.n239 10.6151
R2812 B.n243 B.n242 10.6151
R2813 B.n246 B.n243 10.6151
R2814 B.n247 B.n246 10.6151
R2815 B.n250 B.n247 10.6151
R2816 B.n251 B.n250 10.6151
R2817 B.n254 B.n251 10.6151
R2818 B.n255 B.n254 10.6151
R2819 B.n258 B.n255 10.6151
R2820 B.n259 B.n258 10.6151
R2821 B.n262 B.n259 10.6151
R2822 B.n263 B.n262 10.6151
R2823 B.n267 B.n266 10.6151
R2824 B.n270 B.n267 10.6151
R2825 B.n271 B.n270 10.6151
R2826 B.n274 B.n271 10.6151
R2827 B.n275 B.n274 10.6151
R2828 B.n278 B.n275 10.6151
R2829 B.n279 B.n278 10.6151
R2830 B.n282 B.n279 10.6151
R2831 B.n283 B.n282 10.6151
R2832 B.n287 B.n286 10.6151
R2833 B.n290 B.n287 10.6151
R2834 B.n291 B.n290 10.6151
R2835 B.n294 B.n291 10.6151
R2836 B.n295 B.n294 10.6151
R2837 B.n298 B.n295 10.6151
R2838 B.n299 B.n298 10.6151
R2839 B.n302 B.n299 10.6151
R2840 B.n303 B.n302 10.6151
R2841 B.n306 B.n303 10.6151
R2842 B.n307 B.n306 10.6151
R2843 B.n310 B.n307 10.6151
R2844 B.n311 B.n310 10.6151
R2845 B.n314 B.n311 10.6151
R2846 B.n315 B.n314 10.6151
R2847 B.n318 B.n315 10.6151
R2848 B.n319 B.n318 10.6151
R2849 B.n322 B.n319 10.6151
R2850 B.n323 B.n322 10.6151
R2851 B.n326 B.n323 10.6151
R2852 B.n327 B.n326 10.6151
R2853 B.n330 B.n327 10.6151
R2854 B.n331 B.n330 10.6151
R2855 B.n334 B.n331 10.6151
R2856 B.n335 B.n334 10.6151
R2857 B.n338 B.n335 10.6151
R2858 B.n339 B.n338 10.6151
R2859 B.n342 B.n339 10.6151
R2860 B.n343 B.n342 10.6151
R2861 B.n346 B.n343 10.6151
R2862 B.n347 B.n346 10.6151
R2863 B.n350 B.n347 10.6151
R2864 B.n351 B.n350 10.6151
R2865 B.n354 B.n351 10.6151
R2866 B.n355 B.n354 10.6151
R2867 B.n358 B.n355 10.6151
R2868 B.n360 B.n358 10.6151
R2869 B.n361 B.n360 10.6151
R2870 B.n1049 B.n361 10.6151
R2871 B.n653 B.n652 9.36635
R2872 B.n631 B.n630 9.36635
R2873 B.n263 B.n184 9.36635
R2874 B.n286 B.n181 9.36635
R2875 B.n1202 B.n0 8.11757
R2876 B.n1202 B.n1 8.11757
R2877 B.n652 B.n651 1.24928
R2878 B.n632 B.n631 1.24928
R2879 B.n266 B.n184 1.24928
R2880 B.n283 B.n181 1.24928
R2881 VN.n98 VN.n97 161.3
R2882 VN.n96 VN.n51 161.3
R2883 VN.n95 VN.n94 161.3
R2884 VN.n93 VN.n52 161.3
R2885 VN.n92 VN.n91 161.3
R2886 VN.n90 VN.n53 161.3
R2887 VN.n89 VN.n88 161.3
R2888 VN.n87 VN.n54 161.3
R2889 VN.n86 VN.n85 161.3
R2890 VN.n84 VN.n55 161.3
R2891 VN.n83 VN.n82 161.3
R2892 VN.n81 VN.n57 161.3
R2893 VN.n80 VN.n79 161.3
R2894 VN.n78 VN.n58 161.3
R2895 VN.n77 VN.n76 161.3
R2896 VN.n75 VN.n74 161.3
R2897 VN.n73 VN.n60 161.3
R2898 VN.n72 VN.n71 161.3
R2899 VN.n70 VN.n61 161.3
R2900 VN.n69 VN.n68 161.3
R2901 VN.n67 VN.n62 161.3
R2902 VN.n66 VN.n65 161.3
R2903 VN.n48 VN.n47 161.3
R2904 VN.n46 VN.n1 161.3
R2905 VN.n45 VN.n44 161.3
R2906 VN.n43 VN.n2 161.3
R2907 VN.n42 VN.n41 161.3
R2908 VN.n40 VN.n3 161.3
R2909 VN.n39 VN.n38 161.3
R2910 VN.n37 VN.n4 161.3
R2911 VN.n36 VN.n35 161.3
R2912 VN.n33 VN.n5 161.3
R2913 VN.n32 VN.n31 161.3
R2914 VN.n30 VN.n6 161.3
R2915 VN.n29 VN.n28 161.3
R2916 VN.n27 VN.n7 161.3
R2917 VN.n26 VN.n25 161.3
R2918 VN.n24 VN.n23 161.3
R2919 VN.n22 VN.n9 161.3
R2920 VN.n21 VN.n20 161.3
R2921 VN.n19 VN.n10 161.3
R2922 VN.n18 VN.n17 161.3
R2923 VN.n16 VN.n11 161.3
R2924 VN.n15 VN.n14 161.3
R2925 VN.n64 VN.t6 115.392
R2926 VN.n13 VN.t5 115.392
R2927 VN.n12 VN.t4 82.1111
R2928 VN.n8 VN.t8 82.1111
R2929 VN.n34 VN.t7 82.1111
R2930 VN.n0 VN.t9 82.1111
R2931 VN.n63 VN.t2 82.1111
R2932 VN.n59 VN.t1 82.1111
R2933 VN.n56 VN.t3 82.1111
R2934 VN.n50 VN.t0 82.1111
R2935 VN.n49 VN.n0 80.7699
R2936 VN.n99 VN.n50 80.7699
R2937 VN VN.n99 57.2859
R2938 VN.n41 VN.n2 56.5193
R2939 VN.n91 VN.n52 56.5193
R2940 VN.n13 VN.n12 51.5827
R2941 VN.n64 VN.n63 51.5827
R2942 VN.n17 VN.n10 51.1773
R2943 VN.n32 VN.n6 51.1773
R2944 VN.n68 VN.n61 51.1773
R2945 VN.n83 VN.n57 51.1773
R2946 VN.n21 VN.n10 29.8095
R2947 VN.n28 VN.n6 29.8095
R2948 VN.n72 VN.n61 29.8095
R2949 VN.n79 VN.n57 29.8095
R2950 VN.n16 VN.n15 24.4675
R2951 VN.n17 VN.n16 24.4675
R2952 VN.n22 VN.n21 24.4675
R2953 VN.n23 VN.n22 24.4675
R2954 VN.n27 VN.n26 24.4675
R2955 VN.n28 VN.n27 24.4675
R2956 VN.n33 VN.n32 24.4675
R2957 VN.n35 VN.n33 24.4675
R2958 VN.n39 VN.n4 24.4675
R2959 VN.n40 VN.n39 24.4675
R2960 VN.n41 VN.n40 24.4675
R2961 VN.n45 VN.n2 24.4675
R2962 VN.n46 VN.n45 24.4675
R2963 VN.n47 VN.n46 24.4675
R2964 VN.n68 VN.n67 24.4675
R2965 VN.n67 VN.n66 24.4675
R2966 VN.n79 VN.n78 24.4675
R2967 VN.n78 VN.n77 24.4675
R2968 VN.n74 VN.n73 24.4675
R2969 VN.n73 VN.n72 24.4675
R2970 VN.n91 VN.n90 24.4675
R2971 VN.n90 VN.n89 24.4675
R2972 VN.n89 VN.n54 24.4675
R2973 VN.n85 VN.n84 24.4675
R2974 VN.n84 VN.n83 24.4675
R2975 VN.n97 VN.n96 24.4675
R2976 VN.n96 VN.n95 24.4675
R2977 VN.n95 VN.n52 24.4675
R2978 VN.n15 VN.n12 22.9995
R2979 VN.n35 VN.n34 22.9995
R2980 VN.n66 VN.n63 22.9995
R2981 VN.n85 VN.n56 22.9995
R2982 VN.n23 VN.n8 12.234
R2983 VN.n26 VN.n8 12.234
R2984 VN.n77 VN.n59 12.234
R2985 VN.n74 VN.n59 12.234
R2986 VN.n47 VN.n0 9.29796
R2987 VN.n97 VN.n50 9.29796
R2988 VN.n65 VN.n64 3.17993
R2989 VN.n14 VN.n13 3.17993
R2990 VN.n34 VN.n4 1.46852
R2991 VN.n56 VN.n54 1.46852
R2992 VN.n99 VN.n98 0.354971
R2993 VN.n49 VN.n48 0.354971
R2994 VN VN.n49 0.26696
R2995 VN.n98 VN.n51 0.189894
R2996 VN.n94 VN.n51 0.189894
R2997 VN.n94 VN.n93 0.189894
R2998 VN.n93 VN.n92 0.189894
R2999 VN.n92 VN.n53 0.189894
R3000 VN.n88 VN.n53 0.189894
R3001 VN.n88 VN.n87 0.189894
R3002 VN.n87 VN.n86 0.189894
R3003 VN.n86 VN.n55 0.189894
R3004 VN.n82 VN.n55 0.189894
R3005 VN.n82 VN.n81 0.189894
R3006 VN.n81 VN.n80 0.189894
R3007 VN.n80 VN.n58 0.189894
R3008 VN.n76 VN.n58 0.189894
R3009 VN.n76 VN.n75 0.189894
R3010 VN.n75 VN.n60 0.189894
R3011 VN.n71 VN.n60 0.189894
R3012 VN.n71 VN.n70 0.189894
R3013 VN.n70 VN.n69 0.189894
R3014 VN.n69 VN.n62 0.189894
R3015 VN.n65 VN.n62 0.189894
R3016 VN.n14 VN.n11 0.189894
R3017 VN.n18 VN.n11 0.189894
R3018 VN.n19 VN.n18 0.189894
R3019 VN.n20 VN.n19 0.189894
R3020 VN.n20 VN.n9 0.189894
R3021 VN.n24 VN.n9 0.189894
R3022 VN.n25 VN.n24 0.189894
R3023 VN.n25 VN.n7 0.189894
R3024 VN.n29 VN.n7 0.189894
R3025 VN.n30 VN.n29 0.189894
R3026 VN.n31 VN.n30 0.189894
R3027 VN.n31 VN.n5 0.189894
R3028 VN.n36 VN.n5 0.189894
R3029 VN.n37 VN.n36 0.189894
R3030 VN.n38 VN.n37 0.189894
R3031 VN.n38 VN.n3 0.189894
R3032 VN.n42 VN.n3 0.189894
R3033 VN.n43 VN.n42 0.189894
R3034 VN.n44 VN.n43 0.189894
R3035 VN.n44 VN.n1 0.189894
R3036 VN.n48 VN.n1 0.189894
R3037 VDD2.n121 VDD2.n65 289.615
R3038 VDD2.n56 VDD2.n0 289.615
R3039 VDD2.n122 VDD2.n121 185
R3040 VDD2.n120 VDD2.n119 185
R3041 VDD2.n69 VDD2.n68 185
R3042 VDD2.n114 VDD2.n113 185
R3043 VDD2.n112 VDD2.n111 185
R3044 VDD2.n73 VDD2.n72 185
R3045 VDD2.n77 VDD2.n75 185
R3046 VDD2.n106 VDD2.n105 185
R3047 VDD2.n104 VDD2.n103 185
R3048 VDD2.n79 VDD2.n78 185
R3049 VDD2.n98 VDD2.n97 185
R3050 VDD2.n96 VDD2.n95 185
R3051 VDD2.n83 VDD2.n82 185
R3052 VDD2.n90 VDD2.n89 185
R3053 VDD2.n88 VDD2.n87 185
R3054 VDD2.n21 VDD2.n20 185
R3055 VDD2.n23 VDD2.n22 185
R3056 VDD2.n16 VDD2.n15 185
R3057 VDD2.n29 VDD2.n28 185
R3058 VDD2.n31 VDD2.n30 185
R3059 VDD2.n12 VDD2.n11 185
R3060 VDD2.n38 VDD2.n37 185
R3061 VDD2.n39 VDD2.n10 185
R3062 VDD2.n41 VDD2.n40 185
R3063 VDD2.n8 VDD2.n7 185
R3064 VDD2.n47 VDD2.n46 185
R3065 VDD2.n49 VDD2.n48 185
R3066 VDD2.n4 VDD2.n3 185
R3067 VDD2.n55 VDD2.n54 185
R3068 VDD2.n57 VDD2.n56 185
R3069 VDD2.n86 VDD2.t9 149.524
R3070 VDD2.n19 VDD2.t4 149.524
R3071 VDD2.n121 VDD2.n120 104.615
R3072 VDD2.n120 VDD2.n68 104.615
R3073 VDD2.n113 VDD2.n68 104.615
R3074 VDD2.n113 VDD2.n112 104.615
R3075 VDD2.n112 VDD2.n72 104.615
R3076 VDD2.n77 VDD2.n72 104.615
R3077 VDD2.n105 VDD2.n77 104.615
R3078 VDD2.n105 VDD2.n104 104.615
R3079 VDD2.n104 VDD2.n78 104.615
R3080 VDD2.n97 VDD2.n78 104.615
R3081 VDD2.n97 VDD2.n96 104.615
R3082 VDD2.n96 VDD2.n82 104.615
R3083 VDD2.n89 VDD2.n82 104.615
R3084 VDD2.n89 VDD2.n88 104.615
R3085 VDD2.n22 VDD2.n21 104.615
R3086 VDD2.n22 VDD2.n15 104.615
R3087 VDD2.n29 VDD2.n15 104.615
R3088 VDD2.n30 VDD2.n29 104.615
R3089 VDD2.n30 VDD2.n11 104.615
R3090 VDD2.n38 VDD2.n11 104.615
R3091 VDD2.n39 VDD2.n38 104.615
R3092 VDD2.n40 VDD2.n39 104.615
R3093 VDD2.n40 VDD2.n7 104.615
R3094 VDD2.n47 VDD2.n7 104.615
R3095 VDD2.n48 VDD2.n47 104.615
R3096 VDD2.n48 VDD2.n3 104.615
R3097 VDD2.n55 VDD2.n3 104.615
R3098 VDD2.n56 VDD2.n55 104.615
R3099 VDD2.n64 VDD2.n63 67.3487
R3100 VDD2 VDD2.n129 67.3458
R3101 VDD2.n128 VDD2.n127 64.999
R3102 VDD2.n62 VDD2.n61 64.9988
R3103 VDD2.n62 VDD2.n60 54.9801
R3104 VDD2.n88 VDD2.t9 52.3082
R3105 VDD2.n21 VDD2.t4 52.3082
R3106 VDD2.n126 VDD2.n125 51.7732
R3107 VDD2.n126 VDD2.n64 48.905
R3108 VDD2.n75 VDD2.n73 13.1884
R3109 VDD2.n41 VDD2.n8 13.1884
R3110 VDD2.n111 VDD2.n110 12.8005
R3111 VDD2.n107 VDD2.n106 12.8005
R3112 VDD2.n42 VDD2.n10 12.8005
R3113 VDD2.n46 VDD2.n45 12.8005
R3114 VDD2.n114 VDD2.n71 12.0247
R3115 VDD2.n103 VDD2.n76 12.0247
R3116 VDD2.n37 VDD2.n36 12.0247
R3117 VDD2.n49 VDD2.n6 12.0247
R3118 VDD2.n115 VDD2.n69 11.249
R3119 VDD2.n102 VDD2.n79 11.249
R3120 VDD2.n35 VDD2.n12 11.249
R3121 VDD2.n50 VDD2.n4 11.249
R3122 VDD2.n119 VDD2.n118 10.4732
R3123 VDD2.n99 VDD2.n98 10.4732
R3124 VDD2.n32 VDD2.n31 10.4732
R3125 VDD2.n54 VDD2.n53 10.4732
R3126 VDD2.n87 VDD2.n86 10.2747
R3127 VDD2.n20 VDD2.n19 10.2747
R3128 VDD2.n122 VDD2.n67 9.69747
R3129 VDD2.n95 VDD2.n81 9.69747
R3130 VDD2.n28 VDD2.n14 9.69747
R3131 VDD2.n57 VDD2.n2 9.69747
R3132 VDD2.n125 VDD2.n124 9.45567
R3133 VDD2.n60 VDD2.n59 9.45567
R3134 VDD2.n85 VDD2.n84 9.3005
R3135 VDD2.n92 VDD2.n91 9.3005
R3136 VDD2.n94 VDD2.n93 9.3005
R3137 VDD2.n81 VDD2.n80 9.3005
R3138 VDD2.n100 VDD2.n99 9.3005
R3139 VDD2.n102 VDD2.n101 9.3005
R3140 VDD2.n76 VDD2.n74 9.3005
R3141 VDD2.n108 VDD2.n107 9.3005
R3142 VDD2.n124 VDD2.n123 9.3005
R3143 VDD2.n67 VDD2.n66 9.3005
R3144 VDD2.n118 VDD2.n117 9.3005
R3145 VDD2.n116 VDD2.n115 9.3005
R3146 VDD2.n71 VDD2.n70 9.3005
R3147 VDD2.n110 VDD2.n109 9.3005
R3148 VDD2.n59 VDD2.n58 9.3005
R3149 VDD2.n2 VDD2.n1 9.3005
R3150 VDD2.n53 VDD2.n52 9.3005
R3151 VDD2.n51 VDD2.n50 9.3005
R3152 VDD2.n6 VDD2.n5 9.3005
R3153 VDD2.n45 VDD2.n44 9.3005
R3154 VDD2.n18 VDD2.n17 9.3005
R3155 VDD2.n25 VDD2.n24 9.3005
R3156 VDD2.n27 VDD2.n26 9.3005
R3157 VDD2.n14 VDD2.n13 9.3005
R3158 VDD2.n33 VDD2.n32 9.3005
R3159 VDD2.n35 VDD2.n34 9.3005
R3160 VDD2.n36 VDD2.n9 9.3005
R3161 VDD2.n43 VDD2.n42 9.3005
R3162 VDD2.n123 VDD2.n65 8.92171
R3163 VDD2.n94 VDD2.n83 8.92171
R3164 VDD2.n27 VDD2.n16 8.92171
R3165 VDD2.n58 VDD2.n0 8.92171
R3166 VDD2.n91 VDD2.n90 8.14595
R3167 VDD2.n24 VDD2.n23 8.14595
R3168 VDD2.n87 VDD2.n85 7.3702
R3169 VDD2.n20 VDD2.n18 7.3702
R3170 VDD2.n90 VDD2.n85 5.81868
R3171 VDD2.n23 VDD2.n18 5.81868
R3172 VDD2.n125 VDD2.n65 5.04292
R3173 VDD2.n91 VDD2.n83 5.04292
R3174 VDD2.n24 VDD2.n16 5.04292
R3175 VDD2.n60 VDD2.n0 5.04292
R3176 VDD2.n123 VDD2.n122 4.26717
R3177 VDD2.n95 VDD2.n94 4.26717
R3178 VDD2.n28 VDD2.n27 4.26717
R3179 VDD2.n58 VDD2.n57 4.26717
R3180 VDD2.n119 VDD2.n67 3.49141
R3181 VDD2.n98 VDD2.n81 3.49141
R3182 VDD2.n31 VDD2.n14 3.49141
R3183 VDD2.n54 VDD2.n2 3.49141
R3184 VDD2.n128 VDD2.n126 3.2074
R3185 VDD2.n86 VDD2.n84 2.84303
R3186 VDD2.n19 VDD2.n17 2.84303
R3187 VDD2.n118 VDD2.n69 2.71565
R3188 VDD2.n99 VDD2.n79 2.71565
R3189 VDD2.n32 VDD2.n12 2.71565
R3190 VDD2.n53 VDD2.n4 2.71565
R3191 VDD2.n115 VDD2.n114 1.93989
R3192 VDD2.n103 VDD2.n102 1.93989
R3193 VDD2.n37 VDD2.n35 1.93989
R3194 VDD2.n50 VDD2.n49 1.93989
R3195 VDD2.n129 VDD2.t7 1.71479
R3196 VDD2.n129 VDD2.t3 1.71479
R3197 VDD2.n127 VDD2.t6 1.71479
R3198 VDD2.n127 VDD2.t8 1.71479
R3199 VDD2.n63 VDD2.t2 1.71479
R3200 VDD2.n63 VDD2.t0 1.71479
R3201 VDD2.n61 VDD2.t5 1.71479
R3202 VDD2.n61 VDD2.t1 1.71479
R3203 VDD2.n111 VDD2.n71 1.16414
R3204 VDD2.n106 VDD2.n76 1.16414
R3205 VDD2.n36 VDD2.n10 1.16414
R3206 VDD2.n46 VDD2.n6 1.16414
R3207 VDD2 VDD2.n128 0.860414
R3208 VDD2.n64 VDD2.n62 0.746878
R3209 VDD2.n110 VDD2.n73 0.388379
R3210 VDD2.n107 VDD2.n75 0.388379
R3211 VDD2.n42 VDD2.n41 0.388379
R3212 VDD2.n45 VDD2.n8 0.388379
R3213 VDD2.n124 VDD2.n66 0.155672
R3214 VDD2.n117 VDD2.n66 0.155672
R3215 VDD2.n117 VDD2.n116 0.155672
R3216 VDD2.n116 VDD2.n70 0.155672
R3217 VDD2.n109 VDD2.n70 0.155672
R3218 VDD2.n109 VDD2.n108 0.155672
R3219 VDD2.n108 VDD2.n74 0.155672
R3220 VDD2.n101 VDD2.n74 0.155672
R3221 VDD2.n101 VDD2.n100 0.155672
R3222 VDD2.n100 VDD2.n80 0.155672
R3223 VDD2.n93 VDD2.n80 0.155672
R3224 VDD2.n93 VDD2.n92 0.155672
R3225 VDD2.n92 VDD2.n84 0.155672
R3226 VDD2.n25 VDD2.n17 0.155672
R3227 VDD2.n26 VDD2.n25 0.155672
R3228 VDD2.n26 VDD2.n13 0.155672
R3229 VDD2.n33 VDD2.n13 0.155672
R3230 VDD2.n34 VDD2.n33 0.155672
R3231 VDD2.n34 VDD2.n9 0.155672
R3232 VDD2.n43 VDD2.n9 0.155672
R3233 VDD2.n44 VDD2.n43 0.155672
R3234 VDD2.n44 VDD2.n5 0.155672
R3235 VDD2.n51 VDD2.n5 0.155672
R3236 VDD2.n52 VDD2.n51 0.155672
R3237 VDD2.n52 VDD2.n1 0.155672
R3238 VDD2.n59 VDD2.n1 0.155672
C0 VDD1 VN 0.155233f
C1 VDD2 VN 10.7803f
C2 VDD1 VTAIL 10.5498f
C3 VDD1 VP 11.305599f
C4 VDD2 VTAIL 10.6068f
C5 VDD2 VP 0.684413f
C6 VN VTAIL 11.782299f
C7 VP VN 9.48308f
C8 VP VTAIL 11.7966f
C9 VDD1 VDD2 2.68943f
C10 VDD2 B 8.058657f
C11 VDD1 B 8.024604f
C12 VTAIL B 8.631427f
C13 VN B 21.8829f
C14 VP B 20.46065f
C15 VDD2.n0 B 0.036627f
C16 VDD2.n1 B 0.024751f
C17 VDD2.n2 B 0.0133f
C18 VDD2.n3 B 0.031437f
C19 VDD2.n4 B 0.014082f
C20 VDD2.n5 B 0.024751f
C21 VDD2.n6 B 0.0133f
C22 VDD2.n7 B 0.031437f
C23 VDD2.n8 B 0.013691f
C24 VDD2.n9 B 0.024751f
C25 VDD2.n10 B 0.014082f
C26 VDD2.n11 B 0.031437f
C27 VDD2.n12 B 0.014082f
C28 VDD2.n13 B 0.024751f
C29 VDD2.n14 B 0.0133f
C30 VDD2.n15 B 0.031437f
C31 VDD2.n16 B 0.014082f
C32 VDD2.n17 B 1.19911f
C33 VDD2.n18 B 0.0133f
C34 VDD2.t4 B 0.053035f
C35 VDD2.n19 B 0.174178f
C36 VDD2.n20 B 0.022223f
C37 VDD2.n21 B 0.023578f
C38 VDD2.n22 B 0.031437f
C39 VDD2.n23 B 0.014082f
C40 VDD2.n24 B 0.0133f
C41 VDD2.n25 B 0.024751f
C42 VDD2.n26 B 0.024751f
C43 VDD2.n27 B 0.0133f
C44 VDD2.n28 B 0.014082f
C45 VDD2.n29 B 0.031437f
C46 VDD2.n30 B 0.031437f
C47 VDD2.n31 B 0.014082f
C48 VDD2.n32 B 0.0133f
C49 VDD2.n33 B 0.024751f
C50 VDD2.n34 B 0.024751f
C51 VDD2.n35 B 0.0133f
C52 VDD2.n36 B 0.0133f
C53 VDD2.n37 B 0.014082f
C54 VDD2.n38 B 0.031437f
C55 VDD2.n39 B 0.031437f
C56 VDD2.n40 B 0.031437f
C57 VDD2.n41 B 0.013691f
C58 VDD2.n42 B 0.0133f
C59 VDD2.n43 B 0.024751f
C60 VDD2.n44 B 0.024751f
C61 VDD2.n45 B 0.0133f
C62 VDD2.n46 B 0.014082f
C63 VDD2.n47 B 0.031437f
C64 VDD2.n48 B 0.031437f
C65 VDD2.n49 B 0.014082f
C66 VDD2.n50 B 0.0133f
C67 VDD2.n51 B 0.024751f
C68 VDD2.n52 B 0.024751f
C69 VDD2.n53 B 0.0133f
C70 VDD2.n54 B 0.014082f
C71 VDD2.n55 B 0.031437f
C72 VDD2.n56 B 0.071304f
C73 VDD2.n57 B 0.014082f
C74 VDD2.n58 B 0.0133f
C75 VDD2.n59 B 0.062283f
C76 VDD2.n60 B 0.075303f
C77 VDD2.t5 B 0.225908f
C78 VDD2.t1 B 0.225908f
C79 VDD2.n61 B 2.01084f
C80 VDD2.n62 B 0.806203f
C81 VDD2.t2 B 0.225908f
C82 VDD2.t0 B 0.225908f
C83 VDD2.n63 B 2.03369f
C84 VDD2.n64 B 3.25487f
C85 VDD2.n65 B 0.036627f
C86 VDD2.n66 B 0.024751f
C87 VDD2.n67 B 0.0133f
C88 VDD2.n68 B 0.031437f
C89 VDD2.n69 B 0.014082f
C90 VDD2.n70 B 0.024751f
C91 VDD2.n71 B 0.0133f
C92 VDD2.n72 B 0.031437f
C93 VDD2.n73 B 0.013691f
C94 VDD2.n74 B 0.024751f
C95 VDD2.n75 B 0.013691f
C96 VDD2.n76 B 0.0133f
C97 VDD2.n77 B 0.031437f
C98 VDD2.n78 B 0.031437f
C99 VDD2.n79 B 0.014082f
C100 VDD2.n80 B 0.024751f
C101 VDD2.n81 B 0.0133f
C102 VDD2.n82 B 0.031437f
C103 VDD2.n83 B 0.014082f
C104 VDD2.n84 B 1.19911f
C105 VDD2.n85 B 0.0133f
C106 VDD2.t9 B 0.053035f
C107 VDD2.n86 B 0.174178f
C108 VDD2.n87 B 0.022223f
C109 VDD2.n88 B 0.023578f
C110 VDD2.n89 B 0.031437f
C111 VDD2.n90 B 0.014082f
C112 VDD2.n91 B 0.0133f
C113 VDD2.n92 B 0.024751f
C114 VDD2.n93 B 0.024751f
C115 VDD2.n94 B 0.0133f
C116 VDD2.n95 B 0.014082f
C117 VDD2.n96 B 0.031437f
C118 VDD2.n97 B 0.031437f
C119 VDD2.n98 B 0.014082f
C120 VDD2.n99 B 0.0133f
C121 VDD2.n100 B 0.024751f
C122 VDD2.n101 B 0.024751f
C123 VDD2.n102 B 0.0133f
C124 VDD2.n103 B 0.014082f
C125 VDD2.n104 B 0.031437f
C126 VDD2.n105 B 0.031437f
C127 VDD2.n106 B 0.014082f
C128 VDD2.n107 B 0.0133f
C129 VDD2.n108 B 0.024751f
C130 VDD2.n109 B 0.024751f
C131 VDD2.n110 B 0.0133f
C132 VDD2.n111 B 0.014082f
C133 VDD2.n112 B 0.031437f
C134 VDD2.n113 B 0.031437f
C135 VDD2.n114 B 0.014082f
C136 VDD2.n115 B 0.0133f
C137 VDD2.n116 B 0.024751f
C138 VDD2.n117 B 0.024751f
C139 VDD2.n118 B 0.0133f
C140 VDD2.n119 B 0.014082f
C141 VDD2.n120 B 0.031437f
C142 VDD2.n121 B 0.071304f
C143 VDD2.n122 B 0.014082f
C144 VDD2.n123 B 0.0133f
C145 VDD2.n124 B 0.062283f
C146 VDD2.n125 B 0.057435f
C147 VDD2.n126 B 3.13512f
C148 VDD2.t6 B 0.225908f
C149 VDD2.t8 B 0.225908f
C150 VDD2.n127 B 2.01084f
C151 VDD2.n128 B 0.526022f
C152 VDD2.t7 B 0.225908f
C153 VDD2.t3 B 0.225908f
C154 VDD2.n129 B 2.03365f
C155 VN.t9 B 1.93907f
C156 VN.n0 B 0.749744f
C157 VN.n1 B 0.018197f
C158 VN.n2 B 0.022507f
C159 VN.n3 B 0.018197f
C160 VN.n4 B 0.018175f
C161 VN.n5 B 0.018197f
C162 VN.n6 B 0.01775f
C163 VN.n7 B 0.018197f
C164 VN.t8 B 1.93907f
C165 VN.n8 B 0.682307f
C166 VN.n9 B 0.018197f
C167 VN.n10 B 0.01775f
C168 VN.n11 B 0.018197f
C169 VN.t4 B 1.93907f
C170 VN.n12 B 0.752684f
C171 VN.t5 B 2.17436f
C172 VN.n13 B 0.710254f
C173 VN.n14 B 0.222681f
C174 VN.n15 B 0.032909f
C175 VN.n16 B 0.033914f
C176 VN.n17 B 0.033038f
C177 VN.n18 B 0.018197f
C178 VN.n19 B 0.018197f
C179 VN.n20 B 0.018197f
C180 VN.n21 B 0.036253f
C181 VN.n22 B 0.033914f
C182 VN.n23 B 0.025542f
C183 VN.n24 B 0.018197f
C184 VN.n25 B 0.018197f
C185 VN.n26 B 0.025542f
C186 VN.n27 B 0.033914f
C187 VN.n28 B 0.036253f
C188 VN.n29 B 0.018197f
C189 VN.n30 B 0.018197f
C190 VN.n31 B 0.018197f
C191 VN.n32 B 0.033038f
C192 VN.n33 B 0.033914f
C193 VN.t7 B 1.93907f
C194 VN.n34 B 0.682307f
C195 VN.n35 B 0.032909f
C196 VN.n36 B 0.018197f
C197 VN.n37 B 0.018197f
C198 VN.n38 B 0.018197f
C199 VN.n39 B 0.033914f
C200 VN.n40 B 0.033914f
C201 VN.n41 B 0.03062f
C202 VN.n42 B 0.018197f
C203 VN.n43 B 0.018197f
C204 VN.n44 B 0.018197f
C205 VN.n45 B 0.033914f
C206 VN.n46 B 0.033914f
C207 VN.n47 B 0.023533f
C208 VN.n48 B 0.029369f
C209 VN.n49 B 0.048354f
C210 VN.t0 B 1.93907f
C211 VN.n50 B 0.749744f
C212 VN.n51 B 0.018197f
C213 VN.n52 B 0.022507f
C214 VN.n53 B 0.018197f
C215 VN.n54 B 0.018175f
C216 VN.n55 B 0.018197f
C217 VN.t3 B 1.93907f
C218 VN.n56 B 0.682307f
C219 VN.n57 B 0.01775f
C220 VN.n58 B 0.018197f
C221 VN.t1 B 1.93907f
C222 VN.n59 B 0.682307f
C223 VN.n60 B 0.018197f
C224 VN.n61 B 0.01775f
C225 VN.n62 B 0.018197f
C226 VN.t2 B 1.93907f
C227 VN.n63 B 0.752684f
C228 VN.t6 B 2.17436f
C229 VN.n64 B 0.710254f
C230 VN.n65 B 0.222681f
C231 VN.n66 B 0.032909f
C232 VN.n67 B 0.033914f
C233 VN.n68 B 0.033038f
C234 VN.n69 B 0.018197f
C235 VN.n70 B 0.018197f
C236 VN.n71 B 0.018197f
C237 VN.n72 B 0.036253f
C238 VN.n73 B 0.033914f
C239 VN.n74 B 0.025542f
C240 VN.n75 B 0.018197f
C241 VN.n76 B 0.018197f
C242 VN.n77 B 0.025542f
C243 VN.n78 B 0.033914f
C244 VN.n79 B 0.036253f
C245 VN.n80 B 0.018197f
C246 VN.n81 B 0.018197f
C247 VN.n82 B 0.018197f
C248 VN.n83 B 0.033038f
C249 VN.n84 B 0.033914f
C250 VN.n85 B 0.032909f
C251 VN.n86 B 0.018197f
C252 VN.n87 B 0.018197f
C253 VN.n88 B 0.018197f
C254 VN.n89 B 0.033914f
C255 VN.n90 B 0.033914f
C256 VN.n91 B 0.03062f
C257 VN.n92 B 0.018197f
C258 VN.n93 B 0.018197f
C259 VN.n94 B 0.018197f
C260 VN.n95 B 0.033914f
C261 VN.n96 B 0.033914f
C262 VN.n97 B 0.023533f
C263 VN.n98 B 0.029369f
C264 VN.n99 B 1.25758f
C265 VTAIL.t2 B 0.234648f
C266 VTAIL.t0 B 0.234648f
C267 VTAIL.n0 B 2.01802f
C268 VTAIL.n1 B 0.620981f
C269 VTAIL.n2 B 0.038044f
C270 VTAIL.n3 B 0.025709f
C271 VTAIL.n4 B 0.013815f
C272 VTAIL.n5 B 0.032653f
C273 VTAIL.n6 B 0.014627f
C274 VTAIL.n7 B 0.025709f
C275 VTAIL.n8 B 0.013815f
C276 VTAIL.n9 B 0.032653f
C277 VTAIL.n10 B 0.014221f
C278 VTAIL.n11 B 0.025709f
C279 VTAIL.n12 B 0.014627f
C280 VTAIL.n13 B 0.032653f
C281 VTAIL.n14 B 0.014627f
C282 VTAIL.n15 B 0.025709f
C283 VTAIL.n16 B 0.013815f
C284 VTAIL.n17 B 0.032653f
C285 VTAIL.n18 B 0.014627f
C286 VTAIL.n19 B 1.2455f
C287 VTAIL.n20 B 0.013815f
C288 VTAIL.t12 B 0.055087f
C289 VTAIL.n21 B 0.180916f
C290 VTAIL.n22 B 0.023083f
C291 VTAIL.n23 B 0.02449f
C292 VTAIL.n24 B 0.032653f
C293 VTAIL.n25 B 0.014627f
C294 VTAIL.n26 B 0.013815f
C295 VTAIL.n27 B 0.025709f
C296 VTAIL.n28 B 0.025709f
C297 VTAIL.n29 B 0.013815f
C298 VTAIL.n30 B 0.014627f
C299 VTAIL.n31 B 0.032653f
C300 VTAIL.n32 B 0.032653f
C301 VTAIL.n33 B 0.014627f
C302 VTAIL.n34 B 0.013815f
C303 VTAIL.n35 B 0.025709f
C304 VTAIL.n36 B 0.025709f
C305 VTAIL.n37 B 0.013815f
C306 VTAIL.n38 B 0.013815f
C307 VTAIL.n39 B 0.014627f
C308 VTAIL.n40 B 0.032653f
C309 VTAIL.n41 B 0.032653f
C310 VTAIL.n42 B 0.032653f
C311 VTAIL.n43 B 0.014221f
C312 VTAIL.n44 B 0.013815f
C313 VTAIL.n45 B 0.025709f
C314 VTAIL.n46 B 0.025709f
C315 VTAIL.n47 B 0.013815f
C316 VTAIL.n48 B 0.014627f
C317 VTAIL.n49 B 0.032653f
C318 VTAIL.n50 B 0.032653f
C319 VTAIL.n51 B 0.014627f
C320 VTAIL.n52 B 0.013815f
C321 VTAIL.n53 B 0.025709f
C322 VTAIL.n54 B 0.025709f
C323 VTAIL.n55 B 0.013815f
C324 VTAIL.n56 B 0.014627f
C325 VTAIL.n57 B 0.032653f
C326 VTAIL.n58 B 0.074063f
C327 VTAIL.n59 B 0.014627f
C328 VTAIL.n60 B 0.013815f
C329 VTAIL.n61 B 0.064693f
C330 VTAIL.n62 B 0.041944f
C331 VTAIL.n63 B 0.462343f
C332 VTAIL.t9 B 0.234648f
C333 VTAIL.t10 B 0.234648f
C334 VTAIL.n64 B 2.01802f
C335 VTAIL.n65 B 0.776483f
C336 VTAIL.t15 B 0.234648f
C337 VTAIL.t8 B 0.234648f
C338 VTAIL.n66 B 2.01802f
C339 VTAIL.n67 B 2.21619f
C340 VTAIL.t6 B 0.234648f
C341 VTAIL.t18 B 0.234648f
C342 VTAIL.n68 B 2.01803f
C343 VTAIL.n69 B 2.21617f
C344 VTAIL.t7 B 0.234648f
C345 VTAIL.t19 B 0.234648f
C346 VTAIL.n70 B 2.01803f
C347 VTAIL.n71 B 0.776472f
C348 VTAIL.n72 B 0.038044f
C349 VTAIL.n73 B 0.025709f
C350 VTAIL.n74 B 0.013815f
C351 VTAIL.n75 B 0.032653f
C352 VTAIL.n76 B 0.014627f
C353 VTAIL.n77 B 0.025709f
C354 VTAIL.n78 B 0.013815f
C355 VTAIL.n79 B 0.032653f
C356 VTAIL.n80 B 0.014221f
C357 VTAIL.n81 B 0.025709f
C358 VTAIL.n82 B 0.014221f
C359 VTAIL.n83 B 0.013815f
C360 VTAIL.n84 B 0.032653f
C361 VTAIL.n85 B 0.032653f
C362 VTAIL.n86 B 0.014627f
C363 VTAIL.n87 B 0.025709f
C364 VTAIL.n88 B 0.013815f
C365 VTAIL.n89 B 0.032653f
C366 VTAIL.n90 B 0.014627f
C367 VTAIL.n91 B 1.2455f
C368 VTAIL.n92 B 0.013815f
C369 VTAIL.t5 B 0.055087f
C370 VTAIL.n93 B 0.180916f
C371 VTAIL.n94 B 0.023083f
C372 VTAIL.n95 B 0.02449f
C373 VTAIL.n96 B 0.032653f
C374 VTAIL.n97 B 0.014627f
C375 VTAIL.n98 B 0.013815f
C376 VTAIL.n99 B 0.025709f
C377 VTAIL.n100 B 0.025709f
C378 VTAIL.n101 B 0.013815f
C379 VTAIL.n102 B 0.014627f
C380 VTAIL.n103 B 0.032653f
C381 VTAIL.n104 B 0.032653f
C382 VTAIL.n105 B 0.014627f
C383 VTAIL.n106 B 0.013815f
C384 VTAIL.n107 B 0.025709f
C385 VTAIL.n108 B 0.025709f
C386 VTAIL.n109 B 0.013815f
C387 VTAIL.n110 B 0.014627f
C388 VTAIL.n111 B 0.032653f
C389 VTAIL.n112 B 0.032653f
C390 VTAIL.n113 B 0.014627f
C391 VTAIL.n114 B 0.013815f
C392 VTAIL.n115 B 0.025709f
C393 VTAIL.n116 B 0.025709f
C394 VTAIL.n117 B 0.013815f
C395 VTAIL.n118 B 0.014627f
C396 VTAIL.n119 B 0.032653f
C397 VTAIL.n120 B 0.032653f
C398 VTAIL.n121 B 0.014627f
C399 VTAIL.n122 B 0.013815f
C400 VTAIL.n123 B 0.025709f
C401 VTAIL.n124 B 0.025709f
C402 VTAIL.n125 B 0.013815f
C403 VTAIL.n126 B 0.014627f
C404 VTAIL.n127 B 0.032653f
C405 VTAIL.n128 B 0.074063f
C406 VTAIL.n129 B 0.014627f
C407 VTAIL.n130 B 0.013815f
C408 VTAIL.n131 B 0.064693f
C409 VTAIL.n132 B 0.041944f
C410 VTAIL.n133 B 0.462343f
C411 VTAIL.t13 B 0.234648f
C412 VTAIL.t16 B 0.234648f
C413 VTAIL.n134 B 2.01803f
C414 VTAIL.n135 B 0.682563f
C415 VTAIL.t11 B 0.234648f
C416 VTAIL.t17 B 0.234648f
C417 VTAIL.n136 B 2.01803f
C418 VTAIL.n137 B 0.776472f
C419 VTAIL.n138 B 0.038044f
C420 VTAIL.n139 B 0.025709f
C421 VTAIL.n140 B 0.013815f
C422 VTAIL.n141 B 0.032653f
C423 VTAIL.n142 B 0.014627f
C424 VTAIL.n143 B 0.025709f
C425 VTAIL.n144 B 0.013815f
C426 VTAIL.n145 B 0.032653f
C427 VTAIL.n146 B 0.014221f
C428 VTAIL.n147 B 0.025709f
C429 VTAIL.n148 B 0.014221f
C430 VTAIL.n149 B 0.013815f
C431 VTAIL.n150 B 0.032653f
C432 VTAIL.n151 B 0.032653f
C433 VTAIL.n152 B 0.014627f
C434 VTAIL.n153 B 0.025709f
C435 VTAIL.n154 B 0.013815f
C436 VTAIL.n155 B 0.032653f
C437 VTAIL.n156 B 0.014627f
C438 VTAIL.n157 B 1.2455f
C439 VTAIL.n158 B 0.013815f
C440 VTAIL.t14 B 0.055087f
C441 VTAIL.n159 B 0.180916f
C442 VTAIL.n160 B 0.023083f
C443 VTAIL.n161 B 0.02449f
C444 VTAIL.n162 B 0.032653f
C445 VTAIL.n163 B 0.014627f
C446 VTAIL.n164 B 0.013815f
C447 VTAIL.n165 B 0.025709f
C448 VTAIL.n166 B 0.025709f
C449 VTAIL.n167 B 0.013815f
C450 VTAIL.n168 B 0.014627f
C451 VTAIL.n169 B 0.032653f
C452 VTAIL.n170 B 0.032653f
C453 VTAIL.n171 B 0.014627f
C454 VTAIL.n172 B 0.013815f
C455 VTAIL.n173 B 0.025709f
C456 VTAIL.n174 B 0.025709f
C457 VTAIL.n175 B 0.013815f
C458 VTAIL.n176 B 0.014627f
C459 VTAIL.n177 B 0.032653f
C460 VTAIL.n178 B 0.032653f
C461 VTAIL.n179 B 0.014627f
C462 VTAIL.n180 B 0.013815f
C463 VTAIL.n181 B 0.025709f
C464 VTAIL.n182 B 0.025709f
C465 VTAIL.n183 B 0.013815f
C466 VTAIL.n184 B 0.014627f
C467 VTAIL.n185 B 0.032653f
C468 VTAIL.n186 B 0.032653f
C469 VTAIL.n187 B 0.014627f
C470 VTAIL.n188 B 0.013815f
C471 VTAIL.n189 B 0.025709f
C472 VTAIL.n190 B 0.025709f
C473 VTAIL.n191 B 0.013815f
C474 VTAIL.n192 B 0.014627f
C475 VTAIL.n193 B 0.032653f
C476 VTAIL.n194 B 0.074063f
C477 VTAIL.n195 B 0.014627f
C478 VTAIL.n196 B 0.013815f
C479 VTAIL.n197 B 0.064693f
C480 VTAIL.n198 B 0.041944f
C481 VTAIL.n199 B 1.7303f
C482 VTAIL.n200 B 0.038044f
C483 VTAIL.n201 B 0.025709f
C484 VTAIL.n202 B 0.013815f
C485 VTAIL.n203 B 0.032653f
C486 VTAIL.n204 B 0.014627f
C487 VTAIL.n205 B 0.025709f
C488 VTAIL.n206 B 0.013815f
C489 VTAIL.n207 B 0.032653f
C490 VTAIL.n208 B 0.014221f
C491 VTAIL.n209 B 0.025709f
C492 VTAIL.n210 B 0.014627f
C493 VTAIL.n211 B 0.032653f
C494 VTAIL.n212 B 0.014627f
C495 VTAIL.n213 B 0.025709f
C496 VTAIL.n214 B 0.013815f
C497 VTAIL.n215 B 0.032653f
C498 VTAIL.n216 B 0.014627f
C499 VTAIL.n217 B 1.2455f
C500 VTAIL.n218 B 0.013815f
C501 VTAIL.t3 B 0.055087f
C502 VTAIL.n219 B 0.180916f
C503 VTAIL.n220 B 0.023083f
C504 VTAIL.n221 B 0.02449f
C505 VTAIL.n222 B 0.032653f
C506 VTAIL.n223 B 0.014627f
C507 VTAIL.n224 B 0.013815f
C508 VTAIL.n225 B 0.025709f
C509 VTAIL.n226 B 0.025709f
C510 VTAIL.n227 B 0.013815f
C511 VTAIL.n228 B 0.014627f
C512 VTAIL.n229 B 0.032653f
C513 VTAIL.n230 B 0.032653f
C514 VTAIL.n231 B 0.014627f
C515 VTAIL.n232 B 0.013815f
C516 VTAIL.n233 B 0.025709f
C517 VTAIL.n234 B 0.025709f
C518 VTAIL.n235 B 0.013815f
C519 VTAIL.n236 B 0.013815f
C520 VTAIL.n237 B 0.014627f
C521 VTAIL.n238 B 0.032653f
C522 VTAIL.n239 B 0.032653f
C523 VTAIL.n240 B 0.032653f
C524 VTAIL.n241 B 0.014221f
C525 VTAIL.n242 B 0.013815f
C526 VTAIL.n243 B 0.025709f
C527 VTAIL.n244 B 0.025709f
C528 VTAIL.n245 B 0.013815f
C529 VTAIL.n246 B 0.014627f
C530 VTAIL.n247 B 0.032653f
C531 VTAIL.n248 B 0.032653f
C532 VTAIL.n249 B 0.014627f
C533 VTAIL.n250 B 0.013815f
C534 VTAIL.n251 B 0.025709f
C535 VTAIL.n252 B 0.025709f
C536 VTAIL.n253 B 0.013815f
C537 VTAIL.n254 B 0.014627f
C538 VTAIL.n255 B 0.032653f
C539 VTAIL.n256 B 0.074063f
C540 VTAIL.n257 B 0.014627f
C541 VTAIL.n258 B 0.013815f
C542 VTAIL.n259 B 0.064693f
C543 VTAIL.n260 B 0.041944f
C544 VTAIL.n261 B 1.7303f
C545 VTAIL.t1 B 0.234648f
C546 VTAIL.t4 B 0.234648f
C547 VTAIL.n262 B 2.01802f
C548 VTAIL.n263 B 0.57242f
C549 VDD1.n0 B 0.037094f
C550 VDD1.n1 B 0.025067f
C551 VDD1.n2 B 0.01347f
C552 VDD1.n3 B 0.031838f
C553 VDD1.n4 B 0.014262f
C554 VDD1.n5 B 0.025067f
C555 VDD1.n6 B 0.01347f
C556 VDD1.n7 B 0.031838f
C557 VDD1.n8 B 0.013866f
C558 VDD1.n9 B 0.025067f
C559 VDD1.n10 B 0.013866f
C560 VDD1.n11 B 0.01347f
C561 VDD1.n12 B 0.031838f
C562 VDD1.n13 B 0.031838f
C563 VDD1.n14 B 0.014262f
C564 VDD1.n15 B 0.025067f
C565 VDD1.n16 B 0.01347f
C566 VDD1.n17 B 0.031838f
C567 VDD1.n18 B 0.014262f
C568 VDD1.n19 B 1.21441f
C569 VDD1.n20 B 0.01347f
C570 VDD1.t7 B 0.053712f
C571 VDD1.n21 B 0.176399f
C572 VDD1.n22 B 0.022507f
C573 VDD1.n23 B 0.023878f
C574 VDD1.n24 B 0.031838f
C575 VDD1.n25 B 0.014262f
C576 VDD1.n26 B 0.01347f
C577 VDD1.n27 B 0.025067f
C578 VDD1.n28 B 0.025067f
C579 VDD1.n29 B 0.01347f
C580 VDD1.n30 B 0.014262f
C581 VDD1.n31 B 0.031838f
C582 VDD1.n32 B 0.031838f
C583 VDD1.n33 B 0.014262f
C584 VDD1.n34 B 0.01347f
C585 VDD1.n35 B 0.025067f
C586 VDD1.n36 B 0.025067f
C587 VDD1.n37 B 0.01347f
C588 VDD1.n38 B 0.014262f
C589 VDD1.n39 B 0.031838f
C590 VDD1.n40 B 0.031838f
C591 VDD1.n41 B 0.014262f
C592 VDD1.n42 B 0.01347f
C593 VDD1.n43 B 0.025067f
C594 VDD1.n44 B 0.025067f
C595 VDD1.n45 B 0.01347f
C596 VDD1.n46 B 0.014262f
C597 VDD1.n47 B 0.031838f
C598 VDD1.n48 B 0.031838f
C599 VDD1.n49 B 0.014262f
C600 VDD1.n50 B 0.01347f
C601 VDD1.n51 B 0.025067f
C602 VDD1.n52 B 0.025067f
C603 VDD1.n53 B 0.01347f
C604 VDD1.n54 B 0.014262f
C605 VDD1.n55 B 0.031838f
C606 VDD1.n56 B 0.072213f
C607 VDD1.n57 B 0.014262f
C608 VDD1.n58 B 0.01347f
C609 VDD1.n59 B 0.063077f
C610 VDD1.n60 B 0.076263f
C611 VDD1.t4 B 0.228789f
C612 VDD1.t9 B 0.228789f
C613 VDD1.n61 B 2.0365f
C614 VDD1.n62 B 0.824871f
C615 VDD1.n63 B 0.037094f
C616 VDD1.n64 B 0.025067f
C617 VDD1.n65 B 0.01347f
C618 VDD1.n66 B 0.031838f
C619 VDD1.n67 B 0.014262f
C620 VDD1.n68 B 0.025067f
C621 VDD1.n69 B 0.01347f
C622 VDD1.n70 B 0.031838f
C623 VDD1.n71 B 0.013866f
C624 VDD1.n72 B 0.025067f
C625 VDD1.n73 B 0.014262f
C626 VDD1.n74 B 0.031838f
C627 VDD1.n75 B 0.014262f
C628 VDD1.n76 B 0.025067f
C629 VDD1.n77 B 0.01347f
C630 VDD1.n78 B 0.031838f
C631 VDD1.n79 B 0.014262f
C632 VDD1.n80 B 1.21441f
C633 VDD1.n81 B 0.01347f
C634 VDD1.t1 B 0.053712f
C635 VDD1.n82 B 0.176399f
C636 VDD1.n83 B 0.022507f
C637 VDD1.n84 B 0.023878f
C638 VDD1.n85 B 0.031838f
C639 VDD1.n86 B 0.014262f
C640 VDD1.n87 B 0.01347f
C641 VDD1.n88 B 0.025067f
C642 VDD1.n89 B 0.025067f
C643 VDD1.n90 B 0.01347f
C644 VDD1.n91 B 0.014262f
C645 VDD1.n92 B 0.031838f
C646 VDD1.n93 B 0.031838f
C647 VDD1.n94 B 0.014262f
C648 VDD1.n95 B 0.01347f
C649 VDD1.n96 B 0.025067f
C650 VDD1.n97 B 0.025067f
C651 VDD1.n98 B 0.01347f
C652 VDD1.n99 B 0.01347f
C653 VDD1.n100 B 0.014262f
C654 VDD1.n101 B 0.031838f
C655 VDD1.n102 B 0.031838f
C656 VDD1.n103 B 0.031838f
C657 VDD1.n104 B 0.013866f
C658 VDD1.n105 B 0.01347f
C659 VDD1.n106 B 0.025067f
C660 VDD1.n107 B 0.025067f
C661 VDD1.n108 B 0.01347f
C662 VDD1.n109 B 0.014262f
C663 VDD1.n110 B 0.031838f
C664 VDD1.n111 B 0.031838f
C665 VDD1.n112 B 0.014262f
C666 VDD1.n113 B 0.01347f
C667 VDD1.n114 B 0.025067f
C668 VDD1.n115 B 0.025067f
C669 VDD1.n116 B 0.01347f
C670 VDD1.n117 B 0.014262f
C671 VDD1.n118 B 0.031838f
C672 VDD1.n119 B 0.072213f
C673 VDD1.n120 B 0.014262f
C674 VDD1.n121 B 0.01347f
C675 VDD1.n122 B 0.063077f
C676 VDD1.n123 B 0.076263f
C677 VDD1.t2 B 0.228789f
C678 VDD1.t3 B 0.228789f
C679 VDD1.n124 B 2.03649f
C680 VDD1.n125 B 0.816487f
C681 VDD1.t8 B 0.228789f
C682 VDD1.t6 B 0.228789f
C683 VDD1.n126 B 2.05963f
C684 VDD1.n127 B 3.44312f
C685 VDD1.t5 B 0.228789f
C686 VDD1.t0 B 0.228789f
C687 VDD1.n128 B 2.03649f
C688 VDD1.n129 B 3.47368f
C689 VP.t5 B 1.97084f
C690 VP.n0 B 0.76203f
C691 VP.n1 B 0.018495f
C692 VP.n2 B 0.022876f
C693 VP.n3 B 0.018495f
C694 VP.n4 B 0.018473f
C695 VP.n5 B 0.018495f
C696 VP.n6 B 0.01804f
C697 VP.n7 B 0.018495f
C698 VP.t8 B 1.97084f
C699 VP.n8 B 0.693488f
C700 VP.n9 B 0.018495f
C701 VP.n10 B 0.01804f
C702 VP.n11 B 0.018495f
C703 VP.t9 B 1.97084f
C704 VP.n12 B 0.693488f
C705 VP.n13 B 0.018495f
C706 VP.n14 B 0.031122f
C707 VP.n15 B 0.018495f
C708 VP.n16 B 0.023919f
C709 VP.t3 B 1.97084f
C710 VP.n17 B 0.76203f
C711 VP.n18 B 0.018495f
C712 VP.n19 B 0.022876f
C713 VP.n20 B 0.018495f
C714 VP.n21 B 0.018473f
C715 VP.n22 B 0.018495f
C716 VP.n23 B 0.01804f
C717 VP.n24 B 0.018495f
C718 VP.t6 B 1.97084f
C719 VP.n25 B 0.693488f
C720 VP.n26 B 0.018495f
C721 VP.n27 B 0.01804f
C722 VP.n28 B 0.018495f
C723 VP.t1 B 1.97084f
C724 VP.n29 B 0.765017f
C725 VP.t4 B 2.20999f
C726 VP.n30 B 0.721893f
C727 VP.n31 B 0.22633f
C728 VP.n32 B 0.033448f
C729 VP.n33 B 0.03447f
C730 VP.n34 B 0.03358f
C731 VP.n35 B 0.018495f
C732 VP.n36 B 0.018495f
C733 VP.n37 B 0.018495f
C734 VP.n38 B 0.036847f
C735 VP.n39 B 0.03447f
C736 VP.n40 B 0.025961f
C737 VP.n41 B 0.018495f
C738 VP.n42 B 0.018495f
C739 VP.n43 B 0.025961f
C740 VP.n44 B 0.03447f
C741 VP.n45 B 0.036847f
C742 VP.n46 B 0.018495f
C743 VP.n47 B 0.018495f
C744 VP.n48 B 0.018495f
C745 VP.n49 B 0.03358f
C746 VP.n50 B 0.03447f
C747 VP.t0 B 1.97084f
C748 VP.n51 B 0.693488f
C749 VP.n52 B 0.033448f
C750 VP.n53 B 0.018495f
C751 VP.n54 B 0.018495f
C752 VP.n55 B 0.018495f
C753 VP.n56 B 0.03447f
C754 VP.n57 B 0.03447f
C755 VP.n58 B 0.031122f
C756 VP.n59 B 0.018495f
C757 VP.n60 B 0.018495f
C758 VP.n61 B 0.018495f
C759 VP.n62 B 0.03447f
C760 VP.n63 B 0.03447f
C761 VP.n64 B 0.023919f
C762 VP.n65 B 0.02985f
C763 VP.n66 B 1.27094f
C764 VP.t2 B 1.97084f
C765 VP.n67 B 0.76203f
C766 VP.n68 B 1.28258f
C767 VP.n69 B 0.02985f
C768 VP.n70 B 0.018495f
C769 VP.n71 B 0.03447f
C770 VP.n72 B 0.03447f
C771 VP.n73 B 0.022876f
C772 VP.n74 B 0.018495f
C773 VP.n75 B 0.018495f
C774 VP.n76 B 0.018495f
C775 VP.n77 B 0.03447f
C776 VP.n78 B 0.03447f
C777 VP.n79 B 0.018473f
C778 VP.n80 B 0.018495f
C779 VP.n81 B 0.018495f
C780 VP.n82 B 0.033448f
C781 VP.n83 B 0.03447f
C782 VP.n84 B 0.03358f
C783 VP.n85 B 0.018495f
C784 VP.n86 B 0.018495f
C785 VP.n87 B 0.018495f
C786 VP.n88 B 0.036847f
C787 VP.n89 B 0.03447f
C788 VP.n90 B 0.025961f
C789 VP.n91 B 0.018495f
C790 VP.n92 B 0.018495f
C791 VP.n93 B 0.025961f
C792 VP.n94 B 0.03447f
C793 VP.n95 B 0.036847f
C794 VP.n96 B 0.018495f
C795 VP.n97 B 0.018495f
C796 VP.n98 B 0.018495f
C797 VP.n99 B 0.03358f
C798 VP.n100 B 0.03447f
C799 VP.t7 B 1.97084f
C800 VP.n101 B 0.693488f
C801 VP.n102 B 0.033448f
C802 VP.n103 B 0.018495f
C803 VP.n104 B 0.018495f
C804 VP.n105 B 0.018495f
C805 VP.n106 B 0.03447f
C806 VP.n107 B 0.03447f
C807 VP.n108 B 0.031122f
C808 VP.n109 B 0.018495f
C809 VP.n110 B 0.018495f
C810 VP.n111 B 0.018495f
C811 VP.n112 B 0.03447f
C812 VP.n113 B 0.03447f
C813 VP.n114 B 0.023919f
C814 VP.n115 B 0.02985f
C815 VP.n116 B 0.049146f
.ends

