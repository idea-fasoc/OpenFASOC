* NGSPICE file created from diff_pair_sample_0593.ext - technology: sky130A

.subckt diff_pair_sample_0593 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X1 VTAIL.t13 VP.t1 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=2.29515 ps=14.24 w=13.91 l=3.72
X2 VDD1.t0 VP.t2 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X3 VDD2.t7 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X4 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=0 ps=0 w=13.91 l=3.72
X5 VDD2.t6 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X6 VTAIL.t15 VN.t2 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=2.29515 ps=14.24 w=13.91 l=3.72
X7 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=0 ps=0 w=13.91 l=3.72
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=0 ps=0 w=13.91 l=3.72
X9 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=2.29515 ps=14.24 w=13.91 l=3.72
X10 VDD2.t3 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=5.4249 ps=28.6 w=13.91 l=3.72
X11 VDD2.t2 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=5.4249 ps=28.6 w=13.91 l=3.72
X12 VTAIL.t11 VP.t3 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X13 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X14 VTAIL.t10 VP.t4 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=2.29515 ps=14.24 w=13.91 l=3.72
X15 VDD1.t3 VP.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=5.4249 ps=28.6 w=13.91 l=3.72
X16 VDD1.t2 VP.t6 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.4249 pd=28.6 as=0 ps=0 w=13.91 l=3.72
X18 VTAIL.t6 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=2.29515 ps=14.24 w=13.91 l=3.72
X19 VDD1.t5 VP.t7 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.29515 pd=14.24 as=5.4249 ps=28.6 w=13.91 l=3.72
R0 VP.n25 VP.n24 161.3
R1 VP.n26 VP.n21 161.3
R2 VP.n28 VP.n27 161.3
R3 VP.n29 VP.n20 161.3
R4 VP.n31 VP.n30 161.3
R5 VP.n32 VP.n19 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n18 161.3
R8 VP.n38 VP.n37 161.3
R9 VP.n39 VP.n17 161.3
R10 VP.n41 VP.n40 161.3
R11 VP.n42 VP.n16 161.3
R12 VP.n44 VP.n43 161.3
R13 VP.n45 VP.n15 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n48 VP.n14 161.3
R16 VP.n50 VP.n49 161.3
R17 VP.n93 VP.n92 161.3
R18 VP.n91 VP.n1 161.3
R19 VP.n90 VP.n89 161.3
R20 VP.n88 VP.n2 161.3
R21 VP.n87 VP.n86 161.3
R22 VP.n85 VP.n3 161.3
R23 VP.n84 VP.n83 161.3
R24 VP.n82 VP.n4 161.3
R25 VP.n81 VP.n80 161.3
R26 VP.n78 VP.n5 161.3
R27 VP.n77 VP.n76 161.3
R28 VP.n75 VP.n6 161.3
R29 VP.n74 VP.n73 161.3
R30 VP.n72 VP.n7 161.3
R31 VP.n71 VP.n70 161.3
R32 VP.n69 VP.n8 161.3
R33 VP.n68 VP.n67 161.3
R34 VP.n65 VP.n9 161.3
R35 VP.n64 VP.n63 161.3
R36 VP.n62 VP.n10 161.3
R37 VP.n61 VP.n60 161.3
R38 VP.n59 VP.n11 161.3
R39 VP.n58 VP.n57 161.3
R40 VP.n56 VP.n12 161.3
R41 VP.n55 VP.n54 161.3
R42 VP.n22 VP.t1 122.177
R43 VP.n53 VP.t4 90.1164
R44 VP.n66 VP.t6 90.1164
R45 VP.n79 VP.t0 90.1164
R46 VP.n0 VP.t7 90.1164
R47 VP.n13 VP.t5 90.1164
R48 VP.n36 VP.t3 90.1164
R49 VP.n23 VP.t2 90.1164
R50 VP.n53 VP.n52 86.3974
R51 VP.n94 VP.n0 86.3974
R52 VP.n51 VP.n13 86.3974
R53 VP.n23 VP.n22 73.7323
R54 VP.n52 VP.n51 57.6281
R55 VP.n60 VP.n59 45.3497
R56 VP.n86 VP.n2 45.3497
R57 VP.n43 VP.n15 45.3497
R58 VP.n73 VP.n72 40.4934
R59 VP.n73 VP.n6 40.4934
R60 VP.n30 VP.n19 40.4934
R61 VP.n30 VP.n29 40.4934
R62 VP.n60 VP.n10 35.6371
R63 VP.n86 VP.n85 35.6371
R64 VP.n43 VP.n42 35.6371
R65 VP.n54 VP.n12 24.4675
R66 VP.n58 VP.n12 24.4675
R67 VP.n59 VP.n58 24.4675
R68 VP.n64 VP.n10 24.4675
R69 VP.n65 VP.n64 24.4675
R70 VP.n67 VP.n8 24.4675
R71 VP.n71 VP.n8 24.4675
R72 VP.n72 VP.n71 24.4675
R73 VP.n77 VP.n6 24.4675
R74 VP.n78 VP.n77 24.4675
R75 VP.n80 VP.n78 24.4675
R76 VP.n84 VP.n4 24.4675
R77 VP.n85 VP.n84 24.4675
R78 VP.n90 VP.n2 24.4675
R79 VP.n91 VP.n90 24.4675
R80 VP.n92 VP.n91 24.4675
R81 VP.n47 VP.n15 24.4675
R82 VP.n48 VP.n47 24.4675
R83 VP.n49 VP.n48 24.4675
R84 VP.n34 VP.n19 24.4675
R85 VP.n35 VP.n34 24.4675
R86 VP.n37 VP.n35 24.4675
R87 VP.n41 VP.n17 24.4675
R88 VP.n42 VP.n41 24.4675
R89 VP.n24 VP.n21 24.4675
R90 VP.n28 VP.n21 24.4675
R91 VP.n29 VP.n28 24.4675
R92 VP.n66 VP.n65 23.2442
R93 VP.n79 VP.n4 23.2442
R94 VP.n36 VP.n17 23.2442
R95 VP.n54 VP.n53 3.67055
R96 VP.n92 VP.n0 3.67055
R97 VP.n49 VP.n13 3.67055
R98 VP.n25 VP.n22 3.35318
R99 VP.n67 VP.n66 1.22385
R100 VP.n80 VP.n79 1.22385
R101 VP.n37 VP.n36 1.22385
R102 VP.n24 VP.n23 1.22385
R103 VP.n51 VP.n50 0.354971
R104 VP.n55 VP.n52 0.354971
R105 VP.n94 VP.n93 0.354971
R106 VP VP.n94 0.26696
R107 VP.n26 VP.n25 0.189894
R108 VP.n27 VP.n26 0.189894
R109 VP.n27 VP.n20 0.189894
R110 VP.n31 VP.n20 0.189894
R111 VP.n32 VP.n31 0.189894
R112 VP.n33 VP.n32 0.189894
R113 VP.n33 VP.n18 0.189894
R114 VP.n38 VP.n18 0.189894
R115 VP.n39 VP.n38 0.189894
R116 VP.n40 VP.n39 0.189894
R117 VP.n40 VP.n16 0.189894
R118 VP.n44 VP.n16 0.189894
R119 VP.n45 VP.n44 0.189894
R120 VP.n46 VP.n45 0.189894
R121 VP.n46 VP.n14 0.189894
R122 VP.n50 VP.n14 0.189894
R123 VP.n56 VP.n55 0.189894
R124 VP.n57 VP.n56 0.189894
R125 VP.n57 VP.n11 0.189894
R126 VP.n61 VP.n11 0.189894
R127 VP.n62 VP.n61 0.189894
R128 VP.n63 VP.n62 0.189894
R129 VP.n63 VP.n9 0.189894
R130 VP.n68 VP.n9 0.189894
R131 VP.n69 VP.n68 0.189894
R132 VP.n70 VP.n69 0.189894
R133 VP.n70 VP.n7 0.189894
R134 VP.n74 VP.n7 0.189894
R135 VP.n75 VP.n74 0.189894
R136 VP.n76 VP.n75 0.189894
R137 VP.n76 VP.n5 0.189894
R138 VP.n81 VP.n5 0.189894
R139 VP.n82 VP.n81 0.189894
R140 VP.n83 VP.n82 0.189894
R141 VP.n83 VP.n3 0.189894
R142 VP.n87 VP.n3 0.189894
R143 VP.n88 VP.n87 0.189894
R144 VP.n89 VP.n88 0.189894
R145 VP.n89 VP.n1 0.189894
R146 VP.n93 VP.n1 0.189894
R147 VDD1 VDD1.n0 63.0982
R148 VDD1.n3 VDD1.n2 62.9847
R149 VDD1.n3 VDD1.n1 62.9847
R150 VDD1.n5 VDD1.n4 61.2944
R151 VDD1.n5 VDD1.n3 52.0009
R152 VDD1 VDD1.n5 1.688
R153 VDD1.n4 VDD1.t7 1.42394
R154 VDD1.n4 VDD1.t3 1.42394
R155 VDD1.n0 VDD1.t1 1.42394
R156 VDD1.n0 VDD1.t0 1.42394
R157 VDD1.n2 VDD1.t4 1.42394
R158 VDD1.n2 VDD1.t5 1.42394
R159 VDD1.n1 VDD1.t6 1.42394
R160 VDD1.n1 VDD1.t2 1.42394
R161 VTAIL.n14 VTAIL.t9 46.039
R162 VTAIL.n11 VTAIL.t13 46.039
R163 VTAIL.n10 VTAIL.t2 46.039
R164 VTAIL.n7 VTAIL.t1 46.039
R165 VTAIL.n15 VTAIL.t0 46.0388
R166 VTAIL.n2 VTAIL.t15 46.0388
R167 VTAIL.n3 VTAIL.t7 46.0388
R168 VTAIL.n6 VTAIL.t10 46.0388
R169 VTAIL.n13 VTAIL.n12 44.6156
R170 VTAIL.n9 VTAIL.n8 44.6156
R171 VTAIL.n1 VTAIL.n0 44.6155
R172 VTAIL.n5 VTAIL.n4 44.6155
R173 VTAIL.n15 VTAIL.n14 27.8496
R174 VTAIL.n7 VTAIL.n6 27.8496
R175 VTAIL.n9 VTAIL.n7 3.49188
R176 VTAIL.n10 VTAIL.n9 3.49188
R177 VTAIL.n13 VTAIL.n11 3.49188
R178 VTAIL.n14 VTAIL.n13 3.49188
R179 VTAIL.n6 VTAIL.n5 3.49188
R180 VTAIL.n5 VTAIL.n3 3.49188
R181 VTAIL.n2 VTAIL.n1 3.49188
R182 VTAIL VTAIL.n15 3.43369
R183 VTAIL.n0 VTAIL.t5 1.42394
R184 VTAIL.n0 VTAIL.t4 1.42394
R185 VTAIL.n4 VTAIL.t8 1.42394
R186 VTAIL.n4 VTAIL.t14 1.42394
R187 VTAIL.n12 VTAIL.t12 1.42394
R188 VTAIL.n12 VTAIL.t11 1.42394
R189 VTAIL.n8 VTAIL.t3 1.42394
R190 VTAIL.n8 VTAIL.t6 1.42394
R191 VTAIL.n11 VTAIL.n10 0.470328
R192 VTAIL.n3 VTAIL.n2 0.470328
R193 VTAIL VTAIL.n1 0.0586897
R194 B.n1069 B.n1068 585
R195 B.n383 B.n175 585
R196 B.n382 B.n381 585
R197 B.n380 B.n379 585
R198 B.n378 B.n377 585
R199 B.n376 B.n375 585
R200 B.n374 B.n373 585
R201 B.n372 B.n371 585
R202 B.n370 B.n369 585
R203 B.n368 B.n367 585
R204 B.n366 B.n365 585
R205 B.n364 B.n363 585
R206 B.n362 B.n361 585
R207 B.n360 B.n359 585
R208 B.n358 B.n357 585
R209 B.n356 B.n355 585
R210 B.n354 B.n353 585
R211 B.n352 B.n351 585
R212 B.n350 B.n349 585
R213 B.n348 B.n347 585
R214 B.n346 B.n345 585
R215 B.n344 B.n343 585
R216 B.n342 B.n341 585
R217 B.n340 B.n339 585
R218 B.n338 B.n337 585
R219 B.n336 B.n335 585
R220 B.n334 B.n333 585
R221 B.n332 B.n331 585
R222 B.n330 B.n329 585
R223 B.n328 B.n327 585
R224 B.n326 B.n325 585
R225 B.n324 B.n323 585
R226 B.n322 B.n321 585
R227 B.n320 B.n319 585
R228 B.n318 B.n317 585
R229 B.n316 B.n315 585
R230 B.n314 B.n313 585
R231 B.n312 B.n311 585
R232 B.n310 B.n309 585
R233 B.n308 B.n307 585
R234 B.n306 B.n305 585
R235 B.n304 B.n303 585
R236 B.n302 B.n301 585
R237 B.n300 B.n299 585
R238 B.n298 B.n297 585
R239 B.n296 B.n295 585
R240 B.n294 B.n293 585
R241 B.n291 B.n290 585
R242 B.n289 B.n288 585
R243 B.n287 B.n286 585
R244 B.n285 B.n284 585
R245 B.n283 B.n282 585
R246 B.n281 B.n280 585
R247 B.n279 B.n278 585
R248 B.n277 B.n276 585
R249 B.n275 B.n274 585
R250 B.n273 B.n272 585
R251 B.n270 B.n269 585
R252 B.n268 B.n267 585
R253 B.n266 B.n265 585
R254 B.n264 B.n263 585
R255 B.n262 B.n261 585
R256 B.n260 B.n259 585
R257 B.n258 B.n257 585
R258 B.n256 B.n255 585
R259 B.n254 B.n253 585
R260 B.n252 B.n251 585
R261 B.n250 B.n249 585
R262 B.n248 B.n247 585
R263 B.n246 B.n245 585
R264 B.n244 B.n243 585
R265 B.n242 B.n241 585
R266 B.n240 B.n239 585
R267 B.n238 B.n237 585
R268 B.n236 B.n235 585
R269 B.n234 B.n233 585
R270 B.n232 B.n231 585
R271 B.n230 B.n229 585
R272 B.n228 B.n227 585
R273 B.n226 B.n225 585
R274 B.n224 B.n223 585
R275 B.n222 B.n221 585
R276 B.n220 B.n219 585
R277 B.n218 B.n217 585
R278 B.n216 B.n215 585
R279 B.n214 B.n213 585
R280 B.n212 B.n211 585
R281 B.n210 B.n209 585
R282 B.n208 B.n207 585
R283 B.n206 B.n205 585
R284 B.n204 B.n203 585
R285 B.n202 B.n201 585
R286 B.n200 B.n199 585
R287 B.n198 B.n197 585
R288 B.n196 B.n195 585
R289 B.n194 B.n193 585
R290 B.n192 B.n191 585
R291 B.n190 B.n189 585
R292 B.n188 B.n187 585
R293 B.n186 B.n185 585
R294 B.n184 B.n183 585
R295 B.n182 B.n181 585
R296 B.n124 B.n123 585
R297 B.n1074 B.n1073 585
R298 B.n1067 B.n176 585
R299 B.n176 B.n121 585
R300 B.n1066 B.n120 585
R301 B.n1078 B.n120 585
R302 B.n1065 B.n119 585
R303 B.n1079 B.n119 585
R304 B.n1064 B.n118 585
R305 B.n1080 B.n118 585
R306 B.n1063 B.n1062 585
R307 B.n1062 B.n114 585
R308 B.n1061 B.n113 585
R309 B.n1086 B.n113 585
R310 B.n1060 B.n112 585
R311 B.n1087 B.n112 585
R312 B.n1059 B.n111 585
R313 B.n1088 B.n111 585
R314 B.n1058 B.n1057 585
R315 B.n1057 B.n107 585
R316 B.n1056 B.n106 585
R317 B.n1094 B.n106 585
R318 B.n1055 B.n105 585
R319 B.n1095 B.n105 585
R320 B.n1054 B.n104 585
R321 B.n1096 B.n104 585
R322 B.n1053 B.n1052 585
R323 B.n1052 B.n100 585
R324 B.n1051 B.n99 585
R325 B.n1102 B.n99 585
R326 B.n1050 B.n98 585
R327 B.n1103 B.n98 585
R328 B.n1049 B.n97 585
R329 B.n1104 B.n97 585
R330 B.n1048 B.n1047 585
R331 B.n1047 B.n93 585
R332 B.n1046 B.n92 585
R333 B.n1110 B.n92 585
R334 B.n1045 B.n91 585
R335 B.n1111 B.n91 585
R336 B.n1044 B.n90 585
R337 B.n1112 B.n90 585
R338 B.n1043 B.n1042 585
R339 B.n1042 B.n86 585
R340 B.n1041 B.n85 585
R341 B.n1118 B.n85 585
R342 B.n1040 B.n84 585
R343 B.n1119 B.n84 585
R344 B.n1039 B.n83 585
R345 B.n1120 B.n83 585
R346 B.n1038 B.n1037 585
R347 B.n1037 B.n82 585
R348 B.n1036 B.n78 585
R349 B.n1126 B.n78 585
R350 B.n1035 B.n77 585
R351 B.n1127 B.n77 585
R352 B.n1034 B.n76 585
R353 B.n1128 B.n76 585
R354 B.n1033 B.n1032 585
R355 B.n1032 B.n72 585
R356 B.n1031 B.n71 585
R357 B.n1134 B.n71 585
R358 B.n1030 B.n70 585
R359 B.n1135 B.n70 585
R360 B.n1029 B.n69 585
R361 B.n1136 B.n69 585
R362 B.n1028 B.n1027 585
R363 B.n1027 B.n65 585
R364 B.n1026 B.n64 585
R365 B.n1142 B.n64 585
R366 B.n1025 B.n63 585
R367 B.n1143 B.n63 585
R368 B.n1024 B.n62 585
R369 B.n1144 B.n62 585
R370 B.n1023 B.n1022 585
R371 B.n1022 B.n61 585
R372 B.n1021 B.n57 585
R373 B.n1150 B.n57 585
R374 B.n1020 B.n56 585
R375 B.n1151 B.n56 585
R376 B.n1019 B.n55 585
R377 B.n1152 B.n55 585
R378 B.n1018 B.n1017 585
R379 B.n1017 B.n51 585
R380 B.n1016 B.n50 585
R381 B.n1158 B.n50 585
R382 B.n1015 B.n49 585
R383 B.n1159 B.n49 585
R384 B.n1014 B.n48 585
R385 B.n1160 B.n48 585
R386 B.n1013 B.n1012 585
R387 B.n1012 B.n44 585
R388 B.n1011 B.n43 585
R389 B.n1166 B.n43 585
R390 B.n1010 B.n42 585
R391 B.n1167 B.n42 585
R392 B.n1009 B.n41 585
R393 B.n1168 B.n41 585
R394 B.n1008 B.n1007 585
R395 B.n1007 B.n40 585
R396 B.n1006 B.n36 585
R397 B.n1174 B.n36 585
R398 B.n1005 B.n35 585
R399 B.n1175 B.n35 585
R400 B.n1004 B.n34 585
R401 B.n1176 B.n34 585
R402 B.n1003 B.n1002 585
R403 B.n1002 B.n30 585
R404 B.n1001 B.n29 585
R405 B.n1182 B.n29 585
R406 B.n1000 B.n28 585
R407 B.n1183 B.n28 585
R408 B.n999 B.n27 585
R409 B.n1184 B.n27 585
R410 B.n998 B.n997 585
R411 B.n997 B.n23 585
R412 B.n996 B.n22 585
R413 B.n1190 B.n22 585
R414 B.n995 B.n21 585
R415 B.n1191 B.n21 585
R416 B.n994 B.n20 585
R417 B.n1192 B.n20 585
R418 B.n993 B.n992 585
R419 B.n992 B.n16 585
R420 B.n991 B.n15 585
R421 B.n1198 B.n15 585
R422 B.n990 B.n14 585
R423 B.n1199 B.n14 585
R424 B.n989 B.n13 585
R425 B.n1200 B.n13 585
R426 B.n988 B.n987 585
R427 B.n987 B.n12 585
R428 B.n986 B.n985 585
R429 B.n986 B.n8 585
R430 B.n984 B.n7 585
R431 B.n1207 B.n7 585
R432 B.n983 B.n6 585
R433 B.n1208 B.n6 585
R434 B.n982 B.n5 585
R435 B.n1209 B.n5 585
R436 B.n981 B.n980 585
R437 B.n980 B.n4 585
R438 B.n979 B.n384 585
R439 B.n979 B.n978 585
R440 B.n969 B.n385 585
R441 B.n386 B.n385 585
R442 B.n971 B.n970 585
R443 B.n972 B.n971 585
R444 B.n968 B.n391 585
R445 B.n391 B.n390 585
R446 B.n967 B.n966 585
R447 B.n966 B.n965 585
R448 B.n393 B.n392 585
R449 B.n394 B.n393 585
R450 B.n958 B.n957 585
R451 B.n959 B.n958 585
R452 B.n956 B.n399 585
R453 B.n399 B.n398 585
R454 B.n955 B.n954 585
R455 B.n954 B.n953 585
R456 B.n401 B.n400 585
R457 B.n402 B.n401 585
R458 B.n946 B.n945 585
R459 B.n947 B.n946 585
R460 B.n944 B.n407 585
R461 B.n407 B.n406 585
R462 B.n943 B.n942 585
R463 B.n942 B.n941 585
R464 B.n409 B.n408 585
R465 B.n410 B.n409 585
R466 B.n934 B.n933 585
R467 B.n935 B.n934 585
R468 B.n932 B.n415 585
R469 B.n415 B.n414 585
R470 B.n931 B.n930 585
R471 B.n930 B.n929 585
R472 B.n417 B.n416 585
R473 B.n922 B.n417 585
R474 B.n921 B.n920 585
R475 B.n923 B.n921 585
R476 B.n919 B.n422 585
R477 B.n422 B.n421 585
R478 B.n918 B.n917 585
R479 B.n917 B.n916 585
R480 B.n424 B.n423 585
R481 B.n425 B.n424 585
R482 B.n909 B.n908 585
R483 B.n910 B.n909 585
R484 B.n907 B.n430 585
R485 B.n430 B.n429 585
R486 B.n906 B.n905 585
R487 B.n905 B.n904 585
R488 B.n432 B.n431 585
R489 B.n433 B.n432 585
R490 B.n897 B.n896 585
R491 B.n898 B.n897 585
R492 B.n895 B.n438 585
R493 B.n438 B.n437 585
R494 B.n894 B.n893 585
R495 B.n893 B.n892 585
R496 B.n440 B.n439 585
R497 B.n885 B.n440 585
R498 B.n884 B.n883 585
R499 B.n886 B.n884 585
R500 B.n882 B.n445 585
R501 B.n445 B.n444 585
R502 B.n881 B.n880 585
R503 B.n880 B.n879 585
R504 B.n447 B.n446 585
R505 B.n448 B.n447 585
R506 B.n872 B.n871 585
R507 B.n873 B.n872 585
R508 B.n870 B.n453 585
R509 B.n453 B.n452 585
R510 B.n869 B.n868 585
R511 B.n868 B.n867 585
R512 B.n455 B.n454 585
R513 B.n456 B.n455 585
R514 B.n860 B.n859 585
R515 B.n861 B.n860 585
R516 B.n858 B.n461 585
R517 B.n461 B.n460 585
R518 B.n857 B.n856 585
R519 B.n856 B.n855 585
R520 B.n463 B.n462 585
R521 B.n848 B.n463 585
R522 B.n847 B.n846 585
R523 B.n849 B.n847 585
R524 B.n845 B.n468 585
R525 B.n468 B.n467 585
R526 B.n844 B.n843 585
R527 B.n843 B.n842 585
R528 B.n470 B.n469 585
R529 B.n471 B.n470 585
R530 B.n835 B.n834 585
R531 B.n836 B.n835 585
R532 B.n833 B.n476 585
R533 B.n476 B.n475 585
R534 B.n832 B.n831 585
R535 B.n831 B.n830 585
R536 B.n478 B.n477 585
R537 B.n479 B.n478 585
R538 B.n823 B.n822 585
R539 B.n824 B.n823 585
R540 B.n821 B.n484 585
R541 B.n484 B.n483 585
R542 B.n820 B.n819 585
R543 B.n819 B.n818 585
R544 B.n486 B.n485 585
R545 B.n487 B.n486 585
R546 B.n811 B.n810 585
R547 B.n812 B.n811 585
R548 B.n809 B.n492 585
R549 B.n492 B.n491 585
R550 B.n808 B.n807 585
R551 B.n807 B.n806 585
R552 B.n494 B.n493 585
R553 B.n495 B.n494 585
R554 B.n799 B.n798 585
R555 B.n800 B.n799 585
R556 B.n797 B.n500 585
R557 B.n500 B.n499 585
R558 B.n796 B.n795 585
R559 B.n795 B.n794 585
R560 B.n502 B.n501 585
R561 B.n503 B.n502 585
R562 B.n787 B.n786 585
R563 B.n788 B.n787 585
R564 B.n785 B.n508 585
R565 B.n508 B.n507 585
R566 B.n784 B.n783 585
R567 B.n783 B.n782 585
R568 B.n510 B.n509 585
R569 B.n511 B.n510 585
R570 B.n778 B.n777 585
R571 B.n514 B.n513 585
R572 B.n774 B.n773 585
R573 B.n775 B.n774 585
R574 B.n772 B.n566 585
R575 B.n771 B.n770 585
R576 B.n769 B.n768 585
R577 B.n767 B.n766 585
R578 B.n765 B.n764 585
R579 B.n763 B.n762 585
R580 B.n761 B.n760 585
R581 B.n759 B.n758 585
R582 B.n757 B.n756 585
R583 B.n755 B.n754 585
R584 B.n753 B.n752 585
R585 B.n751 B.n750 585
R586 B.n749 B.n748 585
R587 B.n747 B.n746 585
R588 B.n745 B.n744 585
R589 B.n743 B.n742 585
R590 B.n741 B.n740 585
R591 B.n739 B.n738 585
R592 B.n737 B.n736 585
R593 B.n735 B.n734 585
R594 B.n733 B.n732 585
R595 B.n731 B.n730 585
R596 B.n729 B.n728 585
R597 B.n727 B.n726 585
R598 B.n725 B.n724 585
R599 B.n723 B.n722 585
R600 B.n721 B.n720 585
R601 B.n719 B.n718 585
R602 B.n717 B.n716 585
R603 B.n715 B.n714 585
R604 B.n713 B.n712 585
R605 B.n711 B.n710 585
R606 B.n709 B.n708 585
R607 B.n707 B.n706 585
R608 B.n705 B.n704 585
R609 B.n703 B.n702 585
R610 B.n701 B.n700 585
R611 B.n699 B.n698 585
R612 B.n697 B.n696 585
R613 B.n695 B.n694 585
R614 B.n693 B.n692 585
R615 B.n691 B.n690 585
R616 B.n689 B.n688 585
R617 B.n687 B.n686 585
R618 B.n685 B.n684 585
R619 B.n683 B.n682 585
R620 B.n681 B.n680 585
R621 B.n679 B.n678 585
R622 B.n677 B.n676 585
R623 B.n675 B.n674 585
R624 B.n673 B.n672 585
R625 B.n671 B.n670 585
R626 B.n669 B.n668 585
R627 B.n667 B.n666 585
R628 B.n665 B.n664 585
R629 B.n663 B.n662 585
R630 B.n661 B.n660 585
R631 B.n659 B.n658 585
R632 B.n657 B.n656 585
R633 B.n655 B.n654 585
R634 B.n653 B.n652 585
R635 B.n651 B.n650 585
R636 B.n649 B.n648 585
R637 B.n647 B.n646 585
R638 B.n645 B.n644 585
R639 B.n643 B.n642 585
R640 B.n641 B.n640 585
R641 B.n639 B.n638 585
R642 B.n637 B.n636 585
R643 B.n635 B.n634 585
R644 B.n633 B.n632 585
R645 B.n631 B.n630 585
R646 B.n629 B.n628 585
R647 B.n627 B.n626 585
R648 B.n625 B.n624 585
R649 B.n623 B.n622 585
R650 B.n621 B.n620 585
R651 B.n619 B.n618 585
R652 B.n617 B.n616 585
R653 B.n615 B.n614 585
R654 B.n613 B.n612 585
R655 B.n611 B.n610 585
R656 B.n609 B.n608 585
R657 B.n607 B.n606 585
R658 B.n605 B.n604 585
R659 B.n603 B.n602 585
R660 B.n601 B.n600 585
R661 B.n599 B.n598 585
R662 B.n597 B.n596 585
R663 B.n595 B.n594 585
R664 B.n593 B.n592 585
R665 B.n591 B.n590 585
R666 B.n589 B.n588 585
R667 B.n587 B.n586 585
R668 B.n585 B.n584 585
R669 B.n583 B.n582 585
R670 B.n581 B.n580 585
R671 B.n579 B.n578 585
R672 B.n577 B.n576 585
R673 B.n575 B.n574 585
R674 B.n573 B.n565 585
R675 B.n775 B.n565 585
R676 B.n779 B.n512 585
R677 B.n512 B.n511 585
R678 B.n781 B.n780 585
R679 B.n782 B.n781 585
R680 B.n506 B.n505 585
R681 B.n507 B.n506 585
R682 B.n790 B.n789 585
R683 B.n789 B.n788 585
R684 B.n791 B.n504 585
R685 B.n504 B.n503 585
R686 B.n793 B.n792 585
R687 B.n794 B.n793 585
R688 B.n498 B.n497 585
R689 B.n499 B.n498 585
R690 B.n802 B.n801 585
R691 B.n801 B.n800 585
R692 B.n803 B.n496 585
R693 B.n496 B.n495 585
R694 B.n805 B.n804 585
R695 B.n806 B.n805 585
R696 B.n490 B.n489 585
R697 B.n491 B.n490 585
R698 B.n814 B.n813 585
R699 B.n813 B.n812 585
R700 B.n815 B.n488 585
R701 B.n488 B.n487 585
R702 B.n817 B.n816 585
R703 B.n818 B.n817 585
R704 B.n482 B.n481 585
R705 B.n483 B.n482 585
R706 B.n826 B.n825 585
R707 B.n825 B.n824 585
R708 B.n827 B.n480 585
R709 B.n480 B.n479 585
R710 B.n829 B.n828 585
R711 B.n830 B.n829 585
R712 B.n474 B.n473 585
R713 B.n475 B.n474 585
R714 B.n838 B.n837 585
R715 B.n837 B.n836 585
R716 B.n839 B.n472 585
R717 B.n472 B.n471 585
R718 B.n841 B.n840 585
R719 B.n842 B.n841 585
R720 B.n466 B.n465 585
R721 B.n467 B.n466 585
R722 B.n851 B.n850 585
R723 B.n850 B.n849 585
R724 B.n852 B.n464 585
R725 B.n848 B.n464 585
R726 B.n854 B.n853 585
R727 B.n855 B.n854 585
R728 B.n459 B.n458 585
R729 B.n460 B.n459 585
R730 B.n863 B.n862 585
R731 B.n862 B.n861 585
R732 B.n864 B.n457 585
R733 B.n457 B.n456 585
R734 B.n866 B.n865 585
R735 B.n867 B.n866 585
R736 B.n451 B.n450 585
R737 B.n452 B.n451 585
R738 B.n875 B.n874 585
R739 B.n874 B.n873 585
R740 B.n876 B.n449 585
R741 B.n449 B.n448 585
R742 B.n878 B.n877 585
R743 B.n879 B.n878 585
R744 B.n443 B.n442 585
R745 B.n444 B.n443 585
R746 B.n888 B.n887 585
R747 B.n887 B.n886 585
R748 B.n889 B.n441 585
R749 B.n885 B.n441 585
R750 B.n891 B.n890 585
R751 B.n892 B.n891 585
R752 B.n436 B.n435 585
R753 B.n437 B.n436 585
R754 B.n900 B.n899 585
R755 B.n899 B.n898 585
R756 B.n901 B.n434 585
R757 B.n434 B.n433 585
R758 B.n903 B.n902 585
R759 B.n904 B.n903 585
R760 B.n428 B.n427 585
R761 B.n429 B.n428 585
R762 B.n912 B.n911 585
R763 B.n911 B.n910 585
R764 B.n913 B.n426 585
R765 B.n426 B.n425 585
R766 B.n915 B.n914 585
R767 B.n916 B.n915 585
R768 B.n420 B.n419 585
R769 B.n421 B.n420 585
R770 B.n925 B.n924 585
R771 B.n924 B.n923 585
R772 B.n926 B.n418 585
R773 B.n922 B.n418 585
R774 B.n928 B.n927 585
R775 B.n929 B.n928 585
R776 B.n413 B.n412 585
R777 B.n414 B.n413 585
R778 B.n937 B.n936 585
R779 B.n936 B.n935 585
R780 B.n938 B.n411 585
R781 B.n411 B.n410 585
R782 B.n940 B.n939 585
R783 B.n941 B.n940 585
R784 B.n405 B.n404 585
R785 B.n406 B.n405 585
R786 B.n949 B.n948 585
R787 B.n948 B.n947 585
R788 B.n950 B.n403 585
R789 B.n403 B.n402 585
R790 B.n952 B.n951 585
R791 B.n953 B.n952 585
R792 B.n397 B.n396 585
R793 B.n398 B.n397 585
R794 B.n961 B.n960 585
R795 B.n960 B.n959 585
R796 B.n962 B.n395 585
R797 B.n395 B.n394 585
R798 B.n964 B.n963 585
R799 B.n965 B.n964 585
R800 B.n389 B.n388 585
R801 B.n390 B.n389 585
R802 B.n974 B.n973 585
R803 B.n973 B.n972 585
R804 B.n975 B.n387 585
R805 B.n387 B.n386 585
R806 B.n977 B.n976 585
R807 B.n978 B.n977 585
R808 B.n3 B.n0 585
R809 B.n4 B.n3 585
R810 B.n1206 B.n1 585
R811 B.n1207 B.n1206 585
R812 B.n1205 B.n1204 585
R813 B.n1205 B.n8 585
R814 B.n1203 B.n9 585
R815 B.n12 B.n9 585
R816 B.n1202 B.n1201 585
R817 B.n1201 B.n1200 585
R818 B.n11 B.n10 585
R819 B.n1199 B.n11 585
R820 B.n1197 B.n1196 585
R821 B.n1198 B.n1197 585
R822 B.n1195 B.n17 585
R823 B.n17 B.n16 585
R824 B.n1194 B.n1193 585
R825 B.n1193 B.n1192 585
R826 B.n19 B.n18 585
R827 B.n1191 B.n19 585
R828 B.n1189 B.n1188 585
R829 B.n1190 B.n1189 585
R830 B.n1187 B.n24 585
R831 B.n24 B.n23 585
R832 B.n1186 B.n1185 585
R833 B.n1185 B.n1184 585
R834 B.n26 B.n25 585
R835 B.n1183 B.n26 585
R836 B.n1181 B.n1180 585
R837 B.n1182 B.n1181 585
R838 B.n1179 B.n31 585
R839 B.n31 B.n30 585
R840 B.n1178 B.n1177 585
R841 B.n1177 B.n1176 585
R842 B.n33 B.n32 585
R843 B.n1175 B.n33 585
R844 B.n1173 B.n1172 585
R845 B.n1174 B.n1173 585
R846 B.n1171 B.n37 585
R847 B.n40 B.n37 585
R848 B.n1170 B.n1169 585
R849 B.n1169 B.n1168 585
R850 B.n39 B.n38 585
R851 B.n1167 B.n39 585
R852 B.n1165 B.n1164 585
R853 B.n1166 B.n1165 585
R854 B.n1163 B.n45 585
R855 B.n45 B.n44 585
R856 B.n1162 B.n1161 585
R857 B.n1161 B.n1160 585
R858 B.n47 B.n46 585
R859 B.n1159 B.n47 585
R860 B.n1157 B.n1156 585
R861 B.n1158 B.n1157 585
R862 B.n1155 B.n52 585
R863 B.n52 B.n51 585
R864 B.n1154 B.n1153 585
R865 B.n1153 B.n1152 585
R866 B.n54 B.n53 585
R867 B.n1151 B.n54 585
R868 B.n1149 B.n1148 585
R869 B.n1150 B.n1149 585
R870 B.n1147 B.n58 585
R871 B.n61 B.n58 585
R872 B.n1146 B.n1145 585
R873 B.n1145 B.n1144 585
R874 B.n60 B.n59 585
R875 B.n1143 B.n60 585
R876 B.n1141 B.n1140 585
R877 B.n1142 B.n1141 585
R878 B.n1139 B.n66 585
R879 B.n66 B.n65 585
R880 B.n1138 B.n1137 585
R881 B.n1137 B.n1136 585
R882 B.n68 B.n67 585
R883 B.n1135 B.n68 585
R884 B.n1133 B.n1132 585
R885 B.n1134 B.n1133 585
R886 B.n1131 B.n73 585
R887 B.n73 B.n72 585
R888 B.n1130 B.n1129 585
R889 B.n1129 B.n1128 585
R890 B.n75 B.n74 585
R891 B.n1127 B.n75 585
R892 B.n1125 B.n1124 585
R893 B.n1126 B.n1125 585
R894 B.n1123 B.n79 585
R895 B.n82 B.n79 585
R896 B.n1122 B.n1121 585
R897 B.n1121 B.n1120 585
R898 B.n81 B.n80 585
R899 B.n1119 B.n81 585
R900 B.n1117 B.n1116 585
R901 B.n1118 B.n1117 585
R902 B.n1115 B.n87 585
R903 B.n87 B.n86 585
R904 B.n1114 B.n1113 585
R905 B.n1113 B.n1112 585
R906 B.n89 B.n88 585
R907 B.n1111 B.n89 585
R908 B.n1109 B.n1108 585
R909 B.n1110 B.n1109 585
R910 B.n1107 B.n94 585
R911 B.n94 B.n93 585
R912 B.n1106 B.n1105 585
R913 B.n1105 B.n1104 585
R914 B.n96 B.n95 585
R915 B.n1103 B.n96 585
R916 B.n1101 B.n1100 585
R917 B.n1102 B.n1101 585
R918 B.n1099 B.n101 585
R919 B.n101 B.n100 585
R920 B.n1098 B.n1097 585
R921 B.n1097 B.n1096 585
R922 B.n103 B.n102 585
R923 B.n1095 B.n103 585
R924 B.n1093 B.n1092 585
R925 B.n1094 B.n1093 585
R926 B.n1091 B.n108 585
R927 B.n108 B.n107 585
R928 B.n1090 B.n1089 585
R929 B.n1089 B.n1088 585
R930 B.n110 B.n109 585
R931 B.n1087 B.n110 585
R932 B.n1085 B.n1084 585
R933 B.n1086 B.n1085 585
R934 B.n1083 B.n115 585
R935 B.n115 B.n114 585
R936 B.n1082 B.n1081 585
R937 B.n1081 B.n1080 585
R938 B.n117 B.n116 585
R939 B.n1079 B.n117 585
R940 B.n1077 B.n1076 585
R941 B.n1078 B.n1077 585
R942 B.n1075 B.n122 585
R943 B.n122 B.n121 585
R944 B.n1210 B.n1209 585
R945 B.n1208 B.n2 585
R946 B.n1073 B.n122 530.939
R947 B.n1069 B.n176 530.939
R948 B.n565 B.n510 530.939
R949 B.n777 B.n512 530.939
R950 B.n179 B.t16 299.397
R951 B.n177 B.t12 299.397
R952 B.n570 B.t8 299.397
R953 B.n567 B.t19 299.397
R954 B.n1071 B.n1070 256.663
R955 B.n1071 B.n174 256.663
R956 B.n1071 B.n173 256.663
R957 B.n1071 B.n172 256.663
R958 B.n1071 B.n171 256.663
R959 B.n1071 B.n170 256.663
R960 B.n1071 B.n169 256.663
R961 B.n1071 B.n168 256.663
R962 B.n1071 B.n167 256.663
R963 B.n1071 B.n166 256.663
R964 B.n1071 B.n165 256.663
R965 B.n1071 B.n164 256.663
R966 B.n1071 B.n163 256.663
R967 B.n1071 B.n162 256.663
R968 B.n1071 B.n161 256.663
R969 B.n1071 B.n160 256.663
R970 B.n1071 B.n159 256.663
R971 B.n1071 B.n158 256.663
R972 B.n1071 B.n157 256.663
R973 B.n1071 B.n156 256.663
R974 B.n1071 B.n155 256.663
R975 B.n1071 B.n154 256.663
R976 B.n1071 B.n153 256.663
R977 B.n1071 B.n152 256.663
R978 B.n1071 B.n151 256.663
R979 B.n1071 B.n150 256.663
R980 B.n1071 B.n149 256.663
R981 B.n1071 B.n148 256.663
R982 B.n1071 B.n147 256.663
R983 B.n1071 B.n146 256.663
R984 B.n1071 B.n145 256.663
R985 B.n1071 B.n144 256.663
R986 B.n1071 B.n143 256.663
R987 B.n1071 B.n142 256.663
R988 B.n1071 B.n141 256.663
R989 B.n1071 B.n140 256.663
R990 B.n1071 B.n139 256.663
R991 B.n1071 B.n138 256.663
R992 B.n1071 B.n137 256.663
R993 B.n1071 B.n136 256.663
R994 B.n1071 B.n135 256.663
R995 B.n1071 B.n134 256.663
R996 B.n1071 B.n133 256.663
R997 B.n1071 B.n132 256.663
R998 B.n1071 B.n131 256.663
R999 B.n1071 B.n130 256.663
R1000 B.n1071 B.n129 256.663
R1001 B.n1071 B.n128 256.663
R1002 B.n1071 B.n127 256.663
R1003 B.n1071 B.n126 256.663
R1004 B.n1071 B.n125 256.663
R1005 B.n1072 B.n1071 256.663
R1006 B.n776 B.n775 256.663
R1007 B.n775 B.n515 256.663
R1008 B.n775 B.n516 256.663
R1009 B.n775 B.n517 256.663
R1010 B.n775 B.n518 256.663
R1011 B.n775 B.n519 256.663
R1012 B.n775 B.n520 256.663
R1013 B.n775 B.n521 256.663
R1014 B.n775 B.n522 256.663
R1015 B.n775 B.n523 256.663
R1016 B.n775 B.n524 256.663
R1017 B.n775 B.n525 256.663
R1018 B.n775 B.n526 256.663
R1019 B.n775 B.n527 256.663
R1020 B.n775 B.n528 256.663
R1021 B.n775 B.n529 256.663
R1022 B.n775 B.n530 256.663
R1023 B.n775 B.n531 256.663
R1024 B.n775 B.n532 256.663
R1025 B.n775 B.n533 256.663
R1026 B.n775 B.n534 256.663
R1027 B.n775 B.n535 256.663
R1028 B.n775 B.n536 256.663
R1029 B.n775 B.n537 256.663
R1030 B.n775 B.n538 256.663
R1031 B.n775 B.n539 256.663
R1032 B.n775 B.n540 256.663
R1033 B.n775 B.n541 256.663
R1034 B.n775 B.n542 256.663
R1035 B.n775 B.n543 256.663
R1036 B.n775 B.n544 256.663
R1037 B.n775 B.n545 256.663
R1038 B.n775 B.n546 256.663
R1039 B.n775 B.n547 256.663
R1040 B.n775 B.n548 256.663
R1041 B.n775 B.n549 256.663
R1042 B.n775 B.n550 256.663
R1043 B.n775 B.n551 256.663
R1044 B.n775 B.n552 256.663
R1045 B.n775 B.n553 256.663
R1046 B.n775 B.n554 256.663
R1047 B.n775 B.n555 256.663
R1048 B.n775 B.n556 256.663
R1049 B.n775 B.n557 256.663
R1050 B.n775 B.n558 256.663
R1051 B.n775 B.n559 256.663
R1052 B.n775 B.n560 256.663
R1053 B.n775 B.n561 256.663
R1054 B.n775 B.n562 256.663
R1055 B.n775 B.n563 256.663
R1056 B.n775 B.n564 256.663
R1057 B.n1212 B.n1211 256.663
R1058 B.n181 B.n124 163.367
R1059 B.n185 B.n184 163.367
R1060 B.n189 B.n188 163.367
R1061 B.n193 B.n192 163.367
R1062 B.n197 B.n196 163.367
R1063 B.n201 B.n200 163.367
R1064 B.n205 B.n204 163.367
R1065 B.n209 B.n208 163.367
R1066 B.n213 B.n212 163.367
R1067 B.n217 B.n216 163.367
R1068 B.n221 B.n220 163.367
R1069 B.n225 B.n224 163.367
R1070 B.n229 B.n228 163.367
R1071 B.n233 B.n232 163.367
R1072 B.n237 B.n236 163.367
R1073 B.n241 B.n240 163.367
R1074 B.n245 B.n244 163.367
R1075 B.n249 B.n248 163.367
R1076 B.n253 B.n252 163.367
R1077 B.n257 B.n256 163.367
R1078 B.n261 B.n260 163.367
R1079 B.n265 B.n264 163.367
R1080 B.n269 B.n268 163.367
R1081 B.n274 B.n273 163.367
R1082 B.n278 B.n277 163.367
R1083 B.n282 B.n281 163.367
R1084 B.n286 B.n285 163.367
R1085 B.n290 B.n289 163.367
R1086 B.n295 B.n294 163.367
R1087 B.n299 B.n298 163.367
R1088 B.n303 B.n302 163.367
R1089 B.n307 B.n306 163.367
R1090 B.n311 B.n310 163.367
R1091 B.n315 B.n314 163.367
R1092 B.n319 B.n318 163.367
R1093 B.n323 B.n322 163.367
R1094 B.n327 B.n326 163.367
R1095 B.n331 B.n330 163.367
R1096 B.n335 B.n334 163.367
R1097 B.n339 B.n338 163.367
R1098 B.n343 B.n342 163.367
R1099 B.n347 B.n346 163.367
R1100 B.n351 B.n350 163.367
R1101 B.n355 B.n354 163.367
R1102 B.n359 B.n358 163.367
R1103 B.n363 B.n362 163.367
R1104 B.n367 B.n366 163.367
R1105 B.n371 B.n370 163.367
R1106 B.n375 B.n374 163.367
R1107 B.n379 B.n378 163.367
R1108 B.n381 B.n175 163.367
R1109 B.n783 B.n510 163.367
R1110 B.n783 B.n508 163.367
R1111 B.n787 B.n508 163.367
R1112 B.n787 B.n502 163.367
R1113 B.n795 B.n502 163.367
R1114 B.n795 B.n500 163.367
R1115 B.n799 B.n500 163.367
R1116 B.n799 B.n494 163.367
R1117 B.n807 B.n494 163.367
R1118 B.n807 B.n492 163.367
R1119 B.n811 B.n492 163.367
R1120 B.n811 B.n486 163.367
R1121 B.n819 B.n486 163.367
R1122 B.n819 B.n484 163.367
R1123 B.n823 B.n484 163.367
R1124 B.n823 B.n478 163.367
R1125 B.n831 B.n478 163.367
R1126 B.n831 B.n476 163.367
R1127 B.n835 B.n476 163.367
R1128 B.n835 B.n470 163.367
R1129 B.n843 B.n470 163.367
R1130 B.n843 B.n468 163.367
R1131 B.n847 B.n468 163.367
R1132 B.n847 B.n463 163.367
R1133 B.n856 B.n463 163.367
R1134 B.n856 B.n461 163.367
R1135 B.n860 B.n461 163.367
R1136 B.n860 B.n455 163.367
R1137 B.n868 B.n455 163.367
R1138 B.n868 B.n453 163.367
R1139 B.n872 B.n453 163.367
R1140 B.n872 B.n447 163.367
R1141 B.n880 B.n447 163.367
R1142 B.n880 B.n445 163.367
R1143 B.n884 B.n445 163.367
R1144 B.n884 B.n440 163.367
R1145 B.n893 B.n440 163.367
R1146 B.n893 B.n438 163.367
R1147 B.n897 B.n438 163.367
R1148 B.n897 B.n432 163.367
R1149 B.n905 B.n432 163.367
R1150 B.n905 B.n430 163.367
R1151 B.n909 B.n430 163.367
R1152 B.n909 B.n424 163.367
R1153 B.n917 B.n424 163.367
R1154 B.n917 B.n422 163.367
R1155 B.n921 B.n422 163.367
R1156 B.n921 B.n417 163.367
R1157 B.n930 B.n417 163.367
R1158 B.n930 B.n415 163.367
R1159 B.n934 B.n415 163.367
R1160 B.n934 B.n409 163.367
R1161 B.n942 B.n409 163.367
R1162 B.n942 B.n407 163.367
R1163 B.n946 B.n407 163.367
R1164 B.n946 B.n401 163.367
R1165 B.n954 B.n401 163.367
R1166 B.n954 B.n399 163.367
R1167 B.n958 B.n399 163.367
R1168 B.n958 B.n393 163.367
R1169 B.n966 B.n393 163.367
R1170 B.n966 B.n391 163.367
R1171 B.n971 B.n391 163.367
R1172 B.n971 B.n385 163.367
R1173 B.n979 B.n385 163.367
R1174 B.n980 B.n979 163.367
R1175 B.n980 B.n5 163.367
R1176 B.n6 B.n5 163.367
R1177 B.n7 B.n6 163.367
R1178 B.n986 B.n7 163.367
R1179 B.n987 B.n986 163.367
R1180 B.n987 B.n13 163.367
R1181 B.n14 B.n13 163.367
R1182 B.n15 B.n14 163.367
R1183 B.n992 B.n15 163.367
R1184 B.n992 B.n20 163.367
R1185 B.n21 B.n20 163.367
R1186 B.n22 B.n21 163.367
R1187 B.n997 B.n22 163.367
R1188 B.n997 B.n27 163.367
R1189 B.n28 B.n27 163.367
R1190 B.n29 B.n28 163.367
R1191 B.n1002 B.n29 163.367
R1192 B.n1002 B.n34 163.367
R1193 B.n35 B.n34 163.367
R1194 B.n36 B.n35 163.367
R1195 B.n1007 B.n36 163.367
R1196 B.n1007 B.n41 163.367
R1197 B.n42 B.n41 163.367
R1198 B.n43 B.n42 163.367
R1199 B.n1012 B.n43 163.367
R1200 B.n1012 B.n48 163.367
R1201 B.n49 B.n48 163.367
R1202 B.n50 B.n49 163.367
R1203 B.n1017 B.n50 163.367
R1204 B.n1017 B.n55 163.367
R1205 B.n56 B.n55 163.367
R1206 B.n57 B.n56 163.367
R1207 B.n1022 B.n57 163.367
R1208 B.n1022 B.n62 163.367
R1209 B.n63 B.n62 163.367
R1210 B.n64 B.n63 163.367
R1211 B.n1027 B.n64 163.367
R1212 B.n1027 B.n69 163.367
R1213 B.n70 B.n69 163.367
R1214 B.n71 B.n70 163.367
R1215 B.n1032 B.n71 163.367
R1216 B.n1032 B.n76 163.367
R1217 B.n77 B.n76 163.367
R1218 B.n78 B.n77 163.367
R1219 B.n1037 B.n78 163.367
R1220 B.n1037 B.n83 163.367
R1221 B.n84 B.n83 163.367
R1222 B.n85 B.n84 163.367
R1223 B.n1042 B.n85 163.367
R1224 B.n1042 B.n90 163.367
R1225 B.n91 B.n90 163.367
R1226 B.n92 B.n91 163.367
R1227 B.n1047 B.n92 163.367
R1228 B.n1047 B.n97 163.367
R1229 B.n98 B.n97 163.367
R1230 B.n99 B.n98 163.367
R1231 B.n1052 B.n99 163.367
R1232 B.n1052 B.n104 163.367
R1233 B.n105 B.n104 163.367
R1234 B.n106 B.n105 163.367
R1235 B.n1057 B.n106 163.367
R1236 B.n1057 B.n111 163.367
R1237 B.n112 B.n111 163.367
R1238 B.n113 B.n112 163.367
R1239 B.n1062 B.n113 163.367
R1240 B.n1062 B.n118 163.367
R1241 B.n119 B.n118 163.367
R1242 B.n120 B.n119 163.367
R1243 B.n176 B.n120 163.367
R1244 B.n774 B.n514 163.367
R1245 B.n774 B.n566 163.367
R1246 B.n770 B.n769 163.367
R1247 B.n766 B.n765 163.367
R1248 B.n762 B.n761 163.367
R1249 B.n758 B.n757 163.367
R1250 B.n754 B.n753 163.367
R1251 B.n750 B.n749 163.367
R1252 B.n746 B.n745 163.367
R1253 B.n742 B.n741 163.367
R1254 B.n738 B.n737 163.367
R1255 B.n734 B.n733 163.367
R1256 B.n730 B.n729 163.367
R1257 B.n726 B.n725 163.367
R1258 B.n722 B.n721 163.367
R1259 B.n718 B.n717 163.367
R1260 B.n714 B.n713 163.367
R1261 B.n710 B.n709 163.367
R1262 B.n706 B.n705 163.367
R1263 B.n702 B.n701 163.367
R1264 B.n698 B.n697 163.367
R1265 B.n694 B.n693 163.367
R1266 B.n690 B.n689 163.367
R1267 B.n686 B.n685 163.367
R1268 B.n682 B.n681 163.367
R1269 B.n678 B.n677 163.367
R1270 B.n674 B.n673 163.367
R1271 B.n670 B.n669 163.367
R1272 B.n666 B.n665 163.367
R1273 B.n662 B.n661 163.367
R1274 B.n658 B.n657 163.367
R1275 B.n654 B.n653 163.367
R1276 B.n650 B.n649 163.367
R1277 B.n646 B.n645 163.367
R1278 B.n642 B.n641 163.367
R1279 B.n638 B.n637 163.367
R1280 B.n634 B.n633 163.367
R1281 B.n630 B.n629 163.367
R1282 B.n626 B.n625 163.367
R1283 B.n622 B.n621 163.367
R1284 B.n618 B.n617 163.367
R1285 B.n614 B.n613 163.367
R1286 B.n610 B.n609 163.367
R1287 B.n606 B.n605 163.367
R1288 B.n602 B.n601 163.367
R1289 B.n598 B.n597 163.367
R1290 B.n594 B.n593 163.367
R1291 B.n590 B.n589 163.367
R1292 B.n586 B.n585 163.367
R1293 B.n582 B.n581 163.367
R1294 B.n578 B.n577 163.367
R1295 B.n574 B.n565 163.367
R1296 B.n781 B.n512 163.367
R1297 B.n781 B.n506 163.367
R1298 B.n789 B.n506 163.367
R1299 B.n789 B.n504 163.367
R1300 B.n793 B.n504 163.367
R1301 B.n793 B.n498 163.367
R1302 B.n801 B.n498 163.367
R1303 B.n801 B.n496 163.367
R1304 B.n805 B.n496 163.367
R1305 B.n805 B.n490 163.367
R1306 B.n813 B.n490 163.367
R1307 B.n813 B.n488 163.367
R1308 B.n817 B.n488 163.367
R1309 B.n817 B.n482 163.367
R1310 B.n825 B.n482 163.367
R1311 B.n825 B.n480 163.367
R1312 B.n829 B.n480 163.367
R1313 B.n829 B.n474 163.367
R1314 B.n837 B.n474 163.367
R1315 B.n837 B.n472 163.367
R1316 B.n841 B.n472 163.367
R1317 B.n841 B.n466 163.367
R1318 B.n850 B.n466 163.367
R1319 B.n850 B.n464 163.367
R1320 B.n854 B.n464 163.367
R1321 B.n854 B.n459 163.367
R1322 B.n862 B.n459 163.367
R1323 B.n862 B.n457 163.367
R1324 B.n866 B.n457 163.367
R1325 B.n866 B.n451 163.367
R1326 B.n874 B.n451 163.367
R1327 B.n874 B.n449 163.367
R1328 B.n878 B.n449 163.367
R1329 B.n878 B.n443 163.367
R1330 B.n887 B.n443 163.367
R1331 B.n887 B.n441 163.367
R1332 B.n891 B.n441 163.367
R1333 B.n891 B.n436 163.367
R1334 B.n899 B.n436 163.367
R1335 B.n899 B.n434 163.367
R1336 B.n903 B.n434 163.367
R1337 B.n903 B.n428 163.367
R1338 B.n911 B.n428 163.367
R1339 B.n911 B.n426 163.367
R1340 B.n915 B.n426 163.367
R1341 B.n915 B.n420 163.367
R1342 B.n924 B.n420 163.367
R1343 B.n924 B.n418 163.367
R1344 B.n928 B.n418 163.367
R1345 B.n928 B.n413 163.367
R1346 B.n936 B.n413 163.367
R1347 B.n936 B.n411 163.367
R1348 B.n940 B.n411 163.367
R1349 B.n940 B.n405 163.367
R1350 B.n948 B.n405 163.367
R1351 B.n948 B.n403 163.367
R1352 B.n952 B.n403 163.367
R1353 B.n952 B.n397 163.367
R1354 B.n960 B.n397 163.367
R1355 B.n960 B.n395 163.367
R1356 B.n964 B.n395 163.367
R1357 B.n964 B.n389 163.367
R1358 B.n973 B.n389 163.367
R1359 B.n973 B.n387 163.367
R1360 B.n977 B.n387 163.367
R1361 B.n977 B.n3 163.367
R1362 B.n1210 B.n3 163.367
R1363 B.n1206 B.n2 163.367
R1364 B.n1206 B.n1205 163.367
R1365 B.n1205 B.n9 163.367
R1366 B.n1201 B.n9 163.367
R1367 B.n1201 B.n11 163.367
R1368 B.n1197 B.n11 163.367
R1369 B.n1197 B.n17 163.367
R1370 B.n1193 B.n17 163.367
R1371 B.n1193 B.n19 163.367
R1372 B.n1189 B.n19 163.367
R1373 B.n1189 B.n24 163.367
R1374 B.n1185 B.n24 163.367
R1375 B.n1185 B.n26 163.367
R1376 B.n1181 B.n26 163.367
R1377 B.n1181 B.n31 163.367
R1378 B.n1177 B.n31 163.367
R1379 B.n1177 B.n33 163.367
R1380 B.n1173 B.n33 163.367
R1381 B.n1173 B.n37 163.367
R1382 B.n1169 B.n37 163.367
R1383 B.n1169 B.n39 163.367
R1384 B.n1165 B.n39 163.367
R1385 B.n1165 B.n45 163.367
R1386 B.n1161 B.n45 163.367
R1387 B.n1161 B.n47 163.367
R1388 B.n1157 B.n47 163.367
R1389 B.n1157 B.n52 163.367
R1390 B.n1153 B.n52 163.367
R1391 B.n1153 B.n54 163.367
R1392 B.n1149 B.n54 163.367
R1393 B.n1149 B.n58 163.367
R1394 B.n1145 B.n58 163.367
R1395 B.n1145 B.n60 163.367
R1396 B.n1141 B.n60 163.367
R1397 B.n1141 B.n66 163.367
R1398 B.n1137 B.n66 163.367
R1399 B.n1137 B.n68 163.367
R1400 B.n1133 B.n68 163.367
R1401 B.n1133 B.n73 163.367
R1402 B.n1129 B.n73 163.367
R1403 B.n1129 B.n75 163.367
R1404 B.n1125 B.n75 163.367
R1405 B.n1125 B.n79 163.367
R1406 B.n1121 B.n79 163.367
R1407 B.n1121 B.n81 163.367
R1408 B.n1117 B.n81 163.367
R1409 B.n1117 B.n87 163.367
R1410 B.n1113 B.n87 163.367
R1411 B.n1113 B.n89 163.367
R1412 B.n1109 B.n89 163.367
R1413 B.n1109 B.n94 163.367
R1414 B.n1105 B.n94 163.367
R1415 B.n1105 B.n96 163.367
R1416 B.n1101 B.n96 163.367
R1417 B.n1101 B.n101 163.367
R1418 B.n1097 B.n101 163.367
R1419 B.n1097 B.n103 163.367
R1420 B.n1093 B.n103 163.367
R1421 B.n1093 B.n108 163.367
R1422 B.n1089 B.n108 163.367
R1423 B.n1089 B.n110 163.367
R1424 B.n1085 B.n110 163.367
R1425 B.n1085 B.n115 163.367
R1426 B.n1081 B.n115 163.367
R1427 B.n1081 B.n117 163.367
R1428 B.n1077 B.n117 163.367
R1429 B.n1077 B.n122 163.367
R1430 B.n177 B.t14 152.124
R1431 B.n570 B.t11 152.124
R1432 B.n179 B.t17 152.106
R1433 B.n567 B.t21 152.106
R1434 B.n180 B.n179 78.546
R1435 B.n178 B.n177 78.546
R1436 B.n571 B.n570 78.546
R1437 B.n568 B.n567 78.546
R1438 B.n775 B.n511 77.4047
R1439 B.n1071 B.n121 77.4047
R1440 B.n178 B.t15 73.5779
R1441 B.n571 B.t10 73.5779
R1442 B.n180 B.t18 73.5602
R1443 B.n568 B.t20 73.5602
R1444 B.n1073 B.n1072 71.676
R1445 B.n181 B.n125 71.676
R1446 B.n185 B.n126 71.676
R1447 B.n189 B.n127 71.676
R1448 B.n193 B.n128 71.676
R1449 B.n197 B.n129 71.676
R1450 B.n201 B.n130 71.676
R1451 B.n205 B.n131 71.676
R1452 B.n209 B.n132 71.676
R1453 B.n213 B.n133 71.676
R1454 B.n217 B.n134 71.676
R1455 B.n221 B.n135 71.676
R1456 B.n225 B.n136 71.676
R1457 B.n229 B.n137 71.676
R1458 B.n233 B.n138 71.676
R1459 B.n237 B.n139 71.676
R1460 B.n241 B.n140 71.676
R1461 B.n245 B.n141 71.676
R1462 B.n249 B.n142 71.676
R1463 B.n253 B.n143 71.676
R1464 B.n257 B.n144 71.676
R1465 B.n261 B.n145 71.676
R1466 B.n265 B.n146 71.676
R1467 B.n269 B.n147 71.676
R1468 B.n274 B.n148 71.676
R1469 B.n278 B.n149 71.676
R1470 B.n282 B.n150 71.676
R1471 B.n286 B.n151 71.676
R1472 B.n290 B.n152 71.676
R1473 B.n295 B.n153 71.676
R1474 B.n299 B.n154 71.676
R1475 B.n303 B.n155 71.676
R1476 B.n307 B.n156 71.676
R1477 B.n311 B.n157 71.676
R1478 B.n315 B.n158 71.676
R1479 B.n319 B.n159 71.676
R1480 B.n323 B.n160 71.676
R1481 B.n327 B.n161 71.676
R1482 B.n331 B.n162 71.676
R1483 B.n335 B.n163 71.676
R1484 B.n339 B.n164 71.676
R1485 B.n343 B.n165 71.676
R1486 B.n347 B.n166 71.676
R1487 B.n351 B.n167 71.676
R1488 B.n355 B.n168 71.676
R1489 B.n359 B.n169 71.676
R1490 B.n363 B.n170 71.676
R1491 B.n367 B.n171 71.676
R1492 B.n371 B.n172 71.676
R1493 B.n375 B.n173 71.676
R1494 B.n379 B.n174 71.676
R1495 B.n1070 B.n175 71.676
R1496 B.n1070 B.n1069 71.676
R1497 B.n381 B.n174 71.676
R1498 B.n378 B.n173 71.676
R1499 B.n374 B.n172 71.676
R1500 B.n370 B.n171 71.676
R1501 B.n366 B.n170 71.676
R1502 B.n362 B.n169 71.676
R1503 B.n358 B.n168 71.676
R1504 B.n354 B.n167 71.676
R1505 B.n350 B.n166 71.676
R1506 B.n346 B.n165 71.676
R1507 B.n342 B.n164 71.676
R1508 B.n338 B.n163 71.676
R1509 B.n334 B.n162 71.676
R1510 B.n330 B.n161 71.676
R1511 B.n326 B.n160 71.676
R1512 B.n322 B.n159 71.676
R1513 B.n318 B.n158 71.676
R1514 B.n314 B.n157 71.676
R1515 B.n310 B.n156 71.676
R1516 B.n306 B.n155 71.676
R1517 B.n302 B.n154 71.676
R1518 B.n298 B.n153 71.676
R1519 B.n294 B.n152 71.676
R1520 B.n289 B.n151 71.676
R1521 B.n285 B.n150 71.676
R1522 B.n281 B.n149 71.676
R1523 B.n277 B.n148 71.676
R1524 B.n273 B.n147 71.676
R1525 B.n268 B.n146 71.676
R1526 B.n264 B.n145 71.676
R1527 B.n260 B.n144 71.676
R1528 B.n256 B.n143 71.676
R1529 B.n252 B.n142 71.676
R1530 B.n248 B.n141 71.676
R1531 B.n244 B.n140 71.676
R1532 B.n240 B.n139 71.676
R1533 B.n236 B.n138 71.676
R1534 B.n232 B.n137 71.676
R1535 B.n228 B.n136 71.676
R1536 B.n224 B.n135 71.676
R1537 B.n220 B.n134 71.676
R1538 B.n216 B.n133 71.676
R1539 B.n212 B.n132 71.676
R1540 B.n208 B.n131 71.676
R1541 B.n204 B.n130 71.676
R1542 B.n200 B.n129 71.676
R1543 B.n196 B.n128 71.676
R1544 B.n192 B.n127 71.676
R1545 B.n188 B.n126 71.676
R1546 B.n184 B.n125 71.676
R1547 B.n1072 B.n124 71.676
R1548 B.n777 B.n776 71.676
R1549 B.n566 B.n515 71.676
R1550 B.n769 B.n516 71.676
R1551 B.n765 B.n517 71.676
R1552 B.n761 B.n518 71.676
R1553 B.n757 B.n519 71.676
R1554 B.n753 B.n520 71.676
R1555 B.n749 B.n521 71.676
R1556 B.n745 B.n522 71.676
R1557 B.n741 B.n523 71.676
R1558 B.n737 B.n524 71.676
R1559 B.n733 B.n525 71.676
R1560 B.n729 B.n526 71.676
R1561 B.n725 B.n527 71.676
R1562 B.n721 B.n528 71.676
R1563 B.n717 B.n529 71.676
R1564 B.n713 B.n530 71.676
R1565 B.n709 B.n531 71.676
R1566 B.n705 B.n532 71.676
R1567 B.n701 B.n533 71.676
R1568 B.n697 B.n534 71.676
R1569 B.n693 B.n535 71.676
R1570 B.n689 B.n536 71.676
R1571 B.n685 B.n537 71.676
R1572 B.n681 B.n538 71.676
R1573 B.n677 B.n539 71.676
R1574 B.n673 B.n540 71.676
R1575 B.n669 B.n541 71.676
R1576 B.n665 B.n542 71.676
R1577 B.n661 B.n543 71.676
R1578 B.n657 B.n544 71.676
R1579 B.n653 B.n545 71.676
R1580 B.n649 B.n546 71.676
R1581 B.n645 B.n547 71.676
R1582 B.n641 B.n548 71.676
R1583 B.n637 B.n549 71.676
R1584 B.n633 B.n550 71.676
R1585 B.n629 B.n551 71.676
R1586 B.n625 B.n552 71.676
R1587 B.n621 B.n553 71.676
R1588 B.n617 B.n554 71.676
R1589 B.n613 B.n555 71.676
R1590 B.n609 B.n556 71.676
R1591 B.n605 B.n557 71.676
R1592 B.n601 B.n558 71.676
R1593 B.n597 B.n559 71.676
R1594 B.n593 B.n560 71.676
R1595 B.n589 B.n561 71.676
R1596 B.n585 B.n562 71.676
R1597 B.n581 B.n563 71.676
R1598 B.n577 B.n564 71.676
R1599 B.n776 B.n514 71.676
R1600 B.n770 B.n515 71.676
R1601 B.n766 B.n516 71.676
R1602 B.n762 B.n517 71.676
R1603 B.n758 B.n518 71.676
R1604 B.n754 B.n519 71.676
R1605 B.n750 B.n520 71.676
R1606 B.n746 B.n521 71.676
R1607 B.n742 B.n522 71.676
R1608 B.n738 B.n523 71.676
R1609 B.n734 B.n524 71.676
R1610 B.n730 B.n525 71.676
R1611 B.n726 B.n526 71.676
R1612 B.n722 B.n527 71.676
R1613 B.n718 B.n528 71.676
R1614 B.n714 B.n529 71.676
R1615 B.n710 B.n530 71.676
R1616 B.n706 B.n531 71.676
R1617 B.n702 B.n532 71.676
R1618 B.n698 B.n533 71.676
R1619 B.n694 B.n534 71.676
R1620 B.n690 B.n535 71.676
R1621 B.n686 B.n536 71.676
R1622 B.n682 B.n537 71.676
R1623 B.n678 B.n538 71.676
R1624 B.n674 B.n539 71.676
R1625 B.n670 B.n540 71.676
R1626 B.n666 B.n541 71.676
R1627 B.n662 B.n542 71.676
R1628 B.n658 B.n543 71.676
R1629 B.n654 B.n544 71.676
R1630 B.n650 B.n545 71.676
R1631 B.n646 B.n546 71.676
R1632 B.n642 B.n547 71.676
R1633 B.n638 B.n548 71.676
R1634 B.n634 B.n549 71.676
R1635 B.n630 B.n550 71.676
R1636 B.n626 B.n551 71.676
R1637 B.n622 B.n552 71.676
R1638 B.n618 B.n553 71.676
R1639 B.n614 B.n554 71.676
R1640 B.n610 B.n555 71.676
R1641 B.n606 B.n556 71.676
R1642 B.n602 B.n557 71.676
R1643 B.n598 B.n558 71.676
R1644 B.n594 B.n559 71.676
R1645 B.n590 B.n560 71.676
R1646 B.n586 B.n561 71.676
R1647 B.n582 B.n562 71.676
R1648 B.n578 B.n563 71.676
R1649 B.n574 B.n564 71.676
R1650 B.n1211 B.n1210 71.676
R1651 B.n1211 B.n2 71.676
R1652 B.n271 B.n180 59.5399
R1653 B.n292 B.n178 59.5399
R1654 B.n572 B.n571 59.5399
R1655 B.n569 B.n568 59.5399
R1656 B.n782 B.n511 38.9893
R1657 B.n782 B.n507 38.9893
R1658 B.n788 B.n507 38.9893
R1659 B.n788 B.n503 38.9893
R1660 B.n794 B.n503 38.9893
R1661 B.n794 B.n499 38.9893
R1662 B.n800 B.n499 38.9893
R1663 B.n800 B.n495 38.9893
R1664 B.n806 B.n495 38.9893
R1665 B.n812 B.n491 38.9893
R1666 B.n812 B.n487 38.9893
R1667 B.n818 B.n487 38.9893
R1668 B.n818 B.n483 38.9893
R1669 B.n824 B.n483 38.9893
R1670 B.n824 B.n479 38.9893
R1671 B.n830 B.n479 38.9893
R1672 B.n830 B.n475 38.9893
R1673 B.n836 B.n475 38.9893
R1674 B.n836 B.n471 38.9893
R1675 B.n842 B.n471 38.9893
R1676 B.n842 B.n467 38.9893
R1677 B.n849 B.n467 38.9893
R1678 B.n849 B.n848 38.9893
R1679 B.n855 B.n460 38.9893
R1680 B.n861 B.n460 38.9893
R1681 B.n861 B.n456 38.9893
R1682 B.n867 B.n456 38.9893
R1683 B.n867 B.n452 38.9893
R1684 B.n873 B.n452 38.9893
R1685 B.n873 B.n448 38.9893
R1686 B.n879 B.n448 38.9893
R1687 B.n879 B.n444 38.9893
R1688 B.n886 B.n444 38.9893
R1689 B.n886 B.n885 38.9893
R1690 B.n892 B.n437 38.9893
R1691 B.n898 B.n437 38.9893
R1692 B.n898 B.n433 38.9893
R1693 B.n904 B.n433 38.9893
R1694 B.n904 B.n429 38.9893
R1695 B.n910 B.n429 38.9893
R1696 B.n910 B.n425 38.9893
R1697 B.n916 B.n425 38.9893
R1698 B.n916 B.n421 38.9893
R1699 B.n923 B.n421 38.9893
R1700 B.n923 B.n922 38.9893
R1701 B.n929 B.n414 38.9893
R1702 B.n935 B.n414 38.9893
R1703 B.n935 B.n410 38.9893
R1704 B.n941 B.n410 38.9893
R1705 B.n941 B.n406 38.9893
R1706 B.n947 B.n406 38.9893
R1707 B.n947 B.n402 38.9893
R1708 B.n953 B.n402 38.9893
R1709 B.n953 B.n398 38.9893
R1710 B.n959 B.n398 38.9893
R1711 B.n965 B.n394 38.9893
R1712 B.n965 B.n390 38.9893
R1713 B.n972 B.n390 38.9893
R1714 B.n972 B.n386 38.9893
R1715 B.n978 B.n386 38.9893
R1716 B.n978 B.n4 38.9893
R1717 B.n1209 B.n4 38.9893
R1718 B.n1209 B.n1208 38.9893
R1719 B.n1208 B.n1207 38.9893
R1720 B.n1207 B.n8 38.9893
R1721 B.n12 B.n8 38.9893
R1722 B.n1200 B.n12 38.9893
R1723 B.n1200 B.n1199 38.9893
R1724 B.n1199 B.n1198 38.9893
R1725 B.n1198 B.n16 38.9893
R1726 B.n1192 B.n1191 38.9893
R1727 B.n1191 B.n1190 38.9893
R1728 B.n1190 B.n23 38.9893
R1729 B.n1184 B.n23 38.9893
R1730 B.n1184 B.n1183 38.9893
R1731 B.n1183 B.n1182 38.9893
R1732 B.n1182 B.n30 38.9893
R1733 B.n1176 B.n30 38.9893
R1734 B.n1176 B.n1175 38.9893
R1735 B.n1175 B.n1174 38.9893
R1736 B.n1168 B.n40 38.9893
R1737 B.n1168 B.n1167 38.9893
R1738 B.n1167 B.n1166 38.9893
R1739 B.n1166 B.n44 38.9893
R1740 B.n1160 B.n44 38.9893
R1741 B.n1160 B.n1159 38.9893
R1742 B.n1159 B.n1158 38.9893
R1743 B.n1158 B.n51 38.9893
R1744 B.n1152 B.n51 38.9893
R1745 B.n1152 B.n1151 38.9893
R1746 B.n1151 B.n1150 38.9893
R1747 B.n1144 B.n61 38.9893
R1748 B.n1144 B.n1143 38.9893
R1749 B.n1143 B.n1142 38.9893
R1750 B.n1142 B.n65 38.9893
R1751 B.n1136 B.n65 38.9893
R1752 B.n1136 B.n1135 38.9893
R1753 B.n1135 B.n1134 38.9893
R1754 B.n1134 B.n72 38.9893
R1755 B.n1128 B.n72 38.9893
R1756 B.n1128 B.n1127 38.9893
R1757 B.n1127 B.n1126 38.9893
R1758 B.n1120 B.n82 38.9893
R1759 B.n1120 B.n1119 38.9893
R1760 B.n1119 B.n1118 38.9893
R1761 B.n1118 B.n86 38.9893
R1762 B.n1112 B.n86 38.9893
R1763 B.n1112 B.n1111 38.9893
R1764 B.n1111 B.n1110 38.9893
R1765 B.n1110 B.n93 38.9893
R1766 B.n1104 B.n93 38.9893
R1767 B.n1104 B.n1103 38.9893
R1768 B.n1103 B.n1102 38.9893
R1769 B.n1102 B.n100 38.9893
R1770 B.n1096 B.n100 38.9893
R1771 B.n1096 B.n1095 38.9893
R1772 B.n1094 B.n107 38.9893
R1773 B.n1088 B.n107 38.9893
R1774 B.n1088 B.n1087 38.9893
R1775 B.n1087 B.n1086 38.9893
R1776 B.n1086 B.n114 38.9893
R1777 B.n1080 B.n114 38.9893
R1778 B.n1080 B.n1079 38.9893
R1779 B.n1079 B.n1078 38.9893
R1780 B.n1078 B.n121 38.9893
R1781 B.n929 B.t6 37.8426
R1782 B.n1174 B.t5 37.8426
R1783 B.n959 B.t2 36.6958
R1784 B.n1192 B.t7 36.6958
R1785 B.t9 B.n491 35.5491
R1786 B.n1095 B.t13 35.5491
R1787 B.n779 B.n778 34.4981
R1788 B.n573 B.n509 34.4981
R1789 B.n1068 B.n1067 34.4981
R1790 B.n1075 B.n1074 34.4981
R1791 B.n892 B.t3 34.4024
R1792 B.n1150 B.t4 34.4024
R1793 B.n855 B.t1 30.9622
R1794 B.n1126 B.t0 30.9622
R1795 B B.n1212 18.0485
R1796 B.n780 B.n779 10.6151
R1797 B.n780 B.n505 10.6151
R1798 B.n790 B.n505 10.6151
R1799 B.n791 B.n790 10.6151
R1800 B.n792 B.n791 10.6151
R1801 B.n792 B.n497 10.6151
R1802 B.n802 B.n497 10.6151
R1803 B.n803 B.n802 10.6151
R1804 B.n804 B.n803 10.6151
R1805 B.n804 B.n489 10.6151
R1806 B.n814 B.n489 10.6151
R1807 B.n815 B.n814 10.6151
R1808 B.n816 B.n815 10.6151
R1809 B.n816 B.n481 10.6151
R1810 B.n826 B.n481 10.6151
R1811 B.n827 B.n826 10.6151
R1812 B.n828 B.n827 10.6151
R1813 B.n828 B.n473 10.6151
R1814 B.n838 B.n473 10.6151
R1815 B.n839 B.n838 10.6151
R1816 B.n840 B.n839 10.6151
R1817 B.n840 B.n465 10.6151
R1818 B.n851 B.n465 10.6151
R1819 B.n852 B.n851 10.6151
R1820 B.n853 B.n852 10.6151
R1821 B.n853 B.n458 10.6151
R1822 B.n863 B.n458 10.6151
R1823 B.n864 B.n863 10.6151
R1824 B.n865 B.n864 10.6151
R1825 B.n865 B.n450 10.6151
R1826 B.n875 B.n450 10.6151
R1827 B.n876 B.n875 10.6151
R1828 B.n877 B.n876 10.6151
R1829 B.n877 B.n442 10.6151
R1830 B.n888 B.n442 10.6151
R1831 B.n889 B.n888 10.6151
R1832 B.n890 B.n889 10.6151
R1833 B.n890 B.n435 10.6151
R1834 B.n900 B.n435 10.6151
R1835 B.n901 B.n900 10.6151
R1836 B.n902 B.n901 10.6151
R1837 B.n902 B.n427 10.6151
R1838 B.n912 B.n427 10.6151
R1839 B.n913 B.n912 10.6151
R1840 B.n914 B.n913 10.6151
R1841 B.n914 B.n419 10.6151
R1842 B.n925 B.n419 10.6151
R1843 B.n926 B.n925 10.6151
R1844 B.n927 B.n926 10.6151
R1845 B.n927 B.n412 10.6151
R1846 B.n937 B.n412 10.6151
R1847 B.n938 B.n937 10.6151
R1848 B.n939 B.n938 10.6151
R1849 B.n939 B.n404 10.6151
R1850 B.n949 B.n404 10.6151
R1851 B.n950 B.n949 10.6151
R1852 B.n951 B.n950 10.6151
R1853 B.n951 B.n396 10.6151
R1854 B.n961 B.n396 10.6151
R1855 B.n962 B.n961 10.6151
R1856 B.n963 B.n962 10.6151
R1857 B.n963 B.n388 10.6151
R1858 B.n974 B.n388 10.6151
R1859 B.n975 B.n974 10.6151
R1860 B.n976 B.n975 10.6151
R1861 B.n976 B.n0 10.6151
R1862 B.n778 B.n513 10.6151
R1863 B.n773 B.n513 10.6151
R1864 B.n773 B.n772 10.6151
R1865 B.n772 B.n771 10.6151
R1866 B.n771 B.n768 10.6151
R1867 B.n768 B.n767 10.6151
R1868 B.n767 B.n764 10.6151
R1869 B.n764 B.n763 10.6151
R1870 B.n763 B.n760 10.6151
R1871 B.n760 B.n759 10.6151
R1872 B.n759 B.n756 10.6151
R1873 B.n756 B.n755 10.6151
R1874 B.n755 B.n752 10.6151
R1875 B.n752 B.n751 10.6151
R1876 B.n751 B.n748 10.6151
R1877 B.n748 B.n747 10.6151
R1878 B.n747 B.n744 10.6151
R1879 B.n744 B.n743 10.6151
R1880 B.n743 B.n740 10.6151
R1881 B.n740 B.n739 10.6151
R1882 B.n739 B.n736 10.6151
R1883 B.n736 B.n735 10.6151
R1884 B.n735 B.n732 10.6151
R1885 B.n732 B.n731 10.6151
R1886 B.n731 B.n728 10.6151
R1887 B.n728 B.n727 10.6151
R1888 B.n727 B.n724 10.6151
R1889 B.n724 B.n723 10.6151
R1890 B.n723 B.n720 10.6151
R1891 B.n720 B.n719 10.6151
R1892 B.n719 B.n716 10.6151
R1893 B.n716 B.n715 10.6151
R1894 B.n715 B.n712 10.6151
R1895 B.n712 B.n711 10.6151
R1896 B.n711 B.n708 10.6151
R1897 B.n708 B.n707 10.6151
R1898 B.n707 B.n704 10.6151
R1899 B.n704 B.n703 10.6151
R1900 B.n703 B.n700 10.6151
R1901 B.n700 B.n699 10.6151
R1902 B.n699 B.n696 10.6151
R1903 B.n696 B.n695 10.6151
R1904 B.n695 B.n692 10.6151
R1905 B.n692 B.n691 10.6151
R1906 B.n691 B.n688 10.6151
R1907 B.n688 B.n687 10.6151
R1908 B.n684 B.n683 10.6151
R1909 B.n683 B.n680 10.6151
R1910 B.n680 B.n679 10.6151
R1911 B.n679 B.n676 10.6151
R1912 B.n676 B.n675 10.6151
R1913 B.n675 B.n672 10.6151
R1914 B.n672 B.n671 10.6151
R1915 B.n671 B.n668 10.6151
R1916 B.n668 B.n667 10.6151
R1917 B.n664 B.n663 10.6151
R1918 B.n663 B.n660 10.6151
R1919 B.n660 B.n659 10.6151
R1920 B.n659 B.n656 10.6151
R1921 B.n656 B.n655 10.6151
R1922 B.n655 B.n652 10.6151
R1923 B.n652 B.n651 10.6151
R1924 B.n651 B.n648 10.6151
R1925 B.n648 B.n647 10.6151
R1926 B.n647 B.n644 10.6151
R1927 B.n644 B.n643 10.6151
R1928 B.n643 B.n640 10.6151
R1929 B.n640 B.n639 10.6151
R1930 B.n639 B.n636 10.6151
R1931 B.n636 B.n635 10.6151
R1932 B.n635 B.n632 10.6151
R1933 B.n632 B.n631 10.6151
R1934 B.n631 B.n628 10.6151
R1935 B.n628 B.n627 10.6151
R1936 B.n627 B.n624 10.6151
R1937 B.n624 B.n623 10.6151
R1938 B.n623 B.n620 10.6151
R1939 B.n620 B.n619 10.6151
R1940 B.n619 B.n616 10.6151
R1941 B.n616 B.n615 10.6151
R1942 B.n615 B.n612 10.6151
R1943 B.n612 B.n611 10.6151
R1944 B.n611 B.n608 10.6151
R1945 B.n608 B.n607 10.6151
R1946 B.n607 B.n604 10.6151
R1947 B.n604 B.n603 10.6151
R1948 B.n603 B.n600 10.6151
R1949 B.n600 B.n599 10.6151
R1950 B.n599 B.n596 10.6151
R1951 B.n596 B.n595 10.6151
R1952 B.n595 B.n592 10.6151
R1953 B.n592 B.n591 10.6151
R1954 B.n591 B.n588 10.6151
R1955 B.n588 B.n587 10.6151
R1956 B.n587 B.n584 10.6151
R1957 B.n584 B.n583 10.6151
R1958 B.n583 B.n580 10.6151
R1959 B.n580 B.n579 10.6151
R1960 B.n579 B.n576 10.6151
R1961 B.n576 B.n575 10.6151
R1962 B.n575 B.n573 10.6151
R1963 B.n784 B.n509 10.6151
R1964 B.n785 B.n784 10.6151
R1965 B.n786 B.n785 10.6151
R1966 B.n786 B.n501 10.6151
R1967 B.n796 B.n501 10.6151
R1968 B.n797 B.n796 10.6151
R1969 B.n798 B.n797 10.6151
R1970 B.n798 B.n493 10.6151
R1971 B.n808 B.n493 10.6151
R1972 B.n809 B.n808 10.6151
R1973 B.n810 B.n809 10.6151
R1974 B.n810 B.n485 10.6151
R1975 B.n820 B.n485 10.6151
R1976 B.n821 B.n820 10.6151
R1977 B.n822 B.n821 10.6151
R1978 B.n822 B.n477 10.6151
R1979 B.n832 B.n477 10.6151
R1980 B.n833 B.n832 10.6151
R1981 B.n834 B.n833 10.6151
R1982 B.n834 B.n469 10.6151
R1983 B.n844 B.n469 10.6151
R1984 B.n845 B.n844 10.6151
R1985 B.n846 B.n845 10.6151
R1986 B.n846 B.n462 10.6151
R1987 B.n857 B.n462 10.6151
R1988 B.n858 B.n857 10.6151
R1989 B.n859 B.n858 10.6151
R1990 B.n859 B.n454 10.6151
R1991 B.n869 B.n454 10.6151
R1992 B.n870 B.n869 10.6151
R1993 B.n871 B.n870 10.6151
R1994 B.n871 B.n446 10.6151
R1995 B.n881 B.n446 10.6151
R1996 B.n882 B.n881 10.6151
R1997 B.n883 B.n882 10.6151
R1998 B.n883 B.n439 10.6151
R1999 B.n894 B.n439 10.6151
R2000 B.n895 B.n894 10.6151
R2001 B.n896 B.n895 10.6151
R2002 B.n896 B.n431 10.6151
R2003 B.n906 B.n431 10.6151
R2004 B.n907 B.n906 10.6151
R2005 B.n908 B.n907 10.6151
R2006 B.n908 B.n423 10.6151
R2007 B.n918 B.n423 10.6151
R2008 B.n919 B.n918 10.6151
R2009 B.n920 B.n919 10.6151
R2010 B.n920 B.n416 10.6151
R2011 B.n931 B.n416 10.6151
R2012 B.n932 B.n931 10.6151
R2013 B.n933 B.n932 10.6151
R2014 B.n933 B.n408 10.6151
R2015 B.n943 B.n408 10.6151
R2016 B.n944 B.n943 10.6151
R2017 B.n945 B.n944 10.6151
R2018 B.n945 B.n400 10.6151
R2019 B.n955 B.n400 10.6151
R2020 B.n956 B.n955 10.6151
R2021 B.n957 B.n956 10.6151
R2022 B.n957 B.n392 10.6151
R2023 B.n967 B.n392 10.6151
R2024 B.n968 B.n967 10.6151
R2025 B.n970 B.n968 10.6151
R2026 B.n970 B.n969 10.6151
R2027 B.n969 B.n384 10.6151
R2028 B.n981 B.n384 10.6151
R2029 B.n982 B.n981 10.6151
R2030 B.n983 B.n982 10.6151
R2031 B.n984 B.n983 10.6151
R2032 B.n985 B.n984 10.6151
R2033 B.n988 B.n985 10.6151
R2034 B.n989 B.n988 10.6151
R2035 B.n990 B.n989 10.6151
R2036 B.n991 B.n990 10.6151
R2037 B.n993 B.n991 10.6151
R2038 B.n994 B.n993 10.6151
R2039 B.n995 B.n994 10.6151
R2040 B.n996 B.n995 10.6151
R2041 B.n998 B.n996 10.6151
R2042 B.n999 B.n998 10.6151
R2043 B.n1000 B.n999 10.6151
R2044 B.n1001 B.n1000 10.6151
R2045 B.n1003 B.n1001 10.6151
R2046 B.n1004 B.n1003 10.6151
R2047 B.n1005 B.n1004 10.6151
R2048 B.n1006 B.n1005 10.6151
R2049 B.n1008 B.n1006 10.6151
R2050 B.n1009 B.n1008 10.6151
R2051 B.n1010 B.n1009 10.6151
R2052 B.n1011 B.n1010 10.6151
R2053 B.n1013 B.n1011 10.6151
R2054 B.n1014 B.n1013 10.6151
R2055 B.n1015 B.n1014 10.6151
R2056 B.n1016 B.n1015 10.6151
R2057 B.n1018 B.n1016 10.6151
R2058 B.n1019 B.n1018 10.6151
R2059 B.n1020 B.n1019 10.6151
R2060 B.n1021 B.n1020 10.6151
R2061 B.n1023 B.n1021 10.6151
R2062 B.n1024 B.n1023 10.6151
R2063 B.n1025 B.n1024 10.6151
R2064 B.n1026 B.n1025 10.6151
R2065 B.n1028 B.n1026 10.6151
R2066 B.n1029 B.n1028 10.6151
R2067 B.n1030 B.n1029 10.6151
R2068 B.n1031 B.n1030 10.6151
R2069 B.n1033 B.n1031 10.6151
R2070 B.n1034 B.n1033 10.6151
R2071 B.n1035 B.n1034 10.6151
R2072 B.n1036 B.n1035 10.6151
R2073 B.n1038 B.n1036 10.6151
R2074 B.n1039 B.n1038 10.6151
R2075 B.n1040 B.n1039 10.6151
R2076 B.n1041 B.n1040 10.6151
R2077 B.n1043 B.n1041 10.6151
R2078 B.n1044 B.n1043 10.6151
R2079 B.n1045 B.n1044 10.6151
R2080 B.n1046 B.n1045 10.6151
R2081 B.n1048 B.n1046 10.6151
R2082 B.n1049 B.n1048 10.6151
R2083 B.n1050 B.n1049 10.6151
R2084 B.n1051 B.n1050 10.6151
R2085 B.n1053 B.n1051 10.6151
R2086 B.n1054 B.n1053 10.6151
R2087 B.n1055 B.n1054 10.6151
R2088 B.n1056 B.n1055 10.6151
R2089 B.n1058 B.n1056 10.6151
R2090 B.n1059 B.n1058 10.6151
R2091 B.n1060 B.n1059 10.6151
R2092 B.n1061 B.n1060 10.6151
R2093 B.n1063 B.n1061 10.6151
R2094 B.n1064 B.n1063 10.6151
R2095 B.n1065 B.n1064 10.6151
R2096 B.n1066 B.n1065 10.6151
R2097 B.n1067 B.n1066 10.6151
R2098 B.n1204 B.n1 10.6151
R2099 B.n1204 B.n1203 10.6151
R2100 B.n1203 B.n1202 10.6151
R2101 B.n1202 B.n10 10.6151
R2102 B.n1196 B.n10 10.6151
R2103 B.n1196 B.n1195 10.6151
R2104 B.n1195 B.n1194 10.6151
R2105 B.n1194 B.n18 10.6151
R2106 B.n1188 B.n18 10.6151
R2107 B.n1188 B.n1187 10.6151
R2108 B.n1187 B.n1186 10.6151
R2109 B.n1186 B.n25 10.6151
R2110 B.n1180 B.n25 10.6151
R2111 B.n1180 B.n1179 10.6151
R2112 B.n1179 B.n1178 10.6151
R2113 B.n1178 B.n32 10.6151
R2114 B.n1172 B.n32 10.6151
R2115 B.n1172 B.n1171 10.6151
R2116 B.n1171 B.n1170 10.6151
R2117 B.n1170 B.n38 10.6151
R2118 B.n1164 B.n38 10.6151
R2119 B.n1164 B.n1163 10.6151
R2120 B.n1163 B.n1162 10.6151
R2121 B.n1162 B.n46 10.6151
R2122 B.n1156 B.n46 10.6151
R2123 B.n1156 B.n1155 10.6151
R2124 B.n1155 B.n1154 10.6151
R2125 B.n1154 B.n53 10.6151
R2126 B.n1148 B.n53 10.6151
R2127 B.n1148 B.n1147 10.6151
R2128 B.n1147 B.n1146 10.6151
R2129 B.n1146 B.n59 10.6151
R2130 B.n1140 B.n59 10.6151
R2131 B.n1140 B.n1139 10.6151
R2132 B.n1139 B.n1138 10.6151
R2133 B.n1138 B.n67 10.6151
R2134 B.n1132 B.n67 10.6151
R2135 B.n1132 B.n1131 10.6151
R2136 B.n1131 B.n1130 10.6151
R2137 B.n1130 B.n74 10.6151
R2138 B.n1124 B.n74 10.6151
R2139 B.n1124 B.n1123 10.6151
R2140 B.n1123 B.n1122 10.6151
R2141 B.n1122 B.n80 10.6151
R2142 B.n1116 B.n80 10.6151
R2143 B.n1116 B.n1115 10.6151
R2144 B.n1115 B.n1114 10.6151
R2145 B.n1114 B.n88 10.6151
R2146 B.n1108 B.n88 10.6151
R2147 B.n1108 B.n1107 10.6151
R2148 B.n1107 B.n1106 10.6151
R2149 B.n1106 B.n95 10.6151
R2150 B.n1100 B.n95 10.6151
R2151 B.n1100 B.n1099 10.6151
R2152 B.n1099 B.n1098 10.6151
R2153 B.n1098 B.n102 10.6151
R2154 B.n1092 B.n102 10.6151
R2155 B.n1092 B.n1091 10.6151
R2156 B.n1091 B.n1090 10.6151
R2157 B.n1090 B.n109 10.6151
R2158 B.n1084 B.n109 10.6151
R2159 B.n1084 B.n1083 10.6151
R2160 B.n1083 B.n1082 10.6151
R2161 B.n1082 B.n116 10.6151
R2162 B.n1076 B.n116 10.6151
R2163 B.n1076 B.n1075 10.6151
R2164 B.n1074 B.n123 10.6151
R2165 B.n182 B.n123 10.6151
R2166 B.n183 B.n182 10.6151
R2167 B.n186 B.n183 10.6151
R2168 B.n187 B.n186 10.6151
R2169 B.n190 B.n187 10.6151
R2170 B.n191 B.n190 10.6151
R2171 B.n194 B.n191 10.6151
R2172 B.n195 B.n194 10.6151
R2173 B.n198 B.n195 10.6151
R2174 B.n199 B.n198 10.6151
R2175 B.n202 B.n199 10.6151
R2176 B.n203 B.n202 10.6151
R2177 B.n206 B.n203 10.6151
R2178 B.n207 B.n206 10.6151
R2179 B.n210 B.n207 10.6151
R2180 B.n211 B.n210 10.6151
R2181 B.n214 B.n211 10.6151
R2182 B.n215 B.n214 10.6151
R2183 B.n218 B.n215 10.6151
R2184 B.n219 B.n218 10.6151
R2185 B.n222 B.n219 10.6151
R2186 B.n223 B.n222 10.6151
R2187 B.n226 B.n223 10.6151
R2188 B.n227 B.n226 10.6151
R2189 B.n230 B.n227 10.6151
R2190 B.n231 B.n230 10.6151
R2191 B.n234 B.n231 10.6151
R2192 B.n235 B.n234 10.6151
R2193 B.n238 B.n235 10.6151
R2194 B.n239 B.n238 10.6151
R2195 B.n242 B.n239 10.6151
R2196 B.n243 B.n242 10.6151
R2197 B.n246 B.n243 10.6151
R2198 B.n247 B.n246 10.6151
R2199 B.n250 B.n247 10.6151
R2200 B.n251 B.n250 10.6151
R2201 B.n254 B.n251 10.6151
R2202 B.n255 B.n254 10.6151
R2203 B.n258 B.n255 10.6151
R2204 B.n259 B.n258 10.6151
R2205 B.n262 B.n259 10.6151
R2206 B.n263 B.n262 10.6151
R2207 B.n266 B.n263 10.6151
R2208 B.n267 B.n266 10.6151
R2209 B.n270 B.n267 10.6151
R2210 B.n275 B.n272 10.6151
R2211 B.n276 B.n275 10.6151
R2212 B.n279 B.n276 10.6151
R2213 B.n280 B.n279 10.6151
R2214 B.n283 B.n280 10.6151
R2215 B.n284 B.n283 10.6151
R2216 B.n287 B.n284 10.6151
R2217 B.n288 B.n287 10.6151
R2218 B.n291 B.n288 10.6151
R2219 B.n296 B.n293 10.6151
R2220 B.n297 B.n296 10.6151
R2221 B.n300 B.n297 10.6151
R2222 B.n301 B.n300 10.6151
R2223 B.n304 B.n301 10.6151
R2224 B.n305 B.n304 10.6151
R2225 B.n308 B.n305 10.6151
R2226 B.n309 B.n308 10.6151
R2227 B.n312 B.n309 10.6151
R2228 B.n313 B.n312 10.6151
R2229 B.n316 B.n313 10.6151
R2230 B.n317 B.n316 10.6151
R2231 B.n320 B.n317 10.6151
R2232 B.n321 B.n320 10.6151
R2233 B.n324 B.n321 10.6151
R2234 B.n325 B.n324 10.6151
R2235 B.n328 B.n325 10.6151
R2236 B.n329 B.n328 10.6151
R2237 B.n332 B.n329 10.6151
R2238 B.n333 B.n332 10.6151
R2239 B.n336 B.n333 10.6151
R2240 B.n337 B.n336 10.6151
R2241 B.n340 B.n337 10.6151
R2242 B.n341 B.n340 10.6151
R2243 B.n344 B.n341 10.6151
R2244 B.n345 B.n344 10.6151
R2245 B.n348 B.n345 10.6151
R2246 B.n349 B.n348 10.6151
R2247 B.n352 B.n349 10.6151
R2248 B.n353 B.n352 10.6151
R2249 B.n356 B.n353 10.6151
R2250 B.n357 B.n356 10.6151
R2251 B.n360 B.n357 10.6151
R2252 B.n361 B.n360 10.6151
R2253 B.n364 B.n361 10.6151
R2254 B.n365 B.n364 10.6151
R2255 B.n368 B.n365 10.6151
R2256 B.n369 B.n368 10.6151
R2257 B.n372 B.n369 10.6151
R2258 B.n373 B.n372 10.6151
R2259 B.n376 B.n373 10.6151
R2260 B.n377 B.n376 10.6151
R2261 B.n380 B.n377 10.6151
R2262 B.n382 B.n380 10.6151
R2263 B.n383 B.n382 10.6151
R2264 B.n1068 B.n383 10.6151
R2265 B.n687 B.n569 9.36635
R2266 B.n664 B.n572 9.36635
R2267 B.n271 B.n270 9.36635
R2268 B.n293 B.n292 9.36635
R2269 B.n1212 B.n0 8.11757
R2270 B.n1212 B.n1 8.11757
R2271 B.n848 B.t1 8.0276
R2272 B.n82 B.t0 8.0276
R2273 B.n885 B.t3 4.58742
R2274 B.n61 B.t4 4.58742
R2275 B.n806 B.t9 3.44069
R2276 B.t13 B.n1094 3.44069
R2277 B.t2 B.n394 2.29396
R2278 B.t7 B.n16 2.29396
R2279 B.n684 B.n569 1.24928
R2280 B.n667 B.n572 1.24928
R2281 B.n272 B.n271 1.24928
R2282 B.n292 B.n291 1.24928
R2283 B.n922 B.t6 1.14723
R2284 B.n40 B.t5 1.14723
R2285 VN.n76 VN.n75 161.3
R2286 VN.n74 VN.n40 161.3
R2287 VN.n73 VN.n72 161.3
R2288 VN.n71 VN.n41 161.3
R2289 VN.n70 VN.n69 161.3
R2290 VN.n68 VN.n42 161.3
R2291 VN.n67 VN.n66 161.3
R2292 VN.n65 VN.n43 161.3
R2293 VN.n64 VN.n63 161.3
R2294 VN.n62 VN.n44 161.3
R2295 VN.n61 VN.n60 161.3
R2296 VN.n59 VN.n46 161.3
R2297 VN.n58 VN.n57 161.3
R2298 VN.n56 VN.n47 161.3
R2299 VN.n55 VN.n54 161.3
R2300 VN.n53 VN.n48 161.3
R2301 VN.n52 VN.n51 161.3
R2302 VN.n37 VN.n36 161.3
R2303 VN.n35 VN.n1 161.3
R2304 VN.n34 VN.n33 161.3
R2305 VN.n32 VN.n2 161.3
R2306 VN.n31 VN.n30 161.3
R2307 VN.n29 VN.n3 161.3
R2308 VN.n28 VN.n27 161.3
R2309 VN.n26 VN.n4 161.3
R2310 VN.n25 VN.n24 161.3
R2311 VN.n22 VN.n5 161.3
R2312 VN.n21 VN.n20 161.3
R2313 VN.n19 VN.n6 161.3
R2314 VN.n18 VN.n17 161.3
R2315 VN.n16 VN.n7 161.3
R2316 VN.n15 VN.n14 161.3
R2317 VN.n13 VN.n8 161.3
R2318 VN.n12 VN.n11 161.3
R2319 VN.n49 VN.t4 122.177
R2320 VN.n9 VN.t2 122.177
R2321 VN.n10 VN.t1 90.1164
R2322 VN.n23 VN.t6 90.1164
R2323 VN.n0 VN.t5 90.1164
R2324 VN.n50 VN.t7 90.1164
R2325 VN.n45 VN.t0 90.1164
R2326 VN.n39 VN.t3 90.1164
R2327 VN.n38 VN.n0 86.3974
R2328 VN.n77 VN.n39 86.3974
R2329 VN.n50 VN.n49 73.7323
R2330 VN.n10 VN.n9 73.7323
R2331 VN VN.n77 57.7935
R2332 VN.n30 VN.n2 45.3497
R2333 VN.n69 VN.n41 45.3497
R2334 VN.n17 VN.n16 40.4934
R2335 VN.n17 VN.n6 40.4934
R2336 VN.n57 VN.n56 40.4934
R2337 VN.n57 VN.n46 40.4934
R2338 VN.n30 VN.n29 35.6371
R2339 VN.n69 VN.n68 35.6371
R2340 VN.n11 VN.n8 24.4675
R2341 VN.n15 VN.n8 24.4675
R2342 VN.n16 VN.n15 24.4675
R2343 VN.n21 VN.n6 24.4675
R2344 VN.n22 VN.n21 24.4675
R2345 VN.n24 VN.n22 24.4675
R2346 VN.n28 VN.n4 24.4675
R2347 VN.n29 VN.n28 24.4675
R2348 VN.n34 VN.n2 24.4675
R2349 VN.n35 VN.n34 24.4675
R2350 VN.n36 VN.n35 24.4675
R2351 VN.n56 VN.n55 24.4675
R2352 VN.n55 VN.n48 24.4675
R2353 VN.n51 VN.n48 24.4675
R2354 VN.n68 VN.n67 24.4675
R2355 VN.n67 VN.n43 24.4675
R2356 VN.n63 VN.n62 24.4675
R2357 VN.n62 VN.n61 24.4675
R2358 VN.n61 VN.n46 24.4675
R2359 VN.n75 VN.n74 24.4675
R2360 VN.n74 VN.n73 24.4675
R2361 VN.n73 VN.n41 24.4675
R2362 VN.n23 VN.n4 23.2442
R2363 VN.n45 VN.n43 23.2442
R2364 VN.n36 VN.n0 3.67055
R2365 VN.n75 VN.n39 3.67055
R2366 VN.n52 VN.n49 3.35319
R2367 VN.n12 VN.n9 3.35319
R2368 VN.n11 VN.n10 1.22385
R2369 VN.n24 VN.n23 1.22385
R2370 VN.n51 VN.n50 1.22385
R2371 VN.n63 VN.n45 1.22385
R2372 VN.n77 VN.n76 0.354971
R2373 VN.n38 VN.n37 0.354971
R2374 VN VN.n38 0.26696
R2375 VN.n76 VN.n40 0.189894
R2376 VN.n72 VN.n40 0.189894
R2377 VN.n72 VN.n71 0.189894
R2378 VN.n71 VN.n70 0.189894
R2379 VN.n70 VN.n42 0.189894
R2380 VN.n66 VN.n42 0.189894
R2381 VN.n66 VN.n65 0.189894
R2382 VN.n65 VN.n64 0.189894
R2383 VN.n64 VN.n44 0.189894
R2384 VN.n60 VN.n44 0.189894
R2385 VN.n60 VN.n59 0.189894
R2386 VN.n59 VN.n58 0.189894
R2387 VN.n58 VN.n47 0.189894
R2388 VN.n54 VN.n47 0.189894
R2389 VN.n54 VN.n53 0.189894
R2390 VN.n53 VN.n52 0.189894
R2391 VN.n13 VN.n12 0.189894
R2392 VN.n14 VN.n13 0.189894
R2393 VN.n14 VN.n7 0.189894
R2394 VN.n18 VN.n7 0.189894
R2395 VN.n19 VN.n18 0.189894
R2396 VN.n20 VN.n19 0.189894
R2397 VN.n20 VN.n5 0.189894
R2398 VN.n25 VN.n5 0.189894
R2399 VN.n26 VN.n25 0.189894
R2400 VN.n27 VN.n26 0.189894
R2401 VN.n27 VN.n3 0.189894
R2402 VN.n31 VN.n3 0.189894
R2403 VN.n32 VN.n31 0.189894
R2404 VN.n33 VN.n32 0.189894
R2405 VN.n33 VN.n1 0.189894
R2406 VN.n37 VN.n1 0.189894
R2407 VDD2.n2 VDD2.n1 62.9847
R2408 VDD2.n2 VDD2.n0 62.9847
R2409 VDD2 VDD2.n5 62.9819
R2410 VDD2.n4 VDD2.n3 61.2944
R2411 VDD2.n4 VDD2.n2 51.4179
R2412 VDD2 VDD2.n4 1.80438
R2413 VDD2.n5 VDD2.t0 1.42394
R2414 VDD2.n5 VDD2.t3 1.42394
R2415 VDD2.n3 VDD2.t4 1.42394
R2416 VDD2.n3 VDD2.t7 1.42394
R2417 VDD2.n1 VDD2.t1 1.42394
R2418 VDD2.n1 VDD2.t2 1.42394
R2419 VDD2.n0 VDD2.t5 1.42394
R2420 VDD2.n0 VDD2.t6 1.42394
C0 VN VTAIL 11.308701f
C1 VN VDD2 10.6301f
C2 VP VN 9.387879f
C3 VN VDD1 0.153473f
C4 VTAIL VDD2 9.15276f
C5 VP VTAIL 11.322801f
C6 VTAIL VDD1 9.09083f
C7 VP VDD2 0.638571f
C8 VDD1 VDD2 2.35657f
C9 VP VDD1 11.1132f
C10 VDD2 B 6.665161f
C11 VDD1 B 7.222494f
C12 VTAIL B 12.38758f
C13 VN B 19.97461f
C14 VP B 18.622849f
C15 VDD2.t5 B 0.296637f
C16 VDD2.t6 B 0.296637f
C17 VDD2.n0 B 2.68323f
C18 VDD2.t1 B 0.296637f
C19 VDD2.t2 B 0.296637f
C20 VDD2.n1 B 2.68323f
C21 VDD2.n2 B 4.37535f
C22 VDD2.t4 B 0.296637f
C23 VDD2.t7 B 0.296637f
C24 VDD2.n3 B 2.66476f
C25 VDD2.n4 B 3.76434f
C26 VDD2.t0 B 0.296637f
C27 VDD2.t3 B 0.296637f
C28 VDD2.n5 B 2.68318f
C29 VN.t5 B 2.42458f
C30 VN.n0 B 0.907519f
C31 VN.n1 B 0.01713f
C32 VN.n2 B 0.032941f
C33 VN.n3 B 0.01713f
C34 VN.n4 B 0.031137f
C35 VN.n5 B 0.01713f
C36 VN.n6 B 0.034046f
C37 VN.n7 B 0.01713f
C38 VN.n8 B 0.031926f
C39 VN.t2 B 2.68035f
C40 VN.n9 B 0.857436f
C41 VN.t1 B 2.42458f
C42 VN.n10 B 0.898331f
C43 VN.n11 B 0.016951f
C44 VN.n12 B 0.217989f
C45 VN.n13 B 0.01713f
C46 VN.n14 B 0.01713f
C47 VN.n15 B 0.031926f
C48 VN.n16 B 0.034046f
C49 VN.n17 B 0.013848f
C50 VN.n18 B 0.01713f
C51 VN.n19 B 0.01713f
C52 VN.n20 B 0.01713f
C53 VN.n21 B 0.031926f
C54 VN.n22 B 0.031926f
C55 VN.t6 B 2.42458f
C56 VN.n23 B 0.843798f
C57 VN.n24 B 0.016951f
C58 VN.n25 B 0.01713f
C59 VN.n26 B 0.01713f
C60 VN.n27 B 0.01713f
C61 VN.n28 B 0.031926f
C62 VN.n29 B 0.034593f
C63 VN.n30 B 0.014406f
C64 VN.n31 B 0.01713f
C65 VN.n32 B 0.01713f
C66 VN.n33 B 0.01713f
C67 VN.n34 B 0.031926f
C68 VN.n35 B 0.031926f
C69 VN.n36 B 0.018528f
C70 VN.n37 B 0.027648f
C71 VN.n38 B 0.051468f
C72 VN.t3 B 2.42458f
C73 VN.n39 B 0.907519f
C74 VN.n40 B 0.01713f
C75 VN.n41 B 0.032941f
C76 VN.n42 B 0.01713f
C77 VN.n43 B 0.031137f
C78 VN.n44 B 0.01713f
C79 VN.t0 B 2.42458f
C80 VN.n45 B 0.843798f
C81 VN.n46 B 0.034046f
C82 VN.n47 B 0.01713f
C83 VN.n48 B 0.031926f
C84 VN.t4 B 2.68035f
C85 VN.n49 B 0.857436f
C86 VN.t7 B 2.42458f
C87 VN.n50 B 0.898331f
C88 VN.n51 B 0.016951f
C89 VN.n52 B 0.217989f
C90 VN.n53 B 0.01713f
C91 VN.n54 B 0.01713f
C92 VN.n55 B 0.031926f
C93 VN.n56 B 0.034046f
C94 VN.n57 B 0.013848f
C95 VN.n58 B 0.01713f
C96 VN.n59 B 0.01713f
C97 VN.n60 B 0.01713f
C98 VN.n61 B 0.031926f
C99 VN.n62 B 0.031926f
C100 VN.n63 B 0.016951f
C101 VN.n64 B 0.01713f
C102 VN.n65 B 0.01713f
C103 VN.n66 B 0.01713f
C104 VN.n67 B 0.031926f
C105 VN.n68 B 0.034593f
C106 VN.n69 B 0.014406f
C107 VN.n70 B 0.01713f
C108 VN.n71 B 0.01713f
C109 VN.n72 B 0.01713f
C110 VN.n73 B 0.031926f
C111 VN.n74 B 0.031926f
C112 VN.n75 B 0.018528f
C113 VN.n76 B 0.027648f
C114 VN.n77 B 1.20459f
C115 VTAIL.t5 B 0.220702f
C116 VTAIL.t4 B 0.220702f
C117 VTAIL.n0 B 1.92106f
C118 VTAIL.n1 B 0.432396f
C119 VTAIL.t15 B 2.45178f
C120 VTAIL.n2 B 0.530221f
C121 VTAIL.t7 B 2.45178f
C122 VTAIL.n3 B 0.530221f
C123 VTAIL.t8 B 0.220702f
C124 VTAIL.t14 B 0.220702f
C125 VTAIL.n4 B 1.92106f
C126 VTAIL.n5 B 0.654511f
C127 VTAIL.t10 B 2.45178f
C128 VTAIL.n6 B 1.77424f
C129 VTAIL.t1 B 2.4518f
C130 VTAIL.n7 B 1.77423f
C131 VTAIL.t3 B 0.220702f
C132 VTAIL.t6 B 0.220702f
C133 VTAIL.n8 B 1.92106f
C134 VTAIL.n9 B 0.654512f
C135 VTAIL.t2 B 2.4518f
C136 VTAIL.n10 B 0.530207f
C137 VTAIL.t13 B 2.4518f
C138 VTAIL.n11 B 0.530207f
C139 VTAIL.t12 B 0.220702f
C140 VTAIL.t11 B 0.220702f
C141 VTAIL.n12 B 1.92106f
C142 VTAIL.n13 B 0.654512f
C143 VTAIL.t9 B 2.45179f
C144 VTAIL.n14 B 1.77423f
C145 VTAIL.t0 B 2.45178f
C146 VTAIL.n15 B 1.77048f
C147 VDD1.t1 B 0.300632f
C148 VDD1.t0 B 0.300632f
C149 VDD1.n0 B 2.72086f
C150 VDD1.t6 B 0.300632f
C151 VDD1.t2 B 0.300632f
C152 VDD1.n1 B 2.71937f
C153 VDD1.t4 B 0.300632f
C154 VDD1.t5 B 0.300632f
C155 VDD1.n2 B 2.71937f
C156 VDD1.n3 B 4.49054f
C157 VDD1.t7 B 0.300632f
C158 VDD1.t3 B 0.300632f
C159 VDD1.n4 B 2.70064f
C160 VDD1.n5 B 3.84953f
C161 VP.t7 B 2.46521f
C162 VP.n0 B 0.922726f
C163 VP.n1 B 0.017417f
C164 VP.n2 B 0.033493f
C165 VP.n3 B 0.017417f
C166 VP.n4 B 0.031659f
C167 VP.n5 B 0.017417f
C168 VP.n6 B 0.034617f
C169 VP.n7 B 0.017417f
C170 VP.n8 B 0.032461f
C171 VP.n9 B 0.017417f
C172 VP.t6 B 2.46521f
C173 VP.n10 B 0.035172f
C174 VP.n11 B 0.017417f
C175 VP.n12 B 0.032461f
C176 VP.t5 B 2.46521f
C177 VP.n13 B 0.922726f
C178 VP.n14 B 0.017417f
C179 VP.n15 B 0.033493f
C180 VP.n16 B 0.017417f
C181 VP.n17 B 0.031659f
C182 VP.n18 B 0.017417f
C183 VP.n19 B 0.034617f
C184 VP.n20 B 0.017417f
C185 VP.n21 B 0.032461f
C186 VP.t1 B 2.72527f
C187 VP.n22 B 0.871805f
C188 VP.t2 B 2.46521f
C189 VP.n23 B 0.913384f
C190 VP.n24 B 0.017235f
C191 VP.n25 B 0.221642f
C192 VP.n26 B 0.017417f
C193 VP.n27 B 0.017417f
C194 VP.n28 B 0.032461f
C195 VP.n29 B 0.034617f
C196 VP.n30 B 0.01408f
C197 VP.n31 B 0.017417f
C198 VP.n32 B 0.017417f
C199 VP.n33 B 0.017417f
C200 VP.n34 B 0.032461f
C201 VP.n35 B 0.032461f
C202 VP.t3 B 2.46521f
C203 VP.n36 B 0.857937f
C204 VP.n37 B 0.017235f
C205 VP.n38 B 0.017417f
C206 VP.n39 B 0.017417f
C207 VP.n40 B 0.017417f
C208 VP.n41 B 0.032461f
C209 VP.n42 B 0.035172f
C210 VP.n43 B 0.014648f
C211 VP.n44 B 0.017417f
C212 VP.n45 B 0.017417f
C213 VP.n46 B 0.017417f
C214 VP.n47 B 0.032461f
C215 VP.n48 B 0.032461f
C216 VP.n49 B 0.018838f
C217 VP.n50 B 0.028111f
C218 VP.n51 B 1.21798f
C219 VP.n52 B 1.22884f
C220 VP.t4 B 2.46521f
C221 VP.n53 B 0.922726f
C222 VP.n54 B 0.018838f
C223 VP.n55 B 0.028111f
C224 VP.n56 B 0.017417f
C225 VP.n57 B 0.017417f
C226 VP.n58 B 0.032461f
C227 VP.n59 B 0.033493f
C228 VP.n60 B 0.014648f
C229 VP.n61 B 0.017417f
C230 VP.n62 B 0.017417f
C231 VP.n63 B 0.017417f
C232 VP.n64 B 0.032461f
C233 VP.n65 B 0.031659f
C234 VP.n66 B 0.857937f
C235 VP.n67 B 0.017235f
C236 VP.n68 B 0.017417f
C237 VP.n69 B 0.017417f
C238 VP.n70 B 0.017417f
C239 VP.n71 B 0.032461f
C240 VP.n72 B 0.034617f
C241 VP.n73 B 0.01408f
C242 VP.n74 B 0.017417f
C243 VP.n75 B 0.017417f
C244 VP.n76 B 0.017417f
C245 VP.n77 B 0.032461f
C246 VP.n78 B 0.032461f
C247 VP.t0 B 2.46521f
C248 VP.n79 B 0.857937f
C249 VP.n80 B 0.017235f
C250 VP.n81 B 0.017417f
C251 VP.n82 B 0.017417f
C252 VP.n83 B 0.017417f
C253 VP.n84 B 0.032461f
C254 VP.n85 B 0.035172f
C255 VP.n86 B 0.014648f
C256 VP.n87 B 0.017417f
C257 VP.n88 B 0.017417f
C258 VP.n89 B 0.017417f
C259 VP.n90 B 0.032461f
C260 VP.n91 B 0.032461f
C261 VP.n92 B 0.018838f
C262 VP.n93 B 0.028111f
C263 VP.n94 B 0.05233f
.ends

