* NGSPICE file created from diff_pair_sample_1551.ext - technology: sky130A

.subckt diff_pair_sample_1551 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X1 VDD1.t6 VP.t1 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X2 VTAIL.t13 VP.t2 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=1.9866 ps=12.37 w=12.04 l=1.34
X3 VTAIL.t7 VN.t0 VDD2.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=1.9866 ps=12.37 w=12.04 l=1.34
X4 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=0 ps=0 w=12.04 l=1.34
X5 VTAIL.t5 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=1.9866 ps=12.37 w=12.04 l=1.34
X6 VDD1.t1 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=4.6956 ps=24.86 w=12.04 l=1.34
X7 VDD1.t4 VP.t4 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X8 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=4.6956 ps=24.86 w=12.04 l=1.34
X9 VTAIL.t10 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X10 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X11 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=4.6956 ps=24.86 w=12.04 l=1.34
X12 VDD1.t5 VP.t6 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=4.6956 ps=24.86 w=12.04 l=1.34
X13 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X14 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=0 ps=0 w=12.04 l=1.34
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=0 ps=0 w=12.04 l=1.34
X16 VDD2.t1 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=0 ps=0 w=12.04 l=1.34
X18 VDD2.t0 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9866 pd=12.37 as=1.9866 ps=12.37 w=12.04 l=1.34
X19 VTAIL.t8 VP.t7 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6956 pd=24.86 as=1.9866 ps=12.37 w=12.04 l=1.34
R0 VP.n11 VP.t2 245.733
R1 VP.n5 VP.t7 216.541
R2 VP.n29 VP.t4 216.541
R3 VP.n36 VP.t5 216.541
R4 VP.n43 VP.t6 216.541
R5 VP.n23 VP.t3 216.541
R6 VP.n16 VP.t0 216.541
R7 VP.n10 VP.t1 216.541
R8 VP.n25 VP.n5 173.351
R9 VP.n44 VP.n43 173.351
R10 VP.n24 VP.n23 173.351
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n42 VP.n0 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n1 161.3
R21 VP.n38 VP.n37 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n11 VP.n10 61.2741
R29 VP.n35 VP.n34 56.5617
R30 VP.n15 VP.n14 56.5617
R31 VP.n30 VP.n28 48.3272
R32 VP.n41 VP.n1 48.3272
R33 VP.n21 VP.n7 48.3272
R34 VP.n25 VP.n24 44.955
R35 VP.n28 VP.n27 32.8269
R36 VP.n42 VP.n41 32.8269
R37 VP.n22 VP.n21 32.8269
R38 VP.n12 VP.n11 27.186
R39 VP.n34 VP.n3 24.5923
R40 VP.n37 VP.n35 24.5923
R41 VP.n17 VP.n15 24.5923
R42 VP.n14 VP.n9 24.5923
R43 VP.n30 VP.n29 20.4117
R44 VP.n36 VP.n1 20.4117
R45 VP.n16 VP.n7 20.4117
R46 VP.n27 VP.n5 12.5423
R47 VP.n43 VP.n42 12.5423
R48 VP.n23 VP.n22 12.5423
R49 VP.n29 VP.n3 4.18111
R50 VP.n37 VP.n36 4.18111
R51 VP.n17 VP.n16 4.18111
R52 VP.n10 VP.n9 4.18111
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VDD1 VDD1.n0 61.1065
R73 VDD1.n3 VDD1.n2 60.9927
R74 VDD1.n3 VDD1.n1 60.9927
R75 VDD1.n5 VDD1.n4 60.3283
R76 VDD1.n5 VDD1.n3 41.1561
R77 VDD1.n4 VDD1.t7 1.64502
R78 VDD1.n4 VDD1.t1 1.64502
R79 VDD1.n0 VDD1.t0 1.64502
R80 VDD1.n0 VDD1.t6 1.64502
R81 VDD1.n2 VDD1.t2 1.64502
R82 VDD1.n2 VDD1.t5 1.64502
R83 VDD1.n1 VDD1.t3 1.64502
R84 VDD1.n1 VDD1.t4 1.64502
R85 VDD1 VDD1.n5 0.662138
R86 VTAIL.n530 VTAIL.n470 289.615
R87 VTAIL.n62 VTAIL.n2 289.615
R88 VTAIL.n128 VTAIL.n68 289.615
R89 VTAIL.n196 VTAIL.n136 289.615
R90 VTAIL.n464 VTAIL.n404 289.615
R91 VTAIL.n396 VTAIL.n336 289.615
R92 VTAIL.n330 VTAIL.n270 289.615
R93 VTAIL.n262 VTAIL.n202 289.615
R94 VTAIL.n490 VTAIL.n489 185
R95 VTAIL.n495 VTAIL.n494 185
R96 VTAIL.n497 VTAIL.n496 185
R97 VTAIL.n486 VTAIL.n485 185
R98 VTAIL.n503 VTAIL.n502 185
R99 VTAIL.n505 VTAIL.n504 185
R100 VTAIL.n482 VTAIL.n481 185
R101 VTAIL.n512 VTAIL.n511 185
R102 VTAIL.n513 VTAIL.n480 185
R103 VTAIL.n515 VTAIL.n514 185
R104 VTAIL.n478 VTAIL.n477 185
R105 VTAIL.n521 VTAIL.n520 185
R106 VTAIL.n523 VTAIL.n522 185
R107 VTAIL.n474 VTAIL.n473 185
R108 VTAIL.n529 VTAIL.n528 185
R109 VTAIL.n531 VTAIL.n530 185
R110 VTAIL.n22 VTAIL.n21 185
R111 VTAIL.n27 VTAIL.n26 185
R112 VTAIL.n29 VTAIL.n28 185
R113 VTAIL.n18 VTAIL.n17 185
R114 VTAIL.n35 VTAIL.n34 185
R115 VTAIL.n37 VTAIL.n36 185
R116 VTAIL.n14 VTAIL.n13 185
R117 VTAIL.n44 VTAIL.n43 185
R118 VTAIL.n45 VTAIL.n12 185
R119 VTAIL.n47 VTAIL.n46 185
R120 VTAIL.n10 VTAIL.n9 185
R121 VTAIL.n53 VTAIL.n52 185
R122 VTAIL.n55 VTAIL.n54 185
R123 VTAIL.n6 VTAIL.n5 185
R124 VTAIL.n61 VTAIL.n60 185
R125 VTAIL.n63 VTAIL.n62 185
R126 VTAIL.n88 VTAIL.n87 185
R127 VTAIL.n93 VTAIL.n92 185
R128 VTAIL.n95 VTAIL.n94 185
R129 VTAIL.n84 VTAIL.n83 185
R130 VTAIL.n101 VTAIL.n100 185
R131 VTAIL.n103 VTAIL.n102 185
R132 VTAIL.n80 VTAIL.n79 185
R133 VTAIL.n110 VTAIL.n109 185
R134 VTAIL.n111 VTAIL.n78 185
R135 VTAIL.n113 VTAIL.n112 185
R136 VTAIL.n76 VTAIL.n75 185
R137 VTAIL.n119 VTAIL.n118 185
R138 VTAIL.n121 VTAIL.n120 185
R139 VTAIL.n72 VTAIL.n71 185
R140 VTAIL.n127 VTAIL.n126 185
R141 VTAIL.n129 VTAIL.n128 185
R142 VTAIL.n156 VTAIL.n155 185
R143 VTAIL.n161 VTAIL.n160 185
R144 VTAIL.n163 VTAIL.n162 185
R145 VTAIL.n152 VTAIL.n151 185
R146 VTAIL.n169 VTAIL.n168 185
R147 VTAIL.n171 VTAIL.n170 185
R148 VTAIL.n148 VTAIL.n147 185
R149 VTAIL.n178 VTAIL.n177 185
R150 VTAIL.n179 VTAIL.n146 185
R151 VTAIL.n181 VTAIL.n180 185
R152 VTAIL.n144 VTAIL.n143 185
R153 VTAIL.n187 VTAIL.n186 185
R154 VTAIL.n189 VTAIL.n188 185
R155 VTAIL.n140 VTAIL.n139 185
R156 VTAIL.n195 VTAIL.n194 185
R157 VTAIL.n197 VTAIL.n196 185
R158 VTAIL.n465 VTAIL.n464 185
R159 VTAIL.n463 VTAIL.n462 185
R160 VTAIL.n408 VTAIL.n407 185
R161 VTAIL.n457 VTAIL.n456 185
R162 VTAIL.n455 VTAIL.n454 185
R163 VTAIL.n412 VTAIL.n411 185
R164 VTAIL.n449 VTAIL.n448 185
R165 VTAIL.n447 VTAIL.n414 185
R166 VTAIL.n446 VTAIL.n445 185
R167 VTAIL.n417 VTAIL.n415 185
R168 VTAIL.n440 VTAIL.n439 185
R169 VTAIL.n438 VTAIL.n437 185
R170 VTAIL.n421 VTAIL.n420 185
R171 VTAIL.n432 VTAIL.n431 185
R172 VTAIL.n430 VTAIL.n429 185
R173 VTAIL.n425 VTAIL.n424 185
R174 VTAIL.n397 VTAIL.n396 185
R175 VTAIL.n395 VTAIL.n394 185
R176 VTAIL.n340 VTAIL.n339 185
R177 VTAIL.n389 VTAIL.n388 185
R178 VTAIL.n387 VTAIL.n386 185
R179 VTAIL.n344 VTAIL.n343 185
R180 VTAIL.n381 VTAIL.n380 185
R181 VTAIL.n379 VTAIL.n346 185
R182 VTAIL.n378 VTAIL.n377 185
R183 VTAIL.n349 VTAIL.n347 185
R184 VTAIL.n372 VTAIL.n371 185
R185 VTAIL.n370 VTAIL.n369 185
R186 VTAIL.n353 VTAIL.n352 185
R187 VTAIL.n364 VTAIL.n363 185
R188 VTAIL.n362 VTAIL.n361 185
R189 VTAIL.n357 VTAIL.n356 185
R190 VTAIL.n331 VTAIL.n330 185
R191 VTAIL.n329 VTAIL.n328 185
R192 VTAIL.n274 VTAIL.n273 185
R193 VTAIL.n323 VTAIL.n322 185
R194 VTAIL.n321 VTAIL.n320 185
R195 VTAIL.n278 VTAIL.n277 185
R196 VTAIL.n315 VTAIL.n314 185
R197 VTAIL.n313 VTAIL.n280 185
R198 VTAIL.n312 VTAIL.n311 185
R199 VTAIL.n283 VTAIL.n281 185
R200 VTAIL.n306 VTAIL.n305 185
R201 VTAIL.n304 VTAIL.n303 185
R202 VTAIL.n287 VTAIL.n286 185
R203 VTAIL.n298 VTAIL.n297 185
R204 VTAIL.n296 VTAIL.n295 185
R205 VTAIL.n291 VTAIL.n290 185
R206 VTAIL.n263 VTAIL.n262 185
R207 VTAIL.n261 VTAIL.n260 185
R208 VTAIL.n206 VTAIL.n205 185
R209 VTAIL.n255 VTAIL.n254 185
R210 VTAIL.n253 VTAIL.n252 185
R211 VTAIL.n210 VTAIL.n209 185
R212 VTAIL.n247 VTAIL.n246 185
R213 VTAIL.n245 VTAIL.n212 185
R214 VTAIL.n244 VTAIL.n243 185
R215 VTAIL.n215 VTAIL.n213 185
R216 VTAIL.n238 VTAIL.n237 185
R217 VTAIL.n236 VTAIL.n235 185
R218 VTAIL.n219 VTAIL.n218 185
R219 VTAIL.n230 VTAIL.n229 185
R220 VTAIL.n228 VTAIL.n227 185
R221 VTAIL.n223 VTAIL.n222 185
R222 VTAIL.n491 VTAIL.t2 149.524
R223 VTAIL.n23 VTAIL.t5 149.524
R224 VTAIL.n89 VTAIL.t9 149.524
R225 VTAIL.n157 VTAIL.t8 149.524
R226 VTAIL.n426 VTAIL.t12 149.524
R227 VTAIL.n358 VTAIL.t13 149.524
R228 VTAIL.n292 VTAIL.t3 149.524
R229 VTAIL.n224 VTAIL.t7 149.524
R230 VTAIL.n495 VTAIL.n489 104.615
R231 VTAIL.n496 VTAIL.n495 104.615
R232 VTAIL.n496 VTAIL.n485 104.615
R233 VTAIL.n503 VTAIL.n485 104.615
R234 VTAIL.n504 VTAIL.n503 104.615
R235 VTAIL.n504 VTAIL.n481 104.615
R236 VTAIL.n512 VTAIL.n481 104.615
R237 VTAIL.n513 VTAIL.n512 104.615
R238 VTAIL.n514 VTAIL.n513 104.615
R239 VTAIL.n514 VTAIL.n477 104.615
R240 VTAIL.n521 VTAIL.n477 104.615
R241 VTAIL.n522 VTAIL.n521 104.615
R242 VTAIL.n522 VTAIL.n473 104.615
R243 VTAIL.n529 VTAIL.n473 104.615
R244 VTAIL.n530 VTAIL.n529 104.615
R245 VTAIL.n27 VTAIL.n21 104.615
R246 VTAIL.n28 VTAIL.n27 104.615
R247 VTAIL.n28 VTAIL.n17 104.615
R248 VTAIL.n35 VTAIL.n17 104.615
R249 VTAIL.n36 VTAIL.n35 104.615
R250 VTAIL.n36 VTAIL.n13 104.615
R251 VTAIL.n44 VTAIL.n13 104.615
R252 VTAIL.n45 VTAIL.n44 104.615
R253 VTAIL.n46 VTAIL.n45 104.615
R254 VTAIL.n46 VTAIL.n9 104.615
R255 VTAIL.n53 VTAIL.n9 104.615
R256 VTAIL.n54 VTAIL.n53 104.615
R257 VTAIL.n54 VTAIL.n5 104.615
R258 VTAIL.n61 VTAIL.n5 104.615
R259 VTAIL.n62 VTAIL.n61 104.615
R260 VTAIL.n93 VTAIL.n87 104.615
R261 VTAIL.n94 VTAIL.n93 104.615
R262 VTAIL.n94 VTAIL.n83 104.615
R263 VTAIL.n101 VTAIL.n83 104.615
R264 VTAIL.n102 VTAIL.n101 104.615
R265 VTAIL.n102 VTAIL.n79 104.615
R266 VTAIL.n110 VTAIL.n79 104.615
R267 VTAIL.n111 VTAIL.n110 104.615
R268 VTAIL.n112 VTAIL.n111 104.615
R269 VTAIL.n112 VTAIL.n75 104.615
R270 VTAIL.n119 VTAIL.n75 104.615
R271 VTAIL.n120 VTAIL.n119 104.615
R272 VTAIL.n120 VTAIL.n71 104.615
R273 VTAIL.n127 VTAIL.n71 104.615
R274 VTAIL.n128 VTAIL.n127 104.615
R275 VTAIL.n161 VTAIL.n155 104.615
R276 VTAIL.n162 VTAIL.n161 104.615
R277 VTAIL.n162 VTAIL.n151 104.615
R278 VTAIL.n169 VTAIL.n151 104.615
R279 VTAIL.n170 VTAIL.n169 104.615
R280 VTAIL.n170 VTAIL.n147 104.615
R281 VTAIL.n178 VTAIL.n147 104.615
R282 VTAIL.n179 VTAIL.n178 104.615
R283 VTAIL.n180 VTAIL.n179 104.615
R284 VTAIL.n180 VTAIL.n143 104.615
R285 VTAIL.n187 VTAIL.n143 104.615
R286 VTAIL.n188 VTAIL.n187 104.615
R287 VTAIL.n188 VTAIL.n139 104.615
R288 VTAIL.n195 VTAIL.n139 104.615
R289 VTAIL.n196 VTAIL.n195 104.615
R290 VTAIL.n464 VTAIL.n463 104.615
R291 VTAIL.n463 VTAIL.n407 104.615
R292 VTAIL.n456 VTAIL.n407 104.615
R293 VTAIL.n456 VTAIL.n455 104.615
R294 VTAIL.n455 VTAIL.n411 104.615
R295 VTAIL.n448 VTAIL.n411 104.615
R296 VTAIL.n448 VTAIL.n447 104.615
R297 VTAIL.n447 VTAIL.n446 104.615
R298 VTAIL.n446 VTAIL.n415 104.615
R299 VTAIL.n439 VTAIL.n415 104.615
R300 VTAIL.n439 VTAIL.n438 104.615
R301 VTAIL.n438 VTAIL.n420 104.615
R302 VTAIL.n431 VTAIL.n420 104.615
R303 VTAIL.n431 VTAIL.n430 104.615
R304 VTAIL.n430 VTAIL.n424 104.615
R305 VTAIL.n396 VTAIL.n395 104.615
R306 VTAIL.n395 VTAIL.n339 104.615
R307 VTAIL.n388 VTAIL.n339 104.615
R308 VTAIL.n388 VTAIL.n387 104.615
R309 VTAIL.n387 VTAIL.n343 104.615
R310 VTAIL.n380 VTAIL.n343 104.615
R311 VTAIL.n380 VTAIL.n379 104.615
R312 VTAIL.n379 VTAIL.n378 104.615
R313 VTAIL.n378 VTAIL.n347 104.615
R314 VTAIL.n371 VTAIL.n347 104.615
R315 VTAIL.n371 VTAIL.n370 104.615
R316 VTAIL.n370 VTAIL.n352 104.615
R317 VTAIL.n363 VTAIL.n352 104.615
R318 VTAIL.n363 VTAIL.n362 104.615
R319 VTAIL.n362 VTAIL.n356 104.615
R320 VTAIL.n330 VTAIL.n329 104.615
R321 VTAIL.n329 VTAIL.n273 104.615
R322 VTAIL.n322 VTAIL.n273 104.615
R323 VTAIL.n322 VTAIL.n321 104.615
R324 VTAIL.n321 VTAIL.n277 104.615
R325 VTAIL.n314 VTAIL.n277 104.615
R326 VTAIL.n314 VTAIL.n313 104.615
R327 VTAIL.n313 VTAIL.n312 104.615
R328 VTAIL.n312 VTAIL.n281 104.615
R329 VTAIL.n305 VTAIL.n281 104.615
R330 VTAIL.n305 VTAIL.n304 104.615
R331 VTAIL.n304 VTAIL.n286 104.615
R332 VTAIL.n297 VTAIL.n286 104.615
R333 VTAIL.n297 VTAIL.n296 104.615
R334 VTAIL.n296 VTAIL.n290 104.615
R335 VTAIL.n262 VTAIL.n261 104.615
R336 VTAIL.n261 VTAIL.n205 104.615
R337 VTAIL.n254 VTAIL.n205 104.615
R338 VTAIL.n254 VTAIL.n253 104.615
R339 VTAIL.n253 VTAIL.n209 104.615
R340 VTAIL.n246 VTAIL.n209 104.615
R341 VTAIL.n246 VTAIL.n245 104.615
R342 VTAIL.n245 VTAIL.n244 104.615
R343 VTAIL.n244 VTAIL.n213 104.615
R344 VTAIL.n237 VTAIL.n213 104.615
R345 VTAIL.n237 VTAIL.n236 104.615
R346 VTAIL.n236 VTAIL.n218 104.615
R347 VTAIL.n229 VTAIL.n218 104.615
R348 VTAIL.n229 VTAIL.n228 104.615
R349 VTAIL.n228 VTAIL.n222 104.615
R350 VTAIL.t2 VTAIL.n489 52.3082
R351 VTAIL.t5 VTAIL.n21 52.3082
R352 VTAIL.t9 VTAIL.n87 52.3082
R353 VTAIL.t8 VTAIL.n155 52.3082
R354 VTAIL.t12 VTAIL.n424 52.3082
R355 VTAIL.t13 VTAIL.n356 52.3082
R356 VTAIL.t3 VTAIL.n290 52.3082
R357 VTAIL.t7 VTAIL.n222 52.3082
R358 VTAIL.n403 VTAIL.n402 43.6496
R359 VTAIL.n269 VTAIL.n268 43.6496
R360 VTAIL.n1 VTAIL.n0 43.6495
R361 VTAIL.n135 VTAIL.n134 43.6495
R362 VTAIL.n535 VTAIL.n534 30.6338
R363 VTAIL.n67 VTAIL.n66 30.6338
R364 VTAIL.n133 VTAIL.n132 30.6338
R365 VTAIL.n201 VTAIL.n200 30.6338
R366 VTAIL.n469 VTAIL.n468 30.6338
R367 VTAIL.n401 VTAIL.n400 30.6338
R368 VTAIL.n335 VTAIL.n334 30.6338
R369 VTAIL.n267 VTAIL.n266 30.6338
R370 VTAIL.n535 VTAIL.n469 24.1858
R371 VTAIL.n267 VTAIL.n201 24.1858
R372 VTAIL.n515 VTAIL.n480 13.1884
R373 VTAIL.n47 VTAIL.n12 13.1884
R374 VTAIL.n113 VTAIL.n78 13.1884
R375 VTAIL.n181 VTAIL.n146 13.1884
R376 VTAIL.n449 VTAIL.n414 13.1884
R377 VTAIL.n381 VTAIL.n346 13.1884
R378 VTAIL.n315 VTAIL.n280 13.1884
R379 VTAIL.n247 VTAIL.n212 13.1884
R380 VTAIL.n511 VTAIL.n510 12.8005
R381 VTAIL.n516 VTAIL.n478 12.8005
R382 VTAIL.n43 VTAIL.n42 12.8005
R383 VTAIL.n48 VTAIL.n10 12.8005
R384 VTAIL.n109 VTAIL.n108 12.8005
R385 VTAIL.n114 VTAIL.n76 12.8005
R386 VTAIL.n177 VTAIL.n176 12.8005
R387 VTAIL.n182 VTAIL.n144 12.8005
R388 VTAIL.n450 VTAIL.n412 12.8005
R389 VTAIL.n445 VTAIL.n416 12.8005
R390 VTAIL.n382 VTAIL.n344 12.8005
R391 VTAIL.n377 VTAIL.n348 12.8005
R392 VTAIL.n316 VTAIL.n278 12.8005
R393 VTAIL.n311 VTAIL.n282 12.8005
R394 VTAIL.n248 VTAIL.n210 12.8005
R395 VTAIL.n243 VTAIL.n214 12.8005
R396 VTAIL.n509 VTAIL.n482 12.0247
R397 VTAIL.n520 VTAIL.n519 12.0247
R398 VTAIL.n41 VTAIL.n14 12.0247
R399 VTAIL.n52 VTAIL.n51 12.0247
R400 VTAIL.n107 VTAIL.n80 12.0247
R401 VTAIL.n118 VTAIL.n117 12.0247
R402 VTAIL.n175 VTAIL.n148 12.0247
R403 VTAIL.n186 VTAIL.n185 12.0247
R404 VTAIL.n454 VTAIL.n453 12.0247
R405 VTAIL.n444 VTAIL.n417 12.0247
R406 VTAIL.n386 VTAIL.n385 12.0247
R407 VTAIL.n376 VTAIL.n349 12.0247
R408 VTAIL.n320 VTAIL.n319 12.0247
R409 VTAIL.n310 VTAIL.n283 12.0247
R410 VTAIL.n252 VTAIL.n251 12.0247
R411 VTAIL.n242 VTAIL.n215 12.0247
R412 VTAIL.n506 VTAIL.n505 11.249
R413 VTAIL.n523 VTAIL.n476 11.249
R414 VTAIL.n38 VTAIL.n37 11.249
R415 VTAIL.n55 VTAIL.n8 11.249
R416 VTAIL.n104 VTAIL.n103 11.249
R417 VTAIL.n121 VTAIL.n74 11.249
R418 VTAIL.n172 VTAIL.n171 11.249
R419 VTAIL.n189 VTAIL.n142 11.249
R420 VTAIL.n457 VTAIL.n410 11.249
R421 VTAIL.n441 VTAIL.n440 11.249
R422 VTAIL.n389 VTAIL.n342 11.249
R423 VTAIL.n373 VTAIL.n372 11.249
R424 VTAIL.n323 VTAIL.n276 11.249
R425 VTAIL.n307 VTAIL.n306 11.249
R426 VTAIL.n255 VTAIL.n208 11.249
R427 VTAIL.n239 VTAIL.n238 11.249
R428 VTAIL.n502 VTAIL.n484 10.4732
R429 VTAIL.n524 VTAIL.n474 10.4732
R430 VTAIL.n34 VTAIL.n16 10.4732
R431 VTAIL.n56 VTAIL.n6 10.4732
R432 VTAIL.n100 VTAIL.n82 10.4732
R433 VTAIL.n122 VTAIL.n72 10.4732
R434 VTAIL.n168 VTAIL.n150 10.4732
R435 VTAIL.n190 VTAIL.n140 10.4732
R436 VTAIL.n458 VTAIL.n408 10.4732
R437 VTAIL.n437 VTAIL.n419 10.4732
R438 VTAIL.n390 VTAIL.n340 10.4732
R439 VTAIL.n369 VTAIL.n351 10.4732
R440 VTAIL.n324 VTAIL.n274 10.4732
R441 VTAIL.n303 VTAIL.n285 10.4732
R442 VTAIL.n256 VTAIL.n206 10.4732
R443 VTAIL.n235 VTAIL.n217 10.4732
R444 VTAIL.n491 VTAIL.n490 10.2747
R445 VTAIL.n23 VTAIL.n22 10.2747
R446 VTAIL.n89 VTAIL.n88 10.2747
R447 VTAIL.n157 VTAIL.n156 10.2747
R448 VTAIL.n426 VTAIL.n425 10.2747
R449 VTAIL.n358 VTAIL.n357 10.2747
R450 VTAIL.n292 VTAIL.n291 10.2747
R451 VTAIL.n224 VTAIL.n223 10.2747
R452 VTAIL.n501 VTAIL.n486 9.69747
R453 VTAIL.n528 VTAIL.n527 9.69747
R454 VTAIL.n33 VTAIL.n18 9.69747
R455 VTAIL.n60 VTAIL.n59 9.69747
R456 VTAIL.n99 VTAIL.n84 9.69747
R457 VTAIL.n126 VTAIL.n125 9.69747
R458 VTAIL.n167 VTAIL.n152 9.69747
R459 VTAIL.n194 VTAIL.n193 9.69747
R460 VTAIL.n462 VTAIL.n461 9.69747
R461 VTAIL.n436 VTAIL.n421 9.69747
R462 VTAIL.n394 VTAIL.n393 9.69747
R463 VTAIL.n368 VTAIL.n353 9.69747
R464 VTAIL.n328 VTAIL.n327 9.69747
R465 VTAIL.n302 VTAIL.n287 9.69747
R466 VTAIL.n260 VTAIL.n259 9.69747
R467 VTAIL.n234 VTAIL.n219 9.69747
R468 VTAIL.n534 VTAIL.n533 9.45567
R469 VTAIL.n66 VTAIL.n65 9.45567
R470 VTAIL.n132 VTAIL.n131 9.45567
R471 VTAIL.n200 VTAIL.n199 9.45567
R472 VTAIL.n468 VTAIL.n467 9.45567
R473 VTAIL.n400 VTAIL.n399 9.45567
R474 VTAIL.n334 VTAIL.n333 9.45567
R475 VTAIL.n266 VTAIL.n265 9.45567
R476 VTAIL.n533 VTAIL.n532 9.3005
R477 VTAIL.n472 VTAIL.n471 9.3005
R478 VTAIL.n527 VTAIL.n526 9.3005
R479 VTAIL.n525 VTAIL.n524 9.3005
R480 VTAIL.n476 VTAIL.n475 9.3005
R481 VTAIL.n519 VTAIL.n518 9.3005
R482 VTAIL.n517 VTAIL.n516 9.3005
R483 VTAIL.n493 VTAIL.n492 9.3005
R484 VTAIL.n488 VTAIL.n487 9.3005
R485 VTAIL.n499 VTAIL.n498 9.3005
R486 VTAIL.n501 VTAIL.n500 9.3005
R487 VTAIL.n484 VTAIL.n483 9.3005
R488 VTAIL.n507 VTAIL.n506 9.3005
R489 VTAIL.n509 VTAIL.n508 9.3005
R490 VTAIL.n510 VTAIL.n479 9.3005
R491 VTAIL.n65 VTAIL.n64 9.3005
R492 VTAIL.n4 VTAIL.n3 9.3005
R493 VTAIL.n59 VTAIL.n58 9.3005
R494 VTAIL.n57 VTAIL.n56 9.3005
R495 VTAIL.n8 VTAIL.n7 9.3005
R496 VTAIL.n51 VTAIL.n50 9.3005
R497 VTAIL.n49 VTAIL.n48 9.3005
R498 VTAIL.n25 VTAIL.n24 9.3005
R499 VTAIL.n20 VTAIL.n19 9.3005
R500 VTAIL.n31 VTAIL.n30 9.3005
R501 VTAIL.n33 VTAIL.n32 9.3005
R502 VTAIL.n16 VTAIL.n15 9.3005
R503 VTAIL.n39 VTAIL.n38 9.3005
R504 VTAIL.n41 VTAIL.n40 9.3005
R505 VTAIL.n42 VTAIL.n11 9.3005
R506 VTAIL.n131 VTAIL.n130 9.3005
R507 VTAIL.n70 VTAIL.n69 9.3005
R508 VTAIL.n125 VTAIL.n124 9.3005
R509 VTAIL.n123 VTAIL.n122 9.3005
R510 VTAIL.n74 VTAIL.n73 9.3005
R511 VTAIL.n117 VTAIL.n116 9.3005
R512 VTAIL.n115 VTAIL.n114 9.3005
R513 VTAIL.n91 VTAIL.n90 9.3005
R514 VTAIL.n86 VTAIL.n85 9.3005
R515 VTAIL.n97 VTAIL.n96 9.3005
R516 VTAIL.n99 VTAIL.n98 9.3005
R517 VTAIL.n82 VTAIL.n81 9.3005
R518 VTAIL.n105 VTAIL.n104 9.3005
R519 VTAIL.n107 VTAIL.n106 9.3005
R520 VTAIL.n108 VTAIL.n77 9.3005
R521 VTAIL.n199 VTAIL.n198 9.3005
R522 VTAIL.n138 VTAIL.n137 9.3005
R523 VTAIL.n193 VTAIL.n192 9.3005
R524 VTAIL.n191 VTAIL.n190 9.3005
R525 VTAIL.n142 VTAIL.n141 9.3005
R526 VTAIL.n185 VTAIL.n184 9.3005
R527 VTAIL.n183 VTAIL.n182 9.3005
R528 VTAIL.n159 VTAIL.n158 9.3005
R529 VTAIL.n154 VTAIL.n153 9.3005
R530 VTAIL.n165 VTAIL.n164 9.3005
R531 VTAIL.n167 VTAIL.n166 9.3005
R532 VTAIL.n150 VTAIL.n149 9.3005
R533 VTAIL.n173 VTAIL.n172 9.3005
R534 VTAIL.n175 VTAIL.n174 9.3005
R535 VTAIL.n176 VTAIL.n145 9.3005
R536 VTAIL.n428 VTAIL.n427 9.3005
R537 VTAIL.n423 VTAIL.n422 9.3005
R538 VTAIL.n434 VTAIL.n433 9.3005
R539 VTAIL.n436 VTAIL.n435 9.3005
R540 VTAIL.n419 VTAIL.n418 9.3005
R541 VTAIL.n442 VTAIL.n441 9.3005
R542 VTAIL.n444 VTAIL.n443 9.3005
R543 VTAIL.n416 VTAIL.n413 9.3005
R544 VTAIL.n467 VTAIL.n466 9.3005
R545 VTAIL.n406 VTAIL.n405 9.3005
R546 VTAIL.n461 VTAIL.n460 9.3005
R547 VTAIL.n459 VTAIL.n458 9.3005
R548 VTAIL.n410 VTAIL.n409 9.3005
R549 VTAIL.n453 VTAIL.n452 9.3005
R550 VTAIL.n451 VTAIL.n450 9.3005
R551 VTAIL.n360 VTAIL.n359 9.3005
R552 VTAIL.n355 VTAIL.n354 9.3005
R553 VTAIL.n366 VTAIL.n365 9.3005
R554 VTAIL.n368 VTAIL.n367 9.3005
R555 VTAIL.n351 VTAIL.n350 9.3005
R556 VTAIL.n374 VTAIL.n373 9.3005
R557 VTAIL.n376 VTAIL.n375 9.3005
R558 VTAIL.n348 VTAIL.n345 9.3005
R559 VTAIL.n399 VTAIL.n398 9.3005
R560 VTAIL.n338 VTAIL.n337 9.3005
R561 VTAIL.n393 VTAIL.n392 9.3005
R562 VTAIL.n391 VTAIL.n390 9.3005
R563 VTAIL.n342 VTAIL.n341 9.3005
R564 VTAIL.n385 VTAIL.n384 9.3005
R565 VTAIL.n383 VTAIL.n382 9.3005
R566 VTAIL.n294 VTAIL.n293 9.3005
R567 VTAIL.n289 VTAIL.n288 9.3005
R568 VTAIL.n300 VTAIL.n299 9.3005
R569 VTAIL.n302 VTAIL.n301 9.3005
R570 VTAIL.n285 VTAIL.n284 9.3005
R571 VTAIL.n308 VTAIL.n307 9.3005
R572 VTAIL.n310 VTAIL.n309 9.3005
R573 VTAIL.n282 VTAIL.n279 9.3005
R574 VTAIL.n333 VTAIL.n332 9.3005
R575 VTAIL.n272 VTAIL.n271 9.3005
R576 VTAIL.n327 VTAIL.n326 9.3005
R577 VTAIL.n325 VTAIL.n324 9.3005
R578 VTAIL.n276 VTAIL.n275 9.3005
R579 VTAIL.n319 VTAIL.n318 9.3005
R580 VTAIL.n317 VTAIL.n316 9.3005
R581 VTAIL.n226 VTAIL.n225 9.3005
R582 VTAIL.n221 VTAIL.n220 9.3005
R583 VTAIL.n232 VTAIL.n231 9.3005
R584 VTAIL.n234 VTAIL.n233 9.3005
R585 VTAIL.n217 VTAIL.n216 9.3005
R586 VTAIL.n240 VTAIL.n239 9.3005
R587 VTAIL.n242 VTAIL.n241 9.3005
R588 VTAIL.n214 VTAIL.n211 9.3005
R589 VTAIL.n265 VTAIL.n264 9.3005
R590 VTAIL.n204 VTAIL.n203 9.3005
R591 VTAIL.n259 VTAIL.n258 9.3005
R592 VTAIL.n257 VTAIL.n256 9.3005
R593 VTAIL.n208 VTAIL.n207 9.3005
R594 VTAIL.n251 VTAIL.n250 9.3005
R595 VTAIL.n249 VTAIL.n248 9.3005
R596 VTAIL.n498 VTAIL.n497 8.92171
R597 VTAIL.n531 VTAIL.n472 8.92171
R598 VTAIL.n30 VTAIL.n29 8.92171
R599 VTAIL.n63 VTAIL.n4 8.92171
R600 VTAIL.n96 VTAIL.n95 8.92171
R601 VTAIL.n129 VTAIL.n70 8.92171
R602 VTAIL.n164 VTAIL.n163 8.92171
R603 VTAIL.n197 VTAIL.n138 8.92171
R604 VTAIL.n465 VTAIL.n406 8.92171
R605 VTAIL.n433 VTAIL.n432 8.92171
R606 VTAIL.n397 VTAIL.n338 8.92171
R607 VTAIL.n365 VTAIL.n364 8.92171
R608 VTAIL.n331 VTAIL.n272 8.92171
R609 VTAIL.n299 VTAIL.n298 8.92171
R610 VTAIL.n263 VTAIL.n204 8.92171
R611 VTAIL.n231 VTAIL.n230 8.92171
R612 VTAIL.n494 VTAIL.n488 8.14595
R613 VTAIL.n532 VTAIL.n470 8.14595
R614 VTAIL.n26 VTAIL.n20 8.14595
R615 VTAIL.n64 VTAIL.n2 8.14595
R616 VTAIL.n92 VTAIL.n86 8.14595
R617 VTAIL.n130 VTAIL.n68 8.14595
R618 VTAIL.n160 VTAIL.n154 8.14595
R619 VTAIL.n198 VTAIL.n136 8.14595
R620 VTAIL.n466 VTAIL.n404 8.14595
R621 VTAIL.n429 VTAIL.n423 8.14595
R622 VTAIL.n398 VTAIL.n336 8.14595
R623 VTAIL.n361 VTAIL.n355 8.14595
R624 VTAIL.n332 VTAIL.n270 8.14595
R625 VTAIL.n295 VTAIL.n289 8.14595
R626 VTAIL.n264 VTAIL.n202 8.14595
R627 VTAIL.n227 VTAIL.n221 8.14595
R628 VTAIL.n493 VTAIL.n490 7.3702
R629 VTAIL.n25 VTAIL.n22 7.3702
R630 VTAIL.n91 VTAIL.n88 7.3702
R631 VTAIL.n159 VTAIL.n156 7.3702
R632 VTAIL.n428 VTAIL.n425 7.3702
R633 VTAIL.n360 VTAIL.n357 7.3702
R634 VTAIL.n294 VTAIL.n291 7.3702
R635 VTAIL.n226 VTAIL.n223 7.3702
R636 VTAIL.n494 VTAIL.n493 5.81868
R637 VTAIL.n534 VTAIL.n470 5.81868
R638 VTAIL.n26 VTAIL.n25 5.81868
R639 VTAIL.n66 VTAIL.n2 5.81868
R640 VTAIL.n92 VTAIL.n91 5.81868
R641 VTAIL.n132 VTAIL.n68 5.81868
R642 VTAIL.n160 VTAIL.n159 5.81868
R643 VTAIL.n200 VTAIL.n136 5.81868
R644 VTAIL.n468 VTAIL.n404 5.81868
R645 VTAIL.n429 VTAIL.n428 5.81868
R646 VTAIL.n400 VTAIL.n336 5.81868
R647 VTAIL.n361 VTAIL.n360 5.81868
R648 VTAIL.n334 VTAIL.n270 5.81868
R649 VTAIL.n295 VTAIL.n294 5.81868
R650 VTAIL.n266 VTAIL.n202 5.81868
R651 VTAIL.n227 VTAIL.n226 5.81868
R652 VTAIL.n497 VTAIL.n488 5.04292
R653 VTAIL.n532 VTAIL.n531 5.04292
R654 VTAIL.n29 VTAIL.n20 5.04292
R655 VTAIL.n64 VTAIL.n63 5.04292
R656 VTAIL.n95 VTAIL.n86 5.04292
R657 VTAIL.n130 VTAIL.n129 5.04292
R658 VTAIL.n163 VTAIL.n154 5.04292
R659 VTAIL.n198 VTAIL.n197 5.04292
R660 VTAIL.n466 VTAIL.n465 5.04292
R661 VTAIL.n432 VTAIL.n423 5.04292
R662 VTAIL.n398 VTAIL.n397 5.04292
R663 VTAIL.n364 VTAIL.n355 5.04292
R664 VTAIL.n332 VTAIL.n331 5.04292
R665 VTAIL.n298 VTAIL.n289 5.04292
R666 VTAIL.n264 VTAIL.n263 5.04292
R667 VTAIL.n230 VTAIL.n221 5.04292
R668 VTAIL.n498 VTAIL.n486 4.26717
R669 VTAIL.n528 VTAIL.n472 4.26717
R670 VTAIL.n30 VTAIL.n18 4.26717
R671 VTAIL.n60 VTAIL.n4 4.26717
R672 VTAIL.n96 VTAIL.n84 4.26717
R673 VTAIL.n126 VTAIL.n70 4.26717
R674 VTAIL.n164 VTAIL.n152 4.26717
R675 VTAIL.n194 VTAIL.n138 4.26717
R676 VTAIL.n462 VTAIL.n406 4.26717
R677 VTAIL.n433 VTAIL.n421 4.26717
R678 VTAIL.n394 VTAIL.n338 4.26717
R679 VTAIL.n365 VTAIL.n353 4.26717
R680 VTAIL.n328 VTAIL.n272 4.26717
R681 VTAIL.n299 VTAIL.n287 4.26717
R682 VTAIL.n260 VTAIL.n204 4.26717
R683 VTAIL.n231 VTAIL.n219 4.26717
R684 VTAIL.n502 VTAIL.n501 3.49141
R685 VTAIL.n527 VTAIL.n474 3.49141
R686 VTAIL.n34 VTAIL.n33 3.49141
R687 VTAIL.n59 VTAIL.n6 3.49141
R688 VTAIL.n100 VTAIL.n99 3.49141
R689 VTAIL.n125 VTAIL.n72 3.49141
R690 VTAIL.n168 VTAIL.n167 3.49141
R691 VTAIL.n193 VTAIL.n140 3.49141
R692 VTAIL.n461 VTAIL.n408 3.49141
R693 VTAIL.n437 VTAIL.n436 3.49141
R694 VTAIL.n393 VTAIL.n340 3.49141
R695 VTAIL.n369 VTAIL.n368 3.49141
R696 VTAIL.n327 VTAIL.n274 3.49141
R697 VTAIL.n303 VTAIL.n302 3.49141
R698 VTAIL.n259 VTAIL.n206 3.49141
R699 VTAIL.n235 VTAIL.n234 3.49141
R700 VTAIL.n492 VTAIL.n491 2.84303
R701 VTAIL.n24 VTAIL.n23 2.84303
R702 VTAIL.n90 VTAIL.n89 2.84303
R703 VTAIL.n158 VTAIL.n157 2.84303
R704 VTAIL.n427 VTAIL.n426 2.84303
R705 VTAIL.n359 VTAIL.n358 2.84303
R706 VTAIL.n293 VTAIL.n292 2.84303
R707 VTAIL.n225 VTAIL.n224 2.84303
R708 VTAIL.n505 VTAIL.n484 2.71565
R709 VTAIL.n524 VTAIL.n523 2.71565
R710 VTAIL.n37 VTAIL.n16 2.71565
R711 VTAIL.n56 VTAIL.n55 2.71565
R712 VTAIL.n103 VTAIL.n82 2.71565
R713 VTAIL.n122 VTAIL.n121 2.71565
R714 VTAIL.n171 VTAIL.n150 2.71565
R715 VTAIL.n190 VTAIL.n189 2.71565
R716 VTAIL.n458 VTAIL.n457 2.71565
R717 VTAIL.n440 VTAIL.n419 2.71565
R718 VTAIL.n390 VTAIL.n389 2.71565
R719 VTAIL.n372 VTAIL.n351 2.71565
R720 VTAIL.n324 VTAIL.n323 2.71565
R721 VTAIL.n306 VTAIL.n285 2.71565
R722 VTAIL.n256 VTAIL.n255 2.71565
R723 VTAIL.n238 VTAIL.n217 2.71565
R724 VTAIL.n506 VTAIL.n482 1.93989
R725 VTAIL.n520 VTAIL.n476 1.93989
R726 VTAIL.n38 VTAIL.n14 1.93989
R727 VTAIL.n52 VTAIL.n8 1.93989
R728 VTAIL.n104 VTAIL.n80 1.93989
R729 VTAIL.n118 VTAIL.n74 1.93989
R730 VTAIL.n172 VTAIL.n148 1.93989
R731 VTAIL.n186 VTAIL.n142 1.93989
R732 VTAIL.n454 VTAIL.n410 1.93989
R733 VTAIL.n441 VTAIL.n417 1.93989
R734 VTAIL.n386 VTAIL.n342 1.93989
R735 VTAIL.n373 VTAIL.n349 1.93989
R736 VTAIL.n320 VTAIL.n276 1.93989
R737 VTAIL.n307 VTAIL.n283 1.93989
R738 VTAIL.n252 VTAIL.n208 1.93989
R739 VTAIL.n239 VTAIL.n215 1.93989
R740 VTAIL.n0 VTAIL.t6 1.64502
R741 VTAIL.n0 VTAIL.t4 1.64502
R742 VTAIL.n134 VTAIL.t11 1.64502
R743 VTAIL.n134 VTAIL.t10 1.64502
R744 VTAIL.n402 VTAIL.t14 1.64502
R745 VTAIL.n402 VTAIL.t15 1.64502
R746 VTAIL.n268 VTAIL.t1 1.64502
R747 VTAIL.n268 VTAIL.t0 1.64502
R748 VTAIL.n269 VTAIL.n267 1.44016
R749 VTAIL.n335 VTAIL.n269 1.44016
R750 VTAIL.n403 VTAIL.n401 1.44016
R751 VTAIL.n469 VTAIL.n403 1.44016
R752 VTAIL.n201 VTAIL.n135 1.44016
R753 VTAIL.n135 VTAIL.n133 1.44016
R754 VTAIL.n67 VTAIL.n1 1.44016
R755 VTAIL VTAIL.n535 1.38197
R756 VTAIL.n511 VTAIL.n509 1.16414
R757 VTAIL.n519 VTAIL.n478 1.16414
R758 VTAIL.n43 VTAIL.n41 1.16414
R759 VTAIL.n51 VTAIL.n10 1.16414
R760 VTAIL.n109 VTAIL.n107 1.16414
R761 VTAIL.n117 VTAIL.n76 1.16414
R762 VTAIL.n177 VTAIL.n175 1.16414
R763 VTAIL.n185 VTAIL.n144 1.16414
R764 VTAIL.n453 VTAIL.n412 1.16414
R765 VTAIL.n445 VTAIL.n444 1.16414
R766 VTAIL.n385 VTAIL.n344 1.16414
R767 VTAIL.n377 VTAIL.n376 1.16414
R768 VTAIL.n319 VTAIL.n278 1.16414
R769 VTAIL.n311 VTAIL.n310 1.16414
R770 VTAIL.n251 VTAIL.n210 1.16414
R771 VTAIL.n243 VTAIL.n242 1.16414
R772 VTAIL.n401 VTAIL.n335 0.470328
R773 VTAIL.n133 VTAIL.n67 0.470328
R774 VTAIL.n510 VTAIL.n480 0.388379
R775 VTAIL.n516 VTAIL.n515 0.388379
R776 VTAIL.n42 VTAIL.n12 0.388379
R777 VTAIL.n48 VTAIL.n47 0.388379
R778 VTAIL.n108 VTAIL.n78 0.388379
R779 VTAIL.n114 VTAIL.n113 0.388379
R780 VTAIL.n176 VTAIL.n146 0.388379
R781 VTAIL.n182 VTAIL.n181 0.388379
R782 VTAIL.n450 VTAIL.n449 0.388379
R783 VTAIL.n416 VTAIL.n414 0.388379
R784 VTAIL.n382 VTAIL.n381 0.388379
R785 VTAIL.n348 VTAIL.n346 0.388379
R786 VTAIL.n316 VTAIL.n315 0.388379
R787 VTAIL.n282 VTAIL.n280 0.388379
R788 VTAIL.n248 VTAIL.n247 0.388379
R789 VTAIL.n214 VTAIL.n212 0.388379
R790 VTAIL.n492 VTAIL.n487 0.155672
R791 VTAIL.n499 VTAIL.n487 0.155672
R792 VTAIL.n500 VTAIL.n499 0.155672
R793 VTAIL.n500 VTAIL.n483 0.155672
R794 VTAIL.n507 VTAIL.n483 0.155672
R795 VTAIL.n508 VTAIL.n507 0.155672
R796 VTAIL.n508 VTAIL.n479 0.155672
R797 VTAIL.n517 VTAIL.n479 0.155672
R798 VTAIL.n518 VTAIL.n517 0.155672
R799 VTAIL.n518 VTAIL.n475 0.155672
R800 VTAIL.n525 VTAIL.n475 0.155672
R801 VTAIL.n526 VTAIL.n525 0.155672
R802 VTAIL.n526 VTAIL.n471 0.155672
R803 VTAIL.n533 VTAIL.n471 0.155672
R804 VTAIL.n24 VTAIL.n19 0.155672
R805 VTAIL.n31 VTAIL.n19 0.155672
R806 VTAIL.n32 VTAIL.n31 0.155672
R807 VTAIL.n32 VTAIL.n15 0.155672
R808 VTAIL.n39 VTAIL.n15 0.155672
R809 VTAIL.n40 VTAIL.n39 0.155672
R810 VTAIL.n40 VTAIL.n11 0.155672
R811 VTAIL.n49 VTAIL.n11 0.155672
R812 VTAIL.n50 VTAIL.n49 0.155672
R813 VTAIL.n50 VTAIL.n7 0.155672
R814 VTAIL.n57 VTAIL.n7 0.155672
R815 VTAIL.n58 VTAIL.n57 0.155672
R816 VTAIL.n58 VTAIL.n3 0.155672
R817 VTAIL.n65 VTAIL.n3 0.155672
R818 VTAIL.n90 VTAIL.n85 0.155672
R819 VTAIL.n97 VTAIL.n85 0.155672
R820 VTAIL.n98 VTAIL.n97 0.155672
R821 VTAIL.n98 VTAIL.n81 0.155672
R822 VTAIL.n105 VTAIL.n81 0.155672
R823 VTAIL.n106 VTAIL.n105 0.155672
R824 VTAIL.n106 VTAIL.n77 0.155672
R825 VTAIL.n115 VTAIL.n77 0.155672
R826 VTAIL.n116 VTAIL.n115 0.155672
R827 VTAIL.n116 VTAIL.n73 0.155672
R828 VTAIL.n123 VTAIL.n73 0.155672
R829 VTAIL.n124 VTAIL.n123 0.155672
R830 VTAIL.n124 VTAIL.n69 0.155672
R831 VTAIL.n131 VTAIL.n69 0.155672
R832 VTAIL.n158 VTAIL.n153 0.155672
R833 VTAIL.n165 VTAIL.n153 0.155672
R834 VTAIL.n166 VTAIL.n165 0.155672
R835 VTAIL.n166 VTAIL.n149 0.155672
R836 VTAIL.n173 VTAIL.n149 0.155672
R837 VTAIL.n174 VTAIL.n173 0.155672
R838 VTAIL.n174 VTAIL.n145 0.155672
R839 VTAIL.n183 VTAIL.n145 0.155672
R840 VTAIL.n184 VTAIL.n183 0.155672
R841 VTAIL.n184 VTAIL.n141 0.155672
R842 VTAIL.n191 VTAIL.n141 0.155672
R843 VTAIL.n192 VTAIL.n191 0.155672
R844 VTAIL.n192 VTAIL.n137 0.155672
R845 VTAIL.n199 VTAIL.n137 0.155672
R846 VTAIL.n467 VTAIL.n405 0.155672
R847 VTAIL.n460 VTAIL.n405 0.155672
R848 VTAIL.n460 VTAIL.n459 0.155672
R849 VTAIL.n459 VTAIL.n409 0.155672
R850 VTAIL.n452 VTAIL.n409 0.155672
R851 VTAIL.n452 VTAIL.n451 0.155672
R852 VTAIL.n451 VTAIL.n413 0.155672
R853 VTAIL.n443 VTAIL.n413 0.155672
R854 VTAIL.n443 VTAIL.n442 0.155672
R855 VTAIL.n442 VTAIL.n418 0.155672
R856 VTAIL.n435 VTAIL.n418 0.155672
R857 VTAIL.n435 VTAIL.n434 0.155672
R858 VTAIL.n434 VTAIL.n422 0.155672
R859 VTAIL.n427 VTAIL.n422 0.155672
R860 VTAIL.n399 VTAIL.n337 0.155672
R861 VTAIL.n392 VTAIL.n337 0.155672
R862 VTAIL.n392 VTAIL.n391 0.155672
R863 VTAIL.n391 VTAIL.n341 0.155672
R864 VTAIL.n384 VTAIL.n341 0.155672
R865 VTAIL.n384 VTAIL.n383 0.155672
R866 VTAIL.n383 VTAIL.n345 0.155672
R867 VTAIL.n375 VTAIL.n345 0.155672
R868 VTAIL.n375 VTAIL.n374 0.155672
R869 VTAIL.n374 VTAIL.n350 0.155672
R870 VTAIL.n367 VTAIL.n350 0.155672
R871 VTAIL.n367 VTAIL.n366 0.155672
R872 VTAIL.n366 VTAIL.n354 0.155672
R873 VTAIL.n359 VTAIL.n354 0.155672
R874 VTAIL.n333 VTAIL.n271 0.155672
R875 VTAIL.n326 VTAIL.n271 0.155672
R876 VTAIL.n326 VTAIL.n325 0.155672
R877 VTAIL.n325 VTAIL.n275 0.155672
R878 VTAIL.n318 VTAIL.n275 0.155672
R879 VTAIL.n318 VTAIL.n317 0.155672
R880 VTAIL.n317 VTAIL.n279 0.155672
R881 VTAIL.n309 VTAIL.n279 0.155672
R882 VTAIL.n309 VTAIL.n308 0.155672
R883 VTAIL.n308 VTAIL.n284 0.155672
R884 VTAIL.n301 VTAIL.n284 0.155672
R885 VTAIL.n301 VTAIL.n300 0.155672
R886 VTAIL.n300 VTAIL.n288 0.155672
R887 VTAIL.n293 VTAIL.n288 0.155672
R888 VTAIL.n265 VTAIL.n203 0.155672
R889 VTAIL.n258 VTAIL.n203 0.155672
R890 VTAIL.n258 VTAIL.n257 0.155672
R891 VTAIL.n257 VTAIL.n207 0.155672
R892 VTAIL.n250 VTAIL.n207 0.155672
R893 VTAIL.n250 VTAIL.n249 0.155672
R894 VTAIL.n249 VTAIL.n211 0.155672
R895 VTAIL.n241 VTAIL.n211 0.155672
R896 VTAIL.n241 VTAIL.n240 0.155672
R897 VTAIL.n240 VTAIL.n216 0.155672
R898 VTAIL.n233 VTAIL.n216 0.155672
R899 VTAIL.n233 VTAIL.n232 0.155672
R900 VTAIL.n232 VTAIL.n220 0.155672
R901 VTAIL.n225 VTAIL.n220 0.155672
R902 VTAIL VTAIL.n1 0.0586897
R903 B.n737 B.n736 585
R904 B.n738 B.n737 585
R905 B.n295 B.n108 585
R906 B.n294 B.n293 585
R907 B.n292 B.n291 585
R908 B.n290 B.n289 585
R909 B.n288 B.n287 585
R910 B.n286 B.n285 585
R911 B.n284 B.n283 585
R912 B.n282 B.n281 585
R913 B.n280 B.n279 585
R914 B.n278 B.n277 585
R915 B.n276 B.n275 585
R916 B.n274 B.n273 585
R917 B.n272 B.n271 585
R918 B.n270 B.n269 585
R919 B.n268 B.n267 585
R920 B.n266 B.n265 585
R921 B.n264 B.n263 585
R922 B.n262 B.n261 585
R923 B.n260 B.n259 585
R924 B.n258 B.n257 585
R925 B.n256 B.n255 585
R926 B.n254 B.n253 585
R927 B.n252 B.n251 585
R928 B.n250 B.n249 585
R929 B.n248 B.n247 585
R930 B.n246 B.n245 585
R931 B.n244 B.n243 585
R932 B.n242 B.n241 585
R933 B.n240 B.n239 585
R934 B.n238 B.n237 585
R935 B.n236 B.n235 585
R936 B.n234 B.n233 585
R937 B.n232 B.n231 585
R938 B.n230 B.n229 585
R939 B.n228 B.n227 585
R940 B.n226 B.n225 585
R941 B.n224 B.n223 585
R942 B.n222 B.n221 585
R943 B.n220 B.n219 585
R944 B.n218 B.n217 585
R945 B.n216 B.n215 585
R946 B.n213 B.n212 585
R947 B.n211 B.n210 585
R948 B.n209 B.n208 585
R949 B.n207 B.n206 585
R950 B.n205 B.n204 585
R951 B.n203 B.n202 585
R952 B.n201 B.n200 585
R953 B.n199 B.n198 585
R954 B.n197 B.n196 585
R955 B.n195 B.n194 585
R956 B.n193 B.n192 585
R957 B.n191 B.n190 585
R958 B.n189 B.n188 585
R959 B.n187 B.n186 585
R960 B.n185 B.n184 585
R961 B.n183 B.n182 585
R962 B.n181 B.n180 585
R963 B.n179 B.n178 585
R964 B.n177 B.n176 585
R965 B.n175 B.n174 585
R966 B.n173 B.n172 585
R967 B.n171 B.n170 585
R968 B.n169 B.n168 585
R969 B.n167 B.n166 585
R970 B.n165 B.n164 585
R971 B.n163 B.n162 585
R972 B.n161 B.n160 585
R973 B.n159 B.n158 585
R974 B.n157 B.n156 585
R975 B.n155 B.n154 585
R976 B.n153 B.n152 585
R977 B.n151 B.n150 585
R978 B.n149 B.n148 585
R979 B.n147 B.n146 585
R980 B.n145 B.n144 585
R981 B.n143 B.n142 585
R982 B.n141 B.n140 585
R983 B.n139 B.n138 585
R984 B.n137 B.n136 585
R985 B.n135 B.n134 585
R986 B.n133 B.n132 585
R987 B.n131 B.n130 585
R988 B.n129 B.n128 585
R989 B.n127 B.n126 585
R990 B.n125 B.n124 585
R991 B.n123 B.n122 585
R992 B.n121 B.n120 585
R993 B.n119 B.n118 585
R994 B.n117 B.n116 585
R995 B.n115 B.n114 585
R996 B.n60 B.n59 585
R997 B.n735 B.n61 585
R998 B.n739 B.n61 585
R999 B.n734 B.n733 585
R1000 B.n733 B.n57 585
R1001 B.n732 B.n56 585
R1002 B.n745 B.n56 585
R1003 B.n731 B.n55 585
R1004 B.n746 B.n55 585
R1005 B.n730 B.n54 585
R1006 B.n747 B.n54 585
R1007 B.n729 B.n728 585
R1008 B.n728 B.n53 585
R1009 B.n727 B.n49 585
R1010 B.n753 B.n49 585
R1011 B.n726 B.n48 585
R1012 B.n754 B.n48 585
R1013 B.n725 B.n47 585
R1014 B.n755 B.n47 585
R1015 B.n724 B.n723 585
R1016 B.n723 B.n43 585
R1017 B.n722 B.n42 585
R1018 B.n761 B.n42 585
R1019 B.n721 B.n41 585
R1020 B.n762 B.n41 585
R1021 B.n720 B.n40 585
R1022 B.n763 B.n40 585
R1023 B.n719 B.n718 585
R1024 B.n718 B.n39 585
R1025 B.n717 B.n35 585
R1026 B.n769 B.n35 585
R1027 B.n716 B.n34 585
R1028 B.n770 B.n34 585
R1029 B.n715 B.n33 585
R1030 B.n771 B.n33 585
R1031 B.n714 B.n713 585
R1032 B.n713 B.n29 585
R1033 B.n712 B.n28 585
R1034 B.n777 B.n28 585
R1035 B.n711 B.n27 585
R1036 B.n778 B.n27 585
R1037 B.n710 B.n26 585
R1038 B.n779 B.n26 585
R1039 B.n709 B.n708 585
R1040 B.n708 B.n22 585
R1041 B.n707 B.n21 585
R1042 B.n785 B.n21 585
R1043 B.n706 B.n20 585
R1044 B.n786 B.n20 585
R1045 B.n705 B.n19 585
R1046 B.n787 B.n19 585
R1047 B.n704 B.n703 585
R1048 B.n703 B.n15 585
R1049 B.n702 B.n14 585
R1050 B.n793 B.n14 585
R1051 B.n701 B.n13 585
R1052 B.n794 B.n13 585
R1053 B.n700 B.n12 585
R1054 B.n795 B.n12 585
R1055 B.n699 B.n698 585
R1056 B.n698 B.n697 585
R1057 B.n696 B.n695 585
R1058 B.n696 B.n8 585
R1059 B.n694 B.n7 585
R1060 B.n802 B.n7 585
R1061 B.n693 B.n6 585
R1062 B.n803 B.n6 585
R1063 B.n692 B.n5 585
R1064 B.n804 B.n5 585
R1065 B.n691 B.n690 585
R1066 B.n690 B.n4 585
R1067 B.n689 B.n296 585
R1068 B.n689 B.n688 585
R1069 B.n679 B.n297 585
R1070 B.n298 B.n297 585
R1071 B.n681 B.n680 585
R1072 B.n682 B.n681 585
R1073 B.n678 B.n303 585
R1074 B.n303 B.n302 585
R1075 B.n677 B.n676 585
R1076 B.n676 B.n675 585
R1077 B.n305 B.n304 585
R1078 B.n306 B.n305 585
R1079 B.n668 B.n667 585
R1080 B.n669 B.n668 585
R1081 B.n666 B.n310 585
R1082 B.n314 B.n310 585
R1083 B.n665 B.n664 585
R1084 B.n664 B.n663 585
R1085 B.n312 B.n311 585
R1086 B.n313 B.n312 585
R1087 B.n656 B.n655 585
R1088 B.n657 B.n656 585
R1089 B.n654 B.n319 585
R1090 B.n319 B.n318 585
R1091 B.n653 B.n652 585
R1092 B.n652 B.n651 585
R1093 B.n321 B.n320 585
R1094 B.n322 B.n321 585
R1095 B.n644 B.n643 585
R1096 B.n645 B.n644 585
R1097 B.n642 B.n327 585
R1098 B.n327 B.n326 585
R1099 B.n641 B.n640 585
R1100 B.n640 B.n639 585
R1101 B.n329 B.n328 585
R1102 B.n632 B.n329 585
R1103 B.n631 B.n630 585
R1104 B.n633 B.n631 585
R1105 B.n629 B.n334 585
R1106 B.n334 B.n333 585
R1107 B.n628 B.n627 585
R1108 B.n627 B.n626 585
R1109 B.n336 B.n335 585
R1110 B.n337 B.n336 585
R1111 B.n619 B.n618 585
R1112 B.n620 B.n619 585
R1113 B.n617 B.n342 585
R1114 B.n342 B.n341 585
R1115 B.n616 B.n615 585
R1116 B.n615 B.n614 585
R1117 B.n344 B.n343 585
R1118 B.n607 B.n344 585
R1119 B.n606 B.n605 585
R1120 B.n608 B.n606 585
R1121 B.n604 B.n349 585
R1122 B.n349 B.n348 585
R1123 B.n603 B.n602 585
R1124 B.n602 B.n601 585
R1125 B.n351 B.n350 585
R1126 B.n352 B.n351 585
R1127 B.n594 B.n593 585
R1128 B.n595 B.n594 585
R1129 B.n355 B.n354 585
R1130 B.n408 B.n406 585
R1131 B.n409 B.n405 585
R1132 B.n409 B.n356 585
R1133 B.n412 B.n411 585
R1134 B.n413 B.n404 585
R1135 B.n415 B.n414 585
R1136 B.n417 B.n403 585
R1137 B.n420 B.n419 585
R1138 B.n421 B.n402 585
R1139 B.n423 B.n422 585
R1140 B.n425 B.n401 585
R1141 B.n428 B.n427 585
R1142 B.n429 B.n400 585
R1143 B.n431 B.n430 585
R1144 B.n433 B.n399 585
R1145 B.n436 B.n435 585
R1146 B.n437 B.n398 585
R1147 B.n439 B.n438 585
R1148 B.n441 B.n397 585
R1149 B.n444 B.n443 585
R1150 B.n445 B.n396 585
R1151 B.n447 B.n446 585
R1152 B.n449 B.n395 585
R1153 B.n452 B.n451 585
R1154 B.n453 B.n394 585
R1155 B.n455 B.n454 585
R1156 B.n457 B.n393 585
R1157 B.n460 B.n459 585
R1158 B.n461 B.n392 585
R1159 B.n463 B.n462 585
R1160 B.n465 B.n391 585
R1161 B.n468 B.n467 585
R1162 B.n469 B.n390 585
R1163 B.n471 B.n470 585
R1164 B.n473 B.n389 585
R1165 B.n476 B.n475 585
R1166 B.n477 B.n388 585
R1167 B.n479 B.n478 585
R1168 B.n481 B.n387 585
R1169 B.n484 B.n483 585
R1170 B.n485 B.n386 585
R1171 B.n490 B.n489 585
R1172 B.n492 B.n385 585
R1173 B.n495 B.n494 585
R1174 B.n496 B.n384 585
R1175 B.n498 B.n497 585
R1176 B.n500 B.n383 585
R1177 B.n503 B.n502 585
R1178 B.n504 B.n382 585
R1179 B.n506 B.n505 585
R1180 B.n508 B.n381 585
R1181 B.n511 B.n510 585
R1182 B.n512 B.n377 585
R1183 B.n514 B.n513 585
R1184 B.n516 B.n376 585
R1185 B.n519 B.n518 585
R1186 B.n520 B.n375 585
R1187 B.n522 B.n521 585
R1188 B.n524 B.n374 585
R1189 B.n527 B.n526 585
R1190 B.n528 B.n373 585
R1191 B.n530 B.n529 585
R1192 B.n532 B.n372 585
R1193 B.n535 B.n534 585
R1194 B.n536 B.n371 585
R1195 B.n538 B.n537 585
R1196 B.n540 B.n370 585
R1197 B.n543 B.n542 585
R1198 B.n544 B.n369 585
R1199 B.n546 B.n545 585
R1200 B.n548 B.n368 585
R1201 B.n551 B.n550 585
R1202 B.n552 B.n367 585
R1203 B.n554 B.n553 585
R1204 B.n556 B.n366 585
R1205 B.n559 B.n558 585
R1206 B.n560 B.n365 585
R1207 B.n562 B.n561 585
R1208 B.n564 B.n364 585
R1209 B.n567 B.n566 585
R1210 B.n568 B.n363 585
R1211 B.n570 B.n569 585
R1212 B.n572 B.n362 585
R1213 B.n575 B.n574 585
R1214 B.n576 B.n361 585
R1215 B.n578 B.n577 585
R1216 B.n580 B.n360 585
R1217 B.n583 B.n582 585
R1218 B.n584 B.n359 585
R1219 B.n586 B.n585 585
R1220 B.n588 B.n358 585
R1221 B.n591 B.n590 585
R1222 B.n592 B.n357 585
R1223 B.n597 B.n596 585
R1224 B.n596 B.n595 585
R1225 B.n598 B.n353 585
R1226 B.n353 B.n352 585
R1227 B.n600 B.n599 585
R1228 B.n601 B.n600 585
R1229 B.n347 B.n346 585
R1230 B.n348 B.n347 585
R1231 B.n610 B.n609 585
R1232 B.n609 B.n608 585
R1233 B.n611 B.n345 585
R1234 B.n607 B.n345 585
R1235 B.n613 B.n612 585
R1236 B.n614 B.n613 585
R1237 B.n340 B.n339 585
R1238 B.n341 B.n340 585
R1239 B.n622 B.n621 585
R1240 B.n621 B.n620 585
R1241 B.n623 B.n338 585
R1242 B.n338 B.n337 585
R1243 B.n625 B.n624 585
R1244 B.n626 B.n625 585
R1245 B.n332 B.n331 585
R1246 B.n333 B.n332 585
R1247 B.n635 B.n634 585
R1248 B.n634 B.n633 585
R1249 B.n636 B.n330 585
R1250 B.n632 B.n330 585
R1251 B.n638 B.n637 585
R1252 B.n639 B.n638 585
R1253 B.n325 B.n324 585
R1254 B.n326 B.n325 585
R1255 B.n647 B.n646 585
R1256 B.n646 B.n645 585
R1257 B.n648 B.n323 585
R1258 B.n323 B.n322 585
R1259 B.n650 B.n649 585
R1260 B.n651 B.n650 585
R1261 B.n317 B.n316 585
R1262 B.n318 B.n317 585
R1263 B.n659 B.n658 585
R1264 B.n658 B.n657 585
R1265 B.n660 B.n315 585
R1266 B.n315 B.n313 585
R1267 B.n662 B.n661 585
R1268 B.n663 B.n662 585
R1269 B.n309 B.n308 585
R1270 B.n314 B.n309 585
R1271 B.n671 B.n670 585
R1272 B.n670 B.n669 585
R1273 B.n672 B.n307 585
R1274 B.n307 B.n306 585
R1275 B.n674 B.n673 585
R1276 B.n675 B.n674 585
R1277 B.n301 B.n300 585
R1278 B.n302 B.n301 585
R1279 B.n684 B.n683 585
R1280 B.n683 B.n682 585
R1281 B.n685 B.n299 585
R1282 B.n299 B.n298 585
R1283 B.n687 B.n686 585
R1284 B.n688 B.n687 585
R1285 B.n3 B.n0 585
R1286 B.n4 B.n3 585
R1287 B.n801 B.n1 585
R1288 B.n802 B.n801 585
R1289 B.n800 B.n799 585
R1290 B.n800 B.n8 585
R1291 B.n798 B.n9 585
R1292 B.n697 B.n9 585
R1293 B.n797 B.n796 585
R1294 B.n796 B.n795 585
R1295 B.n11 B.n10 585
R1296 B.n794 B.n11 585
R1297 B.n792 B.n791 585
R1298 B.n793 B.n792 585
R1299 B.n790 B.n16 585
R1300 B.n16 B.n15 585
R1301 B.n789 B.n788 585
R1302 B.n788 B.n787 585
R1303 B.n18 B.n17 585
R1304 B.n786 B.n18 585
R1305 B.n784 B.n783 585
R1306 B.n785 B.n784 585
R1307 B.n782 B.n23 585
R1308 B.n23 B.n22 585
R1309 B.n781 B.n780 585
R1310 B.n780 B.n779 585
R1311 B.n25 B.n24 585
R1312 B.n778 B.n25 585
R1313 B.n776 B.n775 585
R1314 B.n777 B.n776 585
R1315 B.n774 B.n30 585
R1316 B.n30 B.n29 585
R1317 B.n773 B.n772 585
R1318 B.n772 B.n771 585
R1319 B.n32 B.n31 585
R1320 B.n770 B.n32 585
R1321 B.n768 B.n767 585
R1322 B.n769 B.n768 585
R1323 B.n766 B.n36 585
R1324 B.n39 B.n36 585
R1325 B.n765 B.n764 585
R1326 B.n764 B.n763 585
R1327 B.n38 B.n37 585
R1328 B.n762 B.n38 585
R1329 B.n760 B.n759 585
R1330 B.n761 B.n760 585
R1331 B.n758 B.n44 585
R1332 B.n44 B.n43 585
R1333 B.n757 B.n756 585
R1334 B.n756 B.n755 585
R1335 B.n46 B.n45 585
R1336 B.n754 B.n46 585
R1337 B.n752 B.n751 585
R1338 B.n753 B.n752 585
R1339 B.n750 B.n50 585
R1340 B.n53 B.n50 585
R1341 B.n749 B.n748 585
R1342 B.n748 B.n747 585
R1343 B.n52 B.n51 585
R1344 B.n746 B.n52 585
R1345 B.n744 B.n743 585
R1346 B.n745 B.n744 585
R1347 B.n742 B.n58 585
R1348 B.n58 B.n57 585
R1349 B.n741 B.n740 585
R1350 B.n740 B.n739 585
R1351 B.n805 B.n804 585
R1352 B.n803 B.n2 585
R1353 B.n740 B.n60 530.939
R1354 B.n737 B.n61 530.939
R1355 B.n594 B.n357 530.939
R1356 B.n596 B.n355 530.939
R1357 B.n111 B.t8 421.33
R1358 B.n109 B.t19 421.33
R1359 B.n378 B.t12 421.33
R1360 B.n486 B.t16 421.33
R1361 B.n109 B.t20 315.171
R1362 B.n378 B.t15 315.171
R1363 B.n111 B.t10 315.171
R1364 B.n486 B.t18 315.171
R1365 B.n110 B.t21 282.784
R1366 B.n379 B.t14 282.784
R1367 B.n112 B.t11 282.784
R1368 B.n487 B.t17 282.784
R1369 B.n738 B.n107 256.663
R1370 B.n738 B.n106 256.663
R1371 B.n738 B.n105 256.663
R1372 B.n738 B.n104 256.663
R1373 B.n738 B.n103 256.663
R1374 B.n738 B.n102 256.663
R1375 B.n738 B.n101 256.663
R1376 B.n738 B.n100 256.663
R1377 B.n738 B.n99 256.663
R1378 B.n738 B.n98 256.663
R1379 B.n738 B.n97 256.663
R1380 B.n738 B.n96 256.663
R1381 B.n738 B.n95 256.663
R1382 B.n738 B.n94 256.663
R1383 B.n738 B.n93 256.663
R1384 B.n738 B.n92 256.663
R1385 B.n738 B.n91 256.663
R1386 B.n738 B.n90 256.663
R1387 B.n738 B.n89 256.663
R1388 B.n738 B.n88 256.663
R1389 B.n738 B.n87 256.663
R1390 B.n738 B.n86 256.663
R1391 B.n738 B.n85 256.663
R1392 B.n738 B.n84 256.663
R1393 B.n738 B.n83 256.663
R1394 B.n738 B.n82 256.663
R1395 B.n738 B.n81 256.663
R1396 B.n738 B.n80 256.663
R1397 B.n738 B.n79 256.663
R1398 B.n738 B.n78 256.663
R1399 B.n738 B.n77 256.663
R1400 B.n738 B.n76 256.663
R1401 B.n738 B.n75 256.663
R1402 B.n738 B.n74 256.663
R1403 B.n738 B.n73 256.663
R1404 B.n738 B.n72 256.663
R1405 B.n738 B.n71 256.663
R1406 B.n738 B.n70 256.663
R1407 B.n738 B.n69 256.663
R1408 B.n738 B.n68 256.663
R1409 B.n738 B.n67 256.663
R1410 B.n738 B.n66 256.663
R1411 B.n738 B.n65 256.663
R1412 B.n738 B.n64 256.663
R1413 B.n738 B.n63 256.663
R1414 B.n738 B.n62 256.663
R1415 B.n407 B.n356 256.663
R1416 B.n410 B.n356 256.663
R1417 B.n416 B.n356 256.663
R1418 B.n418 B.n356 256.663
R1419 B.n424 B.n356 256.663
R1420 B.n426 B.n356 256.663
R1421 B.n432 B.n356 256.663
R1422 B.n434 B.n356 256.663
R1423 B.n440 B.n356 256.663
R1424 B.n442 B.n356 256.663
R1425 B.n448 B.n356 256.663
R1426 B.n450 B.n356 256.663
R1427 B.n456 B.n356 256.663
R1428 B.n458 B.n356 256.663
R1429 B.n464 B.n356 256.663
R1430 B.n466 B.n356 256.663
R1431 B.n472 B.n356 256.663
R1432 B.n474 B.n356 256.663
R1433 B.n480 B.n356 256.663
R1434 B.n482 B.n356 256.663
R1435 B.n491 B.n356 256.663
R1436 B.n493 B.n356 256.663
R1437 B.n499 B.n356 256.663
R1438 B.n501 B.n356 256.663
R1439 B.n507 B.n356 256.663
R1440 B.n509 B.n356 256.663
R1441 B.n515 B.n356 256.663
R1442 B.n517 B.n356 256.663
R1443 B.n523 B.n356 256.663
R1444 B.n525 B.n356 256.663
R1445 B.n531 B.n356 256.663
R1446 B.n533 B.n356 256.663
R1447 B.n539 B.n356 256.663
R1448 B.n541 B.n356 256.663
R1449 B.n547 B.n356 256.663
R1450 B.n549 B.n356 256.663
R1451 B.n555 B.n356 256.663
R1452 B.n557 B.n356 256.663
R1453 B.n563 B.n356 256.663
R1454 B.n565 B.n356 256.663
R1455 B.n571 B.n356 256.663
R1456 B.n573 B.n356 256.663
R1457 B.n579 B.n356 256.663
R1458 B.n581 B.n356 256.663
R1459 B.n587 B.n356 256.663
R1460 B.n589 B.n356 256.663
R1461 B.n807 B.n806 256.663
R1462 B.n116 B.n115 163.367
R1463 B.n120 B.n119 163.367
R1464 B.n124 B.n123 163.367
R1465 B.n128 B.n127 163.367
R1466 B.n132 B.n131 163.367
R1467 B.n136 B.n135 163.367
R1468 B.n140 B.n139 163.367
R1469 B.n144 B.n143 163.367
R1470 B.n148 B.n147 163.367
R1471 B.n152 B.n151 163.367
R1472 B.n156 B.n155 163.367
R1473 B.n160 B.n159 163.367
R1474 B.n164 B.n163 163.367
R1475 B.n168 B.n167 163.367
R1476 B.n172 B.n171 163.367
R1477 B.n176 B.n175 163.367
R1478 B.n180 B.n179 163.367
R1479 B.n184 B.n183 163.367
R1480 B.n188 B.n187 163.367
R1481 B.n192 B.n191 163.367
R1482 B.n196 B.n195 163.367
R1483 B.n200 B.n199 163.367
R1484 B.n204 B.n203 163.367
R1485 B.n208 B.n207 163.367
R1486 B.n212 B.n211 163.367
R1487 B.n217 B.n216 163.367
R1488 B.n221 B.n220 163.367
R1489 B.n225 B.n224 163.367
R1490 B.n229 B.n228 163.367
R1491 B.n233 B.n232 163.367
R1492 B.n237 B.n236 163.367
R1493 B.n241 B.n240 163.367
R1494 B.n245 B.n244 163.367
R1495 B.n249 B.n248 163.367
R1496 B.n253 B.n252 163.367
R1497 B.n257 B.n256 163.367
R1498 B.n261 B.n260 163.367
R1499 B.n265 B.n264 163.367
R1500 B.n269 B.n268 163.367
R1501 B.n273 B.n272 163.367
R1502 B.n277 B.n276 163.367
R1503 B.n281 B.n280 163.367
R1504 B.n285 B.n284 163.367
R1505 B.n289 B.n288 163.367
R1506 B.n293 B.n292 163.367
R1507 B.n737 B.n108 163.367
R1508 B.n594 B.n351 163.367
R1509 B.n602 B.n351 163.367
R1510 B.n602 B.n349 163.367
R1511 B.n606 B.n349 163.367
R1512 B.n606 B.n344 163.367
R1513 B.n615 B.n344 163.367
R1514 B.n615 B.n342 163.367
R1515 B.n619 B.n342 163.367
R1516 B.n619 B.n336 163.367
R1517 B.n627 B.n336 163.367
R1518 B.n627 B.n334 163.367
R1519 B.n631 B.n334 163.367
R1520 B.n631 B.n329 163.367
R1521 B.n640 B.n329 163.367
R1522 B.n640 B.n327 163.367
R1523 B.n644 B.n327 163.367
R1524 B.n644 B.n321 163.367
R1525 B.n652 B.n321 163.367
R1526 B.n652 B.n319 163.367
R1527 B.n656 B.n319 163.367
R1528 B.n656 B.n312 163.367
R1529 B.n664 B.n312 163.367
R1530 B.n664 B.n310 163.367
R1531 B.n668 B.n310 163.367
R1532 B.n668 B.n305 163.367
R1533 B.n676 B.n305 163.367
R1534 B.n676 B.n303 163.367
R1535 B.n681 B.n303 163.367
R1536 B.n681 B.n297 163.367
R1537 B.n689 B.n297 163.367
R1538 B.n690 B.n689 163.367
R1539 B.n690 B.n5 163.367
R1540 B.n6 B.n5 163.367
R1541 B.n7 B.n6 163.367
R1542 B.n696 B.n7 163.367
R1543 B.n698 B.n696 163.367
R1544 B.n698 B.n12 163.367
R1545 B.n13 B.n12 163.367
R1546 B.n14 B.n13 163.367
R1547 B.n703 B.n14 163.367
R1548 B.n703 B.n19 163.367
R1549 B.n20 B.n19 163.367
R1550 B.n21 B.n20 163.367
R1551 B.n708 B.n21 163.367
R1552 B.n708 B.n26 163.367
R1553 B.n27 B.n26 163.367
R1554 B.n28 B.n27 163.367
R1555 B.n713 B.n28 163.367
R1556 B.n713 B.n33 163.367
R1557 B.n34 B.n33 163.367
R1558 B.n35 B.n34 163.367
R1559 B.n718 B.n35 163.367
R1560 B.n718 B.n40 163.367
R1561 B.n41 B.n40 163.367
R1562 B.n42 B.n41 163.367
R1563 B.n723 B.n42 163.367
R1564 B.n723 B.n47 163.367
R1565 B.n48 B.n47 163.367
R1566 B.n49 B.n48 163.367
R1567 B.n728 B.n49 163.367
R1568 B.n728 B.n54 163.367
R1569 B.n55 B.n54 163.367
R1570 B.n56 B.n55 163.367
R1571 B.n733 B.n56 163.367
R1572 B.n733 B.n61 163.367
R1573 B.n409 B.n408 163.367
R1574 B.n411 B.n409 163.367
R1575 B.n415 B.n404 163.367
R1576 B.n419 B.n417 163.367
R1577 B.n423 B.n402 163.367
R1578 B.n427 B.n425 163.367
R1579 B.n431 B.n400 163.367
R1580 B.n435 B.n433 163.367
R1581 B.n439 B.n398 163.367
R1582 B.n443 B.n441 163.367
R1583 B.n447 B.n396 163.367
R1584 B.n451 B.n449 163.367
R1585 B.n455 B.n394 163.367
R1586 B.n459 B.n457 163.367
R1587 B.n463 B.n392 163.367
R1588 B.n467 B.n465 163.367
R1589 B.n471 B.n390 163.367
R1590 B.n475 B.n473 163.367
R1591 B.n479 B.n388 163.367
R1592 B.n483 B.n481 163.367
R1593 B.n490 B.n386 163.367
R1594 B.n494 B.n492 163.367
R1595 B.n498 B.n384 163.367
R1596 B.n502 B.n500 163.367
R1597 B.n506 B.n382 163.367
R1598 B.n510 B.n508 163.367
R1599 B.n514 B.n377 163.367
R1600 B.n518 B.n516 163.367
R1601 B.n522 B.n375 163.367
R1602 B.n526 B.n524 163.367
R1603 B.n530 B.n373 163.367
R1604 B.n534 B.n532 163.367
R1605 B.n538 B.n371 163.367
R1606 B.n542 B.n540 163.367
R1607 B.n546 B.n369 163.367
R1608 B.n550 B.n548 163.367
R1609 B.n554 B.n367 163.367
R1610 B.n558 B.n556 163.367
R1611 B.n562 B.n365 163.367
R1612 B.n566 B.n564 163.367
R1613 B.n570 B.n363 163.367
R1614 B.n574 B.n572 163.367
R1615 B.n578 B.n361 163.367
R1616 B.n582 B.n580 163.367
R1617 B.n586 B.n359 163.367
R1618 B.n590 B.n588 163.367
R1619 B.n596 B.n353 163.367
R1620 B.n600 B.n353 163.367
R1621 B.n600 B.n347 163.367
R1622 B.n609 B.n347 163.367
R1623 B.n609 B.n345 163.367
R1624 B.n613 B.n345 163.367
R1625 B.n613 B.n340 163.367
R1626 B.n621 B.n340 163.367
R1627 B.n621 B.n338 163.367
R1628 B.n625 B.n338 163.367
R1629 B.n625 B.n332 163.367
R1630 B.n634 B.n332 163.367
R1631 B.n634 B.n330 163.367
R1632 B.n638 B.n330 163.367
R1633 B.n638 B.n325 163.367
R1634 B.n646 B.n325 163.367
R1635 B.n646 B.n323 163.367
R1636 B.n650 B.n323 163.367
R1637 B.n650 B.n317 163.367
R1638 B.n658 B.n317 163.367
R1639 B.n658 B.n315 163.367
R1640 B.n662 B.n315 163.367
R1641 B.n662 B.n309 163.367
R1642 B.n670 B.n309 163.367
R1643 B.n670 B.n307 163.367
R1644 B.n674 B.n307 163.367
R1645 B.n674 B.n301 163.367
R1646 B.n683 B.n301 163.367
R1647 B.n683 B.n299 163.367
R1648 B.n687 B.n299 163.367
R1649 B.n687 B.n3 163.367
R1650 B.n805 B.n3 163.367
R1651 B.n801 B.n2 163.367
R1652 B.n801 B.n800 163.367
R1653 B.n800 B.n9 163.367
R1654 B.n796 B.n9 163.367
R1655 B.n796 B.n11 163.367
R1656 B.n792 B.n11 163.367
R1657 B.n792 B.n16 163.367
R1658 B.n788 B.n16 163.367
R1659 B.n788 B.n18 163.367
R1660 B.n784 B.n18 163.367
R1661 B.n784 B.n23 163.367
R1662 B.n780 B.n23 163.367
R1663 B.n780 B.n25 163.367
R1664 B.n776 B.n25 163.367
R1665 B.n776 B.n30 163.367
R1666 B.n772 B.n30 163.367
R1667 B.n772 B.n32 163.367
R1668 B.n768 B.n32 163.367
R1669 B.n768 B.n36 163.367
R1670 B.n764 B.n36 163.367
R1671 B.n764 B.n38 163.367
R1672 B.n760 B.n38 163.367
R1673 B.n760 B.n44 163.367
R1674 B.n756 B.n44 163.367
R1675 B.n756 B.n46 163.367
R1676 B.n752 B.n46 163.367
R1677 B.n752 B.n50 163.367
R1678 B.n748 B.n50 163.367
R1679 B.n748 B.n52 163.367
R1680 B.n744 B.n52 163.367
R1681 B.n744 B.n58 163.367
R1682 B.n740 B.n58 163.367
R1683 B.n595 B.n356 85.7643
R1684 B.n739 B.n738 85.7643
R1685 B.n62 B.n60 71.676
R1686 B.n116 B.n63 71.676
R1687 B.n120 B.n64 71.676
R1688 B.n124 B.n65 71.676
R1689 B.n128 B.n66 71.676
R1690 B.n132 B.n67 71.676
R1691 B.n136 B.n68 71.676
R1692 B.n140 B.n69 71.676
R1693 B.n144 B.n70 71.676
R1694 B.n148 B.n71 71.676
R1695 B.n152 B.n72 71.676
R1696 B.n156 B.n73 71.676
R1697 B.n160 B.n74 71.676
R1698 B.n164 B.n75 71.676
R1699 B.n168 B.n76 71.676
R1700 B.n172 B.n77 71.676
R1701 B.n176 B.n78 71.676
R1702 B.n180 B.n79 71.676
R1703 B.n184 B.n80 71.676
R1704 B.n188 B.n81 71.676
R1705 B.n192 B.n82 71.676
R1706 B.n196 B.n83 71.676
R1707 B.n200 B.n84 71.676
R1708 B.n204 B.n85 71.676
R1709 B.n208 B.n86 71.676
R1710 B.n212 B.n87 71.676
R1711 B.n217 B.n88 71.676
R1712 B.n221 B.n89 71.676
R1713 B.n225 B.n90 71.676
R1714 B.n229 B.n91 71.676
R1715 B.n233 B.n92 71.676
R1716 B.n237 B.n93 71.676
R1717 B.n241 B.n94 71.676
R1718 B.n245 B.n95 71.676
R1719 B.n249 B.n96 71.676
R1720 B.n253 B.n97 71.676
R1721 B.n257 B.n98 71.676
R1722 B.n261 B.n99 71.676
R1723 B.n265 B.n100 71.676
R1724 B.n269 B.n101 71.676
R1725 B.n273 B.n102 71.676
R1726 B.n277 B.n103 71.676
R1727 B.n281 B.n104 71.676
R1728 B.n285 B.n105 71.676
R1729 B.n289 B.n106 71.676
R1730 B.n293 B.n107 71.676
R1731 B.n108 B.n107 71.676
R1732 B.n292 B.n106 71.676
R1733 B.n288 B.n105 71.676
R1734 B.n284 B.n104 71.676
R1735 B.n280 B.n103 71.676
R1736 B.n276 B.n102 71.676
R1737 B.n272 B.n101 71.676
R1738 B.n268 B.n100 71.676
R1739 B.n264 B.n99 71.676
R1740 B.n260 B.n98 71.676
R1741 B.n256 B.n97 71.676
R1742 B.n252 B.n96 71.676
R1743 B.n248 B.n95 71.676
R1744 B.n244 B.n94 71.676
R1745 B.n240 B.n93 71.676
R1746 B.n236 B.n92 71.676
R1747 B.n232 B.n91 71.676
R1748 B.n228 B.n90 71.676
R1749 B.n224 B.n89 71.676
R1750 B.n220 B.n88 71.676
R1751 B.n216 B.n87 71.676
R1752 B.n211 B.n86 71.676
R1753 B.n207 B.n85 71.676
R1754 B.n203 B.n84 71.676
R1755 B.n199 B.n83 71.676
R1756 B.n195 B.n82 71.676
R1757 B.n191 B.n81 71.676
R1758 B.n187 B.n80 71.676
R1759 B.n183 B.n79 71.676
R1760 B.n179 B.n78 71.676
R1761 B.n175 B.n77 71.676
R1762 B.n171 B.n76 71.676
R1763 B.n167 B.n75 71.676
R1764 B.n163 B.n74 71.676
R1765 B.n159 B.n73 71.676
R1766 B.n155 B.n72 71.676
R1767 B.n151 B.n71 71.676
R1768 B.n147 B.n70 71.676
R1769 B.n143 B.n69 71.676
R1770 B.n139 B.n68 71.676
R1771 B.n135 B.n67 71.676
R1772 B.n131 B.n66 71.676
R1773 B.n127 B.n65 71.676
R1774 B.n123 B.n64 71.676
R1775 B.n119 B.n63 71.676
R1776 B.n115 B.n62 71.676
R1777 B.n407 B.n355 71.676
R1778 B.n411 B.n410 71.676
R1779 B.n416 B.n415 71.676
R1780 B.n419 B.n418 71.676
R1781 B.n424 B.n423 71.676
R1782 B.n427 B.n426 71.676
R1783 B.n432 B.n431 71.676
R1784 B.n435 B.n434 71.676
R1785 B.n440 B.n439 71.676
R1786 B.n443 B.n442 71.676
R1787 B.n448 B.n447 71.676
R1788 B.n451 B.n450 71.676
R1789 B.n456 B.n455 71.676
R1790 B.n459 B.n458 71.676
R1791 B.n464 B.n463 71.676
R1792 B.n467 B.n466 71.676
R1793 B.n472 B.n471 71.676
R1794 B.n475 B.n474 71.676
R1795 B.n480 B.n479 71.676
R1796 B.n483 B.n482 71.676
R1797 B.n491 B.n490 71.676
R1798 B.n494 B.n493 71.676
R1799 B.n499 B.n498 71.676
R1800 B.n502 B.n501 71.676
R1801 B.n507 B.n506 71.676
R1802 B.n510 B.n509 71.676
R1803 B.n515 B.n514 71.676
R1804 B.n518 B.n517 71.676
R1805 B.n523 B.n522 71.676
R1806 B.n526 B.n525 71.676
R1807 B.n531 B.n530 71.676
R1808 B.n534 B.n533 71.676
R1809 B.n539 B.n538 71.676
R1810 B.n542 B.n541 71.676
R1811 B.n547 B.n546 71.676
R1812 B.n550 B.n549 71.676
R1813 B.n555 B.n554 71.676
R1814 B.n558 B.n557 71.676
R1815 B.n563 B.n562 71.676
R1816 B.n566 B.n565 71.676
R1817 B.n571 B.n570 71.676
R1818 B.n574 B.n573 71.676
R1819 B.n579 B.n578 71.676
R1820 B.n582 B.n581 71.676
R1821 B.n587 B.n586 71.676
R1822 B.n590 B.n589 71.676
R1823 B.n408 B.n407 71.676
R1824 B.n410 B.n404 71.676
R1825 B.n417 B.n416 71.676
R1826 B.n418 B.n402 71.676
R1827 B.n425 B.n424 71.676
R1828 B.n426 B.n400 71.676
R1829 B.n433 B.n432 71.676
R1830 B.n434 B.n398 71.676
R1831 B.n441 B.n440 71.676
R1832 B.n442 B.n396 71.676
R1833 B.n449 B.n448 71.676
R1834 B.n450 B.n394 71.676
R1835 B.n457 B.n456 71.676
R1836 B.n458 B.n392 71.676
R1837 B.n465 B.n464 71.676
R1838 B.n466 B.n390 71.676
R1839 B.n473 B.n472 71.676
R1840 B.n474 B.n388 71.676
R1841 B.n481 B.n480 71.676
R1842 B.n482 B.n386 71.676
R1843 B.n492 B.n491 71.676
R1844 B.n493 B.n384 71.676
R1845 B.n500 B.n499 71.676
R1846 B.n501 B.n382 71.676
R1847 B.n508 B.n507 71.676
R1848 B.n509 B.n377 71.676
R1849 B.n516 B.n515 71.676
R1850 B.n517 B.n375 71.676
R1851 B.n524 B.n523 71.676
R1852 B.n525 B.n373 71.676
R1853 B.n532 B.n531 71.676
R1854 B.n533 B.n371 71.676
R1855 B.n540 B.n539 71.676
R1856 B.n541 B.n369 71.676
R1857 B.n548 B.n547 71.676
R1858 B.n549 B.n367 71.676
R1859 B.n556 B.n555 71.676
R1860 B.n557 B.n365 71.676
R1861 B.n564 B.n563 71.676
R1862 B.n565 B.n363 71.676
R1863 B.n572 B.n571 71.676
R1864 B.n573 B.n361 71.676
R1865 B.n580 B.n579 71.676
R1866 B.n581 B.n359 71.676
R1867 B.n588 B.n587 71.676
R1868 B.n589 B.n357 71.676
R1869 B.n806 B.n805 71.676
R1870 B.n806 B.n2 71.676
R1871 B.n113 B.n112 59.5399
R1872 B.n214 B.n110 59.5399
R1873 B.n380 B.n379 59.5399
R1874 B.n488 B.n487 59.5399
R1875 B.n595 B.n352 43.2
R1876 B.n601 B.n352 43.2
R1877 B.n601 B.n348 43.2
R1878 B.n608 B.n348 43.2
R1879 B.n608 B.n607 43.2
R1880 B.n614 B.n341 43.2
R1881 B.n620 B.n341 43.2
R1882 B.n620 B.n337 43.2
R1883 B.n626 B.n337 43.2
R1884 B.n626 B.n333 43.2
R1885 B.n633 B.n333 43.2
R1886 B.n633 B.n632 43.2
R1887 B.n639 B.n326 43.2
R1888 B.n645 B.n326 43.2
R1889 B.n645 B.n322 43.2
R1890 B.n651 B.n322 43.2
R1891 B.n657 B.n318 43.2
R1892 B.n657 B.n313 43.2
R1893 B.n663 B.n313 43.2
R1894 B.n663 B.n314 43.2
R1895 B.n669 B.n306 43.2
R1896 B.n675 B.n306 43.2
R1897 B.n675 B.n302 43.2
R1898 B.n682 B.n302 43.2
R1899 B.n688 B.n298 43.2
R1900 B.n688 B.n4 43.2
R1901 B.n804 B.n4 43.2
R1902 B.n804 B.n803 43.2
R1903 B.n803 B.n802 43.2
R1904 B.n802 B.n8 43.2
R1905 B.n697 B.n8 43.2
R1906 B.n795 B.n794 43.2
R1907 B.n794 B.n793 43.2
R1908 B.n793 B.n15 43.2
R1909 B.n787 B.n15 43.2
R1910 B.n786 B.n785 43.2
R1911 B.n785 B.n22 43.2
R1912 B.n779 B.n22 43.2
R1913 B.n779 B.n778 43.2
R1914 B.n777 B.n29 43.2
R1915 B.n771 B.n29 43.2
R1916 B.n771 B.n770 43.2
R1917 B.n770 B.n769 43.2
R1918 B.n763 B.n39 43.2
R1919 B.n763 B.n762 43.2
R1920 B.n762 B.n761 43.2
R1921 B.n761 B.n43 43.2
R1922 B.n755 B.n43 43.2
R1923 B.n755 B.n754 43.2
R1924 B.n754 B.n753 43.2
R1925 B.n747 B.n53 43.2
R1926 B.n747 B.n746 43.2
R1927 B.n746 B.n745 43.2
R1928 B.n745 B.n57 43.2
R1929 B.n739 B.n57 43.2
R1930 B.n597 B.n354 34.4981
R1931 B.n593 B.n592 34.4981
R1932 B.n736 B.n735 34.4981
R1933 B.n741 B.n59 34.4981
R1934 B.n112 B.n111 32.3884
R1935 B.n110 B.n109 32.3884
R1936 B.n379 B.n378 32.3884
R1937 B.n487 B.n486 32.3884
R1938 B.n632 B.t7 30.4943
R1939 B.n39 B.t2 30.4943
R1940 B.n651 B.t1 26.6826
R1941 B.t4 B.n777 26.6826
R1942 B.n607 B.t13 25.412
R1943 B.n53 B.t9 25.412
R1944 B.t3 B.n298 24.1414
R1945 B.n697 B.t5 24.1414
R1946 B.n314 B.t0 22.8708
R1947 B.t6 B.n786 22.8708
R1948 B.n669 B.t0 20.3297
R1949 B.n787 B.t6 20.3297
R1950 B.n682 B.t3 19.0591
R1951 B.n795 B.t5 19.0591
R1952 B B.n807 18.0485
R1953 B.n614 B.t13 17.7885
R1954 B.n753 B.t9 17.7885
R1955 B.t1 B.n318 16.518
R1956 B.n778 B.t4 16.518
R1957 B.n639 B.t7 12.7062
R1958 B.n769 B.t2 12.7062
R1959 B.n598 B.n597 10.6151
R1960 B.n599 B.n598 10.6151
R1961 B.n599 B.n346 10.6151
R1962 B.n610 B.n346 10.6151
R1963 B.n611 B.n610 10.6151
R1964 B.n612 B.n611 10.6151
R1965 B.n612 B.n339 10.6151
R1966 B.n622 B.n339 10.6151
R1967 B.n623 B.n622 10.6151
R1968 B.n624 B.n623 10.6151
R1969 B.n624 B.n331 10.6151
R1970 B.n635 B.n331 10.6151
R1971 B.n636 B.n635 10.6151
R1972 B.n637 B.n636 10.6151
R1973 B.n637 B.n324 10.6151
R1974 B.n647 B.n324 10.6151
R1975 B.n648 B.n647 10.6151
R1976 B.n649 B.n648 10.6151
R1977 B.n649 B.n316 10.6151
R1978 B.n659 B.n316 10.6151
R1979 B.n660 B.n659 10.6151
R1980 B.n661 B.n660 10.6151
R1981 B.n661 B.n308 10.6151
R1982 B.n671 B.n308 10.6151
R1983 B.n672 B.n671 10.6151
R1984 B.n673 B.n672 10.6151
R1985 B.n673 B.n300 10.6151
R1986 B.n684 B.n300 10.6151
R1987 B.n685 B.n684 10.6151
R1988 B.n686 B.n685 10.6151
R1989 B.n686 B.n0 10.6151
R1990 B.n406 B.n354 10.6151
R1991 B.n406 B.n405 10.6151
R1992 B.n412 B.n405 10.6151
R1993 B.n413 B.n412 10.6151
R1994 B.n414 B.n413 10.6151
R1995 B.n414 B.n403 10.6151
R1996 B.n420 B.n403 10.6151
R1997 B.n421 B.n420 10.6151
R1998 B.n422 B.n421 10.6151
R1999 B.n422 B.n401 10.6151
R2000 B.n428 B.n401 10.6151
R2001 B.n429 B.n428 10.6151
R2002 B.n430 B.n429 10.6151
R2003 B.n430 B.n399 10.6151
R2004 B.n436 B.n399 10.6151
R2005 B.n437 B.n436 10.6151
R2006 B.n438 B.n437 10.6151
R2007 B.n438 B.n397 10.6151
R2008 B.n444 B.n397 10.6151
R2009 B.n445 B.n444 10.6151
R2010 B.n446 B.n445 10.6151
R2011 B.n446 B.n395 10.6151
R2012 B.n452 B.n395 10.6151
R2013 B.n453 B.n452 10.6151
R2014 B.n454 B.n453 10.6151
R2015 B.n454 B.n393 10.6151
R2016 B.n460 B.n393 10.6151
R2017 B.n461 B.n460 10.6151
R2018 B.n462 B.n461 10.6151
R2019 B.n462 B.n391 10.6151
R2020 B.n468 B.n391 10.6151
R2021 B.n469 B.n468 10.6151
R2022 B.n470 B.n469 10.6151
R2023 B.n470 B.n389 10.6151
R2024 B.n476 B.n389 10.6151
R2025 B.n477 B.n476 10.6151
R2026 B.n478 B.n477 10.6151
R2027 B.n478 B.n387 10.6151
R2028 B.n484 B.n387 10.6151
R2029 B.n485 B.n484 10.6151
R2030 B.n489 B.n485 10.6151
R2031 B.n495 B.n385 10.6151
R2032 B.n496 B.n495 10.6151
R2033 B.n497 B.n496 10.6151
R2034 B.n497 B.n383 10.6151
R2035 B.n503 B.n383 10.6151
R2036 B.n504 B.n503 10.6151
R2037 B.n505 B.n504 10.6151
R2038 B.n505 B.n381 10.6151
R2039 B.n512 B.n511 10.6151
R2040 B.n513 B.n512 10.6151
R2041 B.n513 B.n376 10.6151
R2042 B.n519 B.n376 10.6151
R2043 B.n520 B.n519 10.6151
R2044 B.n521 B.n520 10.6151
R2045 B.n521 B.n374 10.6151
R2046 B.n527 B.n374 10.6151
R2047 B.n528 B.n527 10.6151
R2048 B.n529 B.n528 10.6151
R2049 B.n529 B.n372 10.6151
R2050 B.n535 B.n372 10.6151
R2051 B.n536 B.n535 10.6151
R2052 B.n537 B.n536 10.6151
R2053 B.n537 B.n370 10.6151
R2054 B.n543 B.n370 10.6151
R2055 B.n544 B.n543 10.6151
R2056 B.n545 B.n544 10.6151
R2057 B.n545 B.n368 10.6151
R2058 B.n551 B.n368 10.6151
R2059 B.n552 B.n551 10.6151
R2060 B.n553 B.n552 10.6151
R2061 B.n553 B.n366 10.6151
R2062 B.n559 B.n366 10.6151
R2063 B.n560 B.n559 10.6151
R2064 B.n561 B.n560 10.6151
R2065 B.n561 B.n364 10.6151
R2066 B.n567 B.n364 10.6151
R2067 B.n568 B.n567 10.6151
R2068 B.n569 B.n568 10.6151
R2069 B.n569 B.n362 10.6151
R2070 B.n575 B.n362 10.6151
R2071 B.n576 B.n575 10.6151
R2072 B.n577 B.n576 10.6151
R2073 B.n577 B.n360 10.6151
R2074 B.n583 B.n360 10.6151
R2075 B.n584 B.n583 10.6151
R2076 B.n585 B.n584 10.6151
R2077 B.n585 B.n358 10.6151
R2078 B.n591 B.n358 10.6151
R2079 B.n592 B.n591 10.6151
R2080 B.n593 B.n350 10.6151
R2081 B.n603 B.n350 10.6151
R2082 B.n604 B.n603 10.6151
R2083 B.n605 B.n604 10.6151
R2084 B.n605 B.n343 10.6151
R2085 B.n616 B.n343 10.6151
R2086 B.n617 B.n616 10.6151
R2087 B.n618 B.n617 10.6151
R2088 B.n618 B.n335 10.6151
R2089 B.n628 B.n335 10.6151
R2090 B.n629 B.n628 10.6151
R2091 B.n630 B.n629 10.6151
R2092 B.n630 B.n328 10.6151
R2093 B.n641 B.n328 10.6151
R2094 B.n642 B.n641 10.6151
R2095 B.n643 B.n642 10.6151
R2096 B.n643 B.n320 10.6151
R2097 B.n653 B.n320 10.6151
R2098 B.n654 B.n653 10.6151
R2099 B.n655 B.n654 10.6151
R2100 B.n655 B.n311 10.6151
R2101 B.n665 B.n311 10.6151
R2102 B.n666 B.n665 10.6151
R2103 B.n667 B.n666 10.6151
R2104 B.n667 B.n304 10.6151
R2105 B.n677 B.n304 10.6151
R2106 B.n678 B.n677 10.6151
R2107 B.n680 B.n678 10.6151
R2108 B.n680 B.n679 10.6151
R2109 B.n679 B.n296 10.6151
R2110 B.n691 B.n296 10.6151
R2111 B.n692 B.n691 10.6151
R2112 B.n693 B.n692 10.6151
R2113 B.n694 B.n693 10.6151
R2114 B.n695 B.n694 10.6151
R2115 B.n699 B.n695 10.6151
R2116 B.n700 B.n699 10.6151
R2117 B.n701 B.n700 10.6151
R2118 B.n702 B.n701 10.6151
R2119 B.n704 B.n702 10.6151
R2120 B.n705 B.n704 10.6151
R2121 B.n706 B.n705 10.6151
R2122 B.n707 B.n706 10.6151
R2123 B.n709 B.n707 10.6151
R2124 B.n710 B.n709 10.6151
R2125 B.n711 B.n710 10.6151
R2126 B.n712 B.n711 10.6151
R2127 B.n714 B.n712 10.6151
R2128 B.n715 B.n714 10.6151
R2129 B.n716 B.n715 10.6151
R2130 B.n717 B.n716 10.6151
R2131 B.n719 B.n717 10.6151
R2132 B.n720 B.n719 10.6151
R2133 B.n721 B.n720 10.6151
R2134 B.n722 B.n721 10.6151
R2135 B.n724 B.n722 10.6151
R2136 B.n725 B.n724 10.6151
R2137 B.n726 B.n725 10.6151
R2138 B.n727 B.n726 10.6151
R2139 B.n729 B.n727 10.6151
R2140 B.n730 B.n729 10.6151
R2141 B.n731 B.n730 10.6151
R2142 B.n732 B.n731 10.6151
R2143 B.n734 B.n732 10.6151
R2144 B.n735 B.n734 10.6151
R2145 B.n799 B.n1 10.6151
R2146 B.n799 B.n798 10.6151
R2147 B.n798 B.n797 10.6151
R2148 B.n797 B.n10 10.6151
R2149 B.n791 B.n10 10.6151
R2150 B.n791 B.n790 10.6151
R2151 B.n790 B.n789 10.6151
R2152 B.n789 B.n17 10.6151
R2153 B.n783 B.n17 10.6151
R2154 B.n783 B.n782 10.6151
R2155 B.n782 B.n781 10.6151
R2156 B.n781 B.n24 10.6151
R2157 B.n775 B.n24 10.6151
R2158 B.n775 B.n774 10.6151
R2159 B.n774 B.n773 10.6151
R2160 B.n773 B.n31 10.6151
R2161 B.n767 B.n31 10.6151
R2162 B.n767 B.n766 10.6151
R2163 B.n766 B.n765 10.6151
R2164 B.n765 B.n37 10.6151
R2165 B.n759 B.n37 10.6151
R2166 B.n759 B.n758 10.6151
R2167 B.n758 B.n757 10.6151
R2168 B.n757 B.n45 10.6151
R2169 B.n751 B.n45 10.6151
R2170 B.n751 B.n750 10.6151
R2171 B.n750 B.n749 10.6151
R2172 B.n749 B.n51 10.6151
R2173 B.n743 B.n51 10.6151
R2174 B.n743 B.n742 10.6151
R2175 B.n742 B.n741 10.6151
R2176 B.n114 B.n59 10.6151
R2177 B.n117 B.n114 10.6151
R2178 B.n118 B.n117 10.6151
R2179 B.n121 B.n118 10.6151
R2180 B.n122 B.n121 10.6151
R2181 B.n125 B.n122 10.6151
R2182 B.n126 B.n125 10.6151
R2183 B.n129 B.n126 10.6151
R2184 B.n130 B.n129 10.6151
R2185 B.n133 B.n130 10.6151
R2186 B.n134 B.n133 10.6151
R2187 B.n137 B.n134 10.6151
R2188 B.n138 B.n137 10.6151
R2189 B.n141 B.n138 10.6151
R2190 B.n142 B.n141 10.6151
R2191 B.n145 B.n142 10.6151
R2192 B.n146 B.n145 10.6151
R2193 B.n149 B.n146 10.6151
R2194 B.n150 B.n149 10.6151
R2195 B.n153 B.n150 10.6151
R2196 B.n154 B.n153 10.6151
R2197 B.n157 B.n154 10.6151
R2198 B.n158 B.n157 10.6151
R2199 B.n161 B.n158 10.6151
R2200 B.n162 B.n161 10.6151
R2201 B.n165 B.n162 10.6151
R2202 B.n166 B.n165 10.6151
R2203 B.n169 B.n166 10.6151
R2204 B.n170 B.n169 10.6151
R2205 B.n173 B.n170 10.6151
R2206 B.n174 B.n173 10.6151
R2207 B.n177 B.n174 10.6151
R2208 B.n178 B.n177 10.6151
R2209 B.n181 B.n178 10.6151
R2210 B.n182 B.n181 10.6151
R2211 B.n185 B.n182 10.6151
R2212 B.n186 B.n185 10.6151
R2213 B.n189 B.n186 10.6151
R2214 B.n190 B.n189 10.6151
R2215 B.n193 B.n190 10.6151
R2216 B.n194 B.n193 10.6151
R2217 B.n198 B.n197 10.6151
R2218 B.n201 B.n198 10.6151
R2219 B.n202 B.n201 10.6151
R2220 B.n205 B.n202 10.6151
R2221 B.n206 B.n205 10.6151
R2222 B.n209 B.n206 10.6151
R2223 B.n210 B.n209 10.6151
R2224 B.n213 B.n210 10.6151
R2225 B.n218 B.n215 10.6151
R2226 B.n219 B.n218 10.6151
R2227 B.n222 B.n219 10.6151
R2228 B.n223 B.n222 10.6151
R2229 B.n226 B.n223 10.6151
R2230 B.n227 B.n226 10.6151
R2231 B.n230 B.n227 10.6151
R2232 B.n231 B.n230 10.6151
R2233 B.n234 B.n231 10.6151
R2234 B.n235 B.n234 10.6151
R2235 B.n238 B.n235 10.6151
R2236 B.n239 B.n238 10.6151
R2237 B.n242 B.n239 10.6151
R2238 B.n243 B.n242 10.6151
R2239 B.n246 B.n243 10.6151
R2240 B.n247 B.n246 10.6151
R2241 B.n250 B.n247 10.6151
R2242 B.n251 B.n250 10.6151
R2243 B.n254 B.n251 10.6151
R2244 B.n255 B.n254 10.6151
R2245 B.n258 B.n255 10.6151
R2246 B.n259 B.n258 10.6151
R2247 B.n262 B.n259 10.6151
R2248 B.n263 B.n262 10.6151
R2249 B.n266 B.n263 10.6151
R2250 B.n267 B.n266 10.6151
R2251 B.n270 B.n267 10.6151
R2252 B.n271 B.n270 10.6151
R2253 B.n274 B.n271 10.6151
R2254 B.n275 B.n274 10.6151
R2255 B.n278 B.n275 10.6151
R2256 B.n279 B.n278 10.6151
R2257 B.n282 B.n279 10.6151
R2258 B.n283 B.n282 10.6151
R2259 B.n286 B.n283 10.6151
R2260 B.n287 B.n286 10.6151
R2261 B.n290 B.n287 10.6151
R2262 B.n291 B.n290 10.6151
R2263 B.n294 B.n291 10.6151
R2264 B.n295 B.n294 10.6151
R2265 B.n736 B.n295 10.6151
R2266 B.n807 B.n0 8.11757
R2267 B.n807 B.n1 8.11757
R2268 B.n488 B.n385 6.5566
R2269 B.n381 B.n380 6.5566
R2270 B.n197 B.n113 6.5566
R2271 B.n214 B.n213 6.5566
R2272 B.n489 B.n488 4.05904
R2273 B.n511 B.n380 4.05904
R2274 B.n194 B.n113 4.05904
R2275 B.n215 B.n214 4.05904
R2276 VN.n5 VN.t1 245.733
R2277 VN.n25 VN.t4 245.733
R2278 VN.n4 VN.t6 216.541
R2279 VN.n10 VN.t3 216.541
R2280 VN.n17 VN.t2 216.541
R2281 VN.n24 VN.t5 216.541
R2282 VN.n22 VN.t7 216.541
R2283 VN.n36 VN.t0 216.541
R2284 VN.n18 VN.n17 173.351
R2285 VN.n37 VN.n36 173.351
R2286 VN.n35 VN.n19 161.3
R2287 VN.n34 VN.n33 161.3
R2288 VN.n32 VN.n20 161.3
R2289 VN.n31 VN.n30 161.3
R2290 VN.n29 VN.n21 161.3
R2291 VN.n28 VN.n27 161.3
R2292 VN.n26 VN.n23 161.3
R2293 VN.n16 VN.n0 161.3
R2294 VN.n15 VN.n14 161.3
R2295 VN.n13 VN.n1 161.3
R2296 VN.n12 VN.n11 161.3
R2297 VN.n9 VN.n2 161.3
R2298 VN.n8 VN.n7 161.3
R2299 VN.n6 VN.n3 161.3
R2300 VN.n5 VN.n4 61.2741
R2301 VN.n25 VN.n24 61.2741
R2302 VN.n9 VN.n8 56.5617
R2303 VN.n29 VN.n28 56.5617
R2304 VN.n15 VN.n1 48.3272
R2305 VN.n34 VN.n20 48.3272
R2306 VN VN.n37 45.3357
R2307 VN.n16 VN.n15 32.8269
R2308 VN.n35 VN.n34 32.8269
R2309 VN.n26 VN.n25 27.186
R2310 VN.n6 VN.n5 27.186
R2311 VN.n8 VN.n3 24.5923
R2312 VN.n11 VN.n9 24.5923
R2313 VN.n28 VN.n23 24.5923
R2314 VN.n30 VN.n29 24.5923
R2315 VN.n10 VN.n1 20.4117
R2316 VN.n22 VN.n20 20.4117
R2317 VN.n17 VN.n16 12.5423
R2318 VN.n36 VN.n35 12.5423
R2319 VN.n4 VN.n3 4.18111
R2320 VN.n11 VN.n10 4.18111
R2321 VN.n24 VN.n23 4.18111
R2322 VN.n30 VN.n22 4.18111
R2323 VN.n37 VN.n19 0.189894
R2324 VN.n33 VN.n19 0.189894
R2325 VN.n33 VN.n32 0.189894
R2326 VN.n32 VN.n31 0.189894
R2327 VN.n31 VN.n21 0.189894
R2328 VN.n27 VN.n21 0.189894
R2329 VN.n27 VN.n26 0.189894
R2330 VN.n7 VN.n6 0.189894
R2331 VN.n7 VN.n2 0.189894
R2332 VN.n12 VN.n2 0.189894
R2333 VN.n13 VN.n12 0.189894
R2334 VN.n14 VN.n13 0.189894
R2335 VN.n14 VN.n0 0.189894
R2336 VN.n18 VN.n0 0.189894
R2337 VN VN.n18 0.0516364
R2338 VDD2.n2 VDD2.n1 60.9927
R2339 VDD2.n2 VDD2.n0 60.9927
R2340 VDD2 VDD2.n5 60.9899
R2341 VDD2.n4 VDD2.n3 60.3284
R2342 VDD2.n4 VDD2.n2 40.5731
R2343 VDD2.n5 VDD2.t2 1.64502
R2344 VDD2.n5 VDD2.t3 1.64502
R2345 VDD2.n3 VDD2.t7 1.64502
R2346 VDD2.n3 VDD2.t0 1.64502
R2347 VDD2.n1 VDD2.t4 1.64502
R2348 VDD2.n1 VDD2.t5 1.64502
R2349 VDD2.n0 VDD2.t6 1.64502
R2350 VDD2.n0 VDD2.t1 1.64502
R2351 VDD2 VDD2.n4 0.778517
C0 VN VP 6.12554f
C1 VDD1 VDD2 1.14581f
C2 VTAIL VDD1 8.728661f
C3 VDD2 VP 0.385672f
C4 VTAIL VP 7.31169f
C5 VN VDD2 7.31369f
C6 VN VTAIL 7.29758f
C7 VTAIL VDD2 8.774631f
C8 VDD1 VP 7.54907f
C9 VN VDD1 0.149528f
C10 VDD2 B 4.111149f
C11 VDD1 B 4.410226f
C12 VTAIL B 9.54366f
C13 VN B 10.797339f
C14 VP B 9.137655f
C15 VDD2.t6 B 0.239943f
C16 VDD2.t1 B 0.239943f
C17 VDD2.n0 B 2.14079f
C18 VDD2.t4 B 0.239943f
C19 VDD2.t5 B 0.239943f
C20 VDD2.n1 B 2.14079f
C21 VDD2.n2 B 2.57638f
C22 VDD2.t7 B 0.239943f
C23 VDD2.t0 B 0.239943f
C24 VDD2.n3 B 2.13652f
C25 VDD2.n4 B 2.54081f
C26 VDD2.t2 B 0.239943f
C27 VDD2.t3 B 0.239943f
C28 VDD2.n5 B 2.14076f
C29 VN.n0 B 0.032785f
C30 VN.t2 B 1.44128f
C31 VN.n1 B 0.055989f
C32 VN.n2 B 0.032785f
C33 VN.n3 B 0.035885f
C34 VN.t1 B 1.5162f
C35 VN.t6 B 1.44128f
C36 VN.n4 B 0.569216f
C37 VN.n5 B 0.603947f
C38 VN.n6 B 0.173954f
C39 VN.n7 B 0.032785f
C40 VN.n8 B 0.047658f
C41 VN.n9 B 0.047658f
C42 VN.t3 B 1.44128f
C43 VN.n10 B 0.52412f
C44 VN.n11 B 0.035885f
C45 VN.n12 B 0.032785f
C46 VN.n13 B 0.032785f
C47 VN.n14 B 0.032785f
C48 VN.n15 B 0.029255f
C49 VN.n16 B 0.051058f
C50 VN.n17 B 0.585996f
C51 VN.n18 B 0.030029f
C52 VN.n19 B 0.032785f
C53 VN.t0 B 1.44128f
C54 VN.n20 B 0.055989f
C55 VN.n21 B 0.032785f
C56 VN.t7 B 1.44128f
C57 VN.n22 B 0.52412f
C58 VN.n23 B 0.035885f
C59 VN.t4 B 1.5162f
C60 VN.t5 B 1.44128f
C61 VN.n24 B 0.569216f
C62 VN.n25 B 0.603947f
C63 VN.n26 B 0.173954f
C64 VN.n27 B 0.032785f
C65 VN.n28 B 0.047658f
C66 VN.n29 B 0.047658f
C67 VN.n30 B 0.035885f
C68 VN.n31 B 0.032785f
C69 VN.n32 B 0.032785f
C70 VN.n33 B 0.032785f
C71 VN.n34 B 0.029255f
C72 VN.n35 B 0.051058f
C73 VN.n36 B 0.585996f
C74 VN.n37 B 1.53788f
C75 VTAIL.t6 B 0.182745f
C76 VTAIL.t4 B 0.182745f
C77 VTAIL.n0 B 1.56727f
C78 VTAIL.n1 B 0.28705f
C79 VTAIL.n2 B 0.025961f
C80 VTAIL.n3 B 0.019207f
C81 VTAIL.n4 B 0.010321f
C82 VTAIL.n5 B 0.024395f
C83 VTAIL.n6 B 0.010928f
C84 VTAIL.n7 B 0.019207f
C85 VTAIL.n8 B 0.010321f
C86 VTAIL.n9 B 0.024395f
C87 VTAIL.n10 B 0.010928f
C88 VTAIL.n11 B 0.019207f
C89 VTAIL.n12 B 0.010625f
C90 VTAIL.n13 B 0.024395f
C91 VTAIL.n14 B 0.010928f
C92 VTAIL.n15 B 0.019207f
C93 VTAIL.n16 B 0.010321f
C94 VTAIL.n17 B 0.024395f
C95 VTAIL.n18 B 0.010928f
C96 VTAIL.n19 B 0.019207f
C97 VTAIL.n20 B 0.010321f
C98 VTAIL.n21 B 0.018297f
C99 VTAIL.n22 B 0.017246f
C100 VTAIL.t5 B 0.041207f
C101 VTAIL.n23 B 0.138777f
C102 VTAIL.n24 B 0.972392f
C103 VTAIL.n25 B 0.010321f
C104 VTAIL.n26 B 0.010928f
C105 VTAIL.n27 B 0.024395f
C106 VTAIL.n28 B 0.024395f
C107 VTAIL.n29 B 0.010928f
C108 VTAIL.n30 B 0.010321f
C109 VTAIL.n31 B 0.019207f
C110 VTAIL.n32 B 0.019207f
C111 VTAIL.n33 B 0.010321f
C112 VTAIL.n34 B 0.010928f
C113 VTAIL.n35 B 0.024395f
C114 VTAIL.n36 B 0.024395f
C115 VTAIL.n37 B 0.010928f
C116 VTAIL.n38 B 0.010321f
C117 VTAIL.n39 B 0.019207f
C118 VTAIL.n40 B 0.019207f
C119 VTAIL.n41 B 0.010321f
C120 VTAIL.n42 B 0.010321f
C121 VTAIL.n43 B 0.010928f
C122 VTAIL.n44 B 0.024395f
C123 VTAIL.n45 B 0.024395f
C124 VTAIL.n46 B 0.024395f
C125 VTAIL.n47 B 0.010625f
C126 VTAIL.n48 B 0.010321f
C127 VTAIL.n49 B 0.019207f
C128 VTAIL.n50 B 0.019207f
C129 VTAIL.n51 B 0.010321f
C130 VTAIL.n52 B 0.010928f
C131 VTAIL.n53 B 0.024395f
C132 VTAIL.n54 B 0.024395f
C133 VTAIL.n55 B 0.010928f
C134 VTAIL.n56 B 0.010321f
C135 VTAIL.n57 B 0.019207f
C136 VTAIL.n58 B 0.019207f
C137 VTAIL.n59 B 0.010321f
C138 VTAIL.n60 B 0.010928f
C139 VTAIL.n61 B 0.024395f
C140 VTAIL.n62 B 0.050979f
C141 VTAIL.n63 B 0.010928f
C142 VTAIL.n64 B 0.010321f
C143 VTAIL.n65 B 0.042298f
C144 VTAIL.n66 B 0.02827f
C145 VTAIL.n67 B 0.133399f
C146 VTAIL.n68 B 0.025961f
C147 VTAIL.n69 B 0.019207f
C148 VTAIL.n70 B 0.010321f
C149 VTAIL.n71 B 0.024395f
C150 VTAIL.n72 B 0.010928f
C151 VTAIL.n73 B 0.019207f
C152 VTAIL.n74 B 0.010321f
C153 VTAIL.n75 B 0.024395f
C154 VTAIL.n76 B 0.010928f
C155 VTAIL.n77 B 0.019207f
C156 VTAIL.n78 B 0.010625f
C157 VTAIL.n79 B 0.024395f
C158 VTAIL.n80 B 0.010928f
C159 VTAIL.n81 B 0.019207f
C160 VTAIL.n82 B 0.010321f
C161 VTAIL.n83 B 0.024395f
C162 VTAIL.n84 B 0.010928f
C163 VTAIL.n85 B 0.019207f
C164 VTAIL.n86 B 0.010321f
C165 VTAIL.n87 B 0.018297f
C166 VTAIL.n88 B 0.017246f
C167 VTAIL.t9 B 0.041207f
C168 VTAIL.n89 B 0.138777f
C169 VTAIL.n90 B 0.972392f
C170 VTAIL.n91 B 0.010321f
C171 VTAIL.n92 B 0.010928f
C172 VTAIL.n93 B 0.024395f
C173 VTAIL.n94 B 0.024395f
C174 VTAIL.n95 B 0.010928f
C175 VTAIL.n96 B 0.010321f
C176 VTAIL.n97 B 0.019207f
C177 VTAIL.n98 B 0.019207f
C178 VTAIL.n99 B 0.010321f
C179 VTAIL.n100 B 0.010928f
C180 VTAIL.n101 B 0.024395f
C181 VTAIL.n102 B 0.024395f
C182 VTAIL.n103 B 0.010928f
C183 VTAIL.n104 B 0.010321f
C184 VTAIL.n105 B 0.019207f
C185 VTAIL.n106 B 0.019207f
C186 VTAIL.n107 B 0.010321f
C187 VTAIL.n108 B 0.010321f
C188 VTAIL.n109 B 0.010928f
C189 VTAIL.n110 B 0.024395f
C190 VTAIL.n111 B 0.024395f
C191 VTAIL.n112 B 0.024395f
C192 VTAIL.n113 B 0.010625f
C193 VTAIL.n114 B 0.010321f
C194 VTAIL.n115 B 0.019207f
C195 VTAIL.n116 B 0.019207f
C196 VTAIL.n117 B 0.010321f
C197 VTAIL.n118 B 0.010928f
C198 VTAIL.n119 B 0.024395f
C199 VTAIL.n120 B 0.024395f
C200 VTAIL.n121 B 0.010928f
C201 VTAIL.n122 B 0.010321f
C202 VTAIL.n123 B 0.019207f
C203 VTAIL.n124 B 0.019207f
C204 VTAIL.n125 B 0.010321f
C205 VTAIL.n126 B 0.010928f
C206 VTAIL.n127 B 0.024395f
C207 VTAIL.n128 B 0.050979f
C208 VTAIL.n129 B 0.010928f
C209 VTAIL.n130 B 0.010321f
C210 VTAIL.n131 B 0.042298f
C211 VTAIL.n132 B 0.02827f
C212 VTAIL.n133 B 0.133399f
C213 VTAIL.t11 B 0.182745f
C214 VTAIL.t10 B 0.182745f
C215 VTAIL.n134 B 1.56727f
C216 VTAIL.n135 B 0.372549f
C217 VTAIL.n136 B 0.025961f
C218 VTAIL.n137 B 0.019207f
C219 VTAIL.n138 B 0.010321f
C220 VTAIL.n139 B 0.024395f
C221 VTAIL.n140 B 0.010928f
C222 VTAIL.n141 B 0.019207f
C223 VTAIL.n142 B 0.010321f
C224 VTAIL.n143 B 0.024395f
C225 VTAIL.n144 B 0.010928f
C226 VTAIL.n145 B 0.019207f
C227 VTAIL.n146 B 0.010625f
C228 VTAIL.n147 B 0.024395f
C229 VTAIL.n148 B 0.010928f
C230 VTAIL.n149 B 0.019207f
C231 VTAIL.n150 B 0.010321f
C232 VTAIL.n151 B 0.024395f
C233 VTAIL.n152 B 0.010928f
C234 VTAIL.n153 B 0.019207f
C235 VTAIL.n154 B 0.010321f
C236 VTAIL.n155 B 0.018297f
C237 VTAIL.n156 B 0.017246f
C238 VTAIL.t8 B 0.041207f
C239 VTAIL.n157 B 0.138777f
C240 VTAIL.n158 B 0.972392f
C241 VTAIL.n159 B 0.010321f
C242 VTAIL.n160 B 0.010928f
C243 VTAIL.n161 B 0.024395f
C244 VTAIL.n162 B 0.024395f
C245 VTAIL.n163 B 0.010928f
C246 VTAIL.n164 B 0.010321f
C247 VTAIL.n165 B 0.019207f
C248 VTAIL.n166 B 0.019207f
C249 VTAIL.n167 B 0.010321f
C250 VTAIL.n168 B 0.010928f
C251 VTAIL.n169 B 0.024395f
C252 VTAIL.n170 B 0.024395f
C253 VTAIL.n171 B 0.010928f
C254 VTAIL.n172 B 0.010321f
C255 VTAIL.n173 B 0.019207f
C256 VTAIL.n174 B 0.019207f
C257 VTAIL.n175 B 0.010321f
C258 VTAIL.n176 B 0.010321f
C259 VTAIL.n177 B 0.010928f
C260 VTAIL.n178 B 0.024395f
C261 VTAIL.n179 B 0.024395f
C262 VTAIL.n180 B 0.024395f
C263 VTAIL.n181 B 0.010625f
C264 VTAIL.n182 B 0.010321f
C265 VTAIL.n183 B 0.019207f
C266 VTAIL.n184 B 0.019207f
C267 VTAIL.n185 B 0.010321f
C268 VTAIL.n186 B 0.010928f
C269 VTAIL.n187 B 0.024395f
C270 VTAIL.n188 B 0.024395f
C271 VTAIL.n189 B 0.010928f
C272 VTAIL.n190 B 0.010321f
C273 VTAIL.n191 B 0.019207f
C274 VTAIL.n192 B 0.019207f
C275 VTAIL.n193 B 0.010321f
C276 VTAIL.n194 B 0.010928f
C277 VTAIL.n195 B 0.024395f
C278 VTAIL.n196 B 0.050979f
C279 VTAIL.n197 B 0.010928f
C280 VTAIL.n198 B 0.010321f
C281 VTAIL.n199 B 0.042298f
C282 VTAIL.n200 B 0.02827f
C283 VTAIL.n201 B 1.09671f
C284 VTAIL.n202 B 0.025961f
C285 VTAIL.n203 B 0.019207f
C286 VTAIL.n204 B 0.010321f
C287 VTAIL.n205 B 0.024395f
C288 VTAIL.n206 B 0.010928f
C289 VTAIL.n207 B 0.019207f
C290 VTAIL.n208 B 0.010321f
C291 VTAIL.n209 B 0.024395f
C292 VTAIL.n210 B 0.010928f
C293 VTAIL.n211 B 0.019207f
C294 VTAIL.n212 B 0.010625f
C295 VTAIL.n213 B 0.024395f
C296 VTAIL.n214 B 0.010321f
C297 VTAIL.n215 B 0.010928f
C298 VTAIL.n216 B 0.019207f
C299 VTAIL.n217 B 0.010321f
C300 VTAIL.n218 B 0.024395f
C301 VTAIL.n219 B 0.010928f
C302 VTAIL.n220 B 0.019207f
C303 VTAIL.n221 B 0.010321f
C304 VTAIL.n222 B 0.018297f
C305 VTAIL.n223 B 0.017246f
C306 VTAIL.t7 B 0.041207f
C307 VTAIL.n224 B 0.138777f
C308 VTAIL.n225 B 0.972392f
C309 VTAIL.n226 B 0.010321f
C310 VTAIL.n227 B 0.010928f
C311 VTAIL.n228 B 0.024395f
C312 VTAIL.n229 B 0.024395f
C313 VTAIL.n230 B 0.010928f
C314 VTAIL.n231 B 0.010321f
C315 VTAIL.n232 B 0.019207f
C316 VTAIL.n233 B 0.019207f
C317 VTAIL.n234 B 0.010321f
C318 VTAIL.n235 B 0.010928f
C319 VTAIL.n236 B 0.024395f
C320 VTAIL.n237 B 0.024395f
C321 VTAIL.n238 B 0.010928f
C322 VTAIL.n239 B 0.010321f
C323 VTAIL.n240 B 0.019207f
C324 VTAIL.n241 B 0.019207f
C325 VTAIL.n242 B 0.010321f
C326 VTAIL.n243 B 0.010928f
C327 VTAIL.n244 B 0.024395f
C328 VTAIL.n245 B 0.024395f
C329 VTAIL.n246 B 0.024395f
C330 VTAIL.n247 B 0.010625f
C331 VTAIL.n248 B 0.010321f
C332 VTAIL.n249 B 0.019207f
C333 VTAIL.n250 B 0.019207f
C334 VTAIL.n251 B 0.010321f
C335 VTAIL.n252 B 0.010928f
C336 VTAIL.n253 B 0.024395f
C337 VTAIL.n254 B 0.024395f
C338 VTAIL.n255 B 0.010928f
C339 VTAIL.n256 B 0.010321f
C340 VTAIL.n257 B 0.019207f
C341 VTAIL.n258 B 0.019207f
C342 VTAIL.n259 B 0.010321f
C343 VTAIL.n260 B 0.010928f
C344 VTAIL.n261 B 0.024395f
C345 VTAIL.n262 B 0.050979f
C346 VTAIL.n263 B 0.010928f
C347 VTAIL.n264 B 0.010321f
C348 VTAIL.n265 B 0.042298f
C349 VTAIL.n266 B 0.02827f
C350 VTAIL.n267 B 1.09671f
C351 VTAIL.t1 B 0.182745f
C352 VTAIL.t0 B 0.182745f
C353 VTAIL.n268 B 1.56728f
C354 VTAIL.n269 B 0.37254f
C355 VTAIL.n270 B 0.025961f
C356 VTAIL.n271 B 0.019207f
C357 VTAIL.n272 B 0.010321f
C358 VTAIL.n273 B 0.024395f
C359 VTAIL.n274 B 0.010928f
C360 VTAIL.n275 B 0.019207f
C361 VTAIL.n276 B 0.010321f
C362 VTAIL.n277 B 0.024395f
C363 VTAIL.n278 B 0.010928f
C364 VTAIL.n279 B 0.019207f
C365 VTAIL.n280 B 0.010625f
C366 VTAIL.n281 B 0.024395f
C367 VTAIL.n282 B 0.010321f
C368 VTAIL.n283 B 0.010928f
C369 VTAIL.n284 B 0.019207f
C370 VTAIL.n285 B 0.010321f
C371 VTAIL.n286 B 0.024395f
C372 VTAIL.n287 B 0.010928f
C373 VTAIL.n288 B 0.019207f
C374 VTAIL.n289 B 0.010321f
C375 VTAIL.n290 B 0.018297f
C376 VTAIL.n291 B 0.017246f
C377 VTAIL.t3 B 0.041207f
C378 VTAIL.n292 B 0.138777f
C379 VTAIL.n293 B 0.972392f
C380 VTAIL.n294 B 0.010321f
C381 VTAIL.n295 B 0.010928f
C382 VTAIL.n296 B 0.024395f
C383 VTAIL.n297 B 0.024395f
C384 VTAIL.n298 B 0.010928f
C385 VTAIL.n299 B 0.010321f
C386 VTAIL.n300 B 0.019207f
C387 VTAIL.n301 B 0.019207f
C388 VTAIL.n302 B 0.010321f
C389 VTAIL.n303 B 0.010928f
C390 VTAIL.n304 B 0.024395f
C391 VTAIL.n305 B 0.024395f
C392 VTAIL.n306 B 0.010928f
C393 VTAIL.n307 B 0.010321f
C394 VTAIL.n308 B 0.019207f
C395 VTAIL.n309 B 0.019207f
C396 VTAIL.n310 B 0.010321f
C397 VTAIL.n311 B 0.010928f
C398 VTAIL.n312 B 0.024395f
C399 VTAIL.n313 B 0.024395f
C400 VTAIL.n314 B 0.024395f
C401 VTAIL.n315 B 0.010625f
C402 VTAIL.n316 B 0.010321f
C403 VTAIL.n317 B 0.019207f
C404 VTAIL.n318 B 0.019207f
C405 VTAIL.n319 B 0.010321f
C406 VTAIL.n320 B 0.010928f
C407 VTAIL.n321 B 0.024395f
C408 VTAIL.n322 B 0.024395f
C409 VTAIL.n323 B 0.010928f
C410 VTAIL.n324 B 0.010321f
C411 VTAIL.n325 B 0.019207f
C412 VTAIL.n326 B 0.019207f
C413 VTAIL.n327 B 0.010321f
C414 VTAIL.n328 B 0.010928f
C415 VTAIL.n329 B 0.024395f
C416 VTAIL.n330 B 0.050979f
C417 VTAIL.n331 B 0.010928f
C418 VTAIL.n332 B 0.010321f
C419 VTAIL.n333 B 0.042298f
C420 VTAIL.n334 B 0.02827f
C421 VTAIL.n335 B 0.133399f
C422 VTAIL.n336 B 0.025961f
C423 VTAIL.n337 B 0.019207f
C424 VTAIL.n338 B 0.010321f
C425 VTAIL.n339 B 0.024395f
C426 VTAIL.n340 B 0.010928f
C427 VTAIL.n341 B 0.019207f
C428 VTAIL.n342 B 0.010321f
C429 VTAIL.n343 B 0.024395f
C430 VTAIL.n344 B 0.010928f
C431 VTAIL.n345 B 0.019207f
C432 VTAIL.n346 B 0.010625f
C433 VTAIL.n347 B 0.024395f
C434 VTAIL.n348 B 0.010321f
C435 VTAIL.n349 B 0.010928f
C436 VTAIL.n350 B 0.019207f
C437 VTAIL.n351 B 0.010321f
C438 VTAIL.n352 B 0.024395f
C439 VTAIL.n353 B 0.010928f
C440 VTAIL.n354 B 0.019207f
C441 VTAIL.n355 B 0.010321f
C442 VTAIL.n356 B 0.018297f
C443 VTAIL.n357 B 0.017246f
C444 VTAIL.t13 B 0.041207f
C445 VTAIL.n358 B 0.138777f
C446 VTAIL.n359 B 0.972392f
C447 VTAIL.n360 B 0.010321f
C448 VTAIL.n361 B 0.010928f
C449 VTAIL.n362 B 0.024395f
C450 VTAIL.n363 B 0.024395f
C451 VTAIL.n364 B 0.010928f
C452 VTAIL.n365 B 0.010321f
C453 VTAIL.n366 B 0.019207f
C454 VTAIL.n367 B 0.019207f
C455 VTAIL.n368 B 0.010321f
C456 VTAIL.n369 B 0.010928f
C457 VTAIL.n370 B 0.024395f
C458 VTAIL.n371 B 0.024395f
C459 VTAIL.n372 B 0.010928f
C460 VTAIL.n373 B 0.010321f
C461 VTAIL.n374 B 0.019207f
C462 VTAIL.n375 B 0.019207f
C463 VTAIL.n376 B 0.010321f
C464 VTAIL.n377 B 0.010928f
C465 VTAIL.n378 B 0.024395f
C466 VTAIL.n379 B 0.024395f
C467 VTAIL.n380 B 0.024395f
C468 VTAIL.n381 B 0.010625f
C469 VTAIL.n382 B 0.010321f
C470 VTAIL.n383 B 0.019207f
C471 VTAIL.n384 B 0.019207f
C472 VTAIL.n385 B 0.010321f
C473 VTAIL.n386 B 0.010928f
C474 VTAIL.n387 B 0.024395f
C475 VTAIL.n388 B 0.024395f
C476 VTAIL.n389 B 0.010928f
C477 VTAIL.n390 B 0.010321f
C478 VTAIL.n391 B 0.019207f
C479 VTAIL.n392 B 0.019207f
C480 VTAIL.n393 B 0.010321f
C481 VTAIL.n394 B 0.010928f
C482 VTAIL.n395 B 0.024395f
C483 VTAIL.n396 B 0.050979f
C484 VTAIL.n397 B 0.010928f
C485 VTAIL.n398 B 0.010321f
C486 VTAIL.n399 B 0.042298f
C487 VTAIL.n400 B 0.02827f
C488 VTAIL.n401 B 0.133399f
C489 VTAIL.t14 B 0.182745f
C490 VTAIL.t15 B 0.182745f
C491 VTAIL.n402 B 1.56728f
C492 VTAIL.n403 B 0.37254f
C493 VTAIL.n404 B 0.025961f
C494 VTAIL.n405 B 0.019207f
C495 VTAIL.n406 B 0.010321f
C496 VTAIL.n407 B 0.024395f
C497 VTAIL.n408 B 0.010928f
C498 VTAIL.n409 B 0.019207f
C499 VTAIL.n410 B 0.010321f
C500 VTAIL.n411 B 0.024395f
C501 VTAIL.n412 B 0.010928f
C502 VTAIL.n413 B 0.019207f
C503 VTAIL.n414 B 0.010625f
C504 VTAIL.n415 B 0.024395f
C505 VTAIL.n416 B 0.010321f
C506 VTAIL.n417 B 0.010928f
C507 VTAIL.n418 B 0.019207f
C508 VTAIL.n419 B 0.010321f
C509 VTAIL.n420 B 0.024395f
C510 VTAIL.n421 B 0.010928f
C511 VTAIL.n422 B 0.019207f
C512 VTAIL.n423 B 0.010321f
C513 VTAIL.n424 B 0.018297f
C514 VTAIL.n425 B 0.017246f
C515 VTAIL.t12 B 0.041207f
C516 VTAIL.n426 B 0.138777f
C517 VTAIL.n427 B 0.972392f
C518 VTAIL.n428 B 0.010321f
C519 VTAIL.n429 B 0.010928f
C520 VTAIL.n430 B 0.024395f
C521 VTAIL.n431 B 0.024395f
C522 VTAIL.n432 B 0.010928f
C523 VTAIL.n433 B 0.010321f
C524 VTAIL.n434 B 0.019207f
C525 VTAIL.n435 B 0.019207f
C526 VTAIL.n436 B 0.010321f
C527 VTAIL.n437 B 0.010928f
C528 VTAIL.n438 B 0.024395f
C529 VTAIL.n439 B 0.024395f
C530 VTAIL.n440 B 0.010928f
C531 VTAIL.n441 B 0.010321f
C532 VTAIL.n442 B 0.019207f
C533 VTAIL.n443 B 0.019207f
C534 VTAIL.n444 B 0.010321f
C535 VTAIL.n445 B 0.010928f
C536 VTAIL.n446 B 0.024395f
C537 VTAIL.n447 B 0.024395f
C538 VTAIL.n448 B 0.024395f
C539 VTAIL.n449 B 0.010625f
C540 VTAIL.n450 B 0.010321f
C541 VTAIL.n451 B 0.019207f
C542 VTAIL.n452 B 0.019207f
C543 VTAIL.n453 B 0.010321f
C544 VTAIL.n454 B 0.010928f
C545 VTAIL.n455 B 0.024395f
C546 VTAIL.n456 B 0.024395f
C547 VTAIL.n457 B 0.010928f
C548 VTAIL.n458 B 0.010321f
C549 VTAIL.n459 B 0.019207f
C550 VTAIL.n460 B 0.019207f
C551 VTAIL.n461 B 0.010321f
C552 VTAIL.n462 B 0.010928f
C553 VTAIL.n463 B 0.024395f
C554 VTAIL.n464 B 0.050979f
C555 VTAIL.n465 B 0.010928f
C556 VTAIL.n466 B 0.010321f
C557 VTAIL.n467 B 0.042298f
C558 VTAIL.n468 B 0.02827f
C559 VTAIL.n469 B 1.09671f
C560 VTAIL.n470 B 0.025961f
C561 VTAIL.n471 B 0.019207f
C562 VTAIL.n472 B 0.010321f
C563 VTAIL.n473 B 0.024395f
C564 VTAIL.n474 B 0.010928f
C565 VTAIL.n475 B 0.019207f
C566 VTAIL.n476 B 0.010321f
C567 VTAIL.n477 B 0.024395f
C568 VTAIL.n478 B 0.010928f
C569 VTAIL.n479 B 0.019207f
C570 VTAIL.n480 B 0.010625f
C571 VTAIL.n481 B 0.024395f
C572 VTAIL.n482 B 0.010928f
C573 VTAIL.n483 B 0.019207f
C574 VTAIL.n484 B 0.010321f
C575 VTAIL.n485 B 0.024395f
C576 VTAIL.n486 B 0.010928f
C577 VTAIL.n487 B 0.019207f
C578 VTAIL.n488 B 0.010321f
C579 VTAIL.n489 B 0.018297f
C580 VTAIL.n490 B 0.017246f
C581 VTAIL.t2 B 0.041207f
C582 VTAIL.n491 B 0.138777f
C583 VTAIL.n492 B 0.972392f
C584 VTAIL.n493 B 0.010321f
C585 VTAIL.n494 B 0.010928f
C586 VTAIL.n495 B 0.024395f
C587 VTAIL.n496 B 0.024395f
C588 VTAIL.n497 B 0.010928f
C589 VTAIL.n498 B 0.010321f
C590 VTAIL.n499 B 0.019207f
C591 VTAIL.n500 B 0.019207f
C592 VTAIL.n501 B 0.010321f
C593 VTAIL.n502 B 0.010928f
C594 VTAIL.n503 B 0.024395f
C595 VTAIL.n504 B 0.024395f
C596 VTAIL.n505 B 0.010928f
C597 VTAIL.n506 B 0.010321f
C598 VTAIL.n507 B 0.019207f
C599 VTAIL.n508 B 0.019207f
C600 VTAIL.n509 B 0.010321f
C601 VTAIL.n510 B 0.010321f
C602 VTAIL.n511 B 0.010928f
C603 VTAIL.n512 B 0.024395f
C604 VTAIL.n513 B 0.024395f
C605 VTAIL.n514 B 0.024395f
C606 VTAIL.n515 B 0.010625f
C607 VTAIL.n516 B 0.010321f
C608 VTAIL.n517 B 0.019207f
C609 VTAIL.n518 B 0.019207f
C610 VTAIL.n519 B 0.010321f
C611 VTAIL.n520 B 0.010928f
C612 VTAIL.n521 B 0.024395f
C613 VTAIL.n522 B 0.024395f
C614 VTAIL.n523 B 0.010928f
C615 VTAIL.n524 B 0.010321f
C616 VTAIL.n525 B 0.019207f
C617 VTAIL.n526 B 0.019207f
C618 VTAIL.n527 B 0.010321f
C619 VTAIL.n528 B 0.010928f
C620 VTAIL.n529 B 0.024395f
C621 VTAIL.n530 B 0.050979f
C622 VTAIL.n531 B 0.010928f
C623 VTAIL.n532 B 0.010321f
C624 VTAIL.n533 B 0.042298f
C625 VTAIL.n534 B 0.02827f
C626 VTAIL.n535 B 1.09311f
C627 VDD1.t0 B 0.240045f
C628 VDD1.t6 B 0.240045f
C629 VDD1.n0 B 2.14253f
C630 VDD1.t3 B 0.240045f
C631 VDD1.t4 B 0.240045f
C632 VDD1.n1 B 2.1417f
C633 VDD1.t2 B 0.240045f
C634 VDD1.t5 B 0.240045f
C635 VDD1.n2 B 2.1417f
C636 VDD1.n3 B 2.63082f
C637 VDD1.t7 B 0.240045f
C638 VDD1.t1 B 0.240045f
C639 VDD1.n4 B 2.13742f
C640 VDD1.n5 B 2.57226f
C641 VP.n0 B 0.033175f
C642 VP.t6 B 1.45845f
C643 VP.n1 B 0.056656f
C644 VP.n2 B 0.033175f
C645 VP.n3 B 0.036312f
C646 VP.n4 B 0.033175f
C647 VP.t7 B 1.45845f
C648 VP.n5 B 0.592978f
C649 VP.n6 B 0.033175f
C650 VP.t3 B 1.45845f
C651 VP.n7 B 0.056656f
C652 VP.n8 B 0.033175f
C653 VP.n9 B 0.036312f
C654 VP.t2 B 1.53427f
C655 VP.t1 B 1.45845f
C656 VP.n10 B 0.575998f
C657 VP.n11 B 0.611143f
C658 VP.n12 B 0.176026f
C659 VP.n13 B 0.033175f
C660 VP.n14 B 0.048225f
C661 VP.n15 B 0.048225f
C662 VP.t0 B 1.45845f
C663 VP.n16 B 0.530365f
C664 VP.n17 B 0.036312f
C665 VP.n18 B 0.033175f
C666 VP.n19 B 0.033175f
C667 VP.n20 B 0.033175f
C668 VP.n21 B 0.029604f
C669 VP.n22 B 0.051667f
C670 VP.n23 B 0.592978f
C671 VP.n24 B 1.53451f
C672 VP.n25 B 1.56111f
C673 VP.n26 B 0.033175f
C674 VP.n27 B 0.051667f
C675 VP.n28 B 0.029604f
C676 VP.t4 B 1.45845f
C677 VP.n29 B 0.530365f
C678 VP.n30 B 0.056656f
C679 VP.n31 B 0.033175f
C680 VP.n32 B 0.033175f
C681 VP.n33 B 0.033175f
C682 VP.n34 B 0.048225f
C683 VP.n35 B 0.048225f
C684 VP.t5 B 1.45845f
C685 VP.n36 B 0.530365f
C686 VP.n37 B 0.036312f
C687 VP.n38 B 0.033175f
C688 VP.n39 B 0.033175f
C689 VP.n40 B 0.033175f
C690 VP.n41 B 0.029604f
C691 VP.n42 B 0.051667f
C692 VP.n43 B 0.592978f
C693 VP.n44 B 0.030387f
.ends

