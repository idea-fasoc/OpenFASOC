* NGSPICE file created from diff_pair_sample_0588.ext - technology: sky130A

.subckt diff_pair_sample_0588 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X1 VDD1.t9 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=1.65495 ps=10.36 w=10.03 l=3.98
X2 VDD2.t5 VN.t1 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=3.9117 ps=20.84 w=10.03 l=3.98
X3 VDD1.t8 VP.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X4 VDD2.t7 VN.t2 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=1.65495 ps=10.36 w=10.03 l=3.98
X5 VDD1.t7 VP.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=3.9117 ps=20.84 w=10.03 l=3.98
X6 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X7 VTAIL.t15 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X8 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=0 ps=0 w=10.03 l=3.98
X9 VTAIL.t14 VN.t4 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X10 VDD2.t2 VN.t5 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=1.65495 ps=10.36 w=10.03 l=3.98
X11 VTAIL.t12 VN.t6 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X12 VDD1.t5 VP.t4 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=1.65495 ps=10.36 w=10.03 l=3.98
X13 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=0 ps=0 w=10.03 l=3.98
X14 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=0 ps=0 w=10.03 l=3.98
X15 VTAIL.t3 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X16 VDD2.t1 VN.t7 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X17 VTAIL.t0 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X18 VDD2.t9 VN.t8 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=3.9117 ps=20.84 w=10.03 l=3.98
X19 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.9117 pd=20.84 as=0 ps=0 w=10.03 l=3.98
X21 VTAIL.t8 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
X22 VDD1.t0 VP.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=3.9117 ps=20.84 w=10.03 l=3.98
X23 VDD2.t3 VN.t9 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.65495 pd=10.36 as=1.65495 ps=10.36 w=10.03 l=3.98
R0 VN.n113 VN.n58 161.3
R1 VN.n112 VN.n111 161.3
R2 VN.n110 VN.n59 161.3
R3 VN.n109 VN.n108 161.3
R4 VN.n107 VN.n60 161.3
R5 VN.n106 VN.n105 161.3
R6 VN.n104 VN.n61 161.3
R7 VN.n103 VN.n102 161.3
R8 VN.n100 VN.n62 161.3
R9 VN.n99 VN.n98 161.3
R10 VN.n97 VN.n63 161.3
R11 VN.n96 VN.n95 161.3
R12 VN.n94 VN.n64 161.3
R13 VN.n93 VN.n92 161.3
R14 VN.n91 VN.n65 161.3
R15 VN.n90 VN.n89 161.3
R16 VN.n88 VN.n66 161.3
R17 VN.n86 VN.n85 161.3
R18 VN.n84 VN.n67 161.3
R19 VN.n83 VN.n82 161.3
R20 VN.n81 VN.n68 161.3
R21 VN.n80 VN.n79 161.3
R22 VN.n78 VN.n69 161.3
R23 VN.n77 VN.n76 161.3
R24 VN.n75 VN.n70 161.3
R25 VN.n74 VN.n73 161.3
R26 VN.n55 VN.n0 161.3
R27 VN.n54 VN.n53 161.3
R28 VN.n52 VN.n1 161.3
R29 VN.n51 VN.n50 161.3
R30 VN.n49 VN.n2 161.3
R31 VN.n48 VN.n47 161.3
R32 VN.n46 VN.n3 161.3
R33 VN.n45 VN.n44 161.3
R34 VN.n42 VN.n4 161.3
R35 VN.n41 VN.n40 161.3
R36 VN.n39 VN.n5 161.3
R37 VN.n38 VN.n37 161.3
R38 VN.n36 VN.n6 161.3
R39 VN.n35 VN.n34 161.3
R40 VN.n33 VN.n7 161.3
R41 VN.n32 VN.n31 161.3
R42 VN.n30 VN.n8 161.3
R43 VN.n28 VN.n27 161.3
R44 VN.n26 VN.n9 161.3
R45 VN.n25 VN.n24 161.3
R46 VN.n23 VN.n10 161.3
R47 VN.n22 VN.n21 161.3
R48 VN.n20 VN.n11 161.3
R49 VN.n19 VN.n18 161.3
R50 VN.n17 VN.n12 161.3
R51 VN.n16 VN.n15 161.3
R52 VN.n14 VN.t2 93.0545
R53 VN.n72 VN.t8 93.0545
R54 VN.n14 VN.n13 72.0574
R55 VN.n72 VN.n71 72.0574
R56 VN.n57 VN.n56 64.0762
R57 VN.n115 VN.n114 64.0762
R58 VN.n13 VN.t6 60.7349
R59 VN.n29 VN.t7 60.7349
R60 VN.n43 VN.t0 60.7349
R61 VN.n56 VN.t1 60.7349
R62 VN.n71 VN.t4 60.7349
R63 VN.n87 VN.t9 60.7349
R64 VN.n101 VN.t3 60.7349
R65 VN.n114 VN.t5 60.7349
R66 VN VN.n115 59.3716
R67 VN.n50 VN.n49 56.5193
R68 VN.n108 VN.n107 56.5193
R69 VN.n23 VN.n22 49.7204
R70 VN.n36 VN.n35 49.7204
R71 VN.n81 VN.n80 49.7204
R72 VN.n94 VN.n93 49.7204
R73 VN.n22 VN.n11 31.2664
R74 VN.n37 VN.n36 31.2664
R75 VN.n80 VN.n69 31.2664
R76 VN.n95 VN.n94 31.2664
R77 VN.n17 VN.n16 24.4675
R78 VN.n18 VN.n17 24.4675
R79 VN.n18 VN.n11 24.4675
R80 VN.n24 VN.n23 24.4675
R81 VN.n24 VN.n9 24.4675
R82 VN.n28 VN.n9 24.4675
R83 VN.n31 VN.n30 24.4675
R84 VN.n31 VN.n7 24.4675
R85 VN.n35 VN.n7 24.4675
R86 VN.n37 VN.n5 24.4675
R87 VN.n41 VN.n5 24.4675
R88 VN.n42 VN.n41 24.4675
R89 VN.n44 VN.n3 24.4675
R90 VN.n48 VN.n3 24.4675
R91 VN.n49 VN.n48 24.4675
R92 VN.n50 VN.n1 24.4675
R93 VN.n54 VN.n1 24.4675
R94 VN.n55 VN.n54 24.4675
R95 VN.n76 VN.n69 24.4675
R96 VN.n76 VN.n75 24.4675
R97 VN.n75 VN.n74 24.4675
R98 VN.n93 VN.n65 24.4675
R99 VN.n89 VN.n65 24.4675
R100 VN.n89 VN.n88 24.4675
R101 VN.n86 VN.n67 24.4675
R102 VN.n82 VN.n67 24.4675
R103 VN.n82 VN.n81 24.4675
R104 VN.n107 VN.n106 24.4675
R105 VN.n106 VN.n61 24.4675
R106 VN.n102 VN.n61 24.4675
R107 VN.n100 VN.n99 24.4675
R108 VN.n99 VN.n63 24.4675
R109 VN.n95 VN.n63 24.4675
R110 VN.n113 VN.n112 24.4675
R111 VN.n112 VN.n59 24.4675
R112 VN.n108 VN.n59 24.4675
R113 VN.n44 VN.n43 21.5315
R114 VN.n102 VN.n101 21.5315
R115 VN.n56 VN.n55 18.1061
R116 VN.n114 VN.n113 18.1061
R117 VN.n29 VN.n28 12.234
R118 VN.n30 VN.n29 12.234
R119 VN.n88 VN.n87 12.234
R120 VN.n87 VN.n86 12.234
R121 VN.n16 VN.n13 2.93654
R122 VN.n43 VN.n42 2.93654
R123 VN.n74 VN.n71 2.93654
R124 VN.n101 VN.n100 2.93654
R125 VN.n73 VN.n72 2.75934
R126 VN.n15 VN.n14 2.75934
R127 VN.n115 VN.n58 0.417535
R128 VN.n57 VN.n0 0.417535
R129 VN VN.n57 0.394291
R130 VN.n111 VN.n58 0.189894
R131 VN.n111 VN.n110 0.189894
R132 VN.n110 VN.n109 0.189894
R133 VN.n109 VN.n60 0.189894
R134 VN.n105 VN.n60 0.189894
R135 VN.n105 VN.n104 0.189894
R136 VN.n104 VN.n103 0.189894
R137 VN.n103 VN.n62 0.189894
R138 VN.n98 VN.n62 0.189894
R139 VN.n98 VN.n97 0.189894
R140 VN.n97 VN.n96 0.189894
R141 VN.n96 VN.n64 0.189894
R142 VN.n92 VN.n64 0.189894
R143 VN.n92 VN.n91 0.189894
R144 VN.n91 VN.n90 0.189894
R145 VN.n90 VN.n66 0.189894
R146 VN.n85 VN.n66 0.189894
R147 VN.n85 VN.n84 0.189894
R148 VN.n84 VN.n83 0.189894
R149 VN.n83 VN.n68 0.189894
R150 VN.n79 VN.n68 0.189894
R151 VN.n79 VN.n78 0.189894
R152 VN.n78 VN.n77 0.189894
R153 VN.n77 VN.n70 0.189894
R154 VN.n73 VN.n70 0.189894
R155 VN.n15 VN.n12 0.189894
R156 VN.n19 VN.n12 0.189894
R157 VN.n20 VN.n19 0.189894
R158 VN.n21 VN.n20 0.189894
R159 VN.n21 VN.n10 0.189894
R160 VN.n25 VN.n10 0.189894
R161 VN.n26 VN.n25 0.189894
R162 VN.n27 VN.n26 0.189894
R163 VN.n27 VN.n8 0.189894
R164 VN.n32 VN.n8 0.189894
R165 VN.n33 VN.n32 0.189894
R166 VN.n34 VN.n33 0.189894
R167 VN.n34 VN.n6 0.189894
R168 VN.n38 VN.n6 0.189894
R169 VN.n39 VN.n38 0.189894
R170 VN.n40 VN.n39 0.189894
R171 VN.n40 VN.n4 0.189894
R172 VN.n45 VN.n4 0.189894
R173 VN.n46 VN.n45 0.189894
R174 VN.n47 VN.n46 0.189894
R175 VN.n47 VN.n2 0.189894
R176 VN.n51 VN.n2 0.189894
R177 VN.n52 VN.n51 0.189894
R178 VN.n53 VN.n52 0.189894
R179 VN.n53 VN.n0 0.189894
R180 VDD2.n105 VDD2.n57 289.615
R181 VDD2.n48 VDD2.n0 289.615
R182 VDD2.n106 VDD2.n105 185
R183 VDD2.n104 VDD2.n103 185
R184 VDD2.n61 VDD2.n60 185
R185 VDD2.n98 VDD2.n97 185
R186 VDD2.n96 VDD2.n63 185
R187 VDD2.n95 VDD2.n94 185
R188 VDD2.n66 VDD2.n64 185
R189 VDD2.n89 VDD2.n88 185
R190 VDD2.n87 VDD2.n86 185
R191 VDD2.n70 VDD2.n69 185
R192 VDD2.n81 VDD2.n80 185
R193 VDD2.n79 VDD2.n78 185
R194 VDD2.n74 VDD2.n73 185
R195 VDD2.n16 VDD2.n15 185
R196 VDD2.n21 VDD2.n20 185
R197 VDD2.n23 VDD2.n22 185
R198 VDD2.n12 VDD2.n11 185
R199 VDD2.n29 VDD2.n28 185
R200 VDD2.n31 VDD2.n30 185
R201 VDD2.n8 VDD2.n7 185
R202 VDD2.n38 VDD2.n37 185
R203 VDD2.n39 VDD2.n6 185
R204 VDD2.n41 VDD2.n40 185
R205 VDD2.n4 VDD2.n3 185
R206 VDD2.n47 VDD2.n46 185
R207 VDD2.n49 VDD2.n48 185
R208 VDD2.n75 VDD2.t2 149.524
R209 VDD2.n17 VDD2.t7 149.524
R210 VDD2.n105 VDD2.n104 104.615
R211 VDD2.n104 VDD2.n60 104.615
R212 VDD2.n97 VDD2.n60 104.615
R213 VDD2.n97 VDD2.n96 104.615
R214 VDD2.n96 VDD2.n95 104.615
R215 VDD2.n95 VDD2.n64 104.615
R216 VDD2.n88 VDD2.n64 104.615
R217 VDD2.n88 VDD2.n87 104.615
R218 VDD2.n87 VDD2.n69 104.615
R219 VDD2.n80 VDD2.n69 104.615
R220 VDD2.n80 VDD2.n79 104.615
R221 VDD2.n79 VDD2.n73 104.615
R222 VDD2.n21 VDD2.n15 104.615
R223 VDD2.n22 VDD2.n21 104.615
R224 VDD2.n22 VDD2.n11 104.615
R225 VDD2.n29 VDD2.n11 104.615
R226 VDD2.n30 VDD2.n29 104.615
R227 VDD2.n30 VDD2.n7 104.615
R228 VDD2.n38 VDD2.n7 104.615
R229 VDD2.n39 VDD2.n38 104.615
R230 VDD2.n40 VDD2.n39 104.615
R231 VDD2.n40 VDD2.n3 104.615
R232 VDD2.n47 VDD2.n3 104.615
R233 VDD2.n48 VDD2.n47 104.615
R234 VDD2.n56 VDD2.n55 66.729
R235 VDD2 VDD2.n113 66.7262
R236 VDD2.n112 VDD2.n111 63.9979
R237 VDD2.n54 VDD2.n53 63.9977
R238 VDD2.n54 VDD2.n52 53.9372
R239 VDD2.t2 VDD2.n73 52.3082
R240 VDD2.t7 VDD2.n15 52.3082
R241 VDD2.n110 VDD2.n109 50.2217
R242 VDD2.n110 VDD2.n56 50.0106
R243 VDD2.n98 VDD2.n63 13.1884
R244 VDD2.n41 VDD2.n6 13.1884
R245 VDD2.n99 VDD2.n61 12.8005
R246 VDD2.n94 VDD2.n65 12.8005
R247 VDD2.n37 VDD2.n36 12.8005
R248 VDD2.n42 VDD2.n4 12.8005
R249 VDD2.n103 VDD2.n102 12.0247
R250 VDD2.n93 VDD2.n66 12.0247
R251 VDD2.n35 VDD2.n8 12.0247
R252 VDD2.n46 VDD2.n45 12.0247
R253 VDD2.n106 VDD2.n59 11.249
R254 VDD2.n90 VDD2.n89 11.249
R255 VDD2.n32 VDD2.n31 11.249
R256 VDD2.n49 VDD2.n2 11.249
R257 VDD2.n107 VDD2.n57 10.4732
R258 VDD2.n86 VDD2.n68 10.4732
R259 VDD2.n28 VDD2.n10 10.4732
R260 VDD2.n50 VDD2.n0 10.4732
R261 VDD2.n75 VDD2.n74 10.2747
R262 VDD2.n17 VDD2.n16 10.2747
R263 VDD2.n85 VDD2.n70 9.69747
R264 VDD2.n27 VDD2.n12 9.69747
R265 VDD2.n109 VDD2.n108 9.45567
R266 VDD2.n52 VDD2.n51 9.45567
R267 VDD2.n77 VDD2.n76 9.3005
R268 VDD2.n72 VDD2.n71 9.3005
R269 VDD2.n83 VDD2.n82 9.3005
R270 VDD2.n85 VDD2.n84 9.3005
R271 VDD2.n68 VDD2.n67 9.3005
R272 VDD2.n91 VDD2.n90 9.3005
R273 VDD2.n93 VDD2.n92 9.3005
R274 VDD2.n65 VDD2.n62 9.3005
R275 VDD2.n108 VDD2.n107 9.3005
R276 VDD2.n59 VDD2.n58 9.3005
R277 VDD2.n102 VDD2.n101 9.3005
R278 VDD2.n100 VDD2.n99 9.3005
R279 VDD2.n51 VDD2.n50 9.3005
R280 VDD2.n2 VDD2.n1 9.3005
R281 VDD2.n45 VDD2.n44 9.3005
R282 VDD2.n43 VDD2.n42 9.3005
R283 VDD2.n19 VDD2.n18 9.3005
R284 VDD2.n14 VDD2.n13 9.3005
R285 VDD2.n25 VDD2.n24 9.3005
R286 VDD2.n27 VDD2.n26 9.3005
R287 VDD2.n10 VDD2.n9 9.3005
R288 VDD2.n33 VDD2.n32 9.3005
R289 VDD2.n35 VDD2.n34 9.3005
R290 VDD2.n36 VDD2.n5 9.3005
R291 VDD2.n82 VDD2.n81 8.92171
R292 VDD2.n24 VDD2.n23 8.92171
R293 VDD2.n78 VDD2.n72 8.14595
R294 VDD2.n20 VDD2.n14 8.14595
R295 VDD2.n77 VDD2.n74 7.3702
R296 VDD2.n19 VDD2.n16 7.3702
R297 VDD2.n78 VDD2.n77 5.81868
R298 VDD2.n20 VDD2.n19 5.81868
R299 VDD2.n81 VDD2.n72 5.04292
R300 VDD2.n23 VDD2.n14 5.04292
R301 VDD2.n82 VDD2.n70 4.26717
R302 VDD2.n24 VDD2.n12 4.26717
R303 VDD2.n112 VDD2.n110 3.71602
R304 VDD2.n109 VDD2.n57 3.49141
R305 VDD2.n86 VDD2.n85 3.49141
R306 VDD2.n28 VDD2.n27 3.49141
R307 VDD2.n52 VDD2.n0 3.49141
R308 VDD2.n76 VDD2.n75 2.84303
R309 VDD2.n18 VDD2.n17 2.84303
R310 VDD2.n107 VDD2.n106 2.71565
R311 VDD2.n89 VDD2.n68 2.71565
R312 VDD2.n31 VDD2.n10 2.71565
R313 VDD2.n50 VDD2.n49 2.71565
R314 VDD2.n113 VDD2.t8 1.97458
R315 VDD2.n113 VDD2.t9 1.97458
R316 VDD2.n111 VDD2.t6 1.97458
R317 VDD2.n111 VDD2.t3 1.97458
R318 VDD2.n55 VDD2.t0 1.97458
R319 VDD2.n55 VDD2.t5 1.97458
R320 VDD2.n53 VDD2.t4 1.97458
R321 VDD2.n53 VDD2.t1 1.97458
R322 VDD2.n103 VDD2.n59 1.93989
R323 VDD2.n90 VDD2.n66 1.93989
R324 VDD2.n32 VDD2.n8 1.93989
R325 VDD2.n46 VDD2.n2 1.93989
R326 VDD2.n102 VDD2.n61 1.16414
R327 VDD2.n94 VDD2.n93 1.16414
R328 VDD2.n37 VDD2.n35 1.16414
R329 VDD2.n45 VDD2.n4 1.16414
R330 VDD2 VDD2.n112 0.987569
R331 VDD2.n56 VDD2.n54 0.874033
R332 VDD2.n99 VDD2.n98 0.388379
R333 VDD2.n65 VDD2.n63 0.388379
R334 VDD2.n36 VDD2.n6 0.388379
R335 VDD2.n42 VDD2.n41 0.388379
R336 VDD2.n108 VDD2.n58 0.155672
R337 VDD2.n101 VDD2.n58 0.155672
R338 VDD2.n101 VDD2.n100 0.155672
R339 VDD2.n100 VDD2.n62 0.155672
R340 VDD2.n92 VDD2.n62 0.155672
R341 VDD2.n92 VDD2.n91 0.155672
R342 VDD2.n91 VDD2.n67 0.155672
R343 VDD2.n84 VDD2.n67 0.155672
R344 VDD2.n84 VDD2.n83 0.155672
R345 VDD2.n83 VDD2.n71 0.155672
R346 VDD2.n76 VDD2.n71 0.155672
R347 VDD2.n18 VDD2.n13 0.155672
R348 VDD2.n25 VDD2.n13 0.155672
R349 VDD2.n26 VDD2.n25 0.155672
R350 VDD2.n26 VDD2.n9 0.155672
R351 VDD2.n33 VDD2.n9 0.155672
R352 VDD2.n34 VDD2.n33 0.155672
R353 VDD2.n34 VDD2.n5 0.155672
R354 VDD2.n43 VDD2.n5 0.155672
R355 VDD2.n44 VDD2.n43 0.155672
R356 VDD2.n44 VDD2.n1 0.155672
R357 VDD2.n51 VDD2.n1 0.155672
R358 VTAIL.n224 VTAIL.n176 289.615
R359 VTAIL.n50 VTAIL.n2 289.615
R360 VTAIL.n170 VTAIL.n122 289.615
R361 VTAIL.n112 VTAIL.n64 289.615
R362 VTAIL.n192 VTAIL.n191 185
R363 VTAIL.n197 VTAIL.n196 185
R364 VTAIL.n199 VTAIL.n198 185
R365 VTAIL.n188 VTAIL.n187 185
R366 VTAIL.n205 VTAIL.n204 185
R367 VTAIL.n207 VTAIL.n206 185
R368 VTAIL.n184 VTAIL.n183 185
R369 VTAIL.n214 VTAIL.n213 185
R370 VTAIL.n215 VTAIL.n182 185
R371 VTAIL.n217 VTAIL.n216 185
R372 VTAIL.n180 VTAIL.n179 185
R373 VTAIL.n223 VTAIL.n222 185
R374 VTAIL.n225 VTAIL.n224 185
R375 VTAIL.n18 VTAIL.n17 185
R376 VTAIL.n23 VTAIL.n22 185
R377 VTAIL.n25 VTAIL.n24 185
R378 VTAIL.n14 VTAIL.n13 185
R379 VTAIL.n31 VTAIL.n30 185
R380 VTAIL.n33 VTAIL.n32 185
R381 VTAIL.n10 VTAIL.n9 185
R382 VTAIL.n40 VTAIL.n39 185
R383 VTAIL.n41 VTAIL.n8 185
R384 VTAIL.n43 VTAIL.n42 185
R385 VTAIL.n6 VTAIL.n5 185
R386 VTAIL.n49 VTAIL.n48 185
R387 VTAIL.n51 VTAIL.n50 185
R388 VTAIL.n171 VTAIL.n170 185
R389 VTAIL.n169 VTAIL.n168 185
R390 VTAIL.n126 VTAIL.n125 185
R391 VTAIL.n163 VTAIL.n162 185
R392 VTAIL.n161 VTAIL.n128 185
R393 VTAIL.n160 VTAIL.n159 185
R394 VTAIL.n131 VTAIL.n129 185
R395 VTAIL.n154 VTAIL.n153 185
R396 VTAIL.n152 VTAIL.n151 185
R397 VTAIL.n135 VTAIL.n134 185
R398 VTAIL.n146 VTAIL.n145 185
R399 VTAIL.n144 VTAIL.n143 185
R400 VTAIL.n139 VTAIL.n138 185
R401 VTAIL.n113 VTAIL.n112 185
R402 VTAIL.n111 VTAIL.n110 185
R403 VTAIL.n68 VTAIL.n67 185
R404 VTAIL.n105 VTAIL.n104 185
R405 VTAIL.n103 VTAIL.n70 185
R406 VTAIL.n102 VTAIL.n101 185
R407 VTAIL.n73 VTAIL.n71 185
R408 VTAIL.n96 VTAIL.n95 185
R409 VTAIL.n94 VTAIL.n93 185
R410 VTAIL.n77 VTAIL.n76 185
R411 VTAIL.n88 VTAIL.n87 185
R412 VTAIL.n86 VTAIL.n85 185
R413 VTAIL.n81 VTAIL.n80 185
R414 VTAIL.n193 VTAIL.t17 149.524
R415 VTAIL.n19 VTAIL.t7 149.524
R416 VTAIL.n140 VTAIL.t4 149.524
R417 VTAIL.n82 VTAIL.t10 149.524
R418 VTAIL.n197 VTAIL.n191 104.615
R419 VTAIL.n198 VTAIL.n197 104.615
R420 VTAIL.n198 VTAIL.n187 104.615
R421 VTAIL.n205 VTAIL.n187 104.615
R422 VTAIL.n206 VTAIL.n205 104.615
R423 VTAIL.n206 VTAIL.n183 104.615
R424 VTAIL.n214 VTAIL.n183 104.615
R425 VTAIL.n215 VTAIL.n214 104.615
R426 VTAIL.n216 VTAIL.n215 104.615
R427 VTAIL.n216 VTAIL.n179 104.615
R428 VTAIL.n223 VTAIL.n179 104.615
R429 VTAIL.n224 VTAIL.n223 104.615
R430 VTAIL.n23 VTAIL.n17 104.615
R431 VTAIL.n24 VTAIL.n23 104.615
R432 VTAIL.n24 VTAIL.n13 104.615
R433 VTAIL.n31 VTAIL.n13 104.615
R434 VTAIL.n32 VTAIL.n31 104.615
R435 VTAIL.n32 VTAIL.n9 104.615
R436 VTAIL.n40 VTAIL.n9 104.615
R437 VTAIL.n41 VTAIL.n40 104.615
R438 VTAIL.n42 VTAIL.n41 104.615
R439 VTAIL.n42 VTAIL.n5 104.615
R440 VTAIL.n49 VTAIL.n5 104.615
R441 VTAIL.n50 VTAIL.n49 104.615
R442 VTAIL.n170 VTAIL.n169 104.615
R443 VTAIL.n169 VTAIL.n125 104.615
R444 VTAIL.n162 VTAIL.n125 104.615
R445 VTAIL.n162 VTAIL.n161 104.615
R446 VTAIL.n161 VTAIL.n160 104.615
R447 VTAIL.n160 VTAIL.n129 104.615
R448 VTAIL.n153 VTAIL.n129 104.615
R449 VTAIL.n153 VTAIL.n152 104.615
R450 VTAIL.n152 VTAIL.n134 104.615
R451 VTAIL.n145 VTAIL.n134 104.615
R452 VTAIL.n145 VTAIL.n144 104.615
R453 VTAIL.n144 VTAIL.n138 104.615
R454 VTAIL.n112 VTAIL.n111 104.615
R455 VTAIL.n111 VTAIL.n67 104.615
R456 VTAIL.n104 VTAIL.n67 104.615
R457 VTAIL.n104 VTAIL.n103 104.615
R458 VTAIL.n103 VTAIL.n102 104.615
R459 VTAIL.n102 VTAIL.n71 104.615
R460 VTAIL.n95 VTAIL.n71 104.615
R461 VTAIL.n95 VTAIL.n94 104.615
R462 VTAIL.n94 VTAIL.n76 104.615
R463 VTAIL.n87 VTAIL.n76 104.615
R464 VTAIL.n87 VTAIL.n86 104.615
R465 VTAIL.n86 VTAIL.n80 104.615
R466 VTAIL.t17 VTAIL.n191 52.3082
R467 VTAIL.t7 VTAIL.n17 52.3082
R468 VTAIL.t4 VTAIL.n138 52.3082
R469 VTAIL.t10 VTAIL.n80 52.3082
R470 VTAIL.n121 VTAIL.n120 47.3191
R471 VTAIL.n119 VTAIL.n118 47.3191
R472 VTAIL.n63 VTAIL.n62 47.3191
R473 VTAIL.n61 VTAIL.n60 47.3191
R474 VTAIL.n231 VTAIL.n230 47.3189
R475 VTAIL.n1 VTAIL.n0 47.3189
R476 VTAIL.n57 VTAIL.n56 47.3189
R477 VTAIL.n59 VTAIL.n58 47.3189
R478 VTAIL.n229 VTAIL.n228 33.5429
R479 VTAIL.n55 VTAIL.n54 33.5429
R480 VTAIL.n175 VTAIL.n174 33.5429
R481 VTAIL.n117 VTAIL.n116 33.5429
R482 VTAIL.n61 VTAIL.n59 28.4445
R483 VTAIL.n229 VTAIL.n175 24.7289
R484 VTAIL.n217 VTAIL.n182 13.1884
R485 VTAIL.n43 VTAIL.n8 13.1884
R486 VTAIL.n163 VTAIL.n128 13.1884
R487 VTAIL.n105 VTAIL.n70 13.1884
R488 VTAIL.n213 VTAIL.n212 12.8005
R489 VTAIL.n218 VTAIL.n180 12.8005
R490 VTAIL.n39 VTAIL.n38 12.8005
R491 VTAIL.n44 VTAIL.n6 12.8005
R492 VTAIL.n164 VTAIL.n126 12.8005
R493 VTAIL.n159 VTAIL.n130 12.8005
R494 VTAIL.n106 VTAIL.n68 12.8005
R495 VTAIL.n101 VTAIL.n72 12.8005
R496 VTAIL.n211 VTAIL.n184 12.0247
R497 VTAIL.n222 VTAIL.n221 12.0247
R498 VTAIL.n37 VTAIL.n10 12.0247
R499 VTAIL.n48 VTAIL.n47 12.0247
R500 VTAIL.n168 VTAIL.n167 12.0247
R501 VTAIL.n158 VTAIL.n131 12.0247
R502 VTAIL.n110 VTAIL.n109 12.0247
R503 VTAIL.n100 VTAIL.n73 12.0247
R504 VTAIL.n208 VTAIL.n207 11.249
R505 VTAIL.n225 VTAIL.n178 11.249
R506 VTAIL.n34 VTAIL.n33 11.249
R507 VTAIL.n51 VTAIL.n4 11.249
R508 VTAIL.n171 VTAIL.n124 11.249
R509 VTAIL.n155 VTAIL.n154 11.249
R510 VTAIL.n113 VTAIL.n66 11.249
R511 VTAIL.n97 VTAIL.n96 11.249
R512 VTAIL.n204 VTAIL.n186 10.4732
R513 VTAIL.n226 VTAIL.n176 10.4732
R514 VTAIL.n30 VTAIL.n12 10.4732
R515 VTAIL.n52 VTAIL.n2 10.4732
R516 VTAIL.n172 VTAIL.n122 10.4732
R517 VTAIL.n151 VTAIL.n133 10.4732
R518 VTAIL.n114 VTAIL.n64 10.4732
R519 VTAIL.n93 VTAIL.n75 10.4732
R520 VTAIL.n193 VTAIL.n192 10.2747
R521 VTAIL.n19 VTAIL.n18 10.2747
R522 VTAIL.n140 VTAIL.n139 10.2747
R523 VTAIL.n82 VTAIL.n81 10.2747
R524 VTAIL.n203 VTAIL.n188 9.69747
R525 VTAIL.n29 VTAIL.n14 9.69747
R526 VTAIL.n150 VTAIL.n135 9.69747
R527 VTAIL.n92 VTAIL.n77 9.69747
R528 VTAIL.n228 VTAIL.n227 9.45567
R529 VTAIL.n54 VTAIL.n53 9.45567
R530 VTAIL.n174 VTAIL.n173 9.45567
R531 VTAIL.n116 VTAIL.n115 9.45567
R532 VTAIL.n227 VTAIL.n226 9.3005
R533 VTAIL.n178 VTAIL.n177 9.3005
R534 VTAIL.n221 VTAIL.n220 9.3005
R535 VTAIL.n219 VTAIL.n218 9.3005
R536 VTAIL.n195 VTAIL.n194 9.3005
R537 VTAIL.n190 VTAIL.n189 9.3005
R538 VTAIL.n201 VTAIL.n200 9.3005
R539 VTAIL.n203 VTAIL.n202 9.3005
R540 VTAIL.n186 VTAIL.n185 9.3005
R541 VTAIL.n209 VTAIL.n208 9.3005
R542 VTAIL.n211 VTAIL.n210 9.3005
R543 VTAIL.n212 VTAIL.n181 9.3005
R544 VTAIL.n53 VTAIL.n52 9.3005
R545 VTAIL.n4 VTAIL.n3 9.3005
R546 VTAIL.n47 VTAIL.n46 9.3005
R547 VTAIL.n45 VTAIL.n44 9.3005
R548 VTAIL.n21 VTAIL.n20 9.3005
R549 VTAIL.n16 VTAIL.n15 9.3005
R550 VTAIL.n27 VTAIL.n26 9.3005
R551 VTAIL.n29 VTAIL.n28 9.3005
R552 VTAIL.n12 VTAIL.n11 9.3005
R553 VTAIL.n35 VTAIL.n34 9.3005
R554 VTAIL.n37 VTAIL.n36 9.3005
R555 VTAIL.n38 VTAIL.n7 9.3005
R556 VTAIL.n142 VTAIL.n141 9.3005
R557 VTAIL.n137 VTAIL.n136 9.3005
R558 VTAIL.n148 VTAIL.n147 9.3005
R559 VTAIL.n150 VTAIL.n149 9.3005
R560 VTAIL.n133 VTAIL.n132 9.3005
R561 VTAIL.n156 VTAIL.n155 9.3005
R562 VTAIL.n158 VTAIL.n157 9.3005
R563 VTAIL.n130 VTAIL.n127 9.3005
R564 VTAIL.n173 VTAIL.n172 9.3005
R565 VTAIL.n124 VTAIL.n123 9.3005
R566 VTAIL.n167 VTAIL.n166 9.3005
R567 VTAIL.n165 VTAIL.n164 9.3005
R568 VTAIL.n84 VTAIL.n83 9.3005
R569 VTAIL.n79 VTAIL.n78 9.3005
R570 VTAIL.n90 VTAIL.n89 9.3005
R571 VTAIL.n92 VTAIL.n91 9.3005
R572 VTAIL.n75 VTAIL.n74 9.3005
R573 VTAIL.n98 VTAIL.n97 9.3005
R574 VTAIL.n100 VTAIL.n99 9.3005
R575 VTAIL.n72 VTAIL.n69 9.3005
R576 VTAIL.n115 VTAIL.n114 9.3005
R577 VTAIL.n66 VTAIL.n65 9.3005
R578 VTAIL.n109 VTAIL.n108 9.3005
R579 VTAIL.n107 VTAIL.n106 9.3005
R580 VTAIL.n200 VTAIL.n199 8.92171
R581 VTAIL.n26 VTAIL.n25 8.92171
R582 VTAIL.n147 VTAIL.n146 8.92171
R583 VTAIL.n89 VTAIL.n88 8.92171
R584 VTAIL.n196 VTAIL.n190 8.14595
R585 VTAIL.n22 VTAIL.n16 8.14595
R586 VTAIL.n143 VTAIL.n137 8.14595
R587 VTAIL.n85 VTAIL.n79 8.14595
R588 VTAIL.n195 VTAIL.n192 7.3702
R589 VTAIL.n21 VTAIL.n18 7.3702
R590 VTAIL.n142 VTAIL.n139 7.3702
R591 VTAIL.n84 VTAIL.n81 7.3702
R592 VTAIL.n196 VTAIL.n195 5.81868
R593 VTAIL.n22 VTAIL.n21 5.81868
R594 VTAIL.n143 VTAIL.n142 5.81868
R595 VTAIL.n85 VTAIL.n84 5.81868
R596 VTAIL.n199 VTAIL.n190 5.04292
R597 VTAIL.n25 VTAIL.n16 5.04292
R598 VTAIL.n146 VTAIL.n137 5.04292
R599 VTAIL.n88 VTAIL.n79 5.04292
R600 VTAIL.n200 VTAIL.n188 4.26717
R601 VTAIL.n26 VTAIL.n14 4.26717
R602 VTAIL.n147 VTAIL.n135 4.26717
R603 VTAIL.n89 VTAIL.n77 4.26717
R604 VTAIL.n63 VTAIL.n61 3.71602
R605 VTAIL.n117 VTAIL.n63 3.71602
R606 VTAIL.n121 VTAIL.n119 3.71602
R607 VTAIL.n175 VTAIL.n121 3.71602
R608 VTAIL.n59 VTAIL.n57 3.71602
R609 VTAIL.n57 VTAIL.n55 3.71602
R610 VTAIL.n231 VTAIL.n229 3.71602
R611 VTAIL.n204 VTAIL.n203 3.49141
R612 VTAIL.n228 VTAIL.n176 3.49141
R613 VTAIL.n30 VTAIL.n29 3.49141
R614 VTAIL.n54 VTAIL.n2 3.49141
R615 VTAIL.n174 VTAIL.n122 3.49141
R616 VTAIL.n151 VTAIL.n150 3.49141
R617 VTAIL.n116 VTAIL.n64 3.49141
R618 VTAIL.n93 VTAIL.n92 3.49141
R619 VTAIL VTAIL.n1 2.84533
R620 VTAIL.n194 VTAIL.n193 2.84303
R621 VTAIL.n20 VTAIL.n19 2.84303
R622 VTAIL.n141 VTAIL.n140 2.84303
R623 VTAIL.n83 VTAIL.n82 2.84303
R624 VTAIL.n207 VTAIL.n186 2.71565
R625 VTAIL.n226 VTAIL.n225 2.71565
R626 VTAIL.n33 VTAIL.n12 2.71565
R627 VTAIL.n52 VTAIL.n51 2.71565
R628 VTAIL.n172 VTAIL.n171 2.71565
R629 VTAIL.n154 VTAIL.n133 2.71565
R630 VTAIL.n114 VTAIL.n113 2.71565
R631 VTAIL.n96 VTAIL.n75 2.71565
R632 VTAIL.n119 VTAIL.n117 2.32809
R633 VTAIL.n55 VTAIL.n1 2.32809
R634 VTAIL.n230 VTAIL.t11 1.97458
R635 VTAIL.n230 VTAIL.t18 1.97458
R636 VTAIL.n0 VTAIL.t16 1.97458
R637 VTAIL.n0 VTAIL.t12 1.97458
R638 VTAIL.n56 VTAIL.t1 1.97458
R639 VTAIL.n56 VTAIL.t3 1.97458
R640 VTAIL.n58 VTAIL.t2 1.97458
R641 VTAIL.n58 VTAIL.t5 1.97458
R642 VTAIL.n120 VTAIL.t6 1.97458
R643 VTAIL.n120 VTAIL.t0 1.97458
R644 VTAIL.n118 VTAIL.t19 1.97458
R645 VTAIL.n118 VTAIL.t8 1.97458
R646 VTAIL.n62 VTAIL.t9 1.97458
R647 VTAIL.n62 VTAIL.t14 1.97458
R648 VTAIL.n60 VTAIL.t13 1.97458
R649 VTAIL.n60 VTAIL.t15 1.97458
R650 VTAIL.n208 VTAIL.n184 1.93989
R651 VTAIL.n222 VTAIL.n178 1.93989
R652 VTAIL.n34 VTAIL.n10 1.93989
R653 VTAIL.n48 VTAIL.n4 1.93989
R654 VTAIL.n168 VTAIL.n124 1.93989
R655 VTAIL.n155 VTAIL.n131 1.93989
R656 VTAIL.n110 VTAIL.n66 1.93989
R657 VTAIL.n97 VTAIL.n73 1.93989
R658 VTAIL.n213 VTAIL.n211 1.16414
R659 VTAIL.n221 VTAIL.n180 1.16414
R660 VTAIL.n39 VTAIL.n37 1.16414
R661 VTAIL.n47 VTAIL.n6 1.16414
R662 VTAIL.n167 VTAIL.n126 1.16414
R663 VTAIL.n159 VTAIL.n158 1.16414
R664 VTAIL.n109 VTAIL.n68 1.16414
R665 VTAIL.n101 VTAIL.n100 1.16414
R666 VTAIL VTAIL.n231 0.87119
R667 VTAIL.n212 VTAIL.n182 0.388379
R668 VTAIL.n218 VTAIL.n217 0.388379
R669 VTAIL.n38 VTAIL.n8 0.388379
R670 VTAIL.n44 VTAIL.n43 0.388379
R671 VTAIL.n164 VTAIL.n163 0.388379
R672 VTAIL.n130 VTAIL.n128 0.388379
R673 VTAIL.n106 VTAIL.n105 0.388379
R674 VTAIL.n72 VTAIL.n70 0.388379
R675 VTAIL.n194 VTAIL.n189 0.155672
R676 VTAIL.n201 VTAIL.n189 0.155672
R677 VTAIL.n202 VTAIL.n201 0.155672
R678 VTAIL.n202 VTAIL.n185 0.155672
R679 VTAIL.n209 VTAIL.n185 0.155672
R680 VTAIL.n210 VTAIL.n209 0.155672
R681 VTAIL.n210 VTAIL.n181 0.155672
R682 VTAIL.n219 VTAIL.n181 0.155672
R683 VTAIL.n220 VTAIL.n219 0.155672
R684 VTAIL.n220 VTAIL.n177 0.155672
R685 VTAIL.n227 VTAIL.n177 0.155672
R686 VTAIL.n20 VTAIL.n15 0.155672
R687 VTAIL.n27 VTAIL.n15 0.155672
R688 VTAIL.n28 VTAIL.n27 0.155672
R689 VTAIL.n28 VTAIL.n11 0.155672
R690 VTAIL.n35 VTAIL.n11 0.155672
R691 VTAIL.n36 VTAIL.n35 0.155672
R692 VTAIL.n36 VTAIL.n7 0.155672
R693 VTAIL.n45 VTAIL.n7 0.155672
R694 VTAIL.n46 VTAIL.n45 0.155672
R695 VTAIL.n46 VTAIL.n3 0.155672
R696 VTAIL.n53 VTAIL.n3 0.155672
R697 VTAIL.n173 VTAIL.n123 0.155672
R698 VTAIL.n166 VTAIL.n123 0.155672
R699 VTAIL.n166 VTAIL.n165 0.155672
R700 VTAIL.n165 VTAIL.n127 0.155672
R701 VTAIL.n157 VTAIL.n127 0.155672
R702 VTAIL.n157 VTAIL.n156 0.155672
R703 VTAIL.n156 VTAIL.n132 0.155672
R704 VTAIL.n149 VTAIL.n132 0.155672
R705 VTAIL.n149 VTAIL.n148 0.155672
R706 VTAIL.n148 VTAIL.n136 0.155672
R707 VTAIL.n141 VTAIL.n136 0.155672
R708 VTAIL.n115 VTAIL.n65 0.155672
R709 VTAIL.n108 VTAIL.n65 0.155672
R710 VTAIL.n108 VTAIL.n107 0.155672
R711 VTAIL.n107 VTAIL.n69 0.155672
R712 VTAIL.n99 VTAIL.n69 0.155672
R713 VTAIL.n99 VTAIL.n98 0.155672
R714 VTAIL.n98 VTAIL.n74 0.155672
R715 VTAIL.n91 VTAIL.n74 0.155672
R716 VTAIL.n91 VTAIL.n90 0.155672
R717 VTAIL.n90 VTAIL.n78 0.155672
R718 VTAIL.n83 VTAIL.n78 0.155672
R719 B.n1090 B.n1089 585
R720 B.n1091 B.n1090 585
R721 B.n356 B.n193 585
R722 B.n355 B.n354 585
R723 B.n353 B.n352 585
R724 B.n351 B.n350 585
R725 B.n349 B.n348 585
R726 B.n347 B.n346 585
R727 B.n345 B.n344 585
R728 B.n343 B.n342 585
R729 B.n341 B.n340 585
R730 B.n339 B.n338 585
R731 B.n337 B.n336 585
R732 B.n335 B.n334 585
R733 B.n333 B.n332 585
R734 B.n331 B.n330 585
R735 B.n329 B.n328 585
R736 B.n327 B.n326 585
R737 B.n325 B.n324 585
R738 B.n323 B.n322 585
R739 B.n321 B.n320 585
R740 B.n319 B.n318 585
R741 B.n317 B.n316 585
R742 B.n315 B.n314 585
R743 B.n313 B.n312 585
R744 B.n311 B.n310 585
R745 B.n309 B.n308 585
R746 B.n307 B.n306 585
R747 B.n305 B.n304 585
R748 B.n303 B.n302 585
R749 B.n301 B.n300 585
R750 B.n299 B.n298 585
R751 B.n297 B.n296 585
R752 B.n295 B.n294 585
R753 B.n293 B.n292 585
R754 B.n291 B.n290 585
R755 B.n289 B.n288 585
R756 B.n286 B.n285 585
R757 B.n284 B.n283 585
R758 B.n282 B.n281 585
R759 B.n280 B.n279 585
R760 B.n278 B.n277 585
R761 B.n276 B.n275 585
R762 B.n274 B.n273 585
R763 B.n272 B.n271 585
R764 B.n270 B.n269 585
R765 B.n268 B.n267 585
R766 B.n266 B.n265 585
R767 B.n264 B.n263 585
R768 B.n262 B.n261 585
R769 B.n260 B.n259 585
R770 B.n258 B.n257 585
R771 B.n256 B.n255 585
R772 B.n254 B.n253 585
R773 B.n252 B.n251 585
R774 B.n250 B.n249 585
R775 B.n248 B.n247 585
R776 B.n246 B.n245 585
R777 B.n244 B.n243 585
R778 B.n242 B.n241 585
R779 B.n240 B.n239 585
R780 B.n238 B.n237 585
R781 B.n236 B.n235 585
R782 B.n234 B.n233 585
R783 B.n232 B.n231 585
R784 B.n230 B.n229 585
R785 B.n228 B.n227 585
R786 B.n226 B.n225 585
R787 B.n224 B.n223 585
R788 B.n222 B.n221 585
R789 B.n220 B.n219 585
R790 B.n218 B.n217 585
R791 B.n216 B.n215 585
R792 B.n214 B.n213 585
R793 B.n212 B.n211 585
R794 B.n210 B.n209 585
R795 B.n208 B.n207 585
R796 B.n206 B.n205 585
R797 B.n204 B.n203 585
R798 B.n202 B.n201 585
R799 B.n200 B.n199 585
R800 B.n151 B.n150 585
R801 B.n1088 B.n152 585
R802 B.n1092 B.n152 585
R803 B.n1087 B.n1086 585
R804 B.n1086 B.n148 585
R805 B.n1085 B.n147 585
R806 B.n1098 B.n147 585
R807 B.n1084 B.n146 585
R808 B.n1099 B.n146 585
R809 B.n1083 B.n145 585
R810 B.n1100 B.n145 585
R811 B.n1082 B.n1081 585
R812 B.n1081 B.n141 585
R813 B.n1080 B.n140 585
R814 B.n1106 B.n140 585
R815 B.n1079 B.n139 585
R816 B.n1107 B.n139 585
R817 B.n1078 B.n138 585
R818 B.n1108 B.n138 585
R819 B.n1077 B.n1076 585
R820 B.n1076 B.n137 585
R821 B.n1075 B.n133 585
R822 B.n1114 B.n133 585
R823 B.n1074 B.n132 585
R824 B.n1115 B.n132 585
R825 B.n1073 B.n131 585
R826 B.n1116 B.n131 585
R827 B.n1072 B.n1071 585
R828 B.n1071 B.n127 585
R829 B.n1070 B.n126 585
R830 B.n1122 B.n126 585
R831 B.n1069 B.n125 585
R832 B.n1123 B.n125 585
R833 B.n1068 B.n124 585
R834 B.n1124 B.n124 585
R835 B.n1067 B.n1066 585
R836 B.n1066 B.n120 585
R837 B.n1065 B.n119 585
R838 B.n1130 B.n119 585
R839 B.n1064 B.n118 585
R840 B.n1131 B.n118 585
R841 B.n1063 B.n117 585
R842 B.n1132 B.n117 585
R843 B.n1062 B.n1061 585
R844 B.n1061 B.n113 585
R845 B.n1060 B.n112 585
R846 B.n1138 B.n112 585
R847 B.n1059 B.n111 585
R848 B.n1139 B.n111 585
R849 B.n1058 B.n110 585
R850 B.n1140 B.n110 585
R851 B.n1057 B.n1056 585
R852 B.n1056 B.n109 585
R853 B.n1055 B.n105 585
R854 B.n1146 B.n105 585
R855 B.n1054 B.n104 585
R856 B.n1147 B.n104 585
R857 B.n1053 B.n103 585
R858 B.n1148 B.n103 585
R859 B.n1052 B.n1051 585
R860 B.n1051 B.n99 585
R861 B.n1050 B.n98 585
R862 B.n1154 B.n98 585
R863 B.n1049 B.n97 585
R864 B.n1155 B.n97 585
R865 B.n1048 B.n96 585
R866 B.n1156 B.n96 585
R867 B.n1047 B.n1046 585
R868 B.n1046 B.n92 585
R869 B.n1045 B.n91 585
R870 B.n1162 B.n91 585
R871 B.n1044 B.n90 585
R872 B.n1163 B.n90 585
R873 B.n1043 B.n89 585
R874 B.n1164 B.n89 585
R875 B.n1042 B.n1041 585
R876 B.n1041 B.n85 585
R877 B.n1040 B.n84 585
R878 B.n1170 B.n84 585
R879 B.n1039 B.n83 585
R880 B.n1171 B.n83 585
R881 B.n1038 B.n82 585
R882 B.n1172 B.n82 585
R883 B.n1037 B.n1036 585
R884 B.n1036 B.n78 585
R885 B.n1035 B.n77 585
R886 B.n1178 B.n77 585
R887 B.n1034 B.n76 585
R888 B.n1179 B.n76 585
R889 B.n1033 B.n75 585
R890 B.n1180 B.n75 585
R891 B.n1032 B.n1031 585
R892 B.n1031 B.n71 585
R893 B.n1030 B.n70 585
R894 B.n1186 B.n70 585
R895 B.n1029 B.n69 585
R896 B.n1187 B.n69 585
R897 B.n1028 B.n68 585
R898 B.n1188 B.n68 585
R899 B.n1027 B.n1026 585
R900 B.n1026 B.n64 585
R901 B.n1025 B.n63 585
R902 B.n1194 B.n63 585
R903 B.n1024 B.n62 585
R904 B.n1195 B.n62 585
R905 B.n1023 B.n61 585
R906 B.n1196 B.n61 585
R907 B.n1022 B.n1021 585
R908 B.n1021 B.n57 585
R909 B.n1020 B.n56 585
R910 B.n1202 B.n56 585
R911 B.n1019 B.n55 585
R912 B.n1203 B.n55 585
R913 B.n1018 B.n54 585
R914 B.n1204 B.n54 585
R915 B.n1017 B.n1016 585
R916 B.n1016 B.n50 585
R917 B.n1015 B.n49 585
R918 B.n1210 B.n49 585
R919 B.n1014 B.n48 585
R920 B.n1211 B.n48 585
R921 B.n1013 B.n47 585
R922 B.n1212 B.n47 585
R923 B.n1012 B.n1011 585
R924 B.n1011 B.n43 585
R925 B.n1010 B.n42 585
R926 B.n1218 B.n42 585
R927 B.n1009 B.n41 585
R928 B.n1219 B.n41 585
R929 B.n1008 B.n40 585
R930 B.n1220 B.n40 585
R931 B.n1007 B.n1006 585
R932 B.n1006 B.n36 585
R933 B.n1005 B.n35 585
R934 B.n1226 B.n35 585
R935 B.n1004 B.n34 585
R936 B.n1227 B.n34 585
R937 B.n1003 B.n33 585
R938 B.n1228 B.n33 585
R939 B.n1002 B.n1001 585
R940 B.n1001 B.n29 585
R941 B.n1000 B.n28 585
R942 B.n1234 B.n28 585
R943 B.n999 B.n27 585
R944 B.n1235 B.n27 585
R945 B.n998 B.n26 585
R946 B.n1236 B.n26 585
R947 B.n997 B.n996 585
R948 B.n996 B.n22 585
R949 B.n995 B.n21 585
R950 B.n1242 B.n21 585
R951 B.n994 B.n20 585
R952 B.n1243 B.n20 585
R953 B.n993 B.n19 585
R954 B.n1244 B.n19 585
R955 B.n992 B.n991 585
R956 B.n991 B.n15 585
R957 B.n990 B.n14 585
R958 B.n1250 B.n14 585
R959 B.n989 B.n13 585
R960 B.n1251 B.n13 585
R961 B.n988 B.n12 585
R962 B.n1252 B.n12 585
R963 B.n987 B.n986 585
R964 B.n986 B.n8 585
R965 B.n985 B.n7 585
R966 B.n1258 B.n7 585
R967 B.n984 B.n6 585
R968 B.n1259 B.n6 585
R969 B.n983 B.n5 585
R970 B.n1260 B.n5 585
R971 B.n982 B.n981 585
R972 B.n981 B.n4 585
R973 B.n980 B.n357 585
R974 B.n980 B.n979 585
R975 B.n970 B.n358 585
R976 B.n359 B.n358 585
R977 B.n972 B.n971 585
R978 B.n973 B.n972 585
R979 B.n969 B.n364 585
R980 B.n364 B.n363 585
R981 B.n968 B.n967 585
R982 B.n967 B.n966 585
R983 B.n366 B.n365 585
R984 B.n367 B.n366 585
R985 B.n959 B.n958 585
R986 B.n960 B.n959 585
R987 B.n957 B.n372 585
R988 B.n372 B.n371 585
R989 B.n956 B.n955 585
R990 B.n955 B.n954 585
R991 B.n374 B.n373 585
R992 B.n375 B.n374 585
R993 B.n947 B.n946 585
R994 B.n948 B.n947 585
R995 B.n945 B.n380 585
R996 B.n380 B.n379 585
R997 B.n944 B.n943 585
R998 B.n943 B.n942 585
R999 B.n382 B.n381 585
R1000 B.n383 B.n382 585
R1001 B.n935 B.n934 585
R1002 B.n936 B.n935 585
R1003 B.n933 B.n388 585
R1004 B.n388 B.n387 585
R1005 B.n932 B.n931 585
R1006 B.n931 B.n930 585
R1007 B.n390 B.n389 585
R1008 B.n391 B.n390 585
R1009 B.n923 B.n922 585
R1010 B.n924 B.n923 585
R1011 B.n921 B.n395 585
R1012 B.n399 B.n395 585
R1013 B.n920 B.n919 585
R1014 B.n919 B.n918 585
R1015 B.n397 B.n396 585
R1016 B.n398 B.n397 585
R1017 B.n911 B.n910 585
R1018 B.n912 B.n911 585
R1019 B.n909 B.n404 585
R1020 B.n404 B.n403 585
R1021 B.n908 B.n907 585
R1022 B.n907 B.n906 585
R1023 B.n406 B.n405 585
R1024 B.n407 B.n406 585
R1025 B.n899 B.n898 585
R1026 B.n900 B.n899 585
R1027 B.n897 B.n412 585
R1028 B.n412 B.n411 585
R1029 B.n896 B.n895 585
R1030 B.n895 B.n894 585
R1031 B.n414 B.n413 585
R1032 B.n415 B.n414 585
R1033 B.n887 B.n886 585
R1034 B.n888 B.n887 585
R1035 B.n885 B.n420 585
R1036 B.n420 B.n419 585
R1037 B.n884 B.n883 585
R1038 B.n883 B.n882 585
R1039 B.n422 B.n421 585
R1040 B.n423 B.n422 585
R1041 B.n875 B.n874 585
R1042 B.n876 B.n875 585
R1043 B.n873 B.n428 585
R1044 B.n428 B.n427 585
R1045 B.n872 B.n871 585
R1046 B.n871 B.n870 585
R1047 B.n430 B.n429 585
R1048 B.n431 B.n430 585
R1049 B.n863 B.n862 585
R1050 B.n864 B.n863 585
R1051 B.n861 B.n436 585
R1052 B.n436 B.n435 585
R1053 B.n860 B.n859 585
R1054 B.n859 B.n858 585
R1055 B.n438 B.n437 585
R1056 B.n439 B.n438 585
R1057 B.n851 B.n850 585
R1058 B.n852 B.n851 585
R1059 B.n849 B.n444 585
R1060 B.n444 B.n443 585
R1061 B.n848 B.n847 585
R1062 B.n847 B.n846 585
R1063 B.n446 B.n445 585
R1064 B.n447 B.n446 585
R1065 B.n839 B.n838 585
R1066 B.n840 B.n839 585
R1067 B.n837 B.n452 585
R1068 B.n452 B.n451 585
R1069 B.n836 B.n835 585
R1070 B.n835 B.n834 585
R1071 B.n454 B.n453 585
R1072 B.n455 B.n454 585
R1073 B.n827 B.n826 585
R1074 B.n828 B.n827 585
R1075 B.n825 B.n460 585
R1076 B.n460 B.n459 585
R1077 B.n824 B.n823 585
R1078 B.n823 B.n822 585
R1079 B.n462 B.n461 585
R1080 B.n463 B.n462 585
R1081 B.n815 B.n814 585
R1082 B.n816 B.n815 585
R1083 B.n813 B.n468 585
R1084 B.n468 B.n467 585
R1085 B.n812 B.n811 585
R1086 B.n811 B.n810 585
R1087 B.n470 B.n469 585
R1088 B.n803 B.n470 585
R1089 B.n802 B.n801 585
R1090 B.n804 B.n802 585
R1091 B.n800 B.n475 585
R1092 B.n475 B.n474 585
R1093 B.n799 B.n798 585
R1094 B.n798 B.n797 585
R1095 B.n477 B.n476 585
R1096 B.n478 B.n477 585
R1097 B.n790 B.n789 585
R1098 B.n791 B.n790 585
R1099 B.n788 B.n483 585
R1100 B.n483 B.n482 585
R1101 B.n787 B.n786 585
R1102 B.n786 B.n785 585
R1103 B.n485 B.n484 585
R1104 B.n486 B.n485 585
R1105 B.n778 B.n777 585
R1106 B.n779 B.n778 585
R1107 B.n776 B.n491 585
R1108 B.n491 B.n490 585
R1109 B.n775 B.n774 585
R1110 B.n774 B.n773 585
R1111 B.n493 B.n492 585
R1112 B.n494 B.n493 585
R1113 B.n766 B.n765 585
R1114 B.n767 B.n766 585
R1115 B.n764 B.n499 585
R1116 B.n499 B.n498 585
R1117 B.n763 B.n762 585
R1118 B.n762 B.n761 585
R1119 B.n501 B.n500 585
R1120 B.n754 B.n501 585
R1121 B.n753 B.n752 585
R1122 B.n755 B.n753 585
R1123 B.n751 B.n506 585
R1124 B.n506 B.n505 585
R1125 B.n750 B.n749 585
R1126 B.n749 B.n748 585
R1127 B.n508 B.n507 585
R1128 B.n509 B.n508 585
R1129 B.n741 B.n740 585
R1130 B.n742 B.n741 585
R1131 B.n739 B.n514 585
R1132 B.n514 B.n513 585
R1133 B.n738 B.n737 585
R1134 B.n737 B.n736 585
R1135 B.n516 B.n515 585
R1136 B.n517 B.n516 585
R1137 B.n729 B.n728 585
R1138 B.n730 B.n729 585
R1139 B.n520 B.n519 585
R1140 B.n568 B.n566 585
R1141 B.n569 B.n565 585
R1142 B.n569 B.n521 585
R1143 B.n572 B.n571 585
R1144 B.n573 B.n564 585
R1145 B.n575 B.n574 585
R1146 B.n577 B.n563 585
R1147 B.n580 B.n579 585
R1148 B.n581 B.n562 585
R1149 B.n583 B.n582 585
R1150 B.n585 B.n561 585
R1151 B.n588 B.n587 585
R1152 B.n589 B.n560 585
R1153 B.n591 B.n590 585
R1154 B.n593 B.n559 585
R1155 B.n596 B.n595 585
R1156 B.n597 B.n558 585
R1157 B.n599 B.n598 585
R1158 B.n601 B.n557 585
R1159 B.n604 B.n603 585
R1160 B.n605 B.n556 585
R1161 B.n607 B.n606 585
R1162 B.n609 B.n555 585
R1163 B.n612 B.n611 585
R1164 B.n613 B.n554 585
R1165 B.n615 B.n614 585
R1166 B.n617 B.n553 585
R1167 B.n620 B.n619 585
R1168 B.n621 B.n552 585
R1169 B.n623 B.n622 585
R1170 B.n625 B.n551 585
R1171 B.n628 B.n627 585
R1172 B.n629 B.n550 585
R1173 B.n631 B.n630 585
R1174 B.n633 B.n549 585
R1175 B.n636 B.n635 585
R1176 B.n638 B.n546 585
R1177 B.n640 B.n639 585
R1178 B.n642 B.n545 585
R1179 B.n645 B.n644 585
R1180 B.n646 B.n544 585
R1181 B.n648 B.n647 585
R1182 B.n650 B.n543 585
R1183 B.n653 B.n652 585
R1184 B.n654 B.n540 585
R1185 B.n657 B.n656 585
R1186 B.n659 B.n539 585
R1187 B.n662 B.n661 585
R1188 B.n663 B.n538 585
R1189 B.n665 B.n664 585
R1190 B.n667 B.n537 585
R1191 B.n670 B.n669 585
R1192 B.n671 B.n536 585
R1193 B.n673 B.n672 585
R1194 B.n675 B.n535 585
R1195 B.n678 B.n677 585
R1196 B.n679 B.n534 585
R1197 B.n681 B.n680 585
R1198 B.n683 B.n533 585
R1199 B.n686 B.n685 585
R1200 B.n687 B.n532 585
R1201 B.n689 B.n688 585
R1202 B.n691 B.n531 585
R1203 B.n694 B.n693 585
R1204 B.n695 B.n530 585
R1205 B.n697 B.n696 585
R1206 B.n699 B.n529 585
R1207 B.n702 B.n701 585
R1208 B.n703 B.n528 585
R1209 B.n705 B.n704 585
R1210 B.n707 B.n527 585
R1211 B.n710 B.n709 585
R1212 B.n711 B.n526 585
R1213 B.n713 B.n712 585
R1214 B.n715 B.n525 585
R1215 B.n718 B.n717 585
R1216 B.n719 B.n524 585
R1217 B.n721 B.n720 585
R1218 B.n723 B.n523 585
R1219 B.n726 B.n725 585
R1220 B.n727 B.n522 585
R1221 B.n732 B.n731 585
R1222 B.n731 B.n730 585
R1223 B.n733 B.n518 585
R1224 B.n518 B.n517 585
R1225 B.n735 B.n734 585
R1226 B.n736 B.n735 585
R1227 B.n512 B.n511 585
R1228 B.n513 B.n512 585
R1229 B.n744 B.n743 585
R1230 B.n743 B.n742 585
R1231 B.n745 B.n510 585
R1232 B.n510 B.n509 585
R1233 B.n747 B.n746 585
R1234 B.n748 B.n747 585
R1235 B.n504 B.n503 585
R1236 B.n505 B.n504 585
R1237 B.n757 B.n756 585
R1238 B.n756 B.n755 585
R1239 B.n758 B.n502 585
R1240 B.n754 B.n502 585
R1241 B.n760 B.n759 585
R1242 B.n761 B.n760 585
R1243 B.n497 B.n496 585
R1244 B.n498 B.n497 585
R1245 B.n769 B.n768 585
R1246 B.n768 B.n767 585
R1247 B.n770 B.n495 585
R1248 B.n495 B.n494 585
R1249 B.n772 B.n771 585
R1250 B.n773 B.n772 585
R1251 B.n489 B.n488 585
R1252 B.n490 B.n489 585
R1253 B.n781 B.n780 585
R1254 B.n780 B.n779 585
R1255 B.n782 B.n487 585
R1256 B.n487 B.n486 585
R1257 B.n784 B.n783 585
R1258 B.n785 B.n784 585
R1259 B.n481 B.n480 585
R1260 B.n482 B.n481 585
R1261 B.n793 B.n792 585
R1262 B.n792 B.n791 585
R1263 B.n794 B.n479 585
R1264 B.n479 B.n478 585
R1265 B.n796 B.n795 585
R1266 B.n797 B.n796 585
R1267 B.n473 B.n472 585
R1268 B.n474 B.n473 585
R1269 B.n806 B.n805 585
R1270 B.n805 B.n804 585
R1271 B.n807 B.n471 585
R1272 B.n803 B.n471 585
R1273 B.n809 B.n808 585
R1274 B.n810 B.n809 585
R1275 B.n466 B.n465 585
R1276 B.n467 B.n466 585
R1277 B.n818 B.n817 585
R1278 B.n817 B.n816 585
R1279 B.n819 B.n464 585
R1280 B.n464 B.n463 585
R1281 B.n821 B.n820 585
R1282 B.n822 B.n821 585
R1283 B.n458 B.n457 585
R1284 B.n459 B.n458 585
R1285 B.n830 B.n829 585
R1286 B.n829 B.n828 585
R1287 B.n831 B.n456 585
R1288 B.n456 B.n455 585
R1289 B.n833 B.n832 585
R1290 B.n834 B.n833 585
R1291 B.n450 B.n449 585
R1292 B.n451 B.n450 585
R1293 B.n842 B.n841 585
R1294 B.n841 B.n840 585
R1295 B.n843 B.n448 585
R1296 B.n448 B.n447 585
R1297 B.n845 B.n844 585
R1298 B.n846 B.n845 585
R1299 B.n442 B.n441 585
R1300 B.n443 B.n442 585
R1301 B.n854 B.n853 585
R1302 B.n853 B.n852 585
R1303 B.n855 B.n440 585
R1304 B.n440 B.n439 585
R1305 B.n857 B.n856 585
R1306 B.n858 B.n857 585
R1307 B.n434 B.n433 585
R1308 B.n435 B.n434 585
R1309 B.n866 B.n865 585
R1310 B.n865 B.n864 585
R1311 B.n867 B.n432 585
R1312 B.n432 B.n431 585
R1313 B.n869 B.n868 585
R1314 B.n870 B.n869 585
R1315 B.n426 B.n425 585
R1316 B.n427 B.n426 585
R1317 B.n878 B.n877 585
R1318 B.n877 B.n876 585
R1319 B.n879 B.n424 585
R1320 B.n424 B.n423 585
R1321 B.n881 B.n880 585
R1322 B.n882 B.n881 585
R1323 B.n418 B.n417 585
R1324 B.n419 B.n418 585
R1325 B.n890 B.n889 585
R1326 B.n889 B.n888 585
R1327 B.n891 B.n416 585
R1328 B.n416 B.n415 585
R1329 B.n893 B.n892 585
R1330 B.n894 B.n893 585
R1331 B.n410 B.n409 585
R1332 B.n411 B.n410 585
R1333 B.n902 B.n901 585
R1334 B.n901 B.n900 585
R1335 B.n903 B.n408 585
R1336 B.n408 B.n407 585
R1337 B.n905 B.n904 585
R1338 B.n906 B.n905 585
R1339 B.n402 B.n401 585
R1340 B.n403 B.n402 585
R1341 B.n914 B.n913 585
R1342 B.n913 B.n912 585
R1343 B.n915 B.n400 585
R1344 B.n400 B.n398 585
R1345 B.n917 B.n916 585
R1346 B.n918 B.n917 585
R1347 B.n394 B.n393 585
R1348 B.n399 B.n394 585
R1349 B.n926 B.n925 585
R1350 B.n925 B.n924 585
R1351 B.n927 B.n392 585
R1352 B.n392 B.n391 585
R1353 B.n929 B.n928 585
R1354 B.n930 B.n929 585
R1355 B.n386 B.n385 585
R1356 B.n387 B.n386 585
R1357 B.n938 B.n937 585
R1358 B.n937 B.n936 585
R1359 B.n939 B.n384 585
R1360 B.n384 B.n383 585
R1361 B.n941 B.n940 585
R1362 B.n942 B.n941 585
R1363 B.n378 B.n377 585
R1364 B.n379 B.n378 585
R1365 B.n950 B.n949 585
R1366 B.n949 B.n948 585
R1367 B.n951 B.n376 585
R1368 B.n376 B.n375 585
R1369 B.n953 B.n952 585
R1370 B.n954 B.n953 585
R1371 B.n370 B.n369 585
R1372 B.n371 B.n370 585
R1373 B.n962 B.n961 585
R1374 B.n961 B.n960 585
R1375 B.n963 B.n368 585
R1376 B.n368 B.n367 585
R1377 B.n965 B.n964 585
R1378 B.n966 B.n965 585
R1379 B.n362 B.n361 585
R1380 B.n363 B.n362 585
R1381 B.n975 B.n974 585
R1382 B.n974 B.n973 585
R1383 B.n976 B.n360 585
R1384 B.n360 B.n359 585
R1385 B.n978 B.n977 585
R1386 B.n979 B.n978 585
R1387 B.n2 B.n0 585
R1388 B.n4 B.n2 585
R1389 B.n3 B.n1 585
R1390 B.n1259 B.n3 585
R1391 B.n1257 B.n1256 585
R1392 B.n1258 B.n1257 585
R1393 B.n1255 B.n9 585
R1394 B.n9 B.n8 585
R1395 B.n1254 B.n1253 585
R1396 B.n1253 B.n1252 585
R1397 B.n11 B.n10 585
R1398 B.n1251 B.n11 585
R1399 B.n1249 B.n1248 585
R1400 B.n1250 B.n1249 585
R1401 B.n1247 B.n16 585
R1402 B.n16 B.n15 585
R1403 B.n1246 B.n1245 585
R1404 B.n1245 B.n1244 585
R1405 B.n18 B.n17 585
R1406 B.n1243 B.n18 585
R1407 B.n1241 B.n1240 585
R1408 B.n1242 B.n1241 585
R1409 B.n1239 B.n23 585
R1410 B.n23 B.n22 585
R1411 B.n1238 B.n1237 585
R1412 B.n1237 B.n1236 585
R1413 B.n25 B.n24 585
R1414 B.n1235 B.n25 585
R1415 B.n1233 B.n1232 585
R1416 B.n1234 B.n1233 585
R1417 B.n1231 B.n30 585
R1418 B.n30 B.n29 585
R1419 B.n1230 B.n1229 585
R1420 B.n1229 B.n1228 585
R1421 B.n32 B.n31 585
R1422 B.n1227 B.n32 585
R1423 B.n1225 B.n1224 585
R1424 B.n1226 B.n1225 585
R1425 B.n1223 B.n37 585
R1426 B.n37 B.n36 585
R1427 B.n1222 B.n1221 585
R1428 B.n1221 B.n1220 585
R1429 B.n39 B.n38 585
R1430 B.n1219 B.n39 585
R1431 B.n1217 B.n1216 585
R1432 B.n1218 B.n1217 585
R1433 B.n1215 B.n44 585
R1434 B.n44 B.n43 585
R1435 B.n1214 B.n1213 585
R1436 B.n1213 B.n1212 585
R1437 B.n46 B.n45 585
R1438 B.n1211 B.n46 585
R1439 B.n1209 B.n1208 585
R1440 B.n1210 B.n1209 585
R1441 B.n1207 B.n51 585
R1442 B.n51 B.n50 585
R1443 B.n1206 B.n1205 585
R1444 B.n1205 B.n1204 585
R1445 B.n53 B.n52 585
R1446 B.n1203 B.n53 585
R1447 B.n1201 B.n1200 585
R1448 B.n1202 B.n1201 585
R1449 B.n1199 B.n58 585
R1450 B.n58 B.n57 585
R1451 B.n1198 B.n1197 585
R1452 B.n1197 B.n1196 585
R1453 B.n60 B.n59 585
R1454 B.n1195 B.n60 585
R1455 B.n1193 B.n1192 585
R1456 B.n1194 B.n1193 585
R1457 B.n1191 B.n65 585
R1458 B.n65 B.n64 585
R1459 B.n1190 B.n1189 585
R1460 B.n1189 B.n1188 585
R1461 B.n67 B.n66 585
R1462 B.n1187 B.n67 585
R1463 B.n1185 B.n1184 585
R1464 B.n1186 B.n1185 585
R1465 B.n1183 B.n72 585
R1466 B.n72 B.n71 585
R1467 B.n1182 B.n1181 585
R1468 B.n1181 B.n1180 585
R1469 B.n74 B.n73 585
R1470 B.n1179 B.n74 585
R1471 B.n1177 B.n1176 585
R1472 B.n1178 B.n1177 585
R1473 B.n1175 B.n79 585
R1474 B.n79 B.n78 585
R1475 B.n1174 B.n1173 585
R1476 B.n1173 B.n1172 585
R1477 B.n81 B.n80 585
R1478 B.n1171 B.n81 585
R1479 B.n1169 B.n1168 585
R1480 B.n1170 B.n1169 585
R1481 B.n1167 B.n86 585
R1482 B.n86 B.n85 585
R1483 B.n1166 B.n1165 585
R1484 B.n1165 B.n1164 585
R1485 B.n88 B.n87 585
R1486 B.n1163 B.n88 585
R1487 B.n1161 B.n1160 585
R1488 B.n1162 B.n1161 585
R1489 B.n1159 B.n93 585
R1490 B.n93 B.n92 585
R1491 B.n1158 B.n1157 585
R1492 B.n1157 B.n1156 585
R1493 B.n95 B.n94 585
R1494 B.n1155 B.n95 585
R1495 B.n1153 B.n1152 585
R1496 B.n1154 B.n1153 585
R1497 B.n1151 B.n100 585
R1498 B.n100 B.n99 585
R1499 B.n1150 B.n1149 585
R1500 B.n1149 B.n1148 585
R1501 B.n102 B.n101 585
R1502 B.n1147 B.n102 585
R1503 B.n1145 B.n1144 585
R1504 B.n1146 B.n1145 585
R1505 B.n1143 B.n106 585
R1506 B.n109 B.n106 585
R1507 B.n1142 B.n1141 585
R1508 B.n1141 B.n1140 585
R1509 B.n108 B.n107 585
R1510 B.n1139 B.n108 585
R1511 B.n1137 B.n1136 585
R1512 B.n1138 B.n1137 585
R1513 B.n1135 B.n114 585
R1514 B.n114 B.n113 585
R1515 B.n1134 B.n1133 585
R1516 B.n1133 B.n1132 585
R1517 B.n116 B.n115 585
R1518 B.n1131 B.n116 585
R1519 B.n1129 B.n1128 585
R1520 B.n1130 B.n1129 585
R1521 B.n1127 B.n121 585
R1522 B.n121 B.n120 585
R1523 B.n1126 B.n1125 585
R1524 B.n1125 B.n1124 585
R1525 B.n123 B.n122 585
R1526 B.n1123 B.n123 585
R1527 B.n1121 B.n1120 585
R1528 B.n1122 B.n1121 585
R1529 B.n1119 B.n128 585
R1530 B.n128 B.n127 585
R1531 B.n1118 B.n1117 585
R1532 B.n1117 B.n1116 585
R1533 B.n130 B.n129 585
R1534 B.n1115 B.n130 585
R1535 B.n1113 B.n1112 585
R1536 B.n1114 B.n1113 585
R1537 B.n1111 B.n134 585
R1538 B.n137 B.n134 585
R1539 B.n1110 B.n1109 585
R1540 B.n1109 B.n1108 585
R1541 B.n136 B.n135 585
R1542 B.n1107 B.n136 585
R1543 B.n1105 B.n1104 585
R1544 B.n1106 B.n1105 585
R1545 B.n1103 B.n142 585
R1546 B.n142 B.n141 585
R1547 B.n1102 B.n1101 585
R1548 B.n1101 B.n1100 585
R1549 B.n144 B.n143 585
R1550 B.n1099 B.n144 585
R1551 B.n1097 B.n1096 585
R1552 B.n1098 B.n1097 585
R1553 B.n1095 B.n149 585
R1554 B.n149 B.n148 585
R1555 B.n1094 B.n1093 585
R1556 B.n1093 B.n1092 585
R1557 B.n1262 B.n1261 585
R1558 B.n1261 B.n1260 585
R1559 B.n731 B.n520 545.355
R1560 B.n1093 B.n151 545.355
R1561 B.n729 B.n522 545.355
R1562 B.n1090 B.n152 545.355
R1563 B.n541 B.t20 331.817
R1564 B.n194 B.t15 331.817
R1565 B.n547 B.t23 331.817
R1566 B.n196 B.t12 331.817
R1567 B.n541 B.t17 270.212
R1568 B.n547 B.t21 270.212
R1569 B.n196 B.t10 270.212
R1570 B.n194 B.t14 270.212
R1571 B.n1091 B.n192 256.663
R1572 B.n1091 B.n191 256.663
R1573 B.n1091 B.n190 256.663
R1574 B.n1091 B.n189 256.663
R1575 B.n1091 B.n188 256.663
R1576 B.n1091 B.n187 256.663
R1577 B.n1091 B.n186 256.663
R1578 B.n1091 B.n185 256.663
R1579 B.n1091 B.n184 256.663
R1580 B.n1091 B.n183 256.663
R1581 B.n1091 B.n182 256.663
R1582 B.n1091 B.n181 256.663
R1583 B.n1091 B.n180 256.663
R1584 B.n1091 B.n179 256.663
R1585 B.n1091 B.n178 256.663
R1586 B.n1091 B.n177 256.663
R1587 B.n1091 B.n176 256.663
R1588 B.n1091 B.n175 256.663
R1589 B.n1091 B.n174 256.663
R1590 B.n1091 B.n173 256.663
R1591 B.n1091 B.n172 256.663
R1592 B.n1091 B.n171 256.663
R1593 B.n1091 B.n170 256.663
R1594 B.n1091 B.n169 256.663
R1595 B.n1091 B.n168 256.663
R1596 B.n1091 B.n167 256.663
R1597 B.n1091 B.n166 256.663
R1598 B.n1091 B.n165 256.663
R1599 B.n1091 B.n164 256.663
R1600 B.n1091 B.n163 256.663
R1601 B.n1091 B.n162 256.663
R1602 B.n1091 B.n161 256.663
R1603 B.n1091 B.n160 256.663
R1604 B.n1091 B.n159 256.663
R1605 B.n1091 B.n158 256.663
R1606 B.n1091 B.n157 256.663
R1607 B.n1091 B.n156 256.663
R1608 B.n1091 B.n155 256.663
R1609 B.n1091 B.n154 256.663
R1610 B.n1091 B.n153 256.663
R1611 B.n567 B.n521 256.663
R1612 B.n570 B.n521 256.663
R1613 B.n576 B.n521 256.663
R1614 B.n578 B.n521 256.663
R1615 B.n584 B.n521 256.663
R1616 B.n586 B.n521 256.663
R1617 B.n592 B.n521 256.663
R1618 B.n594 B.n521 256.663
R1619 B.n600 B.n521 256.663
R1620 B.n602 B.n521 256.663
R1621 B.n608 B.n521 256.663
R1622 B.n610 B.n521 256.663
R1623 B.n616 B.n521 256.663
R1624 B.n618 B.n521 256.663
R1625 B.n624 B.n521 256.663
R1626 B.n626 B.n521 256.663
R1627 B.n632 B.n521 256.663
R1628 B.n634 B.n521 256.663
R1629 B.n641 B.n521 256.663
R1630 B.n643 B.n521 256.663
R1631 B.n649 B.n521 256.663
R1632 B.n651 B.n521 256.663
R1633 B.n658 B.n521 256.663
R1634 B.n660 B.n521 256.663
R1635 B.n666 B.n521 256.663
R1636 B.n668 B.n521 256.663
R1637 B.n674 B.n521 256.663
R1638 B.n676 B.n521 256.663
R1639 B.n682 B.n521 256.663
R1640 B.n684 B.n521 256.663
R1641 B.n690 B.n521 256.663
R1642 B.n692 B.n521 256.663
R1643 B.n698 B.n521 256.663
R1644 B.n700 B.n521 256.663
R1645 B.n706 B.n521 256.663
R1646 B.n708 B.n521 256.663
R1647 B.n714 B.n521 256.663
R1648 B.n716 B.n521 256.663
R1649 B.n722 B.n521 256.663
R1650 B.n724 B.n521 256.663
R1651 B.n542 B.t19 248.23
R1652 B.n195 B.t16 248.23
R1653 B.n548 B.t22 248.228
R1654 B.n197 B.t13 248.228
R1655 B.n731 B.n518 163.367
R1656 B.n735 B.n518 163.367
R1657 B.n735 B.n512 163.367
R1658 B.n743 B.n512 163.367
R1659 B.n743 B.n510 163.367
R1660 B.n747 B.n510 163.367
R1661 B.n747 B.n504 163.367
R1662 B.n756 B.n504 163.367
R1663 B.n756 B.n502 163.367
R1664 B.n760 B.n502 163.367
R1665 B.n760 B.n497 163.367
R1666 B.n768 B.n497 163.367
R1667 B.n768 B.n495 163.367
R1668 B.n772 B.n495 163.367
R1669 B.n772 B.n489 163.367
R1670 B.n780 B.n489 163.367
R1671 B.n780 B.n487 163.367
R1672 B.n784 B.n487 163.367
R1673 B.n784 B.n481 163.367
R1674 B.n792 B.n481 163.367
R1675 B.n792 B.n479 163.367
R1676 B.n796 B.n479 163.367
R1677 B.n796 B.n473 163.367
R1678 B.n805 B.n473 163.367
R1679 B.n805 B.n471 163.367
R1680 B.n809 B.n471 163.367
R1681 B.n809 B.n466 163.367
R1682 B.n817 B.n466 163.367
R1683 B.n817 B.n464 163.367
R1684 B.n821 B.n464 163.367
R1685 B.n821 B.n458 163.367
R1686 B.n829 B.n458 163.367
R1687 B.n829 B.n456 163.367
R1688 B.n833 B.n456 163.367
R1689 B.n833 B.n450 163.367
R1690 B.n841 B.n450 163.367
R1691 B.n841 B.n448 163.367
R1692 B.n845 B.n448 163.367
R1693 B.n845 B.n442 163.367
R1694 B.n853 B.n442 163.367
R1695 B.n853 B.n440 163.367
R1696 B.n857 B.n440 163.367
R1697 B.n857 B.n434 163.367
R1698 B.n865 B.n434 163.367
R1699 B.n865 B.n432 163.367
R1700 B.n869 B.n432 163.367
R1701 B.n869 B.n426 163.367
R1702 B.n877 B.n426 163.367
R1703 B.n877 B.n424 163.367
R1704 B.n881 B.n424 163.367
R1705 B.n881 B.n418 163.367
R1706 B.n889 B.n418 163.367
R1707 B.n889 B.n416 163.367
R1708 B.n893 B.n416 163.367
R1709 B.n893 B.n410 163.367
R1710 B.n901 B.n410 163.367
R1711 B.n901 B.n408 163.367
R1712 B.n905 B.n408 163.367
R1713 B.n905 B.n402 163.367
R1714 B.n913 B.n402 163.367
R1715 B.n913 B.n400 163.367
R1716 B.n917 B.n400 163.367
R1717 B.n917 B.n394 163.367
R1718 B.n925 B.n394 163.367
R1719 B.n925 B.n392 163.367
R1720 B.n929 B.n392 163.367
R1721 B.n929 B.n386 163.367
R1722 B.n937 B.n386 163.367
R1723 B.n937 B.n384 163.367
R1724 B.n941 B.n384 163.367
R1725 B.n941 B.n378 163.367
R1726 B.n949 B.n378 163.367
R1727 B.n949 B.n376 163.367
R1728 B.n953 B.n376 163.367
R1729 B.n953 B.n370 163.367
R1730 B.n961 B.n370 163.367
R1731 B.n961 B.n368 163.367
R1732 B.n965 B.n368 163.367
R1733 B.n965 B.n362 163.367
R1734 B.n974 B.n362 163.367
R1735 B.n974 B.n360 163.367
R1736 B.n978 B.n360 163.367
R1737 B.n978 B.n2 163.367
R1738 B.n1261 B.n2 163.367
R1739 B.n1261 B.n3 163.367
R1740 B.n1257 B.n3 163.367
R1741 B.n1257 B.n9 163.367
R1742 B.n1253 B.n9 163.367
R1743 B.n1253 B.n11 163.367
R1744 B.n1249 B.n11 163.367
R1745 B.n1249 B.n16 163.367
R1746 B.n1245 B.n16 163.367
R1747 B.n1245 B.n18 163.367
R1748 B.n1241 B.n18 163.367
R1749 B.n1241 B.n23 163.367
R1750 B.n1237 B.n23 163.367
R1751 B.n1237 B.n25 163.367
R1752 B.n1233 B.n25 163.367
R1753 B.n1233 B.n30 163.367
R1754 B.n1229 B.n30 163.367
R1755 B.n1229 B.n32 163.367
R1756 B.n1225 B.n32 163.367
R1757 B.n1225 B.n37 163.367
R1758 B.n1221 B.n37 163.367
R1759 B.n1221 B.n39 163.367
R1760 B.n1217 B.n39 163.367
R1761 B.n1217 B.n44 163.367
R1762 B.n1213 B.n44 163.367
R1763 B.n1213 B.n46 163.367
R1764 B.n1209 B.n46 163.367
R1765 B.n1209 B.n51 163.367
R1766 B.n1205 B.n51 163.367
R1767 B.n1205 B.n53 163.367
R1768 B.n1201 B.n53 163.367
R1769 B.n1201 B.n58 163.367
R1770 B.n1197 B.n58 163.367
R1771 B.n1197 B.n60 163.367
R1772 B.n1193 B.n60 163.367
R1773 B.n1193 B.n65 163.367
R1774 B.n1189 B.n65 163.367
R1775 B.n1189 B.n67 163.367
R1776 B.n1185 B.n67 163.367
R1777 B.n1185 B.n72 163.367
R1778 B.n1181 B.n72 163.367
R1779 B.n1181 B.n74 163.367
R1780 B.n1177 B.n74 163.367
R1781 B.n1177 B.n79 163.367
R1782 B.n1173 B.n79 163.367
R1783 B.n1173 B.n81 163.367
R1784 B.n1169 B.n81 163.367
R1785 B.n1169 B.n86 163.367
R1786 B.n1165 B.n86 163.367
R1787 B.n1165 B.n88 163.367
R1788 B.n1161 B.n88 163.367
R1789 B.n1161 B.n93 163.367
R1790 B.n1157 B.n93 163.367
R1791 B.n1157 B.n95 163.367
R1792 B.n1153 B.n95 163.367
R1793 B.n1153 B.n100 163.367
R1794 B.n1149 B.n100 163.367
R1795 B.n1149 B.n102 163.367
R1796 B.n1145 B.n102 163.367
R1797 B.n1145 B.n106 163.367
R1798 B.n1141 B.n106 163.367
R1799 B.n1141 B.n108 163.367
R1800 B.n1137 B.n108 163.367
R1801 B.n1137 B.n114 163.367
R1802 B.n1133 B.n114 163.367
R1803 B.n1133 B.n116 163.367
R1804 B.n1129 B.n116 163.367
R1805 B.n1129 B.n121 163.367
R1806 B.n1125 B.n121 163.367
R1807 B.n1125 B.n123 163.367
R1808 B.n1121 B.n123 163.367
R1809 B.n1121 B.n128 163.367
R1810 B.n1117 B.n128 163.367
R1811 B.n1117 B.n130 163.367
R1812 B.n1113 B.n130 163.367
R1813 B.n1113 B.n134 163.367
R1814 B.n1109 B.n134 163.367
R1815 B.n1109 B.n136 163.367
R1816 B.n1105 B.n136 163.367
R1817 B.n1105 B.n142 163.367
R1818 B.n1101 B.n142 163.367
R1819 B.n1101 B.n144 163.367
R1820 B.n1097 B.n144 163.367
R1821 B.n1097 B.n149 163.367
R1822 B.n1093 B.n149 163.367
R1823 B.n569 B.n568 163.367
R1824 B.n571 B.n569 163.367
R1825 B.n575 B.n564 163.367
R1826 B.n579 B.n577 163.367
R1827 B.n583 B.n562 163.367
R1828 B.n587 B.n585 163.367
R1829 B.n591 B.n560 163.367
R1830 B.n595 B.n593 163.367
R1831 B.n599 B.n558 163.367
R1832 B.n603 B.n601 163.367
R1833 B.n607 B.n556 163.367
R1834 B.n611 B.n609 163.367
R1835 B.n615 B.n554 163.367
R1836 B.n619 B.n617 163.367
R1837 B.n623 B.n552 163.367
R1838 B.n627 B.n625 163.367
R1839 B.n631 B.n550 163.367
R1840 B.n635 B.n633 163.367
R1841 B.n640 B.n546 163.367
R1842 B.n644 B.n642 163.367
R1843 B.n648 B.n544 163.367
R1844 B.n652 B.n650 163.367
R1845 B.n657 B.n540 163.367
R1846 B.n661 B.n659 163.367
R1847 B.n665 B.n538 163.367
R1848 B.n669 B.n667 163.367
R1849 B.n673 B.n536 163.367
R1850 B.n677 B.n675 163.367
R1851 B.n681 B.n534 163.367
R1852 B.n685 B.n683 163.367
R1853 B.n689 B.n532 163.367
R1854 B.n693 B.n691 163.367
R1855 B.n697 B.n530 163.367
R1856 B.n701 B.n699 163.367
R1857 B.n705 B.n528 163.367
R1858 B.n709 B.n707 163.367
R1859 B.n713 B.n526 163.367
R1860 B.n717 B.n715 163.367
R1861 B.n721 B.n524 163.367
R1862 B.n725 B.n723 163.367
R1863 B.n729 B.n516 163.367
R1864 B.n737 B.n516 163.367
R1865 B.n737 B.n514 163.367
R1866 B.n741 B.n514 163.367
R1867 B.n741 B.n508 163.367
R1868 B.n749 B.n508 163.367
R1869 B.n749 B.n506 163.367
R1870 B.n753 B.n506 163.367
R1871 B.n753 B.n501 163.367
R1872 B.n762 B.n501 163.367
R1873 B.n762 B.n499 163.367
R1874 B.n766 B.n499 163.367
R1875 B.n766 B.n493 163.367
R1876 B.n774 B.n493 163.367
R1877 B.n774 B.n491 163.367
R1878 B.n778 B.n491 163.367
R1879 B.n778 B.n485 163.367
R1880 B.n786 B.n485 163.367
R1881 B.n786 B.n483 163.367
R1882 B.n790 B.n483 163.367
R1883 B.n790 B.n477 163.367
R1884 B.n798 B.n477 163.367
R1885 B.n798 B.n475 163.367
R1886 B.n802 B.n475 163.367
R1887 B.n802 B.n470 163.367
R1888 B.n811 B.n470 163.367
R1889 B.n811 B.n468 163.367
R1890 B.n815 B.n468 163.367
R1891 B.n815 B.n462 163.367
R1892 B.n823 B.n462 163.367
R1893 B.n823 B.n460 163.367
R1894 B.n827 B.n460 163.367
R1895 B.n827 B.n454 163.367
R1896 B.n835 B.n454 163.367
R1897 B.n835 B.n452 163.367
R1898 B.n839 B.n452 163.367
R1899 B.n839 B.n446 163.367
R1900 B.n847 B.n446 163.367
R1901 B.n847 B.n444 163.367
R1902 B.n851 B.n444 163.367
R1903 B.n851 B.n438 163.367
R1904 B.n859 B.n438 163.367
R1905 B.n859 B.n436 163.367
R1906 B.n863 B.n436 163.367
R1907 B.n863 B.n430 163.367
R1908 B.n871 B.n430 163.367
R1909 B.n871 B.n428 163.367
R1910 B.n875 B.n428 163.367
R1911 B.n875 B.n422 163.367
R1912 B.n883 B.n422 163.367
R1913 B.n883 B.n420 163.367
R1914 B.n887 B.n420 163.367
R1915 B.n887 B.n414 163.367
R1916 B.n895 B.n414 163.367
R1917 B.n895 B.n412 163.367
R1918 B.n899 B.n412 163.367
R1919 B.n899 B.n406 163.367
R1920 B.n907 B.n406 163.367
R1921 B.n907 B.n404 163.367
R1922 B.n911 B.n404 163.367
R1923 B.n911 B.n397 163.367
R1924 B.n919 B.n397 163.367
R1925 B.n919 B.n395 163.367
R1926 B.n923 B.n395 163.367
R1927 B.n923 B.n390 163.367
R1928 B.n931 B.n390 163.367
R1929 B.n931 B.n388 163.367
R1930 B.n935 B.n388 163.367
R1931 B.n935 B.n382 163.367
R1932 B.n943 B.n382 163.367
R1933 B.n943 B.n380 163.367
R1934 B.n947 B.n380 163.367
R1935 B.n947 B.n374 163.367
R1936 B.n955 B.n374 163.367
R1937 B.n955 B.n372 163.367
R1938 B.n959 B.n372 163.367
R1939 B.n959 B.n366 163.367
R1940 B.n967 B.n366 163.367
R1941 B.n967 B.n364 163.367
R1942 B.n972 B.n364 163.367
R1943 B.n972 B.n358 163.367
R1944 B.n980 B.n358 163.367
R1945 B.n981 B.n980 163.367
R1946 B.n981 B.n5 163.367
R1947 B.n6 B.n5 163.367
R1948 B.n7 B.n6 163.367
R1949 B.n986 B.n7 163.367
R1950 B.n986 B.n12 163.367
R1951 B.n13 B.n12 163.367
R1952 B.n14 B.n13 163.367
R1953 B.n991 B.n14 163.367
R1954 B.n991 B.n19 163.367
R1955 B.n20 B.n19 163.367
R1956 B.n21 B.n20 163.367
R1957 B.n996 B.n21 163.367
R1958 B.n996 B.n26 163.367
R1959 B.n27 B.n26 163.367
R1960 B.n28 B.n27 163.367
R1961 B.n1001 B.n28 163.367
R1962 B.n1001 B.n33 163.367
R1963 B.n34 B.n33 163.367
R1964 B.n35 B.n34 163.367
R1965 B.n1006 B.n35 163.367
R1966 B.n1006 B.n40 163.367
R1967 B.n41 B.n40 163.367
R1968 B.n42 B.n41 163.367
R1969 B.n1011 B.n42 163.367
R1970 B.n1011 B.n47 163.367
R1971 B.n48 B.n47 163.367
R1972 B.n49 B.n48 163.367
R1973 B.n1016 B.n49 163.367
R1974 B.n1016 B.n54 163.367
R1975 B.n55 B.n54 163.367
R1976 B.n56 B.n55 163.367
R1977 B.n1021 B.n56 163.367
R1978 B.n1021 B.n61 163.367
R1979 B.n62 B.n61 163.367
R1980 B.n63 B.n62 163.367
R1981 B.n1026 B.n63 163.367
R1982 B.n1026 B.n68 163.367
R1983 B.n69 B.n68 163.367
R1984 B.n70 B.n69 163.367
R1985 B.n1031 B.n70 163.367
R1986 B.n1031 B.n75 163.367
R1987 B.n76 B.n75 163.367
R1988 B.n77 B.n76 163.367
R1989 B.n1036 B.n77 163.367
R1990 B.n1036 B.n82 163.367
R1991 B.n83 B.n82 163.367
R1992 B.n84 B.n83 163.367
R1993 B.n1041 B.n84 163.367
R1994 B.n1041 B.n89 163.367
R1995 B.n90 B.n89 163.367
R1996 B.n91 B.n90 163.367
R1997 B.n1046 B.n91 163.367
R1998 B.n1046 B.n96 163.367
R1999 B.n97 B.n96 163.367
R2000 B.n98 B.n97 163.367
R2001 B.n1051 B.n98 163.367
R2002 B.n1051 B.n103 163.367
R2003 B.n104 B.n103 163.367
R2004 B.n105 B.n104 163.367
R2005 B.n1056 B.n105 163.367
R2006 B.n1056 B.n110 163.367
R2007 B.n111 B.n110 163.367
R2008 B.n112 B.n111 163.367
R2009 B.n1061 B.n112 163.367
R2010 B.n1061 B.n117 163.367
R2011 B.n118 B.n117 163.367
R2012 B.n119 B.n118 163.367
R2013 B.n1066 B.n119 163.367
R2014 B.n1066 B.n124 163.367
R2015 B.n125 B.n124 163.367
R2016 B.n126 B.n125 163.367
R2017 B.n1071 B.n126 163.367
R2018 B.n1071 B.n131 163.367
R2019 B.n132 B.n131 163.367
R2020 B.n133 B.n132 163.367
R2021 B.n1076 B.n133 163.367
R2022 B.n1076 B.n138 163.367
R2023 B.n139 B.n138 163.367
R2024 B.n140 B.n139 163.367
R2025 B.n1081 B.n140 163.367
R2026 B.n1081 B.n145 163.367
R2027 B.n146 B.n145 163.367
R2028 B.n147 B.n146 163.367
R2029 B.n1086 B.n147 163.367
R2030 B.n1086 B.n152 163.367
R2031 B.n201 B.n200 163.367
R2032 B.n205 B.n204 163.367
R2033 B.n209 B.n208 163.367
R2034 B.n213 B.n212 163.367
R2035 B.n217 B.n216 163.367
R2036 B.n221 B.n220 163.367
R2037 B.n225 B.n224 163.367
R2038 B.n229 B.n228 163.367
R2039 B.n233 B.n232 163.367
R2040 B.n237 B.n236 163.367
R2041 B.n241 B.n240 163.367
R2042 B.n245 B.n244 163.367
R2043 B.n249 B.n248 163.367
R2044 B.n253 B.n252 163.367
R2045 B.n257 B.n256 163.367
R2046 B.n261 B.n260 163.367
R2047 B.n265 B.n264 163.367
R2048 B.n269 B.n268 163.367
R2049 B.n273 B.n272 163.367
R2050 B.n277 B.n276 163.367
R2051 B.n281 B.n280 163.367
R2052 B.n285 B.n284 163.367
R2053 B.n290 B.n289 163.367
R2054 B.n294 B.n293 163.367
R2055 B.n298 B.n297 163.367
R2056 B.n302 B.n301 163.367
R2057 B.n306 B.n305 163.367
R2058 B.n310 B.n309 163.367
R2059 B.n314 B.n313 163.367
R2060 B.n318 B.n317 163.367
R2061 B.n322 B.n321 163.367
R2062 B.n326 B.n325 163.367
R2063 B.n330 B.n329 163.367
R2064 B.n334 B.n333 163.367
R2065 B.n338 B.n337 163.367
R2066 B.n342 B.n341 163.367
R2067 B.n346 B.n345 163.367
R2068 B.n350 B.n349 163.367
R2069 B.n354 B.n353 163.367
R2070 B.n1090 B.n193 163.367
R2071 B.n730 B.n521 97.0276
R2072 B.n1092 B.n1091 97.0276
R2073 B.n542 B.n541 83.5884
R2074 B.n548 B.n547 83.5884
R2075 B.n197 B.n196 83.5884
R2076 B.n195 B.n194 83.5884
R2077 B.n567 B.n520 71.676
R2078 B.n571 B.n570 71.676
R2079 B.n576 B.n575 71.676
R2080 B.n579 B.n578 71.676
R2081 B.n584 B.n583 71.676
R2082 B.n587 B.n586 71.676
R2083 B.n592 B.n591 71.676
R2084 B.n595 B.n594 71.676
R2085 B.n600 B.n599 71.676
R2086 B.n603 B.n602 71.676
R2087 B.n608 B.n607 71.676
R2088 B.n611 B.n610 71.676
R2089 B.n616 B.n615 71.676
R2090 B.n619 B.n618 71.676
R2091 B.n624 B.n623 71.676
R2092 B.n627 B.n626 71.676
R2093 B.n632 B.n631 71.676
R2094 B.n635 B.n634 71.676
R2095 B.n641 B.n640 71.676
R2096 B.n644 B.n643 71.676
R2097 B.n649 B.n648 71.676
R2098 B.n652 B.n651 71.676
R2099 B.n658 B.n657 71.676
R2100 B.n661 B.n660 71.676
R2101 B.n666 B.n665 71.676
R2102 B.n669 B.n668 71.676
R2103 B.n674 B.n673 71.676
R2104 B.n677 B.n676 71.676
R2105 B.n682 B.n681 71.676
R2106 B.n685 B.n684 71.676
R2107 B.n690 B.n689 71.676
R2108 B.n693 B.n692 71.676
R2109 B.n698 B.n697 71.676
R2110 B.n701 B.n700 71.676
R2111 B.n706 B.n705 71.676
R2112 B.n709 B.n708 71.676
R2113 B.n714 B.n713 71.676
R2114 B.n717 B.n716 71.676
R2115 B.n722 B.n721 71.676
R2116 B.n725 B.n724 71.676
R2117 B.n153 B.n151 71.676
R2118 B.n201 B.n154 71.676
R2119 B.n205 B.n155 71.676
R2120 B.n209 B.n156 71.676
R2121 B.n213 B.n157 71.676
R2122 B.n217 B.n158 71.676
R2123 B.n221 B.n159 71.676
R2124 B.n225 B.n160 71.676
R2125 B.n229 B.n161 71.676
R2126 B.n233 B.n162 71.676
R2127 B.n237 B.n163 71.676
R2128 B.n241 B.n164 71.676
R2129 B.n245 B.n165 71.676
R2130 B.n249 B.n166 71.676
R2131 B.n253 B.n167 71.676
R2132 B.n257 B.n168 71.676
R2133 B.n261 B.n169 71.676
R2134 B.n265 B.n170 71.676
R2135 B.n269 B.n171 71.676
R2136 B.n273 B.n172 71.676
R2137 B.n277 B.n173 71.676
R2138 B.n281 B.n174 71.676
R2139 B.n285 B.n175 71.676
R2140 B.n290 B.n176 71.676
R2141 B.n294 B.n177 71.676
R2142 B.n298 B.n178 71.676
R2143 B.n302 B.n179 71.676
R2144 B.n306 B.n180 71.676
R2145 B.n310 B.n181 71.676
R2146 B.n314 B.n182 71.676
R2147 B.n318 B.n183 71.676
R2148 B.n322 B.n184 71.676
R2149 B.n326 B.n185 71.676
R2150 B.n330 B.n186 71.676
R2151 B.n334 B.n187 71.676
R2152 B.n338 B.n188 71.676
R2153 B.n342 B.n189 71.676
R2154 B.n346 B.n190 71.676
R2155 B.n350 B.n191 71.676
R2156 B.n354 B.n192 71.676
R2157 B.n193 B.n192 71.676
R2158 B.n353 B.n191 71.676
R2159 B.n349 B.n190 71.676
R2160 B.n345 B.n189 71.676
R2161 B.n341 B.n188 71.676
R2162 B.n337 B.n187 71.676
R2163 B.n333 B.n186 71.676
R2164 B.n329 B.n185 71.676
R2165 B.n325 B.n184 71.676
R2166 B.n321 B.n183 71.676
R2167 B.n317 B.n182 71.676
R2168 B.n313 B.n181 71.676
R2169 B.n309 B.n180 71.676
R2170 B.n305 B.n179 71.676
R2171 B.n301 B.n178 71.676
R2172 B.n297 B.n177 71.676
R2173 B.n293 B.n176 71.676
R2174 B.n289 B.n175 71.676
R2175 B.n284 B.n174 71.676
R2176 B.n280 B.n173 71.676
R2177 B.n276 B.n172 71.676
R2178 B.n272 B.n171 71.676
R2179 B.n268 B.n170 71.676
R2180 B.n264 B.n169 71.676
R2181 B.n260 B.n168 71.676
R2182 B.n256 B.n167 71.676
R2183 B.n252 B.n166 71.676
R2184 B.n248 B.n165 71.676
R2185 B.n244 B.n164 71.676
R2186 B.n240 B.n163 71.676
R2187 B.n236 B.n162 71.676
R2188 B.n232 B.n161 71.676
R2189 B.n228 B.n160 71.676
R2190 B.n224 B.n159 71.676
R2191 B.n220 B.n158 71.676
R2192 B.n216 B.n157 71.676
R2193 B.n212 B.n156 71.676
R2194 B.n208 B.n155 71.676
R2195 B.n204 B.n154 71.676
R2196 B.n200 B.n153 71.676
R2197 B.n568 B.n567 71.676
R2198 B.n570 B.n564 71.676
R2199 B.n577 B.n576 71.676
R2200 B.n578 B.n562 71.676
R2201 B.n585 B.n584 71.676
R2202 B.n586 B.n560 71.676
R2203 B.n593 B.n592 71.676
R2204 B.n594 B.n558 71.676
R2205 B.n601 B.n600 71.676
R2206 B.n602 B.n556 71.676
R2207 B.n609 B.n608 71.676
R2208 B.n610 B.n554 71.676
R2209 B.n617 B.n616 71.676
R2210 B.n618 B.n552 71.676
R2211 B.n625 B.n624 71.676
R2212 B.n626 B.n550 71.676
R2213 B.n633 B.n632 71.676
R2214 B.n634 B.n546 71.676
R2215 B.n642 B.n641 71.676
R2216 B.n643 B.n544 71.676
R2217 B.n650 B.n649 71.676
R2218 B.n651 B.n540 71.676
R2219 B.n659 B.n658 71.676
R2220 B.n660 B.n538 71.676
R2221 B.n667 B.n666 71.676
R2222 B.n668 B.n536 71.676
R2223 B.n675 B.n674 71.676
R2224 B.n676 B.n534 71.676
R2225 B.n683 B.n682 71.676
R2226 B.n684 B.n532 71.676
R2227 B.n691 B.n690 71.676
R2228 B.n692 B.n530 71.676
R2229 B.n699 B.n698 71.676
R2230 B.n700 B.n528 71.676
R2231 B.n707 B.n706 71.676
R2232 B.n708 B.n526 71.676
R2233 B.n715 B.n714 71.676
R2234 B.n716 B.n524 71.676
R2235 B.n723 B.n722 71.676
R2236 B.n724 B.n522 71.676
R2237 B.n655 B.n542 59.5399
R2238 B.n637 B.n548 59.5399
R2239 B.n198 B.n197 59.5399
R2240 B.n287 B.n195 59.5399
R2241 B.n730 B.n517 48.8734
R2242 B.n736 B.n517 48.8734
R2243 B.n736 B.n513 48.8734
R2244 B.n742 B.n513 48.8734
R2245 B.n742 B.n509 48.8734
R2246 B.n748 B.n509 48.8734
R2247 B.n748 B.n505 48.8734
R2248 B.n755 B.n505 48.8734
R2249 B.n755 B.n754 48.8734
R2250 B.n761 B.n498 48.8734
R2251 B.n767 B.n498 48.8734
R2252 B.n767 B.n494 48.8734
R2253 B.n773 B.n494 48.8734
R2254 B.n773 B.n490 48.8734
R2255 B.n779 B.n490 48.8734
R2256 B.n779 B.n486 48.8734
R2257 B.n785 B.n486 48.8734
R2258 B.n785 B.n482 48.8734
R2259 B.n791 B.n482 48.8734
R2260 B.n791 B.n478 48.8734
R2261 B.n797 B.n478 48.8734
R2262 B.n797 B.n474 48.8734
R2263 B.n804 B.n474 48.8734
R2264 B.n804 B.n803 48.8734
R2265 B.n810 B.n467 48.8734
R2266 B.n816 B.n467 48.8734
R2267 B.n816 B.n463 48.8734
R2268 B.n822 B.n463 48.8734
R2269 B.n822 B.n459 48.8734
R2270 B.n828 B.n459 48.8734
R2271 B.n828 B.n455 48.8734
R2272 B.n834 B.n455 48.8734
R2273 B.n834 B.n451 48.8734
R2274 B.n840 B.n451 48.8734
R2275 B.n840 B.n447 48.8734
R2276 B.n846 B.n447 48.8734
R2277 B.n852 B.n443 48.8734
R2278 B.n852 B.n439 48.8734
R2279 B.n858 B.n439 48.8734
R2280 B.n858 B.n435 48.8734
R2281 B.n864 B.n435 48.8734
R2282 B.n864 B.n431 48.8734
R2283 B.n870 B.n431 48.8734
R2284 B.n870 B.n427 48.8734
R2285 B.n876 B.n427 48.8734
R2286 B.n876 B.n423 48.8734
R2287 B.n882 B.n423 48.8734
R2288 B.n888 B.n419 48.8734
R2289 B.n888 B.n415 48.8734
R2290 B.n894 B.n415 48.8734
R2291 B.n894 B.n411 48.8734
R2292 B.n900 B.n411 48.8734
R2293 B.n900 B.n407 48.8734
R2294 B.n906 B.n407 48.8734
R2295 B.n906 B.n403 48.8734
R2296 B.n912 B.n403 48.8734
R2297 B.n912 B.n398 48.8734
R2298 B.n918 B.n398 48.8734
R2299 B.n918 B.n399 48.8734
R2300 B.n924 B.n391 48.8734
R2301 B.n930 B.n391 48.8734
R2302 B.n930 B.n387 48.8734
R2303 B.n936 B.n387 48.8734
R2304 B.n936 B.n383 48.8734
R2305 B.n942 B.n383 48.8734
R2306 B.n942 B.n379 48.8734
R2307 B.n948 B.n379 48.8734
R2308 B.n948 B.n375 48.8734
R2309 B.n954 B.n375 48.8734
R2310 B.n954 B.n371 48.8734
R2311 B.n960 B.n371 48.8734
R2312 B.n966 B.n367 48.8734
R2313 B.n966 B.n363 48.8734
R2314 B.n973 B.n363 48.8734
R2315 B.n973 B.n359 48.8734
R2316 B.n979 B.n359 48.8734
R2317 B.n979 B.n4 48.8734
R2318 B.n1260 B.n4 48.8734
R2319 B.n1260 B.n1259 48.8734
R2320 B.n1259 B.n1258 48.8734
R2321 B.n1258 B.n8 48.8734
R2322 B.n1252 B.n8 48.8734
R2323 B.n1252 B.n1251 48.8734
R2324 B.n1251 B.n1250 48.8734
R2325 B.n1250 B.n15 48.8734
R2326 B.n1244 B.n1243 48.8734
R2327 B.n1243 B.n1242 48.8734
R2328 B.n1242 B.n22 48.8734
R2329 B.n1236 B.n22 48.8734
R2330 B.n1236 B.n1235 48.8734
R2331 B.n1235 B.n1234 48.8734
R2332 B.n1234 B.n29 48.8734
R2333 B.n1228 B.n29 48.8734
R2334 B.n1228 B.n1227 48.8734
R2335 B.n1227 B.n1226 48.8734
R2336 B.n1226 B.n36 48.8734
R2337 B.n1220 B.n36 48.8734
R2338 B.n1219 B.n1218 48.8734
R2339 B.n1218 B.n43 48.8734
R2340 B.n1212 B.n43 48.8734
R2341 B.n1212 B.n1211 48.8734
R2342 B.n1211 B.n1210 48.8734
R2343 B.n1210 B.n50 48.8734
R2344 B.n1204 B.n50 48.8734
R2345 B.n1204 B.n1203 48.8734
R2346 B.n1203 B.n1202 48.8734
R2347 B.n1202 B.n57 48.8734
R2348 B.n1196 B.n57 48.8734
R2349 B.n1196 B.n1195 48.8734
R2350 B.n1194 B.n64 48.8734
R2351 B.n1188 B.n64 48.8734
R2352 B.n1188 B.n1187 48.8734
R2353 B.n1187 B.n1186 48.8734
R2354 B.n1186 B.n71 48.8734
R2355 B.n1180 B.n71 48.8734
R2356 B.n1180 B.n1179 48.8734
R2357 B.n1179 B.n1178 48.8734
R2358 B.n1178 B.n78 48.8734
R2359 B.n1172 B.n78 48.8734
R2360 B.n1172 B.n1171 48.8734
R2361 B.n1170 B.n85 48.8734
R2362 B.n1164 B.n85 48.8734
R2363 B.n1164 B.n1163 48.8734
R2364 B.n1163 B.n1162 48.8734
R2365 B.n1162 B.n92 48.8734
R2366 B.n1156 B.n92 48.8734
R2367 B.n1156 B.n1155 48.8734
R2368 B.n1155 B.n1154 48.8734
R2369 B.n1154 B.n99 48.8734
R2370 B.n1148 B.n99 48.8734
R2371 B.n1148 B.n1147 48.8734
R2372 B.n1147 B.n1146 48.8734
R2373 B.n1140 B.n109 48.8734
R2374 B.n1140 B.n1139 48.8734
R2375 B.n1139 B.n1138 48.8734
R2376 B.n1138 B.n113 48.8734
R2377 B.n1132 B.n113 48.8734
R2378 B.n1132 B.n1131 48.8734
R2379 B.n1131 B.n1130 48.8734
R2380 B.n1130 B.n120 48.8734
R2381 B.n1124 B.n120 48.8734
R2382 B.n1124 B.n1123 48.8734
R2383 B.n1123 B.n1122 48.8734
R2384 B.n1122 B.n127 48.8734
R2385 B.n1116 B.n127 48.8734
R2386 B.n1116 B.n1115 48.8734
R2387 B.n1115 B.n1114 48.8734
R2388 B.n1108 B.n137 48.8734
R2389 B.n1108 B.n1107 48.8734
R2390 B.n1107 B.n1106 48.8734
R2391 B.n1106 B.n141 48.8734
R2392 B.n1100 B.n141 48.8734
R2393 B.n1100 B.n1099 48.8734
R2394 B.n1099 B.n1098 48.8734
R2395 B.n1098 B.n148 48.8734
R2396 B.n1092 B.n148 48.8734
R2397 B.t5 B.n443 47.436
R2398 B.n1171 B.t0 47.436
R2399 B.t7 B.n367 45.9985
R2400 B.t9 B.n15 45.9985
R2401 B.n1089 B.n1088 35.4346
R2402 B.n1094 B.n150 35.4346
R2403 B.n728 B.n727 35.4346
R2404 B.n732 B.n519 35.4346
R2405 B.n882 B.t1 34.499
R2406 B.t6 B.n1194 34.499
R2407 B.n810 B.t2 31.6242
R2408 B.n1146 B.t4 31.6242
R2409 B.n924 B.t3 30.1867
R2410 B.n1220 B.t8 30.1867
R2411 B.n761 B.t18 25.8744
R2412 B.n1114 B.t11 25.8744
R2413 B.n754 B.t18 22.9995
R2414 B.n137 B.t11 22.9995
R2415 B.n399 B.t3 18.6872
R2416 B.t8 B.n1219 18.6872
R2417 B B.n1262 18.0485
R2418 B.n803 B.t2 17.2498
R2419 B.n109 B.t4 17.2498
R2420 B.t1 B.n419 14.3749
R2421 B.n1195 B.t6 14.3749
R2422 B.n199 B.n150 10.6151
R2423 B.n202 B.n199 10.6151
R2424 B.n203 B.n202 10.6151
R2425 B.n206 B.n203 10.6151
R2426 B.n207 B.n206 10.6151
R2427 B.n210 B.n207 10.6151
R2428 B.n211 B.n210 10.6151
R2429 B.n214 B.n211 10.6151
R2430 B.n215 B.n214 10.6151
R2431 B.n218 B.n215 10.6151
R2432 B.n219 B.n218 10.6151
R2433 B.n222 B.n219 10.6151
R2434 B.n223 B.n222 10.6151
R2435 B.n226 B.n223 10.6151
R2436 B.n227 B.n226 10.6151
R2437 B.n230 B.n227 10.6151
R2438 B.n231 B.n230 10.6151
R2439 B.n234 B.n231 10.6151
R2440 B.n235 B.n234 10.6151
R2441 B.n238 B.n235 10.6151
R2442 B.n239 B.n238 10.6151
R2443 B.n242 B.n239 10.6151
R2444 B.n243 B.n242 10.6151
R2445 B.n246 B.n243 10.6151
R2446 B.n247 B.n246 10.6151
R2447 B.n250 B.n247 10.6151
R2448 B.n251 B.n250 10.6151
R2449 B.n254 B.n251 10.6151
R2450 B.n255 B.n254 10.6151
R2451 B.n258 B.n255 10.6151
R2452 B.n259 B.n258 10.6151
R2453 B.n262 B.n259 10.6151
R2454 B.n263 B.n262 10.6151
R2455 B.n266 B.n263 10.6151
R2456 B.n267 B.n266 10.6151
R2457 B.n271 B.n270 10.6151
R2458 B.n274 B.n271 10.6151
R2459 B.n275 B.n274 10.6151
R2460 B.n278 B.n275 10.6151
R2461 B.n279 B.n278 10.6151
R2462 B.n282 B.n279 10.6151
R2463 B.n283 B.n282 10.6151
R2464 B.n286 B.n283 10.6151
R2465 B.n291 B.n288 10.6151
R2466 B.n292 B.n291 10.6151
R2467 B.n295 B.n292 10.6151
R2468 B.n296 B.n295 10.6151
R2469 B.n299 B.n296 10.6151
R2470 B.n300 B.n299 10.6151
R2471 B.n303 B.n300 10.6151
R2472 B.n304 B.n303 10.6151
R2473 B.n307 B.n304 10.6151
R2474 B.n308 B.n307 10.6151
R2475 B.n311 B.n308 10.6151
R2476 B.n312 B.n311 10.6151
R2477 B.n315 B.n312 10.6151
R2478 B.n316 B.n315 10.6151
R2479 B.n319 B.n316 10.6151
R2480 B.n320 B.n319 10.6151
R2481 B.n323 B.n320 10.6151
R2482 B.n324 B.n323 10.6151
R2483 B.n327 B.n324 10.6151
R2484 B.n328 B.n327 10.6151
R2485 B.n331 B.n328 10.6151
R2486 B.n332 B.n331 10.6151
R2487 B.n335 B.n332 10.6151
R2488 B.n336 B.n335 10.6151
R2489 B.n339 B.n336 10.6151
R2490 B.n340 B.n339 10.6151
R2491 B.n343 B.n340 10.6151
R2492 B.n344 B.n343 10.6151
R2493 B.n347 B.n344 10.6151
R2494 B.n348 B.n347 10.6151
R2495 B.n351 B.n348 10.6151
R2496 B.n352 B.n351 10.6151
R2497 B.n355 B.n352 10.6151
R2498 B.n356 B.n355 10.6151
R2499 B.n1089 B.n356 10.6151
R2500 B.n728 B.n515 10.6151
R2501 B.n738 B.n515 10.6151
R2502 B.n739 B.n738 10.6151
R2503 B.n740 B.n739 10.6151
R2504 B.n740 B.n507 10.6151
R2505 B.n750 B.n507 10.6151
R2506 B.n751 B.n750 10.6151
R2507 B.n752 B.n751 10.6151
R2508 B.n752 B.n500 10.6151
R2509 B.n763 B.n500 10.6151
R2510 B.n764 B.n763 10.6151
R2511 B.n765 B.n764 10.6151
R2512 B.n765 B.n492 10.6151
R2513 B.n775 B.n492 10.6151
R2514 B.n776 B.n775 10.6151
R2515 B.n777 B.n776 10.6151
R2516 B.n777 B.n484 10.6151
R2517 B.n787 B.n484 10.6151
R2518 B.n788 B.n787 10.6151
R2519 B.n789 B.n788 10.6151
R2520 B.n789 B.n476 10.6151
R2521 B.n799 B.n476 10.6151
R2522 B.n800 B.n799 10.6151
R2523 B.n801 B.n800 10.6151
R2524 B.n801 B.n469 10.6151
R2525 B.n812 B.n469 10.6151
R2526 B.n813 B.n812 10.6151
R2527 B.n814 B.n813 10.6151
R2528 B.n814 B.n461 10.6151
R2529 B.n824 B.n461 10.6151
R2530 B.n825 B.n824 10.6151
R2531 B.n826 B.n825 10.6151
R2532 B.n826 B.n453 10.6151
R2533 B.n836 B.n453 10.6151
R2534 B.n837 B.n836 10.6151
R2535 B.n838 B.n837 10.6151
R2536 B.n838 B.n445 10.6151
R2537 B.n848 B.n445 10.6151
R2538 B.n849 B.n848 10.6151
R2539 B.n850 B.n849 10.6151
R2540 B.n850 B.n437 10.6151
R2541 B.n860 B.n437 10.6151
R2542 B.n861 B.n860 10.6151
R2543 B.n862 B.n861 10.6151
R2544 B.n862 B.n429 10.6151
R2545 B.n872 B.n429 10.6151
R2546 B.n873 B.n872 10.6151
R2547 B.n874 B.n873 10.6151
R2548 B.n874 B.n421 10.6151
R2549 B.n884 B.n421 10.6151
R2550 B.n885 B.n884 10.6151
R2551 B.n886 B.n885 10.6151
R2552 B.n886 B.n413 10.6151
R2553 B.n896 B.n413 10.6151
R2554 B.n897 B.n896 10.6151
R2555 B.n898 B.n897 10.6151
R2556 B.n898 B.n405 10.6151
R2557 B.n908 B.n405 10.6151
R2558 B.n909 B.n908 10.6151
R2559 B.n910 B.n909 10.6151
R2560 B.n910 B.n396 10.6151
R2561 B.n920 B.n396 10.6151
R2562 B.n921 B.n920 10.6151
R2563 B.n922 B.n921 10.6151
R2564 B.n922 B.n389 10.6151
R2565 B.n932 B.n389 10.6151
R2566 B.n933 B.n932 10.6151
R2567 B.n934 B.n933 10.6151
R2568 B.n934 B.n381 10.6151
R2569 B.n944 B.n381 10.6151
R2570 B.n945 B.n944 10.6151
R2571 B.n946 B.n945 10.6151
R2572 B.n946 B.n373 10.6151
R2573 B.n956 B.n373 10.6151
R2574 B.n957 B.n956 10.6151
R2575 B.n958 B.n957 10.6151
R2576 B.n958 B.n365 10.6151
R2577 B.n968 B.n365 10.6151
R2578 B.n969 B.n968 10.6151
R2579 B.n971 B.n969 10.6151
R2580 B.n971 B.n970 10.6151
R2581 B.n970 B.n357 10.6151
R2582 B.n982 B.n357 10.6151
R2583 B.n983 B.n982 10.6151
R2584 B.n984 B.n983 10.6151
R2585 B.n985 B.n984 10.6151
R2586 B.n987 B.n985 10.6151
R2587 B.n988 B.n987 10.6151
R2588 B.n989 B.n988 10.6151
R2589 B.n990 B.n989 10.6151
R2590 B.n992 B.n990 10.6151
R2591 B.n993 B.n992 10.6151
R2592 B.n994 B.n993 10.6151
R2593 B.n995 B.n994 10.6151
R2594 B.n997 B.n995 10.6151
R2595 B.n998 B.n997 10.6151
R2596 B.n999 B.n998 10.6151
R2597 B.n1000 B.n999 10.6151
R2598 B.n1002 B.n1000 10.6151
R2599 B.n1003 B.n1002 10.6151
R2600 B.n1004 B.n1003 10.6151
R2601 B.n1005 B.n1004 10.6151
R2602 B.n1007 B.n1005 10.6151
R2603 B.n1008 B.n1007 10.6151
R2604 B.n1009 B.n1008 10.6151
R2605 B.n1010 B.n1009 10.6151
R2606 B.n1012 B.n1010 10.6151
R2607 B.n1013 B.n1012 10.6151
R2608 B.n1014 B.n1013 10.6151
R2609 B.n1015 B.n1014 10.6151
R2610 B.n1017 B.n1015 10.6151
R2611 B.n1018 B.n1017 10.6151
R2612 B.n1019 B.n1018 10.6151
R2613 B.n1020 B.n1019 10.6151
R2614 B.n1022 B.n1020 10.6151
R2615 B.n1023 B.n1022 10.6151
R2616 B.n1024 B.n1023 10.6151
R2617 B.n1025 B.n1024 10.6151
R2618 B.n1027 B.n1025 10.6151
R2619 B.n1028 B.n1027 10.6151
R2620 B.n1029 B.n1028 10.6151
R2621 B.n1030 B.n1029 10.6151
R2622 B.n1032 B.n1030 10.6151
R2623 B.n1033 B.n1032 10.6151
R2624 B.n1034 B.n1033 10.6151
R2625 B.n1035 B.n1034 10.6151
R2626 B.n1037 B.n1035 10.6151
R2627 B.n1038 B.n1037 10.6151
R2628 B.n1039 B.n1038 10.6151
R2629 B.n1040 B.n1039 10.6151
R2630 B.n1042 B.n1040 10.6151
R2631 B.n1043 B.n1042 10.6151
R2632 B.n1044 B.n1043 10.6151
R2633 B.n1045 B.n1044 10.6151
R2634 B.n1047 B.n1045 10.6151
R2635 B.n1048 B.n1047 10.6151
R2636 B.n1049 B.n1048 10.6151
R2637 B.n1050 B.n1049 10.6151
R2638 B.n1052 B.n1050 10.6151
R2639 B.n1053 B.n1052 10.6151
R2640 B.n1054 B.n1053 10.6151
R2641 B.n1055 B.n1054 10.6151
R2642 B.n1057 B.n1055 10.6151
R2643 B.n1058 B.n1057 10.6151
R2644 B.n1059 B.n1058 10.6151
R2645 B.n1060 B.n1059 10.6151
R2646 B.n1062 B.n1060 10.6151
R2647 B.n1063 B.n1062 10.6151
R2648 B.n1064 B.n1063 10.6151
R2649 B.n1065 B.n1064 10.6151
R2650 B.n1067 B.n1065 10.6151
R2651 B.n1068 B.n1067 10.6151
R2652 B.n1069 B.n1068 10.6151
R2653 B.n1070 B.n1069 10.6151
R2654 B.n1072 B.n1070 10.6151
R2655 B.n1073 B.n1072 10.6151
R2656 B.n1074 B.n1073 10.6151
R2657 B.n1075 B.n1074 10.6151
R2658 B.n1077 B.n1075 10.6151
R2659 B.n1078 B.n1077 10.6151
R2660 B.n1079 B.n1078 10.6151
R2661 B.n1080 B.n1079 10.6151
R2662 B.n1082 B.n1080 10.6151
R2663 B.n1083 B.n1082 10.6151
R2664 B.n1084 B.n1083 10.6151
R2665 B.n1085 B.n1084 10.6151
R2666 B.n1087 B.n1085 10.6151
R2667 B.n1088 B.n1087 10.6151
R2668 B.n566 B.n519 10.6151
R2669 B.n566 B.n565 10.6151
R2670 B.n572 B.n565 10.6151
R2671 B.n573 B.n572 10.6151
R2672 B.n574 B.n573 10.6151
R2673 B.n574 B.n563 10.6151
R2674 B.n580 B.n563 10.6151
R2675 B.n581 B.n580 10.6151
R2676 B.n582 B.n581 10.6151
R2677 B.n582 B.n561 10.6151
R2678 B.n588 B.n561 10.6151
R2679 B.n589 B.n588 10.6151
R2680 B.n590 B.n589 10.6151
R2681 B.n590 B.n559 10.6151
R2682 B.n596 B.n559 10.6151
R2683 B.n597 B.n596 10.6151
R2684 B.n598 B.n597 10.6151
R2685 B.n598 B.n557 10.6151
R2686 B.n604 B.n557 10.6151
R2687 B.n605 B.n604 10.6151
R2688 B.n606 B.n605 10.6151
R2689 B.n606 B.n555 10.6151
R2690 B.n612 B.n555 10.6151
R2691 B.n613 B.n612 10.6151
R2692 B.n614 B.n613 10.6151
R2693 B.n614 B.n553 10.6151
R2694 B.n620 B.n553 10.6151
R2695 B.n621 B.n620 10.6151
R2696 B.n622 B.n621 10.6151
R2697 B.n622 B.n551 10.6151
R2698 B.n628 B.n551 10.6151
R2699 B.n629 B.n628 10.6151
R2700 B.n630 B.n629 10.6151
R2701 B.n630 B.n549 10.6151
R2702 B.n636 B.n549 10.6151
R2703 B.n639 B.n638 10.6151
R2704 B.n639 B.n545 10.6151
R2705 B.n645 B.n545 10.6151
R2706 B.n646 B.n645 10.6151
R2707 B.n647 B.n646 10.6151
R2708 B.n647 B.n543 10.6151
R2709 B.n653 B.n543 10.6151
R2710 B.n654 B.n653 10.6151
R2711 B.n656 B.n539 10.6151
R2712 B.n662 B.n539 10.6151
R2713 B.n663 B.n662 10.6151
R2714 B.n664 B.n663 10.6151
R2715 B.n664 B.n537 10.6151
R2716 B.n670 B.n537 10.6151
R2717 B.n671 B.n670 10.6151
R2718 B.n672 B.n671 10.6151
R2719 B.n672 B.n535 10.6151
R2720 B.n678 B.n535 10.6151
R2721 B.n679 B.n678 10.6151
R2722 B.n680 B.n679 10.6151
R2723 B.n680 B.n533 10.6151
R2724 B.n686 B.n533 10.6151
R2725 B.n687 B.n686 10.6151
R2726 B.n688 B.n687 10.6151
R2727 B.n688 B.n531 10.6151
R2728 B.n694 B.n531 10.6151
R2729 B.n695 B.n694 10.6151
R2730 B.n696 B.n695 10.6151
R2731 B.n696 B.n529 10.6151
R2732 B.n702 B.n529 10.6151
R2733 B.n703 B.n702 10.6151
R2734 B.n704 B.n703 10.6151
R2735 B.n704 B.n527 10.6151
R2736 B.n710 B.n527 10.6151
R2737 B.n711 B.n710 10.6151
R2738 B.n712 B.n711 10.6151
R2739 B.n712 B.n525 10.6151
R2740 B.n718 B.n525 10.6151
R2741 B.n719 B.n718 10.6151
R2742 B.n720 B.n719 10.6151
R2743 B.n720 B.n523 10.6151
R2744 B.n726 B.n523 10.6151
R2745 B.n727 B.n726 10.6151
R2746 B.n733 B.n732 10.6151
R2747 B.n734 B.n733 10.6151
R2748 B.n734 B.n511 10.6151
R2749 B.n744 B.n511 10.6151
R2750 B.n745 B.n744 10.6151
R2751 B.n746 B.n745 10.6151
R2752 B.n746 B.n503 10.6151
R2753 B.n757 B.n503 10.6151
R2754 B.n758 B.n757 10.6151
R2755 B.n759 B.n758 10.6151
R2756 B.n759 B.n496 10.6151
R2757 B.n769 B.n496 10.6151
R2758 B.n770 B.n769 10.6151
R2759 B.n771 B.n770 10.6151
R2760 B.n771 B.n488 10.6151
R2761 B.n781 B.n488 10.6151
R2762 B.n782 B.n781 10.6151
R2763 B.n783 B.n782 10.6151
R2764 B.n783 B.n480 10.6151
R2765 B.n793 B.n480 10.6151
R2766 B.n794 B.n793 10.6151
R2767 B.n795 B.n794 10.6151
R2768 B.n795 B.n472 10.6151
R2769 B.n806 B.n472 10.6151
R2770 B.n807 B.n806 10.6151
R2771 B.n808 B.n807 10.6151
R2772 B.n808 B.n465 10.6151
R2773 B.n818 B.n465 10.6151
R2774 B.n819 B.n818 10.6151
R2775 B.n820 B.n819 10.6151
R2776 B.n820 B.n457 10.6151
R2777 B.n830 B.n457 10.6151
R2778 B.n831 B.n830 10.6151
R2779 B.n832 B.n831 10.6151
R2780 B.n832 B.n449 10.6151
R2781 B.n842 B.n449 10.6151
R2782 B.n843 B.n842 10.6151
R2783 B.n844 B.n843 10.6151
R2784 B.n844 B.n441 10.6151
R2785 B.n854 B.n441 10.6151
R2786 B.n855 B.n854 10.6151
R2787 B.n856 B.n855 10.6151
R2788 B.n856 B.n433 10.6151
R2789 B.n866 B.n433 10.6151
R2790 B.n867 B.n866 10.6151
R2791 B.n868 B.n867 10.6151
R2792 B.n868 B.n425 10.6151
R2793 B.n878 B.n425 10.6151
R2794 B.n879 B.n878 10.6151
R2795 B.n880 B.n879 10.6151
R2796 B.n880 B.n417 10.6151
R2797 B.n890 B.n417 10.6151
R2798 B.n891 B.n890 10.6151
R2799 B.n892 B.n891 10.6151
R2800 B.n892 B.n409 10.6151
R2801 B.n902 B.n409 10.6151
R2802 B.n903 B.n902 10.6151
R2803 B.n904 B.n903 10.6151
R2804 B.n904 B.n401 10.6151
R2805 B.n914 B.n401 10.6151
R2806 B.n915 B.n914 10.6151
R2807 B.n916 B.n915 10.6151
R2808 B.n916 B.n393 10.6151
R2809 B.n926 B.n393 10.6151
R2810 B.n927 B.n926 10.6151
R2811 B.n928 B.n927 10.6151
R2812 B.n928 B.n385 10.6151
R2813 B.n938 B.n385 10.6151
R2814 B.n939 B.n938 10.6151
R2815 B.n940 B.n939 10.6151
R2816 B.n940 B.n377 10.6151
R2817 B.n950 B.n377 10.6151
R2818 B.n951 B.n950 10.6151
R2819 B.n952 B.n951 10.6151
R2820 B.n952 B.n369 10.6151
R2821 B.n962 B.n369 10.6151
R2822 B.n963 B.n962 10.6151
R2823 B.n964 B.n963 10.6151
R2824 B.n964 B.n361 10.6151
R2825 B.n975 B.n361 10.6151
R2826 B.n976 B.n975 10.6151
R2827 B.n977 B.n976 10.6151
R2828 B.n977 B.n0 10.6151
R2829 B.n1256 B.n1 10.6151
R2830 B.n1256 B.n1255 10.6151
R2831 B.n1255 B.n1254 10.6151
R2832 B.n1254 B.n10 10.6151
R2833 B.n1248 B.n10 10.6151
R2834 B.n1248 B.n1247 10.6151
R2835 B.n1247 B.n1246 10.6151
R2836 B.n1246 B.n17 10.6151
R2837 B.n1240 B.n17 10.6151
R2838 B.n1240 B.n1239 10.6151
R2839 B.n1239 B.n1238 10.6151
R2840 B.n1238 B.n24 10.6151
R2841 B.n1232 B.n24 10.6151
R2842 B.n1232 B.n1231 10.6151
R2843 B.n1231 B.n1230 10.6151
R2844 B.n1230 B.n31 10.6151
R2845 B.n1224 B.n31 10.6151
R2846 B.n1224 B.n1223 10.6151
R2847 B.n1223 B.n1222 10.6151
R2848 B.n1222 B.n38 10.6151
R2849 B.n1216 B.n38 10.6151
R2850 B.n1216 B.n1215 10.6151
R2851 B.n1215 B.n1214 10.6151
R2852 B.n1214 B.n45 10.6151
R2853 B.n1208 B.n45 10.6151
R2854 B.n1208 B.n1207 10.6151
R2855 B.n1207 B.n1206 10.6151
R2856 B.n1206 B.n52 10.6151
R2857 B.n1200 B.n52 10.6151
R2858 B.n1200 B.n1199 10.6151
R2859 B.n1199 B.n1198 10.6151
R2860 B.n1198 B.n59 10.6151
R2861 B.n1192 B.n59 10.6151
R2862 B.n1192 B.n1191 10.6151
R2863 B.n1191 B.n1190 10.6151
R2864 B.n1190 B.n66 10.6151
R2865 B.n1184 B.n66 10.6151
R2866 B.n1184 B.n1183 10.6151
R2867 B.n1183 B.n1182 10.6151
R2868 B.n1182 B.n73 10.6151
R2869 B.n1176 B.n73 10.6151
R2870 B.n1176 B.n1175 10.6151
R2871 B.n1175 B.n1174 10.6151
R2872 B.n1174 B.n80 10.6151
R2873 B.n1168 B.n80 10.6151
R2874 B.n1168 B.n1167 10.6151
R2875 B.n1167 B.n1166 10.6151
R2876 B.n1166 B.n87 10.6151
R2877 B.n1160 B.n87 10.6151
R2878 B.n1160 B.n1159 10.6151
R2879 B.n1159 B.n1158 10.6151
R2880 B.n1158 B.n94 10.6151
R2881 B.n1152 B.n94 10.6151
R2882 B.n1152 B.n1151 10.6151
R2883 B.n1151 B.n1150 10.6151
R2884 B.n1150 B.n101 10.6151
R2885 B.n1144 B.n101 10.6151
R2886 B.n1144 B.n1143 10.6151
R2887 B.n1143 B.n1142 10.6151
R2888 B.n1142 B.n107 10.6151
R2889 B.n1136 B.n107 10.6151
R2890 B.n1136 B.n1135 10.6151
R2891 B.n1135 B.n1134 10.6151
R2892 B.n1134 B.n115 10.6151
R2893 B.n1128 B.n115 10.6151
R2894 B.n1128 B.n1127 10.6151
R2895 B.n1127 B.n1126 10.6151
R2896 B.n1126 B.n122 10.6151
R2897 B.n1120 B.n122 10.6151
R2898 B.n1120 B.n1119 10.6151
R2899 B.n1119 B.n1118 10.6151
R2900 B.n1118 B.n129 10.6151
R2901 B.n1112 B.n129 10.6151
R2902 B.n1112 B.n1111 10.6151
R2903 B.n1111 B.n1110 10.6151
R2904 B.n1110 B.n135 10.6151
R2905 B.n1104 B.n135 10.6151
R2906 B.n1104 B.n1103 10.6151
R2907 B.n1103 B.n1102 10.6151
R2908 B.n1102 B.n143 10.6151
R2909 B.n1096 B.n143 10.6151
R2910 B.n1096 B.n1095 10.6151
R2911 B.n1095 B.n1094 10.6151
R2912 B.n270 B.n198 6.5566
R2913 B.n287 B.n286 6.5566
R2914 B.n638 B.n637 6.5566
R2915 B.n655 B.n654 6.5566
R2916 B.n267 B.n198 4.05904
R2917 B.n288 B.n287 4.05904
R2918 B.n637 B.n636 4.05904
R2919 B.n656 B.n655 4.05904
R2920 B.n960 B.t7 2.87538
R2921 B.n1244 B.t9 2.87538
R2922 B.n1262 B.n0 2.81026
R2923 B.n1262 B.n1 2.81026
R2924 B.n846 B.t5 1.43794
R2925 B.t0 B.n1170 1.43794
R2926 VP.n34 VP.n33 161.3
R2927 VP.n35 VP.n30 161.3
R2928 VP.n37 VP.n36 161.3
R2929 VP.n38 VP.n29 161.3
R2930 VP.n40 VP.n39 161.3
R2931 VP.n41 VP.n28 161.3
R2932 VP.n43 VP.n42 161.3
R2933 VP.n44 VP.n27 161.3
R2934 VP.n46 VP.n45 161.3
R2935 VP.n48 VP.n26 161.3
R2936 VP.n50 VP.n49 161.3
R2937 VP.n51 VP.n25 161.3
R2938 VP.n53 VP.n52 161.3
R2939 VP.n54 VP.n24 161.3
R2940 VP.n56 VP.n55 161.3
R2941 VP.n57 VP.n23 161.3
R2942 VP.n59 VP.n58 161.3
R2943 VP.n60 VP.n22 161.3
R2944 VP.n63 VP.n62 161.3
R2945 VP.n64 VP.n21 161.3
R2946 VP.n66 VP.n65 161.3
R2947 VP.n67 VP.n20 161.3
R2948 VP.n69 VP.n68 161.3
R2949 VP.n70 VP.n19 161.3
R2950 VP.n72 VP.n71 161.3
R2951 VP.n73 VP.n18 161.3
R2952 VP.n130 VP.n0 161.3
R2953 VP.n129 VP.n128 161.3
R2954 VP.n127 VP.n1 161.3
R2955 VP.n126 VP.n125 161.3
R2956 VP.n124 VP.n2 161.3
R2957 VP.n123 VP.n122 161.3
R2958 VP.n121 VP.n3 161.3
R2959 VP.n120 VP.n119 161.3
R2960 VP.n117 VP.n4 161.3
R2961 VP.n116 VP.n115 161.3
R2962 VP.n114 VP.n5 161.3
R2963 VP.n113 VP.n112 161.3
R2964 VP.n111 VP.n6 161.3
R2965 VP.n110 VP.n109 161.3
R2966 VP.n108 VP.n7 161.3
R2967 VP.n107 VP.n106 161.3
R2968 VP.n105 VP.n8 161.3
R2969 VP.n103 VP.n102 161.3
R2970 VP.n101 VP.n9 161.3
R2971 VP.n100 VP.n99 161.3
R2972 VP.n98 VP.n10 161.3
R2973 VP.n97 VP.n96 161.3
R2974 VP.n95 VP.n11 161.3
R2975 VP.n94 VP.n93 161.3
R2976 VP.n92 VP.n12 161.3
R2977 VP.n91 VP.n90 161.3
R2978 VP.n89 VP.n88 161.3
R2979 VP.n87 VP.n14 161.3
R2980 VP.n86 VP.n85 161.3
R2981 VP.n84 VP.n15 161.3
R2982 VP.n83 VP.n82 161.3
R2983 VP.n81 VP.n16 161.3
R2984 VP.n80 VP.n79 161.3
R2985 VP.n78 VP.n17 161.3
R2986 VP.n32 VP.t4 93.0541
R2987 VP.n32 VP.n31 72.0574
R2988 VP.n77 VP.n76 64.0762
R2989 VP.n132 VP.n131 64.0762
R2990 VP.n75 VP.n74 64.0762
R2991 VP.n76 VP.t0 60.7349
R2992 VP.n13 VP.t3 60.7349
R2993 VP.n104 VP.t7 60.7349
R2994 VP.n118 VP.t5 60.7349
R2995 VP.n131 VP.t2 60.7349
R2996 VP.n74 VP.t9 60.7349
R2997 VP.n61 VP.t6 60.7349
R2998 VP.n47 VP.t1 60.7349
R2999 VP.n31 VP.t8 60.7349
R3000 VP.n77 VP.n75 59.3335
R3001 VP.n82 VP.n15 56.5193
R3002 VP.n125 VP.n124 56.5193
R3003 VP.n68 VP.n67 56.5193
R3004 VP.n98 VP.n97 49.7204
R3005 VP.n111 VP.n110 49.7204
R3006 VP.n54 VP.n53 49.7204
R3007 VP.n41 VP.n40 49.7204
R3008 VP.n97 VP.n11 31.2664
R3009 VP.n112 VP.n111 31.2664
R3010 VP.n55 VP.n54 31.2664
R3011 VP.n40 VP.n29 31.2664
R3012 VP.n80 VP.n17 24.4675
R3013 VP.n81 VP.n80 24.4675
R3014 VP.n82 VP.n81 24.4675
R3015 VP.n86 VP.n15 24.4675
R3016 VP.n87 VP.n86 24.4675
R3017 VP.n88 VP.n87 24.4675
R3018 VP.n92 VP.n91 24.4675
R3019 VP.n93 VP.n92 24.4675
R3020 VP.n93 VP.n11 24.4675
R3021 VP.n99 VP.n98 24.4675
R3022 VP.n99 VP.n9 24.4675
R3023 VP.n103 VP.n9 24.4675
R3024 VP.n106 VP.n105 24.4675
R3025 VP.n106 VP.n7 24.4675
R3026 VP.n110 VP.n7 24.4675
R3027 VP.n112 VP.n5 24.4675
R3028 VP.n116 VP.n5 24.4675
R3029 VP.n117 VP.n116 24.4675
R3030 VP.n119 VP.n3 24.4675
R3031 VP.n123 VP.n3 24.4675
R3032 VP.n124 VP.n123 24.4675
R3033 VP.n125 VP.n1 24.4675
R3034 VP.n129 VP.n1 24.4675
R3035 VP.n130 VP.n129 24.4675
R3036 VP.n68 VP.n19 24.4675
R3037 VP.n72 VP.n19 24.4675
R3038 VP.n73 VP.n72 24.4675
R3039 VP.n55 VP.n23 24.4675
R3040 VP.n59 VP.n23 24.4675
R3041 VP.n60 VP.n59 24.4675
R3042 VP.n62 VP.n21 24.4675
R3043 VP.n66 VP.n21 24.4675
R3044 VP.n67 VP.n66 24.4675
R3045 VP.n42 VP.n41 24.4675
R3046 VP.n42 VP.n27 24.4675
R3047 VP.n46 VP.n27 24.4675
R3048 VP.n49 VP.n48 24.4675
R3049 VP.n49 VP.n25 24.4675
R3050 VP.n53 VP.n25 24.4675
R3051 VP.n35 VP.n34 24.4675
R3052 VP.n36 VP.n35 24.4675
R3053 VP.n36 VP.n29 24.4675
R3054 VP.n88 VP.n13 21.5315
R3055 VP.n119 VP.n118 21.5315
R3056 VP.n62 VP.n61 21.5315
R3057 VP.n76 VP.n17 18.1061
R3058 VP.n131 VP.n130 18.1061
R3059 VP.n74 VP.n73 18.1061
R3060 VP.n104 VP.n103 12.234
R3061 VP.n105 VP.n104 12.234
R3062 VP.n47 VP.n46 12.234
R3063 VP.n48 VP.n47 12.234
R3064 VP.n91 VP.n13 2.93654
R3065 VP.n118 VP.n117 2.93654
R3066 VP.n61 VP.n60 2.93654
R3067 VP.n34 VP.n31 2.93654
R3068 VP.n33 VP.n32 2.75932
R3069 VP.n75 VP.n18 0.417535
R3070 VP.n78 VP.n77 0.417535
R3071 VP.n132 VP.n0 0.417535
R3072 VP VP.n132 0.394291
R3073 VP.n33 VP.n30 0.189894
R3074 VP.n37 VP.n30 0.189894
R3075 VP.n38 VP.n37 0.189894
R3076 VP.n39 VP.n38 0.189894
R3077 VP.n39 VP.n28 0.189894
R3078 VP.n43 VP.n28 0.189894
R3079 VP.n44 VP.n43 0.189894
R3080 VP.n45 VP.n44 0.189894
R3081 VP.n45 VP.n26 0.189894
R3082 VP.n50 VP.n26 0.189894
R3083 VP.n51 VP.n50 0.189894
R3084 VP.n52 VP.n51 0.189894
R3085 VP.n52 VP.n24 0.189894
R3086 VP.n56 VP.n24 0.189894
R3087 VP.n57 VP.n56 0.189894
R3088 VP.n58 VP.n57 0.189894
R3089 VP.n58 VP.n22 0.189894
R3090 VP.n63 VP.n22 0.189894
R3091 VP.n64 VP.n63 0.189894
R3092 VP.n65 VP.n64 0.189894
R3093 VP.n65 VP.n20 0.189894
R3094 VP.n69 VP.n20 0.189894
R3095 VP.n70 VP.n69 0.189894
R3096 VP.n71 VP.n70 0.189894
R3097 VP.n71 VP.n18 0.189894
R3098 VP.n79 VP.n78 0.189894
R3099 VP.n79 VP.n16 0.189894
R3100 VP.n83 VP.n16 0.189894
R3101 VP.n84 VP.n83 0.189894
R3102 VP.n85 VP.n84 0.189894
R3103 VP.n85 VP.n14 0.189894
R3104 VP.n89 VP.n14 0.189894
R3105 VP.n90 VP.n89 0.189894
R3106 VP.n90 VP.n12 0.189894
R3107 VP.n94 VP.n12 0.189894
R3108 VP.n95 VP.n94 0.189894
R3109 VP.n96 VP.n95 0.189894
R3110 VP.n96 VP.n10 0.189894
R3111 VP.n100 VP.n10 0.189894
R3112 VP.n101 VP.n100 0.189894
R3113 VP.n102 VP.n101 0.189894
R3114 VP.n102 VP.n8 0.189894
R3115 VP.n107 VP.n8 0.189894
R3116 VP.n108 VP.n107 0.189894
R3117 VP.n109 VP.n108 0.189894
R3118 VP.n109 VP.n6 0.189894
R3119 VP.n113 VP.n6 0.189894
R3120 VP.n114 VP.n113 0.189894
R3121 VP.n115 VP.n114 0.189894
R3122 VP.n115 VP.n4 0.189894
R3123 VP.n120 VP.n4 0.189894
R3124 VP.n121 VP.n120 0.189894
R3125 VP.n122 VP.n121 0.189894
R3126 VP.n122 VP.n2 0.189894
R3127 VP.n126 VP.n2 0.189894
R3128 VP.n127 VP.n126 0.189894
R3129 VP.n128 VP.n127 0.189894
R3130 VP.n128 VP.n0 0.189894
R3131 VDD1.n48 VDD1.n0 289.615
R3132 VDD1.n103 VDD1.n55 289.615
R3133 VDD1.n49 VDD1.n48 185
R3134 VDD1.n47 VDD1.n46 185
R3135 VDD1.n4 VDD1.n3 185
R3136 VDD1.n41 VDD1.n40 185
R3137 VDD1.n39 VDD1.n6 185
R3138 VDD1.n38 VDD1.n37 185
R3139 VDD1.n9 VDD1.n7 185
R3140 VDD1.n32 VDD1.n31 185
R3141 VDD1.n30 VDD1.n29 185
R3142 VDD1.n13 VDD1.n12 185
R3143 VDD1.n24 VDD1.n23 185
R3144 VDD1.n22 VDD1.n21 185
R3145 VDD1.n17 VDD1.n16 185
R3146 VDD1.n71 VDD1.n70 185
R3147 VDD1.n76 VDD1.n75 185
R3148 VDD1.n78 VDD1.n77 185
R3149 VDD1.n67 VDD1.n66 185
R3150 VDD1.n84 VDD1.n83 185
R3151 VDD1.n86 VDD1.n85 185
R3152 VDD1.n63 VDD1.n62 185
R3153 VDD1.n93 VDD1.n92 185
R3154 VDD1.n94 VDD1.n61 185
R3155 VDD1.n96 VDD1.n95 185
R3156 VDD1.n59 VDD1.n58 185
R3157 VDD1.n102 VDD1.n101 185
R3158 VDD1.n104 VDD1.n103 185
R3159 VDD1.n18 VDD1.t5 149.524
R3160 VDD1.n72 VDD1.t9 149.524
R3161 VDD1.n48 VDD1.n47 104.615
R3162 VDD1.n47 VDD1.n3 104.615
R3163 VDD1.n40 VDD1.n3 104.615
R3164 VDD1.n40 VDD1.n39 104.615
R3165 VDD1.n39 VDD1.n38 104.615
R3166 VDD1.n38 VDD1.n7 104.615
R3167 VDD1.n31 VDD1.n7 104.615
R3168 VDD1.n31 VDD1.n30 104.615
R3169 VDD1.n30 VDD1.n12 104.615
R3170 VDD1.n23 VDD1.n12 104.615
R3171 VDD1.n23 VDD1.n22 104.615
R3172 VDD1.n22 VDD1.n16 104.615
R3173 VDD1.n76 VDD1.n70 104.615
R3174 VDD1.n77 VDD1.n76 104.615
R3175 VDD1.n77 VDD1.n66 104.615
R3176 VDD1.n84 VDD1.n66 104.615
R3177 VDD1.n85 VDD1.n84 104.615
R3178 VDD1.n85 VDD1.n62 104.615
R3179 VDD1.n93 VDD1.n62 104.615
R3180 VDD1.n94 VDD1.n93 104.615
R3181 VDD1.n95 VDD1.n94 104.615
R3182 VDD1.n95 VDD1.n58 104.615
R3183 VDD1.n102 VDD1.n58 104.615
R3184 VDD1.n103 VDD1.n102 104.615
R3185 VDD1.n111 VDD1.n110 66.729
R3186 VDD1.n54 VDD1.n53 63.9979
R3187 VDD1.n113 VDD1.n112 63.9977
R3188 VDD1.n109 VDD1.n108 63.9977
R3189 VDD1.n54 VDD1.n52 53.9372
R3190 VDD1.n109 VDD1.n107 53.9372
R3191 VDD1.n113 VDD1.n111 52.4513
R3192 VDD1.t5 VDD1.n16 52.3082
R3193 VDD1.t9 VDD1.n70 52.3082
R3194 VDD1.n41 VDD1.n6 13.1884
R3195 VDD1.n96 VDD1.n61 13.1884
R3196 VDD1.n42 VDD1.n4 12.8005
R3197 VDD1.n37 VDD1.n8 12.8005
R3198 VDD1.n92 VDD1.n91 12.8005
R3199 VDD1.n97 VDD1.n59 12.8005
R3200 VDD1.n46 VDD1.n45 12.0247
R3201 VDD1.n36 VDD1.n9 12.0247
R3202 VDD1.n90 VDD1.n63 12.0247
R3203 VDD1.n101 VDD1.n100 12.0247
R3204 VDD1.n49 VDD1.n2 11.249
R3205 VDD1.n33 VDD1.n32 11.249
R3206 VDD1.n87 VDD1.n86 11.249
R3207 VDD1.n104 VDD1.n57 11.249
R3208 VDD1.n50 VDD1.n0 10.4732
R3209 VDD1.n29 VDD1.n11 10.4732
R3210 VDD1.n83 VDD1.n65 10.4732
R3211 VDD1.n105 VDD1.n55 10.4732
R3212 VDD1.n18 VDD1.n17 10.2747
R3213 VDD1.n72 VDD1.n71 10.2747
R3214 VDD1.n28 VDD1.n13 9.69747
R3215 VDD1.n82 VDD1.n67 9.69747
R3216 VDD1.n52 VDD1.n51 9.45567
R3217 VDD1.n107 VDD1.n106 9.45567
R3218 VDD1.n20 VDD1.n19 9.3005
R3219 VDD1.n15 VDD1.n14 9.3005
R3220 VDD1.n26 VDD1.n25 9.3005
R3221 VDD1.n28 VDD1.n27 9.3005
R3222 VDD1.n11 VDD1.n10 9.3005
R3223 VDD1.n34 VDD1.n33 9.3005
R3224 VDD1.n36 VDD1.n35 9.3005
R3225 VDD1.n8 VDD1.n5 9.3005
R3226 VDD1.n51 VDD1.n50 9.3005
R3227 VDD1.n2 VDD1.n1 9.3005
R3228 VDD1.n45 VDD1.n44 9.3005
R3229 VDD1.n43 VDD1.n42 9.3005
R3230 VDD1.n106 VDD1.n105 9.3005
R3231 VDD1.n57 VDD1.n56 9.3005
R3232 VDD1.n100 VDD1.n99 9.3005
R3233 VDD1.n98 VDD1.n97 9.3005
R3234 VDD1.n74 VDD1.n73 9.3005
R3235 VDD1.n69 VDD1.n68 9.3005
R3236 VDD1.n80 VDD1.n79 9.3005
R3237 VDD1.n82 VDD1.n81 9.3005
R3238 VDD1.n65 VDD1.n64 9.3005
R3239 VDD1.n88 VDD1.n87 9.3005
R3240 VDD1.n90 VDD1.n89 9.3005
R3241 VDD1.n91 VDD1.n60 9.3005
R3242 VDD1.n25 VDD1.n24 8.92171
R3243 VDD1.n79 VDD1.n78 8.92171
R3244 VDD1.n21 VDD1.n15 8.14595
R3245 VDD1.n75 VDD1.n69 8.14595
R3246 VDD1.n20 VDD1.n17 7.3702
R3247 VDD1.n74 VDD1.n71 7.3702
R3248 VDD1.n21 VDD1.n20 5.81868
R3249 VDD1.n75 VDD1.n74 5.81868
R3250 VDD1.n24 VDD1.n15 5.04292
R3251 VDD1.n78 VDD1.n69 5.04292
R3252 VDD1.n25 VDD1.n13 4.26717
R3253 VDD1.n79 VDD1.n67 4.26717
R3254 VDD1.n52 VDD1.n0 3.49141
R3255 VDD1.n29 VDD1.n28 3.49141
R3256 VDD1.n83 VDD1.n82 3.49141
R3257 VDD1.n107 VDD1.n55 3.49141
R3258 VDD1.n19 VDD1.n18 2.84303
R3259 VDD1.n73 VDD1.n72 2.84303
R3260 VDD1 VDD1.n113 2.72895
R3261 VDD1.n50 VDD1.n49 2.71565
R3262 VDD1.n32 VDD1.n11 2.71565
R3263 VDD1.n86 VDD1.n65 2.71565
R3264 VDD1.n105 VDD1.n104 2.71565
R3265 VDD1.n112 VDD1.t3 1.97458
R3266 VDD1.n112 VDD1.t0 1.97458
R3267 VDD1.n53 VDD1.t1 1.97458
R3268 VDD1.n53 VDD1.t8 1.97458
R3269 VDD1.n110 VDD1.t4 1.97458
R3270 VDD1.n110 VDD1.t7 1.97458
R3271 VDD1.n108 VDD1.t6 1.97458
R3272 VDD1.n108 VDD1.t2 1.97458
R3273 VDD1.n46 VDD1.n2 1.93989
R3274 VDD1.n33 VDD1.n9 1.93989
R3275 VDD1.n87 VDD1.n63 1.93989
R3276 VDD1.n101 VDD1.n57 1.93989
R3277 VDD1.n45 VDD1.n4 1.16414
R3278 VDD1.n37 VDD1.n36 1.16414
R3279 VDD1.n92 VDD1.n90 1.16414
R3280 VDD1.n100 VDD1.n59 1.16414
R3281 VDD1 VDD1.n54 0.987569
R3282 VDD1.n111 VDD1.n109 0.874033
R3283 VDD1.n42 VDD1.n41 0.388379
R3284 VDD1.n8 VDD1.n6 0.388379
R3285 VDD1.n91 VDD1.n61 0.388379
R3286 VDD1.n97 VDD1.n96 0.388379
R3287 VDD1.n51 VDD1.n1 0.155672
R3288 VDD1.n44 VDD1.n1 0.155672
R3289 VDD1.n44 VDD1.n43 0.155672
R3290 VDD1.n43 VDD1.n5 0.155672
R3291 VDD1.n35 VDD1.n5 0.155672
R3292 VDD1.n35 VDD1.n34 0.155672
R3293 VDD1.n34 VDD1.n10 0.155672
R3294 VDD1.n27 VDD1.n10 0.155672
R3295 VDD1.n27 VDD1.n26 0.155672
R3296 VDD1.n26 VDD1.n14 0.155672
R3297 VDD1.n19 VDD1.n14 0.155672
R3298 VDD1.n73 VDD1.n68 0.155672
R3299 VDD1.n80 VDD1.n68 0.155672
R3300 VDD1.n81 VDD1.n80 0.155672
R3301 VDD1.n81 VDD1.n64 0.155672
R3302 VDD1.n88 VDD1.n64 0.155672
R3303 VDD1.n89 VDD1.n88 0.155672
R3304 VDD1.n89 VDD1.n60 0.155672
R3305 VDD1.n98 VDD1.n60 0.155672
R3306 VDD1.n99 VDD1.n98 0.155672
R3307 VDD1.n99 VDD1.n56 0.155672
R3308 VDD1.n106 VDD1.n56 0.155672
C0 VP VN 10.072599f
C1 VP VDD1 10.255199f
C2 VP VTAIL 11.0002f
C3 VP VDD2 0.759073f
C4 VN VDD1 0.156566f
C5 VN VTAIL 10.985499f
C6 VTAIL VDD1 10.4002f
C7 VN VDD2 9.655959f
C8 VDD1 VDD2 3.07381f
C9 VTAIL VDD2 10.4618f
C10 VDD2 B 8.50315f
C11 VDD1 B 8.461293f
C12 VTAIL B 8.439853f
C13 VN B 24.63158f
C14 VP B 23.218887f
C15 VDD1.n0 B 0.035638f
C16 VDD1.n1 B 0.025978f
C17 VDD1.n2 B 0.013959f
C18 VDD1.n3 B 0.032995f
C19 VDD1.n4 B 0.01478f
C20 VDD1.n5 B 0.025978f
C21 VDD1.n6 B 0.01437f
C22 VDD1.n7 B 0.032995f
C23 VDD1.n8 B 0.013959f
C24 VDD1.n9 B 0.01478f
C25 VDD1.n10 B 0.025978f
C26 VDD1.n11 B 0.013959f
C27 VDD1.n12 B 0.032995f
C28 VDD1.n13 B 0.01478f
C29 VDD1.n14 B 0.025978f
C30 VDD1.n15 B 0.013959f
C31 VDD1.n16 B 0.024746f
C32 VDD1.n17 B 0.023325f
C33 VDD1.t5 B 0.055453f
C34 VDD1.n18 B 0.167653f
C35 VDD1.n19 B 1.08291f
C36 VDD1.n20 B 0.013959f
C37 VDD1.n21 B 0.01478f
C38 VDD1.n22 B 0.032995f
C39 VDD1.n23 B 0.032995f
C40 VDD1.n24 B 0.01478f
C41 VDD1.n25 B 0.013959f
C42 VDD1.n26 B 0.025978f
C43 VDD1.n27 B 0.025978f
C44 VDD1.n28 B 0.013959f
C45 VDD1.n29 B 0.01478f
C46 VDD1.n30 B 0.032995f
C47 VDD1.n31 B 0.032995f
C48 VDD1.n32 B 0.01478f
C49 VDD1.n33 B 0.013959f
C50 VDD1.n34 B 0.025978f
C51 VDD1.n35 B 0.025978f
C52 VDD1.n36 B 0.013959f
C53 VDD1.n37 B 0.01478f
C54 VDD1.n38 B 0.032995f
C55 VDD1.n39 B 0.032995f
C56 VDD1.n40 B 0.032995f
C57 VDD1.n41 B 0.01437f
C58 VDD1.n42 B 0.013959f
C59 VDD1.n43 B 0.025978f
C60 VDD1.n44 B 0.025978f
C61 VDD1.n45 B 0.013959f
C62 VDD1.n46 B 0.01478f
C63 VDD1.n47 B 0.032995f
C64 VDD1.n48 B 0.069879f
C65 VDD1.n49 B 0.01478f
C66 VDD1.n50 B 0.013959f
C67 VDD1.n51 B 0.062531f
C68 VDD1.n52 B 0.081902f
C69 VDD1.t1 B 0.205901f
C70 VDD1.t8 B 0.205901f
C71 VDD1.n53 B 1.81456f
C72 VDD1.n54 B 0.94184f
C73 VDD1.n55 B 0.035638f
C74 VDD1.n56 B 0.025978f
C75 VDD1.n57 B 0.013959f
C76 VDD1.n58 B 0.032995f
C77 VDD1.n59 B 0.01478f
C78 VDD1.n60 B 0.025978f
C79 VDD1.n61 B 0.01437f
C80 VDD1.n62 B 0.032995f
C81 VDD1.n63 B 0.01478f
C82 VDD1.n64 B 0.025978f
C83 VDD1.n65 B 0.013959f
C84 VDD1.n66 B 0.032995f
C85 VDD1.n67 B 0.01478f
C86 VDD1.n68 B 0.025978f
C87 VDD1.n69 B 0.013959f
C88 VDD1.n70 B 0.024746f
C89 VDD1.n71 B 0.023325f
C90 VDD1.t9 B 0.055453f
C91 VDD1.n72 B 0.167653f
C92 VDD1.n73 B 1.08291f
C93 VDD1.n74 B 0.013959f
C94 VDD1.n75 B 0.01478f
C95 VDD1.n76 B 0.032995f
C96 VDD1.n77 B 0.032995f
C97 VDD1.n78 B 0.01478f
C98 VDD1.n79 B 0.013959f
C99 VDD1.n80 B 0.025978f
C100 VDD1.n81 B 0.025978f
C101 VDD1.n82 B 0.013959f
C102 VDD1.n83 B 0.01478f
C103 VDD1.n84 B 0.032995f
C104 VDD1.n85 B 0.032995f
C105 VDD1.n86 B 0.01478f
C106 VDD1.n87 B 0.013959f
C107 VDD1.n88 B 0.025978f
C108 VDD1.n89 B 0.025978f
C109 VDD1.n90 B 0.013959f
C110 VDD1.n91 B 0.013959f
C111 VDD1.n92 B 0.01478f
C112 VDD1.n93 B 0.032995f
C113 VDD1.n94 B 0.032995f
C114 VDD1.n95 B 0.032995f
C115 VDD1.n96 B 0.01437f
C116 VDD1.n97 B 0.013959f
C117 VDD1.n98 B 0.025978f
C118 VDD1.n99 B 0.025978f
C119 VDD1.n100 B 0.013959f
C120 VDD1.n101 B 0.01478f
C121 VDD1.n102 B 0.032995f
C122 VDD1.n103 B 0.069879f
C123 VDD1.n104 B 0.01478f
C124 VDD1.n105 B 0.013959f
C125 VDD1.n106 B 0.062531f
C126 VDD1.n107 B 0.081902f
C127 VDD1.t6 B 0.205901f
C128 VDD1.t2 B 0.205901f
C129 VDD1.n108 B 1.81456f
C130 VDD1.n109 B 0.933033f
C131 VDD1.t4 B 0.205901f
C132 VDD1.t7 B 0.205901f
C133 VDD1.n110 B 1.84571f
C134 VDD1.n111 B 3.80223f
C135 VDD1.t3 B 0.205901f
C136 VDD1.t0 B 0.205901f
C137 VDD1.n112 B 1.81456f
C138 VDD1.n113 B 3.73366f
C139 VP.n0 B 0.032345f
C140 VP.t2 B 1.85979f
C141 VP.n1 B 0.032048f
C142 VP.n2 B 0.017196f
C143 VP.n3 B 0.032048f
C144 VP.n4 B 0.017196f
C145 VP.t5 B 1.85979f
C146 VP.n5 B 0.032048f
C147 VP.n6 B 0.017196f
C148 VP.n7 B 0.032048f
C149 VP.n8 B 0.017196f
C150 VP.t7 B 1.85979f
C151 VP.n9 B 0.032048f
C152 VP.n10 B 0.017196f
C153 VP.n11 B 0.034525f
C154 VP.n12 B 0.017196f
C155 VP.t3 B 1.85979f
C156 VP.n13 B 0.657063f
C157 VP.n14 B 0.017196f
C158 VP.n15 B 0.023427f
C159 VP.n16 B 0.017196f
C160 VP.n17 B 0.027934f
C161 VP.n18 B 0.032345f
C162 VP.t9 B 1.85979f
C163 VP.n19 B 0.032048f
C164 VP.n20 B 0.017196f
C165 VP.n21 B 0.032048f
C166 VP.n22 B 0.017196f
C167 VP.t6 B 1.85979f
C168 VP.n23 B 0.032048f
C169 VP.n24 B 0.017196f
C170 VP.n25 B 0.032048f
C171 VP.n26 B 0.017196f
C172 VP.t1 B 1.85979f
C173 VP.n27 B 0.032048f
C174 VP.n28 B 0.017196f
C175 VP.n29 B 0.034525f
C176 VP.n30 B 0.017196f
C177 VP.t8 B 1.85979f
C178 VP.n31 B 0.71424f
C179 VP.t4 B 2.13467f
C180 VP.n32 B 0.679866f
C181 VP.n33 B 0.230949f
C182 VP.n34 B 0.018125f
C183 VP.n35 B 0.032048f
C184 VP.n36 B 0.032048f
C185 VP.n37 B 0.017196f
C186 VP.n38 B 0.017196f
C187 VP.n39 B 0.017196f
C188 VP.n40 B 0.016004f
C189 VP.n41 B 0.031727f
C190 VP.n42 B 0.032048f
C191 VP.n43 B 0.017196f
C192 VP.n44 B 0.017196f
C193 VP.n45 B 0.017196f
C194 VP.n46 B 0.024137f
C195 VP.n47 B 0.657063f
C196 VP.n48 B 0.024137f
C197 VP.n49 B 0.032048f
C198 VP.n50 B 0.017196f
C199 VP.n51 B 0.017196f
C200 VP.n52 B 0.017196f
C201 VP.n53 B 0.031727f
C202 VP.n54 B 0.016004f
C203 VP.n55 B 0.034525f
C204 VP.n56 B 0.017196f
C205 VP.n57 B 0.017196f
C206 VP.n58 B 0.017196f
C207 VP.n59 B 0.032048f
C208 VP.n60 B 0.018125f
C209 VP.n61 B 0.657063f
C210 VP.n62 B 0.03015f
C211 VP.n63 B 0.017196f
C212 VP.n64 B 0.017196f
C213 VP.n65 B 0.017196f
C214 VP.n66 B 0.032048f
C215 VP.n67 B 0.023427f
C216 VP.n68 B 0.026781f
C217 VP.n69 B 0.017196f
C218 VP.n70 B 0.017196f
C219 VP.n71 B 0.017196f
C220 VP.n72 B 0.032048f
C221 VP.n73 B 0.027934f
C222 VP.n74 B 0.730101f
C223 VP.n75 B 1.26474f
C224 VP.t0 B 1.85979f
C225 VP.n76 B 0.730101f
C226 VP.n77 B 1.27516f
C227 VP.n78 B 0.032345f
C228 VP.n79 B 0.017196f
C229 VP.n80 B 0.032048f
C230 VP.n81 B 0.032048f
C231 VP.n82 B 0.026781f
C232 VP.n83 B 0.017196f
C233 VP.n84 B 0.017196f
C234 VP.n85 B 0.017196f
C235 VP.n86 B 0.032048f
C236 VP.n87 B 0.032048f
C237 VP.n88 B 0.03015f
C238 VP.n89 B 0.017196f
C239 VP.n90 B 0.017196f
C240 VP.n91 B 0.018125f
C241 VP.n92 B 0.032048f
C242 VP.n93 B 0.032048f
C243 VP.n94 B 0.017196f
C244 VP.n95 B 0.017196f
C245 VP.n96 B 0.017196f
C246 VP.n97 B 0.016004f
C247 VP.n98 B 0.031727f
C248 VP.n99 B 0.032048f
C249 VP.n100 B 0.017196f
C250 VP.n101 B 0.017196f
C251 VP.n102 B 0.017196f
C252 VP.n103 B 0.024137f
C253 VP.n104 B 0.657063f
C254 VP.n105 B 0.024137f
C255 VP.n106 B 0.032048f
C256 VP.n107 B 0.017196f
C257 VP.n108 B 0.017196f
C258 VP.n109 B 0.017196f
C259 VP.n110 B 0.031727f
C260 VP.n111 B 0.016004f
C261 VP.n112 B 0.034525f
C262 VP.n113 B 0.017196f
C263 VP.n114 B 0.017196f
C264 VP.n115 B 0.017196f
C265 VP.n116 B 0.032048f
C266 VP.n117 B 0.018125f
C267 VP.n118 B 0.657063f
C268 VP.n119 B 0.03015f
C269 VP.n120 B 0.017196f
C270 VP.n121 B 0.017196f
C271 VP.n122 B 0.017196f
C272 VP.n123 B 0.032048f
C273 VP.n124 B 0.023427f
C274 VP.n125 B 0.026781f
C275 VP.n126 B 0.017196f
C276 VP.n127 B 0.017196f
C277 VP.n128 B 0.017196f
C278 VP.n129 B 0.032048f
C279 VP.n130 B 0.027934f
C280 VP.n131 B 0.730101f
C281 VP.n132 B 0.056788f
C282 VTAIL.t16 B 0.213627f
C283 VTAIL.t12 B 0.213627f
C284 VTAIL.n0 B 1.80739f
C285 VTAIL.n1 B 0.706459f
C286 VTAIL.n2 B 0.036975f
C287 VTAIL.n3 B 0.026953f
C288 VTAIL.n4 B 0.014483f
C289 VTAIL.n5 B 0.034233f
C290 VTAIL.n6 B 0.015335f
C291 VTAIL.n7 B 0.026953f
C292 VTAIL.n8 B 0.014909f
C293 VTAIL.n9 B 0.034233f
C294 VTAIL.n10 B 0.015335f
C295 VTAIL.n11 B 0.026953f
C296 VTAIL.n12 B 0.014483f
C297 VTAIL.n13 B 0.034233f
C298 VTAIL.n14 B 0.015335f
C299 VTAIL.n15 B 0.026953f
C300 VTAIL.n16 B 0.014483f
C301 VTAIL.n17 B 0.025675f
C302 VTAIL.n18 B 0.0242f
C303 VTAIL.t7 B 0.057533f
C304 VTAIL.n19 B 0.173944f
C305 VTAIL.n20 B 1.12354f
C306 VTAIL.n21 B 0.014483f
C307 VTAIL.n22 B 0.015335f
C308 VTAIL.n23 B 0.034233f
C309 VTAIL.n24 B 0.034233f
C310 VTAIL.n25 B 0.015335f
C311 VTAIL.n26 B 0.014483f
C312 VTAIL.n27 B 0.026953f
C313 VTAIL.n28 B 0.026953f
C314 VTAIL.n29 B 0.014483f
C315 VTAIL.n30 B 0.015335f
C316 VTAIL.n31 B 0.034233f
C317 VTAIL.n32 B 0.034233f
C318 VTAIL.n33 B 0.015335f
C319 VTAIL.n34 B 0.014483f
C320 VTAIL.n35 B 0.026953f
C321 VTAIL.n36 B 0.026953f
C322 VTAIL.n37 B 0.014483f
C323 VTAIL.n38 B 0.014483f
C324 VTAIL.n39 B 0.015335f
C325 VTAIL.n40 B 0.034233f
C326 VTAIL.n41 B 0.034233f
C327 VTAIL.n42 B 0.034233f
C328 VTAIL.n43 B 0.014909f
C329 VTAIL.n44 B 0.014483f
C330 VTAIL.n45 B 0.026953f
C331 VTAIL.n46 B 0.026953f
C332 VTAIL.n47 B 0.014483f
C333 VTAIL.n48 B 0.015335f
C334 VTAIL.n49 B 0.034233f
C335 VTAIL.n50 B 0.072501f
C336 VTAIL.n51 B 0.015335f
C337 VTAIL.n52 B 0.014483f
C338 VTAIL.n53 B 0.064877f
C339 VTAIL.n54 B 0.040479f
C340 VTAIL.n55 B 0.549304f
C341 VTAIL.t1 B 0.213627f
C342 VTAIL.t3 B 0.213627f
C343 VTAIL.n56 B 1.80739f
C344 VTAIL.n57 B 0.902614f
C345 VTAIL.t2 B 0.213627f
C346 VTAIL.t5 B 0.213627f
C347 VTAIL.n58 B 1.80739f
C348 VTAIL.n59 B 2.34235f
C349 VTAIL.t13 B 0.213627f
C350 VTAIL.t15 B 0.213627f
C351 VTAIL.n60 B 1.8074f
C352 VTAIL.n61 B 2.34234f
C353 VTAIL.t9 B 0.213627f
C354 VTAIL.t14 B 0.213627f
C355 VTAIL.n62 B 1.8074f
C356 VTAIL.n63 B 0.902603f
C357 VTAIL.n64 B 0.036975f
C358 VTAIL.n65 B 0.026953f
C359 VTAIL.n66 B 0.014483f
C360 VTAIL.n67 B 0.034233f
C361 VTAIL.n68 B 0.015335f
C362 VTAIL.n69 B 0.026953f
C363 VTAIL.n70 B 0.014909f
C364 VTAIL.n71 B 0.034233f
C365 VTAIL.n72 B 0.014483f
C366 VTAIL.n73 B 0.015335f
C367 VTAIL.n74 B 0.026953f
C368 VTAIL.n75 B 0.014483f
C369 VTAIL.n76 B 0.034233f
C370 VTAIL.n77 B 0.015335f
C371 VTAIL.n78 B 0.026953f
C372 VTAIL.n79 B 0.014483f
C373 VTAIL.n80 B 0.025675f
C374 VTAIL.n81 B 0.0242f
C375 VTAIL.t10 B 0.057533f
C376 VTAIL.n82 B 0.173944f
C377 VTAIL.n83 B 1.12354f
C378 VTAIL.n84 B 0.014483f
C379 VTAIL.n85 B 0.015335f
C380 VTAIL.n86 B 0.034233f
C381 VTAIL.n87 B 0.034233f
C382 VTAIL.n88 B 0.015335f
C383 VTAIL.n89 B 0.014483f
C384 VTAIL.n90 B 0.026953f
C385 VTAIL.n91 B 0.026953f
C386 VTAIL.n92 B 0.014483f
C387 VTAIL.n93 B 0.015335f
C388 VTAIL.n94 B 0.034233f
C389 VTAIL.n95 B 0.034233f
C390 VTAIL.n96 B 0.015335f
C391 VTAIL.n97 B 0.014483f
C392 VTAIL.n98 B 0.026953f
C393 VTAIL.n99 B 0.026953f
C394 VTAIL.n100 B 0.014483f
C395 VTAIL.n101 B 0.015335f
C396 VTAIL.n102 B 0.034233f
C397 VTAIL.n103 B 0.034233f
C398 VTAIL.n104 B 0.034233f
C399 VTAIL.n105 B 0.014909f
C400 VTAIL.n106 B 0.014483f
C401 VTAIL.n107 B 0.026953f
C402 VTAIL.n108 B 0.026953f
C403 VTAIL.n109 B 0.014483f
C404 VTAIL.n110 B 0.015335f
C405 VTAIL.n111 B 0.034233f
C406 VTAIL.n112 B 0.072501f
C407 VTAIL.n113 B 0.015335f
C408 VTAIL.n114 B 0.014483f
C409 VTAIL.n115 B 0.064877f
C410 VTAIL.n116 B 0.040479f
C411 VTAIL.n117 B 0.549304f
C412 VTAIL.t19 B 0.213627f
C413 VTAIL.t8 B 0.213627f
C414 VTAIL.n118 B 1.8074f
C415 VTAIL.n119 B 0.782065f
C416 VTAIL.t6 B 0.213627f
C417 VTAIL.t0 B 0.213627f
C418 VTAIL.n120 B 1.8074f
C419 VTAIL.n121 B 0.902603f
C420 VTAIL.n122 B 0.036975f
C421 VTAIL.n123 B 0.026953f
C422 VTAIL.n124 B 0.014483f
C423 VTAIL.n125 B 0.034233f
C424 VTAIL.n126 B 0.015335f
C425 VTAIL.n127 B 0.026953f
C426 VTAIL.n128 B 0.014909f
C427 VTAIL.n129 B 0.034233f
C428 VTAIL.n130 B 0.014483f
C429 VTAIL.n131 B 0.015335f
C430 VTAIL.n132 B 0.026953f
C431 VTAIL.n133 B 0.014483f
C432 VTAIL.n134 B 0.034233f
C433 VTAIL.n135 B 0.015335f
C434 VTAIL.n136 B 0.026953f
C435 VTAIL.n137 B 0.014483f
C436 VTAIL.n138 B 0.025675f
C437 VTAIL.n139 B 0.0242f
C438 VTAIL.t4 B 0.057533f
C439 VTAIL.n140 B 0.173944f
C440 VTAIL.n141 B 1.12354f
C441 VTAIL.n142 B 0.014483f
C442 VTAIL.n143 B 0.015335f
C443 VTAIL.n144 B 0.034233f
C444 VTAIL.n145 B 0.034233f
C445 VTAIL.n146 B 0.015335f
C446 VTAIL.n147 B 0.014483f
C447 VTAIL.n148 B 0.026953f
C448 VTAIL.n149 B 0.026953f
C449 VTAIL.n150 B 0.014483f
C450 VTAIL.n151 B 0.015335f
C451 VTAIL.n152 B 0.034233f
C452 VTAIL.n153 B 0.034233f
C453 VTAIL.n154 B 0.015335f
C454 VTAIL.n155 B 0.014483f
C455 VTAIL.n156 B 0.026953f
C456 VTAIL.n157 B 0.026953f
C457 VTAIL.n158 B 0.014483f
C458 VTAIL.n159 B 0.015335f
C459 VTAIL.n160 B 0.034233f
C460 VTAIL.n161 B 0.034233f
C461 VTAIL.n162 B 0.034233f
C462 VTAIL.n163 B 0.014909f
C463 VTAIL.n164 B 0.014483f
C464 VTAIL.n165 B 0.026953f
C465 VTAIL.n166 B 0.026953f
C466 VTAIL.n167 B 0.014483f
C467 VTAIL.n168 B 0.015335f
C468 VTAIL.n169 B 0.034233f
C469 VTAIL.n170 B 0.072501f
C470 VTAIL.n171 B 0.015335f
C471 VTAIL.n172 B 0.014483f
C472 VTAIL.n173 B 0.064877f
C473 VTAIL.n174 B 0.040479f
C474 VTAIL.n175 B 1.78689f
C475 VTAIL.n176 B 0.036975f
C476 VTAIL.n177 B 0.026953f
C477 VTAIL.n178 B 0.014483f
C478 VTAIL.n179 B 0.034233f
C479 VTAIL.n180 B 0.015335f
C480 VTAIL.n181 B 0.026953f
C481 VTAIL.n182 B 0.014909f
C482 VTAIL.n183 B 0.034233f
C483 VTAIL.n184 B 0.015335f
C484 VTAIL.n185 B 0.026953f
C485 VTAIL.n186 B 0.014483f
C486 VTAIL.n187 B 0.034233f
C487 VTAIL.n188 B 0.015335f
C488 VTAIL.n189 B 0.026953f
C489 VTAIL.n190 B 0.014483f
C490 VTAIL.n191 B 0.025675f
C491 VTAIL.n192 B 0.0242f
C492 VTAIL.t17 B 0.057533f
C493 VTAIL.n193 B 0.173944f
C494 VTAIL.n194 B 1.12354f
C495 VTAIL.n195 B 0.014483f
C496 VTAIL.n196 B 0.015335f
C497 VTAIL.n197 B 0.034233f
C498 VTAIL.n198 B 0.034233f
C499 VTAIL.n199 B 0.015335f
C500 VTAIL.n200 B 0.014483f
C501 VTAIL.n201 B 0.026953f
C502 VTAIL.n202 B 0.026953f
C503 VTAIL.n203 B 0.014483f
C504 VTAIL.n204 B 0.015335f
C505 VTAIL.n205 B 0.034233f
C506 VTAIL.n206 B 0.034233f
C507 VTAIL.n207 B 0.015335f
C508 VTAIL.n208 B 0.014483f
C509 VTAIL.n209 B 0.026953f
C510 VTAIL.n210 B 0.026953f
C511 VTAIL.n211 B 0.014483f
C512 VTAIL.n212 B 0.014483f
C513 VTAIL.n213 B 0.015335f
C514 VTAIL.n214 B 0.034233f
C515 VTAIL.n215 B 0.034233f
C516 VTAIL.n216 B 0.034233f
C517 VTAIL.n217 B 0.014909f
C518 VTAIL.n218 B 0.014483f
C519 VTAIL.n219 B 0.026953f
C520 VTAIL.n220 B 0.026953f
C521 VTAIL.n221 B 0.014483f
C522 VTAIL.n222 B 0.015335f
C523 VTAIL.n223 B 0.034233f
C524 VTAIL.n224 B 0.072501f
C525 VTAIL.n225 B 0.015335f
C526 VTAIL.n226 B 0.014483f
C527 VTAIL.n227 B 0.064877f
C528 VTAIL.n228 B 0.040479f
C529 VTAIL.n229 B 1.78689f
C530 VTAIL.t11 B 0.213627f
C531 VTAIL.t18 B 0.213627f
C532 VTAIL.n230 B 1.80739f
C533 VTAIL.n231 B 0.655548f
C534 VDD2.n0 B 0.03503f
C535 VDD2.n1 B 0.025535f
C536 VDD2.n2 B 0.013721f
C537 VDD2.n3 B 0.032432f
C538 VDD2.n4 B 0.014529f
C539 VDD2.n5 B 0.025535f
C540 VDD2.n6 B 0.014125f
C541 VDD2.n7 B 0.032432f
C542 VDD2.n8 B 0.014529f
C543 VDD2.n9 B 0.025535f
C544 VDD2.n10 B 0.013721f
C545 VDD2.n11 B 0.032432f
C546 VDD2.n12 B 0.014529f
C547 VDD2.n13 B 0.025535f
C548 VDD2.n14 B 0.013721f
C549 VDD2.n15 B 0.024324f
C550 VDD2.n16 B 0.022927f
C551 VDD2.t7 B 0.054507f
C552 VDD2.n17 B 0.164796f
C553 VDD2.n18 B 1.06445f
C554 VDD2.n19 B 0.013721f
C555 VDD2.n20 B 0.014529f
C556 VDD2.n21 B 0.032432f
C557 VDD2.n22 B 0.032432f
C558 VDD2.n23 B 0.014529f
C559 VDD2.n24 B 0.013721f
C560 VDD2.n25 B 0.025535f
C561 VDD2.n26 B 0.025535f
C562 VDD2.n27 B 0.013721f
C563 VDD2.n28 B 0.014529f
C564 VDD2.n29 B 0.032432f
C565 VDD2.n30 B 0.032432f
C566 VDD2.n31 B 0.014529f
C567 VDD2.n32 B 0.013721f
C568 VDD2.n33 B 0.025535f
C569 VDD2.n34 B 0.025535f
C570 VDD2.n35 B 0.013721f
C571 VDD2.n36 B 0.013721f
C572 VDD2.n37 B 0.014529f
C573 VDD2.n38 B 0.032432f
C574 VDD2.n39 B 0.032432f
C575 VDD2.n40 B 0.032432f
C576 VDD2.n41 B 0.014125f
C577 VDD2.n42 B 0.013721f
C578 VDD2.n43 B 0.025535f
C579 VDD2.n44 B 0.025535f
C580 VDD2.n45 B 0.013721f
C581 VDD2.n46 B 0.014529f
C582 VDD2.n47 B 0.032432f
C583 VDD2.n48 B 0.068688f
C584 VDD2.n49 B 0.014529f
C585 VDD2.n50 B 0.013721f
C586 VDD2.n51 B 0.061465f
C587 VDD2.n52 B 0.080506f
C588 VDD2.t4 B 0.202391f
C589 VDD2.t1 B 0.202391f
C590 VDD2.n53 B 1.78363f
C591 VDD2.n54 B 0.917129f
C592 VDD2.t0 B 0.202391f
C593 VDD2.t5 B 0.202391f
C594 VDD2.n55 B 1.81425f
C595 VDD2.n56 B 3.57234f
C596 VDD2.n57 B 0.03503f
C597 VDD2.n58 B 0.025535f
C598 VDD2.n59 B 0.013721f
C599 VDD2.n60 B 0.032432f
C600 VDD2.n61 B 0.014529f
C601 VDD2.n62 B 0.025535f
C602 VDD2.n63 B 0.014125f
C603 VDD2.n64 B 0.032432f
C604 VDD2.n65 B 0.013721f
C605 VDD2.n66 B 0.014529f
C606 VDD2.n67 B 0.025535f
C607 VDD2.n68 B 0.013721f
C608 VDD2.n69 B 0.032432f
C609 VDD2.n70 B 0.014529f
C610 VDD2.n71 B 0.025535f
C611 VDD2.n72 B 0.013721f
C612 VDD2.n73 B 0.024324f
C613 VDD2.n74 B 0.022927f
C614 VDD2.t2 B 0.054507f
C615 VDD2.n75 B 0.164796f
C616 VDD2.n76 B 1.06445f
C617 VDD2.n77 B 0.013721f
C618 VDD2.n78 B 0.014529f
C619 VDD2.n79 B 0.032432f
C620 VDD2.n80 B 0.032432f
C621 VDD2.n81 B 0.014529f
C622 VDD2.n82 B 0.013721f
C623 VDD2.n83 B 0.025535f
C624 VDD2.n84 B 0.025535f
C625 VDD2.n85 B 0.013721f
C626 VDD2.n86 B 0.014529f
C627 VDD2.n87 B 0.032432f
C628 VDD2.n88 B 0.032432f
C629 VDD2.n89 B 0.014529f
C630 VDD2.n90 B 0.013721f
C631 VDD2.n91 B 0.025535f
C632 VDD2.n92 B 0.025535f
C633 VDD2.n93 B 0.013721f
C634 VDD2.n94 B 0.014529f
C635 VDD2.n95 B 0.032432f
C636 VDD2.n96 B 0.032432f
C637 VDD2.n97 B 0.032432f
C638 VDD2.n98 B 0.014125f
C639 VDD2.n99 B 0.013721f
C640 VDD2.n100 B 0.025535f
C641 VDD2.n101 B 0.025535f
C642 VDD2.n102 B 0.013721f
C643 VDD2.n103 B 0.014529f
C644 VDD2.n104 B 0.032432f
C645 VDD2.n105 B 0.068688f
C646 VDD2.n106 B 0.014529f
C647 VDD2.n107 B 0.013721f
C648 VDD2.n108 B 0.061465f
C649 VDD2.n109 B 0.055963f
C650 VDD2.n110 B 3.34945f
C651 VDD2.t6 B 0.202391f
C652 VDD2.t3 B 0.202391f
C653 VDD2.n111 B 1.78363f
C654 VDD2.n112 B 0.594049f
C655 VDD2.t8 B 0.202391f
C656 VDD2.t9 B 0.202391f
C657 VDD2.n113 B 1.8142f
C658 VN.n0 B 0.031702f
C659 VN.t1 B 1.82285f
C660 VN.n1 B 0.031412f
C661 VN.n2 B 0.016854f
C662 VN.n3 B 0.031412f
C663 VN.n4 B 0.016854f
C664 VN.t0 B 1.82285f
C665 VN.n5 B 0.031412f
C666 VN.n6 B 0.016854f
C667 VN.n7 B 0.031412f
C668 VN.n8 B 0.016854f
C669 VN.t7 B 1.82285f
C670 VN.n9 B 0.031412f
C671 VN.n10 B 0.016854f
C672 VN.n11 B 0.03384f
C673 VN.n12 B 0.016854f
C674 VN.t6 B 1.82285f
C675 VN.n13 B 0.700053f
C676 VN.t2 B 2.09227f
C677 VN.n14 B 0.66636f
C678 VN.n15 B 0.226362f
C679 VN.n16 B 0.017764f
C680 VN.n17 B 0.031412f
C681 VN.n18 B 0.031412f
C682 VN.n19 B 0.016854f
C683 VN.n20 B 0.016854f
C684 VN.n21 B 0.016854f
C685 VN.n22 B 0.015686f
C686 VN.n23 B 0.031097f
C687 VN.n24 B 0.031412f
C688 VN.n25 B 0.016854f
C689 VN.n26 B 0.016854f
C690 VN.n27 B 0.016854f
C691 VN.n28 B 0.023658f
C692 VN.n29 B 0.644012f
C693 VN.n30 B 0.023658f
C694 VN.n31 B 0.031412f
C695 VN.n32 B 0.016854f
C696 VN.n33 B 0.016854f
C697 VN.n34 B 0.016854f
C698 VN.n35 B 0.031097f
C699 VN.n36 B 0.015686f
C700 VN.n37 B 0.03384f
C701 VN.n38 B 0.016854f
C702 VN.n39 B 0.016854f
C703 VN.n40 B 0.016854f
C704 VN.n41 B 0.031412f
C705 VN.n42 B 0.017764f
C706 VN.n43 B 0.644012f
C707 VN.n44 B 0.029551f
C708 VN.n45 B 0.016854f
C709 VN.n46 B 0.016854f
C710 VN.n47 B 0.016854f
C711 VN.n48 B 0.031412f
C712 VN.n49 B 0.022962f
C713 VN.n50 B 0.026249f
C714 VN.n51 B 0.016854f
C715 VN.n52 B 0.016854f
C716 VN.n53 B 0.016854f
C717 VN.n54 B 0.031412f
C718 VN.n55 B 0.02738f
C719 VN.n56 B 0.715599f
C720 VN.n57 B 0.05566f
C721 VN.n58 B 0.031702f
C722 VN.t5 B 1.82285f
C723 VN.n59 B 0.031412f
C724 VN.n60 B 0.016854f
C725 VN.n61 B 0.031412f
C726 VN.n62 B 0.016854f
C727 VN.t3 B 1.82285f
C728 VN.n63 B 0.031412f
C729 VN.n64 B 0.016854f
C730 VN.n65 B 0.031412f
C731 VN.n66 B 0.016854f
C732 VN.t9 B 1.82285f
C733 VN.n67 B 0.031412f
C734 VN.n68 B 0.016854f
C735 VN.n69 B 0.03384f
C736 VN.n70 B 0.016854f
C737 VN.t4 B 1.82285f
C738 VN.n71 B 0.700053f
C739 VN.t8 B 2.09227f
C740 VN.n72 B 0.66636f
C741 VN.n73 B 0.226362f
C742 VN.n74 B 0.017764f
C743 VN.n75 B 0.031412f
C744 VN.n76 B 0.031412f
C745 VN.n77 B 0.016854f
C746 VN.n78 B 0.016854f
C747 VN.n79 B 0.016854f
C748 VN.n80 B 0.015686f
C749 VN.n81 B 0.031097f
C750 VN.n82 B 0.031412f
C751 VN.n83 B 0.016854f
C752 VN.n84 B 0.016854f
C753 VN.n85 B 0.016854f
C754 VN.n86 B 0.023658f
C755 VN.n87 B 0.644012f
C756 VN.n88 B 0.023658f
C757 VN.n89 B 0.031412f
C758 VN.n90 B 0.016854f
C759 VN.n91 B 0.016854f
C760 VN.n92 B 0.016854f
C761 VN.n93 B 0.031097f
C762 VN.n94 B 0.015686f
C763 VN.n95 B 0.03384f
C764 VN.n96 B 0.016854f
C765 VN.n97 B 0.016854f
C766 VN.n98 B 0.016854f
C767 VN.n99 B 0.031412f
C768 VN.n100 B 0.017764f
C769 VN.n101 B 0.644012f
C770 VN.n102 B 0.029551f
C771 VN.n103 B 0.016854f
C772 VN.n104 B 0.016854f
C773 VN.n105 B 0.016854f
C774 VN.n106 B 0.031412f
C775 VN.n107 B 0.022962f
C776 VN.n108 B 0.026249f
C777 VN.n109 B 0.016854f
C778 VN.n110 B 0.016854f
C779 VN.n111 B 0.016854f
C780 VN.n112 B 0.031412f
C781 VN.n113 B 0.02738f
C782 VN.n114 B 0.715599f
C783 VN.n115 B 1.2435f
.ends

