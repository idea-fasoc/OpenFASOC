* NGSPICE file created from diff_pair_sample_0955.ext - technology: sky130A

.subckt diff_pair_sample_0955 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.1419 ps=1.19 w=0.86 l=3.09
X1 VDD1.t4 VP.t1 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0.1419 ps=1.19 w=0.86 l=3.09
X2 VDD1.t1 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.3354 ps=2.5 w=0.86 l=3.09
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0 ps=0 w=0.86 l=3.09
X4 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0 ps=0 w=0.86 l=3.09
X5 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0.1419 ps=1.19 w=0.86 l=3.09
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0 ps=0 w=0.86 l=3.09
X7 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.3354 ps=2.5 w=0.86 l=3.09
X8 VTAIL.t3 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.1419 ps=1.19 w=0.86 l=3.09
X9 VTAIL.t5 VN.t3 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.1419 ps=1.19 w=0.86 l=3.09
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0 ps=0 w=0.86 l=3.09
X11 VDD1.t3 VP.t3 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.3354 ps=2.5 w=0.86 l=3.09
X12 VDD1.t0 VP.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0.1419 ps=1.19 w=0.86 l=3.09
X13 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.3354 ps=2.5 w=0.86 l=3.09
X14 VTAIL.t6 VP.t5 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.1419 pd=1.19 as=0.1419 ps=1.19 w=0.86 l=3.09
X15 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.3354 pd=2.5 as=0.1419 ps=1.19 w=0.86 l=3.09
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n44 VP.n43 161.3
R7 VP.n42 VP.n1 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n39 VP.n2 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n36 VP.n3 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n4 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n5 161.3
R16 VP.n29 VP.n28 161.3
R17 VP.n27 VP.n6 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n24 VP.n23 69.5884
R20 VP.n45 VP.n0 69.5884
R21 VP.n22 VP.n7 69.5884
R22 VP.n30 VP.n29 56.5617
R23 VP.n41 VP.n2 56.5617
R24 VP.n18 VP.n9 56.5617
R25 VP.n12 VP.n11 49.5352
R26 VP.n23 VP.n22 42.3102
R27 VP.n11 VP.t4 40.1966
R28 VP.n25 VP.n6 24.5923
R29 VP.n29 VP.n6 24.5923
R30 VP.n31 VP.n30 24.5923
R31 VP.n31 VP.n4 24.5923
R32 VP.n35 VP.n4 24.5923
R33 VP.n36 VP.n35 24.5923
R34 VP.n37 VP.n36 24.5923
R35 VP.n37 VP.n2 24.5923
R36 VP.n42 VP.n41 24.5923
R37 VP.n43 VP.n42 24.5923
R38 VP.n19 VP.n18 24.5923
R39 VP.n20 VP.n19 24.5923
R40 VP.n13 VP.n12 24.5923
R41 VP.n14 VP.n13 24.5923
R42 VP.n14 VP.n9 24.5923
R43 VP.n25 VP.n24 20.6576
R44 VP.n43 VP.n0 20.6576
R45 VP.n20 VP.n7 20.6576
R46 VP.n35 VP.t0 6.70794
R47 VP.n24 VP.t1 6.70794
R48 VP.n0 VP.t2 6.70794
R49 VP.n12 VP.t5 6.70794
R50 VP.n7 VP.t3 6.70794
R51 VP.n11 VP.n10 3.87328
R52 VP.n22 VP.n21 0.354861
R53 VP.n26 VP.n23 0.354861
R54 VP.n45 VP.n44 0.354861
R55 VP VP.n45 0.267071
R56 VP.n15 VP.n10 0.189894
R57 VP.n16 VP.n15 0.189894
R58 VP.n17 VP.n16 0.189894
R59 VP.n17 VP.n8 0.189894
R60 VP.n21 VP.n8 0.189894
R61 VP.n27 VP.n26 0.189894
R62 VP.n28 VP.n27 0.189894
R63 VP.n28 VP.n5 0.189894
R64 VP.n32 VP.n5 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n34 VP.n3 0.189894
R68 VP.n38 VP.n3 0.189894
R69 VP.n39 VP.n38 0.189894
R70 VP.n40 VP.n39 0.189894
R71 VP.n40 VP.n1 0.189894
R72 VP.n44 VP.n1 0.189894
R73 VDD1 VDD1.t0 262.711
R74 VDD1.n1 VDD1.t4 262.596
R75 VDD1.n1 VDD1.n0 238.099
R76 VDD1.n3 VDD1.n2 237.417
R77 VDD1.n3 VDD1.n1 36.0957
R78 VDD1.n2 VDD1.t2 23.0238
R79 VDD1.n2 VDD1.t3 23.0238
R80 VDD1.n0 VDD1.t5 23.0238
R81 VDD1.n0 VDD1.t1 23.0238
R82 VDD1 VDD1.n3 0.679379
R83 VTAIL.n10 VTAIL.t8 243.762
R84 VTAIL.n7 VTAIL.t4 243.762
R85 VTAIL.n11 VTAIL.t0 243.762
R86 VTAIL.n2 VTAIL.t9 243.762
R87 VTAIL.n9 VTAIL.n8 220.738
R88 VTAIL.n6 VTAIL.n5 220.738
R89 VTAIL.n1 VTAIL.n0 220.738
R90 VTAIL.n4 VTAIL.n3 220.738
R91 VTAIL.n0 VTAIL.t1 23.0238
R92 VTAIL.n0 VTAIL.t3 23.0238
R93 VTAIL.n3 VTAIL.t10 23.0238
R94 VTAIL.n3 VTAIL.t11 23.0238
R95 VTAIL.n8 VTAIL.t7 23.0238
R96 VTAIL.n8 VTAIL.t6 23.0238
R97 VTAIL.n5 VTAIL.t2 23.0238
R98 VTAIL.n5 VTAIL.t5 23.0238
R99 VTAIL.n6 VTAIL.n4 19.0048
R100 VTAIL.n11 VTAIL.n10 16.0565
R101 VTAIL.n7 VTAIL.n6 2.94878
R102 VTAIL.n10 VTAIL.n9 2.94878
R103 VTAIL.n4 VTAIL.n2 2.94878
R104 VTAIL VTAIL.n11 2.15352
R105 VTAIL.n9 VTAIL.n7 1.94447
R106 VTAIL.n2 VTAIL.n1 1.94447
R107 VTAIL VTAIL.n1 0.795759
R108 B.n535 B.n534 585
R109 B.n536 B.n535 585
R110 B.n159 B.n104 585
R111 B.n158 B.n157 585
R112 B.n156 B.n155 585
R113 B.n154 B.n153 585
R114 B.n152 B.n151 585
R115 B.n150 B.n149 585
R116 B.n148 B.n147 585
R117 B.n146 B.n145 585
R118 B.n144 B.n143 585
R119 B.n142 B.n141 585
R120 B.n140 B.n139 585
R121 B.n138 B.n137 585
R122 B.n136 B.n135 585
R123 B.n134 B.n133 585
R124 B.n132 B.n131 585
R125 B.n130 B.n129 585
R126 B.n128 B.n127 585
R127 B.n125 B.n124 585
R128 B.n123 B.n122 585
R129 B.n121 B.n120 585
R130 B.n119 B.n118 585
R131 B.n117 B.n116 585
R132 B.n115 B.n114 585
R133 B.n113 B.n112 585
R134 B.n111 B.n110 585
R135 B.n89 B.n88 585
R136 B.n533 B.n90 585
R137 B.n537 B.n90 585
R138 B.n532 B.n531 585
R139 B.n531 B.n86 585
R140 B.n530 B.n85 585
R141 B.n543 B.n85 585
R142 B.n529 B.n84 585
R143 B.n544 B.n84 585
R144 B.n528 B.n83 585
R145 B.n545 B.n83 585
R146 B.n527 B.n526 585
R147 B.n526 B.n79 585
R148 B.n525 B.n78 585
R149 B.n551 B.n78 585
R150 B.n524 B.n77 585
R151 B.n552 B.n77 585
R152 B.n523 B.n76 585
R153 B.n553 B.n76 585
R154 B.n522 B.n521 585
R155 B.n521 B.n72 585
R156 B.n520 B.n71 585
R157 B.n559 B.n71 585
R158 B.n519 B.n70 585
R159 B.n560 B.n70 585
R160 B.n518 B.n69 585
R161 B.n561 B.n69 585
R162 B.n517 B.n516 585
R163 B.n516 B.n65 585
R164 B.n515 B.n64 585
R165 B.n567 B.n64 585
R166 B.n514 B.n63 585
R167 B.n568 B.n63 585
R168 B.n513 B.n62 585
R169 B.n569 B.n62 585
R170 B.n512 B.n511 585
R171 B.n511 B.n58 585
R172 B.n510 B.n57 585
R173 B.n575 B.n57 585
R174 B.n509 B.n56 585
R175 B.n576 B.n56 585
R176 B.n508 B.n55 585
R177 B.n577 B.n55 585
R178 B.n507 B.n506 585
R179 B.n506 B.n54 585
R180 B.n505 B.n50 585
R181 B.n583 B.n50 585
R182 B.n504 B.n49 585
R183 B.n584 B.n49 585
R184 B.n503 B.n48 585
R185 B.n585 B.n48 585
R186 B.n502 B.n501 585
R187 B.n501 B.n44 585
R188 B.n500 B.n43 585
R189 B.n591 B.n43 585
R190 B.n499 B.n42 585
R191 B.n592 B.n42 585
R192 B.n498 B.n41 585
R193 B.n593 B.n41 585
R194 B.n497 B.n496 585
R195 B.n496 B.n37 585
R196 B.n495 B.n36 585
R197 B.n599 B.n36 585
R198 B.n494 B.n35 585
R199 B.n600 B.n35 585
R200 B.n493 B.n34 585
R201 B.n601 B.n34 585
R202 B.n492 B.n491 585
R203 B.n491 B.n30 585
R204 B.n490 B.n29 585
R205 B.n607 B.n29 585
R206 B.n489 B.n28 585
R207 B.n608 B.n28 585
R208 B.n488 B.n27 585
R209 B.n609 B.n27 585
R210 B.n487 B.n486 585
R211 B.n486 B.n23 585
R212 B.n485 B.n22 585
R213 B.n615 B.n22 585
R214 B.n484 B.n21 585
R215 B.n616 B.n21 585
R216 B.n483 B.n20 585
R217 B.n617 B.n20 585
R218 B.n482 B.n481 585
R219 B.n481 B.n19 585
R220 B.n480 B.n15 585
R221 B.n623 B.n15 585
R222 B.n479 B.n14 585
R223 B.n624 B.n14 585
R224 B.n478 B.n13 585
R225 B.n625 B.n13 585
R226 B.n477 B.n476 585
R227 B.n476 B.n12 585
R228 B.n475 B.n474 585
R229 B.n475 B.n8 585
R230 B.n473 B.n7 585
R231 B.n632 B.n7 585
R232 B.n472 B.n6 585
R233 B.n633 B.n6 585
R234 B.n471 B.n5 585
R235 B.n634 B.n5 585
R236 B.n470 B.n469 585
R237 B.n469 B.n4 585
R238 B.n468 B.n160 585
R239 B.n468 B.n467 585
R240 B.n458 B.n161 585
R241 B.n162 B.n161 585
R242 B.n460 B.n459 585
R243 B.n461 B.n460 585
R244 B.n457 B.n167 585
R245 B.n167 B.n166 585
R246 B.n456 B.n455 585
R247 B.n455 B.n454 585
R248 B.n169 B.n168 585
R249 B.n447 B.n169 585
R250 B.n446 B.n445 585
R251 B.n448 B.n446 585
R252 B.n444 B.n174 585
R253 B.n174 B.n173 585
R254 B.n443 B.n442 585
R255 B.n442 B.n441 585
R256 B.n176 B.n175 585
R257 B.n177 B.n176 585
R258 B.n434 B.n433 585
R259 B.n435 B.n434 585
R260 B.n432 B.n182 585
R261 B.n182 B.n181 585
R262 B.n431 B.n430 585
R263 B.n430 B.n429 585
R264 B.n184 B.n183 585
R265 B.n185 B.n184 585
R266 B.n422 B.n421 585
R267 B.n423 B.n422 585
R268 B.n420 B.n189 585
R269 B.n193 B.n189 585
R270 B.n419 B.n418 585
R271 B.n418 B.n417 585
R272 B.n191 B.n190 585
R273 B.n192 B.n191 585
R274 B.n410 B.n409 585
R275 B.n411 B.n410 585
R276 B.n408 B.n198 585
R277 B.n198 B.n197 585
R278 B.n407 B.n406 585
R279 B.n406 B.n405 585
R280 B.n200 B.n199 585
R281 B.n201 B.n200 585
R282 B.n398 B.n397 585
R283 B.n399 B.n398 585
R284 B.n396 B.n206 585
R285 B.n206 B.n205 585
R286 B.n395 B.n394 585
R287 B.n394 B.n393 585
R288 B.n208 B.n207 585
R289 B.n386 B.n208 585
R290 B.n385 B.n384 585
R291 B.n387 B.n385 585
R292 B.n383 B.n213 585
R293 B.n213 B.n212 585
R294 B.n382 B.n381 585
R295 B.n381 B.n380 585
R296 B.n215 B.n214 585
R297 B.n216 B.n215 585
R298 B.n373 B.n372 585
R299 B.n374 B.n373 585
R300 B.n371 B.n221 585
R301 B.n221 B.n220 585
R302 B.n370 B.n369 585
R303 B.n369 B.n368 585
R304 B.n223 B.n222 585
R305 B.n224 B.n223 585
R306 B.n361 B.n360 585
R307 B.n362 B.n361 585
R308 B.n359 B.n229 585
R309 B.n229 B.n228 585
R310 B.n358 B.n357 585
R311 B.n357 B.n356 585
R312 B.n231 B.n230 585
R313 B.n232 B.n231 585
R314 B.n349 B.n348 585
R315 B.n350 B.n349 585
R316 B.n347 B.n237 585
R317 B.n237 B.n236 585
R318 B.n346 B.n345 585
R319 B.n345 B.n344 585
R320 B.n239 B.n238 585
R321 B.n240 B.n239 585
R322 B.n337 B.n336 585
R323 B.n338 B.n337 585
R324 B.n335 B.n245 585
R325 B.n245 B.n244 585
R326 B.n334 B.n333 585
R327 B.n333 B.n332 585
R328 B.n247 B.n246 585
R329 B.n248 B.n247 585
R330 B.n325 B.n324 585
R331 B.n326 B.n325 585
R332 B.n251 B.n250 585
R333 B.n273 B.n272 585
R334 B.n274 B.n270 585
R335 B.n270 B.n252 585
R336 B.n276 B.n275 585
R337 B.n278 B.n269 585
R338 B.n281 B.n280 585
R339 B.n282 B.n268 585
R340 B.n284 B.n283 585
R341 B.n286 B.n267 585
R342 B.n289 B.n288 585
R343 B.n290 B.n263 585
R344 B.n292 B.n291 585
R345 B.n294 B.n262 585
R346 B.n297 B.n296 585
R347 B.n298 B.n261 585
R348 B.n300 B.n299 585
R349 B.n302 B.n260 585
R350 B.n305 B.n304 585
R351 B.n307 B.n257 585
R352 B.n309 B.n308 585
R353 B.n311 B.n256 585
R354 B.n314 B.n313 585
R355 B.n315 B.n255 585
R356 B.n317 B.n316 585
R357 B.n319 B.n254 585
R358 B.n322 B.n321 585
R359 B.n323 B.n253 585
R360 B.n328 B.n327 585
R361 B.n327 B.n326 585
R362 B.n329 B.n249 585
R363 B.n249 B.n248 585
R364 B.n331 B.n330 585
R365 B.n332 B.n331 585
R366 B.n243 B.n242 585
R367 B.n244 B.n243 585
R368 B.n340 B.n339 585
R369 B.n339 B.n338 585
R370 B.n341 B.n241 585
R371 B.n241 B.n240 585
R372 B.n343 B.n342 585
R373 B.n344 B.n343 585
R374 B.n235 B.n234 585
R375 B.n236 B.n235 585
R376 B.n352 B.n351 585
R377 B.n351 B.n350 585
R378 B.n353 B.n233 585
R379 B.n233 B.n232 585
R380 B.n355 B.n354 585
R381 B.n356 B.n355 585
R382 B.n227 B.n226 585
R383 B.n228 B.n227 585
R384 B.n364 B.n363 585
R385 B.n363 B.n362 585
R386 B.n365 B.n225 585
R387 B.n225 B.n224 585
R388 B.n367 B.n366 585
R389 B.n368 B.n367 585
R390 B.n219 B.n218 585
R391 B.n220 B.n219 585
R392 B.n376 B.n375 585
R393 B.n375 B.n374 585
R394 B.n377 B.n217 585
R395 B.n217 B.n216 585
R396 B.n379 B.n378 585
R397 B.n380 B.n379 585
R398 B.n211 B.n210 585
R399 B.n212 B.n211 585
R400 B.n389 B.n388 585
R401 B.n388 B.n387 585
R402 B.n390 B.n209 585
R403 B.n386 B.n209 585
R404 B.n392 B.n391 585
R405 B.n393 B.n392 585
R406 B.n204 B.n203 585
R407 B.n205 B.n204 585
R408 B.n401 B.n400 585
R409 B.n400 B.n399 585
R410 B.n402 B.n202 585
R411 B.n202 B.n201 585
R412 B.n404 B.n403 585
R413 B.n405 B.n404 585
R414 B.n196 B.n195 585
R415 B.n197 B.n196 585
R416 B.n413 B.n412 585
R417 B.n412 B.n411 585
R418 B.n414 B.n194 585
R419 B.n194 B.n192 585
R420 B.n416 B.n415 585
R421 B.n417 B.n416 585
R422 B.n188 B.n187 585
R423 B.n193 B.n188 585
R424 B.n425 B.n424 585
R425 B.n424 B.n423 585
R426 B.n426 B.n186 585
R427 B.n186 B.n185 585
R428 B.n428 B.n427 585
R429 B.n429 B.n428 585
R430 B.n180 B.n179 585
R431 B.n181 B.n180 585
R432 B.n437 B.n436 585
R433 B.n436 B.n435 585
R434 B.n438 B.n178 585
R435 B.n178 B.n177 585
R436 B.n440 B.n439 585
R437 B.n441 B.n440 585
R438 B.n172 B.n171 585
R439 B.n173 B.n172 585
R440 B.n450 B.n449 585
R441 B.n449 B.n448 585
R442 B.n451 B.n170 585
R443 B.n447 B.n170 585
R444 B.n453 B.n452 585
R445 B.n454 B.n453 585
R446 B.n165 B.n164 585
R447 B.n166 B.n165 585
R448 B.n463 B.n462 585
R449 B.n462 B.n461 585
R450 B.n464 B.n163 585
R451 B.n163 B.n162 585
R452 B.n466 B.n465 585
R453 B.n467 B.n466 585
R454 B.n3 B.n0 585
R455 B.n4 B.n3 585
R456 B.n631 B.n1 585
R457 B.n632 B.n631 585
R458 B.n630 B.n629 585
R459 B.n630 B.n8 585
R460 B.n628 B.n9 585
R461 B.n12 B.n9 585
R462 B.n627 B.n626 585
R463 B.n626 B.n625 585
R464 B.n11 B.n10 585
R465 B.n624 B.n11 585
R466 B.n622 B.n621 585
R467 B.n623 B.n622 585
R468 B.n620 B.n16 585
R469 B.n19 B.n16 585
R470 B.n619 B.n618 585
R471 B.n618 B.n617 585
R472 B.n18 B.n17 585
R473 B.n616 B.n18 585
R474 B.n614 B.n613 585
R475 B.n615 B.n614 585
R476 B.n612 B.n24 585
R477 B.n24 B.n23 585
R478 B.n611 B.n610 585
R479 B.n610 B.n609 585
R480 B.n26 B.n25 585
R481 B.n608 B.n26 585
R482 B.n606 B.n605 585
R483 B.n607 B.n606 585
R484 B.n604 B.n31 585
R485 B.n31 B.n30 585
R486 B.n603 B.n602 585
R487 B.n602 B.n601 585
R488 B.n33 B.n32 585
R489 B.n600 B.n33 585
R490 B.n598 B.n597 585
R491 B.n599 B.n598 585
R492 B.n596 B.n38 585
R493 B.n38 B.n37 585
R494 B.n595 B.n594 585
R495 B.n594 B.n593 585
R496 B.n40 B.n39 585
R497 B.n592 B.n40 585
R498 B.n590 B.n589 585
R499 B.n591 B.n590 585
R500 B.n588 B.n45 585
R501 B.n45 B.n44 585
R502 B.n587 B.n586 585
R503 B.n586 B.n585 585
R504 B.n47 B.n46 585
R505 B.n584 B.n47 585
R506 B.n582 B.n581 585
R507 B.n583 B.n582 585
R508 B.n580 B.n51 585
R509 B.n54 B.n51 585
R510 B.n579 B.n578 585
R511 B.n578 B.n577 585
R512 B.n53 B.n52 585
R513 B.n576 B.n53 585
R514 B.n574 B.n573 585
R515 B.n575 B.n574 585
R516 B.n572 B.n59 585
R517 B.n59 B.n58 585
R518 B.n571 B.n570 585
R519 B.n570 B.n569 585
R520 B.n61 B.n60 585
R521 B.n568 B.n61 585
R522 B.n566 B.n565 585
R523 B.n567 B.n566 585
R524 B.n564 B.n66 585
R525 B.n66 B.n65 585
R526 B.n563 B.n562 585
R527 B.n562 B.n561 585
R528 B.n68 B.n67 585
R529 B.n560 B.n68 585
R530 B.n558 B.n557 585
R531 B.n559 B.n558 585
R532 B.n556 B.n73 585
R533 B.n73 B.n72 585
R534 B.n555 B.n554 585
R535 B.n554 B.n553 585
R536 B.n75 B.n74 585
R537 B.n552 B.n75 585
R538 B.n550 B.n549 585
R539 B.n551 B.n550 585
R540 B.n548 B.n80 585
R541 B.n80 B.n79 585
R542 B.n547 B.n546 585
R543 B.n546 B.n545 585
R544 B.n82 B.n81 585
R545 B.n544 B.n82 585
R546 B.n542 B.n541 585
R547 B.n543 B.n542 585
R548 B.n540 B.n87 585
R549 B.n87 B.n86 585
R550 B.n539 B.n538 585
R551 B.n538 B.n537 585
R552 B.n635 B.n634 585
R553 B.n633 B.n2 585
R554 B.n538 B.n89 497.305
R555 B.n535 B.n90 497.305
R556 B.n325 B.n253 497.305
R557 B.n327 B.n251 497.305
R558 B.n108 B.t18 300.726
R559 B.n105 B.t12 300.726
R560 B.n258 B.t9 300.726
R561 B.n264 B.t16 300.726
R562 B.n536 B.n103 256.663
R563 B.n536 B.n102 256.663
R564 B.n536 B.n101 256.663
R565 B.n536 B.n100 256.663
R566 B.n536 B.n99 256.663
R567 B.n536 B.n98 256.663
R568 B.n536 B.n97 256.663
R569 B.n536 B.n96 256.663
R570 B.n536 B.n95 256.663
R571 B.n536 B.n94 256.663
R572 B.n536 B.n93 256.663
R573 B.n536 B.n92 256.663
R574 B.n536 B.n91 256.663
R575 B.n271 B.n252 256.663
R576 B.n277 B.n252 256.663
R577 B.n279 B.n252 256.663
R578 B.n285 B.n252 256.663
R579 B.n287 B.n252 256.663
R580 B.n293 B.n252 256.663
R581 B.n295 B.n252 256.663
R582 B.n301 B.n252 256.663
R583 B.n303 B.n252 256.663
R584 B.n310 B.n252 256.663
R585 B.n312 B.n252 256.663
R586 B.n318 B.n252 256.663
R587 B.n320 B.n252 256.663
R588 B.n637 B.n636 256.663
R589 B.n109 B.t19 234.399
R590 B.n106 B.t13 234.399
R591 B.n259 B.t8 234.399
R592 B.n265 B.t15 234.399
R593 B.n108 B.t17 209.549
R594 B.n105 B.t10 209.549
R595 B.n258 B.t6 209.549
R596 B.n264 B.t14 209.549
R597 B.n326 B.n252 202.608
R598 B.n537 B.n536 202.608
R599 B.n112 B.n111 163.367
R600 B.n116 B.n115 163.367
R601 B.n120 B.n119 163.367
R602 B.n124 B.n123 163.367
R603 B.n129 B.n128 163.367
R604 B.n133 B.n132 163.367
R605 B.n137 B.n136 163.367
R606 B.n141 B.n140 163.367
R607 B.n145 B.n144 163.367
R608 B.n149 B.n148 163.367
R609 B.n153 B.n152 163.367
R610 B.n157 B.n156 163.367
R611 B.n535 B.n104 163.367
R612 B.n325 B.n247 163.367
R613 B.n333 B.n247 163.367
R614 B.n333 B.n245 163.367
R615 B.n337 B.n245 163.367
R616 B.n337 B.n239 163.367
R617 B.n345 B.n239 163.367
R618 B.n345 B.n237 163.367
R619 B.n349 B.n237 163.367
R620 B.n349 B.n231 163.367
R621 B.n357 B.n231 163.367
R622 B.n357 B.n229 163.367
R623 B.n361 B.n229 163.367
R624 B.n361 B.n223 163.367
R625 B.n369 B.n223 163.367
R626 B.n369 B.n221 163.367
R627 B.n373 B.n221 163.367
R628 B.n373 B.n215 163.367
R629 B.n381 B.n215 163.367
R630 B.n381 B.n213 163.367
R631 B.n385 B.n213 163.367
R632 B.n385 B.n208 163.367
R633 B.n394 B.n208 163.367
R634 B.n394 B.n206 163.367
R635 B.n398 B.n206 163.367
R636 B.n398 B.n200 163.367
R637 B.n406 B.n200 163.367
R638 B.n406 B.n198 163.367
R639 B.n410 B.n198 163.367
R640 B.n410 B.n191 163.367
R641 B.n418 B.n191 163.367
R642 B.n418 B.n189 163.367
R643 B.n422 B.n189 163.367
R644 B.n422 B.n184 163.367
R645 B.n430 B.n184 163.367
R646 B.n430 B.n182 163.367
R647 B.n434 B.n182 163.367
R648 B.n434 B.n176 163.367
R649 B.n442 B.n176 163.367
R650 B.n442 B.n174 163.367
R651 B.n446 B.n174 163.367
R652 B.n446 B.n169 163.367
R653 B.n455 B.n169 163.367
R654 B.n455 B.n167 163.367
R655 B.n460 B.n167 163.367
R656 B.n460 B.n161 163.367
R657 B.n468 B.n161 163.367
R658 B.n469 B.n468 163.367
R659 B.n469 B.n5 163.367
R660 B.n6 B.n5 163.367
R661 B.n7 B.n6 163.367
R662 B.n475 B.n7 163.367
R663 B.n476 B.n475 163.367
R664 B.n476 B.n13 163.367
R665 B.n14 B.n13 163.367
R666 B.n15 B.n14 163.367
R667 B.n481 B.n15 163.367
R668 B.n481 B.n20 163.367
R669 B.n21 B.n20 163.367
R670 B.n22 B.n21 163.367
R671 B.n486 B.n22 163.367
R672 B.n486 B.n27 163.367
R673 B.n28 B.n27 163.367
R674 B.n29 B.n28 163.367
R675 B.n491 B.n29 163.367
R676 B.n491 B.n34 163.367
R677 B.n35 B.n34 163.367
R678 B.n36 B.n35 163.367
R679 B.n496 B.n36 163.367
R680 B.n496 B.n41 163.367
R681 B.n42 B.n41 163.367
R682 B.n43 B.n42 163.367
R683 B.n501 B.n43 163.367
R684 B.n501 B.n48 163.367
R685 B.n49 B.n48 163.367
R686 B.n50 B.n49 163.367
R687 B.n506 B.n50 163.367
R688 B.n506 B.n55 163.367
R689 B.n56 B.n55 163.367
R690 B.n57 B.n56 163.367
R691 B.n511 B.n57 163.367
R692 B.n511 B.n62 163.367
R693 B.n63 B.n62 163.367
R694 B.n64 B.n63 163.367
R695 B.n516 B.n64 163.367
R696 B.n516 B.n69 163.367
R697 B.n70 B.n69 163.367
R698 B.n71 B.n70 163.367
R699 B.n521 B.n71 163.367
R700 B.n521 B.n76 163.367
R701 B.n77 B.n76 163.367
R702 B.n78 B.n77 163.367
R703 B.n526 B.n78 163.367
R704 B.n526 B.n83 163.367
R705 B.n84 B.n83 163.367
R706 B.n85 B.n84 163.367
R707 B.n531 B.n85 163.367
R708 B.n531 B.n90 163.367
R709 B.n272 B.n270 163.367
R710 B.n276 B.n270 163.367
R711 B.n280 B.n278 163.367
R712 B.n284 B.n268 163.367
R713 B.n288 B.n286 163.367
R714 B.n292 B.n263 163.367
R715 B.n296 B.n294 163.367
R716 B.n300 B.n261 163.367
R717 B.n304 B.n302 163.367
R718 B.n309 B.n257 163.367
R719 B.n313 B.n311 163.367
R720 B.n317 B.n255 163.367
R721 B.n321 B.n319 163.367
R722 B.n327 B.n249 163.367
R723 B.n331 B.n249 163.367
R724 B.n331 B.n243 163.367
R725 B.n339 B.n243 163.367
R726 B.n339 B.n241 163.367
R727 B.n343 B.n241 163.367
R728 B.n343 B.n235 163.367
R729 B.n351 B.n235 163.367
R730 B.n351 B.n233 163.367
R731 B.n355 B.n233 163.367
R732 B.n355 B.n227 163.367
R733 B.n363 B.n227 163.367
R734 B.n363 B.n225 163.367
R735 B.n367 B.n225 163.367
R736 B.n367 B.n219 163.367
R737 B.n375 B.n219 163.367
R738 B.n375 B.n217 163.367
R739 B.n379 B.n217 163.367
R740 B.n379 B.n211 163.367
R741 B.n388 B.n211 163.367
R742 B.n388 B.n209 163.367
R743 B.n392 B.n209 163.367
R744 B.n392 B.n204 163.367
R745 B.n400 B.n204 163.367
R746 B.n400 B.n202 163.367
R747 B.n404 B.n202 163.367
R748 B.n404 B.n196 163.367
R749 B.n412 B.n196 163.367
R750 B.n412 B.n194 163.367
R751 B.n416 B.n194 163.367
R752 B.n416 B.n188 163.367
R753 B.n424 B.n188 163.367
R754 B.n424 B.n186 163.367
R755 B.n428 B.n186 163.367
R756 B.n428 B.n180 163.367
R757 B.n436 B.n180 163.367
R758 B.n436 B.n178 163.367
R759 B.n440 B.n178 163.367
R760 B.n440 B.n172 163.367
R761 B.n449 B.n172 163.367
R762 B.n449 B.n170 163.367
R763 B.n453 B.n170 163.367
R764 B.n453 B.n165 163.367
R765 B.n462 B.n165 163.367
R766 B.n462 B.n163 163.367
R767 B.n466 B.n163 163.367
R768 B.n466 B.n3 163.367
R769 B.n635 B.n3 163.367
R770 B.n631 B.n2 163.367
R771 B.n631 B.n630 163.367
R772 B.n630 B.n9 163.367
R773 B.n626 B.n9 163.367
R774 B.n626 B.n11 163.367
R775 B.n622 B.n11 163.367
R776 B.n622 B.n16 163.367
R777 B.n618 B.n16 163.367
R778 B.n618 B.n18 163.367
R779 B.n614 B.n18 163.367
R780 B.n614 B.n24 163.367
R781 B.n610 B.n24 163.367
R782 B.n610 B.n26 163.367
R783 B.n606 B.n26 163.367
R784 B.n606 B.n31 163.367
R785 B.n602 B.n31 163.367
R786 B.n602 B.n33 163.367
R787 B.n598 B.n33 163.367
R788 B.n598 B.n38 163.367
R789 B.n594 B.n38 163.367
R790 B.n594 B.n40 163.367
R791 B.n590 B.n40 163.367
R792 B.n590 B.n45 163.367
R793 B.n586 B.n45 163.367
R794 B.n586 B.n47 163.367
R795 B.n582 B.n47 163.367
R796 B.n582 B.n51 163.367
R797 B.n578 B.n51 163.367
R798 B.n578 B.n53 163.367
R799 B.n574 B.n53 163.367
R800 B.n574 B.n59 163.367
R801 B.n570 B.n59 163.367
R802 B.n570 B.n61 163.367
R803 B.n566 B.n61 163.367
R804 B.n566 B.n66 163.367
R805 B.n562 B.n66 163.367
R806 B.n562 B.n68 163.367
R807 B.n558 B.n68 163.367
R808 B.n558 B.n73 163.367
R809 B.n554 B.n73 163.367
R810 B.n554 B.n75 163.367
R811 B.n550 B.n75 163.367
R812 B.n550 B.n80 163.367
R813 B.n546 B.n80 163.367
R814 B.n546 B.n82 163.367
R815 B.n542 B.n82 163.367
R816 B.n542 B.n87 163.367
R817 B.n538 B.n87 163.367
R818 B.n326 B.n248 121.924
R819 B.n332 B.n248 121.924
R820 B.n332 B.n244 121.924
R821 B.n338 B.n244 121.924
R822 B.n338 B.n240 121.924
R823 B.n344 B.n240 121.924
R824 B.n344 B.n236 121.924
R825 B.n350 B.n236 121.924
R826 B.n356 B.n232 121.924
R827 B.n356 B.n228 121.924
R828 B.n362 B.n228 121.924
R829 B.n362 B.n224 121.924
R830 B.n368 B.n224 121.924
R831 B.n368 B.n220 121.924
R832 B.n374 B.n220 121.924
R833 B.n374 B.n216 121.924
R834 B.n380 B.n216 121.924
R835 B.n380 B.n212 121.924
R836 B.n387 B.n212 121.924
R837 B.n387 B.n386 121.924
R838 B.n393 B.n205 121.924
R839 B.n399 B.n205 121.924
R840 B.n399 B.n201 121.924
R841 B.n405 B.n201 121.924
R842 B.n405 B.n197 121.924
R843 B.n411 B.n197 121.924
R844 B.n411 B.n192 121.924
R845 B.n417 B.n192 121.924
R846 B.n417 B.n193 121.924
R847 B.n423 B.n185 121.924
R848 B.n429 B.n185 121.924
R849 B.n429 B.n181 121.924
R850 B.n435 B.n181 121.924
R851 B.n435 B.n177 121.924
R852 B.n441 B.n177 121.924
R853 B.n441 B.n173 121.924
R854 B.n448 B.n173 121.924
R855 B.n448 B.n447 121.924
R856 B.n454 B.n166 121.924
R857 B.n461 B.n166 121.924
R858 B.n461 B.n162 121.924
R859 B.n467 B.n162 121.924
R860 B.n467 B.n4 121.924
R861 B.n634 B.n4 121.924
R862 B.n634 B.n633 121.924
R863 B.n633 B.n632 121.924
R864 B.n632 B.n8 121.924
R865 B.n12 B.n8 121.924
R866 B.n625 B.n12 121.924
R867 B.n625 B.n624 121.924
R868 B.n624 B.n623 121.924
R869 B.n617 B.n19 121.924
R870 B.n617 B.n616 121.924
R871 B.n616 B.n615 121.924
R872 B.n615 B.n23 121.924
R873 B.n609 B.n23 121.924
R874 B.n609 B.n608 121.924
R875 B.n608 B.n607 121.924
R876 B.n607 B.n30 121.924
R877 B.n601 B.n30 121.924
R878 B.n600 B.n599 121.924
R879 B.n599 B.n37 121.924
R880 B.n593 B.n37 121.924
R881 B.n593 B.n592 121.924
R882 B.n592 B.n591 121.924
R883 B.n591 B.n44 121.924
R884 B.n585 B.n44 121.924
R885 B.n585 B.n584 121.924
R886 B.n584 B.n583 121.924
R887 B.n577 B.n54 121.924
R888 B.n577 B.n576 121.924
R889 B.n576 B.n575 121.924
R890 B.n575 B.n58 121.924
R891 B.n569 B.n58 121.924
R892 B.n569 B.n568 121.924
R893 B.n568 B.n567 121.924
R894 B.n567 B.n65 121.924
R895 B.n561 B.n65 121.924
R896 B.n561 B.n560 121.924
R897 B.n560 B.n559 121.924
R898 B.n559 B.n72 121.924
R899 B.n553 B.n552 121.924
R900 B.n552 B.n551 121.924
R901 B.n551 B.n79 121.924
R902 B.n545 B.n79 121.924
R903 B.n545 B.n544 121.924
R904 B.n544 B.n543 121.924
R905 B.n543 B.n86 121.924
R906 B.n537 B.n86 121.924
R907 B.n447 B.t4 105.787
R908 B.n19 B.t1 105.787
R909 B.n193 B.t5 98.615
R910 B.t3 B.n600 98.615
R911 B.n386 B.t2 91.443
R912 B.n54 B.t0 91.443
R913 B.n91 B.n89 71.676
R914 B.n112 B.n92 71.676
R915 B.n116 B.n93 71.676
R916 B.n120 B.n94 71.676
R917 B.n124 B.n95 71.676
R918 B.n129 B.n96 71.676
R919 B.n133 B.n97 71.676
R920 B.n137 B.n98 71.676
R921 B.n141 B.n99 71.676
R922 B.n145 B.n100 71.676
R923 B.n149 B.n101 71.676
R924 B.n153 B.n102 71.676
R925 B.n157 B.n103 71.676
R926 B.n104 B.n103 71.676
R927 B.n156 B.n102 71.676
R928 B.n152 B.n101 71.676
R929 B.n148 B.n100 71.676
R930 B.n144 B.n99 71.676
R931 B.n140 B.n98 71.676
R932 B.n136 B.n97 71.676
R933 B.n132 B.n96 71.676
R934 B.n128 B.n95 71.676
R935 B.n123 B.n94 71.676
R936 B.n119 B.n93 71.676
R937 B.n115 B.n92 71.676
R938 B.n111 B.n91 71.676
R939 B.n271 B.n251 71.676
R940 B.n277 B.n276 71.676
R941 B.n280 B.n279 71.676
R942 B.n285 B.n284 71.676
R943 B.n288 B.n287 71.676
R944 B.n293 B.n292 71.676
R945 B.n296 B.n295 71.676
R946 B.n301 B.n300 71.676
R947 B.n304 B.n303 71.676
R948 B.n310 B.n309 71.676
R949 B.n313 B.n312 71.676
R950 B.n318 B.n317 71.676
R951 B.n321 B.n320 71.676
R952 B.n272 B.n271 71.676
R953 B.n278 B.n277 71.676
R954 B.n279 B.n268 71.676
R955 B.n286 B.n285 71.676
R956 B.n287 B.n263 71.676
R957 B.n294 B.n293 71.676
R958 B.n295 B.n261 71.676
R959 B.n302 B.n301 71.676
R960 B.n303 B.n257 71.676
R961 B.n311 B.n310 71.676
R962 B.n312 B.n255 71.676
R963 B.n319 B.n318 71.676
R964 B.n320 B.n253 71.676
R965 B.n636 B.n635 71.676
R966 B.n636 B.n2 71.676
R967 B.n109 B.n108 66.3278
R968 B.n106 B.n105 66.3278
R969 B.n259 B.n258 66.3278
R970 B.n265 B.n264 66.3278
R971 B.t7 B.n232 62.7552
R972 B.t11 B.n72 62.7552
R973 B.n126 B.n109 59.5399
R974 B.n107 B.n106 59.5399
R975 B.n306 B.n259 59.5399
R976 B.n266 B.n265 59.5399
R977 B.n350 B.t7 59.1692
R978 B.n553 B.t11 59.1692
R979 B.n328 B.n250 32.3127
R980 B.n324 B.n323 32.3127
R981 B.n534 B.n533 32.3127
R982 B.n539 B.n88 32.3127
R983 B.n393 B.t2 30.4813
R984 B.n583 B.t0 30.4813
R985 B.n423 B.t5 23.3094
R986 B.n601 B.t3 23.3094
R987 B B.n637 18.0485
R988 B.n454 B.t4 16.1374
R989 B.n623 B.t1 16.1374
R990 B.n329 B.n328 10.6151
R991 B.n330 B.n329 10.6151
R992 B.n330 B.n242 10.6151
R993 B.n340 B.n242 10.6151
R994 B.n341 B.n340 10.6151
R995 B.n342 B.n341 10.6151
R996 B.n342 B.n234 10.6151
R997 B.n352 B.n234 10.6151
R998 B.n353 B.n352 10.6151
R999 B.n354 B.n353 10.6151
R1000 B.n354 B.n226 10.6151
R1001 B.n364 B.n226 10.6151
R1002 B.n365 B.n364 10.6151
R1003 B.n366 B.n365 10.6151
R1004 B.n366 B.n218 10.6151
R1005 B.n376 B.n218 10.6151
R1006 B.n377 B.n376 10.6151
R1007 B.n378 B.n377 10.6151
R1008 B.n378 B.n210 10.6151
R1009 B.n389 B.n210 10.6151
R1010 B.n390 B.n389 10.6151
R1011 B.n391 B.n390 10.6151
R1012 B.n391 B.n203 10.6151
R1013 B.n401 B.n203 10.6151
R1014 B.n402 B.n401 10.6151
R1015 B.n403 B.n402 10.6151
R1016 B.n403 B.n195 10.6151
R1017 B.n413 B.n195 10.6151
R1018 B.n414 B.n413 10.6151
R1019 B.n415 B.n414 10.6151
R1020 B.n415 B.n187 10.6151
R1021 B.n425 B.n187 10.6151
R1022 B.n426 B.n425 10.6151
R1023 B.n427 B.n426 10.6151
R1024 B.n427 B.n179 10.6151
R1025 B.n437 B.n179 10.6151
R1026 B.n438 B.n437 10.6151
R1027 B.n439 B.n438 10.6151
R1028 B.n439 B.n171 10.6151
R1029 B.n450 B.n171 10.6151
R1030 B.n451 B.n450 10.6151
R1031 B.n452 B.n451 10.6151
R1032 B.n452 B.n164 10.6151
R1033 B.n463 B.n164 10.6151
R1034 B.n464 B.n463 10.6151
R1035 B.n465 B.n464 10.6151
R1036 B.n465 B.n0 10.6151
R1037 B.n273 B.n250 10.6151
R1038 B.n274 B.n273 10.6151
R1039 B.n275 B.n274 10.6151
R1040 B.n275 B.n269 10.6151
R1041 B.n281 B.n269 10.6151
R1042 B.n282 B.n281 10.6151
R1043 B.n283 B.n282 10.6151
R1044 B.n283 B.n267 10.6151
R1045 B.n290 B.n289 10.6151
R1046 B.n291 B.n290 10.6151
R1047 B.n291 B.n262 10.6151
R1048 B.n297 B.n262 10.6151
R1049 B.n298 B.n297 10.6151
R1050 B.n299 B.n298 10.6151
R1051 B.n299 B.n260 10.6151
R1052 B.n305 B.n260 10.6151
R1053 B.n308 B.n307 10.6151
R1054 B.n308 B.n256 10.6151
R1055 B.n314 B.n256 10.6151
R1056 B.n315 B.n314 10.6151
R1057 B.n316 B.n315 10.6151
R1058 B.n316 B.n254 10.6151
R1059 B.n322 B.n254 10.6151
R1060 B.n323 B.n322 10.6151
R1061 B.n324 B.n246 10.6151
R1062 B.n334 B.n246 10.6151
R1063 B.n335 B.n334 10.6151
R1064 B.n336 B.n335 10.6151
R1065 B.n336 B.n238 10.6151
R1066 B.n346 B.n238 10.6151
R1067 B.n347 B.n346 10.6151
R1068 B.n348 B.n347 10.6151
R1069 B.n348 B.n230 10.6151
R1070 B.n358 B.n230 10.6151
R1071 B.n359 B.n358 10.6151
R1072 B.n360 B.n359 10.6151
R1073 B.n360 B.n222 10.6151
R1074 B.n370 B.n222 10.6151
R1075 B.n371 B.n370 10.6151
R1076 B.n372 B.n371 10.6151
R1077 B.n372 B.n214 10.6151
R1078 B.n382 B.n214 10.6151
R1079 B.n383 B.n382 10.6151
R1080 B.n384 B.n383 10.6151
R1081 B.n384 B.n207 10.6151
R1082 B.n395 B.n207 10.6151
R1083 B.n396 B.n395 10.6151
R1084 B.n397 B.n396 10.6151
R1085 B.n397 B.n199 10.6151
R1086 B.n407 B.n199 10.6151
R1087 B.n408 B.n407 10.6151
R1088 B.n409 B.n408 10.6151
R1089 B.n409 B.n190 10.6151
R1090 B.n419 B.n190 10.6151
R1091 B.n420 B.n419 10.6151
R1092 B.n421 B.n420 10.6151
R1093 B.n421 B.n183 10.6151
R1094 B.n431 B.n183 10.6151
R1095 B.n432 B.n431 10.6151
R1096 B.n433 B.n432 10.6151
R1097 B.n433 B.n175 10.6151
R1098 B.n443 B.n175 10.6151
R1099 B.n444 B.n443 10.6151
R1100 B.n445 B.n444 10.6151
R1101 B.n445 B.n168 10.6151
R1102 B.n456 B.n168 10.6151
R1103 B.n457 B.n456 10.6151
R1104 B.n459 B.n457 10.6151
R1105 B.n459 B.n458 10.6151
R1106 B.n458 B.n160 10.6151
R1107 B.n470 B.n160 10.6151
R1108 B.n471 B.n470 10.6151
R1109 B.n472 B.n471 10.6151
R1110 B.n473 B.n472 10.6151
R1111 B.n474 B.n473 10.6151
R1112 B.n477 B.n474 10.6151
R1113 B.n478 B.n477 10.6151
R1114 B.n479 B.n478 10.6151
R1115 B.n480 B.n479 10.6151
R1116 B.n482 B.n480 10.6151
R1117 B.n483 B.n482 10.6151
R1118 B.n484 B.n483 10.6151
R1119 B.n485 B.n484 10.6151
R1120 B.n487 B.n485 10.6151
R1121 B.n488 B.n487 10.6151
R1122 B.n489 B.n488 10.6151
R1123 B.n490 B.n489 10.6151
R1124 B.n492 B.n490 10.6151
R1125 B.n493 B.n492 10.6151
R1126 B.n494 B.n493 10.6151
R1127 B.n495 B.n494 10.6151
R1128 B.n497 B.n495 10.6151
R1129 B.n498 B.n497 10.6151
R1130 B.n499 B.n498 10.6151
R1131 B.n500 B.n499 10.6151
R1132 B.n502 B.n500 10.6151
R1133 B.n503 B.n502 10.6151
R1134 B.n504 B.n503 10.6151
R1135 B.n505 B.n504 10.6151
R1136 B.n507 B.n505 10.6151
R1137 B.n508 B.n507 10.6151
R1138 B.n509 B.n508 10.6151
R1139 B.n510 B.n509 10.6151
R1140 B.n512 B.n510 10.6151
R1141 B.n513 B.n512 10.6151
R1142 B.n514 B.n513 10.6151
R1143 B.n515 B.n514 10.6151
R1144 B.n517 B.n515 10.6151
R1145 B.n518 B.n517 10.6151
R1146 B.n519 B.n518 10.6151
R1147 B.n520 B.n519 10.6151
R1148 B.n522 B.n520 10.6151
R1149 B.n523 B.n522 10.6151
R1150 B.n524 B.n523 10.6151
R1151 B.n525 B.n524 10.6151
R1152 B.n527 B.n525 10.6151
R1153 B.n528 B.n527 10.6151
R1154 B.n529 B.n528 10.6151
R1155 B.n530 B.n529 10.6151
R1156 B.n532 B.n530 10.6151
R1157 B.n533 B.n532 10.6151
R1158 B.n629 B.n1 10.6151
R1159 B.n629 B.n628 10.6151
R1160 B.n628 B.n627 10.6151
R1161 B.n627 B.n10 10.6151
R1162 B.n621 B.n10 10.6151
R1163 B.n621 B.n620 10.6151
R1164 B.n620 B.n619 10.6151
R1165 B.n619 B.n17 10.6151
R1166 B.n613 B.n17 10.6151
R1167 B.n613 B.n612 10.6151
R1168 B.n612 B.n611 10.6151
R1169 B.n611 B.n25 10.6151
R1170 B.n605 B.n25 10.6151
R1171 B.n605 B.n604 10.6151
R1172 B.n604 B.n603 10.6151
R1173 B.n603 B.n32 10.6151
R1174 B.n597 B.n32 10.6151
R1175 B.n597 B.n596 10.6151
R1176 B.n596 B.n595 10.6151
R1177 B.n595 B.n39 10.6151
R1178 B.n589 B.n39 10.6151
R1179 B.n589 B.n588 10.6151
R1180 B.n588 B.n587 10.6151
R1181 B.n587 B.n46 10.6151
R1182 B.n581 B.n46 10.6151
R1183 B.n581 B.n580 10.6151
R1184 B.n580 B.n579 10.6151
R1185 B.n579 B.n52 10.6151
R1186 B.n573 B.n52 10.6151
R1187 B.n573 B.n572 10.6151
R1188 B.n572 B.n571 10.6151
R1189 B.n571 B.n60 10.6151
R1190 B.n565 B.n60 10.6151
R1191 B.n565 B.n564 10.6151
R1192 B.n564 B.n563 10.6151
R1193 B.n563 B.n67 10.6151
R1194 B.n557 B.n67 10.6151
R1195 B.n557 B.n556 10.6151
R1196 B.n556 B.n555 10.6151
R1197 B.n555 B.n74 10.6151
R1198 B.n549 B.n74 10.6151
R1199 B.n549 B.n548 10.6151
R1200 B.n548 B.n547 10.6151
R1201 B.n547 B.n81 10.6151
R1202 B.n541 B.n81 10.6151
R1203 B.n541 B.n540 10.6151
R1204 B.n540 B.n539 10.6151
R1205 B.n110 B.n88 10.6151
R1206 B.n113 B.n110 10.6151
R1207 B.n114 B.n113 10.6151
R1208 B.n117 B.n114 10.6151
R1209 B.n118 B.n117 10.6151
R1210 B.n121 B.n118 10.6151
R1211 B.n122 B.n121 10.6151
R1212 B.n125 B.n122 10.6151
R1213 B.n130 B.n127 10.6151
R1214 B.n131 B.n130 10.6151
R1215 B.n134 B.n131 10.6151
R1216 B.n135 B.n134 10.6151
R1217 B.n138 B.n135 10.6151
R1218 B.n139 B.n138 10.6151
R1219 B.n142 B.n139 10.6151
R1220 B.n143 B.n142 10.6151
R1221 B.n147 B.n146 10.6151
R1222 B.n150 B.n147 10.6151
R1223 B.n151 B.n150 10.6151
R1224 B.n154 B.n151 10.6151
R1225 B.n155 B.n154 10.6151
R1226 B.n158 B.n155 10.6151
R1227 B.n159 B.n158 10.6151
R1228 B.n534 B.n159 10.6151
R1229 B.n637 B.n0 8.11757
R1230 B.n637 B.n1 8.11757
R1231 B.n289 B.n266 6.5566
R1232 B.n306 B.n305 6.5566
R1233 B.n127 B.n126 6.5566
R1234 B.n143 B.n107 6.5566
R1235 B.n267 B.n266 4.05904
R1236 B.n307 B.n306 4.05904
R1237 B.n126 B.n125 4.05904
R1238 B.n146 B.n107 4.05904
R1239 VN.n30 VN.n29 161.3
R1240 VN.n28 VN.n17 161.3
R1241 VN.n27 VN.n26 161.3
R1242 VN.n25 VN.n18 161.3
R1243 VN.n24 VN.n23 161.3
R1244 VN.n22 VN.n19 161.3
R1245 VN.n14 VN.n13 161.3
R1246 VN.n12 VN.n1 161.3
R1247 VN.n11 VN.n10 161.3
R1248 VN.n9 VN.n2 161.3
R1249 VN.n8 VN.n7 161.3
R1250 VN.n6 VN.n3 161.3
R1251 VN.n15 VN.n0 69.5884
R1252 VN.n31 VN.n16 69.5884
R1253 VN.n11 VN.n2 56.5617
R1254 VN.n27 VN.n18 56.5617
R1255 VN.n5 VN.n4 49.5351
R1256 VN.n21 VN.n20 49.5351
R1257 VN VN.n31 42.4754
R1258 VN.n20 VN.t1 40.1968
R1259 VN.n4 VN.t0 40.1968
R1260 VN.n6 VN.n5 24.5923
R1261 VN.n7 VN.n6 24.5923
R1262 VN.n7 VN.n2 24.5923
R1263 VN.n12 VN.n11 24.5923
R1264 VN.n13 VN.n12 24.5923
R1265 VN.n23 VN.n18 24.5923
R1266 VN.n23 VN.n22 24.5923
R1267 VN.n22 VN.n21 24.5923
R1268 VN.n29 VN.n28 24.5923
R1269 VN.n28 VN.n27 24.5923
R1270 VN.n13 VN.n0 20.6576
R1271 VN.n29 VN.n16 20.6576
R1272 VN.n5 VN.t2 6.70794
R1273 VN.n0 VN.t4 6.70794
R1274 VN.n21 VN.t3 6.70794
R1275 VN.n16 VN.t5 6.70794
R1276 VN.n4 VN.n3 3.87331
R1277 VN.n20 VN.n19 3.87331
R1278 VN.n31 VN.n30 0.354861
R1279 VN.n15 VN.n14 0.354861
R1280 VN VN.n15 0.267071
R1281 VN.n30 VN.n17 0.189894
R1282 VN.n26 VN.n17 0.189894
R1283 VN.n26 VN.n25 0.189894
R1284 VN.n25 VN.n24 0.189894
R1285 VN.n24 VN.n19 0.189894
R1286 VN.n8 VN.n3 0.189894
R1287 VN.n9 VN.n8 0.189894
R1288 VN.n10 VN.n9 0.189894
R1289 VN.n10 VN.n1 0.189894
R1290 VN.n14 VN.n1 0.189894
R1291 VDD2.n1 VDD2.t5 262.596
R1292 VDD2.n2 VDD2.t0 260.44
R1293 VDD2.n1 VDD2.n0 238.099
R1294 VDD2 VDD2.n3 238.096
R1295 VDD2.n2 VDD2.n1 34.0386
R1296 VDD2.n3 VDD2.t2 23.0238
R1297 VDD2.n3 VDD2.t4 23.0238
R1298 VDD2.n0 VDD2.t3 23.0238
R1299 VDD2.n0 VDD2.t1 23.0238
R1300 VDD2 VDD2.n2 2.2699
C0 VDD2 VN 0.868671f
C1 VDD1 VDD2 1.59767f
C2 VTAIL VN 2.07724f
C3 VDD1 VTAIL 4.06049f
C4 VP VN 5.34417f
C5 VDD2 VTAIL 4.11725f
C6 VDD1 VP 1.21452f
C7 VP VDD2 0.509517f
C8 VDD1 VN 0.159888f
C9 VP VTAIL 2.09136f
C10 VDD2 B 4.252586f
C11 VDD1 B 4.553049f
C12 VTAIL B 3.118198f
C13 VN B 13.47079f
C14 VP B 11.960118f
C15 VDD2.t5 B 0.081465f
C16 VDD2.t3 B 0.012967f
C17 VDD2.t1 B 0.012967f
C18 VDD2.n0 B 0.051335f
C19 VDD2.n1 B 1.76937f
C20 VDD2.t0 B 0.079261f
C21 VDD2.n2 B 1.4828f
C22 VDD2.t2 B 0.012967f
C23 VDD2.t4 B 0.012967f
C24 VDD2.n3 B 0.051329f
C25 VN.t4 B 0.144462f
C26 VN.n0 B 0.236507f
C27 VN.n1 B 0.031675f
C28 VN.n2 B 0.042539f
C29 VN.n3 B 0.360256f
C30 VN.t2 B 0.144462f
C31 VN.t0 B 0.420978f
C32 VN.n4 B 0.238326f
C33 VN.n5 B 0.225921f
C34 VN.n6 B 0.058738f
C35 VN.n7 B 0.058738f
C36 VN.n8 B 0.031675f
C37 VN.n9 B 0.031675f
C38 VN.n10 B 0.031675f
C39 VN.n11 B 0.04955f
C40 VN.n12 B 0.058738f
C41 VN.n13 B 0.054099f
C42 VN.n14 B 0.051115f
C43 VN.n15 B 0.06598f
C44 VN.t5 B 0.144462f
C45 VN.n16 B 0.236507f
C46 VN.n17 B 0.031675f
C47 VN.n18 B 0.042539f
C48 VN.n19 B 0.360256f
C49 VN.t3 B 0.144462f
C50 VN.t1 B 0.420978f
C51 VN.n20 B 0.238326f
C52 VN.n21 B 0.225921f
C53 VN.n22 B 0.058738f
C54 VN.n23 B 0.058738f
C55 VN.n24 B 0.031675f
C56 VN.n25 B 0.031675f
C57 VN.n26 B 0.031675f
C58 VN.n27 B 0.04955f
C59 VN.n28 B 0.058738f
C60 VN.n29 B 0.054099f
C61 VN.n30 B 0.051115f
C62 VN.n31 B 1.40687f
C63 VTAIL.t1 B 0.028468f
C64 VTAIL.t3 B 0.028468f
C65 VTAIL.n0 B 0.090912f
C66 VTAIL.n1 B 0.599365f
C67 VTAIL.t9 B 0.155322f
C68 VTAIL.n2 B 0.90321f
C69 VTAIL.t10 B 0.028468f
C70 VTAIL.t11 B 0.028468f
C71 VTAIL.n3 B 0.090912f
C72 VTAIL.n4 B 2.0926f
C73 VTAIL.t2 B 0.028468f
C74 VTAIL.t5 B 0.028468f
C75 VTAIL.n5 B 0.090912f
C76 VTAIL.n6 B 2.0926f
C77 VTAIL.t4 B 0.155322f
C78 VTAIL.n7 B 0.903209f
C79 VTAIL.t7 B 0.028468f
C80 VTAIL.t6 B 0.028468f
C81 VTAIL.n8 B 0.090912f
C82 VTAIL.n9 B 0.889978f
C83 VTAIL.t8 B 0.155322f
C84 VTAIL.n10 B 1.70787f
C85 VTAIL.t0 B 0.155322f
C86 VTAIL.n11 B 1.60053f
C87 VDD1.t0 B 0.080259f
C88 VDD1.t4 B 0.080088f
C89 VDD1.t5 B 0.012748f
C90 VDD1.t1 B 0.012748f
C91 VDD1.n0 B 0.050468f
C92 VDD1.n1 B 1.83224f
C93 VDD1.t2 B 0.012748f
C94 VDD1.t3 B 0.012748f
C95 VDD1.n2 B 0.049474f
C96 VDD1.n3 B 1.51001f
C97 VP.t2 B 0.145336f
C98 VP.n0 B 0.237939f
C99 VP.n1 B 0.031867f
C100 VP.n2 B 0.042797f
C101 VP.n3 B 0.031867f
C102 VP.t0 B 0.145336f
C103 VP.n4 B 0.059094f
C104 VP.n5 B 0.031867f
C105 VP.n6 B 0.059094f
C106 VP.t3 B 0.145336f
C107 VP.n7 B 0.237939f
C108 VP.n8 B 0.031867f
C109 VP.n9 B 0.042797f
C110 VP.n10 B 0.362437f
C111 VP.t5 B 0.145336f
C112 VP.t4 B 0.423526f
C113 VP.n11 B 0.239769f
C114 VP.n12 B 0.227289f
C115 VP.n13 B 0.059094f
C116 VP.n14 B 0.059094f
C117 VP.n15 B 0.031867f
C118 VP.n16 B 0.031867f
C119 VP.n17 B 0.031867f
C120 VP.n18 B 0.04985f
C121 VP.n19 B 0.059094f
C122 VP.n20 B 0.054426f
C123 VP.n21 B 0.051424f
C124 VP.n22 B 1.40155f
C125 VP.n23 B 1.4287f
C126 VP.t1 B 0.145336f
C127 VP.n24 B 0.237939f
C128 VP.n25 B 0.054426f
C129 VP.n26 B 0.051424f
C130 VP.n27 B 0.031867f
C131 VP.n28 B 0.031867f
C132 VP.n29 B 0.04985f
C133 VP.n30 B 0.042797f
C134 VP.n31 B 0.059094f
C135 VP.n32 B 0.031867f
C136 VP.n33 B 0.031867f
C137 VP.n34 B 0.031867f
C138 VP.n35 B 0.138201f
C139 VP.n36 B 0.059094f
C140 VP.n37 B 0.059094f
C141 VP.n38 B 0.031867f
C142 VP.n39 B 0.031867f
C143 VP.n40 B 0.031867f
C144 VP.n41 B 0.04985f
C145 VP.n42 B 0.059094f
C146 VP.n43 B 0.054426f
C147 VP.n44 B 0.051424f
C148 VP.n45 B 0.06638f
.ends

