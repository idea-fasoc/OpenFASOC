* NGSPICE file created from diff_pair_sample_1189.ext - technology: sky130A

.subckt diff_pair_sample_1189 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=0 ps=0 w=17.06 l=1.91
X1 VDD1.t5 VP.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=2.8149 ps=17.39 w=17.06 l=1.91
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=0 ps=0 w=17.06 l=1.91
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=0 ps=0 w=17.06 l=1.91
X4 VTAIL.t6 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=2.8149 ps=17.39 w=17.06 l=1.91
X5 VDD2.t5 VN.t0 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=2.8149 ps=17.39 w=17.06 l=1.91
X6 VDD2.t4 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=6.6534 ps=34.9 w=17.06 l=1.91
X7 VDD1.t3 VP.t2 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=2.8149 ps=17.39 w=17.06 l=1.91
X8 VDD2.t3 VN.t2 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=6.6534 ps=34.9 w=17.06 l=1.91
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=0 ps=0 w=17.06 l=1.91
X10 VDD1.t2 VP.t3 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=6.6534 ps=34.9 w=17.06 l=1.91
X11 VDD2.t2 VN.t3 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.6534 pd=34.9 as=2.8149 ps=17.39 w=17.06 l=1.91
X12 VTAIL.t3 VN.t4 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=2.8149 ps=17.39 w=17.06 l=1.91
X13 VTAIL.t4 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=2.8149 ps=17.39 w=17.06 l=1.91
X14 VDD1.t1 VP.t4 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=6.6534 ps=34.9 w=17.06 l=1.91
X15 VTAIL.t5 VP.t5 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8149 pd=17.39 as=2.8149 ps=17.39 w=17.06 l=1.91
R0 B.n659 B.n132 585
R1 B.n132 B.n65 585
R2 B.n661 B.n660 585
R3 B.n663 B.n131 585
R4 B.n666 B.n665 585
R5 B.n667 B.n130 585
R6 B.n669 B.n668 585
R7 B.n671 B.n129 585
R8 B.n674 B.n673 585
R9 B.n675 B.n128 585
R10 B.n677 B.n676 585
R11 B.n679 B.n127 585
R12 B.n682 B.n681 585
R13 B.n683 B.n126 585
R14 B.n685 B.n684 585
R15 B.n687 B.n125 585
R16 B.n690 B.n689 585
R17 B.n691 B.n124 585
R18 B.n693 B.n692 585
R19 B.n695 B.n123 585
R20 B.n698 B.n697 585
R21 B.n699 B.n122 585
R22 B.n701 B.n700 585
R23 B.n703 B.n121 585
R24 B.n706 B.n705 585
R25 B.n707 B.n120 585
R26 B.n709 B.n708 585
R27 B.n711 B.n119 585
R28 B.n714 B.n713 585
R29 B.n715 B.n118 585
R30 B.n717 B.n716 585
R31 B.n719 B.n117 585
R32 B.n722 B.n721 585
R33 B.n723 B.n116 585
R34 B.n725 B.n724 585
R35 B.n727 B.n115 585
R36 B.n730 B.n729 585
R37 B.n731 B.n114 585
R38 B.n733 B.n732 585
R39 B.n735 B.n113 585
R40 B.n738 B.n737 585
R41 B.n739 B.n112 585
R42 B.n741 B.n740 585
R43 B.n743 B.n111 585
R44 B.n746 B.n745 585
R45 B.n747 B.n110 585
R46 B.n749 B.n748 585
R47 B.n751 B.n109 585
R48 B.n754 B.n753 585
R49 B.n755 B.n108 585
R50 B.n757 B.n756 585
R51 B.n759 B.n107 585
R52 B.n762 B.n761 585
R53 B.n763 B.n106 585
R54 B.n765 B.n764 585
R55 B.n767 B.n105 585
R56 B.n769 B.n768 585
R57 B.n771 B.n770 585
R58 B.n774 B.n773 585
R59 B.n775 B.n100 585
R60 B.n777 B.n776 585
R61 B.n779 B.n99 585
R62 B.n782 B.n781 585
R63 B.n783 B.n98 585
R64 B.n785 B.n784 585
R65 B.n787 B.n97 585
R66 B.n790 B.n789 585
R67 B.n792 B.n94 585
R68 B.n794 B.n793 585
R69 B.n796 B.n93 585
R70 B.n799 B.n798 585
R71 B.n800 B.n92 585
R72 B.n802 B.n801 585
R73 B.n804 B.n91 585
R74 B.n807 B.n806 585
R75 B.n808 B.n90 585
R76 B.n810 B.n809 585
R77 B.n812 B.n89 585
R78 B.n815 B.n814 585
R79 B.n816 B.n88 585
R80 B.n818 B.n817 585
R81 B.n820 B.n87 585
R82 B.n823 B.n822 585
R83 B.n824 B.n86 585
R84 B.n826 B.n825 585
R85 B.n828 B.n85 585
R86 B.n831 B.n830 585
R87 B.n832 B.n84 585
R88 B.n834 B.n833 585
R89 B.n836 B.n83 585
R90 B.n839 B.n838 585
R91 B.n840 B.n82 585
R92 B.n842 B.n841 585
R93 B.n844 B.n81 585
R94 B.n847 B.n846 585
R95 B.n848 B.n80 585
R96 B.n850 B.n849 585
R97 B.n852 B.n79 585
R98 B.n855 B.n854 585
R99 B.n856 B.n78 585
R100 B.n858 B.n857 585
R101 B.n860 B.n77 585
R102 B.n863 B.n862 585
R103 B.n864 B.n76 585
R104 B.n866 B.n865 585
R105 B.n868 B.n75 585
R106 B.n871 B.n870 585
R107 B.n872 B.n74 585
R108 B.n874 B.n873 585
R109 B.n876 B.n73 585
R110 B.n879 B.n878 585
R111 B.n880 B.n72 585
R112 B.n882 B.n881 585
R113 B.n884 B.n71 585
R114 B.n887 B.n886 585
R115 B.n888 B.n70 585
R116 B.n890 B.n889 585
R117 B.n892 B.n69 585
R118 B.n895 B.n894 585
R119 B.n896 B.n68 585
R120 B.n898 B.n897 585
R121 B.n900 B.n67 585
R122 B.n903 B.n902 585
R123 B.n904 B.n66 585
R124 B.n658 B.n64 585
R125 B.n907 B.n64 585
R126 B.n657 B.n63 585
R127 B.n908 B.n63 585
R128 B.n656 B.n62 585
R129 B.n909 B.n62 585
R130 B.n655 B.n654 585
R131 B.n654 B.n58 585
R132 B.n653 B.n57 585
R133 B.n915 B.n57 585
R134 B.n652 B.n56 585
R135 B.n916 B.n56 585
R136 B.n651 B.n55 585
R137 B.n917 B.n55 585
R138 B.n650 B.n649 585
R139 B.n649 B.n51 585
R140 B.n648 B.n50 585
R141 B.n923 B.n50 585
R142 B.n647 B.n49 585
R143 B.n924 B.n49 585
R144 B.n646 B.n48 585
R145 B.n925 B.n48 585
R146 B.n645 B.n644 585
R147 B.n644 B.n44 585
R148 B.n643 B.n43 585
R149 B.n931 B.n43 585
R150 B.n642 B.n42 585
R151 B.n932 B.n42 585
R152 B.n641 B.n41 585
R153 B.n933 B.n41 585
R154 B.n640 B.n639 585
R155 B.n639 B.n37 585
R156 B.n638 B.n36 585
R157 B.n939 B.n36 585
R158 B.n637 B.n35 585
R159 B.n940 B.n35 585
R160 B.n636 B.n34 585
R161 B.n941 B.n34 585
R162 B.n635 B.n634 585
R163 B.n634 B.n30 585
R164 B.n633 B.n29 585
R165 B.n947 B.n29 585
R166 B.n632 B.n28 585
R167 B.n948 B.n28 585
R168 B.n631 B.n27 585
R169 B.n949 B.n27 585
R170 B.n630 B.n629 585
R171 B.n629 B.n26 585
R172 B.n628 B.n22 585
R173 B.n955 B.n22 585
R174 B.n627 B.n21 585
R175 B.n956 B.n21 585
R176 B.n626 B.n20 585
R177 B.n957 B.n20 585
R178 B.n625 B.n624 585
R179 B.n624 B.n16 585
R180 B.n623 B.n15 585
R181 B.n963 B.n15 585
R182 B.n622 B.n14 585
R183 B.n964 B.n14 585
R184 B.n621 B.n13 585
R185 B.n965 B.n13 585
R186 B.n620 B.n619 585
R187 B.n619 B.n12 585
R188 B.n618 B.n617 585
R189 B.n618 B.n8 585
R190 B.n616 B.n7 585
R191 B.n972 B.n7 585
R192 B.n615 B.n6 585
R193 B.n973 B.n6 585
R194 B.n614 B.n5 585
R195 B.n974 B.n5 585
R196 B.n613 B.n612 585
R197 B.n612 B.n4 585
R198 B.n611 B.n133 585
R199 B.n611 B.n610 585
R200 B.n601 B.n134 585
R201 B.n135 B.n134 585
R202 B.n603 B.n602 585
R203 B.n604 B.n603 585
R204 B.n600 B.n139 585
R205 B.n143 B.n139 585
R206 B.n599 B.n598 585
R207 B.n598 B.n597 585
R208 B.n141 B.n140 585
R209 B.n142 B.n141 585
R210 B.n590 B.n589 585
R211 B.n591 B.n590 585
R212 B.n588 B.n148 585
R213 B.n148 B.n147 585
R214 B.n587 B.n586 585
R215 B.n586 B.n585 585
R216 B.n150 B.n149 585
R217 B.n578 B.n150 585
R218 B.n577 B.n576 585
R219 B.n579 B.n577 585
R220 B.n575 B.n155 585
R221 B.n155 B.n154 585
R222 B.n574 B.n573 585
R223 B.n573 B.n572 585
R224 B.n157 B.n156 585
R225 B.n158 B.n157 585
R226 B.n565 B.n564 585
R227 B.n566 B.n565 585
R228 B.n563 B.n163 585
R229 B.n163 B.n162 585
R230 B.n562 B.n561 585
R231 B.n561 B.n560 585
R232 B.n165 B.n164 585
R233 B.n166 B.n165 585
R234 B.n553 B.n552 585
R235 B.n554 B.n553 585
R236 B.n551 B.n171 585
R237 B.n171 B.n170 585
R238 B.n550 B.n549 585
R239 B.n549 B.n548 585
R240 B.n173 B.n172 585
R241 B.n174 B.n173 585
R242 B.n541 B.n540 585
R243 B.n542 B.n541 585
R244 B.n539 B.n179 585
R245 B.n179 B.n178 585
R246 B.n538 B.n537 585
R247 B.n537 B.n536 585
R248 B.n181 B.n180 585
R249 B.n182 B.n181 585
R250 B.n529 B.n528 585
R251 B.n530 B.n529 585
R252 B.n527 B.n187 585
R253 B.n187 B.n186 585
R254 B.n526 B.n525 585
R255 B.n525 B.n524 585
R256 B.n189 B.n188 585
R257 B.n190 B.n189 585
R258 B.n517 B.n516 585
R259 B.n518 B.n517 585
R260 B.n515 B.n195 585
R261 B.n195 B.n194 585
R262 B.n514 B.n513 585
R263 B.n513 B.n512 585
R264 B.n509 B.n199 585
R265 B.n508 B.n507 585
R266 B.n505 B.n200 585
R267 B.n505 B.n198 585
R268 B.n504 B.n503 585
R269 B.n502 B.n501 585
R270 B.n500 B.n202 585
R271 B.n498 B.n497 585
R272 B.n496 B.n203 585
R273 B.n495 B.n494 585
R274 B.n492 B.n204 585
R275 B.n490 B.n489 585
R276 B.n488 B.n205 585
R277 B.n487 B.n486 585
R278 B.n484 B.n206 585
R279 B.n482 B.n481 585
R280 B.n480 B.n207 585
R281 B.n479 B.n478 585
R282 B.n476 B.n208 585
R283 B.n474 B.n473 585
R284 B.n472 B.n209 585
R285 B.n471 B.n470 585
R286 B.n468 B.n210 585
R287 B.n466 B.n465 585
R288 B.n464 B.n211 585
R289 B.n463 B.n462 585
R290 B.n460 B.n212 585
R291 B.n458 B.n457 585
R292 B.n456 B.n213 585
R293 B.n455 B.n454 585
R294 B.n452 B.n214 585
R295 B.n450 B.n449 585
R296 B.n448 B.n215 585
R297 B.n447 B.n446 585
R298 B.n444 B.n216 585
R299 B.n442 B.n441 585
R300 B.n440 B.n217 585
R301 B.n439 B.n438 585
R302 B.n436 B.n218 585
R303 B.n434 B.n433 585
R304 B.n432 B.n219 585
R305 B.n431 B.n430 585
R306 B.n428 B.n220 585
R307 B.n426 B.n425 585
R308 B.n424 B.n221 585
R309 B.n423 B.n422 585
R310 B.n420 B.n222 585
R311 B.n418 B.n417 585
R312 B.n416 B.n223 585
R313 B.n415 B.n414 585
R314 B.n412 B.n224 585
R315 B.n410 B.n409 585
R316 B.n408 B.n225 585
R317 B.n407 B.n406 585
R318 B.n404 B.n226 585
R319 B.n402 B.n401 585
R320 B.n400 B.n227 585
R321 B.n399 B.n398 585
R322 B.n396 B.n395 585
R323 B.n394 B.n393 585
R324 B.n392 B.n232 585
R325 B.n390 B.n389 585
R326 B.n388 B.n233 585
R327 B.n387 B.n386 585
R328 B.n384 B.n234 585
R329 B.n382 B.n381 585
R330 B.n380 B.n235 585
R331 B.n378 B.n377 585
R332 B.n375 B.n238 585
R333 B.n373 B.n372 585
R334 B.n371 B.n239 585
R335 B.n370 B.n369 585
R336 B.n367 B.n240 585
R337 B.n365 B.n364 585
R338 B.n363 B.n241 585
R339 B.n362 B.n361 585
R340 B.n359 B.n242 585
R341 B.n357 B.n356 585
R342 B.n355 B.n243 585
R343 B.n354 B.n353 585
R344 B.n351 B.n244 585
R345 B.n349 B.n348 585
R346 B.n347 B.n245 585
R347 B.n346 B.n345 585
R348 B.n343 B.n246 585
R349 B.n341 B.n340 585
R350 B.n339 B.n247 585
R351 B.n338 B.n337 585
R352 B.n335 B.n248 585
R353 B.n333 B.n332 585
R354 B.n331 B.n249 585
R355 B.n330 B.n329 585
R356 B.n327 B.n250 585
R357 B.n325 B.n324 585
R358 B.n323 B.n251 585
R359 B.n322 B.n321 585
R360 B.n319 B.n252 585
R361 B.n317 B.n316 585
R362 B.n315 B.n253 585
R363 B.n314 B.n313 585
R364 B.n311 B.n254 585
R365 B.n309 B.n308 585
R366 B.n307 B.n255 585
R367 B.n306 B.n305 585
R368 B.n303 B.n256 585
R369 B.n301 B.n300 585
R370 B.n299 B.n257 585
R371 B.n298 B.n297 585
R372 B.n295 B.n258 585
R373 B.n293 B.n292 585
R374 B.n291 B.n259 585
R375 B.n290 B.n289 585
R376 B.n287 B.n260 585
R377 B.n285 B.n284 585
R378 B.n283 B.n261 585
R379 B.n282 B.n281 585
R380 B.n279 B.n262 585
R381 B.n277 B.n276 585
R382 B.n275 B.n263 585
R383 B.n274 B.n273 585
R384 B.n271 B.n264 585
R385 B.n269 B.n268 585
R386 B.n267 B.n266 585
R387 B.n197 B.n196 585
R388 B.n511 B.n510 585
R389 B.n512 B.n511 585
R390 B.n193 B.n192 585
R391 B.n194 B.n193 585
R392 B.n520 B.n519 585
R393 B.n519 B.n518 585
R394 B.n521 B.n191 585
R395 B.n191 B.n190 585
R396 B.n523 B.n522 585
R397 B.n524 B.n523 585
R398 B.n185 B.n184 585
R399 B.n186 B.n185 585
R400 B.n532 B.n531 585
R401 B.n531 B.n530 585
R402 B.n533 B.n183 585
R403 B.n183 B.n182 585
R404 B.n535 B.n534 585
R405 B.n536 B.n535 585
R406 B.n177 B.n176 585
R407 B.n178 B.n177 585
R408 B.n544 B.n543 585
R409 B.n543 B.n542 585
R410 B.n545 B.n175 585
R411 B.n175 B.n174 585
R412 B.n547 B.n546 585
R413 B.n548 B.n547 585
R414 B.n169 B.n168 585
R415 B.n170 B.n169 585
R416 B.n556 B.n555 585
R417 B.n555 B.n554 585
R418 B.n557 B.n167 585
R419 B.n167 B.n166 585
R420 B.n559 B.n558 585
R421 B.n560 B.n559 585
R422 B.n161 B.n160 585
R423 B.n162 B.n161 585
R424 B.n568 B.n567 585
R425 B.n567 B.n566 585
R426 B.n569 B.n159 585
R427 B.n159 B.n158 585
R428 B.n571 B.n570 585
R429 B.n572 B.n571 585
R430 B.n153 B.n152 585
R431 B.n154 B.n153 585
R432 B.n581 B.n580 585
R433 B.n580 B.n579 585
R434 B.n582 B.n151 585
R435 B.n578 B.n151 585
R436 B.n584 B.n583 585
R437 B.n585 B.n584 585
R438 B.n146 B.n145 585
R439 B.n147 B.n146 585
R440 B.n593 B.n592 585
R441 B.n592 B.n591 585
R442 B.n594 B.n144 585
R443 B.n144 B.n142 585
R444 B.n596 B.n595 585
R445 B.n597 B.n596 585
R446 B.n138 B.n137 585
R447 B.n143 B.n138 585
R448 B.n606 B.n605 585
R449 B.n605 B.n604 585
R450 B.n607 B.n136 585
R451 B.n136 B.n135 585
R452 B.n609 B.n608 585
R453 B.n610 B.n609 585
R454 B.n3 B.n0 585
R455 B.n4 B.n3 585
R456 B.n971 B.n1 585
R457 B.n972 B.n971 585
R458 B.n970 B.n969 585
R459 B.n970 B.n8 585
R460 B.n968 B.n9 585
R461 B.n12 B.n9 585
R462 B.n967 B.n966 585
R463 B.n966 B.n965 585
R464 B.n11 B.n10 585
R465 B.n964 B.n11 585
R466 B.n962 B.n961 585
R467 B.n963 B.n962 585
R468 B.n960 B.n17 585
R469 B.n17 B.n16 585
R470 B.n959 B.n958 585
R471 B.n958 B.n957 585
R472 B.n19 B.n18 585
R473 B.n956 B.n19 585
R474 B.n954 B.n953 585
R475 B.n955 B.n954 585
R476 B.n952 B.n23 585
R477 B.n26 B.n23 585
R478 B.n951 B.n950 585
R479 B.n950 B.n949 585
R480 B.n25 B.n24 585
R481 B.n948 B.n25 585
R482 B.n946 B.n945 585
R483 B.n947 B.n946 585
R484 B.n944 B.n31 585
R485 B.n31 B.n30 585
R486 B.n943 B.n942 585
R487 B.n942 B.n941 585
R488 B.n33 B.n32 585
R489 B.n940 B.n33 585
R490 B.n938 B.n937 585
R491 B.n939 B.n938 585
R492 B.n936 B.n38 585
R493 B.n38 B.n37 585
R494 B.n935 B.n934 585
R495 B.n934 B.n933 585
R496 B.n40 B.n39 585
R497 B.n932 B.n40 585
R498 B.n930 B.n929 585
R499 B.n931 B.n930 585
R500 B.n928 B.n45 585
R501 B.n45 B.n44 585
R502 B.n927 B.n926 585
R503 B.n926 B.n925 585
R504 B.n47 B.n46 585
R505 B.n924 B.n47 585
R506 B.n922 B.n921 585
R507 B.n923 B.n922 585
R508 B.n920 B.n52 585
R509 B.n52 B.n51 585
R510 B.n919 B.n918 585
R511 B.n918 B.n917 585
R512 B.n54 B.n53 585
R513 B.n916 B.n54 585
R514 B.n914 B.n913 585
R515 B.n915 B.n914 585
R516 B.n912 B.n59 585
R517 B.n59 B.n58 585
R518 B.n911 B.n910 585
R519 B.n910 B.n909 585
R520 B.n61 B.n60 585
R521 B.n908 B.n61 585
R522 B.n906 B.n905 585
R523 B.n907 B.n906 585
R524 B.n975 B.n974 585
R525 B.n973 B.n2 585
R526 B.n906 B.n66 458.866
R527 B.n132 B.n64 458.866
R528 B.n513 B.n197 458.866
R529 B.n511 B.n199 458.866
R530 B.n95 B.t17 421.959
R531 B.n101 B.t13 421.959
R532 B.n236 B.t6 421.959
R533 B.n228 B.t10 421.959
R534 B.n662 B.n65 256.663
R535 B.n664 B.n65 256.663
R536 B.n670 B.n65 256.663
R537 B.n672 B.n65 256.663
R538 B.n678 B.n65 256.663
R539 B.n680 B.n65 256.663
R540 B.n686 B.n65 256.663
R541 B.n688 B.n65 256.663
R542 B.n694 B.n65 256.663
R543 B.n696 B.n65 256.663
R544 B.n702 B.n65 256.663
R545 B.n704 B.n65 256.663
R546 B.n710 B.n65 256.663
R547 B.n712 B.n65 256.663
R548 B.n718 B.n65 256.663
R549 B.n720 B.n65 256.663
R550 B.n726 B.n65 256.663
R551 B.n728 B.n65 256.663
R552 B.n734 B.n65 256.663
R553 B.n736 B.n65 256.663
R554 B.n742 B.n65 256.663
R555 B.n744 B.n65 256.663
R556 B.n750 B.n65 256.663
R557 B.n752 B.n65 256.663
R558 B.n758 B.n65 256.663
R559 B.n760 B.n65 256.663
R560 B.n766 B.n65 256.663
R561 B.n104 B.n65 256.663
R562 B.n772 B.n65 256.663
R563 B.n778 B.n65 256.663
R564 B.n780 B.n65 256.663
R565 B.n786 B.n65 256.663
R566 B.n788 B.n65 256.663
R567 B.n795 B.n65 256.663
R568 B.n797 B.n65 256.663
R569 B.n803 B.n65 256.663
R570 B.n805 B.n65 256.663
R571 B.n811 B.n65 256.663
R572 B.n813 B.n65 256.663
R573 B.n819 B.n65 256.663
R574 B.n821 B.n65 256.663
R575 B.n827 B.n65 256.663
R576 B.n829 B.n65 256.663
R577 B.n835 B.n65 256.663
R578 B.n837 B.n65 256.663
R579 B.n843 B.n65 256.663
R580 B.n845 B.n65 256.663
R581 B.n851 B.n65 256.663
R582 B.n853 B.n65 256.663
R583 B.n859 B.n65 256.663
R584 B.n861 B.n65 256.663
R585 B.n867 B.n65 256.663
R586 B.n869 B.n65 256.663
R587 B.n875 B.n65 256.663
R588 B.n877 B.n65 256.663
R589 B.n883 B.n65 256.663
R590 B.n885 B.n65 256.663
R591 B.n891 B.n65 256.663
R592 B.n893 B.n65 256.663
R593 B.n899 B.n65 256.663
R594 B.n901 B.n65 256.663
R595 B.n506 B.n198 256.663
R596 B.n201 B.n198 256.663
R597 B.n499 B.n198 256.663
R598 B.n493 B.n198 256.663
R599 B.n491 B.n198 256.663
R600 B.n485 B.n198 256.663
R601 B.n483 B.n198 256.663
R602 B.n477 B.n198 256.663
R603 B.n475 B.n198 256.663
R604 B.n469 B.n198 256.663
R605 B.n467 B.n198 256.663
R606 B.n461 B.n198 256.663
R607 B.n459 B.n198 256.663
R608 B.n453 B.n198 256.663
R609 B.n451 B.n198 256.663
R610 B.n445 B.n198 256.663
R611 B.n443 B.n198 256.663
R612 B.n437 B.n198 256.663
R613 B.n435 B.n198 256.663
R614 B.n429 B.n198 256.663
R615 B.n427 B.n198 256.663
R616 B.n421 B.n198 256.663
R617 B.n419 B.n198 256.663
R618 B.n413 B.n198 256.663
R619 B.n411 B.n198 256.663
R620 B.n405 B.n198 256.663
R621 B.n403 B.n198 256.663
R622 B.n397 B.n198 256.663
R623 B.n231 B.n198 256.663
R624 B.n391 B.n198 256.663
R625 B.n385 B.n198 256.663
R626 B.n383 B.n198 256.663
R627 B.n376 B.n198 256.663
R628 B.n374 B.n198 256.663
R629 B.n368 B.n198 256.663
R630 B.n366 B.n198 256.663
R631 B.n360 B.n198 256.663
R632 B.n358 B.n198 256.663
R633 B.n352 B.n198 256.663
R634 B.n350 B.n198 256.663
R635 B.n344 B.n198 256.663
R636 B.n342 B.n198 256.663
R637 B.n336 B.n198 256.663
R638 B.n334 B.n198 256.663
R639 B.n328 B.n198 256.663
R640 B.n326 B.n198 256.663
R641 B.n320 B.n198 256.663
R642 B.n318 B.n198 256.663
R643 B.n312 B.n198 256.663
R644 B.n310 B.n198 256.663
R645 B.n304 B.n198 256.663
R646 B.n302 B.n198 256.663
R647 B.n296 B.n198 256.663
R648 B.n294 B.n198 256.663
R649 B.n288 B.n198 256.663
R650 B.n286 B.n198 256.663
R651 B.n280 B.n198 256.663
R652 B.n278 B.n198 256.663
R653 B.n272 B.n198 256.663
R654 B.n270 B.n198 256.663
R655 B.n265 B.n198 256.663
R656 B.n977 B.n976 256.663
R657 B.n902 B.n900 163.367
R658 B.n898 B.n68 163.367
R659 B.n894 B.n892 163.367
R660 B.n890 B.n70 163.367
R661 B.n886 B.n884 163.367
R662 B.n882 B.n72 163.367
R663 B.n878 B.n876 163.367
R664 B.n874 B.n74 163.367
R665 B.n870 B.n868 163.367
R666 B.n866 B.n76 163.367
R667 B.n862 B.n860 163.367
R668 B.n858 B.n78 163.367
R669 B.n854 B.n852 163.367
R670 B.n850 B.n80 163.367
R671 B.n846 B.n844 163.367
R672 B.n842 B.n82 163.367
R673 B.n838 B.n836 163.367
R674 B.n834 B.n84 163.367
R675 B.n830 B.n828 163.367
R676 B.n826 B.n86 163.367
R677 B.n822 B.n820 163.367
R678 B.n818 B.n88 163.367
R679 B.n814 B.n812 163.367
R680 B.n810 B.n90 163.367
R681 B.n806 B.n804 163.367
R682 B.n802 B.n92 163.367
R683 B.n798 B.n796 163.367
R684 B.n794 B.n94 163.367
R685 B.n789 B.n787 163.367
R686 B.n785 B.n98 163.367
R687 B.n781 B.n779 163.367
R688 B.n777 B.n100 163.367
R689 B.n773 B.n771 163.367
R690 B.n768 B.n767 163.367
R691 B.n765 B.n106 163.367
R692 B.n761 B.n759 163.367
R693 B.n757 B.n108 163.367
R694 B.n753 B.n751 163.367
R695 B.n749 B.n110 163.367
R696 B.n745 B.n743 163.367
R697 B.n741 B.n112 163.367
R698 B.n737 B.n735 163.367
R699 B.n733 B.n114 163.367
R700 B.n729 B.n727 163.367
R701 B.n725 B.n116 163.367
R702 B.n721 B.n719 163.367
R703 B.n717 B.n118 163.367
R704 B.n713 B.n711 163.367
R705 B.n709 B.n120 163.367
R706 B.n705 B.n703 163.367
R707 B.n701 B.n122 163.367
R708 B.n697 B.n695 163.367
R709 B.n693 B.n124 163.367
R710 B.n689 B.n687 163.367
R711 B.n685 B.n126 163.367
R712 B.n681 B.n679 163.367
R713 B.n677 B.n128 163.367
R714 B.n673 B.n671 163.367
R715 B.n669 B.n130 163.367
R716 B.n665 B.n663 163.367
R717 B.n661 B.n132 163.367
R718 B.n513 B.n195 163.367
R719 B.n517 B.n195 163.367
R720 B.n517 B.n189 163.367
R721 B.n525 B.n189 163.367
R722 B.n525 B.n187 163.367
R723 B.n529 B.n187 163.367
R724 B.n529 B.n181 163.367
R725 B.n537 B.n181 163.367
R726 B.n537 B.n179 163.367
R727 B.n541 B.n179 163.367
R728 B.n541 B.n173 163.367
R729 B.n549 B.n173 163.367
R730 B.n549 B.n171 163.367
R731 B.n553 B.n171 163.367
R732 B.n553 B.n165 163.367
R733 B.n561 B.n165 163.367
R734 B.n561 B.n163 163.367
R735 B.n565 B.n163 163.367
R736 B.n565 B.n157 163.367
R737 B.n573 B.n157 163.367
R738 B.n573 B.n155 163.367
R739 B.n577 B.n155 163.367
R740 B.n577 B.n150 163.367
R741 B.n586 B.n150 163.367
R742 B.n586 B.n148 163.367
R743 B.n590 B.n148 163.367
R744 B.n590 B.n141 163.367
R745 B.n598 B.n141 163.367
R746 B.n598 B.n139 163.367
R747 B.n603 B.n139 163.367
R748 B.n603 B.n134 163.367
R749 B.n611 B.n134 163.367
R750 B.n612 B.n611 163.367
R751 B.n612 B.n5 163.367
R752 B.n6 B.n5 163.367
R753 B.n7 B.n6 163.367
R754 B.n618 B.n7 163.367
R755 B.n619 B.n618 163.367
R756 B.n619 B.n13 163.367
R757 B.n14 B.n13 163.367
R758 B.n15 B.n14 163.367
R759 B.n624 B.n15 163.367
R760 B.n624 B.n20 163.367
R761 B.n21 B.n20 163.367
R762 B.n22 B.n21 163.367
R763 B.n629 B.n22 163.367
R764 B.n629 B.n27 163.367
R765 B.n28 B.n27 163.367
R766 B.n29 B.n28 163.367
R767 B.n634 B.n29 163.367
R768 B.n634 B.n34 163.367
R769 B.n35 B.n34 163.367
R770 B.n36 B.n35 163.367
R771 B.n639 B.n36 163.367
R772 B.n639 B.n41 163.367
R773 B.n42 B.n41 163.367
R774 B.n43 B.n42 163.367
R775 B.n644 B.n43 163.367
R776 B.n644 B.n48 163.367
R777 B.n49 B.n48 163.367
R778 B.n50 B.n49 163.367
R779 B.n649 B.n50 163.367
R780 B.n649 B.n55 163.367
R781 B.n56 B.n55 163.367
R782 B.n57 B.n56 163.367
R783 B.n654 B.n57 163.367
R784 B.n654 B.n62 163.367
R785 B.n63 B.n62 163.367
R786 B.n64 B.n63 163.367
R787 B.n507 B.n505 163.367
R788 B.n505 B.n504 163.367
R789 B.n501 B.n500 163.367
R790 B.n498 B.n203 163.367
R791 B.n494 B.n492 163.367
R792 B.n490 B.n205 163.367
R793 B.n486 B.n484 163.367
R794 B.n482 B.n207 163.367
R795 B.n478 B.n476 163.367
R796 B.n474 B.n209 163.367
R797 B.n470 B.n468 163.367
R798 B.n466 B.n211 163.367
R799 B.n462 B.n460 163.367
R800 B.n458 B.n213 163.367
R801 B.n454 B.n452 163.367
R802 B.n450 B.n215 163.367
R803 B.n446 B.n444 163.367
R804 B.n442 B.n217 163.367
R805 B.n438 B.n436 163.367
R806 B.n434 B.n219 163.367
R807 B.n430 B.n428 163.367
R808 B.n426 B.n221 163.367
R809 B.n422 B.n420 163.367
R810 B.n418 B.n223 163.367
R811 B.n414 B.n412 163.367
R812 B.n410 B.n225 163.367
R813 B.n406 B.n404 163.367
R814 B.n402 B.n227 163.367
R815 B.n398 B.n396 163.367
R816 B.n393 B.n392 163.367
R817 B.n390 B.n233 163.367
R818 B.n386 B.n384 163.367
R819 B.n382 B.n235 163.367
R820 B.n377 B.n375 163.367
R821 B.n373 B.n239 163.367
R822 B.n369 B.n367 163.367
R823 B.n365 B.n241 163.367
R824 B.n361 B.n359 163.367
R825 B.n357 B.n243 163.367
R826 B.n353 B.n351 163.367
R827 B.n349 B.n245 163.367
R828 B.n345 B.n343 163.367
R829 B.n341 B.n247 163.367
R830 B.n337 B.n335 163.367
R831 B.n333 B.n249 163.367
R832 B.n329 B.n327 163.367
R833 B.n325 B.n251 163.367
R834 B.n321 B.n319 163.367
R835 B.n317 B.n253 163.367
R836 B.n313 B.n311 163.367
R837 B.n309 B.n255 163.367
R838 B.n305 B.n303 163.367
R839 B.n301 B.n257 163.367
R840 B.n297 B.n295 163.367
R841 B.n293 B.n259 163.367
R842 B.n289 B.n287 163.367
R843 B.n285 B.n261 163.367
R844 B.n281 B.n279 163.367
R845 B.n277 B.n263 163.367
R846 B.n273 B.n271 163.367
R847 B.n269 B.n266 163.367
R848 B.n511 B.n193 163.367
R849 B.n519 B.n193 163.367
R850 B.n519 B.n191 163.367
R851 B.n523 B.n191 163.367
R852 B.n523 B.n185 163.367
R853 B.n531 B.n185 163.367
R854 B.n531 B.n183 163.367
R855 B.n535 B.n183 163.367
R856 B.n535 B.n177 163.367
R857 B.n543 B.n177 163.367
R858 B.n543 B.n175 163.367
R859 B.n547 B.n175 163.367
R860 B.n547 B.n169 163.367
R861 B.n555 B.n169 163.367
R862 B.n555 B.n167 163.367
R863 B.n559 B.n167 163.367
R864 B.n559 B.n161 163.367
R865 B.n567 B.n161 163.367
R866 B.n567 B.n159 163.367
R867 B.n571 B.n159 163.367
R868 B.n571 B.n153 163.367
R869 B.n580 B.n153 163.367
R870 B.n580 B.n151 163.367
R871 B.n584 B.n151 163.367
R872 B.n584 B.n146 163.367
R873 B.n592 B.n146 163.367
R874 B.n592 B.n144 163.367
R875 B.n596 B.n144 163.367
R876 B.n596 B.n138 163.367
R877 B.n605 B.n138 163.367
R878 B.n605 B.n136 163.367
R879 B.n609 B.n136 163.367
R880 B.n609 B.n3 163.367
R881 B.n975 B.n3 163.367
R882 B.n971 B.n2 163.367
R883 B.n971 B.n970 163.367
R884 B.n970 B.n9 163.367
R885 B.n966 B.n9 163.367
R886 B.n966 B.n11 163.367
R887 B.n962 B.n11 163.367
R888 B.n962 B.n17 163.367
R889 B.n958 B.n17 163.367
R890 B.n958 B.n19 163.367
R891 B.n954 B.n19 163.367
R892 B.n954 B.n23 163.367
R893 B.n950 B.n23 163.367
R894 B.n950 B.n25 163.367
R895 B.n946 B.n25 163.367
R896 B.n946 B.n31 163.367
R897 B.n942 B.n31 163.367
R898 B.n942 B.n33 163.367
R899 B.n938 B.n33 163.367
R900 B.n938 B.n38 163.367
R901 B.n934 B.n38 163.367
R902 B.n934 B.n40 163.367
R903 B.n930 B.n40 163.367
R904 B.n930 B.n45 163.367
R905 B.n926 B.n45 163.367
R906 B.n926 B.n47 163.367
R907 B.n922 B.n47 163.367
R908 B.n922 B.n52 163.367
R909 B.n918 B.n52 163.367
R910 B.n918 B.n54 163.367
R911 B.n914 B.n54 163.367
R912 B.n914 B.n59 163.367
R913 B.n910 B.n59 163.367
R914 B.n910 B.n61 163.367
R915 B.n906 B.n61 163.367
R916 B.n101 B.t15 111.915
R917 B.n236 B.t9 111.915
R918 B.n95 B.t18 111.891
R919 B.n228 B.t12 111.891
R920 B.n901 B.n66 71.676
R921 B.n900 B.n899 71.676
R922 B.n893 B.n68 71.676
R923 B.n892 B.n891 71.676
R924 B.n885 B.n70 71.676
R925 B.n884 B.n883 71.676
R926 B.n877 B.n72 71.676
R927 B.n876 B.n875 71.676
R928 B.n869 B.n74 71.676
R929 B.n868 B.n867 71.676
R930 B.n861 B.n76 71.676
R931 B.n860 B.n859 71.676
R932 B.n853 B.n78 71.676
R933 B.n852 B.n851 71.676
R934 B.n845 B.n80 71.676
R935 B.n844 B.n843 71.676
R936 B.n837 B.n82 71.676
R937 B.n836 B.n835 71.676
R938 B.n829 B.n84 71.676
R939 B.n828 B.n827 71.676
R940 B.n821 B.n86 71.676
R941 B.n820 B.n819 71.676
R942 B.n813 B.n88 71.676
R943 B.n812 B.n811 71.676
R944 B.n805 B.n90 71.676
R945 B.n804 B.n803 71.676
R946 B.n797 B.n92 71.676
R947 B.n796 B.n795 71.676
R948 B.n788 B.n94 71.676
R949 B.n787 B.n786 71.676
R950 B.n780 B.n98 71.676
R951 B.n779 B.n778 71.676
R952 B.n772 B.n100 71.676
R953 B.n771 B.n104 71.676
R954 B.n767 B.n766 71.676
R955 B.n760 B.n106 71.676
R956 B.n759 B.n758 71.676
R957 B.n752 B.n108 71.676
R958 B.n751 B.n750 71.676
R959 B.n744 B.n110 71.676
R960 B.n743 B.n742 71.676
R961 B.n736 B.n112 71.676
R962 B.n735 B.n734 71.676
R963 B.n728 B.n114 71.676
R964 B.n727 B.n726 71.676
R965 B.n720 B.n116 71.676
R966 B.n719 B.n718 71.676
R967 B.n712 B.n118 71.676
R968 B.n711 B.n710 71.676
R969 B.n704 B.n120 71.676
R970 B.n703 B.n702 71.676
R971 B.n696 B.n122 71.676
R972 B.n695 B.n694 71.676
R973 B.n688 B.n124 71.676
R974 B.n687 B.n686 71.676
R975 B.n680 B.n126 71.676
R976 B.n679 B.n678 71.676
R977 B.n672 B.n128 71.676
R978 B.n671 B.n670 71.676
R979 B.n664 B.n130 71.676
R980 B.n663 B.n662 71.676
R981 B.n662 B.n661 71.676
R982 B.n665 B.n664 71.676
R983 B.n670 B.n669 71.676
R984 B.n673 B.n672 71.676
R985 B.n678 B.n677 71.676
R986 B.n681 B.n680 71.676
R987 B.n686 B.n685 71.676
R988 B.n689 B.n688 71.676
R989 B.n694 B.n693 71.676
R990 B.n697 B.n696 71.676
R991 B.n702 B.n701 71.676
R992 B.n705 B.n704 71.676
R993 B.n710 B.n709 71.676
R994 B.n713 B.n712 71.676
R995 B.n718 B.n717 71.676
R996 B.n721 B.n720 71.676
R997 B.n726 B.n725 71.676
R998 B.n729 B.n728 71.676
R999 B.n734 B.n733 71.676
R1000 B.n737 B.n736 71.676
R1001 B.n742 B.n741 71.676
R1002 B.n745 B.n744 71.676
R1003 B.n750 B.n749 71.676
R1004 B.n753 B.n752 71.676
R1005 B.n758 B.n757 71.676
R1006 B.n761 B.n760 71.676
R1007 B.n766 B.n765 71.676
R1008 B.n768 B.n104 71.676
R1009 B.n773 B.n772 71.676
R1010 B.n778 B.n777 71.676
R1011 B.n781 B.n780 71.676
R1012 B.n786 B.n785 71.676
R1013 B.n789 B.n788 71.676
R1014 B.n795 B.n794 71.676
R1015 B.n798 B.n797 71.676
R1016 B.n803 B.n802 71.676
R1017 B.n806 B.n805 71.676
R1018 B.n811 B.n810 71.676
R1019 B.n814 B.n813 71.676
R1020 B.n819 B.n818 71.676
R1021 B.n822 B.n821 71.676
R1022 B.n827 B.n826 71.676
R1023 B.n830 B.n829 71.676
R1024 B.n835 B.n834 71.676
R1025 B.n838 B.n837 71.676
R1026 B.n843 B.n842 71.676
R1027 B.n846 B.n845 71.676
R1028 B.n851 B.n850 71.676
R1029 B.n854 B.n853 71.676
R1030 B.n859 B.n858 71.676
R1031 B.n862 B.n861 71.676
R1032 B.n867 B.n866 71.676
R1033 B.n870 B.n869 71.676
R1034 B.n875 B.n874 71.676
R1035 B.n878 B.n877 71.676
R1036 B.n883 B.n882 71.676
R1037 B.n886 B.n885 71.676
R1038 B.n891 B.n890 71.676
R1039 B.n894 B.n893 71.676
R1040 B.n899 B.n898 71.676
R1041 B.n902 B.n901 71.676
R1042 B.n506 B.n199 71.676
R1043 B.n504 B.n201 71.676
R1044 B.n500 B.n499 71.676
R1045 B.n493 B.n203 71.676
R1046 B.n492 B.n491 71.676
R1047 B.n485 B.n205 71.676
R1048 B.n484 B.n483 71.676
R1049 B.n477 B.n207 71.676
R1050 B.n476 B.n475 71.676
R1051 B.n469 B.n209 71.676
R1052 B.n468 B.n467 71.676
R1053 B.n461 B.n211 71.676
R1054 B.n460 B.n459 71.676
R1055 B.n453 B.n213 71.676
R1056 B.n452 B.n451 71.676
R1057 B.n445 B.n215 71.676
R1058 B.n444 B.n443 71.676
R1059 B.n437 B.n217 71.676
R1060 B.n436 B.n435 71.676
R1061 B.n429 B.n219 71.676
R1062 B.n428 B.n427 71.676
R1063 B.n421 B.n221 71.676
R1064 B.n420 B.n419 71.676
R1065 B.n413 B.n223 71.676
R1066 B.n412 B.n411 71.676
R1067 B.n405 B.n225 71.676
R1068 B.n404 B.n403 71.676
R1069 B.n397 B.n227 71.676
R1070 B.n396 B.n231 71.676
R1071 B.n392 B.n391 71.676
R1072 B.n385 B.n233 71.676
R1073 B.n384 B.n383 71.676
R1074 B.n376 B.n235 71.676
R1075 B.n375 B.n374 71.676
R1076 B.n368 B.n239 71.676
R1077 B.n367 B.n366 71.676
R1078 B.n360 B.n241 71.676
R1079 B.n359 B.n358 71.676
R1080 B.n352 B.n243 71.676
R1081 B.n351 B.n350 71.676
R1082 B.n344 B.n245 71.676
R1083 B.n343 B.n342 71.676
R1084 B.n336 B.n247 71.676
R1085 B.n335 B.n334 71.676
R1086 B.n328 B.n249 71.676
R1087 B.n327 B.n326 71.676
R1088 B.n320 B.n251 71.676
R1089 B.n319 B.n318 71.676
R1090 B.n312 B.n253 71.676
R1091 B.n311 B.n310 71.676
R1092 B.n304 B.n255 71.676
R1093 B.n303 B.n302 71.676
R1094 B.n296 B.n257 71.676
R1095 B.n295 B.n294 71.676
R1096 B.n288 B.n259 71.676
R1097 B.n287 B.n286 71.676
R1098 B.n280 B.n261 71.676
R1099 B.n279 B.n278 71.676
R1100 B.n272 B.n263 71.676
R1101 B.n271 B.n270 71.676
R1102 B.n266 B.n265 71.676
R1103 B.n507 B.n506 71.676
R1104 B.n501 B.n201 71.676
R1105 B.n499 B.n498 71.676
R1106 B.n494 B.n493 71.676
R1107 B.n491 B.n490 71.676
R1108 B.n486 B.n485 71.676
R1109 B.n483 B.n482 71.676
R1110 B.n478 B.n477 71.676
R1111 B.n475 B.n474 71.676
R1112 B.n470 B.n469 71.676
R1113 B.n467 B.n466 71.676
R1114 B.n462 B.n461 71.676
R1115 B.n459 B.n458 71.676
R1116 B.n454 B.n453 71.676
R1117 B.n451 B.n450 71.676
R1118 B.n446 B.n445 71.676
R1119 B.n443 B.n442 71.676
R1120 B.n438 B.n437 71.676
R1121 B.n435 B.n434 71.676
R1122 B.n430 B.n429 71.676
R1123 B.n427 B.n426 71.676
R1124 B.n422 B.n421 71.676
R1125 B.n419 B.n418 71.676
R1126 B.n414 B.n413 71.676
R1127 B.n411 B.n410 71.676
R1128 B.n406 B.n405 71.676
R1129 B.n403 B.n402 71.676
R1130 B.n398 B.n397 71.676
R1131 B.n393 B.n231 71.676
R1132 B.n391 B.n390 71.676
R1133 B.n386 B.n385 71.676
R1134 B.n383 B.n382 71.676
R1135 B.n377 B.n376 71.676
R1136 B.n374 B.n373 71.676
R1137 B.n369 B.n368 71.676
R1138 B.n366 B.n365 71.676
R1139 B.n361 B.n360 71.676
R1140 B.n358 B.n357 71.676
R1141 B.n353 B.n352 71.676
R1142 B.n350 B.n349 71.676
R1143 B.n345 B.n344 71.676
R1144 B.n342 B.n341 71.676
R1145 B.n337 B.n336 71.676
R1146 B.n334 B.n333 71.676
R1147 B.n329 B.n328 71.676
R1148 B.n326 B.n325 71.676
R1149 B.n321 B.n320 71.676
R1150 B.n318 B.n317 71.676
R1151 B.n313 B.n312 71.676
R1152 B.n310 B.n309 71.676
R1153 B.n305 B.n304 71.676
R1154 B.n302 B.n301 71.676
R1155 B.n297 B.n296 71.676
R1156 B.n294 B.n293 71.676
R1157 B.n289 B.n288 71.676
R1158 B.n286 B.n285 71.676
R1159 B.n281 B.n280 71.676
R1160 B.n278 B.n277 71.676
R1161 B.n273 B.n272 71.676
R1162 B.n270 B.n269 71.676
R1163 B.n265 B.n197 71.676
R1164 B.n976 B.n975 71.676
R1165 B.n976 B.n2 71.676
R1166 B.n102 B.t16 68.4716
R1167 B.n237 B.t8 68.4716
R1168 B.n96 B.t19 68.4489
R1169 B.n229 B.t11 68.4489
R1170 B.n512 B.n198 59.5931
R1171 B.n907 B.n65 59.5931
R1172 B.n791 B.n96 59.5399
R1173 B.n103 B.n102 59.5399
R1174 B.n379 B.n237 59.5399
R1175 B.n230 B.n229 59.5399
R1176 B.n96 B.n95 43.4429
R1177 B.n102 B.n101 43.4429
R1178 B.n237 B.n236 43.4429
R1179 B.n229 B.n228 43.4429
R1180 B.n512 B.n194 33.4905
R1181 B.n518 B.n194 33.4905
R1182 B.n518 B.n190 33.4905
R1183 B.n524 B.n190 33.4905
R1184 B.n524 B.n186 33.4905
R1185 B.n530 B.n186 33.4905
R1186 B.n536 B.n182 33.4905
R1187 B.n536 B.n178 33.4905
R1188 B.n542 B.n178 33.4905
R1189 B.n542 B.n174 33.4905
R1190 B.n548 B.n174 33.4905
R1191 B.n548 B.n170 33.4905
R1192 B.n554 B.n170 33.4905
R1193 B.n554 B.n166 33.4905
R1194 B.n560 B.n166 33.4905
R1195 B.n566 B.n162 33.4905
R1196 B.n566 B.n158 33.4905
R1197 B.n572 B.n158 33.4905
R1198 B.n572 B.n154 33.4905
R1199 B.n579 B.n154 33.4905
R1200 B.n579 B.n578 33.4905
R1201 B.n585 B.n147 33.4905
R1202 B.n591 B.n147 33.4905
R1203 B.n591 B.n142 33.4905
R1204 B.n597 B.n142 33.4905
R1205 B.n597 B.n143 33.4905
R1206 B.n604 B.n135 33.4905
R1207 B.n610 B.n135 33.4905
R1208 B.n610 B.n4 33.4905
R1209 B.n974 B.n4 33.4905
R1210 B.n974 B.n973 33.4905
R1211 B.n973 B.n972 33.4905
R1212 B.n972 B.n8 33.4905
R1213 B.n12 B.n8 33.4905
R1214 B.n965 B.n12 33.4905
R1215 B.n964 B.n963 33.4905
R1216 B.n963 B.n16 33.4905
R1217 B.n957 B.n16 33.4905
R1218 B.n957 B.n956 33.4905
R1219 B.n956 B.n955 33.4905
R1220 B.n949 B.n26 33.4905
R1221 B.n949 B.n948 33.4905
R1222 B.n948 B.n947 33.4905
R1223 B.n947 B.n30 33.4905
R1224 B.n941 B.n30 33.4905
R1225 B.n941 B.n940 33.4905
R1226 B.n939 B.n37 33.4905
R1227 B.n933 B.n37 33.4905
R1228 B.n933 B.n932 33.4905
R1229 B.n932 B.n931 33.4905
R1230 B.n931 B.n44 33.4905
R1231 B.n925 B.n44 33.4905
R1232 B.n925 B.n924 33.4905
R1233 B.n924 B.n923 33.4905
R1234 B.n923 B.n51 33.4905
R1235 B.n917 B.n916 33.4905
R1236 B.n916 B.n915 33.4905
R1237 B.n915 B.n58 33.4905
R1238 B.n909 B.n58 33.4905
R1239 B.n909 B.n908 33.4905
R1240 B.n908 B.n907 33.4905
R1241 B.n585 B.t4 32.998
R1242 B.n955 B.t2 32.998
R1243 B.n659 B.n658 29.8151
R1244 B.n510 B.n509 29.8151
R1245 B.n514 B.n196 29.8151
R1246 B.n905 B.n904 29.8151
R1247 B.n530 B.t7 21.178
R1248 B.n917 B.t14 21.178
R1249 B.n143 B.t3 20.193
R1250 B.t1 B.n964 20.193
R1251 B.t5 B.n162 19.208
R1252 B.n940 B.t0 19.208
R1253 B B.n977 18.0485
R1254 B.n560 B.t5 14.283
R1255 B.t0 B.n939 14.283
R1256 B.n604 B.t3 13.298
R1257 B.n965 B.t1 13.298
R1258 B.t7 B.n182 12.313
R1259 B.t14 B.n51 12.313
R1260 B.n510 B.n192 10.6151
R1261 B.n520 B.n192 10.6151
R1262 B.n521 B.n520 10.6151
R1263 B.n522 B.n521 10.6151
R1264 B.n522 B.n184 10.6151
R1265 B.n532 B.n184 10.6151
R1266 B.n533 B.n532 10.6151
R1267 B.n534 B.n533 10.6151
R1268 B.n534 B.n176 10.6151
R1269 B.n544 B.n176 10.6151
R1270 B.n545 B.n544 10.6151
R1271 B.n546 B.n545 10.6151
R1272 B.n546 B.n168 10.6151
R1273 B.n556 B.n168 10.6151
R1274 B.n557 B.n556 10.6151
R1275 B.n558 B.n557 10.6151
R1276 B.n558 B.n160 10.6151
R1277 B.n568 B.n160 10.6151
R1278 B.n569 B.n568 10.6151
R1279 B.n570 B.n569 10.6151
R1280 B.n570 B.n152 10.6151
R1281 B.n581 B.n152 10.6151
R1282 B.n582 B.n581 10.6151
R1283 B.n583 B.n582 10.6151
R1284 B.n583 B.n145 10.6151
R1285 B.n593 B.n145 10.6151
R1286 B.n594 B.n593 10.6151
R1287 B.n595 B.n594 10.6151
R1288 B.n595 B.n137 10.6151
R1289 B.n606 B.n137 10.6151
R1290 B.n607 B.n606 10.6151
R1291 B.n608 B.n607 10.6151
R1292 B.n608 B.n0 10.6151
R1293 B.n509 B.n508 10.6151
R1294 B.n508 B.n200 10.6151
R1295 B.n503 B.n200 10.6151
R1296 B.n503 B.n502 10.6151
R1297 B.n502 B.n202 10.6151
R1298 B.n497 B.n202 10.6151
R1299 B.n497 B.n496 10.6151
R1300 B.n496 B.n495 10.6151
R1301 B.n495 B.n204 10.6151
R1302 B.n489 B.n204 10.6151
R1303 B.n489 B.n488 10.6151
R1304 B.n488 B.n487 10.6151
R1305 B.n487 B.n206 10.6151
R1306 B.n481 B.n206 10.6151
R1307 B.n481 B.n480 10.6151
R1308 B.n480 B.n479 10.6151
R1309 B.n479 B.n208 10.6151
R1310 B.n473 B.n208 10.6151
R1311 B.n473 B.n472 10.6151
R1312 B.n472 B.n471 10.6151
R1313 B.n471 B.n210 10.6151
R1314 B.n465 B.n210 10.6151
R1315 B.n465 B.n464 10.6151
R1316 B.n464 B.n463 10.6151
R1317 B.n463 B.n212 10.6151
R1318 B.n457 B.n212 10.6151
R1319 B.n457 B.n456 10.6151
R1320 B.n456 B.n455 10.6151
R1321 B.n455 B.n214 10.6151
R1322 B.n449 B.n214 10.6151
R1323 B.n449 B.n448 10.6151
R1324 B.n448 B.n447 10.6151
R1325 B.n447 B.n216 10.6151
R1326 B.n441 B.n216 10.6151
R1327 B.n441 B.n440 10.6151
R1328 B.n440 B.n439 10.6151
R1329 B.n439 B.n218 10.6151
R1330 B.n433 B.n218 10.6151
R1331 B.n433 B.n432 10.6151
R1332 B.n432 B.n431 10.6151
R1333 B.n431 B.n220 10.6151
R1334 B.n425 B.n220 10.6151
R1335 B.n425 B.n424 10.6151
R1336 B.n424 B.n423 10.6151
R1337 B.n423 B.n222 10.6151
R1338 B.n417 B.n222 10.6151
R1339 B.n417 B.n416 10.6151
R1340 B.n416 B.n415 10.6151
R1341 B.n415 B.n224 10.6151
R1342 B.n409 B.n224 10.6151
R1343 B.n409 B.n408 10.6151
R1344 B.n408 B.n407 10.6151
R1345 B.n407 B.n226 10.6151
R1346 B.n401 B.n226 10.6151
R1347 B.n401 B.n400 10.6151
R1348 B.n400 B.n399 10.6151
R1349 B.n395 B.n394 10.6151
R1350 B.n394 B.n232 10.6151
R1351 B.n389 B.n232 10.6151
R1352 B.n389 B.n388 10.6151
R1353 B.n388 B.n387 10.6151
R1354 B.n387 B.n234 10.6151
R1355 B.n381 B.n234 10.6151
R1356 B.n381 B.n380 10.6151
R1357 B.n378 B.n238 10.6151
R1358 B.n372 B.n238 10.6151
R1359 B.n372 B.n371 10.6151
R1360 B.n371 B.n370 10.6151
R1361 B.n370 B.n240 10.6151
R1362 B.n364 B.n240 10.6151
R1363 B.n364 B.n363 10.6151
R1364 B.n363 B.n362 10.6151
R1365 B.n362 B.n242 10.6151
R1366 B.n356 B.n242 10.6151
R1367 B.n356 B.n355 10.6151
R1368 B.n355 B.n354 10.6151
R1369 B.n354 B.n244 10.6151
R1370 B.n348 B.n244 10.6151
R1371 B.n348 B.n347 10.6151
R1372 B.n347 B.n346 10.6151
R1373 B.n346 B.n246 10.6151
R1374 B.n340 B.n246 10.6151
R1375 B.n340 B.n339 10.6151
R1376 B.n339 B.n338 10.6151
R1377 B.n338 B.n248 10.6151
R1378 B.n332 B.n248 10.6151
R1379 B.n332 B.n331 10.6151
R1380 B.n331 B.n330 10.6151
R1381 B.n330 B.n250 10.6151
R1382 B.n324 B.n250 10.6151
R1383 B.n324 B.n323 10.6151
R1384 B.n323 B.n322 10.6151
R1385 B.n322 B.n252 10.6151
R1386 B.n316 B.n252 10.6151
R1387 B.n316 B.n315 10.6151
R1388 B.n315 B.n314 10.6151
R1389 B.n314 B.n254 10.6151
R1390 B.n308 B.n254 10.6151
R1391 B.n308 B.n307 10.6151
R1392 B.n307 B.n306 10.6151
R1393 B.n306 B.n256 10.6151
R1394 B.n300 B.n256 10.6151
R1395 B.n300 B.n299 10.6151
R1396 B.n299 B.n298 10.6151
R1397 B.n298 B.n258 10.6151
R1398 B.n292 B.n258 10.6151
R1399 B.n292 B.n291 10.6151
R1400 B.n291 B.n290 10.6151
R1401 B.n290 B.n260 10.6151
R1402 B.n284 B.n260 10.6151
R1403 B.n284 B.n283 10.6151
R1404 B.n283 B.n282 10.6151
R1405 B.n282 B.n262 10.6151
R1406 B.n276 B.n262 10.6151
R1407 B.n276 B.n275 10.6151
R1408 B.n275 B.n274 10.6151
R1409 B.n274 B.n264 10.6151
R1410 B.n268 B.n264 10.6151
R1411 B.n268 B.n267 10.6151
R1412 B.n267 B.n196 10.6151
R1413 B.n515 B.n514 10.6151
R1414 B.n516 B.n515 10.6151
R1415 B.n516 B.n188 10.6151
R1416 B.n526 B.n188 10.6151
R1417 B.n527 B.n526 10.6151
R1418 B.n528 B.n527 10.6151
R1419 B.n528 B.n180 10.6151
R1420 B.n538 B.n180 10.6151
R1421 B.n539 B.n538 10.6151
R1422 B.n540 B.n539 10.6151
R1423 B.n540 B.n172 10.6151
R1424 B.n550 B.n172 10.6151
R1425 B.n551 B.n550 10.6151
R1426 B.n552 B.n551 10.6151
R1427 B.n552 B.n164 10.6151
R1428 B.n562 B.n164 10.6151
R1429 B.n563 B.n562 10.6151
R1430 B.n564 B.n563 10.6151
R1431 B.n564 B.n156 10.6151
R1432 B.n574 B.n156 10.6151
R1433 B.n575 B.n574 10.6151
R1434 B.n576 B.n575 10.6151
R1435 B.n576 B.n149 10.6151
R1436 B.n587 B.n149 10.6151
R1437 B.n588 B.n587 10.6151
R1438 B.n589 B.n588 10.6151
R1439 B.n589 B.n140 10.6151
R1440 B.n599 B.n140 10.6151
R1441 B.n600 B.n599 10.6151
R1442 B.n602 B.n600 10.6151
R1443 B.n602 B.n601 10.6151
R1444 B.n601 B.n133 10.6151
R1445 B.n613 B.n133 10.6151
R1446 B.n614 B.n613 10.6151
R1447 B.n615 B.n614 10.6151
R1448 B.n616 B.n615 10.6151
R1449 B.n617 B.n616 10.6151
R1450 B.n620 B.n617 10.6151
R1451 B.n621 B.n620 10.6151
R1452 B.n622 B.n621 10.6151
R1453 B.n623 B.n622 10.6151
R1454 B.n625 B.n623 10.6151
R1455 B.n626 B.n625 10.6151
R1456 B.n627 B.n626 10.6151
R1457 B.n628 B.n627 10.6151
R1458 B.n630 B.n628 10.6151
R1459 B.n631 B.n630 10.6151
R1460 B.n632 B.n631 10.6151
R1461 B.n633 B.n632 10.6151
R1462 B.n635 B.n633 10.6151
R1463 B.n636 B.n635 10.6151
R1464 B.n637 B.n636 10.6151
R1465 B.n638 B.n637 10.6151
R1466 B.n640 B.n638 10.6151
R1467 B.n641 B.n640 10.6151
R1468 B.n642 B.n641 10.6151
R1469 B.n643 B.n642 10.6151
R1470 B.n645 B.n643 10.6151
R1471 B.n646 B.n645 10.6151
R1472 B.n647 B.n646 10.6151
R1473 B.n648 B.n647 10.6151
R1474 B.n650 B.n648 10.6151
R1475 B.n651 B.n650 10.6151
R1476 B.n652 B.n651 10.6151
R1477 B.n653 B.n652 10.6151
R1478 B.n655 B.n653 10.6151
R1479 B.n656 B.n655 10.6151
R1480 B.n657 B.n656 10.6151
R1481 B.n658 B.n657 10.6151
R1482 B.n969 B.n1 10.6151
R1483 B.n969 B.n968 10.6151
R1484 B.n968 B.n967 10.6151
R1485 B.n967 B.n10 10.6151
R1486 B.n961 B.n10 10.6151
R1487 B.n961 B.n960 10.6151
R1488 B.n960 B.n959 10.6151
R1489 B.n959 B.n18 10.6151
R1490 B.n953 B.n18 10.6151
R1491 B.n953 B.n952 10.6151
R1492 B.n952 B.n951 10.6151
R1493 B.n951 B.n24 10.6151
R1494 B.n945 B.n24 10.6151
R1495 B.n945 B.n944 10.6151
R1496 B.n944 B.n943 10.6151
R1497 B.n943 B.n32 10.6151
R1498 B.n937 B.n32 10.6151
R1499 B.n937 B.n936 10.6151
R1500 B.n936 B.n935 10.6151
R1501 B.n935 B.n39 10.6151
R1502 B.n929 B.n39 10.6151
R1503 B.n929 B.n928 10.6151
R1504 B.n928 B.n927 10.6151
R1505 B.n927 B.n46 10.6151
R1506 B.n921 B.n46 10.6151
R1507 B.n921 B.n920 10.6151
R1508 B.n920 B.n919 10.6151
R1509 B.n919 B.n53 10.6151
R1510 B.n913 B.n53 10.6151
R1511 B.n913 B.n912 10.6151
R1512 B.n912 B.n911 10.6151
R1513 B.n911 B.n60 10.6151
R1514 B.n905 B.n60 10.6151
R1515 B.n904 B.n903 10.6151
R1516 B.n903 B.n67 10.6151
R1517 B.n897 B.n67 10.6151
R1518 B.n897 B.n896 10.6151
R1519 B.n896 B.n895 10.6151
R1520 B.n895 B.n69 10.6151
R1521 B.n889 B.n69 10.6151
R1522 B.n889 B.n888 10.6151
R1523 B.n888 B.n887 10.6151
R1524 B.n887 B.n71 10.6151
R1525 B.n881 B.n71 10.6151
R1526 B.n881 B.n880 10.6151
R1527 B.n880 B.n879 10.6151
R1528 B.n879 B.n73 10.6151
R1529 B.n873 B.n73 10.6151
R1530 B.n873 B.n872 10.6151
R1531 B.n872 B.n871 10.6151
R1532 B.n871 B.n75 10.6151
R1533 B.n865 B.n75 10.6151
R1534 B.n865 B.n864 10.6151
R1535 B.n864 B.n863 10.6151
R1536 B.n863 B.n77 10.6151
R1537 B.n857 B.n77 10.6151
R1538 B.n857 B.n856 10.6151
R1539 B.n856 B.n855 10.6151
R1540 B.n855 B.n79 10.6151
R1541 B.n849 B.n79 10.6151
R1542 B.n849 B.n848 10.6151
R1543 B.n848 B.n847 10.6151
R1544 B.n847 B.n81 10.6151
R1545 B.n841 B.n81 10.6151
R1546 B.n841 B.n840 10.6151
R1547 B.n840 B.n839 10.6151
R1548 B.n839 B.n83 10.6151
R1549 B.n833 B.n83 10.6151
R1550 B.n833 B.n832 10.6151
R1551 B.n832 B.n831 10.6151
R1552 B.n831 B.n85 10.6151
R1553 B.n825 B.n85 10.6151
R1554 B.n825 B.n824 10.6151
R1555 B.n824 B.n823 10.6151
R1556 B.n823 B.n87 10.6151
R1557 B.n817 B.n87 10.6151
R1558 B.n817 B.n816 10.6151
R1559 B.n816 B.n815 10.6151
R1560 B.n815 B.n89 10.6151
R1561 B.n809 B.n89 10.6151
R1562 B.n809 B.n808 10.6151
R1563 B.n808 B.n807 10.6151
R1564 B.n807 B.n91 10.6151
R1565 B.n801 B.n91 10.6151
R1566 B.n801 B.n800 10.6151
R1567 B.n800 B.n799 10.6151
R1568 B.n799 B.n93 10.6151
R1569 B.n793 B.n93 10.6151
R1570 B.n793 B.n792 10.6151
R1571 B.n790 B.n97 10.6151
R1572 B.n784 B.n97 10.6151
R1573 B.n784 B.n783 10.6151
R1574 B.n783 B.n782 10.6151
R1575 B.n782 B.n99 10.6151
R1576 B.n776 B.n99 10.6151
R1577 B.n776 B.n775 10.6151
R1578 B.n775 B.n774 10.6151
R1579 B.n770 B.n769 10.6151
R1580 B.n769 B.n105 10.6151
R1581 B.n764 B.n105 10.6151
R1582 B.n764 B.n763 10.6151
R1583 B.n763 B.n762 10.6151
R1584 B.n762 B.n107 10.6151
R1585 B.n756 B.n107 10.6151
R1586 B.n756 B.n755 10.6151
R1587 B.n755 B.n754 10.6151
R1588 B.n754 B.n109 10.6151
R1589 B.n748 B.n109 10.6151
R1590 B.n748 B.n747 10.6151
R1591 B.n747 B.n746 10.6151
R1592 B.n746 B.n111 10.6151
R1593 B.n740 B.n111 10.6151
R1594 B.n740 B.n739 10.6151
R1595 B.n739 B.n738 10.6151
R1596 B.n738 B.n113 10.6151
R1597 B.n732 B.n113 10.6151
R1598 B.n732 B.n731 10.6151
R1599 B.n731 B.n730 10.6151
R1600 B.n730 B.n115 10.6151
R1601 B.n724 B.n115 10.6151
R1602 B.n724 B.n723 10.6151
R1603 B.n723 B.n722 10.6151
R1604 B.n722 B.n117 10.6151
R1605 B.n716 B.n117 10.6151
R1606 B.n716 B.n715 10.6151
R1607 B.n715 B.n714 10.6151
R1608 B.n714 B.n119 10.6151
R1609 B.n708 B.n119 10.6151
R1610 B.n708 B.n707 10.6151
R1611 B.n707 B.n706 10.6151
R1612 B.n706 B.n121 10.6151
R1613 B.n700 B.n121 10.6151
R1614 B.n700 B.n699 10.6151
R1615 B.n699 B.n698 10.6151
R1616 B.n698 B.n123 10.6151
R1617 B.n692 B.n123 10.6151
R1618 B.n692 B.n691 10.6151
R1619 B.n691 B.n690 10.6151
R1620 B.n690 B.n125 10.6151
R1621 B.n684 B.n125 10.6151
R1622 B.n684 B.n683 10.6151
R1623 B.n683 B.n682 10.6151
R1624 B.n682 B.n127 10.6151
R1625 B.n676 B.n127 10.6151
R1626 B.n676 B.n675 10.6151
R1627 B.n675 B.n674 10.6151
R1628 B.n674 B.n129 10.6151
R1629 B.n668 B.n129 10.6151
R1630 B.n668 B.n667 10.6151
R1631 B.n667 B.n666 10.6151
R1632 B.n666 B.n131 10.6151
R1633 B.n660 B.n131 10.6151
R1634 B.n660 B.n659 10.6151
R1635 B.n977 B.n0 8.11757
R1636 B.n977 B.n1 8.11757
R1637 B.n395 B.n230 6.5566
R1638 B.n380 B.n379 6.5566
R1639 B.n791 B.n790 6.5566
R1640 B.n774 B.n103 6.5566
R1641 B.n399 B.n230 4.05904
R1642 B.n379 B.n378 4.05904
R1643 B.n792 B.n791 4.05904
R1644 B.n770 B.n103 4.05904
R1645 B.n578 B.t4 0.493001
R1646 B.n26 B.t2 0.493001
R1647 VP.n6 VP.t0 246.653
R1648 VP.n17 VP.t2 215.261
R1649 VP.n24 VP.t5 215.261
R1650 VP.n31 VP.t4 215.261
R1651 VP.n14 VP.t3 215.261
R1652 VP.n7 VP.t1 215.261
R1653 VP.n9 VP.n8 161.3
R1654 VP.n10 VP.n5 161.3
R1655 VP.n12 VP.n11 161.3
R1656 VP.n13 VP.n4 161.3
R1657 VP.n30 VP.n0 161.3
R1658 VP.n29 VP.n28 161.3
R1659 VP.n27 VP.n1 161.3
R1660 VP.n26 VP.n25 161.3
R1661 VP.n23 VP.n2 161.3
R1662 VP.n22 VP.n21 161.3
R1663 VP.n20 VP.n3 161.3
R1664 VP.n19 VP.n18 161.3
R1665 VP.n17 VP.n16 86.8082
R1666 VP.n32 VP.n31 86.8082
R1667 VP.n15 VP.n14 86.8082
R1668 VP.n7 VP.n6 58.0461
R1669 VP.n22 VP.n3 53.171
R1670 VP.n29 VP.n1 53.171
R1671 VP.n12 VP.n5 53.171
R1672 VP.n16 VP.n15 49.8709
R1673 VP.n18 VP.n3 27.983
R1674 VP.n30 VP.n29 27.983
R1675 VP.n13 VP.n12 27.983
R1676 VP.n23 VP.n22 24.5923
R1677 VP.n25 VP.n1 24.5923
R1678 VP.n8 VP.n5 24.5923
R1679 VP.n18 VP.n17 24.1005
R1680 VP.n31 VP.n30 24.1005
R1681 VP.n14 VP.n13 24.1005
R1682 VP.n9 VP.n6 12.6777
R1683 VP.n24 VP.n23 12.2964
R1684 VP.n25 VP.n24 12.2964
R1685 VP.n8 VP.n7 12.2964
R1686 VP.n15 VP.n4 0.278335
R1687 VP.n19 VP.n16 0.278335
R1688 VP.n32 VP.n0 0.278335
R1689 VP.n10 VP.n9 0.189894
R1690 VP.n11 VP.n10 0.189894
R1691 VP.n11 VP.n4 0.189894
R1692 VP.n20 VP.n19 0.189894
R1693 VP.n21 VP.n20 0.189894
R1694 VP.n21 VP.n2 0.189894
R1695 VP.n26 VP.n2 0.189894
R1696 VP.n27 VP.n26 0.189894
R1697 VP.n28 VP.n27 0.189894
R1698 VP.n28 VP.n0 0.189894
R1699 VP VP.n32 0.153485
R1700 VTAIL.n7 VTAIL.t2 43.2444
R1701 VTAIL.n11 VTAIL.t1 43.2443
R1702 VTAIL.n2 VTAIL.t7 43.2443
R1703 VTAIL.n10 VTAIL.t9 43.2443
R1704 VTAIL.n9 VTAIL.n8 42.0839
R1705 VTAIL.n6 VTAIL.n5 42.0839
R1706 VTAIL.n1 VTAIL.n0 42.0836
R1707 VTAIL.n4 VTAIL.n3 42.0836
R1708 VTAIL.n6 VTAIL.n4 30.9358
R1709 VTAIL.n11 VTAIL.n10 29.0048
R1710 VTAIL.n7 VTAIL.n6 1.93153
R1711 VTAIL.n10 VTAIL.n9 1.93153
R1712 VTAIL.n4 VTAIL.n2 1.93153
R1713 VTAIL.n9 VTAIL.n7 1.43584
R1714 VTAIL.n2 VTAIL.n1 1.43584
R1715 VTAIL VTAIL.n11 1.39059
R1716 VTAIL.n0 VTAIL.t0 1.16111
R1717 VTAIL.n0 VTAIL.t4 1.16111
R1718 VTAIL.n3 VTAIL.t8 1.16111
R1719 VTAIL.n3 VTAIL.t5 1.16111
R1720 VTAIL.n8 VTAIL.t10 1.16111
R1721 VTAIL.n8 VTAIL.t6 1.16111
R1722 VTAIL.n5 VTAIL.t11 1.16111
R1723 VTAIL.n5 VTAIL.t3 1.16111
R1724 VTAIL VTAIL.n1 0.541448
R1725 VDD1 VDD1.t5 61.4297
R1726 VDD1.n1 VDD1.t3 61.316
R1727 VDD1.n1 VDD1.n0 59.1898
R1728 VDD1.n3 VDD1.n2 58.7625
R1729 VDD1.n3 VDD1.n1 46.2466
R1730 VDD1.n2 VDD1.t4 1.16111
R1731 VDD1.n2 VDD1.t2 1.16111
R1732 VDD1.n0 VDD1.t0 1.16111
R1733 VDD1.n0 VDD1.t1 1.16111
R1734 VDD1 VDD1.n3 0.425069
R1735 VN.n2 VN.t3 246.653
R1736 VN.n14 VN.t2 246.653
R1737 VN.n3 VN.t5 215.261
R1738 VN.n10 VN.t1 215.261
R1739 VN.n15 VN.t4 215.261
R1740 VN.n22 VN.t0 215.261
R1741 VN.n21 VN.n12 161.3
R1742 VN.n20 VN.n19 161.3
R1743 VN.n18 VN.n13 161.3
R1744 VN.n17 VN.n16 161.3
R1745 VN.n9 VN.n0 161.3
R1746 VN.n8 VN.n7 161.3
R1747 VN.n6 VN.n1 161.3
R1748 VN.n5 VN.n4 161.3
R1749 VN.n11 VN.n10 86.8082
R1750 VN.n23 VN.n22 86.8082
R1751 VN.n3 VN.n2 58.0461
R1752 VN.n15 VN.n14 58.0461
R1753 VN.n8 VN.n1 53.171
R1754 VN.n20 VN.n13 53.171
R1755 VN VN.n23 50.1497
R1756 VN.n9 VN.n8 27.983
R1757 VN.n21 VN.n20 27.983
R1758 VN.n4 VN.n1 24.5923
R1759 VN.n16 VN.n13 24.5923
R1760 VN.n10 VN.n9 24.1005
R1761 VN.n22 VN.n21 24.1005
R1762 VN.n17 VN.n14 12.6777
R1763 VN.n5 VN.n2 12.6777
R1764 VN.n4 VN.n3 12.2964
R1765 VN.n16 VN.n15 12.2964
R1766 VN.n23 VN.n12 0.278335
R1767 VN.n11 VN.n0 0.278335
R1768 VN.n19 VN.n12 0.189894
R1769 VN.n19 VN.n18 0.189894
R1770 VN.n18 VN.n17 0.189894
R1771 VN.n6 VN.n5 0.189894
R1772 VN.n7 VN.n6 0.189894
R1773 VN.n7 VN.n0 0.189894
R1774 VN VN.n11 0.153485
R1775 VDD2.n1 VDD2.t2 61.316
R1776 VDD2.n2 VDD2.t5 59.9232
R1777 VDD2.n1 VDD2.n0 59.1898
R1778 VDD2 VDD2.n3 59.1871
R1779 VDD2.n2 VDD2.n1 44.6981
R1780 VDD2 VDD2.n2 1.50697
R1781 VDD2.n3 VDD2.t1 1.16111
R1782 VDD2.n3 VDD2.t3 1.16111
R1783 VDD2.n0 VDD2.t0 1.16111
R1784 VDD2.n0 VDD2.t4 1.16111
C0 VDD1 VDD2 1.1633f
C1 VDD2 VTAIL 9.8776f
C2 VDD1 VTAIL 9.83386f
C3 VP VN 7.18937f
C4 VN VDD2 8.779281f
C5 VDD1 VN 0.15013f
C6 VN VTAIL 8.568081f
C7 VP VDD2 0.400707f
C8 VDD1 VP 9.02531f
C9 VP VTAIL 8.582549f
C10 VDD2 B 6.33739f
C11 VDD1 B 6.627405f
C12 VTAIL B 9.33319f
C13 VN B 11.39893f
C14 VP B 9.771539f
C15 VDD2.t2 B 3.36071f
C16 VDD2.t0 B 0.289047f
C17 VDD2.t4 B 0.289047f
C18 VDD2.n0 B 2.62762f
C19 VDD2.n1 B 2.51692f
C20 VDD2.t5 B 3.35287f
C21 VDD2.n2 B 2.57603f
C22 VDD2.t1 B 0.289047f
C23 VDD2.t3 B 0.289047f
C24 VDD2.n3 B 2.62758f
C25 VN.n0 B 0.036185f
C26 VN.t1 B 2.45749f
C27 VN.n1 B 0.048468f
C28 VN.t3 B 2.584f
C29 VN.n2 B 0.931657f
C30 VN.t5 B 2.45749f
C31 VN.n3 B 0.923974f
C32 VN.n4 B 0.038336f
C33 VN.n5 B 0.203131f
C34 VN.n6 B 0.027448f
C35 VN.n7 B 0.027448f
C36 VN.n8 B 0.028713f
C37 VN.n9 B 0.053015f
C38 VN.n10 B 0.947568f
C39 VN.n11 B 0.029433f
C40 VN.n12 B 0.036185f
C41 VN.t0 B 2.45749f
C42 VN.n13 B 0.048468f
C43 VN.t2 B 2.584f
C44 VN.n14 B 0.931657f
C45 VN.t4 B 2.45749f
C46 VN.n15 B 0.923974f
C47 VN.n16 B 0.038336f
C48 VN.n17 B 0.203131f
C49 VN.n18 B 0.027448f
C50 VN.n19 B 0.027448f
C51 VN.n20 B 0.028713f
C52 VN.n21 B 0.053015f
C53 VN.n22 B 0.947568f
C54 VN.n23 B 1.52061f
C55 VDD1.t5 B 3.36526f
C56 VDD1.t3 B 3.36443f
C57 VDD1.t0 B 0.289367f
C58 VDD1.t1 B 0.289367f
C59 VDD1.n0 B 2.63053f
C60 VDD1.n1 B 2.61352f
C61 VDD1.t4 B 0.289367f
C62 VDD1.t2 B 0.289367f
C63 VDD1.n2 B 2.62797f
C64 VDD1.n3 B 2.56252f
C65 VTAIL.t0 B 0.303308f
C66 VTAIL.t4 B 0.303308f
C67 VTAIL.n0 B 2.6815f
C68 VTAIL.n1 B 0.374454f
C69 VTAIL.t7 B 3.42267f
C70 VTAIL.n2 B 0.561266f
C71 VTAIL.t8 B 0.303308f
C72 VTAIL.t5 B 0.303308f
C73 VTAIL.n3 B 2.6815f
C74 VTAIL.n4 B 2.02294f
C75 VTAIL.t11 B 0.303308f
C76 VTAIL.t3 B 0.303308f
C77 VTAIL.n5 B 2.68151f
C78 VTAIL.n6 B 2.02294f
C79 VTAIL.t2 B 3.42269f
C80 VTAIL.n7 B 0.561244f
C81 VTAIL.t10 B 0.303308f
C82 VTAIL.t6 B 0.303308f
C83 VTAIL.n8 B 2.68151f
C84 VTAIL.n9 B 0.475224f
C85 VTAIL.t9 B 3.42267f
C86 VTAIL.n10 B 1.96899f
C87 VTAIL.t1 B 3.42267f
C88 VTAIL.n11 B 1.92977f
C89 VP.n0 B 0.036537f
C90 VP.t4 B 2.48136f
C91 VP.n1 B 0.048939f
C92 VP.n2 B 0.027715f
C93 VP.t5 B 2.48136f
C94 VP.n3 B 0.028991f
C95 VP.n4 B 0.036537f
C96 VP.t3 B 2.48136f
C97 VP.n5 B 0.048939f
C98 VP.t0 B 2.6091f
C99 VP.n6 B 0.940707f
C100 VP.t1 B 2.48136f
C101 VP.n7 B 0.932949f
C102 VP.n8 B 0.038708f
C103 VP.n9 B 0.205105f
C104 VP.n10 B 0.027715f
C105 VP.n11 B 0.027715f
C106 VP.n12 B 0.028991f
C107 VP.n13 B 0.05353f
C108 VP.n14 B 0.956772f
C109 VP.n15 B 1.52049f
C110 VP.n16 B 1.54052f
C111 VP.t2 B 2.48136f
C112 VP.n17 B 0.956772f
C113 VP.n18 B 0.05353f
C114 VP.n19 B 0.036537f
C115 VP.n20 B 0.027715f
C116 VP.n21 B 0.027715f
C117 VP.n22 B 0.048939f
C118 VP.n23 B 0.038708f
C119 VP.n24 B 0.868976f
C120 VP.n25 B 0.038708f
C121 VP.n26 B 0.027715f
C122 VP.n27 B 0.027715f
C123 VP.n28 B 0.027715f
C124 VP.n29 B 0.028991f
C125 VP.n30 B 0.05353f
C126 VP.n31 B 0.956772f
C127 VP.n32 B 0.029719f
.ends

