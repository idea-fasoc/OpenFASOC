* NGSPICE file created from diff_pair_sample_0296.ext - technology: sky130A

.subckt diff_pair_sample_0296 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=0.62
X2 VDD1.t7 VP.t0 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X3 VDD2.t3 VN.t1 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=0.62
X4 VTAIL.t8 VN.t2 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X5 VDD1.t6 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=0.62
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=0.62
X7 VDD1.t5 VP.t2 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=0.62
X8 VTAIL.t15 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=0.62
X9 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X10 VDD1.t2 VP.t5 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=0.62
X12 VTAIL.t13 VP.t6 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=0.62
X13 VTAIL.t7 VN.t3 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=0.62
X14 VDD2.t7 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=0.62
X15 VTAIL.t2 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=0.62
X17 VTAIL.t5 VN.t5 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=0.62
X18 VDD2.t1 VN.t6 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
X19 VDD2.t0 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=0.62
R0 VN.n1 VN.t5 653.811
R1 VN.n7 VN.t4 653.811
R2 VN.n2 VN.t7 626.99
R3 VN.n3 VN.t0 626.99
R4 VN.n4 VN.t1 626.99
R5 VN.n8 VN.t2 626.99
R6 VN.n9 VN.t6 626.99
R7 VN.n10 VN.t3 626.99
R8 VN.n5 VN.n4 161.3
R9 VN.n11 VN.n10 161.3
R10 VN.n9 VN.n6 80.6037
R11 VN.n3 VN.n0 80.6037
R12 VN.n3 VN.n2 48.2005
R13 VN.n4 VN.n3 48.2005
R14 VN.n9 VN.n8 48.2005
R15 VN.n10 VN.n9 48.2005
R16 VN.n7 VN.n6 45.2318
R17 VN.n1 VN.n0 45.2318
R18 VN VN.n11 43.9721
R19 VN.n8 VN.n7 13.3799
R20 VN.n2 VN.n1 13.3799
R21 VN.n11 VN.n6 0.285035
R22 VN.n5 VN.n0 0.285035
R23 VN VN.n5 0.0516364
R24 VDD2.n2 VDD2.n1 65.5865
R25 VDD2.n2 VDD2.n0 65.5865
R26 VDD2 VDD2.n5 65.5837
R27 VDD2.n4 VDD2.n3 65.2326
R28 VDD2.n4 VDD2.n2 39.9006
R29 VDD2.n5 VDD2.t2 1.36602
R30 VDD2.n5 VDD2.t7 1.36602
R31 VDD2.n3 VDD2.t5 1.36602
R32 VDD2.n3 VDD2.t1 1.36602
R33 VDD2.n1 VDD2.t4 1.36602
R34 VDD2.n1 VDD2.t3 1.36602
R35 VDD2.n0 VDD2.t6 1.36602
R36 VDD2.n0 VDD2.t0 1.36602
R37 VDD2 VDD2.n4 0.468172
R38 VTAIL.n11 VTAIL.t15 49.9192
R39 VTAIL.n10 VTAIL.t6 49.9192
R40 VTAIL.n7 VTAIL.t7 49.9192
R41 VTAIL.n15 VTAIL.t9 49.9191
R42 VTAIL.n2 VTAIL.t5 49.9191
R43 VTAIL.n3 VTAIL.t0 49.9191
R44 VTAIL.n6 VTAIL.t13 49.9191
R45 VTAIL.n14 VTAIL.t12 49.9191
R46 VTAIL.n13 VTAIL.n12 48.5538
R47 VTAIL.n9 VTAIL.n8 48.5538
R48 VTAIL.n1 VTAIL.n0 48.5535
R49 VTAIL.n5 VTAIL.n4 48.5535
R50 VTAIL.n15 VTAIL.n14 25.6858
R51 VTAIL.n7 VTAIL.n6 25.6858
R52 VTAIL.n0 VTAIL.t3 1.36602
R53 VTAIL.n0 VTAIL.t10 1.36602
R54 VTAIL.n4 VTAIL.t14 1.36602
R55 VTAIL.n4 VTAIL.t1 1.36602
R56 VTAIL.n12 VTAIL.t11 1.36602
R57 VTAIL.n12 VTAIL.t2 1.36602
R58 VTAIL.n8 VTAIL.t4 1.36602
R59 VTAIL.n8 VTAIL.t8 1.36602
R60 VTAIL.n9 VTAIL.n7 0.819465
R61 VTAIL.n10 VTAIL.n9 0.819465
R62 VTAIL.n13 VTAIL.n11 0.819465
R63 VTAIL.n14 VTAIL.n13 0.819465
R64 VTAIL.n6 VTAIL.n5 0.819465
R65 VTAIL.n5 VTAIL.n3 0.819465
R66 VTAIL.n2 VTAIL.n1 0.819465
R67 VTAIL VTAIL.n15 0.761276
R68 VTAIL.n11 VTAIL.n10 0.470328
R69 VTAIL.n3 VTAIL.n2 0.470328
R70 VTAIL VTAIL.n1 0.0586897
R71 B.n177 B.t16 767.705
R72 B.n169 B.t8 767.705
R73 B.n68 B.t12 767.705
R74 B.n76 B.t19 767.705
R75 B.n513 B.n512 585
R76 B.n515 B.n101 585
R77 B.n518 B.n517 585
R78 B.n519 B.n100 585
R79 B.n521 B.n520 585
R80 B.n523 B.n99 585
R81 B.n526 B.n525 585
R82 B.n527 B.n98 585
R83 B.n529 B.n528 585
R84 B.n531 B.n97 585
R85 B.n534 B.n533 585
R86 B.n535 B.n96 585
R87 B.n537 B.n536 585
R88 B.n539 B.n95 585
R89 B.n542 B.n541 585
R90 B.n543 B.n94 585
R91 B.n545 B.n544 585
R92 B.n547 B.n93 585
R93 B.n550 B.n549 585
R94 B.n551 B.n92 585
R95 B.n553 B.n552 585
R96 B.n555 B.n91 585
R97 B.n558 B.n557 585
R98 B.n559 B.n90 585
R99 B.n561 B.n560 585
R100 B.n563 B.n89 585
R101 B.n566 B.n565 585
R102 B.n567 B.n88 585
R103 B.n569 B.n568 585
R104 B.n571 B.n87 585
R105 B.n574 B.n573 585
R106 B.n575 B.n86 585
R107 B.n577 B.n576 585
R108 B.n579 B.n85 585
R109 B.n582 B.n581 585
R110 B.n583 B.n84 585
R111 B.n585 B.n584 585
R112 B.n587 B.n83 585
R113 B.n590 B.n589 585
R114 B.n591 B.n82 585
R115 B.n593 B.n592 585
R116 B.n595 B.n81 585
R117 B.n598 B.n597 585
R118 B.n599 B.n80 585
R119 B.n601 B.n600 585
R120 B.n603 B.n79 585
R121 B.n606 B.n605 585
R122 B.n607 B.n75 585
R123 B.n609 B.n608 585
R124 B.n611 B.n74 585
R125 B.n614 B.n613 585
R126 B.n615 B.n73 585
R127 B.n617 B.n616 585
R128 B.n619 B.n72 585
R129 B.n622 B.n621 585
R130 B.n623 B.n71 585
R131 B.n625 B.n624 585
R132 B.n627 B.n70 585
R133 B.n630 B.n629 585
R134 B.n632 B.n67 585
R135 B.n634 B.n633 585
R136 B.n636 B.n66 585
R137 B.n639 B.n638 585
R138 B.n640 B.n65 585
R139 B.n642 B.n641 585
R140 B.n644 B.n64 585
R141 B.n647 B.n646 585
R142 B.n648 B.n63 585
R143 B.n650 B.n649 585
R144 B.n652 B.n62 585
R145 B.n655 B.n654 585
R146 B.n656 B.n61 585
R147 B.n658 B.n657 585
R148 B.n660 B.n60 585
R149 B.n663 B.n662 585
R150 B.n664 B.n59 585
R151 B.n666 B.n665 585
R152 B.n668 B.n58 585
R153 B.n671 B.n670 585
R154 B.n672 B.n57 585
R155 B.n674 B.n673 585
R156 B.n676 B.n56 585
R157 B.n679 B.n678 585
R158 B.n680 B.n55 585
R159 B.n682 B.n681 585
R160 B.n684 B.n54 585
R161 B.n687 B.n686 585
R162 B.n688 B.n53 585
R163 B.n690 B.n689 585
R164 B.n692 B.n52 585
R165 B.n695 B.n694 585
R166 B.n696 B.n51 585
R167 B.n698 B.n697 585
R168 B.n700 B.n50 585
R169 B.n703 B.n702 585
R170 B.n704 B.n49 585
R171 B.n706 B.n705 585
R172 B.n708 B.n48 585
R173 B.n711 B.n710 585
R174 B.n712 B.n47 585
R175 B.n714 B.n713 585
R176 B.n716 B.n46 585
R177 B.n719 B.n718 585
R178 B.n720 B.n45 585
R179 B.n722 B.n721 585
R180 B.n724 B.n44 585
R181 B.n727 B.n726 585
R182 B.n728 B.n43 585
R183 B.n511 B.n41 585
R184 B.n731 B.n41 585
R185 B.n510 B.n40 585
R186 B.n732 B.n40 585
R187 B.n509 B.n39 585
R188 B.n733 B.n39 585
R189 B.n508 B.n507 585
R190 B.n507 B.n35 585
R191 B.n506 B.n34 585
R192 B.n739 B.n34 585
R193 B.n505 B.n33 585
R194 B.n740 B.n33 585
R195 B.n504 B.n32 585
R196 B.n741 B.n32 585
R197 B.n503 B.n502 585
R198 B.n502 B.n28 585
R199 B.n501 B.n27 585
R200 B.n747 B.n27 585
R201 B.n500 B.n26 585
R202 B.n748 B.n26 585
R203 B.n499 B.n25 585
R204 B.n749 B.n25 585
R205 B.n498 B.n497 585
R206 B.n497 B.n21 585
R207 B.n496 B.n20 585
R208 B.n755 B.n20 585
R209 B.n495 B.n19 585
R210 B.n756 B.n19 585
R211 B.n494 B.n18 585
R212 B.n757 B.n18 585
R213 B.n493 B.n492 585
R214 B.n492 B.n14 585
R215 B.n491 B.n13 585
R216 B.n763 B.n13 585
R217 B.n490 B.n12 585
R218 B.n764 B.n12 585
R219 B.n489 B.n11 585
R220 B.n765 B.n11 585
R221 B.n488 B.n487 585
R222 B.n487 B.t5 585
R223 B.n486 B.n7 585
R224 B.n771 B.n7 585
R225 B.n485 B.n6 585
R226 B.n772 B.n6 585
R227 B.n484 B.n5 585
R228 B.n773 B.n5 585
R229 B.n483 B.n482 585
R230 B.n482 B.n4 585
R231 B.n481 B.n102 585
R232 B.n481 B.n480 585
R233 B.n471 B.n103 585
R234 B.t0 B.n103 585
R235 B.n473 B.n472 585
R236 B.n474 B.n473 585
R237 B.n470 B.n108 585
R238 B.n108 B.n107 585
R239 B.n469 B.n468 585
R240 B.n468 B.n467 585
R241 B.n110 B.n109 585
R242 B.n111 B.n110 585
R243 B.n460 B.n459 585
R244 B.n461 B.n460 585
R245 B.n458 B.n115 585
R246 B.n119 B.n115 585
R247 B.n457 B.n456 585
R248 B.n456 B.n455 585
R249 B.n117 B.n116 585
R250 B.n118 B.n117 585
R251 B.n448 B.n447 585
R252 B.n449 B.n448 585
R253 B.n446 B.n124 585
R254 B.n124 B.n123 585
R255 B.n445 B.n444 585
R256 B.n444 B.n443 585
R257 B.n126 B.n125 585
R258 B.n127 B.n126 585
R259 B.n436 B.n435 585
R260 B.n437 B.n436 585
R261 B.n434 B.n132 585
R262 B.n132 B.n131 585
R263 B.n433 B.n432 585
R264 B.n432 B.n431 585
R265 B.n134 B.n133 585
R266 B.n135 B.n134 585
R267 B.n424 B.n423 585
R268 B.n425 B.n424 585
R269 B.n422 B.n140 585
R270 B.n140 B.n139 585
R271 B.n421 B.n420 585
R272 B.n420 B.n419 585
R273 B.n416 B.n144 585
R274 B.n415 B.n414 585
R275 B.n412 B.n145 585
R276 B.n412 B.n143 585
R277 B.n411 B.n410 585
R278 B.n409 B.n408 585
R279 B.n407 B.n147 585
R280 B.n405 B.n404 585
R281 B.n403 B.n148 585
R282 B.n402 B.n401 585
R283 B.n399 B.n149 585
R284 B.n397 B.n396 585
R285 B.n395 B.n150 585
R286 B.n394 B.n393 585
R287 B.n391 B.n151 585
R288 B.n389 B.n388 585
R289 B.n387 B.n152 585
R290 B.n386 B.n385 585
R291 B.n383 B.n153 585
R292 B.n381 B.n380 585
R293 B.n379 B.n154 585
R294 B.n378 B.n377 585
R295 B.n375 B.n155 585
R296 B.n373 B.n372 585
R297 B.n371 B.n156 585
R298 B.n370 B.n369 585
R299 B.n367 B.n157 585
R300 B.n365 B.n364 585
R301 B.n363 B.n158 585
R302 B.n362 B.n361 585
R303 B.n359 B.n159 585
R304 B.n357 B.n356 585
R305 B.n355 B.n160 585
R306 B.n354 B.n353 585
R307 B.n351 B.n161 585
R308 B.n349 B.n348 585
R309 B.n347 B.n162 585
R310 B.n346 B.n345 585
R311 B.n343 B.n163 585
R312 B.n341 B.n340 585
R313 B.n339 B.n164 585
R314 B.n338 B.n337 585
R315 B.n335 B.n165 585
R316 B.n333 B.n332 585
R317 B.n331 B.n166 585
R318 B.n330 B.n329 585
R319 B.n327 B.n167 585
R320 B.n325 B.n324 585
R321 B.n323 B.n168 585
R322 B.n322 B.n321 585
R323 B.n319 B.n318 585
R324 B.n317 B.n316 585
R325 B.n315 B.n173 585
R326 B.n313 B.n312 585
R327 B.n311 B.n174 585
R328 B.n310 B.n309 585
R329 B.n307 B.n175 585
R330 B.n305 B.n304 585
R331 B.n303 B.n176 585
R332 B.n302 B.n301 585
R333 B.n299 B.n298 585
R334 B.n297 B.n296 585
R335 B.n295 B.n181 585
R336 B.n293 B.n292 585
R337 B.n291 B.n182 585
R338 B.n290 B.n289 585
R339 B.n287 B.n183 585
R340 B.n285 B.n284 585
R341 B.n283 B.n184 585
R342 B.n282 B.n281 585
R343 B.n279 B.n185 585
R344 B.n277 B.n276 585
R345 B.n275 B.n186 585
R346 B.n274 B.n273 585
R347 B.n271 B.n187 585
R348 B.n269 B.n268 585
R349 B.n267 B.n188 585
R350 B.n266 B.n265 585
R351 B.n263 B.n189 585
R352 B.n261 B.n260 585
R353 B.n259 B.n190 585
R354 B.n258 B.n257 585
R355 B.n255 B.n191 585
R356 B.n253 B.n252 585
R357 B.n251 B.n192 585
R358 B.n250 B.n249 585
R359 B.n247 B.n193 585
R360 B.n245 B.n244 585
R361 B.n243 B.n194 585
R362 B.n242 B.n241 585
R363 B.n239 B.n195 585
R364 B.n237 B.n236 585
R365 B.n235 B.n196 585
R366 B.n234 B.n233 585
R367 B.n231 B.n197 585
R368 B.n229 B.n228 585
R369 B.n227 B.n198 585
R370 B.n226 B.n225 585
R371 B.n223 B.n199 585
R372 B.n221 B.n220 585
R373 B.n219 B.n200 585
R374 B.n218 B.n217 585
R375 B.n215 B.n201 585
R376 B.n213 B.n212 585
R377 B.n211 B.n202 585
R378 B.n210 B.n209 585
R379 B.n207 B.n203 585
R380 B.n205 B.n204 585
R381 B.n142 B.n141 585
R382 B.n143 B.n142 585
R383 B.n418 B.n417 585
R384 B.n419 B.n418 585
R385 B.n138 B.n137 585
R386 B.n139 B.n138 585
R387 B.n427 B.n426 585
R388 B.n426 B.n425 585
R389 B.n428 B.n136 585
R390 B.n136 B.n135 585
R391 B.n430 B.n429 585
R392 B.n431 B.n430 585
R393 B.n130 B.n129 585
R394 B.n131 B.n130 585
R395 B.n439 B.n438 585
R396 B.n438 B.n437 585
R397 B.n440 B.n128 585
R398 B.n128 B.n127 585
R399 B.n442 B.n441 585
R400 B.n443 B.n442 585
R401 B.n122 B.n121 585
R402 B.n123 B.n122 585
R403 B.n451 B.n450 585
R404 B.n450 B.n449 585
R405 B.n452 B.n120 585
R406 B.n120 B.n118 585
R407 B.n454 B.n453 585
R408 B.n455 B.n454 585
R409 B.n114 B.n113 585
R410 B.n119 B.n114 585
R411 B.n463 B.n462 585
R412 B.n462 B.n461 585
R413 B.n464 B.n112 585
R414 B.n112 B.n111 585
R415 B.n466 B.n465 585
R416 B.n467 B.n466 585
R417 B.n106 B.n105 585
R418 B.n107 B.n106 585
R419 B.n476 B.n475 585
R420 B.n475 B.n474 585
R421 B.n477 B.n104 585
R422 B.n104 B.t0 585
R423 B.n479 B.n478 585
R424 B.n480 B.n479 585
R425 B.n2 B.n0 585
R426 B.n4 B.n2 585
R427 B.n3 B.n1 585
R428 B.n772 B.n3 585
R429 B.n770 B.n769 585
R430 B.n771 B.n770 585
R431 B.n768 B.n8 585
R432 B.n8 B.t5 585
R433 B.n767 B.n766 585
R434 B.n766 B.n765 585
R435 B.n10 B.n9 585
R436 B.n764 B.n10 585
R437 B.n762 B.n761 585
R438 B.n763 B.n762 585
R439 B.n760 B.n15 585
R440 B.n15 B.n14 585
R441 B.n759 B.n758 585
R442 B.n758 B.n757 585
R443 B.n17 B.n16 585
R444 B.n756 B.n17 585
R445 B.n754 B.n753 585
R446 B.n755 B.n754 585
R447 B.n752 B.n22 585
R448 B.n22 B.n21 585
R449 B.n751 B.n750 585
R450 B.n750 B.n749 585
R451 B.n24 B.n23 585
R452 B.n748 B.n24 585
R453 B.n746 B.n745 585
R454 B.n747 B.n746 585
R455 B.n744 B.n29 585
R456 B.n29 B.n28 585
R457 B.n743 B.n742 585
R458 B.n742 B.n741 585
R459 B.n31 B.n30 585
R460 B.n740 B.n31 585
R461 B.n738 B.n737 585
R462 B.n739 B.n738 585
R463 B.n736 B.n36 585
R464 B.n36 B.n35 585
R465 B.n735 B.n734 585
R466 B.n734 B.n733 585
R467 B.n38 B.n37 585
R468 B.n732 B.n38 585
R469 B.n730 B.n729 585
R470 B.n731 B.n730 585
R471 B.n775 B.n774 585
R472 B.n774 B.n773 585
R473 B.n418 B.n144 473.281
R474 B.n730 B.n43 473.281
R475 B.n420 B.n142 473.281
R476 B.n513 B.n41 473.281
R477 B.n514 B.n42 256.663
R478 B.n516 B.n42 256.663
R479 B.n522 B.n42 256.663
R480 B.n524 B.n42 256.663
R481 B.n530 B.n42 256.663
R482 B.n532 B.n42 256.663
R483 B.n538 B.n42 256.663
R484 B.n540 B.n42 256.663
R485 B.n546 B.n42 256.663
R486 B.n548 B.n42 256.663
R487 B.n554 B.n42 256.663
R488 B.n556 B.n42 256.663
R489 B.n562 B.n42 256.663
R490 B.n564 B.n42 256.663
R491 B.n570 B.n42 256.663
R492 B.n572 B.n42 256.663
R493 B.n578 B.n42 256.663
R494 B.n580 B.n42 256.663
R495 B.n586 B.n42 256.663
R496 B.n588 B.n42 256.663
R497 B.n594 B.n42 256.663
R498 B.n596 B.n42 256.663
R499 B.n602 B.n42 256.663
R500 B.n604 B.n42 256.663
R501 B.n610 B.n42 256.663
R502 B.n612 B.n42 256.663
R503 B.n618 B.n42 256.663
R504 B.n620 B.n42 256.663
R505 B.n626 B.n42 256.663
R506 B.n628 B.n42 256.663
R507 B.n635 B.n42 256.663
R508 B.n637 B.n42 256.663
R509 B.n643 B.n42 256.663
R510 B.n645 B.n42 256.663
R511 B.n651 B.n42 256.663
R512 B.n653 B.n42 256.663
R513 B.n659 B.n42 256.663
R514 B.n661 B.n42 256.663
R515 B.n667 B.n42 256.663
R516 B.n669 B.n42 256.663
R517 B.n675 B.n42 256.663
R518 B.n677 B.n42 256.663
R519 B.n683 B.n42 256.663
R520 B.n685 B.n42 256.663
R521 B.n691 B.n42 256.663
R522 B.n693 B.n42 256.663
R523 B.n699 B.n42 256.663
R524 B.n701 B.n42 256.663
R525 B.n707 B.n42 256.663
R526 B.n709 B.n42 256.663
R527 B.n715 B.n42 256.663
R528 B.n717 B.n42 256.663
R529 B.n723 B.n42 256.663
R530 B.n725 B.n42 256.663
R531 B.n413 B.n143 256.663
R532 B.n146 B.n143 256.663
R533 B.n406 B.n143 256.663
R534 B.n400 B.n143 256.663
R535 B.n398 B.n143 256.663
R536 B.n392 B.n143 256.663
R537 B.n390 B.n143 256.663
R538 B.n384 B.n143 256.663
R539 B.n382 B.n143 256.663
R540 B.n376 B.n143 256.663
R541 B.n374 B.n143 256.663
R542 B.n368 B.n143 256.663
R543 B.n366 B.n143 256.663
R544 B.n360 B.n143 256.663
R545 B.n358 B.n143 256.663
R546 B.n352 B.n143 256.663
R547 B.n350 B.n143 256.663
R548 B.n344 B.n143 256.663
R549 B.n342 B.n143 256.663
R550 B.n336 B.n143 256.663
R551 B.n334 B.n143 256.663
R552 B.n328 B.n143 256.663
R553 B.n326 B.n143 256.663
R554 B.n320 B.n143 256.663
R555 B.n172 B.n143 256.663
R556 B.n314 B.n143 256.663
R557 B.n308 B.n143 256.663
R558 B.n306 B.n143 256.663
R559 B.n300 B.n143 256.663
R560 B.n180 B.n143 256.663
R561 B.n294 B.n143 256.663
R562 B.n288 B.n143 256.663
R563 B.n286 B.n143 256.663
R564 B.n280 B.n143 256.663
R565 B.n278 B.n143 256.663
R566 B.n272 B.n143 256.663
R567 B.n270 B.n143 256.663
R568 B.n264 B.n143 256.663
R569 B.n262 B.n143 256.663
R570 B.n256 B.n143 256.663
R571 B.n254 B.n143 256.663
R572 B.n248 B.n143 256.663
R573 B.n246 B.n143 256.663
R574 B.n240 B.n143 256.663
R575 B.n238 B.n143 256.663
R576 B.n232 B.n143 256.663
R577 B.n230 B.n143 256.663
R578 B.n224 B.n143 256.663
R579 B.n222 B.n143 256.663
R580 B.n216 B.n143 256.663
R581 B.n214 B.n143 256.663
R582 B.n208 B.n143 256.663
R583 B.n206 B.n143 256.663
R584 B.n418 B.n138 163.367
R585 B.n426 B.n138 163.367
R586 B.n426 B.n136 163.367
R587 B.n430 B.n136 163.367
R588 B.n430 B.n130 163.367
R589 B.n438 B.n130 163.367
R590 B.n438 B.n128 163.367
R591 B.n442 B.n128 163.367
R592 B.n442 B.n122 163.367
R593 B.n450 B.n122 163.367
R594 B.n450 B.n120 163.367
R595 B.n454 B.n120 163.367
R596 B.n454 B.n114 163.367
R597 B.n462 B.n114 163.367
R598 B.n462 B.n112 163.367
R599 B.n466 B.n112 163.367
R600 B.n466 B.n106 163.367
R601 B.n475 B.n106 163.367
R602 B.n475 B.n104 163.367
R603 B.n479 B.n104 163.367
R604 B.n479 B.n2 163.367
R605 B.n774 B.n2 163.367
R606 B.n774 B.n3 163.367
R607 B.n770 B.n3 163.367
R608 B.n770 B.n8 163.367
R609 B.n766 B.n8 163.367
R610 B.n766 B.n10 163.367
R611 B.n762 B.n10 163.367
R612 B.n762 B.n15 163.367
R613 B.n758 B.n15 163.367
R614 B.n758 B.n17 163.367
R615 B.n754 B.n17 163.367
R616 B.n754 B.n22 163.367
R617 B.n750 B.n22 163.367
R618 B.n750 B.n24 163.367
R619 B.n746 B.n24 163.367
R620 B.n746 B.n29 163.367
R621 B.n742 B.n29 163.367
R622 B.n742 B.n31 163.367
R623 B.n738 B.n31 163.367
R624 B.n738 B.n36 163.367
R625 B.n734 B.n36 163.367
R626 B.n734 B.n38 163.367
R627 B.n730 B.n38 163.367
R628 B.n414 B.n412 163.367
R629 B.n412 B.n411 163.367
R630 B.n408 B.n407 163.367
R631 B.n405 B.n148 163.367
R632 B.n401 B.n399 163.367
R633 B.n397 B.n150 163.367
R634 B.n393 B.n391 163.367
R635 B.n389 B.n152 163.367
R636 B.n385 B.n383 163.367
R637 B.n381 B.n154 163.367
R638 B.n377 B.n375 163.367
R639 B.n373 B.n156 163.367
R640 B.n369 B.n367 163.367
R641 B.n365 B.n158 163.367
R642 B.n361 B.n359 163.367
R643 B.n357 B.n160 163.367
R644 B.n353 B.n351 163.367
R645 B.n349 B.n162 163.367
R646 B.n345 B.n343 163.367
R647 B.n341 B.n164 163.367
R648 B.n337 B.n335 163.367
R649 B.n333 B.n166 163.367
R650 B.n329 B.n327 163.367
R651 B.n325 B.n168 163.367
R652 B.n321 B.n319 163.367
R653 B.n316 B.n315 163.367
R654 B.n313 B.n174 163.367
R655 B.n309 B.n307 163.367
R656 B.n305 B.n176 163.367
R657 B.n301 B.n299 163.367
R658 B.n296 B.n295 163.367
R659 B.n293 B.n182 163.367
R660 B.n289 B.n287 163.367
R661 B.n285 B.n184 163.367
R662 B.n281 B.n279 163.367
R663 B.n277 B.n186 163.367
R664 B.n273 B.n271 163.367
R665 B.n269 B.n188 163.367
R666 B.n265 B.n263 163.367
R667 B.n261 B.n190 163.367
R668 B.n257 B.n255 163.367
R669 B.n253 B.n192 163.367
R670 B.n249 B.n247 163.367
R671 B.n245 B.n194 163.367
R672 B.n241 B.n239 163.367
R673 B.n237 B.n196 163.367
R674 B.n233 B.n231 163.367
R675 B.n229 B.n198 163.367
R676 B.n225 B.n223 163.367
R677 B.n221 B.n200 163.367
R678 B.n217 B.n215 163.367
R679 B.n213 B.n202 163.367
R680 B.n209 B.n207 163.367
R681 B.n205 B.n142 163.367
R682 B.n420 B.n140 163.367
R683 B.n424 B.n140 163.367
R684 B.n424 B.n134 163.367
R685 B.n432 B.n134 163.367
R686 B.n432 B.n132 163.367
R687 B.n436 B.n132 163.367
R688 B.n436 B.n126 163.367
R689 B.n444 B.n126 163.367
R690 B.n444 B.n124 163.367
R691 B.n448 B.n124 163.367
R692 B.n448 B.n117 163.367
R693 B.n456 B.n117 163.367
R694 B.n456 B.n115 163.367
R695 B.n460 B.n115 163.367
R696 B.n460 B.n110 163.367
R697 B.n468 B.n110 163.367
R698 B.n468 B.n108 163.367
R699 B.n473 B.n108 163.367
R700 B.n473 B.n103 163.367
R701 B.n481 B.n103 163.367
R702 B.n482 B.n481 163.367
R703 B.n482 B.n5 163.367
R704 B.n6 B.n5 163.367
R705 B.n7 B.n6 163.367
R706 B.n487 B.n7 163.367
R707 B.n487 B.n11 163.367
R708 B.n12 B.n11 163.367
R709 B.n13 B.n12 163.367
R710 B.n492 B.n13 163.367
R711 B.n492 B.n18 163.367
R712 B.n19 B.n18 163.367
R713 B.n20 B.n19 163.367
R714 B.n497 B.n20 163.367
R715 B.n497 B.n25 163.367
R716 B.n26 B.n25 163.367
R717 B.n27 B.n26 163.367
R718 B.n502 B.n27 163.367
R719 B.n502 B.n32 163.367
R720 B.n33 B.n32 163.367
R721 B.n34 B.n33 163.367
R722 B.n507 B.n34 163.367
R723 B.n507 B.n39 163.367
R724 B.n40 B.n39 163.367
R725 B.n41 B.n40 163.367
R726 B.n726 B.n724 163.367
R727 B.n722 B.n45 163.367
R728 B.n718 B.n716 163.367
R729 B.n714 B.n47 163.367
R730 B.n710 B.n708 163.367
R731 B.n706 B.n49 163.367
R732 B.n702 B.n700 163.367
R733 B.n698 B.n51 163.367
R734 B.n694 B.n692 163.367
R735 B.n690 B.n53 163.367
R736 B.n686 B.n684 163.367
R737 B.n682 B.n55 163.367
R738 B.n678 B.n676 163.367
R739 B.n674 B.n57 163.367
R740 B.n670 B.n668 163.367
R741 B.n666 B.n59 163.367
R742 B.n662 B.n660 163.367
R743 B.n658 B.n61 163.367
R744 B.n654 B.n652 163.367
R745 B.n650 B.n63 163.367
R746 B.n646 B.n644 163.367
R747 B.n642 B.n65 163.367
R748 B.n638 B.n636 163.367
R749 B.n634 B.n67 163.367
R750 B.n629 B.n627 163.367
R751 B.n625 B.n71 163.367
R752 B.n621 B.n619 163.367
R753 B.n617 B.n73 163.367
R754 B.n613 B.n611 163.367
R755 B.n609 B.n75 163.367
R756 B.n605 B.n603 163.367
R757 B.n601 B.n80 163.367
R758 B.n597 B.n595 163.367
R759 B.n593 B.n82 163.367
R760 B.n589 B.n587 163.367
R761 B.n585 B.n84 163.367
R762 B.n581 B.n579 163.367
R763 B.n577 B.n86 163.367
R764 B.n573 B.n571 163.367
R765 B.n569 B.n88 163.367
R766 B.n565 B.n563 163.367
R767 B.n561 B.n90 163.367
R768 B.n557 B.n555 163.367
R769 B.n553 B.n92 163.367
R770 B.n549 B.n547 163.367
R771 B.n545 B.n94 163.367
R772 B.n541 B.n539 163.367
R773 B.n537 B.n96 163.367
R774 B.n533 B.n531 163.367
R775 B.n529 B.n98 163.367
R776 B.n525 B.n523 163.367
R777 B.n521 B.n100 163.367
R778 B.n517 B.n515 163.367
R779 B.n177 B.t18 90.1998
R780 B.n76 B.t20 90.1998
R781 B.n169 B.t11 90.1811
R782 B.n68 B.t14 90.1811
R783 B.n178 B.t17 71.7756
R784 B.n77 B.t21 71.7756
R785 B.n419 B.n143 71.7578
R786 B.n731 B.n42 71.7578
R787 B.n170 B.t10 71.7568
R788 B.n69 B.t15 71.7568
R789 B.n413 B.n144 71.676
R790 B.n411 B.n146 71.676
R791 B.n407 B.n406 71.676
R792 B.n400 B.n148 71.676
R793 B.n399 B.n398 71.676
R794 B.n392 B.n150 71.676
R795 B.n391 B.n390 71.676
R796 B.n384 B.n152 71.676
R797 B.n383 B.n382 71.676
R798 B.n376 B.n154 71.676
R799 B.n375 B.n374 71.676
R800 B.n368 B.n156 71.676
R801 B.n367 B.n366 71.676
R802 B.n360 B.n158 71.676
R803 B.n359 B.n358 71.676
R804 B.n352 B.n160 71.676
R805 B.n351 B.n350 71.676
R806 B.n344 B.n162 71.676
R807 B.n343 B.n342 71.676
R808 B.n336 B.n164 71.676
R809 B.n335 B.n334 71.676
R810 B.n328 B.n166 71.676
R811 B.n327 B.n326 71.676
R812 B.n320 B.n168 71.676
R813 B.n319 B.n172 71.676
R814 B.n315 B.n314 71.676
R815 B.n308 B.n174 71.676
R816 B.n307 B.n306 71.676
R817 B.n300 B.n176 71.676
R818 B.n299 B.n180 71.676
R819 B.n295 B.n294 71.676
R820 B.n288 B.n182 71.676
R821 B.n287 B.n286 71.676
R822 B.n280 B.n184 71.676
R823 B.n279 B.n278 71.676
R824 B.n272 B.n186 71.676
R825 B.n271 B.n270 71.676
R826 B.n264 B.n188 71.676
R827 B.n263 B.n262 71.676
R828 B.n256 B.n190 71.676
R829 B.n255 B.n254 71.676
R830 B.n248 B.n192 71.676
R831 B.n247 B.n246 71.676
R832 B.n240 B.n194 71.676
R833 B.n239 B.n238 71.676
R834 B.n232 B.n196 71.676
R835 B.n231 B.n230 71.676
R836 B.n224 B.n198 71.676
R837 B.n223 B.n222 71.676
R838 B.n216 B.n200 71.676
R839 B.n215 B.n214 71.676
R840 B.n208 B.n202 71.676
R841 B.n207 B.n206 71.676
R842 B.n725 B.n43 71.676
R843 B.n724 B.n723 71.676
R844 B.n717 B.n45 71.676
R845 B.n716 B.n715 71.676
R846 B.n709 B.n47 71.676
R847 B.n708 B.n707 71.676
R848 B.n701 B.n49 71.676
R849 B.n700 B.n699 71.676
R850 B.n693 B.n51 71.676
R851 B.n692 B.n691 71.676
R852 B.n685 B.n53 71.676
R853 B.n684 B.n683 71.676
R854 B.n677 B.n55 71.676
R855 B.n676 B.n675 71.676
R856 B.n669 B.n57 71.676
R857 B.n668 B.n667 71.676
R858 B.n661 B.n59 71.676
R859 B.n660 B.n659 71.676
R860 B.n653 B.n61 71.676
R861 B.n652 B.n651 71.676
R862 B.n645 B.n63 71.676
R863 B.n644 B.n643 71.676
R864 B.n637 B.n65 71.676
R865 B.n636 B.n635 71.676
R866 B.n628 B.n67 71.676
R867 B.n627 B.n626 71.676
R868 B.n620 B.n71 71.676
R869 B.n619 B.n618 71.676
R870 B.n612 B.n73 71.676
R871 B.n611 B.n610 71.676
R872 B.n604 B.n75 71.676
R873 B.n603 B.n602 71.676
R874 B.n596 B.n80 71.676
R875 B.n595 B.n594 71.676
R876 B.n588 B.n82 71.676
R877 B.n587 B.n586 71.676
R878 B.n580 B.n84 71.676
R879 B.n579 B.n578 71.676
R880 B.n572 B.n86 71.676
R881 B.n571 B.n570 71.676
R882 B.n564 B.n88 71.676
R883 B.n563 B.n562 71.676
R884 B.n556 B.n90 71.676
R885 B.n555 B.n554 71.676
R886 B.n548 B.n92 71.676
R887 B.n547 B.n546 71.676
R888 B.n540 B.n94 71.676
R889 B.n539 B.n538 71.676
R890 B.n532 B.n96 71.676
R891 B.n531 B.n530 71.676
R892 B.n524 B.n98 71.676
R893 B.n523 B.n522 71.676
R894 B.n516 B.n100 71.676
R895 B.n515 B.n514 71.676
R896 B.n514 B.n513 71.676
R897 B.n517 B.n516 71.676
R898 B.n522 B.n521 71.676
R899 B.n525 B.n524 71.676
R900 B.n530 B.n529 71.676
R901 B.n533 B.n532 71.676
R902 B.n538 B.n537 71.676
R903 B.n541 B.n540 71.676
R904 B.n546 B.n545 71.676
R905 B.n549 B.n548 71.676
R906 B.n554 B.n553 71.676
R907 B.n557 B.n556 71.676
R908 B.n562 B.n561 71.676
R909 B.n565 B.n564 71.676
R910 B.n570 B.n569 71.676
R911 B.n573 B.n572 71.676
R912 B.n578 B.n577 71.676
R913 B.n581 B.n580 71.676
R914 B.n586 B.n585 71.676
R915 B.n589 B.n588 71.676
R916 B.n594 B.n593 71.676
R917 B.n597 B.n596 71.676
R918 B.n602 B.n601 71.676
R919 B.n605 B.n604 71.676
R920 B.n610 B.n609 71.676
R921 B.n613 B.n612 71.676
R922 B.n618 B.n617 71.676
R923 B.n621 B.n620 71.676
R924 B.n626 B.n625 71.676
R925 B.n629 B.n628 71.676
R926 B.n635 B.n634 71.676
R927 B.n638 B.n637 71.676
R928 B.n643 B.n642 71.676
R929 B.n646 B.n645 71.676
R930 B.n651 B.n650 71.676
R931 B.n654 B.n653 71.676
R932 B.n659 B.n658 71.676
R933 B.n662 B.n661 71.676
R934 B.n667 B.n666 71.676
R935 B.n670 B.n669 71.676
R936 B.n675 B.n674 71.676
R937 B.n678 B.n677 71.676
R938 B.n683 B.n682 71.676
R939 B.n686 B.n685 71.676
R940 B.n691 B.n690 71.676
R941 B.n694 B.n693 71.676
R942 B.n699 B.n698 71.676
R943 B.n702 B.n701 71.676
R944 B.n707 B.n706 71.676
R945 B.n710 B.n709 71.676
R946 B.n715 B.n714 71.676
R947 B.n718 B.n717 71.676
R948 B.n723 B.n722 71.676
R949 B.n726 B.n725 71.676
R950 B.n414 B.n413 71.676
R951 B.n408 B.n146 71.676
R952 B.n406 B.n405 71.676
R953 B.n401 B.n400 71.676
R954 B.n398 B.n397 71.676
R955 B.n393 B.n392 71.676
R956 B.n390 B.n389 71.676
R957 B.n385 B.n384 71.676
R958 B.n382 B.n381 71.676
R959 B.n377 B.n376 71.676
R960 B.n374 B.n373 71.676
R961 B.n369 B.n368 71.676
R962 B.n366 B.n365 71.676
R963 B.n361 B.n360 71.676
R964 B.n358 B.n357 71.676
R965 B.n353 B.n352 71.676
R966 B.n350 B.n349 71.676
R967 B.n345 B.n344 71.676
R968 B.n342 B.n341 71.676
R969 B.n337 B.n336 71.676
R970 B.n334 B.n333 71.676
R971 B.n329 B.n328 71.676
R972 B.n326 B.n325 71.676
R973 B.n321 B.n320 71.676
R974 B.n316 B.n172 71.676
R975 B.n314 B.n313 71.676
R976 B.n309 B.n308 71.676
R977 B.n306 B.n305 71.676
R978 B.n301 B.n300 71.676
R979 B.n296 B.n180 71.676
R980 B.n294 B.n293 71.676
R981 B.n289 B.n288 71.676
R982 B.n286 B.n285 71.676
R983 B.n281 B.n280 71.676
R984 B.n278 B.n277 71.676
R985 B.n273 B.n272 71.676
R986 B.n270 B.n269 71.676
R987 B.n265 B.n264 71.676
R988 B.n262 B.n261 71.676
R989 B.n257 B.n256 71.676
R990 B.n254 B.n253 71.676
R991 B.n249 B.n248 71.676
R992 B.n246 B.n245 71.676
R993 B.n241 B.n240 71.676
R994 B.n238 B.n237 71.676
R995 B.n233 B.n232 71.676
R996 B.n230 B.n229 71.676
R997 B.n225 B.n224 71.676
R998 B.n222 B.n221 71.676
R999 B.n217 B.n216 71.676
R1000 B.n214 B.n213 71.676
R1001 B.n209 B.n208 71.676
R1002 B.n206 B.n205 71.676
R1003 B.n179 B.n178 59.5399
R1004 B.n171 B.n170 59.5399
R1005 B.n631 B.n69 59.5399
R1006 B.n78 B.n77 59.5399
R1007 B.n419 B.n139 37.826
R1008 B.n425 B.n139 37.826
R1009 B.n425 B.n135 37.826
R1010 B.n431 B.n135 37.826
R1011 B.n437 B.n131 37.826
R1012 B.n437 B.n127 37.826
R1013 B.n443 B.n127 37.826
R1014 B.n443 B.n123 37.826
R1015 B.n449 B.n123 37.826
R1016 B.n455 B.n118 37.826
R1017 B.n455 B.n119 37.826
R1018 B.n461 B.n111 37.826
R1019 B.n467 B.n111 37.826
R1020 B.n474 B.n107 37.826
R1021 B.n474 B.t0 37.826
R1022 B.n480 B.t0 37.826
R1023 B.n480 B.n4 37.826
R1024 B.n773 B.n4 37.826
R1025 B.n773 B.n772 37.826
R1026 B.n772 B.n771 37.826
R1027 B.n771 B.t5 37.826
R1028 B.n765 B.t5 37.826
R1029 B.n765 B.n764 37.826
R1030 B.n763 B.n14 37.826
R1031 B.n757 B.n14 37.826
R1032 B.n756 B.n755 37.826
R1033 B.n755 B.n21 37.826
R1034 B.n749 B.n748 37.826
R1035 B.n748 B.n747 37.826
R1036 B.n747 B.n28 37.826
R1037 B.n741 B.n28 37.826
R1038 B.n741 B.n740 37.826
R1039 B.n739 B.n35 37.826
R1040 B.n733 B.n35 37.826
R1041 B.n733 B.n732 37.826
R1042 B.n732 B.n731 37.826
R1043 B.n729 B.n728 30.7517
R1044 B.n512 B.n511 30.7517
R1045 B.n421 B.n141 30.7517
R1046 B.n417 B.n416 30.7517
R1047 B.t1 B.n107 30.0384
R1048 B.n764 B.t3 30.0384
R1049 B.n431 B.t9 23.3633
R1050 B.n449 B.t6 23.3633
R1051 B.n749 B.t7 23.3633
R1052 B.t13 B.n739 23.3633
R1053 B.n461 B.t4 22.2508
R1054 B.n757 B.t2 22.2508
R1055 B.n178 B.n177 18.4247
R1056 B.n170 B.n169 18.4247
R1057 B.n69 B.n68 18.4247
R1058 B.n77 B.n76 18.4247
R1059 B B.n775 18.0485
R1060 B.n119 B.t4 15.5757
R1061 B.t2 B.n756 15.5757
R1062 B.t9 B.n131 14.4632
R1063 B.t6 B.n118 14.4632
R1064 B.t7 B.n21 14.4632
R1065 B.n740 B.t13 14.4632
R1066 B.n728 B.n727 10.6151
R1067 B.n727 B.n44 10.6151
R1068 B.n721 B.n44 10.6151
R1069 B.n721 B.n720 10.6151
R1070 B.n720 B.n719 10.6151
R1071 B.n719 B.n46 10.6151
R1072 B.n713 B.n46 10.6151
R1073 B.n713 B.n712 10.6151
R1074 B.n712 B.n711 10.6151
R1075 B.n711 B.n48 10.6151
R1076 B.n705 B.n48 10.6151
R1077 B.n705 B.n704 10.6151
R1078 B.n704 B.n703 10.6151
R1079 B.n703 B.n50 10.6151
R1080 B.n697 B.n50 10.6151
R1081 B.n697 B.n696 10.6151
R1082 B.n696 B.n695 10.6151
R1083 B.n695 B.n52 10.6151
R1084 B.n689 B.n52 10.6151
R1085 B.n689 B.n688 10.6151
R1086 B.n688 B.n687 10.6151
R1087 B.n687 B.n54 10.6151
R1088 B.n681 B.n54 10.6151
R1089 B.n681 B.n680 10.6151
R1090 B.n680 B.n679 10.6151
R1091 B.n679 B.n56 10.6151
R1092 B.n673 B.n56 10.6151
R1093 B.n673 B.n672 10.6151
R1094 B.n672 B.n671 10.6151
R1095 B.n671 B.n58 10.6151
R1096 B.n665 B.n58 10.6151
R1097 B.n665 B.n664 10.6151
R1098 B.n664 B.n663 10.6151
R1099 B.n663 B.n60 10.6151
R1100 B.n657 B.n60 10.6151
R1101 B.n657 B.n656 10.6151
R1102 B.n656 B.n655 10.6151
R1103 B.n655 B.n62 10.6151
R1104 B.n649 B.n62 10.6151
R1105 B.n649 B.n648 10.6151
R1106 B.n648 B.n647 10.6151
R1107 B.n647 B.n64 10.6151
R1108 B.n641 B.n64 10.6151
R1109 B.n641 B.n640 10.6151
R1110 B.n640 B.n639 10.6151
R1111 B.n639 B.n66 10.6151
R1112 B.n633 B.n66 10.6151
R1113 B.n633 B.n632 10.6151
R1114 B.n630 B.n70 10.6151
R1115 B.n624 B.n70 10.6151
R1116 B.n624 B.n623 10.6151
R1117 B.n623 B.n622 10.6151
R1118 B.n622 B.n72 10.6151
R1119 B.n616 B.n72 10.6151
R1120 B.n616 B.n615 10.6151
R1121 B.n615 B.n614 10.6151
R1122 B.n614 B.n74 10.6151
R1123 B.n608 B.n607 10.6151
R1124 B.n607 B.n606 10.6151
R1125 B.n606 B.n79 10.6151
R1126 B.n600 B.n79 10.6151
R1127 B.n600 B.n599 10.6151
R1128 B.n599 B.n598 10.6151
R1129 B.n598 B.n81 10.6151
R1130 B.n592 B.n81 10.6151
R1131 B.n592 B.n591 10.6151
R1132 B.n591 B.n590 10.6151
R1133 B.n590 B.n83 10.6151
R1134 B.n584 B.n83 10.6151
R1135 B.n584 B.n583 10.6151
R1136 B.n583 B.n582 10.6151
R1137 B.n582 B.n85 10.6151
R1138 B.n576 B.n85 10.6151
R1139 B.n576 B.n575 10.6151
R1140 B.n575 B.n574 10.6151
R1141 B.n574 B.n87 10.6151
R1142 B.n568 B.n87 10.6151
R1143 B.n568 B.n567 10.6151
R1144 B.n567 B.n566 10.6151
R1145 B.n566 B.n89 10.6151
R1146 B.n560 B.n89 10.6151
R1147 B.n560 B.n559 10.6151
R1148 B.n559 B.n558 10.6151
R1149 B.n558 B.n91 10.6151
R1150 B.n552 B.n91 10.6151
R1151 B.n552 B.n551 10.6151
R1152 B.n551 B.n550 10.6151
R1153 B.n550 B.n93 10.6151
R1154 B.n544 B.n93 10.6151
R1155 B.n544 B.n543 10.6151
R1156 B.n543 B.n542 10.6151
R1157 B.n542 B.n95 10.6151
R1158 B.n536 B.n95 10.6151
R1159 B.n536 B.n535 10.6151
R1160 B.n535 B.n534 10.6151
R1161 B.n534 B.n97 10.6151
R1162 B.n528 B.n97 10.6151
R1163 B.n528 B.n527 10.6151
R1164 B.n527 B.n526 10.6151
R1165 B.n526 B.n99 10.6151
R1166 B.n520 B.n99 10.6151
R1167 B.n520 B.n519 10.6151
R1168 B.n519 B.n518 10.6151
R1169 B.n518 B.n101 10.6151
R1170 B.n512 B.n101 10.6151
R1171 B.n422 B.n421 10.6151
R1172 B.n423 B.n422 10.6151
R1173 B.n423 B.n133 10.6151
R1174 B.n433 B.n133 10.6151
R1175 B.n434 B.n433 10.6151
R1176 B.n435 B.n434 10.6151
R1177 B.n435 B.n125 10.6151
R1178 B.n445 B.n125 10.6151
R1179 B.n446 B.n445 10.6151
R1180 B.n447 B.n446 10.6151
R1181 B.n447 B.n116 10.6151
R1182 B.n457 B.n116 10.6151
R1183 B.n458 B.n457 10.6151
R1184 B.n459 B.n458 10.6151
R1185 B.n459 B.n109 10.6151
R1186 B.n469 B.n109 10.6151
R1187 B.n470 B.n469 10.6151
R1188 B.n472 B.n470 10.6151
R1189 B.n472 B.n471 10.6151
R1190 B.n471 B.n102 10.6151
R1191 B.n483 B.n102 10.6151
R1192 B.n484 B.n483 10.6151
R1193 B.n485 B.n484 10.6151
R1194 B.n486 B.n485 10.6151
R1195 B.n488 B.n486 10.6151
R1196 B.n489 B.n488 10.6151
R1197 B.n490 B.n489 10.6151
R1198 B.n491 B.n490 10.6151
R1199 B.n493 B.n491 10.6151
R1200 B.n494 B.n493 10.6151
R1201 B.n495 B.n494 10.6151
R1202 B.n496 B.n495 10.6151
R1203 B.n498 B.n496 10.6151
R1204 B.n499 B.n498 10.6151
R1205 B.n500 B.n499 10.6151
R1206 B.n501 B.n500 10.6151
R1207 B.n503 B.n501 10.6151
R1208 B.n504 B.n503 10.6151
R1209 B.n505 B.n504 10.6151
R1210 B.n506 B.n505 10.6151
R1211 B.n508 B.n506 10.6151
R1212 B.n509 B.n508 10.6151
R1213 B.n510 B.n509 10.6151
R1214 B.n511 B.n510 10.6151
R1215 B.n416 B.n415 10.6151
R1216 B.n415 B.n145 10.6151
R1217 B.n410 B.n145 10.6151
R1218 B.n410 B.n409 10.6151
R1219 B.n409 B.n147 10.6151
R1220 B.n404 B.n147 10.6151
R1221 B.n404 B.n403 10.6151
R1222 B.n403 B.n402 10.6151
R1223 B.n402 B.n149 10.6151
R1224 B.n396 B.n149 10.6151
R1225 B.n396 B.n395 10.6151
R1226 B.n395 B.n394 10.6151
R1227 B.n394 B.n151 10.6151
R1228 B.n388 B.n151 10.6151
R1229 B.n388 B.n387 10.6151
R1230 B.n387 B.n386 10.6151
R1231 B.n386 B.n153 10.6151
R1232 B.n380 B.n153 10.6151
R1233 B.n380 B.n379 10.6151
R1234 B.n379 B.n378 10.6151
R1235 B.n378 B.n155 10.6151
R1236 B.n372 B.n155 10.6151
R1237 B.n372 B.n371 10.6151
R1238 B.n371 B.n370 10.6151
R1239 B.n370 B.n157 10.6151
R1240 B.n364 B.n157 10.6151
R1241 B.n364 B.n363 10.6151
R1242 B.n363 B.n362 10.6151
R1243 B.n362 B.n159 10.6151
R1244 B.n356 B.n159 10.6151
R1245 B.n356 B.n355 10.6151
R1246 B.n355 B.n354 10.6151
R1247 B.n354 B.n161 10.6151
R1248 B.n348 B.n161 10.6151
R1249 B.n348 B.n347 10.6151
R1250 B.n347 B.n346 10.6151
R1251 B.n346 B.n163 10.6151
R1252 B.n340 B.n163 10.6151
R1253 B.n340 B.n339 10.6151
R1254 B.n339 B.n338 10.6151
R1255 B.n338 B.n165 10.6151
R1256 B.n332 B.n165 10.6151
R1257 B.n332 B.n331 10.6151
R1258 B.n331 B.n330 10.6151
R1259 B.n330 B.n167 10.6151
R1260 B.n324 B.n167 10.6151
R1261 B.n324 B.n323 10.6151
R1262 B.n323 B.n322 10.6151
R1263 B.n318 B.n317 10.6151
R1264 B.n317 B.n173 10.6151
R1265 B.n312 B.n173 10.6151
R1266 B.n312 B.n311 10.6151
R1267 B.n311 B.n310 10.6151
R1268 B.n310 B.n175 10.6151
R1269 B.n304 B.n175 10.6151
R1270 B.n304 B.n303 10.6151
R1271 B.n303 B.n302 10.6151
R1272 B.n298 B.n297 10.6151
R1273 B.n297 B.n181 10.6151
R1274 B.n292 B.n181 10.6151
R1275 B.n292 B.n291 10.6151
R1276 B.n291 B.n290 10.6151
R1277 B.n290 B.n183 10.6151
R1278 B.n284 B.n183 10.6151
R1279 B.n284 B.n283 10.6151
R1280 B.n283 B.n282 10.6151
R1281 B.n282 B.n185 10.6151
R1282 B.n276 B.n185 10.6151
R1283 B.n276 B.n275 10.6151
R1284 B.n275 B.n274 10.6151
R1285 B.n274 B.n187 10.6151
R1286 B.n268 B.n187 10.6151
R1287 B.n268 B.n267 10.6151
R1288 B.n267 B.n266 10.6151
R1289 B.n266 B.n189 10.6151
R1290 B.n260 B.n189 10.6151
R1291 B.n260 B.n259 10.6151
R1292 B.n259 B.n258 10.6151
R1293 B.n258 B.n191 10.6151
R1294 B.n252 B.n191 10.6151
R1295 B.n252 B.n251 10.6151
R1296 B.n251 B.n250 10.6151
R1297 B.n250 B.n193 10.6151
R1298 B.n244 B.n193 10.6151
R1299 B.n244 B.n243 10.6151
R1300 B.n243 B.n242 10.6151
R1301 B.n242 B.n195 10.6151
R1302 B.n236 B.n195 10.6151
R1303 B.n236 B.n235 10.6151
R1304 B.n235 B.n234 10.6151
R1305 B.n234 B.n197 10.6151
R1306 B.n228 B.n197 10.6151
R1307 B.n228 B.n227 10.6151
R1308 B.n227 B.n226 10.6151
R1309 B.n226 B.n199 10.6151
R1310 B.n220 B.n199 10.6151
R1311 B.n220 B.n219 10.6151
R1312 B.n219 B.n218 10.6151
R1313 B.n218 B.n201 10.6151
R1314 B.n212 B.n201 10.6151
R1315 B.n212 B.n211 10.6151
R1316 B.n211 B.n210 10.6151
R1317 B.n210 B.n203 10.6151
R1318 B.n204 B.n203 10.6151
R1319 B.n204 B.n141 10.6151
R1320 B.n417 B.n137 10.6151
R1321 B.n427 B.n137 10.6151
R1322 B.n428 B.n427 10.6151
R1323 B.n429 B.n428 10.6151
R1324 B.n429 B.n129 10.6151
R1325 B.n439 B.n129 10.6151
R1326 B.n440 B.n439 10.6151
R1327 B.n441 B.n440 10.6151
R1328 B.n441 B.n121 10.6151
R1329 B.n451 B.n121 10.6151
R1330 B.n452 B.n451 10.6151
R1331 B.n453 B.n452 10.6151
R1332 B.n453 B.n113 10.6151
R1333 B.n463 B.n113 10.6151
R1334 B.n464 B.n463 10.6151
R1335 B.n465 B.n464 10.6151
R1336 B.n465 B.n105 10.6151
R1337 B.n476 B.n105 10.6151
R1338 B.n477 B.n476 10.6151
R1339 B.n478 B.n477 10.6151
R1340 B.n478 B.n0 10.6151
R1341 B.n769 B.n1 10.6151
R1342 B.n769 B.n768 10.6151
R1343 B.n768 B.n767 10.6151
R1344 B.n767 B.n9 10.6151
R1345 B.n761 B.n9 10.6151
R1346 B.n761 B.n760 10.6151
R1347 B.n760 B.n759 10.6151
R1348 B.n759 B.n16 10.6151
R1349 B.n753 B.n16 10.6151
R1350 B.n753 B.n752 10.6151
R1351 B.n752 B.n751 10.6151
R1352 B.n751 B.n23 10.6151
R1353 B.n745 B.n23 10.6151
R1354 B.n745 B.n744 10.6151
R1355 B.n744 B.n743 10.6151
R1356 B.n743 B.n30 10.6151
R1357 B.n737 B.n30 10.6151
R1358 B.n737 B.n736 10.6151
R1359 B.n736 B.n735 10.6151
R1360 B.n735 B.n37 10.6151
R1361 B.n729 B.n37 10.6151
R1362 B.n632 B.n631 9.36635
R1363 B.n608 B.n78 9.36635
R1364 B.n322 B.n171 9.36635
R1365 B.n298 B.n179 9.36635
R1366 B.n467 B.t1 7.78811
R1367 B.t3 B.n763 7.78811
R1368 B.n775 B.n0 2.81026
R1369 B.n775 B.n1 2.81026
R1370 B.n631 B.n630 1.24928
R1371 B.n78 B.n74 1.24928
R1372 B.n318 B.n171 1.24928
R1373 B.n302 B.n179 1.24928
R1374 VP.n3 VP.t3 653.811
R1375 VP.n1 VP.t6 626.99
R1376 VP.n10 VP.t5 626.99
R1377 VP.n11 VP.t4 626.99
R1378 VP.n12 VP.t1 626.99
R1379 VP.n6 VP.t2 626.99
R1380 VP.n5 VP.t7 626.99
R1381 VP.n4 VP.t0 626.99
R1382 VP.n13 VP.n12 161.3
R1383 VP.n7 VP.n6 161.3
R1384 VP.n8 VP.n1 161.3
R1385 VP.n5 VP.n2 80.6037
R1386 VP.n11 VP.n0 80.6037
R1387 VP.n10 VP.n9 80.6037
R1388 VP.n10 VP.n1 48.2005
R1389 VP.n11 VP.n10 48.2005
R1390 VP.n12 VP.n11 48.2005
R1391 VP.n6 VP.n5 48.2005
R1392 VP.n5 VP.n4 48.2005
R1393 VP.n3 VP.n2 45.2318
R1394 VP.n8 VP.n7 43.5914
R1395 VP.n4 VP.n3 13.3799
R1396 VP.n9 VP.n0 0.380177
R1397 VP.n7 VP.n2 0.285035
R1398 VP.n9 VP.n8 0.285035
R1399 VP.n13 VP.n0 0.285035
R1400 VP VP.n13 0.0516364
R1401 VDD1 VDD1.n0 65.7002
R1402 VDD1.n3 VDD1.n2 65.5865
R1403 VDD1.n3 VDD1.n1 65.5865
R1404 VDD1.n5 VDD1.n4 65.2324
R1405 VDD1.n5 VDD1.n3 40.4836
R1406 VDD1.n4 VDD1.t0 1.36602
R1407 VDD1.n4 VDD1.t5 1.36602
R1408 VDD1.n0 VDD1.t4 1.36602
R1409 VDD1.n0 VDD1.t7 1.36602
R1410 VDD1.n2 VDD1.t3 1.36602
R1411 VDD1.n2 VDD1.t6 1.36602
R1412 VDD1.n1 VDD1.t1 1.36602
R1413 VDD1.n1 VDD1.t2 1.36602
R1414 VDD1 VDD1.n5 0.351793
C0 VDD1 VDD2 0.787055f
C1 VP VDD1 6.32083f
C2 VTAIL VDD1 13.714299f
C3 VP VDD2 0.30935f
C4 VTAIL VDD2 13.7554f
C5 VN VDD1 0.148521f
C6 VTAIL VP 5.80181f
C7 VN VDD2 6.1604f
C8 VN VP 5.69914f
C9 VN VTAIL 5.78771f
C10 VDD2 B 3.610105f
C11 VDD1 B 3.834013f
C12 VTAIL B 10.245727f
C13 VN B 8.62262f
C14 VP B 6.481054f
C15 VDD1.t4 B 0.321274f
C16 VDD1.t7 B 0.321274f
C17 VDD1.n0 B 2.90672f
C18 VDD1.t1 B 0.321274f
C19 VDD1.t2 B 0.321274f
C20 VDD1.n1 B 2.90606f
C21 VDD1.t3 B 0.321274f
C22 VDD1.t6 B 0.321274f
C23 VDD1.n2 B 2.90606f
C24 VDD1.n3 B 2.60272f
C25 VDD1.t0 B 0.321274f
C26 VDD1.t5 B 0.321274f
C27 VDD1.n4 B 2.9042f
C28 VDD1.n5 B 2.78092f
C29 VP.n0 B 0.077176f
C30 VP.t6 B 1.18427f
C31 VP.n1 B 0.461091f
C32 VP.n2 B 0.228197f
C33 VP.t2 B 1.18427f
C34 VP.t7 B 1.18427f
C35 VP.t0 B 1.18427f
C36 VP.t3 B 1.2032f
C37 VP.n3 B 0.443582f
C38 VP.n4 B 0.471606f
C39 VP.n5 B 0.471606f
C40 VP.n6 B 0.461091f
C41 VP.n7 B 2.04874f
C42 VP.n8 B 2.08706f
C43 VP.n9 B 0.077176f
C44 VP.t5 B 1.18427f
C45 VP.n10 B 0.471606f
C46 VP.t4 B 1.18427f
C47 VP.n11 B 0.471606f
C48 VP.t1 B 1.18427f
C49 VP.n12 B 0.461091f
C50 VP.n13 B 0.051401f
C51 VTAIL.t3 B 0.231117f
C52 VTAIL.t10 B 0.231117f
C53 VTAIL.n0 B 2.03516f
C54 VTAIL.n1 B 0.244868f
C55 VTAIL.t5 B 2.59888f
C56 VTAIL.n2 B 0.33822f
C57 VTAIL.t0 B 2.59888f
C58 VTAIL.n3 B 0.33822f
C59 VTAIL.t14 B 0.231117f
C60 VTAIL.t1 B 0.231117f
C61 VTAIL.n4 B 2.03516f
C62 VTAIL.n5 B 0.294313f
C63 VTAIL.t13 B 2.59888f
C64 VTAIL.n6 B 1.44731f
C65 VTAIL.t7 B 2.5989f
C66 VTAIL.n7 B 1.44729f
C67 VTAIL.t4 B 0.231117f
C68 VTAIL.t8 B 0.231117f
C69 VTAIL.n8 B 2.03516f
C70 VTAIL.n9 B 0.29431f
C71 VTAIL.t6 B 2.5989f
C72 VTAIL.n10 B 0.338203f
C73 VTAIL.t15 B 2.5989f
C74 VTAIL.n11 B 0.338203f
C75 VTAIL.t11 B 0.231117f
C76 VTAIL.t2 B 0.231117f
C77 VTAIL.n12 B 2.03516f
C78 VTAIL.n13 B 0.29431f
C79 VTAIL.t12 B 2.59888f
C80 VTAIL.n14 B 1.44731f
C81 VTAIL.t9 B 2.59888f
C82 VTAIL.n15 B 1.44353f
C83 VDD2.t6 B 0.322946f
C84 VDD2.t0 B 0.322946f
C85 VDD2.n0 B 2.92119f
C86 VDD2.t4 B 0.322946f
C87 VDD2.t3 B 0.322946f
C88 VDD2.n1 B 2.92119f
C89 VDD2.n2 B 2.55621f
C90 VDD2.t5 B 0.322946f
C91 VDD2.t1 B 0.322946f
C92 VDD2.n3 B 2.91933f
C93 VDD2.n4 B 2.76191f
C94 VDD2.t2 B 0.322946f
C95 VDD2.t7 B 0.322946f
C96 VDD2.n5 B 2.92116f
C97 VN.n0 B 0.226087f
C98 VN.t5 B 1.19207f
C99 VN.n1 B 0.439481f
C100 VN.t7 B 1.17333f
C101 VN.n2 B 0.467247f
C102 VN.t0 B 1.17333f
C103 VN.n3 B 0.467247f
C104 VN.t1 B 1.17333f
C105 VN.n4 B 0.456829f
C106 VN.n5 B 0.050926f
C107 VN.n6 B 0.226087f
C108 VN.t2 B 1.17333f
C109 VN.t4 B 1.19207f
C110 VN.n7 B 0.439481f
C111 VN.n8 B 0.467247f
C112 VN.t6 B 1.17333f
C113 VN.n9 B 0.467247f
C114 VN.t3 B 1.17333f
C115 VN.n10 B 0.456829f
C116 VN.n11 B 2.05987f
.ends

