* NGSPICE file created from diff_pair_sample_0195.ext - technology: sky130A

.subckt diff_pair_sample_0195 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t8 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=3.83
X1 VDD2.t9 VN.t0 VTAIL.t1 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=3.83
X2 VDD1.t8 VP.t1 VTAIL.t11 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=3.83
X3 VDD1.t7 VP.t2 VTAIL.t9 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X4 VTAIL.t18 VN.t1 VDD2.t8 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X5 B.t11 B.t9 B.t10 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=3.83
X6 VTAIL.t10 VP.t3 VDD1.t6 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X7 VDD2.t7 VN.t2 VTAIL.t19 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X8 VDD1.t5 VP.t4 VTAIL.t15 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=3.83
X9 VTAIL.t0 VN.t3 VDD2.t6 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X10 VTAIL.t14 VP.t5 VDD1.t4 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X11 VDD2.t5 VN.t4 VTAIL.t7 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=3.2208 ps=19.85 w=19.52 l=3.83
X12 VDD2.t4 VN.t5 VTAIL.t6 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=3.83
X13 VTAIL.t12 VP.t6 VDD1.t3 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X14 VTAIL.t13 VP.t7 VDD1.t2 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X15 VDD1.t1 VP.t8 VTAIL.t16 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=3.83
X16 B.t8 B.t6 B.t7 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=3.83
X17 VDD1.t0 VP.t9 VTAIL.t17 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X18 VTAIL.t5 VN.t6 VDD2.t3 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X19 B.t5 B.t3 B.t4 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=3.83
X20 B.t2 B.t0 B.t1 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=7.6128 pd=39.82 as=0 ps=0 w=19.52 l=3.83
X21 VDD2.t2 VN.t7 VTAIL.t2 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=7.6128 ps=39.82 w=19.52 l=3.83
X22 VDD2.t1 VN.t8 VTAIL.t4 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
X23 VTAIL.t3 VN.t9 VDD2.t0 w_n5962_n4872# sky130_fd_pr__pfet_01v8 ad=3.2208 pd=19.85 as=3.2208 ps=19.85 w=19.52 l=3.83
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n31 VP.t0 155.917
R60 VP.n75 VP.t1 122.829
R61 VP.n89 VP.t6 122.829
R62 VP.n102 VP.t9 122.829
R63 VP.n115 VP.t7 122.829
R64 VP.n0 VP.t8 122.829
R65 VP.n18 VP.t4 122.829
R66 VP.n58 VP.t5 122.829
R67 VP.n45 VP.t2 122.829
R68 VP.n32 VP.t3 122.829
R69 VP.n75 VP.n74 86.8027
R70 VP.n130 VP.n0 86.8027
R71 VP.n73 VP.n18 86.8027
R72 VP.n74 VP.n73 65.5677
R73 VP.n96 VP.n95 56.5617
R74 VP.n109 VP.n108 56.5617
R75 VP.n52 VP.n51 56.5617
R76 VP.n39 VP.n38 56.5617
R77 VP.n32 VP.n31 55.106
R78 VP.n83 VP.n82 41.5458
R79 VP.n122 VP.n121 41.5458
R80 VP.n65 VP.n64 41.5458
R81 VP.n82 VP.n81 39.6083
R82 VP.n122 VP.n2 39.6083
R83 VP.n65 VP.n20 39.6083
R84 VP.n77 VP.n76 24.5923
R85 VP.n77 VP.n16 24.5923
R86 VP.n81 VP.n16 24.5923
R87 VP.n83 VP.n14 24.5923
R88 VP.n87 VP.n14 24.5923
R89 VP.n88 VP.n87 24.5923
R90 VP.n90 VP.n12 24.5923
R91 VP.n94 VP.n12 24.5923
R92 VP.n95 VP.n94 24.5923
R93 VP.n96 VP.n10 24.5923
R94 VP.n100 VP.n10 24.5923
R95 VP.n101 VP.n100 24.5923
R96 VP.n103 VP.n8 24.5923
R97 VP.n107 VP.n8 24.5923
R98 VP.n108 VP.n107 24.5923
R99 VP.n109 VP.n6 24.5923
R100 VP.n113 VP.n6 24.5923
R101 VP.n114 VP.n113 24.5923
R102 VP.n116 VP.n4 24.5923
R103 VP.n120 VP.n4 24.5923
R104 VP.n121 VP.n120 24.5923
R105 VP.n126 VP.n2 24.5923
R106 VP.n127 VP.n126 24.5923
R107 VP.n128 VP.n127 24.5923
R108 VP.n69 VP.n20 24.5923
R109 VP.n70 VP.n69 24.5923
R110 VP.n71 VP.n70 24.5923
R111 VP.n52 VP.n24 24.5923
R112 VP.n56 VP.n24 24.5923
R113 VP.n57 VP.n56 24.5923
R114 VP.n59 VP.n22 24.5923
R115 VP.n63 VP.n22 24.5923
R116 VP.n64 VP.n63 24.5923
R117 VP.n39 VP.n28 24.5923
R118 VP.n43 VP.n28 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n46 VP.n26 24.5923
R121 VP.n50 VP.n26 24.5923
R122 VP.n51 VP.n50 24.5923
R123 VP.n33 VP.n30 24.5923
R124 VP.n37 VP.n30 24.5923
R125 VP.n38 VP.n37 24.5923
R126 VP.n90 VP.n89 20.1658
R127 VP.n115 VP.n114 20.1658
R128 VP.n58 VP.n57 20.1658
R129 VP.n33 VP.n32 20.1658
R130 VP.n102 VP.n101 12.2964
R131 VP.n103 VP.n102 12.2964
R132 VP.n45 VP.n44 12.2964
R133 VP.n46 VP.n45 12.2964
R134 VP.n89 VP.n88 4.42703
R135 VP.n116 VP.n115 4.42703
R136 VP.n59 VP.n58 4.42703
R137 VP.n76 VP.n75 3.44336
R138 VP.n128 VP.n0 3.44336
R139 VP.n71 VP.n18 3.44336
R140 VP.n34 VP.n31 2.44068
R141 VP.n73 VP.n72 0.354861
R142 VP.n74 VP.n17 0.354861
R143 VP.n130 VP.n129 0.354861
R144 VP VP.n130 0.267071
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n367 VTAIL.n366 585
R203 VTAIL.n364 VTAIL.n363 585
R204 VTAIL.n373 VTAIL.n372 585
R205 VTAIL.n375 VTAIL.n374 585
R206 VTAIL.n360 VTAIL.n359 585
R207 VTAIL.n381 VTAIL.n380 585
R208 VTAIL.n384 VTAIL.n383 585
R209 VTAIL.n382 VTAIL.n356 585
R210 VTAIL.n389 VTAIL.n355 585
R211 VTAIL.n391 VTAIL.n390 585
R212 VTAIL.n393 VTAIL.n392 585
R213 VTAIL.n352 VTAIL.n351 585
R214 VTAIL.n399 VTAIL.n398 585
R215 VTAIL.n401 VTAIL.n400 585
R216 VTAIL.n348 VTAIL.n347 585
R217 VTAIL.n407 VTAIL.n406 585
R218 VTAIL.n409 VTAIL.n408 585
R219 VTAIL.n344 VTAIL.n343 585
R220 VTAIL.n415 VTAIL.n414 585
R221 VTAIL.n417 VTAIL.n416 585
R222 VTAIL.n340 VTAIL.n339 585
R223 VTAIL.n423 VTAIL.n422 585
R224 VTAIL.n425 VTAIL.n424 585
R225 VTAIL.n336 VTAIL.n335 585
R226 VTAIL.n431 VTAIL.n430 585
R227 VTAIL.n433 VTAIL.n432 585
R228 VTAIL.n37 VTAIL.n36 585
R229 VTAIL.n34 VTAIL.n33 585
R230 VTAIL.n43 VTAIL.n42 585
R231 VTAIL.n45 VTAIL.n44 585
R232 VTAIL.n30 VTAIL.n29 585
R233 VTAIL.n51 VTAIL.n50 585
R234 VTAIL.n54 VTAIL.n53 585
R235 VTAIL.n52 VTAIL.n26 585
R236 VTAIL.n59 VTAIL.n25 585
R237 VTAIL.n61 VTAIL.n60 585
R238 VTAIL.n63 VTAIL.n62 585
R239 VTAIL.n22 VTAIL.n21 585
R240 VTAIL.n69 VTAIL.n68 585
R241 VTAIL.n71 VTAIL.n70 585
R242 VTAIL.n18 VTAIL.n17 585
R243 VTAIL.n77 VTAIL.n76 585
R244 VTAIL.n79 VTAIL.n78 585
R245 VTAIL.n14 VTAIL.n13 585
R246 VTAIL.n85 VTAIL.n84 585
R247 VTAIL.n87 VTAIL.n86 585
R248 VTAIL.n10 VTAIL.n9 585
R249 VTAIL.n93 VTAIL.n92 585
R250 VTAIL.n95 VTAIL.n94 585
R251 VTAIL.n6 VTAIL.n5 585
R252 VTAIL.n101 VTAIL.n100 585
R253 VTAIL.n103 VTAIL.n102 585
R254 VTAIL.n327 VTAIL.n326 585
R255 VTAIL.n325 VTAIL.n324 585
R256 VTAIL.n230 VTAIL.n229 585
R257 VTAIL.n319 VTAIL.n318 585
R258 VTAIL.n317 VTAIL.n316 585
R259 VTAIL.n234 VTAIL.n233 585
R260 VTAIL.n311 VTAIL.n310 585
R261 VTAIL.n309 VTAIL.n308 585
R262 VTAIL.n238 VTAIL.n237 585
R263 VTAIL.n303 VTAIL.n302 585
R264 VTAIL.n301 VTAIL.n300 585
R265 VTAIL.n242 VTAIL.n241 585
R266 VTAIL.n295 VTAIL.n294 585
R267 VTAIL.n293 VTAIL.n292 585
R268 VTAIL.n246 VTAIL.n245 585
R269 VTAIL.n287 VTAIL.n286 585
R270 VTAIL.n285 VTAIL.n284 585
R271 VTAIL.n283 VTAIL.n249 585
R272 VTAIL.n253 VTAIL.n250 585
R273 VTAIL.n278 VTAIL.n277 585
R274 VTAIL.n276 VTAIL.n275 585
R275 VTAIL.n255 VTAIL.n254 585
R276 VTAIL.n270 VTAIL.n269 585
R277 VTAIL.n268 VTAIL.n267 585
R278 VTAIL.n259 VTAIL.n258 585
R279 VTAIL.n262 VTAIL.n261 585
R280 VTAIL.n217 VTAIL.n216 585
R281 VTAIL.n215 VTAIL.n214 585
R282 VTAIL.n120 VTAIL.n119 585
R283 VTAIL.n209 VTAIL.n208 585
R284 VTAIL.n207 VTAIL.n206 585
R285 VTAIL.n124 VTAIL.n123 585
R286 VTAIL.n201 VTAIL.n200 585
R287 VTAIL.n199 VTAIL.n198 585
R288 VTAIL.n128 VTAIL.n127 585
R289 VTAIL.n193 VTAIL.n192 585
R290 VTAIL.n191 VTAIL.n190 585
R291 VTAIL.n132 VTAIL.n131 585
R292 VTAIL.n185 VTAIL.n184 585
R293 VTAIL.n183 VTAIL.n182 585
R294 VTAIL.n136 VTAIL.n135 585
R295 VTAIL.n177 VTAIL.n176 585
R296 VTAIL.n175 VTAIL.n174 585
R297 VTAIL.n173 VTAIL.n139 585
R298 VTAIL.n143 VTAIL.n140 585
R299 VTAIL.n168 VTAIL.n167 585
R300 VTAIL.n166 VTAIL.n165 585
R301 VTAIL.n145 VTAIL.n144 585
R302 VTAIL.n160 VTAIL.n159 585
R303 VTAIL.n158 VTAIL.n157 585
R304 VTAIL.n149 VTAIL.n148 585
R305 VTAIL.n152 VTAIL.n151 585
R306 VTAIL.n432 VTAIL.n332 498.474
R307 VTAIL.n102 VTAIL.n2 498.474
R308 VTAIL.n326 VTAIL.n226 498.474
R309 VTAIL.n216 VTAIL.n116 498.474
R310 VTAIL.t2 VTAIL.n365 329.036
R311 VTAIL.t16 VTAIL.n35 329.036
R312 VTAIL.t15 VTAIL.n260 329.036
R313 VTAIL.t6 VTAIL.n150 329.036
R314 VTAIL.n366 VTAIL.n363 171.744
R315 VTAIL.n373 VTAIL.n363 171.744
R316 VTAIL.n374 VTAIL.n373 171.744
R317 VTAIL.n374 VTAIL.n359 171.744
R318 VTAIL.n381 VTAIL.n359 171.744
R319 VTAIL.n383 VTAIL.n381 171.744
R320 VTAIL.n383 VTAIL.n382 171.744
R321 VTAIL.n382 VTAIL.n355 171.744
R322 VTAIL.n391 VTAIL.n355 171.744
R323 VTAIL.n392 VTAIL.n391 171.744
R324 VTAIL.n392 VTAIL.n351 171.744
R325 VTAIL.n399 VTAIL.n351 171.744
R326 VTAIL.n400 VTAIL.n399 171.744
R327 VTAIL.n400 VTAIL.n347 171.744
R328 VTAIL.n407 VTAIL.n347 171.744
R329 VTAIL.n408 VTAIL.n407 171.744
R330 VTAIL.n408 VTAIL.n343 171.744
R331 VTAIL.n415 VTAIL.n343 171.744
R332 VTAIL.n416 VTAIL.n415 171.744
R333 VTAIL.n416 VTAIL.n339 171.744
R334 VTAIL.n423 VTAIL.n339 171.744
R335 VTAIL.n424 VTAIL.n423 171.744
R336 VTAIL.n424 VTAIL.n335 171.744
R337 VTAIL.n431 VTAIL.n335 171.744
R338 VTAIL.n432 VTAIL.n431 171.744
R339 VTAIL.n36 VTAIL.n33 171.744
R340 VTAIL.n43 VTAIL.n33 171.744
R341 VTAIL.n44 VTAIL.n43 171.744
R342 VTAIL.n44 VTAIL.n29 171.744
R343 VTAIL.n51 VTAIL.n29 171.744
R344 VTAIL.n53 VTAIL.n51 171.744
R345 VTAIL.n53 VTAIL.n52 171.744
R346 VTAIL.n52 VTAIL.n25 171.744
R347 VTAIL.n61 VTAIL.n25 171.744
R348 VTAIL.n62 VTAIL.n61 171.744
R349 VTAIL.n62 VTAIL.n21 171.744
R350 VTAIL.n69 VTAIL.n21 171.744
R351 VTAIL.n70 VTAIL.n69 171.744
R352 VTAIL.n70 VTAIL.n17 171.744
R353 VTAIL.n77 VTAIL.n17 171.744
R354 VTAIL.n78 VTAIL.n77 171.744
R355 VTAIL.n78 VTAIL.n13 171.744
R356 VTAIL.n85 VTAIL.n13 171.744
R357 VTAIL.n86 VTAIL.n85 171.744
R358 VTAIL.n86 VTAIL.n9 171.744
R359 VTAIL.n93 VTAIL.n9 171.744
R360 VTAIL.n94 VTAIL.n93 171.744
R361 VTAIL.n94 VTAIL.n5 171.744
R362 VTAIL.n101 VTAIL.n5 171.744
R363 VTAIL.n102 VTAIL.n101 171.744
R364 VTAIL.n326 VTAIL.n325 171.744
R365 VTAIL.n325 VTAIL.n229 171.744
R366 VTAIL.n318 VTAIL.n229 171.744
R367 VTAIL.n318 VTAIL.n317 171.744
R368 VTAIL.n317 VTAIL.n233 171.744
R369 VTAIL.n310 VTAIL.n233 171.744
R370 VTAIL.n310 VTAIL.n309 171.744
R371 VTAIL.n309 VTAIL.n237 171.744
R372 VTAIL.n302 VTAIL.n237 171.744
R373 VTAIL.n302 VTAIL.n301 171.744
R374 VTAIL.n301 VTAIL.n241 171.744
R375 VTAIL.n294 VTAIL.n241 171.744
R376 VTAIL.n294 VTAIL.n293 171.744
R377 VTAIL.n293 VTAIL.n245 171.744
R378 VTAIL.n286 VTAIL.n245 171.744
R379 VTAIL.n286 VTAIL.n285 171.744
R380 VTAIL.n285 VTAIL.n249 171.744
R381 VTAIL.n253 VTAIL.n249 171.744
R382 VTAIL.n277 VTAIL.n253 171.744
R383 VTAIL.n277 VTAIL.n276 171.744
R384 VTAIL.n276 VTAIL.n254 171.744
R385 VTAIL.n269 VTAIL.n254 171.744
R386 VTAIL.n269 VTAIL.n268 171.744
R387 VTAIL.n268 VTAIL.n258 171.744
R388 VTAIL.n261 VTAIL.n258 171.744
R389 VTAIL.n216 VTAIL.n215 171.744
R390 VTAIL.n215 VTAIL.n119 171.744
R391 VTAIL.n208 VTAIL.n119 171.744
R392 VTAIL.n208 VTAIL.n207 171.744
R393 VTAIL.n207 VTAIL.n123 171.744
R394 VTAIL.n200 VTAIL.n123 171.744
R395 VTAIL.n200 VTAIL.n199 171.744
R396 VTAIL.n199 VTAIL.n127 171.744
R397 VTAIL.n192 VTAIL.n127 171.744
R398 VTAIL.n192 VTAIL.n191 171.744
R399 VTAIL.n191 VTAIL.n131 171.744
R400 VTAIL.n184 VTAIL.n131 171.744
R401 VTAIL.n184 VTAIL.n183 171.744
R402 VTAIL.n183 VTAIL.n135 171.744
R403 VTAIL.n176 VTAIL.n135 171.744
R404 VTAIL.n176 VTAIL.n175 171.744
R405 VTAIL.n175 VTAIL.n139 171.744
R406 VTAIL.n143 VTAIL.n139 171.744
R407 VTAIL.n167 VTAIL.n143 171.744
R408 VTAIL.n167 VTAIL.n166 171.744
R409 VTAIL.n166 VTAIL.n144 171.744
R410 VTAIL.n159 VTAIL.n144 171.744
R411 VTAIL.n159 VTAIL.n158 171.744
R412 VTAIL.n158 VTAIL.n148 171.744
R413 VTAIL.n151 VTAIL.n148 171.744
R414 VTAIL.n366 VTAIL.t2 85.8723
R415 VTAIL.n36 VTAIL.t16 85.8723
R416 VTAIL.n261 VTAIL.t15 85.8723
R417 VTAIL.n151 VTAIL.t6 85.8723
R418 VTAIL.n225 VTAIL.n224 55.0433
R419 VTAIL.n223 VTAIL.n222 55.0433
R420 VTAIL.n115 VTAIL.n114 55.0433
R421 VTAIL.n113 VTAIL.n112 55.0433
R422 VTAIL.n439 VTAIL.n438 55.0431
R423 VTAIL.n1 VTAIL.n0 55.0431
R424 VTAIL.n109 VTAIL.n108 55.0431
R425 VTAIL.n111 VTAIL.n110 55.0431
R426 VTAIL.n113 VTAIL.n111 36.3669
R427 VTAIL.n437 VTAIL.n436 36.0641
R428 VTAIL.n107 VTAIL.n106 36.0641
R429 VTAIL.n331 VTAIL.n330 36.0641
R430 VTAIL.n221 VTAIL.n220 36.0641
R431 VTAIL.n437 VTAIL.n331 32.7807
R432 VTAIL.n390 VTAIL.n389 13.1884
R433 VTAIL.n60 VTAIL.n59 13.1884
R434 VTAIL.n284 VTAIL.n283 13.1884
R435 VTAIL.n174 VTAIL.n173 13.1884
R436 VTAIL.n388 VTAIL.n356 12.8005
R437 VTAIL.n393 VTAIL.n354 12.8005
R438 VTAIL.n434 VTAIL.n433 12.8005
R439 VTAIL.n58 VTAIL.n26 12.8005
R440 VTAIL.n63 VTAIL.n24 12.8005
R441 VTAIL.n104 VTAIL.n103 12.8005
R442 VTAIL.n328 VTAIL.n327 12.8005
R443 VTAIL.n287 VTAIL.n248 12.8005
R444 VTAIL.n282 VTAIL.n250 12.8005
R445 VTAIL.n218 VTAIL.n217 12.8005
R446 VTAIL.n177 VTAIL.n138 12.8005
R447 VTAIL.n172 VTAIL.n140 12.8005
R448 VTAIL.n385 VTAIL.n384 12.0247
R449 VTAIL.n394 VTAIL.n352 12.0247
R450 VTAIL.n430 VTAIL.n334 12.0247
R451 VTAIL.n55 VTAIL.n54 12.0247
R452 VTAIL.n64 VTAIL.n22 12.0247
R453 VTAIL.n100 VTAIL.n4 12.0247
R454 VTAIL.n324 VTAIL.n228 12.0247
R455 VTAIL.n288 VTAIL.n246 12.0247
R456 VTAIL.n279 VTAIL.n278 12.0247
R457 VTAIL.n214 VTAIL.n118 12.0247
R458 VTAIL.n178 VTAIL.n136 12.0247
R459 VTAIL.n169 VTAIL.n168 12.0247
R460 VTAIL.n380 VTAIL.n358 11.249
R461 VTAIL.n398 VTAIL.n397 11.249
R462 VTAIL.n429 VTAIL.n336 11.249
R463 VTAIL.n50 VTAIL.n28 11.249
R464 VTAIL.n68 VTAIL.n67 11.249
R465 VTAIL.n99 VTAIL.n6 11.249
R466 VTAIL.n323 VTAIL.n230 11.249
R467 VTAIL.n292 VTAIL.n291 11.249
R468 VTAIL.n275 VTAIL.n252 11.249
R469 VTAIL.n213 VTAIL.n120 11.249
R470 VTAIL.n182 VTAIL.n181 11.249
R471 VTAIL.n165 VTAIL.n142 11.249
R472 VTAIL.n367 VTAIL.n365 10.7239
R473 VTAIL.n37 VTAIL.n35 10.7239
R474 VTAIL.n262 VTAIL.n260 10.7239
R475 VTAIL.n152 VTAIL.n150 10.7239
R476 VTAIL.n379 VTAIL.n360 10.4732
R477 VTAIL.n401 VTAIL.n350 10.4732
R478 VTAIL.n426 VTAIL.n425 10.4732
R479 VTAIL.n49 VTAIL.n30 10.4732
R480 VTAIL.n71 VTAIL.n20 10.4732
R481 VTAIL.n96 VTAIL.n95 10.4732
R482 VTAIL.n320 VTAIL.n319 10.4732
R483 VTAIL.n295 VTAIL.n244 10.4732
R484 VTAIL.n274 VTAIL.n255 10.4732
R485 VTAIL.n210 VTAIL.n209 10.4732
R486 VTAIL.n185 VTAIL.n134 10.4732
R487 VTAIL.n164 VTAIL.n145 10.4732
R488 VTAIL.n376 VTAIL.n375 9.69747
R489 VTAIL.n402 VTAIL.n348 9.69747
R490 VTAIL.n422 VTAIL.n338 9.69747
R491 VTAIL.n46 VTAIL.n45 9.69747
R492 VTAIL.n72 VTAIL.n18 9.69747
R493 VTAIL.n92 VTAIL.n8 9.69747
R494 VTAIL.n316 VTAIL.n232 9.69747
R495 VTAIL.n296 VTAIL.n242 9.69747
R496 VTAIL.n271 VTAIL.n270 9.69747
R497 VTAIL.n206 VTAIL.n122 9.69747
R498 VTAIL.n186 VTAIL.n132 9.69747
R499 VTAIL.n161 VTAIL.n160 9.69747
R500 VTAIL.n436 VTAIL.n435 9.45567
R501 VTAIL.n106 VTAIL.n105 9.45567
R502 VTAIL.n330 VTAIL.n329 9.45567
R503 VTAIL.n220 VTAIL.n219 9.45567
R504 VTAIL.n411 VTAIL.n410 9.3005
R505 VTAIL.n346 VTAIL.n345 9.3005
R506 VTAIL.n405 VTAIL.n404 9.3005
R507 VTAIL.n403 VTAIL.n402 9.3005
R508 VTAIL.n350 VTAIL.n349 9.3005
R509 VTAIL.n397 VTAIL.n396 9.3005
R510 VTAIL.n395 VTAIL.n394 9.3005
R511 VTAIL.n354 VTAIL.n353 9.3005
R512 VTAIL.n369 VTAIL.n368 9.3005
R513 VTAIL.n371 VTAIL.n370 9.3005
R514 VTAIL.n362 VTAIL.n361 9.3005
R515 VTAIL.n377 VTAIL.n376 9.3005
R516 VTAIL.n379 VTAIL.n378 9.3005
R517 VTAIL.n358 VTAIL.n357 9.3005
R518 VTAIL.n386 VTAIL.n385 9.3005
R519 VTAIL.n388 VTAIL.n387 9.3005
R520 VTAIL.n413 VTAIL.n412 9.3005
R521 VTAIL.n342 VTAIL.n341 9.3005
R522 VTAIL.n419 VTAIL.n418 9.3005
R523 VTAIL.n421 VTAIL.n420 9.3005
R524 VTAIL.n338 VTAIL.n337 9.3005
R525 VTAIL.n427 VTAIL.n426 9.3005
R526 VTAIL.n429 VTAIL.n428 9.3005
R527 VTAIL.n334 VTAIL.n333 9.3005
R528 VTAIL.n435 VTAIL.n434 9.3005
R529 VTAIL.n81 VTAIL.n80 9.3005
R530 VTAIL.n16 VTAIL.n15 9.3005
R531 VTAIL.n75 VTAIL.n74 9.3005
R532 VTAIL.n73 VTAIL.n72 9.3005
R533 VTAIL.n20 VTAIL.n19 9.3005
R534 VTAIL.n67 VTAIL.n66 9.3005
R535 VTAIL.n65 VTAIL.n64 9.3005
R536 VTAIL.n24 VTAIL.n23 9.3005
R537 VTAIL.n39 VTAIL.n38 9.3005
R538 VTAIL.n41 VTAIL.n40 9.3005
R539 VTAIL.n32 VTAIL.n31 9.3005
R540 VTAIL.n47 VTAIL.n46 9.3005
R541 VTAIL.n49 VTAIL.n48 9.3005
R542 VTAIL.n28 VTAIL.n27 9.3005
R543 VTAIL.n56 VTAIL.n55 9.3005
R544 VTAIL.n58 VTAIL.n57 9.3005
R545 VTAIL.n83 VTAIL.n82 9.3005
R546 VTAIL.n12 VTAIL.n11 9.3005
R547 VTAIL.n89 VTAIL.n88 9.3005
R548 VTAIL.n91 VTAIL.n90 9.3005
R549 VTAIL.n8 VTAIL.n7 9.3005
R550 VTAIL.n97 VTAIL.n96 9.3005
R551 VTAIL.n99 VTAIL.n98 9.3005
R552 VTAIL.n4 VTAIL.n3 9.3005
R553 VTAIL.n105 VTAIL.n104 9.3005
R554 VTAIL.n264 VTAIL.n263 9.3005
R555 VTAIL.n266 VTAIL.n265 9.3005
R556 VTAIL.n257 VTAIL.n256 9.3005
R557 VTAIL.n272 VTAIL.n271 9.3005
R558 VTAIL.n274 VTAIL.n273 9.3005
R559 VTAIL.n252 VTAIL.n251 9.3005
R560 VTAIL.n280 VTAIL.n279 9.3005
R561 VTAIL.n282 VTAIL.n281 9.3005
R562 VTAIL.n236 VTAIL.n235 9.3005
R563 VTAIL.n313 VTAIL.n312 9.3005
R564 VTAIL.n315 VTAIL.n314 9.3005
R565 VTAIL.n232 VTAIL.n231 9.3005
R566 VTAIL.n321 VTAIL.n320 9.3005
R567 VTAIL.n323 VTAIL.n322 9.3005
R568 VTAIL.n228 VTAIL.n227 9.3005
R569 VTAIL.n329 VTAIL.n328 9.3005
R570 VTAIL.n307 VTAIL.n306 9.3005
R571 VTAIL.n305 VTAIL.n304 9.3005
R572 VTAIL.n240 VTAIL.n239 9.3005
R573 VTAIL.n299 VTAIL.n298 9.3005
R574 VTAIL.n297 VTAIL.n296 9.3005
R575 VTAIL.n244 VTAIL.n243 9.3005
R576 VTAIL.n291 VTAIL.n290 9.3005
R577 VTAIL.n289 VTAIL.n288 9.3005
R578 VTAIL.n248 VTAIL.n247 9.3005
R579 VTAIL.n154 VTAIL.n153 9.3005
R580 VTAIL.n156 VTAIL.n155 9.3005
R581 VTAIL.n147 VTAIL.n146 9.3005
R582 VTAIL.n162 VTAIL.n161 9.3005
R583 VTAIL.n164 VTAIL.n163 9.3005
R584 VTAIL.n142 VTAIL.n141 9.3005
R585 VTAIL.n170 VTAIL.n169 9.3005
R586 VTAIL.n172 VTAIL.n171 9.3005
R587 VTAIL.n126 VTAIL.n125 9.3005
R588 VTAIL.n203 VTAIL.n202 9.3005
R589 VTAIL.n205 VTAIL.n204 9.3005
R590 VTAIL.n122 VTAIL.n121 9.3005
R591 VTAIL.n211 VTAIL.n210 9.3005
R592 VTAIL.n213 VTAIL.n212 9.3005
R593 VTAIL.n118 VTAIL.n117 9.3005
R594 VTAIL.n219 VTAIL.n218 9.3005
R595 VTAIL.n197 VTAIL.n196 9.3005
R596 VTAIL.n195 VTAIL.n194 9.3005
R597 VTAIL.n130 VTAIL.n129 9.3005
R598 VTAIL.n189 VTAIL.n188 9.3005
R599 VTAIL.n187 VTAIL.n186 9.3005
R600 VTAIL.n134 VTAIL.n133 9.3005
R601 VTAIL.n181 VTAIL.n180 9.3005
R602 VTAIL.n179 VTAIL.n178 9.3005
R603 VTAIL.n138 VTAIL.n137 9.3005
R604 VTAIL.n372 VTAIL.n362 8.92171
R605 VTAIL.n406 VTAIL.n405 8.92171
R606 VTAIL.n421 VTAIL.n340 8.92171
R607 VTAIL.n42 VTAIL.n32 8.92171
R608 VTAIL.n76 VTAIL.n75 8.92171
R609 VTAIL.n91 VTAIL.n10 8.92171
R610 VTAIL.n315 VTAIL.n234 8.92171
R611 VTAIL.n300 VTAIL.n299 8.92171
R612 VTAIL.n267 VTAIL.n257 8.92171
R613 VTAIL.n205 VTAIL.n124 8.92171
R614 VTAIL.n190 VTAIL.n189 8.92171
R615 VTAIL.n157 VTAIL.n147 8.92171
R616 VTAIL.n371 VTAIL.n364 8.14595
R617 VTAIL.n409 VTAIL.n346 8.14595
R618 VTAIL.n418 VTAIL.n417 8.14595
R619 VTAIL.n41 VTAIL.n34 8.14595
R620 VTAIL.n79 VTAIL.n16 8.14595
R621 VTAIL.n88 VTAIL.n87 8.14595
R622 VTAIL.n312 VTAIL.n311 8.14595
R623 VTAIL.n303 VTAIL.n240 8.14595
R624 VTAIL.n266 VTAIL.n259 8.14595
R625 VTAIL.n202 VTAIL.n201 8.14595
R626 VTAIL.n193 VTAIL.n130 8.14595
R627 VTAIL.n156 VTAIL.n149 8.14595
R628 VTAIL.n436 VTAIL.n332 7.75445
R629 VTAIL.n106 VTAIL.n2 7.75445
R630 VTAIL.n330 VTAIL.n226 7.75445
R631 VTAIL.n220 VTAIL.n116 7.75445
R632 VTAIL.n368 VTAIL.n367 7.3702
R633 VTAIL.n410 VTAIL.n344 7.3702
R634 VTAIL.n414 VTAIL.n342 7.3702
R635 VTAIL.n38 VTAIL.n37 7.3702
R636 VTAIL.n80 VTAIL.n14 7.3702
R637 VTAIL.n84 VTAIL.n12 7.3702
R638 VTAIL.n308 VTAIL.n236 7.3702
R639 VTAIL.n304 VTAIL.n238 7.3702
R640 VTAIL.n263 VTAIL.n262 7.3702
R641 VTAIL.n198 VTAIL.n126 7.3702
R642 VTAIL.n194 VTAIL.n128 7.3702
R643 VTAIL.n153 VTAIL.n152 7.3702
R644 VTAIL.n413 VTAIL.n344 6.59444
R645 VTAIL.n414 VTAIL.n413 6.59444
R646 VTAIL.n83 VTAIL.n14 6.59444
R647 VTAIL.n84 VTAIL.n83 6.59444
R648 VTAIL.n308 VTAIL.n307 6.59444
R649 VTAIL.n307 VTAIL.n238 6.59444
R650 VTAIL.n198 VTAIL.n197 6.59444
R651 VTAIL.n197 VTAIL.n128 6.59444
R652 VTAIL.n434 VTAIL.n332 6.08283
R653 VTAIL.n104 VTAIL.n2 6.08283
R654 VTAIL.n328 VTAIL.n226 6.08283
R655 VTAIL.n218 VTAIL.n116 6.08283
R656 VTAIL.n368 VTAIL.n364 5.81868
R657 VTAIL.n410 VTAIL.n409 5.81868
R658 VTAIL.n417 VTAIL.n342 5.81868
R659 VTAIL.n38 VTAIL.n34 5.81868
R660 VTAIL.n80 VTAIL.n79 5.81868
R661 VTAIL.n87 VTAIL.n12 5.81868
R662 VTAIL.n311 VTAIL.n236 5.81868
R663 VTAIL.n304 VTAIL.n303 5.81868
R664 VTAIL.n263 VTAIL.n259 5.81868
R665 VTAIL.n201 VTAIL.n126 5.81868
R666 VTAIL.n194 VTAIL.n193 5.81868
R667 VTAIL.n153 VTAIL.n149 5.81868
R668 VTAIL.n372 VTAIL.n371 5.04292
R669 VTAIL.n406 VTAIL.n346 5.04292
R670 VTAIL.n418 VTAIL.n340 5.04292
R671 VTAIL.n42 VTAIL.n41 5.04292
R672 VTAIL.n76 VTAIL.n16 5.04292
R673 VTAIL.n88 VTAIL.n10 5.04292
R674 VTAIL.n312 VTAIL.n234 5.04292
R675 VTAIL.n300 VTAIL.n240 5.04292
R676 VTAIL.n267 VTAIL.n266 5.04292
R677 VTAIL.n202 VTAIL.n124 5.04292
R678 VTAIL.n190 VTAIL.n130 5.04292
R679 VTAIL.n157 VTAIL.n156 5.04292
R680 VTAIL.n375 VTAIL.n362 4.26717
R681 VTAIL.n405 VTAIL.n348 4.26717
R682 VTAIL.n422 VTAIL.n421 4.26717
R683 VTAIL.n45 VTAIL.n32 4.26717
R684 VTAIL.n75 VTAIL.n18 4.26717
R685 VTAIL.n92 VTAIL.n91 4.26717
R686 VTAIL.n316 VTAIL.n315 4.26717
R687 VTAIL.n299 VTAIL.n242 4.26717
R688 VTAIL.n270 VTAIL.n257 4.26717
R689 VTAIL.n206 VTAIL.n205 4.26717
R690 VTAIL.n189 VTAIL.n132 4.26717
R691 VTAIL.n160 VTAIL.n147 4.26717
R692 VTAIL.n115 VTAIL.n113 3.58671
R693 VTAIL.n221 VTAIL.n115 3.58671
R694 VTAIL.n225 VTAIL.n223 3.58671
R695 VTAIL.n331 VTAIL.n225 3.58671
R696 VTAIL.n111 VTAIL.n109 3.58671
R697 VTAIL.n109 VTAIL.n107 3.58671
R698 VTAIL.n439 VTAIL.n437 3.58671
R699 VTAIL.n376 VTAIL.n360 3.49141
R700 VTAIL.n402 VTAIL.n401 3.49141
R701 VTAIL.n425 VTAIL.n338 3.49141
R702 VTAIL.n46 VTAIL.n30 3.49141
R703 VTAIL.n72 VTAIL.n71 3.49141
R704 VTAIL.n95 VTAIL.n8 3.49141
R705 VTAIL.n319 VTAIL.n232 3.49141
R706 VTAIL.n296 VTAIL.n295 3.49141
R707 VTAIL.n271 VTAIL.n255 3.49141
R708 VTAIL.n209 VTAIL.n122 3.49141
R709 VTAIL.n186 VTAIL.n185 3.49141
R710 VTAIL.n161 VTAIL.n145 3.49141
R711 VTAIL VTAIL.n1 2.74834
R712 VTAIL.n380 VTAIL.n379 2.71565
R713 VTAIL.n398 VTAIL.n350 2.71565
R714 VTAIL.n426 VTAIL.n336 2.71565
R715 VTAIL.n50 VTAIL.n49 2.71565
R716 VTAIL.n68 VTAIL.n20 2.71565
R717 VTAIL.n96 VTAIL.n6 2.71565
R718 VTAIL.n320 VTAIL.n230 2.71565
R719 VTAIL.n292 VTAIL.n244 2.71565
R720 VTAIL.n275 VTAIL.n274 2.71565
R721 VTAIL.n210 VTAIL.n120 2.71565
R722 VTAIL.n182 VTAIL.n134 2.71565
R723 VTAIL.n165 VTAIL.n164 2.71565
R724 VTAIL.n264 VTAIL.n260 2.41282
R725 VTAIL.n154 VTAIL.n150 2.41282
R726 VTAIL.n369 VTAIL.n365 2.41282
R727 VTAIL.n39 VTAIL.n35 2.41282
R728 VTAIL.n223 VTAIL.n221 2.26343
R729 VTAIL.n107 VTAIL.n1 2.26343
R730 VTAIL.n384 VTAIL.n358 1.93989
R731 VTAIL.n397 VTAIL.n352 1.93989
R732 VTAIL.n430 VTAIL.n429 1.93989
R733 VTAIL.n54 VTAIL.n28 1.93989
R734 VTAIL.n67 VTAIL.n22 1.93989
R735 VTAIL.n100 VTAIL.n99 1.93989
R736 VTAIL.n324 VTAIL.n323 1.93989
R737 VTAIL.n291 VTAIL.n246 1.93989
R738 VTAIL.n278 VTAIL.n252 1.93989
R739 VTAIL.n214 VTAIL.n213 1.93989
R740 VTAIL.n181 VTAIL.n136 1.93989
R741 VTAIL.n168 VTAIL.n142 1.93989
R742 VTAIL.n438 VTAIL.t4 1.66572
R743 VTAIL.n438 VTAIL.t3 1.66572
R744 VTAIL.n0 VTAIL.t7 1.66572
R745 VTAIL.n0 VTAIL.t0 1.66572
R746 VTAIL.n108 VTAIL.t17 1.66572
R747 VTAIL.n108 VTAIL.t13 1.66572
R748 VTAIL.n110 VTAIL.t11 1.66572
R749 VTAIL.n110 VTAIL.t12 1.66572
R750 VTAIL.n224 VTAIL.t9 1.66572
R751 VTAIL.n224 VTAIL.t14 1.66572
R752 VTAIL.n222 VTAIL.t8 1.66572
R753 VTAIL.n222 VTAIL.t10 1.66572
R754 VTAIL.n114 VTAIL.t19 1.66572
R755 VTAIL.n114 VTAIL.t5 1.66572
R756 VTAIL.n112 VTAIL.t1 1.66572
R757 VTAIL.n112 VTAIL.t18 1.66572
R758 VTAIL.n385 VTAIL.n356 1.16414
R759 VTAIL.n394 VTAIL.n393 1.16414
R760 VTAIL.n433 VTAIL.n334 1.16414
R761 VTAIL.n55 VTAIL.n26 1.16414
R762 VTAIL.n64 VTAIL.n63 1.16414
R763 VTAIL.n103 VTAIL.n4 1.16414
R764 VTAIL.n327 VTAIL.n228 1.16414
R765 VTAIL.n288 VTAIL.n287 1.16414
R766 VTAIL.n279 VTAIL.n250 1.16414
R767 VTAIL.n217 VTAIL.n118 1.16414
R768 VTAIL.n178 VTAIL.n177 1.16414
R769 VTAIL.n169 VTAIL.n140 1.16414
R770 VTAIL VTAIL.n439 0.838862
R771 VTAIL.n389 VTAIL.n388 0.388379
R772 VTAIL.n390 VTAIL.n354 0.388379
R773 VTAIL.n59 VTAIL.n58 0.388379
R774 VTAIL.n60 VTAIL.n24 0.388379
R775 VTAIL.n284 VTAIL.n248 0.388379
R776 VTAIL.n283 VTAIL.n282 0.388379
R777 VTAIL.n174 VTAIL.n138 0.388379
R778 VTAIL.n173 VTAIL.n172 0.388379
R779 VTAIL.n370 VTAIL.n369 0.155672
R780 VTAIL.n370 VTAIL.n361 0.155672
R781 VTAIL.n377 VTAIL.n361 0.155672
R782 VTAIL.n378 VTAIL.n377 0.155672
R783 VTAIL.n378 VTAIL.n357 0.155672
R784 VTAIL.n386 VTAIL.n357 0.155672
R785 VTAIL.n387 VTAIL.n386 0.155672
R786 VTAIL.n387 VTAIL.n353 0.155672
R787 VTAIL.n395 VTAIL.n353 0.155672
R788 VTAIL.n396 VTAIL.n395 0.155672
R789 VTAIL.n396 VTAIL.n349 0.155672
R790 VTAIL.n403 VTAIL.n349 0.155672
R791 VTAIL.n404 VTAIL.n403 0.155672
R792 VTAIL.n404 VTAIL.n345 0.155672
R793 VTAIL.n411 VTAIL.n345 0.155672
R794 VTAIL.n412 VTAIL.n411 0.155672
R795 VTAIL.n412 VTAIL.n341 0.155672
R796 VTAIL.n419 VTAIL.n341 0.155672
R797 VTAIL.n420 VTAIL.n419 0.155672
R798 VTAIL.n420 VTAIL.n337 0.155672
R799 VTAIL.n427 VTAIL.n337 0.155672
R800 VTAIL.n428 VTAIL.n427 0.155672
R801 VTAIL.n428 VTAIL.n333 0.155672
R802 VTAIL.n435 VTAIL.n333 0.155672
R803 VTAIL.n40 VTAIL.n39 0.155672
R804 VTAIL.n40 VTAIL.n31 0.155672
R805 VTAIL.n47 VTAIL.n31 0.155672
R806 VTAIL.n48 VTAIL.n47 0.155672
R807 VTAIL.n48 VTAIL.n27 0.155672
R808 VTAIL.n56 VTAIL.n27 0.155672
R809 VTAIL.n57 VTAIL.n56 0.155672
R810 VTAIL.n57 VTAIL.n23 0.155672
R811 VTAIL.n65 VTAIL.n23 0.155672
R812 VTAIL.n66 VTAIL.n65 0.155672
R813 VTAIL.n66 VTAIL.n19 0.155672
R814 VTAIL.n73 VTAIL.n19 0.155672
R815 VTAIL.n74 VTAIL.n73 0.155672
R816 VTAIL.n74 VTAIL.n15 0.155672
R817 VTAIL.n81 VTAIL.n15 0.155672
R818 VTAIL.n82 VTAIL.n81 0.155672
R819 VTAIL.n82 VTAIL.n11 0.155672
R820 VTAIL.n89 VTAIL.n11 0.155672
R821 VTAIL.n90 VTAIL.n89 0.155672
R822 VTAIL.n90 VTAIL.n7 0.155672
R823 VTAIL.n97 VTAIL.n7 0.155672
R824 VTAIL.n98 VTAIL.n97 0.155672
R825 VTAIL.n98 VTAIL.n3 0.155672
R826 VTAIL.n105 VTAIL.n3 0.155672
R827 VTAIL.n329 VTAIL.n227 0.155672
R828 VTAIL.n322 VTAIL.n227 0.155672
R829 VTAIL.n322 VTAIL.n321 0.155672
R830 VTAIL.n321 VTAIL.n231 0.155672
R831 VTAIL.n314 VTAIL.n231 0.155672
R832 VTAIL.n314 VTAIL.n313 0.155672
R833 VTAIL.n313 VTAIL.n235 0.155672
R834 VTAIL.n306 VTAIL.n235 0.155672
R835 VTAIL.n306 VTAIL.n305 0.155672
R836 VTAIL.n305 VTAIL.n239 0.155672
R837 VTAIL.n298 VTAIL.n239 0.155672
R838 VTAIL.n298 VTAIL.n297 0.155672
R839 VTAIL.n297 VTAIL.n243 0.155672
R840 VTAIL.n290 VTAIL.n243 0.155672
R841 VTAIL.n290 VTAIL.n289 0.155672
R842 VTAIL.n289 VTAIL.n247 0.155672
R843 VTAIL.n281 VTAIL.n247 0.155672
R844 VTAIL.n281 VTAIL.n280 0.155672
R845 VTAIL.n280 VTAIL.n251 0.155672
R846 VTAIL.n273 VTAIL.n251 0.155672
R847 VTAIL.n273 VTAIL.n272 0.155672
R848 VTAIL.n272 VTAIL.n256 0.155672
R849 VTAIL.n265 VTAIL.n256 0.155672
R850 VTAIL.n265 VTAIL.n264 0.155672
R851 VTAIL.n219 VTAIL.n117 0.155672
R852 VTAIL.n212 VTAIL.n117 0.155672
R853 VTAIL.n212 VTAIL.n211 0.155672
R854 VTAIL.n211 VTAIL.n121 0.155672
R855 VTAIL.n204 VTAIL.n121 0.155672
R856 VTAIL.n204 VTAIL.n203 0.155672
R857 VTAIL.n203 VTAIL.n125 0.155672
R858 VTAIL.n196 VTAIL.n125 0.155672
R859 VTAIL.n196 VTAIL.n195 0.155672
R860 VTAIL.n195 VTAIL.n129 0.155672
R861 VTAIL.n188 VTAIL.n129 0.155672
R862 VTAIL.n188 VTAIL.n187 0.155672
R863 VTAIL.n187 VTAIL.n133 0.155672
R864 VTAIL.n180 VTAIL.n133 0.155672
R865 VTAIL.n180 VTAIL.n179 0.155672
R866 VTAIL.n179 VTAIL.n137 0.155672
R867 VTAIL.n171 VTAIL.n137 0.155672
R868 VTAIL.n171 VTAIL.n170 0.155672
R869 VTAIL.n170 VTAIL.n141 0.155672
R870 VTAIL.n163 VTAIL.n141 0.155672
R871 VTAIL.n163 VTAIL.n162 0.155672
R872 VTAIL.n162 VTAIL.n146 0.155672
R873 VTAIL.n155 VTAIL.n146 0.155672
R874 VTAIL.n155 VTAIL.n154 0.155672
R875 VDD1.n101 VDD1.n100 585
R876 VDD1.n99 VDD1.n98 585
R877 VDD1.n4 VDD1.n3 585
R878 VDD1.n93 VDD1.n92 585
R879 VDD1.n91 VDD1.n90 585
R880 VDD1.n8 VDD1.n7 585
R881 VDD1.n85 VDD1.n84 585
R882 VDD1.n83 VDD1.n82 585
R883 VDD1.n12 VDD1.n11 585
R884 VDD1.n77 VDD1.n76 585
R885 VDD1.n75 VDD1.n74 585
R886 VDD1.n16 VDD1.n15 585
R887 VDD1.n69 VDD1.n68 585
R888 VDD1.n67 VDD1.n66 585
R889 VDD1.n20 VDD1.n19 585
R890 VDD1.n61 VDD1.n60 585
R891 VDD1.n59 VDD1.n58 585
R892 VDD1.n57 VDD1.n23 585
R893 VDD1.n27 VDD1.n24 585
R894 VDD1.n52 VDD1.n51 585
R895 VDD1.n50 VDD1.n49 585
R896 VDD1.n29 VDD1.n28 585
R897 VDD1.n44 VDD1.n43 585
R898 VDD1.n42 VDD1.n41 585
R899 VDD1.n33 VDD1.n32 585
R900 VDD1.n36 VDD1.n35 585
R901 VDD1.n142 VDD1.n141 585
R902 VDD1.n139 VDD1.n138 585
R903 VDD1.n148 VDD1.n147 585
R904 VDD1.n150 VDD1.n149 585
R905 VDD1.n135 VDD1.n134 585
R906 VDD1.n156 VDD1.n155 585
R907 VDD1.n159 VDD1.n158 585
R908 VDD1.n157 VDD1.n131 585
R909 VDD1.n164 VDD1.n130 585
R910 VDD1.n166 VDD1.n165 585
R911 VDD1.n168 VDD1.n167 585
R912 VDD1.n127 VDD1.n126 585
R913 VDD1.n174 VDD1.n173 585
R914 VDD1.n176 VDD1.n175 585
R915 VDD1.n123 VDD1.n122 585
R916 VDD1.n182 VDD1.n181 585
R917 VDD1.n184 VDD1.n183 585
R918 VDD1.n119 VDD1.n118 585
R919 VDD1.n190 VDD1.n189 585
R920 VDD1.n192 VDD1.n191 585
R921 VDD1.n115 VDD1.n114 585
R922 VDD1.n198 VDD1.n197 585
R923 VDD1.n200 VDD1.n199 585
R924 VDD1.n111 VDD1.n110 585
R925 VDD1.n206 VDD1.n205 585
R926 VDD1.n208 VDD1.n207 585
R927 VDD1.n100 VDD1.n0 498.474
R928 VDD1.n207 VDD1.n107 498.474
R929 VDD1.t9 VDD1.n34 329.036
R930 VDD1.t8 VDD1.n140 329.036
R931 VDD1.n100 VDD1.n99 171.744
R932 VDD1.n99 VDD1.n3 171.744
R933 VDD1.n92 VDD1.n3 171.744
R934 VDD1.n92 VDD1.n91 171.744
R935 VDD1.n91 VDD1.n7 171.744
R936 VDD1.n84 VDD1.n7 171.744
R937 VDD1.n84 VDD1.n83 171.744
R938 VDD1.n83 VDD1.n11 171.744
R939 VDD1.n76 VDD1.n11 171.744
R940 VDD1.n76 VDD1.n75 171.744
R941 VDD1.n75 VDD1.n15 171.744
R942 VDD1.n68 VDD1.n15 171.744
R943 VDD1.n68 VDD1.n67 171.744
R944 VDD1.n67 VDD1.n19 171.744
R945 VDD1.n60 VDD1.n19 171.744
R946 VDD1.n60 VDD1.n59 171.744
R947 VDD1.n59 VDD1.n23 171.744
R948 VDD1.n27 VDD1.n23 171.744
R949 VDD1.n51 VDD1.n27 171.744
R950 VDD1.n51 VDD1.n50 171.744
R951 VDD1.n50 VDD1.n28 171.744
R952 VDD1.n43 VDD1.n28 171.744
R953 VDD1.n43 VDD1.n42 171.744
R954 VDD1.n42 VDD1.n32 171.744
R955 VDD1.n35 VDD1.n32 171.744
R956 VDD1.n141 VDD1.n138 171.744
R957 VDD1.n148 VDD1.n138 171.744
R958 VDD1.n149 VDD1.n148 171.744
R959 VDD1.n149 VDD1.n134 171.744
R960 VDD1.n156 VDD1.n134 171.744
R961 VDD1.n158 VDD1.n156 171.744
R962 VDD1.n158 VDD1.n157 171.744
R963 VDD1.n157 VDD1.n130 171.744
R964 VDD1.n166 VDD1.n130 171.744
R965 VDD1.n167 VDD1.n166 171.744
R966 VDD1.n167 VDD1.n126 171.744
R967 VDD1.n174 VDD1.n126 171.744
R968 VDD1.n175 VDD1.n174 171.744
R969 VDD1.n175 VDD1.n122 171.744
R970 VDD1.n182 VDD1.n122 171.744
R971 VDD1.n183 VDD1.n182 171.744
R972 VDD1.n183 VDD1.n118 171.744
R973 VDD1.n190 VDD1.n118 171.744
R974 VDD1.n191 VDD1.n190 171.744
R975 VDD1.n191 VDD1.n114 171.744
R976 VDD1.n198 VDD1.n114 171.744
R977 VDD1.n199 VDD1.n198 171.744
R978 VDD1.n199 VDD1.n110 171.744
R979 VDD1.n206 VDD1.n110 171.744
R980 VDD1.n207 VDD1.n206 171.744
R981 VDD1.n35 VDD1.t9 85.8723
R982 VDD1.n141 VDD1.t8 85.8723
R983 VDD1.n215 VDD1.n214 74.3562
R984 VDD1.n106 VDD1.n105 71.722
R985 VDD1.n217 VDD1.n216 71.7219
R986 VDD1.n213 VDD1.n212 71.7219
R987 VDD1.n217 VDD1.n215 59.9535
R988 VDD1.n106 VDD1.n104 56.3291
R989 VDD1.n213 VDD1.n211 56.3291
R990 VDD1.n58 VDD1.n57 13.1884
R991 VDD1.n165 VDD1.n164 13.1884
R992 VDD1.n102 VDD1.n101 12.8005
R993 VDD1.n61 VDD1.n22 12.8005
R994 VDD1.n56 VDD1.n24 12.8005
R995 VDD1.n163 VDD1.n131 12.8005
R996 VDD1.n168 VDD1.n129 12.8005
R997 VDD1.n209 VDD1.n208 12.8005
R998 VDD1.n98 VDD1.n2 12.0247
R999 VDD1.n62 VDD1.n20 12.0247
R1000 VDD1.n53 VDD1.n52 12.0247
R1001 VDD1.n160 VDD1.n159 12.0247
R1002 VDD1.n169 VDD1.n127 12.0247
R1003 VDD1.n205 VDD1.n109 12.0247
R1004 VDD1.n97 VDD1.n4 11.249
R1005 VDD1.n66 VDD1.n65 11.249
R1006 VDD1.n49 VDD1.n26 11.249
R1007 VDD1.n155 VDD1.n133 11.249
R1008 VDD1.n173 VDD1.n172 11.249
R1009 VDD1.n204 VDD1.n111 11.249
R1010 VDD1.n36 VDD1.n34 10.7239
R1011 VDD1.n142 VDD1.n140 10.7239
R1012 VDD1.n94 VDD1.n93 10.4732
R1013 VDD1.n69 VDD1.n18 10.4732
R1014 VDD1.n48 VDD1.n29 10.4732
R1015 VDD1.n154 VDD1.n135 10.4732
R1016 VDD1.n176 VDD1.n125 10.4732
R1017 VDD1.n201 VDD1.n200 10.4732
R1018 VDD1.n90 VDD1.n6 9.69747
R1019 VDD1.n70 VDD1.n16 9.69747
R1020 VDD1.n45 VDD1.n44 9.69747
R1021 VDD1.n151 VDD1.n150 9.69747
R1022 VDD1.n177 VDD1.n123 9.69747
R1023 VDD1.n197 VDD1.n113 9.69747
R1024 VDD1.n104 VDD1.n103 9.45567
R1025 VDD1.n211 VDD1.n210 9.45567
R1026 VDD1.n38 VDD1.n37 9.3005
R1027 VDD1.n40 VDD1.n39 9.3005
R1028 VDD1.n31 VDD1.n30 9.3005
R1029 VDD1.n46 VDD1.n45 9.3005
R1030 VDD1.n48 VDD1.n47 9.3005
R1031 VDD1.n26 VDD1.n25 9.3005
R1032 VDD1.n54 VDD1.n53 9.3005
R1033 VDD1.n56 VDD1.n55 9.3005
R1034 VDD1.n10 VDD1.n9 9.3005
R1035 VDD1.n87 VDD1.n86 9.3005
R1036 VDD1.n89 VDD1.n88 9.3005
R1037 VDD1.n6 VDD1.n5 9.3005
R1038 VDD1.n95 VDD1.n94 9.3005
R1039 VDD1.n97 VDD1.n96 9.3005
R1040 VDD1.n2 VDD1.n1 9.3005
R1041 VDD1.n103 VDD1.n102 9.3005
R1042 VDD1.n81 VDD1.n80 9.3005
R1043 VDD1.n79 VDD1.n78 9.3005
R1044 VDD1.n14 VDD1.n13 9.3005
R1045 VDD1.n73 VDD1.n72 9.3005
R1046 VDD1.n71 VDD1.n70 9.3005
R1047 VDD1.n18 VDD1.n17 9.3005
R1048 VDD1.n65 VDD1.n64 9.3005
R1049 VDD1.n63 VDD1.n62 9.3005
R1050 VDD1.n22 VDD1.n21 9.3005
R1051 VDD1.n186 VDD1.n185 9.3005
R1052 VDD1.n121 VDD1.n120 9.3005
R1053 VDD1.n180 VDD1.n179 9.3005
R1054 VDD1.n178 VDD1.n177 9.3005
R1055 VDD1.n125 VDD1.n124 9.3005
R1056 VDD1.n172 VDD1.n171 9.3005
R1057 VDD1.n170 VDD1.n169 9.3005
R1058 VDD1.n129 VDD1.n128 9.3005
R1059 VDD1.n144 VDD1.n143 9.3005
R1060 VDD1.n146 VDD1.n145 9.3005
R1061 VDD1.n137 VDD1.n136 9.3005
R1062 VDD1.n152 VDD1.n151 9.3005
R1063 VDD1.n154 VDD1.n153 9.3005
R1064 VDD1.n133 VDD1.n132 9.3005
R1065 VDD1.n161 VDD1.n160 9.3005
R1066 VDD1.n163 VDD1.n162 9.3005
R1067 VDD1.n188 VDD1.n187 9.3005
R1068 VDD1.n117 VDD1.n116 9.3005
R1069 VDD1.n194 VDD1.n193 9.3005
R1070 VDD1.n196 VDD1.n195 9.3005
R1071 VDD1.n113 VDD1.n112 9.3005
R1072 VDD1.n202 VDD1.n201 9.3005
R1073 VDD1.n204 VDD1.n203 9.3005
R1074 VDD1.n109 VDD1.n108 9.3005
R1075 VDD1.n210 VDD1.n209 9.3005
R1076 VDD1.n89 VDD1.n8 8.92171
R1077 VDD1.n74 VDD1.n73 8.92171
R1078 VDD1.n41 VDD1.n31 8.92171
R1079 VDD1.n147 VDD1.n137 8.92171
R1080 VDD1.n181 VDD1.n180 8.92171
R1081 VDD1.n196 VDD1.n115 8.92171
R1082 VDD1.n86 VDD1.n85 8.14595
R1083 VDD1.n77 VDD1.n14 8.14595
R1084 VDD1.n40 VDD1.n33 8.14595
R1085 VDD1.n146 VDD1.n139 8.14595
R1086 VDD1.n184 VDD1.n121 8.14595
R1087 VDD1.n193 VDD1.n192 8.14595
R1088 VDD1.n104 VDD1.n0 7.75445
R1089 VDD1.n211 VDD1.n107 7.75445
R1090 VDD1.n82 VDD1.n10 7.3702
R1091 VDD1.n78 VDD1.n12 7.3702
R1092 VDD1.n37 VDD1.n36 7.3702
R1093 VDD1.n143 VDD1.n142 7.3702
R1094 VDD1.n185 VDD1.n119 7.3702
R1095 VDD1.n189 VDD1.n117 7.3702
R1096 VDD1.n82 VDD1.n81 6.59444
R1097 VDD1.n81 VDD1.n12 6.59444
R1098 VDD1.n188 VDD1.n119 6.59444
R1099 VDD1.n189 VDD1.n188 6.59444
R1100 VDD1.n102 VDD1.n0 6.08283
R1101 VDD1.n209 VDD1.n107 6.08283
R1102 VDD1.n85 VDD1.n10 5.81868
R1103 VDD1.n78 VDD1.n77 5.81868
R1104 VDD1.n37 VDD1.n33 5.81868
R1105 VDD1.n143 VDD1.n139 5.81868
R1106 VDD1.n185 VDD1.n184 5.81868
R1107 VDD1.n192 VDD1.n117 5.81868
R1108 VDD1.n86 VDD1.n8 5.04292
R1109 VDD1.n74 VDD1.n14 5.04292
R1110 VDD1.n41 VDD1.n40 5.04292
R1111 VDD1.n147 VDD1.n146 5.04292
R1112 VDD1.n181 VDD1.n121 5.04292
R1113 VDD1.n193 VDD1.n115 5.04292
R1114 VDD1.n90 VDD1.n89 4.26717
R1115 VDD1.n73 VDD1.n16 4.26717
R1116 VDD1.n44 VDD1.n31 4.26717
R1117 VDD1.n150 VDD1.n137 4.26717
R1118 VDD1.n180 VDD1.n123 4.26717
R1119 VDD1.n197 VDD1.n196 4.26717
R1120 VDD1.n93 VDD1.n6 3.49141
R1121 VDD1.n70 VDD1.n69 3.49141
R1122 VDD1.n45 VDD1.n29 3.49141
R1123 VDD1.n151 VDD1.n135 3.49141
R1124 VDD1.n177 VDD1.n176 3.49141
R1125 VDD1.n200 VDD1.n113 3.49141
R1126 VDD1.n94 VDD1.n4 2.71565
R1127 VDD1.n66 VDD1.n18 2.71565
R1128 VDD1.n49 VDD1.n48 2.71565
R1129 VDD1.n155 VDD1.n154 2.71565
R1130 VDD1.n173 VDD1.n125 2.71565
R1131 VDD1.n201 VDD1.n111 2.71565
R1132 VDD1 VDD1.n217 2.63197
R1133 VDD1.n38 VDD1.n34 2.41282
R1134 VDD1.n144 VDD1.n140 2.41282
R1135 VDD1.n98 VDD1.n97 1.93989
R1136 VDD1.n65 VDD1.n20 1.93989
R1137 VDD1.n52 VDD1.n26 1.93989
R1138 VDD1.n159 VDD1.n133 1.93989
R1139 VDD1.n172 VDD1.n127 1.93989
R1140 VDD1.n205 VDD1.n204 1.93989
R1141 VDD1.n216 VDD1.t4 1.66572
R1142 VDD1.n216 VDD1.t5 1.66572
R1143 VDD1.n105 VDD1.t6 1.66572
R1144 VDD1.n105 VDD1.t7 1.66572
R1145 VDD1.n214 VDD1.t2 1.66572
R1146 VDD1.n214 VDD1.t1 1.66572
R1147 VDD1.n212 VDD1.t3 1.66572
R1148 VDD1.n212 VDD1.t0 1.66572
R1149 VDD1.n101 VDD1.n2 1.16414
R1150 VDD1.n62 VDD1.n61 1.16414
R1151 VDD1.n53 VDD1.n24 1.16414
R1152 VDD1.n160 VDD1.n131 1.16414
R1153 VDD1.n169 VDD1.n168 1.16414
R1154 VDD1.n208 VDD1.n109 1.16414
R1155 VDD1 VDD1.n106 0.955241
R1156 VDD1.n215 VDD1.n213 0.841706
R1157 VDD1.n58 VDD1.n22 0.388379
R1158 VDD1.n57 VDD1.n56 0.388379
R1159 VDD1.n164 VDD1.n163 0.388379
R1160 VDD1.n165 VDD1.n129 0.388379
R1161 VDD1.n103 VDD1.n1 0.155672
R1162 VDD1.n96 VDD1.n1 0.155672
R1163 VDD1.n96 VDD1.n95 0.155672
R1164 VDD1.n95 VDD1.n5 0.155672
R1165 VDD1.n88 VDD1.n5 0.155672
R1166 VDD1.n88 VDD1.n87 0.155672
R1167 VDD1.n87 VDD1.n9 0.155672
R1168 VDD1.n80 VDD1.n9 0.155672
R1169 VDD1.n80 VDD1.n79 0.155672
R1170 VDD1.n79 VDD1.n13 0.155672
R1171 VDD1.n72 VDD1.n13 0.155672
R1172 VDD1.n72 VDD1.n71 0.155672
R1173 VDD1.n71 VDD1.n17 0.155672
R1174 VDD1.n64 VDD1.n17 0.155672
R1175 VDD1.n64 VDD1.n63 0.155672
R1176 VDD1.n63 VDD1.n21 0.155672
R1177 VDD1.n55 VDD1.n21 0.155672
R1178 VDD1.n55 VDD1.n54 0.155672
R1179 VDD1.n54 VDD1.n25 0.155672
R1180 VDD1.n47 VDD1.n25 0.155672
R1181 VDD1.n47 VDD1.n46 0.155672
R1182 VDD1.n46 VDD1.n30 0.155672
R1183 VDD1.n39 VDD1.n30 0.155672
R1184 VDD1.n39 VDD1.n38 0.155672
R1185 VDD1.n145 VDD1.n144 0.155672
R1186 VDD1.n145 VDD1.n136 0.155672
R1187 VDD1.n152 VDD1.n136 0.155672
R1188 VDD1.n153 VDD1.n152 0.155672
R1189 VDD1.n153 VDD1.n132 0.155672
R1190 VDD1.n161 VDD1.n132 0.155672
R1191 VDD1.n162 VDD1.n161 0.155672
R1192 VDD1.n162 VDD1.n128 0.155672
R1193 VDD1.n170 VDD1.n128 0.155672
R1194 VDD1.n171 VDD1.n170 0.155672
R1195 VDD1.n171 VDD1.n124 0.155672
R1196 VDD1.n178 VDD1.n124 0.155672
R1197 VDD1.n179 VDD1.n178 0.155672
R1198 VDD1.n179 VDD1.n120 0.155672
R1199 VDD1.n186 VDD1.n120 0.155672
R1200 VDD1.n187 VDD1.n186 0.155672
R1201 VDD1.n187 VDD1.n116 0.155672
R1202 VDD1.n194 VDD1.n116 0.155672
R1203 VDD1.n195 VDD1.n194 0.155672
R1204 VDD1.n195 VDD1.n112 0.155672
R1205 VDD1.n202 VDD1.n112 0.155672
R1206 VDD1.n203 VDD1.n202 0.155672
R1207 VDD1.n203 VDD1.n108 0.155672
R1208 VDD1.n210 VDD1.n108 0.155672
R1209 VN.n110 VN.n109 161.3
R1210 VN.n108 VN.n57 161.3
R1211 VN.n107 VN.n106 161.3
R1212 VN.n105 VN.n58 161.3
R1213 VN.n104 VN.n103 161.3
R1214 VN.n102 VN.n59 161.3
R1215 VN.n101 VN.n100 161.3
R1216 VN.n99 VN.n60 161.3
R1217 VN.n98 VN.n97 161.3
R1218 VN.n95 VN.n61 161.3
R1219 VN.n94 VN.n93 161.3
R1220 VN.n92 VN.n62 161.3
R1221 VN.n91 VN.n90 161.3
R1222 VN.n89 VN.n63 161.3
R1223 VN.n88 VN.n87 161.3
R1224 VN.n86 VN.n64 161.3
R1225 VN.n85 VN.n84 161.3
R1226 VN.n82 VN.n65 161.3
R1227 VN.n81 VN.n80 161.3
R1228 VN.n79 VN.n66 161.3
R1229 VN.n78 VN.n77 161.3
R1230 VN.n76 VN.n67 161.3
R1231 VN.n75 VN.n74 161.3
R1232 VN.n73 VN.n68 161.3
R1233 VN.n72 VN.n71 161.3
R1234 VN.n54 VN.n53 161.3
R1235 VN.n52 VN.n1 161.3
R1236 VN.n51 VN.n50 161.3
R1237 VN.n49 VN.n2 161.3
R1238 VN.n48 VN.n47 161.3
R1239 VN.n46 VN.n3 161.3
R1240 VN.n45 VN.n44 161.3
R1241 VN.n43 VN.n4 161.3
R1242 VN.n42 VN.n41 161.3
R1243 VN.n39 VN.n5 161.3
R1244 VN.n38 VN.n37 161.3
R1245 VN.n36 VN.n6 161.3
R1246 VN.n35 VN.n34 161.3
R1247 VN.n33 VN.n7 161.3
R1248 VN.n32 VN.n31 161.3
R1249 VN.n30 VN.n8 161.3
R1250 VN.n29 VN.n28 161.3
R1251 VN.n26 VN.n9 161.3
R1252 VN.n25 VN.n24 161.3
R1253 VN.n23 VN.n10 161.3
R1254 VN.n22 VN.n21 161.3
R1255 VN.n20 VN.n11 161.3
R1256 VN.n19 VN.n18 161.3
R1257 VN.n17 VN.n12 161.3
R1258 VN.n16 VN.n15 161.3
R1259 VN.n69 VN.t5 155.917
R1260 VN.n13 VN.t4 155.917
R1261 VN.n14 VN.t3 122.829
R1262 VN.n27 VN.t8 122.829
R1263 VN.n40 VN.t9 122.829
R1264 VN.n0 VN.t7 122.829
R1265 VN.n70 VN.t6 122.829
R1266 VN.n83 VN.t2 122.829
R1267 VN.n96 VN.t1 122.829
R1268 VN.n56 VN.t0 122.829
R1269 VN.n55 VN.n0 86.8027
R1270 VN.n111 VN.n56 86.8027
R1271 VN VN.n111 65.733
R1272 VN.n21 VN.n20 56.5617
R1273 VN.n34 VN.n33 56.5617
R1274 VN.n77 VN.n76 56.5617
R1275 VN.n90 VN.n89 56.5617
R1276 VN.n14 VN.n13 55.106
R1277 VN.n70 VN.n69 55.106
R1278 VN.n47 VN.n46 41.5458
R1279 VN.n103 VN.n102 41.5458
R1280 VN.n47 VN.n2 39.6083
R1281 VN.n103 VN.n58 39.6083
R1282 VN.n15 VN.n12 24.5923
R1283 VN.n19 VN.n12 24.5923
R1284 VN.n20 VN.n19 24.5923
R1285 VN.n21 VN.n10 24.5923
R1286 VN.n25 VN.n10 24.5923
R1287 VN.n26 VN.n25 24.5923
R1288 VN.n28 VN.n8 24.5923
R1289 VN.n32 VN.n8 24.5923
R1290 VN.n33 VN.n32 24.5923
R1291 VN.n34 VN.n6 24.5923
R1292 VN.n38 VN.n6 24.5923
R1293 VN.n39 VN.n38 24.5923
R1294 VN.n41 VN.n4 24.5923
R1295 VN.n45 VN.n4 24.5923
R1296 VN.n46 VN.n45 24.5923
R1297 VN.n51 VN.n2 24.5923
R1298 VN.n52 VN.n51 24.5923
R1299 VN.n53 VN.n52 24.5923
R1300 VN.n76 VN.n75 24.5923
R1301 VN.n75 VN.n68 24.5923
R1302 VN.n71 VN.n68 24.5923
R1303 VN.n89 VN.n88 24.5923
R1304 VN.n88 VN.n64 24.5923
R1305 VN.n84 VN.n64 24.5923
R1306 VN.n82 VN.n81 24.5923
R1307 VN.n81 VN.n66 24.5923
R1308 VN.n77 VN.n66 24.5923
R1309 VN.n102 VN.n101 24.5923
R1310 VN.n101 VN.n60 24.5923
R1311 VN.n97 VN.n60 24.5923
R1312 VN.n95 VN.n94 24.5923
R1313 VN.n94 VN.n62 24.5923
R1314 VN.n90 VN.n62 24.5923
R1315 VN.n109 VN.n108 24.5923
R1316 VN.n108 VN.n107 24.5923
R1317 VN.n107 VN.n58 24.5923
R1318 VN.n15 VN.n14 20.1658
R1319 VN.n40 VN.n39 20.1658
R1320 VN.n71 VN.n70 20.1658
R1321 VN.n96 VN.n95 20.1658
R1322 VN.n27 VN.n26 12.2964
R1323 VN.n28 VN.n27 12.2964
R1324 VN.n84 VN.n83 12.2964
R1325 VN.n83 VN.n82 12.2964
R1326 VN.n41 VN.n40 4.42703
R1327 VN.n97 VN.n96 4.42703
R1328 VN.n53 VN.n0 3.44336
R1329 VN.n109 VN.n56 3.44336
R1330 VN.n16 VN.n13 2.44069
R1331 VN.n72 VN.n69 2.44069
R1332 VN.n111 VN.n110 0.354861
R1333 VN.n55 VN.n54 0.354861
R1334 VN VN.n55 0.267071
R1335 VN.n110 VN.n57 0.189894
R1336 VN.n106 VN.n57 0.189894
R1337 VN.n106 VN.n105 0.189894
R1338 VN.n105 VN.n104 0.189894
R1339 VN.n104 VN.n59 0.189894
R1340 VN.n100 VN.n59 0.189894
R1341 VN.n100 VN.n99 0.189894
R1342 VN.n99 VN.n98 0.189894
R1343 VN.n98 VN.n61 0.189894
R1344 VN.n93 VN.n61 0.189894
R1345 VN.n93 VN.n92 0.189894
R1346 VN.n92 VN.n91 0.189894
R1347 VN.n91 VN.n63 0.189894
R1348 VN.n87 VN.n63 0.189894
R1349 VN.n87 VN.n86 0.189894
R1350 VN.n86 VN.n85 0.189894
R1351 VN.n85 VN.n65 0.189894
R1352 VN.n80 VN.n65 0.189894
R1353 VN.n80 VN.n79 0.189894
R1354 VN.n79 VN.n78 0.189894
R1355 VN.n78 VN.n67 0.189894
R1356 VN.n74 VN.n67 0.189894
R1357 VN.n74 VN.n73 0.189894
R1358 VN.n73 VN.n72 0.189894
R1359 VN.n17 VN.n16 0.189894
R1360 VN.n18 VN.n17 0.189894
R1361 VN.n18 VN.n11 0.189894
R1362 VN.n22 VN.n11 0.189894
R1363 VN.n23 VN.n22 0.189894
R1364 VN.n24 VN.n23 0.189894
R1365 VN.n24 VN.n9 0.189894
R1366 VN.n29 VN.n9 0.189894
R1367 VN.n30 VN.n29 0.189894
R1368 VN.n31 VN.n30 0.189894
R1369 VN.n31 VN.n7 0.189894
R1370 VN.n35 VN.n7 0.189894
R1371 VN.n36 VN.n35 0.189894
R1372 VN.n37 VN.n36 0.189894
R1373 VN.n37 VN.n5 0.189894
R1374 VN.n42 VN.n5 0.189894
R1375 VN.n43 VN.n42 0.189894
R1376 VN.n44 VN.n43 0.189894
R1377 VN.n44 VN.n3 0.189894
R1378 VN.n48 VN.n3 0.189894
R1379 VN.n49 VN.n48 0.189894
R1380 VN.n50 VN.n49 0.189894
R1381 VN.n50 VN.n1 0.189894
R1382 VN.n54 VN.n1 0.189894
R1383 VDD2.n210 VDD2.n209 585
R1384 VDD2.n208 VDD2.n207 585
R1385 VDD2.n113 VDD2.n112 585
R1386 VDD2.n202 VDD2.n201 585
R1387 VDD2.n200 VDD2.n199 585
R1388 VDD2.n117 VDD2.n116 585
R1389 VDD2.n194 VDD2.n193 585
R1390 VDD2.n192 VDD2.n191 585
R1391 VDD2.n121 VDD2.n120 585
R1392 VDD2.n186 VDD2.n185 585
R1393 VDD2.n184 VDD2.n183 585
R1394 VDD2.n125 VDD2.n124 585
R1395 VDD2.n178 VDD2.n177 585
R1396 VDD2.n176 VDD2.n175 585
R1397 VDD2.n129 VDD2.n128 585
R1398 VDD2.n170 VDD2.n169 585
R1399 VDD2.n168 VDD2.n167 585
R1400 VDD2.n166 VDD2.n132 585
R1401 VDD2.n136 VDD2.n133 585
R1402 VDD2.n161 VDD2.n160 585
R1403 VDD2.n159 VDD2.n158 585
R1404 VDD2.n138 VDD2.n137 585
R1405 VDD2.n153 VDD2.n152 585
R1406 VDD2.n151 VDD2.n150 585
R1407 VDD2.n142 VDD2.n141 585
R1408 VDD2.n145 VDD2.n144 585
R1409 VDD2.n35 VDD2.n34 585
R1410 VDD2.n32 VDD2.n31 585
R1411 VDD2.n41 VDD2.n40 585
R1412 VDD2.n43 VDD2.n42 585
R1413 VDD2.n28 VDD2.n27 585
R1414 VDD2.n49 VDD2.n48 585
R1415 VDD2.n52 VDD2.n51 585
R1416 VDD2.n50 VDD2.n24 585
R1417 VDD2.n57 VDD2.n23 585
R1418 VDD2.n59 VDD2.n58 585
R1419 VDD2.n61 VDD2.n60 585
R1420 VDD2.n20 VDD2.n19 585
R1421 VDD2.n67 VDD2.n66 585
R1422 VDD2.n69 VDD2.n68 585
R1423 VDD2.n16 VDD2.n15 585
R1424 VDD2.n75 VDD2.n74 585
R1425 VDD2.n77 VDD2.n76 585
R1426 VDD2.n12 VDD2.n11 585
R1427 VDD2.n83 VDD2.n82 585
R1428 VDD2.n85 VDD2.n84 585
R1429 VDD2.n8 VDD2.n7 585
R1430 VDD2.n91 VDD2.n90 585
R1431 VDD2.n93 VDD2.n92 585
R1432 VDD2.n4 VDD2.n3 585
R1433 VDD2.n99 VDD2.n98 585
R1434 VDD2.n101 VDD2.n100 585
R1435 VDD2.n209 VDD2.n109 498.474
R1436 VDD2.n100 VDD2.n0 498.474
R1437 VDD2.t9 VDD2.n143 329.036
R1438 VDD2.t5 VDD2.n33 329.036
R1439 VDD2.n209 VDD2.n208 171.744
R1440 VDD2.n208 VDD2.n112 171.744
R1441 VDD2.n201 VDD2.n112 171.744
R1442 VDD2.n201 VDD2.n200 171.744
R1443 VDD2.n200 VDD2.n116 171.744
R1444 VDD2.n193 VDD2.n116 171.744
R1445 VDD2.n193 VDD2.n192 171.744
R1446 VDD2.n192 VDD2.n120 171.744
R1447 VDD2.n185 VDD2.n120 171.744
R1448 VDD2.n185 VDD2.n184 171.744
R1449 VDD2.n184 VDD2.n124 171.744
R1450 VDD2.n177 VDD2.n124 171.744
R1451 VDD2.n177 VDD2.n176 171.744
R1452 VDD2.n176 VDD2.n128 171.744
R1453 VDD2.n169 VDD2.n128 171.744
R1454 VDD2.n169 VDD2.n168 171.744
R1455 VDD2.n168 VDD2.n132 171.744
R1456 VDD2.n136 VDD2.n132 171.744
R1457 VDD2.n160 VDD2.n136 171.744
R1458 VDD2.n160 VDD2.n159 171.744
R1459 VDD2.n159 VDD2.n137 171.744
R1460 VDD2.n152 VDD2.n137 171.744
R1461 VDD2.n152 VDD2.n151 171.744
R1462 VDD2.n151 VDD2.n141 171.744
R1463 VDD2.n144 VDD2.n141 171.744
R1464 VDD2.n34 VDD2.n31 171.744
R1465 VDD2.n41 VDD2.n31 171.744
R1466 VDD2.n42 VDD2.n41 171.744
R1467 VDD2.n42 VDD2.n27 171.744
R1468 VDD2.n49 VDD2.n27 171.744
R1469 VDD2.n51 VDD2.n49 171.744
R1470 VDD2.n51 VDD2.n50 171.744
R1471 VDD2.n50 VDD2.n23 171.744
R1472 VDD2.n59 VDD2.n23 171.744
R1473 VDD2.n60 VDD2.n59 171.744
R1474 VDD2.n60 VDD2.n19 171.744
R1475 VDD2.n67 VDD2.n19 171.744
R1476 VDD2.n68 VDD2.n67 171.744
R1477 VDD2.n68 VDD2.n15 171.744
R1478 VDD2.n75 VDD2.n15 171.744
R1479 VDD2.n76 VDD2.n75 171.744
R1480 VDD2.n76 VDD2.n11 171.744
R1481 VDD2.n83 VDD2.n11 171.744
R1482 VDD2.n84 VDD2.n83 171.744
R1483 VDD2.n84 VDD2.n7 171.744
R1484 VDD2.n91 VDD2.n7 171.744
R1485 VDD2.n92 VDD2.n91 171.744
R1486 VDD2.n92 VDD2.n3 171.744
R1487 VDD2.n99 VDD2.n3 171.744
R1488 VDD2.n100 VDD2.n99 171.744
R1489 VDD2.n144 VDD2.t9 85.8723
R1490 VDD2.n34 VDD2.t5 85.8723
R1491 VDD2.n108 VDD2.n107 74.3562
R1492 VDD2 VDD2.n217 74.3533
R1493 VDD2.n216 VDD2.n215 71.722
R1494 VDD2.n106 VDD2.n105 71.7219
R1495 VDD2.n214 VDD2.n108 57.5774
R1496 VDD2.n106 VDD2.n104 56.3291
R1497 VDD2.n214 VDD2.n213 52.7429
R1498 VDD2.n167 VDD2.n166 13.1884
R1499 VDD2.n58 VDD2.n57 13.1884
R1500 VDD2.n211 VDD2.n210 12.8005
R1501 VDD2.n170 VDD2.n131 12.8005
R1502 VDD2.n165 VDD2.n133 12.8005
R1503 VDD2.n56 VDD2.n24 12.8005
R1504 VDD2.n61 VDD2.n22 12.8005
R1505 VDD2.n102 VDD2.n101 12.8005
R1506 VDD2.n207 VDD2.n111 12.0247
R1507 VDD2.n171 VDD2.n129 12.0247
R1508 VDD2.n162 VDD2.n161 12.0247
R1509 VDD2.n53 VDD2.n52 12.0247
R1510 VDD2.n62 VDD2.n20 12.0247
R1511 VDD2.n98 VDD2.n2 12.0247
R1512 VDD2.n206 VDD2.n113 11.249
R1513 VDD2.n175 VDD2.n174 11.249
R1514 VDD2.n158 VDD2.n135 11.249
R1515 VDD2.n48 VDD2.n26 11.249
R1516 VDD2.n66 VDD2.n65 11.249
R1517 VDD2.n97 VDD2.n4 11.249
R1518 VDD2.n145 VDD2.n143 10.7239
R1519 VDD2.n35 VDD2.n33 10.7239
R1520 VDD2.n203 VDD2.n202 10.4732
R1521 VDD2.n178 VDD2.n127 10.4732
R1522 VDD2.n157 VDD2.n138 10.4732
R1523 VDD2.n47 VDD2.n28 10.4732
R1524 VDD2.n69 VDD2.n18 10.4732
R1525 VDD2.n94 VDD2.n93 10.4732
R1526 VDD2.n199 VDD2.n115 9.69747
R1527 VDD2.n179 VDD2.n125 9.69747
R1528 VDD2.n154 VDD2.n153 9.69747
R1529 VDD2.n44 VDD2.n43 9.69747
R1530 VDD2.n70 VDD2.n16 9.69747
R1531 VDD2.n90 VDD2.n6 9.69747
R1532 VDD2.n213 VDD2.n212 9.45567
R1533 VDD2.n104 VDD2.n103 9.45567
R1534 VDD2.n147 VDD2.n146 9.3005
R1535 VDD2.n149 VDD2.n148 9.3005
R1536 VDD2.n140 VDD2.n139 9.3005
R1537 VDD2.n155 VDD2.n154 9.3005
R1538 VDD2.n157 VDD2.n156 9.3005
R1539 VDD2.n135 VDD2.n134 9.3005
R1540 VDD2.n163 VDD2.n162 9.3005
R1541 VDD2.n165 VDD2.n164 9.3005
R1542 VDD2.n119 VDD2.n118 9.3005
R1543 VDD2.n196 VDD2.n195 9.3005
R1544 VDD2.n198 VDD2.n197 9.3005
R1545 VDD2.n115 VDD2.n114 9.3005
R1546 VDD2.n204 VDD2.n203 9.3005
R1547 VDD2.n206 VDD2.n205 9.3005
R1548 VDD2.n111 VDD2.n110 9.3005
R1549 VDD2.n212 VDD2.n211 9.3005
R1550 VDD2.n190 VDD2.n189 9.3005
R1551 VDD2.n188 VDD2.n187 9.3005
R1552 VDD2.n123 VDD2.n122 9.3005
R1553 VDD2.n182 VDD2.n181 9.3005
R1554 VDD2.n180 VDD2.n179 9.3005
R1555 VDD2.n127 VDD2.n126 9.3005
R1556 VDD2.n174 VDD2.n173 9.3005
R1557 VDD2.n172 VDD2.n171 9.3005
R1558 VDD2.n131 VDD2.n130 9.3005
R1559 VDD2.n79 VDD2.n78 9.3005
R1560 VDD2.n14 VDD2.n13 9.3005
R1561 VDD2.n73 VDD2.n72 9.3005
R1562 VDD2.n71 VDD2.n70 9.3005
R1563 VDD2.n18 VDD2.n17 9.3005
R1564 VDD2.n65 VDD2.n64 9.3005
R1565 VDD2.n63 VDD2.n62 9.3005
R1566 VDD2.n22 VDD2.n21 9.3005
R1567 VDD2.n37 VDD2.n36 9.3005
R1568 VDD2.n39 VDD2.n38 9.3005
R1569 VDD2.n30 VDD2.n29 9.3005
R1570 VDD2.n45 VDD2.n44 9.3005
R1571 VDD2.n47 VDD2.n46 9.3005
R1572 VDD2.n26 VDD2.n25 9.3005
R1573 VDD2.n54 VDD2.n53 9.3005
R1574 VDD2.n56 VDD2.n55 9.3005
R1575 VDD2.n81 VDD2.n80 9.3005
R1576 VDD2.n10 VDD2.n9 9.3005
R1577 VDD2.n87 VDD2.n86 9.3005
R1578 VDD2.n89 VDD2.n88 9.3005
R1579 VDD2.n6 VDD2.n5 9.3005
R1580 VDD2.n95 VDD2.n94 9.3005
R1581 VDD2.n97 VDD2.n96 9.3005
R1582 VDD2.n2 VDD2.n1 9.3005
R1583 VDD2.n103 VDD2.n102 9.3005
R1584 VDD2.n198 VDD2.n117 8.92171
R1585 VDD2.n183 VDD2.n182 8.92171
R1586 VDD2.n150 VDD2.n140 8.92171
R1587 VDD2.n40 VDD2.n30 8.92171
R1588 VDD2.n74 VDD2.n73 8.92171
R1589 VDD2.n89 VDD2.n8 8.92171
R1590 VDD2.n195 VDD2.n194 8.14595
R1591 VDD2.n186 VDD2.n123 8.14595
R1592 VDD2.n149 VDD2.n142 8.14595
R1593 VDD2.n39 VDD2.n32 8.14595
R1594 VDD2.n77 VDD2.n14 8.14595
R1595 VDD2.n86 VDD2.n85 8.14595
R1596 VDD2.n213 VDD2.n109 7.75445
R1597 VDD2.n104 VDD2.n0 7.75445
R1598 VDD2.n191 VDD2.n119 7.3702
R1599 VDD2.n187 VDD2.n121 7.3702
R1600 VDD2.n146 VDD2.n145 7.3702
R1601 VDD2.n36 VDD2.n35 7.3702
R1602 VDD2.n78 VDD2.n12 7.3702
R1603 VDD2.n82 VDD2.n10 7.3702
R1604 VDD2.n191 VDD2.n190 6.59444
R1605 VDD2.n190 VDD2.n121 6.59444
R1606 VDD2.n81 VDD2.n12 6.59444
R1607 VDD2.n82 VDD2.n81 6.59444
R1608 VDD2.n211 VDD2.n109 6.08283
R1609 VDD2.n102 VDD2.n0 6.08283
R1610 VDD2.n194 VDD2.n119 5.81868
R1611 VDD2.n187 VDD2.n186 5.81868
R1612 VDD2.n146 VDD2.n142 5.81868
R1613 VDD2.n36 VDD2.n32 5.81868
R1614 VDD2.n78 VDD2.n77 5.81868
R1615 VDD2.n85 VDD2.n10 5.81868
R1616 VDD2.n195 VDD2.n117 5.04292
R1617 VDD2.n183 VDD2.n123 5.04292
R1618 VDD2.n150 VDD2.n149 5.04292
R1619 VDD2.n40 VDD2.n39 5.04292
R1620 VDD2.n74 VDD2.n14 5.04292
R1621 VDD2.n86 VDD2.n8 5.04292
R1622 VDD2.n199 VDD2.n198 4.26717
R1623 VDD2.n182 VDD2.n125 4.26717
R1624 VDD2.n153 VDD2.n140 4.26717
R1625 VDD2.n43 VDD2.n30 4.26717
R1626 VDD2.n73 VDD2.n16 4.26717
R1627 VDD2.n90 VDD2.n89 4.26717
R1628 VDD2.n216 VDD2.n214 3.58671
R1629 VDD2.n202 VDD2.n115 3.49141
R1630 VDD2.n179 VDD2.n178 3.49141
R1631 VDD2.n154 VDD2.n138 3.49141
R1632 VDD2.n44 VDD2.n28 3.49141
R1633 VDD2.n70 VDD2.n69 3.49141
R1634 VDD2.n93 VDD2.n6 3.49141
R1635 VDD2.n203 VDD2.n113 2.71565
R1636 VDD2.n175 VDD2.n127 2.71565
R1637 VDD2.n158 VDD2.n157 2.71565
R1638 VDD2.n48 VDD2.n47 2.71565
R1639 VDD2.n66 VDD2.n18 2.71565
R1640 VDD2.n94 VDD2.n4 2.71565
R1641 VDD2.n147 VDD2.n143 2.41282
R1642 VDD2.n37 VDD2.n33 2.41282
R1643 VDD2.n207 VDD2.n206 1.93989
R1644 VDD2.n174 VDD2.n129 1.93989
R1645 VDD2.n161 VDD2.n135 1.93989
R1646 VDD2.n52 VDD2.n26 1.93989
R1647 VDD2.n65 VDD2.n20 1.93989
R1648 VDD2.n98 VDD2.n97 1.93989
R1649 VDD2.n217 VDD2.t3 1.66572
R1650 VDD2.n217 VDD2.t4 1.66572
R1651 VDD2.n215 VDD2.t8 1.66572
R1652 VDD2.n215 VDD2.t7 1.66572
R1653 VDD2.n107 VDD2.t0 1.66572
R1654 VDD2.n107 VDD2.t2 1.66572
R1655 VDD2.n105 VDD2.t6 1.66572
R1656 VDD2.n105 VDD2.t1 1.66572
R1657 VDD2.n210 VDD2.n111 1.16414
R1658 VDD2.n171 VDD2.n170 1.16414
R1659 VDD2.n162 VDD2.n133 1.16414
R1660 VDD2.n53 VDD2.n24 1.16414
R1661 VDD2.n62 VDD2.n61 1.16414
R1662 VDD2.n101 VDD2.n2 1.16414
R1663 VDD2 VDD2.n216 0.955241
R1664 VDD2.n108 VDD2.n106 0.841706
R1665 VDD2.n167 VDD2.n131 0.388379
R1666 VDD2.n166 VDD2.n165 0.388379
R1667 VDD2.n57 VDD2.n56 0.388379
R1668 VDD2.n58 VDD2.n22 0.388379
R1669 VDD2.n212 VDD2.n110 0.155672
R1670 VDD2.n205 VDD2.n110 0.155672
R1671 VDD2.n205 VDD2.n204 0.155672
R1672 VDD2.n204 VDD2.n114 0.155672
R1673 VDD2.n197 VDD2.n114 0.155672
R1674 VDD2.n197 VDD2.n196 0.155672
R1675 VDD2.n196 VDD2.n118 0.155672
R1676 VDD2.n189 VDD2.n118 0.155672
R1677 VDD2.n189 VDD2.n188 0.155672
R1678 VDD2.n188 VDD2.n122 0.155672
R1679 VDD2.n181 VDD2.n122 0.155672
R1680 VDD2.n181 VDD2.n180 0.155672
R1681 VDD2.n180 VDD2.n126 0.155672
R1682 VDD2.n173 VDD2.n126 0.155672
R1683 VDD2.n173 VDD2.n172 0.155672
R1684 VDD2.n172 VDD2.n130 0.155672
R1685 VDD2.n164 VDD2.n130 0.155672
R1686 VDD2.n164 VDD2.n163 0.155672
R1687 VDD2.n163 VDD2.n134 0.155672
R1688 VDD2.n156 VDD2.n134 0.155672
R1689 VDD2.n156 VDD2.n155 0.155672
R1690 VDD2.n155 VDD2.n139 0.155672
R1691 VDD2.n148 VDD2.n139 0.155672
R1692 VDD2.n148 VDD2.n147 0.155672
R1693 VDD2.n38 VDD2.n37 0.155672
R1694 VDD2.n38 VDD2.n29 0.155672
R1695 VDD2.n45 VDD2.n29 0.155672
R1696 VDD2.n46 VDD2.n45 0.155672
R1697 VDD2.n46 VDD2.n25 0.155672
R1698 VDD2.n54 VDD2.n25 0.155672
R1699 VDD2.n55 VDD2.n54 0.155672
R1700 VDD2.n55 VDD2.n21 0.155672
R1701 VDD2.n63 VDD2.n21 0.155672
R1702 VDD2.n64 VDD2.n63 0.155672
R1703 VDD2.n64 VDD2.n17 0.155672
R1704 VDD2.n71 VDD2.n17 0.155672
R1705 VDD2.n72 VDD2.n71 0.155672
R1706 VDD2.n72 VDD2.n13 0.155672
R1707 VDD2.n79 VDD2.n13 0.155672
R1708 VDD2.n80 VDD2.n79 0.155672
R1709 VDD2.n80 VDD2.n9 0.155672
R1710 VDD2.n87 VDD2.n9 0.155672
R1711 VDD2.n88 VDD2.n87 0.155672
R1712 VDD2.n88 VDD2.n5 0.155672
R1713 VDD2.n95 VDD2.n5 0.155672
R1714 VDD2.n96 VDD2.n95 0.155672
R1715 VDD2.n96 VDD2.n1 0.155672
R1716 VDD2.n103 VDD2.n1 0.155672
R1717 B.n231 B.t7 591.712
R1718 B.n83 B.t11 591.712
R1719 B.n237 B.t4 591.712
R1720 B.n76 B.t2 591.712
R1721 B.n637 B.n198 585
R1722 B.n636 B.n635 585
R1723 B.n634 B.n199 585
R1724 B.n633 B.n632 585
R1725 B.n631 B.n200 585
R1726 B.n630 B.n629 585
R1727 B.n628 B.n201 585
R1728 B.n627 B.n626 585
R1729 B.n625 B.n202 585
R1730 B.n624 B.n623 585
R1731 B.n622 B.n203 585
R1732 B.n621 B.n620 585
R1733 B.n619 B.n204 585
R1734 B.n618 B.n617 585
R1735 B.n616 B.n205 585
R1736 B.n615 B.n614 585
R1737 B.n613 B.n206 585
R1738 B.n612 B.n611 585
R1739 B.n610 B.n207 585
R1740 B.n609 B.n608 585
R1741 B.n607 B.n208 585
R1742 B.n606 B.n605 585
R1743 B.n604 B.n209 585
R1744 B.n603 B.n602 585
R1745 B.n601 B.n210 585
R1746 B.n600 B.n599 585
R1747 B.n598 B.n211 585
R1748 B.n597 B.n596 585
R1749 B.n595 B.n212 585
R1750 B.n594 B.n593 585
R1751 B.n592 B.n213 585
R1752 B.n591 B.n590 585
R1753 B.n589 B.n214 585
R1754 B.n588 B.n587 585
R1755 B.n586 B.n215 585
R1756 B.n585 B.n584 585
R1757 B.n583 B.n216 585
R1758 B.n582 B.n581 585
R1759 B.n580 B.n217 585
R1760 B.n579 B.n578 585
R1761 B.n577 B.n218 585
R1762 B.n576 B.n575 585
R1763 B.n574 B.n219 585
R1764 B.n573 B.n572 585
R1765 B.n571 B.n220 585
R1766 B.n570 B.n569 585
R1767 B.n568 B.n221 585
R1768 B.n567 B.n566 585
R1769 B.n565 B.n222 585
R1770 B.n564 B.n563 585
R1771 B.n562 B.n223 585
R1772 B.n561 B.n560 585
R1773 B.n559 B.n224 585
R1774 B.n558 B.n557 585
R1775 B.n556 B.n225 585
R1776 B.n555 B.n554 585
R1777 B.n553 B.n226 585
R1778 B.n552 B.n551 585
R1779 B.n550 B.n227 585
R1780 B.n549 B.n548 585
R1781 B.n547 B.n228 585
R1782 B.n546 B.n545 585
R1783 B.n544 B.n229 585
R1784 B.n543 B.n542 585
R1785 B.n540 B.n230 585
R1786 B.n539 B.n538 585
R1787 B.n537 B.n233 585
R1788 B.n536 B.n535 585
R1789 B.n534 B.n234 585
R1790 B.n533 B.n532 585
R1791 B.n531 B.n235 585
R1792 B.n530 B.n529 585
R1793 B.n528 B.n236 585
R1794 B.n526 B.n525 585
R1795 B.n524 B.n239 585
R1796 B.n523 B.n522 585
R1797 B.n521 B.n240 585
R1798 B.n520 B.n519 585
R1799 B.n518 B.n241 585
R1800 B.n517 B.n516 585
R1801 B.n515 B.n242 585
R1802 B.n514 B.n513 585
R1803 B.n512 B.n243 585
R1804 B.n511 B.n510 585
R1805 B.n509 B.n244 585
R1806 B.n508 B.n507 585
R1807 B.n506 B.n245 585
R1808 B.n505 B.n504 585
R1809 B.n503 B.n246 585
R1810 B.n502 B.n501 585
R1811 B.n500 B.n247 585
R1812 B.n499 B.n498 585
R1813 B.n497 B.n248 585
R1814 B.n496 B.n495 585
R1815 B.n494 B.n249 585
R1816 B.n493 B.n492 585
R1817 B.n491 B.n250 585
R1818 B.n490 B.n489 585
R1819 B.n488 B.n251 585
R1820 B.n487 B.n486 585
R1821 B.n485 B.n252 585
R1822 B.n484 B.n483 585
R1823 B.n482 B.n253 585
R1824 B.n481 B.n480 585
R1825 B.n479 B.n254 585
R1826 B.n478 B.n477 585
R1827 B.n476 B.n255 585
R1828 B.n475 B.n474 585
R1829 B.n473 B.n256 585
R1830 B.n472 B.n471 585
R1831 B.n470 B.n257 585
R1832 B.n469 B.n468 585
R1833 B.n467 B.n258 585
R1834 B.n466 B.n465 585
R1835 B.n464 B.n259 585
R1836 B.n463 B.n462 585
R1837 B.n461 B.n260 585
R1838 B.n460 B.n459 585
R1839 B.n458 B.n261 585
R1840 B.n457 B.n456 585
R1841 B.n455 B.n262 585
R1842 B.n454 B.n453 585
R1843 B.n452 B.n263 585
R1844 B.n451 B.n450 585
R1845 B.n449 B.n264 585
R1846 B.n448 B.n447 585
R1847 B.n446 B.n265 585
R1848 B.n445 B.n444 585
R1849 B.n443 B.n266 585
R1850 B.n442 B.n441 585
R1851 B.n440 B.n267 585
R1852 B.n439 B.n438 585
R1853 B.n437 B.n268 585
R1854 B.n436 B.n435 585
R1855 B.n434 B.n269 585
R1856 B.n433 B.n432 585
R1857 B.n431 B.n270 585
R1858 B.n639 B.n638 585
R1859 B.n640 B.n197 585
R1860 B.n642 B.n641 585
R1861 B.n643 B.n196 585
R1862 B.n645 B.n644 585
R1863 B.n646 B.n195 585
R1864 B.n648 B.n647 585
R1865 B.n649 B.n194 585
R1866 B.n651 B.n650 585
R1867 B.n652 B.n193 585
R1868 B.n654 B.n653 585
R1869 B.n655 B.n192 585
R1870 B.n657 B.n656 585
R1871 B.n658 B.n191 585
R1872 B.n660 B.n659 585
R1873 B.n661 B.n190 585
R1874 B.n663 B.n662 585
R1875 B.n664 B.n189 585
R1876 B.n666 B.n665 585
R1877 B.n667 B.n188 585
R1878 B.n669 B.n668 585
R1879 B.n670 B.n187 585
R1880 B.n672 B.n671 585
R1881 B.n673 B.n186 585
R1882 B.n675 B.n674 585
R1883 B.n676 B.n185 585
R1884 B.n678 B.n677 585
R1885 B.n679 B.n184 585
R1886 B.n681 B.n680 585
R1887 B.n682 B.n183 585
R1888 B.n684 B.n683 585
R1889 B.n685 B.n182 585
R1890 B.n687 B.n686 585
R1891 B.n688 B.n181 585
R1892 B.n690 B.n689 585
R1893 B.n691 B.n180 585
R1894 B.n693 B.n692 585
R1895 B.n694 B.n179 585
R1896 B.n696 B.n695 585
R1897 B.n697 B.n178 585
R1898 B.n699 B.n698 585
R1899 B.n700 B.n177 585
R1900 B.n702 B.n701 585
R1901 B.n703 B.n176 585
R1902 B.n705 B.n704 585
R1903 B.n706 B.n175 585
R1904 B.n708 B.n707 585
R1905 B.n709 B.n174 585
R1906 B.n711 B.n710 585
R1907 B.n712 B.n173 585
R1908 B.n714 B.n713 585
R1909 B.n715 B.n172 585
R1910 B.n717 B.n716 585
R1911 B.n718 B.n171 585
R1912 B.n720 B.n719 585
R1913 B.n721 B.n170 585
R1914 B.n723 B.n722 585
R1915 B.n724 B.n169 585
R1916 B.n726 B.n725 585
R1917 B.n727 B.n168 585
R1918 B.n729 B.n728 585
R1919 B.n730 B.n167 585
R1920 B.n732 B.n731 585
R1921 B.n733 B.n166 585
R1922 B.n735 B.n734 585
R1923 B.n736 B.n165 585
R1924 B.n738 B.n737 585
R1925 B.n739 B.n164 585
R1926 B.n741 B.n740 585
R1927 B.n742 B.n163 585
R1928 B.n744 B.n743 585
R1929 B.n745 B.n162 585
R1930 B.n747 B.n746 585
R1931 B.n748 B.n161 585
R1932 B.n750 B.n749 585
R1933 B.n751 B.n160 585
R1934 B.n753 B.n752 585
R1935 B.n754 B.n159 585
R1936 B.n756 B.n755 585
R1937 B.n757 B.n158 585
R1938 B.n759 B.n758 585
R1939 B.n760 B.n157 585
R1940 B.n762 B.n761 585
R1941 B.n763 B.n156 585
R1942 B.n765 B.n764 585
R1943 B.n766 B.n155 585
R1944 B.n768 B.n767 585
R1945 B.n769 B.n154 585
R1946 B.n771 B.n770 585
R1947 B.n772 B.n153 585
R1948 B.n774 B.n773 585
R1949 B.n775 B.n152 585
R1950 B.n777 B.n776 585
R1951 B.n778 B.n151 585
R1952 B.n780 B.n779 585
R1953 B.n781 B.n150 585
R1954 B.n783 B.n782 585
R1955 B.n784 B.n149 585
R1956 B.n786 B.n785 585
R1957 B.n787 B.n148 585
R1958 B.n789 B.n788 585
R1959 B.n790 B.n147 585
R1960 B.n792 B.n791 585
R1961 B.n793 B.n146 585
R1962 B.n795 B.n794 585
R1963 B.n796 B.n145 585
R1964 B.n798 B.n797 585
R1965 B.n799 B.n144 585
R1966 B.n801 B.n800 585
R1967 B.n802 B.n143 585
R1968 B.n804 B.n803 585
R1969 B.n805 B.n142 585
R1970 B.n807 B.n806 585
R1971 B.n808 B.n141 585
R1972 B.n810 B.n809 585
R1973 B.n811 B.n140 585
R1974 B.n813 B.n812 585
R1975 B.n814 B.n139 585
R1976 B.n816 B.n815 585
R1977 B.n817 B.n138 585
R1978 B.n819 B.n818 585
R1979 B.n820 B.n137 585
R1980 B.n822 B.n821 585
R1981 B.n823 B.n136 585
R1982 B.n825 B.n824 585
R1983 B.n826 B.n135 585
R1984 B.n828 B.n827 585
R1985 B.n829 B.n134 585
R1986 B.n831 B.n830 585
R1987 B.n832 B.n133 585
R1988 B.n834 B.n833 585
R1989 B.n835 B.n132 585
R1990 B.n837 B.n836 585
R1991 B.n838 B.n131 585
R1992 B.n840 B.n839 585
R1993 B.n841 B.n130 585
R1994 B.n843 B.n842 585
R1995 B.n844 B.n129 585
R1996 B.n846 B.n845 585
R1997 B.n847 B.n128 585
R1998 B.n849 B.n848 585
R1999 B.n850 B.n127 585
R2000 B.n852 B.n851 585
R2001 B.n853 B.n126 585
R2002 B.n855 B.n854 585
R2003 B.n856 B.n125 585
R2004 B.n858 B.n857 585
R2005 B.n859 B.n124 585
R2006 B.n861 B.n860 585
R2007 B.n862 B.n123 585
R2008 B.n864 B.n863 585
R2009 B.n865 B.n122 585
R2010 B.n867 B.n866 585
R2011 B.n868 B.n121 585
R2012 B.n870 B.n869 585
R2013 B.n871 B.n120 585
R2014 B.n873 B.n872 585
R2015 B.n874 B.n119 585
R2016 B.n876 B.n875 585
R2017 B.n877 B.n118 585
R2018 B.n879 B.n878 585
R2019 B.n880 B.n117 585
R2020 B.n882 B.n881 585
R2021 B.n883 B.n116 585
R2022 B.n1090 B.n1089 585
R2023 B.n1088 B.n43 585
R2024 B.n1087 B.n1086 585
R2025 B.n1085 B.n44 585
R2026 B.n1084 B.n1083 585
R2027 B.n1082 B.n45 585
R2028 B.n1081 B.n1080 585
R2029 B.n1079 B.n46 585
R2030 B.n1078 B.n1077 585
R2031 B.n1076 B.n47 585
R2032 B.n1075 B.n1074 585
R2033 B.n1073 B.n48 585
R2034 B.n1072 B.n1071 585
R2035 B.n1070 B.n49 585
R2036 B.n1069 B.n1068 585
R2037 B.n1067 B.n50 585
R2038 B.n1066 B.n1065 585
R2039 B.n1064 B.n51 585
R2040 B.n1063 B.n1062 585
R2041 B.n1061 B.n52 585
R2042 B.n1060 B.n1059 585
R2043 B.n1058 B.n53 585
R2044 B.n1057 B.n1056 585
R2045 B.n1055 B.n54 585
R2046 B.n1054 B.n1053 585
R2047 B.n1052 B.n55 585
R2048 B.n1051 B.n1050 585
R2049 B.n1049 B.n56 585
R2050 B.n1048 B.n1047 585
R2051 B.n1046 B.n57 585
R2052 B.n1045 B.n1044 585
R2053 B.n1043 B.n58 585
R2054 B.n1042 B.n1041 585
R2055 B.n1040 B.n59 585
R2056 B.n1039 B.n1038 585
R2057 B.n1037 B.n60 585
R2058 B.n1036 B.n1035 585
R2059 B.n1034 B.n61 585
R2060 B.n1033 B.n1032 585
R2061 B.n1031 B.n62 585
R2062 B.n1030 B.n1029 585
R2063 B.n1028 B.n63 585
R2064 B.n1027 B.n1026 585
R2065 B.n1025 B.n64 585
R2066 B.n1024 B.n1023 585
R2067 B.n1022 B.n65 585
R2068 B.n1021 B.n1020 585
R2069 B.n1019 B.n66 585
R2070 B.n1018 B.n1017 585
R2071 B.n1016 B.n67 585
R2072 B.n1015 B.n1014 585
R2073 B.n1013 B.n68 585
R2074 B.n1012 B.n1011 585
R2075 B.n1010 B.n69 585
R2076 B.n1009 B.n1008 585
R2077 B.n1007 B.n70 585
R2078 B.n1006 B.n1005 585
R2079 B.n1004 B.n71 585
R2080 B.n1003 B.n1002 585
R2081 B.n1001 B.n72 585
R2082 B.n1000 B.n999 585
R2083 B.n998 B.n73 585
R2084 B.n997 B.n996 585
R2085 B.n995 B.n74 585
R2086 B.n994 B.n993 585
R2087 B.n992 B.n75 585
R2088 B.n991 B.n990 585
R2089 B.n989 B.n79 585
R2090 B.n988 B.n987 585
R2091 B.n986 B.n80 585
R2092 B.n985 B.n984 585
R2093 B.n983 B.n81 585
R2094 B.n982 B.n981 585
R2095 B.n979 B.n82 585
R2096 B.n978 B.n977 585
R2097 B.n976 B.n85 585
R2098 B.n975 B.n974 585
R2099 B.n973 B.n86 585
R2100 B.n972 B.n971 585
R2101 B.n970 B.n87 585
R2102 B.n969 B.n968 585
R2103 B.n967 B.n88 585
R2104 B.n966 B.n965 585
R2105 B.n964 B.n89 585
R2106 B.n963 B.n962 585
R2107 B.n961 B.n90 585
R2108 B.n960 B.n959 585
R2109 B.n958 B.n91 585
R2110 B.n957 B.n956 585
R2111 B.n955 B.n92 585
R2112 B.n954 B.n953 585
R2113 B.n952 B.n93 585
R2114 B.n951 B.n950 585
R2115 B.n949 B.n94 585
R2116 B.n948 B.n947 585
R2117 B.n946 B.n95 585
R2118 B.n945 B.n944 585
R2119 B.n943 B.n96 585
R2120 B.n942 B.n941 585
R2121 B.n940 B.n97 585
R2122 B.n939 B.n938 585
R2123 B.n937 B.n98 585
R2124 B.n936 B.n935 585
R2125 B.n934 B.n99 585
R2126 B.n933 B.n932 585
R2127 B.n931 B.n100 585
R2128 B.n930 B.n929 585
R2129 B.n928 B.n101 585
R2130 B.n927 B.n926 585
R2131 B.n925 B.n102 585
R2132 B.n924 B.n923 585
R2133 B.n922 B.n103 585
R2134 B.n921 B.n920 585
R2135 B.n919 B.n104 585
R2136 B.n918 B.n917 585
R2137 B.n916 B.n105 585
R2138 B.n915 B.n914 585
R2139 B.n913 B.n106 585
R2140 B.n912 B.n911 585
R2141 B.n910 B.n107 585
R2142 B.n909 B.n908 585
R2143 B.n907 B.n108 585
R2144 B.n906 B.n905 585
R2145 B.n904 B.n109 585
R2146 B.n903 B.n902 585
R2147 B.n901 B.n110 585
R2148 B.n900 B.n899 585
R2149 B.n898 B.n111 585
R2150 B.n897 B.n896 585
R2151 B.n895 B.n112 585
R2152 B.n894 B.n893 585
R2153 B.n892 B.n113 585
R2154 B.n891 B.n890 585
R2155 B.n889 B.n114 585
R2156 B.n888 B.n887 585
R2157 B.n886 B.n115 585
R2158 B.n885 B.n884 585
R2159 B.n1091 B.n42 585
R2160 B.n1093 B.n1092 585
R2161 B.n1094 B.n41 585
R2162 B.n1096 B.n1095 585
R2163 B.n1097 B.n40 585
R2164 B.n1099 B.n1098 585
R2165 B.n1100 B.n39 585
R2166 B.n1102 B.n1101 585
R2167 B.n1103 B.n38 585
R2168 B.n1105 B.n1104 585
R2169 B.n1106 B.n37 585
R2170 B.n1108 B.n1107 585
R2171 B.n1109 B.n36 585
R2172 B.n1111 B.n1110 585
R2173 B.n1112 B.n35 585
R2174 B.n1114 B.n1113 585
R2175 B.n1115 B.n34 585
R2176 B.n1117 B.n1116 585
R2177 B.n1118 B.n33 585
R2178 B.n1120 B.n1119 585
R2179 B.n1121 B.n32 585
R2180 B.n1123 B.n1122 585
R2181 B.n1124 B.n31 585
R2182 B.n1126 B.n1125 585
R2183 B.n1127 B.n30 585
R2184 B.n1129 B.n1128 585
R2185 B.n1130 B.n29 585
R2186 B.n1132 B.n1131 585
R2187 B.n1133 B.n28 585
R2188 B.n1135 B.n1134 585
R2189 B.n1136 B.n27 585
R2190 B.n1138 B.n1137 585
R2191 B.n1139 B.n26 585
R2192 B.n1141 B.n1140 585
R2193 B.n1142 B.n25 585
R2194 B.n1144 B.n1143 585
R2195 B.n1145 B.n24 585
R2196 B.n1147 B.n1146 585
R2197 B.n1148 B.n23 585
R2198 B.n1150 B.n1149 585
R2199 B.n1151 B.n22 585
R2200 B.n1153 B.n1152 585
R2201 B.n1154 B.n21 585
R2202 B.n1156 B.n1155 585
R2203 B.n1157 B.n20 585
R2204 B.n1159 B.n1158 585
R2205 B.n1160 B.n19 585
R2206 B.n1162 B.n1161 585
R2207 B.n1163 B.n18 585
R2208 B.n1165 B.n1164 585
R2209 B.n1166 B.n17 585
R2210 B.n1168 B.n1167 585
R2211 B.n1169 B.n16 585
R2212 B.n1171 B.n1170 585
R2213 B.n1172 B.n15 585
R2214 B.n1174 B.n1173 585
R2215 B.n1175 B.n14 585
R2216 B.n1177 B.n1176 585
R2217 B.n1178 B.n13 585
R2218 B.n1180 B.n1179 585
R2219 B.n1181 B.n12 585
R2220 B.n1183 B.n1182 585
R2221 B.n1184 B.n11 585
R2222 B.n1186 B.n1185 585
R2223 B.n1187 B.n10 585
R2224 B.n1189 B.n1188 585
R2225 B.n1190 B.n9 585
R2226 B.n1192 B.n1191 585
R2227 B.n1193 B.n8 585
R2228 B.n1195 B.n1194 585
R2229 B.n1196 B.n7 585
R2230 B.n1198 B.n1197 585
R2231 B.n1199 B.n6 585
R2232 B.n1201 B.n1200 585
R2233 B.n1202 B.n5 585
R2234 B.n1204 B.n1203 585
R2235 B.n1205 B.n4 585
R2236 B.n1207 B.n1206 585
R2237 B.n1208 B.n3 585
R2238 B.n1210 B.n1209 585
R2239 B.n1211 B.n0 585
R2240 B.n2 B.n1 585
R2241 B.n311 B.n310 585
R2242 B.n313 B.n312 585
R2243 B.n314 B.n309 585
R2244 B.n316 B.n315 585
R2245 B.n317 B.n308 585
R2246 B.n319 B.n318 585
R2247 B.n320 B.n307 585
R2248 B.n322 B.n321 585
R2249 B.n323 B.n306 585
R2250 B.n325 B.n324 585
R2251 B.n326 B.n305 585
R2252 B.n328 B.n327 585
R2253 B.n329 B.n304 585
R2254 B.n331 B.n330 585
R2255 B.n332 B.n303 585
R2256 B.n334 B.n333 585
R2257 B.n335 B.n302 585
R2258 B.n337 B.n336 585
R2259 B.n338 B.n301 585
R2260 B.n340 B.n339 585
R2261 B.n341 B.n300 585
R2262 B.n343 B.n342 585
R2263 B.n344 B.n299 585
R2264 B.n346 B.n345 585
R2265 B.n347 B.n298 585
R2266 B.n349 B.n348 585
R2267 B.n350 B.n297 585
R2268 B.n352 B.n351 585
R2269 B.n353 B.n296 585
R2270 B.n355 B.n354 585
R2271 B.n356 B.n295 585
R2272 B.n358 B.n357 585
R2273 B.n359 B.n294 585
R2274 B.n361 B.n360 585
R2275 B.n362 B.n293 585
R2276 B.n364 B.n363 585
R2277 B.n365 B.n292 585
R2278 B.n367 B.n366 585
R2279 B.n368 B.n291 585
R2280 B.n370 B.n369 585
R2281 B.n371 B.n290 585
R2282 B.n373 B.n372 585
R2283 B.n374 B.n289 585
R2284 B.n376 B.n375 585
R2285 B.n377 B.n288 585
R2286 B.n379 B.n378 585
R2287 B.n380 B.n287 585
R2288 B.n382 B.n381 585
R2289 B.n383 B.n286 585
R2290 B.n385 B.n384 585
R2291 B.n386 B.n285 585
R2292 B.n388 B.n387 585
R2293 B.n389 B.n284 585
R2294 B.n391 B.n390 585
R2295 B.n392 B.n283 585
R2296 B.n394 B.n393 585
R2297 B.n395 B.n282 585
R2298 B.n397 B.n396 585
R2299 B.n398 B.n281 585
R2300 B.n400 B.n399 585
R2301 B.n401 B.n280 585
R2302 B.n403 B.n402 585
R2303 B.n404 B.n279 585
R2304 B.n406 B.n405 585
R2305 B.n407 B.n278 585
R2306 B.n409 B.n408 585
R2307 B.n410 B.n277 585
R2308 B.n412 B.n411 585
R2309 B.n413 B.n276 585
R2310 B.n415 B.n414 585
R2311 B.n416 B.n275 585
R2312 B.n418 B.n417 585
R2313 B.n419 B.n274 585
R2314 B.n421 B.n420 585
R2315 B.n422 B.n273 585
R2316 B.n424 B.n423 585
R2317 B.n425 B.n272 585
R2318 B.n427 B.n426 585
R2319 B.n428 B.n271 585
R2320 B.n430 B.n429 585
R2321 B.n232 B.t8 511.034
R2322 B.n84 B.t10 511.034
R2323 B.n238 B.t5 511.034
R2324 B.n77 B.t1 511.034
R2325 B.n429 B.n270 506.916
R2326 B.n639 B.n198 506.916
R2327 B.n885 B.n116 506.916
R2328 B.n1091 B.n1090 506.916
R2329 B.n237 B.t3 332.195
R2330 B.n231 B.t6 332.195
R2331 B.n83 B.t9 332.195
R2332 B.n76 B.t0 332.195
R2333 B.n1213 B.n1212 256.663
R2334 B.n1212 B.n1211 235.042
R2335 B.n1212 B.n2 235.042
R2336 B.n433 B.n270 163.367
R2337 B.n434 B.n433 163.367
R2338 B.n435 B.n434 163.367
R2339 B.n435 B.n268 163.367
R2340 B.n439 B.n268 163.367
R2341 B.n440 B.n439 163.367
R2342 B.n441 B.n440 163.367
R2343 B.n441 B.n266 163.367
R2344 B.n445 B.n266 163.367
R2345 B.n446 B.n445 163.367
R2346 B.n447 B.n446 163.367
R2347 B.n447 B.n264 163.367
R2348 B.n451 B.n264 163.367
R2349 B.n452 B.n451 163.367
R2350 B.n453 B.n452 163.367
R2351 B.n453 B.n262 163.367
R2352 B.n457 B.n262 163.367
R2353 B.n458 B.n457 163.367
R2354 B.n459 B.n458 163.367
R2355 B.n459 B.n260 163.367
R2356 B.n463 B.n260 163.367
R2357 B.n464 B.n463 163.367
R2358 B.n465 B.n464 163.367
R2359 B.n465 B.n258 163.367
R2360 B.n469 B.n258 163.367
R2361 B.n470 B.n469 163.367
R2362 B.n471 B.n470 163.367
R2363 B.n471 B.n256 163.367
R2364 B.n475 B.n256 163.367
R2365 B.n476 B.n475 163.367
R2366 B.n477 B.n476 163.367
R2367 B.n477 B.n254 163.367
R2368 B.n481 B.n254 163.367
R2369 B.n482 B.n481 163.367
R2370 B.n483 B.n482 163.367
R2371 B.n483 B.n252 163.367
R2372 B.n487 B.n252 163.367
R2373 B.n488 B.n487 163.367
R2374 B.n489 B.n488 163.367
R2375 B.n489 B.n250 163.367
R2376 B.n493 B.n250 163.367
R2377 B.n494 B.n493 163.367
R2378 B.n495 B.n494 163.367
R2379 B.n495 B.n248 163.367
R2380 B.n499 B.n248 163.367
R2381 B.n500 B.n499 163.367
R2382 B.n501 B.n500 163.367
R2383 B.n501 B.n246 163.367
R2384 B.n505 B.n246 163.367
R2385 B.n506 B.n505 163.367
R2386 B.n507 B.n506 163.367
R2387 B.n507 B.n244 163.367
R2388 B.n511 B.n244 163.367
R2389 B.n512 B.n511 163.367
R2390 B.n513 B.n512 163.367
R2391 B.n513 B.n242 163.367
R2392 B.n517 B.n242 163.367
R2393 B.n518 B.n517 163.367
R2394 B.n519 B.n518 163.367
R2395 B.n519 B.n240 163.367
R2396 B.n523 B.n240 163.367
R2397 B.n524 B.n523 163.367
R2398 B.n525 B.n524 163.367
R2399 B.n525 B.n236 163.367
R2400 B.n530 B.n236 163.367
R2401 B.n531 B.n530 163.367
R2402 B.n532 B.n531 163.367
R2403 B.n532 B.n234 163.367
R2404 B.n536 B.n234 163.367
R2405 B.n537 B.n536 163.367
R2406 B.n538 B.n537 163.367
R2407 B.n538 B.n230 163.367
R2408 B.n543 B.n230 163.367
R2409 B.n544 B.n543 163.367
R2410 B.n545 B.n544 163.367
R2411 B.n545 B.n228 163.367
R2412 B.n549 B.n228 163.367
R2413 B.n550 B.n549 163.367
R2414 B.n551 B.n550 163.367
R2415 B.n551 B.n226 163.367
R2416 B.n555 B.n226 163.367
R2417 B.n556 B.n555 163.367
R2418 B.n557 B.n556 163.367
R2419 B.n557 B.n224 163.367
R2420 B.n561 B.n224 163.367
R2421 B.n562 B.n561 163.367
R2422 B.n563 B.n562 163.367
R2423 B.n563 B.n222 163.367
R2424 B.n567 B.n222 163.367
R2425 B.n568 B.n567 163.367
R2426 B.n569 B.n568 163.367
R2427 B.n569 B.n220 163.367
R2428 B.n573 B.n220 163.367
R2429 B.n574 B.n573 163.367
R2430 B.n575 B.n574 163.367
R2431 B.n575 B.n218 163.367
R2432 B.n579 B.n218 163.367
R2433 B.n580 B.n579 163.367
R2434 B.n581 B.n580 163.367
R2435 B.n581 B.n216 163.367
R2436 B.n585 B.n216 163.367
R2437 B.n586 B.n585 163.367
R2438 B.n587 B.n586 163.367
R2439 B.n587 B.n214 163.367
R2440 B.n591 B.n214 163.367
R2441 B.n592 B.n591 163.367
R2442 B.n593 B.n592 163.367
R2443 B.n593 B.n212 163.367
R2444 B.n597 B.n212 163.367
R2445 B.n598 B.n597 163.367
R2446 B.n599 B.n598 163.367
R2447 B.n599 B.n210 163.367
R2448 B.n603 B.n210 163.367
R2449 B.n604 B.n603 163.367
R2450 B.n605 B.n604 163.367
R2451 B.n605 B.n208 163.367
R2452 B.n609 B.n208 163.367
R2453 B.n610 B.n609 163.367
R2454 B.n611 B.n610 163.367
R2455 B.n611 B.n206 163.367
R2456 B.n615 B.n206 163.367
R2457 B.n616 B.n615 163.367
R2458 B.n617 B.n616 163.367
R2459 B.n617 B.n204 163.367
R2460 B.n621 B.n204 163.367
R2461 B.n622 B.n621 163.367
R2462 B.n623 B.n622 163.367
R2463 B.n623 B.n202 163.367
R2464 B.n627 B.n202 163.367
R2465 B.n628 B.n627 163.367
R2466 B.n629 B.n628 163.367
R2467 B.n629 B.n200 163.367
R2468 B.n633 B.n200 163.367
R2469 B.n634 B.n633 163.367
R2470 B.n635 B.n634 163.367
R2471 B.n635 B.n198 163.367
R2472 B.n881 B.n116 163.367
R2473 B.n881 B.n880 163.367
R2474 B.n880 B.n879 163.367
R2475 B.n879 B.n118 163.367
R2476 B.n875 B.n118 163.367
R2477 B.n875 B.n874 163.367
R2478 B.n874 B.n873 163.367
R2479 B.n873 B.n120 163.367
R2480 B.n869 B.n120 163.367
R2481 B.n869 B.n868 163.367
R2482 B.n868 B.n867 163.367
R2483 B.n867 B.n122 163.367
R2484 B.n863 B.n122 163.367
R2485 B.n863 B.n862 163.367
R2486 B.n862 B.n861 163.367
R2487 B.n861 B.n124 163.367
R2488 B.n857 B.n124 163.367
R2489 B.n857 B.n856 163.367
R2490 B.n856 B.n855 163.367
R2491 B.n855 B.n126 163.367
R2492 B.n851 B.n126 163.367
R2493 B.n851 B.n850 163.367
R2494 B.n850 B.n849 163.367
R2495 B.n849 B.n128 163.367
R2496 B.n845 B.n128 163.367
R2497 B.n845 B.n844 163.367
R2498 B.n844 B.n843 163.367
R2499 B.n843 B.n130 163.367
R2500 B.n839 B.n130 163.367
R2501 B.n839 B.n838 163.367
R2502 B.n838 B.n837 163.367
R2503 B.n837 B.n132 163.367
R2504 B.n833 B.n132 163.367
R2505 B.n833 B.n832 163.367
R2506 B.n832 B.n831 163.367
R2507 B.n831 B.n134 163.367
R2508 B.n827 B.n134 163.367
R2509 B.n827 B.n826 163.367
R2510 B.n826 B.n825 163.367
R2511 B.n825 B.n136 163.367
R2512 B.n821 B.n136 163.367
R2513 B.n821 B.n820 163.367
R2514 B.n820 B.n819 163.367
R2515 B.n819 B.n138 163.367
R2516 B.n815 B.n138 163.367
R2517 B.n815 B.n814 163.367
R2518 B.n814 B.n813 163.367
R2519 B.n813 B.n140 163.367
R2520 B.n809 B.n140 163.367
R2521 B.n809 B.n808 163.367
R2522 B.n808 B.n807 163.367
R2523 B.n807 B.n142 163.367
R2524 B.n803 B.n142 163.367
R2525 B.n803 B.n802 163.367
R2526 B.n802 B.n801 163.367
R2527 B.n801 B.n144 163.367
R2528 B.n797 B.n144 163.367
R2529 B.n797 B.n796 163.367
R2530 B.n796 B.n795 163.367
R2531 B.n795 B.n146 163.367
R2532 B.n791 B.n146 163.367
R2533 B.n791 B.n790 163.367
R2534 B.n790 B.n789 163.367
R2535 B.n789 B.n148 163.367
R2536 B.n785 B.n148 163.367
R2537 B.n785 B.n784 163.367
R2538 B.n784 B.n783 163.367
R2539 B.n783 B.n150 163.367
R2540 B.n779 B.n150 163.367
R2541 B.n779 B.n778 163.367
R2542 B.n778 B.n777 163.367
R2543 B.n777 B.n152 163.367
R2544 B.n773 B.n152 163.367
R2545 B.n773 B.n772 163.367
R2546 B.n772 B.n771 163.367
R2547 B.n771 B.n154 163.367
R2548 B.n767 B.n154 163.367
R2549 B.n767 B.n766 163.367
R2550 B.n766 B.n765 163.367
R2551 B.n765 B.n156 163.367
R2552 B.n761 B.n156 163.367
R2553 B.n761 B.n760 163.367
R2554 B.n760 B.n759 163.367
R2555 B.n759 B.n158 163.367
R2556 B.n755 B.n158 163.367
R2557 B.n755 B.n754 163.367
R2558 B.n754 B.n753 163.367
R2559 B.n753 B.n160 163.367
R2560 B.n749 B.n160 163.367
R2561 B.n749 B.n748 163.367
R2562 B.n748 B.n747 163.367
R2563 B.n747 B.n162 163.367
R2564 B.n743 B.n162 163.367
R2565 B.n743 B.n742 163.367
R2566 B.n742 B.n741 163.367
R2567 B.n741 B.n164 163.367
R2568 B.n737 B.n164 163.367
R2569 B.n737 B.n736 163.367
R2570 B.n736 B.n735 163.367
R2571 B.n735 B.n166 163.367
R2572 B.n731 B.n166 163.367
R2573 B.n731 B.n730 163.367
R2574 B.n730 B.n729 163.367
R2575 B.n729 B.n168 163.367
R2576 B.n725 B.n168 163.367
R2577 B.n725 B.n724 163.367
R2578 B.n724 B.n723 163.367
R2579 B.n723 B.n170 163.367
R2580 B.n719 B.n170 163.367
R2581 B.n719 B.n718 163.367
R2582 B.n718 B.n717 163.367
R2583 B.n717 B.n172 163.367
R2584 B.n713 B.n172 163.367
R2585 B.n713 B.n712 163.367
R2586 B.n712 B.n711 163.367
R2587 B.n711 B.n174 163.367
R2588 B.n707 B.n174 163.367
R2589 B.n707 B.n706 163.367
R2590 B.n706 B.n705 163.367
R2591 B.n705 B.n176 163.367
R2592 B.n701 B.n176 163.367
R2593 B.n701 B.n700 163.367
R2594 B.n700 B.n699 163.367
R2595 B.n699 B.n178 163.367
R2596 B.n695 B.n178 163.367
R2597 B.n695 B.n694 163.367
R2598 B.n694 B.n693 163.367
R2599 B.n693 B.n180 163.367
R2600 B.n689 B.n180 163.367
R2601 B.n689 B.n688 163.367
R2602 B.n688 B.n687 163.367
R2603 B.n687 B.n182 163.367
R2604 B.n683 B.n182 163.367
R2605 B.n683 B.n682 163.367
R2606 B.n682 B.n681 163.367
R2607 B.n681 B.n184 163.367
R2608 B.n677 B.n184 163.367
R2609 B.n677 B.n676 163.367
R2610 B.n676 B.n675 163.367
R2611 B.n675 B.n186 163.367
R2612 B.n671 B.n186 163.367
R2613 B.n671 B.n670 163.367
R2614 B.n670 B.n669 163.367
R2615 B.n669 B.n188 163.367
R2616 B.n665 B.n188 163.367
R2617 B.n665 B.n664 163.367
R2618 B.n664 B.n663 163.367
R2619 B.n663 B.n190 163.367
R2620 B.n659 B.n190 163.367
R2621 B.n659 B.n658 163.367
R2622 B.n658 B.n657 163.367
R2623 B.n657 B.n192 163.367
R2624 B.n653 B.n192 163.367
R2625 B.n653 B.n652 163.367
R2626 B.n652 B.n651 163.367
R2627 B.n651 B.n194 163.367
R2628 B.n647 B.n194 163.367
R2629 B.n647 B.n646 163.367
R2630 B.n646 B.n645 163.367
R2631 B.n645 B.n196 163.367
R2632 B.n641 B.n196 163.367
R2633 B.n641 B.n640 163.367
R2634 B.n640 B.n639 163.367
R2635 B.n1090 B.n43 163.367
R2636 B.n1086 B.n43 163.367
R2637 B.n1086 B.n1085 163.367
R2638 B.n1085 B.n1084 163.367
R2639 B.n1084 B.n45 163.367
R2640 B.n1080 B.n45 163.367
R2641 B.n1080 B.n1079 163.367
R2642 B.n1079 B.n1078 163.367
R2643 B.n1078 B.n47 163.367
R2644 B.n1074 B.n47 163.367
R2645 B.n1074 B.n1073 163.367
R2646 B.n1073 B.n1072 163.367
R2647 B.n1072 B.n49 163.367
R2648 B.n1068 B.n49 163.367
R2649 B.n1068 B.n1067 163.367
R2650 B.n1067 B.n1066 163.367
R2651 B.n1066 B.n51 163.367
R2652 B.n1062 B.n51 163.367
R2653 B.n1062 B.n1061 163.367
R2654 B.n1061 B.n1060 163.367
R2655 B.n1060 B.n53 163.367
R2656 B.n1056 B.n53 163.367
R2657 B.n1056 B.n1055 163.367
R2658 B.n1055 B.n1054 163.367
R2659 B.n1054 B.n55 163.367
R2660 B.n1050 B.n55 163.367
R2661 B.n1050 B.n1049 163.367
R2662 B.n1049 B.n1048 163.367
R2663 B.n1048 B.n57 163.367
R2664 B.n1044 B.n57 163.367
R2665 B.n1044 B.n1043 163.367
R2666 B.n1043 B.n1042 163.367
R2667 B.n1042 B.n59 163.367
R2668 B.n1038 B.n59 163.367
R2669 B.n1038 B.n1037 163.367
R2670 B.n1037 B.n1036 163.367
R2671 B.n1036 B.n61 163.367
R2672 B.n1032 B.n61 163.367
R2673 B.n1032 B.n1031 163.367
R2674 B.n1031 B.n1030 163.367
R2675 B.n1030 B.n63 163.367
R2676 B.n1026 B.n63 163.367
R2677 B.n1026 B.n1025 163.367
R2678 B.n1025 B.n1024 163.367
R2679 B.n1024 B.n65 163.367
R2680 B.n1020 B.n65 163.367
R2681 B.n1020 B.n1019 163.367
R2682 B.n1019 B.n1018 163.367
R2683 B.n1018 B.n67 163.367
R2684 B.n1014 B.n67 163.367
R2685 B.n1014 B.n1013 163.367
R2686 B.n1013 B.n1012 163.367
R2687 B.n1012 B.n69 163.367
R2688 B.n1008 B.n69 163.367
R2689 B.n1008 B.n1007 163.367
R2690 B.n1007 B.n1006 163.367
R2691 B.n1006 B.n71 163.367
R2692 B.n1002 B.n71 163.367
R2693 B.n1002 B.n1001 163.367
R2694 B.n1001 B.n1000 163.367
R2695 B.n1000 B.n73 163.367
R2696 B.n996 B.n73 163.367
R2697 B.n996 B.n995 163.367
R2698 B.n995 B.n994 163.367
R2699 B.n994 B.n75 163.367
R2700 B.n990 B.n75 163.367
R2701 B.n990 B.n989 163.367
R2702 B.n989 B.n988 163.367
R2703 B.n988 B.n80 163.367
R2704 B.n984 B.n80 163.367
R2705 B.n984 B.n983 163.367
R2706 B.n983 B.n982 163.367
R2707 B.n982 B.n82 163.367
R2708 B.n977 B.n82 163.367
R2709 B.n977 B.n976 163.367
R2710 B.n976 B.n975 163.367
R2711 B.n975 B.n86 163.367
R2712 B.n971 B.n86 163.367
R2713 B.n971 B.n970 163.367
R2714 B.n970 B.n969 163.367
R2715 B.n969 B.n88 163.367
R2716 B.n965 B.n88 163.367
R2717 B.n965 B.n964 163.367
R2718 B.n964 B.n963 163.367
R2719 B.n963 B.n90 163.367
R2720 B.n959 B.n90 163.367
R2721 B.n959 B.n958 163.367
R2722 B.n958 B.n957 163.367
R2723 B.n957 B.n92 163.367
R2724 B.n953 B.n92 163.367
R2725 B.n953 B.n952 163.367
R2726 B.n952 B.n951 163.367
R2727 B.n951 B.n94 163.367
R2728 B.n947 B.n94 163.367
R2729 B.n947 B.n946 163.367
R2730 B.n946 B.n945 163.367
R2731 B.n945 B.n96 163.367
R2732 B.n941 B.n96 163.367
R2733 B.n941 B.n940 163.367
R2734 B.n940 B.n939 163.367
R2735 B.n939 B.n98 163.367
R2736 B.n935 B.n98 163.367
R2737 B.n935 B.n934 163.367
R2738 B.n934 B.n933 163.367
R2739 B.n933 B.n100 163.367
R2740 B.n929 B.n100 163.367
R2741 B.n929 B.n928 163.367
R2742 B.n928 B.n927 163.367
R2743 B.n927 B.n102 163.367
R2744 B.n923 B.n102 163.367
R2745 B.n923 B.n922 163.367
R2746 B.n922 B.n921 163.367
R2747 B.n921 B.n104 163.367
R2748 B.n917 B.n104 163.367
R2749 B.n917 B.n916 163.367
R2750 B.n916 B.n915 163.367
R2751 B.n915 B.n106 163.367
R2752 B.n911 B.n106 163.367
R2753 B.n911 B.n910 163.367
R2754 B.n910 B.n909 163.367
R2755 B.n909 B.n108 163.367
R2756 B.n905 B.n108 163.367
R2757 B.n905 B.n904 163.367
R2758 B.n904 B.n903 163.367
R2759 B.n903 B.n110 163.367
R2760 B.n899 B.n110 163.367
R2761 B.n899 B.n898 163.367
R2762 B.n898 B.n897 163.367
R2763 B.n897 B.n112 163.367
R2764 B.n893 B.n112 163.367
R2765 B.n893 B.n892 163.367
R2766 B.n892 B.n891 163.367
R2767 B.n891 B.n114 163.367
R2768 B.n887 B.n114 163.367
R2769 B.n887 B.n886 163.367
R2770 B.n886 B.n885 163.367
R2771 B.n1092 B.n1091 163.367
R2772 B.n1092 B.n41 163.367
R2773 B.n1096 B.n41 163.367
R2774 B.n1097 B.n1096 163.367
R2775 B.n1098 B.n1097 163.367
R2776 B.n1098 B.n39 163.367
R2777 B.n1102 B.n39 163.367
R2778 B.n1103 B.n1102 163.367
R2779 B.n1104 B.n1103 163.367
R2780 B.n1104 B.n37 163.367
R2781 B.n1108 B.n37 163.367
R2782 B.n1109 B.n1108 163.367
R2783 B.n1110 B.n1109 163.367
R2784 B.n1110 B.n35 163.367
R2785 B.n1114 B.n35 163.367
R2786 B.n1115 B.n1114 163.367
R2787 B.n1116 B.n1115 163.367
R2788 B.n1116 B.n33 163.367
R2789 B.n1120 B.n33 163.367
R2790 B.n1121 B.n1120 163.367
R2791 B.n1122 B.n1121 163.367
R2792 B.n1122 B.n31 163.367
R2793 B.n1126 B.n31 163.367
R2794 B.n1127 B.n1126 163.367
R2795 B.n1128 B.n1127 163.367
R2796 B.n1128 B.n29 163.367
R2797 B.n1132 B.n29 163.367
R2798 B.n1133 B.n1132 163.367
R2799 B.n1134 B.n1133 163.367
R2800 B.n1134 B.n27 163.367
R2801 B.n1138 B.n27 163.367
R2802 B.n1139 B.n1138 163.367
R2803 B.n1140 B.n1139 163.367
R2804 B.n1140 B.n25 163.367
R2805 B.n1144 B.n25 163.367
R2806 B.n1145 B.n1144 163.367
R2807 B.n1146 B.n1145 163.367
R2808 B.n1146 B.n23 163.367
R2809 B.n1150 B.n23 163.367
R2810 B.n1151 B.n1150 163.367
R2811 B.n1152 B.n1151 163.367
R2812 B.n1152 B.n21 163.367
R2813 B.n1156 B.n21 163.367
R2814 B.n1157 B.n1156 163.367
R2815 B.n1158 B.n1157 163.367
R2816 B.n1158 B.n19 163.367
R2817 B.n1162 B.n19 163.367
R2818 B.n1163 B.n1162 163.367
R2819 B.n1164 B.n1163 163.367
R2820 B.n1164 B.n17 163.367
R2821 B.n1168 B.n17 163.367
R2822 B.n1169 B.n1168 163.367
R2823 B.n1170 B.n1169 163.367
R2824 B.n1170 B.n15 163.367
R2825 B.n1174 B.n15 163.367
R2826 B.n1175 B.n1174 163.367
R2827 B.n1176 B.n1175 163.367
R2828 B.n1176 B.n13 163.367
R2829 B.n1180 B.n13 163.367
R2830 B.n1181 B.n1180 163.367
R2831 B.n1182 B.n1181 163.367
R2832 B.n1182 B.n11 163.367
R2833 B.n1186 B.n11 163.367
R2834 B.n1187 B.n1186 163.367
R2835 B.n1188 B.n1187 163.367
R2836 B.n1188 B.n9 163.367
R2837 B.n1192 B.n9 163.367
R2838 B.n1193 B.n1192 163.367
R2839 B.n1194 B.n1193 163.367
R2840 B.n1194 B.n7 163.367
R2841 B.n1198 B.n7 163.367
R2842 B.n1199 B.n1198 163.367
R2843 B.n1200 B.n1199 163.367
R2844 B.n1200 B.n5 163.367
R2845 B.n1204 B.n5 163.367
R2846 B.n1205 B.n1204 163.367
R2847 B.n1206 B.n1205 163.367
R2848 B.n1206 B.n3 163.367
R2849 B.n1210 B.n3 163.367
R2850 B.n1211 B.n1210 163.367
R2851 B.n310 B.n2 163.367
R2852 B.n313 B.n310 163.367
R2853 B.n314 B.n313 163.367
R2854 B.n315 B.n314 163.367
R2855 B.n315 B.n308 163.367
R2856 B.n319 B.n308 163.367
R2857 B.n320 B.n319 163.367
R2858 B.n321 B.n320 163.367
R2859 B.n321 B.n306 163.367
R2860 B.n325 B.n306 163.367
R2861 B.n326 B.n325 163.367
R2862 B.n327 B.n326 163.367
R2863 B.n327 B.n304 163.367
R2864 B.n331 B.n304 163.367
R2865 B.n332 B.n331 163.367
R2866 B.n333 B.n332 163.367
R2867 B.n333 B.n302 163.367
R2868 B.n337 B.n302 163.367
R2869 B.n338 B.n337 163.367
R2870 B.n339 B.n338 163.367
R2871 B.n339 B.n300 163.367
R2872 B.n343 B.n300 163.367
R2873 B.n344 B.n343 163.367
R2874 B.n345 B.n344 163.367
R2875 B.n345 B.n298 163.367
R2876 B.n349 B.n298 163.367
R2877 B.n350 B.n349 163.367
R2878 B.n351 B.n350 163.367
R2879 B.n351 B.n296 163.367
R2880 B.n355 B.n296 163.367
R2881 B.n356 B.n355 163.367
R2882 B.n357 B.n356 163.367
R2883 B.n357 B.n294 163.367
R2884 B.n361 B.n294 163.367
R2885 B.n362 B.n361 163.367
R2886 B.n363 B.n362 163.367
R2887 B.n363 B.n292 163.367
R2888 B.n367 B.n292 163.367
R2889 B.n368 B.n367 163.367
R2890 B.n369 B.n368 163.367
R2891 B.n369 B.n290 163.367
R2892 B.n373 B.n290 163.367
R2893 B.n374 B.n373 163.367
R2894 B.n375 B.n374 163.367
R2895 B.n375 B.n288 163.367
R2896 B.n379 B.n288 163.367
R2897 B.n380 B.n379 163.367
R2898 B.n381 B.n380 163.367
R2899 B.n381 B.n286 163.367
R2900 B.n385 B.n286 163.367
R2901 B.n386 B.n385 163.367
R2902 B.n387 B.n386 163.367
R2903 B.n387 B.n284 163.367
R2904 B.n391 B.n284 163.367
R2905 B.n392 B.n391 163.367
R2906 B.n393 B.n392 163.367
R2907 B.n393 B.n282 163.367
R2908 B.n397 B.n282 163.367
R2909 B.n398 B.n397 163.367
R2910 B.n399 B.n398 163.367
R2911 B.n399 B.n280 163.367
R2912 B.n403 B.n280 163.367
R2913 B.n404 B.n403 163.367
R2914 B.n405 B.n404 163.367
R2915 B.n405 B.n278 163.367
R2916 B.n409 B.n278 163.367
R2917 B.n410 B.n409 163.367
R2918 B.n411 B.n410 163.367
R2919 B.n411 B.n276 163.367
R2920 B.n415 B.n276 163.367
R2921 B.n416 B.n415 163.367
R2922 B.n417 B.n416 163.367
R2923 B.n417 B.n274 163.367
R2924 B.n421 B.n274 163.367
R2925 B.n422 B.n421 163.367
R2926 B.n423 B.n422 163.367
R2927 B.n423 B.n272 163.367
R2928 B.n427 B.n272 163.367
R2929 B.n428 B.n427 163.367
R2930 B.n429 B.n428 163.367
R2931 B.n238 B.n237 80.6793
R2932 B.n232 B.n231 80.6793
R2933 B.n84 B.n83 80.6793
R2934 B.n77 B.n76 80.6793
R2935 B.n527 B.n238 59.5399
R2936 B.n541 B.n232 59.5399
R2937 B.n980 B.n84 59.5399
R2938 B.n78 B.n77 59.5399
R2939 B.n1089 B.n42 32.9371
R2940 B.n884 B.n883 32.9371
R2941 B.n638 B.n637 32.9371
R2942 B.n431 B.n430 32.9371
R2943 B B.n1213 18.0485
R2944 B.n1093 B.n42 10.6151
R2945 B.n1094 B.n1093 10.6151
R2946 B.n1095 B.n1094 10.6151
R2947 B.n1095 B.n40 10.6151
R2948 B.n1099 B.n40 10.6151
R2949 B.n1100 B.n1099 10.6151
R2950 B.n1101 B.n1100 10.6151
R2951 B.n1101 B.n38 10.6151
R2952 B.n1105 B.n38 10.6151
R2953 B.n1106 B.n1105 10.6151
R2954 B.n1107 B.n1106 10.6151
R2955 B.n1107 B.n36 10.6151
R2956 B.n1111 B.n36 10.6151
R2957 B.n1112 B.n1111 10.6151
R2958 B.n1113 B.n1112 10.6151
R2959 B.n1113 B.n34 10.6151
R2960 B.n1117 B.n34 10.6151
R2961 B.n1118 B.n1117 10.6151
R2962 B.n1119 B.n1118 10.6151
R2963 B.n1119 B.n32 10.6151
R2964 B.n1123 B.n32 10.6151
R2965 B.n1124 B.n1123 10.6151
R2966 B.n1125 B.n1124 10.6151
R2967 B.n1125 B.n30 10.6151
R2968 B.n1129 B.n30 10.6151
R2969 B.n1130 B.n1129 10.6151
R2970 B.n1131 B.n1130 10.6151
R2971 B.n1131 B.n28 10.6151
R2972 B.n1135 B.n28 10.6151
R2973 B.n1136 B.n1135 10.6151
R2974 B.n1137 B.n1136 10.6151
R2975 B.n1137 B.n26 10.6151
R2976 B.n1141 B.n26 10.6151
R2977 B.n1142 B.n1141 10.6151
R2978 B.n1143 B.n1142 10.6151
R2979 B.n1143 B.n24 10.6151
R2980 B.n1147 B.n24 10.6151
R2981 B.n1148 B.n1147 10.6151
R2982 B.n1149 B.n1148 10.6151
R2983 B.n1149 B.n22 10.6151
R2984 B.n1153 B.n22 10.6151
R2985 B.n1154 B.n1153 10.6151
R2986 B.n1155 B.n1154 10.6151
R2987 B.n1155 B.n20 10.6151
R2988 B.n1159 B.n20 10.6151
R2989 B.n1160 B.n1159 10.6151
R2990 B.n1161 B.n1160 10.6151
R2991 B.n1161 B.n18 10.6151
R2992 B.n1165 B.n18 10.6151
R2993 B.n1166 B.n1165 10.6151
R2994 B.n1167 B.n1166 10.6151
R2995 B.n1167 B.n16 10.6151
R2996 B.n1171 B.n16 10.6151
R2997 B.n1172 B.n1171 10.6151
R2998 B.n1173 B.n1172 10.6151
R2999 B.n1173 B.n14 10.6151
R3000 B.n1177 B.n14 10.6151
R3001 B.n1178 B.n1177 10.6151
R3002 B.n1179 B.n1178 10.6151
R3003 B.n1179 B.n12 10.6151
R3004 B.n1183 B.n12 10.6151
R3005 B.n1184 B.n1183 10.6151
R3006 B.n1185 B.n1184 10.6151
R3007 B.n1185 B.n10 10.6151
R3008 B.n1189 B.n10 10.6151
R3009 B.n1190 B.n1189 10.6151
R3010 B.n1191 B.n1190 10.6151
R3011 B.n1191 B.n8 10.6151
R3012 B.n1195 B.n8 10.6151
R3013 B.n1196 B.n1195 10.6151
R3014 B.n1197 B.n1196 10.6151
R3015 B.n1197 B.n6 10.6151
R3016 B.n1201 B.n6 10.6151
R3017 B.n1202 B.n1201 10.6151
R3018 B.n1203 B.n1202 10.6151
R3019 B.n1203 B.n4 10.6151
R3020 B.n1207 B.n4 10.6151
R3021 B.n1208 B.n1207 10.6151
R3022 B.n1209 B.n1208 10.6151
R3023 B.n1209 B.n0 10.6151
R3024 B.n1089 B.n1088 10.6151
R3025 B.n1088 B.n1087 10.6151
R3026 B.n1087 B.n44 10.6151
R3027 B.n1083 B.n44 10.6151
R3028 B.n1083 B.n1082 10.6151
R3029 B.n1082 B.n1081 10.6151
R3030 B.n1081 B.n46 10.6151
R3031 B.n1077 B.n46 10.6151
R3032 B.n1077 B.n1076 10.6151
R3033 B.n1076 B.n1075 10.6151
R3034 B.n1075 B.n48 10.6151
R3035 B.n1071 B.n48 10.6151
R3036 B.n1071 B.n1070 10.6151
R3037 B.n1070 B.n1069 10.6151
R3038 B.n1069 B.n50 10.6151
R3039 B.n1065 B.n50 10.6151
R3040 B.n1065 B.n1064 10.6151
R3041 B.n1064 B.n1063 10.6151
R3042 B.n1063 B.n52 10.6151
R3043 B.n1059 B.n52 10.6151
R3044 B.n1059 B.n1058 10.6151
R3045 B.n1058 B.n1057 10.6151
R3046 B.n1057 B.n54 10.6151
R3047 B.n1053 B.n54 10.6151
R3048 B.n1053 B.n1052 10.6151
R3049 B.n1052 B.n1051 10.6151
R3050 B.n1051 B.n56 10.6151
R3051 B.n1047 B.n56 10.6151
R3052 B.n1047 B.n1046 10.6151
R3053 B.n1046 B.n1045 10.6151
R3054 B.n1045 B.n58 10.6151
R3055 B.n1041 B.n58 10.6151
R3056 B.n1041 B.n1040 10.6151
R3057 B.n1040 B.n1039 10.6151
R3058 B.n1039 B.n60 10.6151
R3059 B.n1035 B.n60 10.6151
R3060 B.n1035 B.n1034 10.6151
R3061 B.n1034 B.n1033 10.6151
R3062 B.n1033 B.n62 10.6151
R3063 B.n1029 B.n62 10.6151
R3064 B.n1029 B.n1028 10.6151
R3065 B.n1028 B.n1027 10.6151
R3066 B.n1027 B.n64 10.6151
R3067 B.n1023 B.n64 10.6151
R3068 B.n1023 B.n1022 10.6151
R3069 B.n1022 B.n1021 10.6151
R3070 B.n1021 B.n66 10.6151
R3071 B.n1017 B.n66 10.6151
R3072 B.n1017 B.n1016 10.6151
R3073 B.n1016 B.n1015 10.6151
R3074 B.n1015 B.n68 10.6151
R3075 B.n1011 B.n68 10.6151
R3076 B.n1011 B.n1010 10.6151
R3077 B.n1010 B.n1009 10.6151
R3078 B.n1009 B.n70 10.6151
R3079 B.n1005 B.n70 10.6151
R3080 B.n1005 B.n1004 10.6151
R3081 B.n1004 B.n1003 10.6151
R3082 B.n1003 B.n72 10.6151
R3083 B.n999 B.n72 10.6151
R3084 B.n999 B.n998 10.6151
R3085 B.n998 B.n997 10.6151
R3086 B.n997 B.n74 10.6151
R3087 B.n993 B.n992 10.6151
R3088 B.n992 B.n991 10.6151
R3089 B.n991 B.n79 10.6151
R3090 B.n987 B.n79 10.6151
R3091 B.n987 B.n986 10.6151
R3092 B.n986 B.n985 10.6151
R3093 B.n985 B.n81 10.6151
R3094 B.n981 B.n81 10.6151
R3095 B.n979 B.n978 10.6151
R3096 B.n978 B.n85 10.6151
R3097 B.n974 B.n85 10.6151
R3098 B.n974 B.n973 10.6151
R3099 B.n973 B.n972 10.6151
R3100 B.n972 B.n87 10.6151
R3101 B.n968 B.n87 10.6151
R3102 B.n968 B.n967 10.6151
R3103 B.n967 B.n966 10.6151
R3104 B.n966 B.n89 10.6151
R3105 B.n962 B.n89 10.6151
R3106 B.n962 B.n961 10.6151
R3107 B.n961 B.n960 10.6151
R3108 B.n960 B.n91 10.6151
R3109 B.n956 B.n91 10.6151
R3110 B.n956 B.n955 10.6151
R3111 B.n955 B.n954 10.6151
R3112 B.n954 B.n93 10.6151
R3113 B.n950 B.n93 10.6151
R3114 B.n950 B.n949 10.6151
R3115 B.n949 B.n948 10.6151
R3116 B.n948 B.n95 10.6151
R3117 B.n944 B.n95 10.6151
R3118 B.n944 B.n943 10.6151
R3119 B.n943 B.n942 10.6151
R3120 B.n942 B.n97 10.6151
R3121 B.n938 B.n97 10.6151
R3122 B.n938 B.n937 10.6151
R3123 B.n937 B.n936 10.6151
R3124 B.n936 B.n99 10.6151
R3125 B.n932 B.n99 10.6151
R3126 B.n932 B.n931 10.6151
R3127 B.n931 B.n930 10.6151
R3128 B.n930 B.n101 10.6151
R3129 B.n926 B.n101 10.6151
R3130 B.n926 B.n925 10.6151
R3131 B.n925 B.n924 10.6151
R3132 B.n924 B.n103 10.6151
R3133 B.n920 B.n103 10.6151
R3134 B.n920 B.n919 10.6151
R3135 B.n919 B.n918 10.6151
R3136 B.n918 B.n105 10.6151
R3137 B.n914 B.n105 10.6151
R3138 B.n914 B.n913 10.6151
R3139 B.n913 B.n912 10.6151
R3140 B.n912 B.n107 10.6151
R3141 B.n908 B.n107 10.6151
R3142 B.n908 B.n907 10.6151
R3143 B.n907 B.n906 10.6151
R3144 B.n906 B.n109 10.6151
R3145 B.n902 B.n109 10.6151
R3146 B.n902 B.n901 10.6151
R3147 B.n901 B.n900 10.6151
R3148 B.n900 B.n111 10.6151
R3149 B.n896 B.n111 10.6151
R3150 B.n896 B.n895 10.6151
R3151 B.n895 B.n894 10.6151
R3152 B.n894 B.n113 10.6151
R3153 B.n890 B.n113 10.6151
R3154 B.n890 B.n889 10.6151
R3155 B.n889 B.n888 10.6151
R3156 B.n888 B.n115 10.6151
R3157 B.n884 B.n115 10.6151
R3158 B.n883 B.n882 10.6151
R3159 B.n882 B.n117 10.6151
R3160 B.n878 B.n117 10.6151
R3161 B.n878 B.n877 10.6151
R3162 B.n877 B.n876 10.6151
R3163 B.n876 B.n119 10.6151
R3164 B.n872 B.n119 10.6151
R3165 B.n872 B.n871 10.6151
R3166 B.n871 B.n870 10.6151
R3167 B.n870 B.n121 10.6151
R3168 B.n866 B.n121 10.6151
R3169 B.n866 B.n865 10.6151
R3170 B.n865 B.n864 10.6151
R3171 B.n864 B.n123 10.6151
R3172 B.n860 B.n123 10.6151
R3173 B.n860 B.n859 10.6151
R3174 B.n859 B.n858 10.6151
R3175 B.n858 B.n125 10.6151
R3176 B.n854 B.n125 10.6151
R3177 B.n854 B.n853 10.6151
R3178 B.n853 B.n852 10.6151
R3179 B.n852 B.n127 10.6151
R3180 B.n848 B.n127 10.6151
R3181 B.n848 B.n847 10.6151
R3182 B.n847 B.n846 10.6151
R3183 B.n846 B.n129 10.6151
R3184 B.n842 B.n129 10.6151
R3185 B.n842 B.n841 10.6151
R3186 B.n841 B.n840 10.6151
R3187 B.n840 B.n131 10.6151
R3188 B.n836 B.n131 10.6151
R3189 B.n836 B.n835 10.6151
R3190 B.n835 B.n834 10.6151
R3191 B.n834 B.n133 10.6151
R3192 B.n830 B.n133 10.6151
R3193 B.n830 B.n829 10.6151
R3194 B.n829 B.n828 10.6151
R3195 B.n828 B.n135 10.6151
R3196 B.n824 B.n135 10.6151
R3197 B.n824 B.n823 10.6151
R3198 B.n823 B.n822 10.6151
R3199 B.n822 B.n137 10.6151
R3200 B.n818 B.n137 10.6151
R3201 B.n818 B.n817 10.6151
R3202 B.n817 B.n816 10.6151
R3203 B.n816 B.n139 10.6151
R3204 B.n812 B.n139 10.6151
R3205 B.n812 B.n811 10.6151
R3206 B.n811 B.n810 10.6151
R3207 B.n810 B.n141 10.6151
R3208 B.n806 B.n141 10.6151
R3209 B.n806 B.n805 10.6151
R3210 B.n805 B.n804 10.6151
R3211 B.n804 B.n143 10.6151
R3212 B.n800 B.n143 10.6151
R3213 B.n800 B.n799 10.6151
R3214 B.n799 B.n798 10.6151
R3215 B.n798 B.n145 10.6151
R3216 B.n794 B.n145 10.6151
R3217 B.n794 B.n793 10.6151
R3218 B.n793 B.n792 10.6151
R3219 B.n792 B.n147 10.6151
R3220 B.n788 B.n147 10.6151
R3221 B.n788 B.n787 10.6151
R3222 B.n787 B.n786 10.6151
R3223 B.n786 B.n149 10.6151
R3224 B.n782 B.n149 10.6151
R3225 B.n782 B.n781 10.6151
R3226 B.n781 B.n780 10.6151
R3227 B.n780 B.n151 10.6151
R3228 B.n776 B.n151 10.6151
R3229 B.n776 B.n775 10.6151
R3230 B.n775 B.n774 10.6151
R3231 B.n774 B.n153 10.6151
R3232 B.n770 B.n153 10.6151
R3233 B.n770 B.n769 10.6151
R3234 B.n769 B.n768 10.6151
R3235 B.n768 B.n155 10.6151
R3236 B.n764 B.n155 10.6151
R3237 B.n764 B.n763 10.6151
R3238 B.n763 B.n762 10.6151
R3239 B.n762 B.n157 10.6151
R3240 B.n758 B.n157 10.6151
R3241 B.n758 B.n757 10.6151
R3242 B.n757 B.n756 10.6151
R3243 B.n756 B.n159 10.6151
R3244 B.n752 B.n159 10.6151
R3245 B.n752 B.n751 10.6151
R3246 B.n751 B.n750 10.6151
R3247 B.n750 B.n161 10.6151
R3248 B.n746 B.n161 10.6151
R3249 B.n746 B.n745 10.6151
R3250 B.n745 B.n744 10.6151
R3251 B.n744 B.n163 10.6151
R3252 B.n740 B.n163 10.6151
R3253 B.n740 B.n739 10.6151
R3254 B.n739 B.n738 10.6151
R3255 B.n738 B.n165 10.6151
R3256 B.n734 B.n165 10.6151
R3257 B.n734 B.n733 10.6151
R3258 B.n733 B.n732 10.6151
R3259 B.n732 B.n167 10.6151
R3260 B.n728 B.n167 10.6151
R3261 B.n728 B.n727 10.6151
R3262 B.n727 B.n726 10.6151
R3263 B.n726 B.n169 10.6151
R3264 B.n722 B.n169 10.6151
R3265 B.n722 B.n721 10.6151
R3266 B.n721 B.n720 10.6151
R3267 B.n720 B.n171 10.6151
R3268 B.n716 B.n171 10.6151
R3269 B.n716 B.n715 10.6151
R3270 B.n715 B.n714 10.6151
R3271 B.n714 B.n173 10.6151
R3272 B.n710 B.n173 10.6151
R3273 B.n710 B.n709 10.6151
R3274 B.n709 B.n708 10.6151
R3275 B.n708 B.n175 10.6151
R3276 B.n704 B.n175 10.6151
R3277 B.n704 B.n703 10.6151
R3278 B.n703 B.n702 10.6151
R3279 B.n702 B.n177 10.6151
R3280 B.n698 B.n177 10.6151
R3281 B.n698 B.n697 10.6151
R3282 B.n697 B.n696 10.6151
R3283 B.n696 B.n179 10.6151
R3284 B.n692 B.n179 10.6151
R3285 B.n692 B.n691 10.6151
R3286 B.n691 B.n690 10.6151
R3287 B.n690 B.n181 10.6151
R3288 B.n686 B.n181 10.6151
R3289 B.n686 B.n685 10.6151
R3290 B.n685 B.n684 10.6151
R3291 B.n684 B.n183 10.6151
R3292 B.n680 B.n183 10.6151
R3293 B.n680 B.n679 10.6151
R3294 B.n679 B.n678 10.6151
R3295 B.n678 B.n185 10.6151
R3296 B.n674 B.n185 10.6151
R3297 B.n674 B.n673 10.6151
R3298 B.n673 B.n672 10.6151
R3299 B.n672 B.n187 10.6151
R3300 B.n668 B.n187 10.6151
R3301 B.n668 B.n667 10.6151
R3302 B.n667 B.n666 10.6151
R3303 B.n666 B.n189 10.6151
R3304 B.n662 B.n189 10.6151
R3305 B.n662 B.n661 10.6151
R3306 B.n661 B.n660 10.6151
R3307 B.n660 B.n191 10.6151
R3308 B.n656 B.n191 10.6151
R3309 B.n656 B.n655 10.6151
R3310 B.n655 B.n654 10.6151
R3311 B.n654 B.n193 10.6151
R3312 B.n650 B.n193 10.6151
R3313 B.n650 B.n649 10.6151
R3314 B.n649 B.n648 10.6151
R3315 B.n648 B.n195 10.6151
R3316 B.n644 B.n195 10.6151
R3317 B.n644 B.n643 10.6151
R3318 B.n643 B.n642 10.6151
R3319 B.n642 B.n197 10.6151
R3320 B.n638 B.n197 10.6151
R3321 B.n311 B.n1 10.6151
R3322 B.n312 B.n311 10.6151
R3323 B.n312 B.n309 10.6151
R3324 B.n316 B.n309 10.6151
R3325 B.n317 B.n316 10.6151
R3326 B.n318 B.n317 10.6151
R3327 B.n318 B.n307 10.6151
R3328 B.n322 B.n307 10.6151
R3329 B.n323 B.n322 10.6151
R3330 B.n324 B.n323 10.6151
R3331 B.n324 B.n305 10.6151
R3332 B.n328 B.n305 10.6151
R3333 B.n329 B.n328 10.6151
R3334 B.n330 B.n329 10.6151
R3335 B.n330 B.n303 10.6151
R3336 B.n334 B.n303 10.6151
R3337 B.n335 B.n334 10.6151
R3338 B.n336 B.n335 10.6151
R3339 B.n336 B.n301 10.6151
R3340 B.n340 B.n301 10.6151
R3341 B.n341 B.n340 10.6151
R3342 B.n342 B.n341 10.6151
R3343 B.n342 B.n299 10.6151
R3344 B.n346 B.n299 10.6151
R3345 B.n347 B.n346 10.6151
R3346 B.n348 B.n347 10.6151
R3347 B.n348 B.n297 10.6151
R3348 B.n352 B.n297 10.6151
R3349 B.n353 B.n352 10.6151
R3350 B.n354 B.n353 10.6151
R3351 B.n354 B.n295 10.6151
R3352 B.n358 B.n295 10.6151
R3353 B.n359 B.n358 10.6151
R3354 B.n360 B.n359 10.6151
R3355 B.n360 B.n293 10.6151
R3356 B.n364 B.n293 10.6151
R3357 B.n365 B.n364 10.6151
R3358 B.n366 B.n365 10.6151
R3359 B.n366 B.n291 10.6151
R3360 B.n370 B.n291 10.6151
R3361 B.n371 B.n370 10.6151
R3362 B.n372 B.n371 10.6151
R3363 B.n372 B.n289 10.6151
R3364 B.n376 B.n289 10.6151
R3365 B.n377 B.n376 10.6151
R3366 B.n378 B.n377 10.6151
R3367 B.n378 B.n287 10.6151
R3368 B.n382 B.n287 10.6151
R3369 B.n383 B.n382 10.6151
R3370 B.n384 B.n383 10.6151
R3371 B.n384 B.n285 10.6151
R3372 B.n388 B.n285 10.6151
R3373 B.n389 B.n388 10.6151
R3374 B.n390 B.n389 10.6151
R3375 B.n390 B.n283 10.6151
R3376 B.n394 B.n283 10.6151
R3377 B.n395 B.n394 10.6151
R3378 B.n396 B.n395 10.6151
R3379 B.n396 B.n281 10.6151
R3380 B.n400 B.n281 10.6151
R3381 B.n401 B.n400 10.6151
R3382 B.n402 B.n401 10.6151
R3383 B.n402 B.n279 10.6151
R3384 B.n406 B.n279 10.6151
R3385 B.n407 B.n406 10.6151
R3386 B.n408 B.n407 10.6151
R3387 B.n408 B.n277 10.6151
R3388 B.n412 B.n277 10.6151
R3389 B.n413 B.n412 10.6151
R3390 B.n414 B.n413 10.6151
R3391 B.n414 B.n275 10.6151
R3392 B.n418 B.n275 10.6151
R3393 B.n419 B.n418 10.6151
R3394 B.n420 B.n419 10.6151
R3395 B.n420 B.n273 10.6151
R3396 B.n424 B.n273 10.6151
R3397 B.n425 B.n424 10.6151
R3398 B.n426 B.n425 10.6151
R3399 B.n426 B.n271 10.6151
R3400 B.n430 B.n271 10.6151
R3401 B.n432 B.n431 10.6151
R3402 B.n432 B.n269 10.6151
R3403 B.n436 B.n269 10.6151
R3404 B.n437 B.n436 10.6151
R3405 B.n438 B.n437 10.6151
R3406 B.n438 B.n267 10.6151
R3407 B.n442 B.n267 10.6151
R3408 B.n443 B.n442 10.6151
R3409 B.n444 B.n443 10.6151
R3410 B.n444 B.n265 10.6151
R3411 B.n448 B.n265 10.6151
R3412 B.n449 B.n448 10.6151
R3413 B.n450 B.n449 10.6151
R3414 B.n450 B.n263 10.6151
R3415 B.n454 B.n263 10.6151
R3416 B.n455 B.n454 10.6151
R3417 B.n456 B.n455 10.6151
R3418 B.n456 B.n261 10.6151
R3419 B.n460 B.n261 10.6151
R3420 B.n461 B.n460 10.6151
R3421 B.n462 B.n461 10.6151
R3422 B.n462 B.n259 10.6151
R3423 B.n466 B.n259 10.6151
R3424 B.n467 B.n466 10.6151
R3425 B.n468 B.n467 10.6151
R3426 B.n468 B.n257 10.6151
R3427 B.n472 B.n257 10.6151
R3428 B.n473 B.n472 10.6151
R3429 B.n474 B.n473 10.6151
R3430 B.n474 B.n255 10.6151
R3431 B.n478 B.n255 10.6151
R3432 B.n479 B.n478 10.6151
R3433 B.n480 B.n479 10.6151
R3434 B.n480 B.n253 10.6151
R3435 B.n484 B.n253 10.6151
R3436 B.n485 B.n484 10.6151
R3437 B.n486 B.n485 10.6151
R3438 B.n486 B.n251 10.6151
R3439 B.n490 B.n251 10.6151
R3440 B.n491 B.n490 10.6151
R3441 B.n492 B.n491 10.6151
R3442 B.n492 B.n249 10.6151
R3443 B.n496 B.n249 10.6151
R3444 B.n497 B.n496 10.6151
R3445 B.n498 B.n497 10.6151
R3446 B.n498 B.n247 10.6151
R3447 B.n502 B.n247 10.6151
R3448 B.n503 B.n502 10.6151
R3449 B.n504 B.n503 10.6151
R3450 B.n504 B.n245 10.6151
R3451 B.n508 B.n245 10.6151
R3452 B.n509 B.n508 10.6151
R3453 B.n510 B.n509 10.6151
R3454 B.n510 B.n243 10.6151
R3455 B.n514 B.n243 10.6151
R3456 B.n515 B.n514 10.6151
R3457 B.n516 B.n515 10.6151
R3458 B.n516 B.n241 10.6151
R3459 B.n520 B.n241 10.6151
R3460 B.n521 B.n520 10.6151
R3461 B.n522 B.n521 10.6151
R3462 B.n522 B.n239 10.6151
R3463 B.n526 B.n239 10.6151
R3464 B.n529 B.n528 10.6151
R3465 B.n529 B.n235 10.6151
R3466 B.n533 B.n235 10.6151
R3467 B.n534 B.n533 10.6151
R3468 B.n535 B.n534 10.6151
R3469 B.n535 B.n233 10.6151
R3470 B.n539 B.n233 10.6151
R3471 B.n540 B.n539 10.6151
R3472 B.n542 B.n229 10.6151
R3473 B.n546 B.n229 10.6151
R3474 B.n547 B.n546 10.6151
R3475 B.n548 B.n547 10.6151
R3476 B.n548 B.n227 10.6151
R3477 B.n552 B.n227 10.6151
R3478 B.n553 B.n552 10.6151
R3479 B.n554 B.n553 10.6151
R3480 B.n554 B.n225 10.6151
R3481 B.n558 B.n225 10.6151
R3482 B.n559 B.n558 10.6151
R3483 B.n560 B.n559 10.6151
R3484 B.n560 B.n223 10.6151
R3485 B.n564 B.n223 10.6151
R3486 B.n565 B.n564 10.6151
R3487 B.n566 B.n565 10.6151
R3488 B.n566 B.n221 10.6151
R3489 B.n570 B.n221 10.6151
R3490 B.n571 B.n570 10.6151
R3491 B.n572 B.n571 10.6151
R3492 B.n572 B.n219 10.6151
R3493 B.n576 B.n219 10.6151
R3494 B.n577 B.n576 10.6151
R3495 B.n578 B.n577 10.6151
R3496 B.n578 B.n217 10.6151
R3497 B.n582 B.n217 10.6151
R3498 B.n583 B.n582 10.6151
R3499 B.n584 B.n583 10.6151
R3500 B.n584 B.n215 10.6151
R3501 B.n588 B.n215 10.6151
R3502 B.n589 B.n588 10.6151
R3503 B.n590 B.n589 10.6151
R3504 B.n590 B.n213 10.6151
R3505 B.n594 B.n213 10.6151
R3506 B.n595 B.n594 10.6151
R3507 B.n596 B.n595 10.6151
R3508 B.n596 B.n211 10.6151
R3509 B.n600 B.n211 10.6151
R3510 B.n601 B.n600 10.6151
R3511 B.n602 B.n601 10.6151
R3512 B.n602 B.n209 10.6151
R3513 B.n606 B.n209 10.6151
R3514 B.n607 B.n606 10.6151
R3515 B.n608 B.n607 10.6151
R3516 B.n608 B.n207 10.6151
R3517 B.n612 B.n207 10.6151
R3518 B.n613 B.n612 10.6151
R3519 B.n614 B.n613 10.6151
R3520 B.n614 B.n205 10.6151
R3521 B.n618 B.n205 10.6151
R3522 B.n619 B.n618 10.6151
R3523 B.n620 B.n619 10.6151
R3524 B.n620 B.n203 10.6151
R3525 B.n624 B.n203 10.6151
R3526 B.n625 B.n624 10.6151
R3527 B.n626 B.n625 10.6151
R3528 B.n626 B.n201 10.6151
R3529 B.n630 B.n201 10.6151
R3530 B.n631 B.n630 10.6151
R3531 B.n632 B.n631 10.6151
R3532 B.n632 B.n199 10.6151
R3533 B.n636 B.n199 10.6151
R3534 B.n637 B.n636 10.6151
R3535 B.n1213 B.n0 8.11757
R3536 B.n1213 B.n1 8.11757
R3537 B.n993 B.n78 6.5566
R3538 B.n981 B.n980 6.5566
R3539 B.n528 B.n527 6.5566
R3540 B.n541 B.n540 6.5566
R3541 B.n78 B.n74 4.05904
R3542 B.n980 B.n979 4.05904
R3543 B.n527 B.n526 4.05904
R3544 B.n542 B.n541 4.05904
C0 VDD2 VP 0.74029f
C1 B VDD1 3.56539f
C2 VDD2 VN 18.179699f
C3 VTAIL VP 19.0026f
C4 VDD2 w_n5962_n4872# 3.96958f
C5 VTAIL VN 18.9874f
C6 VDD1 VP 18.7595f
C7 VDD1 VN 0.156403f
C8 w_n5962_n4872# VTAIL 4.39256f
C9 B VP 3.0078f
C10 w_n5962_n4872# VDD1 3.76211f
C11 B VN 1.68937f
C12 VDD2 VTAIL 13.9952f
C13 VDD2 VDD1 2.97566f
C14 w_n5962_n4872# B 14.722899f
C15 VP VN 11.5956f
C16 VDD2 B 3.73121f
C17 VTAIL VDD1 13.9362f
C18 w_n5962_n4872# VP 14.03f
C19 B VTAIL 5.990911f
C20 w_n5962_n4872# VN 13.25f
C21 VDD2 VSUBS 2.73109f
C22 VDD1 VSUBS 2.658582f
C23 VTAIL VSUBS 1.849654f
C24 VN VSUBS 9.97886f
C25 VP VSUBS 6.074316f
C26 B VSUBS 7.525259f
C27 w_n5962_n4872# VSUBS 0.354787p
C28 B.n0 VSUBS 0.006447f
C29 B.n1 VSUBS 0.006447f
C30 B.n2 VSUBS 0.009535f
C31 B.n3 VSUBS 0.007307f
C32 B.n4 VSUBS 0.007307f
C33 B.n5 VSUBS 0.007307f
C34 B.n6 VSUBS 0.007307f
C35 B.n7 VSUBS 0.007307f
C36 B.n8 VSUBS 0.007307f
C37 B.n9 VSUBS 0.007307f
C38 B.n10 VSUBS 0.007307f
C39 B.n11 VSUBS 0.007307f
C40 B.n12 VSUBS 0.007307f
C41 B.n13 VSUBS 0.007307f
C42 B.n14 VSUBS 0.007307f
C43 B.n15 VSUBS 0.007307f
C44 B.n16 VSUBS 0.007307f
C45 B.n17 VSUBS 0.007307f
C46 B.n18 VSUBS 0.007307f
C47 B.n19 VSUBS 0.007307f
C48 B.n20 VSUBS 0.007307f
C49 B.n21 VSUBS 0.007307f
C50 B.n22 VSUBS 0.007307f
C51 B.n23 VSUBS 0.007307f
C52 B.n24 VSUBS 0.007307f
C53 B.n25 VSUBS 0.007307f
C54 B.n26 VSUBS 0.007307f
C55 B.n27 VSUBS 0.007307f
C56 B.n28 VSUBS 0.007307f
C57 B.n29 VSUBS 0.007307f
C58 B.n30 VSUBS 0.007307f
C59 B.n31 VSUBS 0.007307f
C60 B.n32 VSUBS 0.007307f
C61 B.n33 VSUBS 0.007307f
C62 B.n34 VSUBS 0.007307f
C63 B.n35 VSUBS 0.007307f
C64 B.n36 VSUBS 0.007307f
C65 B.n37 VSUBS 0.007307f
C66 B.n38 VSUBS 0.007307f
C67 B.n39 VSUBS 0.007307f
C68 B.n40 VSUBS 0.007307f
C69 B.n41 VSUBS 0.007307f
C70 B.n42 VSUBS 0.016785f
C71 B.n43 VSUBS 0.007307f
C72 B.n44 VSUBS 0.007307f
C73 B.n45 VSUBS 0.007307f
C74 B.n46 VSUBS 0.007307f
C75 B.n47 VSUBS 0.007307f
C76 B.n48 VSUBS 0.007307f
C77 B.n49 VSUBS 0.007307f
C78 B.n50 VSUBS 0.007307f
C79 B.n51 VSUBS 0.007307f
C80 B.n52 VSUBS 0.007307f
C81 B.n53 VSUBS 0.007307f
C82 B.n54 VSUBS 0.007307f
C83 B.n55 VSUBS 0.007307f
C84 B.n56 VSUBS 0.007307f
C85 B.n57 VSUBS 0.007307f
C86 B.n58 VSUBS 0.007307f
C87 B.n59 VSUBS 0.007307f
C88 B.n60 VSUBS 0.007307f
C89 B.n61 VSUBS 0.007307f
C90 B.n62 VSUBS 0.007307f
C91 B.n63 VSUBS 0.007307f
C92 B.n64 VSUBS 0.007307f
C93 B.n65 VSUBS 0.007307f
C94 B.n66 VSUBS 0.007307f
C95 B.n67 VSUBS 0.007307f
C96 B.n68 VSUBS 0.007307f
C97 B.n69 VSUBS 0.007307f
C98 B.n70 VSUBS 0.007307f
C99 B.n71 VSUBS 0.007307f
C100 B.n72 VSUBS 0.007307f
C101 B.n73 VSUBS 0.007307f
C102 B.n74 VSUBS 0.00505f
C103 B.n75 VSUBS 0.007307f
C104 B.t1 VSUBS 0.405038f
C105 B.t2 VSUBS 0.453688f
C106 B.t0 VSUBS 3.53993f
C107 B.n76 VSUBS 0.72865f
C108 B.n77 VSUBS 0.367234f
C109 B.n78 VSUBS 0.016929f
C110 B.n79 VSUBS 0.007307f
C111 B.n80 VSUBS 0.007307f
C112 B.n81 VSUBS 0.007307f
C113 B.n82 VSUBS 0.007307f
C114 B.t10 VSUBS 0.405041f
C115 B.t11 VSUBS 0.453691f
C116 B.t9 VSUBS 3.53993f
C117 B.n83 VSUBS 0.728646f
C118 B.n84 VSUBS 0.36723f
C119 B.n85 VSUBS 0.007307f
C120 B.n86 VSUBS 0.007307f
C121 B.n87 VSUBS 0.007307f
C122 B.n88 VSUBS 0.007307f
C123 B.n89 VSUBS 0.007307f
C124 B.n90 VSUBS 0.007307f
C125 B.n91 VSUBS 0.007307f
C126 B.n92 VSUBS 0.007307f
C127 B.n93 VSUBS 0.007307f
C128 B.n94 VSUBS 0.007307f
C129 B.n95 VSUBS 0.007307f
C130 B.n96 VSUBS 0.007307f
C131 B.n97 VSUBS 0.007307f
C132 B.n98 VSUBS 0.007307f
C133 B.n99 VSUBS 0.007307f
C134 B.n100 VSUBS 0.007307f
C135 B.n101 VSUBS 0.007307f
C136 B.n102 VSUBS 0.007307f
C137 B.n103 VSUBS 0.007307f
C138 B.n104 VSUBS 0.007307f
C139 B.n105 VSUBS 0.007307f
C140 B.n106 VSUBS 0.007307f
C141 B.n107 VSUBS 0.007307f
C142 B.n108 VSUBS 0.007307f
C143 B.n109 VSUBS 0.007307f
C144 B.n110 VSUBS 0.007307f
C145 B.n111 VSUBS 0.007307f
C146 B.n112 VSUBS 0.007307f
C147 B.n113 VSUBS 0.007307f
C148 B.n114 VSUBS 0.007307f
C149 B.n115 VSUBS 0.007307f
C150 B.n116 VSUBS 0.016785f
C151 B.n117 VSUBS 0.007307f
C152 B.n118 VSUBS 0.007307f
C153 B.n119 VSUBS 0.007307f
C154 B.n120 VSUBS 0.007307f
C155 B.n121 VSUBS 0.007307f
C156 B.n122 VSUBS 0.007307f
C157 B.n123 VSUBS 0.007307f
C158 B.n124 VSUBS 0.007307f
C159 B.n125 VSUBS 0.007307f
C160 B.n126 VSUBS 0.007307f
C161 B.n127 VSUBS 0.007307f
C162 B.n128 VSUBS 0.007307f
C163 B.n129 VSUBS 0.007307f
C164 B.n130 VSUBS 0.007307f
C165 B.n131 VSUBS 0.007307f
C166 B.n132 VSUBS 0.007307f
C167 B.n133 VSUBS 0.007307f
C168 B.n134 VSUBS 0.007307f
C169 B.n135 VSUBS 0.007307f
C170 B.n136 VSUBS 0.007307f
C171 B.n137 VSUBS 0.007307f
C172 B.n138 VSUBS 0.007307f
C173 B.n139 VSUBS 0.007307f
C174 B.n140 VSUBS 0.007307f
C175 B.n141 VSUBS 0.007307f
C176 B.n142 VSUBS 0.007307f
C177 B.n143 VSUBS 0.007307f
C178 B.n144 VSUBS 0.007307f
C179 B.n145 VSUBS 0.007307f
C180 B.n146 VSUBS 0.007307f
C181 B.n147 VSUBS 0.007307f
C182 B.n148 VSUBS 0.007307f
C183 B.n149 VSUBS 0.007307f
C184 B.n150 VSUBS 0.007307f
C185 B.n151 VSUBS 0.007307f
C186 B.n152 VSUBS 0.007307f
C187 B.n153 VSUBS 0.007307f
C188 B.n154 VSUBS 0.007307f
C189 B.n155 VSUBS 0.007307f
C190 B.n156 VSUBS 0.007307f
C191 B.n157 VSUBS 0.007307f
C192 B.n158 VSUBS 0.007307f
C193 B.n159 VSUBS 0.007307f
C194 B.n160 VSUBS 0.007307f
C195 B.n161 VSUBS 0.007307f
C196 B.n162 VSUBS 0.007307f
C197 B.n163 VSUBS 0.007307f
C198 B.n164 VSUBS 0.007307f
C199 B.n165 VSUBS 0.007307f
C200 B.n166 VSUBS 0.007307f
C201 B.n167 VSUBS 0.007307f
C202 B.n168 VSUBS 0.007307f
C203 B.n169 VSUBS 0.007307f
C204 B.n170 VSUBS 0.007307f
C205 B.n171 VSUBS 0.007307f
C206 B.n172 VSUBS 0.007307f
C207 B.n173 VSUBS 0.007307f
C208 B.n174 VSUBS 0.007307f
C209 B.n175 VSUBS 0.007307f
C210 B.n176 VSUBS 0.007307f
C211 B.n177 VSUBS 0.007307f
C212 B.n178 VSUBS 0.007307f
C213 B.n179 VSUBS 0.007307f
C214 B.n180 VSUBS 0.007307f
C215 B.n181 VSUBS 0.007307f
C216 B.n182 VSUBS 0.007307f
C217 B.n183 VSUBS 0.007307f
C218 B.n184 VSUBS 0.007307f
C219 B.n185 VSUBS 0.007307f
C220 B.n186 VSUBS 0.007307f
C221 B.n187 VSUBS 0.007307f
C222 B.n188 VSUBS 0.007307f
C223 B.n189 VSUBS 0.007307f
C224 B.n190 VSUBS 0.007307f
C225 B.n191 VSUBS 0.007307f
C226 B.n192 VSUBS 0.007307f
C227 B.n193 VSUBS 0.007307f
C228 B.n194 VSUBS 0.007307f
C229 B.n195 VSUBS 0.007307f
C230 B.n196 VSUBS 0.007307f
C231 B.n197 VSUBS 0.007307f
C232 B.n198 VSUBS 0.0176f
C233 B.n199 VSUBS 0.007307f
C234 B.n200 VSUBS 0.007307f
C235 B.n201 VSUBS 0.007307f
C236 B.n202 VSUBS 0.007307f
C237 B.n203 VSUBS 0.007307f
C238 B.n204 VSUBS 0.007307f
C239 B.n205 VSUBS 0.007307f
C240 B.n206 VSUBS 0.007307f
C241 B.n207 VSUBS 0.007307f
C242 B.n208 VSUBS 0.007307f
C243 B.n209 VSUBS 0.007307f
C244 B.n210 VSUBS 0.007307f
C245 B.n211 VSUBS 0.007307f
C246 B.n212 VSUBS 0.007307f
C247 B.n213 VSUBS 0.007307f
C248 B.n214 VSUBS 0.007307f
C249 B.n215 VSUBS 0.007307f
C250 B.n216 VSUBS 0.007307f
C251 B.n217 VSUBS 0.007307f
C252 B.n218 VSUBS 0.007307f
C253 B.n219 VSUBS 0.007307f
C254 B.n220 VSUBS 0.007307f
C255 B.n221 VSUBS 0.007307f
C256 B.n222 VSUBS 0.007307f
C257 B.n223 VSUBS 0.007307f
C258 B.n224 VSUBS 0.007307f
C259 B.n225 VSUBS 0.007307f
C260 B.n226 VSUBS 0.007307f
C261 B.n227 VSUBS 0.007307f
C262 B.n228 VSUBS 0.007307f
C263 B.n229 VSUBS 0.007307f
C264 B.n230 VSUBS 0.007307f
C265 B.t8 VSUBS 0.405041f
C266 B.t7 VSUBS 0.453691f
C267 B.t6 VSUBS 3.53993f
C268 B.n231 VSUBS 0.728646f
C269 B.n232 VSUBS 0.36723f
C270 B.n233 VSUBS 0.007307f
C271 B.n234 VSUBS 0.007307f
C272 B.n235 VSUBS 0.007307f
C273 B.n236 VSUBS 0.007307f
C274 B.t5 VSUBS 0.405038f
C275 B.t4 VSUBS 0.453688f
C276 B.t3 VSUBS 3.53993f
C277 B.n237 VSUBS 0.72865f
C278 B.n238 VSUBS 0.367234f
C279 B.n239 VSUBS 0.007307f
C280 B.n240 VSUBS 0.007307f
C281 B.n241 VSUBS 0.007307f
C282 B.n242 VSUBS 0.007307f
C283 B.n243 VSUBS 0.007307f
C284 B.n244 VSUBS 0.007307f
C285 B.n245 VSUBS 0.007307f
C286 B.n246 VSUBS 0.007307f
C287 B.n247 VSUBS 0.007307f
C288 B.n248 VSUBS 0.007307f
C289 B.n249 VSUBS 0.007307f
C290 B.n250 VSUBS 0.007307f
C291 B.n251 VSUBS 0.007307f
C292 B.n252 VSUBS 0.007307f
C293 B.n253 VSUBS 0.007307f
C294 B.n254 VSUBS 0.007307f
C295 B.n255 VSUBS 0.007307f
C296 B.n256 VSUBS 0.007307f
C297 B.n257 VSUBS 0.007307f
C298 B.n258 VSUBS 0.007307f
C299 B.n259 VSUBS 0.007307f
C300 B.n260 VSUBS 0.007307f
C301 B.n261 VSUBS 0.007307f
C302 B.n262 VSUBS 0.007307f
C303 B.n263 VSUBS 0.007307f
C304 B.n264 VSUBS 0.007307f
C305 B.n265 VSUBS 0.007307f
C306 B.n266 VSUBS 0.007307f
C307 B.n267 VSUBS 0.007307f
C308 B.n268 VSUBS 0.007307f
C309 B.n269 VSUBS 0.007307f
C310 B.n270 VSUBS 0.0176f
C311 B.n271 VSUBS 0.007307f
C312 B.n272 VSUBS 0.007307f
C313 B.n273 VSUBS 0.007307f
C314 B.n274 VSUBS 0.007307f
C315 B.n275 VSUBS 0.007307f
C316 B.n276 VSUBS 0.007307f
C317 B.n277 VSUBS 0.007307f
C318 B.n278 VSUBS 0.007307f
C319 B.n279 VSUBS 0.007307f
C320 B.n280 VSUBS 0.007307f
C321 B.n281 VSUBS 0.007307f
C322 B.n282 VSUBS 0.007307f
C323 B.n283 VSUBS 0.007307f
C324 B.n284 VSUBS 0.007307f
C325 B.n285 VSUBS 0.007307f
C326 B.n286 VSUBS 0.007307f
C327 B.n287 VSUBS 0.007307f
C328 B.n288 VSUBS 0.007307f
C329 B.n289 VSUBS 0.007307f
C330 B.n290 VSUBS 0.007307f
C331 B.n291 VSUBS 0.007307f
C332 B.n292 VSUBS 0.007307f
C333 B.n293 VSUBS 0.007307f
C334 B.n294 VSUBS 0.007307f
C335 B.n295 VSUBS 0.007307f
C336 B.n296 VSUBS 0.007307f
C337 B.n297 VSUBS 0.007307f
C338 B.n298 VSUBS 0.007307f
C339 B.n299 VSUBS 0.007307f
C340 B.n300 VSUBS 0.007307f
C341 B.n301 VSUBS 0.007307f
C342 B.n302 VSUBS 0.007307f
C343 B.n303 VSUBS 0.007307f
C344 B.n304 VSUBS 0.007307f
C345 B.n305 VSUBS 0.007307f
C346 B.n306 VSUBS 0.007307f
C347 B.n307 VSUBS 0.007307f
C348 B.n308 VSUBS 0.007307f
C349 B.n309 VSUBS 0.007307f
C350 B.n310 VSUBS 0.007307f
C351 B.n311 VSUBS 0.007307f
C352 B.n312 VSUBS 0.007307f
C353 B.n313 VSUBS 0.007307f
C354 B.n314 VSUBS 0.007307f
C355 B.n315 VSUBS 0.007307f
C356 B.n316 VSUBS 0.007307f
C357 B.n317 VSUBS 0.007307f
C358 B.n318 VSUBS 0.007307f
C359 B.n319 VSUBS 0.007307f
C360 B.n320 VSUBS 0.007307f
C361 B.n321 VSUBS 0.007307f
C362 B.n322 VSUBS 0.007307f
C363 B.n323 VSUBS 0.007307f
C364 B.n324 VSUBS 0.007307f
C365 B.n325 VSUBS 0.007307f
C366 B.n326 VSUBS 0.007307f
C367 B.n327 VSUBS 0.007307f
C368 B.n328 VSUBS 0.007307f
C369 B.n329 VSUBS 0.007307f
C370 B.n330 VSUBS 0.007307f
C371 B.n331 VSUBS 0.007307f
C372 B.n332 VSUBS 0.007307f
C373 B.n333 VSUBS 0.007307f
C374 B.n334 VSUBS 0.007307f
C375 B.n335 VSUBS 0.007307f
C376 B.n336 VSUBS 0.007307f
C377 B.n337 VSUBS 0.007307f
C378 B.n338 VSUBS 0.007307f
C379 B.n339 VSUBS 0.007307f
C380 B.n340 VSUBS 0.007307f
C381 B.n341 VSUBS 0.007307f
C382 B.n342 VSUBS 0.007307f
C383 B.n343 VSUBS 0.007307f
C384 B.n344 VSUBS 0.007307f
C385 B.n345 VSUBS 0.007307f
C386 B.n346 VSUBS 0.007307f
C387 B.n347 VSUBS 0.007307f
C388 B.n348 VSUBS 0.007307f
C389 B.n349 VSUBS 0.007307f
C390 B.n350 VSUBS 0.007307f
C391 B.n351 VSUBS 0.007307f
C392 B.n352 VSUBS 0.007307f
C393 B.n353 VSUBS 0.007307f
C394 B.n354 VSUBS 0.007307f
C395 B.n355 VSUBS 0.007307f
C396 B.n356 VSUBS 0.007307f
C397 B.n357 VSUBS 0.007307f
C398 B.n358 VSUBS 0.007307f
C399 B.n359 VSUBS 0.007307f
C400 B.n360 VSUBS 0.007307f
C401 B.n361 VSUBS 0.007307f
C402 B.n362 VSUBS 0.007307f
C403 B.n363 VSUBS 0.007307f
C404 B.n364 VSUBS 0.007307f
C405 B.n365 VSUBS 0.007307f
C406 B.n366 VSUBS 0.007307f
C407 B.n367 VSUBS 0.007307f
C408 B.n368 VSUBS 0.007307f
C409 B.n369 VSUBS 0.007307f
C410 B.n370 VSUBS 0.007307f
C411 B.n371 VSUBS 0.007307f
C412 B.n372 VSUBS 0.007307f
C413 B.n373 VSUBS 0.007307f
C414 B.n374 VSUBS 0.007307f
C415 B.n375 VSUBS 0.007307f
C416 B.n376 VSUBS 0.007307f
C417 B.n377 VSUBS 0.007307f
C418 B.n378 VSUBS 0.007307f
C419 B.n379 VSUBS 0.007307f
C420 B.n380 VSUBS 0.007307f
C421 B.n381 VSUBS 0.007307f
C422 B.n382 VSUBS 0.007307f
C423 B.n383 VSUBS 0.007307f
C424 B.n384 VSUBS 0.007307f
C425 B.n385 VSUBS 0.007307f
C426 B.n386 VSUBS 0.007307f
C427 B.n387 VSUBS 0.007307f
C428 B.n388 VSUBS 0.007307f
C429 B.n389 VSUBS 0.007307f
C430 B.n390 VSUBS 0.007307f
C431 B.n391 VSUBS 0.007307f
C432 B.n392 VSUBS 0.007307f
C433 B.n393 VSUBS 0.007307f
C434 B.n394 VSUBS 0.007307f
C435 B.n395 VSUBS 0.007307f
C436 B.n396 VSUBS 0.007307f
C437 B.n397 VSUBS 0.007307f
C438 B.n398 VSUBS 0.007307f
C439 B.n399 VSUBS 0.007307f
C440 B.n400 VSUBS 0.007307f
C441 B.n401 VSUBS 0.007307f
C442 B.n402 VSUBS 0.007307f
C443 B.n403 VSUBS 0.007307f
C444 B.n404 VSUBS 0.007307f
C445 B.n405 VSUBS 0.007307f
C446 B.n406 VSUBS 0.007307f
C447 B.n407 VSUBS 0.007307f
C448 B.n408 VSUBS 0.007307f
C449 B.n409 VSUBS 0.007307f
C450 B.n410 VSUBS 0.007307f
C451 B.n411 VSUBS 0.007307f
C452 B.n412 VSUBS 0.007307f
C453 B.n413 VSUBS 0.007307f
C454 B.n414 VSUBS 0.007307f
C455 B.n415 VSUBS 0.007307f
C456 B.n416 VSUBS 0.007307f
C457 B.n417 VSUBS 0.007307f
C458 B.n418 VSUBS 0.007307f
C459 B.n419 VSUBS 0.007307f
C460 B.n420 VSUBS 0.007307f
C461 B.n421 VSUBS 0.007307f
C462 B.n422 VSUBS 0.007307f
C463 B.n423 VSUBS 0.007307f
C464 B.n424 VSUBS 0.007307f
C465 B.n425 VSUBS 0.007307f
C466 B.n426 VSUBS 0.007307f
C467 B.n427 VSUBS 0.007307f
C468 B.n428 VSUBS 0.007307f
C469 B.n429 VSUBS 0.016785f
C470 B.n430 VSUBS 0.016785f
C471 B.n431 VSUBS 0.0176f
C472 B.n432 VSUBS 0.007307f
C473 B.n433 VSUBS 0.007307f
C474 B.n434 VSUBS 0.007307f
C475 B.n435 VSUBS 0.007307f
C476 B.n436 VSUBS 0.007307f
C477 B.n437 VSUBS 0.007307f
C478 B.n438 VSUBS 0.007307f
C479 B.n439 VSUBS 0.007307f
C480 B.n440 VSUBS 0.007307f
C481 B.n441 VSUBS 0.007307f
C482 B.n442 VSUBS 0.007307f
C483 B.n443 VSUBS 0.007307f
C484 B.n444 VSUBS 0.007307f
C485 B.n445 VSUBS 0.007307f
C486 B.n446 VSUBS 0.007307f
C487 B.n447 VSUBS 0.007307f
C488 B.n448 VSUBS 0.007307f
C489 B.n449 VSUBS 0.007307f
C490 B.n450 VSUBS 0.007307f
C491 B.n451 VSUBS 0.007307f
C492 B.n452 VSUBS 0.007307f
C493 B.n453 VSUBS 0.007307f
C494 B.n454 VSUBS 0.007307f
C495 B.n455 VSUBS 0.007307f
C496 B.n456 VSUBS 0.007307f
C497 B.n457 VSUBS 0.007307f
C498 B.n458 VSUBS 0.007307f
C499 B.n459 VSUBS 0.007307f
C500 B.n460 VSUBS 0.007307f
C501 B.n461 VSUBS 0.007307f
C502 B.n462 VSUBS 0.007307f
C503 B.n463 VSUBS 0.007307f
C504 B.n464 VSUBS 0.007307f
C505 B.n465 VSUBS 0.007307f
C506 B.n466 VSUBS 0.007307f
C507 B.n467 VSUBS 0.007307f
C508 B.n468 VSUBS 0.007307f
C509 B.n469 VSUBS 0.007307f
C510 B.n470 VSUBS 0.007307f
C511 B.n471 VSUBS 0.007307f
C512 B.n472 VSUBS 0.007307f
C513 B.n473 VSUBS 0.007307f
C514 B.n474 VSUBS 0.007307f
C515 B.n475 VSUBS 0.007307f
C516 B.n476 VSUBS 0.007307f
C517 B.n477 VSUBS 0.007307f
C518 B.n478 VSUBS 0.007307f
C519 B.n479 VSUBS 0.007307f
C520 B.n480 VSUBS 0.007307f
C521 B.n481 VSUBS 0.007307f
C522 B.n482 VSUBS 0.007307f
C523 B.n483 VSUBS 0.007307f
C524 B.n484 VSUBS 0.007307f
C525 B.n485 VSUBS 0.007307f
C526 B.n486 VSUBS 0.007307f
C527 B.n487 VSUBS 0.007307f
C528 B.n488 VSUBS 0.007307f
C529 B.n489 VSUBS 0.007307f
C530 B.n490 VSUBS 0.007307f
C531 B.n491 VSUBS 0.007307f
C532 B.n492 VSUBS 0.007307f
C533 B.n493 VSUBS 0.007307f
C534 B.n494 VSUBS 0.007307f
C535 B.n495 VSUBS 0.007307f
C536 B.n496 VSUBS 0.007307f
C537 B.n497 VSUBS 0.007307f
C538 B.n498 VSUBS 0.007307f
C539 B.n499 VSUBS 0.007307f
C540 B.n500 VSUBS 0.007307f
C541 B.n501 VSUBS 0.007307f
C542 B.n502 VSUBS 0.007307f
C543 B.n503 VSUBS 0.007307f
C544 B.n504 VSUBS 0.007307f
C545 B.n505 VSUBS 0.007307f
C546 B.n506 VSUBS 0.007307f
C547 B.n507 VSUBS 0.007307f
C548 B.n508 VSUBS 0.007307f
C549 B.n509 VSUBS 0.007307f
C550 B.n510 VSUBS 0.007307f
C551 B.n511 VSUBS 0.007307f
C552 B.n512 VSUBS 0.007307f
C553 B.n513 VSUBS 0.007307f
C554 B.n514 VSUBS 0.007307f
C555 B.n515 VSUBS 0.007307f
C556 B.n516 VSUBS 0.007307f
C557 B.n517 VSUBS 0.007307f
C558 B.n518 VSUBS 0.007307f
C559 B.n519 VSUBS 0.007307f
C560 B.n520 VSUBS 0.007307f
C561 B.n521 VSUBS 0.007307f
C562 B.n522 VSUBS 0.007307f
C563 B.n523 VSUBS 0.007307f
C564 B.n524 VSUBS 0.007307f
C565 B.n525 VSUBS 0.007307f
C566 B.n526 VSUBS 0.00505f
C567 B.n527 VSUBS 0.016929f
C568 B.n528 VSUBS 0.00591f
C569 B.n529 VSUBS 0.007307f
C570 B.n530 VSUBS 0.007307f
C571 B.n531 VSUBS 0.007307f
C572 B.n532 VSUBS 0.007307f
C573 B.n533 VSUBS 0.007307f
C574 B.n534 VSUBS 0.007307f
C575 B.n535 VSUBS 0.007307f
C576 B.n536 VSUBS 0.007307f
C577 B.n537 VSUBS 0.007307f
C578 B.n538 VSUBS 0.007307f
C579 B.n539 VSUBS 0.007307f
C580 B.n540 VSUBS 0.00591f
C581 B.n541 VSUBS 0.016929f
C582 B.n542 VSUBS 0.00505f
C583 B.n543 VSUBS 0.007307f
C584 B.n544 VSUBS 0.007307f
C585 B.n545 VSUBS 0.007307f
C586 B.n546 VSUBS 0.007307f
C587 B.n547 VSUBS 0.007307f
C588 B.n548 VSUBS 0.007307f
C589 B.n549 VSUBS 0.007307f
C590 B.n550 VSUBS 0.007307f
C591 B.n551 VSUBS 0.007307f
C592 B.n552 VSUBS 0.007307f
C593 B.n553 VSUBS 0.007307f
C594 B.n554 VSUBS 0.007307f
C595 B.n555 VSUBS 0.007307f
C596 B.n556 VSUBS 0.007307f
C597 B.n557 VSUBS 0.007307f
C598 B.n558 VSUBS 0.007307f
C599 B.n559 VSUBS 0.007307f
C600 B.n560 VSUBS 0.007307f
C601 B.n561 VSUBS 0.007307f
C602 B.n562 VSUBS 0.007307f
C603 B.n563 VSUBS 0.007307f
C604 B.n564 VSUBS 0.007307f
C605 B.n565 VSUBS 0.007307f
C606 B.n566 VSUBS 0.007307f
C607 B.n567 VSUBS 0.007307f
C608 B.n568 VSUBS 0.007307f
C609 B.n569 VSUBS 0.007307f
C610 B.n570 VSUBS 0.007307f
C611 B.n571 VSUBS 0.007307f
C612 B.n572 VSUBS 0.007307f
C613 B.n573 VSUBS 0.007307f
C614 B.n574 VSUBS 0.007307f
C615 B.n575 VSUBS 0.007307f
C616 B.n576 VSUBS 0.007307f
C617 B.n577 VSUBS 0.007307f
C618 B.n578 VSUBS 0.007307f
C619 B.n579 VSUBS 0.007307f
C620 B.n580 VSUBS 0.007307f
C621 B.n581 VSUBS 0.007307f
C622 B.n582 VSUBS 0.007307f
C623 B.n583 VSUBS 0.007307f
C624 B.n584 VSUBS 0.007307f
C625 B.n585 VSUBS 0.007307f
C626 B.n586 VSUBS 0.007307f
C627 B.n587 VSUBS 0.007307f
C628 B.n588 VSUBS 0.007307f
C629 B.n589 VSUBS 0.007307f
C630 B.n590 VSUBS 0.007307f
C631 B.n591 VSUBS 0.007307f
C632 B.n592 VSUBS 0.007307f
C633 B.n593 VSUBS 0.007307f
C634 B.n594 VSUBS 0.007307f
C635 B.n595 VSUBS 0.007307f
C636 B.n596 VSUBS 0.007307f
C637 B.n597 VSUBS 0.007307f
C638 B.n598 VSUBS 0.007307f
C639 B.n599 VSUBS 0.007307f
C640 B.n600 VSUBS 0.007307f
C641 B.n601 VSUBS 0.007307f
C642 B.n602 VSUBS 0.007307f
C643 B.n603 VSUBS 0.007307f
C644 B.n604 VSUBS 0.007307f
C645 B.n605 VSUBS 0.007307f
C646 B.n606 VSUBS 0.007307f
C647 B.n607 VSUBS 0.007307f
C648 B.n608 VSUBS 0.007307f
C649 B.n609 VSUBS 0.007307f
C650 B.n610 VSUBS 0.007307f
C651 B.n611 VSUBS 0.007307f
C652 B.n612 VSUBS 0.007307f
C653 B.n613 VSUBS 0.007307f
C654 B.n614 VSUBS 0.007307f
C655 B.n615 VSUBS 0.007307f
C656 B.n616 VSUBS 0.007307f
C657 B.n617 VSUBS 0.007307f
C658 B.n618 VSUBS 0.007307f
C659 B.n619 VSUBS 0.007307f
C660 B.n620 VSUBS 0.007307f
C661 B.n621 VSUBS 0.007307f
C662 B.n622 VSUBS 0.007307f
C663 B.n623 VSUBS 0.007307f
C664 B.n624 VSUBS 0.007307f
C665 B.n625 VSUBS 0.007307f
C666 B.n626 VSUBS 0.007307f
C667 B.n627 VSUBS 0.007307f
C668 B.n628 VSUBS 0.007307f
C669 B.n629 VSUBS 0.007307f
C670 B.n630 VSUBS 0.007307f
C671 B.n631 VSUBS 0.007307f
C672 B.n632 VSUBS 0.007307f
C673 B.n633 VSUBS 0.007307f
C674 B.n634 VSUBS 0.007307f
C675 B.n635 VSUBS 0.007307f
C676 B.n636 VSUBS 0.007307f
C677 B.n637 VSUBS 0.016744f
C678 B.n638 VSUBS 0.017642f
C679 B.n639 VSUBS 0.016785f
C680 B.n640 VSUBS 0.007307f
C681 B.n641 VSUBS 0.007307f
C682 B.n642 VSUBS 0.007307f
C683 B.n643 VSUBS 0.007307f
C684 B.n644 VSUBS 0.007307f
C685 B.n645 VSUBS 0.007307f
C686 B.n646 VSUBS 0.007307f
C687 B.n647 VSUBS 0.007307f
C688 B.n648 VSUBS 0.007307f
C689 B.n649 VSUBS 0.007307f
C690 B.n650 VSUBS 0.007307f
C691 B.n651 VSUBS 0.007307f
C692 B.n652 VSUBS 0.007307f
C693 B.n653 VSUBS 0.007307f
C694 B.n654 VSUBS 0.007307f
C695 B.n655 VSUBS 0.007307f
C696 B.n656 VSUBS 0.007307f
C697 B.n657 VSUBS 0.007307f
C698 B.n658 VSUBS 0.007307f
C699 B.n659 VSUBS 0.007307f
C700 B.n660 VSUBS 0.007307f
C701 B.n661 VSUBS 0.007307f
C702 B.n662 VSUBS 0.007307f
C703 B.n663 VSUBS 0.007307f
C704 B.n664 VSUBS 0.007307f
C705 B.n665 VSUBS 0.007307f
C706 B.n666 VSUBS 0.007307f
C707 B.n667 VSUBS 0.007307f
C708 B.n668 VSUBS 0.007307f
C709 B.n669 VSUBS 0.007307f
C710 B.n670 VSUBS 0.007307f
C711 B.n671 VSUBS 0.007307f
C712 B.n672 VSUBS 0.007307f
C713 B.n673 VSUBS 0.007307f
C714 B.n674 VSUBS 0.007307f
C715 B.n675 VSUBS 0.007307f
C716 B.n676 VSUBS 0.007307f
C717 B.n677 VSUBS 0.007307f
C718 B.n678 VSUBS 0.007307f
C719 B.n679 VSUBS 0.007307f
C720 B.n680 VSUBS 0.007307f
C721 B.n681 VSUBS 0.007307f
C722 B.n682 VSUBS 0.007307f
C723 B.n683 VSUBS 0.007307f
C724 B.n684 VSUBS 0.007307f
C725 B.n685 VSUBS 0.007307f
C726 B.n686 VSUBS 0.007307f
C727 B.n687 VSUBS 0.007307f
C728 B.n688 VSUBS 0.007307f
C729 B.n689 VSUBS 0.007307f
C730 B.n690 VSUBS 0.007307f
C731 B.n691 VSUBS 0.007307f
C732 B.n692 VSUBS 0.007307f
C733 B.n693 VSUBS 0.007307f
C734 B.n694 VSUBS 0.007307f
C735 B.n695 VSUBS 0.007307f
C736 B.n696 VSUBS 0.007307f
C737 B.n697 VSUBS 0.007307f
C738 B.n698 VSUBS 0.007307f
C739 B.n699 VSUBS 0.007307f
C740 B.n700 VSUBS 0.007307f
C741 B.n701 VSUBS 0.007307f
C742 B.n702 VSUBS 0.007307f
C743 B.n703 VSUBS 0.007307f
C744 B.n704 VSUBS 0.007307f
C745 B.n705 VSUBS 0.007307f
C746 B.n706 VSUBS 0.007307f
C747 B.n707 VSUBS 0.007307f
C748 B.n708 VSUBS 0.007307f
C749 B.n709 VSUBS 0.007307f
C750 B.n710 VSUBS 0.007307f
C751 B.n711 VSUBS 0.007307f
C752 B.n712 VSUBS 0.007307f
C753 B.n713 VSUBS 0.007307f
C754 B.n714 VSUBS 0.007307f
C755 B.n715 VSUBS 0.007307f
C756 B.n716 VSUBS 0.007307f
C757 B.n717 VSUBS 0.007307f
C758 B.n718 VSUBS 0.007307f
C759 B.n719 VSUBS 0.007307f
C760 B.n720 VSUBS 0.007307f
C761 B.n721 VSUBS 0.007307f
C762 B.n722 VSUBS 0.007307f
C763 B.n723 VSUBS 0.007307f
C764 B.n724 VSUBS 0.007307f
C765 B.n725 VSUBS 0.007307f
C766 B.n726 VSUBS 0.007307f
C767 B.n727 VSUBS 0.007307f
C768 B.n728 VSUBS 0.007307f
C769 B.n729 VSUBS 0.007307f
C770 B.n730 VSUBS 0.007307f
C771 B.n731 VSUBS 0.007307f
C772 B.n732 VSUBS 0.007307f
C773 B.n733 VSUBS 0.007307f
C774 B.n734 VSUBS 0.007307f
C775 B.n735 VSUBS 0.007307f
C776 B.n736 VSUBS 0.007307f
C777 B.n737 VSUBS 0.007307f
C778 B.n738 VSUBS 0.007307f
C779 B.n739 VSUBS 0.007307f
C780 B.n740 VSUBS 0.007307f
C781 B.n741 VSUBS 0.007307f
C782 B.n742 VSUBS 0.007307f
C783 B.n743 VSUBS 0.007307f
C784 B.n744 VSUBS 0.007307f
C785 B.n745 VSUBS 0.007307f
C786 B.n746 VSUBS 0.007307f
C787 B.n747 VSUBS 0.007307f
C788 B.n748 VSUBS 0.007307f
C789 B.n749 VSUBS 0.007307f
C790 B.n750 VSUBS 0.007307f
C791 B.n751 VSUBS 0.007307f
C792 B.n752 VSUBS 0.007307f
C793 B.n753 VSUBS 0.007307f
C794 B.n754 VSUBS 0.007307f
C795 B.n755 VSUBS 0.007307f
C796 B.n756 VSUBS 0.007307f
C797 B.n757 VSUBS 0.007307f
C798 B.n758 VSUBS 0.007307f
C799 B.n759 VSUBS 0.007307f
C800 B.n760 VSUBS 0.007307f
C801 B.n761 VSUBS 0.007307f
C802 B.n762 VSUBS 0.007307f
C803 B.n763 VSUBS 0.007307f
C804 B.n764 VSUBS 0.007307f
C805 B.n765 VSUBS 0.007307f
C806 B.n766 VSUBS 0.007307f
C807 B.n767 VSUBS 0.007307f
C808 B.n768 VSUBS 0.007307f
C809 B.n769 VSUBS 0.007307f
C810 B.n770 VSUBS 0.007307f
C811 B.n771 VSUBS 0.007307f
C812 B.n772 VSUBS 0.007307f
C813 B.n773 VSUBS 0.007307f
C814 B.n774 VSUBS 0.007307f
C815 B.n775 VSUBS 0.007307f
C816 B.n776 VSUBS 0.007307f
C817 B.n777 VSUBS 0.007307f
C818 B.n778 VSUBS 0.007307f
C819 B.n779 VSUBS 0.007307f
C820 B.n780 VSUBS 0.007307f
C821 B.n781 VSUBS 0.007307f
C822 B.n782 VSUBS 0.007307f
C823 B.n783 VSUBS 0.007307f
C824 B.n784 VSUBS 0.007307f
C825 B.n785 VSUBS 0.007307f
C826 B.n786 VSUBS 0.007307f
C827 B.n787 VSUBS 0.007307f
C828 B.n788 VSUBS 0.007307f
C829 B.n789 VSUBS 0.007307f
C830 B.n790 VSUBS 0.007307f
C831 B.n791 VSUBS 0.007307f
C832 B.n792 VSUBS 0.007307f
C833 B.n793 VSUBS 0.007307f
C834 B.n794 VSUBS 0.007307f
C835 B.n795 VSUBS 0.007307f
C836 B.n796 VSUBS 0.007307f
C837 B.n797 VSUBS 0.007307f
C838 B.n798 VSUBS 0.007307f
C839 B.n799 VSUBS 0.007307f
C840 B.n800 VSUBS 0.007307f
C841 B.n801 VSUBS 0.007307f
C842 B.n802 VSUBS 0.007307f
C843 B.n803 VSUBS 0.007307f
C844 B.n804 VSUBS 0.007307f
C845 B.n805 VSUBS 0.007307f
C846 B.n806 VSUBS 0.007307f
C847 B.n807 VSUBS 0.007307f
C848 B.n808 VSUBS 0.007307f
C849 B.n809 VSUBS 0.007307f
C850 B.n810 VSUBS 0.007307f
C851 B.n811 VSUBS 0.007307f
C852 B.n812 VSUBS 0.007307f
C853 B.n813 VSUBS 0.007307f
C854 B.n814 VSUBS 0.007307f
C855 B.n815 VSUBS 0.007307f
C856 B.n816 VSUBS 0.007307f
C857 B.n817 VSUBS 0.007307f
C858 B.n818 VSUBS 0.007307f
C859 B.n819 VSUBS 0.007307f
C860 B.n820 VSUBS 0.007307f
C861 B.n821 VSUBS 0.007307f
C862 B.n822 VSUBS 0.007307f
C863 B.n823 VSUBS 0.007307f
C864 B.n824 VSUBS 0.007307f
C865 B.n825 VSUBS 0.007307f
C866 B.n826 VSUBS 0.007307f
C867 B.n827 VSUBS 0.007307f
C868 B.n828 VSUBS 0.007307f
C869 B.n829 VSUBS 0.007307f
C870 B.n830 VSUBS 0.007307f
C871 B.n831 VSUBS 0.007307f
C872 B.n832 VSUBS 0.007307f
C873 B.n833 VSUBS 0.007307f
C874 B.n834 VSUBS 0.007307f
C875 B.n835 VSUBS 0.007307f
C876 B.n836 VSUBS 0.007307f
C877 B.n837 VSUBS 0.007307f
C878 B.n838 VSUBS 0.007307f
C879 B.n839 VSUBS 0.007307f
C880 B.n840 VSUBS 0.007307f
C881 B.n841 VSUBS 0.007307f
C882 B.n842 VSUBS 0.007307f
C883 B.n843 VSUBS 0.007307f
C884 B.n844 VSUBS 0.007307f
C885 B.n845 VSUBS 0.007307f
C886 B.n846 VSUBS 0.007307f
C887 B.n847 VSUBS 0.007307f
C888 B.n848 VSUBS 0.007307f
C889 B.n849 VSUBS 0.007307f
C890 B.n850 VSUBS 0.007307f
C891 B.n851 VSUBS 0.007307f
C892 B.n852 VSUBS 0.007307f
C893 B.n853 VSUBS 0.007307f
C894 B.n854 VSUBS 0.007307f
C895 B.n855 VSUBS 0.007307f
C896 B.n856 VSUBS 0.007307f
C897 B.n857 VSUBS 0.007307f
C898 B.n858 VSUBS 0.007307f
C899 B.n859 VSUBS 0.007307f
C900 B.n860 VSUBS 0.007307f
C901 B.n861 VSUBS 0.007307f
C902 B.n862 VSUBS 0.007307f
C903 B.n863 VSUBS 0.007307f
C904 B.n864 VSUBS 0.007307f
C905 B.n865 VSUBS 0.007307f
C906 B.n866 VSUBS 0.007307f
C907 B.n867 VSUBS 0.007307f
C908 B.n868 VSUBS 0.007307f
C909 B.n869 VSUBS 0.007307f
C910 B.n870 VSUBS 0.007307f
C911 B.n871 VSUBS 0.007307f
C912 B.n872 VSUBS 0.007307f
C913 B.n873 VSUBS 0.007307f
C914 B.n874 VSUBS 0.007307f
C915 B.n875 VSUBS 0.007307f
C916 B.n876 VSUBS 0.007307f
C917 B.n877 VSUBS 0.007307f
C918 B.n878 VSUBS 0.007307f
C919 B.n879 VSUBS 0.007307f
C920 B.n880 VSUBS 0.007307f
C921 B.n881 VSUBS 0.007307f
C922 B.n882 VSUBS 0.007307f
C923 B.n883 VSUBS 0.016785f
C924 B.n884 VSUBS 0.0176f
C925 B.n885 VSUBS 0.0176f
C926 B.n886 VSUBS 0.007307f
C927 B.n887 VSUBS 0.007307f
C928 B.n888 VSUBS 0.007307f
C929 B.n889 VSUBS 0.007307f
C930 B.n890 VSUBS 0.007307f
C931 B.n891 VSUBS 0.007307f
C932 B.n892 VSUBS 0.007307f
C933 B.n893 VSUBS 0.007307f
C934 B.n894 VSUBS 0.007307f
C935 B.n895 VSUBS 0.007307f
C936 B.n896 VSUBS 0.007307f
C937 B.n897 VSUBS 0.007307f
C938 B.n898 VSUBS 0.007307f
C939 B.n899 VSUBS 0.007307f
C940 B.n900 VSUBS 0.007307f
C941 B.n901 VSUBS 0.007307f
C942 B.n902 VSUBS 0.007307f
C943 B.n903 VSUBS 0.007307f
C944 B.n904 VSUBS 0.007307f
C945 B.n905 VSUBS 0.007307f
C946 B.n906 VSUBS 0.007307f
C947 B.n907 VSUBS 0.007307f
C948 B.n908 VSUBS 0.007307f
C949 B.n909 VSUBS 0.007307f
C950 B.n910 VSUBS 0.007307f
C951 B.n911 VSUBS 0.007307f
C952 B.n912 VSUBS 0.007307f
C953 B.n913 VSUBS 0.007307f
C954 B.n914 VSUBS 0.007307f
C955 B.n915 VSUBS 0.007307f
C956 B.n916 VSUBS 0.007307f
C957 B.n917 VSUBS 0.007307f
C958 B.n918 VSUBS 0.007307f
C959 B.n919 VSUBS 0.007307f
C960 B.n920 VSUBS 0.007307f
C961 B.n921 VSUBS 0.007307f
C962 B.n922 VSUBS 0.007307f
C963 B.n923 VSUBS 0.007307f
C964 B.n924 VSUBS 0.007307f
C965 B.n925 VSUBS 0.007307f
C966 B.n926 VSUBS 0.007307f
C967 B.n927 VSUBS 0.007307f
C968 B.n928 VSUBS 0.007307f
C969 B.n929 VSUBS 0.007307f
C970 B.n930 VSUBS 0.007307f
C971 B.n931 VSUBS 0.007307f
C972 B.n932 VSUBS 0.007307f
C973 B.n933 VSUBS 0.007307f
C974 B.n934 VSUBS 0.007307f
C975 B.n935 VSUBS 0.007307f
C976 B.n936 VSUBS 0.007307f
C977 B.n937 VSUBS 0.007307f
C978 B.n938 VSUBS 0.007307f
C979 B.n939 VSUBS 0.007307f
C980 B.n940 VSUBS 0.007307f
C981 B.n941 VSUBS 0.007307f
C982 B.n942 VSUBS 0.007307f
C983 B.n943 VSUBS 0.007307f
C984 B.n944 VSUBS 0.007307f
C985 B.n945 VSUBS 0.007307f
C986 B.n946 VSUBS 0.007307f
C987 B.n947 VSUBS 0.007307f
C988 B.n948 VSUBS 0.007307f
C989 B.n949 VSUBS 0.007307f
C990 B.n950 VSUBS 0.007307f
C991 B.n951 VSUBS 0.007307f
C992 B.n952 VSUBS 0.007307f
C993 B.n953 VSUBS 0.007307f
C994 B.n954 VSUBS 0.007307f
C995 B.n955 VSUBS 0.007307f
C996 B.n956 VSUBS 0.007307f
C997 B.n957 VSUBS 0.007307f
C998 B.n958 VSUBS 0.007307f
C999 B.n959 VSUBS 0.007307f
C1000 B.n960 VSUBS 0.007307f
C1001 B.n961 VSUBS 0.007307f
C1002 B.n962 VSUBS 0.007307f
C1003 B.n963 VSUBS 0.007307f
C1004 B.n964 VSUBS 0.007307f
C1005 B.n965 VSUBS 0.007307f
C1006 B.n966 VSUBS 0.007307f
C1007 B.n967 VSUBS 0.007307f
C1008 B.n968 VSUBS 0.007307f
C1009 B.n969 VSUBS 0.007307f
C1010 B.n970 VSUBS 0.007307f
C1011 B.n971 VSUBS 0.007307f
C1012 B.n972 VSUBS 0.007307f
C1013 B.n973 VSUBS 0.007307f
C1014 B.n974 VSUBS 0.007307f
C1015 B.n975 VSUBS 0.007307f
C1016 B.n976 VSUBS 0.007307f
C1017 B.n977 VSUBS 0.007307f
C1018 B.n978 VSUBS 0.007307f
C1019 B.n979 VSUBS 0.00505f
C1020 B.n980 VSUBS 0.016929f
C1021 B.n981 VSUBS 0.00591f
C1022 B.n982 VSUBS 0.007307f
C1023 B.n983 VSUBS 0.007307f
C1024 B.n984 VSUBS 0.007307f
C1025 B.n985 VSUBS 0.007307f
C1026 B.n986 VSUBS 0.007307f
C1027 B.n987 VSUBS 0.007307f
C1028 B.n988 VSUBS 0.007307f
C1029 B.n989 VSUBS 0.007307f
C1030 B.n990 VSUBS 0.007307f
C1031 B.n991 VSUBS 0.007307f
C1032 B.n992 VSUBS 0.007307f
C1033 B.n993 VSUBS 0.00591f
C1034 B.n994 VSUBS 0.007307f
C1035 B.n995 VSUBS 0.007307f
C1036 B.n996 VSUBS 0.007307f
C1037 B.n997 VSUBS 0.007307f
C1038 B.n998 VSUBS 0.007307f
C1039 B.n999 VSUBS 0.007307f
C1040 B.n1000 VSUBS 0.007307f
C1041 B.n1001 VSUBS 0.007307f
C1042 B.n1002 VSUBS 0.007307f
C1043 B.n1003 VSUBS 0.007307f
C1044 B.n1004 VSUBS 0.007307f
C1045 B.n1005 VSUBS 0.007307f
C1046 B.n1006 VSUBS 0.007307f
C1047 B.n1007 VSUBS 0.007307f
C1048 B.n1008 VSUBS 0.007307f
C1049 B.n1009 VSUBS 0.007307f
C1050 B.n1010 VSUBS 0.007307f
C1051 B.n1011 VSUBS 0.007307f
C1052 B.n1012 VSUBS 0.007307f
C1053 B.n1013 VSUBS 0.007307f
C1054 B.n1014 VSUBS 0.007307f
C1055 B.n1015 VSUBS 0.007307f
C1056 B.n1016 VSUBS 0.007307f
C1057 B.n1017 VSUBS 0.007307f
C1058 B.n1018 VSUBS 0.007307f
C1059 B.n1019 VSUBS 0.007307f
C1060 B.n1020 VSUBS 0.007307f
C1061 B.n1021 VSUBS 0.007307f
C1062 B.n1022 VSUBS 0.007307f
C1063 B.n1023 VSUBS 0.007307f
C1064 B.n1024 VSUBS 0.007307f
C1065 B.n1025 VSUBS 0.007307f
C1066 B.n1026 VSUBS 0.007307f
C1067 B.n1027 VSUBS 0.007307f
C1068 B.n1028 VSUBS 0.007307f
C1069 B.n1029 VSUBS 0.007307f
C1070 B.n1030 VSUBS 0.007307f
C1071 B.n1031 VSUBS 0.007307f
C1072 B.n1032 VSUBS 0.007307f
C1073 B.n1033 VSUBS 0.007307f
C1074 B.n1034 VSUBS 0.007307f
C1075 B.n1035 VSUBS 0.007307f
C1076 B.n1036 VSUBS 0.007307f
C1077 B.n1037 VSUBS 0.007307f
C1078 B.n1038 VSUBS 0.007307f
C1079 B.n1039 VSUBS 0.007307f
C1080 B.n1040 VSUBS 0.007307f
C1081 B.n1041 VSUBS 0.007307f
C1082 B.n1042 VSUBS 0.007307f
C1083 B.n1043 VSUBS 0.007307f
C1084 B.n1044 VSUBS 0.007307f
C1085 B.n1045 VSUBS 0.007307f
C1086 B.n1046 VSUBS 0.007307f
C1087 B.n1047 VSUBS 0.007307f
C1088 B.n1048 VSUBS 0.007307f
C1089 B.n1049 VSUBS 0.007307f
C1090 B.n1050 VSUBS 0.007307f
C1091 B.n1051 VSUBS 0.007307f
C1092 B.n1052 VSUBS 0.007307f
C1093 B.n1053 VSUBS 0.007307f
C1094 B.n1054 VSUBS 0.007307f
C1095 B.n1055 VSUBS 0.007307f
C1096 B.n1056 VSUBS 0.007307f
C1097 B.n1057 VSUBS 0.007307f
C1098 B.n1058 VSUBS 0.007307f
C1099 B.n1059 VSUBS 0.007307f
C1100 B.n1060 VSUBS 0.007307f
C1101 B.n1061 VSUBS 0.007307f
C1102 B.n1062 VSUBS 0.007307f
C1103 B.n1063 VSUBS 0.007307f
C1104 B.n1064 VSUBS 0.007307f
C1105 B.n1065 VSUBS 0.007307f
C1106 B.n1066 VSUBS 0.007307f
C1107 B.n1067 VSUBS 0.007307f
C1108 B.n1068 VSUBS 0.007307f
C1109 B.n1069 VSUBS 0.007307f
C1110 B.n1070 VSUBS 0.007307f
C1111 B.n1071 VSUBS 0.007307f
C1112 B.n1072 VSUBS 0.007307f
C1113 B.n1073 VSUBS 0.007307f
C1114 B.n1074 VSUBS 0.007307f
C1115 B.n1075 VSUBS 0.007307f
C1116 B.n1076 VSUBS 0.007307f
C1117 B.n1077 VSUBS 0.007307f
C1118 B.n1078 VSUBS 0.007307f
C1119 B.n1079 VSUBS 0.007307f
C1120 B.n1080 VSUBS 0.007307f
C1121 B.n1081 VSUBS 0.007307f
C1122 B.n1082 VSUBS 0.007307f
C1123 B.n1083 VSUBS 0.007307f
C1124 B.n1084 VSUBS 0.007307f
C1125 B.n1085 VSUBS 0.007307f
C1126 B.n1086 VSUBS 0.007307f
C1127 B.n1087 VSUBS 0.007307f
C1128 B.n1088 VSUBS 0.007307f
C1129 B.n1089 VSUBS 0.0176f
C1130 B.n1090 VSUBS 0.0176f
C1131 B.n1091 VSUBS 0.016785f
C1132 B.n1092 VSUBS 0.007307f
C1133 B.n1093 VSUBS 0.007307f
C1134 B.n1094 VSUBS 0.007307f
C1135 B.n1095 VSUBS 0.007307f
C1136 B.n1096 VSUBS 0.007307f
C1137 B.n1097 VSUBS 0.007307f
C1138 B.n1098 VSUBS 0.007307f
C1139 B.n1099 VSUBS 0.007307f
C1140 B.n1100 VSUBS 0.007307f
C1141 B.n1101 VSUBS 0.007307f
C1142 B.n1102 VSUBS 0.007307f
C1143 B.n1103 VSUBS 0.007307f
C1144 B.n1104 VSUBS 0.007307f
C1145 B.n1105 VSUBS 0.007307f
C1146 B.n1106 VSUBS 0.007307f
C1147 B.n1107 VSUBS 0.007307f
C1148 B.n1108 VSUBS 0.007307f
C1149 B.n1109 VSUBS 0.007307f
C1150 B.n1110 VSUBS 0.007307f
C1151 B.n1111 VSUBS 0.007307f
C1152 B.n1112 VSUBS 0.007307f
C1153 B.n1113 VSUBS 0.007307f
C1154 B.n1114 VSUBS 0.007307f
C1155 B.n1115 VSUBS 0.007307f
C1156 B.n1116 VSUBS 0.007307f
C1157 B.n1117 VSUBS 0.007307f
C1158 B.n1118 VSUBS 0.007307f
C1159 B.n1119 VSUBS 0.007307f
C1160 B.n1120 VSUBS 0.007307f
C1161 B.n1121 VSUBS 0.007307f
C1162 B.n1122 VSUBS 0.007307f
C1163 B.n1123 VSUBS 0.007307f
C1164 B.n1124 VSUBS 0.007307f
C1165 B.n1125 VSUBS 0.007307f
C1166 B.n1126 VSUBS 0.007307f
C1167 B.n1127 VSUBS 0.007307f
C1168 B.n1128 VSUBS 0.007307f
C1169 B.n1129 VSUBS 0.007307f
C1170 B.n1130 VSUBS 0.007307f
C1171 B.n1131 VSUBS 0.007307f
C1172 B.n1132 VSUBS 0.007307f
C1173 B.n1133 VSUBS 0.007307f
C1174 B.n1134 VSUBS 0.007307f
C1175 B.n1135 VSUBS 0.007307f
C1176 B.n1136 VSUBS 0.007307f
C1177 B.n1137 VSUBS 0.007307f
C1178 B.n1138 VSUBS 0.007307f
C1179 B.n1139 VSUBS 0.007307f
C1180 B.n1140 VSUBS 0.007307f
C1181 B.n1141 VSUBS 0.007307f
C1182 B.n1142 VSUBS 0.007307f
C1183 B.n1143 VSUBS 0.007307f
C1184 B.n1144 VSUBS 0.007307f
C1185 B.n1145 VSUBS 0.007307f
C1186 B.n1146 VSUBS 0.007307f
C1187 B.n1147 VSUBS 0.007307f
C1188 B.n1148 VSUBS 0.007307f
C1189 B.n1149 VSUBS 0.007307f
C1190 B.n1150 VSUBS 0.007307f
C1191 B.n1151 VSUBS 0.007307f
C1192 B.n1152 VSUBS 0.007307f
C1193 B.n1153 VSUBS 0.007307f
C1194 B.n1154 VSUBS 0.007307f
C1195 B.n1155 VSUBS 0.007307f
C1196 B.n1156 VSUBS 0.007307f
C1197 B.n1157 VSUBS 0.007307f
C1198 B.n1158 VSUBS 0.007307f
C1199 B.n1159 VSUBS 0.007307f
C1200 B.n1160 VSUBS 0.007307f
C1201 B.n1161 VSUBS 0.007307f
C1202 B.n1162 VSUBS 0.007307f
C1203 B.n1163 VSUBS 0.007307f
C1204 B.n1164 VSUBS 0.007307f
C1205 B.n1165 VSUBS 0.007307f
C1206 B.n1166 VSUBS 0.007307f
C1207 B.n1167 VSUBS 0.007307f
C1208 B.n1168 VSUBS 0.007307f
C1209 B.n1169 VSUBS 0.007307f
C1210 B.n1170 VSUBS 0.007307f
C1211 B.n1171 VSUBS 0.007307f
C1212 B.n1172 VSUBS 0.007307f
C1213 B.n1173 VSUBS 0.007307f
C1214 B.n1174 VSUBS 0.007307f
C1215 B.n1175 VSUBS 0.007307f
C1216 B.n1176 VSUBS 0.007307f
C1217 B.n1177 VSUBS 0.007307f
C1218 B.n1178 VSUBS 0.007307f
C1219 B.n1179 VSUBS 0.007307f
C1220 B.n1180 VSUBS 0.007307f
C1221 B.n1181 VSUBS 0.007307f
C1222 B.n1182 VSUBS 0.007307f
C1223 B.n1183 VSUBS 0.007307f
C1224 B.n1184 VSUBS 0.007307f
C1225 B.n1185 VSUBS 0.007307f
C1226 B.n1186 VSUBS 0.007307f
C1227 B.n1187 VSUBS 0.007307f
C1228 B.n1188 VSUBS 0.007307f
C1229 B.n1189 VSUBS 0.007307f
C1230 B.n1190 VSUBS 0.007307f
C1231 B.n1191 VSUBS 0.007307f
C1232 B.n1192 VSUBS 0.007307f
C1233 B.n1193 VSUBS 0.007307f
C1234 B.n1194 VSUBS 0.007307f
C1235 B.n1195 VSUBS 0.007307f
C1236 B.n1196 VSUBS 0.007307f
C1237 B.n1197 VSUBS 0.007307f
C1238 B.n1198 VSUBS 0.007307f
C1239 B.n1199 VSUBS 0.007307f
C1240 B.n1200 VSUBS 0.007307f
C1241 B.n1201 VSUBS 0.007307f
C1242 B.n1202 VSUBS 0.007307f
C1243 B.n1203 VSUBS 0.007307f
C1244 B.n1204 VSUBS 0.007307f
C1245 B.n1205 VSUBS 0.007307f
C1246 B.n1206 VSUBS 0.007307f
C1247 B.n1207 VSUBS 0.007307f
C1248 B.n1208 VSUBS 0.007307f
C1249 B.n1209 VSUBS 0.007307f
C1250 B.n1210 VSUBS 0.007307f
C1251 B.n1211 VSUBS 0.009535f
C1252 B.n1212 VSUBS 0.010157f
C1253 B.n1213 VSUBS 0.020199f
C1254 VDD2.n0 VSUBS 0.031819f
C1255 VDD2.n1 VSUBS 0.028867f
C1256 VDD2.n2 VSUBS 0.015512f
C1257 VDD2.n3 VSUBS 0.036665f
C1258 VDD2.n4 VSUBS 0.016424f
C1259 VDD2.n5 VSUBS 0.028867f
C1260 VDD2.n6 VSUBS 0.015512f
C1261 VDD2.n7 VSUBS 0.036665f
C1262 VDD2.n8 VSUBS 0.016424f
C1263 VDD2.n9 VSUBS 0.028867f
C1264 VDD2.n10 VSUBS 0.015512f
C1265 VDD2.n11 VSUBS 0.036665f
C1266 VDD2.n12 VSUBS 0.016424f
C1267 VDD2.n13 VSUBS 0.028867f
C1268 VDD2.n14 VSUBS 0.015512f
C1269 VDD2.n15 VSUBS 0.036665f
C1270 VDD2.n16 VSUBS 0.016424f
C1271 VDD2.n17 VSUBS 0.028867f
C1272 VDD2.n18 VSUBS 0.015512f
C1273 VDD2.n19 VSUBS 0.036665f
C1274 VDD2.n20 VSUBS 0.016424f
C1275 VDD2.n21 VSUBS 0.028867f
C1276 VDD2.n22 VSUBS 0.015512f
C1277 VDD2.n23 VSUBS 0.036665f
C1278 VDD2.n24 VSUBS 0.016424f
C1279 VDD2.n25 VSUBS 0.028867f
C1280 VDD2.n26 VSUBS 0.015512f
C1281 VDD2.n27 VSUBS 0.036665f
C1282 VDD2.n28 VSUBS 0.016424f
C1283 VDD2.n29 VSUBS 0.028867f
C1284 VDD2.n30 VSUBS 0.015512f
C1285 VDD2.n31 VSUBS 0.036665f
C1286 VDD2.n32 VSUBS 0.016424f
C1287 VDD2.n33 VSUBS 0.325503f
C1288 VDD2.t5 VSUBS 0.079742f
C1289 VDD2.n34 VSUBS 0.027499f
C1290 VDD2.n35 VSUBS 0.027581f
C1291 VDD2.n36 VSUBS 0.015512f
C1292 VDD2.n37 VSUBS 2.36952f
C1293 VDD2.n38 VSUBS 0.028867f
C1294 VDD2.n39 VSUBS 0.015512f
C1295 VDD2.n40 VSUBS 0.016424f
C1296 VDD2.n41 VSUBS 0.036665f
C1297 VDD2.n42 VSUBS 0.036665f
C1298 VDD2.n43 VSUBS 0.016424f
C1299 VDD2.n44 VSUBS 0.015512f
C1300 VDD2.n45 VSUBS 0.028867f
C1301 VDD2.n46 VSUBS 0.028867f
C1302 VDD2.n47 VSUBS 0.015512f
C1303 VDD2.n48 VSUBS 0.016424f
C1304 VDD2.n49 VSUBS 0.036665f
C1305 VDD2.n50 VSUBS 0.036665f
C1306 VDD2.n51 VSUBS 0.036665f
C1307 VDD2.n52 VSUBS 0.016424f
C1308 VDD2.n53 VSUBS 0.015512f
C1309 VDD2.n54 VSUBS 0.028867f
C1310 VDD2.n55 VSUBS 0.028867f
C1311 VDD2.n56 VSUBS 0.015512f
C1312 VDD2.n57 VSUBS 0.015968f
C1313 VDD2.n58 VSUBS 0.015968f
C1314 VDD2.n59 VSUBS 0.036665f
C1315 VDD2.n60 VSUBS 0.036665f
C1316 VDD2.n61 VSUBS 0.016424f
C1317 VDD2.n62 VSUBS 0.015512f
C1318 VDD2.n63 VSUBS 0.028867f
C1319 VDD2.n64 VSUBS 0.028867f
C1320 VDD2.n65 VSUBS 0.015512f
C1321 VDD2.n66 VSUBS 0.016424f
C1322 VDD2.n67 VSUBS 0.036665f
C1323 VDD2.n68 VSUBS 0.036665f
C1324 VDD2.n69 VSUBS 0.016424f
C1325 VDD2.n70 VSUBS 0.015512f
C1326 VDD2.n71 VSUBS 0.028867f
C1327 VDD2.n72 VSUBS 0.028867f
C1328 VDD2.n73 VSUBS 0.015512f
C1329 VDD2.n74 VSUBS 0.016424f
C1330 VDD2.n75 VSUBS 0.036665f
C1331 VDD2.n76 VSUBS 0.036665f
C1332 VDD2.n77 VSUBS 0.016424f
C1333 VDD2.n78 VSUBS 0.015512f
C1334 VDD2.n79 VSUBS 0.028867f
C1335 VDD2.n80 VSUBS 0.028867f
C1336 VDD2.n81 VSUBS 0.015512f
C1337 VDD2.n82 VSUBS 0.016424f
C1338 VDD2.n83 VSUBS 0.036665f
C1339 VDD2.n84 VSUBS 0.036665f
C1340 VDD2.n85 VSUBS 0.016424f
C1341 VDD2.n86 VSUBS 0.015512f
C1342 VDD2.n87 VSUBS 0.028867f
C1343 VDD2.n88 VSUBS 0.028867f
C1344 VDD2.n89 VSUBS 0.015512f
C1345 VDD2.n90 VSUBS 0.016424f
C1346 VDD2.n91 VSUBS 0.036665f
C1347 VDD2.n92 VSUBS 0.036665f
C1348 VDD2.n93 VSUBS 0.016424f
C1349 VDD2.n94 VSUBS 0.015512f
C1350 VDD2.n95 VSUBS 0.028867f
C1351 VDD2.n96 VSUBS 0.028867f
C1352 VDD2.n97 VSUBS 0.015512f
C1353 VDD2.n98 VSUBS 0.016424f
C1354 VDD2.n99 VSUBS 0.036665f
C1355 VDD2.n100 VSUBS 0.092389f
C1356 VDD2.n101 VSUBS 0.016424f
C1357 VDD2.n102 VSUBS 0.030462f
C1358 VDD2.n103 VSUBS 0.074613f
C1359 VDD2.n104 VSUBS 0.116414f
C1360 VDD2.t6 VSUBS 0.445287f
C1361 VDD2.t1 VSUBS 0.445287f
C1362 VDD2.n105 VSUBS 3.76292f
C1363 VDD2.n106 VSUBS 1.32875f
C1364 VDD2.t0 VSUBS 0.445287f
C1365 VDD2.t2 VSUBS 0.445287f
C1366 VDD2.n107 VSUBS 3.80323f
C1367 VDD2.n108 VSUBS 4.94504f
C1368 VDD2.n109 VSUBS 0.031819f
C1369 VDD2.n110 VSUBS 0.028867f
C1370 VDD2.n111 VSUBS 0.015512f
C1371 VDD2.n112 VSUBS 0.036665f
C1372 VDD2.n113 VSUBS 0.016424f
C1373 VDD2.n114 VSUBS 0.028867f
C1374 VDD2.n115 VSUBS 0.015512f
C1375 VDD2.n116 VSUBS 0.036665f
C1376 VDD2.n117 VSUBS 0.016424f
C1377 VDD2.n118 VSUBS 0.028867f
C1378 VDD2.n119 VSUBS 0.015512f
C1379 VDD2.n120 VSUBS 0.036665f
C1380 VDD2.n121 VSUBS 0.016424f
C1381 VDD2.n122 VSUBS 0.028867f
C1382 VDD2.n123 VSUBS 0.015512f
C1383 VDD2.n124 VSUBS 0.036665f
C1384 VDD2.n125 VSUBS 0.016424f
C1385 VDD2.n126 VSUBS 0.028867f
C1386 VDD2.n127 VSUBS 0.015512f
C1387 VDD2.n128 VSUBS 0.036665f
C1388 VDD2.n129 VSUBS 0.016424f
C1389 VDD2.n130 VSUBS 0.028867f
C1390 VDD2.n131 VSUBS 0.015512f
C1391 VDD2.n132 VSUBS 0.036665f
C1392 VDD2.n133 VSUBS 0.016424f
C1393 VDD2.n134 VSUBS 0.028867f
C1394 VDD2.n135 VSUBS 0.015512f
C1395 VDD2.n136 VSUBS 0.036665f
C1396 VDD2.n137 VSUBS 0.036665f
C1397 VDD2.n138 VSUBS 0.016424f
C1398 VDD2.n139 VSUBS 0.028867f
C1399 VDD2.n140 VSUBS 0.015512f
C1400 VDD2.n141 VSUBS 0.036665f
C1401 VDD2.n142 VSUBS 0.016424f
C1402 VDD2.n143 VSUBS 0.325502f
C1403 VDD2.t9 VSUBS 0.079742f
C1404 VDD2.n144 VSUBS 0.027499f
C1405 VDD2.n145 VSUBS 0.027581f
C1406 VDD2.n146 VSUBS 0.015512f
C1407 VDD2.n147 VSUBS 2.36952f
C1408 VDD2.n148 VSUBS 0.028867f
C1409 VDD2.n149 VSUBS 0.015512f
C1410 VDD2.n150 VSUBS 0.016424f
C1411 VDD2.n151 VSUBS 0.036665f
C1412 VDD2.n152 VSUBS 0.036665f
C1413 VDD2.n153 VSUBS 0.016424f
C1414 VDD2.n154 VSUBS 0.015512f
C1415 VDD2.n155 VSUBS 0.028867f
C1416 VDD2.n156 VSUBS 0.028867f
C1417 VDD2.n157 VSUBS 0.015512f
C1418 VDD2.n158 VSUBS 0.016424f
C1419 VDD2.n159 VSUBS 0.036665f
C1420 VDD2.n160 VSUBS 0.036665f
C1421 VDD2.n161 VSUBS 0.016424f
C1422 VDD2.n162 VSUBS 0.015512f
C1423 VDD2.n163 VSUBS 0.028867f
C1424 VDD2.n164 VSUBS 0.028867f
C1425 VDD2.n165 VSUBS 0.015512f
C1426 VDD2.n166 VSUBS 0.015968f
C1427 VDD2.n167 VSUBS 0.015968f
C1428 VDD2.n168 VSUBS 0.036665f
C1429 VDD2.n169 VSUBS 0.036665f
C1430 VDD2.n170 VSUBS 0.016424f
C1431 VDD2.n171 VSUBS 0.015512f
C1432 VDD2.n172 VSUBS 0.028867f
C1433 VDD2.n173 VSUBS 0.028867f
C1434 VDD2.n174 VSUBS 0.015512f
C1435 VDD2.n175 VSUBS 0.016424f
C1436 VDD2.n176 VSUBS 0.036665f
C1437 VDD2.n177 VSUBS 0.036665f
C1438 VDD2.n178 VSUBS 0.016424f
C1439 VDD2.n179 VSUBS 0.015512f
C1440 VDD2.n180 VSUBS 0.028867f
C1441 VDD2.n181 VSUBS 0.028867f
C1442 VDD2.n182 VSUBS 0.015512f
C1443 VDD2.n183 VSUBS 0.016424f
C1444 VDD2.n184 VSUBS 0.036665f
C1445 VDD2.n185 VSUBS 0.036665f
C1446 VDD2.n186 VSUBS 0.016424f
C1447 VDD2.n187 VSUBS 0.015512f
C1448 VDD2.n188 VSUBS 0.028867f
C1449 VDD2.n189 VSUBS 0.028867f
C1450 VDD2.n190 VSUBS 0.015512f
C1451 VDD2.n191 VSUBS 0.016424f
C1452 VDD2.n192 VSUBS 0.036665f
C1453 VDD2.n193 VSUBS 0.036665f
C1454 VDD2.n194 VSUBS 0.016424f
C1455 VDD2.n195 VSUBS 0.015512f
C1456 VDD2.n196 VSUBS 0.028867f
C1457 VDD2.n197 VSUBS 0.028867f
C1458 VDD2.n198 VSUBS 0.015512f
C1459 VDD2.n199 VSUBS 0.016424f
C1460 VDD2.n200 VSUBS 0.036665f
C1461 VDD2.n201 VSUBS 0.036665f
C1462 VDD2.n202 VSUBS 0.016424f
C1463 VDD2.n203 VSUBS 0.015512f
C1464 VDD2.n204 VSUBS 0.028867f
C1465 VDD2.n205 VSUBS 0.028867f
C1466 VDD2.n206 VSUBS 0.015512f
C1467 VDD2.n207 VSUBS 0.016424f
C1468 VDD2.n208 VSUBS 0.036665f
C1469 VDD2.n209 VSUBS 0.092389f
C1470 VDD2.n210 VSUBS 0.016424f
C1471 VDD2.n211 VSUBS 0.030462f
C1472 VDD2.n212 VSUBS 0.074613f
C1473 VDD2.n213 VSUBS 0.09135f
C1474 VDD2.n214 VSUBS 4.55316f
C1475 VDD2.t8 VSUBS 0.445287f
C1476 VDD2.t7 VSUBS 0.445287f
C1477 VDD2.n215 VSUBS 3.76293f
C1478 VDD2.n216 VSUBS 0.969882f
C1479 VDD2.t3 VSUBS 0.445287f
C1480 VDD2.t4 VSUBS 0.445287f
C1481 VDD2.n217 VSUBS 3.80317f
C1482 VN.t7 VSUBS 4.06388f
C1483 VN.n0 VSUBS 1.4709f
C1484 VN.n1 VSUBS 0.019733f
C1485 VN.n2 VSUBS 0.039196f
C1486 VN.n3 VSUBS 0.019733f
C1487 VN.n4 VSUBS 0.036594f
C1488 VN.n5 VSUBS 0.019733f
C1489 VN.t9 VSUBS 4.06388f
C1490 VN.n6 VSUBS 0.036594f
C1491 VN.n7 VSUBS 0.019733f
C1492 VN.n8 VSUBS 0.036594f
C1493 VN.n9 VSUBS 0.019733f
C1494 VN.t8 VSUBS 4.06388f
C1495 VN.n10 VSUBS 0.036594f
C1496 VN.n11 VSUBS 0.019733f
C1497 VN.n12 VSUBS 0.036594f
C1498 VN.t4 VSUBS 4.39354f
C1499 VN.n13 VSUBS 1.40549f
C1500 VN.t3 VSUBS 4.06388f
C1501 VN.n14 VSUBS 1.47305f
C1502 VN.n15 VSUBS 0.033342f
C1503 VN.n16 VSUBS 0.253914f
C1504 VN.n17 VSUBS 0.019733f
C1505 VN.n18 VSUBS 0.019733f
C1506 VN.n19 VSUBS 0.036594f
C1507 VN.n20 VSUBS 0.024318f
C1508 VN.n21 VSUBS 0.033053f
C1509 VN.n22 VSUBS 0.019733f
C1510 VN.n23 VSUBS 0.019733f
C1511 VN.n24 VSUBS 0.019733f
C1512 VN.n25 VSUBS 0.036594f
C1513 VN.n26 VSUBS 0.027561f
C1514 VN.n27 VSUBS 1.39623f
C1515 VN.n28 VSUBS 0.027561f
C1516 VN.n29 VSUBS 0.019733f
C1517 VN.n30 VSUBS 0.019733f
C1518 VN.n31 VSUBS 0.019733f
C1519 VN.n32 VSUBS 0.036594f
C1520 VN.n33 VSUBS 0.033053f
C1521 VN.n34 VSUBS 0.024318f
C1522 VN.n35 VSUBS 0.019733f
C1523 VN.n36 VSUBS 0.019733f
C1524 VN.n37 VSUBS 0.019733f
C1525 VN.n38 VSUBS 0.036594f
C1526 VN.n39 VSUBS 0.033342f
C1527 VN.n40 VSUBS 1.39623f
C1528 VN.n41 VSUBS 0.02178f
C1529 VN.n42 VSUBS 0.019733f
C1530 VN.n43 VSUBS 0.019733f
C1531 VN.n44 VSUBS 0.019733f
C1532 VN.n45 VSUBS 0.036594f
C1533 VN.n46 VSUBS 0.038805f
C1534 VN.n47 VSUBS 0.015963f
C1535 VN.n48 VSUBS 0.019733f
C1536 VN.n49 VSUBS 0.019733f
C1537 VN.n50 VSUBS 0.019733f
C1538 VN.n51 VSUBS 0.036594f
C1539 VN.n52 VSUBS 0.036594f
C1540 VN.n53 VSUBS 0.021057f
C1541 VN.n54 VSUBS 0.031844f
C1542 VN.n55 VSUBS 0.060543f
C1543 VN.t0 VSUBS 4.06388f
C1544 VN.n56 VSUBS 1.4709f
C1545 VN.n57 VSUBS 0.019733f
C1546 VN.n58 VSUBS 0.039196f
C1547 VN.n59 VSUBS 0.019733f
C1548 VN.n60 VSUBS 0.036594f
C1549 VN.n61 VSUBS 0.019733f
C1550 VN.t1 VSUBS 4.06388f
C1551 VN.n62 VSUBS 0.036594f
C1552 VN.n63 VSUBS 0.019733f
C1553 VN.n64 VSUBS 0.036594f
C1554 VN.n65 VSUBS 0.019733f
C1555 VN.t2 VSUBS 4.06388f
C1556 VN.n66 VSUBS 0.036594f
C1557 VN.n67 VSUBS 0.019733f
C1558 VN.n68 VSUBS 0.036594f
C1559 VN.t5 VSUBS 4.39354f
C1560 VN.n69 VSUBS 1.40549f
C1561 VN.t6 VSUBS 4.06388f
C1562 VN.n70 VSUBS 1.47305f
C1563 VN.n71 VSUBS 0.033342f
C1564 VN.n72 VSUBS 0.253914f
C1565 VN.n73 VSUBS 0.019733f
C1566 VN.n74 VSUBS 0.019733f
C1567 VN.n75 VSUBS 0.036594f
C1568 VN.n76 VSUBS 0.024318f
C1569 VN.n77 VSUBS 0.033053f
C1570 VN.n78 VSUBS 0.019733f
C1571 VN.n79 VSUBS 0.019733f
C1572 VN.n80 VSUBS 0.019733f
C1573 VN.n81 VSUBS 0.036594f
C1574 VN.n82 VSUBS 0.027561f
C1575 VN.n83 VSUBS 1.39623f
C1576 VN.n84 VSUBS 0.027561f
C1577 VN.n85 VSUBS 0.019733f
C1578 VN.n86 VSUBS 0.019733f
C1579 VN.n87 VSUBS 0.019733f
C1580 VN.n88 VSUBS 0.036594f
C1581 VN.n89 VSUBS 0.033053f
C1582 VN.n90 VSUBS 0.024318f
C1583 VN.n91 VSUBS 0.019733f
C1584 VN.n92 VSUBS 0.019733f
C1585 VN.n93 VSUBS 0.019733f
C1586 VN.n94 VSUBS 0.036594f
C1587 VN.n95 VSUBS 0.033342f
C1588 VN.n96 VSUBS 1.39623f
C1589 VN.n97 VSUBS 0.02178f
C1590 VN.n98 VSUBS 0.019733f
C1591 VN.n99 VSUBS 0.019733f
C1592 VN.n100 VSUBS 0.019733f
C1593 VN.n101 VSUBS 0.036594f
C1594 VN.n102 VSUBS 0.038805f
C1595 VN.n103 VSUBS 0.015963f
C1596 VN.n104 VSUBS 0.019733f
C1597 VN.n105 VSUBS 0.019733f
C1598 VN.n106 VSUBS 0.019733f
C1599 VN.n107 VSUBS 0.036594f
C1600 VN.n108 VSUBS 0.036594f
C1601 VN.n109 VSUBS 0.021057f
C1602 VN.n110 VSUBS 0.031844f
C1603 VN.n111 VSUBS 1.64503f
C1604 VDD1.n0 VSUBS 0.031888f
C1605 VDD1.n1 VSUBS 0.02893f
C1606 VDD1.n2 VSUBS 0.015546f
C1607 VDD1.n3 VSUBS 0.036744f
C1608 VDD1.n4 VSUBS 0.01646f
C1609 VDD1.n5 VSUBS 0.02893f
C1610 VDD1.n6 VSUBS 0.015546f
C1611 VDD1.n7 VSUBS 0.036744f
C1612 VDD1.n8 VSUBS 0.01646f
C1613 VDD1.n9 VSUBS 0.02893f
C1614 VDD1.n10 VSUBS 0.015546f
C1615 VDD1.n11 VSUBS 0.036744f
C1616 VDD1.n12 VSUBS 0.01646f
C1617 VDD1.n13 VSUBS 0.02893f
C1618 VDD1.n14 VSUBS 0.015546f
C1619 VDD1.n15 VSUBS 0.036744f
C1620 VDD1.n16 VSUBS 0.01646f
C1621 VDD1.n17 VSUBS 0.02893f
C1622 VDD1.n18 VSUBS 0.015546f
C1623 VDD1.n19 VSUBS 0.036744f
C1624 VDD1.n20 VSUBS 0.01646f
C1625 VDD1.n21 VSUBS 0.02893f
C1626 VDD1.n22 VSUBS 0.015546f
C1627 VDD1.n23 VSUBS 0.036744f
C1628 VDD1.n24 VSUBS 0.01646f
C1629 VDD1.n25 VSUBS 0.02893f
C1630 VDD1.n26 VSUBS 0.015546f
C1631 VDD1.n27 VSUBS 0.036744f
C1632 VDD1.n28 VSUBS 0.036744f
C1633 VDD1.n29 VSUBS 0.01646f
C1634 VDD1.n30 VSUBS 0.02893f
C1635 VDD1.n31 VSUBS 0.015546f
C1636 VDD1.n32 VSUBS 0.036744f
C1637 VDD1.n33 VSUBS 0.01646f
C1638 VDD1.n34 VSUBS 0.326209f
C1639 VDD1.t9 VSUBS 0.079915f
C1640 VDD1.n35 VSUBS 0.027558f
C1641 VDD1.n36 VSUBS 0.027641f
C1642 VDD1.n37 VSUBS 0.015546f
C1643 VDD1.n38 VSUBS 2.37466f
C1644 VDD1.n39 VSUBS 0.02893f
C1645 VDD1.n40 VSUBS 0.015546f
C1646 VDD1.n41 VSUBS 0.01646f
C1647 VDD1.n42 VSUBS 0.036744f
C1648 VDD1.n43 VSUBS 0.036744f
C1649 VDD1.n44 VSUBS 0.01646f
C1650 VDD1.n45 VSUBS 0.015546f
C1651 VDD1.n46 VSUBS 0.02893f
C1652 VDD1.n47 VSUBS 0.02893f
C1653 VDD1.n48 VSUBS 0.015546f
C1654 VDD1.n49 VSUBS 0.01646f
C1655 VDD1.n50 VSUBS 0.036744f
C1656 VDD1.n51 VSUBS 0.036744f
C1657 VDD1.n52 VSUBS 0.01646f
C1658 VDD1.n53 VSUBS 0.015546f
C1659 VDD1.n54 VSUBS 0.02893f
C1660 VDD1.n55 VSUBS 0.02893f
C1661 VDD1.n56 VSUBS 0.015546f
C1662 VDD1.n57 VSUBS 0.016003f
C1663 VDD1.n58 VSUBS 0.016003f
C1664 VDD1.n59 VSUBS 0.036744f
C1665 VDD1.n60 VSUBS 0.036744f
C1666 VDD1.n61 VSUBS 0.01646f
C1667 VDD1.n62 VSUBS 0.015546f
C1668 VDD1.n63 VSUBS 0.02893f
C1669 VDD1.n64 VSUBS 0.02893f
C1670 VDD1.n65 VSUBS 0.015546f
C1671 VDD1.n66 VSUBS 0.01646f
C1672 VDD1.n67 VSUBS 0.036744f
C1673 VDD1.n68 VSUBS 0.036744f
C1674 VDD1.n69 VSUBS 0.01646f
C1675 VDD1.n70 VSUBS 0.015546f
C1676 VDD1.n71 VSUBS 0.02893f
C1677 VDD1.n72 VSUBS 0.02893f
C1678 VDD1.n73 VSUBS 0.015546f
C1679 VDD1.n74 VSUBS 0.01646f
C1680 VDD1.n75 VSUBS 0.036744f
C1681 VDD1.n76 VSUBS 0.036744f
C1682 VDD1.n77 VSUBS 0.01646f
C1683 VDD1.n78 VSUBS 0.015546f
C1684 VDD1.n79 VSUBS 0.02893f
C1685 VDD1.n80 VSUBS 0.02893f
C1686 VDD1.n81 VSUBS 0.015546f
C1687 VDD1.n82 VSUBS 0.01646f
C1688 VDD1.n83 VSUBS 0.036744f
C1689 VDD1.n84 VSUBS 0.036744f
C1690 VDD1.n85 VSUBS 0.01646f
C1691 VDD1.n86 VSUBS 0.015546f
C1692 VDD1.n87 VSUBS 0.02893f
C1693 VDD1.n88 VSUBS 0.02893f
C1694 VDD1.n89 VSUBS 0.015546f
C1695 VDD1.n90 VSUBS 0.01646f
C1696 VDD1.n91 VSUBS 0.036744f
C1697 VDD1.n92 VSUBS 0.036744f
C1698 VDD1.n93 VSUBS 0.01646f
C1699 VDD1.n94 VSUBS 0.015546f
C1700 VDD1.n95 VSUBS 0.02893f
C1701 VDD1.n96 VSUBS 0.02893f
C1702 VDD1.n97 VSUBS 0.015546f
C1703 VDD1.n98 VSUBS 0.01646f
C1704 VDD1.n99 VSUBS 0.036744f
C1705 VDD1.n100 VSUBS 0.09259f
C1706 VDD1.n101 VSUBS 0.01646f
C1707 VDD1.n102 VSUBS 0.030528f
C1708 VDD1.n103 VSUBS 0.074775f
C1709 VDD1.n104 VSUBS 0.116667f
C1710 VDD1.t6 VSUBS 0.446254f
C1711 VDD1.t7 VSUBS 0.446254f
C1712 VDD1.n105 VSUBS 3.7711f
C1713 VDD1.n106 VSUBS 1.34141f
C1714 VDD1.n107 VSUBS 0.031888f
C1715 VDD1.n108 VSUBS 0.02893f
C1716 VDD1.n109 VSUBS 0.015546f
C1717 VDD1.n110 VSUBS 0.036744f
C1718 VDD1.n111 VSUBS 0.01646f
C1719 VDD1.n112 VSUBS 0.02893f
C1720 VDD1.n113 VSUBS 0.015546f
C1721 VDD1.n114 VSUBS 0.036744f
C1722 VDD1.n115 VSUBS 0.01646f
C1723 VDD1.n116 VSUBS 0.02893f
C1724 VDD1.n117 VSUBS 0.015546f
C1725 VDD1.n118 VSUBS 0.036744f
C1726 VDD1.n119 VSUBS 0.01646f
C1727 VDD1.n120 VSUBS 0.02893f
C1728 VDD1.n121 VSUBS 0.015546f
C1729 VDD1.n122 VSUBS 0.036744f
C1730 VDD1.n123 VSUBS 0.01646f
C1731 VDD1.n124 VSUBS 0.02893f
C1732 VDD1.n125 VSUBS 0.015546f
C1733 VDD1.n126 VSUBS 0.036744f
C1734 VDD1.n127 VSUBS 0.01646f
C1735 VDD1.n128 VSUBS 0.02893f
C1736 VDD1.n129 VSUBS 0.015546f
C1737 VDD1.n130 VSUBS 0.036744f
C1738 VDD1.n131 VSUBS 0.01646f
C1739 VDD1.n132 VSUBS 0.02893f
C1740 VDD1.n133 VSUBS 0.015546f
C1741 VDD1.n134 VSUBS 0.036744f
C1742 VDD1.n135 VSUBS 0.01646f
C1743 VDD1.n136 VSUBS 0.02893f
C1744 VDD1.n137 VSUBS 0.015546f
C1745 VDD1.n138 VSUBS 0.036744f
C1746 VDD1.n139 VSUBS 0.01646f
C1747 VDD1.n140 VSUBS 0.326209f
C1748 VDD1.t8 VSUBS 0.079915f
C1749 VDD1.n141 VSUBS 0.027558f
C1750 VDD1.n142 VSUBS 0.027641f
C1751 VDD1.n143 VSUBS 0.015546f
C1752 VDD1.n144 VSUBS 2.37466f
C1753 VDD1.n145 VSUBS 0.02893f
C1754 VDD1.n146 VSUBS 0.015546f
C1755 VDD1.n147 VSUBS 0.01646f
C1756 VDD1.n148 VSUBS 0.036744f
C1757 VDD1.n149 VSUBS 0.036744f
C1758 VDD1.n150 VSUBS 0.01646f
C1759 VDD1.n151 VSUBS 0.015546f
C1760 VDD1.n152 VSUBS 0.02893f
C1761 VDD1.n153 VSUBS 0.02893f
C1762 VDD1.n154 VSUBS 0.015546f
C1763 VDD1.n155 VSUBS 0.01646f
C1764 VDD1.n156 VSUBS 0.036744f
C1765 VDD1.n157 VSUBS 0.036744f
C1766 VDD1.n158 VSUBS 0.036744f
C1767 VDD1.n159 VSUBS 0.01646f
C1768 VDD1.n160 VSUBS 0.015546f
C1769 VDD1.n161 VSUBS 0.02893f
C1770 VDD1.n162 VSUBS 0.02893f
C1771 VDD1.n163 VSUBS 0.015546f
C1772 VDD1.n164 VSUBS 0.016003f
C1773 VDD1.n165 VSUBS 0.016003f
C1774 VDD1.n166 VSUBS 0.036744f
C1775 VDD1.n167 VSUBS 0.036744f
C1776 VDD1.n168 VSUBS 0.01646f
C1777 VDD1.n169 VSUBS 0.015546f
C1778 VDD1.n170 VSUBS 0.02893f
C1779 VDD1.n171 VSUBS 0.02893f
C1780 VDD1.n172 VSUBS 0.015546f
C1781 VDD1.n173 VSUBS 0.01646f
C1782 VDD1.n174 VSUBS 0.036744f
C1783 VDD1.n175 VSUBS 0.036744f
C1784 VDD1.n176 VSUBS 0.01646f
C1785 VDD1.n177 VSUBS 0.015546f
C1786 VDD1.n178 VSUBS 0.02893f
C1787 VDD1.n179 VSUBS 0.02893f
C1788 VDD1.n180 VSUBS 0.015546f
C1789 VDD1.n181 VSUBS 0.01646f
C1790 VDD1.n182 VSUBS 0.036744f
C1791 VDD1.n183 VSUBS 0.036744f
C1792 VDD1.n184 VSUBS 0.01646f
C1793 VDD1.n185 VSUBS 0.015546f
C1794 VDD1.n186 VSUBS 0.02893f
C1795 VDD1.n187 VSUBS 0.02893f
C1796 VDD1.n188 VSUBS 0.015546f
C1797 VDD1.n189 VSUBS 0.01646f
C1798 VDD1.n190 VSUBS 0.036744f
C1799 VDD1.n191 VSUBS 0.036744f
C1800 VDD1.n192 VSUBS 0.01646f
C1801 VDD1.n193 VSUBS 0.015546f
C1802 VDD1.n194 VSUBS 0.02893f
C1803 VDD1.n195 VSUBS 0.02893f
C1804 VDD1.n196 VSUBS 0.015546f
C1805 VDD1.n197 VSUBS 0.01646f
C1806 VDD1.n198 VSUBS 0.036744f
C1807 VDD1.n199 VSUBS 0.036744f
C1808 VDD1.n200 VSUBS 0.01646f
C1809 VDD1.n201 VSUBS 0.015546f
C1810 VDD1.n202 VSUBS 0.02893f
C1811 VDD1.n203 VSUBS 0.02893f
C1812 VDD1.n204 VSUBS 0.015546f
C1813 VDD1.n205 VSUBS 0.01646f
C1814 VDD1.n206 VSUBS 0.036744f
C1815 VDD1.n207 VSUBS 0.09259f
C1816 VDD1.n208 VSUBS 0.01646f
C1817 VDD1.n209 VSUBS 0.030528f
C1818 VDD1.n210 VSUBS 0.074775f
C1819 VDD1.n211 VSUBS 0.116667f
C1820 VDD1.t3 VSUBS 0.446254f
C1821 VDD1.t0 VSUBS 0.446254f
C1822 VDD1.n212 VSUBS 3.77109f
C1823 VDD1.n213 VSUBS 1.33164f
C1824 VDD1.t2 VSUBS 0.446254f
C1825 VDD1.t1 VSUBS 0.446254f
C1826 VDD1.n214 VSUBS 3.81149f
C1827 VDD1.n215 VSUBS 5.14583f
C1828 VDD1.t4 VSUBS 0.446254f
C1829 VDD1.t5 VSUBS 0.446254f
C1830 VDD1.n216 VSUBS 3.77109f
C1831 VDD1.n217 VSUBS 5.22527f
C1832 VTAIL.t7 VSUBS 0.428729f
C1833 VTAIL.t0 VSUBS 0.428729f
C1834 VTAIL.n0 VSUBS 3.46486f
C1835 VTAIL.n1 VSUBS 1.09626f
C1836 VTAIL.n2 VSUBS 0.030635f
C1837 VTAIL.n3 VSUBS 0.027794f
C1838 VTAIL.n4 VSUBS 0.014935f
C1839 VTAIL.n5 VSUBS 0.035301f
C1840 VTAIL.n6 VSUBS 0.015814f
C1841 VTAIL.n7 VSUBS 0.027794f
C1842 VTAIL.n8 VSUBS 0.014935f
C1843 VTAIL.n9 VSUBS 0.035301f
C1844 VTAIL.n10 VSUBS 0.015814f
C1845 VTAIL.n11 VSUBS 0.027794f
C1846 VTAIL.n12 VSUBS 0.014935f
C1847 VTAIL.n13 VSUBS 0.035301f
C1848 VTAIL.n14 VSUBS 0.015814f
C1849 VTAIL.n15 VSUBS 0.027794f
C1850 VTAIL.n16 VSUBS 0.014935f
C1851 VTAIL.n17 VSUBS 0.035301f
C1852 VTAIL.n18 VSUBS 0.015814f
C1853 VTAIL.n19 VSUBS 0.027794f
C1854 VTAIL.n20 VSUBS 0.014935f
C1855 VTAIL.n21 VSUBS 0.035301f
C1856 VTAIL.n22 VSUBS 0.015814f
C1857 VTAIL.n23 VSUBS 0.027794f
C1858 VTAIL.n24 VSUBS 0.014935f
C1859 VTAIL.n25 VSUBS 0.035301f
C1860 VTAIL.n26 VSUBS 0.015814f
C1861 VTAIL.n27 VSUBS 0.027794f
C1862 VTAIL.n28 VSUBS 0.014935f
C1863 VTAIL.n29 VSUBS 0.035301f
C1864 VTAIL.n30 VSUBS 0.015814f
C1865 VTAIL.n31 VSUBS 0.027794f
C1866 VTAIL.n32 VSUBS 0.014935f
C1867 VTAIL.n33 VSUBS 0.035301f
C1868 VTAIL.n34 VSUBS 0.015814f
C1869 VTAIL.n35 VSUBS 0.313399f
C1870 VTAIL.t16 VSUBS 0.076777f
C1871 VTAIL.n36 VSUBS 0.026476f
C1872 VTAIL.n37 VSUBS 0.026556f
C1873 VTAIL.n38 VSUBS 0.014935f
C1874 VTAIL.n39 VSUBS 2.28141f
C1875 VTAIL.n40 VSUBS 0.027794f
C1876 VTAIL.n41 VSUBS 0.014935f
C1877 VTAIL.n42 VSUBS 0.015814f
C1878 VTAIL.n43 VSUBS 0.035301f
C1879 VTAIL.n44 VSUBS 0.035301f
C1880 VTAIL.n45 VSUBS 0.015814f
C1881 VTAIL.n46 VSUBS 0.014935f
C1882 VTAIL.n47 VSUBS 0.027794f
C1883 VTAIL.n48 VSUBS 0.027794f
C1884 VTAIL.n49 VSUBS 0.014935f
C1885 VTAIL.n50 VSUBS 0.015814f
C1886 VTAIL.n51 VSUBS 0.035301f
C1887 VTAIL.n52 VSUBS 0.035301f
C1888 VTAIL.n53 VSUBS 0.035301f
C1889 VTAIL.n54 VSUBS 0.015814f
C1890 VTAIL.n55 VSUBS 0.014935f
C1891 VTAIL.n56 VSUBS 0.027794f
C1892 VTAIL.n57 VSUBS 0.027794f
C1893 VTAIL.n58 VSUBS 0.014935f
C1894 VTAIL.n59 VSUBS 0.015375f
C1895 VTAIL.n60 VSUBS 0.015375f
C1896 VTAIL.n61 VSUBS 0.035301f
C1897 VTAIL.n62 VSUBS 0.035301f
C1898 VTAIL.n63 VSUBS 0.015814f
C1899 VTAIL.n64 VSUBS 0.014935f
C1900 VTAIL.n65 VSUBS 0.027794f
C1901 VTAIL.n66 VSUBS 0.027794f
C1902 VTAIL.n67 VSUBS 0.014935f
C1903 VTAIL.n68 VSUBS 0.015814f
C1904 VTAIL.n69 VSUBS 0.035301f
C1905 VTAIL.n70 VSUBS 0.035301f
C1906 VTAIL.n71 VSUBS 0.015814f
C1907 VTAIL.n72 VSUBS 0.014935f
C1908 VTAIL.n73 VSUBS 0.027794f
C1909 VTAIL.n74 VSUBS 0.027794f
C1910 VTAIL.n75 VSUBS 0.014935f
C1911 VTAIL.n76 VSUBS 0.015814f
C1912 VTAIL.n77 VSUBS 0.035301f
C1913 VTAIL.n78 VSUBS 0.035301f
C1914 VTAIL.n79 VSUBS 0.015814f
C1915 VTAIL.n80 VSUBS 0.014935f
C1916 VTAIL.n81 VSUBS 0.027794f
C1917 VTAIL.n82 VSUBS 0.027794f
C1918 VTAIL.n83 VSUBS 0.014935f
C1919 VTAIL.n84 VSUBS 0.015814f
C1920 VTAIL.n85 VSUBS 0.035301f
C1921 VTAIL.n86 VSUBS 0.035301f
C1922 VTAIL.n87 VSUBS 0.015814f
C1923 VTAIL.n88 VSUBS 0.014935f
C1924 VTAIL.n89 VSUBS 0.027794f
C1925 VTAIL.n90 VSUBS 0.027794f
C1926 VTAIL.n91 VSUBS 0.014935f
C1927 VTAIL.n92 VSUBS 0.015814f
C1928 VTAIL.n93 VSUBS 0.035301f
C1929 VTAIL.n94 VSUBS 0.035301f
C1930 VTAIL.n95 VSUBS 0.015814f
C1931 VTAIL.n96 VSUBS 0.014935f
C1932 VTAIL.n97 VSUBS 0.027794f
C1933 VTAIL.n98 VSUBS 0.027794f
C1934 VTAIL.n99 VSUBS 0.014935f
C1935 VTAIL.n100 VSUBS 0.015814f
C1936 VTAIL.n101 VSUBS 0.035301f
C1937 VTAIL.n102 VSUBS 0.088954f
C1938 VTAIL.n103 VSUBS 0.015814f
C1939 VTAIL.n104 VSUBS 0.029329f
C1940 VTAIL.n105 VSUBS 0.071838f
C1941 VTAIL.n106 VSUBS 0.068815f
C1942 VTAIL.n107 VSUBS 0.551874f
C1943 VTAIL.t17 VSUBS 0.428729f
C1944 VTAIL.t13 VSUBS 0.428729f
C1945 VTAIL.n108 VSUBS 3.46486f
C1946 VTAIL.n109 VSUBS 1.28986f
C1947 VTAIL.t11 VSUBS 0.428729f
C1948 VTAIL.t12 VSUBS 0.428729f
C1949 VTAIL.n110 VSUBS 3.46486f
C1950 VTAIL.n111 VSUBS 3.49563f
C1951 VTAIL.t1 VSUBS 0.428729f
C1952 VTAIL.t18 VSUBS 0.428729f
C1953 VTAIL.n112 VSUBS 3.46488f
C1954 VTAIL.n113 VSUBS 3.49561f
C1955 VTAIL.t19 VSUBS 0.428729f
C1956 VTAIL.t5 VSUBS 0.428729f
C1957 VTAIL.n114 VSUBS 3.46488f
C1958 VTAIL.n115 VSUBS 1.28984f
C1959 VTAIL.n116 VSUBS 0.030635f
C1960 VTAIL.n117 VSUBS 0.027794f
C1961 VTAIL.n118 VSUBS 0.014935f
C1962 VTAIL.n119 VSUBS 0.035301f
C1963 VTAIL.n120 VSUBS 0.015814f
C1964 VTAIL.n121 VSUBS 0.027794f
C1965 VTAIL.n122 VSUBS 0.014935f
C1966 VTAIL.n123 VSUBS 0.035301f
C1967 VTAIL.n124 VSUBS 0.015814f
C1968 VTAIL.n125 VSUBS 0.027794f
C1969 VTAIL.n126 VSUBS 0.014935f
C1970 VTAIL.n127 VSUBS 0.035301f
C1971 VTAIL.n128 VSUBS 0.015814f
C1972 VTAIL.n129 VSUBS 0.027794f
C1973 VTAIL.n130 VSUBS 0.014935f
C1974 VTAIL.n131 VSUBS 0.035301f
C1975 VTAIL.n132 VSUBS 0.015814f
C1976 VTAIL.n133 VSUBS 0.027794f
C1977 VTAIL.n134 VSUBS 0.014935f
C1978 VTAIL.n135 VSUBS 0.035301f
C1979 VTAIL.n136 VSUBS 0.015814f
C1980 VTAIL.n137 VSUBS 0.027794f
C1981 VTAIL.n138 VSUBS 0.014935f
C1982 VTAIL.n139 VSUBS 0.035301f
C1983 VTAIL.n140 VSUBS 0.015814f
C1984 VTAIL.n141 VSUBS 0.027794f
C1985 VTAIL.n142 VSUBS 0.014935f
C1986 VTAIL.n143 VSUBS 0.035301f
C1987 VTAIL.n144 VSUBS 0.035301f
C1988 VTAIL.n145 VSUBS 0.015814f
C1989 VTAIL.n146 VSUBS 0.027794f
C1990 VTAIL.n147 VSUBS 0.014935f
C1991 VTAIL.n148 VSUBS 0.035301f
C1992 VTAIL.n149 VSUBS 0.015814f
C1993 VTAIL.n150 VSUBS 0.313399f
C1994 VTAIL.t6 VSUBS 0.076777f
C1995 VTAIL.n151 VSUBS 0.026476f
C1996 VTAIL.n152 VSUBS 0.026556f
C1997 VTAIL.n153 VSUBS 0.014935f
C1998 VTAIL.n154 VSUBS 2.28141f
C1999 VTAIL.n155 VSUBS 0.027794f
C2000 VTAIL.n156 VSUBS 0.014935f
C2001 VTAIL.n157 VSUBS 0.015814f
C2002 VTAIL.n158 VSUBS 0.035301f
C2003 VTAIL.n159 VSUBS 0.035301f
C2004 VTAIL.n160 VSUBS 0.015814f
C2005 VTAIL.n161 VSUBS 0.014935f
C2006 VTAIL.n162 VSUBS 0.027794f
C2007 VTAIL.n163 VSUBS 0.027794f
C2008 VTAIL.n164 VSUBS 0.014935f
C2009 VTAIL.n165 VSUBS 0.015814f
C2010 VTAIL.n166 VSUBS 0.035301f
C2011 VTAIL.n167 VSUBS 0.035301f
C2012 VTAIL.n168 VSUBS 0.015814f
C2013 VTAIL.n169 VSUBS 0.014935f
C2014 VTAIL.n170 VSUBS 0.027794f
C2015 VTAIL.n171 VSUBS 0.027794f
C2016 VTAIL.n172 VSUBS 0.014935f
C2017 VTAIL.n173 VSUBS 0.015375f
C2018 VTAIL.n174 VSUBS 0.015375f
C2019 VTAIL.n175 VSUBS 0.035301f
C2020 VTAIL.n176 VSUBS 0.035301f
C2021 VTAIL.n177 VSUBS 0.015814f
C2022 VTAIL.n178 VSUBS 0.014935f
C2023 VTAIL.n179 VSUBS 0.027794f
C2024 VTAIL.n180 VSUBS 0.027794f
C2025 VTAIL.n181 VSUBS 0.014935f
C2026 VTAIL.n182 VSUBS 0.015814f
C2027 VTAIL.n183 VSUBS 0.035301f
C2028 VTAIL.n184 VSUBS 0.035301f
C2029 VTAIL.n185 VSUBS 0.015814f
C2030 VTAIL.n186 VSUBS 0.014935f
C2031 VTAIL.n187 VSUBS 0.027794f
C2032 VTAIL.n188 VSUBS 0.027794f
C2033 VTAIL.n189 VSUBS 0.014935f
C2034 VTAIL.n190 VSUBS 0.015814f
C2035 VTAIL.n191 VSUBS 0.035301f
C2036 VTAIL.n192 VSUBS 0.035301f
C2037 VTAIL.n193 VSUBS 0.015814f
C2038 VTAIL.n194 VSUBS 0.014935f
C2039 VTAIL.n195 VSUBS 0.027794f
C2040 VTAIL.n196 VSUBS 0.027794f
C2041 VTAIL.n197 VSUBS 0.014935f
C2042 VTAIL.n198 VSUBS 0.015814f
C2043 VTAIL.n199 VSUBS 0.035301f
C2044 VTAIL.n200 VSUBS 0.035301f
C2045 VTAIL.n201 VSUBS 0.015814f
C2046 VTAIL.n202 VSUBS 0.014935f
C2047 VTAIL.n203 VSUBS 0.027794f
C2048 VTAIL.n204 VSUBS 0.027794f
C2049 VTAIL.n205 VSUBS 0.014935f
C2050 VTAIL.n206 VSUBS 0.015814f
C2051 VTAIL.n207 VSUBS 0.035301f
C2052 VTAIL.n208 VSUBS 0.035301f
C2053 VTAIL.n209 VSUBS 0.015814f
C2054 VTAIL.n210 VSUBS 0.014935f
C2055 VTAIL.n211 VSUBS 0.027794f
C2056 VTAIL.n212 VSUBS 0.027794f
C2057 VTAIL.n213 VSUBS 0.014935f
C2058 VTAIL.n214 VSUBS 0.015814f
C2059 VTAIL.n215 VSUBS 0.035301f
C2060 VTAIL.n216 VSUBS 0.088954f
C2061 VTAIL.n217 VSUBS 0.015814f
C2062 VTAIL.n218 VSUBS 0.029329f
C2063 VTAIL.n219 VSUBS 0.071838f
C2064 VTAIL.n220 VSUBS 0.068815f
C2065 VTAIL.n221 VSUBS 0.551874f
C2066 VTAIL.t8 VSUBS 0.428729f
C2067 VTAIL.t10 VSUBS 0.428729f
C2068 VTAIL.n222 VSUBS 3.46488f
C2069 VTAIL.n223 VSUBS 1.17133f
C2070 VTAIL.t9 VSUBS 0.428729f
C2071 VTAIL.t14 VSUBS 0.428729f
C2072 VTAIL.n224 VSUBS 3.46488f
C2073 VTAIL.n225 VSUBS 1.28984f
C2074 VTAIL.n226 VSUBS 0.030635f
C2075 VTAIL.n227 VSUBS 0.027794f
C2076 VTAIL.n228 VSUBS 0.014935f
C2077 VTAIL.n229 VSUBS 0.035301f
C2078 VTAIL.n230 VSUBS 0.015814f
C2079 VTAIL.n231 VSUBS 0.027794f
C2080 VTAIL.n232 VSUBS 0.014935f
C2081 VTAIL.n233 VSUBS 0.035301f
C2082 VTAIL.n234 VSUBS 0.015814f
C2083 VTAIL.n235 VSUBS 0.027794f
C2084 VTAIL.n236 VSUBS 0.014935f
C2085 VTAIL.n237 VSUBS 0.035301f
C2086 VTAIL.n238 VSUBS 0.015814f
C2087 VTAIL.n239 VSUBS 0.027794f
C2088 VTAIL.n240 VSUBS 0.014935f
C2089 VTAIL.n241 VSUBS 0.035301f
C2090 VTAIL.n242 VSUBS 0.015814f
C2091 VTAIL.n243 VSUBS 0.027794f
C2092 VTAIL.n244 VSUBS 0.014935f
C2093 VTAIL.n245 VSUBS 0.035301f
C2094 VTAIL.n246 VSUBS 0.015814f
C2095 VTAIL.n247 VSUBS 0.027794f
C2096 VTAIL.n248 VSUBS 0.014935f
C2097 VTAIL.n249 VSUBS 0.035301f
C2098 VTAIL.n250 VSUBS 0.015814f
C2099 VTAIL.n251 VSUBS 0.027794f
C2100 VTAIL.n252 VSUBS 0.014935f
C2101 VTAIL.n253 VSUBS 0.035301f
C2102 VTAIL.n254 VSUBS 0.035301f
C2103 VTAIL.n255 VSUBS 0.015814f
C2104 VTAIL.n256 VSUBS 0.027794f
C2105 VTAIL.n257 VSUBS 0.014935f
C2106 VTAIL.n258 VSUBS 0.035301f
C2107 VTAIL.n259 VSUBS 0.015814f
C2108 VTAIL.n260 VSUBS 0.313399f
C2109 VTAIL.t15 VSUBS 0.076777f
C2110 VTAIL.n261 VSUBS 0.026476f
C2111 VTAIL.n262 VSUBS 0.026556f
C2112 VTAIL.n263 VSUBS 0.014935f
C2113 VTAIL.n264 VSUBS 2.28141f
C2114 VTAIL.n265 VSUBS 0.027794f
C2115 VTAIL.n266 VSUBS 0.014935f
C2116 VTAIL.n267 VSUBS 0.015814f
C2117 VTAIL.n268 VSUBS 0.035301f
C2118 VTAIL.n269 VSUBS 0.035301f
C2119 VTAIL.n270 VSUBS 0.015814f
C2120 VTAIL.n271 VSUBS 0.014935f
C2121 VTAIL.n272 VSUBS 0.027794f
C2122 VTAIL.n273 VSUBS 0.027794f
C2123 VTAIL.n274 VSUBS 0.014935f
C2124 VTAIL.n275 VSUBS 0.015814f
C2125 VTAIL.n276 VSUBS 0.035301f
C2126 VTAIL.n277 VSUBS 0.035301f
C2127 VTAIL.n278 VSUBS 0.015814f
C2128 VTAIL.n279 VSUBS 0.014935f
C2129 VTAIL.n280 VSUBS 0.027794f
C2130 VTAIL.n281 VSUBS 0.027794f
C2131 VTAIL.n282 VSUBS 0.014935f
C2132 VTAIL.n283 VSUBS 0.015375f
C2133 VTAIL.n284 VSUBS 0.015375f
C2134 VTAIL.n285 VSUBS 0.035301f
C2135 VTAIL.n286 VSUBS 0.035301f
C2136 VTAIL.n287 VSUBS 0.015814f
C2137 VTAIL.n288 VSUBS 0.014935f
C2138 VTAIL.n289 VSUBS 0.027794f
C2139 VTAIL.n290 VSUBS 0.027794f
C2140 VTAIL.n291 VSUBS 0.014935f
C2141 VTAIL.n292 VSUBS 0.015814f
C2142 VTAIL.n293 VSUBS 0.035301f
C2143 VTAIL.n294 VSUBS 0.035301f
C2144 VTAIL.n295 VSUBS 0.015814f
C2145 VTAIL.n296 VSUBS 0.014935f
C2146 VTAIL.n297 VSUBS 0.027794f
C2147 VTAIL.n298 VSUBS 0.027794f
C2148 VTAIL.n299 VSUBS 0.014935f
C2149 VTAIL.n300 VSUBS 0.015814f
C2150 VTAIL.n301 VSUBS 0.035301f
C2151 VTAIL.n302 VSUBS 0.035301f
C2152 VTAIL.n303 VSUBS 0.015814f
C2153 VTAIL.n304 VSUBS 0.014935f
C2154 VTAIL.n305 VSUBS 0.027794f
C2155 VTAIL.n306 VSUBS 0.027794f
C2156 VTAIL.n307 VSUBS 0.014935f
C2157 VTAIL.n308 VSUBS 0.015814f
C2158 VTAIL.n309 VSUBS 0.035301f
C2159 VTAIL.n310 VSUBS 0.035301f
C2160 VTAIL.n311 VSUBS 0.015814f
C2161 VTAIL.n312 VSUBS 0.014935f
C2162 VTAIL.n313 VSUBS 0.027794f
C2163 VTAIL.n314 VSUBS 0.027794f
C2164 VTAIL.n315 VSUBS 0.014935f
C2165 VTAIL.n316 VSUBS 0.015814f
C2166 VTAIL.n317 VSUBS 0.035301f
C2167 VTAIL.n318 VSUBS 0.035301f
C2168 VTAIL.n319 VSUBS 0.015814f
C2169 VTAIL.n320 VSUBS 0.014935f
C2170 VTAIL.n321 VSUBS 0.027794f
C2171 VTAIL.n322 VSUBS 0.027794f
C2172 VTAIL.n323 VSUBS 0.014935f
C2173 VTAIL.n324 VSUBS 0.015814f
C2174 VTAIL.n325 VSUBS 0.035301f
C2175 VTAIL.n326 VSUBS 0.088954f
C2176 VTAIL.n327 VSUBS 0.015814f
C2177 VTAIL.n328 VSUBS 0.029329f
C2178 VTAIL.n329 VSUBS 0.071838f
C2179 VTAIL.n330 VSUBS 0.068815f
C2180 VTAIL.n331 VSUBS 2.55498f
C2181 VTAIL.n332 VSUBS 0.030635f
C2182 VTAIL.n333 VSUBS 0.027794f
C2183 VTAIL.n334 VSUBS 0.014935f
C2184 VTAIL.n335 VSUBS 0.035301f
C2185 VTAIL.n336 VSUBS 0.015814f
C2186 VTAIL.n337 VSUBS 0.027794f
C2187 VTAIL.n338 VSUBS 0.014935f
C2188 VTAIL.n339 VSUBS 0.035301f
C2189 VTAIL.n340 VSUBS 0.015814f
C2190 VTAIL.n341 VSUBS 0.027794f
C2191 VTAIL.n342 VSUBS 0.014935f
C2192 VTAIL.n343 VSUBS 0.035301f
C2193 VTAIL.n344 VSUBS 0.015814f
C2194 VTAIL.n345 VSUBS 0.027794f
C2195 VTAIL.n346 VSUBS 0.014935f
C2196 VTAIL.n347 VSUBS 0.035301f
C2197 VTAIL.n348 VSUBS 0.015814f
C2198 VTAIL.n349 VSUBS 0.027794f
C2199 VTAIL.n350 VSUBS 0.014935f
C2200 VTAIL.n351 VSUBS 0.035301f
C2201 VTAIL.n352 VSUBS 0.015814f
C2202 VTAIL.n353 VSUBS 0.027794f
C2203 VTAIL.n354 VSUBS 0.014935f
C2204 VTAIL.n355 VSUBS 0.035301f
C2205 VTAIL.n356 VSUBS 0.015814f
C2206 VTAIL.n357 VSUBS 0.027794f
C2207 VTAIL.n358 VSUBS 0.014935f
C2208 VTAIL.n359 VSUBS 0.035301f
C2209 VTAIL.n360 VSUBS 0.015814f
C2210 VTAIL.n361 VSUBS 0.027794f
C2211 VTAIL.n362 VSUBS 0.014935f
C2212 VTAIL.n363 VSUBS 0.035301f
C2213 VTAIL.n364 VSUBS 0.015814f
C2214 VTAIL.n365 VSUBS 0.313399f
C2215 VTAIL.t2 VSUBS 0.076777f
C2216 VTAIL.n366 VSUBS 0.026476f
C2217 VTAIL.n367 VSUBS 0.026556f
C2218 VTAIL.n368 VSUBS 0.014935f
C2219 VTAIL.n369 VSUBS 2.28141f
C2220 VTAIL.n370 VSUBS 0.027794f
C2221 VTAIL.n371 VSUBS 0.014935f
C2222 VTAIL.n372 VSUBS 0.015814f
C2223 VTAIL.n373 VSUBS 0.035301f
C2224 VTAIL.n374 VSUBS 0.035301f
C2225 VTAIL.n375 VSUBS 0.015814f
C2226 VTAIL.n376 VSUBS 0.014935f
C2227 VTAIL.n377 VSUBS 0.027794f
C2228 VTAIL.n378 VSUBS 0.027794f
C2229 VTAIL.n379 VSUBS 0.014935f
C2230 VTAIL.n380 VSUBS 0.015814f
C2231 VTAIL.n381 VSUBS 0.035301f
C2232 VTAIL.n382 VSUBS 0.035301f
C2233 VTAIL.n383 VSUBS 0.035301f
C2234 VTAIL.n384 VSUBS 0.015814f
C2235 VTAIL.n385 VSUBS 0.014935f
C2236 VTAIL.n386 VSUBS 0.027794f
C2237 VTAIL.n387 VSUBS 0.027794f
C2238 VTAIL.n388 VSUBS 0.014935f
C2239 VTAIL.n389 VSUBS 0.015375f
C2240 VTAIL.n390 VSUBS 0.015375f
C2241 VTAIL.n391 VSUBS 0.035301f
C2242 VTAIL.n392 VSUBS 0.035301f
C2243 VTAIL.n393 VSUBS 0.015814f
C2244 VTAIL.n394 VSUBS 0.014935f
C2245 VTAIL.n395 VSUBS 0.027794f
C2246 VTAIL.n396 VSUBS 0.027794f
C2247 VTAIL.n397 VSUBS 0.014935f
C2248 VTAIL.n398 VSUBS 0.015814f
C2249 VTAIL.n399 VSUBS 0.035301f
C2250 VTAIL.n400 VSUBS 0.035301f
C2251 VTAIL.n401 VSUBS 0.015814f
C2252 VTAIL.n402 VSUBS 0.014935f
C2253 VTAIL.n403 VSUBS 0.027794f
C2254 VTAIL.n404 VSUBS 0.027794f
C2255 VTAIL.n405 VSUBS 0.014935f
C2256 VTAIL.n406 VSUBS 0.015814f
C2257 VTAIL.n407 VSUBS 0.035301f
C2258 VTAIL.n408 VSUBS 0.035301f
C2259 VTAIL.n409 VSUBS 0.015814f
C2260 VTAIL.n410 VSUBS 0.014935f
C2261 VTAIL.n411 VSUBS 0.027794f
C2262 VTAIL.n412 VSUBS 0.027794f
C2263 VTAIL.n413 VSUBS 0.014935f
C2264 VTAIL.n414 VSUBS 0.015814f
C2265 VTAIL.n415 VSUBS 0.035301f
C2266 VTAIL.n416 VSUBS 0.035301f
C2267 VTAIL.n417 VSUBS 0.015814f
C2268 VTAIL.n418 VSUBS 0.014935f
C2269 VTAIL.n419 VSUBS 0.027794f
C2270 VTAIL.n420 VSUBS 0.027794f
C2271 VTAIL.n421 VSUBS 0.014935f
C2272 VTAIL.n422 VSUBS 0.015814f
C2273 VTAIL.n423 VSUBS 0.035301f
C2274 VTAIL.n424 VSUBS 0.035301f
C2275 VTAIL.n425 VSUBS 0.015814f
C2276 VTAIL.n426 VSUBS 0.014935f
C2277 VTAIL.n427 VSUBS 0.027794f
C2278 VTAIL.n428 VSUBS 0.027794f
C2279 VTAIL.n429 VSUBS 0.014935f
C2280 VTAIL.n430 VSUBS 0.015814f
C2281 VTAIL.n431 VSUBS 0.035301f
C2282 VTAIL.n432 VSUBS 0.088954f
C2283 VTAIL.n433 VSUBS 0.015814f
C2284 VTAIL.n434 VSUBS 0.029329f
C2285 VTAIL.n435 VSUBS 0.071838f
C2286 VTAIL.n436 VSUBS 0.068815f
C2287 VTAIL.n437 VSUBS 2.55498f
C2288 VTAIL.t4 VSUBS 0.428729f
C2289 VTAIL.t3 VSUBS 0.428729f
C2290 VTAIL.n438 VSUBS 3.46486f
C2291 VTAIL.n439 VSUBS 1.04376f
C2292 VP.t8 VSUBS 4.35424f
C2293 VP.n0 VSUBS 1.57599f
C2294 VP.n1 VSUBS 0.021143f
C2295 VP.n2 VSUBS 0.041997f
C2296 VP.n3 VSUBS 0.021143f
C2297 VP.n4 VSUBS 0.039208f
C2298 VP.n5 VSUBS 0.021143f
C2299 VP.t7 VSUBS 4.35424f
C2300 VP.n6 VSUBS 0.039208f
C2301 VP.n7 VSUBS 0.021143f
C2302 VP.n8 VSUBS 0.039208f
C2303 VP.n9 VSUBS 0.021143f
C2304 VP.t9 VSUBS 4.35424f
C2305 VP.n10 VSUBS 0.039208f
C2306 VP.n11 VSUBS 0.021143f
C2307 VP.n12 VSUBS 0.039208f
C2308 VP.n13 VSUBS 0.021143f
C2309 VP.t6 VSUBS 4.35424f
C2310 VP.n14 VSUBS 0.039208f
C2311 VP.n15 VSUBS 0.021143f
C2312 VP.n16 VSUBS 0.039208f
C2313 VP.n17 VSUBS 0.034119f
C2314 VP.t1 VSUBS 4.35424f
C2315 VP.t4 VSUBS 4.35424f
C2316 VP.n18 VSUBS 1.57599f
C2317 VP.n19 VSUBS 0.021143f
C2318 VP.n20 VSUBS 0.041997f
C2319 VP.n21 VSUBS 0.021143f
C2320 VP.n22 VSUBS 0.039208f
C2321 VP.n23 VSUBS 0.021143f
C2322 VP.t5 VSUBS 4.35424f
C2323 VP.n24 VSUBS 0.039208f
C2324 VP.n25 VSUBS 0.021143f
C2325 VP.n26 VSUBS 0.039208f
C2326 VP.n27 VSUBS 0.021143f
C2327 VP.t2 VSUBS 4.35424f
C2328 VP.n28 VSUBS 0.039208f
C2329 VP.n29 VSUBS 0.021143f
C2330 VP.n30 VSUBS 0.039208f
C2331 VP.t0 VSUBS 4.70745f
C2332 VP.n31 VSUBS 1.50591f
C2333 VP.t3 VSUBS 4.35424f
C2334 VP.n32 VSUBS 1.5783f
C2335 VP.n33 VSUBS 0.035724f
C2336 VP.n34 VSUBS 0.272055f
C2337 VP.n35 VSUBS 0.021143f
C2338 VP.n36 VSUBS 0.021143f
C2339 VP.n37 VSUBS 0.039208f
C2340 VP.n38 VSUBS 0.026055f
C2341 VP.n39 VSUBS 0.035415f
C2342 VP.n40 VSUBS 0.021143f
C2343 VP.n41 VSUBS 0.021143f
C2344 VP.n42 VSUBS 0.021143f
C2345 VP.n43 VSUBS 0.039208f
C2346 VP.n44 VSUBS 0.02953f
C2347 VP.n45 VSUBS 1.49598f
C2348 VP.n46 VSUBS 0.02953f
C2349 VP.n47 VSUBS 0.021143f
C2350 VP.n48 VSUBS 0.021143f
C2351 VP.n49 VSUBS 0.021143f
C2352 VP.n50 VSUBS 0.039208f
C2353 VP.n51 VSUBS 0.035415f
C2354 VP.n52 VSUBS 0.026055f
C2355 VP.n53 VSUBS 0.021143f
C2356 VP.n54 VSUBS 0.021143f
C2357 VP.n55 VSUBS 0.021143f
C2358 VP.n56 VSUBS 0.039208f
C2359 VP.n57 VSUBS 0.035724f
C2360 VP.n58 VSUBS 1.49598f
C2361 VP.n59 VSUBS 0.023336f
C2362 VP.n60 VSUBS 0.021143f
C2363 VP.n61 VSUBS 0.021143f
C2364 VP.n62 VSUBS 0.021143f
C2365 VP.n63 VSUBS 0.039208f
C2366 VP.n64 VSUBS 0.041578f
C2367 VP.n65 VSUBS 0.017104f
C2368 VP.n66 VSUBS 0.021143f
C2369 VP.n67 VSUBS 0.021143f
C2370 VP.n68 VSUBS 0.021143f
C2371 VP.n69 VSUBS 0.039208f
C2372 VP.n70 VSUBS 0.039208f
C2373 VP.n71 VSUBS 0.022562f
C2374 VP.n72 VSUBS 0.034119f
C2375 VP.n73 VSUBS 1.75462f
C2376 VP.n74 VSUBS 1.76625f
C2377 VP.n75 VSUBS 1.57599f
C2378 VP.n76 VSUBS 0.022562f
C2379 VP.n77 VSUBS 0.039208f
C2380 VP.n78 VSUBS 0.021143f
C2381 VP.n79 VSUBS 0.021143f
C2382 VP.n80 VSUBS 0.021143f
C2383 VP.n81 VSUBS 0.041997f
C2384 VP.n82 VSUBS 0.017104f
C2385 VP.n83 VSUBS 0.041578f
C2386 VP.n84 VSUBS 0.021143f
C2387 VP.n85 VSUBS 0.021143f
C2388 VP.n86 VSUBS 0.021143f
C2389 VP.n87 VSUBS 0.039208f
C2390 VP.n88 VSUBS 0.023336f
C2391 VP.n89 VSUBS 1.49598f
C2392 VP.n90 VSUBS 0.035724f
C2393 VP.n91 VSUBS 0.021143f
C2394 VP.n92 VSUBS 0.021143f
C2395 VP.n93 VSUBS 0.021143f
C2396 VP.n94 VSUBS 0.039208f
C2397 VP.n95 VSUBS 0.026055f
C2398 VP.n96 VSUBS 0.035415f
C2399 VP.n97 VSUBS 0.021143f
C2400 VP.n98 VSUBS 0.021143f
C2401 VP.n99 VSUBS 0.021143f
C2402 VP.n100 VSUBS 0.039208f
C2403 VP.n101 VSUBS 0.02953f
C2404 VP.n102 VSUBS 1.49598f
C2405 VP.n103 VSUBS 0.02953f
C2406 VP.n104 VSUBS 0.021143f
C2407 VP.n105 VSUBS 0.021143f
C2408 VP.n106 VSUBS 0.021143f
C2409 VP.n107 VSUBS 0.039208f
C2410 VP.n108 VSUBS 0.035415f
C2411 VP.n109 VSUBS 0.026055f
C2412 VP.n110 VSUBS 0.021143f
C2413 VP.n111 VSUBS 0.021143f
C2414 VP.n112 VSUBS 0.021143f
C2415 VP.n113 VSUBS 0.039208f
C2416 VP.n114 VSUBS 0.035724f
C2417 VP.n115 VSUBS 1.49598f
C2418 VP.n116 VSUBS 0.023336f
C2419 VP.n117 VSUBS 0.021143f
C2420 VP.n118 VSUBS 0.021143f
C2421 VP.n119 VSUBS 0.021143f
C2422 VP.n120 VSUBS 0.039208f
C2423 VP.n121 VSUBS 0.041578f
C2424 VP.n122 VSUBS 0.017104f
C2425 VP.n123 VSUBS 0.021143f
C2426 VP.n124 VSUBS 0.021143f
C2427 VP.n125 VSUBS 0.021143f
C2428 VP.n126 VSUBS 0.039208f
C2429 VP.n127 VSUBS 0.039208f
C2430 VP.n128 VSUBS 0.022562f
C2431 VP.n129 VSUBS 0.034119f
C2432 VP.n130 VSUBS 0.064869f
.ends

