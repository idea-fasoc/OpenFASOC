* NGSPICE file created from diff_pair_sample_1567.ext - technology: sky130A

.subckt diff_pair_sample_1567 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t1 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=1.188 ps=7.53 w=7.2 l=2.2
X1 VTAIL.t0 VP.t0 VDD1.t3 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=1.188 ps=7.53 w=7.2 l=2.2
X2 B.t11 B.t9 B.t10 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=0 ps=0 w=7.2 l=2.2
X3 VTAIL.t6 VN.t1 VDD2.t0 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=1.188 ps=7.53 w=7.2 l=2.2
X4 VDD1.t2 VP.t1 VTAIL.t3 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=1.188 pd=7.53 as=2.808 ps=15.18 w=7.2 l=2.2
X5 B.t8 B.t6 B.t7 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=0 ps=0 w=7.2 l=2.2
X6 VDD2.t3 VN.t2 VTAIL.t5 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=1.188 pd=7.53 as=2.808 ps=15.18 w=7.2 l=2.2
X7 VDD1.t1 VP.t2 VTAIL.t1 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=1.188 pd=7.53 as=2.808 ps=15.18 w=7.2 l=2.2
X8 B.t5 B.t3 B.t4 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=0 ps=0 w=7.2 l=2.2
X9 B.t2 B.t0 B.t1 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=0 ps=0 w=7.2 l=2.2
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=1.188 pd=7.53 as=2.808 ps=15.18 w=7.2 l=2.2
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2488_n2408# sky130_fd_pr__pfet_01v8 ad=2.808 pd=15.18 as=1.188 ps=7.53 w=7.2 l=2.2
R0 VN.n0 VN.t1 114.632
R1 VN.n1 VN.t2 114.632
R2 VN.n0 VN.t3 113.996
R3 VN.n1 VN.t0 113.996
R4 VN VN.n1 47.4734
R5 VN VN.n0 5.82565
R6 VDD2.n2 VDD2.n0 123.63
R7 VDD2.n2 VDD2.n1 87.166
R8 VDD2.n1 VDD2.t1 4.51508
R9 VDD2.n1 VDD2.t3 4.51508
R10 VDD2.n0 VDD2.t0 4.51508
R11 VDD2.n0 VDD2.t2 4.51508
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n265 VTAIL.n264 585
R14 VTAIL.n267 VTAIL.n266 585
R15 VTAIL.n260 VTAIL.n259 585
R16 VTAIL.n273 VTAIL.n272 585
R17 VTAIL.n275 VTAIL.n274 585
R18 VTAIL.n256 VTAIL.n255 585
R19 VTAIL.n281 VTAIL.n280 585
R20 VTAIL.n283 VTAIL.n282 585
R21 VTAIL.n13 VTAIL.n12 585
R22 VTAIL.n15 VTAIL.n14 585
R23 VTAIL.n8 VTAIL.n7 585
R24 VTAIL.n21 VTAIL.n20 585
R25 VTAIL.n23 VTAIL.n22 585
R26 VTAIL.n4 VTAIL.n3 585
R27 VTAIL.n29 VTAIL.n28 585
R28 VTAIL.n31 VTAIL.n30 585
R29 VTAIL.n49 VTAIL.n48 585
R30 VTAIL.n51 VTAIL.n50 585
R31 VTAIL.n44 VTAIL.n43 585
R32 VTAIL.n57 VTAIL.n56 585
R33 VTAIL.n59 VTAIL.n58 585
R34 VTAIL.n40 VTAIL.n39 585
R35 VTAIL.n65 VTAIL.n64 585
R36 VTAIL.n67 VTAIL.n66 585
R37 VTAIL.n85 VTAIL.n84 585
R38 VTAIL.n87 VTAIL.n86 585
R39 VTAIL.n80 VTAIL.n79 585
R40 VTAIL.n93 VTAIL.n92 585
R41 VTAIL.n95 VTAIL.n94 585
R42 VTAIL.n76 VTAIL.n75 585
R43 VTAIL.n101 VTAIL.n100 585
R44 VTAIL.n103 VTAIL.n102 585
R45 VTAIL.n247 VTAIL.n246 585
R46 VTAIL.n245 VTAIL.n244 585
R47 VTAIL.n220 VTAIL.n219 585
R48 VTAIL.n239 VTAIL.n238 585
R49 VTAIL.n237 VTAIL.n236 585
R50 VTAIL.n224 VTAIL.n223 585
R51 VTAIL.n231 VTAIL.n230 585
R52 VTAIL.n229 VTAIL.n228 585
R53 VTAIL.n211 VTAIL.n210 585
R54 VTAIL.n209 VTAIL.n208 585
R55 VTAIL.n184 VTAIL.n183 585
R56 VTAIL.n203 VTAIL.n202 585
R57 VTAIL.n201 VTAIL.n200 585
R58 VTAIL.n188 VTAIL.n187 585
R59 VTAIL.n195 VTAIL.n194 585
R60 VTAIL.n193 VTAIL.n192 585
R61 VTAIL.n175 VTAIL.n174 585
R62 VTAIL.n173 VTAIL.n172 585
R63 VTAIL.n148 VTAIL.n147 585
R64 VTAIL.n167 VTAIL.n166 585
R65 VTAIL.n165 VTAIL.n164 585
R66 VTAIL.n152 VTAIL.n151 585
R67 VTAIL.n159 VTAIL.n158 585
R68 VTAIL.n157 VTAIL.n156 585
R69 VTAIL.n139 VTAIL.n138 585
R70 VTAIL.n137 VTAIL.n136 585
R71 VTAIL.n112 VTAIL.n111 585
R72 VTAIL.n131 VTAIL.n130 585
R73 VTAIL.n129 VTAIL.n128 585
R74 VTAIL.n116 VTAIL.n115 585
R75 VTAIL.n123 VTAIL.n122 585
R76 VTAIL.n121 VTAIL.n120 585
R77 VTAIL.n282 VTAIL.n252 498.474
R78 VTAIL.n30 VTAIL.n0 498.474
R79 VTAIL.n66 VTAIL.n36 498.474
R80 VTAIL.n102 VTAIL.n72 498.474
R81 VTAIL.n246 VTAIL.n216 498.474
R82 VTAIL.n210 VTAIL.n180 498.474
R83 VTAIL.n174 VTAIL.n144 498.474
R84 VTAIL.n138 VTAIL.n108 498.474
R85 VTAIL.n263 VTAIL.t4 329.053
R86 VTAIL.n11 VTAIL.t6 329.053
R87 VTAIL.n47 VTAIL.t3 329.053
R88 VTAIL.n83 VTAIL.t2 329.053
R89 VTAIL.n227 VTAIL.t1 329.053
R90 VTAIL.n191 VTAIL.t0 329.053
R91 VTAIL.n155 VTAIL.t5 329.053
R92 VTAIL.n119 VTAIL.t7 329.053
R93 VTAIL.n266 VTAIL.n265 171.744
R94 VTAIL.n266 VTAIL.n259 171.744
R95 VTAIL.n273 VTAIL.n259 171.744
R96 VTAIL.n274 VTAIL.n273 171.744
R97 VTAIL.n274 VTAIL.n255 171.744
R98 VTAIL.n281 VTAIL.n255 171.744
R99 VTAIL.n282 VTAIL.n281 171.744
R100 VTAIL.n14 VTAIL.n13 171.744
R101 VTAIL.n14 VTAIL.n7 171.744
R102 VTAIL.n21 VTAIL.n7 171.744
R103 VTAIL.n22 VTAIL.n21 171.744
R104 VTAIL.n22 VTAIL.n3 171.744
R105 VTAIL.n29 VTAIL.n3 171.744
R106 VTAIL.n30 VTAIL.n29 171.744
R107 VTAIL.n50 VTAIL.n49 171.744
R108 VTAIL.n50 VTAIL.n43 171.744
R109 VTAIL.n57 VTAIL.n43 171.744
R110 VTAIL.n58 VTAIL.n57 171.744
R111 VTAIL.n58 VTAIL.n39 171.744
R112 VTAIL.n65 VTAIL.n39 171.744
R113 VTAIL.n66 VTAIL.n65 171.744
R114 VTAIL.n86 VTAIL.n85 171.744
R115 VTAIL.n86 VTAIL.n79 171.744
R116 VTAIL.n93 VTAIL.n79 171.744
R117 VTAIL.n94 VTAIL.n93 171.744
R118 VTAIL.n94 VTAIL.n75 171.744
R119 VTAIL.n101 VTAIL.n75 171.744
R120 VTAIL.n102 VTAIL.n101 171.744
R121 VTAIL.n246 VTAIL.n245 171.744
R122 VTAIL.n245 VTAIL.n219 171.744
R123 VTAIL.n238 VTAIL.n219 171.744
R124 VTAIL.n238 VTAIL.n237 171.744
R125 VTAIL.n237 VTAIL.n223 171.744
R126 VTAIL.n230 VTAIL.n223 171.744
R127 VTAIL.n230 VTAIL.n229 171.744
R128 VTAIL.n210 VTAIL.n209 171.744
R129 VTAIL.n209 VTAIL.n183 171.744
R130 VTAIL.n202 VTAIL.n183 171.744
R131 VTAIL.n202 VTAIL.n201 171.744
R132 VTAIL.n201 VTAIL.n187 171.744
R133 VTAIL.n194 VTAIL.n187 171.744
R134 VTAIL.n194 VTAIL.n193 171.744
R135 VTAIL.n174 VTAIL.n173 171.744
R136 VTAIL.n173 VTAIL.n147 171.744
R137 VTAIL.n166 VTAIL.n147 171.744
R138 VTAIL.n166 VTAIL.n165 171.744
R139 VTAIL.n165 VTAIL.n151 171.744
R140 VTAIL.n158 VTAIL.n151 171.744
R141 VTAIL.n158 VTAIL.n157 171.744
R142 VTAIL.n138 VTAIL.n137 171.744
R143 VTAIL.n137 VTAIL.n111 171.744
R144 VTAIL.n130 VTAIL.n111 171.744
R145 VTAIL.n130 VTAIL.n129 171.744
R146 VTAIL.n129 VTAIL.n115 171.744
R147 VTAIL.n122 VTAIL.n115 171.744
R148 VTAIL.n122 VTAIL.n121 171.744
R149 VTAIL.n265 VTAIL.t4 85.8723
R150 VTAIL.n13 VTAIL.t6 85.8723
R151 VTAIL.n49 VTAIL.t3 85.8723
R152 VTAIL.n85 VTAIL.t2 85.8723
R153 VTAIL.n229 VTAIL.t1 85.8723
R154 VTAIL.n193 VTAIL.t0 85.8723
R155 VTAIL.n157 VTAIL.t5 85.8723
R156 VTAIL.n121 VTAIL.t7 85.8723
R157 VTAIL.n287 VTAIL.n286 34.5126
R158 VTAIL.n35 VTAIL.n34 34.5126
R159 VTAIL.n71 VTAIL.n70 34.5126
R160 VTAIL.n107 VTAIL.n106 34.5126
R161 VTAIL.n251 VTAIL.n250 34.5126
R162 VTAIL.n215 VTAIL.n214 34.5126
R163 VTAIL.n179 VTAIL.n178 34.5126
R164 VTAIL.n143 VTAIL.n142 34.5126
R165 VTAIL.n287 VTAIL.n251 20.7548
R166 VTAIL.n143 VTAIL.n107 20.7548
R167 VTAIL.n284 VTAIL.n283 12.8005
R168 VTAIL.n32 VTAIL.n31 12.8005
R169 VTAIL.n68 VTAIL.n67 12.8005
R170 VTAIL.n104 VTAIL.n103 12.8005
R171 VTAIL.n248 VTAIL.n247 12.8005
R172 VTAIL.n212 VTAIL.n211 12.8005
R173 VTAIL.n176 VTAIL.n175 12.8005
R174 VTAIL.n140 VTAIL.n139 12.8005
R175 VTAIL.n280 VTAIL.n254 12.0247
R176 VTAIL.n28 VTAIL.n2 12.0247
R177 VTAIL.n64 VTAIL.n38 12.0247
R178 VTAIL.n100 VTAIL.n74 12.0247
R179 VTAIL.n244 VTAIL.n218 12.0247
R180 VTAIL.n208 VTAIL.n182 12.0247
R181 VTAIL.n172 VTAIL.n146 12.0247
R182 VTAIL.n136 VTAIL.n110 12.0247
R183 VTAIL.n279 VTAIL.n256 11.249
R184 VTAIL.n27 VTAIL.n4 11.249
R185 VTAIL.n63 VTAIL.n40 11.249
R186 VTAIL.n99 VTAIL.n76 11.249
R187 VTAIL.n243 VTAIL.n220 11.249
R188 VTAIL.n207 VTAIL.n184 11.249
R189 VTAIL.n171 VTAIL.n148 11.249
R190 VTAIL.n135 VTAIL.n112 11.249
R191 VTAIL.n264 VTAIL.n263 10.7237
R192 VTAIL.n12 VTAIL.n11 10.7237
R193 VTAIL.n48 VTAIL.n47 10.7237
R194 VTAIL.n84 VTAIL.n83 10.7237
R195 VTAIL.n228 VTAIL.n227 10.7237
R196 VTAIL.n192 VTAIL.n191 10.7237
R197 VTAIL.n156 VTAIL.n155 10.7237
R198 VTAIL.n120 VTAIL.n119 10.7237
R199 VTAIL.n276 VTAIL.n275 10.4732
R200 VTAIL.n24 VTAIL.n23 10.4732
R201 VTAIL.n60 VTAIL.n59 10.4732
R202 VTAIL.n96 VTAIL.n95 10.4732
R203 VTAIL.n240 VTAIL.n239 10.4732
R204 VTAIL.n204 VTAIL.n203 10.4732
R205 VTAIL.n168 VTAIL.n167 10.4732
R206 VTAIL.n132 VTAIL.n131 10.4732
R207 VTAIL.n272 VTAIL.n258 9.69747
R208 VTAIL.n20 VTAIL.n6 9.69747
R209 VTAIL.n56 VTAIL.n42 9.69747
R210 VTAIL.n92 VTAIL.n78 9.69747
R211 VTAIL.n236 VTAIL.n222 9.69747
R212 VTAIL.n200 VTAIL.n186 9.69747
R213 VTAIL.n164 VTAIL.n150 9.69747
R214 VTAIL.n128 VTAIL.n114 9.69747
R215 VTAIL.n286 VTAIL.n285 9.45567
R216 VTAIL.n34 VTAIL.n33 9.45567
R217 VTAIL.n70 VTAIL.n69 9.45567
R218 VTAIL.n106 VTAIL.n105 9.45567
R219 VTAIL.n250 VTAIL.n249 9.45567
R220 VTAIL.n214 VTAIL.n213 9.45567
R221 VTAIL.n178 VTAIL.n177 9.45567
R222 VTAIL.n142 VTAIL.n141 9.45567
R223 VTAIL.n262 VTAIL.n261 9.3005
R224 VTAIL.n269 VTAIL.n268 9.3005
R225 VTAIL.n271 VTAIL.n270 9.3005
R226 VTAIL.n258 VTAIL.n257 9.3005
R227 VTAIL.n277 VTAIL.n276 9.3005
R228 VTAIL.n279 VTAIL.n278 9.3005
R229 VTAIL.n254 VTAIL.n253 9.3005
R230 VTAIL.n285 VTAIL.n284 9.3005
R231 VTAIL.n10 VTAIL.n9 9.3005
R232 VTAIL.n17 VTAIL.n16 9.3005
R233 VTAIL.n19 VTAIL.n18 9.3005
R234 VTAIL.n6 VTAIL.n5 9.3005
R235 VTAIL.n25 VTAIL.n24 9.3005
R236 VTAIL.n27 VTAIL.n26 9.3005
R237 VTAIL.n2 VTAIL.n1 9.3005
R238 VTAIL.n33 VTAIL.n32 9.3005
R239 VTAIL.n46 VTAIL.n45 9.3005
R240 VTAIL.n53 VTAIL.n52 9.3005
R241 VTAIL.n55 VTAIL.n54 9.3005
R242 VTAIL.n42 VTAIL.n41 9.3005
R243 VTAIL.n61 VTAIL.n60 9.3005
R244 VTAIL.n63 VTAIL.n62 9.3005
R245 VTAIL.n38 VTAIL.n37 9.3005
R246 VTAIL.n69 VTAIL.n68 9.3005
R247 VTAIL.n82 VTAIL.n81 9.3005
R248 VTAIL.n89 VTAIL.n88 9.3005
R249 VTAIL.n91 VTAIL.n90 9.3005
R250 VTAIL.n78 VTAIL.n77 9.3005
R251 VTAIL.n97 VTAIL.n96 9.3005
R252 VTAIL.n99 VTAIL.n98 9.3005
R253 VTAIL.n74 VTAIL.n73 9.3005
R254 VTAIL.n105 VTAIL.n104 9.3005
R255 VTAIL.n226 VTAIL.n225 9.3005
R256 VTAIL.n233 VTAIL.n232 9.3005
R257 VTAIL.n235 VTAIL.n234 9.3005
R258 VTAIL.n222 VTAIL.n221 9.3005
R259 VTAIL.n241 VTAIL.n240 9.3005
R260 VTAIL.n243 VTAIL.n242 9.3005
R261 VTAIL.n218 VTAIL.n217 9.3005
R262 VTAIL.n249 VTAIL.n248 9.3005
R263 VTAIL.n190 VTAIL.n189 9.3005
R264 VTAIL.n197 VTAIL.n196 9.3005
R265 VTAIL.n199 VTAIL.n198 9.3005
R266 VTAIL.n186 VTAIL.n185 9.3005
R267 VTAIL.n205 VTAIL.n204 9.3005
R268 VTAIL.n207 VTAIL.n206 9.3005
R269 VTAIL.n182 VTAIL.n181 9.3005
R270 VTAIL.n213 VTAIL.n212 9.3005
R271 VTAIL.n154 VTAIL.n153 9.3005
R272 VTAIL.n161 VTAIL.n160 9.3005
R273 VTAIL.n163 VTAIL.n162 9.3005
R274 VTAIL.n150 VTAIL.n149 9.3005
R275 VTAIL.n169 VTAIL.n168 9.3005
R276 VTAIL.n171 VTAIL.n170 9.3005
R277 VTAIL.n146 VTAIL.n145 9.3005
R278 VTAIL.n177 VTAIL.n176 9.3005
R279 VTAIL.n118 VTAIL.n117 9.3005
R280 VTAIL.n125 VTAIL.n124 9.3005
R281 VTAIL.n127 VTAIL.n126 9.3005
R282 VTAIL.n114 VTAIL.n113 9.3005
R283 VTAIL.n133 VTAIL.n132 9.3005
R284 VTAIL.n135 VTAIL.n134 9.3005
R285 VTAIL.n110 VTAIL.n109 9.3005
R286 VTAIL.n141 VTAIL.n140 9.3005
R287 VTAIL.n271 VTAIL.n260 8.92171
R288 VTAIL.n19 VTAIL.n8 8.92171
R289 VTAIL.n55 VTAIL.n44 8.92171
R290 VTAIL.n91 VTAIL.n80 8.92171
R291 VTAIL.n235 VTAIL.n224 8.92171
R292 VTAIL.n199 VTAIL.n188 8.92171
R293 VTAIL.n163 VTAIL.n152 8.92171
R294 VTAIL.n127 VTAIL.n116 8.92171
R295 VTAIL.n268 VTAIL.n267 8.14595
R296 VTAIL.n16 VTAIL.n15 8.14595
R297 VTAIL.n52 VTAIL.n51 8.14595
R298 VTAIL.n88 VTAIL.n87 8.14595
R299 VTAIL.n232 VTAIL.n231 8.14595
R300 VTAIL.n196 VTAIL.n195 8.14595
R301 VTAIL.n160 VTAIL.n159 8.14595
R302 VTAIL.n124 VTAIL.n123 8.14595
R303 VTAIL.n286 VTAIL.n252 7.75445
R304 VTAIL.n34 VTAIL.n0 7.75445
R305 VTAIL.n70 VTAIL.n36 7.75445
R306 VTAIL.n106 VTAIL.n72 7.75445
R307 VTAIL.n250 VTAIL.n216 7.75445
R308 VTAIL.n214 VTAIL.n180 7.75445
R309 VTAIL.n178 VTAIL.n144 7.75445
R310 VTAIL.n142 VTAIL.n108 7.75445
R311 VTAIL.n264 VTAIL.n262 7.3702
R312 VTAIL.n12 VTAIL.n10 7.3702
R313 VTAIL.n48 VTAIL.n46 7.3702
R314 VTAIL.n84 VTAIL.n82 7.3702
R315 VTAIL.n228 VTAIL.n226 7.3702
R316 VTAIL.n192 VTAIL.n190 7.3702
R317 VTAIL.n156 VTAIL.n154 7.3702
R318 VTAIL.n120 VTAIL.n118 7.3702
R319 VTAIL.n284 VTAIL.n252 6.08283
R320 VTAIL.n32 VTAIL.n0 6.08283
R321 VTAIL.n68 VTAIL.n36 6.08283
R322 VTAIL.n104 VTAIL.n72 6.08283
R323 VTAIL.n248 VTAIL.n216 6.08283
R324 VTAIL.n212 VTAIL.n180 6.08283
R325 VTAIL.n176 VTAIL.n144 6.08283
R326 VTAIL.n140 VTAIL.n108 6.08283
R327 VTAIL.n267 VTAIL.n262 5.81868
R328 VTAIL.n15 VTAIL.n10 5.81868
R329 VTAIL.n51 VTAIL.n46 5.81868
R330 VTAIL.n87 VTAIL.n82 5.81868
R331 VTAIL.n231 VTAIL.n226 5.81868
R332 VTAIL.n195 VTAIL.n190 5.81868
R333 VTAIL.n159 VTAIL.n154 5.81868
R334 VTAIL.n123 VTAIL.n118 5.81868
R335 VTAIL.n268 VTAIL.n260 5.04292
R336 VTAIL.n16 VTAIL.n8 5.04292
R337 VTAIL.n52 VTAIL.n44 5.04292
R338 VTAIL.n88 VTAIL.n80 5.04292
R339 VTAIL.n232 VTAIL.n224 5.04292
R340 VTAIL.n196 VTAIL.n188 5.04292
R341 VTAIL.n160 VTAIL.n152 5.04292
R342 VTAIL.n124 VTAIL.n116 5.04292
R343 VTAIL.n272 VTAIL.n271 4.26717
R344 VTAIL.n20 VTAIL.n19 4.26717
R345 VTAIL.n56 VTAIL.n55 4.26717
R346 VTAIL.n92 VTAIL.n91 4.26717
R347 VTAIL.n236 VTAIL.n235 4.26717
R348 VTAIL.n200 VTAIL.n199 4.26717
R349 VTAIL.n164 VTAIL.n163 4.26717
R350 VTAIL.n128 VTAIL.n127 4.26717
R351 VTAIL.n275 VTAIL.n258 3.49141
R352 VTAIL.n23 VTAIL.n6 3.49141
R353 VTAIL.n59 VTAIL.n42 3.49141
R354 VTAIL.n95 VTAIL.n78 3.49141
R355 VTAIL.n239 VTAIL.n222 3.49141
R356 VTAIL.n203 VTAIL.n186 3.49141
R357 VTAIL.n167 VTAIL.n150 3.49141
R358 VTAIL.n131 VTAIL.n114 3.49141
R359 VTAIL.n276 VTAIL.n256 2.71565
R360 VTAIL.n24 VTAIL.n4 2.71565
R361 VTAIL.n60 VTAIL.n40 2.71565
R362 VTAIL.n96 VTAIL.n76 2.71565
R363 VTAIL.n240 VTAIL.n220 2.71565
R364 VTAIL.n204 VTAIL.n184 2.71565
R365 VTAIL.n168 VTAIL.n148 2.71565
R366 VTAIL.n132 VTAIL.n112 2.71565
R367 VTAIL.n263 VTAIL.n261 2.41305
R368 VTAIL.n11 VTAIL.n9 2.41305
R369 VTAIL.n47 VTAIL.n45 2.41305
R370 VTAIL.n83 VTAIL.n81 2.41305
R371 VTAIL.n227 VTAIL.n225 2.41305
R372 VTAIL.n191 VTAIL.n189 2.41305
R373 VTAIL.n155 VTAIL.n153 2.41305
R374 VTAIL.n119 VTAIL.n117 2.41305
R375 VTAIL.n179 VTAIL.n143 2.18153
R376 VTAIL.n251 VTAIL.n215 2.18153
R377 VTAIL.n107 VTAIL.n71 2.18153
R378 VTAIL.n280 VTAIL.n279 1.93989
R379 VTAIL.n28 VTAIL.n27 1.93989
R380 VTAIL.n64 VTAIL.n63 1.93989
R381 VTAIL.n100 VTAIL.n99 1.93989
R382 VTAIL.n244 VTAIL.n243 1.93989
R383 VTAIL.n208 VTAIL.n207 1.93989
R384 VTAIL.n172 VTAIL.n171 1.93989
R385 VTAIL.n136 VTAIL.n135 1.93989
R386 VTAIL.n283 VTAIL.n254 1.16414
R387 VTAIL.n31 VTAIL.n2 1.16414
R388 VTAIL.n67 VTAIL.n38 1.16414
R389 VTAIL.n103 VTAIL.n74 1.16414
R390 VTAIL.n247 VTAIL.n218 1.16414
R391 VTAIL.n211 VTAIL.n182 1.16414
R392 VTAIL.n175 VTAIL.n146 1.16414
R393 VTAIL.n139 VTAIL.n110 1.16414
R394 VTAIL VTAIL.n35 1.14921
R395 VTAIL VTAIL.n287 1.03283
R396 VTAIL.n215 VTAIL.n179 0.470328
R397 VTAIL.n71 VTAIL.n35 0.470328
R398 VTAIL.n269 VTAIL.n261 0.155672
R399 VTAIL.n270 VTAIL.n269 0.155672
R400 VTAIL.n270 VTAIL.n257 0.155672
R401 VTAIL.n277 VTAIL.n257 0.155672
R402 VTAIL.n278 VTAIL.n277 0.155672
R403 VTAIL.n278 VTAIL.n253 0.155672
R404 VTAIL.n285 VTAIL.n253 0.155672
R405 VTAIL.n17 VTAIL.n9 0.155672
R406 VTAIL.n18 VTAIL.n17 0.155672
R407 VTAIL.n18 VTAIL.n5 0.155672
R408 VTAIL.n25 VTAIL.n5 0.155672
R409 VTAIL.n26 VTAIL.n25 0.155672
R410 VTAIL.n26 VTAIL.n1 0.155672
R411 VTAIL.n33 VTAIL.n1 0.155672
R412 VTAIL.n53 VTAIL.n45 0.155672
R413 VTAIL.n54 VTAIL.n53 0.155672
R414 VTAIL.n54 VTAIL.n41 0.155672
R415 VTAIL.n61 VTAIL.n41 0.155672
R416 VTAIL.n62 VTAIL.n61 0.155672
R417 VTAIL.n62 VTAIL.n37 0.155672
R418 VTAIL.n69 VTAIL.n37 0.155672
R419 VTAIL.n89 VTAIL.n81 0.155672
R420 VTAIL.n90 VTAIL.n89 0.155672
R421 VTAIL.n90 VTAIL.n77 0.155672
R422 VTAIL.n97 VTAIL.n77 0.155672
R423 VTAIL.n98 VTAIL.n97 0.155672
R424 VTAIL.n98 VTAIL.n73 0.155672
R425 VTAIL.n105 VTAIL.n73 0.155672
R426 VTAIL.n249 VTAIL.n217 0.155672
R427 VTAIL.n242 VTAIL.n217 0.155672
R428 VTAIL.n242 VTAIL.n241 0.155672
R429 VTAIL.n241 VTAIL.n221 0.155672
R430 VTAIL.n234 VTAIL.n221 0.155672
R431 VTAIL.n234 VTAIL.n233 0.155672
R432 VTAIL.n233 VTAIL.n225 0.155672
R433 VTAIL.n213 VTAIL.n181 0.155672
R434 VTAIL.n206 VTAIL.n181 0.155672
R435 VTAIL.n206 VTAIL.n205 0.155672
R436 VTAIL.n205 VTAIL.n185 0.155672
R437 VTAIL.n198 VTAIL.n185 0.155672
R438 VTAIL.n198 VTAIL.n197 0.155672
R439 VTAIL.n197 VTAIL.n189 0.155672
R440 VTAIL.n177 VTAIL.n145 0.155672
R441 VTAIL.n170 VTAIL.n145 0.155672
R442 VTAIL.n170 VTAIL.n169 0.155672
R443 VTAIL.n169 VTAIL.n149 0.155672
R444 VTAIL.n162 VTAIL.n149 0.155672
R445 VTAIL.n162 VTAIL.n161 0.155672
R446 VTAIL.n161 VTAIL.n153 0.155672
R447 VTAIL.n141 VTAIL.n109 0.155672
R448 VTAIL.n134 VTAIL.n109 0.155672
R449 VTAIL.n134 VTAIL.n133 0.155672
R450 VTAIL.n133 VTAIL.n113 0.155672
R451 VTAIL.n126 VTAIL.n113 0.155672
R452 VTAIL.n126 VTAIL.n125 0.155672
R453 VTAIL.n125 VTAIL.n117 0.155672
R454 VP.n12 VP.n0 161.3
R455 VP.n11 VP.n10 161.3
R456 VP.n9 VP.n1 161.3
R457 VP.n8 VP.n7 161.3
R458 VP.n6 VP.n2 161.3
R459 VP.n3 VP.t0 114.632
R460 VP.n3 VP.t2 113.996
R461 VP.n5 VP.n4 97.8746
R462 VP.n14 VP.n13 97.8746
R463 VP.n5 VP.t3 78.8732
R464 VP.n13 VP.t1 78.8732
R465 VP.n4 VP.n3 47.1945
R466 VP.n7 VP.n1 40.577
R467 VP.n11 VP.n1 40.577
R468 VP.n7 VP.n6 24.5923
R469 VP.n12 VP.n11 24.5923
R470 VP.n6 VP.n5 13.0342
R471 VP.n13 VP.n12 13.0342
R472 VP.n4 VP.n2 0.278335
R473 VP.n14 VP.n0 0.278335
R474 VP.n8 VP.n2 0.189894
R475 VP.n9 VP.n8 0.189894
R476 VP.n10 VP.n9 0.189894
R477 VP.n10 VP.n0 0.189894
R478 VP VP.n14 0.153485
R479 VDD1 VDD1.n1 124.156
R480 VDD1 VDD1.n0 87.2242
R481 VDD1.n0 VDD1.t3 4.51508
R482 VDD1.n0 VDD1.t1 4.51508
R483 VDD1.n1 VDD1.t0 4.51508
R484 VDD1.n1 VDD1.t2 4.51508
R485 B.n278 B.n277 585
R486 B.n276 B.n85 585
R487 B.n275 B.n274 585
R488 B.n273 B.n86 585
R489 B.n272 B.n271 585
R490 B.n270 B.n87 585
R491 B.n269 B.n268 585
R492 B.n267 B.n88 585
R493 B.n266 B.n265 585
R494 B.n264 B.n89 585
R495 B.n263 B.n262 585
R496 B.n261 B.n90 585
R497 B.n260 B.n259 585
R498 B.n258 B.n91 585
R499 B.n257 B.n256 585
R500 B.n255 B.n92 585
R501 B.n254 B.n253 585
R502 B.n252 B.n93 585
R503 B.n251 B.n250 585
R504 B.n249 B.n94 585
R505 B.n248 B.n247 585
R506 B.n246 B.n95 585
R507 B.n245 B.n244 585
R508 B.n243 B.n96 585
R509 B.n242 B.n241 585
R510 B.n240 B.n97 585
R511 B.n239 B.n238 585
R512 B.n237 B.n98 585
R513 B.n236 B.n235 585
R514 B.n231 B.n99 585
R515 B.n230 B.n229 585
R516 B.n228 B.n100 585
R517 B.n227 B.n226 585
R518 B.n225 B.n101 585
R519 B.n224 B.n223 585
R520 B.n222 B.n102 585
R521 B.n221 B.n220 585
R522 B.n218 B.n103 585
R523 B.n217 B.n216 585
R524 B.n215 B.n106 585
R525 B.n214 B.n213 585
R526 B.n212 B.n107 585
R527 B.n211 B.n210 585
R528 B.n209 B.n108 585
R529 B.n208 B.n207 585
R530 B.n206 B.n109 585
R531 B.n205 B.n204 585
R532 B.n203 B.n110 585
R533 B.n202 B.n201 585
R534 B.n200 B.n111 585
R535 B.n199 B.n198 585
R536 B.n197 B.n112 585
R537 B.n196 B.n195 585
R538 B.n194 B.n113 585
R539 B.n193 B.n192 585
R540 B.n191 B.n114 585
R541 B.n190 B.n189 585
R542 B.n188 B.n115 585
R543 B.n187 B.n186 585
R544 B.n185 B.n116 585
R545 B.n184 B.n183 585
R546 B.n182 B.n117 585
R547 B.n181 B.n180 585
R548 B.n179 B.n118 585
R549 B.n178 B.n177 585
R550 B.n279 B.n84 585
R551 B.n281 B.n280 585
R552 B.n282 B.n83 585
R553 B.n284 B.n283 585
R554 B.n285 B.n82 585
R555 B.n287 B.n286 585
R556 B.n288 B.n81 585
R557 B.n290 B.n289 585
R558 B.n291 B.n80 585
R559 B.n293 B.n292 585
R560 B.n294 B.n79 585
R561 B.n296 B.n295 585
R562 B.n297 B.n78 585
R563 B.n299 B.n298 585
R564 B.n300 B.n77 585
R565 B.n302 B.n301 585
R566 B.n303 B.n76 585
R567 B.n305 B.n304 585
R568 B.n306 B.n75 585
R569 B.n308 B.n307 585
R570 B.n309 B.n74 585
R571 B.n311 B.n310 585
R572 B.n312 B.n73 585
R573 B.n314 B.n313 585
R574 B.n315 B.n72 585
R575 B.n317 B.n316 585
R576 B.n318 B.n71 585
R577 B.n320 B.n319 585
R578 B.n321 B.n70 585
R579 B.n323 B.n322 585
R580 B.n324 B.n69 585
R581 B.n326 B.n325 585
R582 B.n327 B.n68 585
R583 B.n329 B.n328 585
R584 B.n330 B.n67 585
R585 B.n332 B.n331 585
R586 B.n333 B.n66 585
R587 B.n335 B.n334 585
R588 B.n336 B.n65 585
R589 B.n338 B.n337 585
R590 B.n339 B.n64 585
R591 B.n341 B.n340 585
R592 B.n342 B.n63 585
R593 B.n344 B.n343 585
R594 B.n345 B.n62 585
R595 B.n347 B.n346 585
R596 B.n348 B.n61 585
R597 B.n350 B.n349 585
R598 B.n351 B.n60 585
R599 B.n353 B.n352 585
R600 B.n354 B.n59 585
R601 B.n356 B.n355 585
R602 B.n357 B.n58 585
R603 B.n359 B.n358 585
R604 B.n360 B.n57 585
R605 B.n362 B.n361 585
R606 B.n363 B.n56 585
R607 B.n365 B.n364 585
R608 B.n366 B.n55 585
R609 B.n368 B.n367 585
R610 B.n369 B.n54 585
R611 B.n371 B.n370 585
R612 B.n470 B.n17 585
R613 B.n469 B.n468 585
R614 B.n467 B.n18 585
R615 B.n466 B.n465 585
R616 B.n464 B.n19 585
R617 B.n463 B.n462 585
R618 B.n461 B.n20 585
R619 B.n460 B.n459 585
R620 B.n458 B.n21 585
R621 B.n457 B.n456 585
R622 B.n455 B.n22 585
R623 B.n454 B.n453 585
R624 B.n452 B.n23 585
R625 B.n451 B.n450 585
R626 B.n449 B.n24 585
R627 B.n448 B.n447 585
R628 B.n446 B.n25 585
R629 B.n445 B.n444 585
R630 B.n443 B.n26 585
R631 B.n442 B.n441 585
R632 B.n440 B.n27 585
R633 B.n439 B.n438 585
R634 B.n437 B.n28 585
R635 B.n436 B.n435 585
R636 B.n434 B.n29 585
R637 B.n433 B.n432 585
R638 B.n431 B.n30 585
R639 B.n430 B.n429 585
R640 B.n427 B.n31 585
R641 B.n426 B.n425 585
R642 B.n424 B.n34 585
R643 B.n423 B.n422 585
R644 B.n421 B.n35 585
R645 B.n420 B.n419 585
R646 B.n418 B.n36 585
R647 B.n417 B.n416 585
R648 B.n415 B.n37 585
R649 B.n413 B.n412 585
R650 B.n411 B.n40 585
R651 B.n410 B.n409 585
R652 B.n408 B.n41 585
R653 B.n407 B.n406 585
R654 B.n405 B.n42 585
R655 B.n404 B.n403 585
R656 B.n402 B.n43 585
R657 B.n401 B.n400 585
R658 B.n399 B.n44 585
R659 B.n398 B.n397 585
R660 B.n396 B.n45 585
R661 B.n395 B.n394 585
R662 B.n393 B.n46 585
R663 B.n392 B.n391 585
R664 B.n390 B.n47 585
R665 B.n389 B.n388 585
R666 B.n387 B.n48 585
R667 B.n386 B.n385 585
R668 B.n384 B.n49 585
R669 B.n383 B.n382 585
R670 B.n381 B.n50 585
R671 B.n380 B.n379 585
R672 B.n378 B.n51 585
R673 B.n377 B.n376 585
R674 B.n375 B.n52 585
R675 B.n374 B.n373 585
R676 B.n372 B.n53 585
R677 B.n472 B.n471 585
R678 B.n473 B.n16 585
R679 B.n475 B.n474 585
R680 B.n476 B.n15 585
R681 B.n478 B.n477 585
R682 B.n479 B.n14 585
R683 B.n481 B.n480 585
R684 B.n482 B.n13 585
R685 B.n484 B.n483 585
R686 B.n485 B.n12 585
R687 B.n487 B.n486 585
R688 B.n488 B.n11 585
R689 B.n490 B.n489 585
R690 B.n491 B.n10 585
R691 B.n493 B.n492 585
R692 B.n494 B.n9 585
R693 B.n496 B.n495 585
R694 B.n497 B.n8 585
R695 B.n499 B.n498 585
R696 B.n500 B.n7 585
R697 B.n502 B.n501 585
R698 B.n503 B.n6 585
R699 B.n505 B.n504 585
R700 B.n506 B.n5 585
R701 B.n508 B.n507 585
R702 B.n509 B.n4 585
R703 B.n511 B.n510 585
R704 B.n512 B.n3 585
R705 B.n514 B.n513 585
R706 B.n515 B.n0 585
R707 B.n2 B.n1 585
R708 B.n134 B.n133 585
R709 B.n136 B.n135 585
R710 B.n137 B.n132 585
R711 B.n139 B.n138 585
R712 B.n140 B.n131 585
R713 B.n142 B.n141 585
R714 B.n143 B.n130 585
R715 B.n145 B.n144 585
R716 B.n146 B.n129 585
R717 B.n148 B.n147 585
R718 B.n149 B.n128 585
R719 B.n151 B.n150 585
R720 B.n152 B.n127 585
R721 B.n154 B.n153 585
R722 B.n155 B.n126 585
R723 B.n157 B.n156 585
R724 B.n158 B.n125 585
R725 B.n160 B.n159 585
R726 B.n161 B.n124 585
R727 B.n163 B.n162 585
R728 B.n164 B.n123 585
R729 B.n166 B.n165 585
R730 B.n167 B.n122 585
R731 B.n169 B.n168 585
R732 B.n170 B.n121 585
R733 B.n172 B.n171 585
R734 B.n173 B.n120 585
R735 B.n175 B.n174 585
R736 B.n176 B.n119 585
R737 B.n178 B.n119 454.062
R738 B.n279 B.n278 454.062
R739 B.n370 B.n53 454.062
R740 B.n472 B.n17 454.062
R741 B.n232 B.t4 338.26
R742 B.n38 B.t8 338.26
R743 B.n104 B.t1 338.26
R744 B.n32 B.t11 338.26
R745 B.n233 B.t5 289.192
R746 B.n39 B.t7 289.192
R747 B.n105 B.t2 289.192
R748 B.n33 B.t10 289.192
R749 B.n104 B.t0 286.224
R750 B.n232 B.t3 286.224
R751 B.n38 B.t6 286.224
R752 B.n32 B.t9 286.224
R753 B.n517 B.n516 256.663
R754 B.n516 B.n515 235.042
R755 B.n516 B.n2 235.042
R756 B.n179 B.n178 163.367
R757 B.n180 B.n179 163.367
R758 B.n180 B.n117 163.367
R759 B.n184 B.n117 163.367
R760 B.n185 B.n184 163.367
R761 B.n186 B.n185 163.367
R762 B.n186 B.n115 163.367
R763 B.n190 B.n115 163.367
R764 B.n191 B.n190 163.367
R765 B.n192 B.n191 163.367
R766 B.n192 B.n113 163.367
R767 B.n196 B.n113 163.367
R768 B.n197 B.n196 163.367
R769 B.n198 B.n197 163.367
R770 B.n198 B.n111 163.367
R771 B.n202 B.n111 163.367
R772 B.n203 B.n202 163.367
R773 B.n204 B.n203 163.367
R774 B.n204 B.n109 163.367
R775 B.n208 B.n109 163.367
R776 B.n209 B.n208 163.367
R777 B.n210 B.n209 163.367
R778 B.n210 B.n107 163.367
R779 B.n214 B.n107 163.367
R780 B.n215 B.n214 163.367
R781 B.n216 B.n215 163.367
R782 B.n216 B.n103 163.367
R783 B.n221 B.n103 163.367
R784 B.n222 B.n221 163.367
R785 B.n223 B.n222 163.367
R786 B.n223 B.n101 163.367
R787 B.n227 B.n101 163.367
R788 B.n228 B.n227 163.367
R789 B.n229 B.n228 163.367
R790 B.n229 B.n99 163.367
R791 B.n236 B.n99 163.367
R792 B.n237 B.n236 163.367
R793 B.n238 B.n237 163.367
R794 B.n238 B.n97 163.367
R795 B.n242 B.n97 163.367
R796 B.n243 B.n242 163.367
R797 B.n244 B.n243 163.367
R798 B.n244 B.n95 163.367
R799 B.n248 B.n95 163.367
R800 B.n249 B.n248 163.367
R801 B.n250 B.n249 163.367
R802 B.n250 B.n93 163.367
R803 B.n254 B.n93 163.367
R804 B.n255 B.n254 163.367
R805 B.n256 B.n255 163.367
R806 B.n256 B.n91 163.367
R807 B.n260 B.n91 163.367
R808 B.n261 B.n260 163.367
R809 B.n262 B.n261 163.367
R810 B.n262 B.n89 163.367
R811 B.n266 B.n89 163.367
R812 B.n267 B.n266 163.367
R813 B.n268 B.n267 163.367
R814 B.n268 B.n87 163.367
R815 B.n272 B.n87 163.367
R816 B.n273 B.n272 163.367
R817 B.n274 B.n273 163.367
R818 B.n274 B.n85 163.367
R819 B.n278 B.n85 163.367
R820 B.n370 B.n369 163.367
R821 B.n369 B.n368 163.367
R822 B.n368 B.n55 163.367
R823 B.n364 B.n55 163.367
R824 B.n364 B.n363 163.367
R825 B.n363 B.n362 163.367
R826 B.n362 B.n57 163.367
R827 B.n358 B.n57 163.367
R828 B.n358 B.n357 163.367
R829 B.n357 B.n356 163.367
R830 B.n356 B.n59 163.367
R831 B.n352 B.n59 163.367
R832 B.n352 B.n351 163.367
R833 B.n351 B.n350 163.367
R834 B.n350 B.n61 163.367
R835 B.n346 B.n61 163.367
R836 B.n346 B.n345 163.367
R837 B.n345 B.n344 163.367
R838 B.n344 B.n63 163.367
R839 B.n340 B.n63 163.367
R840 B.n340 B.n339 163.367
R841 B.n339 B.n338 163.367
R842 B.n338 B.n65 163.367
R843 B.n334 B.n65 163.367
R844 B.n334 B.n333 163.367
R845 B.n333 B.n332 163.367
R846 B.n332 B.n67 163.367
R847 B.n328 B.n67 163.367
R848 B.n328 B.n327 163.367
R849 B.n327 B.n326 163.367
R850 B.n326 B.n69 163.367
R851 B.n322 B.n69 163.367
R852 B.n322 B.n321 163.367
R853 B.n321 B.n320 163.367
R854 B.n320 B.n71 163.367
R855 B.n316 B.n71 163.367
R856 B.n316 B.n315 163.367
R857 B.n315 B.n314 163.367
R858 B.n314 B.n73 163.367
R859 B.n310 B.n73 163.367
R860 B.n310 B.n309 163.367
R861 B.n309 B.n308 163.367
R862 B.n308 B.n75 163.367
R863 B.n304 B.n75 163.367
R864 B.n304 B.n303 163.367
R865 B.n303 B.n302 163.367
R866 B.n302 B.n77 163.367
R867 B.n298 B.n77 163.367
R868 B.n298 B.n297 163.367
R869 B.n297 B.n296 163.367
R870 B.n296 B.n79 163.367
R871 B.n292 B.n79 163.367
R872 B.n292 B.n291 163.367
R873 B.n291 B.n290 163.367
R874 B.n290 B.n81 163.367
R875 B.n286 B.n81 163.367
R876 B.n286 B.n285 163.367
R877 B.n285 B.n284 163.367
R878 B.n284 B.n83 163.367
R879 B.n280 B.n83 163.367
R880 B.n280 B.n279 163.367
R881 B.n468 B.n17 163.367
R882 B.n468 B.n467 163.367
R883 B.n467 B.n466 163.367
R884 B.n466 B.n19 163.367
R885 B.n462 B.n19 163.367
R886 B.n462 B.n461 163.367
R887 B.n461 B.n460 163.367
R888 B.n460 B.n21 163.367
R889 B.n456 B.n21 163.367
R890 B.n456 B.n455 163.367
R891 B.n455 B.n454 163.367
R892 B.n454 B.n23 163.367
R893 B.n450 B.n23 163.367
R894 B.n450 B.n449 163.367
R895 B.n449 B.n448 163.367
R896 B.n448 B.n25 163.367
R897 B.n444 B.n25 163.367
R898 B.n444 B.n443 163.367
R899 B.n443 B.n442 163.367
R900 B.n442 B.n27 163.367
R901 B.n438 B.n27 163.367
R902 B.n438 B.n437 163.367
R903 B.n437 B.n436 163.367
R904 B.n436 B.n29 163.367
R905 B.n432 B.n29 163.367
R906 B.n432 B.n431 163.367
R907 B.n431 B.n430 163.367
R908 B.n430 B.n31 163.367
R909 B.n425 B.n31 163.367
R910 B.n425 B.n424 163.367
R911 B.n424 B.n423 163.367
R912 B.n423 B.n35 163.367
R913 B.n419 B.n35 163.367
R914 B.n419 B.n418 163.367
R915 B.n418 B.n417 163.367
R916 B.n417 B.n37 163.367
R917 B.n412 B.n37 163.367
R918 B.n412 B.n411 163.367
R919 B.n411 B.n410 163.367
R920 B.n410 B.n41 163.367
R921 B.n406 B.n41 163.367
R922 B.n406 B.n405 163.367
R923 B.n405 B.n404 163.367
R924 B.n404 B.n43 163.367
R925 B.n400 B.n43 163.367
R926 B.n400 B.n399 163.367
R927 B.n399 B.n398 163.367
R928 B.n398 B.n45 163.367
R929 B.n394 B.n45 163.367
R930 B.n394 B.n393 163.367
R931 B.n393 B.n392 163.367
R932 B.n392 B.n47 163.367
R933 B.n388 B.n47 163.367
R934 B.n388 B.n387 163.367
R935 B.n387 B.n386 163.367
R936 B.n386 B.n49 163.367
R937 B.n382 B.n49 163.367
R938 B.n382 B.n381 163.367
R939 B.n381 B.n380 163.367
R940 B.n380 B.n51 163.367
R941 B.n376 B.n51 163.367
R942 B.n376 B.n375 163.367
R943 B.n375 B.n374 163.367
R944 B.n374 B.n53 163.367
R945 B.n473 B.n472 163.367
R946 B.n474 B.n473 163.367
R947 B.n474 B.n15 163.367
R948 B.n478 B.n15 163.367
R949 B.n479 B.n478 163.367
R950 B.n480 B.n479 163.367
R951 B.n480 B.n13 163.367
R952 B.n484 B.n13 163.367
R953 B.n485 B.n484 163.367
R954 B.n486 B.n485 163.367
R955 B.n486 B.n11 163.367
R956 B.n490 B.n11 163.367
R957 B.n491 B.n490 163.367
R958 B.n492 B.n491 163.367
R959 B.n492 B.n9 163.367
R960 B.n496 B.n9 163.367
R961 B.n497 B.n496 163.367
R962 B.n498 B.n497 163.367
R963 B.n498 B.n7 163.367
R964 B.n502 B.n7 163.367
R965 B.n503 B.n502 163.367
R966 B.n504 B.n503 163.367
R967 B.n504 B.n5 163.367
R968 B.n508 B.n5 163.367
R969 B.n509 B.n508 163.367
R970 B.n510 B.n509 163.367
R971 B.n510 B.n3 163.367
R972 B.n514 B.n3 163.367
R973 B.n515 B.n514 163.367
R974 B.n133 B.n2 163.367
R975 B.n136 B.n133 163.367
R976 B.n137 B.n136 163.367
R977 B.n138 B.n137 163.367
R978 B.n138 B.n131 163.367
R979 B.n142 B.n131 163.367
R980 B.n143 B.n142 163.367
R981 B.n144 B.n143 163.367
R982 B.n144 B.n129 163.367
R983 B.n148 B.n129 163.367
R984 B.n149 B.n148 163.367
R985 B.n150 B.n149 163.367
R986 B.n150 B.n127 163.367
R987 B.n154 B.n127 163.367
R988 B.n155 B.n154 163.367
R989 B.n156 B.n155 163.367
R990 B.n156 B.n125 163.367
R991 B.n160 B.n125 163.367
R992 B.n161 B.n160 163.367
R993 B.n162 B.n161 163.367
R994 B.n162 B.n123 163.367
R995 B.n166 B.n123 163.367
R996 B.n167 B.n166 163.367
R997 B.n168 B.n167 163.367
R998 B.n168 B.n121 163.367
R999 B.n172 B.n121 163.367
R1000 B.n173 B.n172 163.367
R1001 B.n174 B.n173 163.367
R1002 B.n174 B.n119 163.367
R1003 B.n219 B.n105 59.5399
R1004 B.n234 B.n233 59.5399
R1005 B.n414 B.n39 59.5399
R1006 B.n428 B.n33 59.5399
R1007 B.n105 B.n104 49.0672
R1008 B.n233 B.n232 49.0672
R1009 B.n39 B.n38 49.0672
R1010 B.n33 B.n32 49.0672
R1011 B.n277 B.n84 29.5029
R1012 B.n471 B.n470 29.5029
R1013 B.n372 B.n371 29.5029
R1014 B.n177 B.n176 29.5029
R1015 B B.n517 18.0485
R1016 B.n471 B.n16 10.6151
R1017 B.n475 B.n16 10.6151
R1018 B.n476 B.n475 10.6151
R1019 B.n477 B.n476 10.6151
R1020 B.n477 B.n14 10.6151
R1021 B.n481 B.n14 10.6151
R1022 B.n482 B.n481 10.6151
R1023 B.n483 B.n482 10.6151
R1024 B.n483 B.n12 10.6151
R1025 B.n487 B.n12 10.6151
R1026 B.n488 B.n487 10.6151
R1027 B.n489 B.n488 10.6151
R1028 B.n489 B.n10 10.6151
R1029 B.n493 B.n10 10.6151
R1030 B.n494 B.n493 10.6151
R1031 B.n495 B.n494 10.6151
R1032 B.n495 B.n8 10.6151
R1033 B.n499 B.n8 10.6151
R1034 B.n500 B.n499 10.6151
R1035 B.n501 B.n500 10.6151
R1036 B.n501 B.n6 10.6151
R1037 B.n505 B.n6 10.6151
R1038 B.n506 B.n505 10.6151
R1039 B.n507 B.n506 10.6151
R1040 B.n507 B.n4 10.6151
R1041 B.n511 B.n4 10.6151
R1042 B.n512 B.n511 10.6151
R1043 B.n513 B.n512 10.6151
R1044 B.n513 B.n0 10.6151
R1045 B.n470 B.n469 10.6151
R1046 B.n469 B.n18 10.6151
R1047 B.n465 B.n18 10.6151
R1048 B.n465 B.n464 10.6151
R1049 B.n464 B.n463 10.6151
R1050 B.n463 B.n20 10.6151
R1051 B.n459 B.n20 10.6151
R1052 B.n459 B.n458 10.6151
R1053 B.n458 B.n457 10.6151
R1054 B.n457 B.n22 10.6151
R1055 B.n453 B.n22 10.6151
R1056 B.n453 B.n452 10.6151
R1057 B.n452 B.n451 10.6151
R1058 B.n451 B.n24 10.6151
R1059 B.n447 B.n24 10.6151
R1060 B.n447 B.n446 10.6151
R1061 B.n446 B.n445 10.6151
R1062 B.n445 B.n26 10.6151
R1063 B.n441 B.n26 10.6151
R1064 B.n441 B.n440 10.6151
R1065 B.n440 B.n439 10.6151
R1066 B.n439 B.n28 10.6151
R1067 B.n435 B.n28 10.6151
R1068 B.n435 B.n434 10.6151
R1069 B.n434 B.n433 10.6151
R1070 B.n433 B.n30 10.6151
R1071 B.n429 B.n30 10.6151
R1072 B.n427 B.n426 10.6151
R1073 B.n426 B.n34 10.6151
R1074 B.n422 B.n34 10.6151
R1075 B.n422 B.n421 10.6151
R1076 B.n421 B.n420 10.6151
R1077 B.n420 B.n36 10.6151
R1078 B.n416 B.n36 10.6151
R1079 B.n416 B.n415 10.6151
R1080 B.n413 B.n40 10.6151
R1081 B.n409 B.n40 10.6151
R1082 B.n409 B.n408 10.6151
R1083 B.n408 B.n407 10.6151
R1084 B.n407 B.n42 10.6151
R1085 B.n403 B.n42 10.6151
R1086 B.n403 B.n402 10.6151
R1087 B.n402 B.n401 10.6151
R1088 B.n401 B.n44 10.6151
R1089 B.n397 B.n44 10.6151
R1090 B.n397 B.n396 10.6151
R1091 B.n396 B.n395 10.6151
R1092 B.n395 B.n46 10.6151
R1093 B.n391 B.n46 10.6151
R1094 B.n391 B.n390 10.6151
R1095 B.n390 B.n389 10.6151
R1096 B.n389 B.n48 10.6151
R1097 B.n385 B.n48 10.6151
R1098 B.n385 B.n384 10.6151
R1099 B.n384 B.n383 10.6151
R1100 B.n383 B.n50 10.6151
R1101 B.n379 B.n50 10.6151
R1102 B.n379 B.n378 10.6151
R1103 B.n378 B.n377 10.6151
R1104 B.n377 B.n52 10.6151
R1105 B.n373 B.n52 10.6151
R1106 B.n373 B.n372 10.6151
R1107 B.n371 B.n54 10.6151
R1108 B.n367 B.n54 10.6151
R1109 B.n367 B.n366 10.6151
R1110 B.n366 B.n365 10.6151
R1111 B.n365 B.n56 10.6151
R1112 B.n361 B.n56 10.6151
R1113 B.n361 B.n360 10.6151
R1114 B.n360 B.n359 10.6151
R1115 B.n359 B.n58 10.6151
R1116 B.n355 B.n58 10.6151
R1117 B.n355 B.n354 10.6151
R1118 B.n354 B.n353 10.6151
R1119 B.n353 B.n60 10.6151
R1120 B.n349 B.n60 10.6151
R1121 B.n349 B.n348 10.6151
R1122 B.n348 B.n347 10.6151
R1123 B.n347 B.n62 10.6151
R1124 B.n343 B.n62 10.6151
R1125 B.n343 B.n342 10.6151
R1126 B.n342 B.n341 10.6151
R1127 B.n341 B.n64 10.6151
R1128 B.n337 B.n64 10.6151
R1129 B.n337 B.n336 10.6151
R1130 B.n336 B.n335 10.6151
R1131 B.n335 B.n66 10.6151
R1132 B.n331 B.n66 10.6151
R1133 B.n331 B.n330 10.6151
R1134 B.n330 B.n329 10.6151
R1135 B.n329 B.n68 10.6151
R1136 B.n325 B.n68 10.6151
R1137 B.n325 B.n324 10.6151
R1138 B.n324 B.n323 10.6151
R1139 B.n323 B.n70 10.6151
R1140 B.n319 B.n70 10.6151
R1141 B.n319 B.n318 10.6151
R1142 B.n318 B.n317 10.6151
R1143 B.n317 B.n72 10.6151
R1144 B.n313 B.n72 10.6151
R1145 B.n313 B.n312 10.6151
R1146 B.n312 B.n311 10.6151
R1147 B.n311 B.n74 10.6151
R1148 B.n307 B.n74 10.6151
R1149 B.n307 B.n306 10.6151
R1150 B.n306 B.n305 10.6151
R1151 B.n305 B.n76 10.6151
R1152 B.n301 B.n76 10.6151
R1153 B.n301 B.n300 10.6151
R1154 B.n300 B.n299 10.6151
R1155 B.n299 B.n78 10.6151
R1156 B.n295 B.n78 10.6151
R1157 B.n295 B.n294 10.6151
R1158 B.n294 B.n293 10.6151
R1159 B.n293 B.n80 10.6151
R1160 B.n289 B.n80 10.6151
R1161 B.n289 B.n288 10.6151
R1162 B.n288 B.n287 10.6151
R1163 B.n287 B.n82 10.6151
R1164 B.n283 B.n82 10.6151
R1165 B.n283 B.n282 10.6151
R1166 B.n282 B.n281 10.6151
R1167 B.n281 B.n84 10.6151
R1168 B.n134 B.n1 10.6151
R1169 B.n135 B.n134 10.6151
R1170 B.n135 B.n132 10.6151
R1171 B.n139 B.n132 10.6151
R1172 B.n140 B.n139 10.6151
R1173 B.n141 B.n140 10.6151
R1174 B.n141 B.n130 10.6151
R1175 B.n145 B.n130 10.6151
R1176 B.n146 B.n145 10.6151
R1177 B.n147 B.n146 10.6151
R1178 B.n147 B.n128 10.6151
R1179 B.n151 B.n128 10.6151
R1180 B.n152 B.n151 10.6151
R1181 B.n153 B.n152 10.6151
R1182 B.n153 B.n126 10.6151
R1183 B.n157 B.n126 10.6151
R1184 B.n158 B.n157 10.6151
R1185 B.n159 B.n158 10.6151
R1186 B.n159 B.n124 10.6151
R1187 B.n163 B.n124 10.6151
R1188 B.n164 B.n163 10.6151
R1189 B.n165 B.n164 10.6151
R1190 B.n165 B.n122 10.6151
R1191 B.n169 B.n122 10.6151
R1192 B.n170 B.n169 10.6151
R1193 B.n171 B.n170 10.6151
R1194 B.n171 B.n120 10.6151
R1195 B.n175 B.n120 10.6151
R1196 B.n176 B.n175 10.6151
R1197 B.n177 B.n118 10.6151
R1198 B.n181 B.n118 10.6151
R1199 B.n182 B.n181 10.6151
R1200 B.n183 B.n182 10.6151
R1201 B.n183 B.n116 10.6151
R1202 B.n187 B.n116 10.6151
R1203 B.n188 B.n187 10.6151
R1204 B.n189 B.n188 10.6151
R1205 B.n189 B.n114 10.6151
R1206 B.n193 B.n114 10.6151
R1207 B.n194 B.n193 10.6151
R1208 B.n195 B.n194 10.6151
R1209 B.n195 B.n112 10.6151
R1210 B.n199 B.n112 10.6151
R1211 B.n200 B.n199 10.6151
R1212 B.n201 B.n200 10.6151
R1213 B.n201 B.n110 10.6151
R1214 B.n205 B.n110 10.6151
R1215 B.n206 B.n205 10.6151
R1216 B.n207 B.n206 10.6151
R1217 B.n207 B.n108 10.6151
R1218 B.n211 B.n108 10.6151
R1219 B.n212 B.n211 10.6151
R1220 B.n213 B.n212 10.6151
R1221 B.n213 B.n106 10.6151
R1222 B.n217 B.n106 10.6151
R1223 B.n218 B.n217 10.6151
R1224 B.n220 B.n102 10.6151
R1225 B.n224 B.n102 10.6151
R1226 B.n225 B.n224 10.6151
R1227 B.n226 B.n225 10.6151
R1228 B.n226 B.n100 10.6151
R1229 B.n230 B.n100 10.6151
R1230 B.n231 B.n230 10.6151
R1231 B.n235 B.n231 10.6151
R1232 B.n239 B.n98 10.6151
R1233 B.n240 B.n239 10.6151
R1234 B.n241 B.n240 10.6151
R1235 B.n241 B.n96 10.6151
R1236 B.n245 B.n96 10.6151
R1237 B.n246 B.n245 10.6151
R1238 B.n247 B.n246 10.6151
R1239 B.n247 B.n94 10.6151
R1240 B.n251 B.n94 10.6151
R1241 B.n252 B.n251 10.6151
R1242 B.n253 B.n252 10.6151
R1243 B.n253 B.n92 10.6151
R1244 B.n257 B.n92 10.6151
R1245 B.n258 B.n257 10.6151
R1246 B.n259 B.n258 10.6151
R1247 B.n259 B.n90 10.6151
R1248 B.n263 B.n90 10.6151
R1249 B.n264 B.n263 10.6151
R1250 B.n265 B.n264 10.6151
R1251 B.n265 B.n88 10.6151
R1252 B.n269 B.n88 10.6151
R1253 B.n270 B.n269 10.6151
R1254 B.n271 B.n270 10.6151
R1255 B.n271 B.n86 10.6151
R1256 B.n275 B.n86 10.6151
R1257 B.n276 B.n275 10.6151
R1258 B.n277 B.n276 10.6151
R1259 B.n517 B.n0 8.11757
R1260 B.n517 B.n1 8.11757
R1261 B.n428 B.n427 6.5566
R1262 B.n415 B.n414 6.5566
R1263 B.n220 B.n219 6.5566
R1264 B.n235 B.n234 6.5566
R1265 B.n429 B.n428 4.05904
R1266 B.n414 B.n413 4.05904
R1267 B.n219 B.n218 4.05904
R1268 B.n234 B.n98 4.05904
C0 VN w_n2488_n2408# 4.05583f
C1 w_n2488_n2408# VDD2 1.29126f
C2 VN VP 5.01317f
C3 VP VDD2 0.369015f
C4 VN B 0.979789f
C5 VDD2 B 1.10872f
C6 VN VTAIL 3.03845f
C7 VDD2 VTAIL 4.20345f
C8 VN VDD2 2.88702f
C9 w_n2488_n2408# VDD1 1.2441f
C10 VP VDD1 3.10659f
C11 B VDD1 1.06314f
C12 VP w_n2488_n2408# 4.37466f
C13 VTAIL VDD1 4.15192f
C14 w_n2488_n2408# B 7.40992f
C15 VP B 1.50701f
C16 w_n2488_n2408# VTAIL 2.87717f
C17 VN VDD1 0.148801f
C18 VDD2 VDD1 0.931855f
C19 VP VTAIL 3.05256f
C20 VTAIL B 3.22225f
C21 VDD2 VSUBS 0.761833f
C22 VDD1 VSUBS 4.87066f
C23 VTAIL VSUBS 0.722561f
C24 VN VSUBS 5.08206f
C25 VP VSUBS 1.793447f
C26 B VSUBS 3.521306f
C27 w_n2488_n2408# VSUBS 74.4907f
C28 B.n0 VSUBS 0.007039f
C29 B.n1 VSUBS 0.007039f
C30 B.n2 VSUBS 0.01041f
C31 B.n3 VSUBS 0.007977f
C32 B.n4 VSUBS 0.007977f
C33 B.n5 VSUBS 0.007977f
C34 B.n6 VSUBS 0.007977f
C35 B.n7 VSUBS 0.007977f
C36 B.n8 VSUBS 0.007977f
C37 B.n9 VSUBS 0.007977f
C38 B.n10 VSUBS 0.007977f
C39 B.n11 VSUBS 0.007977f
C40 B.n12 VSUBS 0.007977f
C41 B.n13 VSUBS 0.007977f
C42 B.n14 VSUBS 0.007977f
C43 B.n15 VSUBS 0.007977f
C44 B.n16 VSUBS 0.007977f
C45 B.n17 VSUBS 0.018103f
C46 B.n18 VSUBS 0.007977f
C47 B.n19 VSUBS 0.007977f
C48 B.n20 VSUBS 0.007977f
C49 B.n21 VSUBS 0.007977f
C50 B.n22 VSUBS 0.007977f
C51 B.n23 VSUBS 0.007977f
C52 B.n24 VSUBS 0.007977f
C53 B.n25 VSUBS 0.007977f
C54 B.n26 VSUBS 0.007977f
C55 B.n27 VSUBS 0.007977f
C56 B.n28 VSUBS 0.007977f
C57 B.n29 VSUBS 0.007977f
C58 B.n30 VSUBS 0.007977f
C59 B.n31 VSUBS 0.007977f
C60 B.t10 VSUBS 0.126507f
C61 B.t11 VSUBS 0.154057f
C62 B.t9 VSUBS 0.838229f
C63 B.n32 VSUBS 0.260717f
C64 B.n33 VSUBS 0.201308f
C65 B.n34 VSUBS 0.007977f
C66 B.n35 VSUBS 0.007977f
C67 B.n36 VSUBS 0.007977f
C68 B.n37 VSUBS 0.007977f
C69 B.t7 VSUBS 0.126509f
C70 B.t8 VSUBS 0.15406f
C71 B.t6 VSUBS 0.838229f
C72 B.n38 VSUBS 0.260715f
C73 B.n39 VSUBS 0.201305f
C74 B.n40 VSUBS 0.007977f
C75 B.n41 VSUBS 0.007977f
C76 B.n42 VSUBS 0.007977f
C77 B.n43 VSUBS 0.007977f
C78 B.n44 VSUBS 0.007977f
C79 B.n45 VSUBS 0.007977f
C80 B.n46 VSUBS 0.007977f
C81 B.n47 VSUBS 0.007977f
C82 B.n48 VSUBS 0.007977f
C83 B.n49 VSUBS 0.007977f
C84 B.n50 VSUBS 0.007977f
C85 B.n51 VSUBS 0.007977f
C86 B.n52 VSUBS 0.007977f
C87 B.n53 VSUBS 0.018103f
C88 B.n54 VSUBS 0.007977f
C89 B.n55 VSUBS 0.007977f
C90 B.n56 VSUBS 0.007977f
C91 B.n57 VSUBS 0.007977f
C92 B.n58 VSUBS 0.007977f
C93 B.n59 VSUBS 0.007977f
C94 B.n60 VSUBS 0.007977f
C95 B.n61 VSUBS 0.007977f
C96 B.n62 VSUBS 0.007977f
C97 B.n63 VSUBS 0.007977f
C98 B.n64 VSUBS 0.007977f
C99 B.n65 VSUBS 0.007977f
C100 B.n66 VSUBS 0.007977f
C101 B.n67 VSUBS 0.007977f
C102 B.n68 VSUBS 0.007977f
C103 B.n69 VSUBS 0.007977f
C104 B.n70 VSUBS 0.007977f
C105 B.n71 VSUBS 0.007977f
C106 B.n72 VSUBS 0.007977f
C107 B.n73 VSUBS 0.007977f
C108 B.n74 VSUBS 0.007977f
C109 B.n75 VSUBS 0.007977f
C110 B.n76 VSUBS 0.007977f
C111 B.n77 VSUBS 0.007977f
C112 B.n78 VSUBS 0.007977f
C113 B.n79 VSUBS 0.007977f
C114 B.n80 VSUBS 0.007977f
C115 B.n81 VSUBS 0.007977f
C116 B.n82 VSUBS 0.007977f
C117 B.n83 VSUBS 0.007977f
C118 B.n84 VSUBS 0.017899f
C119 B.n85 VSUBS 0.007977f
C120 B.n86 VSUBS 0.007977f
C121 B.n87 VSUBS 0.007977f
C122 B.n88 VSUBS 0.007977f
C123 B.n89 VSUBS 0.007977f
C124 B.n90 VSUBS 0.007977f
C125 B.n91 VSUBS 0.007977f
C126 B.n92 VSUBS 0.007977f
C127 B.n93 VSUBS 0.007977f
C128 B.n94 VSUBS 0.007977f
C129 B.n95 VSUBS 0.007977f
C130 B.n96 VSUBS 0.007977f
C131 B.n97 VSUBS 0.007977f
C132 B.n98 VSUBS 0.005514f
C133 B.n99 VSUBS 0.007977f
C134 B.n100 VSUBS 0.007977f
C135 B.n101 VSUBS 0.007977f
C136 B.n102 VSUBS 0.007977f
C137 B.n103 VSUBS 0.007977f
C138 B.t2 VSUBS 0.126507f
C139 B.t1 VSUBS 0.154057f
C140 B.t0 VSUBS 0.838229f
C141 B.n104 VSUBS 0.260717f
C142 B.n105 VSUBS 0.201308f
C143 B.n106 VSUBS 0.007977f
C144 B.n107 VSUBS 0.007977f
C145 B.n108 VSUBS 0.007977f
C146 B.n109 VSUBS 0.007977f
C147 B.n110 VSUBS 0.007977f
C148 B.n111 VSUBS 0.007977f
C149 B.n112 VSUBS 0.007977f
C150 B.n113 VSUBS 0.007977f
C151 B.n114 VSUBS 0.007977f
C152 B.n115 VSUBS 0.007977f
C153 B.n116 VSUBS 0.007977f
C154 B.n117 VSUBS 0.007977f
C155 B.n118 VSUBS 0.007977f
C156 B.n119 VSUBS 0.016856f
C157 B.n120 VSUBS 0.007977f
C158 B.n121 VSUBS 0.007977f
C159 B.n122 VSUBS 0.007977f
C160 B.n123 VSUBS 0.007977f
C161 B.n124 VSUBS 0.007977f
C162 B.n125 VSUBS 0.007977f
C163 B.n126 VSUBS 0.007977f
C164 B.n127 VSUBS 0.007977f
C165 B.n128 VSUBS 0.007977f
C166 B.n129 VSUBS 0.007977f
C167 B.n130 VSUBS 0.007977f
C168 B.n131 VSUBS 0.007977f
C169 B.n132 VSUBS 0.007977f
C170 B.n133 VSUBS 0.007977f
C171 B.n134 VSUBS 0.007977f
C172 B.n135 VSUBS 0.007977f
C173 B.n136 VSUBS 0.007977f
C174 B.n137 VSUBS 0.007977f
C175 B.n138 VSUBS 0.007977f
C176 B.n139 VSUBS 0.007977f
C177 B.n140 VSUBS 0.007977f
C178 B.n141 VSUBS 0.007977f
C179 B.n142 VSUBS 0.007977f
C180 B.n143 VSUBS 0.007977f
C181 B.n144 VSUBS 0.007977f
C182 B.n145 VSUBS 0.007977f
C183 B.n146 VSUBS 0.007977f
C184 B.n147 VSUBS 0.007977f
C185 B.n148 VSUBS 0.007977f
C186 B.n149 VSUBS 0.007977f
C187 B.n150 VSUBS 0.007977f
C188 B.n151 VSUBS 0.007977f
C189 B.n152 VSUBS 0.007977f
C190 B.n153 VSUBS 0.007977f
C191 B.n154 VSUBS 0.007977f
C192 B.n155 VSUBS 0.007977f
C193 B.n156 VSUBS 0.007977f
C194 B.n157 VSUBS 0.007977f
C195 B.n158 VSUBS 0.007977f
C196 B.n159 VSUBS 0.007977f
C197 B.n160 VSUBS 0.007977f
C198 B.n161 VSUBS 0.007977f
C199 B.n162 VSUBS 0.007977f
C200 B.n163 VSUBS 0.007977f
C201 B.n164 VSUBS 0.007977f
C202 B.n165 VSUBS 0.007977f
C203 B.n166 VSUBS 0.007977f
C204 B.n167 VSUBS 0.007977f
C205 B.n168 VSUBS 0.007977f
C206 B.n169 VSUBS 0.007977f
C207 B.n170 VSUBS 0.007977f
C208 B.n171 VSUBS 0.007977f
C209 B.n172 VSUBS 0.007977f
C210 B.n173 VSUBS 0.007977f
C211 B.n174 VSUBS 0.007977f
C212 B.n175 VSUBS 0.007977f
C213 B.n176 VSUBS 0.016856f
C214 B.n177 VSUBS 0.018103f
C215 B.n178 VSUBS 0.018103f
C216 B.n179 VSUBS 0.007977f
C217 B.n180 VSUBS 0.007977f
C218 B.n181 VSUBS 0.007977f
C219 B.n182 VSUBS 0.007977f
C220 B.n183 VSUBS 0.007977f
C221 B.n184 VSUBS 0.007977f
C222 B.n185 VSUBS 0.007977f
C223 B.n186 VSUBS 0.007977f
C224 B.n187 VSUBS 0.007977f
C225 B.n188 VSUBS 0.007977f
C226 B.n189 VSUBS 0.007977f
C227 B.n190 VSUBS 0.007977f
C228 B.n191 VSUBS 0.007977f
C229 B.n192 VSUBS 0.007977f
C230 B.n193 VSUBS 0.007977f
C231 B.n194 VSUBS 0.007977f
C232 B.n195 VSUBS 0.007977f
C233 B.n196 VSUBS 0.007977f
C234 B.n197 VSUBS 0.007977f
C235 B.n198 VSUBS 0.007977f
C236 B.n199 VSUBS 0.007977f
C237 B.n200 VSUBS 0.007977f
C238 B.n201 VSUBS 0.007977f
C239 B.n202 VSUBS 0.007977f
C240 B.n203 VSUBS 0.007977f
C241 B.n204 VSUBS 0.007977f
C242 B.n205 VSUBS 0.007977f
C243 B.n206 VSUBS 0.007977f
C244 B.n207 VSUBS 0.007977f
C245 B.n208 VSUBS 0.007977f
C246 B.n209 VSUBS 0.007977f
C247 B.n210 VSUBS 0.007977f
C248 B.n211 VSUBS 0.007977f
C249 B.n212 VSUBS 0.007977f
C250 B.n213 VSUBS 0.007977f
C251 B.n214 VSUBS 0.007977f
C252 B.n215 VSUBS 0.007977f
C253 B.n216 VSUBS 0.007977f
C254 B.n217 VSUBS 0.007977f
C255 B.n218 VSUBS 0.005514f
C256 B.n219 VSUBS 0.018482f
C257 B.n220 VSUBS 0.006452f
C258 B.n221 VSUBS 0.007977f
C259 B.n222 VSUBS 0.007977f
C260 B.n223 VSUBS 0.007977f
C261 B.n224 VSUBS 0.007977f
C262 B.n225 VSUBS 0.007977f
C263 B.n226 VSUBS 0.007977f
C264 B.n227 VSUBS 0.007977f
C265 B.n228 VSUBS 0.007977f
C266 B.n229 VSUBS 0.007977f
C267 B.n230 VSUBS 0.007977f
C268 B.n231 VSUBS 0.007977f
C269 B.t5 VSUBS 0.126509f
C270 B.t4 VSUBS 0.15406f
C271 B.t3 VSUBS 0.838229f
C272 B.n232 VSUBS 0.260715f
C273 B.n233 VSUBS 0.201305f
C274 B.n234 VSUBS 0.018482f
C275 B.n235 VSUBS 0.006452f
C276 B.n236 VSUBS 0.007977f
C277 B.n237 VSUBS 0.007977f
C278 B.n238 VSUBS 0.007977f
C279 B.n239 VSUBS 0.007977f
C280 B.n240 VSUBS 0.007977f
C281 B.n241 VSUBS 0.007977f
C282 B.n242 VSUBS 0.007977f
C283 B.n243 VSUBS 0.007977f
C284 B.n244 VSUBS 0.007977f
C285 B.n245 VSUBS 0.007977f
C286 B.n246 VSUBS 0.007977f
C287 B.n247 VSUBS 0.007977f
C288 B.n248 VSUBS 0.007977f
C289 B.n249 VSUBS 0.007977f
C290 B.n250 VSUBS 0.007977f
C291 B.n251 VSUBS 0.007977f
C292 B.n252 VSUBS 0.007977f
C293 B.n253 VSUBS 0.007977f
C294 B.n254 VSUBS 0.007977f
C295 B.n255 VSUBS 0.007977f
C296 B.n256 VSUBS 0.007977f
C297 B.n257 VSUBS 0.007977f
C298 B.n258 VSUBS 0.007977f
C299 B.n259 VSUBS 0.007977f
C300 B.n260 VSUBS 0.007977f
C301 B.n261 VSUBS 0.007977f
C302 B.n262 VSUBS 0.007977f
C303 B.n263 VSUBS 0.007977f
C304 B.n264 VSUBS 0.007977f
C305 B.n265 VSUBS 0.007977f
C306 B.n266 VSUBS 0.007977f
C307 B.n267 VSUBS 0.007977f
C308 B.n268 VSUBS 0.007977f
C309 B.n269 VSUBS 0.007977f
C310 B.n270 VSUBS 0.007977f
C311 B.n271 VSUBS 0.007977f
C312 B.n272 VSUBS 0.007977f
C313 B.n273 VSUBS 0.007977f
C314 B.n274 VSUBS 0.007977f
C315 B.n275 VSUBS 0.007977f
C316 B.n276 VSUBS 0.007977f
C317 B.n277 VSUBS 0.017059f
C318 B.n278 VSUBS 0.018103f
C319 B.n279 VSUBS 0.016856f
C320 B.n280 VSUBS 0.007977f
C321 B.n281 VSUBS 0.007977f
C322 B.n282 VSUBS 0.007977f
C323 B.n283 VSUBS 0.007977f
C324 B.n284 VSUBS 0.007977f
C325 B.n285 VSUBS 0.007977f
C326 B.n286 VSUBS 0.007977f
C327 B.n287 VSUBS 0.007977f
C328 B.n288 VSUBS 0.007977f
C329 B.n289 VSUBS 0.007977f
C330 B.n290 VSUBS 0.007977f
C331 B.n291 VSUBS 0.007977f
C332 B.n292 VSUBS 0.007977f
C333 B.n293 VSUBS 0.007977f
C334 B.n294 VSUBS 0.007977f
C335 B.n295 VSUBS 0.007977f
C336 B.n296 VSUBS 0.007977f
C337 B.n297 VSUBS 0.007977f
C338 B.n298 VSUBS 0.007977f
C339 B.n299 VSUBS 0.007977f
C340 B.n300 VSUBS 0.007977f
C341 B.n301 VSUBS 0.007977f
C342 B.n302 VSUBS 0.007977f
C343 B.n303 VSUBS 0.007977f
C344 B.n304 VSUBS 0.007977f
C345 B.n305 VSUBS 0.007977f
C346 B.n306 VSUBS 0.007977f
C347 B.n307 VSUBS 0.007977f
C348 B.n308 VSUBS 0.007977f
C349 B.n309 VSUBS 0.007977f
C350 B.n310 VSUBS 0.007977f
C351 B.n311 VSUBS 0.007977f
C352 B.n312 VSUBS 0.007977f
C353 B.n313 VSUBS 0.007977f
C354 B.n314 VSUBS 0.007977f
C355 B.n315 VSUBS 0.007977f
C356 B.n316 VSUBS 0.007977f
C357 B.n317 VSUBS 0.007977f
C358 B.n318 VSUBS 0.007977f
C359 B.n319 VSUBS 0.007977f
C360 B.n320 VSUBS 0.007977f
C361 B.n321 VSUBS 0.007977f
C362 B.n322 VSUBS 0.007977f
C363 B.n323 VSUBS 0.007977f
C364 B.n324 VSUBS 0.007977f
C365 B.n325 VSUBS 0.007977f
C366 B.n326 VSUBS 0.007977f
C367 B.n327 VSUBS 0.007977f
C368 B.n328 VSUBS 0.007977f
C369 B.n329 VSUBS 0.007977f
C370 B.n330 VSUBS 0.007977f
C371 B.n331 VSUBS 0.007977f
C372 B.n332 VSUBS 0.007977f
C373 B.n333 VSUBS 0.007977f
C374 B.n334 VSUBS 0.007977f
C375 B.n335 VSUBS 0.007977f
C376 B.n336 VSUBS 0.007977f
C377 B.n337 VSUBS 0.007977f
C378 B.n338 VSUBS 0.007977f
C379 B.n339 VSUBS 0.007977f
C380 B.n340 VSUBS 0.007977f
C381 B.n341 VSUBS 0.007977f
C382 B.n342 VSUBS 0.007977f
C383 B.n343 VSUBS 0.007977f
C384 B.n344 VSUBS 0.007977f
C385 B.n345 VSUBS 0.007977f
C386 B.n346 VSUBS 0.007977f
C387 B.n347 VSUBS 0.007977f
C388 B.n348 VSUBS 0.007977f
C389 B.n349 VSUBS 0.007977f
C390 B.n350 VSUBS 0.007977f
C391 B.n351 VSUBS 0.007977f
C392 B.n352 VSUBS 0.007977f
C393 B.n353 VSUBS 0.007977f
C394 B.n354 VSUBS 0.007977f
C395 B.n355 VSUBS 0.007977f
C396 B.n356 VSUBS 0.007977f
C397 B.n357 VSUBS 0.007977f
C398 B.n358 VSUBS 0.007977f
C399 B.n359 VSUBS 0.007977f
C400 B.n360 VSUBS 0.007977f
C401 B.n361 VSUBS 0.007977f
C402 B.n362 VSUBS 0.007977f
C403 B.n363 VSUBS 0.007977f
C404 B.n364 VSUBS 0.007977f
C405 B.n365 VSUBS 0.007977f
C406 B.n366 VSUBS 0.007977f
C407 B.n367 VSUBS 0.007977f
C408 B.n368 VSUBS 0.007977f
C409 B.n369 VSUBS 0.007977f
C410 B.n370 VSUBS 0.016856f
C411 B.n371 VSUBS 0.016856f
C412 B.n372 VSUBS 0.018103f
C413 B.n373 VSUBS 0.007977f
C414 B.n374 VSUBS 0.007977f
C415 B.n375 VSUBS 0.007977f
C416 B.n376 VSUBS 0.007977f
C417 B.n377 VSUBS 0.007977f
C418 B.n378 VSUBS 0.007977f
C419 B.n379 VSUBS 0.007977f
C420 B.n380 VSUBS 0.007977f
C421 B.n381 VSUBS 0.007977f
C422 B.n382 VSUBS 0.007977f
C423 B.n383 VSUBS 0.007977f
C424 B.n384 VSUBS 0.007977f
C425 B.n385 VSUBS 0.007977f
C426 B.n386 VSUBS 0.007977f
C427 B.n387 VSUBS 0.007977f
C428 B.n388 VSUBS 0.007977f
C429 B.n389 VSUBS 0.007977f
C430 B.n390 VSUBS 0.007977f
C431 B.n391 VSUBS 0.007977f
C432 B.n392 VSUBS 0.007977f
C433 B.n393 VSUBS 0.007977f
C434 B.n394 VSUBS 0.007977f
C435 B.n395 VSUBS 0.007977f
C436 B.n396 VSUBS 0.007977f
C437 B.n397 VSUBS 0.007977f
C438 B.n398 VSUBS 0.007977f
C439 B.n399 VSUBS 0.007977f
C440 B.n400 VSUBS 0.007977f
C441 B.n401 VSUBS 0.007977f
C442 B.n402 VSUBS 0.007977f
C443 B.n403 VSUBS 0.007977f
C444 B.n404 VSUBS 0.007977f
C445 B.n405 VSUBS 0.007977f
C446 B.n406 VSUBS 0.007977f
C447 B.n407 VSUBS 0.007977f
C448 B.n408 VSUBS 0.007977f
C449 B.n409 VSUBS 0.007977f
C450 B.n410 VSUBS 0.007977f
C451 B.n411 VSUBS 0.007977f
C452 B.n412 VSUBS 0.007977f
C453 B.n413 VSUBS 0.005514f
C454 B.n414 VSUBS 0.018482f
C455 B.n415 VSUBS 0.006452f
C456 B.n416 VSUBS 0.007977f
C457 B.n417 VSUBS 0.007977f
C458 B.n418 VSUBS 0.007977f
C459 B.n419 VSUBS 0.007977f
C460 B.n420 VSUBS 0.007977f
C461 B.n421 VSUBS 0.007977f
C462 B.n422 VSUBS 0.007977f
C463 B.n423 VSUBS 0.007977f
C464 B.n424 VSUBS 0.007977f
C465 B.n425 VSUBS 0.007977f
C466 B.n426 VSUBS 0.007977f
C467 B.n427 VSUBS 0.006452f
C468 B.n428 VSUBS 0.018482f
C469 B.n429 VSUBS 0.005514f
C470 B.n430 VSUBS 0.007977f
C471 B.n431 VSUBS 0.007977f
C472 B.n432 VSUBS 0.007977f
C473 B.n433 VSUBS 0.007977f
C474 B.n434 VSUBS 0.007977f
C475 B.n435 VSUBS 0.007977f
C476 B.n436 VSUBS 0.007977f
C477 B.n437 VSUBS 0.007977f
C478 B.n438 VSUBS 0.007977f
C479 B.n439 VSUBS 0.007977f
C480 B.n440 VSUBS 0.007977f
C481 B.n441 VSUBS 0.007977f
C482 B.n442 VSUBS 0.007977f
C483 B.n443 VSUBS 0.007977f
C484 B.n444 VSUBS 0.007977f
C485 B.n445 VSUBS 0.007977f
C486 B.n446 VSUBS 0.007977f
C487 B.n447 VSUBS 0.007977f
C488 B.n448 VSUBS 0.007977f
C489 B.n449 VSUBS 0.007977f
C490 B.n450 VSUBS 0.007977f
C491 B.n451 VSUBS 0.007977f
C492 B.n452 VSUBS 0.007977f
C493 B.n453 VSUBS 0.007977f
C494 B.n454 VSUBS 0.007977f
C495 B.n455 VSUBS 0.007977f
C496 B.n456 VSUBS 0.007977f
C497 B.n457 VSUBS 0.007977f
C498 B.n458 VSUBS 0.007977f
C499 B.n459 VSUBS 0.007977f
C500 B.n460 VSUBS 0.007977f
C501 B.n461 VSUBS 0.007977f
C502 B.n462 VSUBS 0.007977f
C503 B.n463 VSUBS 0.007977f
C504 B.n464 VSUBS 0.007977f
C505 B.n465 VSUBS 0.007977f
C506 B.n466 VSUBS 0.007977f
C507 B.n467 VSUBS 0.007977f
C508 B.n468 VSUBS 0.007977f
C509 B.n469 VSUBS 0.007977f
C510 B.n470 VSUBS 0.018103f
C511 B.n471 VSUBS 0.016856f
C512 B.n472 VSUBS 0.016856f
C513 B.n473 VSUBS 0.007977f
C514 B.n474 VSUBS 0.007977f
C515 B.n475 VSUBS 0.007977f
C516 B.n476 VSUBS 0.007977f
C517 B.n477 VSUBS 0.007977f
C518 B.n478 VSUBS 0.007977f
C519 B.n479 VSUBS 0.007977f
C520 B.n480 VSUBS 0.007977f
C521 B.n481 VSUBS 0.007977f
C522 B.n482 VSUBS 0.007977f
C523 B.n483 VSUBS 0.007977f
C524 B.n484 VSUBS 0.007977f
C525 B.n485 VSUBS 0.007977f
C526 B.n486 VSUBS 0.007977f
C527 B.n487 VSUBS 0.007977f
C528 B.n488 VSUBS 0.007977f
C529 B.n489 VSUBS 0.007977f
C530 B.n490 VSUBS 0.007977f
C531 B.n491 VSUBS 0.007977f
C532 B.n492 VSUBS 0.007977f
C533 B.n493 VSUBS 0.007977f
C534 B.n494 VSUBS 0.007977f
C535 B.n495 VSUBS 0.007977f
C536 B.n496 VSUBS 0.007977f
C537 B.n497 VSUBS 0.007977f
C538 B.n498 VSUBS 0.007977f
C539 B.n499 VSUBS 0.007977f
C540 B.n500 VSUBS 0.007977f
C541 B.n501 VSUBS 0.007977f
C542 B.n502 VSUBS 0.007977f
C543 B.n503 VSUBS 0.007977f
C544 B.n504 VSUBS 0.007977f
C545 B.n505 VSUBS 0.007977f
C546 B.n506 VSUBS 0.007977f
C547 B.n507 VSUBS 0.007977f
C548 B.n508 VSUBS 0.007977f
C549 B.n509 VSUBS 0.007977f
C550 B.n510 VSUBS 0.007977f
C551 B.n511 VSUBS 0.007977f
C552 B.n512 VSUBS 0.007977f
C553 B.n513 VSUBS 0.007977f
C554 B.n514 VSUBS 0.007977f
C555 B.n515 VSUBS 0.01041f
C556 B.n516 VSUBS 0.011089f
C557 B.n517 VSUBS 0.022052f
C558 VDD1.t3 VSUBS 0.156963f
C559 VDD1.t1 VSUBS 0.156963f
C560 VDD1.n0 VSUBS 1.11072f
C561 VDD1.t0 VSUBS 0.156963f
C562 VDD1.t2 VSUBS 0.156963f
C563 VDD1.n1 VSUBS 1.60171f
C564 VP.n0 VSUBS 0.057212f
C565 VP.t1 VSUBS 1.83727f
C566 VP.n1 VSUBS 0.035051f
C567 VP.n2 VSUBS 0.057212f
C568 VP.t3 VSUBS 1.83727f
C569 VP.t2 VSUBS 2.12075f
C570 VP.t0 VSUBS 2.12587f
C571 VP.n3 VSUBS 3.27745f
C572 VP.n4 VSUBS 2.09747f
C573 VP.n5 VSUBS 0.809855f
C574 VP.n6 VSUBS 0.061804f
C575 VP.n7 VSUBS 0.085798f
C576 VP.n8 VSUBS 0.043397f
C577 VP.n9 VSUBS 0.043397f
C578 VP.n10 VSUBS 0.043397f
C579 VP.n11 VSUBS 0.085798f
C580 VP.n12 VSUBS 0.061804f
C581 VP.n13 VSUBS 0.809855f
C582 VP.n14 VSUBS 0.062327f
C583 VTAIL.n0 VSUBS 0.027609f
C584 VTAIL.n1 VSUBS 0.026028f
C585 VTAIL.n2 VSUBS 0.013986f
C586 VTAIL.n3 VSUBS 0.033059f
C587 VTAIL.n4 VSUBS 0.014809f
C588 VTAIL.n5 VSUBS 0.026028f
C589 VTAIL.n6 VSUBS 0.013986f
C590 VTAIL.n7 VSUBS 0.033059f
C591 VTAIL.n8 VSUBS 0.014809f
C592 VTAIL.n9 VSUBS 0.7311f
C593 VTAIL.n10 VSUBS 0.013986f
C594 VTAIL.t6 VSUBS 0.070997f
C595 VTAIL.n11 VSUBS 0.148646f
C596 VTAIL.n12 VSUBS 0.024867f
C597 VTAIL.n13 VSUBS 0.024794f
C598 VTAIL.n14 VSUBS 0.033059f
C599 VTAIL.n15 VSUBS 0.014809f
C600 VTAIL.n16 VSUBS 0.013986f
C601 VTAIL.n17 VSUBS 0.026028f
C602 VTAIL.n18 VSUBS 0.026028f
C603 VTAIL.n19 VSUBS 0.013986f
C604 VTAIL.n20 VSUBS 0.014809f
C605 VTAIL.n21 VSUBS 0.033059f
C606 VTAIL.n22 VSUBS 0.033059f
C607 VTAIL.n23 VSUBS 0.014809f
C608 VTAIL.n24 VSUBS 0.013986f
C609 VTAIL.n25 VSUBS 0.026028f
C610 VTAIL.n26 VSUBS 0.026028f
C611 VTAIL.n27 VSUBS 0.013986f
C612 VTAIL.n28 VSUBS 0.014809f
C613 VTAIL.n29 VSUBS 0.033059f
C614 VTAIL.n30 VSUBS 0.081332f
C615 VTAIL.n31 VSUBS 0.014809f
C616 VTAIL.n32 VSUBS 0.027466f
C617 VTAIL.n33 VSUBS 0.06443f
C618 VTAIL.n34 VSUBS 0.061878f
C619 VTAIL.n35 VSUBS 0.160387f
C620 VTAIL.n36 VSUBS 0.027609f
C621 VTAIL.n37 VSUBS 0.026028f
C622 VTAIL.n38 VSUBS 0.013986f
C623 VTAIL.n39 VSUBS 0.033059f
C624 VTAIL.n40 VSUBS 0.014809f
C625 VTAIL.n41 VSUBS 0.026028f
C626 VTAIL.n42 VSUBS 0.013986f
C627 VTAIL.n43 VSUBS 0.033059f
C628 VTAIL.n44 VSUBS 0.014809f
C629 VTAIL.n45 VSUBS 0.7311f
C630 VTAIL.n46 VSUBS 0.013986f
C631 VTAIL.t3 VSUBS 0.070997f
C632 VTAIL.n47 VSUBS 0.148646f
C633 VTAIL.n48 VSUBS 0.024867f
C634 VTAIL.n49 VSUBS 0.024794f
C635 VTAIL.n50 VSUBS 0.033059f
C636 VTAIL.n51 VSUBS 0.014809f
C637 VTAIL.n52 VSUBS 0.013986f
C638 VTAIL.n53 VSUBS 0.026028f
C639 VTAIL.n54 VSUBS 0.026028f
C640 VTAIL.n55 VSUBS 0.013986f
C641 VTAIL.n56 VSUBS 0.014809f
C642 VTAIL.n57 VSUBS 0.033059f
C643 VTAIL.n58 VSUBS 0.033059f
C644 VTAIL.n59 VSUBS 0.014809f
C645 VTAIL.n60 VSUBS 0.013986f
C646 VTAIL.n61 VSUBS 0.026028f
C647 VTAIL.n62 VSUBS 0.026028f
C648 VTAIL.n63 VSUBS 0.013986f
C649 VTAIL.n64 VSUBS 0.014809f
C650 VTAIL.n65 VSUBS 0.033059f
C651 VTAIL.n66 VSUBS 0.081332f
C652 VTAIL.n67 VSUBS 0.014809f
C653 VTAIL.n68 VSUBS 0.027466f
C654 VTAIL.n69 VSUBS 0.06443f
C655 VTAIL.n70 VSUBS 0.061878f
C656 VTAIL.n71 VSUBS 0.246967f
C657 VTAIL.n72 VSUBS 0.027609f
C658 VTAIL.n73 VSUBS 0.026028f
C659 VTAIL.n74 VSUBS 0.013986f
C660 VTAIL.n75 VSUBS 0.033059f
C661 VTAIL.n76 VSUBS 0.014809f
C662 VTAIL.n77 VSUBS 0.026028f
C663 VTAIL.n78 VSUBS 0.013986f
C664 VTAIL.n79 VSUBS 0.033059f
C665 VTAIL.n80 VSUBS 0.014809f
C666 VTAIL.n81 VSUBS 0.7311f
C667 VTAIL.n82 VSUBS 0.013986f
C668 VTAIL.t2 VSUBS 0.070997f
C669 VTAIL.n83 VSUBS 0.148646f
C670 VTAIL.n84 VSUBS 0.024867f
C671 VTAIL.n85 VSUBS 0.024794f
C672 VTAIL.n86 VSUBS 0.033059f
C673 VTAIL.n87 VSUBS 0.014809f
C674 VTAIL.n88 VSUBS 0.013986f
C675 VTAIL.n89 VSUBS 0.026028f
C676 VTAIL.n90 VSUBS 0.026028f
C677 VTAIL.n91 VSUBS 0.013986f
C678 VTAIL.n92 VSUBS 0.014809f
C679 VTAIL.n93 VSUBS 0.033059f
C680 VTAIL.n94 VSUBS 0.033059f
C681 VTAIL.n95 VSUBS 0.014809f
C682 VTAIL.n96 VSUBS 0.013986f
C683 VTAIL.n97 VSUBS 0.026028f
C684 VTAIL.n98 VSUBS 0.026028f
C685 VTAIL.n99 VSUBS 0.013986f
C686 VTAIL.n100 VSUBS 0.014809f
C687 VTAIL.n101 VSUBS 0.033059f
C688 VTAIL.n102 VSUBS 0.081332f
C689 VTAIL.n103 VSUBS 0.014809f
C690 VTAIL.n104 VSUBS 0.027466f
C691 VTAIL.n105 VSUBS 0.06443f
C692 VTAIL.n106 VSUBS 0.061878f
C693 VTAIL.n107 VSUBS 1.26461f
C694 VTAIL.n108 VSUBS 0.027609f
C695 VTAIL.n109 VSUBS 0.026028f
C696 VTAIL.n110 VSUBS 0.013986f
C697 VTAIL.n111 VSUBS 0.033059f
C698 VTAIL.n112 VSUBS 0.014809f
C699 VTAIL.n113 VSUBS 0.026028f
C700 VTAIL.n114 VSUBS 0.013986f
C701 VTAIL.n115 VSUBS 0.033059f
C702 VTAIL.n116 VSUBS 0.014809f
C703 VTAIL.n117 VSUBS 0.7311f
C704 VTAIL.n118 VSUBS 0.013986f
C705 VTAIL.t7 VSUBS 0.070997f
C706 VTAIL.n119 VSUBS 0.148646f
C707 VTAIL.n120 VSUBS 0.024867f
C708 VTAIL.n121 VSUBS 0.024794f
C709 VTAIL.n122 VSUBS 0.033059f
C710 VTAIL.n123 VSUBS 0.014809f
C711 VTAIL.n124 VSUBS 0.013986f
C712 VTAIL.n125 VSUBS 0.026028f
C713 VTAIL.n126 VSUBS 0.026028f
C714 VTAIL.n127 VSUBS 0.013986f
C715 VTAIL.n128 VSUBS 0.014809f
C716 VTAIL.n129 VSUBS 0.033059f
C717 VTAIL.n130 VSUBS 0.033059f
C718 VTAIL.n131 VSUBS 0.014809f
C719 VTAIL.n132 VSUBS 0.013986f
C720 VTAIL.n133 VSUBS 0.026028f
C721 VTAIL.n134 VSUBS 0.026028f
C722 VTAIL.n135 VSUBS 0.013986f
C723 VTAIL.n136 VSUBS 0.014809f
C724 VTAIL.n137 VSUBS 0.033059f
C725 VTAIL.n138 VSUBS 0.081332f
C726 VTAIL.n139 VSUBS 0.014809f
C727 VTAIL.n140 VSUBS 0.027466f
C728 VTAIL.n141 VSUBS 0.06443f
C729 VTAIL.n142 VSUBS 0.061878f
C730 VTAIL.n143 VSUBS 1.26461f
C731 VTAIL.n144 VSUBS 0.027609f
C732 VTAIL.n145 VSUBS 0.026028f
C733 VTAIL.n146 VSUBS 0.013986f
C734 VTAIL.n147 VSUBS 0.033059f
C735 VTAIL.n148 VSUBS 0.014809f
C736 VTAIL.n149 VSUBS 0.026028f
C737 VTAIL.n150 VSUBS 0.013986f
C738 VTAIL.n151 VSUBS 0.033059f
C739 VTAIL.n152 VSUBS 0.014809f
C740 VTAIL.n153 VSUBS 0.7311f
C741 VTAIL.n154 VSUBS 0.013986f
C742 VTAIL.t5 VSUBS 0.070997f
C743 VTAIL.n155 VSUBS 0.148646f
C744 VTAIL.n156 VSUBS 0.024867f
C745 VTAIL.n157 VSUBS 0.024794f
C746 VTAIL.n158 VSUBS 0.033059f
C747 VTAIL.n159 VSUBS 0.014809f
C748 VTAIL.n160 VSUBS 0.013986f
C749 VTAIL.n161 VSUBS 0.026028f
C750 VTAIL.n162 VSUBS 0.026028f
C751 VTAIL.n163 VSUBS 0.013986f
C752 VTAIL.n164 VSUBS 0.014809f
C753 VTAIL.n165 VSUBS 0.033059f
C754 VTAIL.n166 VSUBS 0.033059f
C755 VTAIL.n167 VSUBS 0.014809f
C756 VTAIL.n168 VSUBS 0.013986f
C757 VTAIL.n169 VSUBS 0.026028f
C758 VTAIL.n170 VSUBS 0.026028f
C759 VTAIL.n171 VSUBS 0.013986f
C760 VTAIL.n172 VSUBS 0.014809f
C761 VTAIL.n173 VSUBS 0.033059f
C762 VTAIL.n174 VSUBS 0.081332f
C763 VTAIL.n175 VSUBS 0.014809f
C764 VTAIL.n176 VSUBS 0.027466f
C765 VTAIL.n177 VSUBS 0.06443f
C766 VTAIL.n178 VSUBS 0.061878f
C767 VTAIL.n179 VSUBS 0.246967f
C768 VTAIL.n180 VSUBS 0.027609f
C769 VTAIL.n181 VSUBS 0.026028f
C770 VTAIL.n182 VSUBS 0.013986f
C771 VTAIL.n183 VSUBS 0.033059f
C772 VTAIL.n184 VSUBS 0.014809f
C773 VTAIL.n185 VSUBS 0.026028f
C774 VTAIL.n186 VSUBS 0.013986f
C775 VTAIL.n187 VSUBS 0.033059f
C776 VTAIL.n188 VSUBS 0.014809f
C777 VTAIL.n189 VSUBS 0.7311f
C778 VTAIL.n190 VSUBS 0.013986f
C779 VTAIL.t0 VSUBS 0.070997f
C780 VTAIL.n191 VSUBS 0.148646f
C781 VTAIL.n192 VSUBS 0.024867f
C782 VTAIL.n193 VSUBS 0.024794f
C783 VTAIL.n194 VSUBS 0.033059f
C784 VTAIL.n195 VSUBS 0.014809f
C785 VTAIL.n196 VSUBS 0.013986f
C786 VTAIL.n197 VSUBS 0.026028f
C787 VTAIL.n198 VSUBS 0.026028f
C788 VTAIL.n199 VSUBS 0.013986f
C789 VTAIL.n200 VSUBS 0.014809f
C790 VTAIL.n201 VSUBS 0.033059f
C791 VTAIL.n202 VSUBS 0.033059f
C792 VTAIL.n203 VSUBS 0.014809f
C793 VTAIL.n204 VSUBS 0.013986f
C794 VTAIL.n205 VSUBS 0.026028f
C795 VTAIL.n206 VSUBS 0.026028f
C796 VTAIL.n207 VSUBS 0.013986f
C797 VTAIL.n208 VSUBS 0.014809f
C798 VTAIL.n209 VSUBS 0.033059f
C799 VTAIL.n210 VSUBS 0.081332f
C800 VTAIL.n211 VSUBS 0.014809f
C801 VTAIL.n212 VSUBS 0.027466f
C802 VTAIL.n213 VSUBS 0.06443f
C803 VTAIL.n214 VSUBS 0.061878f
C804 VTAIL.n215 VSUBS 0.246967f
C805 VTAIL.n216 VSUBS 0.027609f
C806 VTAIL.n217 VSUBS 0.026028f
C807 VTAIL.n218 VSUBS 0.013986f
C808 VTAIL.n219 VSUBS 0.033059f
C809 VTAIL.n220 VSUBS 0.014809f
C810 VTAIL.n221 VSUBS 0.026028f
C811 VTAIL.n222 VSUBS 0.013986f
C812 VTAIL.n223 VSUBS 0.033059f
C813 VTAIL.n224 VSUBS 0.014809f
C814 VTAIL.n225 VSUBS 0.7311f
C815 VTAIL.n226 VSUBS 0.013986f
C816 VTAIL.t1 VSUBS 0.070997f
C817 VTAIL.n227 VSUBS 0.148646f
C818 VTAIL.n228 VSUBS 0.024867f
C819 VTAIL.n229 VSUBS 0.024794f
C820 VTAIL.n230 VSUBS 0.033059f
C821 VTAIL.n231 VSUBS 0.014809f
C822 VTAIL.n232 VSUBS 0.013986f
C823 VTAIL.n233 VSUBS 0.026028f
C824 VTAIL.n234 VSUBS 0.026028f
C825 VTAIL.n235 VSUBS 0.013986f
C826 VTAIL.n236 VSUBS 0.014809f
C827 VTAIL.n237 VSUBS 0.033059f
C828 VTAIL.n238 VSUBS 0.033059f
C829 VTAIL.n239 VSUBS 0.014809f
C830 VTAIL.n240 VSUBS 0.013986f
C831 VTAIL.n241 VSUBS 0.026028f
C832 VTAIL.n242 VSUBS 0.026028f
C833 VTAIL.n243 VSUBS 0.013986f
C834 VTAIL.n244 VSUBS 0.014809f
C835 VTAIL.n245 VSUBS 0.033059f
C836 VTAIL.n246 VSUBS 0.081332f
C837 VTAIL.n247 VSUBS 0.014809f
C838 VTAIL.n248 VSUBS 0.027466f
C839 VTAIL.n249 VSUBS 0.06443f
C840 VTAIL.n250 VSUBS 0.061878f
C841 VTAIL.n251 VSUBS 1.26461f
C842 VTAIL.n252 VSUBS 0.027609f
C843 VTAIL.n253 VSUBS 0.026028f
C844 VTAIL.n254 VSUBS 0.013986f
C845 VTAIL.n255 VSUBS 0.033059f
C846 VTAIL.n256 VSUBS 0.014809f
C847 VTAIL.n257 VSUBS 0.026028f
C848 VTAIL.n258 VSUBS 0.013986f
C849 VTAIL.n259 VSUBS 0.033059f
C850 VTAIL.n260 VSUBS 0.014809f
C851 VTAIL.n261 VSUBS 0.7311f
C852 VTAIL.n262 VSUBS 0.013986f
C853 VTAIL.t4 VSUBS 0.070997f
C854 VTAIL.n263 VSUBS 0.148646f
C855 VTAIL.n264 VSUBS 0.024867f
C856 VTAIL.n265 VSUBS 0.024794f
C857 VTAIL.n266 VSUBS 0.033059f
C858 VTAIL.n267 VSUBS 0.014809f
C859 VTAIL.n268 VSUBS 0.013986f
C860 VTAIL.n269 VSUBS 0.026028f
C861 VTAIL.n270 VSUBS 0.026028f
C862 VTAIL.n271 VSUBS 0.013986f
C863 VTAIL.n272 VSUBS 0.014809f
C864 VTAIL.n273 VSUBS 0.033059f
C865 VTAIL.n274 VSUBS 0.033059f
C866 VTAIL.n275 VSUBS 0.014809f
C867 VTAIL.n276 VSUBS 0.013986f
C868 VTAIL.n277 VSUBS 0.026028f
C869 VTAIL.n278 VSUBS 0.026028f
C870 VTAIL.n279 VSUBS 0.013986f
C871 VTAIL.n280 VSUBS 0.014809f
C872 VTAIL.n281 VSUBS 0.033059f
C873 VTAIL.n282 VSUBS 0.081332f
C874 VTAIL.n283 VSUBS 0.014809f
C875 VTAIL.n284 VSUBS 0.027466f
C876 VTAIL.n285 VSUBS 0.06443f
C877 VTAIL.n286 VSUBS 0.061878f
C878 VTAIL.n287 VSUBS 1.16827f
C879 VDD2.t0 VSUBS 0.154824f
C880 VDD2.t2 VSUBS 0.154824f
C881 VDD2.n0 VSUBS 1.55884f
C882 VDD2.t1 VSUBS 0.154824f
C883 VDD2.t3 VSUBS 0.154824f
C884 VDD2.n1 VSUBS 1.09515f
C885 VDD2.n2 VSUBS 3.62962f
C886 VN.t1 VSUBS 2.03615f
C887 VN.t3 VSUBS 2.03124f
C888 VN.n0 VSUBS 1.34664f
C889 VN.t2 VSUBS 2.03615f
C890 VN.t0 VSUBS 2.03124f
C891 VN.n1 VSUBS 3.16087f
.ends

