* NGSPICE file created from diff_pair_sample_0413.ext - technology: sky130A

.subckt diff_pair_sample_0413 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.4017 ps=2.84 w=1.03 l=3.49
X1 VTAIL.t6 VN.t0 VDD2.t7 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0.16995 ps=1.36 w=1.03 l=3.49
X2 VDD1.t6 VP.t1 VTAIL.t15 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X3 VTAIL.t2 VN.t1 VDD2.t6 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0.16995 ps=1.36 w=1.03 l=3.49
X4 B.t11 B.t9 B.t10 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0 ps=0 w=1.03 l=3.49
X5 VDD2.t5 VN.t2 VTAIL.t3 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.4017 ps=2.84 w=1.03 l=3.49
X6 VDD1.t5 VP.t2 VTAIL.t11 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X7 VDD2.t4 VN.t3 VTAIL.t4 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.4017 ps=2.84 w=1.03 l=3.49
X8 VDD1.t4 VP.t3 VTAIL.t8 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.4017 ps=2.84 w=1.03 l=3.49
X9 VTAIL.t0 VN.t4 VDD2.t3 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X10 B.t8 B.t6 B.t7 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0 ps=0 w=1.03 l=3.49
X11 B.t5 B.t3 B.t4 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0 ps=0 w=1.03 l=3.49
X12 VTAIL.t9 VP.t4 VDD1.t3 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X13 VDD2.t2 VN.t5 VTAIL.t1 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X14 VTAIL.t5 VN.t6 VDD2.t1 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X15 VTAIL.t10 VP.t5 VDD1.t2 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0.16995 ps=1.36 w=1.03 l=3.49
X16 VDD2.t0 VN.t7 VTAIL.t7 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
X17 VTAIL.t12 VP.t6 VDD1.t1 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0.16995 ps=1.36 w=1.03 l=3.49
X18 B.t2 B.t0 B.t1 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.4017 pd=2.84 as=0 ps=0 w=1.03 l=3.49
X19 VTAIL.t13 VP.t7 VDD1.t0 w_n4790_n1174# sky130_fd_pr__pfet_01v8 ad=0.16995 pd=1.36 as=0.16995 ps=1.36 w=1.03 l=3.49
R0 VP.n24 VP.n23 161.3
R1 VP.n25 VP.n20 161.3
R2 VP.n27 VP.n26 161.3
R3 VP.n28 VP.n19 161.3
R4 VP.n30 VP.n29 161.3
R5 VP.n31 VP.n18 161.3
R6 VP.n34 VP.n33 161.3
R7 VP.n35 VP.n17 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n85 VP.n84 161.3
R16 VP.n83 VP.n1 161.3
R17 VP.n82 VP.n81 161.3
R18 VP.n80 VP.n2 161.3
R19 VP.n79 VP.n78 161.3
R20 VP.n77 VP.n3 161.3
R21 VP.n76 VP.n75 161.3
R22 VP.n74 VP.n4 161.3
R23 VP.n73 VP.n72 161.3
R24 VP.n70 VP.n5 161.3
R25 VP.n69 VP.n68 161.3
R26 VP.n67 VP.n6 161.3
R27 VP.n66 VP.n65 161.3
R28 VP.n64 VP.n7 161.3
R29 VP.n63 VP.n62 161.3
R30 VP.n61 VP.n60 161.3
R31 VP.n59 VP.n9 161.3
R32 VP.n58 VP.n57 161.3
R33 VP.n56 VP.n10 161.3
R34 VP.n55 VP.n54 161.3
R35 VP.n53 VP.n11 161.3
R36 VP.n52 VP.n51 161.3
R37 VP.n50 VP.n12 161.3
R38 VP.n49 VP.n48 78.8126
R39 VP.n86 VP.n0 78.8126
R40 VP.n47 VP.n13 78.8126
R41 VP.n54 VP.n10 56.5193
R42 VP.n39 VP.n15 56.5193
R43 VP.n78 VP.n2 56.5193
R44 VP.n22 VP.n21 54.5826
R45 VP.n49 VP.n47 46.8554
R46 VP.n22 VP.t5 40.6937
R47 VP.n65 VP.n6 40.4934
R48 VP.n69 VP.n6 40.4934
R49 VP.n30 VP.n19 40.4934
R50 VP.n26 VP.n19 40.4934
R51 VP.n52 VP.n12 24.4675
R52 VP.n53 VP.n52 24.4675
R53 VP.n54 VP.n53 24.4675
R54 VP.n58 VP.n10 24.4675
R55 VP.n59 VP.n58 24.4675
R56 VP.n60 VP.n59 24.4675
R57 VP.n64 VP.n63 24.4675
R58 VP.n65 VP.n64 24.4675
R59 VP.n70 VP.n69 24.4675
R60 VP.n72 VP.n70 24.4675
R61 VP.n76 VP.n4 24.4675
R62 VP.n77 VP.n76 24.4675
R63 VP.n78 VP.n77 24.4675
R64 VP.n82 VP.n2 24.4675
R65 VP.n83 VP.n82 24.4675
R66 VP.n84 VP.n83 24.4675
R67 VP.n43 VP.n15 24.4675
R68 VP.n44 VP.n43 24.4675
R69 VP.n45 VP.n44 24.4675
R70 VP.n31 VP.n30 24.4675
R71 VP.n33 VP.n31 24.4675
R72 VP.n37 VP.n17 24.4675
R73 VP.n38 VP.n37 24.4675
R74 VP.n39 VP.n38 24.4675
R75 VP.n25 VP.n24 24.4675
R76 VP.n26 VP.n25 24.4675
R77 VP.n63 VP.n8 20.0634
R78 VP.n72 VP.n71 20.0634
R79 VP.n33 VP.n32 20.0634
R80 VP.n24 VP.n21 20.0634
R81 VP.n48 VP.n12 11.2553
R82 VP.n84 VP.n0 11.2553
R83 VP.n45 VP.n13 11.2553
R84 VP.n48 VP.t6 7.11311
R85 VP.n8 VP.t2 7.11311
R86 VP.n71 VP.t4 7.11311
R87 VP.n0 VP.t3 7.11311
R88 VP.n13 VP.t0 7.11311
R89 VP.n32 VP.t7 7.11311
R90 VP.n21 VP.t1 7.11311
R91 VP.n60 VP.n8 4.40456
R92 VP.n71 VP.n4 4.40456
R93 VP.n32 VP.n17 4.40456
R94 VP.n23 VP.n22 3.11608
R95 VP.n47 VP.n46 0.354971
R96 VP.n50 VP.n49 0.354971
R97 VP.n86 VP.n85 0.354971
R98 VP VP.n86 0.26696
R99 VP.n23 VP.n20 0.189894
R100 VP.n27 VP.n20 0.189894
R101 VP.n28 VP.n27 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n29 VP.n18 0.189894
R104 VP.n34 VP.n18 0.189894
R105 VP.n35 VP.n34 0.189894
R106 VP.n36 VP.n35 0.189894
R107 VP.n36 VP.n16 0.189894
R108 VP.n40 VP.n16 0.189894
R109 VP.n41 VP.n40 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n42 VP.n14 0.189894
R112 VP.n46 VP.n14 0.189894
R113 VP.n51 VP.n50 0.189894
R114 VP.n51 VP.n11 0.189894
R115 VP.n55 VP.n11 0.189894
R116 VP.n56 VP.n55 0.189894
R117 VP.n57 VP.n56 0.189894
R118 VP.n57 VP.n9 0.189894
R119 VP.n61 VP.n9 0.189894
R120 VP.n62 VP.n61 0.189894
R121 VP.n62 VP.n7 0.189894
R122 VP.n66 VP.n7 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n68 VP.n67 0.189894
R125 VP.n68 VP.n5 0.189894
R126 VP.n73 VP.n5 0.189894
R127 VP.n74 VP.n73 0.189894
R128 VP.n75 VP.n74 0.189894
R129 VP.n75 VP.n3 0.189894
R130 VP.n79 VP.n3 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n81 VP.n80 0.189894
R133 VP.n81 VP.n1 0.189894
R134 VP.n85 VP.n1 0.189894
R135 VTAIL.n15 VTAIL.t3 371.166
R136 VTAIL.n2 VTAIL.t2 371.166
R137 VTAIL.n3 VTAIL.t8 371.166
R138 VTAIL.n6 VTAIL.t12 371.166
R139 VTAIL.n14 VTAIL.t14 371.166
R140 VTAIL.n11 VTAIL.t10 371.166
R141 VTAIL.n10 VTAIL.t4 371.166
R142 VTAIL.n7 VTAIL.t6 371.166
R143 VTAIL.n1 VTAIL.n0 328.228
R144 VTAIL.n5 VTAIL.n4 328.228
R145 VTAIL.n13 VTAIL.n12 328.226
R146 VTAIL.n9 VTAIL.n8 328.226
R147 VTAIL.n0 VTAIL.t1 31.5588
R148 VTAIL.n0 VTAIL.t0 31.5588
R149 VTAIL.n4 VTAIL.t11 31.5588
R150 VTAIL.n4 VTAIL.t9 31.5588
R151 VTAIL.n12 VTAIL.t15 31.5588
R152 VTAIL.n12 VTAIL.t13 31.5588
R153 VTAIL.n8 VTAIL.t7 31.5588
R154 VTAIL.n8 VTAIL.t5 31.5588
R155 VTAIL.n15 VTAIL.n14 16.5479
R156 VTAIL.n7 VTAIL.n6 16.5479
R157 VTAIL.n9 VTAIL.n7 3.2936
R158 VTAIL.n10 VTAIL.n9 3.2936
R159 VTAIL.n13 VTAIL.n11 3.2936
R160 VTAIL.n14 VTAIL.n13 3.2936
R161 VTAIL.n6 VTAIL.n5 3.2936
R162 VTAIL.n5 VTAIL.n3 3.2936
R163 VTAIL.n2 VTAIL.n1 3.2936
R164 VTAIL VTAIL.n15 3.23541
R165 VTAIL.n11 VTAIL.n10 0.470328
R166 VTAIL.n3 VTAIL.n2 0.470328
R167 VTAIL VTAIL.n1 0.0586897
R168 VDD1 VDD1.n0 346.611
R169 VDD1.n3 VDD1.n2 346.498
R170 VDD1.n3 VDD1.n1 346.498
R171 VDD1.n5 VDD1.n4 344.906
R172 VDD1.n5 VDD1.n3 40.0052
R173 VDD1.n4 VDD1.t0 31.5588
R174 VDD1.n4 VDD1.t7 31.5588
R175 VDD1.n0 VDD1.t2 31.5588
R176 VDD1.n0 VDD1.t6 31.5588
R177 VDD1.n2 VDD1.t3 31.5588
R178 VDD1.n2 VDD1.t4 31.5588
R179 VDD1.n1 VDD1.t1 31.5588
R180 VDD1.n1 VDD1.t5 31.5588
R181 VDD1 VDD1.n5 1.58886
R182 VN.n68 VN.n67 161.3
R183 VN.n66 VN.n36 161.3
R184 VN.n65 VN.n64 161.3
R185 VN.n63 VN.n37 161.3
R186 VN.n62 VN.n61 161.3
R187 VN.n60 VN.n38 161.3
R188 VN.n59 VN.n58 161.3
R189 VN.n57 VN.n39 161.3
R190 VN.n56 VN.n55 161.3
R191 VN.n54 VN.n40 161.3
R192 VN.n53 VN.n52 161.3
R193 VN.n51 VN.n42 161.3
R194 VN.n50 VN.n49 161.3
R195 VN.n48 VN.n43 161.3
R196 VN.n47 VN.n46 161.3
R197 VN.n33 VN.n32 161.3
R198 VN.n31 VN.n1 161.3
R199 VN.n30 VN.n29 161.3
R200 VN.n28 VN.n2 161.3
R201 VN.n27 VN.n26 161.3
R202 VN.n25 VN.n3 161.3
R203 VN.n24 VN.n23 161.3
R204 VN.n22 VN.n4 161.3
R205 VN.n21 VN.n20 161.3
R206 VN.n18 VN.n5 161.3
R207 VN.n17 VN.n16 161.3
R208 VN.n15 VN.n6 161.3
R209 VN.n14 VN.n13 161.3
R210 VN.n12 VN.n7 161.3
R211 VN.n11 VN.n10 161.3
R212 VN.n34 VN.n0 78.8126
R213 VN.n69 VN.n35 78.8126
R214 VN.n26 VN.n2 56.5193
R215 VN.n61 VN.n37 56.5193
R216 VN.n45 VN.n44 54.5825
R217 VN.n9 VN.n8 54.5825
R218 VN VN.n69 47.0207
R219 VN.n45 VN.t3 40.6939
R220 VN.n9 VN.t1 40.6939
R221 VN.n13 VN.n6 40.4934
R222 VN.n17 VN.n6 40.4934
R223 VN.n49 VN.n42 40.4934
R224 VN.n53 VN.n42 40.4934
R225 VN.n12 VN.n11 24.4675
R226 VN.n13 VN.n12 24.4675
R227 VN.n18 VN.n17 24.4675
R228 VN.n20 VN.n18 24.4675
R229 VN.n24 VN.n4 24.4675
R230 VN.n25 VN.n24 24.4675
R231 VN.n26 VN.n25 24.4675
R232 VN.n30 VN.n2 24.4675
R233 VN.n31 VN.n30 24.4675
R234 VN.n32 VN.n31 24.4675
R235 VN.n49 VN.n48 24.4675
R236 VN.n48 VN.n47 24.4675
R237 VN.n61 VN.n60 24.4675
R238 VN.n60 VN.n59 24.4675
R239 VN.n59 VN.n39 24.4675
R240 VN.n55 VN.n54 24.4675
R241 VN.n54 VN.n53 24.4675
R242 VN.n67 VN.n66 24.4675
R243 VN.n66 VN.n65 24.4675
R244 VN.n65 VN.n37 24.4675
R245 VN.n11 VN.n8 20.0634
R246 VN.n20 VN.n19 20.0634
R247 VN.n47 VN.n44 20.0634
R248 VN.n55 VN.n41 20.0634
R249 VN.n32 VN.n0 11.2553
R250 VN.n67 VN.n35 11.2553
R251 VN.n8 VN.t5 7.11311
R252 VN.n19 VN.t4 7.11311
R253 VN.n0 VN.t2 7.11311
R254 VN.n44 VN.t6 7.11311
R255 VN.n41 VN.t7 7.11311
R256 VN.n35 VN.t0 7.11311
R257 VN.n19 VN.n4 4.40456
R258 VN.n41 VN.n39 4.40456
R259 VN.n46 VN.n45 3.1161
R260 VN.n10 VN.n9 3.1161
R261 VN.n69 VN.n68 0.354971
R262 VN.n34 VN.n33 0.354971
R263 VN VN.n34 0.26696
R264 VN.n68 VN.n36 0.189894
R265 VN.n64 VN.n36 0.189894
R266 VN.n64 VN.n63 0.189894
R267 VN.n63 VN.n62 0.189894
R268 VN.n62 VN.n38 0.189894
R269 VN.n58 VN.n38 0.189894
R270 VN.n58 VN.n57 0.189894
R271 VN.n57 VN.n56 0.189894
R272 VN.n56 VN.n40 0.189894
R273 VN.n52 VN.n40 0.189894
R274 VN.n52 VN.n51 0.189894
R275 VN.n51 VN.n50 0.189894
R276 VN.n50 VN.n43 0.189894
R277 VN.n46 VN.n43 0.189894
R278 VN.n10 VN.n7 0.189894
R279 VN.n14 VN.n7 0.189894
R280 VN.n15 VN.n14 0.189894
R281 VN.n16 VN.n15 0.189894
R282 VN.n16 VN.n5 0.189894
R283 VN.n21 VN.n5 0.189894
R284 VN.n22 VN.n21 0.189894
R285 VN.n23 VN.n22 0.189894
R286 VN.n23 VN.n3 0.189894
R287 VN.n27 VN.n3 0.189894
R288 VN.n28 VN.n27 0.189894
R289 VN.n29 VN.n28 0.189894
R290 VN.n29 VN.n1 0.189894
R291 VN.n33 VN.n1 0.189894
R292 VDD2.n2 VDD2.n1 346.498
R293 VDD2.n2 VDD2.n0 346.498
R294 VDD2 VDD2.n5 346.495
R295 VDD2.n4 VDD2.n3 344.906
R296 VDD2.n4 VDD2.n2 39.4222
R297 VDD2.n5 VDD2.t1 31.5588
R298 VDD2.n5 VDD2.t4 31.5588
R299 VDD2.n3 VDD2.t7 31.5588
R300 VDD2.n3 VDD2.t0 31.5588
R301 VDD2.n1 VDD2.t3 31.5588
R302 VDD2.n1 VDD2.t5 31.5588
R303 VDD2.n0 VDD2.t6 31.5588
R304 VDD2.n0 VDD2.t2 31.5588
R305 VDD2 VDD2.n4 1.70524
R306 B.n305 B.n118 585
R307 B.n304 B.n303 585
R308 B.n302 B.n119 585
R309 B.n301 B.n300 585
R310 B.n299 B.n120 585
R311 B.n298 B.n297 585
R312 B.n296 B.n121 585
R313 B.n295 B.n294 585
R314 B.n293 B.n122 585
R315 B.n291 B.n290 585
R316 B.n289 B.n125 585
R317 B.n288 B.n287 585
R318 B.n286 B.n126 585
R319 B.n285 B.n284 585
R320 B.n283 B.n127 585
R321 B.n282 B.n281 585
R322 B.n280 B.n128 585
R323 B.n279 B.n278 585
R324 B.n277 B.n129 585
R325 B.n276 B.n275 585
R326 B.n271 B.n130 585
R327 B.n270 B.n269 585
R328 B.n268 B.n131 585
R329 B.n267 B.n266 585
R330 B.n265 B.n132 585
R331 B.n264 B.n263 585
R332 B.n262 B.n133 585
R333 B.n261 B.n260 585
R334 B.n307 B.n306 585
R335 B.n308 B.n117 585
R336 B.n310 B.n309 585
R337 B.n311 B.n116 585
R338 B.n313 B.n312 585
R339 B.n314 B.n115 585
R340 B.n316 B.n315 585
R341 B.n317 B.n114 585
R342 B.n319 B.n318 585
R343 B.n320 B.n113 585
R344 B.n322 B.n321 585
R345 B.n323 B.n112 585
R346 B.n325 B.n324 585
R347 B.n326 B.n111 585
R348 B.n328 B.n327 585
R349 B.n329 B.n110 585
R350 B.n331 B.n330 585
R351 B.n332 B.n109 585
R352 B.n334 B.n333 585
R353 B.n335 B.n108 585
R354 B.n337 B.n336 585
R355 B.n338 B.n107 585
R356 B.n340 B.n339 585
R357 B.n341 B.n106 585
R358 B.n343 B.n342 585
R359 B.n344 B.n105 585
R360 B.n346 B.n345 585
R361 B.n347 B.n104 585
R362 B.n349 B.n348 585
R363 B.n350 B.n103 585
R364 B.n352 B.n351 585
R365 B.n353 B.n102 585
R366 B.n355 B.n354 585
R367 B.n356 B.n101 585
R368 B.n358 B.n357 585
R369 B.n359 B.n100 585
R370 B.n361 B.n360 585
R371 B.n362 B.n99 585
R372 B.n364 B.n363 585
R373 B.n365 B.n98 585
R374 B.n367 B.n366 585
R375 B.n368 B.n97 585
R376 B.n370 B.n369 585
R377 B.n371 B.n96 585
R378 B.n373 B.n372 585
R379 B.n374 B.n95 585
R380 B.n376 B.n375 585
R381 B.n377 B.n94 585
R382 B.n379 B.n378 585
R383 B.n380 B.n93 585
R384 B.n382 B.n381 585
R385 B.n383 B.n92 585
R386 B.n385 B.n384 585
R387 B.n386 B.n91 585
R388 B.n388 B.n387 585
R389 B.n389 B.n90 585
R390 B.n391 B.n390 585
R391 B.n392 B.n89 585
R392 B.n394 B.n393 585
R393 B.n395 B.n88 585
R394 B.n397 B.n396 585
R395 B.n398 B.n87 585
R396 B.n400 B.n399 585
R397 B.n401 B.n86 585
R398 B.n403 B.n402 585
R399 B.n404 B.n85 585
R400 B.n406 B.n405 585
R401 B.n407 B.n84 585
R402 B.n409 B.n408 585
R403 B.n410 B.n83 585
R404 B.n412 B.n411 585
R405 B.n413 B.n82 585
R406 B.n415 B.n414 585
R407 B.n416 B.n81 585
R408 B.n418 B.n417 585
R409 B.n419 B.n80 585
R410 B.n421 B.n420 585
R411 B.n422 B.n79 585
R412 B.n424 B.n423 585
R413 B.n425 B.n78 585
R414 B.n427 B.n426 585
R415 B.n428 B.n77 585
R416 B.n430 B.n429 585
R417 B.n431 B.n76 585
R418 B.n433 B.n432 585
R419 B.n434 B.n75 585
R420 B.n436 B.n435 585
R421 B.n437 B.n74 585
R422 B.n439 B.n438 585
R423 B.n440 B.n73 585
R424 B.n442 B.n441 585
R425 B.n443 B.n72 585
R426 B.n445 B.n444 585
R427 B.n446 B.n71 585
R428 B.n448 B.n447 585
R429 B.n449 B.n70 585
R430 B.n451 B.n450 585
R431 B.n452 B.n69 585
R432 B.n454 B.n453 585
R433 B.n455 B.n68 585
R434 B.n457 B.n456 585
R435 B.n458 B.n67 585
R436 B.n460 B.n459 585
R437 B.n461 B.n66 585
R438 B.n463 B.n462 585
R439 B.n464 B.n65 585
R440 B.n466 B.n465 585
R441 B.n467 B.n64 585
R442 B.n469 B.n468 585
R443 B.n470 B.n63 585
R444 B.n472 B.n471 585
R445 B.n473 B.n62 585
R446 B.n475 B.n474 585
R447 B.n476 B.n61 585
R448 B.n478 B.n477 585
R449 B.n479 B.n60 585
R450 B.n481 B.n480 585
R451 B.n482 B.n59 585
R452 B.n484 B.n483 585
R453 B.n485 B.n58 585
R454 B.n487 B.n486 585
R455 B.n488 B.n57 585
R456 B.n490 B.n489 585
R457 B.n491 B.n56 585
R458 B.n493 B.n492 585
R459 B.n494 B.n55 585
R460 B.n496 B.n495 585
R461 B.n497 B.n54 585
R462 B.n499 B.n498 585
R463 B.n500 B.n53 585
R464 B.n543 B.n34 585
R465 B.n542 B.n541 585
R466 B.n540 B.n35 585
R467 B.n539 B.n538 585
R468 B.n537 B.n36 585
R469 B.n536 B.n535 585
R470 B.n534 B.n37 585
R471 B.n533 B.n532 585
R472 B.n531 B.n38 585
R473 B.n530 B.n529 585
R474 B.n528 B.n39 585
R475 B.n527 B.n526 585
R476 B.n525 B.n43 585
R477 B.n524 B.n523 585
R478 B.n522 B.n44 585
R479 B.n521 B.n520 585
R480 B.n519 B.n45 585
R481 B.n518 B.n517 585
R482 B.n516 B.n46 585
R483 B.n514 B.n513 585
R484 B.n512 B.n49 585
R485 B.n511 B.n510 585
R486 B.n509 B.n50 585
R487 B.n508 B.n507 585
R488 B.n506 B.n51 585
R489 B.n505 B.n504 585
R490 B.n503 B.n52 585
R491 B.n502 B.n501 585
R492 B.n545 B.n544 585
R493 B.n546 B.n33 585
R494 B.n548 B.n547 585
R495 B.n549 B.n32 585
R496 B.n551 B.n550 585
R497 B.n552 B.n31 585
R498 B.n554 B.n553 585
R499 B.n555 B.n30 585
R500 B.n557 B.n556 585
R501 B.n558 B.n29 585
R502 B.n560 B.n559 585
R503 B.n561 B.n28 585
R504 B.n563 B.n562 585
R505 B.n564 B.n27 585
R506 B.n566 B.n565 585
R507 B.n567 B.n26 585
R508 B.n569 B.n568 585
R509 B.n570 B.n25 585
R510 B.n572 B.n571 585
R511 B.n573 B.n24 585
R512 B.n575 B.n574 585
R513 B.n576 B.n23 585
R514 B.n578 B.n577 585
R515 B.n579 B.n22 585
R516 B.n581 B.n580 585
R517 B.n582 B.n21 585
R518 B.n584 B.n583 585
R519 B.n585 B.n20 585
R520 B.n587 B.n586 585
R521 B.n588 B.n19 585
R522 B.n590 B.n589 585
R523 B.n591 B.n18 585
R524 B.n593 B.n592 585
R525 B.n594 B.n17 585
R526 B.n596 B.n595 585
R527 B.n597 B.n16 585
R528 B.n599 B.n598 585
R529 B.n600 B.n15 585
R530 B.n602 B.n601 585
R531 B.n603 B.n14 585
R532 B.n605 B.n604 585
R533 B.n606 B.n13 585
R534 B.n608 B.n607 585
R535 B.n609 B.n12 585
R536 B.n611 B.n610 585
R537 B.n612 B.n11 585
R538 B.n614 B.n613 585
R539 B.n615 B.n10 585
R540 B.n617 B.n616 585
R541 B.n618 B.n9 585
R542 B.n620 B.n619 585
R543 B.n621 B.n8 585
R544 B.n623 B.n622 585
R545 B.n624 B.n7 585
R546 B.n626 B.n625 585
R547 B.n627 B.n6 585
R548 B.n629 B.n628 585
R549 B.n630 B.n5 585
R550 B.n632 B.n631 585
R551 B.n633 B.n4 585
R552 B.n635 B.n634 585
R553 B.n636 B.n3 585
R554 B.n638 B.n637 585
R555 B.n639 B.n0 585
R556 B.n2 B.n1 585
R557 B.n166 B.n165 585
R558 B.n168 B.n167 585
R559 B.n169 B.n164 585
R560 B.n171 B.n170 585
R561 B.n172 B.n163 585
R562 B.n174 B.n173 585
R563 B.n175 B.n162 585
R564 B.n177 B.n176 585
R565 B.n178 B.n161 585
R566 B.n180 B.n179 585
R567 B.n181 B.n160 585
R568 B.n183 B.n182 585
R569 B.n184 B.n159 585
R570 B.n186 B.n185 585
R571 B.n187 B.n158 585
R572 B.n189 B.n188 585
R573 B.n190 B.n157 585
R574 B.n192 B.n191 585
R575 B.n193 B.n156 585
R576 B.n195 B.n194 585
R577 B.n196 B.n155 585
R578 B.n198 B.n197 585
R579 B.n199 B.n154 585
R580 B.n201 B.n200 585
R581 B.n202 B.n153 585
R582 B.n204 B.n203 585
R583 B.n205 B.n152 585
R584 B.n207 B.n206 585
R585 B.n208 B.n151 585
R586 B.n210 B.n209 585
R587 B.n211 B.n150 585
R588 B.n213 B.n212 585
R589 B.n214 B.n149 585
R590 B.n216 B.n215 585
R591 B.n217 B.n148 585
R592 B.n219 B.n218 585
R593 B.n220 B.n147 585
R594 B.n222 B.n221 585
R595 B.n223 B.n146 585
R596 B.n225 B.n224 585
R597 B.n226 B.n145 585
R598 B.n228 B.n227 585
R599 B.n229 B.n144 585
R600 B.n231 B.n230 585
R601 B.n232 B.n143 585
R602 B.n234 B.n233 585
R603 B.n235 B.n142 585
R604 B.n237 B.n236 585
R605 B.n238 B.n141 585
R606 B.n240 B.n239 585
R607 B.n241 B.n140 585
R608 B.n243 B.n242 585
R609 B.n244 B.n139 585
R610 B.n246 B.n245 585
R611 B.n247 B.n138 585
R612 B.n249 B.n248 585
R613 B.n250 B.n137 585
R614 B.n252 B.n251 585
R615 B.n253 B.n136 585
R616 B.n255 B.n254 585
R617 B.n256 B.n135 585
R618 B.n258 B.n257 585
R619 B.n259 B.n134 585
R620 B.n261 B.n134 487.695
R621 B.n307 B.n118 487.695
R622 B.n501 B.n500 487.695
R623 B.n544 B.n543 487.695
R624 B.n272 B.t7 435.865
R625 B.n123 B.t10 435.865
R626 B.n47 B.t2 435.865
R627 B.n40 B.t5 435.865
R628 B.n273 B.t8 361.781
R629 B.n124 B.t11 361.781
R630 B.n48 B.t1 361.781
R631 B.n41 B.t4 361.781
R632 B.n641 B.n640 256.663
R633 B.n640 B.n639 235.042
R634 B.n640 B.n2 235.042
R635 B.n272 B.t6 209.761
R636 B.n123 B.t9 209.761
R637 B.n47 B.t0 209.761
R638 B.n40 B.t3 209.761
R639 B.n262 B.n261 163.367
R640 B.n263 B.n262 163.367
R641 B.n263 B.n132 163.367
R642 B.n267 B.n132 163.367
R643 B.n268 B.n267 163.367
R644 B.n269 B.n268 163.367
R645 B.n269 B.n130 163.367
R646 B.n276 B.n130 163.367
R647 B.n277 B.n276 163.367
R648 B.n278 B.n277 163.367
R649 B.n278 B.n128 163.367
R650 B.n282 B.n128 163.367
R651 B.n283 B.n282 163.367
R652 B.n284 B.n283 163.367
R653 B.n284 B.n126 163.367
R654 B.n288 B.n126 163.367
R655 B.n289 B.n288 163.367
R656 B.n290 B.n289 163.367
R657 B.n290 B.n122 163.367
R658 B.n295 B.n122 163.367
R659 B.n296 B.n295 163.367
R660 B.n297 B.n296 163.367
R661 B.n297 B.n120 163.367
R662 B.n301 B.n120 163.367
R663 B.n302 B.n301 163.367
R664 B.n303 B.n302 163.367
R665 B.n303 B.n118 163.367
R666 B.n500 B.n499 163.367
R667 B.n499 B.n54 163.367
R668 B.n495 B.n54 163.367
R669 B.n495 B.n494 163.367
R670 B.n494 B.n493 163.367
R671 B.n493 B.n56 163.367
R672 B.n489 B.n56 163.367
R673 B.n489 B.n488 163.367
R674 B.n488 B.n487 163.367
R675 B.n487 B.n58 163.367
R676 B.n483 B.n58 163.367
R677 B.n483 B.n482 163.367
R678 B.n482 B.n481 163.367
R679 B.n481 B.n60 163.367
R680 B.n477 B.n60 163.367
R681 B.n477 B.n476 163.367
R682 B.n476 B.n475 163.367
R683 B.n475 B.n62 163.367
R684 B.n471 B.n62 163.367
R685 B.n471 B.n470 163.367
R686 B.n470 B.n469 163.367
R687 B.n469 B.n64 163.367
R688 B.n465 B.n64 163.367
R689 B.n465 B.n464 163.367
R690 B.n464 B.n463 163.367
R691 B.n463 B.n66 163.367
R692 B.n459 B.n66 163.367
R693 B.n459 B.n458 163.367
R694 B.n458 B.n457 163.367
R695 B.n457 B.n68 163.367
R696 B.n453 B.n68 163.367
R697 B.n453 B.n452 163.367
R698 B.n452 B.n451 163.367
R699 B.n451 B.n70 163.367
R700 B.n447 B.n70 163.367
R701 B.n447 B.n446 163.367
R702 B.n446 B.n445 163.367
R703 B.n445 B.n72 163.367
R704 B.n441 B.n72 163.367
R705 B.n441 B.n440 163.367
R706 B.n440 B.n439 163.367
R707 B.n439 B.n74 163.367
R708 B.n435 B.n74 163.367
R709 B.n435 B.n434 163.367
R710 B.n434 B.n433 163.367
R711 B.n433 B.n76 163.367
R712 B.n429 B.n76 163.367
R713 B.n429 B.n428 163.367
R714 B.n428 B.n427 163.367
R715 B.n427 B.n78 163.367
R716 B.n423 B.n78 163.367
R717 B.n423 B.n422 163.367
R718 B.n422 B.n421 163.367
R719 B.n421 B.n80 163.367
R720 B.n417 B.n80 163.367
R721 B.n417 B.n416 163.367
R722 B.n416 B.n415 163.367
R723 B.n415 B.n82 163.367
R724 B.n411 B.n82 163.367
R725 B.n411 B.n410 163.367
R726 B.n410 B.n409 163.367
R727 B.n409 B.n84 163.367
R728 B.n405 B.n84 163.367
R729 B.n405 B.n404 163.367
R730 B.n404 B.n403 163.367
R731 B.n403 B.n86 163.367
R732 B.n399 B.n86 163.367
R733 B.n399 B.n398 163.367
R734 B.n398 B.n397 163.367
R735 B.n397 B.n88 163.367
R736 B.n393 B.n88 163.367
R737 B.n393 B.n392 163.367
R738 B.n392 B.n391 163.367
R739 B.n391 B.n90 163.367
R740 B.n387 B.n90 163.367
R741 B.n387 B.n386 163.367
R742 B.n386 B.n385 163.367
R743 B.n385 B.n92 163.367
R744 B.n381 B.n92 163.367
R745 B.n381 B.n380 163.367
R746 B.n380 B.n379 163.367
R747 B.n379 B.n94 163.367
R748 B.n375 B.n94 163.367
R749 B.n375 B.n374 163.367
R750 B.n374 B.n373 163.367
R751 B.n373 B.n96 163.367
R752 B.n369 B.n96 163.367
R753 B.n369 B.n368 163.367
R754 B.n368 B.n367 163.367
R755 B.n367 B.n98 163.367
R756 B.n363 B.n98 163.367
R757 B.n363 B.n362 163.367
R758 B.n362 B.n361 163.367
R759 B.n361 B.n100 163.367
R760 B.n357 B.n100 163.367
R761 B.n357 B.n356 163.367
R762 B.n356 B.n355 163.367
R763 B.n355 B.n102 163.367
R764 B.n351 B.n102 163.367
R765 B.n351 B.n350 163.367
R766 B.n350 B.n349 163.367
R767 B.n349 B.n104 163.367
R768 B.n345 B.n104 163.367
R769 B.n345 B.n344 163.367
R770 B.n344 B.n343 163.367
R771 B.n343 B.n106 163.367
R772 B.n339 B.n106 163.367
R773 B.n339 B.n338 163.367
R774 B.n338 B.n337 163.367
R775 B.n337 B.n108 163.367
R776 B.n333 B.n108 163.367
R777 B.n333 B.n332 163.367
R778 B.n332 B.n331 163.367
R779 B.n331 B.n110 163.367
R780 B.n327 B.n110 163.367
R781 B.n327 B.n326 163.367
R782 B.n326 B.n325 163.367
R783 B.n325 B.n112 163.367
R784 B.n321 B.n112 163.367
R785 B.n321 B.n320 163.367
R786 B.n320 B.n319 163.367
R787 B.n319 B.n114 163.367
R788 B.n315 B.n114 163.367
R789 B.n315 B.n314 163.367
R790 B.n314 B.n313 163.367
R791 B.n313 B.n116 163.367
R792 B.n309 B.n116 163.367
R793 B.n309 B.n308 163.367
R794 B.n308 B.n307 163.367
R795 B.n543 B.n542 163.367
R796 B.n542 B.n35 163.367
R797 B.n538 B.n35 163.367
R798 B.n538 B.n537 163.367
R799 B.n537 B.n536 163.367
R800 B.n536 B.n37 163.367
R801 B.n532 B.n37 163.367
R802 B.n532 B.n531 163.367
R803 B.n531 B.n530 163.367
R804 B.n530 B.n39 163.367
R805 B.n526 B.n39 163.367
R806 B.n526 B.n525 163.367
R807 B.n525 B.n524 163.367
R808 B.n524 B.n44 163.367
R809 B.n520 B.n44 163.367
R810 B.n520 B.n519 163.367
R811 B.n519 B.n518 163.367
R812 B.n518 B.n46 163.367
R813 B.n513 B.n46 163.367
R814 B.n513 B.n512 163.367
R815 B.n512 B.n511 163.367
R816 B.n511 B.n50 163.367
R817 B.n507 B.n50 163.367
R818 B.n507 B.n506 163.367
R819 B.n506 B.n505 163.367
R820 B.n505 B.n52 163.367
R821 B.n501 B.n52 163.367
R822 B.n544 B.n33 163.367
R823 B.n548 B.n33 163.367
R824 B.n549 B.n548 163.367
R825 B.n550 B.n549 163.367
R826 B.n550 B.n31 163.367
R827 B.n554 B.n31 163.367
R828 B.n555 B.n554 163.367
R829 B.n556 B.n555 163.367
R830 B.n556 B.n29 163.367
R831 B.n560 B.n29 163.367
R832 B.n561 B.n560 163.367
R833 B.n562 B.n561 163.367
R834 B.n562 B.n27 163.367
R835 B.n566 B.n27 163.367
R836 B.n567 B.n566 163.367
R837 B.n568 B.n567 163.367
R838 B.n568 B.n25 163.367
R839 B.n572 B.n25 163.367
R840 B.n573 B.n572 163.367
R841 B.n574 B.n573 163.367
R842 B.n574 B.n23 163.367
R843 B.n578 B.n23 163.367
R844 B.n579 B.n578 163.367
R845 B.n580 B.n579 163.367
R846 B.n580 B.n21 163.367
R847 B.n584 B.n21 163.367
R848 B.n585 B.n584 163.367
R849 B.n586 B.n585 163.367
R850 B.n586 B.n19 163.367
R851 B.n590 B.n19 163.367
R852 B.n591 B.n590 163.367
R853 B.n592 B.n591 163.367
R854 B.n592 B.n17 163.367
R855 B.n596 B.n17 163.367
R856 B.n597 B.n596 163.367
R857 B.n598 B.n597 163.367
R858 B.n598 B.n15 163.367
R859 B.n602 B.n15 163.367
R860 B.n603 B.n602 163.367
R861 B.n604 B.n603 163.367
R862 B.n604 B.n13 163.367
R863 B.n608 B.n13 163.367
R864 B.n609 B.n608 163.367
R865 B.n610 B.n609 163.367
R866 B.n610 B.n11 163.367
R867 B.n614 B.n11 163.367
R868 B.n615 B.n614 163.367
R869 B.n616 B.n615 163.367
R870 B.n616 B.n9 163.367
R871 B.n620 B.n9 163.367
R872 B.n621 B.n620 163.367
R873 B.n622 B.n621 163.367
R874 B.n622 B.n7 163.367
R875 B.n626 B.n7 163.367
R876 B.n627 B.n626 163.367
R877 B.n628 B.n627 163.367
R878 B.n628 B.n5 163.367
R879 B.n632 B.n5 163.367
R880 B.n633 B.n632 163.367
R881 B.n634 B.n633 163.367
R882 B.n634 B.n3 163.367
R883 B.n638 B.n3 163.367
R884 B.n639 B.n638 163.367
R885 B.n166 B.n2 163.367
R886 B.n167 B.n166 163.367
R887 B.n167 B.n164 163.367
R888 B.n171 B.n164 163.367
R889 B.n172 B.n171 163.367
R890 B.n173 B.n172 163.367
R891 B.n173 B.n162 163.367
R892 B.n177 B.n162 163.367
R893 B.n178 B.n177 163.367
R894 B.n179 B.n178 163.367
R895 B.n179 B.n160 163.367
R896 B.n183 B.n160 163.367
R897 B.n184 B.n183 163.367
R898 B.n185 B.n184 163.367
R899 B.n185 B.n158 163.367
R900 B.n189 B.n158 163.367
R901 B.n190 B.n189 163.367
R902 B.n191 B.n190 163.367
R903 B.n191 B.n156 163.367
R904 B.n195 B.n156 163.367
R905 B.n196 B.n195 163.367
R906 B.n197 B.n196 163.367
R907 B.n197 B.n154 163.367
R908 B.n201 B.n154 163.367
R909 B.n202 B.n201 163.367
R910 B.n203 B.n202 163.367
R911 B.n203 B.n152 163.367
R912 B.n207 B.n152 163.367
R913 B.n208 B.n207 163.367
R914 B.n209 B.n208 163.367
R915 B.n209 B.n150 163.367
R916 B.n213 B.n150 163.367
R917 B.n214 B.n213 163.367
R918 B.n215 B.n214 163.367
R919 B.n215 B.n148 163.367
R920 B.n219 B.n148 163.367
R921 B.n220 B.n219 163.367
R922 B.n221 B.n220 163.367
R923 B.n221 B.n146 163.367
R924 B.n225 B.n146 163.367
R925 B.n226 B.n225 163.367
R926 B.n227 B.n226 163.367
R927 B.n227 B.n144 163.367
R928 B.n231 B.n144 163.367
R929 B.n232 B.n231 163.367
R930 B.n233 B.n232 163.367
R931 B.n233 B.n142 163.367
R932 B.n237 B.n142 163.367
R933 B.n238 B.n237 163.367
R934 B.n239 B.n238 163.367
R935 B.n239 B.n140 163.367
R936 B.n243 B.n140 163.367
R937 B.n244 B.n243 163.367
R938 B.n245 B.n244 163.367
R939 B.n245 B.n138 163.367
R940 B.n249 B.n138 163.367
R941 B.n250 B.n249 163.367
R942 B.n251 B.n250 163.367
R943 B.n251 B.n136 163.367
R944 B.n255 B.n136 163.367
R945 B.n256 B.n255 163.367
R946 B.n257 B.n256 163.367
R947 B.n257 B.n134 163.367
R948 B.n273 B.n272 74.0854
R949 B.n124 B.n123 74.0854
R950 B.n48 B.n47 74.0854
R951 B.n41 B.n40 74.0854
R952 B.n274 B.n273 59.5399
R953 B.n292 B.n124 59.5399
R954 B.n515 B.n48 59.5399
R955 B.n42 B.n41 59.5399
R956 B.n545 B.n34 31.6883
R957 B.n502 B.n53 31.6883
R958 B.n306 B.n305 31.6883
R959 B.n260 B.n259 31.6883
R960 B B.n641 18.0485
R961 B.n546 B.n545 10.6151
R962 B.n547 B.n546 10.6151
R963 B.n547 B.n32 10.6151
R964 B.n551 B.n32 10.6151
R965 B.n552 B.n551 10.6151
R966 B.n553 B.n552 10.6151
R967 B.n553 B.n30 10.6151
R968 B.n557 B.n30 10.6151
R969 B.n558 B.n557 10.6151
R970 B.n559 B.n558 10.6151
R971 B.n559 B.n28 10.6151
R972 B.n563 B.n28 10.6151
R973 B.n564 B.n563 10.6151
R974 B.n565 B.n564 10.6151
R975 B.n565 B.n26 10.6151
R976 B.n569 B.n26 10.6151
R977 B.n570 B.n569 10.6151
R978 B.n571 B.n570 10.6151
R979 B.n571 B.n24 10.6151
R980 B.n575 B.n24 10.6151
R981 B.n576 B.n575 10.6151
R982 B.n577 B.n576 10.6151
R983 B.n577 B.n22 10.6151
R984 B.n581 B.n22 10.6151
R985 B.n582 B.n581 10.6151
R986 B.n583 B.n582 10.6151
R987 B.n583 B.n20 10.6151
R988 B.n587 B.n20 10.6151
R989 B.n588 B.n587 10.6151
R990 B.n589 B.n588 10.6151
R991 B.n589 B.n18 10.6151
R992 B.n593 B.n18 10.6151
R993 B.n594 B.n593 10.6151
R994 B.n595 B.n594 10.6151
R995 B.n595 B.n16 10.6151
R996 B.n599 B.n16 10.6151
R997 B.n600 B.n599 10.6151
R998 B.n601 B.n600 10.6151
R999 B.n601 B.n14 10.6151
R1000 B.n605 B.n14 10.6151
R1001 B.n606 B.n605 10.6151
R1002 B.n607 B.n606 10.6151
R1003 B.n607 B.n12 10.6151
R1004 B.n611 B.n12 10.6151
R1005 B.n612 B.n611 10.6151
R1006 B.n613 B.n612 10.6151
R1007 B.n613 B.n10 10.6151
R1008 B.n617 B.n10 10.6151
R1009 B.n618 B.n617 10.6151
R1010 B.n619 B.n618 10.6151
R1011 B.n619 B.n8 10.6151
R1012 B.n623 B.n8 10.6151
R1013 B.n624 B.n623 10.6151
R1014 B.n625 B.n624 10.6151
R1015 B.n625 B.n6 10.6151
R1016 B.n629 B.n6 10.6151
R1017 B.n630 B.n629 10.6151
R1018 B.n631 B.n630 10.6151
R1019 B.n631 B.n4 10.6151
R1020 B.n635 B.n4 10.6151
R1021 B.n636 B.n635 10.6151
R1022 B.n637 B.n636 10.6151
R1023 B.n637 B.n0 10.6151
R1024 B.n541 B.n34 10.6151
R1025 B.n541 B.n540 10.6151
R1026 B.n540 B.n539 10.6151
R1027 B.n539 B.n36 10.6151
R1028 B.n535 B.n36 10.6151
R1029 B.n535 B.n534 10.6151
R1030 B.n534 B.n533 10.6151
R1031 B.n533 B.n38 10.6151
R1032 B.n529 B.n528 10.6151
R1033 B.n528 B.n527 10.6151
R1034 B.n527 B.n43 10.6151
R1035 B.n523 B.n43 10.6151
R1036 B.n523 B.n522 10.6151
R1037 B.n522 B.n521 10.6151
R1038 B.n521 B.n45 10.6151
R1039 B.n517 B.n45 10.6151
R1040 B.n517 B.n516 10.6151
R1041 B.n514 B.n49 10.6151
R1042 B.n510 B.n49 10.6151
R1043 B.n510 B.n509 10.6151
R1044 B.n509 B.n508 10.6151
R1045 B.n508 B.n51 10.6151
R1046 B.n504 B.n51 10.6151
R1047 B.n504 B.n503 10.6151
R1048 B.n503 B.n502 10.6151
R1049 B.n498 B.n53 10.6151
R1050 B.n498 B.n497 10.6151
R1051 B.n497 B.n496 10.6151
R1052 B.n496 B.n55 10.6151
R1053 B.n492 B.n55 10.6151
R1054 B.n492 B.n491 10.6151
R1055 B.n491 B.n490 10.6151
R1056 B.n490 B.n57 10.6151
R1057 B.n486 B.n57 10.6151
R1058 B.n486 B.n485 10.6151
R1059 B.n485 B.n484 10.6151
R1060 B.n484 B.n59 10.6151
R1061 B.n480 B.n59 10.6151
R1062 B.n480 B.n479 10.6151
R1063 B.n479 B.n478 10.6151
R1064 B.n478 B.n61 10.6151
R1065 B.n474 B.n61 10.6151
R1066 B.n474 B.n473 10.6151
R1067 B.n473 B.n472 10.6151
R1068 B.n472 B.n63 10.6151
R1069 B.n468 B.n63 10.6151
R1070 B.n468 B.n467 10.6151
R1071 B.n467 B.n466 10.6151
R1072 B.n466 B.n65 10.6151
R1073 B.n462 B.n65 10.6151
R1074 B.n462 B.n461 10.6151
R1075 B.n461 B.n460 10.6151
R1076 B.n460 B.n67 10.6151
R1077 B.n456 B.n67 10.6151
R1078 B.n456 B.n455 10.6151
R1079 B.n455 B.n454 10.6151
R1080 B.n454 B.n69 10.6151
R1081 B.n450 B.n69 10.6151
R1082 B.n450 B.n449 10.6151
R1083 B.n449 B.n448 10.6151
R1084 B.n448 B.n71 10.6151
R1085 B.n444 B.n71 10.6151
R1086 B.n444 B.n443 10.6151
R1087 B.n443 B.n442 10.6151
R1088 B.n442 B.n73 10.6151
R1089 B.n438 B.n73 10.6151
R1090 B.n438 B.n437 10.6151
R1091 B.n437 B.n436 10.6151
R1092 B.n436 B.n75 10.6151
R1093 B.n432 B.n75 10.6151
R1094 B.n432 B.n431 10.6151
R1095 B.n431 B.n430 10.6151
R1096 B.n430 B.n77 10.6151
R1097 B.n426 B.n77 10.6151
R1098 B.n426 B.n425 10.6151
R1099 B.n425 B.n424 10.6151
R1100 B.n424 B.n79 10.6151
R1101 B.n420 B.n79 10.6151
R1102 B.n420 B.n419 10.6151
R1103 B.n419 B.n418 10.6151
R1104 B.n418 B.n81 10.6151
R1105 B.n414 B.n81 10.6151
R1106 B.n414 B.n413 10.6151
R1107 B.n413 B.n412 10.6151
R1108 B.n412 B.n83 10.6151
R1109 B.n408 B.n83 10.6151
R1110 B.n408 B.n407 10.6151
R1111 B.n407 B.n406 10.6151
R1112 B.n406 B.n85 10.6151
R1113 B.n402 B.n85 10.6151
R1114 B.n402 B.n401 10.6151
R1115 B.n401 B.n400 10.6151
R1116 B.n400 B.n87 10.6151
R1117 B.n396 B.n87 10.6151
R1118 B.n396 B.n395 10.6151
R1119 B.n395 B.n394 10.6151
R1120 B.n394 B.n89 10.6151
R1121 B.n390 B.n89 10.6151
R1122 B.n390 B.n389 10.6151
R1123 B.n389 B.n388 10.6151
R1124 B.n388 B.n91 10.6151
R1125 B.n384 B.n91 10.6151
R1126 B.n384 B.n383 10.6151
R1127 B.n383 B.n382 10.6151
R1128 B.n382 B.n93 10.6151
R1129 B.n378 B.n93 10.6151
R1130 B.n378 B.n377 10.6151
R1131 B.n377 B.n376 10.6151
R1132 B.n376 B.n95 10.6151
R1133 B.n372 B.n95 10.6151
R1134 B.n372 B.n371 10.6151
R1135 B.n371 B.n370 10.6151
R1136 B.n370 B.n97 10.6151
R1137 B.n366 B.n97 10.6151
R1138 B.n366 B.n365 10.6151
R1139 B.n365 B.n364 10.6151
R1140 B.n364 B.n99 10.6151
R1141 B.n360 B.n99 10.6151
R1142 B.n360 B.n359 10.6151
R1143 B.n359 B.n358 10.6151
R1144 B.n358 B.n101 10.6151
R1145 B.n354 B.n101 10.6151
R1146 B.n354 B.n353 10.6151
R1147 B.n353 B.n352 10.6151
R1148 B.n352 B.n103 10.6151
R1149 B.n348 B.n103 10.6151
R1150 B.n348 B.n347 10.6151
R1151 B.n347 B.n346 10.6151
R1152 B.n346 B.n105 10.6151
R1153 B.n342 B.n105 10.6151
R1154 B.n342 B.n341 10.6151
R1155 B.n341 B.n340 10.6151
R1156 B.n340 B.n107 10.6151
R1157 B.n336 B.n107 10.6151
R1158 B.n336 B.n335 10.6151
R1159 B.n335 B.n334 10.6151
R1160 B.n334 B.n109 10.6151
R1161 B.n330 B.n109 10.6151
R1162 B.n330 B.n329 10.6151
R1163 B.n329 B.n328 10.6151
R1164 B.n328 B.n111 10.6151
R1165 B.n324 B.n111 10.6151
R1166 B.n324 B.n323 10.6151
R1167 B.n323 B.n322 10.6151
R1168 B.n322 B.n113 10.6151
R1169 B.n318 B.n113 10.6151
R1170 B.n318 B.n317 10.6151
R1171 B.n317 B.n316 10.6151
R1172 B.n316 B.n115 10.6151
R1173 B.n312 B.n115 10.6151
R1174 B.n312 B.n311 10.6151
R1175 B.n311 B.n310 10.6151
R1176 B.n310 B.n117 10.6151
R1177 B.n306 B.n117 10.6151
R1178 B.n165 B.n1 10.6151
R1179 B.n168 B.n165 10.6151
R1180 B.n169 B.n168 10.6151
R1181 B.n170 B.n169 10.6151
R1182 B.n170 B.n163 10.6151
R1183 B.n174 B.n163 10.6151
R1184 B.n175 B.n174 10.6151
R1185 B.n176 B.n175 10.6151
R1186 B.n176 B.n161 10.6151
R1187 B.n180 B.n161 10.6151
R1188 B.n181 B.n180 10.6151
R1189 B.n182 B.n181 10.6151
R1190 B.n182 B.n159 10.6151
R1191 B.n186 B.n159 10.6151
R1192 B.n187 B.n186 10.6151
R1193 B.n188 B.n187 10.6151
R1194 B.n188 B.n157 10.6151
R1195 B.n192 B.n157 10.6151
R1196 B.n193 B.n192 10.6151
R1197 B.n194 B.n193 10.6151
R1198 B.n194 B.n155 10.6151
R1199 B.n198 B.n155 10.6151
R1200 B.n199 B.n198 10.6151
R1201 B.n200 B.n199 10.6151
R1202 B.n200 B.n153 10.6151
R1203 B.n204 B.n153 10.6151
R1204 B.n205 B.n204 10.6151
R1205 B.n206 B.n205 10.6151
R1206 B.n206 B.n151 10.6151
R1207 B.n210 B.n151 10.6151
R1208 B.n211 B.n210 10.6151
R1209 B.n212 B.n211 10.6151
R1210 B.n212 B.n149 10.6151
R1211 B.n216 B.n149 10.6151
R1212 B.n217 B.n216 10.6151
R1213 B.n218 B.n217 10.6151
R1214 B.n218 B.n147 10.6151
R1215 B.n222 B.n147 10.6151
R1216 B.n223 B.n222 10.6151
R1217 B.n224 B.n223 10.6151
R1218 B.n224 B.n145 10.6151
R1219 B.n228 B.n145 10.6151
R1220 B.n229 B.n228 10.6151
R1221 B.n230 B.n229 10.6151
R1222 B.n230 B.n143 10.6151
R1223 B.n234 B.n143 10.6151
R1224 B.n235 B.n234 10.6151
R1225 B.n236 B.n235 10.6151
R1226 B.n236 B.n141 10.6151
R1227 B.n240 B.n141 10.6151
R1228 B.n241 B.n240 10.6151
R1229 B.n242 B.n241 10.6151
R1230 B.n242 B.n139 10.6151
R1231 B.n246 B.n139 10.6151
R1232 B.n247 B.n246 10.6151
R1233 B.n248 B.n247 10.6151
R1234 B.n248 B.n137 10.6151
R1235 B.n252 B.n137 10.6151
R1236 B.n253 B.n252 10.6151
R1237 B.n254 B.n253 10.6151
R1238 B.n254 B.n135 10.6151
R1239 B.n258 B.n135 10.6151
R1240 B.n259 B.n258 10.6151
R1241 B.n260 B.n133 10.6151
R1242 B.n264 B.n133 10.6151
R1243 B.n265 B.n264 10.6151
R1244 B.n266 B.n265 10.6151
R1245 B.n266 B.n131 10.6151
R1246 B.n270 B.n131 10.6151
R1247 B.n271 B.n270 10.6151
R1248 B.n275 B.n271 10.6151
R1249 B.n279 B.n129 10.6151
R1250 B.n280 B.n279 10.6151
R1251 B.n281 B.n280 10.6151
R1252 B.n281 B.n127 10.6151
R1253 B.n285 B.n127 10.6151
R1254 B.n286 B.n285 10.6151
R1255 B.n287 B.n286 10.6151
R1256 B.n287 B.n125 10.6151
R1257 B.n291 B.n125 10.6151
R1258 B.n294 B.n293 10.6151
R1259 B.n294 B.n121 10.6151
R1260 B.n298 B.n121 10.6151
R1261 B.n299 B.n298 10.6151
R1262 B.n300 B.n299 10.6151
R1263 B.n300 B.n119 10.6151
R1264 B.n304 B.n119 10.6151
R1265 B.n305 B.n304 10.6151
R1266 B.n42 B.n38 9.36635
R1267 B.n515 B.n514 9.36635
R1268 B.n275 B.n274 9.36635
R1269 B.n293 B.n292 9.36635
R1270 B.n641 B.n0 8.11757
R1271 B.n641 B.n1 8.11757
R1272 B.n529 B.n42 1.24928
R1273 B.n516 B.n515 1.24928
R1274 B.n274 B.n129 1.24928
R1275 B.n292 B.n291 1.24928
C0 VDD2 w_n4790_n1174# 2.09194f
C1 VDD2 VN 1.22355f
C2 VDD1 B 1.6254f
C3 VTAIL VDD1 5.25178f
C4 VDD1 VP 1.68215f
C5 VTAIL B 1.39167f
C6 B VP 2.3166f
C7 VDD1 w_n4790_n1174# 1.94096f
C8 VTAIL VP 2.94417f
C9 VDD1 VN 0.160544f
C10 w_n4790_n1174# B 8.525041f
C11 B VN 1.26626f
C12 VTAIL w_n4790_n1174# 1.8057f
C13 VTAIL VN 2.93007f
C14 w_n4790_n1174# VP 10.462299f
C15 VDD2 VDD1 2.23955f
C16 VN VP 6.72904f
C17 VDD2 B 1.7502f
C18 VDD2 VTAIL 5.31216f
C19 w_n4790_n1174# VN 9.84544f
C20 VDD2 VP 0.623766f
C21 VDD2 VSUBS 1.872669f
C22 VDD1 VSUBS 2.393644f
C23 VTAIL VSUBS 0.644828f
C24 VN VSUBS 8.467221f
C25 VP VSUBS 3.82728f
C26 B VSUBS 4.750171f
C27 w_n4790_n1174# VSUBS 72.4823f
C28 B.n0 VSUBS 0.011076f
C29 B.n1 VSUBS 0.011076f
C30 B.n2 VSUBS 0.016381f
C31 B.n3 VSUBS 0.012553f
C32 B.n4 VSUBS 0.012553f
C33 B.n5 VSUBS 0.012553f
C34 B.n6 VSUBS 0.012553f
C35 B.n7 VSUBS 0.012553f
C36 B.n8 VSUBS 0.012553f
C37 B.n9 VSUBS 0.012553f
C38 B.n10 VSUBS 0.012553f
C39 B.n11 VSUBS 0.012553f
C40 B.n12 VSUBS 0.012553f
C41 B.n13 VSUBS 0.012553f
C42 B.n14 VSUBS 0.012553f
C43 B.n15 VSUBS 0.012553f
C44 B.n16 VSUBS 0.012553f
C45 B.n17 VSUBS 0.012553f
C46 B.n18 VSUBS 0.012553f
C47 B.n19 VSUBS 0.012553f
C48 B.n20 VSUBS 0.012553f
C49 B.n21 VSUBS 0.012553f
C50 B.n22 VSUBS 0.012553f
C51 B.n23 VSUBS 0.012553f
C52 B.n24 VSUBS 0.012553f
C53 B.n25 VSUBS 0.012553f
C54 B.n26 VSUBS 0.012553f
C55 B.n27 VSUBS 0.012553f
C56 B.n28 VSUBS 0.012553f
C57 B.n29 VSUBS 0.012553f
C58 B.n30 VSUBS 0.012553f
C59 B.n31 VSUBS 0.012553f
C60 B.n32 VSUBS 0.012553f
C61 B.n33 VSUBS 0.012553f
C62 B.n34 VSUBS 0.029078f
C63 B.n35 VSUBS 0.012553f
C64 B.n36 VSUBS 0.012553f
C65 B.n37 VSUBS 0.012553f
C66 B.n38 VSUBS 0.011815f
C67 B.n39 VSUBS 0.012553f
C68 B.t4 VSUBS 0.034728f
C69 B.t5 VSUBS 0.047096f
C70 B.t3 VSUBS 0.324415f
C71 B.n40 VSUBS 0.126259f
C72 B.n41 VSUBS 0.090672f
C73 B.n42 VSUBS 0.029084f
C74 B.n43 VSUBS 0.012553f
C75 B.n44 VSUBS 0.012553f
C76 B.n45 VSUBS 0.012553f
C77 B.n46 VSUBS 0.012553f
C78 B.t1 VSUBS 0.034728f
C79 B.t2 VSUBS 0.047096f
C80 B.t0 VSUBS 0.324415f
C81 B.n47 VSUBS 0.126259f
C82 B.n48 VSUBS 0.090672f
C83 B.n49 VSUBS 0.012553f
C84 B.n50 VSUBS 0.012553f
C85 B.n51 VSUBS 0.012553f
C86 B.n52 VSUBS 0.012553f
C87 B.n53 VSUBS 0.028519f
C88 B.n54 VSUBS 0.012553f
C89 B.n55 VSUBS 0.012553f
C90 B.n56 VSUBS 0.012553f
C91 B.n57 VSUBS 0.012553f
C92 B.n58 VSUBS 0.012553f
C93 B.n59 VSUBS 0.012553f
C94 B.n60 VSUBS 0.012553f
C95 B.n61 VSUBS 0.012553f
C96 B.n62 VSUBS 0.012553f
C97 B.n63 VSUBS 0.012553f
C98 B.n64 VSUBS 0.012553f
C99 B.n65 VSUBS 0.012553f
C100 B.n66 VSUBS 0.012553f
C101 B.n67 VSUBS 0.012553f
C102 B.n68 VSUBS 0.012553f
C103 B.n69 VSUBS 0.012553f
C104 B.n70 VSUBS 0.012553f
C105 B.n71 VSUBS 0.012553f
C106 B.n72 VSUBS 0.012553f
C107 B.n73 VSUBS 0.012553f
C108 B.n74 VSUBS 0.012553f
C109 B.n75 VSUBS 0.012553f
C110 B.n76 VSUBS 0.012553f
C111 B.n77 VSUBS 0.012553f
C112 B.n78 VSUBS 0.012553f
C113 B.n79 VSUBS 0.012553f
C114 B.n80 VSUBS 0.012553f
C115 B.n81 VSUBS 0.012553f
C116 B.n82 VSUBS 0.012553f
C117 B.n83 VSUBS 0.012553f
C118 B.n84 VSUBS 0.012553f
C119 B.n85 VSUBS 0.012553f
C120 B.n86 VSUBS 0.012553f
C121 B.n87 VSUBS 0.012553f
C122 B.n88 VSUBS 0.012553f
C123 B.n89 VSUBS 0.012553f
C124 B.n90 VSUBS 0.012553f
C125 B.n91 VSUBS 0.012553f
C126 B.n92 VSUBS 0.012553f
C127 B.n93 VSUBS 0.012553f
C128 B.n94 VSUBS 0.012553f
C129 B.n95 VSUBS 0.012553f
C130 B.n96 VSUBS 0.012553f
C131 B.n97 VSUBS 0.012553f
C132 B.n98 VSUBS 0.012553f
C133 B.n99 VSUBS 0.012553f
C134 B.n100 VSUBS 0.012553f
C135 B.n101 VSUBS 0.012553f
C136 B.n102 VSUBS 0.012553f
C137 B.n103 VSUBS 0.012553f
C138 B.n104 VSUBS 0.012553f
C139 B.n105 VSUBS 0.012553f
C140 B.n106 VSUBS 0.012553f
C141 B.n107 VSUBS 0.012553f
C142 B.n108 VSUBS 0.012553f
C143 B.n109 VSUBS 0.012553f
C144 B.n110 VSUBS 0.012553f
C145 B.n111 VSUBS 0.012553f
C146 B.n112 VSUBS 0.012553f
C147 B.n113 VSUBS 0.012553f
C148 B.n114 VSUBS 0.012553f
C149 B.n115 VSUBS 0.012553f
C150 B.n116 VSUBS 0.012553f
C151 B.n117 VSUBS 0.012553f
C152 B.n118 VSUBS 0.029078f
C153 B.n119 VSUBS 0.012553f
C154 B.n120 VSUBS 0.012553f
C155 B.n121 VSUBS 0.012553f
C156 B.n122 VSUBS 0.012553f
C157 B.t11 VSUBS 0.034728f
C158 B.t10 VSUBS 0.047096f
C159 B.t9 VSUBS 0.324415f
C160 B.n123 VSUBS 0.126259f
C161 B.n124 VSUBS 0.090672f
C162 B.n125 VSUBS 0.012553f
C163 B.n126 VSUBS 0.012553f
C164 B.n127 VSUBS 0.012553f
C165 B.n128 VSUBS 0.012553f
C166 B.n129 VSUBS 0.007015f
C167 B.n130 VSUBS 0.012553f
C168 B.n131 VSUBS 0.012553f
C169 B.n132 VSUBS 0.012553f
C170 B.n133 VSUBS 0.012553f
C171 B.n134 VSUBS 0.028519f
C172 B.n135 VSUBS 0.012553f
C173 B.n136 VSUBS 0.012553f
C174 B.n137 VSUBS 0.012553f
C175 B.n138 VSUBS 0.012553f
C176 B.n139 VSUBS 0.012553f
C177 B.n140 VSUBS 0.012553f
C178 B.n141 VSUBS 0.012553f
C179 B.n142 VSUBS 0.012553f
C180 B.n143 VSUBS 0.012553f
C181 B.n144 VSUBS 0.012553f
C182 B.n145 VSUBS 0.012553f
C183 B.n146 VSUBS 0.012553f
C184 B.n147 VSUBS 0.012553f
C185 B.n148 VSUBS 0.012553f
C186 B.n149 VSUBS 0.012553f
C187 B.n150 VSUBS 0.012553f
C188 B.n151 VSUBS 0.012553f
C189 B.n152 VSUBS 0.012553f
C190 B.n153 VSUBS 0.012553f
C191 B.n154 VSUBS 0.012553f
C192 B.n155 VSUBS 0.012553f
C193 B.n156 VSUBS 0.012553f
C194 B.n157 VSUBS 0.012553f
C195 B.n158 VSUBS 0.012553f
C196 B.n159 VSUBS 0.012553f
C197 B.n160 VSUBS 0.012553f
C198 B.n161 VSUBS 0.012553f
C199 B.n162 VSUBS 0.012553f
C200 B.n163 VSUBS 0.012553f
C201 B.n164 VSUBS 0.012553f
C202 B.n165 VSUBS 0.012553f
C203 B.n166 VSUBS 0.012553f
C204 B.n167 VSUBS 0.012553f
C205 B.n168 VSUBS 0.012553f
C206 B.n169 VSUBS 0.012553f
C207 B.n170 VSUBS 0.012553f
C208 B.n171 VSUBS 0.012553f
C209 B.n172 VSUBS 0.012553f
C210 B.n173 VSUBS 0.012553f
C211 B.n174 VSUBS 0.012553f
C212 B.n175 VSUBS 0.012553f
C213 B.n176 VSUBS 0.012553f
C214 B.n177 VSUBS 0.012553f
C215 B.n178 VSUBS 0.012553f
C216 B.n179 VSUBS 0.012553f
C217 B.n180 VSUBS 0.012553f
C218 B.n181 VSUBS 0.012553f
C219 B.n182 VSUBS 0.012553f
C220 B.n183 VSUBS 0.012553f
C221 B.n184 VSUBS 0.012553f
C222 B.n185 VSUBS 0.012553f
C223 B.n186 VSUBS 0.012553f
C224 B.n187 VSUBS 0.012553f
C225 B.n188 VSUBS 0.012553f
C226 B.n189 VSUBS 0.012553f
C227 B.n190 VSUBS 0.012553f
C228 B.n191 VSUBS 0.012553f
C229 B.n192 VSUBS 0.012553f
C230 B.n193 VSUBS 0.012553f
C231 B.n194 VSUBS 0.012553f
C232 B.n195 VSUBS 0.012553f
C233 B.n196 VSUBS 0.012553f
C234 B.n197 VSUBS 0.012553f
C235 B.n198 VSUBS 0.012553f
C236 B.n199 VSUBS 0.012553f
C237 B.n200 VSUBS 0.012553f
C238 B.n201 VSUBS 0.012553f
C239 B.n202 VSUBS 0.012553f
C240 B.n203 VSUBS 0.012553f
C241 B.n204 VSUBS 0.012553f
C242 B.n205 VSUBS 0.012553f
C243 B.n206 VSUBS 0.012553f
C244 B.n207 VSUBS 0.012553f
C245 B.n208 VSUBS 0.012553f
C246 B.n209 VSUBS 0.012553f
C247 B.n210 VSUBS 0.012553f
C248 B.n211 VSUBS 0.012553f
C249 B.n212 VSUBS 0.012553f
C250 B.n213 VSUBS 0.012553f
C251 B.n214 VSUBS 0.012553f
C252 B.n215 VSUBS 0.012553f
C253 B.n216 VSUBS 0.012553f
C254 B.n217 VSUBS 0.012553f
C255 B.n218 VSUBS 0.012553f
C256 B.n219 VSUBS 0.012553f
C257 B.n220 VSUBS 0.012553f
C258 B.n221 VSUBS 0.012553f
C259 B.n222 VSUBS 0.012553f
C260 B.n223 VSUBS 0.012553f
C261 B.n224 VSUBS 0.012553f
C262 B.n225 VSUBS 0.012553f
C263 B.n226 VSUBS 0.012553f
C264 B.n227 VSUBS 0.012553f
C265 B.n228 VSUBS 0.012553f
C266 B.n229 VSUBS 0.012553f
C267 B.n230 VSUBS 0.012553f
C268 B.n231 VSUBS 0.012553f
C269 B.n232 VSUBS 0.012553f
C270 B.n233 VSUBS 0.012553f
C271 B.n234 VSUBS 0.012553f
C272 B.n235 VSUBS 0.012553f
C273 B.n236 VSUBS 0.012553f
C274 B.n237 VSUBS 0.012553f
C275 B.n238 VSUBS 0.012553f
C276 B.n239 VSUBS 0.012553f
C277 B.n240 VSUBS 0.012553f
C278 B.n241 VSUBS 0.012553f
C279 B.n242 VSUBS 0.012553f
C280 B.n243 VSUBS 0.012553f
C281 B.n244 VSUBS 0.012553f
C282 B.n245 VSUBS 0.012553f
C283 B.n246 VSUBS 0.012553f
C284 B.n247 VSUBS 0.012553f
C285 B.n248 VSUBS 0.012553f
C286 B.n249 VSUBS 0.012553f
C287 B.n250 VSUBS 0.012553f
C288 B.n251 VSUBS 0.012553f
C289 B.n252 VSUBS 0.012553f
C290 B.n253 VSUBS 0.012553f
C291 B.n254 VSUBS 0.012553f
C292 B.n255 VSUBS 0.012553f
C293 B.n256 VSUBS 0.012553f
C294 B.n257 VSUBS 0.012553f
C295 B.n258 VSUBS 0.012553f
C296 B.n259 VSUBS 0.028519f
C297 B.n260 VSUBS 0.029078f
C298 B.n261 VSUBS 0.029078f
C299 B.n262 VSUBS 0.012553f
C300 B.n263 VSUBS 0.012553f
C301 B.n264 VSUBS 0.012553f
C302 B.n265 VSUBS 0.012553f
C303 B.n266 VSUBS 0.012553f
C304 B.n267 VSUBS 0.012553f
C305 B.n268 VSUBS 0.012553f
C306 B.n269 VSUBS 0.012553f
C307 B.n270 VSUBS 0.012553f
C308 B.n271 VSUBS 0.012553f
C309 B.t8 VSUBS 0.034728f
C310 B.t7 VSUBS 0.047096f
C311 B.t6 VSUBS 0.324415f
C312 B.n272 VSUBS 0.126259f
C313 B.n273 VSUBS 0.090672f
C314 B.n274 VSUBS 0.029084f
C315 B.n275 VSUBS 0.011815f
C316 B.n276 VSUBS 0.012553f
C317 B.n277 VSUBS 0.012553f
C318 B.n278 VSUBS 0.012553f
C319 B.n279 VSUBS 0.012553f
C320 B.n280 VSUBS 0.012553f
C321 B.n281 VSUBS 0.012553f
C322 B.n282 VSUBS 0.012553f
C323 B.n283 VSUBS 0.012553f
C324 B.n284 VSUBS 0.012553f
C325 B.n285 VSUBS 0.012553f
C326 B.n286 VSUBS 0.012553f
C327 B.n287 VSUBS 0.012553f
C328 B.n288 VSUBS 0.012553f
C329 B.n289 VSUBS 0.012553f
C330 B.n290 VSUBS 0.012553f
C331 B.n291 VSUBS 0.007015f
C332 B.n292 VSUBS 0.029084f
C333 B.n293 VSUBS 0.011815f
C334 B.n294 VSUBS 0.012553f
C335 B.n295 VSUBS 0.012553f
C336 B.n296 VSUBS 0.012553f
C337 B.n297 VSUBS 0.012553f
C338 B.n298 VSUBS 0.012553f
C339 B.n299 VSUBS 0.012553f
C340 B.n300 VSUBS 0.012553f
C341 B.n301 VSUBS 0.012553f
C342 B.n302 VSUBS 0.012553f
C343 B.n303 VSUBS 0.012553f
C344 B.n304 VSUBS 0.012553f
C345 B.n305 VSUBS 0.02755f
C346 B.n306 VSUBS 0.030048f
C347 B.n307 VSUBS 0.028519f
C348 B.n308 VSUBS 0.012553f
C349 B.n309 VSUBS 0.012553f
C350 B.n310 VSUBS 0.012553f
C351 B.n311 VSUBS 0.012553f
C352 B.n312 VSUBS 0.012553f
C353 B.n313 VSUBS 0.012553f
C354 B.n314 VSUBS 0.012553f
C355 B.n315 VSUBS 0.012553f
C356 B.n316 VSUBS 0.012553f
C357 B.n317 VSUBS 0.012553f
C358 B.n318 VSUBS 0.012553f
C359 B.n319 VSUBS 0.012553f
C360 B.n320 VSUBS 0.012553f
C361 B.n321 VSUBS 0.012553f
C362 B.n322 VSUBS 0.012553f
C363 B.n323 VSUBS 0.012553f
C364 B.n324 VSUBS 0.012553f
C365 B.n325 VSUBS 0.012553f
C366 B.n326 VSUBS 0.012553f
C367 B.n327 VSUBS 0.012553f
C368 B.n328 VSUBS 0.012553f
C369 B.n329 VSUBS 0.012553f
C370 B.n330 VSUBS 0.012553f
C371 B.n331 VSUBS 0.012553f
C372 B.n332 VSUBS 0.012553f
C373 B.n333 VSUBS 0.012553f
C374 B.n334 VSUBS 0.012553f
C375 B.n335 VSUBS 0.012553f
C376 B.n336 VSUBS 0.012553f
C377 B.n337 VSUBS 0.012553f
C378 B.n338 VSUBS 0.012553f
C379 B.n339 VSUBS 0.012553f
C380 B.n340 VSUBS 0.012553f
C381 B.n341 VSUBS 0.012553f
C382 B.n342 VSUBS 0.012553f
C383 B.n343 VSUBS 0.012553f
C384 B.n344 VSUBS 0.012553f
C385 B.n345 VSUBS 0.012553f
C386 B.n346 VSUBS 0.012553f
C387 B.n347 VSUBS 0.012553f
C388 B.n348 VSUBS 0.012553f
C389 B.n349 VSUBS 0.012553f
C390 B.n350 VSUBS 0.012553f
C391 B.n351 VSUBS 0.012553f
C392 B.n352 VSUBS 0.012553f
C393 B.n353 VSUBS 0.012553f
C394 B.n354 VSUBS 0.012553f
C395 B.n355 VSUBS 0.012553f
C396 B.n356 VSUBS 0.012553f
C397 B.n357 VSUBS 0.012553f
C398 B.n358 VSUBS 0.012553f
C399 B.n359 VSUBS 0.012553f
C400 B.n360 VSUBS 0.012553f
C401 B.n361 VSUBS 0.012553f
C402 B.n362 VSUBS 0.012553f
C403 B.n363 VSUBS 0.012553f
C404 B.n364 VSUBS 0.012553f
C405 B.n365 VSUBS 0.012553f
C406 B.n366 VSUBS 0.012553f
C407 B.n367 VSUBS 0.012553f
C408 B.n368 VSUBS 0.012553f
C409 B.n369 VSUBS 0.012553f
C410 B.n370 VSUBS 0.012553f
C411 B.n371 VSUBS 0.012553f
C412 B.n372 VSUBS 0.012553f
C413 B.n373 VSUBS 0.012553f
C414 B.n374 VSUBS 0.012553f
C415 B.n375 VSUBS 0.012553f
C416 B.n376 VSUBS 0.012553f
C417 B.n377 VSUBS 0.012553f
C418 B.n378 VSUBS 0.012553f
C419 B.n379 VSUBS 0.012553f
C420 B.n380 VSUBS 0.012553f
C421 B.n381 VSUBS 0.012553f
C422 B.n382 VSUBS 0.012553f
C423 B.n383 VSUBS 0.012553f
C424 B.n384 VSUBS 0.012553f
C425 B.n385 VSUBS 0.012553f
C426 B.n386 VSUBS 0.012553f
C427 B.n387 VSUBS 0.012553f
C428 B.n388 VSUBS 0.012553f
C429 B.n389 VSUBS 0.012553f
C430 B.n390 VSUBS 0.012553f
C431 B.n391 VSUBS 0.012553f
C432 B.n392 VSUBS 0.012553f
C433 B.n393 VSUBS 0.012553f
C434 B.n394 VSUBS 0.012553f
C435 B.n395 VSUBS 0.012553f
C436 B.n396 VSUBS 0.012553f
C437 B.n397 VSUBS 0.012553f
C438 B.n398 VSUBS 0.012553f
C439 B.n399 VSUBS 0.012553f
C440 B.n400 VSUBS 0.012553f
C441 B.n401 VSUBS 0.012553f
C442 B.n402 VSUBS 0.012553f
C443 B.n403 VSUBS 0.012553f
C444 B.n404 VSUBS 0.012553f
C445 B.n405 VSUBS 0.012553f
C446 B.n406 VSUBS 0.012553f
C447 B.n407 VSUBS 0.012553f
C448 B.n408 VSUBS 0.012553f
C449 B.n409 VSUBS 0.012553f
C450 B.n410 VSUBS 0.012553f
C451 B.n411 VSUBS 0.012553f
C452 B.n412 VSUBS 0.012553f
C453 B.n413 VSUBS 0.012553f
C454 B.n414 VSUBS 0.012553f
C455 B.n415 VSUBS 0.012553f
C456 B.n416 VSUBS 0.012553f
C457 B.n417 VSUBS 0.012553f
C458 B.n418 VSUBS 0.012553f
C459 B.n419 VSUBS 0.012553f
C460 B.n420 VSUBS 0.012553f
C461 B.n421 VSUBS 0.012553f
C462 B.n422 VSUBS 0.012553f
C463 B.n423 VSUBS 0.012553f
C464 B.n424 VSUBS 0.012553f
C465 B.n425 VSUBS 0.012553f
C466 B.n426 VSUBS 0.012553f
C467 B.n427 VSUBS 0.012553f
C468 B.n428 VSUBS 0.012553f
C469 B.n429 VSUBS 0.012553f
C470 B.n430 VSUBS 0.012553f
C471 B.n431 VSUBS 0.012553f
C472 B.n432 VSUBS 0.012553f
C473 B.n433 VSUBS 0.012553f
C474 B.n434 VSUBS 0.012553f
C475 B.n435 VSUBS 0.012553f
C476 B.n436 VSUBS 0.012553f
C477 B.n437 VSUBS 0.012553f
C478 B.n438 VSUBS 0.012553f
C479 B.n439 VSUBS 0.012553f
C480 B.n440 VSUBS 0.012553f
C481 B.n441 VSUBS 0.012553f
C482 B.n442 VSUBS 0.012553f
C483 B.n443 VSUBS 0.012553f
C484 B.n444 VSUBS 0.012553f
C485 B.n445 VSUBS 0.012553f
C486 B.n446 VSUBS 0.012553f
C487 B.n447 VSUBS 0.012553f
C488 B.n448 VSUBS 0.012553f
C489 B.n449 VSUBS 0.012553f
C490 B.n450 VSUBS 0.012553f
C491 B.n451 VSUBS 0.012553f
C492 B.n452 VSUBS 0.012553f
C493 B.n453 VSUBS 0.012553f
C494 B.n454 VSUBS 0.012553f
C495 B.n455 VSUBS 0.012553f
C496 B.n456 VSUBS 0.012553f
C497 B.n457 VSUBS 0.012553f
C498 B.n458 VSUBS 0.012553f
C499 B.n459 VSUBS 0.012553f
C500 B.n460 VSUBS 0.012553f
C501 B.n461 VSUBS 0.012553f
C502 B.n462 VSUBS 0.012553f
C503 B.n463 VSUBS 0.012553f
C504 B.n464 VSUBS 0.012553f
C505 B.n465 VSUBS 0.012553f
C506 B.n466 VSUBS 0.012553f
C507 B.n467 VSUBS 0.012553f
C508 B.n468 VSUBS 0.012553f
C509 B.n469 VSUBS 0.012553f
C510 B.n470 VSUBS 0.012553f
C511 B.n471 VSUBS 0.012553f
C512 B.n472 VSUBS 0.012553f
C513 B.n473 VSUBS 0.012553f
C514 B.n474 VSUBS 0.012553f
C515 B.n475 VSUBS 0.012553f
C516 B.n476 VSUBS 0.012553f
C517 B.n477 VSUBS 0.012553f
C518 B.n478 VSUBS 0.012553f
C519 B.n479 VSUBS 0.012553f
C520 B.n480 VSUBS 0.012553f
C521 B.n481 VSUBS 0.012553f
C522 B.n482 VSUBS 0.012553f
C523 B.n483 VSUBS 0.012553f
C524 B.n484 VSUBS 0.012553f
C525 B.n485 VSUBS 0.012553f
C526 B.n486 VSUBS 0.012553f
C527 B.n487 VSUBS 0.012553f
C528 B.n488 VSUBS 0.012553f
C529 B.n489 VSUBS 0.012553f
C530 B.n490 VSUBS 0.012553f
C531 B.n491 VSUBS 0.012553f
C532 B.n492 VSUBS 0.012553f
C533 B.n493 VSUBS 0.012553f
C534 B.n494 VSUBS 0.012553f
C535 B.n495 VSUBS 0.012553f
C536 B.n496 VSUBS 0.012553f
C537 B.n497 VSUBS 0.012553f
C538 B.n498 VSUBS 0.012553f
C539 B.n499 VSUBS 0.012553f
C540 B.n500 VSUBS 0.028519f
C541 B.n501 VSUBS 0.029078f
C542 B.n502 VSUBS 0.029078f
C543 B.n503 VSUBS 0.012553f
C544 B.n504 VSUBS 0.012553f
C545 B.n505 VSUBS 0.012553f
C546 B.n506 VSUBS 0.012553f
C547 B.n507 VSUBS 0.012553f
C548 B.n508 VSUBS 0.012553f
C549 B.n509 VSUBS 0.012553f
C550 B.n510 VSUBS 0.012553f
C551 B.n511 VSUBS 0.012553f
C552 B.n512 VSUBS 0.012553f
C553 B.n513 VSUBS 0.012553f
C554 B.n514 VSUBS 0.011815f
C555 B.n515 VSUBS 0.029084f
C556 B.n516 VSUBS 0.007015f
C557 B.n517 VSUBS 0.012553f
C558 B.n518 VSUBS 0.012553f
C559 B.n519 VSUBS 0.012553f
C560 B.n520 VSUBS 0.012553f
C561 B.n521 VSUBS 0.012553f
C562 B.n522 VSUBS 0.012553f
C563 B.n523 VSUBS 0.012553f
C564 B.n524 VSUBS 0.012553f
C565 B.n525 VSUBS 0.012553f
C566 B.n526 VSUBS 0.012553f
C567 B.n527 VSUBS 0.012553f
C568 B.n528 VSUBS 0.012553f
C569 B.n529 VSUBS 0.007015f
C570 B.n530 VSUBS 0.012553f
C571 B.n531 VSUBS 0.012553f
C572 B.n532 VSUBS 0.012553f
C573 B.n533 VSUBS 0.012553f
C574 B.n534 VSUBS 0.012553f
C575 B.n535 VSUBS 0.012553f
C576 B.n536 VSUBS 0.012553f
C577 B.n537 VSUBS 0.012553f
C578 B.n538 VSUBS 0.012553f
C579 B.n539 VSUBS 0.012553f
C580 B.n540 VSUBS 0.012553f
C581 B.n541 VSUBS 0.012553f
C582 B.n542 VSUBS 0.012553f
C583 B.n543 VSUBS 0.029078f
C584 B.n544 VSUBS 0.028519f
C585 B.n545 VSUBS 0.028519f
C586 B.n546 VSUBS 0.012553f
C587 B.n547 VSUBS 0.012553f
C588 B.n548 VSUBS 0.012553f
C589 B.n549 VSUBS 0.012553f
C590 B.n550 VSUBS 0.012553f
C591 B.n551 VSUBS 0.012553f
C592 B.n552 VSUBS 0.012553f
C593 B.n553 VSUBS 0.012553f
C594 B.n554 VSUBS 0.012553f
C595 B.n555 VSUBS 0.012553f
C596 B.n556 VSUBS 0.012553f
C597 B.n557 VSUBS 0.012553f
C598 B.n558 VSUBS 0.012553f
C599 B.n559 VSUBS 0.012553f
C600 B.n560 VSUBS 0.012553f
C601 B.n561 VSUBS 0.012553f
C602 B.n562 VSUBS 0.012553f
C603 B.n563 VSUBS 0.012553f
C604 B.n564 VSUBS 0.012553f
C605 B.n565 VSUBS 0.012553f
C606 B.n566 VSUBS 0.012553f
C607 B.n567 VSUBS 0.012553f
C608 B.n568 VSUBS 0.012553f
C609 B.n569 VSUBS 0.012553f
C610 B.n570 VSUBS 0.012553f
C611 B.n571 VSUBS 0.012553f
C612 B.n572 VSUBS 0.012553f
C613 B.n573 VSUBS 0.012553f
C614 B.n574 VSUBS 0.012553f
C615 B.n575 VSUBS 0.012553f
C616 B.n576 VSUBS 0.012553f
C617 B.n577 VSUBS 0.012553f
C618 B.n578 VSUBS 0.012553f
C619 B.n579 VSUBS 0.012553f
C620 B.n580 VSUBS 0.012553f
C621 B.n581 VSUBS 0.012553f
C622 B.n582 VSUBS 0.012553f
C623 B.n583 VSUBS 0.012553f
C624 B.n584 VSUBS 0.012553f
C625 B.n585 VSUBS 0.012553f
C626 B.n586 VSUBS 0.012553f
C627 B.n587 VSUBS 0.012553f
C628 B.n588 VSUBS 0.012553f
C629 B.n589 VSUBS 0.012553f
C630 B.n590 VSUBS 0.012553f
C631 B.n591 VSUBS 0.012553f
C632 B.n592 VSUBS 0.012553f
C633 B.n593 VSUBS 0.012553f
C634 B.n594 VSUBS 0.012553f
C635 B.n595 VSUBS 0.012553f
C636 B.n596 VSUBS 0.012553f
C637 B.n597 VSUBS 0.012553f
C638 B.n598 VSUBS 0.012553f
C639 B.n599 VSUBS 0.012553f
C640 B.n600 VSUBS 0.012553f
C641 B.n601 VSUBS 0.012553f
C642 B.n602 VSUBS 0.012553f
C643 B.n603 VSUBS 0.012553f
C644 B.n604 VSUBS 0.012553f
C645 B.n605 VSUBS 0.012553f
C646 B.n606 VSUBS 0.012553f
C647 B.n607 VSUBS 0.012553f
C648 B.n608 VSUBS 0.012553f
C649 B.n609 VSUBS 0.012553f
C650 B.n610 VSUBS 0.012553f
C651 B.n611 VSUBS 0.012553f
C652 B.n612 VSUBS 0.012553f
C653 B.n613 VSUBS 0.012553f
C654 B.n614 VSUBS 0.012553f
C655 B.n615 VSUBS 0.012553f
C656 B.n616 VSUBS 0.012553f
C657 B.n617 VSUBS 0.012553f
C658 B.n618 VSUBS 0.012553f
C659 B.n619 VSUBS 0.012553f
C660 B.n620 VSUBS 0.012553f
C661 B.n621 VSUBS 0.012553f
C662 B.n622 VSUBS 0.012553f
C663 B.n623 VSUBS 0.012553f
C664 B.n624 VSUBS 0.012553f
C665 B.n625 VSUBS 0.012553f
C666 B.n626 VSUBS 0.012553f
C667 B.n627 VSUBS 0.012553f
C668 B.n628 VSUBS 0.012553f
C669 B.n629 VSUBS 0.012553f
C670 B.n630 VSUBS 0.012553f
C671 B.n631 VSUBS 0.012553f
C672 B.n632 VSUBS 0.012553f
C673 B.n633 VSUBS 0.012553f
C674 B.n634 VSUBS 0.012553f
C675 B.n635 VSUBS 0.012553f
C676 B.n636 VSUBS 0.012553f
C677 B.n637 VSUBS 0.012553f
C678 B.n638 VSUBS 0.012553f
C679 B.n639 VSUBS 0.016381f
C680 B.n640 VSUBS 0.01745f
C681 B.n641 VSUBS 0.034702f
C682 VDD2.t6 VSUBS 0.028722f
C683 VDD2.t2 VSUBS 0.028722f
C684 VDD2.n0 VSUBS 0.098958f
C685 VDD2.t3 VSUBS 0.028722f
C686 VDD2.t5 VSUBS 0.028722f
C687 VDD2.n1 VSUBS 0.098958f
C688 VDD2.n2 VSUBS 4.39153f
C689 VDD2.t7 VSUBS 0.028722f
C690 VDD2.t0 VSUBS 0.028722f
C691 VDD2.n3 VSUBS 0.095109f
C692 VDD2.n4 VSUBS 3.37888f
C693 VDD2.t1 VSUBS 0.028722f
C694 VDD2.t4 VSUBS 0.028722f
C695 VDD2.n5 VSUBS 0.098948f
C696 VN.t2 VSUBS 0.38459f
C697 VN.n0 VSUBS 0.462913f
C698 VN.n1 VSUBS 0.056443f
C699 VN.n2 VSUBS 0.071386f
C700 VN.n3 VSUBS 0.056443f
C701 VN.n4 VSUBS 0.062608f
C702 VN.n5 VSUBS 0.056443f
C703 VN.n6 VSUBS 0.045629f
C704 VN.n7 VSUBS 0.056443f
C705 VN.t5 VSUBS 0.38459f
C706 VN.n8 VSUBS 0.454085f
C707 VN.t1 VSUBS 0.93381f
C708 VN.n9 VSUBS 0.540872f
C709 VN.n10 VSUBS 0.695501f
C710 VN.n11 VSUBS 0.095846f
C711 VN.n12 VSUBS 0.105195f
C712 VN.n13 VSUBS 0.112179f
C713 VN.n14 VSUBS 0.056443f
C714 VN.n15 VSUBS 0.056443f
C715 VN.n16 VSUBS 0.056443f
C716 VN.n17 VSUBS 0.112179f
C717 VN.n18 VSUBS 0.105195f
C718 VN.t4 VSUBS 0.38459f
C719 VN.n19 VSUBS 0.24147f
C720 VN.n20 VSUBS 0.095846f
C721 VN.n21 VSUBS 0.056443f
C722 VN.n22 VSUBS 0.056443f
C723 VN.n23 VSUBS 0.056443f
C724 VN.n24 VSUBS 0.105195f
C725 VN.n25 VSUBS 0.105195f
C726 VN.n26 VSUBS 0.093406f
C727 VN.n27 VSUBS 0.056443f
C728 VN.n28 VSUBS 0.056443f
C729 VN.n29 VSUBS 0.056443f
C730 VN.n30 VSUBS 0.105195f
C731 VN.n31 VSUBS 0.105195f
C732 VN.n32 VSUBS 0.07715f
C733 VN.n33 VSUBS 0.091097f
C734 VN.n34 VSUBS 0.148746f
C735 VN.t0 VSUBS 0.38459f
C736 VN.n35 VSUBS 0.462913f
C737 VN.n36 VSUBS 0.056443f
C738 VN.n37 VSUBS 0.071386f
C739 VN.n38 VSUBS 0.056443f
C740 VN.n39 VSUBS 0.062608f
C741 VN.n40 VSUBS 0.056443f
C742 VN.t7 VSUBS 0.38459f
C743 VN.n41 VSUBS 0.24147f
C744 VN.n42 VSUBS 0.045629f
C745 VN.n43 VSUBS 0.056443f
C746 VN.t6 VSUBS 0.38459f
C747 VN.n44 VSUBS 0.454085f
C748 VN.t3 VSUBS 0.93381f
C749 VN.n45 VSUBS 0.540872f
C750 VN.n46 VSUBS 0.695501f
C751 VN.n47 VSUBS 0.095846f
C752 VN.n48 VSUBS 0.105195f
C753 VN.n49 VSUBS 0.112179f
C754 VN.n50 VSUBS 0.056443f
C755 VN.n51 VSUBS 0.056443f
C756 VN.n52 VSUBS 0.056443f
C757 VN.n53 VSUBS 0.112179f
C758 VN.n54 VSUBS 0.105195f
C759 VN.n55 VSUBS 0.095846f
C760 VN.n56 VSUBS 0.056443f
C761 VN.n57 VSUBS 0.056443f
C762 VN.n58 VSUBS 0.056443f
C763 VN.n59 VSUBS 0.105195f
C764 VN.n60 VSUBS 0.105195f
C765 VN.n61 VSUBS 0.093406f
C766 VN.n62 VSUBS 0.056443f
C767 VN.n63 VSUBS 0.056443f
C768 VN.n64 VSUBS 0.056443f
C769 VN.n65 VSUBS 0.105195f
C770 VN.n66 VSUBS 0.105195f
C771 VN.n67 VSUBS 0.07715f
C772 VN.n68 VSUBS 0.091097f
C773 VN.n69 VSUBS 2.95762f
C774 VDD1.t2 VSUBS 0.022139f
C775 VDD1.t6 VSUBS 0.022139f
C776 VDD1.n0 VSUBS 0.076533f
C777 VDD1.t1 VSUBS 0.022139f
C778 VDD1.t5 VSUBS 0.022139f
C779 VDD1.n1 VSUBS 0.076276f
C780 VDD1.t3 VSUBS 0.022139f
C781 VDD1.t4 VSUBS 0.022139f
C782 VDD1.n2 VSUBS 0.076276f
C783 VDD1.n3 VSUBS 3.44128f
C784 VDD1.t0 VSUBS 0.022139f
C785 VDD1.t7 VSUBS 0.022139f
C786 VDD1.n4 VSUBS 0.073309f
C787 VDD1.n5 VSUBS 2.63829f
C788 VTAIL.t1 VSUBS 0.032127f
C789 VTAIL.t0 VSUBS 0.032127f
C790 VTAIL.n0 VSUBS 0.091536f
C791 VTAIL.n1 VSUBS 0.687187f
C792 VTAIL.t2 VSUBS 0.161332f
C793 VTAIL.n2 VSUBS 0.757366f
C794 VTAIL.t8 VSUBS 0.161332f
C795 VTAIL.n3 VSUBS 0.757366f
C796 VTAIL.t11 VSUBS 0.032127f
C797 VTAIL.t9 VSUBS 0.032127f
C798 VTAIL.n4 VSUBS 0.091536f
C799 VTAIL.n5 VSUBS 1.09862f
C800 VTAIL.t12 VSUBS 0.161332f
C801 VTAIL.n6 VSUBS 1.76556f
C802 VTAIL.t6 VSUBS 0.161332f
C803 VTAIL.n7 VSUBS 1.76556f
C804 VTAIL.t7 VSUBS 0.032127f
C805 VTAIL.t5 VSUBS 0.032127f
C806 VTAIL.n8 VSUBS 0.091536f
C807 VTAIL.n9 VSUBS 1.09862f
C808 VTAIL.t4 VSUBS 0.161332f
C809 VTAIL.n10 VSUBS 0.757366f
C810 VTAIL.t10 VSUBS 0.161332f
C811 VTAIL.n11 VSUBS 0.757366f
C812 VTAIL.t15 VSUBS 0.032127f
C813 VTAIL.t13 VSUBS 0.032127f
C814 VTAIL.n12 VSUBS 0.091536f
C815 VTAIL.n13 VSUBS 1.09862f
C816 VTAIL.t14 VSUBS 0.161332f
C817 VTAIL.n14 VSUBS 1.76556f
C818 VTAIL.t3 VSUBS 0.161332f
C819 VTAIL.n15 VSUBS 1.75815f
C820 VP.t3 VSUBS 0.445887f
C821 VP.n0 VSUBS 0.536693f
C822 VP.n1 VSUBS 0.065438f
C823 VP.n2 VSUBS 0.082764f
C824 VP.n3 VSUBS 0.065438f
C825 VP.n4 VSUBS 0.072586f
C826 VP.n5 VSUBS 0.065438f
C827 VP.n6 VSUBS 0.052901f
C828 VP.n7 VSUBS 0.065438f
C829 VP.t2 VSUBS 0.445887f
C830 VP.n8 VSUBS 0.279956f
C831 VP.n9 VSUBS 0.065438f
C832 VP.n10 VSUBS 0.108293f
C833 VP.n11 VSUBS 0.065438f
C834 VP.n12 VSUBS 0.089446f
C835 VP.t0 VSUBS 0.445887f
C836 VP.n13 VSUBS 0.536693f
C837 VP.n14 VSUBS 0.065438f
C838 VP.n15 VSUBS 0.082764f
C839 VP.n16 VSUBS 0.065438f
C840 VP.n17 VSUBS 0.072586f
C841 VP.n18 VSUBS 0.065438f
C842 VP.n19 VSUBS 0.052901f
C843 VP.n20 VSUBS 0.065438f
C844 VP.t1 VSUBS 0.445887f
C845 VP.n21 VSUBS 0.526457f
C846 VP.t5 VSUBS 1.08264f
C847 VP.n22 VSUBS 0.627077f
C848 VP.n23 VSUBS 0.806352f
C849 VP.n24 VSUBS 0.111123f
C850 VP.n25 VSUBS 0.121961f
C851 VP.n26 VSUBS 0.130058f
C852 VP.n27 VSUBS 0.065438f
C853 VP.n28 VSUBS 0.065438f
C854 VP.n29 VSUBS 0.065438f
C855 VP.n30 VSUBS 0.130058f
C856 VP.n31 VSUBS 0.121961f
C857 VP.t7 VSUBS 0.445887f
C858 VP.n32 VSUBS 0.279956f
C859 VP.n33 VSUBS 0.111123f
C860 VP.n34 VSUBS 0.065438f
C861 VP.n35 VSUBS 0.065438f
C862 VP.n36 VSUBS 0.065438f
C863 VP.n37 VSUBS 0.121961f
C864 VP.n38 VSUBS 0.121961f
C865 VP.n39 VSUBS 0.108293f
C866 VP.n40 VSUBS 0.065438f
C867 VP.n41 VSUBS 0.065438f
C868 VP.n42 VSUBS 0.065438f
C869 VP.n43 VSUBS 0.121961f
C870 VP.n44 VSUBS 0.121961f
C871 VP.n45 VSUBS 0.089446f
C872 VP.n46 VSUBS 0.105616f
C873 VP.n47 VSUBS 3.40163f
C874 VP.t6 VSUBS 0.445887f
C875 VP.n48 VSUBS 0.536693f
C876 VP.n49 VSUBS 3.45183f
C877 VP.n50 VSUBS 0.105616f
C878 VP.n51 VSUBS 0.065438f
C879 VP.n52 VSUBS 0.121961f
C880 VP.n53 VSUBS 0.121961f
C881 VP.n54 VSUBS 0.082764f
C882 VP.n55 VSUBS 0.065438f
C883 VP.n56 VSUBS 0.065438f
C884 VP.n57 VSUBS 0.065438f
C885 VP.n58 VSUBS 0.121961f
C886 VP.n59 VSUBS 0.121961f
C887 VP.n60 VSUBS 0.072586f
C888 VP.n61 VSUBS 0.065438f
C889 VP.n62 VSUBS 0.065438f
C890 VP.n63 VSUBS 0.111123f
C891 VP.n64 VSUBS 0.121961f
C892 VP.n65 VSUBS 0.130058f
C893 VP.n66 VSUBS 0.065438f
C894 VP.n67 VSUBS 0.065438f
C895 VP.n68 VSUBS 0.065438f
C896 VP.n69 VSUBS 0.130058f
C897 VP.n70 VSUBS 0.121961f
C898 VP.t4 VSUBS 0.445887f
C899 VP.n71 VSUBS 0.279956f
C900 VP.n72 VSUBS 0.111123f
C901 VP.n73 VSUBS 0.065438f
C902 VP.n74 VSUBS 0.065438f
C903 VP.n75 VSUBS 0.065438f
C904 VP.n76 VSUBS 0.121961f
C905 VP.n77 VSUBS 0.121961f
C906 VP.n78 VSUBS 0.108293f
C907 VP.n79 VSUBS 0.065438f
C908 VP.n80 VSUBS 0.065438f
C909 VP.n81 VSUBS 0.065438f
C910 VP.n82 VSUBS 0.121961f
C911 VP.n83 VSUBS 0.121961f
C912 VP.n84 VSUBS 0.089446f
C913 VP.n85 VSUBS 0.105616f
C914 VP.n86 VSUBS 0.172453f
.ends

