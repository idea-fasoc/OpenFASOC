* NGSPICE file created from diff_pair_sample_1190.ext - technology: sky130A

.subckt diff_pair_sample_1190 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0.31185 ps=2.22 w=1.89 l=0.82
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0 ps=0 w=1.89 l=0.82
X2 VTAIL.t10 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.31185 ps=2.22 w=1.89 l=0.82
X3 VTAIL.t5 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.31185 ps=2.22 w=1.89 l=0.82
X4 VTAIL.t7 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.31185 ps=2.22 w=1.89 l=0.82
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0 ps=0 w=1.89 l=0.82
X6 VTAIL.t4 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.31185 ps=2.22 w=1.89 l=0.82
X7 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0.31185 ps=2.22 w=1.89 l=0.82
X8 VDD2.t2 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.7371 ps=4.56 w=1.89 l=0.82
X9 VDD2.t1 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0.31185 ps=2.22 w=1.89 l=0.82
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0 ps=0 w=1.89 l=0.82
X11 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0.31185 ps=2.22 w=1.89 l=0.82
X12 VDD1.t1 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.7371 ps=4.56 w=1.89 l=0.82
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7371 pd=4.56 as=0 ps=0 w=1.89 l=0.82
X14 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.7371 ps=4.56 w=1.89 l=0.82
X15 VDD2.t0 VN.t5 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.31185 pd=2.22 as=0.7371 ps=4.56 w=1.89 l=0.82
R0 VN.n9 VN.n6 161.3
R1 VN.n3 VN.n0 161.3
R2 VN.n1 VN.t4 118.945
R3 VN.n7 VN.t3 118.945
R4 VN.n4 VN.t5 103.749
R5 VN.n10 VN.t0 103.749
R6 VN.n11 VN.n10 80.6037
R7 VN.n5 VN.n4 80.6037
R8 VN.n4 VN.n3 56.0299
R9 VN.n10 VN.n9 56.0299
R10 VN.n2 VN.t2 55.5481
R11 VN.n8 VN.t1 55.5481
R12 VN.n7 VN.n6 43.941
R13 VN.n1 VN.n0 43.941
R14 VN.n2 VN.n1 42.5398
R15 VN.n8 VN.n7 42.5398
R16 VN VN.n11 34.4195
R17 VN.n3 VN.n2 12.234
R18 VN.n9 VN.n8 12.234
R19 VN.n11 VN.n6 0.285035
R20 VN.n5 VN.n0 0.285035
R21 VN VN.n5 0.146778
R22 VTAIL.n34 VTAIL.n32 289.615
R23 VTAIL.n4 VTAIL.n2 289.615
R24 VTAIL.n26 VTAIL.n24 289.615
R25 VTAIL.n16 VTAIL.n14 289.615
R26 VTAIL.n35 VTAIL.n34 185
R27 VTAIL.n5 VTAIL.n4 185
R28 VTAIL.n27 VTAIL.n26 185
R29 VTAIL.n17 VTAIL.n16 185
R30 VTAIL.t9 VTAIL.n33 164.876
R31 VTAIL.t2 VTAIL.n3 164.876
R32 VTAIL.t3 VTAIL.n25 164.876
R33 VTAIL.t8 VTAIL.n15 164.876
R34 VTAIL.n23 VTAIL.n22 86.8776
R35 VTAIL.n13 VTAIL.n12 86.8776
R36 VTAIL.n1 VTAIL.n0 86.8776
R37 VTAIL.n11 VTAIL.n10 86.8776
R38 VTAIL.n34 VTAIL.t9 52.3082
R39 VTAIL.n4 VTAIL.t2 52.3082
R40 VTAIL.n26 VTAIL.t3 52.3082
R41 VTAIL.n16 VTAIL.t8 52.3082
R42 VTAIL.n39 VTAIL.n38 36.2581
R43 VTAIL.n9 VTAIL.n8 36.2581
R44 VTAIL.n31 VTAIL.n30 36.2581
R45 VTAIL.n21 VTAIL.n20 36.2581
R46 VTAIL.n13 VTAIL.n11 15.9789
R47 VTAIL.n39 VTAIL.n31 14.9876
R48 VTAIL.n35 VTAIL.n33 14.7318
R49 VTAIL.n5 VTAIL.n3 14.7318
R50 VTAIL.n27 VTAIL.n25 14.7318
R51 VTAIL.n17 VTAIL.n15 14.7318
R52 VTAIL.n36 VTAIL.n32 12.8005
R53 VTAIL.n6 VTAIL.n2 12.8005
R54 VTAIL.n28 VTAIL.n24 12.8005
R55 VTAIL.n18 VTAIL.n14 12.8005
R56 VTAIL.n0 VTAIL.t6 10.4767
R57 VTAIL.n0 VTAIL.t7 10.4767
R58 VTAIL.n10 VTAIL.t1 10.4767
R59 VTAIL.n10 VTAIL.t4 10.4767
R60 VTAIL.n22 VTAIL.t0 10.4767
R61 VTAIL.n22 VTAIL.t5 10.4767
R62 VTAIL.n12 VTAIL.t11 10.4767
R63 VTAIL.n12 VTAIL.t10 10.4767
R64 VTAIL.n38 VTAIL.n37 9.45567
R65 VTAIL.n8 VTAIL.n7 9.45567
R66 VTAIL.n30 VTAIL.n29 9.45567
R67 VTAIL.n20 VTAIL.n19 9.45567
R68 VTAIL.n37 VTAIL.n36 9.3005
R69 VTAIL.n7 VTAIL.n6 9.3005
R70 VTAIL.n29 VTAIL.n28 9.3005
R71 VTAIL.n19 VTAIL.n18 9.3005
R72 VTAIL.n37 VTAIL.n33 5.62509
R73 VTAIL.n7 VTAIL.n3 5.62509
R74 VTAIL.n29 VTAIL.n25 5.62509
R75 VTAIL.n19 VTAIL.n15 5.62509
R76 VTAIL.n38 VTAIL.n32 1.16414
R77 VTAIL.n8 VTAIL.n2 1.16414
R78 VTAIL.n30 VTAIL.n24 1.16414
R79 VTAIL.n20 VTAIL.n14 1.16414
R80 VTAIL.n21 VTAIL.n13 0.991879
R81 VTAIL.n31 VTAIL.n23 0.991879
R82 VTAIL.n11 VTAIL.n9 0.991879
R83 VTAIL.n23 VTAIL.n21 0.966017
R84 VTAIL.n9 VTAIL.n1 0.966017
R85 VTAIL VTAIL.n39 0.685845
R86 VTAIL.n36 VTAIL.n35 0.388379
R87 VTAIL.n6 VTAIL.n5 0.388379
R88 VTAIL.n28 VTAIL.n27 0.388379
R89 VTAIL.n18 VTAIL.n17 0.388379
R90 VTAIL VTAIL.n1 0.306534
R91 VDD2.n11 VDD2.n9 289.615
R92 VDD2.n2 VDD2.n0 289.615
R93 VDD2.n12 VDD2.n11 185
R94 VDD2.n3 VDD2.n2 185
R95 VDD2.t5 VDD2.n10 164.876
R96 VDD2.t1 VDD2.n1 164.876
R97 VDD2.n8 VDD2.n7 103.749
R98 VDD2 VDD2.n17 103.746
R99 VDD2.n8 VDD2.n6 53.625
R100 VDD2.n16 VDD2.n15 52.9369
R101 VDD2.n11 VDD2.t5 52.3082
R102 VDD2.n2 VDD2.t1 52.3082
R103 VDD2.n16 VDD2.n8 28.5666
R104 VDD2.n12 VDD2.n10 14.7318
R105 VDD2.n3 VDD2.n1 14.7318
R106 VDD2.n13 VDD2.n9 12.8005
R107 VDD2.n4 VDD2.n0 12.8005
R108 VDD2.n17 VDD2.t4 10.4767
R109 VDD2.n17 VDD2.t2 10.4767
R110 VDD2.n7 VDD2.t3 10.4767
R111 VDD2.n7 VDD2.t0 10.4767
R112 VDD2.n15 VDD2.n14 9.45567
R113 VDD2.n6 VDD2.n5 9.45567
R114 VDD2.n14 VDD2.n13 9.3005
R115 VDD2.n5 VDD2.n4 9.3005
R116 VDD2.n14 VDD2.n10 5.62509
R117 VDD2.n5 VDD2.n1 5.62509
R118 VDD2.n15 VDD2.n9 1.16414
R119 VDD2.n6 VDD2.n0 1.16414
R120 VDD2 VDD2.n16 0.802224
R121 VDD2.n13 VDD2.n12 0.388379
R122 VDD2.n4 VDD2.n3 0.388379
R123 B.n350 B.n349 585
R124 B.n351 B.n350 585
R125 B.n128 B.n59 585
R126 B.n127 B.n126 585
R127 B.n125 B.n124 585
R128 B.n123 B.n122 585
R129 B.n121 B.n120 585
R130 B.n119 B.n118 585
R131 B.n117 B.n116 585
R132 B.n115 B.n114 585
R133 B.n113 B.n112 585
R134 B.n111 B.n110 585
R135 B.n109 B.n108 585
R136 B.n106 B.n105 585
R137 B.n104 B.n103 585
R138 B.n102 B.n101 585
R139 B.n100 B.n99 585
R140 B.n98 B.n97 585
R141 B.n96 B.n95 585
R142 B.n94 B.n93 585
R143 B.n92 B.n91 585
R144 B.n90 B.n89 585
R145 B.n88 B.n87 585
R146 B.n86 B.n85 585
R147 B.n84 B.n83 585
R148 B.n82 B.n81 585
R149 B.n80 B.n79 585
R150 B.n78 B.n77 585
R151 B.n76 B.n75 585
R152 B.n74 B.n73 585
R153 B.n72 B.n71 585
R154 B.n70 B.n69 585
R155 B.n68 B.n67 585
R156 B.n66 B.n65 585
R157 B.n348 B.n42 585
R158 B.n352 B.n42 585
R159 B.n347 B.n41 585
R160 B.n353 B.n41 585
R161 B.n346 B.n345 585
R162 B.n345 B.n37 585
R163 B.n344 B.n36 585
R164 B.n359 B.n36 585
R165 B.n343 B.n35 585
R166 B.n360 B.n35 585
R167 B.n342 B.n34 585
R168 B.n361 B.n34 585
R169 B.n341 B.n340 585
R170 B.n340 B.n30 585
R171 B.n339 B.n29 585
R172 B.n367 B.n29 585
R173 B.n338 B.n28 585
R174 B.n368 B.n28 585
R175 B.n337 B.n27 585
R176 B.n369 B.n27 585
R177 B.n336 B.n335 585
R178 B.n335 B.n23 585
R179 B.n334 B.n22 585
R180 B.n375 B.n22 585
R181 B.n333 B.n21 585
R182 B.n376 B.n21 585
R183 B.n332 B.n20 585
R184 B.n377 B.n20 585
R185 B.n331 B.n330 585
R186 B.n330 B.n19 585
R187 B.n329 B.n15 585
R188 B.n383 B.n15 585
R189 B.n328 B.n14 585
R190 B.n384 B.n14 585
R191 B.n327 B.n13 585
R192 B.n385 B.n13 585
R193 B.n326 B.n325 585
R194 B.n325 B.n12 585
R195 B.n324 B.n323 585
R196 B.n324 B.n8 585
R197 B.n322 B.n7 585
R198 B.n392 B.n7 585
R199 B.n321 B.n6 585
R200 B.n393 B.n6 585
R201 B.n320 B.n5 585
R202 B.n394 B.n5 585
R203 B.n319 B.n318 585
R204 B.n318 B.n4 585
R205 B.n317 B.n129 585
R206 B.n317 B.n316 585
R207 B.n306 B.n130 585
R208 B.n309 B.n130 585
R209 B.n308 B.n307 585
R210 B.n310 B.n308 585
R211 B.n305 B.n135 585
R212 B.n135 B.n134 585
R213 B.n304 B.n303 585
R214 B.n303 B.n302 585
R215 B.n137 B.n136 585
R216 B.n295 B.n137 585
R217 B.n294 B.n293 585
R218 B.n296 B.n294 585
R219 B.n292 B.n142 585
R220 B.n142 B.n141 585
R221 B.n291 B.n290 585
R222 B.n290 B.n289 585
R223 B.n144 B.n143 585
R224 B.n145 B.n144 585
R225 B.n282 B.n281 585
R226 B.n283 B.n282 585
R227 B.n280 B.n150 585
R228 B.n150 B.n149 585
R229 B.n279 B.n278 585
R230 B.n278 B.n277 585
R231 B.n152 B.n151 585
R232 B.n153 B.n152 585
R233 B.n270 B.n269 585
R234 B.n271 B.n270 585
R235 B.n268 B.n157 585
R236 B.n161 B.n157 585
R237 B.n267 B.n266 585
R238 B.n266 B.n265 585
R239 B.n159 B.n158 585
R240 B.n160 B.n159 585
R241 B.n258 B.n257 585
R242 B.n259 B.n258 585
R243 B.n256 B.n166 585
R244 B.n166 B.n165 585
R245 B.n250 B.n249 585
R246 B.n248 B.n184 585
R247 B.n247 B.n183 585
R248 B.n252 B.n183 585
R249 B.n246 B.n245 585
R250 B.n244 B.n243 585
R251 B.n242 B.n241 585
R252 B.n240 B.n239 585
R253 B.n238 B.n237 585
R254 B.n236 B.n235 585
R255 B.n234 B.n233 585
R256 B.n232 B.n231 585
R257 B.n230 B.n229 585
R258 B.n227 B.n226 585
R259 B.n225 B.n224 585
R260 B.n223 B.n222 585
R261 B.n221 B.n220 585
R262 B.n219 B.n218 585
R263 B.n217 B.n216 585
R264 B.n215 B.n214 585
R265 B.n213 B.n212 585
R266 B.n211 B.n210 585
R267 B.n209 B.n208 585
R268 B.n207 B.n206 585
R269 B.n205 B.n204 585
R270 B.n203 B.n202 585
R271 B.n201 B.n200 585
R272 B.n199 B.n198 585
R273 B.n197 B.n196 585
R274 B.n195 B.n194 585
R275 B.n193 B.n192 585
R276 B.n191 B.n190 585
R277 B.n168 B.n167 585
R278 B.n255 B.n254 585
R279 B.n164 B.n163 585
R280 B.n165 B.n164 585
R281 B.n261 B.n260 585
R282 B.n260 B.n259 585
R283 B.n262 B.n162 585
R284 B.n162 B.n160 585
R285 B.n264 B.n263 585
R286 B.n265 B.n264 585
R287 B.n156 B.n155 585
R288 B.n161 B.n156 585
R289 B.n273 B.n272 585
R290 B.n272 B.n271 585
R291 B.n274 B.n154 585
R292 B.n154 B.n153 585
R293 B.n276 B.n275 585
R294 B.n277 B.n276 585
R295 B.n148 B.n147 585
R296 B.n149 B.n148 585
R297 B.n285 B.n284 585
R298 B.n284 B.n283 585
R299 B.n286 B.n146 585
R300 B.n146 B.n145 585
R301 B.n288 B.n287 585
R302 B.n289 B.n288 585
R303 B.n140 B.n139 585
R304 B.n141 B.n140 585
R305 B.n298 B.n297 585
R306 B.n297 B.n296 585
R307 B.n299 B.n138 585
R308 B.n295 B.n138 585
R309 B.n301 B.n300 585
R310 B.n302 B.n301 585
R311 B.n133 B.n132 585
R312 B.n134 B.n133 585
R313 B.n312 B.n311 585
R314 B.n311 B.n310 585
R315 B.n313 B.n131 585
R316 B.n309 B.n131 585
R317 B.n315 B.n314 585
R318 B.n316 B.n315 585
R319 B.n3 B.n0 585
R320 B.n4 B.n3 585
R321 B.n391 B.n1 585
R322 B.n392 B.n391 585
R323 B.n390 B.n389 585
R324 B.n390 B.n8 585
R325 B.n388 B.n9 585
R326 B.n12 B.n9 585
R327 B.n387 B.n386 585
R328 B.n386 B.n385 585
R329 B.n11 B.n10 585
R330 B.n384 B.n11 585
R331 B.n382 B.n381 585
R332 B.n383 B.n382 585
R333 B.n380 B.n16 585
R334 B.n19 B.n16 585
R335 B.n379 B.n378 585
R336 B.n378 B.n377 585
R337 B.n18 B.n17 585
R338 B.n376 B.n18 585
R339 B.n374 B.n373 585
R340 B.n375 B.n374 585
R341 B.n372 B.n24 585
R342 B.n24 B.n23 585
R343 B.n371 B.n370 585
R344 B.n370 B.n369 585
R345 B.n26 B.n25 585
R346 B.n368 B.n26 585
R347 B.n366 B.n365 585
R348 B.n367 B.n366 585
R349 B.n364 B.n31 585
R350 B.n31 B.n30 585
R351 B.n363 B.n362 585
R352 B.n362 B.n361 585
R353 B.n33 B.n32 585
R354 B.n360 B.n33 585
R355 B.n358 B.n357 585
R356 B.n359 B.n358 585
R357 B.n356 B.n38 585
R358 B.n38 B.n37 585
R359 B.n355 B.n354 585
R360 B.n354 B.n353 585
R361 B.n40 B.n39 585
R362 B.n352 B.n40 585
R363 B.n395 B.n394 585
R364 B.n393 B.n2 585
R365 B.n65 B.n40 550.159
R366 B.n350 B.n42 550.159
R367 B.n254 B.n166 550.159
R368 B.n250 B.n164 550.159
R369 B.n62 B.t17 257.209
R370 B.n60 B.t10 257.209
R371 B.n187 B.t6 257.209
R372 B.n185 B.t14 257.209
R373 B.n351 B.n58 256.663
R374 B.n351 B.n57 256.663
R375 B.n351 B.n56 256.663
R376 B.n351 B.n55 256.663
R377 B.n351 B.n54 256.663
R378 B.n351 B.n53 256.663
R379 B.n351 B.n52 256.663
R380 B.n351 B.n51 256.663
R381 B.n351 B.n50 256.663
R382 B.n351 B.n49 256.663
R383 B.n351 B.n48 256.663
R384 B.n351 B.n47 256.663
R385 B.n351 B.n46 256.663
R386 B.n351 B.n45 256.663
R387 B.n351 B.n44 256.663
R388 B.n351 B.n43 256.663
R389 B.n252 B.n251 256.663
R390 B.n252 B.n169 256.663
R391 B.n252 B.n170 256.663
R392 B.n252 B.n171 256.663
R393 B.n252 B.n172 256.663
R394 B.n252 B.n173 256.663
R395 B.n252 B.n174 256.663
R396 B.n252 B.n175 256.663
R397 B.n252 B.n176 256.663
R398 B.n252 B.n177 256.663
R399 B.n252 B.n178 256.663
R400 B.n252 B.n179 256.663
R401 B.n252 B.n180 256.663
R402 B.n252 B.n181 256.663
R403 B.n252 B.n182 256.663
R404 B.n253 B.n252 256.663
R405 B.n397 B.n396 256.663
R406 B.n252 B.n165 204.188
R407 B.n352 B.n351 204.188
R408 B.n69 B.n68 163.367
R409 B.n73 B.n72 163.367
R410 B.n77 B.n76 163.367
R411 B.n81 B.n80 163.367
R412 B.n85 B.n84 163.367
R413 B.n89 B.n88 163.367
R414 B.n93 B.n92 163.367
R415 B.n97 B.n96 163.367
R416 B.n101 B.n100 163.367
R417 B.n105 B.n104 163.367
R418 B.n110 B.n109 163.367
R419 B.n114 B.n113 163.367
R420 B.n118 B.n117 163.367
R421 B.n122 B.n121 163.367
R422 B.n126 B.n125 163.367
R423 B.n350 B.n59 163.367
R424 B.n258 B.n166 163.367
R425 B.n258 B.n159 163.367
R426 B.n266 B.n159 163.367
R427 B.n266 B.n157 163.367
R428 B.n270 B.n157 163.367
R429 B.n270 B.n152 163.367
R430 B.n278 B.n152 163.367
R431 B.n278 B.n150 163.367
R432 B.n282 B.n150 163.367
R433 B.n282 B.n144 163.367
R434 B.n290 B.n144 163.367
R435 B.n290 B.n142 163.367
R436 B.n294 B.n142 163.367
R437 B.n294 B.n137 163.367
R438 B.n303 B.n137 163.367
R439 B.n303 B.n135 163.367
R440 B.n308 B.n135 163.367
R441 B.n308 B.n130 163.367
R442 B.n317 B.n130 163.367
R443 B.n318 B.n317 163.367
R444 B.n318 B.n5 163.367
R445 B.n6 B.n5 163.367
R446 B.n7 B.n6 163.367
R447 B.n324 B.n7 163.367
R448 B.n325 B.n324 163.367
R449 B.n325 B.n13 163.367
R450 B.n14 B.n13 163.367
R451 B.n15 B.n14 163.367
R452 B.n330 B.n15 163.367
R453 B.n330 B.n20 163.367
R454 B.n21 B.n20 163.367
R455 B.n22 B.n21 163.367
R456 B.n335 B.n22 163.367
R457 B.n335 B.n27 163.367
R458 B.n28 B.n27 163.367
R459 B.n29 B.n28 163.367
R460 B.n340 B.n29 163.367
R461 B.n340 B.n34 163.367
R462 B.n35 B.n34 163.367
R463 B.n36 B.n35 163.367
R464 B.n345 B.n36 163.367
R465 B.n345 B.n41 163.367
R466 B.n42 B.n41 163.367
R467 B.n184 B.n183 163.367
R468 B.n245 B.n183 163.367
R469 B.n243 B.n242 163.367
R470 B.n239 B.n238 163.367
R471 B.n235 B.n234 163.367
R472 B.n231 B.n230 163.367
R473 B.n226 B.n225 163.367
R474 B.n222 B.n221 163.367
R475 B.n218 B.n217 163.367
R476 B.n214 B.n213 163.367
R477 B.n210 B.n209 163.367
R478 B.n206 B.n205 163.367
R479 B.n202 B.n201 163.367
R480 B.n198 B.n197 163.367
R481 B.n194 B.n193 163.367
R482 B.n190 B.n168 163.367
R483 B.n260 B.n164 163.367
R484 B.n260 B.n162 163.367
R485 B.n264 B.n162 163.367
R486 B.n264 B.n156 163.367
R487 B.n272 B.n156 163.367
R488 B.n272 B.n154 163.367
R489 B.n276 B.n154 163.367
R490 B.n276 B.n148 163.367
R491 B.n284 B.n148 163.367
R492 B.n284 B.n146 163.367
R493 B.n288 B.n146 163.367
R494 B.n288 B.n140 163.367
R495 B.n297 B.n140 163.367
R496 B.n297 B.n138 163.367
R497 B.n301 B.n138 163.367
R498 B.n301 B.n133 163.367
R499 B.n311 B.n133 163.367
R500 B.n311 B.n131 163.367
R501 B.n315 B.n131 163.367
R502 B.n315 B.n3 163.367
R503 B.n395 B.n3 163.367
R504 B.n391 B.n2 163.367
R505 B.n391 B.n390 163.367
R506 B.n390 B.n9 163.367
R507 B.n386 B.n9 163.367
R508 B.n386 B.n11 163.367
R509 B.n382 B.n11 163.367
R510 B.n382 B.n16 163.367
R511 B.n378 B.n16 163.367
R512 B.n378 B.n18 163.367
R513 B.n374 B.n18 163.367
R514 B.n374 B.n24 163.367
R515 B.n370 B.n24 163.367
R516 B.n370 B.n26 163.367
R517 B.n366 B.n26 163.367
R518 B.n366 B.n31 163.367
R519 B.n362 B.n31 163.367
R520 B.n362 B.n33 163.367
R521 B.n358 B.n33 163.367
R522 B.n358 B.n38 163.367
R523 B.n354 B.n38 163.367
R524 B.n354 B.n40 163.367
R525 B.n60 B.t12 143.189
R526 B.n187 B.t9 143.189
R527 B.n62 B.t18 143.189
R528 B.n185 B.t16 143.189
R529 B.n61 B.t13 120.885
R530 B.n188 B.t8 120.885
R531 B.n63 B.t19 120.885
R532 B.n186 B.t15 120.885
R533 B.n259 B.n165 104.397
R534 B.n259 B.n160 104.397
R535 B.n265 B.n160 104.397
R536 B.n265 B.n161 104.397
R537 B.n271 B.n153 104.397
R538 B.n277 B.n153 104.397
R539 B.n277 B.n149 104.397
R540 B.n283 B.n149 104.397
R541 B.n283 B.n145 104.397
R542 B.n289 B.n145 104.397
R543 B.n296 B.n141 104.397
R544 B.n296 B.n295 104.397
R545 B.n302 B.n134 104.397
R546 B.n310 B.n134 104.397
R547 B.n310 B.n309 104.397
R548 B.n316 B.n4 104.397
R549 B.n394 B.n4 104.397
R550 B.n394 B.n393 104.397
R551 B.n393 B.n392 104.397
R552 B.n392 B.n8 104.397
R553 B.n385 B.n12 104.397
R554 B.n385 B.n384 104.397
R555 B.n384 B.n383 104.397
R556 B.n377 B.n19 104.397
R557 B.n377 B.n376 104.397
R558 B.n375 B.n23 104.397
R559 B.n369 B.n23 104.397
R560 B.n369 B.n368 104.397
R561 B.n368 B.n367 104.397
R562 B.n367 B.n30 104.397
R563 B.n361 B.n30 104.397
R564 B.n360 B.n359 104.397
R565 B.n359 B.n37 104.397
R566 B.n353 B.n37 104.397
R567 B.n353 B.n352 104.397
R568 B.n161 B.t7 89.0445
R569 B.t11 B.n360 89.0445
R570 B.n295 B.t4 85.974
R571 B.n19 B.t5 85.974
R572 B.n316 B.t2 82.9035
R573 B.t0 B.n8 82.9035
R574 B.n65 B.n43 71.676
R575 B.n69 B.n44 71.676
R576 B.n73 B.n45 71.676
R577 B.n77 B.n46 71.676
R578 B.n81 B.n47 71.676
R579 B.n85 B.n48 71.676
R580 B.n89 B.n49 71.676
R581 B.n93 B.n50 71.676
R582 B.n97 B.n51 71.676
R583 B.n101 B.n52 71.676
R584 B.n105 B.n53 71.676
R585 B.n110 B.n54 71.676
R586 B.n114 B.n55 71.676
R587 B.n118 B.n56 71.676
R588 B.n122 B.n57 71.676
R589 B.n126 B.n58 71.676
R590 B.n59 B.n58 71.676
R591 B.n125 B.n57 71.676
R592 B.n121 B.n56 71.676
R593 B.n117 B.n55 71.676
R594 B.n113 B.n54 71.676
R595 B.n109 B.n53 71.676
R596 B.n104 B.n52 71.676
R597 B.n100 B.n51 71.676
R598 B.n96 B.n50 71.676
R599 B.n92 B.n49 71.676
R600 B.n88 B.n48 71.676
R601 B.n84 B.n47 71.676
R602 B.n80 B.n46 71.676
R603 B.n76 B.n45 71.676
R604 B.n72 B.n44 71.676
R605 B.n68 B.n43 71.676
R606 B.n251 B.n250 71.676
R607 B.n245 B.n169 71.676
R608 B.n242 B.n170 71.676
R609 B.n238 B.n171 71.676
R610 B.n234 B.n172 71.676
R611 B.n230 B.n173 71.676
R612 B.n225 B.n174 71.676
R613 B.n221 B.n175 71.676
R614 B.n217 B.n176 71.676
R615 B.n213 B.n177 71.676
R616 B.n209 B.n178 71.676
R617 B.n205 B.n179 71.676
R618 B.n201 B.n180 71.676
R619 B.n197 B.n181 71.676
R620 B.n193 B.n182 71.676
R621 B.n253 B.n168 71.676
R622 B.n251 B.n184 71.676
R623 B.n243 B.n169 71.676
R624 B.n239 B.n170 71.676
R625 B.n235 B.n171 71.676
R626 B.n231 B.n172 71.676
R627 B.n226 B.n173 71.676
R628 B.n222 B.n174 71.676
R629 B.n218 B.n175 71.676
R630 B.n214 B.n176 71.676
R631 B.n210 B.n177 71.676
R632 B.n206 B.n178 71.676
R633 B.n202 B.n179 71.676
R634 B.n198 B.n180 71.676
R635 B.n194 B.n181 71.676
R636 B.n190 B.n182 71.676
R637 B.n254 B.n253 71.676
R638 B.n396 B.n395 71.676
R639 B.n396 B.n2 71.676
R640 B.n64 B.n63 59.5399
R641 B.n107 B.n61 59.5399
R642 B.n189 B.n188 59.5399
R643 B.n228 B.n186 59.5399
R644 B.t1 B.n141 58.3396
R645 B.n376 B.t3 58.3396
R646 B.n289 B.t1 46.0577
R647 B.t3 B.n375 46.0577
R648 B.n249 B.n163 35.7468
R649 B.n256 B.n255 35.7468
R650 B.n66 B.n39 35.7468
R651 B.n349 B.n348 35.7468
R652 B.n63 B.n62 22.3035
R653 B.n61 B.n60 22.3035
R654 B.n188 B.n187 22.3035
R655 B.n186 B.n185 22.3035
R656 B.n309 B.t2 21.4939
R657 B.n12 B.t0 21.4939
R658 B.n302 B.t4 18.4234
R659 B.n383 B.t5 18.4234
R660 B B.n397 18.0485
R661 B.n271 B.t7 15.3529
R662 B.n361 B.t11 15.3529
R663 B.n261 B.n163 10.6151
R664 B.n262 B.n261 10.6151
R665 B.n263 B.n262 10.6151
R666 B.n263 B.n155 10.6151
R667 B.n273 B.n155 10.6151
R668 B.n274 B.n273 10.6151
R669 B.n275 B.n274 10.6151
R670 B.n275 B.n147 10.6151
R671 B.n285 B.n147 10.6151
R672 B.n286 B.n285 10.6151
R673 B.n287 B.n286 10.6151
R674 B.n287 B.n139 10.6151
R675 B.n298 B.n139 10.6151
R676 B.n299 B.n298 10.6151
R677 B.n300 B.n299 10.6151
R678 B.n300 B.n132 10.6151
R679 B.n312 B.n132 10.6151
R680 B.n313 B.n312 10.6151
R681 B.n314 B.n313 10.6151
R682 B.n314 B.n0 10.6151
R683 B.n249 B.n248 10.6151
R684 B.n248 B.n247 10.6151
R685 B.n247 B.n246 10.6151
R686 B.n246 B.n244 10.6151
R687 B.n244 B.n241 10.6151
R688 B.n241 B.n240 10.6151
R689 B.n240 B.n237 10.6151
R690 B.n237 B.n236 10.6151
R691 B.n236 B.n233 10.6151
R692 B.n233 B.n232 10.6151
R693 B.n232 B.n229 10.6151
R694 B.n227 B.n224 10.6151
R695 B.n224 B.n223 10.6151
R696 B.n223 B.n220 10.6151
R697 B.n220 B.n219 10.6151
R698 B.n219 B.n216 10.6151
R699 B.n216 B.n215 10.6151
R700 B.n215 B.n212 10.6151
R701 B.n212 B.n211 10.6151
R702 B.n208 B.n207 10.6151
R703 B.n207 B.n204 10.6151
R704 B.n204 B.n203 10.6151
R705 B.n203 B.n200 10.6151
R706 B.n200 B.n199 10.6151
R707 B.n199 B.n196 10.6151
R708 B.n196 B.n195 10.6151
R709 B.n195 B.n192 10.6151
R710 B.n192 B.n191 10.6151
R711 B.n191 B.n167 10.6151
R712 B.n255 B.n167 10.6151
R713 B.n257 B.n256 10.6151
R714 B.n257 B.n158 10.6151
R715 B.n267 B.n158 10.6151
R716 B.n268 B.n267 10.6151
R717 B.n269 B.n268 10.6151
R718 B.n269 B.n151 10.6151
R719 B.n279 B.n151 10.6151
R720 B.n280 B.n279 10.6151
R721 B.n281 B.n280 10.6151
R722 B.n281 B.n143 10.6151
R723 B.n291 B.n143 10.6151
R724 B.n292 B.n291 10.6151
R725 B.n293 B.n292 10.6151
R726 B.n293 B.n136 10.6151
R727 B.n304 B.n136 10.6151
R728 B.n305 B.n304 10.6151
R729 B.n307 B.n305 10.6151
R730 B.n307 B.n306 10.6151
R731 B.n306 B.n129 10.6151
R732 B.n319 B.n129 10.6151
R733 B.n320 B.n319 10.6151
R734 B.n321 B.n320 10.6151
R735 B.n322 B.n321 10.6151
R736 B.n323 B.n322 10.6151
R737 B.n326 B.n323 10.6151
R738 B.n327 B.n326 10.6151
R739 B.n328 B.n327 10.6151
R740 B.n329 B.n328 10.6151
R741 B.n331 B.n329 10.6151
R742 B.n332 B.n331 10.6151
R743 B.n333 B.n332 10.6151
R744 B.n334 B.n333 10.6151
R745 B.n336 B.n334 10.6151
R746 B.n337 B.n336 10.6151
R747 B.n338 B.n337 10.6151
R748 B.n339 B.n338 10.6151
R749 B.n341 B.n339 10.6151
R750 B.n342 B.n341 10.6151
R751 B.n343 B.n342 10.6151
R752 B.n344 B.n343 10.6151
R753 B.n346 B.n344 10.6151
R754 B.n347 B.n346 10.6151
R755 B.n348 B.n347 10.6151
R756 B.n389 B.n1 10.6151
R757 B.n389 B.n388 10.6151
R758 B.n388 B.n387 10.6151
R759 B.n387 B.n10 10.6151
R760 B.n381 B.n10 10.6151
R761 B.n381 B.n380 10.6151
R762 B.n380 B.n379 10.6151
R763 B.n379 B.n17 10.6151
R764 B.n373 B.n17 10.6151
R765 B.n373 B.n372 10.6151
R766 B.n372 B.n371 10.6151
R767 B.n371 B.n25 10.6151
R768 B.n365 B.n25 10.6151
R769 B.n365 B.n364 10.6151
R770 B.n364 B.n363 10.6151
R771 B.n363 B.n32 10.6151
R772 B.n357 B.n32 10.6151
R773 B.n357 B.n356 10.6151
R774 B.n356 B.n355 10.6151
R775 B.n355 B.n39 10.6151
R776 B.n67 B.n66 10.6151
R777 B.n70 B.n67 10.6151
R778 B.n71 B.n70 10.6151
R779 B.n74 B.n71 10.6151
R780 B.n75 B.n74 10.6151
R781 B.n78 B.n75 10.6151
R782 B.n79 B.n78 10.6151
R783 B.n82 B.n79 10.6151
R784 B.n83 B.n82 10.6151
R785 B.n86 B.n83 10.6151
R786 B.n87 B.n86 10.6151
R787 B.n91 B.n90 10.6151
R788 B.n94 B.n91 10.6151
R789 B.n95 B.n94 10.6151
R790 B.n98 B.n95 10.6151
R791 B.n99 B.n98 10.6151
R792 B.n102 B.n99 10.6151
R793 B.n103 B.n102 10.6151
R794 B.n106 B.n103 10.6151
R795 B.n111 B.n108 10.6151
R796 B.n112 B.n111 10.6151
R797 B.n115 B.n112 10.6151
R798 B.n116 B.n115 10.6151
R799 B.n119 B.n116 10.6151
R800 B.n120 B.n119 10.6151
R801 B.n123 B.n120 10.6151
R802 B.n124 B.n123 10.6151
R803 B.n127 B.n124 10.6151
R804 B.n128 B.n127 10.6151
R805 B.n349 B.n128 10.6151
R806 B.n397 B.n0 8.11757
R807 B.n397 B.n1 8.11757
R808 B.n228 B.n227 6.5566
R809 B.n211 B.n189 6.5566
R810 B.n90 B.n64 6.5566
R811 B.n107 B.n106 6.5566
R812 B.n229 B.n228 4.05904
R813 B.n208 B.n189 4.05904
R814 B.n87 B.n64 4.05904
R815 B.n108 B.n107 4.05904
R816 VP.n5 VP.n2 161.3
R817 VP.n12 VP.n0 161.3
R818 VP.n10 VP.n9 161.3
R819 VP.n3 VP.t2 118.945
R820 VP.n1 VP.t3 103.749
R821 VP.n13 VP.t4 103.749
R822 VP.n6 VP.t5 103.749
R823 VP.n7 VP.n6 80.6037
R824 VP.n14 VP.n13 80.6037
R825 VP.n8 VP.n1 80.6037
R826 VP.n10 VP.n1 56.0299
R827 VP.n13 VP.n12 56.0299
R828 VP.n6 VP.n5 56.0299
R829 VP.n11 VP.t1 55.5481
R830 VP.n4 VP.t0 55.5481
R831 VP.n3 VP.n2 43.941
R832 VP.n4 VP.n3 42.5398
R833 VP.n8 VP.n7 34.134
R834 VP.n11 VP.n10 12.234
R835 VP.n12 VP.n11 12.234
R836 VP.n5 VP.n4 12.234
R837 VP.n7 VP.n2 0.285035
R838 VP.n9 VP.n8 0.285035
R839 VP.n14 VP.n0 0.285035
R840 VP.n9 VP.n0 0.189894
R841 VP VP.n14 0.146778
R842 VDD1.n2 VDD1.n0 289.615
R843 VDD1.n9 VDD1.n7 289.615
R844 VDD1.n3 VDD1.n2 185
R845 VDD1.n10 VDD1.n9 185
R846 VDD1.t3 VDD1.n1 164.876
R847 VDD1.t2 VDD1.n8 164.876
R848 VDD1.n15 VDD1.n14 103.749
R849 VDD1.n17 VDD1.n16 103.556
R850 VDD1 VDD1.n6 53.7386
R851 VDD1.n15 VDD1.n13 53.625
R852 VDD1.n2 VDD1.t3 52.3082
R853 VDD1.n9 VDD1.t2 52.3082
R854 VDD1.n17 VDD1.n15 29.6453
R855 VDD1.n3 VDD1.n1 14.7318
R856 VDD1.n10 VDD1.n8 14.7318
R857 VDD1.n4 VDD1.n0 12.8005
R858 VDD1.n11 VDD1.n7 12.8005
R859 VDD1.n16 VDD1.t5 10.4767
R860 VDD1.n16 VDD1.t0 10.4767
R861 VDD1.n14 VDD1.t4 10.4767
R862 VDD1.n14 VDD1.t1 10.4767
R863 VDD1.n6 VDD1.n5 9.45567
R864 VDD1.n13 VDD1.n12 9.45567
R865 VDD1.n5 VDD1.n4 9.3005
R866 VDD1.n12 VDD1.n11 9.3005
R867 VDD1.n5 VDD1.n1 5.62509
R868 VDD1.n12 VDD1.n8 5.62509
R869 VDD1.n6 VDD1.n0 1.16414
R870 VDD1.n13 VDD1.n7 1.16414
R871 VDD1.n4 VDD1.n3 0.388379
R872 VDD1.n11 VDD1.n10 0.388379
R873 VDD1 VDD1.n17 0.190155
C0 VTAIL VP 1.2828f
C1 VDD2 VTAIL 3.17271f
C2 VDD1 VTAIL 3.13211f
C3 VN VP 3.33641f
C4 VN VDD2 1.02183f
C5 VDD1 VN 0.154895f
C6 VDD2 VP 0.313669f
C7 VDD1 VDD2 0.752107f
C8 VDD1 VP 1.17868f
C9 VN VTAIL 1.26862f
C10 VDD2 B 2.660418f
C11 VDD1 B 2.743344f
C12 VTAIL B 2.506894f
C13 VN B 6.235289f
C14 VP B 5.294965f
C15 VDD1.n0 B 0.023322f
C16 VDD1.n1 B 0.054683f
C17 VDD1.t3 B 0.038654f
C18 VDD1.n2 B 0.04034f
C19 VDD1.n3 B 0.011144f
C20 VDD1.n4 B 0.009046f
C21 VDD1.n5 B 0.107822f
C22 VDD1.n6 B 0.038406f
C23 VDD1.n7 B 0.023322f
C24 VDD1.n8 B 0.054683f
C25 VDD1.t2 B 0.038654f
C26 VDD1.n9 B 0.04034f
C27 VDD1.n10 B 0.011144f
C28 VDD1.n11 B 0.009046f
C29 VDD1.n12 B 0.107822f
C30 VDD1.n13 B 0.03817f
C31 VDD1.t4 B 0.025143f
C32 VDD1.t1 B 0.025143f
C33 VDD1.n14 B 0.161903f
C34 VDD1.n15 B 0.921428f
C35 VDD1.t5 B 0.025143f
C36 VDD1.t0 B 0.025143f
C37 VDD1.n16 B 0.161545f
C38 VDD1.n17 B 0.976684f
C39 VP.n0 B 0.037476f
C40 VP.t1 B 0.100468f
C41 VP.t3 B 0.13575f
C42 VP.n1 B 0.099128f
C43 VP.n2 B 0.123267f
C44 VP.t5 B 0.13575f
C45 VP.t0 B 0.100468f
C46 VP.t2 B 0.148438f
C47 VP.n3 B 0.096727f
C48 VP.n4 B 0.09064f
C49 VP.n5 B 0.033879f
C50 VP.n6 B 0.099128f
C51 VP.n7 B 0.806914f
C52 VP.n8 B 0.836491f
C53 VP.n9 B 0.037476f
C54 VP.n10 B 0.033879f
C55 VP.n11 B 0.066503f
C56 VP.n12 B 0.033879f
C57 VP.t4 B 0.13575f
C58 VP.n13 B 0.099128f
C59 VP.n14 B 0.026303f
C60 VDD2.n0 B 0.024566f
C61 VDD2.n1 B 0.057602f
C62 VDD2.t1 B 0.040717f
C63 VDD2.n2 B 0.042493f
C64 VDD2.n3 B 0.011739f
C65 VDD2.n4 B 0.009529f
C66 VDD2.n5 B 0.113578f
C67 VDD2.n6 B 0.040208f
C68 VDD2.t3 B 0.026485f
C69 VDD2.t0 B 0.026485f
C70 VDD2.n7 B 0.170547f
C71 VDD2.n8 B 0.917989f
C72 VDD2.n9 B 0.024566f
C73 VDD2.n10 B 0.057602f
C74 VDD2.t5 B 0.040717f
C75 VDD2.n11 B 0.042493f
C76 VDD2.n12 B 0.011739f
C77 VDD2.n13 B 0.009529f
C78 VDD2.n14 B 0.113578f
C79 VDD2.n15 B 0.03922f
C80 VDD2.n16 B 0.897241f
C81 VDD2.t4 B 0.026485f
C82 VDD2.t2 B 0.026485f
C83 VDD2.n17 B 0.170538f
C84 VTAIL.t6 B 0.033141f
C85 VTAIL.t7 B 0.033141f
C86 VTAIL.n0 B 0.183245f
C87 VTAIL.n1 B 0.249316f
C88 VTAIL.n2 B 0.03074f
C89 VTAIL.n3 B 0.072079f
C90 VTAIL.t2 B 0.05095f
C91 VTAIL.n4 B 0.053172f
C92 VTAIL.n5 B 0.01469f
C93 VTAIL.n6 B 0.011924f
C94 VTAIL.n7 B 0.142122f
C95 VTAIL.n8 B 0.033798f
C96 VTAIL.n9 B 0.162473f
C97 VTAIL.t1 B 0.033141f
C98 VTAIL.t4 B 0.033141f
C99 VTAIL.n10 B 0.183245f
C100 VTAIL.n11 B 0.788967f
C101 VTAIL.t11 B 0.033141f
C102 VTAIL.t10 B 0.033141f
C103 VTAIL.n12 B 0.183246f
C104 VTAIL.n13 B 0.788966f
C105 VTAIL.n14 B 0.03074f
C106 VTAIL.n15 B 0.072079f
C107 VTAIL.t8 B 0.05095f
C108 VTAIL.n16 B 0.053172f
C109 VTAIL.n17 B 0.01469f
C110 VTAIL.n18 B 0.011924f
C111 VTAIL.n19 B 0.142122f
C112 VTAIL.n20 B 0.033798f
C113 VTAIL.n21 B 0.162473f
C114 VTAIL.t0 B 0.033141f
C115 VTAIL.t5 B 0.033141f
C116 VTAIL.n22 B 0.183246f
C117 VTAIL.n23 B 0.298317f
C118 VTAIL.n24 B 0.03074f
C119 VTAIL.n25 B 0.072079f
C120 VTAIL.t3 B 0.05095f
C121 VTAIL.n26 B 0.053172f
C122 VTAIL.n27 B 0.01469f
C123 VTAIL.n28 B 0.011924f
C124 VTAIL.n29 B 0.142122f
C125 VTAIL.n30 B 0.033798f
C126 VTAIL.n31 B 0.582238f
C127 VTAIL.n32 B 0.03074f
C128 VTAIL.n33 B 0.072079f
C129 VTAIL.t9 B 0.05095f
C130 VTAIL.n34 B 0.053172f
C131 VTAIL.n35 B 0.01469f
C132 VTAIL.n36 B 0.011924f
C133 VTAIL.n37 B 0.142122f
C134 VTAIL.n38 B 0.033798f
C135 VTAIL.n39 B 0.560357f
C136 VN.n0 B 0.121809f
C137 VN.t2 B 0.09928f
C138 VN.t4 B 0.146683f
C139 VN.n1 B 0.095583f
C140 VN.n2 B 0.089568f
C141 VN.n3 B 0.033479f
C142 VN.t5 B 0.134146f
C143 VN.n4 B 0.097956f
C144 VN.n5 B 0.025992f
C145 VN.n6 B 0.121809f
C146 VN.t1 B 0.09928f
C147 VN.t3 B 0.146683f
C148 VN.n7 B 0.095583f
C149 VN.n8 B 0.089568f
C150 VN.n9 B 0.033479f
C151 VN.t0 B 0.134146f
C152 VN.n10 B 0.097956f
C153 VN.n11 B 0.813579f
.ends

