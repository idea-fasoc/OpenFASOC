* NGSPICE file created from diff_pair_sample_0627.ext - technology: sky130A

.subckt diff_pair_sample_0627 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t6 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=0.99
X1 B.t11 B.t9 B.t10 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=0.99
X2 VTAIL.t1 VN.t0 VDD2.t3 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=0.99
X3 VTAIL.t2 VN.t1 VDD2.t2 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=0.99
X4 B.t8 B.t6 B.t7 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=0.99
X5 VDD1.t2 VP.t1 VTAIL.t7 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=0.99
X6 VTAIL.t5 VP.t2 VDD1.t1 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=0.99
X7 VDD2.t1 VN.t2 VTAIL.t0 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=0.99
X8 VDD2.t0 VN.t3 VTAIL.t3 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=2.57565 pd=15.94 as=6.0879 ps=32 w=15.61 l=0.99
X9 B.t5 B.t3 B.t4 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=0.99
X10 VTAIL.t4 VP.t3 VDD1.t0 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=2.57565 ps=15.94 w=15.61 l=0.99
X11 B.t2 B.t0 B.t1 w_n1762_n4090# sky130_fd_pr__pfet_01v8 ad=6.0879 pd=32 as=0 ps=0 w=15.61 l=0.99
R0 VP.n0 VP.t2 438.531
R1 VP.n0 VP.t0 438.445
R2 VP.n2 VP.t3 419.925
R3 VP.n3 VP.t1 419.925
R4 VP.n4 VP.n3 80.6037
R5 VP.n2 VP.n1 80.6037
R6 VP.n1 VP.n0 75.3592
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.380177
R9 VP VP.n4 0.146778
R10 VTAIL.n682 VTAIL.n602 756.745
R11 VTAIL.n80 VTAIL.n0 756.745
R12 VTAIL.n166 VTAIL.n86 756.745
R13 VTAIL.n252 VTAIL.n172 756.745
R14 VTAIL.n596 VTAIL.n516 756.745
R15 VTAIL.n510 VTAIL.n430 756.745
R16 VTAIL.n424 VTAIL.n344 756.745
R17 VTAIL.n338 VTAIL.n258 756.745
R18 VTAIL.n631 VTAIL.n630 585
R19 VTAIL.n633 VTAIL.n632 585
R20 VTAIL.n626 VTAIL.n625 585
R21 VTAIL.n639 VTAIL.n638 585
R22 VTAIL.n641 VTAIL.n640 585
R23 VTAIL.n622 VTAIL.n621 585
R24 VTAIL.n648 VTAIL.n647 585
R25 VTAIL.n649 VTAIL.n620 585
R26 VTAIL.n651 VTAIL.n650 585
R27 VTAIL.n618 VTAIL.n617 585
R28 VTAIL.n657 VTAIL.n656 585
R29 VTAIL.n659 VTAIL.n658 585
R30 VTAIL.n614 VTAIL.n613 585
R31 VTAIL.n665 VTAIL.n664 585
R32 VTAIL.n667 VTAIL.n666 585
R33 VTAIL.n610 VTAIL.n609 585
R34 VTAIL.n673 VTAIL.n672 585
R35 VTAIL.n675 VTAIL.n674 585
R36 VTAIL.n606 VTAIL.n605 585
R37 VTAIL.n681 VTAIL.n680 585
R38 VTAIL.n683 VTAIL.n682 585
R39 VTAIL.n29 VTAIL.n28 585
R40 VTAIL.n31 VTAIL.n30 585
R41 VTAIL.n24 VTAIL.n23 585
R42 VTAIL.n37 VTAIL.n36 585
R43 VTAIL.n39 VTAIL.n38 585
R44 VTAIL.n20 VTAIL.n19 585
R45 VTAIL.n46 VTAIL.n45 585
R46 VTAIL.n47 VTAIL.n18 585
R47 VTAIL.n49 VTAIL.n48 585
R48 VTAIL.n16 VTAIL.n15 585
R49 VTAIL.n55 VTAIL.n54 585
R50 VTAIL.n57 VTAIL.n56 585
R51 VTAIL.n12 VTAIL.n11 585
R52 VTAIL.n63 VTAIL.n62 585
R53 VTAIL.n65 VTAIL.n64 585
R54 VTAIL.n8 VTAIL.n7 585
R55 VTAIL.n71 VTAIL.n70 585
R56 VTAIL.n73 VTAIL.n72 585
R57 VTAIL.n4 VTAIL.n3 585
R58 VTAIL.n79 VTAIL.n78 585
R59 VTAIL.n81 VTAIL.n80 585
R60 VTAIL.n115 VTAIL.n114 585
R61 VTAIL.n117 VTAIL.n116 585
R62 VTAIL.n110 VTAIL.n109 585
R63 VTAIL.n123 VTAIL.n122 585
R64 VTAIL.n125 VTAIL.n124 585
R65 VTAIL.n106 VTAIL.n105 585
R66 VTAIL.n132 VTAIL.n131 585
R67 VTAIL.n133 VTAIL.n104 585
R68 VTAIL.n135 VTAIL.n134 585
R69 VTAIL.n102 VTAIL.n101 585
R70 VTAIL.n141 VTAIL.n140 585
R71 VTAIL.n143 VTAIL.n142 585
R72 VTAIL.n98 VTAIL.n97 585
R73 VTAIL.n149 VTAIL.n148 585
R74 VTAIL.n151 VTAIL.n150 585
R75 VTAIL.n94 VTAIL.n93 585
R76 VTAIL.n157 VTAIL.n156 585
R77 VTAIL.n159 VTAIL.n158 585
R78 VTAIL.n90 VTAIL.n89 585
R79 VTAIL.n165 VTAIL.n164 585
R80 VTAIL.n167 VTAIL.n166 585
R81 VTAIL.n201 VTAIL.n200 585
R82 VTAIL.n203 VTAIL.n202 585
R83 VTAIL.n196 VTAIL.n195 585
R84 VTAIL.n209 VTAIL.n208 585
R85 VTAIL.n211 VTAIL.n210 585
R86 VTAIL.n192 VTAIL.n191 585
R87 VTAIL.n218 VTAIL.n217 585
R88 VTAIL.n219 VTAIL.n190 585
R89 VTAIL.n221 VTAIL.n220 585
R90 VTAIL.n188 VTAIL.n187 585
R91 VTAIL.n227 VTAIL.n226 585
R92 VTAIL.n229 VTAIL.n228 585
R93 VTAIL.n184 VTAIL.n183 585
R94 VTAIL.n235 VTAIL.n234 585
R95 VTAIL.n237 VTAIL.n236 585
R96 VTAIL.n180 VTAIL.n179 585
R97 VTAIL.n243 VTAIL.n242 585
R98 VTAIL.n245 VTAIL.n244 585
R99 VTAIL.n176 VTAIL.n175 585
R100 VTAIL.n251 VTAIL.n250 585
R101 VTAIL.n253 VTAIL.n252 585
R102 VTAIL.n597 VTAIL.n596 585
R103 VTAIL.n595 VTAIL.n594 585
R104 VTAIL.n520 VTAIL.n519 585
R105 VTAIL.n589 VTAIL.n588 585
R106 VTAIL.n587 VTAIL.n586 585
R107 VTAIL.n524 VTAIL.n523 585
R108 VTAIL.n581 VTAIL.n580 585
R109 VTAIL.n579 VTAIL.n578 585
R110 VTAIL.n528 VTAIL.n527 585
R111 VTAIL.n573 VTAIL.n572 585
R112 VTAIL.n571 VTAIL.n570 585
R113 VTAIL.n532 VTAIL.n531 585
R114 VTAIL.n536 VTAIL.n534 585
R115 VTAIL.n565 VTAIL.n564 585
R116 VTAIL.n563 VTAIL.n562 585
R117 VTAIL.n538 VTAIL.n537 585
R118 VTAIL.n557 VTAIL.n556 585
R119 VTAIL.n555 VTAIL.n554 585
R120 VTAIL.n542 VTAIL.n541 585
R121 VTAIL.n549 VTAIL.n548 585
R122 VTAIL.n547 VTAIL.n546 585
R123 VTAIL.n511 VTAIL.n510 585
R124 VTAIL.n509 VTAIL.n508 585
R125 VTAIL.n434 VTAIL.n433 585
R126 VTAIL.n503 VTAIL.n502 585
R127 VTAIL.n501 VTAIL.n500 585
R128 VTAIL.n438 VTAIL.n437 585
R129 VTAIL.n495 VTAIL.n494 585
R130 VTAIL.n493 VTAIL.n492 585
R131 VTAIL.n442 VTAIL.n441 585
R132 VTAIL.n487 VTAIL.n486 585
R133 VTAIL.n485 VTAIL.n484 585
R134 VTAIL.n446 VTAIL.n445 585
R135 VTAIL.n450 VTAIL.n448 585
R136 VTAIL.n479 VTAIL.n478 585
R137 VTAIL.n477 VTAIL.n476 585
R138 VTAIL.n452 VTAIL.n451 585
R139 VTAIL.n471 VTAIL.n470 585
R140 VTAIL.n469 VTAIL.n468 585
R141 VTAIL.n456 VTAIL.n455 585
R142 VTAIL.n463 VTAIL.n462 585
R143 VTAIL.n461 VTAIL.n460 585
R144 VTAIL.n425 VTAIL.n424 585
R145 VTAIL.n423 VTAIL.n422 585
R146 VTAIL.n348 VTAIL.n347 585
R147 VTAIL.n417 VTAIL.n416 585
R148 VTAIL.n415 VTAIL.n414 585
R149 VTAIL.n352 VTAIL.n351 585
R150 VTAIL.n409 VTAIL.n408 585
R151 VTAIL.n407 VTAIL.n406 585
R152 VTAIL.n356 VTAIL.n355 585
R153 VTAIL.n401 VTAIL.n400 585
R154 VTAIL.n399 VTAIL.n398 585
R155 VTAIL.n360 VTAIL.n359 585
R156 VTAIL.n364 VTAIL.n362 585
R157 VTAIL.n393 VTAIL.n392 585
R158 VTAIL.n391 VTAIL.n390 585
R159 VTAIL.n366 VTAIL.n365 585
R160 VTAIL.n385 VTAIL.n384 585
R161 VTAIL.n383 VTAIL.n382 585
R162 VTAIL.n370 VTAIL.n369 585
R163 VTAIL.n377 VTAIL.n376 585
R164 VTAIL.n375 VTAIL.n374 585
R165 VTAIL.n339 VTAIL.n338 585
R166 VTAIL.n337 VTAIL.n336 585
R167 VTAIL.n262 VTAIL.n261 585
R168 VTAIL.n331 VTAIL.n330 585
R169 VTAIL.n329 VTAIL.n328 585
R170 VTAIL.n266 VTAIL.n265 585
R171 VTAIL.n323 VTAIL.n322 585
R172 VTAIL.n321 VTAIL.n320 585
R173 VTAIL.n270 VTAIL.n269 585
R174 VTAIL.n315 VTAIL.n314 585
R175 VTAIL.n313 VTAIL.n312 585
R176 VTAIL.n274 VTAIL.n273 585
R177 VTAIL.n278 VTAIL.n276 585
R178 VTAIL.n307 VTAIL.n306 585
R179 VTAIL.n305 VTAIL.n304 585
R180 VTAIL.n280 VTAIL.n279 585
R181 VTAIL.n299 VTAIL.n298 585
R182 VTAIL.n297 VTAIL.n296 585
R183 VTAIL.n284 VTAIL.n283 585
R184 VTAIL.n291 VTAIL.n290 585
R185 VTAIL.n289 VTAIL.n288 585
R186 VTAIL.n629 VTAIL.t3 329.036
R187 VTAIL.n27 VTAIL.t2 329.036
R188 VTAIL.n113 VTAIL.t7 329.036
R189 VTAIL.n199 VTAIL.t4 329.036
R190 VTAIL.n545 VTAIL.t6 329.036
R191 VTAIL.n459 VTAIL.t5 329.036
R192 VTAIL.n373 VTAIL.t0 329.036
R193 VTAIL.n287 VTAIL.t1 329.036
R194 VTAIL.n632 VTAIL.n631 171.744
R195 VTAIL.n632 VTAIL.n625 171.744
R196 VTAIL.n639 VTAIL.n625 171.744
R197 VTAIL.n640 VTAIL.n639 171.744
R198 VTAIL.n640 VTAIL.n621 171.744
R199 VTAIL.n648 VTAIL.n621 171.744
R200 VTAIL.n649 VTAIL.n648 171.744
R201 VTAIL.n650 VTAIL.n649 171.744
R202 VTAIL.n650 VTAIL.n617 171.744
R203 VTAIL.n657 VTAIL.n617 171.744
R204 VTAIL.n658 VTAIL.n657 171.744
R205 VTAIL.n658 VTAIL.n613 171.744
R206 VTAIL.n665 VTAIL.n613 171.744
R207 VTAIL.n666 VTAIL.n665 171.744
R208 VTAIL.n666 VTAIL.n609 171.744
R209 VTAIL.n673 VTAIL.n609 171.744
R210 VTAIL.n674 VTAIL.n673 171.744
R211 VTAIL.n674 VTAIL.n605 171.744
R212 VTAIL.n681 VTAIL.n605 171.744
R213 VTAIL.n682 VTAIL.n681 171.744
R214 VTAIL.n30 VTAIL.n29 171.744
R215 VTAIL.n30 VTAIL.n23 171.744
R216 VTAIL.n37 VTAIL.n23 171.744
R217 VTAIL.n38 VTAIL.n37 171.744
R218 VTAIL.n38 VTAIL.n19 171.744
R219 VTAIL.n46 VTAIL.n19 171.744
R220 VTAIL.n47 VTAIL.n46 171.744
R221 VTAIL.n48 VTAIL.n47 171.744
R222 VTAIL.n48 VTAIL.n15 171.744
R223 VTAIL.n55 VTAIL.n15 171.744
R224 VTAIL.n56 VTAIL.n55 171.744
R225 VTAIL.n56 VTAIL.n11 171.744
R226 VTAIL.n63 VTAIL.n11 171.744
R227 VTAIL.n64 VTAIL.n63 171.744
R228 VTAIL.n64 VTAIL.n7 171.744
R229 VTAIL.n71 VTAIL.n7 171.744
R230 VTAIL.n72 VTAIL.n71 171.744
R231 VTAIL.n72 VTAIL.n3 171.744
R232 VTAIL.n79 VTAIL.n3 171.744
R233 VTAIL.n80 VTAIL.n79 171.744
R234 VTAIL.n116 VTAIL.n115 171.744
R235 VTAIL.n116 VTAIL.n109 171.744
R236 VTAIL.n123 VTAIL.n109 171.744
R237 VTAIL.n124 VTAIL.n123 171.744
R238 VTAIL.n124 VTAIL.n105 171.744
R239 VTAIL.n132 VTAIL.n105 171.744
R240 VTAIL.n133 VTAIL.n132 171.744
R241 VTAIL.n134 VTAIL.n133 171.744
R242 VTAIL.n134 VTAIL.n101 171.744
R243 VTAIL.n141 VTAIL.n101 171.744
R244 VTAIL.n142 VTAIL.n141 171.744
R245 VTAIL.n142 VTAIL.n97 171.744
R246 VTAIL.n149 VTAIL.n97 171.744
R247 VTAIL.n150 VTAIL.n149 171.744
R248 VTAIL.n150 VTAIL.n93 171.744
R249 VTAIL.n157 VTAIL.n93 171.744
R250 VTAIL.n158 VTAIL.n157 171.744
R251 VTAIL.n158 VTAIL.n89 171.744
R252 VTAIL.n165 VTAIL.n89 171.744
R253 VTAIL.n166 VTAIL.n165 171.744
R254 VTAIL.n202 VTAIL.n201 171.744
R255 VTAIL.n202 VTAIL.n195 171.744
R256 VTAIL.n209 VTAIL.n195 171.744
R257 VTAIL.n210 VTAIL.n209 171.744
R258 VTAIL.n210 VTAIL.n191 171.744
R259 VTAIL.n218 VTAIL.n191 171.744
R260 VTAIL.n219 VTAIL.n218 171.744
R261 VTAIL.n220 VTAIL.n219 171.744
R262 VTAIL.n220 VTAIL.n187 171.744
R263 VTAIL.n227 VTAIL.n187 171.744
R264 VTAIL.n228 VTAIL.n227 171.744
R265 VTAIL.n228 VTAIL.n183 171.744
R266 VTAIL.n235 VTAIL.n183 171.744
R267 VTAIL.n236 VTAIL.n235 171.744
R268 VTAIL.n236 VTAIL.n179 171.744
R269 VTAIL.n243 VTAIL.n179 171.744
R270 VTAIL.n244 VTAIL.n243 171.744
R271 VTAIL.n244 VTAIL.n175 171.744
R272 VTAIL.n251 VTAIL.n175 171.744
R273 VTAIL.n252 VTAIL.n251 171.744
R274 VTAIL.n596 VTAIL.n595 171.744
R275 VTAIL.n595 VTAIL.n519 171.744
R276 VTAIL.n588 VTAIL.n519 171.744
R277 VTAIL.n588 VTAIL.n587 171.744
R278 VTAIL.n587 VTAIL.n523 171.744
R279 VTAIL.n580 VTAIL.n523 171.744
R280 VTAIL.n580 VTAIL.n579 171.744
R281 VTAIL.n579 VTAIL.n527 171.744
R282 VTAIL.n572 VTAIL.n527 171.744
R283 VTAIL.n572 VTAIL.n571 171.744
R284 VTAIL.n571 VTAIL.n531 171.744
R285 VTAIL.n536 VTAIL.n531 171.744
R286 VTAIL.n564 VTAIL.n536 171.744
R287 VTAIL.n564 VTAIL.n563 171.744
R288 VTAIL.n563 VTAIL.n537 171.744
R289 VTAIL.n556 VTAIL.n537 171.744
R290 VTAIL.n556 VTAIL.n555 171.744
R291 VTAIL.n555 VTAIL.n541 171.744
R292 VTAIL.n548 VTAIL.n541 171.744
R293 VTAIL.n548 VTAIL.n547 171.744
R294 VTAIL.n510 VTAIL.n509 171.744
R295 VTAIL.n509 VTAIL.n433 171.744
R296 VTAIL.n502 VTAIL.n433 171.744
R297 VTAIL.n502 VTAIL.n501 171.744
R298 VTAIL.n501 VTAIL.n437 171.744
R299 VTAIL.n494 VTAIL.n437 171.744
R300 VTAIL.n494 VTAIL.n493 171.744
R301 VTAIL.n493 VTAIL.n441 171.744
R302 VTAIL.n486 VTAIL.n441 171.744
R303 VTAIL.n486 VTAIL.n485 171.744
R304 VTAIL.n485 VTAIL.n445 171.744
R305 VTAIL.n450 VTAIL.n445 171.744
R306 VTAIL.n478 VTAIL.n450 171.744
R307 VTAIL.n478 VTAIL.n477 171.744
R308 VTAIL.n477 VTAIL.n451 171.744
R309 VTAIL.n470 VTAIL.n451 171.744
R310 VTAIL.n470 VTAIL.n469 171.744
R311 VTAIL.n469 VTAIL.n455 171.744
R312 VTAIL.n462 VTAIL.n455 171.744
R313 VTAIL.n462 VTAIL.n461 171.744
R314 VTAIL.n424 VTAIL.n423 171.744
R315 VTAIL.n423 VTAIL.n347 171.744
R316 VTAIL.n416 VTAIL.n347 171.744
R317 VTAIL.n416 VTAIL.n415 171.744
R318 VTAIL.n415 VTAIL.n351 171.744
R319 VTAIL.n408 VTAIL.n351 171.744
R320 VTAIL.n408 VTAIL.n407 171.744
R321 VTAIL.n407 VTAIL.n355 171.744
R322 VTAIL.n400 VTAIL.n355 171.744
R323 VTAIL.n400 VTAIL.n399 171.744
R324 VTAIL.n399 VTAIL.n359 171.744
R325 VTAIL.n364 VTAIL.n359 171.744
R326 VTAIL.n392 VTAIL.n364 171.744
R327 VTAIL.n392 VTAIL.n391 171.744
R328 VTAIL.n391 VTAIL.n365 171.744
R329 VTAIL.n384 VTAIL.n365 171.744
R330 VTAIL.n384 VTAIL.n383 171.744
R331 VTAIL.n383 VTAIL.n369 171.744
R332 VTAIL.n376 VTAIL.n369 171.744
R333 VTAIL.n376 VTAIL.n375 171.744
R334 VTAIL.n338 VTAIL.n337 171.744
R335 VTAIL.n337 VTAIL.n261 171.744
R336 VTAIL.n330 VTAIL.n261 171.744
R337 VTAIL.n330 VTAIL.n329 171.744
R338 VTAIL.n329 VTAIL.n265 171.744
R339 VTAIL.n322 VTAIL.n265 171.744
R340 VTAIL.n322 VTAIL.n321 171.744
R341 VTAIL.n321 VTAIL.n269 171.744
R342 VTAIL.n314 VTAIL.n269 171.744
R343 VTAIL.n314 VTAIL.n313 171.744
R344 VTAIL.n313 VTAIL.n273 171.744
R345 VTAIL.n278 VTAIL.n273 171.744
R346 VTAIL.n306 VTAIL.n278 171.744
R347 VTAIL.n306 VTAIL.n305 171.744
R348 VTAIL.n305 VTAIL.n279 171.744
R349 VTAIL.n298 VTAIL.n279 171.744
R350 VTAIL.n298 VTAIL.n297 171.744
R351 VTAIL.n297 VTAIL.n283 171.744
R352 VTAIL.n290 VTAIL.n283 171.744
R353 VTAIL.n290 VTAIL.n289 171.744
R354 VTAIL.n631 VTAIL.t3 85.8723
R355 VTAIL.n29 VTAIL.t2 85.8723
R356 VTAIL.n115 VTAIL.t7 85.8723
R357 VTAIL.n201 VTAIL.t4 85.8723
R358 VTAIL.n547 VTAIL.t6 85.8723
R359 VTAIL.n461 VTAIL.t5 85.8723
R360 VTAIL.n375 VTAIL.t0 85.8723
R361 VTAIL.n289 VTAIL.t1 85.8723
R362 VTAIL.n687 VTAIL.n686 30.052
R363 VTAIL.n85 VTAIL.n84 30.052
R364 VTAIL.n171 VTAIL.n170 30.052
R365 VTAIL.n257 VTAIL.n256 30.052
R366 VTAIL.n601 VTAIL.n600 30.052
R367 VTAIL.n515 VTAIL.n514 30.052
R368 VTAIL.n429 VTAIL.n428 30.052
R369 VTAIL.n343 VTAIL.n342 30.052
R370 VTAIL.n687 VTAIL.n601 26.9617
R371 VTAIL.n343 VTAIL.n257 26.9617
R372 VTAIL.n651 VTAIL.n618 13.1884
R373 VTAIL.n49 VTAIL.n16 13.1884
R374 VTAIL.n135 VTAIL.n102 13.1884
R375 VTAIL.n221 VTAIL.n188 13.1884
R376 VTAIL.n534 VTAIL.n532 13.1884
R377 VTAIL.n448 VTAIL.n446 13.1884
R378 VTAIL.n362 VTAIL.n360 13.1884
R379 VTAIL.n276 VTAIL.n274 13.1884
R380 VTAIL.n652 VTAIL.n620 12.8005
R381 VTAIL.n656 VTAIL.n655 12.8005
R382 VTAIL.n50 VTAIL.n18 12.8005
R383 VTAIL.n54 VTAIL.n53 12.8005
R384 VTAIL.n136 VTAIL.n104 12.8005
R385 VTAIL.n140 VTAIL.n139 12.8005
R386 VTAIL.n222 VTAIL.n190 12.8005
R387 VTAIL.n226 VTAIL.n225 12.8005
R388 VTAIL.n570 VTAIL.n569 12.8005
R389 VTAIL.n566 VTAIL.n565 12.8005
R390 VTAIL.n484 VTAIL.n483 12.8005
R391 VTAIL.n480 VTAIL.n479 12.8005
R392 VTAIL.n398 VTAIL.n397 12.8005
R393 VTAIL.n394 VTAIL.n393 12.8005
R394 VTAIL.n312 VTAIL.n311 12.8005
R395 VTAIL.n308 VTAIL.n307 12.8005
R396 VTAIL.n647 VTAIL.n646 12.0247
R397 VTAIL.n659 VTAIL.n616 12.0247
R398 VTAIL.n45 VTAIL.n44 12.0247
R399 VTAIL.n57 VTAIL.n14 12.0247
R400 VTAIL.n131 VTAIL.n130 12.0247
R401 VTAIL.n143 VTAIL.n100 12.0247
R402 VTAIL.n217 VTAIL.n216 12.0247
R403 VTAIL.n229 VTAIL.n186 12.0247
R404 VTAIL.n573 VTAIL.n530 12.0247
R405 VTAIL.n562 VTAIL.n535 12.0247
R406 VTAIL.n487 VTAIL.n444 12.0247
R407 VTAIL.n476 VTAIL.n449 12.0247
R408 VTAIL.n401 VTAIL.n358 12.0247
R409 VTAIL.n390 VTAIL.n363 12.0247
R410 VTAIL.n315 VTAIL.n272 12.0247
R411 VTAIL.n304 VTAIL.n277 12.0247
R412 VTAIL.n645 VTAIL.n622 11.249
R413 VTAIL.n660 VTAIL.n614 11.249
R414 VTAIL.n43 VTAIL.n20 11.249
R415 VTAIL.n58 VTAIL.n12 11.249
R416 VTAIL.n129 VTAIL.n106 11.249
R417 VTAIL.n144 VTAIL.n98 11.249
R418 VTAIL.n215 VTAIL.n192 11.249
R419 VTAIL.n230 VTAIL.n184 11.249
R420 VTAIL.n574 VTAIL.n528 11.249
R421 VTAIL.n561 VTAIL.n538 11.249
R422 VTAIL.n488 VTAIL.n442 11.249
R423 VTAIL.n475 VTAIL.n452 11.249
R424 VTAIL.n402 VTAIL.n356 11.249
R425 VTAIL.n389 VTAIL.n366 11.249
R426 VTAIL.n316 VTAIL.n270 11.249
R427 VTAIL.n303 VTAIL.n280 11.249
R428 VTAIL.n630 VTAIL.n629 10.7239
R429 VTAIL.n28 VTAIL.n27 10.7239
R430 VTAIL.n114 VTAIL.n113 10.7239
R431 VTAIL.n200 VTAIL.n199 10.7239
R432 VTAIL.n546 VTAIL.n545 10.7239
R433 VTAIL.n460 VTAIL.n459 10.7239
R434 VTAIL.n374 VTAIL.n373 10.7239
R435 VTAIL.n288 VTAIL.n287 10.7239
R436 VTAIL.n642 VTAIL.n641 10.4732
R437 VTAIL.n664 VTAIL.n663 10.4732
R438 VTAIL.n40 VTAIL.n39 10.4732
R439 VTAIL.n62 VTAIL.n61 10.4732
R440 VTAIL.n126 VTAIL.n125 10.4732
R441 VTAIL.n148 VTAIL.n147 10.4732
R442 VTAIL.n212 VTAIL.n211 10.4732
R443 VTAIL.n234 VTAIL.n233 10.4732
R444 VTAIL.n578 VTAIL.n577 10.4732
R445 VTAIL.n558 VTAIL.n557 10.4732
R446 VTAIL.n492 VTAIL.n491 10.4732
R447 VTAIL.n472 VTAIL.n471 10.4732
R448 VTAIL.n406 VTAIL.n405 10.4732
R449 VTAIL.n386 VTAIL.n385 10.4732
R450 VTAIL.n320 VTAIL.n319 10.4732
R451 VTAIL.n300 VTAIL.n299 10.4732
R452 VTAIL.n638 VTAIL.n624 9.69747
R453 VTAIL.n667 VTAIL.n612 9.69747
R454 VTAIL.n686 VTAIL.n602 9.69747
R455 VTAIL.n36 VTAIL.n22 9.69747
R456 VTAIL.n65 VTAIL.n10 9.69747
R457 VTAIL.n84 VTAIL.n0 9.69747
R458 VTAIL.n122 VTAIL.n108 9.69747
R459 VTAIL.n151 VTAIL.n96 9.69747
R460 VTAIL.n170 VTAIL.n86 9.69747
R461 VTAIL.n208 VTAIL.n194 9.69747
R462 VTAIL.n237 VTAIL.n182 9.69747
R463 VTAIL.n256 VTAIL.n172 9.69747
R464 VTAIL.n600 VTAIL.n516 9.69747
R465 VTAIL.n581 VTAIL.n526 9.69747
R466 VTAIL.n554 VTAIL.n540 9.69747
R467 VTAIL.n514 VTAIL.n430 9.69747
R468 VTAIL.n495 VTAIL.n440 9.69747
R469 VTAIL.n468 VTAIL.n454 9.69747
R470 VTAIL.n428 VTAIL.n344 9.69747
R471 VTAIL.n409 VTAIL.n354 9.69747
R472 VTAIL.n382 VTAIL.n368 9.69747
R473 VTAIL.n342 VTAIL.n258 9.69747
R474 VTAIL.n323 VTAIL.n268 9.69747
R475 VTAIL.n296 VTAIL.n282 9.69747
R476 VTAIL.n686 VTAIL.n685 9.45567
R477 VTAIL.n84 VTAIL.n83 9.45567
R478 VTAIL.n170 VTAIL.n169 9.45567
R479 VTAIL.n256 VTAIL.n255 9.45567
R480 VTAIL.n600 VTAIL.n599 9.45567
R481 VTAIL.n514 VTAIL.n513 9.45567
R482 VTAIL.n428 VTAIL.n427 9.45567
R483 VTAIL.n342 VTAIL.n341 9.45567
R484 VTAIL.n677 VTAIL.n676 9.3005
R485 VTAIL.n679 VTAIL.n678 9.3005
R486 VTAIL.n604 VTAIL.n603 9.3005
R487 VTAIL.n685 VTAIL.n684 9.3005
R488 VTAIL.n671 VTAIL.n670 9.3005
R489 VTAIL.n669 VTAIL.n668 9.3005
R490 VTAIL.n612 VTAIL.n611 9.3005
R491 VTAIL.n663 VTAIL.n662 9.3005
R492 VTAIL.n661 VTAIL.n660 9.3005
R493 VTAIL.n616 VTAIL.n615 9.3005
R494 VTAIL.n655 VTAIL.n654 9.3005
R495 VTAIL.n628 VTAIL.n627 9.3005
R496 VTAIL.n635 VTAIL.n634 9.3005
R497 VTAIL.n637 VTAIL.n636 9.3005
R498 VTAIL.n624 VTAIL.n623 9.3005
R499 VTAIL.n643 VTAIL.n642 9.3005
R500 VTAIL.n645 VTAIL.n644 9.3005
R501 VTAIL.n646 VTAIL.n619 9.3005
R502 VTAIL.n653 VTAIL.n652 9.3005
R503 VTAIL.n608 VTAIL.n607 9.3005
R504 VTAIL.n75 VTAIL.n74 9.3005
R505 VTAIL.n77 VTAIL.n76 9.3005
R506 VTAIL.n2 VTAIL.n1 9.3005
R507 VTAIL.n83 VTAIL.n82 9.3005
R508 VTAIL.n69 VTAIL.n68 9.3005
R509 VTAIL.n67 VTAIL.n66 9.3005
R510 VTAIL.n10 VTAIL.n9 9.3005
R511 VTAIL.n61 VTAIL.n60 9.3005
R512 VTAIL.n59 VTAIL.n58 9.3005
R513 VTAIL.n14 VTAIL.n13 9.3005
R514 VTAIL.n53 VTAIL.n52 9.3005
R515 VTAIL.n26 VTAIL.n25 9.3005
R516 VTAIL.n33 VTAIL.n32 9.3005
R517 VTAIL.n35 VTAIL.n34 9.3005
R518 VTAIL.n22 VTAIL.n21 9.3005
R519 VTAIL.n41 VTAIL.n40 9.3005
R520 VTAIL.n43 VTAIL.n42 9.3005
R521 VTAIL.n44 VTAIL.n17 9.3005
R522 VTAIL.n51 VTAIL.n50 9.3005
R523 VTAIL.n6 VTAIL.n5 9.3005
R524 VTAIL.n161 VTAIL.n160 9.3005
R525 VTAIL.n163 VTAIL.n162 9.3005
R526 VTAIL.n88 VTAIL.n87 9.3005
R527 VTAIL.n169 VTAIL.n168 9.3005
R528 VTAIL.n155 VTAIL.n154 9.3005
R529 VTAIL.n153 VTAIL.n152 9.3005
R530 VTAIL.n96 VTAIL.n95 9.3005
R531 VTAIL.n147 VTAIL.n146 9.3005
R532 VTAIL.n145 VTAIL.n144 9.3005
R533 VTAIL.n100 VTAIL.n99 9.3005
R534 VTAIL.n139 VTAIL.n138 9.3005
R535 VTAIL.n112 VTAIL.n111 9.3005
R536 VTAIL.n119 VTAIL.n118 9.3005
R537 VTAIL.n121 VTAIL.n120 9.3005
R538 VTAIL.n108 VTAIL.n107 9.3005
R539 VTAIL.n127 VTAIL.n126 9.3005
R540 VTAIL.n129 VTAIL.n128 9.3005
R541 VTAIL.n130 VTAIL.n103 9.3005
R542 VTAIL.n137 VTAIL.n136 9.3005
R543 VTAIL.n92 VTAIL.n91 9.3005
R544 VTAIL.n247 VTAIL.n246 9.3005
R545 VTAIL.n249 VTAIL.n248 9.3005
R546 VTAIL.n174 VTAIL.n173 9.3005
R547 VTAIL.n255 VTAIL.n254 9.3005
R548 VTAIL.n241 VTAIL.n240 9.3005
R549 VTAIL.n239 VTAIL.n238 9.3005
R550 VTAIL.n182 VTAIL.n181 9.3005
R551 VTAIL.n233 VTAIL.n232 9.3005
R552 VTAIL.n231 VTAIL.n230 9.3005
R553 VTAIL.n186 VTAIL.n185 9.3005
R554 VTAIL.n225 VTAIL.n224 9.3005
R555 VTAIL.n198 VTAIL.n197 9.3005
R556 VTAIL.n205 VTAIL.n204 9.3005
R557 VTAIL.n207 VTAIL.n206 9.3005
R558 VTAIL.n194 VTAIL.n193 9.3005
R559 VTAIL.n213 VTAIL.n212 9.3005
R560 VTAIL.n215 VTAIL.n214 9.3005
R561 VTAIL.n216 VTAIL.n189 9.3005
R562 VTAIL.n223 VTAIL.n222 9.3005
R563 VTAIL.n178 VTAIL.n177 9.3005
R564 VTAIL.n518 VTAIL.n517 9.3005
R565 VTAIL.n593 VTAIL.n592 9.3005
R566 VTAIL.n591 VTAIL.n590 9.3005
R567 VTAIL.n522 VTAIL.n521 9.3005
R568 VTAIL.n585 VTAIL.n584 9.3005
R569 VTAIL.n583 VTAIL.n582 9.3005
R570 VTAIL.n526 VTAIL.n525 9.3005
R571 VTAIL.n577 VTAIL.n576 9.3005
R572 VTAIL.n575 VTAIL.n574 9.3005
R573 VTAIL.n530 VTAIL.n529 9.3005
R574 VTAIL.n569 VTAIL.n568 9.3005
R575 VTAIL.n567 VTAIL.n566 9.3005
R576 VTAIL.n535 VTAIL.n533 9.3005
R577 VTAIL.n561 VTAIL.n560 9.3005
R578 VTAIL.n559 VTAIL.n558 9.3005
R579 VTAIL.n540 VTAIL.n539 9.3005
R580 VTAIL.n553 VTAIL.n552 9.3005
R581 VTAIL.n551 VTAIL.n550 9.3005
R582 VTAIL.n544 VTAIL.n543 9.3005
R583 VTAIL.n599 VTAIL.n598 9.3005
R584 VTAIL.n458 VTAIL.n457 9.3005
R585 VTAIL.n465 VTAIL.n464 9.3005
R586 VTAIL.n467 VTAIL.n466 9.3005
R587 VTAIL.n454 VTAIL.n453 9.3005
R588 VTAIL.n473 VTAIL.n472 9.3005
R589 VTAIL.n475 VTAIL.n474 9.3005
R590 VTAIL.n449 VTAIL.n447 9.3005
R591 VTAIL.n481 VTAIL.n480 9.3005
R592 VTAIL.n507 VTAIL.n506 9.3005
R593 VTAIL.n432 VTAIL.n431 9.3005
R594 VTAIL.n513 VTAIL.n512 9.3005
R595 VTAIL.n505 VTAIL.n504 9.3005
R596 VTAIL.n436 VTAIL.n435 9.3005
R597 VTAIL.n499 VTAIL.n498 9.3005
R598 VTAIL.n497 VTAIL.n496 9.3005
R599 VTAIL.n440 VTAIL.n439 9.3005
R600 VTAIL.n491 VTAIL.n490 9.3005
R601 VTAIL.n489 VTAIL.n488 9.3005
R602 VTAIL.n444 VTAIL.n443 9.3005
R603 VTAIL.n483 VTAIL.n482 9.3005
R604 VTAIL.n372 VTAIL.n371 9.3005
R605 VTAIL.n379 VTAIL.n378 9.3005
R606 VTAIL.n381 VTAIL.n380 9.3005
R607 VTAIL.n368 VTAIL.n367 9.3005
R608 VTAIL.n387 VTAIL.n386 9.3005
R609 VTAIL.n389 VTAIL.n388 9.3005
R610 VTAIL.n363 VTAIL.n361 9.3005
R611 VTAIL.n395 VTAIL.n394 9.3005
R612 VTAIL.n421 VTAIL.n420 9.3005
R613 VTAIL.n346 VTAIL.n345 9.3005
R614 VTAIL.n427 VTAIL.n426 9.3005
R615 VTAIL.n419 VTAIL.n418 9.3005
R616 VTAIL.n350 VTAIL.n349 9.3005
R617 VTAIL.n413 VTAIL.n412 9.3005
R618 VTAIL.n411 VTAIL.n410 9.3005
R619 VTAIL.n354 VTAIL.n353 9.3005
R620 VTAIL.n405 VTAIL.n404 9.3005
R621 VTAIL.n403 VTAIL.n402 9.3005
R622 VTAIL.n358 VTAIL.n357 9.3005
R623 VTAIL.n397 VTAIL.n396 9.3005
R624 VTAIL.n286 VTAIL.n285 9.3005
R625 VTAIL.n293 VTAIL.n292 9.3005
R626 VTAIL.n295 VTAIL.n294 9.3005
R627 VTAIL.n282 VTAIL.n281 9.3005
R628 VTAIL.n301 VTAIL.n300 9.3005
R629 VTAIL.n303 VTAIL.n302 9.3005
R630 VTAIL.n277 VTAIL.n275 9.3005
R631 VTAIL.n309 VTAIL.n308 9.3005
R632 VTAIL.n335 VTAIL.n334 9.3005
R633 VTAIL.n260 VTAIL.n259 9.3005
R634 VTAIL.n341 VTAIL.n340 9.3005
R635 VTAIL.n333 VTAIL.n332 9.3005
R636 VTAIL.n264 VTAIL.n263 9.3005
R637 VTAIL.n327 VTAIL.n326 9.3005
R638 VTAIL.n325 VTAIL.n324 9.3005
R639 VTAIL.n268 VTAIL.n267 9.3005
R640 VTAIL.n319 VTAIL.n318 9.3005
R641 VTAIL.n317 VTAIL.n316 9.3005
R642 VTAIL.n272 VTAIL.n271 9.3005
R643 VTAIL.n311 VTAIL.n310 9.3005
R644 VTAIL.n637 VTAIL.n626 8.92171
R645 VTAIL.n668 VTAIL.n610 8.92171
R646 VTAIL.n684 VTAIL.n683 8.92171
R647 VTAIL.n35 VTAIL.n24 8.92171
R648 VTAIL.n66 VTAIL.n8 8.92171
R649 VTAIL.n82 VTAIL.n81 8.92171
R650 VTAIL.n121 VTAIL.n110 8.92171
R651 VTAIL.n152 VTAIL.n94 8.92171
R652 VTAIL.n168 VTAIL.n167 8.92171
R653 VTAIL.n207 VTAIL.n196 8.92171
R654 VTAIL.n238 VTAIL.n180 8.92171
R655 VTAIL.n254 VTAIL.n253 8.92171
R656 VTAIL.n598 VTAIL.n597 8.92171
R657 VTAIL.n582 VTAIL.n524 8.92171
R658 VTAIL.n553 VTAIL.n542 8.92171
R659 VTAIL.n512 VTAIL.n511 8.92171
R660 VTAIL.n496 VTAIL.n438 8.92171
R661 VTAIL.n467 VTAIL.n456 8.92171
R662 VTAIL.n426 VTAIL.n425 8.92171
R663 VTAIL.n410 VTAIL.n352 8.92171
R664 VTAIL.n381 VTAIL.n370 8.92171
R665 VTAIL.n340 VTAIL.n339 8.92171
R666 VTAIL.n324 VTAIL.n266 8.92171
R667 VTAIL.n295 VTAIL.n284 8.92171
R668 VTAIL.n634 VTAIL.n633 8.14595
R669 VTAIL.n672 VTAIL.n671 8.14595
R670 VTAIL.n680 VTAIL.n604 8.14595
R671 VTAIL.n32 VTAIL.n31 8.14595
R672 VTAIL.n70 VTAIL.n69 8.14595
R673 VTAIL.n78 VTAIL.n2 8.14595
R674 VTAIL.n118 VTAIL.n117 8.14595
R675 VTAIL.n156 VTAIL.n155 8.14595
R676 VTAIL.n164 VTAIL.n88 8.14595
R677 VTAIL.n204 VTAIL.n203 8.14595
R678 VTAIL.n242 VTAIL.n241 8.14595
R679 VTAIL.n250 VTAIL.n174 8.14595
R680 VTAIL.n594 VTAIL.n518 8.14595
R681 VTAIL.n586 VTAIL.n585 8.14595
R682 VTAIL.n550 VTAIL.n549 8.14595
R683 VTAIL.n508 VTAIL.n432 8.14595
R684 VTAIL.n500 VTAIL.n499 8.14595
R685 VTAIL.n464 VTAIL.n463 8.14595
R686 VTAIL.n422 VTAIL.n346 8.14595
R687 VTAIL.n414 VTAIL.n413 8.14595
R688 VTAIL.n378 VTAIL.n377 8.14595
R689 VTAIL.n336 VTAIL.n260 8.14595
R690 VTAIL.n328 VTAIL.n327 8.14595
R691 VTAIL.n292 VTAIL.n291 8.14595
R692 VTAIL.n630 VTAIL.n628 7.3702
R693 VTAIL.n675 VTAIL.n608 7.3702
R694 VTAIL.n679 VTAIL.n606 7.3702
R695 VTAIL.n28 VTAIL.n26 7.3702
R696 VTAIL.n73 VTAIL.n6 7.3702
R697 VTAIL.n77 VTAIL.n4 7.3702
R698 VTAIL.n114 VTAIL.n112 7.3702
R699 VTAIL.n159 VTAIL.n92 7.3702
R700 VTAIL.n163 VTAIL.n90 7.3702
R701 VTAIL.n200 VTAIL.n198 7.3702
R702 VTAIL.n245 VTAIL.n178 7.3702
R703 VTAIL.n249 VTAIL.n176 7.3702
R704 VTAIL.n593 VTAIL.n520 7.3702
R705 VTAIL.n589 VTAIL.n522 7.3702
R706 VTAIL.n546 VTAIL.n544 7.3702
R707 VTAIL.n507 VTAIL.n434 7.3702
R708 VTAIL.n503 VTAIL.n436 7.3702
R709 VTAIL.n460 VTAIL.n458 7.3702
R710 VTAIL.n421 VTAIL.n348 7.3702
R711 VTAIL.n417 VTAIL.n350 7.3702
R712 VTAIL.n374 VTAIL.n372 7.3702
R713 VTAIL.n335 VTAIL.n262 7.3702
R714 VTAIL.n331 VTAIL.n264 7.3702
R715 VTAIL.n288 VTAIL.n286 7.3702
R716 VTAIL.n676 VTAIL.n675 6.59444
R717 VTAIL.n676 VTAIL.n606 6.59444
R718 VTAIL.n74 VTAIL.n73 6.59444
R719 VTAIL.n74 VTAIL.n4 6.59444
R720 VTAIL.n160 VTAIL.n159 6.59444
R721 VTAIL.n160 VTAIL.n90 6.59444
R722 VTAIL.n246 VTAIL.n245 6.59444
R723 VTAIL.n246 VTAIL.n176 6.59444
R724 VTAIL.n590 VTAIL.n520 6.59444
R725 VTAIL.n590 VTAIL.n589 6.59444
R726 VTAIL.n504 VTAIL.n434 6.59444
R727 VTAIL.n504 VTAIL.n503 6.59444
R728 VTAIL.n418 VTAIL.n348 6.59444
R729 VTAIL.n418 VTAIL.n417 6.59444
R730 VTAIL.n332 VTAIL.n262 6.59444
R731 VTAIL.n332 VTAIL.n331 6.59444
R732 VTAIL.n633 VTAIL.n628 5.81868
R733 VTAIL.n672 VTAIL.n608 5.81868
R734 VTAIL.n680 VTAIL.n679 5.81868
R735 VTAIL.n31 VTAIL.n26 5.81868
R736 VTAIL.n70 VTAIL.n6 5.81868
R737 VTAIL.n78 VTAIL.n77 5.81868
R738 VTAIL.n117 VTAIL.n112 5.81868
R739 VTAIL.n156 VTAIL.n92 5.81868
R740 VTAIL.n164 VTAIL.n163 5.81868
R741 VTAIL.n203 VTAIL.n198 5.81868
R742 VTAIL.n242 VTAIL.n178 5.81868
R743 VTAIL.n250 VTAIL.n249 5.81868
R744 VTAIL.n594 VTAIL.n593 5.81868
R745 VTAIL.n586 VTAIL.n522 5.81868
R746 VTAIL.n549 VTAIL.n544 5.81868
R747 VTAIL.n508 VTAIL.n507 5.81868
R748 VTAIL.n500 VTAIL.n436 5.81868
R749 VTAIL.n463 VTAIL.n458 5.81868
R750 VTAIL.n422 VTAIL.n421 5.81868
R751 VTAIL.n414 VTAIL.n350 5.81868
R752 VTAIL.n377 VTAIL.n372 5.81868
R753 VTAIL.n336 VTAIL.n335 5.81868
R754 VTAIL.n328 VTAIL.n264 5.81868
R755 VTAIL.n291 VTAIL.n286 5.81868
R756 VTAIL.n634 VTAIL.n626 5.04292
R757 VTAIL.n671 VTAIL.n610 5.04292
R758 VTAIL.n683 VTAIL.n604 5.04292
R759 VTAIL.n32 VTAIL.n24 5.04292
R760 VTAIL.n69 VTAIL.n8 5.04292
R761 VTAIL.n81 VTAIL.n2 5.04292
R762 VTAIL.n118 VTAIL.n110 5.04292
R763 VTAIL.n155 VTAIL.n94 5.04292
R764 VTAIL.n167 VTAIL.n88 5.04292
R765 VTAIL.n204 VTAIL.n196 5.04292
R766 VTAIL.n241 VTAIL.n180 5.04292
R767 VTAIL.n253 VTAIL.n174 5.04292
R768 VTAIL.n597 VTAIL.n518 5.04292
R769 VTAIL.n585 VTAIL.n524 5.04292
R770 VTAIL.n550 VTAIL.n542 5.04292
R771 VTAIL.n511 VTAIL.n432 5.04292
R772 VTAIL.n499 VTAIL.n438 5.04292
R773 VTAIL.n464 VTAIL.n456 5.04292
R774 VTAIL.n425 VTAIL.n346 5.04292
R775 VTAIL.n413 VTAIL.n352 5.04292
R776 VTAIL.n378 VTAIL.n370 5.04292
R777 VTAIL.n339 VTAIL.n260 5.04292
R778 VTAIL.n327 VTAIL.n266 5.04292
R779 VTAIL.n292 VTAIL.n284 5.04292
R780 VTAIL.n638 VTAIL.n637 4.26717
R781 VTAIL.n668 VTAIL.n667 4.26717
R782 VTAIL.n684 VTAIL.n602 4.26717
R783 VTAIL.n36 VTAIL.n35 4.26717
R784 VTAIL.n66 VTAIL.n65 4.26717
R785 VTAIL.n82 VTAIL.n0 4.26717
R786 VTAIL.n122 VTAIL.n121 4.26717
R787 VTAIL.n152 VTAIL.n151 4.26717
R788 VTAIL.n168 VTAIL.n86 4.26717
R789 VTAIL.n208 VTAIL.n207 4.26717
R790 VTAIL.n238 VTAIL.n237 4.26717
R791 VTAIL.n254 VTAIL.n172 4.26717
R792 VTAIL.n598 VTAIL.n516 4.26717
R793 VTAIL.n582 VTAIL.n581 4.26717
R794 VTAIL.n554 VTAIL.n553 4.26717
R795 VTAIL.n512 VTAIL.n430 4.26717
R796 VTAIL.n496 VTAIL.n495 4.26717
R797 VTAIL.n468 VTAIL.n467 4.26717
R798 VTAIL.n426 VTAIL.n344 4.26717
R799 VTAIL.n410 VTAIL.n409 4.26717
R800 VTAIL.n382 VTAIL.n381 4.26717
R801 VTAIL.n340 VTAIL.n258 4.26717
R802 VTAIL.n324 VTAIL.n323 4.26717
R803 VTAIL.n296 VTAIL.n295 4.26717
R804 VTAIL.n641 VTAIL.n624 3.49141
R805 VTAIL.n664 VTAIL.n612 3.49141
R806 VTAIL.n39 VTAIL.n22 3.49141
R807 VTAIL.n62 VTAIL.n10 3.49141
R808 VTAIL.n125 VTAIL.n108 3.49141
R809 VTAIL.n148 VTAIL.n96 3.49141
R810 VTAIL.n211 VTAIL.n194 3.49141
R811 VTAIL.n234 VTAIL.n182 3.49141
R812 VTAIL.n578 VTAIL.n526 3.49141
R813 VTAIL.n557 VTAIL.n540 3.49141
R814 VTAIL.n492 VTAIL.n440 3.49141
R815 VTAIL.n471 VTAIL.n454 3.49141
R816 VTAIL.n406 VTAIL.n354 3.49141
R817 VTAIL.n385 VTAIL.n368 3.49141
R818 VTAIL.n320 VTAIL.n268 3.49141
R819 VTAIL.n299 VTAIL.n282 3.49141
R820 VTAIL.n642 VTAIL.n622 2.71565
R821 VTAIL.n663 VTAIL.n614 2.71565
R822 VTAIL.n40 VTAIL.n20 2.71565
R823 VTAIL.n61 VTAIL.n12 2.71565
R824 VTAIL.n126 VTAIL.n106 2.71565
R825 VTAIL.n147 VTAIL.n98 2.71565
R826 VTAIL.n212 VTAIL.n192 2.71565
R827 VTAIL.n233 VTAIL.n184 2.71565
R828 VTAIL.n577 VTAIL.n528 2.71565
R829 VTAIL.n558 VTAIL.n538 2.71565
R830 VTAIL.n491 VTAIL.n442 2.71565
R831 VTAIL.n472 VTAIL.n452 2.71565
R832 VTAIL.n405 VTAIL.n356 2.71565
R833 VTAIL.n386 VTAIL.n366 2.71565
R834 VTAIL.n319 VTAIL.n270 2.71565
R835 VTAIL.n300 VTAIL.n280 2.71565
R836 VTAIL.n629 VTAIL.n627 2.41282
R837 VTAIL.n27 VTAIL.n25 2.41282
R838 VTAIL.n113 VTAIL.n111 2.41282
R839 VTAIL.n199 VTAIL.n197 2.41282
R840 VTAIL.n545 VTAIL.n543 2.41282
R841 VTAIL.n459 VTAIL.n457 2.41282
R842 VTAIL.n373 VTAIL.n371 2.41282
R843 VTAIL.n287 VTAIL.n285 2.41282
R844 VTAIL.n647 VTAIL.n645 1.93989
R845 VTAIL.n660 VTAIL.n659 1.93989
R846 VTAIL.n45 VTAIL.n43 1.93989
R847 VTAIL.n58 VTAIL.n57 1.93989
R848 VTAIL.n131 VTAIL.n129 1.93989
R849 VTAIL.n144 VTAIL.n143 1.93989
R850 VTAIL.n217 VTAIL.n215 1.93989
R851 VTAIL.n230 VTAIL.n229 1.93989
R852 VTAIL.n574 VTAIL.n573 1.93989
R853 VTAIL.n562 VTAIL.n561 1.93989
R854 VTAIL.n488 VTAIL.n487 1.93989
R855 VTAIL.n476 VTAIL.n475 1.93989
R856 VTAIL.n402 VTAIL.n401 1.93989
R857 VTAIL.n390 VTAIL.n389 1.93989
R858 VTAIL.n316 VTAIL.n315 1.93989
R859 VTAIL.n304 VTAIL.n303 1.93989
R860 VTAIL.n646 VTAIL.n620 1.16414
R861 VTAIL.n656 VTAIL.n616 1.16414
R862 VTAIL.n44 VTAIL.n18 1.16414
R863 VTAIL.n54 VTAIL.n14 1.16414
R864 VTAIL.n130 VTAIL.n104 1.16414
R865 VTAIL.n140 VTAIL.n100 1.16414
R866 VTAIL.n216 VTAIL.n190 1.16414
R867 VTAIL.n226 VTAIL.n186 1.16414
R868 VTAIL.n570 VTAIL.n530 1.16414
R869 VTAIL.n565 VTAIL.n535 1.16414
R870 VTAIL.n484 VTAIL.n444 1.16414
R871 VTAIL.n479 VTAIL.n449 1.16414
R872 VTAIL.n398 VTAIL.n358 1.16414
R873 VTAIL.n393 VTAIL.n363 1.16414
R874 VTAIL.n312 VTAIL.n272 1.16414
R875 VTAIL.n307 VTAIL.n277 1.16414
R876 VTAIL.n429 VTAIL.n343 1.13843
R877 VTAIL.n601 VTAIL.n515 1.13843
R878 VTAIL.n257 VTAIL.n171 1.13843
R879 VTAIL VTAIL.n85 0.627655
R880 VTAIL VTAIL.n687 0.511276
R881 VTAIL.n515 VTAIL.n429 0.470328
R882 VTAIL.n171 VTAIL.n85 0.470328
R883 VTAIL.n652 VTAIL.n651 0.388379
R884 VTAIL.n655 VTAIL.n618 0.388379
R885 VTAIL.n50 VTAIL.n49 0.388379
R886 VTAIL.n53 VTAIL.n16 0.388379
R887 VTAIL.n136 VTAIL.n135 0.388379
R888 VTAIL.n139 VTAIL.n102 0.388379
R889 VTAIL.n222 VTAIL.n221 0.388379
R890 VTAIL.n225 VTAIL.n188 0.388379
R891 VTAIL.n569 VTAIL.n532 0.388379
R892 VTAIL.n566 VTAIL.n534 0.388379
R893 VTAIL.n483 VTAIL.n446 0.388379
R894 VTAIL.n480 VTAIL.n448 0.388379
R895 VTAIL.n397 VTAIL.n360 0.388379
R896 VTAIL.n394 VTAIL.n362 0.388379
R897 VTAIL.n311 VTAIL.n274 0.388379
R898 VTAIL.n308 VTAIL.n276 0.388379
R899 VTAIL.n635 VTAIL.n627 0.155672
R900 VTAIL.n636 VTAIL.n635 0.155672
R901 VTAIL.n636 VTAIL.n623 0.155672
R902 VTAIL.n643 VTAIL.n623 0.155672
R903 VTAIL.n644 VTAIL.n643 0.155672
R904 VTAIL.n644 VTAIL.n619 0.155672
R905 VTAIL.n653 VTAIL.n619 0.155672
R906 VTAIL.n654 VTAIL.n653 0.155672
R907 VTAIL.n654 VTAIL.n615 0.155672
R908 VTAIL.n661 VTAIL.n615 0.155672
R909 VTAIL.n662 VTAIL.n661 0.155672
R910 VTAIL.n662 VTAIL.n611 0.155672
R911 VTAIL.n669 VTAIL.n611 0.155672
R912 VTAIL.n670 VTAIL.n669 0.155672
R913 VTAIL.n670 VTAIL.n607 0.155672
R914 VTAIL.n677 VTAIL.n607 0.155672
R915 VTAIL.n678 VTAIL.n677 0.155672
R916 VTAIL.n678 VTAIL.n603 0.155672
R917 VTAIL.n685 VTAIL.n603 0.155672
R918 VTAIL.n33 VTAIL.n25 0.155672
R919 VTAIL.n34 VTAIL.n33 0.155672
R920 VTAIL.n34 VTAIL.n21 0.155672
R921 VTAIL.n41 VTAIL.n21 0.155672
R922 VTAIL.n42 VTAIL.n41 0.155672
R923 VTAIL.n42 VTAIL.n17 0.155672
R924 VTAIL.n51 VTAIL.n17 0.155672
R925 VTAIL.n52 VTAIL.n51 0.155672
R926 VTAIL.n52 VTAIL.n13 0.155672
R927 VTAIL.n59 VTAIL.n13 0.155672
R928 VTAIL.n60 VTAIL.n59 0.155672
R929 VTAIL.n60 VTAIL.n9 0.155672
R930 VTAIL.n67 VTAIL.n9 0.155672
R931 VTAIL.n68 VTAIL.n67 0.155672
R932 VTAIL.n68 VTAIL.n5 0.155672
R933 VTAIL.n75 VTAIL.n5 0.155672
R934 VTAIL.n76 VTAIL.n75 0.155672
R935 VTAIL.n76 VTAIL.n1 0.155672
R936 VTAIL.n83 VTAIL.n1 0.155672
R937 VTAIL.n119 VTAIL.n111 0.155672
R938 VTAIL.n120 VTAIL.n119 0.155672
R939 VTAIL.n120 VTAIL.n107 0.155672
R940 VTAIL.n127 VTAIL.n107 0.155672
R941 VTAIL.n128 VTAIL.n127 0.155672
R942 VTAIL.n128 VTAIL.n103 0.155672
R943 VTAIL.n137 VTAIL.n103 0.155672
R944 VTAIL.n138 VTAIL.n137 0.155672
R945 VTAIL.n138 VTAIL.n99 0.155672
R946 VTAIL.n145 VTAIL.n99 0.155672
R947 VTAIL.n146 VTAIL.n145 0.155672
R948 VTAIL.n146 VTAIL.n95 0.155672
R949 VTAIL.n153 VTAIL.n95 0.155672
R950 VTAIL.n154 VTAIL.n153 0.155672
R951 VTAIL.n154 VTAIL.n91 0.155672
R952 VTAIL.n161 VTAIL.n91 0.155672
R953 VTAIL.n162 VTAIL.n161 0.155672
R954 VTAIL.n162 VTAIL.n87 0.155672
R955 VTAIL.n169 VTAIL.n87 0.155672
R956 VTAIL.n205 VTAIL.n197 0.155672
R957 VTAIL.n206 VTAIL.n205 0.155672
R958 VTAIL.n206 VTAIL.n193 0.155672
R959 VTAIL.n213 VTAIL.n193 0.155672
R960 VTAIL.n214 VTAIL.n213 0.155672
R961 VTAIL.n214 VTAIL.n189 0.155672
R962 VTAIL.n223 VTAIL.n189 0.155672
R963 VTAIL.n224 VTAIL.n223 0.155672
R964 VTAIL.n224 VTAIL.n185 0.155672
R965 VTAIL.n231 VTAIL.n185 0.155672
R966 VTAIL.n232 VTAIL.n231 0.155672
R967 VTAIL.n232 VTAIL.n181 0.155672
R968 VTAIL.n239 VTAIL.n181 0.155672
R969 VTAIL.n240 VTAIL.n239 0.155672
R970 VTAIL.n240 VTAIL.n177 0.155672
R971 VTAIL.n247 VTAIL.n177 0.155672
R972 VTAIL.n248 VTAIL.n247 0.155672
R973 VTAIL.n248 VTAIL.n173 0.155672
R974 VTAIL.n255 VTAIL.n173 0.155672
R975 VTAIL.n599 VTAIL.n517 0.155672
R976 VTAIL.n592 VTAIL.n517 0.155672
R977 VTAIL.n592 VTAIL.n591 0.155672
R978 VTAIL.n591 VTAIL.n521 0.155672
R979 VTAIL.n584 VTAIL.n521 0.155672
R980 VTAIL.n584 VTAIL.n583 0.155672
R981 VTAIL.n583 VTAIL.n525 0.155672
R982 VTAIL.n576 VTAIL.n525 0.155672
R983 VTAIL.n576 VTAIL.n575 0.155672
R984 VTAIL.n575 VTAIL.n529 0.155672
R985 VTAIL.n568 VTAIL.n529 0.155672
R986 VTAIL.n568 VTAIL.n567 0.155672
R987 VTAIL.n567 VTAIL.n533 0.155672
R988 VTAIL.n560 VTAIL.n533 0.155672
R989 VTAIL.n560 VTAIL.n559 0.155672
R990 VTAIL.n559 VTAIL.n539 0.155672
R991 VTAIL.n552 VTAIL.n539 0.155672
R992 VTAIL.n552 VTAIL.n551 0.155672
R993 VTAIL.n551 VTAIL.n543 0.155672
R994 VTAIL.n513 VTAIL.n431 0.155672
R995 VTAIL.n506 VTAIL.n431 0.155672
R996 VTAIL.n506 VTAIL.n505 0.155672
R997 VTAIL.n505 VTAIL.n435 0.155672
R998 VTAIL.n498 VTAIL.n435 0.155672
R999 VTAIL.n498 VTAIL.n497 0.155672
R1000 VTAIL.n497 VTAIL.n439 0.155672
R1001 VTAIL.n490 VTAIL.n439 0.155672
R1002 VTAIL.n490 VTAIL.n489 0.155672
R1003 VTAIL.n489 VTAIL.n443 0.155672
R1004 VTAIL.n482 VTAIL.n443 0.155672
R1005 VTAIL.n482 VTAIL.n481 0.155672
R1006 VTAIL.n481 VTAIL.n447 0.155672
R1007 VTAIL.n474 VTAIL.n447 0.155672
R1008 VTAIL.n474 VTAIL.n473 0.155672
R1009 VTAIL.n473 VTAIL.n453 0.155672
R1010 VTAIL.n466 VTAIL.n453 0.155672
R1011 VTAIL.n466 VTAIL.n465 0.155672
R1012 VTAIL.n465 VTAIL.n457 0.155672
R1013 VTAIL.n427 VTAIL.n345 0.155672
R1014 VTAIL.n420 VTAIL.n345 0.155672
R1015 VTAIL.n420 VTAIL.n419 0.155672
R1016 VTAIL.n419 VTAIL.n349 0.155672
R1017 VTAIL.n412 VTAIL.n349 0.155672
R1018 VTAIL.n412 VTAIL.n411 0.155672
R1019 VTAIL.n411 VTAIL.n353 0.155672
R1020 VTAIL.n404 VTAIL.n353 0.155672
R1021 VTAIL.n404 VTAIL.n403 0.155672
R1022 VTAIL.n403 VTAIL.n357 0.155672
R1023 VTAIL.n396 VTAIL.n357 0.155672
R1024 VTAIL.n396 VTAIL.n395 0.155672
R1025 VTAIL.n395 VTAIL.n361 0.155672
R1026 VTAIL.n388 VTAIL.n361 0.155672
R1027 VTAIL.n388 VTAIL.n387 0.155672
R1028 VTAIL.n387 VTAIL.n367 0.155672
R1029 VTAIL.n380 VTAIL.n367 0.155672
R1030 VTAIL.n380 VTAIL.n379 0.155672
R1031 VTAIL.n379 VTAIL.n371 0.155672
R1032 VTAIL.n341 VTAIL.n259 0.155672
R1033 VTAIL.n334 VTAIL.n259 0.155672
R1034 VTAIL.n334 VTAIL.n333 0.155672
R1035 VTAIL.n333 VTAIL.n263 0.155672
R1036 VTAIL.n326 VTAIL.n263 0.155672
R1037 VTAIL.n326 VTAIL.n325 0.155672
R1038 VTAIL.n325 VTAIL.n267 0.155672
R1039 VTAIL.n318 VTAIL.n267 0.155672
R1040 VTAIL.n318 VTAIL.n317 0.155672
R1041 VTAIL.n317 VTAIL.n271 0.155672
R1042 VTAIL.n310 VTAIL.n271 0.155672
R1043 VTAIL.n310 VTAIL.n309 0.155672
R1044 VTAIL.n309 VTAIL.n275 0.155672
R1045 VTAIL.n302 VTAIL.n275 0.155672
R1046 VTAIL.n302 VTAIL.n301 0.155672
R1047 VTAIL.n301 VTAIL.n281 0.155672
R1048 VTAIL.n294 VTAIL.n281 0.155672
R1049 VTAIL.n294 VTAIL.n293 0.155672
R1050 VTAIL.n293 VTAIL.n285 0.155672
R1051 VDD1 VDD1.n1 109.516
R1052 VDD1 VDD1.n0 68.4639
R1053 VDD1.n0 VDD1.t1 2.08282
R1054 VDD1.n0 VDD1.t3 2.08282
R1055 VDD1.n1 VDD1.t0 2.08282
R1056 VDD1.n1 VDD1.t2 2.08282
R1057 B.n363 B.n362 585
R1058 B.n361 B.n94 585
R1059 B.n360 B.n359 585
R1060 B.n358 B.n95 585
R1061 B.n357 B.n356 585
R1062 B.n355 B.n96 585
R1063 B.n354 B.n353 585
R1064 B.n352 B.n97 585
R1065 B.n351 B.n350 585
R1066 B.n349 B.n98 585
R1067 B.n348 B.n347 585
R1068 B.n346 B.n99 585
R1069 B.n345 B.n344 585
R1070 B.n343 B.n100 585
R1071 B.n342 B.n341 585
R1072 B.n340 B.n101 585
R1073 B.n339 B.n338 585
R1074 B.n337 B.n102 585
R1075 B.n336 B.n335 585
R1076 B.n334 B.n103 585
R1077 B.n333 B.n332 585
R1078 B.n331 B.n104 585
R1079 B.n330 B.n329 585
R1080 B.n328 B.n105 585
R1081 B.n327 B.n326 585
R1082 B.n325 B.n106 585
R1083 B.n324 B.n323 585
R1084 B.n322 B.n107 585
R1085 B.n321 B.n320 585
R1086 B.n319 B.n108 585
R1087 B.n318 B.n317 585
R1088 B.n316 B.n109 585
R1089 B.n315 B.n314 585
R1090 B.n313 B.n110 585
R1091 B.n312 B.n311 585
R1092 B.n310 B.n111 585
R1093 B.n309 B.n308 585
R1094 B.n307 B.n112 585
R1095 B.n306 B.n305 585
R1096 B.n304 B.n113 585
R1097 B.n303 B.n302 585
R1098 B.n301 B.n114 585
R1099 B.n300 B.n299 585
R1100 B.n298 B.n115 585
R1101 B.n297 B.n296 585
R1102 B.n295 B.n116 585
R1103 B.n294 B.n293 585
R1104 B.n292 B.n117 585
R1105 B.n291 B.n290 585
R1106 B.n289 B.n118 585
R1107 B.n288 B.n287 585
R1108 B.n286 B.n119 585
R1109 B.n285 B.n284 585
R1110 B.n280 B.n120 585
R1111 B.n279 B.n278 585
R1112 B.n277 B.n121 585
R1113 B.n276 B.n275 585
R1114 B.n274 B.n122 585
R1115 B.n273 B.n272 585
R1116 B.n271 B.n123 585
R1117 B.n270 B.n269 585
R1118 B.n268 B.n124 585
R1119 B.n266 B.n265 585
R1120 B.n264 B.n127 585
R1121 B.n263 B.n262 585
R1122 B.n261 B.n128 585
R1123 B.n260 B.n259 585
R1124 B.n258 B.n129 585
R1125 B.n257 B.n256 585
R1126 B.n255 B.n130 585
R1127 B.n254 B.n253 585
R1128 B.n252 B.n131 585
R1129 B.n251 B.n250 585
R1130 B.n249 B.n132 585
R1131 B.n248 B.n247 585
R1132 B.n246 B.n133 585
R1133 B.n245 B.n244 585
R1134 B.n243 B.n134 585
R1135 B.n242 B.n241 585
R1136 B.n240 B.n135 585
R1137 B.n239 B.n238 585
R1138 B.n237 B.n136 585
R1139 B.n236 B.n235 585
R1140 B.n234 B.n137 585
R1141 B.n233 B.n232 585
R1142 B.n231 B.n138 585
R1143 B.n230 B.n229 585
R1144 B.n228 B.n139 585
R1145 B.n227 B.n226 585
R1146 B.n225 B.n140 585
R1147 B.n224 B.n223 585
R1148 B.n222 B.n141 585
R1149 B.n221 B.n220 585
R1150 B.n219 B.n142 585
R1151 B.n218 B.n217 585
R1152 B.n216 B.n143 585
R1153 B.n215 B.n214 585
R1154 B.n213 B.n144 585
R1155 B.n212 B.n211 585
R1156 B.n210 B.n145 585
R1157 B.n209 B.n208 585
R1158 B.n207 B.n146 585
R1159 B.n206 B.n205 585
R1160 B.n204 B.n147 585
R1161 B.n203 B.n202 585
R1162 B.n201 B.n148 585
R1163 B.n200 B.n199 585
R1164 B.n198 B.n149 585
R1165 B.n197 B.n196 585
R1166 B.n195 B.n150 585
R1167 B.n194 B.n193 585
R1168 B.n192 B.n151 585
R1169 B.n191 B.n190 585
R1170 B.n189 B.n152 585
R1171 B.n364 B.n93 585
R1172 B.n366 B.n365 585
R1173 B.n367 B.n92 585
R1174 B.n369 B.n368 585
R1175 B.n370 B.n91 585
R1176 B.n372 B.n371 585
R1177 B.n373 B.n90 585
R1178 B.n375 B.n374 585
R1179 B.n376 B.n89 585
R1180 B.n378 B.n377 585
R1181 B.n379 B.n88 585
R1182 B.n381 B.n380 585
R1183 B.n382 B.n87 585
R1184 B.n384 B.n383 585
R1185 B.n385 B.n86 585
R1186 B.n387 B.n386 585
R1187 B.n388 B.n85 585
R1188 B.n390 B.n389 585
R1189 B.n391 B.n84 585
R1190 B.n393 B.n392 585
R1191 B.n394 B.n83 585
R1192 B.n396 B.n395 585
R1193 B.n397 B.n82 585
R1194 B.n399 B.n398 585
R1195 B.n400 B.n81 585
R1196 B.n402 B.n401 585
R1197 B.n403 B.n80 585
R1198 B.n405 B.n404 585
R1199 B.n406 B.n79 585
R1200 B.n408 B.n407 585
R1201 B.n409 B.n78 585
R1202 B.n411 B.n410 585
R1203 B.n412 B.n77 585
R1204 B.n414 B.n413 585
R1205 B.n415 B.n76 585
R1206 B.n417 B.n416 585
R1207 B.n418 B.n75 585
R1208 B.n420 B.n419 585
R1209 B.n421 B.n74 585
R1210 B.n423 B.n422 585
R1211 B.n595 B.n594 585
R1212 B.n593 B.n12 585
R1213 B.n592 B.n591 585
R1214 B.n590 B.n13 585
R1215 B.n589 B.n588 585
R1216 B.n587 B.n14 585
R1217 B.n586 B.n585 585
R1218 B.n584 B.n15 585
R1219 B.n583 B.n582 585
R1220 B.n581 B.n16 585
R1221 B.n580 B.n579 585
R1222 B.n578 B.n17 585
R1223 B.n577 B.n576 585
R1224 B.n575 B.n18 585
R1225 B.n574 B.n573 585
R1226 B.n572 B.n19 585
R1227 B.n571 B.n570 585
R1228 B.n569 B.n20 585
R1229 B.n568 B.n567 585
R1230 B.n566 B.n21 585
R1231 B.n565 B.n564 585
R1232 B.n563 B.n22 585
R1233 B.n562 B.n561 585
R1234 B.n560 B.n23 585
R1235 B.n559 B.n558 585
R1236 B.n557 B.n24 585
R1237 B.n556 B.n555 585
R1238 B.n554 B.n25 585
R1239 B.n553 B.n552 585
R1240 B.n551 B.n26 585
R1241 B.n550 B.n549 585
R1242 B.n548 B.n27 585
R1243 B.n547 B.n546 585
R1244 B.n545 B.n28 585
R1245 B.n544 B.n543 585
R1246 B.n542 B.n29 585
R1247 B.n541 B.n540 585
R1248 B.n539 B.n30 585
R1249 B.n538 B.n537 585
R1250 B.n536 B.n31 585
R1251 B.n535 B.n534 585
R1252 B.n533 B.n32 585
R1253 B.n532 B.n531 585
R1254 B.n530 B.n33 585
R1255 B.n529 B.n528 585
R1256 B.n527 B.n34 585
R1257 B.n526 B.n525 585
R1258 B.n524 B.n35 585
R1259 B.n523 B.n522 585
R1260 B.n521 B.n36 585
R1261 B.n520 B.n519 585
R1262 B.n518 B.n37 585
R1263 B.n516 B.n515 585
R1264 B.n514 B.n40 585
R1265 B.n513 B.n512 585
R1266 B.n511 B.n41 585
R1267 B.n510 B.n509 585
R1268 B.n508 B.n42 585
R1269 B.n507 B.n506 585
R1270 B.n505 B.n43 585
R1271 B.n504 B.n503 585
R1272 B.n502 B.n44 585
R1273 B.n501 B.n500 585
R1274 B.n499 B.n45 585
R1275 B.n498 B.n497 585
R1276 B.n496 B.n49 585
R1277 B.n495 B.n494 585
R1278 B.n493 B.n50 585
R1279 B.n492 B.n491 585
R1280 B.n490 B.n51 585
R1281 B.n489 B.n488 585
R1282 B.n487 B.n52 585
R1283 B.n486 B.n485 585
R1284 B.n484 B.n53 585
R1285 B.n483 B.n482 585
R1286 B.n481 B.n54 585
R1287 B.n480 B.n479 585
R1288 B.n478 B.n55 585
R1289 B.n477 B.n476 585
R1290 B.n475 B.n56 585
R1291 B.n474 B.n473 585
R1292 B.n472 B.n57 585
R1293 B.n471 B.n470 585
R1294 B.n469 B.n58 585
R1295 B.n468 B.n467 585
R1296 B.n466 B.n59 585
R1297 B.n465 B.n464 585
R1298 B.n463 B.n60 585
R1299 B.n462 B.n461 585
R1300 B.n460 B.n61 585
R1301 B.n459 B.n458 585
R1302 B.n457 B.n62 585
R1303 B.n456 B.n455 585
R1304 B.n454 B.n63 585
R1305 B.n453 B.n452 585
R1306 B.n451 B.n64 585
R1307 B.n450 B.n449 585
R1308 B.n448 B.n65 585
R1309 B.n447 B.n446 585
R1310 B.n445 B.n66 585
R1311 B.n444 B.n443 585
R1312 B.n442 B.n67 585
R1313 B.n441 B.n440 585
R1314 B.n439 B.n68 585
R1315 B.n438 B.n437 585
R1316 B.n436 B.n69 585
R1317 B.n435 B.n434 585
R1318 B.n433 B.n70 585
R1319 B.n432 B.n431 585
R1320 B.n430 B.n71 585
R1321 B.n429 B.n428 585
R1322 B.n427 B.n72 585
R1323 B.n426 B.n425 585
R1324 B.n424 B.n73 585
R1325 B.n596 B.n11 585
R1326 B.n598 B.n597 585
R1327 B.n599 B.n10 585
R1328 B.n601 B.n600 585
R1329 B.n602 B.n9 585
R1330 B.n604 B.n603 585
R1331 B.n605 B.n8 585
R1332 B.n607 B.n606 585
R1333 B.n608 B.n7 585
R1334 B.n610 B.n609 585
R1335 B.n611 B.n6 585
R1336 B.n613 B.n612 585
R1337 B.n614 B.n5 585
R1338 B.n616 B.n615 585
R1339 B.n617 B.n4 585
R1340 B.n619 B.n618 585
R1341 B.n620 B.n3 585
R1342 B.n622 B.n621 585
R1343 B.n623 B.n0 585
R1344 B.n2 B.n1 585
R1345 B.n162 B.n161 585
R1346 B.n164 B.n163 585
R1347 B.n165 B.n160 585
R1348 B.n167 B.n166 585
R1349 B.n168 B.n159 585
R1350 B.n170 B.n169 585
R1351 B.n171 B.n158 585
R1352 B.n173 B.n172 585
R1353 B.n174 B.n157 585
R1354 B.n176 B.n175 585
R1355 B.n177 B.n156 585
R1356 B.n179 B.n178 585
R1357 B.n180 B.n155 585
R1358 B.n182 B.n181 585
R1359 B.n183 B.n154 585
R1360 B.n185 B.n184 585
R1361 B.n186 B.n153 585
R1362 B.n188 B.n187 585
R1363 B.n125 B.t9 582.86
R1364 B.n281 B.t3 582.86
R1365 B.n46 B.t0 582.86
R1366 B.n38 B.t6 582.86
R1367 B.n187 B.n152 545.355
R1368 B.n364 B.n363 545.355
R1369 B.n424 B.n423 545.355
R1370 B.n594 B.n11 545.355
R1371 B.n281 B.t4 466.442
R1372 B.n46 B.t2 466.442
R1373 B.n125 B.t10 466.442
R1374 B.n38 B.t8 466.442
R1375 B.n282 B.t5 440.841
R1376 B.n47 B.t1 440.841
R1377 B.n126 B.t11 440.841
R1378 B.n39 B.t7 440.841
R1379 B.n625 B.n624 256.663
R1380 B.n624 B.n623 235.042
R1381 B.n624 B.n2 235.042
R1382 B.n191 B.n152 163.367
R1383 B.n192 B.n191 163.367
R1384 B.n193 B.n192 163.367
R1385 B.n193 B.n150 163.367
R1386 B.n197 B.n150 163.367
R1387 B.n198 B.n197 163.367
R1388 B.n199 B.n198 163.367
R1389 B.n199 B.n148 163.367
R1390 B.n203 B.n148 163.367
R1391 B.n204 B.n203 163.367
R1392 B.n205 B.n204 163.367
R1393 B.n205 B.n146 163.367
R1394 B.n209 B.n146 163.367
R1395 B.n210 B.n209 163.367
R1396 B.n211 B.n210 163.367
R1397 B.n211 B.n144 163.367
R1398 B.n215 B.n144 163.367
R1399 B.n216 B.n215 163.367
R1400 B.n217 B.n216 163.367
R1401 B.n217 B.n142 163.367
R1402 B.n221 B.n142 163.367
R1403 B.n222 B.n221 163.367
R1404 B.n223 B.n222 163.367
R1405 B.n223 B.n140 163.367
R1406 B.n227 B.n140 163.367
R1407 B.n228 B.n227 163.367
R1408 B.n229 B.n228 163.367
R1409 B.n229 B.n138 163.367
R1410 B.n233 B.n138 163.367
R1411 B.n234 B.n233 163.367
R1412 B.n235 B.n234 163.367
R1413 B.n235 B.n136 163.367
R1414 B.n239 B.n136 163.367
R1415 B.n240 B.n239 163.367
R1416 B.n241 B.n240 163.367
R1417 B.n241 B.n134 163.367
R1418 B.n245 B.n134 163.367
R1419 B.n246 B.n245 163.367
R1420 B.n247 B.n246 163.367
R1421 B.n247 B.n132 163.367
R1422 B.n251 B.n132 163.367
R1423 B.n252 B.n251 163.367
R1424 B.n253 B.n252 163.367
R1425 B.n253 B.n130 163.367
R1426 B.n257 B.n130 163.367
R1427 B.n258 B.n257 163.367
R1428 B.n259 B.n258 163.367
R1429 B.n259 B.n128 163.367
R1430 B.n263 B.n128 163.367
R1431 B.n264 B.n263 163.367
R1432 B.n265 B.n264 163.367
R1433 B.n265 B.n124 163.367
R1434 B.n270 B.n124 163.367
R1435 B.n271 B.n270 163.367
R1436 B.n272 B.n271 163.367
R1437 B.n272 B.n122 163.367
R1438 B.n276 B.n122 163.367
R1439 B.n277 B.n276 163.367
R1440 B.n278 B.n277 163.367
R1441 B.n278 B.n120 163.367
R1442 B.n285 B.n120 163.367
R1443 B.n286 B.n285 163.367
R1444 B.n287 B.n286 163.367
R1445 B.n287 B.n118 163.367
R1446 B.n291 B.n118 163.367
R1447 B.n292 B.n291 163.367
R1448 B.n293 B.n292 163.367
R1449 B.n293 B.n116 163.367
R1450 B.n297 B.n116 163.367
R1451 B.n298 B.n297 163.367
R1452 B.n299 B.n298 163.367
R1453 B.n299 B.n114 163.367
R1454 B.n303 B.n114 163.367
R1455 B.n304 B.n303 163.367
R1456 B.n305 B.n304 163.367
R1457 B.n305 B.n112 163.367
R1458 B.n309 B.n112 163.367
R1459 B.n310 B.n309 163.367
R1460 B.n311 B.n310 163.367
R1461 B.n311 B.n110 163.367
R1462 B.n315 B.n110 163.367
R1463 B.n316 B.n315 163.367
R1464 B.n317 B.n316 163.367
R1465 B.n317 B.n108 163.367
R1466 B.n321 B.n108 163.367
R1467 B.n322 B.n321 163.367
R1468 B.n323 B.n322 163.367
R1469 B.n323 B.n106 163.367
R1470 B.n327 B.n106 163.367
R1471 B.n328 B.n327 163.367
R1472 B.n329 B.n328 163.367
R1473 B.n329 B.n104 163.367
R1474 B.n333 B.n104 163.367
R1475 B.n334 B.n333 163.367
R1476 B.n335 B.n334 163.367
R1477 B.n335 B.n102 163.367
R1478 B.n339 B.n102 163.367
R1479 B.n340 B.n339 163.367
R1480 B.n341 B.n340 163.367
R1481 B.n341 B.n100 163.367
R1482 B.n345 B.n100 163.367
R1483 B.n346 B.n345 163.367
R1484 B.n347 B.n346 163.367
R1485 B.n347 B.n98 163.367
R1486 B.n351 B.n98 163.367
R1487 B.n352 B.n351 163.367
R1488 B.n353 B.n352 163.367
R1489 B.n353 B.n96 163.367
R1490 B.n357 B.n96 163.367
R1491 B.n358 B.n357 163.367
R1492 B.n359 B.n358 163.367
R1493 B.n359 B.n94 163.367
R1494 B.n363 B.n94 163.367
R1495 B.n423 B.n74 163.367
R1496 B.n419 B.n74 163.367
R1497 B.n419 B.n418 163.367
R1498 B.n418 B.n417 163.367
R1499 B.n417 B.n76 163.367
R1500 B.n413 B.n76 163.367
R1501 B.n413 B.n412 163.367
R1502 B.n412 B.n411 163.367
R1503 B.n411 B.n78 163.367
R1504 B.n407 B.n78 163.367
R1505 B.n407 B.n406 163.367
R1506 B.n406 B.n405 163.367
R1507 B.n405 B.n80 163.367
R1508 B.n401 B.n80 163.367
R1509 B.n401 B.n400 163.367
R1510 B.n400 B.n399 163.367
R1511 B.n399 B.n82 163.367
R1512 B.n395 B.n82 163.367
R1513 B.n395 B.n394 163.367
R1514 B.n394 B.n393 163.367
R1515 B.n393 B.n84 163.367
R1516 B.n389 B.n84 163.367
R1517 B.n389 B.n388 163.367
R1518 B.n388 B.n387 163.367
R1519 B.n387 B.n86 163.367
R1520 B.n383 B.n86 163.367
R1521 B.n383 B.n382 163.367
R1522 B.n382 B.n381 163.367
R1523 B.n381 B.n88 163.367
R1524 B.n377 B.n88 163.367
R1525 B.n377 B.n376 163.367
R1526 B.n376 B.n375 163.367
R1527 B.n375 B.n90 163.367
R1528 B.n371 B.n90 163.367
R1529 B.n371 B.n370 163.367
R1530 B.n370 B.n369 163.367
R1531 B.n369 B.n92 163.367
R1532 B.n365 B.n92 163.367
R1533 B.n365 B.n364 163.367
R1534 B.n594 B.n593 163.367
R1535 B.n593 B.n592 163.367
R1536 B.n592 B.n13 163.367
R1537 B.n588 B.n13 163.367
R1538 B.n588 B.n587 163.367
R1539 B.n587 B.n586 163.367
R1540 B.n586 B.n15 163.367
R1541 B.n582 B.n15 163.367
R1542 B.n582 B.n581 163.367
R1543 B.n581 B.n580 163.367
R1544 B.n580 B.n17 163.367
R1545 B.n576 B.n17 163.367
R1546 B.n576 B.n575 163.367
R1547 B.n575 B.n574 163.367
R1548 B.n574 B.n19 163.367
R1549 B.n570 B.n19 163.367
R1550 B.n570 B.n569 163.367
R1551 B.n569 B.n568 163.367
R1552 B.n568 B.n21 163.367
R1553 B.n564 B.n21 163.367
R1554 B.n564 B.n563 163.367
R1555 B.n563 B.n562 163.367
R1556 B.n562 B.n23 163.367
R1557 B.n558 B.n23 163.367
R1558 B.n558 B.n557 163.367
R1559 B.n557 B.n556 163.367
R1560 B.n556 B.n25 163.367
R1561 B.n552 B.n25 163.367
R1562 B.n552 B.n551 163.367
R1563 B.n551 B.n550 163.367
R1564 B.n550 B.n27 163.367
R1565 B.n546 B.n27 163.367
R1566 B.n546 B.n545 163.367
R1567 B.n545 B.n544 163.367
R1568 B.n544 B.n29 163.367
R1569 B.n540 B.n29 163.367
R1570 B.n540 B.n539 163.367
R1571 B.n539 B.n538 163.367
R1572 B.n538 B.n31 163.367
R1573 B.n534 B.n31 163.367
R1574 B.n534 B.n533 163.367
R1575 B.n533 B.n532 163.367
R1576 B.n532 B.n33 163.367
R1577 B.n528 B.n33 163.367
R1578 B.n528 B.n527 163.367
R1579 B.n527 B.n526 163.367
R1580 B.n526 B.n35 163.367
R1581 B.n522 B.n35 163.367
R1582 B.n522 B.n521 163.367
R1583 B.n521 B.n520 163.367
R1584 B.n520 B.n37 163.367
R1585 B.n515 B.n37 163.367
R1586 B.n515 B.n514 163.367
R1587 B.n514 B.n513 163.367
R1588 B.n513 B.n41 163.367
R1589 B.n509 B.n41 163.367
R1590 B.n509 B.n508 163.367
R1591 B.n508 B.n507 163.367
R1592 B.n507 B.n43 163.367
R1593 B.n503 B.n43 163.367
R1594 B.n503 B.n502 163.367
R1595 B.n502 B.n501 163.367
R1596 B.n501 B.n45 163.367
R1597 B.n497 B.n45 163.367
R1598 B.n497 B.n496 163.367
R1599 B.n496 B.n495 163.367
R1600 B.n495 B.n50 163.367
R1601 B.n491 B.n50 163.367
R1602 B.n491 B.n490 163.367
R1603 B.n490 B.n489 163.367
R1604 B.n489 B.n52 163.367
R1605 B.n485 B.n52 163.367
R1606 B.n485 B.n484 163.367
R1607 B.n484 B.n483 163.367
R1608 B.n483 B.n54 163.367
R1609 B.n479 B.n54 163.367
R1610 B.n479 B.n478 163.367
R1611 B.n478 B.n477 163.367
R1612 B.n477 B.n56 163.367
R1613 B.n473 B.n56 163.367
R1614 B.n473 B.n472 163.367
R1615 B.n472 B.n471 163.367
R1616 B.n471 B.n58 163.367
R1617 B.n467 B.n58 163.367
R1618 B.n467 B.n466 163.367
R1619 B.n466 B.n465 163.367
R1620 B.n465 B.n60 163.367
R1621 B.n461 B.n60 163.367
R1622 B.n461 B.n460 163.367
R1623 B.n460 B.n459 163.367
R1624 B.n459 B.n62 163.367
R1625 B.n455 B.n62 163.367
R1626 B.n455 B.n454 163.367
R1627 B.n454 B.n453 163.367
R1628 B.n453 B.n64 163.367
R1629 B.n449 B.n64 163.367
R1630 B.n449 B.n448 163.367
R1631 B.n448 B.n447 163.367
R1632 B.n447 B.n66 163.367
R1633 B.n443 B.n66 163.367
R1634 B.n443 B.n442 163.367
R1635 B.n442 B.n441 163.367
R1636 B.n441 B.n68 163.367
R1637 B.n437 B.n68 163.367
R1638 B.n437 B.n436 163.367
R1639 B.n436 B.n435 163.367
R1640 B.n435 B.n70 163.367
R1641 B.n431 B.n70 163.367
R1642 B.n431 B.n430 163.367
R1643 B.n430 B.n429 163.367
R1644 B.n429 B.n72 163.367
R1645 B.n425 B.n72 163.367
R1646 B.n425 B.n424 163.367
R1647 B.n598 B.n11 163.367
R1648 B.n599 B.n598 163.367
R1649 B.n600 B.n599 163.367
R1650 B.n600 B.n9 163.367
R1651 B.n604 B.n9 163.367
R1652 B.n605 B.n604 163.367
R1653 B.n606 B.n605 163.367
R1654 B.n606 B.n7 163.367
R1655 B.n610 B.n7 163.367
R1656 B.n611 B.n610 163.367
R1657 B.n612 B.n611 163.367
R1658 B.n612 B.n5 163.367
R1659 B.n616 B.n5 163.367
R1660 B.n617 B.n616 163.367
R1661 B.n618 B.n617 163.367
R1662 B.n618 B.n3 163.367
R1663 B.n622 B.n3 163.367
R1664 B.n623 B.n622 163.367
R1665 B.n162 B.n2 163.367
R1666 B.n163 B.n162 163.367
R1667 B.n163 B.n160 163.367
R1668 B.n167 B.n160 163.367
R1669 B.n168 B.n167 163.367
R1670 B.n169 B.n168 163.367
R1671 B.n169 B.n158 163.367
R1672 B.n173 B.n158 163.367
R1673 B.n174 B.n173 163.367
R1674 B.n175 B.n174 163.367
R1675 B.n175 B.n156 163.367
R1676 B.n179 B.n156 163.367
R1677 B.n180 B.n179 163.367
R1678 B.n181 B.n180 163.367
R1679 B.n181 B.n154 163.367
R1680 B.n185 B.n154 163.367
R1681 B.n186 B.n185 163.367
R1682 B.n187 B.n186 163.367
R1683 B.n267 B.n126 59.5399
R1684 B.n283 B.n282 59.5399
R1685 B.n48 B.n47 59.5399
R1686 B.n517 B.n39 59.5399
R1687 B.n596 B.n595 35.4346
R1688 B.n422 B.n73 35.4346
R1689 B.n362 B.n93 35.4346
R1690 B.n189 B.n188 35.4346
R1691 B.n126 B.n125 25.6005
R1692 B.n282 B.n281 25.6005
R1693 B.n47 B.n46 25.6005
R1694 B.n39 B.n38 25.6005
R1695 B B.n625 18.0485
R1696 B.n597 B.n596 10.6151
R1697 B.n597 B.n10 10.6151
R1698 B.n601 B.n10 10.6151
R1699 B.n602 B.n601 10.6151
R1700 B.n603 B.n602 10.6151
R1701 B.n603 B.n8 10.6151
R1702 B.n607 B.n8 10.6151
R1703 B.n608 B.n607 10.6151
R1704 B.n609 B.n608 10.6151
R1705 B.n609 B.n6 10.6151
R1706 B.n613 B.n6 10.6151
R1707 B.n614 B.n613 10.6151
R1708 B.n615 B.n614 10.6151
R1709 B.n615 B.n4 10.6151
R1710 B.n619 B.n4 10.6151
R1711 B.n620 B.n619 10.6151
R1712 B.n621 B.n620 10.6151
R1713 B.n621 B.n0 10.6151
R1714 B.n595 B.n12 10.6151
R1715 B.n591 B.n12 10.6151
R1716 B.n591 B.n590 10.6151
R1717 B.n590 B.n589 10.6151
R1718 B.n589 B.n14 10.6151
R1719 B.n585 B.n14 10.6151
R1720 B.n585 B.n584 10.6151
R1721 B.n584 B.n583 10.6151
R1722 B.n583 B.n16 10.6151
R1723 B.n579 B.n16 10.6151
R1724 B.n579 B.n578 10.6151
R1725 B.n578 B.n577 10.6151
R1726 B.n577 B.n18 10.6151
R1727 B.n573 B.n18 10.6151
R1728 B.n573 B.n572 10.6151
R1729 B.n572 B.n571 10.6151
R1730 B.n571 B.n20 10.6151
R1731 B.n567 B.n20 10.6151
R1732 B.n567 B.n566 10.6151
R1733 B.n566 B.n565 10.6151
R1734 B.n565 B.n22 10.6151
R1735 B.n561 B.n22 10.6151
R1736 B.n561 B.n560 10.6151
R1737 B.n560 B.n559 10.6151
R1738 B.n559 B.n24 10.6151
R1739 B.n555 B.n24 10.6151
R1740 B.n555 B.n554 10.6151
R1741 B.n554 B.n553 10.6151
R1742 B.n553 B.n26 10.6151
R1743 B.n549 B.n26 10.6151
R1744 B.n549 B.n548 10.6151
R1745 B.n548 B.n547 10.6151
R1746 B.n547 B.n28 10.6151
R1747 B.n543 B.n28 10.6151
R1748 B.n543 B.n542 10.6151
R1749 B.n542 B.n541 10.6151
R1750 B.n541 B.n30 10.6151
R1751 B.n537 B.n30 10.6151
R1752 B.n537 B.n536 10.6151
R1753 B.n536 B.n535 10.6151
R1754 B.n535 B.n32 10.6151
R1755 B.n531 B.n32 10.6151
R1756 B.n531 B.n530 10.6151
R1757 B.n530 B.n529 10.6151
R1758 B.n529 B.n34 10.6151
R1759 B.n525 B.n34 10.6151
R1760 B.n525 B.n524 10.6151
R1761 B.n524 B.n523 10.6151
R1762 B.n523 B.n36 10.6151
R1763 B.n519 B.n36 10.6151
R1764 B.n519 B.n518 10.6151
R1765 B.n516 B.n40 10.6151
R1766 B.n512 B.n40 10.6151
R1767 B.n512 B.n511 10.6151
R1768 B.n511 B.n510 10.6151
R1769 B.n510 B.n42 10.6151
R1770 B.n506 B.n42 10.6151
R1771 B.n506 B.n505 10.6151
R1772 B.n505 B.n504 10.6151
R1773 B.n504 B.n44 10.6151
R1774 B.n500 B.n499 10.6151
R1775 B.n499 B.n498 10.6151
R1776 B.n498 B.n49 10.6151
R1777 B.n494 B.n49 10.6151
R1778 B.n494 B.n493 10.6151
R1779 B.n493 B.n492 10.6151
R1780 B.n492 B.n51 10.6151
R1781 B.n488 B.n51 10.6151
R1782 B.n488 B.n487 10.6151
R1783 B.n487 B.n486 10.6151
R1784 B.n486 B.n53 10.6151
R1785 B.n482 B.n53 10.6151
R1786 B.n482 B.n481 10.6151
R1787 B.n481 B.n480 10.6151
R1788 B.n480 B.n55 10.6151
R1789 B.n476 B.n55 10.6151
R1790 B.n476 B.n475 10.6151
R1791 B.n475 B.n474 10.6151
R1792 B.n474 B.n57 10.6151
R1793 B.n470 B.n57 10.6151
R1794 B.n470 B.n469 10.6151
R1795 B.n469 B.n468 10.6151
R1796 B.n468 B.n59 10.6151
R1797 B.n464 B.n59 10.6151
R1798 B.n464 B.n463 10.6151
R1799 B.n463 B.n462 10.6151
R1800 B.n462 B.n61 10.6151
R1801 B.n458 B.n61 10.6151
R1802 B.n458 B.n457 10.6151
R1803 B.n457 B.n456 10.6151
R1804 B.n456 B.n63 10.6151
R1805 B.n452 B.n63 10.6151
R1806 B.n452 B.n451 10.6151
R1807 B.n451 B.n450 10.6151
R1808 B.n450 B.n65 10.6151
R1809 B.n446 B.n65 10.6151
R1810 B.n446 B.n445 10.6151
R1811 B.n445 B.n444 10.6151
R1812 B.n444 B.n67 10.6151
R1813 B.n440 B.n67 10.6151
R1814 B.n440 B.n439 10.6151
R1815 B.n439 B.n438 10.6151
R1816 B.n438 B.n69 10.6151
R1817 B.n434 B.n69 10.6151
R1818 B.n434 B.n433 10.6151
R1819 B.n433 B.n432 10.6151
R1820 B.n432 B.n71 10.6151
R1821 B.n428 B.n71 10.6151
R1822 B.n428 B.n427 10.6151
R1823 B.n427 B.n426 10.6151
R1824 B.n426 B.n73 10.6151
R1825 B.n422 B.n421 10.6151
R1826 B.n421 B.n420 10.6151
R1827 B.n420 B.n75 10.6151
R1828 B.n416 B.n75 10.6151
R1829 B.n416 B.n415 10.6151
R1830 B.n415 B.n414 10.6151
R1831 B.n414 B.n77 10.6151
R1832 B.n410 B.n77 10.6151
R1833 B.n410 B.n409 10.6151
R1834 B.n409 B.n408 10.6151
R1835 B.n408 B.n79 10.6151
R1836 B.n404 B.n79 10.6151
R1837 B.n404 B.n403 10.6151
R1838 B.n403 B.n402 10.6151
R1839 B.n402 B.n81 10.6151
R1840 B.n398 B.n81 10.6151
R1841 B.n398 B.n397 10.6151
R1842 B.n397 B.n396 10.6151
R1843 B.n396 B.n83 10.6151
R1844 B.n392 B.n83 10.6151
R1845 B.n392 B.n391 10.6151
R1846 B.n391 B.n390 10.6151
R1847 B.n390 B.n85 10.6151
R1848 B.n386 B.n85 10.6151
R1849 B.n386 B.n385 10.6151
R1850 B.n385 B.n384 10.6151
R1851 B.n384 B.n87 10.6151
R1852 B.n380 B.n87 10.6151
R1853 B.n380 B.n379 10.6151
R1854 B.n379 B.n378 10.6151
R1855 B.n378 B.n89 10.6151
R1856 B.n374 B.n89 10.6151
R1857 B.n374 B.n373 10.6151
R1858 B.n373 B.n372 10.6151
R1859 B.n372 B.n91 10.6151
R1860 B.n368 B.n91 10.6151
R1861 B.n368 B.n367 10.6151
R1862 B.n367 B.n366 10.6151
R1863 B.n366 B.n93 10.6151
R1864 B.n161 B.n1 10.6151
R1865 B.n164 B.n161 10.6151
R1866 B.n165 B.n164 10.6151
R1867 B.n166 B.n165 10.6151
R1868 B.n166 B.n159 10.6151
R1869 B.n170 B.n159 10.6151
R1870 B.n171 B.n170 10.6151
R1871 B.n172 B.n171 10.6151
R1872 B.n172 B.n157 10.6151
R1873 B.n176 B.n157 10.6151
R1874 B.n177 B.n176 10.6151
R1875 B.n178 B.n177 10.6151
R1876 B.n178 B.n155 10.6151
R1877 B.n182 B.n155 10.6151
R1878 B.n183 B.n182 10.6151
R1879 B.n184 B.n183 10.6151
R1880 B.n184 B.n153 10.6151
R1881 B.n188 B.n153 10.6151
R1882 B.n190 B.n189 10.6151
R1883 B.n190 B.n151 10.6151
R1884 B.n194 B.n151 10.6151
R1885 B.n195 B.n194 10.6151
R1886 B.n196 B.n195 10.6151
R1887 B.n196 B.n149 10.6151
R1888 B.n200 B.n149 10.6151
R1889 B.n201 B.n200 10.6151
R1890 B.n202 B.n201 10.6151
R1891 B.n202 B.n147 10.6151
R1892 B.n206 B.n147 10.6151
R1893 B.n207 B.n206 10.6151
R1894 B.n208 B.n207 10.6151
R1895 B.n208 B.n145 10.6151
R1896 B.n212 B.n145 10.6151
R1897 B.n213 B.n212 10.6151
R1898 B.n214 B.n213 10.6151
R1899 B.n214 B.n143 10.6151
R1900 B.n218 B.n143 10.6151
R1901 B.n219 B.n218 10.6151
R1902 B.n220 B.n219 10.6151
R1903 B.n220 B.n141 10.6151
R1904 B.n224 B.n141 10.6151
R1905 B.n225 B.n224 10.6151
R1906 B.n226 B.n225 10.6151
R1907 B.n226 B.n139 10.6151
R1908 B.n230 B.n139 10.6151
R1909 B.n231 B.n230 10.6151
R1910 B.n232 B.n231 10.6151
R1911 B.n232 B.n137 10.6151
R1912 B.n236 B.n137 10.6151
R1913 B.n237 B.n236 10.6151
R1914 B.n238 B.n237 10.6151
R1915 B.n238 B.n135 10.6151
R1916 B.n242 B.n135 10.6151
R1917 B.n243 B.n242 10.6151
R1918 B.n244 B.n243 10.6151
R1919 B.n244 B.n133 10.6151
R1920 B.n248 B.n133 10.6151
R1921 B.n249 B.n248 10.6151
R1922 B.n250 B.n249 10.6151
R1923 B.n250 B.n131 10.6151
R1924 B.n254 B.n131 10.6151
R1925 B.n255 B.n254 10.6151
R1926 B.n256 B.n255 10.6151
R1927 B.n256 B.n129 10.6151
R1928 B.n260 B.n129 10.6151
R1929 B.n261 B.n260 10.6151
R1930 B.n262 B.n261 10.6151
R1931 B.n262 B.n127 10.6151
R1932 B.n266 B.n127 10.6151
R1933 B.n269 B.n268 10.6151
R1934 B.n269 B.n123 10.6151
R1935 B.n273 B.n123 10.6151
R1936 B.n274 B.n273 10.6151
R1937 B.n275 B.n274 10.6151
R1938 B.n275 B.n121 10.6151
R1939 B.n279 B.n121 10.6151
R1940 B.n280 B.n279 10.6151
R1941 B.n284 B.n280 10.6151
R1942 B.n288 B.n119 10.6151
R1943 B.n289 B.n288 10.6151
R1944 B.n290 B.n289 10.6151
R1945 B.n290 B.n117 10.6151
R1946 B.n294 B.n117 10.6151
R1947 B.n295 B.n294 10.6151
R1948 B.n296 B.n295 10.6151
R1949 B.n296 B.n115 10.6151
R1950 B.n300 B.n115 10.6151
R1951 B.n301 B.n300 10.6151
R1952 B.n302 B.n301 10.6151
R1953 B.n302 B.n113 10.6151
R1954 B.n306 B.n113 10.6151
R1955 B.n307 B.n306 10.6151
R1956 B.n308 B.n307 10.6151
R1957 B.n308 B.n111 10.6151
R1958 B.n312 B.n111 10.6151
R1959 B.n313 B.n312 10.6151
R1960 B.n314 B.n313 10.6151
R1961 B.n314 B.n109 10.6151
R1962 B.n318 B.n109 10.6151
R1963 B.n319 B.n318 10.6151
R1964 B.n320 B.n319 10.6151
R1965 B.n320 B.n107 10.6151
R1966 B.n324 B.n107 10.6151
R1967 B.n325 B.n324 10.6151
R1968 B.n326 B.n325 10.6151
R1969 B.n326 B.n105 10.6151
R1970 B.n330 B.n105 10.6151
R1971 B.n331 B.n330 10.6151
R1972 B.n332 B.n331 10.6151
R1973 B.n332 B.n103 10.6151
R1974 B.n336 B.n103 10.6151
R1975 B.n337 B.n336 10.6151
R1976 B.n338 B.n337 10.6151
R1977 B.n338 B.n101 10.6151
R1978 B.n342 B.n101 10.6151
R1979 B.n343 B.n342 10.6151
R1980 B.n344 B.n343 10.6151
R1981 B.n344 B.n99 10.6151
R1982 B.n348 B.n99 10.6151
R1983 B.n349 B.n348 10.6151
R1984 B.n350 B.n349 10.6151
R1985 B.n350 B.n97 10.6151
R1986 B.n354 B.n97 10.6151
R1987 B.n355 B.n354 10.6151
R1988 B.n356 B.n355 10.6151
R1989 B.n356 B.n95 10.6151
R1990 B.n360 B.n95 10.6151
R1991 B.n361 B.n360 10.6151
R1992 B.n362 B.n361 10.6151
R1993 B.n518 B.n517 9.36635
R1994 B.n500 B.n48 9.36635
R1995 B.n267 B.n266 9.36635
R1996 B.n283 B.n119 9.36635
R1997 B.n625 B.n0 8.11757
R1998 B.n625 B.n1 8.11757
R1999 B.n517 B.n516 1.24928
R2000 B.n48 B.n44 1.24928
R2001 B.n268 B.n267 1.24928
R2002 B.n284 B.n283 1.24928
R2003 VN.n0 VN.t1 438.531
R2004 VN.n1 VN.t2 438.531
R2005 VN.n1 VN.t0 438.445
R2006 VN.n0 VN.t3 438.445
R2007 VN VN.n1 75.6448
R2008 VN VN.n0 31.2622
R2009 VDD2.n2 VDD2.n0 108.992
R2010 VDD2.n2 VDD2.n1 68.4058
R2011 VDD2.n1 VDD2.t3 2.08282
R2012 VDD2.n1 VDD2.t1 2.08282
R2013 VDD2.n0 VDD2.t2 2.08282
R2014 VDD2.n0 VDD2.t0 2.08282
R2015 VDD2 VDD2.n2 0.0586897
C0 VTAIL B 5.05672f
C1 VDD1 VTAIL 7.40388f
C2 VTAIL VP 4.1882f
C3 w_n1762_n4090# B 8.27662f
C4 VTAIL VDD2 7.44729f
C5 VDD1 w_n1762_n4090# 1.2272f
C6 VP w_n1762_n4090# 2.97746f
C7 VDD1 B 1.07485f
C8 VDD2 w_n1762_n4090# 1.24773f
C9 VP B 1.20648f
C10 VDD1 VP 4.79733f
C11 VDD2 B 1.1008f
C12 VDD1 VDD2 0.636212f
C13 VP VDD2 0.291969f
C14 VTAIL VN 4.17409f
C15 w_n1762_n4090# VN 2.75501f
C16 VN B 0.844846f
C17 VDD1 VN 0.147656f
C18 VP VN 5.70034f
C19 VTAIL w_n1762_n4090# 4.96623f
C20 VDD2 VN 4.65335f
C21 VDD2 VSUBS 0.800765f
C22 VDD1 VSUBS 5.511486f
C23 VTAIL VSUBS 1.099068f
C24 VN VSUBS 5.78619f
C25 VP VSUBS 1.598879f
C26 B VSUBS 3.184022f
C27 w_n1762_n4090# VSUBS 88.3185f
C28 VDD2.t2 VSUBS 0.336252f
C29 VDD2.t0 VSUBS 0.336252f
C30 VDD2.n0 VSUBS 3.52541f
C31 VDD2.t3 VSUBS 0.336252f
C32 VDD2.t1 VSUBS 0.336252f
C33 VDD2.n1 VSUBS 2.72153f
C34 VDD2.n2 VSUBS 4.40223f
C35 VN.t1 VSUBS 2.27826f
C36 VN.t3 VSUBS 2.27807f
C37 VN.n0 VSUBS 1.64583f
C38 VN.t2 VSUBS 2.27826f
C39 VN.t0 VSUBS 2.27807f
C40 VN.n1 VSUBS 3.09925f
C41 B.n0 VSUBS 0.006694f
C42 B.n1 VSUBS 0.006694f
C43 B.n2 VSUBS 0.0099f
C44 B.n3 VSUBS 0.007587f
C45 B.n4 VSUBS 0.007587f
C46 B.n5 VSUBS 0.007587f
C47 B.n6 VSUBS 0.007587f
C48 B.n7 VSUBS 0.007587f
C49 B.n8 VSUBS 0.007587f
C50 B.n9 VSUBS 0.007587f
C51 B.n10 VSUBS 0.007587f
C52 B.n11 VSUBS 0.01819f
C53 B.n12 VSUBS 0.007587f
C54 B.n13 VSUBS 0.007587f
C55 B.n14 VSUBS 0.007587f
C56 B.n15 VSUBS 0.007587f
C57 B.n16 VSUBS 0.007587f
C58 B.n17 VSUBS 0.007587f
C59 B.n18 VSUBS 0.007587f
C60 B.n19 VSUBS 0.007587f
C61 B.n20 VSUBS 0.007587f
C62 B.n21 VSUBS 0.007587f
C63 B.n22 VSUBS 0.007587f
C64 B.n23 VSUBS 0.007587f
C65 B.n24 VSUBS 0.007587f
C66 B.n25 VSUBS 0.007587f
C67 B.n26 VSUBS 0.007587f
C68 B.n27 VSUBS 0.007587f
C69 B.n28 VSUBS 0.007587f
C70 B.n29 VSUBS 0.007587f
C71 B.n30 VSUBS 0.007587f
C72 B.n31 VSUBS 0.007587f
C73 B.n32 VSUBS 0.007587f
C74 B.n33 VSUBS 0.007587f
C75 B.n34 VSUBS 0.007587f
C76 B.n35 VSUBS 0.007587f
C77 B.n36 VSUBS 0.007587f
C78 B.n37 VSUBS 0.007587f
C79 B.t7 VSUBS 0.318825f
C80 B.t8 VSUBS 0.335633f
C81 B.t6 VSUBS 0.696695f
C82 B.n38 VSUBS 0.451597f
C83 B.n39 VSUBS 0.317067f
C84 B.n40 VSUBS 0.007587f
C85 B.n41 VSUBS 0.007587f
C86 B.n42 VSUBS 0.007587f
C87 B.n43 VSUBS 0.007587f
C88 B.n44 VSUBS 0.00424f
C89 B.n45 VSUBS 0.007587f
C90 B.t1 VSUBS 0.318829f
C91 B.t2 VSUBS 0.335636f
C92 B.t0 VSUBS 0.696695f
C93 B.n46 VSUBS 0.451594f
C94 B.n47 VSUBS 0.317063f
C95 B.n48 VSUBS 0.017578f
C96 B.n49 VSUBS 0.007587f
C97 B.n50 VSUBS 0.007587f
C98 B.n51 VSUBS 0.007587f
C99 B.n52 VSUBS 0.007587f
C100 B.n53 VSUBS 0.007587f
C101 B.n54 VSUBS 0.007587f
C102 B.n55 VSUBS 0.007587f
C103 B.n56 VSUBS 0.007587f
C104 B.n57 VSUBS 0.007587f
C105 B.n58 VSUBS 0.007587f
C106 B.n59 VSUBS 0.007587f
C107 B.n60 VSUBS 0.007587f
C108 B.n61 VSUBS 0.007587f
C109 B.n62 VSUBS 0.007587f
C110 B.n63 VSUBS 0.007587f
C111 B.n64 VSUBS 0.007587f
C112 B.n65 VSUBS 0.007587f
C113 B.n66 VSUBS 0.007587f
C114 B.n67 VSUBS 0.007587f
C115 B.n68 VSUBS 0.007587f
C116 B.n69 VSUBS 0.007587f
C117 B.n70 VSUBS 0.007587f
C118 B.n71 VSUBS 0.007587f
C119 B.n72 VSUBS 0.007587f
C120 B.n73 VSUBS 0.019298f
C121 B.n74 VSUBS 0.007587f
C122 B.n75 VSUBS 0.007587f
C123 B.n76 VSUBS 0.007587f
C124 B.n77 VSUBS 0.007587f
C125 B.n78 VSUBS 0.007587f
C126 B.n79 VSUBS 0.007587f
C127 B.n80 VSUBS 0.007587f
C128 B.n81 VSUBS 0.007587f
C129 B.n82 VSUBS 0.007587f
C130 B.n83 VSUBS 0.007587f
C131 B.n84 VSUBS 0.007587f
C132 B.n85 VSUBS 0.007587f
C133 B.n86 VSUBS 0.007587f
C134 B.n87 VSUBS 0.007587f
C135 B.n88 VSUBS 0.007587f
C136 B.n89 VSUBS 0.007587f
C137 B.n90 VSUBS 0.007587f
C138 B.n91 VSUBS 0.007587f
C139 B.n92 VSUBS 0.007587f
C140 B.n93 VSUBS 0.019016f
C141 B.n94 VSUBS 0.007587f
C142 B.n95 VSUBS 0.007587f
C143 B.n96 VSUBS 0.007587f
C144 B.n97 VSUBS 0.007587f
C145 B.n98 VSUBS 0.007587f
C146 B.n99 VSUBS 0.007587f
C147 B.n100 VSUBS 0.007587f
C148 B.n101 VSUBS 0.007587f
C149 B.n102 VSUBS 0.007587f
C150 B.n103 VSUBS 0.007587f
C151 B.n104 VSUBS 0.007587f
C152 B.n105 VSUBS 0.007587f
C153 B.n106 VSUBS 0.007587f
C154 B.n107 VSUBS 0.007587f
C155 B.n108 VSUBS 0.007587f
C156 B.n109 VSUBS 0.007587f
C157 B.n110 VSUBS 0.007587f
C158 B.n111 VSUBS 0.007587f
C159 B.n112 VSUBS 0.007587f
C160 B.n113 VSUBS 0.007587f
C161 B.n114 VSUBS 0.007587f
C162 B.n115 VSUBS 0.007587f
C163 B.n116 VSUBS 0.007587f
C164 B.n117 VSUBS 0.007587f
C165 B.n118 VSUBS 0.007587f
C166 B.n119 VSUBS 0.007141f
C167 B.n120 VSUBS 0.007587f
C168 B.n121 VSUBS 0.007587f
C169 B.n122 VSUBS 0.007587f
C170 B.n123 VSUBS 0.007587f
C171 B.n124 VSUBS 0.007587f
C172 B.t11 VSUBS 0.318825f
C173 B.t10 VSUBS 0.335633f
C174 B.t9 VSUBS 0.696695f
C175 B.n125 VSUBS 0.451597f
C176 B.n126 VSUBS 0.317067f
C177 B.n127 VSUBS 0.007587f
C178 B.n128 VSUBS 0.007587f
C179 B.n129 VSUBS 0.007587f
C180 B.n130 VSUBS 0.007587f
C181 B.n131 VSUBS 0.007587f
C182 B.n132 VSUBS 0.007587f
C183 B.n133 VSUBS 0.007587f
C184 B.n134 VSUBS 0.007587f
C185 B.n135 VSUBS 0.007587f
C186 B.n136 VSUBS 0.007587f
C187 B.n137 VSUBS 0.007587f
C188 B.n138 VSUBS 0.007587f
C189 B.n139 VSUBS 0.007587f
C190 B.n140 VSUBS 0.007587f
C191 B.n141 VSUBS 0.007587f
C192 B.n142 VSUBS 0.007587f
C193 B.n143 VSUBS 0.007587f
C194 B.n144 VSUBS 0.007587f
C195 B.n145 VSUBS 0.007587f
C196 B.n146 VSUBS 0.007587f
C197 B.n147 VSUBS 0.007587f
C198 B.n148 VSUBS 0.007587f
C199 B.n149 VSUBS 0.007587f
C200 B.n150 VSUBS 0.007587f
C201 B.n151 VSUBS 0.007587f
C202 B.n152 VSUBS 0.019298f
C203 B.n153 VSUBS 0.007587f
C204 B.n154 VSUBS 0.007587f
C205 B.n155 VSUBS 0.007587f
C206 B.n156 VSUBS 0.007587f
C207 B.n157 VSUBS 0.007587f
C208 B.n158 VSUBS 0.007587f
C209 B.n159 VSUBS 0.007587f
C210 B.n160 VSUBS 0.007587f
C211 B.n161 VSUBS 0.007587f
C212 B.n162 VSUBS 0.007587f
C213 B.n163 VSUBS 0.007587f
C214 B.n164 VSUBS 0.007587f
C215 B.n165 VSUBS 0.007587f
C216 B.n166 VSUBS 0.007587f
C217 B.n167 VSUBS 0.007587f
C218 B.n168 VSUBS 0.007587f
C219 B.n169 VSUBS 0.007587f
C220 B.n170 VSUBS 0.007587f
C221 B.n171 VSUBS 0.007587f
C222 B.n172 VSUBS 0.007587f
C223 B.n173 VSUBS 0.007587f
C224 B.n174 VSUBS 0.007587f
C225 B.n175 VSUBS 0.007587f
C226 B.n176 VSUBS 0.007587f
C227 B.n177 VSUBS 0.007587f
C228 B.n178 VSUBS 0.007587f
C229 B.n179 VSUBS 0.007587f
C230 B.n180 VSUBS 0.007587f
C231 B.n181 VSUBS 0.007587f
C232 B.n182 VSUBS 0.007587f
C233 B.n183 VSUBS 0.007587f
C234 B.n184 VSUBS 0.007587f
C235 B.n185 VSUBS 0.007587f
C236 B.n186 VSUBS 0.007587f
C237 B.n187 VSUBS 0.01819f
C238 B.n188 VSUBS 0.01819f
C239 B.n189 VSUBS 0.019298f
C240 B.n190 VSUBS 0.007587f
C241 B.n191 VSUBS 0.007587f
C242 B.n192 VSUBS 0.007587f
C243 B.n193 VSUBS 0.007587f
C244 B.n194 VSUBS 0.007587f
C245 B.n195 VSUBS 0.007587f
C246 B.n196 VSUBS 0.007587f
C247 B.n197 VSUBS 0.007587f
C248 B.n198 VSUBS 0.007587f
C249 B.n199 VSUBS 0.007587f
C250 B.n200 VSUBS 0.007587f
C251 B.n201 VSUBS 0.007587f
C252 B.n202 VSUBS 0.007587f
C253 B.n203 VSUBS 0.007587f
C254 B.n204 VSUBS 0.007587f
C255 B.n205 VSUBS 0.007587f
C256 B.n206 VSUBS 0.007587f
C257 B.n207 VSUBS 0.007587f
C258 B.n208 VSUBS 0.007587f
C259 B.n209 VSUBS 0.007587f
C260 B.n210 VSUBS 0.007587f
C261 B.n211 VSUBS 0.007587f
C262 B.n212 VSUBS 0.007587f
C263 B.n213 VSUBS 0.007587f
C264 B.n214 VSUBS 0.007587f
C265 B.n215 VSUBS 0.007587f
C266 B.n216 VSUBS 0.007587f
C267 B.n217 VSUBS 0.007587f
C268 B.n218 VSUBS 0.007587f
C269 B.n219 VSUBS 0.007587f
C270 B.n220 VSUBS 0.007587f
C271 B.n221 VSUBS 0.007587f
C272 B.n222 VSUBS 0.007587f
C273 B.n223 VSUBS 0.007587f
C274 B.n224 VSUBS 0.007587f
C275 B.n225 VSUBS 0.007587f
C276 B.n226 VSUBS 0.007587f
C277 B.n227 VSUBS 0.007587f
C278 B.n228 VSUBS 0.007587f
C279 B.n229 VSUBS 0.007587f
C280 B.n230 VSUBS 0.007587f
C281 B.n231 VSUBS 0.007587f
C282 B.n232 VSUBS 0.007587f
C283 B.n233 VSUBS 0.007587f
C284 B.n234 VSUBS 0.007587f
C285 B.n235 VSUBS 0.007587f
C286 B.n236 VSUBS 0.007587f
C287 B.n237 VSUBS 0.007587f
C288 B.n238 VSUBS 0.007587f
C289 B.n239 VSUBS 0.007587f
C290 B.n240 VSUBS 0.007587f
C291 B.n241 VSUBS 0.007587f
C292 B.n242 VSUBS 0.007587f
C293 B.n243 VSUBS 0.007587f
C294 B.n244 VSUBS 0.007587f
C295 B.n245 VSUBS 0.007587f
C296 B.n246 VSUBS 0.007587f
C297 B.n247 VSUBS 0.007587f
C298 B.n248 VSUBS 0.007587f
C299 B.n249 VSUBS 0.007587f
C300 B.n250 VSUBS 0.007587f
C301 B.n251 VSUBS 0.007587f
C302 B.n252 VSUBS 0.007587f
C303 B.n253 VSUBS 0.007587f
C304 B.n254 VSUBS 0.007587f
C305 B.n255 VSUBS 0.007587f
C306 B.n256 VSUBS 0.007587f
C307 B.n257 VSUBS 0.007587f
C308 B.n258 VSUBS 0.007587f
C309 B.n259 VSUBS 0.007587f
C310 B.n260 VSUBS 0.007587f
C311 B.n261 VSUBS 0.007587f
C312 B.n262 VSUBS 0.007587f
C313 B.n263 VSUBS 0.007587f
C314 B.n264 VSUBS 0.007587f
C315 B.n265 VSUBS 0.007587f
C316 B.n266 VSUBS 0.007141f
C317 B.n267 VSUBS 0.017578f
C318 B.n268 VSUBS 0.00424f
C319 B.n269 VSUBS 0.007587f
C320 B.n270 VSUBS 0.007587f
C321 B.n271 VSUBS 0.007587f
C322 B.n272 VSUBS 0.007587f
C323 B.n273 VSUBS 0.007587f
C324 B.n274 VSUBS 0.007587f
C325 B.n275 VSUBS 0.007587f
C326 B.n276 VSUBS 0.007587f
C327 B.n277 VSUBS 0.007587f
C328 B.n278 VSUBS 0.007587f
C329 B.n279 VSUBS 0.007587f
C330 B.n280 VSUBS 0.007587f
C331 B.t5 VSUBS 0.318829f
C332 B.t4 VSUBS 0.335636f
C333 B.t3 VSUBS 0.696695f
C334 B.n281 VSUBS 0.451594f
C335 B.n282 VSUBS 0.317063f
C336 B.n283 VSUBS 0.017578f
C337 B.n284 VSUBS 0.00424f
C338 B.n285 VSUBS 0.007587f
C339 B.n286 VSUBS 0.007587f
C340 B.n287 VSUBS 0.007587f
C341 B.n288 VSUBS 0.007587f
C342 B.n289 VSUBS 0.007587f
C343 B.n290 VSUBS 0.007587f
C344 B.n291 VSUBS 0.007587f
C345 B.n292 VSUBS 0.007587f
C346 B.n293 VSUBS 0.007587f
C347 B.n294 VSUBS 0.007587f
C348 B.n295 VSUBS 0.007587f
C349 B.n296 VSUBS 0.007587f
C350 B.n297 VSUBS 0.007587f
C351 B.n298 VSUBS 0.007587f
C352 B.n299 VSUBS 0.007587f
C353 B.n300 VSUBS 0.007587f
C354 B.n301 VSUBS 0.007587f
C355 B.n302 VSUBS 0.007587f
C356 B.n303 VSUBS 0.007587f
C357 B.n304 VSUBS 0.007587f
C358 B.n305 VSUBS 0.007587f
C359 B.n306 VSUBS 0.007587f
C360 B.n307 VSUBS 0.007587f
C361 B.n308 VSUBS 0.007587f
C362 B.n309 VSUBS 0.007587f
C363 B.n310 VSUBS 0.007587f
C364 B.n311 VSUBS 0.007587f
C365 B.n312 VSUBS 0.007587f
C366 B.n313 VSUBS 0.007587f
C367 B.n314 VSUBS 0.007587f
C368 B.n315 VSUBS 0.007587f
C369 B.n316 VSUBS 0.007587f
C370 B.n317 VSUBS 0.007587f
C371 B.n318 VSUBS 0.007587f
C372 B.n319 VSUBS 0.007587f
C373 B.n320 VSUBS 0.007587f
C374 B.n321 VSUBS 0.007587f
C375 B.n322 VSUBS 0.007587f
C376 B.n323 VSUBS 0.007587f
C377 B.n324 VSUBS 0.007587f
C378 B.n325 VSUBS 0.007587f
C379 B.n326 VSUBS 0.007587f
C380 B.n327 VSUBS 0.007587f
C381 B.n328 VSUBS 0.007587f
C382 B.n329 VSUBS 0.007587f
C383 B.n330 VSUBS 0.007587f
C384 B.n331 VSUBS 0.007587f
C385 B.n332 VSUBS 0.007587f
C386 B.n333 VSUBS 0.007587f
C387 B.n334 VSUBS 0.007587f
C388 B.n335 VSUBS 0.007587f
C389 B.n336 VSUBS 0.007587f
C390 B.n337 VSUBS 0.007587f
C391 B.n338 VSUBS 0.007587f
C392 B.n339 VSUBS 0.007587f
C393 B.n340 VSUBS 0.007587f
C394 B.n341 VSUBS 0.007587f
C395 B.n342 VSUBS 0.007587f
C396 B.n343 VSUBS 0.007587f
C397 B.n344 VSUBS 0.007587f
C398 B.n345 VSUBS 0.007587f
C399 B.n346 VSUBS 0.007587f
C400 B.n347 VSUBS 0.007587f
C401 B.n348 VSUBS 0.007587f
C402 B.n349 VSUBS 0.007587f
C403 B.n350 VSUBS 0.007587f
C404 B.n351 VSUBS 0.007587f
C405 B.n352 VSUBS 0.007587f
C406 B.n353 VSUBS 0.007587f
C407 B.n354 VSUBS 0.007587f
C408 B.n355 VSUBS 0.007587f
C409 B.n356 VSUBS 0.007587f
C410 B.n357 VSUBS 0.007587f
C411 B.n358 VSUBS 0.007587f
C412 B.n359 VSUBS 0.007587f
C413 B.n360 VSUBS 0.007587f
C414 B.n361 VSUBS 0.007587f
C415 B.n362 VSUBS 0.018472f
C416 B.n363 VSUBS 0.019298f
C417 B.n364 VSUBS 0.01819f
C418 B.n365 VSUBS 0.007587f
C419 B.n366 VSUBS 0.007587f
C420 B.n367 VSUBS 0.007587f
C421 B.n368 VSUBS 0.007587f
C422 B.n369 VSUBS 0.007587f
C423 B.n370 VSUBS 0.007587f
C424 B.n371 VSUBS 0.007587f
C425 B.n372 VSUBS 0.007587f
C426 B.n373 VSUBS 0.007587f
C427 B.n374 VSUBS 0.007587f
C428 B.n375 VSUBS 0.007587f
C429 B.n376 VSUBS 0.007587f
C430 B.n377 VSUBS 0.007587f
C431 B.n378 VSUBS 0.007587f
C432 B.n379 VSUBS 0.007587f
C433 B.n380 VSUBS 0.007587f
C434 B.n381 VSUBS 0.007587f
C435 B.n382 VSUBS 0.007587f
C436 B.n383 VSUBS 0.007587f
C437 B.n384 VSUBS 0.007587f
C438 B.n385 VSUBS 0.007587f
C439 B.n386 VSUBS 0.007587f
C440 B.n387 VSUBS 0.007587f
C441 B.n388 VSUBS 0.007587f
C442 B.n389 VSUBS 0.007587f
C443 B.n390 VSUBS 0.007587f
C444 B.n391 VSUBS 0.007587f
C445 B.n392 VSUBS 0.007587f
C446 B.n393 VSUBS 0.007587f
C447 B.n394 VSUBS 0.007587f
C448 B.n395 VSUBS 0.007587f
C449 B.n396 VSUBS 0.007587f
C450 B.n397 VSUBS 0.007587f
C451 B.n398 VSUBS 0.007587f
C452 B.n399 VSUBS 0.007587f
C453 B.n400 VSUBS 0.007587f
C454 B.n401 VSUBS 0.007587f
C455 B.n402 VSUBS 0.007587f
C456 B.n403 VSUBS 0.007587f
C457 B.n404 VSUBS 0.007587f
C458 B.n405 VSUBS 0.007587f
C459 B.n406 VSUBS 0.007587f
C460 B.n407 VSUBS 0.007587f
C461 B.n408 VSUBS 0.007587f
C462 B.n409 VSUBS 0.007587f
C463 B.n410 VSUBS 0.007587f
C464 B.n411 VSUBS 0.007587f
C465 B.n412 VSUBS 0.007587f
C466 B.n413 VSUBS 0.007587f
C467 B.n414 VSUBS 0.007587f
C468 B.n415 VSUBS 0.007587f
C469 B.n416 VSUBS 0.007587f
C470 B.n417 VSUBS 0.007587f
C471 B.n418 VSUBS 0.007587f
C472 B.n419 VSUBS 0.007587f
C473 B.n420 VSUBS 0.007587f
C474 B.n421 VSUBS 0.007587f
C475 B.n422 VSUBS 0.01819f
C476 B.n423 VSUBS 0.01819f
C477 B.n424 VSUBS 0.019298f
C478 B.n425 VSUBS 0.007587f
C479 B.n426 VSUBS 0.007587f
C480 B.n427 VSUBS 0.007587f
C481 B.n428 VSUBS 0.007587f
C482 B.n429 VSUBS 0.007587f
C483 B.n430 VSUBS 0.007587f
C484 B.n431 VSUBS 0.007587f
C485 B.n432 VSUBS 0.007587f
C486 B.n433 VSUBS 0.007587f
C487 B.n434 VSUBS 0.007587f
C488 B.n435 VSUBS 0.007587f
C489 B.n436 VSUBS 0.007587f
C490 B.n437 VSUBS 0.007587f
C491 B.n438 VSUBS 0.007587f
C492 B.n439 VSUBS 0.007587f
C493 B.n440 VSUBS 0.007587f
C494 B.n441 VSUBS 0.007587f
C495 B.n442 VSUBS 0.007587f
C496 B.n443 VSUBS 0.007587f
C497 B.n444 VSUBS 0.007587f
C498 B.n445 VSUBS 0.007587f
C499 B.n446 VSUBS 0.007587f
C500 B.n447 VSUBS 0.007587f
C501 B.n448 VSUBS 0.007587f
C502 B.n449 VSUBS 0.007587f
C503 B.n450 VSUBS 0.007587f
C504 B.n451 VSUBS 0.007587f
C505 B.n452 VSUBS 0.007587f
C506 B.n453 VSUBS 0.007587f
C507 B.n454 VSUBS 0.007587f
C508 B.n455 VSUBS 0.007587f
C509 B.n456 VSUBS 0.007587f
C510 B.n457 VSUBS 0.007587f
C511 B.n458 VSUBS 0.007587f
C512 B.n459 VSUBS 0.007587f
C513 B.n460 VSUBS 0.007587f
C514 B.n461 VSUBS 0.007587f
C515 B.n462 VSUBS 0.007587f
C516 B.n463 VSUBS 0.007587f
C517 B.n464 VSUBS 0.007587f
C518 B.n465 VSUBS 0.007587f
C519 B.n466 VSUBS 0.007587f
C520 B.n467 VSUBS 0.007587f
C521 B.n468 VSUBS 0.007587f
C522 B.n469 VSUBS 0.007587f
C523 B.n470 VSUBS 0.007587f
C524 B.n471 VSUBS 0.007587f
C525 B.n472 VSUBS 0.007587f
C526 B.n473 VSUBS 0.007587f
C527 B.n474 VSUBS 0.007587f
C528 B.n475 VSUBS 0.007587f
C529 B.n476 VSUBS 0.007587f
C530 B.n477 VSUBS 0.007587f
C531 B.n478 VSUBS 0.007587f
C532 B.n479 VSUBS 0.007587f
C533 B.n480 VSUBS 0.007587f
C534 B.n481 VSUBS 0.007587f
C535 B.n482 VSUBS 0.007587f
C536 B.n483 VSUBS 0.007587f
C537 B.n484 VSUBS 0.007587f
C538 B.n485 VSUBS 0.007587f
C539 B.n486 VSUBS 0.007587f
C540 B.n487 VSUBS 0.007587f
C541 B.n488 VSUBS 0.007587f
C542 B.n489 VSUBS 0.007587f
C543 B.n490 VSUBS 0.007587f
C544 B.n491 VSUBS 0.007587f
C545 B.n492 VSUBS 0.007587f
C546 B.n493 VSUBS 0.007587f
C547 B.n494 VSUBS 0.007587f
C548 B.n495 VSUBS 0.007587f
C549 B.n496 VSUBS 0.007587f
C550 B.n497 VSUBS 0.007587f
C551 B.n498 VSUBS 0.007587f
C552 B.n499 VSUBS 0.007587f
C553 B.n500 VSUBS 0.007141f
C554 B.n501 VSUBS 0.007587f
C555 B.n502 VSUBS 0.007587f
C556 B.n503 VSUBS 0.007587f
C557 B.n504 VSUBS 0.007587f
C558 B.n505 VSUBS 0.007587f
C559 B.n506 VSUBS 0.007587f
C560 B.n507 VSUBS 0.007587f
C561 B.n508 VSUBS 0.007587f
C562 B.n509 VSUBS 0.007587f
C563 B.n510 VSUBS 0.007587f
C564 B.n511 VSUBS 0.007587f
C565 B.n512 VSUBS 0.007587f
C566 B.n513 VSUBS 0.007587f
C567 B.n514 VSUBS 0.007587f
C568 B.n515 VSUBS 0.007587f
C569 B.n516 VSUBS 0.00424f
C570 B.n517 VSUBS 0.017578f
C571 B.n518 VSUBS 0.007141f
C572 B.n519 VSUBS 0.007587f
C573 B.n520 VSUBS 0.007587f
C574 B.n521 VSUBS 0.007587f
C575 B.n522 VSUBS 0.007587f
C576 B.n523 VSUBS 0.007587f
C577 B.n524 VSUBS 0.007587f
C578 B.n525 VSUBS 0.007587f
C579 B.n526 VSUBS 0.007587f
C580 B.n527 VSUBS 0.007587f
C581 B.n528 VSUBS 0.007587f
C582 B.n529 VSUBS 0.007587f
C583 B.n530 VSUBS 0.007587f
C584 B.n531 VSUBS 0.007587f
C585 B.n532 VSUBS 0.007587f
C586 B.n533 VSUBS 0.007587f
C587 B.n534 VSUBS 0.007587f
C588 B.n535 VSUBS 0.007587f
C589 B.n536 VSUBS 0.007587f
C590 B.n537 VSUBS 0.007587f
C591 B.n538 VSUBS 0.007587f
C592 B.n539 VSUBS 0.007587f
C593 B.n540 VSUBS 0.007587f
C594 B.n541 VSUBS 0.007587f
C595 B.n542 VSUBS 0.007587f
C596 B.n543 VSUBS 0.007587f
C597 B.n544 VSUBS 0.007587f
C598 B.n545 VSUBS 0.007587f
C599 B.n546 VSUBS 0.007587f
C600 B.n547 VSUBS 0.007587f
C601 B.n548 VSUBS 0.007587f
C602 B.n549 VSUBS 0.007587f
C603 B.n550 VSUBS 0.007587f
C604 B.n551 VSUBS 0.007587f
C605 B.n552 VSUBS 0.007587f
C606 B.n553 VSUBS 0.007587f
C607 B.n554 VSUBS 0.007587f
C608 B.n555 VSUBS 0.007587f
C609 B.n556 VSUBS 0.007587f
C610 B.n557 VSUBS 0.007587f
C611 B.n558 VSUBS 0.007587f
C612 B.n559 VSUBS 0.007587f
C613 B.n560 VSUBS 0.007587f
C614 B.n561 VSUBS 0.007587f
C615 B.n562 VSUBS 0.007587f
C616 B.n563 VSUBS 0.007587f
C617 B.n564 VSUBS 0.007587f
C618 B.n565 VSUBS 0.007587f
C619 B.n566 VSUBS 0.007587f
C620 B.n567 VSUBS 0.007587f
C621 B.n568 VSUBS 0.007587f
C622 B.n569 VSUBS 0.007587f
C623 B.n570 VSUBS 0.007587f
C624 B.n571 VSUBS 0.007587f
C625 B.n572 VSUBS 0.007587f
C626 B.n573 VSUBS 0.007587f
C627 B.n574 VSUBS 0.007587f
C628 B.n575 VSUBS 0.007587f
C629 B.n576 VSUBS 0.007587f
C630 B.n577 VSUBS 0.007587f
C631 B.n578 VSUBS 0.007587f
C632 B.n579 VSUBS 0.007587f
C633 B.n580 VSUBS 0.007587f
C634 B.n581 VSUBS 0.007587f
C635 B.n582 VSUBS 0.007587f
C636 B.n583 VSUBS 0.007587f
C637 B.n584 VSUBS 0.007587f
C638 B.n585 VSUBS 0.007587f
C639 B.n586 VSUBS 0.007587f
C640 B.n587 VSUBS 0.007587f
C641 B.n588 VSUBS 0.007587f
C642 B.n589 VSUBS 0.007587f
C643 B.n590 VSUBS 0.007587f
C644 B.n591 VSUBS 0.007587f
C645 B.n592 VSUBS 0.007587f
C646 B.n593 VSUBS 0.007587f
C647 B.n594 VSUBS 0.019298f
C648 B.n595 VSUBS 0.019298f
C649 B.n596 VSUBS 0.01819f
C650 B.n597 VSUBS 0.007587f
C651 B.n598 VSUBS 0.007587f
C652 B.n599 VSUBS 0.007587f
C653 B.n600 VSUBS 0.007587f
C654 B.n601 VSUBS 0.007587f
C655 B.n602 VSUBS 0.007587f
C656 B.n603 VSUBS 0.007587f
C657 B.n604 VSUBS 0.007587f
C658 B.n605 VSUBS 0.007587f
C659 B.n606 VSUBS 0.007587f
C660 B.n607 VSUBS 0.007587f
C661 B.n608 VSUBS 0.007587f
C662 B.n609 VSUBS 0.007587f
C663 B.n610 VSUBS 0.007587f
C664 B.n611 VSUBS 0.007587f
C665 B.n612 VSUBS 0.007587f
C666 B.n613 VSUBS 0.007587f
C667 B.n614 VSUBS 0.007587f
C668 B.n615 VSUBS 0.007587f
C669 B.n616 VSUBS 0.007587f
C670 B.n617 VSUBS 0.007587f
C671 B.n618 VSUBS 0.007587f
C672 B.n619 VSUBS 0.007587f
C673 B.n620 VSUBS 0.007587f
C674 B.n621 VSUBS 0.007587f
C675 B.n622 VSUBS 0.007587f
C676 B.n623 VSUBS 0.0099f
C677 B.n624 VSUBS 0.010546f
C678 B.n625 VSUBS 0.020973f
C679 VDD1.t1 VSUBS 0.336233f
C680 VDD1.t3 VSUBS 0.336233f
C681 VDD1.n0 VSUBS 2.72194f
C682 VDD1.t0 VSUBS 0.336233f
C683 VDD1.t2 VSUBS 0.336233f
C684 VDD1.n1 VSUBS 3.55223f
C685 VTAIL.n0 VSUBS 0.025224f
C686 VTAIL.n1 VSUBS 0.022268f
C687 VTAIL.n2 VSUBS 0.011966f
C688 VTAIL.n3 VSUBS 0.028282f
C689 VTAIL.n4 VSUBS 0.012669f
C690 VTAIL.n5 VSUBS 0.022268f
C691 VTAIL.n6 VSUBS 0.011966f
C692 VTAIL.n7 VSUBS 0.028282f
C693 VTAIL.n8 VSUBS 0.012669f
C694 VTAIL.n9 VSUBS 0.022268f
C695 VTAIL.n10 VSUBS 0.011966f
C696 VTAIL.n11 VSUBS 0.028282f
C697 VTAIL.n12 VSUBS 0.012669f
C698 VTAIL.n13 VSUBS 0.022268f
C699 VTAIL.n14 VSUBS 0.011966f
C700 VTAIL.n15 VSUBS 0.028282f
C701 VTAIL.n16 VSUBS 0.012318f
C702 VTAIL.n17 VSUBS 0.022268f
C703 VTAIL.n18 VSUBS 0.012669f
C704 VTAIL.n19 VSUBS 0.028282f
C705 VTAIL.n20 VSUBS 0.012669f
C706 VTAIL.n21 VSUBS 0.022268f
C707 VTAIL.n22 VSUBS 0.011966f
C708 VTAIL.n23 VSUBS 0.028282f
C709 VTAIL.n24 VSUBS 0.012669f
C710 VTAIL.n25 VSUBS 1.4463f
C711 VTAIL.n26 VSUBS 0.011966f
C712 VTAIL.t2 VSUBS 0.061215f
C713 VTAIL.n27 VSUBS 0.211715f
C714 VTAIL.n28 VSUBS 0.021275f
C715 VTAIL.n29 VSUBS 0.021212f
C716 VTAIL.n30 VSUBS 0.028282f
C717 VTAIL.n31 VSUBS 0.012669f
C718 VTAIL.n32 VSUBS 0.011966f
C719 VTAIL.n33 VSUBS 0.022268f
C720 VTAIL.n34 VSUBS 0.022268f
C721 VTAIL.n35 VSUBS 0.011966f
C722 VTAIL.n36 VSUBS 0.012669f
C723 VTAIL.n37 VSUBS 0.028282f
C724 VTAIL.n38 VSUBS 0.028282f
C725 VTAIL.n39 VSUBS 0.012669f
C726 VTAIL.n40 VSUBS 0.011966f
C727 VTAIL.n41 VSUBS 0.022268f
C728 VTAIL.n42 VSUBS 0.022268f
C729 VTAIL.n43 VSUBS 0.011966f
C730 VTAIL.n44 VSUBS 0.011966f
C731 VTAIL.n45 VSUBS 0.012669f
C732 VTAIL.n46 VSUBS 0.028282f
C733 VTAIL.n47 VSUBS 0.028282f
C734 VTAIL.n48 VSUBS 0.028282f
C735 VTAIL.n49 VSUBS 0.012318f
C736 VTAIL.n50 VSUBS 0.011966f
C737 VTAIL.n51 VSUBS 0.022268f
C738 VTAIL.n52 VSUBS 0.022268f
C739 VTAIL.n53 VSUBS 0.011966f
C740 VTAIL.n54 VSUBS 0.012669f
C741 VTAIL.n55 VSUBS 0.028282f
C742 VTAIL.n56 VSUBS 0.028282f
C743 VTAIL.n57 VSUBS 0.012669f
C744 VTAIL.n58 VSUBS 0.011966f
C745 VTAIL.n59 VSUBS 0.022268f
C746 VTAIL.n60 VSUBS 0.022268f
C747 VTAIL.n61 VSUBS 0.011966f
C748 VTAIL.n62 VSUBS 0.012669f
C749 VTAIL.n63 VSUBS 0.028282f
C750 VTAIL.n64 VSUBS 0.028282f
C751 VTAIL.n65 VSUBS 0.012669f
C752 VTAIL.n66 VSUBS 0.011966f
C753 VTAIL.n67 VSUBS 0.022268f
C754 VTAIL.n68 VSUBS 0.022268f
C755 VTAIL.n69 VSUBS 0.011966f
C756 VTAIL.n70 VSUBS 0.012669f
C757 VTAIL.n71 VSUBS 0.028282f
C758 VTAIL.n72 VSUBS 0.028282f
C759 VTAIL.n73 VSUBS 0.012669f
C760 VTAIL.n74 VSUBS 0.011966f
C761 VTAIL.n75 VSUBS 0.022268f
C762 VTAIL.n76 VSUBS 0.022268f
C763 VTAIL.n77 VSUBS 0.011966f
C764 VTAIL.n78 VSUBS 0.012669f
C765 VTAIL.n79 VSUBS 0.028282f
C766 VTAIL.n80 VSUBS 0.071045f
C767 VTAIL.n81 VSUBS 0.012669f
C768 VTAIL.n82 VSUBS 0.011966f
C769 VTAIL.n83 VSUBS 0.048124f
C770 VTAIL.n84 VSUBS 0.035736f
C771 VTAIL.n85 VSUBS 0.095842f
C772 VTAIL.n86 VSUBS 0.025224f
C773 VTAIL.n87 VSUBS 0.022268f
C774 VTAIL.n88 VSUBS 0.011966f
C775 VTAIL.n89 VSUBS 0.028282f
C776 VTAIL.n90 VSUBS 0.012669f
C777 VTAIL.n91 VSUBS 0.022268f
C778 VTAIL.n92 VSUBS 0.011966f
C779 VTAIL.n93 VSUBS 0.028282f
C780 VTAIL.n94 VSUBS 0.012669f
C781 VTAIL.n95 VSUBS 0.022268f
C782 VTAIL.n96 VSUBS 0.011966f
C783 VTAIL.n97 VSUBS 0.028282f
C784 VTAIL.n98 VSUBS 0.012669f
C785 VTAIL.n99 VSUBS 0.022268f
C786 VTAIL.n100 VSUBS 0.011966f
C787 VTAIL.n101 VSUBS 0.028282f
C788 VTAIL.n102 VSUBS 0.012318f
C789 VTAIL.n103 VSUBS 0.022268f
C790 VTAIL.n104 VSUBS 0.012669f
C791 VTAIL.n105 VSUBS 0.028282f
C792 VTAIL.n106 VSUBS 0.012669f
C793 VTAIL.n107 VSUBS 0.022268f
C794 VTAIL.n108 VSUBS 0.011966f
C795 VTAIL.n109 VSUBS 0.028282f
C796 VTAIL.n110 VSUBS 0.012669f
C797 VTAIL.n111 VSUBS 1.4463f
C798 VTAIL.n112 VSUBS 0.011966f
C799 VTAIL.t7 VSUBS 0.061215f
C800 VTAIL.n113 VSUBS 0.211715f
C801 VTAIL.n114 VSUBS 0.021275f
C802 VTAIL.n115 VSUBS 0.021212f
C803 VTAIL.n116 VSUBS 0.028282f
C804 VTAIL.n117 VSUBS 0.012669f
C805 VTAIL.n118 VSUBS 0.011966f
C806 VTAIL.n119 VSUBS 0.022268f
C807 VTAIL.n120 VSUBS 0.022268f
C808 VTAIL.n121 VSUBS 0.011966f
C809 VTAIL.n122 VSUBS 0.012669f
C810 VTAIL.n123 VSUBS 0.028282f
C811 VTAIL.n124 VSUBS 0.028282f
C812 VTAIL.n125 VSUBS 0.012669f
C813 VTAIL.n126 VSUBS 0.011966f
C814 VTAIL.n127 VSUBS 0.022268f
C815 VTAIL.n128 VSUBS 0.022268f
C816 VTAIL.n129 VSUBS 0.011966f
C817 VTAIL.n130 VSUBS 0.011966f
C818 VTAIL.n131 VSUBS 0.012669f
C819 VTAIL.n132 VSUBS 0.028282f
C820 VTAIL.n133 VSUBS 0.028282f
C821 VTAIL.n134 VSUBS 0.028282f
C822 VTAIL.n135 VSUBS 0.012318f
C823 VTAIL.n136 VSUBS 0.011966f
C824 VTAIL.n137 VSUBS 0.022268f
C825 VTAIL.n138 VSUBS 0.022268f
C826 VTAIL.n139 VSUBS 0.011966f
C827 VTAIL.n140 VSUBS 0.012669f
C828 VTAIL.n141 VSUBS 0.028282f
C829 VTAIL.n142 VSUBS 0.028282f
C830 VTAIL.n143 VSUBS 0.012669f
C831 VTAIL.n144 VSUBS 0.011966f
C832 VTAIL.n145 VSUBS 0.022268f
C833 VTAIL.n146 VSUBS 0.022268f
C834 VTAIL.n147 VSUBS 0.011966f
C835 VTAIL.n148 VSUBS 0.012669f
C836 VTAIL.n149 VSUBS 0.028282f
C837 VTAIL.n150 VSUBS 0.028282f
C838 VTAIL.n151 VSUBS 0.012669f
C839 VTAIL.n152 VSUBS 0.011966f
C840 VTAIL.n153 VSUBS 0.022268f
C841 VTAIL.n154 VSUBS 0.022268f
C842 VTAIL.n155 VSUBS 0.011966f
C843 VTAIL.n156 VSUBS 0.012669f
C844 VTAIL.n157 VSUBS 0.028282f
C845 VTAIL.n158 VSUBS 0.028282f
C846 VTAIL.n159 VSUBS 0.012669f
C847 VTAIL.n160 VSUBS 0.011966f
C848 VTAIL.n161 VSUBS 0.022268f
C849 VTAIL.n162 VSUBS 0.022268f
C850 VTAIL.n163 VSUBS 0.011966f
C851 VTAIL.n164 VSUBS 0.012669f
C852 VTAIL.n165 VSUBS 0.028282f
C853 VTAIL.n166 VSUBS 0.071045f
C854 VTAIL.n167 VSUBS 0.012669f
C855 VTAIL.n168 VSUBS 0.011966f
C856 VTAIL.n169 VSUBS 0.048124f
C857 VTAIL.n170 VSUBS 0.035736f
C858 VTAIL.n171 VSUBS 0.132491f
C859 VTAIL.n172 VSUBS 0.025224f
C860 VTAIL.n173 VSUBS 0.022268f
C861 VTAIL.n174 VSUBS 0.011966f
C862 VTAIL.n175 VSUBS 0.028282f
C863 VTAIL.n176 VSUBS 0.012669f
C864 VTAIL.n177 VSUBS 0.022268f
C865 VTAIL.n178 VSUBS 0.011966f
C866 VTAIL.n179 VSUBS 0.028282f
C867 VTAIL.n180 VSUBS 0.012669f
C868 VTAIL.n181 VSUBS 0.022268f
C869 VTAIL.n182 VSUBS 0.011966f
C870 VTAIL.n183 VSUBS 0.028282f
C871 VTAIL.n184 VSUBS 0.012669f
C872 VTAIL.n185 VSUBS 0.022268f
C873 VTAIL.n186 VSUBS 0.011966f
C874 VTAIL.n187 VSUBS 0.028282f
C875 VTAIL.n188 VSUBS 0.012318f
C876 VTAIL.n189 VSUBS 0.022268f
C877 VTAIL.n190 VSUBS 0.012669f
C878 VTAIL.n191 VSUBS 0.028282f
C879 VTAIL.n192 VSUBS 0.012669f
C880 VTAIL.n193 VSUBS 0.022268f
C881 VTAIL.n194 VSUBS 0.011966f
C882 VTAIL.n195 VSUBS 0.028282f
C883 VTAIL.n196 VSUBS 0.012669f
C884 VTAIL.n197 VSUBS 1.4463f
C885 VTAIL.n198 VSUBS 0.011966f
C886 VTAIL.t4 VSUBS 0.061215f
C887 VTAIL.n199 VSUBS 0.211715f
C888 VTAIL.n200 VSUBS 0.021275f
C889 VTAIL.n201 VSUBS 0.021212f
C890 VTAIL.n202 VSUBS 0.028282f
C891 VTAIL.n203 VSUBS 0.012669f
C892 VTAIL.n204 VSUBS 0.011966f
C893 VTAIL.n205 VSUBS 0.022268f
C894 VTAIL.n206 VSUBS 0.022268f
C895 VTAIL.n207 VSUBS 0.011966f
C896 VTAIL.n208 VSUBS 0.012669f
C897 VTAIL.n209 VSUBS 0.028282f
C898 VTAIL.n210 VSUBS 0.028282f
C899 VTAIL.n211 VSUBS 0.012669f
C900 VTAIL.n212 VSUBS 0.011966f
C901 VTAIL.n213 VSUBS 0.022268f
C902 VTAIL.n214 VSUBS 0.022268f
C903 VTAIL.n215 VSUBS 0.011966f
C904 VTAIL.n216 VSUBS 0.011966f
C905 VTAIL.n217 VSUBS 0.012669f
C906 VTAIL.n218 VSUBS 0.028282f
C907 VTAIL.n219 VSUBS 0.028282f
C908 VTAIL.n220 VSUBS 0.028282f
C909 VTAIL.n221 VSUBS 0.012318f
C910 VTAIL.n222 VSUBS 0.011966f
C911 VTAIL.n223 VSUBS 0.022268f
C912 VTAIL.n224 VSUBS 0.022268f
C913 VTAIL.n225 VSUBS 0.011966f
C914 VTAIL.n226 VSUBS 0.012669f
C915 VTAIL.n227 VSUBS 0.028282f
C916 VTAIL.n228 VSUBS 0.028282f
C917 VTAIL.n229 VSUBS 0.012669f
C918 VTAIL.n230 VSUBS 0.011966f
C919 VTAIL.n231 VSUBS 0.022268f
C920 VTAIL.n232 VSUBS 0.022268f
C921 VTAIL.n233 VSUBS 0.011966f
C922 VTAIL.n234 VSUBS 0.012669f
C923 VTAIL.n235 VSUBS 0.028282f
C924 VTAIL.n236 VSUBS 0.028282f
C925 VTAIL.n237 VSUBS 0.012669f
C926 VTAIL.n238 VSUBS 0.011966f
C927 VTAIL.n239 VSUBS 0.022268f
C928 VTAIL.n240 VSUBS 0.022268f
C929 VTAIL.n241 VSUBS 0.011966f
C930 VTAIL.n242 VSUBS 0.012669f
C931 VTAIL.n243 VSUBS 0.028282f
C932 VTAIL.n244 VSUBS 0.028282f
C933 VTAIL.n245 VSUBS 0.012669f
C934 VTAIL.n246 VSUBS 0.011966f
C935 VTAIL.n247 VSUBS 0.022268f
C936 VTAIL.n248 VSUBS 0.022268f
C937 VTAIL.n249 VSUBS 0.011966f
C938 VTAIL.n250 VSUBS 0.012669f
C939 VTAIL.n251 VSUBS 0.028282f
C940 VTAIL.n252 VSUBS 0.071045f
C941 VTAIL.n253 VSUBS 0.012669f
C942 VTAIL.n254 VSUBS 0.011966f
C943 VTAIL.n255 VSUBS 0.048124f
C944 VTAIL.n256 VSUBS 0.035736f
C945 VTAIL.n257 VSUBS 1.44845f
C946 VTAIL.n258 VSUBS 0.025224f
C947 VTAIL.n259 VSUBS 0.022268f
C948 VTAIL.n260 VSUBS 0.011966f
C949 VTAIL.n261 VSUBS 0.028282f
C950 VTAIL.n262 VSUBS 0.012669f
C951 VTAIL.n263 VSUBS 0.022268f
C952 VTAIL.n264 VSUBS 0.011966f
C953 VTAIL.n265 VSUBS 0.028282f
C954 VTAIL.n266 VSUBS 0.012669f
C955 VTAIL.n267 VSUBS 0.022268f
C956 VTAIL.n268 VSUBS 0.011966f
C957 VTAIL.n269 VSUBS 0.028282f
C958 VTAIL.n270 VSUBS 0.012669f
C959 VTAIL.n271 VSUBS 0.022268f
C960 VTAIL.n272 VSUBS 0.011966f
C961 VTAIL.n273 VSUBS 0.028282f
C962 VTAIL.n274 VSUBS 0.012318f
C963 VTAIL.n275 VSUBS 0.022268f
C964 VTAIL.n276 VSUBS 0.012318f
C965 VTAIL.n277 VSUBS 0.011966f
C966 VTAIL.n278 VSUBS 0.028282f
C967 VTAIL.n279 VSUBS 0.028282f
C968 VTAIL.n280 VSUBS 0.012669f
C969 VTAIL.n281 VSUBS 0.022268f
C970 VTAIL.n282 VSUBS 0.011966f
C971 VTAIL.n283 VSUBS 0.028282f
C972 VTAIL.n284 VSUBS 0.012669f
C973 VTAIL.n285 VSUBS 1.4463f
C974 VTAIL.n286 VSUBS 0.011966f
C975 VTAIL.t1 VSUBS 0.061215f
C976 VTAIL.n287 VSUBS 0.211715f
C977 VTAIL.n288 VSUBS 0.021275f
C978 VTAIL.n289 VSUBS 0.021212f
C979 VTAIL.n290 VSUBS 0.028282f
C980 VTAIL.n291 VSUBS 0.012669f
C981 VTAIL.n292 VSUBS 0.011966f
C982 VTAIL.n293 VSUBS 0.022268f
C983 VTAIL.n294 VSUBS 0.022268f
C984 VTAIL.n295 VSUBS 0.011966f
C985 VTAIL.n296 VSUBS 0.012669f
C986 VTAIL.n297 VSUBS 0.028282f
C987 VTAIL.n298 VSUBS 0.028282f
C988 VTAIL.n299 VSUBS 0.012669f
C989 VTAIL.n300 VSUBS 0.011966f
C990 VTAIL.n301 VSUBS 0.022268f
C991 VTAIL.n302 VSUBS 0.022268f
C992 VTAIL.n303 VSUBS 0.011966f
C993 VTAIL.n304 VSUBS 0.012669f
C994 VTAIL.n305 VSUBS 0.028282f
C995 VTAIL.n306 VSUBS 0.028282f
C996 VTAIL.n307 VSUBS 0.012669f
C997 VTAIL.n308 VSUBS 0.011966f
C998 VTAIL.n309 VSUBS 0.022268f
C999 VTAIL.n310 VSUBS 0.022268f
C1000 VTAIL.n311 VSUBS 0.011966f
C1001 VTAIL.n312 VSUBS 0.012669f
C1002 VTAIL.n313 VSUBS 0.028282f
C1003 VTAIL.n314 VSUBS 0.028282f
C1004 VTAIL.n315 VSUBS 0.012669f
C1005 VTAIL.n316 VSUBS 0.011966f
C1006 VTAIL.n317 VSUBS 0.022268f
C1007 VTAIL.n318 VSUBS 0.022268f
C1008 VTAIL.n319 VSUBS 0.011966f
C1009 VTAIL.n320 VSUBS 0.012669f
C1010 VTAIL.n321 VSUBS 0.028282f
C1011 VTAIL.n322 VSUBS 0.028282f
C1012 VTAIL.n323 VSUBS 0.012669f
C1013 VTAIL.n324 VSUBS 0.011966f
C1014 VTAIL.n325 VSUBS 0.022268f
C1015 VTAIL.n326 VSUBS 0.022268f
C1016 VTAIL.n327 VSUBS 0.011966f
C1017 VTAIL.n328 VSUBS 0.012669f
C1018 VTAIL.n329 VSUBS 0.028282f
C1019 VTAIL.n330 VSUBS 0.028282f
C1020 VTAIL.n331 VSUBS 0.012669f
C1021 VTAIL.n332 VSUBS 0.011966f
C1022 VTAIL.n333 VSUBS 0.022268f
C1023 VTAIL.n334 VSUBS 0.022268f
C1024 VTAIL.n335 VSUBS 0.011966f
C1025 VTAIL.n336 VSUBS 0.012669f
C1026 VTAIL.n337 VSUBS 0.028282f
C1027 VTAIL.n338 VSUBS 0.071045f
C1028 VTAIL.n339 VSUBS 0.012669f
C1029 VTAIL.n340 VSUBS 0.011966f
C1030 VTAIL.n341 VSUBS 0.048124f
C1031 VTAIL.n342 VSUBS 0.035736f
C1032 VTAIL.n343 VSUBS 1.44845f
C1033 VTAIL.n344 VSUBS 0.025224f
C1034 VTAIL.n345 VSUBS 0.022268f
C1035 VTAIL.n346 VSUBS 0.011966f
C1036 VTAIL.n347 VSUBS 0.028282f
C1037 VTAIL.n348 VSUBS 0.012669f
C1038 VTAIL.n349 VSUBS 0.022268f
C1039 VTAIL.n350 VSUBS 0.011966f
C1040 VTAIL.n351 VSUBS 0.028282f
C1041 VTAIL.n352 VSUBS 0.012669f
C1042 VTAIL.n353 VSUBS 0.022268f
C1043 VTAIL.n354 VSUBS 0.011966f
C1044 VTAIL.n355 VSUBS 0.028282f
C1045 VTAIL.n356 VSUBS 0.012669f
C1046 VTAIL.n357 VSUBS 0.022268f
C1047 VTAIL.n358 VSUBS 0.011966f
C1048 VTAIL.n359 VSUBS 0.028282f
C1049 VTAIL.n360 VSUBS 0.012318f
C1050 VTAIL.n361 VSUBS 0.022268f
C1051 VTAIL.n362 VSUBS 0.012318f
C1052 VTAIL.n363 VSUBS 0.011966f
C1053 VTAIL.n364 VSUBS 0.028282f
C1054 VTAIL.n365 VSUBS 0.028282f
C1055 VTAIL.n366 VSUBS 0.012669f
C1056 VTAIL.n367 VSUBS 0.022268f
C1057 VTAIL.n368 VSUBS 0.011966f
C1058 VTAIL.n369 VSUBS 0.028282f
C1059 VTAIL.n370 VSUBS 0.012669f
C1060 VTAIL.n371 VSUBS 1.4463f
C1061 VTAIL.n372 VSUBS 0.011966f
C1062 VTAIL.t0 VSUBS 0.061215f
C1063 VTAIL.n373 VSUBS 0.211715f
C1064 VTAIL.n374 VSUBS 0.021275f
C1065 VTAIL.n375 VSUBS 0.021212f
C1066 VTAIL.n376 VSUBS 0.028282f
C1067 VTAIL.n377 VSUBS 0.012669f
C1068 VTAIL.n378 VSUBS 0.011966f
C1069 VTAIL.n379 VSUBS 0.022268f
C1070 VTAIL.n380 VSUBS 0.022268f
C1071 VTAIL.n381 VSUBS 0.011966f
C1072 VTAIL.n382 VSUBS 0.012669f
C1073 VTAIL.n383 VSUBS 0.028282f
C1074 VTAIL.n384 VSUBS 0.028282f
C1075 VTAIL.n385 VSUBS 0.012669f
C1076 VTAIL.n386 VSUBS 0.011966f
C1077 VTAIL.n387 VSUBS 0.022268f
C1078 VTAIL.n388 VSUBS 0.022268f
C1079 VTAIL.n389 VSUBS 0.011966f
C1080 VTAIL.n390 VSUBS 0.012669f
C1081 VTAIL.n391 VSUBS 0.028282f
C1082 VTAIL.n392 VSUBS 0.028282f
C1083 VTAIL.n393 VSUBS 0.012669f
C1084 VTAIL.n394 VSUBS 0.011966f
C1085 VTAIL.n395 VSUBS 0.022268f
C1086 VTAIL.n396 VSUBS 0.022268f
C1087 VTAIL.n397 VSUBS 0.011966f
C1088 VTAIL.n398 VSUBS 0.012669f
C1089 VTAIL.n399 VSUBS 0.028282f
C1090 VTAIL.n400 VSUBS 0.028282f
C1091 VTAIL.n401 VSUBS 0.012669f
C1092 VTAIL.n402 VSUBS 0.011966f
C1093 VTAIL.n403 VSUBS 0.022268f
C1094 VTAIL.n404 VSUBS 0.022268f
C1095 VTAIL.n405 VSUBS 0.011966f
C1096 VTAIL.n406 VSUBS 0.012669f
C1097 VTAIL.n407 VSUBS 0.028282f
C1098 VTAIL.n408 VSUBS 0.028282f
C1099 VTAIL.n409 VSUBS 0.012669f
C1100 VTAIL.n410 VSUBS 0.011966f
C1101 VTAIL.n411 VSUBS 0.022268f
C1102 VTAIL.n412 VSUBS 0.022268f
C1103 VTAIL.n413 VSUBS 0.011966f
C1104 VTAIL.n414 VSUBS 0.012669f
C1105 VTAIL.n415 VSUBS 0.028282f
C1106 VTAIL.n416 VSUBS 0.028282f
C1107 VTAIL.n417 VSUBS 0.012669f
C1108 VTAIL.n418 VSUBS 0.011966f
C1109 VTAIL.n419 VSUBS 0.022268f
C1110 VTAIL.n420 VSUBS 0.022268f
C1111 VTAIL.n421 VSUBS 0.011966f
C1112 VTAIL.n422 VSUBS 0.012669f
C1113 VTAIL.n423 VSUBS 0.028282f
C1114 VTAIL.n424 VSUBS 0.071045f
C1115 VTAIL.n425 VSUBS 0.012669f
C1116 VTAIL.n426 VSUBS 0.011966f
C1117 VTAIL.n427 VSUBS 0.048124f
C1118 VTAIL.n428 VSUBS 0.035736f
C1119 VTAIL.n429 VSUBS 0.132491f
C1120 VTAIL.n430 VSUBS 0.025224f
C1121 VTAIL.n431 VSUBS 0.022268f
C1122 VTAIL.n432 VSUBS 0.011966f
C1123 VTAIL.n433 VSUBS 0.028282f
C1124 VTAIL.n434 VSUBS 0.012669f
C1125 VTAIL.n435 VSUBS 0.022268f
C1126 VTAIL.n436 VSUBS 0.011966f
C1127 VTAIL.n437 VSUBS 0.028282f
C1128 VTAIL.n438 VSUBS 0.012669f
C1129 VTAIL.n439 VSUBS 0.022268f
C1130 VTAIL.n440 VSUBS 0.011966f
C1131 VTAIL.n441 VSUBS 0.028282f
C1132 VTAIL.n442 VSUBS 0.012669f
C1133 VTAIL.n443 VSUBS 0.022268f
C1134 VTAIL.n444 VSUBS 0.011966f
C1135 VTAIL.n445 VSUBS 0.028282f
C1136 VTAIL.n446 VSUBS 0.012318f
C1137 VTAIL.n447 VSUBS 0.022268f
C1138 VTAIL.n448 VSUBS 0.012318f
C1139 VTAIL.n449 VSUBS 0.011966f
C1140 VTAIL.n450 VSUBS 0.028282f
C1141 VTAIL.n451 VSUBS 0.028282f
C1142 VTAIL.n452 VSUBS 0.012669f
C1143 VTAIL.n453 VSUBS 0.022268f
C1144 VTAIL.n454 VSUBS 0.011966f
C1145 VTAIL.n455 VSUBS 0.028282f
C1146 VTAIL.n456 VSUBS 0.012669f
C1147 VTAIL.n457 VSUBS 1.4463f
C1148 VTAIL.n458 VSUBS 0.011966f
C1149 VTAIL.t5 VSUBS 0.061215f
C1150 VTAIL.n459 VSUBS 0.211715f
C1151 VTAIL.n460 VSUBS 0.021275f
C1152 VTAIL.n461 VSUBS 0.021212f
C1153 VTAIL.n462 VSUBS 0.028282f
C1154 VTAIL.n463 VSUBS 0.012669f
C1155 VTAIL.n464 VSUBS 0.011966f
C1156 VTAIL.n465 VSUBS 0.022268f
C1157 VTAIL.n466 VSUBS 0.022268f
C1158 VTAIL.n467 VSUBS 0.011966f
C1159 VTAIL.n468 VSUBS 0.012669f
C1160 VTAIL.n469 VSUBS 0.028282f
C1161 VTAIL.n470 VSUBS 0.028282f
C1162 VTAIL.n471 VSUBS 0.012669f
C1163 VTAIL.n472 VSUBS 0.011966f
C1164 VTAIL.n473 VSUBS 0.022268f
C1165 VTAIL.n474 VSUBS 0.022268f
C1166 VTAIL.n475 VSUBS 0.011966f
C1167 VTAIL.n476 VSUBS 0.012669f
C1168 VTAIL.n477 VSUBS 0.028282f
C1169 VTAIL.n478 VSUBS 0.028282f
C1170 VTAIL.n479 VSUBS 0.012669f
C1171 VTAIL.n480 VSUBS 0.011966f
C1172 VTAIL.n481 VSUBS 0.022268f
C1173 VTAIL.n482 VSUBS 0.022268f
C1174 VTAIL.n483 VSUBS 0.011966f
C1175 VTAIL.n484 VSUBS 0.012669f
C1176 VTAIL.n485 VSUBS 0.028282f
C1177 VTAIL.n486 VSUBS 0.028282f
C1178 VTAIL.n487 VSUBS 0.012669f
C1179 VTAIL.n488 VSUBS 0.011966f
C1180 VTAIL.n489 VSUBS 0.022268f
C1181 VTAIL.n490 VSUBS 0.022268f
C1182 VTAIL.n491 VSUBS 0.011966f
C1183 VTAIL.n492 VSUBS 0.012669f
C1184 VTAIL.n493 VSUBS 0.028282f
C1185 VTAIL.n494 VSUBS 0.028282f
C1186 VTAIL.n495 VSUBS 0.012669f
C1187 VTAIL.n496 VSUBS 0.011966f
C1188 VTAIL.n497 VSUBS 0.022268f
C1189 VTAIL.n498 VSUBS 0.022268f
C1190 VTAIL.n499 VSUBS 0.011966f
C1191 VTAIL.n500 VSUBS 0.012669f
C1192 VTAIL.n501 VSUBS 0.028282f
C1193 VTAIL.n502 VSUBS 0.028282f
C1194 VTAIL.n503 VSUBS 0.012669f
C1195 VTAIL.n504 VSUBS 0.011966f
C1196 VTAIL.n505 VSUBS 0.022268f
C1197 VTAIL.n506 VSUBS 0.022268f
C1198 VTAIL.n507 VSUBS 0.011966f
C1199 VTAIL.n508 VSUBS 0.012669f
C1200 VTAIL.n509 VSUBS 0.028282f
C1201 VTAIL.n510 VSUBS 0.071045f
C1202 VTAIL.n511 VSUBS 0.012669f
C1203 VTAIL.n512 VSUBS 0.011966f
C1204 VTAIL.n513 VSUBS 0.048124f
C1205 VTAIL.n514 VSUBS 0.035736f
C1206 VTAIL.n515 VSUBS 0.132491f
C1207 VTAIL.n516 VSUBS 0.025224f
C1208 VTAIL.n517 VSUBS 0.022268f
C1209 VTAIL.n518 VSUBS 0.011966f
C1210 VTAIL.n519 VSUBS 0.028282f
C1211 VTAIL.n520 VSUBS 0.012669f
C1212 VTAIL.n521 VSUBS 0.022268f
C1213 VTAIL.n522 VSUBS 0.011966f
C1214 VTAIL.n523 VSUBS 0.028282f
C1215 VTAIL.n524 VSUBS 0.012669f
C1216 VTAIL.n525 VSUBS 0.022268f
C1217 VTAIL.n526 VSUBS 0.011966f
C1218 VTAIL.n527 VSUBS 0.028282f
C1219 VTAIL.n528 VSUBS 0.012669f
C1220 VTAIL.n529 VSUBS 0.022268f
C1221 VTAIL.n530 VSUBS 0.011966f
C1222 VTAIL.n531 VSUBS 0.028282f
C1223 VTAIL.n532 VSUBS 0.012318f
C1224 VTAIL.n533 VSUBS 0.022268f
C1225 VTAIL.n534 VSUBS 0.012318f
C1226 VTAIL.n535 VSUBS 0.011966f
C1227 VTAIL.n536 VSUBS 0.028282f
C1228 VTAIL.n537 VSUBS 0.028282f
C1229 VTAIL.n538 VSUBS 0.012669f
C1230 VTAIL.n539 VSUBS 0.022268f
C1231 VTAIL.n540 VSUBS 0.011966f
C1232 VTAIL.n541 VSUBS 0.028282f
C1233 VTAIL.n542 VSUBS 0.012669f
C1234 VTAIL.n543 VSUBS 1.4463f
C1235 VTAIL.n544 VSUBS 0.011966f
C1236 VTAIL.t6 VSUBS 0.061215f
C1237 VTAIL.n545 VSUBS 0.211715f
C1238 VTAIL.n546 VSUBS 0.021275f
C1239 VTAIL.n547 VSUBS 0.021212f
C1240 VTAIL.n548 VSUBS 0.028282f
C1241 VTAIL.n549 VSUBS 0.012669f
C1242 VTAIL.n550 VSUBS 0.011966f
C1243 VTAIL.n551 VSUBS 0.022268f
C1244 VTAIL.n552 VSUBS 0.022268f
C1245 VTAIL.n553 VSUBS 0.011966f
C1246 VTAIL.n554 VSUBS 0.012669f
C1247 VTAIL.n555 VSUBS 0.028282f
C1248 VTAIL.n556 VSUBS 0.028282f
C1249 VTAIL.n557 VSUBS 0.012669f
C1250 VTAIL.n558 VSUBS 0.011966f
C1251 VTAIL.n559 VSUBS 0.022268f
C1252 VTAIL.n560 VSUBS 0.022268f
C1253 VTAIL.n561 VSUBS 0.011966f
C1254 VTAIL.n562 VSUBS 0.012669f
C1255 VTAIL.n563 VSUBS 0.028282f
C1256 VTAIL.n564 VSUBS 0.028282f
C1257 VTAIL.n565 VSUBS 0.012669f
C1258 VTAIL.n566 VSUBS 0.011966f
C1259 VTAIL.n567 VSUBS 0.022268f
C1260 VTAIL.n568 VSUBS 0.022268f
C1261 VTAIL.n569 VSUBS 0.011966f
C1262 VTAIL.n570 VSUBS 0.012669f
C1263 VTAIL.n571 VSUBS 0.028282f
C1264 VTAIL.n572 VSUBS 0.028282f
C1265 VTAIL.n573 VSUBS 0.012669f
C1266 VTAIL.n574 VSUBS 0.011966f
C1267 VTAIL.n575 VSUBS 0.022268f
C1268 VTAIL.n576 VSUBS 0.022268f
C1269 VTAIL.n577 VSUBS 0.011966f
C1270 VTAIL.n578 VSUBS 0.012669f
C1271 VTAIL.n579 VSUBS 0.028282f
C1272 VTAIL.n580 VSUBS 0.028282f
C1273 VTAIL.n581 VSUBS 0.012669f
C1274 VTAIL.n582 VSUBS 0.011966f
C1275 VTAIL.n583 VSUBS 0.022268f
C1276 VTAIL.n584 VSUBS 0.022268f
C1277 VTAIL.n585 VSUBS 0.011966f
C1278 VTAIL.n586 VSUBS 0.012669f
C1279 VTAIL.n587 VSUBS 0.028282f
C1280 VTAIL.n588 VSUBS 0.028282f
C1281 VTAIL.n589 VSUBS 0.012669f
C1282 VTAIL.n590 VSUBS 0.011966f
C1283 VTAIL.n591 VSUBS 0.022268f
C1284 VTAIL.n592 VSUBS 0.022268f
C1285 VTAIL.n593 VSUBS 0.011966f
C1286 VTAIL.n594 VSUBS 0.012669f
C1287 VTAIL.n595 VSUBS 0.028282f
C1288 VTAIL.n596 VSUBS 0.071045f
C1289 VTAIL.n597 VSUBS 0.012669f
C1290 VTAIL.n598 VSUBS 0.011966f
C1291 VTAIL.n599 VSUBS 0.048124f
C1292 VTAIL.n600 VSUBS 0.035736f
C1293 VTAIL.n601 VSUBS 1.44845f
C1294 VTAIL.n602 VSUBS 0.025224f
C1295 VTAIL.n603 VSUBS 0.022268f
C1296 VTAIL.n604 VSUBS 0.011966f
C1297 VTAIL.n605 VSUBS 0.028282f
C1298 VTAIL.n606 VSUBS 0.012669f
C1299 VTAIL.n607 VSUBS 0.022268f
C1300 VTAIL.n608 VSUBS 0.011966f
C1301 VTAIL.n609 VSUBS 0.028282f
C1302 VTAIL.n610 VSUBS 0.012669f
C1303 VTAIL.n611 VSUBS 0.022268f
C1304 VTAIL.n612 VSUBS 0.011966f
C1305 VTAIL.n613 VSUBS 0.028282f
C1306 VTAIL.n614 VSUBS 0.012669f
C1307 VTAIL.n615 VSUBS 0.022268f
C1308 VTAIL.n616 VSUBS 0.011966f
C1309 VTAIL.n617 VSUBS 0.028282f
C1310 VTAIL.n618 VSUBS 0.012318f
C1311 VTAIL.n619 VSUBS 0.022268f
C1312 VTAIL.n620 VSUBS 0.012669f
C1313 VTAIL.n621 VSUBS 0.028282f
C1314 VTAIL.n622 VSUBS 0.012669f
C1315 VTAIL.n623 VSUBS 0.022268f
C1316 VTAIL.n624 VSUBS 0.011966f
C1317 VTAIL.n625 VSUBS 0.028282f
C1318 VTAIL.n626 VSUBS 0.012669f
C1319 VTAIL.n627 VSUBS 1.4463f
C1320 VTAIL.n628 VSUBS 0.011966f
C1321 VTAIL.t3 VSUBS 0.061215f
C1322 VTAIL.n629 VSUBS 0.211715f
C1323 VTAIL.n630 VSUBS 0.021275f
C1324 VTAIL.n631 VSUBS 0.021212f
C1325 VTAIL.n632 VSUBS 0.028282f
C1326 VTAIL.n633 VSUBS 0.012669f
C1327 VTAIL.n634 VSUBS 0.011966f
C1328 VTAIL.n635 VSUBS 0.022268f
C1329 VTAIL.n636 VSUBS 0.022268f
C1330 VTAIL.n637 VSUBS 0.011966f
C1331 VTAIL.n638 VSUBS 0.012669f
C1332 VTAIL.n639 VSUBS 0.028282f
C1333 VTAIL.n640 VSUBS 0.028282f
C1334 VTAIL.n641 VSUBS 0.012669f
C1335 VTAIL.n642 VSUBS 0.011966f
C1336 VTAIL.n643 VSUBS 0.022268f
C1337 VTAIL.n644 VSUBS 0.022268f
C1338 VTAIL.n645 VSUBS 0.011966f
C1339 VTAIL.n646 VSUBS 0.011966f
C1340 VTAIL.n647 VSUBS 0.012669f
C1341 VTAIL.n648 VSUBS 0.028282f
C1342 VTAIL.n649 VSUBS 0.028282f
C1343 VTAIL.n650 VSUBS 0.028282f
C1344 VTAIL.n651 VSUBS 0.012318f
C1345 VTAIL.n652 VSUBS 0.011966f
C1346 VTAIL.n653 VSUBS 0.022268f
C1347 VTAIL.n654 VSUBS 0.022268f
C1348 VTAIL.n655 VSUBS 0.011966f
C1349 VTAIL.n656 VSUBS 0.012669f
C1350 VTAIL.n657 VSUBS 0.028282f
C1351 VTAIL.n658 VSUBS 0.028282f
C1352 VTAIL.n659 VSUBS 0.012669f
C1353 VTAIL.n660 VSUBS 0.011966f
C1354 VTAIL.n661 VSUBS 0.022268f
C1355 VTAIL.n662 VSUBS 0.022268f
C1356 VTAIL.n663 VSUBS 0.011966f
C1357 VTAIL.n664 VSUBS 0.012669f
C1358 VTAIL.n665 VSUBS 0.028282f
C1359 VTAIL.n666 VSUBS 0.028282f
C1360 VTAIL.n667 VSUBS 0.012669f
C1361 VTAIL.n668 VSUBS 0.011966f
C1362 VTAIL.n669 VSUBS 0.022268f
C1363 VTAIL.n670 VSUBS 0.022268f
C1364 VTAIL.n671 VSUBS 0.011966f
C1365 VTAIL.n672 VSUBS 0.012669f
C1366 VTAIL.n673 VSUBS 0.028282f
C1367 VTAIL.n674 VSUBS 0.028282f
C1368 VTAIL.n675 VSUBS 0.012669f
C1369 VTAIL.n676 VSUBS 0.011966f
C1370 VTAIL.n677 VSUBS 0.022268f
C1371 VTAIL.n678 VSUBS 0.022268f
C1372 VTAIL.n679 VSUBS 0.011966f
C1373 VTAIL.n680 VSUBS 0.012669f
C1374 VTAIL.n681 VSUBS 0.028282f
C1375 VTAIL.n682 VSUBS 0.071045f
C1376 VTAIL.n683 VSUBS 0.012669f
C1377 VTAIL.n684 VSUBS 0.011966f
C1378 VTAIL.n685 VSUBS 0.048124f
C1379 VTAIL.n686 VSUBS 0.035736f
C1380 VTAIL.n687 VSUBS 1.40345f
C1381 VP.t0 VSUBS 2.32695f
C1382 VP.t2 VSUBS 2.32714f
C1383 VP.n0 VSUBS 3.14478f
C1384 VP.n1 VSUBS 3.45299f
C1385 VP.t3 VSUBS 2.2899f
C1386 VP.n2 VSUBS 0.87702f
C1387 VP.t1 VSUBS 2.2899f
C1388 VP.n3 VSUBS 0.87702f
C1389 VP.n4 VSUBS 0.066292f
.ends

