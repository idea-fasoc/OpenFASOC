* NGSPICE file created from diff_pair_sample_0782.ext - technology: sky130A

.subckt diff_pair_sample_0782 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=0.63
X1 B.t8 B.t6 B.t7 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=0.63
X2 VTAIL.t11 VP.t0 VDD1.t4 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=1.96185 ps=12.22 w=11.89 l=0.63
X3 VDD2.t5 VN.t0 VTAIL.t3 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=4.6371 ps=24.56 w=11.89 l=0.63
X4 VDD2.t4 VN.t1 VTAIL.t4 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=4.6371 ps=24.56 w=11.89 l=0.63
X5 VTAIL.t5 VN.t2 VDD2.t3 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=1.96185 ps=12.22 w=11.89 l=0.63
X6 VDD2.t2 VN.t3 VTAIL.t2 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=1.96185 ps=12.22 w=11.89 l=0.63
X7 VDD2.t1 VN.t4 VTAIL.t0 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=1.96185 ps=12.22 w=11.89 l=0.63
X8 VDD1.t2 VP.t1 VTAIL.t10 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=1.96185 ps=12.22 w=11.89 l=0.63
X9 VDD1.t0 VP.t2 VTAIL.t9 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=4.6371 ps=24.56 w=11.89 l=0.63
X10 VDD1.t5 VP.t3 VTAIL.t8 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=1.96185 ps=12.22 w=11.89 l=0.63
X11 B.t5 B.t3 B.t4 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=0.63
X12 VTAIL.t7 VP.t4 VDD1.t3 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=1.96185 ps=12.22 w=11.89 l=0.63
X13 VDD1.t1 VP.t5 VTAIL.t6 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=4.6371 ps=24.56 w=11.89 l=0.63
X14 B.t2 B.t0 B.t1 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=4.6371 pd=24.56 as=0 ps=0 w=11.89 l=0.63
X15 VTAIL.t1 VN.t5 VDD2.t0 w_n1738_n3346# sky130_fd_pr__pfet_01v8 ad=1.96185 pd=12.22 as=1.96185 ps=12.22 w=11.89 l=0.63
R0 B.n108 B.t6 658.761
R1 B.n242 B.t3 658.761
R2 B.n40 B.t0 658.761
R3 B.n32 B.t9 658.761
R4 B.n307 B.n82 585
R5 B.n306 B.n305 585
R6 B.n304 B.n83 585
R7 B.n303 B.n302 585
R8 B.n301 B.n84 585
R9 B.n300 B.n299 585
R10 B.n298 B.n85 585
R11 B.n297 B.n296 585
R12 B.n295 B.n86 585
R13 B.n294 B.n293 585
R14 B.n292 B.n87 585
R15 B.n291 B.n290 585
R16 B.n289 B.n88 585
R17 B.n288 B.n287 585
R18 B.n286 B.n89 585
R19 B.n285 B.n284 585
R20 B.n283 B.n90 585
R21 B.n282 B.n281 585
R22 B.n280 B.n91 585
R23 B.n279 B.n278 585
R24 B.n277 B.n92 585
R25 B.n276 B.n275 585
R26 B.n274 B.n93 585
R27 B.n273 B.n272 585
R28 B.n271 B.n94 585
R29 B.n270 B.n269 585
R30 B.n268 B.n95 585
R31 B.n267 B.n266 585
R32 B.n265 B.n96 585
R33 B.n264 B.n263 585
R34 B.n262 B.n97 585
R35 B.n261 B.n260 585
R36 B.n259 B.n98 585
R37 B.n258 B.n257 585
R38 B.n256 B.n99 585
R39 B.n255 B.n254 585
R40 B.n253 B.n100 585
R41 B.n252 B.n251 585
R42 B.n250 B.n101 585
R43 B.n249 B.n248 585
R44 B.n247 B.n102 585
R45 B.n246 B.n245 585
R46 B.n241 B.n103 585
R47 B.n240 B.n239 585
R48 B.n238 B.n104 585
R49 B.n237 B.n236 585
R50 B.n235 B.n105 585
R51 B.n234 B.n233 585
R52 B.n232 B.n106 585
R53 B.n231 B.n230 585
R54 B.n229 B.n107 585
R55 B.n227 B.n226 585
R56 B.n225 B.n110 585
R57 B.n224 B.n223 585
R58 B.n222 B.n111 585
R59 B.n221 B.n220 585
R60 B.n219 B.n112 585
R61 B.n218 B.n217 585
R62 B.n216 B.n113 585
R63 B.n215 B.n214 585
R64 B.n213 B.n114 585
R65 B.n212 B.n211 585
R66 B.n210 B.n115 585
R67 B.n209 B.n208 585
R68 B.n207 B.n116 585
R69 B.n206 B.n205 585
R70 B.n204 B.n117 585
R71 B.n203 B.n202 585
R72 B.n201 B.n118 585
R73 B.n200 B.n199 585
R74 B.n198 B.n119 585
R75 B.n197 B.n196 585
R76 B.n195 B.n120 585
R77 B.n194 B.n193 585
R78 B.n192 B.n121 585
R79 B.n191 B.n190 585
R80 B.n189 B.n122 585
R81 B.n188 B.n187 585
R82 B.n186 B.n123 585
R83 B.n185 B.n184 585
R84 B.n183 B.n124 585
R85 B.n182 B.n181 585
R86 B.n180 B.n125 585
R87 B.n179 B.n178 585
R88 B.n177 B.n126 585
R89 B.n176 B.n175 585
R90 B.n174 B.n127 585
R91 B.n173 B.n172 585
R92 B.n171 B.n128 585
R93 B.n170 B.n169 585
R94 B.n168 B.n129 585
R95 B.n167 B.n166 585
R96 B.n309 B.n308 585
R97 B.n310 B.n81 585
R98 B.n312 B.n311 585
R99 B.n313 B.n80 585
R100 B.n315 B.n314 585
R101 B.n316 B.n79 585
R102 B.n318 B.n317 585
R103 B.n319 B.n78 585
R104 B.n321 B.n320 585
R105 B.n322 B.n77 585
R106 B.n324 B.n323 585
R107 B.n325 B.n76 585
R108 B.n327 B.n326 585
R109 B.n328 B.n75 585
R110 B.n330 B.n329 585
R111 B.n331 B.n74 585
R112 B.n333 B.n332 585
R113 B.n334 B.n73 585
R114 B.n336 B.n335 585
R115 B.n337 B.n72 585
R116 B.n339 B.n338 585
R117 B.n340 B.n71 585
R118 B.n342 B.n341 585
R119 B.n343 B.n70 585
R120 B.n345 B.n344 585
R121 B.n346 B.n69 585
R122 B.n348 B.n347 585
R123 B.n349 B.n68 585
R124 B.n351 B.n350 585
R125 B.n352 B.n67 585
R126 B.n354 B.n353 585
R127 B.n355 B.n66 585
R128 B.n357 B.n356 585
R129 B.n358 B.n65 585
R130 B.n360 B.n359 585
R131 B.n361 B.n64 585
R132 B.n363 B.n362 585
R133 B.n364 B.n63 585
R134 B.n366 B.n365 585
R135 B.n367 B.n62 585
R136 B.n507 B.n506 585
R137 B.n505 B.n12 585
R138 B.n504 B.n503 585
R139 B.n502 B.n13 585
R140 B.n501 B.n500 585
R141 B.n499 B.n14 585
R142 B.n498 B.n497 585
R143 B.n496 B.n15 585
R144 B.n495 B.n494 585
R145 B.n493 B.n16 585
R146 B.n492 B.n491 585
R147 B.n490 B.n17 585
R148 B.n489 B.n488 585
R149 B.n487 B.n18 585
R150 B.n486 B.n485 585
R151 B.n484 B.n19 585
R152 B.n483 B.n482 585
R153 B.n481 B.n20 585
R154 B.n480 B.n479 585
R155 B.n478 B.n21 585
R156 B.n477 B.n476 585
R157 B.n475 B.n22 585
R158 B.n474 B.n473 585
R159 B.n472 B.n23 585
R160 B.n471 B.n470 585
R161 B.n469 B.n24 585
R162 B.n468 B.n467 585
R163 B.n466 B.n25 585
R164 B.n465 B.n464 585
R165 B.n463 B.n26 585
R166 B.n462 B.n461 585
R167 B.n460 B.n27 585
R168 B.n459 B.n458 585
R169 B.n457 B.n28 585
R170 B.n456 B.n455 585
R171 B.n454 B.n29 585
R172 B.n453 B.n452 585
R173 B.n451 B.n30 585
R174 B.n450 B.n449 585
R175 B.n448 B.n31 585
R176 B.n447 B.n446 585
R177 B.n445 B.n444 585
R178 B.n443 B.n35 585
R179 B.n442 B.n441 585
R180 B.n440 B.n36 585
R181 B.n439 B.n438 585
R182 B.n437 B.n37 585
R183 B.n436 B.n435 585
R184 B.n434 B.n38 585
R185 B.n433 B.n432 585
R186 B.n431 B.n39 585
R187 B.n429 B.n428 585
R188 B.n427 B.n42 585
R189 B.n426 B.n425 585
R190 B.n424 B.n43 585
R191 B.n423 B.n422 585
R192 B.n421 B.n44 585
R193 B.n420 B.n419 585
R194 B.n418 B.n45 585
R195 B.n417 B.n416 585
R196 B.n415 B.n46 585
R197 B.n414 B.n413 585
R198 B.n412 B.n47 585
R199 B.n411 B.n410 585
R200 B.n409 B.n48 585
R201 B.n408 B.n407 585
R202 B.n406 B.n49 585
R203 B.n405 B.n404 585
R204 B.n403 B.n50 585
R205 B.n402 B.n401 585
R206 B.n400 B.n51 585
R207 B.n399 B.n398 585
R208 B.n397 B.n52 585
R209 B.n396 B.n395 585
R210 B.n394 B.n53 585
R211 B.n393 B.n392 585
R212 B.n391 B.n54 585
R213 B.n390 B.n389 585
R214 B.n388 B.n55 585
R215 B.n387 B.n386 585
R216 B.n385 B.n56 585
R217 B.n384 B.n383 585
R218 B.n382 B.n57 585
R219 B.n381 B.n380 585
R220 B.n379 B.n58 585
R221 B.n378 B.n377 585
R222 B.n376 B.n59 585
R223 B.n375 B.n374 585
R224 B.n373 B.n60 585
R225 B.n372 B.n371 585
R226 B.n370 B.n61 585
R227 B.n369 B.n368 585
R228 B.n508 B.n11 585
R229 B.n510 B.n509 585
R230 B.n511 B.n10 585
R231 B.n513 B.n512 585
R232 B.n514 B.n9 585
R233 B.n516 B.n515 585
R234 B.n517 B.n8 585
R235 B.n519 B.n518 585
R236 B.n520 B.n7 585
R237 B.n522 B.n521 585
R238 B.n523 B.n6 585
R239 B.n525 B.n524 585
R240 B.n526 B.n5 585
R241 B.n528 B.n527 585
R242 B.n529 B.n4 585
R243 B.n531 B.n530 585
R244 B.n532 B.n3 585
R245 B.n534 B.n533 585
R246 B.n535 B.n0 585
R247 B.n2 B.n1 585
R248 B.n140 B.n139 585
R249 B.n141 B.n138 585
R250 B.n143 B.n142 585
R251 B.n144 B.n137 585
R252 B.n146 B.n145 585
R253 B.n147 B.n136 585
R254 B.n149 B.n148 585
R255 B.n150 B.n135 585
R256 B.n152 B.n151 585
R257 B.n153 B.n134 585
R258 B.n155 B.n154 585
R259 B.n156 B.n133 585
R260 B.n158 B.n157 585
R261 B.n159 B.n132 585
R262 B.n161 B.n160 585
R263 B.n162 B.n131 585
R264 B.n164 B.n163 585
R265 B.n165 B.n130 585
R266 B.n166 B.n165 497.305
R267 B.n308 B.n307 497.305
R268 B.n368 B.n367 497.305
R269 B.n506 B.n11 497.305
R270 B.n537 B.n536 256.663
R271 B.n536 B.n535 235.042
R272 B.n536 B.n2 235.042
R273 B.n166 B.n129 163.367
R274 B.n170 B.n129 163.367
R275 B.n171 B.n170 163.367
R276 B.n172 B.n171 163.367
R277 B.n172 B.n127 163.367
R278 B.n176 B.n127 163.367
R279 B.n177 B.n176 163.367
R280 B.n178 B.n177 163.367
R281 B.n178 B.n125 163.367
R282 B.n182 B.n125 163.367
R283 B.n183 B.n182 163.367
R284 B.n184 B.n183 163.367
R285 B.n184 B.n123 163.367
R286 B.n188 B.n123 163.367
R287 B.n189 B.n188 163.367
R288 B.n190 B.n189 163.367
R289 B.n190 B.n121 163.367
R290 B.n194 B.n121 163.367
R291 B.n195 B.n194 163.367
R292 B.n196 B.n195 163.367
R293 B.n196 B.n119 163.367
R294 B.n200 B.n119 163.367
R295 B.n201 B.n200 163.367
R296 B.n202 B.n201 163.367
R297 B.n202 B.n117 163.367
R298 B.n206 B.n117 163.367
R299 B.n207 B.n206 163.367
R300 B.n208 B.n207 163.367
R301 B.n208 B.n115 163.367
R302 B.n212 B.n115 163.367
R303 B.n213 B.n212 163.367
R304 B.n214 B.n213 163.367
R305 B.n214 B.n113 163.367
R306 B.n218 B.n113 163.367
R307 B.n219 B.n218 163.367
R308 B.n220 B.n219 163.367
R309 B.n220 B.n111 163.367
R310 B.n224 B.n111 163.367
R311 B.n225 B.n224 163.367
R312 B.n226 B.n225 163.367
R313 B.n226 B.n107 163.367
R314 B.n231 B.n107 163.367
R315 B.n232 B.n231 163.367
R316 B.n233 B.n232 163.367
R317 B.n233 B.n105 163.367
R318 B.n237 B.n105 163.367
R319 B.n238 B.n237 163.367
R320 B.n239 B.n238 163.367
R321 B.n239 B.n103 163.367
R322 B.n246 B.n103 163.367
R323 B.n247 B.n246 163.367
R324 B.n248 B.n247 163.367
R325 B.n248 B.n101 163.367
R326 B.n252 B.n101 163.367
R327 B.n253 B.n252 163.367
R328 B.n254 B.n253 163.367
R329 B.n254 B.n99 163.367
R330 B.n258 B.n99 163.367
R331 B.n259 B.n258 163.367
R332 B.n260 B.n259 163.367
R333 B.n260 B.n97 163.367
R334 B.n264 B.n97 163.367
R335 B.n265 B.n264 163.367
R336 B.n266 B.n265 163.367
R337 B.n266 B.n95 163.367
R338 B.n270 B.n95 163.367
R339 B.n271 B.n270 163.367
R340 B.n272 B.n271 163.367
R341 B.n272 B.n93 163.367
R342 B.n276 B.n93 163.367
R343 B.n277 B.n276 163.367
R344 B.n278 B.n277 163.367
R345 B.n278 B.n91 163.367
R346 B.n282 B.n91 163.367
R347 B.n283 B.n282 163.367
R348 B.n284 B.n283 163.367
R349 B.n284 B.n89 163.367
R350 B.n288 B.n89 163.367
R351 B.n289 B.n288 163.367
R352 B.n290 B.n289 163.367
R353 B.n290 B.n87 163.367
R354 B.n294 B.n87 163.367
R355 B.n295 B.n294 163.367
R356 B.n296 B.n295 163.367
R357 B.n296 B.n85 163.367
R358 B.n300 B.n85 163.367
R359 B.n301 B.n300 163.367
R360 B.n302 B.n301 163.367
R361 B.n302 B.n83 163.367
R362 B.n306 B.n83 163.367
R363 B.n307 B.n306 163.367
R364 B.n367 B.n366 163.367
R365 B.n366 B.n63 163.367
R366 B.n362 B.n63 163.367
R367 B.n362 B.n361 163.367
R368 B.n361 B.n360 163.367
R369 B.n360 B.n65 163.367
R370 B.n356 B.n65 163.367
R371 B.n356 B.n355 163.367
R372 B.n355 B.n354 163.367
R373 B.n354 B.n67 163.367
R374 B.n350 B.n67 163.367
R375 B.n350 B.n349 163.367
R376 B.n349 B.n348 163.367
R377 B.n348 B.n69 163.367
R378 B.n344 B.n69 163.367
R379 B.n344 B.n343 163.367
R380 B.n343 B.n342 163.367
R381 B.n342 B.n71 163.367
R382 B.n338 B.n71 163.367
R383 B.n338 B.n337 163.367
R384 B.n337 B.n336 163.367
R385 B.n336 B.n73 163.367
R386 B.n332 B.n73 163.367
R387 B.n332 B.n331 163.367
R388 B.n331 B.n330 163.367
R389 B.n330 B.n75 163.367
R390 B.n326 B.n75 163.367
R391 B.n326 B.n325 163.367
R392 B.n325 B.n324 163.367
R393 B.n324 B.n77 163.367
R394 B.n320 B.n77 163.367
R395 B.n320 B.n319 163.367
R396 B.n319 B.n318 163.367
R397 B.n318 B.n79 163.367
R398 B.n314 B.n79 163.367
R399 B.n314 B.n313 163.367
R400 B.n313 B.n312 163.367
R401 B.n312 B.n81 163.367
R402 B.n308 B.n81 163.367
R403 B.n506 B.n505 163.367
R404 B.n505 B.n504 163.367
R405 B.n504 B.n13 163.367
R406 B.n500 B.n13 163.367
R407 B.n500 B.n499 163.367
R408 B.n499 B.n498 163.367
R409 B.n498 B.n15 163.367
R410 B.n494 B.n15 163.367
R411 B.n494 B.n493 163.367
R412 B.n493 B.n492 163.367
R413 B.n492 B.n17 163.367
R414 B.n488 B.n17 163.367
R415 B.n488 B.n487 163.367
R416 B.n487 B.n486 163.367
R417 B.n486 B.n19 163.367
R418 B.n482 B.n19 163.367
R419 B.n482 B.n481 163.367
R420 B.n481 B.n480 163.367
R421 B.n480 B.n21 163.367
R422 B.n476 B.n21 163.367
R423 B.n476 B.n475 163.367
R424 B.n475 B.n474 163.367
R425 B.n474 B.n23 163.367
R426 B.n470 B.n23 163.367
R427 B.n470 B.n469 163.367
R428 B.n469 B.n468 163.367
R429 B.n468 B.n25 163.367
R430 B.n464 B.n25 163.367
R431 B.n464 B.n463 163.367
R432 B.n463 B.n462 163.367
R433 B.n462 B.n27 163.367
R434 B.n458 B.n27 163.367
R435 B.n458 B.n457 163.367
R436 B.n457 B.n456 163.367
R437 B.n456 B.n29 163.367
R438 B.n452 B.n29 163.367
R439 B.n452 B.n451 163.367
R440 B.n451 B.n450 163.367
R441 B.n450 B.n31 163.367
R442 B.n446 B.n31 163.367
R443 B.n446 B.n445 163.367
R444 B.n445 B.n35 163.367
R445 B.n441 B.n35 163.367
R446 B.n441 B.n440 163.367
R447 B.n440 B.n439 163.367
R448 B.n439 B.n37 163.367
R449 B.n435 B.n37 163.367
R450 B.n435 B.n434 163.367
R451 B.n434 B.n433 163.367
R452 B.n433 B.n39 163.367
R453 B.n428 B.n39 163.367
R454 B.n428 B.n427 163.367
R455 B.n427 B.n426 163.367
R456 B.n426 B.n43 163.367
R457 B.n422 B.n43 163.367
R458 B.n422 B.n421 163.367
R459 B.n421 B.n420 163.367
R460 B.n420 B.n45 163.367
R461 B.n416 B.n45 163.367
R462 B.n416 B.n415 163.367
R463 B.n415 B.n414 163.367
R464 B.n414 B.n47 163.367
R465 B.n410 B.n47 163.367
R466 B.n410 B.n409 163.367
R467 B.n409 B.n408 163.367
R468 B.n408 B.n49 163.367
R469 B.n404 B.n49 163.367
R470 B.n404 B.n403 163.367
R471 B.n403 B.n402 163.367
R472 B.n402 B.n51 163.367
R473 B.n398 B.n51 163.367
R474 B.n398 B.n397 163.367
R475 B.n397 B.n396 163.367
R476 B.n396 B.n53 163.367
R477 B.n392 B.n53 163.367
R478 B.n392 B.n391 163.367
R479 B.n391 B.n390 163.367
R480 B.n390 B.n55 163.367
R481 B.n386 B.n55 163.367
R482 B.n386 B.n385 163.367
R483 B.n385 B.n384 163.367
R484 B.n384 B.n57 163.367
R485 B.n380 B.n57 163.367
R486 B.n380 B.n379 163.367
R487 B.n379 B.n378 163.367
R488 B.n378 B.n59 163.367
R489 B.n374 B.n59 163.367
R490 B.n374 B.n373 163.367
R491 B.n373 B.n372 163.367
R492 B.n372 B.n61 163.367
R493 B.n368 B.n61 163.367
R494 B.n510 B.n11 163.367
R495 B.n511 B.n510 163.367
R496 B.n512 B.n511 163.367
R497 B.n512 B.n9 163.367
R498 B.n516 B.n9 163.367
R499 B.n517 B.n516 163.367
R500 B.n518 B.n517 163.367
R501 B.n518 B.n7 163.367
R502 B.n522 B.n7 163.367
R503 B.n523 B.n522 163.367
R504 B.n524 B.n523 163.367
R505 B.n524 B.n5 163.367
R506 B.n528 B.n5 163.367
R507 B.n529 B.n528 163.367
R508 B.n530 B.n529 163.367
R509 B.n530 B.n3 163.367
R510 B.n534 B.n3 163.367
R511 B.n535 B.n534 163.367
R512 B.n140 B.n2 163.367
R513 B.n141 B.n140 163.367
R514 B.n142 B.n141 163.367
R515 B.n142 B.n137 163.367
R516 B.n146 B.n137 163.367
R517 B.n147 B.n146 163.367
R518 B.n148 B.n147 163.367
R519 B.n148 B.n135 163.367
R520 B.n152 B.n135 163.367
R521 B.n153 B.n152 163.367
R522 B.n154 B.n153 163.367
R523 B.n154 B.n133 163.367
R524 B.n158 B.n133 163.367
R525 B.n159 B.n158 163.367
R526 B.n160 B.n159 163.367
R527 B.n160 B.n131 163.367
R528 B.n164 B.n131 163.367
R529 B.n165 B.n164 163.367
R530 B.n242 B.t4 132.149
R531 B.n40 B.t2 132.149
R532 B.n108 B.t7 132.136
R533 B.n32 B.t11 132.136
R534 B.n243 B.t5 113.531
R535 B.n41 B.t1 113.531
R536 B.n109 B.t8 113.517
R537 B.n33 B.t10 113.517
R538 B.n228 B.n109 59.5399
R539 B.n244 B.n243 59.5399
R540 B.n430 B.n41 59.5399
R541 B.n34 B.n33 59.5399
R542 B.n508 B.n507 32.3127
R543 B.n369 B.n62 32.3127
R544 B.n309 B.n82 32.3127
R545 B.n167 B.n130 32.3127
R546 B.n109 B.n108 18.6187
R547 B.n243 B.n242 18.6187
R548 B.n41 B.n40 18.6187
R549 B.n33 B.n32 18.6187
R550 B B.n537 18.0485
R551 B.n509 B.n508 10.6151
R552 B.n509 B.n10 10.6151
R553 B.n513 B.n10 10.6151
R554 B.n514 B.n513 10.6151
R555 B.n515 B.n514 10.6151
R556 B.n515 B.n8 10.6151
R557 B.n519 B.n8 10.6151
R558 B.n520 B.n519 10.6151
R559 B.n521 B.n520 10.6151
R560 B.n521 B.n6 10.6151
R561 B.n525 B.n6 10.6151
R562 B.n526 B.n525 10.6151
R563 B.n527 B.n526 10.6151
R564 B.n527 B.n4 10.6151
R565 B.n531 B.n4 10.6151
R566 B.n532 B.n531 10.6151
R567 B.n533 B.n532 10.6151
R568 B.n533 B.n0 10.6151
R569 B.n507 B.n12 10.6151
R570 B.n503 B.n12 10.6151
R571 B.n503 B.n502 10.6151
R572 B.n502 B.n501 10.6151
R573 B.n501 B.n14 10.6151
R574 B.n497 B.n14 10.6151
R575 B.n497 B.n496 10.6151
R576 B.n496 B.n495 10.6151
R577 B.n495 B.n16 10.6151
R578 B.n491 B.n16 10.6151
R579 B.n491 B.n490 10.6151
R580 B.n490 B.n489 10.6151
R581 B.n489 B.n18 10.6151
R582 B.n485 B.n18 10.6151
R583 B.n485 B.n484 10.6151
R584 B.n484 B.n483 10.6151
R585 B.n483 B.n20 10.6151
R586 B.n479 B.n20 10.6151
R587 B.n479 B.n478 10.6151
R588 B.n478 B.n477 10.6151
R589 B.n477 B.n22 10.6151
R590 B.n473 B.n22 10.6151
R591 B.n473 B.n472 10.6151
R592 B.n472 B.n471 10.6151
R593 B.n471 B.n24 10.6151
R594 B.n467 B.n24 10.6151
R595 B.n467 B.n466 10.6151
R596 B.n466 B.n465 10.6151
R597 B.n465 B.n26 10.6151
R598 B.n461 B.n26 10.6151
R599 B.n461 B.n460 10.6151
R600 B.n460 B.n459 10.6151
R601 B.n459 B.n28 10.6151
R602 B.n455 B.n28 10.6151
R603 B.n455 B.n454 10.6151
R604 B.n454 B.n453 10.6151
R605 B.n453 B.n30 10.6151
R606 B.n449 B.n30 10.6151
R607 B.n449 B.n448 10.6151
R608 B.n448 B.n447 10.6151
R609 B.n444 B.n443 10.6151
R610 B.n443 B.n442 10.6151
R611 B.n442 B.n36 10.6151
R612 B.n438 B.n36 10.6151
R613 B.n438 B.n437 10.6151
R614 B.n437 B.n436 10.6151
R615 B.n436 B.n38 10.6151
R616 B.n432 B.n38 10.6151
R617 B.n432 B.n431 10.6151
R618 B.n429 B.n42 10.6151
R619 B.n425 B.n42 10.6151
R620 B.n425 B.n424 10.6151
R621 B.n424 B.n423 10.6151
R622 B.n423 B.n44 10.6151
R623 B.n419 B.n44 10.6151
R624 B.n419 B.n418 10.6151
R625 B.n418 B.n417 10.6151
R626 B.n417 B.n46 10.6151
R627 B.n413 B.n46 10.6151
R628 B.n413 B.n412 10.6151
R629 B.n412 B.n411 10.6151
R630 B.n411 B.n48 10.6151
R631 B.n407 B.n48 10.6151
R632 B.n407 B.n406 10.6151
R633 B.n406 B.n405 10.6151
R634 B.n405 B.n50 10.6151
R635 B.n401 B.n50 10.6151
R636 B.n401 B.n400 10.6151
R637 B.n400 B.n399 10.6151
R638 B.n399 B.n52 10.6151
R639 B.n395 B.n52 10.6151
R640 B.n395 B.n394 10.6151
R641 B.n394 B.n393 10.6151
R642 B.n393 B.n54 10.6151
R643 B.n389 B.n54 10.6151
R644 B.n389 B.n388 10.6151
R645 B.n388 B.n387 10.6151
R646 B.n387 B.n56 10.6151
R647 B.n383 B.n56 10.6151
R648 B.n383 B.n382 10.6151
R649 B.n382 B.n381 10.6151
R650 B.n381 B.n58 10.6151
R651 B.n377 B.n58 10.6151
R652 B.n377 B.n376 10.6151
R653 B.n376 B.n375 10.6151
R654 B.n375 B.n60 10.6151
R655 B.n371 B.n60 10.6151
R656 B.n371 B.n370 10.6151
R657 B.n370 B.n369 10.6151
R658 B.n365 B.n62 10.6151
R659 B.n365 B.n364 10.6151
R660 B.n364 B.n363 10.6151
R661 B.n363 B.n64 10.6151
R662 B.n359 B.n64 10.6151
R663 B.n359 B.n358 10.6151
R664 B.n358 B.n357 10.6151
R665 B.n357 B.n66 10.6151
R666 B.n353 B.n66 10.6151
R667 B.n353 B.n352 10.6151
R668 B.n352 B.n351 10.6151
R669 B.n351 B.n68 10.6151
R670 B.n347 B.n68 10.6151
R671 B.n347 B.n346 10.6151
R672 B.n346 B.n345 10.6151
R673 B.n345 B.n70 10.6151
R674 B.n341 B.n70 10.6151
R675 B.n341 B.n340 10.6151
R676 B.n340 B.n339 10.6151
R677 B.n339 B.n72 10.6151
R678 B.n335 B.n72 10.6151
R679 B.n335 B.n334 10.6151
R680 B.n334 B.n333 10.6151
R681 B.n333 B.n74 10.6151
R682 B.n329 B.n74 10.6151
R683 B.n329 B.n328 10.6151
R684 B.n328 B.n327 10.6151
R685 B.n327 B.n76 10.6151
R686 B.n323 B.n76 10.6151
R687 B.n323 B.n322 10.6151
R688 B.n322 B.n321 10.6151
R689 B.n321 B.n78 10.6151
R690 B.n317 B.n78 10.6151
R691 B.n317 B.n316 10.6151
R692 B.n316 B.n315 10.6151
R693 B.n315 B.n80 10.6151
R694 B.n311 B.n80 10.6151
R695 B.n311 B.n310 10.6151
R696 B.n310 B.n309 10.6151
R697 B.n139 B.n1 10.6151
R698 B.n139 B.n138 10.6151
R699 B.n143 B.n138 10.6151
R700 B.n144 B.n143 10.6151
R701 B.n145 B.n144 10.6151
R702 B.n145 B.n136 10.6151
R703 B.n149 B.n136 10.6151
R704 B.n150 B.n149 10.6151
R705 B.n151 B.n150 10.6151
R706 B.n151 B.n134 10.6151
R707 B.n155 B.n134 10.6151
R708 B.n156 B.n155 10.6151
R709 B.n157 B.n156 10.6151
R710 B.n157 B.n132 10.6151
R711 B.n161 B.n132 10.6151
R712 B.n162 B.n161 10.6151
R713 B.n163 B.n162 10.6151
R714 B.n163 B.n130 10.6151
R715 B.n168 B.n167 10.6151
R716 B.n169 B.n168 10.6151
R717 B.n169 B.n128 10.6151
R718 B.n173 B.n128 10.6151
R719 B.n174 B.n173 10.6151
R720 B.n175 B.n174 10.6151
R721 B.n175 B.n126 10.6151
R722 B.n179 B.n126 10.6151
R723 B.n180 B.n179 10.6151
R724 B.n181 B.n180 10.6151
R725 B.n181 B.n124 10.6151
R726 B.n185 B.n124 10.6151
R727 B.n186 B.n185 10.6151
R728 B.n187 B.n186 10.6151
R729 B.n187 B.n122 10.6151
R730 B.n191 B.n122 10.6151
R731 B.n192 B.n191 10.6151
R732 B.n193 B.n192 10.6151
R733 B.n193 B.n120 10.6151
R734 B.n197 B.n120 10.6151
R735 B.n198 B.n197 10.6151
R736 B.n199 B.n198 10.6151
R737 B.n199 B.n118 10.6151
R738 B.n203 B.n118 10.6151
R739 B.n204 B.n203 10.6151
R740 B.n205 B.n204 10.6151
R741 B.n205 B.n116 10.6151
R742 B.n209 B.n116 10.6151
R743 B.n210 B.n209 10.6151
R744 B.n211 B.n210 10.6151
R745 B.n211 B.n114 10.6151
R746 B.n215 B.n114 10.6151
R747 B.n216 B.n215 10.6151
R748 B.n217 B.n216 10.6151
R749 B.n217 B.n112 10.6151
R750 B.n221 B.n112 10.6151
R751 B.n222 B.n221 10.6151
R752 B.n223 B.n222 10.6151
R753 B.n223 B.n110 10.6151
R754 B.n227 B.n110 10.6151
R755 B.n230 B.n229 10.6151
R756 B.n230 B.n106 10.6151
R757 B.n234 B.n106 10.6151
R758 B.n235 B.n234 10.6151
R759 B.n236 B.n235 10.6151
R760 B.n236 B.n104 10.6151
R761 B.n240 B.n104 10.6151
R762 B.n241 B.n240 10.6151
R763 B.n245 B.n241 10.6151
R764 B.n249 B.n102 10.6151
R765 B.n250 B.n249 10.6151
R766 B.n251 B.n250 10.6151
R767 B.n251 B.n100 10.6151
R768 B.n255 B.n100 10.6151
R769 B.n256 B.n255 10.6151
R770 B.n257 B.n256 10.6151
R771 B.n257 B.n98 10.6151
R772 B.n261 B.n98 10.6151
R773 B.n262 B.n261 10.6151
R774 B.n263 B.n262 10.6151
R775 B.n263 B.n96 10.6151
R776 B.n267 B.n96 10.6151
R777 B.n268 B.n267 10.6151
R778 B.n269 B.n268 10.6151
R779 B.n269 B.n94 10.6151
R780 B.n273 B.n94 10.6151
R781 B.n274 B.n273 10.6151
R782 B.n275 B.n274 10.6151
R783 B.n275 B.n92 10.6151
R784 B.n279 B.n92 10.6151
R785 B.n280 B.n279 10.6151
R786 B.n281 B.n280 10.6151
R787 B.n281 B.n90 10.6151
R788 B.n285 B.n90 10.6151
R789 B.n286 B.n285 10.6151
R790 B.n287 B.n286 10.6151
R791 B.n287 B.n88 10.6151
R792 B.n291 B.n88 10.6151
R793 B.n292 B.n291 10.6151
R794 B.n293 B.n292 10.6151
R795 B.n293 B.n86 10.6151
R796 B.n297 B.n86 10.6151
R797 B.n298 B.n297 10.6151
R798 B.n299 B.n298 10.6151
R799 B.n299 B.n84 10.6151
R800 B.n303 B.n84 10.6151
R801 B.n304 B.n303 10.6151
R802 B.n305 B.n304 10.6151
R803 B.n305 B.n82 10.6151
R804 B.n447 B.n34 9.36635
R805 B.n430 B.n429 9.36635
R806 B.n228 B.n227 9.36635
R807 B.n244 B.n102 9.36635
R808 B.n537 B.n0 8.11757
R809 B.n537 B.n1 8.11757
R810 B.n444 B.n34 1.24928
R811 B.n431 B.n430 1.24928
R812 B.n229 B.n228 1.24928
R813 B.n245 B.n244 1.24928
R814 VP.n1 VP.t3 544.398
R815 VP.n6 VP.t1 517.577
R816 VP.n7 VP.t0 517.577
R817 VP.n8 VP.t5 517.577
R818 VP.n3 VP.t2 517.577
R819 VP.n2 VP.t4 517.577
R820 VP.n9 VP.n8 161.3
R821 VP.n4 VP.n3 161.3
R822 VP.n6 VP.n5 161.3
R823 VP.n7 VP.n0 80.6037
R824 VP.n7 VP.n6 48.2005
R825 VP.n8 VP.n7 48.2005
R826 VP.n3 VP.n2 48.2005
R827 VP.n4 VP.n1 45.1367
R828 VP.n5 VP.n4 40.9626
R829 VP.n2 VP.n1 13.3799
R830 VP.n5 VP.n0 0.285035
R831 VP.n9 VP.n0 0.285035
R832 VP VP.n9 0.0516364
R833 VDD1 VDD1.t5 80.2288
R834 VDD1.n1 VDD1.t2 80.115
R835 VDD1.n1 VDD1.n0 76.9674
R836 VDD1.n3 VDD1.n2 76.816
R837 VDD1.n3 VDD1.n1 37.6518
R838 VDD1.n2 VDD1.t3 2.73431
R839 VDD1.n2 VDD1.t0 2.73431
R840 VDD1.n0 VDD1.t4 2.73431
R841 VDD1.n0 VDD1.t1 2.73431
R842 VDD1 VDD1.n3 0.149207
R843 VTAIL.n7 VTAIL.t4 62.8712
R844 VTAIL.n11 VTAIL.t3 62.8709
R845 VTAIL.n2 VTAIL.t6 62.8709
R846 VTAIL.n10 VTAIL.t9 62.8709
R847 VTAIL.n9 VTAIL.n8 60.1374
R848 VTAIL.n6 VTAIL.n5 60.1374
R849 VTAIL.n1 VTAIL.n0 60.1371
R850 VTAIL.n4 VTAIL.n3 60.1371
R851 VTAIL.n6 VTAIL.n4 24.2721
R852 VTAIL.n11 VTAIL.n10 23.4445
R853 VTAIL.n0 VTAIL.t0 2.73431
R854 VTAIL.n0 VTAIL.t1 2.73431
R855 VTAIL.n3 VTAIL.t10 2.73431
R856 VTAIL.n3 VTAIL.t11 2.73431
R857 VTAIL.n8 VTAIL.t8 2.73431
R858 VTAIL.n8 VTAIL.t7 2.73431
R859 VTAIL.n5 VTAIL.t2 2.73431
R860 VTAIL.n5 VTAIL.t5 2.73431
R861 VTAIL.n9 VTAIL.n7 0.884121
R862 VTAIL.n2 VTAIL.n1 0.884121
R863 VTAIL.n7 VTAIL.n6 0.828086
R864 VTAIL.n10 VTAIL.n9 0.828086
R865 VTAIL.n4 VTAIL.n2 0.828086
R866 VTAIL VTAIL.n11 0.563
R867 VTAIL VTAIL.n1 0.265586
R868 VN.n0 VN.t4 544.398
R869 VN.n4 VN.t1 544.398
R870 VN.n1 VN.t5 517.577
R871 VN.n2 VN.t0 517.577
R872 VN.n5 VN.t2 517.577
R873 VN.n6 VN.t3 517.577
R874 VN.n3 VN.n2 161.3
R875 VN.n7 VN.n6 161.3
R876 VN.n2 VN.n1 48.2005
R877 VN.n6 VN.n5 48.2005
R878 VN.n7 VN.n4 45.1367
R879 VN.n3 VN.n0 45.1367
R880 VN VN.n7 41.3433
R881 VN.n5 VN.n4 13.3799
R882 VN.n1 VN.n0 13.3799
R883 VN VN.n3 0.0516364
R884 VDD2.n1 VDD2.t1 80.115
R885 VDD2.n2 VDD2.t2 79.55
R886 VDD2.n1 VDD2.n0 76.9674
R887 VDD2 VDD2.n3 76.9647
R888 VDD2.n2 VDD2.n1 36.6549
R889 VDD2.n3 VDD2.t3 2.73431
R890 VDD2.n3 VDD2.t4 2.73431
R891 VDD2.n0 VDD2.t0 2.73431
R892 VDD2.n0 VDD2.t5 2.73431
R893 VDD2 VDD2.n2 0.679379
C0 B VDD2 1.55727f
C1 w_n1738_n3346# VN 2.80256f
C2 B VDD1 1.52994f
C3 VN VDD2 4.07633f
C4 B VTAIL 2.64151f
C5 VN VDD1 0.148102f
C6 VN VTAIL 3.74469f
C7 w_n1738_n3346# VP 3.02177f
C8 VP VDD2 0.291766f
C9 VP VDD1 4.21541f
C10 VTAIL VP 3.75931f
C11 B VN 0.747875f
C12 w_n1738_n3346# VDD2 1.80658f
C13 w_n1738_n3346# VDD1 1.7847f
C14 w_n1738_n3346# VTAIL 2.93f
C15 VDD1 VDD2 0.686074f
C16 VTAIL VDD2 10.2921f
C17 B VP 1.10395f
C18 VTAIL VDD1 10.2588f
C19 VN VP 4.98877f
C20 B w_n1738_n3346# 6.92615f
C21 VDD2 VSUBS 1.301013f
C22 VDD1 VSUBS 1.591829f
C23 VTAIL VSUBS 0.727136f
C24 VN VSUBS 4.42087f
C25 VP VSUBS 1.420005f
C26 B VSUBS 2.674959f
C27 w_n1738_n3346# VSUBS 71.5986f
C28 VDD2.t1 VSUBS 2.29093f
C29 VDD2.t0 VSUBS 0.223677f
C30 VDD2.t5 VSUBS 0.223677f
C31 VDD2.n0 VSUBS 1.75138f
C32 VDD2.n1 VSUBS 2.44335f
C33 VDD2.t2 VSUBS 2.28694f
C34 VDD2.n2 VSUBS 2.39584f
C35 VDD2.t3 VSUBS 0.223677f
C36 VDD2.t4 VSUBS 0.223677f
C37 VDD2.n3 VSUBS 1.75135f
C38 VN.t4 VSUBS 1.26729f
C39 VN.n0 VSUBS 0.475532f
C40 VN.t5 VSUBS 1.2427f
C41 VN.n1 VSUBS 0.512042f
C42 VN.t0 VSUBS 1.2427f
C43 VN.n2 VSUBS 0.498845f
C44 VN.n3 VSUBS 0.237977f
C45 VN.t1 VSUBS 1.26729f
C46 VN.n4 VSUBS 0.475532f
C47 VN.t2 VSUBS 1.2427f
C48 VN.n5 VSUBS 0.512042f
C49 VN.t3 VSUBS 1.2427f
C50 VN.n6 VSUBS 0.498845f
C51 VN.n7 VSUBS 2.53274f
C52 VTAIL.t0 VSUBS 0.277529f
C53 VTAIL.t1 VSUBS 0.277529f
C54 VTAIL.n0 VSUBS 2.02239f
C55 VTAIL.n1 VSUBS 0.762675f
C56 VTAIL.t6 VSUBS 2.67051f
C57 VTAIL.n2 VSUBS 0.924996f
C58 VTAIL.t10 VSUBS 0.277529f
C59 VTAIL.t11 VSUBS 0.277529f
C60 VTAIL.n3 VSUBS 2.02239f
C61 VTAIL.n4 VSUBS 2.26643f
C62 VTAIL.t2 VSUBS 0.277529f
C63 VTAIL.t5 VSUBS 0.277529f
C64 VTAIL.n5 VSUBS 2.0224f
C65 VTAIL.n6 VSUBS 2.26642f
C66 VTAIL.t4 VSUBS 2.67051f
C67 VTAIL.n7 VSUBS 0.924988f
C68 VTAIL.t8 VSUBS 0.277529f
C69 VTAIL.t7 VSUBS 0.277529f
C70 VTAIL.n8 VSUBS 2.0224f
C71 VTAIL.n9 VSUBS 0.816203f
C72 VTAIL.t9 VSUBS 2.67051f
C73 VTAIL.n10 VSUBS 2.29645f
C74 VTAIL.t3 VSUBS 2.67051f
C75 VTAIL.n11 VSUBS 2.27122f
C76 VDD1.t5 VSUBS 2.29371f
C77 VDD1.t2 VSUBS 2.29284f
C78 VDD1.t4 VSUBS 0.223863f
C79 VDD1.t1 VSUBS 0.223863f
C80 VDD1.n0 VSUBS 1.75284f
C81 VDD1.n1 VSUBS 2.51731f
C82 VDD1.t3 VSUBS 0.223863f
C83 VDD1.t0 VSUBS 0.223863f
C84 VDD1.n2 VSUBS 1.7518f
C85 VDD1.n3 VSUBS 2.36326f
C86 VP.n0 VSUBS 0.079821f
C87 VP.t3 VSUBS 1.30663f
C88 VP.n1 VSUBS 0.490294f
C89 VP.t2 VSUBS 1.28128f
C90 VP.t4 VSUBS 1.28128f
C91 VP.n2 VSUBS 0.527937f
C92 VP.n3 VSUBS 0.514331f
C93 VP.n4 VSUBS 2.57195f
C94 VP.n5 VSUBS 2.44571f
C95 VP.t1 VSUBS 1.28128f
C96 VP.n6 VSUBS 0.514331f
C97 VP.t0 VSUBS 1.28128f
C98 VP.n7 VSUBS 0.527937f
C99 VP.t5 VSUBS 1.28128f
C100 VP.n8 VSUBS 0.514331f
C101 VP.n9 VSUBS 0.066515f
C102 B.n0 VSUBS 0.006497f
C103 B.n1 VSUBS 0.006497f
C104 B.n2 VSUBS 0.009608f
C105 B.n3 VSUBS 0.007363f
C106 B.n4 VSUBS 0.007363f
C107 B.n5 VSUBS 0.007363f
C108 B.n6 VSUBS 0.007363f
C109 B.n7 VSUBS 0.007363f
C110 B.n8 VSUBS 0.007363f
C111 B.n9 VSUBS 0.007363f
C112 B.n10 VSUBS 0.007363f
C113 B.n11 VSUBS 0.016818f
C114 B.n12 VSUBS 0.007363f
C115 B.n13 VSUBS 0.007363f
C116 B.n14 VSUBS 0.007363f
C117 B.n15 VSUBS 0.007363f
C118 B.n16 VSUBS 0.007363f
C119 B.n17 VSUBS 0.007363f
C120 B.n18 VSUBS 0.007363f
C121 B.n19 VSUBS 0.007363f
C122 B.n20 VSUBS 0.007363f
C123 B.n21 VSUBS 0.007363f
C124 B.n22 VSUBS 0.007363f
C125 B.n23 VSUBS 0.007363f
C126 B.n24 VSUBS 0.007363f
C127 B.n25 VSUBS 0.007363f
C128 B.n26 VSUBS 0.007363f
C129 B.n27 VSUBS 0.007363f
C130 B.n28 VSUBS 0.007363f
C131 B.n29 VSUBS 0.007363f
C132 B.n30 VSUBS 0.007363f
C133 B.n31 VSUBS 0.007363f
C134 B.t10 VSUBS 0.407157f
C135 B.t11 VSUBS 0.415108f
C136 B.t9 VSUBS 0.322869f
C137 B.n32 VSUBS 0.135374f
C138 B.n33 VSUBS 0.06693f
C139 B.n34 VSUBS 0.017059f
C140 B.n35 VSUBS 0.007363f
C141 B.n36 VSUBS 0.007363f
C142 B.n37 VSUBS 0.007363f
C143 B.n38 VSUBS 0.007363f
C144 B.n39 VSUBS 0.007363f
C145 B.t1 VSUBS 0.40715f
C146 B.t2 VSUBS 0.415101f
C147 B.t0 VSUBS 0.322869f
C148 B.n40 VSUBS 0.135381f
C149 B.n41 VSUBS 0.066937f
C150 B.n42 VSUBS 0.007363f
C151 B.n43 VSUBS 0.007363f
C152 B.n44 VSUBS 0.007363f
C153 B.n45 VSUBS 0.007363f
C154 B.n46 VSUBS 0.007363f
C155 B.n47 VSUBS 0.007363f
C156 B.n48 VSUBS 0.007363f
C157 B.n49 VSUBS 0.007363f
C158 B.n50 VSUBS 0.007363f
C159 B.n51 VSUBS 0.007363f
C160 B.n52 VSUBS 0.007363f
C161 B.n53 VSUBS 0.007363f
C162 B.n54 VSUBS 0.007363f
C163 B.n55 VSUBS 0.007363f
C164 B.n56 VSUBS 0.007363f
C165 B.n57 VSUBS 0.007363f
C166 B.n58 VSUBS 0.007363f
C167 B.n59 VSUBS 0.007363f
C168 B.n60 VSUBS 0.007363f
C169 B.n61 VSUBS 0.007363f
C170 B.n62 VSUBS 0.016818f
C171 B.n63 VSUBS 0.007363f
C172 B.n64 VSUBS 0.007363f
C173 B.n65 VSUBS 0.007363f
C174 B.n66 VSUBS 0.007363f
C175 B.n67 VSUBS 0.007363f
C176 B.n68 VSUBS 0.007363f
C177 B.n69 VSUBS 0.007363f
C178 B.n70 VSUBS 0.007363f
C179 B.n71 VSUBS 0.007363f
C180 B.n72 VSUBS 0.007363f
C181 B.n73 VSUBS 0.007363f
C182 B.n74 VSUBS 0.007363f
C183 B.n75 VSUBS 0.007363f
C184 B.n76 VSUBS 0.007363f
C185 B.n77 VSUBS 0.007363f
C186 B.n78 VSUBS 0.007363f
C187 B.n79 VSUBS 0.007363f
C188 B.n80 VSUBS 0.007363f
C189 B.n81 VSUBS 0.007363f
C190 B.n82 VSUBS 0.016518f
C191 B.n83 VSUBS 0.007363f
C192 B.n84 VSUBS 0.007363f
C193 B.n85 VSUBS 0.007363f
C194 B.n86 VSUBS 0.007363f
C195 B.n87 VSUBS 0.007363f
C196 B.n88 VSUBS 0.007363f
C197 B.n89 VSUBS 0.007363f
C198 B.n90 VSUBS 0.007363f
C199 B.n91 VSUBS 0.007363f
C200 B.n92 VSUBS 0.007363f
C201 B.n93 VSUBS 0.007363f
C202 B.n94 VSUBS 0.007363f
C203 B.n95 VSUBS 0.007363f
C204 B.n96 VSUBS 0.007363f
C205 B.n97 VSUBS 0.007363f
C206 B.n98 VSUBS 0.007363f
C207 B.n99 VSUBS 0.007363f
C208 B.n100 VSUBS 0.007363f
C209 B.n101 VSUBS 0.007363f
C210 B.n102 VSUBS 0.00693f
C211 B.n103 VSUBS 0.007363f
C212 B.n104 VSUBS 0.007363f
C213 B.n105 VSUBS 0.007363f
C214 B.n106 VSUBS 0.007363f
C215 B.n107 VSUBS 0.007363f
C216 B.t8 VSUBS 0.407157f
C217 B.t7 VSUBS 0.415108f
C218 B.t6 VSUBS 0.322869f
C219 B.n108 VSUBS 0.135374f
C220 B.n109 VSUBS 0.06693f
C221 B.n110 VSUBS 0.007363f
C222 B.n111 VSUBS 0.007363f
C223 B.n112 VSUBS 0.007363f
C224 B.n113 VSUBS 0.007363f
C225 B.n114 VSUBS 0.007363f
C226 B.n115 VSUBS 0.007363f
C227 B.n116 VSUBS 0.007363f
C228 B.n117 VSUBS 0.007363f
C229 B.n118 VSUBS 0.007363f
C230 B.n119 VSUBS 0.007363f
C231 B.n120 VSUBS 0.007363f
C232 B.n121 VSUBS 0.007363f
C233 B.n122 VSUBS 0.007363f
C234 B.n123 VSUBS 0.007363f
C235 B.n124 VSUBS 0.007363f
C236 B.n125 VSUBS 0.007363f
C237 B.n126 VSUBS 0.007363f
C238 B.n127 VSUBS 0.007363f
C239 B.n128 VSUBS 0.007363f
C240 B.n129 VSUBS 0.007363f
C241 B.n130 VSUBS 0.016818f
C242 B.n131 VSUBS 0.007363f
C243 B.n132 VSUBS 0.007363f
C244 B.n133 VSUBS 0.007363f
C245 B.n134 VSUBS 0.007363f
C246 B.n135 VSUBS 0.007363f
C247 B.n136 VSUBS 0.007363f
C248 B.n137 VSUBS 0.007363f
C249 B.n138 VSUBS 0.007363f
C250 B.n139 VSUBS 0.007363f
C251 B.n140 VSUBS 0.007363f
C252 B.n141 VSUBS 0.007363f
C253 B.n142 VSUBS 0.007363f
C254 B.n143 VSUBS 0.007363f
C255 B.n144 VSUBS 0.007363f
C256 B.n145 VSUBS 0.007363f
C257 B.n146 VSUBS 0.007363f
C258 B.n147 VSUBS 0.007363f
C259 B.n148 VSUBS 0.007363f
C260 B.n149 VSUBS 0.007363f
C261 B.n150 VSUBS 0.007363f
C262 B.n151 VSUBS 0.007363f
C263 B.n152 VSUBS 0.007363f
C264 B.n153 VSUBS 0.007363f
C265 B.n154 VSUBS 0.007363f
C266 B.n155 VSUBS 0.007363f
C267 B.n156 VSUBS 0.007363f
C268 B.n157 VSUBS 0.007363f
C269 B.n158 VSUBS 0.007363f
C270 B.n159 VSUBS 0.007363f
C271 B.n160 VSUBS 0.007363f
C272 B.n161 VSUBS 0.007363f
C273 B.n162 VSUBS 0.007363f
C274 B.n163 VSUBS 0.007363f
C275 B.n164 VSUBS 0.007363f
C276 B.n165 VSUBS 0.016818f
C277 B.n166 VSUBS 0.017397f
C278 B.n167 VSUBS 0.017397f
C279 B.n168 VSUBS 0.007363f
C280 B.n169 VSUBS 0.007363f
C281 B.n170 VSUBS 0.007363f
C282 B.n171 VSUBS 0.007363f
C283 B.n172 VSUBS 0.007363f
C284 B.n173 VSUBS 0.007363f
C285 B.n174 VSUBS 0.007363f
C286 B.n175 VSUBS 0.007363f
C287 B.n176 VSUBS 0.007363f
C288 B.n177 VSUBS 0.007363f
C289 B.n178 VSUBS 0.007363f
C290 B.n179 VSUBS 0.007363f
C291 B.n180 VSUBS 0.007363f
C292 B.n181 VSUBS 0.007363f
C293 B.n182 VSUBS 0.007363f
C294 B.n183 VSUBS 0.007363f
C295 B.n184 VSUBS 0.007363f
C296 B.n185 VSUBS 0.007363f
C297 B.n186 VSUBS 0.007363f
C298 B.n187 VSUBS 0.007363f
C299 B.n188 VSUBS 0.007363f
C300 B.n189 VSUBS 0.007363f
C301 B.n190 VSUBS 0.007363f
C302 B.n191 VSUBS 0.007363f
C303 B.n192 VSUBS 0.007363f
C304 B.n193 VSUBS 0.007363f
C305 B.n194 VSUBS 0.007363f
C306 B.n195 VSUBS 0.007363f
C307 B.n196 VSUBS 0.007363f
C308 B.n197 VSUBS 0.007363f
C309 B.n198 VSUBS 0.007363f
C310 B.n199 VSUBS 0.007363f
C311 B.n200 VSUBS 0.007363f
C312 B.n201 VSUBS 0.007363f
C313 B.n202 VSUBS 0.007363f
C314 B.n203 VSUBS 0.007363f
C315 B.n204 VSUBS 0.007363f
C316 B.n205 VSUBS 0.007363f
C317 B.n206 VSUBS 0.007363f
C318 B.n207 VSUBS 0.007363f
C319 B.n208 VSUBS 0.007363f
C320 B.n209 VSUBS 0.007363f
C321 B.n210 VSUBS 0.007363f
C322 B.n211 VSUBS 0.007363f
C323 B.n212 VSUBS 0.007363f
C324 B.n213 VSUBS 0.007363f
C325 B.n214 VSUBS 0.007363f
C326 B.n215 VSUBS 0.007363f
C327 B.n216 VSUBS 0.007363f
C328 B.n217 VSUBS 0.007363f
C329 B.n218 VSUBS 0.007363f
C330 B.n219 VSUBS 0.007363f
C331 B.n220 VSUBS 0.007363f
C332 B.n221 VSUBS 0.007363f
C333 B.n222 VSUBS 0.007363f
C334 B.n223 VSUBS 0.007363f
C335 B.n224 VSUBS 0.007363f
C336 B.n225 VSUBS 0.007363f
C337 B.n226 VSUBS 0.007363f
C338 B.n227 VSUBS 0.00693f
C339 B.n228 VSUBS 0.017059f
C340 B.n229 VSUBS 0.004115f
C341 B.n230 VSUBS 0.007363f
C342 B.n231 VSUBS 0.007363f
C343 B.n232 VSUBS 0.007363f
C344 B.n233 VSUBS 0.007363f
C345 B.n234 VSUBS 0.007363f
C346 B.n235 VSUBS 0.007363f
C347 B.n236 VSUBS 0.007363f
C348 B.n237 VSUBS 0.007363f
C349 B.n238 VSUBS 0.007363f
C350 B.n239 VSUBS 0.007363f
C351 B.n240 VSUBS 0.007363f
C352 B.n241 VSUBS 0.007363f
C353 B.t5 VSUBS 0.40715f
C354 B.t4 VSUBS 0.415101f
C355 B.t3 VSUBS 0.322869f
C356 B.n242 VSUBS 0.135381f
C357 B.n243 VSUBS 0.066937f
C358 B.n244 VSUBS 0.017059f
C359 B.n245 VSUBS 0.004115f
C360 B.n246 VSUBS 0.007363f
C361 B.n247 VSUBS 0.007363f
C362 B.n248 VSUBS 0.007363f
C363 B.n249 VSUBS 0.007363f
C364 B.n250 VSUBS 0.007363f
C365 B.n251 VSUBS 0.007363f
C366 B.n252 VSUBS 0.007363f
C367 B.n253 VSUBS 0.007363f
C368 B.n254 VSUBS 0.007363f
C369 B.n255 VSUBS 0.007363f
C370 B.n256 VSUBS 0.007363f
C371 B.n257 VSUBS 0.007363f
C372 B.n258 VSUBS 0.007363f
C373 B.n259 VSUBS 0.007363f
C374 B.n260 VSUBS 0.007363f
C375 B.n261 VSUBS 0.007363f
C376 B.n262 VSUBS 0.007363f
C377 B.n263 VSUBS 0.007363f
C378 B.n264 VSUBS 0.007363f
C379 B.n265 VSUBS 0.007363f
C380 B.n266 VSUBS 0.007363f
C381 B.n267 VSUBS 0.007363f
C382 B.n268 VSUBS 0.007363f
C383 B.n269 VSUBS 0.007363f
C384 B.n270 VSUBS 0.007363f
C385 B.n271 VSUBS 0.007363f
C386 B.n272 VSUBS 0.007363f
C387 B.n273 VSUBS 0.007363f
C388 B.n274 VSUBS 0.007363f
C389 B.n275 VSUBS 0.007363f
C390 B.n276 VSUBS 0.007363f
C391 B.n277 VSUBS 0.007363f
C392 B.n278 VSUBS 0.007363f
C393 B.n279 VSUBS 0.007363f
C394 B.n280 VSUBS 0.007363f
C395 B.n281 VSUBS 0.007363f
C396 B.n282 VSUBS 0.007363f
C397 B.n283 VSUBS 0.007363f
C398 B.n284 VSUBS 0.007363f
C399 B.n285 VSUBS 0.007363f
C400 B.n286 VSUBS 0.007363f
C401 B.n287 VSUBS 0.007363f
C402 B.n288 VSUBS 0.007363f
C403 B.n289 VSUBS 0.007363f
C404 B.n290 VSUBS 0.007363f
C405 B.n291 VSUBS 0.007363f
C406 B.n292 VSUBS 0.007363f
C407 B.n293 VSUBS 0.007363f
C408 B.n294 VSUBS 0.007363f
C409 B.n295 VSUBS 0.007363f
C410 B.n296 VSUBS 0.007363f
C411 B.n297 VSUBS 0.007363f
C412 B.n298 VSUBS 0.007363f
C413 B.n299 VSUBS 0.007363f
C414 B.n300 VSUBS 0.007363f
C415 B.n301 VSUBS 0.007363f
C416 B.n302 VSUBS 0.007363f
C417 B.n303 VSUBS 0.007363f
C418 B.n304 VSUBS 0.007363f
C419 B.n305 VSUBS 0.007363f
C420 B.n306 VSUBS 0.007363f
C421 B.n307 VSUBS 0.017397f
C422 B.n308 VSUBS 0.016818f
C423 B.n309 VSUBS 0.017698f
C424 B.n310 VSUBS 0.007363f
C425 B.n311 VSUBS 0.007363f
C426 B.n312 VSUBS 0.007363f
C427 B.n313 VSUBS 0.007363f
C428 B.n314 VSUBS 0.007363f
C429 B.n315 VSUBS 0.007363f
C430 B.n316 VSUBS 0.007363f
C431 B.n317 VSUBS 0.007363f
C432 B.n318 VSUBS 0.007363f
C433 B.n319 VSUBS 0.007363f
C434 B.n320 VSUBS 0.007363f
C435 B.n321 VSUBS 0.007363f
C436 B.n322 VSUBS 0.007363f
C437 B.n323 VSUBS 0.007363f
C438 B.n324 VSUBS 0.007363f
C439 B.n325 VSUBS 0.007363f
C440 B.n326 VSUBS 0.007363f
C441 B.n327 VSUBS 0.007363f
C442 B.n328 VSUBS 0.007363f
C443 B.n329 VSUBS 0.007363f
C444 B.n330 VSUBS 0.007363f
C445 B.n331 VSUBS 0.007363f
C446 B.n332 VSUBS 0.007363f
C447 B.n333 VSUBS 0.007363f
C448 B.n334 VSUBS 0.007363f
C449 B.n335 VSUBS 0.007363f
C450 B.n336 VSUBS 0.007363f
C451 B.n337 VSUBS 0.007363f
C452 B.n338 VSUBS 0.007363f
C453 B.n339 VSUBS 0.007363f
C454 B.n340 VSUBS 0.007363f
C455 B.n341 VSUBS 0.007363f
C456 B.n342 VSUBS 0.007363f
C457 B.n343 VSUBS 0.007363f
C458 B.n344 VSUBS 0.007363f
C459 B.n345 VSUBS 0.007363f
C460 B.n346 VSUBS 0.007363f
C461 B.n347 VSUBS 0.007363f
C462 B.n348 VSUBS 0.007363f
C463 B.n349 VSUBS 0.007363f
C464 B.n350 VSUBS 0.007363f
C465 B.n351 VSUBS 0.007363f
C466 B.n352 VSUBS 0.007363f
C467 B.n353 VSUBS 0.007363f
C468 B.n354 VSUBS 0.007363f
C469 B.n355 VSUBS 0.007363f
C470 B.n356 VSUBS 0.007363f
C471 B.n357 VSUBS 0.007363f
C472 B.n358 VSUBS 0.007363f
C473 B.n359 VSUBS 0.007363f
C474 B.n360 VSUBS 0.007363f
C475 B.n361 VSUBS 0.007363f
C476 B.n362 VSUBS 0.007363f
C477 B.n363 VSUBS 0.007363f
C478 B.n364 VSUBS 0.007363f
C479 B.n365 VSUBS 0.007363f
C480 B.n366 VSUBS 0.007363f
C481 B.n367 VSUBS 0.016818f
C482 B.n368 VSUBS 0.017397f
C483 B.n369 VSUBS 0.017397f
C484 B.n370 VSUBS 0.007363f
C485 B.n371 VSUBS 0.007363f
C486 B.n372 VSUBS 0.007363f
C487 B.n373 VSUBS 0.007363f
C488 B.n374 VSUBS 0.007363f
C489 B.n375 VSUBS 0.007363f
C490 B.n376 VSUBS 0.007363f
C491 B.n377 VSUBS 0.007363f
C492 B.n378 VSUBS 0.007363f
C493 B.n379 VSUBS 0.007363f
C494 B.n380 VSUBS 0.007363f
C495 B.n381 VSUBS 0.007363f
C496 B.n382 VSUBS 0.007363f
C497 B.n383 VSUBS 0.007363f
C498 B.n384 VSUBS 0.007363f
C499 B.n385 VSUBS 0.007363f
C500 B.n386 VSUBS 0.007363f
C501 B.n387 VSUBS 0.007363f
C502 B.n388 VSUBS 0.007363f
C503 B.n389 VSUBS 0.007363f
C504 B.n390 VSUBS 0.007363f
C505 B.n391 VSUBS 0.007363f
C506 B.n392 VSUBS 0.007363f
C507 B.n393 VSUBS 0.007363f
C508 B.n394 VSUBS 0.007363f
C509 B.n395 VSUBS 0.007363f
C510 B.n396 VSUBS 0.007363f
C511 B.n397 VSUBS 0.007363f
C512 B.n398 VSUBS 0.007363f
C513 B.n399 VSUBS 0.007363f
C514 B.n400 VSUBS 0.007363f
C515 B.n401 VSUBS 0.007363f
C516 B.n402 VSUBS 0.007363f
C517 B.n403 VSUBS 0.007363f
C518 B.n404 VSUBS 0.007363f
C519 B.n405 VSUBS 0.007363f
C520 B.n406 VSUBS 0.007363f
C521 B.n407 VSUBS 0.007363f
C522 B.n408 VSUBS 0.007363f
C523 B.n409 VSUBS 0.007363f
C524 B.n410 VSUBS 0.007363f
C525 B.n411 VSUBS 0.007363f
C526 B.n412 VSUBS 0.007363f
C527 B.n413 VSUBS 0.007363f
C528 B.n414 VSUBS 0.007363f
C529 B.n415 VSUBS 0.007363f
C530 B.n416 VSUBS 0.007363f
C531 B.n417 VSUBS 0.007363f
C532 B.n418 VSUBS 0.007363f
C533 B.n419 VSUBS 0.007363f
C534 B.n420 VSUBS 0.007363f
C535 B.n421 VSUBS 0.007363f
C536 B.n422 VSUBS 0.007363f
C537 B.n423 VSUBS 0.007363f
C538 B.n424 VSUBS 0.007363f
C539 B.n425 VSUBS 0.007363f
C540 B.n426 VSUBS 0.007363f
C541 B.n427 VSUBS 0.007363f
C542 B.n428 VSUBS 0.007363f
C543 B.n429 VSUBS 0.00693f
C544 B.n430 VSUBS 0.017059f
C545 B.n431 VSUBS 0.004115f
C546 B.n432 VSUBS 0.007363f
C547 B.n433 VSUBS 0.007363f
C548 B.n434 VSUBS 0.007363f
C549 B.n435 VSUBS 0.007363f
C550 B.n436 VSUBS 0.007363f
C551 B.n437 VSUBS 0.007363f
C552 B.n438 VSUBS 0.007363f
C553 B.n439 VSUBS 0.007363f
C554 B.n440 VSUBS 0.007363f
C555 B.n441 VSUBS 0.007363f
C556 B.n442 VSUBS 0.007363f
C557 B.n443 VSUBS 0.007363f
C558 B.n444 VSUBS 0.004115f
C559 B.n445 VSUBS 0.007363f
C560 B.n446 VSUBS 0.007363f
C561 B.n447 VSUBS 0.00693f
C562 B.n448 VSUBS 0.007363f
C563 B.n449 VSUBS 0.007363f
C564 B.n450 VSUBS 0.007363f
C565 B.n451 VSUBS 0.007363f
C566 B.n452 VSUBS 0.007363f
C567 B.n453 VSUBS 0.007363f
C568 B.n454 VSUBS 0.007363f
C569 B.n455 VSUBS 0.007363f
C570 B.n456 VSUBS 0.007363f
C571 B.n457 VSUBS 0.007363f
C572 B.n458 VSUBS 0.007363f
C573 B.n459 VSUBS 0.007363f
C574 B.n460 VSUBS 0.007363f
C575 B.n461 VSUBS 0.007363f
C576 B.n462 VSUBS 0.007363f
C577 B.n463 VSUBS 0.007363f
C578 B.n464 VSUBS 0.007363f
C579 B.n465 VSUBS 0.007363f
C580 B.n466 VSUBS 0.007363f
C581 B.n467 VSUBS 0.007363f
C582 B.n468 VSUBS 0.007363f
C583 B.n469 VSUBS 0.007363f
C584 B.n470 VSUBS 0.007363f
C585 B.n471 VSUBS 0.007363f
C586 B.n472 VSUBS 0.007363f
C587 B.n473 VSUBS 0.007363f
C588 B.n474 VSUBS 0.007363f
C589 B.n475 VSUBS 0.007363f
C590 B.n476 VSUBS 0.007363f
C591 B.n477 VSUBS 0.007363f
C592 B.n478 VSUBS 0.007363f
C593 B.n479 VSUBS 0.007363f
C594 B.n480 VSUBS 0.007363f
C595 B.n481 VSUBS 0.007363f
C596 B.n482 VSUBS 0.007363f
C597 B.n483 VSUBS 0.007363f
C598 B.n484 VSUBS 0.007363f
C599 B.n485 VSUBS 0.007363f
C600 B.n486 VSUBS 0.007363f
C601 B.n487 VSUBS 0.007363f
C602 B.n488 VSUBS 0.007363f
C603 B.n489 VSUBS 0.007363f
C604 B.n490 VSUBS 0.007363f
C605 B.n491 VSUBS 0.007363f
C606 B.n492 VSUBS 0.007363f
C607 B.n493 VSUBS 0.007363f
C608 B.n494 VSUBS 0.007363f
C609 B.n495 VSUBS 0.007363f
C610 B.n496 VSUBS 0.007363f
C611 B.n497 VSUBS 0.007363f
C612 B.n498 VSUBS 0.007363f
C613 B.n499 VSUBS 0.007363f
C614 B.n500 VSUBS 0.007363f
C615 B.n501 VSUBS 0.007363f
C616 B.n502 VSUBS 0.007363f
C617 B.n503 VSUBS 0.007363f
C618 B.n504 VSUBS 0.007363f
C619 B.n505 VSUBS 0.007363f
C620 B.n506 VSUBS 0.017397f
C621 B.n507 VSUBS 0.017397f
C622 B.n508 VSUBS 0.016818f
C623 B.n509 VSUBS 0.007363f
C624 B.n510 VSUBS 0.007363f
C625 B.n511 VSUBS 0.007363f
C626 B.n512 VSUBS 0.007363f
C627 B.n513 VSUBS 0.007363f
C628 B.n514 VSUBS 0.007363f
C629 B.n515 VSUBS 0.007363f
C630 B.n516 VSUBS 0.007363f
C631 B.n517 VSUBS 0.007363f
C632 B.n518 VSUBS 0.007363f
C633 B.n519 VSUBS 0.007363f
C634 B.n520 VSUBS 0.007363f
C635 B.n521 VSUBS 0.007363f
C636 B.n522 VSUBS 0.007363f
C637 B.n523 VSUBS 0.007363f
C638 B.n524 VSUBS 0.007363f
C639 B.n525 VSUBS 0.007363f
C640 B.n526 VSUBS 0.007363f
C641 B.n527 VSUBS 0.007363f
C642 B.n528 VSUBS 0.007363f
C643 B.n529 VSUBS 0.007363f
C644 B.n530 VSUBS 0.007363f
C645 B.n531 VSUBS 0.007363f
C646 B.n532 VSUBS 0.007363f
C647 B.n533 VSUBS 0.007363f
C648 B.n534 VSUBS 0.007363f
C649 B.n535 VSUBS 0.009608f
C650 B.n536 VSUBS 0.010235f
C651 B.n537 VSUBS 0.020354f
.ends

