* NGSPICE file created from diff_pair_sample_0725.ext - technology: sky130A

.subckt diff_pair_sample_0725 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t3 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=3.13665 ps=19.34 w=19.01 l=3.59
X1 VDD2.t5 VN.t0 VTAIL.t10 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=3.13665 ps=19.34 w=19.01 l=3.59
X2 VDD2.t4 VN.t1 VTAIL.t0 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=3.13665 ps=19.34 w=19.01 l=3.59
X3 VDD1.t2 VP.t1 VTAIL.t8 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=7.4139 ps=38.8 w=19.01 l=3.59
X4 B.t11 B.t9 B.t10 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=0 ps=0 w=19.01 l=3.59
X5 VTAIL.t11 VN.t2 VDD2.t3 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=3.13665 ps=19.34 w=19.01 l=3.59
X6 B.t8 B.t6 B.t7 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=0 ps=0 w=19.01 l=3.59
X7 B.t5 B.t3 B.t4 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=0 ps=0 w=19.01 l=3.59
X8 VDD1.t5 VP.t2 VTAIL.t7 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=3.13665 ps=19.34 w=19.01 l=3.59
X9 VDD2.t2 VN.t3 VTAIL.t1 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=7.4139 ps=38.8 w=19.01 l=3.59
X10 VTAIL.t3 VN.t4 VDD2.t1 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=3.13665 ps=19.34 w=19.01 l=3.59
X11 VDD1.t4 VP.t3 VTAIL.t6 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=7.4139 ps=38.8 w=19.01 l=3.59
X12 VTAIL.t5 VP.t4 VDD1.t1 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=3.13665 ps=19.34 w=19.01 l=3.59
X13 B.t2 B.t0 B.t1 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=0 ps=0 w=19.01 l=3.59
X14 VDD1.t0 VP.t5 VTAIL.t4 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=7.4139 pd=38.8 as=3.13665 ps=19.34 w=19.01 l=3.59
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n4106_n4770# sky130_fd_pr__pfet_01v8 ad=3.13665 pd=19.34 as=7.4139 ps=38.8 w=19.01 l=3.59
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n55 VP.n54 161.3
R9 VP.n53 VP.n1 161.3
R10 VP.n52 VP.n51 161.3
R11 VP.n50 VP.n2 161.3
R12 VP.n49 VP.n48 161.3
R13 VP.n47 VP.n3 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n4 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n40 VP.n5 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n6 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n7 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n31 VP.n8 161.3
R24 VP.n15 VP.t2 160.728
R25 VP.n29 VP.t5 127.617
R26 VP.n41 VP.t4 127.617
R27 VP.n0 VP.t1 127.617
R28 VP.n9 VP.t3 127.617
R29 VP.n14 VP.t0 127.617
R30 VP.n30 VP.n29 81.7486
R31 VP.n56 VP.n0 81.7486
R32 VP.n28 VP.n9 81.7486
R33 VP.n15 VP.n14 62.3163
R34 VP.n30 VP.n28 57.9539
R35 VP.n35 VP.n6 56.5193
R36 VP.n48 VP.n2 56.5193
R37 VP.n20 VP.n11 56.5193
R38 VP.n33 VP.n8 24.4675
R39 VP.n34 VP.n33 24.4675
R40 VP.n35 VP.n34 24.4675
R41 VP.n39 VP.n6 24.4675
R42 VP.n40 VP.n39 24.4675
R43 VP.n42 VP.n40 24.4675
R44 VP.n46 VP.n4 24.4675
R45 VP.n47 VP.n46 24.4675
R46 VP.n48 VP.n47 24.4675
R47 VP.n52 VP.n2 24.4675
R48 VP.n53 VP.n52 24.4675
R49 VP.n54 VP.n53 24.4675
R50 VP.n24 VP.n11 24.4675
R51 VP.n25 VP.n24 24.4675
R52 VP.n26 VP.n25 24.4675
R53 VP.n18 VP.n13 24.4675
R54 VP.n19 VP.n18 24.4675
R55 VP.n20 VP.n19 24.4675
R56 VP.n42 VP.n41 12.234
R57 VP.n41 VP.n4 12.234
R58 VP.n14 VP.n13 12.234
R59 VP.n29 VP.n8 8.31928
R60 VP.n54 VP.n0 8.31928
R61 VP.n26 VP.n9 8.31928
R62 VP.n16 VP.n15 3.21182
R63 VP.n28 VP.n27 0.354971
R64 VP.n31 VP.n30 0.354971
R65 VP.n56 VP.n55 0.354971
R66 VP VP.n56 0.26696
R67 VP.n17 VP.n16 0.189894
R68 VP.n17 VP.n12 0.189894
R69 VP.n21 VP.n12 0.189894
R70 VP.n22 VP.n21 0.189894
R71 VP.n23 VP.n22 0.189894
R72 VP.n23 VP.n10 0.189894
R73 VP.n27 VP.n10 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n32 VP.n7 0.189894
R76 VP.n36 VP.n7 0.189894
R77 VP.n37 VP.n36 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n38 VP.n5 0.189894
R80 VP.n43 VP.n5 0.189894
R81 VP.n44 VP.n43 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n45 VP.n3 0.189894
R84 VP.n49 VP.n3 0.189894
R85 VP.n50 VP.n49 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n51 VP.n1 0.189894
R88 VP.n55 VP.n1 0.189894
R89 VDD1.n100 VDD1.n0 756.745
R90 VDD1.n205 VDD1.n105 756.745
R91 VDD1.n101 VDD1.n100 585
R92 VDD1.n99 VDD1.n98 585
R93 VDD1.n4 VDD1.n3 585
R94 VDD1.n93 VDD1.n92 585
R95 VDD1.n91 VDD1.n90 585
R96 VDD1.n8 VDD1.n7 585
R97 VDD1.n85 VDD1.n84 585
R98 VDD1.n83 VDD1.n82 585
R99 VDD1.n81 VDD1.n11 585
R100 VDD1.n15 VDD1.n12 585
R101 VDD1.n76 VDD1.n75 585
R102 VDD1.n74 VDD1.n73 585
R103 VDD1.n17 VDD1.n16 585
R104 VDD1.n68 VDD1.n67 585
R105 VDD1.n66 VDD1.n65 585
R106 VDD1.n21 VDD1.n20 585
R107 VDD1.n60 VDD1.n59 585
R108 VDD1.n58 VDD1.n57 585
R109 VDD1.n25 VDD1.n24 585
R110 VDD1.n52 VDD1.n51 585
R111 VDD1.n50 VDD1.n49 585
R112 VDD1.n29 VDD1.n28 585
R113 VDD1.n44 VDD1.n43 585
R114 VDD1.n42 VDD1.n41 585
R115 VDD1.n33 VDD1.n32 585
R116 VDD1.n36 VDD1.n35 585
R117 VDD1.n140 VDD1.n139 585
R118 VDD1.n137 VDD1.n136 585
R119 VDD1.n146 VDD1.n145 585
R120 VDD1.n148 VDD1.n147 585
R121 VDD1.n133 VDD1.n132 585
R122 VDD1.n154 VDD1.n153 585
R123 VDD1.n156 VDD1.n155 585
R124 VDD1.n129 VDD1.n128 585
R125 VDD1.n162 VDD1.n161 585
R126 VDD1.n164 VDD1.n163 585
R127 VDD1.n125 VDD1.n124 585
R128 VDD1.n170 VDD1.n169 585
R129 VDD1.n172 VDD1.n171 585
R130 VDD1.n121 VDD1.n120 585
R131 VDD1.n178 VDD1.n177 585
R132 VDD1.n181 VDD1.n180 585
R133 VDD1.n179 VDD1.n117 585
R134 VDD1.n186 VDD1.n116 585
R135 VDD1.n188 VDD1.n187 585
R136 VDD1.n190 VDD1.n189 585
R137 VDD1.n113 VDD1.n112 585
R138 VDD1.n196 VDD1.n195 585
R139 VDD1.n198 VDD1.n197 585
R140 VDD1.n109 VDD1.n108 585
R141 VDD1.n204 VDD1.n203 585
R142 VDD1.n206 VDD1.n205 585
R143 VDD1.t5 VDD1.n34 327.466
R144 VDD1.t0 VDD1.n138 327.466
R145 VDD1.n100 VDD1.n99 171.744
R146 VDD1.n99 VDD1.n3 171.744
R147 VDD1.n92 VDD1.n3 171.744
R148 VDD1.n92 VDD1.n91 171.744
R149 VDD1.n91 VDD1.n7 171.744
R150 VDD1.n84 VDD1.n7 171.744
R151 VDD1.n84 VDD1.n83 171.744
R152 VDD1.n83 VDD1.n11 171.744
R153 VDD1.n15 VDD1.n11 171.744
R154 VDD1.n75 VDD1.n15 171.744
R155 VDD1.n75 VDD1.n74 171.744
R156 VDD1.n74 VDD1.n16 171.744
R157 VDD1.n67 VDD1.n16 171.744
R158 VDD1.n67 VDD1.n66 171.744
R159 VDD1.n66 VDD1.n20 171.744
R160 VDD1.n59 VDD1.n20 171.744
R161 VDD1.n59 VDD1.n58 171.744
R162 VDD1.n58 VDD1.n24 171.744
R163 VDD1.n51 VDD1.n24 171.744
R164 VDD1.n51 VDD1.n50 171.744
R165 VDD1.n50 VDD1.n28 171.744
R166 VDD1.n43 VDD1.n28 171.744
R167 VDD1.n43 VDD1.n42 171.744
R168 VDD1.n42 VDD1.n32 171.744
R169 VDD1.n35 VDD1.n32 171.744
R170 VDD1.n139 VDD1.n136 171.744
R171 VDD1.n146 VDD1.n136 171.744
R172 VDD1.n147 VDD1.n146 171.744
R173 VDD1.n147 VDD1.n132 171.744
R174 VDD1.n154 VDD1.n132 171.744
R175 VDD1.n155 VDD1.n154 171.744
R176 VDD1.n155 VDD1.n128 171.744
R177 VDD1.n162 VDD1.n128 171.744
R178 VDD1.n163 VDD1.n162 171.744
R179 VDD1.n163 VDD1.n124 171.744
R180 VDD1.n170 VDD1.n124 171.744
R181 VDD1.n171 VDD1.n170 171.744
R182 VDD1.n171 VDD1.n120 171.744
R183 VDD1.n178 VDD1.n120 171.744
R184 VDD1.n180 VDD1.n178 171.744
R185 VDD1.n180 VDD1.n179 171.744
R186 VDD1.n179 VDD1.n116 171.744
R187 VDD1.n188 VDD1.n116 171.744
R188 VDD1.n189 VDD1.n188 171.744
R189 VDD1.n189 VDD1.n112 171.744
R190 VDD1.n196 VDD1.n112 171.744
R191 VDD1.n197 VDD1.n196 171.744
R192 VDD1.n197 VDD1.n108 171.744
R193 VDD1.n204 VDD1.n108 171.744
R194 VDD1.n205 VDD1.n204 171.744
R195 VDD1.n35 VDD1.t5 85.8723
R196 VDD1.n139 VDD1.t0 85.8723
R197 VDD1.n211 VDD1.n210 70.1441
R198 VDD1.n213 VDD1.n212 69.3544
R199 VDD1.n213 VDD1.n211 53.3587
R200 VDD1 VDD1.n104 52.4265
R201 VDD1.n211 VDD1.n209 52.313
R202 VDD1.n36 VDD1.n34 16.3895
R203 VDD1.n140 VDD1.n138 16.3895
R204 VDD1.n82 VDD1.n81 13.1884
R205 VDD1.n187 VDD1.n186 13.1884
R206 VDD1.n85 VDD1.n10 12.8005
R207 VDD1.n80 VDD1.n12 12.8005
R208 VDD1.n37 VDD1.n33 12.8005
R209 VDD1.n141 VDD1.n137 12.8005
R210 VDD1.n185 VDD1.n117 12.8005
R211 VDD1.n190 VDD1.n115 12.8005
R212 VDD1.n86 VDD1.n8 12.0247
R213 VDD1.n77 VDD1.n76 12.0247
R214 VDD1.n41 VDD1.n40 12.0247
R215 VDD1.n145 VDD1.n144 12.0247
R216 VDD1.n182 VDD1.n181 12.0247
R217 VDD1.n191 VDD1.n113 12.0247
R218 VDD1.n90 VDD1.n89 11.249
R219 VDD1.n73 VDD1.n14 11.249
R220 VDD1.n44 VDD1.n31 11.249
R221 VDD1.n148 VDD1.n135 11.249
R222 VDD1.n177 VDD1.n119 11.249
R223 VDD1.n195 VDD1.n194 11.249
R224 VDD1.n93 VDD1.n6 10.4732
R225 VDD1.n72 VDD1.n17 10.4732
R226 VDD1.n45 VDD1.n29 10.4732
R227 VDD1.n149 VDD1.n133 10.4732
R228 VDD1.n176 VDD1.n121 10.4732
R229 VDD1.n198 VDD1.n111 10.4732
R230 VDD1.n94 VDD1.n4 9.69747
R231 VDD1.n69 VDD1.n68 9.69747
R232 VDD1.n49 VDD1.n48 9.69747
R233 VDD1.n153 VDD1.n152 9.69747
R234 VDD1.n173 VDD1.n172 9.69747
R235 VDD1.n199 VDD1.n109 9.69747
R236 VDD1.n104 VDD1.n103 9.45567
R237 VDD1.n209 VDD1.n208 9.45567
R238 VDD1.n62 VDD1.n61 9.3005
R239 VDD1.n64 VDD1.n63 9.3005
R240 VDD1.n19 VDD1.n18 9.3005
R241 VDD1.n70 VDD1.n69 9.3005
R242 VDD1.n72 VDD1.n71 9.3005
R243 VDD1.n14 VDD1.n13 9.3005
R244 VDD1.n78 VDD1.n77 9.3005
R245 VDD1.n80 VDD1.n79 9.3005
R246 VDD1.n103 VDD1.n102 9.3005
R247 VDD1.n2 VDD1.n1 9.3005
R248 VDD1.n97 VDD1.n96 9.3005
R249 VDD1.n95 VDD1.n94 9.3005
R250 VDD1.n6 VDD1.n5 9.3005
R251 VDD1.n89 VDD1.n88 9.3005
R252 VDD1.n87 VDD1.n86 9.3005
R253 VDD1.n10 VDD1.n9 9.3005
R254 VDD1.n23 VDD1.n22 9.3005
R255 VDD1.n56 VDD1.n55 9.3005
R256 VDD1.n54 VDD1.n53 9.3005
R257 VDD1.n27 VDD1.n26 9.3005
R258 VDD1.n48 VDD1.n47 9.3005
R259 VDD1.n46 VDD1.n45 9.3005
R260 VDD1.n31 VDD1.n30 9.3005
R261 VDD1.n40 VDD1.n39 9.3005
R262 VDD1.n38 VDD1.n37 9.3005
R263 VDD1.n107 VDD1.n106 9.3005
R264 VDD1.n202 VDD1.n201 9.3005
R265 VDD1.n200 VDD1.n199 9.3005
R266 VDD1.n111 VDD1.n110 9.3005
R267 VDD1.n194 VDD1.n193 9.3005
R268 VDD1.n192 VDD1.n191 9.3005
R269 VDD1.n115 VDD1.n114 9.3005
R270 VDD1.n160 VDD1.n159 9.3005
R271 VDD1.n158 VDD1.n157 9.3005
R272 VDD1.n131 VDD1.n130 9.3005
R273 VDD1.n152 VDD1.n151 9.3005
R274 VDD1.n150 VDD1.n149 9.3005
R275 VDD1.n135 VDD1.n134 9.3005
R276 VDD1.n144 VDD1.n143 9.3005
R277 VDD1.n142 VDD1.n141 9.3005
R278 VDD1.n127 VDD1.n126 9.3005
R279 VDD1.n166 VDD1.n165 9.3005
R280 VDD1.n168 VDD1.n167 9.3005
R281 VDD1.n123 VDD1.n122 9.3005
R282 VDD1.n174 VDD1.n173 9.3005
R283 VDD1.n176 VDD1.n175 9.3005
R284 VDD1.n119 VDD1.n118 9.3005
R285 VDD1.n183 VDD1.n182 9.3005
R286 VDD1.n185 VDD1.n184 9.3005
R287 VDD1.n208 VDD1.n207 9.3005
R288 VDD1.n98 VDD1.n97 8.92171
R289 VDD1.n65 VDD1.n19 8.92171
R290 VDD1.n52 VDD1.n27 8.92171
R291 VDD1.n156 VDD1.n131 8.92171
R292 VDD1.n169 VDD1.n123 8.92171
R293 VDD1.n203 VDD1.n202 8.92171
R294 VDD1.n101 VDD1.n2 8.14595
R295 VDD1.n64 VDD1.n21 8.14595
R296 VDD1.n53 VDD1.n25 8.14595
R297 VDD1.n157 VDD1.n129 8.14595
R298 VDD1.n168 VDD1.n125 8.14595
R299 VDD1.n206 VDD1.n107 8.14595
R300 VDD1.n102 VDD1.n0 7.3702
R301 VDD1.n61 VDD1.n60 7.3702
R302 VDD1.n57 VDD1.n56 7.3702
R303 VDD1.n161 VDD1.n160 7.3702
R304 VDD1.n165 VDD1.n164 7.3702
R305 VDD1.n207 VDD1.n105 7.3702
R306 VDD1.n104 VDD1.n0 6.59444
R307 VDD1.n60 VDD1.n23 6.59444
R308 VDD1.n57 VDD1.n23 6.59444
R309 VDD1.n161 VDD1.n127 6.59444
R310 VDD1.n164 VDD1.n127 6.59444
R311 VDD1.n209 VDD1.n105 6.59444
R312 VDD1.n102 VDD1.n101 5.81868
R313 VDD1.n61 VDD1.n21 5.81868
R314 VDD1.n56 VDD1.n25 5.81868
R315 VDD1.n160 VDD1.n129 5.81868
R316 VDD1.n165 VDD1.n125 5.81868
R317 VDD1.n207 VDD1.n206 5.81868
R318 VDD1.n98 VDD1.n2 5.04292
R319 VDD1.n65 VDD1.n64 5.04292
R320 VDD1.n53 VDD1.n52 5.04292
R321 VDD1.n157 VDD1.n156 5.04292
R322 VDD1.n169 VDD1.n168 5.04292
R323 VDD1.n203 VDD1.n107 5.04292
R324 VDD1.n97 VDD1.n4 4.26717
R325 VDD1.n68 VDD1.n19 4.26717
R326 VDD1.n49 VDD1.n27 4.26717
R327 VDD1.n153 VDD1.n131 4.26717
R328 VDD1.n172 VDD1.n123 4.26717
R329 VDD1.n202 VDD1.n109 4.26717
R330 VDD1.n38 VDD1.n34 3.70982
R331 VDD1.n142 VDD1.n138 3.70982
R332 VDD1.n94 VDD1.n93 3.49141
R333 VDD1.n69 VDD1.n17 3.49141
R334 VDD1.n48 VDD1.n29 3.49141
R335 VDD1.n152 VDD1.n133 3.49141
R336 VDD1.n173 VDD1.n121 3.49141
R337 VDD1.n199 VDD1.n198 3.49141
R338 VDD1.n90 VDD1.n6 2.71565
R339 VDD1.n73 VDD1.n72 2.71565
R340 VDD1.n45 VDD1.n44 2.71565
R341 VDD1.n149 VDD1.n148 2.71565
R342 VDD1.n177 VDD1.n176 2.71565
R343 VDD1.n195 VDD1.n111 2.71565
R344 VDD1.n89 VDD1.n8 1.93989
R345 VDD1.n76 VDD1.n14 1.93989
R346 VDD1.n41 VDD1.n31 1.93989
R347 VDD1.n145 VDD1.n135 1.93989
R348 VDD1.n181 VDD1.n119 1.93989
R349 VDD1.n194 VDD1.n113 1.93989
R350 VDD1.n212 VDD1.t3 1.71039
R351 VDD1.n212 VDD1.t4 1.71039
R352 VDD1.n210 VDD1.t1 1.71039
R353 VDD1.n210 VDD1.t2 1.71039
R354 VDD1.n86 VDD1.n85 1.16414
R355 VDD1.n77 VDD1.n12 1.16414
R356 VDD1.n40 VDD1.n33 1.16414
R357 VDD1.n144 VDD1.n137 1.16414
R358 VDD1.n182 VDD1.n117 1.16414
R359 VDD1.n191 VDD1.n190 1.16414
R360 VDD1 VDD1.n213 0.787138
R361 VDD1.n82 VDD1.n10 0.388379
R362 VDD1.n81 VDD1.n80 0.388379
R363 VDD1.n37 VDD1.n36 0.388379
R364 VDD1.n141 VDD1.n140 0.388379
R365 VDD1.n186 VDD1.n185 0.388379
R366 VDD1.n187 VDD1.n115 0.388379
R367 VDD1.n103 VDD1.n1 0.155672
R368 VDD1.n96 VDD1.n1 0.155672
R369 VDD1.n96 VDD1.n95 0.155672
R370 VDD1.n95 VDD1.n5 0.155672
R371 VDD1.n88 VDD1.n5 0.155672
R372 VDD1.n88 VDD1.n87 0.155672
R373 VDD1.n87 VDD1.n9 0.155672
R374 VDD1.n79 VDD1.n9 0.155672
R375 VDD1.n79 VDD1.n78 0.155672
R376 VDD1.n78 VDD1.n13 0.155672
R377 VDD1.n71 VDD1.n13 0.155672
R378 VDD1.n71 VDD1.n70 0.155672
R379 VDD1.n70 VDD1.n18 0.155672
R380 VDD1.n63 VDD1.n18 0.155672
R381 VDD1.n63 VDD1.n62 0.155672
R382 VDD1.n62 VDD1.n22 0.155672
R383 VDD1.n55 VDD1.n22 0.155672
R384 VDD1.n55 VDD1.n54 0.155672
R385 VDD1.n54 VDD1.n26 0.155672
R386 VDD1.n47 VDD1.n26 0.155672
R387 VDD1.n47 VDD1.n46 0.155672
R388 VDD1.n46 VDD1.n30 0.155672
R389 VDD1.n39 VDD1.n30 0.155672
R390 VDD1.n39 VDD1.n38 0.155672
R391 VDD1.n143 VDD1.n142 0.155672
R392 VDD1.n143 VDD1.n134 0.155672
R393 VDD1.n150 VDD1.n134 0.155672
R394 VDD1.n151 VDD1.n150 0.155672
R395 VDD1.n151 VDD1.n130 0.155672
R396 VDD1.n158 VDD1.n130 0.155672
R397 VDD1.n159 VDD1.n158 0.155672
R398 VDD1.n159 VDD1.n126 0.155672
R399 VDD1.n166 VDD1.n126 0.155672
R400 VDD1.n167 VDD1.n166 0.155672
R401 VDD1.n167 VDD1.n122 0.155672
R402 VDD1.n174 VDD1.n122 0.155672
R403 VDD1.n175 VDD1.n174 0.155672
R404 VDD1.n175 VDD1.n118 0.155672
R405 VDD1.n183 VDD1.n118 0.155672
R406 VDD1.n184 VDD1.n183 0.155672
R407 VDD1.n184 VDD1.n114 0.155672
R408 VDD1.n192 VDD1.n114 0.155672
R409 VDD1.n193 VDD1.n192 0.155672
R410 VDD1.n193 VDD1.n110 0.155672
R411 VDD1.n200 VDD1.n110 0.155672
R412 VDD1.n201 VDD1.n200 0.155672
R413 VDD1.n201 VDD1.n106 0.155672
R414 VDD1.n208 VDD1.n106 0.155672
R415 VTAIL.n426 VTAIL.n326 756.745
R416 VTAIL.n102 VTAIL.n2 756.745
R417 VTAIL.n320 VTAIL.n220 756.745
R418 VTAIL.n212 VTAIL.n112 756.745
R419 VTAIL.n361 VTAIL.n360 585
R420 VTAIL.n358 VTAIL.n357 585
R421 VTAIL.n367 VTAIL.n366 585
R422 VTAIL.n369 VTAIL.n368 585
R423 VTAIL.n354 VTAIL.n353 585
R424 VTAIL.n375 VTAIL.n374 585
R425 VTAIL.n377 VTAIL.n376 585
R426 VTAIL.n350 VTAIL.n349 585
R427 VTAIL.n383 VTAIL.n382 585
R428 VTAIL.n385 VTAIL.n384 585
R429 VTAIL.n346 VTAIL.n345 585
R430 VTAIL.n391 VTAIL.n390 585
R431 VTAIL.n393 VTAIL.n392 585
R432 VTAIL.n342 VTAIL.n341 585
R433 VTAIL.n399 VTAIL.n398 585
R434 VTAIL.n402 VTAIL.n401 585
R435 VTAIL.n400 VTAIL.n338 585
R436 VTAIL.n407 VTAIL.n337 585
R437 VTAIL.n409 VTAIL.n408 585
R438 VTAIL.n411 VTAIL.n410 585
R439 VTAIL.n334 VTAIL.n333 585
R440 VTAIL.n417 VTAIL.n416 585
R441 VTAIL.n419 VTAIL.n418 585
R442 VTAIL.n330 VTAIL.n329 585
R443 VTAIL.n425 VTAIL.n424 585
R444 VTAIL.n427 VTAIL.n426 585
R445 VTAIL.n37 VTAIL.n36 585
R446 VTAIL.n34 VTAIL.n33 585
R447 VTAIL.n43 VTAIL.n42 585
R448 VTAIL.n45 VTAIL.n44 585
R449 VTAIL.n30 VTAIL.n29 585
R450 VTAIL.n51 VTAIL.n50 585
R451 VTAIL.n53 VTAIL.n52 585
R452 VTAIL.n26 VTAIL.n25 585
R453 VTAIL.n59 VTAIL.n58 585
R454 VTAIL.n61 VTAIL.n60 585
R455 VTAIL.n22 VTAIL.n21 585
R456 VTAIL.n67 VTAIL.n66 585
R457 VTAIL.n69 VTAIL.n68 585
R458 VTAIL.n18 VTAIL.n17 585
R459 VTAIL.n75 VTAIL.n74 585
R460 VTAIL.n78 VTAIL.n77 585
R461 VTAIL.n76 VTAIL.n14 585
R462 VTAIL.n83 VTAIL.n13 585
R463 VTAIL.n85 VTAIL.n84 585
R464 VTAIL.n87 VTAIL.n86 585
R465 VTAIL.n10 VTAIL.n9 585
R466 VTAIL.n93 VTAIL.n92 585
R467 VTAIL.n95 VTAIL.n94 585
R468 VTAIL.n6 VTAIL.n5 585
R469 VTAIL.n101 VTAIL.n100 585
R470 VTAIL.n103 VTAIL.n102 585
R471 VTAIL.n321 VTAIL.n320 585
R472 VTAIL.n319 VTAIL.n318 585
R473 VTAIL.n224 VTAIL.n223 585
R474 VTAIL.n313 VTAIL.n312 585
R475 VTAIL.n311 VTAIL.n310 585
R476 VTAIL.n228 VTAIL.n227 585
R477 VTAIL.n305 VTAIL.n304 585
R478 VTAIL.n303 VTAIL.n302 585
R479 VTAIL.n301 VTAIL.n231 585
R480 VTAIL.n235 VTAIL.n232 585
R481 VTAIL.n296 VTAIL.n295 585
R482 VTAIL.n294 VTAIL.n293 585
R483 VTAIL.n237 VTAIL.n236 585
R484 VTAIL.n288 VTAIL.n287 585
R485 VTAIL.n286 VTAIL.n285 585
R486 VTAIL.n241 VTAIL.n240 585
R487 VTAIL.n280 VTAIL.n279 585
R488 VTAIL.n278 VTAIL.n277 585
R489 VTAIL.n245 VTAIL.n244 585
R490 VTAIL.n272 VTAIL.n271 585
R491 VTAIL.n270 VTAIL.n269 585
R492 VTAIL.n249 VTAIL.n248 585
R493 VTAIL.n264 VTAIL.n263 585
R494 VTAIL.n262 VTAIL.n261 585
R495 VTAIL.n253 VTAIL.n252 585
R496 VTAIL.n256 VTAIL.n255 585
R497 VTAIL.n213 VTAIL.n212 585
R498 VTAIL.n211 VTAIL.n210 585
R499 VTAIL.n116 VTAIL.n115 585
R500 VTAIL.n205 VTAIL.n204 585
R501 VTAIL.n203 VTAIL.n202 585
R502 VTAIL.n120 VTAIL.n119 585
R503 VTAIL.n197 VTAIL.n196 585
R504 VTAIL.n195 VTAIL.n194 585
R505 VTAIL.n193 VTAIL.n123 585
R506 VTAIL.n127 VTAIL.n124 585
R507 VTAIL.n188 VTAIL.n187 585
R508 VTAIL.n186 VTAIL.n185 585
R509 VTAIL.n129 VTAIL.n128 585
R510 VTAIL.n180 VTAIL.n179 585
R511 VTAIL.n178 VTAIL.n177 585
R512 VTAIL.n133 VTAIL.n132 585
R513 VTAIL.n172 VTAIL.n171 585
R514 VTAIL.n170 VTAIL.n169 585
R515 VTAIL.n137 VTAIL.n136 585
R516 VTAIL.n164 VTAIL.n163 585
R517 VTAIL.n162 VTAIL.n161 585
R518 VTAIL.n141 VTAIL.n140 585
R519 VTAIL.n156 VTAIL.n155 585
R520 VTAIL.n154 VTAIL.n153 585
R521 VTAIL.n145 VTAIL.n144 585
R522 VTAIL.n148 VTAIL.n147 585
R523 VTAIL.t6 VTAIL.n254 327.466
R524 VTAIL.t1 VTAIL.n146 327.466
R525 VTAIL.t2 VTAIL.n359 327.466
R526 VTAIL.t8 VTAIL.n35 327.466
R527 VTAIL.n360 VTAIL.n357 171.744
R528 VTAIL.n367 VTAIL.n357 171.744
R529 VTAIL.n368 VTAIL.n367 171.744
R530 VTAIL.n368 VTAIL.n353 171.744
R531 VTAIL.n375 VTAIL.n353 171.744
R532 VTAIL.n376 VTAIL.n375 171.744
R533 VTAIL.n376 VTAIL.n349 171.744
R534 VTAIL.n383 VTAIL.n349 171.744
R535 VTAIL.n384 VTAIL.n383 171.744
R536 VTAIL.n384 VTAIL.n345 171.744
R537 VTAIL.n391 VTAIL.n345 171.744
R538 VTAIL.n392 VTAIL.n391 171.744
R539 VTAIL.n392 VTAIL.n341 171.744
R540 VTAIL.n399 VTAIL.n341 171.744
R541 VTAIL.n401 VTAIL.n399 171.744
R542 VTAIL.n401 VTAIL.n400 171.744
R543 VTAIL.n400 VTAIL.n337 171.744
R544 VTAIL.n409 VTAIL.n337 171.744
R545 VTAIL.n410 VTAIL.n409 171.744
R546 VTAIL.n410 VTAIL.n333 171.744
R547 VTAIL.n417 VTAIL.n333 171.744
R548 VTAIL.n418 VTAIL.n417 171.744
R549 VTAIL.n418 VTAIL.n329 171.744
R550 VTAIL.n425 VTAIL.n329 171.744
R551 VTAIL.n426 VTAIL.n425 171.744
R552 VTAIL.n36 VTAIL.n33 171.744
R553 VTAIL.n43 VTAIL.n33 171.744
R554 VTAIL.n44 VTAIL.n43 171.744
R555 VTAIL.n44 VTAIL.n29 171.744
R556 VTAIL.n51 VTAIL.n29 171.744
R557 VTAIL.n52 VTAIL.n51 171.744
R558 VTAIL.n52 VTAIL.n25 171.744
R559 VTAIL.n59 VTAIL.n25 171.744
R560 VTAIL.n60 VTAIL.n59 171.744
R561 VTAIL.n60 VTAIL.n21 171.744
R562 VTAIL.n67 VTAIL.n21 171.744
R563 VTAIL.n68 VTAIL.n67 171.744
R564 VTAIL.n68 VTAIL.n17 171.744
R565 VTAIL.n75 VTAIL.n17 171.744
R566 VTAIL.n77 VTAIL.n75 171.744
R567 VTAIL.n77 VTAIL.n76 171.744
R568 VTAIL.n76 VTAIL.n13 171.744
R569 VTAIL.n85 VTAIL.n13 171.744
R570 VTAIL.n86 VTAIL.n85 171.744
R571 VTAIL.n86 VTAIL.n9 171.744
R572 VTAIL.n93 VTAIL.n9 171.744
R573 VTAIL.n94 VTAIL.n93 171.744
R574 VTAIL.n94 VTAIL.n5 171.744
R575 VTAIL.n101 VTAIL.n5 171.744
R576 VTAIL.n102 VTAIL.n101 171.744
R577 VTAIL.n320 VTAIL.n319 171.744
R578 VTAIL.n319 VTAIL.n223 171.744
R579 VTAIL.n312 VTAIL.n223 171.744
R580 VTAIL.n312 VTAIL.n311 171.744
R581 VTAIL.n311 VTAIL.n227 171.744
R582 VTAIL.n304 VTAIL.n227 171.744
R583 VTAIL.n304 VTAIL.n303 171.744
R584 VTAIL.n303 VTAIL.n231 171.744
R585 VTAIL.n235 VTAIL.n231 171.744
R586 VTAIL.n295 VTAIL.n235 171.744
R587 VTAIL.n295 VTAIL.n294 171.744
R588 VTAIL.n294 VTAIL.n236 171.744
R589 VTAIL.n287 VTAIL.n236 171.744
R590 VTAIL.n287 VTAIL.n286 171.744
R591 VTAIL.n286 VTAIL.n240 171.744
R592 VTAIL.n279 VTAIL.n240 171.744
R593 VTAIL.n279 VTAIL.n278 171.744
R594 VTAIL.n278 VTAIL.n244 171.744
R595 VTAIL.n271 VTAIL.n244 171.744
R596 VTAIL.n271 VTAIL.n270 171.744
R597 VTAIL.n270 VTAIL.n248 171.744
R598 VTAIL.n263 VTAIL.n248 171.744
R599 VTAIL.n263 VTAIL.n262 171.744
R600 VTAIL.n262 VTAIL.n252 171.744
R601 VTAIL.n255 VTAIL.n252 171.744
R602 VTAIL.n212 VTAIL.n211 171.744
R603 VTAIL.n211 VTAIL.n115 171.744
R604 VTAIL.n204 VTAIL.n115 171.744
R605 VTAIL.n204 VTAIL.n203 171.744
R606 VTAIL.n203 VTAIL.n119 171.744
R607 VTAIL.n196 VTAIL.n119 171.744
R608 VTAIL.n196 VTAIL.n195 171.744
R609 VTAIL.n195 VTAIL.n123 171.744
R610 VTAIL.n127 VTAIL.n123 171.744
R611 VTAIL.n187 VTAIL.n127 171.744
R612 VTAIL.n187 VTAIL.n186 171.744
R613 VTAIL.n186 VTAIL.n128 171.744
R614 VTAIL.n179 VTAIL.n128 171.744
R615 VTAIL.n179 VTAIL.n178 171.744
R616 VTAIL.n178 VTAIL.n132 171.744
R617 VTAIL.n171 VTAIL.n132 171.744
R618 VTAIL.n171 VTAIL.n170 171.744
R619 VTAIL.n170 VTAIL.n136 171.744
R620 VTAIL.n163 VTAIL.n136 171.744
R621 VTAIL.n163 VTAIL.n162 171.744
R622 VTAIL.n162 VTAIL.n140 171.744
R623 VTAIL.n155 VTAIL.n140 171.744
R624 VTAIL.n155 VTAIL.n154 171.744
R625 VTAIL.n154 VTAIL.n144 171.744
R626 VTAIL.n147 VTAIL.n144 171.744
R627 VTAIL.n360 VTAIL.t2 85.8723
R628 VTAIL.n36 VTAIL.t8 85.8723
R629 VTAIL.n255 VTAIL.t6 85.8723
R630 VTAIL.n147 VTAIL.t1 85.8723
R631 VTAIL.n1 VTAIL.n0 52.6758
R632 VTAIL.n109 VTAIL.n108 52.6758
R633 VTAIL.n219 VTAIL.n218 52.6758
R634 VTAIL.n111 VTAIL.n110 52.6758
R635 VTAIL.n111 VTAIL.n109 35.5134
R636 VTAIL.n431 VTAIL.n430 33.155
R637 VTAIL.n107 VTAIL.n106 33.155
R638 VTAIL.n325 VTAIL.n324 33.155
R639 VTAIL.n217 VTAIL.n216 33.155
R640 VTAIL.n431 VTAIL.n325 32.1341
R641 VTAIL.n361 VTAIL.n359 16.3895
R642 VTAIL.n37 VTAIL.n35 16.3895
R643 VTAIL.n256 VTAIL.n254 16.3895
R644 VTAIL.n148 VTAIL.n146 16.3895
R645 VTAIL.n408 VTAIL.n407 13.1884
R646 VTAIL.n84 VTAIL.n83 13.1884
R647 VTAIL.n302 VTAIL.n301 13.1884
R648 VTAIL.n194 VTAIL.n193 13.1884
R649 VTAIL.n362 VTAIL.n358 12.8005
R650 VTAIL.n406 VTAIL.n338 12.8005
R651 VTAIL.n411 VTAIL.n336 12.8005
R652 VTAIL.n38 VTAIL.n34 12.8005
R653 VTAIL.n82 VTAIL.n14 12.8005
R654 VTAIL.n87 VTAIL.n12 12.8005
R655 VTAIL.n305 VTAIL.n230 12.8005
R656 VTAIL.n300 VTAIL.n232 12.8005
R657 VTAIL.n257 VTAIL.n253 12.8005
R658 VTAIL.n197 VTAIL.n122 12.8005
R659 VTAIL.n192 VTAIL.n124 12.8005
R660 VTAIL.n149 VTAIL.n145 12.8005
R661 VTAIL.n366 VTAIL.n365 12.0247
R662 VTAIL.n403 VTAIL.n402 12.0247
R663 VTAIL.n412 VTAIL.n334 12.0247
R664 VTAIL.n42 VTAIL.n41 12.0247
R665 VTAIL.n79 VTAIL.n78 12.0247
R666 VTAIL.n88 VTAIL.n10 12.0247
R667 VTAIL.n306 VTAIL.n228 12.0247
R668 VTAIL.n297 VTAIL.n296 12.0247
R669 VTAIL.n261 VTAIL.n260 12.0247
R670 VTAIL.n198 VTAIL.n120 12.0247
R671 VTAIL.n189 VTAIL.n188 12.0247
R672 VTAIL.n153 VTAIL.n152 12.0247
R673 VTAIL.n369 VTAIL.n356 11.249
R674 VTAIL.n398 VTAIL.n340 11.249
R675 VTAIL.n416 VTAIL.n415 11.249
R676 VTAIL.n45 VTAIL.n32 11.249
R677 VTAIL.n74 VTAIL.n16 11.249
R678 VTAIL.n92 VTAIL.n91 11.249
R679 VTAIL.n310 VTAIL.n309 11.249
R680 VTAIL.n293 VTAIL.n234 11.249
R681 VTAIL.n264 VTAIL.n251 11.249
R682 VTAIL.n202 VTAIL.n201 11.249
R683 VTAIL.n185 VTAIL.n126 11.249
R684 VTAIL.n156 VTAIL.n143 11.249
R685 VTAIL.n370 VTAIL.n354 10.4732
R686 VTAIL.n397 VTAIL.n342 10.4732
R687 VTAIL.n419 VTAIL.n332 10.4732
R688 VTAIL.n46 VTAIL.n30 10.4732
R689 VTAIL.n73 VTAIL.n18 10.4732
R690 VTAIL.n95 VTAIL.n8 10.4732
R691 VTAIL.n313 VTAIL.n226 10.4732
R692 VTAIL.n292 VTAIL.n237 10.4732
R693 VTAIL.n265 VTAIL.n249 10.4732
R694 VTAIL.n205 VTAIL.n118 10.4732
R695 VTAIL.n184 VTAIL.n129 10.4732
R696 VTAIL.n157 VTAIL.n141 10.4732
R697 VTAIL.n374 VTAIL.n373 9.69747
R698 VTAIL.n394 VTAIL.n393 9.69747
R699 VTAIL.n420 VTAIL.n330 9.69747
R700 VTAIL.n50 VTAIL.n49 9.69747
R701 VTAIL.n70 VTAIL.n69 9.69747
R702 VTAIL.n96 VTAIL.n6 9.69747
R703 VTAIL.n314 VTAIL.n224 9.69747
R704 VTAIL.n289 VTAIL.n288 9.69747
R705 VTAIL.n269 VTAIL.n268 9.69747
R706 VTAIL.n206 VTAIL.n116 9.69747
R707 VTAIL.n181 VTAIL.n180 9.69747
R708 VTAIL.n161 VTAIL.n160 9.69747
R709 VTAIL.n430 VTAIL.n429 9.45567
R710 VTAIL.n106 VTAIL.n105 9.45567
R711 VTAIL.n324 VTAIL.n323 9.45567
R712 VTAIL.n216 VTAIL.n215 9.45567
R713 VTAIL.n328 VTAIL.n327 9.3005
R714 VTAIL.n423 VTAIL.n422 9.3005
R715 VTAIL.n421 VTAIL.n420 9.3005
R716 VTAIL.n332 VTAIL.n331 9.3005
R717 VTAIL.n415 VTAIL.n414 9.3005
R718 VTAIL.n413 VTAIL.n412 9.3005
R719 VTAIL.n336 VTAIL.n335 9.3005
R720 VTAIL.n381 VTAIL.n380 9.3005
R721 VTAIL.n379 VTAIL.n378 9.3005
R722 VTAIL.n352 VTAIL.n351 9.3005
R723 VTAIL.n373 VTAIL.n372 9.3005
R724 VTAIL.n371 VTAIL.n370 9.3005
R725 VTAIL.n356 VTAIL.n355 9.3005
R726 VTAIL.n365 VTAIL.n364 9.3005
R727 VTAIL.n363 VTAIL.n362 9.3005
R728 VTAIL.n348 VTAIL.n347 9.3005
R729 VTAIL.n387 VTAIL.n386 9.3005
R730 VTAIL.n389 VTAIL.n388 9.3005
R731 VTAIL.n344 VTAIL.n343 9.3005
R732 VTAIL.n395 VTAIL.n394 9.3005
R733 VTAIL.n397 VTAIL.n396 9.3005
R734 VTAIL.n340 VTAIL.n339 9.3005
R735 VTAIL.n404 VTAIL.n403 9.3005
R736 VTAIL.n406 VTAIL.n405 9.3005
R737 VTAIL.n429 VTAIL.n428 9.3005
R738 VTAIL.n4 VTAIL.n3 9.3005
R739 VTAIL.n99 VTAIL.n98 9.3005
R740 VTAIL.n97 VTAIL.n96 9.3005
R741 VTAIL.n8 VTAIL.n7 9.3005
R742 VTAIL.n91 VTAIL.n90 9.3005
R743 VTAIL.n89 VTAIL.n88 9.3005
R744 VTAIL.n12 VTAIL.n11 9.3005
R745 VTAIL.n57 VTAIL.n56 9.3005
R746 VTAIL.n55 VTAIL.n54 9.3005
R747 VTAIL.n28 VTAIL.n27 9.3005
R748 VTAIL.n49 VTAIL.n48 9.3005
R749 VTAIL.n47 VTAIL.n46 9.3005
R750 VTAIL.n32 VTAIL.n31 9.3005
R751 VTAIL.n41 VTAIL.n40 9.3005
R752 VTAIL.n39 VTAIL.n38 9.3005
R753 VTAIL.n24 VTAIL.n23 9.3005
R754 VTAIL.n63 VTAIL.n62 9.3005
R755 VTAIL.n65 VTAIL.n64 9.3005
R756 VTAIL.n20 VTAIL.n19 9.3005
R757 VTAIL.n71 VTAIL.n70 9.3005
R758 VTAIL.n73 VTAIL.n72 9.3005
R759 VTAIL.n16 VTAIL.n15 9.3005
R760 VTAIL.n80 VTAIL.n79 9.3005
R761 VTAIL.n82 VTAIL.n81 9.3005
R762 VTAIL.n105 VTAIL.n104 9.3005
R763 VTAIL.n282 VTAIL.n281 9.3005
R764 VTAIL.n284 VTAIL.n283 9.3005
R765 VTAIL.n239 VTAIL.n238 9.3005
R766 VTAIL.n290 VTAIL.n289 9.3005
R767 VTAIL.n292 VTAIL.n291 9.3005
R768 VTAIL.n234 VTAIL.n233 9.3005
R769 VTAIL.n298 VTAIL.n297 9.3005
R770 VTAIL.n300 VTAIL.n299 9.3005
R771 VTAIL.n323 VTAIL.n322 9.3005
R772 VTAIL.n222 VTAIL.n221 9.3005
R773 VTAIL.n317 VTAIL.n316 9.3005
R774 VTAIL.n315 VTAIL.n314 9.3005
R775 VTAIL.n226 VTAIL.n225 9.3005
R776 VTAIL.n309 VTAIL.n308 9.3005
R777 VTAIL.n307 VTAIL.n306 9.3005
R778 VTAIL.n230 VTAIL.n229 9.3005
R779 VTAIL.n243 VTAIL.n242 9.3005
R780 VTAIL.n276 VTAIL.n275 9.3005
R781 VTAIL.n274 VTAIL.n273 9.3005
R782 VTAIL.n247 VTAIL.n246 9.3005
R783 VTAIL.n268 VTAIL.n267 9.3005
R784 VTAIL.n266 VTAIL.n265 9.3005
R785 VTAIL.n251 VTAIL.n250 9.3005
R786 VTAIL.n260 VTAIL.n259 9.3005
R787 VTAIL.n258 VTAIL.n257 9.3005
R788 VTAIL.n174 VTAIL.n173 9.3005
R789 VTAIL.n176 VTAIL.n175 9.3005
R790 VTAIL.n131 VTAIL.n130 9.3005
R791 VTAIL.n182 VTAIL.n181 9.3005
R792 VTAIL.n184 VTAIL.n183 9.3005
R793 VTAIL.n126 VTAIL.n125 9.3005
R794 VTAIL.n190 VTAIL.n189 9.3005
R795 VTAIL.n192 VTAIL.n191 9.3005
R796 VTAIL.n215 VTAIL.n214 9.3005
R797 VTAIL.n114 VTAIL.n113 9.3005
R798 VTAIL.n209 VTAIL.n208 9.3005
R799 VTAIL.n207 VTAIL.n206 9.3005
R800 VTAIL.n118 VTAIL.n117 9.3005
R801 VTAIL.n201 VTAIL.n200 9.3005
R802 VTAIL.n199 VTAIL.n198 9.3005
R803 VTAIL.n122 VTAIL.n121 9.3005
R804 VTAIL.n135 VTAIL.n134 9.3005
R805 VTAIL.n168 VTAIL.n167 9.3005
R806 VTAIL.n166 VTAIL.n165 9.3005
R807 VTAIL.n139 VTAIL.n138 9.3005
R808 VTAIL.n160 VTAIL.n159 9.3005
R809 VTAIL.n158 VTAIL.n157 9.3005
R810 VTAIL.n143 VTAIL.n142 9.3005
R811 VTAIL.n152 VTAIL.n151 9.3005
R812 VTAIL.n150 VTAIL.n149 9.3005
R813 VTAIL.n377 VTAIL.n352 8.92171
R814 VTAIL.n390 VTAIL.n344 8.92171
R815 VTAIL.n424 VTAIL.n423 8.92171
R816 VTAIL.n53 VTAIL.n28 8.92171
R817 VTAIL.n66 VTAIL.n20 8.92171
R818 VTAIL.n100 VTAIL.n99 8.92171
R819 VTAIL.n318 VTAIL.n317 8.92171
R820 VTAIL.n285 VTAIL.n239 8.92171
R821 VTAIL.n272 VTAIL.n247 8.92171
R822 VTAIL.n210 VTAIL.n209 8.92171
R823 VTAIL.n177 VTAIL.n131 8.92171
R824 VTAIL.n164 VTAIL.n139 8.92171
R825 VTAIL.n378 VTAIL.n350 8.14595
R826 VTAIL.n389 VTAIL.n346 8.14595
R827 VTAIL.n427 VTAIL.n328 8.14595
R828 VTAIL.n54 VTAIL.n26 8.14595
R829 VTAIL.n65 VTAIL.n22 8.14595
R830 VTAIL.n103 VTAIL.n4 8.14595
R831 VTAIL.n321 VTAIL.n222 8.14595
R832 VTAIL.n284 VTAIL.n241 8.14595
R833 VTAIL.n273 VTAIL.n245 8.14595
R834 VTAIL.n213 VTAIL.n114 8.14595
R835 VTAIL.n176 VTAIL.n133 8.14595
R836 VTAIL.n165 VTAIL.n137 8.14595
R837 VTAIL.n382 VTAIL.n381 7.3702
R838 VTAIL.n386 VTAIL.n385 7.3702
R839 VTAIL.n428 VTAIL.n326 7.3702
R840 VTAIL.n58 VTAIL.n57 7.3702
R841 VTAIL.n62 VTAIL.n61 7.3702
R842 VTAIL.n104 VTAIL.n2 7.3702
R843 VTAIL.n322 VTAIL.n220 7.3702
R844 VTAIL.n281 VTAIL.n280 7.3702
R845 VTAIL.n277 VTAIL.n276 7.3702
R846 VTAIL.n214 VTAIL.n112 7.3702
R847 VTAIL.n173 VTAIL.n172 7.3702
R848 VTAIL.n169 VTAIL.n168 7.3702
R849 VTAIL.n382 VTAIL.n348 6.59444
R850 VTAIL.n385 VTAIL.n348 6.59444
R851 VTAIL.n430 VTAIL.n326 6.59444
R852 VTAIL.n58 VTAIL.n24 6.59444
R853 VTAIL.n61 VTAIL.n24 6.59444
R854 VTAIL.n106 VTAIL.n2 6.59444
R855 VTAIL.n324 VTAIL.n220 6.59444
R856 VTAIL.n280 VTAIL.n243 6.59444
R857 VTAIL.n277 VTAIL.n243 6.59444
R858 VTAIL.n216 VTAIL.n112 6.59444
R859 VTAIL.n172 VTAIL.n135 6.59444
R860 VTAIL.n169 VTAIL.n135 6.59444
R861 VTAIL.n381 VTAIL.n350 5.81868
R862 VTAIL.n386 VTAIL.n346 5.81868
R863 VTAIL.n428 VTAIL.n427 5.81868
R864 VTAIL.n57 VTAIL.n26 5.81868
R865 VTAIL.n62 VTAIL.n22 5.81868
R866 VTAIL.n104 VTAIL.n103 5.81868
R867 VTAIL.n322 VTAIL.n321 5.81868
R868 VTAIL.n281 VTAIL.n241 5.81868
R869 VTAIL.n276 VTAIL.n245 5.81868
R870 VTAIL.n214 VTAIL.n213 5.81868
R871 VTAIL.n173 VTAIL.n133 5.81868
R872 VTAIL.n168 VTAIL.n137 5.81868
R873 VTAIL.n378 VTAIL.n377 5.04292
R874 VTAIL.n390 VTAIL.n389 5.04292
R875 VTAIL.n424 VTAIL.n328 5.04292
R876 VTAIL.n54 VTAIL.n53 5.04292
R877 VTAIL.n66 VTAIL.n65 5.04292
R878 VTAIL.n100 VTAIL.n4 5.04292
R879 VTAIL.n318 VTAIL.n222 5.04292
R880 VTAIL.n285 VTAIL.n284 5.04292
R881 VTAIL.n273 VTAIL.n272 5.04292
R882 VTAIL.n210 VTAIL.n114 5.04292
R883 VTAIL.n177 VTAIL.n176 5.04292
R884 VTAIL.n165 VTAIL.n164 5.04292
R885 VTAIL.n374 VTAIL.n352 4.26717
R886 VTAIL.n393 VTAIL.n344 4.26717
R887 VTAIL.n423 VTAIL.n330 4.26717
R888 VTAIL.n50 VTAIL.n28 4.26717
R889 VTAIL.n69 VTAIL.n20 4.26717
R890 VTAIL.n99 VTAIL.n6 4.26717
R891 VTAIL.n317 VTAIL.n224 4.26717
R892 VTAIL.n288 VTAIL.n239 4.26717
R893 VTAIL.n269 VTAIL.n247 4.26717
R894 VTAIL.n209 VTAIL.n116 4.26717
R895 VTAIL.n180 VTAIL.n131 4.26717
R896 VTAIL.n161 VTAIL.n139 4.26717
R897 VTAIL.n363 VTAIL.n359 3.70982
R898 VTAIL.n39 VTAIL.n35 3.70982
R899 VTAIL.n258 VTAIL.n254 3.70982
R900 VTAIL.n150 VTAIL.n146 3.70982
R901 VTAIL.n373 VTAIL.n354 3.49141
R902 VTAIL.n394 VTAIL.n342 3.49141
R903 VTAIL.n420 VTAIL.n419 3.49141
R904 VTAIL.n49 VTAIL.n30 3.49141
R905 VTAIL.n70 VTAIL.n18 3.49141
R906 VTAIL.n96 VTAIL.n95 3.49141
R907 VTAIL.n314 VTAIL.n313 3.49141
R908 VTAIL.n289 VTAIL.n237 3.49141
R909 VTAIL.n268 VTAIL.n249 3.49141
R910 VTAIL.n206 VTAIL.n205 3.49141
R911 VTAIL.n181 VTAIL.n129 3.49141
R912 VTAIL.n160 VTAIL.n141 3.49141
R913 VTAIL.n217 VTAIL.n111 3.37981
R914 VTAIL.n325 VTAIL.n219 3.37981
R915 VTAIL.n109 VTAIL.n107 3.37981
R916 VTAIL.n370 VTAIL.n369 2.71565
R917 VTAIL.n398 VTAIL.n397 2.71565
R918 VTAIL.n416 VTAIL.n332 2.71565
R919 VTAIL.n46 VTAIL.n45 2.71565
R920 VTAIL.n74 VTAIL.n73 2.71565
R921 VTAIL.n92 VTAIL.n8 2.71565
R922 VTAIL.n310 VTAIL.n226 2.71565
R923 VTAIL.n293 VTAIL.n292 2.71565
R924 VTAIL.n265 VTAIL.n264 2.71565
R925 VTAIL.n202 VTAIL.n118 2.71565
R926 VTAIL.n185 VTAIL.n184 2.71565
R927 VTAIL.n157 VTAIL.n156 2.71565
R928 VTAIL VTAIL.n431 2.47679
R929 VTAIL.n219 VTAIL.n217 2.15998
R930 VTAIL.n107 VTAIL.n1 2.15998
R931 VTAIL.n366 VTAIL.n356 1.93989
R932 VTAIL.n402 VTAIL.n340 1.93989
R933 VTAIL.n415 VTAIL.n334 1.93989
R934 VTAIL.n42 VTAIL.n32 1.93989
R935 VTAIL.n78 VTAIL.n16 1.93989
R936 VTAIL.n91 VTAIL.n10 1.93989
R937 VTAIL.n309 VTAIL.n228 1.93989
R938 VTAIL.n296 VTAIL.n234 1.93989
R939 VTAIL.n261 VTAIL.n251 1.93989
R940 VTAIL.n201 VTAIL.n120 1.93989
R941 VTAIL.n188 VTAIL.n126 1.93989
R942 VTAIL.n153 VTAIL.n143 1.93989
R943 VTAIL.n0 VTAIL.t0 1.71039
R944 VTAIL.n0 VTAIL.t3 1.71039
R945 VTAIL.n108 VTAIL.t4 1.71039
R946 VTAIL.n108 VTAIL.t5 1.71039
R947 VTAIL.n218 VTAIL.t7 1.71039
R948 VTAIL.n218 VTAIL.t9 1.71039
R949 VTAIL.n110 VTAIL.t10 1.71039
R950 VTAIL.n110 VTAIL.t11 1.71039
R951 VTAIL.n365 VTAIL.n358 1.16414
R952 VTAIL.n403 VTAIL.n338 1.16414
R953 VTAIL.n412 VTAIL.n411 1.16414
R954 VTAIL.n41 VTAIL.n34 1.16414
R955 VTAIL.n79 VTAIL.n14 1.16414
R956 VTAIL.n88 VTAIL.n87 1.16414
R957 VTAIL.n306 VTAIL.n305 1.16414
R958 VTAIL.n297 VTAIL.n232 1.16414
R959 VTAIL.n260 VTAIL.n253 1.16414
R960 VTAIL.n198 VTAIL.n197 1.16414
R961 VTAIL.n189 VTAIL.n124 1.16414
R962 VTAIL.n152 VTAIL.n145 1.16414
R963 VTAIL VTAIL.n1 0.903517
R964 VTAIL.n362 VTAIL.n361 0.388379
R965 VTAIL.n407 VTAIL.n406 0.388379
R966 VTAIL.n408 VTAIL.n336 0.388379
R967 VTAIL.n38 VTAIL.n37 0.388379
R968 VTAIL.n83 VTAIL.n82 0.388379
R969 VTAIL.n84 VTAIL.n12 0.388379
R970 VTAIL.n302 VTAIL.n230 0.388379
R971 VTAIL.n301 VTAIL.n300 0.388379
R972 VTAIL.n257 VTAIL.n256 0.388379
R973 VTAIL.n194 VTAIL.n122 0.388379
R974 VTAIL.n193 VTAIL.n192 0.388379
R975 VTAIL.n149 VTAIL.n148 0.388379
R976 VTAIL.n364 VTAIL.n363 0.155672
R977 VTAIL.n364 VTAIL.n355 0.155672
R978 VTAIL.n371 VTAIL.n355 0.155672
R979 VTAIL.n372 VTAIL.n371 0.155672
R980 VTAIL.n372 VTAIL.n351 0.155672
R981 VTAIL.n379 VTAIL.n351 0.155672
R982 VTAIL.n380 VTAIL.n379 0.155672
R983 VTAIL.n380 VTAIL.n347 0.155672
R984 VTAIL.n387 VTAIL.n347 0.155672
R985 VTAIL.n388 VTAIL.n387 0.155672
R986 VTAIL.n388 VTAIL.n343 0.155672
R987 VTAIL.n395 VTAIL.n343 0.155672
R988 VTAIL.n396 VTAIL.n395 0.155672
R989 VTAIL.n396 VTAIL.n339 0.155672
R990 VTAIL.n404 VTAIL.n339 0.155672
R991 VTAIL.n405 VTAIL.n404 0.155672
R992 VTAIL.n405 VTAIL.n335 0.155672
R993 VTAIL.n413 VTAIL.n335 0.155672
R994 VTAIL.n414 VTAIL.n413 0.155672
R995 VTAIL.n414 VTAIL.n331 0.155672
R996 VTAIL.n421 VTAIL.n331 0.155672
R997 VTAIL.n422 VTAIL.n421 0.155672
R998 VTAIL.n422 VTAIL.n327 0.155672
R999 VTAIL.n429 VTAIL.n327 0.155672
R1000 VTAIL.n40 VTAIL.n39 0.155672
R1001 VTAIL.n40 VTAIL.n31 0.155672
R1002 VTAIL.n47 VTAIL.n31 0.155672
R1003 VTAIL.n48 VTAIL.n47 0.155672
R1004 VTAIL.n48 VTAIL.n27 0.155672
R1005 VTAIL.n55 VTAIL.n27 0.155672
R1006 VTAIL.n56 VTAIL.n55 0.155672
R1007 VTAIL.n56 VTAIL.n23 0.155672
R1008 VTAIL.n63 VTAIL.n23 0.155672
R1009 VTAIL.n64 VTAIL.n63 0.155672
R1010 VTAIL.n64 VTAIL.n19 0.155672
R1011 VTAIL.n71 VTAIL.n19 0.155672
R1012 VTAIL.n72 VTAIL.n71 0.155672
R1013 VTAIL.n72 VTAIL.n15 0.155672
R1014 VTAIL.n80 VTAIL.n15 0.155672
R1015 VTAIL.n81 VTAIL.n80 0.155672
R1016 VTAIL.n81 VTAIL.n11 0.155672
R1017 VTAIL.n89 VTAIL.n11 0.155672
R1018 VTAIL.n90 VTAIL.n89 0.155672
R1019 VTAIL.n90 VTAIL.n7 0.155672
R1020 VTAIL.n97 VTAIL.n7 0.155672
R1021 VTAIL.n98 VTAIL.n97 0.155672
R1022 VTAIL.n98 VTAIL.n3 0.155672
R1023 VTAIL.n105 VTAIL.n3 0.155672
R1024 VTAIL.n323 VTAIL.n221 0.155672
R1025 VTAIL.n316 VTAIL.n221 0.155672
R1026 VTAIL.n316 VTAIL.n315 0.155672
R1027 VTAIL.n315 VTAIL.n225 0.155672
R1028 VTAIL.n308 VTAIL.n225 0.155672
R1029 VTAIL.n308 VTAIL.n307 0.155672
R1030 VTAIL.n307 VTAIL.n229 0.155672
R1031 VTAIL.n299 VTAIL.n229 0.155672
R1032 VTAIL.n299 VTAIL.n298 0.155672
R1033 VTAIL.n298 VTAIL.n233 0.155672
R1034 VTAIL.n291 VTAIL.n233 0.155672
R1035 VTAIL.n291 VTAIL.n290 0.155672
R1036 VTAIL.n290 VTAIL.n238 0.155672
R1037 VTAIL.n283 VTAIL.n238 0.155672
R1038 VTAIL.n283 VTAIL.n282 0.155672
R1039 VTAIL.n282 VTAIL.n242 0.155672
R1040 VTAIL.n275 VTAIL.n242 0.155672
R1041 VTAIL.n275 VTAIL.n274 0.155672
R1042 VTAIL.n274 VTAIL.n246 0.155672
R1043 VTAIL.n267 VTAIL.n246 0.155672
R1044 VTAIL.n267 VTAIL.n266 0.155672
R1045 VTAIL.n266 VTAIL.n250 0.155672
R1046 VTAIL.n259 VTAIL.n250 0.155672
R1047 VTAIL.n259 VTAIL.n258 0.155672
R1048 VTAIL.n215 VTAIL.n113 0.155672
R1049 VTAIL.n208 VTAIL.n113 0.155672
R1050 VTAIL.n208 VTAIL.n207 0.155672
R1051 VTAIL.n207 VTAIL.n117 0.155672
R1052 VTAIL.n200 VTAIL.n117 0.155672
R1053 VTAIL.n200 VTAIL.n199 0.155672
R1054 VTAIL.n199 VTAIL.n121 0.155672
R1055 VTAIL.n191 VTAIL.n121 0.155672
R1056 VTAIL.n191 VTAIL.n190 0.155672
R1057 VTAIL.n190 VTAIL.n125 0.155672
R1058 VTAIL.n183 VTAIL.n125 0.155672
R1059 VTAIL.n183 VTAIL.n182 0.155672
R1060 VTAIL.n182 VTAIL.n130 0.155672
R1061 VTAIL.n175 VTAIL.n130 0.155672
R1062 VTAIL.n175 VTAIL.n174 0.155672
R1063 VTAIL.n174 VTAIL.n134 0.155672
R1064 VTAIL.n167 VTAIL.n134 0.155672
R1065 VTAIL.n167 VTAIL.n166 0.155672
R1066 VTAIL.n166 VTAIL.n138 0.155672
R1067 VTAIL.n159 VTAIL.n138 0.155672
R1068 VTAIL.n159 VTAIL.n158 0.155672
R1069 VTAIL.n158 VTAIL.n142 0.155672
R1070 VTAIL.n151 VTAIL.n142 0.155672
R1071 VTAIL.n151 VTAIL.n150 0.155672
R1072 VN.n38 VN.n37 161.3
R1073 VN.n36 VN.n21 161.3
R1074 VN.n35 VN.n34 161.3
R1075 VN.n33 VN.n22 161.3
R1076 VN.n32 VN.n31 161.3
R1077 VN.n30 VN.n23 161.3
R1078 VN.n29 VN.n28 161.3
R1079 VN.n27 VN.n24 161.3
R1080 VN.n18 VN.n17 161.3
R1081 VN.n16 VN.n1 161.3
R1082 VN.n15 VN.n14 161.3
R1083 VN.n13 VN.n2 161.3
R1084 VN.n12 VN.n11 161.3
R1085 VN.n10 VN.n3 161.3
R1086 VN.n9 VN.n8 161.3
R1087 VN.n7 VN.n4 161.3
R1088 VN.n26 VN.t3 160.728
R1089 VN.n6 VN.t1 160.728
R1090 VN.n5 VN.t4 127.617
R1091 VN.n0 VN.t5 127.617
R1092 VN.n25 VN.t2 127.617
R1093 VN.n20 VN.t0 127.617
R1094 VN.n19 VN.n0 81.7486
R1095 VN.n39 VN.n20 81.7486
R1096 VN.n26 VN.n25 62.3163
R1097 VN.n6 VN.n5 62.3162
R1098 VN VN.n39 58.1192
R1099 VN.n11 VN.n2 56.5193
R1100 VN.n31 VN.n22 56.5193
R1101 VN.n9 VN.n4 24.4675
R1102 VN.n10 VN.n9 24.4675
R1103 VN.n11 VN.n10 24.4675
R1104 VN.n15 VN.n2 24.4675
R1105 VN.n16 VN.n15 24.4675
R1106 VN.n17 VN.n16 24.4675
R1107 VN.n31 VN.n30 24.4675
R1108 VN.n30 VN.n29 24.4675
R1109 VN.n29 VN.n24 24.4675
R1110 VN.n37 VN.n36 24.4675
R1111 VN.n36 VN.n35 24.4675
R1112 VN.n35 VN.n22 24.4675
R1113 VN.n5 VN.n4 12.234
R1114 VN.n25 VN.n24 12.234
R1115 VN.n17 VN.n0 8.31928
R1116 VN.n37 VN.n20 8.31928
R1117 VN.n7 VN.n6 3.21184
R1118 VN.n27 VN.n26 3.21184
R1119 VN.n39 VN.n38 0.354971
R1120 VN.n19 VN.n18 0.354971
R1121 VN VN.n19 0.26696
R1122 VN.n38 VN.n21 0.189894
R1123 VN.n34 VN.n21 0.189894
R1124 VN.n34 VN.n33 0.189894
R1125 VN.n33 VN.n32 0.189894
R1126 VN.n32 VN.n23 0.189894
R1127 VN.n28 VN.n23 0.189894
R1128 VN.n28 VN.n27 0.189894
R1129 VN.n8 VN.n7 0.189894
R1130 VN.n8 VN.n3 0.189894
R1131 VN.n12 VN.n3 0.189894
R1132 VN.n13 VN.n12 0.189894
R1133 VN.n14 VN.n13 0.189894
R1134 VN.n14 VN.n1 0.189894
R1135 VN.n18 VN.n1 0.189894
R1136 VDD2.n207 VDD2.n107 756.745
R1137 VDD2.n100 VDD2.n0 756.745
R1138 VDD2.n208 VDD2.n207 585
R1139 VDD2.n206 VDD2.n205 585
R1140 VDD2.n111 VDD2.n110 585
R1141 VDD2.n200 VDD2.n199 585
R1142 VDD2.n198 VDD2.n197 585
R1143 VDD2.n115 VDD2.n114 585
R1144 VDD2.n192 VDD2.n191 585
R1145 VDD2.n190 VDD2.n189 585
R1146 VDD2.n188 VDD2.n118 585
R1147 VDD2.n122 VDD2.n119 585
R1148 VDD2.n183 VDD2.n182 585
R1149 VDD2.n181 VDD2.n180 585
R1150 VDD2.n124 VDD2.n123 585
R1151 VDD2.n175 VDD2.n174 585
R1152 VDD2.n173 VDD2.n172 585
R1153 VDD2.n128 VDD2.n127 585
R1154 VDD2.n167 VDD2.n166 585
R1155 VDD2.n165 VDD2.n164 585
R1156 VDD2.n132 VDD2.n131 585
R1157 VDD2.n159 VDD2.n158 585
R1158 VDD2.n157 VDD2.n156 585
R1159 VDD2.n136 VDD2.n135 585
R1160 VDD2.n151 VDD2.n150 585
R1161 VDD2.n149 VDD2.n148 585
R1162 VDD2.n140 VDD2.n139 585
R1163 VDD2.n143 VDD2.n142 585
R1164 VDD2.n35 VDD2.n34 585
R1165 VDD2.n32 VDD2.n31 585
R1166 VDD2.n41 VDD2.n40 585
R1167 VDD2.n43 VDD2.n42 585
R1168 VDD2.n28 VDD2.n27 585
R1169 VDD2.n49 VDD2.n48 585
R1170 VDD2.n51 VDD2.n50 585
R1171 VDD2.n24 VDD2.n23 585
R1172 VDD2.n57 VDD2.n56 585
R1173 VDD2.n59 VDD2.n58 585
R1174 VDD2.n20 VDD2.n19 585
R1175 VDD2.n65 VDD2.n64 585
R1176 VDD2.n67 VDD2.n66 585
R1177 VDD2.n16 VDD2.n15 585
R1178 VDD2.n73 VDD2.n72 585
R1179 VDD2.n76 VDD2.n75 585
R1180 VDD2.n74 VDD2.n12 585
R1181 VDD2.n81 VDD2.n11 585
R1182 VDD2.n83 VDD2.n82 585
R1183 VDD2.n85 VDD2.n84 585
R1184 VDD2.n8 VDD2.n7 585
R1185 VDD2.n91 VDD2.n90 585
R1186 VDD2.n93 VDD2.n92 585
R1187 VDD2.n4 VDD2.n3 585
R1188 VDD2.n99 VDD2.n98 585
R1189 VDD2.n101 VDD2.n100 585
R1190 VDD2.t5 VDD2.n141 327.466
R1191 VDD2.t4 VDD2.n33 327.466
R1192 VDD2.n207 VDD2.n206 171.744
R1193 VDD2.n206 VDD2.n110 171.744
R1194 VDD2.n199 VDD2.n110 171.744
R1195 VDD2.n199 VDD2.n198 171.744
R1196 VDD2.n198 VDD2.n114 171.744
R1197 VDD2.n191 VDD2.n114 171.744
R1198 VDD2.n191 VDD2.n190 171.744
R1199 VDD2.n190 VDD2.n118 171.744
R1200 VDD2.n122 VDD2.n118 171.744
R1201 VDD2.n182 VDD2.n122 171.744
R1202 VDD2.n182 VDD2.n181 171.744
R1203 VDD2.n181 VDD2.n123 171.744
R1204 VDD2.n174 VDD2.n123 171.744
R1205 VDD2.n174 VDD2.n173 171.744
R1206 VDD2.n173 VDD2.n127 171.744
R1207 VDD2.n166 VDD2.n127 171.744
R1208 VDD2.n166 VDD2.n165 171.744
R1209 VDD2.n165 VDD2.n131 171.744
R1210 VDD2.n158 VDD2.n131 171.744
R1211 VDD2.n158 VDD2.n157 171.744
R1212 VDD2.n157 VDD2.n135 171.744
R1213 VDD2.n150 VDD2.n135 171.744
R1214 VDD2.n150 VDD2.n149 171.744
R1215 VDD2.n149 VDD2.n139 171.744
R1216 VDD2.n142 VDD2.n139 171.744
R1217 VDD2.n34 VDD2.n31 171.744
R1218 VDD2.n41 VDD2.n31 171.744
R1219 VDD2.n42 VDD2.n41 171.744
R1220 VDD2.n42 VDD2.n27 171.744
R1221 VDD2.n49 VDD2.n27 171.744
R1222 VDD2.n50 VDD2.n49 171.744
R1223 VDD2.n50 VDD2.n23 171.744
R1224 VDD2.n57 VDD2.n23 171.744
R1225 VDD2.n58 VDD2.n57 171.744
R1226 VDD2.n58 VDD2.n19 171.744
R1227 VDD2.n65 VDD2.n19 171.744
R1228 VDD2.n66 VDD2.n65 171.744
R1229 VDD2.n66 VDD2.n15 171.744
R1230 VDD2.n73 VDD2.n15 171.744
R1231 VDD2.n75 VDD2.n73 171.744
R1232 VDD2.n75 VDD2.n74 171.744
R1233 VDD2.n74 VDD2.n11 171.744
R1234 VDD2.n83 VDD2.n11 171.744
R1235 VDD2.n84 VDD2.n83 171.744
R1236 VDD2.n84 VDD2.n7 171.744
R1237 VDD2.n91 VDD2.n7 171.744
R1238 VDD2.n92 VDD2.n91 171.744
R1239 VDD2.n92 VDD2.n3 171.744
R1240 VDD2.n99 VDD2.n3 171.744
R1241 VDD2.n100 VDD2.n99 171.744
R1242 VDD2.n142 VDD2.t5 85.8723
R1243 VDD2.n34 VDD2.t4 85.8723
R1244 VDD2.n106 VDD2.n105 70.1441
R1245 VDD2 VDD2.n213 70.1411
R1246 VDD2.n106 VDD2.n104 52.313
R1247 VDD2.n212 VDD2.n106 51.086
R1248 VDD2.n212 VDD2.n211 49.8338
R1249 VDD2.n143 VDD2.n141 16.3895
R1250 VDD2.n35 VDD2.n33 16.3895
R1251 VDD2.n189 VDD2.n188 13.1884
R1252 VDD2.n82 VDD2.n81 13.1884
R1253 VDD2.n192 VDD2.n117 12.8005
R1254 VDD2.n187 VDD2.n119 12.8005
R1255 VDD2.n144 VDD2.n140 12.8005
R1256 VDD2.n36 VDD2.n32 12.8005
R1257 VDD2.n80 VDD2.n12 12.8005
R1258 VDD2.n85 VDD2.n10 12.8005
R1259 VDD2.n193 VDD2.n115 12.0247
R1260 VDD2.n184 VDD2.n183 12.0247
R1261 VDD2.n148 VDD2.n147 12.0247
R1262 VDD2.n40 VDD2.n39 12.0247
R1263 VDD2.n77 VDD2.n76 12.0247
R1264 VDD2.n86 VDD2.n8 12.0247
R1265 VDD2.n197 VDD2.n196 11.249
R1266 VDD2.n180 VDD2.n121 11.249
R1267 VDD2.n151 VDD2.n138 11.249
R1268 VDD2.n43 VDD2.n30 11.249
R1269 VDD2.n72 VDD2.n14 11.249
R1270 VDD2.n90 VDD2.n89 11.249
R1271 VDD2.n200 VDD2.n113 10.4732
R1272 VDD2.n179 VDD2.n124 10.4732
R1273 VDD2.n152 VDD2.n136 10.4732
R1274 VDD2.n44 VDD2.n28 10.4732
R1275 VDD2.n71 VDD2.n16 10.4732
R1276 VDD2.n93 VDD2.n6 10.4732
R1277 VDD2.n201 VDD2.n111 9.69747
R1278 VDD2.n176 VDD2.n175 9.69747
R1279 VDD2.n156 VDD2.n155 9.69747
R1280 VDD2.n48 VDD2.n47 9.69747
R1281 VDD2.n68 VDD2.n67 9.69747
R1282 VDD2.n94 VDD2.n4 9.69747
R1283 VDD2.n211 VDD2.n210 9.45567
R1284 VDD2.n104 VDD2.n103 9.45567
R1285 VDD2.n169 VDD2.n168 9.3005
R1286 VDD2.n171 VDD2.n170 9.3005
R1287 VDD2.n126 VDD2.n125 9.3005
R1288 VDD2.n177 VDD2.n176 9.3005
R1289 VDD2.n179 VDD2.n178 9.3005
R1290 VDD2.n121 VDD2.n120 9.3005
R1291 VDD2.n185 VDD2.n184 9.3005
R1292 VDD2.n187 VDD2.n186 9.3005
R1293 VDD2.n210 VDD2.n209 9.3005
R1294 VDD2.n109 VDD2.n108 9.3005
R1295 VDD2.n204 VDD2.n203 9.3005
R1296 VDD2.n202 VDD2.n201 9.3005
R1297 VDD2.n113 VDD2.n112 9.3005
R1298 VDD2.n196 VDD2.n195 9.3005
R1299 VDD2.n194 VDD2.n193 9.3005
R1300 VDD2.n117 VDD2.n116 9.3005
R1301 VDD2.n130 VDD2.n129 9.3005
R1302 VDD2.n163 VDD2.n162 9.3005
R1303 VDD2.n161 VDD2.n160 9.3005
R1304 VDD2.n134 VDD2.n133 9.3005
R1305 VDD2.n155 VDD2.n154 9.3005
R1306 VDD2.n153 VDD2.n152 9.3005
R1307 VDD2.n138 VDD2.n137 9.3005
R1308 VDD2.n147 VDD2.n146 9.3005
R1309 VDD2.n145 VDD2.n144 9.3005
R1310 VDD2.n2 VDD2.n1 9.3005
R1311 VDD2.n97 VDD2.n96 9.3005
R1312 VDD2.n95 VDD2.n94 9.3005
R1313 VDD2.n6 VDD2.n5 9.3005
R1314 VDD2.n89 VDD2.n88 9.3005
R1315 VDD2.n87 VDD2.n86 9.3005
R1316 VDD2.n10 VDD2.n9 9.3005
R1317 VDD2.n55 VDD2.n54 9.3005
R1318 VDD2.n53 VDD2.n52 9.3005
R1319 VDD2.n26 VDD2.n25 9.3005
R1320 VDD2.n47 VDD2.n46 9.3005
R1321 VDD2.n45 VDD2.n44 9.3005
R1322 VDD2.n30 VDD2.n29 9.3005
R1323 VDD2.n39 VDD2.n38 9.3005
R1324 VDD2.n37 VDD2.n36 9.3005
R1325 VDD2.n22 VDD2.n21 9.3005
R1326 VDD2.n61 VDD2.n60 9.3005
R1327 VDD2.n63 VDD2.n62 9.3005
R1328 VDD2.n18 VDD2.n17 9.3005
R1329 VDD2.n69 VDD2.n68 9.3005
R1330 VDD2.n71 VDD2.n70 9.3005
R1331 VDD2.n14 VDD2.n13 9.3005
R1332 VDD2.n78 VDD2.n77 9.3005
R1333 VDD2.n80 VDD2.n79 9.3005
R1334 VDD2.n103 VDD2.n102 9.3005
R1335 VDD2.n205 VDD2.n204 8.92171
R1336 VDD2.n172 VDD2.n126 8.92171
R1337 VDD2.n159 VDD2.n134 8.92171
R1338 VDD2.n51 VDD2.n26 8.92171
R1339 VDD2.n64 VDD2.n18 8.92171
R1340 VDD2.n98 VDD2.n97 8.92171
R1341 VDD2.n208 VDD2.n109 8.14595
R1342 VDD2.n171 VDD2.n128 8.14595
R1343 VDD2.n160 VDD2.n132 8.14595
R1344 VDD2.n52 VDD2.n24 8.14595
R1345 VDD2.n63 VDD2.n20 8.14595
R1346 VDD2.n101 VDD2.n2 8.14595
R1347 VDD2.n209 VDD2.n107 7.3702
R1348 VDD2.n168 VDD2.n167 7.3702
R1349 VDD2.n164 VDD2.n163 7.3702
R1350 VDD2.n56 VDD2.n55 7.3702
R1351 VDD2.n60 VDD2.n59 7.3702
R1352 VDD2.n102 VDD2.n0 7.3702
R1353 VDD2.n211 VDD2.n107 6.59444
R1354 VDD2.n167 VDD2.n130 6.59444
R1355 VDD2.n164 VDD2.n130 6.59444
R1356 VDD2.n56 VDD2.n22 6.59444
R1357 VDD2.n59 VDD2.n22 6.59444
R1358 VDD2.n104 VDD2.n0 6.59444
R1359 VDD2.n209 VDD2.n208 5.81868
R1360 VDD2.n168 VDD2.n128 5.81868
R1361 VDD2.n163 VDD2.n132 5.81868
R1362 VDD2.n55 VDD2.n24 5.81868
R1363 VDD2.n60 VDD2.n20 5.81868
R1364 VDD2.n102 VDD2.n101 5.81868
R1365 VDD2.n205 VDD2.n109 5.04292
R1366 VDD2.n172 VDD2.n171 5.04292
R1367 VDD2.n160 VDD2.n159 5.04292
R1368 VDD2.n52 VDD2.n51 5.04292
R1369 VDD2.n64 VDD2.n63 5.04292
R1370 VDD2.n98 VDD2.n2 5.04292
R1371 VDD2.n204 VDD2.n111 4.26717
R1372 VDD2.n175 VDD2.n126 4.26717
R1373 VDD2.n156 VDD2.n134 4.26717
R1374 VDD2.n48 VDD2.n26 4.26717
R1375 VDD2.n67 VDD2.n18 4.26717
R1376 VDD2.n97 VDD2.n4 4.26717
R1377 VDD2.n145 VDD2.n141 3.70982
R1378 VDD2.n37 VDD2.n33 3.70982
R1379 VDD2.n201 VDD2.n200 3.49141
R1380 VDD2.n176 VDD2.n124 3.49141
R1381 VDD2.n155 VDD2.n136 3.49141
R1382 VDD2.n47 VDD2.n28 3.49141
R1383 VDD2.n68 VDD2.n16 3.49141
R1384 VDD2.n94 VDD2.n93 3.49141
R1385 VDD2.n197 VDD2.n113 2.71565
R1386 VDD2.n180 VDD2.n179 2.71565
R1387 VDD2.n152 VDD2.n151 2.71565
R1388 VDD2.n44 VDD2.n43 2.71565
R1389 VDD2.n72 VDD2.n71 2.71565
R1390 VDD2.n90 VDD2.n6 2.71565
R1391 VDD2 VDD2.n212 2.59317
R1392 VDD2.n196 VDD2.n115 1.93989
R1393 VDD2.n183 VDD2.n121 1.93989
R1394 VDD2.n148 VDD2.n138 1.93989
R1395 VDD2.n40 VDD2.n30 1.93989
R1396 VDD2.n76 VDD2.n14 1.93989
R1397 VDD2.n89 VDD2.n8 1.93989
R1398 VDD2.n213 VDD2.t3 1.71039
R1399 VDD2.n213 VDD2.t2 1.71039
R1400 VDD2.n105 VDD2.t1 1.71039
R1401 VDD2.n105 VDD2.t0 1.71039
R1402 VDD2.n193 VDD2.n192 1.16414
R1403 VDD2.n184 VDD2.n119 1.16414
R1404 VDD2.n147 VDD2.n140 1.16414
R1405 VDD2.n39 VDD2.n32 1.16414
R1406 VDD2.n77 VDD2.n12 1.16414
R1407 VDD2.n86 VDD2.n85 1.16414
R1408 VDD2.n189 VDD2.n117 0.388379
R1409 VDD2.n188 VDD2.n187 0.388379
R1410 VDD2.n144 VDD2.n143 0.388379
R1411 VDD2.n36 VDD2.n35 0.388379
R1412 VDD2.n81 VDD2.n80 0.388379
R1413 VDD2.n82 VDD2.n10 0.388379
R1414 VDD2.n210 VDD2.n108 0.155672
R1415 VDD2.n203 VDD2.n108 0.155672
R1416 VDD2.n203 VDD2.n202 0.155672
R1417 VDD2.n202 VDD2.n112 0.155672
R1418 VDD2.n195 VDD2.n112 0.155672
R1419 VDD2.n195 VDD2.n194 0.155672
R1420 VDD2.n194 VDD2.n116 0.155672
R1421 VDD2.n186 VDD2.n116 0.155672
R1422 VDD2.n186 VDD2.n185 0.155672
R1423 VDD2.n185 VDD2.n120 0.155672
R1424 VDD2.n178 VDD2.n120 0.155672
R1425 VDD2.n178 VDD2.n177 0.155672
R1426 VDD2.n177 VDD2.n125 0.155672
R1427 VDD2.n170 VDD2.n125 0.155672
R1428 VDD2.n170 VDD2.n169 0.155672
R1429 VDD2.n169 VDD2.n129 0.155672
R1430 VDD2.n162 VDD2.n129 0.155672
R1431 VDD2.n162 VDD2.n161 0.155672
R1432 VDD2.n161 VDD2.n133 0.155672
R1433 VDD2.n154 VDD2.n133 0.155672
R1434 VDD2.n154 VDD2.n153 0.155672
R1435 VDD2.n153 VDD2.n137 0.155672
R1436 VDD2.n146 VDD2.n137 0.155672
R1437 VDD2.n146 VDD2.n145 0.155672
R1438 VDD2.n38 VDD2.n37 0.155672
R1439 VDD2.n38 VDD2.n29 0.155672
R1440 VDD2.n45 VDD2.n29 0.155672
R1441 VDD2.n46 VDD2.n45 0.155672
R1442 VDD2.n46 VDD2.n25 0.155672
R1443 VDD2.n53 VDD2.n25 0.155672
R1444 VDD2.n54 VDD2.n53 0.155672
R1445 VDD2.n54 VDD2.n21 0.155672
R1446 VDD2.n61 VDD2.n21 0.155672
R1447 VDD2.n62 VDD2.n61 0.155672
R1448 VDD2.n62 VDD2.n17 0.155672
R1449 VDD2.n69 VDD2.n17 0.155672
R1450 VDD2.n70 VDD2.n69 0.155672
R1451 VDD2.n70 VDD2.n13 0.155672
R1452 VDD2.n78 VDD2.n13 0.155672
R1453 VDD2.n79 VDD2.n78 0.155672
R1454 VDD2.n79 VDD2.n9 0.155672
R1455 VDD2.n87 VDD2.n9 0.155672
R1456 VDD2.n88 VDD2.n87 0.155672
R1457 VDD2.n88 VDD2.n5 0.155672
R1458 VDD2.n95 VDD2.n5 0.155672
R1459 VDD2.n96 VDD2.n95 0.155672
R1460 VDD2.n96 VDD2.n1 0.155672
R1461 VDD2.n103 VDD2.n1 0.155672
R1462 B.n699 B.n100 585
R1463 B.n701 B.n700 585
R1464 B.n702 B.n99 585
R1465 B.n704 B.n703 585
R1466 B.n705 B.n98 585
R1467 B.n707 B.n706 585
R1468 B.n708 B.n97 585
R1469 B.n710 B.n709 585
R1470 B.n711 B.n96 585
R1471 B.n713 B.n712 585
R1472 B.n714 B.n95 585
R1473 B.n716 B.n715 585
R1474 B.n717 B.n94 585
R1475 B.n719 B.n718 585
R1476 B.n720 B.n93 585
R1477 B.n722 B.n721 585
R1478 B.n723 B.n92 585
R1479 B.n725 B.n724 585
R1480 B.n726 B.n91 585
R1481 B.n728 B.n727 585
R1482 B.n729 B.n90 585
R1483 B.n731 B.n730 585
R1484 B.n732 B.n89 585
R1485 B.n734 B.n733 585
R1486 B.n735 B.n88 585
R1487 B.n737 B.n736 585
R1488 B.n738 B.n87 585
R1489 B.n740 B.n739 585
R1490 B.n741 B.n86 585
R1491 B.n743 B.n742 585
R1492 B.n744 B.n85 585
R1493 B.n746 B.n745 585
R1494 B.n747 B.n84 585
R1495 B.n749 B.n748 585
R1496 B.n750 B.n83 585
R1497 B.n752 B.n751 585
R1498 B.n753 B.n82 585
R1499 B.n755 B.n754 585
R1500 B.n756 B.n81 585
R1501 B.n758 B.n757 585
R1502 B.n759 B.n80 585
R1503 B.n761 B.n760 585
R1504 B.n762 B.n79 585
R1505 B.n764 B.n763 585
R1506 B.n765 B.n78 585
R1507 B.n767 B.n766 585
R1508 B.n768 B.n77 585
R1509 B.n770 B.n769 585
R1510 B.n771 B.n76 585
R1511 B.n773 B.n772 585
R1512 B.n774 B.n75 585
R1513 B.n776 B.n775 585
R1514 B.n777 B.n74 585
R1515 B.n779 B.n778 585
R1516 B.n780 B.n73 585
R1517 B.n782 B.n781 585
R1518 B.n783 B.n72 585
R1519 B.n785 B.n784 585
R1520 B.n786 B.n71 585
R1521 B.n788 B.n787 585
R1522 B.n789 B.n70 585
R1523 B.n791 B.n790 585
R1524 B.n793 B.n67 585
R1525 B.n795 B.n794 585
R1526 B.n796 B.n66 585
R1527 B.n798 B.n797 585
R1528 B.n799 B.n65 585
R1529 B.n801 B.n800 585
R1530 B.n802 B.n64 585
R1531 B.n804 B.n803 585
R1532 B.n805 B.n63 585
R1533 B.n807 B.n806 585
R1534 B.n809 B.n808 585
R1535 B.n810 B.n59 585
R1536 B.n812 B.n811 585
R1537 B.n813 B.n58 585
R1538 B.n815 B.n814 585
R1539 B.n816 B.n57 585
R1540 B.n818 B.n817 585
R1541 B.n819 B.n56 585
R1542 B.n821 B.n820 585
R1543 B.n822 B.n55 585
R1544 B.n824 B.n823 585
R1545 B.n825 B.n54 585
R1546 B.n827 B.n826 585
R1547 B.n828 B.n53 585
R1548 B.n830 B.n829 585
R1549 B.n831 B.n52 585
R1550 B.n833 B.n832 585
R1551 B.n834 B.n51 585
R1552 B.n836 B.n835 585
R1553 B.n837 B.n50 585
R1554 B.n839 B.n838 585
R1555 B.n840 B.n49 585
R1556 B.n842 B.n841 585
R1557 B.n843 B.n48 585
R1558 B.n845 B.n844 585
R1559 B.n846 B.n47 585
R1560 B.n848 B.n847 585
R1561 B.n849 B.n46 585
R1562 B.n851 B.n850 585
R1563 B.n852 B.n45 585
R1564 B.n854 B.n853 585
R1565 B.n855 B.n44 585
R1566 B.n857 B.n856 585
R1567 B.n858 B.n43 585
R1568 B.n860 B.n859 585
R1569 B.n861 B.n42 585
R1570 B.n863 B.n862 585
R1571 B.n864 B.n41 585
R1572 B.n866 B.n865 585
R1573 B.n867 B.n40 585
R1574 B.n869 B.n868 585
R1575 B.n870 B.n39 585
R1576 B.n872 B.n871 585
R1577 B.n873 B.n38 585
R1578 B.n875 B.n874 585
R1579 B.n876 B.n37 585
R1580 B.n878 B.n877 585
R1581 B.n879 B.n36 585
R1582 B.n881 B.n880 585
R1583 B.n882 B.n35 585
R1584 B.n884 B.n883 585
R1585 B.n885 B.n34 585
R1586 B.n887 B.n886 585
R1587 B.n888 B.n33 585
R1588 B.n890 B.n889 585
R1589 B.n891 B.n32 585
R1590 B.n893 B.n892 585
R1591 B.n894 B.n31 585
R1592 B.n896 B.n895 585
R1593 B.n897 B.n30 585
R1594 B.n899 B.n898 585
R1595 B.n900 B.n29 585
R1596 B.n698 B.n697 585
R1597 B.n696 B.n101 585
R1598 B.n695 B.n694 585
R1599 B.n693 B.n102 585
R1600 B.n692 B.n691 585
R1601 B.n690 B.n103 585
R1602 B.n689 B.n688 585
R1603 B.n687 B.n104 585
R1604 B.n686 B.n685 585
R1605 B.n684 B.n105 585
R1606 B.n683 B.n682 585
R1607 B.n681 B.n106 585
R1608 B.n680 B.n679 585
R1609 B.n678 B.n107 585
R1610 B.n677 B.n676 585
R1611 B.n675 B.n108 585
R1612 B.n674 B.n673 585
R1613 B.n672 B.n109 585
R1614 B.n671 B.n670 585
R1615 B.n669 B.n110 585
R1616 B.n668 B.n667 585
R1617 B.n666 B.n111 585
R1618 B.n665 B.n664 585
R1619 B.n663 B.n112 585
R1620 B.n662 B.n661 585
R1621 B.n660 B.n113 585
R1622 B.n659 B.n658 585
R1623 B.n657 B.n114 585
R1624 B.n656 B.n655 585
R1625 B.n654 B.n115 585
R1626 B.n653 B.n652 585
R1627 B.n651 B.n116 585
R1628 B.n650 B.n649 585
R1629 B.n648 B.n117 585
R1630 B.n647 B.n646 585
R1631 B.n645 B.n118 585
R1632 B.n644 B.n643 585
R1633 B.n642 B.n119 585
R1634 B.n641 B.n640 585
R1635 B.n639 B.n120 585
R1636 B.n638 B.n637 585
R1637 B.n636 B.n121 585
R1638 B.n635 B.n634 585
R1639 B.n633 B.n122 585
R1640 B.n632 B.n631 585
R1641 B.n630 B.n123 585
R1642 B.n629 B.n628 585
R1643 B.n627 B.n124 585
R1644 B.n626 B.n625 585
R1645 B.n624 B.n125 585
R1646 B.n623 B.n622 585
R1647 B.n621 B.n126 585
R1648 B.n620 B.n619 585
R1649 B.n618 B.n127 585
R1650 B.n617 B.n616 585
R1651 B.n615 B.n128 585
R1652 B.n614 B.n613 585
R1653 B.n612 B.n129 585
R1654 B.n611 B.n610 585
R1655 B.n609 B.n130 585
R1656 B.n608 B.n607 585
R1657 B.n606 B.n131 585
R1658 B.n605 B.n604 585
R1659 B.n603 B.n132 585
R1660 B.n602 B.n601 585
R1661 B.n600 B.n133 585
R1662 B.n599 B.n598 585
R1663 B.n597 B.n134 585
R1664 B.n596 B.n595 585
R1665 B.n594 B.n135 585
R1666 B.n593 B.n592 585
R1667 B.n591 B.n136 585
R1668 B.n590 B.n589 585
R1669 B.n588 B.n137 585
R1670 B.n587 B.n586 585
R1671 B.n585 B.n138 585
R1672 B.n584 B.n583 585
R1673 B.n582 B.n139 585
R1674 B.n581 B.n580 585
R1675 B.n579 B.n140 585
R1676 B.n578 B.n577 585
R1677 B.n576 B.n141 585
R1678 B.n575 B.n574 585
R1679 B.n573 B.n142 585
R1680 B.n572 B.n571 585
R1681 B.n570 B.n143 585
R1682 B.n569 B.n568 585
R1683 B.n567 B.n144 585
R1684 B.n566 B.n565 585
R1685 B.n564 B.n145 585
R1686 B.n563 B.n562 585
R1687 B.n561 B.n146 585
R1688 B.n560 B.n559 585
R1689 B.n558 B.n147 585
R1690 B.n557 B.n556 585
R1691 B.n555 B.n148 585
R1692 B.n554 B.n553 585
R1693 B.n552 B.n149 585
R1694 B.n551 B.n550 585
R1695 B.n549 B.n150 585
R1696 B.n548 B.n547 585
R1697 B.n546 B.n151 585
R1698 B.n545 B.n544 585
R1699 B.n543 B.n152 585
R1700 B.n542 B.n541 585
R1701 B.n540 B.n153 585
R1702 B.n539 B.n538 585
R1703 B.n537 B.n154 585
R1704 B.n536 B.n535 585
R1705 B.n333 B.n226 585
R1706 B.n335 B.n334 585
R1707 B.n336 B.n225 585
R1708 B.n338 B.n337 585
R1709 B.n339 B.n224 585
R1710 B.n341 B.n340 585
R1711 B.n342 B.n223 585
R1712 B.n344 B.n343 585
R1713 B.n345 B.n222 585
R1714 B.n347 B.n346 585
R1715 B.n348 B.n221 585
R1716 B.n350 B.n349 585
R1717 B.n351 B.n220 585
R1718 B.n353 B.n352 585
R1719 B.n354 B.n219 585
R1720 B.n356 B.n355 585
R1721 B.n357 B.n218 585
R1722 B.n359 B.n358 585
R1723 B.n360 B.n217 585
R1724 B.n362 B.n361 585
R1725 B.n363 B.n216 585
R1726 B.n365 B.n364 585
R1727 B.n366 B.n215 585
R1728 B.n368 B.n367 585
R1729 B.n369 B.n214 585
R1730 B.n371 B.n370 585
R1731 B.n372 B.n213 585
R1732 B.n374 B.n373 585
R1733 B.n375 B.n212 585
R1734 B.n377 B.n376 585
R1735 B.n378 B.n211 585
R1736 B.n380 B.n379 585
R1737 B.n381 B.n210 585
R1738 B.n383 B.n382 585
R1739 B.n384 B.n209 585
R1740 B.n386 B.n385 585
R1741 B.n387 B.n208 585
R1742 B.n389 B.n388 585
R1743 B.n390 B.n207 585
R1744 B.n392 B.n391 585
R1745 B.n393 B.n206 585
R1746 B.n395 B.n394 585
R1747 B.n396 B.n205 585
R1748 B.n398 B.n397 585
R1749 B.n399 B.n204 585
R1750 B.n401 B.n400 585
R1751 B.n402 B.n203 585
R1752 B.n404 B.n403 585
R1753 B.n405 B.n202 585
R1754 B.n407 B.n406 585
R1755 B.n408 B.n201 585
R1756 B.n410 B.n409 585
R1757 B.n411 B.n200 585
R1758 B.n413 B.n412 585
R1759 B.n414 B.n199 585
R1760 B.n416 B.n415 585
R1761 B.n417 B.n198 585
R1762 B.n419 B.n418 585
R1763 B.n420 B.n197 585
R1764 B.n422 B.n421 585
R1765 B.n423 B.n196 585
R1766 B.n425 B.n424 585
R1767 B.n427 B.n193 585
R1768 B.n429 B.n428 585
R1769 B.n430 B.n192 585
R1770 B.n432 B.n431 585
R1771 B.n433 B.n191 585
R1772 B.n435 B.n434 585
R1773 B.n436 B.n190 585
R1774 B.n438 B.n437 585
R1775 B.n439 B.n189 585
R1776 B.n441 B.n440 585
R1777 B.n443 B.n442 585
R1778 B.n444 B.n185 585
R1779 B.n446 B.n445 585
R1780 B.n447 B.n184 585
R1781 B.n449 B.n448 585
R1782 B.n450 B.n183 585
R1783 B.n452 B.n451 585
R1784 B.n453 B.n182 585
R1785 B.n455 B.n454 585
R1786 B.n456 B.n181 585
R1787 B.n458 B.n457 585
R1788 B.n459 B.n180 585
R1789 B.n461 B.n460 585
R1790 B.n462 B.n179 585
R1791 B.n464 B.n463 585
R1792 B.n465 B.n178 585
R1793 B.n467 B.n466 585
R1794 B.n468 B.n177 585
R1795 B.n470 B.n469 585
R1796 B.n471 B.n176 585
R1797 B.n473 B.n472 585
R1798 B.n474 B.n175 585
R1799 B.n476 B.n475 585
R1800 B.n477 B.n174 585
R1801 B.n479 B.n478 585
R1802 B.n480 B.n173 585
R1803 B.n482 B.n481 585
R1804 B.n483 B.n172 585
R1805 B.n485 B.n484 585
R1806 B.n486 B.n171 585
R1807 B.n488 B.n487 585
R1808 B.n489 B.n170 585
R1809 B.n491 B.n490 585
R1810 B.n492 B.n169 585
R1811 B.n494 B.n493 585
R1812 B.n495 B.n168 585
R1813 B.n497 B.n496 585
R1814 B.n498 B.n167 585
R1815 B.n500 B.n499 585
R1816 B.n501 B.n166 585
R1817 B.n503 B.n502 585
R1818 B.n504 B.n165 585
R1819 B.n506 B.n505 585
R1820 B.n507 B.n164 585
R1821 B.n509 B.n508 585
R1822 B.n510 B.n163 585
R1823 B.n512 B.n511 585
R1824 B.n513 B.n162 585
R1825 B.n515 B.n514 585
R1826 B.n516 B.n161 585
R1827 B.n518 B.n517 585
R1828 B.n519 B.n160 585
R1829 B.n521 B.n520 585
R1830 B.n522 B.n159 585
R1831 B.n524 B.n523 585
R1832 B.n525 B.n158 585
R1833 B.n527 B.n526 585
R1834 B.n528 B.n157 585
R1835 B.n530 B.n529 585
R1836 B.n531 B.n156 585
R1837 B.n533 B.n532 585
R1838 B.n534 B.n155 585
R1839 B.n332 B.n331 585
R1840 B.n330 B.n227 585
R1841 B.n329 B.n328 585
R1842 B.n327 B.n228 585
R1843 B.n326 B.n325 585
R1844 B.n324 B.n229 585
R1845 B.n323 B.n322 585
R1846 B.n321 B.n230 585
R1847 B.n320 B.n319 585
R1848 B.n318 B.n231 585
R1849 B.n317 B.n316 585
R1850 B.n315 B.n232 585
R1851 B.n314 B.n313 585
R1852 B.n312 B.n233 585
R1853 B.n311 B.n310 585
R1854 B.n309 B.n234 585
R1855 B.n308 B.n307 585
R1856 B.n306 B.n235 585
R1857 B.n305 B.n304 585
R1858 B.n303 B.n236 585
R1859 B.n302 B.n301 585
R1860 B.n300 B.n237 585
R1861 B.n299 B.n298 585
R1862 B.n297 B.n238 585
R1863 B.n296 B.n295 585
R1864 B.n294 B.n239 585
R1865 B.n293 B.n292 585
R1866 B.n291 B.n240 585
R1867 B.n290 B.n289 585
R1868 B.n288 B.n241 585
R1869 B.n287 B.n286 585
R1870 B.n285 B.n242 585
R1871 B.n284 B.n283 585
R1872 B.n282 B.n243 585
R1873 B.n281 B.n280 585
R1874 B.n279 B.n244 585
R1875 B.n278 B.n277 585
R1876 B.n276 B.n245 585
R1877 B.n275 B.n274 585
R1878 B.n273 B.n246 585
R1879 B.n272 B.n271 585
R1880 B.n270 B.n247 585
R1881 B.n269 B.n268 585
R1882 B.n267 B.n248 585
R1883 B.n266 B.n265 585
R1884 B.n264 B.n249 585
R1885 B.n263 B.n262 585
R1886 B.n261 B.n250 585
R1887 B.n260 B.n259 585
R1888 B.n258 B.n251 585
R1889 B.n257 B.n256 585
R1890 B.n255 B.n252 585
R1891 B.n254 B.n253 585
R1892 B.n2 B.n0 585
R1893 B.n981 B.n1 585
R1894 B.n980 B.n979 585
R1895 B.n978 B.n3 585
R1896 B.n977 B.n976 585
R1897 B.n975 B.n4 585
R1898 B.n974 B.n973 585
R1899 B.n972 B.n5 585
R1900 B.n971 B.n970 585
R1901 B.n969 B.n6 585
R1902 B.n968 B.n967 585
R1903 B.n966 B.n7 585
R1904 B.n965 B.n964 585
R1905 B.n963 B.n8 585
R1906 B.n962 B.n961 585
R1907 B.n960 B.n9 585
R1908 B.n959 B.n958 585
R1909 B.n957 B.n10 585
R1910 B.n956 B.n955 585
R1911 B.n954 B.n11 585
R1912 B.n953 B.n952 585
R1913 B.n951 B.n12 585
R1914 B.n950 B.n949 585
R1915 B.n948 B.n13 585
R1916 B.n947 B.n946 585
R1917 B.n945 B.n14 585
R1918 B.n944 B.n943 585
R1919 B.n942 B.n15 585
R1920 B.n941 B.n940 585
R1921 B.n939 B.n16 585
R1922 B.n938 B.n937 585
R1923 B.n936 B.n17 585
R1924 B.n935 B.n934 585
R1925 B.n933 B.n18 585
R1926 B.n932 B.n931 585
R1927 B.n930 B.n19 585
R1928 B.n929 B.n928 585
R1929 B.n927 B.n20 585
R1930 B.n926 B.n925 585
R1931 B.n924 B.n21 585
R1932 B.n923 B.n922 585
R1933 B.n921 B.n22 585
R1934 B.n920 B.n919 585
R1935 B.n918 B.n23 585
R1936 B.n917 B.n916 585
R1937 B.n915 B.n24 585
R1938 B.n914 B.n913 585
R1939 B.n912 B.n25 585
R1940 B.n911 B.n910 585
R1941 B.n909 B.n26 585
R1942 B.n908 B.n907 585
R1943 B.n906 B.n27 585
R1944 B.n905 B.n904 585
R1945 B.n903 B.n28 585
R1946 B.n902 B.n901 585
R1947 B.n983 B.n982 585
R1948 B.n186 B.t11 578.106
R1949 B.n68 B.t4 578.106
R1950 B.n194 B.t8 578.106
R1951 B.n60 B.t1 578.106
R1952 B.n333 B.n332 540.549
R1953 B.n902 B.n29 540.549
R1954 B.n536 B.n155 540.549
R1955 B.n699 B.n698 540.549
R1956 B.n187 B.t10 502.082
R1957 B.n69 B.t5 502.082
R1958 B.n195 B.t7 502.082
R1959 B.n61 B.t2 502.082
R1960 B.n186 B.t9 336.788
R1961 B.n194 B.t6 336.788
R1962 B.n60 B.t0 336.788
R1963 B.n68 B.t3 336.788
R1964 B.n332 B.n227 163.367
R1965 B.n328 B.n227 163.367
R1966 B.n328 B.n327 163.367
R1967 B.n327 B.n326 163.367
R1968 B.n326 B.n229 163.367
R1969 B.n322 B.n229 163.367
R1970 B.n322 B.n321 163.367
R1971 B.n321 B.n320 163.367
R1972 B.n320 B.n231 163.367
R1973 B.n316 B.n231 163.367
R1974 B.n316 B.n315 163.367
R1975 B.n315 B.n314 163.367
R1976 B.n314 B.n233 163.367
R1977 B.n310 B.n233 163.367
R1978 B.n310 B.n309 163.367
R1979 B.n309 B.n308 163.367
R1980 B.n308 B.n235 163.367
R1981 B.n304 B.n235 163.367
R1982 B.n304 B.n303 163.367
R1983 B.n303 B.n302 163.367
R1984 B.n302 B.n237 163.367
R1985 B.n298 B.n237 163.367
R1986 B.n298 B.n297 163.367
R1987 B.n297 B.n296 163.367
R1988 B.n296 B.n239 163.367
R1989 B.n292 B.n239 163.367
R1990 B.n292 B.n291 163.367
R1991 B.n291 B.n290 163.367
R1992 B.n290 B.n241 163.367
R1993 B.n286 B.n241 163.367
R1994 B.n286 B.n285 163.367
R1995 B.n285 B.n284 163.367
R1996 B.n284 B.n243 163.367
R1997 B.n280 B.n243 163.367
R1998 B.n280 B.n279 163.367
R1999 B.n279 B.n278 163.367
R2000 B.n278 B.n245 163.367
R2001 B.n274 B.n245 163.367
R2002 B.n274 B.n273 163.367
R2003 B.n273 B.n272 163.367
R2004 B.n272 B.n247 163.367
R2005 B.n268 B.n247 163.367
R2006 B.n268 B.n267 163.367
R2007 B.n267 B.n266 163.367
R2008 B.n266 B.n249 163.367
R2009 B.n262 B.n249 163.367
R2010 B.n262 B.n261 163.367
R2011 B.n261 B.n260 163.367
R2012 B.n260 B.n251 163.367
R2013 B.n256 B.n251 163.367
R2014 B.n256 B.n255 163.367
R2015 B.n255 B.n254 163.367
R2016 B.n254 B.n2 163.367
R2017 B.n982 B.n2 163.367
R2018 B.n982 B.n981 163.367
R2019 B.n981 B.n980 163.367
R2020 B.n980 B.n3 163.367
R2021 B.n976 B.n3 163.367
R2022 B.n976 B.n975 163.367
R2023 B.n975 B.n974 163.367
R2024 B.n974 B.n5 163.367
R2025 B.n970 B.n5 163.367
R2026 B.n970 B.n969 163.367
R2027 B.n969 B.n968 163.367
R2028 B.n968 B.n7 163.367
R2029 B.n964 B.n7 163.367
R2030 B.n964 B.n963 163.367
R2031 B.n963 B.n962 163.367
R2032 B.n962 B.n9 163.367
R2033 B.n958 B.n9 163.367
R2034 B.n958 B.n957 163.367
R2035 B.n957 B.n956 163.367
R2036 B.n956 B.n11 163.367
R2037 B.n952 B.n11 163.367
R2038 B.n952 B.n951 163.367
R2039 B.n951 B.n950 163.367
R2040 B.n950 B.n13 163.367
R2041 B.n946 B.n13 163.367
R2042 B.n946 B.n945 163.367
R2043 B.n945 B.n944 163.367
R2044 B.n944 B.n15 163.367
R2045 B.n940 B.n15 163.367
R2046 B.n940 B.n939 163.367
R2047 B.n939 B.n938 163.367
R2048 B.n938 B.n17 163.367
R2049 B.n934 B.n17 163.367
R2050 B.n934 B.n933 163.367
R2051 B.n933 B.n932 163.367
R2052 B.n932 B.n19 163.367
R2053 B.n928 B.n19 163.367
R2054 B.n928 B.n927 163.367
R2055 B.n927 B.n926 163.367
R2056 B.n926 B.n21 163.367
R2057 B.n922 B.n21 163.367
R2058 B.n922 B.n921 163.367
R2059 B.n921 B.n920 163.367
R2060 B.n920 B.n23 163.367
R2061 B.n916 B.n23 163.367
R2062 B.n916 B.n915 163.367
R2063 B.n915 B.n914 163.367
R2064 B.n914 B.n25 163.367
R2065 B.n910 B.n25 163.367
R2066 B.n910 B.n909 163.367
R2067 B.n909 B.n908 163.367
R2068 B.n908 B.n27 163.367
R2069 B.n904 B.n27 163.367
R2070 B.n904 B.n903 163.367
R2071 B.n903 B.n902 163.367
R2072 B.n334 B.n333 163.367
R2073 B.n334 B.n225 163.367
R2074 B.n338 B.n225 163.367
R2075 B.n339 B.n338 163.367
R2076 B.n340 B.n339 163.367
R2077 B.n340 B.n223 163.367
R2078 B.n344 B.n223 163.367
R2079 B.n345 B.n344 163.367
R2080 B.n346 B.n345 163.367
R2081 B.n346 B.n221 163.367
R2082 B.n350 B.n221 163.367
R2083 B.n351 B.n350 163.367
R2084 B.n352 B.n351 163.367
R2085 B.n352 B.n219 163.367
R2086 B.n356 B.n219 163.367
R2087 B.n357 B.n356 163.367
R2088 B.n358 B.n357 163.367
R2089 B.n358 B.n217 163.367
R2090 B.n362 B.n217 163.367
R2091 B.n363 B.n362 163.367
R2092 B.n364 B.n363 163.367
R2093 B.n364 B.n215 163.367
R2094 B.n368 B.n215 163.367
R2095 B.n369 B.n368 163.367
R2096 B.n370 B.n369 163.367
R2097 B.n370 B.n213 163.367
R2098 B.n374 B.n213 163.367
R2099 B.n375 B.n374 163.367
R2100 B.n376 B.n375 163.367
R2101 B.n376 B.n211 163.367
R2102 B.n380 B.n211 163.367
R2103 B.n381 B.n380 163.367
R2104 B.n382 B.n381 163.367
R2105 B.n382 B.n209 163.367
R2106 B.n386 B.n209 163.367
R2107 B.n387 B.n386 163.367
R2108 B.n388 B.n387 163.367
R2109 B.n388 B.n207 163.367
R2110 B.n392 B.n207 163.367
R2111 B.n393 B.n392 163.367
R2112 B.n394 B.n393 163.367
R2113 B.n394 B.n205 163.367
R2114 B.n398 B.n205 163.367
R2115 B.n399 B.n398 163.367
R2116 B.n400 B.n399 163.367
R2117 B.n400 B.n203 163.367
R2118 B.n404 B.n203 163.367
R2119 B.n405 B.n404 163.367
R2120 B.n406 B.n405 163.367
R2121 B.n406 B.n201 163.367
R2122 B.n410 B.n201 163.367
R2123 B.n411 B.n410 163.367
R2124 B.n412 B.n411 163.367
R2125 B.n412 B.n199 163.367
R2126 B.n416 B.n199 163.367
R2127 B.n417 B.n416 163.367
R2128 B.n418 B.n417 163.367
R2129 B.n418 B.n197 163.367
R2130 B.n422 B.n197 163.367
R2131 B.n423 B.n422 163.367
R2132 B.n424 B.n423 163.367
R2133 B.n424 B.n193 163.367
R2134 B.n429 B.n193 163.367
R2135 B.n430 B.n429 163.367
R2136 B.n431 B.n430 163.367
R2137 B.n431 B.n191 163.367
R2138 B.n435 B.n191 163.367
R2139 B.n436 B.n435 163.367
R2140 B.n437 B.n436 163.367
R2141 B.n437 B.n189 163.367
R2142 B.n441 B.n189 163.367
R2143 B.n442 B.n441 163.367
R2144 B.n442 B.n185 163.367
R2145 B.n446 B.n185 163.367
R2146 B.n447 B.n446 163.367
R2147 B.n448 B.n447 163.367
R2148 B.n448 B.n183 163.367
R2149 B.n452 B.n183 163.367
R2150 B.n453 B.n452 163.367
R2151 B.n454 B.n453 163.367
R2152 B.n454 B.n181 163.367
R2153 B.n458 B.n181 163.367
R2154 B.n459 B.n458 163.367
R2155 B.n460 B.n459 163.367
R2156 B.n460 B.n179 163.367
R2157 B.n464 B.n179 163.367
R2158 B.n465 B.n464 163.367
R2159 B.n466 B.n465 163.367
R2160 B.n466 B.n177 163.367
R2161 B.n470 B.n177 163.367
R2162 B.n471 B.n470 163.367
R2163 B.n472 B.n471 163.367
R2164 B.n472 B.n175 163.367
R2165 B.n476 B.n175 163.367
R2166 B.n477 B.n476 163.367
R2167 B.n478 B.n477 163.367
R2168 B.n478 B.n173 163.367
R2169 B.n482 B.n173 163.367
R2170 B.n483 B.n482 163.367
R2171 B.n484 B.n483 163.367
R2172 B.n484 B.n171 163.367
R2173 B.n488 B.n171 163.367
R2174 B.n489 B.n488 163.367
R2175 B.n490 B.n489 163.367
R2176 B.n490 B.n169 163.367
R2177 B.n494 B.n169 163.367
R2178 B.n495 B.n494 163.367
R2179 B.n496 B.n495 163.367
R2180 B.n496 B.n167 163.367
R2181 B.n500 B.n167 163.367
R2182 B.n501 B.n500 163.367
R2183 B.n502 B.n501 163.367
R2184 B.n502 B.n165 163.367
R2185 B.n506 B.n165 163.367
R2186 B.n507 B.n506 163.367
R2187 B.n508 B.n507 163.367
R2188 B.n508 B.n163 163.367
R2189 B.n512 B.n163 163.367
R2190 B.n513 B.n512 163.367
R2191 B.n514 B.n513 163.367
R2192 B.n514 B.n161 163.367
R2193 B.n518 B.n161 163.367
R2194 B.n519 B.n518 163.367
R2195 B.n520 B.n519 163.367
R2196 B.n520 B.n159 163.367
R2197 B.n524 B.n159 163.367
R2198 B.n525 B.n524 163.367
R2199 B.n526 B.n525 163.367
R2200 B.n526 B.n157 163.367
R2201 B.n530 B.n157 163.367
R2202 B.n531 B.n530 163.367
R2203 B.n532 B.n531 163.367
R2204 B.n532 B.n155 163.367
R2205 B.n537 B.n536 163.367
R2206 B.n538 B.n537 163.367
R2207 B.n538 B.n153 163.367
R2208 B.n542 B.n153 163.367
R2209 B.n543 B.n542 163.367
R2210 B.n544 B.n543 163.367
R2211 B.n544 B.n151 163.367
R2212 B.n548 B.n151 163.367
R2213 B.n549 B.n548 163.367
R2214 B.n550 B.n549 163.367
R2215 B.n550 B.n149 163.367
R2216 B.n554 B.n149 163.367
R2217 B.n555 B.n554 163.367
R2218 B.n556 B.n555 163.367
R2219 B.n556 B.n147 163.367
R2220 B.n560 B.n147 163.367
R2221 B.n561 B.n560 163.367
R2222 B.n562 B.n561 163.367
R2223 B.n562 B.n145 163.367
R2224 B.n566 B.n145 163.367
R2225 B.n567 B.n566 163.367
R2226 B.n568 B.n567 163.367
R2227 B.n568 B.n143 163.367
R2228 B.n572 B.n143 163.367
R2229 B.n573 B.n572 163.367
R2230 B.n574 B.n573 163.367
R2231 B.n574 B.n141 163.367
R2232 B.n578 B.n141 163.367
R2233 B.n579 B.n578 163.367
R2234 B.n580 B.n579 163.367
R2235 B.n580 B.n139 163.367
R2236 B.n584 B.n139 163.367
R2237 B.n585 B.n584 163.367
R2238 B.n586 B.n585 163.367
R2239 B.n586 B.n137 163.367
R2240 B.n590 B.n137 163.367
R2241 B.n591 B.n590 163.367
R2242 B.n592 B.n591 163.367
R2243 B.n592 B.n135 163.367
R2244 B.n596 B.n135 163.367
R2245 B.n597 B.n596 163.367
R2246 B.n598 B.n597 163.367
R2247 B.n598 B.n133 163.367
R2248 B.n602 B.n133 163.367
R2249 B.n603 B.n602 163.367
R2250 B.n604 B.n603 163.367
R2251 B.n604 B.n131 163.367
R2252 B.n608 B.n131 163.367
R2253 B.n609 B.n608 163.367
R2254 B.n610 B.n609 163.367
R2255 B.n610 B.n129 163.367
R2256 B.n614 B.n129 163.367
R2257 B.n615 B.n614 163.367
R2258 B.n616 B.n615 163.367
R2259 B.n616 B.n127 163.367
R2260 B.n620 B.n127 163.367
R2261 B.n621 B.n620 163.367
R2262 B.n622 B.n621 163.367
R2263 B.n622 B.n125 163.367
R2264 B.n626 B.n125 163.367
R2265 B.n627 B.n626 163.367
R2266 B.n628 B.n627 163.367
R2267 B.n628 B.n123 163.367
R2268 B.n632 B.n123 163.367
R2269 B.n633 B.n632 163.367
R2270 B.n634 B.n633 163.367
R2271 B.n634 B.n121 163.367
R2272 B.n638 B.n121 163.367
R2273 B.n639 B.n638 163.367
R2274 B.n640 B.n639 163.367
R2275 B.n640 B.n119 163.367
R2276 B.n644 B.n119 163.367
R2277 B.n645 B.n644 163.367
R2278 B.n646 B.n645 163.367
R2279 B.n646 B.n117 163.367
R2280 B.n650 B.n117 163.367
R2281 B.n651 B.n650 163.367
R2282 B.n652 B.n651 163.367
R2283 B.n652 B.n115 163.367
R2284 B.n656 B.n115 163.367
R2285 B.n657 B.n656 163.367
R2286 B.n658 B.n657 163.367
R2287 B.n658 B.n113 163.367
R2288 B.n662 B.n113 163.367
R2289 B.n663 B.n662 163.367
R2290 B.n664 B.n663 163.367
R2291 B.n664 B.n111 163.367
R2292 B.n668 B.n111 163.367
R2293 B.n669 B.n668 163.367
R2294 B.n670 B.n669 163.367
R2295 B.n670 B.n109 163.367
R2296 B.n674 B.n109 163.367
R2297 B.n675 B.n674 163.367
R2298 B.n676 B.n675 163.367
R2299 B.n676 B.n107 163.367
R2300 B.n680 B.n107 163.367
R2301 B.n681 B.n680 163.367
R2302 B.n682 B.n681 163.367
R2303 B.n682 B.n105 163.367
R2304 B.n686 B.n105 163.367
R2305 B.n687 B.n686 163.367
R2306 B.n688 B.n687 163.367
R2307 B.n688 B.n103 163.367
R2308 B.n692 B.n103 163.367
R2309 B.n693 B.n692 163.367
R2310 B.n694 B.n693 163.367
R2311 B.n694 B.n101 163.367
R2312 B.n698 B.n101 163.367
R2313 B.n898 B.n29 163.367
R2314 B.n898 B.n897 163.367
R2315 B.n897 B.n896 163.367
R2316 B.n896 B.n31 163.367
R2317 B.n892 B.n31 163.367
R2318 B.n892 B.n891 163.367
R2319 B.n891 B.n890 163.367
R2320 B.n890 B.n33 163.367
R2321 B.n886 B.n33 163.367
R2322 B.n886 B.n885 163.367
R2323 B.n885 B.n884 163.367
R2324 B.n884 B.n35 163.367
R2325 B.n880 B.n35 163.367
R2326 B.n880 B.n879 163.367
R2327 B.n879 B.n878 163.367
R2328 B.n878 B.n37 163.367
R2329 B.n874 B.n37 163.367
R2330 B.n874 B.n873 163.367
R2331 B.n873 B.n872 163.367
R2332 B.n872 B.n39 163.367
R2333 B.n868 B.n39 163.367
R2334 B.n868 B.n867 163.367
R2335 B.n867 B.n866 163.367
R2336 B.n866 B.n41 163.367
R2337 B.n862 B.n41 163.367
R2338 B.n862 B.n861 163.367
R2339 B.n861 B.n860 163.367
R2340 B.n860 B.n43 163.367
R2341 B.n856 B.n43 163.367
R2342 B.n856 B.n855 163.367
R2343 B.n855 B.n854 163.367
R2344 B.n854 B.n45 163.367
R2345 B.n850 B.n45 163.367
R2346 B.n850 B.n849 163.367
R2347 B.n849 B.n848 163.367
R2348 B.n848 B.n47 163.367
R2349 B.n844 B.n47 163.367
R2350 B.n844 B.n843 163.367
R2351 B.n843 B.n842 163.367
R2352 B.n842 B.n49 163.367
R2353 B.n838 B.n49 163.367
R2354 B.n838 B.n837 163.367
R2355 B.n837 B.n836 163.367
R2356 B.n836 B.n51 163.367
R2357 B.n832 B.n51 163.367
R2358 B.n832 B.n831 163.367
R2359 B.n831 B.n830 163.367
R2360 B.n830 B.n53 163.367
R2361 B.n826 B.n53 163.367
R2362 B.n826 B.n825 163.367
R2363 B.n825 B.n824 163.367
R2364 B.n824 B.n55 163.367
R2365 B.n820 B.n55 163.367
R2366 B.n820 B.n819 163.367
R2367 B.n819 B.n818 163.367
R2368 B.n818 B.n57 163.367
R2369 B.n814 B.n57 163.367
R2370 B.n814 B.n813 163.367
R2371 B.n813 B.n812 163.367
R2372 B.n812 B.n59 163.367
R2373 B.n808 B.n59 163.367
R2374 B.n808 B.n807 163.367
R2375 B.n807 B.n63 163.367
R2376 B.n803 B.n63 163.367
R2377 B.n803 B.n802 163.367
R2378 B.n802 B.n801 163.367
R2379 B.n801 B.n65 163.367
R2380 B.n797 B.n65 163.367
R2381 B.n797 B.n796 163.367
R2382 B.n796 B.n795 163.367
R2383 B.n795 B.n67 163.367
R2384 B.n790 B.n67 163.367
R2385 B.n790 B.n789 163.367
R2386 B.n789 B.n788 163.367
R2387 B.n788 B.n71 163.367
R2388 B.n784 B.n71 163.367
R2389 B.n784 B.n783 163.367
R2390 B.n783 B.n782 163.367
R2391 B.n782 B.n73 163.367
R2392 B.n778 B.n73 163.367
R2393 B.n778 B.n777 163.367
R2394 B.n777 B.n776 163.367
R2395 B.n776 B.n75 163.367
R2396 B.n772 B.n75 163.367
R2397 B.n772 B.n771 163.367
R2398 B.n771 B.n770 163.367
R2399 B.n770 B.n77 163.367
R2400 B.n766 B.n77 163.367
R2401 B.n766 B.n765 163.367
R2402 B.n765 B.n764 163.367
R2403 B.n764 B.n79 163.367
R2404 B.n760 B.n79 163.367
R2405 B.n760 B.n759 163.367
R2406 B.n759 B.n758 163.367
R2407 B.n758 B.n81 163.367
R2408 B.n754 B.n81 163.367
R2409 B.n754 B.n753 163.367
R2410 B.n753 B.n752 163.367
R2411 B.n752 B.n83 163.367
R2412 B.n748 B.n83 163.367
R2413 B.n748 B.n747 163.367
R2414 B.n747 B.n746 163.367
R2415 B.n746 B.n85 163.367
R2416 B.n742 B.n85 163.367
R2417 B.n742 B.n741 163.367
R2418 B.n741 B.n740 163.367
R2419 B.n740 B.n87 163.367
R2420 B.n736 B.n87 163.367
R2421 B.n736 B.n735 163.367
R2422 B.n735 B.n734 163.367
R2423 B.n734 B.n89 163.367
R2424 B.n730 B.n89 163.367
R2425 B.n730 B.n729 163.367
R2426 B.n729 B.n728 163.367
R2427 B.n728 B.n91 163.367
R2428 B.n724 B.n91 163.367
R2429 B.n724 B.n723 163.367
R2430 B.n723 B.n722 163.367
R2431 B.n722 B.n93 163.367
R2432 B.n718 B.n93 163.367
R2433 B.n718 B.n717 163.367
R2434 B.n717 B.n716 163.367
R2435 B.n716 B.n95 163.367
R2436 B.n712 B.n95 163.367
R2437 B.n712 B.n711 163.367
R2438 B.n711 B.n710 163.367
R2439 B.n710 B.n97 163.367
R2440 B.n706 B.n97 163.367
R2441 B.n706 B.n705 163.367
R2442 B.n705 B.n704 163.367
R2443 B.n704 B.n99 163.367
R2444 B.n700 B.n99 163.367
R2445 B.n700 B.n699 163.367
R2446 B.n187 B.n186 76.0247
R2447 B.n195 B.n194 76.0247
R2448 B.n61 B.n60 76.0247
R2449 B.n69 B.n68 76.0247
R2450 B.n188 B.n187 59.5399
R2451 B.n426 B.n195 59.5399
R2452 B.n62 B.n61 59.5399
R2453 B.n792 B.n69 59.5399
R2454 B.n901 B.n900 35.1225
R2455 B.n697 B.n100 35.1225
R2456 B.n535 B.n534 35.1225
R2457 B.n331 B.n226 35.1225
R2458 B B.n983 18.0485
R2459 B.n900 B.n899 10.6151
R2460 B.n899 B.n30 10.6151
R2461 B.n895 B.n30 10.6151
R2462 B.n895 B.n894 10.6151
R2463 B.n894 B.n893 10.6151
R2464 B.n893 B.n32 10.6151
R2465 B.n889 B.n32 10.6151
R2466 B.n889 B.n888 10.6151
R2467 B.n888 B.n887 10.6151
R2468 B.n887 B.n34 10.6151
R2469 B.n883 B.n34 10.6151
R2470 B.n883 B.n882 10.6151
R2471 B.n882 B.n881 10.6151
R2472 B.n881 B.n36 10.6151
R2473 B.n877 B.n36 10.6151
R2474 B.n877 B.n876 10.6151
R2475 B.n876 B.n875 10.6151
R2476 B.n875 B.n38 10.6151
R2477 B.n871 B.n38 10.6151
R2478 B.n871 B.n870 10.6151
R2479 B.n870 B.n869 10.6151
R2480 B.n869 B.n40 10.6151
R2481 B.n865 B.n40 10.6151
R2482 B.n865 B.n864 10.6151
R2483 B.n864 B.n863 10.6151
R2484 B.n863 B.n42 10.6151
R2485 B.n859 B.n42 10.6151
R2486 B.n859 B.n858 10.6151
R2487 B.n858 B.n857 10.6151
R2488 B.n857 B.n44 10.6151
R2489 B.n853 B.n44 10.6151
R2490 B.n853 B.n852 10.6151
R2491 B.n852 B.n851 10.6151
R2492 B.n851 B.n46 10.6151
R2493 B.n847 B.n46 10.6151
R2494 B.n847 B.n846 10.6151
R2495 B.n846 B.n845 10.6151
R2496 B.n845 B.n48 10.6151
R2497 B.n841 B.n48 10.6151
R2498 B.n841 B.n840 10.6151
R2499 B.n840 B.n839 10.6151
R2500 B.n839 B.n50 10.6151
R2501 B.n835 B.n50 10.6151
R2502 B.n835 B.n834 10.6151
R2503 B.n834 B.n833 10.6151
R2504 B.n833 B.n52 10.6151
R2505 B.n829 B.n52 10.6151
R2506 B.n829 B.n828 10.6151
R2507 B.n828 B.n827 10.6151
R2508 B.n827 B.n54 10.6151
R2509 B.n823 B.n54 10.6151
R2510 B.n823 B.n822 10.6151
R2511 B.n822 B.n821 10.6151
R2512 B.n821 B.n56 10.6151
R2513 B.n817 B.n56 10.6151
R2514 B.n817 B.n816 10.6151
R2515 B.n816 B.n815 10.6151
R2516 B.n815 B.n58 10.6151
R2517 B.n811 B.n58 10.6151
R2518 B.n811 B.n810 10.6151
R2519 B.n810 B.n809 10.6151
R2520 B.n806 B.n805 10.6151
R2521 B.n805 B.n804 10.6151
R2522 B.n804 B.n64 10.6151
R2523 B.n800 B.n64 10.6151
R2524 B.n800 B.n799 10.6151
R2525 B.n799 B.n798 10.6151
R2526 B.n798 B.n66 10.6151
R2527 B.n794 B.n66 10.6151
R2528 B.n794 B.n793 10.6151
R2529 B.n791 B.n70 10.6151
R2530 B.n787 B.n70 10.6151
R2531 B.n787 B.n786 10.6151
R2532 B.n786 B.n785 10.6151
R2533 B.n785 B.n72 10.6151
R2534 B.n781 B.n72 10.6151
R2535 B.n781 B.n780 10.6151
R2536 B.n780 B.n779 10.6151
R2537 B.n779 B.n74 10.6151
R2538 B.n775 B.n74 10.6151
R2539 B.n775 B.n774 10.6151
R2540 B.n774 B.n773 10.6151
R2541 B.n773 B.n76 10.6151
R2542 B.n769 B.n76 10.6151
R2543 B.n769 B.n768 10.6151
R2544 B.n768 B.n767 10.6151
R2545 B.n767 B.n78 10.6151
R2546 B.n763 B.n78 10.6151
R2547 B.n763 B.n762 10.6151
R2548 B.n762 B.n761 10.6151
R2549 B.n761 B.n80 10.6151
R2550 B.n757 B.n80 10.6151
R2551 B.n757 B.n756 10.6151
R2552 B.n756 B.n755 10.6151
R2553 B.n755 B.n82 10.6151
R2554 B.n751 B.n82 10.6151
R2555 B.n751 B.n750 10.6151
R2556 B.n750 B.n749 10.6151
R2557 B.n749 B.n84 10.6151
R2558 B.n745 B.n84 10.6151
R2559 B.n745 B.n744 10.6151
R2560 B.n744 B.n743 10.6151
R2561 B.n743 B.n86 10.6151
R2562 B.n739 B.n86 10.6151
R2563 B.n739 B.n738 10.6151
R2564 B.n738 B.n737 10.6151
R2565 B.n737 B.n88 10.6151
R2566 B.n733 B.n88 10.6151
R2567 B.n733 B.n732 10.6151
R2568 B.n732 B.n731 10.6151
R2569 B.n731 B.n90 10.6151
R2570 B.n727 B.n90 10.6151
R2571 B.n727 B.n726 10.6151
R2572 B.n726 B.n725 10.6151
R2573 B.n725 B.n92 10.6151
R2574 B.n721 B.n92 10.6151
R2575 B.n721 B.n720 10.6151
R2576 B.n720 B.n719 10.6151
R2577 B.n719 B.n94 10.6151
R2578 B.n715 B.n94 10.6151
R2579 B.n715 B.n714 10.6151
R2580 B.n714 B.n713 10.6151
R2581 B.n713 B.n96 10.6151
R2582 B.n709 B.n96 10.6151
R2583 B.n709 B.n708 10.6151
R2584 B.n708 B.n707 10.6151
R2585 B.n707 B.n98 10.6151
R2586 B.n703 B.n98 10.6151
R2587 B.n703 B.n702 10.6151
R2588 B.n702 B.n701 10.6151
R2589 B.n701 B.n100 10.6151
R2590 B.n535 B.n154 10.6151
R2591 B.n539 B.n154 10.6151
R2592 B.n540 B.n539 10.6151
R2593 B.n541 B.n540 10.6151
R2594 B.n541 B.n152 10.6151
R2595 B.n545 B.n152 10.6151
R2596 B.n546 B.n545 10.6151
R2597 B.n547 B.n546 10.6151
R2598 B.n547 B.n150 10.6151
R2599 B.n551 B.n150 10.6151
R2600 B.n552 B.n551 10.6151
R2601 B.n553 B.n552 10.6151
R2602 B.n553 B.n148 10.6151
R2603 B.n557 B.n148 10.6151
R2604 B.n558 B.n557 10.6151
R2605 B.n559 B.n558 10.6151
R2606 B.n559 B.n146 10.6151
R2607 B.n563 B.n146 10.6151
R2608 B.n564 B.n563 10.6151
R2609 B.n565 B.n564 10.6151
R2610 B.n565 B.n144 10.6151
R2611 B.n569 B.n144 10.6151
R2612 B.n570 B.n569 10.6151
R2613 B.n571 B.n570 10.6151
R2614 B.n571 B.n142 10.6151
R2615 B.n575 B.n142 10.6151
R2616 B.n576 B.n575 10.6151
R2617 B.n577 B.n576 10.6151
R2618 B.n577 B.n140 10.6151
R2619 B.n581 B.n140 10.6151
R2620 B.n582 B.n581 10.6151
R2621 B.n583 B.n582 10.6151
R2622 B.n583 B.n138 10.6151
R2623 B.n587 B.n138 10.6151
R2624 B.n588 B.n587 10.6151
R2625 B.n589 B.n588 10.6151
R2626 B.n589 B.n136 10.6151
R2627 B.n593 B.n136 10.6151
R2628 B.n594 B.n593 10.6151
R2629 B.n595 B.n594 10.6151
R2630 B.n595 B.n134 10.6151
R2631 B.n599 B.n134 10.6151
R2632 B.n600 B.n599 10.6151
R2633 B.n601 B.n600 10.6151
R2634 B.n601 B.n132 10.6151
R2635 B.n605 B.n132 10.6151
R2636 B.n606 B.n605 10.6151
R2637 B.n607 B.n606 10.6151
R2638 B.n607 B.n130 10.6151
R2639 B.n611 B.n130 10.6151
R2640 B.n612 B.n611 10.6151
R2641 B.n613 B.n612 10.6151
R2642 B.n613 B.n128 10.6151
R2643 B.n617 B.n128 10.6151
R2644 B.n618 B.n617 10.6151
R2645 B.n619 B.n618 10.6151
R2646 B.n619 B.n126 10.6151
R2647 B.n623 B.n126 10.6151
R2648 B.n624 B.n623 10.6151
R2649 B.n625 B.n624 10.6151
R2650 B.n625 B.n124 10.6151
R2651 B.n629 B.n124 10.6151
R2652 B.n630 B.n629 10.6151
R2653 B.n631 B.n630 10.6151
R2654 B.n631 B.n122 10.6151
R2655 B.n635 B.n122 10.6151
R2656 B.n636 B.n635 10.6151
R2657 B.n637 B.n636 10.6151
R2658 B.n637 B.n120 10.6151
R2659 B.n641 B.n120 10.6151
R2660 B.n642 B.n641 10.6151
R2661 B.n643 B.n642 10.6151
R2662 B.n643 B.n118 10.6151
R2663 B.n647 B.n118 10.6151
R2664 B.n648 B.n647 10.6151
R2665 B.n649 B.n648 10.6151
R2666 B.n649 B.n116 10.6151
R2667 B.n653 B.n116 10.6151
R2668 B.n654 B.n653 10.6151
R2669 B.n655 B.n654 10.6151
R2670 B.n655 B.n114 10.6151
R2671 B.n659 B.n114 10.6151
R2672 B.n660 B.n659 10.6151
R2673 B.n661 B.n660 10.6151
R2674 B.n661 B.n112 10.6151
R2675 B.n665 B.n112 10.6151
R2676 B.n666 B.n665 10.6151
R2677 B.n667 B.n666 10.6151
R2678 B.n667 B.n110 10.6151
R2679 B.n671 B.n110 10.6151
R2680 B.n672 B.n671 10.6151
R2681 B.n673 B.n672 10.6151
R2682 B.n673 B.n108 10.6151
R2683 B.n677 B.n108 10.6151
R2684 B.n678 B.n677 10.6151
R2685 B.n679 B.n678 10.6151
R2686 B.n679 B.n106 10.6151
R2687 B.n683 B.n106 10.6151
R2688 B.n684 B.n683 10.6151
R2689 B.n685 B.n684 10.6151
R2690 B.n685 B.n104 10.6151
R2691 B.n689 B.n104 10.6151
R2692 B.n690 B.n689 10.6151
R2693 B.n691 B.n690 10.6151
R2694 B.n691 B.n102 10.6151
R2695 B.n695 B.n102 10.6151
R2696 B.n696 B.n695 10.6151
R2697 B.n697 B.n696 10.6151
R2698 B.n335 B.n226 10.6151
R2699 B.n336 B.n335 10.6151
R2700 B.n337 B.n336 10.6151
R2701 B.n337 B.n224 10.6151
R2702 B.n341 B.n224 10.6151
R2703 B.n342 B.n341 10.6151
R2704 B.n343 B.n342 10.6151
R2705 B.n343 B.n222 10.6151
R2706 B.n347 B.n222 10.6151
R2707 B.n348 B.n347 10.6151
R2708 B.n349 B.n348 10.6151
R2709 B.n349 B.n220 10.6151
R2710 B.n353 B.n220 10.6151
R2711 B.n354 B.n353 10.6151
R2712 B.n355 B.n354 10.6151
R2713 B.n355 B.n218 10.6151
R2714 B.n359 B.n218 10.6151
R2715 B.n360 B.n359 10.6151
R2716 B.n361 B.n360 10.6151
R2717 B.n361 B.n216 10.6151
R2718 B.n365 B.n216 10.6151
R2719 B.n366 B.n365 10.6151
R2720 B.n367 B.n366 10.6151
R2721 B.n367 B.n214 10.6151
R2722 B.n371 B.n214 10.6151
R2723 B.n372 B.n371 10.6151
R2724 B.n373 B.n372 10.6151
R2725 B.n373 B.n212 10.6151
R2726 B.n377 B.n212 10.6151
R2727 B.n378 B.n377 10.6151
R2728 B.n379 B.n378 10.6151
R2729 B.n379 B.n210 10.6151
R2730 B.n383 B.n210 10.6151
R2731 B.n384 B.n383 10.6151
R2732 B.n385 B.n384 10.6151
R2733 B.n385 B.n208 10.6151
R2734 B.n389 B.n208 10.6151
R2735 B.n390 B.n389 10.6151
R2736 B.n391 B.n390 10.6151
R2737 B.n391 B.n206 10.6151
R2738 B.n395 B.n206 10.6151
R2739 B.n396 B.n395 10.6151
R2740 B.n397 B.n396 10.6151
R2741 B.n397 B.n204 10.6151
R2742 B.n401 B.n204 10.6151
R2743 B.n402 B.n401 10.6151
R2744 B.n403 B.n402 10.6151
R2745 B.n403 B.n202 10.6151
R2746 B.n407 B.n202 10.6151
R2747 B.n408 B.n407 10.6151
R2748 B.n409 B.n408 10.6151
R2749 B.n409 B.n200 10.6151
R2750 B.n413 B.n200 10.6151
R2751 B.n414 B.n413 10.6151
R2752 B.n415 B.n414 10.6151
R2753 B.n415 B.n198 10.6151
R2754 B.n419 B.n198 10.6151
R2755 B.n420 B.n419 10.6151
R2756 B.n421 B.n420 10.6151
R2757 B.n421 B.n196 10.6151
R2758 B.n425 B.n196 10.6151
R2759 B.n428 B.n427 10.6151
R2760 B.n428 B.n192 10.6151
R2761 B.n432 B.n192 10.6151
R2762 B.n433 B.n432 10.6151
R2763 B.n434 B.n433 10.6151
R2764 B.n434 B.n190 10.6151
R2765 B.n438 B.n190 10.6151
R2766 B.n439 B.n438 10.6151
R2767 B.n440 B.n439 10.6151
R2768 B.n444 B.n443 10.6151
R2769 B.n445 B.n444 10.6151
R2770 B.n445 B.n184 10.6151
R2771 B.n449 B.n184 10.6151
R2772 B.n450 B.n449 10.6151
R2773 B.n451 B.n450 10.6151
R2774 B.n451 B.n182 10.6151
R2775 B.n455 B.n182 10.6151
R2776 B.n456 B.n455 10.6151
R2777 B.n457 B.n456 10.6151
R2778 B.n457 B.n180 10.6151
R2779 B.n461 B.n180 10.6151
R2780 B.n462 B.n461 10.6151
R2781 B.n463 B.n462 10.6151
R2782 B.n463 B.n178 10.6151
R2783 B.n467 B.n178 10.6151
R2784 B.n468 B.n467 10.6151
R2785 B.n469 B.n468 10.6151
R2786 B.n469 B.n176 10.6151
R2787 B.n473 B.n176 10.6151
R2788 B.n474 B.n473 10.6151
R2789 B.n475 B.n474 10.6151
R2790 B.n475 B.n174 10.6151
R2791 B.n479 B.n174 10.6151
R2792 B.n480 B.n479 10.6151
R2793 B.n481 B.n480 10.6151
R2794 B.n481 B.n172 10.6151
R2795 B.n485 B.n172 10.6151
R2796 B.n486 B.n485 10.6151
R2797 B.n487 B.n486 10.6151
R2798 B.n487 B.n170 10.6151
R2799 B.n491 B.n170 10.6151
R2800 B.n492 B.n491 10.6151
R2801 B.n493 B.n492 10.6151
R2802 B.n493 B.n168 10.6151
R2803 B.n497 B.n168 10.6151
R2804 B.n498 B.n497 10.6151
R2805 B.n499 B.n498 10.6151
R2806 B.n499 B.n166 10.6151
R2807 B.n503 B.n166 10.6151
R2808 B.n504 B.n503 10.6151
R2809 B.n505 B.n504 10.6151
R2810 B.n505 B.n164 10.6151
R2811 B.n509 B.n164 10.6151
R2812 B.n510 B.n509 10.6151
R2813 B.n511 B.n510 10.6151
R2814 B.n511 B.n162 10.6151
R2815 B.n515 B.n162 10.6151
R2816 B.n516 B.n515 10.6151
R2817 B.n517 B.n516 10.6151
R2818 B.n517 B.n160 10.6151
R2819 B.n521 B.n160 10.6151
R2820 B.n522 B.n521 10.6151
R2821 B.n523 B.n522 10.6151
R2822 B.n523 B.n158 10.6151
R2823 B.n527 B.n158 10.6151
R2824 B.n528 B.n527 10.6151
R2825 B.n529 B.n528 10.6151
R2826 B.n529 B.n156 10.6151
R2827 B.n533 B.n156 10.6151
R2828 B.n534 B.n533 10.6151
R2829 B.n331 B.n330 10.6151
R2830 B.n330 B.n329 10.6151
R2831 B.n329 B.n228 10.6151
R2832 B.n325 B.n228 10.6151
R2833 B.n325 B.n324 10.6151
R2834 B.n324 B.n323 10.6151
R2835 B.n323 B.n230 10.6151
R2836 B.n319 B.n230 10.6151
R2837 B.n319 B.n318 10.6151
R2838 B.n318 B.n317 10.6151
R2839 B.n317 B.n232 10.6151
R2840 B.n313 B.n232 10.6151
R2841 B.n313 B.n312 10.6151
R2842 B.n312 B.n311 10.6151
R2843 B.n311 B.n234 10.6151
R2844 B.n307 B.n234 10.6151
R2845 B.n307 B.n306 10.6151
R2846 B.n306 B.n305 10.6151
R2847 B.n305 B.n236 10.6151
R2848 B.n301 B.n236 10.6151
R2849 B.n301 B.n300 10.6151
R2850 B.n300 B.n299 10.6151
R2851 B.n299 B.n238 10.6151
R2852 B.n295 B.n238 10.6151
R2853 B.n295 B.n294 10.6151
R2854 B.n294 B.n293 10.6151
R2855 B.n293 B.n240 10.6151
R2856 B.n289 B.n240 10.6151
R2857 B.n289 B.n288 10.6151
R2858 B.n288 B.n287 10.6151
R2859 B.n287 B.n242 10.6151
R2860 B.n283 B.n242 10.6151
R2861 B.n283 B.n282 10.6151
R2862 B.n282 B.n281 10.6151
R2863 B.n281 B.n244 10.6151
R2864 B.n277 B.n244 10.6151
R2865 B.n277 B.n276 10.6151
R2866 B.n276 B.n275 10.6151
R2867 B.n275 B.n246 10.6151
R2868 B.n271 B.n246 10.6151
R2869 B.n271 B.n270 10.6151
R2870 B.n270 B.n269 10.6151
R2871 B.n269 B.n248 10.6151
R2872 B.n265 B.n248 10.6151
R2873 B.n265 B.n264 10.6151
R2874 B.n264 B.n263 10.6151
R2875 B.n263 B.n250 10.6151
R2876 B.n259 B.n250 10.6151
R2877 B.n259 B.n258 10.6151
R2878 B.n258 B.n257 10.6151
R2879 B.n257 B.n252 10.6151
R2880 B.n253 B.n252 10.6151
R2881 B.n253 B.n0 10.6151
R2882 B.n979 B.n1 10.6151
R2883 B.n979 B.n978 10.6151
R2884 B.n978 B.n977 10.6151
R2885 B.n977 B.n4 10.6151
R2886 B.n973 B.n4 10.6151
R2887 B.n973 B.n972 10.6151
R2888 B.n972 B.n971 10.6151
R2889 B.n971 B.n6 10.6151
R2890 B.n967 B.n6 10.6151
R2891 B.n967 B.n966 10.6151
R2892 B.n966 B.n965 10.6151
R2893 B.n965 B.n8 10.6151
R2894 B.n961 B.n8 10.6151
R2895 B.n961 B.n960 10.6151
R2896 B.n960 B.n959 10.6151
R2897 B.n959 B.n10 10.6151
R2898 B.n955 B.n10 10.6151
R2899 B.n955 B.n954 10.6151
R2900 B.n954 B.n953 10.6151
R2901 B.n953 B.n12 10.6151
R2902 B.n949 B.n12 10.6151
R2903 B.n949 B.n948 10.6151
R2904 B.n948 B.n947 10.6151
R2905 B.n947 B.n14 10.6151
R2906 B.n943 B.n14 10.6151
R2907 B.n943 B.n942 10.6151
R2908 B.n942 B.n941 10.6151
R2909 B.n941 B.n16 10.6151
R2910 B.n937 B.n16 10.6151
R2911 B.n937 B.n936 10.6151
R2912 B.n936 B.n935 10.6151
R2913 B.n935 B.n18 10.6151
R2914 B.n931 B.n18 10.6151
R2915 B.n931 B.n930 10.6151
R2916 B.n930 B.n929 10.6151
R2917 B.n929 B.n20 10.6151
R2918 B.n925 B.n20 10.6151
R2919 B.n925 B.n924 10.6151
R2920 B.n924 B.n923 10.6151
R2921 B.n923 B.n22 10.6151
R2922 B.n919 B.n22 10.6151
R2923 B.n919 B.n918 10.6151
R2924 B.n918 B.n917 10.6151
R2925 B.n917 B.n24 10.6151
R2926 B.n913 B.n24 10.6151
R2927 B.n913 B.n912 10.6151
R2928 B.n912 B.n911 10.6151
R2929 B.n911 B.n26 10.6151
R2930 B.n907 B.n26 10.6151
R2931 B.n907 B.n906 10.6151
R2932 B.n906 B.n905 10.6151
R2933 B.n905 B.n28 10.6151
R2934 B.n901 B.n28 10.6151
R2935 B.n809 B.n62 9.36635
R2936 B.n792 B.n791 9.36635
R2937 B.n426 B.n425 9.36635
R2938 B.n443 B.n188 9.36635
R2939 B.n983 B.n0 2.81026
R2940 B.n983 B.n1 2.81026
R2941 B.n806 B.n62 1.24928
R2942 B.n793 B.n792 1.24928
R2943 B.n427 B.n426 1.24928
R2944 B.n440 B.n188 1.24928
C0 VP B 2.35432f
C1 VDD1 VDD2 1.79451f
C2 VN B 1.45842f
C3 VTAIL B 5.72478f
C4 VDD2 w_n4106_n4770# 3.12849f
C5 VP VN 9.18762f
C6 VDD1 B 2.91524f
C7 VTAIL VP 11.0783f
C8 VDD1 VP 11.385201f
C9 VTAIL VN 11.0639f
C10 w_n4106_n4770# B 13.0088f
C11 VDD1 VN 0.152188f
C12 VP w_n4106_n4770# 8.68005f
C13 VTAIL VDD1 10.3325f
C14 VN w_n4106_n4770# 8.146441f
C15 VTAIL w_n4106_n4770# 4.01335f
C16 VDD2 B 3.01307f
C17 VDD1 w_n4106_n4770# 3.01177f
C18 VP VDD2 0.5427f
C19 VN VDD2 10.9986f
C20 VTAIL VDD2 10.3897f
C21 VDD2 VSUBS 2.34577f
C22 VDD1 VSUBS 2.351966f
C23 VTAIL VSUBS 1.63051f
C24 VN VSUBS 7.061f
C25 VP VSUBS 3.959883f
C26 B VSUBS 6.207049f
C27 w_n4106_n4770# VSUBS 0.239314p
C28 B.n0 VSUBS 0.004491f
C29 B.n1 VSUBS 0.004491f
C30 B.n2 VSUBS 0.007102f
C31 B.n3 VSUBS 0.007102f
C32 B.n4 VSUBS 0.007102f
C33 B.n5 VSUBS 0.007102f
C34 B.n6 VSUBS 0.007102f
C35 B.n7 VSUBS 0.007102f
C36 B.n8 VSUBS 0.007102f
C37 B.n9 VSUBS 0.007102f
C38 B.n10 VSUBS 0.007102f
C39 B.n11 VSUBS 0.007102f
C40 B.n12 VSUBS 0.007102f
C41 B.n13 VSUBS 0.007102f
C42 B.n14 VSUBS 0.007102f
C43 B.n15 VSUBS 0.007102f
C44 B.n16 VSUBS 0.007102f
C45 B.n17 VSUBS 0.007102f
C46 B.n18 VSUBS 0.007102f
C47 B.n19 VSUBS 0.007102f
C48 B.n20 VSUBS 0.007102f
C49 B.n21 VSUBS 0.007102f
C50 B.n22 VSUBS 0.007102f
C51 B.n23 VSUBS 0.007102f
C52 B.n24 VSUBS 0.007102f
C53 B.n25 VSUBS 0.007102f
C54 B.n26 VSUBS 0.007102f
C55 B.n27 VSUBS 0.007102f
C56 B.n28 VSUBS 0.007102f
C57 B.n29 VSUBS 0.017945f
C58 B.n30 VSUBS 0.007102f
C59 B.n31 VSUBS 0.007102f
C60 B.n32 VSUBS 0.007102f
C61 B.n33 VSUBS 0.007102f
C62 B.n34 VSUBS 0.007102f
C63 B.n35 VSUBS 0.007102f
C64 B.n36 VSUBS 0.007102f
C65 B.n37 VSUBS 0.007102f
C66 B.n38 VSUBS 0.007102f
C67 B.n39 VSUBS 0.007102f
C68 B.n40 VSUBS 0.007102f
C69 B.n41 VSUBS 0.007102f
C70 B.n42 VSUBS 0.007102f
C71 B.n43 VSUBS 0.007102f
C72 B.n44 VSUBS 0.007102f
C73 B.n45 VSUBS 0.007102f
C74 B.n46 VSUBS 0.007102f
C75 B.n47 VSUBS 0.007102f
C76 B.n48 VSUBS 0.007102f
C77 B.n49 VSUBS 0.007102f
C78 B.n50 VSUBS 0.007102f
C79 B.n51 VSUBS 0.007102f
C80 B.n52 VSUBS 0.007102f
C81 B.n53 VSUBS 0.007102f
C82 B.n54 VSUBS 0.007102f
C83 B.n55 VSUBS 0.007102f
C84 B.n56 VSUBS 0.007102f
C85 B.n57 VSUBS 0.007102f
C86 B.n58 VSUBS 0.007102f
C87 B.n59 VSUBS 0.007102f
C88 B.t2 VSUBS 0.381267f
C89 B.t1 VSUBS 0.425909f
C90 B.t0 VSUBS 3.13202f
C91 B.n60 VSUBS 0.678055f
C92 B.n61 VSUBS 0.349601f
C93 B.n62 VSUBS 0.016454f
C94 B.n63 VSUBS 0.007102f
C95 B.n64 VSUBS 0.007102f
C96 B.n65 VSUBS 0.007102f
C97 B.n66 VSUBS 0.007102f
C98 B.n67 VSUBS 0.007102f
C99 B.t5 VSUBS 0.38127f
C100 B.t4 VSUBS 0.425912f
C101 B.t3 VSUBS 3.13202f
C102 B.n68 VSUBS 0.678052f
C103 B.n69 VSUBS 0.349597f
C104 B.n70 VSUBS 0.007102f
C105 B.n71 VSUBS 0.007102f
C106 B.n72 VSUBS 0.007102f
C107 B.n73 VSUBS 0.007102f
C108 B.n74 VSUBS 0.007102f
C109 B.n75 VSUBS 0.007102f
C110 B.n76 VSUBS 0.007102f
C111 B.n77 VSUBS 0.007102f
C112 B.n78 VSUBS 0.007102f
C113 B.n79 VSUBS 0.007102f
C114 B.n80 VSUBS 0.007102f
C115 B.n81 VSUBS 0.007102f
C116 B.n82 VSUBS 0.007102f
C117 B.n83 VSUBS 0.007102f
C118 B.n84 VSUBS 0.007102f
C119 B.n85 VSUBS 0.007102f
C120 B.n86 VSUBS 0.007102f
C121 B.n87 VSUBS 0.007102f
C122 B.n88 VSUBS 0.007102f
C123 B.n89 VSUBS 0.007102f
C124 B.n90 VSUBS 0.007102f
C125 B.n91 VSUBS 0.007102f
C126 B.n92 VSUBS 0.007102f
C127 B.n93 VSUBS 0.007102f
C128 B.n94 VSUBS 0.007102f
C129 B.n95 VSUBS 0.007102f
C130 B.n96 VSUBS 0.007102f
C131 B.n97 VSUBS 0.007102f
C132 B.n98 VSUBS 0.007102f
C133 B.n99 VSUBS 0.007102f
C134 B.n100 VSUBS 0.017165f
C135 B.n101 VSUBS 0.007102f
C136 B.n102 VSUBS 0.007102f
C137 B.n103 VSUBS 0.007102f
C138 B.n104 VSUBS 0.007102f
C139 B.n105 VSUBS 0.007102f
C140 B.n106 VSUBS 0.007102f
C141 B.n107 VSUBS 0.007102f
C142 B.n108 VSUBS 0.007102f
C143 B.n109 VSUBS 0.007102f
C144 B.n110 VSUBS 0.007102f
C145 B.n111 VSUBS 0.007102f
C146 B.n112 VSUBS 0.007102f
C147 B.n113 VSUBS 0.007102f
C148 B.n114 VSUBS 0.007102f
C149 B.n115 VSUBS 0.007102f
C150 B.n116 VSUBS 0.007102f
C151 B.n117 VSUBS 0.007102f
C152 B.n118 VSUBS 0.007102f
C153 B.n119 VSUBS 0.007102f
C154 B.n120 VSUBS 0.007102f
C155 B.n121 VSUBS 0.007102f
C156 B.n122 VSUBS 0.007102f
C157 B.n123 VSUBS 0.007102f
C158 B.n124 VSUBS 0.007102f
C159 B.n125 VSUBS 0.007102f
C160 B.n126 VSUBS 0.007102f
C161 B.n127 VSUBS 0.007102f
C162 B.n128 VSUBS 0.007102f
C163 B.n129 VSUBS 0.007102f
C164 B.n130 VSUBS 0.007102f
C165 B.n131 VSUBS 0.007102f
C166 B.n132 VSUBS 0.007102f
C167 B.n133 VSUBS 0.007102f
C168 B.n134 VSUBS 0.007102f
C169 B.n135 VSUBS 0.007102f
C170 B.n136 VSUBS 0.007102f
C171 B.n137 VSUBS 0.007102f
C172 B.n138 VSUBS 0.007102f
C173 B.n139 VSUBS 0.007102f
C174 B.n140 VSUBS 0.007102f
C175 B.n141 VSUBS 0.007102f
C176 B.n142 VSUBS 0.007102f
C177 B.n143 VSUBS 0.007102f
C178 B.n144 VSUBS 0.007102f
C179 B.n145 VSUBS 0.007102f
C180 B.n146 VSUBS 0.007102f
C181 B.n147 VSUBS 0.007102f
C182 B.n148 VSUBS 0.007102f
C183 B.n149 VSUBS 0.007102f
C184 B.n150 VSUBS 0.007102f
C185 B.n151 VSUBS 0.007102f
C186 B.n152 VSUBS 0.007102f
C187 B.n153 VSUBS 0.007102f
C188 B.n154 VSUBS 0.007102f
C189 B.n155 VSUBS 0.017945f
C190 B.n156 VSUBS 0.007102f
C191 B.n157 VSUBS 0.007102f
C192 B.n158 VSUBS 0.007102f
C193 B.n159 VSUBS 0.007102f
C194 B.n160 VSUBS 0.007102f
C195 B.n161 VSUBS 0.007102f
C196 B.n162 VSUBS 0.007102f
C197 B.n163 VSUBS 0.007102f
C198 B.n164 VSUBS 0.007102f
C199 B.n165 VSUBS 0.007102f
C200 B.n166 VSUBS 0.007102f
C201 B.n167 VSUBS 0.007102f
C202 B.n168 VSUBS 0.007102f
C203 B.n169 VSUBS 0.007102f
C204 B.n170 VSUBS 0.007102f
C205 B.n171 VSUBS 0.007102f
C206 B.n172 VSUBS 0.007102f
C207 B.n173 VSUBS 0.007102f
C208 B.n174 VSUBS 0.007102f
C209 B.n175 VSUBS 0.007102f
C210 B.n176 VSUBS 0.007102f
C211 B.n177 VSUBS 0.007102f
C212 B.n178 VSUBS 0.007102f
C213 B.n179 VSUBS 0.007102f
C214 B.n180 VSUBS 0.007102f
C215 B.n181 VSUBS 0.007102f
C216 B.n182 VSUBS 0.007102f
C217 B.n183 VSUBS 0.007102f
C218 B.n184 VSUBS 0.007102f
C219 B.n185 VSUBS 0.007102f
C220 B.t10 VSUBS 0.38127f
C221 B.t11 VSUBS 0.425912f
C222 B.t9 VSUBS 3.13202f
C223 B.n186 VSUBS 0.678052f
C224 B.n187 VSUBS 0.349597f
C225 B.n188 VSUBS 0.016454f
C226 B.n189 VSUBS 0.007102f
C227 B.n190 VSUBS 0.007102f
C228 B.n191 VSUBS 0.007102f
C229 B.n192 VSUBS 0.007102f
C230 B.n193 VSUBS 0.007102f
C231 B.t7 VSUBS 0.381267f
C232 B.t8 VSUBS 0.425909f
C233 B.t6 VSUBS 3.13202f
C234 B.n194 VSUBS 0.678055f
C235 B.n195 VSUBS 0.349601f
C236 B.n196 VSUBS 0.007102f
C237 B.n197 VSUBS 0.007102f
C238 B.n198 VSUBS 0.007102f
C239 B.n199 VSUBS 0.007102f
C240 B.n200 VSUBS 0.007102f
C241 B.n201 VSUBS 0.007102f
C242 B.n202 VSUBS 0.007102f
C243 B.n203 VSUBS 0.007102f
C244 B.n204 VSUBS 0.007102f
C245 B.n205 VSUBS 0.007102f
C246 B.n206 VSUBS 0.007102f
C247 B.n207 VSUBS 0.007102f
C248 B.n208 VSUBS 0.007102f
C249 B.n209 VSUBS 0.007102f
C250 B.n210 VSUBS 0.007102f
C251 B.n211 VSUBS 0.007102f
C252 B.n212 VSUBS 0.007102f
C253 B.n213 VSUBS 0.007102f
C254 B.n214 VSUBS 0.007102f
C255 B.n215 VSUBS 0.007102f
C256 B.n216 VSUBS 0.007102f
C257 B.n217 VSUBS 0.007102f
C258 B.n218 VSUBS 0.007102f
C259 B.n219 VSUBS 0.007102f
C260 B.n220 VSUBS 0.007102f
C261 B.n221 VSUBS 0.007102f
C262 B.n222 VSUBS 0.007102f
C263 B.n223 VSUBS 0.007102f
C264 B.n224 VSUBS 0.007102f
C265 B.n225 VSUBS 0.007102f
C266 B.n226 VSUBS 0.017945f
C267 B.n227 VSUBS 0.007102f
C268 B.n228 VSUBS 0.007102f
C269 B.n229 VSUBS 0.007102f
C270 B.n230 VSUBS 0.007102f
C271 B.n231 VSUBS 0.007102f
C272 B.n232 VSUBS 0.007102f
C273 B.n233 VSUBS 0.007102f
C274 B.n234 VSUBS 0.007102f
C275 B.n235 VSUBS 0.007102f
C276 B.n236 VSUBS 0.007102f
C277 B.n237 VSUBS 0.007102f
C278 B.n238 VSUBS 0.007102f
C279 B.n239 VSUBS 0.007102f
C280 B.n240 VSUBS 0.007102f
C281 B.n241 VSUBS 0.007102f
C282 B.n242 VSUBS 0.007102f
C283 B.n243 VSUBS 0.007102f
C284 B.n244 VSUBS 0.007102f
C285 B.n245 VSUBS 0.007102f
C286 B.n246 VSUBS 0.007102f
C287 B.n247 VSUBS 0.007102f
C288 B.n248 VSUBS 0.007102f
C289 B.n249 VSUBS 0.007102f
C290 B.n250 VSUBS 0.007102f
C291 B.n251 VSUBS 0.007102f
C292 B.n252 VSUBS 0.007102f
C293 B.n253 VSUBS 0.007102f
C294 B.n254 VSUBS 0.007102f
C295 B.n255 VSUBS 0.007102f
C296 B.n256 VSUBS 0.007102f
C297 B.n257 VSUBS 0.007102f
C298 B.n258 VSUBS 0.007102f
C299 B.n259 VSUBS 0.007102f
C300 B.n260 VSUBS 0.007102f
C301 B.n261 VSUBS 0.007102f
C302 B.n262 VSUBS 0.007102f
C303 B.n263 VSUBS 0.007102f
C304 B.n264 VSUBS 0.007102f
C305 B.n265 VSUBS 0.007102f
C306 B.n266 VSUBS 0.007102f
C307 B.n267 VSUBS 0.007102f
C308 B.n268 VSUBS 0.007102f
C309 B.n269 VSUBS 0.007102f
C310 B.n270 VSUBS 0.007102f
C311 B.n271 VSUBS 0.007102f
C312 B.n272 VSUBS 0.007102f
C313 B.n273 VSUBS 0.007102f
C314 B.n274 VSUBS 0.007102f
C315 B.n275 VSUBS 0.007102f
C316 B.n276 VSUBS 0.007102f
C317 B.n277 VSUBS 0.007102f
C318 B.n278 VSUBS 0.007102f
C319 B.n279 VSUBS 0.007102f
C320 B.n280 VSUBS 0.007102f
C321 B.n281 VSUBS 0.007102f
C322 B.n282 VSUBS 0.007102f
C323 B.n283 VSUBS 0.007102f
C324 B.n284 VSUBS 0.007102f
C325 B.n285 VSUBS 0.007102f
C326 B.n286 VSUBS 0.007102f
C327 B.n287 VSUBS 0.007102f
C328 B.n288 VSUBS 0.007102f
C329 B.n289 VSUBS 0.007102f
C330 B.n290 VSUBS 0.007102f
C331 B.n291 VSUBS 0.007102f
C332 B.n292 VSUBS 0.007102f
C333 B.n293 VSUBS 0.007102f
C334 B.n294 VSUBS 0.007102f
C335 B.n295 VSUBS 0.007102f
C336 B.n296 VSUBS 0.007102f
C337 B.n297 VSUBS 0.007102f
C338 B.n298 VSUBS 0.007102f
C339 B.n299 VSUBS 0.007102f
C340 B.n300 VSUBS 0.007102f
C341 B.n301 VSUBS 0.007102f
C342 B.n302 VSUBS 0.007102f
C343 B.n303 VSUBS 0.007102f
C344 B.n304 VSUBS 0.007102f
C345 B.n305 VSUBS 0.007102f
C346 B.n306 VSUBS 0.007102f
C347 B.n307 VSUBS 0.007102f
C348 B.n308 VSUBS 0.007102f
C349 B.n309 VSUBS 0.007102f
C350 B.n310 VSUBS 0.007102f
C351 B.n311 VSUBS 0.007102f
C352 B.n312 VSUBS 0.007102f
C353 B.n313 VSUBS 0.007102f
C354 B.n314 VSUBS 0.007102f
C355 B.n315 VSUBS 0.007102f
C356 B.n316 VSUBS 0.007102f
C357 B.n317 VSUBS 0.007102f
C358 B.n318 VSUBS 0.007102f
C359 B.n319 VSUBS 0.007102f
C360 B.n320 VSUBS 0.007102f
C361 B.n321 VSUBS 0.007102f
C362 B.n322 VSUBS 0.007102f
C363 B.n323 VSUBS 0.007102f
C364 B.n324 VSUBS 0.007102f
C365 B.n325 VSUBS 0.007102f
C366 B.n326 VSUBS 0.007102f
C367 B.n327 VSUBS 0.007102f
C368 B.n328 VSUBS 0.007102f
C369 B.n329 VSUBS 0.007102f
C370 B.n330 VSUBS 0.007102f
C371 B.n331 VSUBS 0.016936f
C372 B.n332 VSUBS 0.016936f
C373 B.n333 VSUBS 0.017945f
C374 B.n334 VSUBS 0.007102f
C375 B.n335 VSUBS 0.007102f
C376 B.n336 VSUBS 0.007102f
C377 B.n337 VSUBS 0.007102f
C378 B.n338 VSUBS 0.007102f
C379 B.n339 VSUBS 0.007102f
C380 B.n340 VSUBS 0.007102f
C381 B.n341 VSUBS 0.007102f
C382 B.n342 VSUBS 0.007102f
C383 B.n343 VSUBS 0.007102f
C384 B.n344 VSUBS 0.007102f
C385 B.n345 VSUBS 0.007102f
C386 B.n346 VSUBS 0.007102f
C387 B.n347 VSUBS 0.007102f
C388 B.n348 VSUBS 0.007102f
C389 B.n349 VSUBS 0.007102f
C390 B.n350 VSUBS 0.007102f
C391 B.n351 VSUBS 0.007102f
C392 B.n352 VSUBS 0.007102f
C393 B.n353 VSUBS 0.007102f
C394 B.n354 VSUBS 0.007102f
C395 B.n355 VSUBS 0.007102f
C396 B.n356 VSUBS 0.007102f
C397 B.n357 VSUBS 0.007102f
C398 B.n358 VSUBS 0.007102f
C399 B.n359 VSUBS 0.007102f
C400 B.n360 VSUBS 0.007102f
C401 B.n361 VSUBS 0.007102f
C402 B.n362 VSUBS 0.007102f
C403 B.n363 VSUBS 0.007102f
C404 B.n364 VSUBS 0.007102f
C405 B.n365 VSUBS 0.007102f
C406 B.n366 VSUBS 0.007102f
C407 B.n367 VSUBS 0.007102f
C408 B.n368 VSUBS 0.007102f
C409 B.n369 VSUBS 0.007102f
C410 B.n370 VSUBS 0.007102f
C411 B.n371 VSUBS 0.007102f
C412 B.n372 VSUBS 0.007102f
C413 B.n373 VSUBS 0.007102f
C414 B.n374 VSUBS 0.007102f
C415 B.n375 VSUBS 0.007102f
C416 B.n376 VSUBS 0.007102f
C417 B.n377 VSUBS 0.007102f
C418 B.n378 VSUBS 0.007102f
C419 B.n379 VSUBS 0.007102f
C420 B.n380 VSUBS 0.007102f
C421 B.n381 VSUBS 0.007102f
C422 B.n382 VSUBS 0.007102f
C423 B.n383 VSUBS 0.007102f
C424 B.n384 VSUBS 0.007102f
C425 B.n385 VSUBS 0.007102f
C426 B.n386 VSUBS 0.007102f
C427 B.n387 VSUBS 0.007102f
C428 B.n388 VSUBS 0.007102f
C429 B.n389 VSUBS 0.007102f
C430 B.n390 VSUBS 0.007102f
C431 B.n391 VSUBS 0.007102f
C432 B.n392 VSUBS 0.007102f
C433 B.n393 VSUBS 0.007102f
C434 B.n394 VSUBS 0.007102f
C435 B.n395 VSUBS 0.007102f
C436 B.n396 VSUBS 0.007102f
C437 B.n397 VSUBS 0.007102f
C438 B.n398 VSUBS 0.007102f
C439 B.n399 VSUBS 0.007102f
C440 B.n400 VSUBS 0.007102f
C441 B.n401 VSUBS 0.007102f
C442 B.n402 VSUBS 0.007102f
C443 B.n403 VSUBS 0.007102f
C444 B.n404 VSUBS 0.007102f
C445 B.n405 VSUBS 0.007102f
C446 B.n406 VSUBS 0.007102f
C447 B.n407 VSUBS 0.007102f
C448 B.n408 VSUBS 0.007102f
C449 B.n409 VSUBS 0.007102f
C450 B.n410 VSUBS 0.007102f
C451 B.n411 VSUBS 0.007102f
C452 B.n412 VSUBS 0.007102f
C453 B.n413 VSUBS 0.007102f
C454 B.n414 VSUBS 0.007102f
C455 B.n415 VSUBS 0.007102f
C456 B.n416 VSUBS 0.007102f
C457 B.n417 VSUBS 0.007102f
C458 B.n418 VSUBS 0.007102f
C459 B.n419 VSUBS 0.007102f
C460 B.n420 VSUBS 0.007102f
C461 B.n421 VSUBS 0.007102f
C462 B.n422 VSUBS 0.007102f
C463 B.n423 VSUBS 0.007102f
C464 B.n424 VSUBS 0.007102f
C465 B.n425 VSUBS 0.006684f
C466 B.n426 VSUBS 0.016454f
C467 B.n427 VSUBS 0.003969f
C468 B.n428 VSUBS 0.007102f
C469 B.n429 VSUBS 0.007102f
C470 B.n430 VSUBS 0.007102f
C471 B.n431 VSUBS 0.007102f
C472 B.n432 VSUBS 0.007102f
C473 B.n433 VSUBS 0.007102f
C474 B.n434 VSUBS 0.007102f
C475 B.n435 VSUBS 0.007102f
C476 B.n436 VSUBS 0.007102f
C477 B.n437 VSUBS 0.007102f
C478 B.n438 VSUBS 0.007102f
C479 B.n439 VSUBS 0.007102f
C480 B.n440 VSUBS 0.003969f
C481 B.n441 VSUBS 0.007102f
C482 B.n442 VSUBS 0.007102f
C483 B.n443 VSUBS 0.006684f
C484 B.n444 VSUBS 0.007102f
C485 B.n445 VSUBS 0.007102f
C486 B.n446 VSUBS 0.007102f
C487 B.n447 VSUBS 0.007102f
C488 B.n448 VSUBS 0.007102f
C489 B.n449 VSUBS 0.007102f
C490 B.n450 VSUBS 0.007102f
C491 B.n451 VSUBS 0.007102f
C492 B.n452 VSUBS 0.007102f
C493 B.n453 VSUBS 0.007102f
C494 B.n454 VSUBS 0.007102f
C495 B.n455 VSUBS 0.007102f
C496 B.n456 VSUBS 0.007102f
C497 B.n457 VSUBS 0.007102f
C498 B.n458 VSUBS 0.007102f
C499 B.n459 VSUBS 0.007102f
C500 B.n460 VSUBS 0.007102f
C501 B.n461 VSUBS 0.007102f
C502 B.n462 VSUBS 0.007102f
C503 B.n463 VSUBS 0.007102f
C504 B.n464 VSUBS 0.007102f
C505 B.n465 VSUBS 0.007102f
C506 B.n466 VSUBS 0.007102f
C507 B.n467 VSUBS 0.007102f
C508 B.n468 VSUBS 0.007102f
C509 B.n469 VSUBS 0.007102f
C510 B.n470 VSUBS 0.007102f
C511 B.n471 VSUBS 0.007102f
C512 B.n472 VSUBS 0.007102f
C513 B.n473 VSUBS 0.007102f
C514 B.n474 VSUBS 0.007102f
C515 B.n475 VSUBS 0.007102f
C516 B.n476 VSUBS 0.007102f
C517 B.n477 VSUBS 0.007102f
C518 B.n478 VSUBS 0.007102f
C519 B.n479 VSUBS 0.007102f
C520 B.n480 VSUBS 0.007102f
C521 B.n481 VSUBS 0.007102f
C522 B.n482 VSUBS 0.007102f
C523 B.n483 VSUBS 0.007102f
C524 B.n484 VSUBS 0.007102f
C525 B.n485 VSUBS 0.007102f
C526 B.n486 VSUBS 0.007102f
C527 B.n487 VSUBS 0.007102f
C528 B.n488 VSUBS 0.007102f
C529 B.n489 VSUBS 0.007102f
C530 B.n490 VSUBS 0.007102f
C531 B.n491 VSUBS 0.007102f
C532 B.n492 VSUBS 0.007102f
C533 B.n493 VSUBS 0.007102f
C534 B.n494 VSUBS 0.007102f
C535 B.n495 VSUBS 0.007102f
C536 B.n496 VSUBS 0.007102f
C537 B.n497 VSUBS 0.007102f
C538 B.n498 VSUBS 0.007102f
C539 B.n499 VSUBS 0.007102f
C540 B.n500 VSUBS 0.007102f
C541 B.n501 VSUBS 0.007102f
C542 B.n502 VSUBS 0.007102f
C543 B.n503 VSUBS 0.007102f
C544 B.n504 VSUBS 0.007102f
C545 B.n505 VSUBS 0.007102f
C546 B.n506 VSUBS 0.007102f
C547 B.n507 VSUBS 0.007102f
C548 B.n508 VSUBS 0.007102f
C549 B.n509 VSUBS 0.007102f
C550 B.n510 VSUBS 0.007102f
C551 B.n511 VSUBS 0.007102f
C552 B.n512 VSUBS 0.007102f
C553 B.n513 VSUBS 0.007102f
C554 B.n514 VSUBS 0.007102f
C555 B.n515 VSUBS 0.007102f
C556 B.n516 VSUBS 0.007102f
C557 B.n517 VSUBS 0.007102f
C558 B.n518 VSUBS 0.007102f
C559 B.n519 VSUBS 0.007102f
C560 B.n520 VSUBS 0.007102f
C561 B.n521 VSUBS 0.007102f
C562 B.n522 VSUBS 0.007102f
C563 B.n523 VSUBS 0.007102f
C564 B.n524 VSUBS 0.007102f
C565 B.n525 VSUBS 0.007102f
C566 B.n526 VSUBS 0.007102f
C567 B.n527 VSUBS 0.007102f
C568 B.n528 VSUBS 0.007102f
C569 B.n529 VSUBS 0.007102f
C570 B.n530 VSUBS 0.007102f
C571 B.n531 VSUBS 0.007102f
C572 B.n532 VSUBS 0.007102f
C573 B.n533 VSUBS 0.007102f
C574 B.n534 VSUBS 0.017945f
C575 B.n535 VSUBS 0.016936f
C576 B.n536 VSUBS 0.016936f
C577 B.n537 VSUBS 0.007102f
C578 B.n538 VSUBS 0.007102f
C579 B.n539 VSUBS 0.007102f
C580 B.n540 VSUBS 0.007102f
C581 B.n541 VSUBS 0.007102f
C582 B.n542 VSUBS 0.007102f
C583 B.n543 VSUBS 0.007102f
C584 B.n544 VSUBS 0.007102f
C585 B.n545 VSUBS 0.007102f
C586 B.n546 VSUBS 0.007102f
C587 B.n547 VSUBS 0.007102f
C588 B.n548 VSUBS 0.007102f
C589 B.n549 VSUBS 0.007102f
C590 B.n550 VSUBS 0.007102f
C591 B.n551 VSUBS 0.007102f
C592 B.n552 VSUBS 0.007102f
C593 B.n553 VSUBS 0.007102f
C594 B.n554 VSUBS 0.007102f
C595 B.n555 VSUBS 0.007102f
C596 B.n556 VSUBS 0.007102f
C597 B.n557 VSUBS 0.007102f
C598 B.n558 VSUBS 0.007102f
C599 B.n559 VSUBS 0.007102f
C600 B.n560 VSUBS 0.007102f
C601 B.n561 VSUBS 0.007102f
C602 B.n562 VSUBS 0.007102f
C603 B.n563 VSUBS 0.007102f
C604 B.n564 VSUBS 0.007102f
C605 B.n565 VSUBS 0.007102f
C606 B.n566 VSUBS 0.007102f
C607 B.n567 VSUBS 0.007102f
C608 B.n568 VSUBS 0.007102f
C609 B.n569 VSUBS 0.007102f
C610 B.n570 VSUBS 0.007102f
C611 B.n571 VSUBS 0.007102f
C612 B.n572 VSUBS 0.007102f
C613 B.n573 VSUBS 0.007102f
C614 B.n574 VSUBS 0.007102f
C615 B.n575 VSUBS 0.007102f
C616 B.n576 VSUBS 0.007102f
C617 B.n577 VSUBS 0.007102f
C618 B.n578 VSUBS 0.007102f
C619 B.n579 VSUBS 0.007102f
C620 B.n580 VSUBS 0.007102f
C621 B.n581 VSUBS 0.007102f
C622 B.n582 VSUBS 0.007102f
C623 B.n583 VSUBS 0.007102f
C624 B.n584 VSUBS 0.007102f
C625 B.n585 VSUBS 0.007102f
C626 B.n586 VSUBS 0.007102f
C627 B.n587 VSUBS 0.007102f
C628 B.n588 VSUBS 0.007102f
C629 B.n589 VSUBS 0.007102f
C630 B.n590 VSUBS 0.007102f
C631 B.n591 VSUBS 0.007102f
C632 B.n592 VSUBS 0.007102f
C633 B.n593 VSUBS 0.007102f
C634 B.n594 VSUBS 0.007102f
C635 B.n595 VSUBS 0.007102f
C636 B.n596 VSUBS 0.007102f
C637 B.n597 VSUBS 0.007102f
C638 B.n598 VSUBS 0.007102f
C639 B.n599 VSUBS 0.007102f
C640 B.n600 VSUBS 0.007102f
C641 B.n601 VSUBS 0.007102f
C642 B.n602 VSUBS 0.007102f
C643 B.n603 VSUBS 0.007102f
C644 B.n604 VSUBS 0.007102f
C645 B.n605 VSUBS 0.007102f
C646 B.n606 VSUBS 0.007102f
C647 B.n607 VSUBS 0.007102f
C648 B.n608 VSUBS 0.007102f
C649 B.n609 VSUBS 0.007102f
C650 B.n610 VSUBS 0.007102f
C651 B.n611 VSUBS 0.007102f
C652 B.n612 VSUBS 0.007102f
C653 B.n613 VSUBS 0.007102f
C654 B.n614 VSUBS 0.007102f
C655 B.n615 VSUBS 0.007102f
C656 B.n616 VSUBS 0.007102f
C657 B.n617 VSUBS 0.007102f
C658 B.n618 VSUBS 0.007102f
C659 B.n619 VSUBS 0.007102f
C660 B.n620 VSUBS 0.007102f
C661 B.n621 VSUBS 0.007102f
C662 B.n622 VSUBS 0.007102f
C663 B.n623 VSUBS 0.007102f
C664 B.n624 VSUBS 0.007102f
C665 B.n625 VSUBS 0.007102f
C666 B.n626 VSUBS 0.007102f
C667 B.n627 VSUBS 0.007102f
C668 B.n628 VSUBS 0.007102f
C669 B.n629 VSUBS 0.007102f
C670 B.n630 VSUBS 0.007102f
C671 B.n631 VSUBS 0.007102f
C672 B.n632 VSUBS 0.007102f
C673 B.n633 VSUBS 0.007102f
C674 B.n634 VSUBS 0.007102f
C675 B.n635 VSUBS 0.007102f
C676 B.n636 VSUBS 0.007102f
C677 B.n637 VSUBS 0.007102f
C678 B.n638 VSUBS 0.007102f
C679 B.n639 VSUBS 0.007102f
C680 B.n640 VSUBS 0.007102f
C681 B.n641 VSUBS 0.007102f
C682 B.n642 VSUBS 0.007102f
C683 B.n643 VSUBS 0.007102f
C684 B.n644 VSUBS 0.007102f
C685 B.n645 VSUBS 0.007102f
C686 B.n646 VSUBS 0.007102f
C687 B.n647 VSUBS 0.007102f
C688 B.n648 VSUBS 0.007102f
C689 B.n649 VSUBS 0.007102f
C690 B.n650 VSUBS 0.007102f
C691 B.n651 VSUBS 0.007102f
C692 B.n652 VSUBS 0.007102f
C693 B.n653 VSUBS 0.007102f
C694 B.n654 VSUBS 0.007102f
C695 B.n655 VSUBS 0.007102f
C696 B.n656 VSUBS 0.007102f
C697 B.n657 VSUBS 0.007102f
C698 B.n658 VSUBS 0.007102f
C699 B.n659 VSUBS 0.007102f
C700 B.n660 VSUBS 0.007102f
C701 B.n661 VSUBS 0.007102f
C702 B.n662 VSUBS 0.007102f
C703 B.n663 VSUBS 0.007102f
C704 B.n664 VSUBS 0.007102f
C705 B.n665 VSUBS 0.007102f
C706 B.n666 VSUBS 0.007102f
C707 B.n667 VSUBS 0.007102f
C708 B.n668 VSUBS 0.007102f
C709 B.n669 VSUBS 0.007102f
C710 B.n670 VSUBS 0.007102f
C711 B.n671 VSUBS 0.007102f
C712 B.n672 VSUBS 0.007102f
C713 B.n673 VSUBS 0.007102f
C714 B.n674 VSUBS 0.007102f
C715 B.n675 VSUBS 0.007102f
C716 B.n676 VSUBS 0.007102f
C717 B.n677 VSUBS 0.007102f
C718 B.n678 VSUBS 0.007102f
C719 B.n679 VSUBS 0.007102f
C720 B.n680 VSUBS 0.007102f
C721 B.n681 VSUBS 0.007102f
C722 B.n682 VSUBS 0.007102f
C723 B.n683 VSUBS 0.007102f
C724 B.n684 VSUBS 0.007102f
C725 B.n685 VSUBS 0.007102f
C726 B.n686 VSUBS 0.007102f
C727 B.n687 VSUBS 0.007102f
C728 B.n688 VSUBS 0.007102f
C729 B.n689 VSUBS 0.007102f
C730 B.n690 VSUBS 0.007102f
C731 B.n691 VSUBS 0.007102f
C732 B.n692 VSUBS 0.007102f
C733 B.n693 VSUBS 0.007102f
C734 B.n694 VSUBS 0.007102f
C735 B.n695 VSUBS 0.007102f
C736 B.n696 VSUBS 0.007102f
C737 B.n697 VSUBS 0.017717f
C738 B.n698 VSUBS 0.016936f
C739 B.n699 VSUBS 0.017945f
C740 B.n700 VSUBS 0.007102f
C741 B.n701 VSUBS 0.007102f
C742 B.n702 VSUBS 0.007102f
C743 B.n703 VSUBS 0.007102f
C744 B.n704 VSUBS 0.007102f
C745 B.n705 VSUBS 0.007102f
C746 B.n706 VSUBS 0.007102f
C747 B.n707 VSUBS 0.007102f
C748 B.n708 VSUBS 0.007102f
C749 B.n709 VSUBS 0.007102f
C750 B.n710 VSUBS 0.007102f
C751 B.n711 VSUBS 0.007102f
C752 B.n712 VSUBS 0.007102f
C753 B.n713 VSUBS 0.007102f
C754 B.n714 VSUBS 0.007102f
C755 B.n715 VSUBS 0.007102f
C756 B.n716 VSUBS 0.007102f
C757 B.n717 VSUBS 0.007102f
C758 B.n718 VSUBS 0.007102f
C759 B.n719 VSUBS 0.007102f
C760 B.n720 VSUBS 0.007102f
C761 B.n721 VSUBS 0.007102f
C762 B.n722 VSUBS 0.007102f
C763 B.n723 VSUBS 0.007102f
C764 B.n724 VSUBS 0.007102f
C765 B.n725 VSUBS 0.007102f
C766 B.n726 VSUBS 0.007102f
C767 B.n727 VSUBS 0.007102f
C768 B.n728 VSUBS 0.007102f
C769 B.n729 VSUBS 0.007102f
C770 B.n730 VSUBS 0.007102f
C771 B.n731 VSUBS 0.007102f
C772 B.n732 VSUBS 0.007102f
C773 B.n733 VSUBS 0.007102f
C774 B.n734 VSUBS 0.007102f
C775 B.n735 VSUBS 0.007102f
C776 B.n736 VSUBS 0.007102f
C777 B.n737 VSUBS 0.007102f
C778 B.n738 VSUBS 0.007102f
C779 B.n739 VSUBS 0.007102f
C780 B.n740 VSUBS 0.007102f
C781 B.n741 VSUBS 0.007102f
C782 B.n742 VSUBS 0.007102f
C783 B.n743 VSUBS 0.007102f
C784 B.n744 VSUBS 0.007102f
C785 B.n745 VSUBS 0.007102f
C786 B.n746 VSUBS 0.007102f
C787 B.n747 VSUBS 0.007102f
C788 B.n748 VSUBS 0.007102f
C789 B.n749 VSUBS 0.007102f
C790 B.n750 VSUBS 0.007102f
C791 B.n751 VSUBS 0.007102f
C792 B.n752 VSUBS 0.007102f
C793 B.n753 VSUBS 0.007102f
C794 B.n754 VSUBS 0.007102f
C795 B.n755 VSUBS 0.007102f
C796 B.n756 VSUBS 0.007102f
C797 B.n757 VSUBS 0.007102f
C798 B.n758 VSUBS 0.007102f
C799 B.n759 VSUBS 0.007102f
C800 B.n760 VSUBS 0.007102f
C801 B.n761 VSUBS 0.007102f
C802 B.n762 VSUBS 0.007102f
C803 B.n763 VSUBS 0.007102f
C804 B.n764 VSUBS 0.007102f
C805 B.n765 VSUBS 0.007102f
C806 B.n766 VSUBS 0.007102f
C807 B.n767 VSUBS 0.007102f
C808 B.n768 VSUBS 0.007102f
C809 B.n769 VSUBS 0.007102f
C810 B.n770 VSUBS 0.007102f
C811 B.n771 VSUBS 0.007102f
C812 B.n772 VSUBS 0.007102f
C813 B.n773 VSUBS 0.007102f
C814 B.n774 VSUBS 0.007102f
C815 B.n775 VSUBS 0.007102f
C816 B.n776 VSUBS 0.007102f
C817 B.n777 VSUBS 0.007102f
C818 B.n778 VSUBS 0.007102f
C819 B.n779 VSUBS 0.007102f
C820 B.n780 VSUBS 0.007102f
C821 B.n781 VSUBS 0.007102f
C822 B.n782 VSUBS 0.007102f
C823 B.n783 VSUBS 0.007102f
C824 B.n784 VSUBS 0.007102f
C825 B.n785 VSUBS 0.007102f
C826 B.n786 VSUBS 0.007102f
C827 B.n787 VSUBS 0.007102f
C828 B.n788 VSUBS 0.007102f
C829 B.n789 VSUBS 0.007102f
C830 B.n790 VSUBS 0.007102f
C831 B.n791 VSUBS 0.006684f
C832 B.n792 VSUBS 0.016454f
C833 B.n793 VSUBS 0.003969f
C834 B.n794 VSUBS 0.007102f
C835 B.n795 VSUBS 0.007102f
C836 B.n796 VSUBS 0.007102f
C837 B.n797 VSUBS 0.007102f
C838 B.n798 VSUBS 0.007102f
C839 B.n799 VSUBS 0.007102f
C840 B.n800 VSUBS 0.007102f
C841 B.n801 VSUBS 0.007102f
C842 B.n802 VSUBS 0.007102f
C843 B.n803 VSUBS 0.007102f
C844 B.n804 VSUBS 0.007102f
C845 B.n805 VSUBS 0.007102f
C846 B.n806 VSUBS 0.003969f
C847 B.n807 VSUBS 0.007102f
C848 B.n808 VSUBS 0.007102f
C849 B.n809 VSUBS 0.006684f
C850 B.n810 VSUBS 0.007102f
C851 B.n811 VSUBS 0.007102f
C852 B.n812 VSUBS 0.007102f
C853 B.n813 VSUBS 0.007102f
C854 B.n814 VSUBS 0.007102f
C855 B.n815 VSUBS 0.007102f
C856 B.n816 VSUBS 0.007102f
C857 B.n817 VSUBS 0.007102f
C858 B.n818 VSUBS 0.007102f
C859 B.n819 VSUBS 0.007102f
C860 B.n820 VSUBS 0.007102f
C861 B.n821 VSUBS 0.007102f
C862 B.n822 VSUBS 0.007102f
C863 B.n823 VSUBS 0.007102f
C864 B.n824 VSUBS 0.007102f
C865 B.n825 VSUBS 0.007102f
C866 B.n826 VSUBS 0.007102f
C867 B.n827 VSUBS 0.007102f
C868 B.n828 VSUBS 0.007102f
C869 B.n829 VSUBS 0.007102f
C870 B.n830 VSUBS 0.007102f
C871 B.n831 VSUBS 0.007102f
C872 B.n832 VSUBS 0.007102f
C873 B.n833 VSUBS 0.007102f
C874 B.n834 VSUBS 0.007102f
C875 B.n835 VSUBS 0.007102f
C876 B.n836 VSUBS 0.007102f
C877 B.n837 VSUBS 0.007102f
C878 B.n838 VSUBS 0.007102f
C879 B.n839 VSUBS 0.007102f
C880 B.n840 VSUBS 0.007102f
C881 B.n841 VSUBS 0.007102f
C882 B.n842 VSUBS 0.007102f
C883 B.n843 VSUBS 0.007102f
C884 B.n844 VSUBS 0.007102f
C885 B.n845 VSUBS 0.007102f
C886 B.n846 VSUBS 0.007102f
C887 B.n847 VSUBS 0.007102f
C888 B.n848 VSUBS 0.007102f
C889 B.n849 VSUBS 0.007102f
C890 B.n850 VSUBS 0.007102f
C891 B.n851 VSUBS 0.007102f
C892 B.n852 VSUBS 0.007102f
C893 B.n853 VSUBS 0.007102f
C894 B.n854 VSUBS 0.007102f
C895 B.n855 VSUBS 0.007102f
C896 B.n856 VSUBS 0.007102f
C897 B.n857 VSUBS 0.007102f
C898 B.n858 VSUBS 0.007102f
C899 B.n859 VSUBS 0.007102f
C900 B.n860 VSUBS 0.007102f
C901 B.n861 VSUBS 0.007102f
C902 B.n862 VSUBS 0.007102f
C903 B.n863 VSUBS 0.007102f
C904 B.n864 VSUBS 0.007102f
C905 B.n865 VSUBS 0.007102f
C906 B.n866 VSUBS 0.007102f
C907 B.n867 VSUBS 0.007102f
C908 B.n868 VSUBS 0.007102f
C909 B.n869 VSUBS 0.007102f
C910 B.n870 VSUBS 0.007102f
C911 B.n871 VSUBS 0.007102f
C912 B.n872 VSUBS 0.007102f
C913 B.n873 VSUBS 0.007102f
C914 B.n874 VSUBS 0.007102f
C915 B.n875 VSUBS 0.007102f
C916 B.n876 VSUBS 0.007102f
C917 B.n877 VSUBS 0.007102f
C918 B.n878 VSUBS 0.007102f
C919 B.n879 VSUBS 0.007102f
C920 B.n880 VSUBS 0.007102f
C921 B.n881 VSUBS 0.007102f
C922 B.n882 VSUBS 0.007102f
C923 B.n883 VSUBS 0.007102f
C924 B.n884 VSUBS 0.007102f
C925 B.n885 VSUBS 0.007102f
C926 B.n886 VSUBS 0.007102f
C927 B.n887 VSUBS 0.007102f
C928 B.n888 VSUBS 0.007102f
C929 B.n889 VSUBS 0.007102f
C930 B.n890 VSUBS 0.007102f
C931 B.n891 VSUBS 0.007102f
C932 B.n892 VSUBS 0.007102f
C933 B.n893 VSUBS 0.007102f
C934 B.n894 VSUBS 0.007102f
C935 B.n895 VSUBS 0.007102f
C936 B.n896 VSUBS 0.007102f
C937 B.n897 VSUBS 0.007102f
C938 B.n898 VSUBS 0.007102f
C939 B.n899 VSUBS 0.007102f
C940 B.n900 VSUBS 0.017945f
C941 B.n901 VSUBS 0.016936f
C942 B.n902 VSUBS 0.016936f
C943 B.n903 VSUBS 0.007102f
C944 B.n904 VSUBS 0.007102f
C945 B.n905 VSUBS 0.007102f
C946 B.n906 VSUBS 0.007102f
C947 B.n907 VSUBS 0.007102f
C948 B.n908 VSUBS 0.007102f
C949 B.n909 VSUBS 0.007102f
C950 B.n910 VSUBS 0.007102f
C951 B.n911 VSUBS 0.007102f
C952 B.n912 VSUBS 0.007102f
C953 B.n913 VSUBS 0.007102f
C954 B.n914 VSUBS 0.007102f
C955 B.n915 VSUBS 0.007102f
C956 B.n916 VSUBS 0.007102f
C957 B.n917 VSUBS 0.007102f
C958 B.n918 VSUBS 0.007102f
C959 B.n919 VSUBS 0.007102f
C960 B.n920 VSUBS 0.007102f
C961 B.n921 VSUBS 0.007102f
C962 B.n922 VSUBS 0.007102f
C963 B.n923 VSUBS 0.007102f
C964 B.n924 VSUBS 0.007102f
C965 B.n925 VSUBS 0.007102f
C966 B.n926 VSUBS 0.007102f
C967 B.n927 VSUBS 0.007102f
C968 B.n928 VSUBS 0.007102f
C969 B.n929 VSUBS 0.007102f
C970 B.n930 VSUBS 0.007102f
C971 B.n931 VSUBS 0.007102f
C972 B.n932 VSUBS 0.007102f
C973 B.n933 VSUBS 0.007102f
C974 B.n934 VSUBS 0.007102f
C975 B.n935 VSUBS 0.007102f
C976 B.n936 VSUBS 0.007102f
C977 B.n937 VSUBS 0.007102f
C978 B.n938 VSUBS 0.007102f
C979 B.n939 VSUBS 0.007102f
C980 B.n940 VSUBS 0.007102f
C981 B.n941 VSUBS 0.007102f
C982 B.n942 VSUBS 0.007102f
C983 B.n943 VSUBS 0.007102f
C984 B.n944 VSUBS 0.007102f
C985 B.n945 VSUBS 0.007102f
C986 B.n946 VSUBS 0.007102f
C987 B.n947 VSUBS 0.007102f
C988 B.n948 VSUBS 0.007102f
C989 B.n949 VSUBS 0.007102f
C990 B.n950 VSUBS 0.007102f
C991 B.n951 VSUBS 0.007102f
C992 B.n952 VSUBS 0.007102f
C993 B.n953 VSUBS 0.007102f
C994 B.n954 VSUBS 0.007102f
C995 B.n955 VSUBS 0.007102f
C996 B.n956 VSUBS 0.007102f
C997 B.n957 VSUBS 0.007102f
C998 B.n958 VSUBS 0.007102f
C999 B.n959 VSUBS 0.007102f
C1000 B.n960 VSUBS 0.007102f
C1001 B.n961 VSUBS 0.007102f
C1002 B.n962 VSUBS 0.007102f
C1003 B.n963 VSUBS 0.007102f
C1004 B.n964 VSUBS 0.007102f
C1005 B.n965 VSUBS 0.007102f
C1006 B.n966 VSUBS 0.007102f
C1007 B.n967 VSUBS 0.007102f
C1008 B.n968 VSUBS 0.007102f
C1009 B.n969 VSUBS 0.007102f
C1010 B.n970 VSUBS 0.007102f
C1011 B.n971 VSUBS 0.007102f
C1012 B.n972 VSUBS 0.007102f
C1013 B.n973 VSUBS 0.007102f
C1014 B.n974 VSUBS 0.007102f
C1015 B.n975 VSUBS 0.007102f
C1016 B.n976 VSUBS 0.007102f
C1017 B.n977 VSUBS 0.007102f
C1018 B.n978 VSUBS 0.007102f
C1019 B.n979 VSUBS 0.007102f
C1020 B.n980 VSUBS 0.007102f
C1021 B.n981 VSUBS 0.007102f
C1022 B.n982 VSUBS 0.007102f
C1023 B.n983 VSUBS 0.016081f
C1024 VDD2.n0 VSUBS 0.030704f
C1025 VDD2.n1 VSUBS 0.027105f
C1026 VDD2.n2 VSUBS 0.014565f
C1027 VDD2.n3 VSUBS 0.034427f
C1028 VDD2.n4 VSUBS 0.015422f
C1029 VDD2.n5 VSUBS 0.027105f
C1030 VDD2.n6 VSUBS 0.014565f
C1031 VDD2.n7 VSUBS 0.034427f
C1032 VDD2.n8 VSUBS 0.015422f
C1033 VDD2.n9 VSUBS 0.027105f
C1034 VDD2.n10 VSUBS 0.014565f
C1035 VDD2.n11 VSUBS 0.034427f
C1036 VDD2.n12 VSUBS 0.015422f
C1037 VDD2.n13 VSUBS 0.027105f
C1038 VDD2.n14 VSUBS 0.014565f
C1039 VDD2.n15 VSUBS 0.034427f
C1040 VDD2.n16 VSUBS 0.015422f
C1041 VDD2.n17 VSUBS 0.027105f
C1042 VDD2.n18 VSUBS 0.014565f
C1043 VDD2.n19 VSUBS 0.034427f
C1044 VDD2.n20 VSUBS 0.015422f
C1045 VDD2.n21 VSUBS 0.027105f
C1046 VDD2.n22 VSUBS 0.014565f
C1047 VDD2.n23 VSUBS 0.034427f
C1048 VDD2.n24 VSUBS 0.015422f
C1049 VDD2.n25 VSUBS 0.027105f
C1050 VDD2.n26 VSUBS 0.014565f
C1051 VDD2.n27 VSUBS 0.034427f
C1052 VDD2.n28 VSUBS 0.015422f
C1053 VDD2.n29 VSUBS 0.027105f
C1054 VDD2.n30 VSUBS 0.014565f
C1055 VDD2.n31 VSUBS 0.034427f
C1056 VDD2.n32 VSUBS 0.015422f
C1057 VDD2.n33 VSUBS 0.223128f
C1058 VDD2.t4 VSUBS 0.073971f
C1059 VDD2.n34 VSUBS 0.02582f
C1060 VDD2.n35 VSUBS 0.021901f
C1061 VDD2.n36 VSUBS 0.014565f
C1062 VDD2.n37 VSUBS 2.22415f
C1063 VDD2.n38 VSUBS 0.027105f
C1064 VDD2.n39 VSUBS 0.014565f
C1065 VDD2.n40 VSUBS 0.015422f
C1066 VDD2.n41 VSUBS 0.034427f
C1067 VDD2.n42 VSUBS 0.034427f
C1068 VDD2.n43 VSUBS 0.015422f
C1069 VDD2.n44 VSUBS 0.014565f
C1070 VDD2.n45 VSUBS 0.027105f
C1071 VDD2.n46 VSUBS 0.027105f
C1072 VDD2.n47 VSUBS 0.014565f
C1073 VDD2.n48 VSUBS 0.015422f
C1074 VDD2.n49 VSUBS 0.034427f
C1075 VDD2.n50 VSUBS 0.034427f
C1076 VDD2.n51 VSUBS 0.015422f
C1077 VDD2.n52 VSUBS 0.014565f
C1078 VDD2.n53 VSUBS 0.027105f
C1079 VDD2.n54 VSUBS 0.027105f
C1080 VDD2.n55 VSUBS 0.014565f
C1081 VDD2.n56 VSUBS 0.015422f
C1082 VDD2.n57 VSUBS 0.034427f
C1083 VDD2.n58 VSUBS 0.034427f
C1084 VDD2.n59 VSUBS 0.015422f
C1085 VDD2.n60 VSUBS 0.014565f
C1086 VDD2.n61 VSUBS 0.027105f
C1087 VDD2.n62 VSUBS 0.027105f
C1088 VDD2.n63 VSUBS 0.014565f
C1089 VDD2.n64 VSUBS 0.015422f
C1090 VDD2.n65 VSUBS 0.034427f
C1091 VDD2.n66 VSUBS 0.034427f
C1092 VDD2.n67 VSUBS 0.015422f
C1093 VDD2.n68 VSUBS 0.014565f
C1094 VDD2.n69 VSUBS 0.027105f
C1095 VDD2.n70 VSUBS 0.027105f
C1096 VDD2.n71 VSUBS 0.014565f
C1097 VDD2.n72 VSUBS 0.015422f
C1098 VDD2.n73 VSUBS 0.034427f
C1099 VDD2.n74 VSUBS 0.034427f
C1100 VDD2.n75 VSUBS 0.034427f
C1101 VDD2.n76 VSUBS 0.015422f
C1102 VDD2.n77 VSUBS 0.014565f
C1103 VDD2.n78 VSUBS 0.027105f
C1104 VDD2.n79 VSUBS 0.027105f
C1105 VDD2.n80 VSUBS 0.014565f
C1106 VDD2.n81 VSUBS 0.014993f
C1107 VDD2.n82 VSUBS 0.014993f
C1108 VDD2.n83 VSUBS 0.034427f
C1109 VDD2.n84 VSUBS 0.034427f
C1110 VDD2.n85 VSUBS 0.015422f
C1111 VDD2.n86 VSUBS 0.014565f
C1112 VDD2.n87 VSUBS 0.027105f
C1113 VDD2.n88 VSUBS 0.027105f
C1114 VDD2.n89 VSUBS 0.014565f
C1115 VDD2.n90 VSUBS 0.015422f
C1116 VDD2.n91 VSUBS 0.034427f
C1117 VDD2.n92 VSUBS 0.034427f
C1118 VDD2.n93 VSUBS 0.015422f
C1119 VDD2.n94 VSUBS 0.014565f
C1120 VDD2.n95 VSUBS 0.027105f
C1121 VDD2.n96 VSUBS 0.027105f
C1122 VDD2.n97 VSUBS 0.014565f
C1123 VDD2.n98 VSUBS 0.015422f
C1124 VDD2.n99 VSUBS 0.034427f
C1125 VDD2.n100 VSUBS 0.08648f
C1126 VDD2.n101 VSUBS 0.015422f
C1127 VDD2.n102 VSUBS 0.014565f
C1128 VDD2.n103 VSUBS 0.064504f
C1129 VDD2.n104 VSUBS 0.075184f
C1130 VDD2.t1 VSUBS 0.407182f
C1131 VDD2.t0 VSUBS 0.407182f
C1132 VDD2.n105 VSUBS 3.41872f
C1133 VDD2.n106 VSUBS 4.15453f
C1134 VDD2.n107 VSUBS 0.030704f
C1135 VDD2.n108 VSUBS 0.027105f
C1136 VDD2.n109 VSUBS 0.014565f
C1137 VDD2.n110 VSUBS 0.034427f
C1138 VDD2.n111 VSUBS 0.015422f
C1139 VDD2.n112 VSUBS 0.027105f
C1140 VDD2.n113 VSUBS 0.014565f
C1141 VDD2.n114 VSUBS 0.034427f
C1142 VDD2.n115 VSUBS 0.015422f
C1143 VDD2.n116 VSUBS 0.027105f
C1144 VDD2.n117 VSUBS 0.014565f
C1145 VDD2.n118 VSUBS 0.034427f
C1146 VDD2.n119 VSUBS 0.015422f
C1147 VDD2.n120 VSUBS 0.027105f
C1148 VDD2.n121 VSUBS 0.014565f
C1149 VDD2.n122 VSUBS 0.034427f
C1150 VDD2.n123 VSUBS 0.034427f
C1151 VDD2.n124 VSUBS 0.015422f
C1152 VDD2.n125 VSUBS 0.027105f
C1153 VDD2.n126 VSUBS 0.014565f
C1154 VDD2.n127 VSUBS 0.034427f
C1155 VDD2.n128 VSUBS 0.015422f
C1156 VDD2.n129 VSUBS 0.027105f
C1157 VDD2.n130 VSUBS 0.014565f
C1158 VDD2.n131 VSUBS 0.034427f
C1159 VDD2.n132 VSUBS 0.015422f
C1160 VDD2.n133 VSUBS 0.027105f
C1161 VDD2.n134 VSUBS 0.014565f
C1162 VDD2.n135 VSUBS 0.034427f
C1163 VDD2.n136 VSUBS 0.015422f
C1164 VDD2.n137 VSUBS 0.027105f
C1165 VDD2.n138 VSUBS 0.014565f
C1166 VDD2.n139 VSUBS 0.034427f
C1167 VDD2.n140 VSUBS 0.015422f
C1168 VDD2.n141 VSUBS 0.223128f
C1169 VDD2.t5 VSUBS 0.073971f
C1170 VDD2.n142 VSUBS 0.02582f
C1171 VDD2.n143 VSUBS 0.021901f
C1172 VDD2.n144 VSUBS 0.014565f
C1173 VDD2.n145 VSUBS 2.22415f
C1174 VDD2.n146 VSUBS 0.027105f
C1175 VDD2.n147 VSUBS 0.014565f
C1176 VDD2.n148 VSUBS 0.015422f
C1177 VDD2.n149 VSUBS 0.034427f
C1178 VDD2.n150 VSUBS 0.034427f
C1179 VDD2.n151 VSUBS 0.015422f
C1180 VDD2.n152 VSUBS 0.014565f
C1181 VDD2.n153 VSUBS 0.027105f
C1182 VDD2.n154 VSUBS 0.027105f
C1183 VDD2.n155 VSUBS 0.014565f
C1184 VDD2.n156 VSUBS 0.015422f
C1185 VDD2.n157 VSUBS 0.034427f
C1186 VDD2.n158 VSUBS 0.034427f
C1187 VDD2.n159 VSUBS 0.015422f
C1188 VDD2.n160 VSUBS 0.014565f
C1189 VDD2.n161 VSUBS 0.027105f
C1190 VDD2.n162 VSUBS 0.027105f
C1191 VDD2.n163 VSUBS 0.014565f
C1192 VDD2.n164 VSUBS 0.015422f
C1193 VDD2.n165 VSUBS 0.034427f
C1194 VDD2.n166 VSUBS 0.034427f
C1195 VDD2.n167 VSUBS 0.015422f
C1196 VDD2.n168 VSUBS 0.014565f
C1197 VDD2.n169 VSUBS 0.027105f
C1198 VDD2.n170 VSUBS 0.027105f
C1199 VDD2.n171 VSUBS 0.014565f
C1200 VDD2.n172 VSUBS 0.015422f
C1201 VDD2.n173 VSUBS 0.034427f
C1202 VDD2.n174 VSUBS 0.034427f
C1203 VDD2.n175 VSUBS 0.015422f
C1204 VDD2.n176 VSUBS 0.014565f
C1205 VDD2.n177 VSUBS 0.027105f
C1206 VDD2.n178 VSUBS 0.027105f
C1207 VDD2.n179 VSUBS 0.014565f
C1208 VDD2.n180 VSUBS 0.015422f
C1209 VDD2.n181 VSUBS 0.034427f
C1210 VDD2.n182 VSUBS 0.034427f
C1211 VDD2.n183 VSUBS 0.015422f
C1212 VDD2.n184 VSUBS 0.014565f
C1213 VDD2.n185 VSUBS 0.027105f
C1214 VDD2.n186 VSUBS 0.027105f
C1215 VDD2.n187 VSUBS 0.014565f
C1216 VDD2.n188 VSUBS 0.014993f
C1217 VDD2.n189 VSUBS 0.014993f
C1218 VDD2.n190 VSUBS 0.034427f
C1219 VDD2.n191 VSUBS 0.034427f
C1220 VDD2.n192 VSUBS 0.015422f
C1221 VDD2.n193 VSUBS 0.014565f
C1222 VDD2.n194 VSUBS 0.027105f
C1223 VDD2.n195 VSUBS 0.027105f
C1224 VDD2.n196 VSUBS 0.014565f
C1225 VDD2.n197 VSUBS 0.015422f
C1226 VDD2.n198 VSUBS 0.034427f
C1227 VDD2.n199 VSUBS 0.034427f
C1228 VDD2.n200 VSUBS 0.015422f
C1229 VDD2.n201 VSUBS 0.014565f
C1230 VDD2.n202 VSUBS 0.027105f
C1231 VDD2.n203 VSUBS 0.027105f
C1232 VDD2.n204 VSUBS 0.014565f
C1233 VDD2.n205 VSUBS 0.015422f
C1234 VDD2.n206 VSUBS 0.034427f
C1235 VDD2.n207 VSUBS 0.08648f
C1236 VDD2.n208 VSUBS 0.015422f
C1237 VDD2.n209 VSUBS 0.014565f
C1238 VDD2.n210 VSUBS 0.064504f
C1239 VDD2.n211 VSUBS 0.062387f
C1240 VDD2.n212 VSUBS 3.64889f
C1241 VDD2.t3 VSUBS 0.407182f
C1242 VDD2.t2 VSUBS 0.407182f
C1243 VDD2.n213 VSUBS 3.41866f
C1244 VN.t5 VSUBS 4.18329f
C1245 VN.n0 VSUBS 1.52554f
C1246 VN.n1 VSUBS 0.022263f
C1247 VN.n2 VSUBS 0.034981f
C1248 VN.n3 VSUBS 0.022263f
C1249 VN.n4 VSUBS 0.03125f
C1250 VN.t4 VSUBS 4.18329f
C1251 VN.n5 VSUBS 1.51702f
C1252 VN.t1 VSUBS 4.51463f
C1253 VN.n6 VSUBS 1.45148f
C1254 VN.n7 VSUBS 0.278146f
C1255 VN.n8 VSUBS 0.022263f
C1256 VN.n9 VSUBS 0.041493f
C1257 VN.n10 VSUBS 0.041493f
C1258 VN.n11 VSUBS 0.030018f
C1259 VN.n12 VSUBS 0.022263f
C1260 VN.n13 VSUBS 0.022263f
C1261 VN.n14 VSUBS 0.022263f
C1262 VN.n15 VSUBS 0.041493f
C1263 VN.n16 VSUBS 0.041493f
C1264 VN.n17 VSUBS 0.027972f
C1265 VN.n18 VSUBS 0.035932f
C1266 VN.n19 VSUBS 0.062073f
C1267 VN.t0 VSUBS 4.18329f
C1268 VN.n20 VSUBS 1.52554f
C1269 VN.n21 VSUBS 0.022263f
C1270 VN.n22 VSUBS 0.034981f
C1271 VN.n23 VSUBS 0.022263f
C1272 VN.n24 VSUBS 0.03125f
C1273 VN.t3 VSUBS 4.51463f
C1274 VN.t2 VSUBS 4.18329f
C1275 VN.n25 VSUBS 1.51702f
C1276 VN.n26 VSUBS 1.45148f
C1277 VN.n27 VSUBS 0.278146f
C1278 VN.n28 VSUBS 0.022263f
C1279 VN.n29 VSUBS 0.041493f
C1280 VN.n30 VSUBS 0.041493f
C1281 VN.n31 VSUBS 0.030018f
C1282 VN.n32 VSUBS 0.022263f
C1283 VN.n33 VSUBS 0.022263f
C1284 VN.n34 VSUBS 0.022263f
C1285 VN.n35 VSUBS 0.041493f
C1286 VN.n36 VSUBS 0.041493f
C1287 VN.n37 VSUBS 0.027972f
C1288 VN.n38 VSUBS 0.035932f
C1289 VN.n39 VSUBS 1.57301f
C1290 VTAIL.t0 VSUBS 0.419659f
C1291 VTAIL.t3 VSUBS 0.419659f
C1292 VTAIL.n0 VSUBS 3.34004f
C1293 VTAIL.n1 VSUBS 0.961864f
C1294 VTAIL.n2 VSUBS 0.031644f
C1295 VTAIL.n3 VSUBS 0.027936f
C1296 VTAIL.n4 VSUBS 0.015011f
C1297 VTAIL.n5 VSUBS 0.035482f
C1298 VTAIL.n6 VSUBS 0.015895f
C1299 VTAIL.n7 VSUBS 0.027936f
C1300 VTAIL.n8 VSUBS 0.015011f
C1301 VTAIL.n9 VSUBS 0.035482f
C1302 VTAIL.n10 VSUBS 0.015895f
C1303 VTAIL.n11 VSUBS 0.027936f
C1304 VTAIL.n12 VSUBS 0.015011f
C1305 VTAIL.n13 VSUBS 0.035482f
C1306 VTAIL.n14 VSUBS 0.015895f
C1307 VTAIL.n15 VSUBS 0.027936f
C1308 VTAIL.n16 VSUBS 0.015011f
C1309 VTAIL.n17 VSUBS 0.035482f
C1310 VTAIL.n18 VSUBS 0.015895f
C1311 VTAIL.n19 VSUBS 0.027936f
C1312 VTAIL.n20 VSUBS 0.015011f
C1313 VTAIL.n21 VSUBS 0.035482f
C1314 VTAIL.n22 VSUBS 0.015895f
C1315 VTAIL.n23 VSUBS 0.027936f
C1316 VTAIL.n24 VSUBS 0.015011f
C1317 VTAIL.n25 VSUBS 0.035482f
C1318 VTAIL.n26 VSUBS 0.015895f
C1319 VTAIL.n27 VSUBS 0.027936f
C1320 VTAIL.n28 VSUBS 0.015011f
C1321 VTAIL.n29 VSUBS 0.035482f
C1322 VTAIL.n30 VSUBS 0.015895f
C1323 VTAIL.n31 VSUBS 0.027936f
C1324 VTAIL.n32 VSUBS 0.015011f
C1325 VTAIL.n33 VSUBS 0.035482f
C1326 VTAIL.n34 VSUBS 0.015895f
C1327 VTAIL.n35 VSUBS 0.229965f
C1328 VTAIL.t8 VSUBS 0.076238f
C1329 VTAIL.n36 VSUBS 0.026611f
C1330 VTAIL.n37 VSUBS 0.022572f
C1331 VTAIL.n38 VSUBS 0.015011f
C1332 VTAIL.n39 VSUBS 2.29231f
C1333 VTAIL.n40 VSUBS 0.027936f
C1334 VTAIL.n41 VSUBS 0.015011f
C1335 VTAIL.n42 VSUBS 0.015895f
C1336 VTAIL.n43 VSUBS 0.035482f
C1337 VTAIL.n44 VSUBS 0.035482f
C1338 VTAIL.n45 VSUBS 0.015895f
C1339 VTAIL.n46 VSUBS 0.015011f
C1340 VTAIL.n47 VSUBS 0.027936f
C1341 VTAIL.n48 VSUBS 0.027936f
C1342 VTAIL.n49 VSUBS 0.015011f
C1343 VTAIL.n50 VSUBS 0.015895f
C1344 VTAIL.n51 VSUBS 0.035482f
C1345 VTAIL.n52 VSUBS 0.035482f
C1346 VTAIL.n53 VSUBS 0.015895f
C1347 VTAIL.n54 VSUBS 0.015011f
C1348 VTAIL.n55 VSUBS 0.027936f
C1349 VTAIL.n56 VSUBS 0.027936f
C1350 VTAIL.n57 VSUBS 0.015011f
C1351 VTAIL.n58 VSUBS 0.015895f
C1352 VTAIL.n59 VSUBS 0.035482f
C1353 VTAIL.n60 VSUBS 0.035482f
C1354 VTAIL.n61 VSUBS 0.015895f
C1355 VTAIL.n62 VSUBS 0.015011f
C1356 VTAIL.n63 VSUBS 0.027936f
C1357 VTAIL.n64 VSUBS 0.027936f
C1358 VTAIL.n65 VSUBS 0.015011f
C1359 VTAIL.n66 VSUBS 0.015895f
C1360 VTAIL.n67 VSUBS 0.035482f
C1361 VTAIL.n68 VSUBS 0.035482f
C1362 VTAIL.n69 VSUBS 0.015895f
C1363 VTAIL.n70 VSUBS 0.015011f
C1364 VTAIL.n71 VSUBS 0.027936f
C1365 VTAIL.n72 VSUBS 0.027936f
C1366 VTAIL.n73 VSUBS 0.015011f
C1367 VTAIL.n74 VSUBS 0.015895f
C1368 VTAIL.n75 VSUBS 0.035482f
C1369 VTAIL.n76 VSUBS 0.035482f
C1370 VTAIL.n77 VSUBS 0.035482f
C1371 VTAIL.n78 VSUBS 0.015895f
C1372 VTAIL.n79 VSUBS 0.015011f
C1373 VTAIL.n80 VSUBS 0.027936f
C1374 VTAIL.n81 VSUBS 0.027936f
C1375 VTAIL.n82 VSUBS 0.015011f
C1376 VTAIL.n83 VSUBS 0.015453f
C1377 VTAIL.n84 VSUBS 0.015453f
C1378 VTAIL.n85 VSUBS 0.035482f
C1379 VTAIL.n86 VSUBS 0.035482f
C1380 VTAIL.n87 VSUBS 0.015895f
C1381 VTAIL.n88 VSUBS 0.015011f
C1382 VTAIL.n89 VSUBS 0.027936f
C1383 VTAIL.n90 VSUBS 0.027936f
C1384 VTAIL.n91 VSUBS 0.015011f
C1385 VTAIL.n92 VSUBS 0.015895f
C1386 VTAIL.n93 VSUBS 0.035482f
C1387 VTAIL.n94 VSUBS 0.035482f
C1388 VTAIL.n95 VSUBS 0.015895f
C1389 VTAIL.n96 VSUBS 0.015011f
C1390 VTAIL.n97 VSUBS 0.027936f
C1391 VTAIL.n98 VSUBS 0.027936f
C1392 VTAIL.n99 VSUBS 0.015011f
C1393 VTAIL.n100 VSUBS 0.015895f
C1394 VTAIL.n101 VSUBS 0.035482f
C1395 VTAIL.n102 VSUBS 0.08913f
C1396 VTAIL.n103 VSUBS 0.015895f
C1397 VTAIL.n104 VSUBS 0.015011f
C1398 VTAIL.n105 VSUBS 0.06648f
C1399 VTAIL.n106 VSUBS 0.045024f
C1400 VTAIL.n107 VSUBS 0.523513f
C1401 VTAIL.t4 VSUBS 0.419659f
C1402 VTAIL.t5 VSUBS 0.419659f
C1403 VTAIL.n108 VSUBS 3.34004f
C1404 VTAIL.n109 VSUBS 3.4534f
C1405 VTAIL.t10 VSUBS 0.419659f
C1406 VTAIL.t11 VSUBS 0.419659f
C1407 VTAIL.n110 VSUBS 3.34005f
C1408 VTAIL.n111 VSUBS 3.45339f
C1409 VTAIL.n112 VSUBS 0.031644f
C1410 VTAIL.n113 VSUBS 0.027936f
C1411 VTAIL.n114 VSUBS 0.015011f
C1412 VTAIL.n115 VSUBS 0.035482f
C1413 VTAIL.n116 VSUBS 0.015895f
C1414 VTAIL.n117 VSUBS 0.027936f
C1415 VTAIL.n118 VSUBS 0.015011f
C1416 VTAIL.n119 VSUBS 0.035482f
C1417 VTAIL.n120 VSUBS 0.015895f
C1418 VTAIL.n121 VSUBS 0.027936f
C1419 VTAIL.n122 VSUBS 0.015011f
C1420 VTAIL.n123 VSUBS 0.035482f
C1421 VTAIL.n124 VSUBS 0.015895f
C1422 VTAIL.n125 VSUBS 0.027936f
C1423 VTAIL.n126 VSUBS 0.015011f
C1424 VTAIL.n127 VSUBS 0.035482f
C1425 VTAIL.n128 VSUBS 0.035482f
C1426 VTAIL.n129 VSUBS 0.015895f
C1427 VTAIL.n130 VSUBS 0.027936f
C1428 VTAIL.n131 VSUBS 0.015011f
C1429 VTAIL.n132 VSUBS 0.035482f
C1430 VTAIL.n133 VSUBS 0.015895f
C1431 VTAIL.n134 VSUBS 0.027936f
C1432 VTAIL.n135 VSUBS 0.015011f
C1433 VTAIL.n136 VSUBS 0.035482f
C1434 VTAIL.n137 VSUBS 0.015895f
C1435 VTAIL.n138 VSUBS 0.027936f
C1436 VTAIL.n139 VSUBS 0.015011f
C1437 VTAIL.n140 VSUBS 0.035482f
C1438 VTAIL.n141 VSUBS 0.015895f
C1439 VTAIL.n142 VSUBS 0.027936f
C1440 VTAIL.n143 VSUBS 0.015011f
C1441 VTAIL.n144 VSUBS 0.035482f
C1442 VTAIL.n145 VSUBS 0.015895f
C1443 VTAIL.n146 VSUBS 0.229965f
C1444 VTAIL.t1 VSUBS 0.076238f
C1445 VTAIL.n147 VSUBS 0.026611f
C1446 VTAIL.n148 VSUBS 0.022572f
C1447 VTAIL.n149 VSUBS 0.015011f
C1448 VTAIL.n150 VSUBS 2.29231f
C1449 VTAIL.n151 VSUBS 0.027936f
C1450 VTAIL.n152 VSUBS 0.015011f
C1451 VTAIL.n153 VSUBS 0.015895f
C1452 VTAIL.n154 VSUBS 0.035482f
C1453 VTAIL.n155 VSUBS 0.035482f
C1454 VTAIL.n156 VSUBS 0.015895f
C1455 VTAIL.n157 VSUBS 0.015011f
C1456 VTAIL.n158 VSUBS 0.027936f
C1457 VTAIL.n159 VSUBS 0.027936f
C1458 VTAIL.n160 VSUBS 0.015011f
C1459 VTAIL.n161 VSUBS 0.015895f
C1460 VTAIL.n162 VSUBS 0.035482f
C1461 VTAIL.n163 VSUBS 0.035482f
C1462 VTAIL.n164 VSUBS 0.015895f
C1463 VTAIL.n165 VSUBS 0.015011f
C1464 VTAIL.n166 VSUBS 0.027936f
C1465 VTAIL.n167 VSUBS 0.027936f
C1466 VTAIL.n168 VSUBS 0.015011f
C1467 VTAIL.n169 VSUBS 0.015895f
C1468 VTAIL.n170 VSUBS 0.035482f
C1469 VTAIL.n171 VSUBS 0.035482f
C1470 VTAIL.n172 VSUBS 0.015895f
C1471 VTAIL.n173 VSUBS 0.015011f
C1472 VTAIL.n174 VSUBS 0.027936f
C1473 VTAIL.n175 VSUBS 0.027936f
C1474 VTAIL.n176 VSUBS 0.015011f
C1475 VTAIL.n177 VSUBS 0.015895f
C1476 VTAIL.n178 VSUBS 0.035482f
C1477 VTAIL.n179 VSUBS 0.035482f
C1478 VTAIL.n180 VSUBS 0.015895f
C1479 VTAIL.n181 VSUBS 0.015011f
C1480 VTAIL.n182 VSUBS 0.027936f
C1481 VTAIL.n183 VSUBS 0.027936f
C1482 VTAIL.n184 VSUBS 0.015011f
C1483 VTAIL.n185 VSUBS 0.015895f
C1484 VTAIL.n186 VSUBS 0.035482f
C1485 VTAIL.n187 VSUBS 0.035482f
C1486 VTAIL.n188 VSUBS 0.015895f
C1487 VTAIL.n189 VSUBS 0.015011f
C1488 VTAIL.n190 VSUBS 0.027936f
C1489 VTAIL.n191 VSUBS 0.027936f
C1490 VTAIL.n192 VSUBS 0.015011f
C1491 VTAIL.n193 VSUBS 0.015453f
C1492 VTAIL.n194 VSUBS 0.015453f
C1493 VTAIL.n195 VSUBS 0.035482f
C1494 VTAIL.n196 VSUBS 0.035482f
C1495 VTAIL.n197 VSUBS 0.015895f
C1496 VTAIL.n198 VSUBS 0.015011f
C1497 VTAIL.n199 VSUBS 0.027936f
C1498 VTAIL.n200 VSUBS 0.027936f
C1499 VTAIL.n201 VSUBS 0.015011f
C1500 VTAIL.n202 VSUBS 0.015895f
C1501 VTAIL.n203 VSUBS 0.035482f
C1502 VTAIL.n204 VSUBS 0.035482f
C1503 VTAIL.n205 VSUBS 0.015895f
C1504 VTAIL.n206 VSUBS 0.015011f
C1505 VTAIL.n207 VSUBS 0.027936f
C1506 VTAIL.n208 VSUBS 0.027936f
C1507 VTAIL.n209 VSUBS 0.015011f
C1508 VTAIL.n210 VSUBS 0.015895f
C1509 VTAIL.n211 VSUBS 0.035482f
C1510 VTAIL.n212 VSUBS 0.08913f
C1511 VTAIL.n213 VSUBS 0.015895f
C1512 VTAIL.n214 VSUBS 0.015011f
C1513 VTAIL.n215 VSUBS 0.06648f
C1514 VTAIL.n216 VSUBS 0.045024f
C1515 VTAIL.n217 VSUBS 0.523513f
C1516 VTAIL.t7 VSUBS 0.419659f
C1517 VTAIL.t9 VSUBS 0.419659f
C1518 VTAIL.n218 VSUBS 3.34005f
C1519 VTAIL.n219 VSUBS 1.18476f
C1520 VTAIL.n220 VSUBS 0.031644f
C1521 VTAIL.n221 VSUBS 0.027936f
C1522 VTAIL.n222 VSUBS 0.015011f
C1523 VTAIL.n223 VSUBS 0.035482f
C1524 VTAIL.n224 VSUBS 0.015895f
C1525 VTAIL.n225 VSUBS 0.027936f
C1526 VTAIL.n226 VSUBS 0.015011f
C1527 VTAIL.n227 VSUBS 0.035482f
C1528 VTAIL.n228 VSUBS 0.015895f
C1529 VTAIL.n229 VSUBS 0.027936f
C1530 VTAIL.n230 VSUBS 0.015011f
C1531 VTAIL.n231 VSUBS 0.035482f
C1532 VTAIL.n232 VSUBS 0.015895f
C1533 VTAIL.n233 VSUBS 0.027936f
C1534 VTAIL.n234 VSUBS 0.015011f
C1535 VTAIL.n235 VSUBS 0.035482f
C1536 VTAIL.n236 VSUBS 0.035482f
C1537 VTAIL.n237 VSUBS 0.015895f
C1538 VTAIL.n238 VSUBS 0.027936f
C1539 VTAIL.n239 VSUBS 0.015011f
C1540 VTAIL.n240 VSUBS 0.035482f
C1541 VTAIL.n241 VSUBS 0.015895f
C1542 VTAIL.n242 VSUBS 0.027936f
C1543 VTAIL.n243 VSUBS 0.015011f
C1544 VTAIL.n244 VSUBS 0.035482f
C1545 VTAIL.n245 VSUBS 0.015895f
C1546 VTAIL.n246 VSUBS 0.027936f
C1547 VTAIL.n247 VSUBS 0.015011f
C1548 VTAIL.n248 VSUBS 0.035482f
C1549 VTAIL.n249 VSUBS 0.015895f
C1550 VTAIL.n250 VSUBS 0.027936f
C1551 VTAIL.n251 VSUBS 0.015011f
C1552 VTAIL.n252 VSUBS 0.035482f
C1553 VTAIL.n253 VSUBS 0.015895f
C1554 VTAIL.n254 VSUBS 0.229965f
C1555 VTAIL.t6 VSUBS 0.076238f
C1556 VTAIL.n255 VSUBS 0.026611f
C1557 VTAIL.n256 VSUBS 0.022572f
C1558 VTAIL.n257 VSUBS 0.015011f
C1559 VTAIL.n258 VSUBS 2.29231f
C1560 VTAIL.n259 VSUBS 0.027936f
C1561 VTAIL.n260 VSUBS 0.015011f
C1562 VTAIL.n261 VSUBS 0.015895f
C1563 VTAIL.n262 VSUBS 0.035482f
C1564 VTAIL.n263 VSUBS 0.035482f
C1565 VTAIL.n264 VSUBS 0.015895f
C1566 VTAIL.n265 VSUBS 0.015011f
C1567 VTAIL.n266 VSUBS 0.027936f
C1568 VTAIL.n267 VSUBS 0.027936f
C1569 VTAIL.n268 VSUBS 0.015011f
C1570 VTAIL.n269 VSUBS 0.015895f
C1571 VTAIL.n270 VSUBS 0.035482f
C1572 VTAIL.n271 VSUBS 0.035482f
C1573 VTAIL.n272 VSUBS 0.015895f
C1574 VTAIL.n273 VSUBS 0.015011f
C1575 VTAIL.n274 VSUBS 0.027936f
C1576 VTAIL.n275 VSUBS 0.027936f
C1577 VTAIL.n276 VSUBS 0.015011f
C1578 VTAIL.n277 VSUBS 0.015895f
C1579 VTAIL.n278 VSUBS 0.035482f
C1580 VTAIL.n279 VSUBS 0.035482f
C1581 VTAIL.n280 VSUBS 0.015895f
C1582 VTAIL.n281 VSUBS 0.015011f
C1583 VTAIL.n282 VSUBS 0.027936f
C1584 VTAIL.n283 VSUBS 0.027936f
C1585 VTAIL.n284 VSUBS 0.015011f
C1586 VTAIL.n285 VSUBS 0.015895f
C1587 VTAIL.n286 VSUBS 0.035482f
C1588 VTAIL.n287 VSUBS 0.035482f
C1589 VTAIL.n288 VSUBS 0.015895f
C1590 VTAIL.n289 VSUBS 0.015011f
C1591 VTAIL.n290 VSUBS 0.027936f
C1592 VTAIL.n291 VSUBS 0.027936f
C1593 VTAIL.n292 VSUBS 0.015011f
C1594 VTAIL.n293 VSUBS 0.015895f
C1595 VTAIL.n294 VSUBS 0.035482f
C1596 VTAIL.n295 VSUBS 0.035482f
C1597 VTAIL.n296 VSUBS 0.015895f
C1598 VTAIL.n297 VSUBS 0.015011f
C1599 VTAIL.n298 VSUBS 0.027936f
C1600 VTAIL.n299 VSUBS 0.027936f
C1601 VTAIL.n300 VSUBS 0.015011f
C1602 VTAIL.n301 VSUBS 0.015453f
C1603 VTAIL.n302 VSUBS 0.015453f
C1604 VTAIL.n303 VSUBS 0.035482f
C1605 VTAIL.n304 VSUBS 0.035482f
C1606 VTAIL.n305 VSUBS 0.015895f
C1607 VTAIL.n306 VSUBS 0.015011f
C1608 VTAIL.n307 VSUBS 0.027936f
C1609 VTAIL.n308 VSUBS 0.027936f
C1610 VTAIL.n309 VSUBS 0.015011f
C1611 VTAIL.n310 VSUBS 0.015895f
C1612 VTAIL.n311 VSUBS 0.035482f
C1613 VTAIL.n312 VSUBS 0.035482f
C1614 VTAIL.n313 VSUBS 0.015895f
C1615 VTAIL.n314 VSUBS 0.015011f
C1616 VTAIL.n315 VSUBS 0.027936f
C1617 VTAIL.n316 VSUBS 0.027936f
C1618 VTAIL.n317 VSUBS 0.015011f
C1619 VTAIL.n318 VSUBS 0.015895f
C1620 VTAIL.n319 VSUBS 0.035482f
C1621 VTAIL.n320 VSUBS 0.08913f
C1622 VTAIL.n321 VSUBS 0.015895f
C1623 VTAIL.n322 VSUBS 0.015011f
C1624 VTAIL.n323 VSUBS 0.06648f
C1625 VTAIL.n324 VSUBS 0.045024f
C1626 VTAIL.n325 VSUBS 2.48796f
C1627 VTAIL.n326 VSUBS 0.031644f
C1628 VTAIL.n327 VSUBS 0.027936f
C1629 VTAIL.n328 VSUBS 0.015011f
C1630 VTAIL.n329 VSUBS 0.035482f
C1631 VTAIL.n330 VSUBS 0.015895f
C1632 VTAIL.n331 VSUBS 0.027936f
C1633 VTAIL.n332 VSUBS 0.015011f
C1634 VTAIL.n333 VSUBS 0.035482f
C1635 VTAIL.n334 VSUBS 0.015895f
C1636 VTAIL.n335 VSUBS 0.027936f
C1637 VTAIL.n336 VSUBS 0.015011f
C1638 VTAIL.n337 VSUBS 0.035482f
C1639 VTAIL.n338 VSUBS 0.015895f
C1640 VTAIL.n339 VSUBS 0.027936f
C1641 VTAIL.n340 VSUBS 0.015011f
C1642 VTAIL.n341 VSUBS 0.035482f
C1643 VTAIL.n342 VSUBS 0.015895f
C1644 VTAIL.n343 VSUBS 0.027936f
C1645 VTAIL.n344 VSUBS 0.015011f
C1646 VTAIL.n345 VSUBS 0.035482f
C1647 VTAIL.n346 VSUBS 0.015895f
C1648 VTAIL.n347 VSUBS 0.027936f
C1649 VTAIL.n348 VSUBS 0.015011f
C1650 VTAIL.n349 VSUBS 0.035482f
C1651 VTAIL.n350 VSUBS 0.015895f
C1652 VTAIL.n351 VSUBS 0.027936f
C1653 VTAIL.n352 VSUBS 0.015011f
C1654 VTAIL.n353 VSUBS 0.035482f
C1655 VTAIL.n354 VSUBS 0.015895f
C1656 VTAIL.n355 VSUBS 0.027936f
C1657 VTAIL.n356 VSUBS 0.015011f
C1658 VTAIL.n357 VSUBS 0.035482f
C1659 VTAIL.n358 VSUBS 0.015895f
C1660 VTAIL.n359 VSUBS 0.229965f
C1661 VTAIL.t2 VSUBS 0.076238f
C1662 VTAIL.n360 VSUBS 0.026611f
C1663 VTAIL.n361 VSUBS 0.022572f
C1664 VTAIL.n362 VSUBS 0.015011f
C1665 VTAIL.n363 VSUBS 2.29231f
C1666 VTAIL.n364 VSUBS 0.027936f
C1667 VTAIL.n365 VSUBS 0.015011f
C1668 VTAIL.n366 VSUBS 0.015895f
C1669 VTAIL.n367 VSUBS 0.035482f
C1670 VTAIL.n368 VSUBS 0.035482f
C1671 VTAIL.n369 VSUBS 0.015895f
C1672 VTAIL.n370 VSUBS 0.015011f
C1673 VTAIL.n371 VSUBS 0.027936f
C1674 VTAIL.n372 VSUBS 0.027936f
C1675 VTAIL.n373 VSUBS 0.015011f
C1676 VTAIL.n374 VSUBS 0.015895f
C1677 VTAIL.n375 VSUBS 0.035482f
C1678 VTAIL.n376 VSUBS 0.035482f
C1679 VTAIL.n377 VSUBS 0.015895f
C1680 VTAIL.n378 VSUBS 0.015011f
C1681 VTAIL.n379 VSUBS 0.027936f
C1682 VTAIL.n380 VSUBS 0.027936f
C1683 VTAIL.n381 VSUBS 0.015011f
C1684 VTAIL.n382 VSUBS 0.015895f
C1685 VTAIL.n383 VSUBS 0.035482f
C1686 VTAIL.n384 VSUBS 0.035482f
C1687 VTAIL.n385 VSUBS 0.015895f
C1688 VTAIL.n386 VSUBS 0.015011f
C1689 VTAIL.n387 VSUBS 0.027936f
C1690 VTAIL.n388 VSUBS 0.027936f
C1691 VTAIL.n389 VSUBS 0.015011f
C1692 VTAIL.n390 VSUBS 0.015895f
C1693 VTAIL.n391 VSUBS 0.035482f
C1694 VTAIL.n392 VSUBS 0.035482f
C1695 VTAIL.n393 VSUBS 0.015895f
C1696 VTAIL.n394 VSUBS 0.015011f
C1697 VTAIL.n395 VSUBS 0.027936f
C1698 VTAIL.n396 VSUBS 0.027936f
C1699 VTAIL.n397 VSUBS 0.015011f
C1700 VTAIL.n398 VSUBS 0.015895f
C1701 VTAIL.n399 VSUBS 0.035482f
C1702 VTAIL.n400 VSUBS 0.035482f
C1703 VTAIL.n401 VSUBS 0.035482f
C1704 VTAIL.n402 VSUBS 0.015895f
C1705 VTAIL.n403 VSUBS 0.015011f
C1706 VTAIL.n404 VSUBS 0.027936f
C1707 VTAIL.n405 VSUBS 0.027936f
C1708 VTAIL.n406 VSUBS 0.015011f
C1709 VTAIL.n407 VSUBS 0.015453f
C1710 VTAIL.n408 VSUBS 0.015453f
C1711 VTAIL.n409 VSUBS 0.035482f
C1712 VTAIL.n410 VSUBS 0.035482f
C1713 VTAIL.n411 VSUBS 0.015895f
C1714 VTAIL.n412 VSUBS 0.015011f
C1715 VTAIL.n413 VSUBS 0.027936f
C1716 VTAIL.n414 VSUBS 0.027936f
C1717 VTAIL.n415 VSUBS 0.015011f
C1718 VTAIL.n416 VSUBS 0.015895f
C1719 VTAIL.n417 VSUBS 0.035482f
C1720 VTAIL.n418 VSUBS 0.035482f
C1721 VTAIL.n419 VSUBS 0.015895f
C1722 VTAIL.n420 VSUBS 0.015011f
C1723 VTAIL.n421 VSUBS 0.027936f
C1724 VTAIL.n422 VSUBS 0.027936f
C1725 VTAIL.n423 VSUBS 0.015011f
C1726 VTAIL.n424 VSUBS 0.015895f
C1727 VTAIL.n425 VSUBS 0.035482f
C1728 VTAIL.n426 VSUBS 0.08913f
C1729 VTAIL.n427 VSUBS 0.015895f
C1730 VTAIL.n428 VSUBS 0.015011f
C1731 VTAIL.n429 VSUBS 0.06648f
C1732 VTAIL.n430 VSUBS 0.045024f
C1733 VTAIL.n431 VSUBS 2.40667f
C1734 VDD1.n0 VSUBS 0.030703f
C1735 VDD1.n1 VSUBS 0.027105f
C1736 VDD1.n2 VSUBS 0.014565f
C1737 VDD1.n3 VSUBS 0.034427f
C1738 VDD1.n4 VSUBS 0.015422f
C1739 VDD1.n5 VSUBS 0.027105f
C1740 VDD1.n6 VSUBS 0.014565f
C1741 VDD1.n7 VSUBS 0.034427f
C1742 VDD1.n8 VSUBS 0.015422f
C1743 VDD1.n9 VSUBS 0.027105f
C1744 VDD1.n10 VSUBS 0.014565f
C1745 VDD1.n11 VSUBS 0.034427f
C1746 VDD1.n12 VSUBS 0.015422f
C1747 VDD1.n13 VSUBS 0.027105f
C1748 VDD1.n14 VSUBS 0.014565f
C1749 VDD1.n15 VSUBS 0.034427f
C1750 VDD1.n16 VSUBS 0.034427f
C1751 VDD1.n17 VSUBS 0.015422f
C1752 VDD1.n18 VSUBS 0.027105f
C1753 VDD1.n19 VSUBS 0.014565f
C1754 VDD1.n20 VSUBS 0.034427f
C1755 VDD1.n21 VSUBS 0.015422f
C1756 VDD1.n22 VSUBS 0.027105f
C1757 VDD1.n23 VSUBS 0.014565f
C1758 VDD1.n24 VSUBS 0.034427f
C1759 VDD1.n25 VSUBS 0.015422f
C1760 VDD1.n26 VSUBS 0.027105f
C1761 VDD1.n27 VSUBS 0.014565f
C1762 VDD1.n28 VSUBS 0.034427f
C1763 VDD1.n29 VSUBS 0.015422f
C1764 VDD1.n30 VSUBS 0.027105f
C1765 VDD1.n31 VSUBS 0.014565f
C1766 VDD1.n32 VSUBS 0.034427f
C1767 VDD1.n33 VSUBS 0.015422f
C1768 VDD1.n34 VSUBS 0.223127f
C1769 VDD1.t5 VSUBS 0.073971f
C1770 VDD1.n35 VSUBS 0.02582f
C1771 VDD1.n36 VSUBS 0.021901f
C1772 VDD1.n37 VSUBS 0.014565f
C1773 VDD1.n38 VSUBS 2.22414f
C1774 VDD1.n39 VSUBS 0.027105f
C1775 VDD1.n40 VSUBS 0.014565f
C1776 VDD1.n41 VSUBS 0.015422f
C1777 VDD1.n42 VSUBS 0.034427f
C1778 VDD1.n43 VSUBS 0.034427f
C1779 VDD1.n44 VSUBS 0.015422f
C1780 VDD1.n45 VSUBS 0.014565f
C1781 VDD1.n46 VSUBS 0.027105f
C1782 VDD1.n47 VSUBS 0.027105f
C1783 VDD1.n48 VSUBS 0.014565f
C1784 VDD1.n49 VSUBS 0.015422f
C1785 VDD1.n50 VSUBS 0.034427f
C1786 VDD1.n51 VSUBS 0.034427f
C1787 VDD1.n52 VSUBS 0.015422f
C1788 VDD1.n53 VSUBS 0.014565f
C1789 VDD1.n54 VSUBS 0.027105f
C1790 VDD1.n55 VSUBS 0.027105f
C1791 VDD1.n56 VSUBS 0.014565f
C1792 VDD1.n57 VSUBS 0.015422f
C1793 VDD1.n58 VSUBS 0.034427f
C1794 VDD1.n59 VSUBS 0.034427f
C1795 VDD1.n60 VSUBS 0.015422f
C1796 VDD1.n61 VSUBS 0.014565f
C1797 VDD1.n62 VSUBS 0.027105f
C1798 VDD1.n63 VSUBS 0.027105f
C1799 VDD1.n64 VSUBS 0.014565f
C1800 VDD1.n65 VSUBS 0.015422f
C1801 VDD1.n66 VSUBS 0.034427f
C1802 VDD1.n67 VSUBS 0.034427f
C1803 VDD1.n68 VSUBS 0.015422f
C1804 VDD1.n69 VSUBS 0.014565f
C1805 VDD1.n70 VSUBS 0.027105f
C1806 VDD1.n71 VSUBS 0.027105f
C1807 VDD1.n72 VSUBS 0.014565f
C1808 VDD1.n73 VSUBS 0.015422f
C1809 VDD1.n74 VSUBS 0.034427f
C1810 VDD1.n75 VSUBS 0.034427f
C1811 VDD1.n76 VSUBS 0.015422f
C1812 VDD1.n77 VSUBS 0.014565f
C1813 VDD1.n78 VSUBS 0.027105f
C1814 VDD1.n79 VSUBS 0.027105f
C1815 VDD1.n80 VSUBS 0.014565f
C1816 VDD1.n81 VSUBS 0.014993f
C1817 VDD1.n82 VSUBS 0.014993f
C1818 VDD1.n83 VSUBS 0.034427f
C1819 VDD1.n84 VSUBS 0.034427f
C1820 VDD1.n85 VSUBS 0.015422f
C1821 VDD1.n86 VSUBS 0.014565f
C1822 VDD1.n87 VSUBS 0.027105f
C1823 VDD1.n88 VSUBS 0.027105f
C1824 VDD1.n89 VSUBS 0.014565f
C1825 VDD1.n90 VSUBS 0.015422f
C1826 VDD1.n91 VSUBS 0.034427f
C1827 VDD1.n92 VSUBS 0.034427f
C1828 VDD1.n93 VSUBS 0.015422f
C1829 VDD1.n94 VSUBS 0.014565f
C1830 VDD1.n95 VSUBS 0.027105f
C1831 VDD1.n96 VSUBS 0.027105f
C1832 VDD1.n97 VSUBS 0.014565f
C1833 VDD1.n98 VSUBS 0.015422f
C1834 VDD1.n99 VSUBS 0.034427f
C1835 VDD1.n100 VSUBS 0.086479f
C1836 VDD1.n101 VSUBS 0.015422f
C1837 VDD1.n102 VSUBS 0.014565f
C1838 VDD1.n103 VSUBS 0.064504f
C1839 VDD1.n104 VSUBS 0.076218f
C1840 VDD1.n105 VSUBS 0.030703f
C1841 VDD1.n106 VSUBS 0.027105f
C1842 VDD1.n107 VSUBS 0.014565f
C1843 VDD1.n108 VSUBS 0.034427f
C1844 VDD1.n109 VSUBS 0.015422f
C1845 VDD1.n110 VSUBS 0.027105f
C1846 VDD1.n111 VSUBS 0.014565f
C1847 VDD1.n112 VSUBS 0.034427f
C1848 VDD1.n113 VSUBS 0.015422f
C1849 VDD1.n114 VSUBS 0.027105f
C1850 VDD1.n115 VSUBS 0.014565f
C1851 VDD1.n116 VSUBS 0.034427f
C1852 VDD1.n117 VSUBS 0.015422f
C1853 VDD1.n118 VSUBS 0.027105f
C1854 VDD1.n119 VSUBS 0.014565f
C1855 VDD1.n120 VSUBS 0.034427f
C1856 VDD1.n121 VSUBS 0.015422f
C1857 VDD1.n122 VSUBS 0.027105f
C1858 VDD1.n123 VSUBS 0.014565f
C1859 VDD1.n124 VSUBS 0.034427f
C1860 VDD1.n125 VSUBS 0.015422f
C1861 VDD1.n126 VSUBS 0.027105f
C1862 VDD1.n127 VSUBS 0.014565f
C1863 VDD1.n128 VSUBS 0.034427f
C1864 VDD1.n129 VSUBS 0.015422f
C1865 VDD1.n130 VSUBS 0.027105f
C1866 VDD1.n131 VSUBS 0.014565f
C1867 VDD1.n132 VSUBS 0.034427f
C1868 VDD1.n133 VSUBS 0.015422f
C1869 VDD1.n134 VSUBS 0.027105f
C1870 VDD1.n135 VSUBS 0.014565f
C1871 VDD1.n136 VSUBS 0.034427f
C1872 VDD1.n137 VSUBS 0.015422f
C1873 VDD1.n138 VSUBS 0.223127f
C1874 VDD1.t0 VSUBS 0.073971f
C1875 VDD1.n139 VSUBS 0.02582f
C1876 VDD1.n140 VSUBS 0.021901f
C1877 VDD1.n141 VSUBS 0.014565f
C1878 VDD1.n142 VSUBS 2.22414f
C1879 VDD1.n143 VSUBS 0.027105f
C1880 VDD1.n144 VSUBS 0.014565f
C1881 VDD1.n145 VSUBS 0.015422f
C1882 VDD1.n146 VSUBS 0.034427f
C1883 VDD1.n147 VSUBS 0.034427f
C1884 VDD1.n148 VSUBS 0.015422f
C1885 VDD1.n149 VSUBS 0.014565f
C1886 VDD1.n150 VSUBS 0.027105f
C1887 VDD1.n151 VSUBS 0.027105f
C1888 VDD1.n152 VSUBS 0.014565f
C1889 VDD1.n153 VSUBS 0.015422f
C1890 VDD1.n154 VSUBS 0.034427f
C1891 VDD1.n155 VSUBS 0.034427f
C1892 VDD1.n156 VSUBS 0.015422f
C1893 VDD1.n157 VSUBS 0.014565f
C1894 VDD1.n158 VSUBS 0.027105f
C1895 VDD1.n159 VSUBS 0.027105f
C1896 VDD1.n160 VSUBS 0.014565f
C1897 VDD1.n161 VSUBS 0.015422f
C1898 VDD1.n162 VSUBS 0.034427f
C1899 VDD1.n163 VSUBS 0.034427f
C1900 VDD1.n164 VSUBS 0.015422f
C1901 VDD1.n165 VSUBS 0.014565f
C1902 VDD1.n166 VSUBS 0.027105f
C1903 VDD1.n167 VSUBS 0.027105f
C1904 VDD1.n168 VSUBS 0.014565f
C1905 VDD1.n169 VSUBS 0.015422f
C1906 VDD1.n170 VSUBS 0.034427f
C1907 VDD1.n171 VSUBS 0.034427f
C1908 VDD1.n172 VSUBS 0.015422f
C1909 VDD1.n173 VSUBS 0.014565f
C1910 VDD1.n174 VSUBS 0.027105f
C1911 VDD1.n175 VSUBS 0.027105f
C1912 VDD1.n176 VSUBS 0.014565f
C1913 VDD1.n177 VSUBS 0.015422f
C1914 VDD1.n178 VSUBS 0.034427f
C1915 VDD1.n179 VSUBS 0.034427f
C1916 VDD1.n180 VSUBS 0.034427f
C1917 VDD1.n181 VSUBS 0.015422f
C1918 VDD1.n182 VSUBS 0.014565f
C1919 VDD1.n183 VSUBS 0.027105f
C1920 VDD1.n184 VSUBS 0.027105f
C1921 VDD1.n185 VSUBS 0.014565f
C1922 VDD1.n186 VSUBS 0.014993f
C1923 VDD1.n187 VSUBS 0.014993f
C1924 VDD1.n188 VSUBS 0.034427f
C1925 VDD1.n189 VSUBS 0.034427f
C1926 VDD1.n190 VSUBS 0.015422f
C1927 VDD1.n191 VSUBS 0.014565f
C1928 VDD1.n192 VSUBS 0.027105f
C1929 VDD1.n193 VSUBS 0.027105f
C1930 VDD1.n194 VSUBS 0.014565f
C1931 VDD1.n195 VSUBS 0.015422f
C1932 VDD1.n196 VSUBS 0.034427f
C1933 VDD1.n197 VSUBS 0.034427f
C1934 VDD1.n198 VSUBS 0.015422f
C1935 VDD1.n199 VSUBS 0.014565f
C1936 VDD1.n200 VSUBS 0.027105f
C1937 VDD1.n201 VSUBS 0.027105f
C1938 VDD1.n202 VSUBS 0.014565f
C1939 VDD1.n203 VSUBS 0.015422f
C1940 VDD1.n204 VSUBS 0.034427f
C1941 VDD1.n205 VSUBS 0.086479f
C1942 VDD1.n206 VSUBS 0.015422f
C1943 VDD1.n207 VSUBS 0.014565f
C1944 VDD1.n208 VSUBS 0.064504f
C1945 VDD1.n209 VSUBS 0.075183f
C1946 VDD1.t1 VSUBS 0.40718f
C1947 VDD1.t2 VSUBS 0.40718f
C1948 VDD1.n210 VSUBS 3.4187f
C1949 VDD1.n211 VSUBS 4.32358f
C1950 VDD1.t3 VSUBS 0.40718f
C1951 VDD1.t4 VSUBS 0.40718f
C1952 VDD1.n212 VSUBS 3.40845f
C1953 VDD1.n213 VSUBS 4.2099f
C1954 VP.t1 VSUBS 4.5479f
C1955 VP.n0 VSUBS 1.6585f
C1956 VP.n1 VSUBS 0.024203f
C1957 VP.n2 VSUBS 0.03803f
C1958 VP.n3 VSUBS 0.024203f
C1959 VP.n4 VSUBS 0.033974f
C1960 VP.n5 VSUBS 0.024203f
C1961 VP.n6 VSUBS 0.032635f
C1962 VP.n7 VSUBS 0.024203f
C1963 VP.n8 VSUBS 0.030411f
C1964 VP.t3 VSUBS 4.5479f
C1965 VP.n9 VSUBS 1.6585f
C1966 VP.n10 VSUBS 0.024203f
C1967 VP.n11 VSUBS 0.03803f
C1968 VP.n12 VSUBS 0.024203f
C1969 VP.n13 VSUBS 0.033974f
C1970 VP.t2 VSUBS 4.90812f
C1971 VP.t0 VSUBS 4.5479f
C1972 VP.n14 VSUBS 1.64924f
C1973 VP.n15 VSUBS 1.57799f
C1974 VP.n16 VSUBS 0.302389f
C1975 VP.n17 VSUBS 0.024203f
C1976 VP.n18 VSUBS 0.045109f
C1977 VP.n19 VSUBS 0.045109f
C1978 VP.n20 VSUBS 0.032635f
C1979 VP.n21 VSUBS 0.024203f
C1980 VP.n22 VSUBS 0.024203f
C1981 VP.n23 VSUBS 0.024203f
C1982 VP.n24 VSUBS 0.045109f
C1983 VP.n25 VSUBS 0.045109f
C1984 VP.n26 VSUBS 0.030411f
C1985 VP.n27 VSUBS 0.039064f
C1986 VP.n28 VSUBS 1.70068f
C1987 VP.t5 VSUBS 4.5479f
C1988 VP.n29 VSUBS 1.6585f
C1989 VP.n30 VSUBS 1.71569f
C1990 VP.n31 VSUBS 0.039064f
C1991 VP.n32 VSUBS 0.024203f
C1992 VP.n33 VSUBS 0.045109f
C1993 VP.n34 VSUBS 0.045109f
C1994 VP.n35 VSUBS 0.03803f
C1995 VP.n36 VSUBS 0.024203f
C1996 VP.n37 VSUBS 0.024203f
C1997 VP.n38 VSUBS 0.024203f
C1998 VP.n39 VSUBS 0.045109f
C1999 VP.n40 VSUBS 0.045109f
C2000 VP.t4 VSUBS 4.5479f
C2001 VP.n41 VSUBS 1.56529f
C2002 VP.n42 VSUBS 0.033974f
C2003 VP.n43 VSUBS 0.024203f
C2004 VP.n44 VSUBS 0.024203f
C2005 VP.n45 VSUBS 0.024203f
C2006 VP.n46 VSUBS 0.045109f
C2007 VP.n47 VSUBS 0.045109f
C2008 VP.n48 VSUBS 0.032635f
C2009 VP.n49 VSUBS 0.024203f
C2010 VP.n50 VSUBS 0.024203f
C2011 VP.n51 VSUBS 0.024203f
C2012 VP.n52 VSUBS 0.045109f
C2013 VP.n53 VSUBS 0.045109f
C2014 VP.n54 VSUBS 0.030411f
C2015 VP.n55 VSUBS 0.039064f
C2016 VP.n56 VSUBS 0.067483f
.ends

