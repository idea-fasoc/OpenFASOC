// Module definition for lc-dco
`timescale 1ns/1ps
module lc_dco(sw, outp, outn, div_clk, Ibias);
    output outp, outn, div_clk;
    inout Ibias;
    input [7:0] sw;
    real Freq;
    parameter DivReg=4;
    reg outpwire, outnwire;
    reg [DivReg-1:0]div_reg;
    // Freq LUT
    initial begin
        outpwire <= 1'b1;
        outnwire <= 1'b0;
    end
    always @ (*)
        begin
        case (sw)
            1  : Freq = 3.287149;
            2  : Freq = 3.280689;
            3  : Freq = 3.274255;
            4  : Freq = 3.267224;
            5  : Freq = 3.260223;
            6  : Freq = 3.253252;
            7  : Freq = 3.246311;
            8  : Freq = 3.238598;
            9  : Freq = 3.230921;
            10 : Freq = 3.223281;
            11 : Freq = 3.215677;
            12 : Freq = 3.208109;
            13 : Freq = 3.200576;
            14 : Freq = 3.193079;
            15 : Freq = 3.185616;
            16 : Freq = 3.177806;
            17 : Freq = 3.170033;
            18 : Freq = 3.162298;
            19 : Freq = 3.154601;
            20 : Freq = 3.146942;
            21 : Freq = 3.139319;
            22 : Freq = 3.131734;
            23 : Freq = 3.124185;
            24 : Freq = 3.116672;
            25 : Freq = 3.109195;
            26 : Freq = 3.101754;
            27 : Freq = 3.094349;
            28 : Freq = 3.086979;
            29 : Freq = 3.079644;
            30 : Freq = 3.072344;
            31 : Freq = 3.065078;
            32 : Freq = 3.058144;
            33 : Freq = 3.051241;
            34 : Freq = 3.044369;
            35 : Freq = 3.037529;
            36 : Freq = 3.030719;
            37 : Freq = 3.023939;
            38 : Freq = 3.017190;
            39 : Freq = 3.010470;
            40 : Freq = 3.003781;
            41 : Freq = 2.997121;
            42 : Freq = 2.990491;
            43 : Freq = 2.983890;
            44 : Freq = 2.977318;
            45 : Freq = 2.970775;
            46 : Freq = 2.964261;
            47 : Freq = 2.957775;
            48 : Freq = 2.951317;
            49 : Freq = 2.944888;
            50 : Freq = 2.938486;
            51 : Freq = 2.932113;
            52 : Freq = 2.925767;
            53 : Freq = 2.919448;
            54 : Freq = 2.913157;
            55 : Freq = 2.906892;
            56 : Freq = 2.900655;
            57 : Freq = 2.894444;
            58 : Freq = 2.888260;
            59 : Freq = 2.882102;
            60 : Freq = 2.875970;
            61 : Freq = 2.869865;
            62 : Freq = 2.863785;
            63 : Freq = 2.857731;
            64 : Freq = 2.852320;
            65 : Freq = 2.846929;
            66 : Freq = 2.841559;
            67 : Freq = 2.836209;
            68 : Freq = 2.830879;
            69 : Freq = 2.825569;
            70 : Freq = 2.820279;
            71 : Freq = 2.815009;
            72 : Freq = 2.809759;
            73 : Freq = 2.804528;
            74 : Freq = 2.799316;
            75 : Freq = 2.794124;
            76 : Freq = 2.788951;
            77 : Freq = 2.783797;
            78 : Freq = 2.778662;
            79 : Freq = 2.773546;
            80 : Freq = 2.768449;
            81 : Freq = 2.763371;
            82 : Freq = 2.758311;
            83 : Freq = 2.753269;
            84 : Freq = 2.748246;
            85 : Freq = 2.743242;
            86 : Freq = 2.738255;
            87 : Freq = 2.733287;
            88 : Freq = 2.728337;
            89 : Freq = 2.723404;
            90 : Freq = 2.718489;
            91 : Freq = 2.713592;
            92 : Freq = 2.708713;
            93 : Freq = 2.703851;
            94 : Freq = 2.699007;
            95 : Freq = 2.694180;
            96 : Freq = 2.689370;
            97 : Freq = 2.684577;
            98 : Freq = 2.679801;
            99 : Freq = 2.675043;
            100: Freq = 2.670301;
            101: Freq = 2.665576;
            102: Freq = 2.660867;
            103: Freq = 2.656176;
            104: Freq = 2.651500;
            105: Freq = 2.646842;
            106: Freq = 2.642199;
            107: Freq = 2.637573;
            108: Freq = 2.632963;
            109: Freq = 2.628369;
            110: Freq = 2.623791;
            111: Freq = 2.619229;
            112: Freq = 2.614683;
            113: Freq = 2.610152;
            114: Freq = 2.605638;
            115: Freq = 2.601138;
            116: Freq = 2.596655;
            117: Freq = 2.592186;
            118: Freq = 2.587734;
            119: Freq = 2.583296;
            120: Freq = 2.578874;
            121: Freq = 2.574466;
            122: Freq = 2.570074;
            123: Freq = 2.565697;
            124: Freq = 2.561334;
            125: Freq = 2.556987;
            126: Freq = 2.552654;
            127: Freq = 2.548336;
            128: Freq = 2.544632;
            129: Freq = 2.540939;
            130: Freq = 2.537257;
            131: Freq = 2.533586;
            132: Freq = 2.529925;
            133: Freq = 2.526275;
            134: Freq = 2.522635;
            135: Freq = 2.519006;
            136: Freq = 2.515388;
            137: Freq = 2.511779;
            138: Freq = 2.508181;
            139: Freq = 2.504593;
            140: Freq = 2.501016;
            141: Freq = 2.497449;
            142: Freq = 2.493891;
            143: Freq = 2.490344;
            144: Freq = 2.486808;
            145: Freq = 2.483281;
            146: Freq = 2.479764;
            147: Freq = 2.476257;
            148: Freq = 2.472760;
            149: Freq = 2.469273;
            150: Freq = 2.465795;
            151: Freq = 2.462328;
            152: Freq = 2.458870;
            153: Freq = 2.455422;
            154: Freq = 2.451983;
            155: Freq = 2.448554;
            156: Freq = 2.445135;
            157: Freq = 2.441725;
            158: Freq = 2.438325;
            159: Freq = 2.434934;
            160: Freq = 2.431553;
            161: Freq = 2.428181;
            162: Freq = 2.424818;
            163: Freq = 2.421465;
            164: Freq = 2.418120;
            165: Freq = 2.414786;
            166: Freq = 2.411460;
            167: Freq = 2.408143;
            168: Freq = 2.404836;
            169: Freq = 2.401537;
            170: Freq = 2.398248;
            171: Freq = 2.394968;
            172: Freq = 2.391696;
            173: Freq = 2.388434;
            174: Freq = 2.385180;
            175: Freq = 2.381936;
            176: Freq = 2.378700;
            177: Freq = 2.375473;
            178: Freq = 2.372254;
            179: Freq = 2.369045;
            180: Freq = 2.365844;
            181: Freq = 2.362651;
            182: Freq = 2.359467;
            183: Freq = 2.356292;
            184: Freq = 2.353126;
            185: Freq = 2.349968;
            186: Freq = 2.346818;
            187: Freq = 2.343677;
            188: Freq = 2.340544;
            189: Freq = 2.337419;
            190: Freq = 2.334303;
            191: Freq = 2.331195;
            192: Freq = 2.328096;
            193: Freq = 2.325004;
            194: Freq = 2.321921;
            195: Freq = 2.318846;
            196: Freq = 2.315779;
            197: Freq = 2.312721;
            198: Freq = 2.309670;
            199: Freq = 2.306627;
            200: Freq = 2.303593;
            201: Freq = 2.300566;
            202: Freq = 2.297547;
            203: Freq = 2.294536;
            204: Freq = 2.291533;
            205: Freq = 2.288538;
            206: Freq = 2.285551;
            207: Freq = 2.282572;
            208: Freq = 2.279600;
            209: Freq = 2.276636;
            210: Freq = 2.273679;
            211: Freq = 2.270731;
            212: Freq = 2.267790;
            213: Freq = 2.264856;
            214: Freq = 2.261931;
            215: Freq = 2.259012;
            216: Freq = 2.256102;
            217: Freq = 2.253198;
            218: Freq = 2.250303;
            219: Freq = 2.247414;
            220: Freq = 2.244533;
            221: Freq = 2.241660;
            222: Freq = 2.238794;
            223: Freq = 2.235935;
            224: Freq = 2.233083;
            225: Freq = 2.230239;
            226: Freq = 2.227402;
            227: Freq = 2.224572;
            228: Freq = 2.221749;
            229: Freq = 2.218934;
            230: Freq = 2.216125;
            231: Freq = 2.213324;
            232: Freq = 2.210529;
            233: Freq = 2.207742;
            234: Freq = 2.204962;
            235: Freq = 2.202189;
            236: Freq = 2.199423;
            237: Freq = 2.196663;
            238: Freq = 2.193911;
            239: Freq = 2.191165;
            240: Freq = 2.188427;
            241: Freq = 2.185695;
            242: Freq = 2.182970;
            243: Freq = 2.180252;
            244: Freq = 2.177540;
            245: Freq = 2.174836;
            246: Freq = 2.172138;
            247: Freq = 2.169447;
            248: Freq = 2.166762;
            249: Freq = 2.164084;
            250: Freq = 2.161412;
            251: Freq = 2.158748;
            252: Freq = 2.156089;
            253: Freq = 2.153438;
            254: Freq = 2.150793;
            255: Freq = 2.148154;
	    default: Freq = 1; // Catch for not oscillating
        endcase
    end
    // NOTE:
    // Only this assignment works in verilator, doesn like delay on RHS
	always @(*) begin
		//$display("Freq is %d",Freq);
		#(1/(2*Freq)) outpwire <= ~outpwire;
	end
	//forever begin
	//	outpwire = 1'b0;
	//	#(1/(2*Freq));
	//	outpwire =1'b1;
	//	#(1/(2*Freq));
	//end
	assign outp = outpwire;
	assign outn = ~outpwire;

    initial begin
        div_reg =1'b0;
    end
    always @(posedge outp) begin
        div_reg = div_reg+1;
    end
    // Divider Module (Programmable??)
    assign div_clk = div_reg[DivReg-1];
endmodule
