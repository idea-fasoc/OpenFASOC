* NGSPICE file created from diff_pair_sample_0524.ext - technology: sky130A

.subckt diff_pair_sample_0524 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=1.6467 ps=10.31 w=9.98 l=3.21
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=0 ps=0 w=9.98 l=3.21
X2 VDD1.t4 VP.t1 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=1.6467 ps=10.31 w=9.98 l=3.21
X3 VTAIL.t8 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=1.6467 ps=10.31 w=9.98 l=3.21
X4 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=1.6467 ps=10.31 w=9.98 l=3.21
X5 VDD1.t2 VP.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=3.8922 ps=20.74 w=9.98 l=3.21
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=0 ps=0 w=9.98 l=3.21
X7 VTAIL.t10 VP.t4 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=1.6467 ps=10.31 w=9.98 l=3.21
X8 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=3.8922 ps=20.74 w=9.98 l=3.21
X9 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=1.6467 ps=10.31 w=9.98 l=3.21
X10 VDD2.t2 VN.t3 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=3.8922 ps=20.74 w=9.98 l=3.21
X11 VDD1.t0 VP.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=3.8922 ps=20.74 w=9.98 l=3.21
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=0 ps=0 w=9.98 l=3.21
X13 VTAIL.t0 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6467 pd=10.31 as=1.6467 ps=10.31 w=9.98 l=3.21
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=0 ps=0 w=9.98 l=3.21
X15 VDD2.t0 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.8922 pd=20.74 as=1.6467 ps=10.31 w=9.98 l=3.21
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t0 107.742
R22 VP.n27 VP.n8 75.7718
R23 VP.n50 VP.n0 75.7718
R24 VP.n26 VP.n9 75.7718
R25 VP.n8 VP.t1 74.9282
R26 VP.n4 VP.t4 74.9282
R27 VP.n0 VP.t5 74.9282
R28 VP.n9 VP.t3 74.9282
R29 VP.n13 VP.t2 74.9282
R30 VP.n14 VP.n13 61.8768
R31 VP.n27 VP.n26 49.6203
R32 VP.n31 VP.n6 42.3581
R33 VP.n46 VP.n2 42.3581
R34 VP.n22 VP.n11 42.3581
R35 VP.n35 VP.n6 38.4631
R36 VP.n42 VP.n2 38.4631
R37 VP.n18 VP.n11 38.4631
R38 VP.n30 VP.n29 24.3439
R39 VP.n31 VP.n30 24.3439
R40 VP.n36 VP.n35 24.3439
R41 VP.n37 VP.n36 24.3439
R42 VP.n41 VP.n40 24.3439
R43 VP.n42 VP.n41 24.3439
R44 VP.n47 VP.n46 24.3439
R45 VP.n48 VP.n47 24.3439
R46 VP.n23 VP.n22 24.3439
R47 VP.n24 VP.n23 24.3439
R48 VP.n17 VP.n16 24.3439
R49 VP.n18 VP.n17 24.3439
R50 VP.n29 VP.n8 14.1197
R51 VP.n48 VP.n0 14.1197
R52 VP.n24 VP.n9 14.1197
R53 VP.n37 VP.n4 12.1722
R54 VP.n40 VP.n4 12.1722
R55 VP.n16 VP.n13 12.1722
R56 VP.n15 VP.n14 4.19698
R57 VP.n26 VP.n25 0.355081
R58 VP.n28 VP.n27 0.355081
R59 VP.n50 VP.n49 0.355081
R60 VP VP.n50 0.26685
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VTAIL.n218 VTAIL.n170 289.615
R81 VTAIL.n50 VTAIL.n2 289.615
R82 VTAIL.n164 VTAIL.n116 289.615
R83 VTAIL.n108 VTAIL.n60 289.615
R84 VTAIL.n186 VTAIL.n185 185
R85 VTAIL.n191 VTAIL.n190 185
R86 VTAIL.n193 VTAIL.n192 185
R87 VTAIL.n182 VTAIL.n181 185
R88 VTAIL.n199 VTAIL.n198 185
R89 VTAIL.n201 VTAIL.n200 185
R90 VTAIL.n178 VTAIL.n177 185
R91 VTAIL.n208 VTAIL.n207 185
R92 VTAIL.n209 VTAIL.n176 185
R93 VTAIL.n211 VTAIL.n210 185
R94 VTAIL.n174 VTAIL.n173 185
R95 VTAIL.n217 VTAIL.n216 185
R96 VTAIL.n219 VTAIL.n218 185
R97 VTAIL.n18 VTAIL.n17 185
R98 VTAIL.n23 VTAIL.n22 185
R99 VTAIL.n25 VTAIL.n24 185
R100 VTAIL.n14 VTAIL.n13 185
R101 VTAIL.n31 VTAIL.n30 185
R102 VTAIL.n33 VTAIL.n32 185
R103 VTAIL.n10 VTAIL.n9 185
R104 VTAIL.n40 VTAIL.n39 185
R105 VTAIL.n41 VTAIL.n8 185
R106 VTAIL.n43 VTAIL.n42 185
R107 VTAIL.n6 VTAIL.n5 185
R108 VTAIL.n49 VTAIL.n48 185
R109 VTAIL.n51 VTAIL.n50 185
R110 VTAIL.n165 VTAIL.n164 185
R111 VTAIL.n163 VTAIL.n162 185
R112 VTAIL.n120 VTAIL.n119 185
R113 VTAIL.n157 VTAIL.n156 185
R114 VTAIL.n155 VTAIL.n122 185
R115 VTAIL.n154 VTAIL.n153 185
R116 VTAIL.n125 VTAIL.n123 185
R117 VTAIL.n148 VTAIL.n147 185
R118 VTAIL.n146 VTAIL.n145 185
R119 VTAIL.n129 VTAIL.n128 185
R120 VTAIL.n140 VTAIL.n139 185
R121 VTAIL.n138 VTAIL.n137 185
R122 VTAIL.n133 VTAIL.n132 185
R123 VTAIL.n109 VTAIL.n108 185
R124 VTAIL.n107 VTAIL.n106 185
R125 VTAIL.n64 VTAIL.n63 185
R126 VTAIL.n101 VTAIL.n100 185
R127 VTAIL.n99 VTAIL.n66 185
R128 VTAIL.n98 VTAIL.n97 185
R129 VTAIL.n69 VTAIL.n67 185
R130 VTAIL.n92 VTAIL.n91 185
R131 VTAIL.n90 VTAIL.n89 185
R132 VTAIL.n73 VTAIL.n72 185
R133 VTAIL.n84 VTAIL.n83 185
R134 VTAIL.n82 VTAIL.n81 185
R135 VTAIL.n77 VTAIL.n76 185
R136 VTAIL.n187 VTAIL.t3 149.524
R137 VTAIL.n19 VTAIL.t6 149.524
R138 VTAIL.n134 VTAIL.t11 149.524
R139 VTAIL.n78 VTAIL.t5 149.524
R140 VTAIL.n191 VTAIL.n185 104.615
R141 VTAIL.n192 VTAIL.n191 104.615
R142 VTAIL.n192 VTAIL.n181 104.615
R143 VTAIL.n199 VTAIL.n181 104.615
R144 VTAIL.n200 VTAIL.n199 104.615
R145 VTAIL.n200 VTAIL.n177 104.615
R146 VTAIL.n208 VTAIL.n177 104.615
R147 VTAIL.n209 VTAIL.n208 104.615
R148 VTAIL.n210 VTAIL.n209 104.615
R149 VTAIL.n210 VTAIL.n173 104.615
R150 VTAIL.n217 VTAIL.n173 104.615
R151 VTAIL.n218 VTAIL.n217 104.615
R152 VTAIL.n23 VTAIL.n17 104.615
R153 VTAIL.n24 VTAIL.n23 104.615
R154 VTAIL.n24 VTAIL.n13 104.615
R155 VTAIL.n31 VTAIL.n13 104.615
R156 VTAIL.n32 VTAIL.n31 104.615
R157 VTAIL.n32 VTAIL.n9 104.615
R158 VTAIL.n40 VTAIL.n9 104.615
R159 VTAIL.n41 VTAIL.n40 104.615
R160 VTAIL.n42 VTAIL.n41 104.615
R161 VTAIL.n42 VTAIL.n5 104.615
R162 VTAIL.n49 VTAIL.n5 104.615
R163 VTAIL.n50 VTAIL.n49 104.615
R164 VTAIL.n164 VTAIL.n163 104.615
R165 VTAIL.n163 VTAIL.n119 104.615
R166 VTAIL.n156 VTAIL.n119 104.615
R167 VTAIL.n156 VTAIL.n155 104.615
R168 VTAIL.n155 VTAIL.n154 104.615
R169 VTAIL.n154 VTAIL.n123 104.615
R170 VTAIL.n147 VTAIL.n123 104.615
R171 VTAIL.n147 VTAIL.n146 104.615
R172 VTAIL.n146 VTAIL.n128 104.615
R173 VTAIL.n139 VTAIL.n128 104.615
R174 VTAIL.n139 VTAIL.n138 104.615
R175 VTAIL.n138 VTAIL.n132 104.615
R176 VTAIL.n108 VTAIL.n107 104.615
R177 VTAIL.n107 VTAIL.n63 104.615
R178 VTAIL.n100 VTAIL.n63 104.615
R179 VTAIL.n100 VTAIL.n99 104.615
R180 VTAIL.n99 VTAIL.n98 104.615
R181 VTAIL.n98 VTAIL.n67 104.615
R182 VTAIL.n91 VTAIL.n67 104.615
R183 VTAIL.n91 VTAIL.n90 104.615
R184 VTAIL.n90 VTAIL.n72 104.615
R185 VTAIL.n83 VTAIL.n72 104.615
R186 VTAIL.n83 VTAIL.n82 104.615
R187 VTAIL.n82 VTAIL.n76 104.615
R188 VTAIL.t3 VTAIL.n185 52.3082
R189 VTAIL.t6 VTAIL.n17 52.3082
R190 VTAIL.t11 VTAIL.n132 52.3082
R191 VTAIL.t5 VTAIL.n76 52.3082
R192 VTAIL.n115 VTAIL.n114 46.3494
R193 VTAIL.n59 VTAIL.n58 46.3494
R194 VTAIL.n1 VTAIL.n0 46.3492
R195 VTAIL.n57 VTAIL.n56 46.3492
R196 VTAIL.n223 VTAIL.n222 32.5732
R197 VTAIL.n55 VTAIL.n54 32.5732
R198 VTAIL.n169 VTAIL.n168 32.5732
R199 VTAIL.n113 VTAIL.n112 32.5732
R200 VTAIL.n59 VTAIL.n57 27.0738
R201 VTAIL.n223 VTAIL.n169 24.0221
R202 VTAIL.n211 VTAIL.n176 13.1884
R203 VTAIL.n43 VTAIL.n8 13.1884
R204 VTAIL.n157 VTAIL.n122 13.1884
R205 VTAIL.n101 VTAIL.n66 13.1884
R206 VTAIL.n207 VTAIL.n206 12.8005
R207 VTAIL.n212 VTAIL.n174 12.8005
R208 VTAIL.n39 VTAIL.n38 12.8005
R209 VTAIL.n44 VTAIL.n6 12.8005
R210 VTAIL.n158 VTAIL.n120 12.8005
R211 VTAIL.n153 VTAIL.n124 12.8005
R212 VTAIL.n102 VTAIL.n64 12.8005
R213 VTAIL.n97 VTAIL.n68 12.8005
R214 VTAIL.n205 VTAIL.n178 12.0247
R215 VTAIL.n216 VTAIL.n215 12.0247
R216 VTAIL.n37 VTAIL.n10 12.0247
R217 VTAIL.n48 VTAIL.n47 12.0247
R218 VTAIL.n162 VTAIL.n161 12.0247
R219 VTAIL.n152 VTAIL.n125 12.0247
R220 VTAIL.n106 VTAIL.n105 12.0247
R221 VTAIL.n96 VTAIL.n69 12.0247
R222 VTAIL.n202 VTAIL.n201 11.249
R223 VTAIL.n219 VTAIL.n172 11.249
R224 VTAIL.n34 VTAIL.n33 11.249
R225 VTAIL.n51 VTAIL.n4 11.249
R226 VTAIL.n165 VTAIL.n118 11.249
R227 VTAIL.n149 VTAIL.n148 11.249
R228 VTAIL.n109 VTAIL.n62 11.249
R229 VTAIL.n93 VTAIL.n92 11.249
R230 VTAIL.n198 VTAIL.n180 10.4732
R231 VTAIL.n220 VTAIL.n170 10.4732
R232 VTAIL.n30 VTAIL.n12 10.4732
R233 VTAIL.n52 VTAIL.n2 10.4732
R234 VTAIL.n166 VTAIL.n116 10.4732
R235 VTAIL.n145 VTAIL.n127 10.4732
R236 VTAIL.n110 VTAIL.n60 10.4732
R237 VTAIL.n89 VTAIL.n71 10.4732
R238 VTAIL.n187 VTAIL.n186 10.2747
R239 VTAIL.n19 VTAIL.n18 10.2747
R240 VTAIL.n134 VTAIL.n133 10.2747
R241 VTAIL.n78 VTAIL.n77 10.2747
R242 VTAIL.n197 VTAIL.n182 9.69747
R243 VTAIL.n29 VTAIL.n14 9.69747
R244 VTAIL.n144 VTAIL.n129 9.69747
R245 VTAIL.n88 VTAIL.n73 9.69747
R246 VTAIL.n222 VTAIL.n221 9.45567
R247 VTAIL.n54 VTAIL.n53 9.45567
R248 VTAIL.n168 VTAIL.n167 9.45567
R249 VTAIL.n112 VTAIL.n111 9.45567
R250 VTAIL.n221 VTAIL.n220 9.3005
R251 VTAIL.n172 VTAIL.n171 9.3005
R252 VTAIL.n215 VTAIL.n214 9.3005
R253 VTAIL.n213 VTAIL.n212 9.3005
R254 VTAIL.n189 VTAIL.n188 9.3005
R255 VTAIL.n184 VTAIL.n183 9.3005
R256 VTAIL.n195 VTAIL.n194 9.3005
R257 VTAIL.n197 VTAIL.n196 9.3005
R258 VTAIL.n180 VTAIL.n179 9.3005
R259 VTAIL.n203 VTAIL.n202 9.3005
R260 VTAIL.n205 VTAIL.n204 9.3005
R261 VTAIL.n206 VTAIL.n175 9.3005
R262 VTAIL.n53 VTAIL.n52 9.3005
R263 VTAIL.n4 VTAIL.n3 9.3005
R264 VTAIL.n47 VTAIL.n46 9.3005
R265 VTAIL.n45 VTAIL.n44 9.3005
R266 VTAIL.n21 VTAIL.n20 9.3005
R267 VTAIL.n16 VTAIL.n15 9.3005
R268 VTAIL.n27 VTAIL.n26 9.3005
R269 VTAIL.n29 VTAIL.n28 9.3005
R270 VTAIL.n12 VTAIL.n11 9.3005
R271 VTAIL.n35 VTAIL.n34 9.3005
R272 VTAIL.n37 VTAIL.n36 9.3005
R273 VTAIL.n38 VTAIL.n7 9.3005
R274 VTAIL.n136 VTAIL.n135 9.3005
R275 VTAIL.n131 VTAIL.n130 9.3005
R276 VTAIL.n142 VTAIL.n141 9.3005
R277 VTAIL.n144 VTAIL.n143 9.3005
R278 VTAIL.n127 VTAIL.n126 9.3005
R279 VTAIL.n150 VTAIL.n149 9.3005
R280 VTAIL.n152 VTAIL.n151 9.3005
R281 VTAIL.n124 VTAIL.n121 9.3005
R282 VTAIL.n167 VTAIL.n166 9.3005
R283 VTAIL.n118 VTAIL.n117 9.3005
R284 VTAIL.n161 VTAIL.n160 9.3005
R285 VTAIL.n159 VTAIL.n158 9.3005
R286 VTAIL.n80 VTAIL.n79 9.3005
R287 VTAIL.n75 VTAIL.n74 9.3005
R288 VTAIL.n86 VTAIL.n85 9.3005
R289 VTAIL.n88 VTAIL.n87 9.3005
R290 VTAIL.n71 VTAIL.n70 9.3005
R291 VTAIL.n94 VTAIL.n93 9.3005
R292 VTAIL.n96 VTAIL.n95 9.3005
R293 VTAIL.n68 VTAIL.n65 9.3005
R294 VTAIL.n111 VTAIL.n110 9.3005
R295 VTAIL.n62 VTAIL.n61 9.3005
R296 VTAIL.n105 VTAIL.n104 9.3005
R297 VTAIL.n103 VTAIL.n102 9.3005
R298 VTAIL.n194 VTAIL.n193 8.92171
R299 VTAIL.n26 VTAIL.n25 8.92171
R300 VTAIL.n141 VTAIL.n140 8.92171
R301 VTAIL.n85 VTAIL.n84 8.92171
R302 VTAIL.n190 VTAIL.n184 8.14595
R303 VTAIL.n22 VTAIL.n16 8.14595
R304 VTAIL.n137 VTAIL.n131 8.14595
R305 VTAIL.n81 VTAIL.n75 8.14595
R306 VTAIL.n189 VTAIL.n186 7.3702
R307 VTAIL.n21 VTAIL.n18 7.3702
R308 VTAIL.n136 VTAIL.n133 7.3702
R309 VTAIL.n80 VTAIL.n77 7.3702
R310 VTAIL.n190 VTAIL.n189 5.81868
R311 VTAIL.n22 VTAIL.n21 5.81868
R312 VTAIL.n137 VTAIL.n136 5.81868
R313 VTAIL.n81 VTAIL.n80 5.81868
R314 VTAIL.n193 VTAIL.n184 5.04292
R315 VTAIL.n25 VTAIL.n16 5.04292
R316 VTAIL.n140 VTAIL.n131 5.04292
R317 VTAIL.n84 VTAIL.n75 5.04292
R318 VTAIL.n194 VTAIL.n182 4.26717
R319 VTAIL.n26 VTAIL.n14 4.26717
R320 VTAIL.n141 VTAIL.n129 4.26717
R321 VTAIL.n85 VTAIL.n73 4.26717
R322 VTAIL.n198 VTAIL.n197 3.49141
R323 VTAIL.n222 VTAIL.n170 3.49141
R324 VTAIL.n30 VTAIL.n29 3.49141
R325 VTAIL.n54 VTAIL.n2 3.49141
R326 VTAIL.n168 VTAIL.n116 3.49141
R327 VTAIL.n145 VTAIL.n144 3.49141
R328 VTAIL.n112 VTAIL.n60 3.49141
R329 VTAIL.n89 VTAIL.n88 3.49141
R330 VTAIL.n113 VTAIL.n59 3.05222
R331 VTAIL.n169 VTAIL.n115 3.05222
R332 VTAIL.n57 VTAIL.n55 3.05222
R333 VTAIL.n188 VTAIL.n187 2.84303
R334 VTAIL.n20 VTAIL.n19 2.84303
R335 VTAIL.n135 VTAIL.n134 2.84303
R336 VTAIL.n79 VTAIL.n78 2.84303
R337 VTAIL.n201 VTAIL.n180 2.71565
R338 VTAIL.n220 VTAIL.n219 2.71565
R339 VTAIL.n33 VTAIL.n12 2.71565
R340 VTAIL.n52 VTAIL.n51 2.71565
R341 VTAIL.n166 VTAIL.n165 2.71565
R342 VTAIL.n148 VTAIL.n127 2.71565
R343 VTAIL.n110 VTAIL.n109 2.71565
R344 VTAIL.n92 VTAIL.n71 2.71565
R345 VTAIL VTAIL.n223 2.2311
R346 VTAIL.n115 VTAIL.n113 1.99619
R347 VTAIL.n55 VTAIL.n1 1.99619
R348 VTAIL.n0 VTAIL.t2 1.98447
R349 VTAIL.n0 VTAIL.t1 1.98447
R350 VTAIL.n56 VTAIL.t9 1.98447
R351 VTAIL.n56 VTAIL.t10 1.98447
R352 VTAIL.n114 VTAIL.t7 1.98447
R353 VTAIL.n114 VTAIL.t8 1.98447
R354 VTAIL.n58 VTAIL.t4 1.98447
R355 VTAIL.n58 VTAIL.t0 1.98447
R356 VTAIL.n202 VTAIL.n178 1.93989
R357 VTAIL.n216 VTAIL.n172 1.93989
R358 VTAIL.n34 VTAIL.n10 1.93989
R359 VTAIL.n48 VTAIL.n4 1.93989
R360 VTAIL.n162 VTAIL.n118 1.93989
R361 VTAIL.n149 VTAIL.n125 1.93989
R362 VTAIL.n106 VTAIL.n62 1.93989
R363 VTAIL.n93 VTAIL.n69 1.93989
R364 VTAIL.n207 VTAIL.n205 1.16414
R365 VTAIL.n215 VTAIL.n174 1.16414
R366 VTAIL.n39 VTAIL.n37 1.16414
R367 VTAIL.n47 VTAIL.n6 1.16414
R368 VTAIL.n161 VTAIL.n120 1.16414
R369 VTAIL.n153 VTAIL.n152 1.16414
R370 VTAIL.n105 VTAIL.n64 1.16414
R371 VTAIL.n97 VTAIL.n96 1.16414
R372 VTAIL VTAIL.n1 0.821621
R373 VTAIL.n206 VTAIL.n176 0.388379
R374 VTAIL.n212 VTAIL.n211 0.388379
R375 VTAIL.n38 VTAIL.n8 0.388379
R376 VTAIL.n44 VTAIL.n43 0.388379
R377 VTAIL.n158 VTAIL.n157 0.388379
R378 VTAIL.n124 VTAIL.n122 0.388379
R379 VTAIL.n102 VTAIL.n101 0.388379
R380 VTAIL.n68 VTAIL.n66 0.388379
R381 VTAIL.n188 VTAIL.n183 0.155672
R382 VTAIL.n195 VTAIL.n183 0.155672
R383 VTAIL.n196 VTAIL.n195 0.155672
R384 VTAIL.n196 VTAIL.n179 0.155672
R385 VTAIL.n203 VTAIL.n179 0.155672
R386 VTAIL.n204 VTAIL.n203 0.155672
R387 VTAIL.n204 VTAIL.n175 0.155672
R388 VTAIL.n213 VTAIL.n175 0.155672
R389 VTAIL.n214 VTAIL.n213 0.155672
R390 VTAIL.n214 VTAIL.n171 0.155672
R391 VTAIL.n221 VTAIL.n171 0.155672
R392 VTAIL.n20 VTAIL.n15 0.155672
R393 VTAIL.n27 VTAIL.n15 0.155672
R394 VTAIL.n28 VTAIL.n27 0.155672
R395 VTAIL.n28 VTAIL.n11 0.155672
R396 VTAIL.n35 VTAIL.n11 0.155672
R397 VTAIL.n36 VTAIL.n35 0.155672
R398 VTAIL.n36 VTAIL.n7 0.155672
R399 VTAIL.n45 VTAIL.n7 0.155672
R400 VTAIL.n46 VTAIL.n45 0.155672
R401 VTAIL.n46 VTAIL.n3 0.155672
R402 VTAIL.n53 VTAIL.n3 0.155672
R403 VTAIL.n167 VTAIL.n117 0.155672
R404 VTAIL.n160 VTAIL.n117 0.155672
R405 VTAIL.n160 VTAIL.n159 0.155672
R406 VTAIL.n159 VTAIL.n121 0.155672
R407 VTAIL.n151 VTAIL.n121 0.155672
R408 VTAIL.n151 VTAIL.n150 0.155672
R409 VTAIL.n150 VTAIL.n126 0.155672
R410 VTAIL.n143 VTAIL.n126 0.155672
R411 VTAIL.n143 VTAIL.n142 0.155672
R412 VTAIL.n142 VTAIL.n130 0.155672
R413 VTAIL.n135 VTAIL.n130 0.155672
R414 VTAIL.n111 VTAIL.n61 0.155672
R415 VTAIL.n104 VTAIL.n61 0.155672
R416 VTAIL.n104 VTAIL.n103 0.155672
R417 VTAIL.n103 VTAIL.n65 0.155672
R418 VTAIL.n95 VTAIL.n65 0.155672
R419 VTAIL.n95 VTAIL.n94 0.155672
R420 VTAIL.n94 VTAIL.n70 0.155672
R421 VTAIL.n87 VTAIL.n70 0.155672
R422 VTAIL.n87 VTAIL.n86 0.155672
R423 VTAIL.n86 VTAIL.n74 0.155672
R424 VTAIL.n79 VTAIL.n74 0.155672
R425 VDD1.n48 VDD1.n0 289.615
R426 VDD1.n101 VDD1.n53 289.615
R427 VDD1.n49 VDD1.n48 185
R428 VDD1.n47 VDD1.n46 185
R429 VDD1.n4 VDD1.n3 185
R430 VDD1.n41 VDD1.n40 185
R431 VDD1.n39 VDD1.n6 185
R432 VDD1.n38 VDD1.n37 185
R433 VDD1.n9 VDD1.n7 185
R434 VDD1.n32 VDD1.n31 185
R435 VDD1.n30 VDD1.n29 185
R436 VDD1.n13 VDD1.n12 185
R437 VDD1.n24 VDD1.n23 185
R438 VDD1.n22 VDD1.n21 185
R439 VDD1.n17 VDD1.n16 185
R440 VDD1.n69 VDD1.n68 185
R441 VDD1.n74 VDD1.n73 185
R442 VDD1.n76 VDD1.n75 185
R443 VDD1.n65 VDD1.n64 185
R444 VDD1.n82 VDD1.n81 185
R445 VDD1.n84 VDD1.n83 185
R446 VDD1.n61 VDD1.n60 185
R447 VDD1.n91 VDD1.n90 185
R448 VDD1.n92 VDD1.n59 185
R449 VDD1.n94 VDD1.n93 185
R450 VDD1.n57 VDD1.n56 185
R451 VDD1.n100 VDD1.n99 185
R452 VDD1.n102 VDD1.n101 185
R453 VDD1.n18 VDD1.t5 149.524
R454 VDD1.n70 VDD1.t4 149.524
R455 VDD1.n48 VDD1.n47 104.615
R456 VDD1.n47 VDD1.n3 104.615
R457 VDD1.n40 VDD1.n3 104.615
R458 VDD1.n40 VDD1.n39 104.615
R459 VDD1.n39 VDD1.n38 104.615
R460 VDD1.n38 VDD1.n7 104.615
R461 VDD1.n31 VDD1.n7 104.615
R462 VDD1.n31 VDD1.n30 104.615
R463 VDD1.n30 VDD1.n12 104.615
R464 VDD1.n23 VDD1.n12 104.615
R465 VDD1.n23 VDD1.n22 104.615
R466 VDD1.n22 VDD1.n16 104.615
R467 VDD1.n74 VDD1.n68 104.615
R468 VDD1.n75 VDD1.n74 104.615
R469 VDD1.n75 VDD1.n64 104.615
R470 VDD1.n82 VDD1.n64 104.615
R471 VDD1.n83 VDD1.n82 104.615
R472 VDD1.n83 VDD1.n60 104.615
R473 VDD1.n91 VDD1.n60 104.615
R474 VDD1.n92 VDD1.n91 104.615
R475 VDD1.n93 VDD1.n92 104.615
R476 VDD1.n93 VDD1.n56 104.615
R477 VDD1.n100 VDD1.n56 104.615
R478 VDD1.n101 VDD1.n100 104.615
R479 VDD1.n107 VDD1.n106 63.7356
R480 VDD1.n109 VDD1.n108 63.028
R481 VDD1.t5 VDD1.n16 52.3082
R482 VDD1.t4 VDD1.n68 52.3082
R483 VDD1 VDD1.n52 51.599
R484 VDD1.n107 VDD1.n105 51.4855
R485 VDD1.n109 VDD1.n107 44.3457
R486 VDD1.n41 VDD1.n6 13.1884
R487 VDD1.n94 VDD1.n59 13.1884
R488 VDD1.n42 VDD1.n4 12.8005
R489 VDD1.n37 VDD1.n8 12.8005
R490 VDD1.n90 VDD1.n89 12.8005
R491 VDD1.n95 VDD1.n57 12.8005
R492 VDD1.n46 VDD1.n45 12.0247
R493 VDD1.n36 VDD1.n9 12.0247
R494 VDD1.n88 VDD1.n61 12.0247
R495 VDD1.n99 VDD1.n98 12.0247
R496 VDD1.n49 VDD1.n2 11.249
R497 VDD1.n33 VDD1.n32 11.249
R498 VDD1.n85 VDD1.n84 11.249
R499 VDD1.n102 VDD1.n55 11.249
R500 VDD1.n50 VDD1.n0 10.4732
R501 VDD1.n29 VDD1.n11 10.4732
R502 VDD1.n81 VDD1.n63 10.4732
R503 VDD1.n103 VDD1.n53 10.4732
R504 VDD1.n18 VDD1.n17 10.2747
R505 VDD1.n70 VDD1.n69 10.2747
R506 VDD1.n28 VDD1.n13 9.69747
R507 VDD1.n80 VDD1.n65 9.69747
R508 VDD1.n52 VDD1.n51 9.45567
R509 VDD1.n105 VDD1.n104 9.45567
R510 VDD1.n20 VDD1.n19 9.3005
R511 VDD1.n15 VDD1.n14 9.3005
R512 VDD1.n26 VDD1.n25 9.3005
R513 VDD1.n28 VDD1.n27 9.3005
R514 VDD1.n11 VDD1.n10 9.3005
R515 VDD1.n34 VDD1.n33 9.3005
R516 VDD1.n36 VDD1.n35 9.3005
R517 VDD1.n8 VDD1.n5 9.3005
R518 VDD1.n51 VDD1.n50 9.3005
R519 VDD1.n2 VDD1.n1 9.3005
R520 VDD1.n45 VDD1.n44 9.3005
R521 VDD1.n43 VDD1.n42 9.3005
R522 VDD1.n104 VDD1.n103 9.3005
R523 VDD1.n55 VDD1.n54 9.3005
R524 VDD1.n98 VDD1.n97 9.3005
R525 VDD1.n96 VDD1.n95 9.3005
R526 VDD1.n72 VDD1.n71 9.3005
R527 VDD1.n67 VDD1.n66 9.3005
R528 VDD1.n78 VDD1.n77 9.3005
R529 VDD1.n80 VDD1.n79 9.3005
R530 VDD1.n63 VDD1.n62 9.3005
R531 VDD1.n86 VDD1.n85 9.3005
R532 VDD1.n88 VDD1.n87 9.3005
R533 VDD1.n89 VDD1.n58 9.3005
R534 VDD1.n25 VDD1.n24 8.92171
R535 VDD1.n77 VDD1.n76 8.92171
R536 VDD1.n21 VDD1.n15 8.14595
R537 VDD1.n73 VDD1.n67 8.14595
R538 VDD1.n20 VDD1.n17 7.3702
R539 VDD1.n72 VDD1.n69 7.3702
R540 VDD1.n21 VDD1.n20 5.81868
R541 VDD1.n73 VDD1.n72 5.81868
R542 VDD1.n24 VDD1.n15 5.04292
R543 VDD1.n76 VDD1.n67 5.04292
R544 VDD1.n25 VDD1.n13 4.26717
R545 VDD1.n77 VDD1.n65 4.26717
R546 VDD1.n52 VDD1.n0 3.49141
R547 VDD1.n29 VDD1.n28 3.49141
R548 VDD1.n81 VDD1.n80 3.49141
R549 VDD1.n105 VDD1.n53 3.49141
R550 VDD1.n19 VDD1.n18 2.84303
R551 VDD1.n71 VDD1.n70 2.84303
R552 VDD1.n50 VDD1.n49 2.71565
R553 VDD1.n32 VDD1.n11 2.71565
R554 VDD1.n84 VDD1.n63 2.71565
R555 VDD1.n103 VDD1.n102 2.71565
R556 VDD1.n108 VDD1.t3 1.98447
R557 VDD1.n108 VDD1.t2 1.98447
R558 VDD1.n106 VDD1.t1 1.98447
R559 VDD1.n106 VDD1.t0 1.98447
R560 VDD1.n46 VDD1.n2 1.93989
R561 VDD1.n33 VDD1.n9 1.93989
R562 VDD1.n85 VDD1.n61 1.93989
R563 VDD1.n99 VDD1.n55 1.93989
R564 VDD1.n45 VDD1.n4 1.16414
R565 VDD1.n37 VDD1.n36 1.16414
R566 VDD1.n90 VDD1.n88 1.16414
R567 VDD1.n98 VDD1.n57 1.16414
R568 VDD1 VDD1.n109 0.705241
R569 VDD1.n42 VDD1.n41 0.388379
R570 VDD1.n8 VDD1.n6 0.388379
R571 VDD1.n89 VDD1.n59 0.388379
R572 VDD1.n95 VDD1.n94 0.388379
R573 VDD1.n51 VDD1.n1 0.155672
R574 VDD1.n44 VDD1.n1 0.155672
R575 VDD1.n44 VDD1.n43 0.155672
R576 VDD1.n43 VDD1.n5 0.155672
R577 VDD1.n35 VDD1.n5 0.155672
R578 VDD1.n35 VDD1.n34 0.155672
R579 VDD1.n34 VDD1.n10 0.155672
R580 VDD1.n27 VDD1.n10 0.155672
R581 VDD1.n27 VDD1.n26 0.155672
R582 VDD1.n26 VDD1.n14 0.155672
R583 VDD1.n19 VDD1.n14 0.155672
R584 VDD1.n71 VDD1.n66 0.155672
R585 VDD1.n78 VDD1.n66 0.155672
R586 VDD1.n79 VDD1.n78 0.155672
R587 VDD1.n79 VDD1.n62 0.155672
R588 VDD1.n86 VDD1.n62 0.155672
R589 VDD1.n87 VDD1.n86 0.155672
R590 VDD1.n87 VDD1.n58 0.155672
R591 VDD1.n96 VDD1.n58 0.155672
R592 VDD1.n97 VDD1.n96 0.155672
R593 VDD1.n97 VDD1.n54 0.155672
R594 VDD1.n104 VDD1.n54 0.155672
R595 B.n814 B.n813 585
R596 B.n815 B.n814 585
R597 B.n297 B.n132 585
R598 B.n296 B.n295 585
R599 B.n294 B.n293 585
R600 B.n292 B.n291 585
R601 B.n290 B.n289 585
R602 B.n288 B.n287 585
R603 B.n286 B.n285 585
R604 B.n284 B.n283 585
R605 B.n282 B.n281 585
R606 B.n280 B.n279 585
R607 B.n278 B.n277 585
R608 B.n276 B.n275 585
R609 B.n274 B.n273 585
R610 B.n272 B.n271 585
R611 B.n270 B.n269 585
R612 B.n268 B.n267 585
R613 B.n266 B.n265 585
R614 B.n264 B.n263 585
R615 B.n262 B.n261 585
R616 B.n260 B.n259 585
R617 B.n258 B.n257 585
R618 B.n256 B.n255 585
R619 B.n254 B.n253 585
R620 B.n252 B.n251 585
R621 B.n250 B.n249 585
R622 B.n248 B.n247 585
R623 B.n246 B.n245 585
R624 B.n244 B.n243 585
R625 B.n242 B.n241 585
R626 B.n240 B.n239 585
R627 B.n238 B.n237 585
R628 B.n236 B.n235 585
R629 B.n234 B.n233 585
R630 B.n232 B.n231 585
R631 B.n230 B.n229 585
R632 B.n227 B.n226 585
R633 B.n225 B.n224 585
R634 B.n223 B.n222 585
R635 B.n221 B.n220 585
R636 B.n219 B.n218 585
R637 B.n217 B.n216 585
R638 B.n215 B.n214 585
R639 B.n213 B.n212 585
R640 B.n211 B.n210 585
R641 B.n209 B.n208 585
R642 B.n207 B.n206 585
R643 B.n205 B.n204 585
R644 B.n203 B.n202 585
R645 B.n201 B.n200 585
R646 B.n199 B.n198 585
R647 B.n197 B.n196 585
R648 B.n195 B.n194 585
R649 B.n193 B.n192 585
R650 B.n191 B.n190 585
R651 B.n189 B.n188 585
R652 B.n187 B.n186 585
R653 B.n185 B.n184 585
R654 B.n183 B.n182 585
R655 B.n181 B.n180 585
R656 B.n179 B.n178 585
R657 B.n177 B.n176 585
R658 B.n175 B.n174 585
R659 B.n173 B.n172 585
R660 B.n171 B.n170 585
R661 B.n169 B.n168 585
R662 B.n167 B.n166 585
R663 B.n165 B.n164 585
R664 B.n163 B.n162 585
R665 B.n161 B.n160 585
R666 B.n159 B.n158 585
R667 B.n157 B.n156 585
R668 B.n155 B.n154 585
R669 B.n153 B.n152 585
R670 B.n151 B.n150 585
R671 B.n149 B.n148 585
R672 B.n147 B.n146 585
R673 B.n145 B.n144 585
R674 B.n143 B.n142 585
R675 B.n141 B.n140 585
R676 B.n139 B.n138 585
R677 B.n812 B.n91 585
R678 B.n816 B.n91 585
R679 B.n811 B.n90 585
R680 B.n817 B.n90 585
R681 B.n810 B.n809 585
R682 B.n809 B.n86 585
R683 B.n808 B.n85 585
R684 B.n823 B.n85 585
R685 B.n807 B.n84 585
R686 B.n824 B.n84 585
R687 B.n806 B.n83 585
R688 B.n825 B.n83 585
R689 B.n805 B.n804 585
R690 B.n804 B.n79 585
R691 B.n803 B.n78 585
R692 B.n831 B.n78 585
R693 B.n802 B.n77 585
R694 B.n832 B.n77 585
R695 B.n801 B.n76 585
R696 B.n833 B.n76 585
R697 B.n800 B.n799 585
R698 B.n799 B.n72 585
R699 B.n798 B.n71 585
R700 B.n839 B.n71 585
R701 B.n797 B.n70 585
R702 B.n840 B.n70 585
R703 B.n796 B.n69 585
R704 B.n841 B.n69 585
R705 B.n795 B.n794 585
R706 B.n794 B.n65 585
R707 B.n793 B.n64 585
R708 B.n847 B.n64 585
R709 B.n792 B.n63 585
R710 B.n848 B.n63 585
R711 B.n791 B.n62 585
R712 B.n849 B.n62 585
R713 B.n790 B.n789 585
R714 B.n789 B.n58 585
R715 B.n788 B.n57 585
R716 B.n855 B.n57 585
R717 B.n787 B.n56 585
R718 B.n856 B.n56 585
R719 B.n786 B.n55 585
R720 B.n857 B.n55 585
R721 B.n785 B.n784 585
R722 B.n784 B.n51 585
R723 B.n783 B.n50 585
R724 B.n863 B.n50 585
R725 B.n782 B.n49 585
R726 B.n864 B.n49 585
R727 B.n781 B.n48 585
R728 B.n865 B.n48 585
R729 B.n780 B.n779 585
R730 B.n779 B.n44 585
R731 B.n778 B.n43 585
R732 B.n871 B.n43 585
R733 B.n777 B.n42 585
R734 B.n872 B.n42 585
R735 B.n776 B.n41 585
R736 B.n873 B.n41 585
R737 B.n775 B.n774 585
R738 B.n774 B.n37 585
R739 B.n773 B.n36 585
R740 B.n879 B.n36 585
R741 B.n772 B.n35 585
R742 B.n880 B.n35 585
R743 B.n771 B.n34 585
R744 B.n881 B.n34 585
R745 B.n770 B.n769 585
R746 B.n769 B.n30 585
R747 B.n768 B.n29 585
R748 B.n887 B.n29 585
R749 B.n767 B.n28 585
R750 B.n888 B.n28 585
R751 B.n766 B.n27 585
R752 B.n889 B.n27 585
R753 B.n765 B.n764 585
R754 B.n764 B.n23 585
R755 B.n763 B.n22 585
R756 B.n895 B.n22 585
R757 B.n762 B.n21 585
R758 B.n896 B.n21 585
R759 B.n761 B.n20 585
R760 B.n897 B.n20 585
R761 B.n760 B.n759 585
R762 B.n759 B.n19 585
R763 B.n758 B.n15 585
R764 B.n903 B.n15 585
R765 B.n757 B.n14 585
R766 B.n904 B.n14 585
R767 B.n756 B.n13 585
R768 B.n905 B.n13 585
R769 B.n755 B.n754 585
R770 B.n754 B.n12 585
R771 B.n753 B.n752 585
R772 B.n753 B.n8 585
R773 B.n751 B.n7 585
R774 B.n912 B.n7 585
R775 B.n750 B.n6 585
R776 B.n913 B.n6 585
R777 B.n749 B.n5 585
R778 B.n914 B.n5 585
R779 B.n748 B.n747 585
R780 B.n747 B.n4 585
R781 B.n746 B.n298 585
R782 B.n746 B.n745 585
R783 B.n736 B.n299 585
R784 B.n300 B.n299 585
R785 B.n738 B.n737 585
R786 B.n739 B.n738 585
R787 B.n735 B.n305 585
R788 B.n305 B.n304 585
R789 B.n734 B.n733 585
R790 B.n733 B.n732 585
R791 B.n307 B.n306 585
R792 B.n725 B.n307 585
R793 B.n724 B.n723 585
R794 B.n726 B.n724 585
R795 B.n722 B.n312 585
R796 B.n312 B.n311 585
R797 B.n721 B.n720 585
R798 B.n720 B.n719 585
R799 B.n314 B.n313 585
R800 B.n315 B.n314 585
R801 B.n712 B.n711 585
R802 B.n713 B.n712 585
R803 B.n710 B.n320 585
R804 B.n320 B.n319 585
R805 B.n709 B.n708 585
R806 B.n708 B.n707 585
R807 B.n322 B.n321 585
R808 B.n323 B.n322 585
R809 B.n700 B.n699 585
R810 B.n701 B.n700 585
R811 B.n698 B.n327 585
R812 B.n331 B.n327 585
R813 B.n697 B.n696 585
R814 B.n696 B.n695 585
R815 B.n329 B.n328 585
R816 B.n330 B.n329 585
R817 B.n688 B.n687 585
R818 B.n689 B.n688 585
R819 B.n686 B.n336 585
R820 B.n336 B.n335 585
R821 B.n685 B.n684 585
R822 B.n684 B.n683 585
R823 B.n338 B.n337 585
R824 B.n339 B.n338 585
R825 B.n676 B.n675 585
R826 B.n677 B.n676 585
R827 B.n674 B.n344 585
R828 B.n344 B.n343 585
R829 B.n673 B.n672 585
R830 B.n672 B.n671 585
R831 B.n346 B.n345 585
R832 B.n347 B.n346 585
R833 B.n664 B.n663 585
R834 B.n665 B.n664 585
R835 B.n662 B.n352 585
R836 B.n352 B.n351 585
R837 B.n661 B.n660 585
R838 B.n660 B.n659 585
R839 B.n354 B.n353 585
R840 B.n355 B.n354 585
R841 B.n652 B.n651 585
R842 B.n653 B.n652 585
R843 B.n650 B.n360 585
R844 B.n360 B.n359 585
R845 B.n649 B.n648 585
R846 B.n648 B.n647 585
R847 B.n362 B.n361 585
R848 B.n363 B.n362 585
R849 B.n640 B.n639 585
R850 B.n641 B.n640 585
R851 B.n638 B.n368 585
R852 B.n368 B.n367 585
R853 B.n637 B.n636 585
R854 B.n636 B.n635 585
R855 B.n370 B.n369 585
R856 B.n371 B.n370 585
R857 B.n628 B.n627 585
R858 B.n629 B.n628 585
R859 B.n626 B.n375 585
R860 B.n379 B.n375 585
R861 B.n625 B.n624 585
R862 B.n624 B.n623 585
R863 B.n377 B.n376 585
R864 B.n378 B.n377 585
R865 B.n616 B.n615 585
R866 B.n617 B.n616 585
R867 B.n614 B.n384 585
R868 B.n384 B.n383 585
R869 B.n613 B.n612 585
R870 B.n612 B.n611 585
R871 B.n386 B.n385 585
R872 B.n387 B.n386 585
R873 B.n604 B.n603 585
R874 B.n605 B.n604 585
R875 B.n602 B.n392 585
R876 B.n392 B.n391 585
R877 B.n596 B.n595 585
R878 B.n594 B.n434 585
R879 B.n593 B.n433 585
R880 B.n598 B.n433 585
R881 B.n592 B.n591 585
R882 B.n590 B.n589 585
R883 B.n588 B.n587 585
R884 B.n586 B.n585 585
R885 B.n584 B.n583 585
R886 B.n582 B.n581 585
R887 B.n580 B.n579 585
R888 B.n578 B.n577 585
R889 B.n576 B.n575 585
R890 B.n574 B.n573 585
R891 B.n572 B.n571 585
R892 B.n570 B.n569 585
R893 B.n568 B.n567 585
R894 B.n566 B.n565 585
R895 B.n564 B.n563 585
R896 B.n562 B.n561 585
R897 B.n560 B.n559 585
R898 B.n558 B.n557 585
R899 B.n556 B.n555 585
R900 B.n554 B.n553 585
R901 B.n552 B.n551 585
R902 B.n550 B.n549 585
R903 B.n548 B.n547 585
R904 B.n546 B.n545 585
R905 B.n544 B.n543 585
R906 B.n542 B.n541 585
R907 B.n540 B.n539 585
R908 B.n538 B.n537 585
R909 B.n536 B.n535 585
R910 B.n534 B.n533 585
R911 B.n532 B.n531 585
R912 B.n530 B.n529 585
R913 B.n528 B.n527 585
R914 B.n525 B.n524 585
R915 B.n523 B.n522 585
R916 B.n521 B.n520 585
R917 B.n519 B.n518 585
R918 B.n517 B.n516 585
R919 B.n515 B.n514 585
R920 B.n513 B.n512 585
R921 B.n511 B.n510 585
R922 B.n509 B.n508 585
R923 B.n507 B.n506 585
R924 B.n505 B.n504 585
R925 B.n503 B.n502 585
R926 B.n501 B.n500 585
R927 B.n499 B.n498 585
R928 B.n497 B.n496 585
R929 B.n495 B.n494 585
R930 B.n493 B.n492 585
R931 B.n491 B.n490 585
R932 B.n489 B.n488 585
R933 B.n487 B.n486 585
R934 B.n485 B.n484 585
R935 B.n483 B.n482 585
R936 B.n481 B.n480 585
R937 B.n479 B.n478 585
R938 B.n477 B.n476 585
R939 B.n475 B.n474 585
R940 B.n473 B.n472 585
R941 B.n471 B.n470 585
R942 B.n469 B.n468 585
R943 B.n467 B.n466 585
R944 B.n465 B.n464 585
R945 B.n463 B.n462 585
R946 B.n461 B.n460 585
R947 B.n459 B.n458 585
R948 B.n457 B.n456 585
R949 B.n455 B.n454 585
R950 B.n453 B.n452 585
R951 B.n451 B.n450 585
R952 B.n449 B.n448 585
R953 B.n447 B.n446 585
R954 B.n445 B.n444 585
R955 B.n443 B.n442 585
R956 B.n441 B.n440 585
R957 B.n394 B.n393 585
R958 B.n601 B.n600 585
R959 B.n390 B.n389 585
R960 B.n391 B.n390 585
R961 B.n607 B.n606 585
R962 B.n606 B.n605 585
R963 B.n608 B.n388 585
R964 B.n388 B.n387 585
R965 B.n610 B.n609 585
R966 B.n611 B.n610 585
R967 B.n382 B.n381 585
R968 B.n383 B.n382 585
R969 B.n619 B.n618 585
R970 B.n618 B.n617 585
R971 B.n620 B.n380 585
R972 B.n380 B.n378 585
R973 B.n622 B.n621 585
R974 B.n623 B.n622 585
R975 B.n374 B.n373 585
R976 B.n379 B.n374 585
R977 B.n631 B.n630 585
R978 B.n630 B.n629 585
R979 B.n632 B.n372 585
R980 B.n372 B.n371 585
R981 B.n634 B.n633 585
R982 B.n635 B.n634 585
R983 B.n366 B.n365 585
R984 B.n367 B.n366 585
R985 B.n643 B.n642 585
R986 B.n642 B.n641 585
R987 B.n644 B.n364 585
R988 B.n364 B.n363 585
R989 B.n646 B.n645 585
R990 B.n647 B.n646 585
R991 B.n358 B.n357 585
R992 B.n359 B.n358 585
R993 B.n655 B.n654 585
R994 B.n654 B.n653 585
R995 B.n656 B.n356 585
R996 B.n356 B.n355 585
R997 B.n658 B.n657 585
R998 B.n659 B.n658 585
R999 B.n350 B.n349 585
R1000 B.n351 B.n350 585
R1001 B.n667 B.n666 585
R1002 B.n666 B.n665 585
R1003 B.n668 B.n348 585
R1004 B.n348 B.n347 585
R1005 B.n670 B.n669 585
R1006 B.n671 B.n670 585
R1007 B.n342 B.n341 585
R1008 B.n343 B.n342 585
R1009 B.n679 B.n678 585
R1010 B.n678 B.n677 585
R1011 B.n680 B.n340 585
R1012 B.n340 B.n339 585
R1013 B.n682 B.n681 585
R1014 B.n683 B.n682 585
R1015 B.n334 B.n333 585
R1016 B.n335 B.n334 585
R1017 B.n691 B.n690 585
R1018 B.n690 B.n689 585
R1019 B.n692 B.n332 585
R1020 B.n332 B.n330 585
R1021 B.n694 B.n693 585
R1022 B.n695 B.n694 585
R1023 B.n326 B.n325 585
R1024 B.n331 B.n326 585
R1025 B.n703 B.n702 585
R1026 B.n702 B.n701 585
R1027 B.n704 B.n324 585
R1028 B.n324 B.n323 585
R1029 B.n706 B.n705 585
R1030 B.n707 B.n706 585
R1031 B.n318 B.n317 585
R1032 B.n319 B.n318 585
R1033 B.n715 B.n714 585
R1034 B.n714 B.n713 585
R1035 B.n716 B.n316 585
R1036 B.n316 B.n315 585
R1037 B.n718 B.n717 585
R1038 B.n719 B.n718 585
R1039 B.n310 B.n309 585
R1040 B.n311 B.n310 585
R1041 B.n728 B.n727 585
R1042 B.n727 B.n726 585
R1043 B.n729 B.n308 585
R1044 B.n725 B.n308 585
R1045 B.n731 B.n730 585
R1046 B.n732 B.n731 585
R1047 B.n303 B.n302 585
R1048 B.n304 B.n303 585
R1049 B.n741 B.n740 585
R1050 B.n740 B.n739 585
R1051 B.n742 B.n301 585
R1052 B.n301 B.n300 585
R1053 B.n744 B.n743 585
R1054 B.n745 B.n744 585
R1055 B.n3 B.n0 585
R1056 B.n4 B.n3 585
R1057 B.n911 B.n1 585
R1058 B.n912 B.n911 585
R1059 B.n910 B.n909 585
R1060 B.n910 B.n8 585
R1061 B.n908 B.n9 585
R1062 B.n12 B.n9 585
R1063 B.n907 B.n906 585
R1064 B.n906 B.n905 585
R1065 B.n11 B.n10 585
R1066 B.n904 B.n11 585
R1067 B.n902 B.n901 585
R1068 B.n903 B.n902 585
R1069 B.n900 B.n16 585
R1070 B.n19 B.n16 585
R1071 B.n899 B.n898 585
R1072 B.n898 B.n897 585
R1073 B.n18 B.n17 585
R1074 B.n896 B.n18 585
R1075 B.n894 B.n893 585
R1076 B.n895 B.n894 585
R1077 B.n892 B.n24 585
R1078 B.n24 B.n23 585
R1079 B.n891 B.n890 585
R1080 B.n890 B.n889 585
R1081 B.n26 B.n25 585
R1082 B.n888 B.n26 585
R1083 B.n886 B.n885 585
R1084 B.n887 B.n886 585
R1085 B.n884 B.n31 585
R1086 B.n31 B.n30 585
R1087 B.n883 B.n882 585
R1088 B.n882 B.n881 585
R1089 B.n33 B.n32 585
R1090 B.n880 B.n33 585
R1091 B.n878 B.n877 585
R1092 B.n879 B.n878 585
R1093 B.n876 B.n38 585
R1094 B.n38 B.n37 585
R1095 B.n875 B.n874 585
R1096 B.n874 B.n873 585
R1097 B.n40 B.n39 585
R1098 B.n872 B.n40 585
R1099 B.n870 B.n869 585
R1100 B.n871 B.n870 585
R1101 B.n868 B.n45 585
R1102 B.n45 B.n44 585
R1103 B.n867 B.n866 585
R1104 B.n866 B.n865 585
R1105 B.n47 B.n46 585
R1106 B.n864 B.n47 585
R1107 B.n862 B.n861 585
R1108 B.n863 B.n862 585
R1109 B.n860 B.n52 585
R1110 B.n52 B.n51 585
R1111 B.n859 B.n858 585
R1112 B.n858 B.n857 585
R1113 B.n54 B.n53 585
R1114 B.n856 B.n54 585
R1115 B.n854 B.n853 585
R1116 B.n855 B.n854 585
R1117 B.n852 B.n59 585
R1118 B.n59 B.n58 585
R1119 B.n851 B.n850 585
R1120 B.n850 B.n849 585
R1121 B.n61 B.n60 585
R1122 B.n848 B.n61 585
R1123 B.n846 B.n845 585
R1124 B.n847 B.n846 585
R1125 B.n844 B.n66 585
R1126 B.n66 B.n65 585
R1127 B.n843 B.n842 585
R1128 B.n842 B.n841 585
R1129 B.n68 B.n67 585
R1130 B.n840 B.n68 585
R1131 B.n838 B.n837 585
R1132 B.n839 B.n838 585
R1133 B.n836 B.n73 585
R1134 B.n73 B.n72 585
R1135 B.n835 B.n834 585
R1136 B.n834 B.n833 585
R1137 B.n75 B.n74 585
R1138 B.n832 B.n75 585
R1139 B.n830 B.n829 585
R1140 B.n831 B.n830 585
R1141 B.n828 B.n80 585
R1142 B.n80 B.n79 585
R1143 B.n827 B.n826 585
R1144 B.n826 B.n825 585
R1145 B.n82 B.n81 585
R1146 B.n824 B.n82 585
R1147 B.n822 B.n821 585
R1148 B.n823 B.n822 585
R1149 B.n820 B.n87 585
R1150 B.n87 B.n86 585
R1151 B.n819 B.n818 585
R1152 B.n818 B.n817 585
R1153 B.n89 B.n88 585
R1154 B.n816 B.n89 585
R1155 B.n915 B.n914 585
R1156 B.n913 B.n2 585
R1157 B.n138 B.n89 535.745
R1158 B.n814 B.n91 535.745
R1159 B.n600 B.n392 535.745
R1160 B.n596 B.n390 535.745
R1161 B.n133 B.t15 315.913
R1162 B.n437 B.t12 315.913
R1163 B.n135 B.t18 315.913
R1164 B.n435 B.t9 315.913
R1165 B.n135 B.t17 283.741
R1166 B.n133 B.t13 283.741
R1167 B.n437 B.t10 283.741
R1168 B.n435 B.t6 283.741
R1169 B.n815 B.n131 256.663
R1170 B.n815 B.n130 256.663
R1171 B.n815 B.n129 256.663
R1172 B.n815 B.n128 256.663
R1173 B.n815 B.n127 256.663
R1174 B.n815 B.n126 256.663
R1175 B.n815 B.n125 256.663
R1176 B.n815 B.n124 256.663
R1177 B.n815 B.n123 256.663
R1178 B.n815 B.n122 256.663
R1179 B.n815 B.n121 256.663
R1180 B.n815 B.n120 256.663
R1181 B.n815 B.n119 256.663
R1182 B.n815 B.n118 256.663
R1183 B.n815 B.n117 256.663
R1184 B.n815 B.n116 256.663
R1185 B.n815 B.n115 256.663
R1186 B.n815 B.n114 256.663
R1187 B.n815 B.n113 256.663
R1188 B.n815 B.n112 256.663
R1189 B.n815 B.n111 256.663
R1190 B.n815 B.n110 256.663
R1191 B.n815 B.n109 256.663
R1192 B.n815 B.n108 256.663
R1193 B.n815 B.n107 256.663
R1194 B.n815 B.n106 256.663
R1195 B.n815 B.n105 256.663
R1196 B.n815 B.n104 256.663
R1197 B.n815 B.n103 256.663
R1198 B.n815 B.n102 256.663
R1199 B.n815 B.n101 256.663
R1200 B.n815 B.n100 256.663
R1201 B.n815 B.n99 256.663
R1202 B.n815 B.n98 256.663
R1203 B.n815 B.n97 256.663
R1204 B.n815 B.n96 256.663
R1205 B.n815 B.n95 256.663
R1206 B.n815 B.n94 256.663
R1207 B.n815 B.n93 256.663
R1208 B.n815 B.n92 256.663
R1209 B.n598 B.n597 256.663
R1210 B.n598 B.n395 256.663
R1211 B.n598 B.n396 256.663
R1212 B.n598 B.n397 256.663
R1213 B.n598 B.n398 256.663
R1214 B.n598 B.n399 256.663
R1215 B.n598 B.n400 256.663
R1216 B.n598 B.n401 256.663
R1217 B.n598 B.n402 256.663
R1218 B.n598 B.n403 256.663
R1219 B.n598 B.n404 256.663
R1220 B.n598 B.n405 256.663
R1221 B.n598 B.n406 256.663
R1222 B.n598 B.n407 256.663
R1223 B.n598 B.n408 256.663
R1224 B.n598 B.n409 256.663
R1225 B.n598 B.n410 256.663
R1226 B.n598 B.n411 256.663
R1227 B.n598 B.n412 256.663
R1228 B.n598 B.n413 256.663
R1229 B.n598 B.n414 256.663
R1230 B.n598 B.n415 256.663
R1231 B.n598 B.n416 256.663
R1232 B.n598 B.n417 256.663
R1233 B.n598 B.n418 256.663
R1234 B.n598 B.n419 256.663
R1235 B.n598 B.n420 256.663
R1236 B.n598 B.n421 256.663
R1237 B.n598 B.n422 256.663
R1238 B.n598 B.n423 256.663
R1239 B.n598 B.n424 256.663
R1240 B.n598 B.n425 256.663
R1241 B.n598 B.n426 256.663
R1242 B.n598 B.n427 256.663
R1243 B.n598 B.n428 256.663
R1244 B.n598 B.n429 256.663
R1245 B.n598 B.n430 256.663
R1246 B.n598 B.n431 256.663
R1247 B.n598 B.n432 256.663
R1248 B.n599 B.n598 256.663
R1249 B.n917 B.n916 256.663
R1250 B.n134 B.t16 247.26
R1251 B.n438 B.t11 247.26
R1252 B.n136 B.t19 247.26
R1253 B.n436 B.t8 247.26
R1254 B.n142 B.n141 163.367
R1255 B.n146 B.n145 163.367
R1256 B.n150 B.n149 163.367
R1257 B.n154 B.n153 163.367
R1258 B.n158 B.n157 163.367
R1259 B.n162 B.n161 163.367
R1260 B.n166 B.n165 163.367
R1261 B.n170 B.n169 163.367
R1262 B.n174 B.n173 163.367
R1263 B.n178 B.n177 163.367
R1264 B.n182 B.n181 163.367
R1265 B.n186 B.n185 163.367
R1266 B.n190 B.n189 163.367
R1267 B.n194 B.n193 163.367
R1268 B.n198 B.n197 163.367
R1269 B.n202 B.n201 163.367
R1270 B.n206 B.n205 163.367
R1271 B.n210 B.n209 163.367
R1272 B.n214 B.n213 163.367
R1273 B.n218 B.n217 163.367
R1274 B.n222 B.n221 163.367
R1275 B.n226 B.n225 163.367
R1276 B.n231 B.n230 163.367
R1277 B.n235 B.n234 163.367
R1278 B.n239 B.n238 163.367
R1279 B.n243 B.n242 163.367
R1280 B.n247 B.n246 163.367
R1281 B.n251 B.n250 163.367
R1282 B.n255 B.n254 163.367
R1283 B.n259 B.n258 163.367
R1284 B.n263 B.n262 163.367
R1285 B.n267 B.n266 163.367
R1286 B.n271 B.n270 163.367
R1287 B.n275 B.n274 163.367
R1288 B.n279 B.n278 163.367
R1289 B.n283 B.n282 163.367
R1290 B.n287 B.n286 163.367
R1291 B.n291 B.n290 163.367
R1292 B.n295 B.n294 163.367
R1293 B.n814 B.n132 163.367
R1294 B.n604 B.n392 163.367
R1295 B.n604 B.n386 163.367
R1296 B.n612 B.n386 163.367
R1297 B.n612 B.n384 163.367
R1298 B.n616 B.n384 163.367
R1299 B.n616 B.n377 163.367
R1300 B.n624 B.n377 163.367
R1301 B.n624 B.n375 163.367
R1302 B.n628 B.n375 163.367
R1303 B.n628 B.n370 163.367
R1304 B.n636 B.n370 163.367
R1305 B.n636 B.n368 163.367
R1306 B.n640 B.n368 163.367
R1307 B.n640 B.n362 163.367
R1308 B.n648 B.n362 163.367
R1309 B.n648 B.n360 163.367
R1310 B.n652 B.n360 163.367
R1311 B.n652 B.n354 163.367
R1312 B.n660 B.n354 163.367
R1313 B.n660 B.n352 163.367
R1314 B.n664 B.n352 163.367
R1315 B.n664 B.n346 163.367
R1316 B.n672 B.n346 163.367
R1317 B.n672 B.n344 163.367
R1318 B.n676 B.n344 163.367
R1319 B.n676 B.n338 163.367
R1320 B.n684 B.n338 163.367
R1321 B.n684 B.n336 163.367
R1322 B.n688 B.n336 163.367
R1323 B.n688 B.n329 163.367
R1324 B.n696 B.n329 163.367
R1325 B.n696 B.n327 163.367
R1326 B.n700 B.n327 163.367
R1327 B.n700 B.n322 163.367
R1328 B.n708 B.n322 163.367
R1329 B.n708 B.n320 163.367
R1330 B.n712 B.n320 163.367
R1331 B.n712 B.n314 163.367
R1332 B.n720 B.n314 163.367
R1333 B.n720 B.n312 163.367
R1334 B.n724 B.n312 163.367
R1335 B.n724 B.n307 163.367
R1336 B.n733 B.n307 163.367
R1337 B.n733 B.n305 163.367
R1338 B.n738 B.n305 163.367
R1339 B.n738 B.n299 163.367
R1340 B.n746 B.n299 163.367
R1341 B.n747 B.n746 163.367
R1342 B.n747 B.n5 163.367
R1343 B.n6 B.n5 163.367
R1344 B.n7 B.n6 163.367
R1345 B.n753 B.n7 163.367
R1346 B.n754 B.n753 163.367
R1347 B.n754 B.n13 163.367
R1348 B.n14 B.n13 163.367
R1349 B.n15 B.n14 163.367
R1350 B.n759 B.n15 163.367
R1351 B.n759 B.n20 163.367
R1352 B.n21 B.n20 163.367
R1353 B.n22 B.n21 163.367
R1354 B.n764 B.n22 163.367
R1355 B.n764 B.n27 163.367
R1356 B.n28 B.n27 163.367
R1357 B.n29 B.n28 163.367
R1358 B.n769 B.n29 163.367
R1359 B.n769 B.n34 163.367
R1360 B.n35 B.n34 163.367
R1361 B.n36 B.n35 163.367
R1362 B.n774 B.n36 163.367
R1363 B.n774 B.n41 163.367
R1364 B.n42 B.n41 163.367
R1365 B.n43 B.n42 163.367
R1366 B.n779 B.n43 163.367
R1367 B.n779 B.n48 163.367
R1368 B.n49 B.n48 163.367
R1369 B.n50 B.n49 163.367
R1370 B.n784 B.n50 163.367
R1371 B.n784 B.n55 163.367
R1372 B.n56 B.n55 163.367
R1373 B.n57 B.n56 163.367
R1374 B.n789 B.n57 163.367
R1375 B.n789 B.n62 163.367
R1376 B.n63 B.n62 163.367
R1377 B.n64 B.n63 163.367
R1378 B.n794 B.n64 163.367
R1379 B.n794 B.n69 163.367
R1380 B.n70 B.n69 163.367
R1381 B.n71 B.n70 163.367
R1382 B.n799 B.n71 163.367
R1383 B.n799 B.n76 163.367
R1384 B.n77 B.n76 163.367
R1385 B.n78 B.n77 163.367
R1386 B.n804 B.n78 163.367
R1387 B.n804 B.n83 163.367
R1388 B.n84 B.n83 163.367
R1389 B.n85 B.n84 163.367
R1390 B.n809 B.n85 163.367
R1391 B.n809 B.n90 163.367
R1392 B.n91 B.n90 163.367
R1393 B.n434 B.n433 163.367
R1394 B.n591 B.n433 163.367
R1395 B.n589 B.n588 163.367
R1396 B.n585 B.n584 163.367
R1397 B.n581 B.n580 163.367
R1398 B.n577 B.n576 163.367
R1399 B.n573 B.n572 163.367
R1400 B.n569 B.n568 163.367
R1401 B.n565 B.n564 163.367
R1402 B.n561 B.n560 163.367
R1403 B.n557 B.n556 163.367
R1404 B.n553 B.n552 163.367
R1405 B.n549 B.n548 163.367
R1406 B.n545 B.n544 163.367
R1407 B.n541 B.n540 163.367
R1408 B.n537 B.n536 163.367
R1409 B.n533 B.n532 163.367
R1410 B.n529 B.n528 163.367
R1411 B.n524 B.n523 163.367
R1412 B.n520 B.n519 163.367
R1413 B.n516 B.n515 163.367
R1414 B.n512 B.n511 163.367
R1415 B.n508 B.n507 163.367
R1416 B.n504 B.n503 163.367
R1417 B.n500 B.n499 163.367
R1418 B.n496 B.n495 163.367
R1419 B.n492 B.n491 163.367
R1420 B.n488 B.n487 163.367
R1421 B.n484 B.n483 163.367
R1422 B.n480 B.n479 163.367
R1423 B.n476 B.n475 163.367
R1424 B.n472 B.n471 163.367
R1425 B.n468 B.n467 163.367
R1426 B.n464 B.n463 163.367
R1427 B.n460 B.n459 163.367
R1428 B.n456 B.n455 163.367
R1429 B.n452 B.n451 163.367
R1430 B.n448 B.n447 163.367
R1431 B.n444 B.n443 163.367
R1432 B.n440 B.n394 163.367
R1433 B.n606 B.n390 163.367
R1434 B.n606 B.n388 163.367
R1435 B.n610 B.n388 163.367
R1436 B.n610 B.n382 163.367
R1437 B.n618 B.n382 163.367
R1438 B.n618 B.n380 163.367
R1439 B.n622 B.n380 163.367
R1440 B.n622 B.n374 163.367
R1441 B.n630 B.n374 163.367
R1442 B.n630 B.n372 163.367
R1443 B.n634 B.n372 163.367
R1444 B.n634 B.n366 163.367
R1445 B.n642 B.n366 163.367
R1446 B.n642 B.n364 163.367
R1447 B.n646 B.n364 163.367
R1448 B.n646 B.n358 163.367
R1449 B.n654 B.n358 163.367
R1450 B.n654 B.n356 163.367
R1451 B.n658 B.n356 163.367
R1452 B.n658 B.n350 163.367
R1453 B.n666 B.n350 163.367
R1454 B.n666 B.n348 163.367
R1455 B.n670 B.n348 163.367
R1456 B.n670 B.n342 163.367
R1457 B.n678 B.n342 163.367
R1458 B.n678 B.n340 163.367
R1459 B.n682 B.n340 163.367
R1460 B.n682 B.n334 163.367
R1461 B.n690 B.n334 163.367
R1462 B.n690 B.n332 163.367
R1463 B.n694 B.n332 163.367
R1464 B.n694 B.n326 163.367
R1465 B.n702 B.n326 163.367
R1466 B.n702 B.n324 163.367
R1467 B.n706 B.n324 163.367
R1468 B.n706 B.n318 163.367
R1469 B.n714 B.n318 163.367
R1470 B.n714 B.n316 163.367
R1471 B.n718 B.n316 163.367
R1472 B.n718 B.n310 163.367
R1473 B.n727 B.n310 163.367
R1474 B.n727 B.n308 163.367
R1475 B.n731 B.n308 163.367
R1476 B.n731 B.n303 163.367
R1477 B.n740 B.n303 163.367
R1478 B.n740 B.n301 163.367
R1479 B.n744 B.n301 163.367
R1480 B.n744 B.n3 163.367
R1481 B.n915 B.n3 163.367
R1482 B.n911 B.n2 163.367
R1483 B.n911 B.n910 163.367
R1484 B.n910 B.n9 163.367
R1485 B.n906 B.n9 163.367
R1486 B.n906 B.n11 163.367
R1487 B.n902 B.n11 163.367
R1488 B.n902 B.n16 163.367
R1489 B.n898 B.n16 163.367
R1490 B.n898 B.n18 163.367
R1491 B.n894 B.n18 163.367
R1492 B.n894 B.n24 163.367
R1493 B.n890 B.n24 163.367
R1494 B.n890 B.n26 163.367
R1495 B.n886 B.n26 163.367
R1496 B.n886 B.n31 163.367
R1497 B.n882 B.n31 163.367
R1498 B.n882 B.n33 163.367
R1499 B.n878 B.n33 163.367
R1500 B.n878 B.n38 163.367
R1501 B.n874 B.n38 163.367
R1502 B.n874 B.n40 163.367
R1503 B.n870 B.n40 163.367
R1504 B.n870 B.n45 163.367
R1505 B.n866 B.n45 163.367
R1506 B.n866 B.n47 163.367
R1507 B.n862 B.n47 163.367
R1508 B.n862 B.n52 163.367
R1509 B.n858 B.n52 163.367
R1510 B.n858 B.n54 163.367
R1511 B.n854 B.n54 163.367
R1512 B.n854 B.n59 163.367
R1513 B.n850 B.n59 163.367
R1514 B.n850 B.n61 163.367
R1515 B.n846 B.n61 163.367
R1516 B.n846 B.n66 163.367
R1517 B.n842 B.n66 163.367
R1518 B.n842 B.n68 163.367
R1519 B.n838 B.n68 163.367
R1520 B.n838 B.n73 163.367
R1521 B.n834 B.n73 163.367
R1522 B.n834 B.n75 163.367
R1523 B.n830 B.n75 163.367
R1524 B.n830 B.n80 163.367
R1525 B.n826 B.n80 163.367
R1526 B.n826 B.n82 163.367
R1527 B.n822 B.n82 163.367
R1528 B.n822 B.n87 163.367
R1529 B.n818 B.n87 163.367
R1530 B.n818 B.n89 163.367
R1531 B.n598 B.n391 101.672
R1532 B.n816 B.n815 101.672
R1533 B.n138 B.n92 71.676
R1534 B.n142 B.n93 71.676
R1535 B.n146 B.n94 71.676
R1536 B.n150 B.n95 71.676
R1537 B.n154 B.n96 71.676
R1538 B.n158 B.n97 71.676
R1539 B.n162 B.n98 71.676
R1540 B.n166 B.n99 71.676
R1541 B.n170 B.n100 71.676
R1542 B.n174 B.n101 71.676
R1543 B.n178 B.n102 71.676
R1544 B.n182 B.n103 71.676
R1545 B.n186 B.n104 71.676
R1546 B.n190 B.n105 71.676
R1547 B.n194 B.n106 71.676
R1548 B.n198 B.n107 71.676
R1549 B.n202 B.n108 71.676
R1550 B.n206 B.n109 71.676
R1551 B.n210 B.n110 71.676
R1552 B.n214 B.n111 71.676
R1553 B.n218 B.n112 71.676
R1554 B.n222 B.n113 71.676
R1555 B.n226 B.n114 71.676
R1556 B.n231 B.n115 71.676
R1557 B.n235 B.n116 71.676
R1558 B.n239 B.n117 71.676
R1559 B.n243 B.n118 71.676
R1560 B.n247 B.n119 71.676
R1561 B.n251 B.n120 71.676
R1562 B.n255 B.n121 71.676
R1563 B.n259 B.n122 71.676
R1564 B.n263 B.n123 71.676
R1565 B.n267 B.n124 71.676
R1566 B.n271 B.n125 71.676
R1567 B.n275 B.n126 71.676
R1568 B.n279 B.n127 71.676
R1569 B.n283 B.n128 71.676
R1570 B.n287 B.n129 71.676
R1571 B.n291 B.n130 71.676
R1572 B.n295 B.n131 71.676
R1573 B.n132 B.n131 71.676
R1574 B.n294 B.n130 71.676
R1575 B.n290 B.n129 71.676
R1576 B.n286 B.n128 71.676
R1577 B.n282 B.n127 71.676
R1578 B.n278 B.n126 71.676
R1579 B.n274 B.n125 71.676
R1580 B.n270 B.n124 71.676
R1581 B.n266 B.n123 71.676
R1582 B.n262 B.n122 71.676
R1583 B.n258 B.n121 71.676
R1584 B.n254 B.n120 71.676
R1585 B.n250 B.n119 71.676
R1586 B.n246 B.n118 71.676
R1587 B.n242 B.n117 71.676
R1588 B.n238 B.n116 71.676
R1589 B.n234 B.n115 71.676
R1590 B.n230 B.n114 71.676
R1591 B.n225 B.n113 71.676
R1592 B.n221 B.n112 71.676
R1593 B.n217 B.n111 71.676
R1594 B.n213 B.n110 71.676
R1595 B.n209 B.n109 71.676
R1596 B.n205 B.n108 71.676
R1597 B.n201 B.n107 71.676
R1598 B.n197 B.n106 71.676
R1599 B.n193 B.n105 71.676
R1600 B.n189 B.n104 71.676
R1601 B.n185 B.n103 71.676
R1602 B.n181 B.n102 71.676
R1603 B.n177 B.n101 71.676
R1604 B.n173 B.n100 71.676
R1605 B.n169 B.n99 71.676
R1606 B.n165 B.n98 71.676
R1607 B.n161 B.n97 71.676
R1608 B.n157 B.n96 71.676
R1609 B.n153 B.n95 71.676
R1610 B.n149 B.n94 71.676
R1611 B.n145 B.n93 71.676
R1612 B.n141 B.n92 71.676
R1613 B.n597 B.n596 71.676
R1614 B.n591 B.n395 71.676
R1615 B.n588 B.n396 71.676
R1616 B.n584 B.n397 71.676
R1617 B.n580 B.n398 71.676
R1618 B.n576 B.n399 71.676
R1619 B.n572 B.n400 71.676
R1620 B.n568 B.n401 71.676
R1621 B.n564 B.n402 71.676
R1622 B.n560 B.n403 71.676
R1623 B.n556 B.n404 71.676
R1624 B.n552 B.n405 71.676
R1625 B.n548 B.n406 71.676
R1626 B.n544 B.n407 71.676
R1627 B.n540 B.n408 71.676
R1628 B.n536 B.n409 71.676
R1629 B.n532 B.n410 71.676
R1630 B.n528 B.n411 71.676
R1631 B.n523 B.n412 71.676
R1632 B.n519 B.n413 71.676
R1633 B.n515 B.n414 71.676
R1634 B.n511 B.n415 71.676
R1635 B.n507 B.n416 71.676
R1636 B.n503 B.n417 71.676
R1637 B.n499 B.n418 71.676
R1638 B.n495 B.n419 71.676
R1639 B.n491 B.n420 71.676
R1640 B.n487 B.n421 71.676
R1641 B.n483 B.n422 71.676
R1642 B.n479 B.n423 71.676
R1643 B.n475 B.n424 71.676
R1644 B.n471 B.n425 71.676
R1645 B.n467 B.n426 71.676
R1646 B.n463 B.n427 71.676
R1647 B.n459 B.n428 71.676
R1648 B.n455 B.n429 71.676
R1649 B.n451 B.n430 71.676
R1650 B.n447 B.n431 71.676
R1651 B.n443 B.n432 71.676
R1652 B.n599 B.n394 71.676
R1653 B.n597 B.n434 71.676
R1654 B.n589 B.n395 71.676
R1655 B.n585 B.n396 71.676
R1656 B.n581 B.n397 71.676
R1657 B.n577 B.n398 71.676
R1658 B.n573 B.n399 71.676
R1659 B.n569 B.n400 71.676
R1660 B.n565 B.n401 71.676
R1661 B.n561 B.n402 71.676
R1662 B.n557 B.n403 71.676
R1663 B.n553 B.n404 71.676
R1664 B.n549 B.n405 71.676
R1665 B.n545 B.n406 71.676
R1666 B.n541 B.n407 71.676
R1667 B.n537 B.n408 71.676
R1668 B.n533 B.n409 71.676
R1669 B.n529 B.n410 71.676
R1670 B.n524 B.n411 71.676
R1671 B.n520 B.n412 71.676
R1672 B.n516 B.n413 71.676
R1673 B.n512 B.n414 71.676
R1674 B.n508 B.n415 71.676
R1675 B.n504 B.n416 71.676
R1676 B.n500 B.n417 71.676
R1677 B.n496 B.n418 71.676
R1678 B.n492 B.n419 71.676
R1679 B.n488 B.n420 71.676
R1680 B.n484 B.n421 71.676
R1681 B.n480 B.n422 71.676
R1682 B.n476 B.n423 71.676
R1683 B.n472 B.n424 71.676
R1684 B.n468 B.n425 71.676
R1685 B.n464 B.n426 71.676
R1686 B.n460 B.n427 71.676
R1687 B.n456 B.n428 71.676
R1688 B.n452 B.n429 71.676
R1689 B.n448 B.n430 71.676
R1690 B.n444 B.n431 71.676
R1691 B.n440 B.n432 71.676
R1692 B.n600 B.n599 71.676
R1693 B.n916 B.n915 71.676
R1694 B.n916 B.n2 71.676
R1695 B.n136 B.n135 68.655
R1696 B.n134 B.n133 68.655
R1697 B.n438 B.n437 68.655
R1698 B.n436 B.n435 68.655
R1699 B.n137 B.n136 59.5399
R1700 B.n228 B.n134 59.5399
R1701 B.n439 B.n438 59.5399
R1702 B.n526 B.n436 59.5399
R1703 B.n605 B.n391 49.0336
R1704 B.n605 B.n387 49.0336
R1705 B.n611 B.n387 49.0336
R1706 B.n611 B.n383 49.0336
R1707 B.n617 B.n383 49.0336
R1708 B.n617 B.n378 49.0336
R1709 B.n623 B.n378 49.0336
R1710 B.n623 B.n379 49.0336
R1711 B.n629 B.n371 49.0336
R1712 B.n635 B.n371 49.0336
R1713 B.n635 B.n367 49.0336
R1714 B.n641 B.n367 49.0336
R1715 B.n641 B.n363 49.0336
R1716 B.n647 B.n363 49.0336
R1717 B.n647 B.n359 49.0336
R1718 B.n653 B.n359 49.0336
R1719 B.n653 B.n355 49.0336
R1720 B.n659 B.n355 49.0336
R1721 B.n659 B.n351 49.0336
R1722 B.n665 B.n351 49.0336
R1723 B.n671 B.n347 49.0336
R1724 B.n671 B.n343 49.0336
R1725 B.n677 B.n343 49.0336
R1726 B.n677 B.n339 49.0336
R1727 B.n683 B.n339 49.0336
R1728 B.n683 B.n335 49.0336
R1729 B.n689 B.n335 49.0336
R1730 B.n689 B.n330 49.0336
R1731 B.n695 B.n330 49.0336
R1732 B.n695 B.n331 49.0336
R1733 B.n701 B.n323 49.0336
R1734 B.n707 B.n323 49.0336
R1735 B.n707 B.n319 49.0336
R1736 B.n713 B.n319 49.0336
R1737 B.n713 B.n315 49.0336
R1738 B.n719 B.n315 49.0336
R1739 B.n719 B.n311 49.0336
R1740 B.n726 B.n311 49.0336
R1741 B.n726 B.n725 49.0336
R1742 B.n732 B.n304 49.0336
R1743 B.n739 B.n304 49.0336
R1744 B.n739 B.n300 49.0336
R1745 B.n745 B.n300 49.0336
R1746 B.n745 B.n4 49.0336
R1747 B.n914 B.n4 49.0336
R1748 B.n914 B.n913 49.0336
R1749 B.n913 B.n912 49.0336
R1750 B.n912 B.n8 49.0336
R1751 B.n12 B.n8 49.0336
R1752 B.n905 B.n12 49.0336
R1753 B.n905 B.n904 49.0336
R1754 B.n904 B.n903 49.0336
R1755 B.n897 B.n19 49.0336
R1756 B.n897 B.n896 49.0336
R1757 B.n896 B.n895 49.0336
R1758 B.n895 B.n23 49.0336
R1759 B.n889 B.n23 49.0336
R1760 B.n889 B.n888 49.0336
R1761 B.n888 B.n887 49.0336
R1762 B.n887 B.n30 49.0336
R1763 B.n881 B.n30 49.0336
R1764 B.n880 B.n879 49.0336
R1765 B.n879 B.n37 49.0336
R1766 B.n873 B.n37 49.0336
R1767 B.n873 B.n872 49.0336
R1768 B.n872 B.n871 49.0336
R1769 B.n871 B.n44 49.0336
R1770 B.n865 B.n44 49.0336
R1771 B.n865 B.n864 49.0336
R1772 B.n864 B.n863 49.0336
R1773 B.n863 B.n51 49.0336
R1774 B.n857 B.n856 49.0336
R1775 B.n856 B.n855 49.0336
R1776 B.n855 B.n58 49.0336
R1777 B.n849 B.n58 49.0336
R1778 B.n849 B.n848 49.0336
R1779 B.n848 B.n847 49.0336
R1780 B.n847 B.n65 49.0336
R1781 B.n841 B.n65 49.0336
R1782 B.n841 B.n840 49.0336
R1783 B.n840 B.n839 49.0336
R1784 B.n839 B.n72 49.0336
R1785 B.n833 B.n72 49.0336
R1786 B.n832 B.n831 49.0336
R1787 B.n831 B.n79 49.0336
R1788 B.n825 B.n79 49.0336
R1789 B.n825 B.n824 49.0336
R1790 B.n824 B.n823 49.0336
R1791 B.n823 B.n86 49.0336
R1792 B.n817 B.n86 49.0336
R1793 B.n817 B.n816 49.0336
R1794 B.n665 B.t4 42.5439
R1795 B.n857 B.t3 42.5439
R1796 B.n629 B.t7 36.7753
R1797 B.n833 B.t14 36.7753
R1798 B.n701 B.t0 35.3332
R1799 B.n881 B.t1 35.3332
R1800 B.n595 B.n389 34.8103
R1801 B.n602 B.n601 34.8103
R1802 B.n813 B.n812 34.8103
R1803 B.n139 B.n88 34.8103
R1804 B.n725 B.t5 33.891
R1805 B.n19 B.t2 33.891
R1806 B B.n917 18.0485
R1807 B.n732 B.t5 15.1431
R1808 B.n903 B.t2 15.1431
R1809 B.n331 B.t0 13.7009
R1810 B.t1 B.n880 13.7009
R1811 B.n379 B.t7 12.2588
R1812 B.t14 B.n832 12.2588
R1813 B.n607 B.n389 10.6151
R1814 B.n608 B.n607 10.6151
R1815 B.n609 B.n608 10.6151
R1816 B.n609 B.n381 10.6151
R1817 B.n619 B.n381 10.6151
R1818 B.n620 B.n619 10.6151
R1819 B.n621 B.n620 10.6151
R1820 B.n621 B.n373 10.6151
R1821 B.n631 B.n373 10.6151
R1822 B.n632 B.n631 10.6151
R1823 B.n633 B.n632 10.6151
R1824 B.n633 B.n365 10.6151
R1825 B.n643 B.n365 10.6151
R1826 B.n644 B.n643 10.6151
R1827 B.n645 B.n644 10.6151
R1828 B.n645 B.n357 10.6151
R1829 B.n655 B.n357 10.6151
R1830 B.n656 B.n655 10.6151
R1831 B.n657 B.n656 10.6151
R1832 B.n657 B.n349 10.6151
R1833 B.n667 B.n349 10.6151
R1834 B.n668 B.n667 10.6151
R1835 B.n669 B.n668 10.6151
R1836 B.n669 B.n341 10.6151
R1837 B.n679 B.n341 10.6151
R1838 B.n680 B.n679 10.6151
R1839 B.n681 B.n680 10.6151
R1840 B.n681 B.n333 10.6151
R1841 B.n691 B.n333 10.6151
R1842 B.n692 B.n691 10.6151
R1843 B.n693 B.n692 10.6151
R1844 B.n693 B.n325 10.6151
R1845 B.n703 B.n325 10.6151
R1846 B.n704 B.n703 10.6151
R1847 B.n705 B.n704 10.6151
R1848 B.n705 B.n317 10.6151
R1849 B.n715 B.n317 10.6151
R1850 B.n716 B.n715 10.6151
R1851 B.n717 B.n716 10.6151
R1852 B.n717 B.n309 10.6151
R1853 B.n728 B.n309 10.6151
R1854 B.n729 B.n728 10.6151
R1855 B.n730 B.n729 10.6151
R1856 B.n730 B.n302 10.6151
R1857 B.n741 B.n302 10.6151
R1858 B.n742 B.n741 10.6151
R1859 B.n743 B.n742 10.6151
R1860 B.n743 B.n0 10.6151
R1861 B.n595 B.n594 10.6151
R1862 B.n594 B.n593 10.6151
R1863 B.n593 B.n592 10.6151
R1864 B.n592 B.n590 10.6151
R1865 B.n590 B.n587 10.6151
R1866 B.n587 B.n586 10.6151
R1867 B.n586 B.n583 10.6151
R1868 B.n583 B.n582 10.6151
R1869 B.n582 B.n579 10.6151
R1870 B.n579 B.n578 10.6151
R1871 B.n578 B.n575 10.6151
R1872 B.n575 B.n574 10.6151
R1873 B.n574 B.n571 10.6151
R1874 B.n571 B.n570 10.6151
R1875 B.n570 B.n567 10.6151
R1876 B.n567 B.n566 10.6151
R1877 B.n566 B.n563 10.6151
R1878 B.n563 B.n562 10.6151
R1879 B.n562 B.n559 10.6151
R1880 B.n559 B.n558 10.6151
R1881 B.n558 B.n555 10.6151
R1882 B.n555 B.n554 10.6151
R1883 B.n554 B.n551 10.6151
R1884 B.n551 B.n550 10.6151
R1885 B.n550 B.n547 10.6151
R1886 B.n547 B.n546 10.6151
R1887 B.n546 B.n543 10.6151
R1888 B.n543 B.n542 10.6151
R1889 B.n542 B.n539 10.6151
R1890 B.n539 B.n538 10.6151
R1891 B.n538 B.n535 10.6151
R1892 B.n535 B.n534 10.6151
R1893 B.n534 B.n531 10.6151
R1894 B.n531 B.n530 10.6151
R1895 B.n530 B.n527 10.6151
R1896 B.n525 B.n522 10.6151
R1897 B.n522 B.n521 10.6151
R1898 B.n521 B.n518 10.6151
R1899 B.n518 B.n517 10.6151
R1900 B.n517 B.n514 10.6151
R1901 B.n514 B.n513 10.6151
R1902 B.n513 B.n510 10.6151
R1903 B.n510 B.n509 10.6151
R1904 B.n506 B.n505 10.6151
R1905 B.n505 B.n502 10.6151
R1906 B.n502 B.n501 10.6151
R1907 B.n501 B.n498 10.6151
R1908 B.n498 B.n497 10.6151
R1909 B.n497 B.n494 10.6151
R1910 B.n494 B.n493 10.6151
R1911 B.n493 B.n490 10.6151
R1912 B.n490 B.n489 10.6151
R1913 B.n489 B.n486 10.6151
R1914 B.n486 B.n485 10.6151
R1915 B.n485 B.n482 10.6151
R1916 B.n482 B.n481 10.6151
R1917 B.n481 B.n478 10.6151
R1918 B.n478 B.n477 10.6151
R1919 B.n477 B.n474 10.6151
R1920 B.n474 B.n473 10.6151
R1921 B.n473 B.n470 10.6151
R1922 B.n470 B.n469 10.6151
R1923 B.n469 B.n466 10.6151
R1924 B.n466 B.n465 10.6151
R1925 B.n465 B.n462 10.6151
R1926 B.n462 B.n461 10.6151
R1927 B.n461 B.n458 10.6151
R1928 B.n458 B.n457 10.6151
R1929 B.n457 B.n454 10.6151
R1930 B.n454 B.n453 10.6151
R1931 B.n453 B.n450 10.6151
R1932 B.n450 B.n449 10.6151
R1933 B.n449 B.n446 10.6151
R1934 B.n446 B.n445 10.6151
R1935 B.n445 B.n442 10.6151
R1936 B.n442 B.n441 10.6151
R1937 B.n441 B.n393 10.6151
R1938 B.n601 B.n393 10.6151
R1939 B.n603 B.n602 10.6151
R1940 B.n603 B.n385 10.6151
R1941 B.n613 B.n385 10.6151
R1942 B.n614 B.n613 10.6151
R1943 B.n615 B.n614 10.6151
R1944 B.n615 B.n376 10.6151
R1945 B.n625 B.n376 10.6151
R1946 B.n626 B.n625 10.6151
R1947 B.n627 B.n626 10.6151
R1948 B.n627 B.n369 10.6151
R1949 B.n637 B.n369 10.6151
R1950 B.n638 B.n637 10.6151
R1951 B.n639 B.n638 10.6151
R1952 B.n639 B.n361 10.6151
R1953 B.n649 B.n361 10.6151
R1954 B.n650 B.n649 10.6151
R1955 B.n651 B.n650 10.6151
R1956 B.n651 B.n353 10.6151
R1957 B.n661 B.n353 10.6151
R1958 B.n662 B.n661 10.6151
R1959 B.n663 B.n662 10.6151
R1960 B.n663 B.n345 10.6151
R1961 B.n673 B.n345 10.6151
R1962 B.n674 B.n673 10.6151
R1963 B.n675 B.n674 10.6151
R1964 B.n675 B.n337 10.6151
R1965 B.n685 B.n337 10.6151
R1966 B.n686 B.n685 10.6151
R1967 B.n687 B.n686 10.6151
R1968 B.n687 B.n328 10.6151
R1969 B.n697 B.n328 10.6151
R1970 B.n698 B.n697 10.6151
R1971 B.n699 B.n698 10.6151
R1972 B.n699 B.n321 10.6151
R1973 B.n709 B.n321 10.6151
R1974 B.n710 B.n709 10.6151
R1975 B.n711 B.n710 10.6151
R1976 B.n711 B.n313 10.6151
R1977 B.n721 B.n313 10.6151
R1978 B.n722 B.n721 10.6151
R1979 B.n723 B.n722 10.6151
R1980 B.n723 B.n306 10.6151
R1981 B.n734 B.n306 10.6151
R1982 B.n735 B.n734 10.6151
R1983 B.n737 B.n735 10.6151
R1984 B.n737 B.n736 10.6151
R1985 B.n736 B.n298 10.6151
R1986 B.n748 B.n298 10.6151
R1987 B.n749 B.n748 10.6151
R1988 B.n750 B.n749 10.6151
R1989 B.n751 B.n750 10.6151
R1990 B.n752 B.n751 10.6151
R1991 B.n755 B.n752 10.6151
R1992 B.n756 B.n755 10.6151
R1993 B.n757 B.n756 10.6151
R1994 B.n758 B.n757 10.6151
R1995 B.n760 B.n758 10.6151
R1996 B.n761 B.n760 10.6151
R1997 B.n762 B.n761 10.6151
R1998 B.n763 B.n762 10.6151
R1999 B.n765 B.n763 10.6151
R2000 B.n766 B.n765 10.6151
R2001 B.n767 B.n766 10.6151
R2002 B.n768 B.n767 10.6151
R2003 B.n770 B.n768 10.6151
R2004 B.n771 B.n770 10.6151
R2005 B.n772 B.n771 10.6151
R2006 B.n773 B.n772 10.6151
R2007 B.n775 B.n773 10.6151
R2008 B.n776 B.n775 10.6151
R2009 B.n777 B.n776 10.6151
R2010 B.n778 B.n777 10.6151
R2011 B.n780 B.n778 10.6151
R2012 B.n781 B.n780 10.6151
R2013 B.n782 B.n781 10.6151
R2014 B.n783 B.n782 10.6151
R2015 B.n785 B.n783 10.6151
R2016 B.n786 B.n785 10.6151
R2017 B.n787 B.n786 10.6151
R2018 B.n788 B.n787 10.6151
R2019 B.n790 B.n788 10.6151
R2020 B.n791 B.n790 10.6151
R2021 B.n792 B.n791 10.6151
R2022 B.n793 B.n792 10.6151
R2023 B.n795 B.n793 10.6151
R2024 B.n796 B.n795 10.6151
R2025 B.n797 B.n796 10.6151
R2026 B.n798 B.n797 10.6151
R2027 B.n800 B.n798 10.6151
R2028 B.n801 B.n800 10.6151
R2029 B.n802 B.n801 10.6151
R2030 B.n803 B.n802 10.6151
R2031 B.n805 B.n803 10.6151
R2032 B.n806 B.n805 10.6151
R2033 B.n807 B.n806 10.6151
R2034 B.n808 B.n807 10.6151
R2035 B.n810 B.n808 10.6151
R2036 B.n811 B.n810 10.6151
R2037 B.n812 B.n811 10.6151
R2038 B.n909 B.n1 10.6151
R2039 B.n909 B.n908 10.6151
R2040 B.n908 B.n907 10.6151
R2041 B.n907 B.n10 10.6151
R2042 B.n901 B.n10 10.6151
R2043 B.n901 B.n900 10.6151
R2044 B.n900 B.n899 10.6151
R2045 B.n899 B.n17 10.6151
R2046 B.n893 B.n17 10.6151
R2047 B.n893 B.n892 10.6151
R2048 B.n892 B.n891 10.6151
R2049 B.n891 B.n25 10.6151
R2050 B.n885 B.n25 10.6151
R2051 B.n885 B.n884 10.6151
R2052 B.n884 B.n883 10.6151
R2053 B.n883 B.n32 10.6151
R2054 B.n877 B.n32 10.6151
R2055 B.n877 B.n876 10.6151
R2056 B.n876 B.n875 10.6151
R2057 B.n875 B.n39 10.6151
R2058 B.n869 B.n39 10.6151
R2059 B.n869 B.n868 10.6151
R2060 B.n868 B.n867 10.6151
R2061 B.n867 B.n46 10.6151
R2062 B.n861 B.n46 10.6151
R2063 B.n861 B.n860 10.6151
R2064 B.n860 B.n859 10.6151
R2065 B.n859 B.n53 10.6151
R2066 B.n853 B.n53 10.6151
R2067 B.n853 B.n852 10.6151
R2068 B.n852 B.n851 10.6151
R2069 B.n851 B.n60 10.6151
R2070 B.n845 B.n60 10.6151
R2071 B.n845 B.n844 10.6151
R2072 B.n844 B.n843 10.6151
R2073 B.n843 B.n67 10.6151
R2074 B.n837 B.n67 10.6151
R2075 B.n837 B.n836 10.6151
R2076 B.n836 B.n835 10.6151
R2077 B.n835 B.n74 10.6151
R2078 B.n829 B.n74 10.6151
R2079 B.n829 B.n828 10.6151
R2080 B.n828 B.n827 10.6151
R2081 B.n827 B.n81 10.6151
R2082 B.n821 B.n81 10.6151
R2083 B.n821 B.n820 10.6151
R2084 B.n820 B.n819 10.6151
R2085 B.n819 B.n88 10.6151
R2086 B.n140 B.n139 10.6151
R2087 B.n143 B.n140 10.6151
R2088 B.n144 B.n143 10.6151
R2089 B.n147 B.n144 10.6151
R2090 B.n148 B.n147 10.6151
R2091 B.n151 B.n148 10.6151
R2092 B.n152 B.n151 10.6151
R2093 B.n155 B.n152 10.6151
R2094 B.n156 B.n155 10.6151
R2095 B.n159 B.n156 10.6151
R2096 B.n160 B.n159 10.6151
R2097 B.n163 B.n160 10.6151
R2098 B.n164 B.n163 10.6151
R2099 B.n167 B.n164 10.6151
R2100 B.n168 B.n167 10.6151
R2101 B.n171 B.n168 10.6151
R2102 B.n172 B.n171 10.6151
R2103 B.n175 B.n172 10.6151
R2104 B.n176 B.n175 10.6151
R2105 B.n179 B.n176 10.6151
R2106 B.n180 B.n179 10.6151
R2107 B.n183 B.n180 10.6151
R2108 B.n184 B.n183 10.6151
R2109 B.n187 B.n184 10.6151
R2110 B.n188 B.n187 10.6151
R2111 B.n191 B.n188 10.6151
R2112 B.n192 B.n191 10.6151
R2113 B.n195 B.n192 10.6151
R2114 B.n196 B.n195 10.6151
R2115 B.n199 B.n196 10.6151
R2116 B.n200 B.n199 10.6151
R2117 B.n203 B.n200 10.6151
R2118 B.n204 B.n203 10.6151
R2119 B.n207 B.n204 10.6151
R2120 B.n208 B.n207 10.6151
R2121 B.n212 B.n211 10.6151
R2122 B.n215 B.n212 10.6151
R2123 B.n216 B.n215 10.6151
R2124 B.n219 B.n216 10.6151
R2125 B.n220 B.n219 10.6151
R2126 B.n223 B.n220 10.6151
R2127 B.n224 B.n223 10.6151
R2128 B.n227 B.n224 10.6151
R2129 B.n232 B.n229 10.6151
R2130 B.n233 B.n232 10.6151
R2131 B.n236 B.n233 10.6151
R2132 B.n237 B.n236 10.6151
R2133 B.n240 B.n237 10.6151
R2134 B.n241 B.n240 10.6151
R2135 B.n244 B.n241 10.6151
R2136 B.n245 B.n244 10.6151
R2137 B.n248 B.n245 10.6151
R2138 B.n249 B.n248 10.6151
R2139 B.n252 B.n249 10.6151
R2140 B.n253 B.n252 10.6151
R2141 B.n256 B.n253 10.6151
R2142 B.n257 B.n256 10.6151
R2143 B.n260 B.n257 10.6151
R2144 B.n261 B.n260 10.6151
R2145 B.n264 B.n261 10.6151
R2146 B.n265 B.n264 10.6151
R2147 B.n268 B.n265 10.6151
R2148 B.n269 B.n268 10.6151
R2149 B.n272 B.n269 10.6151
R2150 B.n273 B.n272 10.6151
R2151 B.n276 B.n273 10.6151
R2152 B.n277 B.n276 10.6151
R2153 B.n280 B.n277 10.6151
R2154 B.n281 B.n280 10.6151
R2155 B.n284 B.n281 10.6151
R2156 B.n285 B.n284 10.6151
R2157 B.n288 B.n285 10.6151
R2158 B.n289 B.n288 10.6151
R2159 B.n292 B.n289 10.6151
R2160 B.n293 B.n292 10.6151
R2161 B.n296 B.n293 10.6151
R2162 B.n297 B.n296 10.6151
R2163 B.n813 B.n297 10.6151
R2164 B.n917 B.n0 8.11757
R2165 B.n917 B.n1 8.11757
R2166 B.n526 B.n525 6.5566
R2167 B.n509 B.n439 6.5566
R2168 B.n211 B.n137 6.5566
R2169 B.n228 B.n227 6.5566
R2170 B.t4 B.n347 6.49018
R2171 B.t3 B.n51 6.49018
R2172 B.n527 B.n526 4.05904
R2173 B.n506 B.n439 4.05904
R2174 B.n208 B.n137 4.05904
R2175 B.n229 B.n228 4.05904
R2176 VN.n34 VN.n33 161.3
R2177 VN.n32 VN.n19 161.3
R2178 VN.n31 VN.n30 161.3
R2179 VN.n29 VN.n20 161.3
R2180 VN.n28 VN.n27 161.3
R2181 VN.n26 VN.n21 161.3
R2182 VN.n25 VN.n24 161.3
R2183 VN.n16 VN.n15 161.3
R2184 VN.n14 VN.n1 161.3
R2185 VN.n13 VN.n12 161.3
R2186 VN.n11 VN.n2 161.3
R2187 VN.n10 VN.n9 161.3
R2188 VN.n8 VN.n3 161.3
R2189 VN.n7 VN.n6 161.3
R2190 VN.n23 VN.t3 107.742
R2191 VN.n5 VN.t5 107.742
R2192 VN.n17 VN.n0 75.7718
R2193 VN.n35 VN.n18 75.7718
R2194 VN.n4 VN.t2 74.9282
R2195 VN.n0 VN.t1 74.9282
R2196 VN.n22 VN.t4 74.9282
R2197 VN.n18 VN.t0 74.9282
R2198 VN.n5 VN.n4 61.8768
R2199 VN.n23 VN.n22 61.8768
R2200 VN VN.n35 49.7858
R2201 VN.n13 VN.n2 42.3581
R2202 VN.n31 VN.n20 42.3581
R2203 VN.n9 VN.n2 38.4631
R2204 VN.n27 VN.n20 38.4631
R2205 VN.n8 VN.n7 24.3439
R2206 VN.n9 VN.n8 24.3439
R2207 VN.n14 VN.n13 24.3439
R2208 VN.n15 VN.n14 24.3439
R2209 VN.n27 VN.n26 24.3439
R2210 VN.n26 VN.n25 24.3439
R2211 VN.n33 VN.n32 24.3439
R2212 VN.n32 VN.n31 24.3439
R2213 VN.n15 VN.n0 14.1197
R2214 VN.n33 VN.n18 14.1197
R2215 VN.n7 VN.n4 12.1722
R2216 VN.n25 VN.n22 12.1722
R2217 VN.n6 VN.n5 4.197
R2218 VN.n24 VN.n23 4.197
R2219 VN.n35 VN.n34 0.355081
R2220 VN.n17 VN.n16 0.355081
R2221 VN VN.n17 0.26685
R2222 VN.n34 VN.n19 0.189894
R2223 VN.n30 VN.n19 0.189894
R2224 VN.n30 VN.n29 0.189894
R2225 VN.n29 VN.n28 0.189894
R2226 VN.n28 VN.n21 0.189894
R2227 VN.n24 VN.n21 0.189894
R2228 VN.n6 VN.n3 0.189894
R2229 VN.n10 VN.n3 0.189894
R2230 VN.n11 VN.n10 0.189894
R2231 VN.n12 VN.n11 0.189894
R2232 VN.n12 VN.n1 0.189894
R2233 VN.n16 VN.n1 0.189894
R2234 VDD2.n103 VDD2.n55 289.615
R2235 VDD2.n48 VDD2.n0 289.615
R2236 VDD2.n104 VDD2.n103 185
R2237 VDD2.n102 VDD2.n101 185
R2238 VDD2.n59 VDD2.n58 185
R2239 VDD2.n96 VDD2.n95 185
R2240 VDD2.n94 VDD2.n61 185
R2241 VDD2.n93 VDD2.n92 185
R2242 VDD2.n64 VDD2.n62 185
R2243 VDD2.n87 VDD2.n86 185
R2244 VDD2.n85 VDD2.n84 185
R2245 VDD2.n68 VDD2.n67 185
R2246 VDD2.n79 VDD2.n78 185
R2247 VDD2.n77 VDD2.n76 185
R2248 VDD2.n72 VDD2.n71 185
R2249 VDD2.n16 VDD2.n15 185
R2250 VDD2.n21 VDD2.n20 185
R2251 VDD2.n23 VDD2.n22 185
R2252 VDD2.n12 VDD2.n11 185
R2253 VDD2.n29 VDD2.n28 185
R2254 VDD2.n31 VDD2.n30 185
R2255 VDD2.n8 VDD2.n7 185
R2256 VDD2.n38 VDD2.n37 185
R2257 VDD2.n39 VDD2.n6 185
R2258 VDD2.n41 VDD2.n40 185
R2259 VDD2.n4 VDD2.n3 185
R2260 VDD2.n47 VDD2.n46 185
R2261 VDD2.n49 VDD2.n48 185
R2262 VDD2.n73 VDD2.t5 149.524
R2263 VDD2.n17 VDD2.t0 149.524
R2264 VDD2.n103 VDD2.n102 104.615
R2265 VDD2.n102 VDD2.n58 104.615
R2266 VDD2.n95 VDD2.n58 104.615
R2267 VDD2.n95 VDD2.n94 104.615
R2268 VDD2.n94 VDD2.n93 104.615
R2269 VDD2.n93 VDD2.n62 104.615
R2270 VDD2.n86 VDD2.n62 104.615
R2271 VDD2.n86 VDD2.n85 104.615
R2272 VDD2.n85 VDD2.n67 104.615
R2273 VDD2.n78 VDD2.n67 104.615
R2274 VDD2.n78 VDD2.n77 104.615
R2275 VDD2.n77 VDD2.n71 104.615
R2276 VDD2.n21 VDD2.n15 104.615
R2277 VDD2.n22 VDD2.n21 104.615
R2278 VDD2.n22 VDD2.n11 104.615
R2279 VDD2.n29 VDD2.n11 104.615
R2280 VDD2.n30 VDD2.n29 104.615
R2281 VDD2.n30 VDD2.n7 104.615
R2282 VDD2.n38 VDD2.n7 104.615
R2283 VDD2.n39 VDD2.n38 104.615
R2284 VDD2.n40 VDD2.n39 104.615
R2285 VDD2.n40 VDD2.n3 104.615
R2286 VDD2.n47 VDD2.n3 104.615
R2287 VDD2.n48 VDD2.n47 104.615
R2288 VDD2.n54 VDD2.n53 63.7356
R2289 VDD2 VDD2.n109 63.7328
R2290 VDD2.t5 VDD2.n71 52.3082
R2291 VDD2.t0 VDD2.n15 52.3082
R2292 VDD2.n54 VDD2.n52 51.4855
R2293 VDD2.n108 VDD2.n107 49.252
R2294 VDD2.n108 VDD2.n54 42.2369
R2295 VDD2.n96 VDD2.n61 13.1884
R2296 VDD2.n41 VDD2.n6 13.1884
R2297 VDD2.n97 VDD2.n59 12.8005
R2298 VDD2.n92 VDD2.n63 12.8005
R2299 VDD2.n37 VDD2.n36 12.8005
R2300 VDD2.n42 VDD2.n4 12.8005
R2301 VDD2.n101 VDD2.n100 12.0247
R2302 VDD2.n91 VDD2.n64 12.0247
R2303 VDD2.n35 VDD2.n8 12.0247
R2304 VDD2.n46 VDD2.n45 12.0247
R2305 VDD2.n104 VDD2.n57 11.249
R2306 VDD2.n88 VDD2.n87 11.249
R2307 VDD2.n32 VDD2.n31 11.249
R2308 VDD2.n49 VDD2.n2 11.249
R2309 VDD2.n105 VDD2.n55 10.4732
R2310 VDD2.n84 VDD2.n66 10.4732
R2311 VDD2.n28 VDD2.n10 10.4732
R2312 VDD2.n50 VDD2.n0 10.4732
R2313 VDD2.n73 VDD2.n72 10.2747
R2314 VDD2.n17 VDD2.n16 10.2747
R2315 VDD2.n83 VDD2.n68 9.69747
R2316 VDD2.n27 VDD2.n12 9.69747
R2317 VDD2.n107 VDD2.n106 9.45567
R2318 VDD2.n52 VDD2.n51 9.45567
R2319 VDD2.n75 VDD2.n74 9.3005
R2320 VDD2.n70 VDD2.n69 9.3005
R2321 VDD2.n81 VDD2.n80 9.3005
R2322 VDD2.n83 VDD2.n82 9.3005
R2323 VDD2.n66 VDD2.n65 9.3005
R2324 VDD2.n89 VDD2.n88 9.3005
R2325 VDD2.n91 VDD2.n90 9.3005
R2326 VDD2.n63 VDD2.n60 9.3005
R2327 VDD2.n106 VDD2.n105 9.3005
R2328 VDD2.n57 VDD2.n56 9.3005
R2329 VDD2.n100 VDD2.n99 9.3005
R2330 VDD2.n98 VDD2.n97 9.3005
R2331 VDD2.n51 VDD2.n50 9.3005
R2332 VDD2.n2 VDD2.n1 9.3005
R2333 VDD2.n45 VDD2.n44 9.3005
R2334 VDD2.n43 VDD2.n42 9.3005
R2335 VDD2.n19 VDD2.n18 9.3005
R2336 VDD2.n14 VDD2.n13 9.3005
R2337 VDD2.n25 VDD2.n24 9.3005
R2338 VDD2.n27 VDD2.n26 9.3005
R2339 VDD2.n10 VDD2.n9 9.3005
R2340 VDD2.n33 VDD2.n32 9.3005
R2341 VDD2.n35 VDD2.n34 9.3005
R2342 VDD2.n36 VDD2.n5 9.3005
R2343 VDD2.n80 VDD2.n79 8.92171
R2344 VDD2.n24 VDD2.n23 8.92171
R2345 VDD2.n76 VDD2.n70 8.14595
R2346 VDD2.n20 VDD2.n14 8.14595
R2347 VDD2.n75 VDD2.n72 7.3702
R2348 VDD2.n19 VDD2.n16 7.3702
R2349 VDD2.n76 VDD2.n75 5.81868
R2350 VDD2.n20 VDD2.n19 5.81868
R2351 VDD2.n79 VDD2.n70 5.04292
R2352 VDD2.n23 VDD2.n14 5.04292
R2353 VDD2.n80 VDD2.n68 4.26717
R2354 VDD2.n24 VDD2.n12 4.26717
R2355 VDD2.n107 VDD2.n55 3.49141
R2356 VDD2.n84 VDD2.n83 3.49141
R2357 VDD2.n28 VDD2.n27 3.49141
R2358 VDD2.n52 VDD2.n0 3.49141
R2359 VDD2.n74 VDD2.n73 2.84303
R2360 VDD2.n18 VDD2.n17 2.84303
R2361 VDD2.n105 VDD2.n104 2.71565
R2362 VDD2.n87 VDD2.n66 2.71565
R2363 VDD2.n31 VDD2.n10 2.71565
R2364 VDD2.n50 VDD2.n49 2.71565
R2365 VDD2 VDD2.n108 2.34748
R2366 VDD2.n109 VDD2.t1 1.98447
R2367 VDD2.n109 VDD2.t2 1.98447
R2368 VDD2.n53 VDD2.t3 1.98447
R2369 VDD2.n53 VDD2.t4 1.98447
R2370 VDD2.n101 VDD2.n57 1.93989
R2371 VDD2.n88 VDD2.n64 1.93989
R2372 VDD2.n32 VDD2.n8 1.93989
R2373 VDD2.n46 VDD2.n2 1.93989
R2374 VDD2.n100 VDD2.n59 1.16414
R2375 VDD2.n92 VDD2.n91 1.16414
R2376 VDD2.n37 VDD2.n35 1.16414
R2377 VDD2.n45 VDD2.n4 1.16414
R2378 VDD2.n97 VDD2.n96 0.388379
R2379 VDD2.n63 VDD2.n61 0.388379
R2380 VDD2.n36 VDD2.n6 0.388379
R2381 VDD2.n42 VDD2.n41 0.388379
R2382 VDD2.n106 VDD2.n56 0.155672
R2383 VDD2.n99 VDD2.n56 0.155672
R2384 VDD2.n99 VDD2.n98 0.155672
R2385 VDD2.n98 VDD2.n60 0.155672
R2386 VDD2.n90 VDD2.n60 0.155672
R2387 VDD2.n90 VDD2.n89 0.155672
R2388 VDD2.n89 VDD2.n65 0.155672
R2389 VDD2.n82 VDD2.n65 0.155672
R2390 VDD2.n82 VDD2.n81 0.155672
R2391 VDD2.n81 VDD2.n69 0.155672
R2392 VDD2.n74 VDD2.n69 0.155672
R2393 VDD2.n18 VDD2.n13 0.155672
R2394 VDD2.n25 VDD2.n13 0.155672
R2395 VDD2.n26 VDD2.n25 0.155672
R2396 VDD2.n26 VDD2.n9 0.155672
R2397 VDD2.n33 VDD2.n9 0.155672
R2398 VDD2.n34 VDD2.n33 0.155672
R2399 VDD2.n34 VDD2.n5 0.155672
R2400 VDD2.n43 VDD2.n5 0.155672
R2401 VDD2.n44 VDD2.n43 0.155672
R2402 VDD2.n44 VDD2.n1 0.155672
R2403 VDD2.n51 VDD2.n1 0.155672
C0 VN VTAIL 6.26878f
C1 VTAIL VDD2 7.27898f
C2 VP VDD1 6.22514f
C3 VN VDD1 0.151064f
C4 VDD1 VDD2 1.64349f
C5 VTAIL VDD1 7.22312f
C6 VP VN 7.15396f
C7 VP VDD2 0.509396f
C8 VN VDD2 5.8696f
C9 VP VTAIL 6.283f
C10 VDD2 B 6.092057f
C11 VDD1 B 6.246597f
C12 VTAIL B 7.39017f
C13 VN B 14.54401f
C14 VP B 13.241833f
C15 VDD2.n0 B 0.028854f
C16 VDD2.n1 B 0.021564f
C17 VDD2.n2 B 0.011587f
C18 VDD2.n3 B 0.027388f
C19 VDD2.n4 B 0.012269f
C20 VDD2.n5 B 0.021564f
C21 VDD2.n6 B 0.011928f
C22 VDD2.n7 B 0.027388f
C23 VDD2.n8 B 0.012269f
C24 VDD2.n9 B 0.021564f
C25 VDD2.n10 B 0.011587f
C26 VDD2.n11 B 0.027388f
C27 VDD2.n12 B 0.012269f
C28 VDD2.n13 B 0.021564f
C29 VDD2.n14 B 0.011587f
C30 VDD2.n15 B 0.020541f
C31 VDD2.n16 B 0.019361f
C32 VDD2.t0 B 0.046024f
C33 VDD2.n17 B 0.13875f
C34 VDD2.n18 B 0.894094f
C35 VDD2.n19 B 0.011587f
C36 VDD2.n20 B 0.012269f
C37 VDD2.n21 B 0.027388f
C38 VDD2.n22 B 0.027388f
C39 VDD2.n23 B 0.012269f
C40 VDD2.n24 B 0.011587f
C41 VDD2.n25 B 0.021564f
C42 VDD2.n26 B 0.021564f
C43 VDD2.n27 B 0.011587f
C44 VDD2.n28 B 0.012269f
C45 VDD2.n29 B 0.027388f
C46 VDD2.n30 B 0.027388f
C47 VDD2.n31 B 0.012269f
C48 VDD2.n32 B 0.011587f
C49 VDD2.n33 B 0.021564f
C50 VDD2.n34 B 0.021564f
C51 VDD2.n35 B 0.011587f
C52 VDD2.n36 B 0.011587f
C53 VDD2.n37 B 0.012269f
C54 VDD2.n38 B 0.027388f
C55 VDD2.n39 B 0.027388f
C56 VDD2.n40 B 0.027388f
C57 VDD2.n41 B 0.011928f
C58 VDD2.n42 B 0.011587f
C59 VDD2.n43 B 0.021564f
C60 VDD2.n44 B 0.021564f
C61 VDD2.n45 B 0.011587f
C62 VDD2.n46 B 0.012269f
C63 VDD2.n47 B 0.027388f
C64 VDD2.n48 B 0.056718f
C65 VDD2.n49 B 0.012269f
C66 VDD2.n50 B 0.011587f
C67 VDD2.n51 B 0.050432f
C68 VDD2.n52 B 0.054931f
C69 VDD2.t3 B 0.17006f
C70 VDD2.t4 B 0.17006f
C71 VDD2.n53 B 1.50241f
C72 VDD2.n54 B 2.42807f
C73 VDD2.n55 B 0.028854f
C74 VDD2.n56 B 0.021564f
C75 VDD2.n57 B 0.011587f
C76 VDD2.n58 B 0.027388f
C77 VDD2.n59 B 0.012269f
C78 VDD2.n60 B 0.021564f
C79 VDD2.n61 B 0.011928f
C80 VDD2.n62 B 0.027388f
C81 VDD2.n63 B 0.011587f
C82 VDD2.n64 B 0.012269f
C83 VDD2.n65 B 0.021564f
C84 VDD2.n66 B 0.011587f
C85 VDD2.n67 B 0.027388f
C86 VDD2.n68 B 0.012269f
C87 VDD2.n69 B 0.021564f
C88 VDD2.n70 B 0.011587f
C89 VDD2.n71 B 0.020541f
C90 VDD2.n72 B 0.019361f
C91 VDD2.t5 B 0.046024f
C92 VDD2.n73 B 0.13875f
C93 VDD2.n74 B 0.894094f
C94 VDD2.n75 B 0.011587f
C95 VDD2.n76 B 0.012269f
C96 VDD2.n77 B 0.027388f
C97 VDD2.n78 B 0.027388f
C98 VDD2.n79 B 0.012269f
C99 VDD2.n80 B 0.011587f
C100 VDD2.n81 B 0.021564f
C101 VDD2.n82 B 0.021564f
C102 VDD2.n83 B 0.011587f
C103 VDD2.n84 B 0.012269f
C104 VDD2.n85 B 0.027388f
C105 VDD2.n86 B 0.027388f
C106 VDD2.n87 B 0.012269f
C107 VDD2.n88 B 0.011587f
C108 VDD2.n89 B 0.021564f
C109 VDD2.n90 B 0.021564f
C110 VDD2.n91 B 0.011587f
C111 VDD2.n92 B 0.012269f
C112 VDD2.n93 B 0.027388f
C113 VDD2.n94 B 0.027388f
C114 VDD2.n95 B 0.027388f
C115 VDD2.n96 B 0.011928f
C116 VDD2.n97 B 0.011587f
C117 VDD2.n98 B 0.021564f
C118 VDD2.n99 B 0.021564f
C119 VDD2.n100 B 0.011587f
C120 VDD2.n101 B 0.012269f
C121 VDD2.n102 B 0.027388f
C122 VDD2.n103 B 0.056718f
C123 VDD2.n104 B 0.012269f
C124 VDD2.n105 B 0.011587f
C125 VDD2.n106 B 0.050432f
C126 VDD2.n107 B 0.046374f
C127 VDD2.n108 B 2.21868f
C128 VDD2.t1 B 0.17006f
C129 VDD2.t2 B 0.17006f
C130 VDD2.n109 B 1.50238f
C131 VN.t1 B 1.82868f
C132 VN.n0 B 0.73087f
C133 VN.n1 B 0.021072f
C134 VN.n2 B 0.017162f
C135 VN.n3 B 0.021072f
C136 VN.t2 B 1.82868f
C137 VN.n4 B 0.720001f
C138 VN.t5 B 2.07202f
C139 VN.n5 B 0.686468f
C140 VN.n6 B 0.245605f
C141 VN.n7 B 0.029726f
C142 VN.n8 B 0.039471f
C143 VN.n9 B 0.042475f
C144 VN.n10 B 0.021072f
C145 VN.n11 B 0.021072f
C146 VN.n12 B 0.021072f
C147 VN.n13 B 0.041625f
C148 VN.n14 B 0.039471f
C149 VN.n15 B 0.031285f
C150 VN.n16 B 0.034016f
C151 VN.n17 B 0.050658f
C152 VN.t0 B 1.82868f
C153 VN.n18 B 0.73087f
C154 VN.n19 B 0.021072f
C155 VN.n20 B 0.017162f
C156 VN.n21 B 0.021072f
C157 VN.t4 B 1.82868f
C158 VN.n22 B 0.720001f
C159 VN.t3 B 2.07202f
C160 VN.n23 B 0.686468f
C161 VN.n24 B 0.245605f
C162 VN.n25 B 0.029726f
C163 VN.n26 B 0.039471f
C164 VN.n27 B 0.042475f
C165 VN.n28 B 0.021072f
C166 VN.n29 B 0.021072f
C167 VN.n30 B 0.021072f
C168 VN.n31 B 0.041625f
C169 VN.n32 B 0.039471f
C170 VN.n33 B 0.031285f
C171 VN.n34 B 0.034016f
C172 VN.n35 B 1.19332f
C173 VDD1.n0 B 0.029116f
C174 VDD1.n1 B 0.021759f
C175 VDD1.n2 B 0.011692f
C176 VDD1.n3 B 0.027636f
C177 VDD1.n4 B 0.01238f
C178 VDD1.n5 B 0.021759f
C179 VDD1.n6 B 0.012036f
C180 VDD1.n7 B 0.027636f
C181 VDD1.n8 B 0.011692f
C182 VDD1.n9 B 0.01238f
C183 VDD1.n10 B 0.021759f
C184 VDD1.n11 B 0.011692f
C185 VDD1.n12 B 0.027636f
C186 VDD1.n13 B 0.01238f
C187 VDD1.n14 B 0.021759f
C188 VDD1.n15 B 0.011692f
C189 VDD1.n16 B 0.020727f
C190 VDD1.n17 B 0.019537f
C191 VDD1.t5 B 0.046441f
C192 VDD1.n18 B 0.140007f
C193 VDD1.n19 B 0.902197f
C194 VDD1.n20 B 0.011692f
C195 VDD1.n21 B 0.01238f
C196 VDD1.n22 B 0.027636f
C197 VDD1.n23 B 0.027636f
C198 VDD1.n24 B 0.01238f
C199 VDD1.n25 B 0.011692f
C200 VDD1.n26 B 0.021759f
C201 VDD1.n27 B 0.021759f
C202 VDD1.n28 B 0.011692f
C203 VDD1.n29 B 0.01238f
C204 VDD1.n30 B 0.027636f
C205 VDD1.n31 B 0.027636f
C206 VDD1.n32 B 0.01238f
C207 VDD1.n33 B 0.011692f
C208 VDD1.n34 B 0.021759f
C209 VDD1.n35 B 0.021759f
C210 VDD1.n36 B 0.011692f
C211 VDD1.n37 B 0.01238f
C212 VDD1.n38 B 0.027636f
C213 VDD1.n39 B 0.027636f
C214 VDD1.n40 B 0.027636f
C215 VDD1.n41 B 0.012036f
C216 VDD1.n42 B 0.011692f
C217 VDD1.n43 B 0.021759f
C218 VDD1.n44 B 0.021759f
C219 VDD1.n45 B 0.011692f
C220 VDD1.n46 B 0.01238f
C221 VDD1.n47 B 0.027636f
C222 VDD1.n48 B 0.057232f
C223 VDD1.n49 B 0.01238f
C224 VDD1.n50 B 0.011692f
C225 VDD1.n51 B 0.050889f
C226 VDD1.n52 B 0.0562f
C227 VDD1.n53 B 0.029116f
C228 VDD1.n54 B 0.021759f
C229 VDD1.n55 B 0.011692f
C230 VDD1.n56 B 0.027636f
C231 VDD1.n57 B 0.01238f
C232 VDD1.n58 B 0.021759f
C233 VDD1.n59 B 0.012036f
C234 VDD1.n60 B 0.027636f
C235 VDD1.n61 B 0.01238f
C236 VDD1.n62 B 0.021759f
C237 VDD1.n63 B 0.011692f
C238 VDD1.n64 B 0.027636f
C239 VDD1.n65 B 0.01238f
C240 VDD1.n66 B 0.021759f
C241 VDD1.n67 B 0.011692f
C242 VDD1.n68 B 0.020727f
C243 VDD1.n69 B 0.019537f
C244 VDD1.t4 B 0.046441f
C245 VDD1.n70 B 0.140007f
C246 VDD1.n71 B 0.902197f
C247 VDD1.n72 B 0.011692f
C248 VDD1.n73 B 0.01238f
C249 VDD1.n74 B 0.027636f
C250 VDD1.n75 B 0.027636f
C251 VDD1.n76 B 0.01238f
C252 VDD1.n77 B 0.011692f
C253 VDD1.n78 B 0.021759f
C254 VDD1.n79 B 0.021759f
C255 VDD1.n80 B 0.011692f
C256 VDD1.n81 B 0.01238f
C257 VDD1.n82 B 0.027636f
C258 VDD1.n83 B 0.027636f
C259 VDD1.n84 B 0.01238f
C260 VDD1.n85 B 0.011692f
C261 VDD1.n86 B 0.021759f
C262 VDD1.n87 B 0.021759f
C263 VDD1.n88 B 0.011692f
C264 VDD1.n89 B 0.011692f
C265 VDD1.n90 B 0.01238f
C266 VDD1.n91 B 0.027636f
C267 VDD1.n92 B 0.027636f
C268 VDD1.n93 B 0.027636f
C269 VDD1.n94 B 0.012036f
C270 VDD1.n95 B 0.011692f
C271 VDD1.n96 B 0.021759f
C272 VDD1.n97 B 0.021759f
C273 VDD1.n98 B 0.011692f
C274 VDD1.n99 B 0.01238f
C275 VDD1.n100 B 0.027636f
C276 VDD1.n101 B 0.057232f
C277 VDD1.n102 B 0.01238f
C278 VDD1.n103 B 0.011692f
C279 VDD1.n104 B 0.050889f
C280 VDD1.n105 B 0.055429f
C281 VDD1.t1 B 0.171601f
C282 VDD1.t0 B 0.171601f
C283 VDD1.n106 B 1.51603f
C284 VDD1.n107 B 2.57051f
C285 VDD1.t3 B 0.171601f
C286 VDD1.t2 B 0.171601f
C287 VDD1.n108 B 1.51103f
C288 VDD1.n109 B 2.44122f
C289 VTAIL.t2 B 0.196518f
C290 VTAIL.t1 B 0.196518f
C291 VTAIL.n0 B 1.65914f
C292 VTAIL.n1 B 0.466465f
C293 VTAIL.n2 B 0.033344f
C294 VTAIL.n3 B 0.024918f
C295 VTAIL.n4 B 0.01339f
C296 VTAIL.n5 B 0.031649f
C297 VTAIL.n6 B 0.014178f
C298 VTAIL.n7 B 0.024918f
C299 VTAIL.n8 B 0.013784f
C300 VTAIL.n9 B 0.031649f
C301 VTAIL.n10 B 0.014178f
C302 VTAIL.n11 B 0.024918f
C303 VTAIL.n12 B 0.01339f
C304 VTAIL.n13 B 0.031649f
C305 VTAIL.n14 B 0.014178f
C306 VTAIL.n15 B 0.024918f
C307 VTAIL.n16 B 0.01339f
C308 VTAIL.n17 B 0.023737f
C309 VTAIL.n18 B 0.022373f
C310 VTAIL.t6 B 0.053184f
C311 VTAIL.n19 B 0.160337f
C312 VTAIL.n20 B 1.0332f
C313 VTAIL.n21 B 0.01339f
C314 VTAIL.n22 B 0.014178f
C315 VTAIL.n23 B 0.031649f
C316 VTAIL.n24 B 0.031649f
C317 VTAIL.n25 B 0.014178f
C318 VTAIL.n26 B 0.01339f
C319 VTAIL.n27 B 0.024918f
C320 VTAIL.n28 B 0.024918f
C321 VTAIL.n29 B 0.01339f
C322 VTAIL.n30 B 0.014178f
C323 VTAIL.n31 B 0.031649f
C324 VTAIL.n32 B 0.031649f
C325 VTAIL.n33 B 0.014178f
C326 VTAIL.n34 B 0.01339f
C327 VTAIL.n35 B 0.024918f
C328 VTAIL.n36 B 0.024918f
C329 VTAIL.n37 B 0.01339f
C330 VTAIL.n38 B 0.01339f
C331 VTAIL.n39 B 0.014178f
C332 VTAIL.n40 B 0.031649f
C333 VTAIL.n41 B 0.031649f
C334 VTAIL.n42 B 0.031649f
C335 VTAIL.n43 B 0.013784f
C336 VTAIL.n44 B 0.01339f
C337 VTAIL.n45 B 0.024918f
C338 VTAIL.n46 B 0.024918f
C339 VTAIL.n47 B 0.01339f
C340 VTAIL.n48 B 0.014178f
C341 VTAIL.n49 B 0.031649f
C342 VTAIL.n50 B 0.065542f
C343 VTAIL.n51 B 0.014178f
C344 VTAIL.n52 B 0.01339f
C345 VTAIL.n53 B 0.058278f
C346 VTAIL.n54 B 0.036389f
C347 VTAIL.n55 B 0.426936f
C348 VTAIL.t9 B 0.196518f
C349 VTAIL.t10 B 0.196518f
C350 VTAIL.n56 B 1.65914f
C351 VTAIL.n57 B 2.00467f
C352 VTAIL.t4 B 0.196518f
C353 VTAIL.t0 B 0.196518f
C354 VTAIL.n58 B 1.65915f
C355 VTAIL.n59 B 2.00466f
C356 VTAIL.n60 B 0.033344f
C357 VTAIL.n61 B 0.024918f
C358 VTAIL.n62 B 0.01339f
C359 VTAIL.n63 B 0.031649f
C360 VTAIL.n64 B 0.014178f
C361 VTAIL.n65 B 0.024918f
C362 VTAIL.n66 B 0.013784f
C363 VTAIL.n67 B 0.031649f
C364 VTAIL.n68 B 0.01339f
C365 VTAIL.n69 B 0.014178f
C366 VTAIL.n70 B 0.024918f
C367 VTAIL.n71 B 0.01339f
C368 VTAIL.n72 B 0.031649f
C369 VTAIL.n73 B 0.014178f
C370 VTAIL.n74 B 0.024918f
C371 VTAIL.n75 B 0.01339f
C372 VTAIL.n76 B 0.023737f
C373 VTAIL.n77 B 0.022373f
C374 VTAIL.t5 B 0.053184f
C375 VTAIL.n78 B 0.160337f
C376 VTAIL.n79 B 1.0332f
C377 VTAIL.n80 B 0.01339f
C378 VTAIL.n81 B 0.014178f
C379 VTAIL.n82 B 0.031649f
C380 VTAIL.n83 B 0.031649f
C381 VTAIL.n84 B 0.014178f
C382 VTAIL.n85 B 0.01339f
C383 VTAIL.n86 B 0.024918f
C384 VTAIL.n87 B 0.024918f
C385 VTAIL.n88 B 0.01339f
C386 VTAIL.n89 B 0.014178f
C387 VTAIL.n90 B 0.031649f
C388 VTAIL.n91 B 0.031649f
C389 VTAIL.n92 B 0.014178f
C390 VTAIL.n93 B 0.01339f
C391 VTAIL.n94 B 0.024918f
C392 VTAIL.n95 B 0.024918f
C393 VTAIL.n96 B 0.01339f
C394 VTAIL.n97 B 0.014178f
C395 VTAIL.n98 B 0.031649f
C396 VTAIL.n99 B 0.031649f
C397 VTAIL.n100 B 0.031649f
C398 VTAIL.n101 B 0.013784f
C399 VTAIL.n102 B 0.01339f
C400 VTAIL.n103 B 0.024918f
C401 VTAIL.n104 B 0.024918f
C402 VTAIL.n105 B 0.01339f
C403 VTAIL.n106 B 0.014178f
C404 VTAIL.n107 B 0.031649f
C405 VTAIL.n108 B 0.065542f
C406 VTAIL.n109 B 0.014178f
C407 VTAIL.n110 B 0.01339f
C408 VTAIL.n111 B 0.058278f
C409 VTAIL.n112 B 0.036389f
C410 VTAIL.n113 B 0.426936f
C411 VTAIL.t7 B 0.196518f
C412 VTAIL.t8 B 0.196518f
C413 VTAIL.n114 B 1.65915f
C414 VTAIL.n115 B 0.645556f
C415 VTAIL.n116 B 0.033344f
C416 VTAIL.n117 B 0.024918f
C417 VTAIL.n118 B 0.01339f
C418 VTAIL.n119 B 0.031649f
C419 VTAIL.n120 B 0.014178f
C420 VTAIL.n121 B 0.024918f
C421 VTAIL.n122 B 0.013784f
C422 VTAIL.n123 B 0.031649f
C423 VTAIL.n124 B 0.01339f
C424 VTAIL.n125 B 0.014178f
C425 VTAIL.n126 B 0.024918f
C426 VTAIL.n127 B 0.01339f
C427 VTAIL.n128 B 0.031649f
C428 VTAIL.n129 B 0.014178f
C429 VTAIL.n130 B 0.024918f
C430 VTAIL.n131 B 0.01339f
C431 VTAIL.n132 B 0.023737f
C432 VTAIL.n133 B 0.022373f
C433 VTAIL.t11 B 0.053184f
C434 VTAIL.n134 B 0.160337f
C435 VTAIL.n135 B 1.0332f
C436 VTAIL.n136 B 0.01339f
C437 VTAIL.n137 B 0.014178f
C438 VTAIL.n138 B 0.031649f
C439 VTAIL.n139 B 0.031649f
C440 VTAIL.n140 B 0.014178f
C441 VTAIL.n141 B 0.01339f
C442 VTAIL.n142 B 0.024918f
C443 VTAIL.n143 B 0.024918f
C444 VTAIL.n144 B 0.01339f
C445 VTAIL.n145 B 0.014178f
C446 VTAIL.n146 B 0.031649f
C447 VTAIL.n147 B 0.031649f
C448 VTAIL.n148 B 0.014178f
C449 VTAIL.n149 B 0.01339f
C450 VTAIL.n150 B 0.024918f
C451 VTAIL.n151 B 0.024918f
C452 VTAIL.n152 B 0.01339f
C453 VTAIL.n153 B 0.014178f
C454 VTAIL.n154 B 0.031649f
C455 VTAIL.n155 B 0.031649f
C456 VTAIL.n156 B 0.031649f
C457 VTAIL.n157 B 0.013784f
C458 VTAIL.n158 B 0.01339f
C459 VTAIL.n159 B 0.024918f
C460 VTAIL.n160 B 0.024918f
C461 VTAIL.n161 B 0.01339f
C462 VTAIL.n162 B 0.014178f
C463 VTAIL.n163 B 0.031649f
C464 VTAIL.n164 B 0.065542f
C465 VTAIL.n165 B 0.014178f
C466 VTAIL.n166 B 0.01339f
C467 VTAIL.n167 B 0.058278f
C468 VTAIL.n168 B 0.036389f
C469 VTAIL.n169 B 1.54101f
C470 VTAIL.n170 B 0.033344f
C471 VTAIL.n171 B 0.024918f
C472 VTAIL.n172 B 0.01339f
C473 VTAIL.n173 B 0.031649f
C474 VTAIL.n174 B 0.014178f
C475 VTAIL.n175 B 0.024918f
C476 VTAIL.n176 B 0.013784f
C477 VTAIL.n177 B 0.031649f
C478 VTAIL.n178 B 0.014178f
C479 VTAIL.n179 B 0.024918f
C480 VTAIL.n180 B 0.01339f
C481 VTAIL.n181 B 0.031649f
C482 VTAIL.n182 B 0.014178f
C483 VTAIL.n183 B 0.024918f
C484 VTAIL.n184 B 0.01339f
C485 VTAIL.n185 B 0.023737f
C486 VTAIL.n186 B 0.022373f
C487 VTAIL.t3 B 0.053184f
C488 VTAIL.n187 B 0.160337f
C489 VTAIL.n188 B 1.0332f
C490 VTAIL.n189 B 0.01339f
C491 VTAIL.n190 B 0.014178f
C492 VTAIL.n191 B 0.031649f
C493 VTAIL.n192 B 0.031649f
C494 VTAIL.n193 B 0.014178f
C495 VTAIL.n194 B 0.01339f
C496 VTAIL.n195 B 0.024918f
C497 VTAIL.n196 B 0.024918f
C498 VTAIL.n197 B 0.01339f
C499 VTAIL.n198 B 0.014178f
C500 VTAIL.n199 B 0.031649f
C501 VTAIL.n200 B 0.031649f
C502 VTAIL.n201 B 0.014178f
C503 VTAIL.n202 B 0.01339f
C504 VTAIL.n203 B 0.024918f
C505 VTAIL.n204 B 0.024918f
C506 VTAIL.n205 B 0.01339f
C507 VTAIL.n206 B 0.01339f
C508 VTAIL.n207 B 0.014178f
C509 VTAIL.n208 B 0.031649f
C510 VTAIL.n209 B 0.031649f
C511 VTAIL.n210 B 0.031649f
C512 VTAIL.n211 B 0.013784f
C513 VTAIL.n212 B 0.01339f
C514 VTAIL.n213 B 0.024918f
C515 VTAIL.n214 B 0.024918f
C516 VTAIL.n215 B 0.01339f
C517 VTAIL.n216 B 0.014178f
C518 VTAIL.n217 B 0.031649f
C519 VTAIL.n218 B 0.065542f
C520 VTAIL.n219 B 0.014178f
C521 VTAIL.n220 B 0.01339f
C522 VTAIL.n221 B 0.058278f
C523 VTAIL.n222 B 0.036389f
C524 VTAIL.n223 B 1.47508f
C525 VP.t5 B 1.8598f
C526 VP.n0 B 0.743307f
C527 VP.n1 B 0.021431f
C528 VP.n2 B 0.017454f
C529 VP.n3 B 0.021431f
C530 VP.t4 B 1.8598f
C531 VP.n4 B 0.661173f
C532 VP.n5 B 0.021431f
C533 VP.n6 B 0.017454f
C534 VP.n7 B 0.021431f
C535 VP.t1 B 1.8598f
C536 VP.n8 B 0.743307f
C537 VP.t3 B 1.8598f
C538 VP.n9 B 0.743307f
C539 VP.n10 B 0.021431f
C540 VP.n11 B 0.017454f
C541 VP.n12 B 0.021431f
C542 VP.t2 B 1.8598f
C543 VP.n13 B 0.732253f
C544 VP.t0 B 2.10727f
C545 VP.n14 B 0.69815f
C546 VP.n15 B 0.249785f
C547 VP.n16 B 0.030232f
C548 VP.n17 B 0.040142f
C549 VP.n18 B 0.043198f
C550 VP.n19 B 0.021431f
C551 VP.n20 B 0.021431f
C552 VP.n21 B 0.021431f
C553 VP.n22 B 0.042334f
C554 VP.n23 B 0.040142f
C555 VP.n24 B 0.031818f
C556 VP.n25 B 0.034595f
C557 VP.n26 B 1.20483f
C558 VP.n27 B 1.22031f
C559 VP.n28 B 0.034595f
C560 VP.n29 B 0.031818f
C561 VP.n30 B 0.040142f
C562 VP.n31 B 0.042334f
C563 VP.n32 B 0.021431f
C564 VP.n33 B 0.021431f
C565 VP.n34 B 0.021431f
C566 VP.n35 B 0.043198f
C567 VP.n36 B 0.040142f
C568 VP.n37 B 0.030232f
C569 VP.n38 B 0.021431f
C570 VP.n39 B 0.021431f
C571 VP.n40 B 0.030232f
C572 VP.n41 B 0.040142f
C573 VP.n42 B 0.043198f
C574 VP.n43 B 0.021431f
C575 VP.n44 B 0.021431f
C576 VP.n45 B 0.021431f
C577 VP.n46 B 0.042334f
C578 VP.n47 B 0.040142f
C579 VP.n48 B 0.031818f
C580 VP.n49 B 0.034595f
C581 VP.n50 B 0.051521f
.ends

