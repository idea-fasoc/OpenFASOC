* NGSPICE file created from diff_pair_sample_1345.ext - technology: sky130A

.subckt diff_pair_sample_1345 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=0 ps=0 w=17.51 l=3.47
X1 VDD1.t3 VP.t0 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88915 pd=17.84 as=6.8289 ps=35.8 w=17.51 l=3.47
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=0 ps=0 w=17.51 l=3.47
X3 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=2.88915 ps=17.84 w=17.51 l=3.47
X4 VTAIL.t6 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=2.88915 ps=17.84 w=17.51 l=3.47
X5 VTAIL.t5 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=2.88915 ps=17.84 w=17.51 l=3.47
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=0 ps=0 w=17.51 l=3.47
X7 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88915 pd=17.84 as=6.8289 ps=35.8 w=17.51 l=3.47
X8 VDD1.t0 VP.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88915 pd=17.84 as=6.8289 ps=35.8 w=17.51 l=3.47
X9 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88915 pd=17.84 as=6.8289 ps=35.8 w=17.51 l=3.47
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=0 ps=0 w=17.51 l=3.47
X11 VTAIL.t1 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8289 pd=35.8 as=2.88915 ps=17.84 w=17.51 l=3.47
R0 B.n970 B.n969 585
R1 B.n971 B.n970 585
R2 B.n393 B.n140 585
R3 B.n392 B.n391 585
R4 B.n390 B.n389 585
R5 B.n388 B.n387 585
R6 B.n386 B.n385 585
R7 B.n384 B.n383 585
R8 B.n382 B.n381 585
R9 B.n380 B.n379 585
R10 B.n378 B.n377 585
R11 B.n376 B.n375 585
R12 B.n374 B.n373 585
R13 B.n372 B.n371 585
R14 B.n370 B.n369 585
R15 B.n368 B.n367 585
R16 B.n366 B.n365 585
R17 B.n364 B.n363 585
R18 B.n362 B.n361 585
R19 B.n360 B.n359 585
R20 B.n358 B.n357 585
R21 B.n356 B.n355 585
R22 B.n354 B.n353 585
R23 B.n352 B.n351 585
R24 B.n350 B.n349 585
R25 B.n348 B.n347 585
R26 B.n346 B.n345 585
R27 B.n344 B.n343 585
R28 B.n342 B.n341 585
R29 B.n340 B.n339 585
R30 B.n338 B.n337 585
R31 B.n336 B.n335 585
R32 B.n334 B.n333 585
R33 B.n332 B.n331 585
R34 B.n330 B.n329 585
R35 B.n328 B.n327 585
R36 B.n326 B.n325 585
R37 B.n324 B.n323 585
R38 B.n322 B.n321 585
R39 B.n320 B.n319 585
R40 B.n318 B.n317 585
R41 B.n316 B.n315 585
R42 B.n314 B.n313 585
R43 B.n312 B.n311 585
R44 B.n310 B.n309 585
R45 B.n308 B.n307 585
R46 B.n306 B.n305 585
R47 B.n304 B.n303 585
R48 B.n302 B.n301 585
R49 B.n300 B.n299 585
R50 B.n298 B.n297 585
R51 B.n296 B.n295 585
R52 B.n294 B.n293 585
R53 B.n292 B.n291 585
R54 B.n290 B.n289 585
R55 B.n288 B.n287 585
R56 B.n286 B.n285 585
R57 B.n284 B.n283 585
R58 B.n282 B.n281 585
R59 B.n279 B.n278 585
R60 B.n277 B.n276 585
R61 B.n275 B.n274 585
R62 B.n273 B.n272 585
R63 B.n271 B.n270 585
R64 B.n269 B.n268 585
R65 B.n267 B.n266 585
R66 B.n265 B.n264 585
R67 B.n263 B.n262 585
R68 B.n261 B.n260 585
R69 B.n259 B.n258 585
R70 B.n257 B.n256 585
R71 B.n255 B.n254 585
R72 B.n253 B.n252 585
R73 B.n251 B.n250 585
R74 B.n249 B.n248 585
R75 B.n247 B.n246 585
R76 B.n245 B.n244 585
R77 B.n243 B.n242 585
R78 B.n241 B.n240 585
R79 B.n239 B.n238 585
R80 B.n237 B.n236 585
R81 B.n235 B.n234 585
R82 B.n233 B.n232 585
R83 B.n231 B.n230 585
R84 B.n229 B.n228 585
R85 B.n227 B.n226 585
R86 B.n225 B.n224 585
R87 B.n223 B.n222 585
R88 B.n221 B.n220 585
R89 B.n219 B.n218 585
R90 B.n217 B.n216 585
R91 B.n215 B.n214 585
R92 B.n213 B.n212 585
R93 B.n211 B.n210 585
R94 B.n209 B.n208 585
R95 B.n207 B.n206 585
R96 B.n205 B.n204 585
R97 B.n203 B.n202 585
R98 B.n201 B.n200 585
R99 B.n199 B.n198 585
R100 B.n197 B.n196 585
R101 B.n195 B.n194 585
R102 B.n193 B.n192 585
R103 B.n191 B.n190 585
R104 B.n189 B.n188 585
R105 B.n187 B.n186 585
R106 B.n185 B.n184 585
R107 B.n183 B.n182 585
R108 B.n181 B.n180 585
R109 B.n179 B.n178 585
R110 B.n177 B.n176 585
R111 B.n175 B.n174 585
R112 B.n173 B.n172 585
R113 B.n171 B.n170 585
R114 B.n169 B.n168 585
R115 B.n167 B.n166 585
R116 B.n165 B.n164 585
R117 B.n163 B.n162 585
R118 B.n161 B.n160 585
R119 B.n159 B.n158 585
R120 B.n157 B.n156 585
R121 B.n155 B.n154 585
R122 B.n153 B.n152 585
R123 B.n151 B.n150 585
R124 B.n149 B.n148 585
R125 B.n147 B.n146 585
R126 B.n968 B.n77 585
R127 B.n972 B.n77 585
R128 B.n967 B.n76 585
R129 B.n973 B.n76 585
R130 B.n966 B.n965 585
R131 B.n965 B.n72 585
R132 B.n964 B.n71 585
R133 B.n979 B.n71 585
R134 B.n963 B.n70 585
R135 B.n980 B.n70 585
R136 B.n962 B.n69 585
R137 B.n981 B.n69 585
R138 B.n961 B.n960 585
R139 B.n960 B.n65 585
R140 B.n959 B.n64 585
R141 B.n987 B.n64 585
R142 B.n958 B.n63 585
R143 B.n988 B.n63 585
R144 B.n957 B.n62 585
R145 B.n989 B.n62 585
R146 B.n956 B.n955 585
R147 B.n955 B.n58 585
R148 B.n954 B.n57 585
R149 B.n995 B.n57 585
R150 B.n953 B.n56 585
R151 B.n996 B.n56 585
R152 B.n952 B.n55 585
R153 B.n997 B.n55 585
R154 B.n951 B.n950 585
R155 B.n950 B.n51 585
R156 B.n949 B.n50 585
R157 B.n1003 B.n50 585
R158 B.n948 B.n49 585
R159 B.n1004 B.n49 585
R160 B.n947 B.n48 585
R161 B.n1005 B.n48 585
R162 B.n946 B.n945 585
R163 B.n945 B.n44 585
R164 B.n944 B.n43 585
R165 B.n1011 B.n43 585
R166 B.n943 B.n42 585
R167 B.n1012 B.n42 585
R168 B.n942 B.n41 585
R169 B.n1013 B.n41 585
R170 B.n941 B.n940 585
R171 B.n940 B.n37 585
R172 B.n939 B.n36 585
R173 B.n1019 B.n36 585
R174 B.n938 B.n35 585
R175 B.n1020 B.n35 585
R176 B.n937 B.n34 585
R177 B.n1021 B.n34 585
R178 B.n936 B.n935 585
R179 B.n935 B.n30 585
R180 B.n934 B.n29 585
R181 B.n1027 B.n29 585
R182 B.n933 B.n28 585
R183 B.n1028 B.n28 585
R184 B.n932 B.n27 585
R185 B.n1029 B.n27 585
R186 B.n931 B.n930 585
R187 B.n930 B.n23 585
R188 B.n929 B.n22 585
R189 B.n1035 B.n22 585
R190 B.n928 B.n21 585
R191 B.n1036 B.n21 585
R192 B.n927 B.n20 585
R193 B.n1037 B.n20 585
R194 B.n926 B.n925 585
R195 B.n925 B.n19 585
R196 B.n924 B.n15 585
R197 B.n1043 B.n15 585
R198 B.n923 B.n14 585
R199 B.n1044 B.n14 585
R200 B.n922 B.n13 585
R201 B.n1045 B.n13 585
R202 B.n921 B.n920 585
R203 B.n920 B.n12 585
R204 B.n919 B.n918 585
R205 B.n919 B.n8 585
R206 B.n917 B.n7 585
R207 B.n1052 B.n7 585
R208 B.n916 B.n6 585
R209 B.n1053 B.n6 585
R210 B.n915 B.n5 585
R211 B.n1054 B.n5 585
R212 B.n914 B.n913 585
R213 B.n913 B.n4 585
R214 B.n912 B.n394 585
R215 B.n912 B.n911 585
R216 B.n902 B.n395 585
R217 B.n396 B.n395 585
R218 B.n904 B.n903 585
R219 B.n905 B.n904 585
R220 B.n901 B.n401 585
R221 B.n401 B.n400 585
R222 B.n900 B.n899 585
R223 B.n899 B.n898 585
R224 B.n403 B.n402 585
R225 B.n891 B.n403 585
R226 B.n890 B.n889 585
R227 B.n892 B.n890 585
R228 B.n888 B.n408 585
R229 B.n408 B.n407 585
R230 B.n887 B.n886 585
R231 B.n886 B.n885 585
R232 B.n410 B.n409 585
R233 B.n411 B.n410 585
R234 B.n878 B.n877 585
R235 B.n879 B.n878 585
R236 B.n876 B.n416 585
R237 B.n416 B.n415 585
R238 B.n875 B.n874 585
R239 B.n874 B.n873 585
R240 B.n418 B.n417 585
R241 B.n419 B.n418 585
R242 B.n866 B.n865 585
R243 B.n867 B.n866 585
R244 B.n864 B.n424 585
R245 B.n424 B.n423 585
R246 B.n863 B.n862 585
R247 B.n862 B.n861 585
R248 B.n426 B.n425 585
R249 B.n427 B.n426 585
R250 B.n854 B.n853 585
R251 B.n855 B.n854 585
R252 B.n852 B.n432 585
R253 B.n432 B.n431 585
R254 B.n851 B.n850 585
R255 B.n850 B.n849 585
R256 B.n434 B.n433 585
R257 B.n435 B.n434 585
R258 B.n842 B.n841 585
R259 B.n843 B.n842 585
R260 B.n840 B.n440 585
R261 B.n440 B.n439 585
R262 B.n839 B.n838 585
R263 B.n838 B.n837 585
R264 B.n442 B.n441 585
R265 B.n443 B.n442 585
R266 B.n830 B.n829 585
R267 B.n831 B.n830 585
R268 B.n828 B.n448 585
R269 B.n448 B.n447 585
R270 B.n827 B.n826 585
R271 B.n826 B.n825 585
R272 B.n450 B.n449 585
R273 B.n451 B.n450 585
R274 B.n818 B.n817 585
R275 B.n819 B.n818 585
R276 B.n816 B.n455 585
R277 B.n459 B.n455 585
R278 B.n815 B.n814 585
R279 B.n814 B.n813 585
R280 B.n457 B.n456 585
R281 B.n458 B.n457 585
R282 B.n806 B.n805 585
R283 B.n807 B.n806 585
R284 B.n804 B.n464 585
R285 B.n464 B.n463 585
R286 B.n803 B.n802 585
R287 B.n802 B.n801 585
R288 B.n466 B.n465 585
R289 B.n467 B.n466 585
R290 B.n794 B.n793 585
R291 B.n795 B.n794 585
R292 B.n792 B.n472 585
R293 B.n472 B.n471 585
R294 B.n786 B.n785 585
R295 B.n784 B.n536 585
R296 B.n783 B.n535 585
R297 B.n788 B.n535 585
R298 B.n782 B.n781 585
R299 B.n780 B.n779 585
R300 B.n778 B.n777 585
R301 B.n776 B.n775 585
R302 B.n774 B.n773 585
R303 B.n772 B.n771 585
R304 B.n770 B.n769 585
R305 B.n768 B.n767 585
R306 B.n766 B.n765 585
R307 B.n764 B.n763 585
R308 B.n762 B.n761 585
R309 B.n760 B.n759 585
R310 B.n758 B.n757 585
R311 B.n756 B.n755 585
R312 B.n754 B.n753 585
R313 B.n752 B.n751 585
R314 B.n750 B.n749 585
R315 B.n748 B.n747 585
R316 B.n746 B.n745 585
R317 B.n744 B.n743 585
R318 B.n742 B.n741 585
R319 B.n740 B.n739 585
R320 B.n738 B.n737 585
R321 B.n736 B.n735 585
R322 B.n734 B.n733 585
R323 B.n732 B.n731 585
R324 B.n730 B.n729 585
R325 B.n728 B.n727 585
R326 B.n726 B.n725 585
R327 B.n724 B.n723 585
R328 B.n722 B.n721 585
R329 B.n720 B.n719 585
R330 B.n718 B.n717 585
R331 B.n716 B.n715 585
R332 B.n714 B.n713 585
R333 B.n712 B.n711 585
R334 B.n710 B.n709 585
R335 B.n708 B.n707 585
R336 B.n706 B.n705 585
R337 B.n704 B.n703 585
R338 B.n702 B.n701 585
R339 B.n700 B.n699 585
R340 B.n698 B.n697 585
R341 B.n696 B.n695 585
R342 B.n694 B.n693 585
R343 B.n692 B.n691 585
R344 B.n690 B.n689 585
R345 B.n688 B.n687 585
R346 B.n686 B.n685 585
R347 B.n684 B.n683 585
R348 B.n682 B.n681 585
R349 B.n680 B.n679 585
R350 B.n678 B.n677 585
R351 B.n676 B.n675 585
R352 B.n674 B.n673 585
R353 B.n671 B.n670 585
R354 B.n669 B.n668 585
R355 B.n667 B.n666 585
R356 B.n665 B.n664 585
R357 B.n663 B.n662 585
R358 B.n661 B.n660 585
R359 B.n659 B.n658 585
R360 B.n657 B.n656 585
R361 B.n655 B.n654 585
R362 B.n653 B.n652 585
R363 B.n651 B.n650 585
R364 B.n649 B.n648 585
R365 B.n647 B.n646 585
R366 B.n645 B.n644 585
R367 B.n643 B.n642 585
R368 B.n641 B.n640 585
R369 B.n639 B.n638 585
R370 B.n637 B.n636 585
R371 B.n635 B.n634 585
R372 B.n633 B.n632 585
R373 B.n631 B.n630 585
R374 B.n629 B.n628 585
R375 B.n627 B.n626 585
R376 B.n625 B.n624 585
R377 B.n623 B.n622 585
R378 B.n621 B.n620 585
R379 B.n619 B.n618 585
R380 B.n617 B.n616 585
R381 B.n615 B.n614 585
R382 B.n613 B.n612 585
R383 B.n611 B.n610 585
R384 B.n609 B.n608 585
R385 B.n607 B.n606 585
R386 B.n605 B.n604 585
R387 B.n603 B.n602 585
R388 B.n601 B.n600 585
R389 B.n599 B.n598 585
R390 B.n597 B.n596 585
R391 B.n595 B.n594 585
R392 B.n593 B.n592 585
R393 B.n591 B.n590 585
R394 B.n589 B.n588 585
R395 B.n587 B.n586 585
R396 B.n585 B.n584 585
R397 B.n583 B.n582 585
R398 B.n581 B.n580 585
R399 B.n579 B.n578 585
R400 B.n577 B.n576 585
R401 B.n575 B.n574 585
R402 B.n573 B.n572 585
R403 B.n571 B.n570 585
R404 B.n569 B.n568 585
R405 B.n567 B.n566 585
R406 B.n565 B.n564 585
R407 B.n563 B.n562 585
R408 B.n561 B.n560 585
R409 B.n559 B.n558 585
R410 B.n557 B.n556 585
R411 B.n555 B.n554 585
R412 B.n553 B.n552 585
R413 B.n551 B.n550 585
R414 B.n549 B.n548 585
R415 B.n547 B.n546 585
R416 B.n545 B.n544 585
R417 B.n543 B.n542 585
R418 B.n474 B.n473 585
R419 B.n791 B.n790 585
R420 B.n470 B.n469 585
R421 B.n471 B.n470 585
R422 B.n797 B.n796 585
R423 B.n796 B.n795 585
R424 B.n798 B.n468 585
R425 B.n468 B.n467 585
R426 B.n800 B.n799 585
R427 B.n801 B.n800 585
R428 B.n462 B.n461 585
R429 B.n463 B.n462 585
R430 B.n809 B.n808 585
R431 B.n808 B.n807 585
R432 B.n810 B.n460 585
R433 B.n460 B.n458 585
R434 B.n812 B.n811 585
R435 B.n813 B.n812 585
R436 B.n454 B.n453 585
R437 B.n459 B.n454 585
R438 B.n821 B.n820 585
R439 B.n820 B.n819 585
R440 B.n822 B.n452 585
R441 B.n452 B.n451 585
R442 B.n824 B.n823 585
R443 B.n825 B.n824 585
R444 B.n446 B.n445 585
R445 B.n447 B.n446 585
R446 B.n833 B.n832 585
R447 B.n832 B.n831 585
R448 B.n834 B.n444 585
R449 B.n444 B.n443 585
R450 B.n836 B.n835 585
R451 B.n837 B.n836 585
R452 B.n438 B.n437 585
R453 B.n439 B.n438 585
R454 B.n845 B.n844 585
R455 B.n844 B.n843 585
R456 B.n846 B.n436 585
R457 B.n436 B.n435 585
R458 B.n848 B.n847 585
R459 B.n849 B.n848 585
R460 B.n430 B.n429 585
R461 B.n431 B.n430 585
R462 B.n857 B.n856 585
R463 B.n856 B.n855 585
R464 B.n858 B.n428 585
R465 B.n428 B.n427 585
R466 B.n860 B.n859 585
R467 B.n861 B.n860 585
R468 B.n422 B.n421 585
R469 B.n423 B.n422 585
R470 B.n869 B.n868 585
R471 B.n868 B.n867 585
R472 B.n870 B.n420 585
R473 B.n420 B.n419 585
R474 B.n872 B.n871 585
R475 B.n873 B.n872 585
R476 B.n414 B.n413 585
R477 B.n415 B.n414 585
R478 B.n881 B.n880 585
R479 B.n880 B.n879 585
R480 B.n882 B.n412 585
R481 B.n412 B.n411 585
R482 B.n884 B.n883 585
R483 B.n885 B.n884 585
R484 B.n406 B.n405 585
R485 B.n407 B.n406 585
R486 B.n894 B.n893 585
R487 B.n893 B.n892 585
R488 B.n895 B.n404 585
R489 B.n891 B.n404 585
R490 B.n897 B.n896 585
R491 B.n898 B.n897 585
R492 B.n399 B.n398 585
R493 B.n400 B.n399 585
R494 B.n907 B.n906 585
R495 B.n906 B.n905 585
R496 B.n908 B.n397 585
R497 B.n397 B.n396 585
R498 B.n910 B.n909 585
R499 B.n911 B.n910 585
R500 B.n3 B.n0 585
R501 B.n4 B.n3 585
R502 B.n1051 B.n1 585
R503 B.n1052 B.n1051 585
R504 B.n1050 B.n1049 585
R505 B.n1050 B.n8 585
R506 B.n1048 B.n9 585
R507 B.n12 B.n9 585
R508 B.n1047 B.n1046 585
R509 B.n1046 B.n1045 585
R510 B.n11 B.n10 585
R511 B.n1044 B.n11 585
R512 B.n1042 B.n1041 585
R513 B.n1043 B.n1042 585
R514 B.n1040 B.n16 585
R515 B.n19 B.n16 585
R516 B.n1039 B.n1038 585
R517 B.n1038 B.n1037 585
R518 B.n18 B.n17 585
R519 B.n1036 B.n18 585
R520 B.n1034 B.n1033 585
R521 B.n1035 B.n1034 585
R522 B.n1032 B.n24 585
R523 B.n24 B.n23 585
R524 B.n1031 B.n1030 585
R525 B.n1030 B.n1029 585
R526 B.n26 B.n25 585
R527 B.n1028 B.n26 585
R528 B.n1026 B.n1025 585
R529 B.n1027 B.n1026 585
R530 B.n1024 B.n31 585
R531 B.n31 B.n30 585
R532 B.n1023 B.n1022 585
R533 B.n1022 B.n1021 585
R534 B.n33 B.n32 585
R535 B.n1020 B.n33 585
R536 B.n1018 B.n1017 585
R537 B.n1019 B.n1018 585
R538 B.n1016 B.n38 585
R539 B.n38 B.n37 585
R540 B.n1015 B.n1014 585
R541 B.n1014 B.n1013 585
R542 B.n40 B.n39 585
R543 B.n1012 B.n40 585
R544 B.n1010 B.n1009 585
R545 B.n1011 B.n1010 585
R546 B.n1008 B.n45 585
R547 B.n45 B.n44 585
R548 B.n1007 B.n1006 585
R549 B.n1006 B.n1005 585
R550 B.n47 B.n46 585
R551 B.n1004 B.n47 585
R552 B.n1002 B.n1001 585
R553 B.n1003 B.n1002 585
R554 B.n1000 B.n52 585
R555 B.n52 B.n51 585
R556 B.n999 B.n998 585
R557 B.n998 B.n997 585
R558 B.n54 B.n53 585
R559 B.n996 B.n54 585
R560 B.n994 B.n993 585
R561 B.n995 B.n994 585
R562 B.n992 B.n59 585
R563 B.n59 B.n58 585
R564 B.n991 B.n990 585
R565 B.n990 B.n989 585
R566 B.n61 B.n60 585
R567 B.n988 B.n61 585
R568 B.n986 B.n985 585
R569 B.n987 B.n986 585
R570 B.n984 B.n66 585
R571 B.n66 B.n65 585
R572 B.n983 B.n982 585
R573 B.n982 B.n981 585
R574 B.n68 B.n67 585
R575 B.n980 B.n68 585
R576 B.n978 B.n977 585
R577 B.n979 B.n978 585
R578 B.n976 B.n73 585
R579 B.n73 B.n72 585
R580 B.n975 B.n974 585
R581 B.n974 B.n973 585
R582 B.n75 B.n74 585
R583 B.n972 B.n75 585
R584 B.n1055 B.n1054 585
R585 B.n1053 B.n2 585
R586 B.n146 B.n75 540.549
R587 B.n970 B.n77 540.549
R588 B.n790 B.n472 540.549
R589 B.n786 B.n470 540.549
R590 B.n143 B.t9 450.762
R591 B.n141 B.t6 450.762
R592 B.n539 B.t17 450.762
R593 B.n537 B.t14 450.762
R594 B.n142 B.t7 377.065
R595 B.n540 B.t16 377.065
R596 B.n144 B.t10 377.065
R597 B.n538 B.t13 377.065
R598 B.n143 B.t8 330.678
R599 B.n141 B.t4 330.678
R600 B.n539 B.t15 330.678
R601 B.n537 B.t11 330.678
R602 B.n971 B.n139 256.663
R603 B.n971 B.n138 256.663
R604 B.n971 B.n137 256.663
R605 B.n971 B.n136 256.663
R606 B.n971 B.n135 256.663
R607 B.n971 B.n134 256.663
R608 B.n971 B.n133 256.663
R609 B.n971 B.n132 256.663
R610 B.n971 B.n131 256.663
R611 B.n971 B.n130 256.663
R612 B.n971 B.n129 256.663
R613 B.n971 B.n128 256.663
R614 B.n971 B.n127 256.663
R615 B.n971 B.n126 256.663
R616 B.n971 B.n125 256.663
R617 B.n971 B.n124 256.663
R618 B.n971 B.n123 256.663
R619 B.n971 B.n122 256.663
R620 B.n971 B.n121 256.663
R621 B.n971 B.n120 256.663
R622 B.n971 B.n119 256.663
R623 B.n971 B.n118 256.663
R624 B.n971 B.n117 256.663
R625 B.n971 B.n116 256.663
R626 B.n971 B.n115 256.663
R627 B.n971 B.n114 256.663
R628 B.n971 B.n113 256.663
R629 B.n971 B.n112 256.663
R630 B.n971 B.n111 256.663
R631 B.n971 B.n110 256.663
R632 B.n971 B.n109 256.663
R633 B.n971 B.n108 256.663
R634 B.n971 B.n107 256.663
R635 B.n971 B.n106 256.663
R636 B.n971 B.n105 256.663
R637 B.n971 B.n104 256.663
R638 B.n971 B.n103 256.663
R639 B.n971 B.n102 256.663
R640 B.n971 B.n101 256.663
R641 B.n971 B.n100 256.663
R642 B.n971 B.n99 256.663
R643 B.n971 B.n98 256.663
R644 B.n971 B.n97 256.663
R645 B.n971 B.n96 256.663
R646 B.n971 B.n95 256.663
R647 B.n971 B.n94 256.663
R648 B.n971 B.n93 256.663
R649 B.n971 B.n92 256.663
R650 B.n971 B.n91 256.663
R651 B.n971 B.n90 256.663
R652 B.n971 B.n89 256.663
R653 B.n971 B.n88 256.663
R654 B.n971 B.n87 256.663
R655 B.n971 B.n86 256.663
R656 B.n971 B.n85 256.663
R657 B.n971 B.n84 256.663
R658 B.n971 B.n83 256.663
R659 B.n971 B.n82 256.663
R660 B.n971 B.n81 256.663
R661 B.n971 B.n80 256.663
R662 B.n971 B.n79 256.663
R663 B.n971 B.n78 256.663
R664 B.n788 B.n787 256.663
R665 B.n788 B.n475 256.663
R666 B.n788 B.n476 256.663
R667 B.n788 B.n477 256.663
R668 B.n788 B.n478 256.663
R669 B.n788 B.n479 256.663
R670 B.n788 B.n480 256.663
R671 B.n788 B.n481 256.663
R672 B.n788 B.n482 256.663
R673 B.n788 B.n483 256.663
R674 B.n788 B.n484 256.663
R675 B.n788 B.n485 256.663
R676 B.n788 B.n486 256.663
R677 B.n788 B.n487 256.663
R678 B.n788 B.n488 256.663
R679 B.n788 B.n489 256.663
R680 B.n788 B.n490 256.663
R681 B.n788 B.n491 256.663
R682 B.n788 B.n492 256.663
R683 B.n788 B.n493 256.663
R684 B.n788 B.n494 256.663
R685 B.n788 B.n495 256.663
R686 B.n788 B.n496 256.663
R687 B.n788 B.n497 256.663
R688 B.n788 B.n498 256.663
R689 B.n788 B.n499 256.663
R690 B.n788 B.n500 256.663
R691 B.n788 B.n501 256.663
R692 B.n788 B.n502 256.663
R693 B.n788 B.n503 256.663
R694 B.n788 B.n504 256.663
R695 B.n788 B.n505 256.663
R696 B.n788 B.n506 256.663
R697 B.n788 B.n507 256.663
R698 B.n788 B.n508 256.663
R699 B.n788 B.n509 256.663
R700 B.n788 B.n510 256.663
R701 B.n788 B.n511 256.663
R702 B.n788 B.n512 256.663
R703 B.n788 B.n513 256.663
R704 B.n788 B.n514 256.663
R705 B.n788 B.n515 256.663
R706 B.n788 B.n516 256.663
R707 B.n788 B.n517 256.663
R708 B.n788 B.n518 256.663
R709 B.n788 B.n519 256.663
R710 B.n788 B.n520 256.663
R711 B.n788 B.n521 256.663
R712 B.n788 B.n522 256.663
R713 B.n788 B.n523 256.663
R714 B.n788 B.n524 256.663
R715 B.n788 B.n525 256.663
R716 B.n788 B.n526 256.663
R717 B.n788 B.n527 256.663
R718 B.n788 B.n528 256.663
R719 B.n788 B.n529 256.663
R720 B.n788 B.n530 256.663
R721 B.n788 B.n531 256.663
R722 B.n788 B.n532 256.663
R723 B.n788 B.n533 256.663
R724 B.n788 B.n534 256.663
R725 B.n789 B.n788 256.663
R726 B.n1057 B.n1056 256.663
R727 B.n150 B.n149 163.367
R728 B.n154 B.n153 163.367
R729 B.n158 B.n157 163.367
R730 B.n162 B.n161 163.367
R731 B.n166 B.n165 163.367
R732 B.n170 B.n169 163.367
R733 B.n174 B.n173 163.367
R734 B.n178 B.n177 163.367
R735 B.n182 B.n181 163.367
R736 B.n186 B.n185 163.367
R737 B.n190 B.n189 163.367
R738 B.n194 B.n193 163.367
R739 B.n198 B.n197 163.367
R740 B.n202 B.n201 163.367
R741 B.n206 B.n205 163.367
R742 B.n210 B.n209 163.367
R743 B.n214 B.n213 163.367
R744 B.n218 B.n217 163.367
R745 B.n222 B.n221 163.367
R746 B.n226 B.n225 163.367
R747 B.n230 B.n229 163.367
R748 B.n234 B.n233 163.367
R749 B.n238 B.n237 163.367
R750 B.n242 B.n241 163.367
R751 B.n246 B.n245 163.367
R752 B.n250 B.n249 163.367
R753 B.n254 B.n253 163.367
R754 B.n258 B.n257 163.367
R755 B.n262 B.n261 163.367
R756 B.n266 B.n265 163.367
R757 B.n270 B.n269 163.367
R758 B.n274 B.n273 163.367
R759 B.n278 B.n277 163.367
R760 B.n283 B.n282 163.367
R761 B.n287 B.n286 163.367
R762 B.n291 B.n290 163.367
R763 B.n295 B.n294 163.367
R764 B.n299 B.n298 163.367
R765 B.n303 B.n302 163.367
R766 B.n307 B.n306 163.367
R767 B.n311 B.n310 163.367
R768 B.n315 B.n314 163.367
R769 B.n319 B.n318 163.367
R770 B.n323 B.n322 163.367
R771 B.n327 B.n326 163.367
R772 B.n331 B.n330 163.367
R773 B.n335 B.n334 163.367
R774 B.n339 B.n338 163.367
R775 B.n343 B.n342 163.367
R776 B.n347 B.n346 163.367
R777 B.n351 B.n350 163.367
R778 B.n355 B.n354 163.367
R779 B.n359 B.n358 163.367
R780 B.n363 B.n362 163.367
R781 B.n367 B.n366 163.367
R782 B.n371 B.n370 163.367
R783 B.n375 B.n374 163.367
R784 B.n379 B.n378 163.367
R785 B.n383 B.n382 163.367
R786 B.n387 B.n386 163.367
R787 B.n391 B.n390 163.367
R788 B.n970 B.n140 163.367
R789 B.n794 B.n472 163.367
R790 B.n794 B.n466 163.367
R791 B.n802 B.n466 163.367
R792 B.n802 B.n464 163.367
R793 B.n806 B.n464 163.367
R794 B.n806 B.n457 163.367
R795 B.n814 B.n457 163.367
R796 B.n814 B.n455 163.367
R797 B.n818 B.n455 163.367
R798 B.n818 B.n450 163.367
R799 B.n826 B.n450 163.367
R800 B.n826 B.n448 163.367
R801 B.n830 B.n448 163.367
R802 B.n830 B.n442 163.367
R803 B.n838 B.n442 163.367
R804 B.n838 B.n440 163.367
R805 B.n842 B.n440 163.367
R806 B.n842 B.n434 163.367
R807 B.n850 B.n434 163.367
R808 B.n850 B.n432 163.367
R809 B.n854 B.n432 163.367
R810 B.n854 B.n426 163.367
R811 B.n862 B.n426 163.367
R812 B.n862 B.n424 163.367
R813 B.n866 B.n424 163.367
R814 B.n866 B.n418 163.367
R815 B.n874 B.n418 163.367
R816 B.n874 B.n416 163.367
R817 B.n878 B.n416 163.367
R818 B.n878 B.n410 163.367
R819 B.n886 B.n410 163.367
R820 B.n886 B.n408 163.367
R821 B.n890 B.n408 163.367
R822 B.n890 B.n403 163.367
R823 B.n899 B.n403 163.367
R824 B.n899 B.n401 163.367
R825 B.n904 B.n401 163.367
R826 B.n904 B.n395 163.367
R827 B.n912 B.n395 163.367
R828 B.n913 B.n912 163.367
R829 B.n913 B.n5 163.367
R830 B.n6 B.n5 163.367
R831 B.n7 B.n6 163.367
R832 B.n919 B.n7 163.367
R833 B.n920 B.n919 163.367
R834 B.n920 B.n13 163.367
R835 B.n14 B.n13 163.367
R836 B.n15 B.n14 163.367
R837 B.n925 B.n15 163.367
R838 B.n925 B.n20 163.367
R839 B.n21 B.n20 163.367
R840 B.n22 B.n21 163.367
R841 B.n930 B.n22 163.367
R842 B.n930 B.n27 163.367
R843 B.n28 B.n27 163.367
R844 B.n29 B.n28 163.367
R845 B.n935 B.n29 163.367
R846 B.n935 B.n34 163.367
R847 B.n35 B.n34 163.367
R848 B.n36 B.n35 163.367
R849 B.n940 B.n36 163.367
R850 B.n940 B.n41 163.367
R851 B.n42 B.n41 163.367
R852 B.n43 B.n42 163.367
R853 B.n945 B.n43 163.367
R854 B.n945 B.n48 163.367
R855 B.n49 B.n48 163.367
R856 B.n50 B.n49 163.367
R857 B.n950 B.n50 163.367
R858 B.n950 B.n55 163.367
R859 B.n56 B.n55 163.367
R860 B.n57 B.n56 163.367
R861 B.n955 B.n57 163.367
R862 B.n955 B.n62 163.367
R863 B.n63 B.n62 163.367
R864 B.n64 B.n63 163.367
R865 B.n960 B.n64 163.367
R866 B.n960 B.n69 163.367
R867 B.n70 B.n69 163.367
R868 B.n71 B.n70 163.367
R869 B.n965 B.n71 163.367
R870 B.n965 B.n76 163.367
R871 B.n77 B.n76 163.367
R872 B.n536 B.n535 163.367
R873 B.n781 B.n535 163.367
R874 B.n779 B.n778 163.367
R875 B.n775 B.n774 163.367
R876 B.n771 B.n770 163.367
R877 B.n767 B.n766 163.367
R878 B.n763 B.n762 163.367
R879 B.n759 B.n758 163.367
R880 B.n755 B.n754 163.367
R881 B.n751 B.n750 163.367
R882 B.n747 B.n746 163.367
R883 B.n743 B.n742 163.367
R884 B.n739 B.n738 163.367
R885 B.n735 B.n734 163.367
R886 B.n731 B.n730 163.367
R887 B.n727 B.n726 163.367
R888 B.n723 B.n722 163.367
R889 B.n719 B.n718 163.367
R890 B.n715 B.n714 163.367
R891 B.n711 B.n710 163.367
R892 B.n707 B.n706 163.367
R893 B.n703 B.n702 163.367
R894 B.n699 B.n698 163.367
R895 B.n695 B.n694 163.367
R896 B.n691 B.n690 163.367
R897 B.n687 B.n686 163.367
R898 B.n683 B.n682 163.367
R899 B.n679 B.n678 163.367
R900 B.n675 B.n674 163.367
R901 B.n670 B.n669 163.367
R902 B.n666 B.n665 163.367
R903 B.n662 B.n661 163.367
R904 B.n658 B.n657 163.367
R905 B.n654 B.n653 163.367
R906 B.n650 B.n649 163.367
R907 B.n646 B.n645 163.367
R908 B.n642 B.n641 163.367
R909 B.n638 B.n637 163.367
R910 B.n634 B.n633 163.367
R911 B.n630 B.n629 163.367
R912 B.n626 B.n625 163.367
R913 B.n622 B.n621 163.367
R914 B.n618 B.n617 163.367
R915 B.n614 B.n613 163.367
R916 B.n610 B.n609 163.367
R917 B.n606 B.n605 163.367
R918 B.n602 B.n601 163.367
R919 B.n598 B.n597 163.367
R920 B.n594 B.n593 163.367
R921 B.n590 B.n589 163.367
R922 B.n586 B.n585 163.367
R923 B.n582 B.n581 163.367
R924 B.n578 B.n577 163.367
R925 B.n574 B.n573 163.367
R926 B.n570 B.n569 163.367
R927 B.n566 B.n565 163.367
R928 B.n562 B.n561 163.367
R929 B.n558 B.n557 163.367
R930 B.n554 B.n553 163.367
R931 B.n550 B.n549 163.367
R932 B.n546 B.n545 163.367
R933 B.n542 B.n474 163.367
R934 B.n796 B.n470 163.367
R935 B.n796 B.n468 163.367
R936 B.n800 B.n468 163.367
R937 B.n800 B.n462 163.367
R938 B.n808 B.n462 163.367
R939 B.n808 B.n460 163.367
R940 B.n812 B.n460 163.367
R941 B.n812 B.n454 163.367
R942 B.n820 B.n454 163.367
R943 B.n820 B.n452 163.367
R944 B.n824 B.n452 163.367
R945 B.n824 B.n446 163.367
R946 B.n832 B.n446 163.367
R947 B.n832 B.n444 163.367
R948 B.n836 B.n444 163.367
R949 B.n836 B.n438 163.367
R950 B.n844 B.n438 163.367
R951 B.n844 B.n436 163.367
R952 B.n848 B.n436 163.367
R953 B.n848 B.n430 163.367
R954 B.n856 B.n430 163.367
R955 B.n856 B.n428 163.367
R956 B.n860 B.n428 163.367
R957 B.n860 B.n422 163.367
R958 B.n868 B.n422 163.367
R959 B.n868 B.n420 163.367
R960 B.n872 B.n420 163.367
R961 B.n872 B.n414 163.367
R962 B.n880 B.n414 163.367
R963 B.n880 B.n412 163.367
R964 B.n884 B.n412 163.367
R965 B.n884 B.n406 163.367
R966 B.n893 B.n406 163.367
R967 B.n893 B.n404 163.367
R968 B.n897 B.n404 163.367
R969 B.n897 B.n399 163.367
R970 B.n906 B.n399 163.367
R971 B.n906 B.n397 163.367
R972 B.n910 B.n397 163.367
R973 B.n910 B.n3 163.367
R974 B.n1055 B.n3 163.367
R975 B.n1051 B.n2 163.367
R976 B.n1051 B.n1050 163.367
R977 B.n1050 B.n9 163.367
R978 B.n1046 B.n9 163.367
R979 B.n1046 B.n11 163.367
R980 B.n1042 B.n11 163.367
R981 B.n1042 B.n16 163.367
R982 B.n1038 B.n16 163.367
R983 B.n1038 B.n18 163.367
R984 B.n1034 B.n18 163.367
R985 B.n1034 B.n24 163.367
R986 B.n1030 B.n24 163.367
R987 B.n1030 B.n26 163.367
R988 B.n1026 B.n26 163.367
R989 B.n1026 B.n31 163.367
R990 B.n1022 B.n31 163.367
R991 B.n1022 B.n33 163.367
R992 B.n1018 B.n33 163.367
R993 B.n1018 B.n38 163.367
R994 B.n1014 B.n38 163.367
R995 B.n1014 B.n40 163.367
R996 B.n1010 B.n40 163.367
R997 B.n1010 B.n45 163.367
R998 B.n1006 B.n45 163.367
R999 B.n1006 B.n47 163.367
R1000 B.n1002 B.n47 163.367
R1001 B.n1002 B.n52 163.367
R1002 B.n998 B.n52 163.367
R1003 B.n998 B.n54 163.367
R1004 B.n994 B.n54 163.367
R1005 B.n994 B.n59 163.367
R1006 B.n990 B.n59 163.367
R1007 B.n990 B.n61 163.367
R1008 B.n986 B.n61 163.367
R1009 B.n986 B.n66 163.367
R1010 B.n982 B.n66 163.367
R1011 B.n982 B.n68 163.367
R1012 B.n978 B.n68 163.367
R1013 B.n978 B.n73 163.367
R1014 B.n974 B.n73 163.367
R1015 B.n974 B.n75 163.367
R1016 B.n144 B.n143 73.6975
R1017 B.n142 B.n141 73.6975
R1018 B.n540 B.n539 73.6975
R1019 B.n538 B.n537 73.6975
R1020 B.n146 B.n78 71.676
R1021 B.n150 B.n79 71.676
R1022 B.n154 B.n80 71.676
R1023 B.n158 B.n81 71.676
R1024 B.n162 B.n82 71.676
R1025 B.n166 B.n83 71.676
R1026 B.n170 B.n84 71.676
R1027 B.n174 B.n85 71.676
R1028 B.n178 B.n86 71.676
R1029 B.n182 B.n87 71.676
R1030 B.n186 B.n88 71.676
R1031 B.n190 B.n89 71.676
R1032 B.n194 B.n90 71.676
R1033 B.n198 B.n91 71.676
R1034 B.n202 B.n92 71.676
R1035 B.n206 B.n93 71.676
R1036 B.n210 B.n94 71.676
R1037 B.n214 B.n95 71.676
R1038 B.n218 B.n96 71.676
R1039 B.n222 B.n97 71.676
R1040 B.n226 B.n98 71.676
R1041 B.n230 B.n99 71.676
R1042 B.n234 B.n100 71.676
R1043 B.n238 B.n101 71.676
R1044 B.n242 B.n102 71.676
R1045 B.n246 B.n103 71.676
R1046 B.n250 B.n104 71.676
R1047 B.n254 B.n105 71.676
R1048 B.n258 B.n106 71.676
R1049 B.n262 B.n107 71.676
R1050 B.n266 B.n108 71.676
R1051 B.n270 B.n109 71.676
R1052 B.n274 B.n110 71.676
R1053 B.n278 B.n111 71.676
R1054 B.n283 B.n112 71.676
R1055 B.n287 B.n113 71.676
R1056 B.n291 B.n114 71.676
R1057 B.n295 B.n115 71.676
R1058 B.n299 B.n116 71.676
R1059 B.n303 B.n117 71.676
R1060 B.n307 B.n118 71.676
R1061 B.n311 B.n119 71.676
R1062 B.n315 B.n120 71.676
R1063 B.n319 B.n121 71.676
R1064 B.n323 B.n122 71.676
R1065 B.n327 B.n123 71.676
R1066 B.n331 B.n124 71.676
R1067 B.n335 B.n125 71.676
R1068 B.n339 B.n126 71.676
R1069 B.n343 B.n127 71.676
R1070 B.n347 B.n128 71.676
R1071 B.n351 B.n129 71.676
R1072 B.n355 B.n130 71.676
R1073 B.n359 B.n131 71.676
R1074 B.n363 B.n132 71.676
R1075 B.n367 B.n133 71.676
R1076 B.n371 B.n134 71.676
R1077 B.n375 B.n135 71.676
R1078 B.n379 B.n136 71.676
R1079 B.n383 B.n137 71.676
R1080 B.n387 B.n138 71.676
R1081 B.n391 B.n139 71.676
R1082 B.n140 B.n139 71.676
R1083 B.n390 B.n138 71.676
R1084 B.n386 B.n137 71.676
R1085 B.n382 B.n136 71.676
R1086 B.n378 B.n135 71.676
R1087 B.n374 B.n134 71.676
R1088 B.n370 B.n133 71.676
R1089 B.n366 B.n132 71.676
R1090 B.n362 B.n131 71.676
R1091 B.n358 B.n130 71.676
R1092 B.n354 B.n129 71.676
R1093 B.n350 B.n128 71.676
R1094 B.n346 B.n127 71.676
R1095 B.n342 B.n126 71.676
R1096 B.n338 B.n125 71.676
R1097 B.n334 B.n124 71.676
R1098 B.n330 B.n123 71.676
R1099 B.n326 B.n122 71.676
R1100 B.n322 B.n121 71.676
R1101 B.n318 B.n120 71.676
R1102 B.n314 B.n119 71.676
R1103 B.n310 B.n118 71.676
R1104 B.n306 B.n117 71.676
R1105 B.n302 B.n116 71.676
R1106 B.n298 B.n115 71.676
R1107 B.n294 B.n114 71.676
R1108 B.n290 B.n113 71.676
R1109 B.n286 B.n112 71.676
R1110 B.n282 B.n111 71.676
R1111 B.n277 B.n110 71.676
R1112 B.n273 B.n109 71.676
R1113 B.n269 B.n108 71.676
R1114 B.n265 B.n107 71.676
R1115 B.n261 B.n106 71.676
R1116 B.n257 B.n105 71.676
R1117 B.n253 B.n104 71.676
R1118 B.n249 B.n103 71.676
R1119 B.n245 B.n102 71.676
R1120 B.n241 B.n101 71.676
R1121 B.n237 B.n100 71.676
R1122 B.n233 B.n99 71.676
R1123 B.n229 B.n98 71.676
R1124 B.n225 B.n97 71.676
R1125 B.n221 B.n96 71.676
R1126 B.n217 B.n95 71.676
R1127 B.n213 B.n94 71.676
R1128 B.n209 B.n93 71.676
R1129 B.n205 B.n92 71.676
R1130 B.n201 B.n91 71.676
R1131 B.n197 B.n90 71.676
R1132 B.n193 B.n89 71.676
R1133 B.n189 B.n88 71.676
R1134 B.n185 B.n87 71.676
R1135 B.n181 B.n86 71.676
R1136 B.n177 B.n85 71.676
R1137 B.n173 B.n84 71.676
R1138 B.n169 B.n83 71.676
R1139 B.n165 B.n82 71.676
R1140 B.n161 B.n81 71.676
R1141 B.n157 B.n80 71.676
R1142 B.n153 B.n79 71.676
R1143 B.n149 B.n78 71.676
R1144 B.n787 B.n786 71.676
R1145 B.n781 B.n475 71.676
R1146 B.n778 B.n476 71.676
R1147 B.n774 B.n477 71.676
R1148 B.n770 B.n478 71.676
R1149 B.n766 B.n479 71.676
R1150 B.n762 B.n480 71.676
R1151 B.n758 B.n481 71.676
R1152 B.n754 B.n482 71.676
R1153 B.n750 B.n483 71.676
R1154 B.n746 B.n484 71.676
R1155 B.n742 B.n485 71.676
R1156 B.n738 B.n486 71.676
R1157 B.n734 B.n487 71.676
R1158 B.n730 B.n488 71.676
R1159 B.n726 B.n489 71.676
R1160 B.n722 B.n490 71.676
R1161 B.n718 B.n491 71.676
R1162 B.n714 B.n492 71.676
R1163 B.n710 B.n493 71.676
R1164 B.n706 B.n494 71.676
R1165 B.n702 B.n495 71.676
R1166 B.n698 B.n496 71.676
R1167 B.n694 B.n497 71.676
R1168 B.n690 B.n498 71.676
R1169 B.n686 B.n499 71.676
R1170 B.n682 B.n500 71.676
R1171 B.n678 B.n501 71.676
R1172 B.n674 B.n502 71.676
R1173 B.n669 B.n503 71.676
R1174 B.n665 B.n504 71.676
R1175 B.n661 B.n505 71.676
R1176 B.n657 B.n506 71.676
R1177 B.n653 B.n507 71.676
R1178 B.n649 B.n508 71.676
R1179 B.n645 B.n509 71.676
R1180 B.n641 B.n510 71.676
R1181 B.n637 B.n511 71.676
R1182 B.n633 B.n512 71.676
R1183 B.n629 B.n513 71.676
R1184 B.n625 B.n514 71.676
R1185 B.n621 B.n515 71.676
R1186 B.n617 B.n516 71.676
R1187 B.n613 B.n517 71.676
R1188 B.n609 B.n518 71.676
R1189 B.n605 B.n519 71.676
R1190 B.n601 B.n520 71.676
R1191 B.n597 B.n521 71.676
R1192 B.n593 B.n522 71.676
R1193 B.n589 B.n523 71.676
R1194 B.n585 B.n524 71.676
R1195 B.n581 B.n525 71.676
R1196 B.n577 B.n526 71.676
R1197 B.n573 B.n527 71.676
R1198 B.n569 B.n528 71.676
R1199 B.n565 B.n529 71.676
R1200 B.n561 B.n530 71.676
R1201 B.n557 B.n531 71.676
R1202 B.n553 B.n532 71.676
R1203 B.n549 B.n533 71.676
R1204 B.n545 B.n534 71.676
R1205 B.n789 B.n474 71.676
R1206 B.n787 B.n536 71.676
R1207 B.n779 B.n475 71.676
R1208 B.n775 B.n476 71.676
R1209 B.n771 B.n477 71.676
R1210 B.n767 B.n478 71.676
R1211 B.n763 B.n479 71.676
R1212 B.n759 B.n480 71.676
R1213 B.n755 B.n481 71.676
R1214 B.n751 B.n482 71.676
R1215 B.n747 B.n483 71.676
R1216 B.n743 B.n484 71.676
R1217 B.n739 B.n485 71.676
R1218 B.n735 B.n486 71.676
R1219 B.n731 B.n487 71.676
R1220 B.n727 B.n488 71.676
R1221 B.n723 B.n489 71.676
R1222 B.n719 B.n490 71.676
R1223 B.n715 B.n491 71.676
R1224 B.n711 B.n492 71.676
R1225 B.n707 B.n493 71.676
R1226 B.n703 B.n494 71.676
R1227 B.n699 B.n495 71.676
R1228 B.n695 B.n496 71.676
R1229 B.n691 B.n497 71.676
R1230 B.n687 B.n498 71.676
R1231 B.n683 B.n499 71.676
R1232 B.n679 B.n500 71.676
R1233 B.n675 B.n501 71.676
R1234 B.n670 B.n502 71.676
R1235 B.n666 B.n503 71.676
R1236 B.n662 B.n504 71.676
R1237 B.n658 B.n505 71.676
R1238 B.n654 B.n506 71.676
R1239 B.n650 B.n507 71.676
R1240 B.n646 B.n508 71.676
R1241 B.n642 B.n509 71.676
R1242 B.n638 B.n510 71.676
R1243 B.n634 B.n511 71.676
R1244 B.n630 B.n512 71.676
R1245 B.n626 B.n513 71.676
R1246 B.n622 B.n514 71.676
R1247 B.n618 B.n515 71.676
R1248 B.n614 B.n516 71.676
R1249 B.n610 B.n517 71.676
R1250 B.n606 B.n518 71.676
R1251 B.n602 B.n519 71.676
R1252 B.n598 B.n520 71.676
R1253 B.n594 B.n521 71.676
R1254 B.n590 B.n522 71.676
R1255 B.n586 B.n523 71.676
R1256 B.n582 B.n524 71.676
R1257 B.n578 B.n525 71.676
R1258 B.n574 B.n526 71.676
R1259 B.n570 B.n527 71.676
R1260 B.n566 B.n528 71.676
R1261 B.n562 B.n529 71.676
R1262 B.n558 B.n530 71.676
R1263 B.n554 B.n531 71.676
R1264 B.n550 B.n532 71.676
R1265 B.n546 B.n533 71.676
R1266 B.n542 B.n534 71.676
R1267 B.n790 B.n789 71.676
R1268 B.n1056 B.n1055 71.676
R1269 B.n1056 B.n2 71.676
R1270 B.n788 B.n471 64.2094
R1271 B.n972 B.n971 64.2094
R1272 B.n145 B.n144 59.5399
R1273 B.n280 B.n142 59.5399
R1274 B.n541 B.n540 59.5399
R1275 B.n672 B.n538 59.5399
R1276 B.n785 B.n469 35.1225
R1277 B.n792 B.n791 35.1225
R1278 B.n969 B.n968 35.1225
R1279 B.n147 B.n74 35.1225
R1280 B.n795 B.n471 32.8291
R1281 B.n795 B.n467 32.8291
R1282 B.n801 B.n467 32.8291
R1283 B.n801 B.n463 32.8291
R1284 B.n807 B.n463 32.8291
R1285 B.n807 B.n458 32.8291
R1286 B.n813 B.n458 32.8291
R1287 B.n813 B.n459 32.8291
R1288 B.n819 B.n451 32.8291
R1289 B.n825 B.n451 32.8291
R1290 B.n825 B.n447 32.8291
R1291 B.n831 B.n447 32.8291
R1292 B.n831 B.n443 32.8291
R1293 B.n837 B.n443 32.8291
R1294 B.n837 B.n439 32.8291
R1295 B.n843 B.n439 32.8291
R1296 B.n843 B.n435 32.8291
R1297 B.n849 B.n435 32.8291
R1298 B.n849 B.n431 32.8291
R1299 B.n855 B.n431 32.8291
R1300 B.n855 B.n427 32.8291
R1301 B.n861 B.n427 32.8291
R1302 B.n867 B.n423 32.8291
R1303 B.n867 B.n419 32.8291
R1304 B.n873 B.n419 32.8291
R1305 B.n873 B.n415 32.8291
R1306 B.n879 B.n415 32.8291
R1307 B.n879 B.n411 32.8291
R1308 B.n885 B.n411 32.8291
R1309 B.n885 B.n407 32.8291
R1310 B.n892 B.n407 32.8291
R1311 B.n892 B.n891 32.8291
R1312 B.n898 B.n400 32.8291
R1313 B.n905 B.n400 32.8291
R1314 B.n905 B.n396 32.8291
R1315 B.n911 B.n396 32.8291
R1316 B.n911 B.n4 32.8291
R1317 B.n1054 B.n4 32.8291
R1318 B.n1054 B.n1053 32.8291
R1319 B.n1053 B.n1052 32.8291
R1320 B.n1052 B.n8 32.8291
R1321 B.n12 B.n8 32.8291
R1322 B.n1045 B.n12 32.8291
R1323 B.n1045 B.n1044 32.8291
R1324 B.n1044 B.n1043 32.8291
R1325 B.n1037 B.n19 32.8291
R1326 B.n1037 B.n1036 32.8291
R1327 B.n1036 B.n1035 32.8291
R1328 B.n1035 B.n23 32.8291
R1329 B.n1029 B.n23 32.8291
R1330 B.n1029 B.n1028 32.8291
R1331 B.n1028 B.n1027 32.8291
R1332 B.n1027 B.n30 32.8291
R1333 B.n1021 B.n30 32.8291
R1334 B.n1021 B.n1020 32.8291
R1335 B.n1019 B.n37 32.8291
R1336 B.n1013 B.n37 32.8291
R1337 B.n1013 B.n1012 32.8291
R1338 B.n1012 B.n1011 32.8291
R1339 B.n1011 B.n44 32.8291
R1340 B.n1005 B.n44 32.8291
R1341 B.n1005 B.n1004 32.8291
R1342 B.n1004 B.n1003 32.8291
R1343 B.n1003 B.n51 32.8291
R1344 B.n997 B.n51 32.8291
R1345 B.n997 B.n996 32.8291
R1346 B.n996 B.n995 32.8291
R1347 B.n995 B.n58 32.8291
R1348 B.n989 B.n58 32.8291
R1349 B.n988 B.n987 32.8291
R1350 B.n987 B.n65 32.8291
R1351 B.n981 B.n65 32.8291
R1352 B.n981 B.n980 32.8291
R1353 B.n980 B.n979 32.8291
R1354 B.n979 B.n72 32.8291
R1355 B.n973 B.n72 32.8291
R1356 B.n973 B.n972 32.8291
R1357 B.t3 B.n423 28.4842
R1358 B.n1020 B.t0 28.4842
R1359 B.n459 B.t12 24.622
R1360 B.t5 B.n988 24.622
R1361 B.n898 B.t2 22.6909
R1362 B.n1043 B.t1 22.6909
R1363 B B.n1057 18.0485
R1364 B.n797 B.n469 10.6151
R1365 B.n798 B.n797 10.6151
R1366 B.n799 B.n798 10.6151
R1367 B.n799 B.n461 10.6151
R1368 B.n809 B.n461 10.6151
R1369 B.n810 B.n809 10.6151
R1370 B.n811 B.n810 10.6151
R1371 B.n811 B.n453 10.6151
R1372 B.n821 B.n453 10.6151
R1373 B.n822 B.n821 10.6151
R1374 B.n823 B.n822 10.6151
R1375 B.n823 B.n445 10.6151
R1376 B.n833 B.n445 10.6151
R1377 B.n834 B.n833 10.6151
R1378 B.n835 B.n834 10.6151
R1379 B.n835 B.n437 10.6151
R1380 B.n845 B.n437 10.6151
R1381 B.n846 B.n845 10.6151
R1382 B.n847 B.n846 10.6151
R1383 B.n847 B.n429 10.6151
R1384 B.n857 B.n429 10.6151
R1385 B.n858 B.n857 10.6151
R1386 B.n859 B.n858 10.6151
R1387 B.n859 B.n421 10.6151
R1388 B.n869 B.n421 10.6151
R1389 B.n870 B.n869 10.6151
R1390 B.n871 B.n870 10.6151
R1391 B.n871 B.n413 10.6151
R1392 B.n881 B.n413 10.6151
R1393 B.n882 B.n881 10.6151
R1394 B.n883 B.n882 10.6151
R1395 B.n883 B.n405 10.6151
R1396 B.n894 B.n405 10.6151
R1397 B.n895 B.n894 10.6151
R1398 B.n896 B.n895 10.6151
R1399 B.n896 B.n398 10.6151
R1400 B.n907 B.n398 10.6151
R1401 B.n908 B.n907 10.6151
R1402 B.n909 B.n908 10.6151
R1403 B.n909 B.n0 10.6151
R1404 B.n785 B.n784 10.6151
R1405 B.n784 B.n783 10.6151
R1406 B.n783 B.n782 10.6151
R1407 B.n782 B.n780 10.6151
R1408 B.n780 B.n777 10.6151
R1409 B.n777 B.n776 10.6151
R1410 B.n776 B.n773 10.6151
R1411 B.n773 B.n772 10.6151
R1412 B.n772 B.n769 10.6151
R1413 B.n769 B.n768 10.6151
R1414 B.n768 B.n765 10.6151
R1415 B.n765 B.n764 10.6151
R1416 B.n764 B.n761 10.6151
R1417 B.n761 B.n760 10.6151
R1418 B.n760 B.n757 10.6151
R1419 B.n757 B.n756 10.6151
R1420 B.n756 B.n753 10.6151
R1421 B.n753 B.n752 10.6151
R1422 B.n752 B.n749 10.6151
R1423 B.n749 B.n748 10.6151
R1424 B.n748 B.n745 10.6151
R1425 B.n745 B.n744 10.6151
R1426 B.n744 B.n741 10.6151
R1427 B.n741 B.n740 10.6151
R1428 B.n740 B.n737 10.6151
R1429 B.n737 B.n736 10.6151
R1430 B.n736 B.n733 10.6151
R1431 B.n733 B.n732 10.6151
R1432 B.n732 B.n729 10.6151
R1433 B.n729 B.n728 10.6151
R1434 B.n728 B.n725 10.6151
R1435 B.n725 B.n724 10.6151
R1436 B.n724 B.n721 10.6151
R1437 B.n721 B.n720 10.6151
R1438 B.n720 B.n717 10.6151
R1439 B.n717 B.n716 10.6151
R1440 B.n716 B.n713 10.6151
R1441 B.n713 B.n712 10.6151
R1442 B.n712 B.n709 10.6151
R1443 B.n709 B.n708 10.6151
R1444 B.n708 B.n705 10.6151
R1445 B.n705 B.n704 10.6151
R1446 B.n704 B.n701 10.6151
R1447 B.n701 B.n700 10.6151
R1448 B.n700 B.n697 10.6151
R1449 B.n697 B.n696 10.6151
R1450 B.n696 B.n693 10.6151
R1451 B.n693 B.n692 10.6151
R1452 B.n692 B.n689 10.6151
R1453 B.n689 B.n688 10.6151
R1454 B.n688 B.n685 10.6151
R1455 B.n685 B.n684 10.6151
R1456 B.n684 B.n681 10.6151
R1457 B.n681 B.n680 10.6151
R1458 B.n680 B.n677 10.6151
R1459 B.n677 B.n676 10.6151
R1460 B.n676 B.n673 10.6151
R1461 B.n671 B.n668 10.6151
R1462 B.n668 B.n667 10.6151
R1463 B.n667 B.n664 10.6151
R1464 B.n664 B.n663 10.6151
R1465 B.n663 B.n660 10.6151
R1466 B.n660 B.n659 10.6151
R1467 B.n659 B.n656 10.6151
R1468 B.n656 B.n655 10.6151
R1469 B.n652 B.n651 10.6151
R1470 B.n651 B.n648 10.6151
R1471 B.n648 B.n647 10.6151
R1472 B.n647 B.n644 10.6151
R1473 B.n644 B.n643 10.6151
R1474 B.n643 B.n640 10.6151
R1475 B.n640 B.n639 10.6151
R1476 B.n639 B.n636 10.6151
R1477 B.n636 B.n635 10.6151
R1478 B.n635 B.n632 10.6151
R1479 B.n632 B.n631 10.6151
R1480 B.n631 B.n628 10.6151
R1481 B.n628 B.n627 10.6151
R1482 B.n627 B.n624 10.6151
R1483 B.n624 B.n623 10.6151
R1484 B.n623 B.n620 10.6151
R1485 B.n620 B.n619 10.6151
R1486 B.n619 B.n616 10.6151
R1487 B.n616 B.n615 10.6151
R1488 B.n615 B.n612 10.6151
R1489 B.n612 B.n611 10.6151
R1490 B.n611 B.n608 10.6151
R1491 B.n608 B.n607 10.6151
R1492 B.n607 B.n604 10.6151
R1493 B.n604 B.n603 10.6151
R1494 B.n603 B.n600 10.6151
R1495 B.n600 B.n599 10.6151
R1496 B.n599 B.n596 10.6151
R1497 B.n596 B.n595 10.6151
R1498 B.n595 B.n592 10.6151
R1499 B.n592 B.n591 10.6151
R1500 B.n591 B.n588 10.6151
R1501 B.n588 B.n587 10.6151
R1502 B.n587 B.n584 10.6151
R1503 B.n584 B.n583 10.6151
R1504 B.n583 B.n580 10.6151
R1505 B.n580 B.n579 10.6151
R1506 B.n579 B.n576 10.6151
R1507 B.n576 B.n575 10.6151
R1508 B.n575 B.n572 10.6151
R1509 B.n572 B.n571 10.6151
R1510 B.n571 B.n568 10.6151
R1511 B.n568 B.n567 10.6151
R1512 B.n567 B.n564 10.6151
R1513 B.n564 B.n563 10.6151
R1514 B.n563 B.n560 10.6151
R1515 B.n560 B.n559 10.6151
R1516 B.n559 B.n556 10.6151
R1517 B.n556 B.n555 10.6151
R1518 B.n555 B.n552 10.6151
R1519 B.n552 B.n551 10.6151
R1520 B.n551 B.n548 10.6151
R1521 B.n548 B.n547 10.6151
R1522 B.n547 B.n544 10.6151
R1523 B.n544 B.n543 10.6151
R1524 B.n543 B.n473 10.6151
R1525 B.n791 B.n473 10.6151
R1526 B.n793 B.n792 10.6151
R1527 B.n793 B.n465 10.6151
R1528 B.n803 B.n465 10.6151
R1529 B.n804 B.n803 10.6151
R1530 B.n805 B.n804 10.6151
R1531 B.n805 B.n456 10.6151
R1532 B.n815 B.n456 10.6151
R1533 B.n816 B.n815 10.6151
R1534 B.n817 B.n816 10.6151
R1535 B.n817 B.n449 10.6151
R1536 B.n827 B.n449 10.6151
R1537 B.n828 B.n827 10.6151
R1538 B.n829 B.n828 10.6151
R1539 B.n829 B.n441 10.6151
R1540 B.n839 B.n441 10.6151
R1541 B.n840 B.n839 10.6151
R1542 B.n841 B.n840 10.6151
R1543 B.n841 B.n433 10.6151
R1544 B.n851 B.n433 10.6151
R1545 B.n852 B.n851 10.6151
R1546 B.n853 B.n852 10.6151
R1547 B.n853 B.n425 10.6151
R1548 B.n863 B.n425 10.6151
R1549 B.n864 B.n863 10.6151
R1550 B.n865 B.n864 10.6151
R1551 B.n865 B.n417 10.6151
R1552 B.n875 B.n417 10.6151
R1553 B.n876 B.n875 10.6151
R1554 B.n877 B.n876 10.6151
R1555 B.n877 B.n409 10.6151
R1556 B.n887 B.n409 10.6151
R1557 B.n888 B.n887 10.6151
R1558 B.n889 B.n888 10.6151
R1559 B.n889 B.n402 10.6151
R1560 B.n900 B.n402 10.6151
R1561 B.n901 B.n900 10.6151
R1562 B.n903 B.n901 10.6151
R1563 B.n903 B.n902 10.6151
R1564 B.n902 B.n394 10.6151
R1565 B.n914 B.n394 10.6151
R1566 B.n915 B.n914 10.6151
R1567 B.n916 B.n915 10.6151
R1568 B.n917 B.n916 10.6151
R1569 B.n918 B.n917 10.6151
R1570 B.n921 B.n918 10.6151
R1571 B.n922 B.n921 10.6151
R1572 B.n923 B.n922 10.6151
R1573 B.n924 B.n923 10.6151
R1574 B.n926 B.n924 10.6151
R1575 B.n927 B.n926 10.6151
R1576 B.n928 B.n927 10.6151
R1577 B.n929 B.n928 10.6151
R1578 B.n931 B.n929 10.6151
R1579 B.n932 B.n931 10.6151
R1580 B.n933 B.n932 10.6151
R1581 B.n934 B.n933 10.6151
R1582 B.n936 B.n934 10.6151
R1583 B.n937 B.n936 10.6151
R1584 B.n938 B.n937 10.6151
R1585 B.n939 B.n938 10.6151
R1586 B.n941 B.n939 10.6151
R1587 B.n942 B.n941 10.6151
R1588 B.n943 B.n942 10.6151
R1589 B.n944 B.n943 10.6151
R1590 B.n946 B.n944 10.6151
R1591 B.n947 B.n946 10.6151
R1592 B.n948 B.n947 10.6151
R1593 B.n949 B.n948 10.6151
R1594 B.n951 B.n949 10.6151
R1595 B.n952 B.n951 10.6151
R1596 B.n953 B.n952 10.6151
R1597 B.n954 B.n953 10.6151
R1598 B.n956 B.n954 10.6151
R1599 B.n957 B.n956 10.6151
R1600 B.n958 B.n957 10.6151
R1601 B.n959 B.n958 10.6151
R1602 B.n961 B.n959 10.6151
R1603 B.n962 B.n961 10.6151
R1604 B.n963 B.n962 10.6151
R1605 B.n964 B.n963 10.6151
R1606 B.n966 B.n964 10.6151
R1607 B.n967 B.n966 10.6151
R1608 B.n968 B.n967 10.6151
R1609 B.n1049 B.n1 10.6151
R1610 B.n1049 B.n1048 10.6151
R1611 B.n1048 B.n1047 10.6151
R1612 B.n1047 B.n10 10.6151
R1613 B.n1041 B.n10 10.6151
R1614 B.n1041 B.n1040 10.6151
R1615 B.n1040 B.n1039 10.6151
R1616 B.n1039 B.n17 10.6151
R1617 B.n1033 B.n17 10.6151
R1618 B.n1033 B.n1032 10.6151
R1619 B.n1032 B.n1031 10.6151
R1620 B.n1031 B.n25 10.6151
R1621 B.n1025 B.n25 10.6151
R1622 B.n1025 B.n1024 10.6151
R1623 B.n1024 B.n1023 10.6151
R1624 B.n1023 B.n32 10.6151
R1625 B.n1017 B.n32 10.6151
R1626 B.n1017 B.n1016 10.6151
R1627 B.n1016 B.n1015 10.6151
R1628 B.n1015 B.n39 10.6151
R1629 B.n1009 B.n39 10.6151
R1630 B.n1009 B.n1008 10.6151
R1631 B.n1008 B.n1007 10.6151
R1632 B.n1007 B.n46 10.6151
R1633 B.n1001 B.n46 10.6151
R1634 B.n1001 B.n1000 10.6151
R1635 B.n1000 B.n999 10.6151
R1636 B.n999 B.n53 10.6151
R1637 B.n993 B.n53 10.6151
R1638 B.n993 B.n992 10.6151
R1639 B.n992 B.n991 10.6151
R1640 B.n991 B.n60 10.6151
R1641 B.n985 B.n60 10.6151
R1642 B.n985 B.n984 10.6151
R1643 B.n984 B.n983 10.6151
R1644 B.n983 B.n67 10.6151
R1645 B.n977 B.n67 10.6151
R1646 B.n977 B.n976 10.6151
R1647 B.n976 B.n975 10.6151
R1648 B.n975 B.n74 10.6151
R1649 B.n148 B.n147 10.6151
R1650 B.n151 B.n148 10.6151
R1651 B.n152 B.n151 10.6151
R1652 B.n155 B.n152 10.6151
R1653 B.n156 B.n155 10.6151
R1654 B.n159 B.n156 10.6151
R1655 B.n160 B.n159 10.6151
R1656 B.n163 B.n160 10.6151
R1657 B.n164 B.n163 10.6151
R1658 B.n167 B.n164 10.6151
R1659 B.n168 B.n167 10.6151
R1660 B.n171 B.n168 10.6151
R1661 B.n172 B.n171 10.6151
R1662 B.n175 B.n172 10.6151
R1663 B.n176 B.n175 10.6151
R1664 B.n179 B.n176 10.6151
R1665 B.n180 B.n179 10.6151
R1666 B.n183 B.n180 10.6151
R1667 B.n184 B.n183 10.6151
R1668 B.n187 B.n184 10.6151
R1669 B.n188 B.n187 10.6151
R1670 B.n191 B.n188 10.6151
R1671 B.n192 B.n191 10.6151
R1672 B.n195 B.n192 10.6151
R1673 B.n196 B.n195 10.6151
R1674 B.n199 B.n196 10.6151
R1675 B.n200 B.n199 10.6151
R1676 B.n203 B.n200 10.6151
R1677 B.n204 B.n203 10.6151
R1678 B.n207 B.n204 10.6151
R1679 B.n208 B.n207 10.6151
R1680 B.n211 B.n208 10.6151
R1681 B.n212 B.n211 10.6151
R1682 B.n215 B.n212 10.6151
R1683 B.n216 B.n215 10.6151
R1684 B.n219 B.n216 10.6151
R1685 B.n220 B.n219 10.6151
R1686 B.n223 B.n220 10.6151
R1687 B.n224 B.n223 10.6151
R1688 B.n227 B.n224 10.6151
R1689 B.n228 B.n227 10.6151
R1690 B.n231 B.n228 10.6151
R1691 B.n232 B.n231 10.6151
R1692 B.n235 B.n232 10.6151
R1693 B.n236 B.n235 10.6151
R1694 B.n239 B.n236 10.6151
R1695 B.n240 B.n239 10.6151
R1696 B.n243 B.n240 10.6151
R1697 B.n244 B.n243 10.6151
R1698 B.n247 B.n244 10.6151
R1699 B.n248 B.n247 10.6151
R1700 B.n251 B.n248 10.6151
R1701 B.n252 B.n251 10.6151
R1702 B.n255 B.n252 10.6151
R1703 B.n256 B.n255 10.6151
R1704 B.n259 B.n256 10.6151
R1705 B.n260 B.n259 10.6151
R1706 B.n264 B.n263 10.6151
R1707 B.n267 B.n264 10.6151
R1708 B.n268 B.n267 10.6151
R1709 B.n271 B.n268 10.6151
R1710 B.n272 B.n271 10.6151
R1711 B.n275 B.n272 10.6151
R1712 B.n276 B.n275 10.6151
R1713 B.n279 B.n276 10.6151
R1714 B.n284 B.n281 10.6151
R1715 B.n285 B.n284 10.6151
R1716 B.n288 B.n285 10.6151
R1717 B.n289 B.n288 10.6151
R1718 B.n292 B.n289 10.6151
R1719 B.n293 B.n292 10.6151
R1720 B.n296 B.n293 10.6151
R1721 B.n297 B.n296 10.6151
R1722 B.n300 B.n297 10.6151
R1723 B.n301 B.n300 10.6151
R1724 B.n304 B.n301 10.6151
R1725 B.n305 B.n304 10.6151
R1726 B.n308 B.n305 10.6151
R1727 B.n309 B.n308 10.6151
R1728 B.n312 B.n309 10.6151
R1729 B.n313 B.n312 10.6151
R1730 B.n316 B.n313 10.6151
R1731 B.n317 B.n316 10.6151
R1732 B.n320 B.n317 10.6151
R1733 B.n321 B.n320 10.6151
R1734 B.n324 B.n321 10.6151
R1735 B.n325 B.n324 10.6151
R1736 B.n328 B.n325 10.6151
R1737 B.n329 B.n328 10.6151
R1738 B.n332 B.n329 10.6151
R1739 B.n333 B.n332 10.6151
R1740 B.n336 B.n333 10.6151
R1741 B.n337 B.n336 10.6151
R1742 B.n340 B.n337 10.6151
R1743 B.n341 B.n340 10.6151
R1744 B.n344 B.n341 10.6151
R1745 B.n345 B.n344 10.6151
R1746 B.n348 B.n345 10.6151
R1747 B.n349 B.n348 10.6151
R1748 B.n352 B.n349 10.6151
R1749 B.n353 B.n352 10.6151
R1750 B.n356 B.n353 10.6151
R1751 B.n357 B.n356 10.6151
R1752 B.n360 B.n357 10.6151
R1753 B.n361 B.n360 10.6151
R1754 B.n364 B.n361 10.6151
R1755 B.n365 B.n364 10.6151
R1756 B.n368 B.n365 10.6151
R1757 B.n369 B.n368 10.6151
R1758 B.n372 B.n369 10.6151
R1759 B.n373 B.n372 10.6151
R1760 B.n376 B.n373 10.6151
R1761 B.n377 B.n376 10.6151
R1762 B.n380 B.n377 10.6151
R1763 B.n381 B.n380 10.6151
R1764 B.n384 B.n381 10.6151
R1765 B.n385 B.n384 10.6151
R1766 B.n388 B.n385 10.6151
R1767 B.n389 B.n388 10.6151
R1768 B.n392 B.n389 10.6151
R1769 B.n393 B.n392 10.6151
R1770 B.n969 B.n393 10.6151
R1771 B.n891 B.t2 10.1387
R1772 B.n19 B.t1 10.1387
R1773 B.n819 B.t12 8.20765
R1774 B.n989 B.t5 8.20765
R1775 B.n1057 B.n0 8.11757
R1776 B.n1057 B.n1 8.11757
R1777 B.n672 B.n671 6.5566
R1778 B.n655 B.n541 6.5566
R1779 B.n263 B.n145 6.5566
R1780 B.n280 B.n279 6.5566
R1781 B.n861 B.t3 4.34546
R1782 B.t0 B.n1019 4.34546
R1783 B.n673 B.n672 4.05904
R1784 B.n652 B.n541 4.05904
R1785 B.n260 B.n145 4.05904
R1786 B.n281 B.n280 4.05904
R1787 VP.n19 VP.n18 161.3
R1788 VP.n17 VP.n1 161.3
R1789 VP.n16 VP.n15 161.3
R1790 VP.n14 VP.n2 161.3
R1791 VP.n13 VP.n12 161.3
R1792 VP.n11 VP.n3 161.3
R1793 VP.n10 VP.n9 161.3
R1794 VP.n8 VP.n4 161.3
R1795 VP.n5 VP.t1 155.904
R1796 VP.n5 VP.t3 154.691
R1797 VP.n6 VP.t2 121.612
R1798 VP.n0 VP.t0 121.612
R1799 VP.n7 VP.n6 82.7273
R1800 VP.n20 VP.n0 82.7273
R1801 VP.n12 VP.n2 56.5193
R1802 VP.n7 VP.n5 55.3886
R1803 VP.n10 VP.n4 24.4675
R1804 VP.n11 VP.n10 24.4675
R1805 VP.n12 VP.n11 24.4675
R1806 VP.n16 VP.n2 24.4675
R1807 VP.n17 VP.n16 24.4675
R1808 VP.n18 VP.n17 24.4675
R1809 VP.n6 VP.n4 7.3406
R1810 VP.n18 VP.n0 7.3406
R1811 VP.n8 VP.n7 0.354971
R1812 VP.n20 VP.n19 0.354971
R1813 VP VP.n20 0.26696
R1814 VP.n9 VP.n8 0.189894
R1815 VP.n9 VP.n3 0.189894
R1816 VP.n13 VP.n3 0.189894
R1817 VP.n14 VP.n13 0.189894
R1818 VP.n15 VP.n14 0.189894
R1819 VP.n15 VP.n1 0.189894
R1820 VP.n19 VP.n1 0.189894
R1821 VTAIL.n778 VTAIL.n686 289.615
R1822 VTAIL.n92 VTAIL.n0 289.615
R1823 VTAIL.n190 VTAIL.n98 289.615
R1824 VTAIL.n288 VTAIL.n196 289.615
R1825 VTAIL.n680 VTAIL.n588 289.615
R1826 VTAIL.n582 VTAIL.n490 289.615
R1827 VTAIL.n484 VTAIL.n392 289.615
R1828 VTAIL.n386 VTAIL.n294 289.615
R1829 VTAIL.n719 VTAIL.n718 185
R1830 VTAIL.n721 VTAIL.n720 185
R1831 VTAIL.n714 VTAIL.n713 185
R1832 VTAIL.n727 VTAIL.n726 185
R1833 VTAIL.n729 VTAIL.n728 185
R1834 VTAIL.n710 VTAIL.n709 185
R1835 VTAIL.n735 VTAIL.n734 185
R1836 VTAIL.n737 VTAIL.n736 185
R1837 VTAIL.n706 VTAIL.n705 185
R1838 VTAIL.n743 VTAIL.n742 185
R1839 VTAIL.n745 VTAIL.n744 185
R1840 VTAIL.n702 VTAIL.n701 185
R1841 VTAIL.n751 VTAIL.n750 185
R1842 VTAIL.n753 VTAIL.n752 185
R1843 VTAIL.n698 VTAIL.n697 185
R1844 VTAIL.n760 VTAIL.n759 185
R1845 VTAIL.n761 VTAIL.n696 185
R1846 VTAIL.n763 VTAIL.n762 185
R1847 VTAIL.n694 VTAIL.n693 185
R1848 VTAIL.n769 VTAIL.n768 185
R1849 VTAIL.n771 VTAIL.n770 185
R1850 VTAIL.n690 VTAIL.n689 185
R1851 VTAIL.n777 VTAIL.n776 185
R1852 VTAIL.n779 VTAIL.n778 185
R1853 VTAIL.n33 VTAIL.n32 185
R1854 VTAIL.n35 VTAIL.n34 185
R1855 VTAIL.n28 VTAIL.n27 185
R1856 VTAIL.n41 VTAIL.n40 185
R1857 VTAIL.n43 VTAIL.n42 185
R1858 VTAIL.n24 VTAIL.n23 185
R1859 VTAIL.n49 VTAIL.n48 185
R1860 VTAIL.n51 VTAIL.n50 185
R1861 VTAIL.n20 VTAIL.n19 185
R1862 VTAIL.n57 VTAIL.n56 185
R1863 VTAIL.n59 VTAIL.n58 185
R1864 VTAIL.n16 VTAIL.n15 185
R1865 VTAIL.n65 VTAIL.n64 185
R1866 VTAIL.n67 VTAIL.n66 185
R1867 VTAIL.n12 VTAIL.n11 185
R1868 VTAIL.n74 VTAIL.n73 185
R1869 VTAIL.n75 VTAIL.n10 185
R1870 VTAIL.n77 VTAIL.n76 185
R1871 VTAIL.n8 VTAIL.n7 185
R1872 VTAIL.n83 VTAIL.n82 185
R1873 VTAIL.n85 VTAIL.n84 185
R1874 VTAIL.n4 VTAIL.n3 185
R1875 VTAIL.n91 VTAIL.n90 185
R1876 VTAIL.n93 VTAIL.n92 185
R1877 VTAIL.n131 VTAIL.n130 185
R1878 VTAIL.n133 VTAIL.n132 185
R1879 VTAIL.n126 VTAIL.n125 185
R1880 VTAIL.n139 VTAIL.n138 185
R1881 VTAIL.n141 VTAIL.n140 185
R1882 VTAIL.n122 VTAIL.n121 185
R1883 VTAIL.n147 VTAIL.n146 185
R1884 VTAIL.n149 VTAIL.n148 185
R1885 VTAIL.n118 VTAIL.n117 185
R1886 VTAIL.n155 VTAIL.n154 185
R1887 VTAIL.n157 VTAIL.n156 185
R1888 VTAIL.n114 VTAIL.n113 185
R1889 VTAIL.n163 VTAIL.n162 185
R1890 VTAIL.n165 VTAIL.n164 185
R1891 VTAIL.n110 VTAIL.n109 185
R1892 VTAIL.n172 VTAIL.n171 185
R1893 VTAIL.n173 VTAIL.n108 185
R1894 VTAIL.n175 VTAIL.n174 185
R1895 VTAIL.n106 VTAIL.n105 185
R1896 VTAIL.n181 VTAIL.n180 185
R1897 VTAIL.n183 VTAIL.n182 185
R1898 VTAIL.n102 VTAIL.n101 185
R1899 VTAIL.n189 VTAIL.n188 185
R1900 VTAIL.n191 VTAIL.n190 185
R1901 VTAIL.n229 VTAIL.n228 185
R1902 VTAIL.n231 VTAIL.n230 185
R1903 VTAIL.n224 VTAIL.n223 185
R1904 VTAIL.n237 VTAIL.n236 185
R1905 VTAIL.n239 VTAIL.n238 185
R1906 VTAIL.n220 VTAIL.n219 185
R1907 VTAIL.n245 VTAIL.n244 185
R1908 VTAIL.n247 VTAIL.n246 185
R1909 VTAIL.n216 VTAIL.n215 185
R1910 VTAIL.n253 VTAIL.n252 185
R1911 VTAIL.n255 VTAIL.n254 185
R1912 VTAIL.n212 VTAIL.n211 185
R1913 VTAIL.n261 VTAIL.n260 185
R1914 VTAIL.n263 VTAIL.n262 185
R1915 VTAIL.n208 VTAIL.n207 185
R1916 VTAIL.n270 VTAIL.n269 185
R1917 VTAIL.n271 VTAIL.n206 185
R1918 VTAIL.n273 VTAIL.n272 185
R1919 VTAIL.n204 VTAIL.n203 185
R1920 VTAIL.n279 VTAIL.n278 185
R1921 VTAIL.n281 VTAIL.n280 185
R1922 VTAIL.n200 VTAIL.n199 185
R1923 VTAIL.n287 VTAIL.n286 185
R1924 VTAIL.n289 VTAIL.n288 185
R1925 VTAIL.n681 VTAIL.n680 185
R1926 VTAIL.n679 VTAIL.n678 185
R1927 VTAIL.n592 VTAIL.n591 185
R1928 VTAIL.n673 VTAIL.n672 185
R1929 VTAIL.n671 VTAIL.n670 185
R1930 VTAIL.n596 VTAIL.n595 185
R1931 VTAIL.n600 VTAIL.n598 185
R1932 VTAIL.n665 VTAIL.n664 185
R1933 VTAIL.n663 VTAIL.n662 185
R1934 VTAIL.n602 VTAIL.n601 185
R1935 VTAIL.n657 VTAIL.n656 185
R1936 VTAIL.n655 VTAIL.n654 185
R1937 VTAIL.n606 VTAIL.n605 185
R1938 VTAIL.n649 VTAIL.n648 185
R1939 VTAIL.n647 VTAIL.n646 185
R1940 VTAIL.n610 VTAIL.n609 185
R1941 VTAIL.n641 VTAIL.n640 185
R1942 VTAIL.n639 VTAIL.n638 185
R1943 VTAIL.n614 VTAIL.n613 185
R1944 VTAIL.n633 VTAIL.n632 185
R1945 VTAIL.n631 VTAIL.n630 185
R1946 VTAIL.n618 VTAIL.n617 185
R1947 VTAIL.n625 VTAIL.n624 185
R1948 VTAIL.n623 VTAIL.n622 185
R1949 VTAIL.n583 VTAIL.n582 185
R1950 VTAIL.n581 VTAIL.n580 185
R1951 VTAIL.n494 VTAIL.n493 185
R1952 VTAIL.n575 VTAIL.n574 185
R1953 VTAIL.n573 VTAIL.n572 185
R1954 VTAIL.n498 VTAIL.n497 185
R1955 VTAIL.n502 VTAIL.n500 185
R1956 VTAIL.n567 VTAIL.n566 185
R1957 VTAIL.n565 VTAIL.n564 185
R1958 VTAIL.n504 VTAIL.n503 185
R1959 VTAIL.n559 VTAIL.n558 185
R1960 VTAIL.n557 VTAIL.n556 185
R1961 VTAIL.n508 VTAIL.n507 185
R1962 VTAIL.n551 VTAIL.n550 185
R1963 VTAIL.n549 VTAIL.n548 185
R1964 VTAIL.n512 VTAIL.n511 185
R1965 VTAIL.n543 VTAIL.n542 185
R1966 VTAIL.n541 VTAIL.n540 185
R1967 VTAIL.n516 VTAIL.n515 185
R1968 VTAIL.n535 VTAIL.n534 185
R1969 VTAIL.n533 VTAIL.n532 185
R1970 VTAIL.n520 VTAIL.n519 185
R1971 VTAIL.n527 VTAIL.n526 185
R1972 VTAIL.n525 VTAIL.n524 185
R1973 VTAIL.n485 VTAIL.n484 185
R1974 VTAIL.n483 VTAIL.n482 185
R1975 VTAIL.n396 VTAIL.n395 185
R1976 VTAIL.n477 VTAIL.n476 185
R1977 VTAIL.n475 VTAIL.n474 185
R1978 VTAIL.n400 VTAIL.n399 185
R1979 VTAIL.n404 VTAIL.n402 185
R1980 VTAIL.n469 VTAIL.n468 185
R1981 VTAIL.n467 VTAIL.n466 185
R1982 VTAIL.n406 VTAIL.n405 185
R1983 VTAIL.n461 VTAIL.n460 185
R1984 VTAIL.n459 VTAIL.n458 185
R1985 VTAIL.n410 VTAIL.n409 185
R1986 VTAIL.n453 VTAIL.n452 185
R1987 VTAIL.n451 VTAIL.n450 185
R1988 VTAIL.n414 VTAIL.n413 185
R1989 VTAIL.n445 VTAIL.n444 185
R1990 VTAIL.n443 VTAIL.n442 185
R1991 VTAIL.n418 VTAIL.n417 185
R1992 VTAIL.n437 VTAIL.n436 185
R1993 VTAIL.n435 VTAIL.n434 185
R1994 VTAIL.n422 VTAIL.n421 185
R1995 VTAIL.n429 VTAIL.n428 185
R1996 VTAIL.n427 VTAIL.n426 185
R1997 VTAIL.n387 VTAIL.n386 185
R1998 VTAIL.n385 VTAIL.n384 185
R1999 VTAIL.n298 VTAIL.n297 185
R2000 VTAIL.n379 VTAIL.n378 185
R2001 VTAIL.n377 VTAIL.n376 185
R2002 VTAIL.n302 VTAIL.n301 185
R2003 VTAIL.n306 VTAIL.n304 185
R2004 VTAIL.n371 VTAIL.n370 185
R2005 VTAIL.n369 VTAIL.n368 185
R2006 VTAIL.n308 VTAIL.n307 185
R2007 VTAIL.n363 VTAIL.n362 185
R2008 VTAIL.n361 VTAIL.n360 185
R2009 VTAIL.n312 VTAIL.n311 185
R2010 VTAIL.n355 VTAIL.n354 185
R2011 VTAIL.n353 VTAIL.n352 185
R2012 VTAIL.n316 VTAIL.n315 185
R2013 VTAIL.n347 VTAIL.n346 185
R2014 VTAIL.n345 VTAIL.n344 185
R2015 VTAIL.n320 VTAIL.n319 185
R2016 VTAIL.n339 VTAIL.n338 185
R2017 VTAIL.n337 VTAIL.n336 185
R2018 VTAIL.n324 VTAIL.n323 185
R2019 VTAIL.n331 VTAIL.n330 185
R2020 VTAIL.n329 VTAIL.n328 185
R2021 VTAIL.n717 VTAIL.t0 147.659
R2022 VTAIL.n31 VTAIL.t1 147.659
R2023 VTAIL.n129 VTAIL.t7 147.659
R2024 VTAIL.n227 VTAIL.t5 147.659
R2025 VTAIL.n621 VTAIL.t4 147.659
R2026 VTAIL.n523 VTAIL.t6 147.659
R2027 VTAIL.n425 VTAIL.t2 147.659
R2028 VTAIL.n327 VTAIL.t3 147.659
R2029 VTAIL.n720 VTAIL.n719 104.615
R2030 VTAIL.n720 VTAIL.n713 104.615
R2031 VTAIL.n727 VTAIL.n713 104.615
R2032 VTAIL.n728 VTAIL.n727 104.615
R2033 VTAIL.n728 VTAIL.n709 104.615
R2034 VTAIL.n735 VTAIL.n709 104.615
R2035 VTAIL.n736 VTAIL.n735 104.615
R2036 VTAIL.n736 VTAIL.n705 104.615
R2037 VTAIL.n743 VTAIL.n705 104.615
R2038 VTAIL.n744 VTAIL.n743 104.615
R2039 VTAIL.n744 VTAIL.n701 104.615
R2040 VTAIL.n751 VTAIL.n701 104.615
R2041 VTAIL.n752 VTAIL.n751 104.615
R2042 VTAIL.n752 VTAIL.n697 104.615
R2043 VTAIL.n760 VTAIL.n697 104.615
R2044 VTAIL.n761 VTAIL.n760 104.615
R2045 VTAIL.n762 VTAIL.n761 104.615
R2046 VTAIL.n762 VTAIL.n693 104.615
R2047 VTAIL.n769 VTAIL.n693 104.615
R2048 VTAIL.n770 VTAIL.n769 104.615
R2049 VTAIL.n770 VTAIL.n689 104.615
R2050 VTAIL.n777 VTAIL.n689 104.615
R2051 VTAIL.n778 VTAIL.n777 104.615
R2052 VTAIL.n34 VTAIL.n33 104.615
R2053 VTAIL.n34 VTAIL.n27 104.615
R2054 VTAIL.n41 VTAIL.n27 104.615
R2055 VTAIL.n42 VTAIL.n41 104.615
R2056 VTAIL.n42 VTAIL.n23 104.615
R2057 VTAIL.n49 VTAIL.n23 104.615
R2058 VTAIL.n50 VTAIL.n49 104.615
R2059 VTAIL.n50 VTAIL.n19 104.615
R2060 VTAIL.n57 VTAIL.n19 104.615
R2061 VTAIL.n58 VTAIL.n57 104.615
R2062 VTAIL.n58 VTAIL.n15 104.615
R2063 VTAIL.n65 VTAIL.n15 104.615
R2064 VTAIL.n66 VTAIL.n65 104.615
R2065 VTAIL.n66 VTAIL.n11 104.615
R2066 VTAIL.n74 VTAIL.n11 104.615
R2067 VTAIL.n75 VTAIL.n74 104.615
R2068 VTAIL.n76 VTAIL.n75 104.615
R2069 VTAIL.n76 VTAIL.n7 104.615
R2070 VTAIL.n83 VTAIL.n7 104.615
R2071 VTAIL.n84 VTAIL.n83 104.615
R2072 VTAIL.n84 VTAIL.n3 104.615
R2073 VTAIL.n91 VTAIL.n3 104.615
R2074 VTAIL.n92 VTAIL.n91 104.615
R2075 VTAIL.n132 VTAIL.n131 104.615
R2076 VTAIL.n132 VTAIL.n125 104.615
R2077 VTAIL.n139 VTAIL.n125 104.615
R2078 VTAIL.n140 VTAIL.n139 104.615
R2079 VTAIL.n140 VTAIL.n121 104.615
R2080 VTAIL.n147 VTAIL.n121 104.615
R2081 VTAIL.n148 VTAIL.n147 104.615
R2082 VTAIL.n148 VTAIL.n117 104.615
R2083 VTAIL.n155 VTAIL.n117 104.615
R2084 VTAIL.n156 VTAIL.n155 104.615
R2085 VTAIL.n156 VTAIL.n113 104.615
R2086 VTAIL.n163 VTAIL.n113 104.615
R2087 VTAIL.n164 VTAIL.n163 104.615
R2088 VTAIL.n164 VTAIL.n109 104.615
R2089 VTAIL.n172 VTAIL.n109 104.615
R2090 VTAIL.n173 VTAIL.n172 104.615
R2091 VTAIL.n174 VTAIL.n173 104.615
R2092 VTAIL.n174 VTAIL.n105 104.615
R2093 VTAIL.n181 VTAIL.n105 104.615
R2094 VTAIL.n182 VTAIL.n181 104.615
R2095 VTAIL.n182 VTAIL.n101 104.615
R2096 VTAIL.n189 VTAIL.n101 104.615
R2097 VTAIL.n190 VTAIL.n189 104.615
R2098 VTAIL.n230 VTAIL.n229 104.615
R2099 VTAIL.n230 VTAIL.n223 104.615
R2100 VTAIL.n237 VTAIL.n223 104.615
R2101 VTAIL.n238 VTAIL.n237 104.615
R2102 VTAIL.n238 VTAIL.n219 104.615
R2103 VTAIL.n245 VTAIL.n219 104.615
R2104 VTAIL.n246 VTAIL.n245 104.615
R2105 VTAIL.n246 VTAIL.n215 104.615
R2106 VTAIL.n253 VTAIL.n215 104.615
R2107 VTAIL.n254 VTAIL.n253 104.615
R2108 VTAIL.n254 VTAIL.n211 104.615
R2109 VTAIL.n261 VTAIL.n211 104.615
R2110 VTAIL.n262 VTAIL.n261 104.615
R2111 VTAIL.n262 VTAIL.n207 104.615
R2112 VTAIL.n270 VTAIL.n207 104.615
R2113 VTAIL.n271 VTAIL.n270 104.615
R2114 VTAIL.n272 VTAIL.n271 104.615
R2115 VTAIL.n272 VTAIL.n203 104.615
R2116 VTAIL.n279 VTAIL.n203 104.615
R2117 VTAIL.n280 VTAIL.n279 104.615
R2118 VTAIL.n280 VTAIL.n199 104.615
R2119 VTAIL.n287 VTAIL.n199 104.615
R2120 VTAIL.n288 VTAIL.n287 104.615
R2121 VTAIL.n680 VTAIL.n679 104.615
R2122 VTAIL.n679 VTAIL.n591 104.615
R2123 VTAIL.n672 VTAIL.n591 104.615
R2124 VTAIL.n672 VTAIL.n671 104.615
R2125 VTAIL.n671 VTAIL.n595 104.615
R2126 VTAIL.n600 VTAIL.n595 104.615
R2127 VTAIL.n664 VTAIL.n600 104.615
R2128 VTAIL.n664 VTAIL.n663 104.615
R2129 VTAIL.n663 VTAIL.n601 104.615
R2130 VTAIL.n656 VTAIL.n601 104.615
R2131 VTAIL.n656 VTAIL.n655 104.615
R2132 VTAIL.n655 VTAIL.n605 104.615
R2133 VTAIL.n648 VTAIL.n605 104.615
R2134 VTAIL.n648 VTAIL.n647 104.615
R2135 VTAIL.n647 VTAIL.n609 104.615
R2136 VTAIL.n640 VTAIL.n609 104.615
R2137 VTAIL.n640 VTAIL.n639 104.615
R2138 VTAIL.n639 VTAIL.n613 104.615
R2139 VTAIL.n632 VTAIL.n613 104.615
R2140 VTAIL.n632 VTAIL.n631 104.615
R2141 VTAIL.n631 VTAIL.n617 104.615
R2142 VTAIL.n624 VTAIL.n617 104.615
R2143 VTAIL.n624 VTAIL.n623 104.615
R2144 VTAIL.n582 VTAIL.n581 104.615
R2145 VTAIL.n581 VTAIL.n493 104.615
R2146 VTAIL.n574 VTAIL.n493 104.615
R2147 VTAIL.n574 VTAIL.n573 104.615
R2148 VTAIL.n573 VTAIL.n497 104.615
R2149 VTAIL.n502 VTAIL.n497 104.615
R2150 VTAIL.n566 VTAIL.n502 104.615
R2151 VTAIL.n566 VTAIL.n565 104.615
R2152 VTAIL.n565 VTAIL.n503 104.615
R2153 VTAIL.n558 VTAIL.n503 104.615
R2154 VTAIL.n558 VTAIL.n557 104.615
R2155 VTAIL.n557 VTAIL.n507 104.615
R2156 VTAIL.n550 VTAIL.n507 104.615
R2157 VTAIL.n550 VTAIL.n549 104.615
R2158 VTAIL.n549 VTAIL.n511 104.615
R2159 VTAIL.n542 VTAIL.n511 104.615
R2160 VTAIL.n542 VTAIL.n541 104.615
R2161 VTAIL.n541 VTAIL.n515 104.615
R2162 VTAIL.n534 VTAIL.n515 104.615
R2163 VTAIL.n534 VTAIL.n533 104.615
R2164 VTAIL.n533 VTAIL.n519 104.615
R2165 VTAIL.n526 VTAIL.n519 104.615
R2166 VTAIL.n526 VTAIL.n525 104.615
R2167 VTAIL.n484 VTAIL.n483 104.615
R2168 VTAIL.n483 VTAIL.n395 104.615
R2169 VTAIL.n476 VTAIL.n395 104.615
R2170 VTAIL.n476 VTAIL.n475 104.615
R2171 VTAIL.n475 VTAIL.n399 104.615
R2172 VTAIL.n404 VTAIL.n399 104.615
R2173 VTAIL.n468 VTAIL.n404 104.615
R2174 VTAIL.n468 VTAIL.n467 104.615
R2175 VTAIL.n467 VTAIL.n405 104.615
R2176 VTAIL.n460 VTAIL.n405 104.615
R2177 VTAIL.n460 VTAIL.n459 104.615
R2178 VTAIL.n459 VTAIL.n409 104.615
R2179 VTAIL.n452 VTAIL.n409 104.615
R2180 VTAIL.n452 VTAIL.n451 104.615
R2181 VTAIL.n451 VTAIL.n413 104.615
R2182 VTAIL.n444 VTAIL.n413 104.615
R2183 VTAIL.n444 VTAIL.n443 104.615
R2184 VTAIL.n443 VTAIL.n417 104.615
R2185 VTAIL.n436 VTAIL.n417 104.615
R2186 VTAIL.n436 VTAIL.n435 104.615
R2187 VTAIL.n435 VTAIL.n421 104.615
R2188 VTAIL.n428 VTAIL.n421 104.615
R2189 VTAIL.n428 VTAIL.n427 104.615
R2190 VTAIL.n386 VTAIL.n385 104.615
R2191 VTAIL.n385 VTAIL.n297 104.615
R2192 VTAIL.n378 VTAIL.n297 104.615
R2193 VTAIL.n378 VTAIL.n377 104.615
R2194 VTAIL.n377 VTAIL.n301 104.615
R2195 VTAIL.n306 VTAIL.n301 104.615
R2196 VTAIL.n370 VTAIL.n306 104.615
R2197 VTAIL.n370 VTAIL.n369 104.615
R2198 VTAIL.n369 VTAIL.n307 104.615
R2199 VTAIL.n362 VTAIL.n307 104.615
R2200 VTAIL.n362 VTAIL.n361 104.615
R2201 VTAIL.n361 VTAIL.n311 104.615
R2202 VTAIL.n354 VTAIL.n311 104.615
R2203 VTAIL.n354 VTAIL.n353 104.615
R2204 VTAIL.n353 VTAIL.n315 104.615
R2205 VTAIL.n346 VTAIL.n315 104.615
R2206 VTAIL.n346 VTAIL.n345 104.615
R2207 VTAIL.n345 VTAIL.n319 104.615
R2208 VTAIL.n338 VTAIL.n319 104.615
R2209 VTAIL.n338 VTAIL.n337 104.615
R2210 VTAIL.n337 VTAIL.n323 104.615
R2211 VTAIL.n330 VTAIL.n323 104.615
R2212 VTAIL.n330 VTAIL.n329 104.615
R2213 VTAIL.n719 VTAIL.t0 52.3082
R2214 VTAIL.n33 VTAIL.t1 52.3082
R2215 VTAIL.n131 VTAIL.t7 52.3082
R2216 VTAIL.n229 VTAIL.t5 52.3082
R2217 VTAIL.n623 VTAIL.t4 52.3082
R2218 VTAIL.n525 VTAIL.t6 52.3082
R2219 VTAIL.n427 VTAIL.t2 52.3082
R2220 VTAIL.n329 VTAIL.t3 52.3082
R2221 VTAIL.n783 VTAIL.n782 31.9914
R2222 VTAIL.n97 VTAIL.n96 31.9914
R2223 VTAIL.n195 VTAIL.n194 31.9914
R2224 VTAIL.n293 VTAIL.n292 31.9914
R2225 VTAIL.n685 VTAIL.n684 31.9914
R2226 VTAIL.n587 VTAIL.n586 31.9914
R2227 VTAIL.n489 VTAIL.n488 31.9914
R2228 VTAIL.n391 VTAIL.n390 31.9914
R2229 VTAIL.n783 VTAIL.n685 30.7376
R2230 VTAIL.n391 VTAIL.n293 30.7376
R2231 VTAIL.n718 VTAIL.n717 15.6677
R2232 VTAIL.n32 VTAIL.n31 15.6677
R2233 VTAIL.n130 VTAIL.n129 15.6677
R2234 VTAIL.n228 VTAIL.n227 15.6677
R2235 VTAIL.n622 VTAIL.n621 15.6677
R2236 VTAIL.n524 VTAIL.n523 15.6677
R2237 VTAIL.n426 VTAIL.n425 15.6677
R2238 VTAIL.n328 VTAIL.n327 15.6677
R2239 VTAIL.n763 VTAIL.n694 13.1884
R2240 VTAIL.n77 VTAIL.n8 13.1884
R2241 VTAIL.n175 VTAIL.n106 13.1884
R2242 VTAIL.n273 VTAIL.n204 13.1884
R2243 VTAIL.n598 VTAIL.n596 13.1884
R2244 VTAIL.n500 VTAIL.n498 13.1884
R2245 VTAIL.n402 VTAIL.n400 13.1884
R2246 VTAIL.n304 VTAIL.n302 13.1884
R2247 VTAIL.n721 VTAIL.n716 12.8005
R2248 VTAIL.n764 VTAIL.n696 12.8005
R2249 VTAIL.n768 VTAIL.n767 12.8005
R2250 VTAIL.n35 VTAIL.n30 12.8005
R2251 VTAIL.n78 VTAIL.n10 12.8005
R2252 VTAIL.n82 VTAIL.n81 12.8005
R2253 VTAIL.n133 VTAIL.n128 12.8005
R2254 VTAIL.n176 VTAIL.n108 12.8005
R2255 VTAIL.n180 VTAIL.n179 12.8005
R2256 VTAIL.n231 VTAIL.n226 12.8005
R2257 VTAIL.n274 VTAIL.n206 12.8005
R2258 VTAIL.n278 VTAIL.n277 12.8005
R2259 VTAIL.n670 VTAIL.n669 12.8005
R2260 VTAIL.n666 VTAIL.n665 12.8005
R2261 VTAIL.n625 VTAIL.n620 12.8005
R2262 VTAIL.n572 VTAIL.n571 12.8005
R2263 VTAIL.n568 VTAIL.n567 12.8005
R2264 VTAIL.n527 VTAIL.n522 12.8005
R2265 VTAIL.n474 VTAIL.n473 12.8005
R2266 VTAIL.n470 VTAIL.n469 12.8005
R2267 VTAIL.n429 VTAIL.n424 12.8005
R2268 VTAIL.n376 VTAIL.n375 12.8005
R2269 VTAIL.n372 VTAIL.n371 12.8005
R2270 VTAIL.n331 VTAIL.n326 12.8005
R2271 VTAIL.n722 VTAIL.n714 12.0247
R2272 VTAIL.n759 VTAIL.n758 12.0247
R2273 VTAIL.n771 VTAIL.n692 12.0247
R2274 VTAIL.n36 VTAIL.n28 12.0247
R2275 VTAIL.n73 VTAIL.n72 12.0247
R2276 VTAIL.n85 VTAIL.n6 12.0247
R2277 VTAIL.n134 VTAIL.n126 12.0247
R2278 VTAIL.n171 VTAIL.n170 12.0247
R2279 VTAIL.n183 VTAIL.n104 12.0247
R2280 VTAIL.n232 VTAIL.n224 12.0247
R2281 VTAIL.n269 VTAIL.n268 12.0247
R2282 VTAIL.n281 VTAIL.n202 12.0247
R2283 VTAIL.n673 VTAIL.n594 12.0247
R2284 VTAIL.n662 VTAIL.n599 12.0247
R2285 VTAIL.n626 VTAIL.n618 12.0247
R2286 VTAIL.n575 VTAIL.n496 12.0247
R2287 VTAIL.n564 VTAIL.n501 12.0247
R2288 VTAIL.n528 VTAIL.n520 12.0247
R2289 VTAIL.n477 VTAIL.n398 12.0247
R2290 VTAIL.n466 VTAIL.n403 12.0247
R2291 VTAIL.n430 VTAIL.n422 12.0247
R2292 VTAIL.n379 VTAIL.n300 12.0247
R2293 VTAIL.n368 VTAIL.n305 12.0247
R2294 VTAIL.n332 VTAIL.n324 12.0247
R2295 VTAIL.n726 VTAIL.n725 11.249
R2296 VTAIL.n757 VTAIL.n698 11.249
R2297 VTAIL.n772 VTAIL.n690 11.249
R2298 VTAIL.n40 VTAIL.n39 11.249
R2299 VTAIL.n71 VTAIL.n12 11.249
R2300 VTAIL.n86 VTAIL.n4 11.249
R2301 VTAIL.n138 VTAIL.n137 11.249
R2302 VTAIL.n169 VTAIL.n110 11.249
R2303 VTAIL.n184 VTAIL.n102 11.249
R2304 VTAIL.n236 VTAIL.n235 11.249
R2305 VTAIL.n267 VTAIL.n208 11.249
R2306 VTAIL.n282 VTAIL.n200 11.249
R2307 VTAIL.n674 VTAIL.n592 11.249
R2308 VTAIL.n661 VTAIL.n602 11.249
R2309 VTAIL.n630 VTAIL.n629 11.249
R2310 VTAIL.n576 VTAIL.n494 11.249
R2311 VTAIL.n563 VTAIL.n504 11.249
R2312 VTAIL.n532 VTAIL.n531 11.249
R2313 VTAIL.n478 VTAIL.n396 11.249
R2314 VTAIL.n465 VTAIL.n406 11.249
R2315 VTAIL.n434 VTAIL.n433 11.249
R2316 VTAIL.n380 VTAIL.n298 11.249
R2317 VTAIL.n367 VTAIL.n308 11.249
R2318 VTAIL.n336 VTAIL.n335 11.249
R2319 VTAIL.n729 VTAIL.n712 10.4732
R2320 VTAIL.n754 VTAIL.n753 10.4732
R2321 VTAIL.n776 VTAIL.n775 10.4732
R2322 VTAIL.n43 VTAIL.n26 10.4732
R2323 VTAIL.n68 VTAIL.n67 10.4732
R2324 VTAIL.n90 VTAIL.n89 10.4732
R2325 VTAIL.n141 VTAIL.n124 10.4732
R2326 VTAIL.n166 VTAIL.n165 10.4732
R2327 VTAIL.n188 VTAIL.n187 10.4732
R2328 VTAIL.n239 VTAIL.n222 10.4732
R2329 VTAIL.n264 VTAIL.n263 10.4732
R2330 VTAIL.n286 VTAIL.n285 10.4732
R2331 VTAIL.n678 VTAIL.n677 10.4732
R2332 VTAIL.n658 VTAIL.n657 10.4732
R2333 VTAIL.n633 VTAIL.n616 10.4732
R2334 VTAIL.n580 VTAIL.n579 10.4732
R2335 VTAIL.n560 VTAIL.n559 10.4732
R2336 VTAIL.n535 VTAIL.n518 10.4732
R2337 VTAIL.n482 VTAIL.n481 10.4732
R2338 VTAIL.n462 VTAIL.n461 10.4732
R2339 VTAIL.n437 VTAIL.n420 10.4732
R2340 VTAIL.n384 VTAIL.n383 10.4732
R2341 VTAIL.n364 VTAIL.n363 10.4732
R2342 VTAIL.n339 VTAIL.n322 10.4732
R2343 VTAIL.n730 VTAIL.n710 9.69747
R2344 VTAIL.n750 VTAIL.n700 9.69747
R2345 VTAIL.n779 VTAIL.n688 9.69747
R2346 VTAIL.n44 VTAIL.n24 9.69747
R2347 VTAIL.n64 VTAIL.n14 9.69747
R2348 VTAIL.n93 VTAIL.n2 9.69747
R2349 VTAIL.n142 VTAIL.n122 9.69747
R2350 VTAIL.n162 VTAIL.n112 9.69747
R2351 VTAIL.n191 VTAIL.n100 9.69747
R2352 VTAIL.n240 VTAIL.n220 9.69747
R2353 VTAIL.n260 VTAIL.n210 9.69747
R2354 VTAIL.n289 VTAIL.n198 9.69747
R2355 VTAIL.n681 VTAIL.n590 9.69747
R2356 VTAIL.n654 VTAIL.n604 9.69747
R2357 VTAIL.n634 VTAIL.n614 9.69747
R2358 VTAIL.n583 VTAIL.n492 9.69747
R2359 VTAIL.n556 VTAIL.n506 9.69747
R2360 VTAIL.n536 VTAIL.n516 9.69747
R2361 VTAIL.n485 VTAIL.n394 9.69747
R2362 VTAIL.n458 VTAIL.n408 9.69747
R2363 VTAIL.n438 VTAIL.n418 9.69747
R2364 VTAIL.n387 VTAIL.n296 9.69747
R2365 VTAIL.n360 VTAIL.n310 9.69747
R2366 VTAIL.n340 VTAIL.n320 9.69747
R2367 VTAIL.n782 VTAIL.n781 9.45567
R2368 VTAIL.n96 VTAIL.n95 9.45567
R2369 VTAIL.n194 VTAIL.n193 9.45567
R2370 VTAIL.n292 VTAIL.n291 9.45567
R2371 VTAIL.n684 VTAIL.n683 9.45567
R2372 VTAIL.n586 VTAIL.n585 9.45567
R2373 VTAIL.n488 VTAIL.n487 9.45567
R2374 VTAIL.n390 VTAIL.n389 9.45567
R2375 VTAIL.n781 VTAIL.n780 9.3005
R2376 VTAIL.n688 VTAIL.n687 9.3005
R2377 VTAIL.n775 VTAIL.n774 9.3005
R2378 VTAIL.n773 VTAIL.n772 9.3005
R2379 VTAIL.n692 VTAIL.n691 9.3005
R2380 VTAIL.n767 VTAIL.n766 9.3005
R2381 VTAIL.n739 VTAIL.n738 9.3005
R2382 VTAIL.n708 VTAIL.n707 9.3005
R2383 VTAIL.n733 VTAIL.n732 9.3005
R2384 VTAIL.n731 VTAIL.n730 9.3005
R2385 VTAIL.n712 VTAIL.n711 9.3005
R2386 VTAIL.n725 VTAIL.n724 9.3005
R2387 VTAIL.n723 VTAIL.n722 9.3005
R2388 VTAIL.n716 VTAIL.n715 9.3005
R2389 VTAIL.n741 VTAIL.n740 9.3005
R2390 VTAIL.n704 VTAIL.n703 9.3005
R2391 VTAIL.n747 VTAIL.n746 9.3005
R2392 VTAIL.n749 VTAIL.n748 9.3005
R2393 VTAIL.n700 VTAIL.n699 9.3005
R2394 VTAIL.n755 VTAIL.n754 9.3005
R2395 VTAIL.n757 VTAIL.n756 9.3005
R2396 VTAIL.n758 VTAIL.n695 9.3005
R2397 VTAIL.n765 VTAIL.n764 9.3005
R2398 VTAIL.n95 VTAIL.n94 9.3005
R2399 VTAIL.n2 VTAIL.n1 9.3005
R2400 VTAIL.n89 VTAIL.n88 9.3005
R2401 VTAIL.n87 VTAIL.n86 9.3005
R2402 VTAIL.n6 VTAIL.n5 9.3005
R2403 VTAIL.n81 VTAIL.n80 9.3005
R2404 VTAIL.n53 VTAIL.n52 9.3005
R2405 VTAIL.n22 VTAIL.n21 9.3005
R2406 VTAIL.n47 VTAIL.n46 9.3005
R2407 VTAIL.n45 VTAIL.n44 9.3005
R2408 VTAIL.n26 VTAIL.n25 9.3005
R2409 VTAIL.n39 VTAIL.n38 9.3005
R2410 VTAIL.n37 VTAIL.n36 9.3005
R2411 VTAIL.n30 VTAIL.n29 9.3005
R2412 VTAIL.n55 VTAIL.n54 9.3005
R2413 VTAIL.n18 VTAIL.n17 9.3005
R2414 VTAIL.n61 VTAIL.n60 9.3005
R2415 VTAIL.n63 VTAIL.n62 9.3005
R2416 VTAIL.n14 VTAIL.n13 9.3005
R2417 VTAIL.n69 VTAIL.n68 9.3005
R2418 VTAIL.n71 VTAIL.n70 9.3005
R2419 VTAIL.n72 VTAIL.n9 9.3005
R2420 VTAIL.n79 VTAIL.n78 9.3005
R2421 VTAIL.n193 VTAIL.n192 9.3005
R2422 VTAIL.n100 VTAIL.n99 9.3005
R2423 VTAIL.n187 VTAIL.n186 9.3005
R2424 VTAIL.n185 VTAIL.n184 9.3005
R2425 VTAIL.n104 VTAIL.n103 9.3005
R2426 VTAIL.n179 VTAIL.n178 9.3005
R2427 VTAIL.n151 VTAIL.n150 9.3005
R2428 VTAIL.n120 VTAIL.n119 9.3005
R2429 VTAIL.n145 VTAIL.n144 9.3005
R2430 VTAIL.n143 VTAIL.n142 9.3005
R2431 VTAIL.n124 VTAIL.n123 9.3005
R2432 VTAIL.n137 VTAIL.n136 9.3005
R2433 VTAIL.n135 VTAIL.n134 9.3005
R2434 VTAIL.n128 VTAIL.n127 9.3005
R2435 VTAIL.n153 VTAIL.n152 9.3005
R2436 VTAIL.n116 VTAIL.n115 9.3005
R2437 VTAIL.n159 VTAIL.n158 9.3005
R2438 VTAIL.n161 VTAIL.n160 9.3005
R2439 VTAIL.n112 VTAIL.n111 9.3005
R2440 VTAIL.n167 VTAIL.n166 9.3005
R2441 VTAIL.n169 VTAIL.n168 9.3005
R2442 VTAIL.n170 VTAIL.n107 9.3005
R2443 VTAIL.n177 VTAIL.n176 9.3005
R2444 VTAIL.n291 VTAIL.n290 9.3005
R2445 VTAIL.n198 VTAIL.n197 9.3005
R2446 VTAIL.n285 VTAIL.n284 9.3005
R2447 VTAIL.n283 VTAIL.n282 9.3005
R2448 VTAIL.n202 VTAIL.n201 9.3005
R2449 VTAIL.n277 VTAIL.n276 9.3005
R2450 VTAIL.n249 VTAIL.n248 9.3005
R2451 VTAIL.n218 VTAIL.n217 9.3005
R2452 VTAIL.n243 VTAIL.n242 9.3005
R2453 VTAIL.n241 VTAIL.n240 9.3005
R2454 VTAIL.n222 VTAIL.n221 9.3005
R2455 VTAIL.n235 VTAIL.n234 9.3005
R2456 VTAIL.n233 VTAIL.n232 9.3005
R2457 VTAIL.n226 VTAIL.n225 9.3005
R2458 VTAIL.n251 VTAIL.n250 9.3005
R2459 VTAIL.n214 VTAIL.n213 9.3005
R2460 VTAIL.n257 VTAIL.n256 9.3005
R2461 VTAIL.n259 VTAIL.n258 9.3005
R2462 VTAIL.n210 VTAIL.n209 9.3005
R2463 VTAIL.n265 VTAIL.n264 9.3005
R2464 VTAIL.n267 VTAIL.n266 9.3005
R2465 VTAIL.n268 VTAIL.n205 9.3005
R2466 VTAIL.n275 VTAIL.n274 9.3005
R2467 VTAIL.n608 VTAIL.n607 9.3005
R2468 VTAIL.n651 VTAIL.n650 9.3005
R2469 VTAIL.n653 VTAIL.n652 9.3005
R2470 VTAIL.n604 VTAIL.n603 9.3005
R2471 VTAIL.n659 VTAIL.n658 9.3005
R2472 VTAIL.n661 VTAIL.n660 9.3005
R2473 VTAIL.n599 VTAIL.n597 9.3005
R2474 VTAIL.n667 VTAIL.n666 9.3005
R2475 VTAIL.n683 VTAIL.n682 9.3005
R2476 VTAIL.n590 VTAIL.n589 9.3005
R2477 VTAIL.n677 VTAIL.n676 9.3005
R2478 VTAIL.n675 VTAIL.n674 9.3005
R2479 VTAIL.n594 VTAIL.n593 9.3005
R2480 VTAIL.n669 VTAIL.n668 9.3005
R2481 VTAIL.n645 VTAIL.n644 9.3005
R2482 VTAIL.n643 VTAIL.n642 9.3005
R2483 VTAIL.n612 VTAIL.n611 9.3005
R2484 VTAIL.n637 VTAIL.n636 9.3005
R2485 VTAIL.n635 VTAIL.n634 9.3005
R2486 VTAIL.n616 VTAIL.n615 9.3005
R2487 VTAIL.n629 VTAIL.n628 9.3005
R2488 VTAIL.n627 VTAIL.n626 9.3005
R2489 VTAIL.n620 VTAIL.n619 9.3005
R2490 VTAIL.n510 VTAIL.n509 9.3005
R2491 VTAIL.n553 VTAIL.n552 9.3005
R2492 VTAIL.n555 VTAIL.n554 9.3005
R2493 VTAIL.n506 VTAIL.n505 9.3005
R2494 VTAIL.n561 VTAIL.n560 9.3005
R2495 VTAIL.n563 VTAIL.n562 9.3005
R2496 VTAIL.n501 VTAIL.n499 9.3005
R2497 VTAIL.n569 VTAIL.n568 9.3005
R2498 VTAIL.n585 VTAIL.n584 9.3005
R2499 VTAIL.n492 VTAIL.n491 9.3005
R2500 VTAIL.n579 VTAIL.n578 9.3005
R2501 VTAIL.n577 VTAIL.n576 9.3005
R2502 VTAIL.n496 VTAIL.n495 9.3005
R2503 VTAIL.n571 VTAIL.n570 9.3005
R2504 VTAIL.n547 VTAIL.n546 9.3005
R2505 VTAIL.n545 VTAIL.n544 9.3005
R2506 VTAIL.n514 VTAIL.n513 9.3005
R2507 VTAIL.n539 VTAIL.n538 9.3005
R2508 VTAIL.n537 VTAIL.n536 9.3005
R2509 VTAIL.n518 VTAIL.n517 9.3005
R2510 VTAIL.n531 VTAIL.n530 9.3005
R2511 VTAIL.n529 VTAIL.n528 9.3005
R2512 VTAIL.n522 VTAIL.n521 9.3005
R2513 VTAIL.n412 VTAIL.n411 9.3005
R2514 VTAIL.n455 VTAIL.n454 9.3005
R2515 VTAIL.n457 VTAIL.n456 9.3005
R2516 VTAIL.n408 VTAIL.n407 9.3005
R2517 VTAIL.n463 VTAIL.n462 9.3005
R2518 VTAIL.n465 VTAIL.n464 9.3005
R2519 VTAIL.n403 VTAIL.n401 9.3005
R2520 VTAIL.n471 VTAIL.n470 9.3005
R2521 VTAIL.n487 VTAIL.n486 9.3005
R2522 VTAIL.n394 VTAIL.n393 9.3005
R2523 VTAIL.n481 VTAIL.n480 9.3005
R2524 VTAIL.n479 VTAIL.n478 9.3005
R2525 VTAIL.n398 VTAIL.n397 9.3005
R2526 VTAIL.n473 VTAIL.n472 9.3005
R2527 VTAIL.n449 VTAIL.n448 9.3005
R2528 VTAIL.n447 VTAIL.n446 9.3005
R2529 VTAIL.n416 VTAIL.n415 9.3005
R2530 VTAIL.n441 VTAIL.n440 9.3005
R2531 VTAIL.n439 VTAIL.n438 9.3005
R2532 VTAIL.n420 VTAIL.n419 9.3005
R2533 VTAIL.n433 VTAIL.n432 9.3005
R2534 VTAIL.n431 VTAIL.n430 9.3005
R2535 VTAIL.n424 VTAIL.n423 9.3005
R2536 VTAIL.n314 VTAIL.n313 9.3005
R2537 VTAIL.n357 VTAIL.n356 9.3005
R2538 VTAIL.n359 VTAIL.n358 9.3005
R2539 VTAIL.n310 VTAIL.n309 9.3005
R2540 VTAIL.n365 VTAIL.n364 9.3005
R2541 VTAIL.n367 VTAIL.n366 9.3005
R2542 VTAIL.n305 VTAIL.n303 9.3005
R2543 VTAIL.n373 VTAIL.n372 9.3005
R2544 VTAIL.n389 VTAIL.n388 9.3005
R2545 VTAIL.n296 VTAIL.n295 9.3005
R2546 VTAIL.n383 VTAIL.n382 9.3005
R2547 VTAIL.n381 VTAIL.n380 9.3005
R2548 VTAIL.n300 VTAIL.n299 9.3005
R2549 VTAIL.n375 VTAIL.n374 9.3005
R2550 VTAIL.n351 VTAIL.n350 9.3005
R2551 VTAIL.n349 VTAIL.n348 9.3005
R2552 VTAIL.n318 VTAIL.n317 9.3005
R2553 VTAIL.n343 VTAIL.n342 9.3005
R2554 VTAIL.n341 VTAIL.n340 9.3005
R2555 VTAIL.n322 VTAIL.n321 9.3005
R2556 VTAIL.n335 VTAIL.n334 9.3005
R2557 VTAIL.n333 VTAIL.n332 9.3005
R2558 VTAIL.n326 VTAIL.n325 9.3005
R2559 VTAIL.n734 VTAIL.n733 8.92171
R2560 VTAIL.n749 VTAIL.n702 8.92171
R2561 VTAIL.n780 VTAIL.n686 8.92171
R2562 VTAIL.n48 VTAIL.n47 8.92171
R2563 VTAIL.n63 VTAIL.n16 8.92171
R2564 VTAIL.n94 VTAIL.n0 8.92171
R2565 VTAIL.n146 VTAIL.n145 8.92171
R2566 VTAIL.n161 VTAIL.n114 8.92171
R2567 VTAIL.n192 VTAIL.n98 8.92171
R2568 VTAIL.n244 VTAIL.n243 8.92171
R2569 VTAIL.n259 VTAIL.n212 8.92171
R2570 VTAIL.n290 VTAIL.n196 8.92171
R2571 VTAIL.n682 VTAIL.n588 8.92171
R2572 VTAIL.n653 VTAIL.n606 8.92171
R2573 VTAIL.n638 VTAIL.n637 8.92171
R2574 VTAIL.n584 VTAIL.n490 8.92171
R2575 VTAIL.n555 VTAIL.n508 8.92171
R2576 VTAIL.n540 VTAIL.n539 8.92171
R2577 VTAIL.n486 VTAIL.n392 8.92171
R2578 VTAIL.n457 VTAIL.n410 8.92171
R2579 VTAIL.n442 VTAIL.n441 8.92171
R2580 VTAIL.n388 VTAIL.n294 8.92171
R2581 VTAIL.n359 VTAIL.n312 8.92171
R2582 VTAIL.n344 VTAIL.n343 8.92171
R2583 VTAIL.n737 VTAIL.n708 8.14595
R2584 VTAIL.n746 VTAIL.n745 8.14595
R2585 VTAIL.n51 VTAIL.n22 8.14595
R2586 VTAIL.n60 VTAIL.n59 8.14595
R2587 VTAIL.n149 VTAIL.n120 8.14595
R2588 VTAIL.n158 VTAIL.n157 8.14595
R2589 VTAIL.n247 VTAIL.n218 8.14595
R2590 VTAIL.n256 VTAIL.n255 8.14595
R2591 VTAIL.n650 VTAIL.n649 8.14595
R2592 VTAIL.n641 VTAIL.n612 8.14595
R2593 VTAIL.n552 VTAIL.n551 8.14595
R2594 VTAIL.n543 VTAIL.n514 8.14595
R2595 VTAIL.n454 VTAIL.n453 8.14595
R2596 VTAIL.n445 VTAIL.n416 8.14595
R2597 VTAIL.n356 VTAIL.n355 8.14595
R2598 VTAIL.n347 VTAIL.n318 8.14595
R2599 VTAIL.n738 VTAIL.n706 7.3702
R2600 VTAIL.n742 VTAIL.n704 7.3702
R2601 VTAIL.n52 VTAIL.n20 7.3702
R2602 VTAIL.n56 VTAIL.n18 7.3702
R2603 VTAIL.n150 VTAIL.n118 7.3702
R2604 VTAIL.n154 VTAIL.n116 7.3702
R2605 VTAIL.n248 VTAIL.n216 7.3702
R2606 VTAIL.n252 VTAIL.n214 7.3702
R2607 VTAIL.n646 VTAIL.n608 7.3702
R2608 VTAIL.n642 VTAIL.n610 7.3702
R2609 VTAIL.n548 VTAIL.n510 7.3702
R2610 VTAIL.n544 VTAIL.n512 7.3702
R2611 VTAIL.n450 VTAIL.n412 7.3702
R2612 VTAIL.n446 VTAIL.n414 7.3702
R2613 VTAIL.n352 VTAIL.n314 7.3702
R2614 VTAIL.n348 VTAIL.n316 7.3702
R2615 VTAIL.n741 VTAIL.n706 6.59444
R2616 VTAIL.n742 VTAIL.n741 6.59444
R2617 VTAIL.n55 VTAIL.n20 6.59444
R2618 VTAIL.n56 VTAIL.n55 6.59444
R2619 VTAIL.n153 VTAIL.n118 6.59444
R2620 VTAIL.n154 VTAIL.n153 6.59444
R2621 VTAIL.n251 VTAIL.n216 6.59444
R2622 VTAIL.n252 VTAIL.n251 6.59444
R2623 VTAIL.n646 VTAIL.n645 6.59444
R2624 VTAIL.n645 VTAIL.n610 6.59444
R2625 VTAIL.n548 VTAIL.n547 6.59444
R2626 VTAIL.n547 VTAIL.n512 6.59444
R2627 VTAIL.n450 VTAIL.n449 6.59444
R2628 VTAIL.n449 VTAIL.n414 6.59444
R2629 VTAIL.n352 VTAIL.n351 6.59444
R2630 VTAIL.n351 VTAIL.n316 6.59444
R2631 VTAIL.n738 VTAIL.n737 5.81868
R2632 VTAIL.n745 VTAIL.n704 5.81868
R2633 VTAIL.n52 VTAIL.n51 5.81868
R2634 VTAIL.n59 VTAIL.n18 5.81868
R2635 VTAIL.n150 VTAIL.n149 5.81868
R2636 VTAIL.n157 VTAIL.n116 5.81868
R2637 VTAIL.n248 VTAIL.n247 5.81868
R2638 VTAIL.n255 VTAIL.n214 5.81868
R2639 VTAIL.n649 VTAIL.n608 5.81868
R2640 VTAIL.n642 VTAIL.n641 5.81868
R2641 VTAIL.n551 VTAIL.n510 5.81868
R2642 VTAIL.n544 VTAIL.n543 5.81868
R2643 VTAIL.n453 VTAIL.n412 5.81868
R2644 VTAIL.n446 VTAIL.n445 5.81868
R2645 VTAIL.n355 VTAIL.n314 5.81868
R2646 VTAIL.n348 VTAIL.n347 5.81868
R2647 VTAIL.n734 VTAIL.n708 5.04292
R2648 VTAIL.n746 VTAIL.n702 5.04292
R2649 VTAIL.n782 VTAIL.n686 5.04292
R2650 VTAIL.n48 VTAIL.n22 5.04292
R2651 VTAIL.n60 VTAIL.n16 5.04292
R2652 VTAIL.n96 VTAIL.n0 5.04292
R2653 VTAIL.n146 VTAIL.n120 5.04292
R2654 VTAIL.n158 VTAIL.n114 5.04292
R2655 VTAIL.n194 VTAIL.n98 5.04292
R2656 VTAIL.n244 VTAIL.n218 5.04292
R2657 VTAIL.n256 VTAIL.n212 5.04292
R2658 VTAIL.n292 VTAIL.n196 5.04292
R2659 VTAIL.n684 VTAIL.n588 5.04292
R2660 VTAIL.n650 VTAIL.n606 5.04292
R2661 VTAIL.n638 VTAIL.n612 5.04292
R2662 VTAIL.n586 VTAIL.n490 5.04292
R2663 VTAIL.n552 VTAIL.n508 5.04292
R2664 VTAIL.n540 VTAIL.n514 5.04292
R2665 VTAIL.n488 VTAIL.n392 5.04292
R2666 VTAIL.n454 VTAIL.n410 5.04292
R2667 VTAIL.n442 VTAIL.n416 5.04292
R2668 VTAIL.n390 VTAIL.n294 5.04292
R2669 VTAIL.n356 VTAIL.n312 5.04292
R2670 VTAIL.n344 VTAIL.n318 5.04292
R2671 VTAIL.n717 VTAIL.n715 4.38563
R2672 VTAIL.n31 VTAIL.n29 4.38563
R2673 VTAIL.n129 VTAIL.n127 4.38563
R2674 VTAIL.n227 VTAIL.n225 4.38563
R2675 VTAIL.n621 VTAIL.n619 4.38563
R2676 VTAIL.n523 VTAIL.n521 4.38563
R2677 VTAIL.n425 VTAIL.n423 4.38563
R2678 VTAIL.n327 VTAIL.n325 4.38563
R2679 VTAIL.n733 VTAIL.n710 4.26717
R2680 VTAIL.n750 VTAIL.n749 4.26717
R2681 VTAIL.n780 VTAIL.n779 4.26717
R2682 VTAIL.n47 VTAIL.n24 4.26717
R2683 VTAIL.n64 VTAIL.n63 4.26717
R2684 VTAIL.n94 VTAIL.n93 4.26717
R2685 VTAIL.n145 VTAIL.n122 4.26717
R2686 VTAIL.n162 VTAIL.n161 4.26717
R2687 VTAIL.n192 VTAIL.n191 4.26717
R2688 VTAIL.n243 VTAIL.n220 4.26717
R2689 VTAIL.n260 VTAIL.n259 4.26717
R2690 VTAIL.n290 VTAIL.n289 4.26717
R2691 VTAIL.n682 VTAIL.n681 4.26717
R2692 VTAIL.n654 VTAIL.n653 4.26717
R2693 VTAIL.n637 VTAIL.n614 4.26717
R2694 VTAIL.n584 VTAIL.n583 4.26717
R2695 VTAIL.n556 VTAIL.n555 4.26717
R2696 VTAIL.n539 VTAIL.n516 4.26717
R2697 VTAIL.n486 VTAIL.n485 4.26717
R2698 VTAIL.n458 VTAIL.n457 4.26717
R2699 VTAIL.n441 VTAIL.n418 4.26717
R2700 VTAIL.n388 VTAIL.n387 4.26717
R2701 VTAIL.n360 VTAIL.n359 4.26717
R2702 VTAIL.n343 VTAIL.n320 4.26717
R2703 VTAIL.n730 VTAIL.n729 3.49141
R2704 VTAIL.n753 VTAIL.n700 3.49141
R2705 VTAIL.n776 VTAIL.n688 3.49141
R2706 VTAIL.n44 VTAIL.n43 3.49141
R2707 VTAIL.n67 VTAIL.n14 3.49141
R2708 VTAIL.n90 VTAIL.n2 3.49141
R2709 VTAIL.n142 VTAIL.n141 3.49141
R2710 VTAIL.n165 VTAIL.n112 3.49141
R2711 VTAIL.n188 VTAIL.n100 3.49141
R2712 VTAIL.n240 VTAIL.n239 3.49141
R2713 VTAIL.n263 VTAIL.n210 3.49141
R2714 VTAIL.n286 VTAIL.n198 3.49141
R2715 VTAIL.n678 VTAIL.n590 3.49141
R2716 VTAIL.n657 VTAIL.n604 3.49141
R2717 VTAIL.n634 VTAIL.n633 3.49141
R2718 VTAIL.n580 VTAIL.n492 3.49141
R2719 VTAIL.n559 VTAIL.n506 3.49141
R2720 VTAIL.n536 VTAIL.n535 3.49141
R2721 VTAIL.n482 VTAIL.n394 3.49141
R2722 VTAIL.n461 VTAIL.n408 3.49141
R2723 VTAIL.n438 VTAIL.n437 3.49141
R2724 VTAIL.n384 VTAIL.n296 3.49141
R2725 VTAIL.n363 VTAIL.n310 3.49141
R2726 VTAIL.n340 VTAIL.n339 3.49141
R2727 VTAIL.n489 VTAIL.n391 3.27636
R2728 VTAIL.n685 VTAIL.n587 3.27636
R2729 VTAIL.n293 VTAIL.n195 3.27636
R2730 VTAIL.n726 VTAIL.n712 2.71565
R2731 VTAIL.n754 VTAIL.n698 2.71565
R2732 VTAIL.n775 VTAIL.n690 2.71565
R2733 VTAIL.n40 VTAIL.n26 2.71565
R2734 VTAIL.n68 VTAIL.n12 2.71565
R2735 VTAIL.n89 VTAIL.n4 2.71565
R2736 VTAIL.n138 VTAIL.n124 2.71565
R2737 VTAIL.n166 VTAIL.n110 2.71565
R2738 VTAIL.n187 VTAIL.n102 2.71565
R2739 VTAIL.n236 VTAIL.n222 2.71565
R2740 VTAIL.n264 VTAIL.n208 2.71565
R2741 VTAIL.n285 VTAIL.n200 2.71565
R2742 VTAIL.n677 VTAIL.n592 2.71565
R2743 VTAIL.n658 VTAIL.n602 2.71565
R2744 VTAIL.n630 VTAIL.n616 2.71565
R2745 VTAIL.n579 VTAIL.n494 2.71565
R2746 VTAIL.n560 VTAIL.n504 2.71565
R2747 VTAIL.n532 VTAIL.n518 2.71565
R2748 VTAIL.n481 VTAIL.n396 2.71565
R2749 VTAIL.n462 VTAIL.n406 2.71565
R2750 VTAIL.n434 VTAIL.n420 2.71565
R2751 VTAIL.n383 VTAIL.n298 2.71565
R2752 VTAIL.n364 VTAIL.n308 2.71565
R2753 VTAIL.n336 VTAIL.n322 2.71565
R2754 VTAIL.n725 VTAIL.n714 1.93989
R2755 VTAIL.n759 VTAIL.n757 1.93989
R2756 VTAIL.n772 VTAIL.n771 1.93989
R2757 VTAIL.n39 VTAIL.n28 1.93989
R2758 VTAIL.n73 VTAIL.n71 1.93989
R2759 VTAIL.n86 VTAIL.n85 1.93989
R2760 VTAIL.n137 VTAIL.n126 1.93989
R2761 VTAIL.n171 VTAIL.n169 1.93989
R2762 VTAIL.n184 VTAIL.n183 1.93989
R2763 VTAIL.n235 VTAIL.n224 1.93989
R2764 VTAIL.n269 VTAIL.n267 1.93989
R2765 VTAIL.n282 VTAIL.n281 1.93989
R2766 VTAIL.n674 VTAIL.n673 1.93989
R2767 VTAIL.n662 VTAIL.n661 1.93989
R2768 VTAIL.n629 VTAIL.n618 1.93989
R2769 VTAIL.n576 VTAIL.n575 1.93989
R2770 VTAIL.n564 VTAIL.n563 1.93989
R2771 VTAIL.n531 VTAIL.n520 1.93989
R2772 VTAIL.n478 VTAIL.n477 1.93989
R2773 VTAIL.n466 VTAIL.n465 1.93989
R2774 VTAIL.n433 VTAIL.n422 1.93989
R2775 VTAIL.n380 VTAIL.n379 1.93989
R2776 VTAIL.n368 VTAIL.n367 1.93989
R2777 VTAIL.n335 VTAIL.n324 1.93989
R2778 VTAIL VTAIL.n97 1.69662
R2779 VTAIL VTAIL.n783 1.58024
R2780 VTAIL.n722 VTAIL.n721 1.16414
R2781 VTAIL.n758 VTAIL.n696 1.16414
R2782 VTAIL.n768 VTAIL.n692 1.16414
R2783 VTAIL.n36 VTAIL.n35 1.16414
R2784 VTAIL.n72 VTAIL.n10 1.16414
R2785 VTAIL.n82 VTAIL.n6 1.16414
R2786 VTAIL.n134 VTAIL.n133 1.16414
R2787 VTAIL.n170 VTAIL.n108 1.16414
R2788 VTAIL.n180 VTAIL.n104 1.16414
R2789 VTAIL.n232 VTAIL.n231 1.16414
R2790 VTAIL.n268 VTAIL.n206 1.16414
R2791 VTAIL.n278 VTAIL.n202 1.16414
R2792 VTAIL.n670 VTAIL.n594 1.16414
R2793 VTAIL.n665 VTAIL.n599 1.16414
R2794 VTAIL.n626 VTAIL.n625 1.16414
R2795 VTAIL.n572 VTAIL.n496 1.16414
R2796 VTAIL.n567 VTAIL.n501 1.16414
R2797 VTAIL.n528 VTAIL.n527 1.16414
R2798 VTAIL.n474 VTAIL.n398 1.16414
R2799 VTAIL.n469 VTAIL.n403 1.16414
R2800 VTAIL.n430 VTAIL.n429 1.16414
R2801 VTAIL.n376 VTAIL.n300 1.16414
R2802 VTAIL.n371 VTAIL.n305 1.16414
R2803 VTAIL.n332 VTAIL.n331 1.16414
R2804 VTAIL.n587 VTAIL.n489 0.470328
R2805 VTAIL.n195 VTAIL.n97 0.470328
R2806 VTAIL.n718 VTAIL.n716 0.388379
R2807 VTAIL.n764 VTAIL.n763 0.388379
R2808 VTAIL.n767 VTAIL.n694 0.388379
R2809 VTAIL.n32 VTAIL.n30 0.388379
R2810 VTAIL.n78 VTAIL.n77 0.388379
R2811 VTAIL.n81 VTAIL.n8 0.388379
R2812 VTAIL.n130 VTAIL.n128 0.388379
R2813 VTAIL.n176 VTAIL.n175 0.388379
R2814 VTAIL.n179 VTAIL.n106 0.388379
R2815 VTAIL.n228 VTAIL.n226 0.388379
R2816 VTAIL.n274 VTAIL.n273 0.388379
R2817 VTAIL.n277 VTAIL.n204 0.388379
R2818 VTAIL.n669 VTAIL.n596 0.388379
R2819 VTAIL.n666 VTAIL.n598 0.388379
R2820 VTAIL.n622 VTAIL.n620 0.388379
R2821 VTAIL.n571 VTAIL.n498 0.388379
R2822 VTAIL.n568 VTAIL.n500 0.388379
R2823 VTAIL.n524 VTAIL.n522 0.388379
R2824 VTAIL.n473 VTAIL.n400 0.388379
R2825 VTAIL.n470 VTAIL.n402 0.388379
R2826 VTAIL.n426 VTAIL.n424 0.388379
R2827 VTAIL.n375 VTAIL.n302 0.388379
R2828 VTAIL.n372 VTAIL.n304 0.388379
R2829 VTAIL.n328 VTAIL.n326 0.388379
R2830 VTAIL.n723 VTAIL.n715 0.155672
R2831 VTAIL.n724 VTAIL.n723 0.155672
R2832 VTAIL.n724 VTAIL.n711 0.155672
R2833 VTAIL.n731 VTAIL.n711 0.155672
R2834 VTAIL.n732 VTAIL.n731 0.155672
R2835 VTAIL.n732 VTAIL.n707 0.155672
R2836 VTAIL.n739 VTAIL.n707 0.155672
R2837 VTAIL.n740 VTAIL.n739 0.155672
R2838 VTAIL.n740 VTAIL.n703 0.155672
R2839 VTAIL.n747 VTAIL.n703 0.155672
R2840 VTAIL.n748 VTAIL.n747 0.155672
R2841 VTAIL.n748 VTAIL.n699 0.155672
R2842 VTAIL.n755 VTAIL.n699 0.155672
R2843 VTAIL.n756 VTAIL.n755 0.155672
R2844 VTAIL.n756 VTAIL.n695 0.155672
R2845 VTAIL.n765 VTAIL.n695 0.155672
R2846 VTAIL.n766 VTAIL.n765 0.155672
R2847 VTAIL.n766 VTAIL.n691 0.155672
R2848 VTAIL.n773 VTAIL.n691 0.155672
R2849 VTAIL.n774 VTAIL.n773 0.155672
R2850 VTAIL.n774 VTAIL.n687 0.155672
R2851 VTAIL.n781 VTAIL.n687 0.155672
R2852 VTAIL.n37 VTAIL.n29 0.155672
R2853 VTAIL.n38 VTAIL.n37 0.155672
R2854 VTAIL.n38 VTAIL.n25 0.155672
R2855 VTAIL.n45 VTAIL.n25 0.155672
R2856 VTAIL.n46 VTAIL.n45 0.155672
R2857 VTAIL.n46 VTAIL.n21 0.155672
R2858 VTAIL.n53 VTAIL.n21 0.155672
R2859 VTAIL.n54 VTAIL.n53 0.155672
R2860 VTAIL.n54 VTAIL.n17 0.155672
R2861 VTAIL.n61 VTAIL.n17 0.155672
R2862 VTAIL.n62 VTAIL.n61 0.155672
R2863 VTAIL.n62 VTAIL.n13 0.155672
R2864 VTAIL.n69 VTAIL.n13 0.155672
R2865 VTAIL.n70 VTAIL.n69 0.155672
R2866 VTAIL.n70 VTAIL.n9 0.155672
R2867 VTAIL.n79 VTAIL.n9 0.155672
R2868 VTAIL.n80 VTAIL.n79 0.155672
R2869 VTAIL.n80 VTAIL.n5 0.155672
R2870 VTAIL.n87 VTAIL.n5 0.155672
R2871 VTAIL.n88 VTAIL.n87 0.155672
R2872 VTAIL.n88 VTAIL.n1 0.155672
R2873 VTAIL.n95 VTAIL.n1 0.155672
R2874 VTAIL.n135 VTAIL.n127 0.155672
R2875 VTAIL.n136 VTAIL.n135 0.155672
R2876 VTAIL.n136 VTAIL.n123 0.155672
R2877 VTAIL.n143 VTAIL.n123 0.155672
R2878 VTAIL.n144 VTAIL.n143 0.155672
R2879 VTAIL.n144 VTAIL.n119 0.155672
R2880 VTAIL.n151 VTAIL.n119 0.155672
R2881 VTAIL.n152 VTAIL.n151 0.155672
R2882 VTAIL.n152 VTAIL.n115 0.155672
R2883 VTAIL.n159 VTAIL.n115 0.155672
R2884 VTAIL.n160 VTAIL.n159 0.155672
R2885 VTAIL.n160 VTAIL.n111 0.155672
R2886 VTAIL.n167 VTAIL.n111 0.155672
R2887 VTAIL.n168 VTAIL.n167 0.155672
R2888 VTAIL.n168 VTAIL.n107 0.155672
R2889 VTAIL.n177 VTAIL.n107 0.155672
R2890 VTAIL.n178 VTAIL.n177 0.155672
R2891 VTAIL.n178 VTAIL.n103 0.155672
R2892 VTAIL.n185 VTAIL.n103 0.155672
R2893 VTAIL.n186 VTAIL.n185 0.155672
R2894 VTAIL.n186 VTAIL.n99 0.155672
R2895 VTAIL.n193 VTAIL.n99 0.155672
R2896 VTAIL.n233 VTAIL.n225 0.155672
R2897 VTAIL.n234 VTAIL.n233 0.155672
R2898 VTAIL.n234 VTAIL.n221 0.155672
R2899 VTAIL.n241 VTAIL.n221 0.155672
R2900 VTAIL.n242 VTAIL.n241 0.155672
R2901 VTAIL.n242 VTAIL.n217 0.155672
R2902 VTAIL.n249 VTAIL.n217 0.155672
R2903 VTAIL.n250 VTAIL.n249 0.155672
R2904 VTAIL.n250 VTAIL.n213 0.155672
R2905 VTAIL.n257 VTAIL.n213 0.155672
R2906 VTAIL.n258 VTAIL.n257 0.155672
R2907 VTAIL.n258 VTAIL.n209 0.155672
R2908 VTAIL.n265 VTAIL.n209 0.155672
R2909 VTAIL.n266 VTAIL.n265 0.155672
R2910 VTAIL.n266 VTAIL.n205 0.155672
R2911 VTAIL.n275 VTAIL.n205 0.155672
R2912 VTAIL.n276 VTAIL.n275 0.155672
R2913 VTAIL.n276 VTAIL.n201 0.155672
R2914 VTAIL.n283 VTAIL.n201 0.155672
R2915 VTAIL.n284 VTAIL.n283 0.155672
R2916 VTAIL.n284 VTAIL.n197 0.155672
R2917 VTAIL.n291 VTAIL.n197 0.155672
R2918 VTAIL.n683 VTAIL.n589 0.155672
R2919 VTAIL.n676 VTAIL.n589 0.155672
R2920 VTAIL.n676 VTAIL.n675 0.155672
R2921 VTAIL.n675 VTAIL.n593 0.155672
R2922 VTAIL.n668 VTAIL.n593 0.155672
R2923 VTAIL.n668 VTAIL.n667 0.155672
R2924 VTAIL.n667 VTAIL.n597 0.155672
R2925 VTAIL.n660 VTAIL.n597 0.155672
R2926 VTAIL.n660 VTAIL.n659 0.155672
R2927 VTAIL.n659 VTAIL.n603 0.155672
R2928 VTAIL.n652 VTAIL.n603 0.155672
R2929 VTAIL.n652 VTAIL.n651 0.155672
R2930 VTAIL.n651 VTAIL.n607 0.155672
R2931 VTAIL.n644 VTAIL.n607 0.155672
R2932 VTAIL.n644 VTAIL.n643 0.155672
R2933 VTAIL.n643 VTAIL.n611 0.155672
R2934 VTAIL.n636 VTAIL.n611 0.155672
R2935 VTAIL.n636 VTAIL.n635 0.155672
R2936 VTAIL.n635 VTAIL.n615 0.155672
R2937 VTAIL.n628 VTAIL.n615 0.155672
R2938 VTAIL.n628 VTAIL.n627 0.155672
R2939 VTAIL.n627 VTAIL.n619 0.155672
R2940 VTAIL.n585 VTAIL.n491 0.155672
R2941 VTAIL.n578 VTAIL.n491 0.155672
R2942 VTAIL.n578 VTAIL.n577 0.155672
R2943 VTAIL.n577 VTAIL.n495 0.155672
R2944 VTAIL.n570 VTAIL.n495 0.155672
R2945 VTAIL.n570 VTAIL.n569 0.155672
R2946 VTAIL.n569 VTAIL.n499 0.155672
R2947 VTAIL.n562 VTAIL.n499 0.155672
R2948 VTAIL.n562 VTAIL.n561 0.155672
R2949 VTAIL.n561 VTAIL.n505 0.155672
R2950 VTAIL.n554 VTAIL.n505 0.155672
R2951 VTAIL.n554 VTAIL.n553 0.155672
R2952 VTAIL.n553 VTAIL.n509 0.155672
R2953 VTAIL.n546 VTAIL.n509 0.155672
R2954 VTAIL.n546 VTAIL.n545 0.155672
R2955 VTAIL.n545 VTAIL.n513 0.155672
R2956 VTAIL.n538 VTAIL.n513 0.155672
R2957 VTAIL.n538 VTAIL.n537 0.155672
R2958 VTAIL.n537 VTAIL.n517 0.155672
R2959 VTAIL.n530 VTAIL.n517 0.155672
R2960 VTAIL.n530 VTAIL.n529 0.155672
R2961 VTAIL.n529 VTAIL.n521 0.155672
R2962 VTAIL.n487 VTAIL.n393 0.155672
R2963 VTAIL.n480 VTAIL.n393 0.155672
R2964 VTAIL.n480 VTAIL.n479 0.155672
R2965 VTAIL.n479 VTAIL.n397 0.155672
R2966 VTAIL.n472 VTAIL.n397 0.155672
R2967 VTAIL.n472 VTAIL.n471 0.155672
R2968 VTAIL.n471 VTAIL.n401 0.155672
R2969 VTAIL.n464 VTAIL.n401 0.155672
R2970 VTAIL.n464 VTAIL.n463 0.155672
R2971 VTAIL.n463 VTAIL.n407 0.155672
R2972 VTAIL.n456 VTAIL.n407 0.155672
R2973 VTAIL.n456 VTAIL.n455 0.155672
R2974 VTAIL.n455 VTAIL.n411 0.155672
R2975 VTAIL.n448 VTAIL.n411 0.155672
R2976 VTAIL.n448 VTAIL.n447 0.155672
R2977 VTAIL.n447 VTAIL.n415 0.155672
R2978 VTAIL.n440 VTAIL.n415 0.155672
R2979 VTAIL.n440 VTAIL.n439 0.155672
R2980 VTAIL.n439 VTAIL.n419 0.155672
R2981 VTAIL.n432 VTAIL.n419 0.155672
R2982 VTAIL.n432 VTAIL.n431 0.155672
R2983 VTAIL.n431 VTAIL.n423 0.155672
R2984 VTAIL.n389 VTAIL.n295 0.155672
R2985 VTAIL.n382 VTAIL.n295 0.155672
R2986 VTAIL.n382 VTAIL.n381 0.155672
R2987 VTAIL.n381 VTAIL.n299 0.155672
R2988 VTAIL.n374 VTAIL.n299 0.155672
R2989 VTAIL.n374 VTAIL.n373 0.155672
R2990 VTAIL.n373 VTAIL.n303 0.155672
R2991 VTAIL.n366 VTAIL.n303 0.155672
R2992 VTAIL.n366 VTAIL.n365 0.155672
R2993 VTAIL.n365 VTAIL.n309 0.155672
R2994 VTAIL.n358 VTAIL.n309 0.155672
R2995 VTAIL.n358 VTAIL.n357 0.155672
R2996 VTAIL.n357 VTAIL.n313 0.155672
R2997 VTAIL.n350 VTAIL.n313 0.155672
R2998 VTAIL.n350 VTAIL.n349 0.155672
R2999 VTAIL.n349 VTAIL.n317 0.155672
R3000 VTAIL.n342 VTAIL.n317 0.155672
R3001 VTAIL.n342 VTAIL.n341 0.155672
R3002 VTAIL.n341 VTAIL.n321 0.155672
R3003 VTAIL.n334 VTAIL.n321 0.155672
R3004 VTAIL.n334 VTAIL.n333 0.155672
R3005 VTAIL.n333 VTAIL.n325 0.155672
R3006 VDD1 VDD1.n1 109.65
R3007 VDD1 VDD1.n0 60.5462
R3008 VDD1.n0 VDD1.t2 1.13128
R3009 VDD1.n0 VDD1.t0 1.13128
R3010 VDD1.n1 VDD1.t1 1.13128
R3011 VDD1.n1 VDD1.t3 1.13128
R3012 VN.n1 VN.t1 155.905
R3013 VN.n0 VN.t3 155.905
R3014 VN.n0 VN.t2 154.691
R3015 VN.n1 VN.t0 154.691
R3016 VN VN.n1 55.554
R3017 VN VN.n0 2.23199
R3018 VDD2.n2 VDD2.n0 109.126
R3019 VDD2.n2 VDD2.n1 60.488
R3020 VDD2.n1 VDD2.t3 1.13128
R3021 VDD2.n1 VDD2.t2 1.13128
R3022 VDD2.n0 VDD2.t0 1.13128
R3023 VDD2.n0 VDD2.t1 1.13128
R3024 VDD2 VDD2.n2 0.0586897
C0 VDD1 VN 0.149936f
C1 VP VTAIL 6.90155f
C2 VDD1 VTAIL 6.81161f
C3 VDD2 VN 7.10309f
C4 VDD2 VTAIL 6.87165f
C5 VDD1 VP 7.40201f
C6 VDD2 VP 0.449815f
C7 VDD1 VDD2 1.23376f
C8 VN VTAIL 6.88745f
C9 VP VN 7.841331f
C10 VDD2 B 4.695212f
C11 VDD1 B 9.68151f
C12 VTAIL B 13.901127f
C13 VN B 12.809911f
C14 VP B 11.164065f
C15 VDD2.t0 B 0.370063f
C16 VDD2.t1 B 0.370063f
C17 VDD2.n0 B 4.30392f
C18 VDD2.t3 B 0.370063f
C19 VDD2.t2 B 0.370063f
C20 VDD2.n1 B 3.36699f
C21 VDD2.n2 B 4.56078f
C22 VN.t2 B 3.60316f
C23 VN.t3 B 3.61293f
C24 VN.n0 B 2.22023f
C25 VN.t1 B 3.61293f
C26 VN.t0 B 3.60316f
C27 VN.n1 B 3.61867f
C28 VDD1.t2 B 0.37272f
C29 VDD1.t0 B 0.37272f
C30 VDD1.n0 B 3.39167f
C31 VDD1.t1 B 0.37272f
C32 VDD1.t3 B 0.37272f
C33 VDD1.n1 B 4.36404f
C34 VTAIL.n0 B 0.021604f
C35 VTAIL.n1 B 0.015748f
C36 VTAIL.n2 B 0.008462f
C37 VTAIL.n3 B 0.020001f
C38 VTAIL.n4 B 0.00896f
C39 VTAIL.n5 B 0.015748f
C40 VTAIL.n6 B 0.008462f
C41 VTAIL.n7 B 0.020001f
C42 VTAIL.n8 B 0.008711f
C43 VTAIL.n9 B 0.015748f
C44 VTAIL.n10 B 0.00896f
C45 VTAIL.n11 B 0.020001f
C46 VTAIL.n12 B 0.00896f
C47 VTAIL.n13 B 0.015748f
C48 VTAIL.n14 B 0.008462f
C49 VTAIL.n15 B 0.020001f
C50 VTAIL.n16 B 0.00896f
C51 VTAIL.n17 B 0.015748f
C52 VTAIL.n18 B 0.008462f
C53 VTAIL.n19 B 0.020001f
C54 VTAIL.n20 B 0.00896f
C55 VTAIL.n21 B 0.015748f
C56 VTAIL.n22 B 0.008462f
C57 VTAIL.n23 B 0.020001f
C58 VTAIL.n24 B 0.00896f
C59 VTAIL.n25 B 0.015748f
C60 VTAIL.n26 B 0.008462f
C61 VTAIL.n27 B 0.020001f
C62 VTAIL.n28 B 0.00896f
C63 VTAIL.n29 B 1.20573f
C64 VTAIL.n30 B 0.008462f
C65 VTAIL.t1 B 0.033116f
C66 VTAIL.n31 B 0.112621f
C67 VTAIL.n32 B 0.011816f
C68 VTAIL.n33 B 0.015001f
C69 VTAIL.n34 B 0.020001f
C70 VTAIL.n35 B 0.00896f
C71 VTAIL.n36 B 0.008462f
C72 VTAIL.n37 B 0.015748f
C73 VTAIL.n38 B 0.015748f
C74 VTAIL.n39 B 0.008462f
C75 VTAIL.n40 B 0.00896f
C76 VTAIL.n41 B 0.020001f
C77 VTAIL.n42 B 0.020001f
C78 VTAIL.n43 B 0.00896f
C79 VTAIL.n44 B 0.008462f
C80 VTAIL.n45 B 0.015748f
C81 VTAIL.n46 B 0.015748f
C82 VTAIL.n47 B 0.008462f
C83 VTAIL.n48 B 0.00896f
C84 VTAIL.n49 B 0.020001f
C85 VTAIL.n50 B 0.020001f
C86 VTAIL.n51 B 0.00896f
C87 VTAIL.n52 B 0.008462f
C88 VTAIL.n53 B 0.015748f
C89 VTAIL.n54 B 0.015748f
C90 VTAIL.n55 B 0.008462f
C91 VTAIL.n56 B 0.00896f
C92 VTAIL.n57 B 0.020001f
C93 VTAIL.n58 B 0.020001f
C94 VTAIL.n59 B 0.00896f
C95 VTAIL.n60 B 0.008462f
C96 VTAIL.n61 B 0.015748f
C97 VTAIL.n62 B 0.015748f
C98 VTAIL.n63 B 0.008462f
C99 VTAIL.n64 B 0.00896f
C100 VTAIL.n65 B 0.020001f
C101 VTAIL.n66 B 0.020001f
C102 VTAIL.n67 B 0.00896f
C103 VTAIL.n68 B 0.008462f
C104 VTAIL.n69 B 0.015748f
C105 VTAIL.n70 B 0.015748f
C106 VTAIL.n71 B 0.008462f
C107 VTAIL.n72 B 0.008462f
C108 VTAIL.n73 B 0.00896f
C109 VTAIL.n74 B 0.020001f
C110 VTAIL.n75 B 0.020001f
C111 VTAIL.n76 B 0.020001f
C112 VTAIL.n77 B 0.008711f
C113 VTAIL.n78 B 0.008462f
C114 VTAIL.n79 B 0.015748f
C115 VTAIL.n80 B 0.015748f
C116 VTAIL.n81 B 0.008462f
C117 VTAIL.n82 B 0.00896f
C118 VTAIL.n83 B 0.020001f
C119 VTAIL.n84 B 0.020001f
C120 VTAIL.n85 B 0.00896f
C121 VTAIL.n86 B 0.008462f
C122 VTAIL.n87 B 0.015748f
C123 VTAIL.n88 B 0.015748f
C124 VTAIL.n89 B 0.008462f
C125 VTAIL.n90 B 0.00896f
C126 VTAIL.n91 B 0.020001f
C127 VTAIL.n92 B 0.04236f
C128 VTAIL.n93 B 0.00896f
C129 VTAIL.n94 B 0.008462f
C130 VTAIL.n95 B 0.036185f
C131 VTAIL.n96 B 0.023599f
C132 VTAIL.n97 B 0.123235f
C133 VTAIL.n98 B 0.021604f
C134 VTAIL.n99 B 0.015748f
C135 VTAIL.n100 B 0.008462f
C136 VTAIL.n101 B 0.020001f
C137 VTAIL.n102 B 0.00896f
C138 VTAIL.n103 B 0.015748f
C139 VTAIL.n104 B 0.008462f
C140 VTAIL.n105 B 0.020001f
C141 VTAIL.n106 B 0.008711f
C142 VTAIL.n107 B 0.015748f
C143 VTAIL.n108 B 0.00896f
C144 VTAIL.n109 B 0.020001f
C145 VTAIL.n110 B 0.00896f
C146 VTAIL.n111 B 0.015748f
C147 VTAIL.n112 B 0.008462f
C148 VTAIL.n113 B 0.020001f
C149 VTAIL.n114 B 0.00896f
C150 VTAIL.n115 B 0.015748f
C151 VTAIL.n116 B 0.008462f
C152 VTAIL.n117 B 0.020001f
C153 VTAIL.n118 B 0.00896f
C154 VTAIL.n119 B 0.015748f
C155 VTAIL.n120 B 0.008462f
C156 VTAIL.n121 B 0.020001f
C157 VTAIL.n122 B 0.00896f
C158 VTAIL.n123 B 0.015748f
C159 VTAIL.n124 B 0.008462f
C160 VTAIL.n125 B 0.020001f
C161 VTAIL.n126 B 0.00896f
C162 VTAIL.n127 B 1.20573f
C163 VTAIL.n128 B 0.008462f
C164 VTAIL.t7 B 0.033116f
C165 VTAIL.n129 B 0.112621f
C166 VTAIL.n130 B 0.011816f
C167 VTAIL.n131 B 0.015001f
C168 VTAIL.n132 B 0.020001f
C169 VTAIL.n133 B 0.00896f
C170 VTAIL.n134 B 0.008462f
C171 VTAIL.n135 B 0.015748f
C172 VTAIL.n136 B 0.015748f
C173 VTAIL.n137 B 0.008462f
C174 VTAIL.n138 B 0.00896f
C175 VTAIL.n139 B 0.020001f
C176 VTAIL.n140 B 0.020001f
C177 VTAIL.n141 B 0.00896f
C178 VTAIL.n142 B 0.008462f
C179 VTAIL.n143 B 0.015748f
C180 VTAIL.n144 B 0.015748f
C181 VTAIL.n145 B 0.008462f
C182 VTAIL.n146 B 0.00896f
C183 VTAIL.n147 B 0.020001f
C184 VTAIL.n148 B 0.020001f
C185 VTAIL.n149 B 0.00896f
C186 VTAIL.n150 B 0.008462f
C187 VTAIL.n151 B 0.015748f
C188 VTAIL.n152 B 0.015748f
C189 VTAIL.n153 B 0.008462f
C190 VTAIL.n154 B 0.00896f
C191 VTAIL.n155 B 0.020001f
C192 VTAIL.n156 B 0.020001f
C193 VTAIL.n157 B 0.00896f
C194 VTAIL.n158 B 0.008462f
C195 VTAIL.n159 B 0.015748f
C196 VTAIL.n160 B 0.015748f
C197 VTAIL.n161 B 0.008462f
C198 VTAIL.n162 B 0.00896f
C199 VTAIL.n163 B 0.020001f
C200 VTAIL.n164 B 0.020001f
C201 VTAIL.n165 B 0.00896f
C202 VTAIL.n166 B 0.008462f
C203 VTAIL.n167 B 0.015748f
C204 VTAIL.n168 B 0.015748f
C205 VTAIL.n169 B 0.008462f
C206 VTAIL.n170 B 0.008462f
C207 VTAIL.n171 B 0.00896f
C208 VTAIL.n172 B 0.020001f
C209 VTAIL.n173 B 0.020001f
C210 VTAIL.n174 B 0.020001f
C211 VTAIL.n175 B 0.008711f
C212 VTAIL.n176 B 0.008462f
C213 VTAIL.n177 B 0.015748f
C214 VTAIL.n178 B 0.015748f
C215 VTAIL.n179 B 0.008462f
C216 VTAIL.n180 B 0.00896f
C217 VTAIL.n181 B 0.020001f
C218 VTAIL.n182 B 0.020001f
C219 VTAIL.n183 B 0.00896f
C220 VTAIL.n184 B 0.008462f
C221 VTAIL.n185 B 0.015748f
C222 VTAIL.n186 B 0.015748f
C223 VTAIL.n187 B 0.008462f
C224 VTAIL.n188 B 0.00896f
C225 VTAIL.n189 B 0.020001f
C226 VTAIL.n190 B 0.04236f
C227 VTAIL.n191 B 0.00896f
C228 VTAIL.n192 B 0.008462f
C229 VTAIL.n193 B 0.036185f
C230 VTAIL.n194 B 0.023599f
C231 VTAIL.n195 B 0.203395f
C232 VTAIL.n196 B 0.021604f
C233 VTAIL.n197 B 0.015748f
C234 VTAIL.n198 B 0.008462f
C235 VTAIL.n199 B 0.020001f
C236 VTAIL.n200 B 0.00896f
C237 VTAIL.n201 B 0.015748f
C238 VTAIL.n202 B 0.008462f
C239 VTAIL.n203 B 0.020001f
C240 VTAIL.n204 B 0.008711f
C241 VTAIL.n205 B 0.015748f
C242 VTAIL.n206 B 0.00896f
C243 VTAIL.n207 B 0.020001f
C244 VTAIL.n208 B 0.00896f
C245 VTAIL.n209 B 0.015748f
C246 VTAIL.n210 B 0.008462f
C247 VTAIL.n211 B 0.020001f
C248 VTAIL.n212 B 0.00896f
C249 VTAIL.n213 B 0.015748f
C250 VTAIL.n214 B 0.008462f
C251 VTAIL.n215 B 0.020001f
C252 VTAIL.n216 B 0.00896f
C253 VTAIL.n217 B 0.015748f
C254 VTAIL.n218 B 0.008462f
C255 VTAIL.n219 B 0.020001f
C256 VTAIL.n220 B 0.00896f
C257 VTAIL.n221 B 0.015748f
C258 VTAIL.n222 B 0.008462f
C259 VTAIL.n223 B 0.020001f
C260 VTAIL.n224 B 0.00896f
C261 VTAIL.n225 B 1.20573f
C262 VTAIL.n226 B 0.008462f
C263 VTAIL.t5 B 0.033116f
C264 VTAIL.n227 B 0.112621f
C265 VTAIL.n228 B 0.011816f
C266 VTAIL.n229 B 0.015001f
C267 VTAIL.n230 B 0.020001f
C268 VTAIL.n231 B 0.00896f
C269 VTAIL.n232 B 0.008462f
C270 VTAIL.n233 B 0.015748f
C271 VTAIL.n234 B 0.015748f
C272 VTAIL.n235 B 0.008462f
C273 VTAIL.n236 B 0.00896f
C274 VTAIL.n237 B 0.020001f
C275 VTAIL.n238 B 0.020001f
C276 VTAIL.n239 B 0.00896f
C277 VTAIL.n240 B 0.008462f
C278 VTAIL.n241 B 0.015748f
C279 VTAIL.n242 B 0.015748f
C280 VTAIL.n243 B 0.008462f
C281 VTAIL.n244 B 0.00896f
C282 VTAIL.n245 B 0.020001f
C283 VTAIL.n246 B 0.020001f
C284 VTAIL.n247 B 0.00896f
C285 VTAIL.n248 B 0.008462f
C286 VTAIL.n249 B 0.015748f
C287 VTAIL.n250 B 0.015748f
C288 VTAIL.n251 B 0.008462f
C289 VTAIL.n252 B 0.00896f
C290 VTAIL.n253 B 0.020001f
C291 VTAIL.n254 B 0.020001f
C292 VTAIL.n255 B 0.00896f
C293 VTAIL.n256 B 0.008462f
C294 VTAIL.n257 B 0.015748f
C295 VTAIL.n258 B 0.015748f
C296 VTAIL.n259 B 0.008462f
C297 VTAIL.n260 B 0.00896f
C298 VTAIL.n261 B 0.020001f
C299 VTAIL.n262 B 0.020001f
C300 VTAIL.n263 B 0.00896f
C301 VTAIL.n264 B 0.008462f
C302 VTAIL.n265 B 0.015748f
C303 VTAIL.n266 B 0.015748f
C304 VTAIL.n267 B 0.008462f
C305 VTAIL.n268 B 0.008462f
C306 VTAIL.n269 B 0.00896f
C307 VTAIL.n270 B 0.020001f
C308 VTAIL.n271 B 0.020001f
C309 VTAIL.n272 B 0.020001f
C310 VTAIL.n273 B 0.008711f
C311 VTAIL.n274 B 0.008462f
C312 VTAIL.n275 B 0.015748f
C313 VTAIL.n276 B 0.015748f
C314 VTAIL.n277 B 0.008462f
C315 VTAIL.n278 B 0.00896f
C316 VTAIL.n279 B 0.020001f
C317 VTAIL.n280 B 0.020001f
C318 VTAIL.n281 B 0.00896f
C319 VTAIL.n282 B 0.008462f
C320 VTAIL.n283 B 0.015748f
C321 VTAIL.n284 B 0.015748f
C322 VTAIL.n285 B 0.008462f
C323 VTAIL.n286 B 0.00896f
C324 VTAIL.n287 B 0.020001f
C325 VTAIL.n288 B 0.04236f
C326 VTAIL.n289 B 0.00896f
C327 VTAIL.n290 B 0.008462f
C328 VTAIL.n291 B 0.036185f
C329 VTAIL.n292 B 0.023599f
C330 VTAIL.n293 B 1.32565f
C331 VTAIL.n294 B 0.021604f
C332 VTAIL.n295 B 0.015748f
C333 VTAIL.n296 B 0.008462f
C334 VTAIL.n297 B 0.020001f
C335 VTAIL.n298 B 0.00896f
C336 VTAIL.n299 B 0.015748f
C337 VTAIL.n300 B 0.008462f
C338 VTAIL.n301 B 0.020001f
C339 VTAIL.n302 B 0.008711f
C340 VTAIL.n303 B 0.015748f
C341 VTAIL.n304 B 0.008711f
C342 VTAIL.n305 B 0.008462f
C343 VTAIL.n306 B 0.020001f
C344 VTAIL.n307 B 0.020001f
C345 VTAIL.n308 B 0.00896f
C346 VTAIL.n309 B 0.015748f
C347 VTAIL.n310 B 0.008462f
C348 VTAIL.n311 B 0.020001f
C349 VTAIL.n312 B 0.00896f
C350 VTAIL.n313 B 0.015748f
C351 VTAIL.n314 B 0.008462f
C352 VTAIL.n315 B 0.020001f
C353 VTAIL.n316 B 0.00896f
C354 VTAIL.n317 B 0.015748f
C355 VTAIL.n318 B 0.008462f
C356 VTAIL.n319 B 0.020001f
C357 VTAIL.n320 B 0.00896f
C358 VTAIL.n321 B 0.015748f
C359 VTAIL.n322 B 0.008462f
C360 VTAIL.n323 B 0.020001f
C361 VTAIL.n324 B 0.00896f
C362 VTAIL.n325 B 1.20573f
C363 VTAIL.n326 B 0.008462f
C364 VTAIL.t3 B 0.033116f
C365 VTAIL.n327 B 0.112621f
C366 VTAIL.n328 B 0.011816f
C367 VTAIL.n329 B 0.015001f
C368 VTAIL.n330 B 0.020001f
C369 VTAIL.n331 B 0.00896f
C370 VTAIL.n332 B 0.008462f
C371 VTAIL.n333 B 0.015748f
C372 VTAIL.n334 B 0.015748f
C373 VTAIL.n335 B 0.008462f
C374 VTAIL.n336 B 0.00896f
C375 VTAIL.n337 B 0.020001f
C376 VTAIL.n338 B 0.020001f
C377 VTAIL.n339 B 0.00896f
C378 VTAIL.n340 B 0.008462f
C379 VTAIL.n341 B 0.015748f
C380 VTAIL.n342 B 0.015748f
C381 VTAIL.n343 B 0.008462f
C382 VTAIL.n344 B 0.00896f
C383 VTAIL.n345 B 0.020001f
C384 VTAIL.n346 B 0.020001f
C385 VTAIL.n347 B 0.00896f
C386 VTAIL.n348 B 0.008462f
C387 VTAIL.n349 B 0.015748f
C388 VTAIL.n350 B 0.015748f
C389 VTAIL.n351 B 0.008462f
C390 VTAIL.n352 B 0.00896f
C391 VTAIL.n353 B 0.020001f
C392 VTAIL.n354 B 0.020001f
C393 VTAIL.n355 B 0.00896f
C394 VTAIL.n356 B 0.008462f
C395 VTAIL.n357 B 0.015748f
C396 VTAIL.n358 B 0.015748f
C397 VTAIL.n359 B 0.008462f
C398 VTAIL.n360 B 0.00896f
C399 VTAIL.n361 B 0.020001f
C400 VTAIL.n362 B 0.020001f
C401 VTAIL.n363 B 0.00896f
C402 VTAIL.n364 B 0.008462f
C403 VTAIL.n365 B 0.015748f
C404 VTAIL.n366 B 0.015748f
C405 VTAIL.n367 B 0.008462f
C406 VTAIL.n368 B 0.00896f
C407 VTAIL.n369 B 0.020001f
C408 VTAIL.n370 B 0.020001f
C409 VTAIL.n371 B 0.00896f
C410 VTAIL.n372 B 0.008462f
C411 VTAIL.n373 B 0.015748f
C412 VTAIL.n374 B 0.015748f
C413 VTAIL.n375 B 0.008462f
C414 VTAIL.n376 B 0.00896f
C415 VTAIL.n377 B 0.020001f
C416 VTAIL.n378 B 0.020001f
C417 VTAIL.n379 B 0.00896f
C418 VTAIL.n380 B 0.008462f
C419 VTAIL.n381 B 0.015748f
C420 VTAIL.n382 B 0.015748f
C421 VTAIL.n383 B 0.008462f
C422 VTAIL.n384 B 0.00896f
C423 VTAIL.n385 B 0.020001f
C424 VTAIL.n386 B 0.04236f
C425 VTAIL.n387 B 0.00896f
C426 VTAIL.n388 B 0.008462f
C427 VTAIL.n389 B 0.036185f
C428 VTAIL.n390 B 0.023599f
C429 VTAIL.n391 B 1.32565f
C430 VTAIL.n392 B 0.021604f
C431 VTAIL.n393 B 0.015748f
C432 VTAIL.n394 B 0.008462f
C433 VTAIL.n395 B 0.020001f
C434 VTAIL.n396 B 0.00896f
C435 VTAIL.n397 B 0.015748f
C436 VTAIL.n398 B 0.008462f
C437 VTAIL.n399 B 0.020001f
C438 VTAIL.n400 B 0.008711f
C439 VTAIL.n401 B 0.015748f
C440 VTAIL.n402 B 0.008711f
C441 VTAIL.n403 B 0.008462f
C442 VTAIL.n404 B 0.020001f
C443 VTAIL.n405 B 0.020001f
C444 VTAIL.n406 B 0.00896f
C445 VTAIL.n407 B 0.015748f
C446 VTAIL.n408 B 0.008462f
C447 VTAIL.n409 B 0.020001f
C448 VTAIL.n410 B 0.00896f
C449 VTAIL.n411 B 0.015748f
C450 VTAIL.n412 B 0.008462f
C451 VTAIL.n413 B 0.020001f
C452 VTAIL.n414 B 0.00896f
C453 VTAIL.n415 B 0.015748f
C454 VTAIL.n416 B 0.008462f
C455 VTAIL.n417 B 0.020001f
C456 VTAIL.n418 B 0.00896f
C457 VTAIL.n419 B 0.015748f
C458 VTAIL.n420 B 0.008462f
C459 VTAIL.n421 B 0.020001f
C460 VTAIL.n422 B 0.00896f
C461 VTAIL.n423 B 1.20573f
C462 VTAIL.n424 B 0.008462f
C463 VTAIL.t2 B 0.033116f
C464 VTAIL.n425 B 0.112621f
C465 VTAIL.n426 B 0.011816f
C466 VTAIL.n427 B 0.015001f
C467 VTAIL.n428 B 0.020001f
C468 VTAIL.n429 B 0.00896f
C469 VTAIL.n430 B 0.008462f
C470 VTAIL.n431 B 0.015748f
C471 VTAIL.n432 B 0.015748f
C472 VTAIL.n433 B 0.008462f
C473 VTAIL.n434 B 0.00896f
C474 VTAIL.n435 B 0.020001f
C475 VTAIL.n436 B 0.020001f
C476 VTAIL.n437 B 0.00896f
C477 VTAIL.n438 B 0.008462f
C478 VTAIL.n439 B 0.015748f
C479 VTAIL.n440 B 0.015748f
C480 VTAIL.n441 B 0.008462f
C481 VTAIL.n442 B 0.00896f
C482 VTAIL.n443 B 0.020001f
C483 VTAIL.n444 B 0.020001f
C484 VTAIL.n445 B 0.00896f
C485 VTAIL.n446 B 0.008462f
C486 VTAIL.n447 B 0.015748f
C487 VTAIL.n448 B 0.015748f
C488 VTAIL.n449 B 0.008462f
C489 VTAIL.n450 B 0.00896f
C490 VTAIL.n451 B 0.020001f
C491 VTAIL.n452 B 0.020001f
C492 VTAIL.n453 B 0.00896f
C493 VTAIL.n454 B 0.008462f
C494 VTAIL.n455 B 0.015748f
C495 VTAIL.n456 B 0.015748f
C496 VTAIL.n457 B 0.008462f
C497 VTAIL.n458 B 0.00896f
C498 VTAIL.n459 B 0.020001f
C499 VTAIL.n460 B 0.020001f
C500 VTAIL.n461 B 0.00896f
C501 VTAIL.n462 B 0.008462f
C502 VTAIL.n463 B 0.015748f
C503 VTAIL.n464 B 0.015748f
C504 VTAIL.n465 B 0.008462f
C505 VTAIL.n466 B 0.00896f
C506 VTAIL.n467 B 0.020001f
C507 VTAIL.n468 B 0.020001f
C508 VTAIL.n469 B 0.00896f
C509 VTAIL.n470 B 0.008462f
C510 VTAIL.n471 B 0.015748f
C511 VTAIL.n472 B 0.015748f
C512 VTAIL.n473 B 0.008462f
C513 VTAIL.n474 B 0.00896f
C514 VTAIL.n475 B 0.020001f
C515 VTAIL.n476 B 0.020001f
C516 VTAIL.n477 B 0.00896f
C517 VTAIL.n478 B 0.008462f
C518 VTAIL.n479 B 0.015748f
C519 VTAIL.n480 B 0.015748f
C520 VTAIL.n481 B 0.008462f
C521 VTAIL.n482 B 0.00896f
C522 VTAIL.n483 B 0.020001f
C523 VTAIL.n484 B 0.04236f
C524 VTAIL.n485 B 0.00896f
C525 VTAIL.n486 B 0.008462f
C526 VTAIL.n487 B 0.036185f
C527 VTAIL.n488 B 0.023599f
C528 VTAIL.n489 B 0.203395f
C529 VTAIL.n490 B 0.021604f
C530 VTAIL.n491 B 0.015748f
C531 VTAIL.n492 B 0.008462f
C532 VTAIL.n493 B 0.020001f
C533 VTAIL.n494 B 0.00896f
C534 VTAIL.n495 B 0.015748f
C535 VTAIL.n496 B 0.008462f
C536 VTAIL.n497 B 0.020001f
C537 VTAIL.n498 B 0.008711f
C538 VTAIL.n499 B 0.015748f
C539 VTAIL.n500 B 0.008711f
C540 VTAIL.n501 B 0.008462f
C541 VTAIL.n502 B 0.020001f
C542 VTAIL.n503 B 0.020001f
C543 VTAIL.n504 B 0.00896f
C544 VTAIL.n505 B 0.015748f
C545 VTAIL.n506 B 0.008462f
C546 VTAIL.n507 B 0.020001f
C547 VTAIL.n508 B 0.00896f
C548 VTAIL.n509 B 0.015748f
C549 VTAIL.n510 B 0.008462f
C550 VTAIL.n511 B 0.020001f
C551 VTAIL.n512 B 0.00896f
C552 VTAIL.n513 B 0.015748f
C553 VTAIL.n514 B 0.008462f
C554 VTAIL.n515 B 0.020001f
C555 VTAIL.n516 B 0.00896f
C556 VTAIL.n517 B 0.015748f
C557 VTAIL.n518 B 0.008462f
C558 VTAIL.n519 B 0.020001f
C559 VTAIL.n520 B 0.00896f
C560 VTAIL.n521 B 1.20573f
C561 VTAIL.n522 B 0.008462f
C562 VTAIL.t6 B 0.033116f
C563 VTAIL.n523 B 0.112621f
C564 VTAIL.n524 B 0.011816f
C565 VTAIL.n525 B 0.015001f
C566 VTAIL.n526 B 0.020001f
C567 VTAIL.n527 B 0.00896f
C568 VTAIL.n528 B 0.008462f
C569 VTAIL.n529 B 0.015748f
C570 VTAIL.n530 B 0.015748f
C571 VTAIL.n531 B 0.008462f
C572 VTAIL.n532 B 0.00896f
C573 VTAIL.n533 B 0.020001f
C574 VTAIL.n534 B 0.020001f
C575 VTAIL.n535 B 0.00896f
C576 VTAIL.n536 B 0.008462f
C577 VTAIL.n537 B 0.015748f
C578 VTAIL.n538 B 0.015748f
C579 VTAIL.n539 B 0.008462f
C580 VTAIL.n540 B 0.00896f
C581 VTAIL.n541 B 0.020001f
C582 VTAIL.n542 B 0.020001f
C583 VTAIL.n543 B 0.00896f
C584 VTAIL.n544 B 0.008462f
C585 VTAIL.n545 B 0.015748f
C586 VTAIL.n546 B 0.015748f
C587 VTAIL.n547 B 0.008462f
C588 VTAIL.n548 B 0.00896f
C589 VTAIL.n549 B 0.020001f
C590 VTAIL.n550 B 0.020001f
C591 VTAIL.n551 B 0.00896f
C592 VTAIL.n552 B 0.008462f
C593 VTAIL.n553 B 0.015748f
C594 VTAIL.n554 B 0.015748f
C595 VTAIL.n555 B 0.008462f
C596 VTAIL.n556 B 0.00896f
C597 VTAIL.n557 B 0.020001f
C598 VTAIL.n558 B 0.020001f
C599 VTAIL.n559 B 0.00896f
C600 VTAIL.n560 B 0.008462f
C601 VTAIL.n561 B 0.015748f
C602 VTAIL.n562 B 0.015748f
C603 VTAIL.n563 B 0.008462f
C604 VTAIL.n564 B 0.00896f
C605 VTAIL.n565 B 0.020001f
C606 VTAIL.n566 B 0.020001f
C607 VTAIL.n567 B 0.00896f
C608 VTAIL.n568 B 0.008462f
C609 VTAIL.n569 B 0.015748f
C610 VTAIL.n570 B 0.015748f
C611 VTAIL.n571 B 0.008462f
C612 VTAIL.n572 B 0.00896f
C613 VTAIL.n573 B 0.020001f
C614 VTAIL.n574 B 0.020001f
C615 VTAIL.n575 B 0.00896f
C616 VTAIL.n576 B 0.008462f
C617 VTAIL.n577 B 0.015748f
C618 VTAIL.n578 B 0.015748f
C619 VTAIL.n579 B 0.008462f
C620 VTAIL.n580 B 0.00896f
C621 VTAIL.n581 B 0.020001f
C622 VTAIL.n582 B 0.04236f
C623 VTAIL.n583 B 0.00896f
C624 VTAIL.n584 B 0.008462f
C625 VTAIL.n585 B 0.036185f
C626 VTAIL.n586 B 0.023599f
C627 VTAIL.n587 B 0.203395f
C628 VTAIL.n588 B 0.021604f
C629 VTAIL.n589 B 0.015748f
C630 VTAIL.n590 B 0.008462f
C631 VTAIL.n591 B 0.020001f
C632 VTAIL.n592 B 0.00896f
C633 VTAIL.n593 B 0.015748f
C634 VTAIL.n594 B 0.008462f
C635 VTAIL.n595 B 0.020001f
C636 VTAIL.n596 B 0.008711f
C637 VTAIL.n597 B 0.015748f
C638 VTAIL.n598 B 0.008711f
C639 VTAIL.n599 B 0.008462f
C640 VTAIL.n600 B 0.020001f
C641 VTAIL.n601 B 0.020001f
C642 VTAIL.n602 B 0.00896f
C643 VTAIL.n603 B 0.015748f
C644 VTAIL.n604 B 0.008462f
C645 VTAIL.n605 B 0.020001f
C646 VTAIL.n606 B 0.00896f
C647 VTAIL.n607 B 0.015748f
C648 VTAIL.n608 B 0.008462f
C649 VTAIL.n609 B 0.020001f
C650 VTAIL.n610 B 0.00896f
C651 VTAIL.n611 B 0.015748f
C652 VTAIL.n612 B 0.008462f
C653 VTAIL.n613 B 0.020001f
C654 VTAIL.n614 B 0.00896f
C655 VTAIL.n615 B 0.015748f
C656 VTAIL.n616 B 0.008462f
C657 VTAIL.n617 B 0.020001f
C658 VTAIL.n618 B 0.00896f
C659 VTAIL.n619 B 1.20573f
C660 VTAIL.n620 B 0.008462f
C661 VTAIL.t4 B 0.033116f
C662 VTAIL.n621 B 0.112621f
C663 VTAIL.n622 B 0.011816f
C664 VTAIL.n623 B 0.015001f
C665 VTAIL.n624 B 0.020001f
C666 VTAIL.n625 B 0.00896f
C667 VTAIL.n626 B 0.008462f
C668 VTAIL.n627 B 0.015748f
C669 VTAIL.n628 B 0.015748f
C670 VTAIL.n629 B 0.008462f
C671 VTAIL.n630 B 0.00896f
C672 VTAIL.n631 B 0.020001f
C673 VTAIL.n632 B 0.020001f
C674 VTAIL.n633 B 0.00896f
C675 VTAIL.n634 B 0.008462f
C676 VTAIL.n635 B 0.015748f
C677 VTAIL.n636 B 0.015748f
C678 VTAIL.n637 B 0.008462f
C679 VTAIL.n638 B 0.00896f
C680 VTAIL.n639 B 0.020001f
C681 VTAIL.n640 B 0.020001f
C682 VTAIL.n641 B 0.00896f
C683 VTAIL.n642 B 0.008462f
C684 VTAIL.n643 B 0.015748f
C685 VTAIL.n644 B 0.015748f
C686 VTAIL.n645 B 0.008462f
C687 VTAIL.n646 B 0.00896f
C688 VTAIL.n647 B 0.020001f
C689 VTAIL.n648 B 0.020001f
C690 VTAIL.n649 B 0.00896f
C691 VTAIL.n650 B 0.008462f
C692 VTAIL.n651 B 0.015748f
C693 VTAIL.n652 B 0.015748f
C694 VTAIL.n653 B 0.008462f
C695 VTAIL.n654 B 0.00896f
C696 VTAIL.n655 B 0.020001f
C697 VTAIL.n656 B 0.020001f
C698 VTAIL.n657 B 0.00896f
C699 VTAIL.n658 B 0.008462f
C700 VTAIL.n659 B 0.015748f
C701 VTAIL.n660 B 0.015748f
C702 VTAIL.n661 B 0.008462f
C703 VTAIL.n662 B 0.00896f
C704 VTAIL.n663 B 0.020001f
C705 VTAIL.n664 B 0.020001f
C706 VTAIL.n665 B 0.00896f
C707 VTAIL.n666 B 0.008462f
C708 VTAIL.n667 B 0.015748f
C709 VTAIL.n668 B 0.015748f
C710 VTAIL.n669 B 0.008462f
C711 VTAIL.n670 B 0.00896f
C712 VTAIL.n671 B 0.020001f
C713 VTAIL.n672 B 0.020001f
C714 VTAIL.n673 B 0.00896f
C715 VTAIL.n674 B 0.008462f
C716 VTAIL.n675 B 0.015748f
C717 VTAIL.n676 B 0.015748f
C718 VTAIL.n677 B 0.008462f
C719 VTAIL.n678 B 0.00896f
C720 VTAIL.n679 B 0.020001f
C721 VTAIL.n680 B 0.04236f
C722 VTAIL.n681 B 0.00896f
C723 VTAIL.n682 B 0.008462f
C724 VTAIL.n683 B 0.036185f
C725 VTAIL.n684 B 0.023599f
C726 VTAIL.n685 B 1.32565f
C727 VTAIL.n686 B 0.021604f
C728 VTAIL.n687 B 0.015748f
C729 VTAIL.n688 B 0.008462f
C730 VTAIL.n689 B 0.020001f
C731 VTAIL.n690 B 0.00896f
C732 VTAIL.n691 B 0.015748f
C733 VTAIL.n692 B 0.008462f
C734 VTAIL.n693 B 0.020001f
C735 VTAIL.n694 B 0.008711f
C736 VTAIL.n695 B 0.015748f
C737 VTAIL.n696 B 0.00896f
C738 VTAIL.n697 B 0.020001f
C739 VTAIL.n698 B 0.00896f
C740 VTAIL.n699 B 0.015748f
C741 VTAIL.n700 B 0.008462f
C742 VTAIL.n701 B 0.020001f
C743 VTAIL.n702 B 0.00896f
C744 VTAIL.n703 B 0.015748f
C745 VTAIL.n704 B 0.008462f
C746 VTAIL.n705 B 0.020001f
C747 VTAIL.n706 B 0.00896f
C748 VTAIL.n707 B 0.015748f
C749 VTAIL.n708 B 0.008462f
C750 VTAIL.n709 B 0.020001f
C751 VTAIL.n710 B 0.00896f
C752 VTAIL.n711 B 0.015748f
C753 VTAIL.n712 B 0.008462f
C754 VTAIL.n713 B 0.020001f
C755 VTAIL.n714 B 0.00896f
C756 VTAIL.n715 B 1.20573f
C757 VTAIL.n716 B 0.008462f
C758 VTAIL.t0 B 0.033116f
C759 VTAIL.n717 B 0.112621f
C760 VTAIL.n718 B 0.011816f
C761 VTAIL.n719 B 0.015001f
C762 VTAIL.n720 B 0.020001f
C763 VTAIL.n721 B 0.00896f
C764 VTAIL.n722 B 0.008462f
C765 VTAIL.n723 B 0.015748f
C766 VTAIL.n724 B 0.015748f
C767 VTAIL.n725 B 0.008462f
C768 VTAIL.n726 B 0.00896f
C769 VTAIL.n727 B 0.020001f
C770 VTAIL.n728 B 0.020001f
C771 VTAIL.n729 B 0.00896f
C772 VTAIL.n730 B 0.008462f
C773 VTAIL.n731 B 0.015748f
C774 VTAIL.n732 B 0.015748f
C775 VTAIL.n733 B 0.008462f
C776 VTAIL.n734 B 0.00896f
C777 VTAIL.n735 B 0.020001f
C778 VTAIL.n736 B 0.020001f
C779 VTAIL.n737 B 0.00896f
C780 VTAIL.n738 B 0.008462f
C781 VTAIL.n739 B 0.015748f
C782 VTAIL.n740 B 0.015748f
C783 VTAIL.n741 B 0.008462f
C784 VTAIL.n742 B 0.00896f
C785 VTAIL.n743 B 0.020001f
C786 VTAIL.n744 B 0.020001f
C787 VTAIL.n745 B 0.00896f
C788 VTAIL.n746 B 0.008462f
C789 VTAIL.n747 B 0.015748f
C790 VTAIL.n748 B 0.015748f
C791 VTAIL.n749 B 0.008462f
C792 VTAIL.n750 B 0.00896f
C793 VTAIL.n751 B 0.020001f
C794 VTAIL.n752 B 0.020001f
C795 VTAIL.n753 B 0.00896f
C796 VTAIL.n754 B 0.008462f
C797 VTAIL.n755 B 0.015748f
C798 VTAIL.n756 B 0.015748f
C799 VTAIL.n757 B 0.008462f
C800 VTAIL.n758 B 0.008462f
C801 VTAIL.n759 B 0.00896f
C802 VTAIL.n760 B 0.020001f
C803 VTAIL.n761 B 0.020001f
C804 VTAIL.n762 B 0.020001f
C805 VTAIL.n763 B 0.008711f
C806 VTAIL.n764 B 0.008462f
C807 VTAIL.n765 B 0.015748f
C808 VTAIL.n766 B 0.015748f
C809 VTAIL.n767 B 0.008462f
C810 VTAIL.n768 B 0.00896f
C811 VTAIL.n769 B 0.020001f
C812 VTAIL.n770 B 0.020001f
C813 VTAIL.n771 B 0.00896f
C814 VTAIL.n772 B 0.008462f
C815 VTAIL.n773 B 0.015748f
C816 VTAIL.n774 B 0.015748f
C817 VTAIL.n775 B 0.008462f
C818 VTAIL.n776 B 0.00896f
C819 VTAIL.n777 B 0.020001f
C820 VTAIL.n778 B 0.04236f
C821 VTAIL.n779 B 0.00896f
C822 VTAIL.n780 B 0.008462f
C823 VTAIL.n781 B 0.036185f
C824 VTAIL.n782 B 0.023599f
C825 VTAIL.n783 B 1.23959f
C826 VP.t0 B 3.37657f
C827 VP.n0 B 1.24029f
C828 VP.n1 B 0.020215f
C829 VP.n2 B 0.02951f
C830 VP.n3 B 0.020215f
C831 VP.n4 B 0.024655f
C832 VP.t1 B 3.66736f
C833 VP.t3 B 3.65744f
C834 VP.n5 B 3.66522f
C835 VP.t2 B 3.37657f
C836 VP.n6 B 1.24029f
C837 VP.n7 B 1.33591f
C838 VP.n8 B 0.032626f
C839 VP.n9 B 0.020215f
C840 VP.n10 B 0.037675f
C841 VP.n11 B 0.037675f
C842 VP.n12 B 0.02951f
C843 VP.n13 B 0.020215f
C844 VP.n14 B 0.020215f
C845 VP.n15 B 0.020215f
C846 VP.n16 B 0.037675f
C847 VP.n17 B 0.037675f
C848 VP.n18 B 0.024655f
C849 VP.n19 B 0.032626f
C850 VP.n20 B 0.055797f
.ends

