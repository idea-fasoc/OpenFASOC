* NGSPICE file created from diff_pair_sample_0449.ext - technology: sky130A

.subckt diff_pair_sample_0449 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=1.79
X1 VDD2.t7 VN.t0 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=1.79
X2 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=1.79
X3 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=1.79
X4 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=1.79
X5 VTAIL.t11 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X6 VTAIL.t10 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=1.79
X7 VDD2.t4 VN.t3 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X8 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=1.79
X9 VDD2.t3 VN.t4 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X10 VDD2.t2 VN.t5 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=1.79
X11 VTAIL.t12 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X12 VDD1.t6 VP.t1 VTAIL.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X13 VTAIL.t0 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=1.79
X14 VTAIL.t1 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=1.79
X15 VDD1.t3 VP.t4 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=1.79
X16 VTAIL.t3 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X17 VTAIL.t8 VN.t7 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=1.79
X18 VDD1.t1 VP.t6 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
X19 VTAIL.t4 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=1.79
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n20 VP.n19 161.3
R5 VP.n21 VP.n7 161.3
R6 VP.n23 VP.n22 161.3
R7 VP.n24 VP.n6 161.3
R8 VP.n48 VP.n0 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n1 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n41 VP.n2 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n3 161.3
R15 VP.n37 VP.n36 161.3
R16 VP.n34 VP.n4 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n31 VP.n5 161.3
R19 VP.n30 VP.n29 161.3
R20 VP.n10 VP.t2 95.6032
R21 VP.n28 VP.n27 89.7148
R22 VP.n50 VP.n49 89.7148
R23 VP.n26 VP.n25 89.7148
R24 VP.n28 VP.t3 64.7608
R25 VP.n35 VP.t1 64.7608
R26 VP.n42 VP.t7 64.7608
R27 VP.n49 VP.t0 64.7608
R28 VP.n25 VP.t4 64.7608
R29 VP.n18 VP.t5 64.7608
R30 VP.n11 VP.t6 64.7608
R31 VP.n40 VP.n3 56.5193
R32 VP.n16 VP.n9 56.5193
R33 VP.n11 VP.n10 54.5414
R34 VP.n33 VP.n5 53.1199
R35 VP.n47 VP.n1 53.1199
R36 VP.n23 VP.n7 53.1199
R37 VP.n27 VP.n26 41.6511
R38 VP.n29 VP.n5 27.8669
R39 VP.n48 VP.n47 27.8669
R40 VP.n24 VP.n23 27.8669
R41 VP.n34 VP.n33 24.4675
R42 VP.n36 VP.n3 24.4675
R43 VP.n41 VP.n40 24.4675
R44 VP.n43 VP.n1 24.4675
R45 VP.n17 VP.n16 24.4675
R46 VP.n19 VP.n7 24.4675
R47 VP.n12 VP.n9 24.4675
R48 VP.n29 VP.n28 21.0421
R49 VP.n49 VP.n48 21.0421
R50 VP.n25 VP.n24 21.0421
R51 VP.n36 VP.n35 15.17
R52 VP.n42 VP.n41 15.17
R53 VP.n18 VP.n17 15.17
R54 VP.n12 VP.n11 15.17
R55 VP.n13 VP.n10 13.1161
R56 VP.n35 VP.n34 9.29796
R57 VP.n43 VP.n42 9.29796
R58 VP.n19 VP.n18 9.29796
R59 VP.n26 VP.n6 0.278367
R60 VP.n30 VP.n27 0.278367
R61 VP.n50 VP.n0 0.278367
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153454
R81 VTAIL.n11 VTAIL.t0 54.8713
R82 VTAIL.n10 VTAIL.t13 54.8713
R83 VTAIL.n7 VTAIL.t8 54.8713
R84 VTAIL.n15 VTAIL.t14 54.8712
R85 VTAIL.n2 VTAIL.t10 54.8712
R86 VTAIL.n3 VTAIL.t6 54.8712
R87 VTAIL.n6 VTAIL.t1 54.8712
R88 VTAIL.n14 VTAIL.t5 54.8712
R89 VTAIL.n13 VTAIL.n12 50.755
R90 VTAIL.n9 VTAIL.n8 50.755
R91 VTAIL.n1 VTAIL.n0 50.7547
R92 VTAIL.n5 VTAIL.n4 50.7547
R93 VTAIL.n15 VTAIL.n14 18.341
R94 VTAIL.n7 VTAIL.n6 18.341
R95 VTAIL.n0 VTAIL.t9 4.11692
R96 VTAIL.n0 VTAIL.t11 4.11692
R97 VTAIL.n4 VTAIL.t7 4.11692
R98 VTAIL.n4 VTAIL.t4 4.11692
R99 VTAIL.n12 VTAIL.t2 4.11692
R100 VTAIL.n12 VTAIL.t3 4.11692
R101 VTAIL.n8 VTAIL.t15 4.11692
R102 VTAIL.n8 VTAIL.t12 4.11692
R103 VTAIL.n9 VTAIL.n7 1.82809
R104 VTAIL.n10 VTAIL.n9 1.82809
R105 VTAIL.n13 VTAIL.n11 1.82809
R106 VTAIL.n14 VTAIL.n13 1.82809
R107 VTAIL.n6 VTAIL.n5 1.82809
R108 VTAIL.n5 VTAIL.n3 1.82809
R109 VTAIL.n2 VTAIL.n1 1.82809
R110 VTAIL VTAIL.n15 1.7699
R111 VTAIL.n11 VTAIL.n10 0.470328
R112 VTAIL.n3 VTAIL.n2 0.470328
R113 VTAIL VTAIL.n1 0.0586897
R114 VDD1 VDD1.n0 68.4057
R115 VDD1.n3 VDD1.n2 68.292
R116 VDD1.n3 VDD1.n1 68.292
R117 VDD1.n5 VDD1.n4 67.4336
R118 VDD1.n5 VDD1.n3 36.669
R119 VDD1.n4 VDD1.t2 4.11692
R120 VDD1.n4 VDD1.t3 4.11692
R121 VDD1.n0 VDD1.t5 4.11692
R122 VDD1.n0 VDD1.t1 4.11692
R123 VDD1.n2 VDD1.t0 4.11692
R124 VDD1.n2 VDD1.t7 4.11692
R125 VDD1.n1 VDD1.t4 4.11692
R126 VDD1.n1 VDD1.t6 4.11692
R127 VDD1 VDD1.n5 0.856103
R128 B.n403 B.n273 588.598
R129 B.n576 B.n72 588.598
R130 B.n299 B.n271 588.598
R131 B.n572 B.n99 588.598
R132 B.n572 B.n571 585
R133 B.n198 B.n98 585
R134 B.n197 B.n196 585
R135 B.n195 B.n194 585
R136 B.n193 B.n192 585
R137 B.n191 B.n190 585
R138 B.n189 B.n188 585
R139 B.n187 B.n186 585
R140 B.n185 B.n184 585
R141 B.n183 B.n182 585
R142 B.n181 B.n180 585
R143 B.n179 B.n178 585
R144 B.n177 B.n176 585
R145 B.n175 B.n174 585
R146 B.n173 B.n172 585
R147 B.n171 B.n170 585
R148 B.n169 B.n168 585
R149 B.n167 B.n166 585
R150 B.n165 B.n164 585
R151 B.n163 B.n162 585
R152 B.n161 B.n160 585
R153 B.n159 B.n158 585
R154 B.n157 B.n156 585
R155 B.n155 B.n154 585
R156 B.n153 B.n152 585
R157 B.n151 B.n150 585
R158 B.n149 B.n148 585
R159 B.n147 B.n146 585
R160 B.n145 B.n144 585
R161 B.n143 B.n142 585
R162 B.n141 B.n140 585
R163 B.n139 B.n138 585
R164 B.n137 B.n136 585
R165 B.n135 B.n134 585
R166 B.n133 B.n132 585
R167 B.n131 B.n130 585
R168 B.n129 B.n128 585
R169 B.n127 B.n126 585
R170 B.n125 B.n124 585
R171 B.n123 B.n122 585
R172 B.n121 B.n120 585
R173 B.n119 B.n118 585
R174 B.n117 B.n116 585
R175 B.n115 B.n114 585
R176 B.n113 B.n112 585
R177 B.n111 B.n110 585
R178 B.n109 B.n108 585
R179 B.n107 B.n106 585
R180 B.n74 B.n73 585
R181 B.n577 B.n576 585
R182 B.n570 B.n99 585
R183 B.n99 B.n71 585
R184 B.n569 B.n70 585
R185 B.n581 B.n70 585
R186 B.n568 B.n69 585
R187 B.n582 B.n69 585
R188 B.n567 B.n68 585
R189 B.n583 B.n68 585
R190 B.n566 B.n565 585
R191 B.n565 B.n64 585
R192 B.n564 B.n63 585
R193 B.n589 B.n63 585
R194 B.n563 B.n62 585
R195 B.n590 B.n62 585
R196 B.n562 B.n61 585
R197 B.n591 B.n61 585
R198 B.n561 B.n560 585
R199 B.n560 B.n57 585
R200 B.n559 B.n56 585
R201 B.n597 B.n56 585
R202 B.n558 B.n55 585
R203 B.n598 B.n55 585
R204 B.n557 B.n54 585
R205 B.n599 B.n54 585
R206 B.n556 B.n555 585
R207 B.n555 B.n50 585
R208 B.n554 B.n49 585
R209 B.n605 B.n49 585
R210 B.n553 B.n48 585
R211 B.n606 B.n48 585
R212 B.n552 B.n47 585
R213 B.n607 B.n47 585
R214 B.n551 B.n550 585
R215 B.n550 B.n43 585
R216 B.n549 B.n42 585
R217 B.n613 B.n42 585
R218 B.n548 B.n41 585
R219 B.n614 B.n41 585
R220 B.n547 B.n40 585
R221 B.n615 B.n40 585
R222 B.n546 B.n545 585
R223 B.n545 B.n36 585
R224 B.n544 B.n35 585
R225 B.n621 B.n35 585
R226 B.n543 B.n34 585
R227 B.n622 B.n34 585
R228 B.n542 B.n33 585
R229 B.n623 B.n33 585
R230 B.n541 B.n540 585
R231 B.n540 B.n29 585
R232 B.n539 B.n28 585
R233 B.n629 B.n28 585
R234 B.n538 B.n27 585
R235 B.n630 B.n27 585
R236 B.n537 B.n26 585
R237 B.n631 B.n26 585
R238 B.n536 B.n535 585
R239 B.n535 B.n25 585
R240 B.n534 B.n21 585
R241 B.n637 B.n21 585
R242 B.n533 B.n20 585
R243 B.n638 B.n20 585
R244 B.n532 B.n19 585
R245 B.n639 B.n19 585
R246 B.n531 B.n530 585
R247 B.n530 B.n15 585
R248 B.n529 B.n14 585
R249 B.n645 B.n14 585
R250 B.n528 B.n13 585
R251 B.n646 B.n13 585
R252 B.n527 B.n12 585
R253 B.n647 B.n12 585
R254 B.n526 B.n525 585
R255 B.n525 B.n8 585
R256 B.n524 B.n7 585
R257 B.n653 B.n7 585
R258 B.n523 B.n6 585
R259 B.n654 B.n6 585
R260 B.n522 B.n5 585
R261 B.n655 B.n5 585
R262 B.n521 B.n520 585
R263 B.n520 B.n4 585
R264 B.n519 B.n199 585
R265 B.n519 B.n518 585
R266 B.n509 B.n200 585
R267 B.n201 B.n200 585
R268 B.n511 B.n510 585
R269 B.n512 B.n511 585
R270 B.n508 B.n205 585
R271 B.n209 B.n205 585
R272 B.n507 B.n506 585
R273 B.n506 B.n505 585
R274 B.n207 B.n206 585
R275 B.n208 B.n207 585
R276 B.n498 B.n497 585
R277 B.n499 B.n498 585
R278 B.n496 B.n214 585
R279 B.n214 B.n213 585
R280 B.n495 B.n494 585
R281 B.n494 B.n493 585
R282 B.n216 B.n215 585
R283 B.n486 B.n216 585
R284 B.n485 B.n484 585
R285 B.n487 B.n485 585
R286 B.n483 B.n221 585
R287 B.n221 B.n220 585
R288 B.n482 B.n481 585
R289 B.n481 B.n480 585
R290 B.n223 B.n222 585
R291 B.n224 B.n223 585
R292 B.n473 B.n472 585
R293 B.n474 B.n473 585
R294 B.n471 B.n229 585
R295 B.n229 B.n228 585
R296 B.n470 B.n469 585
R297 B.n469 B.n468 585
R298 B.n231 B.n230 585
R299 B.n232 B.n231 585
R300 B.n461 B.n460 585
R301 B.n462 B.n461 585
R302 B.n459 B.n237 585
R303 B.n237 B.n236 585
R304 B.n458 B.n457 585
R305 B.n457 B.n456 585
R306 B.n239 B.n238 585
R307 B.n240 B.n239 585
R308 B.n449 B.n448 585
R309 B.n450 B.n449 585
R310 B.n447 B.n245 585
R311 B.n245 B.n244 585
R312 B.n446 B.n445 585
R313 B.n445 B.n444 585
R314 B.n247 B.n246 585
R315 B.n248 B.n247 585
R316 B.n437 B.n436 585
R317 B.n438 B.n437 585
R318 B.n435 B.n253 585
R319 B.n253 B.n252 585
R320 B.n434 B.n433 585
R321 B.n433 B.n432 585
R322 B.n255 B.n254 585
R323 B.n256 B.n255 585
R324 B.n425 B.n424 585
R325 B.n426 B.n425 585
R326 B.n423 B.n260 585
R327 B.n264 B.n260 585
R328 B.n422 B.n421 585
R329 B.n421 B.n420 585
R330 B.n262 B.n261 585
R331 B.n263 B.n262 585
R332 B.n413 B.n412 585
R333 B.n414 B.n413 585
R334 B.n411 B.n269 585
R335 B.n269 B.n268 585
R336 B.n410 B.n409 585
R337 B.n409 B.n408 585
R338 B.n271 B.n270 585
R339 B.n272 B.n271 585
R340 B.n404 B.n403 585
R341 B.n275 B.n274 585
R342 B.n400 B.n399 585
R343 B.n401 B.n400 585
R344 B.n398 B.n300 585
R345 B.n397 B.n396 585
R346 B.n395 B.n394 585
R347 B.n393 B.n392 585
R348 B.n391 B.n390 585
R349 B.n389 B.n388 585
R350 B.n387 B.n386 585
R351 B.n385 B.n384 585
R352 B.n383 B.n382 585
R353 B.n381 B.n380 585
R354 B.n379 B.n378 585
R355 B.n377 B.n376 585
R356 B.n375 B.n374 585
R357 B.n373 B.n372 585
R358 B.n371 B.n370 585
R359 B.n369 B.n368 585
R360 B.n367 B.n366 585
R361 B.n364 B.n363 585
R362 B.n362 B.n361 585
R363 B.n360 B.n359 585
R364 B.n358 B.n357 585
R365 B.n356 B.n355 585
R366 B.n354 B.n353 585
R367 B.n352 B.n351 585
R368 B.n350 B.n349 585
R369 B.n348 B.n347 585
R370 B.n346 B.n345 585
R371 B.n343 B.n342 585
R372 B.n341 B.n340 585
R373 B.n339 B.n338 585
R374 B.n337 B.n336 585
R375 B.n335 B.n334 585
R376 B.n333 B.n332 585
R377 B.n331 B.n330 585
R378 B.n329 B.n328 585
R379 B.n327 B.n326 585
R380 B.n325 B.n324 585
R381 B.n323 B.n322 585
R382 B.n321 B.n320 585
R383 B.n319 B.n318 585
R384 B.n317 B.n316 585
R385 B.n315 B.n314 585
R386 B.n313 B.n312 585
R387 B.n311 B.n310 585
R388 B.n309 B.n308 585
R389 B.n307 B.n306 585
R390 B.n305 B.n299 585
R391 B.n401 B.n299 585
R392 B.n405 B.n273 585
R393 B.n273 B.n272 585
R394 B.n407 B.n406 585
R395 B.n408 B.n407 585
R396 B.n267 B.n266 585
R397 B.n268 B.n267 585
R398 B.n416 B.n415 585
R399 B.n415 B.n414 585
R400 B.n417 B.n265 585
R401 B.n265 B.n263 585
R402 B.n419 B.n418 585
R403 B.n420 B.n419 585
R404 B.n259 B.n258 585
R405 B.n264 B.n259 585
R406 B.n428 B.n427 585
R407 B.n427 B.n426 585
R408 B.n429 B.n257 585
R409 B.n257 B.n256 585
R410 B.n431 B.n430 585
R411 B.n432 B.n431 585
R412 B.n251 B.n250 585
R413 B.n252 B.n251 585
R414 B.n440 B.n439 585
R415 B.n439 B.n438 585
R416 B.n441 B.n249 585
R417 B.n249 B.n248 585
R418 B.n443 B.n442 585
R419 B.n444 B.n443 585
R420 B.n243 B.n242 585
R421 B.n244 B.n243 585
R422 B.n452 B.n451 585
R423 B.n451 B.n450 585
R424 B.n453 B.n241 585
R425 B.n241 B.n240 585
R426 B.n455 B.n454 585
R427 B.n456 B.n455 585
R428 B.n235 B.n234 585
R429 B.n236 B.n235 585
R430 B.n464 B.n463 585
R431 B.n463 B.n462 585
R432 B.n465 B.n233 585
R433 B.n233 B.n232 585
R434 B.n467 B.n466 585
R435 B.n468 B.n467 585
R436 B.n227 B.n226 585
R437 B.n228 B.n227 585
R438 B.n476 B.n475 585
R439 B.n475 B.n474 585
R440 B.n477 B.n225 585
R441 B.n225 B.n224 585
R442 B.n479 B.n478 585
R443 B.n480 B.n479 585
R444 B.n219 B.n218 585
R445 B.n220 B.n219 585
R446 B.n489 B.n488 585
R447 B.n488 B.n487 585
R448 B.n490 B.n217 585
R449 B.n486 B.n217 585
R450 B.n492 B.n491 585
R451 B.n493 B.n492 585
R452 B.n212 B.n211 585
R453 B.n213 B.n212 585
R454 B.n501 B.n500 585
R455 B.n500 B.n499 585
R456 B.n502 B.n210 585
R457 B.n210 B.n208 585
R458 B.n504 B.n503 585
R459 B.n505 B.n504 585
R460 B.n204 B.n203 585
R461 B.n209 B.n204 585
R462 B.n514 B.n513 585
R463 B.n513 B.n512 585
R464 B.n515 B.n202 585
R465 B.n202 B.n201 585
R466 B.n517 B.n516 585
R467 B.n518 B.n517 585
R468 B.n2 B.n0 585
R469 B.n4 B.n2 585
R470 B.n3 B.n1 585
R471 B.n654 B.n3 585
R472 B.n652 B.n651 585
R473 B.n653 B.n652 585
R474 B.n650 B.n9 585
R475 B.n9 B.n8 585
R476 B.n649 B.n648 585
R477 B.n648 B.n647 585
R478 B.n11 B.n10 585
R479 B.n646 B.n11 585
R480 B.n644 B.n643 585
R481 B.n645 B.n644 585
R482 B.n642 B.n16 585
R483 B.n16 B.n15 585
R484 B.n641 B.n640 585
R485 B.n640 B.n639 585
R486 B.n18 B.n17 585
R487 B.n638 B.n18 585
R488 B.n636 B.n635 585
R489 B.n637 B.n636 585
R490 B.n634 B.n22 585
R491 B.n25 B.n22 585
R492 B.n633 B.n632 585
R493 B.n632 B.n631 585
R494 B.n24 B.n23 585
R495 B.n630 B.n24 585
R496 B.n628 B.n627 585
R497 B.n629 B.n628 585
R498 B.n626 B.n30 585
R499 B.n30 B.n29 585
R500 B.n625 B.n624 585
R501 B.n624 B.n623 585
R502 B.n32 B.n31 585
R503 B.n622 B.n32 585
R504 B.n620 B.n619 585
R505 B.n621 B.n620 585
R506 B.n618 B.n37 585
R507 B.n37 B.n36 585
R508 B.n617 B.n616 585
R509 B.n616 B.n615 585
R510 B.n39 B.n38 585
R511 B.n614 B.n39 585
R512 B.n612 B.n611 585
R513 B.n613 B.n612 585
R514 B.n610 B.n44 585
R515 B.n44 B.n43 585
R516 B.n609 B.n608 585
R517 B.n608 B.n607 585
R518 B.n46 B.n45 585
R519 B.n606 B.n46 585
R520 B.n604 B.n603 585
R521 B.n605 B.n604 585
R522 B.n602 B.n51 585
R523 B.n51 B.n50 585
R524 B.n601 B.n600 585
R525 B.n600 B.n599 585
R526 B.n53 B.n52 585
R527 B.n598 B.n53 585
R528 B.n596 B.n595 585
R529 B.n597 B.n596 585
R530 B.n594 B.n58 585
R531 B.n58 B.n57 585
R532 B.n593 B.n592 585
R533 B.n592 B.n591 585
R534 B.n60 B.n59 585
R535 B.n590 B.n60 585
R536 B.n588 B.n587 585
R537 B.n589 B.n588 585
R538 B.n586 B.n65 585
R539 B.n65 B.n64 585
R540 B.n585 B.n584 585
R541 B.n584 B.n583 585
R542 B.n67 B.n66 585
R543 B.n582 B.n67 585
R544 B.n580 B.n579 585
R545 B.n581 B.n580 585
R546 B.n578 B.n72 585
R547 B.n72 B.n71 585
R548 B.n657 B.n656 585
R549 B.n656 B.n655 585
R550 B.n303 B.t8 271.139
R551 B.n301 B.t19 271.139
R552 B.n103 B.t12 271.139
R553 B.n100 B.t16 271.139
R554 B.n574 B.n573 256.663
R555 B.n574 B.n97 256.663
R556 B.n574 B.n96 256.663
R557 B.n574 B.n95 256.663
R558 B.n574 B.n94 256.663
R559 B.n574 B.n93 256.663
R560 B.n574 B.n92 256.663
R561 B.n574 B.n91 256.663
R562 B.n574 B.n90 256.663
R563 B.n574 B.n89 256.663
R564 B.n574 B.n88 256.663
R565 B.n574 B.n87 256.663
R566 B.n574 B.n86 256.663
R567 B.n574 B.n85 256.663
R568 B.n574 B.n84 256.663
R569 B.n574 B.n83 256.663
R570 B.n574 B.n82 256.663
R571 B.n574 B.n81 256.663
R572 B.n574 B.n80 256.663
R573 B.n574 B.n79 256.663
R574 B.n574 B.n78 256.663
R575 B.n574 B.n77 256.663
R576 B.n574 B.n76 256.663
R577 B.n574 B.n75 256.663
R578 B.n575 B.n574 256.663
R579 B.n402 B.n401 256.663
R580 B.n401 B.n276 256.663
R581 B.n401 B.n277 256.663
R582 B.n401 B.n278 256.663
R583 B.n401 B.n279 256.663
R584 B.n401 B.n280 256.663
R585 B.n401 B.n281 256.663
R586 B.n401 B.n282 256.663
R587 B.n401 B.n283 256.663
R588 B.n401 B.n284 256.663
R589 B.n401 B.n285 256.663
R590 B.n401 B.n286 256.663
R591 B.n401 B.n287 256.663
R592 B.n401 B.n288 256.663
R593 B.n401 B.n289 256.663
R594 B.n401 B.n290 256.663
R595 B.n401 B.n291 256.663
R596 B.n401 B.n292 256.663
R597 B.n401 B.n293 256.663
R598 B.n401 B.n294 256.663
R599 B.n401 B.n295 256.663
R600 B.n401 B.n296 256.663
R601 B.n401 B.n297 256.663
R602 B.n401 B.n298 256.663
R603 B.n407 B.n273 163.367
R604 B.n407 B.n267 163.367
R605 B.n415 B.n267 163.367
R606 B.n415 B.n265 163.367
R607 B.n419 B.n265 163.367
R608 B.n419 B.n259 163.367
R609 B.n427 B.n259 163.367
R610 B.n427 B.n257 163.367
R611 B.n431 B.n257 163.367
R612 B.n431 B.n251 163.367
R613 B.n439 B.n251 163.367
R614 B.n439 B.n249 163.367
R615 B.n443 B.n249 163.367
R616 B.n443 B.n243 163.367
R617 B.n451 B.n243 163.367
R618 B.n451 B.n241 163.367
R619 B.n455 B.n241 163.367
R620 B.n455 B.n235 163.367
R621 B.n463 B.n235 163.367
R622 B.n463 B.n233 163.367
R623 B.n467 B.n233 163.367
R624 B.n467 B.n227 163.367
R625 B.n475 B.n227 163.367
R626 B.n475 B.n225 163.367
R627 B.n479 B.n225 163.367
R628 B.n479 B.n219 163.367
R629 B.n488 B.n219 163.367
R630 B.n488 B.n217 163.367
R631 B.n492 B.n217 163.367
R632 B.n492 B.n212 163.367
R633 B.n500 B.n212 163.367
R634 B.n500 B.n210 163.367
R635 B.n504 B.n210 163.367
R636 B.n504 B.n204 163.367
R637 B.n513 B.n204 163.367
R638 B.n513 B.n202 163.367
R639 B.n517 B.n202 163.367
R640 B.n517 B.n2 163.367
R641 B.n656 B.n2 163.367
R642 B.n656 B.n3 163.367
R643 B.n652 B.n3 163.367
R644 B.n652 B.n9 163.367
R645 B.n648 B.n9 163.367
R646 B.n648 B.n11 163.367
R647 B.n644 B.n11 163.367
R648 B.n644 B.n16 163.367
R649 B.n640 B.n16 163.367
R650 B.n640 B.n18 163.367
R651 B.n636 B.n18 163.367
R652 B.n636 B.n22 163.367
R653 B.n632 B.n22 163.367
R654 B.n632 B.n24 163.367
R655 B.n628 B.n24 163.367
R656 B.n628 B.n30 163.367
R657 B.n624 B.n30 163.367
R658 B.n624 B.n32 163.367
R659 B.n620 B.n32 163.367
R660 B.n620 B.n37 163.367
R661 B.n616 B.n37 163.367
R662 B.n616 B.n39 163.367
R663 B.n612 B.n39 163.367
R664 B.n612 B.n44 163.367
R665 B.n608 B.n44 163.367
R666 B.n608 B.n46 163.367
R667 B.n604 B.n46 163.367
R668 B.n604 B.n51 163.367
R669 B.n600 B.n51 163.367
R670 B.n600 B.n53 163.367
R671 B.n596 B.n53 163.367
R672 B.n596 B.n58 163.367
R673 B.n592 B.n58 163.367
R674 B.n592 B.n60 163.367
R675 B.n588 B.n60 163.367
R676 B.n588 B.n65 163.367
R677 B.n584 B.n65 163.367
R678 B.n584 B.n67 163.367
R679 B.n580 B.n67 163.367
R680 B.n580 B.n72 163.367
R681 B.n400 B.n275 163.367
R682 B.n400 B.n300 163.367
R683 B.n396 B.n395 163.367
R684 B.n392 B.n391 163.367
R685 B.n388 B.n387 163.367
R686 B.n384 B.n383 163.367
R687 B.n380 B.n379 163.367
R688 B.n376 B.n375 163.367
R689 B.n372 B.n371 163.367
R690 B.n368 B.n367 163.367
R691 B.n363 B.n362 163.367
R692 B.n359 B.n358 163.367
R693 B.n355 B.n354 163.367
R694 B.n351 B.n350 163.367
R695 B.n347 B.n346 163.367
R696 B.n342 B.n341 163.367
R697 B.n338 B.n337 163.367
R698 B.n334 B.n333 163.367
R699 B.n330 B.n329 163.367
R700 B.n326 B.n325 163.367
R701 B.n322 B.n321 163.367
R702 B.n318 B.n317 163.367
R703 B.n314 B.n313 163.367
R704 B.n310 B.n309 163.367
R705 B.n306 B.n299 163.367
R706 B.n409 B.n271 163.367
R707 B.n409 B.n269 163.367
R708 B.n413 B.n269 163.367
R709 B.n413 B.n262 163.367
R710 B.n421 B.n262 163.367
R711 B.n421 B.n260 163.367
R712 B.n425 B.n260 163.367
R713 B.n425 B.n255 163.367
R714 B.n433 B.n255 163.367
R715 B.n433 B.n253 163.367
R716 B.n437 B.n253 163.367
R717 B.n437 B.n247 163.367
R718 B.n445 B.n247 163.367
R719 B.n445 B.n245 163.367
R720 B.n449 B.n245 163.367
R721 B.n449 B.n239 163.367
R722 B.n457 B.n239 163.367
R723 B.n457 B.n237 163.367
R724 B.n461 B.n237 163.367
R725 B.n461 B.n231 163.367
R726 B.n469 B.n231 163.367
R727 B.n469 B.n229 163.367
R728 B.n473 B.n229 163.367
R729 B.n473 B.n223 163.367
R730 B.n481 B.n223 163.367
R731 B.n481 B.n221 163.367
R732 B.n485 B.n221 163.367
R733 B.n485 B.n216 163.367
R734 B.n494 B.n216 163.367
R735 B.n494 B.n214 163.367
R736 B.n498 B.n214 163.367
R737 B.n498 B.n207 163.367
R738 B.n506 B.n207 163.367
R739 B.n506 B.n205 163.367
R740 B.n511 B.n205 163.367
R741 B.n511 B.n200 163.367
R742 B.n519 B.n200 163.367
R743 B.n520 B.n519 163.367
R744 B.n520 B.n5 163.367
R745 B.n6 B.n5 163.367
R746 B.n7 B.n6 163.367
R747 B.n525 B.n7 163.367
R748 B.n525 B.n12 163.367
R749 B.n13 B.n12 163.367
R750 B.n14 B.n13 163.367
R751 B.n530 B.n14 163.367
R752 B.n530 B.n19 163.367
R753 B.n20 B.n19 163.367
R754 B.n21 B.n20 163.367
R755 B.n535 B.n21 163.367
R756 B.n535 B.n26 163.367
R757 B.n27 B.n26 163.367
R758 B.n28 B.n27 163.367
R759 B.n540 B.n28 163.367
R760 B.n540 B.n33 163.367
R761 B.n34 B.n33 163.367
R762 B.n35 B.n34 163.367
R763 B.n545 B.n35 163.367
R764 B.n545 B.n40 163.367
R765 B.n41 B.n40 163.367
R766 B.n42 B.n41 163.367
R767 B.n550 B.n42 163.367
R768 B.n550 B.n47 163.367
R769 B.n48 B.n47 163.367
R770 B.n49 B.n48 163.367
R771 B.n555 B.n49 163.367
R772 B.n555 B.n54 163.367
R773 B.n55 B.n54 163.367
R774 B.n56 B.n55 163.367
R775 B.n560 B.n56 163.367
R776 B.n560 B.n61 163.367
R777 B.n62 B.n61 163.367
R778 B.n63 B.n62 163.367
R779 B.n565 B.n63 163.367
R780 B.n565 B.n68 163.367
R781 B.n69 B.n68 163.367
R782 B.n70 B.n69 163.367
R783 B.n99 B.n70 163.367
R784 B.n106 B.n74 163.367
R785 B.n110 B.n109 163.367
R786 B.n114 B.n113 163.367
R787 B.n118 B.n117 163.367
R788 B.n122 B.n121 163.367
R789 B.n126 B.n125 163.367
R790 B.n130 B.n129 163.367
R791 B.n134 B.n133 163.367
R792 B.n138 B.n137 163.367
R793 B.n142 B.n141 163.367
R794 B.n146 B.n145 163.367
R795 B.n150 B.n149 163.367
R796 B.n154 B.n153 163.367
R797 B.n158 B.n157 163.367
R798 B.n162 B.n161 163.367
R799 B.n166 B.n165 163.367
R800 B.n170 B.n169 163.367
R801 B.n174 B.n173 163.367
R802 B.n178 B.n177 163.367
R803 B.n182 B.n181 163.367
R804 B.n186 B.n185 163.367
R805 B.n190 B.n189 163.367
R806 B.n194 B.n193 163.367
R807 B.n196 B.n98 163.367
R808 B.n401 B.n272 155.975
R809 B.n574 B.n71 155.975
R810 B.n303 B.t11 112.43
R811 B.n100 B.t17 112.43
R812 B.n301 B.t21 112.424
R813 B.n103 B.t14 112.424
R814 B.n408 B.n272 74.1701
R815 B.n408 B.n268 74.1701
R816 B.n414 B.n268 74.1701
R817 B.n414 B.n263 74.1701
R818 B.n420 B.n263 74.1701
R819 B.n420 B.n264 74.1701
R820 B.n426 B.n256 74.1701
R821 B.n432 B.n256 74.1701
R822 B.n432 B.n252 74.1701
R823 B.n438 B.n252 74.1701
R824 B.n438 B.n248 74.1701
R825 B.n444 B.n248 74.1701
R826 B.n444 B.n244 74.1701
R827 B.n450 B.n244 74.1701
R828 B.n456 B.n240 74.1701
R829 B.n456 B.n236 74.1701
R830 B.n462 B.n236 74.1701
R831 B.n462 B.n232 74.1701
R832 B.n468 B.n232 74.1701
R833 B.n474 B.n228 74.1701
R834 B.n474 B.n224 74.1701
R835 B.n480 B.n224 74.1701
R836 B.n480 B.n220 74.1701
R837 B.n487 B.n220 74.1701
R838 B.n487 B.n486 74.1701
R839 B.n493 B.n213 74.1701
R840 B.n499 B.n213 74.1701
R841 B.n499 B.n208 74.1701
R842 B.n505 B.n208 74.1701
R843 B.n505 B.n209 74.1701
R844 B.n512 B.n201 74.1701
R845 B.n518 B.n201 74.1701
R846 B.n518 B.n4 74.1701
R847 B.n655 B.n4 74.1701
R848 B.n655 B.n654 74.1701
R849 B.n654 B.n653 74.1701
R850 B.n653 B.n8 74.1701
R851 B.n647 B.n8 74.1701
R852 B.n646 B.n645 74.1701
R853 B.n645 B.n15 74.1701
R854 B.n639 B.n15 74.1701
R855 B.n639 B.n638 74.1701
R856 B.n638 B.n637 74.1701
R857 B.n631 B.n25 74.1701
R858 B.n631 B.n630 74.1701
R859 B.n630 B.n629 74.1701
R860 B.n629 B.n29 74.1701
R861 B.n623 B.n29 74.1701
R862 B.n623 B.n622 74.1701
R863 B.n621 B.n36 74.1701
R864 B.n615 B.n36 74.1701
R865 B.n615 B.n614 74.1701
R866 B.n614 B.n613 74.1701
R867 B.n613 B.n43 74.1701
R868 B.n607 B.n606 74.1701
R869 B.n606 B.n605 74.1701
R870 B.n605 B.n50 74.1701
R871 B.n599 B.n50 74.1701
R872 B.n599 B.n598 74.1701
R873 B.n598 B.n597 74.1701
R874 B.n597 B.n57 74.1701
R875 B.n591 B.n57 74.1701
R876 B.n590 B.n589 74.1701
R877 B.n589 B.n64 74.1701
R878 B.n583 B.n64 74.1701
R879 B.n583 B.n582 74.1701
R880 B.n582 B.n581 74.1701
R881 B.n581 B.n71 74.1701
R882 B.n403 B.n402 71.676
R883 B.n300 B.n276 71.676
R884 B.n395 B.n277 71.676
R885 B.n391 B.n278 71.676
R886 B.n387 B.n279 71.676
R887 B.n383 B.n280 71.676
R888 B.n379 B.n281 71.676
R889 B.n375 B.n282 71.676
R890 B.n371 B.n283 71.676
R891 B.n367 B.n284 71.676
R892 B.n362 B.n285 71.676
R893 B.n358 B.n286 71.676
R894 B.n354 B.n287 71.676
R895 B.n350 B.n288 71.676
R896 B.n346 B.n289 71.676
R897 B.n341 B.n290 71.676
R898 B.n337 B.n291 71.676
R899 B.n333 B.n292 71.676
R900 B.n329 B.n293 71.676
R901 B.n325 B.n294 71.676
R902 B.n321 B.n295 71.676
R903 B.n317 B.n296 71.676
R904 B.n313 B.n297 71.676
R905 B.n309 B.n298 71.676
R906 B.n576 B.n575 71.676
R907 B.n106 B.n75 71.676
R908 B.n110 B.n76 71.676
R909 B.n114 B.n77 71.676
R910 B.n118 B.n78 71.676
R911 B.n122 B.n79 71.676
R912 B.n126 B.n80 71.676
R913 B.n130 B.n81 71.676
R914 B.n134 B.n82 71.676
R915 B.n138 B.n83 71.676
R916 B.n142 B.n84 71.676
R917 B.n146 B.n85 71.676
R918 B.n150 B.n86 71.676
R919 B.n154 B.n87 71.676
R920 B.n158 B.n88 71.676
R921 B.n162 B.n89 71.676
R922 B.n166 B.n90 71.676
R923 B.n170 B.n91 71.676
R924 B.n174 B.n92 71.676
R925 B.n178 B.n93 71.676
R926 B.n182 B.n94 71.676
R927 B.n186 B.n95 71.676
R928 B.n190 B.n96 71.676
R929 B.n194 B.n97 71.676
R930 B.n573 B.n98 71.676
R931 B.n573 B.n572 71.676
R932 B.n196 B.n97 71.676
R933 B.n193 B.n96 71.676
R934 B.n189 B.n95 71.676
R935 B.n185 B.n94 71.676
R936 B.n181 B.n93 71.676
R937 B.n177 B.n92 71.676
R938 B.n173 B.n91 71.676
R939 B.n169 B.n90 71.676
R940 B.n165 B.n89 71.676
R941 B.n161 B.n88 71.676
R942 B.n157 B.n87 71.676
R943 B.n153 B.n86 71.676
R944 B.n149 B.n85 71.676
R945 B.n145 B.n84 71.676
R946 B.n141 B.n83 71.676
R947 B.n137 B.n82 71.676
R948 B.n133 B.n81 71.676
R949 B.n129 B.n80 71.676
R950 B.n125 B.n79 71.676
R951 B.n121 B.n78 71.676
R952 B.n117 B.n77 71.676
R953 B.n113 B.n76 71.676
R954 B.n109 B.n75 71.676
R955 B.n575 B.n74 71.676
R956 B.n402 B.n275 71.676
R957 B.n396 B.n276 71.676
R958 B.n392 B.n277 71.676
R959 B.n388 B.n278 71.676
R960 B.n384 B.n279 71.676
R961 B.n380 B.n280 71.676
R962 B.n376 B.n281 71.676
R963 B.n372 B.n282 71.676
R964 B.n368 B.n283 71.676
R965 B.n363 B.n284 71.676
R966 B.n359 B.n285 71.676
R967 B.n355 B.n286 71.676
R968 B.n351 B.n287 71.676
R969 B.n347 B.n288 71.676
R970 B.n342 B.n289 71.676
R971 B.n338 B.n290 71.676
R972 B.n334 B.n291 71.676
R973 B.n330 B.n292 71.676
R974 B.n326 B.n293 71.676
R975 B.n322 B.n294 71.676
R976 B.n318 B.n295 71.676
R977 B.n314 B.n296 71.676
R978 B.n310 B.n297 71.676
R979 B.n306 B.n298 71.676
R980 B.n304 B.t10 71.314
R981 B.n101 B.t18 71.314
R982 B.n302 B.t20 71.3092
R983 B.n104 B.t15 71.3092
R984 B.n493 B.t0 70.8979
R985 B.n637 B.t1 70.8979
R986 B.n426 B.t9 64.3535
R987 B.n591 B.t13 64.3535
R988 B.n468 B.t6 59.9906
R989 B.t2 B.n621 59.9906
R990 B.n344 B.n304 59.5399
R991 B.n365 B.n302 59.5399
R992 B.n105 B.n104 59.5399
R993 B.n102 B.n101 59.5399
R994 B.n512 B.t7 53.4462
R995 B.n647 B.t5 53.4462
R996 B.n450 B.t4 42.5389
R997 B.n607 B.t3 42.5389
R998 B.n304 B.n303 41.1157
R999 B.n302 B.n301 41.1157
R1000 B.n104 B.n103 41.1157
R1001 B.n101 B.n100 41.1157
R1002 B.n578 B.n577 38.2444
R1003 B.n571 B.n570 38.2444
R1004 B.n305 B.n270 38.2444
R1005 B.n405 B.n404 38.2444
R1006 B.t4 B.n240 31.6316
R1007 B.t3 B.n43 31.6316
R1008 B.n209 B.t7 20.7243
R1009 B.t5 B.n646 20.7243
R1010 B B.n657 18.0485
R1011 B.t6 B.n228 14.18
R1012 B.n622 B.t2 14.18
R1013 B.n577 B.n73 10.6151
R1014 B.n107 B.n73 10.6151
R1015 B.n108 B.n107 10.6151
R1016 B.n111 B.n108 10.6151
R1017 B.n112 B.n111 10.6151
R1018 B.n115 B.n112 10.6151
R1019 B.n116 B.n115 10.6151
R1020 B.n119 B.n116 10.6151
R1021 B.n120 B.n119 10.6151
R1022 B.n123 B.n120 10.6151
R1023 B.n124 B.n123 10.6151
R1024 B.n127 B.n124 10.6151
R1025 B.n128 B.n127 10.6151
R1026 B.n131 B.n128 10.6151
R1027 B.n132 B.n131 10.6151
R1028 B.n135 B.n132 10.6151
R1029 B.n136 B.n135 10.6151
R1030 B.n139 B.n136 10.6151
R1031 B.n140 B.n139 10.6151
R1032 B.n144 B.n143 10.6151
R1033 B.n147 B.n144 10.6151
R1034 B.n148 B.n147 10.6151
R1035 B.n151 B.n148 10.6151
R1036 B.n152 B.n151 10.6151
R1037 B.n155 B.n152 10.6151
R1038 B.n156 B.n155 10.6151
R1039 B.n159 B.n156 10.6151
R1040 B.n160 B.n159 10.6151
R1041 B.n164 B.n163 10.6151
R1042 B.n167 B.n164 10.6151
R1043 B.n168 B.n167 10.6151
R1044 B.n171 B.n168 10.6151
R1045 B.n172 B.n171 10.6151
R1046 B.n175 B.n172 10.6151
R1047 B.n176 B.n175 10.6151
R1048 B.n179 B.n176 10.6151
R1049 B.n180 B.n179 10.6151
R1050 B.n183 B.n180 10.6151
R1051 B.n184 B.n183 10.6151
R1052 B.n187 B.n184 10.6151
R1053 B.n188 B.n187 10.6151
R1054 B.n191 B.n188 10.6151
R1055 B.n192 B.n191 10.6151
R1056 B.n195 B.n192 10.6151
R1057 B.n197 B.n195 10.6151
R1058 B.n198 B.n197 10.6151
R1059 B.n571 B.n198 10.6151
R1060 B.n410 B.n270 10.6151
R1061 B.n411 B.n410 10.6151
R1062 B.n412 B.n411 10.6151
R1063 B.n412 B.n261 10.6151
R1064 B.n422 B.n261 10.6151
R1065 B.n423 B.n422 10.6151
R1066 B.n424 B.n423 10.6151
R1067 B.n424 B.n254 10.6151
R1068 B.n434 B.n254 10.6151
R1069 B.n435 B.n434 10.6151
R1070 B.n436 B.n435 10.6151
R1071 B.n436 B.n246 10.6151
R1072 B.n446 B.n246 10.6151
R1073 B.n447 B.n446 10.6151
R1074 B.n448 B.n447 10.6151
R1075 B.n448 B.n238 10.6151
R1076 B.n458 B.n238 10.6151
R1077 B.n459 B.n458 10.6151
R1078 B.n460 B.n459 10.6151
R1079 B.n460 B.n230 10.6151
R1080 B.n470 B.n230 10.6151
R1081 B.n471 B.n470 10.6151
R1082 B.n472 B.n471 10.6151
R1083 B.n472 B.n222 10.6151
R1084 B.n482 B.n222 10.6151
R1085 B.n483 B.n482 10.6151
R1086 B.n484 B.n483 10.6151
R1087 B.n484 B.n215 10.6151
R1088 B.n495 B.n215 10.6151
R1089 B.n496 B.n495 10.6151
R1090 B.n497 B.n496 10.6151
R1091 B.n497 B.n206 10.6151
R1092 B.n507 B.n206 10.6151
R1093 B.n508 B.n507 10.6151
R1094 B.n510 B.n508 10.6151
R1095 B.n510 B.n509 10.6151
R1096 B.n509 B.n199 10.6151
R1097 B.n521 B.n199 10.6151
R1098 B.n522 B.n521 10.6151
R1099 B.n523 B.n522 10.6151
R1100 B.n524 B.n523 10.6151
R1101 B.n526 B.n524 10.6151
R1102 B.n527 B.n526 10.6151
R1103 B.n528 B.n527 10.6151
R1104 B.n529 B.n528 10.6151
R1105 B.n531 B.n529 10.6151
R1106 B.n532 B.n531 10.6151
R1107 B.n533 B.n532 10.6151
R1108 B.n534 B.n533 10.6151
R1109 B.n536 B.n534 10.6151
R1110 B.n537 B.n536 10.6151
R1111 B.n538 B.n537 10.6151
R1112 B.n539 B.n538 10.6151
R1113 B.n541 B.n539 10.6151
R1114 B.n542 B.n541 10.6151
R1115 B.n543 B.n542 10.6151
R1116 B.n544 B.n543 10.6151
R1117 B.n546 B.n544 10.6151
R1118 B.n547 B.n546 10.6151
R1119 B.n548 B.n547 10.6151
R1120 B.n549 B.n548 10.6151
R1121 B.n551 B.n549 10.6151
R1122 B.n552 B.n551 10.6151
R1123 B.n553 B.n552 10.6151
R1124 B.n554 B.n553 10.6151
R1125 B.n556 B.n554 10.6151
R1126 B.n557 B.n556 10.6151
R1127 B.n558 B.n557 10.6151
R1128 B.n559 B.n558 10.6151
R1129 B.n561 B.n559 10.6151
R1130 B.n562 B.n561 10.6151
R1131 B.n563 B.n562 10.6151
R1132 B.n564 B.n563 10.6151
R1133 B.n566 B.n564 10.6151
R1134 B.n567 B.n566 10.6151
R1135 B.n568 B.n567 10.6151
R1136 B.n569 B.n568 10.6151
R1137 B.n570 B.n569 10.6151
R1138 B.n404 B.n274 10.6151
R1139 B.n399 B.n274 10.6151
R1140 B.n399 B.n398 10.6151
R1141 B.n398 B.n397 10.6151
R1142 B.n397 B.n394 10.6151
R1143 B.n394 B.n393 10.6151
R1144 B.n393 B.n390 10.6151
R1145 B.n390 B.n389 10.6151
R1146 B.n389 B.n386 10.6151
R1147 B.n386 B.n385 10.6151
R1148 B.n385 B.n382 10.6151
R1149 B.n382 B.n381 10.6151
R1150 B.n381 B.n378 10.6151
R1151 B.n378 B.n377 10.6151
R1152 B.n377 B.n374 10.6151
R1153 B.n374 B.n373 10.6151
R1154 B.n373 B.n370 10.6151
R1155 B.n370 B.n369 10.6151
R1156 B.n369 B.n366 10.6151
R1157 B.n364 B.n361 10.6151
R1158 B.n361 B.n360 10.6151
R1159 B.n360 B.n357 10.6151
R1160 B.n357 B.n356 10.6151
R1161 B.n356 B.n353 10.6151
R1162 B.n353 B.n352 10.6151
R1163 B.n352 B.n349 10.6151
R1164 B.n349 B.n348 10.6151
R1165 B.n348 B.n345 10.6151
R1166 B.n343 B.n340 10.6151
R1167 B.n340 B.n339 10.6151
R1168 B.n339 B.n336 10.6151
R1169 B.n336 B.n335 10.6151
R1170 B.n335 B.n332 10.6151
R1171 B.n332 B.n331 10.6151
R1172 B.n331 B.n328 10.6151
R1173 B.n328 B.n327 10.6151
R1174 B.n327 B.n324 10.6151
R1175 B.n324 B.n323 10.6151
R1176 B.n323 B.n320 10.6151
R1177 B.n320 B.n319 10.6151
R1178 B.n319 B.n316 10.6151
R1179 B.n316 B.n315 10.6151
R1180 B.n315 B.n312 10.6151
R1181 B.n312 B.n311 10.6151
R1182 B.n311 B.n308 10.6151
R1183 B.n308 B.n307 10.6151
R1184 B.n307 B.n305 10.6151
R1185 B.n406 B.n405 10.6151
R1186 B.n406 B.n266 10.6151
R1187 B.n416 B.n266 10.6151
R1188 B.n417 B.n416 10.6151
R1189 B.n418 B.n417 10.6151
R1190 B.n418 B.n258 10.6151
R1191 B.n428 B.n258 10.6151
R1192 B.n429 B.n428 10.6151
R1193 B.n430 B.n429 10.6151
R1194 B.n430 B.n250 10.6151
R1195 B.n440 B.n250 10.6151
R1196 B.n441 B.n440 10.6151
R1197 B.n442 B.n441 10.6151
R1198 B.n442 B.n242 10.6151
R1199 B.n452 B.n242 10.6151
R1200 B.n453 B.n452 10.6151
R1201 B.n454 B.n453 10.6151
R1202 B.n454 B.n234 10.6151
R1203 B.n464 B.n234 10.6151
R1204 B.n465 B.n464 10.6151
R1205 B.n466 B.n465 10.6151
R1206 B.n466 B.n226 10.6151
R1207 B.n476 B.n226 10.6151
R1208 B.n477 B.n476 10.6151
R1209 B.n478 B.n477 10.6151
R1210 B.n478 B.n218 10.6151
R1211 B.n489 B.n218 10.6151
R1212 B.n490 B.n489 10.6151
R1213 B.n491 B.n490 10.6151
R1214 B.n491 B.n211 10.6151
R1215 B.n501 B.n211 10.6151
R1216 B.n502 B.n501 10.6151
R1217 B.n503 B.n502 10.6151
R1218 B.n503 B.n203 10.6151
R1219 B.n514 B.n203 10.6151
R1220 B.n515 B.n514 10.6151
R1221 B.n516 B.n515 10.6151
R1222 B.n516 B.n0 10.6151
R1223 B.n651 B.n1 10.6151
R1224 B.n651 B.n650 10.6151
R1225 B.n650 B.n649 10.6151
R1226 B.n649 B.n10 10.6151
R1227 B.n643 B.n10 10.6151
R1228 B.n643 B.n642 10.6151
R1229 B.n642 B.n641 10.6151
R1230 B.n641 B.n17 10.6151
R1231 B.n635 B.n17 10.6151
R1232 B.n635 B.n634 10.6151
R1233 B.n634 B.n633 10.6151
R1234 B.n633 B.n23 10.6151
R1235 B.n627 B.n23 10.6151
R1236 B.n627 B.n626 10.6151
R1237 B.n626 B.n625 10.6151
R1238 B.n625 B.n31 10.6151
R1239 B.n619 B.n31 10.6151
R1240 B.n619 B.n618 10.6151
R1241 B.n618 B.n617 10.6151
R1242 B.n617 B.n38 10.6151
R1243 B.n611 B.n38 10.6151
R1244 B.n611 B.n610 10.6151
R1245 B.n610 B.n609 10.6151
R1246 B.n609 B.n45 10.6151
R1247 B.n603 B.n45 10.6151
R1248 B.n603 B.n602 10.6151
R1249 B.n602 B.n601 10.6151
R1250 B.n601 B.n52 10.6151
R1251 B.n595 B.n52 10.6151
R1252 B.n595 B.n594 10.6151
R1253 B.n594 B.n593 10.6151
R1254 B.n593 B.n59 10.6151
R1255 B.n587 B.n59 10.6151
R1256 B.n587 B.n586 10.6151
R1257 B.n586 B.n585 10.6151
R1258 B.n585 B.n66 10.6151
R1259 B.n579 B.n66 10.6151
R1260 B.n579 B.n578 10.6151
R1261 B.n264 B.t9 9.81706
R1262 B.t13 B.n590 9.81706
R1263 B.n140 B.n105 9.36635
R1264 B.n163 B.n102 9.36635
R1265 B.n366 B.n365 9.36635
R1266 B.n344 B.n343 9.36635
R1267 B.n486 B.t0 3.27269
R1268 B.n25 B.t1 3.27269
R1269 B.n657 B.n0 2.81026
R1270 B.n657 B.n1 2.81026
R1271 B.n143 B.n105 1.24928
R1272 B.n160 B.n102 1.24928
R1273 B.n365 B.n364 1.24928
R1274 B.n345 B.n344 1.24928
R1275 VN.n39 VN.n21 161.3
R1276 VN.n38 VN.n37 161.3
R1277 VN.n36 VN.n22 161.3
R1278 VN.n35 VN.n34 161.3
R1279 VN.n32 VN.n23 161.3
R1280 VN.n31 VN.n30 161.3
R1281 VN.n29 VN.n24 161.3
R1282 VN.n28 VN.n27 161.3
R1283 VN.n18 VN.n0 161.3
R1284 VN.n17 VN.n16 161.3
R1285 VN.n15 VN.n1 161.3
R1286 VN.n14 VN.n13 161.3
R1287 VN.n11 VN.n2 161.3
R1288 VN.n10 VN.n9 161.3
R1289 VN.n8 VN.n3 161.3
R1290 VN.n7 VN.n6 161.3
R1291 VN.n4 VN.t2 95.6032
R1292 VN.n25 VN.t5 95.6032
R1293 VN.n20 VN.n19 89.7148
R1294 VN.n41 VN.n40 89.7148
R1295 VN.n5 VN.t3 64.7608
R1296 VN.n12 VN.t1 64.7608
R1297 VN.n19 VN.t0 64.7608
R1298 VN.n26 VN.t6 64.7608
R1299 VN.n33 VN.t4 64.7608
R1300 VN.n40 VN.t7 64.7608
R1301 VN.n10 VN.n3 56.5193
R1302 VN.n31 VN.n24 56.5193
R1303 VN.n5 VN.n4 54.5414
R1304 VN.n26 VN.n25 54.5414
R1305 VN.n17 VN.n1 53.1199
R1306 VN.n38 VN.n22 53.1199
R1307 VN VN.n41 41.93
R1308 VN.n18 VN.n17 27.8669
R1309 VN.n39 VN.n38 27.8669
R1310 VN.n6 VN.n3 24.4675
R1311 VN.n11 VN.n10 24.4675
R1312 VN.n13 VN.n1 24.4675
R1313 VN.n27 VN.n24 24.4675
R1314 VN.n34 VN.n22 24.4675
R1315 VN.n32 VN.n31 24.4675
R1316 VN.n19 VN.n18 21.0421
R1317 VN.n40 VN.n39 21.0421
R1318 VN.n6 VN.n5 15.17
R1319 VN.n12 VN.n11 15.17
R1320 VN.n27 VN.n26 15.17
R1321 VN.n33 VN.n32 15.17
R1322 VN.n28 VN.n25 13.1161
R1323 VN.n7 VN.n4 13.1161
R1324 VN.n13 VN.n12 9.29796
R1325 VN.n34 VN.n33 9.29796
R1326 VN.n41 VN.n21 0.278367
R1327 VN.n20 VN.n0 0.278367
R1328 VN.n37 VN.n21 0.189894
R1329 VN.n37 VN.n36 0.189894
R1330 VN.n36 VN.n35 0.189894
R1331 VN.n35 VN.n23 0.189894
R1332 VN.n30 VN.n23 0.189894
R1333 VN.n30 VN.n29 0.189894
R1334 VN.n29 VN.n28 0.189894
R1335 VN.n8 VN.n7 0.189894
R1336 VN.n9 VN.n8 0.189894
R1337 VN.n9 VN.n2 0.189894
R1338 VN.n14 VN.n2 0.189894
R1339 VN.n15 VN.n14 0.189894
R1340 VN.n16 VN.n15 0.189894
R1341 VN.n16 VN.n0 0.189894
R1342 VN VN.n20 0.153454
R1343 VDD2.n2 VDD2.n1 68.292
R1344 VDD2.n2 VDD2.n0 68.292
R1345 VDD2 VDD2.n5 68.2892
R1346 VDD2.n4 VDD2.n3 67.4337
R1347 VDD2.n4 VDD2.n2 36.086
R1348 VDD2.n5 VDD2.t1 4.11692
R1349 VDD2.n5 VDD2.t2 4.11692
R1350 VDD2.n3 VDD2.t0 4.11692
R1351 VDD2.n3 VDD2.t3 4.11692
R1352 VDD2.n1 VDD2.t6 4.11692
R1353 VDD2.n1 VDD2.t7 4.11692
R1354 VDD2.n0 VDD2.t5 4.11692
R1355 VDD2.n0 VDD2.t4 4.11692
R1356 VDD2 VDD2.n4 0.972483
C0 VN VDD1 0.154051f
C1 VP VDD2 0.437713f
C2 VP VN 5.34463f
C3 VDD2 VTAIL 5.2618f
C4 VN VTAIL 4.02142f
C5 VP VDD1 3.7336f
C6 VDD1 VTAIL 5.21282f
C7 VN VDD2 3.45148f
C8 VP VTAIL 4.03553f
C9 VDD1 VDD2 1.35554f
C10 VDD2 B 4.00279f
C11 VDD1 B 4.348683f
C12 VTAIL B 5.372451f
C13 VN B 11.701509f
C14 VP B 10.28044f
C15 VDD2.t5 B 0.094201f
C16 VDD2.t4 B 0.094201f
C17 VDD2.n0 B 0.767911f
C18 VDD2.t6 B 0.094201f
C19 VDD2.t7 B 0.094201f
C20 VDD2.n1 B 0.767911f
C21 VDD2.n2 B 2.33705f
C22 VDD2.t0 B 0.094201f
C23 VDD2.t3 B 0.094201f
C24 VDD2.n3 B 0.762609f
C25 VDD2.n4 B 2.08131f
C26 VDD2.t1 B 0.094201f
C27 VDD2.t2 B 0.094201f
C28 VDD2.n5 B 0.767881f
C29 VN.n0 B 0.040851f
C30 VN.t0 B 0.695835f
C31 VN.n1 B 0.054978f
C32 VN.n2 B 0.030985f
C33 VN.t1 B 0.695835f
C34 VN.n3 B 0.045233f
C35 VN.t2 B 0.830702f
C36 VN.n4 B 0.348402f
C37 VN.t3 B 0.695835f
C38 VN.n5 B 0.349612f
C39 VN.n6 B 0.046915f
C40 VN.n7 B 0.226163f
C41 VN.n8 B 0.030985f
C42 VN.n9 B 0.030985f
C43 VN.n10 B 0.045233f
C44 VN.n11 B 0.046915f
C45 VN.n12 B 0.277727f
C46 VN.n13 B 0.040072f
C47 VN.n14 B 0.030985f
C48 VN.n15 B 0.030985f
C49 VN.n16 B 0.030985f
C50 VN.n17 B 0.032499f
C51 VN.n18 B 0.056747f
C52 VN.n19 B 0.365059f
C53 VN.n20 B 0.035534f
C54 VN.n21 B 0.040851f
C55 VN.t7 B 0.695835f
C56 VN.n22 B 0.054978f
C57 VN.n23 B 0.030985f
C58 VN.t4 B 0.695835f
C59 VN.n24 B 0.045233f
C60 VN.t5 B 0.830702f
C61 VN.n25 B 0.348402f
C62 VN.t6 B 0.695835f
C63 VN.n26 B 0.349612f
C64 VN.n27 B 0.046915f
C65 VN.n28 B 0.226163f
C66 VN.n29 B 0.030985f
C67 VN.n30 B 0.030985f
C68 VN.n31 B 0.045233f
C69 VN.n32 B 0.046915f
C70 VN.n33 B 0.277727f
C71 VN.n34 B 0.040072f
C72 VN.n35 B 0.030985f
C73 VN.n36 B 0.030985f
C74 VN.n37 B 0.030985f
C75 VN.n38 B 0.032499f
C76 VN.n39 B 0.056747f
C77 VN.n40 B 0.365059f
C78 VN.n41 B 1.30151f
C79 VDD1.t5 B 0.094291f
C80 VDD1.t1 B 0.094291f
C81 VDD1.n0 B 0.769456f
C82 VDD1.t4 B 0.094291f
C83 VDD1.t6 B 0.094291f
C84 VDD1.n1 B 0.768641f
C85 VDD1.t0 B 0.094291f
C86 VDD1.t7 B 0.094291f
C87 VDD1.n2 B 0.768641f
C88 VDD1.n3 B 2.39165f
C89 VDD1.t2 B 0.094291f
C90 VDD1.t3 B 0.094291f
C91 VDD1.n4 B 0.763331f
C92 VDD1.n5 B 2.11324f
C93 VTAIL.t9 B 0.088654f
C94 VTAIL.t11 B 0.088654f
C95 VTAIL.n0 B 0.658294f
C96 VTAIL.n1 B 0.354631f
C97 VTAIL.t10 B 0.839203f
C98 VTAIL.n2 B 0.446442f
C99 VTAIL.t6 B 0.839203f
C100 VTAIL.n3 B 0.446442f
C101 VTAIL.t7 B 0.088654f
C102 VTAIL.t4 B 0.088654f
C103 VTAIL.n4 B 0.658294f
C104 VTAIL.n5 B 0.487609f
C105 VTAIL.t1 B 0.839203f
C106 VTAIL.n6 B 1.17694f
C107 VTAIL.t8 B 0.839209f
C108 VTAIL.n7 B 1.17694f
C109 VTAIL.t15 B 0.088654f
C110 VTAIL.t12 B 0.088654f
C111 VTAIL.n8 B 0.658298f
C112 VTAIL.n9 B 0.487605f
C113 VTAIL.t13 B 0.839209f
C114 VTAIL.n10 B 0.446436f
C115 VTAIL.t0 B 0.839209f
C116 VTAIL.n11 B 0.446436f
C117 VTAIL.t2 B 0.088654f
C118 VTAIL.t3 B 0.088654f
C119 VTAIL.n12 B 0.658298f
C120 VTAIL.n13 B 0.487605f
C121 VTAIL.t5 B 0.839203f
C122 VTAIL.n14 B 1.17694f
C123 VTAIL.t14 B 0.839203f
C124 VTAIL.n15 B 1.17257f
C125 VP.n0 B 0.041631f
C126 VP.t0 B 0.70912f
C127 VP.n1 B 0.056028f
C128 VP.n2 B 0.031577f
C129 VP.t7 B 0.70912f
C130 VP.n3 B 0.046097f
C131 VP.n4 B 0.031577f
C132 VP.t1 B 0.70912f
C133 VP.n5 B 0.033119f
C134 VP.n6 B 0.041631f
C135 VP.t4 B 0.70912f
C136 VP.n7 B 0.056028f
C137 VP.n8 B 0.031577f
C138 VP.t5 B 0.70912f
C139 VP.n9 B 0.046097f
C140 VP.t2 B 0.846563f
C141 VP.n10 B 0.355054f
C142 VP.t6 B 0.70912f
C143 VP.n11 B 0.356287f
C144 VP.n12 B 0.047811f
C145 VP.n13 B 0.230482f
C146 VP.n14 B 0.031577f
C147 VP.n15 B 0.031577f
C148 VP.n16 B 0.046097f
C149 VP.n17 B 0.047811f
C150 VP.n18 B 0.283029f
C151 VP.n19 B 0.040837f
C152 VP.n20 B 0.031577f
C153 VP.n21 B 0.031577f
C154 VP.n22 B 0.031577f
C155 VP.n23 B 0.033119f
C156 VP.n24 B 0.05783f
C157 VP.n25 B 0.372029f
C158 VP.n26 B 1.30885f
C159 VP.n27 B 1.3361f
C160 VP.t3 B 0.70912f
C161 VP.n28 B 0.372029f
C162 VP.n29 B 0.05783f
C163 VP.n30 B 0.041631f
C164 VP.n31 B 0.031577f
C165 VP.n32 B 0.031577f
C166 VP.n33 B 0.056028f
C167 VP.n34 B 0.040837f
C168 VP.n35 B 0.283029f
C169 VP.n36 B 0.047811f
C170 VP.n37 B 0.031577f
C171 VP.n38 B 0.031577f
C172 VP.n39 B 0.031577f
C173 VP.n40 B 0.046097f
C174 VP.n41 B 0.047811f
C175 VP.n42 B 0.283029f
C176 VP.n43 B 0.040837f
C177 VP.n44 B 0.031577f
C178 VP.n45 B 0.031577f
C179 VP.n46 B 0.031577f
C180 VP.n47 B 0.033119f
C181 VP.n48 B 0.05783f
C182 VP.n49 B 0.372029f
C183 VP.n50 B 0.036212f
.ends

