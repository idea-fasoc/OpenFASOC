* NGSPICE file created from diff_pair_sample_0565.ext - technology: sky130A

.subckt diff_pair_sample_0565 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X1 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0 ps=0 w=5.47 l=1.8
X2 VDD2.t4 VN.t1 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X3 VTAIL.t3 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X4 VDD1.t8 VP.t1 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X5 VTAIL.t5 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X6 VDD1.t6 VP.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0.90255 ps=5.8 w=5.47 l=1.8
X7 VDD2.t1 VN.t2 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X8 VDD2.t6 VN.t3 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0.90255 ps=5.8 w=5.47 l=1.8
X9 VTAIL.t15 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X10 VTAIL.t8 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X11 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0 ps=0 w=5.47 l=1.8
X12 VDD1.t4 VP.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=2.1333 ps=11.72 w=5.47 l=1.8
X13 VDD2.t7 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=2.1333 ps=11.72 w=5.47 l=1.8
X14 VTAIL.t0 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X15 VDD2.t8 VN.t6 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0.90255 ps=5.8 w=5.47 l=1.8
X16 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0 ps=0 w=5.47 l=1.8
X17 VDD2.t9 VN.t7 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=2.1333 ps=11.72 w=5.47 l=1.8
X18 VDD1.t2 VP.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=2.1333 ps=11.72 w=5.47 l=1.8
X19 VDD1.t1 VP.t8 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0.90255 ps=5.8 w=5.47 l=1.8
X20 VDD1.t0 VP.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.1333 pd=11.72 as=0 ps=0 w=5.47 l=1.8
X22 VTAIL.t11 VN.t8 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
X23 VTAIL.t10 VN.t9 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=0.90255 pd=5.8 as=0.90255 ps=5.8 w=5.47 l=1.8
R0 VN.n31 VN.n30 185.279
R1 VN.n63 VN.n62 185.279
R2 VN.n61 VN.n32 161.3
R3 VN.n60 VN.n59 161.3
R4 VN.n58 VN.n33 161.3
R5 VN.n57 VN.n56 161.3
R6 VN.n55 VN.n34 161.3
R7 VN.n53 VN.n52 161.3
R8 VN.n51 VN.n35 161.3
R9 VN.n50 VN.n49 161.3
R10 VN.n48 VN.n36 161.3
R11 VN.n46 VN.n45 161.3
R12 VN.n44 VN.n37 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n41 VN.n38 161.3
R15 VN.n29 VN.n0 161.3
R16 VN.n28 VN.n27 161.3
R17 VN.n26 VN.n1 161.3
R18 VN.n25 VN.n24 161.3
R19 VN.n23 VN.n2 161.3
R20 VN.n21 VN.n20 161.3
R21 VN.n19 VN.n3 161.3
R22 VN.n18 VN.n17 161.3
R23 VN.n16 VN.n4 161.3
R24 VN.n14 VN.n13 161.3
R25 VN.n12 VN.n5 161.3
R26 VN.n11 VN.n10 161.3
R27 VN.n9 VN.n6 161.3
R28 VN.n7 VN.t6 105.445
R29 VN.n39 VN.t5 105.445
R30 VN.n8 VN.t0 73.2377
R31 VN.n15 VN.t1 73.2377
R32 VN.n22 VN.t4 73.2377
R33 VN.n30 VN.t7 73.2377
R34 VN.n40 VN.t8 73.2377
R35 VN.n47 VN.t2 73.2377
R36 VN.n54 VN.t9 73.2377
R37 VN.n62 VN.t3 73.2377
R38 VN.n10 VN.n5 56.5193
R39 VN.n17 VN.n3 56.5193
R40 VN.n42 VN.n37 56.5193
R41 VN.n49 VN.n35 56.5193
R42 VN.n8 VN.n7 51.0503
R43 VN.n40 VN.n39 51.0503
R44 VN.n24 VN.n1 45.8354
R45 VN.n56 VN.n33 45.8354
R46 VN VN.n63 44.0516
R47 VN.n28 VN.n1 35.1514
R48 VN.n60 VN.n33 35.1514
R49 VN.n10 VN.n9 24.4675
R50 VN.n14 VN.n5 24.4675
R51 VN.n17 VN.n16 24.4675
R52 VN.n21 VN.n3 24.4675
R53 VN.n24 VN.n23 24.4675
R54 VN.n29 VN.n28 24.4675
R55 VN.n42 VN.n41 24.4675
R56 VN.n49 VN.n48 24.4675
R57 VN.n46 VN.n37 24.4675
R58 VN.n56 VN.n55 24.4675
R59 VN.n53 VN.n35 24.4675
R60 VN.n61 VN.n60 24.4675
R61 VN.n9 VN.n8 18.5954
R62 VN.n22 VN.n21 18.5954
R63 VN.n41 VN.n40 18.5954
R64 VN.n54 VN.n53 18.5954
R65 VN.n39 VN.n38 12.5362
R66 VN.n7 VN.n6 12.5362
R67 VN.n15 VN.n14 12.234
R68 VN.n16 VN.n15 12.234
R69 VN.n48 VN.n47 12.234
R70 VN.n47 VN.n46 12.234
R71 VN.n23 VN.n22 5.87258
R72 VN.n55 VN.n54 5.87258
R73 VN.n30 VN.n29 0.48984
R74 VN.n62 VN.n61 0.48984
R75 VN.n63 VN.n32 0.189894
R76 VN.n59 VN.n32 0.189894
R77 VN.n59 VN.n58 0.189894
R78 VN.n58 VN.n57 0.189894
R79 VN.n57 VN.n34 0.189894
R80 VN.n52 VN.n34 0.189894
R81 VN.n52 VN.n51 0.189894
R82 VN.n51 VN.n50 0.189894
R83 VN.n50 VN.n36 0.189894
R84 VN.n45 VN.n36 0.189894
R85 VN.n45 VN.n44 0.189894
R86 VN.n44 VN.n43 0.189894
R87 VN.n43 VN.n38 0.189894
R88 VN.n11 VN.n6 0.189894
R89 VN.n12 VN.n11 0.189894
R90 VN.n13 VN.n12 0.189894
R91 VN.n13 VN.n4 0.189894
R92 VN.n18 VN.n4 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n20 VN.n19 0.189894
R95 VN.n20 VN.n2 0.189894
R96 VN.n25 VN.n2 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n27 VN.n26 0.189894
R99 VN.n27 VN.n0 0.189894
R100 VN.n31 VN.n0 0.189894
R101 VN VN.n31 0.0516364
R102 VDD2.n1 VDD2.t8 76.1066
R103 VDD2.n4 VDD2.t6 74.2713
R104 VDD2.n3 VDD2.n2 71.9733
R105 VDD2 VDD2.n7 71.9696
R106 VDD2.n6 VDD2.n5 70.6516
R107 VDD2.n1 VDD2.n0 70.6515
R108 VDD2.n4 VDD2.n3 37.1528
R109 VDD2.n7 VDD2.t2 3.62024
R110 VDD2.n7 VDD2.t7 3.62024
R111 VDD2.n5 VDD2.t5 3.62024
R112 VDD2.n5 VDD2.t1 3.62024
R113 VDD2.n2 VDD2.t3 3.62024
R114 VDD2.n2 VDD2.t9 3.62024
R115 VDD2.n0 VDD2.t0 3.62024
R116 VDD2.n0 VDD2.t4 3.62024
R117 VDD2.n6 VDD2.n4 1.83671
R118 VDD2 VDD2.n6 0.517741
R119 VDD2.n3 VDD2.n1 0.404206
R120 VTAIL.n11 VTAIL.t14 57.5926
R121 VTAIL.n16 VTAIL.t2 57.5916
R122 VTAIL.n17 VTAIL.t12 57.5916
R123 VTAIL.n2 VTAIL.t1 57.5916
R124 VTAIL.n15 VTAIL.n14 53.9728
R125 VTAIL.n13 VTAIL.n12 53.9728
R126 VTAIL.n10 VTAIL.n9 53.9728
R127 VTAIL.n8 VTAIL.n7 53.9728
R128 VTAIL.n19 VTAIL.n18 53.9727
R129 VTAIL.n1 VTAIL.n0 53.9727
R130 VTAIL.n4 VTAIL.n3 53.9727
R131 VTAIL.n6 VTAIL.n5 53.9727
R132 VTAIL.n8 VTAIL.n6 20.7548
R133 VTAIL.n17 VTAIL.n16 18.9186
R134 VTAIL.n18 VTAIL.t18 3.62024
R135 VTAIL.n18 VTAIL.t15 3.62024
R136 VTAIL.n0 VTAIL.t13 3.62024
R137 VTAIL.n0 VTAIL.t19 3.62024
R138 VTAIL.n3 VTAIL.t9 3.62024
R139 VTAIL.n3 VTAIL.t3 3.62024
R140 VTAIL.n5 VTAIL.t4 3.62024
R141 VTAIL.n5 VTAIL.t8 3.62024
R142 VTAIL.n14 VTAIL.t6 3.62024
R143 VTAIL.n14 VTAIL.t5 3.62024
R144 VTAIL.n12 VTAIL.t7 3.62024
R145 VTAIL.n12 VTAIL.t0 3.62024
R146 VTAIL.n9 VTAIL.t17 3.62024
R147 VTAIL.n9 VTAIL.t11 3.62024
R148 VTAIL.n7 VTAIL.t16 3.62024
R149 VTAIL.n7 VTAIL.t10 3.62024
R150 VTAIL.n10 VTAIL.n8 1.83671
R151 VTAIL.n11 VTAIL.n10 1.83671
R152 VTAIL.n15 VTAIL.n13 1.83671
R153 VTAIL.n16 VTAIL.n15 1.83671
R154 VTAIL.n6 VTAIL.n4 1.83671
R155 VTAIL.n4 VTAIL.n2 1.83671
R156 VTAIL.n19 VTAIL.n17 1.83671
R157 VTAIL VTAIL.n1 1.43584
R158 VTAIL.n13 VTAIL.n11 1.38843
R159 VTAIL.n2 VTAIL.n1 1.38843
R160 VTAIL VTAIL.n19 0.401362
R161 B.n646 B.n645 585
R162 B.n222 B.n111 585
R163 B.n221 B.n220 585
R164 B.n219 B.n218 585
R165 B.n217 B.n216 585
R166 B.n215 B.n214 585
R167 B.n213 B.n212 585
R168 B.n211 B.n210 585
R169 B.n209 B.n208 585
R170 B.n207 B.n206 585
R171 B.n205 B.n204 585
R172 B.n203 B.n202 585
R173 B.n201 B.n200 585
R174 B.n199 B.n198 585
R175 B.n197 B.n196 585
R176 B.n195 B.n194 585
R177 B.n193 B.n192 585
R178 B.n191 B.n190 585
R179 B.n189 B.n188 585
R180 B.n187 B.n186 585
R181 B.n185 B.n184 585
R182 B.n183 B.n182 585
R183 B.n181 B.n180 585
R184 B.n179 B.n178 585
R185 B.n177 B.n176 585
R186 B.n175 B.n174 585
R187 B.n173 B.n172 585
R188 B.n171 B.n170 585
R189 B.n169 B.n168 585
R190 B.n167 B.n166 585
R191 B.n165 B.n164 585
R192 B.n163 B.n162 585
R193 B.n161 B.n160 585
R194 B.n159 B.n158 585
R195 B.n157 B.n156 585
R196 B.n155 B.n154 585
R197 B.n153 B.n152 585
R198 B.n151 B.n150 585
R199 B.n149 B.n148 585
R200 B.n147 B.n146 585
R201 B.n145 B.n144 585
R202 B.n143 B.n142 585
R203 B.n141 B.n140 585
R204 B.n139 B.n138 585
R205 B.n137 B.n136 585
R206 B.n135 B.n134 585
R207 B.n133 B.n132 585
R208 B.n131 B.n130 585
R209 B.n129 B.n128 585
R210 B.n127 B.n126 585
R211 B.n125 B.n124 585
R212 B.n123 B.n122 585
R213 B.n121 B.n120 585
R214 B.n119 B.n118 585
R215 B.n644 B.n84 585
R216 B.n649 B.n84 585
R217 B.n643 B.n83 585
R218 B.n650 B.n83 585
R219 B.n642 B.n641 585
R220 B.n641 B.n79 585
R221 B.n640 B.n78 585
R222 B.n656 B.n78 585
R223 B.n639 B.n77 585
R224 B.n657 B.n77 585
R225 B.n638 B.n76 585
R226 B.n658 B.n76 585
R227 B.n637 B.n636 585
R228 B.n636 B.n75 585
R229 B.n635 B.n71 585
R230 B.n664 B.n71 585
R231 B.n634 B.n70 585
R232 B.n665 B.n70 585
R233 B.n633 B.n69 585
R234 B.n666 B.n69 585
R235 B.n632 B.n631 585
R236 B.n631 B.n65 585
R237 B.n630 B.n64 585
R238 B.n672 B.n64 585
R239 B.n629 B.n63 585
R240 B.n673 B.n63 585
R241 B.n628 B.n62 585
R242 B.n674 B.n62 585
R243 B.n627 B.n626 585
R244 B.n626 B.n58 585
R245 B.n625 B.n57 585
R246 B.n680 B.n57 585
R247 B.n624 B.n56 585
R248 B.n681 B.n56 585
R249 B.n623 B.n55 585
R250 B.n682 B.n55 585
R251 B.n622 B.n621 585
R252 B.n621 B.n51 585
R253 B.n620 B.n50 585
R254 B.n688 B.n50 585
R255 B.n619 B.n49 585
R256 B.n689 B.n49 585
R257 B.n618 B.n48 585
R258 B.n690 B.n48 585
R259 B.n617 B.n616 585
R260 B.n616 B.n44 585
R261 B.n615 B.n43 585
R262 B.n696 B.n43 585
R263 B.n614 B.n42 585
R264 B.n697 B.n42 585
R265 B.n613 B.n41 585
R266 B.n698 B.n41 585
R267 B.n612 B.n611 585
R268 B.n611 B.n37 585
R269 B.n610 B.n36 585
R270 B.n704 B.n36 585
R271 B.n609 B.n35 585
R272 B.n705 B.n35 585
R273 B.n608 B.n34 585
R274 B.n706 B.n34 585
R275 B.n607 B.n606 585
R276 B.n606 B.n30 585
R277 B.n605 B.n29 585
R278 B.n712 B.n29 585
R279 B.n604 B.n28 585
R280 B.n713 B.n28 585
R281 B.n603 B.n27 585
R282 B.n714 B.n27 585
R283 B.n602 B.n601 585
R284 B.n601 B.n26 585
R285 B.n600 B.n22 585
R286 B.n720 B.n22 585
R287 B.n599 B.n21 585
R288 B.n721 B.n21 585
R289 B.n598 B.n20 585
R290 B.n722 B.n20 585
R291 B.n597 B.n596 585
R292 B.n596 B.n16 585
R293 B.n595 B.n15 585
R294 B.n728 B.n15 585
R295 B.n594 B.n14 585
R296 B.n729 B.n14 585
R297 B.n593 B.n13 585
R298 B.n730 B.n13 585
R299 B.n592 B.n591 585
R300 B.n591 B.n12 585
R301 B.n590 B.n589 585
R302 B.n590 B.n8 585
R303 B.n588 B.n7 585
R304 B.n737 B.n7 585
R305 B.n587 B.n6 585
R306 B.n738 B.n6 585
R307 B.n586 B.n5 585
R308 B.n739 B.n5 585
R309 B.n585 B.n584 585
R310 B.n584 B.n4 585
R311 B.n583 B.n223 585
R312 B.n583 B.n582 585
R313 B.n573 B.n224 585
R314 B.n225 B.n224 585
R315 B.n575 B.n574 585
R316 B.n576 B.n575 585
R317 B.n572 B.n229 585
R318 B.n233 B.n229 585
R319 B.n571 B.n570 585
R320 B.n570 B.n569 585
R321 B.n231 B.n230 585
R322 B.n232 B.n231 585
R323 B.n562 B.n561 585
R324 B.n563 B.n562 585
R325 B.n560 B.n238 585
R326 B.n238 B.n237 585
R327 B.n559 B.n558 585
R328 B.n558 B.n557 585
R329 B.n240 B.n239 585
R330 B.n550 B.n240 585
R331 B.n549 B.n548 585
R332 B.n551 B.n549 585
R333 B.n547 B.n245 585
R334 B.n245 B.n244 585
R335 B.n546 B.n545 585
R336 B.n545 B.n544 585
R337 B.n247 B.n246 585
R338 B.n248 B.n247 585
R339 B.n537 B.n536 585
R340 B.n538 B.n537 585
R341 B.n535 B.n252 585
R342 B.n256 B.n252 585
R343 B.n534 B.n533 585
R344 B.n533 B.n532 585
R345 B.n254 B.n253 585
R346 B.n255 B.n254 585
R347 B.n525 B.n524 585
R348 B.n526 B.n525 585
R349 B.n523 B.n261 585
R350 B.n261 B.n260 585
R351 B.n522 B.n521 585
R352 B.n521 B.n520 585
R353 B.n263 B.n262 585
R354 B.n264 B.n263 585
R355 B.n513 B.n512 585
R356 B.n514 B.n513 585
R357 B.n511 B.n269 585
R358 B.n269 B.n268 585
R359 B.n510 B.n509 585
R360 B.n509 B.n508 585
R361 B.n271 B.n270 585
R362 B.n272 B.n271 585
R363 B.n501 B.n500 585
R364 B.n502 B.n501 585
R365 B.n499 B.n277 585
R366 B.n277 B.n276 585
R367 B.n498 B.n497 585
R368 B.n497 B.n496 585
R369 B.n279 B.n278 585
R370 B.n280 B.n279 585
R371 B.n489 B.n488 585
R372 B.n490 B.n489 585
R373 B.n487 B.n285 585
R374 B.n285 B.n284 585
R375 B.n486 B.n485 585
R376 B.n485 B.n484 585
R377 B.n287 B.n286 585
R378 B.n288 B.n287 585
R379 B.n477 B.n476 585
R380 B.n478 B.n477 585
R381 B.n475 B.n293 585
R382 B.n293 B.n292 585
R383 B.n474 B.n473 585
R384 B.n473 B.n472 585
R385 B.n295 B.n294 585
R386 B.n465 B.n295 585
R387 B.n464 B.n463 585
R388 B.n466 B.n464 585
R389 B.n462 B.n300 585
R390 B.n300 B.n299 585
R391 B.n461 B.n460 585
R392 B.n460 B.n459 585
R393 B.n302 B.n301 585
R394 B.n303 B.n302 585
R395 B.n452 B.n451 585
R396 B.n453 B.n452 585
R397 B.n450 B.n308 585
R398 B.n308 B.n307 585
R399 B.n445 B.n444 585
R400 B.n443 B.n337 585
R401 B.n442 B.n336 585
R402 B.n447 B.n336 585
R403 B.n441 B.n440 585
R404 B.n439 B.n438 585
R405 B.n437 B.n436 585
R406 B.n435 B.n434 585
R407 B.n433 B.n432 585
R408 B.n431 B.n430 585
R409 B.n429 B.n428 585
R410 B.n427 B.n426 585
R411 B.n425 B.n424 585
R412 B.n423 B.n422 585
R413 B.n421 B.n420 585
R414 B.n419 B.n418 585
R415 B.n417 B.n416 585
R416 B.n415 B.n414 585
R417 B.n413 B.n412 585
R418 B.n411 B.n410 585
R419 B.n409 B.n408 585
R420 B.n407 B.n406 585
R421 B.n405 B.n404 585
R422 B.n402 B.n401 585
R423 B.n400 B.n399 585
R424 B.n398 B.n397 585
R425 B.n396 B.n395 585
R426 B.n394 B.n393 585
R427 B.n392 B.n391 585
R428 B.n390 B.n389 585
R429 B.n388 B.n387 585
R430 B.n386 B.n385 585
R431 B.n384 B.n383 585
R432 B.n381 B.n380 585
R433 B.n379 B.n378 585
R434 B.n377 B.n376 585
R435 B.n375 B.n374 585
R436 B.n373 B.n372 585
R437 B.n371 B.n370 585
R438 B.n369 B.n368 585
R439 B.n367 B.n366 585
R440 B.n365 B.n364 585
R441 B.n363 B.n362 585
R442 B.n361 B.n360 585
R443 B.n359 B.n358 585
R444 B.n357 B.n356 585
R445 B.n355 B.n354 585
R446 B.n353 B.n352 585
R447 B.n351 B.n350 585
R448 B.n349 B.n348 585
R449 B.n347 B.n346 585
R450 B.n345 B.n344 585
R451 B.n343 B.n342 585
R452 B.n310 B.n309 585
R453 B.n449 B.n448 585
R454 B.n448 B.n447 585
R455 B.n306 B.n305 585
R456 B.n307 B.n306 585
R457 B.n455 B.n454 585
R458 B.n454 B.n453 585
R459 B.n456 B.n304 585
R460 B.n304 B.n303 585
R461 B.n458 B.n457 585
R462 B.n459 B.n458 585
R463 B.n298 B.n297 585
R464 B.n299 B.n298 585
R465 B.n468 B.n467 585
R466 B.n467 B.n466 585
R467 B.n469 B.n296 585
R468 B.n465 B.n296 585
R469 B.n471 B.n470 585
R470 B.n472 B.n471 585
R471 B.n291 B.n290 585
R472 B.n292 B.n291 585
R473 B.n480 B.n479 585
R474 B.n479 B.n478 585
R475 B.n481 B.n289 585
R476 B.n289 B.n288 585
R477 B.n483 B.n482 585
R478 B.n484 B.n483 585
R479 B.n283 B.n282 585
R480 B.n284 B.n283 585
R481 B.n492 B.n491 585
R482 B.n491 B.n490 585
R483 B.n493 B.n281 585
R484 B.n281 B.n280 585
R485 B.n495 B.n494 585
R486 B.n496 B.n495 585
R487 B.n275 B.n274 585
R488 B.n276 B.n275 585
R489 B.n504 B.n503 585
R490 B.n503 B.n502 585
R491 B.n505 B.n273 585
R492 B.n273 B.n272 585
R493 B.n507 B.n506 585
R494 B.n508 B.n507 585
R495 B.n267 B.n266 585
R496 B.n268 B.n267 585
R497 B.n516 B.n515 585
R498 B.n515 B.n514 585
R499 B.n517 B.n265 585
R500 B.n265 B.n264 585
R501 B.n519 B.n518 585
R502 B.n520 B.n519 585
R503 B.n259 B.n258 585
R504 B.n260 B.n259 585
R505 B.n528 B.n527 585
R506 B.n527 B.n526 585
R507 B.n529 B.n257 585
R508 B.n257 B.n255 585
R509 B.n531 B.n530 585
R510 B.n532 B.n531 585
R511 B.n251 B.n250 585
R512 B.n256 B.n251 585
R513 B.n540 B.n539 585
R514 B.n539 B.n538 585
R515 B.n541 B.n249 585
R516 B.n249 B.n248 585
R517 B.n543 B.n542 585
R518 B.n544 B.n543 585
R519 B.n243 B.n242 585
R520 B.n244 B.n243 585
R521 B.n553 B.n552 585
R522 B.n552 B.n551 585
R523 B.n554 B.n241 585
R524 B.n550 B.n241 585
R525 B.n556 B.n555 585
R526 B.n557 B.n556 585
R527 B.n236 B.n235 585
R528 B.n237 B.n236 585
R529 B.n565 B.n564 585
R530 B.n564 B.n563 585
R531 B.n566 B.n234 585
R532 B.n234 B.n232 585
R533 B.n568 B.n567 585
R534 B.n569 B.n568 585
R535 B.n228 B.n227 585
R536 B.n233 B.n228 585
R537 B.n578 B.n577 585
R538 B.n577 B.n576 585
R539 B.n579 B.n226 585
R540 B.n226 B.n225 585
R541 B.n581 B.n580 585
R542 B.n582 B.n581 585
R543 B.n3 B.n0 585
R544 B.n4 B.n3 585
R545 B.n736 B.n1 585
R546 B.n737 B.n736 585
R547 B.n735 B.n734 585
R548 B.n735 B.n8 585
R549 B.n733 B.n9 585
R550 B.n12 B.n9 585
R551 B.n732 B.n731 585
R552 B.n731 B.n730 585
R553 B.n11 B.n10 585
R554 B.n729 B.n11 585
R555 B.n727 B.n726 585
R556 B.n728 B.n727 585
R557 B.n725 B.n17 585
R558 B.n17 B.n16 585
R559 B.n724 B.n723 585
R560 B.n723 B.n722 585
R561 B.n19 B.n18 585
R562 B.n721 B.n19 585
R563 B.n719 B.n718 585
R564 B.n720 B.n719 585
R565 B.n717 B.n23 585
R566 B.n26 B.n23 585
R567 B.n716 B.n715 585
R568 B.n715 B.n714 585
R569 B.n25 B.n24 585
R570 B.n713 B.n25 585
R571 B.n711 B.n710 585
R572 B.n712 B.n711 585
R573 B.n709 B.n31 585
R574 B.n31 B.n30 585
R575 B.n708 B.n707 585
R576 B.n707 B.n706 585
R577 B.n33 B.n32 585
R578 B.n705 B.n33 585
R579 B.n703 B.n702 585
R580 B.n704 B.n703 585
R581 B.n701 B.n38 585
R582 B.n38 B.n37 585
R583 B.n700 B.n699 585
R584 B.n699 B.n698 585
R585 B.n40 B.n39 585
R586 B.n697 B.n40 585
R587 B.n695 B.n694 585
R588 B.n696 B.n695 585
R589 B.n693 B.n45 585
R590 B.n45 B.n44 585
R591 B.n692 B.n691 585
R592 B.n691 B.n690 585
R593 B.n47 B.n46 585
R594 B.n689 B.n47 585
R595 B.n687 B.n686 585
R596 B.n688 B.n687 585
R597 B.n685 B.n52 585
R598 B.n52 B.n51 585
R599 B.n684 B.n683 585
R600 B.n683 B.n682 585
R601 B.n54 B.n53 585
R602 B.n681 B.n54 585
R603 B.n679 B.n678 585
R604 B.n680 B.n679 585
R605 B.n677 B.n59 585
R606 B.n59 B.n58 585
R607 B.n676 B.n675 585
R608 B.n675 B.n674 585
R609 B.n61 B.n60 585
R610 B.n673 B.n61 585
R611 B.n671 B.n670 585
R612 B.n672 B.n671 585
R613 B.n669 B.n66 585
R614 B.n66 B.n65 585
R615 B.n668 B.n667 585
R616 B.n667 B.n666 585
R617 B.n68 B.n67 585
R618 B.n665 B.n68 585
R619 B.n663 B.n662 585
R620 B.n664 B.n663 585
R621 B.n661 B.n72 585
R622 B.n75 B.n72 585
R623 B.n660 B.n659 585
R624 B.n659 B.n658 585
R625 B.n74 B.n73 585
R626 B.n657 B.n74 585
R627 B.n655 B.n654 585
R628 B.n656 B.n655 585
R629 B.n653 B.n80 585
R630 B.n80 B.n79 585
R631 B.n652 B.n651 585
R632 B.n651 B.n650 585
R633 B.n82 B.n81 585
R634 B.n649 B.n82 585
R635 B.n740 B.n739 585
R636 B.n738 B.n2 585
R637 B.n118 B.n82 564.573
R638 B.n646 B.n84 564.573
R639 B.n448 B.n308 564.573
R640 B.n445 B.n306 564.573
R641 B.n115 B.t17 279.644
R642 B.n112 B.t21 279.644
R643 B.n340 B.t14 279.644
R644 B.n338 B.t10 279.644
R645 B.n648 B.n647 256.663
R646 B.n648 B.n110 256.663
R647 B.n648 B.n109 256.663
R648 B.n648 B.n108 256.663
R649 B.n648 B.n107 256.663
R650 B.n648 B.n106 256.663
R651 B.n648 B.n105 256.663
R652 B.n648 B.n104 256.663
R653 B.n648 B.n103 256.663
R654 B.n648 B.n102 256.663
R655 B.n648 B.n101 256.663
R656 B.n648 B.n100 256.663
R657 B.n648 B.n99 256.663
R658 B.n648 B.n98 256.663
R659 B.n648 B.n97 256.663
R660 B.n648 B.n96 256.663
R661 B.n648 B.n95 256.663
R662 B.n648 B.n94 256.663
R663 B.n648 B.n93 256.663
R664 B.n648 B.n92 256.663
R665 B.n648 B.n91 256.663
R666 B.n648 B.n90 256.663
R667 B.n648 B.n89 256.663
R668 B.n648 B.n88 256.663
R669 B.n648 B.n87 256.663
R670 B.n648 B.n86 256.663
R671 B.n648 B.n85 256.663
R672 B.n447 B.n446 256.663
R673 B.n447 B.n311 256.663
R674 B.n447 B.n312 256.663
R675 B.n447 B.n313 256.663
R676 B.n447 B.n314 256.663
R677 B.n447 B.n315 256.663
R678 B.n447 B.n316 256.663
R679 B.n447 B.n317 256.663
R680 B.n447 B.n318 256.663
R681 B.n447 B.n319 256.663
R682 B.n447 B.n320 256.663
R683 B.n447 B.n321 256.663
R684 B.n447 B.n322 256.663
R685 B.n447 B.n323 256.663
R686 B.n447 B.n324 256.663
R687 B.n447 B.n325 256.663
R688 B.n447 B.n326 256.663
R689 B.n447 B.n327 256.663
R690 B.n447 B.n328 256.663
R691 B.n447 B.n329 256.663
R692 B.n447 B.n330 256.663
R693 B.n447 B.n331 256.663
R694 B.n447 B.n332 256.663
R695 B.n447 B.n333 256.663
R696 B.n447 B.n334 256.663
R697 B.n447 B.n335 256.663
R698 B.n742 B.n741 256.663
R699 B.n122 B.n121 163.367
R700 B.n126 B.n125 163.367
R701 B.n130 B.n129 163.367
R702 B.n134 B.n133 163.367
R703 B.n138 B.n137 163.367
R704 B.n142 B.n141 163.367
R705 B.n146 B.n145 163.367
R706 B.n150 B.n149 163.367
R707 B.n154 B.n153 163.367
R708 B.n158 B.n157 163.367
R709 B.n162 B.n161 163.367
R710 B.n166 B.n165 163.367
R711 B.n170 B.n169 163.367
R712 B.n174 B.n173 163.367
R713 B.n178 B.n177 163.367
R714 B.n182 B.n181 163.367
R715 B.n186 B.n185 163.367
R716 B.n190 B.n189 163.367
R717 B.n194 B.n193 163.367
R718 B.n198 B.n197 163.367
R719 B.n202 B.n201 163.367
R720 B.n206 B.n205 163.367
R721 B.n210 B.n209 163.367
R722 B.n214 B.n213 163.367
R723 B.n218 B.n217 163.367
R724 B.n220 B.n111 163.367
R725 B.n452 B.n308 163.367
R726 B.n452 B.n302 163.367
R727 B.n460 B.n302 163.367
R728 B.n460 B.n300 163.367
R729 B.n464 B.n300 163.367
R730 B.n464 B.n295 163.367
R731 B.n473 B.n295 163.367
R732 B.n473 B.n293 163.367
R733 B.n477 B.n293 163.367
R734 B.n477 B.n287 163.367
R735 B.n485 B.n287 163.367
R736 B.n485 B.n285 163.367
R737 B.n489 B.n285 163.367
R738 B.n489 B.n279 163.367
R739 B.n497 B.n279 163.367
R740 B.n497 B.n277 163.367
R741 B.n501 B.n277 163.367
R742 B.n501 B.n271 163.367
R743 B.n509 B.n271 163.367
R744 B.n509 B.n269 163.367
R745 B.n513 B.n269 163.367
R746 B.n513 B.n263 163.367
R747 B.n521 B.n263 163.367
R748 B.n521 B.n261 163.367
R749 B.n525 B.n261 163.367
R750 B.n525 B.n254 163.367
R751 B.n533 B.n254 163.367
R752 B.n533 B.n252 163.367
R753 B.n537 B.n252 163.367
R754 B.n537 B.n247 163.367
R755 B.n545 B.n247 163.367
R756 B.n545 B.n245 163.367
R757 B.n549 B.n245 163.367
R758 B.n549 B.n240 163.367
R759 B.n558 B.n240 163.367
R760 B.n558 B.n238 163.367
R761 B.n562 B.n238 163.367
R762 B.n562 B.n231 163.367
R763 B.n570 B.n231 163.367
R764 B.n570 B.n229 163.367
R765 B.n575 B.n229 163.367
R766 B.n575 B.n224 163.367
R767 B.n583 B.n224 163.367
R768 B.n584 B.n583 163.367
R769 B.n584 B.n5 163.367
R770 B.n6 B.n5 163.367
R771 B.n7 B.n6 163.367
R772 B.n590 B.n7 163.367
R773 B.n591 B.n590 163.367
R774 B.n591 B.n13 163.367
R775 B.n14 B.n13 163.367
R776 B.n15 B.n14 163.367
R777 B.n596 B.n15 163.367
R778 B.n596 B.n20 163.367
R779 B.n21 B.n20 163.367
R780 B.n22 B.n21 163.367
R781 B.n601 B.n22 163.367
R782 B.n601 B.n27 163.367
R783 B.n28 B.n27 163.367
R784 B.n29 B.n28 163.367
R785 B.n606 B.n29 163.367
R786 B.n606 B.n34 163.367
R787 B.n35 B.n34 163.367
R788 B.n36 B.n35 163.367
R789 B.n611 B.n36 163.367
R790 B.n611 B.n41 163.367
R791 B.n42 B.n41 163.367
R792 B.n43 B.n42 163.367
R793 B.n616 B.n43 163.367
R794 B.n616 B.n48 163.367
R795 B.n49 B.n48 163.367
R796 B.n50 B.n49 163.367
R797 B.n621 B.n50 163.367
R798 B.n621 B.n55 163.367
R799 B.n56 B.n55 163.367
R800 B.n57 B.n56 163.367
R801 B.n626 B.n57 163.367
R802 B.n626 B.n62 163.367
R803 B.n63 B.n62 163.367
R804 B.n64 B.n63 163.367
R805 B.n631 B.n64 163.367
R806 B.n631 B.n69 163.367
R807 B.n70 B.n69 163.367
R808 B.n71 B.n70 163.367
R809 B.n636 B.n71 163.367
R810 B.n636 B.n76 163.367
R811 B.n77 B.n76 163.367
R812 B.n78 B.n77 163.367
R813 B.n641 B.n78 163.367
R814 B.n641 B.n83 163.367
R815 B.n84 B.n83 163.367
R816 B.n337 B.n336 163.367
R817 B.n440 B.n336 163.367
R818 B.n438 B.n437 163.367
R819 B.n434 B.n433 163.367
R820 B.n430 B.n429 163.367
R821 B.n426 B.n425 163.367
R822 B.n422 B.n421 163.367
R823 B.n418 B.n417 163.367
R824 B.n414 B.n413 163.367
R825 B.n410 B.n409 163.367
R826 B.n406 B.n405 163.367
R827 B.n401 B.n400 163.367
R828 B.n397 B.n396 163.367
R829 B.n393 B.n392 163.367
R830 B.n389 B.n388 163.367
R831 B.n385 B.n384 163.367
R832 B.n380 B.n379 163.367
R833 B.n376 B.n375 163.367
R834 B.n372 B.n371 163.367
R835 B.n368 B.n367 163.367
R836 B.n364 B.n363 163.367
R837 B.n360 B.n359 163.367
R838 B.n356 B.n355 163.367
R839 B.n352 B.n351 163.367
R840 B.n348 B.n347 163.367
R841 B.n344 B.n343 163.367
R842 B.n448 B.n310 163.367
R843 B.n454 B.n306 163.367
R844 B.n454 B.n304 163.367
R845 B.n458 B.n304 163.367
R846 B.n458 B.n298 163.367
R847 B.n467 B.n298 163.367
R848 B.n467 B.n296 163.367
R849 B.n471 B.n296 163.367
R850 B.n471 B.n291 163.367
R851 B.n479 B.n291 163.367
R852 B.n479 B.n289 163.367
R853 B.n483 B.n289 163.367
R854 B.n483 B.n283 163.367
R855 B.n491 B.n283 163.367
R856 B.n491 B.n281 163.367
R857 B.n495 B.n281 163.367
R858 B.n495 B.n275 163.367
R859 B.n503 B.n275 163.367
R860 B.n503 B.n273 163.367
R861 B.n507 B.n273 163.367
R862 B.n507 B.n267 163.367
R863 B.n515 B.n267 163.367
R864 B.n515 B.n265 163.367
R865 B.n519 B.n265 163.367
R866 B.n519 B.n259 163.367
R867 B.n527 B.n259 163.367
R868 B.n527 B.n257 163.367
R869 B.n531 B.n257 163.367
R870 B.n531 B.n251 163.367
R871 B.n539 B.n251 163.367
R872 B.n539 B.n249 163.367
R873 B.n543 B.n249 163.367
R874 B.n543 B.n243 163.367
R875 B.n552 B.n243 163.367
R876 B.n552 B.n241 163.367
R877 B.n556 B.n241 163.367
R878 B.n556 B.n236 163.367
R879 B.n564 B.n236 163.367
R880 B.n564 B.n234 163.367
R881 B.n568 B.n234 163.367
R882 B.n568 B.n228 163.367
R883 B.n577 B.n228 163.367
R884 B.n577 B.n226 163.367
R885 B.n581 B.n226 163.367
R886 B.n581 B.n3 163.367
R887 B.n740 B.n3 163.367
R888 B.n736 B.n2 163.367
R889 B.n736 B.n735 163.367
R890 B.n735 B.n9 163.367
R891 B.n731 B.n9 163.367
R892 B.n731 B.n11 163.367
R893 B.n727 B.n11 163.367
R894 B.n727 B.n17 163.367
R895 B.n723 B.n17 163.367
R896 B.n723 B.n19 163.367
R897 B.n719 B.n19 163.367
R898 B.n719 B.n23 163.367
R899 B.n715 B.n23 163.367
R900 B.n715 B.n25 163.367
R901 B.n711 B.n25 163.367
R902 B.n711 B.n31 163.367
R903 B.n707 B.n31 163.367
R904 B.n707 B.n33 163.367
R905 B.n703 B.n33 163.367
R906 B.n703 B.n38 163.367
R907 B.n699 B.n38 163.367
R908 B.n699 B.n40 163.367
R909 B.n695 B.n40 163.367
R910 B.n695 B.n45 163.367
R911 B.n691 B.n45 163.367
R912 B.n691 B.n47 163.367
R913 B.n687 B.n47 163.367
R914 B.n687 B.n52 163.367
R915 B.n683 B.n52 163.367
R916 B.n683 B.n54 163.367
R917 B.n679 B.n54 163.367
R918 B.n679 B.n59 163.367
R919 B.n675 B.n59 163.367
R920 B.n675 B.n61 163.367
R921 B.n671 B.n61 163.367
R922 B.n671 B.n66 163.367
R923 B.n667 B.n66 163.367
R924 B.n667 B.n68 163.367
R925 B.n663 B.n68 163.367
R926 B.n663 B.n72 163.367
R927 B.n659 B.n72 163.367
R928 B.n659 B.n74 163.367
R929 B.n655 B.n74 163.367
R930 B.n655 B.n80 163.367
R931 B.n651 B.n80 163.367
R932 B.n651 B.n82 163.367
R933 B.n447 B.n307 140.251
R934 B.n649 B.n648 140.251
R935 B.n112 B.t22 111.675
R936 B.n340 B.t16 111.675
R937 B.n115 B.t19 111.669
R938 B.n338 B.t13 111.669
R939 B.n118 B.n85 71.676
R940 B.n122 B.n86 71.676
R941 B.n126 B.n87 71.676
R942 B.n130 B.n88 71.676
R943 B.n134 B.n89 71.676
R944 B.n138 B.n90 71.676
R945 B.n142 B.n91 71.676
R946 B.n146 B.n92 71.676
R947 B.n150 B.n93 71.676
R948 B.n154 B.n94 71.676
R949 B.n158 B.n95 71.676
R950 B.n162 B.n96 71.676
R951 B.n166 B.n97 71.676
R952 B.n170 B.n98 71.676
R953 B.n174 B.n99 71.676
R954 B.n178 B.n100 71.676
R955 B.n182 B.n101 71.676
R956 B.n186 B.n102 71.676
R957 B.n190 B.n103 71.676
R958 B.n194 B.n104 71.676
R959 B.n198 B.n105 71.676
R960 B.n202 B.n106 71.676
R961 B.n206 B.n107 71.676
R962 B.n210 B.n108 71.676
R963 B.n214 B.n109 71.676
R964 B.n218 B.n110 71.676
R965 B.n647 B.n111 71.676
R966 B.n647 B.n646 71.676
R967 B.n220 B.n110 71.676
R968 B.n217 B.n109 71.676
R969 B.n213 B.n108 71.676
R970 B.n209 B.n107 71.676
R971 B.n205 B.n106 71.676
R972 B.n201 B.n105 71.676
R973 B.n197 B.n104 71.676
R974 B.n193 B.n103 71.676
R975 B.n189 B.n102 71.676
R976 B.n185 B.n101 71.676
R977 B.n181 B.n100 71.676
R978 B.n177 B.n99 71.676
R979 B.n173 B.n98 71.676
R980 B.n169 B.n97 71.676
R981 B.n165 B.n96 71.676
R982 B.n161 B.n95 71.676
R983 B.n157 B.n94 71.676
R984 B.n153 B.n93 71.676
R985 B.n149 B.n92 71.676
R986 B.n145 B.n91 71.676
R987 B.n141 B.n90 71.676
R988 B.n137 B.n89 71.676
R989 B.n133 B.n88 71.676
R990 B.n129 B.n87 71.676
R991 B.n125 B.n86 71.676
R992 B.n121 B.n85 71.676
R993 B.n446 B.n445 71.676
R994 B.n440 B.n311 71.676
R995 B.n437 B.n312 71.676
R996 B.n433 B.n313 71.676
R997 B.n429 B.n314 71.676
R998 B.n425 B.n315 71.676
R999 B.n421 B.n316 71.676
R1000 B.n417 B.n317 71.676
R1001 B.n413 B.n318 71.676
R1002 B.n409 B.n319 71.676
R1003 B.n405 B.n320 71.676
R1004 B.n400 B.n321 71.676
R1005 B.n396 B.n322 71.676
R1006 B.n392 B.n323 71.676
R1007 B.n388 B.n324 71.676
R1008 B.n384 B.n325 71.676
R1009 B.n379 B.n326 71.676
R1010 B.n375 B.n327 71.676
R1011 B.n371 B.n328 71.676
R1012 B.n367 B.n329 71.676
R1013 B.n363 B.n330 71.676
R1014 B.n359 B.n331 71.676
R1015 B.n355 B.n332 71.676
R1016 B.n351 B.n333 71.676
R1017 B.n347 B.n334 71.676
R1018 B.n343 B.n335 71.676
R1019 B.n446 B.n337 71.676
R1020 B.n438 B.n311 71.676
R1021 B.n434 B.n312 71.676
R1022 B.n430 B.n313 71.676
R1023 B.n426 B.n314 71.676
R1024 B.n422 B.n315 71.676
R1025 B.n418 B.n316 71.676
R1026 B.n414 B.n317 71.676
R1027 B.n410 B.n318 71.676
R1028 B.n406 B.n319 71.676
R1029 B.n401 B.n320 71.676
R1030 B.n397 B.n321 71.676
R1031 B.n393 B.n322 71.676
R1032 B.n389 B.n323 71.676
R1033 B.n385 B.n324 71.676
R1034 B.n380 B.n325 71.676
R1035 B.n376 B.n326 71.676
R1036 B.n372 B.n327 71.676
R1037 B.n368 B.n328 71.676
R1038 B.n364 B.n329 71.676
R1039 B.n360 B.n330 71.676
R1040 B.n356 B.n331 71.676
R1041 B.n352 B.n332 71.676
R1042 B.n348 B.n333 71.676
R1043 B.n344 B.n334 71.676
R1044 B.n335 B.n310 71.676
R1045 B.n741 B.n740 71.676
R1046 B.n741 B.n2 71.676
R1047 B.n113 B.t23 70.3659
R1048 B.n341 B.t15 70.3659
R1049 B.n116 B.t20 70.3601
R1050 B.n339 B.t12 70.3601
R1051 B.n453 B.n307 69.6143
R1052 B.n453 B.n303 69.6143
R1053 B.n459 B.n303 69.6143
R1054 B.n459 B.n299 69.6143
R1055 B.n466 B.n299 69.6143
R1056 B.n466 B.n465 69.6143
R1057 B.n472 B.n292 69.6143
R1058 B.n478 B.n292 69.6143
R1059 B.n478 B.n288 69.6143
R1060 B.n484 B.n288 69.6143
R1061 B.n484 B.n284 69.6143
R1062 B.n490 B.n284 69.6143
R1063 B.n490 B.n280 69.6143
R1064 B.n496 B.n280 69.6143
R1065 B.n502 B.n276 69.6143
R1066 B.n502 B.n272 69.6143
R1067 B.n508 B.n272 69.6143
R1068 B.n508 B.n268 69.6143
R1069 B.n514 B.n268 69.6143
R1070 B.n520 B.n264 69.6143
R1071 B.n520 B.n260 69.6143
R1072 B.n526 B.n260 69.6143
R1073 B.n526 B.n255 69.6143
R1074 B.n532 B.n255 69.6143
R1075 B.n532 B.n256 69.6143
R1076 B.n538 B.n248 69.6143
R1077 B.n544 B.n248 69.6143
R1078 B.n544 B.n244 69.6143
R1079 B.n551 B.n244 69.6143
R1080 B.n551 B.n550 69.6143
R1081 B.n557 B.n237 69.6143
R1082 B.n563 B.n237 69.6143
R1083 B.n563 B.n232 69.6143
R1084 B.n569 B.n232 69.6143
R1085 B.n569 B.n233 69.6143
R1086 B.n576 B.n225 69.6143
R1087 B.n582 B.n225 69.6143
R1088 B.n582 B.n4 69.6143
R1089 B.n739 B.n4 69.6143
R1090 B.n739 B.n738 69.6143
R1091 B.n738 B.n737 69.6143
R1092 B.n737 B.n8 69.6143
R1093 B.n12 B.n8 69.6143
R1094 B.n730 B.n12 69.6143
R1095 B.n729 B.n728 69.6143
R1096 B.n728 B.n16 69.6143
R1097 B.n722 B.n16 69.6143
R1098 B.n722 B.n721 69.6143
R1099 B.n721 B.n720 69.6143
R1100 B.n714 B.n26 69.6143
R1101 B.n714 B.n713 69.6143
R1102 B.n713 B.n712 69.6143
R1103 B.n712 B.n30 69.6143
R1104 B.n706 B.n30 69.6143
R1105 B.n705 B.n704 69.6143
R1106 B.n704 B.n37 69.6143
R1107 B.n698 B.n37 69.6143
R1108 B.n698 B.n697 69.6143
R1109 B.n697 B.n696 69.6143
R1110 B.n696 B.n44 69.6143
R1111 B.n690 B.n689 69.6143
R1112 B.n689 B.n688 69.6143
R1113 B.n688 B.n51 69.6143
R1114 B.n682 B.n51 69.6143
R1115 B.n682 B.n681 69.6143
R1116 B.n680 B.n58 69.6143
R1117 B.n674 B.n58 69.6143
R1118 B.n674 B.n673 69.6143
R1119 B.n673 B.n672 69.6143
R1120 B.n672 B.n65 69.6143
R1121 B.n666 B.n65 69.6143
R1122 B.n666 B.n665 69.6143
R1123 B.n665 B.n664 69.6143
R1124 B.n658 B.n75 69.6143
R1125 B.n658 B.n657 69.6143
R1126 B.n657 B.n656 69.6143
R1127 B.n656 B.n79 69.6143
R1128 B.n650 B.n79 69.6143
R1129 B.n650 B.n649 69.6143
R1130 B.n514 B.t8 67.5668
R1131 B.n690 B.t5 67.5668
R1132 B.n117 B.n116 59.5399
R1133 B.n114 B.n113 59.5399
R1134 B.n382 B.n341 59.5399
R1135 B.n403 B.n339 59.5399
R1136 B.n472 B.t11 53.2346
R1137 B.n538 B.t9 53.2346
R1138 B.n233 B.t1 53.2346
R1139 B.t7 B.n729 53.2346
R1140 B.n706 B.t6 53.2346
R1141 B.n664 B.t18 53.2346
R1142 B.n496 B.t4 49.1396
R1143 B.t2 B.n680 49.1396
R1144 B.n116 B.n115 41.3096
R1145 B.n113 B.n112 41.3096
R1146 B.n341 B.n340 41.3096
R1147 B.n339 B.n338 41.3096
R1148 B.n444 B.n305 36.6834
R1149 B.n450 B.n449 36.6834
R1150 B.n645 B.n644 36.6834
R1151 B.n119 B.n81 36.6834
R1152 B.n550 B.t3 34.8074
R1153 B.n557 B.t3 34.8074
R1154 B.n720 B.t0 34.8074
R1155 B.n26 B.t0 34.8074
R1156 B.t4 B.n276 20.4751
R1157 B.n681 B.t2 20.4751
R1158 B B.n742 18.0485
R1159 B.n465 B.t11 16.3802
R1160 B.n256 B.t9 16.3802
R1161 B.n576 B.t1 16.3802
R1162 B.n730 B.t7 16.3802
R1163 B.t6 B.n705 16.3802
R1164 B.n75 B.t18 16.3802
R1165 B.n455 B.n305 10.6151
R1166 B.n456 B.n455 10.6151
R1167 B.n457 B.n456 10.6151
R1168 B.n457 B.n297 10.6151
R1169 B.n468 B.n297 10.6151
R1170 B.n469 B.n468 10.6151
R1171 B.n470 B.n469 10.6151
R1172 B.n470 B.n290 10.6151
R1173 B.n480 B.n290 10.6151
R1174 B.n481 B.n480 10.6151
R1175 B.n482 B.n481 10.6151
R1176 B.n482 B.n282 10.6151
R1177 B.n492 B.n282 10.6151
R1178 B.n493 B.n492 10.6151
R1179 B.n494 B.n493 10.6151
R1180 B.n494 B.n274 10.6151
R1181 B.n504 B.n274 10.6151
R1182 B.n505 B.n504 10.6151
R1183 B.n506 B.n505 10.6151
R1184 B.n506 B.n266 10.6151
R1185 B.n516 B.n266 10.6151
R1186 B.n517 B.n516 10.6151
R1187 B.n518 B.n517 10.6151
R1188 B.n518 B.n258 10.6151
R1189 B.n528 B.n258 10.6151
R1190 B.n529 B.n528 10.6151
R1191 B.n530 B.n529 10.6151
R1192 B.n530 B.n250 10.6151
R1193 B.n540 B.n250 10.6151
R1194 B.n541 B.n540 10.6151
R1195 B.n542 B.n541 10.6151
R1196 B.n542 B.n242 10.6151
R1197 B.n553 B.n242 10.6151
R1198 B.n554 B.n553 10.6151
R1199 B.n555 B.n554 10.6151
R1200 B.n555 B.n235 10.6151
R1201 B.n565 B.n235 10.6151
R1202 B.n566 B.n565 10.6151
R1203 B.n567 B.n566 10.6151
R1204 B.n567 B.n227 10.6151
R1205 B.n578 B.n227 10.6151
R1206 B.n579 B.n578 10.6151
R1207 B.n580 B.n579 10.6151
R1208 B.n580 B.n0 10.6151
R1209 B.n444 B.n443 10.6151
R1210 B.n443 B.n442 10.6151
R1211 B.n442 B.n441 10.6151
R1212 B.n441 B.n439 10.6151
R1213 B.n439 B.n436 10.6151
R1214 B.n436 B.n435 10.6151
R1215 B.n435 B.n432 10.6151
R1216 B.n432 B.n431 10.6151
R1217 B.n431 B.n428 10.6151
R1218 B.n428 B.n427 10.6151
R1219 B.n427 B.n424 10.6151
R1220 B.n424 B.n423 10.6151
R1221 B.n423 B.n420 10.6151
R1222 B.n420 B.n419 10.6151
R1223 B.n419 B.n416 10.6151
R1224 B.n416 B.n415 10.6151
R1225 B.n415 B.n412 10.6151
R1226 B.n412 B.n411 10.6151
R1227 B.n411 B.n408 10.6151
R1228 B.n408 B.n407 10.6151
R1229 B.n407 B.n404 10.6151
R1230 B.n402 B.n399 10.6151
R1231 B.n399 B.n398 10.6151
R1232 B.n398 B.n395 10.6151
R1233 B.n395 B.n394 10.6151
R1234 B.n394 B.n391 10.6151
R1235 B.n391 B.n390 10.6151
R1236 B.n390 B.n387 10.6151
R1237 B.n387 B.n386 10.6151
R1238 B.n386 B.n383 10.6151
R1239 B.n381 B.n378 10.6151
R1240 B.n378 B.n377 10.6151
R1241 B.n377 B.n374 10.6151
R1242 B.n374 B.n373 10.6151
R1243 B.n373 B.n370 10.6151
R1244 B.n370 B.n369 10.6151
R1245 B.n369 B.n366 10.6151
R1246 B.n366 B.n365 10.6151
R1247 B.n365 B.n362 10.6151
R1248 B.n362 B.n361 10.6151
R1249 B.n361 B.n358 10.6151
R1250 B.n358 B.n357 10.6151
R1251 B.n357 B.n354 10.6151
R1252 B.n354 B.n353 10.6151
R1253 B.n353 B.n350 10.6151
R1254 B.n350 B.n349 10.6151
R1255 B.n349 B.n346 10.6151
R1256 B.n346 B.n345 10.6151
R1257 B.n345 B.n342 10.6151
R1258 B.n342 B.n309 10.6151
R1259 B.n449 B.n309 10.6151
R1260 B.n451 B.n450 10.6151
R1261 B.n451 B.n301 10.6151
R1262 B.n461 B.n301 10.6151
R1263 B.n462 B.n461 10.6151
R1264 B.n463 B.n462 10.6151
R1265 B.n463 B.n294 10.6151
R1266 B.n474 B.n294 10.6151
R1267 B.n475 B.n474 10.6151
R1268 B.n476 B.n475 10.6151
R1269 B.n476 B.n286 10.6151
R1270 B.n486 B.n286 10.6151
R1271 B.n487 B.n486 10.6151
R1272 B.n488 B.n487 10.6151
R1273 B.n488 B.n278 10.6151
R1274 B.n498 B.n278 10.6151
R1275 B.n499 B.n498 10.6151
R1276 B.n500 B.n499 10.6151
R1277 B.n500 B.n270 10.6151
R1278 B.n510 B.n270 10.6151
R1279 B.n511 B.n510 10.6151
R1280 B.n512 B.n511 10.6151
R1281 B.n512 B.n262 10.6151
R1282 B.n522 B.n262 10.6151
R1283 B.n523 B.n522 10.6151
R1284 B.n524 B.n523 10.6151
R1285 B.n524 B.n253 10.6151
R1286 B.n534 B.n253 10.6151
R1287 B.n535 B.n534 10.6151
R1288 B.n536 B.n535 10.6151
R1289 B.n536 B.n246 10.6151
R1290 B.n546 B.n246 10.6151
R1291 B.n547 B.n546 10.6151
R1292 B.n548 B.n547 10.6151
R1293 B.n548 B.n239 10.6151
R1294 B.n559 B.n239 10.6151
R1295 B.n560 B.n559 10.6151
R1296 B.n561 B.n560 10.6151
R1297 B.n561 B.n230 10.6151
R1298 B.n571 B.n230 10.6151
R1299 B.n572 B.n571 10.6151
R1300 B.n574 B.n572 10.6151
R1301 B.n574 B.n573 10.6151
R1302 B.n573 B.n223 10.6151
R1303 B.n585 B.n223 10.6151
R1304 B.n586 B.n585 10.6151
R1305 B.n587 B.n586 10.6151
R1306 B.n588 B.n587 10.6151
R1307 B.n589 B.n588 10.6151
R1308 B.n592 B.n589 10.6151
R1309 B.n593 B.n592 10.6151
R1310 B.n594 B.n593 10.6151
R1311 B.n595 B.n594 10.6151
R1312 B.n597 B.n595 10.6151
R1313 B.n598 B.n597 10.6151
R1314 B.n599 B.n598 10.6151
R1315 B.n600 B.n599 10.6151
R1316 B.n602 B.n600 10.6151
R1317 B.n603 B.n602 10.6151
R1318 B.n604 B.n603 10.6151
R1319 B.n605 B.n604 10.6151
R1320 B.n607 B.n605 10.6151
R1321 B.n608 B.n607 10.6151
R1322 B.n609 B.n608 10.6151
R1323 B.n610 B.n609 10.6151
R1324 B.n612 B.n610 10.6151
R1325 B.n613 B.n612 10.6151
R1326 B.n614 B.n613 10.6151
R1327 B.n615 B.n614 10.6151
R1328 B.n617 B.n615 10.6151
R1329 B.n618 B.n617 10.6151
R1330 B.n619 B.n618 10.6151
R1331 B.n620 B.n619 10.6151
R1332 B.n622 B.n620 10.6151
R1333 B.n623 B.n622 10.6151
R1334 B.n624 B.n623 10.6151
R1335 B.n625 B.n624 10.6151
R1336 B.n627 B.n625 10.6151
R1337 B.n628 B.n627 10.6151
R1338 B.n629 B.n628 10.6151
R1339 B.n630 B.n629 10.6151
R1340 B.n632 B.n630 10.6151
R1341 B.n633 B.n632 10.6151
R1342 B.n634 B.n633 10.6151
R1343 B.n635 B.n634 10.6151
R1344 B.n637 B.n635 10.6151
R1345 B.n638 B.n637 10.6151
R1346 B.n639 B.n638 10.6151
R1347 B.n640 B.n639 10.6151
R1348 B.n642 B.n640 10.6151
R1349 B.n643 B.n642 10.6151
R1350 B.n644 B.n643 10.6151
R1351 B.n734 B.n1 10.6151
R1352 B.n734 B.n733 10.6151
R1353 B.n733 B.n732 10.6151
R1354 B.n732 B.n10 10.6151
R1355 B.n726 B.n10 10.6151
R1356 B.n726 B.n725 10.6151
R1357 B.n725 B.n724 10.6151
R1358 B.n724 B.n18 10.6151
R1359 B.n718 B.n18 10.6151
R1360 B.n718 B.n717 10.6151
R1361 B.n717 B.n716 10.6151
R1362 B.n716 B.n24 10.6151
R1363 B.n710 B.n24 10.6151
R1364 B.n710 B.n709 10.6151
R1365 B.n709 B.n708 10.6151
R1366 B.n708 B.n32 10.6151
R1367 B.n702 B.n32 10.6151
R1368 B.n702 B.n701 10.6151
R1369 B.n701 B.n700 10.6151
R1370 B.n700 B.n39 10.6151
R1371 B.n694 B.n39 10.6151
R1372 B.n694 B.n693 10.6151
R1373 B.n693 B.n692 10.6151
R1374 B.n692 B.n46 10.6151
R1375 B.n686 B.n46 10.6151
R1376 B.n686 B.n685 10.6151
R1377 B.n685 B.n684 10.6151
R1378 B.n684 B.n53 10.6151
R1379 B.n678 B.n53 10.6151
R1380 B.n678 B.n677 10.6151
R1381 B.n677 B.n676 10.6151
R1382 B.n676 B.n60 10.6151
R1383 B.n670 B.n60 10.6151
R1384 B.n670 B.n669 10.6151
R1385 B.n669 B.n668 10.6151
R1386 B.n668 B.n67 10.6151
R1387 B.n662 B.n67 10.6151
R1388 B.n662 B.n661 10.6151
R1389 B.n661 B.n660 10.6151
R1390 B.n660 B.n73 10.6151
R1391 B.n654 B.n73 10.6151
R1392 B.n654 B.n653 10.6151
R1393 B.n653 B.n652 10.6151
R1394 B.n652 B.n81 10.6151
R1395 B.n120 B.n119 10.6151
R1396 B.n123 B.n120 10.6151
R1397 B.n124 B.n123 10.6151
R1398 B.n127 B.n124 10.6151
R1399 B.n128 B.n127 10.6151
R1400 B.n131 B.n128 10.6151
R1401 B.n132 B.n131 10.6151
R1402 B.n135 B.n132 10.6151
R1403 B.n136 B.n135 10.6151
R1404 B.n139 B.n136 10.6151
R1405 B.n140 B.n139 10.6151
R1406 B.n143 B.n140 10.6151
R1407 B.n144 B.n143 10.6151
R1408 B.n147 B.n144 10.6151
R1409 B.n148 B.n147 10.6151
R1410 B.n151 B.n148 10.6151
R1411 B.n152 B.n151 10.6151
R1412 B.n155 B.n152 10.6151
R1413 B.n156 B.n155 10.6151
R1414 B.n159 B.n156 10.6151
R1415 B.n160 B.n159 10.6151
R1416 B.n164 B.n163 10.6151
R1417 B.n167 B.n164 10.6151
R1418 B.n168 B.n167 10.6151
R1419 B.n171 B.n168 10.6151
R1420 B.n172 B.n171 10.6151
R1421 B.n175 B.n172 10.6151
R1422 B.n176 B.n175 10.6151
R1423 B.n179 B.n176 10.6151
R1424 B.n180 B.n179 10.6151
R1425 B.n184 B.n183 10.6151
R1426 B.n187 B.n184 10.6151
R1427 B.n188 B.n187 10.6151
R1428 B.n191 B.n188 10.6151
R1429 B.n192 B.n191 10.6151
R1430 B.n195 B.n192 10.6151
R1431 B.n196 B.n195 10.6151
R1432 B.n199 B.n196 10.6151
R1433 B.n200 B.n199 10.6151
R1434 B.n203 B.n200 10.6151
R1435 B.n204 B.n203 10.6151
R1436 B.n207 B.n204 10.6151
R1437 B.n208 B.n207 10.6151
R1438 B.n211 B.n208 10.6151
R1439 B.n212 B.n211 10.6151
R1440 B.n215 B.n212 10.6151
R1441 B.n216 B.n215 10.6151
R1442 B.n219 B.n216 10.6151
R1443 B.n221 B.n219 10.6151
R1444 B.n222 B.n221 10.6151
R1445 B.n645 B.n222 10.6151
R1446 B.n404 B.n403 9.36635
R1447 B.n382 B.n381 9.36635
R1448 B.n160 B.n117 9.36635
R1449 B.n183 B.n114 9.36635
R1450 B.n742 B.n0 8.11757
R1451 B.n742 B.n1 8.11757
R1452 B.t8 B.n264 2.04796
R1453 B.t5 B.n44 2.04796
R1454 B.n403 B.n402 1.24928
R1455 B.n383 B.n382 1.24928
R1456 B.n163 B.n117 1.24928
R1457 B.n180 B.n114 1.24928
R1458 VP.n42 VP.n9 185.279
R1459 VP.n74 VP.n73 185.279
R1460 VP.n41 VP.n40 185.279
R1461 VP.n19 VP.n16 161.3
R1462 VP.n21 VP.n20 161.3
R1463 VP.n22 VP.n15 161.3
R1464 VP.n24 VP.n23 161.3
R1465 VP.n26 VP.n14 161.3
R1466 VP.n28 VP.n27 161.3
R1467 VP.n29 VP.n13 161.3
R1468 VP.n31 VP.n30 161.3
R1469 VP.n33 VP.n12 161.3
R1470 VP.n35 VP.n34 161.3
R1471 VP.n36 VP.n11 161.3
R1472 VP.n38 VP.n37 161.3
R1473 VP.n39 VP.n10 161.3
R1474 VP.n72 VP.n0 161.3
R1475 VP.n71 VP.n70 161.3
R1476 VP.n69 VP.n1 161.3
R1477 VP.n68 VP.n67 161.3
R1478 VP.n66 VP.n2 161.3
R1479 VP.n64 VP.n63 161.3
R1480 VP.n62 VP.n3 161.3
R1481 VP.n61 VP.n60 161.3
R1482 VP.n59 VP.n4 161.3
R1483 VP.n57 VP.n56 161.3
R1484 VP.n55 VP.n5 161.3
R1485 VP.n54 VP.n53 161.3
R1486 VP.n52 VP.n6 161.3
R1487 VP.n50 VP.n49 161.3
R1488 VP.n48 VP.n7 161.3
R1489 VP.n47 VP.n46 161.3
R1490 VP.n45 VP.n8 161.3
R1491 VP.n44 VP.n43 161.3
R1492 VP.n17 VP.t3 105.445
R1493 VP.n9 VP.t8 73.2377
R1494 VP.n51 VP.t4 73.2377
R1495 VP.n58 VP.t1 73.2377
R1496 VP.n65 VP.t0 73.2377
R1497 VP.n73 VP.t7 73.2377
R1498 VP.n40 VP.t5 73.2377
R1499 VP.n32 VP.t2 73.2377
R1500 VP.n25 VP.t9 73.2377
R1501 VP.n18 VP.t6 73.2377
R1502 VP.n53 VP.n5 56.5193
R1503 VP.n60 VP.n3 56.5193
R1504 VP.n27 VP.n13 56.5193
R1505 VP.n20 VP.n15 56.5193
R1506 VP.n18 VP.n17 51.0503
R1507 VP.n46 VP.n7 45.8354
R1508 VP.n67 VP.n1 45.8354
R1509 VP.n34 VP.n11 45.8354
R1510 VP.n42 VP.n41 43.671
R1511 VP.n46 VP.n45 35.1514
R1512 VP.n71 VP.n1 35.1514
R1513 VP.n38 VP.n11 35.1514
R1514 VP.n45 VP.n44 24.4675
R1515 VP.n50 VP.n7 24.4675
R1516 VP.n53 VP.n52 24.4675
R1517 VP.n57 VP.n5 24.4675
R1518 VP.n60 VP.n59 24.4675
R1519 VP.n64 VP.n3 24.4675
R1520 VP.n67 VP.n66 24.4675
R1521 VP.n72 VP.n71 24.4675
R1522 VP.n39 VP.n38 24.4675
R1523 VP.n31 VP.n13 24.4675
R1524 VP.n34 VP.n33 24.4675
R1525 VP.n24 VP.n15 24.4675
R1526 VP.n27 VP.n26 24.4675
R1527 VP.n20 VP.n19 24.4675
R1528 VP.n52 VP.n51 18.5954
R1529 VP.n65 VP.n64 18.5954
R1530 VP.n32 VP.n31 18.5954
R1531 VP.n19 VP.n18 18.5954
R1532 VP.n17 VP.n16 12.5362
R1533 VP.n58 VP.n57 12.234
R1534 VP.n59 VP.n58 12.234
R1535 VP.n25 VP.n24 12.234
R1536 VP.n26 VP.n25 12.234
R1537 VP.n51 VP.n50 5.87258
R1538 VP.n66 VP.n65 5.87258
R1539 VP.n33 VP.n32 5.87258
R1540 VP.n44 VP.n9 0.48984
R1541 VP.n73 VP.n72 0.48984
R1542 VP.n40 VP.n39 0.48984
R1543 VP.n21 VP.n16 0.189894
R1544 VP.n22 VP.n21 0.189894
R1545 VP.n23 VP.n22 0.189894
R1546 VP.n23 VP.n14 0.189894
R1547 VP.n28 VP.n14 0.189894
R1548 VP.n29 VP.n28 0.189894
R1549 VP.n30 VP.n29 0.189894
R1550 VP.n30 VP.n12 0.189894
R1551 VP.n35 VP.n12 0.189894
R1552 VP.n36 VP.n35 0.189894
R1553 VP.n37 VP.n36 0.189894
R1554 VP.n37 VP.n10 0.189894
R1555 VP.n41 VP.n10 0.189894
R1556 VP.n43 VP.n42 0.189894
R1557 VP.n43 VP.n8 0.189894
R1558 VP.n47 VP.n8 0.189894
R1559 VP.n48 VP.n47 0.189894
R1560 VP.n49 VP.n48 0.189894
R1561 VP.n49 VP.n6 0.189894
R1562 VP.n54 VP.n6 0.189894
R1563 VP.n55 VP.n54 0.189894
R1564 VP.n56 VP.n55 0.189894
R1565 VP.n56 VP.n4 0.189894
R1566 VP.n61 VP.n4 0.189894
R1567 VP.n62 VP.n61 0.189894
R1568 VP.n63 VP.n62 0.189894
R1569 VP.n63 VP.n2 0.189894
R1570 VP.n68 VP.n2 0.189894
R1571 VP.n69 VP.n68 0.189894
R1572 VP.n70 VP.n69 0.189894
R1573 VP.n70 VP.n0 0.189894
R1574 VP.n74 VP.n0 0.189894
R1575 VP VP.n74 0.0516364
R1576 VDD1.n1 VDD1.t6 76.1076
R1577 VDD1.n3 VDD1.t1 76.1066
R1578 VDD1.n5 VDD1.n4 71.9733
R1579 VDD1.n1 VDD1.n0 70.6516
R1580 VDD1.n3 VDD1.n2 70.6515
R1581 VDD1.n7 VDD1.n6 70.6507
R1582 VDD1.n7 VDD1.n5 38.6539
R1583 VDD1.n6 VDD1.t7 3.62024
R1584 VDD1.n6 VDD1.t4 3.62024
R1585 VDD1.n0 VDD1.t3 3.62024
R1586 VDD1.n0 VDD1.t0 3.62024
R1587 VDD1.n4 VDD1.t9 3.62024
R1588 VDD1.n4 VDD1.t2 3.62024
R1589 VDD1.n2 VDD1.t5 3.62024
R1590 VDD1.n2 VDD1.t8 3.62024
R1591 VDD1 VDD1.n7 1.31947
R1592 VDD1 VDD1.n1 0.517741
R1593 VDD1.n5 VDD1.n3 0.404206
C0 VDD2 VDD1 1.65261f
C1 VN VTAIL 5.46002f
C2 VDD2 VTAIL 6.96593f
C3 VN VP 6.01122f
C4 VDD2 VP 0.484679f
C5 VDD1 VTAIL 6.91935f
C6 VP VDD1 5.05264f
C7 VN VDD2 4.72575f
C8 VN VDD1 0.151473f
C9 VP VTAIL 5.47424f
C10 VDD2 B 5.085109f
C11 VDD1 B 5.077453f
C12 VTAIL B 4.698694f
C13 VN B 13.666069f
C14 VP B 12.189775f
C15 VDD1.t6 B 1.06725f
C16 VDD1.t3 B 0.100032f
C17 VDD1.t0 B 0.100032f
C18 VDD1.n0 B 0.834565f
C19 VDD1.n1 B 0.71415f
C20 VDD1.t1 B 1.06725f
C21 VDD1.t5 B 0.100032f
C22 VDD1.t8 B 0.100032f
C23 VDD1.n2 B 0.834562f
C24 VDD1.n3 B 0.707015f
C25 VDD1.t9 B 0.100032f
C26 VDD1.t2 B 0.100032f
C27 VDD1.n4 B 0.842301f
C28 VDD1.n5 B 2.01613f
C29 VDD1.t7 B 0.100032f
C30 VDD1.t4 B 0.100032f
C31 VDD1.n6 B 0.834563f
C32 VDD1.n7 B 2.14504f
C33 VP.n0 B 0.030249f
C34 VP.t7 B 0.783797f
C35 VP.n1 B 0.025651f
C36 VP.n2 B 0.030249f
C37 VP.t0 B 0.783797f
C38 VP.n3 B 0.038682f
C39 VP.n4 B 0.030249f
C40 VP.t1 B 0.783797f
C41 VP.n5 B 0.04964f
C42 VP.n6 B 0.030249f
C43 VP.t4 B 0.783797f
C44 VP.n7 B 0.057933f
C45 VP.n8 B 0.030249f
C46 VP.t8 B 0.783797f
C47 VP.n9 B 0.370157f
C48 VP.n10 B 0.030249f
C49 VP.t5 B 0.783797f
C50 VP.n11 B 0.025651f
C51 VP.n12 B 0.030249f
C52 VP.t2 B 0.783797f
C53 VP.n13 B 0.038682f
C54 VP.n14 B 0.030249f
C55 VP.t9 B 0.783797f
C56 VP.n15 B 0.04964f
C57 VP.n16 B 0.221262f
C58 VP.t6 B 0.783797f
C59 VP.t3 B 0.920766f
C60 VP.n17 B 0.373524f
C61 VP.n18 B 0.380714f
C62 VP.n19 B 0.049696f
C63 VP.n20 B 0.038682f
C64 VP.n21 B 0.030249f
C65 VP.n22 B 0.030249f
C66 VP.n23 B 0.030249f
C67 VP.n24 B 0.04246f
C68 VP.n25 B 0.306053f
C69 VP.n26 B 0.04246f
C70 VP.n27 B 0.04964f
C71 VP.n28 B 0.030249f
C72 VP.n29 B 0.030249f
C73 VP.n30 B 0.030249f
C74 VP.n31 B 0.049696f
C75 VP.n32 B 0.306053f
C76 VP.n33 B 0.035223f
C77 VP.n34 B 0.057933f
C78 VP.n35 B 0.030249f
C79 VP.n36 B 0.030249f
C80 VP.n37 B 0.030249f
C81 VP.n38 B 0.061114f
C82 VP.n39 B 0.0291f
C83 VP.n40 B 0.370157f
C84 VP.n41 B 1.34087f
C85 VP.n42 B 1.36577f
C86 VP.n43 B 0.030249f
C87 VP.n44 B 0.0291f
C88 VP.n45 B 0.061114f
C89 VP.n46 B 0.025651f
C90 VP.n47 B 0.030249f
C91 VP.n48 B 0.030249f
C92 VP.n49 B 0.030249f
C93 VP.n50 B 0.035223f
C94 VP.n51 B 0.306053f
C95 VP.n52 B 0.049696f
C96 VP.n53 B 0.038682f
C97 VP.n54 B 0.030249f
C98 VP.n55 B 0.030249f
C99 VP.n56 B 0.030249f
C100 VP.n57 B 0.04246f
C101 VP.n58 B 0.306053f
C102 VP.n59 B 0.04246f
C103 VP.n60 B 0.04964f
C104 VP.n61 B 0.030249f
C105 VP.n62 B 0.030249f
C106 VP.n63 B 0.030249f
C107 VP.n64 B 0.049696f
C108 VP.n65 B 0.306053f
C109 VP.n66 B 0.035223f
C110 VP.n67 B 0.057933f
C111 VP.n68 B 0.030249f
C112 VP.n69 B 0.030249f
C113 VP.n70 B 0.030249f
C114 VP.n71 B 0.061114f
C115 VP.n72 B 0.0291f
C116 VP.n73 B 0.370157f
C117 VP.n74 B 0.032971f
C118 VTAIL.t13 B 0.121307f
C119 VTAIL.t19 B 0.121307f
C120 VTAIL.n0 B 0.9477f
C121 VTAIL.n1 B 0.495122f
C122 VTAIL.t1 B 1.20581f
C123 VTAIL.n2 B 0.604101f
C124 VTAIL.t9 B 0.121307f
C125 VTAIL.t3 B 0.121307f
C126 VTAIL.n3 B 0.9477f
C127 VTAIL.n4 B 0.571907f
C128 VTAIL.t4 B 0.121307f
C129 VTAIL.t8 B 0.121307f
C130 VTAIL.n5 B 0.9477f
C131 VTAIL.n6 B 1.54558f
C132 VTAIL.t16 B 0.121307f
C133 VTAIL.t10 B 0.121307f
C134 VTAIL.n7 B 0.947705f
C135 VTAIL.n8 B 1.54557f
C136 VTAIL.t17 B 0.121307f
C137 VTAIL.t11 B 0.121307f
C138 VTAIL.n9 B 0.947705f
C139 VTAIL.n10 B 0.571903f
C140 VTAIL.t14 B 1.20581f
C141 VTAIL.n11 B 0.6041f
C142 VTAIL.t7 B 0.121307f
C143 VTAIL.t0 B 0.121307f
C144 VTAIL.n12 B 0.947705f
C145 VTAIL.n13 B 0.531366f
C146 VTAIL.t6 B 0.121307f
C147 VTAIL.t5 B 0.121307f
C148 VTAIL.n14 B 0.947705f
C149 VTAIL.n15 B 0.571903f
C150 VTAIL.t2 B 1.2058f
C151 VTAIL.n16 B 1.45227f
C152 VTAIL.t12 B 1.20581f
C153 VTAIL.n17 B 1.45226f
C154 VTAIL.t18 B 0.121307f
C155 VTAIL.t15 B 0.121307f
C156 VTAIL.n18 B 0.9477f
C157 VTAIL.n19 B 0.442113f
C158 VDD2.t8 B 1.04803f
C159 VDD2.t0 B 0.098231f
C160 VDD2.t4 B 0.098231f
C161 VDD2.n0 B 0.819536f
C162 VDD2.n1 B 0.694284f
C163 VDD2.t3 B 0.098231f
C164 VDD2.t9 B 0.098231f
C165 VDD2.n2 B 0.827135f
C166 VDD2.n3 B 1.88939f
C167 VDD2.t6 B 1.03923f
C168 VDD2.n4 B 2.06455f
C169 VDD2.t5 B 0.098231f
C170 VDD2.t1 B 0.098231f
C171 VDD2.n5 B 0.819538f
C172 VDD2.n6 B 0.345302f
C173 VDD2.t2 B 0.098231f
C174 VDD2.t7 B 0.098231f
C175 VDD2.n7 B 0.827108f
C176 VN.n0 B 0.029444f
C177 VN.t7 B 0.762956f
C178 VN.n1 B 0.024968f
C179 VN.n2 B 0.029444f
C180 VN.t4 B 0.762956f
C181 VN.n3 B 0.037653f
C182 VN.n4 B 0.029444f
C183 VN.t1 B 0.762956f
C184 VN.n5 B 0.04832f
C185 VN.n6 B 0.215378f
C186 VN.t0 B 0.762956f
C187 VN.t6 B 0.896283f
C188 VN.n7 B 0.363592f
C189 VN.n8 B 0.370591f
C190 VN.n9 B 0.048375f
C191 VN.n10 B 0.037653f
C192 VN.n11 B 0.029444f
C193 VN.n12 B 0.029444f
C194 VN.n13 B 0.029444f
C195 VN.n14 B 0.041331f
C196 VN.n15 B 0.297915f
C197 VN.n16 B 0.041331f
C198 VN.n17 B 0.04832f
C199 VN.n18 B 0.029444f
C200 VN.n19 B 0.029444f
C201 VN.n20 B 0.029444f
C202 VN.n21 B 0.048375f
C203 VN.n22 B 0.297915f
C204 VN.n23 B 0.034286f
C205 VN.n24 B 0.056393f
C206 VN.n25 B 0.029444f
C207 VN.n26 B 0.029444f
C208 VN.n27 B 0.029444f
C209 VN.n28 B 0.059489f
C210 VN.n29 B 0.028326f
C211 VN.n30 B 0.360315f
C212 VN.n31 B 0.032094f
C213 VN.n32 B 0.029444f
C214 VN.t3 B 0.762956f
C215 VN.n33 B 0.024968f
C216 VN.n34 B 0.029444f
C217 VN.t9 B 0.762956f
C218 VN.n35 B 0.037653f
C219 VN.n36 B 0.029444f
C220 VN.t2 B 0.762956f
C221 VN.n37 B 0.04832f
C222 VN.n38 B 0.215378f
C223 VN.t8 B 0.762956f
C224 VN.t5 B 0.896283f
C225 VN.n39 B 0.363592f
C226 VN.n40 B 0.370591f
C227 VN.n41 B 0.048375f
C228 VN.n42 B 0.037653f
C229 VN.n43 B 0.029444f
C230 VN.n44 B 0.029444f
C231 VN.n45 B 0.029444f
C232 VN.n46 B 0.041331f
C233 VN.n47 B 0.297915f
C234 VN.n48 B 0.041331f
C235 VN.n49 B 0.04832f
C236 VN.n50 B 0.029444f
C237 VN.n51 B 0.029444f
C238 VN.n52 B 0.029444f
C239 VN.n53 B 0.048375f
C240 VN.n54 B 0.297915f
C241 VN.n55 B 0.034286f
C242 VN.n56 B 0.056393f
C243 VN.n57 B 0.029444f
C244 VN.n58 B 0.029444f
C245 VN.n59 B 0.029444f
C246 VN.n60 B 0.059489f
C247 VN.n61 B 0.028326f
C248 VN.n62 B 0.360315f
C249 VN.n63 B 1.3245f
.ends

