* NGSPICE file created from diff_pair_sample_1267.ext - technology: sky130A

.subckt diff_pair_sample_1267 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=6.357 ps=33.38 w=16.3 l=3.47
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=0 ps=0 w=16.3 l=3.47
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=6.357 ps=33.38 w=16.3 l=3.47
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=0 ps=0 w=16.3 l=3.47
X4 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=6.357 ps=33.38 w=16.3 l=3.47
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=0 ps=0 w=16.3 l=3.47
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=6.357 ps=33.38 w=16.3 l=3.47
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.357 pd=33.38 as=0 ps=0 w=16.3 l=3.47
R0 VN VN.t1 202.181
R1 VN VN.t0 152.579
R2 VTAIL.n354 VTAIL.n270 289.615
R3 VTAIL.n84 VTAIL.n0 289.615
R4 VTAIL.n264 VTAIL.n180 289.615
R5 VTAIL.n174 VTAIL.n90 289.615
R6 VTAIL.n298 VTAIL.n297 185
R7 VTAIL.n303 VTAIL.n302 185
R8 VTAIL.n305 VTAIL.n304 185
R9 VTAIL.n294 VTAIL.n293 185
R10 VTAIL.n311 VTAIL.n310 185
R11 VTAIL.n313 VTAIL.n312 185
R12 VTAIL.n290 VTAIL.n289 185
R13 VTAIL.n319 VTAIL.n318 185
R14 VTAIL.n321 VTAIL.n320 185
R15 VTAIL.n286 VTAIL.n285 185
R16 VTAIL.n327 VTAIL.n326 185
R17 VTAIL.n329 VTAIL.n328 185
R18 VTAIL.n282 VTAIL.n281 185
R19 VTAIL.n335 VTAIL.n334 185
R20 VTAIL.n337 VTAIL.n336 185
R21 VTAIL.n278 VTAIL.n277 185
R22 VTAIL.n344 VTAIL.n343 185
R23 VTAIL.n345 VTAIL.n276 185
R24 VTAIL.n347 VTAIL.n346 185
R25 VTAIL.n274 VTAIL.n273 185
R26 VTAIL.n353 VTAIL.n352 185
R27 VTAIL.n355 VTAIL.n354 185
R28 VTAIL.n28 VTAIL.n27 185
R29 VTAIL.n33 VTAIL.n32 185
R30 VTAIL.n35 VTAIL.n34 185
R31 VTAIL.n24 VTAIL.n23 185
R32 VTAIL.n41 VTAIL.n40 185
R33 VTAIL.n43 VTAIL.n42 185
R34 VTAIL.n20 VTAIL.n19 185
R35 VTAIL.n49 VTAIL.n48 185
R36 VTAIL.n51 VTAIL.n50 185
R37 VTAIL.n16 VTAIL.n15 185
R38 VTAIL.n57 VTAIL.n56 185
R39 VTAIL.n59 VTAIL.n58 185
R40 VTAIL.n12 VTAIL.n11 185
R41 VTAIL.n65 VTAIL.n64 185
R42 VTAIL.n67 VTAIL.n66 185
R43 VTAIL.n8 VTAIL.n7 185
R44 VTAIL.n74 VTAIL.n73 185
R45 VTAIL.n75 VTAIL.n6 185
R46 VTAIL.n77 VTAIL.n76 185
R47 VTAIL.n4 VTAIL.n3 185
R48 VTAIL.n83 VTAIL.n82 185
R49 VTAIL.n85 VTAIL.n84 185
R50 VTAIL.n265 VTAIL.n264 185
R51 VTAIL.n263 VTAIL.n262 185
R52 VTAIL.n184 VTAIL.n183 185
R53 VTAIL.n257 VTAIL.n256 185
R54 VTAIL.n255 VTAIL.n186 185
R55 VTAIL.n254 VTAIL.n253 185
R56 VTAIL.n189 VTAIL.n187 185
R57 VTAIL.n248 VTAIL.n247 185
R58 VTAIL.n246 VTAIL.n245 185
R59 VTAIL.n193 VTAIL.n192 185
R60 VTAIL.n240 VTAIL.n239 185
R61 VTAIL.n238 VTAIL.n237 185
R62 VTAIL.n197 VTAIL.n196 185
R63 VTAIL.n232 VTAIL.n231 185
R64 VTAIL.n230 VTAIL.n229 185
R65 VTAIL.n201 VTAIL.n200 185
R66 VTAIL.n224 VTAIL.n223 185
R67 VTAIL.n222 VTAIL.n221 185
R68 VTAIL.n205 VTAIL.n204 185
R69 VTAIL.n216 VTAIL.n215 185
R70 VTAIL.n214 VTAIL.n213 185
R71 VTAIL.n209 VTAIL.n208 185
R72 VTAIL.n175 VTAIL.n174 185
R73 VTAIL.n173 VTAIL.n172 185
R74 VTAIL.n94 VTAIL.n93 185
R75 VTAIL.n167 VTAIL.n166 185
R76 VTAIL.n165 VTAIL.n96 185
R77 VTAIL.n164 VTAIL.n163 185
R78 VTAIL.n99 VTAIL.n97 185
R79 VTAIL.n158 VTAIL.n157 185
R80 VTAIL.n156 VTAIL.n155 185
R81 VTAIL.n103 VTAIL.n102 185
R82 VTAIL.n150 VTAIL.n149 185
R83 VTAIL.n148 VTAIL.n147 185
R84 VTAIL.n107 VTAIL.n106 185
R85 VTAIL.n142 VTAIL.n141 185
R86 VTAIL.n140 VTAIL.n139 185
R87 VTAIL.n111 VTAIL.n110 185
R88 VTAIL.n134 VTAIL.n133 185
R89 VTAIL.n132 VTAIL.n131 185
R90 VTAIL.n115 VTAIL.n114 185
R91 VTAIL.n126 VTAIL.n125 185
R92 VTAIL.n124 VTAIL.n123 185
R93 VTAIL.n119 VTAIL.n118 185
R94 VTAIL.n299 VTAIL.t3 147.659
R95 VTAIL.n29 VTAIL.t1 147.659
R96 VTAIL.n210 VTAIL.t0 147.659
R97 VTAIL.n120 VTAIL.t2 147.659
R98 VTAIL.n303 VTAIL.n297 104.615
R99 VTAIL.n304 VTAIL.n303 104.615
R100 VTAIL.n304 VTAIL.n293 104.615
R101 VTAIL.n311 VTAIL.n293 104.615
R102 VTAIL.n312 VTAIL.n311 104.615
R103 VTAIL.n312 VTAIL.n289 104.615
R104 VTAIL.n319 VTAIL.n289 104.615
R105 VTAIL.n320 VTAIL.n319 104.615
R106 VTAIL.n320 VTAIL.n285 104.615
R107 VTAIL.n327 VTAIL.n285 104.615
R108 VTAIL.n328 VTAIL.n327 104.615
R109 VTAIL.n328 VTAIL.n281 104.615
R110 VTAIL.n335 VTAIL.n281 104.615
R111 VTAIL.n336 VTAIL.n335 104.615
R112 VTAIL.n336 VTAIL.n277 104.615
R113 VTAIL.n344 VTAIL.n277 104.615
R114 VTAIL.n345 VTAIL.n344 104.615
R115 VTAIL.n346 VTAIL.n345 104.615
R116 VTAIL.n346 VTAIL.n273 104.615
R117 VTAIL.n353 VTAIL.n273 104.615
R118 VTAIL.n354 VTAIL.n353 104.615
R119 VTAIL.n33 VTAIL.n27 104.615
R120 VTAIL.n34 VTAIL.n33 104.615
R121 VTAIL.n34 VTAIL.n23 104.615
R122 VTAIL.n41 VTAIL.n23 104.615
R123 VTAIL.n42 VTAIL.n41 104.615
R124 VTAIL.n42 VTAIL.n19 104.615
R125 VTAIL.n49 VTAIL.n19 104.615
R126 VTAIL.n50 VTAIL.n49 104.615
R127 VTAIL.n50 VTAIL.n15 104.615
R128 VTAIL.n57 VTAIL.n15 104.615
R129 VTAIL.n58 VTAIL.n57 104.615
R130 VTAIL.n58 VTAIL.n11 104.615
R131 VTAIL.n65 VTAIL.n11 104.615
R132 VTAIL.n66 VTAIL.n65 104.615
R133 VTAIL.n66 VTAIL.n7 104.615
R134 VTAIL.n74 VTAIL.n7 104.615
R135 VTAIL.n75 VTAIL.n74 104.615
R136 VTAIL.n76 VTAIL.n75 104.615
R137 VTAIL.n76 VTAIL.n3 104.615
R138 VTAIL.n83 VTAIL.n3 104.615
R139 VTAIL.n84 VTAIL.n83 104.615
R140 VTAIL.n264 VTAIL.n263 104.615
R141 VTAIL.n263 VTAIL.n183 104.615
R142 VTAIL.n256 VTAIL.n183 104.615
R143 VTAIL.n256 VTAIL.n255 104.615
R144 VTAIL.n255 VTAIL.n254 104.615
R145 VTAIL.n254 VTAIL.n187 104.615
R146 VTAIL.n247 VTAIL.n187 104.615
R147 VTAIL.n247 VTAIL.n246 104.615
R148 VTAIL.n246 VTAIL.n192 104.615
R149 VTAIL.n239 VTAIL.n192 104.615
R150 VTAIL.n239 VTAIL.n238 104.615
R151 VTAIL.n238 VTAIL.n196 104.615
R152 VTAIL.n231 VTAIL.n196 104.615
R153 VTAIL.n231 VTAIL.n230 104.615
R154 VTAIL.n230 VTAIL.n200 104.615
R155 VTAIL.n223 VTAIL.n200 104.615
R156 VTAIL.n223 VTAIL.n222 104.615
R157 VTAIL.n222 VTAIL.n204 104.615
R158 VTAIL.n215 VTAIL.n204 104.615
R159 VTAIL.n215 VTAIL.n214 104.615
R160 VTAIL.n214 VTAIL.n208 104.615
R161 VTAIL.n174 VTAIL.n173 104.615
R162 VTAIL.n173 VTAIL.n93 104.615
R163 VTAIL.n166 VTAIL.n93 104.615
R164 VTAIL.n166 VTAIL.n165 104.615
R165 VTAIL.n165 VTAIL.n164 104.615
R166 VTAIL.n164 VTAIL.n97 104.615
R167 VTAIL.n157 VTAIL.n97 104.615
R168 VTAIL.n157 VTAIL.n156 104.615
R169 VTAIL.n156 VTAIL.n102 104.615
R170 VTAIL.n149 VTAIL.n102 104.615
R171 VTAIL.n149 VTAIL.n148 104.615
R172 VTAIL.n148 VTAIL.n106 104.615
R173 VTAIL.n141 VTAIL.n106 104.615
R174 VTAIL.n141 VTAIL.n140 104.615
R175 VTAIL.n140 VTAIL.n110 104.615
R176 VTAIL.n133 VTAIL.n110 104.615
R177 VTAIL.n133 VTAIL.n132 104.615
R178 VTAIL.n132 VTAIL.n114 104.615
R179 VTAIL.n125 VTAIL.n114 104.615
R180 VTAIL.n125 VTAIL.n124 104.615
R181 VTAIL.n124 VTAIL.n118 104.615
R182 VTAIL.t3 VTAIL.n297 52.3082
R183 VTAIL.t1 VTAIL.n27 52.3082
R184 VTAIL.t0 VTAIL.n208 52.3082
R185 VTAIL.t2 VTAIL.n118 52.3082
R186 VTAIL.n359 VTAIL.n358 36.452
R187 VTAIL.n89 VTAIL.n88 36.452
R188 VTAIL.n269 VTAIL.n268 36.452
R189 VTAIL.n179 VTAIL.n178 36.452
R190 VTAIL.n179 VTAIL.n89 32.9703
R191 VTAIL.n359 VTAIL.n269 29.6945
R192 VTAIL.n299 VTAIL.n298 15.6677
R193 VTAIL.n29 VTAIL.n28 15.6677
R194 VTAIL.n210 VTAIL.n209 15.6677
R195 VTAIL.n120 VTAIL.n119 15.6677
R196 VTAIL.n347 VTAIL.n276 13.1884
R197 VTAIL.n77 VTAIL.n6 13.1884
R198 VTAIL.n257 VTAIL.n186 13.1884
R199 VTAIL.n167 VTAIL.n96 13.1884
R200 VTAIL.n302 VTAIL.n301 12.8005
R201 VTAIL.n343 VTAIL.n342 12.8005
R202 VTAIL.n348 VTAIL.n274 12.8005
R203 VTAIL.n32 VTAIL.n31 12.8005
R204 VTAIL.n73 VTAIL.n72 12.8005
R205 VTAIL.n78 VTAIL.n4 12.8005
R206 VTAIL.n258 VTAIL.n184 12.8005
R207 VTAIL.n253 VTAIL.n188 12.8005
R208 VTAIL.n213 VTAIL.n212 12.8005
R209 VTAIL.n168 VTAIL.n94 12.8005
R210 VTAIL.n163 VTAIL.n98 12.8005
R211 VTAIL.n123 VTAIL.n122 12.8005
R212 VTAIL.n305 VTAIL.n296 12.0247
R213 VTAIL.n341 VTAIL.n278 12.0247
R214 VTAIL.n352 VTAIL.n351 12.0247
R215 VTAIL.n35 VTAIL.n26 12.0247
R216 VTAIL.n71 VTAIL.n8 12.0247
R217 VTAIL.n82 VTAIL.n81 12.0247
R218 VTAIL.n262 VTAIL.n261 12.0247
R219 VTAIL.n252 VTAIL.n189 12.0247
R220 VTAIL.n216 VTAIL.n207 12.0247
R221 VTAIL.n172 VTAIL.n171 12.0247
R222 VTAIL.n162 VTAIL.n99 12.0247
R223 VTAIL.n126 VTAIL.n117 12.0247
R224 VTAIL.n306 VTAIL.n294 11.249
R225 VTAIL.n338 VTAIL.n337 11.249
R226 VTAIL.n355 VTAIL.n272 11.249
R227 VTAIL.n36 VTAIL.n24 11.249
R228 VTAIL.n68 VTAIL.n67 11.249
R229 VTAIL.n85 VTAIL.n2 11.249
R230 VTAIL.n265 VTAIL.n182 11.249
R231 VTAIL.n249 VTAIL.n248 11.249
R232 VTAIL.n217 VTAIL.n205 11.249
R233 VTAIL.n175 VTAIL.n92 11.249
R234 VTAIL.n159 VTAIL.n158 11.249
R235 VTAIL.n127 VTAIL.n115 11.249
R236 VTAIL.n310 VTAIL.n309 10.4732
R237 VTAIL.n334 VTAIL.n280 10.4732
R238 VTAIL.n356 VTAIL.n270 10.4732
R239 VTAIL.n40 VTAIL.n39 10.4732
R240 VTAIL.n64 VTAIL.n10 10.4732
R241 VTAIL.n86 VTAIL.n0 10.4732
R242 VTAIL.n266 VTAIL.n180 10.4732
R243 VTAIL.n245 VTAIL.n191 10.4732
R244 VTAIL.n221 VTAIL.n220 10.4732
R245 VTAIL.n176 VTAIL.n90 10.4732
R246 VTAIL.n155 VTAIL.n101 10.4732
R247 VTAIL.n131 VTAIL.n130 10.4732
R248 VTAIL.n313 VTAIL.n292 9.69747
R249 VTAIL.n333 VTAIL.n282 9.69747
R250 VTAIL.n43 VTAIL.n22 9.69747
R251 VTAIL.n63 VTAIL.n12 9.69747
R252 VTAIL.n244 VTAIL.n193 9.69747
R253 VTAIL.n224 VTAIL.n203 9.69747
R254 VTAIL.n154 VTAIL.n103 9.69747
R255 VTAIL.n134 VTAIL.n113 9.69747
R256 VTAIL.n358 VTAIL.n357 9.45567
R257 VTAIL.n88 VTAIL.n87 9.45567
R258 VTAIL.n268 VTAIL.n267 9.45567
R259 VTAIL.n178 VTAIL.n177 9.45567
R260 VTAIL.n357 VTAIL.n356 9.3005
R261 VTAIL.n272 VTAIL.n271 9.3005
R262 VTAIL.n351 VTAIL.n350 9.3005
R263 VTAIL.n349 VTAIL.n348 9.3005
R264 VTAIL.n288 VTAIL.n287 9.3005
R265 VTAIL.n317 VTAIL.n316 9.3005
R266 VTAIL.n315 VTAIL.n314 9.3005
R267 VTAIL.n292 VTAIL.n291 9.3005
R268 VTAIL.n309 VTAIL.n308 9.3005
R269 VTAIL.n307 VTAIL.n306 9.3005
R270 VTAIL.n296 VTAIL.n295 9.3005
R271 VTAIL.n301 VTAIL.n300 9.3005
R272 VTAIL.n323 VTAIL.n322 9.3005
R273 VTAIL.n325 VTAIL.n324 9.3005
R274 VTAIL.n284 VTAIL.n283 9.3005
R275 VTAIL.n331 VTAIL.n330 9.3005
R276 VTAIL.n333 VTAIL.n332 9.3005
R277 VTAIL.n280 VTAIL.n279 9.3005
R278 VTAIL.n339 VTAIL.n338 9.3005
R279 VTAIL.n341 VTAIL.n340 9.3005
R280 VTAIL.n342 VTAIL.n275 9.3005
R281 VTAIL.n87 VTAIL.n86 9.3005
R282 VTAIL.n2 VTAIL.n1 9.3005
R283 VTAIL.n81 VTAIL.n80 9.3005
R284 VTAIL.n79 VTAIL.n78 9.3005
R285 VTAIL.n18 VTAIL.n17 9.3005
R286 VTAIL.n47 VTAIL.n46 9.3005
R287 VTAIL.n45 VTAIL.n44 9.3005
R288 VTAIL.n22 VTAIL.n21 9.3005
R289 VTAIL.n39 VTAIL.n38 9.3005
R290 VTAIL.n37 VTAIL.n36 9.3005
R291 VTAIL.n26 VTAIL.n25 9.3005
R292 VTAIL.n31 VTAIL.n30 9.3005
R293 VTAIL.n53 VTAIL.n52 9.3005
R294 VTAIL.n55 VTAIL.n54 9.3005
R295 VTAIL.n14 VTAIL.n13 9.3005
R296 VTAIL.n61 VTAIL.n60 9.3005
R297 VTAIL.n63 VTAIL.n62 9.3005
R298 VTAIL.n10 VTAIL.n9 9.3005
R299 VTAIL.n69 VTAIL.n68 9.3005
R300 VTAIL.n71 VTAIL.n70 9.3005
R301 VTAIL.n72 VTAIL.n5 9.3005
R302 VTAIL.n236 VTAIL.n235 9.3005
R303 VTAIL.n195 VTAIL.n194 9.3005
R304 VTAIL.n242 VTAIL.n241 9.3005
R305 VTAIL.n244 VTAIL.n243 9.3005
R306 VTAIL.n191 VTAIL.n190 9.3005
R307 VTAIL.n250 VTAIL.n249 9.3005
R308 VTAIL.n252 VTAIL.n251 9.3005
R309 VTAIL.n188 VTAIL.n185 9.3005
R310 VTAIL.n267 VTAIL.n266 9.3005
R311 VTAIL.n182 VTAIL.n181 9.3005
R312 VTAIL.n261 VTAIL.n260 9.3005
R313 VTAIL.n259 VTAIL.n258 9.3005
R314 VTAIL.n234 VTAIL.n233 9.3005
R315 VTAIL.n199 VTAIL.n198 9.3005
R316 VTAIL.n228 VTAIL.n227 9.3005
R317 VTAIL.n226 VTAIL.n225 9.3005
R318 VTAIL.n203 VTAIL.n202 9.3005
R319 VTAIL.n220 VTAIL.n219 9.3005
R320 VTAIL.n218 VTAIL.n217 9.3005
R321 VTAIL.n207 VTAIL.n206 9.3005
R322 VTAIL.n212 VTAIL.n211 9.3005
R323 VTAIL.n146 VTAIL.n145 9.3005
R324 VTAIL.n105 VTAIL.n104 9.3005
R325 VTAIL.n152 VTAIL.n151 9.3005
R326 VTAIL.n154 VTAIL.n153 9.3005
R327 VTAIL.n101 VTAIL.n100 9.3005
R328 VTAIL.n160 VTAIL.n159 9.3005
R329 VTAIL.n162 VTAIL.n161 9.3005
R330 VTAIL.n98 VTAIL.n95 9.3005
R331 VTAIL.n177 VTAIL.n176 9.3005
R332 VTAIL.n92 VTAIL.n91 9.3005
R333 VTAIL.n171 VTAIL.n170 9.3005
R334 VTAIL.n169 VTAIL.n168 9.3005
R335 VTAIL.n144 VTAIL.n143 9.3005
R336 VTAIL.n109 VTAIL.n108 9.3005
R337 VTAIL.n138 VTAIL.n137 9.3005
R338 VTAIL.n136 VTAIL.n135 9.3005
R339 VTAIL.n113 VTAIL.n112 9.3005
R340 VTAIL.n130 VTAIL.n129 9.3005
R341 VTAIL.n128 VTAIL.n127 9.3005
R342 VTAIL.n117 VTAIL.n116 9.3005
R343 VTAIL.n122 VTAIL.n121 9.3005
R344 VTAIL.n314 VTAIL.n290 8.92171
R345 VTAIL.n330 VTAIL.n329 8.92171
R346 VTAIL.n44 VTAIL.n20 8.92171
R347 VTAIL.n60 VTAIL.n59 8.92171
R348 VTAIL.n241 VTAIL.n240 8.92171
R349 VTAIL.n225 VTAIL.n201 8.92171
R350 VTAIL.n151 VTAIL.n150 8.92171
R351 VTAIL.n135 VTAIL.n111 8.92171
R352 VTAIL.n318 VTAIL.n317 8.14595
R353 VTAIL.n326 VTAIL.n284 8.14595
R354 VTAIL.n48 VTAIL.n47 8.14595
R355 VTAIL.n56 VTAIL.n14 8.14595
R356 VTAIL.n237 VTAIL.n195 8.14595
R357 VTAIL.n229 VTAIL.n228 8.14595
R358 VTAIL.n147 VTAIL.n105 8.14595
R359 VTAIL.n139 VTAIL.n138 8.14595
R360 VTAIL.n321 VTAIL.n288 7.3702
R361 VTAIL.n325 VTAIL.n286 7.3702
R362 VTAIL.n51 VTAIL.n18 7.3702
R363 VTAIL.n55 VTAIL.n16 7.3702
R364 VTAIL.n236 VTAIL.n197 7.3702
R365 VTAIL.n232 VTAIL.n199 7.3702
R366 VTAIL.n146 VTAIL.n107 7.3702
R367 VTAIL.n142 VTAIL.n109 7.3702
R368 VTAIL.n322 VTAIL.n321 6.59444
R369 VTAIL.n322 VTAIL.n286 6.59444
R370 VTAIL.n52 VTAIL.n51 6.59444
R371 VTAIL.n52 VTAIL.n16 6.59444
R372 VTAIL.n233 VTAIL.n197 6.59444
R373 VTAIL.n233 VTAIL.n232 6.59444
R374 VTAIL.n143 VTAIL.n107 6.59444
R375 VTAIL.n143 VTAIL.n142 6.59444
R376 VTAIL.n318 VTAIL.n288 5.81868
R377 VTAIL.n326 VTAIL.n325 5.81868
R378 VTAIL.n48 VTAIL.n18 5.81868
R379 VTAIL.n56 VTAIL.n55 5.81868
R380 VTAIL.n237 VTAIL.n236 5.81868
R381 VTAIL.n229 VTAIL.n199 5.81868
R382 VTAIL.n147 VTAIL.n146 5.81868
R383 VTAIL.n139 VTAIL.n109 5.81868
R384 VTAIL.n317 VTAIL.n290 5.04292
R385 VTAIL.n329 VTAIL.n284 5.04292
R386 VTAIL.n47 VTAIL.n20 5.04292
R387 VTAIL.n59 VTAIL.n14 5.04292
R388 VTAIL.n240 VTAIL.n195 5.04292
R389 VTAIL.n228 VTAIL.n201 5.04292
R390 VTAIL.n150 VTAIL.n105 5.04292
R391 VTAIL.n138 VTAIL.n111 5.04292
R392 VTAIL.n300 VTAIL.n299 4.38563
R393 VTAIL.n30 VTAIL.n29 4.38563
R394 VTAIL.n211 VTAIL.n210 4.38563
R395 VTAIL.n121 VTAIL.n120 4.38563
R396 VTAIL.n314 VTAIL.n313 4.26717
R397 VTAIL.n330 VTAIL.n282 4.26717
R398 VTAIL.n44 VTAIL.n43 4.26717
R399 VTAIL.n60 VTAIL.n12 4.26717
R400 VTAIL.n241 VTAIL.n193 4.26717
R401 VTAIL.n225 VTAIL.n224 4.26717
R402 VTAIL.n151 VTAIL.n103 4.26717
R403 VTAIL.n135 VTAIL.n134 4.26717
R404 VTAIL.n310 VTAIL.n292 3.49141
R405 VTAIL.n334 VTAIL.n333 3.49141
R406 VTAIL.n358 VTAIL.n270 3.49141
R407 VTAIL.n40 VTAIL.n22 3.49141
R408 VTAIL.n64 VTAIL.n63 3.49141
R409 VTAIL.n88 VTAIL.n0 3.49141
R410 VTAIL.n268 VTAIL.n180 3.49141
R411 VTAIL.n245 VTAIL.n244 3.49141
R412 VTAIL.n221 VTAIL.n203 3.49141
R413 VTAIL.n178 VTAIL.n90 3.49141
R414 VTAIL.n155 VTAIL.n154 3.49141
R415 VTAIL.n131 VTAIL.n113 3.49141
R416 VTAIL.n309 VTAIL.n294 2.71565
R417 VTAIL.n337 VTAIL.n280 2.71565
R418 VTAIL.n356 VTAIL.n355 2.71565
R419 VTAIL.n39 VTAIL.n24 2.71565
R420 VTAIL.n67 VTAIL.n10 2.71565
R421 VTAIL.n86 VTAIL.n85 2.71565
R422 VTAIL.n266 VTAIL.n265 2.71565
R423 VTAIL.n248 VTAIL.n191 2.71565
R424 VTAIL.n220 VTAIL.n205 2.71565
R425 VTAIL.n176 VTAIL.n175 2.71565
R426 VTAIL.n158 VTAIL.n101 2.71565
R427 VTAIL.n130 VTAIL.n115 2.71565
R428 VTAIL.n269 VTAIL.n179 2.10826
R429 VTAIL.n306 VTAIL.n305 1.93989
R430 VTAIL.n338 VTAIL.n278 1.93989
R431 VTAIL.n352 VTAIL.n272 1.93989
R432 VTAIL.n36 VTAIL.n35 1.93989
R433 VTAIL.n68 VTAIL.n8 1.93989
R434 VTAIL.n82 VTAIL.n2 1.93989
R435 VTAIL.n262 VTAIL.n182 1.93989
R436 VTAIL.n249 VTAIL.n189 1.93989
R437 VTAIL.n217 VTAIL.n216 1.93989
R438 VTAIL.n172 VTAIL.n92 1.93989
R439 VTAIL.n159 VTAIL.n99 1.93989
R440 VTAIL.n127 VTAIL.n126 1.93989
R441 VTAIL VTAIL.n89 1.34748
R442 VTAIL.n302 VTAIL.n296 1.16414
R443 VTAIL.n343 VTAIL.n341 1.16414
R444 VTAIL.n351 VTAIL.n274 1.16414
R445 VTAIL.n32 VTAIL.n26 1.16414
R446 VTAIL.n73 VTAIL.n71 1.16414
R447 VTAIL.n81 VTAIL.n4 1.16414
R448 VTAIL.n261 VTAIL.n184 1.16414
R449 VTAIL.n253 VTAIL.n252 1.16414
R450 VTAIL.n213 VTAIL.n207 1.16414
R451 VTAIL.n171 VTAIL.n94 1.16414
R452 VTAIL.n163 VTAIL.n162 1.16414
R453 VTAIL.n123 VTAIL.n117 1.16414
R454 VTAIL VTAIL.n359 0.761276
R455 VTAIL.n301 VTAIL.n298 0.388379
R456 VTAIL.n342 VTAIL.n276 0.388379
R457 VTAIL.n348 VTAIL.n347 0.388379
R458 VTAIL.n31 VTAIL.n28 0.388379
R459 VTAIL.n72 VTAIL.n6 0.388379
R460 VTAIL.n78 VTAIL.n77 0.388379
R461 VTAIL.n258 VTAIL.n257 0.388379
R462 VTAIL.n188 VTAIL.n186 0.388379
R463 VTAIL.n212 VTAIL.n209 0.388379
R464 VTAIL.n168 VTAIL.n167 0.388379
R465 VTAIL.n98 VTAIL.n96 0.388379
R466 VTAIL.n122 VTAIL.n119 0.388379
R467 VTAIL.n300 VTAIL.n295 0.155672
R468 VTAIL.n307 VTAIL.n295 0.155672
R469 VTAIL.n308 VTAIL.n307 0.155672
R470 VTAIL.n308 VTAIL.n291 0.155672
R471 VTAIL.n315 VTAIL.n291 0.155672
R472 VTAIL.n316 VTAIL.n315 0.155672
R473 VTAIL.n316 VTAIL.n287 0.155672
R474 VTAIL.n323 VTAIL.n287 0.155672
R475 VTAIL.n324 VTAIL.n323 0.155672
R476 VTAIL.n324 VTAIL.n283 0.155672
R477 VTAIL.n331 VTAIL.n283 0.155672
R478 VTAIL.n332 VTAIL.n331 0.155672
R479 VTAIL.n332 VTAIL.n279 0.155672
R480 VTAIL.n339 VTAIL.n279 0.155672
R481 VTAIL.n340 VTAIL.n339 0.155672
R482 VTAIL.n340 VTAIL.n275 0.155672
R483 VTAIL.n349 VTAIL.n275 0.155672
R484 VTAIL.n350 VTAIL.n349 0.155672
R485 VTAIL.n350 VTAIL.n271 0.155672
R486 VTAIL.n357 VTAIL.n271 0.155672
R487 VTAIL.n30 VTAIL.n25 0.155672
R488 VTAIL.n37 VTAIL.n25 0.155672
R489 VTAIL.n38 VTAIL.n37 0.155672
R490 VTAIL.n38 VTAIL.n21 0.155672
R491 VTAIL.n45 VTAIL.n21 0.155672
R492 VTAIL.n46 VTAIL.n45 0.155672
R493 VTAIL.n46 VTAIL.n17 0.155672
R494 VTAIL.n53 VTAIL.n17 0.155672
R495 VTAIL.n54 VTAIL.n53 0.155672
R496 VTAIL.n54 VTAIL.n13 0.155672
R497 VTAIL.n61 VTAIL.n13 0.155672
R498 VTAIL.n62 VTAIL.n61 0.155672
R499 VTAIL.n62 VTAIL.n9 0.155672
R500 VTAIL.n69 VTAIL.n9 0.155672
R501 VTAIL.n70 VTAIL.n69 0.155672
R502 VTAIL.n70 VTAIL.n5 0.155672
R503 VTAIL.n79 VTAIL.n5 0.155672
R504 VTAIL.n80 VTAIL.n79 0.155672
R505 VTAIL.n80 VTAIL.n1 0.155672
R506 VTAIL.n87 VTAIL.n1 0.155672
R507 VTAIL.n267 VTAIL.n181 0.155672
R508 VTAIL.n260 VTAIL.n181 0.155672
R509 VTAIL.n260 VTAIL.n259 0.155672
R510 VTAIL.n259 VTAIL.n185 0.155672
R511 VTAIL.n251 VTAIL.n185 0.155672
R512 VTAIL.n251 VTAIL.n250 0.155672
R513 VTAIL.n250 VTAIL.n190 0.155672
R514 VTAIL.n243 VTAIL.n190 0.155672
R515 VTAIL.n243 VTAIL.n242 0.155672
R516 VTAIL.n242 VTAIL.n194 0.155672
R517 VTAIL.n235 VTAIL.n194 0.155672
R518 VTAIL.n235 VTAIL.n234 0.155672
R519 VTAIL.n234 VTAIL.n198 0.155672
R520 VTAIL.n227 VTAIL.n198 0.155672
R521 VTAIL.n227 VTAIL.n226 0.155672
R522 VTAIL.n226 VTAIL.n202 0.155672
R523 VTAIL.n219 VTAIL.n202 0.155672
R524 VTAIL.n219 VTAIL.n218 0.155672
R525 VTAIL.n218 VTAIL.n206 0.155672
R526 VTAIL.n211 VTAIL.n206 0.155672
R527 VTAIL.n177 VTAIL.n91 0.155672
R528 VTAIL.n170 VTAIL.n91 0.155672
R529 VTAIL.n170 VTAIL.n169 0.155672
R530 VTAIL.n169 VTAIL.n95 0.155672
R531 VTAIL.n161 VTAIL.n95 0.155672
R532 VTAIL.n161 VTAIL.n160 0.155672
R533 VTAIL.n160 VTAIL.n100 0.155672
R534 VTAIL.n153 VTAIL.n100 0.155672
R535 VTAIL.n153 VTAIL.n152 0.155672
R536 VTAIL.n152 VTAIL.n104 0.155672
R537 VTAIL.n145 VTAIL.n104 0.155672
R538 VTAIL.n145 VTAIL.n144 0.155672
R539 VTAIL.n144 VTAIL.n108 0.155672
R540 VTAIL.n137 VTAIL.n108 0.155672
R541 VTAIL.n137 VTAIL.n136 0.155672
R542 VTAIL.n136 VTAIL.n112 0.155672
R543 VTAIL.n129 VTAIL.n112 0.155672
R544 VTAIL.n129 VTAIL.n128 0.155672
R545 VTAIL.n128 VTAIL.n116 0.155672
R546 VTAIL.n121 VTAIL.n116 0.155672
R547 VDD2.n173 VDD2.n89 289.615
R548 VDD2.n84 VDD2.n0 289.615
R549 VDD2.n174 VDD2.n173 185
R550 VDD2.n172 VDD2.n171 185
R551 VDD2.n93 VDD2.n92 185
R552 VDD2.n166 VDD2.n165 185
R553 VDD2.n164 VDD2.n95 185
R554 VDD2.n163 VDD2.n162 185
R555 VDD2.n98 VDD2.n96 185
R556 VDD2.n157 VDD2.n156 185
R557 VDD2.n155 VDD2.n154 185
R558 VDD2.n102 VDD2.n101 185
R559 VDD2.n149 VDD2.n148 185
R560 VDD2.n147 VDD2.n146 185
R561 VDD2.n106 VDD2.n105 185
R562 VDD2.n141 VDD2.n140 185
R563 VDD2.n139 VDD2.n138 185
R564 VDD2.n110 VDD2.n109 185
R565 VDD2.n133 VDD2.n132 185
R566 VDD2.n131 VDD2.n130 185
R567 VDD2.n114 VDD2.n113 185
R568 VDD2.n125 VDD2.n124 185
R569 VDD2.n123 VDD2.n122 185
R570 VDD2.n118 VDD2.n117 185
R571 VDD2.n28 VDD2.n27 185
R572 VDD2.n33 VDD2.n32 185
R573 VDD2.n35 VDD2.n34 185
R574 VDD2.n24 VDD2.n23 185
R575 VDD2.n41 VDD2.n40 185
R576 VDD2.n43 VDD2.n42 185
R577 VDD2.n20 VDD2.n19 185
R578 VDD2.n49 VDD2.n48 185
R579 VDD2.n51 VDD2.n50 185
R580 VDD2.n16 VDD2.n15 185
R581 VDD2.n57 VDD2.n56 185
R582 VDD2.n59 VDD2.n58 185
R583 VDD2.n12 VDD2.n11 185
R584 VDD2.n65 VDD2.n64 185
R585 VDD2.n67 VDD2.n66 185
R586 VDD2.n8 VDD2.n7 185
R587 VDD2.n74 VDD2.n73 185
R588 VDD2.n75 VDD2.n6 185
R589 VDD2.n77 VDD2.n76 185
R590 VDD2.n4 VDD2.n3 185
R591 VDD2.n83 VDD2.n82 185
R592 VDD2.n85 VDD2.n84 185
R593 VDD2.n119 VDD2.t0 147.659
R594 VDD2.n29 VDD2.t1 147.659
R595 VDD2.n173 VDD2.n172 104.615
R596 VDD2.n172 VDD2.n92 104.615
R597 VDD2.n165 VDD2.n92 104.615
R598 VDD2.n165 VDD2.n164 104.615
R599 VDD2.n164 VDD2.n163 104.615
R600 VDD2.n163 VDD2.n96 104.615
R601 VDD2.n156 VDD2.n96 104.615
R602 VDD2.n156 VDD2.n155 104.615
R603 VDD2.n155 VDD2.n101 104.615
R604 VDD2.n148 VDD2.n101 104.615
R605 VDD2.n148 VDD2.n147 104.615
R606 VDD2.n147 VDD2.n105 104.615
R607 VDD2.n140 VDD2.n105 104.615
R608 VDD2.n140 VDD2.n139 104.615
R609 VDD2.n139 VDD2.n109 104.615
R610 VDD2.n132 VDD2.n109 104.615
R611 VDD2.n132 VDD2.n131 104.615
R612 VDD2.n131 VDD2.n113 104.615
R613 VDD2.n124 VDD2.n113 104.615
R614 VDD2.n124 VDD2.n123 104.615
R615 VDD2.n123 VDD2.n117 104.615
R616 VDD2.n33 VDD2.n27 104.615
R617 VDD2.n34 VDD2.n33 104.615
R618 VDD2.n34 VDD2.n23 104.615
R619 VDD2.n41 VDD2.n23 104.615
R620 VDD2.n42 VDD2.n41 104.615
R621 VDD2.n42 VDD2.n19 104.615
R622 VDD2.n49 VDD2.n19 104.615
R623 VDD2.n50 VDD2.n49 104.615
R624 VDD2.n50 VDD2.n15 104.615
R625 VDD2.n57 VDD2.n15 104.615
R626 VDD2.n58 VDD2.n57 104.615
R627 VDD2.n58 VDD2.n11 104.615
R628 VDD2.n65 VDD2.n11 104.615
R629 VDD2.n66 VDD2.n65 104.615
R630 VDD2.n66 VDD2.n7 104.615
R631 VDD2.n74 VDD2.n7 104.615
R632 VDD2.n75 VDD2.n74 104.615
R633 VDD2.n76 VDD2.n75 104.615
R634 VDD2.n76 VDD2.n3 104.615
R635 VDD2.n83 VDD2.n3 104.615
R636 VDD2.n84 VDD2.n83 104.615
R637 VDD2.n178 VDD2.n88 97.3937
R638 VDD2.n178 VDD2.n177 53.1308
R639 VDD2.t0 VDD2.n117 52.3082
R640 VDD2.t1 VDD2.n27 52.3082
R641 VDD2.n119 VDD2.n118 15.6677
R642 VDD2.n29 VDD2.n28 15.6677
R643 VDD2.n166 VDD2.n95 13.1884
R644 VDD2.n77 VDD2.n6 13.1884
R645 VDD2.n167 VDD2.n93 12.8005
R646 VDD2.n162 VDD2.n97 12.8005
R647 VDD2.n122 VDD2.n121 12.8005
R648 VDD2.n32 VDD2.n31 12.8005
R649 VDD2.n73 VDD2.n72 12.8005
R650 VDD2.n78 VDD2.n4 12.8005
R651 VDD2.n171 VDD2.n170 12.0247
R652 VDD2.n161 VDD2.n98 12.0247
R653 VDD2.n125 VDD2.n116 12.0247
R654 VDD2.n35 VDD2.n26 12.0247
R655 VDD2.n71 VDD2.n8 12.0247
R656 VDD2.n82 VDD2.n81 12.0247
R657 VDD2.n174 VDD2.n91 11.249
R658 VDD2.n158 VDD2.n157 11.249
R659 VDD2.n126 VDD2.n114 11.249
R660 VDD2.n36 VDD2.n24 11.249
R661 VDD2.n68 VDD2.n67 11.249
R662 VDD2.n85 VDD2.n2 11.249
R663 VDD2.n175 VDD2.n89 10.4732
R664 VDD2.n154 VDD2.n100 10.4732
R665 VDD2.n130 VDD2.n129 10.4732
R666 VDD2.n40 VDD2.n39 10.4732
R667 VDD2.n64 VDD2.n10 10.4732
R668 VDD2.n86 VDD2.n0 10.4732
R669 VDD2.n153 VDD2.n102 9.69747
R670 VDD2.n133 VDD2.n112 9.69747
R671 VDD2.n43 VDD2.n22 9.69747
R672 VDD2.n63 VDD2.n12 9.69747
R673 VDD2.n177 VDD2.n176 9.45567
R674 VDD2.n88 VDD2.n87 9.45567
R675 VDD2.n145 VDD2.n144 9.3005
R676 VDD2.n104 VDD2.n103 9.3005
R677 VDD2.n151 VDD2.n150 9.3005
R678 VDD2.n153 VDD2.n152 9.3005
R679 VDD2.n100 VDD2.n99 9.3005
R680 VDD2.n159 VDD2.n158 9.3005
R681 VDD2.n161 VDD2.n160 9.3005
R682 VDD2.n97 VDD2.n94 9.3005
R683 VDD2.n176 VDD2.n175 9.3005
R684 VDD2.n91 VDD2.n90 9.3005
R685 VDD2.n170 VDD2.n169 9.3005
R686 VDD2.n168 VDD2.n167 9.3005
R687 VDD2.n143 VDD2.n142 9.3005
R688 VDD2.n108 VDD2.n107 9.3005
R689 VDD2.n137 VDD2.n136 9.3005
R690 VDD2.n135 VDD2.n134 9.3005
R691 VDD2.n112 VDD2.n111 9.3005
R692 VDD2.n129 VDD2.n128 9.3005
R693 VDD2.n127 VDD2.n126 9.3005
R694 VDD2.n116 VDD2.n115 9.3005
R695 VDD2.n121 VDD2.n120 9.3005
R696 VDD2.n87 VDD2.n86 9.3005
R697 VDD2.n2 VDD2.n1 9.3005
R698 VDD2.n81 VDD2.n80 9.3005
R699 VDD2.n79 VDD2.n78 9.3005
R700 VDD2.n18 VDD2.n17 9.3005
R701 VDD2.n47 VDD2.n46 9.3005
R702 VDD2.n45 VDD2.n44 9.3005
R703 VDD2.n22 VDD2.n21 9.3005
R704 VDD2.n39 VDD2.n38 9.3005
R705 VDD2.n37 VDD2.n36 9.3005
R706 VDD2.n26 VDD2.n25 9.3005
R707 VDD2.n31 VDD2.n30 9.3005
R708 VDD2.n53 VDD2.n52 9.3005
R709 VDD2.n55 VDD2.n54 9.3005
R710 VDD2.n14 VDD2.n13 9.3005
R711 VDD2.n61 VDD2.n60 9.3005
R712 VDD2.n63 VDD2.n62 9.3005
R713 VDD2.n10 VDD2.n9 9.3005
R714 VDD2.n69 VDD2.n68 9.3005
R715 VDD2.n71 VDD2.n70 9.3005
R716 VDD2.n72 VDD2.n5 9.3005
R717 VDD2.n150 VDD2.n149 8.92171
R718 VDD2.n134 VDD2.n110 8.92171
R719 VDD2.n44 VDD2.n20 8.92171
R720 VDD2.n60 VDD2.n59 8.92171
R721 VDD2.n146 VDD2.n104 8.14595
R722 VDD2.n138 VDD2.n137 8.14595
R723 VDD2.n48 VDD2.n47 8.14595
R724 VDD2.n56 VDD2.n14 8.14595
R725 VDD2.n145 VDD2.n106 7.3702
R726 VDD2.n141 VDD2.n108 7.3702
R727 VDD2.n51 VDD2.n18 7.3702
R728 VDD2.n55 VDD2.n16 7.3702
R729 VDD2.n142 VDD2.n106 6.59444
R730 VDD2.n142 VDD2.n141 6.59444
R731 VDD2.n52 VDD2.n51 6.59444
R732 VDD2.n52 VDD2.n16 6.59444
R733 VDD2.n146 VDD2.n145 5.81868
R734 VDD2.n138 VDD2.n108 5.81868
R735 VDD2.n48 VDD2.n18 5.81868
R736 VDD2.n56 VDD2.n55 5.81868
R737 VDD2.n149 VDD2.n104 5.04292
R738 VDD2.n137 VDD2.n110 5.04292
R739 VDD2.n47 VDD2.n20 5.04292
R740 VDD2.n59 VDD2.n14 5.04292
R741 VDD2.n120 VDD2.n119 4.38563
R742 VDD2.n30 VDD2.n29 4.38563
R743 VDD2.n150 VDD2.n102 4.26717
R744 VDD2.n134 VDD2.n133 4.26717
R745 VDD2.n44 VDD2.n43 4.26717
R746 VDD2.n60 VDD2.n12 4.26717
R747 VDD2.n177 VDD2.n89 3.49141
R748 VDD2.n154 VDD2.n153 3.49141
R749 VDD2.n130 VDD2.n112 3.49141
R750 VDD2.n40 VDD2.n22 3.49141
R751 VDD2.n64 VDD2.n63 3.49141
R752 VDD2.n88 VDD2.n0 3.49141
R753 VDD2.n175 VDD2.n174 2.71565
R754 VDD2.n157 VDD2.n100 2.71565
R755 VDD2.n129 VDD2.n114 2.71565
R756 VDD2.n39 VDD2.n24 2.71565
R757 VDD2.n67 VDD2.n10 2.71565
R758 VDD2.n86 VDD2.n85 2.71565
R759 VDD2.n171 VDD2.n91 1.93989
R760 VDD2.n158 VDD2.n98 1.93989
R761 VDD2.n126 VDD2.n125 1.93989
R762 VDD2.n36 VDD2.n35 1.93989
R763 VDD2.n68 VDD2.n8 1.93989
R764 VDD2.n82 VDD2.n2 1.93989
R765 VDD2.n170 VDD2.n93 1.16414
R766 VDD2.n162 VDD2.n161 1.16414
R767 VDD2.n122 VDD2.n116 1.16414
R768 VDD2.n32 VDD2.n26 1.16414
R769 VDD2.n73 VDD2.n71 1.16414
R770 VDD2.n81 VDD2.n4 1.16414
R771 VDD2 VDD2.n178 0.877655
R772 VDD2.n167 VDD2.n166 0.388379
R773 VDD2.n97 VDD2.n95 0.388379
R774 VDD2.n121 VDD2.n118 0.388379
R775 VDD2.n31 VDD2.n28 0.388379
R776 VDD2.n72 VDD2.n6 0.388379
R777 VDD2.n78 VDD2.n77 0.388379
R778 VDD2.n176 VDD2.n90 0.155672
R779 VDD2.n169 VDD2.n90 0.155672
R780 VDD2.n169 VDD2.n168 0.155672
R781 VDD2.n168 VDD2.n94 0.155672
R782 VDD2.n160 VDD2.n94 0.155672
R783 VDD2.n160 VDD2.n159 0.155672
R784 VDD2.n159 VDD2.n99 0.155672
R785 VDD2.n152 VDD2.n99 0.155672
R786 VDD2.n152 VDD2.n151 0.155672
R787 VDD2.n151 VDD2.n103 0.155672
R788 VDD2.n144 VDD2.n103 0.155672
R789 VDD2.n144 VDD2.n143 0.155672
R790 VDD2.n143 VDD2.n107 0.155672
R791 VDD2.n136 VDD2.n107 0.155672
R792 VDD2.n136 VDD2.n135 0.155672
R793 VDD2.n135 VDD2.n111 0.155672
R794 VDD2.n128 VDD2.n111 0.155672
R795 VDD2.n128 VDD2.n127 0.155672
R796 VDD2.n127 VDD2.n115 0.155672
R797 VDD2.n120 VDD2.n115 0.155672
R798 VDD2.n30 VDD2.n25 0.155672
R799 VDD2.n37 VDD2.n25 0.155672
R800 VDD2.n38 VDD2.n37 0.155672
R801 VDD2.n38 VDD2.n21 0.155672
R802 VDD2.n45 VDD2.n21 0.155672
R803 VDD2.n46 VDD2.n45 0.155672
R804 VDD2.n46 VDD2.n17 0.155672
R805 VDD2.n53 VDD2.n17 0.155672
R806 VDD2.n54 VDD2.n53 0.155672
R807 VDD2.n54 VDD2.n13 0.155672
R808 VDD2.n61 VDD2.n13 0.155672
R809 VDD2.n62 VDD2.n61 0.155672
R810 VDD2.n62 VDD2.n9 0.155672
R811 VDD2.n69 VDD2.n9 0.155672
R812 VDD2.n70 VDD2.n69 0.155672
R813 VDD2.n70 VDD2.n5 0.155672
R814 VDD2.n79 VDD2.n5 0.155672
R815 VDD2.n80 VDD2.n79 0.155672
R816 VDD2.n80 VDD2.n1 0.155672
R817 VDD2.n87 VDD2.n1 0.155672
R818 B.n614 B.n613 585
R819 B.n615 B.n123 585
R820 B.n617 B.n616 585
R821 B.n619 B.n122 585
R822 B.n622 B.n621 585
R823 B.n623 B.n121 585
R824 B.n625 B.n624 585
R825 B.n627 B.n120 585
R826 B.n630 B.n629 585
R827 B.n631 B.n119 585
R828 B.n633 B.n632 585
R829 B.n635 B.n118 585
R830 B.n638 B.n637 585
R831 B.n639 B.n117 585
R832 B.n641 B.n640 585
R833 B.n643 B.n116 585
R834 B.n646 B.n645 585
R835 B.n647 B.n115 585
R836 B.n649 B.n648 585
R837 B.n651 B.n114 585
R838 B.n654 B.n653 585
R839 B.n655 B.n113 585
R840 B.n657 B.n656 585
R841 B.n659 B.n112 585
R842 B.n662 B.n661 585
R843 B.n663 B.n111 585
R844 B.n665 B.n664 585
R845 B.n667 B.n110 585
R846 B.n670 B.n669 585
R847 B.n671 B.n109 585
R848 B.n673 B.n672 585
R849 B.n675 B.n108 585
R850 B.n678 B.n677 585
R851 B.n679 B.n107 585
R852 B.n681 B.n680 585
R853 B.n683 B.n106 585
R854 B.n686 B.n685 585
R855 B.n687 B.n105 585
R856 B.n689 B.n688 585
R857 B.n691 B.n104 585
R858 B.n694 B.n693 585
R859 B.n695 B.n103 585
R860 B.n697 B.n696 585
R861 B.n699 B.n102 585
R862 B.n702 B.n701 585
R863 B.n703 B.n101 585
R864 B.n705 B.n704 585
R865 B.n707 B.n100 585
R866 B.n710 B.n709 585
R867 B.n711 B.n99 585
R868 B.n713 B.n712 585
R869 B.n715 B.n98 585
R870 B.n717 B.n716 585
R871 B.n719 B.n718 585
R872 B.n722 B.n721 585
R873 B.n723 B.n93 585
R874 B.n725 B.n724 585
R875 B.n727 B.n92 585
R876 B.n730 B.n729 585
R877 B.n731 B.n91 585
R878 B.n733 B.n732 585
R879 B.n735 B.n90 585
R880 B.n737 B.n736 585
R881 B.n739 B.n738 585
R882 B.n742 B.n741 585
R883 B.n743 B.n85 585
R884 B.n745 B.n744 585
R885 B.n747 B.n84 585
R886 B.n750 B.n749 585
R887 B.n751 B.n83 585
R888 B.n753 B.n752 585
R889 B.n755 B.n82 585
R890 B.n758 B.n757 585
R891 B.n759 B.n81 585
R892 B.n761 B.n760 585
R893 B.n763 B.n80 585
R894 B.n766 B.n765 585
R895 B.n767 B.n79 585
R896 B.n769 B.n768 585
R897 B.n771 B.n78 585
R898 B.n774 B.n773 585
R899 B.n775 B.n77 585
R900 B.n777 B.n776 585
R901 B.n779 B.n76 585
R902 B.n782 B.n781 585
R903 B.n783 B.n75 585
R904 B.n785 B.n784 585
R905 B.n787 B.n74 585
R906 B.n790 B.n789 585
R907 B.n791 B.n73 585
R908 B.n793 B.n792 585
R909 B.n795 B.n72 585
R910 B.n798 B.n797 585
R911 B.n799 B.n71 585
R912 B.n801 B.n800 585
R913 B.n803 B.n70 585
R914 B.n806 B.n805 585
R915 B.n807 B.n69 585
R916 B.n809 B.n808 585
R917 B.n811 B.n68 585
R918 B.n814 B.n813 585
R919 B.n815 B.n67 585
R920 B.n817 B.n816 585
R921 B.n819 B.n66 585
R922 B.n822 B.n821 585
R923 B.n823 B.n65 585
R924 B.n825 B.n824 585
R925 B.n827 B.n64 585
R926 B.n830 B.n829 585
R927 B.n831 B.n63 585
R928 B.n833 B.n832 585
R929 B.n835 B.n62 585
R930 B.n838 B.n837 585
R931 B.n839 B.n61 585
R932 B.n841 B.n840 585
R933 B.n843 B.n60 585
R934 B.n846 B.n845 585
R935 B.n847 B.n59 585
R936 B.n611 B.n57 585
R937 B.n850 B.n57 585
R938 B.n610 B.n56 585
R939 B.n851 B.n56 585
R940 B.n609 B.n55 585
R941 B.n852 B.n55 585
R942 B.n608 B.n607 585
R943 B.n607 B.n51 585
R944 B.n606 B.n50 585
R945 B.n858 B.n50 585
R946 B.n605 B.n49 585
R947 B.n859 B.n49 585
R948 B.n604 B.n48 585
R949 B.n860 B.n48 585
R950 B.n603 B.n602 585
R951 B.n602 B.n44 585
R952 B.n601 B.n43 585
R953 B.n866 B.n43 585
R954 B.n600 B.n42 585
R955 B.n867 B.n42 585
R956 B.n599 B.n41 585
R957 B.n868 B.n41 585
R958 B.n598 B.n597 585
R959 B.n597 B.n37 585
R960 B.n596 B.n36 585
R961 B.n874 B.n36 585
R962 B.n595 B.n35 585
R963 B.n875 B.n35 585
R964 B.n594 B.n34 585
R965 B.n876 B.n34 585
R966 B.n593 B.n592 585
R967 B.n592 B.n30 585
R968 B.n591 B.n29 585
R969 B.n882 B.n29 585
R970 B.n590 B.n28 585
R971 B.n883 B.n28 585
R972 B.n589 B.n27 585
R973 B.n884 B.n27 585
R974 B.n588 B.n587 585
R975 B.n587 B.n23 585
R976 B.n586 B.n22 585
R977 B.n890 B.n22 585
R978 B.n585 B.n21 585
R979 B.n891 B.n21 585
R980 B.n584 B.n20 585
R981 B.n892 B.n20 585
R982 B.n583 B.n582 585
R983 B.n582 B.n19 585
R984 B.n581 B.n15 585
R985 B.n898 B.n15 585
R986 B.n580 B.n14 585
R987 B.n899 B.n14 585
R988 B.n579 B.n13 585
R989 B.n900 B.n13 585
R990 B.n578 B.n577 585
R991 B.n577 B.n12 585
R992 B.n576 B.n575 585
R993 B.n576 B.n8 585
R994 B.n574 B.n7 585
R995 B.n907 B.n7 585
R996 B.n573 B.n6 585
R997 B.n908 B.n6 585
R998 B.n572 B.n5 585
R999 B.n909 B.n5 585
R1000 B.n571 B.n570 585
R1001 B.n570 B.n4 585
R1002 B.n569 B.n124 585
R1003 B.n569 B.n568 585
R1004 B.n559 B.n125 585
R1005 B.n126 B.n125 585
R1006 B.n561 B.n560 585
R1007 B.n562 B.n561 585
R1008 B.n558 B.n131 585
R1009 B.n131 B.n130 585
R1010 B.n557 B.n556 585
R1011 B.n556 B.n555 585
R1012 B.n133 B.n132 585
R1013 B.n548 B.n133 585
R1014 B.n547 B.n546 585
R1015 B.n549 B.n547 585
R1016 B.n545 B.n138 585
R1017 B.n138 B.n137 585
R1018 B.n544 B.n543 585
R1019 B.n543 B.n542 585
R1020 B.n140 B.n139 585
R1021 B.n141 B.n140 585
R1022 B.n535 B.n534 585
R1023 B.n536 B.n535 585
R1024 B.n533 B.n146 585
R1025 B.n146 B.n145 585
R1026 B.n532 B.n531 585
R1027 B.n531 B.n530 585
R1028 B.n148 B.n147 585
R1029 B.n149 B.n148 585
R1030 B.n523 B.n522 585
R1031 B.n524 B.n523 585
R1032 B.n521 B.n154 585
R1033 B.n154 B.n153 585
R1034 B.n520 B.n519 585
R1035 B.n519 B.n518 585
R1036 B.n156 B.n155 585
R1037 B.n157 B.n156 585
R1038 B.n511 B.n510 585
R1039 B.n512 B.n511 585
R1040 B.n509 B.n162 585
R1041 B.n162 B.n161 585
R1042 B.n508 B.n507 585
R1043 B.n507 B.n506 585
R1044 B.n164 B.n163 585
R1045 B.n165 B.n164 585
R1046 B.n499 B.n498 585
R1047 B.n500 B.n499 585
R1048 B.n497 B.n170 585
R1049 B.n170 B.n169 585
R1050 B.n496 B.n495 585
R1051 B.n495 B.n494 585
R1052 B.n172 B.n171 585
R1053 B.n173 B.n172 585
R1054 B.n487 B.n486 585
R1055 B.n488 B.n487 585
R1056 B.n485 B.n178 585
R1057 B.n178 B.n177 585
R1058 B.n484 B.n483 585
R1059 B.n483 B.n482 585
R1060 B.n479 B.n182 585
R1061 B.n478 B.n477 585
R1062 B.n475 B.n183 585
R1063 B.n475 B.n181 585
R1064 B.n474 B.n473 585
R1065 B.n472 B.n471 585
R1066 B.n470 B.n185 585
R1067 B.n468 B.n467 585
R1068 B.n466 B.n186 585
R1069 B.n465 B.n464 585
R1070 B.n462 B.n187 585
R1071 B.n460 B.n459 585
R1072 B.n458 B.n188 585
R1073 B.n457 B.n456 585
R1074 B.n454 B.n189 585
R1075 B.n452 B.n451 585
R1076 B.n450 B.n190 585
R1077 B.n449 B.n448 585
R1078 B.n446 B.n191 585
R1079 B.n444 B.n443 585
R1080 B.n442 B.n192 585
R1081 B.n441 B.n440 585
R1082 B.n438 B.n193 585
R1083 B.n436 B.n435 585
R1084 B.n434 B.n194 585
R1085 B.n433 B.n432 585
R1086 B.n430 B.n195 585
R1087 B.n428 B.n427 585
R1088 B.n426 B.n196 585
R1089 B.n425 B.n424 585
R1090 B.n422 B.n197 585
R1091 B.n420 B.n419 585
R1092 B.n418 B.n198 585
R1093 B.n417 B.n416 585
R1094 B.n414 B.n199 585
R1095 B.n412 B.n411 585
R1096 B.n410 B.n200 585
R1097 B.n409 B.n408 585
R1098 B.n406 B.n201 585
R1099 B.n404 B.n403 585
R1100 B.n402 B.n202 585
R1101 B.n401 B.n400 585
R1102 B.n398 B.n203 585
R1103 B.n396 B.n395 585
R1104 B.n394 B.n204 585
R1105 B.n393 B.n392 585
R1106 B.n390 B.n205 585
R1107 B.n388 B.n387 585
R1108 B.n386 B.n206 585
R1109 B.n385 B.n384 585
R1110 B.n382 B.n207 585
R1111 B.n380 B.n379 585
R1112 B.n378 B.n208 585
R1113 B.n377 B.n376 585
R1114 B.n374 B.n209 585
R1115 B.n372 B.n371 585
R1116 B.n370 B.n210 585
R1117 B.n369 B.n368 585
R1118 B.n366 B.n214 585
R1119 B.n364 B.n363 585
R1120 B.n362 B.n215 585
R1121 B.n361 B.n360 585
R1122 B.n358 B.n216 585
R1123 B.n356 B.n355 585
R1124 B.n354 B.n217 585
R1125 B.n352 B.n351 585
R1126 B.n349 B.n220 585
R1127 B.n347 B.n346 585
R1128 B.n345 B.n221 585
R1129 B.n344 B.n343 585
R1130 B.n341 B.n222 585
R1131 B.n339 B.n338 585
R1132 B.n337 B.n223 585
R1133 B.n336 B.n335 585
R1134 B.n333 B.n224 585
R1135 B.n331 B.n330 585
R1136 B.n329 B.n225 585
R1137 B.n328 B.n327 585
R1138 B.n325 B.n226 585
R1139 B.n323 B.n322 585
R1140 B.n321 B.n227 585
R1141 B.n320 B.n319 585
R1142 B.n317 B.n228 585
R1143 B.n315 B.n314 585
R1144 B.n313 B.n229 585
R1145 B.n312 B.n311 585
R1146 B.n309 B.n230 585
R1147 B.n307 B.n306 585
R1148 B.n305 B.n231 585
R1149 B.n304 B.n303 585
R1150 B.n301 B.n232 585
R1151 B.n299 B.n298 585
R1152 B.n297 B.n233 585
R1153 B.n296 B.n295 585
R1154 B.n293 B.n234 585
R1155 B.n291 B.n290 585
R1156 B.n289 B.n235 585
R1157 B.n288 B.n287 585
R1158 B.n285 B.n236 585
R1159 B.n283 B.n282 585
R1160 B.n281 B.n237 585
R1161 B.n280 B.n279 585
R1162 B.n277 B.n238 585
R1163 B.n275 B.n274 585
R1164 B.n273 B.n239 585
R1165 B.n272 B.n271 585
R1166 B.n269 B.n240 585
R1167 B.n267 B.n266 585
R1168 B.n265 B.n241 585
R1169 B.n264 B.n263 585
R1170 B.n261 B.n242 585
R1171 B.n259 B.n258 585
R1172 B.n257 B.n243 585
R1173 B.n256 B.n255 585
R1174 B.n253 B.n244 585
R1175 B.n251 B.n250 585
R1176 B.n249 B.n245 585
R1177 B.n248 B.n247 585
R1178 B.n180 B.n179 585
R1179 B.n181 B.n180 585
R1180 B.n481 B.n480 585
R1181 B.n482 B.n481 585
R1182 B.n176 B.n175 585
R1183 B.n177 B.n176 585
R1184 B.n490 B.n489 585
R1185 B.n489 B.n488 585
R1186 B.n491 B.n174 585
R1187 B.n174 B.n173 585
R1188 B.n493 B.n492 585
R1189 B.n494 B.n493 585
R1190 B.n168 B.n167 585
R1191 B.n169 B.n168 585
R1192 B.n502 B.n501 585
R1193 B.n501 B.n500 585
R1194 B.n503 B.n166 585
R1195 B.n166 B.n165 585
R1196 B.n505 B.n504 585
R1197 B.n506 B.n505 585
R1198 B.n160 B.n159 585
R1199 B.n161 B.n160 585
R1200 B.n514 B.n513 585
R1201 B.n513 B.n512 585
R1202 B.n515 B.n158 585
R1203 B.n158 B.n157 585
R1204 B.n517 B.n516 585
R1205 B.n518 B.n517 585
R1206 B.n152 B.n151 585
R1207 B.n153 B.n152 585
R1208 B.n526 B.n525 585
R1209 B.n525 B.n524 585
R1210 B.n527 B.n150 585
R1211 B.n150 B.n149 585
R1212 B.n529 B.n528 585
R1213 B.n530 B.n529 585
R1214 B.n144 B.n143 585
R1215 B.n145 B.n144 585
R1216 B.n538 B.n537 585
R1217 B.n537 B.n536 585
R1218 B.n539 B.n142 585
R1219 B.n142 B.n141 585
R1220 B.n541 B.n540 585
R1221 B.n542 B.n541 585
R1222 B.n136 B.n135 585
R1223 B.n137 B.n136 585
R1224 B.n551 B.n550 585
R1225 B.n550 B.n549 585
R1226 B.n552 B.n134 585
R1227 B.n548 B.n134 585
R1228 B.n554 B.n553 585
R1229 B.n555 B.n554 585
R1230 B.n129 B.n128 585
R1231 B.n130 B.n129 585
R1232 B.n564 B.n563 585
R1233 B.n563 B.n562 585
R1234 B.n565 B.n127 585
R1235 B.n127 B.n126 585
R1236 B.n567 B.n566 585
R1237 B.n568 B.n567 585
R1238 B.n3 B.n0 585
R1239 B.n4 B.n3 585
R1240 B.n906 B.n1 585
R1241 B.n907 B.n906 585
R1242 B.n905 B.n904 585
R1243 B.n905 B.n8 585
R1244 B.n903 B.n9 585
R1245 B.n12 B.n9 585
R1246 B.n902 B.n901 585
R1247 B.n901 B.n900 585
R1248 B.n11 B.n10 585
R1249 B.n899 B.n11 585
R1250 B.n897 B.n896 585
R1251 B.n898 B.n897 585
R1252 B.n895 B.n16 585
R1253 B.n19 B.n16 585
R1254 B.n894 B.n893 585
R1255 B.n893 B.n892 585
R1256 B.n18 B.n17 585
R1257 B.n891 B.n18 585
R1258 B.n889 B.n888 585
R1259 B.n890 B.n889 585
R1260 B.n887 B.n24 585
R1261 B.n24 B.n23 585
R1262 B.n886 B.n885 585
R1263 B.n885 B.n884 585
R1264 B.n26 B.n25 585
R1265 B.n883 B.n26 585
R1266 B.n881 B.n880 585
R1267 B.n882 B.n881 585
R1268 B.n879 B.n31 585
R1269 B.n31 B.n30 585
R1270 B.n878 B.n877 585
R1271 B.n877 B.n876 585
R1272 B.n33 B.n32 585
R1273 B.n875 B.n33 585
R1274 B.n873 B.n872 585
R1275 B.n874 B.n873 585
R1276 B.n871 B.n38 585
R1277 B.n38 B.n37 585
R1278 B.n870 B.n869 585
R1279 B.n869 B.n868 585
R1280 B.n40 B.n39 585
R1281 B.n867 B.n40 585
R1282 B.n865 B.n864 585
R1283 B.n866 B.n865 585
R1284 B.n863 B.n45 585
R1285 B.n45 B.n44 585
R1286 B.n862 B.n861 585
R1287 B.n861 B.n860 585
R1288 B.n47 B.n46 585
R1289 B.n859 B.n47 585
R1290 B.n857 B.n856 585
R1291 B.n858 B.n857 585
R1292 B.n855 B.n52 585
R1293 B.n52 B.n51 585
R1294 B.n854 B.n853 585
R1295 B.n853 B.n852 585
R1296 B.n54 B.n53 585
R1297 B.n851 B.n54 585
R1298 B.n849 B.n848 585
R1299 B.n850 B.n849 585
R1300 B.n910 B.n909 585
R1301 B.n908 B.n2 585
R1302 B.n849 B.n59 502.111
R1303 B.n613 B.n57 502.111
R1304 B.n483 B.n180 502.111
R1305 B.n481 B.n182 502.111
R1306 B.n94 B.t14 430.247
R1307 B.n218 B.t12 430.247
R1308 B.n86 B.t8 430.247
R1309 B.n211 B.t5 430.247
R1310 B.n95 B.t15 356.55
R1311 B.n219 B.t11 356.55
R1312 B.n87 B.t9 356.55
R1313 B.n212 B.t4 356.55
R1314 B.n86 B.t6 322.274
R1315 B.n94 B.t13 322.274
R1316 B.n218 B.t10 322.274
R1317 B.n211 B.t2 322.274
R1318 B.n612 B.n58 256.663
R1319 B.n618 B.n58 256.663
R1320 B.n620 B.n58 256.663
R1321 B.n626 B.n58 256.663
R1322 B.n628 B.n58 256.663
R1323 B.n634 B.n58 256.663
R1324 B.n636 B.n58 256.663
R1325 B.n642 B.n58 256.663
R1326 B.n644 B.n58 256.663
R1327 B.n650 B.n58 256.663
R1328 B.n652 B.n58 256.663
R1329 B.n658 B.n58 256.663
R1330 B.n660 B.n58 256.663
R1331 B.n666 B.n58 256.663
R1332 B.n668 B.n58 256.663
R1333 B.n674 B.n58 256.663
R1334 B.n676 B.n58 256.663
R1335 B.n682 B.n58 256.663
R1336 B.n684 B.n58 256.663
R1337 B.n690 B.n58 256.663
R1338 B.n692 B.n58 256.663
R1339 B.n698 B.n58 256.663
R1340 B.n700 B.n58 256.663
R1341 B.n706 B.n58 256.663
R1342 B.n708 B.n58 256.663
R1343 B.n714 B.n58 256.663
R1344 B.n97 B.n58 256.663
R1345 B.n720 B.n58 256.663
R1346 B.n726 B.n58 256.663
R1347 B.n728 B.n58 256.663
R1348 B.n734 B.n58 256.663
R1349 B.n89 B.n58 256.663
R1350 B.n740 B.n58 256.663
R1351 B.n746 B.n58 256.663
R1352 B.n748 B.n58 256.663
R1353 B.n754 B.n58 256.663
R1354 B.n756 B.n58 256.663
R1355 B.n762 B.n58 256.663
R1356 B.n764 B.n58 256.663
R1357 B.n770 B.n58 256.663
R1358 B.n772 B.n58 256.663
R1359 B.n778 B.n58 256.663
R1360 B.n780 B.n58 256.663
R1361 B.n786 B.n58 256.663
R1362 B.n788 B.n58 256.663
R1363 B.n794 B.n58 256.663
R1364 B.n796 B.n58 256.663
R1365 B.n802 B.n58 256.663
R1366 B.n804 B.n58 256.663
R1367 B.n810 B.n58 256.663
R1368 B.n812 B.n58 256.663
R1369 B.n818 B.n58 256.663
R1370 B.n820 B.n58 256.663
R1371 B.n826 B.n58 256.663
R1372 B.n828 B.n58 256.663
R1373 B.n834 B.n58 256.663
R1374 B.n836 B.n58 256.663
R1375 B.n842 B.n58 256.663
R1376 B.n844 B.n58 256.663
R1377 B.n476 B.n181 256.663
R1378 B.n184 B.n181 256.663
R1379 B.n469 B.n181 256.663
R1380 B.n463 B.n181 256.663
R1381 B.n461 B.n181 256.663
R1382 B.n455 B.n181 256.663
R1383 B.n453 B.n181 256.663
R1384 B.n447 B.n181 256.663
R1385 B.n445 B.n181 256.663
R1386 B.n439 B.n181 256.663
R1387 B.n437 B.n181 256.663
R1388 B.n431 B.n181 256.663
R1389 B.n429 B.n181 256.663
R1390 B.n423 B.n181 256.663
R1391 B.n421 B.n181 256.663
R1392 B.n415 B.n181 256.663
R1393 B.n413 B.n181 256.663
R1394 B.n407 B.n181 256.663
R1395 B.n405 B.n181 256.663
R1396 B.n399 B.n181 256.663
R1397 B.n397 B.n181 256.663
R1398 B.n391 B.n181 256.663
R1399 B.n389 B.n181 256.663
R1400 B.n383 B.n181 256.663
R1401 B.n381 B.n181 256.663
R1402 B.n375 B.n181 256.663
R1403 B.n373 B.n181 256.663
R1404 B.n367 B.n181 256.663
R1405 B.n365 B.n181 256.663
R1406 B.n359 B.n181 256.663
R1407 B.n357 B.n181 256.663
R1408 B.n350 B.n181 256.663
R1409 B.n348 B.n181 256.663
R1410 B.n342 B.n181 256.663
R1411 B.n340 B.n181 256.663
R1412 B.n334 B.n181 256.663
R1413 B.n332 B.n181 256.663
R1414 B.n326 B.n181 256.663
R1415 B.n324 B.n181 256.663
R1416 B.n318 B.n181 256.663
R1417 B.n316 B.n181 256.663
R1418 B.n310 B.n181 256.663
R1419 B.n308 B.n181 256.663
R1420 B.n302 B.n181 256.663
R1421 B.n300 B.n181 256.663
R1422 B.n294 B.n181 256.663
R1423 B.n292 B.n181 256.663
R1424 B.n286 B.n181 256.663
R1425 B.n284 B.n181 256.663
R1426 B.n278 B.n181 256.663
R1427 B.n276 B.n181 256.663
R1428 B.n270 B.n181 256.663
R1429 B.n268 B.n181 256.663
R1430 B.n262 B.n181 256.663
R1431 B.n260 B.n181 256.663
R1432 B.n254 B.n181 256.663
R1433 B.n252 B.n181 256.663
R1434 B.n246 B.n181 256.663
R1435 B.n912 B.n911 256.663
R1436 B.n845 B.n843 163.367
R1437 B.n841 B.n61 163.367
R1438 B.n837 B.n835 163.367
R1439 B.n833 B.n63 163.367
R1440 B.n829 B.n827 163.367
R1441 B.n825 B.n65 163.367
R1442 B.n821 B.n819 163.367
R1443 B.n817 B.n67 163.367
R1444 B.n813 B.n811 163.367
R1445 B.n809 B.n69 163.367
R1446 B.n805 B.n803 163.367
R1447 B.n801 B.n71 163.367
R1448 B.n797 B.n795 163.367
R1449 B.n793 B.n73 163.367
R1450 B.n789 B.n787 163.367
R1451 B.n785 B.n75 163.367
R1452 B.n781 B.n779 163.367
R1453 B.n777 B.n77 163.367
R1454 B.n773 B.n771 163.367
R1455 B.n769 B.n79 163.367
R1456 B.n765 B.n763 163.367
R1457 B.n761 B.n81 163.367
R1458 B.n757 B.n755 163.367
R1459 B.n753 B.n83 163.367
R1460 B.n749 B.n747 163.367
R1461 B.n745 B.n85 163.367
R1462 B.n741 B.n739 163.367
R1463 B.n736 B.n735 163.367
R1464 B.n733 B.n91 163.367
R1465 B.n729 B.n727 163.367
R1466 B.n725 B.n93 163.367
R1467 B.n721 B.n719 163.367
R1468 B.n716 B.n715 163.367
R1469 B.n713 B.n99 163.367
R1470 B.n709 B.n707 163.367
R1471 B.n705 B.n101 163.367
R1472 B.n701 B.n699 163.367
R1473 B.n697 B.n103 163.367
R1474 B.n693 B.n691 163.367
R1475 B.n689 B.n105 163.367
R1476 B.n685 B.n683 163.367
R1477 B.n681 B.n107 163.367
R1478 B.n677 B.n675 163.367
R1479 B.n673 B.n109 163.367
R1480 B.n669 B.n667 163.367
R1481 B.n665 B.n111 163.367
R1482 B.n661 B.n659 163.367
R1483 B.n657 B.n113 163.367
R1484 B.n653 B.n651 163.367
R1485 B.n649 B.n115 163.367
R1486 B.n645 B.n643 163.367
R1487 B.n641 B.n117 163.367
R1488 B.n637 B.n635 163.367
R1489 B.n633 B.n119 163.367
R1490 B.n629 B.n627 163.367
R1491 B.n625 B.n121 163.367
R1492 B.n621 B.n619 163.367
R1493 B.n617 B.n123 163.367
R1494 B.n483 B.n178 163.367
R1495 B.n487 B.n178 163.367
R1496 B.n487 B.n172 163.367
R1497 B.n495 B.n172 163.367
R1498 B.n495 B.n170 163.367
R1499 B.n499 B.n170 163.367
R1500 B.n499 B.n164 163.367
R1501 B.n507 B.n164 163.367
R1502 B.n507 B.n162 163.367
R1503 B.n511 B.n162 163.367
R1504 B.n511 B.n156 163.367
R1505 B.n519 B.n156 163.367
R1506 B.n519 B.n154 163.367
R1507 B.n523 B.n154 163.367
R1508 B.n523 B.n148 163.367
R1509 B.n531 B.n148 163.367
R1510 B.n531 B.n146 163.367
R1511 B.n535 B.n146 163.367
R1512 B.n535 B.n140 163.367
R1513 B.n543 B.n140 163.367
R1514 B.n543 B.n138 163.367
R1515 B.n547 B.n138 163.367
R1516 B.n547 B.n133 163.367
R1517 B.n556 B.n133 163.367
R1518 B.n556 B.n131 163.367
R1519 B.n561 B.n131 163.367
R1520 B.n561 B.n125 163.367
R1521 B.n569 B.n125 163.367
R1522 B.n570 B.n569 163.367
R1523 B.n570 B.n5 163.367
R1524 B.n6 B.n5 163.367
R1525 B.n7 B.n6 163.367
R1526 B.n576 B.n7 163.367
R1527 B.n577 B.n576 163.367
R1528 B.n577 B.n13 163.367
R1529 B.n14 B.n13 163.367
R1530 B.n15 B.n14 163.367
R1531 B.n582 B.n15 163.367
R1532 B.n582 B.n20 163.367
R1533 B.n21 B.n20 163.367
R1534 B.n22 B.n21 163.367
R1535 B.n587 B.n22 163.367
R1536 B.n587 B.n27 163.367
R1537 B.n28 B.n27 163.367
R1538 B.n29 B.n28 163.367
R1539 B.n592 B.n29 163.367
R1540 B.n592 B.n34 163.367
R1541 B.n35 B.n34 163.367
R1542 B.n36 B.n35 163.367
R1543 B.n597 B.n36 163.367
R1544 B.n597 B.n41 163.367
R1545 B.n42 B.n41 163.367
R1546 B.n43 B.n42 163.367
R1547 B.n602 B.n43 163.367
R1548 B.n602 B.n48 163.367
R1549 B.n49 B.n48 163.367
R1550 B.n50 B.n49 163.367
R1551 B.n607 B.n50 163.367
R1552 B.n607 B.n55 163.367
R1553 B.n56 B.n55 163.367
R1554 B.n57 B.n56 163.367
R1555 B.n477 B.n475 163.367
R1556 B.n475 B.n474 163.367
R1557 B.n471 B.n470 163.367
R1558 B.n468 B.n186 163.367
R1559 B.n464 B.n462 163.367
R1560 B.n460 B.n188 163.367
R1561 B.n456 B.n454 163.367
R1562 B.n452 B.n190 163.367
R1563 B.n448 B.n446 163.367
R1564 B.n444 B.n192 163.367
R1565 B.n440 B.n438 163.367
R1566 B.n436 B.n194 163.367
R1567 B.n432 B.n430 163.367
R1568 B.n428 B.n196 163.367
R1569 B.n424 B.n422 163.367
R1570 B.n420 B.n198 163.367
R1571 B.n416 B.n414 163.367
R1572 B.n412 B.n200 163.367
R1573 B.n408 B.n406 163.367
R1574 B.n404 B.n202 163.367
R1575 B.n400 B.n398 163.367
R1576 B.n396 B.n204 163.367
R1577 B.n392 B.n390 163.367
R1578 B.n388 B.n206 163.367
R1579 B.n384 B.n382 163.367
R1580 B.n380 B.n208 163.367
R1581 B.n376 B.n374 163.367
R1582 B.n372 B.n210 163.367
R1583 B.n368 B.n366 163.367
R1584 B.n364 B.n215 163.367
R1585 B.n360 B.n358 163.367
R1586 B.n356 B.n217 163.367
R1587 B.n351 B.n349 163.367
R1588 B.n347 B.n221 163.367
R1589 B.n343 B.n341 163.367
R1590 B.n339 B.n223 163.367
R1591 B.n335 B.n333 163.367
R1592 B.n331 B.n225 163.367
R1593 B.n327 B.n325 163.367
R1594 B.n323 B.n227 163.367
R1595 B.n319 B.n317 163.367
R1596 B.n315 B.n229 163.367
R1597 B.n311 B.n309 163.367
R1598 B.n307 B.n231 163.367
R1599 B.n303 B.n301 163.367
R1600 B.n299 B.n233 163.367
R1601 B.n295 B.n293 163.367
R1602 B.n291 B.n235 163.367
R1603 B.n287 B.n285 163.367
R1604 B.n283 B.n237 163.367
R1605 B.n279 B.n277 163.367
R1606 B.n275 B.n239 163.367
R1607 B.n271 B.n269 163.367
R1608 B.n267 B.n241 163.367
R1609 B.n263 B.n261 163.367
R1610 B.n259 B.n243 163.367
R1611 B.n255 B.n253 163.367
R1612 B.n251 B.n245 163.367
R1613 B.n247 B.n180 163.367
R1614 B.n481 B.n176 163.367
R1615 B.n489 B.n176 163.367
R1616 B.n489 B.n174 163.367
R1617 B.n493 B.n174 163.367
R1618 B.n493 B.n168 163.367
R1619 B.n501 B.n168 163.367
R1620 B.n501 B.n166 163.367
R1621 B.n505 B.n166 163.367
R1622 B.n505 B.n160 163.367
R1623 B.n513 B.n160 163.367
R1624 B.n513 B.n158 163.367
R1625 B.n517 B.n158 163.367
R1626 B.n517 B.n152 163.367
R1627 B.n525 B.n152 163.367
R1628 B.n525 B.n150 163.367
R1629 B.n529 B.n150 163.367
R1630 B.n529 B.n144 163.367
R1631 B.n537 B.n144 163.367
R1632 B.n537 B.n142 163.367
R1633 B.n541 B.n142 163.367
R1634 B.n541 B.n136 163.367
R1635 B.n550 B.n136 163.367
R1636 B.n550 B.n134 163.367
R1637 B.n554 B.n134 163.367
R1638 B.n554 B.n129 163.367
R1639 B.n563 B.n129 163.367
R1640 B.n563 B.n127 163.367
R1641 B.n567 B.n127 163.367
R1642 B.n567 B.n3 163.367
R1643 B.n910 B.n3 163.367
R1644 B.n906 B.n2 163.367
R1645 B.n906 B.n905 163.367
R1646 B.n905 B.n9 163.367
R1647 B.n901 B.n9 163.367
R1648 B.n901 B.n11 163.367
R1649 B.n897 B.n11 163.367
R1650 B.n897 B.n16 163.367
R1651 B.n893 B.n16 163.367
R1652 B.n893 B.n18 163.367
R1653 B.n889 B.n18 163.367
R1654 B.n889 B.n24 163.367
R1655 B.n885 B.n24 163.367
R1656 B.n885 B.n26 163.367
R1657 B.n881 B.n26 163.367
R1658 B.n881 B.n31 163.367
R1659 B.n877 B.n31 163.367
R1660 B.n877 B.n33 163.367
R1661 B.n873 B.n33 163.367
R1662 B.n873 B.n38 163.367
R1663 B.n869 B.n38 163.367
R1664 B.n869 B.n40 163.367
R1665 B.n865 B.n40 163.367
R1666 B.n865 B.n45 163.367
R1667 B.n861 B.n45 163.367
R1668 B.n861 B.n47 163.367
R1669 B.n857 B.n47 163.367
R1670 B.n857 B.n52 163.367
R1671 B.n853 B.n52 163.367
R1672 B.n853 B.n54 163.367
R1673 B.n849 B.n54 163.367
R1674 B.n87 B.n86 73.6975
R1675 B.n95 B.n94 73.6975
R1676 B.n219 B.n218 73.6975
R1677 B.n212 B.n211 73.6975
R1678 B.n844 B.n59 71.676
R1679 B.n843 B.n842 71.676
R1680 B.n836 B.n61 71.676
R1681 B.n835 B.n834 71.676
R1682 B.n828 B.n63 71.676
R1683 B.n827 B.n826 71.676
R1684 B.n820 B.n65 71.676
R1685 B.n819 B.n818 71.676
R1686 B.n812 B.n67 71.676
R1687 B.n811 B.n810 71.676
R1688 B.n804 B.n69 71.676
R1689 B.n803 B.n802 71.676
R1690 B.n796 B.n71 71.676
R1691 B.n795 B.n794 71.676
R1692 B.n788 B.n73 71.676
R1693 B.n787 B.n786 71.676
R1694 B.n780 B.n75 71.676
R1695 B.n779 B.n778 71.676
R1696 B.n772 B.n77 71.676
R1697 B.n771 B.n770 71.676
R1698 B.n764 B.n79 71.676
R1699 B.n763 B.n762 71.676
R1700 B.n756 B.n81 71.676
R1701 B.n755 B.n754 71.676
R1702 B.n748 B.n83 71.676
R1703 B.n747 B.n746 71.676
R1704 B.n740 B.n85 71.676
R1705 B.n739 B.n89 71.676
R1706 B.n735 B.n734 71.676
R1707 B.n728 B.n91 71.676
R1708 B.n727 B.n726 71.676
R1709 B.n720 B.n93 71.676
R1710 B.n719 B.n97 71.676
R1711 B.n715 B.n714 71.676
R1712 B.n708 B.n99 71.676
R1713 B.n707 B.n706 71.676
R1714 B.n700 B.n101 71.676
R1715 B.n699 B.n698 71.676
R1716 B.n692 B.n103 71.676
R1717 B.n691 B.n690 71.676
R1718 B.n684 B.n105 71.676
R1719 B.n683 B.n682 71.676
R1720 B.n676 B.n107 71.676
R1721 B.n675 B.n674 71.676
R1722 B.n668 B.n109 71.676
R1723 B.n667 B.n666 71.676
R1724 B.n660 B.n111 71.676
R1725 B.n659 B.n658 71.676
R1726 B.n652 B.n113 71.676
R1727 B.n651 B.n650 71.676
R1728 B.n644 B.n115 71.676
R1729 B.n643 B.n642 71.676
R1730 B.n636 B.n117 71.676
R1731 B.n635 B.n634 71.676
R1732 B.n628 B.n119 71.676
R1733 B.n627 B.n626 71.676
R1734 B.n620 B.n121 71.676
R1735 B.n619 B.n618 71.676
R1736 B.n612 B.n123 71.676
R1737 B.n613 B.n612 71.676
R1738 B.n618 B.n617 71.676
R1739 B.n621 B.n620 71.676
R1740 B.n626 B.n625 71.676
R1741 B.n629 B.n628 71.676
R1742 B.n634 B.n633 71.676
R1743 B.n637 B.n636 71.676
R1744 B.n642 B.n641 71.676
R1745 B.n645 B.n644 71.676
R1746 B.n650 B.n649 71.676
R1747 B.n653 B.n652 71.676
R1748 B.n658 B.n657 71.676
R1749 B.n661 B.n660 71.676
R1750 B.n666 B.n665 71.676
R1751 B.n669 B.n668 71.676
R1752 B.n674 B.n673 71.676
R1753 B.n677 B.n676 71.676
R1754 B.n682 B.n681 71.676
R1755 B.n685 B.n684 71.676
R1756 B.n690 B.n689 71.676
R1757 B.n693 B.n692 71.676
R1758 B.n698 B.n697 71.676
R1759 B.n701 B.n700 71.676
R1760 B.n706 B.n705 71.676
R1761 B.n709 B.n708 71.676
R1762 B.n714 B.n713 71.676
R1763 B.n716 B.n97 71.676
R1764 B.n721 B.n720 71.676
R1765 B.n726 B.n725 71.676
R1766 B.n729 B.n728 71.676
R1767 B.n734 B.n733 71.676
R1768 B.n736 B.n89 71.676
R1769 B.n741 B.n740 71.676
R1770 B.n746 B.n745 71.676
R1771 B.n749 B.n748 71.676
R1772 B.n754 B.n753 71.676
R1773 B.n757 B.n756 71.676
R1774 B.n762 B.n761 71.676
R1775 B.n765 B.n764 71.676
R1776 B.n770 B.n769 71.676
R1777 B.n773 B.n772 71.676
R1778 B.n778 B.n777 71.676
R1779 B.n781 B.n780 71.676
R1780 B.n786 B.n785 71.676
R1781 B.n789 B.n788 71.676
R1782 B.n794 B.n793 71.676
R1783 B.n797 B.n796 71.676
R1784 B.n802 B.n801 71.676
R1785 B.n805 B.n804 71.676
R1786 B.n810 B.n809 71.676
R1787 B.n813 B.n812 71.676
R1788 B.n818 B.n817 71.676
R1789 B.n821 B.n820 71.676
R1790 B.n826 B.n825 71.676
R1791 B.n829 B.n828 71.676
R1792 B.n834 B.n833 71.676
R1793 B.n837 B.n836 71.676
R1794 B.n842 B.n841 71.676
R1795 B.n845 B.n844 71.676
R1796 B.n476 B.n182 71.676
R1797 B.n474 B.n184 71.676
R1798 B.n470 B.n469 71.676
R1799 B.n463 B.n186 71.676
R1800 B.n462 B.n461 71.676
R1801 B.n455 B.n188 71.676
R1802 B.n454 B.n453 71.676
R1803 B.n447 B.n190 71.676
R1804 B.n446 B.n445 71.676
R1805 B.n439 B.n192 71.676
R1806 B.n438 B.n437 71.676
R1807 B.n431 B.n194 71.676
R1808 B.n430 B.n429 71.676
R1809 B.n423 B.n196 71.676
R1810 B.n422 B.n421 71.676
R1811 B.n415 B.n198 71.676
R1812 B.n414 B.n413 71.676
R1813 B.n407 B.n200 71.676
R1814 B.n406 B.n405 71.676
R1815 B.n399 B.n202 71.676
R1816 B.n398 B.n397 71.676
R1817 B.n391 B.n204 71.676
R1818 B.n390 B.n389 71.676
R1819 B.n383 B.n206 71.676
R1820 B.n382 B.n381 71.676
R1821 B.n375 B.n208 71.676
R1822 B.n374 B.n373 71.676
R1823 B.n367 B.n210 71.676
R1824 B.n366 B.n365 71.676
R1825 B.n359 B.n215 71.676
R1826 B.n358 B.n357 71.676
R1827 B.n350 B.n217 71.676
R1828 B.n349 B.n348 71.676
R1829 B.n342 B.n221 71.676
R1830 B.n341 B.n340 71.676
R1831 B.n334 B.n223 71.676
R1832 B.n333 B.n332 71.676
R1833 B.n326 B.n225 71.676
R1834 B.n325 B.n324 71.676
R1835 B.n318 B.n227 71.676
R1836 B.n317 B.n316 71.676
R1837 B.n310 B.n229 71.676
R1838 B.n309 B.n308 71.676
R1839 B.n302 B.n231 71.676
R1840 B.n301 B.n300 71.676
R1841 B.n294 B.n233 71.676
R1842 B.n293 B.n292 71.676
R1843 B.n286 B.n235 71.676
R1844 B.n285 B.n284 71.676
R1845 B.n278 B.n237 71.676
R1846 B.n277 B.n276 71.676
R1847 B.n270 B.n239 71.676
R1848 B.n269 B.n268 71.676
R1849 B.n262 B.n241 71.676
R1850 B.n261 B.n260 71.676
R1851 B.n254 B.n243 71.676
R1852 B.n253 B.n252 71.676
R1853 B.n246 B.n245 71.676
R1854 B.n477 B.n476 71.676
R1855 B.n471 B.n184 71.676
R1856 B.n469 B.n468 71.676
R1857 B.n464 B.n463 71.676
R1858 B.n461 B.n460 71.676
R1859 B.n456 B.n455 71.676
R1860 B.n453 B.n452 71.676
R1861 B.n448 B.n447 71.676
R1862 B.n445 B.n444 71.676
R1863 B.n440 B.n439 71.676
R1864 B.n437 B.n436 71.676
R1865 B.n432 B.n431 71.676
R1866 B.n429 B.n428 71.676
R1867 B.n424 B.n423 71.676
R1868 B.n421 B.n420 71.676
R1869 B.n416 B.n415 71.676
R1870 B.n413 B.n412 71.676
R1871 B.n408 B.n407 71.676
R1872 B.n405 B.n404 71.676
R1873 B.n400 B.n399 71.676
R1874 B.n397 B.n396 71.676
R1875 B.n392 B.n391 71.676
R1876 B.n389 B.n388 71.676
R1877 B.n384 B.n383 71.676
R1878 B.n381 B.n380 71.676
R1879 B.n376 B.n375 71.676
R1880 B.n373 B.n372 71.676
R1881 B.n368 B.n367 71.676
R1882 B.n365 B.n364 71.676
R1883 B.n360 B.n359 71.676
R1884 B.n357 B.n356 71.676
R1885 B.n351 B.n350 71.676
R1886 B.n348 B.n347 71.676
R1887 B.n343 B.n342 71.676
R1888 B.n340 B.n339 71.676
R1889 B.n335 B.n334 71.676
R1890 B.n332 B.n331 71.676
R1891 B.n327 B.n326 71.676
R1892 B.n324 B.n323 71.676
R1893 B.n319 B.n318 71.676
R1894 B.n316 B.n315 71.676
R1895 B.n311 B.n310 71.676
R1896 B.n308 B.n307 71.676
R1897 B.n303 B.n302 71.676
R1898 B.n300 B.n299 71.676
R1899 B.n295 B.n294 71.676
R1900 B.n292 B.n291 71.676
R1901 B.n287 B.n286 71.676
R1902 B.n284 B.n283 71.676
R1903 B.n279 B.n278 71.676
R1904 B.n276 B.n275 71.676
R1905 B.n271 B.n270 71.676
R1906 B.n268 B.n267 71.676
R1907 B.n263 B.n262 71.676
R1908 B.n260 B.n259 71.676
R1909 B.n255 B.n254 71.676
R1910 B.n252 B.n251 71.676
R1911 B.n247 B.n246 71.676
R1912 B.n911 B.n910 71.676
R1913 B.n911 B.n2 71.676
R1914 B.n482 B.n181 61.6923
R1915 B.n850 B.n58 61.6923
R1916 B.n88 B.n87 59.5399
R1917 B.n96 B.n95 59.5399
R1918 B.n353 B.n219 59.5399
R1919 B.n213 B.n212 59.5399
R1920 B.n482 B.n177 34.6703
R1921 B.n488 B.n177 34.6703
R1922 B.n488 B.n173 34.6703
R1923 B.n494 B.n173 34.6703
R1924 B.n494 B.n169 34.6703
R1925 B.n500 B.n169 34.6703
R1926 B.n500 B.n165 34.6703
R1927 B.n506 B.n165 34.6703
R1928 B.n512 B.n161 34.6703
R1929 B.n512 B.n157 34.6703
R1930 B.n518 B.n157 34.6703
R1931 B.n518 B.n153 34.6703
R1932 B.n524 B.n153 34.6703
R1933 B.n524 B.n149 34.6703
R1934 B.n530 B.n149 34.6703
R1935 B.n530 B.n145 34.6703
R1936 B.n536 B.n145 34.6703
R1937 B.n536 B.n141 34.6703
R1938 B.n542 B.n141 34.6703
R1939 B.n542 B.n137 34.6703
R1940 B.n549 B.n137 34.6703
R1941 B.n549 B.n548 34.6703
R1942 B.n555 B.n130 34.6703
R1943 B.n562 B.n130 34.6703
R1944 B.n562 B.n126 34.6703
R1945 B.n568 B.n126 34.6703
R1946 B.n568 B.n4 34.6703
R1947 B.n909 B.n4 34.6703
R1948 B.n909 B.n908 34.6703
R1949 B.n908 B.n907 34.6703
R1950 B.n907 B.n8 34.6703
R1951 B.n12 B.n8 34.6703
R1952 B.n900 B.n12 34.6703
R1953 B.n900 B.n899 34.6703
R1954 B.n899 B.n898 34.6703
R1955 B.n892 B.n19 34.6703
R1956 B.n892 B.n891 34.6703
R1957 B.n891 B.n890 34.6703
R1958 B.n890 B.n23 34.6703
R1959 B.n884 B.n23 34.6703
R1960 B.n884 B.n883 34.6703
R1961 B.n883 B.n882 34.6703
R1962 B.n882 B.n30 34.6703
R1963 B.n876 B.n30 34.6703
R1964 B.n876 B.n875 34.6703
R1965 B.n875 B.n874 34.6703
R1966 B.n874 B.n37 34.6703
R1967 B.n868 B.n37 34.6703
R1968 B.n868 B.n867 34.6703
R1969 B.n866 B.n44 34.6703
R1970 B.n860 B.n44 34.6703
R1971 B.n860 B.n859 34.6703
R1972 B.n859 B.n858 34.6703
R1973 B.n858 B.n51 34.6703
R1974 B.n852 B.n51 34.6703
R1975 B.n852 B.n851 34.6703
R1976 B.n851 B.n850 34.6703
R1977 B.n480 B.n479 32.6249
R1978 B.n484 B.n179 32.6249
R1979 B.n614 B.n611 32.6249
R1980 B.n848 B.n847 32.6249
R1981 B.n506 B.t3 32.121
R1982 B.t7 B.n866 32.121
R1983 B.n555 B.t1 23.9634
R1984 B.n898 B.t0 23.9634
R1985 B B.n912 18.0485
R1986 B.n548 B.t1 10.7073
R1987 B.n19 B.t0 10.7073
R1988 B.n480 B.n175 10.6151
R1989 B.n490 B.n175 10.6151
R1990 B.n491 B.n490 10.6151
R1991 B.n492 B.n491 10.6151
R1992 B.n492 B.n167 10.6151
R1993 B.n502 B.n167 10.6151
R1994 B.n503 B.n502 10.6151
R1995 B.n504 B.n503 10.6151
R1996 B.n504 B.n159 10.6151
R1997 B.n514 B.n159 10.6151
R1998 B.n515 B.n514 10.6151
R1999 B.n516 B.n515 10.6151
R2000 B.n516 B.n151 10.6151
R2001 B.n526 B.n151 10.6151
R2002 B.n527 B.n526 10.6151
R2003 B.n528 B.n527 10.6151
R2004 B.n528 B.n143 10.6151
R2005 B.n538 B.n143 10.6151
R2006 B.n539 B.n538 10.6151
R2007 B.n540 B.n539 10.6151
R2008 B.n540 B.n135 10.6151
R2009 B.n551 B.n135 10.6151
R2010 B.n552 B.n551 10.6151
R2011 B.n553 B.n552 10.6151
R2012 B.n553 B.n128 10.6151
R2013 B.n564 B.n128 10.6151
R2014 B.n565 B.n564 10.6151
R2015 B.n566 B.n565 10.6151
R2016 B.n566 B.n0 10.6151
R2017 B.n479 B.n478 10.6151
R2018 B.n478 B.n183 10.6151
R2019 B.n473 B.n183 10.6151
R2020 B.n473 B.n472 10.6151
R2021 B.n472 B.n185 10.6151
R2022 B.n467 B.n185 10.6151
R2023 B.n467 B.n466 10.6151
R2024 B.n466 B.n465 10.6151
R2025 B.n465 B.n187 10.6151
R2026 B.n459 B.n187 10.6151
R2027 B.n459 B.n458 10.6151
R2028 B.n458 B.n457 10.6151
R2029 B.n457 B.n189 10.6151
R2030 B.n451 B.n189 10.6151
R2031 B.n451 B.n450 10.6151
R2032 B.n450 B.n449 10.6151
R2033 B.n449 B.n191 10.6151
R2034 B.n443 B.n191 10.6151
R2035 B.n443 B.n442 10.6151
R2036 B.n442 B.n441 10.6151
R2037 B.n441 B.n193 10.6151
R2038 B.n435 B.n193 10.6151
R2039 B.n435 B.n434 10.6151
R2040 B.n434 B.n433 10.6151
R2041 B.n433 B.n195 10.6151
R2042 B.n427 B.n195 10.6151
R2043 B.n427 B.n426 10.6151
R2044 B.n426 B.n425 10.6151
R2045 B.n425 B.n197 10.6151
R2046 B.n419 B.n197 10.6151
R2047 B.n419 B.n418 10.6151
R2048 B.n418 B.n417 10.6151
R2049 B.n417 B.n199 10.6151
R2050 B.n411 B.n199 10.6151
R2051 B.n411 B.n410 10.6151
R2052 B.n410 B.n409 10.6151
R2053 B.n409 B.n201 10.6151
R2054 B.n403 B.n201 10.6151
R2055 B.n403 B.n402 10.6151
R2056 B.n402 B.n401 10.6151
R2057 B.n401 B.n203 10.6151
R2058 B.n395 B.n203 10.6151
R2059 B.n395 B.n394 10.6151
R2060 B.n394 B.n393 10.6151
R2061 B.n393 B.n205 10.6151
R2062 B.n387 B.n205 10.6151
R2063 B.n387 B.n386 10.6151
R2064 B.n386 B.n385 10.6151
R2065 B.n385 B.n207 10.6151
R2066 B.n379 B.n207 10.6151
R2067 B.n379 B.n378 10.6151
R2068 B.n378 B.n377 10.6151
R2069 B.n377 B.n209 10.6151
R2070 B.n371 B.n370 10.6151
R2071 B.n370 B.n369 10.6151
R2072 B.n369 B.n214 10.6151
R2073 B.n363 B.n214 10.6151
R2074 B.n363 B.n362 10.6151
R2075 B.n362 B.n361 10.6151
R2076 B.n361 B.n216 10.6151
R2077 B.n355 B.n216 10.6151
R2078 B.n355 B.n354 10.6151
R2079 B.n352 B.n220 10.6151
R2080 B.n346 B.n220 10.6151
R2081 B.n346 B.n345 10.6151
R2082 B.n345 B.n344 10.6151
R2083 B.n344 B.n222 10.6151
R2084 B.n338 B.n222 10.6151
R2085 B.n338 B.n337 10.6151
R2086 B.n337 B.n336 10.6151
R2087 B.n336 B.n224 10.6151
R2088 B.n330 B.n224 10.6151
R2089 B.n330 B.n329 10.6151
R2090 B.n329 B.n328 10.6151
R2091 B.n328 B.n226 10.6151
R2092 B.n322 B.n226 10.6151
R2093 B.n322 B.n321 10.6151
R2094 B.n321 B.n320 10.6151
R2095 B.n320 B.n228 10.6151
R2096 B.n314 B.n228 10.6151
R2097 B.n314 B.n313 10.6151
R2098 B.n313 B.n312 10.6151
R2099 B.n312 B.n230 10.6151
R2100 B.n306 B.n230 10.6151
R2101 B.n306 B.n305 10.6151
R2102 B.n305 B.n304 10.6151
R2103 B.n304 B.n232 10.6151
R2104 B.n298 B.n232 10.6151
R2105 B.n298 B.n297 10.6151
R2106 B.n297 B.n296 10.6151
R2107 B.n296 B.n234 10.6151
R2108 B.n290 B.n234 10.6151
R2109 B.n290 B.n289 10.6151
R2110 B.n289 B.n288 10.6151
R2111 B.n288 B.n236 10.6151
R2112 B.n282 B.n236 10.6151
R2113 B.n282 B.n281 10.6151
R2114 B.n281 B.n280 10.6151
R2115 B.n280 B.n238 10.6151
R2116 B.n274 B.n238 10.6151
R2117 B.n274 B.n273 10.6151
R2118 B.n273 B.n272 10.6151
R2119 B.n272 B.n240 10.6151
R2120 B.n266 B.n240 10.6151
R2121 B.n266 B.n265 10.6151
R2122 B.n265 B.n264 10.6151
R2123 B.n264 B.n242 10.6151
R2124 B.n258 B.n242 10.6151
R2125 B.n258 B.n257 10.6151
R2126 B.n257 B.n256 10.6151
R2127 B.n256 B.n244 10.6151
R2128 B.n250 B.n244 10.6151
R2129 B.n250 B.n249 10.6151
R2130 B.n249 B.n248 10.6151
R2131 B.n248 B.n179 10.6151
R2132 B.n485 B.n484 10.6151
R2133 B.n486 B.n485 10.6151
R2134 B.n486 B.n171 10.6151
R2135 B.n496 B.n171 10.6151
R2136 B.n497 B.n496 10.6151
R2137 B.n498 B.n497 10.6151
R2138 B.n498 B.n163 10.6151
R2139 B.n508 B.n163 10.6151
R2140 B.n509 B.n508 10.6151
R2141 B.n510 B.n509 10.6151
R2142 B.n510 B.n155 10.6151
R2143 B.n520 B.n155 10.6151
R2144 B.n521 B.n520 10.6151
R2145 B.n522 B.n521 10.6151
R2146 B.n522 B.n147 10.6151
R2147 B.n532 B.n147 10.6151
R2148 B.n533 B.n532 10.6151
R2149 B.n534 B.n533 10.6151
R2150 B.n534 B.n139 10.6151
R2151 B.n544 B.n139 10.6151
R2152 B.n545 B.n544 10.6151
R2153 B.n546 B.n545 10.6151
R2154 B.n546 B.n132 10.6151
R2155 B.n557 B.n132 10.6151
R2156 B.n558 B.n557 10.6151
R2157 B.n560 B.n558 10.6151
R2158 B.n560 B.n559 10.6151
R2159 B.n559 B.n124 10.6151
R2160 B.n571 B.n124 10.6151
R2161 B.n572 B.n571 10.6151
R2162 B.n573 B.n572 10.6151
R2163 B.n574 B.n573 10.6151
R2164 B.n575 B.n574 10.6151
R2165 B.n578 B.n575 10.6151
R2166 B.n579 B.n578 10.6151
R2167 B.n580 B.n579 10.6151
R2168 B.n581 B.n580 10.6151
R2169 B.n583 B.n581 10.6151
R2170 B.n584 B.n583 10.6151
R2171 B.n585 B.n584 10.6151
R2172 B.n586 B.n585 10.6151
R2173 B.n588 B.n586 10.6151
R2174 B.n589 B.n588 10.6151
R2175 B.n590 B.n589 10.6151
R2176 B.n591 B.n590 10.6151
R2177 B.n593 B.n591 10.6151
R2178 B.n594 B.n593 10.6151
R2179 B.n595 B.n594 10.6151
R2180 B.n596 B.n595 10.6151
R2181 B.n598 B.n596 10.6151
R2182 B.n599 B.n598 10.6151
R2183 B.n600 B.n599 10.6151
R2184 B.n601 B.n600 10.6151
R2185 B.n603 B.n601 10.6151
R2186 B.n604 B.n603 10.6151
R2187 B.n605 B.n604 10.6151
R2188 B.n606 B.n605 10.6151
R2189 B.n608 B.n606 10.6151
R2190 B.n609 B.n608 10.6151
R2191 B.n610 B.n609 10.6151
R2192 B.n611 B.n610 10.6151
R2193 B.n904 B.n1 10.6151
R2194 B.n904 B.n903 10.6151
R2195 B.n903 B.n902 10.6151
R2196 B.n902 B.n10 10.6151
R2197 B.n896 B.n10 10.6151
R2198 B.n896 B.n895 10.6151
R2199 B.n895 B.n894 10.6151
R2200 B.n894 B.n17 10.6151
R2201 B.n888 B.n17 10.6151
R2202 B.n888 B.n887 10.6151
R2203 B.n887 B.n886 10.6151
R2204 B.n886 B.n25 10.6151
R2205 B.n880 B.n25 10.6151
R2206 B.n880 B.n879 10.6151
R2207 B.n879 B.n878 10.6151
R2208 B.n878 B.n32 10.6151
R2209 B.n872 B.n32 10.6151
R2210 B.n872 B.n871 10.6151
R2211 B.n871 B.n870 10.6151
R2212 B.n870 B.n39 10.6151
R2213 B.n864 B.n39 10.6151
R2214 B.n864 B.n863 10.6151
R2215 B.n863 B.n862 10.6151
R2216 B.n862 B.n46 10.6151
R2217 B.n856 B.n46 10.6151
R2218 B.n856 B.n855 10.6151
R2219 B.n855 B.n854 10.6151
R2220 B.n854 B.n53 10.6151
R2221 B.n848 B.n53 10.6151
R2222 B.n847 B.n846 10.6151
R2223 B.n846 B.n60 10.6151
R2224 B.n840 B.n60 10.6151
R2225 B.n840 B.n839 10.6151
R2226 B.n839 B.n838 10.6151
R2227 B.n838 B.n62 10.6151
R2228 B.n832 B.n62 10.6151
R2229 B.n832 B.n831 10.6151
R2230 B.n831 B.n830 10.6151
R2231 B.n830 B.n64 10.6151
R2232 B.n824 B.n64 10.6151
R2233 B.n824 B.n823 10.6151
R2234 B.n823 B.n822 10.6151
R2235 B.n822 B.n66 10.6151
R2236 B.n816 B.n66 10.6151
R2237 B.n816 B.n815 10.6151
R2238 B.n815 B.n814 10.6151
R2239 B.n814 B.n68 10.6151
R2240 B.n808 B.n68 10.6151
R2241 B.n808 B.n807 10.6151
R2242 B.n807 B.n806 10.6151
R2243 B.n806 B.n70 10.6151
R2244 B.n800 B.n70 10.6151
R2245 B.n800 B.n799 10.6151
R2246 B.n799 B.n798 10.6151
R2247 B.n798 B.n72 10.6151
R2248 B.n792 B.n72 10.6151
R2249 B.n792 B.n791 10.6151
R2250 B.n791 B.n790 10.6151
R2251 B.n790 B.n74 10.6151
R2252 B.n784 B.n74 10.6151
R2253 B.n784 B.n783 10.6151
R2254 B.n783 B.n782 10.6151
R2255 B.n782 B.n76 10.6151
R2256 B.n776 B.n76 10.6151
R2257 B.n776 B.n775 10.6151
R2258 B.n775 B.n774 10.6151
R2259 B.n774 B.n78 10.6151
R2260 B.n768 B.n78 10.6151
R2261 B.n768 B.n767 10.6151
R2262 B.n767 B.n766 10.6151
R2263 B.n766 B.n80 10.6151
R2264 B.n760 B.n80 10.6151
R2265 B.n760 B.n759 10.6151
R2266 B.n759 B.n758 10.6151
R2267 B.n758 B.n82 10.6151
R2268 B.n752 B.n82 10.6151
R2269 B.n752 B.n751 10.6151
R2270 B.n751 B.n750 10.6151
R2271 B.n750 B.n84 10.6151
R2272 B.n744 B.n84 10.6151
R2273 B.n744 B.n743 10.6151
R2274 B.n743 B.n742 10.6151
R2275 B.n738 B.n737 10.6151
R2276 B.n737 B.n90 10.6151
R2277 B.n732 B.n90 10.6151
R2278 B.n732 B.n731 10.6151
R2279 B.n731 B.n730 10.6151
R2280 B.n730 B.n92 10.6151
R2281 B.n724 B.n92 10.6151
R2282 B.n724 B.n723 10.6151
R2283 B.n723 B.n722 10.6151
R2284 B.n718 B.n717 10.6151
R2285 B.n717 B.n98 10.6151
R2286 B.n712 B.n98 10.6151
R2287 B.n712 B.n711 10.6151
R2288 B.n711 B.n710 10.6151
R2289 B.n710 B.n100 10.6151
R2290 B.n704 B.n100 10.6151
R2291 B.n704 B.n703 10.6151
R2292 B.n703 B.n702 10.6151
R2293 B.n702 B.n102 10.6151
R2294 B.n696 B.n102 10.6151
R2295 B.n696 B.n695 10.6151
R2296 B.n695 B.n694 10.6151
R2297 B.n694 B.n104 10.6151
R2298 B.n688 B.n104 10.6151
R2299 B.n688 B.n687 10.6151
R2300 B.n687 B.n686 10.6151
R2301 B.n686 B.n106 10.6151
R2302 B.n680 B.n106 10.6151
R2303 B.n680 B.n679 10.6151
R2304 B.n679 B.n678 10.6151
R2305 B.n678 B.n108 10.6151
R2306 B.n672 B.n108 10.6151
R2307 B.n672 B.n671 10.6151
R2308 B.n671 B.n670 10.6151
R2309 B.n670 B.n110 10.6151
R2310 B.n664 B.n110 10.6151
R2311 B.n664 B.n663 10.6151
R2312 B.n663 B.n662 10.6151
R2313 B.n662 B.n112 10.6151
R2314 B.n656 B.n112 10.6151
R2315 B.n656 B.n655 10.6151
R2316 B.n655 B.n654 10.6151
R2317 B.n654 B.n114 10.6151
R2318 B.n648 B.n114 10.6151
R2319 B.n648 B.n647 10.6151
R2320 B.n647 B.n646 10.6151
R2321 B.n646 B.n116 10.6151
R2322 B.n640 B.n116 10.6151
R2323 B.n640 B.n639 10.6151
R2324 B.n639 B.n638 10.6151
R2325 B.n638 B.n118 10.6151
R2326 B.n632 B.n118 10.6151
R2327 B.n632 B.n631 10.6151
R2328 B.n631 B.n630 10.6151
R2329 B.n630 B.n120 10.6151
R2330 B.n624 B.n120 10.6151
R2331 B.n624 B.n623 10.6151
R2332 B.n623 B.n622 10.6151
R2333 B.n622 B.n122 10.6151
R2334 B.n616 B.n122 10.6151
R2335 B.n616 B.n615 10.6151
R2336 B.n615 B.n614 10.6151
R2337 B.n213 B.n209 9.36635
R2338 B.n353 B.n352 9.36635
R2339 B.n742 B.n88 9.36635
R2340 B.n718 B.n96 9.36635
R2341 B.n912 B.n0 8.11757
R2342 B.n912 B.n1 8.11757
R2343 B.t3 B.n161 2.54975
R2344 B.n867 B.t7 2.54975
R2345 B.n371 B.n213 1.24928
R2346 B.n354 B.n353 1.24928
R2347 B.n738 B.n88 1.24928
R2348 B.n722 B.n96 1.24928
R2349 VP.n0 VP.t1 202.274
R2350 VP.n0 VP.t0 152.054
R2351 VP VP.n0 0.526373
R2352 VDD1.n84 VDD1.n0 289.615
R2353 VDD1.n173 VDD1.n89 289.615
R2354 VDD1.n85 VDD1.n84 185
R2355 VDD1.n83 VDD1.n82 185
R2356 VDD1.n4 VDD1.n3 185
R2357 VDD1.n77 VDD1.n76 185
R2358 VDD1.n75 VDD1.n6 185
R2359 VDD1.n74 VDD1.n73 185
R2360 VDD1.n9 VDD1.n7 185
R2361 VDD1.n68 VDD1.n67 185
R2362 VDD1.n66 VDD1.n65 185
R2363 VDD1.n13 VDD1.n12 185
R2364 VDD1.n60 VDD1.n59 185
R2365 VDD1.n58 VDD1.n57 185
R2366 VDD1.n17 VDD1.n16 185
R2367 VDD1.n52 VDD1.n51 185
R2368 VDD1.n50 VDD1.n49 185
R2369 VDD1.n21 VDD1.n20 185
R2370 VDD1.n44 VDD1.n43 185
R2371 VDD1.n42 VDD1.n41 185
R2372 VDD1.n25 VDD1.n24 185
R2373 VDD1.n36 VDD1.n35 185
R2374 VDD1.n34 VDD1.n33 185
R2375 VDD1.n29 VDD1.n28 185
R2376 VDD1.n117 VDD1.n116 185
R2377 VDD1.n122 VDD1.n121 185
R2378 VDD1.n124 VDD1.n123 185
R2379 VDD1.n113 VDD1.n112 185
R2380 VDD1.n130 VDD1.n129 185
R2381 VDD1.n132 VDD1.n131 185
R2382 VDD1.n109 VDD1.n108 185
R2383 VDD1.n138 VDD1.n137 185
R2384 VDD1.n140 VDD1.n139 185
R2385 VDD1.n105 VDD1.n104 185
R2386 VDD1.n146 VDD1.n145 185
R2387 VDD1.n148 VDD1.n147 185
R2388 VDD1.n101 VDD1.n100 185
R2389 VDD1.n154 VDD1.n153 185
R2390 VDD1.n156 VDD1.n155 185
R2391 VDD1.n97 VDD1.n96 185
R2392 VDD1.n163 VDD1.n162 185
R2393 VDD1.n164 VDD1.n95 185
R2394 VDD1.n166 VDD1.n165 185
R2395 VDD1.n93 VDD1.n92 185
R2396 VDD1.n172 VDD1.n171 185
R2397 VDD1.n174 VDD1.n173 185
R2398 VDD1.n30 VDD1.t0 147.659
R2399 VDD1.n118 VDD1.t1 147.659
R2400 VDD1.n84 VDD1.n83 104.615
R2401 VDD1.n83 VDD1.n3 104.615
R2402 VDD1.n76 VDD1.n3 104.615
R2403 VDD1.n76 VDD1.n75 104.615
R2404 VDD1.n75 VDD1.n74 104.615
R2405 VDD1.n74 VDD1.n7 104.615
R2406 VDD1.n67 VDD1.n7 104.615
R2407 VDD1.n67 VDD1.n66 104.615
R2408 VDD1.n66 VDD1.n12 104.615
R2409 VDD1.n59 VDD1.n12 104.615
R2410 VDD1.n59 VDD1.n58 104.615
R2411 VDD1.n58 VDD1.n16 104.615
R2412 VDD1.n51 VDD1.n16 104.615
R2413 VDD1.n51 VDD1.n50 104.615
R2414 VDD1.n50 VDD1.n20 104.615
R2415 VDD1.n43 VDD1.n20 104.615
R2416 VDD1.n43 VDD1.n42 104.615
R2417 VDD1.n42 VDD1.n24 104.615
R2418 VDD1.n35 VDD1.n24 104.615
R2419 VDD1.n35 VDD1.n34 104.615
R2420 VDD1.n34 VDD1.n28 104.615
R2421 VDD1.n122 VDD1.n116 104.615
R2422 VDD1.n123 VDD1.n122 104.615
R2423 VDD1.n123 VDD1.n112 104.615
R2424 VDD1.n130 VDD1.n112 104.615
R2425 VDD1.n131 VDD1.n130 104.615
R2426 VDD1.n131 VDD1.n108 104.615
R2427 VDD1.n138 VDD1.n108 104.615
R2428 VDD1.n139 VDD1.n138 104.615
R2429 VDD1.n139 VDD1.n104 104.615
R2430 VDD1.n146 VDD1.n104 104.615
R2431 VDD1.n147 VDD1.n146 104.615
R2432 VDD1.n147 VDD1.n100 104.615
R2433 VDD1.n154 VDD1.n100 104.615
R2434 VDD1.n155 VDD1.n154 104.615
R2435 VDD1.n155 VDD1.n96 104.615
R2436 VDD1.n163 VDD1.n96 104.615
R2437 VDD1.n164 VDD1.n163 104.615
R2438 VDD1.n165 VDD1.n164 104.615
R2439 VDD1.n165 VDD1.n92 104.615
R2440 VDD1.n172 VDD1.n92 104.615
R2441 VDD1.n173 VDD1.n172 104.615
R2442 VDD1 VDD1.n177 98.7375
R2443 VDD1 VDD1.n88 54.008
R2444 VDD1.t0 VDD1.n28 52.3082
R2445 VDD1.t1 VDD1.n116 52.3082
R2446 VDD1.n30 VDD1.n29 15.6677
R2447 VDD1.n118 VDD1.n117 15.6677
R2448 VDD1.n77 VDD1.n6 13.1884
R2449 VDD1.n166 VDD1.n95 13.1884
R2450 VDD1.n78 VDD1.n4 12.8005
R2451 VDD1.n73 VDD1.n8 12.8005
R2452 VDD1.n33 VDD1.n32 12.8005
R2453 VDD1.n121 VDD1.n120 12.8005
R2454 VDD1.n162 VDD1.n161 12.8005
R2455 VDD1.n167 VDD1.n93 12.8005
R2456 VDD1.n82 VDD1.n81 12.0247
R2457 VDD1.n72 VDD1.n9 12.0247
R2458 VDD1.n36 VDD1.n27 12.0247
R2459 VDD1.n124 VDD1.n115 12.0247
R2460 VDD1.n160 VDD1.n97 12.0247
R2461 VDD1.n171 VDD1.n170 12.0247
R2462 VDD1.n85 VDD1.n2 11.249
R2463 VDD1.n69 VDD1.n68 11.249
R2464 VDD1.n37 VDD1.n25 11.249
R2465 VDD1.n125 VDD1.n113 11.249
R2466 VDD1.n157 VDD1.n156 11.249
R2467 VDD1.n174 VDD1.n91 11.249
R2468 VDD1.n86 VDD1.n0 10.4732
R2469 VDD1.n65 VDD1.n11 10.4732
R2470 VDD1.n41 VDD1.n40 10.4732
R2471 VDD1.n129 VDD1.n128 10.4732
R2472 VDD1.n153 VDD1.n99 10.4732
R2473 VDD1.n175 VDD1.n89 10.4732
R2474 VDD1.n64 VDD1.n13 9.69747
R2475 VDD1.n44 VDD1.n23 9.69747
R2476 VDD1.n132 VDD1.n111 9.69747
R2477 VDD1.n152 VDD1.n101 9.69747
R2478 VDD1.n88 VDD1.n87 9.45567
R2479 VDD1.n177 VDD1.n176 9.45567
R2480 VDD1.n56 VDD1.n55 9.3005
R2481 VDD1.n15 VDD1.n14 9.3005
R2482 VDD1.n62 VDD1.n61 9.3005
R2483 VDD1.n64 VDD1.n63 9.3005
R2484 VDD1.n11 VDD1.n10 9.3005
R2485 VDD1.n70 VDD1.n69 9.3005
R2486 VDD1.n72 VDD1.n71 9.3005
R2487 VDD1.n8 VDD1.n5 9.3005
R2488 VDD1.n87 VDD1.n86 9.3005
R2489 VDD1.n2 VDD1.n1 9.3005
R2490 VDD1.n81 VDD1.n80 9.3005
R2491 VDD1.n79 VDD1.n78 9.3005
R2492 VDD1.n54 VDD1.n53 9.3005
R2493 VDD1.n19 VDD1.n18 9.3005
R2494 VDD1.n48 VDD1.n47 9.3005
R2495 VDD1.n46 VDD1.n45 9.3005
R2496 VDD1.n23 VDD1.n22 9.3005
R2497 VDD1.n40 VDD1.n39 9.3005
R2498 VDD1.n38 VDD1.n37 9.3005
R2499 VDD1.n27 VDD1.n26 9.3005
R2500 VDD1.n32 VDD1.n31 9.3005
R2501 VDD1.n176 VDD1.n175 9.3005
R2502 VDD1.n91 VDD1.n90 9.3005
R2503 VDD1.n170 VDD1.n169 9.3005
R2504 VDD1.n168 VDD1.n167 9.3005
R2505 VDD1.n107 VDD1.n106 9.3005
R2506 VDD1.n136 VDD1.n135 9.3005
R2507 VDD1.n134 VDD1.n133 9.3005
R2508 VDD1.n111 VDD1.n110 9.3005
R2509 VDD1.n128 VDD1.n127 9.3005
R2510 VDD1.n126 VDD1.n125 9.3005
R2511 VDD1.n115 VDD1.n114 9.3005
R2512 VDD1.n120 VDD1.n119 9.3005
R2513 VDD1.n142 VDD1.n141 9.3005
R2514 VDD1.n144 VDD1.n143 9.3005
R2515 VDD1.n103 VDD1.n102 9.3005
R2516 VDD1.n150 VDD1.n149 9.3005
R2517 VDD1.n152 VDD1.n151 9.3005
R2518 VDD1.n99 VDD1.n98 9.3005
R2519 VDD1.n158 VDD1.n157 9.3005
R2520 VDD1.n160 VDD1.n159 9.3005
R2521 VDD1.n161 VDD1.n94 9.3005
R2522 VDD1.n61 VDD1.n60 8.92171
R2523 VDD1.n45 VDD1.n21 8.92171
R2524 VDD1.n133 VDD1.n109 8.92171
R2525 VDD1.n149 VDD1.n148 8.92171
R2526 VDD1.n57 VDD1.n15 8.14595
R2527 VDD1.n49 VDD1.n48 8.14595
R2528 VDD1.n137 VDD1.n136 8.14595
R2529 VDD1.n145 VDD1.n103 8.14595
R2530 VDD1.n56 VDD1.n17 7.3702
R2531 VDD1.n52 VDD1.n19 7.3702
R2532 VDD1.n140 VDD1.n107 7.3702
R2533 VDD1.n144 VDD1.n105 7.3702
R2534 VDD1.n53 VDD1.n17 6.59444
R2535 VDD1.n53 VDD1.n52 6.59444
R2536 VDD1.n141 VDD1.n140 6.59444
R2537 VDD1.n141 VDD1.n105 6.59444
R2538 VDD1.n57 VDD1.n56 5.81868
R2539 VDD1.n49 VDD1.n19 5.81868
R2540 VDD1.n137 VDD1.n107 5.81868
R2541 VDD1.n145 VDD1.n144 5.81868
R2542 VDD1.n60 VDD1.n15 5.04292
R2543 VDD1.n48 VDD1.n21 5.04292
R2544 VDD1.n136 VDD1.n109 5.04292
R2545 VDD1.n148 VDD1.n103 5.04292
R2546 VDD1.n31 VDD1.n30 4.38563
R2547 VDD1.n119 VDD1.n118 4.38563
R2548 VDD1.n61 VDD1.n13 4.26717
R2549 VDD1.n45 VDD1.n44 4.26717
R2550 VDD1.n133 VDD1.n132 4.26717
R2551 VDD1.n149 VDD1.n101 4.26717
R2552 VDD1.n88 VDD1.n0 3.49141
R2553 VDD1.n65 VDD1.n64 3.49141
R2554 VDD1.n41 VDD1.n23 3.49141
R2555 VDD1.n129 VDD1.n111 3.49141
R2556 VDD1.n153 VDD1.n152 3.49141
R2557 VDD1.n177 VDD1.n89 3.49141
R2558 VDD1.n86 VDD1.n85 2.71565
R2559 VDD1.n68 VDD1.n11 2.71565
R2560 VDD1.n40 VDD1.n25 2.71565
R2561 VDD1.n128 VDD1.n113 2.71565
R2562 VDD1.n156 VDD1.n99 2.71565
R2563 VDD1.n175 VDD1.n174 2.71565
R2564 VDD1.n82 VDD1.n2 1.93989
R2565 VDD1.n69 VDD1.n9 1.93989
R2566 VDD1.n37 VDD1.n36 1.93989
R2567 VDD1.n125 VDD1.n124 1.93989
R2568 VDD1.n157 VDD1.n97 1.93989
R2569 VDD1.n171 VDD1.n91 1.93989
R2570 VDD1.n81 VDD1.n4 1.16414
R2571 VDD1.n73 VDD1.n72 1.16414
R2572 VDD1.n33 VDD1.n27 1.16414
R2573 VDD1.n121 VDD1.n115 1.16414
R2574 VDD1.n162 VDD1.n160 1.16414
R2575 VDD1.n170 VDD1.n93 1.16414
R2576 VDD1.n78 VDD1.n77 0.388379
R2577 VDD1.n8 VDD1.n6 0.388379
R2578 VDD1.n32 VDD1.n29 0.388379
R2579 VDD1.n120 VDD1.n117 0.388379
R2580 VDD1.n161 VDD1.n95 0.388379
R2581 VDD1.n167 VDD1.n166 0.388379
R2582 VDD1.n87 VDD1.n1 0.155672
R2583 VDD1.n80 VDD1.n1 0.155672
R2584 VDD1.n80 VDD1.n79 0.155672
R2585 VDD1.n79 VDD1.n5 0.155672
R2586 VDD1.n71 VDD1.n5 0.155672
R2587 VDD1.n71 VDD1.n70 0.155672
R2588 VDD1.n70 VDD1.n10 0.155672
R2589 VDD1.n63 VDD1.n10 0.155672
R2590 VDD1.n63 VDD1.n62 0.155672
R2591 VDD1.n62 VDD1.n14 0.155672
R2592 VDD1.n55 VDD1.n14 0.155672
R2593 VDD1.n55 VDD1.n54 0.155672
R2594 VDD1.n54 VDD1.n18 0.155672
R2595 VDD1.n47 VDD1.n18 0.155672
R2596 VDD1.n47 VDD1.n46 0.155672
R2597 VDD1.n46 VDD1.n22 0.155672
R2598 VDD1.n39 VDD1.n22 0.155672
R2599 VDD1.n39 VDD1.n38 0.155672
R2600 VDD1.n38 VDD1.n26 0.155672
R2601 VDD1.n31 VDD1.n26 0.155672
R2602 VDD1.n119 VDD1.n114 0.155672
R2603 VDD1.n126 VDD1.n114 0.155672
R2604 VDD1.n127 VDD1.n126 0.155672
R2605 VDD1.n127 VDD1.n110 0.155672
R2606 VDD1.n134 VDD1.n110 0.155672
R2607 VDD1.n135 VDD1.n134 0.155672
R2608 VDD1.n135 VDD1.n106 0.155672
R2609 VDD1.n142 VDD1.n106 0.155672
R2610 VDD1.n143 VDD1.n142 0.155672
R2611 VDD1.n143 VDD1.n102 0.155672
R2612 VDD1.n150 VDD1.n102 0.155672
R2613 VDD1.n151 VDD1.n150 0.155672
R2614 VDD1.n151 VDD1.n98 0.155672
R2615 VDD1.n158 VDD1.n98 0.155672
R2616 VDD1.n159 VDD1.n158 0.155672
R2617 VDD1.n159 VDD1.n94 0.155672
R2618 VDD1.n168 VDD1.n94 0.155672
R2619 VDD1.n169 VDD1.n168 0.155672
R2620 VDD1.n169 VDD1.n90 0.155672
R2621 VDD1.n176 VDD1.n90 0.155672
C0 VDD1 VDD2 0.781239f
C1 VDD2 VN 3.83555f
C2 VDD2 VTAIL 6.37422f
C3 VDD1 VN 0.148856f
C4 VP VDD2 0.370226f
C5 VDD1 VTAIL 6.31776f
C6 VP VDD1 4.05415f
C7 VN VTAIL 3.35542f
C8 VP VN 6.655991f
C9 VP VTAIL 3.36969f
C10 VDD2 B 5.502325f
C11 VDD1 B 8.769401f
C12 VTAIL B 9.544897f
C13 VN B 12.556869f
C14 VP B 7.76504f
C15 VDD1.n0 B 0.029951f
C16 VDD1.n1 B 0.020333f
C17 VDD1.n2 B 0.010926f
C18 VDD1.n3 B 0.025825f
C19 VDD1.n4 B 0.011569f
C20 VDD1.n5 B 0.020333f
C21 VDD1.n6 B 0.011247f
C22 VDD1.n7 B 0.025825f
C23 VDD1.n8 B 0.010926f
C24 VDD1.n9 B 0.011569f
C25 VDD1.n10 B 0.020333f
C26 VDD1.n11 B 0.010926f
C27 VDD1.n12 B 0.025825f
C28 VDD1.n13 B 0.011569f
C29 VDD1.n14 B 0.020333f
C30 VDD1.n15 B 0.010926f
C31 VDD1.n16 B 0.025825f
C32 VDD1.n17 B 0.011569f
C33 VDD1.n18 B 0.020333f
C34 VDD1.n19 B 0.010926f
C35 VDD1.n20 B 0.025825f
C36 VDD1.n21 B 0.011569f
C37 VDD1.n22 B 0.020333f
C38 VDD1.n23 B 0.010926f
C39 VDD1.n24 B 0.025825f
C40 VDD1.n25 B 0.011569f
C41 VDD1.n26 B 0.020333f
C42 VDD1.n27 B 0.010926f
C43 VDD1.n28 B 0.019369f
C44 VDD1.n29 B 0.015256f
C45 VDD1.t0 B 0.042673f
C46 VDD1.n30 B 0.139242f
C47 VDD1.n31 B 1.44402f
C48 VDD1.n32 B 0.010926f
C49 VDD1.n33 B 0.011569f
C50 VDD1.n34 B 0.025825f
C51 VDD1.n35 B 0.025825f
C52 VDD1.n36 B 0.011569f
C53 VDD1.n37 B 0.010926f
C54 VDD1.n38 B 0.020333f
C55 VDD1.n39 B 0.020333f
C56 VDD1.n40 B 0.010926f
C57 VDD1.n41 B 0.011569f
C58 VDD1.n42 B 0.025825f
C59 VDD1.n43 B 0.025825f
C60 VDD1.n44 B 0.011569f
C61 VDD1.n45 B 0.010926f
C62 VDD1.n46 B 0.020333f
C63 VDD1.n47 B 0.020333f
C64 VDD1.n48 B 0.010926f
C65 VDD1.n49 B 0.011569f
C66 VDD1.n50 B 0.025825f
C67 VDD1.n51 B 0.025825f
C68 VDD1.n52 B 0.011569f
C69 VDD1.n53 B 0.010926f
C70 VDD1.n54 B 0.020333f
C71 VDD1.n55 B 0.020333f
C72 VDD1.n56 B 0.010926f
C73 VDD1.n57 B 0.011569f
C74 VDD1.n58 B 0.025825f
C75 VDD1.n59 B 0.025825f
C76 VDD1.n60 B 0.011569f
C77 VDD1.n61 B 0.010926f
C78 VDD1.n62 B 0.020333f
C79 VDD1.n63 B 0.020333f
C80 VDD1.n64 B 0.010926f
C81 VDD1.n65 B 0.011569f
C82 VDD1.n66 B 0.025825f
C83 VDD1.n67 B 0.025825f
C84 VDD1.n68 B 0.011569f
C85 VDD1.n69 B 0.010926f
C86 VDD1.n70 B 0.020333f
C87 VDD1.n71 B 0.020333f
C88 VDD1.n72 B 0.010926f
C89 VDD1.n73 B 0.011569f
C90 VDD1.n74 B 0.025825f
C91 VDD1.n75 B 0.025825f
C92 VDD1.n76 B 0.025825f
C93 VDD1.n77 B 0.011247f
C94 VDD1.n78 B 0.010926f
C95 VDD1.n79 B 0.020333f
C96 VDD1.n80 B 0.020333f
C97 VDD1.n81 B 0.010926f
C98 VDD1.n82 B 0.011569f
C99 VDD1.n83 B 0.025825f
C100 VDD1.n84 B 0.058333f
C101 VDD1.n85 B 0.011569f
C102 VDD1.n86 B 0.010926f
C103 VDD1.n87 B 0.053109f
C104 VDD1.n88 B 0.04869f
C105 VDD1.n89 B 0.029951f
C106 VDD1.n90 B 0.020333f
C107 VDD1.n91 B 0.010926f
C108 VDD1.n92 B 0.025825f
C109 VDD1.n93 B 0.011569f
C110 VDD1.n94 B 0.020333f
C111 VDD1.n95 B 0.011247f
C112 VDD1.n96 B 0.025825f
C113 VDD1.n97 B 0.011569f
C114 VDD1.n98 B 0.020333f
C115 VDD1.n99 B 0.010926f
C116 VDD1.n100 B 0.025825f
C117 VDD1.n101 B 0.011569f
C118 VDD1.n102 B 0.020333f
C119 VDD1.n103 B 0.010926f
C120 VDD1.n104 B 0.025825f
C121 VDD1.n105 B 0.011569f
C122 VDD1.n106 B 0.020333f
C123 VDD1.n107 B 0.010926f
C124 VDD1.n108 B 0.025825f
C125 VDD1.n109 B 0.011569f
C126 VDD1.n110 B 0.020333f
C127 VDD1.n111 B 0.010926f
C128 VDD1.n112 B 0.025825f
C129 VDD1.n113 B 0.011569f
C130 VDD1.n114 B 0.020333f
C131 VDD1.n115 B 0.010926f
C132 VDD1.n116 B 0.019369f
C133 VDD1.n117 B 0.015256f
C134 VDD1.t1 B 0.042673f
C135 VDD1.n118 B 0.139242f
C136 VDD1.n119 B 1.44402f
C137 VDD1.n120 B 0.010926f
C138 VDD1.n121 B 0.011569f
C139 VDD1.n122 B 0.025825f
C140 VDD1.n123 B 0.025825f
C141 VDD1.n124 B 0.011569f
C142 VDD1.n125 B 0.010926f
C143 VDD1.n126 B 0.020333f
C144 VDD1.n127 B 0.020333f
C145 VDD1.n128 B 0.010926f
C146 VDD1.n129 B 0.011569f
C147 VDD1.n130 B 0.025825f
C148 VDD1.n131 B 0.025825f
C149 VDD1.n132 B 0.011569f
C150 VDD1.n133 B 0.010926f
C151 VDD1.n134 B 0.020333f
C152 VDD1.n135 B 0.020333f
C153 VDD1.n136 B 0.010926f
C154 VDD1.n137 B 0.011569f
C155 VDD1.n138 B 0.025825f
C156 VDD1.n139 B 0.025825f
C157 VDD1.n140 B 0.011569f
C158 VDD1.n141 B 0.010926f
C159 VDD1.n142 B 0.020333f
C160 VDD1.n143 B 0.020333f
C161 VDD1.n144 B 0.010926f
C162 VDD1.n145 B 0.011569f
C163 VDD1.n146 B 0.025825f
C164 VDD1.n147 B 0.025825f
C165 VDD1.n148 B 0.011569f
C166 VDD1.n149 B 0.010926f
C167 VDD1.n150 B 0.020333f
C168 VDD1.n151 B 0.020333f
C169 VDD1.n152 B 0.010926f
C170 VDD1.n153 B 0.011569f
C171 VDD1.n154 B 0.025825f
C172 VDD1.n155 B 0.025825f
C173 VDD1.n156 B 0.011569f
C174 VDD1.n157 B 0.010926f
C175 VDD1.n158 B 0.020333f
C176 VDD1.n159 B 0.020333f
C177 VDD1.n160 B 0.010926f
C178 VDD1.n161 B 0.010926f
C179 VDD1.n162 B 0.011569f
C180 VDD1.n163 B 0.025825f
C181 VDD1.n164 B 0.025825f
C182 VDD1.n165 B 0.025825f
C183 VDD1.n166 B 0.011247f
C184 VDD1.n167 B 0.010926f
C185 VDD1.n168 B 0.020333f
C186 VDD1.n169 B 0.020333f
C187 VDD1.n170 B 0.010926f
C188 VDD1.n171 B 0.011569f
C189 VDD1.n172 B 0.025825f
C190 VDD1.n173 B 0.058333f
C191 VDD1.n174 B 0.011569f
C192 VDD1.n175 B 0.010926f
C193 VDD1.n176 B 0.053109f
C194 VDD1.n177 B 0.795516f
C195 VP.t1 B 5.022779f
C196 VP.t0 B 4.3397f
C197 VP.n0 B 4.74369f
C198 VDD2.n0 B 0.029589f
C199 VDD2.n1 B 0.020087f
C200 VDD2.n2 B 0.010794f
C201 VDD2.n3 B 0.025513f
C202 VDD2.n4 B 0.011429f
C203 VDD2.n5 B 0.020087f
C204 VDD2.n6 B 0.011111f
C205 VDD2.n7 B 0.025513f
C206 VDD2.n8 B 0.011429f
C207 VDD2.n9 B 0.020087f
C208 VDD2.n10 B 0.010794f
C209 VDD2.n11 B 0.025513f
C210 VDD2.n12 B 0.011429f
C211 VDD2.n13 B 0.020087f
C212 VDD2.n14 B 0.010794f
C213 VDD2.n15 B 0.025513f
C214 VDD2.n16 B 0.011429f
C215 VDD2.n17 B 0.020087f
C216 VDD2.n18 B 0.010794f
C217 VDD2.n19 B 0.025513f
C218 VDD2.n20 B 0.011429f
C219 VDD2.n21 B 0.020087f
C220 VDD2.n22 B 0.010794f
C221 VDD2.n23 B 0.025513f
C222 VDD2.n24 B 0.011429f
C223 VDD2.n25 B 0.020087f
C224 VDD2.n26 B 0.010794f
C225 VDD2.n27 B 0.019134f
C226 VDD2.n28 B 0.015071f
C227 VDD2.t1 B 0.042157f
C228 VDD2.n29 B 0.137557f
C229 VDD2.n30 B 1.42655f
C230 VDD2.n31 B 0.010794f
C231 VDD2.n32 B 0.011429f
C232 VDD2.n33 B 0.025513f
C233 VDD2.n34 B 0.025513f
C234 VDD2.n35 B 0.011429f
C235 VDD2.n36 B 0.010794f
C236 VDD2.n37 B 0.020087f
C237 VDD2.n38 B 0.020087f
C238 VDD2.n39 B 0.010794f
C239 VDD2.n40 B 0.011429f
C240 VDD2.n41 B 0.025513f
C241 VDD2.n42 B 0.025513f
C242 VDD2.n43 B 0.011429f
C243 VDD2.n44 B 0.010794f
C244 VDD2.n45 B 0.020087f
C245 VDD2.n46 B 0.020087f
C246 VDD2.n47 B 0.010794f
C247 VDD2.n48 B 0.011429f
C248 VDD2.n49 B 0.025513f
C249 VDD2.n50 B 0.025513f
C250 VDD2.n51 B 0.011429f
C251 VDD2.n52 B 0.010794f
C252 VDD2.n53 B 0.020087f
C253 VDD2.n54 B 0.020087f
C254 VDD2.n55 B 0.010794f
C255 VDD2.n56 B 0.011429f
C256 VDD2.n57 B 0.025513f
C257 VDD2.n58 B 0.025513f
C258 VDD2.n59 B 0.011429f
C259 VDD2.n60 B 0.010794f
C260 VDD2.n61 B 0.020087f
C261 VDD2.n62 B 0.020087f
C262 VDD2.n63 B 0.010794f
C263 VDD2.n64 B 0.011429f
C264 VDD2.n65 B 0.025513f
C265 VDD2.n66 B 0.025513f
C266 VDD2.n67 B 0.011429f
C267 VDD2.n68 B 0.010794f
C268 VDD2.n69 B 0.020087f
C269 VDD2.n70 B 0.020087f
C270 VDD2.n71 B 0.010794f
C271 VDD2.n72 B 0.010794f
C272 VDD2.n73 B 0.011429f
C273 VDD2.n74 B 0.025513f
C274 VDD2.n75 B 0.025513f
C275 VDD2.n76 B 0.025513f
C276 VDD2.n77 B 0.011111f
C277 VDD2.n78 B 0.010794f
C278 VDD2.n79 B 0.020087f
C279 VDD2.n80 B 0.020087f
C280 VDD2.n81 B 0.010794f
C281 VDD2.n82 B 0.011429f
C282 VDD2.n83 B 0.025513f
C283 VDD2.n84 B 0.057627f
C284 VDD2.n85 B 0.011429f
C285 VDD2.n86 B 0.010794f
C286 VDD2.n87 B 0.052467f
C287 VDD2.n88 B 0.738678f
C288 VDD2.n89 B 0.029589f
C289 VDD2.n90 B 0.020087f
C290 VDD2.n91 B 0.010794f
C291 VDD2.n92 B 0.025513f
C292 VDD2.n93 B 0.011429f
C293 VDD2.n94 B 0.020087f
C294 VDD2.n95 B 0.011111f
C295 VDD2.n96 B 0.025513f
C296 VDD2.n97 B 0.010794f
C297 VDD2.n98 B 0.011429f
C298 VDD2.n99 B 0.020087f
C299 VDD2.n100 B 0.010794f
C300 VDD2.n101 B 0.025513f
C301 VDD2.n102 B 0.011429f
C302 VDD2.n103 B 0.020087f
C303 VDD2.n104 B 0.010794f
C304 VDD2.n105 B 0.025513f
C305 VDD2.n106 B 0.011429f
C306 VDD2.n107 B 0.020087f
C307 VDD2.n108 B 0.010794f
C308 VDD2.n109 B 0.025513f
C309 VDD2.n110 B 0.011429f
C310 VDD2.n111 B 0.020087f
C311 VDD2.n112 B 0.010794f
C312 VDD2.n113 B 0.025513f
C313 VDD2.n114 B 0.011429f
C314 VDD2.n115 B 0.020087f
C315 VDD2.n116 B 0.010794f
C316 VDD2.n117 B 0.019134f
C317 VDD2.n118 B 0.015071f
C318 VDD2.t0 B 0.042157f
C319 VDD2.n119 B 0.137558f
C320 VDD2.n120 B 1.42655f
C321 VDD2.n121 B 0.010794f
C322 VDD2.n122 B 0.011429f
C323 VDD2.n123 B 0.025513f
C324 VDD2.n124 B 0.025513f
C325 VDD2.n125 B 0.011429f
C326 VDD2.n126 B 0.010794f
C327 VDD2.n127 B 0.020087f
C328 VDD2.n128 B 0.020087f
C329 VDD2.n129 B 0.010794f
C330 VDD2.n130 B 0.011429f
C331 VDD2.n131 B 0.025513f
C332 VDD2.n132 B 0.025513f
C333 VDD2.n133 B 0.011429f
C334 VDD2.n134 B 0.010794f
C335 VDD2.n135 B 0.020087f
C336 VDD2.n136 B 0.020087f
C337 VDD2.n137 B 0.010794f
C338 VDD2.n138 B 0.011429f
C339 VDD2.n139 B 0.025513f
C340 VDD2.n140 B 0.025513f
C341 VDD2.n141 B 0.011429f
C342 VDD2.n142 B 0.010794f
C343 VDD2.n143 B 0.020087f
C344 VDD2.n144 B 0.020087f
C345 VDD2.n145 B 0.010794f
C346 VDD2.n146 B 0.011429f
C347 VDD2.n147 B 0.025513f
C348 VDD2.n148 B 0.025513f
C349 VDD2.n149 B 0.011429f
C350 VDD2.n150 B 0.010794f
C351 VDD2.n151 B 0.020087f
C352 VDD2.n152 B 0.020087f
C353 VDD2.n153 B 0.010794f
C354 VDD2.n154 B 0.011429f
C355 VDD2.n155 B 0.025513f
C356 VDD2.n156 B 0.025513f
C357 VDD2.n157 B 0.011429f
C358 VDD2.n158 B 0.010794f
C359 VDD2.n159 B 0.020087f
C360 VDD2.n160 B 0.020087f
C361 VDD2.n161 B 0.010794f
C362 VDD2.n162 B 0.011429f
C363 VDD2.n163 B 0.025513f
C364 VDD2.n164 B 0.025513f
C365 VDD2.n165 B 0.025513f
C366 VDD2.n166 B 0.011111f
C367 VDD2.n167 B 0.010794f
C368 VDD2.n168 B 0.020087f
C369 VDD2.n169 B 0.020087f
C370 VDD2.n170 B 0.010794f
C371 VDD2.n171 B 0.011429f
C372 VDD2.n172 B 0.025513f
C373 VDD2.n173 B 0.057627f
C374 VDD2.n174 B 0.011429f
C375 VDD2.n175 B 0.010794f
C376 VDD2.n176 B 0.052467f
C377 VDD2.n177 B 0.046495f
C378 VDD2.n178 B 2.9753f
C379 VTAIL.n0 B 0.029876f
C380 VTAIL.n1 B 0.020282f
C381 VTAIL.n2 B 0.010899f
C382 VTAIL.n3 B 0.02576f
C383 VTAIL.n4 B 0.01154f
C384 VTAIL.n5 B 0.020282f
C385 VTAIL.n6 B 0.011219f
C386 VTAIL.n7 B 0.02576f
C387 VTAIL.n8 B 0.01154f
C388 VTAIL.n9 B 0.020282f
C389 VTAIL.n10 B 0.010899f
C390 VTAIL.n11 B 0.02576f
C391 VTAIL.n12 B 0.01154f
C392 VTAIL.n13 B 0.020282f
C393 VTAIL.n14 B 0.010899f
C394 VTAIL.n15 B 0.02576f
C395 VTAIL.n16 B 0.01154f
C396 VTAIL.n17 B 0.020282f
C397 VTAIL.n18 B 0.010899f
C398 VTAIL.n19 B 0.02576f
C399 VTAIL.n20 B 0.01154f
C400 VTAIL.n21 B 0.020282f
C401 VTAIL.n22 B 0.010899f
C402 VTAIL.n23 B 0.02576f
C403 VTAIL.n24 B 0.01154f
C404 VTAIL.n25 B 0.020282f
C405 VTAIL.n26 B 0.010899f
C406 VTAIL.n27 B 0.01932f
C407 VTAIL.n28 B 0.015217f
C408 VTAIL.t1 B 0.042566f
C409 VTAIL.n29 B 0.138893f
C410 VTAIL.n30 B 1.4404f
C411 VTAIL.n31 B 0.010899f
C412 VTAIL.n32 B 0.01154f
C413 VTAIL.n33 B 0.02576f
C414 VTAIL.n34 B 0.02576f
C415 VTAIL.n35 B 0.01154f
C416 VTAIL.n36 B 0.010899f
C417 VTAIL.n37 B 0.020282f
C418 VTAIL.n38 B 0.020282f
C419 VTAIL.n39 B 0.010899f
C420 VTAIL.n40 B 0.01154f
C421 VTAIL.n41 B 0.02576f
C422 VTAIL.n42 B 0.02576f
C423 VTAIL.n43 B 0.01154f
C424 VTAIL.n44 B 0.010899f
C425 VTAIL.n45 B 0.020282f
C426 VTAIL.n46 B 0.020282f
C427 VTAIL.n47 B 0.010899f
C428 VTAIL.n48 B 0.01154f
C429 VTAIL.n49 B 0.02576f
C430 VTAIL.n50 B 0.02576f
C431 VTAIL.n51 B 0.01154f
C432 VTAIL.n52 B 0.010899f
C433 VTAIL.n53 B 0.020282f
C434 VTAIL.n54 B 0.020282f
C435 VTAIL.n55 B 0.010899f
C436 VTAIL.n56 B 0.01154f
C437 VTAIL.n57 B 0.02576f
C438 VTAIL.n58 B 0.02576f
C439 VTAIL.n59 B 0.01154f
C440 VTAIL.n60 B 0.010899f
C441 VTAIL.n61 B 0.020282f
C442 VTAIL.n62 B 0.020282f
C443 VTAIL.n63 B 0.010899f
C444 VTAIL.n64 B 0.01154f
C445 VTAIL.n65 B 0.02576f
C446 VTAIL.n66 B 0.02576f
C447 VTAIL.n67 B 0.01154f
C448 VTAIL.n68 B 0.010899f
C449 VTAIL.n69 B 0.020282f
C450 VTAIL.n70 B 0.020282f
C451 VTAIL.n71 B 0.010899f
C452 VTAIL.n72 B 0.010899f
C453 VTAIL.n73 B 0.01154f
C454 VTAIL.n74 B 0.02576f
C455 VTAIL.n75 B 0.02576f
C456 VTAIL.n76 B 0.02576f
C457 VTAIL.n77 B 0.011219f
C458 VTAIL.n78 B 0.010899f
C459 VTAIL.n79 B 0.020282f
C460 VTAIL.n80 B 0.020282f
C461 VTAIL.n81 B 0.010899f
C462 VTAIL.n82 B 0.01154f
C463 VTAIL.n83 B 0.02576f
C464 VTAIL.n84 B 0.058186f
C465 VTAIL.n85 B 0.01154f
C466 VTAIL.n86 B 0.010899f
C467 VTAIL.n87 B 0.052976f
C468 VTAIL.n88 B 0.032984f
C469 VTAIL.n89 B 1.73079f
C470 VTAIL.n90 B 0.029876f
C471 VTAIL.n91 B 0.020282f
C472 VTAIL.n92 B 0.010899f
C473 VTAIL.n93 B 0.02576f
C474 VTAIL.n94 B 0.01154f
C475 VTAIL.n95 B 0.020282f
C476 VTAIL.n96 B 0.011219f
C477 VTAIL.n97 B 0.02576f
C478 VTAIL.n98 B 0.010899f
C479 VTAIL.n99 B 0.01154f
C480 VTAIL.n100 B 0.020282f
C481 VTAIL.n101 B 0.010899f
C482 VTAIL.n102 B 0.02576f
C483 VTAIL.n103 B 0.01154f
C484 VTAIL.n104 B 0.020282f
C485 VTAIL.n105 B 0.010899f
C486 VTAIL.n106 B 0.02576f
C487 VTAIL.n107 B 0.01154f
C488 VTAIL.n108 B 0.020282f
C489 VTAIL.n109 B 0.010899f
C490 VTAIL.n110 B 0.02576f
C491 VTAIL.n111 B 0.01154f
C492 VTAIL.n112 B 0.020282f
C493 VTAIL.n113 B 0.010899f
C494 VTAIL.n114 B 0.02576f
C495 VTAIL.n115 B 0.01154f
C496 VTAIL.n116 B 0.020282f
C497 VTAIL.n117 B 0.010899f
C498 VTAIL.n118 B 0.01932f
C499 VTAIL.n119 B 0.015217f
C500 VTAIL.t2 B 0.042566f
C501 VTAIL.n120 B 0.138893f
C502 VTAIL.n121 B 1.4404f
C503 VTAIL.n122 B 0.010899f
C504 VTAIL.n123 B 0.01154f
C505 VTAIL.n124 B 0.02576f
C506 VTAIL.n125 B 0.02576f
C507 VTAIL.n126 B 0.01154f
C508 VTAIL.n127 B 0.010899f
C509 VTAIL.n128 B 0.020282f
C510 VTAIL.n129 B 0.020282f
C511 VTAIL.n130 B 0.010899f
C512 VTAIL.n131 B 0.01154f
C513 VTAIL.n132 B 0.02576f
C514 VTAIL.n133 B 0.02576f
C515 VTAIL.n134 B 0.01154f
C516 VTAIL.n135 B 0.010899f
C517 VTAIL.n136 B 0.020282f
C518 VTAIL.n137 B 0.020282f
C519 VTAIL.n138 B 0.010899f
C520 VTAIL.n139 B 0.01154f
C521 VTAIL.n140 B 0.02576f
C522 VTAIL.n141 B 0.02576f
C523 VTAIL.n142 B 0.01154f
C524 VTAIL.n143 B 0.010899f
C525 VTAIL.n144 B 0.020282f
C526 VTAIL.n145 B 0.020282f
C527 VTAIL.n146 B 0.010899f
C528 VTAIL.n147 B 0.01154f
C529 VTAIL.n148 B 0.02576f
C530 VTAIL.n149 B 0.02576f
C531 VTAIL.n150 B 0.01154f
C532 VTAIL.n151 B 0.010899f
C533 VTAIL.n152 B 0.020282f
C534 VTAIL.n153 B 0.020282f
C535 VTAIL.n154 B 0.010899f
C536 VTAIL.n155 B 0.01154f
C537 VTAIL.n156 B 0.02576f
C538 VTAIL.n157 B 0.02576f
C539 VTAIL.n158 B 0.01154f
C540 VTAIL.n159 B 0.010899f
C541 VTAIL.n160 B 0.020282f
C542 VTAIL.n161 B 0.020282f
C543 VTAIL.n162 B 0.010899f
C544 VTAIL.n163 B 0.01154f
C545 VTAIL.n164 B 0.02576f
C546 VTAIL.n165 B 0.02576f
C547 VTAIL.n166 B 0.02576f
C548 VTAIL.n167 B 0.011219f
C549 VTAIL.n168 B 0.010899f
C550 VTAIL.n169 B 0.020282f
C551 VTAIL.n170 B 0.020282f
C552 VTAIL.n171 B 0.010899f
C553 VTAIL.n172 B 0.01154f
C554 VTAIL.n173 B 0.02576f
C555 VTAIL.n174 B 0.058186f
C556 VTAIL.n175 B 0.01154f
C557 VTAIL.n176 B 0.010899f
C558 VTAIL.n177 B 0.052976f
C559 VTAIL.n178 B 0.032984f
C560 VTAIL.n179 B 1.78051f
C561 VTAIL.n180 B 0.029876f
C562 VTAIL.n181 B 0.020282f
C563 VTAIL.n182 B 0.010899f
C564 VTAIL.n183 B 0.02576f
C565 VTAIL.n184 B 0.01154f
C566 VTAIL.n185 B 0.020282f
C567 VTAIL.n186 B 0.011219f
C568 VTAIL.n187 B 0.02576f
C569 VTAIL.n188 B 0.010899f
C570 VTAIL.n189 B 0.01154f
C571 VTAIL.n190 B 0.020282f
C572 VTAIL.n191 B 0.010899f
C573 VTAIL.n192 B 0.02576f
C574 VTAIL.n193 B 0.01154f
C575 VTAIL.n194 B 0.020282f
C576 VTAIL.n195 B 0.010899f
C577 VTAIL.n196 B 0.02576f
C578 VTAIL.n197 B 0.01154f
C579 VTAIL.n198 B 0.020282f
C580 VTAIL.n199 B 0.010899f
C581 VTAIL.n200 B 0.02576f
C582 VTAIL.n201 B 0.01154f
C583 VTAIL.n202 B 0.020282f
C584 VTAIL.n203 B 0.010899f
C585 VTAIL.n204 B 0.02576f
C586 VTAIL.n205 B 0.01154f
C587 VTAIL.n206 B 0.020282f
C588 VTAIL.n207 B 0.010899f
C589 VTAIL.n208 B 0.01932f
C590 VTAIL.n209 B 0.015217f
C591 VTAIL.t0 B 0.042566f
C592 VTAIL.n210 B 0.138893f
C593 VTAIL.n211 B 1.4404f
C594 VTAIL.n212 B 0.010899f
C595 VTAIL.n213 B 0.01154f
C596 VTAIL.n214 B 0.02576f
C597 VTAIL.n215 B 0.02576f
C598 VTAIL.n216 B 0.01154f
C599 VTAIL.n217 B 0.010899f
C600 VTAIL.n218 B 0.020282f
C601 VTAIL.n219 B 0.020282f
C602 VTAIL.n220 B 0.010899f
C603 VTAIL.n221 B 0.01154f
C604 VTAIL.n222 B 0.02576f
C605 VTAIL.n223 B 0.02576f
C606 VTAIL.n224 B 0.01154f
C607 VTAIL.n225 B 0.010899f
C608 VTAIL.n226 B 0.020282f
C609 VTAIL.n227 B 0.020282f
C610 VTAIL.n228 B 0.010899f
C611 VTAIL.n229 B 0.01154f
C612 VTAIL.n230 B 0.02576f
C613 VTAIL.n231 B 0.02576f
C614 VTAIL.n232 B 0.01154f
C615 VTAIL.n233 B 0.010899f
C616 VTAIL.n234 B 0.020282f
C617 VTAIL.n235 B 0.020282f
C618 VTAIL.n236 B 0.010899f
C619 VTAIL.n237 B 0.01154f
C620 VTAIL.n238 B 0.02576f
C621 VTAIL.n239 B 0.02576f
C622 VTAIL.n240 B 0.01154f
C623 VTAIL.n241 B 0.010899f
C624 VTAIL.n242 B 0.020282f
C625 VTAIL.n243 B 0.020282f
C626 VTAIL.n244 B 0.010899f
C627 VTAIL.n245 B 0.01154f
C628 VTAIL.n246 B 0.02576f
C629 VTAIL.n247 B 0.02576f
C630 VTAIL.n248 B 0.01154f
C631 VTAIL.n249 B 0.010899f
C632 VTAIL.n250 B 0.020282f
C633 VTAIL.n251 B 0.020282f
C634 VTAIL.n252 B 0.010899f
C635 VTAIL.n253 B 0.01154f
C636 VTAIL.n254 B 0.02576f
C637 VTAIL.n255 B 0.02576f
C638 VTAIL.n256 B 0.02576f
C639 VTAIL.n257 B 0.011219f
C640 VTAIL.n258 B 0.010899f
C641 VTAIL.n259 B 0.020282f
C642 VTAIL.n260 B 0.020282f
C643 VTAIL.n261 B 0.010899f
C644 VTAIL.n262 B 0.01154f
C645 VTAIL.n263 B 0.02576f
C646 VTAIL.n264 B 0.058186f
C647 VTAIL.n265 B 0.01154f
C648 VTAIL.n266 B 0.010899f
C649 VTAIL.n267 B 0.052976f
C650 VTAIL.n268 B 0.032984f
C651 VTAIL.n269 B 1.56642f
C652 VTAIL.n270 B 0.029876f
C653 VTAIL.n271 B 0.020282f
C654 VTAIL.n272 B 0.010899f
C655 VTAIL.n273 B 0.02576f
C656 VTAIL.n274 B 0.01154f
C657 VTAIL.n275 B 0.020282f
C658 VTAIL.n276 B 0.011219f
C659 VTAIL.n277 B 0.02576f
C660 VTAIL.n278 B 0.01154f
C661 VTAIL.n279 B 0.020282f
C662 VTAIL.n280 B 0.010899f
C663 VTAIL.n281 B 0.02576f
C664 VTAIL.n282 B 0.01154f
C665 VTAIL.n283 B 0.020282f
C666 VTAIL.n284 B 0.010899f
C667 VTAIL.n285 B 0.02576f
C668 VTAIL.n286 B 0.01154f
C669 VTAIL.n287 B 0.020282f
C670 VTAIL.n288 B 0.010899f
C671 VTAIL.n289 B 0.02576f
C672 VTAIL.n290 B 0.01154f
C673 VTAIL.n291 B 0.020282f
C674 VTAIL.n292 B 0.010899f
C675 VTAIL.n293 B 0.02576f
C676 VTAIL.n294 B 0.01154f
C677 VTAIL.n295 B 0.020282f
C678 VTAIL.n296 B 0.010899f
C679 VTAIL.n297 B 0.01932f
C680 VTAIL.n298 B 0.015217f
C681 VTAIL.t3 B 0.042566f
C682 VTAIL.n299 B 0.138893f
C683 VTAIL.n300 B 1.4404f
C684 VTAIL.n301 B 0.010899f
C685 VTAIL.n302 B 0.01154f
C686 VTAIL.n303 B 0.02576f
C687 VTAIL.n304 B 0.02576f
C688 VTAIL.n305 B 0.01154f
C689 VTAIL.n306 B 0.010899f
C690 VTAIL.n307 B 0.020282f
C691 VTAIL.n308 B 0.020282f
C692 VTAIL.n309 B 0.010899f
C693 VTAIL.n310 B 0.01154f
C694 VTAIL.n311 B 0.02576f
C695 VTAIL.n312 B 0.02576f
C696 VTAIL.n313 B 0.01154f
C697 VTAIL.n314 B 0.010899f
C698 VTAIL.n315 B 0.020282f
C699 VTAIL.n316 B 0.020282f
C700 VTAIL.n317 B 0.010899f
C701 VTAIL.n318 B 0.01154f
C702 VTAIL.n319 B 0.02576f
C703 VTAIL.n320 B 0.02576f
C704 VTAIL.n321 B 0.01154f
C705 VTAIL.n322 B 0.010899f
C706 VTAIL.n323 B 0.020282f
C707 VTAIL.n324 B 0.020282f
C708 VTAIL.n325 B 0.010899f
C709 VTAIL.n326 B 0.01154f
C710 VTAIL.n327 B 0.02576f
C711 VTAIL.n328 B 0.02576f
C712 VTAIL.n329 B 0.01154f
C713 VTAIL.n330 B 0.010899f
C714 VTAIL.n331 B 0.020282f
C715 VTAIL.n332 B 0.020282f
C716 VTAIL.n333 B 0.010899f
C717 VTAIL.n334 B 0.01154f
C718 VTAIL.n335 B 0.02576f
C719 VTAIL.n336 B 0.02576f
C720 VTAIL.n337 B 0.01154f
C721 VTAIL.n338 B 0.010899f
C722 VTAIL.n339 B 0.020282f
C723 VTAIL.n340 B 0.020282f
C724 VTAIL.n341 B 0.010899f
C725 VTAIL.n342 B 0.010899f
C726 VTAIL.n343 B 0.01154f
C727 VTAIL.n344 B 0.02576f
C728 VTAIL.n345 B 0.02576f
C729 VTAIL.n346 B 0.02576f
C730 VTAIL.n347 B 0.011219f
C731 VTAIL.n348 B 0.010899f
C732 VTAIL.n349 B 0.020282f
C733 VTAIL.n350 B 0.020282f
C734 VTAIL.n351 B 0.010899f
C735 VTAIL.n352 B 0.01154f
C736 VTAIL.n353 B 0.02576f
C737 VTAIL.n354 B 0.058186f
C738 VTAIL.n355 B 0.01154f
C739 VTAIL.n356 B 0.010899f
C740 VTAIL.n357 B 0.052976f
C741 VTAIL.n358 B 0.032984f
C742 VTAIL.n359 B 1.47839f
C743 VN.t0 B 4.24188f
C744 VN.t1 B 4.904069f
.ends

