* NGSPICE file created from diff_pair_sample_0743.ext - technology: sky130A

.subckt diff_pair_sample_0743 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=1.5639 ps=8.8 w=4.01 l=2.01
X1 B.t11 B.t9 B.t10 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=0 ps=0 w=4.01 l=2.01
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=1.5639 ps=8.8 w=4.01 l=2.01
X3 VDD1.t0 VP.t1 VTAIL.t2 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=1.5639 ps=8.8 w=4.01 l=2.01
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=1.5639 ps=8.8 w=4.01 l=2.01
X5 B.t8 B.t6 B.t7 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=0 ps=0 w=4.01 l=2.01
X6 B.t5 B.t3 B.t4 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=0 ps=0 w=4.01 l=2.01
X7 B.t2 B.t0 B.t1 w_n1906_n1770# sky130_fd_pr__pfet_01v8 ad=1.5639 pd=8.8 as=0 ps=0 w=4.01 l=2.01
R0 VP.n0 VP.t1 143.98
R1 VP.n0 VP.t0 106.942
R2 VP VP.n0 0.241678
R3 VTAIL.n74 VTAIL.n60 756.745
R4 VTAIL.n14 VTAIL.n0 756.745
R5 VTAIL.n54 VTAIL.n40 756.745
R6 VTAIL.n34 VTAIL.n20 756.745
R7 VTAIL.n67 VTAIL.n66 585
R8 VTAIL.n64 VTAIL.n63 585
R9 VTAIL.n73 VTAIL.n72 585
R10 VTAIL.n75 VTAIL.n74 585
R11 VTAIL.n7 VTAIL.n6 585
R12 VTAIL.n4 VTAIL.n3 585
R13 VTAIL.n13 VTAIL.n12 585
R14 VTAIL.n15 VTAIL.n14 585
R15 VTAIL.n55 VTAIL.n54 585
R16 VTAIL.n53 VTAIL.n52 585
R17 VTAIL.n44 VTAIL.n43 585
R18 VTAIL.n47 VTAIL.n46 585
R19 VTAIL.n35 VTAIL.n34 585
R20 VTAIL.n33 VTAIL.n32 585
R21 VTAIL.n24 VTAIL.n23 585
R22 VTAIL.n27 VTAIL.n26 585
R23 VTAIL.t0 VTAIL.n65 330.707
R24 VTAIL.t3 VTAIL.n5 330.707
R25 VTAIL.t2 VTAIL.n45 330.707
R26 VTAIL.t1 VTAIL.n25 330.707
R27 VTAIL.n66 VTAIL.n63 171.744
R28 VTAIL.n73 VTAIL.n63 171.744
R29 VTAIL.n74 VTAIL.n73 171.744
R30 VTAIL.n6 VTAIL.n3 171.744
R31 VTAIL.n13 VTAIL.n3 171.744
R32 VTAIL.n14 VTAIL.n13 171.744
R33 VTAIL.n54 VTAIL.n53 171.744
R34 VTAIL.n53 VTAIL.n43 171.744
R35 VTAIL.n46 VTAIL.n43 171.744
R36 VTAIL.n34 VTAIL.n33 171.744
R37 VTAIL.n33 VTAIL.n23 171.744
R38 VTAIL.n26 VTAIL.n23 171.744
R39 VTAIL.n66 VTAIL.t0 85.8723
R40 VTAIL.n6 VTAIL.t3 85.8723
R41 VTAIL.n46 VTAIL.t2 85.8723
R42 VTAIL.n26 VTAIL.t1 85.8723
R43 VTAIL.n79 VTAIL.n78 35.4823
R44 VTAIL.n19 VTAIL.n18 35.4823
R45 VTAIL.n59 VTAIL.n58 35.4823
R46 VTAIL.n39 VTAIL.n38 35.4823
R47 VTAIL.n39 VTAIL.n19 19.8583
R48 VTAIL.n79 VTAIL.n59 17.841
R49 VTAIL.n67 VTAIL.n65 16.3201
R50 VTAIL.n7 VTAIL.n5 16.3201
R51 VTAIL.n47 VTAIL.n45 16.3201
R52 VTAIL.n27 VTAIL.n25 16.3201
R53 VTAIL.n68 VTAIL.n64 12.8005
R54 VTAIL.n8 VTAIL.n4 12.8005
R55 VTAIL.n48 VTAIL.n44 12.8005
R56 VTAIL.n28 VTAIL.n24 12.8005
R57 VTAIL.n72 VTAIL.n71 12.0247
R58 VTAIL.n12 VTAIL.n11 12.0247
R59 VTAIL.n52 VTAIL.n51 12.0247
R60 VTAIL.n32 VTAIL.n31 12.0247
R61 VTAIL.n75 VTAIL.n62 11.249
R62 VTAIL.n15 VTAIL.n2 11.249
R63 VTAIL.n55 VTAIL.n42 11.249
R64 VTAIL.n35 VTAIL.n22 11.249
R65 VTAIL.n76 VTAIL.n60 10.4732
R66 VTAIL.n16 VTAIL.n0 10.4732
R67 VTAIL.n56 VTAIL.n40 10.4732
R68 VTAIL.n36 VTAIL.n20 10.4732
R69 VTAIL.n78 VTAIL.n77 9.45567
R70 VTAIL.n18 VTAIL.n17 9.45567
R71 VTAIL.n58 VTAIL.n57 9.45567
R72 VTAIL.n38 VTAIL.n37 9.45567
R73 VTAIL.n77 VTAIL.n76 9.3005
R74 VTAIL.n62 VTAIL.n61 9.3005
R75 VTAIL.n71 VTAIL.n70 9.3005
R76 VTAIL.n69 VTAIL.n68 9.3005
R77 VTAIL.n17 VTAIL.n16 9.3005
R78 VTAIL.n2 VTAIL.n1 9.3005
R79 VTAIL.n11 VTAIL.n10 9.3005
R80 VTAIL.n9 VTAIL.n8 9.3005
R81 VTAIL.n57 VTAIL.n56 9.3005
R82 VTAIL.n42 VTAIL.n41 9.3005
R83 VTAIL.n51 VTAIL.n50 9.3005
R84 VTAIL.n49 VTAIL.n48 9.3005
R85 VTAIL.n37 VTAIL.n36 9.3005
R86 VTAIL.n22 VTAIL.n21 9.3005
R87 VTAIL.n31 VTAIL.n30 9.3005
R88 VTAIL.n29 VTAIL.n28 9.3005
R89 VTAIL.n69 VTAIL.n65 3.78097
R90 VTAIL.n9 VTAIL.n5 3.78097
R91 VTAIL.n49 VTAIL.n45 3.78097
R92 VTAIL.n29 VTAIL.n25 3.78097
R93 VTAIL.n78 VTAIL.n60 3.49141
R94 VTAIL.n18 VTAIL.n0 3.49141
R95 VTAIL.n58 VTAIL.n40 3.49141
R96 VTAIL.n38 VTAIL.n20 3.49141
R97 VTAIL.n76 VTAIL.n75 2.71565
R98 VTAIL.n16 VTAIL.n15 2.71565
R99 VTAIL.n56 VTAIL.n55 2.71565
R100 VTAIL.n36 VTAIL.n35 2.71565
R101 VTAIL.n72 VTAIL.n62 1.93989
R102 VTAIL.n12 VTAIL.n2 1.93989
R103 VTAIL.n52 VTAIL.n42 1.93989
R104 VTAIL.n32 VTAIL.n22 1.93989
R105 VTAIL.n59 VTAIL.n39 1.47895
R106 VTAIL.n71 VTAIL.n64 1.16414
R107 VTAIL.n11 VTAIL.n4 1.16414
R108 VTAIL.n51 VTAIL.n44 1.16414
R109 VTAIL.n31 VTAIL.n24 1.16414
R110 VTAIL VTAIL.n19 1.03283
R111 VTAIL VTAIL.n79 0.446621
R112 VTAIL.n68 VTAIL.n67 0.388379
R113 VTAIL.n8 VTAIL.n7 0.388379
R114 VTAIL.n48 VTAIL.n47 0.388379
R115 VTAIL.n28 VTAIL.n27 0.388379
R116 VTAIL.n70 VTAIL.n69 0.155672
R117 VTAIL.n70 VTAIL.n61 0.155672
R118 VTAIL.n77 VTAIL.n61 0.155672
R119 VTAIL.n10 VTAIL.n9 0.155672
R120 VTAIL.n10 VTAIL.n1 0.155672
R121 VTAIL.n17 VTAIL.n1 0.155672
R122 VTAIL.n57 VTAIL.n41 0.155672
R123 VTAIL.n50 VTAIL.n41 0.155672
R124 VTAIL.n50 VTAIL.n49 0.155672
R125 VTAIL.n37 VTAIL.n21 0.155672
R126 VTAIL.n30 VTAIL.n21 0.155672
R127 VTAIL.n30 VTAIL.n29 0.155672
R128 VDD1.n14 VDD1.n0 756.745
R129 VDD1.n33 VDD1.n19 756.745
R130 VDD1.n15 VDD1.n14 585
R131 VDD1.n13 VDD1.n12 585
R132 VDD1.n4 VDD1.n3 585
R133 VDD1.n7 VDD1.n6 585
R134 VDD1.n26 VDD1.n25 585
R135 VDD1.n23 VDD1.n22 585
R136 VDD1.n32 VDD1.n31 585
R137 VDD1.n34 VDD1.n33 585
R138 VDD1.t0 VDD1.n5 330.707
R139 VDD1.t1 VDD1.n24 330.707
R140 VDD1.n14 VDD1.n13 171.744
R141 VDD1.n13 VDD1.n3 171.744
R142 VDD1.n6 VDD1.n3 171.744
R143 VDD1.n25 VDD1.n22 171.744
R144 VDD1.n32 VDD1.n22 171.744
R145 VDD1.n33 VDD1.n32 171.744
R146 VDD1.n6 VDD1.t0 85.8723
R147 VDD1.n25 VDD1.t1 85.8723
R148 VDD1 VDD1.n37 84.3411
R149 VDD1 VDD1.n18 52.7236
R150 VDD1.n7 VDD1.n5 16.3201
R151 VDD1.n26 VDD1.n24 16.3201
R152 VDD1.n8 VDD1.n4 12.8005
R153 VDD1.n27 VDD1.n23 12.8005
R154 VDD1.n12 VDD1.n11 12.0247
R155 VDD1.n31 VDD1.n30 12.0247
R156 VDD1.n15 VDD1.n2 11.249
R157 VDD1.n34 VDD1.n21 11.249
R158 VDD1.n16 VDD1.n0 10.4732
R159 VDD1.n35 VDD1.n19 10.4732
R160 VDD1.n18 VDD1.n17 9.45567
R161 VDD1.n37 VDD1.n36 9.45567
R162 VDD1.n17 VDD1.n16 9.3005
R163 VDD1.n2 VDD1.n1 9.3005
R164 VDD1.n11 VDD1.n10 9.3005
R165 VDD1.n9 VDD1.n8 9.3005
R166 VDD1.n36 VDD1.n35 9.3005
R167 VDD1.n21 VDD1.n20 9.3005
R168 VDD1.n30 VDD1.n29 9.3005
R169 VDD1.n28 VDD1.n27 9.3005
R170 VDD1.n9 VDD1.n5 3.78097
R171 VDD1.n28 VDD1.n24 3.78097
R172 VDD1.n18 VDD1.n0 3.49141
R173 VDD1.n37 VDD1.n19 3.49141
R174 VDD1.n16 VDD1.n15 2.71565
R175 VDD1.n35 VDD1.n34 2.71565
R176 VDD1.n12 VDD1.n2 1.93989
R177 VDD1.n31 VDD1.n21 1.93989
R178 VDD1.n11 VDD1.n4 1.16414
R179 VDD1.n30 VDD1.n23 1.16414
R180 VDD1.n8 VDD1.n7 0.388379
R181 VDD1.n27 VDD1.n26 0.388379
R182 VDD1.n17 VDD1.n1 0.155672
R183 VDD1.n10 VDD1.n1 0.155672
R184 VDD1.n10 VDD1.n9 0.155672
R185 VDD1.n29 VDD1.n28 0.155672
R186 VDD1.n29 VDD1.n20 0.155672
R187 VDD1.n36 VDD1.n20 0.155672
R188 B.n271 B.n40 585
R189 B.n273 B.n272 585
R190 B.n274 B.n39 585
R191 B.n276 B.n275 585
R192 B.n277 B.n38 585
R193 B.n279 B.n278 585
R194 B.n280 B.n37 585
R195 B.n282 B.n281 585
R196 B.n283 B.n36 585
R197 B.n285 B.n284 585
R198 B.n286 B.n35 585
R199 B.n288 B.n287 585
R200 B.n289 B.n34 585
R201 B.n291 B.n290 585
R202 B.n292 B.n33 585
R203 B.n294 B.n293 585
R204 B.n295 B.n32 585
R205 B.n297 B.n296 585
R206 B.n299 B.n29 585
R207 B.n301 B.n300 585
R208 B.n302 B.n28 585
R209 B.n304 B.n303 585
R210 B.n305 B.n27 585
R211 B.n307 B.n306 585
R212 B.n308 B.n26 585
R213 B.n310 B.n309 585
R214 B.n311 B.n25 585
R215 B.n313 B.n312 585
R216 B.n315 B.n314 585
R217 B.n316 B.n21 585
R218 B.n318 B.n317 585
R219 B.n319 B.n20 585
R220 B.n321 B.n320 585
R221 B.n322 B.n19 585
R222 B.n324 B.n323 585
R223 B.n325 B.n18 585
R224 B.n327 B.n326 585
R225 B.n328 B.n17 585
R226 B.n330 B.n329 585
R227 B.n331 B.n16 585
R228 B.n333 B.n332 585
R229 B.n334 B.n15 585
R230 B.n336 B.n335 585
R231 B.n337 B.n14 585
R232 B.n339 B.n338 585
R233 B.n340 B.n13 585
R234 B.n270 B.n269 585
R235 B.n268 B.n41 585
R236 B.n267 B.n266 585
R237 B.n265 B.n42 585
R238 B.n264 B.n263 585
R239 B.n262 B.n43 585
R240 B.n261 B.n260 585
R241 B.n259 B.n44 585
R242 B.n258 B.n257 585
R243 B.n256 B.n45 585
R244 B.n255 B.n254 585
R245 B.n253 B.n46 585
R246 B.n252 B.n251 585
R247 B.n250 B.n47 585
R248 B.n249 B.n248 585
R249 B.n247 B.n48 585
R250 B.n246 B.n245 585
R251 B.n244 B.n49 585
R252 B.n243 B.n242 585
R253 B.n241 B.n50 585
R254 B.n240 B.n239 585
R255 B.n238 B.n51 585
R256 B.n237 B.n236 585
R257 B.n235 B.n52 585
R258 B.n234 B.n233 585
R259 B.n232 B.n53 585
R260 B.n231 B.n230 585
R261 B.n229 B.n54 585
R262 B.n228 B.n227 585
R263 B.n226 B.n55 585
R264 B.n225 B.n224 585
R265 B.n223 B.n56 585
R266 B.n222 B.n221 585
R267 B.n220 B.n57 585
R268 B.n219 B.n218 585
R269 B.n217 B.n58 585
R270 B.n216 B.n215 585
R271 B.n214 B.n59 585
R272 B.n213 B.n212 585
R273 B.n211 B.n60 585
R274 B.n210 B.n209 585
R275 B.n208 B.n61 585
R276 B.n207 B.n206 585
R277 B.n205 B.n62 585
R278 B.n204 B.n203 585
R279 B.n133 B.n90 585
R280 B.n135 B.n134 585
R281 B.n136 B.n89 585
R282 B.n138 B.n137 585
R283 B.n139 B.n88 585
R284 B.n141 B.n140 585
R285 B.n142 B.n87 585
R286 B.n144 B.n143 585
R287 B.n145 B.n86 585
R288 B.n147 B.n146 585
R289 B.n148 B.n85 585
R290 B.n150 B.n149 585
R291 B.n151 B.n84 585
R292 B.n153 B.n152 585
R293 B.n154 B.n83 585
R294 B.n156 B.n155 585
R295 B.n157 B.n82 585
R296 B.n159 B.n158 585
R297 B.n161 B.n79 585
R298 B.n163 B.n162 585
R299 B.n164 B.n78 585
R300 B.n166 B.n165 585
R301 B.n167 B.n77 585
R302 B.n169 B.n168 585
R303 B.n170 B.n76 585
R304 B.n172 B.n171 585
R305 B.n173 B.n75 585
R306 B.n175 B.n174 585
R307 B.n177 B.n176 585
R308 B.n178 B.n71 585
R309 B.n180 B.n179 585
R310 B.n181 B.n70 585
R311 B.n183 B.n182 585
R312 B.n184 B.n69 585
R313 B.n186 B.n185 585
R314 B.n187 B.n68 585
R315 B.n189 B.n188 585
R316 B.n190 B.n67 585
R317 B.n192 B.n191 585
R318 B.n193 B.n66 585
R319 B.n195 B.n194 585
R320 B.n196 B.n65 585
R321 B.n198 B.n197 585
R322 B.n199 B.n64 585
R323 B.n201 B.n200 585
R324 B.n202 B.n63 585
R325 B.n132 B.n131 585
R326 B.n130 B.n91 585
R327 B.n129 B.n128 585
R328 B.n127 B.n92 585
R329 B.n126 B.n125 585
R330 B.n124 B.n93 585
R331 B.n123 B.n122 585
R332 B.n121 B.n94 585
R333 B.n120 B.n119 585
R334 B.n118 B.n95 585
R335 B.n117 B.n116 585
R336 B.n115 B.n96 585
R337 B.n114 B.n113 585
R338 B.n112 B.n97 585
R339 B.n111 B.n110 585
R340 B.n109 B.n98 585
R341 B.n108 B.n107 585
R342 B.n106 B.n99 585
R343 B.n105 B.n104 585
R344 B.n103 B.n100 585
R345 B.n102 B.n101 585
R346 B.n2 B.n0 585
R347 B.n373 B.n1 585
R348 B.n372 B.n371 585
R349 B.n370 B.n3 585
R350 B.n369 B.n368 585
R351 B.n367 B.n4 585
R352 B.n366 B.n365 585
R353 B.n364 B.n5 585
R354 B.n363 B.n362 585
R355 B.n361 B.n6 585
R356 B.n360 B.n359 585
R357 B.n358 B.n7 585
R358 B.n357 B.n356 585
R359 B.n355 B.n8 585
R360 B.n354 B.n353 585
R361 B.n352 B.n9 585
R362 B.n351 B.n350 585
R363 B.n349 B.n10 585
R364 B.n348 B.n347 585
R365 B.n346 B.n11 585
R366 B.n345 B.n344 585
R367 B.n343 B.n12 585
R368 B.n342 B.n341 585
R369 B.n375 B.n374 585
R370 B.n133 B.n132 463.671
R371 B.n342 B.n13 463.671
R372 B.n204 B.n63 463.671
R373 B.n271 B.n270 463.671
R374 B.n72 B.t11 281.205
R375 B.n30 B.t7 281.205
R376 B.n80 B.t2 281.205
R377 B.n22 B.t4 281.205
R378 B.n72 B.t9 255.022
R379 B.n80 B.t0 255.022
R380 B.n22 B.t3 255.022
R381 B.n30 B.t6 255.022
R382 B.n73 B.t10 235.823
R383 B.n31 B.t8 235.823
R384 B.n81 B.t1 235.823
R385 B.n23 B.t5 235.823
R386 B.n132 B.n91 163.367
R387 B.n128 B.n91 163.367
R388 B.n128 B.n127 163.367
R389 B.n127 B.n126 163.367
R390 B.n126 B.n93 163.367
R391 B.n122 B.n93 163.367
R392 B.n122 B.n121 163.367
R393 B.n121 B.n120 163.367
R394 B.n120 B.n95 163.367
R395 B.n116 B.n95 163.367
R396 B.n116 B.n115 163.367
R397 B.n115 B.n114 163.367
R398 B.n114 B.n97 163.367
R399 B.n110 B.n97 163.367
R400 B.n110 B.n109 163.367
R401 B.n109 B.n108 163.367
R402 B.n108 B.n99 163.367
R403 B.n104 B.n99 163.367
R404 B.n104 B.n103 163.367
R405 B.n103 B.n102 163.367
R406 B.n102 B.n2 163.367
R407 B.n374 B.n2 163.367
R408 B.n374 B.n373 163.367
R409 B.n373 B.n372 163.367
R410 B.n372 B.n3 163.367
R411 B.n368 B.n3 163.367
R412 B.n368 B.n367 163.367
R413 B.n367 B.n366 163.367
R414 B.n366 B.n5 163.367
R415 B.n362 B.n5 163.367
R416 B.n362 B.n361 163.367
R417 B.n361 B.n360 163.367
R418 B.n360 B.n7 163.367
R419 B.n356 B.n7 163.367
R420 B.n356 B.n355 163.367
R421 B.n355 B.n354 163.367
R422 B.n354 B.n9 163.367
R423 B.n350 B.n9 163.367
R424 B.n350 B.n349 163.367
R425 B.n349 B.n348 163.367
R426 B.n348 B.n11 163.367
R427 B.n344 B.n11 163.367
R428 B.n344 B.n343 163.367
R429 B.n343 B.n342 163.367
R430 B.n134 B.n133 163.367
R431 B.n134 B.n89 163.367
R432 B.n138 B.n89 163.367
R433 B.n139 B.n138 163.367
R434 B.n140 B.n139 163.367
R435 B.n140 B.n87 163.367
R436 B.n144 B.n87 163.367
R437 B.n145 B.n144 163.367
R438 B.n146 B.n145 163.367
R439 B.n146 B.n85 163.367
R440 B.n150 B.n85 163.367
R441 B.n151 B.n150 163.367
R442 B.n152 B.n151 163.367
R443 B.n152 B.n83 163.367
R444 B.n156 B.n83 163.367
R445 B.n157 B.n156 163.367
R446 B.n158 B.n157 163.367
R447 B.n158 B.n79 163.367
R448 B.n163 B.n79 163.367
R449 B.n164 B.n163 163.367
R450 B.n165 B.n164 163.367
R451 B.n165 B.n77 163.367
R452 B.n169 B.n77 163.367
R453 B.n170 B.n169 163.367
R454 B.n171 B.n170 163.367
R455 B.n171 B.n75 163.367
R456 B.n175 B.n75 163.367
R457 B.n176 B.n175 163.367
R458 B.n176 B.n71 163.367
R459 B.n180 B.n71 163.367
R460 B.n181 B.n180 163.367
R461 B.n182 B.n181 163.367
R462 B.n182 B.n69 163.367
R463 B.n186 B.n69 163.367
R464 B.n187 B.n186 163.367
R465 B.n188 B.n187 163.367
R466 B.n188 B.n67 163.367
R467 B.n192 B.n67 163.367
R468 B.n193 B.n192 163.367
R469 B.n194 B.n193 163.367
R470 B.n194 B.n65 163.367
R471 B.n198 B.n65 163.367
R472 B.n199 B.n198 163.367
R473 B.n200 B.n199 163.367
R474 B.n200 B.n63 163.367
R475 B.n205 B.n204 163.367
R476 B.n206 B.n205 163.367
R477 B.n206 B.n61 163.367
R478 B.n210 B.n61 163.367
R479 B.n211 B.n210 163.367
R480 B.n212 B.n211 163.367
R481 B.n212 B.n59 163.367
R482 B.n216 B.n59 163.367
R483 B.n217 B.n216 163.367
R484 B.n218 B.n217 163.367
R485 B.n218 B.n57 163.367
R486 B.n222 B.n57 163.367
R487 B.n223 B.n222 163.367
R488 B.n224 B.n223 163.367
R489 B.n224 B.n55 163.367
R490 B.n228 B.n55 163.367
R491 B.n229 B.n228 163.367
R492 B.n230 B.n229 163.367
R493 B.n230 B.n53 163.367
R494 B.n234 B.n53 163.367
R495 B.n235 B.n234 163.367
R496 B.n236 B.n235 163.367
R497 B.n236 B.n51 163.367
R498 B.n240 B.n51 163.367
R499 B.n241 B.n240 163.367
R500 B.n242 B.n241 163.367
R501 B.n242 B.n49 163.367
R502 B.n246 B.n49 163.367
R503 B.n247 B.n246 163.367
R504 B.n248 B.n247 163.367
R505 B.n248 B.n47 163.367
R506 B.n252 B.n47 163.367
R507 B.n253 B.n252 163.367
R508 B.n254 B.n253 163.367
R509 B.n254 B.n45 163.367
R510 B.n258 B.n45 163.367
R511 B.n259 B.n258 163.367
R512 B.n260 B.n259 163.367
R513 B.n260 B.n43 163.367
R514 B.n264 B.n43 163.367
R515 B.n265 B.n264 163.367
R516 B.n266 B.n265 163.367
R517 B.n266 B.n41 163.367
R518 B.n270 B.n41 163.367
R519 B.n338 B.n13 163.367
R520 B.n338 B.n337 163.367
R521 B.n337 B.n336 163.367
R522 B.n336 B.n15 163.367
R523 B.n332 B.n15 163.367
R524 B.n332 B.n331 163.367
R525 B.n331 B.n330 163.367
R526 B.n330 B.n17 163.367
R527 B.n326 B.n17 163.367
R528 B.n326 B.n325 163.367
R529 B.n325 B.n324 163.367
R530 B.n324 B.n19 163.367
R531 B.n320 B.n19 163.367
R532 B.n320 B.n319 163.367
R533 B.n319 B.n318 163.367
R534 B.n318 B.n21 163.367
R535 B.n314 B.n21 163.367
R536 B.n314 B.n313 163.367
R537 B.n313 B.n25 163.367
R538 B.n309 B.n25 163.367
R539 B.n309 B.n308 163.367
R540 B.n308 B.n307 163.367
R541 B.n307 B.n27 163.367
R542 B.n303 B.n27 163.367
R543 B.n303 B.n302 163.367
R544 B.n302 B.n301 163.367
R545 B.n301 B.n29 163.367
R546 B.n296 B.n29 163.367
R547 B.n296 B.n295 163.367
R548 B.n295 B.n294 163.367
R549 B.n294 B.n33 163.367
R550 B.n290 B.n33 163.367
R551 B.n290 B.n289 163.367
R552 B.n289 B.n288 163.367
R553 B.n288 B.n35 163.367
R554 B.n284 B.n35 163.367
R555 B.n284 B.n283 163.367
R556 B.n283 B.n282 163.367
R557 B.n282 B.n37 163.367
R558 B.n278 B.n37 163.367
R559 B.n278 B.n277 163.367
R560 B.n277 B.n276 163.367
R561 B.n276 B.n39 163.367
R562 B.n272 B.n39 163.367
R563 B.n272 B.n271 163.367
R564 B.n74 B.n73 59.5399
R565 B.n160 B.n81 59.5399
R566 B.n24 B.n23 59.5399
R567 B.n298 B.n31 59.5399
R568 B.n73 B.n72 45.3823
R569 B.n81 B.n80 45.3823
R570 B.n23 B.n22 45.3823
R571 B.n31 B.n30 45.3823
R572 B.n341 B.n340 30.1273
R573 B.n269 B.n40 30.1273
R574 B.n203 B.n202 30.1273
R575 B.n131 B.n90 30.1273
R576 B B.n375 18.0485
R577 B.n340 B.n339 10.6151
R578 B.n339 B.n14 10.6151
R579 B.n335 B.n14 10.6151
R580 B.n335 B.n334 10.6151
R581 B.n334 B.n333 10.6151
R582 B.n333 B.n16 10.6151
R583 B.n329 B.n16 10.6151
R584 B.n329 B.n328 10.6151
R585 B.n328 B.n327 10.6151
R586 B.n327 B.n18 10.6151
R587 B.n323 B.n18 10.6151
R588 B.n323 B.n322 10.6151
R589 B.n322 B.n321 10.6151
R590 B.n321 B.n20 10.6151
R591 B.n317 B.n20 10.6151
R592 B.n317 B.n316 10.6151
R593 B.n316 B.n315 10.6151
R594 B.n312 B.n311 10.6151
R595 B.n311 B.n310 10.6151
R596 B.n310 B.n26 10.6151
R597 B.n306 B.n26 10.6151
R598 B.n306 B.n305 10.6151
R599 B.n305 B.n304 10.6151
R600 B.n304 B.n28 10.6151
R601 B.n300 B.n28 10.6151
R602 B.n300 B.n299 10.6151
R603 B.n297 B.n32 10.6151
R604 B.n293 B.n32 10.6151
R605 B.n293 B.n292 10.6151
R606 B.n292 B.n291 10.6151
R607 B.n291 B.n34 10.6151
R608 B.n287 B.n34 10.6151
R609 B.n287 B.n286 10.6151
R610 B.n286 B.n285 10.6151
R611 B.n285 B.n36 10.6151
R612 B.n281 B.n36 10.6151
R613 B.n281 B.n280 10.6151
R614 B.n280 B.n279 10.6151
R615 B.n279 B.n38 10.6151
R616 B.n275 B.n38 10.6151
R617 B.n275 B.n274 10.6151
R618 B.n274 B.n273 10.6151
R619 B.n273 B.n40 10.6151
R620 B.n203 B.n62 10.6151
R621 B.n207 B.n62 10.6151
R622 B.n208 B.n207 10.6151
R623 B.n209 B.n208 10.6151
R624 B.n209 B.n60 10.6151
R625 B.n213 B.n60 10.6151
R626 B.n214 B.n213 10.6151
R627 B.n215 B.n214 10.6151
R628 B.n215 B.n58 10.6151
R629 B.n219 B.n58 10.6151
R630 B.n220 B.n219 10.6151
R631 B.n221 B.n220 10.6151
R632 B.n221 B.n56 10.6151
R633 B.n225 B.n56 10.6151
R634 B.n226 B.n225 10.6151
R635 B.n227 B.n226 10.6151
R636 B.n227 B.n54 10.6151
R637 B.n231 B.n54 10.6151
R638 B.n232 B.n231 10.6151
R639 B.n233 B.n232 10.6151
R640 B.n233 B.n52 10.6151
R641 B.n237 B.n52 10.6151
R642 B.n238 B.n237 10.6151
R643 B.n239 B.n238 10.6151
R644 B.n239 B.n50 10.6151
R645 B.n243 B.n50 10.6151
R646 B.n244 B.n243 10.6151
R647 B.n245 B.n244 10.6151
R648 B.n245 B.n48 10.6151
R649 B.n249 B.n48 10.6151
R650 B.n250 B.n249 10.6151
R651 B.n251 B.n250 10.6151
R652 B.n251 B.n46 10.6151
R653 B.n255 B.n46 10.6151
R654 B.n256 B.n255 10.6151
R655 B.n257 B.n256 10.6151
R656 B.n257 B.n44 10.6151
R657 B.n261 B.n44 10.6151
R658 B.n262 B.n261 10.6151
R659 B.n263 B.n262 10.6151
R660 B.n263 B.n42 10.6151
R661 B.n267 B.n42 10.6151
R662 B.n268 B.n267 10.6151
R663 B.n269 B.n268 10.6151
R664 B.n135 B.n90 10.6151
R665 B.n136 B.n135 10.6151
R666 B.n137 B.n136 10.6151
R667 B.n137 B.n88 10.6151
R668 B.n141 B.n88 10.6151
R669 B.n142 B.n141 10.6151
R670 B.n143 B.n142 10.6151
R671 B.n143 B.n86 10.6151
R672 B.n147 B.n86 10.6151
R673 B.n148 B.n147 10.6151
R674 B.n149 B.n148 10.6151
R675 B.n149 B.n84 10.6151
R676 B.n153 B.n84 10.6151
R677 B.n154 B.n153 10.6151
R678 B.n155 B.n154 10.6151
R679 B.n155 B.n82 10.6151
R680 B.n159 B.n82 10.6151
R681 B.n162 B.n161 10.6151
R682 B.n162 B.n78 10.6151
R683 B.n166 B.n78 10.6151
R684 B.n167 B.n166 10.6151
R685 B.n168 B.n167 10.6151
R686 B.n168 B.n76 10.6151
R687 B.n172 B.n76 10.6151
R688 B.n173 B.n172 10.6151
R689 B.n174 B.n173 10.6151
R690 B.n178 B.n177 10.6151
R691 B.n179 B.n178 10.6151
R692 B.n179 B.n70 10.6151
R693 B.n183 B.n70 10.6151
R694 B.n184 B.n183 10.6151
R695 B.n185 B.n184 10.6151
R696 B.n185 B.n68 10.6151
R697 B.n189 B.n68 10.6151
R698 B.n190 B.n189 10.6151
R699 B.n191 B.n190 10.6151
R700 B.n191 B.n66 10.6151
R701 B.n195 B.n66 10.6151
R702 B.n196 B.n195 10.6151
R703 B.n197 B.n196 10.6151
R704 B.n197 B.n64 10.6151
R705 B.n201 B.n64 10.6151
R706 B.n202 B.n201 10.6151
R707 B.n131 B.n130 10.6151
R708 B.n130 B.n129 10.6151
R709 B.n129 B.n92 10.6151
R710 B.n125 B.n92 10.6151
R711 B.n125 B.n124 10.6151
R712 B.n124 B.n123 10.6151
R713 B.n123 B.n94 10.6151
R714 B.n119 B.n94 10.6151
R715 B.n119 B.n118 10.6151
R716 B.n118 B.n117 10.6151
R717 B.n117 B.n96 10.6151
R718 B.n113 B.n96 10.6151
R719 B.n113 B.n112 10.6151
R720 B.n112 B.n111 10.6151
R721 B.n111 B.n98 10.6151
R722 B.n107 B.n98 10.6151
R723 B.n107 B.n106 10.6151
R724 B.n106 B.n105 10.6151
R725 B.n105 B.n100 10.6151
R726 B.n101 B.n100 10.6151
R727 B.n101 B.n0 10.6151
R728 B.n371 B.n1 10.6151
R729 B.n371 B.n370 10.6151
R730 B.n370 B.n369 10.6151
R731 B.n369 B.n4 10.6151
R732 B.n365 B.n4 10.6151
R733 B.n365 B.n364 10.6151
R734 B.n364 B.n363 10.6151
R735 B.n363 B.n6 10.6151
R736 B.n359 B.n6 10.6151
R737 B.n359 B.n358 10.6151
R738 B.n358 B.n357 10.6151
R739 B.n357 B.n8 10.6151
R740 B.n353 B.n8 10.6151
R741 B.n353 B.n352 10.6151
R742 B.n352 B.n351 10.6151
R743 B.n351 B.n10 10.6151
R744 B.n347 B.n10 10.6151
R745 B.n347 B.n346 10.6151
R746 B.n346 B.n345 10.6151
R747 B.n345 B.n12 10.6151
R748 B.n341 B.n12 10.6151
R749 B.n315 B.n24 9.36635
R750 B.n298 B.n297 9.36635
R751 B.n160 B.n159 9.36635
R752 B.n177 B.n74 9.36635
R753 B.n375 B.n0 2.81026
R754 B.n375 B.n1 2.81026
R755 B.n312 B.n24 1.24928
R756 B.n299 B.n298 1.24928
R757 B.n161 B.n160 1.24928
R758 B.n174 B.n74 1.24928
R759 VN VN.t0 144.172
R760 VN VN.t1 107.183
R761 VDD2.n33 VDD2.n19 756.745
R762 VDD2.n14 VDD2.n0 756.745
R763 VDD2.n34 VDD2.n33 585
R764 VDD2.n32 VDD2.n31 585
R765 VDD2.n23 VDD2.n22 585
R766 VDD2.n26 VDD2.n25 585
R767 VDD2.n7 VDD2.n6 585
R768 VDD2.n4 VDD2.n3 585
R769 VDD2.n13 VDD2.n12 585
R770 VDD2.n15 VDD2.n14 585
R771 VDD2.t1 VDD2.n24 330.707
R772 VDD2.t0 VDD2.n5 330.707
R773 VDD2.n33 VDD2.n32 171.744
R774 VDD2.n32 VDD2.n22 171.744
R775 VDD2.n25 VDD2.n22 171.744
R776 VDD2.n6 VDD2.n3 171.744
R777 VDD2.n13 VDD2.n3 171.744
R778 VDD2.n14 VDD2.n13 171.744
R779 VDD2.n25 VDD2.t1 85.8723
R780 VDD2.n6 VDD2.t0 85.8723
R781 VDD2.n38 VDD2.n18 83.3119
R782 VDD2.n38 VDD2.n37 52.1611
R783 VDD2.n26 VDD2.n24 16.3201
R784 VDD2.n7 VDD2.n5 16.3201
R785 VDD2.n27 VDD2.n23 12.8005
R786 VDD2.n8 VDD2.n4 12.8005
R787 VDD2.n31 VDD2.n30 12.0247
R788 VDD2.n12 VDD2.n11 12.0247
R789 VDD2.n34 VDD2.n21 11.249
R790 VDD2.n15 VDD2.n2 11.249
R791 VDD2.n35 VDD2.n19 10.4732
R792 VDD2.n16 VDD2.n0 10.4732
R793 VDD2.n37 VDD2.n36 9.45567
R794 VDD2.n18 VDD2.n17 9.45567
R795 VDD2.n36 VDD2.n35 9.3005
R796 VDD2.n21 VDD2.n20 9.3005
R797 VDD2.n30 VDD2.n29 9.3005
R798 VDD2.n28 VDD2.n27 9.3005
R799 VDD2.n17 VDD2.n16 9.3005
R800 VDD2.n2 VDD2.n1 9.3005
R801 VDD2.n11 VDD2.n10 9.3005
R802 VDD2.n9 VDD2.n8 9.3005
R803 VDD2.n28 VDD2.n24 3.78097
R804 VDD2.n9 VDD2.n5 3.78097
R805 VDD2.n37 VDD2.n19 3.49141
R806 VDD2.n18 VDD2.n0 3.49141
R807 VDD2.n35 VDD2.n34 2.71565
R808 VDD2.n16 VDD2.n15 2.71565
R809 VDD2.n31 VDD2.n21 1.93989
R810 VDD2.n12 VDD2.n2 1.93989
R811 VDD2.n30 VDD2.n23 1.16414
R812 VDD2.n11 VDD2.n4 1.16414
R813 VDD2 VDD2.n38 0.563
R814 VDD2.n27 VDD2.n26 0.388379
R815 VDD2.n8 VDD2.n7 0.388379
R816 VDD2.n36 VDD2.n20 0.155672
R817 VDD2.n29 VDD2.n20 0.155672
R818 VDD2.n29 VDD2.n28 0.155672
R819 VDD2.n10 VDD2.n9 0.155672
R820 VDD2.n10 VDD2.n1 0.155672
R821 VDD2.n17 VDD2.n1 0.155672
C0 B VDD2 1.02776f
C1 VDD1 w_n1906_n1770# 1.15121f
C2 VN VP 3.70237f
C3 VTAIL VP 1.13814f
C4 VN VDD1 0.152088f
C5 B VP 1.24337f
C6 VTAIL VDD1 2.79961f
C7 VP VDD2 0.312162f
C8 B VDD1 1.00278f
C9 VN w_n1906_n1770# 2.41783f
C10 VDD1 VDD2 0.603344f
C11 VTAIL w_n1906_n1770# 1.58954f
C12 B w_n1906_n1770# 5.94068f
C13 w_n1906_n1770# VDD2 1.16966f
C14 VDD1 VP 1.21462f
C15 VN VTAIL 1.12396f
C16 VN B 0.848874f
C17 B VTAIL 1.66769f
C18 VN VDD2 1.05613f
C19 VP w_n1906_n1770# 2.65847f
C20 VTAIL VDD2 2.84786f
C21 VDD2 VSUBS 0.552677f
C22 VDD1 VSUBS 2.072798f
C23 VTAIL VSUBS 0.411594f
C24 VN VSUBS 4.98662f
C25 VP VSUBS 1.097004f
C26 B VSUBS 2.644245f
C27 w_n1906_n1770# VSUBS 42.4733f
C28 VDD2.n0 VSUBS 0.017028f
C29 VDD2.n1 VSUBS 0.015261f
C30 VDD2.n2 VSUBS 0.008201f
C31 VDD2.n3 VSUBS 0.019383f
C32 VDD2.n4 VSUBS 0.008683f
C33 VDD2.n5 VSUBS 0.059701f
C34 VDD2.t0 VSUBS 0.043131f
C35 VDD2.n6 VSUBS 0.014538f
C36 VDD2.n7 VSUBS 0.012192f
C37 VDD2.n8 VSUBS 0.008201f
C38 VDD2.n9 VSUBS 0.209544f
C39 VDD2.n10 VSUBS 0.015261f
C40 VDD2.n11 VSUBS 0.008201f
C41 VDD2.n12 VSUBS 0.008683f
C42 VDD2.n13 VSUBS 0.019383f
C43 VDD2.n14 VSUBS 0.047809f
C44 VDD2.n15 VSUBS 0.008683f
C45 VDD2.n16 VSUBS 0.008201f
C46 VDD2.n17 VSUBS 0.038819f
C47 VDD2.n18 VSUBS 0.26205f
C48 VDD2.n19 VSUBS 0.017028f
C49 VDD2.n20 VSUBS 0.015261f
C50 VDD2.n21 VSUBS 0.008201f
C51 VDD2.n22 VSUBS 0.019383f
C52 VDD2.n23 VSUBS 0.008683f
C53 VDD2.n24 VSUBS 0.059701f
C54 VDD2.t1 VSUBS 0.043131f
C55 VDD2.n25 VSUBS 0.014538f
C56 VDD2.n26 VSUBS 0.012192f
C57 VDD2.n27 VSUBS 0.008201f
C58 VDD2.n28 VSUBS 0.209544f
C59 VDD2.n29 VSUBS 0.015261f
C60 VDD2.n30 VSUBS 0.008201f
C61 VDD2.n31 VSUBS 0.008683f
C62 VDD2.n32 VSUBS 0.019383f
C63 VDD2.n33 VSUBS 0.047809f
C64 VDD2.n34 VSUBS 0.008683f
C65 VDD2.n35 VSUBS 0.008201f
C66 VDD2.n36 VSUBS 0.038819f
C67 VDD2.n37 VSUBS 0.034699f
C68 VDD2.n38 VSUBS 1.28376f
C69 VN.t1 VSUBS 1.21508f
C70 VN.t0 VSUBS 1.68055f
C71 B.n0 VSUBS 0.004504f
C72 B.n1 VSUBS 0.004504f
C73 B.n2 VSUBS 0.007122f
C74 B.n3 VSUBS 0.007122f
C75 B.n4 VSUBS 0.007122f
C76 B.n5 VSUBS 0.007122f
C77 B.n6 VSUBS 0.007122f
C78 B.n7 VSUBS 0.007122f
C79 B.n8 VSUBS 0.007122f
C80 B.n9 VSUBS 0.007122f
C81 B.n10 VSUBS 0.007122f
C82 B.n11 VSUBS 0.007122f
C83 B.n12 VSUBS 0.007122f
C84 B.n13 VSUBS 0.016227f
C85 B.n14 VSUBS 0.007122f
C86 B.n15 VSUBS 0.007122f
C87 B.n16 VSUBS 0.007122f
C88 B.n17 VSUBS 0.007122f
C89 B.n18 VSUBS 0.007122f
C90 B.n19 VSUBS 0.007122f
C91 B.n20 VSUBS 0.007122f
C92 B.n21 VSUBS 0.007122f
C93 B.t5 VSUBS 0.059276f
C94 B.t4 VSUBS 0.076236f
C95 B.t3 VSUBS 0.3905f
C96 B.n22 VSUBS 0.134722f
C97 B.n23 VSUBS 0.115252f
C98 B.n24 VSUBS 0.016501f
C99 B.n25 VSUBS 0.007122f
C100 B.n26 VSUBS 0.007122f
C101 B.n27 VSUBS 0.007122f
C102 B.n28 VSUBS 0.007122f
C103 B.n29 VSUBS 0.007122f
C104 B.t8 VSUBS 0.059277f
C105 B.t7 VSUBS 0.076237f
C106 B.t6 VSUBS 0.3905f
C107 B.n30 VSUBS 0.134721f
C108 B.n31 VSUBS 0.115251f
C109 B.n32 VSUBS 0.007122f
C110 B.n33 VSUBS 0.007122f
C111 B.n34 VSUBS 0.007122f
C112 B.n35 VSUBS 0.007122f
C113 B.n36 VSUBS 0.007122f
C114 B.n37 VSUBS 0.007122f
C115 B.n38 VSUBS 0.007122f
C116 B.n39 VSUBS 0.007122f
C117 B.n40 VSUBS 0.015315f
C118 B.n41 VSUBS 0.007122f
C119 B.n42 VSUBS 0.007122f
C120 B.n43 VSUBS 0.007122f
C121 B.n44 VSUBS 0.007122f
C122 B.n45 VSUBS 0.007122f
C123 B.n46 VSUBS 0.007122f
C124 B.n47 VSUBS 0.007122f
C125 B.n48 VSUBS 0.007122f
C126 B.n49 VSUBS 0.007122f
C127 B.n50 VSUBS 0.007122f
C128 B.n51 VSUBS 0.007122f
C129 B.n52 VSUBS 0.007122f
C130 B.n53 VSUBS 0.007122f
C131 B.n54 VSUBS 0.007122f
C132 B.n55 VSUBS 0.007122f
C133 B.n56 VSUBS 0.007122f
C134 B.n57 VSUBS 0.007122f
C135 B.n58 VSUBS 0.007122f
C136 B.n59 VSUBS 0.007122f
C137 B.n60 VSUBS 0.007122f
C138 B.n61 VSUBS 0.007122f
C139 B.n62 VSUBS 0.007122f
C140 B.n63 VSUBS 0.016227f
C141 B.n64 VSUBS 0.007122f
C142 B.n65 VSUBS 0.007122f
C143 B.n66 VSUBS 0.007122f
C144 B.n67 VSUBS 0.007122f
C145 B.n68 VSUBS 0.007122f
C146 B.n69 VSUBS 0.007122f
C147 B.n70 VSUBS 0.007122f
C148 B.n71 VSUBS 0.007122f
C149 B.t10 VSUBS 0.059277f
C150 B.t11 VSUBS 0.076237f
C151 B.t9 VSUBS 0.3905f
C152 B.n72 VSUBS 0.134721f
C153 B.n73 VSUBS 0.115251f
C154 B.n74 VSUBS 0.016501f
C155 B.n75 VSUBS 0.007122f
C156 B.n76 VSUBS 0.007122f
C157 B.n77 VSUBS 0.007122f
C158 B.n78 VSUBS 0.007122f
C159 B.n79 VSUBS 0.007122f
C160 B.t1 VSUBS 0.059276f
C161 B.t2 VSUBS 0.076236f
C162 B.t0 VSUBS 0.3905f
C163 B.n80 VSUBS 0.134722f
C164 B.n81 VSUBS 0.115252f
C165 B.n82 VSUBS 0.007122f
C166 B.n83 VSUBS 0.007122f
C167 B.n84 VSUBS 0.007122f
C168 B.n85 VSUBS 0.007122f
C169 B.n86 VSUBS 0.007122f
C170 B.n87 VSUBS 0.007122f
C171 B.n88 VSUBS 0.007122f
C172 B.n89 VSUBS 0.007122f
C173 B.n90 VSUBS 0.016227f
C174 B.n91 VSUBS 0.007122f
C175 B.n92 VSUBS 0.007122f
C176 B.n93 VSUBS 0.007122f
C177 B.n94 VSUBS 0.007122f
C178 B.n95 VSUBS 0.007122f
C179 B.n96 VSUBS 0.007122f
C180 B.n97 VSUBS 0.007122f
C181 B.n98 VSUBS 0.007122f
C182 B.n99 VSUBS 0.007122f
C183 B.n100 VSUBS 0.007122f
C184 B.n101 VSUBS 0.007122f
C185 B.n102 VSUBS 0.007122f
C186 B.n103 VSUBS 0.007122f
C187 B.n104 VSUBS 0.007122f
C188 B.n105 VSUBS 0.007122f
C189 B.n106 VSUBS 0.007122f
C190 B.n107 VSUBS 0.007122f
C191 B.n108 VSUBS 0.007122f
C192 B.n109 VSUBS 0.007122f
C193 B.n110 VSUBS 0.007122f
C194 B.n111 VSUBS 0.007122f
C195 B.n112 VSUBS 0.007122f
C196 B.n113 VSUBS 0.007122f
C197 B.n114 VSUBS 0.007122f
C198 B.n115 VSUBS 0.007122f
C199 B.n116 VSUBS 0.007122f
C200 B.n117 VSUBS 0.007122f
C201 B.n118 VSUBS 0.007122f
C202 B.n119 VSUBS 0.007122f
C203 B.n120 VSUBS 0.007122f
C204 B.n121 VSUBS 0.007122f
C205 B.n122 VSUBS 0.007122f
C206 B.n123 VSUBS 0.007122f
C207 B.n124 VSUBS 0.007122f
C208 B.n125 VSUBS 0.007122f
C209 B.n126 VSUBS 0.007122f
C210 B.n127 VSUBS 0.007122f
C211 B.n128 VSUBS 0.007122f
C212 B.n129 VSUBS 0.007122f
C213 B.n130 VSUBS 0.007122f
C214 B.n131 VSUBS 0.015404f
C215 B.n132 VSUBS 0.015404f
C216 B.n133 VSUBS 0.016227f
C217 B.n134 VSUBS 0.007122f
C218 B.n135 VSUBS 0.007122f
C219 B.n136 VSUBS 0.007122f
C220 B.n137 VSUBS 0.007122f
C221 B.n138 VSUBS 0.007122f
C222 B.n139 VSUBS 0.007122f
C223 B.n140 VSUBS 0.007122f
C224 B.n141 VSUBS 0.007122f
C225 B.n142 VSUBS 0.007122f
C226 B.n143 VSUBS 0.007122f
C227 B.n144 VSUBS 0.007122f
C228 B.n145 VSUBS 0.007122f
C229 B.n146 VSUBS 0.007122f
C230 B.n147 VSUBS 0.007122f
C231 B.n148 VSUBS 0.007122f
C232 B.n149 VSUBS 0.007122f
C233 B.n150 VSUBS 0.007122f
C234 B.n151 VSUBS 0.007122f
C235 B.n152 VSUBS 0.007122f
C236 B.n153 VSUBS 0.007122f
C237 B.n154 VSUBS 0.007122f
C238 B.n155 VSUBS 0.007122f
C239 B.n156 VSUBS 0.007122f
C240 B.n157 VSUBS 0.007122f
C241 B.n158 VSUBS 0.007122f
C242 B.n159 VSUBS 0.006703f
C243 B.n160 VSUBS 0.016501f
C244 B.n161 VSUBS 0.00398f
C245 B.n162 VSUBS 0.007122f
C246 B.n163 VSUBS 0.007122f
C247 B.n164 VSUBS 0.007122f
C248 B.n165 VSUBS 0.007122f
C249 B.n166 VSUBS 0.007122f
C250 B.n167 VSUBS 0.007122f
C251 B.n168 VSUBS 0.007122f
C252 B.n169 VSUBS 0.007122f
C253 B.n170 VSUBS 0.007122f
C254 B.n171 VSUBS 0.007122f
C255 B.n172 VSUBS 0.007122f
C256 B.n173 VSUBS 0.007122f
C257 B.n174 VSUBS 0.00398f
C258 B.n175 VSUBS 0.007122f
C259 B.n176 VSUBS 0.007122f
C260 B.n177 VSUBS 0.006703f
C261 B.n178 VSUBS 0.007122f
C262 B.n179 VSUBS 0.007122f
C263 B.n180 VSUBS 0.007122f
C264 B.n181 VSUBS 0.007122f
C265 B.n182 VSUBS 0.007122f
C266 B.n183 VSUBS 0.007122f
C267 B.n184 VSUBS 0.007122f
C268 B.n185 VSUBS 0.007122f
C269 B.n186 VSUBS 0.007122f
C270 B.n187 VSUBS 0.007122f
C271 B.n188 VSUBS 0.007122f
C272 B.n189 VSUBS 0.007122f
C273 B.n190 VSUBS 0.007122f
C274 B.n191 VSUBS 0.007122f
C275 B.n192 VSUBS 0.007122f
C276 B.n193 VSUBS 0.007122f
C277 B.n194 VSUBS 0.007122f
C278 B.n195 VSUBS 0.007122f
C279 B.n196 VSUBS 0.007122f
C280 B.n197 VSUBS 0.007122f
C281 B.n198 VSUBS 0.007122f
C282 B.n199 VSUBS 0.007122f
C283 B.n200 VSUBS 0.007122f
C284 B.n201 VSUBS 0.007122f
C285 B.n202 VSUBS 0.016227f
C286 B.n203 VSUBS 0.015404f
C287 B.n204 VSUBS 0.015404f
C288 B.n205 VSUBS 0.007122f
C289 B.n206 VSUBS 0.007122f
C290 B.n207 VSUBS 0.007122f
C291 B.n208 VSUBS 0.007122f
C292 B.n209 VSUBS 0.007122f
C293 B.n210 VSUBS 0.007122f
C294 B.n211 VSUBS 0.007122f
C295 B.n212 VSUBS 0.007122f
C296 B.n213 VSUBS 0.007122f
C297 B.n214 VSUBS 0.007122f
C298 B.n215 VSUBS 0.007122f
C299 B.n216 VSUBS 0.007122f
C300 B.n217 VSUBS 0.007122f
C301 B.n218 VSUBS 0.007122f
C302 B.n219 VSUBS 0.007122f
C303 B.n220 VSUBS 0.007122f
C304 B.n221 VSUBS 0.007122f
C305 B.n222 VSUBS 0.007122f
C306 B.n223 VSUBS 0.007122f
C307 B.n224 VSUBS 0.007122f
C308 B.n225 VSUBS 0.007122f
C309 B.n226 VSUBS 0.007122f
C310 B.n227 VSUBS 0.007122f
C311 B.n228 VSUBS 0.007122f
C312 B.n229 VSUBS 0.007122f
C313 B.n230 VSUBS 0.007122f
C314 B.n231 VSUBS 0.007122f
C315 B.n232 VSUBS 0.007122f
C316 B.n233 VSUBS 0.007122f
C317 B.n234 VSUBS 0.007122f
C318 B.n235 VSUBS 0.007122f
C319 B.n236 VSUBS 0.007122f
C320 B.n237 VSUBS 0.007122f
C321 B.n238 VSUBS 0.007122f
C322 B.n239 VSUBS 0.007122f
C323 B.n240 VSUBS 0.007122f
C324 B.n241 VSUBS 0.007122f
C325 B.n242 VSUBS 0.007122f
C326 B.n243 VSUBS 0.007122f
C327 B.n244 VSUBS 0.007122f
C328 B.n245 VSUBS 0.007122f
C329 B.n246 VSUBS 0.007122f
C330 B.n247 VSUBS 0.007122f
C331 B.n248 VSUBS 0.007122f
C332 B.n249 VSUBS 0.007122f
C333 B.n250 VSUBS 0.007122f
C334 B.n251 VSUBS 0.007122f
C335 B.n252 VSUBS 0.007122f
C336 B.n253 VSUBS 0.007122f
C337 B.n254 VSUBS 0.007122f
C338 B.n255 VSUBS 0.007122f
C339 B.n256 VSUBS 0.007122f
C340 B.n257 VSUBS 0.007122f
C341 B.n258 VSUBS 0.007122f
C342 B.n259 VSUBS 0.007122f
C343 B.n260 VSUBS 0.007122f
C344 B.n261 VSUBS 0.007122f
C345 B.n262 VSUBS 0.007122f
C346 B.n263 VSUBS 0.007122f
C347 B.n264 VSUBS 0.007122f
C348 B.n265 VSUBS 0.007122f
C349 B.n266 VSUBS 0.007122f
C350 B.n267 VSUBS 0.007122f
C351 B.n268 VSUBS 0.007122f
C352 B.n269 VSUBS 0.016316f
C353 B.n270 VSUBS 0.015404f
C354 B.n271 VSUBS 0.016227f
C355 B.n272 VSUBS 0.007122f
C356 B.n273 VSUBS 0.007122f
C357 B.n274 VSUBS 0.007122f
C358 B.n275 VSUBS 0.007122f
C359 B.n276 VSUBS 0.007122f
C360 B.n277 VSUBS 0.007122f
C361 B.n278 VSUBS 0.007122f
C362 B.n279 VSUBS 0.007122f
C363 B.n280 VSUBS 0.007122f
C364 B.n281 VSUBS 0.007122f
C365 B.n282 VSUBS 0.007122f
C366 B.n283 VSUBS 0.007122f
C367 B.n284 VSUBS 0.007122f
C368 B.n285 VSUBS 0.007122f
C369 B.n286 VSUBS 0.007122f
C370 B.n287 VSUBS 0.007122f
C371 B.n288 VSUBS 0.007122f
C372 B.n289 VSUBS 0.007122f
C373 B.n290 VSUBS 0.007122f
C374 B.n291 VSUBS 0.007122f
C375 B.n292 VSUBS 0.007122f
C376 B.n293 VSUBS 0.007122f
C377 B.n294 VSUBS 0.007122f
C378 B.n295 VSUBS 0.007122f
C379 B.n296 VSUBS 0.007122f
C380 B.n297 VSUBS 0.006703f
C381 B.n298 VSUBS 0.016501f
C382 B.n299 VSUBS 0.00398f
C383 B.n300 VSUBS 0.007122f
C384 B.n301 VSUBS 0.007122f
C385 B.n302 VSUBS 0.007122f
C386 B.n303 VSUBS 0.007122f
C387 B.n304 VSUBS 0.007122f
C388 B.n305 VSUBS 0.007122f
C389 B.n306 VSUBS 0.007122f
C390 B.n307 VSUBS 0.007122f
C391 B.n308 VSUBS 0.007122f
C392 B.n309 VSUBS 0.007122f
C393 B.n310 VSUBS 0.007122f
C394 B.n311 VSUBS 0.007122f
C395 B.n312 VSUBS 0.00398f
C396 B.n313 VSUBS 0.007122f
C397 B.n314 VSUBS 0.007122f
C398 B.n315 VSUBS 0.006703f
C399 B.n316 VSUBS 0.007122f
C400 B.n317 VSUBS 0.007122f
C401 B.n318 VSUBS 0.007122f
C402 B.n319 VSUBS 0.007122f
C403 B.n320 VSUBS 0.007122f
C404 B.n321 VSUBS 0.007122f
C405 B.n322 VSUBS 0.007122f
C406 B.n323 VSUBS 0.007122f
C407 B.n324 VSUBS 0.007122f
C408 B.n325 VSUBS 0.007122f
C409 B.n326 VSUBS 0.007122f
C410 B.n327 VSUBS 0.007122f
C411 B.n328 VSUBS 0.007122f
C412 B.n329 VSUBS 0.007122f
C413 B.n330 VSUBS 0.007122f
C414 B.n331 VSUBS 0.007122f
C415 B.n332 VSUBS 0.007122f
C416 B.n333 VSUBS 0.007122f
C417 B.n334 VSUBS 0.007122f
C418 B.n335 VSUBS 0.007122f
C419 B.n336 VSUBS 0.007122f
C420 B.n337 VSUBS 0.007122f
C421 B.n338 VSUBS 0.007122f
C422 B.n339 VSUBS 0.007122f
C423 B.n340 VSUBS 0.016227f
C424 B.n341 VSUBS 0.015404f
C425 B.n342 VSUBS 0.015404f
C426 B.n343 VSUBS 0.007122f
C427 B.n344 VSUBS 0.007122f
C428 B.n345 VSUBS 0.007122f
C429 B.n346 VSUBS 0.007122f
C430 B.n347 VSUBS 0.007122f
C431 B.n348 VSUBS 0.007122f
C432 B.n349 VSUBS 0.007122f
C433 B.n350 VSUBS 0.007122f
C434 B.n351 VSUBS 0.007122f
C435 B.n352 VSUBS 0.007122f
C436 B.n353 VSUBS 0.007122f
C437 B.n354 VSUBS 0.007122f
C438 B.n355 VSUBS 0.007122f
C439 B.n356 VSUBS 0.007122f
C440 B.n357 VSUBS 0.007122f
C441 B.n358 VSUBS 0.007122f
C442 B.n359 VSUBS 0.007122f
C443 B.n360 VSUBS 0.007122f
C444 B.n361 VSUBS 0.007122f
C445 B.n362 VSUBS 0.007122f
C446 B.n363 VSUBS 0.007122f
C447 B.n364 VSUBS 0.007122f
C448 B.n365 VSUBS 0.007122f
C449 B.n366 VSUBS 0.007122f
C450 B.n367 VSUBS 0.007122f
C451 B.n368 VSUBS 0.007122f
C452 B.n369 VSUBS 0.007122f
C453 B.n370 VSUBS 0.007122f
C454 B.n371 VSUBS 0.007122f
C455 B.n372 VSUBS 0.007122f
C456 B.n373 VSUBS 0.007122f
C457 B.n374 VSUBS 0.007122f
C458 B.n375 VSUBS 0.016127f
C459 VDD1.n0 VSUBS 0.016692f
C460 VDD1.n1 VSUBS 0.01496f
C461 VDD1.n2 VSUBS 0.008039f
C462 VDD1.n3 VSUBS 0.019001f
C463 VDD1.n4 VSUBS 0.008512f
C464 VDD1.n5 VSUBS 0.058523f
C465 VDD1.t0 VSUBS 0.04228f
C466 VDD1.n6 VSUBS 0.014251f
C467 VDD1.n7 VSUBS 0.011951f
C468 VDD1.n8 VSUBS 0.008039f
C469 VDD1.n9 VSUBS 0.205409f
C470 VDD1.n10 VSUBS 0.01496f
C471 VDD1.n11 VSUBS 0.008039f
C472 VDD1.n12 VSUBS 0.008512f
C473 VDD1.n13 VSUBS 0.019001f
C474 VDD1.n14 VSUBS 0.046866f
C475 VDD1.n15 VSUBS 0.008512f
C476 VDD1.n16 VSUBS 0.008039f
C477 VDD1.n17 VSUBS 0.038053f
C478 VDD1.n18 VSUBS 0.034632f
C479 VDD1.n19 VSUBS 0.016692f
C480 VDD1.n20 VSUBS 0.01496f
C481 VDD1.n21 VSUBS 0.008039f
C482 VDD1.n22 VSUBS 0.019001f
C483 VDD1.n23 VSUBS 0.008512f
C484 VDD1.n24 VSUBS 0.058523f
C485 VDD1.t1 VSUBS 0.04228f
C486 VDD1.n25 VSUBS 0.014251f
C487 VDD1.n26 VSUBS 0.011951f
C488 VDD1.n27 VSUBS 0.008039f
C489 VDD1.n28 VSUBS 0.205409f
C490 VDD1.n29 VSUBS 0.01496f
C491 VDD1.n30 VSUBS 0.008039f
C492 VDD1.n31 VSUBS 0.008512f
C493 VDD1.n32 VSUBS 0.019001f
C494 VDD1.n33 VSUBS 0.046866f
C495 VDD1.n34 VSUBS 0.008512f
C496 VDD1.n35 VSUBS 0.008039f
C497 VDD1.n36 VSUBS 0.038053f
C498 VDD1.n37 VSUBS 0.27826f
C499 VTAIL.n0 VSUBS 0.01972f
C500 VTAIL.n1 VSUBS 0.017673f
C501 VTAIL.n2 VSUBS 0.009497f
C502 VTAIL.n3 VSUBS 0.022447f
C503 VTAIL.n4 VSUBS 0.010055f
C504 VTAIL.n5 VSUBS 0.069137f
C505 VTAIL.t3 VSUBS 0.049948f
C506 VTAIL.n6 VSUBS 0.016835f
C507 VTAIL.n7 VSUBS 0.014119f
C508 VTAIL.n8 VSUBS 0.009497f
C509 VTAIL.n9 VSUBS 0.242664f
C510 VTAIL.n10 VSUBS 0.017673f
C511 VTAIL.n11 VSUBS 0.009497f
C512 VTAIL.n12 VSUBS 0.010055f
C513 VTAIL.n13 VSUBS 0.022447f
C514 VTAIL.n14 VSUBS 0.055366f
C515 VTAIL.n15 VSUBS 0.010055f
C516 VTAIL.n16 VSUBS 0.009497f
C517 VTAIL.n17 VSUBS 0.044955f
C518 VTAIL.n18 VSUBS 0.028009f
C519 VTAIL.n19 VSUBS 0.742885f
C520 VTAIL.n20 VSUBS 0.01972f
C521 VTAIL.n21 VSUBS 0.017673f
C522 VTAIL.n22 VSUBS 0.009497f
C523 VTAIL.n23 VSUBS 0.022447f
C524 VTAIL.n24 VSUBS 0.010055f
C525 VTAIL.n25 VSUBS 0.069137f
C526 VTAIL.t1 VSUBS 0.049948f
C527 VTAIL.n26 VSUBS 0.016835f
C528 VTAIL.n27 VSUBS 0.014119f
C529 VTAIL.n28 VSUBS 0.009497f
C530 VTAIL.n29 VSUBS 0.242664f
C531 VTAIL.n30 VSUBS 0.017673f
C532 VTAIL.n31 VSUBS 0.009497f
C533 VTAIL.n32 VSUBS 0.010055f
C534 VTAIL.n33 VSUBS 0.022447f
C535 VTAIL.n34 VSUBS 0.055366f
C536 VTAIL.n35 VSUBS 0.010055f
C537 VTAIL.n36 VSUBS 0.009497f
C538 VTAIL.n37 VSUBS 0.044955f
C539 VTAIL.n38 VSUBS 0.028009f
C540 VTAIL.n39 VSUBS 0.76829f
C541 VTAIL.n40 VSUBS 0.01972f
C542 VTAIL.n41 VSUBS 0.017673f
C543 VTAIL.n42 VSUBS 0.009497f
C544 VTAIL.n43 VSUBS 0.022447f
C545 VTAIL.n44 VSUBS 0.010055f
C546 VTAIL.n45 VSUBS 0.069137f
C547 VTAIL.t2 VSUBS 0.049948f
C548 VTAIL.n46 VSUBS 0.016835f
C549 VTAIL.n47 VSUBS 0.014119f
C550 VTAIL.n48 VSUBS 0.009497f
C551 VTAIL.n49 VSUBS 0.242664f
C552 VTAIL.n50 VSUBS 0.017673f
C553 VTAIL.n51 VSUBS 0.009497f
C554 VTAIL.n52 VSUBS 0.010055f
C555 VTAIL.n53 VSUBS 0.022447f
C556 VTAIL.n54 VSUBS 0.055366f
C557 VTAIL.n55 VSUBS 0.010055f
C558 VTAIL.n56 VSUBS 0.009497f
C559 VTAIL.n57 VSUBS 0.044955f
C560 VTAIL.n58 VSUBS 0.028009f
C561 VTAIL.n59 VSUBS 0.653414f
C562 VTAIL.n60 VSUBS 0.01972f
C563 VTAIL.n61 VSUBS 0.017673f
C564 VTAIL.n62 VSUBS 0.009497f
C565 VTAIL.n63 VSUBS 0.022447f
C566 VTAIL.n64 VSUBS 0.010055f
C567 VTAIL.n65 VSUBS 0.069137f
C568 VTAIL.t0 VSUBS 0.049948f
C569 VTAIL.n66 VSUBS 0.016835f
C570 VTAIL.n67 VSUBS 0.014119f
C571 VTAIL.n68 VSUBS 0.009497f
C572 VTAIL.n69 VSUBS 0.242664f
C573 VTAIL.n70 VSUBS 0.017673f
C574 VTAIL.n71 VSUBS 0.009497f
C575 VTAIL.n72 VSUBS 0.010055f
C576 VTAIL.n73 VSUBS 0.022447f
C577 VTAIL.n74 VSUBS 0.055366f
C578 VTAIL.n75 VSUBS 0.010055f
C579 VTAIL.n76 VSUBS 0.009497f
C580 VTAIL.n77 VSUBS 0.044955f
C581 VTAIL.n78 VSUBS 0.028009f
C582 VTAIL.n79 VSUBS 0.594626f
C583 VP.t1 VSUBS 1.77316f
C584 VP.t0 VSUBS 1.28653f
C585 VP.n0 VSUBS 3.26409f
.ends

