* NGSPICE file created from diff_pair_sample_0119.ext - technology: sky130A

.subckt diff_pair_sample_0119 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=1.2903 ps=8.15 w=7.82 l=0.66
X1 B.t11 B.t9 B.t10 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=0 ps=0 w=7.82 l=0.66
X2 B.t8 B.t6 B.t7 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=0 ps=0 w=7.82 l=0.66
X3 B.t5 B.t3 B.t4 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=0 ps=0 w=7.82 l=0.66
X4 VTAIL.t2 VN.t0 VDD2.t5 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=1.2903 ps=8.15 w=7.82 l=0.66
X5 VTAIL.t10 VP.t1 VDD1.t4 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=1.2903 ps=8.15 w=7.82 l=0.66
X6 B.t2 B.t0 B.t1 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=0 ps=0 w=7.82 l=0.66
X7 VDD2.t4 VN.t1 VTAIL.t1 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=3.0498 ps=16.42 w=7.82 l=0.66
X8 VTAIL.t0 VN.t2 VDD2.t3 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=1.2903 ps=8.15 w=7.82 l=0.66
X9 VDD2.t2 VN.t3 VTAIL.t5 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=1.2903 ps=8.15 w=7.82 l=0.66
X10 VDD1.t3 VP.t2 VTAIL.t7 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=1.2903 ps=8.15 w=7.82 l=0.66
X11 VTAIL.t8 VP.t3 VDD1.t2 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=1.2903 ps=8.15 w=7.82 l=0.66
X12 VDD1.t1 VP.t4 VTAIL.t6 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=3.0498 ps=16.42 w=7.82 l=0.66
X13 VDD2.t1 VN.t4 VTAIL.t4 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=3.0498 pd=16.42 as=1.2903 ps=8.15 w=7.82 l=0.66
X14 VDD2.t0 VN.t5 VTAIL.t3 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=3.0498 ps=16.42 w=7.82 l=0.66
X15 VDD1.t0 VP.t5 VTAIL.t11 w_n1762_n2532# sky130_fd_pr__pfet_01v8 ad=1.2903 pd=8.15 as=3.0498 ps=16.42 w=7.82 l=0.66
R0 VP.n3 VP.t2 366.592
R1 VP.n8 VP.t0 345.798
R2 VP.n12 VP.t1 345.798
R3 VP.n14 VP.t5 345.798
R4 VP.n6 VP.t4 345.798
R5 VP.n4 VP.t3 345.798
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.8515
R14 VP.n9 VP.n7 37.8376
R15 VP.n12 VP.n1 24.8308
R16 VP.n13 VP.n12 24.8308
R17 VP.n5 VP.n4 24.8308
R18 VP.n8 VP.n1 23.3702
R19 VP.n14 VP.n13 23.3702
R20 VP.n6 VP.n5 23.3702
R21 VP.n4 VP.n3 21.148
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VTAIL.n170 VTAIL.n134 756.745
R29 VTAIL.n38 VTAIL.n2 756.745
R30 VTAIL.n128 VTAIL.n92 756.745
R31 VTAIL.n84 VTAIL.n48 756.745
R32 VTAIL.n146 VTAIL.n145 585
R33 VTAIL.n151 VTAIL.n150 585
R34 VTAIL.n153 VTAIL.n152 585
R35 VTAIL.n142 VTAIL.n141 585
R36 VTAIL.n159 VTAIL.n158 585
R37 VTAIL.n161 VTAIL.n160 585
R38 VTAIL.n138 VTAIL.n137 585
R39 VTAIL.n168 VTAIL.n167 585
R40 VTAIL.n169 VTAIL.n136 585
R41 VTAIL.n171 VTAIL.n170 585
R42 VTAIL.n14 VTAIL.n13 585
R43 VTAIL.n19 VTAIL.n18 585
R44 VTAIL.n21 VTAIL.n20 585
R45 VTAIL.n10 VTAIL.n9 585
R46 VTAIL.n27 VTAIL.n26 585
R47 VTAIL.n29 VTAIL.n28 585
R48 VTAIL.n6 VTAIL.n5 585
R49 VTAIL.n36 VTAIL.n35 585
R50 VTAIL.n37 VTAIL.n4 585
R51 VTAIL.n39 VTAIL.n38 585
R52 VTAIL.n129 VTAIL.n128 585
R53 VTAIL.n127 VTAIL.n94 585
R54 VTAIL.n126 VTAIL.n125 585
R55 VTAIL.n97 VTAIL.n95 585
R56 VTAIL.n120 VTAIL.n119 585
R57 VTAIL.n118 VTAIL.n117 585
R58 VTAIL.n101 VTAIL.n100 585
R59 VTAIL.n112 VTAIL.n111 585
R60 VTAIL.n110 VTAIL.n109 585
R61 VTAIL.n105 VTAIL.n104 585
R62 VTAIL.n85 VTAIL.n84 585
R63 VTAIL.n83 VTAIL.n50 585
R64 VTAIL.n82 VTAIL.n81 585
R65 VTAIL.n53 VTAIL.n51 585
R66 VTAIL.n76 VTAIL.n75 585
R67 VTAIL.n74 VTAIL.n73 585
R68 VTAIL.n57 VTAIL.n56 585
R69 VTAIL.n68 VTAIL.n67 585
R70 VTAIL.n66 VTAIL.n65 585
R71 VTAIL.n61 VTAIL.n60 585
R72 VTAIL.n147 VTAIL.t3 329.043
R73 VTAIL.n15 VTAIL.t11 329.043
R74 VTAIL.n106 VTAIL.t6 329.043
R75 VTAIL.n62 VTAIL.t1 329.043
R76 VTAIL.n151 VTAIL.n145 171.744
R77 VTAIL.n152 VTAIL.n151 171.744
R78 VTAIL.n152 VTAIL.n141 171.744
R79 VTAIL.n159 VTAIL.n141 171.744
R80 VTAIL.n160 VTAIL.n159 171.744
R81 VTAIL.n160 VTAIL.n137 171.744
R82 VTAIL.n168 VTAIL.n137 171.744
R83 VTAIL.n169 VTAIL.n168 171.744
R84 VTAIL.n170 VTAIL.n169 171.744
R85 VTAIL.n19 VTAIL.n13 171.744
R86 VTAIL.n20 VTAIL.n19 171.744
R87 VTAIL.n20 VTAIL.n9 171.744
R88 VTAIL.n27 VTAIL.n9 171.744
R89 VTAIL.n28 VTAIL.n27 171.744
R90 VTAIL.n28 VTAIL.n5 171.744
R91 VTAIL.n36 VTAIL.n5 171.744
R92 VTAIL.n37 VTAIL.n36 171.744
R93 VTAIL.n38 VTAIL.n37 171.744
R94 VTAIL.n128 VTAIL.n127 171.744
R95 VTAIL.n127 VTAIL.n126 171.744
R96 VTAIL.n126 VTAIL.n95 171.744
R97 VTAIL.n119 VTAIL.n95 171.744
R98 VTAIL.n119 VTAIL.n118 171.744
R99 VTAIL.n118 VTAIL.n100 171.744
R100 VTAIL.n111 VTAIL.n100 171.744
R101 VTAIL.n111 VTAIL.n110 171.744
R102 VTAIL.n110 VTAIL.n104 171.744
R103 VTAIL.n84 VTAIL.n83 171.744
R104 VTAIL.n83 VTAIL.n82 171.744
R105 VTAIL.n82 VTAIL.n51 171.744
R106 VTAIL.n75 VTAIL.n51 171.744
R107 VTAIL.n75 VTAIL.n74 171.744
R108 VTAIL.n74 VTAIL.n56 171.744
R109 VTAIL.n67 VTAIL.n56 171.744
R110 VTAIL.n67 VTAIL.n66 171.744
R111 VTAIL.n66 VTAIL.n60 171.744
R112 VTAIL.t3 VTAIL.n145 85.8723
R113 VTAIL.t11 VTAIL.n13 85.8723
R114 VTAIL.t6 VTAIL.n104 85.8723
R115 VTAIL.t1 VTAIL.n60 85.8723
R116 VTAIL.n91 VTAIL.n90 66.0683
R117 VTAIL.n47 VTAIL.n46 66.0683
R118 VTAIL.n1 VTAIL.n0 66.0682
R119 VTAIL.n45 VTAIL.n44 66.0682
R120 VTAIL.n175 VTAIL.n174 32.5732
R121 VTAIL.n43 VTAIL.n42 32.5732
R122 VTAIL.n133 VTAIL.n132 32.5732
R123 VTAIL.n89 VTAIL.n88 32.5732
R124 VTAIL.n47 VTAIL.n45 20.8152
R125 VTAIL.n175 VTAIL.n133 19.9617
R126 VTAIL.n171 VTAIL.n136 13.1884
R127 VTAIL.n39 VTAIL.n4 13.1884
R128 VTAIL.n129 VTAIL.n94 13.1884
R129 VTAIL.n85 VTAIL.n50 13.1884
R130 VTAIL.n167 VTAIL.n166 12.8005
R131 VTAIL.n172 VTAIL.n134 12.8005
R132 VTAIL.n35 VTAIL.n34 12.8005
R133 VTAIL.n40 VTAIL.n2 12.8005
R134 VTAIL.n130 VTAIL.n92 12.8005
R135 VTAIL.n125 VTAIL.n96 12.8005
R136 VTAIL.n86 VTAIL.n48 12.8005
R137 VTAIL.n81 VTAIL.n52 12.8005
R138 VTAIL.n165 VTAIL.n138 12.0247
R139 VTAIL.n33 VTAIL.n6 12.0247
R140 VTAIL.n124 VTAIL.n97 12.0247
R141 VTAIL.n80 VTAIL.n53 12.0247
R142 VTAIL.n162 VTAIL.n161 11.249
R143 VTAIL.n30 VTAIL.n29 11.249
R144 VTAIL.n121 VTAIL.n120 11.249
R145 VTAIL.n77 VTAIL.n76 11.249
R146 VTAIL.n147 VTAIL.n146 10.7238
R147 VTAIL.n15 VTAIL.n14 10.7238
R148 VTAIL.n106 VTAIL.n105 10.7238
R149 VTAIL.n62 VTAIL.n61 10.7238
R150 VTAIL.n158 VTAIL.n140 10.4732
R151 VTAIL.n26 VTAIL.n8 10.4732
R152 VTAIL.n117 VTAIL.n99 10.4732
R153 VTAIL.n73 VTAIL.n55 10.4732
R154 VTAIL.n157 VTAIL.n142 9.69747
R155 VTAIL.n25 VTAIL.n10 9.69747
R156 VTAIL.n116 VTAIL.n101 9.69747
R157 VTAIL.n72 VTAIL.n57 9.69747
R158 VTAIL.n174 VTAIL.n173 9.45567
R159 VTAIL.n42 VTAIL.n41 9.45567
R160 VTAIL.n132 VTAIL.n131 9.45567
R161 VTAIL.n88 VTAIL.n87 9.45567
R162 VTAIL.n173 VTAIL.n172 9.3005
R163 VTAIL.n149 VTAIL.n148 9.3005
R164 VTAIL.n144 VTAIL.n143 9.3005
R165 VTAIL.n155 VTAIL.n154 9.3005
R166 VTAIL.n157 VTAIL.n156 9.3005
R167 VTAIL.n140 VTAIL.n139 9.3005
R168 VTAIL.n163 VTAIL.n162 9.3005
R169 VTAIL.n165 VTAIL.n164 9.3005
R170 VTAIL.n166 VTAIL.n135 9.3005
R171 VTAIL.n41 VTAIL.n40 9.3005
R172 VTAIL.n17 VTAIL.n16 9.3005
R173 VTAIL.n12 VTAIL.n11 9.3005
R174 VTAIL.n23 VTAIL.n22 9.3005
R175 VTAIL.n25 VTAIL.n24 9.3005
R176 VTAIL.n8 VTAIL.n7 9.3005
R177 VTAIL.n31 VTAIL.n30 9.3005
R178 VTAIL.n33 VTAIL.n32 9.3005
R179 VTAIL.n34 VTAIL.n3 9.3005
R180 VTAIL.n108 VTAIL.n107 9.3005
R181 VTAIL.n103 VTAIL.n102 9.3005
R182 VTAIL.n114 VTAIL.n113 9.3005
R183 VTAIL.n116 VTAIL.n115 9.3005
R184 VTAIL.n99 VTAIL.n98 9.3005
R185 VTAIL.n122 VTAIL.n121 9.3005
R186 VTAIL.n124 VTAIL.n123 9.3005
R187 VTAIL.n96 VTAIL.n93 9.3005
R188 VTAIL.n131 VTAIL.n130 9.3005
R189 VTAIL.n64 VTAIL.n63 9.3005
R190 VTAIL.n59 VTAIL.n58 9.3005
R191 VTAIL.n70 VTAIL.n69 9.3005
R192 VTAIL.n72 VTAIL.n71 9.3005
R193 VTAIL.n55 VTAIL.n54 9.3005
R194 VTAIL.n78 VTAIL.n77 9.3005
R195 VTAIL.n80 VTAIL.n79 9.3005
R196 VTAIL.n52 VTAIL.n49 9.3005
R197 VTAIL.n87 VTAIL.n86 9.3005
R198 VTAIL.n154 VTAIL.n153 8.92171
R199 VTAIL.n22 VTAIL.n21 8.92171
R200 VTAIL.n113 VTAIL.n112 8.92171
R201 VTAIL.n69 VTAIL.n68 8.92171
R202 VTAIL.n150 VTAIL.n144 8.14595
R203 VTAIL.n18 VTAIL.n12 8.14595
R204 VTAIL.n109 VTAIL.n103 8.14595
R205 VTAIL.n65 VTAIL.n59 8.14595
R206 VTAIL.n149 VTAIL.n146 7.3702
R207 VTAIL.n17 VTAIL.n14 7.3702
R208 VTAIL.n108 VTAIL.n105 7.3702
R209 VTAIL.n64 VTAIL.n61 7.3702
R210 VTAIL.n150 VTAIL.n149 5.81868
R211 VTAIL.n18 VTAIL.n17 5.81868
R212 VTAIL.n109 VTAIL.n108 5.81868
R213 VTAIL.n65 VTAIL.n64 5.81868
R214 VTAIL.n153 VTAIL.n144 5.04292
R215 VTAIL.n21 VTAIL.n12 5.04292
R216 VTAIL.n112 VTAIL.n103 5.04292
R217 VTAIL.n68 VTAIL.n59 5.04292
R218 VTAIL.n154 VTAIL.n142 4.26717
R219 VTAIL.n22 VTAIL.n10 4.26717
R220 VTAIL.n113 VTAIL.n101 4.26717
R221 VTAIL.n69 VTAIL.n57 4.26717
R222 VTAIL.n0 VTAIL.t4 4.15715
R223 VTAIL.n0 VTAIL.t2 4.15715
R224 VTAIL.n44 VTAIL.t9 4.15715
R225 VTAIL.n44 VTAIL.t10 4.15715
R226 VTAIL.n90 VTAIL.t7 4.15715
R227 VTAIL.n90 VTAIL.t8 4.15715
R228 VTAIL.n46 VTAIL.t5 4.15715
R229 VTAIL.n46 VTAIL.t0 4.15715
R230 VTAIL.n158 VTAIL.n157 3.49141
R231 VTAIL.n26 VTAIL.n25 3.49141
R232 VTAIL.n117 VTAIL.n116 3.49141
R233 VTAIL.n73 VTAIL.n72 3.49141
R234 VTAIL.n161 VTAIL.n140 2.71565
R235 VTAIL.n29 VTAIL.n8 2.71565
R236 VTAIL.n120 VTAIL.n99 2.71565
R237 VTAIL.n76 VTAIL.n55 2.71565
R238 VTAIL.n148 VTAIL.n147 2.4129
R239 VTAIL.n16 VTAIL.n15 2.4129
R240 VTAIL.n107 VTAIL.n106 2.4129
R241 VTAIL.n63 VTAIL.n62 2.4129
R242 VTAIL.n162 VTAIL.n138 1.93989
R243 VTAIL.n30 VTAIL.n6 1.93989
R244 VTAIL.n121 VTAIL.n97 1.93989
R245 VTAIL.n77 VTAIL.n53 1.93989
R246 VTAIL.n167 VTAIL.n165 1.16414
R247 VTAIL.n174 VTAIL.n134 1.16414
R248 VTAIL.n35 VTAIL.n33 1.16414
R249 VTAIL.n42 VTAIL.n2 1.16414
R250 VTAIL.n132 VTAIL.n92 1.16414
R251 VTAIL.n125 VTAIL.n124 1.16414
R252 VTAIL.n88 VTAIL.n48 1.16414
R253 VTAIL.n81 VTAIL.n80 1.16414
R254 VTAIL.n91 VTAIL.n89 0.897052
R255 VTAIL.n43 VTAIL.n1 0.897052
R256 VTAIL.n89 VTAIL.n47 0.853948
R257 VTAIL.n133 VTAIL.n91 0.853948
R258 VTAIL.n45 VTAIL.n43 0.853948
R259 VTAIL VTAIL.n175 0.582397
R260 VTAIL.n166 VTAIL.n136 0.388379
R261 VTAIL.n172 VTAIL.n171 0.388379
R262 VTAIL.n34 VTAIL.n4 0.388379
R263 VTAIL.n40 VTAIL.n39 0.388379
R264 VTAIL.n130 VTAIL.n129 0.388379
R265 VTAIL.n96 VTAIL.n94 0.388379
R266 VTAIL.n86 VTAIL.n85 0.388379
R267 VTAIL.n52 VTAIL.n50 0.388379
R268 VTAIL VTAIL.n1 0.272052
R269 VTAIL.n148 VTAIL.n143 0.155672
R270 VTAIL.n155 VTAIL.n143 0.155672
R271 VTAIL.n156 VTAIL.n155 0.155672
R272 VTAIL.n156 VTAIL.n139 0.155672
R273 VTAIL.n163 VTAIL.n139 0.155672
R274 VTAIL.n164 VTAIL.n163 0.155672
R275 VTAIL.n164 VTAIL.n135 0.155672
R276 VTAIL.n173 VTAIL.n135 0.155672
R277 VTAIL.n16 VTAIL.n11 0.155672
R278 VTAIL.n23 VTAIL.n11 0.155672
R279 VTAIL.n24 VTAIL.n23 0.155672
R280 VTAIL.n24 VTAIL.n7 0.155672
R281 VTAIL.n31 VTAIL.n7 0.155672
R282 VTAIL.n32 VTAIL.n31 0.155672
R283 VTAIL.n32 VTAIL.n3 0.155672
R284 VTAIL.n41 VTAIL.n3 0.155672
R285 VTAIL.n131 VTAIL.n93 0.155672
R286 VTAIL.n123 VTAIL.n93 0.155672
R287 VTAIL.n123 VTAIL.n122 0.155672
R288 VTAIL.n122 VTAIL.n98 0.155672
R289 VTAIL.n115 VTAIL.n98 0.155672
R290 VTAIL.n115 VTAIL.n114 0.155672
R291 VTAIL.n114 VTAIL.n102 0.155672
R292 VTAIL.n107 VTAIL.n102 0.155672
R293 VTAIL.n87 VTAIL.n49 0.155672
R294 VTAIL.n79 VTAIL.n49 0.155672
R295 VTAIL.n79 VTAIL.n78 0.155672
R296 VTAIL.n78 VTAIL.n54 0.155672
R297 VTAIL.n71 VTAIL.n54 0.155672
R298 VTAIL.n71 VTAIL.n70 0.155672
R299 VTAIL.n70 VTAIL.n58 0.155672
R300 VTAIL.n63 VTAIL.n58 0.155672
R301 VDD1.n36 VDD1.n0 756.745
R302 VDD1.n77 VDD1.n41 756.745
R303 VDD1.n37 VDD1.n36 585
R304 VDD1.n35 VDD1.n2 585
R305 VDD1.n34 VDD1.n33 585
R306 VDD1.n5 VDD1.n3 585
R307 VDD1.n28 VDD1.n27 585
R308 VDD1.n26 VDD1.n25 585
R309 VDD1.n9 VDD1.n8 585
R310 VDD1.n20 VDD1.n19 585
R311 VDD1.n18 VDD1.n17 585
R312 VDD1.n13 VDD1.n12 585
R313 VDD1.n53 VDD1.n52 585
R314 VDD1.n58 VDD1.n57 585
R315 VDD1.n60 VDD1.n59 585
R316 VDD1.n49 VDD1.n48 585
R317 VDD1.n66 VDD1.n65 585
R318 VDD1.n68 VDD1.n67 585
R319 VDD1.n45 VDD1.n44 585
R320 VDD1.n75 VDD1.n74 585
R321 VDD1.n76 VDD1.n43 585
R322 VDD1.n78 VDD1.n77 585
R323 VDD1.n14 VDD1.t3 329.043
R324 VDD1.n54 VDD1.t5 329.043
R325 VDD1.n36 VDD1.n35 171.744
R326 VDD1.n35 VDD1.n34 171.744
R327 VDD1.n34 VDD1.n3 171.744
R328 VDD1.n27 VDD1.n3 171.744
R329 VDD1.n27 VDD1.n26 171.744
R330 VDD1.n26 VDD1.n8 171.744
R331 VDD1.n19 VDD1.n8 171.744
R332 VDD1.n19 VDD1.n18 171.744
R333 VDD1.n18 VDD1.n12 171.744
R334 VDD1.n58 VDD1.n52 171.744
R335 VDD1.n59 VDD1.n58 171.744
R336 VDD1.n59 VDD1.n48 171.744
R337 VDD1.n66 VDD1.n48 171.744
R338 VDD1.n67 VDD1.n66 171.744
R339 VDD1.n67 VDD1.n44 171.744
R340 VDD1.n75 VDD1.n44 171.744
R341 VDD1.n76 VDD1.n75 171.744
R342 VDD1.n77 VDD1.n76 171.744
R343 VDD1.t3 VDD1.n12 85.8723
R344 VDD1.t5 VDD1.n52 85.8723
R345 VDD1.n83 VDD1.n82 82.9049
R346 VDD1.n85 VDD1.n84 82.7469
R347 VDD1 VDD1.n40 49.9503
R348 VDD1.n83 VDD1.n81 49.8368
R349 VDD1.n85 VDD1.n83 34.2401
R350 VDD1.n37 VDD1.n2 13.1884
R351 VDD1.n78 VDD1.n43 13.1884
R352 VDD1.n38 VDD1.n0 12.8005
R353 VDD1.n33 VDD1.n4 12.8005
R354 VDD1.n74 VDD1.n73 12.8005
R355 VDD1.n79 VDD1.n41 12.8005
R356 VDD1.n32 VDD1.n5 12.0247
R357 VDD1.n72 VDD1.n45 12.0247
R358 VDD1.n29 VDD1.n28 11.249
R359 VDD1.n69 VDD1.n68 11.249
R360 VDD1.n14 VDD1.n13 10.7238
R361 VDD1.n54 VDD1.n53 10.7238
R362 VDD1.n25 VDD1.n7 10.4732
R363 VDD1.n65 VDD1.n47 10.4732
R364 VDD1.n24 VDD1.n9 9.69747
R365 VDD1.n64 VDD1.n49 9.69747
R366 VDD1.n40 VDD1.n39 9.45567
R367 VDD1.n81 VDD1.n80 9.45567
R368 VDD1.n16 VDD1.n15 9.3005
R369 VDD1.n11 VDD1.n10 9.3005
R370 VDD1.n22 VDD1.n21 9.3005
R371 VDD1.n24 VDD1.n23 9.3005
R372 VDD1.n7 VDD1.n6 9.3005
R373 VDD1.n30 VDD1.n29 9.3005
R374 VDD1.n32 VDD1.n31 9.3005
R375 VDD1.n4 VDD1.n1 9.3005
R376 VDD1.n39 VDD1.n38 9.3005
R377 VDD1.n80 VDD1.n79 9.3005
R378 VDD1.n56 VDD1.n55 9.3005
R379 VDD1.n51 VDD1.n50 9.3005
R380 VDD1.n62 VDD1.n61 9.3005
R381 VDD1.n64 VDD1.n63 9.3005
R382 VDD1.n47 VDD1.n46 9.3005
R383 VDD1.n70 VDD1.n69 9.3005
R384 VDD1.n72 VDD1.n71 9.3005
R385 VDD1.n73 VDD1.n42 9.3005
R386 VDD1.n21 VDD1.n20 8.92171
R387 VDD1.n61 VDD1.n60 8.92171
R388 VDD1.n17 VDD1.n11 8.14595
R389 VDD1.n57 VDD1.n51 8.14595
R390 VDD1.n16 VDD1.n13 7.3702
R391 VDD1.n56 VDD1.n53 7.3702
R392 VDD1.n17 VDD1.n16 5.81868
R393 VDD1.n57 VDD1.n56 5.81868
R394 VDD1.n20 VDD1.n11 5.04292
R395 VDD1.n60 VDD1.n51 5.04292
R396 VDD1.n21 VDD1.n9 4.26717
R397 VDD1.n61 VDD1.n49 4.26717
R398 VDD1.n84 VDD1.t2 4.15715
R399 VDD1.n84 VDD1.t1 4.15715
R400 VDD1.n82 VDD1.t4 4.15715
R401 VDD1.n82 VDD1.t0 4.15715
R402 VDD1.n25 VDD1.n24 3.49141
R403 VDD1.n65 VDD1.n64 3.49141
R404 VDD1.n28 VDD1.n7 2.71565
R405 VDD1.n68 VDD1.n47 2.71565
R406 VDD1.n15 VDD1.n14 2.4129
R407 VDD1.n55 VDD1.n54 2.4129
R408 VDD1.n29 VDD1.n5 1.93989
R409 VDD1.n69 VDD1.n45 1.93989
R410 VDD1.n40 VDD1.n0 1.16414
R411 VDD1.n33 VDD1.n32 1.16414
R412 VDD1.n74 VDD1.n72 1.16414
R413 VDD1.n81 VDD1.n41 1.16414
R414 VDD1.n38 VDD1.n37 0.388379
R415 VDD1.n4 VDD1.n2 0.388379
R416 VDD1.n73 VDD1.n43 0.388379
R417 VDD1.n79 VDD1.n78 0.388379
R418 VDD1.n39 VDD1.n1 0.155672
R419 VDD1.n31 VDD1.n1 0.155672
R420 VDD1.n31 VDD1.n30 0.155672
R421 VDD1.n30 VDD1.n6 0.155672
R422 VDD1.n23 VDD1.n6 0.155672
R423 VDD1.n23 VDD1.n22 0.155672
R424 VDD1.n22 VDD1.n10 0.155672
R425 VDD1.n15 VDD1.n10 0.155672
R426 VDD1.n55 VDD1.n50 0.155672
R427 VDD1.n62 VDD1.n50 0.155672
R428 VDD1.n63 VDD1.n62 0.155672
R429 VDD1.n63 VDD1.n46 0.155672
R430 VDD1.n70 VDD1.n46 0.155672
R431 VDD1.n71 VDD1.n70 0.155672
R432 VDD1.n71 VDD1.n42 0.155672
R433 VDD1.n80 VDD1.n42 0.155672
R434 VDD1 VDD1.n85 0.155672
R435 B.n247 B.n70 585
R436 B.n246 B.n245 585
R437 B.n244 B.n71 585
R438 B.n243 B.n242 585
R439 B.n241 B.n72 585
R440 B.n240 B.n239 585
R441 B.n238 B.n73 585
R442 B.n237 B.n236 585
R443 B.n235 B.n74 585
R444 B.n234 B.n233 585
R445 B.n232 B.n75 585
R446 B.n231 B.n230 585
R447 B.n229 B.n76 585
R448 B.n228 B.n227 585
R449 B.n226 B.n77 585
R450 B.n225 B.n224 585
R451 B.n223 B.n78 585
R452 B.n222 B.n221 585
R453 B.n220 B.n79 585
R454 B.n219 B.n218 585
R455 B.n217 B.n80 585
R456 B.n216 B.n215 585
R457 B.n214 B.n81 585
R458 B.n213 B.n212 585
R459 B.n211 B.n82 585
R460 B.n210 B.n209 585
R461 B.n208 B.n83 585
R462 B.n207 B.n206 585
R463 B.n205 B.n84 585
R464 B.n204 B.n203 585
R465 B.n199 B.n85 585
R466 B.n198 B.n197 585
R467 B.n196 B.n86 585
R468 B.n195 B.n194 585
R469 B.n193 B.n87 585
R470 B.n192 B.n191 585
R471 B.n190 B.n88 585
R472 B.n189 B.n188 585
R473 B.n187 B.n89 585
R474 B.n185 B.n184 585
R475 B.n183 B.n92 585
R476 B.n182 B.n181 585
R477 B.n180 B.n93 585
R478 B.n179 B.n178 585
R479 B.n177 B.n94 585
R480 B.n176 B.n175 585
R481 B.n174 B.n95 585
R482 B.n173 B.n172 585
R483 B.n171 B.n96 585
R484 B.n170 B.n169 585
R485 B.n168 B.n97 585
R486 B.n167 B.n166 585
R487 B.n165 B.n98 585
R488 B.n164 B.n163 585
R489 B.n162 B.n99 585
R490 B.n161 B.n160 585
R491 B.n159 B.n100 585
R492 B.n158 B.n157 585
R493 B.n156 B.n101 585
R494 B.n155 B.n154 585
R495 B.n153 B.n102 585
R496 B.n152 B.n151 585
R497 B.n150 B.n103 585
R498 B.n149 B.n148 585
R499 B.n147 B.n104 585
R500 B.n146 B.n145 585
R501 B.n144 B.n105 585
R502 B.n143 B.n142 585
R503 B.n249 B.n248 585
R504 B.n250 B.n69 585
R505 B.n252 B.n251 585
R506 B.n253 B.n68 585
R507 B.n255 B.n254 585
R508 B.n256 B.n67 585
R509 B.n258 B.n257 585
R510 B.n259 B.n66 585
R511 B.n261 B.n260 585
R512 B.n262 B.n65 585
R513 B.n264 B.n263 585
R514 B.n265 B.n64 585
R515 B.n267 B.n266 585
R516 B.n268 B.n63 585
R517 B.n270 B.n269 585
R518 B.n271 B.n62 585
R519 B.n273 B.n272 585
R520 B.n274 B.n61 585
R521 B.n276 B.n275 585
R522 B.n277 B.n60 585
R523 B.n279 B.n278 585
R524 B.n280 B.n59 585
R525 B.n282 B.n281 585
R526 B.n283 B.n58 585
R527 B.n285 B.n284 585
R528 B.n286 B.n57 585
R529 B.n288 B.n287 585
R530 B.n289 B.n56 585
R531 B.n291 B.n290 585
R532 B.n292 B.n55 585
R533 B.n294 B.n293 585
R534 B.n295 B.n54 585
R535 B.n297 B.n296 585
R536 B.n298 B.n53 585
R537 B.n300 B.n299 585
R538 B.n301 B.n52 585
R539 B.n303 B.n302 585
R540 B.n304 B.n51 585
R541 B.n306 B.n305 585
R542 B.n307 B.n50 585
R543 B.n411 B.n410 585
R544 B.n409 B.n12 585
R545 B.n408 B.n407 585
R546 B.n406 B.n13 585
R547 B.n405 B.n404 585
R548 B.n403 B.n14 585
R549 B.n402 B.n401 585
R550 B.n400 B.n15 585
R551 B.n399 B.n398 585
R552 B.n397 B.n16 585
R553 B.n396 B.n395 585
R554 B.n394 B.n17 585
R555 B.n393 B.n392 585
R556 B.n391 B.n18 585
R557 B.n390 B.n389 585
R558 B.n388 B.n19 585
R559 B.n387 B.n386 585
R560 B.n385 B.n20 585
R561 B.n384 B.n383 585
R562 B.n382 B.n21 585
R563 B.n381 B.n380 585
R564 B.n379 B.n22 585
R565 B.n378 B.n377 585
R566 B.n376 B.n23 585
R567 B.n375 B.n374 585
R568 B.n373 B.n24 585
R569 B.n372 B.n371 585
R570 B.n370 B.n25 585
R571 B.n369 B.n368 585
R572 B.n367 B.n366 585
R573 B.n365 B.n29 585
R574 B.n364 B.n363 585
R575 B.n362 B.n30 585
R576 B.n361 B.n360 585
R577 B.n359 B.n31 585
R578 B.n358 B.n357 585
R579 B.n356 B.n32 585
R580 B.n355 B.n354 585
R581 B.n353 B.n33 585
R582 B.n351 B.n350 585
R583 B.n349 B.n36 585
R584 B.n348 B.n347 585
R585 B.n346 B.n37 585
R586 B.n345 B.n344 585
R587 B.n343 B.n38 585
R588 B.n342 B.n341 585
R589 B.n340 B.n39 585
R590 B.n339 B.n338 585
R591 B.n337 B.n40 585
R592 B.n336 B.n335 585
R593 B.n334 B.n41 585
R594 B.n333 B.n332 585
R595 B.n331 B.n42 585
R596 B.n330 B.n329 585
R597 B.n328 B.n43 585
R598 B.n327 B.n326 585
R599 B.n325 B.n44 585
R600 B.n324 B.n323 585
R601 B.n322 B.n45 585
R602 B.n321 B.n320 585
R603 B.n319 B.n46 585
R604 B.n318 B.n317 585
R605 B.n316 B.n47 585
R606 B.n315 B.n314 585
R607 B.n313 B.n48 585
R608 B.n312 B.n311 585
R609 B.n310 B.n49 585
R610 B.n309 B.n308 585
R611 B.n412 B.n11 585
R612 B.n414 B.n413 585
R613 B.n415 B.n10 585
R614 B.n417 B.n416 585
R615 B.n418 B.n9 585
R616 B.n420 B.n419 585
R617 B.n421 B.n8 585
R618 B.n423 B.n422 585
R619 B.n424 B.n7 585
R620 B.n426 B.n425 585
R621 B.n427 B.n6 585
R622 B.n429 B.n428 585
R623 B.n430 B.n5 585
R624 B.n432 B.n431 585
R625 B.n433 B.n4 585
R626 B.n435 B.n434 585
R627 B.n436 B.n3 585
R628 B.n438 B.n437 585
R629 B.n439 B.n0 585
R630 B.n2 B.n1 585
R631 B.n116 B.n115 585
R632 B.n117 B.n114 585
R633 B.n119 B.n118 585
R634 B.n120 B.n113 585
R635 B.n122 B.n121 585
R636 B.n123 B.n112 585
R637 B.n125 B.n124 585
R638 B.n126 B.n111 585
R639 B.n128 B.n127 585
R640 B.n129 B.n110 585
R641 B.n131 B.n130 585
R642 B.n132 B.n109 585
R643 B.n134 B.n133 585
R644 B.n135 B.n108 585
R645 B.n137 B.n136 585
R646 B.n138 B.n107 585
R647 B.n140 B.n139 585
R648 B.n141 B.n106 585
R649 B.n142 B.n141 559.769
R650 B.n248 B.n247 559.769
R651 B.n308 B.n307 559.769
R652 B.n410 B.n11 559.769
R653 B.n90 B.t6 489.036
R654 B.n200 B.t3 489.036
R655 B.n34 B.t0 489.036
R656 B.n26 B.t9 489.036
R657 B.n200 B.t4 319.399
R658 B.n34 B.t2 319.399
R659 B.n90 B.t7 319.399
R660 B.n26 B.t11 319.399
R661 B.n201 B.t5 300.2
R662 B.n35 B.t1 300.2
R663 B.n91 B.t8 300.2
R664 B.n27 B.t10 300.2
R665 B.n441 B.n440 256.663
R666 B.n440 B.n439 235.042
R667 B.n440 B.n2 235.042
R668 B.n142 B.n105 163.367
R669 B.n146 B.n105 163.367
R670 B.n147 B.n146 163.367
R671 B.n148 B.n147 163.367
R672 B.n148 B.n103 163.367
R673 B.n152 B.n103 163.367
R674 B.n153 B.n152 163.367
R675 B.n154 B.n153 163.367
R676 B.n154 B.n101 163.367
R677 B.n158 B.n101 163.367
R678 B.n159 B.n158 163.367
R679 B.n160 B.n159 163.367
R680 B.n160 B.n99 163.367
R681 B.n164 B.n99 163.367
R682 B.n165 B.n164 163.367
R683 B.n166 B.n165 163.367
R684 B.n166 B.n97 163.367
R685 B.n170 B.n97 163.367
R686 B.n171 B.n170 163.367
R687 B.n172 B.n171 163.367
R688 B.n172 B.n95 163.367
R689 B.n176 B.n95 163.367
R690 B.n177 B.n176 163.367
R691 B.n178 B.n177 163.367
R692 B.n178 B.n93 163.367
R693 B.n182 B.n93 163.367
R694 B.n183 B.n182 163.367
R695 B.n184 B.n183 163.367
R696 B.n184 B.n89 163.367
R697 B.n189 B.n89 163.367
R698 B.n190 B.n189 163.367
R699 B.n191 B.n190 163.367
R700 B.n191 B.n87 163.367
R701 B.n195 B.n87 163.367
R702 B.n196 B.n195 163.367
R703 B.n197 B.n196 163.367
R704 B.n197 B.n85 163.367
R705 B.n204 B.n85 163.367
R706 B.n205 B.n204 163.367
R707 B.n206 B.n205 163.367
R708 B.n206 B.n83 163.367
R709 B.n210 B.n83 163.367
R710 B.n211 B.n210 163.367
R711 B.n212 B.n211 163.367
R712 B.n212 B.n81 163.367
R713 B.n216 B.n81 163.367
R714 B.n217 B.n216 163.367
R715 B.n218 B.n217 163.367
R716 B.n218 B.n79 163.367
R717 B.n222 B.n79 163.367
R718 B.n223 B.n222 163.367
R719 B.n224 B.n223 163.367
R720 B.n224 B.n77 163.367
R721 B.n228 B.n77 163.367
R722 B.n229 B.n228 163.367
R723 B.n230 B.n229 163.367
R724 B.n230 B.n75 163.367
R725 B.n234 B.n75 163.367
R726 B.n235 B.n234 163.367
R727 B.n236 B.n235 163.367
R728 B.n236 B.n73 163.367
R729 B.n240 B.n73 163.367
R730 B.n241 B.n240 163.367
R731 B.n242 B.n241 163.367
R732 B.n242 B.n71 163.367
R733 B.n246 B.n71 163.367
R734 B.n247 B.n246 163.367
R735 B.n307 B.n306 163.367
R736 B.n306 B.n51 163.367
R737 B.n302 B.n51 163.367
R738 B.n302 B.n301 163.367
R739 B.n301 B.n300 163.367
R740 B.n300 B.n53 163.367
R741 B.n296 B.n53 163.367
R742 B.n296 B.n295 163.367
R743 B.n295 B.n294 163.367
R744 B.n294 B.n55 163.367
R745 B.n290 B.n55 163.367
R746 B.n290 B.n289 163.367
R747 B.n289 B.n288 163.367
R748 B.n288 B.n57 163.367
R749 B.n284 B.n57 163.367
R750 B.n284 B.n283 163.367
R751 B.n283 B.n282 163.367
R752 B.n282 B.n59 163.367
R753 B.n278 B.n59 163.367
R754 B.n278 B.n277 163.367
R755 B.n277 B.n276 163.367
R756 B.n276 B.n61 163.367
R757 B.n272 B.n61 163.367
R758 B.n272 B.n271 163.367
R759 B.n271 B.n270 163.367
R760 B.n270 B.n63 163.367
R761 B.n266 B.n63 163.367
R762 B.n266 B.n265 163.367
R763 B.n265 B.n264 163.367
R764 B.n264 B.n65 163.367
R765 B.n260 B.n65 163.367
R766 B.n260 B.n259 163.367
R767 B.n259 B.n258 163.367
R768 B.n258 B.n67 163.367
R769 B.n254 B.n67 163.367
R770 B.n254 B.n253 163.367
R771 B.n253 B.n252 163.367
R772 B.n252 B.n69 163.367
R773 B.n248 B.n69 163.367
R774 B.n410 B.n409 163.367
R775 B.n409 B.n408 163.367
R776 B.n408 B.n13 163.367
R777 B.n404 B.n13 163.367
R778 B.n404 B.n403 163.367
R779 B.n403 B.n402 163.367
R780 B.n402 B.n15 163.367
R781 B.n398 B.n15 163.367
R782 B.n398 B.n397 163.367
R783 B.n397 B.n396 163.367
R784 B.n396 B.n17 163.367
R785 B.n392 B.n17 163.367
R786 B.n392 B.n391 163.367
R787 B.n391 B.n390 163.367
R788 B.n390 B.n19 163.367
R789 B.n386 B.n19 163.367
R790 B.n386 B.n385 163.367
R791 B.n385 B.n384 163.367
R792 B.n384 B.n21 163.367
R793 B.n380 B.n21 163.367
R794 B.n380 B.n379 163.367
R795 B.n379 B.n378 163.367
R796 B.n378 B.n23 163.367
R797 B.n374 B.n23 163.367
R798 B.n374 B.n373 163.367
R799 B.n373 B.n372 163.367
R800 B.n372 B.n25 163.367
R801 B.n368 B.n25 163.367
R802 B.n368 B.n367 163.367
R803 B.n367 B.n29 163.367
R804 B.n363 B.n29 163.367
R805 B.n363 B.n362 163.367
R806 B.n362 B.n361 163.367
R807 B.n361 B.n31 163.367
R808 B.n357 B.n31 163.367
R809 B.n357 B.n356 163.367
R810 B.n356 B.n355 163.367
R811 B.n355 B.n33 163.367
R812 B.n350 B.n33 163.367
R813 B.n350 B.n349 163.367
R814 B.n349 B.n348 163.367
R815 B.n348 B.n37 163.367
R816 B.n344 B.n37 163.367
R817 B.n344 B.n343 163.367
R818 B.n343 B.n342 163.367
R819 B.n342 B.n39 163.367
R820 B.n338 B.n39 163.367
R821 B.n338 B.n337 163.367
R822 B.n337 B.n336 163.367
R823 B.n336 B.n41 163.367
R824 B.n332 B.n41 163.367
R825 B.n332 B.n331 163.367
R826 B.n331 B.n330 163.367
R827 B.n330 B.n43 163.367
R828 B.n326 B.n43 163.367
R829 B.n326 B.n325 163.367
R830 B.n325 B.n324 163.367
R831 B.n324 B.n45 163.367
R832 B.n320 B.n45 163.367
R833 B.n320 B.n319 163.367
R834 B.n319 B.n318 163.367
R835 B.n318 B.n47 163.367
R836 B.n314 B.n47 163.367
R837 B.n314 B.n313 163.367
R838 B.n313 B.n312 163.367
R839 B.n312 B.n49 163.367
R840 B.n308 B.n49 163.367
R841 B.n414 B.n11 163.367
R842 B.n415 B.n414 163.367
R843 B.n416 B.n415 163.367
R844 B.n416 B.n9 163.367
R845 B.n420 B.n9 163.367
R846 B.n421 B.n420 163.367
R847 B.n422 B.n421 163.367
R848 B.n422 B.n7 163.367
R849 B.n426 B.n7 163.367
R850 B.n427 B.n426 163.367
R851 B.n428 B.n427 163.367
R852 B.n428 B.n5 163.367
R853 B.n432 B.n5 163.367
R854 B.n433 B.n432 163.367
R855 B.n434 B.n433 163.367
R856 B.n434 B.n3 163.367
R857 B.n438 B.n3 163.367
R858 B.n439 B.n438 163.367
R859 B.n116 B.n2 163.367
R860 B.n117 B.n116 163.367
R861 B.n118 B.n117 163.367
R862 B.n118 B.n113 163.367
R863 B.n122 B.n113 163.367
R864 B.n123 B.n122 163.367
R865 B.n124 B.n123 163.367
R866 B.n124 B.n111 163.367
R867 B.n128 B.n111 163.367
R868 B.n129 B.n128 163.367
R869 B.n130 B.n129 163.367
R870 B.n130 B.n109 163.367
R871 B.n134 B.n109 163.367
R872 B.n135 B.n134 163.367
R873 B.n136 B.n135 163.367
R874 B.n136 B.n107 163.367
R875 B.n140 B.n107 163.367
R876 B.n141 B.n140 163.367
R877 B.n186 B.n91 59.5399
R878 B.n202 B.n201 59.5399
R879 B.n352 B.n35 59.5399
R880 B.n28 B.n27 59.5399
R881 B.n249 B.n70 36.3712
R882 B.n412 B.n411 36.3712
R883 B.n309 B.n50 36.3712
R884 B.n143 B.n106 36.3712
R885 B.n91 B.n90 19.2005
R886 B.n201 B.n200 19.2005
R887 B.n35 B.n34 19.2005
R888 B.n27 B.n26 19.2005
R889 B B.n441 18.0485
R890 B.n413 B.n412 10.6151
R891 B.n413 B.n10 10.6151
R892 B.n417 B.n10 10.6151
R893 B.n418 B.n417 10.6151
R894 B.n419 B.n418 10.6151
R895 B.n419 B.n8 10.6151
R896 B.n423 B.n8 10.6151
R897 B.n424 B.n423 10.6151
R898 B.n425 B.n424 10.6151
R899 B.n425 B.n6 10.6151
R900 B.n429 B.n6 10.6151
R901 B.n430 B.n429 10.6151
R902 B.n431 B.n430 10.6151
R903 B.n431 B.n4 10.6151
R904 B.n435 B.n4 10.6151
R905 B.n436 B.n435 10.6151
R906 B.n437 B.n436 10.6151
R907 B.n437 B.n0 10.6151
R908 B.n411 B.n12 10.6151
R909 B.n407 B.n12 10.6151
R910 B.n407 B.n406 10.6151
R911 B.n406 B.n405 10.6151
R912 B.n405 B.n14 10.6151
R913 B.n401 B.n14 10.6151
R914 B.n401 B.n400 10.6151
R915 B.n400 B.n399 10.6151
R916 B.n399 B.n16 10.6151
R917 B.n395 B.n16 10.6151
R918 B.n395 B.n394 10.6151
R919 B.n394 B.n393 10.6151
R920 B.n393 B.n18 10.6151
R921 B.n389 B.n18 10.6151
R922 B.n389 B.n388 10.6151
R923 B.n388 B.n387 10.6151
R924 B.n387 B.n20 10.6151
R925 B.n383 B.n20 10.6151
R926 B.n383 B.n382 10.6151
R927 B.n382 B.n381 10.6151
R928 B.n381 B.n22 10.6151
R929 B.n377 B.n22 10.6151
R930 B.n377 B.n376 10.6151
R931 B.n376 B.n375 10.6151
R932 B.n375 B.n24 10.6151
R933 B.n371 B.n24 10.6151
R934 B.n371 B.n370 10.6151
R935 B.n370 B.n369 10.6151
R936 B.n366 B.n365 10.6151
R937 B.n365 B.n364 10.6151
R938 B.n364 B.n30 10.6151
R939 B.n360 B.n30 10.6151
R940 B.n360 B.n359 10.6151
R941 B.n359 B.n358 10.6151
R942 B.n358 B.n32 10.6151
R943 B.n354 B.n32 10.6151
R944 B.n354 B.n353 10.6151
R945 B.n351 B.n36 10.6151
R946 B.n347 B.n36 10.6151
R947 B.n347 B.n346 10.6151
R948 B.n346 B.n345 10.6151
R949 B.n345 B.n38 10.6151
R950 B.n341 B.n38 10.6151
R951 B.n341 B.n340 10.6151
R952 B.n340 B.n339 10.6151
R953 B.n339 B.n40 10.6151
R954 B.n335 B.n40 10.6151
R955 B.n335 B.n334 10.6151
R956 B.n334 B.n333 10.6151
R957 B.n333 B.n42 10.6151
R958 B.n329 B.n42 10.6151
R959 B.n329 B.n328 10.6151
R960 B.n328 B.n327 10.6151
R961 B.n327 B.n44 10.6151
R962 B.n323 B.n44 10.6151
R963 B.n323 B.n322 10.6151
R964 B.n322 B.n321 10.6151
R965 B.n321 B.n46 10.6151
R966 B.n317 B.n46 10.6151
R967 B.n317 B.n316 10.6151
R968 B.n316 B.n315 10.6151
R969 B.n315 B.n48 10.6151
R970 B.n311 B.n48 10.6151
R971 B.n311 B.n310 10.6151
R972 B.n310 B.n309 10.6151
R973 B.n305 B.n50 10.6151
R974 B.n305 B.n304 10.6151
R975 B.n304 B.n303 10.6151
R976 B.n303 B.n52 10.6151
R977 B.n299 B.n52 10.6151
R978 B.n299 B.n298 10.6151
R979 B.n298 B.n297 10.6151
R980 B.n297 B.n54 10.6151
R981 B.n293 B.n54 10.6151
R982 B.n293 B.n292 10.6151
R983 B.n292 B.n291 10.6151
R984 B.n291 B.n56 10.6151
R985 B.n287 B.n56 10.6151
R986 B.n287 B.n286 10.6151
R987 B.n286 B.n285 10.6151
R988 B.n285 B.n58 10.6151
R989 B.n281 B.n58 10.6151
R990 B.n281 B.n280 10.6151
R991 B.n280 B.n279 10.6151
R992 B.n279 B.n60 10.6151
R993 B.n275 B.n60 10.6151
R994 B.n275 B.n274 10.6151
R995 B.n274 B.n273 10.6151
R996 B.n273 B.n62 10.6151
R997 B.n269 B.n62 10.6151
R998 B.n269 B.n268 10.6151
R999 B.n268 B.n267 10.6151
R1000 B.n267 B.n64 10.6151
R1001 B.n263 B.n64 10.6151
R1002 B.n263 B.n262 10.6151
R1003 B.n262 B.n261 10.6151
R1004 B.n261 B.n66 10.6151
R1005 B.n257 B.n66 10.6151
R1006 B.n257 B.n256 10.6151
R1007 B.n256 B.n255 10.6151
R1008 B.n255 B.n68 10.6151
R1009 B.n251 B.n68 10.6151
R1010 B.n251 B.n250 10.6151
R1011 B.n250 B.n249 10.6151
R1012 B.n115 B.n1 10.6151
R1013 B.n115 B.n114 10.6151
R1014 B.n119 B.n114 10.6151
R1015 B.n120 B.n119 10.6151
R1016 B.n121 B.n120 10.6151
R1017 B.n121 B.n112 10.6151
R1018 B.n125 B.n112 10.6151
R1019 B.n126 B.n125 10.6151
R1020 B.n127 B.n126 10.6151
R1021 B.n127 B.n110 10.6151
R1022 B.n131 B.n110 10.6151
R1023 B.n132 B.n131 10.6151
R1024 B.n133 B.n132 10.6151
R1025 B.n133 B.n108 10.6151
R1026 B.n137 B.n108 10.6151
R1027 B.n138 B.n137 10.6151
R1028 B.n139 B.n138 10.6151
R1029 B.n139 B.n106 10.6151
R1030 B.n144 B.n143 10.6151
R1031 B.n145 B.n144 10.6151
R1032 B.n145 B.n104 10.6151
R1033 B.n149 B.n104 10.6151
R1034 B.n150 B.n149 10.6151
R1035 B.n151 B.n150 10.6151
R1036 B.n151 B.n102 10.6151
R1037 B.n155 B.n102 10.6151
R1038 B.n156 B.n155 10.6151
R1039 B.n157 B.n156 10.6151
R1040 B.n157 B.n100 10.6151
R1041 B.n161 B.n100 10.6151
R1042 B.n162 B.n161 10.6151
R1043 B.n163 B.n162 10.6151
R1044 B.n163 B.n98 10.6151
R1045 B.n167 B.n98 10.6151
R1046 B.n168 B.n167 10.6151
R1047 B.n169 B.n168 10.6151
R1048 B.n169 B.n96 10.6151
R1049 B.n173 B.n96 10.6151
R1050 B.n174 B.n173 10.6151
R1051 B.n175 B.n174 10.6151
R1052 B.n175 B.n94 10.6151
R1053 B.n179 B.n94 10.6151
R1054 B.n180 B.n179 10.6151
R1055 B.n181 B.n180 10.6151
R1056 B.n181 B.n92 10.6151
R1057 B.n185 B.n92 10.6151
R1058 B.n188 B.n187 10.6151
R1059 B.n188 B.n88 10.6151
R1060 B.n192 B.n88 10.6151
R1061 B.n193 B.n192 10.6151
R1062 B.n194 B.n193 10.6151
R1063 B.n194 B.n86 10.6151
R1064 B.n198 B.n86 10.6151
R1065 B.n199 B.n198 10.6151
R1066 B.n203 B.n199 10.6151
R1067 B.n207 B.n84 10.6151
R1068 B.n208 B.n207 10.6151
R1069 B.n209 B.n208 10.6151
R1070 B.n209 B.n82 10.6151
R1071 B.n213 B.n82 10.6151
R1072 B.n214 B.n213 10.6151
R1073 B.n215 B.n214 10.6151
R1074 B.n215 B.n80 10.6151
R1075 B.n219 B.n80 10.6151
R1076 B.n220 B.n219 10.6151
R1077 B.n221 B.n220 10.6151
R1078 B.n221 B.n78 10.6151
R1079 B.n225 B.n78 10.6151
R1080 B.n226 B.n225 10.6151
R1081 B.n227 B.n226 10.6151
R1082 B.n227 B.n76 10.6151
R1083 B.n231 B.n76 10.6151
R1084 B.n232 B.n231 10.6151
R1085 B.n233 B.n232 10.6151
R1086 B.n233 B.n74 10.6151
R1087 B.n237 B.n74 10.6151
R1088 B.n238 B.n237 10.6151
R1089 B.n239 B.n238 10.6151
R1090 B.n239 B.n72 10.6151
R1091 B.n243 B.n72 10.6151
R1092 B.n244 B.n243 10.6151
R1093 B.n245 B.n244 10.6151
R1094 B.n245 B.n70 10.6151
R1095 B.n369 B.n28 9.36635
R1096 B.n352 B.n351 9.36635
R1097 B.n186 B.n185 9.36635
R1098 B.n202 B.n84 9.36635
R1099 B.n441 B.n0 8.11757
R1100 B.n441 B.n1 8.11757
R1101 B.n366 B.n28 1.24928
R1102 B.n353 B.n352 1.24928
R1103 B.n187 B.n186 1.24928
R1104 B.n203 B.n202 1.24928
R1105 VN.n1 VN.t4 366.592
R1106 VN.n7 VN.t1 366.592
R1107 VN.n2 VN.t0 345.798
R1108 VN.n4 VN.t5 345.798
R1109 VN.n8 VN.t2 345.798
R1110 VN.n10 VN.t3 345.798
R1111 VN.n5 VN.n4 161.3
R1112 VN.n11 VN.n10 161.3
R1113 VN.n9 VN.n6 161.3
R1114 VN.n3 VN.n0 161.3
R1115 VN.n7 VN.n6 44.8515
R1116 VN.n1 VN.n0 44.8515
R1117 VN VN.n11 38.2183
R1118 VN.n3 VN.n2 24.8308
R1119 VN.n9 VN.n8 24.8308
R1120 VN.n4 VN.n3 23.3702
R1121 VN.n10 VN.n9 23.3702
R1122 VN.n2 VN.n1 21.148
R1123 VN.n8 VN.n7 21.148
R1124 VN.n11 VN.n6 0.189894
R1125 VN.n5 VN.n0 0.189894
R1126 VN VN.n5 0.0516364
R1127 VDD2.n79 VDD2.n43 756.745
R1128 VDD2.n36 VDD2.n0 756.745
R1129 VDD2.n80 VDD2.n79 585
R1130 VDD2.n78 VDD2.n45 585
R1131 VDD2.n77 VDD2.n76 585
R1132 VDD2.n48 VDD2.n46 585
R1133 VDD2.n71 VDD2.n70 585
R1134 VDD2.n69 VDD2.n68 585
R1135 VDD2.n52 VDD2.n51 585
R1136 VDD2.n63 VDD2.n62 585
R1137 VDD2.n61 VDD2.n60 585
R1138 VDD2.n56 VDD2.n55 585
R1139 VDD2.n12 VDD2.n11 585
R1140 VDD2.n17 VDD2.n16 585
R1141 VDD2.n19 VDD2.n18 585
R1142 VDD2.n8 VDD2.n7 585
R1143 VDD2.n25 VDD2.n24 585
R1144 VDD2.n27 VDD2.n26 585
R1145 VDD2.n4 VDD2.n3 585
R1146 VDD2.n34 VDD2.n33 585
R1147 VDD2.n35 VDD2.n2 585
R1148 VDD2.n37 VDD2.n36 585
R1149 VDD2.n57 VDD2.t2 329.043
R1150 VDD2.n13 VDD2.t1 329.043
R1151 VDD2.n79 VDD2.n78 171.744
R1152 VDD2.n78 VDD2.n77 171.744
R1153 VDD2.n77 VDD2.n46 171.744
R1154 VDD2.n70 VDD2.n46 171.744
R1155 VDD2.n70 VDD2.n69 171.744
R1156 VDD2.n69 VDD2.n51 171.744
R1157 VDD2.n62 VDD2.n51 171.744
R1158 VDD2.n62 VDD2.n61 171.744
R1159 VDD2.n61 VDD2.n55 171.744
R1160 VDD2.n17 VDD2.n11 171.744
R1161 VDD2.n18 VDD2.n17 171.744
R1162 VDD2.n18 VDD2.n7 171.744
R1163 VDD2.n25 VDD2.n7 171.744
R1164 VDD2.n26 VDD2.n25 171.744
R1165 VDD2.n26 VDD2.n3 171.744
R1166 VDD2.n34 VDD2.n3 171.744
R1167 VDD2.n35 VDD2.n34 171.744
R1168 VDD2.n36 VDD2.n35 171.744
R1169 VDD2.t2 VDD2.n55 85.8723
R1170 VDD2.t1 VDD2.n11 85.8723
R1171 VDD2.n42 VDD2.n41 82.9049
R1172 VDD2 VDD2.n85 82.9021
R1173 VDD2.n42 VDD2.n40 49.8368
R1174 VDD2.n84 VDD2.n83 49.252
R1175 VDD2.n84 VDD2.n42 33.2304
R1176 VDD2.n80 VDD2.n45 13.1884
R1177 VDD2.n37 VDD2.n2 13.1884
R1178 VDD2.n81 VDD2.n43 12.8005
R1179 VDD2.n76 VDD2.n47 12.8005
R1180 VDD2.n33 VDD2.n32 12.8005
R1181 VDD2.n38 VDD2.n0 12.8005
R1182 VDD2.n75 VDD2.n48 12.0247
R1183 VDD2.n31 VDD2.n4 12.0247
R1184 VDD2.n72 VDD2.n71 11.249
R1185 VDD2.n28 VDD2.n27 11.249
R1186 VDD2.n57 VDD2.n56 10.7238
R1187 VDD2.n13 VDD2.n12 10.7238
R1188 VDD2.n68 VDD2.n50 10.4732
R1189 VDD2.n24 VDD2.n6 10.4732
R1190 VDD2.n67 VDD2.n52 9.69747
R1191 VDD2.n23 VDD2.n8 9.69747
R1192 VDD2.n83 VDD2.n82 9.45567
R1193 VDD2.n40 VDD2.n39 9.45567
R1194 VDD2.n59 VDD2.n58 9.3005
R1195 VDD2.n54 VDD2.n53 9.3005
R1196 VDD2.n65 VDD2.n64 9.3005
R1197 VDD2.n67 VDD2.n66 9.3005
R1198 VDD2.n50 VDD2.n49 9.3005
R1199 VDD2.n73 VDD2.n72 9.3005
R1200 VDD2.n75 VDD2.n74 9.3005
R1201 VDD2.n47 VDD2.n44 9.3005
R1202 VDD2.n82 VDD2.n81 9.3005
R1203 VDD2.n39 VDD2.n38 9.3005
R1204 VDD2.n15 VDD2.n14 9.3005
R1205 VDD2.n10 VDD2.n9 9.3005
R1206 VDD2.n21 VDD2.n20 9.3005
R1207 VDD2.n23 VDD2.n22 9.3005
R1208 VDD2.n6 VDD2.n5 9.3005
R1209 VDD2.n29 VDD2.n28 9.3005
R1210 VDD2.n31 VDD2.n30 9.3005
R1211 VDD2.n32 VDD2.n1 9.3005
R1212 VDD2.n64 VDD2.n63 8.92171
R1213 VDD2.n20 VDD2.n19 8.92171
R1214 VDD2.n60 VDD2.n54 8.14595
R1215 VDD2.n16 VDD2.n10 8.14595
R1216 VDD2.n59 VDD2.n56 7.3702
R1217 VDD2.n15 VDD2.n12 7.3702
R1218 VDD2.n60 VDD2.n59 5.81868
R1219 VDD2.n16 VDD2.n15 5.81868
R1220 VDD2.n63 VDD2.n54 5.04292
R1221 VDD2.n19 VDD2.n10 5.04292
R1222 VDD2.n64 VDD2.n52 4.26717
R1223 VDD2.n20 VDD2.n8 4.26717
R1224 VDD2.n85 VDD2.t3 4.15715
R1225 VDD2.n85 VDD2.t4 4.15715
R1226 VDD2.n41 VDD2.t5 4.15715
R1227 VDD2.n41 VDD2.t0 4.15715
R1228 VDD2.n68 VDD2.n67 3.49141
R1229 VDD2.n24 VDD2.n23 3.49141
R1230 VDD2.n71 VDD2.n50 2.71565
R1231 VDD2.n27 VDD2.n6 2.71565
R1232 VDD2.n58 VDD2.n57 2.4129
R1233 VDD2.n14 VDD2.n13 2.4129
R1234 VDD2.n72 VDD2.n48 1.93989
R1235 VDD2.n28 VDD2.n4 1.93989
R1236 VDD2.n83 VDD2.n43 1.16414
R1237 VDD2.n76 VDD2.n75 1.16414
R1238 VDD2.n33 VDD2.n31 1.16414
R1239 VDD2.n40 VDD2.n0 1.16414
R1240 VDD2 VDD2.n84 0.698776
R1241 VDD2.n81 VDD2.n80 0.388379
R1242 VDD2.n47 VDD2.n45 0.388379
R1243 VDD2.n32 VDD2.n2 0.388379
R1244 VDD2.n38 VDD2.n37 0.388379
R1245 VDD2.n82 VDD2.n44 0.155672
R1246 VDD2.n74 VDD2.n44 0.155672
R1247 VDD2.n74 VDD2.n73 0.155672
R1248 VDD2.n73 VDD2.n49 0.155672
R1249 VDD2.n66 VDD2.n49 0.155672
R1250 VDD2.n66 VDD2.n65 0.155672
R1251 VDD2.n65 VDD2.n53 0.155672
R1252 VDD2.n58 VDD2.n53 0.155672
R1253 VDD2.n14 VDD2.n9 0.155672
R1254 VDD2.n21 VDD2.n9 0.155672
R1255 VDD2.n22 VDD2.n21 0.155672
R1256 VDD2.n22 VDD2.n5 0.155672
R1257 VDD2.n29 VDD2.n5 0.155672
R1258 VDD2.n30 VDD2.n29 0.155672
R1259 VDD2.n30 VDD2.n1 0.155672
R1260 VDD2.n39 VDD2.n1 0.155672
C0 VN VDD2 2.86353f
C1 w_n1762_n2532# VDD1 1.4874f
C2 VP VDD1 3.00595f
C3 B VDD1 1.24404f
C4 VP w_n1762_n2532# 3.02994f
C5 VTAIL VDD1 7.26041f
C6 w_n1762_n2532# B 5.8262f
C7 VP B 1.06593f
C8 w_n1762_n2532# VTAIL 2.27209f
C9 VN VDD1 0.147518f
C10 VDD2 VDD1 0.693619f
C11 VP VTAIL 2.71743f
C12 VTAIL B 1.94234f
C13 VN w_n1762_n2532# 2.80755f
C14 w_n1762_n2532# VDD2 1.51023f
C15 VN VP 4.27376f
C16 VP VDD2 0.29304f
C17 VN B 0.704383f
C18 VDD2 B 1.27207f
C19 VN VTAIL 2.70299f
C20 VDD2 VTAIL 7.29643f
C21 VDD2 VSUBS 1.137366f
C22 VDD1 VSUBS 0.995421f
C23 VTAIL VSUBS 0.610321f
C24 VN VSUBS 4.10964f
C25 VP VSUBS 1.276006f
C26 B VSUBS 2.358378f
C27 w_n1762_n2532# VSUBS 55.3761f
C28 VDD2.n0 VSUBS 0.023725f
C29 VDD2.n1 VSUBS 0.023693f
C30 VDD2.n2 VSUBS 0.013106f
C31 VDD2.n3 VSUBS 0.030093f
C32 VDD2.n4 VSUBS 0.013481f
C33 VDD2.n5 VSUBS 0.023693f
C34 VDD2.n6 VSUBS 0.012732f
C35 VDD2.n7 VSUBS 0.030093f
C36 VDD2.n8 VSUBS 0.013481f
C37 VDD2.n9 VSUBS 0.023693f
C38 VDD2.n10 VSUBS 0.012732f
C39 VDD2.n11 VSUBS 0.02257f
C40 VDD2.n12 VSUBS 0.022637f
C41 VDD2.t1 VSUBS 0.064591f
C42 VDD2.n13 VSUBS 0.141882f
C43 VDD2.n14 VSUBS 0.730037f
C44 VDD2.n15 VSUBS 0.012732f
C45 VDD2.n16 VSUBS 0.013481f
C46 VDD2.n17 VSUBS 0.030093f
C47 VDD2.n18 VSUBS 0.030093f
C48 VDD2.n19 VSUBS 0.013481f
C49 VDD2.n20 VSUBS 0.012732f
C50 VDD2.n21 VSUBS 0.023693f
C51 VDD2.n22 VSUBS 0.023693f
C52 VDD2.n23 VSUBS 0.012732f
C53 VDD2.n24 VSUBS 0.013481f
C54 VDD2.n25 VSUBS 0.030093f
C55 VDD2.n26 VSUBS 0.030093f
C56 VDD2.n27 VSUBS 0.013481f
C57 VDD2.n28 VSUBS 0.012732f
C58 VDD2.n29 VSUBS 0.023693f
C59 VDD2.n30 VSUBS 0.023693f
C60 VDD2.n31 VSUBS 0.012732f
C61 VDD2.n32 VSUBS 0.012732f
C62 VDD2.n33 VSUBS 0.013481f
C63 VDD2.n34 VSUBS 0.030093f
C64 VDD2.n35 VSUBS 0.030093f
C65 VDD2.n36 VSUBS 0.064989f
C66 VDD2.n37 VSUBS 0.013106f
C67 VDD2.n38 VSUBS 0.012732f
C68 VDD2.n39 VSUBS 0.055413f
C69 VDD2.n40 VSUBS 0.049782f
C70 VDD2.t5 VSUBS 0.146415f
C71 VDD2.t0 VSUBS 0.146415f
C72 VDD2.n41 VSUBS 1.05246f
C73 VDD2.n42 VSUBS 1.70907f
C74 VDD2.n43 VSUBS 0.023725f
C75 VDD2.n44 VSUBS 0.023693f
C76 VDD2.n45 VSUBS 0.013106f
C77 VDD2.n46 VSUBS 0.030093f
C78 VDD2.n47 VSUBS 0.012732f
C79 VDD2.n48 VSUBS 0.013481f
C80 VDD2.n49 VSUBS 0.023693f
C81 VDD2.n50 VSUBS 0.012732f
C82 VDD2.n51 VSUBS 0.030093f
C83 VDD2.n52 VSUBS 0.013481f
C84 VDD2.n53 VSUBS 0.023693f
C85 VDD2.n54 VSUBS 0.012732f
C86 VDD2.n55 VSUBS 0.02257f
C87 VDD2.n56 VSUBS 0.022637f
C88 VDD2.t2 VSUBS 0.064591f
C89 VDD2.n57 VSUBS 0.141882f
C90 VDD2.n58 VSUBS 0.730037f
C91 VDD2.n59 VSUBS 0.012732f
C92 VDD2.n60 VSUBS 0.013481f
C93 VDD2.n61 VSUBS 0.030093f
C94 VDD2.n62 VSUBS 0.030093f
C95 VDD2.n63 VSUBS 0.013481f
C96 VDD2.n64 VSUBS 0.012732f
C97 VDD2.n65 VSUBS 0.023693f
C98 VDD2.n66 VSUBS 0.023693f
C99 VDD2.n67 VSUBS 0.012732f
C100 VDD2.n68 VSUBS 0.013481f
C101 VDD2.n69 VSUBS 0.030093f
C102 VDD2.n70 VSUBS 0.030093f
C103 VDD2.n71 VSUBS 0.013481f
C104 VDD2.n72 VSUBS 0.012732f
C105 VDD2.n73 VSUBS 0.023693f
C106 VDD2.n74 VSUBS 0.023693f
C107 VDD2.n75 VSUBS 0.012732f
C108 VDD2.n76 VSUBS 0.013481f
C109 VDD2.n77 VSUBS 0.030093f
C110 VDD2.n78 VSUBS 0.030093f
C111 VDD2.n79 VSUBS 0.064989f
C112 VDD2.n80 VSUBS 0.013106f
C113 VDD2.n81 VSUBS 0.012732f
C114 VDD2.n82 VSUBS 0.055413f
C115 VDD2.n83 VSUBS 0.048707f
C116 VDD2.n84 VSUBS 1.61396f
C117 VDD2.t3 VSUBS 0.146415f
C118 VDD2.t4 VSUBS 0.146415f
C119 VDD2.n85 VSUBS 1.05243f
C120 VN.n0 VSUBS 0.248354f
C121 VN.t4 VSUBS 0.930105f
C122 VN.n1 VSUBS 0.37736f
C123 VN.t0 VSUBS 0.907775f
C124 VN.n2 VSUBS 0.399868f
C125 VN.n3 VSUBS 0.013858f
C126 VN.t5 VSUBS 0.907775f
C127 VN.n4 VSUBS 0.388866f
C128 VN.n5 VSUBS 0.047326f
C129 VN.n6 VSUBS 0.248354f
C130 VN.t1 VSUBS 0.930105f
C131 VN.n7 VSUBS 0.37736f
C132 VN.t2 VSUBS 0.907775f
C133 VN.n8 VSUBS 0.399868f
C134 VN.n9 VSUBS 0.013858f
C135 VN.t3 VSUBS 0.907775f
C136 VN.n10 VSUBS 0.388866f
C137 VN.n11 VSUBS 2.14455f
C138 B.n0 VSUBS 0.005317f
C139 B.n1 VSUBS 0.005317f
C140 B.n2 VSUBS 0.007863f
C141 B.n3 VSUBS 0.006025f
C142 B.n4 VSUBS 0.006025f
C143 B.n5 VSUBS 0.006025f
C144 B.n6 VSUBS 0.006025f
C145 B.n7 VSUBS 0.006025f
C146 B.n8 VSUBS 0.006025f
C147 B.n9 VSUBS 0.006025f
C148 B.n10 VSUBS 0.006025f
C149 B.n11 VSUBS 0.01477f
C150 B.n12 VSUBS 0.006025f
C151 B.n13 VSUBS 0.006025f
C152 B.n14 VSUBS 0.006025f
C153 B.n15 VSUBS 0.006025f
C154 B.n16 VSUBS 0.006025f
C155 B.n17 VSUBS 0.006025f
C156 B.n18 VSUBS 0.006025f
C157 B.n19 VSUBS 0.006025f
C158 B.n20 VSUBS 0.006025f
C159 B.n21 VSUBS 0.006025f
C160 B.n22 VSUBS 0.006025f
C161 B.n23 VSUBS 0.006025f
C162 B.n24 VSUBS 0.006025f
C163 B.n25 VSUBS 0.006025f
C164 B.t10 VSUBS 0.105714f
C165 B.t11 VSUBS 0.114557f
C166 B.t9 VSUBS 0.187747f
C167 B.n26 VSUBS 0.185372f
C168 B.n27 VSUBS 0.155701f
C169 B.n28 VSUBS 0.01396f
C170 B.n29 VSUBS 0.006025f
C171 B.n30 VSUBS 0.006025f
C172 B.n31 VSUBS 0.006025f
C173 B.n32 VSUBS 0.006025f
C174 B.n33 VSUBS 0.006025f
C175 B.t1 VSUBS 0.105716f
C176 B.t2 VSUBS 0.114559f
C177 B.t0 VSUBS 0.187747f
C178 B.n34 VSUBS 0.185371f
C179 B.n35 VSUBS 0.155699f
C180 B.n36 VSUBS 0.006025f
C181 B.n37 VSUBS 0.006025f
C182 B.n38 VSUBS 0.006025f
C183 B.n39 VSUBS 0.006025f
C184 B.n40 VSUBS 0.006025f
C185 B.n41 VSUBS 0.006025f
C186 B.n42 VSUBS 0.006025f
C187 B.n43 VSUBS 0.006025f
C188 B.n44 VSUBS 0.006025f
C189 B.n45 VSUBS 0.006025f
C190 B.n46 VSUBS 0.006025f
C191 B.n47 VSUBS 0.006025f
C192 B.n48 VSUBS 0.006025f
C193 B.n49 VSUBS 0.006025f
C194 B.n50 VSUBS 0.01477f
C195 B.n51 VSUBS 0.006025f
C196 B.n52 VSUBS 0.006025f
C197 B.n53 VSUBS 0.006025f
C198 B.n54 VSUBS 0.006025f
C199 B.n55 VSUBS 0.006025f
C200 B.n56 VSUBS 0.006025f
C201 B.n57 VSUBS 0.006025f
C202 B.n58 VSUBS 0.006025f
C203 B.n59 VSUBS 0.006025f
C204 B.n60 VSUBS 0.006025f
C205 B.n61 VSUBS 0.006025f
C206 B.n62 VSUBS 0.006025f
C207 B.n63 VSUBS 0.006025f
C208 B.n64 VSUBS 0.006025f
C209 B.n65 VSUBS 0.006025f
C210 B.n66 VSUBS 0.006025f
C211 B.n67 VSUBS 0.006025f
C212 B.n68 VSUBS 0.006025f
C213 B.n69 VSUBS 0.006025f
C214 B.n70 VSUBS 0.014895f
C215 B.n71 VSUBS 0.006025f
C216 B.n72 VSUBS 0.006025f
C217 B.n73 VSUBS 0.006025f
C218 B.n74 VSUBS 0.006025f
C219 B.n75 VSUBS 0.006025f
C220 B.n76 VSUBS 0.006025f
C221 B.n77 VSUBS 0.006025f
C222 B.n78 VSUBS 0.006025f
C223 B.n79 VSUBS 0.006025f
C224 B.n80 VSUBS 0.006025f
C225 B.n81 VSUBS 0.006025f
C226 B.n82 VSUBS 0.006025f
C227 B.n83 VSUBS 0.006025f
C228 B.n84 VSUBS 0.005671f
C229 B.n85 VSUBS 0.006025f
C230 B.n86 VSUBS 0.006025f
C231 B.n87 VSUBS 0.006025f
C232 B.n88 VSUBS 0.006025f
C233 B.n89 VSUBS 0.006025f
C234 B.t8 VSUBS 0.105714f
C235 B.t7 VSUBS 0.114557f
C236 B.t6 VSUBS 0.187747f
C237 B.n90 VSUBS 0.185372f
C238 B.n91 VSUBS 0.155701f
C239 B.n92 VSUBS 0.006025f
C240 B.n93 VSUBS 0.006025f
C241 B.n94 VSUBS 0.006025f
C242 B.n95 VSUBS 0.006025f
C243 B.n96 VSUBS 0.006025f
C244 B.n97 VSUBS 0.006025f
C245 B.n98 VSUBS 0.006025f
C246 B.n99 VSUBS 0.006025f
C247 B.n100 VSUBS 0.006025f
C248 B.n101 VSUBS 0.006025f
C249 B.n102 VSUBS 0.006025f
C250 B.n103 VSUBS 0.006025f
C251 B.n104 VSUBS 0.006025f
C252 B.n105 VSUBS 0.006025f
C253 B.n106 VSUBS 0.01477f
C254 B.n107 VSUBS 0.006025f
C255 B.n108 VSUBS 0.006025f
C256 B.n109 VSUBS 0.006025f
C257 B.n110 VSUBS 0.006025f
C258 B.n111 VSUBS 0.006025f
C259 B.n112 VSUBS 0.006025f
C260 B.n113 VSUBS 0.006025f
C261 B.n114 VSUBS 0.006025f
C262 B.n115 VSUBS 0.006025f
C263 B.n116 VSUBS 0.006025f
C264 B.n117 VSUBS 0.006025f
C265 B.n118 VSUBS 0.006025f
C266 B.n119 VSUBS 0.006025f
C267 B.n120 VSUBS 0.006025f
C268 B.n121 VSUBS 0.006025f
C269 B.n122 VSUBS 0.006025f
C270 B.n123 VSUBS 0.006025f
C271 B.n124 VSUBS 0.006025f
C272 B.n125 VSUBS 0.006025f
C273 B.n126 VSUBS 0.006025f
C274 B.n127 VSUBS 0.006025f
C275 B.n128 VSUBS 0.006025f
C276 B.n129 VSUBS 0.006025f
C277 B.n130 VSUBS 0.006025f
C278 B.n131 VSUBS 0.006025f
C279 B.n132 VSUBS 0.006025f
C280 B.n133 VSUBS 0.006025f
C281 B.n134 VSUBS 0.006025f
C282 B.n135 VSUBS 0.006025f
C283 B.n136 VSUBS 0.006025f
C284 B.n137 VSUBS 0.006025f
C285 B.n138 VSUBS 0.006025f
C286 B.n139 VSUBS 0.006025f
C287 B.n140 VSUBS 0.006025f
C288 B.n141 VSUBS 0.01477f
C289 B.n142 VSUBS 0.015534f
C290 B.n143 VSUBS 0.015534f
C291 B.n144 VSUBS 0.006025f
C292 B.n145 VSUBS 0.006025f
C293 B.n146 VSUBS 0.006025f
C294 B.n147 VSUBS 0.006025f
C295 B.n148 VSUBS 0.006025f
C296 B.n149 VSUBS 0.006025f
C297 B.n150 VSUBS 0.006025f
C298 B.n151 VSUBS 0.006025f
C299 B.n152 VSUBS 0.006025f
C300 B.n153 VSUBS 0.006025f
C301 B.n154 VSUBS 0.006025f
C302 B.n155 VSUBS 0.006025f
C303 B.n156 VSUBS 0.006025f
C304 B.n157 VSUBS 0.006025f
C305 B.n158 VSUBS 0.006025f
C306 B.n159 VSUBS 0.006025f
C307 B.n160 VSUBS 0.006025f
C308 B.n161 VSUBS 0.006025f
C309 B.n162 VSUBS 0.006025f
C310 B.n163 VSUBS 0.006025f
C311 B.n164 VSUBS 0.006025f
C312 B.n165 VSUBS 0.006025f
C313 B.n166 VSUBS 0.006025f
C314 B.n167 VSUBS 0.006025f
C315 B.n168 VSUBS 0.006025f
C316 B.n169 VSUBS 0.006025f
C317 B.n170 VSUBS 0.006025f
C318 B.n171 VSUBS 0.006025f
C319 B.n172 VSUBS 0.006025f
C320 B.n173 VSUBS 0.006025f
C321 B.n174 VSUBS 0.006025f
C322 B.n175 VSUBS 0.006025f
C323 B.n176 VSUBS 0.006025f
C324 B.n177 VSUBS 0.006025f
C325 B.n178 VSUBS 0.006025f
C326 B.n179 VSUBS 0.006025f
C327 B.n180 VSUBS 0.006025f
C328 B.n181 VSUBS 0.006025f
C329 B.n182 VSUBS 0.006025f
C330 B.n183 VSUBS 0.006025f
C331 B.n184 VSUBS 0.006025f
C332 B.n185 VSUBS 0.005671f
C333 B.n186 VSUBS 0.01396f
C334 B.n187 VSUBS 0.003367f
C335 B.n188 VSUBS 0.006025f
C336 B.n189 VSUBS 0.006025f
C337 B.n190 VSUBS 0.006025f
C338 B.n191 VSUBS 0.006025f
C339 B.n192 VSUBS 0.006025f
C340 B.n193 VSUBS 0.006025f
C341 B.n194 VSUBS 0.006025f
C342 B.n195 VSUBS 0.006025f
C343 B.n196 VSUBS 0.006025f
C344 B.n197 VSUBS 0.006025f
C345 B.n198 VSUBS 0.006025f
C346 B.n199 VSUBS 0.006025f
C347 B.t5 VSUBS 0.105716f
C348 B.t4 VSUBS 0.114559f
C349 B.t3 VSUBS 0.187747f
C350 B.n200 VSUBS 0.185371f
C351 B.n201 VSUBS 0.155699f
C352 B.n202 VSUBS 0.01396f
C353 B.n203 VSUBS 0.003367f
C354 B.n204 VSUBS 0.006025f
C355 B.n205 VSUBS 0.006025f
C356 B.n206 VSUBS 0.006025f
C357 B.n207 VSUBS 0.006025f
C358 B.n208 VSUBS 0.006025f
C359 B.n209 VSUBS 0.006025f
C360 B.n210 VSUBS 0.006025f
C361 B.n211 VSUBS 0.006025f
C362 B.n212 VSUBS 0.006025f
C363 B.n213 VSUBS 0.006025f
C364 B.n214 VSUBS 0.006025f
C365 B.n215 VSUBS 0.006025f
C366 B.n216 VSUBS 0.006025f
C367 B.n217 VSUBS 0.006025f
C368 B.n218 VSUBS 0.006025f
C369 B.n219 VSUBS 0.006025f
C370 B.n220 VSUBS 0.006025f
C371 B.n221 VSUBS 0.006025f
C372 B.n222 VSUBS 0.006025f
C373 B.n223 VSUBS 0.006025f
C374 B.n224 VSUBS 0.006025f
C375 B.n225 VSUBS 0.006025f
C376 B.n226 VSUBS 0.006025f
C377 B.n227 VSUBS 0.006025f
C378 B.n228 VSUBS 0.006025f
C379 B.n229 VSUBS 0.006025f
C380 B.n230 VSUBS 0.006025f
C381 B.n231 VSUBS 0.006025f
C382 B.n232 VSUBS 0.006025f
C383 B.n233 VSUBS 0.006025f
C384 B.n234 VSUBS 0.006025f
C385 B.n235 VSUBS 0.006025f
C386 B.n236 VSUBS 0.006025f
C387 B.n237 VSUBS 0.006025f
C388 B.n238 VSUBS 0.006025f
C389 B.n239 VSUBS 0.006025f
C390 B.n240 VSUBS 0.006025f
C391 B.n241 VSUBS 0.006025f
C392 B.n242 VSUBS 0.006025f
C393 B.n243 VSUBS 0.006025f
C394 B.n244 VSUBS 0.006025f
C395 B.n245 VSUBS 0.006025f
C396 B.n246 VSUBS 0.006025f
C397 B.n247 VSUBS 0.015534f
C398 B.n248 VSUBS 0.01477f
C399 B.n249 VSUBS 0.01541f
C400 B.n250 VSUBS 0.006025f
C401 B.n251 VSUBS 0.006025f
C402 B.n252 VSUBS 0.006025f
C403 B.n253 VSUBS 0.006025f
C404 B.n254 VSUBS 0.006025f
C405 B.n255 VSUBS 0.006025f
C406 B.n256 VSUBS 0.006025f
C407 B.n257 VSUBS 0.006025f
C408 B.n258 VSUBS 0.006025f
C409 B.n259 VSUBS 0.006025f
C410 B.n260 VSUBS 0.006025f
C411 B.n261 VSUBS 0.006025f
C412 B.n262 VSUBS 0.006025f
C413 B.n263 VSUBS 0.006025f
C414 B.n264 VSUBS 0.006025f
C415 B.n265 VSUBS 0.006025f
C416 B.n266 VSUBS 0.006025f
C417 B.n267 VSUBS 0.006025f
C418 B.n268 VSUBS 0.006025f
C419 B.n269 VSUBS 0.006025f
C420 B.n270 VSUBS 0.006025f
C421 B.n271 VSUBS 0.006025f
C422 B.n272 VSUBS 0.006025f
C423 B.n273 VSUBS 0.006025f
C424 B.n274 VSUBS 0.006025f
C425 B.n275 VSUBS 0.006025f
C426 B.n276 VSUBS 0.006025f
C427 B.n277 VSUBS 0.006025f
C428 B.n278 VSUBS 0.006025f
C429 B.n279 VSUBS 0.006025f
C430 B.n280 VSUBS 0.006025f
C431 B.n281 VSUBS 0.006025f
C432 B.n282 VSUBS 0.006025f
C433 B.n283 VSUBS 0.006025f
C434 B.n284 VSUBS 0.006025f
C435 B.n285 VSUBS 0.006025f
C436 B.n286 VSUBS 0.006025f
C437 B.n287 VSUBS 0.006025f
C438 B.n288 VSUBS 0.006025f
C439 B.n289 VSUBS 0.006025f
C440 B.n290 VSUBS 0.006025f
C441 B.n291 VSUBS 0.006025f
C442 B.n292 VSUBS 0.006025f
C443 B.n293 VSUBS 0.006025f
C444 B.n294 VSUBS 0.006025f
C445 B.n295 VSUBS 0.006025f
C446 B.n296 VSUBS 0.006025f
C447 B.n297 VSUBS 0.006025f
C448 B.n298 VSUBS 0.006025f
C449 B.n299 VSUBS 0.006025f
C450 B.n300 VSUBS 0.006025f
C451 B.n301 VSUBS 0.006025f
C452 B.n302 VSUBS 0.006025f
C453 B.n303 VSUBS 0.006025f
C454 B.n304 VSUBS 0.006025f
C455 B.n305 VSUBS 0.006025f
C456 B.n306 VSUBS 0.006025f
C457 B.n307 VSUBS 0.01477f
C458 B.n308 VSUBS 0.015534f
C459 B.n309 VSUBS 0.015534f
C460 B.n310 VSUBS 0.006025f
C461 B.n311 VSUBS 0.006025f
C462 B.n312 VSUBS 0.006025f
C463 B.n313 VSUBS 0.006025f
C464 B.n314 VSUBS 0.006025f
C465 B.n315 VSUBS 0.006025f
C466 B.n316 VSUBS 0.006025f
C467 B.n317 VSUBS 0.006025f
C468 B.n318 VSUBS 0.006025f
C469 B.n319 VSUBS 0.006025f
C470 B.n320 VSUBS 0.006025f
C471 B.n321 VSUBS 0.006025f
C472 B.n322 VSUBS 0.006025f
C473 B.n323 VSUBS 0.006025f
C474 B.n324 VSUBS 0.006025f
C475 B.n325 VSUBS 0.006025f
C476 B.n326 VSUBS 0.006025f
C477 B.n327 VSUBS 0.006025f
C478 B.n328 VSUBS 0.006025f
C479 B.n329 VSUBS 0.006025f
C480 B.n330 VSUBS 0.006025f
C481 B.n331 VSUBS 0.006025f
C482 B.n332 VSUBS 0.006025f
C483 B.n333 VSUBS 0.006025f
C484 B.n334 VSUBS 0.006025f
C485 B.n335 VSUBS 0.006025f
C486 B.n336 VSUBS 0.006025f
C487 B.n337 VSUBS 0.006025f
C488 B.n338 VSUBS 0.006025f
C489 B.n339 VSUBS 0.006025f
C490 B.n340 VSUBS 0.006025f
C491 B.n341 VSUBS 0.006025f
C492 B.n342 VSUBS 0.006025f
C493 B.n343 VSUBS 0.006025f
C494 B.n344 VSUBS 0.006025f
C495 B.n345 VSUBS 0.006025f
C496 B.n346 VSUBS 0.006025f
C497 B.n347 VSUBS 0.006025f
C498 B.n348 VSUBS 0.006025f
C499 B.n349 VSUBS 0.006025f
C500 B.n350 VSUBS 0.006025f
C501 B.n351 VSUBS 0.005671f
C502 B.n352 VSUBS 0.01396f
C503 B.n353 VSUBS 0.003367f
C504 B.n354 VSUBS 0.006025f
C505 B.n355 VSUBS 0.006025f
C506 B.n356 VSUBS 0.006025f
C507 B.n357 VSUBS 0.006025f
C508 B.n358 VSUBS 0.006025f
C509 B.n359 VSUBS 0.006025f
C510 B.n360 VSUBS 0.006025f
C511 B.n361 VSUBS 0.006025f
C512 B.n362 VSUBS 0.006025f
C513 B.n363 VSUBS 0.006025f
C514 B.n364 VSUBS 0.006025f
C515 B.n365 VSUBS 0.006025f
C516 B.n366 VSUBS 0.003367f
C517 B.n367 VSUBS 0.006025f
C518 B.n368 VSUBS 0.006025f
C519 B.n369 VSUBS 0.005671f
C520 B.n370 VSUBS 0.006025f
C521 B.n371 VSUBS 0.006025f
C522 B.n372 VSUBS 0.006025f
C523 B.n373 VSUBS 0.006025f
C524 B.n374 VSUBS 0.006025f
C525 B.n375 VSUBS 0.006025f
C526 B.n376 VSUBS 0.006025f
C527 B.n377 VSUBS 0.006025f
C528 B.n378 VSUBS 0.006025f
C529 B.n379 VSUBS 0.006025f
C530 B.n380 VSUBS 0.006025f
C531 B.n381 VSUBS 0.006025f
C532 B.n382 VSUBS 0.006025f
C533 B.n383 VSUBS 0.006025f
C534 B.n384 VSUBS 0.006025f
C535 B.n385 VSUBS 0.006025f
C536 B.n386 VSUBS 0.006025f
C537 B.n387 VSUBS 0.006025f
C538 B.n388 VSUBS 0.006025f
C539 B.n389 VSUBS 0.006025f
C540 B.n390 VSUBS 0.006025f
C541 B.n391 VSUBS 0.006025f
C542 B.n392 VSUBS 0.006025f
C543 B.n393 VSUBS 0.006025f
C544 B.n394 VSUBS 0.006025f
C545 B.n395 VSUBS 0.006025f
C546 B.n396 VSUBS 0.006025f
C547 B.n397 VSUBS 0.006025f
C548 B.n398 VSUBS 0.006025f
C549 B.n399 VSUBS 0.006025f
C550 B.n400 VSUBS 0.006025f
C551 B.n401 VSUBS 0.006025f
C552 B.n402 VSUBS 0.006025f
C553 B.n403 VSUBS 0.006025f
C554 B.n404 VSUBS 0.006025f
C555 B.n405 VSUBS 0.006025f
C556 B.n406 VSUBS 0.006025f
C557 B.n407 VSUBS 0.006025f
C558 B.n408 VSUBS 0.006025f
C559 B.n409 VSUBS 0.006025f
C560 B.n410 VSUBS 0.015534f
C561 B.n411 VSUBS 0.015534f
C562 B.n412 VSUBS 0.01477f
C563 B.n413 VSUBS 0.006025f
C564 B.n414 VSUBS 0.006025f
C565 B.n415 VSUBS 0.006025f
C566 B.n416 VSUBS 0.006025f
C567 B.n417 VSUBS 0.006025f
C568 B.n418 VSUBS 0.006025f
C569 B.n419 VSUBS 0.006025f
C570 B.n420 VSUBS 0.006025f
C571 B.n421 VSUBS 0.006025f
C572 B.n422 VSUBS 0.006025f
C573 B.n423 VSUBS 0.006025f
C574 B.n424 VSUBS 0.006025f
C575 B.n425 VSUBS 0.006025f
C576 B.n426 VSUBS 0.006025f
C577 B.n427 VSUBS 0.006025f
C578 B.n428 VSUBS 0.006025f
C579 B.n429 VSUBS 0.006025f
C580 B.n430 VSUBS 0.006025f
C581 B.n431 VSUBS 0.006025f
C582 B.n432 VSUBS 0.006025f
C583 B.n433 VSUBS 0.006025f
C584 B.n434 VSUBS 0.006025f
C585 B.n435 VSUBS 0.006025f
C586 B.n436 VSUBS 0.006025f
C587 B.n437 VSUBS 0.006025f
C588 B.n438 VSUBS 0.006025f
C589 B.n439 VSUBS 0.007863f
C590 B.n440 VSUBS 0.008376f
C591 B.n441 VSUBS 0.016656f
C592 VDD1.n0 VSUBS 0.023754f
C593 VDD1.n1 VSUBS 0.023722f
C594 VDD1.n2 VSUBS 0.013122f
C595 VDD1.n3 VSUBS 0.03013f
C596 VDD1.n4 VSUBS 0.012747f
C597 VDD1.n5 VSUBS 0.013497f
C598 VDD1.n6 VSUBS 0.023722f
C599 VDD1.n7 VSUBS 0.012747f
C600 VDD1.n8 VSUBS 0.03013f
C601 VDD1.n9 VSUBS 0.013497f
C602 VDD1.n10 VSUBS 0.023722f
C603 VDD1.n11 VSUBS 0.012747f
C604 VDD1.n12 VSUBS 0.022597f
C605 VDD1.n13 VSUBS 0.022665f
C606 VDD1.t3 VSUBS 0.064669f
C607 VDD1.n14 VSUBS 0.142054f
C608 VDD1.n15 VSUBS 0.730924f
C609 VDD1.n16 VSUBS 0.012747f
C610 VDD1.n17 VSUBS 0.013497f
C611 VDD1.n18 VSUBS 0.03013f
C612 VDD1.n19 VSUBS 0.03013f
C613 VDD1.n20 VSUBS 0.013497f
C614 VDD1.n21 VSUBS 0.012747f
C615 VDD1.n22 VSUBS 0.023722f
C616 VDD1.n23 VSUBS 0.023722f
C617 VDD1.n24 VSUBS 0.012747f
C618 VDD1.n25 VSUBS 0.013497f
C619 VDD1.n26 VSUBS 0.03013f
C620 VDD1.n27 VSUBS 0.03013f
C621 VDD1.n28 VSUBS 0.013497f
C622 VDD1.n29 VSUBS 0.012747f
C623 VDD1.n30 VSUBS 0.023722f
C624 VDD1.n31 VSUBS 0.023722f
C625 VDD1.n32 VSUBS 0.012747f
C626 VDD1.n33 VSUBS 0.013497f
C627 VDD1.n34 VSUBS 0.03013f
C628 VDD1.n35 VSUBS 0.03013f
C629 VDD1.n36 VSUBS 0.065067f
C630 VDD1.n37 VSUBS 0.013122f
C631 VDD1.n38 VSUBS 0.012747f
C632 VDD1.n39 VSUBS 0.05548f
C633 VDD1.n40 VSUBS 0.050156f
C634 VDD1.n41 VSUBS 0.023754f
C635 VDD1.n42 VSUBS 0.023722f
C636 VDD1.n43 VSUBS 0.013122f
C637 VDD1.n44 VSUBS 0.03013f
C638 VDD1.n45 VSUBS 0.013497f
C639 VDD1.n46 VSUBS 0.023722f
C640 VDD1.n47 VSUBS 0.012747f
C641 VDD1.n48 VSUBS 0.03013f
C642 VDD1.n49 VSUBS 0.013497f
C643 VDD1.n50 VSUBS 0.023722f
C644 VDD1.n51 VSUBS 0.012747f
C645 VDD1.n52 VSUBS 0.022597f
C646 VDD1.n53 VSUBS 0.022665f
C647 VDD1.t5 VSUBS 0.064669f
C648 VDD1.n54 VSUBS 0.142054f
C649 VDD1.n55 VSUBS 0.730923f
C650 VDD1.n56 VSUBS 0.012747f
C651 VDD1.n57 VSUBS 0.013497f
C652 VDD1.n58 VSUBS 0.03013f
C653 VDD1.n59 VSUBS 0.03013f
C654 VDD1.n60 VSUBS 0.013497f
C655 VDD1.n61 VSUBS 0.012747f
C656 VDD1.n62 VSUBS 0.023722f
C657 VDD1.n63 VSUBS 0.023722f
C658 VDD1.n64 VSUBS 0.012747f
C659 VDD1.n65 VSUBS 0.013497f
C660 VDD1.n66 VSUBS 0.03013f
C661 VDD1.n67 VSUBS 0.03013f
C662 VDD1.n68 VSUBS 0.013497f
C663 VDD1.n69 VSUBS 0.012747f
C664 VDD1.n70 VSUBS 0.023722f
C665 VDD1.n71 VSUBS 0.023722f
C666 VDD1.n72 VSUBS 0.012747f
C667 VDD1.n73 VSUBS 0.012747f
C668 VDD1.n74 VSUBS 0.013497f
C669 VDD1.n75 VSUBS 0.03013f
C670 VDD1.n76 VSUBS 0.03013f
C671 VDD1.n77 VSUBS 0.065067f
C672 VDD1.n78 VSUBS 0.013122f
C673 VDD1.n79 VSUBS 0.012747f
C674 VDD1.n80 VSUBS 0.05548f
C675 VDD1.n81 VSUBS 0.049842f
C676 VDD1.t4 VSUBS 0.146593f
C677 VDD1.t0 VSUBS 0.146593f
C678 VDD1.n82 VSUBS 1.05373f
C679 VDD1.n83 VSUBS 1.78196f
C680 VDD1.t2 VSUBS 0.146593f
C681 VDD1.t1 VSUBS 0.146593f
C682 VDD1.n84 VSUBS 1.0528f
C683 VDD1.n85 VSUBS 2.02236f
C684 VTAIL.t4 VSUBS 0.174877f
C685 VTAIL.t2 VSUBS 0.174877f
C686 VTAIL.n0 VSUBS 1.13609f
C687 VTAIL.n1 VSUBS 0.667946f
C688 VTAIL.n2 VSUBS 0.028337f
C689 VTAIL.n3 VSUBS 0.028299f
C690 VTAIL.n4 VSUBS 0.015654f
C691 VTAIL.n5 VSUBS 0.035943f
C692 VTAIL.n6 VSUBS 0.016101f
C693 VTAIL.n7 VSUBS 0.028299f
C694 VTAIL.n8 VSUBS 0.015207f
C695 VTAIL.n9 VSUBS 0.035943f
C696 VTAIL.n10 VSUBS 0.016101f
C697 VTAIL.n11 VSUBS 0.028299f
C698 VTAIL.n12 VSUBS 0.015207f
C699 VTAIL.n13 VSUBS 0.026957f
C700 VTAIL.n14 VSUBS 0.027038f
C701 VTAIL.t11 VSUBS 0.077147f
C702 VTAIL.n15 VSUBS 0.169463f
C703 VTAIL.n16 VSUBS 0.87195f
C704 VTAIL.n17 VSUBS 0.015207f
C705 VTAIL.n18 VSUBS 0.016101f
C706 VTAIL.n19 VSUBS 0.035943f
C707 VTAIL.n20 VSUBS 0.035943f
C708 VTAIL.n21 VSUBS 0.016101f
C709 VTAIL.n22 VSUBS 0.015207f
C710 VTAIL.n23 VSUBS 0.028299f
C711 VTAIL.n24 VSUBS 0.028299f
C712 VTAIL.n25 VSUBS 0.015207f
C713 VTAIL.n26 VSUBS 0.016101f
C714 VTAIL.n27 VSUBS 0.035943f
C715 VTAIL.n28 VSUBS 0.035943f
C716 VTAIL.n29 VSUBS 0.016101f
C717 VTAIL.n30 VSUBS 0.015207f
C718 VTAIL.n31 VSUBS 0.028299f
C719 VTAIL.n32 VSUBS 0.028299f
C720 VTAIL.n33 VSUBS 0.015207f
C721 VTAIL.n34 VSUBS 0.015207f
C722 VTAIL.n35 VSUBS 0.016101f
C723 VTAIL.n36 VSUBS 0.035943f
C724 VTAIL.n37 VSUBS 0.035943f
C725 VTAIL.n38 VSUBS 0.077622f
C726 VTAIL.n39 VSUBS 0.015654f
C727 VTAIL.n40 VSUBS 0.015207f
C728 VTAIL.n41 VSUBS 0.066185f
C729 VTAIL.n42 VSUBS 0.038642f
C730 VTAIL.n43 VSUBS 0.184181f
C731 VTAIL.t9 VSUBS 0.174877f
C732 VTAIL.t10 VSUBS 0.174877f
C733 VTAIL.n44 VSUBS 1.13609f
C734 VTAIL.n45 VSUBS 1.79403f
C735 VTAIL.t5 VSUBS 0.174877f
C736 VTAIL.t0 VSUBS 0.174877f
C737 VTAIL.n46 VSUBS 1.1361f
C738 VTAIL.n47 VSUBS 1.79402f
C739 VTAIL.n48 VSUBS 0.028337f
C740 VTAIL.n49 VSUBS 0.028299f
C741 VTAIL.n50 VSUBS 0.015654f
C742 VTAIL.n51 VSUBS 0.035943f
C743 VTAIL.n52 VSUBS 0.015207f
C744 VTAIL.n53 VSUBS 0.016101f
C745 VTAIL.n54 VSUBS 0.028299f
C746 VTAIL.n55 VSUBS 0.015207f
C747 VTAIL.n56 VSUBS 0.035943f
C748 VTAIL.n57 VSUBS 0.016101f
C749 VTAIL.n58 VSUBS 0.028299f
C750 VTAIL.n59 VSUBS 0.015207f
C751 VTAIL.n60 VSUBS 0.026957f
C752 VTAIL.n61 VSUBS 0.027038f
C753 VTAIL.t1 VSUBS 0.077147f
C754 VTAIL.n62 VSUBS 0.169463f
C755 VTAIL.n63 VSUBS 0.87195f
C756 VTAIL.n64 VSUBS 0.015207f
C757 VTAIL.n65 VSUBS 0.016101f
C758 VTAIL.n66 VSUBS 0.035943f
C759 VTAIL.n67 VSUBS 0.035943f
C760 VTAIL.n68 VSUBS 0.016101f
C761 VTAIL.n69 VSUBS 0.015207f
C762 VTAIL.n70 VSUBS 0.028299f
C763 VTAIL.n71 VSUBS 0.028299f
C764 VTAIL.n72 VSUBS 0.015207f
C765 VTAIL.n73 VSUBS 0.016101f
C766 VTAIL.n74 VSUBS 0.035943f
C767 VTAIL.n75 VSUBS 0.035943f
C768 VTAIL.n76 VSUBS 0.016101f
C769 VTAIL.n77 VSUBS 0.015207f
C770 VTAIL.n78 VSUBS 0.028299f
C771 VTAIL.n79 VSUBS 0.028299f
C772 VTAIL.n80 VSUBS 0.015207f
C773 VTAIL.n81 VSUBS 0.016101f
C774 VTAIL.n82 VSUBS 0.035943f
C775 VTAIL.n83 VSUBS 0.035943f
C776 VTAIL.n84 VSUBS 0.077622f
C777 VTAIL.n85 VSUBS 0.015654f
C778 VTAIL.n86 VSUBS 0.015207f
C779 VTAIL.n87 VSUBS 0.066185f
C780 VTAIL.n88 VSUBS 0.038642f
C781 VTAIL.n89 VSUBS 0.184181f
C782 VTAIL.t7 VSUBS 0.174877f
C783 VTAIL.t8 VSUBS 0.174877f
C784 VTAIL.n90 VSUBS 1.1361f
C785 VTAIL.n91 VSUBS 0.720998f
C786 VTAIL.n92 VSUBS 0.028337f
C787 VTAIL.n93 VSUBS 0.028299f
C788 VTAIL.n94 VSUBS 0.015654f
C789 VTAIL.n95 VSUBS 0.035943f
C790 VTAIL.n96 VSUBS 0.015207f
C791 VTAIL.n97 VSUBS 0.016101f
C792 VTAIL.n98 VSUBS 0.028299f
C793 VTAIL.n99 VSUBS 0.015207f
C794 VTAIL.n100 VSUBS 0.035943f
C795 VTAIL.n101 VSUBS 0.016101f
C796 VTAIL.n102 VSUBS 0.028299f
C797 VTAIL.n103 VSUBS 0.015207f
C798 VTAIL.n104 VSUBS 0.026957f
C799 VTAIL.n105 VSUBS 0.027038f
C800 VTAIL.t6 VSUBS 0.077147f
C801 VTAIL.n106 VSUBS 0.169463f
C802 VTAIL.n107 VSUBS 0.87195f
C803 VTAIL.n108 VSUBS 0.015207f
C804 VTAIL.n109 VSUBS 0.016101f
C805 VTAIL.n110 VSUBS 0.035943f
C806 VTAIL.n111 VSUBS 0.035943f
C807 VTAIL.n112 VSUBS 0.016101f
C808 VTAIL.n113 VSUBS 0.015207f
C809 VTAIL.n114 VSUBS 0.028299f
C810 VTAIL.n115 VSUBS 0.028299f
C811 VTAIL.n116 VSUBS 0.015207f
C812 VTAIL.n117 VSUBS 0.016101f
C813 VTAIL.n118 VSUBS 0.035943f
C814 VTAIL.n119 VSUBS 0.035943f
C815 VTAIL.n120 VSUBS 0.016101f
C816 VTAIL.n121 VSUBS 0.015207f
C817 VTAIL.n122 VSUBS 0.028299f
C818 VTAIL.n123 VSUBS 0.028299f
C819 VTAIL.n124 VSUBS 0.015207f
C820 VTAIL.n125 VSUBS 0.016101f
C821 VTAIL.n126 VSUBS 0.035943f
C822 VTAIL.n127 VSUBS 0.035943f
C823 VTAIL.n128 VSUBS 0.077622f
C824 VTAIL.n129 VSUBS 0.015654f
C825 VTAIL.n130 VSUBS 0.015207f
C826 VTAIL.n131 VSUBS 0.066185f
C827 VTAIL.n132 VSUBS 0.038642f
C828 VTAIL.n133 VSUBS 1.17938f
C829 VTAIL.n134 VSUBS 0.028337f
C830 VTAIL.n135 VSUBS 0.028299f
C831 VTAIL.n136 VSUBS 0.015654f
C832 VTAIL.n137 VSUBS 0.035943f
C833 VTAIL.n138 VSUBS 0.016101f
C834 VTAIL.n139 VSUBS 0.028299f
C835 VTAIL.n140 VSUBS 0.015207f
C836 VTAIL.n141 VSUBS 0.035943f
C837 VTAIL.n142 VSUBS 0.016101f
C838 VTAIL.n143 VSUBS 0.028299f
C839 VTAIL.n144 VSUBS 0.015207f
C840 VTAIL.n145 VSUBS 0.026957f
C841 VTAIL.n146 VSUBS 0.027038f
C842 VTAIL.t3 VSUBS 0.077147f
C843 VTAIL.n147 VSUBS 0.169463f
C844 VTAIL.n148 VSUBS 0.87195f
C845 VTAIL.n149 VSUBS 0.015207f
C846 VTAIL.n150 VSUBS 0.016101f
C847 VTAIL.n151 VSUBS 0.035943f
C848 VTAIL.n152 VSUBS 0.035943f
C849 VTAIL.n153 VSUBS 0.016101f
C850 VTAIL.n154 VSUBS 0.015207f
C851 VTAIL.n155 VSUBS 0.028299f
C852 VTAIL.n156 VSUBS 0.028299f
C853 VTAIL.n157 VSUBS 0.015207f
C854 VTAIL.n158 VSUBS 0.016101f
C855 VTAIL.n159 VSUBS 0.035943f
C856 VTAIL.n160 VSUBS 0.035943f
C857 VTAIL.n161 VSUBS 0.016101f
C858 VTAIL.n162 VSUBS 0.015207f
C859 VTAIL.n163 VSUBS 0.028299f
C860 VTAIL.n164 VSUBS 0.028299f
C861 VTAIL.n165 VSUBS 0.015207f
C862 VTAIL.n166 VSUBS 0.015207f
C863 VTAIL.n167 VSUBS 0.016101f
C864 VTAIL.n168 VSUBS 0.035943f
C865 VTAIL.n169 VSUBS 0.035943f
C866 VTAIL.n170 VSUBS 0.077622f
C867 VTAIL.n171 VSUBS 0.015654f
C868 VTAIL.n172 VSUBS 0.015207f
C869 VTAIL.n173 VSUBS 0.066185f
C870 VTAIL.n174 VSUBS 0.038642f
C871 VTAIL.n175 VSUBS 1.15462f
C872 VP.n0 VSUBS 0.062936f
C873 VP.n1 VSUBS 0.014282f
C874 VP.n2 VSUBS 0.25595f
C875 VP.t4 VSUBS 0.935542f
C876 VP.t3 VSUBS 0.935542f
C877 VP.t2 VSUBS 0.958555f
C878 VP.n3 VSUBS 0.388903f
C879 VP.n4 VSUBS 0.412099f
C880 VP.n5 VSUBS 0.014282f
C881 VP.n6 VSUBS 0.40076f
C882 VP.n7 VSUBS 2.16855f
C883 VP.t0 VSUBS 0.935542f
C884 VP.n8 VSUBS 0.40076f
C885 VP.n9 VSUBS 2.22817f
C886 VP.n10 VSUBS 0.062936f
C887 VP.n11 VSUBS 0.062936f
C888 VP.t1 VSUBS 0.935542f
C889 VP.n12 VSUBS 0.407745f
C890 VP.n13 VSUBS 0.014282f
C891 VP.t5 VSUBS 0.935542f
C892 VP.n14 VSUBS 0.40076f
C893 VP.n15 VSUBS 0.048773f
.ends

