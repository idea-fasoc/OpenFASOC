* NGSPICE file created from diff_pair_sample_1200.ext - technology: sky130A

.subckt diff_pair_sample_1200 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0 ps=0 w=4.3 l=3.92
X1 VDD1.t5 VP.t0 VTAIL.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0.7095 ps=4.63 w=4.3 l=3.92
X2 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0 ps=0 w=4.3 l=3.92
X3 VDD2.t5 VN.t0 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0.7095 ps=4.63 w=4.3 l=3.92
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0 ps=0 w=4.3 l=3.92
X5 VTAIL.t9 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=0.7095 ps=4.63 w=4.3 l=3.92
X6 VTAIL.t3 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=0.7095 ps=4.63 w=4.3 l=3.92
X7 VDD2.t3 VN.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=1.677 ps=9.38 w=4.3 l=3.92
X8 VDD2.t2 VN.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0.7095 ps=4.63 w=4.3 l=3.92
X9 VDD1.t3 VP.t2 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=1.677 ps=9.38 w=4.3 l=3.92
X10 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0 ps=0 w=4.3 l=3.92
X11 VTAIL.t5 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=0.7095 ps=4.63 w=4.3 l=3.92
X12 VDD2.t1 VN.t4 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=1.677 ps=9.38 w=4.3 l=3.92
X13 VDD1.t1 VP.t4 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.677 pd=9.38 as=0.7095 ps=4.63 w=4.3 l=3.92
X14 VDD1.t0 VP.t5 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=1.677 ps=9.38 w=4.3 l=3.92
X15 VTAIL.t11 VN.t5 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7095 pd=4.63 as=0.7095 ps=4.63 w=4.3 l=3.92
R0 B.n623 B.n622 585
R1 B.n625 B.n135 585
R2 B.n628 B.n627 585
R3 B.n629 B.n134 585
R4 B.n631 B.n630 585
R5 B.n633 B.n133 585
R6 B.n636 B.n635 585
R7 B.n637 B.n132 585
R8 B.n639 B.n638 585
R9 B.n641 B.n131 585
R10 B.n644 B.n643 585
R11 B.n645 B.n130 585
R12 B.n647 B.n646 585
R13 B.n649 B.n129 585
R14 B.n652 B.n651 585
R15 B.n653 B.n128 585
R16 B.n655 B.n654 585
R17 B.n657 B.n127 585
R18 B.n660 B.n659 585
R19 B.n662 B.n124 585
R20 B.n664 B.n663 585
R21 B.n666 B.n123 585
R22 B.n669 B.n668 585
R23 B.n670 B.n122 585
R24 B.n672 B.n671 585
R25 B.n674 B.n121 585
R26 B.n677 B.n676 585
R27 B.n678 B.n117 585
R28 B.n680 B.n679 585
R29 B.n682 B.n116 585
R30 B.n685 B.n684 585
R31 B.n686 B.n115 585
R32 B.n688 B.n687 585
R33 B.n690 B.n114 585
R34 B.n693 B.n692 585
R35 B.n694 B.n113 585
R36 B.n696 B.n695 585
R37 B.n698 B.n112 585
R38 B.n701 B.n700 585
R39 B.n702 B.n111 585
R40 B.n704 B.n703 585
R41 B.n706 B.n110 585
R42 B.n709 B.n708 585
R43 B.n710 B.n109 585
R44 B.n712 B.n711 585
R45 B.n714 B.n108 585
R46 B.n717 B.n716 585
R47 B.n718 B.n107 585
R48 B.n621 B.n105 585
R49 B.n721 B.n105 585
R50 B.n620 B.n104 585
R51 B.n722 B.n104 585
R52 B.n619 B.n103 585
R53 B.n723 B.n103 585
R54 B.n618 B.n617 585
R55 B.n617 B.n99 585
R56 B.n616 B.n98 585
R57 B.n729 B.n98 585
R58 B.n615 B.n97 585
R59 B.n730 B.n97 585
R60 B.n614 B.n96 585
R61 B.n731 B.n96 585
R62 B.n613 B.n612 585
R63 B.n612 B.n92 585
R64 B.n611 B.n91 585
R65 B.n737 B.n91 585
R66 B.n610 B.n90 585
R67 B.n738 B.n90 585
R68 B.n609 B.n89 585
R69 B.n739 B.n89 585
R70 B.n608 B.n607 585
R71 B.n607 B.n85 585
R72 B.n606 B.n84 585
R73 B.n745 B.n84 585
R74 B.n605 B.n83 585
R75 B.n746 B.n83 585
R76 B.n604 B.n82 585
R77 B.n747 B.n82 585
R78 B.n603 B.n602 585
R79 B.n602 B.n78 585
R80 B.n601 B.n77 585
R81 B.n753 B.n77 585
R82 B.n600 B.n76 585
R83 B.n754 B.n76 585
R84 B.n599 B.n75 585
R85 B.n755 B.n75 585
R86 B.n598 B.n597 585
R87 B.n597 B.n71 585
R88 B.n596 B.n70 585
R89 B.n761 B.n70 585
R90 B.n595 B.n69 585
R91 B.n762 B.n69 585
R92 B.n594 B.n68 585
R93 B.n763 B.n68 585
R94 B.n593 B.n592 585
R95 B.n592 B.n64 585
R96 B.n591 B.n63 585
R97 B.n769 B.n63 585
R98 B.n590 B.n62 585
R99 B.n770 B.n62 585
R100 B.n589 B.n61 585
R101 B.n771 B.n61 585
R102 B.n588 B.n587 585
R103 B.n587 B.n57 585
R104 B.n586 B.n56 585
R105 B.n777 B.n56 585
R106 B.n585 B.n55 585
R107 B.n778 B.n55 585
R108 B.n584 B.n54 585
R109 B.n779 B.n54 585
R110 B.n583 B.n582 585
R111 B.n582 B.n50 585
R112 B.n581 B.n49 585
R113 B.n785 B.n49 585
R114 B.n580 B.n48 585
R115 B.n786 B.n48 585
R116 B.n579 B.n47 585
R117 B.n787 B.n47 585
R118 B.n578 B.n577 585
R119 B.n577 B.n43 585
R120 B.n576 B.n42 585
R121 B.n793 B.n42 585
R122 B.n575 B.n41 585
R123 B.n794 B.n41 585
R124 B.n574 B.n40 585
R125 B.n795 B.n40 585
R126 B.n573 B.n572 585
R127 B.n572 B.n36 585
R128 B.n571 B.n35 585
R129 B.n801 B.n35 585
R130 B.n570 B.n34 585
R131 B.n802 B.n34 585
R132 B.n569 B.n33 585
R133 B.n803 B.n33 585
R134 B.n568 B.n567 585
R135 B.n567 B.n29 585
R136 B.n566 B.n28 585
R137 B.n809 B.n28 585
R138 B.n565 B.n27 585
R139 B.n810 B.n27 585
R140 B.n564 B.n26 585
R141 B.n811 B.n26 585
R142 B.n563 B.n562 585
R143 B.n562 B.n22 585
R144 B.n561 B.n21 585
R145 B.n817 B.n21 585
R146 B.n560 B.n20 585
R147 B.n818 B.n20 585
R148 B.n559 B.n19 585
R149 B.n819 B.n19 585
R150 B.n558 B.n557 585
R151 B.n557 B.n15 585
R152 B.n556 B.n14 585
R153 B.n825 B.n14 585
R154 B.n555 B.n13 585
R155 B.n826 B.n13 585
R156 B.n554 B.n12 585
R157 B.n827 B.n12 585
R158 B.n553 B.n552 585
R159 B.n552 B.n8 585
R160 B.n551 B.n7 585
R161 B.n833 B.n7 585
R162 B.n550 B.n6 585
R163 B.n834 B.n6 585
R164 B.n549 B.n5 585
R165 B.n835 B.n5 585
R166 B.n548 B.n547 585
R167 B.n547 B.n4 585
R168 B.n546 B.n136 585
R169 B.n546 B.n545 585
R170 B.n536 B.n137 585
R171 B.n138 B.n137 585
R172 B.n538 B.n537 585
R173 B.n539 B.n538 585
R174 B.n535 B.n143 585
R175 B.n143 B.n142 585
R176 B.n534 B.n533 585
R177 B.n533 B.n532 585
R178 B.n145 B.n144 585
R179 B.n146 B.n145 585
R180 B.n525 B.n524 585
R181 B.n526 B.n525 585
R182 B.n523 B.n151 585
R183 B.n151 B.n150 585
R184 B.n522 B.n521 585
R185 B.n521 B.n520 585
R186 B.n153 B.n152 585
R187 B.n154 B.n153 585
R188 B.n513 B.n512 585
R189 B.n514 B.n513 585
R190 B.n511 B.n159 585
R191 B.n159 B.n158 585
R192 B.n510 B.n509 585
R193 B.n509 B.n508 585
R194 B.n161 B.n160 585
R195 B.n162 B.n161 585
R196 B.n501 B.n500 585
R197 B.n502 B.n501 585
R198 B.n499 B.n167 585
R199 B.n167 B.n166 585
R200 B.n498 B.n497 585
R201 B.n497 B.n496 585
R202 B.n169 B.n168 585
R203 B.n170 B.n169 585
R204 B.n489 B.n488 585
R205 B.n490 B.n489 585
R206 B.n487 B.n174 585
R207 B.n178 B.n174 585
R208 B.n486 B.n485 585
R209 B.n485 B.n484 585
R210 B.n176 B.n175 585
R211 B.n177 B.n176 585
R212 B.n477 B.n476 585
R213 B.n478 B.n477 585
R214 B.n475 B.n183 585
R215 B.n183 B.n182 585
R216 B.n474 B.n473 585
R217 B.n473 B.n472 585
R218 B.n185 B.n184 585
R219 B.n186 B.n185 585
R220 B.n465 B.n464 585
R221 B.n466 B.n465 585
R222 B.n463 B.n191 585
R223 B.n191 B.n190 585
R224 B.n462 B.n461 585
R225 B.n461 B.n460 585
R226 B.n193 B.n192 585
R227 B.n194 B.n193 585
R228 B.n453 B.n452 585
R229 B.n454 B.n453 585
R230 B.n451 B.n198 585
R231 B.n202 B.n198 585
R232 B.n450 B.n449 585
R233 B.n449 B.n448 585
R234 B.n200 B.n199 585
R235 B.n201 B.n200 585
R236 B.n441 B.n440 585
R237 B.n442 B.n441 585
R238 B.n439 B.n207 585
R239 B.n207 B.n206 585
R240 B.n438 B.n437 585
R241 B.n437 B.n436 585
R242 B.n209 B.n208 585
R243 B.n210 B.n209 585
R244 B.n429 B.n428 585
R245 B.n430 B.n429 585
R246 B.n427 B.n215 585
R247 B.n215 B.n214 585
R248 B.n426 B.n425 585
R249 B.n425 B.n424 585
R250 B.n217 B.n216 585
R251 B.n218 B.n217 585
R252 B.n417 B.n416 585
R253 B.n418 B.n417 585
R254 B.n415 B.n223 585
R255 B.n223 B.n222 585
R256 B.n414 B.n413 585
R257 B.n413 B.n412 585
R258 B.n225 B.n224 585
R259 B.n226 B.n225 585
R260 B.n405 B.n404 585
R261 B.n406 B.n405 585
R262 B.n403 B.n230 585
R263 B.n234 B.n230 585
R264 B.n402 B.n401 585
R265 B.n401 B.n400 585
R266 B.n232 B.n231 585
R267 B.n233 B.n232 585
R268 B.n393 B.n392 585
R269 B.n394 B.n393 585
R270 B.n391 B.n239 585
R271 B.n239 B.n238 585
R272 B.n390 B.n389 585
R273 B.n389 B.n388 585
R274 B.n241 B.n240 585
R275 B.n242 B.n241 585
R276 B.n381 B.n380 585
R277 B.n382 B.n381 585
R278 B.n379 B.n247 585
R279 B.n247 B.n246 585
R280 B.n378 B.n377 585
R281 B.n377 B.n376 585
R282 B.n373 B.n251 585
R283 B.n372 B.n371 585
R284 B.n369 B.n252 585
R285 B.n369 B.n250 585
R286 B.n368 B.n367 585
R287 B.n366 B.n365 585
R288 B.n364 B.n254 585
R289 B.n362 B.n361 585
R290 B.n360 B.n255 585
R291 B.n359 B.n358 585
R292 B.n356 B.n256 585
R293 B.n354 B.n353 585
R294 B.n352 B.n257 585
R295 B.n351 B.n350 585
R296 B.n348 B.n258 585
R297 B.n346 B.n345 585
R298 B.n344 B.n259 585
R299 B.n343 B.n342 585
R300 B.n340 B.n260 585
R301 B.n338 B.n337 585
R302 B.n335 B.n261 585
R303 B.n334 B.n333 585
R304 B.n331 B.n264 585
R305 B.n329 B.n328 585
R306 B.n327 B.n265 585
R307 B.n326 B.n325 585
R308 B.n323 B.n266 585
R309 B.n321 B.n320 585
R310 B.n319 B.n267 585
R311 B.n318 B.n317 585
R312 B.n315 B.n314 585
R313 B.n313 B.n312 585
R314 B.n311 B.n272 585
R315 B.n309 B.n308 585
R316 B.n307 B.n273 585
R317 B.n306 B.n305 585
R318 B.n303 B.n274 585
R319 B.n301 B.n300 585
R320 B.n299 B.n275 585
R321 B.n298 B.n297 585
R322 B.n295 B.n276 585
R323 B.n293 B.n292 585
R324 B.n291 B.n277 585
R325 B.n290 B.n289 585
R326 B.n287 B.n278 585
R327 B.n285 B.n284 585
R328 B.n283 B.n279 585
R329 B.n282 B.n281 585
R330 B.n249 B.n248 585
R331 B.n250 B.n249 585
R332 B.n375 B.n374 585
R333 B.n376 B.n375 585
R334 B.n245 B.n244 585
R335 B.n246 B.n245 585
R336 B.n384 B.n383 585
R337 B.n383 B.n382 585
R338 B.n385 B.n243 585
R339 B.n243 B.n242 585
R340 B.n387 B.n386 585
R341 B.n388 B.n387 585
R342 B.n237 B.n236 585
R343 B.n238 B.n237 585
R344 B.n396 B.n395 585
R345 B.n395 B.n394 585
R346 B.n397 B.n235 585
R347 B.n235 B.n233 585
R348 B.n399 B.n398 585
R349 B.n400 B.n399 585
R350 B.n229 B.n228 585
R351 B.n234 B.n229 585
R352 B.n408 B.n407 585
R353 B.n407 B.n406 585
R354 B.n409 B.n227 585
R355 B.n227 B.n226 585
R356 B.n411 B.n410 585
R357 B.n412 B.n411 585
R358 B.n221 B.n220 585
R359 B.n222 B.n221 585
R360 B.n420 B.n419 585
R361 B.n419 B.n418 585
R362 B.n421 B.n219 585
R363 B.n219 B.n218 585
R364 B.n423 B.n422 585
R365 B.n424 B.n423 585
R366 B.n213 B.n212 585
R367 B.n214 B.n213 585
R368 B.n432 B.n431 585
R369 B.n431 B.n430 585
R370 B.n433 B.n211 585
R371 B.n211 B.n210 585
R372 B.n435 B.n434 585
R373 B.n436 B.n435 585
R374 B.n205 B.n204 585
R375 B.n206 B.n205 585
R376 B.n444 B.n443 585
R377 B.n443 B.n442 585
R378 B.n445 B.n203 585
R379 B.n203 B.n201 585
R380 B.n447 B.n446 585
R381 B.n448 B.n447 585
R382 B.n197 B.n196 585
R383 B.n202 B.n197 585
R384 B.n456 B.n455 585
R385 B.n455 B.n454 585
R386 B.n457 B.n195 585
R387 B.n195 B.n194 585
R388 B.n459 B.n458 585
R389 B.n460 B.n459 585
R390 B.n189 B.n188 585
R391 B.n190 B.n189 585
R392 B.n468 B.n467 585
R393 B.n467 B.n466 585
R394 B.n469 B.n187 585
R395 B.n187 B.n186 585
R396 B.n471 B.n470 585
R397 B.n472 B.n471 585
R398 B.n181 B.n180 585
R399 B.n182 B.n181 585
R400 B.n480 B.n479 585
R401 B.n479 B.n478 585
R402 B.n481 B.n179 585
R403 B.n179 B.n177 585
R404 B.n483 B.n482 585
R405 B.n484 B.n483 585
R406 B.n173 B.n172 585
R407 B.n178 B.n173 585
R408 B.n492 B.n491 585
R409 B.n491 B.n490 585
R410 B.n493 B.n171 585
R411 B.n171 B.n170 585
R412 B.n495 B.n494 585
R413 B.n496 B.n495 585
R414 B.n165 B.n164 585
R415 B.n166 B.n165 585
R416 B.n504 B.n503 585
R417 B.n503 B.n502 585
R418 B.n505 B.n163 585
R419 B.n163 B.n162 585
R420 B.n507 B.n506 585
R421 B.n508 B.n507 585
R422 B.n157 B.n156 585
R423 B.n158 B.n157 585
R424 B.n516 B.n515 585
R425 B.n515 B.n514 585
R426 B.n517 B.n155 585
R427 B.n155 B.n154 585
R428 B.n519 B.n518 585
R429 B.n520 B.n519 585
R430 B.n149 B.n148 585
R431 B.n150 B.n149 585
R432 B.n528 B.n527 585
R433 B.n527 B.n526 585
R434 B.n529 B.n147 585
R435 B.n147 B.n146 585
R436 B.n531 B.n530 585
R437 B.n532 B.n531 585
R438 B.n141 B.n140 585
R439 B.n142 B.n141 585
R440 B.n541 B.n540 585
R441 B.n540 B.n539 585
R442 B.n542 B.n139 585
R443 B.n139 B.n138 585
R444 B.n544 B.n543 585
R445 B.n545 B.n544 585
R446 B.n2 B.n0 585
R447 B.n4 B.n2 585
R448 B.n3 B.n1 585
R449 B.n834 B.n3 585
R450 B.n832 B.n831 585
R451 B.n833 B.n832 585
R452 B.n830 B.n9 585
R453 B.n9 B.n8 585
R454 B.n829 B.n828 585
R455 B.n828 B.n827 585
R456 B.n11 B.n10 585
R457 B.n826 B.n11 585
R458 B.n824 B.n823 585
R459 B.n825 B.n824 585
R460 B.n822 B.n16 585
R461 B.n16 B.n15 585
R462 B.n821 B.n820 585
R463 B.n820 B.n819 585
R464 B.n18 B.n17 585
R465 B.n818 B.n18 585
R466 B.n816 B.n815 585
R467 B.n817 B.n816 585
R468 B.n814 B.n23 585
R469 B.n23 B.n22 585
R470 B.n813 B.n812 585
R471 B.n812 B.n811 585
R472 B.n25 B.n24 585
R473 B.n810 B.n25 585
R474 B.n808 B.n807 585
R475 B.n809 B.n808 585
R476 B.n806 B.n30 585
R477 B.n30 B.n29 585
R478 B.n805 B.n804 585
R479 B.n804 B.n803 585
R480 B.n32 B.n31 585
R481 B.n802 B.n32 585
R482 B.n800 B.n799 585
R483 B.n801 B.n800 585
R484 B.n798 B.n37 585
R485 B.n37 B.n36 585
R486 B.n797 B.n796 585
R487 B.n796 B.n795 585
R488 B.n39 B.n38 585
R489 B.n794 B.n39 585
R490 B.n792 B.n791 585
R491 B.n793 B.n792 585
R492 B.n790 B.n44 585
R493 B.n44 B.n43 585
R494 B.n789 B.n788 585
R495 B.n788 B.n787 585
R496 B.n46 B.n45 585
R497 B.n786 B.n46 585
R498 B.n784 B.n783 585
R499 B.n785 B.n784 585
R500 B.n782 B.n51 585
R501 B.n51 B.n50 585
R502 B.n781 B.n780 585
R503 B.n780 B.n779 585
R504 B.n53 B.n52 585
R505 B.n778 B.n53 585
R506 B.n776 B.n775 585
R507 B.n777 B.n776 585
R508 B.n774 B.n58 585
R509 B.n58 B.n57 585
R510 B.n773 B.n772 585
R511 B.n772 B.n771 585
R512 B.n60 B.n59 585
R513 B.n770 B.n60 585
R514 B.n768 B.n767 585
R515 B.n769 B.n768 585
R516 B.n766 B.n65 585
R517 B.n65 B.n64 585
R518 B.n765 B.n764 585
R519 B.n764 B.n763 585
R520 B.n67 B.n66 585
R521 B.n762 B.n67 585
R522 B.n760 B.n759 585
R523 B.n761 B.n760 585
R524 B.n758 B.n72 585
R525 B.n72 B.n71 585
R526 B.n757 B.n756 585
R527 B.n756 B.n755 585
R528 B.n74 B.n73 585
R529 B.n754 B.n74 585
R530 B.n752 B.n751 585
R531 B.n753 B.n752 585
R532 B.n750 B.n79 585
R533 B.n79 B.n78 585
R534 B.n749 B.n748 585
R535 B.n748 B.n747 585
R536 B.n81 B.n80 585
R537 B.n746 B.n81 585
R538 B.n744 B.n743 585
R539 B.n745 B.n744 585
R540 B.n742 B.n86 585
R541 B.n86 B.n85 585
R542 B.n741 B.n740 585
R543 B.n740 B.n739 585
R544 B.n88 B.n87 585
R545 B.n738 B.n88 585
R546 B.n736 B.n735 585
R547 B.n737 B.n736 585
R548 B.n734 B.n93 585
R549 B.n93 B.n92 585
R550 B.n733 B.n732 585
R551 B.n732 B.n731 585
R552 B.n95 B.n94 585
R553 B.n730 B.n95 585
R554 B.n728 B.n727 585
R555 B.n729 B.n728 585
R556 B.n726 B.n100 585
R557 B.n100 B.n99 585
R558 B.n725 B.n724 585
R559 B.n724 B.n723 585
R560 B.n102 B.n101 585
R561 B.n722 B.n102 585
R562 B.n720 B.n719 585
R563 B.n721 B.n720 585
R564 B.n837 B.n836 585
R565 B.n836 B.n835 585
R566 B.n375 B.n251 478.086
R567 B.n720 B.n107 478.086
R568 B.n377 B.n249 478.086
R569 B.n623 B.n105 478.086
R570 B.n624 B.n106 256.663
R571 B.n626 B.n106 256.663
R572 B.n632 B.n106 256.663
R573 B.n634 B.n106 256.663
R574 B.n640 B.n106 256.663
R575 B.n642 B.n106 256.663
R576 B.n648 B.n106 256.663
R577 B.n650 B.n106 256.663
R578 B.n656 B.n106 256.663
R579 B.n658 B.n106 256.663
R580 B.n665 B.n106 256.663
R581 B.n667 B.n106 256.663
R582 B.n673 B.n106 256.663
R583 B.n675 B.n106 256.663
R584 B.n681 B.n106 256.663
R585 B.n683 B.n106 256.663
R586 B.n689 B.n106 256.663
R587 B.n691 B.n106 256.663
R588 B.n697 B.n106 256.663
R589 B.n699 B.n106 256.663
R590 B.n705 B.n106 256.663
R591 B.n707 B.n106 256.663
R592 B.n713 B.n106 256.663
R593 B.n715 B.n106 256.663
R594 B.n370 B.n250 256.663
R595 B.n253 B.n250 256.663
R596 B.n363 B.n250 256.663
R597 B.n357 B.n250 256.663
R598 B.n355 B.n250 256.663
R599 B.n349 B.n250 256.663
R600 B.n347 B.n250 256.663
R601 B.n341 B.n250 256.663
R602 B.n339 B.n250 256.663
R603 B.n332 B.n250 256.663
R604 B.n330 B.n250 256.663
R605 B.n324 B.n250 256.663
R606 B.n322 B.n250 256.663
R607 B.n316 B.n250 256.663
R608 B.n271 B.n250 256.663
R609 B.n310 B.n250 256.663
R610 B.n304 B.n250 256.663
R611 B.n302 B.n250 256.663
R612 B.n296 B.n250 256.663
R613 B.n294 B.n250 256.663
R614 B.n288 B.n250 256.663
R615 B.n286 B.n250 256.663
R616 B.n280 B.n250 256.663
R617 B.n268 B.t17 235.87
R618 B.n262 B.t13 235.87
R619 B.n118 B.t10 235.87
R620 B.n125 B.t6 235.87
R621 B.n375 B.n245 163.367
R622 B.n383 B.n245 163.367
R623 B.n383 B.n243 163.367
R624 B.n387 B.n243 163.367
R625 B.n387 B.n237 163.367
R626 B.n395 B.n237 163.367
R627 B.n395 B.n235 163.367
R628 B.n399 B.n235 163.367
R629 B.n399 B.n229 163.367
R630 B.n407 B.n229 163.367
R631 B.n407 B.n227 163.367
R632 B.n411 B.n227 163.367
R633 B.n411 B.n221 163.367
R634 B.n419 B.n221 163.367
R635 B.n419 B.n219 163.367
R636 B.n423 B.n219 163.367
R637 B.n423 B.n213 163.367
R638 B.n431 B.n213 163.367
R639 B.n431 B.n211 163.367
R640 B.n435 B.n211 163.367
R641 B.n435 B.n205 163.367
R642 B.n443 B.n205 163.367
R643 B.n443 B.n203 163.367
R644 B.n447 B.n203 163.367
R645 B.n447 B.n197 163.367
R646 B.n455 B.n197 163.367
R647 B.n455 B.n195 163.367
R648 B.n459 B.n195 163.367
R649 B.n459 B.n189 163.367
R650 B.n467 B.n189 163.367
R651 B.n467 B.n187 163.367
R652 B.n471 B.n187 163.367
R653 B.n471 B.n181 163.367
R654 B.n479 B.n181 163.367
R655 B.n479 B.n179 163.367
R656 B.n483 B.n179 163.367
R657 B.n483 B.n173 163.367
R658 B.n491 B.n173 163.367
R659 B.n491 B.n171 163.367
R660 B.n495 B.n171 163.367
R661 B.n495 B.n165 163.367
R662 B.n503 B.n165 163.367
R663 B.n503 B.n163 163.367
R664 B.n507 B.n163 163.367
R665 B.n507 B.n157 163.367
R666 B.n515 B.n157 163.367
R667 B.n515 B.n155 163.367
R668 B.n519 B.n155 163.367
R669 B.n519 B.n149 163.367
R670 B.n527 B.n149 163.367
R671 B.n527 B.n147 163.367
R672 B.n531 B.n147 163.367
R673 B.n531 B.n141 163.367
R674 B.n540 B.n141 163.367
R675 B.n540 B.n139 163.367
R676 B.n544 B.n139 163.367
R677 B.n544 B.n2 163.367
R678 B.n836 B.n2 163.367
R679 B.n836 B.n3 163.367
R680 B.n832 B.n3 163.367
R681 B.n832 B.n9 163.367
R682 B.n828 B.n9 163.367
R683 B.n828 B.n11 163.367
R684 B.n824 B.n11 163.367
R685 B.n824 B.n16 163.367
R686 B.n820 B.n16 163.367
R687 B.n820 B.n18 163.367
R688 B.n816 B.n18 163.367
R689 B.n816 B.n23 163.367
R690 B.n812 B.n23 163.367
R691 B.n812 B.n25 163.367
R692 B.n808 B.n25 163.367
R693 B.n808 B.n30 163.367
R694 B.n804 B.n30 163.367
R695 B.n804 B.n32 163.367
R696 B.n800 B.n32 163.367
R697 B.n800 B.n37 163.367
R698 B.n796 B.n37 163.367
R699 B.n796 B.n39 163.367
R700 B.n792 B.n39 163.367
R701 B.n792 B.n44 163.367
R702 B.n788 B.n44 163.367
R703 B.n788 B.n46 163.367
R704 B.n784 B.n46 163.367
R705 B.n784 B.n51 163.367
R706 B.n780 B.n51 163.367
R707 B.n780 B.n53 163.367
R708 B.n776 B.n53 163.367
R709 B.n776 B.n58 163.367
R710 B.n772 B.n58 163.367
R711 B.n772 B.n60 163.367
R712 B.n768 B.n60 163.367
R713 B.n768 B.n65 163.367
R714 B.n764 B.n65 163.367
R715 B.n764 B.n67 163.367
R716 B.n760 B.n67 163.367
R717 B.n760 B.n72 163.367
R718 B.n756 B.n72 163.367
R719 B.n756 B.n74 163.367
R720 B.n752 B.n74 163.367
R721 B.n752 B.n79 163.367
R722 B.n748 B.n79 163.367
R723 B.n748 B.n81 163.367
R724 B.n744 B.n81 163.367
R725 B.n744 B.n86 163.367
R726 B.n740 B.n86 163.367
R727 B.n740 B.n88 163.367
R728 B.n736 B.n88 163.367
R729 B.n736 B.n93 163.367
R730 B.n732 B.n93 163.367
R731 B.n732 B.n95 163.367
R732 B.n728 B.n95 163.367
R733 B.n728 B.n100 163.367
R734 B.n724 B.n100 163.367
R735 B.n724 B.n102 163.367
R736 B.n720 B.n102 163.367
R737 B.n371 B.n369 163.367
R738 B.n369 B.n368 163.367
R739 B.n365 B.n364 163.367
R740 B.n362 B.n255 163.367
R741 B.n358 B.n356 163.367
R742 B.n354 B.n257 163.367
R743 B.n350 B.n348 163.367
R744 B.n346 B.n259 163.367
R745 B.n342 B.n340 163.367
R746 B.n338 B.n261 163.367
R747 B.n333 B.n331 163.367
R748 B.n329 B.n265 163.367
R749 B.n325 B.n323 163.367
R750 B.n321 B.n267 163.367
R751 B.n317 B.n315 163.367
R752 B.n312 B.n311 163.367
R753 B.n309 B.n273 163.367
R754 B.n305 B.n303 163.367
R755 B.n301 B.n275 163.367
R756 B.n297 B.n295 163.367
R757 B.n293 B.n277 163.367
R758 B.n289 B.n287 163.367
R759 B.n285 B.n279 163.367
R760 B.n281 B.n249 163.367
R761 B.n377 B.n247 163.367
R762 B.n381 B.n247 163.367
R763 B.n381 B.n241 163.367
R764 B.n389 B.n241 163.367
R765 B.n389 B.n239 163.367
R766 B.n393 B.n239 163.367
R767 B.n393 B.n232 163.367
R768 B.n401 B.n232 163.367
R769 B.n401 B.n230 163.367
R770 B.n405 B.n230 163.367
R771 B.n405 B.n225 163.367
R772 B.n413 B.n225 163.367
R773 B.n413 B.n223 163.367
R774 B.n417 B.n223 163.367
R775 B.n417 B.n217 163.367
R776 B.n425 B.n217 163.367
R777 B.n425 B.n215 163.367
R778 B.n429 B.n215 163.367
R779 B.n429 B.n209 163.367
R780 B.n437 B.n209 163.367
R781 B.n437 B.n207 163.367
R782 B.n441 B.n207 163.367
R783 B.n441 B.n200 163.367
R784 B.n449 B.n200 163.367
R785 B.n449 B.n198 163.367
R786 B.n453 B.n198 163.367
R787 B.n453 B.n193 163.367
R788 B.n461 B.n193 163.367
R789 B.n461 B.n191 163.367
R790 B.n465 B.n191 163.367
R791 B.n465 B.n185 163.367
R792 B.n473 B.n185 163.367
R793 B.n473 B.n183 163.367
R794 B.n477 B.n183 163.367
R795 B.n477 B.n176 163.367
R796 B.n485 B.n176 163.367
R797 B.n485 B.n174 163.367
R798 B.n489 B.n174 163.367
R799 B.n489 B.n169 163.367
R800 B.n497 B.n169 163.367
R801 B.n497 B.n167 163.367
R802 B.n501 B.n167 163.367
R803 B.n501 B.n161 163.367
R804 B.n509 B.n161 163.367
R805 B.n509 B.n159 163.367
R806 B.n513 B.n159 163.367
R807 B.n513 B.n153 163.367
R808 B.n521 B.n153 163.367
R809 B.n521 B.n151 163.367
R810 B.n525 B.n151 163.367
R811 B.n525 B.n145 163.367
R812 B.n533 B.n145 163.367
R813 B.n533 B.n143 163.367
R814 B.n538 B.n143 163.367
R815 B.n538 B.n137 163.367
R816 B.n546 B.n137 163.367
R817 B.n547 B.n546 163.367
R818 B.n547 B.n5 163.367
R819 B.n6 B.n5 163.367
R820 B.n7 B.n6 163.367
R821 B.n552 B.n7 163.367
R822 B.n552 B.n12 163.367
R823 B.n13 B.n12 163.367
R824 B.n14 B.n13 163.367
R825 B.n557 B.n14 163.367
R826 B.n557 B.n19 163.367
R827 B.n20 B.n19 163.367
R828 B.n21 B.n20 163.367
R829 B.n562 B.n21 163.367
R830 B.n562 B.n26 163.367
R831 B.n27 B.n26 163.367
R832 B.n28 B.n27 163.367
R833 B.n567 B.n28 163.367
R834 B.n567 B.n33 163.367
R835 B.n34 B.n33 163.367
R836 B.n35 B.n34 163.367
R837 B.n572 B.n35 163.367
R838 B.n572 B.n40 163.367
R839 B.n41 B.n40 163.367
R840 B.n42 B.n41 163.367
R841 B.n577 B.n42 163.367
R842 B.n577 B.n47 163.367
R843 B.n48 B.n47 163.367
R844 B.n49 B.n48 163.367
R845 B.n582 B.n49 163.367
R846 B.n582 B.n54 163.367
R847 B.n55 B.n54 163.367
R848 B.n56 B.n55 163.367
R849 B.n587 B.n56 163.367
R850 B.n587 B.n61 163.367
R851 B.n62 B.n61 163.367
R852 B.n63 B.n62 163.367
R853 B.n592 B.n63 163.367
R854 B.n592 B.n68 163.367
R855 B.n69 B.n68 163.367
R856 B.n70 B.n69 163.367
R857 B.n597 B.n70 163.367
R858 B.n597 B.n75 163.367
R859 B.n76 B.n75 163.367
R860 B.n77 B.n76 163.367
R861 B.n602 B.n77 163.367
R862 B.n602 B.n82 163.367
R863 B.n83 B.n82 163.367
R864 B.n84 B.n83 163.367
R865 B.n607 B.n84 163.367
R866 B.n607 B.n89 163.367
R867 B.n90 B.n89 163.367
R868 B.n91 B.n90 163.367
R869 B.n612 B.n91 163.367
R870 B.n612 B.n96 163.367
R871 B.n97 B.n96 163.367
R872 B.n98 B.n97 163.367
R873 B.n617 B.n98 163.367
R874 B.n617 B.n103 163.367
R875 B.n104 B.n103 163.367
R876 B.n105 B.n104 163.367
R877 B.n716 B.n714 163.367
R878 B.n712 B.n109 163.367
R879 B.n708 B.n706 163.367
R880 B.n704 B.n111 163.367
R881 B.n700 B.n698 163.367
R882 B.n696 B.n113 163.367
R883 B.n692 B.n690 163.367
R884 B.n688 B.n115 163.367
R885 B.n684 B.n682 163.367
R886 B.n680 B.n117 163.367
R887 B.n676 B.n674 163.367
R888 B.n672 B.n122 163.367
R889 B.n668 B.n666 163.367
R890 B.n664 B.n124 163.367
R891 B.n659 B.n657 163.367
R892 B.n655 B.n128 163.367
R893 B.n651 B.n649 163.367
R894 B.n647 B.n130 163.367
R895 B.n643 B.n641 163.367
R896 B.n639 B.n132 163.367
R897 B.n635 B.n633 163.367
R898 B.n631 B.n134 163.367
R899 B.n627 B.n625 163.367
R900 B.n268 B.t19 157.71
R901 B.n125 B.t8 157.71
R902 B.n262 B.t16 157.707
R903 B.n118 B.t11 157.707
R904 B.n376 B.n250 150.496
R905 B.n721 B.n106 150.496
R906 B.n269 B.n268 82.4247
R907 B.n263 B.n262 82.4247
R908 B.n119 B.n118 82.4247
R909 B.n126 B.n125 82.4247
R910 B.n376 B.n246 78.1206
R911 B.n382 B.n246 78.1206
R912 B.n382 B.n242 78.1206
R913 B.n388 B.n242 78.1206
R914 B.n388 B.n238 78.1206
R915 B.n394 B.n238 78.1206
R916 B.n394 B.n233 78.1206
R917 B.n400 B.n233 78.1206
R918 B.n400 B.n234 78.1206
R919 B.n406 B.n226 78.1206
R920 B.n412 B.n226 78.1206
R921 B.n412 B.n222 78.1206
R922 B.n418 B.n222 78.1206
R923 B.n418 B.n218 78.1206
R924 B.n424 B.n218 78.1206
R925 B.n424 B.n214 78.1206
R926 B.n430 B.n214 78.1206
R927 B.n430 B.n210 78.1206
R928 B.n436 B.n210 78.1206
R929 B.n436 B.n206 78.1206
R930 B.n442 B.n206 78.1206
R931 B.n442 B.n201 78.1206
R932 B.n448 B.n201 78.1206
R933 B.n448 B.n202 78.1206
R934 B.n454 B.n194 78.1206
R935 B.n460 B.n194 78.1206
R936 B.n460 B.n190 78.1206
R937 B.n466 B.n190 78.1206
R938 B.n466 B.n186 78.1206
R939 B.n472 B.n186 78.1206
R940 B.n472 B.n182 78.1206
R941 B.n478 B.n182 78.1206
R942 B.n478 B.n177 78.1206
R943 B.n484 B.n177 78.1206
R944 B.n484 B.n178 78.1206
R945 B.n490 B.n170 78.1206
R946 B.n496 B.n170 78.1206
R947 B.n496 B.n166 78.1206
R948 B.n502 B.n166 78.1206
R949 B.n502 B.n162 78.1206
R950 B.n508 B.n162 78.1206
R951 B.n508 B.n158 78.1206
R952 B.n514 B.n158 78.1206
R953 B.n514 B.n154 78.1206
R954 B.n520 B.n154 78.1206
R955 B.n520 B.n150 78.1206
R956 B.n526 B.n150 78.1206
R957 B.n532 B.n146 78.1206
R958 B.n532 B.n142 78.1206
R959 B.n539 B.n142 78.1206
R960 B.n539 B.n138 78.1206
R961 B.n545 B.n138 78.1206
R962 B.n545 B.n4 78.1206
R963 B.n835 B.n4 78.1206
R964 B.n835 B.n834 78.1206
R965 B.n834 B.n833 78.1206
R966 B.n833 B.n8 78.1206
R967 B.n827 B.n8 78.1206
R968 B.n827 B.n826 78.1206
R969 B.n826 B.n825 78.1206
R970 B.n825 B.n15 78.1206
R971 B.n819 B.n818 78.1206
R972 B.n818 B.n817 78.1206
R973 B.n817 B.n22 78.1206
R974 B.n811 B.n22 78.1206
R975 B.n811 B.n810 78.1206
R976 B.n810 B.n809 78.1206
R977 B.n809 B.n29 78.1206
R978 B.n803 B.n29 78.1206
R979 B.n803 B.n802 78.1206
R980 B.n802 B.n801 78.1206
R981 B.n801 B.n36 78.1206
R982 B.n795 B.n36 78.1206
R983 B.n794 B.n793 78.1206
R984 B.n793 B.n43 78.1206
R985 B.n787 B.n43 78.1206
R986 B.n787 B.n786 78.1206
R987 B.n786 B.n785 78.1206
R988 B.n785 B.n50 78.1206
R989 B.n779 B.n50 78.1206
R990 B.n779 B.n778 78.1206
R991 B.n778 B.n777 78.1206
R992 B.n777 B.n57 78.1206
R993 B.n771 B.n57 78.1206
R994 B.n770 B.n769 78.1206
R995 B.n769 B.n64 78.1206
R996 B.n763 B.n64 78.1206
R997 B.n763 B.n762 78.1206
R998 B.n762 B.n761 78.1206
R999 B.n761 B.n71 78.1206
R1000 B.n755 B.n71 78.1206
R1001 B.n755 B.n754 78.1206
R1002 B.n754 B.n753 78.1206
R1003 B.n753 B.n78 78.1206
R1004 B.n747 B.n78 78.1206
R1005 B.n747 B.n746 78.1206
R1006 B.n746 B.n745 78.1206
R1007 B.n745 B.n85 78.1206
R1008 B.n739 B.n85 78.1206
R1009 B.n738 B.n737 78.1206
R1010 B.n737 B.n92 78.1206
R1011 B.n731 B.n92 78.1206
R1012 B.n731 B.n730 78.1206
R1013 B.n730 B.n729 78.1206
R1014 B.n729 B.n99 78.1206
R1015 B.n723 B.n99 78.1206
R1016 B.n723 B.n722 78.1206
R1017 B.n722 B.n721 78.1206
R1018 B.n269 B.t18 75.2858
R1019 B.n126 B.t9 75.2858
R1020 B.n263 B.t15 75.282
R1021 B.n119 B.t12 75.282
R1022 B.n370 B.n251 71.676
R1023 B.n368 B.n253 71.676
R1024 B.n364 B.n363 71.676
R1025 B.n357 B.n255 71.676
R1026 B.n356 B.n355 71.676
R1027 B.n349 B.n257 71.676
R1028 B.n348 B.n347 71.676
R1029 B.n341 B.n259 71.676
R1030 B.n340 B.n339 71.676
R1031 B.n332 B.n261 71.676
R1032 B.n331 B.n330 71.676
R1033 B.n324 B.n265 71.676
R1034 B.n323 B.n322 71.676
R1035 B.n316 B.n267 71.676
R1036 B.n315 B.n271 71.676
R1037 B.n311 B.n310 71.676
R1038 B.n304 B.n273 71.676
R1039 B.n303 B.n302 71.676
R1040 B.n296 B.n275 71.676
R1041 B.n295 B.n294 71.676
R1042 B.n288 B.n277 71.676
R1043 B.n287 B.n286 71.676
R1044 B.n280 B.n279 71.676
R1045 B.n715 B.n107 71.676
R1046 B.n714 B.n713 71.676
R1047 B.n707 B.n109 71.676
R1048 B.n706 B.n705 71.676
R1049 B.n699 B.n111 71.676
R1050 B.n698 B.n697 71.676
R1051 B.n691 B.n113 71.676
R1052 B.n690 B.n689 71.676
R1053 B.n683 B.n115 71.676
R1054 B.n682 B.n681 71.676
R1055 B.n675 B.n117 71.676
R1056 B.n674 B.n673 71.676
R1057 B.n667 B.n122 71.676
R1058 B.n666 B.n665 71.676
R1059 B.n658 B.n124 71.676
R1060 B.n657 B.n656 71.676
R1061 B.n650 B.n128 71.676
R1062 B.n649 B.n648 71.676
R1063 B.n642 B.n130 71.676
R1064 B.n641 B.n640 71.676
R1065 B.n634 B.n132 71.676
R1066 B.n633 B.n632 71.676
R1067 B.n626 B.n134 71.676
R1068 B.n625 B.n624 71.676
R1069 B.n624 B.n623 71.676
R1070 B.n627 B.n626 71.676
R1071 B.n632 B.n631 71.676
R1072 B.n635 B.n634 71.676
R1073 B.n640 B.n639 71.676
R1074 B.n643 B.n642 71.676
R1075 B.n648 B.n647 71.676
R1076 B.n651 B.n650 71.676
R1077 B.n656 B.n655 71.676
R1078 B.n659 B.n658 71.676
R1079 B.n665 B.n664 71.676
R1080 B.n668 B.n667 71.676
R1081 B.n673 B.n672 71.676
R1082 B.n676 B.n675 71.676
R1083 B.n681 B.n680 71.676
R1084 B.n684 B.n683 71.676
R1085 B.n689 B.n688 71.676
R1086 B.n692 B.n691 71.676
R1087 B.n697 B.n696 71.676
R1088 B.n700 B.n699 71.676
R1089 B.n705 B.n704 71.676
R1090 B.n708 B.n707 71.676
R1091 B.n713 B.n712 71.676
R1092 B.n716 B.n715 71.676
R1093 B.n371 B.n370 71.676
R1094 B.n365 B.n253 71.676
R1095 B.n363 B.n362 71.676
R1096 B.n358 B.n357 71.676
R1097 B.n355 B.n354 71.676
R1098 B.n350 B.n349 71.676
R1099 B.n347 B.n346 71.676
R1100 B.n342 B.n341 71.676
R1101 B.n339 B.n338 71.676
R1102 B.n333 B.n332 71.676
R1103 B.n330 B.n329 71.676
R1104 B.n325 B.n324 71.676
R1105 B.n322 B.n321 71.676
R1106 B.n317 B.n316 71.676
R1107 B.n312 B.n271 71.676
R1108 B.n310 B.n309 71.676
R1109 B.n305 B.n304 71.676
R1110 B.n302 B.n301 71.676
R1111 B.n297 B.n296 71.676
R1112 B.n294 B.n293 71.676
R1113 B.n289 B.n288 71.676
R1114 B.n286 B.n285 71.676
R1115 B.n281 B.n280 71.676
R1116 B.n454 B.t2 66.6324
R1117 B.t0 B.n146 66.6324
R1118 B.t3 B.n15 66.6324
R1119 B.n771 B.t5 66.6324
R1120 B.n270 B.n269 59.5399
R1121 B.n336 B.n263 59.5399
R1122 B.n120 B.n119 59.5399
R1123 B.n661 B.n126 59.5399
R1124 B.n178 B.t1 50.5488
R1125 B.t4 B.n794 50.5488
R1126 B.n406 B.t14 43.6558
R1127 B.n739 B.t7 43.6558
R1128 B.n234 B.t14 34.4653
R1129 B.t7 B.n738 34.4653
R1130 B.n719 B.n718 31.0639
R1131 B.n622 B.n621 31.0639
R1132 B.n378 B.n248 31.0639
R1133 B.n374 B.n373 31.0639
R1134 B.n490 B.t1 27.5723
R1135 B.n795 B.t4 27.5723
R1136 B B.n837 18.0485
R1137 B.n202 B.t2 11.4888
R1138 B.n526 B.t0 11.4888
R1139 B.n819 B.t3 11.4888
R1140 B.t5 B.n770 11.4888
R1141 B.n718 B.n717 10.6151
R1142 B.n717 B.n108 10.6151
R1143 B.n711 B.n108 10.6151
R1144 B.n711 B.n710 10.6151
R1145 B.n710 B.n709 10.6151
R1146 B.n709 B.n110 10.6151
R1147 B.n703 B.n110 10.6151
R1148 B.n703 B.n702 10.6151
R1149 B.n702 B.n701 10.6151
R1150 B.n701 B.n112 10.6151
R1151 B.n695 B.n112 10.6151
R1152 B.n695 B.n694 10.6151
R1153 B.n694 B.n693 10.6151
R1154 B.n693 B.n114 10.6151
R1155 B.n687 B.n114 10.6151
R1156 B.n687 B.n686 10.6151
R1157 B.n686 B.n685 10.6151
R1158 B.n685 B.n116 10.6151
R1159 B.n679 B.n678 10.6151
R1160 B.n678 B.n677 10.6151
R1161 B.n677 B.n121 10.6151
R1162 B.n671 B.n121 10.6151
R1163 B.n671 B.n670 10.6151
R1164 B.n670 B.n669 10.6151
R1165 B.n669 B.n123 10.6151
R1166 B.n663 B.n123 10.6151
R1167 B.n663 B.n662 10.6151
R1168 B.n660 B.n127 10.6151
R1169 B.n654 B.n127 10.6151
R1170 B.n654 B.n653 10.6151
R1171 B.n653 B.n652 10.6151
R1172 B.n652 B.n129 10.6151
R1173 B.n646 B.n129 10.6151
R1174 B.n646 B.n645 10.6151
R1175 B.n645 B.n644 10.6151
R1176 B.n644 B.n131 10.6151
R1177 B.n638 B.n131 10.6151
R1178 B.n638 B.n637 10.6151
R1179 B.n637 B.n636 10.6151
R1180 B.n636 B.n133 10.6151
R1181 B.n630 B.n133 10.6151
R1182 B.n630 B.n629 10.6151
R1183 B.n629 B.n628 10.6151
R1184 B.n628 B.n135 10.6151
R1185 B.n622 B.n135 10.6151
R1186 B.n379 B.n378 10.6151
R1187 B.n380 B.n379 10.6151
R1188 B.n380 B.n240 10.6151
R1189 B.n390 B.n240 10.6151
R1190 B.n391 B.n390 10.6151
R1191 B.n392 B.n391 10.6151
R1192 B.n392 B.n231 10.6151
R1193 B.n402 B.n231 10.6151
R1194 B.n403 B.n402 10.6151
R1195 B.n404 B.n403 10.6151
R1196 B.n404 B.n224 10.6151
R1197 B.n414 B.n224 10.6151
R1198 B.n415 B.n414 10.6151
R1199 B.n416 B.n415 10.6151
R1200 B.n416 B.n216 10.6151
R1201 B.n426 B.n216 10.6151
R1202 B.n427 B.n426 10.6151
R1203 B.n428 B.n427 10.6151
R1204 B.n428 B.n208 10.6151
R1205 B.n438 B.n208 10.6151
R1206 B.n439 B.n438 10.6151
R1207 B.n440 B.n439 10.6151
R1208 B.n440 B.n199 10.6151
R1209 B.n450 B.n199 10.6151
R1210 B.n451 B.n450 10.6151
R1211 B.n452 B.n451 10.6151
R1212 B.n452 B.n192 10.6151
R1213 B.n462 B.n192 10.6151
R1214 B.n463 B.n462 10.6151
R1215 B.n464 B.n463 10.6151
R1216 B.n464 B.n184 10.6151
R1217 B.n474 B.n184 10.6151
R1218 B.n475 B.n474 10.6151
R1219 B.n476 B.n475 10.6151
R1220 B.n476 B.n175 10.6151
R1221 B.n486 B.n175 10.6151
R1222 B.n487 B.n486 10.6151
R1223 B.n488 B.n487 10.6151
R1224 B.n488 B.n168 10.6151
R1225 B.n498 B.n168 10.6151
R1226 B.n499 B.n498 10.6151
R1227 B.n500 B.n499 10.6151
R1228 B.n500 B.n160 10.6151
R1229 B.n510 B.n160 10.6151
R1230 B.n511 B.n510 10.6151
R1231 B.n512 B.n511 10.6151
R1232 B.n512 B.n152 10.6151
R1233 B.n522 B.n152 10.6151
R1234 B.n523 B.n522 10.6151
R1235 B.n524 B.n523 10.6151
R1236 B.n524 B.n144 10.6151
R1237 B.n534 B.n144 10.6151
R1238 B.n535 B.n534 10.6151
R1239 B.n537 B.n535 10.6151
R1240 B.n537 B.n536 10.6151
R1241 B.n536 B.n136 10.6151
R1242 B.n548 B.n136 10.6151
R1243 B.n549 B.n548 10.6151
R1244 B.n550 B.n549 10.6151
R1245 B.n551 B.n550 10.6151
R1246 B.n553 B.n551 10.6151
R1247 B.n554 B.n553 10.6151
R1248 B.n555 B.n554 10.6151
R1249 B.n556 B.n555 10.6151
R1250 B.n558 B.n556 10.6151
R1251 B.n559 B.n558 10.6151
R1252 B.n560 B.n559 10.6151
R1253 B.n561 B.n560 10.6151
R1254 B.n563 B.n561 10.6151
R1255 B.n564 B.n563 10.6151
R1256 B.n565 B.n564 10.6151
R1257 B.n566 B.n565 10.6151
R1258 B.n568 B.n566 10.6151
R1259 B.n569 B.n568 10.6151
R1260 B.n570 B.n569 10.6151
R1261 B.n571 B.n570 10.6151
R1262 B.n573 B.n571 10.6151
R1263 B.n574 B.n573 10.6151
R1264 B.n575 B.n574 10.6151
R1265 B.n576 B.n575 10.6151
R1266 B.n578 B.n576 10.6151
R1267 B.n579 B.n578 10.6151
R1268 B.n580 B.n579 10.6151
R1269 B.n581 B.n580 10.6151
R1270 B.n583 B.n581 10.6151
R1271 B.n584 B.n583 10.6151
R1272 B.n585 B.n584 10.6151
R1273 B.n586 B.n585 10.6151
R1274 B.n588 B.n586 10.6151
R1275 B.n589 B.n588 10.6151
R1276 B.n590 B.n589 10.6151
R1277 B.n591 B.n590 10.6151
R1278 B.n593 B.n591 10.6151
R1279 B.n594 B.n593 10.6151
R1280 B.n595 B.n594 10.6151
R1281 B.n596 B.n595 10.6151
R1282 B.n598 B.n596 10.6151
R1283 B.n599 B.n598 10.6151
R1284 B.n600 B.n599 10.6151
R1285 B.n601 B.n600 10.6151
R1286 B.n603 B.n601 10.6151
R1287 B.n604 B.n603 10.6151
R1288 B.n605 B.n604 10.6151
R1289 B.n606 B.n605 10.6151
R1290 B.n608 B.n606 10.6151
R1291 B.n609 B.n608 10.6151
R1292 B.n610 B.n609 10.6151
R1293 B.n611 B.n610 10.6151
R1294 B.n613 B.n611 10.6151
R1295 B.n614 B.n613 10.6151
R1296 B.n615 B.n614 10.6151
R1297 B.n616 B.n615 10.6151
R1298 B.n618 B.n616 10.6151
R1299 B.n619 B.n618 10.6151
R1300 B.n620 B.n619 10.6151
R1301 B.n621 B.n620 10.6151
R1302 B.n373 B.n372 10.6151
R1303 B.n372 B.n252 10.6151
R1304 B.n367 B.n252 10.6151
R1305 B.n367 B.n366 10.6151
R1306 B.n366 B.n254 10.6151
R1307 B.n361 B.n254 10.6151
R1308 B.n361 B.n360 10.6151
R1309 B.n360 B.n359 10.6151
R1310 B.n359 B.n256 10.6151
R1311 B.n353 B.n256 10.6151
R1312 B.n353 B.n352 10.6151
R1313 B.n352 B.n351 10.6151
R1314 B.n351 B.n258 10.6151
R1315 B.n345 B.n258 10.6151
R1316 B.n345 B.n344 10.6151
R1317 B.n344 B.n343 10.6151
R1318 B.n343 B.n260 10.6151
R1319 B.n337 B.n260 10.6151
R1320 B.n335 B.n334 10.6151
R1321 B.n334 B.n264 10.6151
R1322 B.n328 B.n264 10.6151
R1323 B.n328 B.n327 10.6151
R1324 B.n327 B.n326 10.6151
R1325 B.n326 B.n266 10.6151
R1326 B.n320 B.n266 10.6151
R1327 B.n320 B.n319 10.6151
R1328 B.n319 B.n318 10.6151
R1329 B.n314 B.n313 10.6151
R1330 B.n313 B.n272 10.6151
R1331 B.n308 B.n272 10.6151
R1332 B.n308 B.n307 10.6151
R1333 B.n307 B.n306 10.6151
R1334 B.n306 B.n274 10.6151
R1335 B.n300 B.n274 10.6151
R1336 B.n300 B.n299 10.6151
R1337 B.n299 B.n298 10.6151
R1338 B.n298 B.n276 10.6151
R1339 B.n292 B.n276 10.6151
R1340 B.n292 B.n291 10.6151
R1341 B.n291 B.n290 10.6151
R1342 B.n290 B.n278 10.6151
R1343 B.n284 B.n278 10.6151
R1344 B.n284 B.n283 10.6151
R1345 B.n283 B.n282 10.6151
R1346 B.n282 B.n248 10.6151
R1347 B.n374 B.n244 10.6151
R1348 B.n384 B.n244 10.6151
R1349 B.n385 B.n384 10.6151
R1350 B.n386 B.n385 10.6151
R1351 B.n386 B.n236 10.6151
R1352 B.n396 B.n236 10.6151
R1353 B.n397 B.n396 10.6151
R1354 B.n398 B.n397 10.6151
R1355 B.n398 B.n228 10.6151
R1356 B.n408 B.n228 10.6151
R1357 B.n409 B.n408 10.6151
R1358 B.n410 B.n409 10.6151
R1359 B.n410 B.n220 10.6151
R1360 B.n420 B.n220 10.6151
R1361 B.n421 B.n420 10.6151
R1362 B.n422 B.n421 10.6151
R1363 B.n422 B.n212 10.6151
R1364 B.n432 B.n212 10.6151
R1365 B.n433 B.n432 10.6151
R1366 B.n434 B.n433 10.6151
R1367 B.n434 B.n204 10.6151
R1368 B.n444 B.n204 10.6151
R1369 B.n445 B.n444 10.6151
R1370 B.n446 B.n445 10.6151
R1371 B.n446 B.n196 10.6151
R1372 B.n456 B.n196 10.6151
R1373 B.n457 B.n456 10.6151
R1374 B.n458 B.n457 10.6151
R1375 B.n458 B.n188 10.6151
R1376 B.n468 B.n188 10.6151
R1377 B.n469 B.n468 10.6151
R1378 B.n470 B.n469 10.6151
R1379 B.n470 B.n180 10.6151
R1380 B.n480 B.n180 10.6151
R1381 B.n481 B.n480 10.6151
R1382 B.n482 B.n481 10.6151
R1383 B.n482 B.n172 10.6151
R1384 B.n492 B.n172 10.6151
R1385 B.n493 B.n492 10.6151
R1386 B.n494 B.n493 10.6151
R1387 B.n494 B.n164 10.6151
R1388 B.n504 B.n164 10.6151
R1389 B.n505 B.n504 10.6151
R1390 B.n506 B.n505 10.6151
R1391 B.n506 B.n156 10.6151
R1392 B.n516 B.n156 10.6151
R1393 B.n517 B.n516 10.6151
R1394 B.n518 B.n517 10.6151
R1395 B.n518 B.n148 10.6151
R1396 B.n528 B.n148 10.6151
R1397 B.n529 B.n528 10.6151
R1398 B.n530 B.n529 10.6151
R1399 B.n530 B.n140 10.6151
R1400 B.n541 B.n140 10.6151
R1401 B.n542 B.n541 10.6151
R1402 B.n543 B.n542 10.6151
R1403 B.n543 B.n0 10.6151
R1404 B.n831 B.n1 10.6151
R1405 B.n831 B.n830 10.6151
R1406 B.n830 B.n829 10.6151
R1407 B.n829 B.n10 10.6151
R1408 B.n823 B.n10 10.6151
R1409 B.n823 B.n822 10.6151
R1410 B.n822 B.n821 10.6151
R1411 B.n821 B.n17 10.6151
R1412 B.n815 B.n17 10.6151
R1413 B.n815 B.n814 10.6151
R1414 B.n814 B.n813 10.6151
R1415 B.n813 B.n24 10.6151
R1416 B.n807 B.n24 10.6151
R1417 B.n807 B.n806 10.6151
R1418 B.n806 B.n805 10.6151
R1419 B.n805 B.n31 10.6151
R1420 B.n799 B.n31 10.6151
R1421 B.n799 B.n798 10.6151
R1422 B.n798 B.n797 10.6151
R1423 B.n797 B.n38 10.6151
R1424 B.n791 B.n38 10.6151
R1425 B.n791 B.n790 10.6151
R1426 B.n790 B.n789 10.6151
R1427 B.n789 B.n45 10.6151
R1428 B.n783 B.n45 10.6151
R1429 B.n783 B.n782 10.6151
R1430 B.n782 B.n781 10.6151
R1431 B.n781 B.n52 10.6151
R1432 B.n775 B.n52 10.6151
R1433 B.n775 B.n774 10.6151
R1434 B.n774 B.n773 10.6151
R1435 B.n773 B.n59 10.6151
R1436 B.n767 B.n59 10.6151
R1437 B.n767 B.n766 10.6151
R1438 B.n766 B.n765 10.6151
R1439 B.n765 B.n66 10.6151
R1440 B.n759 B.n66 10.6151
R1441 B.n759 B.n758 10.6151
R1442 B.n758 B.n757 10.6151
R1443 B.n757 B.n73 10.6151
R1444 B.n751 B.n73 10.6151
R1445 B.n751 B.n750 10.6151
R1446 B.n750 B.n749 10.6151
R1447 B.n749 B.n80 10.6151
R1448 B.n743 B.n80 10.6151
R1449 B.n743 B.n742 10.6151
R1450 B.n742 B.n741 10.6151
R1451 B.n741 B.n87 10.6151
R1452 B.n735 B.n87 10.6151
R1453 B.n735 B.n734 10.6151
R1454 B.n734 B.n733 10.6151
R1455 B.n733 B.n94 10.6151
R1456 B.n727 B.n94 10.6151
R1457 B.n727 B.n726 10.6151
R1458 B.n726 B.n725 10.6151
R1459 B.n725 B.n101 10.6151
R1460 B.n719 B.n101 10.6151
R1461 B.n120 B.n116 9.36635
R1462 B.n661 B.n660 9.36635
R1463 B.n337 B.n336 9.36635
R1464 B.n314 B.n270 9.36635
R1465 B.n837 B.n0 2.81026
R1466 B.n837 B.n1 2.81026
R1467 B.n679 B.n120 1.24928
R1468 B.n662 B.n661 1.24928
R1469 B.n336 B.n335 1.24928
R1470 B.n318 B.n270 1.24928
R1471 VP.n15 VP.n14 161.3
R1472 VP.n16 VP.n11 161.3
R1473 VP.n18 VP.n17 161.3
R1474 VP.n19 VP.n10 161.3
R1475 VP.n21 VP.n20 161.3
R1476 VP.n22 VP.n9 161.3
R1477 VP.n24 VP.n23 161.3
R1478 VP.n25 VP.n8 161.3
R1479 VP.n54 VP.n0 161.3
R1480 VP.n53 VP.n52 161.3
R1481 VP.n51 VP.n1 161.3
R1482 VP.n50 VP.n49 161.3
R1483 VP.n48 VP.n2 161.3
R1484 VP.n47 VP.n46 161.3
R1485 VP.n45 VP.n3 161.3
R1486 VP.n44 VP.n43 161.3
R1487 VP.n41 VP.n4 161.3
R1488 VP.n40 VP.n39 161.3
R1489 VP.n38 VP.n5 161.3
R1490 VP.n37 VP.n36 161.3
R1491 VP.n35 VP.n6 161.3
R1492 VP.n34 VP.n33 161.3
R1493 VP.n32 VP.n7 161.3
R1494 VP.n31 VP.n30 161.3
R1495 VP.n13 VP.n12 63.0913
R1496 VP.n12 VP.t0 58.5062
R1497 VP.n29 VP.n28 57.7881
R1498 VP.n56 VP.n55 57.7881
R1499 VP.n27 VP.n26 57.7881
R1500 VP.n36 VP.n35 52.6866
R1501 VP.n49 VP.n48 52.6866
R1502 VP.n20 VP.n19 52.6866
R1503 VP.n28 VP.n27 48.3113
R1504 VP.n35 VP.n34 28.4674
R1505 VP.n49 VP.n1 28.4674
R1506 VP.n20 VP.n9 28.4674
R1507 VP.n55 VP.t2 26.4367
R1508 VP.n29 VP.t4 26.4367
R1509 VP.n42 VP.t3 26.4367
R1510 VP.n26 VP.t5 26.4367
R1511 VP.n13 VP.t1 26.4367
R1512 VP.n30 VP.n29 24.5923
R1513 VP.n30 VP.n7 24.5923
R1514 VP.n34 VP.n7 24.5923
R1515 VP.n36 VP.n5 24.5923
R1516 VP.n40 VP.n5 24.5923
R1517 VP.n41 VP.n40 24.5923
R1518 VP.n43 VP.n3 24.5923
R1519 VP.n47 VP.n3 24.5923
R1520 VP.n48 VP.n47 24.5923
R1521 VP.n53 VP.n1 24.5923
R1522 VP.n54 VP.n53 24.5923
R1523 VP.n55 VP.n54 24.5923
R1524 VP.n24 VP.n9 24.5923
R1525 VP.n25 VP.n24 24.5923
R1526 VP.n26 VP.n25 24.5923
R1527 VP.n14 VP.n11 24.5923
R1528 VP.n18 VP.n11 24.5923
R1529 VP.n19 VP.n18 24.5923
R1530 VP.n42 VP.n41 12.2964
R1531 VP.n43 VP.n42 12.2964
R1532 VP.n14 VP.n13 12.2964
R1533 VP.n15 VP.n12 2.52309
R1534 VP.n27 VP.n8 0.417304
R1535 VP.n31 VP.n28 0.417304
R1536 VP.n56 VP.n0 0.417304
R1537 VP VP.n56 0.394524
R1538 VP.n16 VP.n15 0.189894
R1539 VP.n17 VP.n16 0.189894
R1540 VP.n17 VP.n10 0.189894
R1541 VP.n21 VP.n10 0.189894
R1542 VP.n22 VP.n21 0.189894
R1543 VP.n23 VP.n22 0.189894
R1544 VP.n23 VP.n8 0.189894
R1545 VP.n32 VP.n31 0.189894
R1546 VP.n33 VP.n32 0.189894
R1547 VP.n33 VP.n6 0.189894
R1548 VP.n37 VP.n6 0.189894
R1549 VP.n38 VP.n37 0.189894
R1550 VP.n39 VP.n38 0.189894
R1551 VP.n39 VP.n4 0.189894
R1552 VP.n44 VP.n4 0.189894
R1553 VP.n45 VP.n44 0.189894
R1554 VP.n46 VP.n45 0.189894
R1555 VP.n46 VP.n2 0.189894
R1556 VP.n50 VP.n2 0.189894
R1557 VP.n51 VP.n50 0.189894
R1558 VP.n52 VP.n51 0.189894
R1559 VP.n52 VP.n0 0.189894
R1560 VTAIL.n7 VTAIL.t6 61.7837
R1561 VTAIL.n11 VTAIL.t8 61.7835
R1562 VTAIL.n2 VTAIL.t4 61.7835
R1563 VTAIL.n10 VTAIL.t2 61.7835
R1564 VTAIL.n9 VTAIL.n8 57.179
R1565 VTAIL.n6 VTAIL.n5 57.179
R1566 VTAIL.n1 VTAIL.n0 57.1788
R1567 VTAIL.n4 VTAIL.n3 57.1788
R1568 VTAIL.n6 VTAIL.n4 23.4014
R1569 VTAIL.n11 VTAIL.n10 19.7376
R1570 VTAIL.n0 VTAIL.t10 4.60515
R1571 VTAIL.n0 VTAIL.t9 4.60515
R1572 VTAIL.n3 VTAIL.t1 4.60515
R1573 VTAIL.n3 VTAIL.t5 4.60515
R1574 VTAIL.n8 VTAIL.t0 4.60515
R1575 VTAIL.n8 VTAIL.t3 4.60515
R1576 VTAIL.n5 VTAIL.t7 4.60515
R1577 VTAIL.n5 VTAIL.t11 4.60515
R1578 VTAIL.n7 VTAIL.n6 3.66429
R1579 VTAIL.n10 VTAIL.n9 3.66429
R1580 VTAIL.n4 VTAIL.n2 3.66429
R1581 VTAIL VTAIL.n11 2.69016
R1582 VTAIL.n9 VTAIL.n7 2.30222
R1583 VTAIL.n2 VTAIL.n1 2.30222
R1584 VTAIL VTAIL.n1 0.974638
R1585 VDD1 VDD1.t5 81.2685
R1586 VDD1.n1 VDD1.t1 81.1548
R1587 VDD1.n1 VDD1.n0 74.7182
R1588 VDD1.n3 VDD1.n2 73.8577
R1589 VDD1.n3 VDD1.n1 41.7444
R1590 VDD1.n2 VDD1.t4 4.60515
R1591 VDD1.n2 VDD1.t0 4.60515
R1592 VDD1.n0 VDD1.t2 4.60515
R1593 VDD1.n0 VDD1.t3 4.60515
R1594 VDD1 VDD1.n3 0.858259
R1595 VN.n37 VN.n20 161.3
R1596 VN.n36 VN.n35 161.3
R1597 VN.n34 VN.n21 161.3
R1598 VN.n33 VN.n32 161.3
R1599 VN.n31 VN.n22 161.3
R1600 VN.n30 VN.n29 161.3
R1601 VN.n28 VN.n23 161.3
R1602 VN.n27 VN.n26 161.3
R1603 VN.n17 VN.n0 161.3
R1604 VN.n16 VN.n15 161.3
R1605 VN.n14 VN.n1 161.3
R1606 VN.n13 VN.n12 161.3
R1607 VN.n11 VN.n2 161.3
R1608 VN.n10 VN.n9 161.3
R1609 VN.n8 VN.n3 161.3
R1610 VN.n7 VN.n6 161.3
R1611 VN.n5 VN.n4 63.0912
R1612 VN.n25 VN.n24 63.0912
R1613 VN.n4 VN.t0 58.5067
R1614 VN.n24 VN.t2 58.5067
R1615 VN.n19 VN.n18 57.7881
R1616 VN.n39 VN.n38 57.7881
R1617 VN.n12 VN.n11 52.6866
R1618 VN.n32 VN.n31 52.6866
R1619 VN VN.n39 48.3491
R1620 VN.n12 VN.n1 28.4674
R1621 VN.n32 VN.n21 28.4674
R1622 VN.n18 VN.t4 26.4367
R1623 VN.n5 VN.t1 26.4367
R1624 VN.n38 VN.t3 26.4367
R1625 VN.n25 VN.t5 26.4367
R1626 VN.n6 VN.n3 24.5923
R1627 VN.n10 VN.n3 24.5923
R1628 VN.n11 VN.n10 24.5923
R1629 VN.n16 VN.n1 24.5923
R1630 VN.n17 VN.n16 24.5923
R1631 VN.n18 VN.n17 24.5923
R1632 VN.n31 VN.n30 24.5923
R1633 VN.n30 VN.n23 24.5923
R1634 VN.n26 VN.n23 24.5923
R1635 VN.n38 VN.n37 24.5923
R1636 VN.n37 VN.n36 24.5923
R1637 VN.n36 VN.n21 24.5923
R1638 VN.n6 VN.n5 12.2964
R1639 VN.n26 VN.n25 12.2964
R1640 VN.n27 VN.n24 2.52312
R1641 VN.n7 VN.n4 2.52312
R1642 VN.n39 VN.n20 0.417304
R1643 VN.n19 VN.n0 0.417304
R1644 VN VN.n19 0.394524
R1645 VN.n35 VN.n20 0.189894
R1646 VN.n35 VN.n34 0.189894
R1647 VN.n34 VN.n33 0.189894
R1648 VN.n33 VN.n22 0.189894
R1649 VN.n29 VN.n22 0.189894
R1650 VN.n29 VN.n28 0.189894
R1651 VN.n28 VN.n27 0.189894
R1652 VN.n8 VN.n7 0.189894
R1653 VN.n9 VN.n8 0.189894
R1654 VN.n9 VN.n2 0.189894
R1655 VN.n13 VN.n2 0.189894
R1656 VN.n14 VN.n13 0.189894
R1657 VN.n15 VN.n14 0.189894
R1658 VN.n15 VN.n0 0.189894
R1659 VDD2.n1 VDD2.t5 81.1548
R1660 VDD2.n2 VDD2.t2 78.4625
R1661 VDD2.n1 VDD2.n0 74.7182
R1662 VDD2 VDD2.n3 74.7155
R1663 VDD2.n2 VDD2.n1 39.3295
R1664 VDD2.n3 VDD2.t0 4.60515
R1665 VDD2.n3 VDD2.t3 4.60515
R1666 VDD2.n0 VDD2.t4 4.60515
R1667 VDD2.n0 VDD2.t1 4.60515
R1668 VDD2 VDD2.n2 2.80653
C0 VN VDD2 2.83551f
C1 VDD1 VDD2 1.92173f
C2 VTAIL VP 3.93777f
C3 VTAIL VN 3.92339f
C4 VN VP 6.78355f
C5 VDD1 VTAIL 5.79579f
C6 VDD1 VP 3.25055f
C7 VDD1 VN 0.157013f
C8 VTAIL VDD2 5.85766f
C9 VP VDD2 0.574655f
C10 VDD2 B 5.635012f
C11 VDD1 B 6.021833f
C12 VTAIL B 5.039178f
C13 VN B 16.103039f
C14 VP B 14.739175f
C15 VDD2.t5 B 0.776714f
C16 VDD2.t4 B 0.07542f
C17 VDD2.t1 B 0.07542f
C18 VDD2.n0 B 0.605832f
C19 VDD2.n1 B 2.63979f
C20 VDD2.t2 B 0.762826f
C21 VDD2.n2 B 2.24471f
C22 VDD2.t0 B 0.07542f
C23 VDD2.t3 B 0.07542f
C24 VDD2.n3 B 0.605803f
C25 VN.n0 B 0.042704f
C26 VN.t4 B 0.989603f
C27 VN.n1 B 0.04449f
C28 VN.n2 B 0.02271f
C29 VN.n3 B 0.042113f
C30 VN.t0 B 1.29688f
C31 VN.n4 B 0.467198f
C32 VN.t1 B 0.989603f
C33 VN.n5 B 0.460341f
C34 VN.n6 B 0.031718f
C35 VN.n7 B 0.296479f
C36 VN.n8 B 0.02271f
C37 VN.n9 B 0.02271f
C38 VN.n10 B 0.042113f
C39 VN.n11 B 0.040339f
C40 VN.n12 B 0.023307f
C41 VN.n13 B 0.02271f
C42 VN.n14 B 0.02271f
C43 VN.n15 B 0.02271f
C44 VN.n16 B 0.042113f
C45 VN.n17 B 0.042113f
C46 VN.n18 B 0.48345f
C47 VN.n19 B 0.066094f
C48 VN.n20 B 0.042704f
C49 VN.t3 B 0.989603f
C50 VN.n21 B 0.04449f
C51 VN.n22 B 0.02271f
C52 VN.n23 B 0.042113f
C53 VN.t2 B 1.29688f
C54 VN.n24 B 0.467198f
C55 VN.t5 B 0.989603f
C56 VN.n25 B 0.460341f
C57 VN.n26 B 0.031718f
C58 VN.n27 B 0.296479f
C59 VN.n28 B 0.02271f
C60 VN.n29 B 0.02271f
C61 VN.n30 B 0.042113f
C62 VN.n31 B 0.040339f
C63 VN.n32 B 0.023307f
C64 VN.n33 B 0.02271f
C65 VN.n34 B 0.02271f
C66 VN.n35 B 0.02271f
C67 VN.n36 B 0.042113f
C68 VN.n37 B 0.042113f
C69 VN.n38 B 0.48345f
C70 VN.n39 B 1.26083f
C71 VDD1.t5 B 0.805713f
C72 VDD1.t1 B 0.804842f
C73 VDD1.t2 B 0.078151f
C74 VDD1.t3 B 0.078151f
C75 VDD1.n0 B 0.627771f
C76 VDD1.n1 B 2.87371f
C77 VDD1.t4 B 0.078151f
C78 VDD1.t0 B 0.078151f
C79 VDD1.n2 B 0.621716f
C80 VDD1.n3 B 2.35534f
C81 VTAIL.t10 B 0.105267f
C82 VTAIL.t9 B 0.105267f
C83 VTAIL.n0 B 0.768265f
C84 VTAIL.n1 B 0.597095f
C85 VTAIL.t4 B 0.984548f
C86 VTAIL.n2 B 0.936392f
C87 VTAIL.t1 B 0.105267f
C88 VTAIL.t5 B 0.105267f
C89 VTAIL.n3 B 0.768265f
C90 VTAIL.n4 B 2.15812f
C91 VTAIL.t7 B 0.105267f
C92 VTAIL.t11 B 0.105267f
C93 VTAIL.n5 B 0.768269f
C94 VTAIL.n6 B 2.15812f
C95 VTAIL.t6 B 0.984552f
C96 VTAIL.n7 B 0.936389f
C97 VTAIL.t0 B 0.105267f
C98 VTAIL.t3 B 0.105267f
C99 VTAIL.n8 B 0.768269f
C100 VTAIL.n9 B 0.865579f
C101 VTAIL.t2 B 0.984548f
C102 VTAIL.n10 B 1.86321f
C103 VTAIL.t8 B 0.984548f
C104 VTAIL.n11 B 1.76596f
C105 VP.n0 B 0.044391f
C106 VP.t2 B 1.02869f
C107 VP.n1 B 0.046247f
C108 VP.n2 B 0.023606f
C109 VP.n3 B 0.043776f
C110 VP.n4 B 0.023606f
C111 VP.t3 B 1.02869f
C112 VP.n5 B 0.043776f
C113 VP.n6 B 0.023606f
C114 VP.n7 B 0.043776f
C115 VP.n8 B 0.044391f
C116 VP.t5 B 1.02869f
C117 VP.n9 B 0.046247f
C118 VP.n10 B 0.023606f
C119 VP.n11 B 0.043776f
C120 VP.t0 B 1.34809f
C121 VP.n12 B 0.485652f
C122 VP.t1 B 1.02869f
C123 VP.n13 B 0.478522f
C124 VP.n14 B 0.03297f
C125 VP.n15 B 0.308189f
C126 VP.n16 B 0.023606f
C127 VP.n17 B 0.023606f
C128 VP.n18 B 0.043776f
C129 VP.n19 B 0.041932f
C130 VP.n20 B 0.024228f
C131 VP.n21 B 0.023606f
C132 VP.n22 B 0.023606f
C133 VP.n23 B 0.023606f
C134 VP.n24 B 0.043776f
C135 VP.n25 B 0.043776f
C136 VP.n26 B 0.502544f
C137 VP.n27 B 1.30431f
C138 VP.n28 B 1.32192f
C139 VP.t4 B 1.02869f
C140 VP.n29 B 0.502544f
C141 VP.n30 B 0.043776f
C142 VP.n31 B 0.044391f
C143 VP.n32 B 0.023606f
C144 VP.n33 B 0.023606f
C145 VP.n34 B 0.046247f
C146 VP.n35 B 0.024228f
C147 VP.n36 B 0.041932f
C148 VP.n37 B 0.023606f
C149 VP.n38 B 0.023606f
C150 VP.n39 B 0.023606f
C151 VP.n40 B 0.043776f
C152 VP.n41 B 0.03297f
C153 VP.n42 B 0.393322f
C154 VP.n43 B 0.03297f
C155 VP.n44 B 0.023606f
C156 VP.n45 B 0.023606f
C157 VP.n46 B 0.023606f
C158 VP.n47 B 0.043776f
C159 VP.n48 B 0.041932f
C160 VP.n49 B 0.024228f
C161 VP.n50 B 0.023606f
C162 VP.n51 B 0.023606f
C163 VP.n52 B 0.023606f
C164 VP.n53 B 0.043776f
C165 VP.n54 B 0.043776f
C166 VP.n55 B 0.502544f
C167 VP.n56 B 0.068704f
.ends

