* NGSPICE file created from diff_pair_sample_0304.ext - technology: sky130A

.subckt diff_pair_sample_0304 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 B.t23 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=2.2425 ps=12.28 w=5.75 l=0.46
X1 VDD1.t9 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=2.2425 ps=12.28 w=5.75 l=0.46
X2 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0 ps=0 w=5.75 l=0.46
X3 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0 ps=0 w=5.75 l=0.46
X4 VTAIL.t15 VP.t1 VDD1.t8 B.t20 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X5 VDD1.t7 VP.t2 VTAIL.t16 B.t22 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0.94875 ps=6.08 w=5.75 l=0.46
X6 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0 ps=0 w=5.75 l=0.46
X7 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0 ps=0 w=5.75 l=0.46
X8 VDD2.t8 VN.t1 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0.94875 ps=6.08 w=5.75 l=0.46
X9 VTAIL.t17 VP.t3 VDD1.t6 B.t19 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X10 VDD2.t7 VN.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X11 VDD2.t6 VN.t3 VTAIL.t9 B.t21 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X12 VDD1.t5 VP.t4 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=2.2425 ps=12.28 w=5.75 l=0.46
X13 VTAIL.t14 VN.t4 VDD2.t5 B.t20 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X14 VTAIL.t0 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X15 VDD2.t4 VN.t5 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=2.2425 ps=12.28 w=5.75 l=0.46
X16 VTAIL.t6 VN.t6 VDD2.t3 B.t19 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X17 VDD1.t3 VP.t6 VTAIL.t19 B.t21 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X18 VDD1.t2 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X19 VTAIL.t3 VP.t8 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X20 VDD1.t0 VP.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0.94875 ps=6.08 w=5.75 l=0.46
X21 VDD2.t2 VN.t7 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.2425 pd=12.28 as=0.94875 ps=6.08 w=5.75 l=0.46
X22 VTAIL.t13 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
X23 VTAIL.t5 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.94875 pd=6.08 as=0.94875 ps=6.08 w=5.75 l=0.46
R0 VN.n2 VN.t7 408.154
R1 VN.n14 VN.t5 408.154
R2 VN.n3 VN.t8 387.173
R3 VN.n1 VN.t3 387.173
R4 VN.n9 VN.t9 387.173
R5 VN.n10 VN.t0 387.173
R6 VN.n15 VN.t6 387.173
R7 VN.n13 VN.t2 387.173
R8 VN.n21 VN.t4 387.173
R9 VN.n22 VN.t1 387.173
R10 VN.n11 VN.n10 161.3
R11 VN.n23 VN.n22 161.3
R12 VN.n21 VN.n12 161.3
R13 VN.n20 VN.n19 161.3
R14 VN.n18 VN.n13 161.3
R15 VN.n17 VN.n16 161.3
R16 VN.n9 VN.n0 161.3
R17 VN.n8 VN.n7 161.3
R18 VN.n6 VN.n1 161.3
R19 VN.n5 VN.n4 161.3
R20 VN.n17 VN.n14 70.4033
R21 VN.n5 VN.n2 70.4033
R22 VN.n10 VN.n9 48.2005
R23 VN.n22 VN.n21 48.2005
R24 VN.n4 VN.n1 39.4369
R25 VN.n8 VN.n1 39.4369
R26 VN.n16 VN.n13 39.4369
R27 VN.n20 VN.n13 39.4369
R28 VN VN.n23 37.0819
R29 VN.n15 VN.n14 20.9576
R30 VN.n3 VN.n2 20.9576
R31 VN.n4 VN.n3 8.76414
R32 VN.n9 VN.n8 8.76414
R33 VN.n16 VN.n15 8.76414
R34 VN.n21 VN.n20 8.76414
R35 VN.n23 VN.n12 0.189894
R36 VN.n19 VN.n12 0.189894
R37 VN.n19 VN.n18 0.189894
R38 VN.n18 VN.n17 0.189894
R39 VN.n6 VN.n5 0.189894
R40 VN.n7 VN.n6 0.189894
R41 VN.n7 VN.n0 0.189894
R42 VN.n11 VN.n0 0.189894
R43 VN VN.n11 0.0516364
R44 VTAIL.n11 VTAIL.t8 56.768
R45 VTAIL.n17 VTAIL.t10 56.7678
R46 VTAIL.n2 VTAIL.t1 56.7678
R47 VTAIL.n16 VTAIL.t18 56.7678
R48 VTAIL.n15 VTAIL.n14 53.3246
R49 VTAIL.n13 VTAIL.n12 53.3246
R50 VTAIL.n10 VTAIL.n9 53.3246
R51 VTAIL.n8 VTAIL.n7 53.3246
R52 VTAIL.n19 VTAIL.n18 53.3244
R53 VTAIL.n1 VTAIL.n0 53.3244
R54 VTAIL.n4 VTAIL.n3 53.3244
R55 VTAIL.n6 VTAIL.n5 53.3244
R56 VTAIL.n8 VTAIL.n6 18.6858
R57 VTAIL.n17 VTAIL.n16 18.0048
R58 VTAIL.n18 VTAIL.t9 3.44398
R59 VTAIL.n18 VTAIL.t5 3.44398
R60 VTAIL.n0 VTAIL.t12 3.44398
R61 VTAIL.n0 VTAIL.t13 3.44398
R62 VTAIL.n3 VTAIL.t2 3.44398
R63 VTAIL.n3 VTAIL.t17 3.44398
R64 VTAIL.n5 VTAIL.t16 3.44398
R65 VTAIL.n5 VTAIL.t15 3.44398
R66 VTAIL.n14 VTAIL.t19 3.44398
R67 VTAIL.n14 VTAIL.t3 3.44398
R68 VTAIL.n12 VTAIL.t4 3.44398
R69 VTAIL.n12 VTAIL.t0 3.44398
R70 VTAIL.n9 VTAIL.t7 3.44398
R71 VTAIL.n9 VTAIL.t6 3.44398
R72 VTAIL.n7 VTAIL.t11 3.44398
R73 VTAIL.n7 VTAIL.t14 3.44398
R74 VTAIL.n13 VTAIL.n11 0.810845
R75 VTAIL.n2 VTAIL.n1 0.810845
R76 VTAIL.n10 VTAIL.n8 0.681535
R77 VTAIL.n11 VTAIL.n10 0.681535
R78 VTAIL.n15 VTAIL.n13 0.681535
R79 VTAIL.n16 VTAIL.n15 0.681535
R80 VTAIL.n6 VTAIL.n4 0.681535
R81 VTAIL.n4 VTAIL.n2 0.681535
R82 VTAIL.n19 VTAIL.n17 0.681535
R83 VTAIL VTAIL.n1 0.569465
R84 VTAIL VTAIL.n19 0.112569
R85 VDD2.n1 VDD2.t2 74.1277
R86 VDD2.n4 VDD2.t8 73.4468
R87 VDD2.n3 VDD2.n2 70.4586
R88 VDD2 VDD2.n7 70.4558
R89 VDD2.n6 VDD2.n5 70.0034
R90 VDD2.n1 VDD2.n0 70.0031
R91 VDD2.n4 VDD2.n3 31.9071
R92 VDD2.n7 VDD2.t3 3.44398
R93 VDD2.n7 VDD2.t4 3.44398
R94 VDD2.n5 VDD2.t5 3.44398
R95 VDD2.n5 VDD2.t7 3.44398
R96 VDD2.n2 VDD2.t0 3.44398
R97 VDD2.n2 VDD2.t9 3.44398
R98 VDD2.n0 VDD2.t1 3.44398
R99 VDD2.n0 VDD2.t6 3.44398
R100 VDD2.n6 VDD2.n4 0.681535
R101 VDD2 VDD2.n6 0.228948
R102 VDD2.n3 VDD2.n1 0.115413
R103 B.n359 B.n358 585
R104 B.n361 B.n76 585
R105 B.n364 B.n363 585
R106 B.n365 B.n75 585
R107 B.n367 B.n366 585
R108 B.n369 B.n74 585
R109 B.n372 B.n371 585
R110 B.n373 B.n73 585
R111 B.n375 B.n374 585
R112 B.n377 B.n72 585
R113 B.n380 B.n379 585
R114 B.n381 B.n71 585
R115 B.n383 B.n382 585
R116 B.n385 B.n70 585
R117 B.n388 B.n387 585
R118 B.n389 B.n69 585
R119 B.n391 B.n390 585
R120 B.n393 B.n68 585
R121 B.n396 B.n395 585
R122 B.n397 B.n67 585
R123 B.n399 B.n398 585
R124 B.n401 B.n66 585
R125 B.n404 B.n403 585
R126 B.n406 B.n63 585
R127 B.n408 B.n407 585
R128 B.n410 B.n62 585
R129 B.n413 B.n412 585
R130 B.n414 B.n61 585
R131 B.n416 B.n415 585
R132 B.n418 B.n60 585
R133 B.n421 B.n420 585
R134 B.n422 B.n56 585
R135 B.n424 B.n423 585
R136 B.n426 B.n55 585
R137 B.n429 B.n428 585
R138 B.n430 B.n54 585
R139 B.n432 B.n431 585
R140 B.n434 B.n53 585
R141 B.n437 B.n436 585
R142 B.n438 B.n52 585
R143 B.n440 B.n439 585
R144 B.n442 B.n51 585
R145 B.n445 B.n444 585
R146 B.n446 B.n50 585
R147 B.n448 B.n447 585
R148 B.n450 B.n49 585
R149 B.n453 B.n452 585
R150 B.n454 B.n48 585
R151 B.n456 B.n455 585
R152 B.n458 B.n47 585
R153 B.n461 B.n460 585
R154 B.n462 B.n46 585
R155 B.n464 B.n463 585
R156 B.n466 B.n45 585
R157 B.n469 B.n468 585
R158 B.n470 B.n44 585
R159 B.n357 B.n42 585
R160 B.n473 B.n42 585
R161 B.n356 B.n41 585
R162 B.n474 B.n41 585
R163 B.n355 B.n40 585
R164 B.n475 B.n40 585
R165 B.n354 B.n353 585
R166 B.n353 B.n36 585
R167 B.n352 B.n35 585
R168 B.n481 B.n35 585
R169 B.n351 B.n34 585
R170 B.n482 B.n34 585
R171 B.n350 B.n33 585
R172 B.n483 B.n33 585
R173 B.n349 B.n348 585
R174 B.n348 B.n29 585
R175 B.n347 B.n28 585
R176 B.n489 B.n28 585
R177 B.n346 B.n27 585
R178 B.n490 B.n27 585
R179 B.n345 B.n26 585
R180 B.n491 B.n26 585
R181 B.n344 B.n343 585
R182 B.n343 B.n22 585
R183 B.n342 B.n21 585
R184 B.n497 B.n21 585
R185 B.n341 B.n20 585
R186 B.n498 B.n20 585
R187 B.n340 B.n19 585
R188 B.n499 B.n19 585
R189 B.n339 B.n338 585
R190 B.n338 B.n15 585
R191 B.n337 B.n14 585
R192 B.n505 B.n14 585
R193 B.n336 B.n13 585
R194 B.n506 B.n13 585
R195 B.n335 B.n12 585
R196 B.n507 B.n12 585
R197 B.n334 B.n333 585
R198 B.n333 B.n11 585
R199 B.n332 B.n7 585
R200 B.n513 B.n7 585
R201 B.n331 B.n6 585
R202 B.n514 B.n6 585
R203 B.n330 B.n5 585
R204 B.n515 B.n5 585
R205 B.n329 B.n328 585
R206 B.n328 B.n4 585
R207 B.n327 B.n77 585
R208 B.n327 B.n326 585
R209 B.n316 B.n78 585
R210 B.n319 B.n78 585
R211 B.n318 B.n317 585
R212 B.n320 B.n318 585
R213 B.n315 B.n83 585
R214 B.n83 B.n82 585
R215 B.n314 B.n313 585
R216 B.n313 B.n312 585
R217 B.n85 B.n84 585
R218 B.n86 B.n85 585
R219 B.n305 B.n304 585
R220 B.n306 B.n305 585
R221 B.n303 B.n91 585
R222 B.n91 B.n90 585
R223 B.n302 B.n301 585
R224 B.n301 B.n300 585
R225 B.n93 B.n92 585
R226 B.n94 B.n93 585
R227 B.n293 B.n292 585
R228 B.n294 B.n293 585
R229 B.n291 B.n98 585
R230 B.n102 B.n98 585
R231 B.n290 B.n289 585
R232 B.n289 B.n288 585
R233 B.n100 B.n99 585
R234 B.n101 B.n100 585
R235 B.n281 B.n280 585
R236 B.n282 B.n281 585
R237 B.n279 B.n107 585
R238 B.n107 B.n106 585
R239 B.n278 B.n277 585
R240 B.n277 B.n276 585
R241 B.n109 B.n108 585
R242 B.n110 B.n109 585
R243 B.n269 B.n268 585
R244 B.n270 B.n269 585
R245 B.n267 B.n115 585
R246 B.n115 B.n114 585
R247 B.n266 B.n265 585
R248 B.n265 B.n264 585
R249 B.n261 B.n119 585
R250 B.n260 B.n259 585
R251 B.n257 B.n120 585
R252 B.n257 B.n118 585
R253 B.n256 B.n255 585
R254 B.n254 B.n253 585
R255 B.n252 B.n122 585
R256 B.n250 B.n249 585
R257 B.n248 B.n123 585
R258 B.n247 B.n246 585
R259 B.n244 B.n124 585
R260 B.n242 B.n241 585
R261 B.n240 B.n125 585
R262 B.n239 B.n238 585
R263 B.n236 B.n126 585
R264 B.n234 B.n233 585
R265 B.n232 B.n127 585
R266 B.n231 B.n230 585
R267 B.n228 B.n128 585
R268 B.n226 B.n225 585
R269 B.n224 B.n129 585
R270 B.n223 B.n222 585
R271 B.n220 B.n130 585
R272 B.n218 B.n217 585
R273 B.n215 B.n131 585
R274 B.n214 B.n213 585
R275 B.n211 B.n134 585
R276 B.n209 B.n208 585
R277 B.n207 B.n135 585
R278 B.n206 B.n205 585
R279 B.n203 B.n136 585
R280 B.n201 B.n200 585
R281 B.n199 B.n137 585
R282 B.n198 B.n197 585
R283 B.n195 B.n194 585
R284 B.n193 B.n192 585
R285 B.n191 B.n142 585
R286 B.n189 B.n188 585
R287 B.n187 B.n143 585
R288 B.n186 B.n185 585
R289 B.n183 B.n144 585
R290 B.n181 B.n180 585
R291 B.n179 B.n145 585
R292 B.n178 B.n177 585
R293 B.n175 B.n146 585
R294 B.n173 B.n172 585
R295 B.n171 B.n147 585
R296 B.n170 B.n169 585
R297 B.n167 B.n148 585
R298 B.n165 B.n164 585
R299 B.n163 B.n149 585
R300 B.n162 B.n161 585
R301 B.n159 B.n150 585
R302 B.n157 B.n156 585
R303 B.n155 B.n151 585
R304 B.n154 B.n153 585
R305 B.n117 B.n116 585
R306 B.n118 B.n117 585
R307 B.n263 B.n262 585
R308 B.n264 B.n263 585
R309 B.n113 B.n112 585
R310 B.n114 B.n113 585
R311 B.n272 B.n271 585
R312 B.n271 B.n270 585
R313 B.n273 B.n111 585
R314 B.n111 B.n110 585
R315 B.n275 B.n274 585
R316 B.n276 B.n275 585
R317 B.n105 B.n104 585
R318 B.n106 B.n105 585
R319 B.n284 B.n283 585
R320 B.n283 B.n282 585
R321 B.n285 B.n103 585
R322 B.n103 B.n101 585
R323 B.n287 B.n286 585
R324 B.n288 B.n287 585
R325 B.n97 B.n96 585
R326 B.n102 B.n97 585
R327 B.n296 B.n295 585
R328 B.n295 B.n294 585
R329 B.n297 B.n95 585
R330 B.n95 B.n94 585
R331 B.n299 B.n298 585
R332 B.n300 B.n299 585
R333 B.n89 B.n88 585
R334 B.n90 B.n89 585
R335 B.n308 B.n307 585
R336 B.n307 B.n306 585
R337 B.n309 B.n87 585
R338 B.n87 B.n86 585
R339 B.n311 B.n310 585
R340 B.n312 B.n311 585
R341 B.n81 B.n80 585
R342 B.n82 B.n81 585
R343 B.n322 B.n321 585
R344 B.n321 B.n320 585
R345 B.n323 B.n79 585
R346 B.n319 B.n79 585
R347 B.n325 B.n324 585
R348 B.n326 B.n325 585
R349 B.n2 B.n0 585
R350 B.n4 B.n2 585
R351 B.n3 B.n1 585
R352 B.n514 B.n3 585
R353 B.n512 B.n511 585
R354 B.n513 B.n512 585
R355 B.n510 B.n8 585
R356 B.n11 B.n8 585
R357 B.n509 B.n508 585
R358 B.n508 B.n507 585
R359 B.n10 B.n9 585
R360 B.n506 B.n10 585
R361 B.n504 B.n503 585
R362 B.n505 B.n504 585
R363 B.n502 B.n16 585
R364 B.n16 B.n15 585
R365 B.n501 B.n500 585
R366 B.n500 B.n499 585
R367 B.n18 B.n17 585
R368 B.n498 B.n18 585
R369 B.n496 B.n495 585
R370 B.n497 B.n496 585
R371 B.n494 B.n23 585
R372 B.n23 B.n22 585
R373 B.n493 B.n492 585
R374 B.n492 B.n491 585
R375 B.n25 B.n24 585
R376 B.n490 B.n25 585
R377 B.n488 B.n487 585
R378 B.n489 B.n488 585
R379 B.n486 B.n30 585
R380 B.n30 B.n29 585
R381 B.n485 B.n484 585
R382 B.n484 B.n483 585
R383 B.n32 B.n31 585
R384 B.n482 B.n32 585
R385 B.n480 B.n479 585
R386 B.n481 B.n480 585
R387 B.n478 B.n37 585
R388 B.n37 B.n36 585
R389 B.n477 B.n476 585
R390 B.n476 B.n475 585
R391 B.n39 B.n38 585
R392 B.n474 B.n39 585
R393 B.n472 B.n471 585
R394 B.n473 B.n472 585
R395 B.n517 B.n516 585
R396 B.n516 B.n515 585
R397 B.n263 B.n119 511.721
R398 B.n472 B.n44 511.721
R399 B.n265 B.n117 511.721
R400 B.n359 B.n42 511.721
R401 B.n138 B.t9 508.705
R402 B.n132 B.t16 508.705
R403 B.n57 B.t13 508.705
R404 B.n64 B.t5 508.705
R405 B.n360 B.n43 256.663
R406 B.n362 B.n43 256.663
R407 B.n368 B.n43 256.663
R408 B.n370 B.n43 256.663
R409 B.n376 B.n43 256.663
R410 B.n378 B.n43 256.663
R411 B.n384 B.n43 256.663
R412 B.n386 B.n43 256.663
R413 B.n392 B.n43 256.663
R414 B.n394 B.n43 256.663
R415 B.n400 B.n43 256.663
R416 B.n402 B.n43 256.663
R417 B.n409 B.n43 256.663
R418 B.n411 B.n43 256.663
R419 B.n417 B.n43 256.663
R420 B.n419 B.n43 256.663
R421 B.n425 B.n43 256.663
R422 B.n427 B.n43 256.663
R423 B.n433 B.n43 256.663
R424 B.n435 B.n43 256.663
R425 B.n441 B.n43 256.663
R426 B.n443 B.n43 256.663
R427 B.n449 B.n43 256.663
R428 B.n451 B.n43 256.663
R429 B.n457 B.n43 256.663
R430 B.n459 B.n43 256.663
R431 B.n465 B.n43 256.663
R432 B.n467 B.n43 256.663
R433 B.n258 B.n118 256.663
R434 B.n121 B.n118 256.663
R435 B.n251 B.n118 256.663
R436 B.n245 B.n118 256.663
R437 B.n243 B.n118 256.663
R438 B.n237 B.n118 256.663
R439 B.n235 B.n118 256.663
R440 B.n229 B.n118 256.663
R441 B.n227 B.n118 256.663
R442 B.n221 B.n118 256.663
R443 B.n219 B.n118 256.663
R444 B.n212 B.n118 256.663
R445 B.n210 B.n118 256.663
R446 B.n204 B.n118 256.663
R447 B.n202 B.n118 256.663
R448 B.n196 B.n118 256.663
R449 B.n141 B.n118 256.663
R450 B.n190 B.n118 256.663
R451 B.n184 B.n118 256.663
R452 B.n182 B.n118 256.663
R453 B.n176 B.n118 256.663
R454 B.n174 B.n118 256.663
R455 B.n168 B.n118 256.663
R456 B.n166 B.n118 256.663
R457 B.n160 B.n118 256.663
R458 B.n158 B.n118 256.663
R459 B.n152 B.n118 256.663
R460 B.n263 B.n113 163.367
R461 B.n271 B.n113 163.367
R462 B.n271 B.n111 163.367
R463 B.n275 B.n111 163.367
R464 B.n275 B.n105 163.367
R465 B.n283 B.n105 163.367
R466 B.n283 B.n103 163.367
R467 B.n287 B.n103 163.367
R468 B.n287 B.n97 163.367
R469 B.n295 B.n97 163.367
R470 B.n295 B.n95 163.367
R471 B.n299 B.n95 163.367
R472 B.n299 B.n89 163.367
R473 B.n307 B.n89 163.367
R474 B.n307 B.n87 163.367
R475 B.n311 B.n87 163.367
R476 B.n311 B.n81 163.367
R477 B.n321 B.n81 163.367
R478 B.n321 B.n79 163.367
R479 B.n325 B.n79 163.367
R480 B.n325 B.n2 163.367
R481 B.n516 B.n2 163.367
R482 B.n516 B.n3 163.367
R483 B.n512 B.n3 163.367
R484 B.n512 B.n8 163.367
R485 B.n508 B.n8 163.367
R486 B.n508 B.n10 163.367
R487 B.n504 B.n10 163.367
R488 B.n504 B.n16 163.367
R489 B.n500 B.n16 163.367
R490 B.n500 B.n18 163.367
R491 B.n496 B.n18 163.367
R492 B.n496 B.n23 163.367
R493 B.n492 B.n23 163.367
R494 B.n492 B.n25 163.367
R495 B.n488 B.n25 163.367
R496 B.n488 B.n30 163.367
R497 B.n484 B.n30 163.367
R498 B.n484 B.n32 163.367
R499 B.n480 B.n32 163.367
R500 B.n480 B.n37 163.367
R501 B.n476 B.n37 163.367
R502 B.n476 B.n39 163.367
R503 B.n472 B.n39 163.367
R504 B.n259 B.n257 163.367
R505 B.n257 B.n256 163.367
R506 B.n253 B.n252 163.367
R507 B.n250 B.n123 163.367
R508 B.n246 B.n244 163.367
R509 B.n242 B.n125 163.367
R510 B.n238 B.n236 163.367
R511 B.n234 B.n127 163.367
R512 B.n230 B.n228 163.367
R513 B.n226 B.n129 163.367
R514 B.n222 B.n220 163.367
R515 B.n218 B.n131 163.367
R516 B.n213 B.n211 163.367
R517 B.n209 B.n135 163.367
R518 B.n205 B.n203 163.367
R519 B.n201 B.n137 163.367
R520 B.n197 B.n195 163.367
R521 B.n192 B.n191 163.367
R522 B.n189 B.n143 163.367
R523 B.n185 B.n183 163.367
R524 B.n181 B.n145 163.367
R525 B.n177 B.n175 163.367
R526 B.n173 B.n147 163.367
R527 B.n169 B.n167 163.367
R528 B.n165 B.n149 163.367
R529 B.n161 B.n159 163.367
R530 B.n157 B.n151 163.367
R531 B.n153 B.n117 163.367
R532 B.n265 B.n115 163.367
R533 B.n269 B.n115 163.367
R534 B.n269 B.n109 163.367
R535 B.n277 B.n109 163.367
R536 B.n277 B.n107 163.367
R537 B.n281 B.n107 163.367
R538 B.n281 B.n100 163.367
R539 B.n289 B.n100 163.367
R540 B.n289 B.n98 163.367
R541 B.n293 B.n98 163.367
R542 B.n293 B.n93 163.367
R543 B.n301 B.n93 163.367
R544 B.n301 B.n91 163.367
R545 B.n305 B.n91 163.367
R546 B.n305 B.n85 163.367
R547 B.n313 B.n85 163.367
R548 B.n313 B.n83 163.367
R549 B.n318 B.n83 163.367
R550 B.n318 B.n78 163.367
R551 B.n327 B.n78 163.367
R552 B.n328 B.n327 163.367
R553 B.n328 B.n5 163.367
R554 B.n6 B.n5 163.367
R555 B.n7 B.n6 163.367
R556 B.n333 B.n7 163.367
R557 B.n333 B.n12 163.367
R558 B.n13 B.n12 163.367
R559 B.n14 B.n13 163.367
R560 B.n338 B.n14 163.367
R561 B.n338 B.n19 163.367
R562 B.n20 B.n19 163.367
R563 B.n21 B.n20 163.367
R564 B.n343 B.n21 163.367
R565 B.n343 B.n26 163.367
R566 B.n27 B.n26 163.367
R567 B.n28 B.n27 163.367
R568 B.n348 B.n28 163.367
R569 B.n348 B.n33 163.367
R570 B.n34 B.n33 163.367
R571 B.n35 B.n34 163.367
R572 B.n353 B.n35 163.367
R573 B.n353 B.n40 163.367
R574 B.n41 B.n40 163.367
R575 B.n42 B.n41 163.367
R576 B.n468 B.n466 163.367
R577 B.n464 B.n46 163.367
R578 B.n460 B.n458 163.367
R579 B.n456 B.n48 163.367
R580 B.n452 B.n450 163.367
R581 B.n448 B.n50 163.367
R582 B.n444 B.n442 163.367
R583 B.n440 B.n52 163.367
R584 B.n436 B.n434 163.367
R585 B.n432 B.n54 163.367
R586 B.n428 B.n426 163.367
R587 B.n424 B.n56 163.367
R588 B.n420 B.n418 163.367
R589 B.n416 B.n61 163.367
R590 B.n412 B.n410 163.367
R591 B.n408 B.n63 163.367
R592 B.n403 B.n401 163.367
R593 B.n399 B.n67 163.367
R594 B.n395 B.n393 163.367
R595 B.n391 B.n69 163.367
R596 B.n387 B.n385 163.367
R597 B.n383 B.n71 163.367
R598 B.n379 B.n377 163.367
R599 B.n375 B.n73 163.367
R600 B.n371 B.n369 163.367
R601 B.n367 B.n75 163.367
R602 B.n363 B.n361 163.367
R603 B.n264 B.n118 126.713
R604 B.n473 B.n43 126.713
R605 B.n138 B.t12 90.9412
R606 B.n64 B.t7 90.9412
R607 B.n132 B.t18 90.9354
R608 B.n57 B.t14 90.9354
R609 B.n139 B.t11 75.62
R610 B.n65 B.t8 75.62
R611 B.n133 B.t17 75.6142
R612 B.n58 B.t15 75.6142
R613 B.n258 B.n119 71.676
R614 B.n256 B.n121 71.676
R615 B.n252 B.n251 71.676
R616 B.n245 B.n123 71.676
R617 B.n244 B.n243 71.676
R618 B.n237 B.n125 71.676
R619 B.n236 B.n235 71.676
R620 B.n229 B.n127 71.676
R621 B.n228 B.n227 71.676
R622 B.n221 B.n129 71.676
R623 B.n220 B.n219 71.676
R624 B.n212 B.n131 71.676
R625 B.n211 B.n210 71.676
R626 B.n204 B.n135 71.676
R627 B.n203 B.n202 71.676
R628 B.n196 B.n137 71.676
R629 B.n195 B.n141 71.676
R630 B.n191 B.n190 71.676
R631 B.n184 B.n143 71.676
R632 B.n183 B.n182 71.676
R633 B.n176 B.n145 71.676
R634 B.n175 B.n174 71.676
R635 B.n168 B.n147 71.676
R636 B.n167 B.n166 71.676
R637 B.n160 B.n149 71.676
R638 B.n159 B.n158 71.676
R639 B.n152 B.n151 71.676
R640 B.n467 B.n44 71.676
R641 B.n466 B.n465 71.676
R642 B.n459 B.n46 71.676
R643 B.n458 B.n457 71.676
R644 B.n451 B.n48 71.676
R645 B.n450 B.n449 71.676
R646 B.n443 B.n50 71.676
R647 B.n442 B.n441 71.676
R648 B.n435 B.n52 71.676
R649 B.n434 B.n433 71.676
R650 B.n427 B.n54 71.676
R651 B.n426 B.n425 71.676
R652 B.n419 B.n56 71.676
R653 B.n418 B.n417 71.676
R654 B.n411 B.n61 71.676
R655 B.n410 B.n409 71.676
R656 B.n402 B.n63 71.676
R657 B.n401 B.n400 71.676
R658 B.n394 B.n67 71.676
R659 B.n393 B.n392 71.676
R660 B.n386 B.n69 71.676
R661 B.n385 B.n384 71.676
R662 B.n378 B.n71 71.676
R663 B.n377 B.n376 71.676
R664 B.n370 B.n73 71.676
R665 B.n369 B.n368 71.676
R666 B.n362 B.n75 71.676
R667 B.n361 B.n360 71.676
R668 B.n360 B.n359 71.676
R669 B.n363 B.n362 71.676
R670 B.n368 B.n367 71.676
R671 B.n371 B.n370 71.676
R672 B.n376 B.n375 71.676
R673 B.n379 B.n378 71.676
R674 B.n384 B.n383 71.676
R675 B.n387 B.n386 71.676
R676 B.n392 B.n391 71.676
R677 B.n395 B.n394 71.676
R678 B.n400 B.n399 71.676
R679 B.n403 B.n402 71.676
R680 B.n409 B.n408 71.676
R681 B.n412 B.n411 71.676
R682 B.n417 B.n416 71.676
R683 B.n420 B.n419 71.676
R684 B.n425 B.n424 71.676
R685 B.n428 B.n427 71.676
R686 B.n433 B.n432 71.676
R687 B.n436 B.n435 71.676
R688 B.n441 B.n440 71.676
R689 B.n444 B.n443 71.676
R690 B.n449 B.n448 71.676
R691 B.n452 B.n451 71.676
R692 B.n457 B.n456 71.676
R693 B.n460 B.n459 71.676
R694 B.n465 B.n464 71.676
R695 B.n468 B.n467 71.676
R696 B.n259 B.n258 71.676
R697 B.n253 B.n121 71.676
R698 B.n251 B.n250 71.676
R699 B.n246 B.n245 71.676
R700 B.n243 B.n242 71.676
R701 B.n238 B.n237 71.676
R702 B.n235 B.n234 71.676
R703 B.n230 B.n229 71.676
R704 B.n227 B.n226 71.676
R705 B.n222 B.n221 71.676
R706 B.n219 B.n218 71.676
R707 B.n213 B.n212 71.676
R708 B.n210 B.n209 71.676
R709 B.n205 B.n204 71.676
R710 B.n202 B.n201 71.676
R711 B.n197 B.n196 71.676
R712 B.n192 B.n141 71.676
R713 B.n190 B.n189 71.676
R714 B.n185 B.n184 71.676
R715 B.n182 B.n181 71.676
R716 B.n177 B.n176 71.676
R717 B.n174 B.n173 71.676
R718 B.n169 B.n168 71.676
R719 B.n166 B.n165 71.676
R720 B.n161 B.n160 71.676
R721 B.n158 B.n157 71.676
R722 B.n153 B.n152 71.676
R723 B.n264 B.n114 67.8463
R724 B.n270 B.n114 67.8463
R725 B.n270 B.n110 67.8463
R726 B.n276 B.n110 67.8463
R727 B.n282 B.n106 67.8463
R728 B.n282 B.n101 67.8463
R729 B.n288 B.n101 67.8463
R730 B.n288 B.n102 67.8463
R731 B.n294 B.n94 67.8463
R732 B.n300 B.n94 67.8463
R733 B.n306 B.n90 67.8463
R734 B.n312 B.n86 67.8463
R735 B.n320 B.n82 67.8463
R736 B.n320 B.n319 67.8463
R737 B.n326 B.n4 67.8463
R738 B.n515 B.n4 67.8463
R739 B.n515 B.n514 67.8463
R740 B.n514 B.n513 67.8463
R741 B.n507 B.n11 67.8463
R742 B.n507 B.n506 67.8463
R743 B.n505 B.n15 67.8463
R744 B.n499 B.n498 67.8463
R745 B.n497 B.n22 67.8463
R746 B.n491 B.n22 67.8463
R747 B.n490 B.n489 67.8463
R748 B.n489 B.n29 67.8463
R749 B.n483 B.n29 67.8463
R750 B.n483 B.n482 67.8463
R751 B.n481 B.n36 67.8463
R752 B.n475 B.n36 67.8463
R753 B.n475 B.n474 67.8463
R754 B.n474 B.n473 67.8463
R755 B.n102 B.t22 63.8554
R756 B.t23 B.n490 63.8554
R757 B.n312 B.t19 61.8599
R758 B.t0 B.n505 61.8599
R759 B.n140 B.n139 59.5399
R760 B.n216 B.n133 59.5399
R761 B.n59 B.n58 59.5399
R762 B.n405 B.n65 59.5399
R763 B.n326 B.t1 51.8826
R764 B.n513 B.t4 51.8826
R765 B.t20 B.n90 49.8871
R766 B.n498 B.t3 49.8871
R767 B.t10 B.n106 39.9098
R768 B.n306 B.t2 39.9098
R769 B.n499 B.t21 39.9098
R770 B.n482 B.t6 39.9098
R771 B.n471 B.n470 33.2493
R772 B.n358 B.n357 33.2493
R773 B.n266 B.n116 33.2493
R774 B.n262 B.n261 33.2493
R775 B.n276 B.t10 27.937
R776 B.t2 B.n86 27.937
R777 B.t21 B.n15 27.937
R778 B.t6 B.n481 27.937
R779 B B.n517 18.0485
R780 B.n300 B.t20 17.9597
R781 B.t3 B.n497 17.9597
R782 B.n319 B.t1 15.9642
R783 B.n11 B.t4 15.9642
R784 B.n139 B.n138 15.3217
R785 B.n133 B.n132 15.3217
R786 B.n58 B.n57 15.3217
R787 B.n65 B.n64 15.3217
R788 B.n470 B.n469 10.6151
R789 B.n469 B.n45 10.6151
R790 B.n463 B.n45 10.6151
R791 B.n463 B.n462 10.6151
R792 B.n462 B.n461 10.6151
R793 B.n461 B.n47 10.6151
R794 B.n455 B.n47 10.6151
R795 B.n455 B.n454 10.6151
R796 B.n454 B.n453 10.6151
R797 B.n453 B.n49 10.6151
R798 B.n447 B.n49 10.6151
R799 B.n447 B.n446 10.6151
R800 B.n446 B.n445 10.6151
R801 B.n445 B.n51 10.6151
R802 B.n439 B.n51 10.6151
R803 B.n439 B.n438 10.6151
R804 B.n438 B.n437 10.6151
R805 B.n437 B.n53 10.6151
R806 B.n431 B.n53 10.6151
R807 B.n431 B.n430 10.6151
R808 B.n430 B.n429 10.6151
R809 B.n429 B.n55 10.6151
R810 B.n423 B.n422 10.6151
R811 B.n422 B.n421 10.6151
R812 B.n421 B.n60 10.6151
R813 B.n415 B.n60 10.6151
R814 B.n415 B.n414 10.6151
R815 B.n414 B.n413 10.6151
R816 B.n413 B.n62 10.6151
R817 B.n407 B.n62 10.6151
R818 B.n407 B.n406 10.6151
R819 B.n404 B.n66 10.6151
R820 B.n398 B.n66 10.6151
R821 B.n398 B.n397 10.6151
R822 B.n397 B.n396 10.6151
R823 B.n396 B.n68 10.6151
R824 B.n390 B.n68 10.6151
R825 B.n390 B.n389 10.6151
R826 B.n389 B.n388 10.6151
R827 B.n388 B.n70 10.6151
R828 B.n382 B.n70 10.6151
R829 B.n382 B.n381 10.6151
R830 B.n381 B.n380 10.6151
R831 B.n380 B.n72 10.6151
R832 B.n374 B.n72 10.6151
R833 B.n374 B.n373 10.6151
R834 B.n373 B.n372 10.6151
R835 B.n372 B.n74 10.6151
R836 B.n366 B.n74 10.6151
R837 B.n366 B.n365 10.6151
R838 B.n365 B.n364 10.6151
R839 B.n364 B.n76 10.6151
R840 B.n358 B.n76 10.6151
R841 B.n267 B.n266 10.6151
R842 B.n268 B.n267 10.6151
R843 B.n268 B.n108 10.6151
R844 B.n278 B.n108 10.6151
R845 B.n279 B.n278 10.6151
R846 B.n280 B.n279 10.6151
R847 B.n280 B.n99 10.6151
R848 B.n290 B.n99 10.6151
R849 B.n291 B.n290 10.6151
R850 B.n292 B.n291 10.6151
R851 B.n292 B.n92 10.6151
R852 B.n302 B.n92 10.6151
R853 B.n303 B.n302 10.6151
R854 B.n304 B.n303 10.6151
R855 B.n304 B.n84 10.6151
R856 B.n314 B.n84 10.6151
R857 B.n315 B.n314 10.6151
R858 B.n317 B.n315 10.6151
R859 B.n317 B.n316 10.6151
R860 B.n316 B.n77 10.6151
R861 B.n329 B.n77 10.6151
R862 B.n330 B.n329 10.6151
R863 B.n331 B.n330 10.6151
R864 B.n332 B.n331 10.6151
R865 B.n334 B.n332 10.6151
R866 B.n335 B.n334 10.6151
R867 B.n336 B.n335 10.6151
R868 B.n337 B.n336 10.6151
R869 B.n339 B.n337 10.6151
R870 B.n340 B.n339 10.6151
R871 B.n341 B.n340 10.6151
R872 B.n342 B.n341 10.6151
R873 B.n344 B.n342 10.6151
R874 B.n345 B.n344 10.6151
R875 B.n346 B.n345 10.6151
R876 B.n347 B.n346 10.6151
R877 B.n349 B.n347 10.6151
R878 B.n350 B.n349 10.6151
R879 B.n351 B.n350 10.6151
R880 B.n352 B.n351 10.6151
R881 B.n354 B.n352 10.6151
R882 B.n355 B.n354 10.6151
R883 B.n356 B.n355 10.6151
R884 B.n357 B.n356 10.6151
R885 B.n261 B.n260 10.6151
R886 B.n260 B.n120 10.6151
R887 B.n255 B.n120 10.6151
R888 B.n255 B.n254 10.6151
R889 B.n254 B.n122 10.6151
R890 B.n249 B.n122 10.6151
R891 B.n249 B.n248 10.6151
R892 B.n248 B.n247 10.6151
R893 B.n247 B.n124 10.6151
R894 B.n241 B.n124 10.6151
R895 B.n241 B.n240 10.6151
R896 B.n240 B.n239 10.6151
R897 B.n239 B.n126 10.6151
R898 B.n233 B.n126 10.6151
R899 B.n233 B.n232 10.6151
R900 B.n232 B.n231 10.6151
R901 B.n231 B.n128 10.6151
R902 B.n225 B.n128 10.6151
R903 B.n225 B.n224 10.6151
R904 B.n224 B.n223 10.6151
R905 B.n223 B.n130 10.6151
R906 B.n217 B.n130 10.6151
R907 B.n215 B.n214 10.6151
R908 B.n214 B.n134 10.6151
R909 B.n208 B.n134 10.6151
R910 B.n208 B.n207 10.6151
R911 B.n207 B.n206 10.6151
R912 B.n206 B.n136 10.6151
R913 B.n200 B.n136 10.6151
R914 B.n200 B.n199 10.6151
R915 B.n199 B.n198 10.6151
R916 B.n194 B.n193 10.6151
R917 B.n193 B.n142 10.6151
R918 B.n188 B.n142 10.6151
R919 B.n188 B.n187 10.6151
R920 B.n187 B.n186 10.6151
R921 B.n186 B.n144 10.6151
R922 B.n180 B.n144 10.6151
R923 B.n180 B.n179 10.6151
R924 B.n179 B.n178 10.6151
R925 B.n178 B.n146 10.6151
R926 B.n172 B.n146 10.6151
R927 B.n172 B.n171 10.6151
R928 B.n171 B.n170 10.6151
R929 B.n170 B.n148 10.6151
R930 B.n164 B.n148 10.6151
R931 B.n164 B.n163 10.6151
R932 B.n163 B.n162 10.6151
R933 B.n162 B.n150 10.6151
R934 B.n156 B.n150 10.6151
R935 B.n156 B.n155 10.6151
R936 B.n155 B.n154 10.6151
R937 B.n154 B.n116 10.6151
R938 B.n262 B.n112 10.6151
R939 B.n272 B.n112 10.6151
R940 B.n273 B.n272 10.6151
R941 B.n274 B.n273 10.6151
R942 B.n274 B.n104 10.6151
R943 B.n284 B.n104 10.6151
R944 B.n285 B.n284 10.6151
R945 B.n286 B.n285 10.6151
R946 B.n286 B.n96 10.6151
R947 B.n296 B.n96 10.6151
R948 B.n297 B.n296 10.6151
R949 B.n298 B.n297 10.6151
R950 B.n298 B.n88 10.6151
R951 B.n308 B.n88 10.6151
R952 B.n309 B.n308 10.6151
R953 B.n310 B.n309 10.6151
R954 B.n310 B.n80 10.6151
R955 B.n322 B.n80 10.6151
R956 B.n323 B.n322 10.6151
R957 B.n324 B.n323 10.6151
R958 B.n324 B.n0 10.6151
R959 B.n511 B.n1 10.6151
R960 B.n511 B.n510 10.6151
R961 B.n510 B.n509 10.6151
R962 B.n509 B.n9 10.6151
R963 B.n503 B.n9 10.6151
R964 B.n503 B.n502 10.6151
R965 B.n502 B.n501 10.6151
R966 B.n501 B.n17 10.6151
R967 B.n495 B.n17 10.6151
R968 B.n495 B.n494 10.6151
R969 B.n494 B.n493 10.6151
R970 B.n493 B.n24 10.6151
R971 B.n487 B.n24 10.6151
R972 B.n487 B.n486 10.6151
R973 B.n486 B.n485 10.6151
R974 B.n485 B.n31 10.6151
R975 B.n479 B.n31 10.6151
R976 B.n479 B.n478 10.6151
R977 B.n478 B.n477 10.6151
R978 B.n477 B.n38 10.6151
R979 B.n471 B.n38 10.6151
R980 B.n59 B.n55 9.36635
R981 B.n405 B.n404 9.36635
R982 B.n217 B.n216 9.36635
R983 B.n194 B.n140 9.36635
R984 B.t19 B.n82 5.98689
R985 B.n506 B.t0 5.98689
R986 B.n294 B.t22 3.99143
R987 B.n491 B.t23 3.99143
R988 B.n517 B.n0 2.81026
R989 B.n517 B.n1 2.81026
R990 B.n423 B.n59 1.24928
R991 B.n406 B.n405 1.24928
R992 B.n216 B.n215 1.24928
R993 B.n198 B.n140 1.24928
R994 VP.n5 VP.t9 408.154
R995 VP.n16 VP.t2 387.173
R996 VP.n17 VP.t1 387.173
R997 VP.n1 VP.t7 387.173
R998 VP.n23 VP.t3 387.173
R999 VP.n24 VP.t0 387.173
R1000 VP.n13 VP.t4 387.173
R1001 VP.n12 VP.t8 387.173
R1002 VP.n4 VP.t6 387.173
R1003 VP.n6 VP.t5 387.173
R1004 VP.n25 VP.n24 161.3
R1005 VP.n8 VP.n7 161.3
R1006 VP.n9 VP.n4 161.3
R1007 VP.n11 VP.n10 161.3
R1008 VP.n12 VP.n3 161.3
R1009 VP.n14 VP.n13 161.3
R1010 VP.n23 VP.n0 161.3
R1011 VP.n22 VP.n21 161.3
R1012 VP.n20 VP.n1 161.3
R1013 VP.n19 VP.n18 161.3
R1014 VP.n17 VP.n2 161.3
R1015 VP.n16 VP.n15 161.3
R1016 VP.n8 VP.n5 70.4033
R1017 VP.n17 VP.n16 48.2005
R1018 VP.n24 VP.n23 48.2005
R1019 VP.n13 VP.n12 48.2005
R1020 VP.n18 VP.n1 39.4369
R1021 VP.n22 VP.n1 39.4369
R1022 VP.n11 VP.n4 39.4369
R1023 VP.n7 VP.n4 39.4369
R1024 VP.n15 VP.n14 36.7013
R1025 VP.n6 VP.n5 20.9576
R1026 VP.n18 VP.n17 8.76414
R1027 VP.n23 VP.n22 8.76414
R1028 VP.n12 VP.n11 8.76414
R1029 VP.n7 VP.n6 8.76414
R1030 VP.n9 VP.n8 0.189894
R1031 VP.n10 VP.n9 0.189894
R1032 VP.n10 VP.n3 0.189894
R1033 VP.n14 VP.n3 0.189894
R1034 VP.n15 VP.n2 0.189894
R1035 VP.n19 VP.n2 0.189894
R1036 VP.n20 VP.n19 0.189894
R1037 VP.n21 VP.n20 0.189894
R1038 VP.n21 VP.n0 0.189894
R1039 VP.n25 VP.n0 0.189894
R1040 VP VP.n25 0.0516364
R1041 VDD1.n1 VDD1.t0 74.1279
R1042 VDD1.n3 VDD1.t7 74.1277
R1043 VDD1.n5 VDD1.n4 70.4586
R1044 VDD1.n1 VDD1.n0 70.0034
R1045 VDD1.n7 VDD1.n6 70.0032
R1046 VDD1.n3 VDD1.n2 70.0031
R1047 VDD1.n7 VDD1.n5 32.8306
R1048 VDD1.n6 VDD1.t1 3.44398
R1049 VDD1.n6 VDD1.t5 3.44398
R1050 VDD1.n0 VDD1.t4 3.44398
R1051 VDD1.n0 VDD1.t3 3.44398
R1052 VDD1.n4 VDD1.t6 3.44398
R1053 VDD1.n4 VDD1.t9 3.44398
R1054 VDD1.n2 VDD1.t8 3.44398
R1055 VDD1.n2 VDD1.t2 3.44398
R1056 VDD1 VDD1.n7 0.453086
R1057 VDD1 VDD1.n1 0.228948
R1058 VDD1.n5 VDD1.n3 0.115413
C0 VTAIL VDD1 9.41275f
C1 VP VDD2 0.310049f
C2 VP VN 4.08993f
C3 VDD2 VDD1 0.821619f
C4 VN VDD1 0.148478f
C5 VDD2 VTAIL 9.44828f
C6 VTAIL VN 2.73957f
C7 VP VDD1 2.88616f
C8 VP VTAIL 2.75396f
C9 VDD2 VN 2.7272f
C10 VDD2 B 3.582324f
C11 VDD1 B 3.485552f
C12 VTAIL B 3.917662f
C13 VN B 7.58692f
C14 VP B 5.852046f
C15 VDD1.t0 B 1.27723f
C16 VDD1.t4 B 0.120679f
C17 VDD1.t3 B 0.120679f
C18 VDD1.n0 B 1.00173f
C19 VDD1.n1 B 0.628689f
C20 VDD1.t7 B 1.27723f
C21 VDD1.t8 B 0.120679f
C22 VDD1.t2 B 0.120679f
C23 VDD1.n2 B 1.00172f
C24 VDD1.n3 B 0.624338f
C25 VDD1.t6 B 0.120679f
C26 VDD1.t9 B 0.120679f
C27 VDD1.n4 B 1.00381f
C28 VDD1.n5 B 1.56103f
C29 VDD1.t1 B 0.120679f
C30 VDD1.t5 B 0.120679f
C31 VDD1.n6 B 1.00172f
C32 VDD1.n7 B 1.89878f
C33 VP.n0 B 0.050683f
C34 VP.t7 B 0.389626f
C35 VP.n1 B 0.193384f
C36 VP.n2 B 0.050683f
C37 VP.n3 B 0.050683f
C38 VP.t4 B 0.389626f
C39 VP.t8 B 0.389626f
C40 VP.t6 B 0.389626f
C41 VP.n4 B 0.193384f
C42 VP.t9 B 0.399233f
C43 VP.n5 B 0.177561f
C44 VP.t5 B 0.389626f
C45 VP.n6 B 0.188697f
C46 VP.n7 B 0.011501f
C47 VP.n8 B 0.155452f
C48 VP.n9 B 0.050683f
C49 VP.n10 B 0.050683f
C50 VP.n11 B 0.011501f
C51 VP.n12 B 0.188697f
C52 VP.n13 B 0.186822f
C53 VP.n14 B 1.65178f
C54 VP.n15 B 1.70142f
C55 VP.t2 B 0.389626f
C56 VP.n16 B 0.186822f
C57 VP.t1 B 0.389626f
C58 VP.n17 B 0.188697f
C59 VP.n18 B 0.011501f
C60 VP.n19 B 0.050683f
C61 VP.n20 B 0.050683f
C62 VP.n21 B 0.050683f
C63 VP.n22 B 0.011501f
C64 VP.t3 B 0.389626f
C65 VP.n23 B 0.188697f
C66 VP.t0 B 0.389626f
C67 VP.n24 B 0.186822f
C68 VP.n25 B 0.039277f
C69 VDD2.t2 B 1.26656f
C70 VDD2.t1 B 0.119671f
C71 VDD2.t6 B 0.119671f
C72 VDD2.n0 B 0.993356f
C73 VDD2.n1 B 0.619124f
C74 VDD2.t0 B 0.119671f
C75 VDD2.t9 B 0.119671f
C76 VDD2.n2 B 0.995429f
C77 VDD2.n3 B 1.47486f
C78 VDD2.t8 B 1.26347f
C79 VDD2.n4 B 1.87664f
C80 VDD2.t5 B 0.119671f
C81 VDD2.t7 B 0.119671f
C82 VDD2.n5 B 0.99336f
C83 VDD2.n6 B 0.289525f
C84 VDD2.t3 B 0.119671f
C85 VDD2.t4 B 0.119671f
C86 VDD2.n7 B 0.995406f
C87 VTAIL.t12 B 0.132668f
C88 VTAIL.t13 B 0.132668f
C89 VTAIL.n0 B 1.02935f
C90 VTAIL.n1 B 0.397384f
C91 VTAIL.t1 B 1.31483f
C92 VTAIL.n2 B 0.484268f
C93 VTAIL.t2 B 0.132668f
C94 VTAIL.t17 B 0.132668f
C95 VTAIL.n3 B 1.02935f
C96 VTAIL.n4 B 0.395762f
C97 VTAIL.t16 B 0.132668f
C98 VTAIL.t15 B 0.132668f
C99 VTAIL.n5 B 1.02935f
C100 VTAIL.n6 B 1.3228f
C101 VTAIL.t11 B 0.132668f
C102 VTAIL.t14 B 0.132668f
C103 VTAIL.n7 B 1.02936f
C104 VTAIL.n8 B 1.32279f
C105 VTAIL.t7 B 0.132668f
C106 VTAIL.t6 B 0.132668f
C107 VTAIL.n9 B 1.02936f
C108 VTAIL.n10 B 0.395756f
C109 VTAIL.t8 B 1.31484f
C110 VTAIL.n11 B 0.484262f
C111 VTAIL.t4 B 0.132668f
C112 VTAIL.t0 B 0.132668f
C113 VTAIL.n12 B 1.02936f
C114 VTAIL.n13 B 0.407922f
C115 VTAIL.t19 B 0.132668f
C116 VTAIL.t3 B 0.132668f
C117 VTAIL.n14 B 1.02936f
C118 VTAIL.n15 B 0.395756f
C119 VTAIL.t18 B 1.31483f
C120 VTAIL.n16 B 1.33506f
C121 VTAIL.t10 B 1.31483f
C122 VTAIL.n17 B 1.33507f
C123 VTAIL.t9 B 0.132668f
C124 VTAIL.t5 B 0.132668f
C125 VTAIL.n18 B 1.02935f
C126 VTAIL.n19 B 0.342233f
C127 VN.n0 B 0.048777f
C128 VN.t3 B 0.374973f
C129 VN.n1 B 0.186111f
C130 VN.t7 B 0.384219f
C131 VN.n2 B 0.170883f
C132 VN.t8 B 0.374973f
C133 VN.n3 B 0.1816f
C134 VN.n4 B 0.011068f
C135 VN.n5 B 0.149605f
C136 VN.n6 B 0.048777f
C137 VN.n7 B 0.048777f
C138 VN.n8 B 0.011068f
C139 VN.t9 B 0.374973f
C140 VN.n9 B 0.1816f
C141 VN.t0 B 0.374973f
C142 VN.n10 B 0.179796f
C143 VN.n11 B 0.0378f
C144 VN.n12 B 0.048777f
C145 VN.t2 B 0.374973f
C146 VN.n13 B 0.186111f
C147 VN.t5 B 0.384219f
C148 VN.n14 B 0.170883f
C149 VN.t6 B 0.374973f
C150 VN.n15 B 0.1816f
C151 VN.n16 B 0.011068f
C152 VN.n17 B 0.149605f
C153 VN.n18 B 0.048777f
C154 VN.n19 B 0.048777f
C155 VN.n20 B 0.011068f
C156 VN.t4 B 0.374973f
C157 VN.n21 B 0.1816f
C158 VN.t1 B 0.374973f
C159 VN.n22 B 0.179796f
C160 VN.n23 B 1.62196f
.ends

