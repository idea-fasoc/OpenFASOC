* NGSPICE file created from diff_pair_sample_0239.ext - technology: sky130A

.subckt diff_pair_sample_0239 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=4.1496 ps=22.06 w=10.64 l=3.16
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=0 ps=0 w=10.64 l=3.16
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=4.1496 ps=22.06 w=10.64 l=3.16
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=0 ps=0 w=10.64 l=3.16
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=4.1496 ps=22.06 w=10.64 l=3.16
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=0 ps=0 w=10.64 l=3.16
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=0 ps=0 w=10.64 l=3.16
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1496 pd=22.06 as=4.1496 ps=22.06 w=10.64 l=3.16
R0 VP.n0 VP.t0 164.988
R1 VP.n0 VP.t1 119.877
R2 VP VP.n0 0.526368
R3 VTAIL.n226 VTAIL.n174 289.615
R4 VTAIL.n52 VTAIL.n0 289.615
R5 VTAIL.n168 VTAIL.n116 289.615
R6 VTAIL.n110 VTAIL.n58 289.615
R7 VTAIL.n193 VTAIL.n192 185
R8 VTAIL.n190 VTAIL.n189 185
R9 VTAIL.n199 VTAIL.n198 185
R10 VTAIL.n201 VTAIL.n200 185
R11 VTAIL.n186 VTAIL.n185 185
R12 VTAIL.n207 VTAIL.n206 185
R13 VTAIL.n210 VTAIL.n209 185
R14 VTAIL.n208 VTAIL.n182 185
R15 VTAIL.n215 VTAIL.n181 185
R16 VTAIL.n217 VTAIL.n216 185
R17 VTAIL.n219 VTAIL.n218 185
R18 VTAIL.n178 VTAIL.n177 185
R19 VTAIL.n225 VTAIL.n224 185
R20 VTAIL.n227 VTAIL.n226 185
R21 VTAIL.n19 VTAIL.n18 185
R22 VTAIL.n16 VTAIL.n15 185
R23 VTAIL.n25 VTAIL.n24 185
R24 VTAIL.n27 VTAIL.n26 185
R25 VTAIL.n12 VTAIL.n11 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n36 VTAIL.n35 185
R28 VTAIL.n34 VTAIL.n8 185
R29 VTAIL.n41 VTAIL.n7 185
R30 VTAIL.n43 VTAIL.n42 185
R31 VTAIL.n45 VTAIL.n44 185
R32 VTAIL.n4 VTAIL.n3 185
R33 VTAIL.n51 VTAIL.n50 185
R34 VTAIL.n53 VTAIL.n52 185
R35 VTAIL.n169 VTAIL.n168 185
R36 VTAIL.n167 VTAIL.n166 185
R37 VTAIL.n120 VTAIL.n119 185
R38 VTAIL.n161 VTAIL.n160 185
R39 VTAIL.n159 VTAIL.n158 185
R40 VTAIL.n157 VTAIL.n123 185
R41 VTAIL.n127 VTAIL.n124 185
R42 VTAIL.n152 VTAIL.n151 185
R43 VTAIL.n150 VTAIL.n149 185
R44 VTAIL.n129 VTAIL.n128 185
R45 VTAIL.n144 VTAIL.n143 185
R46 VTAIL.n142 VTAIL.n141 185
R47 VTAIL.n133 VTAIL.n132 185
R48 VTAIL.n136 VTAIL.n135 185
R49 VTAIL.n111 VTAIL.n110 185
R50 VTAIL.n109 VTAIL.n108 185
R51 VTAIL.n62 VTAIL.n61 185
R52 VTAIL.n103 VTAIL.n102 185
R53 VTAIL.n101 VTAIL.n100 185
R54 VTAIL.n99 VTAIL.n65 185
R55 VTAIL.n69 VTAIL.n66 185
R56 VTAIL.n94 VTAIL.n93 185
R57 VTAIL.n92 VTAIL.n91 185
R58 VTAIL.n71 VTAIL.n70 185
R59 VTAIL.n86 VTAIL.n85 185
R60 VTAIL.n84 VTAIL.n83 185
R61 VTAIL.n75 VTAIL.n74 185
R62 VTAIL.n78 VTAIL.n77 185
R63 VTAIL.t0 VTAIL.n191 149.524
R64 VTAIL.t3 VTAIL.n17 149.524
R65 VTAIL.t2 VTAIL.n134 149.524
R66 VTAIL.t1 VTAIL.n76 149.524
R67 VTAIL.n192 VTAIL.n189 104.615
R68 VTAIL.n199 VTAIL.n189 104.615
R69 VTAIL.n200 VTAIL.n199 104.615
R70 VTAIL.n200 VTAIL.n185 104.615
R71 VTAIL.n207 VTAIL.n185 104.615
R72 VTAIL.n209 VTAIL.n207 104.615
R73 VTAIL.n209 VTAIL.n208 104.615
R74 VTAIL.n208 VTAIL.n181 104.615
R75 VTAIL.n217 VTAIL.n181 104.615
R76 VTAIL.n218 VTAIL.n217 104.615
R77 VTAIL.n218 VTAIL.n177 104.615
R78 VTAIL.n225 VTAIL.n177 104.615
R79 VTAIL.n226 VTAIL.n225 104.615
R80 VTAIL.n18 VTAIL.n15 104.615
R81 VTAIL.n25 VTAIL.n15 104.615
R82 VTAIL.n26 VTAIL.n25 104.615
R83 VTAIL.n26 VTAIL.n11 104.615
R84 VTAIL.n33 VTAIL.n11 104.615
R85 VTAIL.n35 VTAIL.n33 104.615
R86 VTAIL.n35 VTAIL.n34 104.615
R87 VTAIL.n34 VTAIL.n7 104.615
R88 VTAIL.n43 VTAIL.n7 104.615
R89 VTAIL.n44 VTAIL.n43 104.615
R90 VTAIL.n44 VTAIL.n3 104.615
R91 VTAIL.n51 VTAIL.n3 104.615
R92 VTAIL.n52 VTAIL.n51 104.615
R93 VTAIL.n168 VTAIL.n167 104.615
R94 VTAIL.n167 VTAIL.n119 104.615
R95 VTAIL.n160 VTAIL.n119 104.615
R96 VTAIL.n160 VTAIL.n159 104.615
R97 VTAIL.n159 VTAIL.n123 104.615
R98 VTAIL.n127 VTAIL.n123 104.615
R99 VTAIL.n151 VTAIL.n127 104.615
R100 VTAIL.n151 VTAIL.n150 104.615
R101 VTAIL.n150 VTAIL.n128 104.615
R102 VTAIL.n143 VTAIL.n128 104.615
R103 VTAIL.n143 VTAIL.n142 104.615
R104 VTAIL.n142 VTAIL.n132 104.615
R105 VTAIL.n135 VTAIL.n132 104.615
R106 VTAIL.n110 VTAIL.n109 104.615
R107 VTAIL.n109 VTAIL.n61 104.615
R108 VTAIL.n102 VTAIL.n61 104.615
R109 VTAIL.n102 VTAIL.n101 104.615
R110 VTAIL.n101 VTAIL.n65 104.615
R111 VTAIL.n69 VTAIL.n65 104.615
R112 VTAIL.n93 VTAIL.n69 104.615
R113 VTAIL.n93 VTAIL.n92 104.615
R114 VTAIL.n92 VTAIL.n70 104.615
R115 VTAIL.n85 VTAIL.n70 104.615
R116 VTAIL.n85 VTAIL.n84 104.615
R117 VTAIL.n84 VTAIL.n74 104.615
R118 VTAIL.n77 VTAIL.n74 104.615
R119 VTAIL.n192 VTAIL.t0 52.3082
R120 VTAIL.n18 VTAIL.t3 52.3082
R121 VTAIL.n135 VTAIL.t2 52.3082
R122 VTAIL.n77 VTAIL.t1 52.3082
R123 VTAIL.n231 VTAIL.n230 31.4096
R124 VTAIL.n57 VTAIL.n56 31.4096
R125 VTAIL.n173 VTAIL.n172 31.4096
R126 VTAIL.n115 VTAIL.n114 31.4096
R127 VTAIL.n115 VTAIL.n57 27.5565
R128 VTAIL.n231 VTAIL.n173 24.5479
R129 VTAIL.n216 VTAIL.n215 13.1884
R130 VTAIL.n42 VTAIL.n41 13.1884
R131 VTAIL.n158 VTAIL.n157 13.1884
R132 VTAIL.n100 VTAIL.n99 13.1884
R133 VTAIL.n214 VTAIL.n182 12.8005
R134 VTAIL.n219 VTAIL.n180 12.8005
R135 VTAIL.n40 VTAIL.n8 12.8005
R136 VTAIL.n45 VTAIL.n6 12.8005
R137 VTAIL.n161 VTAIL.n122 12.8005
R138 VTAIL.n156 VTAIL.n124 12.8005
R139 VTAIL.n103 VTAIL.n64 12.8005
R140 VTAIL.n98 VTAIL.n66 12.8005
R141 VTAIL.n211 VTAIL.n210 12.0247
R142 VTAIL.n220 VTAIL.n178 12.0247
R143 VTAIL.n37 VTAIL.n36 12.0247
R144 VTAIL.n46 VTAIL.n4 12.0247
R145 VTAIL.n162 VTAIL.n120 12.0247
R146 VTAIL.n153 VTAIL.n152 12.0247
R147 VTAIL.n104 VTAIL.n62 12.0247
R148 VTAIL.n95 VTAIL.n94 12.0247
R149 VTAIL.n206 VTAIL.n184 11.249
R150 VTAIL.n224 VTAIL.n223 11.249
R151 VTAIL.n32 VTAIL.n10 11.249
R152 VTAIL.n50 VTAIL.n49 11.249
R153 VTAIL.n166 VTAIL.n165 11.249
R154 VTAIL.n149 VTAIL.n126 11.249
R155 VTAIL.n108 VTAIL.n107 11.249
R156 VTAIL.n91 VTAIL.n68 11.249
R157 VTAIL.n205 VTAIL.n186 10.4732
R158 VTAIL.n227 VTAIL.n176 10.4732
R159 VTAIL.n31 VTAIL.n12 10.4732
R160 VTAIL.n53 VTAIL.n2 10.4732
R161 VTAIL.n169 VTAIL.n118 10.4732
R162 VTAIL.n148 VTAIL.n129 10.4732
R163 VTAIL.n111 VTAIL.n60 10.4732
R164 VTAIL.n90 VTAIL.n71 10.4732
R165 VTAIL.n193 VTAIL.n191 10.2747
R166 VTAIL.n19 VTAIL.n17 10.2747
R167 VTAIL.n136 VTAIL.n134 10.2747
R168 VTAIL.n78 VTAIL.n76 10.2747
R169 VTAIL.n202 VTAIL.n201 9.69747
R170 VTAIL.n228 VTAIL.n174 9.69747
R171 VTAIL.n28 VTAIL.n27 9.69747
R172 VTAIL.n54 VTAIL.n0 9.69747
R173 VTAIL.n170 VTAIL.n116 9.69747
R174 VTAIL.n145 VTAIL.n144 9.69747
R175 VTAIL.n112 VTAIL.n58 9.69747
R176 VTAIL.n87 VTAIL.n86 9.69747
R177 VTAIL.n230 VTAIL.n229 9.45567
R178 VTAIL.n56 VTAIL.n55 9.45567
R179 VTAIL.n172 VTAIL.n171 9.45567
R180 VTAIL.n114 VTAIL.n113 9.45567
R181 VTAIL.n229 VTAIL.n228 9.3005
R182 VTAIL.n176 VTAIL.n175 9.3005
R183 VTAIL.n223 VTAIL.n222 9.3005
R184 VTAIL.n221 VTAIL.n220 9.3005
R185 VTAIL.n180 VTAIL.n179 9.3005
R186 VTAIL.n195 VTAIL.n194 9.3005
R187 VTAIL.n197 VTAIL.n196 9.3005
R188 VTAIL.n188 VTAIL.n187 9.3005
R189 VTAIL.n203 VTAIL.n202 9.3005
R190 VTAIL.n205 VTAIL.n204 9.3005
R191 VTAIL.n184 VTAIL.n183 9.3005
R192 VTAIL.n212 VTAIL.n211 9.3005
R193 VTAIL.n214 VTAIL.n213 9.3005
R194 VTAIL.n55 VTAIL.n54 9.3005
R195 VTAIL.n2 VTAIL.n1 9.3005
R196 VTAIL.n49 VTAIL.n48 9.3005
R197 VTAIL.n47 VTAIL.n46 9.3005
R198 VTAIL.n6 VTAIL.n5 9.3005
R199 VTAIL.n21 VTAIL.n20 9.3005
R200 VTAIL.n23 VTAIL.n22 9.3005
R201 VTAIL.n14 VTAIL.n13 9.3005
R202 VTAIL.n29 VTAIL.n28 9.3005
R203 VTAIL.n31 VTAIL.n30 9.3005
R204 VTAIL.n10 VTAIL.n9 9.3005
R205 VTAIL.n38 VTAIL.n37 9.3005
R206 VTAIL.n40 VTAIL.n39 9.3005
R207 VTAIL.n138 VTAIL.n137 9.3005
R208 VTAIL.n140 VTAIL.n139 9.3005
R209 VTAIL.n131 VTAIL.n130 9.3005
R210 VTAIL.n146 VTAIL.n145 9.3005
R211 VTAIL.n148 VTAIL.n147 9.3005
R212 VTAIL.n126 VTAIL.n125 9.3005
R213 VTAIL.n154 VTAIL.n153 9.3005
R214 VTAIL.n156 VTAIL.n155 9.3005
R215 VTAIL.n171 VTAIL.n170 9.3005
R216 VTAIL.n118 VTAIL.n117 9.3005
R217 VTAIL.n165 VTAIL.n164 9.3005
R218 VTAIL.n163 VTAIL.n162 9.3005
R219 VTAIL.n122 VTAIL.n121 9.3005
R220 VTAIL.n80 VTAIL.n79 9.3005
R221 VTAIL.n82 VTAIL.n81 9.3005
R222 VTAIL.n73 VTAIL.n72 9.3005
R223 VTAIL.n88 VTAIL.n87 9.3005
R224 VTAIL.n90 VTAIL.n89 9.3005
R225 VTAIL.n68 VTAIL.n67 9.3005
R226 VTAIL.n96 VTAIL.n95 9.3005
R227 VTAIL.n98 VTAIL.n97 9.3005
R228 VTAIL.n113 VTAIL.n112 9.3005
R229 VTAIL.n60 VTAIL.n59 9.3005
R230 VTAIL.n107 VTAIL.n106 9.3005
R231 VTAIL.n105 VTAIL.n104 9.3005
R232 VTAIL.n64 VTAIL.n63 9.3005
R233 VTAIL.n198 VTAIL.n188 8.92171
R234 VTAIL.n24 VTAIL.n14 8.92171
R235 VTAIL.n141 VTAIL.n131 8.92171
R236 VTAIL.n83 VTAIL.n73 8.92171
R237 VTAIL.n197 VTAIL.n190 8.14595
R238 VTAIL.n23 VTAIL.n16 8.14595
R239 VTAIL.n140 VTAIL.n133 8.14595
R240 VTAIL.n82 VTAIL.n75 8.14595
R241 VTAIL.n194 VTAIL.n193 7.3702
R242 VTAIL.n20 VTAIL.n19 7.3702
R243 VTAIL.n137 VTAIL.n136 7.3702
R244 VTAIL.n79 VTAIL.n78 7.3702
R245 VTAIL.n194 VTAIL.n190 5.81868
R246 VTAIL.n20 VTAIL.n16 5.81868
R247 VTAIL.n137 VTAIL.n133 5.81868
R248 VTAIL.n79 VTAIL.n75 5.81868
R249 VTAIL.n198 VTAIL.n197 5.04292
R250 VTAIL.n24 VTAIL.n23 5.04292
R251 VTAIL.n141 VTAIL.n140 5.04292
R252 VTAIL.n83 VTAIL.n82 5.04292
R253 VTAIL.n201 VTAIL.n188 4.26717
R254 VTAIL.n230 VTAIL.n174 4.26717
R255 VTAIL.n27 VTAIL.n14 4.26717
R256 VTAIL.n56 VTAIL.n0 4.26717
R257 VTAIL.n172 VTAIL.n116 4.26717
R258 VTAIL.n144 VTAIL.n131 4.26717
R259 VTAIL.n114 VTAIL.n58 4.26717
R260 VTAIL.n86 VTAIL.n73 4.26717
R261 VTAIL.n202 VTAIL.n186 3.49141
R262 VTAIL.n228 VTAIL.n227 3.49141
R263 VTAIL.n28 VTAIL.n12 3.49141
R264 VTAIL.n54 VTAIL.n53 3.49141
R265 VTAIL.n170 VTAIL.n169 3.49141
R266 VTAIL.n145 VTAIL.n129 3.49141
R267 VTAIL.n112 VTAIL.n111 3.49141
R268 VTAIL.n87 VTAIL.n71 3.49141
R269 VTAIL.n195 VTAIL.n191 2.84303
R270 VTAIL.n21 VTAIL.n17 2.84303
R271 VTAIL.n138 VTAIL.n134 2.84303
R272 VTAIL.n80 VTAIL.n76 2.84303
R273 VTAIL.n206 VTAIL.n205 2.71565
R274 VTAIL.n224 VTAIL.n176 2.71565
R275 VTAIL.n32 VTAIL.n31 2.71565
R276 VTAIL.n50 VTAIL.n2 2.71565
R277 VTAIL.n166 VTAIL.n118 2.71565
R278 VTAIL.n149 VTAIL.n148 2.71565
R279 VTAIL.n108 VTAIL.n60 2.71565
R280 VTAIL.n91 VTAIL.n90 2.71565
R281 VTAIL.n173 VTAIL.n115 1.97464
R282 VTAIL.n210 VTAIL.n184 1.93989
R283 VTAIL.n223 VTAIL.n178 1.93989
R284 VTAIL.n36 VTAIL.n10 1.93989
R285 VTAIL.n49 VTAIL.n4 1.93989
R286 VTAIL.n165 VTAIL.n120 1.93989
R287 VTAIL.n152 VTAIL.n126 1.93989
R288 VTAIL.n107 VTAIL.n62 1.93989
R289 VTAIL.n94 VTAIL.n68 1.93989
R290 VTAIL VTAIL.n57 1.28067
R291 VTAIL.n211 VTAIL.n182 1.16414
R292 VTAIL.n220 VTAIL.n219 1.16414
R293 VTAIL.n37 VTAIL.n8 1.16414
R294 VTAIL.n46 VTAIL.n45 1.16414
R295 VTAIL.n162 VTAIL.n161 1.16414
R296 VTAIL.n153 VTAIL.n124 1.16414
R297 VTAIL.n104 VTAIL.n103 1.16414
R298 VTAIL.n95 VTAIL.n66 1.16414
R299 VTAIL VTAIL.n231 0.694465
R300 VTAIL.n215 VTAIL.n214 0.388379
R301 VTAIL.n216 VTAIL.n180 0.388379
R302 VTAIL.n41 VTAIL.n40 0.388379
R303 VTAIL.n42 VTAIL.n6 0.388379
R304 VTAIL.n158 VTAIL.n122 0.388379
R305 VTAIL.n157 VTAIL.n156 0.388379
R306 VTAIL.n100 VTAIL.n64 0.388379
R307 VTAIL.n99 VTAIL.n98 0.388379
R308 VTAIL.n196 VTAIL.n195 0.155672
R309 VTAIL.n196 VTAIL.n187 0.155672
R310 VTAIL.n203 VTAIL.n187 0.155672
R311 VTAIL.n204 VTAIL.n203 0.155672
R312 VTAIL.n204 VTAIL.n183 0.155672
R313 VTAIL.n212 VTAIL.n183 0.155672
R314 VTAIL.n213 VTAIL.n212 0.155672
R315 VTAIL.n213 VTAIL.n179 0.155672
R316 VTAIL.n221 VTAIL.n179 0.155672
R317 VTAIL.n222 VTAIL.n221 0.155672
R318 VTAIL.n222 VTAIL.n175 0.155672
R319 VTAIL.n229 VTAIL.n175 0.155672
R320 VTAIL.n22 VTAIL.n21 0.155672
R321 VTAIL.n22 VTAIL.n13 0.155672
R322 VTAIL.n29 VTAIL.n13 0.155672
R323 VTAIL.n30 VTAIL.n29 0.155672
R324 VTAIL.n30 VTAIL.n9 0.155672
R325 VTAIL.n38 VTAIL.n9 0.155672
R326 VTAIL.n39 VTAIL.n38 0.155672
R327 VTAIL.n39 VTAIL.n5 0.155672
R328 VTAIL.n47 VTAIL.n5 0.155672
R329 VTAIL.n48 VTAIL.n47 0.155672
R330 VTAIL.n48 VTAIL.n1 0.155672
R331 VTAIL.n55 VTAIL.n1 0.155672
R332 VTAIL.n171 VTAIL.n117 0.155672
R333 VTAIL.n164 VTAIL.n117 0.155672
R334 VTAIL.n164 VTAIL.n163 0.155672
R335 VTAIL.n163 VTAIL.n121 0.155672
R336 VTAIL.n155 VTAIL.n121 0.155672
R337 VTAIL.n155 VTAIL.n154 0.155672
R338 VTAIL.n154 VTAIL.n125 0.155672
R339 VTAIL.n147 VTAIL.n125 0.155672
R340 VTAIL.n147 VTAIL.n146 0.155672
R341 VTAIL.n146 VTAIL.n130 0.155672
R342 VTAIL.n139 VTAIL.n130 0.155672
R343 VTAIL.n139 VTAIL.n138 0.155672
R344 VTAIL.n113 VTAIL.n59 0.155672
R345 VTAIL.n106 VTAIL.n59 0.155672
R346 VTAIL.n106 VTAIL.n105 0.155672
R347 VTAIL.n105 VTAIL.n63 0.155672
R348 VTAIL.n97 VTAIL.n63 0.155672
R349 VTAIL.n97 VTAIL.n96 0.155672
R350 VTAIL.n96 VTAIL.n67 0.155672
R351 VTAIL.n89 VTAIL.n67 0.155672
R352 VTAIL.n89 VTAIL.n88 0.155672
R353 VTAIL.n88 VTAIL.n72 0.155672
R354 VTAIL.n81 VTAIL.n72 0.155672
R355 VTAIL.n81 VTAIL.n80 0.155672
R356 VDD1.n52 VDD1.n0 289.615
R357 VDD1.n109 VDD1.n57 289.615
R358 VDD1.n53 VDD1.n52 185
R359 VDD1.n51 VDD1.n50 185
R360 VDD1.n4 VDD1.n3 185
R361 VDD1.n45 VDD1.n44 185
R362 VDD1.n43 VDD1.n42 185
R363 VDD1.n41 VDD1.n7 185
R364 VDD1.n11 VDD1.n8 185
R365 VDD1.n36 VDD1.n35 185
R366 VDD1.n34 VDD1.n33 185
R367 VDD1.n13 VDD1.n12 185
R368 VDD1.n28 VDD1.n27 185
R369 VDD1.n26 VDD1.n25 185
R370 VDD1.n17 VDD1.n16 185
R371 VDD1.n20 VDD1.n19 185
R372 VDD1.n76 VDD1.n75 185
R373 VDD1.n73 VDD1.n72 185
R374 VDD1.n82 VDD1.n81 185
R375 VDD1.n84 VDD1.n83 185
R376 VDD1.n69 VDD1.n68 185
R377 VDD1.n90 VDD1.n89 185
R378 VDD1.n93 VDD1.n92 185
R379 VDD1.n91 VDD1.n65 185
R380 VDD1.n98 VDD1.n64 185
R381 VDD1.n100 VDD1.n99 185
R382 VDD1.n102 VDD1.n101 185
R383 VDD1.n61 VDD1.n60 185
R384 VDD1.n108 VDD1.n107 185
R385 VDD1.n110 VDD1.n109 185
R386 VDD1.t1 VDD1.n18 149.524
R387 VDD1.t0 VDD1.n74 149.524
R388 VDD1.n52 VDD1.n51 104.615
R389 VDD1.n51 VDD1.n3 104.615
R390 VDD1.n44 VDD1.n3 104.615
R391 VDD1.n44 VDD1.n43 104.615
R392 VDD1.n43 VDD1.n7 104.615
R393 VDD1.n11 VDD1.n7 104.615
R394 VDD1.n35 VDD1.n11 104.615
R395 VDD1.n35 VDD1.n34 104.615
R396 VDD1.n34 VDD1.n12 104.615
R397 VDD1.n27 VDD1.n12 104.615
R398 VDD1.n27 VDD1.n26 104.615
R399 VDD1.n26 VDD1.n16 104.615
R400 VDD1.n19 VDD1.n16 104.615
R401 VDD1.n75 VDD1.n72 104.615
R402 VDD1.n82 VDD1.n72 104.615
R403 VDD1.n83 VDD1.n82 104.615
R404 VDD1.n83 VDD1.n68 104.615
R405 VDD1.n90 VDD1.n68 104.615
R406 VDD1.n92 VDD1.n90 104.615
R407 VDD1.n92 VDD1.n91 104.615
R408 VDD1.n91 VDD1.n64 104.615
R409 VDD1.n100 VDD1.n64 104.615
R410 VDD1.n101 VDD1.n100 104.615
R411 VDD1.n101 VDD1.n60 104.615
R412 VDD1.n108 VDD1.n60 104.615
R413 VDD1.n109 VDD1.n108 104.615
R414 VDD1 VDD1.n113 88.2145
R415 VDD1.n19 VDD1.t1 52.3082
R416 VDD1.n75 VDD1.t0 52.3082
R417 VDD1 VDD1.n56 48.8987
R418 VDD1.n42 VDD1.n41 13.1884
R419 VDD1.n99 VDD1.n98 13.1884
R420 VDD1.n45 VDD1.n6 12.8005
R421 VDD1.n40 VDD1.n8 12.8005
R422 VDD1.n97 VDD1.n65 12.8005
R423 VDD1.n102 VDD1.n63 12.8005
R424 VDD1.n46 VDD1.n4 12.0247
R425 VDD1.n37 VDD1.n36 12.0247
R426 VDD1.n94 VDD1.n93 12.0247
R427 VDD1.n103 VDD1.n61 12.0247
R428 VDD1.n50 VDD1.n49 11.249
R429 VDD1.n33 VDD1.n10 11.249
R430 VDD1.n89 VDD1.n67 11.249
R431 VDD1.n107 VDD1.n106 11.249
R432 VDD1.n53 VDD1.n2 10.4732
R433 VDD1.n32 VDD1.n13 10.4732
R434 VDD1.n88 VDD1.n69 10.4732
R435 VDD1.n110 VDD1.n59 10.4732
R436 VDD1.n20 VDD1.n18 10.2747
R437 VDD1.n76 VDD1.n74 10.2747
R438 VDD1.n54 VDD1.n0 9.69747
R439 VDD1.n29 VDD1.n28 9.69747
R440 VDD1.n85 VDD1.n84 9.69747
R441 VDD1.n111 VDD1.n57 9.69747
R442 VDD1.n56 VDD1.n55 9.45567
R443 VDD1.n113 VDD1.n112 9.45567
R444 VDD1.n22 VDD1.n21 9.3005
R445 VDD1.n24 VDD1.n23 9.3005
R446 VDD1.n15 VDD1.n14 9.3005
R447 VDD1.n30 VDD1.n29 9.3005
R448 VDD1.n32 VDD1.n31 9.3005
R449 VDD1.n10 VDD1.n9 9.3005
R450 VDD1.n38 VDD1.n37 9.3005
R451 VDD1.n40 VDD1.n39 9.3005
R452 VDD1.n55 VDD1.n54 9.3005
R453 VDD1.n2 VDD1.n1 9.3005
R454 VDD1.n49 VDD1.n48 9.3005
R455 VDD1.n47 VDD1.n46 9.3005
R456 VDD1.n6 VDD1.n5 9.3005
R457 VDD1.n112 VDD1.n111 9.3005
R458 VDD1.n59 VDD1.n58 9.3005
R459 VDD1.n106 VDD1.n105 9.3005
R460 VDD1.n104 VDD1.n103 9.3005
R461 VDD1.n63 VDD1.n62 9.3005
R462 VDD1.n78 VDD1.n77 9.3005
R463 VDD1.n80 VDD1.n79 9.3005
R464 VDD1.n71 VDD1.n70 9.3005
R465 VDD1.n86 VDD1.n85 9.3005
R466 VDD1.n88 VDD1.n87 9.3005
R467 VDD1.n67 VDD1.n66 9.3005
R468 VDD1.n95 VDD1.n94 9.3005
R469 VDD1.n97 VDD1.n96 9.3005
R470 VDD1.n25 VDD1.n15 8.92171
R471 VDD1.n81 VDD1.n71 8.92171
R472 VDD1.n24 VDD1.n17 8.14595
R473 VDD1.n80 VDD1.n73 8.14595
R474 VDD1.n21 VDD1.n20 7.3702
R475 VDD1.n77 VDD1.n76 7.3702
R476 VDD1.n21 VDD1.n17 5.81868
R477 VDD1.n77 VDD1.n73 5.81868
R478 VDD1.n25 VDD1.n24 5.04292
R479 VDD1.n81 VDD1.n80 5.04292
R480 VDD1.n56 VDD1.n0 4.26717
R481 VDD1.n28 VDD1.n15 4.26717
R482 VDD1.n84 VDD1.n71 4.26717
R483 VDD1.n113 VDD1.n57 4.26717
R484 VDD1.n54 VDD1.n53 3.49141
R485 VDD1.n29 VDD1.n13 3.49141
R486 VDD1.n85 VDD1.n69 3.49141
R487 VDD1.n111 VDD1.n110 3.49141
R488 VDD1.n22 VDD1.n18 2.84303
R489 VDD1.n78 VDD1.n74 2.84303
R490 VDD1.n50 VDD1.n2 2.71565
R491 VDD1.n33 VDD1.n32 2.71565
R492 VDD1.n89 VDD1.n88 2.71565
R493 VDD1.n107 VDD1.n59 2.71565
R494 VDD1.n49 VDD1.n4 1.93989
R495 VDD1.n36 VDD1.n10 1.93989
R496 VDD1.n93 VDD1.n67 1.93989
R497 VDD1.n106 VDD1.n61 1.93989
R498 VDD1.n46 VDD1.n45 1.16414
R499 VDD1.n37 VDD1.n8 1.16414
R500 VDD1.n94 VDD1.n65 1.16414
R501 VDD1.n103 VDD1.n102 1.16414
R502 VDD1.n42 VDD1.n6 0.388379
R503 VDD1.n41 VDD1.n40 0.388379
R504 VDD1.n98 VDD1.n97 0.388379
R505 VDD1.n99 VDD1.n63 0.388379
R506 VDD1.n55 VDD1.n1 0.155672
R507 VDD1.n48 VDD1.n1 0.155672
R508 VDD1.n48 VDD1.n47 0.155672
R509 VDD1.n47 VDD1.n5 0.155672
R510 VDD1.n39 VDD1.n5 0.155672
R511 VDD1.n39 VDD1.n38 0.155672
R512 VDD1.n38 VDD1.n9 0.155672
R513 VDD1.n31 VDD1.n9 0.155672
R514 VDD1.n31 VDD1.n30 0.155672
R515 VDD1.n30 VDD1.n14 0.155672
R516 VDD1.n23 VDD1.n14 0.155672
R517 VDD1.n23 VDD1.n22 0.155672
R518 VDD1.n79 VDD1.n78 0.155672
R519 VDD1.n79 VDD1.n70 0.155672
R520 VDD1.n86 VDD1.n70 0.155672
R521 VDD1.n87 VDD1.n86 0.155672
R522 VDD1.n87 VDD1.n66 0.155672
R523 VDD1.n95 VDD1.n66 0.155672
R524 VDD1.n96 VDD1.n95 0.155672
R525 VDD1.n96 VDD1.n62 0.155672
R526 VDD1.n104 VDD1.n62 0.155672
R527 VDD1.n105 VDD1.n104 0.155672
R528 VDD1.n105 VDD1.n58 0.155672
R529 VDD1.n112 VDD1.n58 0.155672
R530 B.n665 B.n664 585
R531 B.n666 B.n665 585
R532 B.n269 B.n98 585
R533 B.n268 B.n267 585
R534 B.n266 B.n265 585
R535 B.n264 B.n263 585
R536 B.n262 B.n261 585
R537 B.n260 B.n259 585
R538 B.n258 B.n257 585
R539 B.n256 B.n255 585
R540 B.n254 B.n253 585
R541 B.n252 B.n251 585
R542 B.n250 B.n249 585
R543 B.n248 B.n247 585
R544 B.n246 B.n245 585
R545 B.n244 B.n243 585
R546 B.n242 B.n241 585
R547 B.n240 B.n239 585
R548 B.n238 B.n237 585
R549 B.n236 B.n235 585
R550 B.n234 B.n233 585
R551 B.n232 B.n231 585
R552 B.n230 B.n229 585
R553 B.n228 B.n227 585
R554 B.n226 B.n225 585
R555 B.n224 B.n223 585
R556 B.n222 B.n221 585
R557 B.n220 B.n219 585
R558 B.n218 B.n217 585
R559 B.n216 B.n215 585
R560 B.n214 B.n213 585
R561 B.n212 B.n211 585
R562 B.n210 B.n209 585
R563 B.n208 B.n207 585
R564 B.n206 B.n205 585
R565 B.n204 B.n203 585
R566 B.n202 B.n201 585
R567 B.n200 B.n199 585
R568 B.n198 B.n197 585
R569 B.n195 B.n194 585
R570 B.n193 B.n192 585
R571 B.n191 B.n190 585
R572 B.n189 B.n188 585
R573 B.n187 B.n186 585
R574 B.n185 B.n184 585
R575 B.n183 B.n182 585
R576 B.n181 B.n180 585
R577 B.n179 B.n178 585
R578 B.n177 B.n176 585
R579 B.n175 B.n174 585
R580 B.n173 B.n172 585
R581 B.n171 B.n170 585
R582 B.n169 B.n168 585
R583 B.n167 B.n166 585
R584 B.n165 B.n164 585
R585 B.n163 B.n162 585
R586 B.n161 B.n160 585
R587 B.n159 B.n158 585
R588 B.n157 B.n156 585
R589 B.n155 B.n154 585
R590 B.n153 B.n152 585
R591 B.n151 B.n150 585
R592 B.n149 B.n148 585
R593 B.n147 B.n146 585
R594 B.n145 B.n144 585
R595 B.n143 B.n142 585
R596 B.n141 B.n140 585
R597 B.n139 B.n138 585
R598 B.n137 B.n136 585
R599 B.n135 B.n134 585
R600 B.n133 B.n132 585
R601 B.n131 B.n130 585
R602 B.n129 B.n128 585
R603 B.n127 B.n126 585
R604 B.n125 B.n124 585
R605 B.n123 B.n122 585
R606 B.n121 B.n120 585
R607 B.n119 B.n118 585
R608 B.n117 B.n116 585
R609 B.n115 B.n114 585
R610 B.n113 B.n112 585
R611 B.n111 B.n110 585
R612 B.n109 B.n108 585
R613 B.n107 B.n106 585
R614 B.n105 B.n104 585
R615 B.n54 B.n53 585
R616 B.n663 B.n55 585
R617 B.n667 B.n55 585
R618 B.n662 B.n661 585
R619 B.n661 B.n51 585
R620 B.n660 B.n50 585
R621 B.n673 B.n50 585
R622 B.n659 B.n49 585
R623 B.n674 B.n49 585
R624 B.n658 B.n48 585
R625 B.n675 B.n48 585
R626 B.n657 B.n656 585
R627 B.n656 B.n44 585
R628 B.n655 B.n43 585
R629 B.n681 B.n43 585
R630 B.n654 B.n42 585
R631 B.n682 B.n42 585
R632 B.n653 B.n41 585
R633 B.n683 B.n41 585
R634 B.n652 B.n651 585
R635 B.n651 B.n37 585
R636 B.n650 B.n36 585
R637 B.n689 B.n36 585
R638 B.n649 B.n35 585
R639 B.n690 B.n35 585
R640 B.n648 B.n34 585
R641 B.n691 B.n34 585
R642 B.n647 B.n646 585
R643 B.n646 B.n30 585
R644 B.n645 B.n29 585
R645 B.n697 B.n29 585
R646 B.n644 B.n28 585
R647 B.n698 B.n28 585
R648 B.n643 B.n27 585
R649 B.n699 B.n27 585
R650 B.n642 B.n641 585
R651 B.n641 B.n23 585
R652 B.n640 B.n22 585
R653 B.n705 B.n22 585
R654 B.n639 B.n21 585
R655 B.n706 B.n21 585
R656 B.n638 B.n20 585
R657 B.n707 B.n20 585
R658 B.n637 B.n636 585
R659 B.n636 B.n19 585
R660 B.n635 B.n15 585
R661 B.n713 B.n15 585
R662 B.n634 B.n14 585
R663 B.n714 B.n14 585
R664 B.n633 B.n13 585
R665 B.n715 B.n13 585
R666 B.n632 B.n631 585
R667 B.n631 B.n12 585
R668 B.n630 B.n629 585
R669 B.n630 B.n8 585
R670 B.n628 B.n7 585
R671 B.n722 B.n7 585
R672 B.n627 B.n6 585
R673 B.n723 B.n6 585
R674 B.n626 B.n5 585
R675 B.n724 B.n5 585
R676 B.n625 B.n624 585
R677 B.n624 B.n4 585
R678 B.n623 B.n270 585
R679 B.n623 B.n622 585
R680 B.n613 B.n271 585
R681 B.n272 B.n271 585
R682 B.n615 B.n614 585
R683 B.n616 B.n615 585
R684 B.n612 B.n277 585
R685 B.n277 B.n276 585
R686 B.n611 B.n610 585
R687 B.n610 B.n609 585
R688 B.n279 B.n278 585
R689 B.n602 B.n279 585
R690 B.n601 B.n600 585
R691 B.n603 B.n601 585
R692 B.n599 B.n284 585
R693 B.n284 B.n283 585
R694 B.n598 B.n597 585
R695 B.n597 B.n596 585
R696 B.n286 B.n285 585
R697 B.n287 B.n286 585
R698 B.n589 B.n588 585
R699 B.n590 B.n589 585
R700 B.n587 B.n292 585
R701 B.n292 B.n291 585
R702 B.n586 B.n585 585
R703 B.n585 B.n584 585
R704 B.n294 B.n293 585
R705 B.n295 B.n294 585
R706 B.n577 B.n576 585
R707 B.n578 B.n577 585
R708 B.n575 B.n300 585
R709 B.n300 B.n299 585
R710 B.n574 B.n573 585
R711 B.n573 B.n572 585
R712 B.n302 B.n301 585
R713 B.n303 B.n302 585
R714 B.n565 B.n564 585
R715 B.n566 B.n565 585
R716 B.n563 B.n308 585
R717 B.n308 B.n307 585
R718 B.n562 B.n561 585
R719 B.n561 B.n560 585
R720 B.n310 B.n309 585
R721 B.n311 B.n310 585
R722 B.n553 B.n552 585
R723 B.n554 B.n553 585
R724 B.n551 B.n316 585
R725 B.n316 B.n315 585
R726 B.n550 B.n549 585
R727 B.n549 B.n548 585
R728 B.n318 B.n317 585
R729 B.n319 B.n318 585
R730 B.n541 B.n540 585
R731 B.n542 B.n541 585
R732 B.n322 B.n321 585
R733 B.n371 B.n369 585
R734 B.n372 B.n368 585
R735 B.n372 B.n323 585
R736 B.n375 B.n374 585
R737 B.n376 B.n367 585
R738 B.n378 B.n377 585
R739 B.n380 B.n366 585
R740 B.n383 B.n382 585
R741 B.n384 B.n365 585
R742 B.n386 B.n385 585
R743 B.n388 B.n364 585
R744 B.n391 B.n390 585
R745 B.n392 B.n363 585
R746 B.n394 B.n393 585
R747 B.n396 B.n362 585
R748 B.n399 B.n398 585
R749 B.n400 B.n361 585
R750 B.n402 B.n401 585
R751 B.n404 B.n360 585
R752 B.n407 B.n406 585
R753 B.n408 B.n359 585
R754 B.n410 B.n409 585
R755 B.n412 B.n358 585
R756 B.n415 B.n414 585
R757 B.n416 B.n357 585
R758 B.n418 B.n417 585
R759 B.n420 B.n356 585
R760 B.n423 B.n422 585
R761 B.n424 B.n355 585
R762 B.n426 B.n425 585
R763 B.n428 B.n354 585
R764 B.n431 B.n430 585
R765 B.n432 B.n353 585
R766 B.n434 B.n433 585
R767 B.n436 B.n352 585
R768 B.n439 B.n438 585
R769 B.n440 B.n351 585
R770 B.n445 B.n444 585
R771 B.n447 B.n350 585
R772 B.n450 B.n449 585
R773 B.n451 B.n349 585
R774 B.n453 B.n452 585
R775 B.n455 B.n348 585
R776 B.n458 B.n457 585
R777 B.n459 B.n347 585
R778 B.n461 B.n460 585
R779 B.n463 B.n346 585
R780 B.n466 B.n465 585
R781 B.n467 B.n342 585
R782 B.n469 B.n468 585
R783 B.n471 B.n341 585
R784 B.n474 B.n473 585
R785 B.n475 B.n340 585
R786 B.n477 B.n476 585
R787 B.n479 B.n339 585
R788 B.n482 B.n481 585
R789 B.n483 B.n338 585
R790 B.n485 B.n484 585
R791 B.n487 B.n337 585
R792 B.n490 B.n489 585
R793 B.n491 B.n336 585
R794 B.n493 B.n492 585
R795 B.n495 B.n335 585
R796 B.n498 B.n497 585
R797 B.n499 B.n334 585
R798 B.n501 B.n500 585
R799 B.n503 B.n333 585
R800 B.n506 B.n505 585
R801 B.n507 B.n332 585
R802 B.n509 B.n508 585
R803 B.n511 B.n331 585
R804 B.n514 B.n513 585
R805 B.n515 B.n330 585
R806 B.n517 B.n516 585
R807 B.n519 B.n329 585
R808 B.n522 B.n521 585
R809 B.n523 B.n328 585
R810 B.n525 B.n524 585
R811 B.n527 B.n327 585
R812 B.n530 B.n529 585
R813 B.n531 B.n326 585
R814 B.n533 B.n532 585
R815 B.n535 B.n325 585
R816 B.n538 B.n537 585
R817 B.n539 B.n324 585
R818 B.n544 B.n543 585
R819 B.n543 B.n542 585
R820 B.n545 B.n320 585
R821 B.n320 B.n319 585
R822 B.n547 B.n546 585
R823 B.n548 B.n547 585
R824 B.n314 B.n313 585
R825 B.n315 B.n314 585
R826 B.n556 B.n555 585
R827 B.n555 B.n554 585
R828 B.n557 B.n312 585
R829 B.n312 B.n311 585
R830 B.n559 B.n558 585
R831 B.n560 B.n559 585
R832 B.n306 B.n305 585
R833 B.n307 B.n306 585
R834 B.n568 B.n567 585
R835 B.n567 B.n566 585
R836 B.n569 B.n304 585
R837 B.n304 B.n303 585
R838 B.n571 B.n570 585
R839 B.n572 B.n571 585
R840 B.n298 B.n297 585
R841 B.n299 B.n298 585
R842 B.n580 B.n579 585
R843 B.n579 B.n578 585
R844 B.n581 B.n296 585
R845 B.n296 B.n295 585
R846 B.n583 B.n582 585
R847 B.n584 B.n583 585
R848 B.n290 B.n289 585
R849 B.n291 B.n290 585
R850 B.n592 B.n591 585
R851 B.n591 B.n590 585
R852 B.n593 B.n288 585
R853 B.n288 B.n287 585
R854 B.n595 B.n594 585
R855 B.n596 B.n595 585
R856 B.n282 B.n281 585
R857 B.n283 B.n282 585
R858 B.n605 B.n604 585
R859 B.n604 B.n603 585
R860 B.n606 B.n280 585
R861 B.n602 B.n280 585
R862 B.n608 B.n607 585
R863 B.n609 B.n608 585
R864 B.n275 B.n274 585
R865 B.n276 B.n275 585
R866 B.n618 B.n617 585
R867 B.n617 B.n616 585
R868 B.n619 B.n273 585
R869 B.n273 B.n272 585
R870 B.n621 B.n620 585
R871 B.n622 B.n621 585
R872 B.n3 B.n0 585
R873 B.n4 B.n3 585
R874 B.n721 B.n1 585
R875 B.n722 B.n721 585
R876 B.n720 B.n719 585
R877 B.n720 B.n8 585
R878 B.n718 B.n9 585
R879 B.n12 B.n9 585
R880 B.n717 B.n716 585
R881 B.n716 B.n715 585
R882 B.n11 B.n10 585
R883 B.n714 B.n11 585
R884 B.n712 B.n711 585
R885 B.n713 B.n712 585
R886 B.n710 B.n16 585
R887 B.n19 B.n16 585
R888 B.n709 B.n708 585
R889 B.n708 B.n707 585
R890 B.n18 B.n17 585
R891 B.n706 B.n18 585
R892 B.n704 B.n703 585
R893 B.n705 B.n704 585
R894 B.n702 B.n24 585
R895 B.n24 B.n23 585
R896 B.n701 B.n700 585
R897 B.n700 B.n699 585
R898 B.n26 B.n25 585
R899 B.n698 B.n26 585
R900 B.n696 B.n695 585
R901 B.n697 B.n696 585
R902 B.n694 B.n31 585
R903 B.n31 B.n30 585
R904 B.n693 B.n692 585
R905 B.n692 B.n691 585
R906 B.n33 B.n32 585
R907 B.n690 B.n33 585
R908 B.n688 B.n687 585
R909 B.n689 B.n688 585
R910 B.n686 B.n38 585
R911 B.n38 B.n37 585
R912 B.n685 B.n684 585
R913 B.n684 B.n683 585
R914 B.n40 B.n39 585
R915 B.n682 B.n40 585
R916 B.n680 B.n679 585
R917 B.n681 B.n680 585
R918 B.n678 B.n45 585
R919 B.n45 B.n44 585
R920 B.n677 B.n676 585
R921 B.n676 B.n675 585
R922 B.n47 B.n46 585
R923 B.n674 B.n47 585
R924 B.n672 B.n671 585
R925 B.n673 B.n672 585
R926 B.n670 B.n52 585
R927 B.n52 B.n51 585
R928 B.n669 B.n668 585
R929 B.n668 B.n667 585
R930 B.n725 B.n724 585
R931 B.n723 B.n2 585
R932 B.n668 B.n54 506.916
R933 B.n665 B.n55 506.916
R934 B.n541 B.n324 506.916
R935 B.n543 B.n322 506.916
R936 B.n99 B.t11 326.269
R937 B.n343 B.t5 326.269
R938 B.n101 B.t14 326.269
R939 B.n441 B.t8 326.269
R940 B.n101 B.t13 289.908
R941 B.n99 B.t9 289.908
R942 B.n343 B.t2 289.908
R943 B.n441 B.t6 289.908
R944 B.n100 B.t12 258.584
R945 B.n344 B.t4 258.584
R946 B.n102 B.t15 258.584
R947 B.n442 B.t7 258.584
R948 B.n666 B.n97 256.663
R949 B.n666 B.n96 256.663
R950 B.n666 B.n95 256.663
R951 B.n666 B.n94 256.663
R952 B.n666 B.n93 256.663
R953 B.n666 B.n92 256.663
R954 B.n666 B.n91 256.663
R955 B.n666 B.n90 256.663
R956 B.n666 B.n89 256.663
R957 B.n666 B.n88 256.663
R958 B.n666 B.n87 256.663
R959 B.n666 B.n86 256.663
R960 B.n666 B.n85 256.663
R961 B.n666 B.n84 256.663
R962 B.n666 B.n83 256.663
R963 B.n666 B.n82 256.663
R964 B.n666 B.n81 256.663
R965 B.n666 B.n80 256.663
R966 B.n666 B.n79 256.663
R967 B.n666 B.n78 256.663
R968 B.n666 B.n77 256.663
R969 B.n666 B.n76 256.663
R970 B.n666 B.n75 256.663
R971 B.n666 B.n74 256.663
R972 B.n666 B.n73 256.663
R973 B.n666 B.n72 256.663
R974 B.n666 B.n71 256.663
R975 B.n666 B.n70 256.663
R976 B.n666 B.n69 256.663
R977 B.n666 B.n68 256.663
R978 B.n666 B.n67 256.663
R979 B.n666 B.n66 256.663
R980 B.n666 B.n65 256.663
R981 B.n666 B.n64 256.663
R982 B.n666 B.n63 256.663
R983 B.n666 B.n62 256.663
R984 B.n666 B.n61 256.663
R985 B.n666 B.n60 256.663
R986 B.n666 B.n59 256.663
R987 B.n666 B.n58 256.663
R988 B.n666 B.n57 256.663
R989 B.n666 B.n56 256.663
R990 B.n370 B.n323 256.663
R991 B.n373 B.n323 256.663
R992 B.n379 B.n323 256.663
R993 B.n381 B.n323 256.663
R994 B.n387 B.n323 256.663
R995 B.n389 B.n323 256.663
R996 B.n395 B.n323 256.663
R997 B.n397 B.n323 256.663
R998 B.n403 B.n323 256.663
R999 B.n405 B.n323 256.663
R1000 B.n411 B.n323 256.663
R1001 B.n413 B.n323 256.663
R1002 B.n419 B.n323 256.663
R1003 B.n421 B.n323 256.663
R1004 B.n427 B.n323 256.663
R1005 B.n429 B.n323 256.663
R1006 B.n435 B.n323 256.663
R1007 B.n437 B.n323 256.663
R1008 B.n446 B.n323 256.663
R1009 B.n448 B.n323 256.663
R1010 B.n454 B.n323 256.663
R1011 B.n456 B.n323 256.663
R1012 B.n462 B.n323 256.663
R1013 B.n464 B.n323 256.663
R1014 B.n470 B.n323 256.663
R1015 B.n472 B.n323 256.663
R1016 B.n478 B.n323 256.663
R1017 B.n480 B.n323 256.663
R1018 B.n486 B.n323 256.663
R1019 B.n488 B.n323 256.663
R1020 B.n494 B.n323 256.663
R1021 B.n496 B.n323 256.663
R1022 B.n502 B.n323 256.663
R1023 B.n504 B.n323 256.663
R1024 B.n510 B.n323 256.663
R1025 B.n512 B.n323 256.663
R1026 B.n518 B.n323 256.663
R1027 B.n520 B.n323 256.663
R1028 B.n526 B.n323 256.663
R1029 B.n528 B.n323 256.663
R1030 B.n534 B.n323 256.663
R1031 B.n536 B.n323 256.663
R1032 B.n727 B.n726 256.663
R1033 B.n106 B.n105 163.367
R1034 B.n110 B.n109 163.367
R1035 B.n114 B.n113 163.367
R1036 B.n118 B.n117 163.367
R1037 B.n122 B.n121 163.367
R1038 B.n126 B.n125 163.367
R1039 B.n130 B.n129 163.367
R1040 B.n134 B.n133 163.367
R1041 B.n138 B.n137 163.367
R1042 B.n142 B.n141 163.367
R1043 B.n146 B.n145 163.367
R1044 B.n150 B.n149 163.367
R1045 B.n154 B.n153 163.367
R1046 B.n158 B.n157 163.367
R1047 B.n162 B.n161 163.367
R1048 B.n166 B.n165 163.367
R1049 B.n170 B.n169 163.367
R1050 B.n174 B.n173 163.367
R1051 B.n178 B.n177 163.367
R1052 B.n182 B.n181 163.367
R1053 B.n186 B.n185 163.367
R1054 B.n190 B.n189 163.367
R1055 B.n194 B.n193 163.367
R1056 B.n199 B.n198 163.367
R1057 B.n203 B.n202 163.367
R1058 B.n207 B.n206 163.367
R1059 B.n211 B.n210 163.367
R1060 B.n215 B.n214 163.367
R1061 B.n219 B.n218 163.367
R1062 B.n223 B.n222 163.367
R1063 B.n227 B.n226 163.367
R1064 B.n231 B.n230 163.367
R1065 B.n235 B.n234 163.367
R1066 B.n239 B.n238 163.367
R1067 B.n243 B.n242 163.367
R1068 B.n247 B.n246 163.367
R1069 B.n251 B.n250 163.367
R1070 B.n255 B.n254 163.367
R1071 B.n259 B.n258 163.367
R1072 B.n263 B.n262 163.367
R1073 B.n267 B.n266 163.367
R1074 B.n665 B.n98 163.367
R1075 B.n541 B.n318 163.367
R1076 B.n549 B.n318 163.367
R1077 B.n549 B.n316 163.367
R1078 B.n553 B.n316 163.367
R1079 B.n553 B.n310 163.367
R1080 B.n561 B.n310 163.367
R1081 B.n561 B.n308 163.367
R1082 B.n565 B.n308 163.367
R1083 B.n565 B.n302 163.367
R1084 B.n573 B.n302 163.367
R1085 B.n573 B.n300 163.367
R1086 B.n577 B.n300 163.367
R1087 B.n577 B.n294 163.367
R1088 B.n585 B.n294 163.367
R1089 B.n585 B.n292 163.367
R1090 B.n589 B.n292 163.367
R1091 B.n589 B.n286 163.367
R1092 B.n597 B.n286 163.367
R1093 B.n597 B.n284 163.367
R1094 B.n601 B.n284 163.367
R1095 B.n601 B.n279 163.367
R1096 B.n610 B.n279 163.367
R1097 B.n610 B.n277 163.367
R1098 B.n615 B.n277 163.367
R1099 B.n615 B.n271 163.367
R1100 B.n623 B.n271 163.367
R1101 B.n624 B.n623 163.367
R1102 B.n624 B.n5 163.367
R1103 B.n6 B.n5 163.367
R1104 B.n7 B.n6 163.367
R1105 B.n630 B.n7 163.367
R1106 B.n631 B.n630 163.367
R1107 B.n631 B.n13 163.367
R1108 B.n14 B.n13 163.367
R1109 B.n15 B.n14 163.367
R1110 B.n636 B.n15 163.367
R1111 B.n636 B.n20 163.367
R1112 B.n21 B.n20 163.367
R1113 B.n22 B.n21 163.367
R1114 B.n641 B.n22 163.367
R1115 B.n641 B.n27 163.367
R1116 B.n28 B.n27 163.367
R1117 B.n29 B.n28 163.367
R1118 B.n646 B.n29 163.367
R1119 B.n646 B.n34 163.367
R1120 B.n35 B.n34 163.367
R1121 B.n36 B.n35 163.367
R1122 B.n651 B.n36 163.367
R1123 B.n651 B.n41 163.367
R1124 B.n42 B.n41 163.367
R1125 B.n43 B.n42 163.367
R1126 B.n656 B.n43 163.367
R1127 B.n656 B.n48 163.367
R1128 B.n49 B.n48 163.367
R1129 B.n50 B.n49 163.367
R1130 B.n661 B.n50 163.367
R1131 B.n661 B.n55 163.367
R1132 B.n372 B.n371 163.367
R1133 B.n374 B.n372 163.367
R1134 B.n378 B.n367 163.367
R1135 B.n382 B.n380 163.367
R1136 B.n386 B.n365 163.367
R1137 B.n390 B.n388 163.367
R1138 B.n394 B.n363 163.367
R1139 B.n398 B.n396 163.367
R1140 B.n402 B.n361 163.367
R1141 B.n406 B.n404 163.367
R1142 B.n410 B.n359 163.367
R1143 B.n414 B.n412 163.367
R1144 B.n418 B.n357 163.367
R1145 B.n422 B.n420 163.367
R1146 B.n426 B.n355 163.367
R1147 B.n430 B.n428 163.367
R1148 B.n434 B.n353 163.367
R1149 B.n438 B.n436 163.367
R1150 B.n445 B.n351 163.367
R1151 B.n449 B.n447 163.367
R1152 B.n453 B.n349 163.367
R1153 B.n457 B.n455 163.367
R1154 B.n461 B.n347 163.367
R1155 B.n465 B.n463 163.367
R1156 B.n469 B.n342 163.367
R1157 B.n473 B.n471 163.367
R1158 B.n477 B.n340 163.367
R1159 B.n481 B.n479 163.367
R1160 B.n485 B.n338 163.367
R1161 B.n489 B.n487 163.367
R1162 B.n493 B.n336 163.367
R1163 B.n497 B.n495 163.367
R1164 B.n501 B.n334 163.367
R1165 B.n505 B.n503 163.367
R1166 B.n509 B.n332 163.367
R1167 B.n513 B.n511 163.367
R1168 B.n517 B.n330 163.367
R1169 B.n521 B.n519 163.367
R1170 B.n525 B.n328 163.367
R1171 B.n529 B.n527 163.367
R1172 B.n533 B.n326 163.367
R1173 B.n537 B.n535 163.367
R1174 B.n543 B.n320 163.367
R1175 B.n547 B.n320 163.367
R1176 B.n547 B.n314 163.367
R1177 B.n555 B.n314 163.367
R1178 B.n555 B.n312 163.367
R1179 B.n559 B.n312 163.367
R1180 B.n559 B.n306 163.367
R1181 B.n567 B.n306 163.367
R1182 B.n567 B.n304 163.367
R1183 B.n571 B.n304 163.367
R1184 B.n571 B.n298 163.367
R1185 B.n579 B.n298 163.367
R1186 B.n579 B.n296 163.367
R1187 B.n583 B.n296 163.367
R1188 B.n583 B.n290 163.367
R1189 B.n591 B.n290 163.367
R1190 B.n591 B.n288 163.367
R1191 B.n595 B.n288 163.367
R1192 B.n595 B.n282 163.367
R1193 B.n604 B.n282 163.367
R1194 B.n604 B.n280 163.367
R1195 B.n608 B.n280 163.367
R1196 B.n608 B.n275 163.367
R1197 B.n617 B.n275 163.367
R1198 B.n617 B.n273 163.367
R1199 B.n621 B.n273 163.367
R1200 B.n621 B.n3 163.367
R1201 B.n725 B.n3 163.367
R1202 B.n721 B.n2 163.367
R1203 B.n721 B.n720 163.367
R1204 B.n720 B.n9 163.367
R1205 B.n716 B.n9 163.367
R1206 B.n716 B.n11 163.367
R1207 B.n712 B.n11 163.367
R1208 B.n712 B.n16 163.367
R1209 B.n708 B.n16 163.367
R1210 B.n708 B.n18 163.367
R1211 B.n704 B.n18 163.367
R1212 B.n704 B.n24 163.367
R1213 B.n700 B.n24 163.367
R1214 B.n700 B.n26 163.367
R1215 B.n696 B.n26 163.367
R1216 B.n696 B.n31 163.367
R1217 B.n692 B.n31 163.367
R1218 B.n692 B.n33 163.367
R1219 B.n688 B.n33 163.367
R1220 B.n688 B.n38 163.367
R1221 B.n684 B.n38 163.367
R1222 B.n684 B.n40 163.367
R1223 B.n680 B.n40 163.367
R1224 B.n680 B.n45 163.367
R1225 B.n676 B.n45 163.367
R1226 B.n676 B.n47 163.367
R1227 B.n672 B.n47 163.367
R1228 B.n672 B.n52 163.367
R1229 B.n668 B.n52 163.367
R1230 B.n542 B.n323 91.9264
R1231 B.n667 B.n666 91.9264
R1232 B.n56 B.n54 71.676
R1233 B.n106 B.n57 71.676
R1234 B.n110 B.n58 71.676
R1235 B.n114 B.n59 71.676
R1236 B.n118 B.n60 71.676
R1237 B.n122 B.n61 71.676
R1238 B.n126 B.n62 71.676
R1239 B.n130 B.n63 71.676
R1240 B.n134 B.n64 71.676
R1241 B.n138 B.n65 71.676
R1242 B.n142 B.n66 71.676
R1243 B.n146 B.n67 71.676
R1244 B.n150 B.n68 71.676
R1245 B.n154 B.n69 71.676
R1246 B.n158 B.n70 71.676
R1247 B.n162 B.n71 71.676
R1248 B.n166 B.n72 71.676
R1249 B.n170 B.n73 71.676
R1250 B.n174 B.n74 71.676
R1251 B.n178 B.n75 71.676
R1252 B.n182 B.n76 71.676
R1253 B.n186 B.n77 71.676
R1254 B.n190 B.n78 71.676
R1255 B.n194 B.n79 71.676
R1256 B.n199 B.n80 71.676
R1257 B.n203 B.n81 71.676
R1258 B.n207 B.n82 71.676
R1259 B.n211 B.n83 71.676
R1260 B.n215 B.n84 71.676
R1261 B.n219 B.n85 71.676
R1262 B.n223 B.n86 71.676
R1263 B.n227 B.n87 71.676
R1264 B.n231 B.n88 71.676
R1265 B.n235 B.n89 71.676
R1266 B.n239 B.n90 71.676
R1267 B.n243 B.n91 71.676
R1268 B.n247 B.n92 71.676
R1269 B.n251 B.n93 71.676
R1270 B.n255 B.n94 71.676
R1271 B.n259 B.n95 71.676
R1272 B.n263 B.n96 71.676
R1273 B.n267 B.n97 71.676
R1274 B.n98 B.n97 71.676
R1275 B.n266 B.n96 71.676
R1276 B.n262 B.n95 71.676
R1277 B.n258 B.n94 71.676
R1278 B.n254 B.n93 71.676
R1279 B.n250 B.n92 71.676
R1280 B.n246 B.n91 71.676
R1281 B.n242 B.n90 71.676
R1282 B.n238 B.n89 71.676
R1283 B.n234 B.n88 71.676
R1284 B.n230 B.n87 71.676
R1285 B.n226 B.n86 71.676
R1286 B.n222 B.n85 71.676
R1287 B.n218 B.n84 71.676
R1288 B.n214 B.n83 71.676
R1289 B.n210 B.n82 71.676
R1290 B.n206 B.n81 71.676
R1291 B.n202 B.n80 71.676
R1292 B.n198 B.n79 71.676
R1293 B.n193 B.n78 71.676
R1294 B.n189 B.n77 71.676
R1295 B.n185 B.n76 71.676
R1296 B.n181 B.n75 71.676
R1297 B.n177 B.n74 71.676
R1298 B.n173 B.n73 71.676
R1299 B.n169 B.n72 71.676
R1300 B.n165 B.n71 71.676
R1301 B.n161 B.n70 71.676
R1302 B.n157 B.n69 71.676
R1303 B.n153 B.n68 71.676
R1304 B.n149 B.n67 71.676
R1305 B.n145 B.n66 71.676
R1306 B.n141 B.n65 71.676
R1307 B.n137 B.n64 71.676
R1308 B.n133 B.n63 71.676
R1309 B.n129 B.n62 71.676
R1310 B.n125 B.n61 71.676
R1311 B.n121 B.n60 71.676
R1312 B.n117 B.n59 71.676
R1313 B.n113 B.n58 71.676
R1314 B.n109 B.n57 71.676
R1315 B.n105 B.n56 71.676
R1316 B.n370 B.n322 71.676
R1317 B.n374 B.n373 71.676
R1318 B.n379 B.n378 71.676
R1319 B.n382 B.n381 71.676
R1320 B.n387 B.n386 71.676
R1321 B.n390 B.n389 71.676
R1322 B.n395 B.n394 71.676
R1323 B.n398 B.n397 71.676
R1324 B.n403 B.n402 71.676
R1325 B.n406 B.n405 71.676
R1326 B.n411 B.n410 71.676
R1327 B.n414 B.n413 71.676
R1328 B.n419 B.n418 71.676
R1329 B.n422 B.n421 71.676
R1330 B.n427 B.n426 71.676
R1331 B.n430 B.n429 71.676
R1332 B.n435 B.n434 71.676
R1333 B.n438 B.n437 71.676
R1334 B.n446 B.n445 71.676
R1335 B.n449 B.n448 71.676
R1336 B.n454 B.n453 71.676
R1337 B.n457 B.n456 71.676
R1338 B.n462 B.n461 71.676
R1339 B.n465 B.n464 71.676
R1340 B.n470 B.n469 71.676
R1341 B.n473 B.n472 71.676
R1342 B.n478 B.n477 71.676
R1343 B.n481 B.n480 71.676
R1344 B.n486 B.n485 71.676
R1345 B.n489 B.n488 71.676
R1346 B.n494 B.n493 71.676
R1347 B.n497 B.n496 71.676
R1348 B.n502 B.n501 71.676
R1349 B.n505 B.n504 71.676
R1350 B.n510 B.n509 71.676
R1351 B.n513 B.n512 71.676
R1352 B.n518 B.n517 71.676
R1353 B.n521 B.n520 71.676
R1354 B.n526 B.n525 71.676
R1355 B.n529 B.n528 71.676
R1356 B.n534 B.n533 71.676
R1357 B.n537 B.n536 71.676
R1358 B.n371 B.n370 71.676
R1359 B.n373 B.n367 71.676
R1360 B.n380 B.n379 71.676
R1361 B.n381 B.n365 71.676
R1362 B.n388 B.n387 71.676
R1363 B.n389 B.n363 71.676
R1364 B.n396 B.n395 71.676
R1365 B.n397 B.n361 71.676
R1366 B.n404 B.n403 71.676
R1367 B.n405 B.n359 71.676
R1368 B.n412 B.n411 71.676
R1369 B.n413 B.n357 71.676
R1370 B.n420 B.n419 71.676
R1371 B.n421 B.n355 71.676
R1372 B.n428 B.n427 71.676
R1373 B.n429 B.n353 71.676
R1374 B.n436 B.n435 71.676
R1375 B.n437 B.n351 71.676
R1376 B.n447 B.n446 71.676
R1377 B.n448 B.n349 71.676
R1378 B.n455 B.n454 71.676
R1379 B.n456 B.n347 71.676
R1380 B.n463 B.n462 71.676
R1381 B.n464 B.n342 71.676
R1382 B.n471 B.n470 71.676
R1383 B.n472 B.n340 71.676
R1384 B.n479 B.n478 71.676
R1385 B.n480 B.n338 71.676
R1386 B.n487 B.n486 71.676
R1387 B.n488 B.n336 71.676
R1388 B.n495 B.n494 71.676
R1389 B.n496 B.n334 71.676
R1390 B.n503 B.n502 71.676
R1391 B.n504 B.n332 71.676
R1392 B.n511 B.n510 71.676
R1393 B.n512 B.n330 71.676
R1394 B.n519 B.n518 71.676
R1395 B.n520 B.n328 71.676
R1396 B.n527 B.n526 71.676
R1397 B.n528 B.n326 71.676
R1398 B.n535 B.n534 71.676
R1399 B.n536 B.n324 71.676
R1400 B.n726 B.n725 71.676
R1401 B.n726 B.n2 71.676
R1402 B.n102 B.n101 67.6854
R1403 B.n100 B.n99 67.6854
R1404 B.n344 B.n343 67.6854
R1405 B.n442 B.n441 67.6854
R1406 B.n103 B.n102 59.5399
R1407 B.n196 B.n100 59.5399
R1408 B.n345 B.n344 59.5399
R1409 B.n443 B.n442 59.5399
R1410 B.n542 B.n319 47.0002
R1411 B.n548 B.n319 47.0002
R1412 B.n548 B.n315 47.0002
R1413 B.n554 B.n315 47.0002
R1414 B.n554 B.n311 47.0002
R1415 B.n560 B.n311 47.0002
R1416 B.n560 B.n307 47.0002
R1417 B.n566 B.n307 47.0002
R1418 B.n572 B.n303 47.0002
R1419 B.n572 B.n299 47.0002
R1420 B.n578 B.n299 47.0002
R1421 B.n578 B.n295 47.0002
R1422 B.n584 B.n295 47.0002
R1423 B.n584 B.n291 47.0002
R1424 B.n590 B.n291 47.0002
R1425 B.n590 B.n287 47.0002
R1426 B.n596 B.n287 47.0002
R1427 B.n596 B.n283 47.0002
R1428 B.n603 B.n283 47.0002
R1429 B.n603 B.n602 47.0002
R1430 B.n609 B.n276 47.0002
R1431 B.n616 B.n276 47.0002
R1432 B.n616 B.n272 47.0002
R1433 B.n622 B.n272 47.0002
R1434 B.n622 B.n4 47.0002
R1435 B.n724 B.n4 47.0002
R1436 B.n724 B.n723 47.0002
R1437 B.n723 B.n722 47.0002
R1438 B.n722 B.n8 47.0002
R1439 B.n12 B.n8 47.0002
R1440 B.n715 B.n12 47.0002
R1441 B.n715 B.n714 47.0002
R1442 B.n714 B.n713 47.0002
R1443 B.n707 B.n19 47.0002
R1444 B.n707 B.n706 47.0002
R1445 B.n706 B.n705 47.0002
R1446 B.n705 B.n23 47.0002
R1447 B.n699 B.n23 47.0002
R1448 B.n699 B.n698 47.0002
R1449 B.n698 B.n697 47.0002
R1450 B.n697 B.n30 47.0002
R1451 B.n691 B.n30 47.0002
R1452 B.n691 B.n690 47.0002
R1453 B.n690 B.n689 47.0002
R1454 B.n689 B.n37 47.0002
R1455 B.n683 B.n682 47.0002
R1456 B.n682 B.n681 47.0002
R1457 B.n681 B.n44 47.0002
R1458 B.n675 B.n44 47.0002
R1459 B.n675 B.n674 47.0002
R1460 B.n674 B.n673 47.0002
R1461 B.n673 B.n51 47.0002
R1462 B.n667 B.n51 47.0002
R1463 B.n602 B.t1 35.9414
R1464 B.n19 B.t0 35.9414
R1465 B.t3 B.n303 33.1768
R1466 B.t10 B.n37 33.1768
R1467 B.n544 B.n321 32.9371
R1468 B.n540 B.n539 32.9371
R1469 B.n664 B.n663 32.9371
R1470 B.n669 B.n53 32.9371
R1471 B B.n727 18.0485
R1472 B.n566 B.t3 13.8239
R1473 B.n683 B.t10 13.8239
R1474 B.n609 B.t1 11.0593
R1475 B.n713 B.t0 11.0593
R1476 B.n545 B.n544 10.6151
R1477 B.n546 B.n545 10.6151
R1478 B.n546 B.n313 10.6151
R1479 B.n556 B.n313 10.6151
R1480 B.n557 B.n556 10.6151
R1481 B.n558 B.n557 10.6151
R1482 B.n558 B.n305 10.6151
R1483 B.n568 B.n305 10.6151
R1484 B.n569 B.n568 10.6151
R1485 B.n570 B.n569 10.6151
R1486 B.n570 B.n297 10.6151
R1487 B.n580 B.n297 10.6151
R1488 B.n581 B.n580 10.6151
R1489 B.n582 B.n581 10.6151
R1490 B.n582 B.n289 10.6151
R1491 B.n592 B.n289 10.6151
R1492 B.n593 B.n592 10.6151
R1493 B.n594 B.n593 10.6151
R1494 B.n594 B.n281 10.6151
R1495 B.n605 B.n281 10.6151
R1496 B.n606 B.n605 10.6151
R1497 B.n607 B.n606 10.6151
R1498 B.n607 B.n274 10.6151
R1499 B.n618 B.n274 10.6151
R1500 B.n619 B.n618 10.6151
R1501 B.n620 B.n619 10.6151
R1502 B.n620 B.n0 10.6151
R1503 B.n369 B.n321 10.6151
R1504 B.n369 B.n368 10.6151
R1505 B.n375 B.n368 10.6151
R1506 B.n376 B.n375 10.6151
R1507 B.n377 B.n376 10.6151
R1508 B.n377 B.n366 10.6151
R1509 B.n383 B.n366 10.6151
R1510 B.n384 B.n383 10.6151
R1511 B.n385 B.n384 10.6151
R1512 B.n385 B.n364 10.6151
R1513 B.n391 B.n364 10.6151
R1514 B.n392 B.n391 10.6151
R1515 B.n393 B.n392 10.6151
R1516 B.n393 B.n362 10.6151
R1517 B.n399 B.n362 10.6151
R1518 B.n400 B.n399 10.6151
R1519 B.n401 B.n400 10.6151
R1520 B.n401 B.n360 10.6151
R1521 B.n407 B.n360 10.6151
R1522 B.n408 B.n407 10.6151
R1523 B.n409 B.n408 10.6151
R1524 B.n409 B.n358 10.6151
R1525 B.n415 B.n358 10.6151
R1526 B.n416 B.n415 10.6151
R1527 B.n417 B.n416 10.6151
R1528 B.n417 B.n356 10.6151
R1529 B.n423 B.n356 10.6151
R1530 B.n424 B.n423 10.6151
R1531 B.n425 B.n424 10.6151
R1532 B.n425 B.n354 10.6151
R1533 B.n431 B.n354 10.6151
R1534 B.n432 B.n431 10.6151
R1535 B.n433 B.n432 10.6151
R1536 B.n433 B.n352 10.6151
R1537 B.n439 B.n352 10.6151
R1538 B.n440 B.n439 10.6151
R1539 B.n444 B.n440 10.6151
R1540 B.n450 B.n350 10.6151
R1541 B.n451 B.n450 10.6151
R1542 B.n452 B.n451 10.6151
R1543 B.n452 B.n348 10.6151
R1544 B.n458 B.n348 10.6151
R1545 B.n459 B.n458 10.6151
R1546 B.n460 B.n459 10.6151
R1547 B.n460 B.n346 10.6151
R1548 B.n467 B.n466 10.6151
R1549 B.n468 B.n467 10.6151
R1550 B.n468 B.n341 10.6151
R1551 B.n474 B.n341 10.6151
R1552 B.n475 B.n474 10.6151
R1553 B.n476 B.n475 10.6151
R1554 B.n476 B.n339 10.6151
R1555 B.n482 B.n339 10.6151
R1556 B.n483 B.n482 10.6151
R1557 B.n484 B.n483 10.6151
R1558 B.n484 B.n337 10.6151
R1559 B.n490 B.n337 10.6151
R1560 B.n491 B.n490 10.6151
R1561 B.n492 B.n491 10.6151
R1562 B.n492 B.n335 10.6151
R1563 B.n498 B.n335 10.6151
R1564 B.n499 B.n498 10.6151
R1565 B.n500 B.n499 10.6151
R1566 B.n500 B.n333 10.6151
R1567 B.n506 B.n333 10.6151
R1568 B.n507 B.n506 10.6151
R1569 B.n508 B.n507 10.6151
R1570 B.n508 B.n331 10.6151
R1571 B.n514 B.n331 10.6151
R1572 B.n515 B.n514 10.6151
R1573 B.n516 B.n515 10.6151
R1574 B.n516 B.n329 10.6151
R1575 B.n522 B.n329 10.6151
R1576 B.n523 B.n522 10.6151
R1577 B.n524 B.n523 10.6151
R1578 B.n524 B.n327 10.6151
R1579 B.n530 B.n327 10.6151
R1580 B.n531 B.n530 10.6151
R1581 B.n532 B.n531 10.6151
R1582 B.n532 B.n325 10.6151
R1583 B.n538 B.n325 10.6151
R1584 B.n539 B.n538 10.6151
R1585 B.n540 B.n317 10.6151
R1586 B.n550 B.n317 10.6151
R1587 B.n551 B.n550 10.6151
R1588 B.n552 B.n551 10.6151
R1589 B.n552 B.n309 10.6151
R1590 B.n562 B.n309 10.6151
R1591 B.n563 B.n562 10.6151
R1592 B.n564 B.n563 10.6151
R1593 B.n564 B.n301 10.6151
R1594 B.n574 B.n301 10.6151
R1595 B.n575 B.n574 10.6151
R1596 B.n576 B.n575 10.6151
R1597 B.n576 B.n293 10.6151
R1598 B.n586 B.n293 10.6151
R1599 B.n587 B.n586 10.6151
R1600 B.n588 B.n587 10.6151
R1601 B.n588 B.n285 10.6151
R1602 B.n598 B.n285 10.6151
R1603 B.n599 B.n598 10.6151
R1604 B.n600 B.n599 10.6151
R1605 B.n600 B.n278 10.6151
R1606 B.n611 B.n278 10.6151
R1607 B.n612 B.n611 10.6151
R1608 B.n614 B.n612 10.6151
R1609 B.n614 B.n613 10.6151
R1610 B.n613 B.n270 10.6151
R1611 B.n625 B.n270 10.6151
R1612 B.n626 B.n625 10.6151
R1613 B.n627 B.n626 10.6151
R1614 B.n628 B.n627 10.6151
R1615 B.n629 B.n628 10.6151
R1616 B.n632 B.n629 10.6151
R1617 B.n633 B.n632 10.6151
R1618 B.n634 B.n633 10.6151
R1619 B.n635 B.n634 10.6151
R1620 B.n637 B.n635 10.6151
R1621 B.n638 B.n637 10.6151
R1622 B.n639 B.n638 10.6151
R1623 B.n640 B.n639 10.6151
R1624 B.n642 B.n640 10.6151
R1625 B.n643 B.n642 10.6151
R1626 B.n644 B.n643 10.6151
R1627 B.n645 B.n644 10.6151
R1628 B.n647 B.n645 10.6151
R1629 B.n648 B.n647 10.6151
R1630 B.n649 B.n648 10.6151
R1631 B.n650 B.n649 10.6151
R1632 B.n652 B.n650 10.6151
R1633 B.n653 B.n652 10.6151
R1634 B.n654 B.n653 10.6151
R1635 B.n655 B.n654 10.6151
R1636 B.n657 B.n655 10.6151
R1637 B.n658 B.n657 10.6151
R1638 B.n659 B.n658 10.6151
R1639 B.n660 B.n659 10.6151
R1640 B.n662 B.n660 10.6151
R1641 B.n663 B.n662 10.6151
R1642 B.n719 B.n1 10.6151
R1643 B.n719 B.n718 10.6151
R1644 B.n718 B.n717 10.6151
R1645 B.n717 B.n10 10.6151
R1646 B.n711 B.n10 10.6151
R1647 B.n711 B.n710 10.6151
R1648 B.n710 B.n709 10.6151
R1649 B.n709 B.n17 10.6151
R1650 B.n703 B.n17 10.6151
R1651 B.n703 B.n702 10.6151
R1652 B.n702 B.n701 10.6151
R1653 B.n701 B.n25 10.6151
R1654 B.n695 B.n25 10.6151
R1655 B.n695 B.n694 10.6151
R1656 B.n694 B.n693 10.6151
R1657 B.n693 B.n32 10.6151
R1658 B.n687 B.n32 10.6151
R1659 B.n687 B.n686 10.6151
R1660 B.n686 B.n685 10.6151
R1661 B.n685 B.n39 10.6151
R1662 B.n679 B.n39 10.6151
R1663 B.n679 B.n678 10.6151
R1664 B.n678 B.n677 10.6151
R1665 B.n677 B.n46 10.6151
R1666 B.n671 B.n46 10.6151
R1667 B.n671 B.n670 10.6151
R1668 B.n670 B.n669 10.6151
R1669 B.n104 B.n53 10.6151
R1670 B.n107 B.n104 10.6151
R1671 B.n108 B.n107 10.6151
R1672 B.n111 B.n108 10.6151
R1673 B.n112 B.n111 10.6151
R1674 B.n115 B.n112 10.6151
R1675 B.n116 B.n115 10.6151
R1676 B.n119 B.n116 10.6151
R1677 B.n120 B.n119 10.6151
R1678 B.n123 B.n120 10.6151
R1679 B.n124 B.n123 10.6151
R1680 B.n127 B.n124 10.6151
R1681 B.n128 B.n127 10.6151
R1682 B.n131 B.n128 10.6151
R1683 B.n132 B.n131 10.6151
R1684 B.n135 B.n132 10.6151
R1685 B.n136 B.n135 10.6151
R1686 B.n139 B.n136 10.6151
R1687 B.n140 B.n139 10.6151
R1688 B.n143 B.n140 10.6151
R1689 B.n144 B.n143 10.6151
R1690 B.n147 B.n144 10.6151
R1691 B.n148 B.n147 10.6151
R1692 B.n151 B.n148 10.6151
R1693 B.n152 B.n151 10.6151
R1694 B.n155 B.n152 10.6151
R1695 B.n156 B.n155 10.6151
R1696 B.n159 B.n156 10.6151
R1697 B.n160 B.n159 10.6151
R1698 B.n163 B.n160 10.6151
R1699 B.n164 B.n163 10.6151
R1700 B.n167 B.n164 10.6151
R1701 B.n168 B.n167 10.6151
R1702 B.n171 B.n168 10.6151
R1703 B.n172 B.n171 10.6151
R1704 B.n175 B.n172 10.6151
R1705 B.n176 B.n175 10.6151
R1706 B.n180 B.n179 10.6151
R1707 B.n183 B.n180 10.6151
R1708 B.n184 B.n183 10.6151
R1709 B.n187 B.n184 10.6151
R1710 B.n188 B.n187 10.6151
R1711 B.n191 B.n188 10.6151
R1712 B.n192 B.n191 10.6151
R1713 B.n195 B.n192 10.6151
R1714 B.n200 B.n197 10.6151
R1715 B.n201 B.n200 10.6151
R1716 B.n204 B.n201 10.6151
R1717 B.n205 B.n204 10.6151
R1718 B.n208 B.n205 10.6151
R1719 B.n209 B.n208 10.6151
R1720 B.n212 B.n209 10.6151
R1721 B.n213 B.n212 10.6151
R1722 B.n216 B.n213 10.6151
R1723 B.n217 B.n216 10.6151
R1724 B.n220 B.n217 10.6151
R1725 B.n221 B.n220 10.6151
R1726 B.n224 B.n221 10.6151
R1727 B.n225 B.n224 10.6151
R1728 B.n228 B.n225 10.6151
R1729 B.n229 B.n228 10.6151
R1730 B.n232 B.n229 10.6151
R1731 B.n233 B.n232 10.6151
R1732 B.n236 B.n233 10.6151
R1733 B.n237 B.n236 10.6151
R1734 B.n240 B.n237 10.6151
R1735 B.n241 B.n240 10.6151
R1736 B.n244 B.n241 10.6151
R1737 B.n245 B.n244 10.6151
R1738 B.n248 B.n245 10.6151
R1739 B.n249 B.n248 10.6151
R1740 B.n252 B.n249 10.6151
R1741 B.n253 B.n252 10.6151
R1742 B.n256 B.n253 10.6151
R1743 B.n257 B.n256 10.6151
R1744 B.n260 B.n257 10.6151
R1745 B.n261 B.n260 10.6151
R1746 B.n264 B.n261 10.6151
R1747 B.n265 B.n264 10.6151
R1748 B.n268 B.n265 10.6151
R1749 B.n269 B.n268 10.6151
R1750 B.n664 B.n269 10.6151
R1751 B.n727 B.n0 8.11757
R1752 B.n727 B.n1 8.11757
R1753 B.n443 B.n350 6.5566
R1754 B.n346 B.n345 6.5566
R1755 B.n179 B.n103 6.5566
R1756 B.n196 B.n195 6.5566
R1757 B.n444 B.n443 4.05904
R1758 B.n466 B.n345 4.05904
R1759 B.n176 B.n103 4.05904
R1760 B.n197 B.n196 4.05904
R1761 VN VN.t1 164.897
R1762 VN VN.t0 120.403
R1763 VDD2.n109 VDD2.n57 289.615
R1764 VDD2.n52 VDD2.n0 289.615
R1765 VDD2.n110 VDD2.n109 185
R1766 VDD2.n108 VDD2.n107 185
R1767 VDD2.n61 VDD2.n60 185
R1768 VDD2.n102 VDD2.n101 185
R1769 VDD2.n100 VDD2.n99 185
R1770 VDD2.n98 VDD2.n64 185
R1771 VDD2.n68 VDD2.n65 185
R1772 VDD2.n93 VDD2.n92 185
R1773 VDD2.n91 VDD2.n90 185
R1774 VDD2.n70 VDD2.n69 185
R1775 VDD2.n85 VDD2.n84 185
R1776 VDD2.n83 VDD2.n82 185
R1777 VDD2.n74 VDD2.n73 185
R1778 VDD2.n77 VDD2.n76 185
R1779 VDD2.n19 VDD2.n18 185
R1780 VDD2.n16 VDD2.n15 185
R1781 VDD2.n25 VDD2.n24 185
R1782 VDD2.n27 VDD2.n26 185
R1783 VDD2.n12 VDD2.n11 185
R1784 VDD2.n33 VDD2.n32 185
R1785 VDD2.n36 VDD2.n35 185
R1786 VDD2.n34 VDD2.n8 185
R1787 VDD2.n41 VDD2.n7 185
R1788 VDD2.n43 VDD2.n42 185
R1789 VDD2.n45 VDD2.n44 185
R1790 VDD2.n4 VDD2.n3 185
R1791 VDD2.n51 VDD2.n50 185
R1792 VDD2.n53 VDD2.n52 185
R1793 VDD2.t0 VDD2.n75 149.524
R1794 VDD2.t1 VDD2.n17 149.524
R1795 VDD2.n109 VDD2.n108 104.615
R1796 VDD2.n108 VDD2.n60 104.615
R1797 VDD2.n101 VDD2.n60 104.615
R1798 VDD2.n101 VDD2.n100 104.615
R1799 VDD2.n100 VDD2.n64 104.615
R1800 VDD2.n68 VDD2.n64 104.615
R1801 VDD2.n92 VDD2.n68 104.615
R1802 VDD2.n92 VDD2.n91 104.615
R1803 VDD2.n91 VDD2.n69 104.615
R1804 VDD2.n84 VDD2.n69 104.615
R1805 VDD2.n84 VDD2.n83 104.615
R1806 VDD2.n83 VDD2.n73 104.615
R1807 VDD2.n76 VDD2.n73 104.615
R1808 VDD2.n18 VDD2.n15 104.615
R1809 VDD2.n25 VDD2.n15 104.615
R1810 VDD2.n26 VDD2.n25 104.615
R1811 VDD2.n26 VDD2.n11 104.615
R1812 VDD2.n33 VDD2.n11 104.615
R1813 VDD2.n35 VDD2.n33 104.615
R1814 VDD2.n35 VDD2.n34 104.615
R1815 VDD2.n34 VDD2.n7 104.615
R1816 VDD2.n43 VDD2.n7 104.615
R1817 VDD2.n44 VDD2.n43 104.615
R1818 VDD2.n44 VDD2.n3 104.615
R1819 VDD2.n51 VDD2.n3 104.615
R1820 VDD2.n52 VDD2.n51 104.615
R1821 VDD2.n114 VDD2.n56 86.9375
R1822 VDD2.n76 VDD2.t0 52.3082
R1823 VDD2.n18 VDD2.t1 52.3082
R1824 VDD2.n114 VDD2.n113 48.0884
R1825 VDD2.n99 VDD2.n98 13.1884
R1826 VDD2.n42 VDD2.n41 13.1884
R1827 VDD2.n102 VDD2.n63 12.8005
R1828 VDD2.n97 VDD2.n65 12.8005
R1829 VDD2.n40 VDD2.n8 12.8005
R1830 VDD2.n45 VDD2.n6 12.8005
R1831 VDD2.n103 VDD2.n61 12.0247
R1832 VDD2.n94 VDD2.n93 12.0247
R1833 VDD2.n37 VDD2.n36 12.0247
R1834 VDD2.n46 VDD2.n4 12.0247
R1835 VDD2.n107 VDD2.n106 11.249
R1836 VDD2.n90 VDD2.n67 11.249
R1837 VDD2.n32 VDD2.n10 11.249
R1838 VDD2.n50 VDD2.n49 11.249
R1839 VDD2.n110 VDD2.n59 10.4732
R1840 VDD2.n89 VDD2.n70 10.4732
R1841 VDD2.n31 VDD2.n12 10.4732
R1842 VDD2.n53 VDD2.n2 10.4732
R1843 VDD2.n77 VDD2.n75 10.2747
R1844 VDD2.n19 VDD2.n17 10.2747
R1845 VDD2.n111 VDD2.n57 9.69747
R1846 VDD2.n86 VDD2.n85 9.69747
R1847 VDD2.n28 VDD2.n27 9.69747
R1848 VDD2.n54 VDD2.n0 9.69747
R1849 VDD2.n113 VDD2.n112 9.45567
R1850 VDD2.n56 VDD2.n55 9.45567
R1851 VDD2.n79 VDD2.n78 9.3005
R1852 VDD2.n81 VDD2.n80 9.3005
R1853 VDD2.n72 VDD2.n71 9.3005
R1854 VDD2.n87 VDD2.n86 9.3005
R1855 VDD2.n89 VDD2.n88 9.3005
R1856 VDD2.n67 VDD2.n66 9.3005
R1857 VDD2.n95 VDD2.n94 9.3005
R1858 VDD2.n97 VDD2.n96 9.3005
R1859 VDD2.n112 VDD2.n111 9.3005
R1860 VDD2.n59 VDD2.n58 9.3005
R1861 VDD2.n106 VDD2.n105 9.3005
R1862 VDD2.n104 VDD2.n103 9.3005
R1863 VDD2.n63 VDD2.n62 9.3005
R1864 VDD2.n55 VDD2.n54 9.3005
R1865 VDD2.n2 VDD2.n1 9.3005
R1866 VDD2.n49 VDD2.n48 9.3005
R1867 VDD2.n47 VDD2.n46 9.3005
R1868 VDD2.n6 VDD2.n5 9.3005
R1869 VDD2.n21 VDD2.n20 9.3005
R1870 VDD2.n23 VDD2.n22 9.3005
R1871 VDD2.n14 VDD2.n13 9.3005
R1872 VDD2.n29 VDD2.n28 9.3005
R1873 VDD2.n31 VDD2.n30 9.3005
R1874 VDD2.n10 VDD2.n9 9.3005
R1875 VDD2.n38 VDD2.n37 9.3005
R1876 VDD2.n40 VDD2.n39 9.3005
R1877 VDD2.n82 VDD2.n72 8.92171
R1878 VDD2.n24 VDD2.n14 8.92171
R1879 VDD2.n81 VDD2.n74 8.14595
R1880 VDD2.n23 VDD2.n16 8.14595
R1881 VDD2.n78 VDD2.n77 7.3702
R1882 VDD2.n20 VDD2.n19 7.3702
R1883 VDD2.n78 VDD2.n74 5.81868
R1884 VDD2.n20 VDD2.n16 5.81868
R1885 VDD2.n82 VDD2.n81 5.04292
R1886 VDD2.n24 VDD2.n23 5.04292
R1887 VDD2.n113 VDD2.n57 4.26717
R1888 VDD2.n85 VDD2.n72 4.26717
R1889 VDD2.n27 VDD2.n14 4.26717
R1890 VDD2.n56 VDD2.n0 4.26717
R1891 VDD2.n111 VDD2.n110 3.49141
R1892 VDD2.n86 VDD2.n70 3.49141
R1893 VDD2.n28 VDD2.n12 3.49141
R1894 VDD2.n54 VDD2.n53 3.49141
R1895 VDD2.n79 VDD2.n75 2.84303
R1896 VDD2.n21 VDD2.n17 2.84303
R1897 VDD2.n107 VDD2.n59 2.71565
R1898 VDD2.n90 VDD2.n89 2.71565
R1899 VDD2.n32 VDD2.n31 2.71565
R1900 VDD2.n50 VDD2.n2 2.71565
R1901 VDD2.n106 VDD2.n61 1.93989
R1902 VDD2.n93 VDD2.n67 1.93989
R1903 VDD2.n36 VDD2.n10 1.93989
R1904 VDD2.n49 VDD2.n4 1.93989
R1905 VDD2.n103 VDD2.n102 1.16414
R1906 VDD2.n94 VDD2.n65 1.16414
R1907 VDD2.n37 VDD2.n8 1.16414
R1908 VDD2.n46 VDD2.n45 1.16414
R1909 VDD2 VDD2.n114 0.810845
R1910 VDD2.n99 VDD2.n63 0.388379
R1911 VDD2.n98 VDD2.n97 0.388379
R1912 VDD2.n41 VDD2.n40 0.388379
R1913 VDD2.n42 VDD2.n6 0.388379
R1914 VDD2.n112 VDD2.n58 0.155672
R1915 VDD2.n105 VDD2.n58 0.155672
R1916 VDD2.n105 VDD2.n104 0.155672
R1917 VDD2.n104 VDD2.n62 0.155672
R1918 VDD2.n96 VDD2.n62 0.155672
R1919 VDD2.n96 VDD2.n95 0.155672
R1920 VDD2.n95 VDD2.n66 0.155672
R1921 VDD2.n88 VDD2.n66 0.155672
R1922 VDD2.n88 VDD2.n87 0.155672
R1923 VDD2.n87 VDD2.n71 0.155672
R1924 VDD2.n80 VDD2.n71 0.155672
R1925 VDD2.n80 VDD2.n79 0.155672
R1926 VDD2.n22 VDD2.n21 0.155672
R1927 VDD2.n22 VDD2.n13 0.155672
R1928 VDD2.n29 VDD2.n13 0.155672
R1929 VDD2.n30 VDD2.n29 0.155672
R1930 VDD2.n30 VDD2.n9 0.155672
R1931 VDD2.n38 VDD2.n9 0.155672
R1932 VDD2.n39 VDD2.n38 0.155672
R1933 VDD2.n39 VDD2.n5 0.155672
R1934 VDD2.n47 VDD2.n5 0.155672
R1935 VDD2.n48 VDD2.n47 0.155672
R1936 VDD2.n48 VDD2.n1 0.155672
R1937 VDD2.n55 VDD2.n1 0.155672
C0 VP VDD2 0.356161f
C1 VDD1 VDD2 0.742601f
C2 VP VDD1 2.76814f
C3 VTAIL VDD2 4.87224f
C4 VN VDD2 2.56211f
C5 VTAIL VP 2.34422f
C6 VTAIL VDD1 4.81709f
C7 VN VP 5.47415f
C8 VN VDD1 0.148045f
C9 VN VTAIL 2.32998f
C10 VDD2 B 4.384187f
C11 VDD1 B 7.13353f
C12 VTAIL B 7.078322f
C13 VN B 10.99576f
C14 VP B 7.01793f
C15 VDD2.n0 B 0.027371f
C16 VDD2.n1 B 0.020663f
C17 VDD2.n2 B 0.011103f
C18 VDD2.n3 B 0.026245f
C19 VDD2.n4 B 0.011757f
C20 VDD2.n5 B 0.020663f
C21 VDD2.n6 B 0.011103f
C22 VDD2.n7 B 0.026245f
C23 VDD2.n8 B 0.011757f
C24 VDD2.n9 B 0.020663f
C25 VDD2.n10 B 0.011103f
C26 VDD2.n11 B 0.026245f
C27 VDD2.n12 B 0.011757f
C28 VDD2.n13 B 0.020663f
C29 VDD2.n14 B 0.011103f
C30 VDD2.n15 B 0.026245f
C31 VDD2.n16 B 0.011757f
C32 VDD2.n17 B 0.138192f
C33 VDD2.t1 B 0.044175f
C34 VDD2.n18 B 0.019684f
C35 VDD2.n19 B 0.018553f
C36 VDD2.n20 B 0.011103f
C37 VDD2.n21 B 0.91743f
C38 VDD2.n22 B 0.020663f
C39 VDD2.n23 B 0.011103f
C40 VDD2.n24 B 0.011757f
C41 VDD2.n25 B 0.026245f
C42 VDD2.n26 B 0.026245f
C43 VDD2.n27 B 0.011757f
C44 VDD2.n28 B 0.011103f
C45 VDD2.n29 B 0.020663f
C46 VDD2.n30 B 0.020663f
C47 VDD2.n31 B 0.011103f
C48 VDD2.n32 B 0.011757f
C49 VDD2.n33 B 0.026245f
C50 VDD2.n34 B 0.026245f
C51 VDD2.n35 B 0.026245f
C52 VDD2.n36 B 0.011757f
C53 VDD2.n37 B 0.011103f
C54 VDD2.n38 B 0.020663f
C55 VDD2.n39 B 0.020663f
C56 VDD2.n40 B 0.011103f
C57 VDD2.n41 B 0.01143f
C58 VDD2.n42 B 0.01143f
C59 VDD2.n43 B 0.026245f
C60 VDD2.n44 B 0.026245f
C61 VDD2.n45 B 0.011757f
C62 VDD2.n46 B 0.011103f
C63 VDD2.n47 B 0.020663f
C64 VDD2.n48 B 0.020663f
C65 VDD2.n49 B 0.011103f
C66 VDD2.n50 B 0.011757f
C67 VDD2.n51 B 0.026245f
C68 VDD2.n52 B 0.053857f
C69 VDD2.n53 B 0.011757f
C70 VDD2.n54 B 0.011103f
C71 VDD2.n55 B 0.046633f
C72 VDD2.n56 B 0.600749f
C73 VDD2.n57 B 0.027371f
C74 VDD2.n58 B 0.020663f
C75 VDD2.n59 B 0.011103f
C76 VDD2.n60 B 0.026245f
C77 VDD2.n61 B 0.011757f
C78 VDD2.n62 B 0.020663f
C79 VDD2.n63 B 0.011103f
C80 VDD2.n64 B 0.026245f
C81 VDD2.n65 B 0.011757f
C82 VDD2.n66 B 0.020663f
C83 VDD2.n67 B 0.011103f
C84 VDD2.n68 B 0.026245f
C85 VDD2.n69 B 0.026245f
C86 VDD2.n70 B 0.011757f
C87 VDD2.n71 B 0.020663f
C88 VDD2.n72 B 0.011103f
C89 VDD2.n73 B 0.026245f
C90 VDD2.n74 B 0.011757f
C91 VDD2.n75 B 0.138192f
C92 VDD2.t0 B 0.044175f
C93 VDD2.n76 B 0.019684f
C94 VDD2.n77 B 0.018553f
C95 VDD2.n78 B 0.011103f
C96 VDD2.n79 B 0.91743f
C97 VDD2.n80 B 0.020663f
C98 VDD2.n81 B 0.011103f
C99 VDD2.n82 B 0.011757f
C100 VDD2.n83 B 0.026245f
C101 VDD2.n84 B 0.026245f
C102 VDD2.n85 B 0.011757f
C103 VDD2.n86 B 0.011103f
C104 VDD2.n87 B 0.020663f
C105 VDD2.n88 B 0.020663f
C106 VDD2.n89 B 0.011103f
C107 VDD2.n90 B 0.011757f
C108 VDD2.n91 B 0.026245f
C109 VDD2.n92 B 0.026245f
C110 VDD2.n93 B 0.011757f
C111 VDD2.n94 B 0.011103f
C112 VDD2.n95 B 0.020663f
C113 VDD2.n96 B 0.020663f
C114 VDD2.n97 B 0.011103f
C115 VDD2.n98 B 0.01143f
C116 VDD2.n99 B 0.01143f
C117 VDD2.n100 B 0.026245f
C118 VDD2.n101 B 0.026245f
C119 VDD2.n102 B 0.011757f
C120 VDD2.n103 B 0.011103f
C121 VDD2.n104 B 0.020663f
C122 VDD2.n105 B 0.020663f
C123 VDD2.n106 B 0.011103f
C124 VDD2.n107 B 0.011757f
C125 VDD2.n108 B 0.026245f
C126 VDD2.n109 B 0.053857f
C127 VDD2.n110 B 0.011757f
C128 VDD2.n111 B 0.011103f
C129 VDD2.n112 B 0.046633f
C130 VDD2.n113 B 0.044073f
C131 VDD2.n114 B 2.49118f
C132 VN.t0 B 2.92122f
C133 VN.t1 B 3.53304f
C134 VDD1.n0 B 0.027457f
C135 VDD1.n1 B 0.020728f
C136 VDD1.n2 B 0.011138f
C137 VDD1.n3 B 0.026327f
C138 VDD1.n4 B 0.011793f
C139 VDD1.n5 B 0.020728f
C140 VDD1.n6 B 0.011138f
C141 VDD1.n7 B 0.026327f
C142 VDD1.n8 B 0.011793f
C143 VDD1.n9 B 0.020728f
C144 VDD1.n10 B 0.011138f
C145 VDD1.n11 B 0.026327f
C146 VDD1.n12 B 0.026327f
C147 VDD1.n13 B 0.011793f
C148 VDD1.n14 B 0.020728f
C149 VDD1.n15 B 0.011138f
C150 VDD1.n16 B 0.026327f
C151 VDD1.n17 B 0.011793f
C152 VDD1.n18 B 0.138624f
C153 VDD1.t1 B 0.044313f
C154 VDD1.n19 B 0.019745f
C155 VDD1.n20 B 0.018611f
C156 VDD1.n21 B 0.011138f
C157 VDD1.n22 B 0.920297f
C158 VDD1.n23 B 0.020728f
C159 VDD1.n24 B 0.011138f
C160 VDD1.n25 B 0.011793f
C161 VDD1.n26 B 0.026327f
C162 VDD1.n27 B 0.026327f
C163 VDD1.n28 B 0.011793f
C164 VDD1.n29 B 0.011138f
C165 VDD1.n30 B 0.020728f
C166 VDD1.n31 B 0.020728f
C167 VDD1.n32 B 0.011138f
C168 VDD1.n33 B 0.011793f
C169 VDD1.n34 B 0.026327f
C170 VDD1.n35 B 0.026327f
C171 VDD1.n36 B 0.011793f
C172 VDD1.n37 B 0.011138f
C173 VDD1.n38 B 0.020728f
C174 VDD1.n39 B 0.020728f
C175 VDD1.n40 B 0.011138f
C176 VDD1.n41 B 0.011466f
C177 VDD1.n42 B 0.011466f
C178 VDD1.n43 B 0.026327f
C179 VDD1.n44 B 0.026327f
C180 VDD1.n45 B 0.011793f
C181 VDD1.n46 B 0.011138f
C182 VDD1.n47 B 0.020728f
C183 VDD1.n48 B 0.020728f
C184 VDD1.n49 B 0.011138f
C185 VDD1.n50 B 0.011793f
C186 VDD1.n51 B 0.026327f
C187 VDD1.n52 B 0.054025f
C188 VDD1.n53 B 0.011793f
C189 VDD1.n54 B 0.011138f
C190 VDD1.n55 B 0.046779f
C191 VDD1.n56 B 0.045758f
C192 VDD1.n57 B 0.027457f
C193 VDD1.n58 B 0.020728f
C194 VDD1.n59 B 0.011138f
C195 VDD1.n60 B 0.026327f
C196 VDD1.n61 B 0.011793f
C197 VDD1.n62 B 0.020728f
C198 VDD1.n63 B 0.011138f
C199 VDD1.n64 B 0.026327f
C200 VDD1.n65 B 0.011793f
C201 VDD1.n66 B 0.020728f
C202 VDD1.n67 B 0.011138f
C203 VDD1.n68 B 0.026327f
C204 VDD1.n69 B 0.011793f
C205 VDD1.n70 B 0.020728f
C206 VDD1.n71 B 0.011138f
C207 VDD1.n72 B 0.026327f
C208 VDD1.n73 B 0.011793f
C209 VDD1.n74 B 0.138624f
C210 VDD1.t0 B 0.044313f
C211 VDD1.n75 B 0.019745f
C212 VDD1.n76 B 0.018611f
C213 VDD1.n77 B 0.011138f
C214 VDD1.n78 B 0.920297f
C215 VDD1.n79 B 0.020728f
C216 VDD1.n80 B 0.011138f
C217 VDD1.n81 B 0.011793f
C218 VDD1.n82 B 0.026327f
C219 VDD1.n83 B 0.026327f
C220 VDD1.n84 B 0.011793f
C221 VDD1.n85 B 0.011138f
C222 VDD1.n86 B 0.020728f
C223 VDD1.n87 B 0.020728f
C224 VDD1.n88 B 0.011138f
C225 VDD1.n89 B 0.011793f
C226 VDD1.n90 B 0.026327f
C227 VDD1.n91 B 0.026327f
C228 VDD1.n92 B 0.026327f
C229 VDD1.n93 B 0.011793f
C230 VDD1.n94 B 0.011138f
C231 VDD1.n95 B 0.020728f
C232 VDD1.n96 B 0.020728f
C233 VDD1.n97 B 0.011138f
C234 VDD1.n98 B 0.011466f
C235 VDD1.n99 B 0.011466f
C236 VDD1.n100 B 0.026327f
C237 VDD1.n101 B 0.026327f
C238 VDD1.n102 B 0.011793f
C239 VDD1.n103 B 0.011138f
C240 VDD1.n104 B 0.020728f
C241 VDD1.n105 B 0.020728f
C242 VDD1.n106 B 0.011138f
C243 VDD1.n107 B 0.011793f
C244 VDD1.n108 B 0.026327f
C245 VDD1.n109 B 0.054025f
C246 VDD1.n110 B 0.011793f
C247 VDD1.n111 B 0.011138f
C248 VDD1.n112 B 0.046779f
C249 VDD1.n113 B 0.646709f
C250 VTAIL.n0 B 0.028161f
C251 VTAIL.n1 B 0.021259f
C252 VTAIL.n2 B 0.011424f
C253 VTAIL.n3 B 0.027002f
C254 VTAIL.n4 B 0.012096f
C255 VTAIL.n5 B 0.021259f
C256 VTAIL.n6 B 0.011424f
C257 VTAIL.n7 B 0.027002f
C258 VTAIL.n8 B 0.012096f
C259 VTAIL.n9 B 0.021259f
C260 VTAIL.n10 B 0.011424f
C261 VTAIL.n11 B 0.027002f
C262 VTAIL.n12 B 0.012096f
C263 VTAIL.n13 B 0.021259f
C264 VTAIL.n14 B 0.011424f
C265 VTAIL.n15 B 0.027002f
C266 VTAIL.n16 B 0.012096f
C267 VTAIL.n17 B 0.142177f
C268 VTAIL.t3 B 0.045449f
C269 VTAIL.n18 B 0.020251f
C270 VTAIL.n19 B 0.019088f
C271 VTAIL.n20 B 0.011424f
C272 VTAIL.n21 B 0.94389f
C273 VTAIL.n22 B 0.021259f
C274 VTAIL.n23 B 0.011424f
C275 VTAIL.n24 B 0.012096f
C276 VTAIL.n25 B 0.027002f
C277 VTAIL.n26 B 0.027002f
C278 VTAIL.n27 B 0.012096f
C279 VTAIL.n28 B 0.011424f
C280 VTAIL.n29 B 0.021259f
C281 VTAIL.n30 B 0.021259f
C282 VTAIL.n31 B 0.011424f
C283 VTAIL.n32 B 0.012096f
C284 VTAIL.n33 B 0.027002f
C285 VTAIL.n34 B 0.027002f
C286 VTAIL.n35 B 0.027002f
C287 VTAIL.n36 B 0.012096f
C288 VTAIL.n37 B 0.011424f
C289 VTAIL.n38 B 0.021259f
C290 VTAIL.n39 B 0.021259f
C291 VTAIL.n40 B 0.011424f
C292 VTAIL.n41 B 0.01176f
C293 VTAIL.n42 B 0.01176f
C294 VTAIL.n43 B 0.027002f
C295 VTAIL.n44 B 0.027002f
C296 VTAIL.n45 B 0.012096f
C297 VTAIL.n46 B 0.011424f
C298 VTAIL.n47 B 0.021259f
C299 VTAIL.n48 B 0.021259f
C300 VTAIL.n49 B 0.011424f
C301 VTAIL.n50 B 0.012096f
C302 VTAIL.n51 B 0.027002f
C303 VTAIL.n52 B 0.05541f
C304 VTAIL.n53 B 0.012096f
C305 VTAIL.n54 B 0.011424f
C306 VTAIL.n55 B 0.047978f
C307 VTAIL.n56 B 0.030655f
C308 VTAIL.n57 B 1.4345f
C309 VTAIL.n58 B 0.028161f
C310 VTAIL.n59 B 0.021259f
C311 VTAIL.n60 B 0.011424f
C312 VTAIL.n61 B 0.027002f
C313 VTAIL.n62 B 0.012096f
C314 VTAIL.n63 B 0.021259f
C315 VTAIL.n64 B 0.011424f
C316 VTAIL.n65 B 0.027002f
C317 VTAIL.n66 B 0.012096f
C318 VTAIL.n67 B 0.021259f
C319 VTAIL.n68 B 0.011424f
C320 VTAIL.n69 B 0.027002f
C321 VTAIL.n70 B 0.027002f
C322 VTAIL.n71 B 0.012096f
C323 VTAIL.n72 B 0.021259f
C324 VTAIL.n73 B 0.011424f
C325 VTAIL.n74 B 0.027002f
C326 VTAIL.n75 B 0.012096f
C327 VTAIL.n76 B 0.142177f
C328 VTAIL.t1 B 0.045449f
C329 VTAIL.n77 B 0.020251f
C330 VTAIL.n78 B 0.019088f
C331 VTAIL.n79 B 0.011424f
C332 VTAIL.n80 B 0.94389f
C333 VTAIL.n81 B 0.021259f
C334 VTAIL.n82 B 0.011424f
C335 VTAIL.n83 B 0.012096f
C336 VTAIL.n84 B 0.027002f
C337 VTAIL.n85 B 0.027002f
C338 VTAIL.n86 B 0.012096f
C339 VTAIL.n87 B 0.011424f
C340 VTAIL.n88 B 0.021259f
C341 VTAIL.n89 B 0.021259f
C342 VTAIL.n90 B 0.011424f
C343 VTAIL.n91 B 0.012096f
C344 VTAIL.n92 B 0.027002f
C345 VTAIL.n93 B 0.027002f
C346 VTAIL.n94 B 0.012096f
C347 VTAIL.n95 B 0.011424f
C348 VTAIL.n96 B 0.021259f
C349 VTAIL.n97 B 0.021259f
C350 VTAIL.n98 B 0.011424f
C351 VTAIL.n99 B 0.01176f
C352 VTAIL.n100 B 0.01176f
C353 VTAIL.n101 B 0.027002f
C354 VTAIL.n102 B 0.027002f
C355 VTAIL.n103 B 0.012096f
C356 VTAIL.n104 B 0.011424f
C357 VTAIL.n105 B 0.021259f
C358 VTAIL.n106 B 0.021259f
C359 VTAIL.n107 B 0.011424f
C360 VTAIL.n108 B 0.012096f
C361 VTAIL.n109 B 0.027002f
C362 VTAIL.n110 B 0.05541f
C363 VTAIL.n111 B 0.012096f
C364 VTAIL.n112 B 0.011424f
C365 VTAIL.n113 B 0.047978f
C366 VTAIL.n114 B 0.030655f
C367 VTAIL.n115 B 1.48204f
C368 VTAIL.n116 B 0.028161f
C369 VTAIL.n117 B 0.021259f
C370 VTAIL.n118 B 0.011424f
C371 VTAIL.n119 B 0.027002f
C372 VTAIL.n120 B 0.012096f
C373 VTAIL.n121 B 0.021259f
C374 VTAIL.n122 B 0.011424f
C375 VTAIL.n123 B 0.027002f
C376 VTAIL.n124 B 0.012096f
C377 VTAIL.n125 B 0.021259f
C378 VTAIL.n126 B 0.011424f
C379 VTAIL.n127 B 0.027002f
C380 VTAIL.n128 B 0.027002f
C381 VTAIL.n129 B 0.012096f
C382 VTAIL.n130 B 0.021259f
C383 VTAIL.n131 B 0.011424f
C384 VTAIL.n132 B 0.027002f
C385 VTAIL.n133 B 0.012096f
C386 VTAIL.n134 B 0.142177f
C387 VTAIL.t2 B 0.045449f
C388 VTAIL.n135 B 0.020251f
C389 VTAIL.n136 B 0.019088f
C390 VTAIL.n137 B 0.011424f
C391 VTAIL.n138 B 0.94389f
C392 VTAIL.n139 B 0.021259f
C393 VTAIL.n140 B 0.011424f
C394 VTAIL.n141 B 0.012096f
C395 VTAIL.n142 B 0.027002f
C396 VTAIL.n143 B 0.027002f
C397 VTAIL.n144 B 0.012096f
C398 VTAIL.n145 B 0.011424f
C399 VTAIL.n146 B 0.021259f
C400 VTAIL.n147 B 0.021259f
C401 VTAIL.n148 B 0.011424f
C402 VTAIL.n149 B 0.012096f
C403 VTAIL.n150 B 0.027002f
C404 VTAIL.n151 B 0.027002f
C405 VTAIL.n152 B 0.012096f
C406 VTAIL.n153 B 0.011424f
C407 VTAIL.n154 B 0.021259f
C408 VTAIL.n155 B 0.021259f
C409 VTAIL.n156 B 0.011424f
C410 VTAIL.n157 B 0.01176f
C411 VTAIL.n158 B 0.01176f
C412 VTAIL.n159 B 0.027002f
C413 VTAIL.n160 B 0.027002f
C414 VTAIL.n161 B 0.012096f
C415 VTAIL.n162 B 0.011424f
C416 VTAIL.n163 B 0.021259f
C417 VTAIL.n164 B 0.021259f
C418 VTAIL.n165 B 0.011424f
C419 VTAIL.n166 B 0.012096f
C420 VTAIL.n167 B 0.027002f
C421 VTAIL.n168 B 0.05541f
C422 VTAIL.n169 B 0.012096f
C423 VTAIL.n170 B 0.011424f
C424 VTAIL.n171 B 0.047978f
C425 VTAIL.n172 B 0.030655f
C426 VTAIL.n173 B 1.27594f
C427 VTAIL.n174 B 0.028161f
C428 VTAIL.n175 B 0.021259f
C429 VTAIL.n176 B 0.011424f
C430 VTAIL.n177 B 0.027002f
C431 VTAIL.n178 B 0.012096f
C432 VTAIL.n179 B 0.021259f
C433 VTAIL.n180 B 0.011424f
C434 VTAIL.n181 B 0.027002f
C435 VTAIL.n182 B 0.012096f
C436 VTAIL.n183 B 0.021259f
C437 VTAIL.n184 B 0.011424f
C438 VTAIL.n185 B 0.027002f
C439 VTAIL.n186 B 0.012096f
C440 VTAIL.n187 B 0.021259f
C441 VTAIL.n188 B 0.011424f
C442 VTAIL.n189 B 0.027002f
C443 VTAIL.n190 B 0.012096f
C444 VTAIL.n191 B 0.142177f
C445 VTAIL.t0 B 0.045449f
C446 VTAIL.n192 B 0.020251f
C447 VTAIL.n193 B 0.019088f
C448 VTAIL.n194 B 0.011424f
C449 VTAIL.n195 B 0.94389f
C450 VTAIL.n196 B 0.021259f
C451 VTAIL.n197 B 0.011424f
C452 VTAIL.n198 B 0.012096f
C453 VTAIL.n199 B 0.027002f
C454 VTAIL.n200 B 0.027002f
C455 VTAIL.n201 B 0.012096f
C456 VTAIL.n202 B 0.011424f
C457 VTAIL.n203 B 0.021259f
C458 VTAIL.n204 B 0.021259f
C459 VTAIL.n205 B 0.011424f
C460 VTAIL.n206 B 0.012096f
C461 VTAIL.n207 B 0.027002f
C462 VTAIL.n208 B 0.027002f
C463 VTAIL.n209 B 0.027002f
C464 VTAIL.n210 B 0.012096f
C465 VTAIL.n211 B 0.011424f
C466 VTAIL.n212 B 0.021259f
C467 VTAIL.n213 B 0.021259f
C468 VTAIL.n214 B 0.011424f
C469 VTAIL.n215 B 0.01176f
C470 VTAIL.n216 B 0.01176f
C471 VTAIL.n217 B 0.027002f
C472 VTAIL.n218 B 0.027002f
C473 VTAIL.n219 B 0.012096f
C474 VTAIL.n220 B 0.011424f
C475 VTAIL.n221 B 0.021259f
C476 VTAIL.n222 B 0.021259f
C477 VTAIL.n223 B 0.011424f
C478 VTAIL.n224 B 0.012096f
C479 VTAIL.n225 B 0.027002f
C480 VTAIL.n226 B 0.05541f
C481 VTAIL.n227 B 0.012096f
C482 VTAIL.n228 B 0.011424f
C483 VTAIL.n229 B 0.047978f
C484 VTAIL.n230 B 0.030655f
C485 VTAIL.n231 B 1.18824f
C486 VP.t0 B 3.61453f
C487 VP.t1 B 2.98455f
C488 VP.n0 B 3.90526f
.ends

