* NGSPICE file created from diff_pair_sample_1074.ext - technology: sky130A

.subckt diff_pair_sample_1074 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X1 VDD2.t9 VN.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X2 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X3 VTAIL.t17 VP.t1 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X4 VDD2.t7 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=1.57245 ps=9.86 w=9.53 l=3.8
X5 VDD2.t6 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=1.57245 ps=9.86 w=9.53 l=3.8
X6 VDD1.t2 VP.t2 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X7 VDD1.t8 VP.t3 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X8 VDD1.t4 VP.t4 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=1.57245 ps=9.86 w=9.53 l=3.8
X9 VTAIL.t5 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X10 VDD1.t7 VP.t5 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=3.7167 ps=19.84 w=9.53 l=3.8
X11 VTAIL.t12 VP.t6 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X12 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=0 ps=0 w=9.53 l=3.8
X13 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=0 ps=0 w=9.53 l=3.8
X14 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=0 ps=0 w=9.53 l=3.8
X15 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=3.7167 ps=19.84 w=9.53 l=3.8
X16 VTAIL.t11 VP.t7 VDD1.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X17 VTAIL.t6 VN.t6 VDD2.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X18 VDD1.t9 VP.t8 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=3.7167 ps=19.84 w=9.53 l=3.8
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=0 ps=0 w=9.53 l=3.8
X20 VDD2.t2 VN.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=3.7167 ps=19.84 w=9.53 l=3.8
X21 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X22 VTAIL.t19 VN.t9 VDD2.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=1.57245 pd=9.86 as=1.57245 ps=9.86 w=9.53 l=3.8
X23 VDD1.t3 VP.t9 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7167 pd=19.84 as=1.57245 ps=9.86 w=9.53 l=3.8
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n31 VP.t4 92.6443
R60 VP.n75 VP.n74 89.5781
R61 VP.n130 VP.n0 89.5781
R62 VP.n73 VP.n18 89.5781
R63 VP.n75 VP.t9 60.4408
R64 VP.n89 VP.t1 60.4408
R65 VP.n102 VP.t2 60.4408
R66 VP.n115 VP.t7 60.4408
R67 VP.n0 VP.t8 60.4408
R68 VP.n18 VP.t5 60.4408
R69 VP.n58 VP.t0 60.4408
R70 VP.n45 VP.t3 60.4408
R71 VP.n32 VP.t6 60.4408
R72 VP.n74 VP.n73 57.7834
R73 VP.n96 VP.n95 56.5193
R74 VP.n109 VP.n108 56.5193
R75 VP.n52 VP.n51 56.5193
R76 VP.n39 VP.n38 56.5193
R77 VP.n32 VP.n31 56.4597
R78 VP.n83 VP.n82 45.8354
R79 VP.n122 VP.n121 45.8354
R80 VP.n65 VP.n64 45.8354
R81 VP.n82 VP.n81 35.1514
R82 VP.n122 VP.n2 35.1514
R83 VP.n65 VP.n20 35.1514
R84 VP.n77 VP.n76 24.4675
R85 VP.n77 VP.n16 24.4675
R86 VP.n81 VP.n16 24.4675
R87 VP.n83 VP.n14 24.4675
R88 VP.n87 VP.n14 24.4675
R89 VP.n88 VP.n87 24.4675
R90 VP.n90 VP.n12 24.4675
R91 VP.n94 VP.n12 24.4675
R92 VP.n95 VP.n94 24.4675
R93 VP.n96 VP.n10 24.4675
R94 VP.n100 VP.n10 24.4675
R95 VP.n101 VP.n100 24.4675
R96 VP.n103 VP.n8 24.4675
R97 VP.n107 VP.n8 24.4675
R98 VP.n108 VP.n107 24.4675
R99 VP.n109 VP.n6 24.4675
R100 VP.n113 VP.n6 24.4675
R101 VP.n114 VP.n113 24.4675
R102 VP.n116 VP.n4 24.4675
R103 VP.n120 VP.n4 24.4675
R104 VP.n121 VP.n120 24.4675
R105 VP.n126 VP.n2 24.4675
R106 VP.n127 VP.n126 24.4675
R107 VP.n128 VP.n127 24.4675
R108 VP.n69 VP.n20 24.4675
R109 VP.n70 VP.n69 24.4675
R110 VP.n71 VP.n70 24.4675
R111 VP.n52 VP.n24 24.4675
R112 VP.n56 VP.n24 24.4675
R113 VP.n57 VP.n56 24.4675
R114 VP.n59 VP.n22 24.4675
R115 VP.n63 VP.n22 24.4675
R116 VP.n64 VP.n63 24.4675
R117 VP.n39 VP.n28 24.4675
R118 VP.n43 VP.n28 24.4675
R119 VP.n44 VP.n43 24.4675
R120 VP.n46 VP.n26 24.4675
R121 VP.n50 VP.n26 24.4675
R122 VP.n51 VP.n50 24.4675
R123 VP.n33 VP.n30 24.4675
R124 VP.n37 VP.n30 24.4675
R125 VP.n38 VP.n37 24.4675
R126 VP.n90 VP.n89 18.5954
R127 VP.n115 VP.n114 18.5954
R128 VP.n58 VP.n57 18.5954
R129 VP.n33 VP.n32 18.5954
R130 VP.n102 VP.n101 12.234
R131 VP.n103 VP.n102 12.234
R132 VP.n45 VP.n44 12.234
R133 VP.n46 VP.n45 12.234
R134 VP.n89 VP.n88 5.87258
R135 VP.n116 VP.n115 5.87258
R136 VP.n59 VP.n58 5.87258
R137 VP.n34 VP.n31 2.51719
R138 VP.n76 VP.n75 0.48984
R139 VP.n128 VP.n0 0.48984
R140 VP.n71 VP.n18 0.48984
R141 VP.n73 VP.n72 0.354971
R142 VP.n74 VP.n17 0.354971
R143 VP.n130 VP.n129 0.354971
R144 VP VP.n130 0.26696
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VDD1.n1 VDD1.t4 67.0925
R203 VDD1.n3 VDD1.t3 67.0924
R204 VDD1.n5 VDD1.n4 64.0692
R205 VDD1.n1 VDD1.n0 61.4545
R206 VDD1.n7 VDD1.n6 61.4544
R207 VDD1.n3 VDD1.n2 61.4543
R208 VDD1.n7 VDD1.n5 51.2056
R209 VDD1 VDD1.n7 2.61257
R210 VDD1.n6 VDD1.t5 2.07815
R211 VDD1.n6 VDD1.t7 2.07815
R212 VDD1.n0 VDD1.t6 2.07815
R213 VDD1.n0 VDD1.t8 2.07815
R214 VDD1.n4 VDD1.t1 2.07815
R215 VDD1.n4 VDD1.t9 2.07815
R216 VDD1.n2 VDD1.t0 2.07815
R217 VDD1.n2 VDD1.t2 2.07815
R218 VDD1 VDD1.n1 0.948776
R219 VDD1.n5 VDD1.n3 0.83524
R220 VTAIL.n11 VTAIL.t4 46.8533
R221 VTAIL.n17 VTAIL.t0 46.8532
R222 VTAIL.n2 VTAIL.t10 46.8532
R223 VTAIL.n16 VTAIL.t13 46.8532
R224 VTAIL.n15 VTAIL.n14 44.7758
R225 VTAIL.n13 VTAIL.n12 44.7758
R226 VTAIL.n10 VTAIL.n9 44.7758
R227 VTAIL.n8 VTAIL.n7 44.7758
R228 VTAIL.n19 VTAIL.n18 44.7755
R229 VTAIL.n1 VTAIL.n0 44.7755
R230 VTAIL.n4 VTAIL.n3 44.7755
R231 VTAIL.n6 VTAIL.n5 44.7755
R232 VTAIL.n8 VTAIL.n6 27.7031
R233 VTAIL.n17 VTAIL.n16 24.1427
R234 VTAIL.n10 VTAIL.n8 3.56084
R235 VTAIL.n11 VTAIL.n10 3.56084
R236 VTAIL.n15 VTAIL.n13 3.56084
R237 VTAIL.n16 VTAIL.n15 3.56084
R238 VTAIL.n6 VTAIL.n4 3.56084
R239 VTAIL.n4 VTAIL.n2 3.56084
R240 VTAIL.n19 VTAIL.n17 3.56084
R241 VTAIL VTAIL.n1 2.72895
R242 VTAIL.n13 VTAIL.n11 2.2505
R243 VTAIL.n2 VTAIL.n1 2.2505
R244 VTAIL.n18 VTAIL.t3 2.07815
R245 VTAIL.n18 VTAIL.t6 2.07815
R246 VTAIL.n0 VTAIL.t1 2.07815
R247 VTAIL.n0 VTAIL.t8 2.07815
R248 VTAIL.n3 VTAIL.t16 2.07815
R249 VTAIL.n3 VTAIL.t11 2.07815
R250 VTAIL.n5 VTAIL.t9 2.07815
R251 VTAIL.n5 VTAIL.t17 2.07815
R252 VTAIL.n14 VTAIL.t15 2.07815
R253 VTAIL.n14 VTAIL.t18 2.07815
R254 VTAIL.n12 VTAIL.t14 2.07815
R255 VTAIL.n12 VTAIL.t12 2.07815
R256 VTAIL.n9 VTAIL.t7 2.07815
R257 VTAIL.n9 VTAIL.t19 2.07815
R258 VTAIL.n7 VTAIL.t2 2.07815
R259 VTAIL.n7 VTAIL.t5 2.07815
R260 VTAIL VTAIL.n19 0.832397
R261 B.n1051 B.n1050 585
R262 B.n344 B.n185 585
R263 B.n343 B.n342 585
R264 B.n341 B.n340 585
R265 B.n339 B.n338 585
R266 B.n337 B.n336 585
R267 B.n335 B.n334 585
R268 B.n333 B.n332 585
R269 B.n331 B.n330 585
R270 B.n329 B.n328 585
R271 B.n327 B.n326 585
R272 B.n325 B.n324 585
R273 B.n323 B.n322 585
R274 B.n321 B.n320 585
R275 B.n319 B.n318 585
R276 B.n317 B.n316 585
R277 B.n315 B.n314 585
R278 B.n313 B.n312 585
R279 B.n311 B.n310 585
R280 B.n309 B.n308 585
R281 B.n307 B.n306 585
R282 B.n305 B.n304 585
R283 B.n303 B.n302 585
R284 B.n301 B.n300 585
R285 B.n299 B.n298 585
R286 B.n297 B.n296 585
R287 B.n295 B.n294 585
R288 B.n293 B.n292 585
R289 B.n291 B.n290 585
R290 B.n289 B.n288 585
R291 B.n287 B.n286 585
R292 B.n285 B.n284 585
R293 B.n283 B.n282 585
R294 B.n281 B.n280 585
R295 B.n279 B.n278 585
R296 B.n277 B.n276 585
R297 B.n275 B.n274 585
R298 B.n273 B.n272 585
R299 B.n271 B.n270 585
R300 B.n269 B.n268 585
R301 B.n267 B.n266 585
R302 B.n265 B.n264 585
R303 B.n263 B.n262 585
R304 B.n261 B.n260 585
R305 B.n259 B.n258 585
R306 B.n257 B.n256 585
R307 B.n255 B.n254 585
R308 B.n253 B.n252 585
R309 B.n251 B.n250 585
R310 B.n249 B.n248 585
R311 B.n247 B.n246 585
R312 B.n245 B.n244 585
R313 B.n243 B.n242 585
R314 B.n241 B.n240 585
R315 B.n239 B.n238 585
R316 B.n237 B.n236 585
R317 B.n235 B.n234 585
R318 B.n233 B.n232 585
R319 B.n231 B.n230 585
R320 B.n229 B.n228 585
R321 B.n227 B.n226 585
R322 B.n225 B.n224 585
R323 B.n223 B.n222 585
R324 B.n221 B.n220 585
R325 B.n219 B.n218 585
R326 B.n217 B.n216 585
R327 B.n215 B.n214 585
R328 B.n213 B.n212 585
R329 B.n211 B.n210 585
R330 B.n209 B.n208 585
R331 B.n207 B.n206 585
R332 B.n205 B.n204 585
R333 B.n203 B.n202 585
R334 B.n201 B.n200 585
R335 B.n199 B.n198 585
R336 B.n197 B.n196 585
R337 B.n195 B.n194 585
R338 B.n193 B.n192 585
R339 B.n1049 B.n146 585
R340 B.n1054 B.n146 585
R341 B.n1048 B.n145 585
R342 B.n1055 B.n145 585
R343 B.n1047 B.n1046 585
R344 B.n1046 B.n141 585
R345 B.n1045 B.n140 585
R346 B.n1061 B.n140 585
R347 B.n1044 B.n139 585
R348 B.n1062 B.n139 585
R349 B.n1043 B.n138 585
R350 B.n1063 B.n138 585
R351 B.n1042 B.n1041 585
R352 B.n1041 B.n134 585
R353 B.n1040 B.n133 585
R354 B.n1069 B.n133 585
R355 B.n1039 B.n132 585
R356 B.n1070 B.n132 585
R357 B.n1038 B.n131 585
R358 B.n1071 B.n131 585
R359 B.n1037 B.n1036 585
R360 B.n1036 B.n127 585
R361 B.n1035 B.n126 585
R362 B.n1077 B.n126 585
R363 B.n1034 B.n125 585
R364 B.n1078 B.n125 585
R365 B.n1033 B.n124 585
R366 B.n1079 B.n124 585
R367 B.n1032 B.n1031 585
R368 B.n1031 B.n120 585
R369 B.n1030 B.n119 585
R370 B.n1085 B.n119 585
R371 B.n1029 B.n118 585
R372 B.n1086 B.n118 585
R373 B.n1028 B.n117 585
R374 B.n1087 B.n117 585
R375 B.n1027 B.n1026 585
R376 B.n1026 B.n113 585
R377 B.n1025 B.n112 585
R378 B.n1093 B.n112 585
R379 B.n1024 B.n111 585
R380 B.n1094 B.n111 585
R381 B.n1023 B.n110 585
R382 B.n1095 B.n110 585
R383 B.n1022 B.n1021 585
R384 B.n1021 B.n106 585
R385 B.n1020 B.n105 585
R386 B.n1101 B.n105 585
R387 B.n1019 B.n104 585
R388 B.n1102 B.n104 585
R389 B.n1018 B.n103 585
R390 B.n1103 B.n103 585
R391 B.n1017 B.n1016 585
R392 B.n1016 B.n99 585
R393 B.n1015 B.n98 585
R394 B.n1109 B.n98 585
R395 B.n1014 B.n97 585
R396 B.n1110 B.n97 585
R397 B.n1013 B.n96 585
R398 B.n1111 B.n96 585
R399 B.n1012 B.n1011 585
R400 B.n1011 B.n92 585
R401 B.n1010 B.n91 585
R402 B.n1117 B.n91 585
R403 B.n1009 B.n90 585
R404 B.n1118 B.n90 585
R405 B.n1008 B.n89 585
R406 B.n1119 B.n89 585
R407 B.n1007 B.n1006 585
R408 B.n1006 B.n85 585
R409 B.n1005 B.n84 585
R410 B.n1125 B.n84 585
R411 B.n1004 B.n83 585
R412 B.n1126 B.n83 585
R413 B.n1003 B.n82 585
R414 B.n1127 B.n82 585
R415 B.n1002 B.n1001 585
R416 B.n1001 B.n78 585
R417 B.n1000 B.n77 585
R418 B.n1133 B.n77 585
R419 B.n999 B.n76 585
R420 B.n1134 B.n76 585
R421 B.n998 B.n75 585
R422 B.n1135 B.n75 585
R423 B.n997 B.n996 585
R424 B.n996 B.n71 585
R425 B.n995 B.n70 585
R426 B.n1141 B.n70 585
R427 B.n994 B.n69 585
R428 B.n1142 B.n69 585
R429 B.n993 B.n68 585
R430 B.n1143 B.n68 585
R431 B.n992 B.n991 585
R432 B.n991 B.n64 585
R433 B.n990 B.n63 585
R434 B.n1149 B.n63 585
R435 B.n989 B.n62 585
R436 B.n1150 B.n62 585
R437 B.n988 B.n61 585
R438 B.n1151 B.n61 585
R439 B.n987 B.n986 585
R440 B.n986 B.n57 585
R441 B.n985 B.n56 585
R442 B.n1157 B.n56 585
R443 B.n984 B.n55 585
R444 B.n1158 B.n55 585
R445 B.n983 B.n54 585
R446 B.n1159 B.n54 585
R447 B.n982 B.n981 585
R448 B.n981 B.n50 585
R449 B.n980 B.n49 585
R450 B.n1165 B.n49 585
R451 B.n979 B.n48 585
R452 B.n1166 B.n48 585
R453 B.n978 B.n47 585
R454 B.n1167 B.n47 585
R455 B.n977 B.n976 585
R456 B.n976 B.n43 585
R457 B.n975 B.n42 585
R458 B.n1173 B.n42 585
R459 B.n974 B.n41 585
R460 B.n1174 B.n41 585
R461 B.n973 B.n40 585
R462 B.n1175 B.n40 585
R463 B.n972 B.n971 585
R464 B.n971 B.n36 585
R465 B.n970 B.n35 585
R466 B.n1181 B.n35 585
R467 B.n969 B.n34 585
R468 B.n1182 B.n34 585
R469 B.n968 B.n33 585
R470 B.n1183 B.n33 585
R471 B.n967 B.n966 585
R472 B.n966 B.n29 585
R473 B.n965 B.n28 585
R474 B.n1189 B.n28 585
R475 B.n964 B.n27 585
R476 B.n1190 B.n27 585
R477 B.n963 B.n26 585
R478 B.n1191 B.n26 585
R479 B.n962 B.n961 585
R480 B.n961 B.n22 585
R481 B.n960 B.n21 585
R482 B.n1197 B.n21 585
R483 B.n959 B.n20 585
R484 B.n1198 B.n20 585
R485 B.n958 B.n19 585
R486 B.n1199 B.n19 585
R487 B.n957 B.n956 585
R488 B.n956 B.n15 585
R489 B.n955 B.n14 585
R490 B.n1205 B.n14 585
R491 B.n954 B.n13 585
R492 B.n1206 B.n13 585
R493 B.n953 B.n12 585
R494 B.n1207 B.n12 585
R495 B.n952 B.n951 585
R496 B.n951 B.n8 585
R497 B.n950 B.n7 585
R498 B.n1213 B.n7 585
R499 B.n949 B.n6 585
R500 B.n1214 B.n6 585
R501 B.n948 B.n5 585
R502 B.n1215 B.n5 585
R503 B.n947 B.n946 585
R504 B.n946 B.n4 585
R505 B.n945 B.n345 585
R506 B.n945 B.n944 585
R507 B.n935 B.n346 585
R508 B.n347 B.n346 585
R509 B.n937 B.n936 585
R510 B.n938 B.n937 585
R511 B.n934 B.n352 585
R512 B.n352 B.n351 585
R513 B.n933 B.n932 585
R514 B.n932 B.n931 585
R515 B.n354 B.n353 585
R516 B.n355 B.n354 585
R517 B.n924 B.n923 585
R518 B.n925 B.n924 585
R519 B.n922 B.n360 585
R520 B.n360 B.n359 585
R521 B.n921 B.n920 585
R522 B.n920 B.n919 585
R523 B.n362 B.n361 585
R524 B.n363 B.n362 585
R525 B.n912 B.n911 585
R526 B.n913 B.n912 585
R527 B.n910 B.n368 585
R528 B.n368 B.n367 585
R529 B.n909 B.n908 585
R530 B.n908 B.n907 585
R531 B.n370 B.n369 585
R532 B.n371 B.n370 585
R533 B.n900 B.n899 585
R534 B.n901 B.n900 585
R535 B.n898 B.n376 585
R536 B.n376 B.n375 585
R537 B.n897 B.n896 585
R538 B.n896 B.n895 585
R539 B.n378 B.n377 585
R540 B.n379 B.n378 585
R541 B.n888 B.n887 585
R542 B.n889 B.n888 585
R543 B.n886 B.n384 585
R544 B.n384 B.n383 585
R545 B.n885 B.n884 585
R546 B.n884 B.n883 585
R547 B.n386 B.n385 585
R548 B.n387 B.n386 585
R549 B.n876 B.n875 585
R550 B.n877 B.n876 585
R551 B.n874 B.n392 585
R552 B.n392 B.n391 585
R553 B.n873 B.n872 585
R554 B.n872 B.n871 585
R555 B.n394 B.n393 585
R556 B.n395 B.n394 585
R557 B.n864 B.n863 585
R558 B.n865 B.n864 585
R559 B.n862 B.n400 585
R560 B.n400 B.n399 585
R561 B.n861 B.n860 585
R562 B.n860 B.n859 585
R563 B.n402 B.n401 585
R564 B.n403 B.n402 585
R565 B.n852 B.n851 585
R566 B.n853 B.n852 585
R567 B.n850 B.n408 585
R568 B.n408 B.n407 585
R569 B.n849 B.n848 585
R570 B.n848 B.n847 585
R571 B.n410 B.n409 585
R572 B.n411 B.n410 585
R573 B.n840 B.n839 585
R574 B.n841 B.n840 585
R575 B.n838 B.n416 585
R576 B.n416 B.n415 585
R577 B.n837 B.n836 585
R578 B.n836 B.n835 585
R579 B.n418 B.n417 585
R580 B.n419 B.n418 585
R581 B.n828 B.n827 585
R582 B.n829 B.n828 585
R583 B.n826 B.n424 585
R584 B.n424 B.n423 585
R585 B.n825 B.n824 585
R586 B.n824 B.n823 585
R587 B.n426 B.n425 585
R588 B.n427 B.n426 585
R589 B.n816 B.n815 585
R590 B.n817 B.n816 585
R591 B.n814 B.n431 585
R592 B.n435 B.n431 585
R593 B.n813 B.n812 585
R594 B.n812 B.n811 585
R595 B.n433 B.n432 585
R596 B.n434 B.n433 585
R597 B.n804 B.n803 585
R598 B.n805 B.n804 585
R599 B.n802 B.n440 585
R600 B.n440 B.n439 585
R601 B.n801 B.n800 585
R602 B.n800 B.n799 585
R603 B.n442 B.n441 585
R604 B.n443 B.n442 585
R605 B.n792 B.n791 585
R606 B.n793 B.n792 585
R607 B.n790 B.n448 585
R608 B.n448 B.n447 585
R609 B.n789 B.n788 585
R610 B.n788 B.n787 585
R611 B.n450 B.n449 585
R612 B.n451 B.n450 585
R613 B.n780 B.n779 585
R614 B.n781 B.n780 585
R615 B.n778 B.n455 585
R616 B.n459 B.n455 585
R617 B.n777 B.n776 585
R618 B.n776 B.n775 585
R619 B.n457 B.n456 585
R620 B.n458 B.n457 585
R621 B.n768 B.n767 585
R622 B.n769 B.n768 585
R623 B.n766 B.n464 585
R624 B.n464 B.n463 585
R625 B.n765 B.n764 585
R626 B.n764 B.n763 585
R627 B.n466 B.n465 585
R628 B.n467 B.n466 585
R629 B.n756 B.n755 585
R630 B.n757 B.n756 585
R631 B.n754 B.n472 585
R632 B.n472 B.n471 585
R633 B.n753 B.n752 585
R634 B.n752 B.n751 585
R635 B.n474 B.n473 585
R636 B.n475 B.n474 585
R637 B.n744 B.n743 585
R638 B.n745 B.n744 585
R639 B.n742 B.n480 585
R640 B.n480 B.n479 585
R641 B.n741 B.n740 585
R642 B.n740 B.n739 585
R643 B.n482 B.n481 585
R644 B.n483 B.n482 585
R645 B.n732 B.n731 585
R646 B.n733 B.n732 585
R647 B.n730 B.n488 585
R648 B.n488 B.n487 585
R649 B.n729 B.n728 585
R650 B.n728 B.n727 585
R651 B.n490 B.n489 585
R652 B.n491 B.n490 585
R653 B.n720 B.n719 585
R654 B.n721 B.n720 585
R655 B.n718 B.n496 585
R656 B.n496 B.n495 585
R657 B.n717 B.n716 585
R658 B.n716 B.n715 585
R659 B.n498 B.n497 585
R660 B.n499 B.n498 585
R661 B.n708 B.n707 585
R662 B.n709 B.n708 585
R663 B.n706 B.n504 585
R664 B.n504 B.n503 585
R665 B.n701 B.n700 585
R666 B.n699 B.n545 585
R667 B.n698 B.n544 585
R668 B.n703 B.n544 585
R669 B.n697 B.n696 585
R670 B.n695 B.n694 585
R671 B.n693 B.n692 585
R672 B.n691 B.n690 585
R673 B.n689 B.n688 585
R674 B.n687 B.n686 585
R675 B.n685 B.n684 585
R676 B.n683 B.n682 585
R677 B.n681 B.n680 585
R678 B.n679 B.n678 585
R679 B.n677 B.n676 585
R680 B.n675 B.n674 585
R681 B.n673 B.n672 585
R682 B.n671 B.n670 585
R683 B.n669 B.n668 585
R684 B.n667 B.n666 585
R685 B.n665 B.n664 585
R686 B.n663 B.n662 585
R687 B.n661 B.n660 585
R688 B.n659 B.n658 585
R689 B.n657 B.n656 585
R690 B.n655 B.n654 585
R691 B.n653 B.n652 585
R692 B.n651 B.n650 585
R693 B.n649 B.n648 585
R694 B.n647 B.n646 585
R695 B.n645 B.n644 585
R696 B.n643 B.n642 585
R697 B.n641 B.n640 585
R698 B.n639 B.n638 585
R699 B.n637 B.n636 585
R700 B.n634 B.n633 585
R701 B.n632 B.n631 585
R702 B.n630 B.n629 585
R703 B.n628 B.n627 585
R704 B.n626 B.n625 585
R705 B.n624 B.n623 585
R706 B.n622 B.n621 585
R707 B.n620 B.n619 585
R708 B.n618 B.n617 585
R709 B.n616 B.n615 585
R710 B.n613 B.n612 585
R711 B.n611 B.n610 585
R712 B.n609 B.n608 585
R713 B.n607 B.n606 585
R714 B.n605 B.n604 585
R715 B.n603 B.n602 585
R716 B.n601 B.n600 585
R717 B.n599 B.n598 585
R718 B.n597 B.n596 585
R719 B.n595 B.n594 585
R720 B.n593 B.n592 585
R721 B.n591 B.n590 585
R722 B.n589 B.n588 585
R723 B.n587 B.n586 585
R724 B.n585 B.n584 585
R725 B.n583 B.n582 585
R726 B.n581 B.n580 585
R727 B.n579 B.n578 585
R728 B.n577 B.n576 585
R729 B.n575 B.n574 585
R730 B.n573 B.n572 585
R731 B.n571 B.n570 585
R732 B.n569 B.n568 585
R733 B.n567 B.n566 585
R734 B.n565 B.n564 585
R735 B.n563 B.n562 585
R736 B.n561 B.n560 585
R737 B.n559 B.n558 585
R738 B.n557 B.n556 585
R739 B.n555 B.n554 585
R740 B.n553 B.n552 585
R741 B.n551 B.n550 585
R742 B.n506 B.n505 585
R743 B.n705 B.n704 585
R744 B.n704 B.n703 585
R745 B.n502 B.n501 585
R746 B.n503 B.n502 585
R747 B.n711 B.n710 585
R748 B.n710 B.n709 585
R749 B.n712 B.n500 585
R750 B.n500 B.n499 585
R751 B.n714 B.n713 585
R752 B.n715 B.n714 585
R753 B.n494 B.n493 585
R754 B.n495 B.n494 585
R755 B.n723 B.n722 585
R756 B.n722 B.n721 585
R757 B.n724 B.n492 585
R758 B.n492 B.n491 585
R759 B.n726 B.n725 585
R760 B.n727 B.n726 585
R761 B.n486 B.n485 585
R762 B.n487 B.n486 585
R763 B.n735 B.n734 585
R764 B.n734 B.n733 585
R765 B.n736 B.n484 585
R766 B.n484 B.n483 585
R767 B.n738 B.n737 585
R768 B.n739 B.n738 585
R769 B.n478 B.n477 585
R770 B.n479 B.n478 585
R771 B.n747 B.n746 585
R772 B.n746 B.n745 585
R773 B.n748 B.n476 585
R774 B.n476 B.n475 585
R775 B.n750 B.n749 585
R776 B.n751 B.n750 585
R777 B.n470 B.n469 585
R778 B.n471 B.n470 585
R779 B.n759 B.n758 585
R780 B.n758 B.n757 585
R781 B.n760 B.n468 585
R782 B.n468 B.n467 585
R783 B.n762 B.n761 585
R784 B.n763 B.n762 585
R785 B.n462 B.n461 585
R786 B.n463 B.n462 585
R787 B.n771 B.n770 585
R788 B.n770 B.n769 585
R789 B.n772 B.n460 585
R790 B.n460 B.n458 585
R791 B.n774 B.n773 585
R792 B.n775 B.n774 585
R793 B.n454 B.n453 585
R794 B.n459 B.n454 585
R795 B.n783 B.n782 585
R796 B.n782 B.n781 585
R797 B.n784 B.n452 585
R798 B.n452 B.n451 585
R799 B.n786 B.n785 585
R800 B.n787 B.n786 585
R801 B.n446 B.n445 585
R802 B.n447 B.n446 585
R803 B.n795 B.n794 585
R804 B.n794 B.n793 585
R805 B.n796 B.n444 585
R806 B.n444 B.n443 585
R807 B.n798 B.n797 585
R808 B.n799 B.n798 585
R809 B.n438 B.n437 585
R810 B.n439 B.n438 585
R811 B.n807 B.n806 585
R812 B.n806 B.n805 585
R813 B.n808 B.n436 585
R814 B.n436 B.n434 585
R815 B.n810 B.n809 585
R816 B.n811 B.n810 585
R817 B.n430 B.n429 585
R818 B.n435 B.n430 585
R819 B.n819 B.n818 585
R820 B.n818 B.n817 585
R821 B.n820 B.n428 585
R822 B.n428 B.n427 585
R823 B.n822 B.n821 585
R824 B.n823 B.n822 585
R825 B.n422 B.n421 585
R826 B.n423 B.n422 585
R827 B.n831 B.n830 585
R828 B.n830 B.n829 585
R829 B.n832 B.n420 585
R830 B.n420 B.n419 585
R831 B.n834 B.n833 585
R832 B.n835 B.n834 585
R833 B.n414 B.n413 585
R834 B.n415 B.n414 585
R835 B.n843 B.n842 585
R836 B.n842 B.n841 585
R837 B.n844 B.n412 585
R838 B.n412 B.n411 585
R839 B.n846 B.n845 585
R840 B.n847 B.n846 585
R841 B.n406 B.n405 585
R842 B.n407 B.n406 585
R843 B.n855 B.n854 585
R844 B.n854 B.n853 585
R845 B.n856 B.n404 585
R846 B.n404 B.n403 585
R847 B.n858 B.n857 585
R848 B.n859 B.n858 585
R849 B.n398 B.n397 585
R850 B.n399 B.n398 585
R851 B.n867 B.n866 585
R852 B.n866 B.n865 585
R853 B.n868 B.n396 585
R854 B.n396 B.n395 585
R855 B.n870 B.n869 585
R856 B.n871 B.n870 585
R857 B.n390 B.n389 585
R858 B.n391 B.n390 585
R859 B.n879 B.n878 585
R860 B.n878 B.n877 585
R861 B.n880 B.n388 585
R862 B.n388 B.n387 585
R863 B.n882 B.n881 585
R864 B.n883 B.n882 585
R865 B.n382 B.n381 585
R866 B.n383 B.n382 585
R867 B.n891 B.n890 585
R868 B.n890 B.n889 585
R869 B.n892 B.n380 585
R870 B.n380 B.n379 585
R871 B.n894 B.n893 585
R872 B.n895 B.n894 585
R873 B.n374 B.n373 585
R874 B.n375 B.n374 585
R875 B.n903 B.n902 585
R876 B.n902 B.n901 585
R877 B.n904 B.n372 585
R878 B.n372 B.n371 585
R879 B.n906 B.n905 585
R880 B.n907 B.n906 585
R881 B.n366 B.n365 585
R882 B.n367 B.n366 585
R883 B.n915 B.n914 585
R884 B.n914 B.n913 585
R885 B.n916 B.n364 585
R886 B.n364 B.n363 585
R887 B.n918 B.n917 585
R888 B.n919 B.n918 585
R889 B.n358 B.n357 585
R890 B.n359 B.n358 585
R891 B.n927 B.n926 585
R892 B.n926 B.n925 585
R893 B.n928 B.n356 585
R894 B.n356 B.n355 585
R895 B.n930 B.n929 585
R896 B.n931 B.n930 585
R897 B.n350 B.n349 585
R898 B.n351 B.n350 585
R899 B.n940 B.n939 585
R900 B.n939 B.n938 585
R901 B.n941 B.n348 585
R902 B.n348 B.n347 585
R903 B.n943 B.n942 585
R904 B.n944 B.n943 585
R905 B.n2 B.n0 585
R906 B.n4 B.n2 585
R907 B.n3 B.n1 585
R908 B.n1214 B.n3 585
R909 B.n1212 B.n1211 585
R910 B.n1213 B.n1212 585
R911 B.n1210 B.n9 585
R912 B.n9 B.n8 585
R913 B.n1209 B.n1208 585
R914 B.n1208 B.n1207 585
R915 B.n11 B.n10 585
R916 B.n1206 B.n11 585
R917 B.n1204 B.n1203 585
R918 B.n1205 B.n1204 585
R919 B.n1202 B.n16 585
R920 B.n16 B.n15 585
R921 B.n1201 B.n1200 585
R922 B.n1200 B.n1199 585
R923 B.n18 B.n17 585
R924 B.n1198 B.n18 585
R925 B.n1196 B.n1195 585
R926 B.n1197 B.n1196 585
R927 B.n1194 B.n23 585
R928 B.n23 B.n22 585
R929 B.n1193 B.n1192 585
R930 B.n1192 B.n1191 585
R931 B.n25 B.n24 585
R932 B.n1190 B.n25 585
R933 B.n1188 B.n1187 585
R934 B.n1189 B.n1188 585
R935 B.n1186 B.n30 585
R936 B.n30 B.n29 585
R937 B.n1185 B.n1184 585
R938 B.n1184 B.n1183 585
R939 B.n32 B.n31 585
R940 B.n1182 B.n32 585
R941 B.n1180 B.n1179 585
R942 B.n1181 B.n1180 585
R943 B.n1178 B.n37 585
R944 B.n37 B.n36 585
R945 B.n1177 B.n1176 585
R946 B.n1176 B.n1175 585
R947 B.n39 B.n38 585
R948 B.n1174 B.n39 585
R949 B.n1172 B.n1171 585
R950 B.n1173 B.n1172 585
R951 B.n1170 B.n44 585
R952 B.n44 B.n43 585
R953 B.n1169 B.n1168 585
R954 B.n1168 B.n1167 585
R955 B.n46 B.n45 585
R956 B.n1166 B.n46 585
R957 B.n1164 B.n1163 585
R958 B.n1165 B.n1164 585
R959 B.n1162 B.n51 585
R960 B.n51 B.n50 585
R961 B.n1161 B.n1160 585
R962 B.n1160 B.n1159 585
R963 B.n53 B.n52 585
R964 B.n1158 B.n53 585
R965 B.n1156 B.n1155 585
R966 B.n1157 B.n1156 585
R967 B.n1154 B.n58 585
R968 B.n58 B.n57 585
R969 B.n1153 B.n1152 585
R970 B.n1152 B.n1151 585
R971 B.n60 B.n59 585
R972 B.n1150 B.n60 585
R973 B.n1148 B.n1147 585
R974 B.n1149 B.n1148 585
R975 B.n1146 B.n65 585
R976 B.n65 B.n64 585
R977 B.n1145 B.n1144 585
R978 B.n1144 B.n1143 585
R979 B.n67 B.n66 585
R980 B.n1142 B.n67 585
R981 B.n1140 B.n1139 585
R982 B.n1141 B.n1140 585
R983 B.n1138 B.n72 585
R984 B.n72 B.n71 585
R985 B.n1137 B.n1136 585
R986 B.n1136 B.n1135 585
R987 B.n74 B.n73 585
R988 B.n1134 B.n74 585
R989 B.n1132 B.n1131 585
R990 B.n1133 B.n1132 585
R991 B.n1130 B.n79 585
R992 B.n79 B.n78 585
R993 B.n1129 B.n1128 585
R994 B.n1128 B.n1127 585
R995 B.n81 B.n80 585
R996 B.n1126 B.n81 585
R997 B.n1124 B.n1123 585
R998 B.n1125 B.n1124 585
R999 B.n1122 B.n86 585
R1000 B.n86 B.n85 585
R1001 B.n1121 B.n1120 585
R1002 B.n1120 B.n1119 585
R1003 B.n88 B.n87 585
R1004 B.n1118 B.n88 585
R1005 B.n1116 B.n1115 585
R1006 B.n1117 B.n1116 585
R1007 B.n1114 B.n93 585
R1008 B.n93 B.n92 585
R1009 B.n1113 B.n1112 585
R1010 B.n1112 B.n1111 585
R1011 B.n95 B.n94 585
R1012 B.n1110 B.n95 585
R1013 B.n1108 B.n1107 585
R1014 B.n1109 B.n1108 585
R1015 B.n1106 B.n100 585
R1016 B.n100 B.n99 585
R1017 B.n1105 B.n1104 585
R1018 B.n1104 B.n1103 585
R1019 B.n102 B.n101 585
R1020 B.n1102 B.n102 585
R1021 B.n1100 B.n1099 585
R1022 B.n1101 B.n1100 585
R1023 B.n1098 B.n107 585
R1024 B.n107 B.n106 585
R1025 B.n1097 B.n1096 585
R1026 B.n1096 B.n1095 585
R1027 B.n109 B.n108 585
R1028 B.n1094 B.n109 585
R1029 B.n1092 B.n1091 585
R1030 B.n1093 B.n1092 585
R1031 B.n1090 B.n114 585
R1032 B.n114 B.n113 585
R1033 B.n1089 B.n1088 585
R1034 B.n1088 B.n1087 585
R1035 B.n116 B.n115 585
R1036 B.n1086 B.n116 585
R1037 B.n1084 B.n1083 585
R1038 B.n1085 B.n1084 585
R1039 B.n1082 B.n121 585
R1040 B.n121 B.n120 585
R1041 B.n1081 B.n1080 585
R1042 B.n1080 B.n1079 585
R1043 B.n123 B.n122 585
R1044 B.n1078 B.n123 585
R1045 B.n1076 B.n1075 585
R1046 B.n1077 B.n1076 585
R1047 B.n1074 B.n128 585
R1048 B.n128 B.n127 585
R1049 B.n1073 B.n1072 585
R1050 B.n1072 B.n1071 585
R1051 B.n130 B.n129 585
R1052 B.n1070 B.n130 585
R1053 B.n1068 B.n1067 585
R1054 B.n1069 B.n1068 585
R1055 B.n1066 B.n135 585
R1056 B.n135 B.n134 585
R1057 B.n1065 B.n1064 585
R1058 B.n1064 B.n1063 585
R1059 B.n137 B.n136 585
R1060 B.n1062 B.n137 585
R1061 B.n1060 B.n1059 585
R1062 B.n1061 B.n1060 585
R1063 B.n1058 B.n142 585
R1064 B.n142 B.n141 585
R1065 B.n1057 B.n1056 585
R1066 B.n1056 B.n1055 585
R1067 B.n144 B.n143 585
R1068 B.n1054 B.n144 585
R1069 B.n1217 B.n1216 585
R1070 B.n1216 B.n1215 585
R1071 B.n701 B.n502 521.33
R1072 B.n192 B.n144 521.33
R1073 B.n704 B.n504 521.33
R1074 B.n1051 B.n146 521.33
R1075 B.n548 B.t14 269.784
R1076 B.n546 B.t18 269.784
R1077 B.n189 B.t10 269.784
R1078 B.n186 B.t21 269.784
R1079 B.n1053 B.n1052 256.663
R1080 B.n1053 B.n184 256.663
R1081 B.n1053 B.n183 256.663
R1082 B.n1053 B.n182 256.663
R1083 B.n1053 B.n181 256.663
R1084 B.n1053 B.n180 256.663
R1085 B.n1053 B.n179 256.663
R1086 B.n1053 B.n178 256.663
R1087 B.n1053 B.n177 256.663
R1088 B.n1053 B.n176 256.663
R1089 B.n1053 B.n175 256.663
R1090 B.n1053 B.n174 256.663
R1091 B.n1053 B.n173 256.663
R1092 B.n1053 B.n172 256.663
R1093 B.n1053 B.n171 256.663
R1094 B.n1053 B.n170 256.663
R1095 B.n1053 B.n169 256.663
R1096 B.n1053 B.n168 256.663
R1097 B.n1053 B.n167 256.663
R1098 B.n1053 B.n166 256.663
R1099 B.n1053 B.n165 256.663
R1100 B.n1053 B.n164 256.663
R1101 B.n1053 B.n163 256.663
R1102 B.n1053 B.n162 256.663
R1103 B.n1053 B.n161 256.663
R1104 B.n1053 B.n160 256.663
R1105 B.n1053 B.n159 256.663
R1106 B.n1053 B.n158 256.663
R1107 B.n1053 B.n157 256.663
R1108 B.n1053 B.n156 256.663
R1109 B.n1053 B.n155 256.663
R1110 B.n1053 B.n154 256.663
R1111 B.n1053 B.n153 256.663
R1112 B.n1053 B.n152 256.663
R1113 B.n1053 B.n151 256.663
R1114 B.n1053 B.n150 256.663
R1115 B.n1053 B.n149 256.663
R1116 B.n1053 B.n148 256.663
R1117 B.n1053 B.n147 256.663
R1118 B.n703 B.n702 256.663
R1119 B.n703 B.n507 256.663
R1120 B.n703 B.n508 256.663
R1121 B.n703 B.n509 256.663
R1122 B.n703 B.n510 256.663
R1123 B.n703 B.n511 256.663
R1124 B.n703 B.n512 256.663
R1125 B.n703 B.n513 256.663
R1126 B.n703 B.n514 256.663
R1127 B.n703 B.n515 256.663
R1128 B.n703 B.n516 256.663
R1129 B.n703 B.n517 256.663
R1130 B.n703 B.n518 256.663
R1131 B.n703 B.n519 256.663
R1132 B.n703 B.n520 256.663
R1133 B.n703 B.n521 256.663
R1134 B.n703 B.n522 256.663
R1135 B.n703 B.n523 256.663
R1136 B.n703 B.n524 256.663
R1137 B.n703 B.n525 256.663
R1138 B.n703 B.n526 256.663
R1139 B.n703 B.n527 256.663
R1140 B.n703 B.n528 256.663
R1141 B.n703 B.n529 256.663
R1142 B.n703 B.n530 256.663
R1143 B.n703 B.n531 256.663
R1144 B.n703 B.n532 256.663
R1145 B.n703 B.n533 256.663
R1146 B.n703 B.n534 256.663
R1147 B.n703 B.n535 256.663
R1148 B.n703 B.n536 256.663
R1149 B.n703 B.n537 256.663
R1150 B.n703 B.n538 256.663
R1151 B.n703 B.n539 256.663
R1152 B.n703 B.n540 256.663
R1153 B.n703 B.n541 256.663
R1154 B.n703 B.n542 256.663
R1155 B.n703 B.n543 256.663
R1156 B.n710 B.n502 163.367
R1157 B.n710 B.n500 163.367
R1158 B.n714 B.n500 163.367
R1159 B.n714 B.n494 163.367
R1160 B.n722 B.n494 163.367
R1161 B.n722 B.n492 163.367
R1162 B.n726 B.n492 163.367
R1163 B.n726 B.n486 163.367
R1164 B.n734 B.n486 163.367
R1165 B.n734 B.n484 163.367
R1166 B.n738 B.n484 163.367
R1167 B.n738 B.n478 163.367
R1168 B.n746 B.n478 163.367
R1169 B.n746 B.n476 163.367
R1170 B.n750 B.n476 163.367
R1171 B.n750 B.n470 163.367
R1172 B.n758 B.n470 163.367
R1173 B.n758 B.n468 163.367
R1174 B.n762 B.n468 163.367
R1175 B.n762 B.n462 163.367
R1176 B.n770 B.n462 163.367
R1177 B.n770 B.n460 163.367
R1178 B.n774 B.n460 163.367
R1179 B.n774 B.n454 163.367
R1180 B.n782 B.n454 163.367
R1181 B.n782 B.n452 163.367
R1182 B.n786 B.n452 163.367
R1183 B.n786 B.n446 163.367
R1184 B.n794 B.n446 163.367
R1185 B.n794 B.n444 163.367
R1186 B.n798 B.n444 163.367
R1187 B.n798 B.n438 163.367
R1188 B.n806 B.n438 163.367
R1189 B.n806 B.n436 163.367
R1190 B.n810 B.n436 163.367
R1191 B.n810 B.n430 163.367
R1192 B.n818 B.n430 163.367
R1193 B.n818 B.n428 163.367
R1194 B.n822 B.n428 163.367
R1195 B.n822 B.n422 163.367
R1196 B.n830 B.n422 163.367
R1197 B.n830 B.n420 163.367
R1198 B.n834 B.n420 163.367
R1199 B.n834 B.n414 163.367
R1200 B.n842 B.n414 163.367
R1201 B.n842 B.n412 163.367
R1202 B.n846 B.n412 163.367
R1203 B.n846 B.n406 163.367
R1204 B.n854 B.n406 163.367
R1205 B.n854 B.n404 163.367
R1206 B.n858 B.n404 163.367
R1207 B.n858 B.n398 163.367
R1208 B.n866 B.n398 163.367
R1209 B.n866 B.n396 163.367
R1210 B.n870 B.n396 163.367
R1211 B.n870 B.n390 163.367
R1212 B.n878 B.n390 163.367
R1213 B.n878 B.n388 163.367
R1214 B.n882 B.n388 163.367
R1215 B.n882 B.n382 163.367
R1216 B.n890 B.n382 163.367
R1217 B.n890 B.n380 163.367
R1218 B.n894 B.n380 163.367
R1219 B.n894 B.n374 163.367
R1220 B.n902 B.n374 163.367
R1221 B.n902 B.n372 163.367
R1222 B.n906 B.n372 163.367
R1223 B.n906 B.n366 163.367
R1224 B.n914 B.n366 163.367
R1225 B.n914 B.n364 163.367
R1226 B.n918 B.n364 163.367
R1227 B.n918 B.n358 163.367
R1228 B.n926 B.n358 163.367
R1229 B.n926 B.n356 163.367
R1230 B.n930 B.n356 163.367
R1231 B.n930 B.n350 163.367
R1232 B.n939 B.n350 163.367
R1233 B.n939 B.n348 163.367
R1234 B.n943 B.n348 163.367
R1235 B.n943 B.n2 163.367
R1236 B.n1216 B.n2 163.367
R1237 B.n1216 B.n3 163.367
R1238 B.n1212 B.n3 163.367
R1239 B.n1212 B.n9 163.367
R1240 B.n1208 B.n9 163.367
R1241 B.n1208 B.n11 163.367
R1242 B.n1204 B.n11 163.367
R1243 B.n1204 B.n16 163.367
R1244 B.n1200 B.n16 163.367
R1245 B.n1200 B.n18 163.367
R1246 B.n1196 B.n18 163.367
R1247 B.n1196 B.n23 163.367
R1248 B.n1192 B.n23 163.367
R1249 B.n1192 B.n25 163.367
R1250 B.n1188 B.n25 163.367
R1251 B.n1188 B.n30 163.367
R1252 B.n1184 B.n30 163.367
R1253 B.n1184 B.n32 163.367
R1254 B.n1180 B.n32 163.367
R1255 B.n1180 B.n37 163.367
R1256 B.n1176 B.n37 163.367
R1257 B.n1176 B.n39 163.367
R1258 B.n1172 B.n39 163.367
R1259 B.n1172 B.n44 163.367
R1260 B.n1168 B.n44 163.367
R1261 B.n1168 B.n46 163.367
R1262 B.n1164 B.n46 163.367
R1263 B.n1164 B.n51 163.367
R1264 B.n1160 B.n51 163.367
R1265 B.n1160 B.n53 163.367
R1266 B.n1156 B.n53 163.367
R1267 B.n1156 B.n58 163.367
R1268 B.n1152 B.n58 163.367
R1269 B.n1152 B.n60 163.367
R1270 B.n1148 B.n60 163.367
R1271 B.n1148 B.n65 163.367
R1272 B.n1144 B.n65 163.367
R1273 B.n1144 B.n67 163.367
R1274 B.n1140 B.n67 163.367
R1275 B.n1140 B.n72 163.367
R1276 B.n1136 B.n72 163.367
R1277 B.n1136 B.n74 163.367
R1278 B.n1132 B.n74 163.367
R1279 B.n1132 B.n79 163.367
R1280 B.n1128 B.n79 163.367
R1281 B.n1128 B.n81 163.367
R1282 B.n1124 B.n81 163.367
R1283 B.n1124 B.n86 163.367
R1284 B.n1120 B.n86 163.367
R1285 B.n1120 B.n88 163.367
R1286 B.n1116 B.n88 163.367
R1287 B.n1116 B.n93 163.367
R1288 B.n1112 B.n93 163.367
R1289 B.n1112 B.n95 163.367
R1290 B.n1108 B.n95 163.367
R1291 B.n1108 B.n100 163.367
R1292 B.n1104 B.n100 163.367
R1293 B.n1104 B.n102 163.367
R1294 B.n1100 B.n102 163.367
R1295 B.n1100 B.n107 163.367
R1296 B.n1096 B.n107 163.367
R1297 B.n1096 B.n109 163.367
R1298 B.n1092 B.n109 163.367
R1299 B.n1092 B.n114 163.367
R1300 B.n1088 B.n114 163.367
R1301 B.n1088 B.n116 163.367
R1302 B.n1084 B.n116 163.367
R1303 B.n1084 B.n121 163.367
R1304 B.n1080 B.n121 163.367
R1305 B.n1080 B.n123 163.367
R1306 B.n1076 B.n123 163.367
R1307 B.n1076 B.n128 163.367
R1308 B.n1072 B.n128 163.367
R1309 B.n1072 B.n130 163.367
R1310 B.n1068 B.n130 163.367
R1311 B.n1068 B.n135 163.367
R1312 B.n1064 B.n135 163.367
R1313 B.n1064 B.n137 163.367
R1314 B.n1060 B.n137 163.367
R1315 B.n1060 B.n142 163.367
R1316 B.n1056 B.n142 163.367
R1317 B.n1056 B.n144 163.367
R1318 B.n545 B.n544 163.367
R1319 B.n696 B.n544 163.367
R1320 B.n694 B.n693 163.367
R1321 B.n690 B.n689 163.367
R1322 B.n686 B.n685 163.367
R1323 B.n682 B.n681 163.367
R1324 B.n678 B.n677 163.367
R1325 B.n674 B.n673 163.367
R1326 B.n670 B.n669 163.367
R1327 B.n666 B.n665 163.367
R1328 B.n662 B.n661 163.367
R1329 B.n658 B.n657 163.367
R1330 B.n654 B.n653 163.367
R1331 B.n650 B.n649 163.367
R1332 B.n646 B.n645 163.367
R1333 B.n642 B.n641 163.367
R1334 B.n638 B.n637 163.367
R1335 B.n633 B.n632 163.367
R1336 B.n629 B.n628 163.367
R1337 B.n625 B.n624 163.367
R1338 B.n621 B.n620 163.367
R1339 B.n617 B.n616 163.367
R1340 B.n612 B.n611 163.367
R1341 B.n608 B.n607 163.367
R1342 B.n604 B.n603 163.367
R1343 B.n600 B.n599 163.367
R1344 B.n596 B.n595 163.367
R1345 B.n592 B.n591 163.367
R1346 B.n588 B.n587 163.367
R1347 B.n584 B.n583 163.367
R1348 B.n580 B.n579 163.367
R1349 B.n576 B.n575 163.367
R1350 B.n572 B.n571 163.367
R1351 B.n568 B.n567 163.367
R1352 B.n564 B.n563 163.367
R1353 B.n560 B.n559 163.367
R1354 B.n556 B.n555 163.367
R1355 B.n552 B.n551 163.367
R1356 B.n704 B.n506 163.367
R1357 B.n708 B.n504 163.367
R1358 B.n708 B.n498 163.367
R1359 B.n716 B.n498 163.367
R1360 B.n716 B.n496 163.367
R1361 B.n720 B.n496 163.367
R1362 B.n720 B.n490 163.367
R1363 B.n728 B.n490 163.367
R1364 B.n728 B.n488 163.367
R1365 B.n732 B.n488 163.367
R1366 B.n732 B.n482 163.367
R1367 B.n740 B.n482 163.367
R1368 B.n740 B.n480 163.367
R1369 B.n744 B.n480 163.367
R1370 B.n744 B.n474 163.367
R1371 B.n752 B.n474 163.367
R1372 B.n752 B.n472 163.367
R1373 B.n756 B.n472 163.367
R1374 B.n756 B.n466 163.367
R1375 B.n764 B.n466 163.367
R1376 B.n764 B.n464 163.367
R1377 B.n768 B.n464 163.367
R1378 B.n768 B.n457 163.367
R1379 B.n776 B.n457 163.367
R1380 B.n776 B.n455 163.367
R1381 B.n780 B.n455 163.367
R1382 B.n780 B.n450 163.367
R1383 B.n788 B.n450 163.367
R1384 B.n788 B.n448 163.367
R1385 B.n792 B.n448 163.367
R1386 B.n792 B.n442 163.367
R1387 B.n800 B.n442 163.367
R1388 B.n800 B.n440 163.367
R1389 B.n804 B.n440 163.367
R1390 B.n804 B.n433 163.367
R1391 B.n812 B.n433 163.367
R1392 B.n812 B.n431 163.367
R1393 B.n816 B.n431 163.367
R1394 B.n816 B.n426 163.367
R1395 B.n824 B.n426 163.367
R1396 B.n824 B.n424 163.367
R1397 B.n828 B.n424 163.367
R1398 B.n828 B.n418 163.367
R1399 B.n836 B.n418 163.367
R1400 B.n836 B.n416 163.367
R1401 B.n840 B.n416 163.367
R1402 B.n840 B.n410 163.367
R1403 B.n848 B.n410 163.367
R1404 B.n848 B.n408 163.367
R1405 B.n852 B.n408 163.367
R1406 B.n852 B.n402 163.367
R1407 B.n860 B.n402 163.367
R1408 B.n860 B.n400 163.367
R1409 B.n864 B.n400 163.367
R1410 B.n864 B.n394 163.367
R1411 B.n872 B.n394 163.367
R1412 B.n872 B.n392 163.367
R1413 B.n876 B.n392 163.367
R1414 B.n876 B.n386 163.367
R1415 B.n884 B.n386 163.367
R1416 B.n884 B.n384 163.367
R1417 B.n888 B.n384 163.367
R1418 B.n888 B.n378 163.367
R1419 B.n896 B.n378 163.367
R1420 B.n896 B.n376 163.367
R1421 B.n900 B.n376 163.367
R1422 B.n900 B.n370 163.367
R1423 B.n908 B.n370 163.367
R1424 B.n908 B.n368 163.367
R1425 B.n912 B.n368 163.367
R1426 B.n912 B.n362 163.367
R1427 B.n920 B.n362 163.367
R1428 B.n920 B.n360 163.367
R1429 B.n924 B.n360 163.367
R1430 B.n924 B.n354 163.367
R1431 B.n932 B.n354 163.367
R1432 B.n932 B.n352 163.367
R1433 B.n937 B.n352 163.367
R1434 B.n937 B.n346 163.367
R1435 B.n945 B.n346 163.367
R1436 B.n946 B.n945 163.367
R1437 B.n946 B.n5 163.367
R1438 B.n6 B.n5 163.367
R1439 B.n7 B.n6 163.367
R1440 B.n951 B.n7 163.367
R1441 B.n951 B.n12 163.367
R1442 B.n13 B.n12 163.367
R1443 B.n14 B.n13 163.367
R1444 B.n956 B.n14 163.367
R1445 B.n956 B.n19 163.367
R1446 B.n20 B.n19 163.367
R1447 B.n21 B.n20 163.367
R1448 B.n961 B.n21 163.367
R1449 B.n961 B.n26 163.367
R1450 B.n27 B.n26 163.367
R1451 B.n28 B.n27 163.367
R1452 B.n966 B.n28 163.367
R1453 B.n966 B.n33 163.367
R1454 B.n34 B.n33 163.367
R1455 B.n35 B.n34 163.367
R1456 B.n971 B.n35 163.367
R1457 B.n971 B.n40 163.367
R1458 B.n41 B.n40 163.367
R1459 B.n42 B.n41 163.367
R1460 B.n976 B.n42 163.367
R1461 B.n976 B.n47 163.367
R1462 B.n48 B.n47 163.367
R1463 B.n49 B.n48 163.367
R1464 B.n981 B.n49 163.367
R1465 B.n981 B.n54 163.367
R1466 B.n55 B.n54 163.367
R1467 B.n56 B.n55 163.367
R1468 B.n986 B.n56 163.367
R1469 B.n986 B.n61 163.367
R1470 B.n62 B.n61 163.367
R1471 B.n63 B.n62 163.367
R1472 B.n991 B.n63 163.367
R1473 B.n991 B.n68 163.367
R1474 B.n69 B.n68 163.367
R1475 B.n70 B.n69 163.367
R1476 B.n996 B.n70 163.367
R1477 B.n996 B.n75 163.367
R1478 B.n76 B.n75 163.367
R1479 B.n77 B.n76 163.367
R1480 B.n1001 B.n77 163.367
R1481 B.n1001 B.n82 163.367
R1482 B.n83 B.n82 163.367
R1483 B.n84 B.n83 163.367
R1484 B.n1006 B.n84 163.367
R1485 B.n1006 B.n89 163.367
R1486 B.n90 B.n89 163.367
R1487 B.n91 B.n90 163.367
R1488 B.n1011 B.n91 163.367
R1489 B.n1011 B.n96 163.367
R1490 B.n97 B.n96 163.367
R1491 B.n98 B.n97 163.367
R1492 B.n1016 B.n98 163.367
R1493 B.n1016 B.n103 163.367
R1494 B.n104 B.n103 163.367
R1495 B.n105 B.n104 163.367
R1496 B.n1021 B.n105 163.367
R1497 B.n1021 B.n110 163.367
R1498 B.n111 B.n110 163.367
R1499 B.n112 B.n111 163.367
R1500 B.n1026 B.n112 163.367
R1501 B.n1026 B.n117 163.367
R1502 B.n118 B.n117 163.367
R1503 B.n119 B.n118 163.367
R1504 B.n1031 B.n119 163.367
R1505 B.n1031 B.n124 163.367
R1506 B.n125 B.n124 163.367
R1507 B.n126 B.n125 163.367
R1508 B.n1036 B.n126 163.367
R1509 B.n1036 B.n131 163.367
R1510 B.n132 B.n131 163.367
R1511 B.n133 B.n132 163.367
R1512 B.n1041 B.n133 163.367
R1513 B.n1041 B.n138 163.367
R1514 B.n139 B.n138 163.367
R1515 B.n140 B.n139 163.367
R1516 B.n1046 B.n140 163.367
R1517 B.n1046 B.n145 163.367
R1518 B.n146 B.n145 163.367
R1519 B.n196 B.n195 163.367
R1520 B.n200 B.n199 163.367
R1521 B.n204 B.n203 163.367
R1522 B.n208 B.n207 163.367
R1523 B.n212 B.n211 163.367
R1524 B.n216 B.n215 163.367
R1525 B.n220 B.n219 163.367
R1526 B.n224 B.n223 163.367
R1527 B.n228 B.n227 163.367
R1528 B.n232 B.n231 163.367
R1529 B.n236 B.n235 163.367
R1530 B.n240 B.n239 163.367
R1531 B.n244 B.n243 163.367
R1532 B.n248 B.n247 163.367
R1533 B.n252 B.n251 163.367
R1534 B.n256 B.n255 163.367
R1535 B.n260 B.n259 163.367
R1536 B.n264 B.n263 163.367
R1537 B.n268 B.n267 163.367
R1538 B.n272 B.n271 163.367
R1539 B.n276 B.n275 163.367
R1540 B.n280 B.n279 163.367
R1541 B.n284 B.n283 163.367
R1542 B.n288 B.n287 163.367
R1543 B.n292 B.n291 163.367
R1544 B.n296 B.n295 163.367
R1545 B.n300 B.n299 163.367
R1546 B.n304 B.n303 163.367
R1547 B.n308 B.n307 163.367
R1548 B.n312 B.n311 163.367
R1549 B.n316 B.n315 163.367
R1550 B.n320 B.n319 163.367
R1551 B.n324 B.n323 163.367
R1552 B.n328 B.n327 163.367
R1553 B.n332 B.n331 163.367
R1554 B.n336 B.n335 163.367
R1555 B.n340 B.n339 163.367
R1556 B.n342 B.n185 163.367
R1557 B.n548 B.t17 148.506
R1558 B.n186 B.t22 148.506
R1559 B.n546 B.t20 148.494
R1560 B.n189 B.t12 148.494
R1561 B.n703 B.n503 91.3885
R1562 B.n1054 B.n1053 91.3885
R1563 B.n549 B.n548 80.0975
R1564 B.n547 B.n546 80.0975
R1565 B.n190 B.n189 80.0975
R1566 B.n187 B.n186 80.0975
R1567 B.n702 B.n701 71.676
R1568 B.n696 B.n507 71.676
R1569 B.n693 B.n508 71.676
R1570 B.n689 B.n509 71.676
R1571 B.n685 B.n510 71.676
R1572 B.n681 B.n511 71.676
R1573 B.n677 B.n512 71.676
R1574 B.n673 B.n513 71.676
R1575 B.n669 B.n514 71.676
R1576 B.n665 B.n515 71.676
R1577 B.n661 B.n516 71.676
R1578 B.n657 B.n517 71.676
R1579 B.n653 B.n518 71.676
R1580 B.n649 B.n519 71.676
R1581 B.n645 B.n520 71.676
R1582 B.n641 B.n521 71.676
R1583 B.n637 B.n522 71.676
R1584 B.n632 B.n523 71.676
R1585 B.n628 B.n524 71.676
R1586 B.n624 B.n525 71.676
R1587 B.n620 B.n526 71.676
R1588 B.n616 B.n527 71.676
R1589 B.n611 B.n528 71.676
R1590 B.n607 B.n529 71.676
R1591 B.n603 B.n530 71.676
R1592 B.n599 B.n531 71.676
R1593 B.n595 B.n532 71.676
R1594 B.n591 B.n533 71.676
R1595 B.n587 B.n534 71.676
R1596 B.n583 B.n535 71.676
R1597 B.n579 B.n536 71.676
R1598 B.n575 B.n537 71.676
R1599 B.n571 B.n538 71.676
R1600 B.n567 B.n539 71.676
R1601 B.n563 B.n540 71.676
R1602 B.n559 B.n541 71.676
R1603 B.n555 B.n542 71.676
R1604 B.n551 B.n543 71.676
R1605 B.n192 B.n147 71.676
R1606 B.n196 B.n148 71.676
R1607 B.n200 B.n149 71.676
R1608 B.n204 B.n150 71.676
R1609 B.n208 B.n151 71.676
R1610 B.n212 B.n152 71.676
R1611 B.n216 B.n153 71.676
R1612 B.n220 B.n154 71.676
R1613 B.n224 B.n155 71.676
R1614 B.n228 B.n156 71.676
R1615 B.n232 B.n157 71.676
R1616 B.n236 B.n158 71.676
R1617 B.n240 B.n159 71.676
R1618 B.n244 B.n160 71.676
R1619 B.n248 B.n161 71.676
R1620 B.n252 B.n162 71.676
R1621 B.n256 B.n163 71.676
R1622 B.n260 B.n164 71.676
R1623 B.n264 B.n165 71.676
R1624 B.n268 B.n166 71.676
R1625 B.n272 B.n167 71.676
R1626 B.n276 B.n168 71.676
R1627 B.n280 B.n169 71.676
R1628 B.n284 B.n170 71.676
R1629 B.n288 B.n171 71.676
R1630 B.n292 B.n172 71.676
R1631 B.n296 B.n173 71.676
R1632 B.n300 B.n174 71.676
R1633 B.n304 B.n175 71.676
R1634 B.n308 B.n176 71.676
R1635 B.n312 B.n177 71.676
R1636 B.n316 B.n178 71.676
R1637 B.n320 B.n179 71.676
R1638 B.n324 B.n180 71.676
R1639 B.n328 B.n181 71.676
R1640 B.n332 B.n182 71.676
R1641 B.n336 B.n183 71.676
R1642 B.n340 B.n184 71.676
R1643 B.n1052 B.n185 71.676
R1644 B.n1052 B.n1051 71.676
R1645 B.n342 B.n184 71.676
R1646 B.n339 B.n183 71.676
R1647 B.n335 B.n182 71.676
R1648 B.n331 B.n181 71.676
R1649 B.n327 B.n180 71.676
R1650 B.n323 B.n179 71.676
R1651 B.n319 B.n178 71.676
R1652 B.n315 B.n177 71.676
R1653 B.n311 B.n176 71.676
R1654 B.n307 B.n175 71.676
R1655 B.n303 B.n174 71.676
R1656 B.n299 B.n173 71.676
R1657 B.n295 B.n172 71.676
R1658 B.n291 B.n171 71.676
R1659 B.n287 B.n170 71.676
R1660 B.n283 B.n169 71.676
R1661 B.n279 B.n168 71.676
R1662 B.n275 B.n167 71.676
R1663 B.n271 B.n166 71.676
R1664 B.n267 B.n165 71.676
R1665 B.n263 B.n164 71.676
R1666 B.n259 B.n163 71.676
R1667 B.n255 B.n162 71.676
R1668 B.n251 B.n161 71.676
R1669 B.n247 B.n160 71.676
R1670 B.n243 B.n159 71.676
R1671 B.n239 B.n158 71.676
R1672 B.n235 B.n157 71.676
R1673 B.n231 B.n156 71.676
R1674 B.n227 B.n155 71.676
R1675 B.n223 B.n154 71.676
R1676 B.n219 B.n153 71.676
R1677 B.n215 B.n152 71.676
R1678 B.n211 B.n151 71.676
R1679 B.n207 B.n150 71.676
R1680 B.n203 B.n149 71.676
R1681 B.n199 B.n148 71.676
R1682 B.n195 B.n147 71.676
R1683 B.n702 B.n545 71.676
R1684 B.n694 B.n507 71.676
R1685 B.n690 B.n508 71.676
R1686 B.n686 B.n509 71.676
R1687 B.n682 B.n510 71.676
R1688 B.n678 B.n511 71.676
R1689 B.n674 B.n512 71.676
R1690 B.n670 B.n513 71.676
R1691 B.n666 B.n514 71.676
R1692 B.n662 B.n515 71.676
R1693 B.n658 B.n516 71.676
R1694 B.n654 B.n517 71.676
R1695 B.n650 B.n518 71.676
R1696 B.n646 B.n519 71.676
R1697 B.n642 B.n520 71.676
R1698 B.n638 B.n521 71.676
R1699 B.n633 B.n522 71.676
R1700 B.n629 B.n523 71.676
R1701 B.n625 B.n524 71.676
R1702 B.n621 B.n525 71.676
R1703 B.n617 B.n526 71.676
R1704 B.n612 B.n527 71.676
R1705 B.n608 B.n528 71.676
R1706 B.n604 B.n529 71.676
R1707 B.n600 B.n530 71.676
R1708 B.n596 B.n531 71.676
R1709 B.n592 B.n532 71.676
R1710 B.n588 B.n533 71.676
R1711 B.n584 B.n534 71.676
R1712 B.n580 B.n535 71.676
R1713 B.n576 B.n536 71.676
R1714 B.n572 B.n537 71.676
R1715 B.n568 B.n538 71.676
R1716 B.n564 B.n539 71.676
R1717 B.n560 B.n540 71.676
R1718 B.n556 B.n541 71.676
R1719 B.n552 B.n542 71.676
R1720 B.n543 B.n506 71.676
R1721 B.n549 B.t16 68.408
R1722 B.n187 B.t23 68.408
R1723 B.n547 B.t19 68.3963
R1724 B.n190 B.t13 68.3963
R1725 B.n614 B.n549 59.5399
R1726 B.n635 B.n547 59.5399
R1727 B.n191 B.n190 59.5399
R1728 B.n188 B.n187 59.5399
R1729 B.n709 B.n503 50.524
R1730 B.n709 B.n499 50.524
R1731 B.n715 B.n499 50.524
R1732 B.n715 B.n495 50.524
R1733 B.n721 B.n495 50.524
R1734 B.n721 B.n491 50.524
R1735 B.n727 B.n491 50.524
R1736 B.n727 B.n487 50.524
R1737 B.n733 B.n487 50.524
R1738 B.n739 B.n483 50.524
R1739 B.n739 B.n479 50.524
R1740 B.n745 B.n479 50.524
R1741 B.n745 B.n475 50.524
R1742 B.n751 B.n475 50.524
R1743 B.n751 B.n471 50.524
R1744 B.n757 B.n471 50.524
R1745 B.n757 B.n467 50.524
R1746 B.n763 B.n467 50.524
R1747 B.n763 B.n463 50.524
R1748 B.n769 B.n463 50.524
R1749 B.n769 B.n458 50.524
R1750 B.n775 B.n458 50.524
R1751 B.n775 B.n459 50.524
R1752 B.n781 B.n451 50.524
R1753 B.n787 B.n451 50.524
R1754 B.n787 B.n447 50.524
R1755 B.n793 B.n447 50.524
R1756 B.n793 B.n443 50.524
R1757 B.n799 B.n443 50.524
R1758 B.n799 B.n439 50.524
R1759 B.n805 B.n439 50.524
R1760 B.n805 B.n434 50.524
R1761 B.n811 B.n434 50.524
R1762 B.n811 B.n435 50.524
R1763 B.n817 B.n427 50.524
R1764 B.n823 B.n427 50.524
R1765 B.n823 B.n423 50.524
R1766 B.n829 B.n423 50.524
R1767 B.n829 B.n419 50.524
R1768 B.n835 B.n419 50.524
R1769 B.n835 B.n415 50.524
R1770 B.n841 B.n415 50.524
R1771 B.n841 B.n411 50.524
R1772 B.n847 B.n411 50.524
R1773 B.n847 B.n407 50.524
R1774 B.n853 B.n407 50.524
R1775 B.n859 B.n403 50.524
R1776 B.n859 B.n399 50.524
R1777 B.n865 B.n399 50.524
R1778 B.n865 B.n395 50.524
R1779 B.n871 B.n395 50.524
R1780 B.n871 B.n391 50.524
R1781 B.n877 B.n391 50.524
R1782 B.n877 B.n387 50.524
R1783 B.n883 B.n387 50.524
R1784 B.n883 B.n383 50.524
R1785 B.n889 B.n383 50.524
R1786 B.n895 B.n379 50.524
R1787 B.n895 B.n375 50.524
R1788 B.n901 B.n375 50.524
R1789 B.n901 B.n371 50.524
R1790 B.n907 B.n371 50.524
R1791 B.n907 B.n367 50.524
R1792 B.n913 B.n367 50.524
R1793 B.n913 B.n363 50.524
R1794 B.n919 B.n363 50.524
R1795 B.n919 B.n359 50.524
R1796 B.n925 B.n359 50.524
R1797 B.n931 B.n355 50.524
R1798 B.n931 B.n351 50.524
R1799 B.n938 B.n351 50.524
R1800 B.n938 B.n347 50.524
R1801 B.n944 B.n347 50.524
R1802 B.n944 B.n4 50.524
R1803 B.n1215 B.n4 50.524
R1804 B.n1215 B.n1214 50.524
R1805 B.n1214 B.n1213 50.524
R1806 B.n1213 B.n8 50.524
R1807 B.n1207 B.n8 50.524
R1808 B.n1207 B.n1206 50.524
R1809 B.n1206 B.n1205 50.524
R1810 B.n1205 B.n15 50.524
R1811 B.n1199 B.n1198 50.524
R1812 B.n1198 B.n1197 50.524
R1813 B.n1197 B.n22 50.524
R1814 B.n1191 B.n22 50.524
R1815 B.n1191 B.n1190 50.524
R1816 B.n1190 B.n1189 50.524
R1817 B.n1189 B.n29 50.524
R1818 B.n1183 B.n29 50.524
R1819 B.n1183 B.n1182 50.524
R1820 B.n1182 B.n1181 50.524
R1821 B.n1181 B.n36 50.524
R1822 B.n1175 B.n1174 50.524
R1823 B.n1174 B.n1173 50.524
R1824 B.n1173 B.n43 50.524
R1825 B.n1167 B.n43 50.524
R1826 B.n1167 B.n1166 50.524
R1827 B.n1166 B.n1165 50.524
R1828 B.n1165 B.n50 50.524
R1829 B.n1159 B.n50 50.524
R1830 B.n1159 B.n1158 50.524
R1831 B.n1158 B.n1157 50.524
R1832 B.n1157 B.n57 50.524
R1833 B.n1151 B.n1150 50.524
R1834 B.n1150 B.n1149 50.524
R1835 B.n1149 B.n64 50.524
R1836 B.n1143 B.n64 50.524
R1837 B.n1143 B.n1142 50.524
R1838 B.n1142 B.n1141 50.524
R1839 B.n1141 B.n71 50.524
R1840 B.n1135 B.n71 50.524
R1841 B.n1135 B.n1134 50.524
R1842 B.n1134 B.n1133 50.524
R1843 B.n1133 B.n78 50.524
R1844 B.n1127 B.n78 50.524
R1845 B.n1126 B.n1125 50.524
R1846 B.n1125 B.n85 50.524
R1847 B.n1119 B.n85 50.524
R1848 B.n1119 B.n1118 50.524
R1849 B.n1118 B.n1117 50.524
R1850 B.n1117 B.n92 50.524
R1851 B.n1111 B.n92 50.524
R1852 B.n1111 B.n1110 50.524
R1853 B.n1110 B.n1109 50.524
R1854 B.n1109 B.n99 50.524
R1855 B.n1103 B.n99 50.524
R1856 B.n1102 B.n1101 50.524
R1857 B.n1101 B.n106 50.524
R1858 B.n1095 B.n106 50.524
R1859 B.n1095 B.n1094 50.524
R1860 B.n1094 B.n1093 50.524
R1861 B.n1093 B.n113 50.524
R1862 B.n1087 B.n113 50.524
R1863 B.n1087 B.n1086 50.524
R1864 B.n1086 B.n1085 50.524
R1865 B.n1085 B.n120 50.524
R1866 B.n1079 B.n120 50.524
R1867 B.n1079 B.n1078 50.524
R1868 B.n1078 B.n1077 50.524
R1869 B.n1077 B.n127 50.524
R1870 B.n1071 B.n1070 50.524
R1871 B.n1070 B.n1069 50.524
R1872 B.n1069 B.n134 50.524
R1873 B.n1063 B.n134 50.524
R1874 B.n1063 B.n1062 50.524
R1875 B.n1062 B.n1061 50.524
R1876 B.n1061 B.n141 50.524
R1877 B.n1055 B.n141 50.524
R1878 B.n1055 B.n1054 50.524
R1879 B.t7 B.n403 49.038
R1880 B.t3 B.n57 49.038
R1881 B.n435 B.t5 44.58
R1882 B.t6 B.n1126 44.58
R1883 B.t9 B.n379 41.6081
R1884 B.t8 B.n36 41.6081
R1885 B.n459 B.t2 37.1501
R1886 B.t0 B.n1102 37.1501
R1887 B.t4 B.n355 34.1781
R1888 B.t1 B.n15 34.1781
R1889 B.n193 B.n143 33.8737
R1890 B.n1050 B.n1049 33.8737
R1891 B.n706 B.n705 33.8737
R1892 B.n700 B.n501 33.8737
R1893 B.t15 B.n483 31.2062
R1894 B.t11 B.n127 31.2062
R1895 B.n733 B.t15 19.3183
R1896 B.n1071 B.t11 19.3183
R1897 B B.n1217 18.0485
R1898 B.n925 B.t4 16.3463
R1899 B.n1199 B.t1 16.3463
R1900 B.n781 B.t2 13.3744
R1901 B.n1103 B.t0 13.3744
R1902 B.n194 B.n193 10.6151
R1903 B.n197 B.n194 10.6151
R1904 B.n198 B.n197 10.6151
R1905 B.n201 B.n198 10.6151
R1906 B.n202 B.n201 10.6151
R1907 B.n205 B.n202 10.6151
R1908 B.n206 B.n205 10.6151
R1909 B.n209 B.n206 10.6151
R1910 B.n210 B.n209 10.6151
R1911 B.n213 B.n210 10.6151
R1912 B.n214 B.n213 10.6151
R1913 B.n217 B.n214 10.6151
R1914 B.n218 B.n217 10.6151
R1915 B.n221 B.n218 10.6151
R1916 B.n222 B.n221 10.6151
R1917 B.n225 B.n222 10.6151
R1918 B.n226 B.n225 10.6151
R1919 B.n229 B.n226 10.6151
R1920 B.n230 B.n229 10.6151
R1921 B.n233 B.n230 10.6151
R1922 B.n234 B.n233 10.6151
R1923 B.n237 B.n234 10.6151
R1924 B.n238 B.n237 10.6151
R1925 B.n241 B.n238 10.6151
R1926 B.n242 B.n241 10.6151
R1927 B.n245 B.n242 10.6151
R1928 B.n246 B.n245 10.6151
R1929 B.n249 B.n246 10.6151
R1930 B.n250 B.n249 10.6151
R1931 B.n253 B.n250 10.6151
R1932 B.n254 B.n253 10.6151
R1933 B.n257 B.n254 10.6151
R1934 B.n258 B.n257 10.6151
R1935 B.n262 B.n261 10.6151
R1936 B.n265 B.n262 10.6151
R1937 B.n266 B.n265 10.6151
R1938 B.n269 B.n266 10.6151
R1939 B.n270 B.n269 10.6151
R1940 B.n273 B.n270 10.6151
R1941 B.n274 B.n273 10.6151
R1942 B.n277 B.n274 10.6151
R1943 B.n278 B.n277 10.6151
R1944 B.n282 B.n281 10.6151
R1945 B.n285 B.n282 10.6151
R1946 B.n286 B.n285 10.6151
R1947 B.n289 B.n286 10.6151
R1948 B.n290 B.n289 10.6151
R1949 B.n293 B.n290 10.6151
R1950 B.n294 B.n293 10.6151
R1951 B.n297 B.n294 10.6151
R1952 B.n298 B.n297 10.6151
R1953 B.n301 B.n298 10.6151
R1954 B.n302 B.n301 10.6151
R1955 B.n305 B.n302 10.6151
R1956 B.n306 B.n305 10.6151
R1957 B.n309 B.n306 10.6151
R1958 B.n310 B.n309 10.6151
R1959 B.n313 B.n310 10.6151
R1960 B.n314 B.n313 10.6151
R1961 B.n317 B.n314 10.6151
R1962 B.n318 B.n317 10.6151
R1963 B.n321 B.n318 10.6151
R1964 B.n322 B.n321 10.6151
R1965 B.n325 B.n322 10.6151
R1966 B.n326 B.n325 10.6151
R1967 B.n329 B.n326 10.6151
R1968 B.n330 B.n329 10.6151
R1969 B.n333 B.n330 10.6151
R1970 B.n334 B.n333 10.6151
R1971 B.n337 B.n334 10.6151
R1972 B.n338 B.n337 10.6151
R1973 B.n341 B.n338 10.6151
R1974 B.n343 B.n341 10.6151
R1975 B.n344 B.n343 10.6151
R1976 B.n1050 B.n344 10.6151
R1977 B.n707 B.n706 10.6151
R1978 B.n707 B.n497 10.6151
R1979 B.n717 B.n497 10.6151
R1980 B.n718 B.n717 10.6151
R1981 B.n719 B.n718 10.6151
R1982 B.n719 B.n489 10.6151
R1983 B.n729 B.n489 10.6151
R1984 B.n730 B.n729 10.6151
R1985 B.n731 B.n730 10.6151
R1986 B.n731 B.n481 10.6151
R1987 B.n741 B.n481 10.6151
R1988 B.n742 B.n741 10.6151
R1989 B.n743 B.n742 10.6151
R1990 B.n743 B.n473 10.6151
R1991 B.n753 B.n473 10.6151
R1992 B.n754 B.n753 10.6151
R1993 B.n755 B.n754 10.6151
R1994 B.n755 B.n465 10.6151
R1995 B.n765 B.n465 10.6151
R1996 B.n766 B.n765 10.6151
R1997 B.n767 B.n766 10.6151
R1998 B.n767 B.n456 10.6151
R1999 B.n777 B.n456 10.6151
R2000 B.n778 B.n777 10.6151
R2001 B.n779 B.n778 10.6151
R2002 B.n779 B.n449 10.6151
R2003 B.n789 B.n449 10.6151
R2004 B.n790 B.n789 10.6151
R2005 B.n791 B.n790 10.6151
R2006 B.n791 B.n441 10.6151
R2007 B.n801 B.n441 10.6151
R2008 B.n802 B.n801 10.6151
R2009 B.n803 B.n802 10.6151
R2010 B.n803 B.n432 10.6151
R2011 B.n813 B.n432 10.6151
R2012 B.n814 B.n813 10.6151
R2013 B.n815 B.n814 10.6151
R2014 B.n815 B.n425 10.6151
R2015 B.n825 B.n425 10.6151
R2016 B.n826 B.n825 10.6151
R2017 B.n827 B.n826 10.6151
R2018 B.n827 B.n417 10.6151
R2019 B.n837 B.n417 10.6151
R2020 B.n838 B.n837 10.6151
R2021 B.n839 B.n838 10.6151
R2022 B.n839 B.n409 10.6151
R2023 B.n849 B.n409 10.6151
R2024 B.n850 B.n849 10.6151
R2025 B.n851 B.n850 10.6151
R2026 B.n851 B.n401 10.6151
R2027 B.n861 B.n401 10.6151
R2028 B.n862 B.n861 10.6151
R2029 B.n863 B.n862 10.6151
R2030 B.n863 B.n393 10.6151
R2031 B.n873 B.n393 10.6151
R2032 B.n874 B.n873 10.6151
R2033 B.n875 B.n874 10.6151
R2034 B.n875 B.n385 10.6151
R2035 B.n885 B.n385 10.6151
R2036 B.n886 B.n885 10.6151
R2037 B.n887 B.n886 10.6151
R2038 B.n887 B.n377 10.6151
R2039 B.n897 B.n377 10.6151
R2040 B.n898 B.n897 10.6151
R2041 B.n899 B.n898 10.6151
R2042 B.n899 B.n369 10.6151
R2043 B.n909 B.n369 10.6151
R2044 B.n910 B.n909 10.6151
R2045 B.n911 B.n910 10.6151
R2046 B.n911 B.n361 10.6151
R2047 B.n921 B.n361 10.6151
R2048 B.n922 B.n921 10.6151
R2049 B.n923 B.n922 10.6151
R2050 B.n923 B.n353 10.6151
R2051 B.n933 B.n353 10.6151
R2052 B.n934 B.n933 10.6151
R2053 B.n936 B.n934 10.6151
R2054 B.n936 B.n935 10.6151
R2055 B.n935 B.n345 10.6151
R2056 B.n947 B.n345 10.6151
R2057 B.n948 B.n947 10.6151
R2058 B.n949 B.n948 10.6151
R2059 B.n950 B.n949 10.6151
R2060 B.n952 B.n950 10.6151
R2061 B.n953 B.n952 10.6151
R2062 B.n954 B.n953 10.6151
R2063 B.n955 B.n954 10.6151
R2064 B.n957 B.n955 10.6151
R2065 B.n958 B.n957 10.6151
R2066 B.n959 B.n958 10.6151
R2067 B.n960 B.n959 10.6151
R2068 B.n962 B.n960 10.6151
R2069 B.n963 B.n962 10.6151
R2070 B.n964 B.n963 10.6151
R2071 B.n965 B.n964 10.6151
R2072 B.n967 B.n965 10.6151
R2073 B.n968 B.n967 10.6151
R2074 B.n969 B.n968 10.6151
R2075 B.n970 B.n969 10.6151
R2076 B.n972 B.n970 10.6151
R2077 B.n973 B.n972 10.6151
R2078 B.n974 B.n973 10.6151
R2079 B.n975 B.n974 10.6151
R2080 B.n977 B.n975 10.6151
R2081 B.n978 B.n977 10.6151
R2082 B.n979 B.n978 10.6151
R2083 B.n980 B.n979 10.6151
R2084 B.n982 B.n980 10.6151
R2085 B.n983 B.n982 10.6151
R2086 B.n984 B.n983 10.6151
R2087 B.n985 B.n984 10.6151
R2088 B.n987 B.n985 10.6151
R2089 B.n988 B.n987 10.6151
R2090 B.n989 B.n988 10.6151
R2091 B.n990 B.n989 10.6151
R2092 B.n992 B.n990 10.6151
R2093 B.n993 B.n992 10.6151
R2094 B.n994 B.n993 10.6151
R2095 B.n995 B.n994 10.6151
R2096 B.n997 B.n995 10.6151
R2097 B.n998 B.n997 10.6151
R2098 B.n999 B.n998 10.6151
R2099 B.n1000 B.n999 10.6151
R2100 B.n1002 B.n1000 10.6151
R2101 B.n1003 B.n1002 10.6151
R2102 B.n1004 B.n1003 10.6151
R2103 B.n1005 B.n1004 10.6151
R2104 B.n1007 B.n1005 10.6151
R2105 B.n1008 B.n1007 10.6151
R2106 B.n1009 B.n1008 10.6151
R2107 B.n1010 B.n1009 10.6151
R2108 B.n1012 B.n1010 10.6151
R2109 B.n1013 B.n1012 10.6151
R2110 B.n1014 B.n1013 10.6151
R2111 B.n1015 B.n1014 10.6151
R2112 B.n1017 B.n1015 10.6151
R2113 B.n1018 B.n1017 10.6151
R2114 B.n1019 B.n1018 10.6151
R2115 B.n1020 B.n1019 10.6151
R2116 B.n1022 B.n1020 10.6151
R2117 B.n1023 B.n1022 10.6151
R2118 B.n1024 B.n1023 10.6151
R2119 B.n1025 B.n1024 10.6151
R2120 B.n1027 B.n1025 10.6151
R2121 B.n1028 B.n1027 10.6151
R2122 B.n1029 B.n1028 10.6151
R2123 B.n1030 B.n1029 10.6151
R2124 B.n1032 B.n1030 10.6151
R2125 B.n1033 B.n1032 10.6151
R2126 B.n1034 B.n1033 10.6151
R2127 B.n1035 B.n1034 10.6151
R2128 B.n1037 B.n1035 10.6151
R2129 B.n1038 B.n1037 10.6151
R2130 B.n1039 B.n1038 10.6151
R2131 B.n1040 B.n1039 10.6151
R2132 B.n1042 B.n1040 10.6151
R2133 B.n1043 B.n1042 10.6151
R2134 B.n1044 B.n1043 10.6151
R2135 B.n1045 B.n1044 10.6151
R2136 B.n1047 B.n1045 10.6151
R2137 B.n1048 B.n1047 10.6151
R2138 B.n1049 B.n1048 10.6151
R2139 B.n700 B.n699 10.6151
R2140 B.n699 B.n698 10.6151
R2141 B.n698 B.n697 10.6151
R2142 B.n697 B.n695 10.6151
R2143 B.n695 B.n692 10.6151
R2144 B.n692 B.n691 10.6151
R2145 B.n691 B.n688 10.6151
R2146 B.n688 B.n687 10.6151
R2147 B.n687 B.n684 10.6151
R2148 B.n684 B.n683 10.6151
R2149 B.n683 B.n680 10.6151
R2150 B.n680 B.n679 10.6151
R2151 B.n679 B.n676 10.6151
R2152 B.n676 B.n675 10.6151
R2153 B.n675 B.n672 10.6151
R2154 B.n672 B.n671 10.6151
R2155 B.n671 B.n668 10.6151
R2156 B.n668 B.n667 10.6151
R2157 B.n667 B.n664 10.6151
R2158 B.n664 B.n663 10.6151
R2159 B.n663 B.n660 10.6151
R2160 B.n660 B.n659 10.6151
R2161 B.n659 B.n656 10.6151
R2162 B.n656 B.n655 10.6151
R2163 B.n655 B.n652 10.6151
R2164 B.n652 B.n651 10.6151
R2165 B.n651 B.n648 10.6151
R2166 B.n648 B.n647 10.6151
R2167 B.n647 B.n644 10.6151
R2168 B.n644 B.n643 10.6151
R2169 B.n643 B.n640 10.6151
R2170 B.n640 B.n639 10.6151
R2171 B.n639 B.n636 10.6151
R2172 B.n634 B.n631 10.6151
R2173 B.n631 B.n630 10.6151
R2174 B.n630 B.n627 10.6151
R2175 B.n627 B.n626 10.6151
R2176 B.n626 B.n623 10.6151
R2177 B.n623 B.n622 10.6151
R2178 B.n622 B.n619 10.6151
R2179 B.n619 B.n618 10.6151
R2180 B.n618 B.n615 10.6151
R2181 B.n613 B.n610 10.6151
R2182 B.n610 B.n609 10.6151
R2183 B.n609 B.n606 10.6151
R2184 B.n606 B.n605 10.6151
R2185 B.n605 B.n602 10.6151
R2186 B.n602 B.n601 10.6151
R2187 B.n601 B.n598 10.6151
R2188 B.n598 B.n597 10.6151
R2189 B.n597 B.n594 10.6151
R2190 B.n594 B.n593 10.6151
R2191 B.n593 B.n590 10.6151
R2192 B.n590 B.n589 10.6151
R2193 B.n589 B.n586 10.6151
R2194 B.n586 B.n585 10.6151
R2195 B.n585 B.n582 10.6151
R2196 B.n582 B.n581 10.6151
R2197 B.n581 B.n578 10.6151
R2198 B.n578 B.n577 10.6151
R2199 B.n577 B.n574 10.6151
R2200 B.n574 B.n573 10.6151
R2201 B.n573 B.n570 10.6151
R2202 B.n570 B.n569 10.6151
R2203 B.n569 B.n566 10.6151
R2204 B.n566 B.n565 10.6151
R2205 B.n565 B.n562 10.6151
R2206 B.n562 B.n561 10.6151
R2207 B.n561 B.n558 10.6151
R2208 B.n558 B.n557 10.6151
R2209 B.n557 B.n554 10.6151
R2210 B.n554 B.n553 10.6151
R2211 B.n553 B.n550 10.6151
R2212 B.n550 B.n505 10.6151
R2213 B.n705 B.n505 10.6151
R2214 B.n711 B.n501 10.6151
R2215 B.n712 B.n711 10.6151
R2216 B.n713 B.n712 10.6151
R2217 B.n713 B.n493 10.6151
R2218 B.n723 B.n493 10.6151
R2219 B.n724 B.n723 10.6151
R2220 B.n725 B.n724 10.6151
R2221 B.n725 B.n485 10.6151
R2222 B.n735 B.n485 10.6151
R2223 B.n736 B.n735 10.6151
R2224 B.n737 B.n736 10.6151
R2225 B.n737 B.n477 10.6151
R2226 B.n747 B.n477 10.6151
R2227 B.n748 B.n747 10.6151
R2228 B.n749 B.n748 10.6151
R2229 B.n749 B.n469 10.6151
R2230 B.n759 B.n469 10.6151
R2231 B.n760 B.n759 10.6151
R2232 B.n761 B.n760 10.6151
R2233 B.n761 B.n461 10.6151
R2234 B.n771 B.n461 10.6151
R2235 B.n772 B.n771 10.6151
R2236 B.n773 B.n772 10.6151
R2237 B.n773 B.n453 10.6151
R2238 B.n783 B.n453 10.6151
R2239 B.n784 B.n783 10.6151
R2240 B.n785 B.n784 10.6151
R2241 B.n785 B.n445 10.6151
R2242 B.n795 B.n445 10.6151
R2243 B.n796 B.n795 10.6151
R2244 B.n797 B.n796 10.6151
R2245 B.n797 B.n437 10.6151
R2246 B.n807 B.n437 10.6151
R2247 B.n808 B.n807 10.6151
R2248 B.n809 B.n808 10.6151
R2249 B.n809 B.n429 10.6151
R2250 B.n819 B.n429 10.6151
R2251 B.n820 B.n819 10.6151
R2252 B.n821 B.n820 10.6151
R2253 B.n821 B.n421 10.6151
R2254 B.n831 B.n421 10.6151
R2255 B.n832 B.n831 10.6151
R2256 B.n833 B.n832 10.6151
R2257 B.n833 B.n413 10.6151
R2258 B.n843 B.n413 10.6151
R2259 B.n844 B.n843 10.6151
R2260 B.n845 B.n844 10.6151
R2261 B.n845 B.n405 10.6151
R2262 B.n855 B.n405 10.6151
R2263 B.n856 B.n855 10.6151
R2264 B.n857 B.n856 10.6151
R2265 B.n857 B.n397 10.6151
R2266 B.n867 B.n397 10.6151
R2267 B.n868 B.n867 10.6151
R2268 B.n869 B.n868 10.6151
R2269 B.n869 B.n389 10.6151
R2270 B.n879 B.n389 10.6151
R2271 B.n880 B.n879 10.6151
R2272 B.n881 B.n880 10.6151
R2273 B.n881 B.n381 10.6151
R2274 B.n891 B.n381 10.6151
R2275 B.n892 B.n891 10.6151
R2276 B.n893 B.n892 10.6151
R2277 B.n893 B.n373 10.6151
R2278 B.n903 B.n373 10.6151
R2279 B.n904 B.n903 10.6151
R2280 B.n905 B.n904 10.6151
R2281 B.n905 B.n365 10.6151
R2282 B.n915 B.n365 10.6151
R2283 B.n916 B.n915 10.6151
R2284 B.n917 B.n916 10.6151
R2285 B.n917 B.n357 10.6151
R2286 B.n927 B.n357 10.6151
R2287 B.n928 B.n927 10.6151
R2288 B.n929 B.n928 10.6151
R2289 B.n929 B.n349 10.6151
R2290 B.n940 B.n349 10.6151
R2291 B.n941 B.n940 10.6151
R2292 B.n942 B.n941 10.6151
R2293 B.n942 B.n0 10.6151
R2294 B.n1211 B.n1 10.6151
R2295 B.n1211 B.n1210 10.6151
R2296 B.n1210 B.n1209 10.6151
R2297 B.n1209 B.n10 10.6151
R2298 B.n1203 B.n10 10.6151
R2299 B.n1203 B.n1202 10.6151
R2300 B.n1202 B.n1201 10.6151
R2301 B.n1201 B.n17 10.6151
R2302 B.n1195 B.n17 10.6151
R2303 B.n1195 B.n1194 10.6151
R2304 B.n1194 B.n1193 10.6151
R2305 B.n1193 B.n24 10.6151
R2306 B.n1187 B.n24 10.6151
R2307 B.n1187 B.n1186 10.6151
R2308 B.n1186 B.n1185 10.6151
R2309 B.n1185 B.n31 10.6151
R2310 B.n1179 B.n31 10.6151
R2311 B.n1179 B.n1178 10.6151
R2312 B.n1178 B.n1177 10.6151
R2313 B.n1177 B.n38 10.6151
R2314 B.n1171 B.n38 10.6151
R2315 B.n1171 B.n1170 10.6151
R2316 B.n1170 B.n1169 10.6151
R2317 B.n1169 B.n45 10.6151
R2318 B.n1163 B.n45 10.6151
R2319 B.n1163 B.n1162 10.6151
R2320 B.n1162 B.n1161 10.6151
R2321 B.n1161 B.n52 10.6151
R2322 B.n1155 B.n52 10.6151
R2323 B.n1155 B.n1154 10.6151
R2324 B.n1154 B.n1153 10.6151
R2325 B.n1153 B.n59 10.6151
R2326 B.n1147 B.n59 10.6151
R2327 B.n1147 B.n1146 10.6151
R2328 B.n1146 B.n1145 10.6151
R2329 B.n1145 B.n66 10.6151
R2330 B.n1139 B.n66 10.6151
R2331 B.n1139 B.n1138 10.6151
R2332 B.n1138 B.n1137 10.6151
R2333 B.n1137 B.n73 10.6151
R2334 B.n1131 B.n73 10.6151
R2335 B.n1131 B.n1130 10.6151
R2336 B.n1130 B.n1129 10.6151
R2337 B.n1129 B.n80 10.6151
R2338 B.n1123 B.n80 10.6151
R2339 B.n1123 B.n1122 10.6151
R2340 B.n1122 B.n1121 10.6151
R2341 B.n1121 B.n87 10.6151
R2342 B.n1115 B.n87 10.6151
R2343 B.n1115 B.n1114 10.6151
R2344 B.n1114 B.n1113 10.6151
R2345 B.n1113 B.n94 10.6151
R2346 B.n1107 B.n94 10.6151
R2347 B.n1107 B.n1106 10.6151
R2348 B.n1106 B.n1105 10.6151
R2349 B.n1105 B.n101 10.6151
R2350 B.n1099 B.n101 10.6151
R2351 B.n1099 B.n1098 10.6151
R2352 B.n1098 B.n1097 10.6151
R2353 B.n1097 B.n108 10.6151
R2354 B.n1091 B.n108 10.6151
R2355 B.n1091 B.n1090 10.6151
R2356 B.n1090 B.n1089 10.6151
R2357 B.n1089 B.n115 10.6151
R2358 B.n1083 B.n115 10.6151
R2359 B.n1083 B.n1082 10.6151
R2360 B.n1082 B.n1081 10.6151
R2361 B.n1081 B.n122 10.6151
R2362 B.n1075 B.n122 10.6151
R2363 B.n1075 B.n1074 10.6151
R2364 B.n1074 B.n1073 10.6151
R2365 B.n1073 B.n129 10.6151
R2366 B.n1067 B.n129 10.6151
R2367 B.n1067 B.n1066 10.6151
R2368 B.n1066 B.n1065 10.6151
R2369 B.n1065 B.n136 10.6151
R2370 B.n1059 B.n136 10.6151
R2371 B.n1059 B.n1058 10.6151
R2372 B.n1058 B.n1057 10.6151
R2373 B.n1057 B.n143 10.6151
R2374 B.n258 B.n191 9.36635
R2375 B.n281 B.n188 9.36635
R2376 B.n636 B.n635 9.36635
R2377 B.n614 B.n613 9.36635
R2378 B.n889 B.t9 8.91641
R2379 B.n1175 B.t8 8.91641
R2380 B.n817 B.t5 5.94444
R2381 B.n1127 B.t6 5.94444
R2382 B.n1217 B.n0 2.81026
R2383 B.n1217 B.n1 2.81026
R2384 B.n853 B.t7 1.48648
R2385 B.n1151 B.t3 1.48648
R2386 B.n261 B.n191 1.24928
R2387 B.n278 B.n188 1.24928
R2388 B.n635 B.n634 1.24928
R2389 B.n615 B.n614 1.24928
R2390 VN.n110 VN.n109 161.3
R2391 VN.n108 VN.n57 161.3
R2392 VN.n107 VN.n106 161.3
R2393 VN.n105 VN.n58 161.3
R2394 VN.n104 VN.n103 161.3
R2395 VN.n102 VN.n59 161.3
R2396 VN.n101 VN.n100 161.3
R2397 VN.n99 VN.n60 161.3
R2398 VN.n98 VN.n97 161.3
R2399 VN.n95 VN.n61 161.3
R2400 VN.n94 VN.n93 161.3
R2401 VN.n92 VN.n62 161.3
R2402 VN.n91 VN.n90 161.3
R2403 VN.n89 VN.n63 161.3
R2404 VN.n88 VN.n87 161.3
R2405 VN.n86 VN.n64 161.3
R2406 VN.n85 VN.n84 161.3
R2407 VN.n82 VN.n65 161.3
R2408 VN.n81 VN.n80 161.3
R2409 VN.n79 VN.n66 161.3
R2410 VN.n78 VN.n77 161.3
R2411 VN.n76 VN.n67 161.3
R2412 VN.n75 VN.n74 161.3
R2413 VN.n73 VN.n68 161.3
R2414 VN.n72 VN.n71 161.3
R2415 VN.n54 VN.n53 161.3
R2416 VN.n52 VN.n1 161.3
R2417 VN.n51 VN.n50 161.3
R2418 VN.n49 VN.n2 161.3
R2419 VN.n48 VN.n47 161.3
R2420 VN.n46 VN.n3 161.3
R2421 VN.n45 VN.n44 161.3
R2422 VN.n43 VN.n4 161.3
R2423 VN.n42 VN.n41 161.3
R2424 VN.n39 VN.n5 161.3
R2425 VN.n38 VN.n37 161.3
R2426 VN.n36 VN.n6 161.3
R2427 VN.n35 VN.n34 161.3
R2428 VN.n33 VN.n7 161.3
R2429 VN.n32 VN.n31 161.3
R2430 VN.n30 VN.n8 161.3
R2431 VN.n29 VN.n28 161.3
R2432 VN.n26 VN.n9 161.3
R2433 VN.n25 VN.n24 161.3
R2434 VN.n23 VN.n10 161.3
R2435 VN.n22 VN.n21 161.3
R2436 VN.n20 VN.n11 161.3
R2437 VN.n19 VN.n18 161.3
R2438 VN.n17 VN.n12 161.3
R2439 VN.n16 VN.n15 161.3
R2440 VN.n69 VN.t7 92.6444
R2441 VN.n13 VN.t3 92.6444
R2442 VN.n55 VN.n0 89.5781
R2443 VN.n111 VN.n56 89.5781
R2444 VN.n14 VN.t1 60.4408
R2445 VN.n27 VN.t8 60.4408
R2446 VN.n40 VN.t6 60.4408
R2447 VN.n0 VN.t5 60.4408
R2448 VN.n70 VN.t9 60.4408
R2449 VN.n83 VN.t0 60.4408
R2450 VN.n96 VN.t4 60.4408
R2451 VN.n56 VN.t2 60.4408
R2452 VN VN.n111 57.9488
R2453 VN.n21 VN.n20 56.5193
R2454 VN.n34 VN.n33 56.5193
R2455 VN.n77 VN.n76 56.5193
R2456 VN.n90 VN.n89 56.5193
R2457 VN.n14 VN.n13 56.4597
R2458 VN.n70 VN.n69 56.4597
R2459 VN.n47 VN.n46 45.8354
R2460 VN.n103 VN.n102 45.8354
R2461 VN.n47 VN.n2 35.1514
R2462 VN.n103 VN.n58 35.1514
R2463 VN.n15 VN.n12 24.4675
R2464 VN.n19 VN.n12 24.4675
R2465 VN.n20 VN.n19 24.4675
R2466 VN.n21 VN.n10 24.4675
R2467 VN.n25 VN.n10 24.4675
R2468 VN.n26 VN.n25 24.4675
R2469 VN.n28 VN.n8 24.4675
R2470 VN.n32 VN.n8 24.4675
R2471 VN.n33 VN.n32 24.4675
R2472 VN.n34 VN.n6 24.4675
R2473 VN.n38 VN.n6 24.4675
R2474 VN.n39 VN.n38 24.4675
R2475 VN.n41 VN.n4 24.4675
R2476 VN.n45 VN.n4 24.4675
R2477 VN.n46 VN.n45 24.4675
R2478 VN.n51 VN.n2 24.4675
R2479 VN.n52 VN.n51 24.4675
R2480 VN.n53 VN.n52 24.4675
R2481 VN.n76 VN.n75 24.4675
R2482 VN.n75 VN.n68 24.4675
R2483 VN.n71 VN.n68 24.4675
R2484 VN.n89 VN.n88 24.4675
R2485 VN.n88 VN.n64 24.4675
R2486 VN.n84 VN.n64 24.4675
R2487 VN.n82 VN.n81 24.4675
R2488 VN.n81 VN.n66 24.4675
R2489 VN.n77 VN.n66 24.4675
R2490 VN.n102 VN.n101 24.4675
R2491 VN.n101 VN.n60 24.4675
R2492 VN.n97 VN.n60 24.4675
R2493 VN.n95 VN.n94 24.4675
R2494 VN.n94 VN.n62 24.4675
R2495 VN.n90 VN.n62 24.4675
R2496 VN.n109 VN.n108 24.4675
R2497 VN.n108 VN.n107 24.4675
R2498 VN.n107 VN.n58 24.4675
R2499 VN.n15 VN.n14 18.5954
R2500 VN.n40 VN.n39 18.5954
R2501 VN.n71 VN.n70 18.5954
R2502 VN.n96 VN.n95 18.5954
R2503 VN.n27 VN.n26 12.234
R2504 VN.n28 VN.n27 12.234
R2505 VN.n84 VN.n83 12.234
R2506 VN.n83 VN.n82 12.234
R2507 VN.n41 VN.n40 5.87258
R2508 VN.n97 VN.n96 5.87258
R2509 VN.n72 VN.n69 2.5172
R2510 VN.n16 VN.n13 2.5172
R2511 VN.n53 VN.n0 0.48984
R2512 VN.n109 VN.n56 0.48984
R2513 VN.n111 VN.n110 0.354971
R2514 VN.n55 VN.n54 0.354971
R2515 VN VN.n55 0.26696
R2516 VN.n110 VN.n57 0.189894
R2517 VN.n106 VN.n57 0.189894
R2518 VN.n106 VN.n105 0.189894
R2519 VN.n105 VN.n104 0.189894
R2520 VN.n104 VN.n59 0.189894
R2521 VN.n100 VN.n59 0.189894
R2522 VN.n100 VN.n99 0.189894
R2523 VN.n99 VN.n98 0.189894
R2524 VN.n98 VN.n61 0.189894
R2525 VN.n93 VN.n61 0.189894
R2526 VN.n93 VN.n92 0.189894
R2527 VN.n92 VN.n91 0.189894
R2528 VN.n91 VN.n63 0.189894
R2529 VN.n87 VN.n63 0.189894
R2530 VN.n87 VN.n86 0.189894
R2531 VN.n86 VN.n85 0.189894
R2532 VN.n85 VN.n65 0.189894
R2533 VN.n80 VN.n65 0.189894
R2534 VN.n80 VN.n79 0.189894
R2535 VN.n79 VN.n78 0.189894
R2536 VN.n78 VN.n67 0.189894
R2537 VN.n74 VN.n67 0.189894
R2538 VN.n74 VN.n73 0.189894
R2539 VN.n73 VN.n72 0.189894
R2540 VN.n17 VN.n16 0.189894
R2541 VN.n18 VN.n17 0.189894
R2542 VN.n18 VN.n11 0.189894
R2543 VN.n22 VN.n11 0.189894
R2544 VN.n23 VN.n22 0.189894
R2545 VN.n24 VN.n23 0.189894
R2546 VN.n24 VN.n9 0.189894
R2547 VN.n29 VN.n9 0.189894
R2548 VN.n30 VN.n29 0.189894
R2549 VN.n31 VN.n30 0.189894
R2550 VN.n31 VN.n7 0.189894
R2551 VN.n35 VN.n7 0.189894
R2552 VN.n36 VN.n35 0.189894
R2553 VN.n37 VN.n36 0.189894
R2554 VN.n37 VN.n5 0.189894
R2555 VN.n42 VN.n5 0.189894
R2556 VN.n43 VN.n42 0.189894
R2557 VN.n44 VN.n43 0.189894
R2558 VN.n44 VN.n3 0.189894
R2559 VN.n48 VN.n3 0.189894
R2560 VN.n49 VN.n48 0.189894
R2561 VN.n50 VN.n49 0.189894
R2562 VN.n50 VN.n1 0.189894
R2563 VN.n54 VN.n1 0.189894
R2564 VDD2.n1 VDD2.t6 67.0924
R2565 VDD2.n3 VDD2.n2 64.0692
R2566 VDD2 VDD2.n7 64.0664
R2567 VDD2.n4 VDD2.t7 63.5321
R2568 VDD2.n6 VDD2.n5 61.4545
R2569 VDD2.n1 VDD2.n0 61.4543
R2570 VDD2.n4 VDD2.n3 48.8424
R2571 VDD2.n6 VDD2.n4 3.56084
R2572 VDD2.n7 VDD2.t0 2.07815
R2573 VDD2.n7 VDD2.t2 2.07815
R2574 VDD2.n5 VDD2.t5 2.07815
R2575 VDD2.n5 VDD2.t9 2.07815
R2576 VDD2.n2 VDD2.t3 2.07815
R2577 VDD2.n2 VDD2.t4 2.07815
R2578 VDD2.n0 VDD2.t8 2.07815
R2579 VDD2.n0 VDD2.t1 2.07815
R2580 VDD2 VDD2.n6 0.948776
R2581 VDD2.n3 VDD2.n1 0.83524
C0 VN VDD1 0.156081f
C1 VN VTAIL 10.4198f
C2 VTAIL VDD1 10.055f
C3 VN VDD2 9.144929f
C4 VN VP 9.71288f
C5 VDD1 VDD2 2.95589f
C6 VDD1 VP 9.72169f
C7 VTAIL VDD2 10.115299f
C8 VTAIL VP 10.434401f
C9 VDD2 VP 0.736145f
C10 VDD2 B 8.191076f
C11 VDD1 B 8.149543f
C12 VTAIL B 8.107109f
C13 VN B 23.704142f
C14 VP B 22.299063f
C15 VDD2.t6 B 2.16855f
C16 VDD2.t8 B 0.191712f
C17 VDD2.t1 B 0.191712f
C18 VDD2.n0 B 1.68093f
C19 VDD2.n1 B 1.11477f
C20 VDD2.t3 B 0.191712f
C21 VDD2.t4 B 0.191712f
C22 VDD2.n2 B 1.71052f
C23 VDD2.n3 B 3.43551f
C24 VDD2.t7 B 2.13799f
C25 VDD2.n4 B 3.46172f
C26 VDD2.t5 B 0.191712f
C27 VDD2.t9 B 0.191712f
C28 VDD2.n5 B 1.68093f
C29 VDD2.n6 B 0.577836f
C30 VDD2.t0 B 0.191712f
C31 VDD2.t2 B 0.191712f
C32 VDD2.n7 B 1.71047f
C33 VN.t5 B 1.70647f
C34 VN.n0 B 0.668717f
C35 VN.n1 B 0.017424f
C36 VN.n2 B 0.035202f
C37 VN.n3 B 0.017424f
C38 VN.n4 B 0.032474f
C39 VN.n5 B 0.017424f
C40 VN.t6 B 1.70647f
C41 VN.n6 B 0.032474f
C42 VN.n7 B 0.017424f
C43 VN.n8 B 0.032474f
C44 VN.n9 B 0.017424f
C45 VN.t8 B 1.70647f
C46 VN.n10 B 0.032474f
C47 VN.n11 B 0.017424f
C48 VN.n12 B 0.032474f
C49 VN.t3 B 1.96512f
C50 VN.n13 B 0.642604f
C51 VN.t1 B 1.70647f
C52 VN.n14 B 0.672487f
C53 VN.n15 B 0.028626f
C54 VN.n16 B 0.2248f
C55 VN.n17 B 0.017424f
C56 VN.n18 B 0.017424f
C57 VN.n19 B 0.032474f
C58 VN.n20 B 0.022281f
C59 VN.n21 B 0.028593f
C60 VN.n22 B 0.017424f
C61 VN.n23 B 0.017424f
C62 VN.n24 B 0.017424f
C63 VN.n25 B 0.032474f
C64 VN.n26 B 0.024457f
C65 VN.n27 B 0.605472f
C66 VN.n28 B 0.024457f
C67 VN.n29 B 0.017424f
C68 VN.n30 B 0.017424f
C69 VN.n31 B 0.017424f
C70 VN.n32 B 0.032474f
C71 VN.n33 B 0.028593f
C72 VN.n34 B 0.022281f
C73 VN.n35 B 0.017424f
C74 VN.n36 B 0.017424f
C75 VN.n37 B 0.017424f
C76 VN.n38 B 0.032474f
C77 VN.n39 B 0.028626f
C78 VN.n40 B 0.605472f
C79 VN.n41 B 0.020289f
C80 VN.n42 B 0.017424f
C81 VN.n43 B 0.017424f
C82 VN.n44 B 0.017424f
C83 VN.n45 B 0.032474f
C84 VN.n46 B 0.03337f
C85 VN.n47 B 0.014775f
C86 VN.n48 B 0.017424f
C87 VN.n49 B 0.017424f
C88 VN.n50 B 0.017424f
C89 VN.n51 B 0.032474f
C90 VN.n52 B 0.032474f
C91 VN.n53 B 0.016762f
C92 VN.n54 B 0.028122f
C93 VN.n55 B 0.054702f
C94 VN.t2 B 1.70647f
C95 VN.n56 B 0.668717f
C96 VN.n57 B 0.017424f
C97 VN.n58 B 0.035202f
C98 VN.n59 B 0.017424f
C99 VN.n60 B 0.032474f
C100 VN.n61 B 0.017424f
C101 VN.t4 B 1.70647f
C102 VN.n62 B 0.032474f
C103 VN.n63 B 0.017424f
C104 VN.n64 B 0.032474f
C105 VN.n65 B 0.017424f
C106 VN.t0 B 1.70647f
C107 VN.n66 B 0.032474f
C108 VN.n67 B 0.017424f
C109 VN.n68 B 0.032474f
C110 VN.t7 B 1.96512f
C111 VN.n69 B 0.642604f
C112 VN.t9 B 1.70647f
C113 VN.n70 B 0.672487f
C114 VN.n71 B 0.028626f
C115 VN.n72 B 0.2248f
C116 VN.n73 B 0.017424f
C117 VN.n74 B 0.017424f
C118 VN.n75 B 0.032474f
C119 VN.n76 B 0.022281f
C120 VN.n77 B 0.028593f
C121 VN.n78 B 0.017424f
C122 VN.n79 B 0.017424f
C123 VN.n80 B 0.017424f
C124 VN.n81 B 0.032474f
C125 VN.n82 B 0.024457f
C126 VN.n83 B 0.605472f
C127 VN.n84 B 0.024457f
C128 VN.n85 B 0.017424f
C129 VN.n86 B 0.017424f
C130 VN.n87 B 0.017424f
C131 VN.n88 B 0.032474f
C132 VN.n89 B 0.028593f
C133 VN.n90 B 0.022281f
C134 VN.n91 B 0.017424f
C135 VN.n92 B 0.017424f
C136 VN.n93 B 0.017424f
C137 VN.n94 B 0.032474f
C138 VN.n95 B 0.028626f
C139 VN.n96 B 0.605472f
C140 VN.n97 B 0.020289f
C141 VN.n98 B 0.017424f
C142 VN.n99 B 0.017424f
C143 VN.n100 B 0.017424f
C144 VN.n101 B 0.032474f
C145 VN.n102 B 0.03337f
C146 VN.n103 B 0.014775f
C147 VN.n104 B 0.017424f
C148 VN.n105 B 0.017424f
C149 VN.n106 B 0.017424f
C150 VN.n107 B 0.032474f
C151 VN.n108 B 0.032474f
C152 VN.n109 B 0.016762f
C153 VN.n110 B 0.028122f
C154 VN.n111 B 1.23171f
C155 VTAIL.t1 B 0.203353f
C156 VTAIL.t8 B 0.203353f
C157 VTAIL.n0 B 1.70273f
C158 VTAIL.n1 B 0.69738f
C159 VTAIL.t10 B 2.16624f
C160 VTAIL.n2 B 0.860849f
C161 VTAIL.t16 B 0.203353f
C162 VTAIL.t11 B 0.203353f
C163 VTAIL.n3 B 1.70273f
C164 VTAIL.n4 B 0.883772f
C165 VTAIL.t9 B 0.203353f
C166 VTAIL.t17 B 0.203353f
C167 VTAIL.n5 B 1.70273f
C168 VTAIL.n6 B 2.27516f
C169 VTAIL.t2 B 0.203353f
C170 VTAIL.t5 B 0.203353f
C171 VTAIL.n7 B 1.70273f
C172 VTAIL.n8 B 2.27516f
C173 VTAIL.t7 B 0.203353f
C174 VTAIL.t19 B 0.203353f
C175 VTAIL.n9 B 1.70273f
C176 VTAIL.n10 B 0.883767f
C177 VTAIL.t4 B 2.16625f
C178 VTAIL.n11 B 0.860833f
C179 VTAIL.t14 B 0.203353f
C180 VTAIL.t12 B 0.203353f
C181 VTAIL.n12 B 1.70273f
C182 VTAIL.n13 B 0.769756f
C183 VTAIL.t15 B 0.203353f
C184 VTAIL.t18 B 0.203353f
C185 VTAIL.n14 B 1.70273f
C186 VTAIL.n15 B 0.883767f
C187 VTAIL.t13 B 2.16624f
C188 VTAIL.n16 B 2.05647f
C189 VTAIL.t0 B 2.16624f
C190 VTAIL.n17 B 2.05647f
C191 VTAIL.t3 B 0.203353f
C192 VTAIL.t6 B 0.203353f
C193 VTAIL.n18 B 1.70273f
C194 VTAIL.n19 B 0.646375f
C195 VDD1.t4 B 2.21777f
C196 VDD1.t6 B 0.196063f
C197 VDD1.t8 B 0.196063f
C198 VDD1.n0 B 1.71908f
C199 VDD1.n1 B 1.14886f
C200 VDD1.t3 B 2.21776f
C201 VDD1.t0 B 0.196063f
C202 VDD1.t2 B 0.196063f
C203 VDD1.n2 B 1.71908f
C204 VDD1.n3 B 1.14007f
C205 VDD1.t1 B 0.196063f
C206 VDD1.t9 B 0.196063f
C207 VDD1.n4 B 1.74934f
C208 VDD1.n5 B 3.67604f
C209 VDD1.t5 B 0.196063f
C210 VDD1.t7 B 0.196063f
C211 VDD1.n6 B 1.71907f
C212 VDD1.n7 B 3.62574f
C213 VP.t8 B 1.743f
C214 VP.n0 B 0.683031f
C215 VP.n1 B 0.017797f
C216 VP.n2 B 0.035956f
C217 VP.n3 B 0.017797f
C218 VP.n4 B 0.033169f
C219 VP.n5 B 0.017797f
C220 VP.t7 B 1.743f
C221 VP.n6 B 0.033169f
C222 VP.n7 B 0.017797f
C223 VP.n8 B 0.033169f
C224 VP.n9 B 0.017797f
C225 VP.t2 B 1.743f
C226 VP.n10 B 0.033169f
C227 VP.n11 B 0.017797f
C228 VP.n12 B 0.033169f
C229 VP.n13 B 0.017797f
C230 VP.t1 B 1.743f
C231 VP.n14 B 0.033169f
C232 VP.n15 B 0.017797f
C233 VP.n16 B 0.033169f
C234 VP.n17 B 0.028724f
C235 VP.t9 B 1.743f
C236 VP.t5 B 1.743f
C237 VP.n18 B 0.683031f
C238 VP.n19 B 0.017797f
C239 VP.n20 B 0.035956f
C240 VP.n21 B 0.017797f
C241 VP.n22 B 0.033169f
C242 VP.n23 B 0.017797f
C243 VP.t0 B 1.743f
C244 VP.n24 B 0.033169f
C245 VP.n25 B 0.017797f
C246 VP.n26 B 0.033169f
C247 VP.n27 B 0.017797f
C248 VP.t3 B 1.743f
C249 VP.n28 B 0.033169f
C250 VP.n29 B 0.017797f
C251 VP.n30 B 0.033169f
C252 VP.t4 B 2.00719f
C253 VP.n31 B 0.656359f
C254 VP.t6 B 1.743f
C255 VP.n32 B 0.686881f
C256 VP.n33 B 0.029239f
C257 VP.n34 B 0.229612f
C258 VP.n35 B 0.017797f
C259 VP.n36 B 0.017797f
C260 VP.n37 B 0.033169f
C261 VP.n38 B 0.022758f
C262 VP.n39 B 0.029205f
C263 VP.n40 B 0.017797f
C264 VP.n41 B 0.017797f
C265 VP.n42 B 0.017797f
C266 VP.n43 B 0.033169f
C267 VP.n44 B 0.024981f
C268 VP.n45 B 0.618432f
C269 VP.n46 B 0.024981f
C270 VP.n47 B 0.017797f
C271 VP.n48 B 0.017797f
C272 VP.n49 B 0.017797f
C273 VP.n50 B 0.033169f
C274 VP.n51 B 0.029205f
C275 VP.n52 B 0.022758f
C276 VP.n53 B 0.017797f
C277 VP.n54 B 0.017797f
C278 VP.n55 B 0.017797f
C279 VP.n56 B 0.033169f
C280 VP.n57 B 0.029239f
C281 VP.n58 B 0.618432f
C282 VP.n59 B 0.020723f
C283 VP.n60 B 0.017797f
C284 VP.n61 B 0.017797f
C285 VP.n62 B 0.017797f
C286 VP.n63 B 0.033169f
C287 VP.n64 B 0.034085f
C288 VP.n65 B 0.015091f
C289 VP.n66 B 0.017797f
C290 VP.n67 B 0.017797f
C291 VP.n68 B 0.017797f
C292 VP.n69 B 0.033169f
C293 VP.n70 B 0.033169f
C294 VP.n71 B 0.017121f
C295 VP.n72 B 0.028724f
C296 VP.n73 B 1.25113f
C297 VP.n74 B 1.2622f
C298 VP.n75 B 0.683031f
C299 VP.n76 B 0.017121f
C300 VP.n77 B 0.033169f
C301 VP.n78 B 0.017797f
C302 VP.n79 B 0.017797f
C303 VP.n80 B 0.017797f
C304 VP.n81 B 0.035956f
C305 VP.n82 B 0.015091f
C306 VP.n83 B 0.034085f
C307 VP.n84 B 0.017797f
C308 VP.n85 B 0.017797f
C309 VP.n86 B 0.017797f
C310 VP.n87 B 0.033169f
C311 VP.n88 B 0.020723f
C312 VP.n89 B 0.618432f
C313 VP.n90 B 0.029239f
C314 VP.n91 B 0.017797f
C315 VP.n92 B 0.017797f
C316 VP.n93 B 0.017797f
C317 VP.n94 B 0.033169f
C318 VP.n95 B 0.022758f
C319 VP.n96 B 0.029205f
C320 VP.n97 B 0.017797f
C321 VP.n98 B 0.017797f
C322 VP.n99 B 0.017797f
C323 VP.n100 B 0.033169f
C324 VP.n101 B 0.024981f
C325 VP.n102 B 0.618432f
C326 VP.n103 B 0.024981f
C327 VP.n104 B 0.017797f
C328 VP.n105 B 0.017797f
C329 VP.n106 B 0.017797f
C330 VP.n107 B 0.033169f
C331 VP.n108 B 0.029205f
C332 VP.n109 B 0.022758f
C333 VP.n110 B 0.017797f
C334 VP.n111 B 0.017797f
C335 VP.n112 B 0.017797f
C336 VP.n113 B 0.033169f
C337 VP.n114 B 0.029239f
C338 VP.n115 B 0.618432f
C339 VP.n116 B 0.020723f
C340 VP.n117 B 0.017797f
C341 VP.n118 B 0.017797f
C342 VP.n119 B 0.017797f
C343 VP.n120 B 0.033169f
C344 VP.n121 B 0.034085f
C345 VP.n122 B 0.015091f
C346 VP.n123 B 0.017797f
C347 VP.n124 B 0.017797f
C348 VP.n125 B 0.017797f
C349 VP.n126 B 0.033169f
C350 VP.n127 B 0.033169f
C351 VP.n128 B 0.017121f
C352 VP.n129 B 0.028724f
C353 VP.n130 B 0.055873f
.ends

