* NGSPICE file created from diff_pair_sample_1467.ext - technology: sky130A

.subckt diff_pair_sample_1467 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=5.538 ps=29.18 w=14.2 l=3.55
X1 VTAIL.t1 VN.t0 VDD2.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X2 VDD1.t8 VP.t1 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=2.343 ps=14.53 w=14.2 l=3.55
X3 VDD1.t7 VP.t2 VTAIL.t19 B.t6 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=5.538 ps=29.18 w=14.2 l=3.55
X4 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=0 ps=0 w=14.2 l=3.55
X6 VDD2.t7 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=5.538 ps=29.18 w=14.2 l=3.55
X7 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=0 ps=0 w=14.2 l=3.55
X8 VTAIL.t7 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X9 VTAIL.t18 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X10 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X11 VTAIL.t11 VP.t4 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X12 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=0 ps=0 w=14.2 l=3.55
X13 VDD2.t4 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=2.343 ps=14.53 w=14.2 l=3.55
X14 VTAIL.t17 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X15 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=5.538 ps=29.18 w=14.2 l=3.55
X16 VDD2.t2 VN.t7 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=2.343 ps=14.53 w=14.2 l=3.55
X17 VDD2.t1 VN.t8 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X18 VDD1.t3 VP.t6 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X19 VTAIL.t15 VP.t7 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=0 ps=0 w=14.2 l=3.55
X21 VTAIL.t5 VN.t9 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
X22 VDD1.t1 VP.t8 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=5.538 pd=29.18 as=2.343 ps=14.53 w=14.2 l=3.55
X23 VDD1.t0 VP.t9 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=2.343 pd=14.53 as=2.343 ps=14.53 w=14.2 l=3.55
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n42 VP.n25 161.3
R8 VP.n44 VP.n43 161.3
R9 VP.n45 VP.n24 161.3
R10 VP.n47 VP.n46 161.3
R11 VP.n48 VP.n23 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n51 VP.n22 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n21 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n20 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n19 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n64 VP.n18 161.3
R22 VP.n66 VP.n65 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n4 161.3
R31 VP.n105 VP.n104 161.3
R32 VP.n102 VP.n5 161.3
R33 VP.n101 VP.n100 161.3
R34 VP.n99 VP.n6 161.3
R35 VP.n98 VP.n97 161.3
R36 VP.n96 VP.n7 161.3
R37 VP.n95 VP.n94 161.3
R38 VP.n93 VP.n8 161.3
R39 VP.n92 VP.n91 161.3
R40 VP.n90 VP.n9 161.3
R41 VP.n89 VP.n88 161.3
R42 VP.n87 VP.n10 161.3
R43 VP.n86 VP.n85 161.3
R44 VP.n84 VP.n11 161.3
R45 VP.n83 VP.n82 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n79 VP.n13 161.3
R48 VP.n78 VP.n77 161.3
R49 VP.n76 VP.n14 161.3
R50 VP.n75 VP.n74 161.3
R51 VP.n73 VP.n15 161.3
R52 VP.n72 VP.n71 161.3
R53 VP.n70 VP.n16 161.3
R54 VP.n30 VP.t1 130.255
R55 VP.n8 VP.t9 96.4005
R56 VP.n68 VP.t8 96.4005
R57 VP.n12 VP.t7 96.4005
R58 VP.n103 VP.t3 96.4005
R59 VP.n0 VP.t2 96.4005
R60 VP.n25 VP.t6 96.4005
R61 VP.n17 VP.t0 96.4005
R62 VP.n52 VP.t5 96.4005
R63 VP.n29 VP.t4 96.4005
R64 VP.n69 VP.n68 77.4578
R65 VP.n118 VP.n0 77.4578
R66 VP.n67 VP.n17 77.4578
R67 VP.n69 VP.n67 60.0905
R68 VP.n74 VP.n14 56.5617
R69 VP.n110 VP.n2 56.5617
R70 VP.n59 VP.n19 56.5617
R71 VP.n30 VP.n29 56.2361
R72 VP.n89 VP.n10 46.3896
R73 VP.n97 VP.n6 46.3896
R74 VP.n46 VP.n23 46.3896
R75 VP.n38 VP.n27 46.3896
R76 VP.n85 VP.n10 34.7644
R77 VP.n101 VP.n6 34.7644
R78 VP.n50 VP.n23 34.7644
R79 VP.n34 VP.n27 34.7644
R80 VP.n72 VP.n16 24.5923
R81 VP.n73 VP.n72 24.5923
R82 VP.n74 VP.n73 24.5923
R83 VP.n78 VP.n14 24.5923
R84 VP.n79 VP.n78 24.5923
R85 VP.n80 VP.n79 24.5923
R86 VP.n84 VP.n83 24.5923
R87 VP.n85 VP.n84 24.5923
R88 VP.n90 VP.n89 24.5923
R89 VP.n91 VP.n90 24.5923
R90 VP.n91 VP.n8 24.5923
R91 VP.n95 VP.n8 24.5923
R92 VP.n96 VP.n95 24.5923
R93 VP.n97 VP.n96 24.5923
R94 VP.n102 VP.n101 24.5923
R95 VP.n104 VP.n102 24.5923
R96 VP.n108 VP.n4 24.5923
R97 VP.n109 VP.n108 24.5923
R98 VP.n110 VP.n109 24.5923
R99 VP.n114 VP.n2 24.5923
R100 VP.n115 VP.n114 24.5923
R101 VP.n116 VP.n115 24.5923
R102 VP.n63 VP.n19 24.5923
R103 VP.n64 VP.n63 24.5923
R104 VP.n65 VP.n64 24.5923
R105 VP.n51 VP.n50 24.5923
R106 VP.n53 VP.n51 24.5923
R107 VP.n57 VP.n21 24.5923
R108 VP.n58 VP.n57 24.5923
R109 VP.n59 VP.n58 24.5923
R110 VP.n39 VP.n38 24.5923
R111 VP.n40 VP.n39 24.5923
R112 VP.n40 VP.n25 24.5923
R113 VP.n44 VP.n25 24.5923
R114 VP.n45 VP.n44 24.5923
R115 VP.n46 VP.n45 24.5923
R116 VP.n33 VP.n32 24.5923
R117 VP.n34 VP.n33 24.5923
R118 VP.n83 VP.n12 18.6903
R119 VP.n104 VP.n103 18.6903
R120 VP.n53 VP.n52 18.6903
R121 VP.n32 VP.n29 18.6903
R122 VP.n68 VP.n16 12.7883
R123 VP.n116 VP.n0 12.7883
R124 VP.n65 VP.n17 12.7883
R125 VP.n80 VP.n12 5.90254
R126 VP.n103 VP.n4 5.90254
R127 VP.n52 VP.n21 5.90254
R128 VP.n31 VP.n30 3.05548
R129 VP.n67 VP.n66 0.354861
R130 VP.n70 VP.n69 0.354861
R131 VP.n118 VP.n117 0.354861
R132 VP VP.n118 0.267071
R133 VP.n31 VP.n28 0.189894
R134 VP.n35 VP.n28 0.189894
R135 VP.n36 VP.n35 0.189894
R136 VP.n37 VP.n36 0.189894
R137 VP.n37 VP.n26 0.189894
R138 VP.n41 VP.n26 0.189894
R139 VP.n42 VP.n41 0.189894
R140 VP.n43 VP.n42 0.189894
R141 VP.n43 VP.n24 0.189894
R142 VP.n47 VP.n24 0.189894
R143 VP.n48 VP.n47 0.189894
R144 VP.n49 VP.n48 0.189894
R145 VP.n49 VP.n22 0.189894
R146 VP.n54 VP.n22 0.189894
R147 VP.n55 VP.n54 0.189894
R148 VP.n56 VP.n55 0.189894
R149 VP.n56 VP.n20 0.189894
R150 VP.n60 VP.n20 0.189894
R151 VP.n61 VP.n60 0.189894
R152 VP.n62 VP.n61 0.189894
R153 VP.n62 VP.n18 0.189894
R154 VP.n66 VP.n18 0.189894
R155 VP.n71 VP.n70 0.189894
R156 VP.n71 VP.n15 0.189894
R157 VP.n75 VP.n15 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n77 VP.n76 0.189894
R160 VP.n77 VP.n13 0.189894
R161 VP.n81 VP.n13 0.189894
R162 VP.n82 VP.n81 0.189894
R163 VP.n82 VP.n11 0.189894
R164 VP.n86 VP.n11 0.189894
R165 VP.n87 VP.n86 0.189894
R166 VP.n88 VP.n87 0.189894
R167 VP.n88 VP.n9 0.189894
R168 VP.n92 VP.n9 0.189894
R169 VP.n93 VP.n92 0.189894
R170 VP.n94 VP.n93 0.189894
R171 VP.n94 VP.n7 0.189894
R172 VP.n98 VP.n7 0.189894
R173 VP.n99 VP.n98 0.189894
R174 VP.n100 VP.n99 0.189894
R175 VP.n100 VP.n5 0.189894
R176 VP.n105 VP.n5 0.189894
R177 VP.n106 VP.n105 0.189894
R178 VP.n107 VP.n106 0.189894
R179 VP.n107 VP.n3 0.189894
R180 VP.n111 VP.n3 0.189894
R181 VP.n112 VP.n111 0.189894
R182 VP.n113 VP.n112 0.189894
R183 VP.n113 VP.n1 0.189894
R184 VP.n117 VP.n1 0.189894
R185 VTAIL.n320 VTAIL.n248 289.615
R186 VTAIL.n74 VTAIL.n2 289.615
R187 VTAIL.n242 VTAIL.n170 289.615
R188 VTAIL.n160 VTAIL.n88 289.615
R189 VTAIL.n272 VTAIL.n271 185
R190 VTAIL.n277 VTAIL.n276 185
R191 VTAIL.n279 VTAIL.n278 185
R192 VTAIL.n268 VTAIL.n267 185
R193 VTAIL.n285 VTAIL.n284 185
R194 VTAIL.n287 VTAIL.n286 185
R195 VTAIL.n264 VTAIL.n263 185
R196 VTAIL.n294 VTAIL.n293 185
R197 VTAIL.n295 VTAIL.n262 185
R198 VTAIL.n297 VTAIL.n296 185
R199 VTAIL.n260 VTAIL.n259 185
R200 VTAIL.n303 VTAIL.n302 185
R201 VTAIL.n305 VTAIL.n304 185
R202 VTAIL.n256 VTAIL.n255 185
R203 VTAIL.n311 VTAIL.n310 185
R204 VTAIL.n313 VTAIL.n312 185
R205 VTAIL.n252 VTAIL.n251 185
R206 VTAIL.n319 VTAIL.n318 185
R207 VTAIL.n321 VTAIL.n320 185
R208 VTAIL.n26 VTAIL.n25 185
R209 VTAIL.n31 VTAIL.n30 185
R210 VTAIL.n33 VTAIL.n32 185
R211 VTAIL.n22 VTAIL.n21 185
R212 VTAIL.n39 VTAIL.n38 185
R213 VTAIL.n41 VTAIL.n40 185
R214 VTAIL.n18 VTAIL.n17 185
R215 VTAIL.n48 VTAIL.n47 185
R216 VTAIL.n49 VTAIL.n16 185
R217 VTAIL.n51 VTAIL.n50 185
R218 VTAIL.n14 VTAIL.n13 185
R219 VTAIL.n57 VTAIL.n56 185
R220 VTAIL.n59 VTAIL.n58 185
R221 VTAIL.n10 VTAIL.n9 185
R222 VTAIL.n65 VTAIL.n64 185
R223 VTAIL.n67 VTAIL.n66 185
R224 VTAIL.n6 VTAIL.n5 185
R225 VTAIL.n73 VTAIL.n72 185
R226 VTAIL.n75 VTAIL.n74 185
R227 VTAIL.n243 VTAIL.n242 185
R228 VTAIL.n241 VTAIL.n240 185
R229 VTAIL.n174 VTAIL.n173 185
R230 VTAIL.n235 VTAIL.n234 185
R231 VTAIL.n233 VTAIL.n232 185
R232 VTAIL.n178 VTAIL.n177 185
R233 VTAIL.n227 VTAIL.n226 185
R234 VTAIL.n225 VTAIL.n224 185
R235 VTAIL.n182 VTAIL.n181 185
R236 VTAIL.n219 VTAIL.n218 185
R237 VTAIL.n217 VTAIL.n184 185
R238 VTAIL.n216 VTAIL.n215 185
R239 VTAIL.n187 VTAIL.n185 185
R240 VTAIL.n210 VTAIL.n209 185
R241 VTAIL.n208 VTAIL.n207 185
R242 VTAIL.n191 VTAIL.n190 185
R243 VTAIL.n202 VTAIL.n201 185
R244 VTAIL.n200 VTAIL.n199 185
R245 VTAIL.n195 VTAIL.n194 185
R246 VTAIL.n161 VTAIL.n160 185
R247 VTAIL.n159 VTAIL.n158 185
R248 VTAIL.n92 VTAIL.n91 185
R249 VTAIL.n153 VTAIL.n152 185
R250 VTAIL.n151 VTAIL.n150 185
R251 VTAIL.n96 VTAIL.n95 185
R252 VTAIL.n145 VTAIL.n144 185
R253 VTAIL.n143 VTAIL.n142 185
R254 VTAIL.n100 VTAIL.n99 185
R255 VTAIL.n137 VTAIL.n136 185
R256 VTAIL.n135 VTAIL.n102 185
R257 VTAIL.n134 VTAIL.n133 185
R258 VTAIL.n105 VTAIL.n103 185
R259 VTAIL.n128 VTAIL.n127 185
R260 VTAIL.n126 VTAIL.n125 185
R261 VTAIL.n109 VTAIL.n108 185
R262 VTAIL.n120 VTAIL.n119 185
R263 VTAIL.n118 VTAIL.n117 185
R264 VTAIL.n113 VTAIL.n112 185
R265 VTAIL.n273 VTAIL.t0 149.524
R266 VTAIL.n27 VTAIL.t19 149.524
R267 VTAIL.n196 VTAIL.t12 149.524
R268 VTAIL.n114 VTAIL.t6 149.524
R269 VTAIL.n277 VTAIL.n271 104.615
R270 VTAIL.n278 VTAIL.n277 104.615
R271 VTAIL.n278 VTAIL.n267 104.615
R272 VTAIL.n285 VTAIL.n267 104.615
R273 VTAIL.n286 VTAIL.n285 104.615
R274 VTAIL.n286 VTAIL.n263 104.615
R275 VTAIL.n294 VTAIL.n263 104.615
R276 VTAIL.n295 VTAIL.n294 104.615
R277 VTAIL.n296 VTAIL.n295 104.615
R278 VTAIL.n296 VTAIL.n259 104.615
R279 VTAIL.n303 VTAIL.n259 104.615
R280 VTAIL.n304 VTAIL.n303 104.615
R281 VTAIL.n304 VTAIL.n255 104.615
R282 VTAIL.n311 VTAIL.n255 104.615
R283 VTAIL.n312 VTAIL.n311 104.615
R284 VTAIL.n312 VTAIL.n251 104.615
R285 VTAIL.n319 VTAIL.n251 104.615
R286 VTAIL.n320 VTAIL.n319 104.615
R287 VTAIL.n31 VTAIL.n25 104.615
R288 VTAIL.n32 VTAIL.n31 104.615
R289 VTAIL.n32 VTAIL.n21 104.615
R290 VTAIL.n39 VTAIL.n21 104.615
R291 VTAIL.n40 VTAIL.n39 104.615
R292 VTAIL.n40 VTAIL.n17 104.615
R293 VTAIL.n48 VTAIL.n17 104.615
R294 VTAIL.n49 VTAIL.n48 104.615
R295 VTAIL.n50 VTAIL.n49 104.615
R296 VTAIL.n50 VTAIL.n13 104.615
R297 VTAIL.n57 VTAIL.n13 104.615
R298 VTAIL.n58 VTAIL.n57 104.615
R299 VTAIL.n58 VTAIL.n9 104.615
R300 VTAIL.n65 VTAIL.n9 104.615
R301 VTAIL.n66 VTAIL.n65 104.615
R302 VTAIL.n66 VTAIL.n5 104.615
R303 VTAIL.n73 VTAIL.n5 104.615
R304 VTAIL.n74 VTAIL.n73 104.615
R305 VTAIL.n242 VTAIL.n241 104.615
R306 VTAIL.n241 VTAIL.n173 104.615
R307 VTAIL.n234 VTAIL.n173 104.615
R308 VTAIL.n234 VTAIL.n233 104.615
R309 VTAIL.n233 VTAIL.n177 104.615
R310 VTAIL.n226 VTAIL.n177 104.615
R311 VTAIL.n226 VTAIL.n225 104.615
R312 VTAIL.n225 VTAIL.n181 104.615
R313 VTAIL.n218 VTAIL.n181 104.615
R314 VTAIL.n218 VTAIL.n217 104.615
R315 VTAIL.n217 VTAIL.n216 104.615
R316 VTAIL.n216 VTAIL.n185 104.615
R317 VTAIL.n209 VTAIL.n185 104.615
R318 VTAIL.n209 VTAIL.n208 104.615
R319 VTAIL.n208 VTAIL.n190 104.615
R320 VTAIL.n201 VTAIL.n190 104.615
R321 VTAIL.n201 VTAIL.n200 104.615
R322 VTAIL.n200 VTAIL.n194 104.615
R323 VTAIL.n160 VTAIL.n159 104.615
R324 VTAIL.n159 VTAIL.n91 104.615
R325 VTAIL.n152 VTAIL.n91 104.615
R326 VTAIL.n152 VTAIL.n151 104.615
R327 VTAIL.n151 VTAIL.n95 104.615
R328 VTAIL.n144 VTAIL.n95 104.615
R329 VTAIL.n144 VTAIL.n143 104.615
R330 VTAIL.n143 VTAIL.n99 104.615
R331 VTAIL.n136 VTAIL.n99 104.615
R332 VTAIL.n136 VTAIL.n135 104.615
R333 VTAIL.n135 VTAIL.n134 104.615
R334 VTAIL.n134 VTAIL.n103 104.615
R335 VTAIL.n127 VTAIL.n103 104.615
R336 VTAIL.n127 VTAIL.n126 104.615
R337 VTAIL.n126 VTAIL.n108 104.615
R338 VTAIL.n119 VTAIL.n108 104.615
R339 VTAIL.n119 VTAIL.n118 104.615
R340 VTAIL.n118 VTAIL.n112 104.615
R341 VTAIL.t0 VTAIL.n271 52.3082
R342 VTAIL.t19 VTAIL.n25 52.3082
R343 VTAIL.t12 VTAIL.n194 52.3082
R344 VTAIL.t6 VTAIL.n112 52.3082
R345 VTAIL.n169 VTAIL.n168 43.1979
R346 VTAIL.n167 VTAIL.n166 43.1979
R347 VTAIL.n87 VTAIL.n86 43.1979
R348 VTAIL.n85 VTAIL.n84 43.1979
R349 VTAIL.n327 VTAIL.n326 43.1979
R350 VTAIL.n1 VTAIL.n0 43.1979
R351 VTAIL.n81 VTAIL.n80 43.1979
R352 VTAIL.n83 VTAIL.n82 43.1979
R353 VTAIL.n85 VTAIL.n83 31.2979
R354 VTAIL.n325 VTAIL.n324 30.6338
R355 VTAIL.n79 VTAIL.n78 30.6338
R356 VTAIL.n247 VTAIL.n246 30.6338
R357 VTAIL.n165 VTAIL.n164 30.6338
R358 VTAIL.n325 VTAIL.n247 27.9531
R359 VTAIL.n297 VTAIL.n262 13.1884
R360 VTAIL.n51 VTAIL.n16 13.1884
R361 VTAIL.n219 VTAIL.n184 13.1884
R362 VTAIL.n137 VTAIL.n102 13.1884
R363 VTAIL.n293 VTAIL.n292 12.8005
R364 VTAIL.n298 VTAIL.n260 12.8005
R365 VTAIL.n47 VTAIL.n46 12.8005
R366 VTAIL.n52 VTAIL.n14 12.8005
R367 VTAIL.n220 VTAIL.n182 12.8005
R368 VTAIL.n215 VTAIL.n186 12.8005
R369 VTAIL.n138 VTAIL.n100 12.8005
R370 VTAIL.n133 VTAIL.n104 12.8005
R371 VTAIL.n291 VTAIL.n264 12.0247
R372 VTAIL.n302 VTAIL.n301 12.0247
R373 VTAIL.n45 VTAIL.n18 12.0247
R374 VTAIL.n56 VTAIL.n55 12.0247
R375 VTAIL.n224 VTAIL.n223 12.0247
R376 VTAIL.n214 VTAIL.n187 12.0247
R377 VTAIL.n142 VTAIL.n141 12.0247
R378 VTAIL.n132 VTAIL.n105 12.0247
R379 VTAIL.n288 VTAIL.n287 11.249
R380 VTAIL.n305 VTAIL.n258 11.249
R381 VTAIL.n42 VTAIL.n41 11.249
R382 VTAIL.n59 VTAIL.n12 11.249
R383 VTAIL.n227 VTAIL.n180 11.249
R384 VTAIL.n211 VTAIL.n210 11.249
R385 VTAIL.n145 VTAIL.n98 11.249
R386 VTAIL.n129 VTAIL.n128 11.249
R387 VTAIL.n284 VTAIL.n266 10.4732
R388 VTAIL.n306 VTAIL.n256 10.4732
R389 VTAIL.n38 VTAIL.n20 10.4732
R390 VTAIL.n60 VTAIL.n10 10.4732
R391 VTAIL.n228 VTAIL.n178 10.4732
R392 VTAIL.n207 VTAIL.n189 10.4732
R393 VTAIL.n146 VTAIL.n96 10.4732
R394 VTAIL.n125 VTAIL.n107 10.4732
R395 VTAIL.n273 VTAIL.n272 10.2747
R396 VTAIL.n27 VTAIL.n26 10.2747
R397 VTAIL.n196 VTAIL.n195 10.2747
R398 VTAIL.n114 VTAIL.n113 10.2747
R399 VTAIL.n283 VTAIL.n268 9.69747
R400 VTAIL.n310 VTAIL.n309 9.69747
R401 VTAIL.n37 VTAIL.n22 9.69747
R402 VTAIL.n64 VTAIL.n63 9.69747
R403 VTAIL.n232 VTAIL.n231 9.69747
R404 VTAIL.n206 VTAIL.n191 9.69747
R405 VTAIL.n150 VTAIL.n149 9.69747
R406 VTAIL.n124 VTAIL.n109 9.69747
R407 VTAIL.n324 VTAIL.n323 9.45567
R408 VTAIL.n78 VTAIL.n77 9.45567
R409 VTAIL.n246 VTAIL.n245 9.45567
R410 VTAIL.n164 VTAIL.n163 9.45567
R411 VTAIL.n250 VTAIL.n249 9.3005
R412 VTAIL.n323 VTAIL.n322 9.3005
R413 VTAIL.n315 VTAIL.n314 9.3005
R414 VTAIL.n254 VTAIL.n253 9.3005
R415 VTAIL.n309 VTAIL.n308 9.3005
R416 VTAIL.n307 VTAIL.n306 9.3005
R417 VTAIL.n258 VTAIL.n257 9.3005
R418 VTAIL.n301 VTAIL.n300 9.3005
R419 VTAIL.n299 VTAIL.n298 9.3005
R420 VTAIL.n275 VTAIL.n274 9.3005
R421 VTAIL.n270 VTAIL.n269 9.3005
R422 VTAIL.n281 VTAIL.n280 9.3005
R423 VTAIL.n283 VTAIL.n282 9.3005
R424 VTAIL.n266 VTAIL.n265 9.3005
R425 VTAIL.n289 VTAIL.n288 9.3005
R426 VTAIL.n291 VTAIL.n290 9.3005
R427 VTAIL.n292 VTAIL.n261 9.3005
R428 VTAIL.n317 VTAIL.n316 9.3005
R429 VTAIL.n4 VTAIL.n3 9.3005
R430 VTAIL.n77 VTAIL.n76 9.3005
R431 VTAIL.n69 VTAIL.n68 9.3005
R432 VTAIL.n8 VTAIL.n7 9.3005
R433 VTAIL.n63 VTAIL.n62 9.3005
R434 VTAIL.n61 VTAIL.n60 9.3005
R435 VTAIL.n12 VTAIL.n11 9.3005
R436 VTAIL.n55 VTAIL.n54 9.3005
R437 VTAIL.n53 VTAIL.n52 9.3005
R438 VTAIL.n29 VTAIL.n28 9.3005
R439 VTAIL.n24 VTAIL.n23 9.3005
R440 VTAIL.n35 VTAIL.n34 9.3005
R441 VTAIL.n37 VTAIL.n36 9.3005
R442 VTAIL.n20 VTAIL.n19 9.3005
R443 VTAIL.n43 VTAIL.n42 9.3005
R444 VTAIL.n45 VTAIL.n44 9.3005
R445 VTAIL.n46 VTAIL.n15 9.3005
R446 VTAIL.n71 VTAIL.n70 9.3005
R447 VTAIL.n172 VTAIL.n171 9.3005
R448 VTAIL.n239 VTAIL.n238 9.3005
R449 VTAIL.n237 VTAIL.n236 9.3005
R450 VTAIL.n176 VTAIL.n175 9.3005
R451 VTAIL.n231 VTAIL.n230 9.3005
R452 VTAIL.n229 VTAIL.n228 9.3005
R453 VTAIL.n180 VTAIL.n179 9.3005
R454 VTAIL.n223 VTAIL.n222 9.3005
R455 VTAIL.n221 VTAIL.n220 9.3005
R456 VTAIL.n186 VTAIL.n183 9.3005
R457 VTAIL.n214 VTAIL.n213 9.3005
R458 VTAIL.n212 VTAIL.n211 9.3005
R459 VTAIL.n189 VTAIL.n188 9.3005
R460 VTAIL.n206 VTAIL.n205 9.3005
R461 VTAIL.n204 VTAIL.n203 9.3005
R462 VTAIL.n193 VTAIL.n192 9.3005
R463 VTAIL.n198 VTAIL.n197 9.3005
R464 VTAIL.n245 VTAIL.n244 9.3005
R465 VTAIL.n116 VTAIL.n115 9.3005
R466 VTAIL.n111 VTAIL.n110 9.3005
R467 VTAIL.n122 VTAIL.n121 9.3005
R468 VTAIL.n124 VTAIL.n123 9.3005
R469 VTAIL.n107 VTAIL.n106 9.3005
R470 VTAIL.n130 VTAIL.n129 9.3005
R471 VTAIL.n132 VTAIL.n131 9.3005
R472 VTAIL.n104 VTAIL.n101 9.3005
R473 VTAIL.n163 VTAIL.n162 9.3005
R474 VTAIL.n90 VTAIL.n89 9.3005
R475 VTAIL.n157 VTAIL.n156 9.3005
R476 VTAIL.n155 VTAIL.n154 9.3005
R477 VTAIL.n94 VTAIL.n93 9.3005
R478 VTAIL.n149 VTAIL.n148 9.3005
R479 VTAIL.n147 VTAIL.n146 9.3005
R480 VTAIL.n98 VTAIL.n97 9.3005
R481 VTAIL.n141 VTAIL.n140 9.3005
R482 VTAIL.n139 VTAIL.n138 9.3005
R483 VTAIL.n280 VTAIL.n279 8.92171
R484 VTAIL.n313 VTAIL.n254 8.92171
R485 VTAIL.n34 VTAIL.n33 8.92171
R486 VTAIL.n67 VTAIL.n8 8.92171
R487 VTAIL.n235 VTAIL.n176 8.92171
R488 VTAIL.n203 VTAIL.n202 8.92171
R489 VTAIL.n153 VTAIL.n94 8.92171
R490 VTAIL.n121 VTAIL.n120 8.92171
R491 VTAIL.n276 VTAIL.n270 8.14595
R492 VTAIL.n314 VTAIL.n252 8.14595
R493 VTAIL.n324 VTAIL.n248 8.14595
R494 VTAIL.n30 VTAIL.n24 8.14595
R495 VTAIL.n68 VTAIL.n6 8.14595
R496 VTAIL.n78 VTAIL.n2 8.14595
R497 VTAIL.n246 VTAIL.n170 8.14595
R498 VTAIL.n236 VTAIL.n174 8.14595
R499 VTAIL.n199 VTAIL.n193 8.14595
R500 VTAIL.n164 VTAIL.n88 8.14595
R501 VTAIL.n154 VTAIL.n92 8.14595
R502 VTAIL.n117 VTAIL.n111 8.14595
R503 VTAIL.n275 VTAIL.n272 7.3702
R504 VTAIL.n318 VTAIL.n317 7.3702
R505 VTAIL.n322 VTAIL.n321 7.3702
R506 VTAIL.n29 VTAIL.n26 7.3702
R507 VTAIL.n72 VTAIL.n71 7.3702
R508 VTAIL.n76 VTAIL.n75 7.3702
R509 VTAIL.n244 VTAIL.n243 7.3702
R510 VTAIL.n240 VTAIL.n239 7.3702
R511 VTAIL.n198 VTAIL.n195 7.3702
R512 VTAIL.n162 VTAIL.n161 7.3702
R513 VTAIL.n158 VTAIL.n157 7.3702
R514 VTAIL.n116 VTAIL.n113 7.3702
R515 VTAIL.n318 VTAIL.n250 6.59444
R516 VTAIL.n321 VTAIL.n250 6.59444
R517 VTAIL.n72 VTAIL.n4 6.59444
R518 VTAIL.n75 VTAIL.n4 6.59444
R519 VTAIL.n243 VTAIL.n172 6.59444
R520 VTAIL.n240 VTAIL.n172 6.59444
R521 VTAIL.n161 VTAIL.n90 6.59444
R522 VTAIL.n158 VTAIL.n90 6.59444
R523 VTAIL.n276 VTAIL.n275 5.81868
R524 VTAIL.n317 VTAIL.n252 5.81868
R525 VTAIL.n322 VTAIL.n248 5.81868
R526 VTAIL.n30 VTAIL.n29 5.81868
R527 VTAIL.n71 VTAIL.n6 5.81868
R528 VTAIL.n76 VTAIL.n2 5.81868
R529 VTAIL.n244 VTAIL.n170 5.81868
R530 VTAIL.n239 VTAIL.n174 5.81868
R531 VTAIL.n199 VTAIL.n198 5.81868
R532 VTAIL.n162 VTAIL.n88 5.81868
R533 VTAIL.n157 VTAIL.n92 5.81868
R534 VTAIL.n117 VTAIL.n116 5.81868
R535 VTAIL.n279 VTAIL.n270 5.04292
R536 VTAIL.n314 VTAIL.n313 5.04292
R537 VTAIL.n33 VTAIL.n24 5.04292
R538 VTAIL.n68 VTAIL.n67 5.04292
R539 VTAIL.n236 VTAIL.n235 5.04292
R540 VTAIL.n202 VTAIL.n193 5.04292
R541 VTAIL.n154 VTAIL.n153 5.04292
R542 VTAIL.n120 VTAIL.n111 5.04292
R543 VTAIL.n280 VTAIL.n268 4.26717
R544 VTAIL.n310 VTAIL.n254 4.26717
R545 VTAIL.n34 VTAIL.n22 4.26717
R546 VTAIL.n64 VTAIL.n8 4.26717
R547 VTAIL.n232 VTAIL.n176 4.26717
R548 VTAIL.n203 VTAIL.n191 4.26717
R549 VTAIL.n150 VTAIL.n94 4.26717
R550 VTAIL.n121 VTAIL.n109 4.26717
R551 VTAIL.n284 VTAIL.n283 3.49141
R552 VTAIL.n309 VTAIL.n256 3.49141
R553 VTAIL.n38 VTAIL.n37 3.49141
R554 VTAIL.n63 VTAIL.n10 3.49141
R555 VTAIL.n231 VTAIL.n178 3.49141
R556 VTAIL.n207 VTAIL.n206 3.49141
R557 VTAIL.n149 VTAIL.n96 3.49141
R558 VTAIL.n125 VTAIL.n124 3.49141
R559 VTAIL.n87 VTAIL.n85 3.34533
R560 VTAIL.n165 VTAIL.n87 3.34533
R561 VTAIL.n169 VTAIL.n167 3.34533
R562 VTAIL.n247 VTAIL.n169 3.34533
R563 VTAIL.n83 VTAIL.n81 3.34533
R564 VTAIL.n81 VTAIL.n79 3.34533
R565 VTAIL.n327 VTAIL.n325 3.34533
R566 VTAIL.n274 VTAIL.n273 2.84303
R567 VTAIL.n28 VTAIL.n27 2.84303
R568 VTAIL.n115 VTAIL.n114 2.84303
R569 VTAIL.n197 VTAIL.n196 2.84303
R570 VTAIL.n287 VTAIL.n266 2.71565
R571 VTAIL.n306 VTAIL.n305 2.71565
R572 VTAIL.n41 VTAIL.n20 2.71565
R573 VTAIL.n60 VTAIL.n59 2.71565
R574 VTAIL.n228 VTAIL.n227 2.71565
R575 VTAIL.n210 VTAIL.n189 2.71565
R576 VTAIL.n146 VTAIL.n145 2.71565
R577 VTAIL.n128 VTAIL.n107 2.71565
R578 VTAIL VTAIL.n1 2.56731
R579 VTAIL.n167 VTAIL.n165 2.14274
R580 VTAIL.n79 VTAIL.n1 2.14274
R581 VTAIL.n288 VTAIL.n264 1.93989
R582 VTAIL.n302 VTAIL.n258 1.93989
R583 VTAIL.n42 VTAIL.n18 1.93989
R584 VTAIL.n56 VTAIL.n12 1.93989
R585 VTAIL.n224 VTAIL.n180 1.93989
R586 VTAIL.n211 VTAIL.n187 1.93989
R587 VTAIL.n142 VTAIL.n98 1.93989
R588 VTAIL.n129 VTAIL.n105 1.93989
R589 VTAIL.n326 VTAIL.t9 1.39487
R590 VTAIL.n326 VTAIL.t7 1.39487
R591 VTAIL.n0 VTAIL.t2 1.39487
R592 VTAIL.n0 VTAIL.t5 1.39487
R593 VTAIL.n80 VTAIL.t14 1.39487
R594 VTAIL.n80 VTAIL.t18 1.39487
R595 VTAIL.n82 VTAIL.t16 1.39487
R596 VTAIL.n82 VTAIL.t15 1.39487
R597 VTAIL.n168 VTAIL.t10 1.39487
R598 VTAIL.n168 VTAIL.t17 1.39487
R599 VTAIL.n166 VTAIL.t13 1.39487
R600 VTAIL.n166 VTAIL.t11 1.39487
R601 VTAIL.n86 VTAIL.t3 1.39487
R602 VTAIL.n86 VTAIL.t1 1.39487
R603 VTAIL.n84 VTAIL.t8 1.39487
R604 VTAIL.n84 VTAIL.t4 1.39487
R605 VTAIL.n293 VTAIL.n291 1.16414
R606 VTAIL.n301 VTAIL.n260 1.16414
R607 VTAIL.n47 VTAIL.n45 1.16414
R608 VTAIL.n55 VTAIL.n14 1.16414
R609 VTAIL.n223 VTAIL.n182 1.16414
R610 VTAIL.n215 VTAIL.n214 1.16414
R611 VTAIL.n141 VTAIL.n100 1.16414
R612 VTAIL.n133 VTAIL.n132 1.16414
R613 VTAIL VTAIL.n327 0.778517
R614 VTAIL.n292 VTAIL.n262 0.388379
R615 VTAIL.n298 VTAIL.n297 0.388379
R616 VTAIL.n46 VTAIL.n16 0.388379
R617 VTAIL.n52 VTAIL.n51 0.388379
R618 VTAIL.n220 VTAIL.n219 0.388379
R619 VTAIL.n186 VTAIL.n184 0.388379
R620 VTAIL.n138 VTAIL.n137 0.388379
R621 VTAIL.n104 VTAIL.n102 0.388379
R622 VTAIL.n274 VTAIL.n269 0.155672
R623 VTAIL.n281 VTAIL.n269 0.155672
R624 VTAIL.n282 VTAIL.n281 0.155672
R625 VTAIL.n282 VTAIL.n265 0.155672
R626 VTAIL.n289 VTAIL.n265 0.155672
R627 VTAIL.n290 VTAIL.n289 0.155672
R628 VTAIL.n290 VTAIL.n261 0.155672
R629 VTAIL.n299 VTAIL.n261 0.155672
R630 VTAIL.n300 VTAIL.n299 0.155672
R631 VTAIL.n300 VTAIL.n257 0.155672
R632 VTAIL.n307 VTAIL.n257 0.155672
R633 VTAIL.n308 VTAIL.n307 0.155672
R634 VTAIL.n308 VTAIL.n253 0.155672
R635 VTAIL.n315 VTAIL.n253 0.155672
R636 VTAIL.n316 VTAIL.n315 0.155672
R637 VTAIL.n316 VTAIL.n249 0.155672
R638 VTAIL.n323 VTAIL.n249 0.155672
R639 VTAIL.n28 VTAIL.n23 0.155672
R640 VTAIL.n35 VTAIL.n23 0.155672
R641 VTAIL.n36 VTAIL.n35 0.155672
R642 VTAIL.n36 VTAIL.n19 0.155672
R643 VTAIL.n43 VTAIL.n19 0.155672
R644 VTAIL.n44 VTAIL.n43 0.155672
R645 VTAIL.n44 VTAIL.n15 0.155672
R646 VTAIL.n53 VTAIL.n15 0.155672
R647 VTAIL.n54 VTAIL.n53 0.155672
R648 VTAIL.n54 VTAIL.n11 0.155672
R649 VTAIL.n61 VTAIL.n11 0.155672
R650 VTAIL.n62 VTAIL.n61 0.155672
R651 VTAIL.n62 VTAIL.n7 0.155672
R652 VTAIL.n69 VTAIL.n7 0.155672
R653 VTAIL.n70 VTAIL.n69 0.155672
R654 VTAIL.n70 VTAIL.n3 0.155672
R655 VTAIL.n77 VTAIL.n3 0.155672
R656 VTAIL.n245 VTAIL.n171 0.155672
R657 VTAIL.n238 VTAIL.n171 0.155672
R658 VTAIL.n238 VTAIL.n237 0.155672
R659 VTAIL.n237 VTAIL.n175 0.155672
R660 VTAIL.n230 VTAIL.n175 0.155672
R661 VTAIL.n230 VTAIL.n229 0.155672
R662 VTAIL.n229 VTAIL.n179 0.155672
R663 VTAIL.n222 VTAIL.n179 0.155672
R664 VTAIL.n222 VTAIL.n221 0.155672
R665 VTAIL.n221 VTAIL.n183 0.155672
R666 VTAIL.n213 VTAIL.n183 0.155672
R667 VTAIL.n213 VTAIL.n212 0.155672
R668 VTAIL.n212 VTAIL.n188 0.155672
R669 VTAIL.n205 VTAIL.n188 0.155672
R670 VTAIL.n205 VTAIL.n204 0.155672
R671 VTAIL.n204 VTAIL.n192 0.155672
R672 VTAIL.n197 VTAIL.n192 0.155672
R673 VTAIL.n163 VTAIL.n89 0.155672
R674 VTAIL.n156 VTAIL.n89 0.155672
R675 VTAIL.n156 VTAIL.n155 0.155672
R676 VTAIL.n155 VTAIL.n93 0.155672
R677 VTAIL.n148 VTAIL.n93 0.155672
R678 VTAIL.n148 VTAIL.n147 0.155672
R679 VTAIL.n147 VTAIL.n97 0.155672
R680 VTAIL.n140 VTAIL.n97 0.155672
R681 VTAIL.n140 VTAIL.n139 0.155672
R682 VTAIL.n139 VTAIL.n101 0.155672
R683 VTAIL.n131 VTAIL.n101 0.155672
R684 VTAIL.n131 VTAIL.n130 0.155672
R685 VTAIL.n130 VTAIL.n106 0.155672
R686 VTAIL.n123 VTAIL.n106 0.155672
R687 VTAIL.n123 VTAIL.n122 0.155672
R688 VTAIL.n122 VTAIL.n110 0.155672
R689 VTAIL.n115 VTAIL.n110 0.155672
R690 VDD1.n72 VDD1.n0 289.615
R691 VDD1.n151 VDD1.n79 289.615
R692 VDD1.n73 VDD1.n72 185
R693 VDD1.n71 VDD1.n70 185
R694 VDD1.n4 VDD1.n3 185
R695 VDD1.n65 VDD1.n64 185
R696 VDD1.n63 VDD1.n62 185
R697 VDD1.n8 VDD1.n7 185
R698 VDD1.n57 VDD1.n56 185
R699 VDD1.n55 VDD1.n54 185
R700 VDD1.n12 VDD1.n11 185
R701 VDD1.n49 VDD1.n48 185
R702 VDD1.n47 VDD1.n14 185
R703 VDD1.n46 VDD1.n45 185
R704 VDD1.n17 VDD1.n15 185
R705 VDD1.n40 VDD1.n39 185
R706 VDD1.n38 VDD1.n37 185
R707 VDD1.n21 VDD1.n20 185
R708 VDD1.n32 VDD1.n31 185
R709 VDD1.n30 VDD1.n29 185
R710 VDD1.n25 VDD1.n24 185
R711 VDD1.n103 VDD1.n102 185
R712 VDD1.n108 VDD1.n107 185
R713 VDD1.n110 VDD1.n109 185
R714 VDD1.n99 VDD1.n98 185
R715 VDD1.n116 VDD1.n115 185
R716 VDD1.n118 VDD1.n117 185
R717 VDD1.n95 VDD1.n94 185
R718 VDD1.n125 VDD1.n124 185
R719 VDD1.n126 VDD1.n93 185
R720 VDD1.n128 VDD1.n127 185
R721 VDD1.n91 VDD1.n90 185
R722 VDD1.n134 VDD1.n133 185
R723 VDD1.n136 VDD1.n135 185
R724 VDD1.n87 VDD1.n86 185
R725 VDD1.n142 VDD1.n141 185
R726 VDD1.n144 VDD1.n143 185
R727 VDD1.n83 VDD1.n82 185
R728 VDD1.n150 VDD1.n149 185
R729 VDD1.n152 VDD1.n151 185
R730 VDD1.n26 VDD1.t8 149.524
R731 VDD1.n104 VDD1.t1 149.524
R732 VDD1.n72 VDD1.n71 104.615
R733 VDD1.n71 VDD1.n3 104.615
R734 VDD1.n64 VDD1.n3 104.615
R735 VDD1.n64 VDD1.n63 104.615
R736 VDD1.n63 VDD1.n7 104.615
R737 VDD1.n56 VDD1.n7 104.615
R738 VDD1.n56 VDD1.n55 104.615
R739 VDD1.n55 VDD1.n11 104.615
R740 VDD1.n48 VDD1.n11 104.615
R741 VDD1.n48 VDD1.n47 104.615
R742 VDD1.n47 VDD1.n46 104.615
R743 VDD1.n46 VDD1.n15 104.615
R744 VDD1.n39 VDD1.n15 104.615
R745 VDD1.n39 VDD1.n38 104.615
R746 VDD1.n38 VDD1.n20 104.615
R747 VDD1.n31 VDD1.n20 104.615
R748 VDD1.n31 VDD1.n30 104.615
R749 VDD1.n30 VDD1.n24 104.615
R750 VDD1.n108 VDD1.n102 104.615
R751 VDD1.n109 VDD1.n108 104.615
R752 VDD1.n109 VDD1.n98 104.615
R753 VDD1.n116 VDD1.n98 104.615
R754 VDD1.n117 VDD1.n116 104.615
R755 VDD1.n117 VDD1.n94 104.615
R756 VDD1.n125 VDD1.n94 104.615
R757 VDD1.n126 VDD1.n125 104.615
R758 VDD1.n127 VDD1.n126 104.615
R759 VDD1.n127 VDD1.n90 104.615
R760 VDD1.n134 VDD1.n90 104.615
R761 VDD1.n135 VDD1.n134 104.615
R762 VDD1.n135 VDD1.n86 104.615
R763 VDD1.n142 VDD1.n86 104.615
R764 VDD1.n143 VDD1.n142 104.615
R765 VDD1.n143 VDD1.n82 104.615
R766 VDD1.n150 VDD1.n82 104.615
R767 VDD1.n151 VDD1.n150 104.615
R768 VDD1.n159 VDD1.n158 62.3299
R769 VDD1.n161 VDD1.n160 59.8767
R770 VDD1.n78 VDD1.n77 59.8767
R771 VDD1.n157 VDD1.n156 59.8767
R772 VDD1.n161 VDD1.n159 54.1
R773 VDD1.t8 VDD1.n24 52.3082
R774 VDD1.t1 VDD1.n102 52.3082
R775 VDD1.n78 VDD1.n76 50.6574
R776 VDD1.n157 VDD1.n155 50.6574
R777 VDD1.n49 VDD1.n14 13.1884
R778 VDD1.n128 VDD1.n93 13.1884
R779 VDD1.n50 VDD1.n12 12.8005
R780 VDD1.n45 VDD1.n16 12.8005
R781 VDD1.n124 VDD1.n123 12.8005
R782 VDD1.n129 VDD1.n91 12.8005
R783 VDD1.n54 VDD1.n53 12.0247
R784 VDD1.n44 VDD1.n17 12.0247
R785 VDD1.n122 VDD1.n95 12.0247
R786 VDD1.n133 VDD1.n132 12.0247
R787 VDD1.n57 VDD1.n10 11.249
R788 VDD1.n41 VDD1.n40 11.249
R789 VDD1.n119 VDD1.n118 11.249
R790 VDD1.n136 VDD1.n89 11.249
R791 VDD1.n58 VDD1.n8 10.4732
R792 VDD1.n37 VDD1.n19 10.4732
R793 VDD1.n115 VDD1.n97 10.4732
R794 VDD1.n137 VDD1.n87 10.4732
R795 VDD1.n26 VDD1.n25 10.2747
R796 VDD1.n104 VDD1.n103 10.2747
R797 VDD1.n62 VDD1.n61 9.69747
R798 VDD1.n36 VDD1.n21 9.69747
R799 VDD1.n114 VDD1.n99 9.69747
R800 VDD1.n141 VDD1.n140 9.69747
R801 VDD1.n76 VDD1.n75 9.45567
R802 VDD1.n155 VDD1.n154 9.45567
R803 VDD1.n28 VDD1.n27 9.3005
R804 VDD1.n23 VDD1.n22 9.3005
R805 VDD1.n34 VDD1.n33 9.3005
R806 VDD1.n36 VDD1.n35 9.3005
R807 VDD1.n19 VDD1.n18 9.3005
R808 VDD1.n42 VDD1.n41 9.3005
R809 VDD1.n44 VDD1.n43 9.3005
R810 VDD1.n16 VDD1.n13 9.3005
R811 VDD1.n75 VDD1.n74 9.3005
R812 VDD1.n2 VDD1.n1 9.3005
R813 VDD1.n69 VDD1.n68 9.3005
R814 VDD1.n67 VDD1.n66 9.3005
R815 VDD1.n6 VDD1.n5 9.3005
R816 VDD1.n61 VDD1.n60 9.3005
R817 VDD1.n59 VDD1.n58 9.3005
R818 VDD1.n10 VDD1.n9 9.3005
R819 VDD1.n53 VDD1.n52 9.3005
R820 VDD1.n51 VDD1.n50 9.3005
R821 VDD1.n81 VDD1.n80 9.3005
R822 VDD1.n154 VDD1.n153 9.3005
R823 VDD1.n146 VDD1.n145 9.3005
R824 VDD1.n85 VDD1.n84 9.3005
R825 VDD1.n140 VDD1.n139 9.3005
R826 VDD1.n138 VDD1.n137 9.3005
R827 VDD1.n89 VDD1.n88 9.3005
R828 VDD1.n132 VDD1.n131 9.3005
R829 VDD1.n130 VDD1.n129 9.3005
R830 VDD1.n106 VDD1.n105 9.3005
R831 VDD1.n101 VDD1.n100 9.3005
R832 VDD1.n112 VDD1.n111 9.3005
R833 VDD1.n114 VDD1.n113 9.3005
R834 VDD1.n97 VDD1.n96 9.3005
R835 VDD1.n120 VDD1.n119 9.3005
R836 VDD1.n122 VDD1.n121 9.3005
R837 VDD1.n123 VDD1.n92 9.3005
R838 VDD1.n148 VDD1.n147 9.3005
R839 VDD1.n65 VDD1.n6 8.92171
R840 VDD1.n33 VDD1.n32 8.92171
R841 VDD1.n111 VDD1.n110 8.92171
R842 VDD1.n144 VDD1.n85 8.92171
R843 VDD1.n76 VDD1.n0 8.14595
R844 VDD1.n66 VDD1.n4 8.14595
R845 VDD1.n29 VDD1.n23 8.14595
R846 VDD1.n107 VDD1.n101 8.14595
R847 VDD1.n145 VDD1.n83 8.14595
R848 VDD1.n155 VDD1.n79 8.14595
R849 VDD1.n74 VDD1.n73 7.3702
R850 VDD1.n70 VDD1.n69 7.3702
R851 VDD1.n28 VDD1.n25 7.3702
R852 VDD1.n106 VDD1.n103 7.3702
R853 VDD1.n149 VDD1.n148 7.3702
R854 VDD1.n153 VDD1.n152 7.3702
R855 VDD1.n73 VDD1.n2 6.59444
R856 VDD1.n70 VDD1.n2 6.59444
R857 VDD1.n149 VDD1.n81 6.59444
R858 VDD1.n152 VDD1.n81 6.59444
R859 VDD1.n74 VDD1.n0 5.81868
R860 VDD1.n69 VDD1.n4 5.81868
R861 VDD1.n29 VDD1.n28 5.81868
R862 VDD1.n107 VDD1.n106 5.81868
R863 VDD1.n148 VDD1.n83 5.81868
R864 VDD1.n153 VDD1.n79 5.81868
R865 VDD1.n66 VDD1.n65 5.04292
R866 VDD1.n32 VDD1.n23 5.04292
R867 VDD1.n110 VDD1.n101 5.04292
R868 VDD1.n145 VDD1.n144 5.04292
R869 VDD1.n62 VDD1.n6 4.26717
R870 VDD1.n33 VDD1.n21 4.26717
R871 VDD1.n111 VDD1.n99 4.26717
R872 VDD1.n141 VDD1.n85 4.26717
R873 VDD1.n61 VDD1.n8 3.49141
R874 VDD1.n37 VDD1.n36 3.49141
R875 VDD1.n115 VDD1.n114 3.49141
R876 VDD1.n140 VDD1.n87 3.49141
R877 VDD1.n27 VDD1.n26 2.84303
R878 VDD1.n105 VDD1.n104 2.84303
R879 VDD1.n58 VDD1.n57 2.71565
R880 VDD1.n40 VDD1.n19 2.71565
R881 VDD1.n118 VDD1.n97 2.71565
R882 VDD1.n137 VDD1.n136 2.71565
R883 VDD1 VDD1.n161 2.45093
R884 VDD1.n54 VDD1.n10 1.93989
R885 VDD1.n41 VDD1.n17 1.93989
R886 VDD1.n119 VDD1.n95 1.93989
R887 VDD1.n133 VDD1.n89 1.93989
R888 VDD1.n160 VDD1.t4 1.39487
R889 VDD1.n160 VDD1.t9 1.39487
R890 VDD1.n77 VDD1.t5 1.39487
R891 VDD1.n77 VDD1.t3 1.39487
R892 VDD1.n158 VDD1.t6 1.39487
R893 VDD1.n158 VDD1.t7 1.39487
R894 VDD1.n156 VDD1.t2 1.39487
R895 VDD1.n156 VDD1.t0 1.39487
R896 VDD1.n53 VDD1.n12 1.16414
R897 VDD1.n45 VDD1.n44 1.16414
R898 VDD1.n124 VDD1.n122 1.16414
R899 VDD1.n132 VDD1.n91 1.16414
R900 VDD1 VDD1.n78 0.894897
R901 VDD1.n159 VDD1.n157 0.781361
R902 VDD1.n50 VDD1.n49 0.388379
R903 VDD1.n16 VDD1.n14 0.388379
R904 VDD1.n123 VDD1.n93 0.388379
R905 VDD1.n129 VDD1.n128 0.388379
R906 VDD1.n75 VDD1.n1 0.155672
R907 VDD1.n68 VDD1.n1 0.155672
R908 VDD1.n68 VDD1.n67 0.155672
R909 VDD1.n67 VDD1.n5 0.155672
R910 VDD1.n60 VDD1.n5 0.155672
R911 VDD1.n60 VDD1.n59 0.155672
R912 VDD1.n59 VDD1.n9 0.155672
R913 VDD1.n52 VDD1.n9 0.155672
R914 VDD1.n52 VDD1.n51 0.155672
R915 VDD1.n51 VDD1.n13 0.155672
R916 VDD1.n43 VDD1.n13 0.155672
R917 VDD1.n43 VDD1.n42 0.155672
R918 VDD1.n42 VDD1.n18 0.155672
R919 VDD1.n35 VDD1.n18 0.155672
R920 VDD1.n35 VDD1.n34 0.155672
R921 VDD1.n34 VDD1.n22 0.155672
R922 VDD1.n27 VDD1.n22 0.155672
R923 VDD1.n105 VDD1.n100 0.155672
R924 VDD1.n112 VDD1.n100 0.155672
R925 VDD1.n113 VDD1.n112 0.155672
R926 VDD1.n113 VDD1.n96 0.155672
R927 VDD1.n120 VDD1.n96 0.155672
R928 VDD1.n121 VDD1.n120 0.155672
R929 VDD1.n121 VDD1.n92 0.155672
R930 VDD1.n130 VDD1.n92 0.155672
R931 VDD1.n131 VDD1.n130 0.155672
R932 VDD1.n131 VDD1.n88 0.155672
R933 VDD1.n138 VDD1.n88 0.155672
R934 VDD1.n139 VDD1.n138 0.155672
R935 VDD1.n139 VDD1.n84 0.155672
R936 VDD1.n146 VDD1.n84 0.155672
R937 VDD1.n147 VDD1.n146 0.155672
R938 VDD1.n147 VDD1.n80 0.155672
R939 VDD1.n154 VDD1.n80 0.155672
R940 B.n1153 B.n1152 585
R941 B.n405 B.n192 585
R942 B.n404 B.n403 585
R943 B.n402 B.n401 585
R944 B.n400 B.n399 585
R945 B.n398 B.n397 585
R946 B.n396 B.n395 585
R947 B.n394 B.n393 585
R948 B.n392 B.n391 585
R949 B.n390 B.n389 585
R950 B.n388 B.n387 585
R951 B.n386 B.n385 585
R952 B.n384 B.n383 585
R953 B.n382 B.n381 585
R954 B.n380 B.n379 585
R955 B.n378 B.n377 585
R956 B.n376 B.n375 585
R957 B.n374 B.n373 585
R958 B.n372 B.n371 585
R959 B.n370 B.n369 585
R960 B.n368 B.n367 585
R961 B.n366 B.n365 585
R962 B.n364 B.n363 585
R963 B.n362 B.n361 585
R964 B.n360 B.n359 585
R965 B.n358 B.n357 585
R966 B.n356 B.n355 585
R967 B.n354 B.n353 585
R968 B.n352 B.n351 585
R969 B.n350 B.n349 585
R970 B.n348 B.n347 585
R971 B.n346 B.n345 585
R972 B.n344 B.n343 585
R973 B.n342 B.n341 585
R974 B.n340 B.n339 585
R975 B.n338 B.n337 585
R976 B.n336 B.n335 585
R977 B.n334 B.n333 585
R978 B.n332 B.n331 585
R979 B.n330 B.n329 585
R980 B.n328 B.n327 585
R981 B.n326 B.n325 585
R982 B.n324 B.n323 585
R983 B.n322 B.n321 585
R984 B.n320 B.n319 585
R985 B.n318 B.n317 585
R986 B.n316 B.n315 585
R987 B.n314 B.n313 585
R988 B.n312 B.n311 585
R989 B.n310 B.n309 585
R990 B.n308 B.n307 585
R991 B.n306 B.n305 585
R992 B.n304 B.n303 585
R993 B.n302 B.n301 585
R994 B.n300 B.n299 585
R995 B.n298 B.n297 585
R996 B.n296 B.n295 585
R997 B.n294 B.n293 585
R998 B.n292 B.n291 585
R999 B.n290 B.n289 585
R1000 B.n288 B.n287 585
R1001 B.n286 B.n285 585
R1002 B.n284 B.n283 585
R1003 B.n282 B.n281 585
R1004 B.n280 B.n279 585
R1005 B.n278 B.n277 585
R1006 B.n276 B.n275 585
R1007 B.n274 B.n273 585
R1008 B.n272 B.n271 585
R1009 B.n270 B.n269 585
R1010 B.n268 B.n267 585
R1011 B.n266 B.n265 585
R1012 B.n264 B.n263 585
R1013 B.n262 B.n261 585
R1014 B.n260 B.n259 585
R1015 B.n258 B.n257 585
R1016 B.n256 B.n255 585
R1017 B.n254 B.n253 585
R1018 B.n252 B.n251 585
R1019 B.n250 B.n249 585
R1020 B.n248 B.n247 585
R1021 B.n246 B.n245 585
R1022 B.n244 B.n243 585
R1023 B.n242 B.n241 585
R1024 B.n240 B.n239 585
R1025 B.n238 B.n237 585
R1026 B.n236 B.n235 585
R1027 B.n234 B.n233 585
R1028 B.n232 B.n231 585
R1029 B.n230 B.n229 585
R1030 B.n228 B.n227 585
R1031 B.n226 B.n225 585
R1032 B.n224 B.n223 585
R1033 B.n222 B.n221 585
R1034 B.n220 B.n219 585
R1035 B.n218 B.n217 585
R1036 B.n216 B.n215 585
R1037 B.n214 B.n213 585
R1038 B.n212 B.n211 585
R1039 B.n210 B.n209 585
R1040 B.n208 B.n207 585
R1041 B.n206 B.n205 585
R1042 B.n204 B.n203 585
R1043 B.n202 B.n201 585
R1044 B.n200 B.n199 585
R1045 B.n138 B.n137 585
R1046 B.n1151 B.n139 585
R1047 B.n1156 B.n139 585
R1048 B.n1150 B.n1149 585
R1049 B.n1149 B.n135 585
R1050 B.n1148 B.n134 585
R1051 B.n1162 B.n134 585
R1052 B.n1147 B.n133 585
R1053 B.n1163 B.n133 585
R1054 B.n1146 B.n132 585
R1055 B.n1164 B.n132 585
R1056 B.n1145 B.n1144 585
R1057 B.n1144 B.n128 585
R1058 B.n1143 B.n127 585
R1059 B.n1170 B.n127 585
R1060 B.n1142 B.n126 585
R1061 B.n1171 B.n126 585
R1062 B.n1141 B.n125 585
R1063 B.n1172 B.n125 585
R1064 B.n1140 B.n1139 585
R1065 B.n1139 B.n121 585
R1066 B.n1138 B.n120 585
R1067 B.n1178 B.n120 585
R1068 B.n1137 B.n119 585
R1069 B.n1179 B.n119 585
R1070 B.n1136 B.n118 585
R1071 B.n1180 B.n118 585
R1072 B.n1135 B.n1134 585
R1073 B.n1134 B.n114 585
R1074 B.n1133 B.n113 585
R1075 B.n1186 B.n113 585
R1076 B.n1132 B.n112 585
R1077 B.n1187 B.n112 585
R1078 B.n1131 B.n111 585
R1079 B.n1188 B.n111 585
R1080 B.n1130 B.n1129 585
R1081 B.n1129 B.n107 585
R1082 B.n1128 B.n106 585
R1083 B.n1194 B.n106 585
R1084 B.n1127 B.n105 585
R1085 B.n1195 B.n105 585
R1086 B.n1126 B.n104 585
R1087 B.n1196 B.n104 585
R1088 B.n1125 B.n1124 585
R1089 B.n1124 B.n100 585
R1090 B.n1123 B.n99 585
R1091 B.n1202 B.n99 585
R1092 B.n1122 B.n98 585
R1093 B.n1203 B.n98 585
R1094 B.n1121 B.n97 585
R1095 B.n1204 B.n97 585
R1096 B.n1120 B.n1119 585
R1097 B.n1119 B.n93 585
R1098 B.n1118 B.n92 585
R1099 B.n1210 B.n92 585
R1100 B.n1117 B.n91 585
R1101 B.n1211 B.n91 585
R1102 B.n1116 B.n90 585
R1103 B.n1212 B.n90 585
R1104 B.n1115 B.n1114 585
R1105 B.n1114 B.n86 585
R1106 B.n1113 B.n85 585
R1107 B.n1218 B.n85 585
R1108 B.n1112 B.n84 585
R1109 B.n1219 B.n84 585
R1110 B.n1111 B.n83 585
R1111 B.n1220 B.n83 585
R1112 B.n1110 B.n1109 585
R1113 B.n1109 B.n79 585
R1114 B.n1108 B.n78 585
R1115 B.n1226 B.n78 585
R1116 B.n1107 B.n77 585
R1117 B.n1227 B.n77 585
R1118 B.n1106 B.n76 585
R1119 B.n1228 B.n76 585
R1120 B.n1105 B.n1104 585
R1121 B.n1104 B.n72 585
R1122 B.n1103 B.n71 585
R1123 B.n1234 B.n71 585
R1124 B.n1102 B.n70 585
R1125 B.n1235 B.n70 585
R1126 B.n1101 B.n69 585
R1127 B.n1236 B.n69 585
R1128 B.n1100 B.n1099 585
R1129 B.n1099 B.n65 585
R1130 B.n1098 B.n64 585
R1131 B.n1242 B.n64 585
R1132 B.n1097 B.n63 585
R1133 B.n1243 B.n63 585
R1134 B.n1096 B.n62 585
R1135 B.n1244 B.n62 585
R1136 B.n1095 B.n1094 585
R1137 B.n1094 B.n58 585
R1138 B.n1093 B.n57 585
R1139 B.n1250 B.n57 585
R1140 B.n1092 B.n56 585
R1141 B.n1251 B.n56 585
R1142 B.n1091 B.n55 585
R1143 B.n1252 B.n55 585
R1144 B.n1090 B.n1089 585
R1145 B.n1089 B.n51 585
R1146 B.n1088 B.n50 585
R1147 B.n1258 B.n50 585
R1148 B.n1087 B.n49 585
R1149 B.n1259 B.n49 585
R1150 B.n1086 B.n48 585
R1151 B.n1260 B.n48 585
R1152 B.n1085 B.n1084 585
R1153 B.n1084 B.n44 585
R1154 B.n1083 B.n43 585
R1155 B.n1266 B.n43 585
R1156 B.n1082 B.n42 585
R1157 B.n1267 B.n42 585
R1158 B.n1081 B.n41 585
R1159 B.n1268 B.n41 585
R1160 B.n1080 B.n1079 585
R1161 B.n1079 B.n40 585
R1162 B.n1078 B.n36 585
R1163 B.n1274 B.n36 585
R1164 B.n1077 B.n35 585
R1165 B.n1275 B.n35 585
R1166 B.n1076 B.n34 585
R1167 B.n1276 B.n34 585
R1168 B.n1075 B.n1074 585
R1169 B.n1074 B.n30 585
R1170 B.n1073 B.n29 585
R1171 B.n1282 B.n29 585
R1172 B.n1072 B.n28 585
R1173 B.n1283 B.n28 585
R1174 B.n1071 B.n27 585
R1175 B.n1284 B.n27 585
R1176 B.n1070 B.n1069 585
R1177 B.n1069 B.n23 585
R1178 B.n1068 B.n22 585
R1179 B.n1290 B.n22 585
R1180 B.n1067 B.n21 585
R1181 B.n1291 B.n21 585
R1182 B.n1066 B.n20 585
R1183 B.n1292 B.n20 585
R1184 B.n1065 B.n1064 585
R1185 B.n1064 B.n19 585
R1186 B.n1063 B.n15 585
R1187 B.n1298 B.n15 585
R1188 B.n1062 B.n14 585
R1189 B.n1299 B.n14 585
R1190 B.n1061 B.n13 585
R1191 B.n1300 B.n13 585
R1192 B.n1060 B.n1059 585
R1193 B.n1059 B.n12 585
R1194 B.n1058 B.n1057 585
R1195 B.n1058 B.n8 585
R1196 B.n1056 B.n7 585
R1197 B.n1307 B.n7 585
R1198 B.n1055 B.n6 585
R1199 B.n1308 B.n6 585
R1200 B.n1054 B.n5 585
R1201 B.n1309 B.n5 585
R1202 B.n1053 B.n1052 585
R1203 B.n1052 B.n4 585
R1204 B.n1051 B.n406 585
R1205 B.n1051 B.n1050 585
R1206 B.n1041 B.n407 585
R1207 B.n408 B.n407 585
R1208 B.n1043 B.n1042 585
R1209 B.n1044 B.n1043 585
R1210 B.n1040 B.n413 585
R1211 B.n413 B.n412 585
R1212 B.n1039 B.n1038 585
R1213 B.n1038 B.n1037 585
R1214 B.n415 B.n414 585
R1215 B.n1030 B.n415 585
R1216 B.n1029 B.n1028 585
R1217 B.n1031 B.n1029 585
R1218 B.n1027 B.n420 585
R1219 B.n420 B.n419 585
R1220 B.n1026 B.n1025 585
R1221 B.n1025 B.n1024 585
R1222 B.n422 B.n421 585
R1223 B.n423 B.n422 585
R1224 B.n1017 B.n1016 585
R1225 B.n1018 B.n1017 585
R1226 B.n1015 B.n428 585
R1227 B.n428 B.n427 585
R1228 B.n1014 B.n1013 585
R1229 B.n1013 B.n1012 585
R1230 B.n430 B.n429 585
R1231 B.n431 B.n430 585
R1232 B.n1005 B.n1004 585
R1233 B.n1006 B.n1005 585
R1234 B.n1003 B.n436 585
R1235 B.n436 B.n435 585
R1236 B.n1002 B.n1001 585
R1237 B.n1001 B.n1000 585
R1238 B.n438 B.n437 585
R1239 B.n993 B.n438 585
R1240 B.n992 B.n991 585
R1241 B.n994 B.n992 585
R1242 B.n990 B.n443 585
R1243 B.n443 B.n442 585
R1244 B.n989 B.n988 585
R1245 B.n988 B.n987 585
R1246 B.n445 B.n444 585
R1247 B.n446 B.n445 585
R1248 B.n980 B.n979 585
R1249 B.n981 B.n980 585
R1250 B.n978 B.n451 585
R1251 B.n451 B.n450 585
R1252 B.n977 B.n976 585
R1253 B.n976 B.n975 585
R1254 B.n453 B.n452 585
R1255 B.n454 B.n453 585
R1256 B.n968 B.n967 585
R1257 B.n969 B.n968 585
R1258 B.n966 B.n459 585
R1259 B.n459 B.n458 585
R1260 B.n965 B.n964 585
R1261 B.n964 B.n963 585
R1262 B.n461 B.n460 585
R1263 B.n462 B.n461 585
R1264 B.n956 B.n955 585
R1265 B.n957 B.n956 585
R1266 B.n954 B.n467 585
R1267 B.n467 B.n466 585
R1268 B.n953 B.n952 585
R1269 B.n952 B.n951 585
R1270 B.n469 B.n468 585
R1271 B.n470 B.n469 585
R1272 B.n944 B.n943 585
R1273 B.n945 B.n944 585
R1274 B.n942 B.n475 585
R1275 B.n475 B.n474 585
R1276 B.n941 B.n940 585
R1277 B.n940 B.n939 585
R1278 B.n477 B.n476 585
R1279 B.n478 B.n477 585
R1280 B.n932 B.n931 585
R1281 B.n933 B.n932 585
R1282 B.n930 B.n483 585
R1283 B.n483 B.n482 585
R1284 B.n929 B.n928 585
R1285 B.n928 B.n927 585
R1286 B.n485 B.n484 585
R1287 B.n486 B.n485 585
R1288 B.n920 B.n919 585
R1289 B.n921 B.n920 585
R1290 B.n918 B.n491 585
R1291 B.n491 B.n490 585
R1292 B.n917 B.n916 585
R1293 B.n916 B.n915 585
R1294 B.n493 B.n492 585
R1295 B.n494 B.n493 585
R1296 B.n908 B.n907 585
R1297 B.n909 B.n908 585
R1298 B.n906 B.n499 585
R1299 B.n499 B.n498 585
R1300 B.n905 B.n904 585
R1301 B.n904 B.n903 585
R1302 B.n501 B.n500 585
R1303 B.n502 B.n501 585
R1304 B.n896 B.n895 585
R1305 B.n897 B.n896 585
R1306 B.n894 B.n506 585
R1307 B.n510 B.n506 585
R1308 B.n893 B.n892 585
R1309 B.n892 B.n891 585
R1310 B.n508 B.n507 585
R1311 B.n509 B.n508 585
R1312 B.n884 B.n883 585
R1313 B.n885 B.n884 585
R1314 B.n882 B.n515 585
R1315 B.n515 B.n514 585
R1316 B.n881 B.n880 585
R1317 B.n880 B.n879 585
R1318 B.n517 B.n516 585
R1319 B.n518 B.n517 585
R1320 B.n872 B.n871 585
R1321 B.n873 B.n872 585
R1322 B.n870 B.n523 585
R1323 B.n523 B.n522 585
R1324 B.n869 B.n868 585
R1325 B.n868 B.n867 585
R1326 B.n525 B.n524 585
R1327 B.n526 B.n525 585
R1328 B.n860 B.n859 585
R1329 B.n861 B.n860 585
R1330 B.n858 B.n531 585
R1331 B.n531 B.n530 585
R1332 B.n857 B.n856 585
R1333 B.n856 B.n855 585
R1334 B.n533 B.n532 585
R1335 B.n534 B.n533 585
R1336 B.n848 B.n847 585
R1337 B.n849 B.n848 585
R1338 B.n846 B.n539 585
R1339 B.n539 B.n538 585
R1340 B.n845 B.n844 585
R1341 B.n844 B.n843 585
R1342 B.n541 B.n540 585
R1343 B.n542 B.n541 585
R1344 B.n836 B.n835 585
R1345 B.n837 B.n836 585
R1346 B.n834 B.n547 585
R1347 B.n547 B.n546 585
R1348 B.n833 B.n832 585
R1349 B.n832 B.n831 585
R1350 B.n549 B.n548 585
R1351 B.n550 B.n549 585
R1352 B.n824 B.n823 585
R1353 B.n825 B.n824 585
R1354 B.n553 B.n552 585
R1355 B.n612 B.n610 585
R1356 B.n613 B.n609 585
R1357 B.n613 B.n554 585
R1358 B.n616 B.n615 585
R1359 B.n617 B.n608 585
R1360 B.n619 B.n618 585
R1361 B.n621 B.n607 585
R1362 B.n624 B.n623 585
R1363 B.n625 B.n606 585
R1364 B.n627 B.n626 585
R1365 B.n629 B.n605 585
R1366 B.n632 B.n631 585
R1367 B.n633 B.n604 585
R1368 B.n635 B.n634 585
R1369 B.n637 B.n603 585
R1370 B.n640 B.n639 585
R1371 B.n641 B.n602 585
R1372 B.n643 B.n642 585
R1373 B.n645 B.n601 585
R1374 B.n648 B.n647 585
R1375 B.n649 B.n600 585
R1376 B.n651 B.n650 585
R1377 B.n653 B.n599 585
R1378 B.n656 B.n655 585
R1379 B.n657 B.n598 585
R1380 B.n659 B.n658 585
R1381 B.n661 B.n597 585
R1382 B.n664 B.n663 585
R1383 B.n665 B.n596 585
R1384 B.n667 B.n666 585
R1385 B.n669 B.n595 585
R1386 B.n672 B.n671 585
R1387 B.n673 B.n594 585
R1388 B.n675 B.n674 585
R1389 B.n677 B.n593 585
R1390 B.n680 B.n679 585
R1391 B.n681 B.n592 585
R1392 B.n683 B.n682 585
R1393 B.n685 B.n591 585
R1394 B.n688 B.n687 585
R1395 B.n689 B.n590 585
R1396 B.n691 B.n690 585
R1397 B.n693 B.n589 585
R1398 B.n696 B.n695 585
R1399 B.n697 B.n588 585
R1400 B.n699 B.n698 585
R1401 B.n701 B.n587 585
R1402 B.n704 B.n703 585
R1403 B.n706 B.n584 585
R1404 B.n708 B.n707 585
R1405 B.n710 B.n583 585
R1406 B.n713 B.n712 585
R1407 B.n714 B.n582 585
R1408 B.n716 B.n715 585
R1409 B.n718 B.n581 585
R1410 B.n721 B.n720 585
R1411 B.n722 B.n580 585
R1412 B.n727 B.n726 585
R1413 B.n729 B.n579 585
R1414 B.n732 B.n731 585
R1415 B.n733 B.n578 585
R1416 B.n735 B.n734 585
R1417 B.n737 B.n577 585
R1418 B.n740 B.n739 585
R1419 B.n741 B.n576 585
R1420 B.n743 B.n742 585
R1421 B.n745 B.n575 585
R1422 B.n748 B.n747 585
R1423 B.n749 B.n574 585
R1424 B.n751 B.n750 585
R1425 B.n753 B.n573 585
R1426 B.n756 B.n755 585
R1427 B.n757 B.n572 585
R1428 B.n759 B.n758 585
R1429 B.n761 B.n571 585
R1430 B.n764 B.n763 585
R1431 B.n765 B.n570 585
R1432 B.n767 B.n766 585
R1433 B.n769 B.n569 585
R1434 B.n772 B.n771 585
R1435 B.n773 B.n568 585
R1436 B.n775 B.n774 585
R1437 B.n777 B.n567 585
R1438 B.n780 B.n779 585
R1439 B.n781 B.n566 585
R1440 B.n783 B.n782 585
R1441 B.n785 B.n565 585
R1442 B.n788 B.n787 585
R1443 B.n789 B.n564 585
R1444 B.n791 B.n790 585
R1445 B.n793 B.n563 585
R1446 B.n796 B.n795 585
R1447 B.n797 B.n562 585
R1448 B.n799 B.n798 585
R1449 B.n801 B.n561 585
R1450 B.n804 B.n803 585
R1451 B.n805 B.n560 585
R1452 B.n807 B.n806 585
R1453 B.n809 B.n559 585
R1454 B.n812 B.n811 585
R1455 B.n813 B.n558 585
R1456 B.n815 B.n814 585
R1457 B.n817 B.n557 585
R1458 B.n818 B.n556 585
R1459 B.n821 B.n820 585
R1460 B.n822 B.n555 585
R1461 B.n555 B.n554 585
R1462 B.n827 B.n826 585
R1463 B.n826 B.n825 585
R1464 B.n828 B.n551 585
R1465 B.n551 B.n550 585
R1466 B.n830 B.n829 585
R1467 B.n831 B.n830 585
R1468 B.n545 B.n544 585
R1469 B.n546 B.n545 585
R1470 B.n839 B.n838 585
R1471 B.n838 B.n837 585
R1472 B.n840 B.n543 585
R1473 B.n543 B.n542 585
R1474 B.n842 B.n841 585
R1475 B.n843 B.n842 585
R1476 B.n537 B.n536 585
R1477 B.n538 B.n537 585
R1478 B.n851 B.n850 585
R1479 B.n850 B.n849 585
R1480 B.n852 B.n535 585
R1481 B.n535 B.n534 585
R1482 B.n854 B.n853 585
R1483 B.n855 B.n854 585
R1484 B.n529 B.n528 585
R1485 B.n530 B.n529 585
R1486 B.n863 B.n862 585
R1487 B.n862 B.n861 585
R1488 B.n864 B.n527 585
R1489 B.n527 B.n526 585
R1490 B.n866 B.n865 585
R1491 B.n867 B.n866 585
R1492 B.n521 B.n520 585
R1493 B.n522 B.n521 585
R1494 B.n875 B.n874 585
R1495 B.n874 B.n873 585
R1496 B.n876 B.n519 585
R1497 B.n519 B.n518 585
R1498 B.n878 B.n877 585
R1499 B.n879 B.n878 585
R1500 B.n513 B.n512 585
R1501 B.n514 B.n513 585
R1502 B.n887 B.n886 585
R1503 B.n886 B.n885 585
R1504 B.n888 B.n511 585
R1505 B.n511 B.n509 585
R1506 B.n890 B.n889 585
R1507 B.n891 B.n890 585
R1508 B.n505 B.n504 585
R1509 B.n510 B.n505 585
R1510 B.n899 B.n898 585
R1511 B.n898 B.n897 585
R1512 B.n900 B.n503 585
R1513 B.n503 B.n502 585
R1514 B.n902 B.n901 585
R1515 B.n903 B.n902 585
R1516 B.n497 B.n496 585
R1517 B.n498 B.n497 585
R1518 B.n911 B.n910 585
R1519 B.n910 B.n909 585
R1520 B.n912 B.n495 585
R1521 B.n495 B.n494 585
R1522 B.n914 B.n913 585
R1523 B.n915 B.n914 585
R1524 B.n489 B.n488 585
R1525 B.n490 B.n489 585
R1526 B.n923 B.n922 585
R1527 B.n922 B.n921 585
R1528 B.n924 B.n487 585
R1529 B.n487 B.n486 585
R1530 B.n926 B.n925 585
R1531 B.n927 B.n926 585
R1532 B.n481 B.n480 585
R1533 B.n482 B.n481 585
R1534 B.n935 B.n934 585
R1535 B.n934 B.n933 585
R1536 B.n936 B.n479 585
R1537 B.n479 B.n478 585
R1538 B.n938 B.n937 585
R1539 B.n939 B.n938 585
R1540 B.n473 B.n472 585
R1541 B.n474 B.n473 585
R1542 B.n947 B.n946 585
R1543 B.n946 B.n945 585
R1544 B.n948 B.n471 585
R1545 B.n471 B.n470 585
R1546 B.n950 B.n949 585
R1547 B.n951 B.n950 585
R1548 B.n465 B.n464 585
R1549 B.n466 B.n465 585
R1550 B.n959 B.n958 585
R1551 B.n958 B.n957 585
R1552 B.n960 B.n463 585
R1553 B.n463 B.n462 585
R1554 B.n962 B.n961 585
R1555 B.n963 B.n962 585
R1556 B.n457 B.n456 585
R1557 B.n458 B.n457 585
R1558 B.n971 B.n970 585
R1559 B.n970 B.n969 585
R1560 B.n972 B.n455 585
R1561 B.n455 B.n454 585
R1562 B.n974 B.n973 585
R1563 B.n975 B.n974 585
R1564 B.n449 B.n448 585
R1565 B.n450 B.n449 585
R1566 B.n983 B.n982 585
R1567 B.n982 B.n981 585
R1568 B.n984 B.n447 585
R1569 B.n447 B.n446 585
R1570 B.n986 B.n985 585
R1571 B.n987 B.n986 585
R1572 B.n441 B.n440 585
R1573 B.n442 B.n441 585
R1574 B.n996 B.n995 585
R1575 B.n995 B.n994 585
R1576 B.n997 B.n439 585
R1577 B.n993 B.n439 585
R1578 B.n999 B.n998 585
R1579 B.n1000 B.n999 585
R1580 B.n434 B.n433 585
R1581 B.n435 B.n434 585
R1582 B.n1008 B.n1007 585
R1583 B.n1007 B.n1006 585
R1584 B.n1009 B.n432 585
R1585 B.n432 B.n431 585
R1586 B.n1011 B.n1010 585
R1587 B.n1012 B.n1011 585
R1588 B.n426 B.n425 585
R1589 B.n427 B.n426 585
R1590 B.n1020 B.n1019 585
R1591 B.n1019 B.n1018 585
R1592 B.n1021 B.n424 585
R1593 B.n424 B.n423 585
R1594 B.n1023 B.n1022 585
R1595 B.n1024 B.n1023 585
R1596 B.n418 B.n417 585
R1597 B.n419 B.n418 585
R1598 B.n1033 B.n1032 585
R1599 B.n1032 B.n1031 585
R1600 B.n1034 B.n416 585
R1601 B.n1030 B.n416 585
R1602 B.n1036 B.n1035 585
R1603 B.n1037 B.n1036 585
R1604 B.n411 B.n410 585
R1605 B.n412 B.n411 585
R1606 B.n1046 B.n1045 585
R1607 B.n1045 B.n1044 585
R1608 B.n1047 B.n409 585
R1609 B.n409 B.n408 585
R1610 B.n1049 B.n1048 585
R1611 B.n1050 B.n1049 585
R1612 B.n3 B.n0 585
R1613 B.n4 B.n3 585
R1614 B.n1306 B.n1 585
R1615 B.n1307 B.n1306 585
R1616 B.n1305 B.n1304 585
R1617 B.n1305 B.n8 585
R1618 B.n1303 B.n9 585
R1619 B.n12 B.n9 585
R1620 B.n1302 B.n1301 585
R1621 B.n1301 B.n1300 585
R1622 B.n11 B.n10 585
R1623 B.n1299 B.n11 585
R1624 B.n1297 B.n1296 585
R1625 B.n1298 B.n1297 585
R1626 B.n1295 B.n16 585
R1627 B.n19 B.n16 585
R1628 B.n1294 B.n1293 585
R1629 B.n1293 B.n1292 585
R1630 B.n18 B.n17 585
R1631 B.n1291 B.n18 585
R1632 B.n1289 B.n1288 585
R1633 B.n1290 B.n1289 585
R1634 B.n1287 B.n24 585
R1635 B.n24 B.n23 585
R1636 B.n1286 B.n1285 585
R1637 B.n1285 B.n1284 585
R1638 B.n26 B.n25 585
R1639 B.n1283 B.n26 585
R1640 B.n1281 B.n1280 585
R1641 B.n1282 B.n1281 585
R1642 B.n1279 B.n31 585
R1643 B.n31 B.n30 585
R1644 B.n1278 B.n1277 585
R1645 B.n1277 B.n1276 585
R1646 B.n33 B.n32 585
R1647 B.n1275 B.n33 585
R1648 B.n1273 B.n1272 585
R1649 B.n1274 B.n1273 585
R1650 B.n1271 B.n37 585
R1651 B.n40 B.n37 585
R1652 B.n1270 B.n1269 585
R1653 B.n1269 B.n1268 585
R1654 B.n39 B.n38 585
R1655 B.n1267 B.n39 585
R1656 B.n1265 B.n1264 585
R1657 B.n1266 B.n1265 585
R1658 B.n1263 B.n45 585
R1659 B.n45 B.n44 585
R1660 B.n1262 B.n1261 585
R1661 B.n1261 B.n1260 585
R1662 B.n47 B.n46 585
R1663 B.n1259 B.n47 585
R1664 B.n1257 B.n1256 585
R1665 B.n1258 B.n1257 585
R1666 B.n1255 B.n52 585
R1667 B.n52 B.n51 585
R1668 B.n1254 B.n1253 585
R1669 B.n1253 B.n1252 585
R1670 B.n54 B.n53 585
R1671 B.n1251 B.n54 585
R1672 B.n1249 B.n1248 585
R1673 B.n1250 B.n1249 585
R1674 B.n1247 B.n59 585
R1675 B.n59 B.n58 585
R1676 B.n1246 B.n1245 585
R1677 B.n1245 B.n1244 585
R1678 B.n61 B.n60 585
R1679 B.n1243 B.n61 585
R1680 B.n1241 B.n1240 585
R1681 B.n1242 B.n1241 585
R1682 B.n1239 B.n66 585
R1683 B.n66 B.n65 585
R1684 B.n1238 B.n1237 585
R1685 B.n1237 B.n1236 585
R1686 B.n68 B.n67 585
R1687 B.n1235 B.n68 585
R1688 B.n1233 B.n1232 585
R1689 B.n1234 B.n1233 585
R1690 B.n1231 B.n73 585
R1691 B.n73 B.n72 585
R1692 B.n1230 B.n1229 585
R1693 B.n1229 B.n1228 585
R1694 B.n75 B.n74 585
R1695 B.n1227 B.n75 585
R1696 B.n1225 B.n1224 585
R1697 B.n1226 B.n1225 585
R1698 B.n1223 B.n80 585
R1699 B.n80 B.n79 585
R1700 B.n1222 B.n1221 585
R1701 B.n1221 B.n1220 585
R1702 B.n82 B.n81 585
R1703 B.n1219 B.n82 585
R1704 B.n1217 B.n1216 585
R1705 B.n1218 B.n1217 585
R1706 B.n1215 B.n87 585
R1707 B.n87 B.n86 585
R1708 B.n1214 B.n1213 585
R1709 B.n1213 B.n1212 585
R1710 B.n89 B.n88 585
R1711 B.n1211 B.n89 585
R1712 B.n1209 B.n1208 585
R1713 B.n1210 B.n1209 585
R1714 B.n1207 B.n94 585
R1715 B.n94 B.n93 585
R1716 B.n1206 B.n1205 585
R1717 B.n1205 B.n1204 585
R1718 B.n96 B.n95 585
R1719 B.n1203 B.n96 585
R1720 B.n1201 B.n1200 585
R1721 B.n1202 B.n1201 585
R1722 B.n1199 B.n101 585
R1723 B.n101 B.n100 585
R1724 B.n1198 B.n1197 585
R1725 B.n1197 B.n1196 585
R1726 B.n103 B.n102 585
R1727 B.n1195 B.n103 585
R1728 B.n1193 B.n1192 585
R1729 B.n1194 B.n1193 585
R1730 B.n1191 B.n108 585
R1731 B.n108 B.n107 585
R1732 B.n1190 B.n1189 585
R1733 B.n1189 B.n1188 585
R1734 B.n110 B.n109 585
R1735 B.n1187 B.n110 585
R1736 B.n1185 B.n1184 585
R1737 B.n1186 B.n1185 585
R1738 B.n1183 B.n115 585
R1739 B.n115 B.n114 585
R1740 B.n1182 B.n1181 585
R1741 B.n1181 B.n1180 585
R1742 B.n117 B.n116 585
R1743 B.n1179 B.n117 585
R1744 B.n1177 B.n1176 585
R1745 B.n1178 B.n1177 585
R1746 B.n1175 B.n122 585
R1747 B.n122 B.n121 585
R1748 B.n1174 B.n1173 585
R1749 B.n1173 B.n1172 585
R1750 B.n124 B.n123 585
R1751 B.n1171 B.n124 585
R1752 B.n1169 B.n1168 585
R1753 B.n1170 B.n1169 585
R1754 B.n1167 B.n129 585
R1755 B.n129 B.n128 585
R1756 B.n1166 B.n1165 585
R1757 B.n1165 B.n1164 585
R1758 B.n131 B.n130 585
R1759 B.n1163 B.n131 585
R1760 B.n1161 B.n1160 585
R1761 B.n1162 B.n1161 585
R1762 B.n1159 B.n136 585
R1763 B.n136 B.n135 585
R1764 B.n1158 B.n1157 585
R1765 B.n1157 B.n1156 585
R1766 B.n1310 B.n1309 585
R1767 B.n1308 B.n2 585
R1768 B.n1157 B.n138 492.5
R1769 B.n1153 B.n139 492.5
R1770 B.n824 B.n555 492.5
R1771 B.n826 B.n553 492.5
R1772 B.n193 B.t19 395.497
R1773 B.n723 B.t17 395.497
R1774 B.n196 B.t12 395.497
R1775 B.n585 B.t23 395.497
R1776 B.n194 B.t20 320.248
R1777 B.n724 B.t16 320.248
R1778 B.n197 B.t13 320.248
R1779 B.n586 B.t22 320.248
R1780 B.n196 B.t10 305.538
R1781 B.n193 B.t18 305.538
R1782 B.n723 B.t14 305.538
R1783 B.n585 B.t21 305.538
R1784 B.n1155 B.n1154 256.663
R1785 B.n1155 B.n191 256.663
R1786 B.n1155 B.n190 256.663
R1787 B.n1155 B.n189 256.663
R1788 B.n1155 B.n188 256.663
R1789 B.n1155 B.n187 256.663
R1790 B.n1155 B.n186 256.663
R1791 B.n1155 B.n185 256.663
R1792 B.n1155 B.n184 256.663
R1793 B.n1155 B.n183 256.663
R1794 B.n1155 B.n182 256.663
R1795 B.n1155 B.n181 256.663
R1796 B.n1155 B.n180 256.663
R1797 B.n1155 B.n179 256.663
R1798 B.n1155 B.n178 256.663
R1799 B.n1155 B.n177 256.663
R1800 B.n1155 B.n176 256.663
R1801 B.n1155 B.n175 256.663
R1802 B.n1155 B.n174 256.663
R1803 B.n1155 B.n173 256.663
R1804 B.n1155 B.n172 256.663
R1805 B.n1155 B.n171 256.663
R1806 B.n1155 B.n170 256.663
R1807 B.n1155 B.n169 256.663
R1808 B.n1155 B.n168 256.663
R1809 B.n1155 B.n167 256.663
R1810 B.n1155 B.n166 256.663
R1811 B.n1155 B.n165 256.663
R1812 B.n1155 B.n164 256.663
R1813 B.n1155 B.n163 256.663
R1814 B.n1155 B.n162 256.663
R1815 B.n1155 B.n161 256.663
R1816 B.n1155 B.n160 256.663
R1817 B.n1155 B.n159 256.663
R1818 B.n1155 B.n158 256.663
R1819 B.n1155 B.n157 256.663
R1820 B.n1155 B.n156 256.663
R1821 B.n1155 B.n155 256.663
R1822 B.n1155 B.n154 256.663
R1823 B.n1155 B.n153 256.663
R1824 B.n1155 B.n152 256.663
R1825 B.n1155 B.n151 256.663
R1826 B.n1155 B.n150 256.663
R1827 B.n1155 B.n149 256.663
R1828 B.n1155 B.n148 256.663
R1829 B.n1155 B.n147 256.663
R1830 B.n1155 B.n146 256.663
R1831 B.n1155 B.n145 256.663
R1832 B.n1155 B.n144 256.663
R1833 B.n1155 B.n143 256.663
R1834 B.n1155 B.n142 256.663
R1835 B.n1155 B.n141 256.663
R1836 B.n1155 B.n140 256.663
R1837 B.n611 B.n554 256.663
R1838 B.n614 B.n554 256.663
R1839 B.n620 B.n554 256.663
R1840 B.n622 B.n554 256.663
R1841 B.n628 B.n554 256.663
R1842 B.n630 B.n554 256.663
R1843 B.n636 B.n554 256.663
R1844 B.n638 B.n554 256.663
R1845 B.n644 B.n554 256.663
R1846 B.n646 B.n554 256.663
R1847 B.n652 B.n554 256.663
R1848 B.n654 B.n554 256.663
R1849 B.n660 B.n554 256.663
R1850 B.n662 B.n554 256.663
R1851 B.n668 B.n554 256.663
R1852 B.n670 B.n554 256.663
R1853 B.n676 B.n554 256.663
R1854 B.n678 B.n554 256.663
R1855 B.n684 B.n554 256.663
R1856 B.n686 B.n554 256.663
R1857 B.n692 B.n554 256.663
R1858 B.n694 B.n554 256.663
R1859 B.n700 B.n554 256.663
R1860 B.n702 B.n554 256.663
R1861 B.n709 B.n554 256.663
R1862 B.n711 B.n554 256.663
R1863 B.n717 B.n554 256.663
R1864 B.n719 B.n554 256.663
R1865 B.n728 B.n554 256.663
R1866 B.n730 B.n554 256.663
R1867 B.n736 B.n554 256.663
R1868 B.n738 B.n554 256.663
R1869 B.n744 B.n554 256.663
R1870 B.n746 B.n554 256.663
R1871 B.n752 B.n554 256.663
R1872 B.n754 B.n554 256.663
R1873 B.n760 B.n554 256.663
R1874 B.n762 B.n554 256.663
R1875 B.n768 B.n554 256.663
R1876 B.n770 B.n554 256.663
R1877 B.n776 B.n554 256.663
R1878 B.n778 B.n554 256.663
R1879 B.n784 B.n554 256.663
R1880 B.n786 B.n554 256.663
R1881 B.n792 B.n554 256.663
R1882 B.n794 B.n554 256.663
R1883 B.n800 B.n554 256.663
R1884 B.n802 B.n554 256.663
R1885 B.n808 B.n554 256.663
R1886 B.n810 B.n554 256.663
R1887 B.n816 B.n554 256.663
R1888 B.n819 B.n554 256.663
R1889 B.n1312 B.n1311 256.663
R1890 B.n201 B.n200 163.367
R1891 B.n205 B.n204 163.367
R1892 B.n209 B.n208 163.367
R1893 B.n213 B.n212 163.367
R1894 B.n217 B.n216 163.367
R1895 B.n221 B.n220 163.367
R1896 B.n225 B.n224 163.367
R1897 B.n229 B.n228 163.367
R1898 B.n233 B.n232 163.367
R1899 B.n237 B.n236 163.367
R1900 B.n241 B.n240 163.367
R1901 B.n245 B.n244 163.367
R1902 B.n249 B.n248 163.367
R1903 B.n253 B.n252 163.367
R1904 B.n257 B.n256 163.367
R1905 B.n261 B.n260 163.367
R1906 B.n265 B.n264 163.367
R1907 B.n269 B.n268 163.367
R1908 B.n273 B.n272 163.367
R1909 B.n277 B.n276 163.367
R1910 B.n281 B.n280 163.367
R1911 B.n285 B.n284 163.367
R1912 B.n289 B.n288 163.367
R1913 B.n293 B.n292 163.367
R1914 B.n297 B.n296 163.367
R1915 B.n301 B.n300 163.367
R1916 B.n305 B.n304 163.367
R1917 B.n309 B.n308 163.367
R1918 B.n313 B.n312 163.367
R1919 B.n317 B.n316 163.367
R1920 B.n321 B.n320 163.367
R1921 B.n325 B.n324 163.367
R1922 B.n329 B.n328 163.367
R1923 B.n333 B.n332 163.367
R1924 B.n337 B.n336 163.367
R1925 B.n341 B.n340 163.367
R1926 B.n345 B.n344 163.367
R1927 B.n349 B.n348 163.367
R1928 B.n353 B.n352 163.367
R1929 B.n357 B.n356 163.367
R1930 B.n361 B.n360 163.367
R1931 B.n365 B.n364 163.367
R1932 B.n369 B.n368 163.367
R1933 B.n373 B.n372 163.367
R1934 B.n377 B.n376 163.367
R1935 B.n381 B.n380 163.367
R1936 B.n385 B.n384 163.367
R1937 B.n389 B.n388 163.367
R1938 B.n393 B.n392 163.367
R1939 B.n397 B.n396 163.367
R1940 B.n401 B.n400 163.367
R1941 B.n403 B.n192 163.367
R1942 B.n824 B.n549 163.367
R1943 B.n832 B.n549 163.367
R1944 B.n832 B.n547 163.367
R1945 B.n836 B.n547 163.367
R1946 B.n836 B.n541 163.367
R1947 B.n844 B.n541 163.367
R1948 B.n844 B.n539 163.367
R1949 B.n848 B.n539 163.367
R1950 B.n848 B.n533 163.367
R1951 B.n856 B.n533 163.367
R1952 B.n856 B.n531 163.367
R1953 B.n860 B.n531 163.367
R1954 B.n860 B.n525 163.367
R1955 B.n868 B.n525 163.367
R1956 B.n868 B.n523 163.367
R1957 B.n872 B.n523 163.367
R1958 B.n872 B.n517 163.367
R1959 B.n880 B.n517 163.367
R1960 B.n880 B.n515 163.367
R1961 B.n884 B.n515 163.367
R1962 B.n884 B.n508 163.367
R1963 B.n892 B.n508 163.367
R1964 B.n892 B.n506 163.367
R1965 B.n896 B.n506 163.367
R1966 B.n896 B.n501 163.367
R1967 B.n904 B.n501 163.367
R1968 B.n904 B.n499 163.367
R1969 B.n908 B.n499 163.367
R1970 B.n908 B.n493 163.367
R1971 B.n916 B.n493 163.367
R1972 B.n916 B.n491 163.367
R1973 B.n920 B.n491 163.367
R1974 B.n920 B.n485 163.367
R1975 B.n928 B.n485 163.367
R1976 B.n928 B.n483 163.367
R1977 B.n932 B.n483 163.367
R1978 B.n932 B.n477 163.367
R1979 B.n940 B.n477 163.367
R1980 B.n940 B.n475 163.367
R1981 B.n944 B.n475 163.367
R1982 B.n944 B.n469 163.367
R1983 B.n952 B.n469 163.367
R1984 B.n952 B.n467 163.367
R1985 B.n956 B.n467 163.367
R1986 B.n956 B.n461 163.367
R1987 B.n964 B.n461 163.367
R1988 B.n964 B.n459 163.367
R1989 B.n968 B.n459 163.367
R1990 B.n968 B.n453 163.367
R1991 B.n976 B.n453 163.367
R1992 B.n976 B.n451 163.367
R1993 B.n980 B.n451 163.367
R1994 B.n980 B.n445 163.367
R1995 B.n988 B.n445 163.367
R1996 B.n988 B.n443 163.367
R1997 B.n992 B.n443 163.367
R1998 B.n992 B.n438 163.367
R1999 B.n1001 B.n438 163.367
R2000 B.n1001 B.n436 163.367
R2001 B.n1005 B.n436 163.367
R2002 B.n1005 B.n430 163.367
R2003 B.n1013 B.n430 163.367
R2004 B.n1013 B.n428 163.367
R2005 B.n1017 B.n428 163.367
R2006 B.n1017 B.n422 163.367
R2007 B.n1025 B.n422 163.367
R2008 B.n1025 B.n420 163.367
R2009 B.n1029 B.n420 163.367
R2010 B.n1029 B.n415 163.367
R2011 B.n1038 B.n415 163.367
R2012 B.n1038 B.n413 163.367
R2013 B.n1043 B.n413 163.367
R2014 B.n1043 B.n407 163.367
R2015 B.n1051 B.n407 163.367
R2016 B.n1052 B.n1051 163.367
R2017 B.n1052 B.n5 163.367
R2018 B.n6 B.n5 163.367
R2019 B.n7 B.n6 163.367
R2020 B.n1058 B.n7 163.367
R2021 B.n1059 B.n1058 163.367
R2022 B.n1059 B.n13 163.367
R2023 B.n14 B.n13 163.367
R2024 B.n15 B.n14 163.367
R2025 B.n1064 B.n15 163.367
R2026 B.n1064 B.n20 163.367
R2027 B.n21 B.n20 163.367
R2028 B.n22 B.n21 163.367
R2029 B.n1069 B.n22 163.367
R2030 B.n1069 B.n27 163.367
R2031 B.n28 B.n27 163.367
R2032 B.n29 B.n28 163.367
R2033 B.n1074 B.n29 163.367
R2034 B.n1074 B.n34 163.367
R2035 B.n35 B.n34 163.367
R2036 B.n36 B.n35 163.367
R2037 B.n1079 B.n36 163.367
R2038 B.n1079 B.n41 163.367
R2039 B.n42 B.n41 163.367
R2040 B.n43 B.n42 163.367
R2041 B.n1084 B.n43 163.367
R2042 B.n1084 B.n48 163.367
R2043 B.n49 B.n48 163.367
R2044 B.n50 B.n49 163.367
R2045 B.n1089 B.n50 163.367
R2046 B.n1089 B.n55 163.367
R2047 B.n56 B.n55 163.367
R2048 B.n57 B.n56 163.367
R2049 B.n1094 B.n57 163.367
R2050 B.n1094 B.n62 163.367
R2051 B.n63 B.n62 163.367
R2052 B.n64 B.n63 163.367
R2053 B.n1099 B.n64 163.367
R2054 B.n1099 B.n69 163.367
R2055 B.n70 B.n69 163.367
R2056 B.n71 B.n70 163.367
R2057 B.n1104 B.n71 163.367
R2058 B.n1104 B.n76 163.367
R2059 B.n77 B.n76 163.367
R2060 B.n78 B.n77 163.367
R2061 B.n1109 B.n78 163.367
R2062 B.n1109 B.n83 163.367
R2063 B.n84 B.n83 163.367
R2064 B.n85 B.n84 163.367
R2065 B.n1114 B.n85 163.367
R2066 B.n1114 B.n90 163.367
R2067 B.n91 B.n90 163.367
R2068 B.n92 B.n91 163.367
R2069 B.n1119 B.n92 163.367
R2070 B.n1119 B.n97 163.367
R2071 B.n98 B.n97 163.367
R2072 B.n99 B.n98 163.367
R2073 B.n1124 B.n99 163.367
R2074 B.n1124 B.n104 163.367
R2075 B.n105 B.n104 163.367
R2076 B.n106 B.n105 163.367
R2077 B.n1129 B.n106 163.367
R2078 B.n1129 B.n111 163.367
R2079 B.n112 B.n111 163.367
R2080 B.n113 B.n112 163.367
R2081 B.n1134 B.n113 163.367
R2082 B.n1134 B.n118 163.367
R2083 B.n119 B.n118 163.367
R2084 B.n120 B.n119 163.367
R2085 B.n1139 B.n120 163.367
R2086 B.n1139 B.n125 163.367
R2087 B.n126 B.n125 163.367
R2088 B.n127 B.n126 163.367
R2089 B.n1144 B.n127 163.367
R2090 B.n1144 B.n132 163.367
R2091 B.n133 B.n132 163.367
R2092 B.n134 B.n133 163.367
R2093 B.n1149 B.n134 163.367
R2094 B.n1149 B.n139 163.367
R2095 B.n613 B.n612 163.367
R2096 B.n615 B.n613 163.367
R2097 B.n619 B.n608 163.367
R2098 B.n623 B.n621 163.367
R2099 B.n627 B.n606 163.367
R2100 B.n631 B.n629 163.367
R2101 B.n635 B.n604 163.367
R2102 B.n639 B.n637 163.367
R2103 B.n643 B.n602 163.367
R2104 B.n647 B.n645 163.367
R2105 B.n651 B.n600 163.367
R2106 B.n655 B.n653 163.367
R2107 B.n659 B.n598 163.367
R2108 B.n663 B.n661 163.367
R2109 B.n667 B.n596 163.367
R2110 B.n671 B.n669 163.367
R2111 B.n675 B.n594 163.367
R2112 B.n679 B.n677 163.367
R2113 B.n683 B.n592 163.367
R2114 B.n687 B.n685 163.367
R2115 B.n691 B.n590 163.367
R2116 B.n695 B.n693 163.367
R2117 B.n699 B.n588 163.367
R2118 B.n703 B.n701 163.367
R2119 B.n708 B.n584 163.367
R2120 B.n712 B.n710 163.367
R2121 B.n716 B.n582 163.367
R2122 B.n720 B.n718 163.367
R2123 B.n727 B.n580 163.367
R2124 B.n731 B.n729 163.367
R2125 B.n735 B.n578 163.367
R2126 B.n739 B.n737 163.367
R2127 B.n743 B.n576 163.367
R2128 B.n747 B.n745 163.367
R2129 B.n751 B.n574 163.367
R2130 B.n755 B.n753 163.367
R2131 B.n759 B.n572 163.367
R2132 B.n763 B.n761 163.367
R2133 B.n767 B.n570 163.367
R2134 B.n771 B.n769 163.367
R2135 B.n775 B.n568 163.367
R2136 B.n779 B.n777 163.367
R2137 B.n783 B.n566 163.367
R2138 B.n787 B.n785 163.367
R2139 B.n791 B.n564 163.367
R2140 B.n795 B.n793 163.367
R2141 B.n799 B.n562 163.367
R2142 B.n803 B.n801 163.367
R2143 B.n807 B.n560 163.367
R2144 B.n811 B.n809 163.367
R2145 B.n815 B.n558 163.367
R2146 B.n818 B.n817 163.367
R2147 B.n820 B.n555 163.367
R2148 B.n826 B.n551 163.367
R2149 B.n830 B.n551 163.367
R2150 B.n830 B.n545 163.367
R2151 B.n838 B.n545 163.367
R2152 B.n838 B.n543 163.367
R2153 B.n842 B.n543 163.367
R2154 B.n842 B.n537 163.367
R2155 B.n850 B.n537 163.367
R2156 B.n850 B.n535 163.367
R2157 B.n854 B.n535 163.367
R2158 B.n854 B.n529 163.367
R2159 B.n862 B.n529 163.367
R2160 B.n862 B.n527 163.367
R2161 B.n866 B.n527 163.367
R2162 B.n866 B.n521 163.367
R2163 B.n874 B.n521 163.367
R2164 B.n874 B.n519 163.367
R2165 B.n878 B.n519 163.367
R2166 B.n878 B.n513 163.367
R2167 B.n886 B.n513 163.367
R2168 B.n886 B.n511 163.367
R2169 B.n890 B.n511 163.367
R2170 B.n890 B.n505 163.367
R2171 B.n898 B.n505 163.367
R2172 B.n898 B.n503 163.367
R2173 B.n902 B.n503 163.367
R2174 B.n902 B.n497 163.367
R2175 B.n910 B.n497 163.367
R2176 B.n910 B.n495 163.367
R2177 B.n914 B.n495 163.367
R2178 B.n914 B.n489 163.367
R2179 B.n922 B.n489 163.367
R2180 B.n922 B.n487 163.367
R2181 B.n926 B.n487 163.367
R2182 B.n926 B.n481 163.367
R2183 B.n934 B.n481 163.367
R2184 B.n934 B.n479 163.367
R2185 B.n938 B.n479 163.367
R2186 B.n938 B.n473 163.367
R2187 B.n946 B.n473 163.367
R2188 B.n946 B.n471 163.367
R2189 B.n950 B.n471 163.367
R2190 B.n950 B.n465 163.367
R2191 B.n958 B.n465 163.367
R2192 B.n958 B.n463 163.367
R2193 B.n962 B.n463 163.367
R2194 B.n962 B.n457 163.367
R2195 B.n970 B.n457 163.367
R2196 B.n970 B.n455 163.367
R2197 B.n974 B.n455 163.367
R2198 B.n974 B.n449 163.367
R2199 B.n982 B.n449 163.367
R2200 B.n982 B.n447 163.367
R2201 B.n986 B.n447 163.367
R2202 B.n986 B.n441 163.367
R2203 B.n995 B.n441 163.367
R2204 B.n995 B.n439 163.367
R2205 B.n999 B.n439 163.367
R2206 B.n999 B.n434 163.367
R2207 B.n1007 B.n434 163.367
R2208 B.n1007 B.n432 163.367
R2209 B.n1011 B.n432 163.367
R2210 B.n1011 B.n426 163.367
R2211 B.n1019 B.n426 163.367
R2212 B.n1019 B.n424 163.367
R2213 B.n1023 B.n424 163.367
R2214 B.n1023 B.n418 163.367
R2215 B.n1032 B.n418 163.367
R2216 B.n1032 B.n416 163.367
R2217 B.n1036 B.n416 163.367
R2218 B.n1036 B.n411 163.367
R2219 B.n1045 B.n411 163.367
R2220 B.n1045 B.n409 163.367
R2221 B.n1049 B.n409 163.367
R2222 B.n1049 B.n3 163.367
R2223 B.n1310 B.n3 163.367
R2224 B.n1306 B.n2 163.367
R2225 B.n1306 B.n1305 163.367
R2226 B.n1305 B.n9 163.367
R2227 B.n1301 B.n9 163.367
R2228 B.n1301 B.n11 163.367
R2229 B.n1297 B.n11 163.367
R2230 B.n1297 B.n16 163.367
R2231 B.n1293 B.n16 163.367
R2232 B.n1293 B.n18 163.367
R2233 B.n1289 B.n18 163.367
R2234 B.n1289 B.n24 163.367
R2235 B.n1285 B.n24 163.367
R2236 B.n1285 B.n26 163.367
R2237 B.n1281 B.n26 163.367
R2238 B.n1281 B.n31 163.367
R2239 B.n1277 B.n31 163.367
R2240 B.n1277 B.n33 163.367
R2241 B.n1273 B.n33 163.367
R2242 B.n1273 B.n37 163.367
R2243 B.n1269 B.n37 163.367
R2244 B.n1269 B.n39 163.367
R2245 B.n1265 B.n39 163.367
R2246 B.n1265 B.n45 163.367
R2247 B.n1261 B.n45 163.367
R2248 B.n1261 B.n47 163.367
R2249 B.n1257 B.n47 163.367
R2250 B.n1257 B.n52 163.367
R2251 B.n1253 B.n52 163.367
R2252 B.n1253 B.n54 163.367
R2253 B.n1249 B.n54 163.367
R2254 B.n1249 B.n59 163.367
R2255 B.n1245 B.n59 163.367
R2256 B.n1245 B.n61 163.367
R2257 B.n1241 B.n61 163.367
R2258 B.n1241 B.n66 163.367
R2259 B.n1237 B.n66 163.367
R2260 B.n1237 B.n68 163.367
R2261 B.n1233 B.n68 163.367
R2262 B.n1233 B.n73 163.367
R2263 B.n1229 B.n73 163.367
R2264 B.n1229 B.n75 163.367
R2265 B.n1225 B.n75 163.367
R2266 B.n1225 B.n80 163.367
R2267 B.n1221 B.n80 163.367
R2268 B.n1221 B.n82 163.367
R2269 B.n1217 B.n82 163.367
R2270 B.n1217 B.n87 163.367
R2271 B.n1213 B.n87 163.367
R2272 B.n1213 B.n89 163.367
R2273 B.n1209 B.n89 163.367
R2274 B.n1209 B.n94 163.367
R2275 B.n1205 B.n94 163.367
R2276 B.n1205 B.n96 163.367
R2277 B.n1201 B.n96 163.367
R2278 B.n1201 B.n101 163.367
R2279 B.n1197 B.n101 163.367
R2280 B.n1197 B.n103 163.367
R2281 B.n1193 B.n103 163.367
R2282 B.n1193 B.n108 163.367
R2283 B.n1189 B.n108 163.367
R2284 B.n1189 B.n110 163.367
R2285 B.n1185 B.n110 163.367
R2286 B.n1185 B.n115 163.367
R2287 B.n1181 B.n115 163.367
R2288 B.n1181 B.n117 163.367
R2289 B.n1177 B.n117 163.367
R2290 B.n1177 B.n122 163.367
R2291 B.n1173 B.n122 163.367
R2292 B.n1173 B.n124 163.367
R2293 B.n1169 B.n124 163.367
R2294 B.n1169 B.n129 163.367
R2295 B.n1165 B.n129 163.367
R2296 B.n1165 B.n131 163.367
R2297 B.n1161 B.n131 163.367
R2298 B.n1161 B.n136 163.367
R2299 B.n1157 B.n136 163.367
R2300 B.n197 B.n196 75.249
R2301 B.n194 B.n193 75.249
R2302 B.n724 B.n723 75.249
R2303 B.n586 B.n585 75.249
R2304 B.n825 B.n554 72.8631
R2305 B.n1156 B.n1155 72.8631
R2306 B.n140 B.n138 71.676
R2307 B.n201 B.n141 71.676
R2308 B.n205 B.n142 71.676
R2309 B.n209 B.n143 71.676
R2310 B.n213 B.n144 71.676
R2311 B.n217 B.n145 71.676
R2312 B.n221 B.n146 71.676
R2313 B.n225 B.n147 71.676
R2314 B.n229 B.n148 71.676
R2315 B.n233 B.n149 71.676
R2316 B.n237 B.n150 71.676
R2317 B.n241 B.n151 71.676
R2318 B.n245 B.n152 71.676
R2319 B.n249 B.n153 71.676
R2320 B.n253 B.n154 71.676
R2321 B.n257 B.n155 71.676
R2322 B.n261 B.n156 71.676
R2323 B.n265 B.n157 71.676
R2324 B.n269 B.n158 71.676
R2325 B.n273 B.n159 71.676
R2326 B.n277 B.n160 71.676
R2327 B.n281 B.n161 71.676
R2328 B.n285 B.n162 71.676
R2329 B.n289 B.n163 71.676
R2330 B.n293 B.n164 71.676
R2331 B.n297 B.n165 71.676
R2332 B.n301 B.n166 71.676
R2333 B.n305 B.n167 71.676
R2334 B.n309 B.n168 71.676
R2335 B.n313 B.n169 71.676
R2336 B.n317 B.n170 71.676
R2337 B.n321 B.n171 71.676
R2338 B.n325 B.n172 71.676
R2339 B.n329 B.n173 71.676
R2340 B.n333 B.n174 71.676
R2341 B.n337 B.n175 71.676
R2342 B.n341 B.n176 71.676
R2343 B.n345 B.n177 71.676
R2344 B.n349 B.n178 71.676
R2345 B.n353 B.n179 71.676
R2346 B.n357 B.n180 71.676
R2347 B.n361 B.n181 71.676
R2348 B.n365 B.n182 71.676
R2349 B.n369 B.n183 71.676
R2350 B.n373 B.n184 71.676
R2351 B.n377 B.n185 71.676
R2352 B.n381 B.n186 71.676
R2353 B.n385 B.n187 71.676
R2354 B.n389 B.n188 71.676
R2355 B.n393 B.n189 71.676
R2356 B.n397 B.n190 71.676
R2357 B.n401 B.n191 71.676
R2358 B.n1154 B.n192 71.676
R2359 B.n1154 B.n1153 71.676
R2360 B.n403 B.n191 71.676
R2361 B.n400 B.n190 71.676
R2362 B.n396 B.n189 71.676
R2363 B.n392 B.n188 71.676
R2364 B.n388 B.n187 71.676
R2365 B.n384 B.n186 71.676
R2366 B.n380 B.n185 71.676
R2367 B.n376 B.n184 71.676
R2368 B.n372 B.n183 71.676
R2369 B.n368 B.n182 71.676
R2370 B.n364 B.n181 71.676
R2371 B.n360 B.n180 71.676
R2372 B.n356 B.n179 71.676
R2373 B.n352 B.n178 71.676
R2374 B.n348 B.n177 71.676
R2375 B.n344 B.n176 71.676
R2376 B.n340 B.n175 71.676
R2377 B.n336 B.n174 71.676
R2378 B.n332 B.n173 71.676
R2379 B.n328 B.n172 71.676
R2380 B.n324 B.n171 71.676
R2381 B.n320 B.n170 71.676
R2382 B.n316 B.n169 71.676
R2383 B.n312 B.n168 71.676
R2384 B.n308 B.n167 71.676
R2385 B.n304 B.n166 71.676
R2386 B.n300 B.n165 71.676
R2387 B.n296 B.n164 71.676
R2388 B.n292 B.n163 71.676
R2389 B.n288 B.n162 71.676
R2390 B.n284 B.n161 71.676
R2391 B.n280 B.n160 71.676
R2392 B.n276 B.n159 71.676
R2393 B.n272 B.n158 71.676
R2394 B.n268 B.n157 71.676
R2395 B.n264 B.n156 71.676
R2396 B.n260 B.n155 71.676
R2397 B.n256 B.n154 71.676
R2398 B.n252 B.n153 71.676
R2399 B.n248 B.n152 71.676
R2400 B.n244 B.n151 71.676
R2401 B.n240 B.n150 71.676
R2402 B.n236 B.n149 71.676
R2403 B.n232 B.n148 71.676
R2404 B.n228 B.n147 71.676
R2405 B.n224 B.n146 71.676
R2406 B.n220 B.n145 71.676
R2407 B.n216 B.n144 71.676
R2408 B.n212 B.n143 71.676
R2409 B.n208 B.n142 71.676
R2410 B.n204 B.n141 71.676
R2411 B.n200 B.n140 71.676
R2412 B.n611 B.n553 71.676
R2413 B.n615 B.n614 71.676
R2414 B.n620 B.n619 71.676
R2415 B.n623 B.n622 71.676
R2416 B.n628 B.n627 71.676
R2417 B.n631 B.n630 71.676
R2418 B.n636 B.n635 71.676
R2419 B.n639 B.n638 71.676
R2420 B.n644 B.n643 71.676
R2421 B.n647 B.n646 71.676
R2422 B.n652 B.n651 71.676
R2423 B.n655 B.n654 71.676
R2424 B.n660 B.n659 71.676
R2425 B.n663 B.n662 71.676
R2426 B.n668 B.n667 71.676
R2427 B.n671 B.n670 71.676
R2428 B.n676 B.n675 71.676
R2429 B.n679 B.n678 71.676
R2430 B.n684 B.n683 71.676
R2431 B.n687 B.n686 71.676
R2432 B.n692 B.n691 71.676
R2433 B.n695 B.n694 71.676
R2434 B.n700 B.n699 71.676
R2435 B.n703 B.n702 71.676
R2436 B.n709 B.n708 71.676
R2437 B.n712 B.n711 71.676
R2438 B.n717 B.n716 71.676
R2439 B.n720 B.n719 71.676
R2440 B.n728 B.n727 71.676
R2441 B.n731 B.n730 71.676
R2442 B.n736 B.n735 71.676
R2443 B.n739 B.n738 71.676
R2444 B.n744 B.n743 71.676
R2445 B.n747 B.n746 71.676
R2446 B.n752 B.n751 71.676
R2447 B.n755 B.n754 71.676
R2448 B.n760 B.n759 71.676
R2449 B.n763 B.n762 71.676
R2450 B.n768 B.n767 71.676
R2451 B.n771 B.n770 71.676
R2452 B.n776 B.n775 71.676
R2453 B.n779 B.n778 71.676
R2454 B.n784 B.n783 71.676
R2455 B.n787 B.n786 71.676
R2456 B.n792 B.n791 71.676
R2457 B.n795 B.n794 71.676
R2458 B.n800 B.n799 71.676
R2459 B.n803 B.n802 71.676
R2460 B.n808 B.n807 71.676
R2461 B.n811 B.n810 71.676
R2462 B.n816 B.n815 71.676
R2463 B.n819 B.n818 71.676
R2464 B.n612 B.n611 71.676
R2465 B.n614 B.n608 71.676
R2466 B.n621 B.n620 71.676
R2467 B.n622 B.n606 71.676
R2468 B.n629 B.n628 71.676
R2469 B.n630 B.n604 71.676
R2470 B.n637 B.n636 71.676
R2471 B.n638 B.n602 71.676
R2472 B.n645 B.n644 71.676
R2473 B.n646 B.n600 71.676
R2474 B.n653 B.n652 71.676
R2475 B.n654 B.n598 71.676
R2476 B.n661 B.n660 71.676
R2477 B.n662 B.n596 71.676
R2478 B.n669 B.n668 71.676
R2479 B.n670 B.n594 71.676
R2480 B.n677 B.n676 71.676
R2481 B.n678 B.n592 71.676
R2482 B.n685 B.n684 71.676
R2483 B.n686 B.n590 71.676
R2484 B.n693 B.n692 71.676
R2485 B.n694 B.n588 71.676
R2486 B.n701 B.n700 71.676
R2487 B.n702 B.n584 71.676
R2488 B.n710 B.n709 71.676
R2489 B.n711 B.n582 71.676
R2490 B.n718 B.n717 71.676
R2491 B.n719 B.n580 71.676
R2492 B.n729 B.n728 71.676
R2493 B.n730 B.n578 71.676
R2494 B.n737 B.n736 71.676
R2495 B.n738 B.n576 71.676
R2496 B.n745 B.n744 71.676
R2497 B.n746 B.n574 71.676
R2498 B.n753 B.n752 71.676
R2499 B.n754 B.n572 71.676
R2500 B.n761 B.n760 71.676
R2501 B.n762 B.n570 71.676
R2502 B.n769 B.n768 71.676
R2503 B.n770 B.n568 71.676
R2504 B.n777 B.n776 71.676
R2505 B.n778 B.n566 71.676
R2506 B.n785 B.n784 71.676
R2507 B.n786 B.n564 71.676
R2508 B.n793 B.n792 71.676
R2509 B.n794 B.n562 71.676
R2510 B.n801 B.n800 71.676
R2511 B.n802 B.n560 71.676
R2512 B.n809 B.n808 71.676
R2513 B.n810 B.n558 71.676
R2514 B.n817 B.n816 71.676
R2515 B.n820 B.n819 71.676
R2516 B.n1311 B.n1310 71.676
R2517 B.n1311 B.n2 71.676
R2518 B.n198 B.n197 59.5399
R2519 B.n195 B.n194 59.5399
R2520 B.n725 B.n724 59.5399
R2521 B.n705 B.n586 59.5399
R2522 B.n825 B.n550 38.4087
R2523 B.n831 B.n550 38.4087
R2524 B.n831 B.n546 38.4087
R2525 B.n837 B.n546 38.4087
R2526 B.n837 B.n542 38.4087
R2527 B.n843 B.n542 38.4087
R2528 B.n843 B.n538 38.4087
R2529 B.n849 B.n538 38.4087
R2530 B.n855 B.n534 38.4087
R2531 B.n855 B.n530 38.4087
R2532 B.n861 B.n530 38.4087
R2533 B.n861 B.n526 38.4087
R2534 B.n867 B.n526 38.4087
R2535 B.n867 B.n522 38.4087
R2536 B.n873 B.n522 38.4087
R2537 B.n873 B.n518 38.4087
R2538 B.n879 B.n518 38.4087
R2539 B.n879 B.n514 38.4087
R2540 B.n885 B.n514 38.4087
R2541 B.n885 B.n509 38.4087
R2542 B.n891 B.n509 38.4087
R2543 B.n891 B.n510 38.4087
R2544 B.n897 B.n502 38.4087
R2545 B.n903 B.n502 38.4087
R2546 B.n903 B.n498 38.4087
R2547 B.n909 B.n498 38.4087
R2548 B.n909 B.n494 38.4087
R2549 B.n915 B.n494 38.4087
R2550 B.n915 B.n490 38.4087
R2551 B.n921 B.n490 38.4087
R2552 B.n921 B.n486 38.4087
R2553 B.n927 B.n486 38.4087
R2554 B.n933 B.n482 38.4087
R2555 B.n933 B.n478 38.4087
R2556 B.n939 B.n478 38.4087
R2557 B.n939 B.n474 38.4087
R2558 B.n945 B.n474 38.4087
R2559 B.n945 B.n470 38.4087
R2560 B.n951 B.n470 38.4087
R2561 B.n951 B.n466 38.4087
R2562 B.n957 B.n466 38.4087
R2563 B.n957 B.n462 38.4087
R2564 B.n963 B.n462 38.4087
R2565 B.n969 B.n458 38.4087
R2566 B.n969 B.n454 38.4087
R2567 B.n975 B.n454 38.4087
R2568 B.n975 B.n450 38.4087
R2569 B.n981 B.n450 38.4087
R2570 B.n981 B.n446 38.4087
R2571 B.n987 B.n446 38.4087
R2572 B.n987 B.n442 38.4087
R2573 B.n994 B.n442 38.4087
R2574 B.n994 B.n993 38.4087
R2575 B.n1000 B.n435 38.4087
R2576 B.n1006 B.n435 38.4087
R2577 B.n1006 B.n431 38.4087
R2578 B.n1012 B.n431 38.4087
R2579 B.n1012 B.n427 38.4087
R2580 B.n1018 B.n427 38.4087
R2581 B.n1018 B.n423 38.4087
R2582 B.n1024 B.n423 38.4087
R2583 B.n1024 B.n419 38.4087
R2584 B.n1031 B.n419 38.4087
R2585 B.n1031 B.n1030 38.4087
R2586 B.n1037 B.n412 38.4087
R2587 B.n1044 B.n412 38.4087
R2588 B.n1044 B.n408 38.4087
R2589 B.n1050 B.n408 38.4087
R2590 B.n1050 B.n4 38.4087
R2591 B.n1309 B.n4 38.4087
R2592 B.n1309 B.n1308 38.4087
R2593 B.n1308 B.n1307 38.4087
R2594 B.n1307 B.n8 38.4087
R2595 B.n12 B.n8 38.4087
R2596 B.n1300 B.n12 38.4087
R2597 B.n1300 B.n1299 38.4087
R2598 B.n1299 B.n1298 38.4087
R2599 B.n1292 B.n19 38.4087
R2600 B.n1292 B.n1291 38.4087
R2601 B.n1291 B.n1290 38.4087
R2602 B.n1290 B.n23 38.4087
R2603 B.n1284 B.n23 38.4087
R2604 B.n1284 B.n1283 38.4087
R2605 B.n1283 B.n1282 38.4087
R2606 B.n1282 B.n30 38.4087
R2607 B.n1276 B.n30 38.4087
R2608 B.n1276 B.n1275 38.4087
R2609 B.n1275 B.n1274 38.4087
R2610 B.n1268 B.n40 38.4087
R2611 B.n1268 B.n1267 38.4087
R2612 B.n1267 B.n1266 38.4087
R2613 B.n1266 B.n44 38.4087
R2614 B.n1260 B.n44 38.4087
R2615 B.n1260 B.n1259 38.4087
R2616 B.n1259 B.n1258 38.4087
R2617 B.n1258 B.n51 38.4087
R2618 B.n1252 B.n51 38.4087
R2619 B.n1252 B.n1251 38.4087
R2620 B.n1250 B.n58 38.4087
R2621 B.n1244 B.n58 38.4087
R2622 B.n1244 B.n1243 38.4087
R2623 B.n1243 B.n1242 38.4087
R2624 B.n1242 B.n65 38.4087
R2625 B.n1236 B.n65 38.4087
R2626 B.n1236 B.n1235 38.4087
R2627 B.n1235 B.n1234 38.4087
R2628 B.n1234 B.n72 38.4087
R2629 B.n1228 B.n72 38.4087
R2630 B.n1228 B.n1227 38.4087
R2631 B.n1226 B.n79 38.4087
R2632 B.n1220 B.n79 38.4087
R2633 B.n1220 B.n1219 38.4087
R2634 B.n1219 B.n1218 38.4087
R2635 B.n1218 B.n86 38.4087
R2636 B.n1212 B.n86 38.4087
R2637 B.n1212 B.n1211 38.4087
R2638 B.n1211 B.n1210 38.4087
R2639 B.n1210 B.n93 38.4087
R2640 B.n1204 B.n93 38.4087
R2641 B.n1203 B.n1202 38.4087
R2642 B.n1202 B.n100 38.4087
R2643 B.n1196 B.n100 38.4087
R2644 B.n1196 B.n1195 38.4087
R2645 B.n1195 B.n1194 38.4087
R2646 B.n1194 B.n107 38.4087
R2647 B.n1188 B.n107 38.4087
R2648 B.n1188 B.n1187 38.4087
R2649 B.n1187 B.n1186 38.4087
R2650 B.n1186 B.n114 38.4087
R2651 B.n1180 B.n114 38.4087
R2652 B.n1180 B.n1179 38.4087
R2653 B.n1179 B.n1178 38.4087
R2654 B.n1178 B.n121 38.4087
R2655 B.n1172 B.n1171 38.4087
R2656 B.n1171 B.n1170 38.4087
R2657 B.n1170 B.n128 38.4087
R2658 B.n1164 B.n128 38.4087
R2659 B.n1164 B.n1163 38.4087
R2660 B.n1163 B.n1162 38.4087
R2661 B.n1162 B.n135 38.4087
R2662 B.n1156 B.n135 38.4087
R2663 B.n927 B.t4 36.7142
R2664 B.t7 B.n1226 36.7142
R2665 B.n849 B.t15 35.5846
R2666 B.n1172 B.t11 35.5846
R2667 B.n827 B.n552 32.0005
R2668 B.n823 B.n822 32.0005
R2669 B.n1152 B.n1151 32.0005
R2670 B.n1158 B.n137 32.0005
R2671 B.n1037 B.t6 31.066
R2672 B.n1298 B.t2 31.066
R2673 B.n993 B.t1 29.9363
R2674 B.n40 B.t5 29.9363
R2675 B.t3 B.n458 24.288
R2676 B.n1251 B.t9 24.288
R2677 B.n510 B.t8 20.8991
R2678 B.t0 B.n1203 20.8991
R2679 B B.n1312 18.0485
R2680 B.n897 B.t8 17.5101
R2681 B.n1204 B.t0 17.5101
R2682 B.n963 B.t3 14.1212
R2683 B.t9 B.n1250 14.1212
R2684 B.n828 B.n827 10.6151
R2685 B.n829 B.n828 10.6151
R2686 B.n829 B.n544 10.6151
R2687 B.n839 B.n544 10.6151
R2688 B.n840 B.n839 10.6151
R2689 B.n841 B.n840 10.6151
R2690 B.n841 B.n536 10.6151
R2691 B.n851 B.n536 10.6151
R2692 B.n852 B.n851 10.6151
R2693 B.n853 B.n852 10.6151
R2694 B.n853 B.n528 10.6151
R2695 B.n863 B.n528 10.6151
R2696 B.n864 B.n863 10.6151
R2697 B.n865 B.n864 10.6151
R2698 B.n865 B.n520 10.6151
R2699 B.n875 B.n520 10.6151
R2700 B.n876 B.n875 10.6151
R2701 B.n877 B.n876 10.6151
R2702 B.n877 B.n512 10.6151
R2703 B.n887 B.n512 10.6151
R2704 B.n888 B.n887 10.6151
R2705 B.n889 B.n888 10.6151
R2706 B.n889 B.n504 10.6151
R2707 B.n899 B.n504 10.6151
R2708 B.n900 B.n899 10.6151
R2709 B.n901 B.n900 10.6151
R2710 B.n901 B.n496 10.6151
R2711 B.n911 B.n496 10.6151
R2712 B.n912 B.n911 10.6151
R2713 B.n913 B.n912 10.6151
R2714 B.n913 B.n488 10.6151
R2715 B.n923 B.n488 10.6151
R2716 B.n924 B.n923 10.6151
R2717 B.n925 B.n924 10.6151
R2718 B.n925 B.n480 10.6151
R2719 B.n935 B.n480 10.6151
R2720 B.n936 B.n935 10.6151
R2721 B.n937 B.n936 10.6151
R2722 B.n937 B.n472 10.6151
R2723 B.n947 B.n472 10.6151
R2724 B.n948 B.n947 10.6151
R2725 B.n949 B.n948 10.6151
R2726 B.n949 B.n464 10.6151
R2727 B.n959 B.n464 10.6151
R2728 B.n960 B.n959 10.6151
R2729 B.n961 B.n960 10.6151
R2730 B.n961 B.n456 10.6151
R2731 B.n971 B.n456 10.6151
R2732 B.n972 B.n971 10.6151
R2733 B.n973 B.n972 10.6151
R2734 B.n973 B.n448 10.6151
R2735 B.n983 B.n448 10.6151
R2736 B.n984 B.n983 10.6151
R2737 B.n985 B.n984 10.6151
R2738 B.n985 B.n440 10.6151
R2739 B.n996 B.n440 10.6151
R2740 B.n997 B.n996 10.6151
R2741 B.n998 B.n997 10.6151
R2742 B.n998 B.n433 10.6151
R2743 B.n1008 B.n433 10.6151
R2744 B.n1009 B.n1008 10.6151
R2745 B.n1010 B.n1009 10.6151
R2746 B.n1010 B.n425 10.6151
R2747 B.n1020 B.n425 10.6151
R2748 B.n1021 B.n1020 10.6151
R2749 B.n1022 B.n1021 10.6151
R2750 B.n1022 B.n417 10.6151
R2751 B.n1033 B.n417 10.6151
R2752 B.n1034 B.n1033 10.6151
R2753 B.n1035 B.n1034 10.6151
R2754 B.n1035 B.n410 10.6151
R2755 B.n1046 B.n410 10.6151
R2756 B.n1047 B.n1046 10.6151
R2757 B.n1048 B.n1047 10.6151
R2758 B.n1048 B.n0 10.6151
R2759 B.n610 B.n552 10.6151
R2760 B.n610 B.n609 10.6151
R2761 B.n616 B.n609 10.6151
R2762 B.n617 B.n616 10.6151
R2763 B.n618 B.n617 10.6151
R2764 B.n618 B.n607 10.6151
R2765 B.n624 B.n607 10.6151
R2766 B.n625 B.n624 10.6151
R2767 B.n626 B.n625 10.6151
R2768 B.n626 B.n605 10.6151
R2769 B.n632 B.n605 10.6151
R2770 B.n633 B.n632 10.6151
R2771 B.n634 B.n633 10.6151
R2772 B.n634 B.n603 10.6151
R2773 B.n640 B.n603 10.6151
R2774 B.n641 B.n640 10.6151
R2775 B.n642 B.n641 10.6151
R2776 B.n642 B.n601 10.6151
R2777 B.n648 B.n601 10.6151
R2778 B.n649 B.n648 10.6151
R2779 B.n650 B.n649 10.6151
R2780 B.n650 B.n599 10.6151
R2781 B.n656 B.n599 10.6151
R2782 B.n657 B.n656 10.6151
R2783 B.n658 B.n657 10.6151
R2784 B.n658 B.n597 10.6151
R2785 B.n664 B.n597 10.6151
R2786 B.n665 B.n664 10.6151
R2787 B.n666 B.n665 10.6151
R2788 B.n666 B.n595 10.6151
R2789 B.n672 B.n595 10.6151
R2790 B.n673 B.n672 10.6151
R2791 B.n674 B.n673 10.6151
R2792 B.n674 B.n593 10.6151
R2793 B.n680 B.n593 10.6151
R2794 B.n681 B.n680 10.6151
R2795 B.n682 B.n681 10.6151
R2796 B.n682 B.n591 10.6151
R2797 B.n688 B.n591 10.6151
R2798 B.n689 B.n688 10.6151
R2799 B.n690 B.n689 10.6151
R2800 B.n690 B.n589 10.6151
R2801 B.n696 B.n589 10.6151
R2802 B.n697 B.n696 10.6151
R2803 B.n698 B.n697 10.6151
R2804 B.n698 B.n587 10.6151
R2805 B.n704 B.n587 10.6151
R2806 B.n707 B.n706 10.6151
R2807 B.n707 B.n583 10.6151
R2808 B.n713 B.n583 10.6151
R2809 B.n714 B.n713 10.6151
R2810 B.n715 B.n714 10.6151
R2811 B.n715 B.n581 10.6151
R2812 B.n721 B.n581 10.6151
R2813 B.n722 B.n721 10.6151
R2814 B.n726 B.n722 10.6151
R2815 B.n732 B.n579 10.6151
R2816 B.n733 B.n732 10.6151
R2817 B.n734 B.n733 10.6151
R2818 B.n734 B.n577 10.6151
R2819 B.n740 B.n577 10.6151
R2820 B.n741 B.n740 10.6151
R2821 B.n742 B.n741 10.6151
R2822 B.n742 B.n575 10.6151
R2823 B.n748 B.n575 10.6151
R2824 B.n749 B.n748 10.6151
R2825 B.n750 B.n749 10.6151
R2826 B.n750 B.n573 10.6151
R2827 B.n756 B.n573 10.6151
R2828 B.n757 B.n756 10.6151
R2829 B.n758 B.n757 10.6151
R2830 B.n758 B.n571 10.6151
R2831 B.n764 B.n571 10.6151
R2832 B.n765 B.n764 10.6151
R2833 B.n766 B.n765 10.6151
R2834 B.n766 B.n569 10.6151
R2835 B.n772 B.n569 10.6151
R2836 B.n773 B.n772 10.6151
R2837 B.n774 B.n773 10.6151
R2838 B.n774 B.n567 10.6151
R2839 B.n780 B.n567 10.6151
R2840 B.n781 B.n780 10.6151
R2841 B.n782 B.n781 10.6151
R2842 B.n782 B.n565 10.6151
R2843 B.n788 B.n565 10.6151
R2844 B.n789 B.n788 10.6151
R2845 B.n790 B.n789 10.6151
R2846 B.n790 B.n563 10.6151
R2847 B.n796 B.n563 10.6151
R2848 B.n797 B.n796 10.6151
R2849 B.n798 B.n797 10.6151
R2850 B.n798 B.n561 10.6151
R2851 B.n804 B.n561 10.6151
R2852 B.n805 B.n804 10.6151
R2853 B.n806 B.n805 10.6151
R2854 B.n806 B.n559 10.6151
R2855 B.n812 B.n559 10.6151
R2856 B.n813 B.n812 10.6151
R2857 B.n814 B.n813 10.6151
R2858 B.n814 B.n557 10.6151
R2859 B.n557 B.n556 10.6151
R2860 B.n821 B.n556 10.6151
R2861 B.n822 B.n821 10.6151
R2862 B.n823 B.n548 10.6151
R2863 B.n833 B.n548 10.6151
R2864 B.n834 B.n833 10.6151
R2865 B.n835 B.n834 10.6151
R2866 B.n835 B.n540 10.6151
R2867 B.n845 B.n540 10.6151
R2868 B.n846 B.n845 10.6151
R2869 B.n847 B.n846 10.6151
R2870 B.n847 B.n532 10.6151
R2871 B.n857 B.n532 10.6151
R2872 B.n858 B.n857 10.6151
R2873 B.n859 B.n858 10.6151
R2874 B.n859 B.n524 10.6151
R2875 B.n869 B.n524 10.6151
R2876 B.n870 B.n869 10.6151
R2877 B.n871 B.n870 10.6151
R2878 B.n871 B.n516 10.6151
R2879 B.n881 B.n516 10.6151
R2880 B.n882 B.n881 10.6151
R2881 B.n883 B.n882 10.6151
R2882 B.n883 B.n507 10.6151
R2883 B.n893 B.n507 10.6151
R2884 B.n894 B.n893 10.6151
R2885 B.n895 B.n894 10.6151
R2886 B.n895 B.n500 10.6151
R2887 B.n905 B.n500 10.6151
R2888 B.n906 B.n905 10.6151
R2889 B.n907 B.n906 10.6151
R2890 B.n907 B.n492 10.6151
R2891 B.n917 B.n492 10.6151
R2892 B.n918 B.n917 10.6151
R2893 B.n919 B.n918 10.6151
R2894 B.n919 B.n484 10.6151
R2895 B.n929 B.n484 10.6151
R2896 B.n930 B.n929 10.6151
R2897 B.n931 B.n930 10.6151
R2898 B.n931 B.n476 10.6151
R2899 B.n941 B.n476 10.6151
R2900 B.n942 B.n941 10.6151
R2901 B.n943 B.n942 10.6151
R2902 B.n943 B.n468 10.6151
R2903 B.n953 B.n468 10.6151
R2904 B.n954 B.n953 10.6151
R2905 B.n955 B.n954 10.6151
R2906 B.n955 B.n460 10.6151
R2907 B.n965 B.n460 10.6151
R2908 B.n966 B.n965 10.6151
R2909 B.n967 B.n966 10.6151
R2910 B.n967 B.n452 10.6151
R2911 B.n977 B.n452 10.6151
R2912 B.n978 B.n977 10.6151
R2913 B.n979 B.n978 10.6151
R2914 B.n979 B.n444 10.6151
R2915 B.n989 B.n444 10.6151
R2916 B.n990 B.n989 10.6151
R2917 B.n991 B.n990 10.6151
R2918 B.n991 B.n437 10.6151
R2919 B.n1002 B.n437 10.6151
R2920 B.n1003 B.n1002 10.6151
R2921 B.n1004 B.n1003 10.6151
R2922 B.n1004 B.n429 10.6151
R2923 B.n1014 B.n429 10.6151
R2924 B.n1015 B.n1014 10.6151
R2925 B.n1016 B.n1015 10.6151
R2926 B.n1016 B.n421 10.6151
R2927 B.n1026 B.n421 10.6151
R2928 B.n1027 B.n1026 10.6151
R2929 B.n1028 B.n1027 10.6151
R2930 B.n1028 B.n414 10.6151
R2931 B.n1039 B.n414 10.6151
R2932 B.n1040 B.n1039 10.6151
R2933 B.n1042 B.n1040 10.6151
R2934 B.n1042 B.n1041 10.6151
R2935 B.n1041 B.n406 10.6151
R2936 B.n1053 B.n406 10.6151
R2937 B.n1054 B.n1053 10.6151
R2938 B.n1055 B.n1054 10.6151
R2939 B.n1056 B.n1055 10.6151
R2940 B.n1057 B.n1056 10.6151
R2941 B.n1060 B.n1057 10.6151
R2942 B.n1061 B.n1060 10.6151
R2943 B.n1062 B.n1061 10.6151
R2944 B.n1063 B.n1062 10.6151
R2945 B.n1065 B.n1063 10.6151
R2946 B.n1066 B.n1065 10.6151
R2947 B.n1067 B.n1066 10.6151
R2948 B.n1068 B.n1067 10.6151
R2949 B.n1070 B.n1068 10.6151
R2950 B.n1071 B.n1070 10.6151
R2951 B.n1072 B.n1071 10.6151
R2952 B.n1073 B.n1072 10.6151
R2953 B.n1075 B.n1073 10.6151
R2954 B.n1076 B.n1075 10.6151
R2955 B.n1077 B.n1076 10.6151
R2956 B.n1078 B.n1077 10.6151
R2957 B.n1080 B.n1078 10.6151
R2958 B.n1081 B.n1080 10.6151
R2959 B.n1082 B.n1081 10.6151
R2960 B.n1083 B.n1082 10.6151
R2961 B.n1085 B.n1083 10.6151
R2962 B.n1086 B.n1085 10.6151
R2963 B.n1087 B.n1086 10.6151
R2964 B.n1088 B.n1087 10.6151
R2965 B.n1090 B.n1088 10.6151
R2966 B.n1091 B.n1090 10.6151
R2967 B.n1092 B.n1091 10.6151
R2968 B.n1093 B.n1092 10.6151
R2969 B.n1095 B.n1093 10.6151
R2970 B.n1096 B.n1095 10.6151
R2971 B.n1097 B.n1096 10.6151
R2972 B.n1098 B.n1097 10.6151
R2973 B.n1100 B.n1098 10.6151
R2974 B.n1101 B.n1100 10.6151
R2975 B.n1102 B.n1101 10.6151
R2976 B.n1103 B.n1102 10.6151
R2977 B.n1105 B.n1103 10.6151
R2978 B.n1106 B.n1105 10.6151
R2979 B.n1107 B.n1106 10.6151
R2980 B.n1108 B.n1107 10.6151
R2981 B.n1110 B.n1108 10.6151
R2982 B.n1111 B.n1110 10.6151
R2983 B.n1112 B.n1111 10.6151
R2984 B.n1113 B.n1112 10.6151
R2985 B.n1115 B.n1113 10.6151
R2986 B.n1116 B.n1115 10.6151
R2987 B.n1117 B.n1116 10.6151
R2988 B.n1118 B.n1117 10.6151
R2989 B.n1120 B.n1118 10.6151
R2990 B.n1121 B.n1120 10.6151
R2991 B.n1122 B.n1121 10.6151
R2992 B.n1123 B.n1122 10.6151
R2993 B.n1125 B.n1123 10.6151
R2994 B.n1126 B.n1125 10.6151
R2995 B.n1127 B.n1126 10.6151
R2996 B.n1128 B.n1127 10.6151
R2997 B.n1130 B.n1128 10.6151
R2998 B.n1131 B.n1130 10.6151
R2999 B.n1132 B.n1131 10.6151
R3000 B.n1133 B.n1132 10.6151
R3001 B.n1135 B.n1133 10.6151
R3002 B.n1136 B.n1135 10.6151
R3003 B.n1137 B.n1136 10.6151
R3004 B.n1138 B.n1137 10.6151
R3005 B.n1140 B.n1138 10.6151
R3006 B.n1141 B.n1140 10.6151
R3007 B.n1142 B.n1141 10.6151
R3008 B.n1143 B.n1142 10.6151
R3009 B.n1145 B.n1143 10.6151
R3010 B.n1146 B.n1145 10.6151
R3011 B.n1147 B.n1146 10.6151
R3012 B.n1148 B.n1147 10.6151
R3013 B.n1150 B.n1148 10.6151
R3014 B.n1151 B.n1150 10.6151
R3015 B.n1304 B.n1 10.6151
R3016 B.n1304 B.n1303 10.6151
R3017 B.n1303 B.n1302 10.6151
R3018 B.n1302 B.n10 10.6151
R3019 B.n1296 B.n10 10.6151
R3020 B.n1296 B.n1295 10.6151
R3021 B.n1295 B.n1294 10.6151
R3022 B.n1294 B.n17 10.6151
R3023 B.n1288 B.n17 10.6151
R3024 B.n1288 B.n1287 10.6151
R3025 B.n1287 B.n1286 10.6151
R3026 B.n1286 B.n25 10.6151
R3027 B.n1280 B.n25 10.6151
R3028 B.n1280 B.n1279 10.6151
R3029 B.n1279 B.n1278 10.6151
R3030 B.n1278 B.n32 10.6151
R3031 B.n1272 B.n32 10.6151
R3032 B.n1272 B.n1271 10.6151
R3033 B.n1271 B.n1270 10.6151
R3034 B.n1270 B.n38 10.6151
R3035 B.n1264 B.n38 10.6151
R3036 B.n1264 B.n1263 10.6151
R3037 B.n1263 B.n1262 10.6151
R3038 B.n1262 B.n46 10.6151
R3039 B.n1256 B.n46 10.6151
R3040 B.n1256 B.n1255 10.6151
R3041 B.n1255 B.n1254 10.6151
R3042 B.n1254 B.n53 10.6151
R3043 B.n1248 B.n53 10.6151
R3044 B.n1248 B.n1247 10.6151
R3045 B.n1247 B.n1246 10.6151
R3046 B.n1246 B.n60 10.6151
R3047 B.n1240 B.n60 10.6151
R3048 B.n1240 B.n1239 10.6151
R3049 B.n1239 B.n1238 10.6151
R3050 B.n1238 B.n67 10.6151
R3051 B.n1232 B.n67 10.6151
R3052 B.n1232 B.n1231 10.6151
R3053 B.n1231 B.n1230 10.6151
R3054 B.n1230 B.n74 10.6151
R3055 B.n1224 B.n74 10.6151
R3056 B.n1224 B.n1223 10.6151
R3057 B.n1223 B.n1222 10.6151
R3058 B.n1222 B.n81 10.6151
R3059 B.n1216 B.n81 10.6151
R3060 B.n1216 B.n1215 10.6151
R3061 B.n1215 B.n1214 10.6151
R3062 B.n1214 B.n88 10.6151
R3063 B.n1208 B.n88 10.6151
R3064 B.n1208 B.n1207 10.6151
R3065 B.n1207 B.n1206 10.6151
R3066 B.n1206 B.n95 10.6151
R3067 B.n1200 B.n95 10.6151
R3068 B.n1200 B.n1199 10.6151
R3069 B.n1199 B.n1198 10.6151
R3070 B.n1198 B.n102 10.6151
R3071 B.n1192 B.n102 10.6151
R3072 B.n1192 B.n1191 10.6151
R3073 B.n1191 B.n1190 10.6151
R3074 B.n1190 B.n109 10.6151
R3075 B.n1184 B.n109 10.6151
R3076 B.n1184 B.n1183 10.6151
R3077 B.n1183 B.n1182 10.6151
R3078 B.n1182 B.n116 10.6151
R3079 B.n1176 B.n116 10.6151
R3080 B.n1176 B.n1175 10.6151
R3081 B.n1175 B.n1174 10.6151
R3082 B.n1174 B.n123 10.6151
R3083 B.n1168 B.n123 10.6151
R3084 B.n1168 B.n1167 10.6151
R3085 B.n1167 B.n1166 10.6151
R3086 B.n1166 B.n130 10.6151
R3087 B.n1160 B.n130 10.6151
R3088 B.n1160 B.n1159 10.6151
R3089 B.n1159 B.n1158 10.6151
R3090 B.n199 B.n137 10.6151
R3091 B.n202 B.n199 10.6151
R3092 B.n203 B.n202 10.6151
R3093 B.n206 B.n203 10.6151
R3094 B.n207 B.n206 10.6151
R3095 B.n210 B.n207 10.6151
R3096 B.n211 B.n210 10.6151
R3097 B.n214 B.n211 10.6151
R3098 B.n215 B.n214 10.6151
R3099 B.n218 B.n215 10.6151
R3100 B.n219 B.n218 10.6151
R3101 B.n222 B.n219 10.6151
R3102 B.n223 B.n222 10.6151
R3103 B.n226 B.n223 10.6151
R3104 B.n227 B.n226 10.6151
R3105 B.n230 B.n227 10.6151
R3106 B.n231 B.n230 10.6151
R3107 B.n234 B.n231 10.6151
R3108 B.n235 B.n234 10.6151
R3109 B.n238 B.n235 10.6151
R3110 B.n239 B.n238 10.6151
R3111 B.n242 B.n239 10.6151
R3112 B.n243 B.n242 10.6151
R3113 B.n246 B.n243 10.6151
R3114 B.n247 B.n246 10.6151
R3115 B.n250 B.n247 10.6151
R3116 B.n251 B.n250 10.6151
R3117 B.n254 B.n251 10.6151
R3118 B.n255 B.n254 10.6151
R3119 B.n258 B.n255 10.6151
R3120 B.n259 B.n258 10.6151
R3121 B.n262 B.n259 10.6151
R3122 B.n263 B.n262 10.6151
R3123 B.n266 B.n263 10.6151
R3124 B.n267 B.n266 10.6151
R3125 B.n270 B.n267 10.6151
R3126 B.n271 B.n270 10.6151
R3127 B.n274 B.n271 10.6151
R3128 B.n275 B.n274 10.6151
R3129 B.n278 B.n275 10.6151
R3130 B.n279 B.n278 10.6151
R3131 B.n282 B.n279 10.6151
R3132 B.n283 B.n282 10.6151
R3133 B.n286 B.n283 10.6151
R3134 B.n287 B.n286 10.6151
R3135 B.n290 B.n287 10.6151
R3136 B.n291 B.n290 10.6151
R3137 B.n295 B.n294 10.6151
R3138 B.n298 B.n295 10.6151
R3139 B.n299 B.n298 10.6151
R3140 B.n302 B.n299 10.6151
R3141 B.n303 B.n302 10.6151
R3142 B.n306 B.n303 10.6151
R3143 B.n307 B.n306 10.6151
R3144 B.n310 B.n307 10.6151
R3145 B.n311 B.n310 10.6151
R3146 B.n315 B.n314 10.6151
R3147 B.n318 B.n315 10.6151
R3148 B.n319 B.n318 10.6151
R3149 B.n322 B.n319 10.6151
R3150 B.n323 B.n322 10.6151
R3151 B.n326 B.n323 10.6151
R3152 B.n327 B.n326 10.6151
R3153 B.n330 B.n327 10.6151
R3154 B.n331 B.n330 10.6151
R3155 B.n334 B.n331 10.6151
R3156 B.n335 B.n334 10.6151
R3157 B.n338 B.n335 10.6151
R3158 B.n339 B.n338 10.6151
R3159 B.n342 B.n339 10.6151
R3160 B.n343 B.n342 10.6151
R3161 B.n346 B.n343 10.6151
R3162 B.n347 B.n346 10.6151
R3163 B.n350 B.n347 10.6151
R3164 B.n351 B.n350 10.6151
R3165 B.n354 B.n351 10.6151
R3166 B.n355 B.n354 10.6151
R3167 B.n358 B.n355 10.6151
R3168 B.n359 B.n358 10.6151
R3169 B.n362 B.n359 10.6151
R3170 B.n363 B.n362 10.6151
R3171 B.n366 B.n363 10.6151
R3172 B.n367 B.n366 10.6151
R3173 B.n370 B.n367 10.6151
R3174 B.n371 B.n370 10.6151
R3175 B.n374 B.n371 10.6151
R3176 B.n375 B.n374 10.6151
R3177 B.n378 B.n375 10.6151
R3178 B.n379 B.n378 10.6151
R3179 B.n382 B.n379 10.6151
R3180 B.n383 B.n382 10.6151
R3181 B.n386 B.n383 10.6151
R3182 B.n387 B.n386 10.6151
R3183 B.n390 B.n387 10.6151
R3184 B.n391 B.n390 10.6151
R3185 B.n394 B.n391 10.6151
R3186 B.n395 B.n394 10.6151
R3187 B.n398 B.n395 10.6151
R3188 B.n399 B.n398 10.6151
R3189 B.n402 B.n399 10.6151
R3190 B.n404 B.n402 10.6151
R3191 B.n405 B.n404 10.6151
R3192 B.n1152 B.n405 10.6151
R3193 B.n705 B.n704 9.36635
R3194 B.n725 B.n579 9.36635
R3195 B.n291 B.n198 9.36635
R3196 B.n314 B.n195 9.36635
R3197 B.n1000 B.t1 8.4729
R3198 B.n1274 B.t5 8.4729
R3199 B.n1312 B.n0 8.11757
R3200 B.n1312 B.n1 8.11757
R3201 B.n1030 B.t6 7.34325
R3202 B.n19 B.t2 7.34325
R3203 B.t15 B.n534 2.82463
R3204 B.t11 B.n121 2.82463
R3205 B.t4 B.n482 1.69498
R3206 B.n1227 B.t7 1.69498
R3207 B.n706 B.n705 1.24928
R3208 B.n726 B.n725 1.24928
R3209 B.n294 B.n198 1.24928
R3210 B.n311 B.n195 1.24928
R3211 VN.n100 VN.n99 161.3
R3212 VN.n98 VN.n52 161.3
R3213 VN.n97 VN.n96 161.3
R3214 VN.n95 VN.n53 161.3
R3215 VN.n94 VN.n93 161.3
R3216 VN.n92 VN.n54 161.3
R3217 VN.n91 VN.n90 161.3
R3218 VN.n89 VN.n55 161.3
R3219 VN.n88 VN.n87 161.3
R3220 VN.n86 VN.n56 161.3
R3221 VN.n85 VN.n84 161.3
R3222 VN.n83 VN.n58 161.3
R3223 VN.n82 VN.n81 161.3
R3224 VN.n80 VN.n59 161.3
R3225 VN.n79 VN.n78 161.3
R3226 VN.n77 VN.n60 161.3
R3227 VN.n76 VN.n75 161.3
R3228 VN.n74 VN.n61 161.3
R3229 VN.n73 VN.n72 161.3
R3230 VN.n71 VN.n62 161.3
R3231 VN.n70 VN.n69 161.3
R3232 VN.n68 VN.n63 161.3
R3233 VN.n67 VN.n66 161.3
R3234 VN.n49 VN.n48 161.3
R3235 VN.n47 VN.n1 161.3
R3236 VN.n46 VN.n45 161.3
R3237 VN.n44 VN.n2 161.3
R3238 VN.n43 VN.n42 161.3
R3239 VN.n41 VN.n3 161.3
R3240 VN.n40 VN.n39 161.3
R3241 VN.n38 VN.n4 161.3
R3242 VN.n37 VN.n36 161.3
R3243 VN.n34 VN.n5 161.3
R3244 VN.n33 VN.n32 161.3
R3245 VN.n31 VN.n6 161.3
R3246 VN.n30 VN.n29 161.3
R3247 VN.n28 VN.n7 161.3
R3248 VN.n27 VN.n26 161.3
R3249 VN.n25 VN.n8 161.3
R3250 VN.n24 VN.n23 161.3
R3251 VN.n22 VN.n9 161.3
R3252 VN.n21 VN.n20 161.3
R3253 VN.n19 VN.n10 161.3
R3254 VN.n18 VN.n17 161.3
R3255 VN.n16 VN.n11 161.3
R3256 VN.n15 VN.n14 161.3
R3257 VN.n65 VN.t6 130.255
R3258 VN.n13 VN.t5 130.255
R3259 VN.n8 VN.t8 96.4005
R3260 VN.n12 VN.t9 96.4005
R3261 VN.n35 VN.t3 96.4005
R3262 VN.n0 VN.t2 96.4005
R3263 VN.n60 VN.t1 96.4005
R3264 VN.n64 VN.t0 96.4005
R3265 VN.n57 VN.t4 96.4005
R3266 VN.n51 VN.t7 96.4005
R3267 VN.n50 VN.n0 77.4578
R3268 VN.n101 VN.n51 77.4578
R3269 VN VN.n101 60.2557
R3270 VN.n42 VN.n2 56.5617
R3271 VN.n93 VN.n53 56.5617
R3272 VN.n13 VN.n12 56.2361
R3273 VN.n65 VN.n64 56.2361
R3274 VN.n21 VN.n10 46.3896
R3275 VN.n29 VN.n6 46.3896
R3276 VN.n73 VN.n62 46.3896
R3277 VN.n81 VN.n58 46.3896
R3278 VN.n17 VN.n10 34.7644
R3279 VN.n33 VN.n6 34.7644
R3280 VN.n69 VN.n62 34.7644
R3281 VN.n85 VN.n58 34.7644
R3282 VN.n16 VN.n15 24.5923
R3283 VN.n17 VN.n16 24.5923
R3284 VN.n22 VN.n21 24.5923
R3285 VN.n23 VN.n22 24.5923
R3286 VN.n23 VN.n8 24.5923
R3287 VN.n27 VN.n8 24.5923
R3288 VN.n28 VN.n27 24.5923
R3289 VN.n29 VN.n28 24.5923
R3290 VN.n34 VN.n33 24.5923
R3291 VN.n36 VN.n34 24.5923
R3292 VN.n40 VN.n4 24.5923
R3293 VN.n41 VN.n40 24.5923
R3294 VN.n42 VN.n41 24.5923
R3295 VN.n46 VN.n2 24.5923
R3296 VN.n47 VN.n46 24.5923
R3297 VN.n48 VN.n47 24.5923
R3298 VN.n69 VN.n68 24.5923
R3299 VN.n68 VN.n67 24.5923
R3300 VN.n81 VN.n80 24.5923
R3301 VN.n80 VN.n79 24.5923
R3302 VN.n79 VN.n60 24.5923
R3303 VN.n75 VN.n60 24.5923
R3304 VN.n75 VN.n74 24.5923
R3305 VN.n74 VN.n73 24.5923
R3306 VN.n93 VN.n92 24.5923
R3307 VN.n92 VN.n91 24.5923
R3308 VN.n91 VN.n55 24.5923
R3309 VN.n87 VN.n86 24.5923
R3310 VN.n86 VN.n85 24.5923
R3311 VN.n99 VN.n98 24.5923
R3312 VN.n98 VN.n97 24.5923
R3313 VN.n97 VN.n53 24.5923
R3314 VN.n15 VN.n12 18.6903
R3315 VN.n36 VN.n35 18.6903
R3316 VN.n67 VN.n64 18.6903
R3317 VN.n87 VN.n57 18.6903
R3318 VN.n48 VN.n0 12.7883
R3319 VN.n99 VN.n51 12.7883
R3320 VN.n35 VN.n4 5.90254
R3321 VN.n57 VN.n55 5.90254
R3322 VN.n66 VN.n65 3.05549
R3323 VN.n14 VN.n13 3.05549
R3324 VN.n101 VN.n100 0.354861
R3325 VN.n50 VN.n49 0.354861
R3326 VN VN.n50 0.267071
R3327 VN.n100 VN.n52 0.189894
R3328 VN.n96 VN.n52 0.189894
R3329 VN.n96 VN.n95 0.189894
R3330 VN.n95 VN.n94 0.189894
R3331 VN.n94 VN.n54 0.189894
R3332 VN.n90 VN.n54 0.189894
R3333 VN.n90 VN.n89 0.189894
R3334 VN.n89 VN.n88 0.189894
R3335 VN.n88 VN.n56 0.189894
R3336 VN.n84 VN.n56 0.189894
R3337 VN.n84 VN.n83 0.189894
R3338 VN.n83 VN.n82 0.189894
R3339 VN.n82 VN.n59 0.189894
R3340 VN.n78 VN.n59 0.189894
R3341 VN.n78 VN.n77 0.189894
R3342 VN.n77 VN.n76 0.189894
R3343 VN.n76 VN.n61 0.189894
R3344 VN.n72 VN.n61 0.189894
R3345 VN.n72 VN.n71 0.189894
R3346 VN.n71 VN.n70 0.189894
R3347 VN.n70 VN.n63 0.189894
R3348 VN.n66 VN.n63 0.189894
R3349 VN.n14 VN.n11 0.189894
R3350 VN.n18 VN.n11 0.189894
R3351 VN.n19 VN.n18 0.189894
R3352 VN.n20 VN.n19 0.189894
R3353 VN.n20 VN.n9 0.189894
R3354 VN.n24 VN.n9 0.189894
R3355 VN.n25 VN.n24 0.189894
R3356 VN.n26 VN.n25 0.189894
R3357 VN.n26 VN.n7 0.189894
R3358 VN.n30 VN.n7 0.189894
R3359 VN.n31 VN.n30 0.189894
R3360 VN.n32 VN.n31 0.189894
R3361 VN.n32 VN.n5 0.189894
R3362 VN.n37 VN.n5 0.189894
R3363 VN.n38 VN.n37 0.189894
R3364 VN.n39 VN.n38 0.189894
R3365 VN.n39 VN.n3 0.189894
R3366 VN.n43 VN.n3 0.189894
R3367 VN.n44 VN.n43 0.189894
R3368 VN.n45 VN.n44 0.189894
R3369 VN.n45 VN.n1 0.189894
R3370 VN.n49 VN.n1 0.189894
R3371 VDD2.n153 VDD2.n81 289.615
R3372 VDD2.n72 VDD2.n0 289.615
R3373 VDD2.n154 VDD2.n153 185
R3374 VDD2.n152 VDD2.n151 185
R3375 VDD2.n85 VDD2.n84 185
R3376 VDD2.n146 VDD2.n145 185
R3377 VDD2.n144 VDD2.n143 185
R3378 VDD2.n89 VDD2.n88 185
R3379 VDD2.n138 VDD2.n137 185
R3380 VDD2.n136 VDD2.n135 185
R3381 VDD2.n93 VDD2.n92 185
R3382 VDD2.n130 VDD2.n129 185
R3383 VDD2.n128 VDD2.n95 185
R3384 VDD2.n127 VDD2.n126 185
R3385 VDD2.n98 VDD2.n96 185
R3386 VDD2.n121 VDD2.n120 185
R3387 VDD2.n119 VDD2.n118 185
R3388 VDD2.n102 VDD2.n101 185
R3389 VDD2.n113 VDD2.n112 185
R3390 VDD2.n111 VDD2.n110 185
R3391 VDD2.n106 VDD2.n105 185
R3392 VDD2.n24 VDD2.n23 185
R3393 VDD2.n29 VDD2.n28 185
R3394 VDD2.n31 VDD2.n30 185
R3395 VDD2.n20 VDD2.n19 185
R3396 VDD2.n37 VDD2.n36 185
R3397 VDD2.n39 VDD2.n38 185
R3398 VDD2.n16 VDD2.n15 185
R3399 VDD2.n46 VDD2.n45 185
R3400 VDD2.n47 VDD2.n14 185
R3401 VDD2.n49 VDD2.n48 185
R3402 VDD2.n12 VDD2.n11 185
R3403 VDD2.n55 VDD2.n54 185
R3404 VDD2.n57 VDD2.n56 185
R3405 VDD2.n8 VDD2.n7 185
R3406 VDD2.n63 VDD2.n62 185
R3407 VDD2.n65 VDD2.n64 185
R3408 VDD2.n4 VDD2.n3 185
R3409 VDD2.n71 VDD2.n70 185
R3410 VDD2.n73 VDD2.n72 185
R3411 VDD2.n107 VDD2.t2 149.524
R3412 VDD2.n25 VDD2.t4 149.524
R3413 VDD2.n153 VDD2.n152 104.615
R3414 VDD2.n152 VDD2.n84 104.615
R3415 VDD2.n145 VDD2.n84 104.615
R3416 VDD2.n145 VDD2.n144 104.615
R3417 VDD2.n144 VDD2.n88 104.615
R3418 VDD2.n137 VDD2.n88 104.615
R3419 VDD2.n137 VDD2.n136 104.615
R3420 VDD2.n136 VDD2.n92 104.615
R3421 VDD2.n129 VDD2.n92 104.615
R3422 VDD2.n129 VDD2.n128 104.615
R3423 VDD2.n128 VDD2.n127 104.615
R3424 VDD2.n127 VDD2.n96 104.615
R3425 VDD2.n120 VDD2.n96 104.615
R3426 VDD2.n120 VDD2.n119 104.615
R3427 VDD2.n119 VDD2.n101 104.615
R3428 VDD2.n112 VDD2.n101 104.615
R3429 VDD2.n112 VDD2.n111 104.615
R3430 VDD2.n111 VDD2.n105 104.615
R3431 VDD2.n29 VDD2.n23 104.615
R3432 VDD2.n30 VDD2.n29 104.615
R3433 VDD2.n30 VDD2.n19 104.615
R3434 VDD2.n37 VDD2.n19 104.615
R3435 VDD2.n38 VDD2.n37 104.615
R3436 VDD2.n38 VDD2.n15 104.615
R3437 VDD2.n46 VDD2.n15 104.615
R3438 VDD2.n47 VDD2.n46 104.615
R3439 VDD2.n48 VDD2.n47 104.615
R3440 VDD2.n48 VDD2.n11 104.615
R3441 VDD2.n55 VDD2.n11 104.615
R3442 VDD2.n56 VDD2.n55 104.615
R3443 VDD2.n56 VDD2.n7 104.615
R3444 VDD2.n63 VDD2.n7 104.615
R3445 VDD2.n64 VDD2.n63 104.615
R3446 VDD2.n64 VDD2.n3 104.615
R3447 VDD2.n71 VDD2.n3 104.615
R3448 VDD2.n72 VDD2.n71 104.615
R3449 VDD2.n80 VDD2.n79 62.3299
R3450 VDD2 VDD2.n161 62.3271
R3451 VDD2.n160 VDD2.n159 59.8767
R3452 VDD2.n78 VDD2.n77 59.8767
R3453 VDD2.t2 VDD2.n105 52.3082
R3454 VDD2.t4 VDD2.n23 52.3082
R3455 VDD2.n158 VDD2.n80 51.8446
R3456 VDD2.n78 VDD2.n76 50.6574
R3457 VDD2.n158 VDD2.n157 47.3126
R3458 VDD2.n130 VDD2.n95 13.1884
R3459 VDD2.n49 VDD2.n14 13.1884
R3460 VDD2.n131 VDD2.n93 12.8005
R3461 VDD2.n126 VDD2.n97 12.8005
R3462 VDD2.n45 VDD2.n44 12.8005
R3463 VDD2.n50 VDD2.n12 12.8005
R3464 VDD2.n135 VDD2.n134 12.0247
R3465 VDD2.n125 VDD2.n98 12.0247
R3466 VDD2.n43 VDD2.n16 12.0247
R3467 VDD2.n54 VDD2.n53 12.0247
R3468 VDD2.n138 VDD2.n91 11.249
R3469 VDD2.n122 VDD2.n121 11.249
R3470 VDD2.n40 VDD2.n39 11.249
R3471 VDD2.n57 VDD2.n10 11.249
R3472 VDD2.n139 VDD2.n89 10.4732
R3473 VDD2.n118 VDD2.n100 10.4732
R3474 VDD2.n36 VDD2.n18 10.4732
R3475 VDD2.n58 VDD2.n8 10.4732
R3476 VDD2.n107 VDD2.n106 10.2747
R3477 VDD2.n25 VDD2.n24 10.2747
R3478 VDD2.n143 VDD2.n142 9.69747
R3479 VDD2.n117 VDD2.n102 9.69747
R3480 VDD2.n35 VDD2.n20 9.69747
R3481 VDD2.n62 VDD2.n61 9.69747
R3482 VDD2.n157 VDD2.n156 9.45567
R3483 VDD2.n76 VDD2.n75 9.45567
R3484 VDD2.n109 VDD2.n108 9.3005
R3485 VDD2.n104 VDD2.n103 9.3005
R3486 VDD2.n115 VDD2.n114 9.3005
R3487 VDD2.n117 VDD2.n116 9.3005
R3488 VDD2.n100 VDD2.n99 9.3005
R3489 VDD2.n123 VDD2.n122 9.3005
R3490 VDD2.n125 VDD2.n124 9.3005
R3491 VDD2.n97 VDD2.n94 9.3005
R3492 VDD2.n156 VDD2.n155 9.3005
R3493 VDD2.n83 VDD2.n82 9.3005
R3494 VDD2.n150 VDD2.n149 9.3005
R3495 VDD2.n148 VDD2.n147 9.3005
R3496 VDD2.n87 VDD2.n86 9.3005
R3497 VDD2.n142 VDD2.n141 9.3005
R3498 VDD2.n140 VDD2.n139 9.3005
R3499 VDD2.n91 VDD2.n90 9.3005
R3500 VDD2.n134 VDD2.n133 9.3005
R3501 VDD2.n132 VDD2.n131 9.3005
R3502 VDD2.n2 VDD2.n1 9.3005
R3503 VDD2.n75 VDD2.n74 9.3005
R3504 VDD2.n67 VDD2.n66 9.3005
R3505 VDD2.n6 VDD2.n5 9.3005
R3506 VDD2.n61 VDD2.n60 9.3005
R3507 VDD2.n59 VDD2.n58 9.3005
R3508 VDD2.n10 VDD2.n9 9.3005
R3509 VDD2.n53 VDD2.n52 9.3005
R3510 VDD2.n51 VDD2.n50 9.3005
R3511 VDD2.n27 VDD2.n26 9.3005
R3512 VDD2.n22 VDD2.n21 9.3005
R3513 VDD2.n33 VDD2.n32 9.3005
R3514 VDD2.n35 VDD2.n34 9.3005
R3515 VDD2.n18 VDD2.n17 9.3005
R3516 VDD2.n41 VDD2.n40 9.3005
R3517 VDD2.n43 VDD2.n42 9.3005
R3518 VDD2.n44 VDD2.n13 9.3005
R3519 VDD2.n69 VDD2.n68 9.3005
R3520 VDD2.n146 VDD2.n87 8.92171
R3521 VDD2.n114 VDD2.n113 8.92171
R3522 VDD2.n32 VDD2.n31 8.92171
R3523 VDD2.n65 VDD2.n6 8.92171
R3524 VDD2.n157 VDD2.n81 8.14595
R3525 VDD2.n147 VDD2.n85 8.14595
R3526 VDD2.n110 VDD2.n104 8.14595
R3527 VDD2.n28 VDD2.n22 8.14595
R3528 VDD2.n66 VDD2.n4 8.14595
R3529 VDD2.n76 VDD2.n0 8.14595
R3530 VDD2.n155 VDD2.n154 7.3702
R3531 VDD2.n151 VDD2.n150 7.3702
R3532 VDD2.n109 VDD2.n106 7.3702
R3533 VDD2.n27 VDD2.n24 7.3702
R3534 VDD2.n70 VDD2.n69 7.3702
R3535 VDD2.n74 VDD2.n73 7.3702
R3536 VDD2.n154 VDD2.n83 6.59444
R3537 VDD2.n151 VDD2.n83 6.59444
R3538 VDD2.n70 VDD2.n2 6.59444
R3539 VDD2.n73 VDD2.n2 6.59444
R3540 VDD2.n155 VDD2.n81 5.81868
R3541 VDD2.n150 VDD2.n85 5.81868
R3542 VDD2.n110 VDD2.n109 5.81868
R3543 VDD2.n28 VDD2.n27 5.81868
R3544 VDD2.n69 VDD2.n4 5.81868
R3545 VDD2.n74 VDD2.n0 5.81868
R3546 VDD2.n147 VDD2.n146 5.04292
R3547 VDD2.n113 VDD2.n104 5.04292
R3548 VDD2.n31 VDD2.n22 5.04292
R3549 VDD2.n66 VDD2.n65 5.04292
R3550 VDD2.n143 VDD2.n87 4.26717
R3551 VDD2.n114 VDD2.n102 4.26717
R3552 VDD2.n32 VDD2.n20 4.26717
R3553 VDD2.n62 VDD2.n6 4.26717
R3554 VDD2.n142 VDD2.n89 3.49141
R3555 VDD2.n118 VDD2.n117 3.49141
R3556 VDD2.n36 VDD2.n35 3.49141
R3557 VDD2.n61 VDD2.n8 3.49141
R3558 VDD2.n160 VDD2.n158 3.34533
R3559 VDD2.n108 VDD2.n107 2.84303
R3560 VDD2.n26 VDD2.n25 2.84303
R3561 VDD2.n139 VDD2.n138 2.71565
R3562 VDD2.n121 VDD2.n100 2.71565
R3563 VDD2.n39 VDD2.n18 2.71565
R3564 VDD2.n58 VDD2.n57 2.71565
R3565 VDD2.n135 VDD2.n91 1.93989
R3566 VDD2.n122 VDD2.n98 1.93989
R3567 VDD2.n40 VDD2.n16 1.93989
R3568 VDD2.n54 VDD2.n10 1.93989
R3569 VDD2.n161 VDD2.t9 1.39487
R3570 VDD2.n161 VDD2.t3 1.39487
R3571 VDD2.n159 VDD2.t5 1.39487
R3572 VDD2.n159 VDD2.t8 1.39487
R3573 VDD2.n79 VDD2.t6 1.39487
R3574 VDD2.n79 VDD2.t7 1.39487
R3575 VDD2.n77 VDD2.t0 1.39487
R3576 VDD2.n77 VDD2.t1 1.39487
R3577 VDD2.n134 VDD2.n93 1.16414
R3578 VDD2.n126 VDD2.n125 1.16414
R3579 VDD2.n45 VDD2.n43 1.16414
R3580 VDD2.n53 VDD2.n12 1.16414
R3581 VDD2 VDD2.n160 0.894897
R3582 VDD2.n80 VDD2.n78 0.781361
R3583 VDD2.n131 VDD2.n130 0.388379
R3584 VDD2.n97 VDD2.n95 0.388379
R3585 VDD2.n44 VDD2.n14 0.388379
R3586 VDD2.n50 VDD2.n49 0.388379
R3587 VDD2.n156 VDD2.n82 0.155672
R3588 VDD2.n149 VDD2.n82 0.155672
R3589 VDD2.n149 VDD2.n148 0.155672
R3590 VDD2.n148 VDD2.n86 0.155672
R3591 VDD2.n141 VDD2.n86 0.155672
R3592 VDD2.n141 VDD2.n140 0.155672
R3593 VDD2.n140 VDD2.n90 0.155672
R3594 VDD2.n133 VDD2.n90 0.155672
R3595 VDD2.n133 VDD2.n132 0.155672
R3596 VDD2.n132 VDD2.n94 0.155672
R3597 VDD2.n124 VDD2.n94 0.155672
R3598 VDD2.n124 VDD2.n123 0.155672
R3599 VDD2.n123 VDD2.n99 0.155672
R3600 VDD2.n116 VDD2.n99 0.155672
R3601 VDD2.n116 VDD2.n115 0.155672
R3602 VDD2.n115 VDD2.n103 0.155672
R3603 VDD2.n108 VDD2.n103 0.155672
R3604 VDD2.n26 VDD2.n21 0.155672
R3605 VDD2.n33 VDD2.n21 0.155672
R3606 VDD2.n34 VDD2.n33 0.155672
R3607 VDD2.n34 VDD2.n17 0.155672
R3608 VDD2.n41 VDD2.n17 0.155672
R3609 VDD2.n42 VDD2.n41 0.155672
R3610 VDD2.n42 VDD2.n13 0.155672
R3611 VDD2.n51 VDD2.n13 0.155672
R3612 VDD2.n52 VDD2.n51 0.155672
R3613 VDD2.n52 VDD2.n9 0.155672
R3614 VDD2.n59 VDD2.n9 0.155672
R3615 VDD2.n60 VDD2.n59 0.155672
R3616 VDD2.n60 VDD2.n5 0.155672
R3617 VDD2.n67 VDD2.n5 0.155672
R3618 VDD2.n68 VDD2.n67 0.155672
R3619 VDD2.n68 VDD2.n1 0.155672
R3620 VDD2.n75 VDD2.n1 0.155672
C0 VN VDD1 0.155846f
C1 VN VTAIL 14.172501f
C2 VTAIL VDD1 11.712701f
C3 VN VDD2 13.226901f
C4 VDD1 VDD2 2.79333f
C5 VTAIL VDD2 11.7705f
C6 VN VP 10.1962f
C7 VDD1 VP 13.772099f
C8 VTAIL VP 14.1867f
C9 VDD2 VP 0.705246f
C10 VDD2 B 8.696749f
C11 VDD1 B 8.672803f
C12 VTAIL B 9.818188f
C13 VN B 22.82462f
C14 VP B 21.389992f
C15 VDD2.n0 B 0.034788f
C16 VDD2.n1 B 0.024284f
C17 VDD2.n2 B 0.013049f
C18 VDD2.n3 B 0.030843f
C19 VDD2.n4 B 0.013816f
C20 VDD2.n5 B 0.024284f
C21 VDD2.n6 B 0.013049f
C22 VDD2.n7 B 0.030843f
C23 VDD2.n8 B 0.013816f
C24 VDD2.n9 B 0.024284f
C25 VDD2.n10 B 0.013049f
C26 VDD2.n11 B 0.030843f
C27 VDD2.n12 B 0.013816f
C28 VDD2.n13 B 0.024284f
C29 VDD2.n14 B 0.013433f
C30 VDD2.n15 B 0.030843f
C31 VDD2.n16 B 0.013816f
C32 VDD2.n17 B 0.024284f
C33 VDD2.n18 B 0.013049f
C34 VDD2.n19 B 0.030843f
C35 VDD2.n20 B 0.013816f
C36 VDD2.n21 B 0.024284f
C37 VDD2.n22 B 0.013049f
C38 VDD2.n23 B 0.023132f
C39 VDD2.n24 B 0.021804f
C40 VDD2.t4 B 0.052379f
C41 VDD2.n25 B 0.195591f
C42 VDD2.n26 B 1.46268f
C43 VDD2.n27 B 0.013049f
C44 VDD2.n28 B 0.013816f
C45 VDD2.n29 B 0.030843f
C46 VDD2.n30 B 0.030843f
C47 VDD2.n31 B 0.013816f
C48 VDD2.n32 B 0.013049f
C49 VDD2.n33 B 0.024284f
C50 VDD2.n34 B 0.024284f
C51 VDD2.n35 B 0.013049f
C52 VDD2.n36 B 0.013816f
C53 VDD2.n37 B 0.030843f
C54 VDD2.n38 B 0.030843f
C55 VDD2.n39 B 0.013816f
C56 VDD2.n40 B 0.013049f
C57 VDD2.n41 B 0.024284f
C58 VDD2.n42 B 0.024284f
C59 VDD2.n43 B 0.013049f
C60 VDD2.n44 B 0.013049f
C61 VDD2.n45 B 0.013816f
C62 VDD2.n46 B 0.030843f
C63 VDD2.n47 B 0.030843f
C64 VDD2.n48 B 0.030843f
C65 VDD2.n49 B 0.013433f
C66 VDD2.n50 B 0.013049f
C67 VDD2.n51 B 0.024284f
C68 VDD2.n52 B 0.024284f
C69 VDD2.n53 B 0.013049f
C70 VDD2.n54 B 0.013816f
C71 VDD2.n55 B 0.030843f
C72 VDD2.n56 B 0.030843f
C73 VDD2.n57 B 0.013816f
C74 VDD2.n58 B 0.013049f
C75 VDD2.n59 B 0.024284f
C76 VDD2.n60 B 0.024284f
C77 VDD2.n61 B 0.013049f
C78 VDD2.n62 B 0.013816f
C79 VDD2.n63 B 0.030843f
C80 VDD2.n64 B 0.030843f
C81 VDD2.n65 B 0.013816f
C82 VDD2.n66 B 0.013049f
C83 VDD2.n67 B 0.024284f
C84 VDD2.n68 B 0.024284f
C85 VDD2.n69 B 0.013049f
C86 VDD2.n70 B 0.013816f
C87 VDD2.n71 B 0.030843f
C88 VDD2.n72 B 0.067928f
C89 VDD2.n73 B 0.013816f
C90 VDD2.n74 B 0.013049f
C91 VDD2.n75 B 0.053476f
C92 VDD2.n76 B 0.075102f
C93 VDD2.t0 B 0.272491f
C94 VDD2.t1 B 0.272491f
C95 VDD2.n77 B 2.4488f
C96 VDD2.n78 B 0.816019f
C97 VDD2.t6 B 0.272491f
C98 VDD2.t7 B 0.272491f
C99 VDD2.n79 B 2.47516f
C100 VDD2.n80 B 3.44055f
C101 VDD2.n81 B 0.034788f
C102 VDD2.n82 B 0.024284f
C103 VDD2.n83 B 0.013049f
C104 VDD2.n84 B 0.030843f
C105 VDD2.n85 B 0.013816f
C106 VDD2.n86 B 0.024284f
C107 VDD2.n87 B 0.013049f
C108 VDD2.n88 B 0.030843f
C109 VDD2.n89 B 0.013816f
C110 VDD2.n90 B 0.024284f
C111 VDD2.n91 B 0.013049f
C112 VDD2.n92 B 0.030843f
C113 VDD2.n93 B 0.013816f
C114 VDD2.n94 B 0.024284f
C115 VDD2.n95 B 0.013433f
C116 VDD2.n96 B 0.030843f
C117 VDD2.n97 B 0.013049f
C118 VDD2.n98 B 0.013816f
C119 VDD2.n99 B 0.024284f
C120 VDD2.n100 B 0.013049f
C121 VDD2.n101 B 0.030843f
C122 VDD2.n102 B 0.013816f
C123 VDD2.n103 B 0.024284f
C124 VDD2.n104 B 0.013049f
C125 VDD2.n105 B 0.023132f
C126 VDD2.n106 B 0.021804f
C127 VDD2.t2 B 0.052379f
C128 VDD2.n107 B 0.195591f
C129 VDD2.n108 B 1.46268f
C130 VDD2.n109 B 0.013049f
C131 VDD2.n110 B 0.013816f
C132 VDD2.n111 B 0.030843f
C133 VDD2.n112 B 0.030843f
C134 VDD2.n113 B 0.013816f
C135 VDD2.n114 B 0.013049f
C136 VDD2.n115 B 0.024284f
C137 VDD2.n116 B 0.024284f
C138 VDD2.n117 B 0.013049f
C139 VDD2.n118 B 0.013816f
C140 VDD2.n119 B 0.030843f
C141 VDD2.n120 B 0.030843f
C142 VDD2.n121 B 0.013816f
C143 VDD2.n122 B 0.013049f
C144 VDD2.n123 B 0.024284f
C145 VDD2.n124 B 0.024284f
C146 VDD2.n125 B 0.013049f
C147 VDD2.n126 B 0.013816f
C148 VDD2.n127 B 0.030843f
C149 VDD2.n128 B 0.030843f
C150 VDD2.n129 B 0.030843f
C151 VDD2.n130 B 0.013433f
C152 VDD2.n131 B 0.013049f
C153 VDD2.n132 B 0.024284f
C154 VDD2.n133 B 0.024284f
C155 VDD2.n134 B 0.013049f
C156 VDD2.n135 B 0.013816f
C157 VDD2.n136 B 0.030843f
C158 VDD2.n137 B 0.030843f
C159 VDD2.n138 B 0.013816f
C160 VDD2.n139 B 0.013049f
C161 VDD2.n140 B 0.024284f
C162 VDD2.n141 B 0.024284f
C163 VDD2.n142 B 0.013049f
C164 VDD2.n143 B 0.013816f
C165 VDD2.n144 B 0.030843f
C166 VDD2.n145 B 0.030843f
C167 VDD2.n146 B 0.013816f
C168 VDD2.n147 B 0.013049f
C169 VDD2.n148 B 0.024284f
C170 VDD2.n149 B 0.024284f
C171 VDD2.n150 B 0.013049f
C172 VDD2.n151 B 0.013816f
C173 VDD2.n152 B 0.030843f
C174 VDD2.n153 B 0.067928f
C175 VDD2.n154 B 0.013816f
C176 VDD2.n155 B 0.013049f
C177 VDD2.n156 B 0.053476f
C178 VDD2.n157 B 0.054834f
C179 VDD2.n158 B 3.32886f
C180 VDD2.t5 B 0.272491f
C181 VDD2.t8 B 0.272491f
C182 VDD2.n159 B 2.44881f
C183 VDD2.n160 B 0.537485f
C184 VDD2.t9 B 0.272491f
C185 VDD2.t3 B 0.272491f
C186 VDD2.n161 B 2.47511f
C187 VN.t2 B 2.3573f
C188 VN.n0 B 0.889508f
C189 VN.n1 B 0.017087f
C190 VN.n2 B 0.02153f
C191 VN.n3 B 0.017087f
C192 VN.n4 B 0.019798f
C193 VN.n5 B 0.017087f
C194 VN.n6 B 0.014601f
C195 VN.n7 B 0.017087f
C196 VN.t8 B 2.3573f
C197 VN.n8 B 0.836341f
C198 VN.n9 B 0.017087f
C199 VN.n10 B 0.014601f
C200 VN.n11 B 0.017087f
C201 VN.t9 B 2.3573f
C202 VN.n12 B 0.883549f
C203 VN.t5 B 2.60419f
C204 VN.n13 B 0.835312f
C205 VN.n14 B 0.211052f
C206 VN.n15 B 0.027933f
C207 VN.n16 B 0.031687f
C208 VN.n17 B 0.034342f
C209 VN.n18 B 0.017087f
C210 VN.n19 B 0.017087f
C211 VN.n20 B 0.017087f
C212 VN.n21 B 0.032422f
C213 VN.n22 B 0.031687f
C214 VN.n23 B 0.031687f
C215 VN.n24 B 0.017087f
C216 VN.n25 B 0.017087f
C217 VN.n26 B 0.017087f
C218 VN.n27 B 0.031687f
C219 VN.n28 B 0.031687f
C220 VN.n29 B 0.032422f
C221 VN.n30 B 0.017087f
C222 VN.n31 B 0.017087f
C223 VN.n32 B 0.017087f
C224 VN.n33 B 0.034342f
C225 VN.n34 B 0.031687f
C226 VN.t3 B 2.3573f
C227 VN.n35 B 0.820298f
C228 VN.n36 B 0.027933f
C229 VN.n37 B 0.017087f
C230 VN.n38 B 0.017087f
C231 VN.n39 B 0.017087f
C232 VN.n40 B 0.031687f
C233 VN.n41 B 0.031687f
C234 VN.n42 B 0.028148f
C235 VN.n43 B 0.017087f
C236 VN.n44 B 0.017087f
C237 VN.n45 B 0.017087f
C238 VN.n46 B 0.031687f
C239 VN.n47 B 0.031687f
C240 VN.n48 B 0.024178f
C241 VN.n49 B 0.027574f
C242 VN.n50 B 0.044465f
C243 VN.t7 B 2.3573f
C244 VN.n51 B 0.889508f
C245 VN.n52 B 0.017087f
C246 VN.n53 B 0.02153f
C247 VN.n54 B 0.017087f
C248 VN.n55 B 0.019798f
C249 VN.n56 B 0.017087f
C250 VN.t4 B 2.3573f
C251 VN.n57 B 0.820298f
C252 VN.n58 B 0.014601f
C253 VN.n59 B 0.017087f
C254 VN.t1 B 2.3573f
C255 VN.n60 B 0.836341f
C256 VN.n61 B 0.017087f
C257 VN.n62 B 0.014601f
C258 VN.n63 B 0.017087f
C259 VN.t0 B 2.3573f
C260 VN.n64 B 0.883549f
C261 VN.t6 B 2.60419f
C262 VN.n65 B 0.835312f
C263 VN.n66 B 0.211052f
C264 VN.n67 B 0.027933f
C265 VN.n68 B 0.031687f
C266 VN.n69 B 0.034342f
C267 VN.n70 B 0.017087f
C268 VN.n71 B 0.017087f
C269 VN.n72 B 0.017087f
C270 VN.n73 B 0.032422f
C271 VN.n74 B 0.031687f
C272 VN.n75 B 0.031687f
C273 VN.n76 B 0.017087f
C274 VN.n77 B 0.017087f
C275 VN.n78 B 0.017087f
C276 VN.n79 B 0.031687f
C277 VN.n80 B 0.031687f
C278 VN.n81 B 0.032422f
C279 VN.n82 B 0.017087f
C280 VN.n83 B 0.017087f
C281 VN.n84 B 0.017087f
C282 VN.n85 B 0.034342f
C283 VN.n86 B 0.031687f
C284 VN.n87 B 0.027933f
C285 VN.n88 B 0.017087f
C286 VN.n89 B 0.017087f
C287 VN.n90 B 0.017087f
C288 VN.n91 B 0.031687f
C289 VN.n92 B 0.031687f
C290 VN.n93 B 0.028148f
C291 VN.n94 B 0.017087f
C292 VN.n95 B 0.017087f
C293 VN.n96 B 0.017087f
C294 VN.n97 B 0.031687f
C295 VN.n98 B 0.031687f
C296 VN.n99 B 0.024178f
C297 VN.n100 B 0.027574f
C298 VN.n101 B 1.26447f
C299 VDD1.n0 B 0.0353f
C300 VDD1.n1 B 0.024641f
C301 VDD1.n2 B 0.013241f
C302 VDD1.n3 B 0.031297f
C303 VDD1.n4 B 0.01402f
C304 VDD1.n5 B 0.024641f
C305 VDD1.n6 B 0.013241f
C306 VDD1.n7 B 0.031297f
C307 VDD1.n8 B 0.01402f
C308 VDD1.n9 B 0.024641f
C309 VDD1.n10 B 0.013241f
C310 VDD1.n11 B 0.031297f
C311 VDD1.n12 B 0.01402f
C312 VDD1.n13 B 0.024641f
C313 VDD1.n14 B 0.01363f
C314 VDD1.n15 B 0.031297f
C315 VDD1.n16 B 0.013241f
C316 VDD1.n17 B 0.01402f
C317 VDD1.n18 B 0.024641f
C318 VDD1.n19 B 0.013241f
C319 VDD1.n20 B 0.031297f
C320 VDD1.n21 B 0.01402f
C321 VDD1.n22 B 0.024641f
C322 VDD1.n23 B 0.013241f
C323 VDD1.n24 B 0.023472f
C324 VDD1.n25 B 0.022124f
C325 VDD1.t8 B 0.05315f
C326 VDD1.n26 B 0.198469f
C327 VDD1.n27 B 1.4842f
C328 VDD1.n28 B 0.013241f
C329 VDD1.n29 B 0.01402f
C330 VDD1.n30 B 0.031297f
C331 VDD1.n31 B 0.031297f
C332 VDD1.n32 B 0.01402f
C333 VDD1.n33 B 0.013241f
C334 VDD1.n34 B 0.024641f
C335 VDD1.n35 B 0.024641f
C336 VDD1.n36 B 0.013241f
C337 VDD1.n37 B 0.01402f
C338 VDD1.n38 B 0.031297f
C339 VDD1.n39 B 0.031297f
C340 VDD1.n40 B 0.01402f
C341 VDD1.n41 B 0.013241f
C342 VDD1.n42 B 0.024641f
C343 VDD1.n43 B 0.024641f
C344 VDD1.n44 B 0.013241f
C345 VDD1.n45 B 0.01402f
C346 VDD1.n46 B 0.031297f
C347 VDD1.n47 B 0.031297f
C348 VDD1.n48 B 0.031297f
C349 VDD1.n49 B 0.01363f
C350 VDD1.n50 B 0.013241f
C351 VDD1.n51 B 0.024641f
C352 VDD1.n52 B 0.024641f
C353 VDD1.n53 B 0.013241f
C354 VDD1.n54 B 0.01402f
C355 VDD1.n55 B 0.031297f
C356 VDD1.n56 B 0.031297f
C357 VDD1.n57 B 0.01402f
C358 VDD1.n58 B 0.013241f
C359 VDD1.n59 B 0.024641f
C360 VDD1.n60 B 0.024641f
C361 VDD1.n61 B 0.013241f
C362 VDD1.n62 B 0.01402f
C363 VDD1.n63 B 0.031297f
C364 VDD1.n64 B 0.031297f
C365 VDD1.n65 B 0.01402f
C366 VDD1.n66 B 0.013241f
C367 VDD1.n67 B 0.024641f
C368 VDD1.n68 B 0.024641f
C369 VDD1.n69 B 0.013241f
C370 VDD1.n70 B 0.01402f
C371 VDD1.n71 B 0.031297f
C372 VDD1.n72 B 0.068928f
C373 VDD1.n73 B 0.01402f
C374 VDD1.n74 B 0.013241f
C375 VDD1.n75 B 0.054263f
C376 VDD1.n76 B 0.076207f
C377 VDD1.t5 B 0.2765f
C378 VDD1.t3 B 0.2765f
C379 VDD1.n77 B 2.48483f
C380 VDD1.n78 B 0.836305f
C381 VDD1.n79 B 0.0353f
C382 VDD1.n80 B 0.024641f
C383 VDD1.n81 B 0.013241f
C384 VDD1.n82 B 0.031297f
C385 VDD1.n83 B 0.01402f
C386 VDD1.n84 B 0.024641f
C387 VDD1.n85 B 0.013241f
C388 VDD1.n86 B 0.031297f
C389 VDD1.n87 B 0.01402f
C390 VDD1.n88 B 0.024641f
C391 VDD1.n89 B 0.013241f
C392 VDD1.n90 B 0.031297f
C393 VDD1.n91 B 0.01402f
C394 VDD1.n92 B 0.024641f
C395 VDD1.n93 B 0.01363f
C396 VDD1.n94 B 0.031297f
C397 VDD1.n95 B 0.01402f
C398 VDD1.n96 B 0.024641f
C399 VDD1.n97 B 0.013241f
C400 VDD1.n98 B 0.031297f
C401 VDD1.n99 B 0.01402f
C402 VDD1.n100 B 0.024641f
C403 VDD1.n101 B 0.013241f
C404 VDD1.n102 B 0.023472f
C405 VDD1.n103 B 0.022124f
C406 VDD1.t1 B 0.05315f
C407 VDD1.n104 B 0.198469f
C408 VDD1.n105 B 1.4842f
C409 VDD1.n106 B 0.013241f
C410 VDD1.n107 B 0.01402f
C411 VDD1.n108 B 0.031297f
C412 VDD1.n109 B 0.031297f
C413 VDD1.n110 B 0.01402f
C414 VDD1.n111 B 0.013241f
C415 VDD1.n112 B 0.024641f
C416 VDD1.n113 B 0.024641f
C417 VDD1.n114 B 0.013241f
C418 VDD1.n115 B 0.01402f
C419 VDD1.n116 B 0.031297f
C420 VDD1.n117 B 0.031297f
C421 VDD1.n118 B 0.01402f
C422 VDD1.n119 B 0.013241f
C423 VDD1.n120 B 0.024641f
C424 VDD1.n121 B 0.024641f
C425 VDD1.n122 B 0.013241f
C426 VDD1.n123 B 0.013241f
C427 VDD1.n124 B 0.01402f
C428 VDD1.n125 B 0.031297f
C429 VDD1.n126 B 0.031297f
C430 VDD1.n127 B 0.031297f
C431 VDD1.n128 B 0.01363f
C432 VDD1.n129 B 0.013241f
C433 VDD1.n130 B 0.024641f
C434 VDD1.n131 B 0.024641f
C435 VDD1.n132 B 0.013241f
C436 VDD1.n133 B 0.01402f
C437 VDD1.n134 B 0.031297f
C438 VDD1.n135 B 0.031297f
C439 VDD1.n136 B 0.01402f
C440 VDD1.n137 B 0.013241f
C441 VDD1.n138 B 0.024641f
C442 VDD1.n139 B 0.024641f
C443 VDD1.n140 B 0.013241f
C444 VDD1.n141 B 0.01402f
C445 VDD1.n142 B 0.031297f
C446 VDD1.n143 B 0.031297f
C447 VDD1.n144 B 0.01402f
C448 VDD1.n145 B 0.013241f
C449 VDD1.n146 B 0.024641f
C450 VDD1.n147 B 0.024641f
C451 VDD1.n148 B 0.013241f
C452 VDD1.n149 B 0.01402f
C453 VDD1.n150 B 0.031297f
C454 VDD1.n151 B 0.068928f
C455 VDD1.n152 B 0.01402f
C456 VDD1.n153 B 0.013241f
C457 VDD1.n154 B 0.054263f
C458 VDD1.n155 B 0.076207f
C459 VDD1.t2 B 0.2765f
C460 VDD1.t0 B 0.2765f
C461 VDD1.n156 B 2.48483f
C462 VDD1.n157 B 0.828024f
C463 VDD1.t6 B 0.2765f
C464 VDD1.t7 B 0.2765f
C465 VDD1.n158 B 2.51157f
C466 VDD1.n159 B 3.64178f
C467 VDD1.t4 B 0.2765f
C468 VDD1.t9 B 0.2765f
C469 VDD1.n160 B 2.48483f
C470 VDD1.n161 B 3.68561f
C471 VTAIL.t2 B 0.280764f
C472 VTAIL.t5 B 0.280764f
C473 VTAIL.n0 B 2.44313f
C474 VTAIL.n1 B 0.637703f
C475 VTAIL.n2 B 0.035844f
C476 VTAIL.n3 B 0.025021f
C477 VTAIL.n4 B 0.013445f
C478 VTAIL.n5 B 0.031779f
C479 VTAIL.n6 B 0.014236f
C480 VTAIL.n7 B 0.025021f
C481 VTAIL.n8 B 0.013445f
C482 VTAIL.n9 B 0.031779f
C483 VTAIL.n10 B 0.014236f
C484 VTAIL.n11 B 0.025021f
C485 VTAIL.n12 B 0.013445f
C486 VTAIL.n13 B 0.031779f
C487 VTAIL.n14 B 0.014236f
C488 VTAIL.n15 B 0.025021f
C489 VTAIL.n16 B 0.013841f
C490 VTAIL.n17 B 0.031779f
C491 VTAIL.n18 B 0.014236f
C492 VTAIL.n19 B 0.025021f
C493 VTAIL.n20 B 0.013445f
C494 VTAIL.n21 B 0.031779f
C495 VTAIL.n22 B 0.014236f
C496 VTAIL.n23 B 0.025021f
C497 VTAIL.n24 B 0.013445f
C498 VTAIL.n25 B 0.023834f
C499 VTAIL.n26 B 0.022465f
C500 VTAIL.t19 B 0.053969f
C501 VTAIL.n27 B 0.201529f
C502 VTAIL.n28 B 1.50709f
C503 VTAIL.n29 B 0.013445f
C504 VTAIL.n30 B 0.014236f
C505 VTAIL.n31 B 0.031779f
C506 VTAIL.n32 B 0.031779f
C507 VTAIL.n33 B 0.014236f
C508 VTAIL.n34 B 0.013445f
C509 VTAIL.n35 B 0.025021f
C510 VTAIL.n36 B 0.025021f
C511 VTAIL.n37 B 0.013445f
C512 VTAIL.n38 B 0.014236f
C513 VTAIL.n39 B 0.031779f
C514 VTAIL.n40 B 0.031779f
C515 VTAIL.n41 B 0.014236f
C516 VTAIL.n42 B 0.013445f
C517 VTAIL.n43 B 0.025021f
C518 VTAIL.n44 B 0.025021f
C519 VTAIL.n45 B 0.013445f
C520 VTAIL.n46 B 0.013445f
C521 VTAIL.n47 B 0.014236f
C522 VTAIL.n48 B 0.031779f
C523 VTAIL.n49 B 0.031779f
C524 VTAIL.n50 B 0.031779f
C525 VTAIL.n51 B 0.013841f
C526 VTAIL.n52 B 0.013445f
C527 VTAIL.n53 B 0.025021f
C528 VTAIL.n54 B 0.025021f
C529 VTAIL.n55 B 0.013445f
C530 VTAIL.n56 B 0.014236f
C531 VTAIL.n57 B 0.031779f
C532 VTAIL.n58 B 0.031779f
C533 VTAIL.n59 B 0.014236f
C534 VTAIL.n60 B 0.013445f
C535 VTAIL.n61 B 0.025021f
C536 VTAIL.n62 B 0.025021f
C537 VTAIL.n63 B 0.013445f
C538 VTAIL.n64 B 0.014236f
C539 VTAIL.n65 B 0.031779f
C540 VTAIL.n66 B 0.031779f
C541 VTAIL.n67 B 0.014236f
C542 VTAIL.n68 B 0.013445f
C543 VTAIL.n69 B 0.025021f
C544 VTAIL.n70 B 0.025021f
C545 VTAIL.n71 B 0.013445f
C546 VTAIL.n72 B 0.014236f
C547 VTAIL.n73 B 0.031779f
C548 VTAIL.n74 B 0.069991f
C549 VTAIL.n75 B 0.014236f
C550 VTAIL.n76 B 0.013445f
C551 VTAIL.n77 B 0.0551f
C552 VTAIL.n78 B 0.039199f
C553 VTAIL.n79 B 0.462209f
C554 VTAIL.t14 B 0.280764f
C555 VTAIL.t18 B 0.280764f
C556 VTAIL.n80 B 2.44313f
C557 VTAIL.n81 B 0.797385f
C558 VTAIL.t16 B 0.280764f
C559 VTAIL.t15 B 0.280764f
C560 VTAIL.n82 B 2.44313f
C561 VTAIL.n83 B 2.39386f
C562 VTAIL.t8 B 0.280764f
C563 VTAIL.t4 B 0.280764f
C564 VTAIL.n84 B 2.44313f
C565 VTAIL.n85 B 2.39386f
C566 VTAIL.t3 B 0.280764f
C567 VTAIL.t1 B 0.280764f
C568 VTAIL.n86 B 2.44313f
C569 VTAIL.n87 B 0.79738f
C570 VTAIL.n88 B 0.035844f
C571 VTAIL.n89 B 0.025021f
C572 VTAIL.n90 B 0.013445f
C573 VTAIL.n91 B 0.031779f
C574 VTAIL.n92 B 0.014236f
C575 VTAIL.n93 B 0.025021f
C576 VTAIL.n94 B 0.013445f
C577 VTAIL.n95 B 0.031779f
C578 VTAIL.n96 B 0.014236f
C579 VTAIL.n97 B 0.025021f
C580 VTAIL.n98 B 0.013445f
C581 VTAIL.n99 B 0.031779f
C582 VTAIL.n100 B 0.014236f
C583 VTAIL.n101 B 0.025021f
C584 VTAIL.n102 B 0.013841f
C585 VTAIL.n103 B 0.031779f
C586 VTAIL.n104 B 0.013445f
C587 VTAIL.n105 B 0.014236f
C588 VTAIL.n106 B 0.025021f
C589 VTAIL.n107 B 0.013445f
C590 VTAIL.n108 B 0.031779f
C591 VTAIL.n109 B 0.014236f
C592 VTAIL.n110 B 0.025021f
C593 VTAIL.n111 B 0.013445f
C594 VTAIL.n112 B 0.023834f
C595 VTAIL.n113 B 0.022465f
C596 VTAIL.t6 B 0.053969f
C597 VTAIL.n114 B 0.201529f
C598 VTAIL.n115 B 1.50709f
C599 VTAIL.n116 B 0.013445f
C600 VTAIL.n117 B 0.014236f
C601 VTAIL.n118 B 0.031779f
C602 VTAIL.n119 B 0.031779f
C603 VTAIL.n120 B 0.014236f
C604 VTAIL.n121 B 0.013445f
C605 VTAIL.n122 B 0.025021f
C606 VTAIL.n123 B 0.025021f
C607 VTAIL.n124 B 0.013445f
C608 VTAIL.n125 B 0.014236f
C609 VTAIL.n126 B 0.031779f
C610 VTAIL.n127 B 0.031779f
C611 VTAIL.n128 B 0.014236f
C612 VTAIL.n129 B 0.013445f
C613 VTAIL.n130 B 0.025021f
C614 VTAIL.n131 B 0.025021f
C615 VTAIL.n132 B 0.013445f
C616 VTAIL.n133 B 0.014236f
C617 VTAIL.n134 B 0.031779f
C618 VTAIL.n135 B 0.031779f
C619 VTAIL.n136 B 0.031779f
C620 VTAIL.n137 B 0.013841f
C621 VTAIL.n138 B 0.013445f
C622 VTAIL.n139 B 0.025021f
C623 VTAIL.n140 B 0.025021f
C624 VTAIL.n141 B 0.013445f
C625 VTAIL.n142 B 0.014236f
C626 VTAIL.n143 B 0.031779f
C627 VTAIL.n144 B 0.031779f
C628 VTAIL.n145 B 0.014236f
C629 VTAIL.n146 B 0.013445f
C630 VTAIL.n147 B 0.025021f
C631 VTAIL.n148 B 0.025021f
C632 VTAIL.n149 B 0.013445f
C633 VTAIL.n150 B 0.014236f
C634 VTAIL.n151 B 0.031779f
C635 VTAIL.n152 B 0.031779f
C636 VTAIL.n153 B 0.014236f
C637 VTAIL.n154 B 0.013445f
C638 VTAIL.n155 B 0.025021f
C639 VTAIL.n156 B 0.025021f
C640 VTAIL.n157 B 0.013445f
C641 VTAIL.n158 B 0.014236f
C642 VTAIL.n159 B 0.031779f
C643 VTAIL.n160 B 0.069991f
C644 VTAIL.n161 B 0.014236f
C645 VTAIL.n162 B 0.013445f
C646 VTAIL.n163 B 0.0551f
C647 VTAIL.n164 B 0.039199f
C648 VTAIL.n165 B 0.462209f
C649 VTAIL.t13 B 0.280764f
C650 VTAIL.t11 B 0.280764f
C651 VTAIL.n166 B 2.44313f
C652 VTAIL.n167 B 0.700425f
C653 VTAIL.t10 B 0.280764f
C654 VTAIL.t17 B 0.280764f
C655 VTAIL.n168 B 2.44313f
C656 VTAIL.n169 B 0.79738f
C657 VTAIL.n170 B 0.035844f
C658 VTAIL.n171 B 0.025021f
C659 VTAIL.n172 B 0.013445f
C660 VTAIL.n173 B 0.031779f
C661 VTAIL.n174 B 0.014236f
C662 VTAIL.n175 B 0.025021f
C663 VTAIL.n176 B 0.013445f
C664 VTAIL.n177 B 0.031779f
C665 VTAIL.n178 B 0.014236f
C666 VTAIL.n179 B 0.025021f
C667 VTAIL.n180 B 0.013445f
C668 VTAIL.n181 B 0.031779f
C669 VTAIL.n182 B 0.014236f
C670 VTAIL.n183 B 0.025021f
C671 VTAIL.n184 B 0.013841f
C672 VTAIL.n185 B 0.031779f
C673 VTAIL.n186 B 0.013445f
C674 VTAIL.n187 B 0.014236f
C675 VTAIL.n188 B 0.025021f
C676 VTAIL.n189 B 0.013445f
C677 VTAIL.n190 B 0.031779f
C678 VTAIL.n191 B 0.014236f
C679 VTAIL.n192 B 0.025021f
C680 VTAIL.n193 B 0.013445f
C681 VTAIL.n194 B 0.023834f
C682 VTAIL.n195 B 0.022465f
C683 VTAIL.t12 B 0.053969f
C684 VTAIL.n196 B 0.201529f
C685 VTAIL.n197 B 1.50709f
C686 VTAIL.n198 B 0.013445f
C687 VTAIL.n199 B 0.014236f
C688 VTAIL.n200 B 0.031779f
C689 VTAIL.n201 B 0.031779f
C690 VTAIL.n202 B 0.014236f
C691 VTAIL.n203 B 0.013445f
C692 VTAIL.n204 B 0.025021f
C693 VTAIL.n205 B 0.025021f
C694 VTAIL.n206 B 0.013445f
C695 VTAIL.n207 B 0.014236f
C696 VTAIL.n208 B 0.031779f
C697 VTAIL.n209 B 0.031779f
C698 VTAIL.n210 B 0.014236f
C699 VTAIL.n211 B 0.013445f
C700 VTAIL.n212 B 0.025021f
C701 VTAIL.n213 B 0.025021f
C702 VTAIL.n214 B 0.013445f
C703 VTAIL.n215 B 0.014236f
C704 VTAIL.n216 B 0.031779f
C705 VTAIL.n217 B 0.031779f
C706 VTAIL.n218 B 0.031779f
C707 VTAIL.n219 B 0.013841f
C708 VTAIL.n220 B 0.013445f
C709 VTAIL.n221 B 0.025021f
C710 VTAIL.n222 B 0.025021f
C711 VTAIL.n223 B 0.013445f
C712 VTAIL.n224 B 0.014236f
C713 VTAIL.n225 B 0.031779f
C714 VTAIL.n226 B 0.031779f
C715 VTAIL.n227 B 0.014236f
C716 VTAIL.n228 B 0.013445f
C717 VTAIL.n229 B 0.025021f
C718 VTAIL.n230 B 0.025021f
C719 VTAIL.n231 B 0.013445f
C720 VTAIL.n232 B 0.014236f
C721 VTAIL.n233 B 0.031779f
C722 VTAIL.n234 B 0.031779f
C723 VTAIL.n235 B 0.014236f
C724 VTAIL.n236 B 0.013445f
C725 VTAIL.n237 B 0.025021f
C726 VTAIL.n238 B 0.025021f
C727 VTAIL.n239 B 0.013445f
C728 VTAIL.n240 B 0.014236f
C729 VTAIL.n241 B 0.031779f
C730 VTAIL.n242 B 0.069991f
C731 VTAIL.n243 B 0.014236f
C732 VTAIL.n244 B 0.013445f
C733 VTAIL.n245 B 0.0551f
C734 VTAIL.n246 B 0.039199f
C735 VTAIL.n247 B 1.88597f
C736 VTAIL.n248 B 0.035844f
C737 VTAIL.n249 B 0.025021f
C738 VTAIL.n250 B 0.013445f
C739 VTAIL.n251 B 0.031779f
C740 VTAIL.n252 B 0.014236f
C741 VTAIL.n253 B 0.025021f
C742 VTAIL.n254 B 0.013445f
C743 VTAIL.n255 B 0.031779f
C744 VTAIL.n256 B 0.014236f
C745 VTAIL.n257 B 0.025021f
C746 VTAIL.n258 B 0.013445f
C747 VTAIL.n259 B 0.031779f
C748 VTAIL.n260 B 0.014236f
C749 VTAIL.n261 B 0.025021f
C750 VTAIL.n262 B 0.013841f
C751 VTAIL.n263 B 0.031779f
C752 VTAIL.n264 B 0.014236f
C753 VTAIL.n265 B 0.025021f
C754 VTAIL.n266 B 0.013445f
C755 VTAIL.n267 B 0.031779f
C756 VTAIL.n268 B 0.014236f
C757 VTAIL.n269 B 0.025021f
C758 VTAIL.n270 B 0.013445f
C759 VTAIL.n271 B 0.023834f
C760 VTAIL.n272 B 0.022465f
C761 VTAIL.t0 B 0.053969f
C762 VTAIL.n273 B 0.201529f
C763 VTAIL.n274 B 1.50709f
C764 VTAIL.n275 B 0.013445f
C765 VTAIL.n276 B 0.014236f
C766 VTAIL.n277 B 0.031779f
C767 VTAIL.n278 B 0.031779f
C768 VTAIL.n279 B 0.014236f
C769 VTAIL.n280 B 0.013445f
C770 VTAIL.n281 B 0.025021f
C771 VTAIL.n282 B 0.025021f
C772 VTAIL.n283 B 0.013445f
C773 VTAIL.n284 B 0.014236f
C774 VTAIL.n285 B 0.031779f
C775 VTAIL.n286 B 0.031779f
C776 VTAIL.n287 B 0.014236f
C777 VTAIL.n288 B 0.013445f
C778 VTAIL.n289 B 0.025021f
C779 VTAIL.n290 B 0.025021f
C780 VTAIL.n291 B 0.013445f
C781 VTAIL.n292 B 0.013445f
C782 VTAIL.n293 B 0.014236f
C783 VTAIL.n294 B 0.031779f
C784 VTAIL.n295 B 0.031779f
C785 VTAIL.n296 B 0.031779f
C786 VTAIL.n297 B 0.013841f
C787 VTAIL.n298 B 0.013445f
C788 VTAIL.n299 B 0.025021f
C789 VTAIL.n300 B 0.025021f
C790 VTAIL.n301 B 0.013445f
C791 VTAIL.n302 B 0.014236f
C792 VTAIL.n303 B 0.031779f
C793 VTAIL.n304 B 0.031779f
C794 VTAIL.n305 B 0.014236f
C795 VTAIL.n306 B 0.013445f
C796 VTAIL.n307 B 0.025021f
C797 VTAIL.n308 B 0.025021f
C798 VTAIL.n309 B 0.013445f
C799 VTAIL.n310 B 0.014236f
C800 VTAIL.n311 B 0.031779f
C801 VTAIL.n312 B 0.031779f
C802 VTAIL.n313 B 0.014236f
C803 VTAIL.n314 B 0.013445f
C804 VTAIL.n315 B 0.025021f
C805 VTAIL.n316 B 0.025021f
C806 VTAIL.n317 B 0.013445f
C807 VTAIL.n318 B 0.014236f
C808 VTAIL.n319 B 0.031779f
C809 VTAIL.n320 B 0.069991f
C810 VTAIL.n321 B 0.014236f
C811 VTAIL.n322 B 0.013445f
C812 VTAIL.n323 B 0.0551f
C813 VTAIL.n324 B 0.039199f
C814 VTAIL.n325 B 1.88597f
C815 VTAIL.t9 B 0.280764f
C816 VTAIL.t7 B 0.280764f
C817 VTAIL.n326 B 2.44313f
C818 VTAIL.n327 B 0.590442f
C819 VP.t2 B 2.39645f
C820 VP.n0 B 0.90428f
C821 VP.n1 B 0.017371f
C822 VP.n2 B 0.021887f
C823 VP.n3 B 0.017371f
C824 VP.n4 B 0.020127f
C825 VP.n5 B 0.017371f
C826 VP.n6 B 0.014844f
C827 VP.n7 B 0.017371f
C828 VP.t9 B 2.39645f
C829 VP.n8 B 0.85023f
C830 VP.n9 B 0.017371f
C831 VP.n10 B 0.014844f
C832 VP.n11 B 0.017371f
C833 VP.t7 B 2.39645f
C834 VP.n12 B 0.83392f
C835 VP.n13 B 0.017371f
C836 VP.n14 B 0.028616f
C837 VP.n15 B 0.017371f
C838 VP.n16 B 0.02458f
C839 VP.t0 B 2.39645f
C840 VP.n17 B 0.90428f
C841 VP.n18 B 0.017371f
C842 VP.n19 B 0.021887f
C843 VP.n20 B 0.017371f
C844 VP.n21 B 0.020127f
C845 VP.n22 B 0.017371f
C846 VP.n23 B 0.014844f
C847 VP.n24 B 0.017371f
C848 VP.t6 B 2.39645f
C849 VP.n25 B 0.85023f
C850 VP.n26 B 0.017371f
C851 VP.n27 B 0.014844f
C852 VP.n28 B 0.017371f
C853 VP.t4 B 2.39645f
C854 VP.n29 B 0.898222f
C855 VP.t1 B 2.64744f
C856 VP.n30 B 0.849185f
C857 VP.n31 B 0.214558f
C858 VP.n32 B 0.028396f
C859 VP.n33 B 0.032213f
C860 VP.n34 B 0.034912f
C861 VP.n35 B 0.017371f
C862 VP.n36 B 0.017371f
C863 VP.n37 B 0.017371f
C864 VP.n38 B 0.03296f
C865 VP.n39 B 0.032213f
C866 VP.n40 B 0.032213f
C867 VP.n41 B 0.017371f
C868 VP.n42 B 0.017371f
C869 VP.n43 B 0.017371f
C870 VP.n44 B 0.032213f
C871 VP.n45 B 0.032213f
C872 VP.n46 B 0.03296f
C873 VP.n47 B 0.017371f
C874 VP.n48 B 0.017371f
C875 VP.n49 B 0.017371f
C876 VP.n50 B 0.034912f
C877 VP.n51 B 0.032213f
C878 VP.t5 B 2.39645f
C879 VP.n52 B 0.83392f
C880 VP.n53 B 0.028396f
C881 VP.n54 B 0.017371f
C882 VP.n55 B 0.017371f
C883 VP.n56 B 0.017371f
C884 VP.n57 B 0.032213f
C885 VP.n58 B 0.032213f
C886 VP.n59 B 0.028616f
C887 VP.n60 B 0.017371f
C888 VP.n61 B 0.017371f
C889 VP.n62 B 0.017371f
C890 VP.n63 B 0.032213f
C891 VP.n64 B 0.032213f
C892 VP.n65 B 0.02458f
C893 VP.n66 B 0.028032f
C894 VP.n67 B 1.27878f
C895 VP.t8 B 2.39645f
C896 VP.n68 B 0.90428f
C897 VP.n69 B 1.2892f
C898 VP.n70 B 0.028032f
C899 VP.n71 B 0.017371f
C900 VP.n72 B 0.032213f
C901 VP.n73 B 0.032213f
C902 VP.n74 B 0.021887f
C903 VP.n75 B 0.017371f
C904 VP.n76 B 0.017371f
C905 VP.n77 B 0.017371f
C906 VP.n78 B 0.032213f
C907 VP.n79 B 0.032213f
C908 VP.n80 B 0.020127f
C909 VP.n81 B 0.017371f
C910 VP.n82 B 0.017371f
C911 VP.n83 B 0.028396f
C912 VP.n84 B 0.032213f
C913 VP.n85 B 0.034912f
C914 VP.n86 B 0.017371f
C915 VP.n87 B 0.017371f
C916 VP.n88 B 0.017371f
C917 VP.n89 B 0.03296f
C918 VP.n90 B 0.032213f
C919 VP.n91 B 0.032213f
C920 VP.n92 B 0.017371f
C921 VP.n93 B 0.017371f
C922 VP.n94 B 0.017371f
C923 VP.n95 B 0.032213f
C924 VP.n96 B 0.032213f
C925 VP.n97 B 0.03296f
C926 VP.n98 B 0.017371f
C927 VP.n99 B 0.017371f
C928 VP.n100 B 0.017371f
C929 VP.n101 B 0.034912f
C930 VP.n102 B 0.032213f
C931 VP.t3 B 2.39645f
C932 VP.n103 B 0.83392f
C933 VP.n104 B 0.028396f
C934 VP.n105 B 0.017371f
C935 VP.n106 B 0.017371f
C936 VP.n107 B 0.017371f
C937 VP.n108 B 0.032213f
C938 VP.n109 B 0.032213f
C939 VP.n110 B 0.028616f
C940 VP.n111 B 0.017371f
C941 VP.n112 B 0.017371f
C942 VP.n113 B 0.017371f
C943 VP.n114 B 0.032213f
C944 VP.n115 B 0.032213f
C945 VP.n116 B 0.02458f
C946 VP.n117 B 0.028032f
C947 VP.n118 B 0.045204f
.ends

