* NGSPICE file created from diff_pair_sample_0343.ext - technology: sky130A

.subckt diff_pair_sample_0343 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X1 VTAIL.t1 VN.t0 VDD2.t9 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X2 VDD2.t8 VN.t1 VTAIL.t3 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X3 VTAIL.t6 VN.t2 VDD2.t7 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X4 VTAIL.t18 VP.t1 VDD1.t0 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X5 B.t11 B.t9 B.t10 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=0 ps=0 w=14.32 l=3.18
X6 VDD1.t9 VP.t2 VTAIL.t17 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=5.5848 ps=29.42 w=14.32 l=3.18
X7 B.t8 B.t6 B.t7 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=0 ps=0 w=14.32 l=3.18
X8 VTAIL.t2 VN.t3 VDD2.t6 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X9 VDD1.t8 VP.t3 VTAIL.t16 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=5.5848 ps=29.42 w=14.32 l=3.18
X10 VTAIL.t15 VP.t4 VDD1.t5 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X11 VDD2.t5 VN.t4 VTAIL.t4 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=2.3628 ps=14.65 w=14.32 l=3.18
X12 VDD2.t4 VN.t5 VTAIL.t9 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=2.3628 ps=14.65 w=14.32 l=3.18
X13 VDD1.t4 VP.t5 VTAIL.t14 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X14 VDD2.t3 VN.t6 VTAIL.t0 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=5.5848 ps=29.42 w=14.32 l=3.18
X15 VDD2.t2 VN.t7 VTAIL.t7 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X16 VDD1.t7 VP.t6 VTAIL.t13 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=2.3628 ps=14.65 w=14.32 l=3.18
X17 VTAIL.t8 VN.t8 VDD2.t1 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X18 B.t5 B.t3 B.t4 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=0 ps=0 w=14.32 l=3.18
X19 VDD1.t6 VP.t7 VTAIL.t12 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=2.3628 ps=14.65 w=14.32 l=3.18
X20 B.t2 B.t0 B.t1 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=5.5848 pd=29.42 as=0 ps=0 w=14.32 l=3.18
X21 VDD2.t0 VN.t9 VTAIL.t5 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=5.5848 ps=29.42 w=14.32 l=3.18
X22 VTAIL.t11 VP.t8 VDD1.t3 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
X23 VDD1.t2 VP.t9 VTAIL.t10 w_n5182_n3832# sky130_fd_pr__pfet_01v8 ad=2.3628 pd=14.65 as=2.3628 ps=14.65 w=14.32 l=3.18
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n52 VP.n51 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n20 161.3
R16 VP.n57 VP.n56 161.3
R17 VP.n58 VP.n19 161.3
R18 VP.n60 VP.n59 161.3
R19 VP.n61 VP.n18 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n109 VP.n108 161.3
R22 VP.n107 VP.n1 161.3
R23 VP.n106 VP.n105 161.3
R24 VP.n104 VP.n2 161.3
R25 VP.n103 VP.n102 161.3
R26 VP.n101 VP.n3 161.3
R27 VP.n100 VP.n99 161.3
R28 VP.n98 VP.n97 161.3
R29 VP.n96 VP.n5 161.3
R30 VP.n95 VP.n94 161.3
R31 VP.n93 VP.n6 161.3
R32 VP.n92 VP.n91 161.3
R33 VP.n90 VP.n7 161.3
R34 VP.n89 VP.n88 161.3
R35 VP.n87 VP.n86 161.3
R36 VP.n85 VP.n9 161.3
R37 VP.n84 VP.n83 161.3
R38 VP.n82 VP.n10 161.3
R39 VP.n81 VP.n80 161.3
R40 VP.n79 VP.n11 161.3
R41 VP.n78 VP.n77 161.3
R42 VP.n76 VP.n75 161.3
R43 VP.n74 VP.n13 161.3
R44 VP.n73 VP.n72 161.3
R45 VP.n71 VP.n14 161.3
R46 VP.n70 VP.n69 161.3
R47 VP.n68 VP.n15 161.3
R48 VP.n67 VP.n66 161.3
R49 VP.n30 VP.t7 141.222
R50 VP.n16 VP.t6 108.526
R51 VP.n12 VP.t1 108.526
R52 VP.n8 VP.t5 108.526
R53 VP.n4 VP.t8 108.526
R54 VP.n0 VP.t2 108.526
R55 VP.n17 VP.t3 108.526
R56 VP.n21 VP.t4 108.526
R57 VP.n25 VP.t9 108.526
R58 VP.n29 VP.t0 108.526
R59 VP.n65 VP.n16 76.7455
R60 VP.n110 VP.n0 76.7455
R61 VP.n64 VP.n17 76.7455
R62 VP.n30 VP.n29 61.3641
R63 VP.n65 VP.n64 58.0862
R64 VP.n69 VP.n14 41.8712
R65 VP.n106 VP.n2 41.8712
R66 VP.n60 VP.n19 41.8712
R67 VP.n80 VP.n10 40.8975
R68 VP.n95 VP.n6 40.8975
R69 VP.n49 VP.n23 40.8975
R70 VP.n34 VP.n27 40.8975
R71 VP.n84 VP.n10 39.9237
R72 VP.n91 VP.n6 39.9237
R73 VP.n45 VP.n23 39.9237
R74 VP.n38 VP.n27 39.9237
R75 VP.n73 VP.n14 38.95
R76 VP.n102 VP.n2 38.95
R77 VP.n56 VP.n19 38.95
R78 VP.n68 VP.n67 24.3439
R79 VP.n69 VP.n68 24.3439
R80 VP.n74 VP.n73 24.3439
R81 VP.n75 VP.n74 24.3439
R82 VP.n79 VP.n78 24.3439
R83 VP.n80 VP.n79 24.3439
R84 VP.n85 VP.n84 24.3439
R85 VP.n86 VP.n85 24.3439
R86 VP.n90 VP.n89 24.3439
R87 VP.n91 VP.n90 24.3439
R88 VP.n96 VP.n95 24.3439
R89 VP.n97 VP.n96 24.3439
R90 VP.n101 VP.n100 24.3439
R91 VP.n102 VP.n101 24.3439
R92 VP.n107 VP.n106 24.3439
R93 VP.n108 VP.n107 24.3439
R94 VP.n61 VP.n60 24.3439
R95 VP.n62 VP.n61 24.3439
R96 VP.n50 VP.n49 24.3439
R97 VP.n51 VP.n50 24.3439
R98 VP.n55 VP.n54 24.3439
R99 VP.n56 VP.n55 24.3439
R100 VP.n39 VP.n38 24.3439
R101 VP.n40 VP.n39 24.3439
R102 VP.n44 VP.n43 24.3439
R103 VP.n45 VP.n44 24.3439
R104 VP.n33 VP.n32 24.3439
R105 VP.n34 VP.n33 24.3439
R106 VP.n67 VP.n16 13.146
R107 VP.n108 VP.n0 13.146
R108 VP.n62 VP.n17 13.146
R109 VP.n78 VP.n12 12.6591
R110 VP.n97 VP.n4 12.6591
R111 VP.n51 VP.n21 12.6591
R112 VP.n32 VP.n29 12.6591
R113 VP.n86 VP.n8 12.1722
R114 VP.n89 VP.n8 12.1722
R115 VP.n40 VP.n25 12.1722
R116 VP.n43 VP.n25 12.1722
R117 VP.n75 VP.n12 11.6853
R118 VP.n100 VP.n4 11.6853
R119 VP.n54 VP.n21 11.6853
R120 VP.n31 VP.n30 4.24426
R121 VP.n64 VP.n63 0.355081
R122 VP.n66 VP.n65 0.355081
R123 VP.n110 VP.n109 0.355081
R124 VP VP.n110 0.26685
R125 VP.n31 VP.n28 0.189894
R126 VP.n35 VP.n28 0.189894
R127 VP.n36 VP.n35 0.189894
R128 VP.n37 VP.n36 0.189894
R129 VP.n37 VP.n26 0.189894
R130 VP.n41 VP.n26 0.189894
R131 VP.n42 VP.n41 0.189894
R132 VP.n42 VP.n24 0.189894
R133 VP.n46 VP.n24 0.189894
R134 VP.n47 VP.n46 0.189894
R135 VP.n48 VP.n47 0.189894
R136 VP.n48 VP.n22 0.189894
R137 VP.n52 VP.n22 0.189894
R138 VP.n53 VP.n52 0.189894
R139 VP.n53 VP.n20 0.189894
R140 VP.n57 VP.n20 0.189894
R141 VP.n58 VP.n57 0.189894
R142 VP.n59 VP.n58 0.189894
R143 VP.n59 VP.n18 0.189894
R144 VP.n63 VP.n18 0.189894
R145 VP.n66 VP.n15 0.189894
R146 VP.n70 VP.n15 0.189894
R147 VP.n71 VP.n70 0.189894
R148 VP.n72 VP.n71 0.189894
R149 VP.n72 VP.n13 0.189894
R150 VP.n76 VP.n13 0.189894
R151 VP.n77 VP.n76 0.189894
R152 VP.n77 VP.n11 0.189894
R153 VP.n81 VP.n11 0.189894
R154 VP.n82 VP.n81 0.189894
R155 VP.n83 VP.n82 0.189894
R156 VP.n83 VP.n9 0.189894
R157 VP.n87 VP.n9 0.189894
R158 VP.n88 VP.n87 0.189894
R159 VP.n88 VP.n7 0.189894
R160 VP.n92 VP.n7 0.189894
R161 VP.n93 VP.n92 0.189894
R162 VP.n94 VP.n93 0.189894
R163 VP.n94 VP.n5 0.189894
R164 VP.n98 VP.n5 0.189894
R165 VP.n99 VP.n98 0.189894
R166 VP.n99 VP.n3 0.189894
R167 VP.n103 VP.n3 0.189894
R168 VP.n104 VP.n103 0.189894
R169 VP.n105 VP.n104 0.189894
R170 VP.n105 VP.n1 0.189894
R171 VP.n109 VP.n1 0.189894
R172 VDD1.n1 VDD1.t6 77.114
R173 VDD1.n3 VDD1.t7 77.1139
R174 VDD1.n5 VDD1.n4 74.0321
R175 VDD1.n1 VDD1.n0 71.8183
R176 VDD1.n7 VDD1.n6 71.8182
R177 VDD1.n3 VDD1.n2 71.8181
R178 VDD1.n7 VDD1.n5 52.5289
R179 VDD1.n6 VDD1.t5 2.2704
R180 VDD1.n6 VDD1.t8 2.2704
R181 VDD1.n0 VDD1.t1 2.2704
R182 VDD1.n0 VDD1.t2 2.2704
R183 VDD1.n4 VDD1.t3 2.2704
R184 VDD1.n4 VDD1.t9 2.2704
R185 VDD1.n2 VDD1.t0 2.2704
R186 VDD1.n2 VDD1.t4 2.2704
R187 VDD1 VDD1.n7 2.21171
R188 VDD1 VDD1.n1 0.815155
R189 VDD1.n5 VDD1.n3 0.701619
R190 VTAIL.n11 VTAIL.t0 57.4094
R191 VTAIL.n17 VTAIL.t5 57.4093
R192 VTAIL.n2 VTAIL.t17 57.4093
R193 VTAIL.n16 VTAIL.t16 57.4093
R194 VTAIL.n15 VTAIL.n14 55.1396
R195 VTAIL.n13 VTAIL.n12 55.1396
R196 VTAIL.n10 VTAIL.n9 55.1396
R197 VTAIL.n8 VTAIL.n7 55.1396
R198 VTAIL.n19 VTAIL.n18 55.1393
R199 VTAIL.n1 VTAIL.n0 55.1393
R200 VTAIL.n4 VTAIL.n3 55.1393
R201 VTAIL.n6 VTAIL.n5 55.1393
R202 VTAIL.n8 VTAIL.n6 30.7634
R203 VTAIL.n17 VTAIL.n16 27.7376
R204 VTAIL.n10 VTAIL.n8 3.02636
R205 VTAIL.n11 VTAIL.n10 3.02636
R206 VTAIL.n15 VTAIL.n13 3.02636
R207 VTAIL.n16 VTAIL.n15 3.02636
R208 VTAIL.n6 VTAIL.n4 3.02636
R209 VTAIL.n4 VTAIL.n2 3.02636
R210 VTAIL.n19 VTAIL.n17 3.02636
R211 VTAIL VTAIL.n1 2.32809
R212 VTAIL.n18 VTAIL.t7 2.2704
R213 VTAIL.n18 VTAIL.t2 2.2704
R214 VTAIL.n0 VTAIL.t9 2.2704
R215 VTAIL.n0 VTAIL.t1 2.2704
R216 VTAIL.n3 VTAIL.t14 2.2704
R217 VTAIL.n3 VTAIL.t11 2.2704
R218 VTAIL.n5 VTAIL.t13 2.2704
R219 VTAIL.n5 VTAIL.t18 2.2704
R220 VTAIL.n14 VTAIL.t10 2.2704
R221 VTAIL.n14 VTAIL.t15 2.2704
R222 VTAIL.n12 VTAIL.t12 2.2704
R223 VTAIL.n12 VTAIL.t19 2.2704
R224 VTAIL.n9 VTAIL.t3 2.2704
R225 VTAIL.n9 VTAIL.t8 2.2704
R226 VTAIL.n7 VTAIL.t4 2.2704
R227 VTAIL.n7 VTAIL.t6 2.2704
R228 VTAIL.n13 VTAIL.n11 1.98326
R229 VTAIL.n2 VTAIL.n1 1.98326
R230 VTAIL VTAIL.n19 0.698776
R231 VN.n94 VN.n93 161.3
R232 VN.n92 VN.n49 161.3
R233 VN.n91 VN.n90 161.3
R234 VN.n89 VN.n50 161.3
R235 VN.n88 VN.n87 161.3
R236 VN.n86 VN.n51 161.3
R237 VN.n85 VN.n84 161.3
R238 VN.n83 VN.n82 161.3
R239 VN.n81 VN.n53 161.3
R240 VN.n80 VN.n79 161.3
R241 VN.n78 VN.n54 161.3
R242 VN.n77 VN.n76 161.3
R243 VN.n75 VN.n55 161.3
R244 VN.n74 VN.n73 161.3
R245 VN.n72 VN.n71 161.3
R246 VN.n70 VN.n57 161.3
R247 VN.n69 VN.n68 161.3
R248 VN.n67 VN.n58 161.3
R249 VN.n66 VN.n65 161.3
R250 VN.n64 VN.n59 161.3
R251 VN.n63 VN.n62 161.3
R252 VN.n46 VN.n45 161.3
R253 VN.n44 VN.n1 161.3
R254 VN.n43 VN.n42 161.3
R255 VN.n41 VN.n2 161.3
R256 VN.n40 VN.n39 161.3
R257 VN.n38 VN.n3 161.3
R258 VN.n37 VN.n36 161.3
R259 VN.n35 VN.n34 161.3
R260 VN.n33 VN.n5 161.3
R261 VN.n32 VN.n31 161.3
R262 VN.n30 VN.n6 161.3
R263 VN.n29 VN.n28 161.3
R264 VN.n27 VN.n7 161.3
R265 VN.n26 VN.n25 161.3
R266 VN.n24 VN.n23 161.3
R267 VN.n22 VN.n9 161.3
R268 VN.n21 VN.n20 161.3
R269 VN.n19 VN.n10 161.3
R270 VN.n18 VN.n17 161.3
R271 VN.n16 VN.n11 161.3
R272 VN.n15 VN.n14 161.3
R273 VN.n61 VN.t6 141.224
R274 VN.n13 VN.t5 141.224
R275 VN.n12 VN.t0 108.526
R276 VN.n8 VN.t7 108.526
R277 VN.n4 VN.t3 108.526
R278 VN.n0 VN.t9 108.526
R279 VN.n60 VN.t8 108.526
R280 VN.n56 VN.t1 108.526
R281 VN.n52 VN.t2 108.526
R282 VN.n48 VN.t4 108.526
R283 VN.n47 VN.n0 76.7455
R284 VN.n95 VN.n48 76.7455
R285 VN.n13 VN.n12 61.3641
R286 VN.n61 VN.n60 61.3641
R287 VN VN.n95 58.2517
R288 VN.n43 VN.n2 41.8712
R289 VN.n91 VN.n50 41.8712
R290 VN.n17 VN.n10 40.8975
R291 VN.n32 VN.n6 40.8975
R292 VN.n65 VN.n58 40.8975
R293 VN.n80 VN.n54 40.8975
R294 VN.n21 VN.n10 39.9237
R295 VN.n28 VN.n6 39.9237
R296 VN.n69 VN.n58 39.9237
R297 VN.n76 VN.n54 39.9237
R298 VN.n39 VN.n2 38.95
R299 VN.n87 VN.n50 38.95
R300 VN.n16 VN.n15 24.3439
R301 VN.n17 VN.n16 24.3439
R302 VN.n22 VN.n21 24.3439
R303 VN.n23 VN.n22 24.3439
R304 VN.n27 VN.n26 24.3439
R305 VN.n28 VN.n27 24.3439
R306 VN.n33 VN.n32 24.3439
R307 VN.n34 VN.n33 24.3439
R308 VN.n38 VN.n37 24.3439
R309 VN.n39 VN.n38 24.3439
R310 VN.n44 VN.n43 24.3439
R311 VN.n45 VN.n44 24.3439
R312 VN.n65 VN.n64 24.3439
R313 VN.n64 VN.n63 24.3439
R314 VN.n76 VN.n75 24.3439
R315 VN.n75 VN.n74 24.3439
R316 VN.n71 VN.n70 24.3439
R317 VN.n70 VN.n69 24.3439
R318 VN.n87 VN.n86 24.3439
R319 VN.n86 VN.n85 24.3439
R320 VN.n82 VN.n81 24.3439
R321 VN.n81 VN.n80 24.3439
R322 VN.n93 VN.n92 24.3439
R323 VN.n92 VN.n91 24.3439
R324 VN.n45 VN.n0 13.146
R325 VN.n93 VN.n48 13.146
R326 VN.n15 VN.n12 12.6591
R327 VN.n34 VN.n4 12.6591
R328 VN.n63 VN.n60 12.6591
R329 VN.n82 VN.n52 12.6591
R330 VN.n23 VN.n8 12.1722
R331 VN.n26 VN.n8 12.1722
R332 VN.n74 VN.n56 12.1722
R333 VN.n71 VN.n56 12.1722
R334 VN.n37 VN.n4 11.6853
R335 VN.n85 VN.n52 11.6853
R336 VN.n62 VN.n61 4.24428
R337 VN.n14 VN.n13 4.24428
R338 VN.n95 VN.n94 0.355081
R339 VN.n47 VN.n46 0.355081
R340 VN VN.n47 0.26685
R341 VN.n94 VN.n49 0.189894
R342 VN.n90 VN.n49 0.189894
R343 VN.n90 VN.n89 0.189894
R344 VN.n89 VN.n88 0.189894
R345 VN.n88 VN.n51 0.189894
R346 VN.n84 VN.n51 0.189894
R347 VN.n84 VN.n83 0.189894
R348 VN.n83 VN.n53 0.189894
R349 VN.n79 VN.n53 0.189894
R350 VN.n79 VN.n78 0.189894
R351 VN.n78 VN.n77 0.189894
R352 VN.n77 VN.n55 0.189894
R353 VN.n73 VN.n55 0.189894
R354 VN.n73 VN.n72 0.189894
R355 VN.n72 VN.n57 0.189894
R356 VN.n68 VN.n57 0.189894
R357 VN.n68 VN.n67 0.189894
R358 VN.n67 VN.n66 0.189894
R359 VN.n66 VN.n59 0.189894
R360 VN.n62 VN.n59 0.189894
R361 VN.n14 VN.n11 0.189894
R362 VN.n18 VN.n11 0.189894
R363 VN.n19 VN.n18 0.189894
R364 VN.n20 VN.n19 0.189894
R365 VN.n20 VN.n9 0.189894
R366 VN.n24 VN.n9 0.189894
R367 VN.n25 VN.n24 0.189894
R368 VN.n25 VN.n7 0.189894
R369 VN.n29 VN.n7 0.189894
R370 VN.n30 VN.n29 0.189894
R371 VN.n31 VN.n30 0.189894
R372 VN.n31 VN.n5 0.189894
R373 VN.n35 VN.n5 0.189894
R374 VN.n36 VN.n35 0.189894
R375 VN.n36 VN.n3 0.189894
R376 VN.n40 VN.n3 0.189894
R377 VN.n41 VN.n40 0.189894
R378 VN.n42 VN.n41 0.189894
R379 VN.n42 VN.n1 0.189894
R380 VN.n46 VN.n1 0.189894
R381 VDD2.n1 VDD2.t4 77.1139
R382 VDD2.n4 VDD2.t5 74.0882
R383 VDD2.n3 VDD2.n2 74.0321
R384 VDD2 VDD2.n7 74.0294
R385 VDD2.n6 VDD2.n5 71.8183
R386 VDD2.n1 VDD2.n0 71.8181
R387 VDD2.n4 VDD2.n3 50.433
R388 VDD2.n6 VDD2.n4 3.02636
R389 VDD2.n7 VDD2.t1 2.2704
R390 VDD2.n7 VDD2.t3 2.2704
R391 VDD2.n5 VDD2.t7 2.2704
R392 VDD2.n5 VDD2.t8 2.2704
R393 VDD2.n2 VDD2.t6 2.2704
R394 VDD2.n2 VDD2.t0 2.2704
R395 VDD2.n0 VDD2.t9 2.2704
R396 VDD2.n0 VDD2.t2 2.2704
R397 VDD2 VDD2.n6 0.815155
R398 VDD2.n3 VDD2.n1 0.701619
R399 B.n733 B.n94 585
R400 B.n735 B.n734 585
R401 B.n736 B.n93 585
R402 B.n738 B.n737 585
R403 B.n739 B.n92 585
R404 B.n741 B.n740 585
R405 B.n742 B.n91 585
R406 B.n744 B.n743 585
R407 B.n745 B.n90 585
R408 B.n747 B.n746 585
R409 B.n748 B.n89 585
R410 B.n750 B.n749 585
R411 B.n751 B.n88 585
R412 B.n753 B.n752 585
R413 B.n754 B.n87 585
R414 B.n756 B.n755 585
R415 B.n757 B.n86 585
R416 B.n759 B.n758 585
R417 B.n760 B.n85 585
R418 B.n762 B.n761 585
R419 B.n763 B.n84 585
R420 B.n765 B.n764 585
R421 B.n766 B.n83 585
R422 B.n768 B.n767 585
R423 B.n769 B.n82 585
R424 B.n771 B.n770 585
R425 B.n772 B.n81 585
R426 B.n774 B.n773 585
R427 B.n775 B.n80 585
R428 B.n777 B.n776 585
R429 B.n778 B.n79 585
R430 B.n780 B.n779 585
R431 B.n781 B.n78 585
R432 B.n783 B.n782 585
R433 B.n784 B.n77 585
R434 B.n786 B.n785 585
R435 B.n787 B.n76 585
R436 B.n789 B.n788 585
R437 B.n790 B.n75 585
R438 B.n792 B.n791 585
R439 B.n793 B.n74 585
R440 B.n795 B.n794 585
R441 B.n796 B.n73 585
R442 B.n798 B.n797 585
R443 B.n799 B.n72 585
R444 B.n801 B.n800 585
R445 B.n802 B.n71 585
R446 B.n804 B.n803 585
R447 B.n806 B.n805 585
R448 B.n807 B.n67 585
R449 B.n809 B.n808 585
R450 B.n810 B.n66 585
R451 B.n812 B.n811 585
R452 B.n813 B.n65 585
R453 B.n815 B.n814 585
R454 B.n816 B.n64 585
R455 B.n818 B.n817 585
R456 B.n819 B.n61 585
R457 B.n822 B.n821 585
R458 B.n823 B.n60 585
R459 B.n825 B.n824 585
R460 B.n826 B.n59 585
R461 B.n828 B.n827 585
R462 B.n829 B.n58 585
R463 B.n831 B.n830 585
R464 B.n832 B.n57 585
R465 B.n834 B.n833 585
R466 B.n835 B.n56 585
R467 B.n837 B.n836 585
R468 B.n838 B.n55 585
R469 B.n840 B.n839 585
R470 B.n841 B.n54 585
R471 B.n843 B.n842 585
R472 B.n844 B.n53 585
R473 B.n846 B.n845 585
R474 B.n847 B.n52 585
R475 B.n849 B.n848 585
R476 B.n850 B.n51 585
R477 B.n852 B.n851 585
R478 B.n853 B.n50 585
R479 B.n855 B.n854 585
R480 B.n856 B.n49 585
R481 B.n858 B.n857 585
R482 B.n859 B.n48 585
R483 B.n861 B.n860 585
R484 B.n862 B.n47 585
R485 B.n864 B.n863 585
R486 B.n865 B.n46 585
R487 B.n867 B.n866 585
R488 B.n868 B.n45 585
R489 B.n870 B.n869 585
R490 B.n871 B.n44 585
R491 B.n873 B.n872 585
R492 B.n874 B.n43 585
R493 B.n876 B.n875 585
R494 B.n877 B.n42 585
R495 B.n879 B.n878 585
R496 B.n880 B.n41 585
R497 B.n882 B.n881 585
R498 B.n883 B.n40 585
R499 B.n885 B.n884 585
R500 B.n886 B.n39 585
R501 B.n888 B.n887 585
R502 B.n889 B.n38 585
R503 B.n891 B.n890 585
R504 B.n892 B.n37 585
R505 B.n732 B.n731 585
R506 B.n730 B.n95 585
R507 B.n729 B.n728 585
R508 B.n727 B.n96 585
R509 B.n726 B.n725 585
R510 B.n724 B.n97 585
R511 B.n723 B.n722 585
R512 B.n721 B.n98 585
R513 B.n720 B.n719 585
R514 B.n718 B.n99 585
R515 B.n717 B.n716 585
R516 B.n715 B.n100 585
R517 B.n714 B.n713 585
R518 B.n712 B.n101 585
R519 B.n711 B.n710 585
R520 B.n709 B.n102 585
R521 B.n708 B.n707 585
R522 B.n706 B.n103 585
R523 B.n705 B.n704 585
R524 B.n703 B.n104 585
R525 B.n702 B.n701 585
R526 B.n700 B.n105 585
R527 B.n699 B.n698 585
R528 B.n697 B.n106 585
R529 B.n696 B.n695 585
R530 B.n694 B.n107 585
R531 B.n693 B.n692 585
R532 B.n691 B.n108 585
R533 B.n690 B.n689 585
R534 B.n688 B.n109 585
R535 B.n687 B.n686 585
R536 B.n685 B.n110 585
R537 B.n684 B.n683 585
R538 B.n682 B.n111 585
R539 B.n681 B.n680 585
R540 B.n679 B.n112 585
R541 B.n678 B.n677 585
R542 B.n676 B.n113 585
R543 B.n675 B.n674 585
R544 B.n673 B.n114 585
R545 B.n672 B.n671 585
R546 B.n670 B.n115 585
R547 B.n669 B.n668 585
R548 B.n667 B.n116 585
R549 B.n666 B.n665 585
R550 B.n664 B.n117 585
R551 B.n663 B.n662 585
R552 B.n661 B.n118 585
R553 B.n660 B.n659 585
R554 B.n658 B.n119 585
R555 B.n657 B.n656 585
R556 B.n655 B.n120 585
R557 B.n654 B.n653 585
R558 B.n652 B.n121 585
R559 B.n651 B.n650 585
R560 B.n649 B.n122 585
R561 B.n648 B.n647 585
R562 B.n646 B.n123 585
R563 B.n645 B.n644 585
R564 B.n643 B.n124 585
R565 B.n642 B.n641 585
R566 B.n640 B.n125 585
R567 B.n639 B.n638 585
R568 B.n637 B.n126 585
R569 B.n636 B.n635 585
R570 B.n634 B.n127 585
R571 B.n633 B.n632 585
R572 B.n631 B.n128 585
R573 B.n630 B.n629 585
R574 B.n628 B.n129 585
R575 B.n627 B.n626 585
R576 B.n625 B.n130 585
R577 B.n624 B.n623 585
R578 B.n622 B.n131 585
R579 B.n621 B.n620 585
R580 B.n619 B.n132 585
R581 B.n618 B.n617 585
R582 B.n616 B.n133 585
R583 B.n615 B.n614 585
R584 B.n613 B.n134 585
R585 B.n612 B.n611 585
R586 B.n610 B.n135 585
R587 B.n609 B.n608 585
R588 B.n607 B.n136 585
R589 B.n606 B.n605 585
R590 B.n604 B.n137 585
R591 B.n603 B.n602 585
R592 B.n601 B.n138 585
R593 B.n600 B.n599 585
R594 B.n598 B.n139 585
R595 B.n597 B.n596 585
R596 B.n595 B.n140 585
R597 B.n594 B.n593 585
R598 B.n592 B.n141 585
R599 B.n591 B.n590 585
R600 B.n589 B.n142 585
R601 B.n588 B.n587 585
R602 B.n586 B.n143 585
R603 B.n585 B.n584 585
R604 B.n583 B.n144 585
R605 B.n582 B.n581 585
R606 B.n580 B.n145 585
R607 B.n579 B.n578 585
R608 B.n577 B.n146 585
R609 B.n576 B.n575 585
R610 B.n574 B.n147 585
R611 B.n573 B.n572 585
R612 B.n571 B.n148 585
R613 B.n570 B.n569 585
R614 B.n568 B.n149 585
R615 B.n567 B.n566 585
R616 B.n565 B.n150 585
R617 B.n564 B.n563 585
R618 B.n562 B.n151 585
R619 B.n561 B.n560 585
R620 B.n559 B.n152 585
R621 B.n558 B.n557 585
R622 B.n556 B.n153 585
R623 B.n555 B.n554 585
R624 B.n553 B.n154 585
R625 B.n552 B.n551 585
R626 B.n550 B.n155 585
R627 B.n549 B.n548 585
R628 B.n547 B.n156 585
R629 B.n546 B.n545 585
R630 B.n544 B.n157 585
R631 B.n543 B.n542 585
R632 B.n541 B.n158 585
R633 B.n540 B.n539 585
R634 B.n538 B.n159 585
R635 B.n537 B.n536 585
R636 B.n535 B.n160 585
R637 B.n534 B.n533 585
R638 B.n532 B.n161 585
R639 B.n531 B.n530 585
R640 B.n529 B.n162 585
R641 B.n528 B.n527 585
R642 B.n526 B.n163 585
R643 B.n525 B.n524 585
R644 B.n523 B.n164 585
R645 B.n522 B.n521 585
R646 B.n361 B.n222 585
R647 B.n363 B.n362 585
R648 B.n364 B.n221 585
R649 B.n366 B.n365 585
R650 B.n367 B.n220 585
R651 B.n369 B.n368 585
R652 B.n370 B.n219 585
R653 B.n372 B.n371 585
R654 B.n373 B.n218 585
R655 B.n375 B.n374 585
R656 B.n376 B.n217 585
R657 B.n378 B.n377 585
R658 B.n379 B.n216 585
R659 B.n381 B.n380 585
R660 B.n382 B.n215 585
R661 B.n384 B.n383 585
R662 B.n385 B.n214 585
R663 B.n387 B.n386 585
R664 B.n388 B.n213 585
R665 B.n390 B.n389 585
R666 B.n391 B.n212 585
R667 B.n393 B.n392 585
R668 B.n394 B.n211 585
R669 B.n396 B.n395 585
R670 B.n397 B.n210 585
R671 B.n399 B.n398 585
R672 B.n400 B.n209 585
R673 B.n402 B.n401 585
R674 B.n403 B.n208 585
R675 B.n405 B.n404 585
R676 B.n406 B.n207 585
R677 B.n408 B.n407 585
R678 B.n409 B.n206 585
R679 B.n411 B.n410 585
R680 B.n412 B.n205 585
R681 B.n414 B.n413 585
R682 B.n415 B.n204 585
R683 B.n417 B.n416 585
R684 B.n418 B.n203 585
R685 B.n420 B.n419 585
R686 B.n421 B.n202 585
R687 B.n423 B.n422 585
R688 B.n424 B.n201 585
R689 B.n426 B.n425 585
R690 B.n427 B.n200 585
R691 B.n429 B.n428 585
R692 B.n430 B.n199 585
R693 B.n432 B.n431 585
R694 B.n434 B.n433 585
R695 B.n435 B.n195 585
R696 B.n437 B.n436 585
R697 B.n438 B.n194 585
R698 B.n440 B.n439 585
R699 B.n441 B.n193 585
R700 B.n443 B.n442 585
R701 B.n444 B.n192 585
R702 B.n446 B.n445 585
R703 B.n447 B.n189 585
R704 B.n450 B.n449 585
R705 B.n451 B.n188 585
R706 B.n453 B.n452 585
R707 B.n454 B.n187 585
R708 B.n456 B.n455 585
R709 B.n457 B.n186 585
R710 B.n459 B.n458 585
R711 B.n460 B.n185 585
R712 B.n462 B.n461 585
R713 B.n463 B.n184 585
R714 B.n465 B.n464 585
R715 B.n466 B.n183 585
R716 B.n468 B.n467 585
R717 B.n469 B.n182 585
R718 B.n471 B.n470 585
R719 B.n472 B.n181 585
R720 B.n474 B.n473 585
R721 B.n475 B.n180 585
R722 B.n477 B.n476 585
R723 B.n478 B.n179 585
R724 B.n480 B.n479 585
R725 B.n481 B.n178 585
R726 B.n483 B.n482 585
R727 B.n484 B.n177 585
R728 B.n486 B.n485 585
R729 B.n487 B.n176 585
R730 B.n489 B.n488 585
R731 B.n490 B.n175 585
R732 B.n492 B.n491 585
R733 B.n493 B.n174 585
R734 B.n495 B.n494 585
R735 B.n496 B.n173 585
R736 B.n498 B.n497 585
R737 B.n499 B.n172 585
R738 B.n501 B.n500 585
R739 B.n502 B.n171 585
R740 B.n504 B.n503 585
R741 B.n505 B.n170 585
R742 B.n507 B.n506 585
R743 B.n508 B.n169 585
R744 B.n510 B.n509 585
R745 B.n511 B.n168 585
R746 B.n513 B.n512 585
R747 B.n514 B.n167 585
R748 B.n516 B.n515 585
R749 B.n517 B.n166 585
R750 B.n519 B.n518 585
R751 B.n520 B.n165 585
R752 B.n360 B.n359 585
R753 B.n358 B.n223 585
R754 B.n357 B.n356 585
R755 B.n355 B.n224 585
R756 B.n354 B.n353 585
R757 B.n352 B.n225 585
R758 B.n351 B.n350 585
R759 B.n349 B.n226 585
R760 B.n348 B.n347 585
R761 B.n346 B.n227 585
R762 B.n345 B.n344 585
R763 B.n343 B.n228 585
R764 B.n342 B.n341 585
R765 B.n340 B.n229 585
R766 B.n339 B.n338 585
R767 B.n337 B.n230 585
R768 B.n336 B.n335 585
R769 B.n334 B.n231 585
R770 B.n333 B.n332 585
R771 B.n331 B.n232 585
R772 B.n330 B.n329 585
R773 B.n328 B.n233 585
R774 B.n327 B.n326 585
R775 B.n325 B.n234 585
R776 B.n324 B.n323 585
R777 B.n322 B.n235 585
R778 B.n321 B.n320 585
R779 B.n319 B.n236 585
R780 B.n318 B.n317 585
R781 B.n316 B.n237 585
R782 B.n315 B.n314 585
R783 B.n313 B.n238 585
R784 B.n312 B.n311 585
R785 B.n310 B.n239 585
R786 B.n309 B.n308 585
R787 B.n307 B.n240 585
R788 B.n306 B.n305 585
R789 B.n304 B.n241 585
R790 B.n303 B.n302 585
R791 B.n301 B.n242 585
R792 B.n300 B.n299 585
R793 B.n298 B.n243 585
R794 B.n297 B.n296 585
R795 B.n295 B.n244 585
R796 B.n294 B.n293 585
R797 B.n292 B.n245 585
R798 B.n291 B.n290 585
R799 B.n289 B.n246 585
R800 B.n288 B.n287 585
R801 B.n286 B.n247 585
R802 B.n285 B.n284 585
R803 B.n283 B.n248 585
R804 B.n282 B.n281 585
R805 B.n280 B.n249 585
R806 B.n279 B.n278 585
R807 B.n277 B.n250 585
R808 B.n276 B.n275 585
R809 B.n274 B.n251 585
R810 B.n273 B.n272 585
R811 B.n271 B.n252 585
R812 B.n270 B.n269 585
R813 B.n268 B.n253 585
R814 B.n267 B.n266 585
R815 B.n265 B.n254 585
R816 B.n264 B.n263 585
R817 B.n262 B.n255 585
R818 B.n261 B.n260 585
R819 B.n259 B.n256 585
R820 B.n258 B.n257 585
R821 B.n2 B.n0 585
R822 B.n997 B.n1 585
R823 B.n996 B.n995 585
R824 B.n994 B.n3 585
R825 B.n993 B.n992 585
R826 B.n991 B.n4 585
R827 B.n990 B.n989 585
R828 B.n988 B.n5 585
R829 B.n987 B.n986 585
R830 B.n985 B.n6 585
R831 B.n984 B.n983 585
R832 B.n982 B.n7 585
R833 B.n981 B.n980 585
R834 B.n979 B.n8 585
R835 B.n978 B.n977 585
R836 B.n976 B.n9 585
R837 B.n975 B.n974 585
R838 B.n973 B.n10 585
R839 B.n972 B.n971 585
R840 B.n970 B.n11 585
R841 B.n969 B.n968 585
R842 B.n967 B.n12 585
R843 B.n966 B.n965 585
R844 B.n964 B.n13 585
R845 B.n963 B.n962 585
R846 B.n961 B.n14 585
R847 B.n960 B.n959 585
R848 B.n958 B.n15 585
R849 B.n957 B.n956 585
R850 B.n955 B.n16 585
R851 B.n954 B.n953 585
R852 B.n952 B.n17 585
R853 B.n951 B.n950 585
R854 B.n949 B.n18 585
R855 B.n948 B.n947 585
R856 B.n946 B.n19 585
R857 B.n945 B.n944 585
R858 B.n943 B.n20 585
R859 B.n942 B.n941 585
R860 B.n940 B.n21 585
R861 B.n939 B.n938 585
R862 B.n937 B.n22 585
R863 B.n936 B.n935 585
R864 B.n934 B.n23 585
R865 B.n933 B.n932 585
R866 B.n931 B.n24 585
R867 B.n930 B.n929 585
R868 B.n928 B.n25 585
R869 B.n927 B.n926 585
R870 B.n925 B.n26 585
R871 B.n924 B.n923 585
R872 B.n922 B.n27 585
R873 B.n921 B.n920 585
R874 B.n919 B.n28 585
R875 B.n918 B.n917 585
R876 B.n916 B.n29 585
R877 B.n915 B.n914 585
R878 B.n913 B.n30 585
R879 B.n912 B.n911 585
R880 B.n910 B.n31 585
R881 B.n909 B.n908 585
R882 B.n907 B.n32 585
R883 B.n906 B.n905 585
R884 B.n904 B.n33 585
R885 B.n903 B.n902 585
R886 B.n901 B.n34 585
R887 B.n900 B.n899 585
R888 B.n898 B.n35 585
R889 B.n897 B.n896 585
R890 B.n895 B.n36 585
R891 B.n894 B.n893 585
R892 B.n999 B.n998 585
R893 B.n361 B.n360 545.355
R894 B.n894 B.n37 545.355
R895 B.n522 B.n165 545.355
R896 B.n733 B.n732 545.355
R897 B.n190 B.t6 317.308
R898 B.n196 B.t0 317.308
R899 B.n62 B.t9 317.308
R900 B.n68 B.t3 317.308
R901 B.n190 B.t8 175.512
R902 B.n68 B.t4 175.512
R903 B.n196 B.t2 175.494
R904 B.n62 B.t10 175.494
R905 B.n360 B.n223 163.367
R906 B.n356 B.n223 163.367
R907 B.n356 B.n355 163.367
R908 B.n355 B.n354 163.367
R909 B.n354 B.n225 163.367
R910 B.n350 B.n225 163.367
R911 B.n350 B.n349 163.367
R912 B.n349 B.n348 163.367
R913 B.n348 B.n227 163.367
R914 B.n344 B.n227 163.367
R915 B.n344 B.n343 163.367
R916 B.n343 B.n342 163.367
R917 B.n342 B.n229 163.367
R918 B.n338 B.n229 163.367
R919 B.n338 B.n337 163.367
R920 B.n337 B.n336 163.367
R921 B.n336 B.n231 163.367
R922 B.n332 B.n231 163.367
R923 B.n332 B.n331 163.367
R924 B.n331 B.n330 163.367
R925 B.n330 B.n233 163.367
R926 B.n326 B.n233 163.367
R927 B.n326 B.n325 163.367
R928 B.n325 B.n324 163.367
R929 B.n324 B.n235 163.367
R930 B.n320 B.n235 163.367
R931 B.n320 B.n319 163.367
R932 B.n319 B.n318 163.367
R933 B.n318 B.n237 163.367
R934 B.n314 B.n237 163.367
R935 B.n314 B.n313 163.367
R936 B.n313 B.n312 163.367
R937 B.n312 B.n239 163.367
R938 B.n308 B.n239 163.367
R939 B.n308 B.n307 163.367
R940 B.n307 B.n306 163.367
R941 B.n306 B.n241 163.367
R942 B.n302 B.n241 163.367
R943 B.n302 B.n301 163.367
R944 B.n301 B.n300 163.367
R945 B.n300 B.n243 163.367
R946 B.n296 B.n243 163.367
R947 B.n296 B.n295 163.367
R948 B.n295 B.n294 163.367
R949 B.n294 B.n245 163.367
R950 B.n290 B.n245 163.367
R951 B.n290 B.n289 163.367
R952 B.n289 B.n288 163.367
R953 B.n288 B.n247 163.367
R954 B.n284 B.n247 163.367
R955 B.n284 B.n283 163.367
R956 B.n283 B.n282 163.367
R957 B.n282 B.n249 163.367
R958 B.n278 B.n249 163.367
R959 B.n278 B.n277 163.367
R960 B.n277 B.n276 163.367
R961 B.n276 B.n251 163.367
R962 B.n272 B.n251 163.367
R963 B.n272 B.n271 163.367
R964 B.n271 B.n270 163.367
R965 B.n270 B.n253 163.367
R966 B.n266 B.n253 163.367
R967 B.n266 B.n265 163.367
R968 B.n265 B.n264 163.367
R969 B.n264 B.n255 163.367
R970 B.n260 B.n255 163.367
R971 B.n260 B.n259 163.367
R972 B.n259 B.n258 163.367
R973 B.n258 B.n2 163.367
R974 B.n998 B.n2 163.367
R975 B.n998 B.n997 163.367
R976 B.n997 B.n996 163.367
R977 B.n996 B.n3 163.367
R978 B.n992 B.n3 163.367
R979 B.n992 B.n991 163.367
R980 B.n991 B.n990 163.367
R981 B.n990 B.n5 163.367
R982 B.n986 B.n5 163.367
R983 B.n986 B.n985 163.367
R984 B.n985 B.n984 163.367
R985 B.n984 B.n7 163.367
R986 B.n980 B.n7 163.367
R987 B.n980 B.n979 163.367
R988 B.n979 B.n978 163.367
R989 B.n978 B.n9 163.367
R990 B.n974 B.n9 163.367
R991 B.n974 B.n973 163.367
R992 B.n973 B.n972 163.367
R993 B.n972 B.n11 163.367
R994 B.n968 B.n11 163.367
R995 B.n968 B.n967 163.367
R996 B.n967 B.n966 163.367
R997 B.n966 B.n13 163.367
R998 B.n962 B.n13 163.367
R999 B.n962 B.n961 163.367
R1000 B.n961 B.n960 163.367
R1001 B.n960 B.n15 163.367
R1002 B.n956 B.n15 163.367
R1003 B.n956 B.n955 163.367
R1004 B.n955 B.n954 163.367
R1005 B.n954 B.n17 163.367
R1006 B.n950 B.n17 163.367
R1007 B.n950 B.n949 163.367
R1008 B.n949 B.n948 163.367
R1009 B.n948 B.n19 163.367
R1010 B.n944 B.n19 163.367
R1011 B.n944 B.n943 163.367
R1012 B.n943 B.n942 163.367
R1013 B.n942 B.n21 163.367
R1014 B.n938 B.n21 163.367
R1015 B.n938 B.n937 163.367
R1016 B.n937 B.n936 163.367
R1017 B.n936 B.n23 163.367
R1018 B.n932 B.n23 163.367
R1019 B.n932 B.n931 163.367
R1020 B.n931 B.n930 163.367
R1021 B.n930 B.n25 163.367
R1022 B.n926 B.n25 163.367
R1023 B.n926 B.n925 163.367
R1024 B.n925 B.n924 163.367
R1025 B.n924 B.n27 163.367
R1026 B.n920 B.n27 163.367
R1027 B.n920 B.n919 163.367
R1028 B.n919 B.n918 163.367
R1029 B.n918 B.n29 163.367
R1030 B.n914 B.n29 163.367
R1031 B.n914 B.n913 163.367
R1032 B.n913 B.n912 163.367
R1033 B.n912 B.n31 163.367
R1034 B.n908 B.n31 163.367
R1035 B.n908 B.n907 163.367
R1036 B.n907 B.n906 163.367
R1037 B.n906 B.n33 163.367
R1038 B.n902 B.n33 163.367
R1039 B.n902 B.n901 163.367
R1040 B.n901 B.n900 163.367
R1041 B.n900 B.n35 163.367
R1042 B.n896 B.n35 163.367
R1043 B.n896 B.n895 163.367
R1044 B.n895 B.n894 163.367
R1045 B.n362 B.n361 163.367
R1046 B.n362 B.n221 163.367
R1047 B.n366 B.n221 163.367
R1048 B.n367 B.n366 163.367
R1049 B.n368 B.n367 163.367
R1050 B.n368 B.n219 163.367
R1051 B.n372 B.n219 163.367
R1052 B.n373 B.n372 163.367
R1053 B.n374 B.n373 163.367
R1054 B.n374 B.n217 163.367
R1055 B.n378 B.n217 163.367
R1056 B.n379 B.n378 163.367
R1057 B.n380 B.n379 163.367
R1058 B.n380 B.n215 163.367
R1059 B.n384 B.n215 163.367
R1060 B.n385 B.n384 163.367
R1061 B.n386 B.n385 163.367
R1062 B.n386 B.n213 163.367
R1063 B.n390 B.n213 163.367
R1064 B.n391 B.n390 163.367
R1065 B.n392 B.n391 163.367
R1066 B.n392 B.n211 163.367
R1067 B.n396 B.n211 163.367
R1068 B.n397 B.n396 163.367
R1069 B.n398 B.n397 163.367
R1070 B.n398 B.n209 163.367
R1071 B.n402 B.n209 163.367
R1072 B.n403 B.n402 163.367
R1073 B.n404 B.n403 163.367
R1074 B.n404 B.n207 163.367
R1075 B.n408 B.n207 163.367
R1076 B.n409 B.n408 163.367
R1077 B.n410 B.n409 163.367
R1078 B.n410 B.n205 163.367
R1079 B.n414 B.n205 163.367
R1080 B.n415 B.n414 163.367
R1081 B.n416 B.n415 163.367
R1082 B.n416 B.n203 163.367
R1083 B.n420 B.n203 163.367
R1084 B.n421 B.n420 163.367
R1085 B.n422 B.n421 163.367
R1086 B.n422 B.n201 163.367
R1087 B.n426 B.n201 163.367
R1088 B.n427 B.n426 163.367
R1089 B.n428 B.n427 163.367
R1090 B.n428 B.n199 163.367
R1091 B.n432 B.n199 163.367
R1092 B.n433 B.n432 163.367
R1093 B.n433 B.n195 163.367
R1094 B.n437 B.n195 163.367
R1095 B.n438 B.n437 163.367
R1096 B.n439 B.n438 163.367
R1097 B.n439 B.n193 163.367
R1098 B.n443 B.n193 163.367
R1099 B.n444 B.n443 163.367
R1100 B.n445 B.n444 163.367
R1101 B.n445 B.n189 163.367
R1102 B.n450 B.n189 163.367
R1103 B.n451 B.n450 163.367
R1104 B.n452 B.n451 163.367
R1105 B.n452 B.n187 163.367
R1106 B.n456 B.n187 163.367
R1107 B.n457 B.n456 163.367
R1108 B.n458 B.n457 163.367
R1109 B.n458 B.n185 163.367
R1110 B.n462 B.n185 163.367
R1111 B.n463 B.n462 163.367
R1112 B.n464 B.n463 163.367
R1113 B.n464 B.n183 163.367
R1114 B.n468 B.n183 163.367
R1115 B.n469 B.n468 163.367
R1116 B.n470 B.n469 163.367
R1117 B.n470 B.n181 163.367
R1118 B.n474 B.n181 163.367
R1119 B.n475 B.n474 163.367
R1120 B.n476 B.n475 163.367
R1121 B.n476 B.n179 163.367
R1122 B.n480 B.n179 163.367
R1123 B.n481 B.n480 163.367
R1124 B.n482 B.n481 163.367
R1125 B.n482 B.n177 163.367
R1126 B.n486 B.n177 163.367
R1127 B.n487 B.n486 163.367
R1128 B.n488 B.n487 163.367
R1129 B.n488 B.n175 163.367
R1130 B.n492 B.n175 163.367
R1131 B.n493 B.n492 163.367
R1132 B.n494 B.n493 163.367
R1133 B.n494 B.n173 163.367
R1134 B.n498 B.n173 163.367
R1135 B.n499 B.n498 163.367
R1136 B.n500 B.n499 163.367
R1137 B.n500 B.n171 163.367
R1138 B.n504 B.n171 163.367
R1139 B.n505 B.n504 163.367
R1140 B.n506 B.n505 163.367
R1141 B.n506 B.n169 163.367
R1142 B.n510 B.n169 163.367
R1143 B.n511 B.n510 163.367
R1144 B.n512 B.n511 163.367
R1145 B.n512 B.n167 163.367
R1146 B.n516 B.n167 163.367
R1147 B.n517 B.n516 163.367
R1148 B.n518 B.n517 163.367
R1149 B.n518 B.n165 163.367
R1150 B.n523 B.n522 163.367
R1151 B.n524 B.n523 163.367
R1152 B.n524 B.n163 163.367
R1153 B.n528 B.n163 163.367
R1154 B.n529 B.n528 163.367
R1155 B.n530 B.n529 163.367
R1156 B.n530 B.n161 163.367
R1157 B.n534 B.n161 163.367
R1158 B.n535 B.n534 163.367
R1159 B.n536 B.n535 163.367
R1160 B.n536 B.n159 163.367
R1161 B.n540 B.n159 163.367
R1162 B.n541 B.n540 163.367
R1163 B.n542 B.n541 163.367
R1164 B.n542 B.n157 163.367
R1165 B.n546 B.n157 163.367
R1166 B.n547 B.n546 163.367
R1167 B.n548 B.n547 163.367
R1168 B.n548 B.n155 163.367
R1169 B.n552 B.n155 163.367
R1170 B.n553 B.n552 163.367
R1171 B.n554 B.n553 163.367
R1172 B.n554 B.n153 163.367
R1173 B.n558 B.n153 163.367
R1174 B.n559 B.n558 163.367
R1175 B.n560 B.n559 163.367
R1176 B.n560 B.n151 163.367
R1177 B.n564 B.n151 163.367
R1178 B.n565 B.n564 163.367
R1179 B.n566 B.n565 163.367
R1180 B.n566 B.n149 163.367
R1181 B.n570 B.n149 163.367
R1182 B.n571 B.n570 163.367
R1183 B.n572 B.n571 163.367
R1184 B.n572 B.n147 163.367
R1185 B.n576 B.n147 163.367
R1186 B.n577 B.n576 163.367
R1187 B.n578 B.n577 163.367
R1188 B.n578 B.n145 163.367
R1189 B.n582 B.n145 163.367
R1190 B.n583 B.n582 163.367
R1191 B.n584 B.n583 163.367
R1192 B.n584 B.n143 163.367
R1193 B.n588 B.n143 163.367
R1194 B.n589 B.n588 163.367
R1195 B.n590 B.n589 163.367
R1196 B.n590 B.n141 163.367
R1197 B.n594 B.n141 163.367
R1198 B.n595 B.n594 163.367
R1199 B.n596 B.n595 163.367
R1200 B.n596 B.n139 163.367
R1201 B.n600 B.n139 163.367
R1202 B.n601 B.n600 163.367
R1203 B.n602 B.n601 163.367
R1204 B.n602 B.n137 163.367
R1205 B.n606 B.n137 163.367
R1206 B.n607 B.n606 163.367
R1207 B.n608 B.n607 163.367
R1208 B.n608 B.n135 163.367
R1209 B.n612 B.n135 163.367
R1210 B.n613 B.n612 163.367
R1211 B.n614 B.n613 163.367
R1212 B.n614 B.n133 163.367
R1213 B.n618 B.n133 163.367
R1214 B.n619 B.n618 163.367
R1215 B.n620 B.n619 163.367
R1216 B.n620 B.n131 163.367
R1217 B.n624 B.n131 163.367
R1218 B.n625 B.n624 163.367
R1219 B.n626 B.n625 163.367
R1220 B.n626 B.n129 163.367
R1221 B.n630 B.n129 163.367
R1222 B.n631 B.n630 163.367
R1223 B.n632 B.n631 163.367
R1224 B.n632 B.n127 163.367
R1225 B.n636 B.n127 163.367
R1226 B.n637 B.n636 163.367
R1227 B.n638 B.n637 163.367
R1228 B.n638 B.n125 163.367
R1229 B.n642 B.n125 163.367
R1230 B.n643 B.n642 163.367
R1231 B.n644 B.n643 163.367
R1232 B.n644 B.n123 163.367
R1233 B.n648 B.n123 163.367
R1234 B.n649 B.n648 163.367
R1235 B.n650 B.n649 163.367
R1236 B.n650 B.n121 163.367
R1237 B.n654 B.n121 163.367
R1238 B.n655 B.n654 163.367
R1239 B.n656 B.n655 163.367
R1240 B.n656 B.n119 163.367
R1241 B.n660 B.n119 163.367
R1242 B.n661 B.n660 163.367
R1243 B.n662 B.n661 163.367
R1244 B.n662 B.n117 163.367
R1245 B.n666 B.n117 163.367
R1246 B.n667 B.n666 163.367
R1247 B.n668 B.n667 163.367
R1248 B.n668 B.n115 163.367
R1249 B.n672 B.n115 163.367
R1250 B.n673 B.n672 163.367
R1251 B.n674 B.n673 163.367
R1252 B.n674 B.n113 163.367
R1253 B.n678 B.n113 163.367
R1254 B.n679 B.n678 163.367
R1255 B.n680 B.n679 163.367
R1256 B.n680 B.n111 163.367
R1257 B.n684 B.n111 163.367
R1258 B.n685 B.n684 163.367
R1259 B.n686 B.n685 163.367
R1260 B.n686 B.n109 163.367
R1261 B.n690 B.n109 163.367
R1262 B.n691 B.n690 163.367
R1263 B.n692 B.n691 163.367
R1264 B.n692 B.n107 163.367
R1265 B.n696 B.n107 163.367
R1266 B.n697 B.n696 163.367
R1267 B.n698 B.n697 163.367
R1268 B.n698 B.n105 163.367
R1269 B.n702 B.n105 163.367
R1270 B.n703 B.n702 163.367
R1271 B.n704 B.n703 163.367
R1272 B.n704 B.n103 163.367
R1273 B.n708 B.n103 163.367
R1274 B.n709 B.n708 163.367
R1275 B.n710 B.n709 163.367
R1276 B.n710 B.n101 163.367
R1277 B.n714 B.n101 163.367
R1278 B.n715 B.n714 163.367
R1279 B.n716 B.n715 163.367
R1280 B.n716 B.n99 163.367
R1281 B.n720 B.n99 163.367
R1282 B.n721 B.n720 163.367
R1283 B.n722 B.n721 163.367
R1284 B.n722 B.n97 163.367
R1285 B.n726 B.n97 163.367
R1286 B.n727 B.n726 163.367
R1287 B.n728 B.n727 163.367
R1288 B.n728 B.n95 163.367
R1289 B.n732 B.n95 163.367
R1290 B.n890 B.n37 163.367
R1291 B.n890 B.n889 163.367
R1292 B.n889 B.n888 163.367
R1293 B.n888 B.n39 163.367
R1294 B.n884 B.n39 163.367
R1295 B.n884 B.n883 163.367
R1296 B.n883 B.n882 163.367
R1297 B.n882 B.n41 163.367
R1298 B.n878 B.n41 163.367
R1299 B.n878 B.n877 163.367
R1300 B.n877 B.n876 163.367
R1301 B.n876 B.n43 163.367
R1302 B.n872 B.n43 163.367
R1303 B.n872 B.n871 163.367
R1304 B.n871 B.n870 163.367
R1305 B.n870 B.n45 163.367
R1306 B.n866 B.n45 163.367
R1307 B.n866 B.n865 163.367
R1308 B.n865 B.n864 163.367
R1309 B.n864 B.n47 163.367
R1310 B.n860 B.n47 163.367
R1311 B.n860 B.n859 163.367
R1312 B.n859 B.n858 163.367
R1313 B.n858 B.n49 163.367
R1314 B.n854 B.n49 163.367
R1315 B.n854 B.n853 163.367
R1316 B.n853 B.n852 163.367
R1317 B.n852 B.n51 163.367
R1318 B.n848 B.n51 163.367
R1319 B.n848 B.n847 163.367
R1320 B.n847 B.n846 163.367
R1321 B.n846 B.n53 163.367
R1322 B.n842 B.n53 163.367
R1323 B.n842 B.n841 163.367
R1324 B.n841 B.n840 163.367
R1325 B.n840 B.n55 163.367
R1326 B.n836 B.n55 163.367
R1327 B.n836 B.n835 163.367
R1328 B.n835 B.n834 163.367
R1329 B.n834 B.n57 163.367
R1330 B.n830 B.n57 163.367
R1331 B.n830 B.n829 163.367
R1332 B.n829 B.n828 163.367
R1333 B.n828 B.n59 163.367
R1334 B.n824 B.n59 163.367
R1335 B.n824 B.n823 163.367
R1336 B.n823 B.n822 163.367
R1337 B.n822 B.n61 163.367
R1338 B.n817 B.n61 163.367
R1339 B.n817 B.n816 163.367
R1340 B.n816 B.n815 163.367
R1341 B.n815 B.n65 163.367
R1342 B.n811 B.n65 163.367
R1343 B.n811 B.n810 163.367
R1344 B.n810 B.n809 163.367
R1345 B.n809 B.n67 163.367
R1346 B.n805 B.n67 163.367
R1347 B.n805 B.n804 163.367
R1348 B.n804 B.n71 163.367
R1349 B.n800 B.n71 163.367
R1350 B.n800 B.n799 163.367
R1351 B.n799 B.n798 163.367
R1352 B.n798 B.n73 163.367
R1353 B.n794 B.n73 163.367
R1354 B.n794 B.n793 163.367
R1355 B.n793 B.n792 163.367
R1356 B.n792 B.n75 163.367
R1357 B.n788 B.n75 163.367
R1358 B.n788 B.n787 163.367
R1359 B.n787 B.n786 163.367
R1360 B.n786 B.n77 163.367
R1361 B.n782 B.n77 163.367
R1362 B.n782 B.n781 163.367
R1363 B.n781 B.n780 163.367
R1364 B.n780 B.n79 163.367
R1365 B.n776 B.n79 163.367
R1366 B.n776 B.n775 163.367
R1367 B.n775 B.n774 163.367
R1368 B.n774 B.n81 163.367
R1369 B.n770 B.n81 163.367
R1370 B.n770 B.n769 163.367
R1371 B.n769 B.n768 163.367
R1372 B.n768 B.n83 163.367
R1373 B.n764 B.n83 163.367
R1374 B.n764 B.n763 163.367
R1375 B.n763 B.n762 163.367
R1376 B.n762 B.n85 163.367
R1377 B.n758 B.n85 163.367
R1378 B.n758 B.n757 163.367
R1379 B.n757 B.n756 163.367
R1380 B.n756 B.n87 163.367
R1381 B.n752 B.n87 163.367
R1382 B.n752 B.n751 163.367
R1383 B.n751 B.n750 163.367
R1384 B.n750 B.n89 163.367
R1385 B.n746 B.n89 163.367
R1386 B.n746 B.n745 163.367
R1387 B.n745 B.n744 163.367
R1388 B.n744 B.n91 163.367
R1389 B.n740 B.n91 163.367
R1390 B.n740 B.n739 163.367
R1391 B.n739 B.n738 163.367
R1392 B.n738 B.n93 163.367
R1393 B.n734 B.n93 163.367
R1394 B.n734 B.n733 163.367
R1395 B.n191 B.t7 107.439
R1396 B.n69 B.t5 107.439
R1397 B.n197 B.t1 107.421
R1398 B.n63 B.t11 107.421
R1399 B.n191 B.n190 68.0732
R1400 B.n197 B.n196 68.0732
R1401 B.n63 B.n62 68.0732
R1402 B.n69 B.n68 68.0732
R1403 B.n448 B.n191 59.5399
R1404 B.n198 B.n197 59.5399
R1405 B.n820 B.n63 59.5399
R1406 B.n70 B.n69 59.5399
R1407 B.n893 B.n892 35.4346
R1408 B.n731 B.n94 35.4346
R1409 B.n521 B.n520 35.4346
R1410 B.n359 B.n222 35.4346
R1411 B B.n999 18.0485
R1412 B.n892 B.n891 10.6151
R1413 B.n891 B.n38 10.6151
R1414 B.n887 B.n38 10.6151
R1415 B.n887 B.n886 10.6151
R1416 B.n886 B.n885 10.6151
R1417 B.n885 B.n40 10.6151
R1418 B.n881 B.n40 10.6151
R1419 B.n881 B.n880 10.6151
R1420 B.n880 B.n879 10.6151
R1421 B.n879 B.n42 10.6151
R1422 B.n875 B.n42 10.6151
R1423 B.n875 B.n874 10.6151
R1424 B.n874 B.n873 10.6151
R1425 B.n873 B.n44 10.6151
R1426 B.n869 B.n44 10.6151
R1427 B.n869 B.n868 10.6151
R1428 B.n868 B.n867 10.6151
R1429 B.n867 B.n46 10.6151
R1430 B.n863 B.n46 10.6151
R1431 B.n863 B.n862 10.6151
R1432 B.n862 B.n861 10.6151
R1433 B.n861 B.n48 10.6151
R1434 B.n857 B.n48 10.6151
R1435 B.n857 B.n856 10.6151
R1436 B.n856 B.n855 10.6151
R1437 B.n855 B.n50 10.6151
R1438 B.n851 B.n50 10.6151
R1439 B.n851 B.n850 10.6151
R1440 B.n850 B.n849 10.6151
R1441 B.n849 B.n52 10.6151
R1442 B.n845 B.n52 10.6151
R1443 B.n845 B.n844 10.6151
R1444 B.n844 B.n843 10.6151
R1445 B.n843 B.n54 10.6151
R1446 B.n839 B.n54 10.6151
R1447 B.n839 B.n838 10.6151
R1448 B.n838 B.n837 10.6151
R1449 B.n837 B.n56 10.6151
R1450 B.n833 B.n56 10.6151
R1451 B.n833 B.n832 10.6151
R1452 B.n832 B.n831 10.6151
R1453 B.n831 B.n58 10.6151
R1454 B.n827 B.n58 10.6151
R1455 B.n827 B.n826 10.6151
R1456 B.n826 B.n825 10.6151
R1457 B.n825 B.n60 10.6151
R1458 B.n821 B.n60 10.6151
R1459 B.n819 B.n818 10.6151
R1460 B.n818 B.n64 10.6151
R1461 B.n814 B.n64 10.6151
R1462 B.n814 B.n813 10.6151
R1463 B.n813 B.n812 10.6151
R1464 B.n812 B.n66 10.6151
R1465 B.n808 B.n66 10.6151
R1466 B.n808 B.n807 10.6151
R1467 B.n807 B.n806 10.6151
R1468 B.n803 B.n802 10.6151
R1469 B.n802 B.n801 10.6151
R1470 B.n801 B.n72 10.6151
R1471 B.n797 B.n72 10.6151
R1472 B.n797 B.n796 10.6151
R1473 B.n796 B.n795 10.6151
R1474 B.n795 B.n74 10.6151
R1475 B.n791 B.n74 10.6151
R1476 B.n791 B.n790 10.6151
R1477 B.n790 B.n789 10.6151
R1478 B.n789 B.n76 10.6151
R1479 B.n785 B.n76 10.6151
R1480 B.n785 B.n784 10.6151
R1481 B.n784 B.n783 10.6151
R1482 B.n783 B.n78 10.6151
R1483 B.n779 B.n78 10.6151
R1484 B.n779 B.n778 10.6151
R1485 B.n778 B.n777 10.6151
R1486 B.n777 B.n80 10.6151
R1487 B.n773 B.n80 10.6151
R1488 B.n773 B.n772 10.6151
R1489 B.n772 B.n771 10.6151
R1490 B.n771 B.n82 10.6151
R1491 B.n767 B.n82 10.6151
R1492 B.n767 B.n766 10.6151
R1493 B.n766 B.n765 10.6151
R1494 B.n765 B.n84 10.6151
R1495 B.n761 B.n84 10.6151
R1496 B.n761 B.n760 10.6151
R1497 B.n760 B.n759 10.6151
R1498 B.n759 B.n86 10.6151
R1499 B.n755 B.n86 10.6151
R1500 B.n755 B.n754 10.6151
R1501 B.n754 B.n753 10.6151
R1502 B.n753 B.n88 10.6151
R1503 B.n749 B.n88 10.6151
R1504 B.n749 B.n748 10.6151
R1505 B.n748 B.n747 10.6151
R1506 B.n747 B.n90 10.6151
R1507 B.n743 B.n90 10.6151
R1508 B.n743 B.n742 10.6151
R1509 B.n742 B.n741 10.6151
R1510 B.n741 B.n92 10.6151
R1511 B.n737 B.n92 10.6151
R1512 B.n737 B.n736 10.6151
R1513 B.n736 B.n735 10.6151
R1514 B.n735 B.n94 10.6151
R1515 B.n521 B.n164 10.6151
R1516 B.n525 B.n164 10.6151
R1517 B.n526 B.n525 10.6151
R1518 B.n527 B.n526 10.6151
R1519 B.n527 B.n162 10.6151
R1520 B.n531 B.n162 10.6151
R1521 B.n532 B.n531 10.6151
R1522 B.n533 B.n532 10.6151
R1523 B.n533 B.n160 10.6151
R1524 B.n537 B.n160 10.6151
R1525 B.n538 B.n537 10.6151
R1526 B.n539 B.n538 10.6151
R1527 B.n539 B.n158 10.6151
R1528 B.n543 B.n158 10.6151
R1529 B.n544 B.n543 10.6151
R1530 B.n545 B.n544 10.6151
R1531 B.n545 B.n156 10.6151
R1532 B.n549 B.n156 10.6151
R1533 B.n550 B.n549 10.6151
R1534 B.n551 B.n550 10.6151
R1535 B.n551 B.n154 10.6151
R1536 B.n555 B.n154 10.6151
R1537 B.n556 B.n555 10.6151
R1538 B.n557 B.n556 10.6151
R1539 B.n557 B.n152 10.6151
R1540 B.n561 B.n152 10.6151
R1541 B.n562 B.n561 10.6151
R1542 B.n563 B.n562 10.6151
R1543 B.n563 B.n150 10.6151
R1544 B.n567 B.n150 10.6151
R1545 B.n568 B.n567 10.6151
R1546 B.n569 B.n568 10.6151
R1547 B.n569 B.n148 10.6151
R1548 B.n573 B.n148 10.6151
R1549 B.n574 B.n573 10.6151
R1550 B.n575 B.n574 10.6151
R1551 B.n575 B.n146 10.6151
R1552 B.n579 B.n146 10.6151
R1553 B.n580 B.n579 10.6151
R1554 B.n581 B.n580 10.6151
R1555 B.n581 B.n144 10.6151
R1556 B.n585 B.n144 10.6151
R1557 B.n586 B.n585 10.6151
R1558 B.n587 B.n586 10.6151
R1559 B.n587 B.n142 10.6151
R1560 B.n591 B.n142 10.6151
R1561 B.n592 B.n591 10.6151
R1562 B.n593 B.n592 10.6151
R1563 B.n593 B.n140 10.6151
R1564 B.n597 B.n140 10.6151
R1565 B.n598 B.n597 10.6151
R1566 B.n599 B.n598 10.6151
R1567 B.n599 B.n138 10.6151
R1568 B.n603 B.n138 10.6151
R1569 B.n604 B.n603 10.6151
R1570 B.n605 B.n604 10.6151
R1571 B.n605 B.n136 10.6151
R1572 B.n609 B.n136 10.6151
R1573 B.n610 B.n609 10.6151
R1574 B.n611 B.n610 10.6151
R1575 B.n611 B.n134 10.6151
R1576 B.n615 B.n134 10.6151
R1577 B.n616 B.n615 10.6151
R1578 B.n617 B.n616 10.6151
R1579 B.n617 B.n132 10.6151
R1580 B.n621 B.n132 10.6151
R1581 B.n622 B.n621 10.6151
R1582 B.n623 B.n622 10.6151
R1583 B.n623 B.n130 10.6151
R1584 B.n627 B.n130 10.6151
R1585 B.n628 B.n627 10.6151
R1586 B.n629 B.n628 10.6151
R1587 B.n629 B.n128 10.6151
R1588 B.n633 B.n128 10.6151
R1589 B.n634 B.n633 10.6151
R1590 B.n635 B.n634 10.6151
R1591 B.n635 B.n126 10.6151
R1592 B.n639 B.n126 10.6151
R1593 B.n640 B.n639 10.6151
R1594 B.n641 B.n640 10.6151
R1595 B.n641 B.n124 10.6151
R1596 B.n645 B.n124 10.6151
R1597 B.n646 B.n645 10.6151
R1598 B.n647 B.n646 10.6151
R1599 B.n647 B.n122 10.6151
R1600 B.n651 B.n122 10.6151
R1601 B.n652 B.n651 10.6151
R1602 B.n653 B.n652 10.6151
R1603 B.n653 B.n120 10.6151
R1604 B.n657 B.n120 10.6151
R1605 B.n658 B.n657 10.6151
R1606 B.n659 B.n658 10.6151
R1607 B.n659 B.n118 10.6151
R1608 B.n663 B.n118 10.6151
R1609 B.n664 B.n663 10.6151
R1610 B.n665 B.n664 10.6151
R1611 B.n665 B.n116 10.6151
R1612 B.n669 B.n116 10.6151
R1613 B.n670 B.n669 10.6151
R1614 B.n671 B.n670 10.6151
R1615 B.n671 B.n114 10.6151
R1616 B.n675 B.n114 10.6151
R1617 B.n676 B.n675 10.6151
R1618 B.n677 B.n676 10.6151
R1619 B.n677 B.n112 10.6151
R1620 B.n681 B.n112 10.6151
R1621 B.n682 B.n681 10.6151
R1622 B.n683 B.n682 10.6151
R1623 B.n683 B.n110 10.6151
R1624 B.n687 B.n110 10.6151
R1625 B.n688 B.n687 10.6151
R1626 B.n689 B.n688 10.6151
R1627 B.n689 B.n108 10.6151
R1628 B.n693 B.n108 10.6151
R1629 B.n694 B.n693 10.6151
R1630 B.n695 B.n694 10.6151
R1631 B.n695 B.n106 10.6151
R1632 B.n699 B.n106 10.6151
R1633 B.n700 B.n699 10.6151
R1634 B.n701 B.n700 10.6151
R1635 B.n701 B.n104 10.6151
R1636 B.n705 B.n104 10.6151
R1637 B.n706 B.n705 10.6151
R1638 B.n707 B.n706 10.6151
R1639 B.n707 B.n102 10.6151
R1640 B.n711 B.n102 10.6151
R1641 B.n712 B.n711 10.6151
R1642 B.n713 B.n712 10.6151
R1643 B.n713 B.n100 10.6151
R1644 B.n717 B.n100 10.6151
R1645 B.n718 B.n717 10.6151
R1646 B.n719 B.n718 10.6151
R1647 B.n719 B.n98 10.6151
R1648 B.n723 B.n98 10.6151
R1649 B.n724 B.n723 10.6151
R1650 B.n725 B.n724 10.6151
R1651 B.n725 B.n96 10.6151
R1652 B.n729 B.n96 10.6151
R1653 B.n730 B.n729 10.6151
R1654 B.n731 B.n730 10.6151
R1655 B.n363 B.n222 10.6151
R1656 B.n364 B.n363 10.6151
R1657 B.n365 B.n364 10.6151
R1658 B.n365 B.n220 10.6151
R1659 B.n369 B.n220 10.6151
R1660 B.n370 B.n369 10.6151
R1661 B.n371 B.n370 10.6151
R1662 B.n371 B.n218 10.6151
R1663 B.n375 B.n218 10.6151
R1664 B.n376 B.n375 10.6151
R1665 B.n377 B.n376 10.6151
R1666 B.n377 B.n216 10.6151
R1667 B.n381 B.n216 10.6151
R1668 B.n382 B.n381 10.6151
R1669 B.n383 B.n382 10.6151
R1670 B.n383 B.n214 10.6151
R1671 B.n387 B.n214 10.6151
R1672 B.n388 B.n387 10.6151
R1673 B.n389 B.n388 10.6151
R1674 B.n389 B.n212 10.6151
R1675 B.n393 B.n212 10.6151
R1676 B.n394 B.n393 10.6151
R1677 B.n395 B.n394 10.6151
R1678 B.n395 B.n210 10.6151
R1679 B.n399 B.n210 10.6151
R1680 B.n400 B.n399 10.6151
R1681 B.n401 B.n400 10.6151
R1682 B.n401 B.n208 10.6151
R1683 B.n405 B.n208 10.6151
R1684 B.n406 B.n405 10.6151
R1685 B.n407 B.n406 10.6151
R1686 B.n407 B.n206 10.6151
R1687 B.n411 B.n206 10.6151
R1688 B.n412 B.n411 10.6151
R1689 B.n413 B.n412 10.6151
R1690 B.n413 B.n204 10.6151
R1691 B.n417 B.n204 10.6151
R1692 B.n418 B.n417 10.6151
R1693 B.n419 B.n418 10.6151
R1694 B.n419 B.n202 10.6151
R1695 B.n423 B.n202 10.6151
R1696 B.n424 B.n423 10.6151
R1697 B.n425 B.n424 10.6151
R1698 B.n425 B.n200 10.6151
R1699 B.n429 B.n200 10.6151
R1700 B.n430 B.n429 10.6151
R1701 B.n431 B.n430 10.6151
R1702 B.n435 B.n434 10.6151
R1703 B.n436 B.n435 10.6151
R1704 B.n436 B.n194 10.6151
R1705 B.n440 B.n194 10.6151
R1706 B.n441 B.n440 10.6151
R1707 B.n442 B.n441 10.6151
R1708 B.n442 B.n192 10.6151
R1709 B.n446 B.n192 10.6151
R1710 B.n447 B.n446 10.6151
R1711 B.n449 B.n188 10.6151
R1712 B.n453 B.n188 10.6151
R1713 B.n454 B.n453 10.6151
R1714 B.n455 B.n454 10.6151
R1715 B.n455 B.n186 10.6151
R1716 B.n459 B.n186 10.6151
R1717 B.n460 B.n459 10.6151
R1718 B.n461 B.n460 10.6151
R1719 B.n461 B.n184 10.6151
R1720 B.n465 B.n184 10.6151
R1721 B.n466 B.n465 10.6151
R1722 B.n467 B.n466 10.6151
R1723 B.n467 B.n182 10.6151
R1724 B.n471 B.n182 10.6151
R1725 B.n472 B.n471 10.6151
R1726 B.n473 B.n472 10.6151
R1727 B.n473 B.n180 10.6151
R1728 B.n477 B.n180 10.6151
R1729 B.n478 B.n477 10.6151
R1730 B.n479 B.n478 10.6151
R1731 B.n479 B.n178 10.6151
R1732 B.n483 B.n178 10.6151
R1733 B.n484 B.n483 10.6151
R1734 B.n485 B.n484 10.6151
R1735 B.n485 B.n176 10.6151
R1736 B.n489 B.n176 10.6151
R1737 B.n490 B.n489 10.6151
R1738 B.n491 B.n490 10.6151
R1739 B.n491 B.n174 10.6151
R1740 B.n495 B.n174 10.6151
R1741 B.n496 B.n495 10.6151
R1742 B.n497 B.n496 10.6151
R1743 B.n497 B.n172 10.6151
R1744 B.n501 B.n172 10.6151
R1745 B.n502 B.n501 10.6151
R1746 B.n503 B.n502 10.6151
R1747 B.n503 B.n170 10.6151
R1748 B.n507 B.n170 10.6151
R1749 B.n508 B.n507 10.6151
R1750 B.n509 B.n508 10.6151
R1751 B.n509 B.n168 10.6151
R1752 B.n513 B.n168 10.6151
R1753 B.n514 B.n513 10.6151
R1754 B.n515 B.n514 10.6151
R1755 B.n515 B.n166 10.6151
R1756 B.n519 B.n166 10.6151
R1757 B.n520 B.n519 10.6151
R1758 B.n359 B.n358 10.6151
R1759 B.n358 B.n357 10.6151
R1760 B.n357 B.n224 10.6151
R1761 B.n353 B.n224 10.6151
R1762 B.n353 B.n352 10.6151
R1763 B.n352 B.n351 10.6151
R1764 B.n351 B.n226 10.6151
R1765 B.n347 B.n226 10.6151
R1766 B.n347 B.n346 10.6151
R1767 B.n346 B.n345 10.6151
R1768 B.n345 B.n228 10.6151
R1769 B.n341 B.n228 10.6151
R1770 B.n341 B.n340 10.6151
R1771 B.n340 B.n339 10.6151
R1772 B.n339 B.n230 10.6151
R1773 B.n335 B.n230 10.6151
R1774 B.n335 B.n334 10.6151
R1775 B.n334 B.n333 10.6151
R1776 B.n333 B.n232 10.6151
R1777 B.n329 B.n232 10.6151
R1778 B.n329 B.n328 10.6151
R1779 B.n328 B.n327 10.6151
R1780 B.n327 B.n234 10.6151
R1781 B.n323 B.n234 10.6151
R1782 B.n323 B.n322 10.6151
R1783 B.n322 B.n321 10.6151
R1784 B.n321 B.n236 10.6151
R1785 B.n317 B.n236 10.6151
R1786 B.n317 B.n316 10.6151
R1787 B.n316 B.n315 10.6151
R1788 B.n315 B.n238 10.6151
R1789 B.n311 B.n238 10.6151
R1790 B.n311 B.n310 10.6151
R1791 B.n310 B.n309 10.6151
R1792 B.n309 B.n240 10.6151
R1793 B.n305 B.n240 10.6151
R1794 B.n305 B.n304 10.6151
R1795 B.n304 B.n303 10.6151
R1796 B.n303 B.n242 10.6151
R1797 B.n299 B.n242 10.6151
R1798 B.n299 B.n298 10.6151
R1799 B.n298 B.n297 10.6151
R1800 B.n297 B.n244 10.6151
R1801 B.n293 B.n244 10.6151
R1802 B.n293 B.n292 10.6151
R1803 B.n292 B.n291 10.6151
R1804 B.n291 B.n246 10.6151
R1805 B.n287 B.n246 10.6151
R1806 B.n287 B.n286 10.6151
R1807 B.n286 B.n285 10.6151
R1808 B.n285 B.n248 10.6151
R1809 B.n281 B.n248 10.6151
R1810 B.n281 B.n280 10.6151
R1811 B.n280 B.n279 10.6151
R1812 B.n279 B.n250 10.6151
R1813 B.n275 B.n250 10.6151
R1814 B.n275 B.n274 10.6151
R1815 B.n274 B.n273 10.6151
R1816 B.n273 B.n252 10.6151
R1817 B.n269 B.n252 10.6151
R1818 B.n269 B.n268 10.6151
R1819 B.n268 B.n267 10.6151
R1820 B.n267 B.n254 10.6151
R1821 B.n263 B.n254 10.6151
R1822 B.n263 B.n262 10.6151
R1823 B.n262 B.n261 10.6151
R1824 B.n261 B.n256 10.6151
R1825 B.n257 B.n256 10.6151
R1826 B.n257 B.n0 10.6151
R1827 B.n995 B.n1 10.6151
R1828 B.n995 B.n994 10.6151
R1829 B.n994 B.n993 10.6151
R1830 B.n993 B.n4 10.6151
R1831 B.n989 B.n4 10.6151
R1832 B.n989 B.n988 10.6151
R1833 B.n988 B.n987 10.6151
R1834 B.n987 B.n6 10.6151
R1835 B.n983 B.n6 10.6151
R1836 B.n983 B.n982 10.6151
R1837 B.n982 B.n981 10.6151
R1838 B.n981 B.n8 10.6151
R1839 B.n977 B.n8 10.6151
R1840 B.n977 B.n976 10.6151
R1841 B.n976 B.n975 10.6151
R1842 B.n975 B.n10 10.6151
R1843 B.n971 B.n10 10.6151
R1844 B.n971 B.n970 10.6151
R1845 B.n970 B.n969 10.6151
R1846 B.n969 B.n12 10.6151
R1847 B.n965 B.n12 10.6151
R1848 B.n965 B.n964 10.6151
R1849 B.n964 B.n963 10.6151
R1850 B.n963 B.n14 10.6151
R1851 B.n959 B.n14 10.6151
R1852 B.n959 B.n958 10.6151
R1853 B.n958 B.n957 10.6151
R1854 B.n957 B.n16 10.6151
R1855 B.n953 B.n16 10.6151
R1856 B.n953 B.n952 10.6151
R1857 B.n952 B.n951 10.6151
R1858 B.n951 B.n18 10.6151
R1859 B.n947 B.n18 10.6151
R1860 B.n947 B.n946 10.6151
R1861 B.n946 B.n945 10.6151
R1862 B.n945 B.n20 10.6151
R1863 B.n941 B.n20 10.6151
R1864 B.n941 B.n940 10.6151
R1865 B.n940 B.n939 10.6151
R1866 B.n939 B.n22 10.6151
R1867 B.n935 B.n22 10.6151
R1868 B.n935 B.n934 10.6151
R1869 B.n934 B.n933 10.6151
R1870 B.n933 B.n24 10.6151
R1871 B.n929 B.n24 10.6151
R1872 B.n929 B.n928 10.6151
R1873 B.n928 B.n927 10.6151
R1874 B.n927 B.n26 10.6151
R1875 B.n923 B.n26 10.6151
R1876 B.n923 B.n922 10.6151
R1877 B.n922 B.n921 10.6151
R1878 B.n921 B.n28 10.6151
R1879 B.n917 B.n28 10.6151
R1880 B.n917 B.n916 10.6151
R1881 B.n916 B.n915 10.6151
R1882 B.n915 B.n30 10.6151
R1883 B.n911 B.n30 10.6151
R1884 B.n911 B.n910 10.6151
R1885 B.n910 B.n909 10.6151
R1886 B.n909 B.n32 10.6151
R1887 B.n905 B.n32 10.6151
R1888 B.n905 B.n904 10.6151
R1889 B.n904 B.n903 10.6151
R1890 B.n903 B.n34 10.6151
R1891 B.n899 B.n34 10.6151
R1892 B.n899 B.n898 10.6151
R1893 B.n898 B.n897 10.6151
R1894 B.n897 B.n36 10.6151
R1895 B.n893 B.n36 10.6151
R1896 B.n821 B.n820 9.36635
R1897 B.n803 B.n70 9.36635
R1898 B.n431 B.n198 9.36635
R1899 B.n449 B.n448 9.36635
R1900 B.n999 B.n0 2.81026
R1901 B.n999 B.n1 2.81026
R1902 B.n820 B.n819 1.24928
R1903 B.n806 B.n70 1.24928
R1904 B.n434 B.n198 1.24928
R1905 B.n448 B.n447 1.24928
C0 VP VDD2 0.657002f
C1 VTAIL w_n5182_n3832# 3.59763f
C2 VDD1 VTAIL 11.5843f
C3 VDD2 VN 13.113f
C4 VTAIL B 4.49802f
C5 w_n5182_n3832# VP 12.0133f
C6 VDD1 VP 13.6118f
C7 B VP 2.59453f
C8 w_n5182_n3832# VN 11.3368f
C9 VDD1 VN 0.153955f
C10 B VN 1.45383f
C11 w_n5182_n3832# VDD2 3.336f
C12 VDD1 VDD2 2.5496f
C13 B VDD2 3.03275f
C14 VTAIL VP 13.9112f
C15 VDD1 w_n5182_n3832# 3.1623f
C16 VTAIL VN 13.8969f
C17 w_n5182_n3832# B 12.172501f
C18 VDD1 B 2.89225f
C19 VTAIL VDD2 11.6392f
C20 VP VN 9.69514f
C21 VDD2 VSUBS 2.41204f
C22 VDD1 VSUBS 2.256973f
C23 VTAIL VSUBS 1.521365f
C24 VN VSUBS 8.712911f
C25 VP VSUBS 5.061552f
C26 B VSUBS 6.281902f
C27 w_n5182_n3832# VSUBS 0.243699p
C28 B.n0 VSUBS 0.005367f
C29 B.n1 VSUBS 0.005367f
C30 B.n2 VSUBS 0.008488f
C31 B.n3 VSUBS 0.008488f
C32 B.n4 VSUBS 0.008488f
C33 B.n5 VSUBS 0.008488f
C34 B.n6 VSUBS 0.008488f
C35 B.n7 VSUBS 0.008488f
C36 B.n8 VSUBS 0.008488f
C37 B.n9 VSUBS 0.008488f
C38 B.n10 VSUBS 0.008488f
C39 B.n11 VSUBS 0.008488f
C40 B.n12 VSUBS 0.008488f
C41 B.n13 VSUBS 0.008488f
C42 B.n14 VSUBS 0.008488f
C43 B.n15 VSUBS 0.008488f
C44 B.n16 VSUBS 0.008488f
C45 B.n17 VSUBS 0.008488f
C46 B.n18 VSUBS 0.008488f
C47 B.n19 VSUBS 0.008488f
C48 B.n20 VSUBS 0.008488f
C49 B.n21 VSUBS 0.008488f
C50 B.n22 VSUBS 0.008488f
C51 B.n23 VSUBS 0.008488f
C52 B.n24 VSUBS 0.008488f
C53 B.n25 VSUBS 0.008488f
C54 B.n26 VSUBS 0.008488f
C55 B.n27 VSUBS 0.008488f
C56 B.n28 VSUBS 0.008488f
C57 B.n29 VSUBS 0.008488f
C58 B.n30 VSUBS 0.008488f
C59 B.n31 VSUBS 0.008488f
C60 B.n32 VSUBS 0.008488f
C61 B.n33 VSUBS 0.008488f
C62 B.n34 VSUBS 0.008488f
C63 B.n35 VSUBS 0.008488f
C64 B.n36 VSUBS 0.008488f
C65 B.n37 VSUBS 0.021275f
C66 B.n38 VSUBS 0.008488f
C67 B.n39 VSUBS 0.008488f
C68 B.n40 VSUBS 0.008488f
C69 B.n41 VSUBS 0.008488f
C70 B.n42 VSUBS 0.008488f
C71 B.n43 VSUBS 0.008488f
C72 B.n44 VSUBS 0.008488f
C73 B.n45 VSUBS 0.008488f
C74 B.n46 VSUBS 0.008488f
C75 B.n47 VSUBS 0.008488f
C76 B.n48 VSUBS 0.008488f
C77 B.n49 VSUBS 0.008488f
C78 B.n50 VSUBS 0.008488f
C79 B.n51 VSUBS 0.008488f
C80 B.n52 VSUBS 0.008488f
C81 B.n53 VSUBS 0.008488f
C82 B.n54 VSUBS 0.008488f
C83 B.n55 VSUBS 0.008488f
C84 B.n56 VSUBS 0.008488f
C85 B.n57 VSUBS 0.008488f
C86 B.n58 VSUBS 0.008488f
C87 B.n59 VSUBS 0.008488f
C88 B.n60 VSUBS 0.008488f
C89 B.n61 VSUBS 0.008488f
C90 B.t11 VSUBS 0.575692f
C91 B.t10 VSUBS 0.605977f
C92 B.t9 VSUBS 2.52169f
C93 B.n62 VSUBS 0.340763f
C94 B.n63 VSUBS 0.090181f
C95 B.n64 VSUBS 0.008488f
C96 B.n65 VSUBS 0.008488f
C97 B.n66 VSUBS 0.008488f
C98 B.n67 VSUBS 0.008488f
C99 B.t5 VSUBS 0.575677f
C100 B.t4 VSUBS 0.605964f
C101 B.t3 VSUBS 2.52169f
C102 B.n68 VSUBS 0.340775f
C103 B.n69 VSUBS 0.090197f
C104 B.n70 VSUBS 0.019666f
C105 B.n71 VSUBS 0.008488f
C106 B.n72 VSUBS 0.008488f
C107 B.n73 VSUBS 0.008488f
C108 B.n74 VSUBS 0.008488f
C109 B.n75 VSUBS 0.008488f
C110 B.n76 VSUBS 0.008488f
C111 B.n77 VSUBS 0.008488f
C112 B.n78 VSUBS 0.008488f
C113 B.n79 VSUBS 0.008488f
C114 B.n80 VSUBS 0.008488f
C115 B.n81 VSUBS 0.008488f
C116 B.n82 VSUBS 0.008488f
C117 B.n83 VSUBS 0.008488f
C118 B.n84 VSUBS 0.008488f
C119 B.n85 VSUBS 0.008488f
C120 B.n86 VSUBS 0.008488f
C121 B.n87 VSUBS 0.008488f
C122 B.n88 VSUBS 0.008488f
C123 B.n89 VSUBS 0.008488f
C124 B.n90 VSUBS 0.008488f
C125 B.n91 VSUBS 0.008488f
C126 B.n92 VSUBS 0.008488f
C127 B.n93 VSUBS 0.008488f
C128 B.n94 VSUBS 0.02035f
C129 B.n95 VSUBS 0.008488f
C130 B.n96 VSUBS 0.008488f
C131 B.n97 VSUBS 0.008488f
C132 B.n98 VSUBS 0.008488f
C133 B.n99 VSUBS 0.008488f
C134 B.n100 VSUBS 0.008488f
C135 B.n101 VSUBS 0.008488f
C136 B.n102 VSUBS 0.008488f
C137 B.n103 VSUBS 0.008488f
C138 B.n104 VSUBS 0.008488f
C139 B.n105 VSUBS 0.008488f
C140 B.n106 VSUBS 0.008488f
C141 B.n107 VSUBS 0.008488f
C142 B.n108 VSUBS 0.008488f
C143 B.n109 VSUBS 0.008488f
C144 B.n110 VSUBS 0.008488f
C145 B.n111 VSUBS 0.008488f
C146 B.n112 VSUBS 0.008488f
C147 B.n113 VSUBS 0.008488f
C148 B.n114 VSUBS 0.008488f
C149 B.n115 VSUBS 0.008488f
C150 B.n116 VSUBS 0.008488f
C151 B.n117 VSUBS 0.008488f
C152 B.n118 VSUBS 0.008488f
C153 B.n119 VSUBS 0.008488f
C154 B.n120 VSUBS 0.008488f
C155 B.n121 VSUBS 0.008488f
C156 B.n122 VSUBS 0.008488f
C157 B.n123 VSUBS 0.008488f
C158 B.n124 VSUBS 0.008488f
C159 B.n125 VSUBS 0.008488f
C160 B.n126 VSUBS 0.008488f
C161 B.n127 VSUBS 0.008488f
C162 B.n128 VSUBS 0.008488f
C163 B.n129 VSUBS 0.008488f
C164 B.n130 VSUBS 0.008488f
C165 B.n131 VSUBS 0.008488f
C166 B.n132 VSUBS 0.008488f
C167 B.n133 VSUBS 0.008488f
C168 B.n134 VSUBS 0.008488f
C169 B.n135 VSUBS 0.008488f
C170 B.n136 VSUBS 0.008488f
C171 B.n137 VSUBS 0.008488f
C172 B.n138 VSUBS 0.008488f
C173 B.n139 VSUBS 0.008488f
C174 B.n140 VSUBS 0.008488f
C175 B.n141 VSUBS 0.008488f
C176 B.n142 VSUBS 0.008488f
C177 B.n143 VSUBS 0.008488f
C178 B.n144 VSUBS 0.008488f
C179 B.n145 VSUBS 0.008488f
C180 B.n146 VSUBS 0.008488f
C181 B.n147 VSUBS 0.008488f
C182 B.n148 VSUBS 0.008488f
C183 B.n149 VSUBS 0.008488f
C184 B.n150 VSUBS 0.008488f
C185 B.n151 VSUBS 0.008488f
C186 B.n152 VSUBS 0.008488f
C187 B.n153 VSUBS 0.008488f
C188 B.n154 VSUBS 0.008488f
C189 B.n155 VSUBS 0.008488f
C190 B.n156 VSUBS 0.008488f
C191 B.n157 VSUBS 0.008488f
C192 B.n158 VSUBS 0.008488f
C193 B.n159 VSUBS 0.008488f
C194 B.n160 VSUBS 0.008488f
C195 B.n161 VSUBS 0.008488f
C196 B.n162 VSUBS 0.008488f
C197 B.n163 VSUBS 0.008488f
C198 B.n164 VSUBS 0.008488f
C199 B.n165 VSUBS 0.021275f
C200 B.n166 VSUBS 0.008488f
C201 B.n167 VSUBS 0.008488f
C202 B.n168 VSUBS 0.008488f
C203 B.n169 VSUBS 0.008488f
C204 B.n170 VSUBS 0.008488f
C205 B.n171 VSUBS 0.008488f
C206 B.n172 VSUBS 0.008488f
C207 B.n173 VSUBS 0.008488f
C208 B.n174 VSUBS 0.008488f
C209 B.n175 VSUBS 0.008488f
C210 B.n176 VSUBS 0.008488f
C211 B.n177 VSUBS 0.008488f
C212 B.n178 VSUBS 0.008488f
C213 B.n179 VSUBS 0.008488f
C214 B.n180 VSUBS 0.008488f
C215 B.n181 VSUBS 0.008488f
C216 B.n182 VSUBS 0.008488f
C217 B.n183 VSUBS 0.008488f
C218 B.n184 VSUBS 0.008488f
C219 B.n185 VSUBS 0.008488f
C220 B.n186 VSUBS 0.008488f
C221 B.n187 VSUBS 0.008488f
C222 B.n188 VSUBS 0.008488f
C223 B.n189 VSUBS 0.008488f
C224 B.t7 VSUBS 0.575677f
C225 B.t8 VSUBS 0.605964f
C226 B.t6 VSUBS 2.52169f
C227 B.n190 VSUBS 0.340775f
C228 B.n191 VSUBS 0.090197f
C229 B.n192 VSUBS 0.008488f
C230 B.n193 VSUBS 0.008488f
C231 B.n194 VSUBS 0.008488f
C232 B.n195 VSUBS 0.008488f
C233 B.t1 VSUBS 0.575692f
C234 B.t2 VSUBS 0.605977f
C235 B.t0 VSUBS 2.52169f
C236 B.n196 VSUBS 0.340763f
C237 B.n197 VSUBS 0.090181f
C238 B.n198 VSUBS 0.019666f
C239 B.n199 VSUBS 0.008488f
C240 B.n200 VSUBS 0.008488f
C241 B.n201 VSUBS 0.008488f
C242 B.n202 VSUBS 0.008488f
C243 B.n203 VSUBS 0.008488f
C244 B.n204 VSUBS 0.008488f
C245 B.n205 VSUBS 0.008488f
C246 B.n206 VSUBS 0.008488f
C247 B.n207 VSUBS 0.008488f
C248 B.n208 VSUBS 0.008488f
C249 B.n209 VSUBS 0.008488f
C250 B.n210 VSUBS 0.008488f
C251 B.n211 VSUBS 0.008488f
C252 B.n212 VSUBS 0.008488f
C253 B.n213 VSUBS 0.008488f
C254 B.n214 VSUBS 0.008488f
C255 B.n215 VSUBS 0.008488f
C256 B.n216 VSUBS 0.008488f
C257 B.n217 VSUBS 0.008488f
C258 B.n218 VSUBS 0.008488f
C259 B.n219 VSUBS 0.008488f
C260 B.n220 VSUBS 0.008488f
C261 B.n221 VSUBS 0.008488f
C262 B.n222 VSUBS 0.021275f
C263 B.n223 VSUBS 0.008488f
C264 B.n224 VSUBS 0.008488f
C265 B.n225 VSUBS 0.008488f
C266 B.n226 VSUBS 0.008488f
C267 B.n227 VSUBS 0.008488f
C268 B.n228 VSUBS 0.008488f
C269 B.n229 VSUBS 0.008488f
C270 B.n230 VSUBS 0.008488f
C271 B.n231 VSUBS 0.008488f
C272 B.n232 VSUBS 0.008488f
C273 B.n233 VSUBS 0.008488f
C274 B.n234 VSUBS 0.008488f
C275 B.n235 VSUBS 0.008488f
C276 B.n236 VSUBS 0.008488f
C277 B.n237 VSUBS 0.008488f
C278 B.n238 VSUBS 0.008488f
C279 B.n239 VSUBS 0.008488f
C280 B.n240 VSUBS 0.008488f
C281 B.n241 VSUBS 0.008488f
C282 B.n242 VSUBS 0.008488f
C283 B.n243 VSUBS 0.008488f
C284 B.n244 VSUBS 0.008488f
C285 B.n245 VSUBS 0.008488f
C286 B.n246 VSUBS 0.008488f
C287 B.n247 VSUBS 0.008488f
C288 B.n248 VSUBS 0.008488f
C289 B.n249 VSUBS 0.008488f
C290 B.n250 VSUBS 0.008488f
C291 B.n251 VSUBS 0.008488f
C292 B.n252 VSUBS 0.008488f
C293 B.n253 VSUBS 0.008488f
C294 B.n254 VSUBS 0.008488f
C295 B.n255 VSUBS 0.008488f
C296 B.n256 VSUBS 0.008488f
C297 B.n257 VSUBS 0.008488f
C298 B.n258 VSUBS 0.008488f
C299 B.n259 VSUBS 0.008488f
C300 B.n260 VSUBS 0.008488f
C301 B.n261 VSUBS 0.008488f
C302 B.n262 VSUBS 0.008488f
C303 B.n263 VSUBS 0.008488f
C304 B.n264 VSUBS 0.008488f
C305 B.n265 VSUBS 0.008488f
C306 B.n266 VSUBS 0.008488f
C307 B.n267 VSUBS 0.008488f
C308 B.n268 VSUBS 0.008488f
C309 B.n269 VSUBS 0.008488f
C310 B.n270 VSUBS 0.008488f
C311 B.n271 VSUBS 0.008488f
C312 B.n272 VSUBS 0.008488f
C313 B.n273 VSUBS 0.008488f
C314 B.n274 VSUBS 0.008488f
C315 B.n275 VSUBS 0.008488f
C316 B.n276 VSUBS 0.008488f
C317 B.n277 VSUBS 0.008488f
C318 B.n278 VSUBS 0.008488f
C319 B.n279 VSUBS 0.008488f
C320 B.n280 VSUBS 0.008488f
C321 B.n281 VSUBS 0.008488f
C322 B.n282 VSUBS 0.008488f
C323 B.n283 VSUBS 0.008488f
C324 B.n284 VSUBS 0.008488f
C325 B.n285 VSUBS 0.008488f
C326 B.n286 VSUBS 0.008488f
C327 B.n287 VSUBS 0.008488f
C328 B.n288 VSUBS 0.008488f
C329 B.n289 VSUBS 0.008488f
C330 B.n290 VSUBS 0.008488f
C331 B.n291 VSUBS 0.008488f
C332 B.n292 VSUBS 0.008488f
C333 B.n293 VSUBS 0.008488f
C334 B.n294 VSUBS 0.008488f
C335 B.n295 VSUBS 0.008488f
C336 B.n296 VSUBS 0.008488f
C337 B.n297 VSUBS 0.008488f
C338 B.n298 VSUBS 0.008488f
C339 B.n299 VSUBS 0.008488f
C340 B.n300 VSUBS 0.008488f
C341 B.n301 VSUBS 0.008488f
C342 B.n302 VSUBS 0.008488f
C343 B.n303 VSUBS 0.008488f
C344 B.n304 VSUBS 0.008488f
C345 B.n305 VSUBS 0.008488f
C346 B.n306 VSUBS 0.008488f
C347 B.n307 VSUBS 0.008488f
C348 B.n308 VSUBS 0.008488f
C349 B.n309 VSUBS 0.008488f
C350 B.n310 VSUBS 0.008488f
C351 B.n311 VSUBS 0.008488f
C352 B.n312 VSUBS 0.008488f
C353 B.n313 VSUBS 0.008488f
C354 B.n314 VSUBS 0.008488f
C355 B.n315 VSUBS 0.008488f
C356 B.n316 VSUBS 0.008488f
C357 B.n317 VSUBS 0.008488f
C358 B.n318 VSUBS 0.008488f
C359 B.n319 VSUBS 0.008488f
C360 B.n320 VSUBS 0.008488f
C361 B.n321 VSUBS 0.008488f
C362 B.n322 VSUBS 0.008488f
C363 B.n323 VSUBS 0.008488f
C364 B.n324 VSUBS 0.008488f
C365 B.n325 VSUBS 0.008488f
C366 B.n326 VSUBS 0.008488f
C367 B.n327 VSUBS 0.008488f
C368 B.n328 VSUBS 0.008488f
C369 B.n329 VSUBS 0.008488f
C370 B.n330 VSUBS 0.008488f
C371 B.n331 VSUBS 0.008488f
C372 B.n332 VSUBS 0.008488f
C373 B.n333 VSUBS 0.008488f
C374 B.n334 VSUBS 0.008488f
C375 B.n335 VSUBS 0.008488f
C376 B.n336 VSUBS 0.008488f
C377 B.n337 VSUBS 0.008488f
C378 B.n338 VSUBS 0.008488f
C379 B.n339 VSUBS 0.008488f
C380 B.n340 VSUBS 0.008488f
C381 B.n341 VSUBS 0.008488f
C382 B.n342 VSUBS 0.008488f
C383 B.n343 VSUBS 0.008488f
C384 B.n344 VSUBS 0.008488f
C385 B.n345 VSUBS 0.008488f
C386 B.n346 VSUBS 0.008488f
C387 B.n347 VSUBS 0.008488f
C388 B.n348 VSUBS 0.008488f
C389 B.n349 VSUBS 0.008488f
C390 B.n350 VSUBS 0.008488f
C391 B.n351 VSUBS 0.008488f
C392 B.n352 VSUBS 0.008488f
C393 B.n353 VSUBS 0.008488f
C394 B.n354 VSUBS 0.008488f
C395 B.n355 VSUBS 0.008488f
C396 B.n356 VSUBS 0.008488f
C397 B.n357 VSUBS 0.008488f
C398 B.n358 VSUBS 0.008488f
C399 B.n359 VSUBS 0.020666f
C400 B.n360 VSUBS 0.020666f
C401 B.n361 VSUBS 0.021275f
C402 B.n362 VSUBS 0.008488f
C403 B.n363 VSUBS 0.008488f
C404 B.n364 VSUBS 0.008488f
C405 B.n365 VSUBS 0.008488f
C406 B.n366 VSUBS 0.008488f
C407 B.n367 VSUBS 0.008488f
C408 B.n368 VSUBS 0.008488f
C409 B.n369 VSUBS 0.008488f
C410 B.n370 VSUBS 0.008488f
C411 B.n371 VSUBS 0.008488f
C412 B.n372 VSUBS 0.008488f
C413 B.n373 VSUBS 0.008488f
C414 B.n374 VSUBS 0.008488f
C415 B.n375 VSUBS 0.008488f
C416 B.n376 VSUBS 0.008488f
C417 B.n377 VSUBS 0.008488f
C418 B.n378 VSUBS 0.008488f
C419 B.n379 VSUBS 0.008488f
C420 B.n380 VSUBS 0.008488f
C421 B.n381 VSUBS 0.008488f
C422 B.n382 VSUBS 0.008488f
C423 B.n383 VSUBS 0.008488f
C424 B.n384 VSUBS 0.008488f
C425 B.n385 VSUBS 0.008488f
C426 B.n386 VSUBS 0.008488f
C427 B.n387 VSUBS 0.008488f
C428 B.n388 VSUBS 0.008488f
C429 B.n389 VSUBS 0.008488f
C430 B.n390 VSUBS 0.008488f
C431 B.n391 VSUBS 0.008488f
C432 B.n392 VSUBS 0.008488f
C433 B.n393 VSUBS 0.008488f
C434 B.n394 VSUBS 0.008488f
C435 B.n395 VSUBS 0.008488f
C436 B.n396 VSUBS 0.008488f
C437 B.n397 VSUBS 0.008488f
C438 B.n398 VSUBS 0.008488f
C439 B.n399 VSUBS 0.008488f
C440 B.n400 VSUBS 0.008488f
C441 B.n401 VSUBS 0.008488f
C442 B.n402 VSUBS 0.008488f
C443 B.n403 VSUBS 0.008488f
C444 B.n404 VSUBS 0.008488f
C445 B.n405 VSUBS 0.008488f
C446 B.n406 VSUBS 0.008488f
C447 B.n407 VSUBS 0.008488f
C448 B.n408 VSUBS 0.008488f
C449 B.n409 VSUBS 0.008488f
C450 B.n410 VSUBS 0.008488f
C451 B.n411 VSUBS 0.008488f
C452 B.n412 VSUBS 0.008488f
C453 B.n413 VSUBS 0.008488f
C454 B.n414 VSUBS 0.008488f
C455 B.n415 VSUBS 0.008488f
C456 B.n416 VSUBS 0.008488f
C457 B.n417 VSUBS 0.008488f
C458 B.n418 VSUBS 0.008488f
C459 B.n419 VSUBS 0.008488f
C460 B.n420 VSUBS 0.008488f
C461 B.n421 VSUBS 0.008488f
C462 B.n422 VSUBS 0.008488f
C463 B.n423 VSUBS 0.008488f
C464 B.n424 VSUBS 0.008488f
C465 B.n425 VSUBS 0.008488f
C466 B.n426 VSUBS 0.008488f
C467 B.n427 VSUBS 0.008488f
C468 B.n428 VSUBS 0.008488f
C469 B.n429 VSUBS 0.008488f
C470 B.n430 VSUBS 0.008488f
C471 B.n431 VSUBS 0.007989f
C472 B.n432 VSUBS 0.008488f
C473 B.n433 VSUBS 0.008488f
C474 B.n434 VSUBS 0.004743f
C475 B.n435 VSUBS 0.008488f
C476 B.n436 VSUBS 0.008488f
C477 B.n437 VSUBS 0.008488f
C478 B.n438 VSUBS 0.008488f
C479 B.n439 VSUBS 0.008488f
C480 B.n440 VSUBS 0.008488f
C481 B.n441 VSUBS 0.008488f
C482 B.n442 VSUBS 0.008488f
C483 B.n443 VSUBS 0.008488f
C484 B.n444 VSUBS 0.008488f
C485 B.n445 VSUBS 0.008488f
C486 B.n446 VSUBS 0.008488f
C487 B.n447 VSUBS 0.004743f
C488 B.n448 VSUBS 0.019666f
C489 B.n449 VSUBS 0.007989f
C490 B.n450 VSUBS 0.008488f
C491 B.n451 VSUBS 0.008488f
C492 B.n452 VSUBS 0.008488f
C493 B.n453 VSUBS 0.008488f
C494 B.n454 VSUBS 0.008488f
C495 B.n455 VSUBS 0.008488f
C496 B.n456 VSUBS 0.008488f
C497 B.n457 VSUBS 0.008488f
C498 B.n458 VSUBS 0.008488f
C499 B.n459 VSUBS 0.008488f
C500 B.n460 VSUBS 0.008488f
C501 B.n461 VSUBS 0.008488f
C502 B.n462 VSUBS 0.008488f
C503 B.n463 VSUBS 0.008488f
C504 B.n464 VSUBS 0.008488f
C505 B.n465 VSUBS 0.008488f
C506 B.n466 VSUBS 0.008488f
C507 B.n467 VSUBS 0.008488f
C508 B.n468 VSUBS 0.008488f
C509 B.n469 VSUBS 0.008488f
C510 B.n470 VSUBS 0.008488f
C511 B.n471 VSUBS 0.008488f
C512 B.n472 VSUBS 0.008488f
C513 B.n473 VSUBS 0.008488f
C514 B.n474 VSUBS 0.008488f
C515 B.n475 VSUBS 0.008488f
C516 B.n476 VSUBS 0.008488f
C517 B.n477 VSUBS 0.008488f
C518 B.n478 VSUBS 0.008488f
C519 B.n479 VSUBS 0.008488f
C520 B.n480 VSUBS 0.008488f
C521 B.n481 VSUBS 0.008488f
C522 B.n482 VSUBS 0.008488f
C523 B.n483 VSUBS 0.008488f
C524 B.n484 VSUBS 0.008488f
C525 B.n485 VSUBS 0.008488f
C526 B.n486 VSUBS 0.008488f
C527 B.n487 VSUBS 0.008488f
C528 B.n488 VSUBS 0.008488f
C529 B.n489 VSUBS 0.008488f
C530 B.n490 VSUBS 0.008488f
C531 B.n491 VSUBS 0.008488f
C532 B.n492 VSUBS 0.008488f
C533 B.n493 VSUBS 0.008488f
C534 B.n494 VSUBS 0.008488f
C535 B.n495 VSUBS 0.008488f
C536 B.n496 VSUBS 0.008488f
C537 B.n497 VSUBS 0.008488f
C538 B.n498 VSUBS 0.008488f
C539 B.n499 VSUBS 0.008488f
C540 B.n500 VSUBS 0.008488f
C541 B.n501 VSUBS 0.008488f
C542 B.n502 VSUBS 0.008488f
C543 B.n503 VSUBS 0.008488f
C544 B.n504 VSUBS 0.008488f
C545 B.n505 VSUBS 0.008488f
C546 B.n506 VSUBS 0.008488f
C547 B.n507 VSUBS 0.008488f
C548 B.n508 VSUBS 0.008488f
C549 B.n509 VSUBS 0.008488f
C550 B.n510 VSUBS 0.008488f
C551 B.n511 VSUBS 0.008488f
C552 B.n512 VSUBS 0.008488f
C553 B.n513 VSUBS 0.008488f
C554 B.n514 VSUBS 0.008488f
C555 B.n515 VSUBS 0.008488f
C556 B.n516 VSUBS 0.008488f
C557 B.n517 VSUBS 0.008488f
C558 B.n518 VSUBS 0.008488f
C559 B.n519 VSUBS 0.008488f
C560 B.n520 VSUBS 0.021275f
C561 B.n521 VSUBS 0.020666f
C562 B.n522 VSUBS 0.020666f
C563 B.n523 VSUBS 0.008488f
C564 B.n524 VSUBS 0.008488f
C565 B.n525 VSUBS 0.008488f
C566 B.n526 VSUBS 0.008488f
C567 B.n527 VSUBS 0.008488f
C568 B.n528 VSUBS 0.008488f
C569 B.n529 VSUBS 0.008488f
C570 B.n530 VSUBS 0.008488f
C571 B.n531 VSUBS 0.008488f
C572 B.n532 VSUBS 0.008488f
C573 B.n533 VSUBS 0.008488f
C574 B.n534 VSUBS 0.008488f
C575 B.n535 VSUBS 0.008488f
C576 B.n536 VSUBS 0.008488f
C577 B.n537 VSUBS 0.008488f
C578 B.n538 VSUBS 0.008488f
C579 B.n539 VSUBS 0.008488f
C580 B.n540 VSUBS 0.008488f
C581 B.n541 VSUBS 0.008488f
C582 B.n542 VSUBS 0.008488f
C583 B.n543 VSUBS 0.008488f
C584 B.n544 VSUBS 0.008488f
C585 B.n545 VSUBS 0.008488f
C586 B.n546 VSUBS 0.008488f
C587 B.n547 VSUBS 0.008488f
C588 B.n548 VSUBS 0.008488f
C589 B.n549 VSUBS 0.008488f
C590 B.n550 VSUBS 0.008488f
C591 B.n551 VSUBS 0.008488f
C592 B.n552 VSUBS 0.008488f
C593 B.n553 VSUBS 0.008488f
C594 B.n554 VSUBS 0.008488f
C595 B.n555 VSUBS 0.008488f
C596 B.n556 VSUBS 0.008488f
C597 B.n557 VSUBS 0.008488f
C598 B.n558 VSUBS 0.008488f
C599 B.n559 VSUBS 0.008488f
C600 B.n560 VSUBS 0.008488f
C601 B.n561 VSUBS 0.008488f
C602 B.n562 VSUBS 0.008488f
C603 B.n563 VSUBS 0.008488f
C604 B.n564 VSUBS 0.008488f
C605 B.n565 VSUBS 0.008488f
C606 B.n566 VSUBS 0.008488f
C607 B.n567 VSUBS 0.008488f
C608 B.n568 VSUBS 0.008488f
C609 B.n569 VSUBS 0.008488f
C610 B.n570 VSUBS 0.008488f
C611 B.n571 VSUBS 0.008488f
C612 B.n572 VSUBS 0.008488f
C613 B.n573 VSUBS 0.008488f
C614 B.n574 VSUBS 0.008488f
C615 B.n575 VSUBS 0.008488f
C616 B.n576 VSUBS 0.008488f
C617 B.n577 VSUBS 0.008488f
C618 B.n578 VSUBS 0.008488f
C619 B.n579 VSUBS 0.008488f
C620 B.n580 VSUBS 0.008488f
C621 B.n581 VSUBS 0.008488f
C622 B.n582 VSUBS 0.008488f
C623 B.n583 VSUBS 0.008488f
C624 B.n584 VSUBS 0.008488f
C625 B.n585 VSUBS 0.008488f
C626 B.n586 VSUBS 0.008488f
C627 B.n587 VSUBS 0.008488f
C628 B.n588 VSUBS 0.008488f
C629 B.n589 VSUBS 0.008488f
C630 B.n590 VSUBS 0.008488f
C631 B.n591 VSUBS 0.008488f
C632 B.n592 VSUBS 0.008488f
C633 B.n593 VSUBS 0.008488f
C634 B.n594 VSUBS 0.008488f
C635 B.n595 VSUBS 0.008488f
C636 B.n596 VSUBS 0.008488f
C637 B.n597 VSUBS 0.008488f
C638 B.n598 VSUBS 0.008488f
C639 B.n599 VSUBS 0.008488f
C640 B.n600 VSUBS 0.008488f
C641 B.n601 VSUBS 0.008488f
C642 B.n602 VSUBS 0.008488f
C643 B.n603 VSUBS 0.008488f
C644 B.n604 VSUBS 0.008488f
C645 B.n605 VSUBS 0.008488f
C646 B.n606 VSUBS 0.008488f
C647 B.n607 VSUBS 0.008488f
C648 B.n608 VSUBS 0.008488f
C649 B.n609 VSUBS 0.008488f
C650 B.n610 VSUBS 0.008488f
C651 B.n611 VSUBS 0.008488f
C652 B.n612 VSUBS 0.008488f
C653 B.n613 VSUBS 0.008488f
C654 B.n614 VSUBS 0.008488f
C655 B.n615 VSUBS 0.008488f
C656 B.n616 VSUBS 0.008488f
C657 B.n617 VSUBS 0.008488f
C658 B.n618 VSUBS 0.008488f
C659 B.n619 VSUBS 0.008488f
C660 B.n620 VSUBS 0.008488f
C661 B.n621 VSUBS 0.008488f
C662 B.n622 VSUBS 0.008488f
C663 B.n623 VSUBS 0.008488f
C664 B.n624 VSUBS 0.008488f
C665 B.n625 VSUBS 0.008488f
C666 B.n626 VSUBS 0.008488f
C667 B.n627 VSUBS 0.008488f
C668 B.n628 VSUBS 0.008488f
C669 B.n629 VSUBS 0.008488f
C670 B.n630 VSUBS 0.008488f
C671 B.n631 VSUBS 0.008488f
C672 B.n632 VSUBS 0.008488f
C673 B.n633 VSUBS 0.008488f
C674 B.n634 VSUBS 0.008488f
C675 B.n635 VSUBS 0.008488f
C676 B.n636 VSUBS 0.008488f
C677 B.n637 VSUBS 0.008488f
C678 B.n638 VSUBS 0.008488f
C679 B.n639 VSUBS 0.008488f
C680 B.n640 VSUBS 0.008488f
C681 B.n641 VSUBS 0.008488f
C682 B.n642 VSUBS 0.008488f
C683 B.n643 VSUBS 0.008488f
C684 B.n644 VSUBS 0.008488f
C685 B.n645 VSUBS 0.008488f
C686 B.n646 VSUBS 0.008488f
C687 B.n647 VSUBS 0.008488f
C688 B.n648 VSUBS 0.008488f
C689 B.n649 VSUBS 0.008488f
C690 B.n650 VSUBS 0.008488f
C691 B.n651 VSUBS 0.008488f
C692 B.n652 VSUBS 0.008488f
C693 B.n653 VSUBS 0.008488f
C694 B.n654 VSUBS 0.008488f
C695 B.n655 VSUBS 0.008488f
C696 B.n656 VSUBS 0.008488f
C697 B.n657 VSUBS 0.008488f
C698 B.n658 VSUBS 0.008488f
C699 B.n659 VSUBS 0.008488f
C700 B.n660 VSUBS 0.008488f
C701 B.n661 VSUBS 0.008488f
C702 B.n662 VSUBS 0.008488f
C703 B.n663 VSUBS 0.008488f
C704 B.n664 VSUBS 0.008488f
C705 B.n665 VSUBS 0.008488f
C706 B.n666 VSUBS 0.008488f
C707 B.n667 VSUBS 0.008488f
C708 B.n668 VSUBS 0.008488f
C709 B.n669 VSUBS 0.008488f
C710 B.n670 VSUBS 0.008488f
C711 B.n671 VSUBS 0.008488f
C712 B.n672 VSUBS 0.008488f
C713 B.n673 VSUBS 0.008488f
C714 B.n674 VSUBS 0.008488f
C715 B.n675 VSUBS 0.008488f
C716 B.n676 VSUBS 0.008488f
C717 B.n677 VSUBS 0.008488f
C718 B.n678 VSUBS 0.008488f
C719 B.n679 VSUBS 0.008488f
C720 B.n680 VSUBS 0.008488f
C721 B.n681 VSUBS 0.008488f
C722 B.n682 VSUBS 0.008488f
C723 B.n683 VSUBS 0.008488f
C724 B.n684 VSUBS 0.008488f
C725 B.n685 VSUBS 0.008488f
C726 B.n686 VSUBS 0.008488f
C727 B.n687 VSUBS 0.008488f
C728 B.n688 VSUBS 0.008488f
C729 B.n689 VSUBS 0.008488f
C730 B.n690 VSUBS 0.008488f
C731 B.n691 VSUBS 0.008488f
C732 B.n692 VSUBS 0.008488f
C733 B.n693 VSUBS 0.008488f
C734 B.n694 VSUBS 0.008488f
C735 B.n695 VSUBS 0.008488f
C736 B.n696 VSUBS 0.008488f
C737 B.n697 VSUBS 0.008488f
C738 B.n698 VSUBS 0.008488f
C739 B.n699 VSUBS 0.008488f
C740 B.n700 VSUBS 0.008488f
C741 B.n701 VSUBS 0.008488f
C742 B.n702 VSUBS 0.008488f
C743 B.n703 VSUBS 0.008488f
C744 B.n704 VSUBS 0.008488f
C745 B.n705 VSUBS 0.008488f
C746 B.n706 VSUBS 0.008488f
C747 B.n707 VSUBS 0.008488f
C748 B.n708 VSUBS 0.008488f
C749 B.n709 VSUBS 0.008488f
C750 B.n710 VSUBS 0.008488f
C751 B.n711 VSUBS 0.008488f
C752 B.n712 VSUBS 0.008488f
C753 B.n713 VSUBS 0.008488f
C754 B.n714 VSUBS 0.008488f
C755 B.n715 VSUBS 0.008488f
C756 B.n716 VSUBS 0.008488f
C757 B.n717 VSUBS 0.008488f
C758 B.n718 VSUBS 0.008488f
C759 B.n719 VSUBS 0.008488f
C760 B.n720 VSUBS 0.008488f
C761 B.n721 VSUBS 0.008488f
C762 B.n722 VSUBS 0.008488f
C763 B.n723 VSUBS 0.008488f
C764 B.n724 VSUBS 0.008488f
C765 B.n725 VSUBS 0.008488f
C766 B.n726 VSUBS 0.008488f
C767 B.n727 VSUBS 0.008488f
C768 B.n728 VSUBS 0.008488f
C769 B.n729 VSUBS 0.008488f
C770 B.n730 VSUBS 0.008488f
C771 B.n731 VSUBS 0.02159f
C772 B.n732 VSUBS 0.020666f
C773 B.n733 VSUBS 0.021275f
C774 B.n734 VSUBS 0.008488f
C775 B.n735 VSUBS 0.008488f
C776 B.n736 VSUBS 0.008488f
C777 B.n737 VSUBS 0.008488f
C778 B.n738 VSUBS 0.008488f
C779 B.n739 VSUBS 0.008488f
C780 B.n740 VSUBS 0.008488f
C781 B.n741 VSUBS 0.008488f
C782 B.n742 VSUBS 0.008488f
C783 B.n743 VSUBS 0.008488f
C784 B.n744 VSUBS 0.008488f
C785 B.n745 VSUBS 0.008488f
C786 B.n746 VSUBS 0.008488f
C787 B.n747 VSUBS 0.008488f
C788 B.n748 VSUBS 0.008488f
C789 B.n749 VSUBS 0.008488f
C790 B.n750 VSUBS 0.008488f
C791 B.n751 VSUBS 0.008488f
C792 B.n752 VSUBS 0.008488f
C793 B.n753 VSUBS 0.008488f
C794 B.n754 VSUBS 0.008488f
C795 B.n755 VSUBS 0.008488f
C796 B.n756 VSUBS 0.008488f
C797 B.n757 VSUBS 0.008488f
C798 B.n758 VSUBS 0.008488f
C799 B.n759 VSUBS 0.008488f
C800 B.n760 VSUBS 0.008488f
C801 B.n761 VSUBS 0.008488f
C802 B.n762 VSUBS 0.008488f
C803 B.n763 VSUBS 0.008488f
C804 B.n764 VSUBS 0.008488f
C805 B.n765 VSUBS 0.008488f
C806 B.n766 VSUBS 0.008488f
C807 B.n767 VSUBS 0.008488f
C808 B.n768 VSUBS 0.008488f
C809 B.n769 VSUBS 0.008488f
C810 B.n770 VSUBS 0.008488f
C811 B.n771 VSUBS 0.008488f
C812 B.n772 VSUBS 0.008488f
C813 B.n773 VSUBS 0.008488f
C814 B.n774 VSUBS 0.008488f
C815 B.n775 VSUBS 0.008488f
C816 B.n776 VSUBS 0.008488f
C817 B.n777 VSUBS 0.008488f
C818 B.n778 VSUBS 0.008488f
C819 B.n779 VSUBS 0.008488f
C820 B.n780 VSUBS 0.008488f
C821 B.n781 VSUBS 0.008488f
C822 B.n782 VSUBS 0.008488f
C823 B.n783 VSUBS 0.008488f
C824 B.n784 VSUBS 0.008488f
C825 B.n785 VSUBS 0.008488f
C826 B.n786 VSUBS 0.008488f
C827 B.n787 VSUBS 0.008488f
C828 B.n788 VSUBS 0.008488f
C829 B.n789 VSUBS 0.008488f
C830 B.n790 VSUBS 0.008488f
C831 B.n791 VSUBS 0.008488f
C832 B.n792 VSUBS 0.008488f
C833 B.n793 VSUBS 0.008488f
C834 B.n794 VSUBS 0.008488f
C835 B.n795 VSUBS 0.008488f
C836 B.n796 VSUBS 0.008488f
C837 B.n797 VSUBS 0.008488f
C838 B.n798 VSUBS 0.008488f
C839 B.n799 VSUBS 0.008488f
C840 B.n800 VSUBS 0.008488f
C841 B.n801 VSUBS 0.008488f
C842 B.n802 VSUBS 0.008488f
C843 B.n803 VSUBS 0.007989f
C844 B.n804 VSUBS 0.008488f
C845 B.n805 VSUBS 0.008488f
C846 B.n806 VSUBS 0.004743f
C847 B.n807 VSUBS 0.008488f
C848 B.n808 VSUBS 0.008488f
C849 B.n809 VSUBS 0.008488f
C850 B.n810 VSUBS 0.008488f
C851 B.n811 VSUBS 0.008488f
C852 B.n812 VSUBS 0.008488f
C853 B.n813 VSUBS 0.008488f
C854 B.n814 VSUBS 0.008488f
C855 B.n815 VSUBS 0.008488f
C856 B.n816 VSUBS 0.008488f
C857 B.n817 VSUBS 0.008488f
C858 B.n818 VSUBS 0.008488f
C859 B.n819 VSUBS 0.004743f
C860 B.n820 VSUBS 0.019666f
C861 B.n821 VSUBS 0.007989f
C862 B.n822 VSUBS 0.008488f
C863 B.n823 VSUBS 0.008488f
C864 B.n824 VSUBS 0.008488f
C865 B.n825 VSUBS 0.008488f
C866 B.n826 VSUBS 0.008488f
C867 B.n827 VSUBS 0.008488f
C868 B.n828 VSUBS 0.008488f
C869 B.n829 VSUBS 0.008488f
C870 B.n830 VSUBS 0.008488f
C871 B.n831 VSUBS 0.008488f
C872 B.n832 VSUBS 0.008488f
C873 B.n833 VSUBS 0.008488f
C874 B.n834 VSUBS 0.008488f
C875 B.n835 VSUBS 0.008488f
C876 B.n836 VSUBS 0.008488f
C877 B.n837 VSUBS 0.008488f
C878 B.n838 VSUBS 0.008488f
C879 B.n839 VSUBS 0.008488f
C880 B.n840 VSUBS 0.008488f
C881 B.n841 VSUBS 0.008488f
C882 B.n842 VSUBS 0.008488f
C883 B.n843 VSUBS 0.008488f
C884 B.n844 VSUBS 0.008488f
C885 B.n845 VSUBS 0.008488f
C886 B.n846 VSUBS 0.008488f
C887 B.n847 VSUBS 0.008488f
C888 B.n848 VSUBS 0.008488f
C889 B.n849 VSUBS 0.008488f
C890 B.n850 VSUBS 0.008488f
C891 B.n851 VSUBS 0.008488f
C892 B.n852 VSUBS 0.008488f
C893 B.n853 VSUBS 0.008488f
C894 B.n854 VSUBS 0.008488f
C895 B.n855 VSUBS 0.008488f
C896 B.n856 VSUBS 0.008488f
C897 B.n857 VSUBS 0.008488f
C898 B.n858 VSUBS 0.008488f
C899 B.n859 VSUBS 0.008488f
C900 B.n860 VSUBS 0.008488f
C901 B.n861 VSUBS 0.008488f
C902 B.n862 VSUBS 0.008488f
C903 B.n863 VSUBS 0.008488f
C904 B.n864 VSUBS 0.008488f
C905 B.n865 VSUBS 0.008488f
C906 B.n866 VSUBS 0.008488f
C907 B.n867 VSUBS 0.008488f
C908 B.n868 VSUBS 0.008488f
C909 B.n869 VSUBS 0.008488f
C910 B.n870 VSUBS 0.008488f
C911 B.n871 VSUBS 0.008488f
C912 B.n872 VSUBS 0.008488f
C913 B.n873 VSUBS 0.008488f
C914 B.n874 VSUBS 0.008488f
C915 B.n875 VSUBS 0.008488f
C916 B.n876 VSUBS 0.008488f
C917 B.n877 VSUBS 0.008488f
C918 B.n878 VSUBS 0.008488f
C919 B.n879 VSUBS 0.008488f
C920 B.n880 VSUBS 0.008488f
C921 B.n881 VSUBS 0.008488f
C922 B.n882 VSUBS 0.008488f
C923 B.n883 VSUBS 0.008488f
C924 B.n884 VSUBS 0.008488f
C925 B.n885 VSUBS 0.008488f
C926 B.n886 VSUBS 0.008488f
C927 B.n887 VSUBS 0.008488f
C928 B.n888 VSUBS 0.008488f
C929 B.n889 VSUBS 0.008488f
C930 B.n890 VSUBS 0.008488f
C931 B.n891 VSUBS 0.008488f
C932 B.n892 VSUBS 0.021275f
C933 B.n893 VSUBS 0.020666f
C934 B.n894 VSUBS 0.020666f
C935 B.n895 VSUBS 0.008488f
C936 B.n896 VSUBS 0.008488f
C937 B.n897 VSUBS 0.008488f
C938 B.n898 VSUBS 0.008488f
C939 B.n899 VSUBS 0.008488f
C940 B.n900 VSUBS 0.008488f
C941 B.n901 VSUBS 0.008488f
C942 B.n902 VSUBS 0.008488f
C943 B.n903 VSUBS 0.008488f
C944 B.n904 VSUBS 0.008488f
C945 B.n905 VSUBS 0.008488f
C946 B.n906 VSUBS 0.008488f
C947 B.n907 VSUBS 0.008488f
C948 B.n908 VSUBS 0.008488f
C949 B.n909 VSUBS 0.008488f
C950 B.n910 VSUBS 0.008488f
C951 B.n911 VSUBS 0.008488f
C952 B.n912 VSUBS 0.008488f
C953 B.n913 VSUBS 0.008488f
C954 B.n914 VSUBS 0.008488f
C955 B.n915 VSUBS 0.008488f
C956 B.n916 VSUBS 0.008488f
C957 B.n917 VSUBS 0.008488f
C958 B.n918 VSUBS 0.008488f
C959 B.n919 VSUBS 0.008488f
C960 B.n920 VSUBS 0.008488f
C961 B.n921 VSUBS 0.008488f
C962 B.n922 VSUBS 0.008488f
C963 B.n923 VSUBS 0.008488f
C964 B.n924 VSUBS 0.008488f
C965 B.n925 VSUBS 0.008488f
C966 B.n926 VSUBS 0.008488f
C967 B.n927 VSUBS 0.008488f
C968 B.n928 VSUBS 0.008488f
C969 B.n929 VSUBS 0.008488f
C970 B.n930 VSUBS 0.008488f
C971 B.n931 VSUBS 0.008488f
C972 B.n932 VSUBS 0.008488f
C973 B.n933 VSUBS 0.008488f
C974 B.n934 VSUBS 0.008488f
C975 B.n935 VSUBS 0.008488f
C976 B.n936 VSUBS 0.008488f
C977 B.n937 VSUBS 0.008488f
C978 B.n938 VSUBS 0.008488f
C979 B.n939 VSUBS 0.008488f
C980 B.n940 VSUBS 0.008488f
C981 B.n941 VSUBS 0.008488f
C982 B.n942 VSUBS 0.008488f
C983 B.n943 VSUBS 0.008488f
C984 B.n944 VSUBS 0.008488f
C985 B.n945 VSUBS 0.008488f
C986 B.n946 VSUBS 0.008488f
C987 B.n947 VSUBS 0.008488f
C988 B.n948 VSUBS 0.008488f
C989 B.n949 VSUBS 0.008488f
C990 B.n950 VSUBS 0.008488f
C991 B.n951 VSUBS 0.008488f
C992 B.n952 VSUBS 0.008488f
C993 B.n953 VSUBS 0.008488f
C994 B.n954 VSUBS 0.008488f
C995 B.n955 VSUBS 0.008488f
C996 B.n956 VSUBS 0.008488f
C997 B.n957 VSUBS 0.008488f
C998 B.n958 VSUBS 0.008488f
C999 B.n959 VSUBS 0.008488f
C1000 B.n960 VSUBS 0.008488f
C1001 B.n961 VSUBS 0.008488f
C1002 B.n962 VSUBS 0.008488f
C1003 B.n963 VSUBS 0.008488f
C1004 B.n964 VSUBS 0.008488f
C1005 B.n965 VSUBS 0.008488f
C1006 B.n966 VSUBS 0.008488f
C1007 B.n967 VSUBS 0.008488f
C1008 B.n968 VSUBS 0.008488f
C1009 B.n969 VSUBS 0.008488f
C1010 B.n970 VSUBS 0.008488f
C1011 B.n971 VSUBS 0.008488f
C1012 B.n972 VSUBS 0.008488f
C1013 B.n973 VSUBS 0.008488f
C1014 B.n974 VSUBS 0.008488f
C1015 B.n975 VSUBS 0.008488f
C1016 B.n976 VSUBS 0.008488f
C1017 B.n977 VSUBS 0.008488f
C1018 B.n978 VSUBS 0.008488f
C1019 B.n979 VSUBS 0.008488f
C1020 B.n980 VSUBS 0.008488f
C1021 B.n981 VSUBS 0.008488f
C1022 B.n982 VSUBS 0.008488f
C1023 B.n983 VSUBS 0.008488f
C1024 B.n984 VSUBS 0.008488f
C1025 B.n985 VSUBS 0.008488f
C1026 B.n986 VSUBS 0.008488f
C1027 B.n987 VSUBS 0.008488f
C1028 B.n988 VSUBS 0.008488f
C1029 B.n989 VSUBS 0.008488f
C1030 B.n990 VSUBS 0.008488f
C1031 B.n991 VSUBS 0.008488f
C1032 B.n992 VSUBS 0.008488f
C1033 B.n993 VSUBS 0.008488f
C1034 B.n994 VSUBS 0.008488f
C1035 B.n995 VSUBS 0.008488f
C1036 B.n996 VSUBS 0.008488f
C1037 B.n997 VSUBS 0.008488f
C1038 B.n998 VSUBS 0.008488f
C1039 B.n999 VSUBS 0.01922f
C1040 VDD2.t4 VSUBS 3.55254f
C1041 VDD2.t9 VSUBS 0.334847f
C1042 VDD2.t2 VSUBS 0.334847f
C1043 VDD2.n0 VSUBS 2.70217f
C1044 VDD2.n1 VSUBS 1.8381f
C1045 VDD2.t6 VSUBS 0.334847f
C1046 VDD2.t0 VSUBS 0.334847f
C1047 VDD2.n2 VSUBS 2.7342f
C1048 VDD2.n3 VSUBS 4.27746f
C1049 VDD2.t5 VSUBS 3.51489f
C1050 VDD2.n4 VSUBS 4.5131f
C1051 VDD2.t7 VSUBS 0.334847f
C1052 VDD2.t8 VSUBS 0.334847f
C1053 VDD2.n5 VSUBS 2.70217f
C1054 VDD2.n6 VSUBS 0.925425f
C1055 VDD2.t1 VSUBS 0.334847f
C1056 VDD2.t3 VSUBS 0.334847f
C1057 VDD2.n7 VSUBS 2.73413f
C1058 VN.t9 VSUBS 2.99692f
C1059 VN.n0 VSUBS 1.13495f
C1060 VN.n1 VSUBS 0.024043f
C1061 VN.n2 VSUBS 0.019526f
C1062 VN.n3 VSUBS 0.024043f
C1063 VN.t3 VSUBS 2.99692f
C1064 VN.n4 VSUBS 1.04502f
C1065 VN.n5 VSUBS 0.024043f
C1066 VN.n6 VSUBS 0.019464f
C1067 VN.n7 VSUBS 0.024043f
C1068 VN.t7 VSUBS 2.99692f
C1069 VN.n8 VSUBS 1.04502f
C1070 VN.n9 VSUBS 0.024043f
C1071 VN.n10 VSUBS 0.019464f
C1072 VN.n11 VSUBS 0.024043f
C1073 VN.t0 VSUBS 2.99692f
C1074 VN.n12 VSUBS 1.12484f
C1075 VN.t5 VSUBS 3.27779f
C1076 VN.n13 VSUBS 1.07915f
C1077 VN.n14 VSUBS 0.279673f
C1078 VN.n15 VSUBS 0.034362f
C1079 VN.n16 VSUBS 0.045035f
C1080 VN.n17 VSUBS 0.047915f
C1081 VN.n18 VSUBS 0.024043f
C1082 VN.n19 VSUBS 0.024043f
C1083 VN.n20 VSUBS 0.024043f
C1084 VN.n21 VSUBS 0.048159f
C1085 VN.n22 VSUBS 0.045035f
C1086 VN.n23 VSUBS 0.033917f
C1087 VN.n24 VSUBS 0.024043f
C1088 VN.n25 VSUBS 0.024043f
C1089 VN.n26 VSUBS 0.033917f
C1090 VN.n27 VSUBS 0.045035f
C1091 VN.n28 VSUBS 0.048159f
C1092 VN.n29 VSUBS 0.024043f
C1093 VN.n30 VSUBS 0.024043f
C1094 VN.n31 VSUBS 0.024043f
C1095 VN.n32 VSUBS 0.047915f
C1096 VN.n33 VSUBS 0.045035f
C1097 VN.n34 VSUBS 0.034362f
C1098 VN.n35 VSUBS 0.024043f
C1099 VN.n36 VSUBS 0.024043f
C1100 VN.n37 VSUBS 0.033473f
C1101 VN.n38 VSUBS 0.045035f
C1102 VN.n39 VSUBS 0.04837f
C1103 VN.n40 VSUBS 0.024043f
C1104 VN.n41 VSUBS 0.024043f
C1105 VN.n42 VSUBS 0.024043f
C1106 VN.n43 VSUBS 0.047641f
C1107 VN.n44 VSUBS 0.045035f
C1108 VN.n45 VSUBS 0.034807f
C1109 VN.n46 VSUBS 0.038811f
C1110 VN.n47 VSUBS 0.058371f
C1111 VN.t4 VSUBS 2.99692f
C1112 VN.n48 VSUBS 1.13495f
C1113 VN.n49 VSUBS 0.024043f
C1114 VN.n50 VSUBS 0.019526f
C1115 VN.n51 VSUBS 0.024043f
C1116 VN.t2 VSUBS 2.99692f
C1117 VN.n52 VSUBS 1.04502f
C1118 VN.n53 VSUBS 0.024043f
C1119 VN.n54 VSUBS 0.019464f
C1120 VN.n55 VSUBS 0.024043f
C1121 VN.t1 VSUBS 2.99692f
C1122 VN.n56 VSUBS 1.04502f
C1123 VN.n57 VSUBS 0.024043f
C1124 VN.n58 VSUBS 0.019464f
C1125 VN.n59 VSUBS 0.024043f
C1126 VN.t8 VSUBS 2.99692f
C1127 VN.n60 VSUBS 1.12484f
C1128 VN.t6 VSUBS 3.27779f
C1129 VN.n61 VSUBS 1.07915f
C1130 VN.n62 VSUBS 0.279673f
C1131 VN.n63 VSUBS 0.034362f
C1132 VN.n64 VSUBS 0.045035f
C1133 VN.n65 VSUBS 0.047915f
C1134 VN.n66 VSUBS 0.024043f
C1135 VN.n67 VSUBS 0.024043f
C1136 VN.n68 VSUBS 0.024043f
C1137 VN.n69 VSUBS 0.048159f
C1138 VN.n70 VSUBS 0.045035f
C1139 VN.n71 VSUBS 0.033917f
C1140 VN.n72 VSUBS 0.024043f
C1141 VN.n73 VSUBS 0.024043f
C1142 VN.n74 VSUBS 0.033917f
C1143 VN.n75 VSUBS 0.045035f
C1144 VN.n76 VSUBS 0.048159f
C1145 VN.n77 VSUBS 0.024043f
C1146 VN.n78 VSUBS 0.024043f
C1147 VN.n79 VSUBS 0.024043f
C1148 VN.n80 VSUBS 0.047915f
C1149 VN.n81 VSUBS 0.045035f
C1150 VN.n82 VSUBS 0.034362f
C1151 VN.n83 VSUBS 0.024043f
C1152 VN.n84 VSUBS 0.024043f
C1153 VN.n85 VSUBS 0.033473f
C1154 VN.n86 VSUBS 0.045035f
C1155 VN.n87 VSUBS 0.04837f
C1156 VN.n88 VSUBS 0.024043f
C1157 VN.n89 VSUBS 0.024043f
C1158 VN.n90 VSUBS 0.024043f
C1159 VN.n91 VSUBS 0.047641f
C1160 VN.n92 VSUBS 0.045035f
C1161 VN.n93 VSUBS 0.034807f
C1162 VN.n94 VSUBS 0.038811f
C1163 VN.n95 VSUBS 1.69363f
C1164 VTAIL.t9 VSUBS 0.323971f
C1165 VTAIL.t1 VSUBS 0.323971f
C1166 VTAIL.n0 VSUBS 2.45238f
C1167 VTAIL.n1 VSUBS 1.06182f
C1168 VTAIL.t17 VSUBS 3.21683f
C1169 VTAIL.n2 VSUBS 1.24534f
C1170 VTAIL.t14 VSUBS 0.323971f
C1171 VTAIL.t11 VSUBS 0.323971f
C1172 VTAIL.n3 VSUBS 2.45238f
C1173 VTAIL.n4 VSUBS 1.22246f
C1174 VTAIL.t13 VSUBS 0.323971f
C1175 VTAIL.t18 VSUBS 0.323971f
C1176 VTAIL.n5 VSUBS 2.45238f
C1177 VTAIL.n6 VSUBS 3.0293f
C1178 VTAIL.t4 VSUBS 0.323971f
C1179 VTAIL.t6 VSUBS 0.323971f
C1180 VTAIL.n7 VSUBS 2.45238f
C1181 VTAIL.n8 VSUBS 3.02929f
C1182 VTAIL.t3 VSUBS 0.323971f
C1183 VTAIL.t8 VSUBS 0.323971f
C1184 VTAIL.n9 VSUBS 2.45238f
C1185 VTAIL.n10 VSUBS 1.22246f
C1186 VTAIL.t0 VSUBS 3.21686f
C1187 VTAIL.n11 VSUBS 1.24531f
C1188 VTAIL.t12 VSUBS 0.323971f
C1189 VTAIL.t19 VSUBS 0.323971f
C1190 VTAIL.n12 VSUBS 2.45238f
C1191 VTAIL.n13 VSUBS 1.12623f
C1192 VTAIL.t10 VSUBS 0.323971f
C1193 VTAIL.t15 VSUBS 0.323971f
C1194 VTAIL.n14 VSUBS 2.45238f
C1195 VTAIL.n15 VSUBS 1.22246f
C1196 VTAIL.t16 VSUBS 3.21683f
C1197 VTAIL.n16 VSUBS 2.86927f
C1198 VTAIL.t5 VSUBS 3.21683f
C1199 VTAIL.n17 VSUBS 2.86927f
C1200 VTAIL.t7 VSUBS 0.323971f
C1201 VTAIL.t2 VSUBS 0.323971f
C1202 VTAIL.n18 VSUBS 2.45238f
C1203 VTAIL.n19 VSUBS 1.00774f
C1204 VDD1.t6 VSUBS 3.57272f
C1205 VDD1.t1 VSUBS 0.336747f
C1206 VDD1.t2 VSUBS 0.336747f
C1207 VDD1.n0 VSUBS 2.7175f
C1208 VDD1.n1 VSUBS 1.85841f
C1209 VDD1.t7 VSUBS 3.5727f
C1210 VDD1.t0 VSUBS 0.336747f
C1211 VDD1.t4 VSUBS 0.336747f
C1212 VDD1.n2 VSUBS 2.7175f
C1213 VDD1.n3 VSUBS 1.84853f
C1214 VDD1.t3 VSUBS 0.336747f
C1215 VDD1.t9 VSUBS 0.336747f
C1216 VDD1.n4 VSUBS 2.74971f
C1217 VDD1.n5 VSUBS 4.47139f
C1218 VDD1.t5 VSUBS 0.336747f
C1219 VDD1.t8 VSUBS 0.336747f
C1220 VDD1.n6 VSUBS 2.71749f
C1221 VDD1.n7 VSUBS 4.58993f
C1222 VP.t2 VSUBS 3.23646f
C1223 VP.n0 VSUBS 1.22566f
C1224 VP.n1 VSUBS 0.025965f
C1225 VP.n2 VSUBS 0.021087f
C1226 VP.n3 VSUBS 0.025965f
C1227 VP.t8 VSUBS 3.23646f
C1228 VP.n4 VSUBS 1.12854f
C1229 VP.n5 VSUBS 0.025965f
C1230 VP.n6 VSUBS 0.02102f
C1231 VP.n7 VSUBS 0.025965f
C1232 VP.t5 VSUBS 3.23646f
C1233 VP.n8 VSUBS 1.12854f
C1234 VP.n9 VSUBS 0.025965f
C1235 VP.n10 VSUBS 0.02102f
C1236 VP.n11 VSUBS 0.025965f
C1237 VP.t1 VSUBS 3.23646f
C1238 VP.n12 VSUBS 1.12854f
C1239 VP.n13 VSUBS 0.025965f
C1240 VP.n14 VSUBS 0.021087f
C1241 VP.n15 VSUBS 0.025965f
C1242 VP.t6 VSUBS 3.23646f
C1243 VP.n16 VSUBS 1.22566f
C1244 VP.t3 VSUBS 3.23646f
C1245 VP.n17 VSUBS 1.22566f
C1246 VP.n18 VSUBS 0.025965f
C1247 VP.n19 VSUBS 0.021087f
C1248 VP.n20 VSUBS 0.025965f
C1249 VP.t4 VSUBS 3.23646f
C1250 VP.n21 VSUBS 1.12854f
C1251 VP.n22 VSUBS 0.025965f
C1252 VP.n23 VSUBS 0.02102f
C1253 VP.n24 VSUBS 0.025965f
C1254 VP.t9 VSUBS 3.23646f
C1255 VP.n25 VSUBS 1.12854f
C1256 VP.n26 VSUBS 0.025965f
C1257 VP.n27 VSUBS 0.02102f
C1258 VP.n28 VSUBS 0.025965f
C1259 VP.t0 VSUBS 3.23646f
C1260 VP.n29 VSUBS 1.21475f
C1261 VP.t7 VSUBS 3.53978f
C1262 VP.n30 VSUBS 1.16541f
C1263 VP.n31 VSUBS 0.302027f
C1264 VP.n32 VSUBS 0.037109f
C1265 VP.n33 VSUBS 0.048635f
C1266 VP.n34 VSUBS 0.051745f
C1267 VP.n35 VSUBS 0.025965f
C1268 VP.n36 VSUBS 0.025965f
C1269 VP.n37 VSUBS 0.025965f
C1270 VP.n38 VSUBS 0.052008f
C1271 VP.n39 VSUBS 0.048635f
C1272 VP.n40 VSUBS 0.036628f
C1273 VP.n41 VSUBS 0.025965f
C1274 VP.n42 VSUBS 0.025965f
C1275 VP.n43 VSUBS 0.036628f
C1276 VP.n44 VSUBS 0.048635f
C1277 VP.n45 VSUBS 0.052008f
C1278 VP.n46 VSUBS 0.025965f
C1279 VP.n47 VSUBS 0.025965f
C1280 VP.n48 VSUBS 0.025965f
C1281 VP.n49 VSUBS 0.051745f
C1282 VP.n50 VSUBS 0.048635f
C1283 VP.n51 VSUBS 0.037109f
C1284 VP.n52 VSUBS 0.025965f
C1285 VP.n53 VSUBS 0.025965f
C1286 VP.n54 VSUBS 0.036148f
C1287 VP.n55 VSUBS 0.048635f
C1288 VP.n56 VSUBS 0.052237f
C1289 VP.n57 VSUBS 0.025965f
C1290 VP.n58 VSUBS 0.025965f
C1291 VP.n59 VSUBS 0.025965f
C1292 VP.n60 VSUBS 0.051449f
C1293 VP.n61 VSUBS 0.048635f
C1294 VP.n62 VSUBS 0.037589f
C1295 VP.n63 VSUBS 0.041914f
C1296 VP.n64 VSUBS 1.81887f
C1297 VP.n65 VSUBS 1.83489f
C1298 VP.n66 VSUBS 0.041914f
C1299 VP.n67 VSUBS 0.037589f
C1300 VP.n68 VSUBS 0.048635f
C1301 VP.n69 VSUBS 0.051449f
C1302 VP.n70 VSUBS 0.025965f
C1303 VP.n71 VSUBS 0.025965f
C1304 VP.n72 VSUBS 0.025965f
C1305 VP.n73 VSUBS 0.052237f
C1306 VP.n74 VSUBS 0.048635f
C1307 VP.n75 VSUBS 0.036148f
C1308 VP.n76 VSUBS 0.025965f
C1309 VP.n77 VSUBS 0.025965f
C1310 VP.n78 VSUBS 0.037109f
C1311 VP.n79 VSUBS 0.048635f
C1312 VP.n80 VSUBS 0.051745f
C1313 VP.n81 VSUBS 0.025965f
C1314 VP.n82 VSUBS 0.025965f
C1315 VP.n83 VSUBS 0.025965f
C1316 VP.n84 VSUBS 0.052008f
C1317 VP.n85 VSUBS 0.048635f
C1318 VP.n86 VSUBS 0.036628f
C1319 VP.n87 VSUBS 0.025965f
C1320 VP.n88 VSUBS 0.025965f
C1321 VP.n89 VSUBS 0.036628f
C1322 VP.n90 VSUBS 0.048635f
C1323 VP.n91 VSUBS 0.052008f
C1324 VP.n92 VSUBS 0.025965f
C1325 VP.n93 VSUBS 0.025965f
C1326 VP.n94 VSUBS 0.025965f
C1327 VP.n95 VSUBS 0.051745f
C1328 VP.n96 VSUBS 0.048635f
C1329 VP.n97 VSUBS 0.037109f
C1330 VP.n98 VSUBS 0.025965f
C1331 VP.n99 VSUBS 0.025965f
C1332 VP.n100 VSUBS 0.036148f
C1333 VP.n101 VSUBS 0.048635f
C1334 VP.n102 VSUBS 0.052237f
C1335 VP.n103 VSUBS 0.025965f
C1336 VP.n104 VSUBS 0.025965f
C1337 VP.n105 VSUBS 0.025965f
C1338 VP.n106 VSUBS 0.051449f
C1339 VP.n107 VSUBS 0.048635f
C1340 VP.n108 VSUBS 0.037589f
C1341 VP.n109 VSUBS 0.041914f
C1342 VP.n110 VSUBS 0.063037f
.ends

