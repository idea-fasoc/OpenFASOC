* NGSPICE file created from diff_pair_sample_0946.ext - technology: sky130A

.subckt diff_pair_sample_0946 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X1 VDD1.t9 VP.t0 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=2.7495 ps=14.88 w=7.05 l=2.94
X2 VTAIL.t3 VP.t1 VDD1.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X3 VDD2.t4 VN.t1 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X4 VDD2.t8 VN.t2 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=1.16325 ps=7.38 w=7.05 l=2.94
X5 VDD2.t1 VN.t3 VTAIL.t15 B.t8 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X6 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.94
X7 VTAIL.t14 VN.t4 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X8 VDD2.t9 VN.t5 VTAIL.t13 B.t23 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=2.7495 ps=14.88 w=7.05 l=2.94
X9 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X10 VDD1.t6 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=2.7495 ps=14.88 w=7.05 l=2.94
X11 VTAIL.t1 VP.t4 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X12 VTAIL.t4 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X13 VDD2.t2 VN.t6 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=1.16325 ps=7.38 w=7.05 l=2.94
X14 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.94
X15 VTAIL.t6 VP.t6 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X16 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.94
X17 VDD2.t0 VN.t7 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=2.7495 ps=14.88 w=7.05 l=2.94
X18 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=0 ps=0 w=7.05 l=2.94
X19 VDD1.t2 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=1.16325 ps=7.38 w=7.05 l=2.94
X20 VDD1.t1 VP.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.7495 pd=14.88 as=1.16325 ps=7.38 w=7.05 l=2.94
X21 VDD1.t0 VP.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X22 VTAIL.t10 VN.t8 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
X23 VTAIL.t9 VN.t9 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.16325 pd=7.38 as=1.16325 ps=7.38 w=7.05 l=2.94
R0 VN.n87 VN.n45 161.3
R1 VN.n86 VN.n85 161.3
R2 VN.n84 VN.n46 161.3
R3 VN.n83 VN.n82 161.3
R4 VN.n81 VN.n47 161.3
R5 VN.n80 VN.n79 161.3
R6 VN.n78 VN.n48 161.3
R7 VN.n77 VN.n76 161.3
R8 VN.n75 VN.n49 161.3
R9 VN.n74 VN.n73 161.3
R10 VN.n72 VN.n51 161.3
R11 VN.n71 VN.n70 161.3
R12 VN.n69 VN.n52 161.3
R13 VN.n68 VN.n67 161.3
R14 VN.n66 VN.n53 161.3
R15 VN.n65 VN.n64 161.3
R16 VN.n63 VN.n54 161.3
R17 VN.n62 VN.n61 161.3
R18 VN.n60 VN.n55 161.3
R19 VN.n59 VN.n58 161.3
R20 VN.n42 VN.n0 161.3
R21 VN.n41 VN.n40 161.3
R22 VN.n39 VN.n1 161.3
R23 VN.n38 VN.n37 161.3
R24 VN.n36 VN.n2 161.3
R25 VN.n35 VN.n34 161.3
R26 VN.n33 VN.n3 161.3
R27 VN.n32 VN.n31 161.3
R28 VN.n29 VN.n4 161.3
R29 VN.n28 VN.n27 161.3
R30 VN.n26 VN.n5 161.3
R31 VN.n25 VN.n24 161.3
R32 VN.n23 VN.n6 161.3
R33 VN.n22 VN.n21 161.3
R34 VN.n20 VN.n7 161.3
R35 VN.n19 VN.n18 161.3
R36 VN.n17 VN.n8 161.3
R37 VN.n16 VN.n15 161.3
R38 VN.n14 VN.n9 161.3
R39 VN.n13 VN.n12 161.3
R40 VN.n44 VN.n43 108.799
R41 VN.n89 VN.n88 108.799
R42 VN.n10 VN.t2 90.4745
R43 VN.n56 VN.t7 90.4745
R44 VN.n11 VN.n10 60.6237
R45 VN.n57 VN.n56 60.6237
R46 VN.n22 VN.t3 57.7913
R47 VN.n11 VN.t9 57.7913
R48 VN.n30 VN.t0 57.7913
R49 VN.n43 VN.t5 57.7913
R50 VN.n68 VN.t1 57.7913
R51 VN.n57 VN.t4 57.7913
R52 VN.n50 VN.t8 57.7913
R53 VN.n88 VN.t6 57.7913
R54 VN.n17 VN.n16 53.6055
R55 VN.n28 VN.n5 53.6055
R56 VN.n63 VN.n62 53.6055
R57 VN.n74 VN.n51 53.6055
R58 VN VN.n89 51.4716
R59 VN.n37 VN.n36 49.7204
R60 VN.n82 VN.n81 49.7204
R61 VN.n37 VN.n1 31.2664
R62 VN.n82 VN.n46 31.2664
R63 VN.n18 VN.n17 27.3813
R64 VN.n24 VN.n5 27.3813
R65 VN.n64 VN.n63 27.3813
R66 VN.n70 VN.n51 27.3813
R67 VN.n12 VN.n9 24.4675
R68 VN.n16 VN.n9 24.4675
R69 VN.n18 VN.n7 24.4675
R70 VN.n22 VN.n7 24.4675
R71 VN.n23 VN.n22 24.4675
R72 VN.n24 VN.n23 24.4675
R73 VN.n29 VN.n28 24.4675
R74 VN.n31 VN.n29 24.4675
R75 VN.n35 VN.n3 24.4675
R76 VN.n36 VN.n35 24.4675
R77 VN.n41 VN.n1 24.4675
R78 VN.n42 VN.n41 24.4675
R79 VN.n62 VN.n55 24.4675
R80 VN.n58 VN.n55 24.4675
R81 VN.n70 VN.n69 24.4675
R82 VN.n69 VN.n68 24.4675
R83 VN.n68 VN.n53 24.4675
R84 VN.n64 VN.n53 24.4675
R85 VN.n81 VN.n80 24.4675
R86 VN.n80 VN.n48 24.4675
R87 VN.n76 VN.n75 24.4675
R88 VN.n75 VN.n74 24.4675
R89 VN.n87 VN.n86 24.4675
R90 VN.n86 VN.n46 24.4675
R91 VN.n12 VN.n11 13.2127
R92 VN.n31 VN.n30 13.2127
R93 VN.n58 VN.n57 13.2127
R94 VN.n76 VN.n50 13.2127
R95 VN.n30 VN.n3 11.2553
R96 VN.n50 VN.n48 11.2553
R97 VN.n59 VN.n56 5.12434
R98 VN.n13 VN.n10 5.12434
R99 VN.n43 VN.n42 1.95786
R100 VN.n88 VN.n87 1.95786
R101 VN.n89 VN.n45 0.278367
R102 VN.n44 VN.n0 0.278367
R103 VN.n85 VN.n45 0.189894
R104 VN.n85 VN.n84 0.189894
R105 VN.n84 VN.n83 0.189894
R106 VN.n83 VN.n47 0.189894
R107 VN.n79 VN.n47 0.189894
R108 VN.n79 VN.n78 0.189894
R109 VN.n78 VN.n77 0.189894
R110 VN.n77 VN.n49 0.189894
R111 VN.n73 VN.n49 0.189894
R112 VN.n73 VN.n72 0.189894
R113 VN.n72 VN.n71 0.189894
R114 VN.n71 VN.n52 0.189894
R115 VN.n67 VN.n52 0.189894
R116 VN.n67 VN.n66 0.189894
R117 VN.n66 VN.n65 0.189894
R118 VN.n65 VN.n54 0.189894
R119 VN.n61 VN.n54 0.189894
R120 VN.n61 VN.n60 0.189894
R121 VN.n60 VN.n59 0.189894
R122 VN.n14 VN.n13 0.189894
R123 VN.n15 VN.n14 0.189894
R124 VN.n15 VN.n8 0.189894
R125 VN.n19 VN.n8 0.189894
R126 VN.n20 VN.n19 0.189894
R127 VN.n21 VN.n20 0.189894
R128 VN.n21 VN.n6 0.189894
R129 VN.n25 VN.n6 0.189894
R130 VN.n26 VN.n25 0.189894
R131 VN.n27 VN.n26 0.189894
R132 VN.n27 VN.n4 0.189894
R133 VN.n32 VN.n4 0.189894
R134 VN.n33 VN.n32 0.189894
R135 VN.n34 VN.n33 0.189894
R136 VN.n34 VN.n2 0.189894
R137 VN.n38 VN.n2 0.189894
R138 VN.n39 VN.n38 0.189894
R139 VN.n40 VN.n39 0.189894
R140 VN.n40 VN.n0 0.189894
R141 VN VN.n44 0.153454
R142 VDD2.n1 VDD2.t8 70.6567
R143 VDD2.n4 VDD2.t2 67.8379
R144 VDD2.n3 VDD2.n2 67.0882
R145 VDD2 VDD2.n7 67.0853
R146 VDD2.n6 VDD2.n5 65.0294
R147 VDD2.n1 VDD2.n0 65.0294
R148 VDD2.n4 VDD2.n3 43.183
R149 VDD2.n6 VDD2.n4 2.81947
R150 VDD2.n7 VDD2.t3 2.80901
R151 VDD2.n7 VDD2.t0 2.80901
R152 VDD2.n5 VDD2.t7 2.80901
R153 VDD2.n5 VDD2.t4 2.80901
R154 VDD2.n2 VDD2.t5 2.80901
R155 VDD2.n2 VDD2.t9 2.80901
R156 VDD2.n0 VDD2.t6 2.80901
R157 VDD2.n0 VDD2.t1 2.80901
R158 VDD2 VDD2.n6 0.763431
R159 VDD2.n3 VDD2.n1 0.649895
R160 VTAIL.n11 VTAIL.t11 51.1591
R161 VTAIL.n17 VTAIL.t13 51.1589
R162 VTAIL.n2 VTAIL.t0 51.1589
R163 VTAIL.n16 VTAIL.t19 51.1589
R164 VTAIL.n15 VTAIL.n14 48.3506
R165 VTAIL.n13 VTAIL.n12 48.3506
R166 VTAIL.n10 VTAIL.n9 48.3506
R167 VTAIL.n8 VTAIL.n7 48.3506
R168 VTAIL.n19 VTAIL.n18 48.3506
R169 VTAIL.n1 VTAIL.n0 48.3506
R170 VTAIL.n4 VTAIL.n3 48.3506
R171 VTAIL.n6 VTAIL.n5 48.3506
R172 VTAIL.n8 VTAIL.n6 24.0824
R173 VTAIL.n17 VTAIL.n16 21.2634
R174 VTAIL.n10 VTAIL.n8 2.81947
R175 VTAIL.n11 VTAIL.n10 2.81947
R176 VTAIL.n15 VTAIL.n13 2.81947
R177 VTAIL.n16 VTAIL.n15 2.81947
R178 VTAIL.n6 VTAIL.n4 2.81947
R179 VTAIL.n4 VTAIL.n2 2.81947
R180 VTAIL.n19 VTAIL.n17 2.81947
R181 VTAIL.n18 VTAIL.t15 2.80901
R182 VTAIL.n18 VTAIL.t18 2.80901
R183 VTAIL.n0 VTAIL.t16 2.80901
R184 VTAIL.n0 VTAIL.t9 2.80901
R185 VTAIL.n3 VTAIL.t2 2.80901
R186 VTAIL.n3 VTAIL.t1 2.80901
R187 VTAIL.n5 VTAIL.t5 2.80901
R188 VTAIL.n5 VTAIL.t6 2.80901
R189 VTAIL.n14 VTAIL.t8 2.80901
R190 VTAIL.n14 VTAIL.t4 2.80901
R191 VTAIL.n12 VTAIL.t7 2.80901
R192 VTAIL.n12 VTAIL.t3 2.80901
R193 VTAIL.n9 VTAIL.t17 2.80901
R194 VTAIL.n9 VTAIL.t14 2.80901
R195 VTAIL.n7 VTAIL.t12 2.80901
R196 VTAIL.n7 VTAIL.t10 2.80901
R197 VTAIL VTAIL.n1 2.17291
R198 VTAIL.n13 VTAIL.n11 1.87981
R199 VTAIL.n2 VTAIL.n1 1.87981
R200 VTAIL VTAIL.n19 0.647052
R201 B.n735 B.n734 585
R202 B.n737 B.n157 585
R203 B.n740 B.n739 585
R204 B.n741 B.n156 585
R205 B.n743 B.n742 585
R206 B.n745 B.n155 585
R207 B.n748 B.n747 585
R208 B.n749 B.n154 585
R209 B.n751 B.n750 585
R210 B.n753 B.n153 585
R211 B.n756 B.n755 585
R212 B.n757 B.n152 585
R213 B.n759 B.n758 585
R214 B.n761 B.n151 585
R215 B.n764 B.n763 585
R216 B.n765 B.n150 585
R217 B.n767 B.n766 585
R218 B.n769 B.n149 585
R219 B.n772 B.n771 585
R220 B.n773 B.n148 585
R221 B.n775 B.n774 585
R222 B.n777 B.n147 585
R223 B.n780 B.n779 585
R224 B.n781 B.n146 585
R225 B.n783 B.n782 585
R226 B.n785 B.n145 585
R227 B.n788 B.n787 585
R228 B.n790 B.n142 585
R229 B.n792 B.n791 585
R230 B.n794 B.n141 585
R231 B.n797 B.n796 585
R232 B.n798 B.n140 585
R233 B.n800 B.n799 585
R234 B.n802 B.n139 585
R235 B.n805 B.n804 585
R236 B.n806 B.n135 585
R237 B.n808 B.n807 585
R238 B.n810 B.n134 585
R239 B.n813 B.n812 585
R240 B.n814 B.n133 585
R241 B.n816 B.n815 585
R242 B.n818 B.n132 585
R243 B.n821 B.n820 585
R244 B.n822 B.n131 585
R245 B.n824 B.n823 585
R246 B.n826 B.n130 585
R247 B.n829 B.n828 585
R248 B.n830 B.n129 585
R249 B.n832 B.n831 585
R250 B.n834 B.n128 585
R251 B.n837 B.n836 585
R252 B.n838 B.n127 585
R253 B.n840 B.n839 585
R254 B.n842 B.n126 585
R255 B.n845 B.n844 585
R256 B.n846 B.n125 585
R257 B.n848 B.n847 585
R258 B.n850 B.n124 585
R259 B.n853 B.n852 585
R260 B.n854 B.n123 585
R261 B.n856 B.n855 585
R262 B.n858 B.n122 585
R263 B.n861 B.n860 585
R264 B.n862 B.n121 585
R265 B.n733 B.n119 585
R266 B.n865 B.n119 585
R267 B.n732 B.n118 585
R268 B.n866 B.n118 585
R269 B.n731 B.n117 585
R270 B.n867 B.n117 585
R271 B.n730 B.n729 585
R272 B.n729 B.n113 585
R273 B.n728 B.n112 585
R274 B.n873 B.n112 585
R275 B.n727 B.n111 585
R276 B.n874 B.n111 585
R277 B.n726 B.n110 585
R278 B.n875 B.n110 585
R279 B.n725 B.n724 585
R280 B.n724 B.n106 585
R281 B.n723 B.n105 585
R282 B.n881 B.n105 585
R283 B.n722 B.n104 585
R284 B.n882 B.n104 585
R285 B.n721 B.n103 585
R286 B.n883 B.n103 585
R287 B.n720 B.n719 585
R288 B.n719 B.n99 585
R289 B.n718 B.n98 585
R290 B.n889 B.n98 585
R291 B.n717 B.n97 585
R292 B.n890 B.n97 585
R293 B.n716 B.n96 585
R294 B.n891 B.n96 585
R295 B.n715 B.n714 585
R296 B.n714 B.n92 585
R297 B.n713 B.n91 585
R298 B.n897 B.n91 585
R299 B.n712 B.n90 585
R300 B.n898 B.n90 585
R301 B.n711 B.n89 585
R302 B.n899 B.n89 585
R303 B.n710 B.n709 585
R304 B.n709 B.n85 585
R305 B.n708 B.n84 585
R306 B.n905 B.n84 585
R307 B.n707 B.n83 585
R308 B.n906 B.n83 585
R309 B.n706 B.n82 585
R310 B.n907 B.n82 585
R311 B.n705 B.n704 585
R312 B.n704 B.n78 585
R313 B.n703 B.n77 585
R314 B.n913 B.n77 585
R315 B.n702 B.n76 585
R316 B.n914 B.n76 585
R317 B.n701 B.n75 585
R318 B.n915 B.n75 585
R319 B.n700 B.n699 585
R320 B.n699 B.n71 585
R321 B.n698 B.n70 585
R322 B.n921 B.n70 585
R323 B.n697 B.n69 585
R324 B.n922 B.n69 585
R325 B.n696 B.n68 585
R326 B.n923 B.n68 585
R327 B.n695 B.n694 585
R328 B.n694 B.n64 585
R329 B.n693 B.n63 585
R330 B.n929 B.n63 585
R331 B.n692 B.n62 585
R332 B.n930 B.n62 585
R333 B.n691 B.n61 585
R334 B.n931 B.n61 585
R335 B.n690 B.n689 585
R336 B.n689 B.n57 585
R337 B.n688 B.n56 585
R338 B.n937 B.n56 585
R339 B.n687 B.n55 585
R340 B.n938 B.n55 585
R341 B.n686 B.n54 585
R342 B.n939 B.n54 585
R343 B.n685 B.n684 585
R344 B.n684 B.n50 585
R345 B.n683 B.n49 585
R346 B.n945 B.n49 585
R347 B.n682 B.n48 585
R348 B.n946 B.n48 585
R349 B.n681 B.n47 585
R350 B.n947 B.n47 585
R351 B.n680 B.n679 585
R352 B.n679 B.n43 585
R353 B.n678 B.n42 585
R354 B.n953 B.n42 585
R355 B.n677 B.n41 585
R356 B.n954 B.n41 585
R357 B.n676 B.n40 585
R358 B.n955 B.n40 585
R359 B.n675 B.n674 585
R360 B.n674 B.n36 585
R361 B.n673 B.n35 585
R362 B.n961 B.n35 585
R363 B.n672 B.n34 585
R364 B.n962 B.n34 585
R365 B.n671 B.n33 585
R366 B.n963 B.n33 585
R367 B.n670 B.n669 585
R368 B.n669 B.n29 585
R369 B.n668 B.n28 585
R370 B.n969 B.n28 585
R371 B.n667 B.n27 585
R372 B.n970 B.n27 585
R373 B.n666 B.n26 585
R374 B.n971 B.n26 585
R375 B.n665 B.n664 585
R376 B.n664 B.n22 585
R377 B.n663 B.n21 585
R378 B.n977 B.n21 585
R379 B.n662 B.n20 585
R380 B.n978 B.n20 585
R381 B.n661 B.n19 585
R382 B.n979 B.n19 585
R383 B.n660 B.n659 585
R384 B.n659 B.n18 585
R385 B.n658 B.n14 585
R386 B.n985 B.n14 585
R387 B.n657 B.n13 585
R388 B.n986 B.n13 585
R389 B.n656 B.n12 585
R390 B.n987 B.n12 585
R391 B.n655 B.n654 585
R392 B.n654 B.n8 585
R393 B.n653 B.n7 585
R394 B.n993 B.n7 585
R395 B.n652 B.n6 585
R396 B.n994 B.n6 585
R397 B.n651 B.n5 585
R398 B.n995 B.n5 585
R399 B.n650 B.n649 585
R400 B.n649 B.n4 585
R401 B.n648 B.n158 585
R402 B.n648 B.n647 585
R403 B.n638 B.n159 585
R404 B.n160 B.n159 585
R405 B.n640 B.n639 585
R406 B.n641 B.n640 585
R407 B.n637 B.n165 585
R408 B.n165 B.n164 585
R409 B.n636 B.n635 585
R410 B.n635 B.n634 585
R411 B.n167 B.n166 585
R412 B.n627 B.n167 585
R413 B.n626 B.n625 585
R414 B.n628 B.n626 585
R415 B.n624 B.n172 585
R416 B.n172 B.n171 585
R417 B.n623 B.n622 585
R418 B.n622 B.n621 585
R419 B.n174 B.n173 585
R420 B.n175 B.n174 585
R421 B.n614 B.n613 585
R422 B.n615 B.n614 585
R423 B.n612 B.n180 585
R424 B.n180 B.n179 585
R425 B.n611 B.n610 585
R426 B.n610 B.n609 585
R427 B.n182 B.n181 585
R428 B.n183 B.n182 585
R429 B.n602 B.n601 585
R430 B.n603 B.n602 585
R431 B.n600 B.n187 585
R432 B.n191 B.n187 585
R433 B.n599 B.n598 585
R434 B.n598 B.n597 585
R435 B.n189 B.n188 585
R436 B.n190 B.n189 585
R437 B.n590 B.n589 585
R438 B.n591 B.n590 585
R439 B.n588 B.n196 585
R440 B.n196 B.n195 585
R441 B.n587 B.n586 585
R442 B.n586 B.n585 585
R443 B.n198 B.n197 585
R444 B.n199 B.n198 585
R445 B.n578 B.n577 585
R446 B.n579 B.n578 585
R447 B.n576 B.n204 585
R448 B.n204 B.n203 585
R449 B.n575 B.n574 585
R450 B.n574 B.n573 585
R451 B.n206 B.n205 585
R452 B.n207 B.n206 585
R453 B.n566 B.n565 585
R454 B.n567 B.n566 585
R455 B.n564 B.n212 585
R456 B.n212 B.n211 585
R457 B.n563 B.n562 585
R458 B.n562 B.n561 585
R459 B.n214 B.n213 585
R460 B.n215 B.n214 585
R461 B.n554 B.n553 585
R462 B.n555 B.n554 585
R463 B.n552 B.n220 585
R464 B.n220 B.n219 585
R465 B.n551 B.n550 585
R466 B.n550 B.n549 585
R467 B.n222 B.n221 585
R468 B.n223 B.n222 585
R469 B.n542 B.n541 585
R470 B.n543 B.n542 585
R471 B.n540 B.n228 585
R472 B.n228 B.n227 585
R473 B.n539 B.n538 585
R474 B.n538 B.n537 585
R475 B.n230 B.n229 585
R476 B.n231 B.n230 585
R477 B.n530 B.n529 585
R478 B.n531 B.n530 585
R479 B.n528 B.n236 585
R480 B.n236 B.n235 585
R481 B.n527 B.n526 585
R482 B.n526 B.n525 585
R483 B.n238 B.n237 585
R484 B.n239 B.n238 585
R485 B.n518 B.n517 585
R486 B.n519 B.n518 585
R487 B.n516 B.n243 585
R488 B.n247 B.n243 585
R489 B.n515 B.n514 585
R490 B.n514 B.n513 585
R491 B.n245 B.n244 585
R492 B.n246 B.n245 585
R493 B.n506 B.n505 585
R494 B.n507 B.n506 585
R495 B.n504 B.n252 585
R496 B.n252 B.n251 585
R497 B.n503 B.n502 585
R498 B.n502 B.n501 585
R499 B.n254 B.n253 585
R500 B.n255 B.n254 585
R501 B.n494 B.n493 585
R502 B.n495 B.n494 585
R503 B.n492 B.n260 585
R504 B.n260 B.n259 585
R505 B.n491 B.n490 585
R506 B.n490 B.n489 585
R507 B.n262 B.n261 585
R508 B.n263 B.n262 585
R509 B.n482 B.n481 585
R510 B.n483 B.n482 585
R511 B.n480 B.n268 585
R512 B.n268 B.n267 585
R513 B.n479 B.n478 585
R514 B.n478 B.n477 585
R515 B.n270 B.n269 585
R516 B.n271 B.n270 585
R517 B.n470 B.n469 585
R518 B.n471 B.n470 585
R519 B.n468 B.n276 585
R520 B.n276 B.n275 585
R521 B.n467 B.n466 585
R522 B.n466 B.n465 585
R523 B.n278 B.n277 585
R524 B.n279 B.n278 585
R525 B.n458 B.n457 585
R526 B.n459 B.n458 585
R527 B.n456 B.n284 585
R528 B.n284 B.n283 585
R529 B.n455 B.n454 585
R530 B.n454 B.n453 585
R531 B.n450 B.n288 585
R532 B.n449 B.n448 585
R533 B.n446 B.n289 585
R534 B.n446 B.n287 585
R535 B.n445 B.n444 585
R536 B.n443 B.n442 585
R537 B.n441 B.n291 585
R538 B.n439 B.n438 585
R539 B.n437 B.n292 585
R540 B.n436 B.n435 585
R541 B.n433 B.n293 585
R542 B.n431 B.n430 585
R543 B.n429 B.n294 585
R544 B.n428 B.n427 585
R545 B.n425 B.n295 585
R546 B.n423 B.n422 585
R547 B.n421 B.n296 585
R548 B.n420 B.n419 585
R549 B.n417 B.n297 585
R550 B.n415 B.n414 585
R551 B.n413 B.n298 585
R552 B.n412 B.n411 585
R553 B.n409 B.n299 585
R554 B.n407 B.n406 585
R555 B.n405 B.n300 585
R556 B.n404 B.n403 585
R557 B.n401 B.n301 585
R558 B.n399 B.n398 585
R559 B.n396 B.n302 585
R560 B.n395 B.n394 585
R561 B.n392 B.n305 585
R562 B.n390 B.n389 585
R563 B.n388 B.n306 585
R564 B.n387 B.n386 585
R565 B.n384 B.n307 585
R566 B.n382 B.n381 585
R567 B.n380 B.n308 585
R568 B.n379 B.n378 585
R569 B.n376 B.n375 585
R570 B.n374 B.n373 585
R571 B.n372 B.n313 585
R572 B.n370 B.n369 585
R573 B.n368 B.n314 585
R574 B.n367 B.n366 585
R575 B.n364 B.n315 585
R576 B.n362 B.n361 585
R577 B.n360 B.n316 585
R578 B.n359 B.n358 585
R579 B.n356 B.n317 585
R580 B.n354 B.n353 585
R581 B.n352 B.n318 585
R582 B.n351 B.n350 585
R583 B.n348 B.n319 585
R584 B.n346 B.n345 585
R585 B.n344 B.n320 585
R586 B.n343 B.n342 585
R587 B.n340 B.n321 585
R588 B.n338 B.n337 585
R589 B.n336 B.n322 585
R590 B.n335 B.n334 585
R591 B.n332 B.n323 585
R592 B.n330 B.n329 585
R593 B.n328 B.n324 585
R594 B.n327 B.n326 585
R595 B.n286 B.n285 585
R596 B.n287 B.n286 585
R597 B.n452 B.n451 585
R598 B.n453 B.n452 585
R599 B.n282 B.n281 585
R600 B.n283 B.n282 585
R601 B.n461 B.n460 585
R602 B.n460 B.n459 585
R603 B.n462 B.n280 585
R604 B.n280 B.n279 585
R605 B.n464 B.n463 585
R606 B.n465 B.n464 585
R607 B.n274 B.n273 585
R608 B.n275 B.n274 585
R609 B.n473 B.n472 585
R610 B.n472 B.n471 585
R611 B.n474 B.n272 585
R612 B.n272 B.n271 585
R613 B.n476 B.n475 585
R614 B.n477 B.n476 585
R615 B.n266 B.n265 585
R616 B.n267 B.n266 585
R617 B.n485 B.n484 585
R618 B.n484 B.n483 585
R619 B.n486 B.n264 585
R620 B.n264 B.n263 585
R621 B.n488 B.n487 585
R622 B.n489 B.n488 585
R623 B.n258 B.n257 585
R624 B.n259 B.n258 585
R625 B.n497 B.n496 585
R626 B.n496 B.n495 585
R627 B.n498 B.n256 585
R628 B.n256 B.n255 585
R629 B.n500 B.n499 585
R630 B.n501 B.n500 585
R631 B.n250 B.n249 585
R632 B.n251 B.n250 585
R633 B.n509 B.n508 585
R634 B.n508 B.n507 585
R635 B.n510 B.n248 585
R636 B.n248 B.n246 585
R637 B.n512 B.n511 585
R638 B.n513 B.n512 585
R639 B.n242 B.n241 585
R640 B.n247 B.n242 585
R641 B.n521 B.n520 585
R642 B.n520 B.n519 585
R643 B.n522 B.n240 585
R644 B.n240 B.n239 585
R645 B.n524 B.n523 585
R646 B.n525 B.n524 585
R647 B.n234 B.n233 585
R648 B.n235 B.n234 585
R649 B.n533 B.n532 585
R650 B.n532 B.n531 585
R651 B.n534 B.n232 585
R652 B.n232 B.n231 585
R653 B.n536 B.n535 585
R654 B.n537 B.n536 585
R655 B.n226 B.n225 585
R656 B.n227 B.n226 585
R657 B.n545 B.n544 585
R658 B.n544 B.n543 585
R659 B.n546 B.n224 585
R660 B.n224 B.n223 585
R661 B.n548 B.n547 585
R662 B.n549 B.n548 585
R663 B.n218 B.n217 585
R664 B.n219 B.n218 585
R665 B.n557 B.n556 585
R666 B.n556 B.n555 585
R667 B.n558 B.n216 585
R668 B.n216 B.n215 585
R669 B.n560 B.n559 585
R670 B.n561 B.n560 585
R671 B.n210 B.n209 585
R672 B.n211 B.n210 585
R673 B.n569 B.n568 585
R674 B.n568 B.n567 585
R675 B.n570 B.n208 585
R676 B.n208 B.n207 585
R677 B.n572 B.n571 585
R678 B.n573 B.n572 585
R679 B.n202 B.n201 585
R680 B.n203 B.n202 585
R681 B.n581 B.n580 585
R682 B.n580 B.n579 585
R683 B.n582 B.n200 585
R684 B.n200 B.n199 585
R685 B.n584 B.n583 585
R686 B.n585 B.n584 585
R687 B.n194 B.n193 585
R688 B.n195 B.n194 585
R689 B.n593 B.n592 585
R690 B.n592 B.n591 585
R691 B.n594 B.n192 585
R692 B.n192 B.n190 585
R693 B.n596 B.n595 585
R694 B.n597 B.n596 585
R695 B.n186 B.n185 585
R696 B.n191 B.n186 585
R697 B.n605 B.n604 585
R698 B.n604 B.n603 585
R699 B.n606 B.n184 585
R700 B.n184 B.n183 585
R701 B.n608 B.n607 585
R702 B.n609 B.n608 585
R703 B.n178 B.n177 585
R704 B.n179 B.n178 585
R705 B.n617 B.n616 585
R706 B.n616 B.n615 585
R707 B.n618 B.n176 585
R708 B.n176 B.n175 585
R709 B.n620 B.n619 585
R710 B.n621 B.n620 585
R711 B.n170 B.n169 585
R712 B.n171 B.n170 585
R713 B.n630 B.n629 585
R714 B.n629 B.n628 585
R715 B.n631 B.n168 585
R716 B.n627 B.n168 585
R717 B.n633 B.n632 585
R718 B.n634 B.n633 585
R719 B.n163 B.n162 585
R720 B.n164 B.n163 585
R721 B.n643 B.n642 585
R722 B.n642 B.n641 585
R723 B.n644 B.n161 585
R724 B.n161 B.n160 585
R725 B.n646 B.n645 585
R726 B.n647 B.n646 585
R727 B.n2 B.n0 585
R728 B.n4 B.n2 585
R729 B.n3 B.n1 585
R730 B.n994 B.n3 585
R731 B.n992 B.n991 585
R732 B.n993 B.n992 585
R733 B.n990 B.n9 585
R734 B.n9 B.n8 585
R735 B.n989 B.n988 585
R736 B.n988 B.n987 585
R737 B.n11 B.n10 585
R738 B.n986 B.n11 585
R739 B.n984 B.n983 585
R740 B.n985 B.n984 585
R741 B.n982 B.n15 585
R742 B.n18 B.n15 585
R743 B.n981 B.n980 585
R744 B.n980 B.n979 585
R745 B.n17 B.n16 585
R746 B.n978 B.n17 585
R747 B.n976 B.n975 585
R748 B.n977 B.n976 585
R749 B.n974 B.n23 585
R750 B.n23 B.n22 585
R751 B.n973 B.n972 585
R752 B.n972 B.n971 585
R753 B.n25 B.n24 585
R754 B.n970 B.n25 585
R755 B.n968 B.n967 585
R756 B.n969 B.n968 585
R757 B.n966 B.n30 585
R758 B.n30 B.n29 585
R759 B.n965 B.n964 585
R760 B.n964 B.n963 585
R761 B.n32 B.n31 585
R762 B.n962 B.n32 585
R763 B.n960 B.n959 585
R764 B.n961 B.n960 585
R765 B.n958 B.n37 585
R766 B.n37 B.n36 585
R767 B.n957 B.n956 585
R768 B.n956 B.n955 585
R769 B.n39 B.n38 585
R770 B.n954 B.n39 585
R771 B.n952 B.n951 585
R772 B.n953 B.n952 585
R773 B.n950 B.n44 585
R774 B.n44 B.n43 585
R775 B.n949 B.n948 585
R776 B.n948 B.n947 585
R777 B.n46 B.n45 585
R778 B.n946 B.n46 585
R779 B.n944 B.n943 585
R780 B.n945 B.n944 585
R781 B.n942 B.n51 585
R782 B.n51 B.n50 585
R783 B.n941 B.n940 585
R784 B.n940 B.n939 585
R785 B.n53 B.n52 585
R786 B.n938 B.n53 585
R787 B.n936 B.n935 585
R788 B.n937 B.n936 585
R789 B.n934 B.n58 585
R790 B.n58 B.n57 585
R791 B.n933 B.n932 585
R792 B.n932 B.n931 585
R793 B.n60 B.n59 585
R794 B.n930 B.n60 585
R795 B.n928 B.n927 585
R796 B.n929 B.n928 585
R797 B.n926 B.n65 585
R798 B.n65 B.n64 585
R799 B.n925 B.n924 585
R800 B.n924 B.n923 585
R801 B.n67 B.n66 585
R802 B.n922 B.n67 585
R803 B.n920 B.n919 585
R804 B.n921 B.n920 585
R805 B.n918 B.n72 585
R806 B.n72 B.n71 585
R807 B.n917 B.n916 585
R808 B.n916 B.n915 585
R809 B.n74 B.n73 585
R810 B.n914 B.n74 585
R811 B.n912 B.n911 585
R812 B.n913 B.n912 585
R813 B.n910 B.n79 585
R814 B.n79 B.n78 585
R815 B.n909 B.n908 585
R816 B.n908 B.n907 585
R817 B.n81 B.n80 585
R818 B.n906 B.n81 585
R819 B.n904 B.n903 585
R820 B.n905 B.n904 585
R821 B.n902 B.n86 585
R822 B.n86 B.n85 585
R823 B.n901 B.n900 585
R824 B.n900 B.n899 585
R825 B.n88 B.n87 585
R826 B.n898 B.n88 585
R827 B.n896 B.n895 585
R828 B.n897 B.n896 585
R829 B.n894 B.n93 585
R830 B.n93 B.n92 585
R831 B.n893 B.n892 585
R832 B.n892 B.n891 585
R833 B.n95 B.n94 585
R834 B.n890 B.n95 585
R835 B.n888 B.n887 585
R836 B.n889 B.n888 585
R837 B.n886 B.n100 585
R838 B.n100 B.n99 585
R839 B.n885 B.n884 585
R840 B.n884 B.n883 585
R841 B.n102 B.n101 585
R842 B.n882 B.n102 585
R843 B.n880 B.n879 585
R844 B.n881 B.n880 585
R845 B.n878 B.n107 585
R846 B.n107 B.n106 585
R847 B.n877 B.n876 585
R848 B.n876 B.n875 585
R849 B.n109 B.n108 585
R850 B.n874 B.n109 585
R851 B.n872 B.n871 585
R852 B.n873 B.n872 585
R853 B.n870 B.n114 585
R854 B.n114 B.n113 585
R855 B.n869 B.n868 585
R856 B.n868 B.n867 585
R857 B.n116 B.n115 585
R858 B.n866 B.n116 585
R859 B.n864 B.n863 585
R860 B.n865 B.n864 585
R861 B.n997 B.n996 585
R862 B.n996 B.n995 585
R863 B.n452 B.n288 444.452
R864 B.n864 B.n121 444.452
R865 B.n454 B.n286 444.452
R866 B.n735 B.n119 444.452
R867 B.n309 B.t13 266.3
R868 B.n303 B.t9 266.3
R869 B.n136 B.t20 266.3
R870 B.n143 B.t16 266.3
R871 B.n736 B.n120 256.663
R872 B.n738 B.n120 256.663
R873 B.n744 B.n120 256.663
R874 B.n746 B.n120 256.663
R875 B.n752 B.n120 256.663
R876 B.n754 B.n120 256.663
R877 B.n760 B.n120 256.663
R878 B.n762 B.n120 256.663
R879 B.n768 B.n120 256.663
R880 B.n770 B.n120 256.663
R881 B.n776 B.n120 256.663
R882 B.n778 B.n120 256.663
R883 B.n784 B.n120 256.663
R884 B.n786 B.n120 256.663
R885 B.n793 B.n120 256.663
R886 B.n795 B.n120 256.663
R887 B.n801 B.n120 256.663
R888 B.n803 B.n120 256.663
R889 B.n809 B.n120 256.663
R890 B.n811 B.n120 256.663
R891 B.n817 B.n120 256.663
R892 B.n819 B.n120 256.663
R893 B.n825 B.n120 256.663
R894 B.n827 B.n120 256.663
R895 B.n833 B.n120 256.663
R896 B.n835 B.n120 256.663
R897 B.n841 B.n120 256.663
R898 B.n843 B.n120 256.663
R899 B.n849 B.n120 256.663
R900 B.n851 B.n120 256.663
R901 B.n857 B.n120 256.663
R902 B.n859 B.n120 256.663
R903 B.n447 B.n287 256.663
R904 B.n290 B.n287 256.663
R905 B.n440 B.n287 256.663
R906 B.n434 B.n287 256.663
R907 B.n432 B.n287 256.663
R908 B.n426 B.n287 256.663
R909 B.n424 B.n287 256.663
R910 B.n418 B.n287 256.663
R911 B.n416 B.n287 256.663
R912 B.n410 B.n287 256.663
R913 B.n408 B.n287 256.663
R914 B.n402 B.n287 256.663
R915 B.n400 B.n287 256.663
R916 B.n393 B.n287 256.663
R917 B.n391 B.n287 256.663
R918 B.n385 B.n287 256.663
R919 B.n383 B.n287 256.663
R920 B.n377 B.n287 256.663
R921 B.n312 B.n287 256.663
R922 B.n371 B.n287 256.663
R923 B.n365 B.n287 256.663
R924 B.n363 B.n287 256.663
R925 B.n357 B.n287 256.663
R926 B.n355 B.n287 256.663
R927 B.n349 B.n287 256.663
R928 B.n347 B.n287 256.663
R929 B.n341 B.n287 256.663
R930 B.n339 B.n287 256.663
R931 B.n333 B.n287 256.663
R932 B.n331 B.n287 256.663
R933 B.n325 B.n287 256.663
R934 B.n452 B.n282 163.367
R935 B.n460 B.n282 163.367
R936 B.n460 B.n280 163.367
R937 B.n464 B.n280 163.367
R938 B.n464 B.n274 163.367
R939 B.n472 B.n274 163.367
R940 B.n472 B.n272 163.367
R941 B.n476 B.n272 163.367
R942 B.n476 B.n266 163.367
R943 B.n484 B.n266 163.367
R944 B.n484 B.n264 163.367
R945 B.n488 B.n264 163.367
R946 B.n488 B.n258 163.367
R947 B.n496 B.n258 163.367
R948 B.n496 B.n256 163.367
R949 B.n500 B.n256 163.367
R950 B.n500 B.n250 163.367
R951 B.n508 B.n250 163.367
R952 B.n508 B.n248 163.367
R953 B.n512 B.n248 163.367
R954 B.n512 B.n242 163.367
R955 B.n520 B.n242 163.367
R956 B.n520 B.n240 163.367
R957 B.n524 B.n240 163.367
R958 B.n524 B.n234 163.367
R959 B.n532 B.n234 163.367
R960 B.n532 B.n232 163.367
R961 B.n536 B.n232 163.367
R962 B.n536 B.n226 163.367
R963 B.n544 B.n226 163.367
R964 B.n544 B.n224 163.367
R965 B.n548 B.n224 163.367
R966 B.n548 B.n218 163.367
R967 B.n556 B.n218 163.367
R968 B.n556 B.n216 163.367
R969 B.n560 B.n216 163.367
R970 B.n560 B.n210 163.367
R971 B.n568 B.n210 163.367
R972 B.n568 B.n208 163.367
R973 B.n572 B.n208 163.367
R974 B.n572 B.n202 163.367
R975 B.n580 B.n202 163.367
R976 B.n580 B.n200 163.367
R977 B.n584 B.n200 163.367
R978 B.n584 B.n194 163.367
R979 B.n592 B.n194 163.367
R980 B.n592 B.n192 163.367
R981 B.n596 B.n192 163.367
R982 B.n596 B.n186 163.367
R983 B.n604 B.n186 163.367
R984 B.n604 B.n184 163.367
R985 B.n608 B.n184 163.367
R986 B.n608 B.n178 163.367
R987 B.n616 B.n178 163.367
R988 B.n616 B.n176 163.367
R989 B.n620 B.n176 163.367
R990 B.n620 B.n170 163.367
R991 B.n629 B.n170 163.367
R992 B.n629 B.n168 163.367
R993 B.n633 B.n168 163.367
R994 B.n633 B.n163 163.367
R995 B.n642 B.n163 163.367
R996 B.n642 B.n161 163.367
R997 B.n646 B.n161 163.367
R998 B.n646 B.n2 163.367
R999 B.n996 B.n2 163.367
R1000 B.n996 B.n3 163.367
R1001 B.n992 B.n3 163.367
R1002 B.n992 B.n9 163.367
R1003 B.n988 B.n9 163.367
R1004 B.n988 B.n11 163.367
R1005 B.n984 B.n11 163.367
R1006 B.n984 B.n15 163.367
R1007 B.n980 B.n15 163.367
R1008 B.n980 B.n17 163.367
R1009 B.n976 B.n17 163.367
R1010 B.n976 B.n23 163.367
R1011 B.n972 B.n23 163.367
R1012 B.n972 B.n25 163.367
R1013 B.n968 B.n25 163.367
R1014 B.n968 B.n30 163.367
R1015 B.n964 B.n30 163.367
R1016 B.n964 B.n32 163.367
R1017 B.n960 B.n32 163.367
R1018 B.n960 B.n37 163.367
R1019 B.n956 B.n37 163.367
R1020 B.n956 B.n39 163.367
R1021 B.n952 B.n39 163.367
R1022 B.n952 B.n44 163.367
R1023 B.n948 B.n44 163.367
R1024 B.n948 B.n46 163.367
R1025 B.n944 B.n46 163.367
R1026 B.n944 B.n51 163.367
R1027 B.n940 B.n51 163.367
R1028 B.n940 B.n53 163.367
R1029 B.n936 B.n53 163.367
R1030 B.n936 B.n58 163.367
R1031 B.n932 B.n58 163.367
R1032 B.n932 B.n60 163.367
R1033 B.n928 B.n60 163.367
R1034 B.n928 B.n65 163.367
R1035 B.n924 B.n65 163.367
R1036 B.n924 B.n67 163.367
R1037 B.n920 B.n67 163.367
R1038 B.n920 B.n72 163.367
R1039 B.n916 B.n72 163.367
R1040 B.n916 B.n74 163.367
R1041 B.n912 B.n74 163.367
R1042 B.n912 B.n79 163.367
R1043 B.n908 B.n79 163.367
R1044 B.n908 B.n81 163.367
R1045 B.n904 B.n81 163.367
R1046 B.n904 B.n86 163.367
R1047 B.n900 B.n86 163.367
R1048 B.n900 B.n88 163.367
R1049 B.n896 B.n88 163.367
R1050 B.n896 B.n93 163.367
R1051 B.n892 B.n93 163.367
R1052 B.n892 B.n95 163.367
R1053 B.n888 B.n95 163.367
R1054 B.n888 B.n100 163.367
R1055 B.n884 B.n100 163.367
R1056 B.n884 B.n102 163.367
R1057 B.n880 B.n102 163.367
R1058 B.n880 B.n107 163.367
R1059 B.n876 B.n107 163.367
R1060 B.n876 B.n109 163.367
R1061 B.n872 B.n109 163.367
R1062 B.n872 B.n114 163.367
R1063 B.n868 B.n114 163.367
R1064 B.n868 B.n116 163.367
R1065 B.n864 B.n116 163.367
R1066 B.n448 B.n446 163.367
R1067 B.n446 B.n445 163.367
R1068 B.n442 B.n441 163.367
R1069 B.n439 B.n292 163.367
R1070 B.n435 B.n433 163.367
R1071 B.n431 B.n294 163.367
R1072 B.n427 B.n425 163.367
R1073 B.n423 B.n296 163.367
R1074 B.n419 B.n417 163.367
R1075 B.n415 B.n298 163.367
R1076 B.n411 B.n409 163.367
R1077 B.n407 B.n300 163.367
R1078 B.n403 B.n401 163.367
R1079 B.n399 B.n302 163.367
R1080 B.n394 B.n392 163.367
R1081 B.n390 B.n306 163.367
R1082 B.n386 B.n384 163.367
R1083 B.n382 B.n308 163.367
R1084 B.n378 B.n376 163.367
R1085 B.n373 B.n372 163.367
R1086 B.n370 B.n314 163.367
R1087 B.n366 B.n364 163.367
R1088 B.n362 B.n316 163.367
R1089 B.n358 B.n356 163.367
R1090 B.n354 B.n318 163.367
R1091 B.n350 B.n348 163.367
R1092 B.n346 B.n320 163.367
R1093 B.n342 B.n340 163.367
R1094 B.n338 B.n322 163.367
R1095 B.n334 B.n332 163.367
R1096 B.n330 B.n324 163.367
R1097 B.n326 B.n286 163.367
R1098 B.n454 B.n284 163.367
R1099 B.n458 B.n284 163.367
R1100 B.n458 B.n278 163.367
R1101 B.n466 B.n278 163.367
R1102 B.n466 B.n276 163.367
R1103 B.n470 B.n276 163.367
R1104 B.n470 B.n270 163.367
R1105 B.n478 B.n270 163.367
R1106 B.n478 B.n268 163.367
R1107 B.n482 B.n268 163.367
R1108 B.n482 B.n262 163.367
R1109 B.n490 B.n262 163.367
R1110 B.n490 B.n260 163.367
R1111 B.n494 B.n260 163.367
R1112 B.n494 B.n254 163.367
R1113 B.n502 B.n254 163.367
R1114 B.n502 B.n252 163.367
R1115 B.n506 B.n252 163.367
R1116 B.n506 B.n245 163.367
R1117 B.n514 B.n245 163.367
R1118 B.n514 B.n243 163.367
R1119 B.n518 B.n243 163.367
R1120 B.n518 B.n238 163.367
R1121 B.n526 B.n238 163.367
R1122 B.n526 B.n236 163.367
R1123 B.n530 B.n236 163.367
R1124 B.n530 B.n230 163.367
R1125 B.n538 B.n230 163.367
R1126 B.n538 B.n228 163.367
R1127 B.n542 B.n228 163.367
R1128 B.n542 B.n222 163.367
R1129 B.n550 B.n222 163.367
R1130 B.n550 B.n220 163.367
R1131 B.n554 B.n220 163.367
R1132 B.n554 B.n214 163.367
R1133 B.n562 B.n214 163.367
R1134 B.n562 B.n212 163.367
R1135 B.n566 B.n212 163.367
R1136 B.n566 B.n206 163.367
R1137 B.n574 B.n206 163.367
R1138 B.n574 B.n204 163.367
R1139 B.n578 B.n204 163.367
R1140 B.n578 B.n198 163.367
R1141 B.n586 B.n198 163.367
R1142 B.n586 B.n196 163.367
R1143 B.n590 B.n196 163.367
R1144 B.n590 B.n189 163.367
R1145 B.n598 B.n189 163.367
R1146 B.n598 B.n187 163.367
R1147 B.n602 B.n187 163.367
R1148 B.n602 B.n182 163.367
R1149 B.n610 B.n182 163.367
R1150 B.n610 B.n180 163.367
R1151 B.n614 B.n180 163.367
R1152 B.n614 B.n174 163.367
R1153 B.n622 B.n174 163.367
R1154 B.n622 B.n172 163.367
R1155 B.n626 B.n172 163.367
R1156 B.n626 B.n167 163.367
R1157 B.n635 B.n167 163.367
R1158 B.n635 B.n165 163.367
R1159 B.n640 B.n165 163.367
R1160 B.n640 B.n159 163.367
R1161 B.n648 B.n159 163.367
R1162 B.n649 B.n648 163.367
R1163 B.n649 B.n5 163.367
R1164 B.n6 B.n5 163.367
R1165 B.n7 B.n6 163.367
R1166 B.n654 B.n7 163.367
R1167 B.n654 B.n12 163.367
R1168 B.n13 B.n12 163.367
R1169 B.n14 B.n13 163.367
R1170 B.n659 B.n14 163.367
R1171 B.n659 B.n19 163.367
R1172 B.n20 B.n19 163.367
R1173 B.n21 B.n20 163.367
R1174 B.n664 B.n21 163.367
R1175 B.n664 B.n26 163.367
R1176 B.n27 B.n26 163.367
R1177 B.n28 B.n27 163.367
R1178 B.n669 B.n28 163.367
R1179 B.n669 B.n33 163.367
R1180 B.n34 B.n33 163.367
R1181 B.n35 B.n34 163.367
R1182 B.n674 B.n35 163.367
R1183 B.n674 B.n40 163.367
R1184 B.n41 B.n40 163.367
R1185 B.n42 B.n41 163.367
R1186 B.n679 B.n42 163.367
R1187 B.n679 B.n47 163.367
R1188 B.n48 B.n47 163.367
R1189 B.n49 B.n48 163.367
R1190 B.n684 B.n49 163.367
R1191 B.n684 B.n54 163.367
R1192 B.n55 B.n54 163.367
R1193 B.n56 B.n55 163.367
R1194 B.n689 B.n56 163.367
R1195 B.n689 B.n61 163.367
R1196 B.n62 B.n61 163.367
R1197 B.n63 B.n62 163.367
R1198 B.n694 B.n63 163.367
R1199 B.n694 B.n68 163.367
R1200 B.n69 B.n68 163.367
R1201 B.n70 B.n69 163.367
R1202 B.n699 B.n70 163.367
R1203 B.n699 B.n75 163.367
R1204 B.n76 B.n75 163.367
R1205 B.n77 B.n76 163.367
R1206 B.n704 B.n77 163.367
R1207 B.n704 B.n82 163.367
R1208 B.n83 B.n82 163.367
R1209 B.n84 B.n83 163.367
R1210 B.n709 B.n84 163.367
R1211 B.n709 B.n89 163.367
R1212 B.n90 B.n89 163.367
R1213 B.n91 B.n90 163.367
R1214 B.n714 B.n91 163.367
R1215 B.n714 B.n96 163.367
R1216 B.n97 B.n96 163.367
R1217 B.n98 B.n97 163.367
R1218 B.n719 B.n98 163.367
R1219 B.n719 B.n103 163.367
R1220 B.n104 B.n103 163.367
R1221 B.n105 B.n104 163.367
R1222 B.n724 B.n105 163.367
R1223 B.n724 B.n110 163.367
R1224 B.n111 B.n110 163.367
R1225 B.n112 B.n111 163.367
R1226 B.n729 B.n112 163.367
R1227 B.n729 B.n117 163.367
R1228 B.n118 B.n117 163.367
R1229 B.n119 B.n118 163.367
R1230 B.n860 B.n858 163.367
R1231 B.n856 B.n123 163.367
R1232 B.n852 B.n850 163.367
R1233 B.n848 B.n125 163.367
R1234 B.n844 B.n842 163.367
R1235 B.n840 B.n127 163.367
R1236 B.n836 B.n834 163.367
R1237 B.n832 B.n129 163.367
R1238 B.n828 B.n826 163.367
R1239 B.n824 B.n131 163.367
R1240 B.n820 B.n818 163.367
R1241 B.n816 B.n133 163.367
R1242 B.n812 B.n810 163.367
R1243 B.n808 B.n135 163.367
R1244 B.n804 B.n802 163.367
R1245 B.n800 B.n140 163.367
R1246 B.n796 B.n794 163.367
R1247 B.n792 B.n142 163.367
R1248 B.n787 B.n785 163.367
R1249 B.n783 B.n146 163.367
R1250 B.n779 B.n777 163.367
R1251 B.n775 B.n148 163.367
R1252 B.n771 B.n769 163.367
R1253 B.n767 B.n150 163.367
R1254 B.n763 B.n761 163.367
R1255 B.n759 B.n152 163.367
R1256 B.n755 B.n753 163.367
R1257 B.n751 B.n154 163.367
R1258 B.n747 B.n745 163.367
R1259 B.n743 B.n156 163.367
R1260 B.n739 B.n737 163.367
R1261 B.n309 B.t15 137.212
R1262 B.n143 B.t18 137.212
R1263 B.n303 B.t12 137.203
R1264 B.n136 B.t21 137.203
R1265 B.n453 B.n287 99.0674
R1266 B.n865 B.n120 99.0674
R1267 B.n310 B.t14 73.7934
R1268 B.n144 B.t19 73.7934
R1269 B.n304 B.t11 73.7857
R1270 B.n137 B.t22 73.7857
R1271 B.n447 B.n288 71.676
R1272 B.n445 B.n290 71.676
R1273 B.n441 B.n440 71.676
R1274 B.n434 B.n292 71.676
R1275 B.n433 B.n432 71.676
R1276 B.n426 B.n294 71.676
R1277 B.n425 B.n424 71.676
R1278 B.n418 B.n296 71.676
R1279 B.n417 B.n416 71.676
R1280 B.n410 B.n298 71.676
R1281 B.n409 B.n408 71.676
R1282 B.n402 B.n300 71.676
R1283 B.n401 B.n400 71.676
R1284 B.n393 B.n302 71.676
R1285 B.n392 B.n391 71.676
R1286 B.n385 B.n306 71.676
R1287 B.n384 B.n383 71.676
R1288 B.n377 B.n308 71.676
R1289 B.n376 B.n312 71.676
R1290 B.n372 B.n371 71.676
R1291 B.n365 B.n314 71.676
R1292 B.n364 B.n363 71.676
R1293 B.n357 B.n316 71.676
R1294 B.n356 B.n355 71.676
R1295 B.n349 B.n318 71.676
R1296 B.n348 B.n347 71.676
R1297 B.n341 B.n320 71.676
R1298 B.n340 B.n339 71.676
R1299 B.n333 B.n322 71.676
R1300 B.n332 B.n331 71.676
R1301 B.n325 B.n324 71.676
R1302 B.n859 B.n121 71.676
R1303 B.n858 B.n857 71.676
R1304 B.n851 B.n123 71.676
R1305 B.n850 B.n849 71.676
R1306 B.n843 B.n125 71.676
R1307 B.n842 B.n841 71.676
R1308 B.n835 B.n127 71.676
R1309 B.n834 B.n833 71.676
R1310 B.n827 B.n129 71.676
R1311 B.n826 B.n825 71.676
R1312 B.n819 B.n131 71.676
R1313 B.n818 B.n817 71.676
R1314 B.n811 B.n133 71.676
R1315 B.n810 B.n809 71.676
R1316 B.n803 B.n135 71.676
R1317 B.n802 B.n801 71.676
R1318 B.n795 B.n140 71.676
R1319 B.n794 B.n793 71.676
R1320 B.n786 B.n142 71.676
R1321 B.n785 B.n784 71.676
R1322 B.n778 B.n146 71.676
R1323 B.n777 B.n776 71.676
R1324 B.n770 B.n148 71.676
R1325 B.n769 B.n768 71.676
R1326 B.n762 B.n150 71.676
R1327 B.n761 B.n760 71.676
R1328 B.n754 B.n152 71.676
R1329 B.n753 B.n752 71.676
R1330 B.n746 B.n154 71.676
R1331 B.n745 B.n744 71.676
R1332 B.n738 B.n156 71.676
R1333 B.n737 B.n736 71.676
R1334 B.n736 B.n735 71.676
R1335 B.n739 B.n738 71.676
R1336 B.n744 B.n743 71.676
R1337 B.n747 B.n746 71.676
R1338 B.n752 B.n751 71.676
R1339 B.n755 B.n754 71.676
R1340 B.n760 B.n759 71.676
R1341 B.n763 B.n762 71.676
R1342 B.n768 B.n767 71.676
R1343 B.n771 B.n770 71.676
R1344 B.n776 B.n775 71.676
R1345 B.n779 B.n778 71.676
R1346 B.n784 B.n783 71.676
R1347 B.n787 B.n786 71.676
R1348 B.n793 B.n792 71.676
R1349 B.n796 B.n795 71.676
R1350 B.n801 B.n800 71.676
R1351 B.n804 B.n803 71.676
R1352 B.n809 B.n808 71.676
R1353 B.n812 B.n811 71.676
R1354 B.n817 B.n816 71.676
R1355 B.n820 B.n819 71.676
R1356 B.n825 B.n824 71.676
R1357 B.n828 B.n827 71.676
R1358 B.n833 B.n832 71.676
R1359 B.n836 B.n835 71.676
R1360 B.n841 B.n840 71.676
R1361 B.n844 B.n843 71.676
R1362 B.n849 B.n848 71.676
R1363 B.n852 B.n851 71.676
R1364 B.n857 B.n856 71.676
R1365 B.n860 B.n859 71.676
R1366 B.n448 B.n447 71.676
R1367 B.n442 B.n290 71.676
R1368 B.n440 B.n439 71.676
R1369 B.n435 B.n434 71.676
R1370 B.n432 B.n431 71.676
R1371 B.n427 B.n426 71.676
R1372 B.n424 B.n423 71.676
R1373 B.n419 B.n418 71.676
R1374 B.n416 B.n415 71.676
R1375 B.n411 B.n410 71.676
R1376 B.n408 B.n407 71.676
R1377 B.n403 B.n402 71.676
R1378 B.n400 B.n399 71.676
R1379 B.n394 B.n393 71.676
R1380 B.n391 B.n390 71.676
R1381 B.n386 B.n385 71.676
R1382 B.n383 B.n382 71.676
R1383 B.n378 B.n377 71.676
R1384 B.n373 B.n312 71.676
R1385 B.n371 B.n370 71.676
R1386 B.n366 B.n365 71.676
R1387 B.n363 B.n362 71.676
R1388 B.n358 B.n357 71.676
R1389 B.n355 B.n354 71.676
R1390 B.n350 B.n349 71.676
R1391 B.n347 B.n346 71.676
R1392 B.n342 B.n341 71.676
R1393 B.n339 B.n338 71.676
R1394 B.n334 B.n333 71.676
R1395 B.n331 B.n330 71.676
R1396 B.n326 B.n325 71.676
R1397 B.n310 B.n309 63.4187
R1398 B.n304 B.n303 63.4187
R1399 B.n137 B.n136 63.4187
R1400 B.n144 B.n143 63.4187
R1401 B.n453 B.n283 60.6902
R1402 B.n459 B.n283 60.6902
R1403 B.n459 B.n279 60.6902
R1404 B.n465 B.n279 60.6902
R1405 B.n465 B.n275 60.6902
R1406 B.n471 B.n275 60.6902
R1407 B.n471 B.n271 60.6902
R1408 B.n477 B.n271 60.6902
R1409 B.n483 B.n267 60.6902
R1410 B.n483 B.n263 60.6902
R1411 B.n489 B.n263 60.6902
R1412 B.n489 B.n259 60.6902
R1413 B.n495 B.n259 60.6902
R1414 B.n495 B.n255 60.6902
R1415 B.n501 B.n255 60.6902
R1416 B.n501 B.n251 60.6902
R1417 B.n507 B.n251 60.6902
R1418 B.n507 B.n246 60.6902
R1419 B.n513 B.n246 60.6902
R1420 B.n513 B.n247 60.6902
R1421 B.n519 B.n239 60.6902
R1422 B.n525 B.n239 60.6902
R1423 B.n525 B.n235 60.6902
R1424 B.n531 B.n235 60.6902
R1425 B.n531 B.n231 60.6902
R1426 B.n537 B.n231 60.6902
R1427 B.n537 B.n227 60.6902
R1428 B.n543 B.n227 60.6902
R1429 B.n549 B.n223 60.6902
R1430 B.n549 B.n219 60.6902
R1431 B.n555 B.n219 60.6902
R1432 B.n555 B.n215 60.6902
R1433 B.n561 B.n215 60.6902
R1434 B.n561 B.n211 60.6902
R1435 B.n567 B.n211 60.6902
R1436 B.n567 B.n207 60.6902
R1437 B.n573 B.n207 60.6902
R1438 B.n579 B.n203 60.6902
R1439 B.n579 B.n199 60.6902
R1440 B.n585 B.n199 60.6902
R1441 B.n585 B.n195 60.6902
R1442 B.n591 B.n195 60.6902
R1443 B.n591 B.n190 60.6902
R1444 B.n597 B.n190 60.6902
R1445 B.n597 B.n191 60.6902
R1446 B.n603 B.n183 60.6902
R1447 B.n609 B.n183 60.6902
R1448 B.n609 B.n179 60.6902
R1449 B.n615 B.n179 60.6902
R1450 B.n615 B.n175 60.6902
R1451 B.n621 B.n175 60.6902
R1452 B.n621 B.n171 60.6902
R1453 B.n628 B.n171 60.6902
R1454 B.n628 B.n627 60.6902
R1455 B.n634 B.n164 60.6902
R1456 B.n641 B.n164 60.6902
R1457 B.n641 B.n160 60.6902
R1458 B.n647 B.n160 60.6902
R1459 B.n647 B.n4 60.6902
R1460 B.n995 B.n4 60.6902
R1461 B.n995 B.n994 60.6902
R1462 B.n994 B.n993 60.6902
R1463 B.n993 B.n8 60.6902
R1464 B.n987 B.n8 60.6902
R1465 B.n987 B.n986 60.6902
R1466 B.n986 B.n985 60.6902
R1467 B.n979 B.n18 60.6902
R1468 B.n979 B.n978 60.6902
R1469 B.n978 B.n977 60.6902
R1470 B.n977 B.n22 60.6902
R1471 B.n971 B.n22 60.6902
R1472 B.n971 B.n970 60.6902
R1473 B.n970 B.n969 60.6902
R1474 B.n969 B.n29 60.6902
R1475 B.n963 B.n29 60.6902
R1476 B.n962 B.n961 60.6902
R1477 B.n961 B.n36 60.6902
R1478 B.n955 B.n36 60.6902
R1479 B.n955 B.n954 60.6902
R1480 B.n954 B.n953 60.6902
R1481 B.n953 B.n43 60.6902
R1482 B.n947 B.n43 60.6902
R1483 B.n947 B.n946 60.6902
R1484 B.n945 B.n50 60.6902
R1485 B.n939 B.n50 60.6902
R1486 B.n939 B.n938 60.6902
R1487 B.n938 B.n937 60.6902
R1488 B.n937 B.n57 60.6902
R1489 B.n931 B.n57 60.6902
R1490 B.n931 B.n930 60.6902
R1491 B.n930 B.n929 60.6902
R1492 B.n929 B.n64 60.6902
R1493 B.n923 B.n922 60.6902
R1494 B.n922 B.n921 60.6902
R1495 B.n921 B.n71 60.6902
R1496 B.n915 B.n71 60.6902
R1497 B.n915 B.n914 60.6902
R1498 B.n914 B.n913 60.6902
R1499 B.n913 B.n78 60.6902
R1500 B.n907 B.n78 60.6902
R1501 B.n906 B.n905 60.6902
R1502 B.n905 B.n85 60.6902
R1503 B.n899 B.n85 60.6902
R1504 B.n899 B.n898 60.6902
R1505 B.n898 B.n897 60.6902
R1506 B.n897 B.n92 60.6902
R1507 B.n891 B.n92 60.6902
R1508 B.n891 B.n890 60.6902
R1509 B.n890 B.n889 60.6902
R1510 B.n889 B.n99 60.6902
R1511 B.n883 B.n99 60.6902
R1512 B.n883 B.n882 60.6902
R1513 B.n881 B.n106 60.6902
R1514 B.n875 B.n106 60.6902
R1515 B.n875 B.n874 60.6902
R1516 B.n874 B.n873 60.6902
R1517 B.n873 B.n113 60.6902
R1518 B.n867 B.n113 60.6902
R1519 B.n867 B.n866 60.6902
R1520 B.n866 B.n865 60.6902
R1521 B.n311 B.n310 59.5399
R1522 B.n397 B.n304 59.5399
R1523 B.n138 B.n137 59.5399
R1524 B.n789 B.n144 59.5399
R1525 B.n191 B.t1 58.9052
R1526 B.t3 B.n962 58.9052
R1527 B.n519 B.t5 53.5502
R1528 B.n907 B.t23 53.5502
R1529 B.n543 B.t6 44.6252
R1530 B.n923 B.t4 44.6252
R1531 B.t10 B.n267 42.8403
R1532 B.n882 B.t17 42.8403
R1533 B.t2 B.n203 39.2703
R1534 B.n946 B.t8 39.2703
R1535 B.n627 B.t0 35.7003
R1536 B.n18 B.t7 35.7003
R1537 B.n863 B.n862 28.8785
R1538 B.n455 B.n285 28.8785
R1539 B.n451 B.n450 28.8785
R1540 B.n734 B.n733 28.8785
R1541 B.n634 B.t0 24.9904
R1542 B.n985 B.t7 24.9904
R1543 B.n573 B.t2 21.4204
R1544 B.t8 B.n945 21.4204
R1545 B B.n997 18.0485
R1546 B.n477 B.t10 17.8504
R1547 B.t17 B.n881 17.8504
R1548 B.t6 B.n223 16.0654
R1549 B.t4 B.n64 16.0654
R1550 B.n862 B.n861 10.6151
R1551 B.n861 B.n122 10.6151
R1552 B.n855 B.n122 10.6151
R1553 B.n855 B.n854 10.6151
R1554 B.n854 B.n853 10.6151
R1555 B.n853 B.n124 10.6151
R1556 B.n847 B.n124 10.6151
R1557 B.n847 B.n846 10.6151
R1558 B.n846 B.n845 10.6151
R1559 B.n845 B.n126 10.6151
R1560 B.n839 B.n126 10.6151
R1561 B.n839 B.n838 10.6151
R1562 B.n838 B.n837 10.6151
R1563 B.n837 B.n128 10.6151
R1564 B.n831 B.n128 10.6151
R1565 B.n831 B.n830 10.6151
R1566 B.n830 B.n829 10.6151
R1567 B.n829 B.n130 10.6151
R1568 B.n823 B.n130 10.6151
R1569 B.n823 B.n822 10.6151
R1570 B.n822 B.n821 10.6151
R1571 B.n821 B.n132 10.6151
R1572 B.n815 B.n132 10.6151
R1573 B.n815 B.n814 10.6151
R1574 B.n814 B.n813 10.6151
R1575 B.n813 B.n134 10.6151
R1576 B.n807 B.n806 10.6151
R1577 B.n806 B.n805 10.6151
R1578 B.n805 B.n139 10.6151
R1579 B.n799 B.n139 10.6151
R1580 B.n799 B.n798 10.6151
R1581 B.n798 B.n797 10.6151
R1582 B.n797 B.n141 10.6151
R1583 B.n791 B.n141 10.6151
R1584 B.n791 B.n790 10.6151
R1585 B.n788 B.n145 10.6151
R1586 B.n782 B.n145 10.6151
R1587 B.n782 B.n781 10.6151
R1588 B.n781 B.n780 10.6151
R1589 B.n780 B.n147 10.6151
R1590 B.n774 B.n147 10.6151
R1591 B.n774 B.n773 10.6151
R1592 B.n773 B.n772 10.6151
R1593 B.n772 B.n149 10.6151
R1594 B.n766 B.n149 10.6151
R1595 B.n766 B.n765 10.6151
R1596 B.n765 B.n764 10.6151
R1597 B.n764 B.n151 10.6151
R1598 B.n758 B.n151 10.6151
R1599 B.n758 B.n757 10.6151
R1600 B.n757 B.n756 10.6151
R1601 B.n756 B.n153 10.6151
R1602 B.n750 B.n153 10.6151
R1603 B.n750 B.n749 10.6151
R1604 B.n749 B.n748 10.6151
R1605 B.n748 B.n155 10.6151
R1606 B.n742 B.n155 10.6151
R1607 B.n742 B.n741 10.6151
R1608 B.n741 B.n740 10.6151
R1609 B.n740 B.n157 10.6151
R1610 B.n734 B.n157 10.6151
R1611 B.n456 B.n455 10.6151
R1612 B.n457 B.n456 10.6151
R1613 B.n457 B.n277 10.6151
R1614 B.n467 B.n277 10.6151
R1615 B.n468 B.n467 10.6151
R1616 B.n469 B.n468 10.6151
R1617 B.n469 B.n269 10.6151
R1618 B.n479 B.n269 10.6151
R1619 B.n480 B.n479 10.6151
R1620 B.n481 B.n480 10.6151
R1621 B.n481 B.n261 10.6151
R1622 B.n491 B.n261 10.6151
R1623 B.n492 B.n491 10.6151
R1624 B.n493 B.n492 10.6151
R1625 B.n493 B.n253 10.6151
R1626 B.n503 B.n253 10.6151
R1627 B.n504 B.n503 10.6151
R1628 B.n505 B.n504 10.6151
R1629 B.n505 B.n244 10.6151
R1630 B.n515 B.n244 10.6151
R1631 B.n516 B.n515 10.6151
R1632 B.n517 B.n516 10.6151
R1633 B.n517 B.n237 10.6151
R1634 B.n527 B.n237 10.6151
R1635 B.n528 B.n527 10.6151
R1636 B.n529 B.n528 10.6151
R1637 B.n529 B.n229 10.6151
R1638 B.n539 B.n229 10.6151
R1639 B.n540 B.n539 10.6151
R1640 B.n541 B.n540 10.6151
R1641 B.n541 B.n221 10.6151
R1642 B.n551 B.n221 10.6151
R1643 B.n552 B.n551 10.6151
R1644 B.n553 B.n552 10.6151
R1645 B.n553 B.n213 10.6151
R1646 B.n563 B.n213 10.6151
R1647 B.n564 B.n563 10.6151
R1648 B.n565 B.n564 10.6151
R1649 B.n565 B.n205 10.6151
R1650 B.n575 B.n205 10.6151
R1651 B.n576 B.n575 10.6151
R1652 B.n577 B.n576 10.6151
R1653 B.n577 B.n197 10.6151
R1654 B.n587 B.n197 10.6151
R1655 B.n588 B.n587 10.6151
R1656 B.n589 B.n588 10.6151
R1657 B.n589 B.n188 10.6151
R1658 B.n599 B.n188 10.6151
R1659 B.n600 B.n599 10.6151
R1660 B.n601 B.n600 10.6151
R1661 B.n601 B.n181 10.6151
R1662 B.n611 B.n181 10.6151
R1663 B.n612 B.n611 10.6151
R1664 B.n613 B.n612 10.6151
R1665 B.n613 B.n173 10.6151
R1666 B.n623 B.n173 10.6151
R1667 B.n624 B.n623 10.6151
R1668 B.n625 B.n624 10.6151
R1669 B.n625 B.n166 10.6151
R1670 B.n636 B.n166 10.6151
R1671 B.n637 B.n636 10.6151
R1672 B.n639 B.n637 10.6151
R1673 B.n639 B.n638 10.6151
R1674 B.n638 B.n158 10.6151
R1675 B.n650 B.n158 10.6151
R1676 B.n651 B.n650 10.6151
R1677 B.n652 B.n651 10.6151
R1678 B.n653 B.n652 10.6151
R1679 B.n655 B.n653 10.6151
R1680 B.n656 B.n655 10.6151
R1681 B.n657 B.n656 10.6151
R1682 B.n658 B.n657 10.6151
R1683 B.n660 B.n658 10.6151
R1684 B.n661 B.n660 10.6151
R1685 B.n662 B.n661 10.6151
R1686 B.n663 B.n662 10.6151
R1687 B.n665 B.n663 10.6151
R1688 B.n666 B.n665 10.6151
R1689 B.n667 B.n666 10.6151
R1690 B.n668 B.n667 10.6151
R1691 B.n670 B.n668 10.6151
R1692 B.n671 B.n670 10.6151
R1693 B.n672 B.n671 10.6151
R1694 B.n673 B.n672 10.6151
R1695 B.n675 B.n673 10.6151
R1696 B.n676 B.n675 10.6151
R1697 B.n677 B.n676 10.6151
R1698 B.n678 B.n677 10.6151
R1699 B.n680 B.n678 10.6151
R1700 B.n681 B.n680 10.6151
R1701 B.n682 B.n681 10.6151
R1702 B.n683 B.n682 10.6151
R1703 B.n685 B.n683 10.6151
R1704 B.n686 B.n685 10.6151
R1705 B.n687 B.n686 10.6151
R1706 B.n688 B.n687 10.6151
R1707 B.n690 B.n688 10.6151
R1708 B.n691 B.n690 10.6151
R1709 B.n692 B.n691 10.6151
R1710 B.n693 B.n692 10.6151
R1711 B.n695 B.n693 10.6151
R1712 B.n696 B.n695 10.6151
R1713 B.n697 B.n696 10.6151
R1714 B.n698 B.n697 10.6151
R1715 B.n700 B.n698 10.6151
R1716 B.n701 B.n700 10.6151
R1717 B.n702 B.n701 10.6151
R1718 B.n703 B.n702 10.6151
R1719 B.n705 B.n703 10.6151
R1720 B.n706 B.n705 10.6151
R1721 B.n707 B.n706 10.6151
R1722 B.n708 B.n707 10.6151
R1723 B.n710 B.n708 10.6151
R1724 B.n711 B.n710 10.6151
R1725 B.n712 B.n711 10.6151
R1726 B.n713 B.n712 10.6151
R1727 B.n715 B.n713 10.6151
R1728 B.n716 B.n715 10.6151
R1729 B.n717 B.n716 10.6151
R1730 B.n718 B.n717 10.6151
R1731 B.n720 B.n718 10.6151
R1732 B.n721 B.n720 10.6151
R1733 B.n722 B.n721 10.6151
R1734 B.n723 B.n722 10.6151
R1735 B.n725 B.n723 10.6151
R1736 B.n726 B.n725 10.6151
R1737 B.n727 B.n726 10.6151
R1738 B.n728 B.n727 10.6151
R1739 B.n730 B.n728 10.6151
R1740 B.n731 B.n730 10.6151
R1741 B.n732 B.n731 10.6151
R1742 B.n733 B.n732 10.6151
R1743 B.n450 B.n449 10.6151
R1744 B.n449 B.n289 10.6151
R1745 B.n444 B.n289 10.6151
R1746 B.n444 B.n443 10.6151
R1747 B.n443 B.n291 10.6151
R1748 B.n438 B.n291 10.6151
R1749 B.n438 B.n437 10.6151
R1750 B.n437 B.n436 10.6151
R1751 B.n436 B.n293 10.6151
R1752 B.n430 B.n293 10.6151
R1753 B.n430 B.n429 10.6151
R1754 B.n429 B.n428 10.6151
R1755 B.n428 B.n295 10.6151
R1756 B.n422 B.n295 10.6151
R1757 B.n422 B.n421 10.6151
R1758 B.n421 B.n420 10.6151
R1759 B.n420 B.n297 10.6151
R1760 B.n414 B.n297 10.6151
R1761 B.n414 B.n413 10.6151
R1762 B.n413 B.n412 10.6151
R1763 B.n412 B.n299 10.6151
R1764 B.n406 B.n299 10.6151
R1765 B.n406 B.n405 10.6151
R1766 B.n405 B.n404 10.6151
R1767 B.n404 B.n301 10.6151
R1768 B.n398 B.n301 10.6151
R1769 B.n396 B.n395 10.6151
R1770 B.n395 B.n305 10.6151
R1771 B.n389 B.n305 10.6151
R1772 B.n389 B.n388 10.6151
R1773 B.n388 B.n387 10.6151
R1774 B.n387 B.n307 10.6151
R1775 B.n381 B.n307 10.6151
R1776 B.n381 B.n380 10.6151
R1777 B.n380 B.n379 10.6151
R1778 B.n375 B.n374 10.6151
R1779 B.n374 B.n313 10.6151
R1780 B.n369 B.n313 10.6151
R1781 B.n369 B.n368 10.6151
R1782 B.n368 B.n367 10.6151
R1783 B.n367 B.n315 10.6151
R1784 B.n361 B.n315 10.6151
R1785 B.n361 B.n360 10.6151
R1786 B.n360 B.n359 10.6151
R1787 B.n359 B.n317 10.6151
R1788 B.n353 B.n317 10.6151
R1789 B.n353 B.n352 10.6151
R1790 B.n352 B.n351 10.6151
R1791 B.n351 B.n319 10.6151
R1792 B.n345 B.n319 10.6151
R1793 B.n345 B.n344 10.6151
R1794 B.n344 B.n343 10.6151
R1795 B.n343 B.n321 10.6151
R1796 B.n337 B.n321 10.6151
R1797 B.n337 B.n336 10.6151
R1798 B.n336 B.n335 10.6151
R1799 B.n335 B.n323 10.6151
R1800 B.n329 B.n323 10.6151
R1801 B.n329 B.n328 10.6151
R1802 B.n328 B.n327 10.6151
R1803 B.n327 B.n285 10.6151
R1804 B.n451 B.n281 10.6151
R1805 B.n461 B.n281 10.6151
R1806 B.n462 B.n461 10.6151
R1807 B.n463 B.n462 10.6151
R1808 B.n463 B.n273 10.6151
R1809 B.n473 B.n273 10.6151
R1810 B.n474 B.n473 10.6151
R1811 B.n475 B.n474 10.6151
R1812 B.n475 B.n265 10.6151
R1813 B.n485 B.n265 10.6151
R1814 B.n486 B.n485 10.6151
R1815 B.n487 B.n486 10.6151
R1816 B.n487 B.n257 10.6151
R1817 B.n497 B.n257 10.6151
R1818 B.n498 B.n497 10.6151
R1819 B.n499 B.n498 10.6151
R1820 B.n499 B.n249 10.6151
R1821 B.n509 B.n249 10.6151
R1822 B.n510 B.n509 10.6151
R1823 B.n511 B.n510 10.6151
R1824 B.n511 B.n241 10.6151
R1825 B.n521 B.n241 10.6151
R1826 B.n522 B.n521 10.6151
R1827 B.n523 B.n522 10.6151
R1828 B.n523 B.n233 10.6151
R1829 B.n533 B.n233 10.6151
R1830 B.n534 B.n533 10.6151
R1831 B.n535 B.n534 10.6151
R1832 B.n535 B.n225 10.6151
R1833 B.n545 B.n225 10.6151
R1834 B.n546 B.n545 10.6151
R1835 B.n547 B.n546 10.6151
R1836 B.n547 B.n217 10.6151
R1837 B.n557 B.n217 10.6151
R1838 B.n558 B.n557 10.6151
R1839 B.n559 B.n558 10.6151
R1840 B.n559 B.n209 10.6151
R1841 B.n569 B.n209 10.6151
R1842 B.n570 B.n569 10.6151
R1843 B.n571 B.n570 10.6151
R1844 B.n571 B.n201 10.6151
R1845 B.n581 B.n201 10.6151
R1846 B.n582 B.n581 10.6151
R1847 B.n583 B.n582 10.6151
R1848 B.n583 B.n193 10.6151
R1849 B.n593 B.n193 10.6151
R1850 B.n594 B.n593 10.6151
R1851 B.n595 B.n594 10.6151
R1852 B.n595 B.n185 10.6151
R1853 B.n605 B.n185 10.6151
R1854 B.n606 B.n605 10.6151
R1855 B.n607 B.n606 10.6151
R1856 B.n607 B.n177 10.6151
R1857 B.n617 B.n177 10.6151
R1858 B.n618 B.n617 10.6151
R1859 B.n619 B.n618 10.6151
R1860 B.n619 B.n169 10.6151
R1861 B.n630 B.n169 10.6151
R1862 B.n631 B.n630 10.6151
R1863 B.n632 B.n631 10.6151
R1864 B.n632 B.n162 10.6151
R1865 B.n643 B.n162 10.6151
R1866 B.n644 B.n643 10.6151
R1867 B.n645 B.n644 10.6151
R1868 B.n645 B.n0 10.6151
R1869 B.n991 B.n1 10.6151
R1870 B.n991 B.n990 10.6151
R1871 B.n990 B.n989 10.6151
R1872 B.n989 B.n10 10.6151
R1873 B.n983 B.n10 10.6151
R1874 B.n983 B.n982 10.6151
R1875 B.n982 B.n981 10.6151
R1876 B.n981 B.n16 10.6151
R1877 B.n975 B.n16 10.6151
R1878 B.n975 B.n974 10.6151
R1879 B.n974 B.n973 10.6151
R1880 B.n973 B.n24 10.6151
R1881 B.n967 B.n24 10.6151
R1882 B.n967 B.n966 10.6151
R1883 B.n966 B.n965 10.6151
R1884 B.n965 B.n31 10.6151
R1885 B.n959 B.n31 10.6151
R1886 B.n959 B.n958 10.6151
R1887 B.n958 B.n957 10.6151
R1888 B.n957 B.n38 10.6151
R1889 B.n951 B.n38 10.6151
R1890 B.n951 B.n950 10.6151
R1891 B.n950 B.n949 10.6151
R1892 B.n949 B.n45 10.6151
R1893 B.n943 B.n45 10.6151
R1894 B.n943 B.n942 10.6151
R1895 B.n942 B.n941 10.6151
R1896 B.n941 B.n52 10.6151
R1897 B.n935 B.n52 10.6151
R1898 B.n935 B.n934 10.6151
R1899 B.n934 B.n933 10.6151
R1900 B.n933 B.n59 10.6151
R1901 B.n927 B.n59 10.6151
R1902 B.n927 B.n926 10.6151
R1903 B.n926 B.n925 10.6151
R1904 B.n925 B.n66 10.6151
R1905 B.n919 B.n66 10.6151
R1906 B.n919 B.n918 10.6151
R1907 B.n918 B.n917 10.6151
R1908 B.n917 B.n73 10.6151
R1909 B.n911 B.n73 10.6151
R1910 B.n911 B.n910 10.6151
R1911 B.n910 B.n909 10.6151
R1912 B.n909 B.n80 10.6151
R1913 B.n903 B.n80 10.6151
R1914 B.n903 B.n902 10.6151
R1915 B.n902 B.n901 10.6151
R1916 B.n901 B.n87 10.6151
R1917 B.n895 B.n87 10.6151
R1918 B.n895 B.n894 10.6151
R1919 B.n894 B.n893 10.6151
R1920 B.n893 B.n94 10.6151
R1921 B.n887 B.n94 10.6151
R1922 B.n887 B.n886 10.6151
R1923 B.n886 B.n885 10.6151
R1924 B.n885 B.n101 10.6151
R1925 B.n879 B.n101 10.6151
R1926 B.n879 B.n878 10.6151
R1927 B.n878 B.n877 10.6151
R1928 B.n877 B.n108 10.6151
R1929 B.n871 B.n108 10.6151
R1930 B.n871 B.n870 10.6151
R1931 B.n870 B.n869 10.6151
R1932 B.n869 B.n115 10.6151
R1933 B.n863 B.n115 10.6151
R1934 B.n138 B.n134 9.36635
R1935 B.n789 B.n788 9.36635
R1936 B.n398 B.n397 9.36635
R1937 B.n375 B.n311 9.36635
R1938 B.n247 B.t5 7.14046
R1939 B.t23 B.n906 7.14046
R1940 B.n997 B.n0 2.81026
R1941 B.n997 B.n1 2.81026
R1942 B.n603 B.t1 1.78549
R1943 B.n963 B.t3 1.78549
R1944 B.n807 B.n138 1.24928
R1945 B.n790 B.n789 1.24928
R1946 B.n397 B.n396 1.24928
R1947 B.n379 B.n311 1.24928
R1948 VP.n27 VP.n26 161.3
R1949 VP.n28 VP.n23 161.3
R1950 VP.n30 VP.n29 161.3
R1951 VP.n31 VP.n22 161.3
R1952 VP.n33 VP.n32 161.3
R1953 VP.n34 VP.n21 161.3
R1954 VP.n36 VP.n35 161.3
R1955 VP.n37 VP.n20 161.3
R1956 VP.n39 VP.n38 161.3
R1957 VP.n40 VP.n19 161.3
R1958 VP.n42 VP.n41 161.3
R1959 VP.n43 VP.n18 161.3
R1960 VP.n46 VP.n45 161.3
R1961 VP.n47 VP.n17 161.3
R1962 VP.n49 VP.n48 161.3
R1963 VP.n50 VP.n16 161.3
R1964 VP.n52 VP.n51 161.3
R1965 VP.n53 VP.n15 161.3
R1966 VP.n55 VP.n54 161.3
R1967 VP.n56 VP.n14 161.3
R1968 VP.n102 VP.n0 161.3
R1969 VP.n101 VP.n100 161.3
R1970 VP.n99 VP.n1 161.3
R1971 VP.n98 VP.n97 161.3
R1972 VP.n96 VP.n2 161.3
R1973 VP.n95 VP.n94 161.3
R1974 VP.n93 VP.n3 161.3
R1975 VP.n92 VP.n91 161.3
R1976 VP.n89 VP.n4 161.3
R1977 VP.n88 VP.n87 161.3
R1978 VP.n86 VP.n5 161.3
R1979 VP.n85 VP.n84 161.3
R1980 VP.n83 VP.n6 161.3
R1981 VP.n82 VP.n81 161.3
R1982 VP.n80 VP.n7 161.3
R1983 VP.n79 VP.n78 161.3
R1984 VP.n77 VP.n8 161.3
R1985 VP.n76 VP.n75 161.3
R1986 VP.n74 VP.n9 161.3
R1987 VP.n73 VP.n72 161.3
R1988 VP.n70 VP.n10 161.3
R1989 VP.n69 VP.n68 161.3
R1990 VP.n67 VP.n11 161.3
R1991 VP.n66 VP.n65 161.3
R1992 VP.n64 VP.n12 161.3
R1993 VP.n63 VP.n62 161.3
R1994 VP.n61 VP.n13 161.3
R1995 VP.n60 VP.n59 108.799
R1996 VP.n104 VP.n103 108.799
R1997 VP.n58 VP.n57 108.799
R1998 VP.n24 VP.t8 90.4745
R1999 VP.n25 VP.n24 60.6237
R2000 VP.n82 VP.t2 57.7913
R2001 VP.n59 VP.t7 57.7913
R2002 VP.n71 VP.t6 57.7913
R2003 VP.n90 VP.t4 57.7913
R2004 VP.n103 VP.t3 57.7913
R2005 VP.n36 VP.t9 57.7913
R2006 VP.n57 VP.t0 57.7913
R2007 VP.n44 VP.t5 57.7913
R2008 VP.n25 VP.t1 57.7913
R2009 VP.n77 VP.n76 53.6055
R2010 VP.n88 VP.n5 53.6055
R2011 VP.n42 VP.n19 53.6055
R2012 VP.n31 VP.n30 53.6055
R2013 VP.n60 VP.n58 51.1928
R2014 VP.n65 VP.n11 49.7204
R2015 VP.n97 VP.n96 49.7204
R2016 VP.n51 VP.n50 49.7204
R2017 VP.n65 VP.n64 31.2664
R2018 VP.n97 VP.n1 31.2664
R2019 VP.n51 VP.n15 31.2664
R2020 VP.n78 VP.n77 27.3813
R2021 VP.n84 VP.n5 27.3813
R2022 VP.n38 VP.n19 27.3813
R2023 VP.n32 VP.n31 27.3813
R2024 VP.n63 VP.n13 24.4675
R2025 VP.n64 VP.n63 24.4675
R2026 VP.n69 VP.n11 24.4675
R2027 VP.n70 VP.n69 24.4675
R2028 VP.n72 VP.n9 24.4675
R2029 VP.n76 VP.n9 24.4675
R2030 VP.n78 VP.n7 24.4675
R2031 VP.n82 VP.n7 24.4675
R2032 VP.n83 VP.n82 24.4675
R2033 VP.n84 VP.n83 24.4675
R2034 VP.n89 VP.n88 24.4675
R2035 VP.n91 VP.n89 24.4675
R2036 VP.n95 VP.n3 24.4675
R2037 VP.n96 VP.n95 24.4675
R2038 VP.n101 VP.n1 24.4675
R2039 VP.n102 VP.n101 24.4675
R2040 VP.n55 VP.n15 24.4675
R2041 VP.n56 VP.n55 24.4675
R2042 VP.n43 VP.n42 24.4675
R2043 VP.n45 VP.n43 24.4675
R2044 VP.n49 VP.n17 24.4675
R2045 VP.n50 VP.n49 24.4675
R2046 VP.n32 VP.n21 24.4675
R2047 VP.n36 VP.n21 24.4675
R2048 VP.n37 VP.n36 24.4675
R2049 VP.n38 VP.n37 24.4675
R2050 VP.n26 VP.n23 24.4675
R2051 VP.n30 VP.n23 24.4675
R2052 VP.n72 VP.n71 13.2127
R2053 VP.n91 VP.n90 13.2127
R2054 VP.n45 VP.n44 13.2127
R2055 VP.n26 VP.n25 13.2127
R2056 VP.n71 VP.n70 11.2553
R2057 VP.n90 VP.n3 11.2553
R2058 VP.n44 VP.n17 11.2553
R2059 VP.n27 VP.n24 5.12434
R2060 VP.n59 VP.n13 1.95786
R2061 VP.n103 VP.n102 1.95786
R2062 VP.n57 VP.n56 1.95786
R2063 VP.n58 VP.n14 0.278367
R2064 VP.n61 VP.n60 0.278367
R2065 VP.n104 VP.n0 0.278367
R2066 VP.n28 VP.n27 0.189894
R2067 VP.n29 VP.n28 0.189894
R2068 VP.n29 VP.n22 0.189894
R2069 VP.n33 VP.n22 0.189894
R2070 VP.n34 VP.n33 0.189894
R2071 VP.n35 VP.n34 0.189894
R2072 VP.n35 VP.n20 0.189894
R2073 VP.n39 VP.n20 0.189894
R2074 VP.n40 VP.n39 0.189894
R2075 VP.n41 VP.n40 0.189894
R2076 VP.n41 VP.n18 0.189894
R2077 VP.n46 VP.n18 0.189894
R2078 VP.n47 VP.n46 0.189894
R2079 VP.n48 VP.n47 0.189894
R2080 VP.n48 VP.n16 0.189894
R2081 VP.n52 VP.n16 0.189894
R2082 VP.n53 VP.n52 0.189894
R2083 VP.n54 VP.n53 0.189894
R2084 VP.n54 VP.n14 0.189894
R2085 VP.n62 VP.n61 0.189894
R2086 VP.n62 VP.n12 0.189894
R2087 VP.n66 VP.n12 0.189894
R2088 VP.n67 VP.n66 0.189894
R2089 VP.n68 VP.n67 0.189894
R2090 VP.n68 VP.n10 0.189894
R2091 VP.n73 VP.n10 0.189894
R2092 VP.n74 VP.n73 0.189894
R2093 VP.n75 VP.n74 0.189894
R2094 VP.n75 VP.n8 0.189894
R2095 VP.n79 VP.n8 0.189894
R2096 VP.n80 VP.n79 0.189894
R2097 VP.n81 VP.n80 0.189894
R2098 VP.n81 VP.n6 0.189894
R2099 VP.n85 VP.n6 0.189894
R2100 VP.n86 VP.n85 0.189894
R2101 VP.n87 VP.n86 0.189894
R2102 VP.n87 VP.n4 0.189894
R2103 VP.n92 VP.n4 0.189894
R2104 VP.n93 VP.n92 0.189894
R2105 VP.n94 VP.n93 0.189894
R2106 VP.n94 VP.n2 0.189894
R2107 VP.n98 VP.n2 0.189894
R2108 VP.n99 VP.n98 0.189894
R2109 VP.n100 VP.n99 0.189894
R2110 VP.n100 VP.n0 0.189894
R2111 VP VP.n104 0.153454
R2112 VDD1.n1 VDD1.t1 70.6569
R2113 VDD1.n3 VDD1.t2 70.6567
R2114 VDD1.n5 VDD1.n4 67.0882
R2115 VDD1.n1 VDD1.n0 65.0294
R2116 VDD1.n3 VDD1.n2 65.0294
R2117 VDD1.n7 VDD1.n6 65.0292
R2118 VDD1.n7 VDD1.n5 45.1755
R2119 VDD1.n6 VDD1.t4 2.80901
R2120 VDD1.n6 VDD1.t9 2.80901
R2121 VDD1.n0 VDD1.t8 2.80901
R2122 VDD1.n0 VDD1.t0 2.80901
R2123 VDD1.n4 VDD1.t5 2.80901
R2124 VDD1.n4 VDD1.t6 2.80901
R2125 VDD1.n2 VDD1.t3 2.80901
R2126 VDD1.n2 VDD1.t7 2.80901
R2127 VDD1 VDD1.n7 2.05653
R2128 VDD1 VDD1.n1 0.763431
R2129 VDD1.n5 VDD1.n3 0.649895
C0 VDD1 VTAIL 8.34786f
C1 VTAIL VP 7.87527f
C2 VTAIL VDD2 8.402441f
C3 VTAIL VN 7.86107f
C4 VDD1 VP 7.09959f
C5 VDD1 VDD2 2.39509f
C6 VDD1 VN 0.154108f
C7 VP VDD2 0.626564f
C8 VN VP 7.9819f
C9 VN VDD2 6.63021f
C10 VDD2 B 6.784275f
C11 VDD1 B 6.715201f
C12 VTAIL B 6.009384f
C13 VN B 19.153109f
C14 VP B 17.722136f
C15 VDD1.t1 B 1.60201f
C16 VDD1.t8 B 0.146446f
C17 VDD1.t0 B 0.146446f
C18 VDD1.n0 B 1.24349f
C19 VDD1.n1 B 1.02734f
C20 VDD1.t2 B 1.60201f
C21 VDD1.t3 B 0.146446f
C22 VDD1.t7 B 0.146446f
C23 VDD1.n2 B 1.24349f
C24 VDD1.n3 B 1.01867f
C25 VDD1.t5 B 0.146446f
C26 VDD1.t6 B 0.146446f
C27 VDD1.n4 B 1.26316f
C28 VDD1.n5 B 3.06044f
C29 VDD1.t4 B 0.146446f
C30 VDD1.t9 B 0.146446f
C31 VDD1.n6 B 1.24349f
C32 VDD1.n7 B 3.08556f
C33 VP.n0 B 0.029347f
C34 VP.t3 B 1.23186f
C35 VP.n1 B 0.044693f
C36 VP.n2 B 0.02226f
C37 VP.n3 B 0.030426f
C38 VP.n4 B 0.02226f
C39 VP.n5 B 0.023816f
C40 VP.n6 B 0.02226f
C41 VP.t2 B 1.23186f
C42 VP.n7 B 0.041486f
C43 VP.n8 B 0.02226f
C44 VP.n9 B 0.041486f
C45 VP.n10 B 0.02226f
C46 VP.t6 B 1.23186f
C47 VP.n11 B 0.04107f
C48 VP.n12 B 0.02226f
C49 VP.n13 B 0.022643f
C50 VP.n14 B 0.029347f
C51 VP.t0 B 1.23186f
C52 VP.n15 B 0.044693f
C53 VP.n16 B 0.02226f
C54 VP.n17 B 0.030426f
C55 VP.n18 B 0.02226f
C56 VP.n19 B 0.023816f
C57 VP.n20 B 0.02226f
C58 VP.t9 B 1.23186f
C59 VP.n21 B 0.041486f
C60 VP.n22 B 0.02226f
C61 VP.n23 B 0.041486f
C62 VP.t8 B 1.4501f
C63 VP.n24 B 0.500199f
C64 VP.t1 B 1.23186f
C65 VP.n25 B 0.522285f
C66 VP.n26 B 0.032065f
C67 VP.n27 B 0.237124f
C68 VP.n28 B 0.02226f
C69 VP.n29 B 0.02226f
C70 VP.n30 B 0.03926f
C71 VP.n31 B 0.023816f
C72 VP.n32 B 0.043405f
C73 VP.n33 B 0.02226f
C74 VP.n34 B 0.02226f
C75 VP.n35 B 0.02226f
C76 VP.n36 B 0.472484f
C77 VP.n37 B 0.041486f
C78 VP.n38 B 0.043405f
C79 VP.n39 B 0.02226f
C80 VP.n40 B 0.02226f
C81 VP.n41 B 0.02226f
C82 VP.n42 B 0.03926f
C83 VP.n43 B 0.041486f
C84 VP.t5 B 1.23186f
C85 VP.n44 B 0.45148f
C86 VP.n45 B 0.032065f
C87 VP.n46 B 0.02226f
C88 VP.n47 B 0.02226f
C89 VP.n48 B 0.02226f
C90 VP.n49 B 0.041486f
C91 VP.n50 B 0.04107f
C92 VP.n51 B 0.020717f
C93 VP.n52 B 0.02226f
C94 VP.n53 B 0.02226f
C95 VP.n54 B 0.02226f
C96 VP.n55 B 0.041486f
C97 VP.n56 B 0.022643f
C98 VP.n57 B 0.526322f
C99 VP.n58 B 1.28918f
C100 VP.t7 B 1.23186f
C101 VP.n59 B 0.526322f
C102 VP.n60 B 1.30481f
C103 VP.n61 B 0.029347f
C104 VP.n62 B 0.02226f
C105 VP.n63 B 0.041486f
C106 VP.n64 B 0.044693f
C107 VP.n65 B 0.020717f
C108 VP.n66 B 0.02226f
C109 VP.n67 B 0.02226f
C110 VP.n68 B 0.02226f
C111 VP.n69 B 0.041486f
C112 VP.n70 B 0.030426f
C113 VP.n71 B 0.45148f
C114 VP.n72 B 0.032065f
C115 VP.n73 B 0.02226f
C116 VP.n74 B 0.02226f
C117 VP.n75 B 0.02226f
C118 VP.n76 B 0.03926f
C119 VP.n77 B 0.023816f
C120 VP.n78 B 0.043405f
C121 VP.n79 B 0.02226f
C122 VP.n80 B 0.02226f
C123 VP.n81 B 0.02226f
C124 VP.n82 B 0.472484f
C125 VP.n83 B 0.041486f
C126 VP.n84 B 0.043405f
C127 VP.n85 B 0.02226f
C128 VP.n86 B 0.02226f
C129 VP.n87 B 0.02226f
C130 VP.n88 B 0.03926f
C131 VP.n89 B 0.041486f
C132 VP.t4 B 1.23186f
C133 VP.n90 B 0.45148f
C134 VP.n91 B 0.032065f
C135 VP.n92 B 0.02226f
C136 VP.n93 B 0.02226f
C137 VP.n94 B 0.02226f
C138 VP.n95 B 0.041486f
C139 VP.n96 B 0.04107f
C140 VP.n97 B 0.020717f
C141 VP.n98 B 0.02226f
C142 VP.n99 B 0.02226f
C143 VP.n100 B 0.02226f
C144 VP.n101 B 0.041486f
C145 VP.n102 B 0.022643f
C146 VP.n103 B 0.526322f
C147 VP.n104 B 0.043228f
C148 VTAIL.t16 B 0.156495f
C149 VTAIL.t9 B 0.156495f
C150 VTAIL.n0 B 1.25072f
C151 VTAIL.n1 B 0.638382f
C152 VTAIL.t0 B 1.59402f
C153 VTAIL.n2 B 0.78041f
C154 VTAIL.t2 B 0.156495f
C155 VTAIL.t1 B 0.156495f
C156 VTAIL.n3 B 1.25072f
C157 VTAIL.n4 B 0.781955f
C158 VTAIL.t5 B 0.156495f
C159 VTAIL.t6 B 0.156495f
C160 VTAIL.n5 B 1.25072f
C161 VTAIL.n6 B 1.96878f
C162 VTAIL.t12 B 0.156495f
C163 VTAIL.t10 B 0.156495f
C164 VTAIL.n7 B 1.25072f
C165 VTAIL.n8 B 1.96878f
C166 VTAIL.t17 B 0.156495f
C167 VTAIL.t14 B 0.156495f
C168 VTAIL.n9 B 1.25072f
C169 VTAIL.n10 B 0.781953f
C170 VTAIL.t11 B 1.59402f
C171 VTAIL.n11 B 0.780403f
C172 VTAIL.t7 B 0.156495f
C173 VTAIL.t3 B 0.156495f
C174 VTAIL.n12 B 1.25072f
C175 VTAIL.n13 B 0.696901f
C176 VTAIL.t8 B 0.156495f
C177 VTAIL.t4 B 0.156495f
C178 VTAIL.n14 B 1.25072f
C179 VTAIL.n15 B 0.781953f
C180 VTAIL.t19 B 1.59401f
C181 VTAIL.n16 B 1.79714f
C182 VTAIL.t13 B 1.59402f
C183 VTAIL.n17 B 1.79714f
C184 VTAIL.t15 B 0.156495f
C185 VTAIL.t18 B 0.156495f
C186 VTAIL.n18 B 1.25072f
C187 VTAIL.n19 B 0.585323f
C188 VDD2.t8 B 1.57459f
C189 VDD2.t6 B 0.14394f
C190 VDD2.t1 B 0.14394f
C191 VDD2.n0 B 1.22221f
C192 VDD2.n1 B 1.00124f
C193 VDD2.t5 B 0.14394f
C194 VDD2.t9 B 0.14394f
C195 VDD2.n2 B 1.24155f
C196 VDD2.n3 B 2.87354f
C197 VDD2.t2 B 1.55389f
C198 VDD2.n4 B 2.96159f
C199 VDD2.t7 B 0.14394f
C200 VDD2.t4 B 0.14394f
C201 VDD2.n5 B 1.22222f
C202 VDD2.n6 B 0.511344f
C203 VDD2.t3 B 0.14394f
C204 VDD2.t0 B 0.14394f
C205 VDD2.n7 B 1.2415f
C206 VN.n0 B 0.02867f
C207 VN.t5 B 1.20344f
C208 VN.n1 B 0.043662f
C209 VN.n2 B 0.021746f
C210 VN.n3 B 0.029724f
C211 VN.n4 B 0.021746f
C212 VN.n5 B 0.023267f
C213 VN.n6 B 0.021746f
C214 VN.t3 B 1.20344f
C215 VN.n7 B 0.040529f
C216 VN.n8 B 0.021746f
C217 VN.n9 B 0.040529f
C218 VN.t2 B 1.41665f
C219 VN.n10 B 0.48866f
C220 VN.t9 B 1.20344f
C221 VN.n11 B 0.510237f
C222 VN.n12 B 0.031325f
C223 VN.n13 B 0.231654f
C224 VN.n14 B 0.021746f
C225 VN.n15 B 0.021746f
C226 VN.n16 B 0.038354f
C227 VN.n17 B 0.023267f
C228 VN.n18 B 0.042403f
C229 VN.n19 B 0.021746f
C230 VN.n20 B 0.021746f
C231 VN.n21 B 0.021746f
C232 VN.n22 B 0.461585f
C233 VN.n23 B 0.040529f
C234 VN.n24 B 0.042403f
C235 VN.n25 B 0.021746f
C236 VN.n26 B 0.021746f
C237 VN.n27 B 0.021746f
C238 VN.n28 B 0.038354f
C239 VN.n29 B 0.040529f
C240 VN.t0 B 1.20344f
C241 VN.n30 B 0.441065f
C242 VN.n31 B 0.031325f
C243 VN.n32 B 0.021746f
C244 VN.n33 B 0.021746f
C245 VN.n34 B 0.021746f
C246 VN.n35 B 0.040529f
C247 VN.n36 B 0.040123f
C248 VN.n37 B 0.020239f
C249 VN.n38 B 0.021746f
C250 VN.n39 B 0.021746f
C251 VN.n40 B 0.021746f
C252 VN.n41 B 0.040529f
C253 VN.n42 B 0.022121f
C254 VN.n43 B 0.514181f
C255 VN.n44 B 0.042231f
C256 VN.n45 B 0.02867f
C257 VN.t6 B 1.20344f
C258 VN.n46 B 0.043662f
C259 VN.n47 B 0.021746f
C260 VN.n48 B 0.029724f
C261 VN.n49 B 0.021746f
C262 VN.t8 B 1.20344f
C263 VN.n50 B 0.441065f
C264 VN.n51 B 0.023267f
C265 VN.n52 B 0.021746f
C266 VN.t1 B 1.20344f
C267 VN.n53 B 0.040529f
C268 VN.n54 B 0.021746f
C269 VN.n55 B 0.040529f
C270 VN.t7 B 1.41665f
C271 VN.n56 B 0.48866f
C272 VN.t4 B 1.20344f
C273 VN.n57 B 0.510237f
C274 VN.n58 B 0.031325f
C275 VN.n59 B 0.231654f
C276 VN.n60 B 0.021746f
C277 VN.n61 B 0.021746f
C278 VN.n62 B 0.038354f
C279 VN.n63 B 0.023267f
C280 VN.n64 B 0.042403f
C281 VN.n65 B 0.021746f
C282 VN.n66 B 0.021746f
C283 VN.n67 B 0.021746f
C284 VN.n68 B 0.461585f
C285 VN.n69 B 0.040529f
C286 VN.n70 B 0.042403f
C287 VN.n71 B 0.021746f
C288 VN.n72 B 0.021746f
C289 VN.n73 B 0.021746f
C290 VN.n74 B 0.038354f
C291 VN.n75 B 0.040529f
C292 VN.n76 B 0.031325f
C293 VN.n77 B 0.021746f
C294 VN.n78 B 0.021746f
C295 VN.n79 B 0.021746f
C296 VN.n80 B 0.040529f
C297 VN.n81 B 0.040123f
C298 VN.n82 B 0.020239f
C299 VN.n83 B 0.021746f
C300 VN.n84 B 0.021746f
C301 VN.n85 B 0.021746f
C302 VN.n86 B 0.040529f
C303 VN.n87 B 0.022121f
C304 VN.n88 B 0.514181f
C305 VN.n89 B 1.27108f
.ends

