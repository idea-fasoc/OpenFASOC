* NGSPICE file created from diff_pair_sample_1731.ext - technology: sky130A

.subckt diff_pair_sample_1731 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t3 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=1.53285 ps=9.62 w=9.29 l=3.93
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=0 ps=0 w=9.29 l=3.93
X2 VDD1.t3 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.53285 pd=9.62 as=3.6231 ps=19.36 w=9.29 l=3.93
X3 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=1.53285 ps=9.62 w=9.29 l=3.93
X4 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=1.53285 ps=9.62 w=9.29 l=3.93
X5 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=0 ps=0 w=9.29 l=3.93
X6 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=0 ps=0 w=9.29 l=3.93
X7 VDD2.t0 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53285 pd=9.62 as=3.6231 ps=19.36 w=9.29 l=3.93
X8 VDD2.t3 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.53285 pd=9.62 as=3.6231 ps=19.36 w=9.29 l=3.93
X9 VTAIL.t5 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=1.53285 ps=9.62 w=9.29 l=3.93
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.6231 pd=19.36 as=0 ps=0 w=9.29 l=3.93
X11 VDD1.t0 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53285 pd=9.62 as=3.6231 ps=19.36 w=9.29 l=3.93
R0 VN.n0 VN.t0 90.7955
R1 VN.n1 VN.t2 90.7955
R2 VN.n0 VN.t3 89.3683
R3 VN.n1 VN.t1 89.3683
R4 VN VN.n1 50.2447
R5 VN VN.n0 1.78636
R6 VDD2.n2 VDD2.n0 106.713
R7 VDD2.n2 VDD2.n1 63.9716
R8 VDD2.n1 VDD2.t2 2.13182
R9 VDD2.n1 VDD2.t0 2.13182
R10 VDD2.n0 VDD2.t1 2.13182
R11 VDD2.n0 VDD2.t3 2.13182
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n394 VTAIL.n350 289.615
R14 VTAIL.n44 VTAIL.n0 289.615
R15 VTAIL.n94 VTAIL.n50 289.615
R16 VTAIL.n144 VTAIL.n100 289.615
R17 VTAIL.n344 VTAIL.n300 289.615
R18 VTAIL.n294 VTAIL.n250 289.615
R19 VTAIL.n244 VTAIL.n200 289.615
R20 VTAIL.n194 VTAIL.n150 289.615
R21 VTAIL.n367 VTAIL.n366 185
R22 VTAIL.n369 VTAIL.n368 185
R23 VTAIL.n362 VTAIL.n361 185
R24 VTAIL.n375 VTAIL.n374 185
R25 VTAIL.n377 VTAIL.n376 185
R26 VTAIL.n358 VTAIL.n357 185
R27 VTAIL.n384 VTAIL.n383 185
R28 VTAIL.n385 VTAIL.n356 185
R29 VTAIL.n387 VTAIL.n386 185
R30 VTAIL.n354 VTAIL.n353 185
R31 VTAIL.n393 VTAIL.n392 185
R32 VTAIL.n395 VTAIL.n394 185
R33 VTAIL.n17 VTAIL.n16 185
R34 VTAIL.n19 VTAIL.n18 185
R35 VTAIL.n12 VTAIL.n11 185
R36 VTAIL.n25 VTAIL.n24 185
R37 VTAIL.n27 VTAIL.n26 185
R38 VTAIL.n8 VTAIL.n7 185
R39 VTAIL.n34 VTAIL.n33 185
R40 VTAIL.n35 VTAIL.n6 185
R41 VTAIL.n37 VTAIL.n36 185
R42 VTAIL.n4 VTAIL.n3 185
R43 VTAIL.n43 VTAIL.n42 185
R44 VTAIL.n45 VTAIL.n44 185
R45 VTAIL.n67 VTAIL.n66 185
R46 VTAIL.n69 VTAIL.n68 185
R47 VTAIL.n62 VTAIL.n61 185
R48 VTAIL.n75 VTAIL.n74 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n58 VTAIL.n57 185
R51 VTAIL.n84 VTAIL.n83 185
R52 VTAIL.n85 VTAIL.n56 185
R53 VTAIL.n87 VTAIL.n86 185
R54 VTAIL.n54 VTAIL.n53 185
R55 VTAIL.n93 VTAIL.n92 185
R56 VTAIL.n95 VTAIL.n94 185
R57 VTAIL.n117 VTAIL.n116 185
R58 VTAIL.n119 VTAIL.n118 185
R59 VTAIL.n112 VTAIL.n111 185
R60 VTAIL.n125 VTAIL.n124 185
R61 VTAIL.n127 VTAIL.n126 185
R62 VTAIL.n108 VTAIL.n107 185
R63 VTAIL.n134 VTAIL.n133 185
R64 VTAIL.n135 VTAIL.n106 185
R65 VTAIL.n137 VTAIL.n136 185
R66 VTAIL.n104 VTAIL.n103 185
R67 VTAIL.n143 VTAIL.n142 185
R68 VTAIL.n145 VTAIL.n144 185
R69 VTAIL.n345 VTAIL.n344 185
R70 VTAIL.n343 VTAIL.n342 185
R71 VTAIL.n304 VTAIL.n303 185
R72 VTAIL.n308 VTAIL.n306 185
R73 VTAIL.n337 VTAIL.n336 185
R74 VTAIL.n335 VTAIL.n334 185
R75 VTAIL.n310 VTAIL.n309 185
R76 VTAIL.n329 VTAIL.n328 185
R77 VTAIL.n327 VTAIL.n326 185
R78 VTAIL.n314 VTAIL.n313 185
R79 VTAIL.n321 VTAIL.n320 185
R80 VTAIL.n319 VTAIL.n318 185
R81 VTAIL.n295 VTAIL.n294 185
R82 VTAIL.n293 VTAIL.n292 185
R83 VTAIL.n254 VTAIL.n253 185
R84 VTAIL.n258 VTAIL.n256 185
R85 VTAIL.n287 VTAIL.n286 185
R86 VTAIL.n285 VTAIL.n284 185
R87 VTAIL.n260 VTAIL.n259 185
R88 VTAIL.n279 VTAIL.n278 185
R89 VTAIL.n277 VTAIL.n276 185
R90 VTAIL.n264 VTAIL.n263 185
R91 VTAIL.n271 VTAIL.n270 185
R92 VTAIL.n269 VTAIL.n268 185
R93 VTAIL.n245 VTAIL.n244 185
R94 VTAIL.n243 VTAIL.n242 185
R95 VTAIL.n204 VTAIL.n203 185
R96 VTAIL.n208 VTAIL.n206 185
R97 VTAIL.n237 VTAIL.n236 185
R98 VTAIL.n235 VTAIL.n234 185
R99 VTAIL.n210 VTAIL.n209 185
R100 VTAIL.n229 VTAIL.n228 185
R101 VTAIL.n227 VTAIL.n226 185
R102 VTAIL.n214 VTAIL.n213 185
R103 VTAIL.n221 VTAIL.n220 185
R104 VTAIL.n219 VTAIL.n218 185
R105 VTAIL.n195 VTAIL.n194 185
R106 VTAIL.n193 VTAIL.n192 185
R107 VTAIL.n154 VTAIL.n153 185
R108 VTAIL.n158 VTAIL.n156 185
R109 VTAIL.n187 VTAIL.n186 185
R110 VTAIL.n185 VTAIL.n184 185
R111 VTAIL.n160 VTAIL.n159 185
R112 VTAIL.n179 VTAIL.n178 185
R113 VTAIL.n177 VTAIL.n176 185
R114 VTAIL.n164 VTAIL.n163 185
R115 VTAIL.n171 VTAIL.n170 185
R116 VTAIL.n169 VTAIL.n168 185
R117 VTAIL.n365 VTAIL.t0 149.524
R118 VTAIL.n15 VTAIL.t3 149.524
R119 VTAIL.n65 VTAIL.t4 149.524
R120 VTAIL.n115 VTAIL.t6 149.524
R121 VTAIL.n317 VTAIL.t7 149.524
R122 VTAIL.n267 VTAIL.t5 149.524
R123 VTAIL.n217 VTAIL.t1 149.524
R124 VTAIL.n167 VTAIL.t2 149.524
R125 VTAIL.n368 VTAIL.n367 104.615
R126 VTAIL.n368 VTAIL.n361 104.615
R127 VTAIL.n375 VTAIL.n361 104.615
R128 VTAIL.n376 VTAIL.n375 104.615
R129 VTAIL.n376 VTAIL.n357 104.615
R130 VTAIL.n384 VTAIL.n357 104.615
R131 VTAIL.n385 VTAIL.n384 104.615
R132 VTAIL.n386 VTAIL.n385 104.615
R133 VTAIL.n386 VTAIL.n353 104.615
R134 VTAIL.n393 VTAIL.n353 104.615
R135 VTAIL.n394 VTAIL.n393 104.615
R136 VTAIL.n18 VTAIL.n17 104.615
R137 VTAIL.n18 VTAIL.n11 104.615
R138 VTAIL.n25 VTAIL.n11 104.615
R139 VTAIL.n26 VTAIL.n25 104.615
R140 VTAIL.n26 VTAIL.n7 104.615
R141 VTAIL.n34 VTAIL.n7 104.615
R142 VTAIL.n35 VTAIL.n34 104.615
R143 VTAIL.n36 VTAIL.n35 104.615
R144 VTAIL.n36 VTAIL.n3 104.615
R145 VTAIL.n43 VTAIL.n3 104.615
R146 VTAIL.n44 VTAIL.n43 104.615
R147 VTAIL.n68 VTAIL.n67 104.615
R148 VTAIL.n68 VTAIL.n61 104.615
R149 VTAIL.n75 VTAIL.n61 104.615
R150 VTAIL.n76 VTAIL.n75 104.615
R151 VTAIL.n76 VTAIL.n57 104.615
R152 VTAIL.n84 VTAIL.n57 104.615
R153 VTAIL.n85 VTAIL.n84 104.615
R154 VTAIL.n86 VTAIL.n85 104.615
R155 VTAIL.n86 VTAIL.n53 104.615
R156 VTAIL.n93 VTAIL.n53 104.615
R157 VTAIL.n94 VTAIL.n93 104.615
R158 VTAIL.n118 VTAIL.n117 104.615
R159 VTAIL.n118 VTAIL.n111 104.615
R160 VTAIL.n125 VTAIL.n111 104.615
R161 VTAIL.n126 VTAIL.n125 104.615
R162 VTAIL.n126 VTAIL.n107 104.615
R163 VTAIL.n134 VTAIL.n107 104.615
R164 VTAIL.n135 VTAIL.n134 104.615
R165 VTAIL.n136 VTAIL.n135 104.615
R166 VTAIL.n136 VTAIL.n103 104.615
R167 VTAIL.n143 VTAIL.n103 104.615
R168 VTAIL.n144 VTAIL.n143 104.615
R169 VTAIL.n344 VTAIL.n343 104.615
R170 VTAIL.n343 VTAIL.n303 104.615
R171 VTAIL.n308 VTAIL.n303 104.615
R172 VTAIL.n336 VTAIL.n308 104.615
R173 VTAIL.n336 VTAIL.n335 104.615
R174 VTAIL.n335 VTAIL.n309 104.615
R175 VTAIL.n328 VTAIL.n309 104.615
R176 VTAIL.n328 VTAIL.n327 104.615
R177 VTAIL.n327 VTAIL.n313 104.615
R178 VTAIL.n320 VTAIL.n313 104.615
R179 VTAIL.n320 VTAIL.n319 104.615
R180 VTAIL.n294 VTAIL.n293 104.615
R181 VTAIL.n293 VTAIL.n253 104.615
R182 VTAIL.n258 VTAIL.n253 104.615
R183 VTAIL.n286 VTAIL.n258 104.615
R184 VTAIL.n286 VTAIL.n285 104.615
R185 VTAIL.n285 VTAIL.n259 104.615
R186 VTAIL.n278 VTAIL.n259 104.615
R187 VTAIL.n278 VTAIL.n277 104.615
R188 VTAIL.n277 VTAIL.n263 104.615
R189 VTAIL.n270 VTAIL.n263 104.615
R190 VTAIL.n270 VTAIL.n269 104.615
R191 VTAIL.n244 VTAIL.n243 104.615
R192 VTAIL.n243 VTAIL.n203 104.615
R193 VTAIL.n208 VTAIL.n203 104.615
R194 VTAIL.n236 VTAIL.n208 104.615
R195 VTAIL.n236 VTAIL.n235 104.615
R196 VTAIL.n235 VTAIL.n209 104.615
R197 VTAIL.n228 VTAIL.n209 104.615
R198 VTAIL.n228 VTAIL.n227 104.615
R199 VTAIL.n227 VTAIL.n213 104.615
R200 VTAIL.n220 VTAIL.n213 104.615
R201 VTAIL.n220 VTAIL.n219 104.615
R202 VTAIL.n194 VTAIL.n193 104.615
R203 VTAIL.n193 VTAIL.n153 104.615
R204 VTAIL.n158 VTAIL.n153 104.615
R205 VTAIL.n186 VTAIL.n158 104.615
R206 VTAIL.n186 VTAIL.n185 104.615
R207 VTAIL.n185 VTAIL.n159 104.615
R208 VTAIL.n178 VTAIL.n159 104.615
R209 VTAIL.n178 VTAIL.n177 104.615
R210 VTAIL.n177 VTAIL.n163 104.615
R211 VTAIL.n170 VTAIL.n163 104.615
R212 VTAIL.n170 VTAIL.n169 104.615
R213 VTAIL.n367 VTAIL.t0 52.3082
R214 VTAIL.n17 VTAIL.t3 52.3082
R215 VTAIL.n67 VTAIL.t4 52.3082
R216 VTAIL.n117 VTAIL.t6 52.3082
R217 VTAIL.n319 VTAIL.t7 52.3082
R218 VTAIL.n269 VTAIL.t5 52.3082
R219 VTAIL.n219 VTAIL.t1 52.3082
R220 VTAIL.n169 VTAIL.t2 52.3082
R221 VTAIL.n399 VTAIL.n398 33.155
R222 VTAIL.n49 VTAIL.n48 33.155
R223 VTAIL.n99 VTAIL.n98 33.155
R224 VTAIL.n149 VTAIL.n148 33.155
R225 VTAIL.n349 VTAIL.n348 33.155
R226 VTAIL.n299 VTAIL.n298 33.155
R227 VTAIL.n249 VTAIL.n248 33.155
R228 VTAIL.n199 VTAIL.n198 33.155
R229 VTAIL.n399 VTAIL.n349 24.0479
R230 VTAIL.n199 VTAIL.n149 24.0479
R231 VTAIL.n387 VTAIL.n354 13.1884
R232 VTAIL.n37 VTAIL.n4 13.1884
R233 VTAIL.n87 VTAIL.n54 13.1884
R234 VTAIL.n137 VTAIL.n104 13.1884
R235 VTAIL.n306 VTAIL.n304 13.1884
R236 VTAIL.n256 VTAIL.n254 13.1884
R237 VTAIL.n206 VTAIL.n204 13.1884
R238 VTAIL.n156 VTAIL.n154 13.1884
R239 VTAIL.n388 VTAIL.n356 12.8005
R240 VTAIL.n392 VTAIL.n391 12.8005
R241 VTAIL.n38 VTAIL.n6 12.8005
R242 VTAIL.n42 VTAIL.n41 12.8005
R243 VTAIL.n88 VTAIL.n56 12.8005
R244 VTAIL.n92 VTAIL.n91 12.8005
R245 VTAIL.n138 VTAIL.n106 12.8005
R246 VTAIL.n142 VTAIL.n141 12.8005
R247 VTAIL.n342 VTAIL.n341 12.8005
R248 VTAIL.n338 VTAIL.n337 12.8005
R249 VTAIL.n292 VTAIL.n291 12.8005
R250 VTAIL.n288 VTAIL.n287 12.8005
R251 VTAIL.n242 VTAIL.n241 12.8005
R252 VTAIL.n238 VTAIL.n237 12.8005
R253 VTAIL.n192 VTAIL.n191 12.8005
R254 VTAIL.n188 VTAIL.n187 12.8005
R255 VTAIL.n383 VTAIL.n382 12.0247
R256 VTAIL.n395 VTAIL.n352 12.0247
R257 VTAIL.n33 VTAIL.n32 12.0247
R258 VTAIL.n45 VTAIL.n2 12.0247
R259 VTAIL.n83 VTAIL.n82 12.0247
R260 VTAIL.n95 VTAIL.n52 12.0247
R261 VTAIL.n133 VTAIL.n132 12.0247
R262 VTAIL.n145 VTAIL.n102 12.0247
R263 VTAIL.n345 VTAIL.n302 12.0247
R264 VTAIL.n334 VTAIL.n307 12.0247
R265 VTAIL.n295 VTAIL.n252 12.0247
R266 VTAIL.n284 VTAIL.n257 12.0247
R267 VTAIL.n245 VTAIL.n202 12.0247
R268 VTAIL.n234 VTAIL.n207 12.0247
R269 VTAIL.n195 VTAIL.n152 12.0247
R270 VTAIL.n184 VTAIL.n157 12.0247
R271 VTAIL.n381 VTAIL.n358 11.249
R272 VTAIL.n396 VTAIL.n350 11.249
R273 VTAIL.n31 VTAIL.n8 11.249
R274 VTAIL.n46 VTAIL.n0 11.249
R275 VTAIL.n81 VTAIL.n58 11.249
R276 VTAIL.n96 VTAIL.n50 11.249
R277 VTAIL.n131 VTAIL.n108 11.249
R278 VTAIL.n146 VTAIL.n100 11.249
R279 VTAIL.n346 VTAIL.n300 11.249
R280 VTAIL.n333 VTAIL.n310 11.249
R281 VTAIL.n296 VTAIL.n250 11.249
R282 VTAIL.n283 VTAIL.n260 11.249
R283 VTAIL.n246 VTAIL.n200 11.249
R284 VTAIL.n233 VTAIL.n210 11.249
R285 VTAIL.n196 VTAIL.n150 11.249
R286 VTAIL.n183 VTAIL.n160 11.249
R287 VTAIL.n378 VTAIL.n377 10.4732
R288 VTAIL.n28 VTAIL.n27 10.4732
R289 VTAIL.n78 VTAIL.n77 10.4732
R290 VTAIL.n128 VTAIL.n127 10.4732
R291 VTAIL.n330 VTAIL.n329 10.4732
R292 VTAIL.n280 VTAIL.n279 10.4732
R293 VTAIL.n230 VTAIL.n229 10.4732
R294 VTAIL.n180 VTAIL.n179 10.4732
R295 VTAIL.n366 VTAIL.n365 10.2747
R296 VTAIL.n16 VTAIL.n15 10.2747
R297 VTAIL.n66 VTAIL.n65 10.2747
R298 VTAIL.n116 VTAIL.n115 10.2747
R299 VTAIL.n318 VTAIL.n317 10.2747
R300 VTAIL.n268 VTAIL.n267 10.2747
R301 VTAIL.n218 VTAIL.n217 10.2747
R302 VTAIL.n168 VTAIL.n167 10.2747
R303 VTAIL.n374 VTAIL.n360 9.69747
R304 VTAIL.n24 VTAIL.n10 9.69747
R305 VTAIL.n74 VTAIL.n60 9.69747
R306 VTAIL.n124 VTAIL.n110 9.69747
R307 VTAIL.n326 VTAIL.n312 9.69747
R308 VTAIL.n276 VTAIL.n262 9.69747
R309 VTAIL.n226 VTAIL.n212 9.69747
R310 VTAIL.n176 VTAIL.n162 9.69747
R311 VTAIL.n398 VTAIL.n397 9.45567
R312 VTAIL.n48 VTAIL.n47 9.45567
R313 VTAIL.n98 VTAIL.n97 9.45567
R314 VTAIL.n148 VTAIL.n147 9.45567
R315 VTAIL.n348 VTAIL.n347 9.45567
R316 VTAIL.n298 VTAIL.n297 9.45567
R317 VTAIL.n248 VTAIL.n247 9.45567
R318 VTAIL.n198 VTAIL.n197 9.45567
R319 VTAIL.n397 VTAIL.n396 9.3005
R320 VTAIL.n352 VTAIL.n351 9.3005
R321 VTAIL.n391 VTAIL.n390 9.3005
R322 VTAIL.n364 VTAIL.n363 9.3005
R323 VTAIL.n371 VTAIL.n370 9.3005
R324 VTAIL.n373 VTAIL.n372 9.3005
R325 VTAIL.n360 VTAIL.n359 9.3005
R326 VTAIL.n379 VTAIL.n378 9.3005
R327 VTAIL.n381 VTAIL.n380 9.3005
R328 VTAIL.n382 VTAIL.n355 9.3005
R329 VTAIL.n389 VTAIL.n388 9.3005
R330 VTAIL.n47 VTAIL.n46 9.3005
R331 VTAIL.n2 VTAIL.n1 9.3005
R332 VTAIL.n41 VTAIL.n40 9.3005
R333 VTAIL.n14 VTAIL.n13 9.3005
R334 VTAIL.n21 VTAIL.n20 9.3005
R335 VTAIL.n23 VTAIL.n22 9.3005
R336 VTAIL.n10 VTAIL.n9 9.3005
R337 VTAIL.n29 VTAIL.n28 9.3005
R338 VTAIL.n31 VTAIL.n30 9.3005
R339 VTAIL.n32 VTAIL.n5 9.3005
R340 VTAIL.n39 VTAIL.n38 9.3005
R341 VTAIL.n97 VTAIL.n96 9.3005
R342 VTAIL.n52 VTAIL.n51 9.3005
R343 VTAIL.n91 VTAIL.n90 9.3005
R344 VTAIL.n64 VTAIL.n63 9.3005
R345 VTAIL.n71 VTAIL.n70 9.3005
R346 VTAIL.n73 VTAIL.n72 9.3005
R347 VTAIL.n60 VTAIL.n59 9.3005
R348 VTAIL.n79 VTAIL.n78 9.3005
R349 VTAIL.n81 VTAIL.n80 9.3005
R350 VTAIL.n82 VTAIL.n55 9.3005
R351 VTAIL.n89 VTAIL.n88 9.3005
R352 VTAIL.n147 VTAIL.n146 9.3005
R353 VTAIL.n102 VTAIL.n101 9.3005
R354 VTAIL.n141 VTAIL.n140 9.3005
R355 VTAIL.n114 VTAIL.n113 9.3005
R356 VTAIL.n121 VTAIL.n120 9.3005
R357 VTAIL.n123 VTAIL.n122 9.3005
R358 VTAIL.n110 VTAIL.n109 9.3005
R359 VTAIL.n129 VTAIL.n128 9.3005
R360 VTAIL.n131 VTAIL.n130 9.3005
R361 VTAIL.n132 VTAIL.n105 9.3005
R362 VTAIL.n139 VTAIL.n138 9.3005
R363 VTAIL.n316 VTAIL.n315 9.3005
R364 VTAIL.n323 VTAIL.n322 9.3005
R365 VTAIL.n325 VTAIL.n324 9.3005
R366 VTAIL.n312 VTAIL.n311 9.3005
R367 VTAIL.n331 VTAIL.n330 9.3005
R368 VTAIL.n333 VTAIL.n332 9.3005
R369 VTAIL.n307 VTAIL.n305 9.3005
R370 VTAIL.n339 VTAIL.n338 9.3005
R371 VTAIL.n347 VTAIL.n346 9.3005
R372 VTAIL.n302 VTAIL.n301 9.3005
R373 VTAIL.n341 VTAIL.n340 9.3005
R374 VTAIL.n266 VTAIL.n265 9.3005
R375 VTAIL.n273 VTAIL.n272 9.3005
R376 VTAIL.n275 VTAIL.n274 9.3005
R377 VTAIL.n262 VTAIL.n261 9.3005
R378 VTAIL.n281 VTAIL.n280 9.3005
R379 VTAIL.n283 VTAIL.n282 9.3005
R380 VTAIL.n257 VTAIL.n255 9.3005
R381 VTAIL.n289 VTAIL.n288 9.3005
R382 VTAIL.n297 VTAIL.n296 9.3005
R383 VTAIL.n252 VTAIL.n251 9.3005
R384 VTAIL.n291 VTAIL.n290 9.3005
R385 VTAIL.n216 VTAIL.n215 9.3005
R386 VTAIL.n223 VTAIL.n222 9.3005
R387 VTAIL.n225 VTAIL.n224 9.3005
R388 VTAIL.n212 VTAIL.n211 9.3005
R389 VTAIL.n231 VTAIL.n230 9.3005
R390 VTAIL.n233 VTAIL.n232 9.3005
R391 VTAIL.n207 VTAIL.n205 9.3005
R392 VTAIL.n239 VTAIL.n238 9.3005
R393 VTAIL.n247 VTAIL.n246 9.3005
R394 VTAIL.n202 VTAIL.n201 9.3005
R395 VTAIL.n241 VTAIL.n240 9.3005
R396 VTAIL.n166 VTAIL.n165 9.3005
R397 VTAIL.n173 VTAIL.n172 9.3005
R398 VTAIL.n175 VTAIL.n174 9.3005
R399 VTAIL.n162 VTAIL.n161 9.3005
R400 VTAIL.n181 VTAIL.n180 9.3005
R401 VTAIL.n183 VTAIL.n182 9.3005
R402 VTAIL.n157 VTAIL.n155 9.3005
R403 VTAIL.n189 VTAIL.n188 9.3005
R404 VTAIL.n197 VTAIL.n196 9.3005
R405 VTAIL.n152 VTAIL.n151 9.3005
R406 VTAIL.n191 VTAIL.n190 9.3005
R407 VTAIL.n373 VTAIL.n362 8.92171
R408 VTAIL.n23 VTAIL.n12 8.92171
R409 VTAIL.n73 VTAIL.n62 8.92171
R410 VTAIL.n123 VTAIL.n112 8.92171
R411 VTAIL.n325 VTAIL.n314 8.92171
R412 VTAIL.n275 VTAIL.n264 8.92171
R413 VTAIL.n225 VTAIL.n214 8.92171
R414 VTAIL.n175 VTAIL.n164 8.92171
R415 VTAIL.n370 VTAIL.n369 8.14595
R416 VTAIL.n20 VTAIL.n19 8.14595
R417 VTAIL.n70 VTAIL.n69 8.14595
R418 VTAIL.n120 VTAIL.n119 8.14595
R419 VTAIL.n322 VTAIL.n321 8.14595
R420 VTAIL.n272 VTAIL.n271 8.14595
R421 VTAIL.n222 VTAIL.n221 8.14595
R422 VTAIL.n172 VTAIL.n171 8.14595
R423 VTAIL.n366 VTAIL.n364 7.3702
R424 VTAIL.n16 VTAIL.n14 7.3702
R425 VTAIL.n66 VTAIL.n64 7.3702
R426 VTAIL.n116 VTAIL.n114 7.3702
R427 VTAIL.n318 VTAIL.n316 7.3702
R428 VTAIL.n268 VTAIL.n266 7.3702
R429 VTAIL.n218 VTAIL.n216 7.3702
R430 VTAIL.n168 VTAIL.n166 7.3702
R431 VTAIL.n369 VTAIL.n364 5.81868
R432 VTAIL.n19 VTAIL.n14 5.81868
R433 VTAIL.n69 VTAIL.n64 5.81868
R434 VTAIL.n119 VTAIL.n114 5.81868
R435 VTAIL.n321 VTAIL.n316 5.81868
R436 VTAIL.n271 VTAIL.n266 5.81868
R437 VTAIL.n221 VTAIL.n216 5.81868
R438 VTAIL.n171 VTAIL.n166 5.81868
R439 VTAIL.n370 VTAIL.n362 5.04292
R440 VTAIL.n20 VTAIL.n12 5.04292
R441 VTAIL.n70 VTAIL.n62 5.04292
R442 VTAIL.n120 VTAIL.n112 5.04292
R443 VTAIL.n322 VTAIL.n314 5.04292
R444 VTAIL.n272 VTAIL.n264 5.04292
R445 VTAIL.n222 VTAIL.n214 5.04292
R446 VTAIL.n172 VTAIL.n164 5.04292
R447 VTAIL.n374 VTAIL.n373 4.26717
R448 VTAIL.n24 VTAIL.n23 4.26717
R449 VTAIL.n74 VTAIL.n73 4.26717
R450 VTAIL.n124 VTAIL.n123 4.26717
R451 VTAIL.n326 VTAIL.n325 4.26717
R452 VTAIL.n276 VTAIL.n275 4.26717
R453 VTAIL.n226 VTAIL.n225 4.26717
R454 VTAIL.n176 VTAIL.n175 4.26717
R455 VTAIL.n249 VTAIL.n199 3.67291
R456 VTAIL.n349 VTAIL.n299 3.67291
R457 VTAIL.n149 VTAIL.n99 3.67291
R458 VTAIL.n377 VTAIL.n360 3.49141
R459 VTAIL.n27 VTAIL.n10 3.49141
R460 VTAIL.n77 VTAIL.n60 3.49141
R461 VTAIL.n127 VTAIL.n110 3.49141
R462 VTAIL.n329 VTAIL.n312 3.49141
R463 VTAIL.n279 VTAIL.n262 3.49141
R464 VTAIL.n229 VTAIL.n212 3.49141
R465 VTAIL.n179 VTAIL.n162 3.49141
R466 VTAIL.n365 VTAIL.n363 2.84303
R467 VTAIL.n15 VTAIL.n13 2.84303
R468 VTAIL.n65 VTAIL.n63 2.84303
R469 VTAIL.n115 VTAIL.n113 2.84303
R470 VTAIL.n317 VTAIL.n315 2.84303
R471 VTAIL.n267 VTAIL.n265 2.84303
R472 VTAIL.n217 VTAIL.n215 2.84303
R473 VTAIL.n167 VTAIL.n165 2.84303
R474 VTAIL.n378 VTAIL.n358 2.71565
R475 VTAIL.n398 VTAIL.n350 2.71565
R476 VTAIL.n28 VTAIL.n8 2.71565
R477 VTAIL.n48 VTAIL.n0 2.71565
R478 VTAIL.n78 VTAIL.n58 2.71565
R479 VTAIL.n98 VTAIL.n50 2.71565
R480 VTAIL.n128 VTAIL.n108 2.71565
R481 VTAIL.n148 VTAIL.n100 2.71565
R482 VTAIL.n348 VTAIL.n300 2.71565
R483 VTAIL.n330 VTAIL.n310 2.71565
R484 VTAIL.n298 VTAIL.n250 2.71565
R485 VTAIL.n280 VTAIL.n260 2.71565
R486 VTAIL.n248 VTAIL.n200 2.71565
R487 VTAIL.n230 VTAIL.n210 2.71565
R488 VTAIL.n198 VTAIL.n150 2.71565
R489 VTAIL.n180 VTAIL.n160 2.71565
R490 VTAIL.n383 VTAIL.n381 1.93989
R491 VTAIL.n396 VTAIL.n395 1.93989
R492 VTAIL.n33 VTAIL.n31 1.93989
R493 VTAIL.n46 VTAIL.n45 1.93989
R494 VTAIL.n83 VTAIL.n81 1.93989
R495 VTAIL.n96 VTAIL.n95 1.93989
R496 VTAIL.n133 VTAIL.n131 1.93989
R497 VTAIL.n146 VTAIL.n145 1.93989
R498 VTAIL.n346 VTAIL.n345 1.93989
R499 VTAIL.n334 VTAIL.n333 1.93989
R500 VTAIL.n296 VTAIL.n295 1.93989
R501 VTAIL.n284 VTAIL.n283 1.93989
R502 VTAIL.n246 VTAIL.n245 1.93989
R503 VTAIL.n234 VTAIL.n233 1.93989
R504 VTAIL.n196 VTAIL.n195 1.93989
R505 VTAIL.n184 VTAIL.n183 1.93989
R506 VTAIL VTAIL.n49 1.8949
R507 VTAIL VTAIL.n399 1.77852
R508 VTAIL.n382 VTAIL.n356 1.16414
R509 VTAIL.n392 VTAIL.n352 1.16414
R510 VTAIL.n32 VTAIL.n6 1.16414
R511 VTAIL.n42 VTAIL.n2 1.16414
R512 VTAIL.n82 VTAIL.n56 1.16414
R513 VTAIL.n92 VTAIL.n52 1.16414
R514 VTAIL.n132 VTAIL.n106 1.16414
R515 VTAIL.n142 VTAIL.n102 1.16414
R516 VTAIL.n342 VTAIL.n302 1.16414
R517 VTAIL.n337 VTAIL.n307 1.16414
R518 VTAIL.n292 VTAIL.n252 1.16414
R519 VTAIL.n287 VTAIL.n257 1.16414
R520 VTAIL.n242 VTAIL.n202 1.16414
R521 VTAIL.n237 VTAIL.n207 1.16414
R522 VTAIL.n192 VTAIL.n152 1.16414
R523 VTAIL.n187 VTAIL.n157 1.16414
R524 VTAIL.n299 VTAIL.n249 0.470328
R525 VTAIL.n99 VTAIL.n49 0.470328
R526 VTAIL.n388 VTAIL.n387 0.388379
R527 VTAIL.n391 VTAIL.n354 0.388379
R528 VTAIL.n38 VTAIL.n37 0.388379
R529 VTAIL.n41 VTAIL.n4 0.388379
R530 VTAIL.n88 VTAIL.n87 0.388379
R531 VTAIL.n91 VTAIL.n54 0.388379
R532 VTAIL.n138 VTAIL.n137 0.388379
R533 VTAIL.n141 VTAIL.n104 0.388379
R534 VTAIL.n341 VTAIL.n304 0.388379
R535 VTAIL.n338 VTAIL.n306 0.388379
R536 VTAIL.n291 VTAIL.n254 0.388379
R537 VTAIL.n288 VTAIL.n256 0.388379
R538 VTAIL.n241 VTAIL.n204 0.388379
R539 VTAIL.n238 VTAIL.n206 0.388379
R540 VTAIL.n191 VTAIL.n154 0.388379
R541 VTAIL.n188 VTAIL.n156 0.388379
R542 VTAIL.n371 VTAIL.n363 0.155672
R543 VTAIL.n372 VTAIL.n371 0.155672
R544 VTAIL.n372 VTAIL.n359 0.155672
R545 VTAIL.n379 VTAIL.n359 0.155672
R546 VTAIL.n380 VTAIL.n379 0.155672
R547 VTAIL.n380 VTAIL.n355 0.155672
R548 VTAIL.n389 VTAIL.n355 0.155672
R549 VTAIL.n390 VTAIL.n389 0.155672
R550 VTAIL.n390 VTAIL.n351 0.155672
R551 VTAIL.n397 VTAIL.n351 0.155672
R552 VTAIL.n21 VTAIL.n13 0.155672
R553 VTAIL.n22 VTAIL.n21 0.155672
R554 VTAIL.n22 VTAIL.n9 0.155672
R555 VTAIL.n29 VTAIL.n9 0.155672
R556 VTAIL.n30 VTAIL.n29 0.155672
R557 VTAIL.n30 VTAIL.n5 0.155672
R558 VTAIL.n39 VTAIL.n5 0.155672
R559 VTAIL.n40 VTAIL.n39 0.155672
R560 VTAIL.n40 VTAIL.n1 0.155672
R561 VTAIL.n47 VTAIL.n1 0.155672
R562 VTAIL.n71 VTAIL.n63 0.155672
R563 VTAIL.n72 VTAIL.n71 0.155672
R564 VTAIL.n72 VTAIL.n59 0.155672
R565 VTAIL.n79 VTAIL.n59 0.155672
R566 VTAIL.n80 VTAIL.n79 0.155672
R567 VTAIL.n80 VTAIL.n55 0.155672
R568 VTAIL.n89 VTAIL.n55 0.155672
R569 VTAIL.n90 VTAIL.n89 0.155672
R570 VTAIL.n90 VTAIL.n51 0.155672
R571 VTAIL.n97 VTAIL.n51 0.155672
R572 VTAIL.n121 VTAIL.n113 0.155672
R573 VTAIL.n122 VTAIL.n121 0.155672
R574 VTAIL.n122 VTAIL.n109 0.155672
R575 VTAIL.n129 VTAIL.n109 0.155672
R576 VTAIL.n130 VTAIL.n129 0.155672
R577 VTAIL.n130 VTAIL.n105 0.155672
R578 VTAIL.n139 VTAIL.n105 0.155672
R579 VTAIL.n140 VTAIL.n139 0.155672
R580 VTAIL.n140 VTAIL.n101 0.155672
R581 VTAIL.n147 VTAIL.n101 0.155672
R582 VTAIL.n347 VTAIL.n301 0.155672
R583 VTAIL.n340 VTAIL.n301 0.155672
R584 VTAIL.n340 VTAIL.n339 0.155672
R585 VTAIL.n339 VTAIL.n305 0.155672
R586 VTAIL.n332 VTAIL.n305 0.155672
R587 VTAIL.n332 VTAIL.n331 0.155672
R588 VTAIL.n331 VTAIL.n311 0.155672
R589 VTAIL.n324 VTAIL.n311 0.155672
R590 VTAIL.n324 VTAIL.n323 0.155672
R591 VTAIL.n323 VTAIL.n315 0.155672
R592 VTAIL.n297 VTAIL.n251 0.155672
R593 VTAIL.n290 VTAIL.n251 0.155672
R594 VTAIL.n290 VTAIL.n289 0.155672
R595 VTAIL.n289 VTAIL.n255 0.155672
R596 VTAIL.n282 VTAIL.n255 0.155672
R597 VTAIL.n282 VTAIL.n281 0.155672
R598 VTAIL.n281 VTAIL.n261 0.155672
R599 VTAIL.n274 VTAIL.n261 0.155672
R600 VTAIL.n274 VTAIL.n273 0.155672
R601 VTAIL.n273 VTAIL.n265 0.155672
R602 VTAIL.n247 VTAIL.n201 0.155672
R603 VTAIL.n240 VTAIL.n201 0.155672
R604 VTAIL.n240 VTAIL.n239 0.155672
R605 VTAIL.n239 VTAIL.n205 0.155672
R606 VTAIL.n232 VTAIL.n205 0.155672
R607 VTAIL.n232 VTAIL.n231 0.155672
R608 VTAIL.n231 VTAIL.n211 0.155672
R609 VTAIL.n224 VTAIL.n211 0.155672
R610 VTAIL.n224 VTAIL.n223 0.155672
R611 VTAIL.n223 VTAIL.n215 0.155672
R612 VTAIL.n197 VTAIL.n151 0.155672
R613 VTAIL.n190 VTAIL.n151 0.155672
R614 VTAIL.n190 VTAIL.n189 0.155672
R615 VTAIL.n189 VTAIL.n155 0.155672
R616 VTAIL.n182 VTAIL.n155 0.155672
R617 VTAIL.n182 VTAIL.n181 0.155672
R618 VTAIL.n181 VTAIL.n161 0.155672
R619 VTAIL.n174 VTAIL.n161 0.155672
R620 VTAIL.n174 VTAIL.n173 0.155672
R621 VTAIL.n173 VTAIL.n165 0.155672
R622 B.n762 B.n761 585
R623 B.n763 B.n762 585
R624 B.n280 B.n123 585
R625 B.n279 B.n278 585
R626 B.n277 B.n276 585
R627 B.n275 B.n274 585
R628 B.n273 B.n272 585
R629 B.n271 B.n270 585
R630 B.n269 B.n268 585
R631 B.n267 B.n266 585
R632 B.n265 B.n264 585
R633 B.n263 B.n262 585
R634 B.n261 B.n260 585
R635 B.n259 B.n258 585
R636 B.n257 B.n256 585
R637 B.n255 B.n254 585
R638 B.n253 B.n252 585
R639 B.n251 B.n250 585
R640 B.n249 B.n248 585
R641 B.n247 B.n246 585
R642 B.n245 B.n244 585
R643 B.n243 B.n242 585
R644 B.n241 B.n240 585
R645 B.n239 B.n238 585
R646 B.n237 B.n236 585
R647 B.n235 B.n234 585
R648 B.n233 B.n232 585
R649 B.n231 B.n230 585
R650 B.n229 B.n228 585
R651 B.n227 B.n226 585
R652 B.n225 B.n224 585
R653 B.n223 B.n222 585
R654 B.n221 B.n220 585
R655 B.n219 B.n218 585
R656 B.n217 B.n216 585
R657 B.n214 B.n213 585
R658 B.n212 B.n211 585
R659 B.n210 B.n209 585
R660 B.n208 B.n207 585
R661 B.n206 B.n205 585
R662 B.n204 B.n203 585
R663 B.n202 B.n201 585
R664 B.n200 B.n199 585
R665 B.n198 B.n197 585
R666 B.n196 B.n195 585
R667 B.n194 B.n193 585
R668 B.n192 B.n191 585
R669 B.n190 B.n189 585
R670 B.n188 B.n187 585
R671 B.n186 B.n185 585
R672 B.n184 B.n183 585
R673 B.n182 B.n181 585
R674 B.n180 B.n179 585
R675 B.n178 B.n177 585
R676 B.n176 B.n175 585
R677 B.n174 B.n173 585
R678 B.n172 B.n171 585
R679 B.n170 B.n169 585
R680 B.n168 B.n167 585
R681 B.n166 B.n165 585
R682 B.n164 B.n163 585
R683 B.n162 B.n161 585
R684 B.n160 B.n159 585
R685 B.n158 B.n157 585
R686 B.n156 B.n155 585
R687 B.n154 B.n153 585
R688 B.n152 B.n151 585
R689 B.n150 B.n149 585
R690 B.n148 B.n147 585
R691 B.n146 B.n145 585
R692 B.n144 B.n143 585
R693 B.n142 B.n141 585
R694 B.n140 B.n139 585
R695 B.n138 B.n137 585
R696 B.n136 B.n135 585
R697 B.n134 B.n133 585
R698 B.n132 B.n131 585
R699 B.n130 B.n129 585
R700 B.n760 B.n84 585
R701 B.n764 B.n84 585
R702 B.n759 B.n83 585
R703 B.n765 B.n83 585
R704 B.n758 B.n757 585
R705 B.n757 B.n79 585
R706 B.n756 B.n78 585
R707 B.n771 B.n78 585
R708 B.n755 B.n77 585
R709 B.n772 B.n77 585
R710 B.n754 B.n76 585
R711 B.n773 B.n76 585
R712 B.n753 B.n752 585
R713 B.n752 B.n72 585
R714 B.n751 B.n71 585
R715 B.n779 B.n71 585
R716 B.n750 B.n70 585
R717 B.n780 B.n70 585
R718 B.n749 B.n69 585
R719 B.n781 B.n69 585
R720 B.n748 B.n747 585
R721 B.n747 B.n65 585
R722 B.n746 B.n64 585
R723 B.n787 B.n64 585
R724 B.n745 B.n63 585
R725 B.n788 B.n63 585
R726 B.n744 B.n62 585
R727 B.n789 B.n62 585
R728 B.n743 B.n742 585
R729 B.n742 B.n58 585
R730 B.n741 B.n57 585
R731 B.n795 B.n57 585
R732 B.n740 B.n56 585
R733 B.n796 B.n56 585
R734 B.n739 B.n55 585
R735 B.n797 B.n55 585
R736 B.n738 B.n737 585
R737 B.n737 B.n51 585
R738 B.n736 B.n50 585
R739 B.n803 B.n50 585
R740 B.n735 B.n49 585
R741 B.n804 B.n49 585
R742 B.n734 B.n48 585
R743 B.n805 B.n48 585
R744 B.n733 B.n732 585
R745 B.n732 B.n44 585
R746 B.n731 B.n43 585
R747 B.n811 B.n43 585
R748 B.n730 B.n42 585
R749 B.n812 B.n42 585
R750 B.n729 B.n41 585
R751 B.n813 B.n41 585
R752 B.n728 B.n727 585
R753 B.n727 B.n37 585
R754 B.n726 B.n36 585
R755 B.n819 B.n36 585
R756 B.n725 B.n35 585
R757 B.n820 B.n35 585
R758 B.n724 B.n34 585
R759 B.n821 B.n34 585
R760 B.n723 B.n722 585
R761 B.n722 B.n30 585
R762 B.n721 B.n29 585
R763 B.n827 B.n29 585
R764 B.n720 B.n28 585
R765 B.n828 B.n28 585
R766 B.n719 B.n27 585
R767 B.n829 B.n27 585
R768 B.n718 B.n717 585
R769 B.n717 B.n23 585
R770 B.n716 B.n22 585
R771 B.n835 B.n22 585
R772 B.n715 B.n21 585
R773 B.n836 B.n21 585
R774 B.n714 B.n20 585
R775 B.n837 B.n20 585
R776 B.n713 B.n712 585
R777 B.n712 B.n16 585
R778 B.n711 B.n15 585
R779 B.n843 B.n15 585
R780 B.n710 B.n14 585
R781 B.n844 B.n14 585
R782 B.n709 B.n13 585
R783 B.n845 B.n13 585
R784 B.n708 B.n707 585
R785 B.n707 B.n12 585
R786 B.n706 B.n705 585
R787 B.n706 B.n8 585
R788 B.n704 B.n7 585
R789 B.n852 B.n7 585
R790 B.n703 B.n6 585
R791 B.n853 B.n6 585
R792 B.n702 B.n5 585
R793 B.n854 B.n5 585
R794 B.n701 B.n700 585
R795 B.n700 B.n4 585
R796 B.n699 B.n281 585
R797 B.n699 B.n698 585
R798 B.n689 B.n282 585
R799 B.n283 B.n282 585
R800 B.n691 B.n690 585
R801 B.n692 B.n691 585
R802 B.n688 B.n288 585
R803 B.n288 B.n287 585
R804 B.n687 B.n686 585
R805 B.n686 B.n685 585
R806 B.n290 B.n289 585
R807 B.n291 B.n290 585
R808 B.n678 B.n677 585
R809 B.n679 B.n678 585
R810 B.n676 B.n296 585
R811 B.n296 B.n295 585
R812 B.n675 B.n674 585
R813 B.n674 B.n673 585
R814 B.n298 B.n297 585
R815 B.n299 B.n298 585
R816 B.n666 B.n665 585
R817 B.n667 B.n666 585
R818 B.n664 B.n304 585
R819 B.n304 B.n303 585
R820 B.n663 B.n662 585
R821 B.n662 B.n661 585
R822 B.n306 B.n305 585
R823 B.n307 B.n306 585
R824 B.n654 B.n653 585
R825 B.n655 B.n654 585
R826 B.n652 B.n312 585
R827 B.n312 B.n311 585
R828 B.n651 B.n650 585
R829 B.n650 B.n649 585
R830 B.n314 B.n313 585
R831 B.n315 B.n314 585
R832 B.n642 B.n641 585
R833 B.n643 B.n642 585
R834 B.n640 B.n320 585
R835 B.n320 B.n319 585
R836 B.n639 B.n638 585
R837 B.n638 B.n637 585
R838 B.n322 B.n321 585
R839 B.n323 B.n322 585
R840 B.n630 B.n629 585
R841 B.n631 B.n630 585
R842 B.n628 B.n328 585
R843 B.n328 B.n327 585
R844 B.n627 B.n626 585
R845 B.n626 B.n625 585
R846 B.n330 B.n329 585
R847 B.n331 B.n330 585
R848 B.n618 B.n617 585
R849 B.n619 B.n618 585
R850 B.n616 B.n336 585
R851 B.n336 B.n335 585
R852 B.n615 B.n614 585
R853 B.n614 B.n613 585
R854 B.n338 B.n337 585
R855 B.n339 B.n338 585
R856 B.n606 B.n605 585
R857 B.n607 B.n606 585
R858 B.n604 B.n344 585
R859 B.n344 B.n343 585
R860 B.n603 B.n602 585
R861 B.n602 B.n601 585
R862 B.n346 B.n345 585
R863 B.n347 B.n346 585
R864 B.n594 B.n593 585
R865 B.n595 B.n594 585
R866 B.n592 B.n352 585
R867 B.n352 B.n351 585
R868 B.n591 B.n590 585
R869 B.n590 B.n589 585
R870 B.n354 B.n353 585
R871 B.n355 B.n354 585
R872 B.n582 B.n581 585
R873 B.n583 B.n582 585
R874 B.n580 B.n360 585
R875 B.n360 B.n359 585
R876 B.n579 B.n578 585
R877 B.n578 B.n577 585
R878 B.n362 B.n361 585
R879 B.n363 B.n362 585
R880 B.n570 B.n569 585
R881 B.n571 B.n570 585
R882 B.n568 B.n368 585
R883 B.n368 B.n367 585
R884 B.n562 B.n561 585
R885 B.n560 B.n408 585
R886 B.n559 B.n407 585
R887 B.n564 B.n407 585
R888 B.n558 B.n557 585
R889 B.n556 B.n555 585
R890 B.n554 B.n553 585
R891 B.n552 B.n551 585
R892 B.n550 B.n549 585
R893 B.n548 B.n547 585
R894 B.n546 B.n545 585
R895 B.n544 B.n543 585
R896 B.n542 B.n541 585
R897 B.n540 B.n539 585
R898 B.n538 B.n537 585
R899 B.n536 B.n535 585
R900 B.n534 B.n533 585
R901 B.n532 B.n531 585
R902 B.n530 B.n529 585
R903 B.n528 B.n527 585
R904 B.n526 B.n525 585
R905 B.n524 B.n523 585
R906 B.n522 B.n521 585
R907 B.n520 B.n519 585
R908 B.n518 B.n517 585
R909 B.n516 B.n515 585
R910 B.n514 B.n513 585
R911 B.n512 B.n511 585
R912 B.n510 B.n509 585
R913 B.n508 B.n507 585
R914 B.n506 B.n505 585
R915 B.n504 B.n503 585
R916 B.n502 B.n501 585
R917 B.n500 B.n499 585
R918 B.n498 B.n497 585
R919 B.n495 B.n494 585
R920 B.n493 B.n492 585
R921 B.n491 B.n490 585
R922 B.n489 B.n488 585
R923 B.n487 B.n486 585
R924 B.n485 B.n484 585
R925 B.n483 B.n482 585
R926 B.n481 B.n480 585
R927 B.n479 B.n478 585
R928 B.n477 B.n476 585
R929 B.n475 B.n474 585
R930 B.n473 B.n472 585
R931 B.n471 B.n470 585
R932 B.n469 B.n468 585
R933 B.n467 B.n466 585
R934 B.n465 B.n464 585
R935 B.n463 B.n462 585
R936 B.n461 B.n460 585
R937 B.n459 B.n458 585
R938 B.n457 B.n456 585
R939 B.n455 B.n454 585
R940 B.n453 B.n452 585
R941 B.n451 B.n450 585
R942 B.n449 B.n448 585
R943 B.n447 B.n446 585
R944 B.n445 B.n444 585
R945 B.n443 B.n442 585
R946 B.n441 B.n440 585
R947 B.n439 B.n438 585
R948 B.n437 B.n436 585
R949 B.n435 B.n434 585
R950 B.n433 B.n432 585
R951 B.n431 B.n430 585
R952 B.n429 B.n428 585
R953 B.n427 B.n426 585
R954 B.n425 B.n424 585
R955 B.n423 B.n422 585
R956 B.n421 B.n420 585
R957 B.n419 B.n418 585
R958 B.n417 B.n416 585
R959 B.n415 B.n414 585
R960 B.n370 B.n369 585
R961 B.n567 B.n566 585
R962 B.n366 B.n365 585
R963 B.n367 B.n366 585
R964 B.n573 B.n572 585
R965 B.n572 B.n571 585
R966 B.n574 B.n364 585
R967 B.n364 B.n363 585
R968 B.n576 B.n575 585
R969 B.n577 B.n576 585
R970 B.n358 B.n357 585
R971 B.n359 B.n358 585
R972 B.n585 B.n584 585
R973 B.n584 B.n583 585
R974 B.n586 B.n356 585
R975 B.n356 B.n355 585
R976 B.n588 B.n587 585
R977 B.n589 B.n588 585
R978 B.n350 B.n349 585
R979 B.n351 B.n350 585
R980 B.n597 B.n596 585
R981 B.n596 B.n595 585
R982 B.n598 B.n348 585
R983 B.n348 B.n347 585
R984 B.n600 B.n599 585
R985 B.n601 B.n600 585
R986 B.n342 B.n341 585
R987 B.n343 B.n342 585
R988 B.n609 B.n608 585
R989 B.n608 B.n607 585
R990 B.n610 B.n340 585
R991 B.n340 B.n339 585
R992 B.n612 B.n611 585
R993 B.n613 B.n612 585
R994 B.n334 B.n333 585
R995 B.n335 B.n334 585
R996 B.n621 B.n620 585
R997 B.n620 B.n619 585
R998 B.n622 B.n332 585
R999 B.n332 B.n331 585
R1000 B.n624 B.n623 585
R1001 B.n625 B.n624 585
R1002 B.n326 B.n325 585
R1003 B.n327 B.n326 585
R1004 B.n633 B.n632 585
R1005 B.n632 B.n631 585
R1006 B.n634 B.n324 585
R1007 B.n324 B.n323 585
R1008 B.n636 B.n635 585
R1009 B.n637 B.n636 585
R1010 B.n318 B.n317 585
R1011 B.n319 B.n318 585
R1012 B.n645 B.n644 585
R1013 B.n644 B.n643 585
R1014 B.n646 B.n316 585
R1015 B.n316 B.n315 585
R1016 B.n648 B.n647 585
R1017 B.n649 B.n648 585
R1018 B.n310 B.n309 585
R1019 B.n311 B.n310 585
R1020 B.n657 B.n656 585
R1021 B.n656 B.n655 585
R1022 B.n658 B.n308 585
R1023 B.n308 B.n307 585
R1024 B.n660 B.n659 585
R1025 B.n661 B.n660 585
R1026 B.n302 B.n301 585
R1027 B.n303 B.n302 585
R1028 B.n669 B.n668 585
R1029 B.n668 B.n667 585
R1030 B.n670 B.n300 585
R1031 B.n300 B.n299 585
R1032 B.n672 B.n671 585
R1033 B.n673 B.n672 585
R1034 B.n294 B.n293 585
R1035 B.n295 B.n294 585
R1036 B.n681 B.n680 585
R1037 B.n680 B.n679 585
R1038 B.n682 B.n292 585
R1039 B.n292 B.n291 585
R1040 B.n684 B.n683 585
R1041 B.n685 B.n684 585
R1042 B.n286 B.n285 585
R1043 B.n287 B.n286 585
R1044 B.n694 B.n693 585
R1045 B.n693 B.n692 585
R1046 B.n695 B.n284 585
R1047 B.n284 B.n283 585
R1048 B.n697 B.n696 585
R1049 B.n698 B.n697 585
R1050 B.n3 B.n0 585
R1051 B.n4 B.n3 585
R1052 B.n851 B.n1 585
R1053 B.n852 B.n851 585
R1054 B.n850 B.n849 585
R1055 B.n850 B.n8 585
R1056 B.n848 B.n9 585
R1057 B.n12 B.n9 585
R1058 B.n847 B.n846 585
R1059 B.n846 B.n845 585
R1060 B.n11 B.n10 585
R1061 B.n844 B.n11 585
R1062 B.n842 B.n841 585
R1063 B.n843 B.n842 585
R1064 B.n840 B.n17 585
R1065 B.n17 B.n16 585
R1066 B.n839 B.n838 585
R1067 B.n838 B.n837 585
R1068 B.n19 B.n18 585
R1069 B.n836 B.n19 585
R1070 B.n834 B.n833 585
R1071 B.n835 B.n834 585
R1072 B.n832 B.n24 585
R1073 B.n24 B.n23 585
R1074 B.n831 B.n830 585
R1075 B.n830 B.n829 585
R1076 B.n26 B.n25 585
R1077 B.n828 B.n26 585
R1078 B.n826 B.n825 585
R1079 B.n827 B.n826 585
R1080 B.n824 B.n31 585
R1081 B.n31 B.n30 585
R1082 B.n823 B.n822 585
R1083 B.n822 B.n821 585
R1084 B.n33 B.n32 585
R1085 B.n820 B.n33 585
R1086 B.n818 B.n817 585
R1087 B.n819 B.n818 585
R1088 B.n816 B.n38 585
R1089 B.n38 B.n37 585
R1090 B.n815 B.n814 585
R1091 B.n814 B.n813 585
R1092 B.n40 B.n39 585
R1093 B.n812 B.n40 585
R1094 B.n810 B.n809 585
R1095 B.n811 B.n810 585
R1096 B.n808 B.n45 585
R1097 B.n45 B.n44 585
R1098 B.n807 B.n806 585
R1099 B.n806 B.n805 585
R1100 B.n47 B.n46 585
R1101 B.n804 B.n47 585
R1102 B.n802 B.n801 585
R1103 B.n803 B.n802 585
R1104 B.n800 B.n52 585
R1105 B.n52 B.n51 585
R1106 B.n799 B.n798 585
R1107 B.n798 B.n797 585
R1108 B.n54 B.n53 585
R1109 B.n796 B.n54 585
R1110 B.n794 B.n793 585
R1111 B.n795 B.n794 585
R1112 B.n792 B.n59 585
R1113 B.n59 B.n58 585
R1114 B.n791 B.n790 585
R1115 B.n790 B.n789 585
R1116 B.n61 B.n60 585
R1117 B.n788 B.n61 585
R1118 B.n786 B.n785 585
R1119 B.n787 B.n786 585
R1120 B.n784 B.n66 585
R1121 B.n66 B.n65 585
R1122 B.n783 B.n782 585
R1123 B.n782 B.n781 585
R1124 B.n68 B.n67 585
R1125 B.n780 B.n68 585
R1126 B.n778 B.n777 585
R1127 B.n779 B.n778 585
R1128 B.n776 B.n73 585
R1129 B.n73 B.n72 585
R1130 B.n775 B.n774 585
R1131 B.n774 B.n773 585
R1132 B.n75 B.n74 585
R1133 B.n772 B.n75 585
R1134 B.n770 B.n769 585
R1135 B.n771 B.n770 585
R1136 B.n768 B.n80 585
R1137 B.n80 B.n79 585
R1138 B.n767 B.n766 585
R1139 B.n766 B.n765 585
R1140 B.n82 B.n81 585
R1141 B.n764 B.n82 585
R1142 B.n855 B.n854 585
R1143 B.n853 B.n2 585
R1144 B.n129 B.n82 521.33
R1145 B.n762 B.n84 521.33
R1146 B.n566 B.n368 521.33
R1147 B.n562 B.n366 521.33
R1148 B.n124 B.t16 317.971
R1149 B.n411 B.t7 317.971
R1150 B.n126 B.t13 317.971
R1151 B.n409 B.t10 317.971
R1152 B.n126 B.t11 266.411
R1153 B.n124 B.t15 266.411
R1154 B.n411 B.t4 266.411
R1155 B.n409 B.t8 266.411
R1156 B.n763 B.n122 256.663
R1157 B.n763 B.n121 256.663
R1158 B.n763 B.n120 256.663
R1159 B.n763 B.n119 256.663
R1160 B.n763 B.n118 256.663
R1161 B.n763 B.n117 256.663
R1162 B.n763 B.n116 256.663
R1163 B.n763 B.n115 256.663
R1164 B.n763 B.n114 256.663
R1165 B.n763 B.n113 256.663
R1166 B.n763 B.n112 256.663
R1167 B.n763 B.n111 256.663
R1168 B.n763 B.n110 256.663
R1169 B.n763 B.n109 256.663
R1170 B.n763 B.n108 256.663
R1171 B.n763 B.n107 256.663
R1172 B.n763 B.n106 256.663
R1173 B.n763 B.n105 256.663
R1174 B.n763 B.n104 256.663
R1175 B.n763 B.n103 256.663
R1176 B.n763 B.n102 256.663
R1177 B.n763 B.n101 256.663
R1178 B.n763 B.n100 256.663
R1179 B.n763 B.n99 256.663
R1180 B.n763 B.n98 256.663
R1181 B.n763 B.n97 256.663
R1182 B.n763 B.n96 256.663
R1183 B.n763 B.n95 256.663
R1184 B.n763 B.n94 256.663
R1185 B.n763 B.n93 256.663
R1186 B.n763 B.n92 256.663
R1187 B.n763 B.n91 256.663
R1188 B.n763 B.n90 256.663
R1189 B.n763 B.n89 256.663
R1190 B.n763 B.n88 256.663
R1191 B.n763 B.n87 256.663
R1192 B.n763 B.n86 256.663
R1193 B.n763 B.n85 256.663
R1194 B.n564 B.n563 256.663
R1195 B.n564 B.n371 256.663
R1196 B.n564 B.n372 256.663
R1197 B.n564 B.n373 256.663
R1198 B.n564 B.n374 256.663
R1199 B.n564 B.n375 256.663
R1200 B.n564 B.n376 256.663
R1201 B.n564 B.n377 256.663
R1202 B.n564 B.n378 256.663
R1203 B.n564 B.n379 256.663
R1204 B.n564 B.n380 256.663
R1205 B.n564 B.n381 256.663
R1206 B.n564 B.n382 256.663
R1207 B.n564 B.n383 256.663
R1208 B.n564 B.n384 256.663
R1209 B.n564 B.n385 256.663
R1210 B.n564 B.n386 256.663
R1211 B.n564 B.n387 256.663
R1212 B.n564 B.n388 256.663
R1213 B.n564 B.n389 256.663
R1214 B.n564 B.n390 256.663
R1215 B.n564 B.n391 256.663
R1216 B.n564 B.n392 256.663
R1217 B.n564 B.n393 256.663
R1218 B.n564 B.n394 256.663
R1219 B.n564 B.n395 256.663
R1220 B.n564 B.n396 256.663
R1221 B.n564 B.n397 256.663
R1222 B.n564 B.n398 256.663
R1223 B.n564 B.n399 256.663
R1224 B.n564 B.n400 256.663
R1225 B.n564 B.n401 256.663
R1226 B.n564 B.n402 256.663
R1227 B.n564 B.n403 256.663
R1228 B.n564 B.n404 256.663
R1229 B.n564 B.n405 256.663
R1230 B.n564 B.n406 256.663
R1231 B.n565 B.n564 256.663
R1232 B.n857 B.n856 256.663
R1233 B.n125 B.t17 235.353
R1234 B.n412 B.t6 235.353
R1235 B.n127 B.t14 235.353
R1236 B.n410 B.t9 235.353
R1237 B.n133 B.n132 163.367
R1238 B.n137 B.n136 163.367
R1239 B.n141 B.n140 163.367
R1240 B.n145 B.n144 163.367
R1241 B.n149 B.n148 163.367
R1242 B.n153 B.n152 163.367
R1243 B.n157 B.n156 163.367
R1244 B.n161 B.n160 163.367
R1245 B.n165 B.n164 163.367
R1246 B.n169 B.n168 163.367
R1247 B.n173 B.n172 163.367
R1248 B.n177 B.n176 163.367
R1249 B.n181 B.n180 163.367
R1250 B.n185 B.n184 163.367
R1251 B.n189 B.n188 163.367
R1252 B.n193 B.n192 163.367
R1253 B.n197 B.n196 163.367
R1254 B.n201 B.n200 163.367
R1255 B.n205 B.n204 163.367
R1256 B.n209 B.n208 163.367
R1257 B.n213 B.n212 163.367
R1258 B.n218 B.n217 163.367
R1259 B.n222 B.n221 163.367
R1260 B.n226 B.n225 163.367
R1261 B.n230 B.n229 163.367
R1262 B.n234 B.n233 163.367
R1263 B.n238 B.n237 163.367
R1264 B.n242 B.n241 163.367
R1265 B.n246 B.n245 163.367
R1266 B.n250 B.n249 163.367
R1267 B.n254 B.n253 163.367
R1268 B.n258 B.n257 163.367
R1269 B.n262 B.n261 163.367
R1270 B.n266 B.n265 163.367
R1271 B.n270 B.n269 163.367
R1272 B.n274 B.n273 163.367
R1273 B.n278 B.n277 163.367
R1274 B.n762 B.n123 163.367
R1275 B.n570 B.n368 163.367
R1276 B.n570 B.n362 163.367
R1277 B.n578 B.n362 163.367
R1278 B.n578 B.n360 163.367
R1279 B.n582 B.n360 163.367
R1280 B.n582 B.n354 163.367
R1281 B.n590 B.n354 163.367
R1282 B.n590 B.n352 163.367
R1283 B.n594 B.n352 163.367
R1284 B.n594 B.n346 163.367
R1285 B.n602 B.n346 163.367
R1286 B.n602 B.n344 163.367
R1287 B.n606 B.n344 163.367
R1288 B.n606 B.n338 163.367
R1289 B.n614 B.n338 163.367
R1290 B.n614 B.n336 163.367
R1291 B.n618 B.n336 163.367
R1292 B.n618 B.n330 163.367
R1293 B.n626 B.n330 163.367
R1294 B.n626 B.n328 163.367
R1295 B.n630 B.n328 163.367
R1296 B.n630 B.n322 163.367
R1297 B.n638 B.n322 163.367
R1298 B.n638 B.n320 163.367
R1299 B.n642 B.n320 163.367
R1300 B.n642 B.n314 163.367
R1301 B.n650 B.n314 163.367
R1302 B.n650 B.n312 163.367
R1303 B.n654 B.n312 163.367
R1304 B.n654 B.n306 163.367
R1305 B.n662 B.n306 163.367
R1306 B.n662 B.n304 163.367
R1307 B.n666 B.n304 163.367
R1308 B.n666 B.n298 163.367
R1309 B.n674 B.n298 163.367
R1310 B.n674 B.n296 163.367
R1311 B.n678 B.n296 163.367
R1312 B.n678 B.n290 163.367
R1313 B.n686 B.n290 163.367
R1314 B.n686 B.n288 163.367
R1315 B.n691 B.n288 163.367
R1316 B.n691 B.n282 163.367
R1317 B.n699 B.n282 163.367
R1318 B.n700 B.n699 163.367
R1319 B.n700 B.n5 163.367
R1320 B.n6 B.n5 163.367
R1321 B.n7 B.n6 163.367
R1322 B.n706 B.n7 163.367
R1323 B.n707 B.n706 163.367
R1324 B.n707 B.n13 163.367
R1325 B.n14 B.n13 163.367
R1326 B.n15 B.n14 163.367
R1327 B.n712 B.n15 163.367
R1328 B.n712 B.n20 163.367
R1329 B.n21 B.n20 163.367
R1330 B.n22 B.n21 163.367
R1331 B.n717 B.n22 163.367
R1332 B.n717 B.n27 163.367
R1333 B.n28 B.n27 163.367
R1334 B.n29 B.n28 163.367
R1335 B.n722 B.n29 163.367
R1336 B.n722 B.n34 163.367
R1337 B.n35 B.n34 163.367
R1338 B.n36 B.n35 163.367
R1339 B.n727 B.n36 163.367
R1340 B.n727 B.n41 163.367
R1341 B.n42 B.n41 163.367
R1342 B.n43 B.n42 163.367
R1343 B.n732 B.n43 163.367
R1344 B.n732 B.n48 163.367
R1345 B.n49 B.n48 163.367
R1346 B.n50 B.n49 163.367
R1347 B.n737 B.n50 163.367
R1348 B.n737 B.n55 163.367
R1349 B.n56 B.n55 163.367
R1350 B.n57 B.n56 163.367
R1351 B.n742 B.n57 163.367
R1352 B.n742 B.n62 163.367
R1353 B.n63 B.n62 163.367
R1354 B.n64 B.n63 163.367
R1355 B.n747 B.n64 163.367
R1356 B.n747 B.n69 163.367
R1357 B.n70 B.n69 163.367
R1358 B.n71 B.n70 163.367
R1359 B.n752 B.n71 163.367
R1360 B.n752 B.n76 163.367
R1361 B.n77 B.n76 163.367
R1362 B.n78 B.n77 163.367
R1363 B.n757 B.n78 163.367
R1364 B.n757 B.n83 163.367
R1365 B.n84 B.n83 163.367
R1366 B.n408 B.n407 163.367
R1367 B.n557 B.n407 163.367
R1368 B.n555 B.n554 163.367
R1369 B.n551 B.n550 163.367
R1370 B.n547 B.n546 163.367
R1371 B.n543 B.n542 163.367
R1372 B.n539 B.n538 163.367
R1373 B.n535 B.n534 163.367
R1374 B.n531 B.n530 163.367
R1375 B.n527 B.n526 163.367
R1376 B.n523 B.n522 163.367
R1377 B.n519 B.n518 163.367
R1378 B.n515 B.n514 163.367
R1379 B.n511 B.n510 163.367
R1380 B.n507 B.n506 163.367
R1381 B.n503 B.n502 163.367
R1382 B.n499 B.n498 163.367
R1383 B.n494 B.n493 163.367
R1384 B.n490 B.n489 163.367
R1385 B.n486 B.n485 163.367
R1386 B.n482 B.n481 163.367
R1387 B.n478 B.n477 163.367
R1388 B.n474 B.n473 163.367
R1389 B.n470 B.n469 163.367
R1390 B.n466 B.n465 163.367
R1391 B.n462 B.n461 163.367
R1392 B.n458 B.n457 163.367
R1393 B.n454 B.n453 163.367
R1394 B.n450 B.n449 163.367
R1395 B.n446 B.n445 163.367
R1396 B.n442 B.n441 163.367
R1397 B.n438 B.n437 163.367
R1398 B.n434 B.n433 163.367
R1399 B.n430 B.n429 163.367
R1400 B.n426 B.n425 163.367
R1401 B.n422 B.n421 163.367
R1402 B.n418 B.n417 163.367
R1403 B.n414 B.n370 163.367
R1404 B.n572 B.n366 163.367
R1405 B.n572 B.n364 163.367
R1406 B.n576 B.n364 163.367
R1407 B.n576 B.n358 163.367
R1408 B.n584 B.n358 163.367
R1409 B.n584 B.n356 163.367
R1410 B.n588 B.n356 163.367
R1411 B.n588 B.n350 163.367
R1412 B.n596 B.n350 163.367
R1413 B.n596 B.n348 163.367
R1414 B.n600 B.n348 163.367
R1415 B.n600 B.n342 163.367
R1416 B.n608 B.n342 163.367
R1417 B.n608 B.n340 163.367
R1418 B.n612 B.n340 163.367
R1419 B.n612 B.n334 163.367
R1420 B.n620 B.n334 163.367
R1421 B.n620 B.n332 163.367
R1422 B.n624 B.n332 163.367
R1423 B.n624 B.n326 163.367
R1424 B.n632 B.n326 163.367
R1425 B.n632 B.n324 163.367
R1426 B.n636 B.n324 163.367
R1427 B.n636 B.n318 163.367
R1428 B.n644 B.n318 163.367
R1429 B.n644 B.n316 163.367
R1430 B.n648 B.n316 163.367
R1431 B.n648 B.n310 163.367
R1432 B.n656 B.n310 163.367
R1433 B.n656 B.n308 163.367
R1434 B.n660 B.n308 163.367
R1435 B.n660 B.n302 163.367
R1436 B.n668 B.n302 163.367
R1437 B.n668 B.n300 163.367
R1438 B.n672 B.n300 163.367
R1439 B.n672 B.n294 163.367
R1440 B.n680 B.n294 163.367
R1441 B.n680 B.n292 163.367
R1442 B.n684 B.n292 163.367
R1443 B.n684 B.n286 163.367
R1444 B.n693 B.n286 163.367
R1445 B.n693 B.n284 163.367
R1446 B.n697 B.n284 163.367
R1447 B.n697 B.n3 163.367
R1448 B.n855 B.n3 163.367
R1449 B.n851 B.n2 163.367
R1450 B.n851 B.n850 163.367
R1451 B.n850 B.n9 163.367
R1452 B.n846 B.n9 163.367
R1453 B.n846 B.n11 163.367
R1454 B.n842 B.n11 163.367
R1455 B.n842 B.n17 163.367
R1456 B.n838 B.n17 163.367
R1457 B.n838 B.n19 163.367
R1458 B.n834 B.n19 163.367
R1459 B.n834 B.n24 163.367
R1460 B.n830 B.n24 163.367
R1461 B.n830 B.n26 163.367
R1462 B.n826 B.n26 163.367
R1463 B.n826 B.n31 163.367
R1464 B.n822 B.n31 163.367
R1465 B.n822 B.n33 163.367
R1466 B.n818 B.n33 163.367
R1467 B.n818 B.n38 163.367
R1468 B.n814 B.n38 163.367
R1469 B.n814 B.n40 163.367
R1470 B.n810 B.n40 163.367
R1471 B.n810 B.n45 163.367
R1472 B.n806 B.n45 163.367
R1473 B.n806 B.n47 163.367
R1474 B.n802 B.n47 163.367
R1475 B.n802 B.n52 163.367
R1476 B.n798 B.n52 163.367
R1477 B.n798 B.n54 163.367
R1478 B.n794 B.n54 163.367
R1479 B.n794 B.n59 163.367
R1480 B.n790 B.n59 163.367
R1481 B.n790 B.n61 163.367
R1482 B.n786 B.n61 163.367
R1483 B.n786 B.n66 163.367
R1484 B.n782 B.n66 163.367
R1485 B.n782 B.n68 163.367
R1486 B.n778 B.n68 163.367
R1487 B.n778 B.n73 163.367
R1488 B.n774 B.n73 163.367
R1489 B.n774 B.n75 163.367
R1490 B.n770 B.n75 163.367
R1491 B.n770 B.n80 163.367
R1492 B.n766 B.n80 163.367
R1493 B.n766 B.n82 163.367
R1494 B.n564 B.n367 103.468
R1495 B.n764 B.n763 103.468
R1496 B.n127 B.n126 82.6187
R1497 B.n125 B.n124 82.6187
R1498 B.n412 B.n411 82.6187
R1499 B.n410 B.n409 82.6187
R1500 B.n129 B.n85 71.676
R1501 B.n133 B.n86 71.676
R1502 B.n137 B.n87 71.676
R1503 B.n141 B.n88 71.676
R1504 B.n145 B.n89 71.676
R1505 B.n149 B.n90 71.676
R1506 B.n153 B.n91 71.676
R1507 B.n157 B.n92 71.676
R1508 B.n161 B.n93 71.676
R1509 B.n165 B.n94 71.676
R1510 B.n169 B.n95 71.676
R1511 B.n173 B.n96 71.676
R1512 B.n177 B.n97 71.676
R1513 B.n181 B.n98 71.676
R1514 B.n185 B.n99 71.676
R1515 B.n189 B.n100 71.676
R1516 B.n193 B.n101 71.676
R1517 B.n197 B.n102 71.676
R1518 B.n201 B.n103 71.676
R1519 B.n205 B.n104 71.676
R1520 B.n209 B.n105 71.676
R1521 B.n213 B.n106 71.676
R1522 B.n218 B.n107 71.676
R1523 B.n222 B.n108 71.676
R1524 B.n226 B.n109 71.676
R1525 B.n230 B.n110 71.676
R1526 B.n234 B.n111 71.676
R1527 B.n238 B.n112 71.676
R1528 B.n242 B.n113 71.676
R1529 B.n246 B.n114 71.676
R1530 B.n250 B.n115 71.676
R1531 B.n254 B.n116 71.676
R1532 B.n258 B.n117 71.676
R1533 B.n262 B.n118 71.676
R1534 B.n266 B.n119 71.676
R1535 B.n270 B.n120 71.676
R1536 B.n274 B.n121 71.676
R1537 B.n278 B.n122 71.676
R1538 B.n123 B.n122 71.676
R1539 B.n277 B.n121 71.676
R1540 B.n273 B.n120 71.676
R1541 B.n269 B.n119 71.676
R1542 B.n265 B.n118 71.676
R1543 B.n261 B.n117 71.676
R1544 B.n257 B.n116 71.676
R1545 B.n253 B.n115 71.676
R1546 B.n249 B.n114 71.676
R1547 B.n245 B.n113 71.676
R1548 B.n241 B.n112 71.676
R1549 B.n237 B.n111 71.676
R1550 B.n233 B.n110 71.676
R1551 B.n229 B.n109 71.676
R1552 B.n225 B.n108 71.676
R1553 B.n221 B.n107 71.676
R1554 B.n217 B.n106 71.676
R1555 B.n212 B.n105 71.676
R1556 B.n208 B.n104 71.676
R1557 B.n204 B.n103 71.676
R1558 B.n200 B.n102 71.676
R1559 B.n196 B.n101 71.676
R1560 B.n192 B.n100 71.676
R1561 B.n188 B.n99 71.676
R1562 B.n184 B.n98 71.676
R1563 B.n180 B.n97 71.676
R1564 B.n176 B.n96 71.676
R1565 B.n172 B.n95 71.676
R1566 B.n168 B.n94 71.676
R1567 B.n164 B.n93 71.676
R1568 B.n160 B.n92 71.676
R1569 B.n156 B.n91 71.676
R1570 B.n152 B.n90 71.676
R1571 B.n148 B.n89 71.676
R1572 B.n144 B.n88 71.676
R1573 B.n140 B.n87 71.676
R1574 B.n136 B.n86 71.676
R1575 B.n132 B.n85 71.676
R1576 B.n563 B.n562 71.676
R1577 B.n557 B.n371 71.676
R1578 B.n554 B.n372 71.676
R1579 B.n550 B.n373 71.676
R1580 B.n546 B.n374 71.676
R1581 B.n542 B.n375 71.676
R1582 B.n538 B.n376 71.676
R1583 B.n534 B.n377 71.676
R1584 B.n530 B.n378 71.676
R1585 B.n526 B.n379 71.676
R1586 B.n522 B.n380 71.676
R1587 B.n518 B.n381 71.676
R1588 B.n514 B.n382 71.676
R1589 B.n510 B.n383 71.676
R1590 B.n506 B.n384 71.676
R1591 B.n502 B.n385 71.676
R1592 B.n498 B.n386 71.676
R1593 B.n493 B.n387 71.676
R1594 B.n489 B.n388 71.676
R1595 B.n485 B.n389 71.676
R1596 B.n481 B.n390 71.676
R1597 B.n477 B.n391 71.676
R1598 B.n473 B.n392 71.676
R1599 B.n469 B.n393 71.676
R1600 B.n465 B.n394 71.676
R1601 B.n461 B.n395 71.676
R1602 B.n457 B.n396 71.676
R1603 B.n453 B.n397 71.676
R1604 B.n449 B.n398 71.676
R1605 B.n445 B.n399 71.676
R1606 B.n441 B.n400 71.676
R1607 B.n437 B.n401 71.676
R1608 B.n433 B.n402 71.676
R1609 B.n429 B.n403 71.676
R1610 B.n425 B.n404 71.676
R1611 B.n421 B.n405 71.676
R1612 B.n417 B.n406 71.676
R1613 B.n565 B.n370 71.676
R1614 B.n563 B.n408 71.676
R1615 B.n555 B.n371 71.676
R1616 B.n551 B.n372 71.676
R1617 B.n547 B.n373 71.676
R1618 B.n543 B.n374 71.676
R1619 B.n539 B.n375 71.676
R1620 B.n535 B.n376 71.676
R1621 B.n531 B.n377 71.676
R1622 B.n527 B.n378 71.676
R1623 B.n523 B.n379 71.676
R1624 B.n519 B.n380 71.676
R1625 B.n515 B.n381 71.676
R1626 B.n511 B.n382 71.676
R1627 B.n507 B.n383 71.676
R1628 B.n503 B.n384 71.676
R1629 B.n499 B.n385 71.676
R1630 B.n494 B.n386 71.676
R1631 B.n490 B.n387 71.676
R1632 B.n486 B.n388 71.676
R1633 B.n482 B.n389 71.676
R1634 B.n478 B.n390 71.676
R1635 B.n474 B.n391 71.676
R1636 B.n470 B.n392 71.676
R1637 B.n466 B.n393 71.676
R1638 B.n462 B.n394 71.676
R1639 B.n458 B.n395 71.676
R1640 B.n454 B.n396 71.676
R1641 B.n450 B.n397 71.676
R1642 B.n446 B.n398 71.676
R1643 B.n442 B.n399 71.676
R1644 B.n438 B.n400 71.676
R1645 B.n434 B.n401 71.676
R1646 B.n430 B.n402 71.676
R1647 B.n426 B.n403 71.676
R1648 B.n422 B.n404 71.676
R1649 B.n418 B.n405 71.676
R1650 B.n414 B.n406 71.676
R1651 B.n566 B.n565 71.676
R1652 B.n856 B.n855 71.676
R1653 B.n856 B.n2 71.676
R1654 B.n128 B.n127 59.5399
R1655 B.n215 B.n125 59.5399
R1656 B.n413 B.n412 59.5399
R1657 B.n496 B.n410 59.5399
R1658 B.n571 B.n367 51.3565
R1659 B.n571 B.n363 51.3565
R1660 B.n577 B.n363 51.3565
R1661 B.n577 B.n359 51.3565
R1662 B.n583 B.n359 51.3565
R1663 B.n583 B.n355 51.3565
R1664 B.n589 B.n355 51.3565
R1665 B.n589 B.n351 51.3565
R1666 B.n595 B.n351 51.3565
R1667 B.n601 B.n347 51.3565
R1668 B.n601 B.n343 51.3565
R1669 B.n607 B.n343 51.3565
R1670 B.n607 B.n339 51.3565
R1671 B.n613 B.n339 51.3565
R1672 B.n613 B.n335 51.3565
R1673 B.n619 B.n335 51.3565
R1674 B.n619 B.n331 51.3565
R1675 B.n625 B.n331 51.3565
R1676 B.n625 B.n327 51.3565
R1677 B.n631 B.n327 51.3565
R1678 B.n631 B.n323 51.3565
R1679 B.n637 B.n323 51.3565
R1680 B.n637 B.n319 51.3565
R1681 B.n643 B.n319 51.3565
R1682 B.n649 B.n315 51.3565
R1683 B.n649 B.n311 51.3565
R1684 B.n655 B.n311 51.3565
R1685 B.n655 B.n307 51.3565
R1686 B.n661 B.n307 51.3565
R1687 B.n661 B.n303 51.3565
R1688 B.n667 B.n303 51.3565
R1689 B.n667 B.n299 51.3565
R1690 B.n673 B.n299 51.3565
R1691 B.n673 B.n295 51.3565
R1692 B.n679 B.n295 51.3565
R1693 B.n685 B.n291 51.3565
R1694 B.n685 B.n287 51.3565
R1695 B.n692 B.n287 51.3565
R1696 B.n692 B.n283 51.3565
R1697 B.n698 B.n283 51.3565
R1698 B.n698 B.n4 51.3565
R1699 B.n854 B.n4 51.3565
R1700 B.n854 B.n853 51.3565
R1701 B.n853 B.n852 51.3565
R1702 B.n852 B.n8 51.3565
R1703 B.n12 B.n8 51.3565
R1704 B.n845 B.n12 51.3565
R1705 B.n845 B.n844 51.3565
R1706 B.n844 B.n843 51.3565
R1707 B.n843 B.n16 51.3565
R1708 B.n837 B.n836 51.3565
R1709 B.n836 B.n835 51.3565
R1710 B.n835 B.n23 51.3565
R1711 B.n829 B.n23 51.3565
R1712 B.n829 B.n828 51.3565
R1713 B.n828 B.n827 51.3565
R1714 B.n827 B.n30 51.3565
R1715 B.n821 B.n30 51.3565
R1716 B.n821 B.n820 51.3565
R1717 B.n820 B.n819 51.3565
R1718 B.n819 B.n37 51.3565
R1719 B.n813 B.n812 51.3565
R1720 B.n812 B.n811 51.3565
R1721 B.n811 B.n44 51.3565
R1722 B.n805 B.n44 51.3565
R1723 B.n805 B.n804 51.3565
R1724 B.n804 B.n803 51.3565
R1725 B.n803 B.n51 51.3565
R1726 B.n797 B.n51 51.3565
R1727 B.n797 B.n796 51.3565
R1728 B.n796 B.n795 51.3565
R1729 B.n795 B.n58 51.3565
R1730 B.n789 B.n58 51.3565
R1731 B.n789 B.n788 51.3565
R1732 B.n788 B.n787 51.3565
R1733 B.n787 B.n65 51.3565
R1734 B.n781 B.n780 51.3565
R1735 B.n780 B.n779 51.3565
R1736 B.n779 B.n72 51.3565
R1737 B.n773 B.n72 51.3565
R1738 B.n773 B.n772 51.3565
R1739 B.n772 B.n771 51.3565
R1740 B.n771 B.n79 51.3565
R1741 B.n765 B.n79 51.3565
R1742 B.n765 B.n764 51.3565
R1743 B.t2 B.n315 46.0698
R1744 B.t0 B.n37 46.0698
R1745 B.n561 B.n365 33.8737
R1746 B.n568 B.n567 33.8737
R1747 B.n761 B.n760 33.8737
R1748 B.n130 B.n81 33.8737
R1749 B.t5 B.n347 32.4756
R1750 B.n679 B.t1 32.4756
R1751 B.n837 B.t3 32.4756
R1752 B.t12 B.n65 32.4756
R1753 B.n595 B.t5 18.8814
R1754 B.t1 B.n291 18.8814
R1755 B.t3 B.n16 18.8814
R1756 B.n781 B.t12 18.8814
R1757 B B.n857 18.0485
R1758 B.n573 B.n365 10.6151
R1759 B.n574 B.n573 10.6151
R1760 B.n575 B.n574 10.6151
R1761 B.n575 B.n357 10.6151
R1762 B.n585 B.n357 10.6151
R1763 B.n586 B.n585 10.6151
R1764 B.n587 B.n586 10.6151
R1765 B.n587 B.n349 10.6151
R1766 B.n597 B.n349 10.6151
R1767 B.n598 B.n597 10.6151
R1768 B.n599 B.n598 10.6151
R1769 B.n599 B.n341 10.6151
R1770 B.n609 B.n341 10.6151
R1771 B.n610 B.n609 10.6151
R1772 B.n611 B.n610 10.6151
R1773 B.n611 B.n333 10.6151
R1774 B.n621 B.n333 10.6151
R1775 B.n622 B.n621 10.6151
R1776 B.n623 B.n622 10.6151
R1777 B.n623 B.n325 10.6151
R1778 B.n633 B.n325 10.6151
R1779 B.n634 B.n633 10.6151
R1780 B.n635 B.n634 10.6151
R1781 B.n635 B.n317 10.6151
R1782 B.n645 B.n317 10.6151
R1783 B.n646 B.n645 10.6151
R1784 B.n647 B.n646 10.6151
R1785 B.n647 B.n309 10.6151
R1786 B.n657 B.n309 10.6151
R1787 B.n658 B.n657 10.6151
R1788 B.n659 B.n658 10.6151
R1789 B.n659 B.n301 10.6151
R1790 B.n669 B.n301 10.6151
R1791 B.n670 B.n669 10.6151
R1792 B.n671 B.n670 10.6151
R1793 B.n671 B.n293 10.6151
R1794 B.n681 B.n293 10.6151
R1795 B.n682 B.n681 10.6151
R1796 B.n683 B.n682 10.6151
R1797 B.n683 B.n285 10.6151
R1798 B.n694 B.n285 10.6151
R1799 B.n695 B.n694 10.6151
R1800 B.n696 B.n695 10.6151
R1801 B.n696 B.n0 10.6151
R1802 B.n561 B.n560 10.6151
R1803 B.n560 B.n559 10.6151
R1804 B.n559 B.n558 10.6151
R1805 B.n558 B.n556 10.6151
R1806 B.n556 B.n553 10.6151
R1807 B.n553 B.n552 10.6151
R1808 B.n552 B.n549 10.6151
R1809 B.n549 B.n548 10.6151
R1810 B.n548 B.n545 10.6151
R1811 B.n545 B.n544 10.6151
R1812 B.n544 B.n541 10.6151
R1813 B.n541 B.n540 10.6151
R1814 B.n540 B.n537 10.6151
R1815 B.n537 B.n536 10.6151
R1816 B.n536 B.n533 10.6151
R1817 B.n533 B.n532 10.6151
R1818 B.n532 B.n529 10.6151
R1819 B.n529 B.n528 10.6151
R1820 B.n528 B.n525 10.6151
R1821 B.n525 B.n524 10.6151
R1822 B.n524 B.n521 10.6151
R1823 B.n521 B.n520 10.6151
R1824 B.n520 B.n517 10.6151
R1825 B.n517 B.n516 10.6151
R1826 B.n516 B.n513 10.6151
R1827 B.n513 B.n512 10.6151
R1828 B.n512 B.n509 10.6151
R1829 B.n509 B.n508 10.6151
R1830 B.n508 B.n505 10.6151
R1831 B.n505 B.n504 10.6151
R1832 B.n504 B.n501 10.6151
R1833 B.n501 B.n500 10.6151
R1834 B.n500 B.n497 10.6151
R1835 B.n495 B.n492 10.6151
R1836 B.n492 B.n491 10.6151
R1837 B.n491 B.n488 10.6151
R1838 B.n488 B.n487 10.6151
R1839 B.n487 B.n484 10.6151
R1840 B.n484 B.n483 10.6151
R1841 B.n483 B.n480 10.6151
R1842 B.n480 B.n479 10.6151
R1843 B.n476 B.n475 10.6151
R1844 B.n475 B.n472 10.6151
R1845 B.n472 B.n471 10.6151
R1846 B.n471 B.n468 10.6151
R1847 B.n468 B.n467 10.6151
R1848 B.n467 B.n464 10.6151
R1849 B.n464 B.n463 10.6151
R1850 B.n463 B.n460 10.6151
R1851 B.n460 B.n459 10.6151
R1852 B.n459 B.n456 10.6151
R1853 B.n456 B.n455 10.6151
R1854 B.n455 B.n452 10.6151
R1855 B.n452 B.n451 10.6151
R1856 B.n451 B.n448 10.6151
R1857 B.n448 B.n447 10.6151
R1858 B.n447 B.n444 10.6151
R1859 B.n444 B.n443 10.6151
R1860 B.n443 B.n440 10.6151
R1861 B.n440 B.n439 10.6151
R1862 B.n439 B.n436 10.6151
R1863 B.n436 B.n435 10.6151
R1864 B.n435 B.n432 10.6151
R1865 B.n432 B.n431 10.6151
R1866 B.n431 B.n428 10.6151
R1867 B.n428 B.n427 10.6151
R1868 B.n427 B.n424 10.6151
R1869 B.n424 B.n423 10.6151
R1870 B.n423 B.n420 10.6151
R1871 B.n420 B.n419 10.6151
R1872 B.n419 B.n416 10.6151
R1873 B.n416 B.n415 10.6151
R1874 B.n415 B.n369 10.6151
R1875 B.n567 B.n369 10.6151
R1876 B.n569 B.n568 10.6151
R1877 B.n569 B.n361 10.6151
R1878 B.n579 B.n361 10.6151
R1879 B.n580 B.n579 10.6151
R1880 B.n581 B.n580 10.6151
R1881 B.n581 B.n353 10.6151
R1882 B.n591 B.n353 10.6151
R1883 B.n592 B.n591 10.6151
R1884 B.n593 B.n592 10.6151
R1885 B.n593 B.n345 10.6151
R1886 B.n603 B.n345 10.6151
R1887 B.n604 B.n603 10.6151
R1888 B.n605 B.n604 10.6151
R1889 B.n605 B.n337 10.6151
R1890 B.n615 B.n337 10.6151
R1891 B.n616 B.n615 10.6151
R1892 B.n617 B.n616 10.6151
R1893 B.n617 B.n329 10.6151
R1894 B.n627 B.n329 10.6151
R1895 B.n628 B.n627 10.6151
R1896 B.n629 B.n628 10.6151
R1897 B.n629 B.n321 10.6151
R1898 B.n639 B.n321 10.6151
R1899 B.n640 B.n639 10.6151
R1900 B.n641 B.n640 10.6151
R1901 B.n641 B.n313 10.6151
R1902 B.n651 B.n313 10.6151
R1903 B.n652 B.n651 10.6151
R1904 B.n653 B.n652 10.6151
R1905 B.n653 B.n305 10.6151
R1906 B.n663 B.n305 10.6151
R1907 B.n664 B.n663 10.6151
R1908 B.n665 B.n664 10.6151
R1909 B.n665 B.n297 10.6151
R1910 B.n675 B.n297 10.6151
R1911 B.n676 B.n675 10.6151
R1912 B.n677 B.n676 10.6151
R1913 B.n677 B.n289 10.6151
R1914 B.n687 B.n289 10.6151
R1915 B.n688 B.n687 10.6151
R1916 B.n690 B.n688 10.6151
R1917 B.n690 B.n689 10.6151
R1918 B.n689 B.n281 10.6151
R1919 B.n701 B.n281 10.6151
R1920 B.n702 B.n701 10.6151
R1921 B.n703 B.n702 10.6151
R1922 B.n704 B.n703 10.6151
R1923 B.n705 B.n704 10.6151
R1924 B.n708 B.n705 10.6151
R1925 B.n709 B.n708 10.6151
R1926 B.n710 B.n709 10.6151
R1927 B.n711 B.n710 10.6151
R1928 B.n713 B.n711 10.6151
R1929 B.n714 B.n713 10.6151
R1930 B.n715 B.n714 10.6151
R1931 B.n716 B.n715 10.6151
R1932 B.n718 B.n716 10.6151
R1933 B.n719 B.n718 10.6151
R1934 B.n720 B.n719 10.6151
R1935 B.n721 B.n720 10.6151
R1936 B.n723 B.n721 10.6151
R1937 B.n724 B.n723 10.6151
R1938 B.n725 B.n724 10.6151
R1939 B.n726 B.n725 10.6151
R1940 B.n728 B.n726 10.6151
R1941 B.n729 B.n728 10.6151
R1942 B.n730 B.n729 10.6151
R1943 B.n731 B.n730 10.6151
R1944 B.n733 B.n731 10.6151
R1945 B.n734 B.n733 10.6151
R1946 B.n735 B.n734 10.6151
R1947 B.n736 B.n735 10.6151
R1948 B.n738 B.n736 10.6151
R1949 B.n739 B.n738 10.6151
R1950 B.n740 B.n739 10.6151
R1951 B.n741 B.n740 10.6151
R1952 B.n743 B.n741 10.6151
R1953 B.n744 B.n743 10.6151
R1954 B.n745 B.n744 10.6151
R1955 B.n746 B.n745 10.6151
R1956 B.n748 B.n746 10.6151
R1957 B.n749 B.n748 10.6151
R1958 B.n750 B.n749 10.6151
R1959 B.n751 B.n750 10.6151
R1960 B.n753 B.n751 10.6151
R1961 B.n754 B.n753 10.6151
R1962 B.n755 B.n754 10.6151
R1963 B.n756 B.n755 10.6151
R1964 B.n758 B.n756 10.6151
R1965 B.n759 B.n758 10.6151
R1966 B.n760 B.n759 10.6151
R1967 B.n849 B.n1 10.6151
R1968 B.n849 B.n848 10.6151
R1969 B.n848 B.n847 10.6151
R1970 B.n847 B.n10 10.6151
R1971 B.n841 B.n10 10.6151
R1972 B.n841 B.n840 10.6151
R1973 B.n840 B.n839 10.6151
R1974 B.n839 B.n18 10.6151
R1975 B.n833 B.n18 10.6151
R1976 B.n833 B.n832 10.6151
R1977 B.n832 B.n831 10.6151
R1978 B.n831 B.n25 10.6151
R1979 B.n825 B.n25 10.6151
R1980 B.n825 B.n824 10.6151
R1981 B.n824 B.n823 10.6151
R1982 B.n823 B.n32 10.6151
R1983 B.n817 B.n32 10.6151
R1984 B.n817 B.n816 10.6151
R1985 B.n816 B.n815 10.6151
R1986 B.n815 B.n39 10.6151
R1987 B.n809 B.n39 10.6151
R1988 B.n809 B.n808 10.6151
R1989 B.n808 B.n807 10.6151
R1990 B.n807 B.n46 10.6151
R1991 B.n801 B.n46 10.6151
R1992 B.n801 B.n800 10.6151
R1993 B.n800 B.n799 10.6151
R1994 B.n799 B.n53 10.6151
R1995 B.n793 B.n53 10.6151
R1996 B.n793 B.n792 10.6151
R1997 B.n792 B.n791 10.6151
R1998 B.n791 B.n60 10.6151
R1999 B.n785 B.n60 10.6151
R2000 B.n785 B.n784 10.6151
R2001 B.n784 B.n783 10.6151
R2002 B.n783 B.n67 10.6151
R2003 B.n777 B.n67 10.6151
R2004 B.n777 B.n776 10.6151
R2005 B.n776 B.n775 10.6151
R2006 B.n775 B.n74 10.6151
R2007 B.n769 B.n74 10.6151
R2008 B.n769 B.n768 10.6151
R2009 B.n768 B.n767 10.6151
R2010 B.n767 B.n81 10.6151
R2011 B.n131 B.n130 10.6151
R2012 B.n134 B.n131 10.6151
R2013 B.n135 B.n134 10.6151
R2014 B.n138 B.n135 10.6151
R2015 B.n139 B.n138 10.6151
R2016 B.n142 B.n139 10.6151
R2017 B.n143 B.n142 10.6151
R2018 B.n146 B.n143 10.6151
R2019 B.n147 B.n146 10.6151
R2020 B.n150 B.n147 10.6151
R2021 B.n151 B.n150 10.6151
R2022 B.n154 B.n151 10.6151
R2023 B.n155 B.n154 10.6151
R2024 B.n158 B.n155 10.6151
R2025 B.n159 B.n158 10.6151
R2026 B.n162 B.n159 10.6151
R2027 B.n163 B.n162 10.6151
R2028 B.n166 B.n163 10.6151
R2029 B.n167 B.n166 10.6151
R2030 B.n170 B.n167 10.6151
R2031 B.n171 B.n170 10.6151
R2032 B.n174 B.n171 10.6151
R2033 B.n175 B.n174 10.6151
R2034 B.n178 B.n175 10.6151
R2035 B.n179 B.n178 10.6151
R2036 B.n182 B.n179 10.6151
R2037 B.n183 B.n182 10.6151
R2038 B.n186 B.n183 10.6151
R2039 B.n187 B.n186 10.6151
R2040 B.n190 B.n187 10.6151
R2041 B.n191 B.n190 10.6151
R2042 B.n194 B.n191 10.6151
R2043 B.n195 B.n194 10.6151
R2044 B.n199 B.n198 10.6151
R2045 B.n202 B.n199 10.6151
R2046 B.n203 B.n202 10.6151
R2047 B.n206 B.n203 10.6151
R2048 B.n207 B.n206 10.6151
R2049 B.n210 B.n207 10.6151
R2050 B.n211 B.n210 10.6151
R2051 B.n214 B.n211 10.6151
R2052 B.n219 B.n216 10.6151
R2053 B.n220 B.n219 10.6151
R2054 B.n223 B.n220 10.6151
R2055 B.n224 B.n223 10.6151
R2056 B.n227 B.n224 10.6151
R2057 B.n228 B.n227 10.6151
R2058 B.n231 B.n228 10.6151
R2059 B.n232 B.n231 10.6151
R2060 B.n235 B.n232 10.6151
R2061 B.n236 B.n235 10.6151
R2062 B.n239 B.n236 10.6151
R2063 B.n240 B.n239 10.6151
R2064 B.n243 B.n240 10.6151
R2065 B.n244 B.n243 10.6151
R2066 B.n247 B.n244 10.6151
R2067 B.n248 B.n247 10.6151
R2068 B.n251 B.n248 10.6151
R2069 B.n252 B.n251 10.6151
R2070 B.n255 B.n252 10.6151
R2071 B.n256 B.n255 10.6151
R2072 B.n259 B.n256 10.6151
R2073 B.n260 B.n259 10.6151
R2074 B.n263 B.n260 10.6151
R2075 B.n264 B.n263 10.6151
R2076 B.n267 B.n264 10.6151
R2077 B.n268 B.n267 10.6151
R2078 B.n271 B.n268 10.6151
R2079 B.n272 B.n271 10.6151
R2080 B.n275 B.n272 10.6151
R2081 B.n276 B.n275 10.6151
R2082 B.n279 B.n276 10.6151
R2083 B.n280 B.n279 10.6151
R2084 B.n761 B.n280 10.6151
R2085 B.n857 B.n0 8.11757
R2086 B.n857 B.n1 8.11757
R2087 B.n496 B.n495 6.5566
R2088 B.n479 B.n413 6.5566
R2089 B.n198 B.n128 6.5566
R2090 B.n215 B.n214 6.5566
R2091 B.n643 B.t2 5.28715
R2092 B.n813 B.t0 5.28715
R2093 B.n497 B.n496 4.05904
R2094 B.n476 B.n413 4.05904
R2095 B.n195 B.n128 4.05904
R2096 B.n216 B.n215 4.05904
R2097 VP.n18 VP.n0 161.3
R2098 VP.n17 VP.n16 161.3
R2099 VP.n15 VP.n1 161.3
R2100 VP.n14 VP.n13 161.3
R2101 VP.n12 VP.n2 161.3
R2102 VP.n11 VP.n10 161.3
R2103 VP.n9 VP.n3 161.3
R2104 VP.n8 VP.n7 161.3
R2105 VP.n4 VP.t2 90.7952
R2106 VP.n4 VP.t0 89.3683
R2107 VP.n6 VP.n5 63.5869
R2108 VP.n20 VP.n19 63.5869
R2109 VP.n6 VP.t1 56.9697
R2110 VP.n19 VP.t3 56.9697
R2111 VP.n13 VP.n12 56.5193
R2112 VP.n5 VP.n4 50.2067
R2113 VP.n7 VP.n3 24.4675
R2114 VP.n11 VP.n3 24.4675
R2115 VP.n12 VP.n11 24.4675
R2116 VP.n13 VP.n1 24.4675
R2117 VP.n17 VP.n1 24.4675
R2118 VP.n18 VP.n17 24.4675
R2119 VP.n7 VP.n6 18.5954
R2120 VP.n19 VP.n18 18.5954
R2121 VP.n8 VP.n5 0.417535
R2122 VP.n20 VP.n0 0.417535
R2123 VP VP.n20 0.394291
R2124 VP.n9 VP.n8 0.189894
R2125 VP.n10 VP.n9 0.189894
R2126 VP.n10 VP.n2 0.189894
R2127 VP.n14 VP.n2 0.189894
R2128 VP.n15 VP.n14 0.189894
R2129 VP.n16 VP.n15 0.189894
R2130 VP.n16 VP.n0 0.189894
R2131 VDD1 VDD1.n1 107.237
R2132 VDD1 VDD1.n0 64.0298
R2133 VDD1.n0 VDD1.t1 2.13182
R2134 VDD1.n0 VDD1.t3 2.13182
R2135 VDD1.n1 VDD1.t2 2.13182
R2136 VDD1.n1 VDD1.t0 2.13182
C0 VTAIL VP 4.23944f
C1 VP VDD2 0.479093f
C2 VP VN 6.65215f
C3 VTAIL VDD1 5.23965f
C4 VDD2 VDD1 1.35367f
C5 VN VDD1 0.15036f
C6 VP VDD1 4.31108f
C7 VTAIL VDD2 5.30278f
C8 VTAIL VN 4.22533f
C9 VDD2 VN 3.98342f
C10 VDD2 B 4.312919f
C11 VDD1 B 8.69796f
C12 VTAIL B 9.150627f
C13 VN B 13.12529f
C14 VP B 11.606611f
C15 VDD1.t1 B 0.206161f
C16 VDD1.t3 B 0.206161f
C17 VDD1.n0 B 1.80696f
C18 VDD1.t2 B 0.206161f
C19 VDD1.t0 B 0.206161f
C20 VDD1.n1 B 2.49395f
C21 VP.n0 B 0.039489f
C22 VP.t3 B 2.07094f
C23 VP.n1 B 0.039127f
C24 VP.n2 B 0.020994f
C25 VP.n3 B 0.039127f
C26 VP.t0 B 2.39567f
C27 VP.t2 B 2.40938f
C28 VP.n4 B 2.74736f
C29 VP.n5 B 1.23723f
C30 VP.t1 B 2.07094f
C31 VP.n6 B 0.824311f
C32 VP.n7 B 0.034491f
C33 VP.n8 B 0.039489f
C34 VP.n9 B 0.020994f
C35 VP.n10 B 0.020994f
C36 VP.n11 B 0.039127f
C37 VP.n12 B 0.030647f
C38 VP.n13 B 0.030647f
C39 VP.n14 B 0.020994f
C40 VP.n15 B 0.020994f
C41 VP.n16 B 0.020994f
C42 VP.n17 B 0.039127f
C43 VP.n18 B 0.034491f
C44 VP.n19 B 0.824311f
C45 VP.n20 B 0.068307f
C46 VTAIL.n0 B 0.024333f
C47 VTAIL.n1 B 0.018277f
C48 VTAIL.n2 B 0.009821f
C49 VTAIL.n3 B 0.023214f
C50 VTAIL.n4 B 0.01011f
C51 VTAIL.n5 B 0.018277f
C52 VTAIL.n6 B 0.010399f
C53 VTAIL.n7 B 0.023214f
C54 VTAIL.n8 B 0.010399f
C55 VTAIL.n9 B 0.018277f
C56 VTAIL.n10 B 0.009821f
C57 VTAIL.n11 B 0.023214f
C58 VTAIL.n12 B 0.010399f
C59 VTAIL.n13 B 0.701726f
C60 VTAIL.n14 B 0.009821f
C61 VTAIL.t3 B 0.038943f
C62 VTAIL.n15 B 0.112764f
C63 VTAIL.n16 B 0.01641f
C64 VTAIL.n17 B 0.01741f
C65 VTAIL.n18 B 0.023214f
C66 VTAIL.n19 B 0.010399f
C67 VTAIL.n20 B 0.009821f
C68 VTAIL.n21 B 0.018277f
C69 VTAIL.n22 B 0.018277f
C70 VTAIL.n23 B 0.009821f
C71 VTAIL.n24 B 0.010399f
C72 VTAIL.n25 B 0.023214f
C73 VTAIL.n26 B 0.023214f
C74 VTAIL.n27 B 0.010399f
C75 VTAIL.n28 B 0.009821f
C76 VTAIL.n29 B 0.018277f
C77 VTAIL.n30 B 0.018277f
C78 VTAIL.n31 B 0.009821f
C79 VTAIL.n32 B 0.009821f
C80 VTAIL.n33 B 0.010399f
C81 VTAIL.n34 B 0.023214f
C82 VTAIL.n35 B 0.023214f
C83 VTAIL.n36 B 0.023214f
C84 VTAIL.n37 B 0.01011f
C85 VTAIL.n38 B 0.009821f
C86 VTAIL.n39 B 0.018277f
C87 VTAIL.n40 B 0.018277f
C88 VTAIL.n41 B 0.009821f
C89 VTAIL.n42 B 0.010399f
C90 VTAIL.n43 B 0.023214f
C91 VTAIL.n44 B 0.047855f
C92 VTAIL.n45 B 0.010399f
C93 VTAIL.n46 B 0.009821f
C94 VTAIL.n47 B 0.043495f
C95 VTAIL.n48 B 0.026568f
C96 VTAIL.n49 B 0.155549f
C97 VTAIL.n50 B 0.024333f
C98 VTAIL.n51 B 0.018277f
C99 VTAIL.n52 B 0.009821f
C100 VTAIL.n53 B 0.023214f
C101 VTAIL.n54 B 0.01011f
C102 VTAIL.n55 B 0.018277f
C103 VTAIL.n56 B 0.010399f
C104 VTAIL.n57 B 0.023214f
C105 VTAIL.n58 B 0.010399f
C106 VTAIL.n59 B 0.018277f
C107 VTAIL.n60 B 0.009821f
C108 VTAIL.n61 B 0.023214f
C109 VTAIL.n62 B 0.010399f
C110 VTAIL.n63 B 0.701726f
C111 VTAIL.n64 B 0.009821f
C112 VTAIL.t4 B 0.038943f
C113 VTAIL.n65 B 0.112764f
C114 VTAIL.n66 B 0.01641f
C115 VTAIL.n67 B 0.01741f
C116 VTAIL.n68 B 0.023214f
C117 VTAIL.n69 B 0.010399f
C118 VTAIL.n70 B 0.009821f
C119 VTAIL.n71 B 0.018277f
C120 VTAIL.n72 B 0.018277f
C121 VTAIL.n73 B 0.009821f
C122 VTAIL.n74 B 0.010399f
C123 VTAIL.n75 B 0.023214f
C124 VTAIL.n76 B 0.023214f
C125 VTAIL.n77 B 0.010399f
C126 VTAIL.n78 B 0.009821f
C127 VTAIL.n79 B 0.018277f
C128 VTAIL.n80 B 0.018277f
C129 VTAIL.n81 B 0.009821f
C130 VTAIL.n82 B 0.009821f
C131 VTAIL.n83 B 0.010399f
C132 VTAIL.n84 B 0.023214f
C133 VTAIL.n85 B 0.023214f
C134 VTAIL.n86 B 0.023214f
C135 VTAIL.n87 B 0.01011f
C136 VTAIL.n88 B 0.009821f
C137 VTAIL.n89 B 0.018277f
C138 VTAIL.n90 B 0.018277f
C139 VTAIL.n91 B 0.009821f
C140 VTAIL.n92 B 0.010399f
C141 VTAIL.n93 B 0.023214f
C142 VTAIL.n94 B 0.047855f
C143 VTAIL.n95 B 0.010399f
C144 VTAIL.n96 B 0.009821f
C145 VTAIL.n97 B 0.043495f
C146 VTAIL.n98 B 0.026568f
C147 VTAIL.n99 B 0.260261f
C148 VTAIL.n100 B 0.024333f
C149 VTAIL.n101 B 0.018277f
C150 VTAIL.n102 B 0.009821f
C151 VTAIL.n103 B 0.023214f
C152 VTAIL.n104 B 0.01011f
C153 VTAIL.n105 B 0.018277f
C154 VTAIL.n106 B 0.010399f
C155 VTAIL.n107 B 0.023214f
C156 VTAIL.n108 B 0.010399f
C157 VTAIL.n109 B 0.018277f
C158 VTAIL.n110 B 0.009821f
C159 VTAIL.n111 B 0.023214f
C160 VTAIL.n112 B 0.010399f
C161 VTAIL.n113 B 0.701726f
C162 VTAIL.n114 B 0.009821f
C163 VTAIL.t6 B 0.038943f
C164 VTAIL.n115 B 0.112764f
C165 VTAIL.n116 B 0.01641f
C166 VTAIL.n117 B 0.01741f
C167 VTAIL.n118 B 0.023214f
C168 VTAIL.n119 B 0.010399f
C169 VTAIL.n120 B 0.009821f
C170 VTAIL.n121 B 0.018277f
C171 VTAIL.n122 B 0.018277f
C172 VTAIL.n123 B 0.009821f
C173 VTAIL.n124 B 0.010399f
C174 VTAIL.n125 B 0.023214f
C175 VTAIL.n126 B 0.023214f
C176 VTAIL.n127 B 0.010399f
C177 VTAIL.n128 B 0.009821f
C178 VTAIL.n129 B 0.018277f
C179 VTAIL.n130 B 0.018277f
C180 VTAIL.n131 B 0.009821f
C181 VTAIL.n132 B 0.009821f
C182 VTAIL.n133 B 0.010399f
C183 VTAIL.n134 B 0.023214f
C184 VTAIL.n135 B 0.023214f
C185 VTAIL.n136 B 0.023214f
C186 VTAIL.n137 B 0.01011f
C187 VTAIL.n138 B 0.009821f
C188 VTAIL.n139 B 0.018277f
C189 VTAIL.n140 B 0.018277f
C190 VTAIL.n141 B 0.009821f
C191 VTAIL.n142 B 0.010399f
C192 VTAIL.n143 B 0.023214f
C193 VTAIL.n144 B 0.047855f
C194 VTAIL.n145 B 0.010399f
C195 VTAIL.n146 B 0.009821f
C196 VTAIL.n147 B 0.043495f
C197 VTAIL.n148 B 0.026568f
C198 VTAIL.n149 B 1.16878f
C199 VTAIL.n150 B 0.024333f
C200 VTAIL.n151 B 0.018277f
C201 VTAIL.n152 B 0.009821f
C202 VTAIL.n153 B 0.023214f
C203 VTAIL.n154 B 0.01011f
C204 VTAIL.n155 B 0.018277f
C205 VTAIL.n156 B 0.01011f
C206 VTAIL.n157 B 0.009821f
C207 VTAIL.n158 B 0.023214f
C208 VTAIL.n159 B 0.023214f
C209 VTAIL.n160 B 0.010399f
C210 VTAIL.n161 B 0.018277f
C211 VTAIL.n162 B 0.009821f
C212 VTAIL.n163 B 0.023214f
C213 VTAIL.n164 B 0.010399f
C214 VTAIL.n165 B 0.701726f
C215 VTAIL.n166 B 0.009821f
C216 VTAIL.t2 B 0.038943f
C217 VTAIL.n167 B 0.112764f
C218 VTAIL.n168 B 0.01641f
C219 VTAIL.n169 B 0.01741f
C220 VTAIL.n170 B 0.023214f
C221 VTAIL.n171 B 0.010399f
C222 VTAIL.n172 B 0.009821f
C223 VTAIL.n173 B 0.018277f
C224 VTAIL.n174 B 0.018277f
C225 VTAIL.n175 B 0.009821f
C226 VTAIL.n176 B 0.010399f
C227 VTAIL.n177 B 0.023214f
C228 VTAIL.n178 B 0.023214f
C229 VTAIL.n179 B 0.010399f
C230 VTAIL.n180 B 0.009821f
C231 VTAIL.n181 B 0.018277f
C232 VTAIL.n182 B 0.018277f
C233 VTAIL.n183 B 0.009821f
C234 VTAIL.n184 B 0.010399f
C235 VTAIL.n185 B 0.023214f
C236 VTAIL.n186 B 0.023214f
C237 VTAIL.n187 B 0.010399f
C238 VTAIL.n188 B 0.009821f
C239 VTAIL.n189 B 0.018277f
C240 VTAIL.n190 B 0.018277f
C241 VTAIL.n191 B 0.009821f
C242 VTAIL.n192 B 0.010399f
C243 VTAIL.n193 B 0.023214f
C244 VTAIL.n194 B 0.047855f
C245 VTAIL.n195 B 0.010399f
C246 VTAIL.n196 B 0.009821f
C247 VTAIL.n197 B 0.043495f
C248 VTAIL.n198 B 0.026568f
C249 VTAIL.n199 B 1.16878f
C250 VTAIL.n200 B 0.024333f
C251 VTAIL.n201 B 0.018277f
C252 VTAIL.n202 B 0.009821f
C253 VTAIL.n203 B 0.023214f
C254 VTAIL.n204 B 0.01011f
C255 VTAIL.n205 B 0.018277f
C256 VTAIL.n206 B 0.01011f
C257 VTAIL.n207 B 0.009821f
C258 VTAIL.n208 B 0.023214f
C259 VTAIL.n209 B 0.023214f
C260 VTAIL.n210 B 0.010399f
C261 VTAIL.n211 B 0.018277f
C262 VTAIL.n212 B 0.009821f
C263 VTAIL.n213 B 0.023214f
C264 VTAIL.n214 B 0.010399f
C265 VTAIL.n215 B 0.701726f
C266 VTAIL.n216 B 0.009821f
C267 VTAIL.t1 B 0.038943f
C268 VTAIL.n217 B 0.112764f
C269 VTAIL.n218 B 0.01641f
C270 VTAIL.n219 B 0.01741f
C271 VTAIL.n220 B 0.023214f
C272 VTAIL.n221 B 0.010399f
C273 VTAIL.n222 B 0.009821f
C274 VTAIL.n223 B 0.018277f
C275 VTAIL.n224 B 0.018277f
C276 VTAIL.n225 B 0.009821f
C277 VTAIL.n226 B 0.010399f
C278 VTAIL.n227 B 0.023214f
C279 VTAIL.n228 B 0.023214f
C280 VTAIL.n229 B 0.010399f
C281 VTAIL.n230 B 0.009821f
C282 VTAIL.n231 B 0.018277f
C283 VTAIL.n232 B 0.018277f
C284 VTAIL.n233 B 0.009821f
C285 VTAIL.n234 B 0.010399f
C286 VTAIL.n235 B 0.023214f
C287 VTAIL.n236 B 0.023214f
C288 VTAIL.n237 B 0.010399f
C289 VTAIL.n238 B 0.009821f
C290 VTAIL.n239 B 0.018277f
C291 VTAIL.n240 B 0.018277f
C292 VTAIL.n241 B 0.009821f
C293 VTAIL.n242 B 0.010399f
C294 VTAIL.n243 B 0.023214f
C295 VTAIL.n244 B 0.047855f
C296 VTAIL.n245 B 0.010399f
C297 VTAIL.n246 B 0.009821f
C298 VTAIL.n247 B 0.043495f
C299 VTAIL.n248 B 0.026568f
C300 VTAIL.n249 B 0.260261f
C301 VTAIL.n250 B 0.024333f
C302 VTAIL.n251 B 0.018277f
C303 VTAIL.n252 B 0.009821f
C304 VTAIL.n253 B 0.023214f
C305 VTAIL.n254 B 0.01011f
C306 VTAIL.n255 B 0.018277f
C307 VTAIL.n256 B 0.01011f
C308 VTAIL.n257 B 0.009821f
C309 VTAIL.n258 B 0.023214f
C310 VTAIL.n259 B 0.023214f
C311 VTAIL.n260 B 0.010399f
C312 VTAIL.n261 B 0.018277f
C313 VTAIL.n262 B 0.009821f
C314 VTAIL.n263 B 0.023214f
C315 VTAIL.n264 B 0.010399f
C316 VTAIL.n265 B 0.701726f
C317 VTAIL.n266 B 0.009821f
C318 VTAIL.t5 B 0.038943f
C319 VTAIL.n267 B 0.112764f
C320 VTAIL.n268 B 0.01641f
C321 VTAIL.n269 B 0.01741f
C322 VTAIL.n270 B 0.023214f
C323 VTAIL.n271 B 0.010399f
C324 VTAIL.n272 B 0.009821f
C325 VTAIL.n273 B 0.018277f
C326 VTAIL.n274 B 0.018277f
C327 VTAIL.n275 B 0.009821f
C328 VTAIL.n276 B 0.010399f
C329 VTAIL.n277 B 0.023214f
C330 VTAIL.n278 B 0.023214f
C331 VTAIL.n279 B 0.010399f
C332 VTAIL.n280 B 0.009821f
C333 VTAIL.n281 B 0.018277f
C334 VTAIL.n282 B 0.018277f
C335 VTAIL.n283 B 0.009821f
C336 VTAIL.n284 B 0.010399f
C337 VTAIL.n285 B 0.023214f
C338 VTAIL.n286 B 0.023214f
C339 VTAIL.n287 B 0.010399f
C340 VTAIL.n288 B 0.009821f
C341 VTAIL.n289 B 0.018277f
C342 VTAIL.n290 B 0.018277f
C343 VTAIL.n291 B 0.009821f
C344 VTAIL.n292 B 0.010399f
C345 VTAIL.n293 B 0.023214f
C346 VTAIL.n294 B 0.047855f
C347 VTAIL.n295 B 0.010399f
C348 VTAIL.n296 B 0.009821f
C349 VTAIL.n297 B 0.043495f
C350 VTAIL.n298 B 0.026568f
C351 VTAIL.n299 B 0.260261f
C352 VTAIL.n300 B 0.024333f
C353 VTAIL.n301 B 0.018277f
C354 VTAIL.n302 B 0.009821f
C355 VTAIL.n303 B 0.023214f
C356 VTAIL.n304 B 0.01011f
C357 VTAIL.n305 B 0.018277f
C358 VTAIL.n306 B 0.01011f
C359 VTAIL.n307 B 0.009821f
C360 VTAIL.n308 B 0.023214f
C361 VTAIL.n309 B 0.023214f
C362 VTAIL.n310 B 0.010399f
C363 VTAIL.n311 B 0.018277f
C364 VTAIL.n312 B 0.009821f
C365 VTAIL.n313 B 0.023214f
C366 VTAIL.n314 B 0.010399f
C367 VTAIL.n315 B 0.701726f
C368 VTAIL.n316 B 0.009821f
C369 VTAIL.t7 B 0.038943f
C370 VTAIL.n317 B 0.112764f
C371 VTAIL.n318 B 0.01641f
C372 VTAIL.n319 B 0.01741f
C373 VTAIL.n320 B 0.023214f
C374 VTAIL.n321 B 0.010399f
C375 VTAIL.n322 B 0.009821f
C376 VTAIL.n323 B 0.018277f
C377 VTAIL.n324 B 0.018277f
C378 VTAIL.n325 B 0.009821f
C379 VTAIL.n326 B 0.010399f
C380 VTAIL.n327 B 0.023214f
C381 VTAIL.n328 B 0.023214f
C382 VTAIL.n329 B 0.010399f
C383 VTAIL.n330 B 0.009821f
C384 VTAIL.n331 B 0.018277f
C385 VTAIL.n332 B 0.018277f
C386 VTAIL.n333 B 0.009821f
C387 VTAIL.n334 B 0.010399f
C388 VTAIL.n335 B 0.023214f
C389 VTAIL.n336 B 0.023214f
C390 VTAIL.n337 B 0.010399f
C391 VTAIL.n338 B 0.009821f
C392 VTAIL.n339 B 0.018277f
C393 VTAIL.n340 B 0.018277f
C394 VTAIL.n341 B 0.009821f
C395 VTAIL.n342 B 0.010399f
C396 VTAIL.n343 B 0.023214f
C397 VTAIL.n344 B 0.047855f
C398 VTAIL.n345 B 0.010399f
C399 VTAIL.n346 B 0.009821f
C400 VTAIL.n347 B 0.043495f
C401 VTAIL.n348 B 0.026568f
C402 VTAIL.n349 B 1.16878f
C403 VTAIL.n350 B 0.024333f
C404 VTAIL.n351 B 0.018277f
C405 VTAIL.n352 B 0.009821f
C406 VTAIL.n353 B 0.023214f
C407 VTAIL.n354 B 0.01011f
C408 VTAIL.n355 B 0.018277f
C409 VTAIL.n356 B 0.010399f
C410 VTAIL.n357 B 0.023214f
C411 VTAIL.n358 B 0.010399f
C412 VTAIL.n359 B 0.018277f
C413 VTAIL.n360 B 0.009821f
C414 VTAIL.n361 B 0.023214f
C415 VTAIL.n362 B 0.010399f
C416 VTAIL.n363 B 0.701726f
C417 VTAIL.n364 B 0.009821f
C418 VTAIL.t0 B 0.038943f
C419 VTAIL.n365 B 0.112764f
C420 VTAIL.n366 B 0.01641f
C421 VTAIL.n367 B 0.01741f
C422 VTAIL.n368 B 0.023214f
C423 VTAIL.n369 B 0.010399f
C424 VTAIL.n370 B 0.009821f
C425 VTAIL.n371 B 0.018277f
C426 VTAIL.n372 B 0.018277f
C427 VTAIL.n373 B 0.009821f
C428 VTAIL.n374 B 0.010399f
C429 VTAIL.n375 B 0.023214f
C430 VTAIL.n376 B 0.023214f
C431 VTAIL.n377 B 0.010399f
C432 VTAIL.n378 B 0.009821f
C433 VTAIL.n379 B 0.018277f
C434 VTAIL.n380 B 0.018277f
C435 VTAIL.n381 B 0.009821f
C436 VTAIL.n382 B 0.009821f
C437 VTAIL.n383 B 0.010399f
C438 VTAIL.n384 B 0.023214f
C439 VTAIL.n385 B 0.023214f
C440 VTAIL.n386 B 0.023214f
C441 VTAIL.n387 B 0.01011f
C442 VTAIL.n388 B 0.009821f
C443 VTAIL.n389 B 0.018277f
C444 VTAIL.n390 B 0.018277f
C445 VTAIL.n391 B 0.009821f
C446 VTAIL.n392 B 0.010399f
C447 VTAIL.n393 B 0.023214f
C448 VTAIL.n394 B 0.047855f
C449 VTAIL.n395 B 0.010399f
C450 VTAIL.n396 B 0.009821f
C451 VTAIL.n397 B 0.043495f
C452 VTAIL.n398 B 0.026568f
C453 VTAIL.n399 B 1.05722f
C454 VDD2.t1 B 0.204048f
C455 VDD2.t3 B 0.204048f
C456 VDD2.n0 B 2.44145f
C457 VDD2.t2 B 0.204048f
C458 VDD2.t0 B 0.204048f
C459 VDD2.n1 B 1.78793f
C460 VDD2.n2 B 3.91954f
C461 VN.t0 B 2.35726f
C462 VN.t3 B 2.34384f
C463 VN.n0 B 1.39063f
C464 VN.t2 B 2.35726f
C465 VN.t1 B 2.34384f
C466 VN.n1 B 2.69328f
.ends

