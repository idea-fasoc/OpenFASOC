* NGSPICE file created from diff_pair_sample_0189.ext - technology: sky130A

.subckt diff_pair_sample_0189 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=2.76
X1 VDD2.t3 VN.t0 VTAIL.t5 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=5.2416 ps=27.66 w=13.44 l=2.76
X2 VDD1.t3 VP.t0 VTAIL.t3 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=5.2416 ps=27.66 w=13.44 l=2.76
X3 VDD2.t2 VN.t1 VTAIL.t4 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=5.2416 ps=27.66 w=13.44 l=2.76
X4 VDD1.t2 VP.t1 VTAIL.t2 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=2.2176 pd=13.77 as=5.2416 ps=27.66 w=13.44 l=2.76
X5 VTAIL.t6 VN.t2 VDD2.t1 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=2.2176 ps=13.77 w=13.44 l=2.76
X6 B.t8 B.t6 B.t7 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=2.76
X7 VTAIL.t7 VN.t3 VDD2.t0 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=2.2176 ps=13.77 w=13.44 l=2.76
X8 B.t5 B.t3 B.t4 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=2.76
X9 VTAIL.t1 VP.t2 VDD1.t1 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=2.2176 ps=13.77 w=13.44 l=2.76
X10 B.t2 B.t0 B.t1 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=0 ps=0 w=13.44 l=2.76
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n2824_n3656# sky130_fd_pr__pfet_01v8 ad=5.2416 pd=27.66 as=2.2176 ps=13.77 w=13.44 l=2.76
R0 B.n386 B.n111 585
R1 B.n385 B.n384 585
R2 B.n383 B.n112 585
R3 B.n382 B.n381 585
R4 B.n380 B.n113 585
R5 B.n379 B.n378 585
R6 B.n377 B.n114 585
R7 B.n376 B.n375 585
R8 B.n374 B.n115 585
R9 B.n373 B.n372 585
R10 B.n371 B.n116 585
R11 B.n370 B.n369 585
R12 B.n368 B.n117 585
R13 B.n367 B.n366 585
R14 B.n365 B.n118 585
R15 B.n364 B.n363 585
R16 B.n362 B.n119 585
R17 B.n361 B.n360 585
R18 B.n359 B.n120 585
R19 B.n358 B.n357 585
R20 B.n356 B.n121 585
R21 B.n355 B.n354 585
R22 B.n353 B.n122 585
R23 B.n352 B.n351 585
R24 B.n350 B.n123 585
R25 B.n349 B.n348 585
R26 B.n347 B.n124 585
R27 B.n346 B.n345 585
R28 B.n344 B.n125 585
R29 B.n343 B.n342 585
R30 B.n341 B.n126 585
R31 B.n340 B.n339 585
R32 B.n338 B.n127 585
R33 B.n337 B.n336 585
R34 B.n335 B.n128 585
R35 B.n334 B.n333 585
R36 B.n332 B.n129 585
R37 B.n331 B.n330 585
R38 B.n329 B.n130 585
R39 B.n328 B.n327 585
R40 B.n326 B.n131 585
R41 B.n325 B.n324 585
R42 B.n323 B.n132 585
R43 B.n322 B.n321 585
R44 B.n320 B.n133 585
R45 B.n319 B.n318 585
R46 B.n316 B.n134 585
R47 B.n315 B.n314 585
R48 B.n313 B.n137 585
R49 B.n312 B.n311 585
R50 B.n310 B.n138 585
R51 B.n309 B.n308 585
R52 B.n307 B.n139 585
R53 B.n306 B.n305 585
R54 B.n304 B.n140 585
R55 B.n302 B.n301 585
R56 B.n300 B.n143 585
R57 B.n299 B.n298 585
R58 B.n297 B.n144 585
R59 B.n296 B.n295 585
R60 B.n294 B.n145 585
R61 B.n293 B.n292 585
R62 B.n291 B.n146 585
R63 B.n290 B.n289 585
R64 B.n288 B.n147 585
R65 B.n287 B.n286 585
R66 B.n285 B.n148 585
R67 B.n284 B.n283 585
R68 B.n282 B.n149 585
R69 B.n281 B.n280 585
R70 B.n279 B.n150 585
R71 B.n278 B.n277 585
R72 B.n276 B.n151 585
R73 B.n275 B.n274 585
R74 B.n273 B.n152 585
R75 B.n272 B.n271 585
R76 B.n270 B.n153 585
R77 B.n269 B.n268 585
R78 B.n267 B.n154 585
R79 B.n266 B.n265 585
R80 B.n264 B.n155 585
R81 B.n263 B.n262 585
R82 B.n261 B.n156 585
R83 B.n260 B.n259 585
R84 B.n258 B.n157 585
R85 B.n257 B.n256 585
R86 B.n255 B.n158 585
R87 B.n254 B.n253 585
R88 B.n252 B.n159 585
R89 B.n251 B.n250 585
R90 B.n249 B.n160 585
R91 B.n248 B.n247 585
R92 B.n246 B.n161 585
R93 B.n245 B.n244 585
R94 B.n243 B.n162 585
R95 B.n242 B.n241 585
R96 B.n240 B.n163 585
R97 B.n239 B.n238 585
R98 B.n237 B.n164 585
R99 B.n236 B.n235 585
R100 B.n234 B.n165 585
R101 B.n388 B.n387 585
R102 B.n389 B.n110 585
R103 B.n391 B.n390 585
R104 B.n392 B.n109 585
R105 B.n394 B.n393 585
R106 B.n395 B.n108 585
R107 B.n397 B.n396 585
R108 B.n398 B.n107 585
R109 B.n400 B.n399 585
R110 B.n401 B.n106 585
R111 B.n403 B.n402 585
R112 B.n404 B.n105 585
R113 B.n406 B.n405 585
R114 B.n407 B.n104 585
R115 B.n409 B.n408 585
R116 B.n410 B.n103 585
R117 B.n412 B.n411 585
R118 B.n413 B.n102 585
R119 B.n415 B.n414 585
R120 B.n416 B.n101 585
R121 B.n418 B.n417 585
R122 B.n419 B.n100 585
R123 B.n421 B.n420 585
R124 B.n422 B.n99 585
R125 B.n424 B.n423 585
R126 B.n425 B.n98 585
R127 B.n427 B.n426 585
R128 B.n428 B.n97 585
R129 B.n430 B.n429 585
R130 B.n431 B.n96 585
R131 B.n433 B.n432 585
R132 B.n434 B.n95 585
R133 B.n436 B.n435 585
R134 B.n437 B.n94 585
R135 B.n439 B.n438 585
R136 B.n440 B.n93 585
R137 B.n442 B.n441 585
R138 B.n443 B.n92 585
R139 B.n445 B.n444 585
R140 B.n446 B.n91 585
R141 B.n448 B.n447 585
R142 B.n449 B.n90 585
R143 B.n451 B.n450 585
R144 B.n452 B.n89 585
R145 B.n454 B.n453 585
R146 B.n455 B.n88 585
R147 B.n457 B.n456 585
R148 B.n458 B.n87 585
R149 B.n460 B.n459 585
R150 B.n461 B.n86 585
R151 B.n463 B.n462 585
R152 B.n464 B.n85 585
R153 B.n466 B.n465 585
R154 B.n467 B.n84 585
R155 B.n469 B.n468 585
R156 B.n470 B.n83 585
R157 B.n472 B.n471 585
R158 B.n473 B.n82 585
R159 B.n475 B.n474 585
R160 B.n476 B.n81 585
R161 B.n478 B.n477 585
R162 B.n479 B.n80 585
R163 B.n481 B.n480 585
R164 B.n482 B.n79 585
R165 B.n484 B.n483 585
R166 B.n485 B.n78 585
R167 B.n487 B.n486 585
R168 B.n488 B.n77 585
R169 B.n490 B.n489 585
R170 B.n491 B.n76 585
R171 B.n493 B.n492 585
R172 B.n494 B.n75 585
R173 B.n647 B.n646 585
R174 B.n645 B.n20 585
R175 B.n644 B.n643 585
R176 B.n642 B.n21 585
R177 B.n641 B.n640 585
R178 B.n639 B.n22 585
R179 B.n638 B.n637 585
R180 B.n636 B.n23 585
R181 B.n635 B.n634 585
R182 B.n633 B.n24 585
R183 B.n632 B.n631 585
R184 B.n630 B.n25 585
R185 B.n629 B.n628 585
R186 B.n627 B.n26 585
R187 B.n626 B.n625 585
R188 B.n624 B.n27 585
R189 B.n623 B.n622 585
R190 B.n621 B.n28 585
R191 B.n620 B.n619 585
R192 B.n618 B.n29 585
R193 B.n617 B.n616 585
R194 B.n615 B.n30 585
R195 B.n614 B.n613 585
R196 B.n612 B.n31 585
R197 B.n611 B.n610 585
R198 B.n609 B.n32 585
R199 B.n608 B.n607 585
R200 B.n606 B.n33 585
R201 B.n605 B.n604 585
R202 B.n603 B.n34 585
R203 B.n602 B.n601 585
R204 B.n600 B.n35 585
R205 B.n599 B.n598 585
R206 B.n597 B.n36 585
R207 B.n596 B.n595 585
R208 B.n594 B.n37 585
R209 B.n593 B.n592 585
R210 B.n591 B.n38 585
R211 B.n590 B.n589 585
R212 B.n588 B.n39 585
R213 B.n587 B.n586 585
R214 B.n585 B.n40 585
R215 B.n584 B.n583 585
R216 B.n582 B.n41 585
R217 B.n581 B.n580 585
R218 B.n579 B.n42 585
R219 B.n578 B.n577 585
R220 B.n576 B.n43 585
R221 B.n575 B.n574 585
R222 B.n573 B.n47 585
R223 B.n572 B.n571 585
R224 B.n570 B.n48 585
R225 B.n569 B.n568 585
R226 B.n567 B.n49 585
R227 B.n566 B.n565 585
R228 B.n563 B.n50 585
R229 B.n562 B.n561 585
R230 B.n560 B.n53 585
R231 B.n559 B.n558 585
R232 B.n557 B.n54 585
R233 B.n556 B.n555 585
R234 B.n554 B.n55 585
R235 B.n553 B.n552 585
R236 B.n551 B.n56 585
R237 B.n550 B.n549 585
R238 B.n548 B.n57 585
R239 B.n547 B.n546 585
R240 B.n545 B.n58 585
R241 B.n544 B.n543 585
R242 B.n542 B.n59 585
R243 B.n541 B.n540 585
R244 B.n539 B.n60 585
R245 B.n538 B.n537 585
R246 B.n536 B.n61 585
R247 B.n535 B.n534 585
R248 B.n533 B.n62 585
R249 B.n532 B.n531 585
R250 B.n530 B.n63 585
R251 B.n529 B.n528 585
R252 B.n527 B.n64 585
R253 B.n526 B.n525 585
R254 B.n524 B.n65 585
R255 B.n523 B.n522 585
R256 B.n521 B.n66 585
R257 B.n520 B.n519 585
R258 B.n518 B.n67 585
R259 B.n517 B.n516 585
R260 B.n515 B.n68 585
R261 B.n514 B.n513 585
R262 B.n512 B.n69 585
R263 B.n511 B.n510 585
R264 B.n509 B.n70 585
R265 B.n508 B.n507 585
R266 B.n506 B.n71 585
R267 B.n505 B.n504 585
R268 B.n503 B.n72 585
R269 B.n502 B.n501 585
R270 B.n500 B.n73 585
R271 B.n499 B.n498 585
R272 B.n497 B.n74 585
R273 B.n496 B.n495 585
R274 B.n648 B.n19 585
R275 B.n650 B.n649 585
R276 B.n651 B.n18 585
R277 B.n653 B.n652 585
R278 B.n654 B.n17 585
R279 B.n656 B.n655 585
R280 B.n657 B.n16 585
R281 B.n659 B.n658 585
R282 B.n660 B.n15 585
R283 B.n662 B.n661 585
R284 B.n663 B.n14 585
R285 B.n665 B.n664 585
R286 B.n666 B.n13 585
R287 B.n668 B.n667 585
R288 B.n669 B.n12 585
R289 B.n671 B.n670 585
R290 B.n672 B.n11 585
R291 B.n674 B.n673 585
R292 B.n675 B.n10 585
R293 B.n677 B.n676 585
R294 B.n678 B.n9 585
R295 B.n680 B.n679 585
R296 B.n681 B.n8 585
R297 B.n683 B.n682 585
R298 B.n684 B.n7 585
R299 B.n686 B.n685 585
R300 B.n687 B.n6 585
R301 B.n689 B.n688 585
R302 B.n690 B.n5 585
R303 B.n692 B.n691 585
R304 B.n693 B.n4 585
R305 B.n695 B.n694 585
R306 B.n696 B.n3 585
R307 B.n698 B.n697 585
R308 B.n699 B.n0 585
R309 B.n2 B.n1 585
R310 B.n183 B.n182 585
R311 B.n185 B.n184 585
R312 B.n186 B.n181 585
R313 B.n188 B.n187 585
R314 B.n189 B.n180 585
R315 B.n191 B.n190 585
R316 B.n192 B.n179 585
R317 B.n194 B.n193 585
R318 B.n195 B.n178 585
R319 B.n197 B.n196 585
R320 B.n198 B.n177 585
R321 B.n200 B.n199 585
R322 B.n201 B.n176 585
R323 B.n203 B.n202 585
R324 B.n204 B.n175 585
R325 B.n206 B.n205 585
R326 B.n207 B.n174 585
R327 B.n209 B.n208 585
R328 B.n210 B.n173 585
R329 B.n212 B.n211 585
R330 B.n213 B.n172 585
R331 B.n215 B.n214 585
R332 B.n216 B.n171 585
R333 B.n218 B.n217 585
R334 B.n219 B.n170 585
R335 B.n221 B.n220 585
R336 B.n222 B.n169 585
R337 B.n224 B.n223 585
R338 B.n225 B.n168 585
R339 B.n227 B.n226 585
R340 B.n228 B.n167 585
R341 B.n230 B.n229 585
R342 B.n231 B.n166 585
R343 B.n233 B.n232 585
R344 B.n234 B.n233 502.111
R345 B.n387 B.n386 502.111
R346 B.n495 B.n494 502.111
R347 B.n646 B.n19 502.111
R348 B.n135 B.t1 461.503
R349 B.n51 B.t8 461.503
R350 B.n141 B.t10 461.503
R351 B.n44 B.t5 461.503
R352 B.n136 B.t2 401.575
R353 B.n52 B.t7 401.575
R354 B.n142 B.t11 401.575
R355 B.n45 B.t4 401.575
R356 B.n141 B.t9 325.632
R357 B.n135 B.t0 325.632
R358 B.n51 B.t6 325.632
R359 B.n44 B.t3 325.632
R360 B.n701 B.n700 256.663
R361 B.n700 B.n699 235.042
R362 B.n700 B.n2 235.042
R363 B.n235 B.n234 163.367
R364 B.n235 B.n164 163.367
R365 B.n239 B.n164 163.367
R366 B.n240 B.n239 163.367
R367 B.n241 B.n240 163.367
R368 B.n241 B.n162 163.367
R369 B.n245 B.n162 163.367
R370 B.n246 B.n245 163.367
R371 B.n247 B.n246 163.367
R372 B.n247 B.n160 163.367
R373 B.n251 B.n160 163.367
R374 B.n252 B.n251 163.367
R375 B.n253 B.n252 163.367
R376 B.n253 B.n158 163.367
R377 B.n257 B.n158 163.367
R378 B.n258 B.n257 163.367
R379 B.n259 B.n258 163.367
R380 B.n259 B.n156 163.367
R381 B.n263 B.n156 163.367
R382 B.n264 B.n263 163.367
R383 B.n265 B.n264 163.367
R384 B.n265 B.n154 163.367
R385 B.n269 B.n154 163.367
R386 B.n270 B.n269 163.367
R387 B.n271 B.n270 163.367
R388 B.n271 B.n152 163.367
R389 B.n275 B.n152 163.367
R390 B.n276 B.n275 163.367
R391 B.n277 B.n276 163.367
R392 B.n277 B.n150 163.367
R393 B.n281 B.n150 163.367
R394 B.n282 B.n281 163.367
R395 B.n283 B.n282 163.367
R396 B.n283 B.n148 163.367
R397 B.n287 B.n148 163.367
R398 B.n288 B.n287 163.367
R399 B.n289 B.n288 163.367
R400 B.n289 B.n146 163.367
R401 B.n293 B.n146 163.367
R402 B.n294 B.n293 163.367
R403 B.n295 B.n294 163.367
R404 B.n295 B.n144 163.367
R405 B.n299 B.n144 163.367
R406 B.n300 B.n299 163.367
R407 B.n301 B.n300 163.367
R408 B.n301 B.n140 163.367
R409 B.n306 B.n140 163.367
R410 B.n307 B.n306 163.367
R411 B.n308 B.n307 163.367
R412 B.n308 B.n138 163.367
R413 B.n312 B.n138 163.367
R414 B.n313 B.n312 163.367
R415 B.n314 B.n313 163.367
R416 B.n314 B.n134 163.367
R417 B.n319 B.n134 163.367
R418 B.n320 B.n319 163.367
R419 B.n321 B.n320 163.367
R420 B.n321 B.n132 163.367
R421 B.n325 B.n132 163.367
R422 B.n326 B.n325 163.367
R423 B.n327 B.n326 163.367
R424 B.n327 B.n130 163.367
R425 B.n331 B.n130 163.367
R426 B.n332 B.n331 163.367
R427 B.n333 B.n332 163.367
R428 B.n333 B.n128 163.367
R429 B.n337 B.n128 163.367
R430 B.n338 B.n337 163.367
R431 B.n339 B.n338 163.367
R432 B.n339 B.n126 163.367
R433 B.n343 B.n126 163.367
R434 B.n344 B.n343 163.367
R435 B.n345 B.n344 163.367
R436 B.n345 B.n124 163.367
R437 B.n349 B.n124 163.367
R438 B.n350 B.n349 163.367
R439 B.n351 B.n350 163.367
R440 B.n351 B.n122 163.367
R441 B.n355 B.n122 163.367
R442 B.n356 B.n355 163.367
R443 B.n357 B.n356 163.367
R444 B.n357 B.n120 163.367
R445 B.n361 B.n120 163.367
R446 B.n362 B.n361 163.367
R447 B.n363 B.n362 163.367
R448 B.n363 B.n118 163.367
R449 B.n367 B.n118 163.367
R450 B.n368 B.n367 163.367
R451 B.n369 B.n368 163.367
R452 B.n369 B.n116 163.367
R453 B.n373 B.n116 163.367
R454 B.n374 B.n373 163.367
R455 B.n375 B.n374 163.367
R456 B.n375 B.n114 163.367
R457 B.n379 B.n114 163.367
R458 B.n380 B.n379 163.367
R459 B.n381 B.n380 163.367
R460 B.n381 B.n112 163.367
R461 B.n385 B.n112 163.367
R462 B.n386 B.n385 163.367
R463 B.n494 B.n493 163.367
R464 B.n493 B.n76 163.367
R465 B.n489 B.n76 163.367
R466 B.n489 B.n488 163.367
R467 B.n488 B.n487 163.367
R468 B.n487 B.n78 163.367
R469 B.n483 B.n78 163.367
R470 B.n483 B.n482 163.367
R471 B.n482 B.n481 163.367
R472 B.n481 B.n80 163.367
R473 B.n477 B.n80 163.367
R474 B.n477 B.n476 163.367
R475 B.n476 B.n475 163.367
R476 B.n475 B.n82 163.367
R477 B.n471 B.n82 163.367
R478 B.n471 B.n470 163.367
R479 B.n470 B.n469 163.367
R480 B.n469 B.n84 163.367
R481 B.n465 B.n84 163.367
R482 B.n465 B.n464 163.367
R483 B.n464 B.n463 163.367
R484 B.n463 B.n86 163.367
R485 B.n459 B.n86 163.367
R486 B.n459 B.n458 163.367
R487 B.n458 B.n457 163.367
R488 B.n457 B.n88 163.367
R489 B.n453 B.n88 163.367
R490 B.n453 B.n452 163.367
R491 B.n452 B.n451 163.367
R492 B.n451 B.n90 163.367
R493 B.n447 B.n90 163.367
R494 B.n447 B.n446 163.367
R495 B.n446 B.n445 163.367
R496 B.n445 B.n92 163.367
R497 B.n441 B.n92 163.367
R498 B.n441 B.n440 163.367
R499 B.n440 B.n439 163.367
R500 B.n439 B.n94 163.367
R501 B.n435 B.n94 163.367
R502 B.n435 B.n434 163.367
R503 B.n434 B.n433 163.367
R504 B.n433 B.n96 163.367
R505 B.n429 B.n96 163.367
R506 B.n429 B.n428 163.367
R507 B.n428 B.n427 163.367
R508 B.n427 B.n98 163.367
R509 B.n423 B.n98 163.367
R510 B.n423 B.n422 163.367
R511 B.n422 B.n421 163.367
R512 B.n421 B.n100 163.367
R513 B.n417 B.n100 163.367
R514 B.n417 B.n416 163.367
R515 B.n416 B.n415 163.367
R516 B.n415 B.n102 163.367
R517 B.n411 B.n102 163.367
R518 B.n411 B.n410 163.367
R519 B.n410 B.n409 163.367
R520 B.n409 B.n104 163.367
R521 B.n405 B.n104 163.367
R522 B.n405 B.n404 163.367
R523 B.n404 B.n403 163.367
R524 B.n403 B.n106 163.367
R525 B.n399 B.n106 163.367
R526 B.n399 B.n398 163.367
R527 B.n398 B.n397 163.367
R528 B.n397 B.n108 163.367
R529 B.n393 B.n108 163.367
R530 B.n393 B.n392 163.367
R531 B.n392 B.n391 163.367
R532 B.n391 B.n110 163.367
R533 B.n387 B.n110 163.367
R534 B.n646 B.n645 163.367
R535 B.n645 B.n644 163.367
R536 B.n644 B.n21 163.367
R537 B.n640 B.n21 163.367
R538 B.n640 B.n639 163.367
R539 B.n639 B.n638 163.367
R540 B.n638 B.n23 163.367
R541 B.n634 B.n23 163.367
R542 B.n634 B.n633 163.367
R543 B.n633 B.n632 163.367
R544 B.n632 B.n25 163.367
R545 B.n628 B.n25 163.367
R546 B.n628 B.n627 163.367
R547 B.n627 B.n626 163.367
R548 B.n626 B.n27 163.367
R549 B.n622 B.n27 163.367
R550 B.n622 B.n621 163.367
R551 B.n621 B.n620 163.367
R552 B.n620 B.n29 163.367
R553 B.n616 B.n29 163.367
R554 B.n616 B.n615 163.367
R555 B.n615 B.n614 163.367
R556 B.n614 B.n31 163.367
R557 B.n610 B.n31 163.367
R558 B.n610 B.n609 163.367
R559 B.n609 B.n608 163.367
R560 B.n608 B.n33 163.367
R561 B.n604 B.n33 163.367
R562 B.n604 B.n603 163.367
R563 B.n603 B.n602 163.367
R564 B.n602 B.n35 163.367
R565 B.n598 B.n35 163.367
R566 B.n598 B.n597 163.367
R567 B.n597 B.n596 163.367
R568 B.n596 B.n37 163.367
R569 B.n592 B.n37 163.367
R570 B.n592 B.n591 163.367
R571 B.n591 B.n590 163.367
R572 B.n590 B.n39 163.367
R573 B.n586 B.n39 163.367
R574 B.n586 B.n585 163.367
R575 B.n585 B.n584 163.367
R576 B.n584 B.n41 163.367
R577 B.n580 B.n41 163.367
R578 B.n580 B.n579 163.367
R579 B.n579 B.n578 163.367
R580 B.n578 B.n43 163.367
R581 B.n574 B.n43 163.367
R582 B.n574 B.n573 163.367
R583 B.n573 B.n572 163.367
R584 B.n572 B.n48 163.367
R585 B.n568 B.n48 163.367
R586 B.n568 B.n567 163.367
R587 B.n567 B.n566 163.367
R588 B.n566 B.n50 163.367
R589 B.n561 B.n50 163.367
R590 B.n561 B.n560 163.367
R591 B.n560 B.n559 163.367
R592 B.n559 B.n54 163.367
R593 B.n555 B.n54 163.367
R594 B.n555 B.n554 163.367
R595 B.n554 B.n553 163.367
R596 B.n553 B.n56 163.367
R597 B.n549 B.n56 163.367
R598 B.n549 B.n548 163.367
R599 B.n548 B.n547 163.367
R600 B.n547 B.n58 163.367
R601 B.n543 B.n58 163.367
R602 B.n543 B.n542 163.367
R603 B.n542 B.n541 163.367
R604 B.n541 B.n60 163.367
R605 B.n537 B.n60 163.367
R606 B.n537 B.n536 163.367
R607 B.n536 B.n535 163.367
R608 B.n535 B.n62 163.367
R609 B.n531 B.n62 163.367
R610 B.n531 B.n530 163.367
R611 B.n530 B.n529 163.367
R612 B.n529 B.n64 163.367
R613 B.n525 B.n64 163.367
R614 B.n525 B.n524 163.367
R615 B.n524 B.n523 163.367
R616 B.n523 B.n66 163.367
R617 B.n519 B.n66 163.367
R618 B.n519 B.n518 163.367
R619 B.n518 B.n517 163.367
R620 B.n517 B.n68 163.367
R621 B.n513 B.n68 163.367
R622 B.n513 B.n512 163.367
R623 B.n512 B.n511 163.367
R624 B.n511 B.n70 163.367
R625 B.n507 B.n70 163.367
R626 B.n507 B.n506 163.367
R627 B.n506 B.n505 163.367
R628 B.n505 B.n72 163.367
R629 B.n501 B.n72 163.367
R630 B.n501 B.n500 163.367
R631 B.n500 B.n499 163.367
R632 B.n499 B.n74 163.367
R633 B.n495 B.n74 163.367
R634 B.n650 B.n19 163.367
R635 B.n651 B.n650 163.367
R636 B.n652 B.n651 163.367
R637 B.n652 B.n17 163.367
R638 B.n656 B.n17 163.367
R639 B.n657 B.n656 163.367
R640 B.n658 B.n657 163.367
R641 B.n658 B.n15 163.367
R642 B.n662 B.n15 163.367
R643 B.n663 B.n662 163.367
R644 B.n664 B.n663 163.367
R645 B.n664 B.n13 163.367
R646 B.n668 B.n13 163.367
R647 B.n669 B.n668 163.367
R648 B.n670 B.n669 163.367
R649 B.n670 B.n11 163.367
R650 B.n674 B.n11 163.367
R651 B.n675 B.n674 163.367
R652 B.n676 B.n675 163.367
R653 B.n676 B.n9 163.367
R654 B.n680 B.n9 163.367
R655 B.n681 B.n680 163.367
R656 B.n682 B.n681 163.367
R657 B.n682 B.n7 163.367
R658 B.n686 B.n7 163.367
R659 B.n687 B.n686 163.367
R660 B.n688 B.n687 163.367
R661 B.n688 B.n5 163.367
R662 B.n692 B.n5 163.367
R663 B.n693 B.n692 163.367
R664 B.n694 B.n693 163.367
R665 B.n694 B.n3 163.367
R666 B.n698 B.n3 163.367
R667 B.n699 B.n698 163.367
R668 B.n182 B.n2 163.367
R669 B.n185 B.n182 163.367
R670 B.n186 B.n185 163.367
R671 B.n187 B.n186 163.367
R672 B.n187 B.n180 163.367
R673 B.n191 B.n180 163.367
R674 B.n192 B.n191 163.367
R675 B.n193 B.n192 163.367
R676 B.n193 B.n178 163.367
R677 B.n197 B.n178 163.367
R678 B.n198 B.n197 163.367
R679 B.n199 B.n198 163.367
R680 B.n199 B.n176 163.367
R681 B.n203 B.n176 163.367
R682 B.n204 B.n203 163.367
R683 B.n205 B.n204 163.367
R684 B.n205 B.n174 163.367
R685 B.n209 B.n174 163.367
R686 B.n210 B.n209 163.367
R687 B.n211 B.n210 163.367
R688 B.n211 B.n172 163.367
R689 B.n215 B.n172 163.367
R690 B.n216 B.n215 163.367
R691 B.n217 B.n216 163.367
R692 B.n217 B.n170 163.367
R693 B.n221 B.n170 163.367
R694 B.n222 B.n221 163.367
R695 B.n223 B.n222 163.367
R696 B.n223 B.n168 163.367
R697 B.n227 B.n168 163.367
R698 B.n228 B.n227 163.367
R699 B.n229 B.n228 163.367
R700 B.n229 B.n166 163.367
R701 B.n233 B.n166 163.367
R702 B.n142 B.n141 59.9278
R703 B.n136 B.n135 59.9278
R704 B.n52 B.n51 59.9278
R705 B.n45 B.n44 59.9278
R706 B.n303 B.n142 59.5399
R707 B.n317 B.n136 59.5399
R708 B.n564 B.n52 59.5399
R709 B.n46 B.n45 59.5399
R710 B.n648 B.n647 32.6249
R711 B.n496 B.n75 32.6249
R712 B.n388 B.n111 32.6249
R713 B.n232 B.n165 32.6249
R714 B B.n701 18.0485
R715 B.n649 B.n648 10.6151
R716 B.n649 B.n18 10.6151
R717 B.n653 B.n18 10.6151
R718 B.n654 B.n653 10.6151
R719 B.n655 B.n654 10.6151
R720 B.n655 B.n16 10.6151
R721 B.n659 B.n16 10.6151
R722 B.n660 B.n659 10.6151
R723 B.n661 B.n660 10.6151
R724 B.n661 B.n14 10.6151
R725 B.n665 B.n14 10.6151
R726 B.n666 B.n665 10.6151
R727 B.n667 B.n666 10.6151
R728 B.n667 B.n12 10.6151
R729 B.n671 B.n12 10.6151
R730 B.n672 B.n671 10.6151
R731 B.n673 B.n672 10.6151
R732 B.n673 B.n10 10.6151
R733 B.n677 B.n10 10.6151
R734 B.n678 B.n677 10.6151
R735 B.n679 B.n678 10.6151
R736 B.n679 B.n8 10.6151
R737 B.n683 B.n8 10.6151
R738 B.n684 B.n683 10.6151
R739 B.n685 B.n684 10.6151
R740 B.n685 B.n6 10.6151
R741 B.n689 B.n6 10.6151
R742 B.n690 B.n689 10.6151
R743 B.n691 B.n690 10.6151
R744 B.n691 B.n4 10.6151
R745 B.n695 B.n4 10.6151
R746 B.n696 B.n695 10.6151
R747 B.n697 B.n696 10.6151
R748 B.n697 B.n0 10.6151
R749 B.n647 B.n20 10.6151
R750 B.n643 B.n20 10.6151
R751 B.n643 B.n642 10.6151
R752 B.n642 B.n641 10.6151
R753 B.n641 B.n22 10.6151
R754 B.n637 B.n22 10.6151
R755 B.n637 B.n636 10.6151
R756 B.n636 B.n635 10.6151
R757 B.n635 B.n24 10.6151
R758 B.n631 B.n24 10.6151
R759 B.n631 B.n630 10.6151
R760 B.n630 B.n629 10.6151
R761 B.n629 B.n26 10.6151
R762 B.n625 B.n26 10.6151
R763 B.n625 B.n624 10.6151
R764 B.n624 B.n623 10.6151
R765 B.n623 B.n28 10.6151
R766 B.n619 B.n28 10.6151
R767 B.n619 B.n618 10.6151
R768 B.n618 B.n617 10.6151
R769 B.n617 B.n30 10.6151
R770 B.n613 B.n30 10.6151
R771 B.n613 B.n612 10.6151
R772 B.n612 B.n611 10.6151
R773 B.n611 B.n32 10.6151
R774 B.n607 B.n32 10.6151
R775 B.n607 B.n606 10.6151
R776 B.n606 B.n605 10.6151
R777 B.n605 B.n34 10.6151
R778 B.n601 B.n34 10.6151
R779 B.n601 B.n600 10.6151
R780 B.n600 B.n599 10.6151
R781 B.n599 B.n36 10.6151
R782 B.n595 B.n36 10.6151
R783 B.n595 B.n594 10.6151
R784 B.n594 B.n593 10.6151
R785 B.n593 B.n38 10.6151
R786 B.n589 B.n38 10.6151
R787 B.n589 B.n588 10.6151
R788 B.n588 B.n587 10.6151
R789 B.n587 B.n40 10.6151
R790 B.n583 B.n40 10.6151
R791 B.n583 B.n582 10.6151
R792 B.n582 B.n581 10.6151
R793 B.n581 B.n42 10.6151
R794 B.n577 B.n576 10.6151
R795 B.n576 B.n575 10.6151
R796 B.n575 B.n47 10.6151
R797 B.n571 B.n47 10.6151
R798 B.n571 B.n570 10.6151
R799 B.n570 B.n569 10.6151
R800 B.n569 B.n49 10.6151
R801 B.n565 B.n49 10.6151
R802 B.n563 B.n562 10.6151
R803 B.n562 B.n53 10.6151
R804 B.n558 B.n53 10.6151
R805 B.n558 B.n557 10.6151
R806 B.n557 B.n556 10.6151
R807 B.n556 B.n55 10.6151
R808 B.n552 B.n55 10.6151
R809 B.n552 B.n551 10.6151
R810 B.n551 B.n550 10.6151
R811 B.n550 B.n57 10.6151
R812 B.n546 B.n57 10.6151
R813 B.n546 B.n545 10.6151
R814 B.n545 B.n544 10.6151
R815 B.n544 B.n59 10.6151
R816 B.n540 B.n59 10.6151
R817 B.n540 B.n539 10.6151
R818 B.n539 B.n538 10.6151
R819 B.n538 B.n61 10.6151
R820 B.n534 B.n61 10.6151
R821 B.n534 B.n533 10.6151
R822 B.n533 B.n532 10.6151
R823 B.n532 B.n63 10.6151
R824 B.n528 B.n63 10.6151
R825 B.n528 B.n527 10.6151
R826 B.n527 B.n526 10.6151
R827 B.n526 B.n65 10.6151
R828 B.n522 B.n65 10.6151
R829 B.n522 B.n521 10.6151
R830 B.n521 B.n520 10.6151
R831 B.n520 B.n67 10.6151
R832 B.n516 B.n67 10.6151
R833 B.n516 B.n515 10.6151
R834 B.n515 B.n514 10.6151
R835 B.n514 B.n69 10.6151
R836 B.n510 B.n69 10.6151
R837 B.n510 B.n509 10.6151
R838 B.n509 B.n508 10.6151
R839 B.n508 B.n71 10.6151
R840 B.n504 B.n71 10.6151
R841 B.n504 B.n503 10.6151
R842 B.n503 B.n502 10.6151
R843 B.n502 B.n73 10.6151
R844 B.n498 B.n73 10.6151
R845 B.n498 B.n497 10.6151
R846 B.n497 B.n496 10.6151
R847 B.n492 B.n75 10.6151
R848 B.n492 B.n491 10.6151
R849 B.n491 B.n490 10.6151
R850 B.n490 B.n77 10.6151
R851 B.n486 B.n77 10.6151
R852 B.n486 B.n485 10.6151
R853 B.n485 B.n484 10.6151
R854 B.n484 B.n79 10.6151
R855 B.n480 B.n79 10.6151
R856 B.n480 B.n479 10.6151
R857 B.n479 B.n478 10.6151
R858 B.n478 B.n81 10.6151
R859 B.n474 B.n81 10.6151
R860 B.n474 B.n473 10.6151
R861 B.n473 B.n472 10.6151
R862 B.n472 B.n83 10.6151
R863 B.n468 B.n83 10.6151
R864 B.n468 B.n467 10.6151
R865 B.n467 B.n466 10.6151
R866 B.n466 B.n85 10.6151
R867 B.n462 B.n85 10.6151
R868 B.n462 B.n461 10.6151
R869 B.n461 B.n460 10.6151
R870 B.n460 B.n87 10.6151
R871 B.n456 B.n87 10.6151
R872 B.n456 B.n455 10.6151
R873 B.n455 B.n454 10.6151
R874 B.n454 B.n89 10.6151
R875 B.n450 B.n89 10.6151
R876 B.n450 B.n449 10.6151
R877 B.n449 B.n448 10.6151
R878 B.n448 B.n91 10.6151
R879 B.n444 B.n91 10.6151
R880 B.n444 B.n443 10.6151
R881 B.n443 B.n442 10.6151
R882 B.n442 B.n93 10.6151
R883 B.n438 B.n93 10.6151
R884 B.n438 B.n437 10.6151
R885 B.n437 B.n436 10.6151
R886 B.n436 B.n95 10.6151
R887 B.n432 B.n95 10.6151
R888 B.n432 B.n431 10.6151
R889 B.n431 B.n430 10.6151
R890 B.n430 B.n97 10.6151
R891 B.n426 B.n97 10.6151
R892 B.n426 B.n425 10.6151
R893 B.n425 B.n424 10.6151
R894 B.n424 B.n99 10.6151
R895 B.n420 B.n99 10.6151
R896 B.n420 B.n419 10.6151
R897 B.n419 B.n418 10.6151
R898 B.n418 B.n101 10.6151
R899 B.n414 B.n101 10.6151
R900 B.n414 B.n413 10.6151
R901 B.n413 B.n412 10.6151
R902 B.n412 B.n103 10.6151
R903 B.n408 B.n103 10.6151
R904 B.n408 B.n407 10.6151
R905 B.n407 B.n406 10.6151
R906 B.n406 B.n105 10.6151
R907 B.n402 B.n105 10.6151
R908 B.n402 B.n401 10.6151
R909 B.n401 B.n400 10.6151
R910 B.n400 B.n107 10.6151
R911 B.n396 B.n107 10.6151
R912 B.n396 B.n395 10.6151
R913 B.n395 B.n394 10.6151
R914 B.n394 B.n109 10.6151
R915 B.n390 B.n109 10.6151
R916 B.n390 B.n389 10.6151
R917 B.n389 B.n388 10.6151
R918 B.n183 B.n1 10.6151
R919 B.n184 B.n183 10.6151
R920 B.n184 B.n181 10.6151
R921 B.n188 B.n181 10.6151
R922 B.n189 B.n188 10.6151
R923 B.n190 B.n189 10.6151
R924 B.n190 B.n179 10.6151
R925 B.n194 B.n179 10.6151
R926 B.n195 B.n194 10.6151
R927 B.n196 B.n195 10.6151
R928 B.n196 B.n177 10.6151
R929 B.n200 B.n177 10.6151
R930 B.n201 B.n200 10.6151
R931 B.n202 B.n201 10.6151
R932 B.n202 B.n175 10.6151
R933 B.n206 B.n175 10.6151
R934 B.n207 B.n206 10.6151
R935 B.n208 B.n207 10.6151
R936 B.n208 B.n173 10.6151
R937 B.n212 B.n173 10.6151
R938 B.n213 B.n212 10.6151
R939 B.n214 B.n213 10.6151
R940 B.n214 B.n171 10.6151
R941 B.n218 B.n171 10.6151
R942 B.n219 B.n218 10.6151
R943 B.n220 B.n219 10.6151
R944 B.n220 B.n169 10.6151
R945 B.n224 B.n169 10.6151
R946 B.n225 B.n224 10.6151
R947 B.n226 B.n225 10.6151
R948 B.n226 B.n167 10.6151
R949 B.n230 B.n167 10.6151
R950 B.n231 B.n230 10.6151
R951 B.n232 B.n231 10.6151
R952 B.n236 B.n165 10.6151
R953 B.n237 B.n236 10.6151
R954 B.n238 B.n237 10.6151
R955 B.n238 B.n163 10.6151
R956 B.n242 B.n163 10.6151
R957 B.n243 B.n242 10.6151
R958 B.n244 B.n243 10.6151
R959 B.n244 B.n161 10.6151
R960 B.n248 B.n161 10.6151
R961 B.n249 B.n248 10.6151
R962 B.n250 B.n249 10.6151
R963 B.n250 B.n159 10.6151
R964 B.n254 B.n159 10.6151
R965 B.n255 B.n254 10.6151
R966 B.n256 B.n255 10.6151
R967 B.n256 B.n157 10.6151
R968 B.n260 B.n157 10.6151
R969 B.n261 B.n260 10.6151
R970 B.n262 B.n261 10.6151
R971 B.n262 B.n155 10.6151
R972 B.n266 B.n155 10.6151
R973 B.n267 B.n266 10.6151
R974 B.n268 B.n267 10.6151
R975 B.n268 B.n153 10.6151
R976 B.n272 B.n153 10.6151
R977 B.n273 B.n272 10.6151
R978 B.n274 B.n273 10.6151
R979 B.n274 B.n151 10.6151
R980 B.n278 B.n151 10.6151
R981 B.n279 B.n278 10.6151
R982 B.n280 B.n279 10.6151
R983 B.n280 B.n149 10.6151
R984 B.n284 B.n149 10.6151
R985 B.n285 B.n284 10.6151
R986 B.n286 B.n285 10.6151
R987 B.n286 B.n147 10.6151
R988 B.n290 B.n147 10.6151
R989 B.n291 B.n290 10.6151
R990 B.n292 B.n291 10.6151
R991 B.n292 B.n145 10.6151
R992 B.n296 B.n145 10.6151
R993 B.n297 B.n296 10.6151
R994 B.n298 B.n297 10.6151
R995 B.n298 B.n143 10.6151
R996 B.n302 B.n143 10.6151
R997 B.n305 B.n304 10.6151
R998 B.n305 B.n139 10.6151
R999 B.n309 B.n139 10.6151
R1000 B.n310 B.n309 10.6151
R1001 B.n311 B.n310 10.6151
R1002 B.n311 B.n137 10.6151
R1003 B.n315 B.n137 10.6151
R1004 B.n316 B.n315 10.6151
R1005 B.n318 B.n133 10.6151
R1006 B.n322 B.n133 10.6151
R1007 B.n323 B.n322 10.6151
R1008 B.n324 B.n323 10.6151
R1009 B.n324 B.n131 10.6151
R1010 B.n328 B.n131 10.6151
R1011 B.n329 B.n328 10.6151
R1012 B.n330 B.n329 10.6151
R1013 B.n330 B.n129 10.6151
R1014 B.n334 B.n129 10.6151
R1015 B.n335 B.n334 10.6151
R1016 B.n336 B.n335 10.6151
R1017 B.n336 B.n127 10.6151
R1018 B.n340 B.n127 10.6151
R1019 B.n341 B.n340 10.6151
R1020 B.n342 B.n341 10.6151
R1021 B.n342 B.n125 10.6151
R1022 B.n346 B.n125 10.6151
R1023 B.n347 B.n346 10.6151
R1024 B.n348 B.n347 10.6151
R1025 B.n348 B.n123 10.6151
R1026 B.n352 B.n123 10.6151
R1027 B.n353 B.n352 10.6151
R1028 B.n354 B.n353 10.6151
R1029 B.n354 B.n121 10.6151
R1030 B.n358 B.n121 10.6151
R1031 B.n359 B.n358 10.6151
R1032 B.n360 B.n359 10.6151
R1033 B.n360 B.n119 10.6151
R1034 B.n364 B.n119 10.6151
R1035 B.n365 B.n364 10.6151
R1036 B.n366 B.n365 10.6151
R1037 B.n366 B.n117 10.6151
R1038 B.n370 B.n117 10.6151
R1039 B.n371 B.n370 10.6151
R1040 B.n372 B.n371 10.6151
R1041 B.n372 B.n115 10.6151
R1042 B.n376 B.n115 10.6151
R1043 B.n377 B.n376 10.6151
R1044 B.n378 B.n377 10.6151
R1045 B.n378 B.n113 10.6151
R1046 B.n382 B.n113 10.6151
R1047 B.n383 B.n382 10.6151
R1048 B.n384 B.n383 10.6151
R1049 B.n384 B.n111 10.6151
R1050 B.n701 B.n0 8.11757
R1051 B.n701 B.n1 8.11757
R1052 B.n577 B.n46 6.5566
R1053 B.n565 B.n564 6.5566
R1054 B.n304 B.n303 6.5566
R1055 B.n317 B.n316 6.5566
R1056 B.n46 B.n42 4.05904
R1057 B.n564 B.n563 4.05904
R1058 B.n303 B.n302 4.05904
R1059 B.n318 B.n317 4.05904
R1060 VN.n0 VN.t2 152.019
R1061 VN.n1 VN.t1 152.019
R1062 VN.n0 VN.t0 151.137
R1063 VN.n1 VN.t3 151.137
R1064 VN VN.n1 51.6713
R1065 VN VN.n0 3.55387
R1066 VTAIL.n586 VTAIL.n518 756.745
R1067 VTAIL.n68 VTAIL.n0 756.745
R1068 VTAIL.n142 VTAIL.n74 756.745
R1069 VTAIL.n216 VTAIL.n148 756.745
R1070 VTAIL.n512 VTAIL.n444 756.745
R1071 VTAIL.n438 VTAIL.n370 756.745
R1072 VTAIL.n364 VTAIL.n296 756.745
R1073 VTAIL.n290 VTAIL.n222 756.745
R1074 VTAIL.n543 VTAIL.n542 585
R1075 VTAIL.n545 VTAIL.n544 585
R1076 VTAIL.n538 VTAIL.n537 585
R1077 VTAIL.n551 VTAIL.n550 585
R1078 VTAIL.n553 VTAIL.n552 585
R1079 VTAIL.n534 VTAIL.n533 585
R1080 VTAIL.n560 VTAIL.n559 585
R1081 VTAIL.n561 VTAIL.n532 585
R1082 VTAIL.n563 VTAIL.n562 585
R1083 VTAIL.n530 VTAIL.n529 585
R1084 VTAIL.n569 VTAIL.n568 585
R1085 VTAIL.n571 VTAIL.n570 585
R1086 VTAIL.n526 VTAIL.n525 585
R1087 VTAIL.n577 VTAIL.n576 585
R1088 VTAIL.n579 VTAIL.n578 585
R1089 VTAIL.n522 VTAIL.n521 585
R1090 VTAIL.n585 VTAIL.n584 585
R1091 VTAIL.n587 VTAIL.n586 585
R1092 VTAIL.n25 VTAIL.n24 585
R1093 VTAIL.n27 VTAIL.n26 585
R1094 VTAIL.n20 VTAIL.n19 585
R1095 VTAIL.n33 VTAIL.n32 585
R1096 VTAIL.n35 VTAIL.n34 585
R1097 VTAIL.n16 VTAIL.n15 585
R1098 VTAIL.n42 VTAIL.n41 585
R1099 VTAIL.n43 VTAIL.n14 585
R1100 VTAIL.n45 VTAIL.n44 585
R1101 VTAIL.n12 VTAIL.n11 585
R1102 VTAIL.n51 VTAIL.n50 585
R1103 VTAIL.n53 VTAIL.n52 585
R1104 VTAIL.n8 VTAIL.n7 585
R1105 VTAIL.n59 VTAIL.n58 585
R1106 VTAIL.n61 VTAIL.n60 585
R1107 VTAIL.n4 VTAIL.n3 585
R1108 VTAIL.n67 VTAIL.n66 585
R1109 VTAIL.n69 VTAIL.n68 585
R1110 VTAIL.n99 VTAIL.n98 585
R1111 VTAIL.n101 VTAIL.n100 585
R1112 VTAIL.n94 VTAIL.n93 585
R1113 VTAIL.n107 VTAIL.n106 585
R1114 VTAIL.n109 VTAIL.n108 585
R1115 VTAIL.n90 VTAIL.n89 585
R1116 VTAIL.n116 VTAIL.n115 585
R1117 VTAIL.n117 VTAIL.n88 585
R1118 VTAIL.n119 VTAIL.n118 585
R1119 VTAIL.n86 VTAIL.n85 585
R1120 VTAIL.n125 VTAIL.n124 585
R1121 VTAIL.n127 VTAIL.n126 585
R1122 VTAIL.n82 VTAIL.n81 585
R1123 VTAIL.n133 VTAIL.n132 585
R1124 VTAIL.n135 VTAIL.n134 585
R1125 VTAIL.n78 VTAIL.n77 585
R1126 VTAIL.n141 VTAIL.n140 585
R1127 VTAIL.n143 VTAIL.n142 585
R1128 VTAIL.n173 VTAIL.n172 585
R1129 VTAIL.n175 VTAIL.n174 585
R1130 VTAIL.n168 VTAIL.n167 585
R1131 VTAIL.n181 VTAIL.n180 585
R1132 VTAIL.n183 VTAIL.n182 585
R1133 VTAIL.n164 VTAIL.n163 585
R1134 VTAIL.n190 VTAIL.n189 585
R1135 VTAIL.n191 VTAIL.n162 585
R1136 VTAIL.n193 VTAIL.n192 585
R1137 VTAIL.n160 VTAIL.n159 585
R1138 VTAIL.n199 VTAIL.n198 585
R1139 VTAIL.n201 VTAIL.n200 585
R1140 VTAIL.n156 VTAIL.n155 585
R1141 VTAIL.n207 VTAIL.n206 585
R1142 VTAIL.n209 VTAIL.n208 585
R1143 VTAIL.n152 VTAIL.n151 585
R1144 VTAIL.n215 VTAIL.n214 585
R1145 VTAIL.n217 VTAIL.n216 585
R1146 VTAIL.n513 VTAIL.n512 585
R1147 VTAIL.n511 VTAIL.n510 585
R1148 VTAIL.n448 VTAIL.n447 585
R1149 VTAIL.n505 VTAIL.n504 585
R1150 VTAIL.n503 VTAIL.n502 585
R1151 VTAIL.n452 VTAIL.n451 585
R1152 VTAIL.n497 VTAIL.n496 585
R1153 VTAIL.n495 VTAIL.n494 585
R1154 VTAIL.n456 VTAIL.n455 585
R1155 VTAIL.n460 VTAIL.n458 585
R1156 VTAIL.n489 VTAIL.n488 585
R1157 VTAIL.n487 VTAIL.n486 585
R1158 VTAIL.n462 VTAIL.n461 585
R1159 VTAIL.n481 VTAIL.n480 585
R1160 VTAIL.n479 VTAIL.n478 585
R1161 VTAIL.n466 VTAIL.n465 585
R1162 VTAIL.n473 VTAIL.n472 585
R1163 VTAIL.n471 VTAIL.n470 585
R1164 VTAIL.n439 VTAIL.n438 585
R1165 VTAIL.n437 VTAIL.n436 585
R1166 VTAIL.n374 VTAIL.n373 585
R1167 VTAIL.n431 VTAIL.n430 585
R1168 VTAIL.n429 VTAIL.n428 585
R1169 VTAIL.n378 VTAIL.n377 585
R1170 VTAIL.n423 VTAIL.n422 585
R1171 VTAIL.n421 VTAIL.n420 585
R1172 VTAIL.n382 VTAIL.n381 585
R1173 VTAIL.n386 VTAIL.n384 585
R1174 VTAIL.n415 VTAIL.n414 585
R1175 VTAIL.n413 VTAIL.n412 585
R1176 VTAIL.n388 VTAIL.n387 585
R1177 VTAIL.n407 VTAIL.n406 585
R1178 VTAIL.n405 VTAIL.n404 585
R1179 VTAIL.n392 VTAIL.n391 585
R1180 VTAIL.n399 VTAIL.n398 585
R1181 VTAIL.n397 VTAIL.n396 585
R1182 VTAIL.n365 VTAIL.n364 585
R1183 VTAIL.n363 VTAIL.n362 585
R1184 VTAIL.n300 VTAIL.n299 585
R1185 VTAIL.n357 VTAIL.n356 585
R1186 VTAIL.n355 VTAIL.n354 585
R1187 VTAIL.n304 VTAIL.n303 585
R1188 VTAIL.n349 VTAIL.n348 585
R1189 VTAIL.n347 VTAIL.n346 585
R1190 VTAIL.n308 VTAIL.n307 585
R1191 VTAIL.n312 VTAIL.n310 585
R1192 VTAIL.n341 VTAIL.n340 585
R1193 VTAIL.n339 VTAIL.n338 585
R1194 VTAIL.n314 VTAIL.n313 585
R1195 VTAIL.n333 VTAIL.n332 585
R1196 VTAIL.n331 VTAIL.n330 585
R1197 VTAIL.n318 VTAIL.n317 585
R1198 VTAIL.n325 VTAIL.n324 585
R1199 VTAIL.n323 VTAIL.n322 585
R1200 VTAIL.n291 VTAIL.n290 585
R1201 VTAIL.n289 VTAIL.n288 585
R1202 VTAIL.n226 VTAIL.n225 585
R1203 VTAIL.n283 VTAIL.n282 585
R1204 VTAIL.n281 VTAIL.n280 585
R1205 VTAIL.n230 VTAIL.n229 585
R1206 VTAIL.n275 VTAIL.n274 585
R1207 VTAIL.n273 VTAIL.n272 585
R1208 VTAIL.n234 VTAIL.n233 585
R1209 VTAIL.n238 VTAIL.n236 585
R1210 VTAIL.n267 VTAIL.n266 585
R1211 VTAIL.n265 VTAIL.n264 585
R1212 VTAIL.n240 VTAIL.n239 585
R1213 VTAIL.n259 VTAIL.n258 585
R1214 VTAIL.n257 VTAIL.n256 585
R1215 VTAIL.n244 VTAIL.n243 585
R1216 VTAIL.n251 VTAIL.n250 585
R1217 VTAIL.n249 VTAIL.n248 585
R1218 VTAIL.n541 VTAIL.t5 329.036
R1219 VTAIL.n23 VTAIL.t6 329.036
R1220 VTAIL.n97 VTAIL.t2 329.036
R1221 VTAIL.n171 VTAIL.t0 329.036
R1222 VTAIL.n469 VTAIL.t3 329.036
R1223 VTAIL.n395 VTAIL.t1 329.036
R1224 VTAIL.n321 VTAIL.t4 329.036
R1225 VTAIL.n247 VTAIL.t7 329.036
R1226 VTAIL.n544 VTAIL.n543 171.744
R1227 VTAIL.n544 VTAIL.n537 171.744
R1228 VTAIL.n551 VTAIL.n537 171.744
R1229 VTAIL.n552 VTAIL.n551 171.744
R1230 VTAIL.n552 VTAIL.n533 171.744
R1231 VTAIL.n560 VTAIL.n533 171.744
R1232 VTAIL.n561 VTAIL.n560 171.744
R1233 VTAIL.n562 VTAIL.n561 171.744
R1234 VTAIL.n562 VTAIL.n529 171.744
R1235 VTAIL.n569 VTAIL.n529 171.744
R1236 VTAIL.n570 VTAIL.n569 171.744
R1237 VTAIL.n570 VTAIL.n525 171.744
R1238 VTAIL.n577 VTAIL.n525 171.744
R1239 VTAIL.n578 VTAIL.n577 171.744
R1240 VTAIL.n578 VTAIL.n521 171.744
R1241 VTAIL.n585 VTAIL.n521 171.744
R1242 VTAIL.n586 VTAIL.n585 171.744
R1243 VTAIL.n26 VTAIL.n25 171.744
R1244 VTAIL.n26 VTAIL.n19 171.744
R1245 VTAIL.n33 VTAIL.n19 171.744
R1246 VTAIL.n34 VTAIL.n33 171.744
R1247 VTAIL.n34 VTAIL.n15 171.744
R1248 VTAIL.n42 VTAIL.n15 171.744
R1249 VTAIL.n43 VTAIL.n42 171.744
R1250 VTAIL.n44 VTAIL.n43 171.744
R1251 VTAIL.n44 VTAIL.n11 171.744
R1252 VTAIL.n51 VTAIL.n11 171.744
R1253 VTAIL.n52 VTAIL.n51 171.744
R1254 VTAIL.n52 VTAIL.n7 171.744
R1255 VTAIL.n59 VTAIL.n7 171.744
R1256 VTAIL.n60 VTAIL.n59 171.744
R1257 VTAIL.n60 VTAIL.n3 171.744
R1258 VTAIL.n67 VTAIL.n3 171.744
R1259 VTAIL.n68 VTAIL.n67 171.744
R1260 VTAIL.n100 VTAIL.n99 171.744
R1261 VTAIL.n100 VTAIL.n93 171.744
R1262 VTAIL.n107 VTAIL.n93 171.744
R1263 VTAIL.n108 VTAIL.n107 171.744
R1264 VTAIL.n108 VTAIL.n89 171.744
R1265 VTAIL.n116 VTAIL.n89 171.744
R1266 VTAIL.n117 VTAIL.n116 171.744
R1267 VTAIL.n118 VTAIL.n117 171.744
R1268 VTAIL.n118 VTAIL.n85 171.744
R1269 VTAIL.n125 VTAIL.n85 171.744
R1270 VTAIL.n126 VTAIL.n125 171.744
R1271 VTAIL.n126 VTAIL.n81 171.744
R1272 VTAIL.n133 VTAIL.n81 171.744
R1273 VTAIL.n134 VTAIL.n133 171.744
R1274 VTAIL.n134 VTAIL.n77 171.744
R1275 VTAIL.n141 VTAIL.n77 171.744
R1276 VTAIL.n142 VTAIL.n141 171.744
R1277 VTAIL.n174 VTAIL.n173 171.744
R1278 VTAIL.n174 VTAIL.n167 171.744
R1279 VTAIL.n181 VTAIL.n167 171.744
R1280 VTAIL.n182 VTAIL.n181 171.744
R1281 VTAIL.n182 VTAIL.n163 171.744
R1282 VTAIL.n190 VTAIL.n163 171.744
R1283 VTAIL.n191 VTAIL.n190 171.744
R1284 VTAIL.n192 VTAIL.n191 171.744
R1285 VTAIL.n192 VTAIL.n159 171.744
R1286 VTAIL.n199 VTAIL.n159 171.744
R1287 VTAIL.n200 VTAIL.n199 171.744
R1288 VTAIL.n200 VTAIL.n155 171.744
R1289 VTAIL.n207 VTAIL.n155 171.744
R1290 VTAIL.n208 VTAIL.n207 171.744
R1291 VTAIL.n208 VTAIL.n151 171.744
R1292 VTAIL.n215 VTAIL.n151 171.744
R1293 VTAIL.n216 VTAIL.n215 171.744
R1294 VTAIL.n512 VTAIL.n511 171.744
R1295 VTAIL.n511 VTAIL.n447 171.744
R1296 VTAIL.n504 VTAIL.n447 171.744
R1297 VTAIL.n504 VTAIL.n503 171.744
R1298 VTAIL.n503 VTAIL.n451 171.744
R1299 VTAIL.n496 VTAIL.n451 171.744
R1300 VTAIL.n496 VTAIL.n495 171.744
R1301 VTAIL.n495 VTAIL.n455 171.744
R1302 VTAIL.n460 VTAIL.n455 171.744
R1303 VTAIL.n488 VTAIL.n460 171.744
R1304 VTAIL.n488 VTAIL.n487 171.744
R1305 VTAIL.n487 VTAIL.n461 171.744
R1306 VTAIL.n480 VTAIL.n461 171.744
R1307 VTAIL.n480 VTAIL.n479 171.744
R1308 VTAIL.n479 VTAIL.n465 171.744
R1309 VTAIL.n472 VTAIL.n465 171.744
R1310 VTAIL.n472 VTAIL.n471 171.744
R1311 VTAIL.n438 VTAIL.n437 171.744
R1312 VTAIL.n437 VTAIL.n373 171.744
R1313 VTAIL.n430 VTAIL.n373 171.744
R1314 VTAIL.n430 VTAIL.n429 171.744
R1315 VTAIL.n429 VTAIL.n377 171.744
R1316 VTAIL.n422 VTAIL.n377 171.744
R1317 VTAIL.n422 VTAIL.n421 171.744
R1318 VTAIL.n421 VTAIL.n381 171.744
R1319 VTAIL.n386 VTAIL.n381 171.744
R1320 VTAIL.n414 VTAIL.n386 171.744
R1321 VTAIL.n414 VTAIL.n413 171.744
R1322 VTAIL.n413 VTAIL.n387 171.744
R1323 VTAIL.n406 VTAIL.n387 171.744
R1324 VTAIL.n406 VTAIL.n405 171.744
R1325 VTAIL.n405 VTAIL.n391 171.744
R1326 VTAIL.n398 VTAIL.n391 171.744
R1327 VTAIL.n398 VTAIL.n397 171.744
R1328 VTAIL.n364 VTAIL.n363 171.744
R1329 VTAIL.n363 VTAIL.n299 171.744
R1330 VTAIL.n356 VTAIL.n299 171.744
R1331 VTAIL.n356 VTAIL.n355 171.744
R1332 VTAIL.n355 VTAIL.n303 171.744
R1333 VTAIL.n348 VTAIL.n303 171.744
R1334 VTAIL.n348 VTAIL.n347 171.744
R1335 VTAIL.n347 VTAIL.n307 171.744
R1336 VTAIL.n312 VTAIL.n307 171.744
R1337 VTAIL.n340 VTAIL.n312 171.744
R1338 VTAIL.n340 VTAIL.n339 171.744
R1339 VTAIL.n339 VTAIL.n313 171.744
R1340 VTAIL.n332 VTAIL.n313 171.744
R1341 VTAIL.n332 VTAIL.n331 171.744
R1342 VTAIL.n331 VTAIL.n317 171.744
R1343 VTAIL.n324 VTAIL.n317 171.744
R1344 VTAIL.n324 VTAIL.n323 171.744
R1345 VTAIL.n290 VTAIL.n289 171.744
R1346 VTAIL.n289 VTAIL.n225 171.744
R1347 VTAIL.n282 VTAIL.n225 171.744
R1348 VTAIL.n282 VTAIL.n281 171.744
R1349 VTAIL.n281 VTAIL.n229 171.744
R1350 VTAIL.n274 VTAIL.n229 171.744
R1351 VTAIL.n274 VTAIL.n273 171.744
R1352 VTAIL.n273 VTAIL.n233 171.744
R1353 VTAIL.n238 VTAIL.n233 171.744
R1354 VTAIL.n266 VTAIL.n238 171.744
R1355 VTAIL.n266 VTAIL.n265 171.744
R1356 VTAIL.n265 VTAIL.n239 171.744
R1357 VTAIL.n258 VTAIL.n239 171.744
R1358 VTAIL.n258 VTAIL.n257 171.744
R1359 VTAIL.n257 VTAIL.n243 171.744
R1360 VTAIL.n250 VTAIL.n243 171.744
R1361 VTAIL.n250 VTAIL.n249 171.744
R1362 VTAIL.n543 VTAIL.t5 85.8723
R1363 VTAIL.n25 VTAIL.t6 85.8723
R1364 VTAIL.n99 VTAIL.t2 85.8723
R1365 VTAIL.n173 VTAIL.t0 85.8723
R1366 VTAIL.n471 VTAIL.t3 85.8723
R1367 VTAIL.n397 VTAIL.t1 85.8723
R1368 VTAIL.n323 VTAIL.t4 85.8723
R1369 VTAIL.n249 VTAIL.t7 85.8723
R1370 VTAIL.n591 VTAIL.n590 29.8581
R1371 VTAIL.n73 VTAIL.n72 29.8581
R1372 VTAIL.n147 VTAIL.n146 29.8581
R1373 VTAIL.n221 VTAIL.n220 29.8581
R1374 VTAIL.n517 VTAIL.n516 29.8581
R1375 VTAIL.n443 VTAIL.n442 29.8581
R1376 VTAIL.n369 VTAIL.n368 29.8581
R1377 VTAIL.n295 VTAIL.n294 29.8581
R1378 VTAIL.n591 VTAIL.n517 26.6169
R1379 VTAIL.n295 VTAIL.n221 26.6169
R1380 VTAIL.n563 VTAIL.n530 13.1884
R1381 VTAIL.n45 VTAIL.n12 13.1884
R1382 VTAIL.n119 VTAIL.n86 13.1884
R1383 VTAIL.n193 VTAIL.n160 13.1884
R1384 VTAIL.n458 VTAIL.n456 13.1884
R1385 VTAIL.n384 VTAIL.n382 13.1884
R1386 VTAIL.n310 VTAIL.n308 13.1884
R1387 VTAIL.n236 VTAIL.n234 13.1884
R1388 VTAIL.n564 VTAIL.n532 12.8005
R1389 VTAIL.n568 VTAIL.n567 12.8005
R1390 VTAIL.n46 VTAIL.n14 12.8005
R1391 VTAIL.n50 VTAIL.n49 12.8005
R1392 VTAIL.n120 VTAIL.n88 12.8005
R1393 VTAIL.n124 VTAIL.n123 12.8005
R1394 VTAIL.n194 VTAIL.n162 12.8005
R1395 VTAIL.n198 VTAIL.n197 12.8005
R1396 VTAIL.n494 VTAIL.n493 12.8005
R1397 VTAIL.n490 VTAIL.n489 12.8005
R1398 VTAIL.n420 VTAIL.n419 12.8005
R1399 VTAIL.n416 VTAIL.n415 12.8005
R1400 VTAIL.n346 VTAIL.n345 12.8005
R1401 VTAIL.n342 VTAIL.n341 12.8005
R1402 VTAIL.n272 VTAIL.n271 12.8005
R1403 VTAIL.n268 VTAIL.n267 12.8005
R1404 VTAIL.n559 VTAIL.n558 12.0247
R1405 VTAIL.n571 VTAIL.n528 12.0247
R1406 VTAIL.n41 VTAIL.n40 12.0247
R1407 VTAIL.n53 VTAIL.n10 12.0247
R1408 VTAIL.n115 VTAIL.n114 12.0247
R1409 VTAIL.n127 VTAIL.n84 12.0247
R1410 VTAIL.n189 VTAIL.n188 12.0247
R1411 VTAIL.n201 VTAIL.n158 12.0247
R1412 VTAIL.n497 VTAIL.n454 12.0247
R1413 VTAIL.n486 VTAIL.n459 12.0247
R1414 VTAIL.n423 VTAIL.n380 12.0247
R1415 VTAIL.n412 VTAIL.n385 12.0247
R1416 VTAIL.n349 VTAIL.n306 12.0247
R1417 VTAIL.n338 VTAIL.n311 12.0247
R1418 VTAIL.n275 VTAIL.n232 12.0247
R1419 VTAIL.n264 VTAIL.n237 12.0247
R1420 VTAIL.n557 VTAIL.n534 11.249
R1421 VTAIL.n572 VTAIL.n526 11.249
R1422 VTAIL.n39 VTAIL.n16 11.249
R1423 VTAIL.n54 VTAIL.n8 11.249
R1424 VTAIL.n113 VTAIL.n90 11.249
R1425 VTAIL.n128 VTAIL.n82 11.249
R1426 VTAIL.n187 VTAIL.n164 11.249
R1427 VTAIL.n202 VTAIL.n156 11.249
R1428 VTAIL.n498 VTAIL.n452 11.249
R1429 VTAIL.n485 VTAIL.n462 11.249
R1430 VTAIL.n424 VTAIL.n378 11.249
R1431 VTAIL.n411 VTAIL.n388 11.249
R1432 VTAIL.n350 VTAIL.n304 11.249
R1433 VTAIL.n337 VTAIL.n314 11.249
R1434 VTAIL.n276 VTAIL.n230 11.249
R1435 VTAIL.n263 VTAIL.n240 11.249
R1436 VTAIL.n542 VTAIL.n541 10.7239
R1437 VTAIL.n24 VTAIL.n23 10.7239
R1438 VTAIL.n98 VTAIL.n97 10.7239
R1439 VTAIL.n172 VTAIL.n171 10.7239
R1440 VTAIL.n470 VTAIL.n469 10.7239
R1441 VTAIL.n396 VTAIL.n395 10.7239
R1442 VTAIL.n322 VTAIL.n321 10.7239
R1443 VTAIL.n248 VTAIL.n247 10.7239
R1444 VTAIL.n554 VTAIL.n553 10.4732
R1445 VTAIL.n576 VTAIL.n575 10.4732
R1446 VTAIL.n36 VTAIL.n35 10.4732
R1447 VTAIL.n58 VTAIL.n57 10.4732
R1448 VTAIL.n110 VTAIL.n109 10.4732
R1449 VTAIL.n132 VTAIL.n131 10.4732
R1450 VTAIL.n184 VTAIL.n183 10.4732
R1451 VTAIL.n206 VTAIL.n205 10.4732
R1452 VTAIL.n502 VTAIL.n501 10.4732
R1453 VTAIL.n482 VTAIL.n481 10.4732
R1454 VTAIL.n428 VTAIL.n427 10.4732
R1455 VTAIL.n408 VTAIL.n407 10.4732
R1456 VTAIL.n354 VTAIL.n353 10.4732
R1457 VTAIL.n334 VTAIL.n333 10.4732
R1458 VTAIL.n280 VTAIL.n279 10.4732
R1459 VTAIL.n260 VTAIL.n259 10.4732
R1460 VTAIL.n550 VTAIL.n536 9.69747
R1461 VTAIL.n579 VTAIL.n524 9.69747
R1462 VTAIL.n32 VTAIL.n18 9.69747
R1463 VTAIL.n61 VTAIL.n6 9.69747
R1464 VTAIL.n106 VTAIL.n92 9.69747
R1465 VTAIL.n135 VTAIL.n80 9.69747
R1466 VTAIL.n180 VTAIL.n166 9.69747
R1467 VTAIL.n209 VTAIL.n154 9.69747
R1468 VTAIL.n505 VTAIL.n450 9.69747
R1469 VTAIL.n478 VTAIL.n464 9.69747
R1470 VTAIL.n431 VTAIL.n376 9.69747
R1471 VTAIL.n404 VTAIL.n390 9.69747
R1472 VTAIL.n357 VTAIL.n302 9.69747
R1473 VTAIL.n330 VTAIL.n316 9.69747
R1474 VTAIL.n283 VTAIL.n228 9.69747
R1475 VTAIL.n256 VTAIL.n242 9.69747
R1476 VTAIL.n590 VTAIL.n589 9.45567
R1477 VTAIL.n72 VTAIL.n71 9.45567
R1478 VTAIL.n146 VTAIL.n145 9.45567
R1479 VTAIL.n220 VTAIL.n219 9.45567
R1480 VTAIL.n516 VTAIL.n515 9.45567
R1481 VTAIL.n442 VTAIL.n441 9.45567
R1482 VTAIL.n368 VTAIL.n367 9.45567
R1483 VTAIL.n294 VTAIL.n293 9.45567
R1484 VTAIL.n589 VTAIL.n588 9.3005
R1485 VTAIL.n583 VTAIL.n582 9.3005
R1486 VTAIL.n581 VTAIL.n580 9.3005
R1487 VTAIL.n524 VTAIL.n523 9.3005
R1488 VTAIL.n575 VTAIL.n574 9.3005
R1489 VTAIL.n573 VTAIL.n572 9.3005
R1490 VTAIL.n528 VTAIL.n527 9.3005
R1491 VTAIL.n567 VTAIL.n566 9.3005
R1492 VTAIL.n540 VTAIL.n539 9.3005
R1493 VTAIL.n547 VTAIL.n546 9.3005
R1494 VTAIL.n549 VTAIL.n548 9.3005
R1495 VTAIL.n536 VTAIL.n535 9.3005
R1496 VTAIL.n555 VTAIL.n554 9.3005
R1497 VTAIL.n557 VTAIL.n556 9.3005
R1498 VTAIL.n558 VTAIL.n531 9.3005
R1499 VTAIL.n565 VTAIL.n564 9.3005
R1500 VTAIL.n520 VTAIL.n519 9.3005
R1501 VTAIL.n71 VTAIL.n70 9.3005
R1502 VTAIL.n65 VTAIL.n64 9.3005
R1503 VTAIL.n63 VTAIL.n62 9.3005
R1504 VTAIL.n6 VTAIL.n5 9.3005
R1505 VTAIL.n57 VTAIL.n56 9.3005
R1506 VTAIL.n55 VTAIL.n54 9.3005
R1507 VTAIL.n10 VTAIL.n9 9.3005
R1508 VTAIL.n49 VTAIL.n48 9.3005
R1509 VTAIL.n22 VTAIL.n21 9.3005
R1510 VTAIL.n29 VTAIL.n28 9.3005
R1511 VTAIL.n31 VTAIL.n30 9.3005
R1512 VTAIL.n18 VTAIL.n17 9.3005
R1513 VTAIL.n37 VTAIL.n36 9.3005
R1514 VTAIL.n39 VTAIL.n38 9.3005
R1515 VTAIL.n40 VTAIL.n13 9.3005
R1516 VTAIL.n47 VTAIL.n46 9.3005
R1517 VTAIL.n2 VTAIL.n1 9.3005
R1518 VTAIL.n145 VTAIL.n144 9.3005
R1519 VTAIL.n139 VTAIL.n138 9.3005
R1520 VTAIL.n137 VTAIL.n136 9.3005
R1521 VTAIL.n80 VTAIL.n79 9.3005
R1522 VTAIL.n131 VTAIL.n130 9.3005
R1523 VTAIL.n129 VTAIL.n128 9.3005
R1524 VTAIL.n84 VTAIL.n83 9.3005
R1525 VTAIL.n123 VTAIL.n122 9.3005
R1526 VTAIL.n96 VTAIL.n95 9.3005
R1527 VTAIL.n103 VTAIL.n102 9.3005
R1528 VTAIL.n105 VTAIL.n104 9.3005
R1529 VTAIL.n92 VTAIL.n91 9.3005
R1530 VTAIL.n111 VTAIL.n110 9.3005
R1531 VTAIL.n113 VTAIL.n112 9.3005
R1532 VTAIL.n114 VTAIL.n87 9.3005
R1533 VTAIL.n121 VTAIL.n120 9.3005
R1534 VTAIL.n76 VTAIL.n75 9.3005
R1535 VTAIL.n219 VTAIL.n218 9.3005
R1536 VTAIL.n213 VTAIL.n212 9.3005
R1537 VTAIL.n211 VTAIL.n210 9.3005
R1538 VTAIL.n154 VTAIL.n153 9.3005
R1539 VTAIL.n205 VTAIL.n204 9.3005
R1540 VTAIL.n203 VTAIL.n202 9.3005
R1541 VTAIL.n158 VTAIL.n157 9.3005
R1542 VTAIL.n197 VTAIL.n196 9.3005
R1543 VTAIL.n170 VTAIL.n169 9.3005
R1544 VTAIL.n177 VTAIL.n176 9.3005
R1545 VTAIL.n179 VTAIL.n178 9.3005
R1546 VTAIL.n166 VTAIL.n165 9.3005
R1547 VTAIL.n185 VTAIL.n184 9.3005
R1548 VTAIL.n187 VTAIL.n186 9.3005
R1549 VTAIL.n188 VTAIL.n161 9.3005
R1550 VTAIL.n195 VTAIL.n194 9.3005
R1551 VTAIL.n150 VTAIL.n149 9.3005
R1552 VTAIL.n468 VTAIL.n467 9.3005
R1553 VTAIL.n475 VTAIL.n474 9.3005
R1554 VTAIL.n477 VTAIL.n476 9.3005
R1555 VTAIL.n464 VTAIL.n463 9.3005
R1556 VTAIL.n483 VTAIL.n482 9.3005
R1557 VTAIL.n485 VTAIL.n484 9.3005
R1558 VTAIL.n459 VTAIL.n457 9.3005
R1559 VTAIL.n491 VTAIL.n490 9.3005
R1560 VTAIL.n515 VTAIL.n514 9.3005
R1561 VTAIL.n446 VTAIL.n445 9.3005
R1562 VTAIL.n509 VTAIL.n508 9.3005
R1563 VTAIL.n507 VTAIL.n506 9.3005
R1564 VTAIL.n450 VTAIL.n449 9.3005
R1565 VTAIL.n501 VTAIL.n500 9.3005
R1566 VTAIL.n499 VTAIL.n498 9.3005
R1567 VTAIL.n454 VTAIL.n453 9.3005
R1568 VTAIL.n493 VTAIL.n492 9.3005
R1569 VTAIL.n394 VTAIL.n393 9.3005
R1570 VTAIL.n401 VTAIL.n400 9.3005
R1571 VTAIL.n403 VTAIL.n402 9.3005
R1572 VTAIL.n390 VTAIL.n389 9.3005
R1573 VTAIL.n409 VTAIL.n408 9.3005
R1574 VTAIL.n411 VTAIL.n410 9.3005
R1575 VTAIL.n385 VTAIL.n383 9.3005
R1576 VTAIL.n417 VTAIL.n416 9.3005
R1577 VTAIL.n441 VTAIL.n440 9.3005
R1578 VTAIL.n372 VTAIL.n371 9.3005
R1579 VTAIL.n435 VTAIL.n434 9.3005
R1580 VTAIL.n433 VTAIL.n432 9.3005
R1581 VTAIL.n376 VTAIL.n375 9.3005
R1582 VTAIL.n427 VTAIL.n426 9.3005
R1583 VTAIL.n425 VTAIL.n424 9.3005
R1584 VTAIL.n380 VTAIL.n379 9.3005
R1585 VTAIL.n419 VTAIL.n418 9.3005
R1586 VTAIL.n320 VTAIL.n319 9.3005
R1587 VTAIL.n327 VTAIL.n326 9.3005
R1588 VTAIL.n329 VTAIL.n328 9.3005
R1589 VTAIL.n316 VTAIL.n315 9.3005
R1590 VTAIL.n335 VTAIL.n334 9.3005
R1591 VTAIL.n337 VTAIL.n336 9.3005
R1592 VTAIL.n311 VTAIL.n309 9.3005
R1593 VTAIL.n343 VTAIL.n342 9.3005
R1594 VTAIL.n367 VTAIL.n366 9.3005
R1595 VTAIL.n298 VTAIL.n297 9.3005
R1596 VTAIL.n361 VTAIL.n360 9.3005
R1597 VTAIL.n359 VTAIL.n358 9.3005
R1598 VTAIL.n302 VTAIL.n301 9.3005
R1599 VTAIL.n353 VTAIL.n352 9.3005
R1600 VTAIL.n351 VTAIL.n350 9.3005
R1601 VTAIL.n306 VTAIL.n305 9.3005
R1602 VTAIL.n345 VTAIL.n344 9.3005
R1603 VTAIL.n246 VTAIL.n245 9.3005
R1604 VTAIL.n253 VTAIL.n252 9.3005
R1605 VTAIL.n255 VTAIL.n254 9.3005
R1606 VTAIL.n242 VTAIL.n241 9.3005
R1607 VTAIL.n261 VTAIL.n260 9.3005
R1608 VTAIL.n263 VTAIL.n262 9.3005
R1609 VTAIL.n237 VTAIL.n235 9.3005
R1610 VTAIL.n269 VTAIL.n268 9.3005
R1611 VTAIL.n293 VTAIL.n292 9.3005
R1612 VTAIL.n224 VTAIL.n223 9.3005
R1613 VTAIL.n287 VTAIL.n286 9.3005
R1614 VTAIL.n285 VTAIL.n284 9.3005
R1615 VTAIL.n228 VTAIL.n227 9.3005
R1616 VTAIL.n279 VTAIL.n278 9.3005
R1617 VTAIL.n277 VTAIL.n276 9.3005
R1618 VTAIL.n232 VTAIL.n231 9.3005
R1619 VTAIL.n271 VTAIL.n270 9.3005
R1620 VTAIL.n549 VTAIL.n538 8.92171
R1621 VTAIL.n580 VTAIL.n522 8.92171
R1622 VTAIL.n31 VTAIL.n20 8.92171
R1623 VTAIL.n62 VTAIL.n4 8.92171
R1624 VTAIL.n105 VTAIL.n94 8.92171
R1625 VTAIL.n136 VTAIL.n78 8.92171
R1626 VTAIL.n179 VTAIL.n168 8.92171
R1627 VTAIL.n210 VTAIL.n152 8.92171
R1628 VTAIL.n506 VTAIL.n448 8.92171
R1629 VTAIL.n477 VTAIL.n466 8.92171
R1630 VTAIL.n432 VTAIL.n374 8.92171
R1631 VTAIL.n403 VTAIL.n392 8.92171
R1632 VTAIL.n358 VTAIL.n300 8.92171
R1633 VTAIL.n329 VTAIL.n318 8.92171
R1634 VTAIL.n284 VTAIL.n226 8.92171
R1635 VTAIL.n255 VTAIL.n244 8.92171
R1636 VTAIL.n546 VTAIL.n545 8.14595
R1637 VTAIL.n584 VTAIL.n583 8.14595
R1638 VTAIL.n28 VTAIL.n27 8.14595
R1639 VTAIL.n66 VTAIL.n65 8.14595
R1640 VTAIL.n102 VTAIL.n101 8.14595
R1641 VTAIL.n140 VTAIL.n139 8.14595
R1642 VTAIL.n176 VTAIL.n175 8.14595
R1643 VTAIL.n214 VTAIL.n213 8.14595
R1644 VTAIL.n510 VTAIL.n509 8.14595
R1645 VTAIL.n474 VTAIL.n473 8.14595
R1646 VTAIL.n436 VTAIL.n435 8.14595
R1647 VTAIL.n400 VTAIL.n399 8.14595
R1648 VTAIL.n362 VTAIL.n361 8.14595
R1649 VTAIL.n326 VTAIL.n325 8.14595
R1650 VTAIL.n288 VTAIL.n287 8.14595
R1651 VTAIL.n252 VTAIL.n251 8.14595
R1652 VTAIL.n542 VTAIL.n540 7.3702
R1653 VTAIL.n587 VTAIL.n520 7.3702
R1654 VTAIL.n590 VTAIL.n518 7.3702
R1655 VTAIL.n24 VTAIL.n22 7.3702
R1656 VTAIL.n69 VTAIL.n2 7.3702
R1657 VTAIL.n72 VTAIL.n0 7.3702
R1658 VTAIL.n98 VTAIL.n96 7.3702
R1659 VTAIL.n143 VTAIL.n76 7.3702
R1660 VTAIL.n146 VTAIL.n74 7.3702
R1661 VTAIL.n172 VTAIL.n170 7.3702
R1662 VTAIL.n217 VTAIL.n150 7.3702
R1663 VTAIL.n220 VTAIL.n148 7.3702
R1664 VTAIL.n516 VTAIL.n444 7.3702
R1665 VTAIL.n513 VTAIL.n446 7.3702
R1666 VTAIL.n470 VTAIL.n468 7.3702
R1667 VTAIL.n442 VTAIL.n370 7.3702
R1668 VTAIL.n439 VTAIL.n372 7.3702
R1669 VTAIL.n396 VTAIL.n394 7.3702
R1670 VTAIL.n368 VTAIL.n296 7.3702
R1671 VTAIL.n365 VTAIL.n298 7.3702
R1672 VTAIL.n322 VTAIL.n320 7.3702
R1673 VTAIL.n294 VTAIL.n222 7.3702
R1674 VTAIL.n291 VTAIL.n224 7.3702
R1675 VTAIL.n248 VTAIL.n246 7.3702
R1676 VTAIL.n588 VTAIL.n587 6.59444
R1677 VTAIL.n588 VTAIL.n518 6.59444
R1678 VTAIL.n70 VTAIL.n69 6.59444
R1679 VTAIL.n70 VTAIL.n0 6.59444
R1680 VTAIL.n144 VTAIL.n143 6.59444
R1681 VTAIL.n144 VTAIL.n74 6.59444
R1682 VTAIL.n218 VTAIL.n217 6.59444
R1683 VTAIL.n218 VTAIL.n148 6.59444
R1684 VTAIL.n514 VTAIL.n444 6.59444
R1685 VTAIL.n514 VTAIL.n513 6.59444
R1686 VTAIL.n440 VTAIL.n370 6.59444
R1687 VTAIL.n440 VTAIL.n439 6.59444
R1688 VTAIL.n366 VTAIL.n296 6.59444
R1689 VTAIL.n366 VTAIL.n365 6.59444
R1690 VTAIL.n292 VTAIL.n222 6.59444
R1691 VTAIL.n292 VTAIL.n291 6.59444
R1692 VTAIL.n545 VTAIL.n540 5.81868
R1693 VTAIL.n584 VTAIL.n520 5.81868
R1694 VTAIL.n27 VTAIL.n22 5.81868
R1695 VTAIL.n66 VTAIL.n2 5.81868
R1696 VTAIL.n101 VTAIL.n96 5.81868
R1697 VTAIL.n140 VTAIL.n76 5.81868
R1698 VTAIL.n175 VTAIL.n170 5.81868
R1699 VTAIL.n214 VTAIL.n150 5.81868
R1700 VTAIL.n510 VTAIL.n446 5.81868
R1701 VTAIL.n473 VTAIL.n468 5.81868
R1702 VTAIL.n436 VTAIL.n372 5.81868
R1703 VTAIL.n399 VTAIL.n394 5.81868
R1704 VTAIL.n362 VTAIL.n298 5.81868
R1705 VTAIL.n325 VTAIL.n320 5.81868
R1706 VTAIL.n288 VTAIL.n224 5.81868
R1707 VTAIL.n251 VTAIL.n246 5.81868
R1708 VTAIL.n546 VTAIL.n538 5.04292
R1709 VTAIL.n583 VTAIL.n522 5.04292
R1710 VTAIL.n28 VTAIL.n20 5.04292
R1711 VTAIL.n65 VTAIL.n4 5.04292
R1712 VTAIL.n102 VTAIL.n94 5.04292
R1713 VTAIL.n139 VTAIL.n78 5.04292
R1714 VTAIL.n176 VTAIL.n168 5.04292
R1715 VTAIL.n213 VTAIL.n152 5.04292
R1716 VTAIL.n509 VTAIL.n448 5.04292
R1717 VTAIL.n474 VTAIL.n466 5.04292
R1718 VTAIL.n435 VTAIL.n374 5.04292
R1719 VTAIL.n400 VTAIL.n392 5.04292
R1720 VTAIL.n361 VTAIL.n300 5.04292
R1721 VTAIL.n326 VTAIL.n318 5.04292
R1722 VTAIL.n287 VTAIL.n226 5.04292
R1723 VTAIL.n252 VTAIL.n244 5.04292
R1724 VTAIL.n550 VTAIL.n549 4.26717
R1725 VTAIL.n580 VTAIL.n579 4.26717
R1726 VTAIL.n32 VTAIL.n31 4.26717
R1727 VTAIL.n62 VTAIL.n61 4.26717
R1728 VTAIL.n106 VTAIL.n105 4.26717
R1729 VTAIL.n136 VTAIL.n135 4.26717
R1730 VTAIL.n180 VTAIL.n179 4.26717
R1731 VTAIL.n210 VTAIL.n209 4.26717
R1732 VTAIL.n506 VTAIL.n505 4.26717
R1733 VTAIL.n478 VTAIL.n477 4.26717
R1734 VTAIL.n432 VTAIL.n431 4.26717
R1735 VTAIL.n404 VTAIL.n403 4.26717
R1736 VTAIL.n358 VTAIL.n357 4.26717
R1737 VTAIL.n330 VTAIL.n329 4.26717
R1738 VTAIL.n284 VTAIL.n283 4.26717
R1739 VTAIL.n256 VTAIL.n255 4.26717
R1740 VTAIL.n553 VTAIL.n536 3.49141
R1741 VTAIL.n576 VTAIL.n524 3.49141
R1742 VTAIL.n35 VTAIL.n18 3.49141
R1743 VTAIL.n58 VTAIL.n6 3.49141
R1744 VTAIL.n109 VTAIL.n92 3.49141
R1745 VTAIL.n132 VTAIL.n80 3.49141
R1746 VTAIL.n183 VTAIL.n166 3.49141
R1747 VTAIL.n206 VTAIL.n154 3.49141
R1748 VTAIL.n502 VTAIL.n450 3.49141
R1749 VTAIL.n481 VTAIL.n464 3.49141
R1750 VTAIL.n428 VTAIL.n376 3.49141
R1751 VTAIL.n407 VTAIL.n390 3.49141
R1752 VTAIL.n354 VTAIL.n302 3.49141
R1753 VTAIL.n333 VTAIL.n316 3.49141
R1754 VTAIL.n280 VTAIL.n228 3.49141
R1755 VTAIL.n259 VTAIL.n242 3.49141
R1756 VTAIL.n554 VTAIL.n534 2.71565
R1757 VTAIL.n575 VTAIL.n526 2.71565
R1758 VTAIL.n36 VTAIL.n16 2.71565
R1759 VTAIL.n57 VTAIL.n8 2.71565
R1760 VTAIL.n110 VTAIL.n90 2.71565
R1761 VTAIL.n131 VTAIL.n82 2.71565
R1762 VTAIL.n184 VTAIL.n164 2.71565
R1763 VTAIL.n205 VTAIL.n156 2.71565
R1764 VTAIL.n501 VTAIL.n452 2.71565
R1765 VTAIL.n482 VTAIL.n462 2.71565
R1766 VTAIL.n427 VTAIL.n378 2.71565
R1767 VTAIL.n408 VTAIL.n388 2.71565
R1768 VTAIL.n353 VTAIL.n304 2.71565
R1769 VTAIL.n334 VTAIL.n314 2.71565
R1770 VTAIL.n279 VTAIL.n230 2.71565
R1771 VTAIL.n260 VTAIL.n240 2.71565
R1772 VTAIL.n369 VTAIL.n295 2.66429
R1773 VTAIL.n517 VTAIL.n443 2.66429
R1774 VTAIL.n221 VTAIL.n147 2.66429
R1775 VTAIL.n541 VTAIL.n539 2.41282
R1776 VTAIL.n23 VTAIL.n21 2.41282
R1777 VTAIL.n97 VTAIL.n95 2.41282
R1778 VTAIL.n171 VTAIL.n169 2.41282
R1779 VTAIL.n469 VTAIL.n467 2.41282
R1780 VTAIL.n395 VTAIL.n393 2.41282
R1781 VTAIL.n321 VTAIL.n319 2.41282
R1782 VTAIL.n247 VTAIL.n245 2.41282
R1783 VTAIL.n559 VTAIL.n557 1.93989
R1784 VTAIL.n572 VTAIL.n571 1.93989
R1785 VTAIL.n41 VTAIL.n39 1.93989
R1786 VTAIL.n54 VTAIL.n53 1.93989
R1787 VTAIL.n115 VTAIL.n113 1.93989
R1788 VTAIL.n128 VTAIL.n127 1.93989
R1789 VTAIL.n189 VTAIL.n187 1.93989
R1790 VTAIL.n202 VTAIL.n201 1.93989
R1791 VTAIL.n498 VTAIL.n497 1.93989
R1792 VTAIL.n486 VTAIL.n485 1.93989
R1793 VTAIL.n424 VTAIL.n423 1.93989
R1794 VTAIL.n412 VTAIL.n411 1.93989
R1795 VTAIL.n350 VTAIL.n349 1.93989
R1796 VTAIL.n338 VTAIL.n337 1.93989
R1797 VTAIL.n276 VTAIL.n275 1.93989
R1798 VTAIL.n264 VTAIL.n263 1.93989
R1799 VTAIL VTAIL.n73 1.39059
R1800 VTAIL VTAIL.n591 1.27421
R1801 VTAIL.n558 VTAIL.n532 1.16414
R1802 VTAIL.n568 VTAIL.n528 1.16414
R1803 VTAIL.n40 VTAIL.n14 1.16414
R1804 VTAIL.n50 VTAIL.n10 1.16414
R1805 VTAIL.n114 VTAIL.n88 1.16414
R1806 VTAIL.n124 VTAIL.n84 1.16414
R1807 VTAIL.n188 VTAIL.n162 1.16414
R1808 VTAIL.n198 VTAIL.n158 1.16414
R1809 VTAIL.n494 VTAIL.n454 1.16414
R1810 VTAIL.n489 VTAIL.n459 1.16414
R1811 VTAIL.n420 VTAIL.n380 1.16414
R1812 VTAIL.n415 VTAIL.n385 1.16414
R1813 VTAIL.n346 VTAIL.n306 1.16414
R1814 VTAIL.n341 VTAIL.n311 1.16414
R1815 VTAIL.n272 VTAIL.n232 1.16414
R1816 VTAIL.n267 VTAIL.n237 1.16414
R1817 VTAIL.n443 VTAIL.n369 0.470328
R1818 VTAIL.n147 VTAIL.n73 0.470328
R1819 VTAIL.n564 VTAIL.n563 0.388379
R1820 VTAIL.n567 VTAIL.n530 0.388379
R1821 VTAIL.n46 VTAIL.n45 0.388379
R1822 VTAIL.n49 VTAIL.n12 0.388379
R1823 VTAIL.n120 VTAIL.n119 0.388379
R1824 VTAIL.n123 VTAIL.n86 0.388379
R1825 VTAIL.n194 VTAIL.n193 0.388379
R1826 VTAIL.n197 VTAIL.n160 0.388379
R1827 VTAIL.n493 VTAIL.n456 0.388379
R1828 VTAIL.n490 VTAIL.n458 0.388379
R1829 VTAIL.n419 VTAIL.n382 0.388379
R1830 VTAIL.n416 VTAIL.n384 0.388379
R1831 VTAIL.n345 VTAIL.n308 0.388379
R1832 VTAIL.n342 VTAIL.n310 0.388379
R1833 VTAIL.n271 VTAIL.n234 0.388379
R1834 VTAIL.n268 VTAIL.n236 0.388379
R1835 VTAIL.n547 VTAIL.n539 0.155672
R1836 VTAIL.n548 VTAIL.n547 0.155672
R1837 VTAIL.n548 VTAIL.n535 0.155672
R1838 VTAIL.n555 VTAIL.n535 0.155672
R1839 VTAIL.n556 VTAIL.n555 0.155672
R1840 VTAIL.n556 VTAIL.n531 0.155672
R1841 VTAIL.n565 VTAIL.n531 0.155672
R1842 VTAIL.n566 VTAIL.n565 0.155672
R1843 VTAIL.n566 VTAIL.n527 0.155672
R1844 VTAIL.n573 VTAIL.n527 0.155672
R1845 VTAIL.n574 VTAIL.n573 0.155672
R1846 VTAIL.n574 VTAIL.n523 0.155672
R1847 VTAIL.n581 VTAIL.n523 0.155672
R1848 VTAIL.n582 VTAIL.n581 0.155672
R1849 VTAIL.n582 VTAIL.n519 0.155672
R1850 VTAIL.n589 VTAIL.n519 0.155672
R1851 VTAIL.n29 VTAIL.n21 0.155672
R1852 VTAIL.n30 VTAIL.n29 0.155672
R1853 VTAIL.n30 VTAIL.n17 0.155672
R1854 VTAIL.n37 VTAIL.n17 0.155672
R1855 VTAIL.n38 VTAIL.n37 0.155672
R1856 VTAIL.n38 VTAIL.n13 0.155672
R1857 VTAIL.n47 VTAIL.n13 0.155672
R1858 VTAIL.n48 VTAIL.n47 0.155672
R1859 VTAIL.n48 VTAIL.n9 0.155672
R1860 VTAIL.n55 VTAIL.n9 0.155672
R1861 VTAIL.n56 VTAIL.n55 0.155672
R1862 VTAIL.n56 VTAIL.n5 0.155672
R1863 VTAIL.n63 VTAIL.n5 0.155672
R1864 VTAIL.n64 VTAIL.n63 0.155672
R1865 VTAIL.n64 VTAIL.n1 0.155672
R1866 VTAIL.n71 VTAIL.n1 0.155672
R1867 VTAIL.n103 VTAIL.n95 0.155672
R1868 VTAIL.n104 VTAIL.n103 0.155672
R1869 VTAIL.n104 VTAIL.n91 0.155672
R1870 VTAIL.n111 VTAIL.n91 0.155672
R1871 VTAIL.n112 VTAIL.n111 0.155672
R1872 VTAIL.n112 VTAIL.n87 0.155672
R1873 VTAIL.n121 VTAIL.n87 0.155672
R1874 VTAIL.n122 VTAIL.n121 0.155672
R1875 VTAIL.n122 VTAIL.n83 0.155672
R1876 VTAIL.n129 VTAIL.n83 0.155672
R1877 VTAIL.n130 VTAIL.n129 0.155672
R1878 VTAIL.n130 VTAIL.n79 0.155672
R1879 VTAIL.n137 VTAIL.n79 0.155672
R1880 VTAIL.n138 VTAIL.n137 0.155672
R1881 VTAIL.n138 VTAIL.n75 0.155672
R1882 VTAIL.n145 VTAIL.n75 0.155672
R1883 VTAIL.n177 VTAIL.n169 0.155672
R1884 VTAIL.n178 VTAIL.n177 0.155672
R1885 VTAIL.n178 VTAIL.n165 0.155672
R1886 VTAIL.n185 VTAIL.n165 0.155672
R1887 VTAIL.n186 VTAIL.n185 0.155672
R1888 VTAIL.n186 VTAIL.n161 0.155672
R1889 VTAIL.n195 VTAIL.n161 0.155672
R1890 VTAIL.n196 VTAIL.n195 0.155672
R1891 VTAIL.n196 VTAIL.n157 0.155672
R1892 VTAIL.n203 VTAIL.n157 0.155672
R1893 VTAIL.n204 VTAIL.n203 0.155672
R1894 VTAIL.n204 VTAIL.n153 0.155672
R1895 VTAIL.n211 VTAIL.n153 0.155672
R1896 VTAIL.n212 VTAIL.n211 0.155672
R1897 VTAIL.n212 VTAIL.n149 0.155672
R1898 VTAIL.n219 VTAIL.n149 0.155672
R1899 VTAIL.n515 VTAIL.n445 0.155672
R1900 VTAIL.n508 VTAIL.n445 0.155672
R1901 VTAIL.n508 VTAIL.n507 0.155672
R1902 VTAIL.n507 VTAIL.n449 0.155672
R1903 VTAIL.n500 VTAIL.n449 0.155672
R1904 VTAIL.n500 VTAIL.n499 0.155672
R1905 VTAIL.n499 VTAIL.n453 0.155672
R1906 VTAIL.n492 VTAIL.n453 0.155672
R1907 VTAIL.n492 VTAIL.n491 0.155672
R1908 VTAIL.n491 VTAIL.n457 0.155672
R1909 VTAIL.n484 VTAIL.n457 0.155672
R1910 VTAIL.n484 VTAIL.n483 0.155672
R1911 VTAIL.n483 VTAIL.n463 0.155672
R1912 VTAIL.n476 VTAIL.n463 0.155672
R1913 VTAIL.n476 VTAIL.n475 0.155672
R1914 VTAIL.n475 VTAIL.n467 0.155672
R1915 VTAIL.n441 VTAIL.n371 0.155672
R1916 VTAIL.n434 VTAIL.n371 0.155672
R1917 VTAIL.n434 VTAIL.n433 0.155672
R1918 VTAIL.n433 VTAIL.n375 0.155672
R1919 VTAIL.n426 VTAIL.n375 0.155672
R1920 VTAIL.n426 VTAIL.n425 0.155672
R1921 VTAIL.n425 VTAIL.n379 0.155672
R1922 VTAIL.n418 VTAIL.n379 0.155672
R1923 VTAIL.n418 VTAIL.n417 0.155672
R1924 VTAIL.n417 VTAIL.n383 0.155672
R1925 VTAIL.n410 VTAIL.n383 0.155672
R1926 VTAIL.n410 VTAIL.n409 0.155672
R1927 VTAIL.n409 VTAIL.n389 0.155672
R1928 VTAIL.n402 VTAIL.n389 0.155672
R1929 VTAIL.n402 VTAIL.n401 0.155672
R1930 VTAIL.n401 VTAIL.n393 0.155672
R1931 VTAIL.n367 VTAIL.n297 0.155672
R1932 VTAIL.n360 VTAIL.n297 0.155672
R1933 VTAIL.n360 VTAIL.n359 0.155672
R1934 VTAIL.n359 VTAIL.n301 0.155672
R1935 VTAIL.n352 VTAIL.n301 0.155672
R1936 VTAIL.n352 VTAIL.n351 0.155672
R1937 VTAIL.n351 VTAIL.n305 0.155672
R1938 VTAIL.n344 VTAIL.n305 0.155672
R1939 VTAIL.n344 VTAIL.n343 0.155672
R1940 VTAIL.n343 VTAIL.n309 0.155672
R1941 VTAIL.n336 VTAIL.n309 0.155672
R1942 VTAIL.n336 VTAIL.n335 0.155672
R1943 VTAIL.n335 VTAIL.n315 0.155672
R1944 VTAIL.n328 VTAIL.n315 0.155672
R1945 VTAIL.n328 VTAIL.n327 0.155672
R1946 VTAIL.n327 VTAIL.n319 0.155672
R1947 VTAIL.n293 VTAIL.n223 0.155672
R1948 VTAIL.n286 VTAIL.n223 0.155672
R1949 VTAIL.n286 VTAIL.n285 0.155672
R1950 VTAIL.n285 VTAIL.n227 0.155672
R1951 VTAIL.n278 VTAIL.n227 0.155672
R1952 VTAIL.n278 VTAIL.n277 0.155672
R1953 VTAIL.n277 VTAIL.n231 0.155672
R1954 VTAIL.n270 VTAIL.n231 0.155672
R1955 VTAIL.n270 VTAIL.n269 0.155672
R1956 VTAIL.n269 VTAIL.n235 0.155672
R1957 VTAIL.n262 VTAIL.n235 0.155672
R1958 VTAIL.n262 VTAIL.n261 0.155672
R1959 VTAIL.n261 VTAIL.n241 0.155672
R1960 VTAIL.n254 VTAIL.n241 0.155672
R1961 VTAIL.n254 VTAIL.n253 0.155672
R1962 VTAIL.n253 VTAIL.n245 0.155672
R1963 VDD2.n2 VDD2.n0 113.246
R1964 VDD2.n2 VDD2.n1 69.9534
R1965 VDD2.n1 VDD2.t0 2.41903
R1966 VDD2.n1 VDD2.t2 2.41903
R1967 VDD2.n0 VDD2.t1 2.41903
R1968 VDD2.n0 VDD2.t3 2.41903
R1969 VDD2 VDD2.n2 0.0586897
R1970 VP.n16 VP.n0 161.3
R1971 VP.n15 VP.n14 161.3
R1972 VP.n13 VP.n1 161.3
R1973 VP.n12 VP.n11 161.3
R1974 VP.n10 VP.n2 161.3
R1975 VP.n9 VP.n8 161.3
R1976 VP.n7 VP.n3 161.3
R1977 VP.n4 VP.t2 152.019
R1978 VP.n4 VP.t0 151.137
R1979 VP.n5 VP.t3 117.358
R1980 VP.n17 VP.t1 117.358
R1981 VP.n6 VP.n5 108.695
R1982 VP.n18 VP.n17 108.695
R1983 VP.n6 VP.n4 51.3925
R1984 VP.n11 VP.n10 40.577
R1985 VP.n11 VP.n1 40.577
R1986 VP.n9 VP.n3 24.5923
R1987 VP.n10 VP.n9 24.5923
R1988 VP.n15 VP.n1 24.5923
R1989 VP.n16 VP.n15 24.5923
R1990 VP.n5 VP.n3 2.21377
R1991 VP.n17 VP.n16 2.21377
R1992 VP.n7 VP.n6 0.278335
R1993 VP.n18 VP.n0 0.278335
R1994 VP.n8 VP.n7 0.189894
R1995 VP.n8 VP.n2 0.189894
R1996 VP.n12 VP.n2 0.189894
R1997 VP.n13 VP.n12 0.189894
R1998 VP.n14 VP.n13 0.189894
R1999 VP.n14 VP.n0 0.189894
R2000 VP VP.n18 0.153485
R2001 VDD1 VDD1.n1 113.77
R2002 VDD1 VDD1.n0 70.0116
R2003 VDD1.n0 VDD1.t1 2.41903
R2004 VDD1.n0 VDD1.t3 2.41903
R2005 VDD1.n1 VDD1.t0 2.41903
R2006 VDD1.n1 VDD1.t2 2.41903
C0 w_n2824_n3656# VDD1 1.51975f
C1 VDD1 VP 5.5971f
C2 B VDD2 1.38286f
C3 VDD2 VN 5.34254f
C4 VDD2 VTAIL 5.82597f
C5 w_n2824_n3656# VDD2 1.57941f
C6 B VN 1.15988f
C7 B VTAIL 5.49432f
C8 VTAIL VN 5.20556f
C9 VDD2 VP 0.404658f
C10 B w_n2824_n3656# 9.84665f
C11 w_n2824_n3656# VN 4.83919f
C12 w_n2824_n3656# VTAIL 4.30071f
C13 B VP 1.76374f
C14 VN VP 6.57016f
C15 VTAIL VP 5.21966f
C16 w_n2824_n3656# VP 5.20263f
C17 VDD2 VDD1 1.05943f
C18 B VDD1 1.32806f
C19 VDD1 VN 0.149316f
C20 VDD1 VTAIL 5.77069f
C21 VDD2 VSUBS 1.009813f
C22 VDD1 VSUBS 6.03504f
C23 VTAIL VSUBS 1.300026f
C24 VN VSUBS 5.5642f
C25 VP VSUBS 2.412526f
C26 B VSUBS 4.53622f
C27 w_n2824_n3656# VSUBS 0.126843p
C28 VDD1.t1 VSUBS 0.28785f
C29 VDD1.t3 VSUBS 0.28785f
C30 VDD1.n0 VSUBS 2.27781f
C31 VDD1.t0 VSUBS 0.28785f
C32 VDD1.t2 VSUBS 0.28785f
C33 VDD1.n1 VSUBS 3.10894f
C34 VP.n0 VSUBS 0.042049f
C35 VP.t1 VSUBS 3.23351f
C36 VP.n1 VSUBS 0.063059f
C37 VP.n2 VSUBS 0.031896f
C38 VP.n3 VSUBS 0.032576f
C39 VP.t0 VSUBS 3.53384f
C40 VP.t2 VSUBS 3.54149f
C41 VP.n4 VSUBS 4.0815f
C42 VP.t3 VSUBS 3.23351f
C43 VP.n5 VSUBS 1.23417f
C44 VP.n6 VSUBS 1.83201f
C45 VP.n7 VSUBS 0.042049f
C46 VP.n8 VSUBS 0.031896f
C47 VP.n9 VSUBS 0.059148f
C48 VP.n10 VSUBS 0.063059f
C49 VP.n11 VSUBS 0.025761f
C50 VP.n12 VSUBS 0.031896f
C51 VP.n13 VSUBS 0.031896f
C52 VP.n14 VSUBS 0.031896f
C53 VP.n15 VSUBS 0.059148f
C54 VP.n16 VSUBS 0.032576f
C55 VP.n17 VSUBS 1.23417f
C56 VP.n18 VSUBS 0.059379f
C57 VDD2.t1 VSUBS 0.282758f
C58 VDD2.t3 VSUBS 0.282758f
C59 VDD2.n0 VSUBS 3.02773f
C60 VDD2.t0 VSUBS 0.282758f
C61 VDD2.t2 VSUBS 0.282758f
C62 VDD2.n1 VSUBS 2.23688f
C63 VDD2.n2 VSUBS 4.470109f
C64 VTAIL.n0 VSUBS 0.025154f
C65 VTAIL.n1 VSUBS 0.023341f
C66 VTAIL.n2 VSUBS 0.012543f
C67 VTAIL.n3 VSUBS 0.029646f
C68 VTAIL.n4 VSUBS 0.01328f
C69 VTAIL.n5 VSUBS 0.023341f
C70 VTAIL.n6 VSUBS 0.012543f
C71 VTAIL.n7 VSUBS 0.029646f
C72 VTAIL.n8 VSUBS 0.01328f
C73 VTAIL.n9 VSUBS 0.023341f
C74 VTAIL.n10 VSUBS 0.012543f
C75 VTAIL.n11 VSUBS 0.029646f
C76 VTAIL.n12 VSUBS 0.012912f
C77 VTAIL.n13 VSUBS 0.023341f
C78 VTAIL.n14 VSUBS 0.01328f
C79 VTAIL.n15 VSUBS 0.029646f
C80 VTAIL.n16 VSUBS 0.01328f
C81 VTAIL.n17 VSUBS 0.023341f
C82 VTAIL.n18 VSUBS 0.012543f
C83 VTAIL.n19 VSUBS 0.029646f
C84 VTAIL.n20 VSUBS 0.01328f
C85 VTAIL.n21 VSUBS 1.29411f
C86 VTAIL.n22 VSUBS 0.012543f
C87 VTAIL.t6 VSUBS 0.063995f
C88 VTAIL.n23 VSUBS 0.199022f
C89 VTAIL.n24 VSUBS 0.022301f
C90 VTAIL.n25 VSUBS 0.022235f
C91 VTAIL.n26 VSUBS 0.029646f
C92 VTAIL.n27 VSUBS 0.01328f
C93 VTAIL.n28 VSUBS 0.012543f
C94 VTAIL.n29 VSUBS 0.023341f
C95 VTAIL.n30 VSUBS 0.023341f
C96 VTAIL.n31 VSUBS 0.012543f
C97 VTAIL.n32 VSUBS 0.01328f
C98 VTAIL.n33 VSUBS 0.029646f
C99 VTAIL.n34 VSUBS 0.029646f
C100 VTAIL.n35 VSUBS 0.01328f
C101 VTAIL.n36 VSUBS 0.012543f
C102 VTAIL.n37 VSUBS 0.023341f
C103 VTAIL.n38 VSUBS 0.023341f
C104 VTAIL.n39 VSUBS 0.012543f
C105 VTAIL.n40 VSUBS 0.012543f
C106 VTAIL.n41 VSUBS 0.01328f
C107 VTAIL.n42 VSUBS 0.029646f
C108 VTAIL.n43 VSUBS 0.029646f
C109 VTAIL.n44 VSUBS 0.029646f
C110 VTAIL.n45 VSUBS 0.012912f
C111 VTAIL.n46 VSUBS 0.012543f
C112 VTAIL.n47 VSUBS 0.023341f
C113 VTAIL.n48 VSUBS 0.023341f
C114 VTAIL.n49 VSUBS 0.012543f
C115 VTAIL.n50 VSUBS 0.01328f
C116 VTAIL.n51 VSUBS 0.029646f
C117 VTAIL.n52 VSUBS 0.029646f
C118 VTAIL.n53 VSUBS 0.01328f
C119 VTAIL.n54 VSUBS 0.012543f
C120 VTAIL.n55 VSUBS 0.023341f
C121 VTAIL.n56 VSUBS 0.023341f
C122 VTAIL.n57 VSUBS 0.012543f
C123 VTAIL.n58 VSUBS 0.01328f
C124 VTAIL.n59 VSUBS 0.029646f
C125 VTAIL.n60 VSUBS 0.029646f
C126 VTAIL.n61 VSUBS 0.01328f
C127 VTAIL.n62 VSUBS 0.012543f
C128 VTAIL.n63 VSUBS 0.023341f
C129 VTAIL.n64 VSUBS 0.023341f
C130 VTAIL.n65 VSUBS 0.012543f
C131 VTAIL.n66 VSUBS 0.01328f
C132 VTAIL.n67 VSUBS 0.029646f
C133 VTAIL.n68 VSUBS 0.07009f
C134 VTAIL.n69 VSUBS 0.01328f
C135 VTAIL.n70 VSUBS 0.012543f
C136 VTAIL.n71 VSUBS 0.050126f
C137 VTAIL.n72 VSUBS 0.035051f
C138 VTAIL.n73 VSUBS 0.157666f
C139 VTAIL.n74 VSUBS 0.025154f
C140 VTAIL.n75 VSUBS 0.023341f
C141 VTAIL.n76 VSUBS 0.012543f
C142 VTAIL.n77 VSUBS 0.029646f
C143 VTAIL.n78 VSUBS 0.01328f
C144 VTAIL.n79 VSUBS 0.023341f
C145 VTAIL.n80 VSUBS 0.012543f
C146 VTAIL.n81 VSUBS 0.029646f
C147 VTAIL.n82 VSUBS 0.01328f
C148 VTAIL.n83 VSUBS 0.023341f
C149 VTAIL.n84 VSUBS 0.012543f
C150 VTAIL.n85 VSUBS 0.029646f
C151 VTAIL.n86 VSUBS 0.012912f
C152 VTAIL.n87 VSUBS 0.023341f
C153 VTAIL.n88 VSUBS 0.01328f
C154 VTAIL.n89 VSUBS 0.029646f
C155 VTAIL.n90 VSUBS 0.01328f
C156 VTAIL.n91 VSUBS 0.023341f
C157 VTAIL.n92 VSUBS 0.012543f
C158 VTAIL.n93 VSUBS 0.029646f
C159 VTAIL.n94 VSUBS 0.01328f
C160 VTAIL.n95 VSUBS 1.29411f
C161 VTAIL.n96 VSUBS 0.012543f
C162 VTAIL.t2 VSUBS 0.063995f
C163 VTAIL.n97 VSUBS 0.199022f
C164 VTAIL.n98 VSUBS 0.022301f
C165 VTAIL.n99 VSUBS 0.022235f
C166 VTAIL.n100 VSUBS 0.029646f
C167 VTAIL.n101 VSUBS 0.01328f
C168 VTAIL.n102 VSUBS 0.012543f
C169 VTAIL.n103 VSUBS 0.023341f
C170 VTAIL.n104 VSUBS 0.023341f
C171 VTAIL.n105 VSUBS 0.012543f
C172 VTAIL.n106 VSUBS 0.01328f
C173 VTAIL.n107 VSUBS 0.029646f
C174 VTAIL.n108 VSUBS 0.029646f
C175 VTAIL.n109 VSUBS 0.01328f
C176 VTAIL.n110 VSUBS 0.012543f
C177 VTAIL.n111 VSUBS 0.023341f
C178 VTAIL.n112 VSUBS 0.023341f
C179 VTAIL.n113 VSUBS 0.012543f
C180 VTAIL.n114 VSUBS 0.012543f
C181 VTAIL.n115 VSUBS 0.01328f
C182 VTAIL.n116 VSUBS 0.029646f
C183 VTAIL.n117 VSUBS 0.029646f
C184 VTAIL.n118 VSUBS 0.029646f
C185 VTAIL.n119 VSUBS 0.012912f
C186 VTAIL.n120 VSUBS 0.012543f
C187 VTAIL.n121 VSUBS 0.023341f
C188 VTAIL.n122 VSUBS 0.023341f
C189 VTAIL.n123 VSUBS 0.012543f
C190 VTAIL.n124 VSUBS 0.01328f
C191 VTAIL.n125 VSUBS 0.029646f
C192 VTAIL.n126 VSUBS 0.029646f
C193 VTAIL.n127 VSUBS 0.01328f
C194 VTAIL.n128 VSUBS 0.012543f
C195 VTAIL.n129 VSUBS 0.023341f
C196 VTAIL.n130 VSUBS 0.023341f
C197 VTAIL.n131 VSUBS 0.012543f
C198 VTAIL.n132 VSUBS 0.01328f
C199 VTAIL.n133 VSUBS 0.029646f
C200 VTAIL.n134 VSUBS 0.029646f
C201 VTAIL.n135 VSUBS 0.01328f
C202 VTAIL.n136 VSUBS 0.012543f
C203 VTAIL.n137 VSUBS 0.023341f
C204 VTAIL.n138 VSUBS 0.023341f
C205 VTAIL.n139 VSUBS 0.012543f
C206 VTAIL.n140 VSUBS 0.01328f
C207 VTAIL.n141 VSUBS 0.029646f
C208 VTAIL.n142 VSUBS 0.07009f
C209 VTAIL.n143 VSUBS 0.01328f
C210 VTAIL.n144 VSUBS 0.012543f
C211 VTAIL.n145 VSUBS 0.050126f
C212 VTAIL.n146 VSUBS 0.035051f
C213 VTAIL.n147 VSUBS 0.253462f
C214 VTAIL.n148 VSUBS 0.025154f
C215 VTAIL.n149 VSUBS 0.023341f
C216 VTAIL.n150 VSUBS 0.012543f
C217 VTAIL.n151 VSUBS 0.029646f
C218 VTAIL.n152 VSUBS 0.01328f
C219 VTAIL.n153 VSUBS 0.023341f
C220 VTAIL.n154 VSUBS 0.012543f
C221 VTAIL.n155 VSUBS 0.029646f
C222 VTAIL.n156 VSUBS 0.01328f
C223 VTAIL.n157 VSUBS 0.023341f
C224 VTAIL.n158 VSUBS 0.012543f
C225 VTAIL.n159 VSUBS 0.029646f
C226 VTAIL.n160 VSUBS 0.012912f
C227 VTAIL.n161 VSUBS 0.023341f
C228 VTAIL.n162 VSUBS 0.01328f
C229 VTAIL.n163 VSUBS 0.029646f
C230 VTAIL.n164 VSUBS 0.01328f
C231 VTAIL.n165 VSUBS 0.023341f
C232 VTAIL.n166 VSUBS 0.012543f
C233 VTAIL.n167 VSUBS 0.029646f
C234 VTAIL.n168 VSUBS 0.01328f
C235 VTAIL.n169 VSUBS 1.29411f
C236 VTAIL.n170 VSUBS 0.012543f
C237 VTAIL.t0 VSUBS 0.063995f
C238 VTAIL.n171 VSUBS 0.199022f
C239 VTAIL.n172 VSUBS 0.022301f
C240 VTAIL.n173 VSUBS 0.022235f
C241 VTAIL.n174 VSUBS 0.029646f
C242 VTAIL.n175 VSUBS 0.01328f
C243 VTAIL.n176 VSUBS 0.012543f
C244 VTAIL.n177 VSUBS 0.023341f
C245 VTAIL.n178 VSUBS 0.023341f
C246 VTAIL.n179 VSUBS 0.012543f
C247 VTAIL.n180 VSUBS 0.01328f
C248 VTAIL.n181 VSUBS 0.029646f
C249 VTAIL.n182 VSUBS 0.029646f
C250 VTAIL.n183 VSUBS 0.01328f
C251 VTAIL.n184 VSUBS 0.012543f
C252 VTAIL.n185 VSUBS 0.023341f
C253 VTAIL.n186 VSUBS 0.023341f
C254 VTAIL.n187 VSUBS 0.012543f
C255 VTAIL.n188 VSUBS 0.012543f
C256 VTAIL.n189 VSUBS 0.01328f
C257 VTAIL.n190 VSUBS 0.029646f
C258 VTAIL.n191 VSUBS 0.029646f
C259 VTAIL.n192 VSUBS 0.029646f
C260 VTAIL.n193 VSUBS 0.012912f
C261 VTAIL.n194 VSUBS 0.012543f
C262 VTAIL.n195 VSUBS 0.023341f
C263 VTAIL.n196 VSUBS 0.023341f
C264 VTAIL.n197 VSUBS 0.012543f
C265 VTAIL.n198 VSUBS 0.01328f
C266 VTAIL.n199 VSUBS 0.029646f
C267 VTAIL.n200 VSUBS 0.029646f
C268 VTAIL.n201 VSUBS 0.01328f
C269 VTAIL.n202 VSUBS 0.012543f
C270 VTAIL.n203 VSUBS 0.023341f
C271 VTAIL.n204 VSUBS 0.023341f
C272 VTAIL.n205 VSUBS 0.012543f
C273 VTAIL.n206 VSUBS 0.01328f
C274 VTAIL.n207 VSUBS 0.029646f
C275 VTAIL.n208 VSUBS 0.029646f
C276 VTAIL.n209 VSUBS 0.01328f
C277 VTAIL.n210 VSUBS 0.012543f
C278 VTAIL.n211 VSUBS 0.023341f
C279 VTAIL.n212 VSUBS 0.023341f
C280 VTAIL.n213 VSUBS 0.012543f
C281 VTAIL.n214 VSUBS 0.01328f
C282 VTAIL.n215 VSUBS 0.029646f
C283 VTAIL.n216 VSUBS 0.07009f
C284 VTAIL.n217 VSUBS 0.01328f
C285 VTAIL.n218 VSUBS 0.012543f
C286 VTAIL.n219 VSUBS 0.050126f
C287 VTAIL.n220 VSUBS 0.035051f
C288 VTAIL.n221 VSUBS 1.60695f
C289 VTAIL.n222 VSUBS 0.025154f
C290 VTAIL.n223 VSUBS 0.023341f
C291 VTAIL.n224 VSUBS 0.012543f
C292 VTAIL.n225 VSUBS 0.029646f
C293 VTAIL.n226 VSUBS 0.01328f
C294 VTAIL.n227 VSUBS 0.023341f
C295 VTAIL.n228 VSUBS 0.012543f
C296 VTAIL.n229 VSUBS 0.029646f
C297 VTAIL.n230 VSUBS 0.01328f
C298 VTAIL.n231 VSUBS 0.023341f
C299 VTAIL.n232 VSUBS 0.012543f
C300 VTAIL.n233 VSUBS 0.029646f
C301 VTAIL.n234 VSUBS 0.012912f
C302 VTAIL.n235 VSUBS 0.023341f
C303 VTAIL.n236 VSUBS 0.012912f
C304 VTAIL.n237 VSUBS 0.012543f
C305 VTAIL.n238 VSUBS 0.029646f
C306 VTAIL.n239 VSUBS 0.029646f
C307 VTAIL.n240 VSUBS 0.01328f
C308 VTAIL.n241 VSUBS 0.023341f
C309 VTAIL.n242 VSUBS 0.012543f
C310 VTAIL.n243 VSUBS 0.029646f
C311 VTAIL.n244 VSUBS 0.01328f
C312 VTAIL.n245 VSUBS 1.29411f
C313 VTAIL.n246 VSUBS 0.012543f
C314 VTAIL.t7 VSUBS 0.063995f
C315 VTAIL.n247 VSUBS 0.199022f
C316 VTAIL.n248 VSUBS 0.022301f
C317 VTAIL.n249 VSUBS 0.022235f
C318 VTAIL.n250 VSUBS 0.029646f
C319 VTAIL.n251 VSUBS 0.01328f
C320 VTAIL.n252 VSUBS 0.012543f
C321 VTAIL.n253 VSUBS 0.023341f
C322 VTAIL.n254 VSUBS 0.023341f
C323 VTAIL.n255 VSUBS 0.012543f
C324 VTAIL.n256 VSUBS 0.01328f
C325 VTAIL.n257 VSUBS 0.029646f
C326 VTAIL.n258 VSUBS 0.029646f
C327 VTAIL.n259 VSUBS 0.01328f
C328 VTAIL.n260 VSUBS 0.012543f
C329 VTAIL.n261 VSUBS 0.023341f
C330 VTAIL.n262 VSUBS 0.023341f
C331 VTAIL.n263 VSUBS 0.012543f
C332 VTAIL.n264 VSUBS 0.01328f
C333 VTAIL.n265 VSUBS 0.029646f
C334 VTAIL.n266 VSUBS 0.029646f
C335 VTAIL.n267 VSUBS 0.01328f
C336 VTAIL.n268 VSUBS 0.012543f
C337 VTAIL.n269 VSUBS 0.023341f
C338 VTAIL.n270 VSUBS 0.023341f
C339 VTAIL.n271 VSUBS 0.012543f
C340 VTAIL.n272 VSUBS 0.01328f
C341 VTAIL.n273 VSUBS 0.029646f
C342 VTAIL.n274 VSUBS 0.029646f
C343 VTAIL.n275 VSUBS 0.01328f
C344 VTAIL.n276 VSUBS 0.012543f
C345 VTAIL.n277 VSUBS 0.023341f
C346 VTAIL.n278 VSUBS 0.023341f
C347 VTAIL.n279 VSUBS 0.012543f
C348 VTAIL.n280 VSUBS 0.01328f
C349 VTAIL.n281 VSUBS 0.029646f
C350 VTAIL.n282 VSUBS 0.029646f
C351 VTAIL.n283 VSUBS 0.01328f
C352 VTAIL.n284 VSUBS 0.012543f
C353 VTAIL.n285 VSUBS 0.023341f
C354 VTAIL.n286 VSUBS 0.023341f
C355 VTAIL.n287 VSUBS 0.012543f
C356 VTAIL.n288 VSUBS 0.01328f
C357 VTAIL.n289 VSUBS 0.029646f
C358 VTAIL.n290 VSUBS 0.07009f
C359 VTAIL.n291 VSUBS 0.01328f
C360 VTAIL.n292 VSUBS 0.012543f
C361 VTAIL.n293 VSUBS 0.050126f
C362 VTAIL.n294 VSUBS 0.035051f
C363 VTAIL.n295 VSUBS 1.60695f
C364 VTAIL.n296 VSUBS 0.025154f
C365 VTAIL.n297 VSUBS 0.023341f
C366 VTAIL.n298 VSUBS 0.012543f
C367 VTAIL.n299 VSUBS 0.029646f
C368 VTAIL.n300 VSUBS 0.01328f
C369 VTAIL.n301 VSUBS 0.023341f
C370 VTAIL.n302 VSUBS 0.012543f
C371 VTAIL.n303 VSUBS 0.029646f
C372 VTAIL.n304 VSUBS 0.01328f
C373 VTAIL.n305 VSUBS 0.023341f
C374 VTAIL.n306 VSUBS 0.012543f
C375 VTAIL.n307 VSUBS 0.029646f
C376 VTAIL.n308 VSUBS 0.012912f
C377 VTAIL.n309 VSUBS 0.023341f
C378 VTAIL.n310 VSUBS 0.012912f
C379 VTAIL.n311 VSUBS 0.012543f
C380 VTAIL.n312 VSUBS 0.029646f
C381 VTAIL.n313 VSUBS 0.029646f
C382 VTAIL.n314 VSUBS 0.01328f
C383 VTAIL.n315 VSUBS 0.023341f
C384 VTAIL.n316 VSUBS 0.012543f
C385 VTAIL.n317 VSUBS 0.029646f
C386 VTAIL.n318 VSUBS 0.01328f
C387 VTAIL.n319 VSUBS 1.29411f
C388 VTAIL.n320 VSUBS 0.012543f
C389 VTAIL.t4 VSUBS 0.063995f
C390 VTAIL.n321 VSUBS 0.199022f
C391 VTAIL.n322 VSUBS 0.022301f
C392 VTAIL.n323 VSUBS 0.022235f
C393 VTAIL.n324 VSUBS 0.029646f
C394 VTAIL.n325 VSUBS 0.01328f
C395 VTAIL.n326 VSUBS 0.012543f
C396 VTAIL.n327 VSUBS 0.023341f
C397 VTAIL.n328 VSUBS 0.023341f
C398 VTAIL.n329 VSUBS 0.012543f
C399 VTAIL.n330 VSUBS 0.01328f
C400 VTAIL.n331 VSUBS 0.029646f
C401 VTAIL.n332 VSUBS 0.029646f
C402 VTAIL.n333 VSUBS 0.01328f
C403 VTAIL.n334 VSUBS 0.012543f
C404 VTAIL.n335 VSUBS 0.023341f
C405 VTAIL.n336 VSUBS 0.023341f
C406 VTAIL.n337 VSUBS 0.012543f
C407 VTAIL.n338 VSUBS 0.01328f
C408 VTAIL.n339 VSUBS 0.029646f
C409 VTAIL.n340 VSUBS 0.029646f
C410 VTAIL.n341 VSUBS 0.01328f
C411 VTAIL.n342 VSUBS 0.012543f
C412 VTAIL.n343 VSUBS 0.023341f
C413 VTAIL.n344 VSUBS 0.023341f
C414 VTAIL.n345 VSUBS 0.012543f
C415 VTAIL.n346 VSUBS 0.01328f
C416 VTAIL.n347 VSUBS 0.029646f
C417 VTAIL.n348 VSUBS 0.029646f
C418 VTAIL.n349 VSUBS 0.01328f
C419 VTAIL.n350 VSUBS 0.012543f
C420 VTAIL.n351 VSUBS 0.023341f
C421 VTAIL.n352 VSUBS 0.023341f
C422 VTAIL.n353 VSUBS 0.012543f
C423 VTAIL.n354 VSUBS 0.01328f
C424 VTAIL.n355 VSUBS 0.029646f
C425 VTAIL.n356 VSUBS 0.029646f
C426 VTAIL.n357 VSUBS 0.01328f
C427 VTAIL.n358 VSUBS 0.012543f
C428 VTAIL.n359 VSUBS 0.023341f
C429 VTAIL.n360 VSUBS 0.023341f
C430 VTAIL.n361 VSUBS 0.012543f
C431 VTAIL.n362 VSUBS 0.01328f
C432 VTAIL.n363 VSUBS 0.029646f
C433 VTAIL.n364 VSUBS 0.07009f
C434 VTAIL.n365 VSUBS 0.01328f
C435 VTAIL.n366 VSUBS 0.012543f
C436 VTAIL.n367 VSUBS 0.050126f
C437 VTAIL.n368 VSUBS 0.035051f
C438 VTAIL.n369 VSUBS 0.253462f
C439 VTAIL.n370 VSUBS 0.025154f
C440 VTAIL.n371 VSUBS 0.023341f
C441 VTAIL.n372 VSUBS 0.012543f
C442 VTAIL.n373 VSUBS 0.029646f
C443 VTAIL.n374 VSUBS 0.01328f
C444 VTAIL.n375 VSUBS 0.023341f
C445 VTAIL.n376 VSUBS 0.012543f
C446 VTAIL.n377 VSUBS 0.029646f
C447 VTAIL.n378 VSUBS 0.01328f
C448 VTAIL.n379 VSUBS 0.023341f
C449 VTAIL.n380 VSUBS 0.012543f
C450 VTAIL.n381 VSUBS 0.029646f
C451 VTAIL.n382 VSUBS 0.012912f
C452 VTAIL.n383 VSUBS 0.023341f
C453 VTAIL.n384 VSUBS 0.012912f
C454 VTAIL.n385 VSUBS 0.012543f
C455 VTAIL.n386 VSUBS 0.029646f
C456 VTAIL.n387 VSUBS 0.029646f
C457 VTAIL.n388 VSUBS 0.01328f
C458 VTAIL.n389 VSUBS 0.023341f
C459 VTAIL.n390 VSUBS 0.012543f
C460 VTAIL.n391 VSUBS 0.029646f
C461 VTAIL.n392 VSUBS 0.01328f
C462 VTAIL.n393 VSUBS 1.29411f
C463 VTAIL.n394 VSUBS 0.012543f
C464 VTAIL.t1 VSUBS 0.063995f
C465 VTAIL.n395 VSUBS 0.199022f
C466 VTAIL.n396 VSUBS 0.022301f
C467 VTAIL.n397 VSUBS 0.022235f
C468 VTAIL.n398 VSUBS 0.029646f
C469 VTAIL.n399 VSUBS 0.01328f
C470 VTAIL.n400 VSUBS 0.012543f
C471 VTAIL.n401 VSUBS 0.023341f
C472 VTAIL.n402 VSUBS 0.023341f
C473 VTAIL.n403 VSUBS 0.012543f
C474 VTAIL.n404 VSUBS 0.01328f
C475 VTAIL.n405 VSUBS 0.029646f
C476 VTAIL.n406 VSUBS 0.029646f
C477 VTAIL.n407 VSUBS 0.01328f
C478 VTAIL.n408 VSUBS 0.012543f
C479 VTAIL.n409 VSUBS 0.023341f
C480 VTAIL.n410 VSUBS 0.023341f
C481 VTAIL.n411 VSUBS 0.012543f
C482 VTAIL.n412 VSUBS 0.01328f
C483 VTAIL.n413 VSUBS 0.029646f
C484 VTAIL.n414 VSUBS 0.029646f
C485 VTAIL.n415 VSUBS 0.01328f
C486 VTAIL.n416 VSUBS 0.012543f
C487 VTAIL.n417 VSUBS 0.023341f
C488 VTAIL.n418 VSUBS 0.023341f
C489 VTAIL.n419 VSUBS 0.012543f
C490 VTAIL.n420 VSUBS 0.01328f
C491 VTAIL.n421 VSUBS 0.029646f
C492 VTAIL.n422 VSUBS 0.029646f
C493 VTAIL.n423 VSUBS 0.01328f
C494 VTAIL.n424 VSUBS 0.012543f
C495 VTAIL.n425 VSUBS 0.023341f
C496 VTAIL.n426 VSUBS 0.023341f
C497 VTAIL.n427 VSUBS 0.012543f
C498 VTAIL.n428 VSUBS 0.01328f
C499 VTAIL.n429 VSUBS 0.029646f
C500 VTAIL.n430 VSUBS 0.029646f
C501 VTAIL.n431 VSUBS 0.01328f
C502 VTAIL.n432 VSUBS 0.012543f
C503 VTAIL.n433 VSUBS 0.023341f
C504 VTAIL.n434 VSUBS 0.023341f
C505 VTAIL.n435 VSUBS 0.012543f
C506 VTAIL.n436 VSUBS 0.01328f
C507 VTAIL.n437 VSUBS 0.029646f
C508 VTAIL.n438 VSUBS 0.07009f
C509 VTAIL.n439 VSUBS 0.01328f
C510 VTAIL.n440 VSUBS 0.012543f
C511 VTAIL.n441 VSUBS 0.050126f
C512 VTAIL.n442 VSUBS 0.035051f
C513 VTAIL.n443 VSUBS 0.253462f
C514 VTAIL.n444 VSUBS 0.025154f
C515 VTAIL.n445 VSUBS 0.023341f
C516 VTAIL.n446 VSUBS 0.012543f
C517 VTAIL.n447 VSUBS 0.029646f
C518 VTAIL.n448 VSUBS 0.01328f
C519 VTAIL.n449 VSUBS 0.023341f
C520 VTAIL.n450 VSUBS 0.012543f
C521 VTAIL.n451 VSUBS 0.029646f
C522 VTAIL.n452 VSUBS 0.01328f
C523 VTAIL.n453 VSUBS 0.023341f
C524 VTAIL.n454 VSUBS 0.012543f
C525 VTAIL.n455 VSUBS 0.029646f
C526 VTAIL.n456 VSUBS 0.012912f
C527 VTAIL.n457 VSUBS 0.023341f
C528 VTAIL.n458 VSUBS 0.012912f
C529 VTAIL.n459 VSUBS 0.012543f
C530 VTAIL.n460 VSUBS 0.029646f
C531 VTAIL.n461 VSUBS 0.029646f
C532 VTAIL.n462 VSUBS 0.01328f
C533 VTAIL.n463 VSUBS 0.023341f
C534 VTAIL.n464 VSUBS 0.012543f
C535 VTAIL.n465 VSUBS 0.029646f
C536 VTAIL.n466 VSUBS 0.01328f
C537 VTAIL.n467 VSUBS 1.29411f
C538 VTAIL.n468 VSUBS 0.012543f
C539 VTAIL.t3 VSUBS 0.063995f
C540 VTAIL.n469 VSUBS 0.199022f
C541 VTAIL.n470 VSUBS 0.022301f
C542 VTAIL.n471 VSUBS 0.022235f
C543 VTAIL.n472 VSUBS 0.029646f
C544 VTAIL.n473 VSUBS 0.01328f
C545 VTAIL.n474 VSUBS 0.012543f
C546 VTAIL.n475 VSUBS 0.023341f
C547 VTAIL.n476 VSUBS 0.023341f
C548 VTAIL.n477 VSUBS 0.012543f
C549 VTAIL.n478 VSUBS 0.01328f
C550 VTAIL.n479 VSUBS 0.029646f
C551 VTAIL.n480 VSUBS 0.029646f
C552 VTAIL.n481 VSUBS 0.01328f
C553 VTAIL.n482 VSUBS 0.012543f
C554 VTAIL.n483 VSUBS 0.023341f
C555 VTAIL.n484 VSUBS 0.023341f
C556 VTAIL.n485 VSUBS 0.012543f
C557 VTAIL.n486 VSUBS 0.01328f
C558 VTAIL.n487 VSUBS 0.029646f
C559 VTAIL.n488 VSUBS 0.029646f
C560 VTAIL.n489 VSUBS 0.01328f
C561 VTAIL.n490 VSUBS 0.012543f
C562 VTAIL.n491 VSUBS 0.023341f
C563 VTAIL.n492 VSUBS 0.023341f
C564 VTAIL.n493 VSUBS 0.012543f
C565 VTAIL.n494 VSUBS 0.01328f
C566 VTAIL.n495 VSUBS 0.029646f
C567 VTAIL.n496 VSUBS 0.029646f
C568 VTAIL.n497 VSUBS 0.01328f
C569 VTAIL.n498 VSUBS 0.012543f
C570 VTAIL.n499 VSUBS 0.023341f
C571 VTAIL.n500 VSUBS 0.023341f
C572 VTAIL.n501 VSUBS 0.012543f
C573 VTAIL.n502 VSUBS 0.01328f
C574 VTAIL.n503 VSUBS 0.029646f
C575 VTAIL.n504 VSUBS 0.029646f
C576 VTAIL.n505 VSUBS 0.01328f
C577 VTAIL.n506 VSUBS 0.012543f
C578 VTAIL.n507 VSUBS 0.023341f
C579 VTAIL.n508 VSUBS 0.023341f
C580 VTAIL.n509 VSUBS 0.012543f
C581 VTAIL.n510 VSUBS 0.01328f
C582 VTAIL.n511 VSUBS 0.029646f
C583 VTAIL.n512 VSUBS 0.07009f
C584 VTAIL.n513 VSUBS 0.01328f
C585 VTAIL.n514 VSUBS 0.012543f
C586 VTAIL.n515 VSUBS 0.050126f
C587 VTAIL.n516 VSUBS 0.035051f
C588 VTAIL.n517 VSUBS 1.60695f
C589 VTAIL.n518 VSUBS 0.025154f
C590 VTAIL.n519 VSUBS 0.023341f
C591 VTAIL.n520 VSUBS 0.012543f
C592 VTAIL.n521 VSUBS 0.029646f
C593 VTAIL.n522 VSUBS 0.01328f
C594 VTAIL.n523 VSUBS 0.023341f
C595 VTAIL.n524 VSUBS 0.012543f
C596 VTAIL.n525 VSUBS 0.029646f
C597 VTAIL.n526 VSUBS 0.01328f
C598 VTAIL.n527 VSUBS 0.023341f
C599 VTAIL.n528 VSUBS 0.012543f
C600 VTAIL.n529 VSUBS 0.029646f
C601 VTAIL.n530 VSUBS 0.012912f
C602 VTAIL.n531 VSUBS 0.023341f
C603 VTAIL.n532 VSUBS 0.01328f
C604 VTAIL.n533 VSUBS 0.029646f
C605 VTAIL.n534 VSUBS 0.01328f
C606 VTAIL.n535 VSUBS 0.023341f
C607 VTAIL.n536 VSUBS 0.012543f
C608 VTAIL.n537 VSUBS 0.029646f
C609 VTAIL.n538 VSUBS 0.01328f
C610 VTAIL.n539 VSUBS 1.29411f
C611 VTAIL.n540 VSUBS 0.012543f
C612 VTAIL.t5 VSUBS 0.063995f
C613 VTAIL.n541 VSUBS 0.199022f
C614 VTAIL.n542 VSUBS 0.022301f
C615 VTAIL.n543 VSUBS 0.022235f
C616 VTAIL.n544 VSUBS 0.029646f
C617 VTAIL.n545 VSUBS 0.01328f
C618 VTAIL.n546 VSUBS 0.012543f
C619 VTAIL.n547 VSUBS 0.023341f
C620 VTAIL.n548 VSUBS 0.023341f
C621 VTAIL.n549 VSUBS 0.012543f
C622 VTAIL.n550 VSUBS 0.01328f
C623 VTAIL.n551 VSUBS 0.029646f
C624 VTAIL.n552 VSUBS 0.029646f
C625 VTAIL.n553 VSUBS 0.01328f
C626 VTAIL.n554 VSUBS 0.012543f
C627 VTAIL.n555 VSUBS 0.023341f
C628 VTAIL.n556 VSUBS 0.023341f
C629 VTAIL.n557 VSUBS 0.012543f
C630 VTAIL.n558 VSUBS 0.012543f
C631 VTAIL.n559 VSUBS 0.01328f
C632 VTAIL.n560 VSUBS 0.029646f
C633 VTAIL.n561 VSUBS 0.029646f
C634 VTAIL.n562 VSUBS 0.029646f
C635 VTAIL.n563 VSUBS 0.012912f
C636 VTAIL.n564 VSUBS 0.012543f
C637 VTAIL.n565 VSUBS 0.023341f
C638 VTAIL.n566 VSUBS 0.023341f
C639 VTAIL.n567 VSUBS 0.012543f
C640 VTAIL.n568 VSUBS 0.01328f
C641 VTAIL.n569 VSUBS 0.029646f
C642 VTAIL.n570 VSUBS 0.029646f
C643 VTAIL.n571 VSUBS 0.01328f
C644 VTAIL.n572 VSUBS 0.012543f
C645 VTAIL.n573 VSUBS 0.023341f
C646 VTAIL.n574 VSUBS 0.023341f
C647 VTAIL.n575 VSUBS 0.012543f
C648 VTAIL.n576 VSUBS 0.01328f
C649 VTAIL.n577 VSUBS 0.029646f
C650 VTAIL.n578 VSUBS 0.029646f
C651 VTAIL.n579 VSUBS 0.01328f
C652 VTAIL.n580 VSUBS 0.012543f
C653 VTAIL.n581 VSUBS 0.023341f
C654 VTAIL.n582 VSUBS 0.023341f
C655 VTAIL.n583 VSUBS 0.012543f
C656 VTAIL.n584 VSUBS 0.01328f
C657 VTAIL.n585 VSUBS 0.029646f
C658 VTAIL.n586 VSUBS 0.07009f
C659 VTAIL.n587 VSUBS 0.01328f
C660 VTAIL.n588 VSUBS 0.012543f
C661 VTAIL.n589 VSUBS 0.050126f
C662 VTAIL.n590 VSUBS 0.035051f
C663 VTAIL.n591 VSUBS 1.5024f
C664 VN.t2 VSUBS 3.42501f
C665 VN.t0 VSUBS 3.4176f
C666 VN.n0 VSUBS 2.17182f
C667 VN.t1 VSUBS 3.42501f
C668 VN.t3 VSUBS 3.4176f
C669 VN.n1 VSUBS 3.96352f
C670 B.n0 VSUBS 0.005653f
C671 B.n1 VSUBS 0.005653f
C672 B.n2 VSUBS 0.00836f
C673 B.n3 VSUBS 0.006407f
C674 B.n4 VSUBS 0.006407f
C675 B.n5 VSUBS 0.006407f
C676 B.n6 VSUBS 0.006407f
C677 B.n7 VSUBS 0.006407f
C678 B.n8 VSUBS 0.006407f
C679 B.n9 VSUBS 0.006407f
C680 B.n10 VSUBS 0.006407f
C681 B.n11 VSUBS 0.006407f
C682 B.n12 VSUBS 0.006407f
C683 B.n13 VSUBS 0.006407f
C684 B.n14 VSUBS 0.006407f
C685 B.n15 VSUBS 0.006407f
C686 B.n16 VSUBS 0.006407f
C687 B.n17 VSUBS 0.006407f
C688 B.n18 VSUBS 0.006407f
C689 B.n19 VSUBS 0.014786f
C690 B.n20 VSUBS 0.006407f
C691 B.n21 VSUBS 0.006407f
C692 B.n22 VSUBS 0.006407f
C693 B.n23 VSUBS 0.006407f
C694 B.n24 VSUBS 0.006407f
C695 B.n25 VSUBS 0.006407f
C696 B.n26 VSUBS 0.006407f
C697 B.n27 VSUBS 0.006407f
C698 B.n28 VSUBS 0.006407f
C699 B.n29 VSUBS 0.006407f
C700 B.n30 VSUBS 0.006407f
C701 B.n31 VSUBS 0.006407f
C702 B.n32 VSUBS 0.006407f
C703 B.n33 VSUBS 0.006407f
C704 B.n34 VSUBS 0.006407f
C705 B.n35 VSUBS 0.006407f
C706 B.n36 VSUBS 0.006407f
C707 B.n37 VSUBS 0.006407f
C708 B.n38 VSUBS 0.006407f
C709 B.n39 VSUBS 0.006407f
C710 B.n40 VSUBS 0.006407f
C711 B.n41 VSUBS 0.006407f
C712 B.n42 VSUBS 0.004428f
C713 B.n43 VSUBS 0.006407f
C714 B.t4 VSUBS 0.222888f
C715 B.t5 VSUBS 0.254033f
C716 B.t3 VSUBS 1.54172f
C717 B.n44 VSUBS 0.400217f
C718 B.n45 VSUBS 0.24899f
C719 B.n46 VSUBS 0.014843f
C720 B.n47 VSUBS 0.006407f
C721 B.n48 VSUBS 0.006407f
C722 B.n49 VSUBS 0.006407f
C723 B.n50 VSUBS 0.006407f
C724 B.t7 VSUBS 0.222891f
C725 B.t8 VSUBS 0.254036f
C726 B.t6 VSUBS 1.54172f
C727 B.n51 VSUBS 0.400214f
C728 B.n52 VSUBS 0.248987f
C729 B.n53 VSUBS 0.006407f
C730 B.n54 VSUBS 0.006407f
C731 B.n55 VSUBS 0.006407f
C732 B.n56 VSUBS 0.006407f
C733 B.n57 VSUBS 0.006407f
C734 B.n58 VSUBS 0.006407f
C735 B.n59 VSUBS 0.006407f
C736 B.n60 VSUBS 0.006407f
C737 B.n61 VSUBS 0.006407f
C738 B.n62 VSUBS 0.006407f
C739 B.n63 VSUBS 0.006407f
C740 B.n64 VSUBS 0.006407f
C741 B.n65 VSUBS 0.006407f
C742 B.n66 VSUBS 0.006407f
C743 B.n67 VSUBS 0.006407f
C744 B.n68 VSUBS 0.006407f
C745 B.n69 VSUBS 0.006407f
C746 B.n70 VSUBS 0.006407f
C747 B.n71 VSUBS 0.006407f
C748 B.n72 VSUBS 0.006407f
C749 B.n73 VSUBS 0.006407f
C750 B.n74 VSUBS 0.006407f
C751 B.n75 VSUBS 0.014786f
C752 B.n76 VSUBS 0.006407f
C753 B.n77 VSUBS 0.006407f
C754 B.n78 VSUBS 0.006407f
C755 B.n79 VSUBS 0.006407f
C756 B.n80 VSUBS 0.006407f
C757 B.n81 VSUBS 0.006407f
C758 B.n82 VSUBS 0.006407f
C759 B.n83 VSUBS 0.006407f
C760 B.n84 VSUBS 0.006407f
C761 B.n85 VSUBS 0.006407f
C762 B.n86 VSUBS 0.006407f
C763 B.n87 VSUBS 0.006407f
C764 B.n88 VSUBS 0.006407f
C765 B.n89 VSUBS 0.006407f
C766 B.n90 VSUBS 0.006407f
C767 B.n91 VSUBS 0.006407f
C768 B.n92 VSUBS 0.006407f
C769 B.n93 VSUBS 0.006407f
C770 B.n94 VSUBS 0.006407f
C771 B.n95 VSUBS 0.006407f
C772 B.n96 VSUBS 0.006407f
C773 B.n97 VSUBS 0.006407f
C774 B.n98 VSUBS 0.006407f
C775 B.n99 VSUBS 0.006407f
C776 B.n100 VSUBS 0.006407f
C777 B.n101 VSUBS 0.006407f
C778 B.n102 VSUBS 0.006407f
C779 B.n103 VSUBS 0.006407f
C780 B.n104 VSUBS 0.006407f
C781 B.n105 VSUBS 0.006407f
C782 B.n106 VSUBS 0.006407f
C783 B.n107 VSUBS 0.006407f
C784 B.n108 VSUBS 0.006407f
C785 B.n109 VSUBS 0.006407f
C786 B.n110 VSUBS 0.006407f
C787 B.n111 VSUBS 0.014416f
C788 B.n112 VSUBS 0.006407f
C789 B.n113 VSUBS 0.006407f
C790 B.n114 VSUBS 0.006407f
C791 B.n115 VSUBS 0.006407f
C792 B.n116 VSUBS 0.006407f
C793 B.n117 VSUBS 0.006407f
C794 B.n118 VSUBS 0.006407f
C795 B.n119 VSUBS 0.006407f
C796 B.n120 VSUBS 0.006407f
C797 B.n121 VSUBS 0.006407f
C798 B.n122 VSUBS 0.006407f
C799 B.n123 VSUBS 0.006407f
C800 B.n124 VSUBS 0.006407f
C801 B.n125 VSUBS 0.006407f
C802 B.n126 VSUBS 0.006407f
C803 B.n127 VSUBS 0.006407f
C804 B.n128 VSUBS 0.006407f
C805 B.n129 VSUBS 0.006407f
C806 B.n130 VSUBS 0.006407f
C807 B.n131 VSUBS 0.006407f
C808 B.n132 VSUBS 0.006407f
C809 B.n133 VSUBS 0.006407f
C810 B.n134 VSUBS 0.006407f
C811 B.t2 VSUBS 0.222891f
C812 B.t1 VSUBS 0.254036f
C813 B.t0 VSUBS 1.54172f
C814 B.n135 VSUBS 0.400214f
C815 B.n136 VSUBS 0.248987f
C816 B.n137 VSUBS 0.006407f
C817 B.n138 VSUBS 0.006407f
C818 B.n139 VSUBS 0.006407f
C819 B.n140 VSUBS 0.006407f
C820 B.t11 VSUBS 0.222888f
C821 B.t10 VSUBS 0.254033f
C822 B.t9 VSUBS 1.54172f
C823 B.n141 VSUBS 0.400217f
C824 B.n142 VSUBS 0.24899f
C825 B.n143 VSUBS 0.006407f
C826 B.n144 VSUBS 0.006407f
C827 B.n145 VSUBS 0.006407f
C828 B.n146 VSUBS 0.006407f
C829 B.n147 VSUBS 0.006407f
C830 B.n148 VSUBS 0.006407f
C831 B.n149 VSUBS 0.006407f
C832 B.n150 VSUBS 0.006407f
C833 B.n151 VSUBS 0.006407f
C834 B.n152 VSUBS 0.006407f
C835 B.n153 VSUBS 0.006407f
C836 B.n154 VSUBS 0.006407f
C837 B.n155 VSUBS 0.006407f
C838 B.n156 VSUBS 0.006407f
C839 B.n157 VSUBS 0.006407f
C840 B.n158 VSUBS 0.006407f
C841 B.n159 VSUBS 0.006407f
C842 B.n160 VSUBS 0.006407f
C843 B.n161 VSUBS 0.006407f
C844 B.n162 VSUBS 0.006407f
C845 B.n163 VSUBS 0.006407f
C846 B.n164 VSUBS 0.006407f
C847 B.n165 VSUBS 0.015174f
C848 B.n166 VSUBS 0.006407f
C849 B.n167 VSUBS 0.006407f
C850 B.n168 VSUBS 0.006407f
C851 B.n169 VSUBS 0.006407f
C852 B.n170 VSUBS 0.006407f
C853 B.n171 VSUBS 0.006407f
C854 B.n172 VSUBS 0.006407f
C855 B.n173 VSUBS 0.006407f
C856 B.n174 VSUBS 0.006407f
C857 B.n175 VSUBS 0.006407f
C858 B.n176 VSUBS 0.006407f
C859 B.n177 VSUBS 0.006407f
C860 B.n178 VSUBS 0.006407f
C861 B.n179 VSUBS 0.006407f
C862 B.n180 VSUBS 0.006407f
C863 B.n181 VSUBS 0.006407f
C864 B.n182 VSUBS 0.006407f
C865 B.n183 VSUBS 0.006407f
C866 B.n184 VSUBS 0.006407f
C867 B.n185 VSUBS 0.006407f
C868 B.n186 VSUBS 0.006407f
C869 B.n187 VSUBS 0.006407f
C870 B.n188 VSUBS 0.006407f
C871 B.n189 VSUBS 0.006407f
C872 B.n190 VSUBS 0.006407f
C873 B.n191 VSUBS 0.006407f
C874 B.n192 VSUBS 0.006407f
C875 B.n193 VSUBS 0.006407f
C876 B.n194 VSUBS 0.006407f
C877 B.n195 VSUBS 0.006407f
C878 B.n196 VSUBS 0.006407f
C879 B.n197 VSUBS 0.006407f
C880 B.n198 VSUBS 0.006407f
C881 B.n199 VSUBS 0.006407f
C882 B.n200 VSUBS 0.006407f
C883 B.n201 VSUBS 0.006407f
C884 B.n202 VSUBS 0.006407f
C885 B.n203 VSUBS 0.006407f
C886 B.n204 VSUBS 0.006407f
C887 B.n205 VSUBS 0.006407f
C888 B.n206 VSUBS 0.006407f
C889 B.n207 VSUBS 0.006407f
C890 B.n208 VSUBS 0.006407f
C891 B.n209 VSUBS 0.006407f
C892 B.n210 VSUBS 0.006407f
C893 B.n211 VSUBS 0.006407f
C894 B.n212 VSUBS 0.006407f
C895 B.n213 VSUBS 0.006407f
C896 B.n214 VSUBS 0.006407f
C897 B.n215 VSUBS 0.006407f
C898 B.n216 VSUBS 0.006407f
C899 B.n217 VSUBS 0.006407f
C900 B.n218 VSUBS 0.006407f
C901 B.n219 VSUBS 0.006407f
C902 B.n220 VSUBS 0.006407f
C903 B.n221 VSUBS 0.006407f
C904 B.n222 VSUBS 0.006407f
C905 B.n223 VSUBS 0.006407f
C906 B.n224 VSUBS 0.006407f
C907 B.n225 VSUBS 0.006407f
C908 B.n226 VSUBS 0.006407f
C909 B.n227 VSUBS 0.006407f
C910 B.n228 VSUBS 0.006407f
C911 B.n229 VSUBS 0.006407f
C912 B.n230 VSUBS 0.006407f
C913 B.n231 VSUBS 0.006407f
C914 B.n232 VSUBS 0.014786f
C915 B.n233 VSUBS 0.014786f
C916 B.n234 VSUBS 0.015174f
C917 B.n235 VSUBS 0.006407f
C918 B.n236 VSUBS 0.006407f
C919 B.n237 VSUBS 0.006407f
C920 B.n238 VSUBS 0.006407f
C921 B.n239 VSUBS 0.006407f
C922 B.n240 VSUBS 0.006407f
C923 B.n241 VSUBS 0.006407f
C924 B.n242 VSUBS 0.006407f
C925 B.n243 VSUBS 0.006407f
C926 B.n244 VSUBS 0.006407f
C927 B.n245 VSUBS 0.006407f
C928 B.n246 VSUBS 0.006407f
C929 B.n247 VSUBS 0.006407f
C930 B.n248 VSUBS 0.006407f
C931 B.n249 VSUBS 0.006407f
C932 B.n250 VSUBS 0.006407f
C933 B.n251 VSUBS 0.006407f
C934 B.n252 VSUBS 0.006407f
C935 B.n253 VSUBS 0.006407f
C936 B.n254 VSUBS 0.006407f
C937 B.n255 VSUBS 0.006407f
C938 B.n256 VSUBS 0.006407f
C939 B.n257 VSUBS 0.006407f
C940 B.n258 VSUBS 0.006407f
C941 B.n259 VSUBS 0.006407f
C942 B.n260 VSUBS 0.006407f
C943 B.n261 VSUBS 0.006407f
C944 B.n262 VSUBS 0.006407f
C945 B.n263 VSUBS 0.006407f
C946 B.n264 VSUBS 0.006407f
C947 B.n265 VSUBS 0.006407f
C948 B.n266 VSUBS 0.006407f
C949 B.n267 VSUBS 0.006407f
C950 B.n268 VSUBS 0.006407f
C951 B.n269 VSUBS 0.006407f
C952 B.n270 VSUBS 0.006407f
C953 B.n271 VSUBS 0.006407f
C954 B.n272 VSUBS 0.006407f
C955 B.n273 VSUBS 0.006407f
C956 B.n274 VSUBS 0.006407f
C957 B.n275 VSUBS 0.006407f
C958 B.n276 VSUBS 0.006407f
C959 B.n277 VSUBS 0.006407f
C960 B.n278 VSUBS 0.006407f
C961 B.n279 VSUBS 0.006407f
C962 B.n280 VSUBS 0.006407f
C963 B.n281 VSUBS 0.006407f
C964 B.n282 VSUBS 0.006407f
C965 B.n283 VSUBS 0.006407f
C966 B.n284 VSUBS 0.006407f
C967 B.n285 VSUBS 0.006407f
C968 B.n286 VSUBS 0.006407f
C969 B.n287 VSUBS 0.006407f
C970 B.n288 VSUBS 0.006407f
C971 B.n289 VSUBS 0.006407f
C972 B.n290 VSUBS 0.006407f
C973 B.n291 VSUBS 0.006407f
C974 B.n292 VSUBS 0.006407f
C975 B.n293 VSUBS 0.006407f
C976 B.n294 VSUBS 0.006407f
C977 B.n295 VSUBS 0.006407f
C978 B.n296 VSUBS 0.006407f
C979 B.n297 VSUBS 0.006407f
C980 B.n298 VSUBS 0.006407f
C981 B.n299 VSUBS 0.006407f
C982 B.n300 VSUBS 0.006407f
C983 B.n301 VSUBS 0.006407f
C984 B.n302 VSUBS 0.004428f
C985 B.n303 VSUBS 0.014843f
C986 B.n304 VSUBS 0.005182f
C987 B.n305 VSUBS 0.006407f
C988 B.n306 VSUBS 0.006407f
C989 B.n307 VSUBS 0.006407f
C990 B.n308 VSUBS 0.006407f
C991 B.n309 VSUBS 0.006407f
C992 B.n310 VSUBS 0.006407f
C993 B.n311 VSUBS 0.006407f
C994 B.n312 VSUBS 0.006407f
C995 B.n313 VSUBS 0.006407f
C996 B.n314 VSUBS 0.006407f
C997 B.n315 VSUBS 0.006407f
C998 B.n316 VSUBS 0.005182f
C999 B.n317 VSUBS 0.014843f
C1000 B.n318 VSUBS 0.004428f
C1001 B.n319 VSUBS 0.006407f
C1002 B.n320 VSUBS 0.006407f
C1003 B.n321 VSUBS 0.006407f
C1004 B.n322 VSUBS 0.006407f
C1005 B.n323 VSUBS 0.006407f
C1006 B.n324 VSUBS 0.006407f
C1007 B.n325 VSUBS 0.006407f
C1008 B.n326 VSUBS 0.006407f
C1009 B.n327 VSUBS 0.006407f
C1010 B.n328 VSUBS 0.006407f
C1011 B.n329 VSUBS 0.006407f
C1012 B.n330 VSUBS 0.006407f
C1013 B.n331 VSUBS 0.006407f
C1014 B.n332 VSUBS 0.006407f
C1015 B.n333 VSUBS 0.006407f
C1016 B.n334 VSUBS 0.006407f
C1017 B.n335 VSUBS 0.006407f
C1018 B.n336 VSUBS 0.006407f
C1019 B.n337 VSUBS 0.006407f
C1020 B.n338 VSUBS 0.006407f
C1021 B.n339 VSUBS 0.006407f
C1022 B.n340 VSUBS 0.006407f
C1023 B.n341 VSUBS 0.006407f
C1024 B.n342 VSUBS 0.006407f
C1025 B.n343 VSUBS 0.006407f
C1026 B.n344 VSUBS 0.006407f
C1027 B.n345 VSUBS 0.006407f
C1028 B.n346 VSUBS 0.006407f
C1029 B.n347 VSUBS 0.006407f
C1030 B.n348 VSUBS 0.006407f
C1031 B.n349 VSUBS 0.006407f
C1032 B.n350 VSUBS 0.006407f
C1033 B.n351 VSUBS 0.006407f
C1034 B.n352 VSUBS 0.006407f
C1035 B.n353 VSUBS 0.006407f
C1036 B.n354 VSUBS 0.006407f
C1037 B.n355 VSUBS 0.006407f
C1038 B.n356 VSUBS 0.006407f
C1039 B.n357 VSUBS 0.006407f
C1040 B.n358 VSUBS 0.006407f
C1041 B.n359 VSUBS 0.006407f
C1042 B.n360 VSUBS 0.006407f
C1043 B.n361 VSUBS 0.006407f
C1044 B.n362 VSUBS 0.006407f
C1045 B.n363 VSUBS 0.006407f
C1046 B.n364 VSUBS 0.006407f
C1047 B.n365 VSUBS 0.006407f
C1048 B.n366 VSUBS 0.006407f
C1049 B.n367 VSUBS 0.006407f
C1050 B.n368 VSUBS 0.006407f
C1051 B.n369 VSUBS 0.006407f
C1052 B.n370 VSUBS 0.006407f
C1053 B.n371 VSUBS 0.006407f
C1054 B.n372 VSUBS 0.006407f
C1055 B.n373 VSUBS 0.006407f
C1056 B.n374 VSUBS 0.006407f
C1057 B.n375 VSUBS 0.006407f
C1058 B.n376 VSUBS 0.006407f
C1059 B.n377 VSUBS 0.006407f
C1060 B.n378 VSUBS 0.006407f
C1061 B.n379 VSUBS 0.006407f
C1062 B.n380 VSUBS 0.006407f
C1063 B.n381 VSUBS 0.006407f
C1064 B.n382 VSUBS 0.006407f
C1065 B.n383 VSUBS 0.006407f
C1066 B.n384 VSUBS 0.006407f
C1067 B.n385 VSUBS 0.006407f
C1068 B.n386 VSUBS 0.015174f
C1069 B.n387 VSUBS 0.014786f
C1070 B.n388 VSUBS 0.015544f
C1071 B.n389 VSUBS 0.006407f
C1072 B.n390 VSUBS 0.006407f
C1073 B.n391 VSUBS 0.006407f
C1074 B.n392 VSUBS 0.006407f
C1075 B.n393 VSUBS 0.006407f
C1076 B.n394 VSUBS 0.006407f
C1077 B.n395 VSUBS 0.006407f
C1078 B.n396 VSUBS 0.006407f
C1079 B.n397 VSUBS 0.006407f
C1080 B.n398 VSUBS 0.006407f
C1081 B.n399 VSUBS 0.006407f
C1082 B.n400 VSUBS 0.006407f
C1083 B.n401 VSUBS 0.006407f
C1084 B.n402 VSUBS 0.006407f
C1085 B.n403 VSUBS 0.006407f
C1086 B.n404 VSUBS 0.006407f
C1087 B.n405 VSUBS 0.006407f
C1088 B.n406 VSUBS 0.006407f
C1089 B.n407 VSUBS 0.006407f
C1090 B.n408 VSUBS 0.006407f
C1091 B.n409 VSUBS 0.006407f
C1092 B.n410 VSUBS 0.006407f
C1093 B.n411 VSUBS 0.006407f
C1094 B.n412 VSUBS 0.006407f
C1095 B.n413 VSUBS 0.006407f
C1096 B.n414 VSUBS 0.006407f
C1097 B.n415 VSUBS 0.006407f
C1098 B.n416 VSUBS 0.006407f
C1099 B.n417 VSUBS 0.006407f
C1100 B.n418 VSUBS 0.006407f
C1101 B.n419 VSUBS 0.006407f
C1102 B.n420 VSUBS 0.006407f
C1103 B.n421 VSUBS 0.006407f
C1104 B.n422 VSUBS 0.006407f
C1105 B.n423 VSUBS 0.006407f
C1106 B.n424 VSUBS 0.006407f
C1107 B.n425 VSUBS 0.006407f
C1108 B.n426 VSUBS 0.006407f
C1109 B.n427 VSUBS 0.006407f
C1110 B.n428 VSUBS 0.006407f
C1111 B.n429 VSUBS 0.006407f
C1112 B.n430 VSUBS 0.006407f
C1113 B.n431 VSUBS 0.006407f
C1114 B.n432 VSUBS 0.006407f
C1115 B.n433 VSUBS 0.006407f
C1116 B.n434 VSUBS 0.006407f
C1117 B.n435 VSUBS 0.006407f
C1118 B.n436 VSUBS 0.006407f
C1119 B.n437 VSUBS 0.006407f
C1120 B.n438 VSUBS 0.006407f
C1121 B.n439 VSUBS 0.006407f
C1122 B.n440 VSUBS 0.006407f
C1123 B.n441 VSUBS 0.006407f
C1124 B.n442 VSUBS 0.006407f
C1125 B.n443 VSUBS 0.006407f
C1126 B.n444 VSUBS 0.006407f
C1127 B.n445 VSUBS 0.006407f
C1128 B.n446 VSUBS 0.006407f
C1129 B.n447 VSUBS 0.006407f
C1130 B.n448 VSUBS 0.006407f
C1131 B.n449 VSUBS 0.006407f
C1132 B.n450 VSUBS 0.006407f
C1133 B.n451 VSUBS 0.006407f
C1134 B.n452 VSUBS 0.006407f
C1135 B.n453 VSUBS 0.006407f
C1136 B.n454 VSUBS 0.006407f
C1137 B.n455 VSUBS 0.006407f
C1138 B.n456 VSUBS 0.006407f
C1139 B.n457 VSUBS 0.006407f
C1140 B.n458 VSUBS 0.006407f
C1141 B.n459 VSUBS 0.006407f
C1142 B.n460 VSUBS 0.006407f
C1143 B.n461 VSUBS 0.006407f
C1144 B.n462 VSUBS 0.006407f
C1145 B.n463 VSUBS 0.006407f
C1146 B.n464 VSUBS 0.006407f
C1147 B.n465 VSUBS 0.006407f
C1148 B.n466 VSUBS 0.006407f
C1149 B.n467 VSUBS 0.006407f
C1150 B.n468 VSUBS 0.006407f
C1151 B.n469 VSUBS 0.006407f
C1152 B.n470 VSUBS 0.006407f
C1153 B.n471 VSUBS 0.006407f
C1154 B.n472 VSUBS 0.006407f
C1155 B.n473 VSUBS 0.006407f
C1156 B.n474 VSUBS 0.006407f
C1157 B.n475 VSUBS 0.006407f
C1158 B.n476 VSUBS 0.006407f
C1159 B.n477 VSUBS 0.006407f
C1160 B.n478 VSUBS 0.006407f
C1161 B.n479 VSUBS 0.006407f
C1162 B.n480 VSUBS 0.006407f
C1163 B.n481 VSUBS 0.006407f
C1164 B.n482 VSUBS 0.006407f
C1165 B.n483 VSUBS 0.006407f
C1166 B.n484 VSUBS 0.006407f
C1167 B.n485 VSUBS 0.006407f
C1168 B.n486 VSUBS 0.006407f
C1169 B.n487 VSUBS 0.006407f
C1170 B.n488 VSUBS 0.006407f
C1171 B.n489 VSUBS 0.006407f
C1172 B.n490 VSUBS 0.006407f
C1173 B.n491 VSUBS 0.006407f
C1174 B.n492 VSUBS 0.006407f
C1175 B.n493 VSUBS 0.006407f
C1176 B.n494 VSUBS 0.014786f
C1177 B.n495 VSUBS 0.015174f
C1178 B.n496 VSUBS 0.015174f
C1179 B.n497 VSUBS 0.006407f
C1180 B.n498 VSUBS 0.006407f
C1181 B.n499 VSUBS 0.006407f
C1182 B.n500 VSUBS 0.006407f
C1183 B.n501 VSUBS 0.006407f
C1184 B.n502 VSUBS 0.006407f
C1185 B.n503 VSUBS 0.006407f
C1186 B.n504 VSUBS 0.006407f
C1187 B.n505 VSUBS 0.006407f
C1188 B.n506 VSUBS 0.006407f
C1189 B.n507 VSUBS 0.006407f
C1190 B.n508 VSUBS 0.006407f
C1191 B.n509 VSUBS 0.006407f
C1192 B.n510 VSUBS 0.006407f
C1193 B.n511 VSUBS 0.006407f
C1194 B.n512 VSUBS 0.006407f
C1195 B.n513 VSUBS 0.006407f
C1196 B.n514 VSUBS 0.006407f
C1197 B.n515 VSUBS 0.006407f
C1198 B.n516 VSUBS 0.006407f
C1199 B.n517 VSUBS 0.006407f
C1200 B.n518 VSUBS 0.006407f
C1201 B.n519 VSUBS 0.006407f
C1202 B.n520 VSUBS 0.006407f
C1203 B.n521 VSUBS 0.006407f
C1204 B.n522 VSUBS 0.006407f
C1205 B.n523 VSUBS 0.006407f
C1206 B.n524 VSUBS 0.006407f
C1207 B.n525 VSUBS 0.006407f
C1208 B.n526 VSUBS 0.006407f
C1209 B.n527 VSUBS 0.006407f
C1210 B.n528 VSUBS 0.006407f
C1211 B.n529 VSUBS 0.006407f
C1212 B.n530 VSUBS 0.006407f
C1213 B.n531 VSUBS 0.006407f
C1214 B.n532 VSUBS 0.006407f
C1215 B.n533 VSUBS 0.006407f
C1216 B.n534 VSUBS 0.006407f
C1217 B.n535 VSUBS 0.006407f
C1218 B.n536 VSUBS 0.006407f
C1219 B.n537 VSUBS 0.006407f
C1220 B.n538 VSUBS 0.006407f
C1221 B.n539 VSUBS 0.006407f
C1222 B.n540 VSUBS 0.006407f
C1223 B.n541 VSUBS 0.006407f
C1224 B.n542 VSUBS 0.006407f
C1225 B.n543 VSUBS 0.006407f
C1226 B.n544 VSUBS 0.006407f
C1227 B.n545 VSUBS 0.006407f
C1228 B.n546 VSUBS 0.006407f
C1229 B.n547 VSUBS 0.006407f
C1230 B.n548 VSUBS 0.006407f
C1231 B.n549 VSUBS 0.006407f
C1232 B.n550 VSUBS 0.006407f
C1233 B.n551 VSUBS 0.006407f
C1234 B.n552 VSUBS 0.006407f
C1235 B.n553 VSUBS 0.006407f
C1236 B.n554 VSUBS 0.006407f
C1237 B.n555 VSUBS 0.006407f
C1238 B.n556 VSUBS 0.006407f
C1239 B.n557 VSUBS 0.006407f
C1240 B.n558 VSUBS 0.006407f
C1241 B.n559 VSUBS 0.006407f
C1242 B.n560 VSUBS 0.006407f
C1243 B.n561 VSUBS 0.006407f
C1244 B.n562 VSUBS 0.006407f
C1245 B.n563 VSUBS 0.004428f
C1246 B.n564 VSUBS 0.014843f
C1247 B.n565 VSUBS 0.005182f
C1248 B.n566 VSUBS 0.006407f
C1249 B.n567 VSUBS 0.006407f
C1250 B.n568 VSUBS 0.006407f
C1251 B.n569 VSUBS 0.006407f
C1252 B.n570 VSUBS 0.006407f
C1253 B.n571 VSUBS 0.006407f
C1254 B.n572 VSUBS 0.006407f
C1255 B.n573 VSUBS 0.006407f
C1256 B.n574 VSUBS 0.006407f
C1257 B.n575 VSUBS 0.006407f
C1258 B.n576 VSUBS 0.006407f
C1259 B.n577 VSUBS 0.005182f
C1260 B.n578 VSUBS 0.006407f
C1261 B.n579 VSUBS 0.006407f
C1262 B.n580 VSUBS 0.006407f
C1263 B.n581 VSUBS 0.006407f
C1264 B.n582 VSUBS 0.006407f
C1265 B.n583 VSUBS 0.006407f
C1266 B.n584 VSUBS 0.006407f
C1267 B.n585 VSUBS 0.006407f
C1268 B.n586 VSUBS 0.006407f
C1269 B.n587 VSUBS 0.006407f
C1270 B.n588 VSUBS 0.006407f
C1271 B.n589 VSUBS 0.006407f
C1272 B.n590 VSUBS 0.006407f
C1273 B.n591 VSUBS 0.006407f
C1274 B.n592 VSUBS 0.006407f
C1275 B.n593 VSUBS 0.006407f
C1276 B.n594 VSUBS 0.006407f
C1277 B.n595 VSUBS 0.006407f
C1278 B.n596 VSUBS 0.006407f
C1279 B.n597 VSUBS 0.006407f
C1280 B.n598 VSUBS 0.006407f
C1281 B.n599 VSUBS 0.006407f
C1282 B.n600 VSUBS 0.006407f
C1283 B.n601 VSUBS 0.006407f
C1284 B.n602 VSUBS 0.006407f
C1285 B.n603 VSUBS 0.006407f
C1286 B.n604 VSUBS 0.006407f
C1287 B.n605 VSUBS 0.006407f
C1288 B.n606 VSUBS 0.006407f
C1289 B.n607 VSUBS 0.006407f
C1290 B.n608 VSUBS 0.006407f
C1291 B.n609 VSUBS 0.006407f
C1292 B.n610 VSUBS 0.006407f
C1293 B.n611 VSUBS 0.006407f
C1294 B.n612 VSUBS 0.006407f
C1295 B.n613 VSUBS 0.006407f
C1296 B.n614 VSUBS 0.006407f
C1297 B.n615 VSUBS 0.006407f
C1298 B.n616 VSUBS 0.006407f
C1299 B.n617 VSUBS 0.006407f
C1300 B.n618 VSUBS 0.006407f
C1301 B.n619 VSUBS 0.006407f
C1302 B.n620 VSUBS 0.006407f
C1303 B.n621 VSUBS 0.006407f
C1304 B.n622 VSUBS 0.006407f
C1305 B.n623 VSUBS 0.006407f
C1306 B.n624 VSUBS 0.006407f
C1307 B.n625 VSUBS 0.006407f
C1308 B.n626 VSUBS 0.006407f
C1309 B.n627 VSUBS 0.006407f
C1310 B.n628 VSUBS 0.006407f
C1311 B.n629 VSUBS 0.006407f
C1312 B.n630 VSUBS 0.006407f
C1313 B.n631 VSUBS 0.006407f
C1314 B.n632 VSUBS 0.006407f
C1315 B.n633 VSUBS 0.006407f
C1316 B.n634 VSUBS 0.006407f
C1317 B.n635 VSUBS 0.006407f
C1318 B.n636 VSUBS 0.006407f
C1319 B.n637 VSUBS 0.006407f
C1320 B.n638 VSUBS 0.006407f
C1321 B.n639 VSUBS 0.006407f
C1322 B.n640 VSUBS 0.006407f
C1323 B.n641 VSUBS 0.006407f
C1324 B.n642 VSUBS 0.006407f
C1325 B.n643 VSUBS 0.006407f
C1326 B.n644 VSUBS 0.006407f
C1327 B.n645 VSUBS 0.006407f
C1328 B.n646 VSUBS 0.015174f
C1329 B.n647 VSUBS 0.015174f
C1330 B.n648 VSUBS 0.014786f
C1331 B.n649 VSUBS 0.006407f
C1332 B.n650 VSUBS 0.006407f
C1333 B.n651 VSUBS 0.006407f
C1334 B.n652 VSUBS 0.006407f
C1335 B.n653 VSUBS 0.006407f
C1336 B.n654 VSUBS 0.006407f
C1337 B.n655 VSUBS 0.006407f
C1338 B.n656 VSUBS 0.006407f
C1339 B.n657 VSUBS 0.006407f
C1340 B.n658 VSUBS 0.006407f
C1341 B.n659 VSUBS 0.006407f
C1342 B.n660 VSUBS 0.006407f
C1343 B.n661 VSUBS 0.006407f
C1344 B.n662 VSUBS 0.006407f
C1345 B.n663 VSUBS 0.006407f
C1346 B.n664 VSUBS 0.006407f
C1347 B.n665 VSUBS 0.006407f
C1348 B.n666 VSUBS 0.006407f
C1349 B.n667 VSUBS 0.006407f
C1350 B.n668 VSUBS 0.006407f
C1351 B.n669 VSUBS 0.006407f
C1352 B.n670 VSUBS 0.006407f
C1353 B.n671 VSUBS 0.006407f
C1354 B.n672 VSUBS 0.006407f
C1355 B.n673 VSUBS 0.006407f
C1356 B.n674 VSUBS 0.006407f
C1357 B.n675 VSUBS 0.006407f
C1358 B.n676 VSUBS 0.006407f
C1359 B.n677 VSUBS 0.006407f
C1360 B.n678 VSUBS 0.006407f
C1361 B.n679 VSUBS 0.006407f
C1362 B.n680 VSUBS 0.006407f
C1363 B.n681 VSUBS 0.006407f
C1364 B.n682 VSUBS 0.006407f
C1365 B.n683 VSUBS 0.006407f
C1366 B.n684 VSUBS 0.006407f
C1367 B.n685 VSUBS 0.006407f
C1368 B.n686 VSUBS 0.006407f
C1369 B.n687 VSUBS 0.006407f
C1370 B.n688 VSUBS 0.006407f
C1371 B.n689 VSUBS 0.006407f
C1372 B.n690 VSUBS 0.006407f
C1373 B.n691 VSUBS 0.006407f
C1374 B.n692 VSUBS 0.006407f
C1375 B.n693 VSUBS 0.006407f
C1376 B.n694 VSUBS 0.006407f
C1377 B.n695 VSUBS 0.006407f
C1378 B.n696 VSUBS 0.006407f
C1379 B.n697 VSUBS 0.006407f
C1380 B.n698 VSUBS 0.006407f
C1381 B.n699 VSUBS 0.00836f
C1382 B.n700 VSUBS 0.008906f
C1383 B.n701 VSUBS 0.01771f
.ends

