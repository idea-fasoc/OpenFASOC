* NGSPICE file created from diff_pair_sample_0716.ext - technology: sky130A

.subckt diff_pair_sample_0716 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=0 ps=0 w=19.55 l=1.33
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=7.6245 ps=39.88 w=19.55 l=1.33
X2 VDD1.t1 VP.t0 VTAIL.t0 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=7.6245 ps=39.88 w=19.55 l=1.33
X3 VDD1.t0 VP.t1 VTAIL.t1 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=7.6245 ps=39.88 w=19.55 l=1.33
X4 B.t8 B.t6 B.t7 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=0 ps=0 w=19.55 l=1.33
X5 B.t5 B.t3 B.t4 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=0 ps=0 w=19.55 l=1.33
X6 VDD2.t0 VN.t1 VTAIL.t3 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=7.6245 ps=39.88 w=19.55 l=1.33
X7 B.t2 B.t0 B.t1 w_n1634_n4878# sky130_fd_pr__pfet_01v8 ad=7.6245 pd=39.88 as=0 ps=0 w=19.55 l=1.33
R0 B.n472 B.n83 585
R1 B.n474 B.n473 585
R2 B.n475 B.n82 585
R3 B.n477 B.n476 585
R4 B.n478 B.n81 585
R5 B.n480 B.n479 585
R6 B.n481 B.n80 585
R7 B.n483 B.n482 585
R8 B.n484 B.n79 585
R9 B.n486 B.n485 585
R10 B.n487 B.n78 585
R11 B.n489 B.n488 585
R12 B.n490 B.n77 585
R13 B.n492 B.n491 585
R14 B.n493 B.n76 585
R15 B.n495 B.n494 585
R16 B.n496 B.n75 585
R17 B.n498 B.n497 585
R18 B.n499 B.n74 585
R19 B.n501 B.n500 585
R20 B.n502 B.n73 585
R21 B.n504 B.n503 585
R22 B.n505 B.n72 585
R23 B.n507 B.n506 585
R24 B.n508 B.n71 585
R25 B.n510 B.n509 585
R26 B.n511 B.n70 585
R27 B.n513 B.n512 585
R28 B.n514 B.n69 585
R29 B.n516 B.n515 585
R30 B.n517 B.n68 585
R31 B.n519 B.n518 585
R32 B.n520 B.n67 585
R33 B.n522 B.n521 585
R34 B.n523 B.n66 585
R35 B.n525 B.n524 585
R36 B.n526 B.n65 585
R37 B.n528 B.n527 585
R38 B.n529 B.n64 585
R39 B.n531 B.n530 585
R40 B.n532 B.n63 585
R41 B.n534 B.n533 585
R42 B.n535 B.n62 585
R43 B.n537 B.n536 585
R44 B.n538 B.n61 585
R45 B.n540 B.n539 585
R46 B.n541 B.n60 585
R47 B.n543 B.n542 585
R48 B.n544 B.n59 585
R49 B.n546 B.n545 585
R50 B.n547 B.n58 585
R51 B.n549 B.n548 585
R52 B.n550 B.n57 585
R53 B.n552 B.n551 585
R54 B.n553 B.n56 585
R55 B.n555 B.n554 585
R56 B.n556 B.n55 585
R57 B.n558 B.n557 585
R58 B.n559 B.n54 585
R59 B.n561 B.n560 585
R60 B.n562 B.n53 585
R61 B.n564 B.n563 585
R62 B.n565 B.n52 585
R63 B.n567 B.n566 585
R64 B.n569 B.n49 585
R65 B.n571 B.n570 585
R66 B.n572 B.n48 585
R67 B.n574 B.n573 585
R68 B.n575 B.n47 585
R69 B.n577 B.n576 585
R70 B.n578 B.n46 585
R71 B.n580 B.n579 585
R72 B.n581 B.n43 585
R73 B.n584 B.n583 585
R74 B.n585 B.n42 585
R75 B.n587 B.n586 585
R76 B.n588 B.n41 585
R77 B.n590 B.n589 585
R78 B.n591 B.n40 585
R79 B.n593 B.n592 585
R80 B.n594 B.n39 585
R81 B.n596 B.n595 585
R82 B.n597 B.n38 585
R83 B.n599 B.n598 585
R84 B.n600 B.n37 585
R85 B.n602 B.n601 585
R86 B.n603 B.n36 585
R87 B.n605 B.n604 585
R88 B.n606 B.n35 585
R89 B.n608 B.n607 585
R90 B.n609 B.n34 585
R91 B.n611 B.n610 585
R92 B.n612 B.n33 585
R93 B.n614 B.n613 585
R94 B.n615 B.n32 585
R95 B.n617 B.n616 585
R96 B.n618 B.n31 585
R97 B.n620 B.n619 585
R98 B.n621 B.n30 585
R99 B.n623 B.n622 585
R100 B.n624 B.n29 585
R101 B.n626 B.n625 585
R102 B.n627 B.n28 585
R103 B.n629 B.n628 585
R104 B.n630 B.n27 585
R105 B.n632 B.n631 585
R106 B.n633 B.n26 585
R107 B.n635 B.n634 585
R108 B.n636 B.n25 585
R109 B.n638 B.n637 585
R110 B.n639 B.n24 585
R111 B.n641 B.n640 585
R112 B.n642 B.n23 585
R113 B.n644 B.n643 585
R114 B.n645 B.n22 585
R115 B.n647 B.n646 585
R116 B.n648 B.n21 585
R117 B.n650 B.n649 585
R118 B.n651 B.n20 585
R119 B.n653 B.n652 585
R120 B.n654 B.n19 585
R121 B.n656 B.n655 585
R122 B.n657 B.n18 585
R123 B.n659 B.n658 585
R124 B.n660 B.n17 585
R125 B.n662 B.n661 585
R126 B.n663 B.n16 585
R127 B.n665 B.n664 585
R128 B.n666 B.n15 585
R129 B.n668 B.n667 585
R130 B.n669 B.n14 585
R131 B.n671 B.n670 585
R132 B.n672 B.n13 585
R133 B.n674 B.n673 585
R134 B.n675 B.n12 585
R135 B.n677 B.n676 585
R136 B.n678 B.n11 585
R137 B.n471 B.n470 585
R138 B.n469 B.n84 585
R139 B.n468 B.n467 585
R140 B.n466 B.n85 585
R141 B.n465 B.n464 585
R142 B.n463 B.n86 585
R143 B.n462 B.n461 585
R144 B.n460 B.n87 585
R145 B.n459 B.n458 585
R146 B.n457 B.n88 585
R147 B.n456 B.n455 585
R148 B.n454 B.n89 585
R149 B.n453 B.n452 585
R150 B.n451 B.n90 585
R151 B.n450 B.n449 585
R152 B.n448 B.n91 585
R153 B.n447 B.n446 585
R154 B.n445 B.n92 585
R155 B.n444 B.n443 585
R156 B.n442 B.n93 585
R157 B.n441 B.n440 585
R158 B.n439 B.n94 585
R159 B.n438 B.n437 585
R160 B.n436 B.n95 585
R161 B.n435 B.n434 585
R162 B.n433 B.n96 585
R163 B.n432 B.n431 585
R164 B.n430 B.n97 585
R165 B.n429 B.n428 585
R166 B.n427 B.n98 585
R167 B.n426 B.n425 585
R168 B.n424 B.n99 585
R169 B.n423 B.n422 585
R170 B.n421 B.n100 585
R171 B.n420 B.n419 585
R172 B.n418 B.n101 585
R173 B.n417 B.n416 585
R174 B.n210 B.n209 585
R175 B.n211 B.n174 585
R176 B.n213 B.n212 585
R177 B.n214 B.n173 585
R178 B.n216 B.n215 585
R179 B.n217 B.n172 585
R180 B.n219 B.n218 585
R181 B.n220 B.n171 585
R182 B.n222 B.n221 585
R183 B.n223 B.n170 585
R184 B.n225 B.n224 585
R185 B.n226 B.n169 585
R186 B.n228 B.n227 585
R187 B.n229 B.n168 585
R188 B.n231 B.n230 585
R189 B.n232 B.n167 585
R190 B.n234 B.n233 585
R191 B.n235 B.n166 585
R192 B.n237 B.n236 585
R193 B.n238 B.n165 585
R194 B.n240 B.n239 585
R195 B.n241 B.n164 585
R196 B.n243 B.n242 585
R197 B.n244 B.n163 585
R198 B.n246 B.n245 585
R199 B.n247 B.n162 585
R200 B.n249 B.n248 585
R201 B.n250 B.n161 585
R202 B.n252 B.n251 585
R203 B.n253 B.n160 585
R204 B.n255 B.n254 585
R205 B.n256 B.n159 585
R206 B.n258 B.n257 585
R207 B.n259 B.n158 585
R208 B.n261 B.n260 585
R209 B.n262 B.n157 585
R210 B.n264 B.n263 585
R211 B.n265 B.n156 585
R212 B.n267 B.n266 585
R213 B.n268 B.n155 585
R214 B.n270 B.n269 585
R215 B.n271 B.n154 585
R216 B.n273 B.n272 585
R217 B.n274 B.n153 585
R218 B.n276 B.n275 585
R219 B.n277 B.n152 585
R220 B.n279 B.n278 585
R221 B.n280 B.n151 585
R222 B.n282 B.n281 585
R223 B.n283 B.n150 585
R224 B.n285 B.n284 585
R225 B.n286 B.n149 585
R226 B.n288 B.n287 585
R227 B.n289 B.n148 585
R228 B.n291 B.n290 585
R229 B.n292 B.n147 585
R230 B.n294 B.n293 585
R231 B.n295 B.n146 585
R232 B.n297 B.n296 585
R233 B.n298 B.n145 585
R234 B.n300 B.n299 585
R235 B.n301 B.n144 585
R236 B.n303 B.n302 585
R237 B.n304 B.n141 585
R238 B.n307 B.n306 585
R239 B.n308 B.n140 585
R240 B.n310 B.n309 585
R241 B.n311 B.n139 585
R242 B.n313 B.n312 585
R243 B.n314 B.n138 585
R244 B.n316 B.n315 585
R245 B.n317 B.n137 585
R246 B.n319 B.n318 585
R247 B.n321 B.n320 585
R248 B.n322 B.n133 585
R249 B.n324 B.n323 585
R250 B.n325 B.n132 585
R251 B.n327 B.n326 585
R252 B.n328 B.n131 585
R253 B.n330 B.n329 585
R254 B.n331 B.n130 585
R255 B.n333 B.n332 585
R256 B.n334 B.n129 585
R257 B.n336 B.n335 585
R258 B.n337 B.n128 585
R259 B.n339 B.n338 585
R260 B.n340 B.n127 585
R261 B.n342 B.n341 585
R262 B.n343 B.n126 585
R263 B.n345 B.n344 585
R264 B.n346 B.n125 585
R265 B.n348 B.n347 585
R266 B.n349 B.n124 585
R267 B.n351 B.n350 585
R268 B.n352 B.n123 585
R269 B.n354 B.n353 585
R270 B.n355 B.n122 585
R271 B.n357 B.n356 585
R272 B.n358 B.n121 585
R273 B.n360 B.n359 585
R274 B.n361 B.n120 585
R275 B.n363 B.n362 585
R276 B.n364 B.n119 585
R277 B.n366 B.n365 585
R278 B.n367 B.n118 585
R279 B.n369 B.n368 585
R280 B.n370 B.n117 585
R281 B.n372 B.n371 585
R282 B.n373 B.n116 585
R283 B.n375 B.n374 585
R284 B.n376 B.n115 585
R285 B.n378 B.n377 585
R286 B.n379 B.n114 585
R287 B.n381 B.n380 585
R288 B.n382 B.n113 585
R289 B.n384 B.n383 585
R290 B.n385 B.n112 585
R291 B.n387 B.n386 585
R292 B.n388 B.n111 585
R293 B.n390 B.n389 585
R294 B.n391 B.n110 585
R295 B.n393 B.n392 585
R296 B.n394 B.n109 585
R297 B.n396 B.n395 585
R298 B.n397 B.n108 585
R299 B.n399 B.n398 585
R300 B.n400 B.n107 585
R301 B.n402 B.n401 585
R302 B.n403 B.n106 585
R303 B.n405 B.n404 585
R304 B.n406 B.n105 585
R305 B.n408 B.n407 585
R306 B.n409 B.n104 585
R307 B.n411 B.n410 585
R308 B.n412 B.n103 585
R309 B.n414 B.n413 585
R310 B.n415 B.n102 585
R311 B.n208 B.n175 585
R312 B.n207 B.n206 585
R313 B.n205 B.n176 585
R314 B.n204 B.n203 585
R315 B.n202 B.n177 585
R316 B.n201 B.n200 585
R317 B.n199 B.n178 585
R318 B.n198 B.n197 585
R319 B.n196 B.n179 585
R320 B.n195 B.n194 585
R321 B.n193 B.n180 585
R322 B.n192 B.n191 585
R323 B.n190 B.n181 585
R324 B.n189 B.n188 585
R325 B.n187 B.n182 585
R326 B.n186 B.n185 585
R327 B.n184 B.n183 585
R328 B.n2 B.n0 585
R329 B.n705 B.n1 585
R330 B.n704 B.n703 585
R331 B.n702 B.n3 585
R332 B.n701 B.n700 585
R333 B.n699 B.n4 585
R334 B.n698 B.n697 585
R335 B.n696 B.n5 585
R336 B.n695 B.n694 585
R337 B.n693 B.n6 585
R338 B.n692 B.n691 585
R339 B.n690 B.n7 585
R340 B.n689 B.n688 585
R341 B.n687 B.n8 585
R342 B.n686 B.n685 585
R343 B.n684 B.n9 585
R344 B.n683 B.n682 585
R345 B.n681 B.n10 585
R346 B.n680 B.n679 585
R347 B.n707 B.n706 585
R348 B.n134 B.t0 558.997
R349 B.n142 B.t6 558.997
R350 B.n44 B.t3 558.997
R351 B.n50 B.t9 558.997
R352 B.n134 B.t2 543.809
R353 B.n50 B.t10 543.809
R354 B.n142 B.t8 543.809
R355 B.n44 B.t4 543.809
R356 B.n135 B.t1 511.615
R357 B.n51 B.t11 511.615
R358 B.n143 B.t7 511.615
R359 B.n45 B.t5 511.615
R360 B.n210 B.n175 497.305
R361 B.n680 B.n11 497.305
R362 B.n416 B.n415 497.305
R363 B.n470 B.n83 497.305
R364 B.n206 B.n175 163.367
R365 B.n206 B.n205 163.367
R366 B.n205 B.n204 163.367
R367 B.n204 B.n177 163.367
R368 B.n200 B.n177 163.367
R369 B.n200 B.n199 163.367
R370 B.n199 B.n198 163.367
R371 B.n198 B.n179 163.367
R372 B.n194 B.n179 163.367
R373 B.n194 B.n193 163.367
R374 B.n193 B.n192 163.367
R375 B.n192 B.n181 163.367
R376 B.n188 B.n181 163.367
R377 B.n188 B.n187 163.367
R378 B.n187 B.n186 163.367
R379 B.n186 B.n183 163.367
R380 B.n183 B.n2 163.367
R381 B.n706 B.n2 163.367
R382 B.n706 B.n705 163.367
R383 B.n705 B.n704 163.367
R384 B.n704 B.n3 163.367
R385 B.n700 B.n3 163.367
R386 B.n700 B.n699 163.367
R387 B.n699 B.n698 163.367
R388 B.n698 B.n5 163.367
R389 B.n694 B.n5 163.367
R390 B.n694 B.n693 163.367
R391 B.n693 B.n692 163.367
R392 B.n692 B.n7 163.367
R393 B.n688 B.n7 163.367
R394 B.n688 B.n687 163.367
R395 B.n687 B.n686 163.367
R396 B.n686 B.n9 163.367
R397 B.n682 B.n9 163.367
R398 B.n682 B.n681 163.367
R399 B.n681 B.n680 163.367
R400 B.n211 B.n210 163.367
R401 B.n212 B.n211 163.367
R402 B.n212 B.n173 163.367
R403 B.n216 B.n173 163.367
R404 B.n217 B.n216 163.367
R405 B.n218 B.n217 163.367
R406 B.n218 B.n171 163.367
R407 B.n222 B.n171 163.367
R408 B.n223 B.n222 163.367
R409 B.n224 B.n223 163.367
R410 B.n224 B.n169 163.367
R411 B.n228 B.n169 163.367
R412 B.n229 B.n228 163.367
R413 B.n230 B.n229 163.367
R414 B.n230 B.n167 163.367
R415 B.n234 B.n167 163.367
R416 B.n235 B.n234 163.367
R417 B.n236 B.n235 163.367
R418 B.n236 B.n165 163.367
R419 B.n240 B.n165 163.367
R420 B.n241 B.n240 163.367
R421 B.n242 B.n241 163.367
R422 B.n242 B.n163 163.367
R423 B.n246 B.n163 163.367
R424 B.n247 B.n246 163.367
R425 B.n248 B.n247 163.367
R426 B.n248 B.n161 163.367
R427 B.n252 B.n161 163.367
R428 B.n253 B.n252 163.367
R429 B.n254 B.n253 163.367
R430 B.n254 B.n159 163.367
R431 B.n258 B.n159 163.367
R432 B.n259 B.n258 163.367
R433 B.n260 B.n259 163.367
R434 B.n260 B.n157 163.367
R435 B.n264 B.n157 163.367
R436 B.n265 B.n264 163.367
R437 B.n266 B.n265 163.367
R438 B.n266 B.n155 163.367
R439 B.n270 B.n155 163.367
R440 B.n271 B.n270 163.367
R441 B.n272 B.n271 163.367
R442 B.n272 B.n153 163.367
R443 B.n276 B.n153 163.367
R444 B.n277 B.n276 163.367
R445 B.n278 B.n277 163.367
R446 B.n278 B.n151 163.367
R447 B.n282 B.n151 163.367
R448 B.n283 B.n282 163.367
R449 B.n284 B.n283 163.367
R450 B.n284 B.n149 163.367
R451 B.n288 B.n149 163.367
R452 B.n289 B.n288 163.367
R453 B.n290 B.n289 163.367
R454 B.n290 B.n147 163.367
R455 B.n294 B.n147 163.367
R456 B.n295 B.n294 163.367
R457 B.n296 B.n295 163.367
R458 B.n296 B.n145 163.367
R459 B.n300 B.n145 163.367
R460 B.n301 B.n300 163.367
R461 B.n302 B.n301 163.367
R462 B.n302 B.n141 163.367
R463 B.n307 B.n141 163.367
R464 B.n308 B.n307 163.367
R465 B.n309 B.n308 163.367
R466 B.n309 B.n139 163.367
R467 B.n313 B.n139 163.367
R468 B.n314 B.n313 163.367
R469 B.n315 B.n314 163.367
R470 B.n315 B.n137 163.367
R471 B.n319 B.n137 163.367
R472 B.n320 B.n319 163.367
R473 B.n320 B.n133 163.367
R474 B.n324 B.n133 163.367
R475 B.n325 B.n324 163.367
R476 B.n326 B.n325 163.367
R477 B.n326 B.n131 163.367
R478 B.n330 B.n131 163.367
R479 B.n331 B.n330 163.367
R480 B.n332 B.n331 163.367
R481 B.n332 B.n129 163.367
R482 B.n336 B.n129 163.367
R483 B.n337 B.n336 163.367
R484 B.n338 B.n337 163.367
R485 B.n338 B.n127 163.367
R486 B.n342 B.n127 163.367
R487 B.n343 B.n342 163.367
R488 B.n344 B.n343 163.367
R489 B.n344 B.n125 163.367
R490 B.n348 B.n125 163.367
R491 B.n349 B.n348 163.367
R492 B.n350 B.n349 163.367
R493 B.n350 B.n123 163.367
R494 B.n354 B.n123 163.367
R495 B.n355 B.n354 163.367
R496 B.n356 B.n355 163.367
R497 B.n356 B.n121 163.367
R498 B.n360 B.n121 163.367
R499 B.n361 B.n360 163.367
R500 B.n362 B.n361 163.367
R501 B.n362 B.n119 163.367
R502 B.n366 B.n119 163.367
R503 B.n367 B.n366 163.367
R504 B.n368 B.n367 163.367
R505 B.n368 B.n117 163.367
R506 B.n372 B.n117 163.367
R507 B.n373 B.n372 163.367
R508 B.n374 B.n373 163.367
R509 B.n374 B.n115 163.367
R510 B.n378 B.n115 163.367
R511 B.n379 B.n378 163.367
R512 B.n380 B.n379 163.367
R513 B.n380 B.n113 163.367
R514 B.n384 B.n113 163.367
R515 B.n385 B.n384 163.367
R516 B.n386 B.n385 163.367
R517 B.n386 B.n111 163.367
R518 B.n390 B.n111 163.367
R519 B.n391 B.n390 163.367
R520 B.n392 B.n391 163.367
R521 B.n392 B.n109 163.367
R522 B.n396 B.n109 163.367
R523 B.n397 B.n396 163.367
R524 B.n398 B.n397 163.367
R525 B.n398 B.n107 163.367
R526 B.n402 B.n107 163.367
R527 B.n403 B.n402 163.367
R528 B.n404 B.n403 163.367
R529 B.n404 B.n105 163.367
R530 B.n408 B.n105 163.367
R531 B.n409 B.n408 163.367
R532 B.n410 B.n409 163.367
R533 B.n410 B.n103 163.367
R534 B.n414 B.n103 163.367
R535 B.n415 B.n414 163.367
R536 B.n416 B.n101 163.367
R537 B.n420 B.n101 163.367
R538 B.n421 B.n420 163.367
R539 B.n422 B.n421 163.367
R540 B.n422 B.n99 163.367
R541 B.n426 B.n99 163.367
R542 B.n427 B.n426 163.367
R543 B.n428 B.n427 163.367
R544 B.n428 B.n97 163.367
R545 B.n432 B.n97 163.367
R546 B.n433 B.n432 163.367
R547 B.n434 B.n433 163.367
R548 B.n434 B.n95 163.367
R549 B.n438 B.n95 163.367
R550 B.n439 B.n438 163.367
R551 B.n440 B.n439 163.367
R552 B.n440 B.n93 163.367
R553 B.n444 B.n93 163.367
R554 B.n445 B.n444 163.367
R555 B.n446 B.n445 163.367
R556 B.n446 B.n91 163.367
R557 B.n450 B.n91 163.367
R558 B.n451 B.n450 163.367
R559 B.n452 B.n451 163.367
R560 B.n452 B.n89 163.367
R561 B.n456 B.n89 163.367
R562 B.n457 B.n456 163.367
R563 B.n458 B.n457 163.367
R564 B.n458 B.n87 163.367
R565 B.n462 B.n87 163.367
R566 B.n463 B.n462 163.367
R567 B.n464 B.n463 163.367
R568 B.n464 B.n85 163.367
R569 B.n468 B.n85 163.367
R570 B.n469 B.n468 163.367
R571 B.n470 B.n469 163.367
R572 B.n676 B.n11 163.367
R573 B.n676 B.n675 163.367
R574 B.n675 B.n674 163.367
R575 B.n674 B.n13 163.367
R576 B.n670 B.n13 163.367
R577 B.n670 B.n669 163.367
R578 B.n669 B.n668 163.367
R579 B.n668 B.n15 163.367
R580 B.n664 B.n15 163.367
R581 B.n664 B.n663 163.367
R582 B.n663 B.n662 163.367
R583 B.n662 B.n17 163.367
R584 B.n658 B.n17 163.367
R585 B.n658 B.n657 163.367
R586 B.n657 B.n656 163.367
R587 B.n656 B.n19 163.367
R588 B.n652 B.n19 163.367
R589 B.n652 B.n651 163.367
R590 B.n651 B.n650 163.367
R591 B.n650 B.n21 163.367
R592 B.n646 B.n21 163.367
R593 B.n646 B.n645 163.367
R594 B.n645 B.n644 163.367
R595 B.n644 B.n23 163.367
R596 B.n640 B.n23 163.367
R597 B.n640 B.n639 163.367
R598 B.n639 B.n638 163.367
R599 B.n638 B.n25 163.367
R600 B.n634 B.n25 163.367
R601 B.n634 B.n633 163.367
R602 B.n633 B.n632 163.367
R603 B.n632 B.n27 163.367
R604 B.n628 B.n27 163.367
R605 B.n628 B.n627 163.367
R606 B.n627 B.n626 163.367
R607 B.n626 B.n29 163.367
R608 B.n622 B.n29 163.367
R609 B.n622 B.n621 163.367
R610 B.n621 B.n620 163.367
R611 B.n620 B.n31 163.367
R612 B.n616 B.n31 163.367
R613 B.n616 B.n615 163.367
R614 B.n615 B.n614 163.367
R615 B.n614 B.n33 163.367
R616 B.n610 B.n33 163.367
R617 B.n610 B.n609 163.367
R618 B.n609 B.n608 163.367
R619 B.n608 B.n35 163.367
R620 B.n604 B.n35 163.367
R621 B.n604 B.n603 163.367
R622 B.n603 B.n602 163.367
R623 B.n602 B.n37 163.367
R624 B.n598 B.n37 163.367
R625 B.n598 B.n597 163.367
R626 B.n597 B.n596 163.367
R627 B.n596 B.n39 163.367
R628 B.n592 B.n39 163.367
R629 B.n592 B.n591 163.367
R630 B.n591 B.n590 163.367
R631 B.n590 B.n41 163.367
R632 B.n586 B.n41 163.367
R633 B.n586 B.n585 163.367
R634 B.n585 B.n584 163.367
R635 B.n584 B.n43 163.367
R636 B.n579 B.n43 163.367
R637 B.n579 B.n578 163.367
R638 B.n578 B.n577 163.367
R639 B.n577 B.n47 163.367
R640 B.n573 B.n47 163.367
R641 B.n573 B.n572 163.367
R642 B.n572 B.n571 163.367
R643 B.n571 B.n49 163.367
R644 B.n566 B.n49 163.367
R645 B.n566 B.n565 163.367
R646 B.n565 B.n564 163.367
R647 B.n564 B.n53 163.367
R648 B.n560 B.n53 163.367
R649 B.n560 B.n559 163.367
R650 B.n559 B.n558 163.367
R651 B.n558 B.n55 163.367
R652 B.n554 B.n55 163.367
R653 B.n554 B.n553 163.367
R654 B.n553 B.n552 163.367
R655 B.n552 B.n57 163.367
R656 B.n548 B.n57 163.367
R657 B.n548 B.n547 163.367
R658 B.n547 B.n546 163.367
R659 B.n546 B.n59 163.367
R660 B.n542 B.n59 163.367
R661 B.n542 B.n541 163.367
R662 B.n541 B.n540 163.367
R663 B.n540 B.n61 163.367
R664 B.n536 B.n61 163.367
R665 B.n536 B.n535 163.367
R666 B.n535 B.n534 163.367
R667 B.n534 B.n63 163.367
R668 B.n530 B.n63 163.367
R669 B.n530 B.n529 163.367
R670 B.n529 B.n528 163.367
R671 B.n528 B.n65 163.367
R672 B.n524 B.n65 163.367
R673 B.n524 B.n523 163.367
R674 B.n523 B.n522 163.367
R675 B.n522 B.n67 163.367
R676 B.n518 B.n67 163.367
R677 B.n518 B.n517 163.367
R678 B.n517 B.n516 163.367
R679 B.n516 B.n69 163.367
R680 B.n512 B.n69 163.367
R681 B.n512 B.n511 163.367
R682 B.n511 B.n510 163.367
R683 B.n510 B.n71 163.367
R684 B.n506 B.n71 163.367
R685 B.n506 B.n505 163.367
R686 B.n505 B.n504 163.367
R687 B.n504 B.n73 163.367
R688 B.n500 B.n73 163.367
R689 B.n500 B.n499 163.367
R690 B.n499 B.n498 163.367
R691 B.n498 B.n75 163.367
R692 B.n494 B.n75 163.367
R693 B.n494 B.n493 163.367
R694 B.n493 B.n492 163.367
R695 B.n492 B.n77 163.367
R696 B.n488 B.n77 163.367
R697 B.n488 B.n487 163.367
R698 B.n487 B.n486 163.367
R699 B.n486 B.n79 163.367
R700 B.n482 B.n79 163.367
R701 B.n482 B.n481 163.367
R702 B.n481 B.n480 163.367
R703 B.n480 B.n81 163.367
R704 B.n476 B.n81 163.367
R705 B.n476 B.n475 163.367
R706 B.n475 B.n474 163.367
R707 B.n474 B.n83 163.367
R708 B.n136 B.n135 59.5399
R709 B.n305 B.n143 59.5399
R710 B.n582 B.n45 59.5399
R711 B.n568 B.n51 59.5399
R712 B.n679 B.n678 32.3127
R713 B.n472 B.n471 32.3127
R714 B.n417 B.n102 32.3127
R715 B.n209 B.n208 32.3127
R716 B.n135 B.n134 32.1944
R717 B.n143 B.n142 32.1944
R718 B.n45 B.n44 32.1944
R719 B.n51 B.n50 32.1944
R720 B B.n707 18.0485
R721 B.n678 B.n677 10.6151
R722 B.n677 B.n12 10.6151
R723 B.n673 B.n12 10.6151
R724 B.n673 B.n672 10.6151
R725 B.n672 B.n671 10.6151
R726 B.n671 B.n14 10.6151
R727 B.n667 B.n14 10.6151
R728 B.n667 B.n666 10.6151
R729 B.n666 B.n665 10.6151
R730 B.n665 B.n16 10.6151
R731 B.n661 B.n16 10.6151
R732 B.n661 B.n660 10.6151
R733 B.n660 B.n659 10.6151
R734 B.n659 B.n18 10.6151
R735 B.n655 B.n18 10.6151
R736 B.n655 B.n654 10.6151
R737 B.n654 B.n653 10.6151
R738 B.n653 B.n20 10.6151
R739 B.n649 B.n20 10.6151
R740 B.n649 B.n648 10.6151
R741 B.n648 B.n647 10.6151
R742 B.n647 B.n22 10.6151
R743 B.n643 B.n22 10.6151
R744 B.n643 B.n642 10.6151
R745 B.n642 B.n641 10.6151
R746 B.n641 B.n24 10.6151
R747 B.n637 B.n24 10.6151
R748 B.n637 B.n636 10.6151
R749 B.n636 B.n635 10.6151
R750 B.n635 B.n26 10.6151
R751 B.n631 B.n26 10.6151
R752 B.n631 B.n630 10.6151
R753 B.n630 B.n629 10.6151
R754 B.n629 B.n28 10.6151
R755 B.n625 B.n28 10.6151
R756 B.n625 B.n624 10.6151
R757 B.n624 B.n623 10.6151
R758 B.n623 B.n30 10.6151
R759 B.n619 B.n30 10.6151
R760 B.n619 B.n618 10.6151
R761 B.n618 B.n617 10.6151
R762 B.n617 B.n32 10.6151
R763 B.n613 B.n32 10.6151
R764 B.n613 B.n612 10.6151
R765 B.n612 B.n611 10.6151
R766 B.n611 B.n34 10.6151
R767 B.n607 B.n34 10.6151
R768 B.n607 B.n606 10.6151
R769 B.n606 B.n605 10.6151
R770 B.n605 B.n36 10.6151
R771 B.n601 B.n36 10.6151
R772 B.n601 B.n600 10.6151
R773 B.n600 B.n599 10.6151
R774 B.n599 B.n38 10.6151
R775 B.n595 B.n38 10.6151
R776 B.n595 B.n594 10.6151
R777 B.n594 B.n593 10.6151
R778 B.n593 B.n40 10.6151
R779 B.n589 B.n40 10.6151
R780 B.n589 B.n588 10.6151
R781 B.n588 B.n587 10.6151
R782 B.n587 B.n42 10.6151
R783 B.n583 B.n42 10.6151
R784 B.n581 B.n580 10.6151
R785 B.n580 B.n46 10.6151
R786 B.n576 B.n46 10.6151
R787 B.n576 B.n575 10.6151
R788 B.n575 B.n574 10.6151
R789 B.n574 B.n48 10.6151
R790 B.n570 B.n48 10.6151
R791 B.n570 B.n569 10.6151
R792 B.n567 B.n52 10.6151
R793 B.n563 B.n52 10.6151
R794 B.n563 B.n562 10.6151
R795 B.n562 B.n561 10.6151
R796 B.n561 B.n54 10.6151
R797 B.n557 B.n54 10.6151
R798 B.n557 B.n556 10.6151
R799 B.n556 B.n555 10.6151
R800 B.n555 B.n56 10.6151
R801 B.n551 B.n56 10.6151
R802 B.n551 B.n550 10.6151
R803 B.n550 B.n549 10.6151
R804 B.n549 B.n58 10.6151
R805 B.n545 B.n58 10.6151
R806 B.n545 B.n544 10.6151
R807 B.n544 B.n543 10.6151
R808 B.n543 B.n60 10.6151
R809 B.n539 B.n60 10.6151
R810 B.n539 B.n538 10.6151
R811 B.n538 B.n537 10.6151
R812 B.n537 B.n62 10.6151
R813 B.n533 B.n62 10.6151
R814 B.n533 B.n532 10.6151
R815 B.n532 B.n531 10.6151
R816 B.n531 B.n64 10.6151
R817 B.n527 B.n64 10.6151
R818 B.n527 B.n526 10.6151
R819 B.n526 B.n525 10.6151
R820 B.n525 B.n66 10.6151
R821 B.n521 B.n66 10.6151
R822 B.n521 B.n520 10.6151
R823 B.n520 B.n519 10.6151
R824 B.n519 B.n68 10.6151
R825 B.n515 B.n68 10.6151
R826 B.n515 B.n514 10.6151
R827 B.n514 B.n513 10.6151
R828 B.n513 B.n70 10.6151
R829 B.n509 B.n70 10.6151
R830 B.n509 B.n508 10.6151
R831 B.n508 B.n507 10.6151
R832 B.n507 B.n72 10.6151
R833 B.n503 B.n72 10.6151
R834 B.n503 B.n502 10.6151
R835 B.n502 B.n501 10.6151
R836 B.n501 B.n74 10.6151
R837 B.n497 B.n74 10.6151
R838 B.n497 B.n496 10.6151
R839 B.n496 B.n495 10.6151
R840 B.n495 B.n76 10.6151
R841 B.n491 B.n76 10.6151
R842 B.n491 B.n490 10.6151
R843 B.n490 B.n489 10.6151
R844 B.n489 B.n78 10.6151
R845 B.n485 B.n78 10.6151
R846 B.n485 B.n484 10.6151
R847 B.n484 B.n483 10.6151
R848 B.n483 B.n80 10.6151
R849 B.n479 B.n80 10.6151
R850 B.n479 B.n478 10.6151
R851 B.n478 B.n477 10.6151
R852 B.n477 B.n82 10.6151
R853 B.n473 B.n82 10.6151
R854 B.n473 B.n472 10.6151
R855 B.n418 B.n417 10.6151
R856 B.n419 B.n418 10.6151
R857 B.n419 B.n100 10.6151
R858 B.n423 B.n100 10.6151
R859 B.n424 B.n423 10.6151
R860 B.n425 B.n424 10.6151
R861 B.n425 B.n98 10.6151
R862 B.n429 B.n98 10.6151
R863 B.n430 B.n429 10.6151
R864 B.n431 B.n430 10.6151
R865 B.n431 B.n96 10.6151
R866 B.n435 B.n96 10.6151
R867 B.n436 B.n435 10.6151
R868 B.n437 B.n436 10.6151
R869 B.n437 B.n94 10.6151
R870 B.n441 B.n94 10.6151
R871 B.n442 B.n441 10.6151
R872 B.n443 B.n442 10.6151
R873 B.n443 B.n92 10.6151
R874 B.n447 B.n92 10.6151
R875 B.n448 B.n447 10.6151
R876 B.n449 B.n448 10.6151
R877 B.n449 B.n90 10.6151
R878 B.n453 B.n90 10.6151
R879 B.n454 B.n453 10.6151
R880 B.n455 B.n454 10.6151
R881 B.n455 B.n88 10.6151
R882 B.n459 B.n88 10.6151
R883 B.n460 B.n459 10.6151
R884 B.n461 B.n460 10.6151
R885 B.n461 B.n86 10.6151
R886 B.n465 B.n86 10.6151
R887 B.n466 B.n465 10.6151
R888 B.n467 B.n466 10.6151
R889 B.n467 B.n84 10.6151
R890 B.n471 B.n84 10.6151
R891 B.n209 B.n174 10.6151
R892 B.n213 B.n174 10.6151
R893 B.n214 B.n213 10.6151
R894 B.n215 B.n214 10.6151
R895 B.n215 B.n172 10.6151
R896 B.n219 B.n172 10.6151
R897 B.n220 B.n219 10.6151
R898 B.n221 B.n220 10.6151
R899 B.n221 B.n170 10.6151
R900 B.n225 B.n170 10.6151
R901 B.n226 B.n225 10.6151
R902 B.n227 B.n226 10.6151
R903 B.n227 B.n168 10.6151
R904 B.n231 B.n168 10.6151
R905 B.n232 B.n231 10.6151
R906 B.n233 B.n232 10.6151
R907 B.n233 B.n166 10.6151
R908 B.n237 B.n166 10.6151
R909 B.n238 B.n237 10.6151
R910 B.n239 B.n238 10.6151
R911 B.n239 B.n164 10.6151
R912 B.n243 B.n164 10.6151
R913 B.n244 B.n243 10.6151
R914 B.n245 B.n244 10.6151
R915 B.n245 B.n162 10.6151
R916 B.n249 B.n162 10.6151
R917 B.n250 B.n249 10.6151
R918 B.n251 B.n250 10.6151
R919 B.n251 B.n160 10.6151
R920 B.n255 B.n160 10.6151
R921 B.n256 B.n255 10.6151
R922 B.n257 B.n256 10.6151
R923 B.n257 B.n158 10.6151
R924 B.n261 B.n158 10.6151
R925 B.n262 B.n261 10.6151
R926 B.n263 B.n262 10.6151
R927 B.n263 B.n156 10.6151
R928 B.n267 B.n156 10.6151
R929 B.n268 B.n267 10.6151
R930 B.n269 B.n268 10.6151
R931 B.n269 B.n154 10.6151
R932 B.n273 B.n154 10.6151
R933 B.n274 B.n273 10.6151
R934 B.n275 B.n274 10.6151
R935 B.n275 B.n152 10.6151
R936 B.n279 B.n152 10.6151
R937 B.n280 B.n279 10.6151
R938 B.n281 B.n280 10.6151
R939 B.n281 B.n150 10.6151
R940 B.n285 B.n150 10.6151
R941 B.n286 B.n285 10.6151
R942 B.n287 B.n286 10.6151
R943 B.n287 B.n148 10.6151
R944 B.n291 B.n148 10.6151
R945 B.n292 B.n291 10.6151
R946 B.n293 B.n292 10.6151
R947 B.n293 B.n146 10.6151
R948 B.n297 B.n146 10.6151
R949 B.n298 B.n297 10.6151
R950 B.n299 B.n298 10.6151
R951 B.n299 B.n144 10.6151
R952 B.n303 B.n144 10.6151
R953 B.n304 B.n303 10.6151
R954 B.n306 B.n140 10.6151
R955 B.n310 B.n140 10.6151
R956 B.n311 B.n310 10.6151
R957 B.n312 B.n311 10.6151
R958 B.n312 B.n138 10.6151
R959 B.n316 B.n138 10.6151
R960 B.n317 B.n316 10.6151
R961 B.n318 B.n317 10.6151
R962 B.n322 B.n321 10.6151
R963 B.n323 B.n322 10.6151
R964 B.n323 B.n132 10.6151
R965 B.n327 B.n132 10.6151
R966 B.n328 B.n327 10.6151
R967 B.n329 B.n328 10.6151
R968 B.n329 B.n130 10.6151
R969 B.n333 B.n130 10.6151
R970 B.n334 B.n333 10.6151
R971 B.n335 B.n334 10.6151
R972 B.n335 B.n128 10.6151
R973 B.n339 B.n128 10.6151
R974 B.n340 B.n339 10.6151
R975 B.n341 B.n340 10.6151
R976 B.n341 B.n126 10.6151
R977 B.n345 B.n126 10.6151
R978 B.n346 B.n345 10.6151
R979 B.n347 B.n346 10.6151
R980 B.n347 B.n124 10.6151
R981 B.n351 B.n124 10.6151
R982 B.n352 B.n351 10.6151
R983 B.n353 B.n352 10.6151
R984 B.n353 B.n122 10.6151
R985 B.n357 B.n122 10.6151
R986 B.n358 B.n357 10.6151
R987 B.n359 B.n358 10.6151
R988 B.n359 B.n120 10.6151
R989 B.n363 B.n120 10.6151
R990 B.n364 B.n363 10.6151
R991 B.n365 B.n364 10.6151
R992 B.n365 B.n118 10.6151
R993 B.n369 B.n118 10.6151
R994 B.n370 B.n369 10.6151
R995 B.n371 B.n370 10.6151
R996 B.n371 B.n116 10.6151
R997 B.n375 B.n116 10.6151
R998 B.n376 B.n375 10.6151
R999 B.n377 B.n376 10.6151
R1000 B.n377 B.n114 10.6151
R1001 B.n381 B.n114 10.6151
R1002 B.n382 B.n381 10.6151
R1003 B.n383 B.n382 10.6151
R1004 B.n383 B.n112 10.6151
R1005 B.n387 B.n112 10.6151
R1006 B.n388 B.n387 10.6151
R1007 B.n389 B.n388 10.6151
R1008 B.n389 B.n110 10.6151
R1009 B.n393 B.n110 10.6151
R1010 B.n394 B.n393 10.6151
R1011 B.n395 B.n394 10.6151
R1012 B.n395 B.n108 10.6151
R1013 B.n399 B.n108 10.6151
R1014 B.n400 B.n399 10.6151
R1015 B.n401 B.n400 10.6151
R1016 B.n401 B.n106 10.6151
R1017 B.n405 B.n106 10.6151
R1018 B.n406 B.n405 10.6151
R1019 B.n407 B.n406 10.6151
R1020 B.n407 B.n104 10.6151
R1021 B.n411 B.n104 10.6151
R1022 B.n412 B.n411 10.6151
R1023 B.n413 B.n412 10.6151
R1024 B.n413 B.n102 10.6151
R1025 B.n208 B.n207 10.6151
R1026 B.n207 B.n176 10.6151
R1027 B.n203 B.n176 10.6151
R1028 B.n203 B.n202 10.6151
R1029 B.n202 B.n201 10.6151
R1030 B.n201 B.n178 10.6151
R1031 B.n197 B.n178 10.6151
R1032 B.n197 B.n196 10.6151
R1033 B.n196 B.n195 10.6151
R1034 B.n195 B.n180 10.6151
R1035 B.n191 B.n180 10.6151
R1036 B.n191 B.n190 10.6151
R1037 B.n190 B.n189 10.6151
R1038 B.n189 B.n182 10.6151
R1039 B.n185 B.n182 10.6151
R1040 B.n185 B.n184 10.6151
R1041 B.n184 B.n0 10.6151
R1042 B.n703 B.n1 10.6151
R1043 B.n703 B.n702 10.6151
R1044 B.n702 B.n701 10.6151
R1045 B.n701 B.n4 10.6151
R1046 B.n697 B.n4 10.6151
R1047 B.n697 B.n696 10.6151
R1048 B.n696 B.n695 10.6151
R1049 B.n695 B.n6 10.6151
R1050 B.n691 B.n6 10.6151
R1051 B.n691 B.n690 10.6151
R1052 B.n690 B.n689 10.6151
R1053 B.n689 B.n8 10.6151
R1054 B.n685 B.n8 10.6151
R1055 B.n685 B.n684 10.6151
R1056 B.n684 B.n683 10.6151
R1057 B.n683 B.n10 10.6151
R1058 B.n679 B.n10 10.6151
R1059 B.n582 B.n581 6.5566
R1060 B.n569 B.n568 6.5566
R1061 B.n306 B.n305 6.5566
R1062 B.n318 B.n136 6.5566
R1063 B.n583 B.n582 4.05904
R1064 B.n568 B.n567 4.05904
R1065 B.n305 B.n304 4.05904
R1066 B.n321 B.n136 4.05904
R1067 B.n707 B.n0 2.81026
R1068 B.n707 B.n1 2.81026
R1069 VN VN.t0 511.866
R1070 VN VN.t1 464.719
R1071 VTAIL.n353 VTAIL.n352 585
R1072 VTAIL.n350 VTAIL.n349 585
R1073 VTAIL.n359 VTAIL.n358 585
R1074 VTAIL.n361 VTAIL.n360 585
R1075 VTAIL.n346 VTAIL.n345 585
R1076 VTAIL.n367 VTAIL.n366 585
R1077 VTAIL.n370 VTAIL.n369 585
R1078 VTAIL.n368 VTAIL.n342 585
R1079 VTAIL.n375 VTAIL.n341 585
R1080 VTAIL.n377 VTAIL.n376 585
R1081 VTAIL.n379 VTAIL.n378 585
R1082 VTAIL.n338 VTAIL.n337 585
R1083 VTAIL.n385 VTAIL.n384 585
R1084 VTAIL.n387 VTAIL.n386 585
R1085 VTAIL.n334 VTAIL.n333 585
R1086 VTAIL.n393 VTAIL.n392 585
R1087 VTAIL.n395 VTAIL.n394 585
R1088 VTAIL.n330 VTAIL.n329 585
R1089 VTAIL.n401 VTAIL.n400 585
R1090 VTAIL.n403 VTAIL.n402 585
R1091 VTAIL.n326 VTAIL.n325 585
R1092 VTAIL.n409 VTAIL.n408 585
R1093 VTAIL.n411 VTAIL.n410 585
R1094 VTAIL.n322 VTAIL.n321 585
R1095 VTAIL.n417 VTAIL.n416 585
R1096 VTAIL.n419 VTAIL.n418 585
R1097 VTAIL.n35 VTAIL.n34 585
R1098 VTAIL.n32 VTAIL.n31 585
R1099 VTAIL.n41 VTAIL.n40 585
R1100 VTAIL.n43 VTAIL.n42 585
R1101 VTAIL.n28 VTAIL.n27 585
R1102 VTAIL.n49 VTAIL.n48 585
R1103 VTAIL.n52 VTAIL.n51 585
R1104 VTAIL.n50 VTAIL.n24 585
R1105 VTAIL.n57 VTAIL.n23 585
R1106 VTAIL.n59 VTAIL.n58 585
R1107 VTAIL.n61 VTAIL.n60 585
R1108 VTAIL.n20 VTAIL.n19 585
R1109 VTAIL.n67 VTAIL.n66 585
R1110 VTAIL.n69 VTAIL.n68 585
R1111 VTAIL.n16 VTAIL.n15 585
R1112 VTAIL.n75 VTAIL.n74 585
R1113 VTAIL.n77 VTAIL.n76 585
R1114 VTAIL.n12 VTAIL.n11 585
R1115 VTAIL.n83 VTAIL.n82 585
R1116 VTAIL.n85 VTAIL.n84 585
R1117 VTAIL.n8 VTAIL.n7 585
R1118 VTAIL.n91 VTAIL.n90 585
R1119 VTAIL.n93 VTAIL.n92 585
R1120 VTAIL.n4 VTAIL.n3 585
R1121 VTAIL.n99 VTAIL.n98 585
R1122 VTAIL.n101 VTAIL.n100 585
R1123 VTAIL.n313 VTAIL.n312 585
R1124 VTAIL.n311 VTAIL.n310 585
R1125 VTAIL.n216 VTAIL.n215 585
R1126 VTAIL.n305 VTAIL.n304 585
R1127 VTAIL.n303 VTAIL.n302 585
R1128 VTAIL.n220 VTAIL.n219 585
R1129 VTAIL.n297 VTAIL.n296 585
R1130 VTAIL.n295 VTAIL.n294 585
R1131 VTAIL.n224 VTAIL.n223 585
R1132 VTAIL.n289 VTAIL.n288 585
R1133 VTAIL.n287 VTAIL.n286 585
R1134 VTAIL.n228 VTAIL.n227 585
R1135 VTAIL.n281 VTAIL.n280 585
R1136 VTAIL.n279 VTAIL.n278 585
R1137 VTAIL.n232 VTAIL.n231 585
R1138 VTAIL.n273 VTAIL.n272 585
R1139 VTAIL.n271 VTAIL.n270 585
R1140 VTAIL.n269 VTAIL.n235 585
R1141 VTAIL.n239 VTAIL.n236 585
R1142 VTAIL.n264 VTAIL.n263 585
R1143 VTAIL.n262 VTAIL.n261 585
R1144 VTAIL.n241 VTAIL.n240 585
R1145 VTAIL.n256 VTAIL.n255 585
R1146 VTAIL.n254 VTAIL.n253 585
R1147 VTAIL.n245 VTAIL.n244 585
R1148 VTAIL.n248 VTAIL.n247 585
R1149 VTAIL.n207 VTAIL.n206 585
R1150 VTAIL.n205 VTAIL.n204 585
R1151 VTAIL.n110 VTAIL.n109 585
R1152 VTAIL.n199 VTAIL.n198 585
R1153 VTAIL.n197 VTAIL.n196 585
R1154 VTAIL.n114 VTAIL.n113 585
R1155 VTAIL.n191 VTAIL.n190 585
R1156 VTAIL.n189 VTAIL.n188 585
R1157 VTAIL.n118 VTAIL.n117 585
R1158 VTAIL.n183 VTAIL.n182 585
R1159 VTAIL.n181 VTAIL.n180 585
R1160 VTAIL.n122 VTAIL.n121 585
R1161 VTAIL.n175 VTAIL.n174 585
R1162 VTAIL.n173 VTAIL.n172 585
R1163 VTAIL.n126 VTAIL.n125 585
R1164 VTAIL.n167 VTAIL.n166 585
R1165 VTAIL.n165 VTAIL.n164 585
R1166 VTAIL.n163 VTAIL.n129 585
R1167 VTAIL.n133 VTAIL.n130 585
R1168 VTAIL.n158 VTAIL.n157 585
R1169 VTAIL.n156 VTAIL.n155 585
R1170 VTAIL.n135 VTAIL.n134 585
R1171 VTAIL.n150 VTAIL.n149 585
R1172 VTAIL.n148 VTAIL.n147 585
R1173 VTAIL.n139 VTAIL.n138 585
R1174 VTAIL.n142 VTAIL.n141 585
R1175 VTAIL.n418 VTAIL.n318 498.474
R1176 VTAIL.n100 VTAIL.n0 498.474
R1177 VTAIL.n312 VTAIL.n212 498.474
R1178 VTAIL.n206 VTAIL.n106 498.474
R1179 VTAIL.t3 VTAIL.n351 329.036
R1180 VTAIL.t1 VTAIL.n33 329.036
R1181 VTAIL.t0 VTAIL.n246 329.036
R1182 VTAIL.t2 VTAIL.n140 329.036
R1183 VTAIL.n352 VTAIL.n349 171.744
R1184 VTAIL.n359 VTAIL.n349 171.744
R1185 VTAIL.n360 VTAIL.n359 171.744
R1186 VTAIL.n360 VTAIL.n345 171.744
R1187 VTAIL.n367 VTAIL.n345 171.744
R1188 VTAIL.n369 VTAIL.n367 171.744
R1189 VTAIL.n369 VTAIL.n368 171.744
R1190 VTAIL.n368 VTAIL.n341 171.744
R1191 VTAIL.n377 VTAIL.n341 171.744
R1192 VTAIL.n378 VTAIL.n377 171.744
R1193 VTAIL.n378 VTAIL.n337 171.744
R1194 VTAIL.n385 VTAIL.n337 171.744
R1195 VTAIL.n386 VTAIL.n385 171.744
R1196 VTAIL.n386 VTAIL.n333 171.744
R1197 VTAIL.n393 VTAIL.n333 171.744
R1198 VTAIL.n394 VTAIL.n393 171.744
R1199 VTAIL.n394 VTAIL.n329 171.744
R1200 VTAIL.n401 VTAIL.n329 171.744
R1201 VTAIL.n402 VTAIL.n401 171.744
R1202 VTAIL.n402 VTAIL.n325 171.744
R1203 VTAIL.n409 VTAIL.n325 171.744
R1204 VTAIL.n410 VTAIL.n409 171.744
R1205 VTAIL.n410 VTAIL.n321 171.744
R1206 VTAIL.n417 VTAIL.n321 171.744
R1207 VTAIL.n418 VTAIL.n417 171.744
R1208 VTAIL.n34 VTAIL.n31 171.744
R1209 VTAIL.n41 VTAIL.n31 171.744
R1210 VTAIL.n42 VTAIL.n41 171.744
R1211 VTAIL.n42 VTAIL.n27 171.744
R1212 VTAIL.n49 VTAIL.n27 171.744
R1213 VTAIL.n51 VTAIL.n49 171.744
R1214 VTAIL.n51 VTAIL.n50 171.744
R1215 VTAIL.n50 VTAIL.n23 171.744
R1216 VTAIL.n59 VTAIL.n23 171.744
R1217 VTAIL.n60 VTAIL.n59 171.744
R1218 VTAIL.n60 VTAIL.n19 171.744
R1219 VTAIL.n67 VTAIL.n19 171.744
R1220 VTAIL.n68 VTAIL.n67 171.744
R1221 VTAIL.n68 VTAIL.n15 171.744
R1222 VTAIL.n75 VTAIL.n15 171.744
R1223 VTAIL.n76 VTAIL.n75 171.744
R1224 VTAIL.n76 VTAIL.n11 171.744
R1225 VTAIL.n83 VTAIL.n11 171.744
R1226 VTAIL.n84 VTAIL.n83 171.744
R1227 VTAIL.n84 VTAIL.n7 171.744
R1228 VTAIL.n91 VTAIL.n7 171.744
R1229 VTAIL.n92 VTAIL.n91 171.744
R1230 VTAIL.n92 VTAIL.n3 171.744
R1231 VTAIL.n99 VTAIL.n3 171.744
R1232 VTAIL.n100 VTAIL.n99 171.744
R1233 VTAIL.n312 VTAIL.n311 171.744
R1234 VTAIL.n311 VTAIL.n215 171.744
R1235 VTAIL.n304 VTAIL.n215 171.744
R1236 VTAIL.n304 VTAIL.n303 171.744
R1237 VTAIL.n303 VTAIL.n219 171.744
R1238 VTAIL.n296 VTAIL.n219 171.744
R1239 VTAIL.n296 VTAIL.n295 171.744
R1240 VTAIL.n295 VTAIL.n223 171.744
R1241 VTAIL.n288 VTAIL.n223 171.744
R1242 VTAIL.n288 VTAIL.n287 171.744
R1243 VTAIL.n287 VTAIL.n227 171.744
R1244 VTAIL.n280 VTAIL.n227 171.744
R1245 VTAIL.n280 VTAIL.n279 171.744
R1246 VTAIL.n279 VTAIL.n231 171.744
R1247 VTAIL.n272 VTAIL.n231 171.744
R1248 VTAIL.n272 VTAIL.n271 171.744
R1249 VTAIL.n271 VTAIL.n235 171.744
R1250 VTAIL.n239 VTAIL.n235 171.744
R1251 VTAIL.n263 VTAIL.n239 171.744
R1252 VTAIL.n263 VTAIL.n262 171.744
R1253 VTAIL.n262 VTAIL.n240 171.744
R1254 VTAIL.n255 VTAIL.n240 171.744
R1255 VTAIL.n255 VTAIL.n254 171.744
R1256 VTAIL.n254 VTAIL.n244 171.744
R1257 VTAIL.n247 VTAIL.n244 171.744
R1258 VTAIL.n206 VTAIL.n205 171.744
R1259 VTAIL.n205 VTAIL.n109 171.744
R1260 VTAIL.n198 VTAIL.n109 171.744
R1261 VTAIL.n198 VTAIL.n197 171.744
R1262 VTAIL.n197 VTAIL.n113 171.744
R1263 VTAIL.n190 VTAIL.n113 171.744
R1264 VTAIL.n190 VTAIL.n189 171.744
R1265 VTAIL.n189 VTAIL.n117 171.744
R1266 VTAIL.n182 VTAIL.n117 171.744
R1267 VTAIL.n182 VTAIL.n181 171.744
R1268 VTAIL.n181 VTAIL.n121 171.744
R1269 VTAIL.n174 VTAIL.n121 171.744
R1270 VTAIL.n174 VTAIL.n173 171.744
R1271 VTAIL.n173 VTAIL.n125 171.744
R1272 VTAIL.n166 VTAIL.n125 171.744
R1273 VTAIL.n166 VTAIL.n165 171.744
R1274 VTAIL.n165 VTAIL.n129 171.744
R1275 VTAIL.n133 VTAIL.n129 171.744
R1276 VTAIL.n157 VTAIL.n133 171.744
R1277 VTAIL.n157 VTAIL.n156 171.744
R1278 VTAIL.n156 VTAIL.n134 171.744
R1279 VTAIL.n149 VTAIL.n134 171.744
R1280 VTAIL.n149 VTAIL.n148 171.744
R1281 VTAIL.n148 VTAIL.n138 171.744
R1282 VTAIL.n141 VTAIL.n138 171.744
R1283 VTAIL.n352 VTAIL.t3 85.8723
R1284 VTAIL.n34 VTAIL.t1 85.8723
R1285 VTAIL.n247 VTAIL.t0 85.8723
R1286 VTAIL.n141 VTAIL.t2 85.8723
R1287 VTAIL.n423 VTAIL.n422 36.646
R1288 VTAIL.n105 VTAIL.n104 36.646
R1289 VTAIL.n317 VTAIL.n316 36.646
R1290 VTAIL.n211 VTAIL.n210 36.646
R1291 VTAIL.n211 VTAIL.n105 32.0824
R1292 VTAIL.n423 VTAIL.n317 30.6514
R1293 VTAIL.n376 VTAIL.n375 13.1884
R1294 VTAIL.n58 VTAIL.n57 13.1884
R1295 VTAIL.n270 VTAIL.n269 13.1884
R1296 VTAIL.n164 VTAIL.n163 13.1884
R1297 VTAIL.n374 VTAIL.n342 12.8005
R1298 VTAIL.n379 VTAIL.n340 12.8005
R1299 VTAIL.n420 VTAIL.n419 12.8005
R1300 VTAIL.n56 VTAIL.n24 12.8005
R1301 VTAIL.n61 VTAIL.n22 12.8005
R1302 VTAIL.n102 VTAIL.n101 12.8005
R1303 VTAIL.n314 VTAIL.n313 12.8005
R1304 VTAIL.n273 VTAIL.n234 12.8005
R1305 VTAIL.n268 VTAIL.n236 12.8005
R1306 VTAIL.n208 VTAIL.n207 12.8005
R1307 VTAIL.n167 VTAIL.n128 12.8005
R1308 VTAIL.n162 VTAIL.n130 12.8005
R1309 VTAIL.n371 VTAIL.n370 12.0247
R1310 VTAIL.n380 VTAIL.n338 12.0247
R1311 VTAIL.n416 VTAIL.n320 12.0247
R1312 VTAIL.n53 VTAIL.n52 12.0247
R1313 VTAIL.n62 VTAIL.n20 12.0247
R1314 VTAIL.n98 VTAIL.n2 12.0247
R1315 VTAIL.n310 VTAIL.n214 12.0247
R1316 VTAIL.n274 VTAIL.n232 12.0247
R1317 VTAIL.n265 VTAIL.n264 12.0247
R1318 VTAIL.n204 VTAIL.n108 12.0247
R1319 VTAIL.n168 VTAIL.n126 12.0247
R1320 VTAIL.n159 VTAIL.n158 12.0247
R1321 VTAIL.n366 VTAIL.n344 11.249
R1322 VTAIL.n384 VTAIL.n383 11.249
R1323 VTAIL.n415 VTAIL.n322 11.249
R1324 VTAIL.n48 VTAIL.n26 11.249
R1325 VTAIL.n66 VTAIL.n65 11.249
R1326 VTAIL.n97 VTAIL.n4 11.249
R1327 VTAIL.n309 VTAIL.n216 11.249
R1328 VTAIL.n278 VTAIL.n277 11.249
R1329 VTAIL.n261 VTAIL.n238 11.249
R1330 VTAIL.n203 VTAIL.n110 11.249
R1331 VTAIL.n172 VTAIL.n171 11.249
R1332 VTAIL.n155 VTAIL.n132 11.249
R1333 VTAIL.n353 VTAIL.n351 10.7239
R1334 VTAIL.n35 VTAIL.n33 10.7239
R1335 VTAIL.n248 VTAIL.n246 10.7239
R1336 VTAIL.n142 VTAIL.n140 10.7239
R1337 VTAIL.n365 VTAIL.n346 10.4732
R1338 VTAIL.n387 VTAIL.n336 10.4732
R1339 VTAIL.n412 VTAIL.n411 10.4732
R1340 VTAIL.n47 VTAIL.n28 10.4732
R1341 VTAIL.n69 VTAIL.n18 10.4732
R1342 VTAIL.n94 VTAIL.n93 10.4732
R1343 VTAIL.n306 VTAIL.n305 10.4732
R1344 VTAIL.n281 VTAIL.n230 10.4732
R1345 VTAIL.n260 VTAIL.n241 10.4732
R1346 VTAIL.n200 VTAIL.n199 10.4732
R1347 VTAIL.n175 VTAIL.n124 10.4732
R1348 VTAIL.n154 VTAIL.n135 10.4732
R1349 VTAIL.n362 VTAIL.n361 9.69747
R1350 VTAIL.n388 VTAIL.n334 9.69747
R1351 VTAIL.n408 VTAIL.n324 9.69747
R1352 VTAIL.n44 VTAIL.n43 9.69747
R1353 VTAIL.n70 VTAIL.n16 9.69747
R1354 VTAIL.n90 VTAIL.n6 9.69747
R1355 VTAIL.n302 VTAIL.n218 9.69747
R1356 VTAIL.n282 VTAIL.n228 9.69747
R1357 VTAIL.n257 VTAIL.n256 9.69747
R1358 VTAIL.n196 VTAIL.n112 9.69747
R1359 VTAIL.n176 VTAIL.n122 9.69747
R1360 VTAIL.n151 VTAIL.n150 9.69747
R1361 VTAIL.n422 VTAIL.n421 9.45567
R1362 VTAIL.n104 VTAIL.n103 9.45567
R1363 VTAIL.n316 VTAIL.n315 9.45567
R1364 VTAIL.n210 VTAIL.n209 9.45567
R1365 VTAIL.n397 VTAIL.n396 9.3005
R1366 VTAIL.n332 VTAIL.n331 9.3005
R1367 VTAIL.n391 VTAIL.n390 9.3005
R1368 VTAIL.n389 VTAIL.n388 9.3005
R1369 VTAIL.n336 VTAIL.n335 9.3005
R1370 VTAIL.n383 VTAIL.n382 9.3005
R1371 VTAIL.n381 VTAIL.n380 9.3005
R1372 VTAIL.n340 VTAIL.n339 9.3005
R1373 VTAIL.n355 VTAIL.n354 9.3005
R1374 VTAIL.n357 VTAIL.n356 9.3005
R1375 VTAIL.n348 VTAIL.n347 9.3005
R1376 VTAIL.n363 VTAIL.n362 9.3005
R1377 VTAIL.n365 VTAIL.n364 9.3005
R1378 VTAIL.n344 VTAIL.n343 9.3005
R1379 VTAIL.n372 VTAIL.n371 9.3005
R1380 VTAIL.n374 VTAIL.n373 9.3005
R1381 VTAIL.n399 VTAIL.n398 9.3005
R1382 VTAIL.n328 VTAIL.n327 9.3005
R1383 VTAIL.n405 VTAIL.n404 9.3005
R1384 VTAIL.n407 VTAIL.n406 9.3005
R1385 VTAIL.n324 VTAIL.n323 9.3005
R1386 VTAIL.n413 VTAIL.n412 9.3005
R1387 VTAIL.n415 VTAIL.n414 9.3005
R1388 VTAIL.n320 VTAIL.n319 9.3005
R1389 VTAIL.n421 VTAIL.n420 9.3005
R1390 VTAIL.n79 VTAIL.n78 9.3005
R1391 VTAIL.n14 VTAIL.n13 9.3005
R1392 VTAIL.n73 VTAIL.n72 9.3005
R1393 VTAIL.n71 VTAIL.n70 9.3005
R1394 VTAIL.n18 VTAIL.n17 9.3005
R1395 VTAIL.n65 VTAIL.n64 9.3005
R1396 VTAIL.n63 VTAIL.n62 9.3005
R1397 VTAIL.n22 VTAIL.n21 9.3005
R1398 VTAIL.n37 VTAIL.n36 9.3005
R1399 VTAIL.n39 VTAIL.n38 9.3005
R1400 VTAIL.n30 VTAIL.n29 9.3005
R1401 VTAIL.n45 VTAIL.n44 9.3005
R1402 VTAIL.n47 VTAIL.n46 9.3005
R1403 VTAIL.n26 VTAIL.n25 9.3005
R1404 VTAIL.n54 VTAIL.n53 9.3005
R1405 VTAIL.n56 VTAIL.n55 9.3005
R1406 VTAIL.n81 VTAIL.n80 9.3005
R1407 VTAIL.n10 VTAIL.n9 9.3005
R1408 VTAIL.n87 VTAIL.n86 9.3005
R1409 VTAIL.n89 VTAIL.n88 9.3005
R1410 VTAIL.n6 VTAIL.n5 9.3005
R1411 VTAIL.n95 VTAIL.n94 9.3005
R1412 VTAIL.n97 VTAIL.n96 9.3005
R1413 VTAIL.n2 VTAIL.n1 9.3005
R1414 VTAIL.n103 VTAIL.n102 9.3005
R1415 VTAIL.n250 VTAIL.n249 9.3005
R1416 VTAIL.n252 VTAIL.n251 9.3005
R1417 VTAIL.n243 VTAIL.n242 9.3005
R1418 VTAIL.n258 VTAIL.n257 9.3005
R1419 VTAIL.n260 VTAIL.n259 9.3005
R1420 VTAIL.n238 VTAIL.n237 9.3005
R1421 VTAIL.n266 VTAIL.n265 9.3005
R1422 VTAIL.n268 VTAIL.n267 9.3005
R1423 VTAIL.n222 VTAIL.n221 9.3005
R1424 VTAIL.n299 VTAIL.n298 9.3005
R1425 VTAIL.n301 VTAIL.n300 9.3005
R1426 VTAIL.n218 VTAIL.n217 9.3005
R1427 VTAIL.n307 VTAIL.n306 9.3005
R1428 VTAIL.n309 VTAIL.n308 9.3005
R1429 VTAIL.n214 VTAIL.n213 9.3005
R1430 VTAIL.n315 VTAIL.n314 9.3005
R1431 VTAIL.n293 VTAIL.n292 9.3005
R1432 VTAIL.n291 VTAIL.n290 9.3005
R1433 VTAIL.n226 VTAIL.n225 9.3005
R1434 VTAIL.n285 VTAIL.n284 9.3005
R1435 VTAIL.n283 VTAIL.n282 9.3005
R1436 VTAIL.n230 VTAIL.n229 9.3005
R1437 VTAIL.n277 VTAIL.n276 9.3005
R1438 VTAIL.n275 VTAIL.n274 9.3005
R1439 VTAIL.n234 VTAIL.n233 9.3005
R1440 VTAIL.n144 VTAIL.n143 9.3005
R1441 VTAIL.n146 VTAIL.n145 9.3005
R1442 VTAIL.n137 VTAIL.n136 9.3005
R1443 VTAIL.n152 VTAIL.n151 9.3005
R1444 VTAIL.n154 VTAIL.n153 9.3005
R1445 VTAIL.n132 VTAIL.n131 9.3005
R1446 VTAIL.n160 VTAIL.n159 9.3005
R1447 VTAIL.n162 VTAIL.n161 9.3005
R1448 VTAIL.n116 VTAIL.n115 9.3005
R1449 VTAIL.n193 VTAIL.n192 9.3005
R1450 VTAIL.n195 VTAIL.n194 9.3005
R1451 VTAIL.n112 VTAIL.n111 9.3005
R1452 VTAIL.n201 VTAIL.n200 9.3005
R1453 VTAIL.n203 VTAIL.n202 9.3005
R1454 VTAIL.n108 VTAIL.n107 9.3005
R1455 VTAIL.n209 VTAIL.n208 9.3005
R1456 VTAIL.n187 VTAIL.n186 9.3005
R1457 VTAIL.n185 VTAIL.n184 9.3005
R1458 VTAIL.n120 VTAIL.n119 9.3005
R1459 VTAIL.n179 VTAIL.n178 9.3005
R1460 VTAIL.n177 VTAIL.n176 9.3005
R1461 VTAIL.n124 VTAIL.n123 9.3005
R1462 VTAIL.n171 VTAIL.n170 9.3005
R1463 VTAIL.n169 VTAIL.n168 9.3005
R1464 VTAIL.n128 VTAIL.n127 9.3005
R1465 VTAIL.n358 VTAIL.n348 8.92171
R1466 VTAIL.n392 VTAIL.n391 8.92171
R1467 VTAIL.n407 VTAIL.n326 8.92171
R1468 VTAIL.n40 VTAIL.n30 8.92171
R1469 VTAIL.n74 VTAIL.n73 8.92171
R1470 VTAIL.n89 VTAIL.n8 8.92171
R1471 VTAIL.n301 VTAIL.n220 8.92171
R1472 VTAIL.n286 VTAIL.n285 8.92171
R1473 VTAIL.n253 VTAIL.n243 8.92171
R1474 VTAIL.n195 VTAIL.n114 8.92171
R1475 VTAIL.n180 VTAIL.n179 8.92171
R1476 VTAIL.n147 VTAIL.n137 8.92171
R1477 VTAIL.n357 VTAIL.n350 8.14595
R1478 VTAIL.n395 VTAIL.n332 8.14595
R1479 VTAIL.n404 VTAIL.n403 8.14595
R1480 VTAIL.n39 VTAIL.n32 8.14595
R1481 VTAIL.n77 VTAIL.n14 8.14595
R1482 VTAIL.n86 VTAIL.n85 8.14595
R1483 VTAIL.n298 VTAIL.n297 8.14595
R1484 VTAIL.n289 VTAIL.n226 8.14595
R1485 VTAIL.n252 VTAIL.n245 8.14595
R1486 VTAIL.n192 VTAIL.n191 8.14595
R1487 VTAIL.n183 VTAIL.n120 8.14595
R1488 VTAIL.n146 VTAIL.n139 8.14595
R1489 VTAIL.n422 VTAIL.n318 7.75445
R1490 VTAIL.n104 VTAIL.n0 7.75445
R1491 VTAIL.n316 VTAIL.n212 7.75445
R1492 VTAIL.n210 VTAIL.n106 7.75445
R1493 VTAIL.n354 VTAIL.n353 7.3702
R1494 VTAIL.n396 VTAIL.n330 7.3702
R1495 VTAIL.n400 VTAIL.n328 7.3702
R1496 VTAIL.n36 VTAIL.n35 7.3702
R1497 VTAIL.n78 VTAIL.n12 7.3702
R1498 VTAIL.n82 VTAIL.n10 7.3702
R1499 VTAIL.n294 VTAIL.n222 7.3702
R1500 VTAIL.n290 VTAIL.n224 7.3702
R1501 VTAIL.n249 VTAIL.n248 7.3702
R1502 VTAIL.n188 VTAIL.n116 7.3702
R1503 VTAIL.n184 VTAIL.n118 7.3702
R1504 VTAIL.n143 VTAIL.n142 7.3702
R1505 VTAIL.n399 VTAIL.n330 6.59444
R1506 VTAIL.n400 VTAIL.n399 6.59444
R1507 VTAIL.n81 VTAIL.n12 6.59444
R1508 VTAIL.n82 VTAIL.n81 6.59444
R1509 VTAIL.n294 VTAIL.n293 6.59444
R1510 VTAIL.n293 VTAIL.n224 6.59444
R1511 VTAIL.n188 VTAIL.n187 6.59444
R1512 VTAIL.n187 VTAIL.n118 6.59444
R1513 VTAIL.n420 VTAIL.n318 6.08283
R1514 VTAIL.n102 VTAIL.n0 6.08283
R1515 VTAIL.n314 VTAIL.n212 6.08283
R1516 VTAIL.n208 VTAIL.n106 6.08283
R1517 VTAIL.n354 VTAIL.n350 5.81868
R1518 VTAIL.n396 VTAIL.n395 5.81868
R1519 VTAIL.n403 VTAIL.n328 5.81868
R1520 VTAIL.n36 VTAIL.n32 5.81868
R1521 VTAIL.n78 VTAIL.n77 5.81868
R1522 VTAIL.n85 VTAIL.n10 5.81868
R1523 VTAIL.n297 VTAIL.n222 5.81868
R1524 VTAIL.n290 VTAIL.n289 5.81868
R1525 VTAIL.n249 VTAIL.n245 5.81868
R1526 VTAIL.n191 VTAIL.n116 5.81868
R1527 VTAIL.n184 VTAIL.n183 5.81868
R1528 VTAIL.n143 VTAIL.n139 5.81868
R1529 VTAIL.n358 VTAIL.n357 5.04292
R1530 VTAIL.n392 VTAIL.n332 5.04292
R1531 VTAIL.n404 VTAIL.n326 5.04292
R1532 VTAIL.n40 VTAIL.n39 5.04292
R1533 VTAIL.n74 VTAIL.n14 5.04292
R1534 VTAIL.n86 VTAIL.n8 5.04292
R1535 VTAIL.n298 VTAIL.n220 5.04292
R1536 VTAIL.n286 VTAIL.n226 5.04292
R1537 VTAIL.n253 VTAIL.n252 5.04292
R1538 VTAIL.n192 VTAIL.n114 5.04292
R1539 VTAIL.n180 VTAIL.n120 5.04292
R1540 VTAIL.n147 VTAIL.n146 5.04292
R1541 VTAIL.n361 VTAIL.n348 4.26717
R1542 VTAIL.n391 VTAIL.n334 4.26717
R1543 VTAIL.n408 VTAIL.n407 4.26717
R1544 VTAIL.n43 VTAIL.n30 4.26717
R1545 VTAIL.n73 VTAIL.n16 4.26717
R1546 VTAIL.n90 VTAIL.n89 4.26717
R1547 VTAIL.n302 VTAIL.n301 4.26717
R1548 VTAIL.n285 VTAIL.n228 4.26717
R1549 VTAIL.n256 VTAIL.n243 4.26717
R1550 VTAIL.n196 VTAIL.n195 4.26717
R1551 VTAIL.n179 VTAIL.n122 4.26717
R1552 VTAIL.n150 VTAIL.n137 4.26717
R1553 VTAIL.n362 VTAIL.n346 3.49141
R1554 VTAIL.n388 VTAIL.n387 3.49141
R1555 VTAIL.n411 VTAIL.n324 3.49141
R1556 VTAIL.n44 VTAIL.n28 3.49141
R1557 VTAIL.n70 VTAIL.n69 3.49141
R1558 VTAIL.n93 VTAIL.n6 3.49141
R1559 VTAIL.n305 VTAIL.n218 3.49141
R1560 VTAIL.n282 VTAIL.n281 3.49141
R1561 VTAIL.n257 VTAIL.n241 3.49141
R1562 VTAIL.n199 VTAIL.n112 3.49141
R1563 VTAIL.n176 VTAIL.n175 3.49141
R1564 VTAIL.n151 VTAIL.n135 3.49141
R1565 VTAIL.n366 VTAIL.n365 2.71565
R1566 VTAIL.n384 VTAIL.n336 2.71565
R1567 VTAIL.n412 VTAIL.n322 2.71565
R1568 VTAIL.n48 VTAIL.n47 2.71565
R1569 VTAIL.n66 VTAIL.n18 2.71565
R1570 VTAIL.n94 VTAIL.n4 2.71565
R1571 VTAIL.n306 VTAIL.n216 2.71565
R1572 VTAIL.n278 VTAIL.n230 2.71565
R1573 VTAIL.n261 VTAIL.n260 2.71565
R1574 VTAIL.n200 VTAIL.n110 2.71565
R1575 VTAIL.n172 VTAIL.n124 2.71565
R1576 VTAIL.n155 VTAIL.n154 2.71565
R1577 VTAIL.n250 VTAIL.n246 2.41282
R1578 VTAIL.n144 VTAIL.n140 2.41282
R1579 VTAIL.n355 VTAIL.n351 2.41282
R1580 VTAIL.n37 VTAIL.n33 2.41282
R1581 VTAIL.n370 VTAIL.n344 1.93989
R1582 VTAIL.n383 VTAIL.n338 1.93989
R1583 VTAIL.n416 VTAIL.n415 1.93989
R1584 VTAIL.n52 VTAIL.n26 1.93989
R1585 VTAIL.n65 VTAIL.n20 1.93989
R1586 VTAIL.n98 VTAIL.n97 1.93989
R1587 VTAIL.n310 VTAIL.n309 1.93989
R1588 VTAIL.n277 VTAIL.n232 1.93989
R1589 VTAIL.n264 VTAIL.n238 1.93989
R1590 VTAIL.n204 VTAIL.n203 1.93989
R1591 VTAIL.n171 VTAIL.n126 1.93989
R1592 VTAIL.n158 VTAIL.n132 1.93989
R1593 VTAIL.n317 VTAIL.n211 1.18584
R1594 VTAIL.n371 VTAIL.n342 1.16414
R1595 VTAIL.n380 VTAIL.n379 1.16414
R1596 VTAIL.n419 VTAIL.n320 1.16414
R1597 VTAIL.n53 VTAIL.n24 1.16414
R1598 VTAIL.n62 VTAIL.n61 1.16414
R1599 VTAIL.n101 VTAIL.n2 1.16414
R1600 VTAIL.n313 VTAIL.n214 1.16414
R1601 VTAIL.n274 VTAIL.n273 1.16414
R1602 VTAIL.n265 VTAIL.n236 1.16414
R1603 VTAIL.n207 VTAIL.n108 1.16414
R1604 VTAIL.n168 VTAIL.n167 1.16414
R1605 VTAIL.n159 VTAIL.n130 1.16414
R1606 VTAIL VTAIL.n105 0.886276
R1607 VTAIL.n375 VTAIL.n374 0.388379
R1608 VTAIL.n376 VTAIL.n340 0.388379
R1609 VTAIL.n57 VTAIL.n56 0.388379
R1610 VTAIL.n58 VTAIL.n22 0.388379
R1611 VTAIL.n270 VTAIL.n234 0.388379
R1612 VTAIL.n269 VTAIL.n268 0.388379
R1613 VTAIL.n164 VTAIL.n128 0.388379
R1614 VTAIL.n163 VTAIL.n162 0.388379
R1615 VTAIL VTAIL.n423 0.300069
R1616 VTAIL.n356 VTAIL.n355 0.155672
R1617 VTAIL.n356 VTAIL.n347 0.155672
R1618 VTAIL.n363 VTAIL.n347 0.155672
R1619 VTAIL.n364 VTAIL.n363 0.155672
R1620 VTAIL.n364 VTAIL.n343 0.155672
R1621 VTAIL.n372 VTAIL.n343 0.155672
R1622 VTAIL.n373 VTAIL.n372 0.155672
R1623 VTAIL.n373 VTAIL.n339 0.155672
R1624 VTAIL.n381 VTAIL.n339 0.155672
R1625 VTAIL.n382 VTAIL.n381 0.155672
R1626 VTAIL.n382 VTAIL.n335 0.155672
R1627 VTAIL.n389 VTAIL.n335 0.155672
R1628 VTAIL.n390 VTAIL.n389 0.155672
R1629 VTAIL.n390 VTAIL.n331 0.155672
R1630 VTAIL.n397 VTAIL.n331 0.155672
R1631 VTAIL.n398 VTAIL.n397 0.155672
R1632 VTAIL.n398 VTAIL.n327 0.155672
R1633 VTAIL.n405 VTAIL.n327 0.155672
R1634 VTAIL.n406 VTAIL.n405 0.155672
R1635 VTAIL.n406 VTAIL.n323 0.155672
R1636 VTAIL.n413 VTAIL.n323 0.155672
R1637 VTAIL.n414 VTAIL.n413 0.155672
R1638 VTAIL.n414 VTAIL.n319 0.155672
R1639 VTAIL.n421 VTAIL.n319 0.155672
R1640 VTAIL.n38 VTAIL.n37 0.155672
R1641 VTAIL.n38 VTAIL.n29 0.155672
R1642 VTAIL.n45 VTAIL.n29 0.155672
R1643 VTAIL.n46 VTAIL.n45 0.155672
R1644 VTAIL.n46 VTAIL.n25 0.155672
R1645 VTAIL.n54 VTAIL.n25 0.155672
R1646 VTAIL.n55 VTAIL.n54 0.155672
R1647 VTAIL.n55 VTAIL.n21 0.155672
R1648 VTAIL.n63 VTAIL.n21 0.155672
R1649 VTAIL.n64 VTAIL.n63 0.155672
R1650 VTAIL.n64 VTAIL.n17 0.155672
R1651 VTAIL.n71 VTAIL.n17 0.155672
R1652 VTAIL.n72 VTAIL.n71 0.155672
R1653 VTAIL.n72 VTAIL.n13 0.155672
R1654 VTAIL.n79 VTAIL.n13 0.155672
R1655 VTAIL.n80 VTAIL.n79 0.155672
R1656 VTAIL.n80 VTAIL.n9 0.155672
R1657 VTAIL.n87 VTAIL.n9 0.155672
R1658 VTAIL.n88 VTAIL.n87 0.155672
R1659 VTAIL.n88 VTAIL.n5 0.155672
R1660 VTAIL.n95 VTAIL.n5 0.155672
R1661 VTAIL.n96 VTAIL.n95 0.155672
R1662 VTAIL.n96 VTAIL.n1 0.155672
R1663 VTAIL.n103 VTAIL.n1 0.155672
R1664 VTAIL.n315 VTAIL.n213 0.155672
R1665 VTAIL.n308 VTAIL.n213 0.155672
R1666 VTAIL.n308 VTAIL.n307 0.155672
R1667 VTAIL.n307 VTAIL.n217 0.155672
R1668 VTAIL.n300 VTAIL.n217 0.155672
R1669 VTAIL.n300 VTAIL.n299 0.155672
R1670 VTAIL.n299 VTAIL.n221 0.155672
R1671 VTAIL.n292 VTAIL.n221 0.155672
R1672 VTAIL.n292 VTAIL.n291 0.155672
R1673 VTAIL.n291 VTAIL.n225 0.155672
R1674 VTAIL.n284 VTAIL.n225 0.155672
R1675 VTAIL.n284 VTAIL.n283 0.155672
R1676 VTAIL.n283 VTAIL.n229 0.155672
R1677 VTAIL.n276 VTAIL.n229 0.155672
R1678 VTAIL.n276 VTAIL.n275 0.155672
R1679 VTAIL.n275 VTAIL.n233 0.155672
R1680 VTAIL.n267 VTAIL.n233 0.155672
R1681 VTAIL.n267 VTAIL.n266 0.155672
R1682 VTAIL.n266 VTAIL.n237 0.155672
R1683 VTAIL.n259 VTAIL.n237 0.155672
R1684 VTAIL.n259 VTAIL.n258 0.155672
R1685 VTAIL.n258 VTAIL.n242 0.155672
R1686 VTAIL.n251 VTAIL.n242 0.155672
R1687 VTAIL.n251 VTAIL.n250 0.155672
R1688 VTAIL.n209 VTAIL.n107 0.155672
R1689 VTAIL.n202 VTAIL.n107 0.155672
R1690 VTAIL.n202 VTAIL.n201 0.155672
R1691 VTAIL.n201 VTAIL.n111 0.155672
R1692 VTAIL.n194 VTAIL.n111 0.155672
R1693 VTAIL.n194 VTAIL.n193 0.155672
R1694 VTAIL.n193 VTAIL.n115 0.155672
R1695 VTAIL.n186 VTAIL.n115 0.155672
R1696 VTAIL.n186 VTAIL.n185 0.155672
R1697 VTAIL.n185 VTAIL.n119 0.155672
R1698 VTAIL.n178 VTAIL.n119 0.155672
R1699 VTAIL.n178 VTAIL.n177 0.155672
R1700 VTAIL.n177 VTAIL.n123 0.155672
R1701 VTAIL.n170 VTAIL.n123 0.155672
R1702 VTAIL.n170 VTAIL.n169 0.155672
R1703 VTAIL.n169 VTAIL.n127 0.155672
R1704 VTAIL.n161 VTAIL.n127 0.155672
R1705 VTAIL.n161 VTAIL.n160 0.155672
R1706 VTAIL.n160 VTAIL.n131 0.155672
R1707 VTAIL.n153 VTAIL.n131 0.155672
R1708 VTAIL.n153 VTAIL.n152 0.155672
R1709 VTAIL.n152 VTAIL.n136 0.155672
R1710 VTAIL.n145 VTAIL.n136 0.155672
R1711 VTAIL.n145 VTAIL.n144 0.155672
R1712 VDD2.n206 VDD2.n205 585
R1713 VDD2.n204 VDD2.n203 585
R1714 VDD2.n109 VDD2.n108 585
R1715 VDD2.n198 VDD2.n197 585
R1716 VDD2.n196 VDD2.n195 585
R1717 VDD2.n113 VDD2.n112 585
R1718 VDD2.n190 VDD2.n189 585
R1719 VDD2.n188 VDD2.n187 585
R1720 VDD2.n117 VDD2.n116 585
R1721 VDD2.n182 VDD2.n181 585
R1722 VDD2.n180 VDD2.n179 585
R1723 VDD2.n121 VDD2.n120 585
R1724 VDD2.n174 VDD2.n173 585
R1725 VDD2.n172 VDD2.n171 585
R1726 VDD2.n125 VDD2.n124 585
R1727 VDD2.n166 VDD2.n165 585
R1728 VDD2.n164 VDD2.n163 585
R1729 VDD2.n162 VDD2.n128 585
R1730 VDD2.n132 VDD2.n129 585
R1731 VDD2.n157 VDD2.n156 585
R1732 VDD2.n155 VDD2.n154 585
R1733 VDD2.n134 VDD2.n133 585
R1734 VDD2.n149 VDD2.n148 585
R1735 VDD2.n147 VDD2.n146 585
R1736 VDD2.n138 VDD2.n137 585
R1737 VDD2.n141 VDD2.n140 585
R1738 VDD2.n35 VDD2.n34 585
R1739 VDD2.n32 VDD2.n31 585
R1740 VDD2.n41 VDD2.n40 585
R1741 VDD2.n43 VDD2.n42 585
R1742 VDD2.n28 VDD2.n27 585
R1743 VDD2.n49 VDD2.n48 585
R1744 VDD2.n52 VDD2.n51 585
R1745 VDD2.n50 VDD2.n24 585
R1746 VDD2.n57 VDD2.n23 585
R1747 VDD2.n59 VDD2.n58 585
R1748 VDD2.n61 VDD2.n60 585
R1749 VDD2.n20 VDD2.n19 585
R1750 VDD2.n67 VDD2.n66 585
R1751 VDD2.n69 VDD2.n68 585
R1752 VDD2.n16 VDD2.n15 585
R1753 VDD2.n75 VDD2.n74 585
R1754 VDD2.n77 VDD2.n76 585
R1755 VDD2.n12 VDD2.n11 585
R1756 VDD2.n83 VDD2.n82 585
R1757 VDD2.n85 VDD2.n84 585
R1758 VDD2.n8 VDD2.n7 585
R1759 VDD2.n91 VDD2.n90 585
R1760 VDD2.n93 VDD2.n92 585
R1761 VDD2.n4 VDD2.n3 585
R1762 VDD2.n99 VDD2.n98 585
R1763 VDD2.n101 VDD2.n100 585
R1764 VDD2.n205 VDD2.n105 498.474
R1765 VDD2.n100 VDD2.n0 498.474
R1766 VDD2.t1 VDD2.n139 329.036
R1767 VDD2.t0 VDD2.n33 329.036
R1768 VDD2.n205 VDD2.n204 171.744
R1769 VDD2.n204 VDD2.n108 171.744
R1770 VDD2.n197 VDD2.n108 171.744
R1771 VDD2.n197 VDD2.n196 171.744
R1772 VDD2.n196 VDD2.n112 171.744
R1773 VDD2.n189 VDD2.n112 171.744
R1774 VDD2.n189 VDD2.n188 171.744
R1775 VDD2.n188 VDD2.n116 171.744
R1776 VDD2.n181 VDD2.n116 171.744
R1777 VDD2.n181 VDD2.n180 171.744
R1778 VDD2.n180 VDD2.n120 171.744
R1779 VDD2.n173 VDD2.n120 171.744
R1780 VDD2.n173 VDD2.n172 171.744
R1781 VDD2.n172 VDD2.n124 171.744
R1782 VDD2.n165 VDD2.n124 171.744
R1783 VDD2.n165 VDD2.n164 171.744
R1784 VDD2.n164 VDD2.n128 171.744
R1785 VDD2.n132 VDD2.n128 171.744
R1786 VDD2.n156 VDD2.n132 171.744
R1787 VDD2.n156 VDD2.n155 171.744
R1788 VDD2.n155 VDD2.n133 171.744
R1789 VDD2.n148 VDD2.n133 171.744
R1790 VDD2.n148 VDD2.n147 171.744
R1791 VDD2.n147 VDD2.n137 171.744
R1792 VDD2.n140 VDD2.n137 171.744
R1793 VDD2.n34 VDD2.n31 171.744
R1794 VDD2.n41 VDD2.n31 171.744
R1795 VDD2.n42 VDD2.n41 171.744
R1796 VDD2.n42 VDD2.n27 171.744
R1797 VDD2.n49 VDD2.n27 171.744
R1798 VDD2.n51 VDD2.n49 171.744
R1799 VDD2.n51 VDD2.n50 171.744
R1800 VDD2.n50 VDD2.n23 171.744
R1801 VDD2.n59 VDD2.n23 171.744
R1802 VDD2.n60 VDD2.n59 171.744
R1803 VDD2.n60 VDD2.n19 171.744
R1804 VDD2.n67 VDD2.n19 171.744
R1805 VDD2.n68 VDD2.n67 171.744
R1806 VDD2.n68 VDD2.n15 171.744
R1807 VDD2.n75 VDD2.n15 171.744
R1808 VDD2.n76 VDD2.n75 171.744
R1809 VDD2.n76 VDD2.n11 171.744
R1810 VDD2.n83 VDD2.n11 171.744
R1811 VDD2.n84 VDD2.n83 171.744
R1812 VDD2.n84 VDD2.n7 171.744
R1813 VDD2.n91 VDD2.n7 171.744
R1814 VDD2.n92 VDD2.n91 171.744
R1815 VDD2.n92 VDD2.n3 171.744
R1816 VDD2.n99 VDD2.n3 171.744
R1817 VDD2.n100 VDD2.n99 171.744
R1818 VDD2.n210 VDD2.n104 96.6997
R1819 VDD2.n140 VDD2.t1 85.8723
R1820 VDD2.n34 VDD2.t0 85.8723
R1821 VDD2.n210 VDD2.n209 53.3247
R1822 VDD2.n163 VDD2.n162 13.1884
R1823 VDD2.n58 VDD2.n57 13.1884
R1824 VDD2.n207 VDD2.n206 12.8005
R1825 VDD2.n166 VDD2.n127 12.8005
R1826 VDD2.n161 VDD2.n129 12.8005
R1827 VDD2.n56 VDD2.n24 12.8005
R1828 VDD2.n61 VDD2.n22 12.8005
R1829 VDD2.n102 VDD2.n101 12.8005
R1830 VDD2.n203 VDD2.n107 12.0247
R1831 VDD2.n167 VDD2.n125 12.0247
R1832 VDD2.n158 VDD2.n157 12.0247
R1833 VDD2.n53 VDD2.n52 12.0247
R1834 VDD2.n62 VDD2.n20 12.0247
R1835 VDD2.n98 VDD2.n2 12.0247
R1836 VDD2.n202 VDD2.n109 11.249
R1837 VDD2.n171 VDD2.n170 11.249
R1838 VDD2.n154 VDD2.n131 11.249
R1839 VDD2.n48 VDD2.n26 11.249
R1840 VDD2.n66 VDD2.n65 11.249
R1841 VDD2.n97 VDD2.n4 11.249
R1842 VDD2.n141 VDD2.n139 10.7239
R1843 VDD2.n35 VDD2.n33 10.7239
R1844 VDD2.n199 VDD2.n198 10.4732
R1845 VDD2.n174 VDD2.n123 10.4732
R1846 VDD2.n153 VDD2.n134 10.4732
R1847 VDD2.n47 VDD2.n28 10.4732
R1848 VDD2.n69 VDD2.n18 10.4732
R1849 VDD2.n94 VDD2.n93 10.4732
R1850 VDD2.n195 VDD2.n111 9.69747
R1851 VDD2.n175 VDD2.n121 9.69747
R1852 VDD2.n150 VDD2.n149 9.69747
R1853 VDD2.n44 VDD2.n43 9.69747
R1854 VDD2.n70 VDD2.n16 9.69747
R1855 VDD2.n90 VDD2.n6 9.69747
R1856 VDD2.n209 VDD2.n208 9.45567
R1857 VDD2.n104 VDD2.n103 9.45567
R1858 VDD2.n143 VDD2.n142 9.3005
R1859 VDD2.n145 VDD2.n144 9.3005
R1860 VDD2.n136 VDD2.n135 9.3005
R1861 VDD2.n151 VDD2.n150 9.3005
R1862 VDD2.n153 VDD2.n152 9.3005
R1863 VDD2.n131 VDD2.n130 9.3005
R1864 VDD2.n159 VDD2.n158 9.3005
R1865 VDD2.n161 VDD2.n160 9.3005
R1866 VDD2.n115 VDD2.n114 9.3005
R1867 VDD2.n192 VDD2.n191 9.3005
R1868 VDD2.n194 VDD2.n193 9.3005
R1869 VDD2.n111 VDD2.n110 9.3005
R1870 VDD2.n200 VDD2.n199 9.3005
R1871 VDD2.n202 VDD2.n201 9.3005
R1872 VDD2.n107 VDD2.n106 9.3005
R1873 VDD2.n208 VDD2.n207 9.3005
R1874 VDD2.n186 VDD2.n185 9.3005
R1875 VDD2.n184 VDD2.n183 9.3005
R1876 VDD2.n119 VDD2.n118 9.3005
R1877 VDD2.n178 VDD2.n177 9.3005
R1878 VDD2.n176 VDD2.n175 9.3005
R1879 VDD2.n123 VDD2.n122 9.3005
R1880 VDD2.n170 VDD2.n169 9.3005
R1881 VDD2.n168 VDD2.n167 9.3005
R1882 VDD2.n127 VDD2.n126 9.3005
R1883 VDD2.n79 VDD2.n78 9.3005
R1884 VDD2.n14 VDD2.n13 9.3005
R1885 VDD2.n73 VDD2.n72 9.3005
R1886 VDD2.n71 VDD2.n70 9.3005
R1887 VDD2.n18 VDD2.n17 9.3005
R1888 VDD2.n65 VDD2.n64 9.3005
R1889 VDD2.n63 VDD2.n62 9.3005
R1890 VDD2.n22 VDD2.n21 9.3005
R1891 VDD2.n37 VDD2.n36 9.3005
R1892 VDD2.n39 VDD2.n38 9.3005
R1893 VDD2.n30 VDD2.n29 9.3005
R1894 VDD2.n45 VDD2.n44 9.3005
R1895 VDD2.n47 VDD2.n46 9.3005
R1896 VDD2.n26 VDD2.n25 9.3005
R1897 VDD2.n54 VDD2.n53 9.3005
R1898 VDD2.n56 VDD2.n55 9.3005
R1899 VDD2.n81 VDD2.n80 9.3005
R1900 VDD2.n10 VDD2.n9 9.3005
R1901 VDD2.n87 VDD2.n86 9.3005
R1902 VDD2.n89 VDD2.n88 9.3005
R1903 VDD2.n6 VDD2.n5 9.3005
R1904 VDD2.n95 VDD2.n94 9.3005
R1905 VDD2.n97 VDD2.n96 9.3005
R1906 VDD2.n2 VDD2.n1 9.3005
R1907 VDD2.n103 VDD2.n102 9.3005
R1908 VDD2.n194 VDD2.n113 8.92171
R1909 VDD2.n179 VDD2.n178 8.92171
R1910 VDD2.n146 VDD2.n136 8.92171
R1911 VDD2.n40 VDD2.n30 8.92171
R1912 VDD2.n74 VDD2.n73 8.92171
R1913 VDD2.n89 VDD2.n8 8.92171
R1914 VDD2.n191 VDD2.n190 8.14595
R1915 VDD2.n182 VDD2.n119 8.14595
R1916 VDD2.n145 VDD2.n138 8.14595
R1917 VDD2.n39 VDD2.n32 8.14595
R1918 VDD2.n77 VDD2.n14 8.14595
R1919 VDD2.n86 VDD2.n85 8.14595
R1920 VDD2.n209 VDD2.n105 7.75445
R1921 VDD2.n104 VDD2.n0 7.75445
R1922 VDD2.n187 VDD2.n115 7.3702
R1923 VDD2.n183 VDD2.n117 7.3702
R1924 VDD2.n142 VDD2.n141 7.3702
R1925 VDD2.n36 VDD2.n35 7.3702
R1926 VDD2.n78 VDD2.n12 7.3702
R1927 VDD2.n82 VDD2.n10 7.3702
R1928 VDD2.n187 VDD2.n186 6.59444
R1929 VDD2.n186 VDD2.n117 6.59444
R1930 VDD2.n81 VDD2.n12 6.59444
R1931 VDD2.n82 VDD2.n81 6.59444
R1932 VDD2.n207 VDD2.n105 6.08283
R1933 VDD2.n102 VDD2.n0 6.08283
R1934 VDD2.n190 VDD2.n115 5.81868
R1935 VDD2.n183 VDD2.n182 5.81868
R1936 VDD2.n142 VDD2.n138 5.81868
R1937 VDD2.n36 VDD2.n32 5.81868
R1938 VDD2.n78 VDD2.n77 5.81868
R1939 VDD2.n85 VDD2.n10 5.81868
R1940 VDD2.n191 VDD2.n113 5.04292
R1941 VDD2.n179 VDD2.n119 5.04292
R1942 VDD2.n146 VDD2.n145 5.04292
R1943 VDD2.n40 VDD2.n39 5.04292
R1944 VDD2.n74 VDD2.n14 5.04292
R1945 VDD2.n86 VDD2.n8 5.04292
R1946 VDD2.n195 VDD2.n194 4.26717
R1947 VDD2.n178 VDD2.n121 4.26717
R1948 VDD2.n149 VDD2.n136 4.26717
R1949 VDD2.n43 VDD2.n30 4.26717
R1950 VDD2.n73 VDD2.n16 4.26717
R1951 VDD2.n90 VDD2.n89 4.26717
R1952 VDD2.n198 VDD2.n111 3.49141
R1953 VDD2.n175 VDD2.n174 3.49141
R1954 VDD2.n150 VDD2.n134 3.49141
R1955 VDD2.n44 VDD2.n28 3.49141
R1956 VDD2.n70 VDD2.n69 3.49141
R1957 VDD2.n93 VDD2.n6 3.49141
R1958 VDD2.n199 VDD2.n109 2.71565
R1959 VDD2.n171 VDD2.n123 2.71565
R1960 VDD2.n154 VDD2.n153 2.71565
R1961 VDD2.n48 VDD2.n47 2.71565
R1962 VDD2.n66 VDD2.n18 2.71565
R1963 VDD2.n94 VDD2.n4 2.71565
R1964 VDD2.n143 VDD2.n139 2.41282
R1965 VDD2.n37 VDD2.n33 2.41282
R1966 VDD2.n203 VDD2.n202 1.93989
R1967 VDD2.n170 VDD2.n125 1.93989
R1968 VDD2.n157 VDD2.n131 1.93989
R1969 VDD2.n52 VDD2.n26 1.93989
R1970 VDD2.n65 VDD2.n20 1.93989
R1971 VDD2.n98 VDD2.n97 1.93989
R1972 VDD2.n206 VDD2.n107 1.16414
R1973 VDD2.n167 VDD2.n166 1.16414
R1974 VDD2.n158 VDD2.n129 1.16414
R1975 VDD2.n53 VDD2.n24 1.16414
R1976 VDD2.n62 VDD2.n61 1.16414
R1977 VDD2.n101 VDD2.n2 1.16414
R1978 VDD2 VDD2.n210 0.416448
R1979 VDD2.n163 VDD2.n127 0.388379
R1980 VDD2.n162 VDD2.n161 0.388379
R1981 VDD2.n57 VDD2.n56 0.388379
R1982 VDD2.n58 VDD2.n22 0.388379
R1983 VDD2.n208 VDD2.n106 0.155672
R1984 VDD2.n201 VDD2.n106 0.155672
R1985 VDD2.n201 VDD2.n200 0.155672
R1986 VDD2.n200 VDD2.n110 0.155672
R1987 VDD2.n193 VDD2.n110 0.155672
R1988 VDD2.n193 VDD2.n192 0.155672
R1989 VDD2.n192 VDD2.n114 0.155672
R1990 VDD2.n185 VDD2.n114 0.155672
R1991 VDD2.n185 VDD2.n184 0.155672
R1992 VDD2.n184 VDD2.n118 0.155672
R1993 VDD2.n177 VDD2.n118 0.155672
R1994 VDD2.n177 VDD2.n176 0.155672
R1995 VDD2.n176 VDD2.n122 0.155672
R1996 VDD2.n169 VDD2.n122 0.155672
R1997 VDD2.n169 VDD2.n168 0.155672
R1998 VDD2.n168 VDD2.n126 0.155672
R1999 VDD2.n160 VDD2.n126 0.155672
R2000 VDD2.n160 VDD2.n159 0.155672
R2001 VDD2.n159 VDD2.n130 0.155672
R2002 VDD2.n152 VDD2.n130 0.155672
R2003 VDD2.n152 VDD2.n151 0.155672
R2004 VDD2.n151 VDD2.n135 0.155672
R2005 VDD2.n144 VDD2.n135 0.155672
R2006 VDD2.n144 VDD2.n143 0.155672
R2007 VDD2.n38 VDD2.n37 0.155672
R2008 VDD2.n38 VDD2.n29 0.155672
R2009 VDD2.n45 VDD2.n29 0.155672
R2010 VDD2.n46 VDD2.n45 0.155672
R2011 VDD2.n46 VDD2.n25 0.155672
R2012 VDD2.n54 VDD2.n25 0.155672
R2013 VDD2.n55 VDD2.n54 0.155672
R2014 VDD2.n55 VDD2.n21 0.155672
R2015 VDD2.n63 VDD2.n21 0.155672
R2016 VDD2.n64 VDD2.n63 0.155672
R2017 VDD2.n64 VDD2.n17 0.155672
R2018 VDD2.n71 VDD2.n17 0.155672
R2019 VDD2.n72 VDD2.n71 0.155672
R2020 VDD2.n72 VDD2.n13 0.155672
R2021 VDD2.n79 VDD2.n13 0.155672
R2022 VDD2.n80 VDD2.n79 0.155672
R2023 VDD2.n80 VDD2.n9 0.155672
R2024 VDD2.n87 VDD2.n9 0.155672
R2025 VDD2.n88 VDD2.n87 0.155672
R2026 VDD2.n88 VDD2.n5 0.155672
R2027 VDD2.n95 VDD2.n5 0.155672
R2028 VDD2.n96 VDD2.n95 0.155672
R2029 VDD2.n96 VDD2.n1 0.155672
R2030 VDD2.n103 VDD2.n1 0.155672
R2031 VP.n0 VP.t0 511.582
R2032 VP.n0 VP.t1 464.572
R2033 VP VP.n0 0.146778
R2034 VDD1.n101 VDD1.n100 585
R2035 VDD1.n99 VDD1.n98 585
R2036 VDD1.n4 VDD1.n3 585
R2037 VDD1.n93 VDD1.n92 585
R2038 VDD1.n91 VDD1.n90 585
R2039 VDD1.n8 VDD1.n7 585
R2040 VDD1.n85 VDD1.n84 585
R2041 VDD1.n83 VDD1.n82 585
R2042 VDD1.n12 VDD1.n11 585
R2043 VDD1.n77 VDD1.n76 585
R2044 VDD1.n75 VDD1.n74 585
R2045 VDD1.n16 VDD1.n15 585
R2046 VDD1.n69 VDD1.n68 585
R2047 VDD1.n67 VDD1.n66 585
R2048 VDD1.n20 VDD1.n19 585
R2049 VDD1.n61 VDD1.n60 585
R2050 VDD1.n59 VDD1.n58 585
R2051 VDD1.n57 VDD1.n23 585
R2052 VDD1.n27 VDD1.n24 585
R2053 VDD1.n52 VDD1.n51 585
R2054 VDD1.n50 VDD1.n49 585
R2055 VDD1.n29 VDD1.n28 585
R2056 VDD1.n44 VDD1.n43 585
R2057 VDD1.n42 VDD1.n41 585
R2058 VDD1.n33 VDD1.n32 585
R2059 VDD1.n36 VDD1.n35 585
R2060 VDD1.n140 VDD1.n139 585
R2061 VDD1.n137 VDD1.n136 585
R2062 VDD1.n146 VDD1.n145 585
R2063 VDD1.n148 VDD1.n147 585
R2064 VDD1.n133 VDD1.n132 585
R2065 VDD1.n154 VDD1.n153 585
R2066 VDD1.n157 VDD1.n156 585
R2067 VDD1.n155 VDD1.n129 585
R2068 VDD1.n162 VDD1.n128 585
R2069 VDD1.n164 VDD1.n163 585
R2070 VDD1.n166 VDD1.n165 585
R2071 VDD1.n125 VDD1.n124 585
R2072 VDD1.n172 VDD1.n171 585
R2073 VDD1.n174 VDD1.n173 585
R2074 VDD1.n121 VDD1.n120 585
R2075 VDD1.n180 VDD1.n179 585
R2076 VDD1.n182 VDD1.n181 585
R2077 VDD1.n117 VDD1.n116 585
R2078 VDD1.n188 VDD1.n187 585
R2079 VDD1.n190 VDD1.n189 585
R2080 VDD1.n113 VDD1.n112 585
R2081 VDD1.n196 VDD1.n195 585
R2082 VDD1.n198 VDD1.n197 585
R2083 VDD1.n109 VDD1.n108 585
R2084 VDD1.n204 VDD1.n203 585
R2085 VDD1.n206 VDD1.n205 585
R2086 VDD1.n100 VDD1.n0 498.474
R2087 VDD1.n205 VDD1.n105 498.474
R2088 VDD1.t1 VDD1.n34 329.036
R2089 VDD1.t0 VDD1.n138 329.036
R2090 VDD1.n100 VDD1.n99 171.744
R2091 VDD1.n99 VDD1.n3 171.744
R2092 VDD1.n92 VDD1.n3 171.744
R2093 VDD1.n92 VDD1.n91 171.744
R2094 VDD1.n91 VDD1.n7 171.744
R2095 VDD1.n84 VDD1.n7 171.744
R2096 VDD1.n84 VDD1.n83 171.744
R2097 VDD1.n83 VDD1.n11 171.744
R2098 VDD1.n76 VDD1.n11 171.744
R2099 VDD1.n76 VDD1.n75 171.744
R2100 VDD1.n75 VDD1.n15 171.744
R2101 VDD1.n68 VDD1.n15 171.744
R2102 VDD1.n68 VDD1.n67 171.744
R2103 VDD1.n67 VDD1.n19 171.744
R2104 VDD1.n60 VDD1.n19 171.744
R2105 VDD1.n60 VDD1.n59 171.744
R2106 VDD1.n59 VDD1.n23 171.744
R2107 VDD1.n27 VDD1.n23 171.744
R2108 VDD1.n51 VDD1.n27 171.744
R2109 VDD1.n51 VDD1.n50 171.744
R2110 VDD1.n50 VDD1.n28 171.744
R2111 VDD1.n43 VDD1.n28 171.744
R2112 VDD1.n43 VDD1.n42 171.744
R2113 VDD1.n42 VDD1.n32 171.744
R2114 VDD1.n35 VDD1.n32 171.744
R2115 VDD1.n139 VDD1.n136 171.744
R2116 VDD1.n146 VDD1.n136 171.744
R2117 VDD1.n147 VDD1.n146 171.744
R2118 VDD1.n147 VDD1.n132 171.744
R2119 VDD1.n154 VDD1.n132 171.744
R2120 VDD1.n156 VDD1.n154 171.744
R2121 VDD1.n156 VDD1.n155 171.744
R2122 VDD1.n155 VDD1.n128 171.744
R2123 VDD1.n164 VDD1.n128 171.744
R2124 VDD1.n165 VDD1.n164 171.744
R2125 VDD1.n165 VDD1.n124 171.744
R2126 VDD1.n172 VDD1.n124 171.744
R2127 VDD1.n173 VDD1.n172 171.744
R2128 VDD1.n173 VDD1.n120 171.744
R2129 VDD1.n180 VDD1.n120 171.744
R2130 VDD1.n181 VDD1.n180 171.744
R2131 VDD1.n181 VDD1.n116 171.744
R2132 VDD1.n188 VDD1.n116 171.744
R2133 VDD1.n189 VDD1.n188 171.744
R2134 VDD1.n189 VDD1.n112 171.744
R2135 VDD1.n196 VDD1.n112 171.744
R2136 VDD1.n197 VDD1.n196 171.744
R2137 VDD1.n197 VDD1.n108 171.744
R2138 VDD1.n204 VDD1.n108 171.744
R2139 VDD1.n205 VDD1.n204 171.744
R2140 VDD1 VDD1.n209 97.5823
R2141 VDD1.n35 VDD1.t1 85.8723
R2142 VDD1.n139 VDD1.t0 85.8723
R2143 VDD1 VDD1.n104 53.7407
R2144 VDD1.n58 VDD1.n57 13.1884
R2145 VDD1.n163 VDD1.n162 13.1884
R2146 VDD1.n102 VDD1.n101 12.8005
R2147 VDD1.n61 VDD1.n22 12.8005
R2148 VDD1.n56 VDD1.n24 12.8005
R2149 VDD1.n161 VDD1.n129 12.8005
R2150 VDD1.n166 VDD1.n127 12.8005
R2151 VDD1.n207 VDD1.n206 12.8005
R2152 VDD1.n98 VDD1.n2 12.0247
R2153 VDD1.n62 VDD1.n20 12.0247
R2154 VDD1.n53 VDD1.n52 12.0247
R2155 VDD1.n158 VDD1.n157 12.0247
R2156 VDD1.n167 VDD1.n125 12.0247
R2157 VDD1.n203 VDD1.n107 12.0247
R2158 VDD1.n97 VDD1.n4 11.249
R2159 VDD1.n66 VDD1.n65 11.249
R2160 VDD1.n49 VDD1.n26 11.249
R2161 VDD1.n153 VDD1.n131 11.249
R2162 VDD1.n171 VDD1.n170 11.249
R2163 VDD1.n202 VDD1.n109 11.249
R2164 VDD1.n36 VDD1.n34 10.7239
R2165 VDD1.n140 VDD1.n138 10.7239
R2166 VDD1.n94 VDD1.n93 10.4732
R2167 VDD1.n69 VDD1.n18 10.4732
R2168 VDD1.n48 VDD1.n29 10.4732
R2169 VDD1.n152 VDD1.n133 10.4732
R2170 VDD1.n174 VDD1.n123 10.4732
R2171 VDD1.n199 VDD1.n198 10.4732
R2172 VDD1.n90 VDD1.n6 9.69747
R2173 VDD1.n70 VDD1.n16 9.69747
R2174 VDD1.n45 VDD1.n44 9.69747
R2175 VDD1.n149 VDD1.n148 9.69747
R2176 VDD1.n175 VDD1.n121 9.69747
R2177 VDD1.n195 VDD1.n111 9.69747
R2178 VDD1.n104 VDD1.n103 9.45567
R2179 VDD1.n209 VDD1.n208 9.45567
R2180 VDD1.n38 VDD1.n37 9.3005
R2181 VDD1.n40 VDD1.n39 9.3005
R2182 VDD1.n31 VDD1.n30 9.3005
R2183 VDD1.n46 VDD1.n45 9.3005
R2184 VDD1.n48 VDD1.n47 9.3005
R2185 VDD1.n26 VDD1.n25 9.3005
R2186 VDD1.n54 VDD1.n53 9.3005
R2187 VDD1.n56 VDD1.n55 9.3005
R2188 VDD1.n10 VDD1.n9 9.3005
R2189 VDD1.n87 VDD1.n86 9.3005
R2190 VDD1.n89 VDD1.n88 9.3005
R2191 VDD1.n6 VDD1.n5 9.3005
R2192 VDD1.n95 VDD1.n94 9.3005
R2193 VDD1.n97 VDD1.n96 9.3005
R2194 VDD1.n2 VDD1.n1 9.3005
R2195 VDD1.n103 VDD1.n102 9.3005
R2196 VDD1.n81 VDD1.n80 9.3005
R2197 VDD1.n79 VDD1.n78 9.3005
R2198 VDD1.n14 VDD1.n13 9.3005
R2199 VDD1.n73 VDD1.n72 9.3005
R2200 VDD1.n71 VDD1.n70 9.3005
R2201 VDD1.n18 VDD1.n17 9.3005
R2202 VDD1.n65 VDD1.n64 9.3005
R2203 VDD1.n63 VDD1.n62 9.3005
R2204 VDD1.n22 VDD1.n21 9.3005
R2205 VDD1.n184 VDD1.n183 9.3005
R2206 VDD1.n119 VDD1.n118 9.3005
R2207 VDD1.n178 VDD1.n177 9.3005
R2208 VDD1.n176 VDD1.n175 9.3005
R2209 VDD1.n123 VDD1.n122 9.3005
R2210 VDD1.n170 VDD1.n169 9.3005
R2211 VDD1.n168 VDD1.n167 9.3005
R2212 VDD1.n127 VDD1.n126 9.3005
R2213 VDD1.n142 VDD1.n141 9.3005
R2214 VDD1.n144 VDD1.n143 9.3005
R2215 VDD1.n135 VDD1.n134 9.3005
R2216 VDD1.n150 VDD1.n149 9.3005
R2217 VDD1.n152 VDD1.n151 9.3005
R2218 VDD1.n131 VDD1.n130 9.3005
R2219 VDD1.n159 VDD1.n158 9.3005
R2220 VDD1.n161 VDD1.n160 9.3005
R2221 VDD1.n186 VDD1.n185 9.3005
R2222 VDD1.n115 VDD1.n114 9.3005
R2223 VDD1.n192 VDD1.n191 9.3005
R2224 VDD1.n194 VDD1.n193 9.3005
R2225 VDD1.n111 VDD1.n110 9.3005
R2226 VDD1.n200 VDD1.n199 9.3005
R2227 VDD1.n202 VDD1.n201 9.3005
R2228 VDD1.n107 VDD1.n106 9.3005
R2229 VDD1.n208 VDD1.n207 9.3005
R2230 VDD1.n89 VDD1.n8 8.92171
R2231 VDD1.n74 VDD1.n73 8.92171
R2232 VDD1.n41 VDD1.n31 8.92171
R2233 VDD1.n145 VDD1.n135 8.92171
R2234 VDD1.n179 VDD1.n178 8.92171
R2235 VDD1.n194 VDD1.n113 8.92171
R2236 VDD1.n86 VDD1.n85 8.14595
R2237 VDD1.n77 VDD1.n14 8.14595
R2238 VDD1.n40 VDD1.n33 8.14595
R2239 VDD1.n144 VDD1.n137 8.14595
R2240 VDD1.n182 VDD1.n119 8.14595
R2241 VDD1.n191 VDD1.n190 8.14595
R2242 VDD1.n104 VDD1.n0 7.75445
R2243 VDD1.n209 VDD1.n105 7.75445
R2244 VDD1.n82 VDD1.n10 7.3702
R2245 VDD1.n78 VDD1.n12 7.3702
R2246 VDD1.n37 VDD1.n36 7.3702
R2247 VDD1.n141 VDD1.n140 7.3702
R2248 VDD1.n183 VDD1.n117 7.3702
R2249 VDD1.n187 VDD1.n115 7.3702
R2250 VDD1.n82 VDD1.n81 6.59444
R2251 VDD1.n81 VDD1.n12 6.59444
R2252 VDD1.n186 VDD1.n117 6.59444
R2253 VDD1.n187 VDD1.n186 6.59444
R2254 VDD1.n102 VDD1.n0 6.08283
R2255 VDD1.n207 VDD1.n105 6.08283
R2256 VDD1.n85 VDD1.n10 5.81868
R2257 VDD1.n78 VDD1.n77 5.81868
R2258 VDD1.n37 VDD1.n33 5.81868
R2259 VDD1.n141 VDD1.n137 5.81868
R2260 VDD1.n183 VDD1.n182 5.81868
R2261 VDD1.n190 VDD1.n115 5.81868
R2262 VDD1.n86 VDD1.n8 5.04292
R2263 VDD1.n74 VDD1.n14 5.04292
R2264 VDD1.n41 VDD1.n40 5.04292
R2265 VDD1.n145 VDD1.n144 5.04292
R2266 VDD1.n179 VDD1.n119 5.04292
R2267 VDD1.n191 VDD1.n113 5.04292
R2268 VDD1.n90 VDD1.n89 4.26717
R2269 VDD1.n73 VDD1.n16 4.26717
R2270 VDD1.n44 VDD1.n31 4.26717
R2271 VDD1.n148 VDD1.n135 4.26717
R2272 VDD1.n178 VDD1.n121 4.26717
R2273 VDD1.n195 VDD1.n194 4.26717
R2274 VDD1.n93 VDD1.n6 3.49141
R2275 VDD1.n70 VDD1.n69 3.49141
R2276 VDD1.n45 VDD1.n29 3.49141
R2277 VDD1.n149 VDD1.n133 3.49141
R2278 VDD1.n175 VDD1.n174 3.49141
R2279 VDD1.n198 VDD1.n111 3.49141
R2280 VDD1.n94 VDD1.n4 2.71565
R2281 VDD1.n66 VDD1.n18 2.71565
R2282 VDD1.n49 VDD1.n48 2.71565
R2283 VDD1.n153 VDD1.n152 2.71565
R2284 VDD1.n171 VDD1.n123 2.71565
R2285 VDD1.n199 VDD1.n109 2.71565
R2286 VDD1.n38 VDD1.n34 2.41282
R2287 VDD1.n142 VDD1.n138 2.41282
R2288 VDD1.n98 VDD1.n97 1.93989
R2289 VDD1.n65 VDD1.n20 1.93989
R2290 VDD1.n52 VDD1.n26 1.93989
R2291 VDD1.n157 VDD1.n131 1.93989
R2292 VDD1.n170 VDD1.n125 1.93989
R2293 VDD1.n203 VDD1.n202 1.93989
R2294 VDD1.n101 VDD1.n2 1.16414
R2295 VDD1.n62 VDD1.n61 1.16414
R2296 VDD1.n53 VDD1.n24 1.16414
R2297 VDD1.n158 VDD1.n129 1.16414
R2298 VDD1.n167 VDD1.n166 1.16414
R2299 VDD1.n206 VDD1.n107 1.16414
R2300 VDD1.n58 VDD1.n22 0.388379
R2301 VDD1.n57 VDD1.n56 0.388379
R2302 VDD1.n162 VDD1.n161 0.388379
R2303 VDD1.n163 VDD1.n127 0.388379
R2304 VDD1.n103 VDD1.n1 0.155672
R2305 VDD1.n96 VDD1.n1 0.155672
R2306 VDD1.n96 VDD1.n95 0.155672
R2307 VDD1.n95 VDD1.n5 0.155672
R2308 VDD1.n88 VDD1.n5 0.155672
R2309 VDD1.n88 VDD1.n87 0.155672
R2310 VDD1.n87 VDD1.n9 0.155672
R2311 VDD1.n80 VDD1.n9 0.155672
R2312 VDD1.n80 VDD1.n79 0.155672
R2313 VDD1.n79 VDD1.n13 0.155672
R2314 VDD1.n72 VDD1.n13 0.155672
R2315 VDD1.n72 VDD1.n71 0.155672
R2316 VDD1.n71 VDD1.n17 0.155672
R2317 VDD1.n64 VDD1.n17 0.155672
R2318 VDD1.n64 VDD1.n63 0.155672
R2319 VDD1.n63 VDD1.n21 0.155672
R2320 VDD1.n55 VDD1.n21 0.155672
R2321 VDD1.n55 VDD1.n54 0.155672
R2322 VDD1.n54 VDD1.n25 0.155672
R2323 VDD1.n47 VDD1.n25 0.155672
R2324 VDD1.n47 VDD1.n46 0.155672
R2325 VDD1.n46 VDD1.n30 0.155672
R2326 VDD1.n39 VDD1.n30 0.155672
R2327 VDD1.n39 VDD1.n38 0.155672
R2328 VDD1.n143 VDD1.n142 0.155672
R2329 VDD1.n143 VDD1.n134 0.155672
R2330 VDD1.n150 VDD1.n134 0.155672
R2331 VDD1.n151 VDD1.n150 0.155672
R2332 VDD1.n151 VDD1.n130 0.155672
R2333 VDD1.n159 VDD1.n130 0.155672
R2334 VDD1.n160 VDD1.n159 0.155672
R2335 VDD1.n160 VDD1.n126 0.155672
R2336 VDD1.n168 VDD1.n126 0.155672
R2337 VDD1.n169 VDD1.n168 0.155672
R2338 VDD1.n169 VDD1.n122 0.155672
R2339 VDD1.n176 VDD1.n122 0.155672
R2340 VDD1.n177 VDD1.n176 0.155672
R2341 VDD1.n177 VDD1.n118 0.155672
R2342 VDD1.n184 VDD1.n118 0.155672
R2343 VDD1.n185 VDD1.n184 0.155672
R2344 VDD1.n185 VDD1.n114 0.155672
R2345 VDD1.n192 VDD1.n114 0.155672
R2346 VDD1.n193 VDD1.n192 0.155672
R2347 VDD1.n193 VDD1.n110 0.155672
R2348 VDD1.n200 VDD1.n110 0.155672
R2349 VDD1.n201 VDD1.n200 0.155672
R2350 VDD1.n201 VDD1.n106 0.155672
R2351 VDD1.n208 VDD1.n106 0.155672
C0 VN VTAIL 3.05537f
C1 B w_n1634_n4878# 9.55231f
C2 VDD1 w_n1634_n4878# 2.1818f
C3 VP w_n1634_n4878# 2.49194f
C4 VDD2 w_n1634_n4878# 2.19278f
C5 VDD1 B 2.09285f
C6 VTAIL w_n1634_n4878# 3.95539f
C7 B VP 1.25629f
C8 VDD2 B 2.11197f
C9 VDD1 VP 3.92722f
C10 VDD1 VDD2 0.528877f
C11 VN w_n1634_n4878# 2.28654f
C12 VDD2 VP 0.280797f
C13 VTAIL B 4.55866f
C14 VDD1 VTAIL 7.425479f
C15 VTAIL VP 3.07004f
C16 VDD2 VTAIL 7.4625f
C17 VN B 0.923699f
C18 VDD1 VN 0.14754f
C19 VN VP 6.25803f
C20 VDD2 VN 3.79949f
C21 VDD2 VSUBS 1.065567f
C22 VDD1 VSUBS 5.29897f
C23 VTAIL VSUBS 1.126377f
C24 VN VSUBS 9.357861f
C25 VP VSUBS 1.585583f
C26 B VSUBS 3.59634f
C27 w_n1634_n4878# VSUBS 97.35371f
C28 VDD1.n0 VSUBS 0.030826f
C29 VDD1.n1 VSUBS 0.027578f
C30 VDD1.n2 VSUBS 0.014819f
C31 VDD1.n3 VSUBS 0.035027f
C32 VDD1.n4 VSUBS 0.015691f
C33 VDD1.n5 VSUBS 0.027578f
C34 VDD1.n6 VSUBS 0.014819f
C35 VDD1.n7 VSUBS 0.035027f
C36 VDD1.n8 VSUBS 0.015691f
C37 VDD1.n9 VSUBS 0.027578f
C38 VDD1.n10 VSUBS 0.014819f
C39 VDD1.n11 VSUBS 0.035027f
C40 VDD1.n12 VSUBS 0.015691f
C41 VDD1.n13 VSUBS 0.027578f
C42 VDD1.n14 VSUBS 0.014819f
C43 VDD1.n15 VSUBS 0.035027f
C44 VDD1.n16 VSUBS 0.015691f
C45 VDD1.n17 VSUBS 0.027578f
C46 VDD1.n18 VSUBS 0.014819f
C47 VDD1.n19 VSUBS 0.035027f
C48 VDD1.n20 VSUBS 0.015691f
C49 VDD1.n21 VSUBS 0.027578f
C50 VDD1.n22 VSUBS 0.014819f
C51 VDD1.n23 VSUBS 0.035027f
C52 VDD1.n24 VSUBS 0.015691f
C53 VDD1.n25 VSUBS 0.027578f
C54 VDD1.n26 VSUBS 0.014819f
C55 VDD1.n27 VSUBS 0.035027f
C56 VDD1.n28 VSUBS 0.035027f
C57 VDD1.n29 VSUBS 0.015691f
C58 VDD1.n30 VSUBS 0.027578f
C59 VDD1.n31 VSUBS 0.014819f
C60 VDD1.n32 VSUBS 0.035027f
C61 VDD1.n33 VSUBS 0.015691f
C62 VDD1.n34 VSUBS 0.311333f
C63 VDD1.t1 VSUBS 0.076182f
C64 VDD1.n35 VSUBS 0.02627f
C65 VDD1.n36 VSUBS 0.026349f
C66 VDD1.n37 VSUBS 0.014819f
C67 VDD1.n38 VSUBS 2.26727f
C68 VDD1.n39 VSUBS 0.027578f
C69 VDD1.n40 VSUBS 0.014819f
C70 VDD1.n41 VSUBS 0.015691f
C71 VDD1.n42 VSUBS 0.035027f
C72 VDD1.n43 VSUBS 0.035027f
C73 VDD1.n44 VSUBS 0.015691f
C74 VDD1.n45 VSUBS 0.014819f
C75 VDD1.n46 VSUBS 0.027578f
C76 VDD1.n47 VSUBS 0.027578f
C77 VDD1.n48 VSUBS 0.014819f
C78 VDD1.n49 VSUBS 0.015691f
C79 VDD1.n50 VSUBS 0.035027f
C80 VDD1.n51 VSUBS 0.035027f
C81 VDD1.n52 VSUBS 0.015691f
C82 VDD1.n53 VSUBS 0.014819f
C83 VDD1.n54 VSUBS 0.027578f
C84 VDD1.n55 VSUBS 0.027578f
C85 VDD1.n56 VSUBS 0.014819f
C86 VDD1.n57 VSUBS 0.015255f
C87 VDD1.n58 VSUBS 0.015255f
C88 VDD1.n59 VSUBS 0.035027f
C89 VDD1.n60 VSUBS 0.035027f
C90 VDD1.n61 VSUBS 0.015691f
C91 VDD1.n62 VSUBS 0.014819f
C92 VDD1.n63 VSUBS 0.027578f
C93 VDD1.n64 VSUBS 0.027578f
C94 VDD1.n65 VSUBS 0.014819f
C95 VDD1.n66 VSUBS 0.015691f
C96 VDD1.n67 VSUBS 0.035027f
C97 VDD1.n68 VSUBS 0.035027f
C98 VDD1.n69 VSUBS 0.015691f
C99 VDD1.n70 VSUBS 0.014819f
C100 VDD1.n71 VSUBS 0.027578f
C101 VDD1.n72 VSUBS 0.027578f
C102 VDD1.n73 VSUBS 0.014819f
C103 VDD1.n74 VSUBS 0.015691f
C104 VDD1.n75 VSUBS 0.035027f
C105 VDD1.n76 VSUBS 0.035027f
C106 VDD1.n77 VSUBS 0.015691f
C107 VDD1.n78 VSUBS 0.014819f
C108 VDD1.n79 VSUBS 0.027578f
C109 VDD1.n80 VSUBS 0.027578f
C110 VDD1.n81 VSUBS 0.014819f
C111 VDD1.n82 VSUBS 0.015691f
C112 VDD1.n83 VSUBS 0.035027f
C113 VDD1.n84 VSUBS 0.035027f
C114 VDD1.n85 VSUBS 0.015691f
C115 VDD1.n86 VSUBS 0.014819f
C116 VDD1.n87 VSUBS 0.027578f
C117 VDD1.n88 VSUBS 0.027578f
C118 VDD1.n89 VSUBS 0.014819f
C119 VDD1.n90 VSUBS 0.015691f
C120 VDD1.n91 VSUBS 0.035027f
C121 VDD1.n92 VSUBS 0.035027f
C122 VDD1.n93 VSUBS 0.015691f
C123 VDD1.n94 VSUBS 0.014819f
C124 VDD1.n95 VSUBS 0.027578f
C125 VDD1.n96 VSUBS 0.027578f
C126 VDD1.n97 VSUBS 0.014819f
C127 VDD1.n98 VSUBS 0.015691f
C128 VDD1.n99 VSUBS 0.035027f
C129 VDD1.n100 VSUBS 0.089044f
C130 VDD1.n101 VSUBS 0.015691f
C131 VDD1.n102 VSUBS 0.029101f
C132 VDD1.n103 VSUBS 0.072409f
C133 VDD1.n104 VSUBS 0.089016f
C134 VDD1.n105 VSUBS 0.030826f
C135 VDD1.n106 VSUBS 0.027578f
C136 VDD1.n107 VSUBS 0.014819f
C137 VDD1.n108 VSUBS 0.035027f
C138 VDD1.n109 VSUBS 0.015691f
C139 VDD1.n110 VSUBS 0.027578f
C140 VDD1.n111 VSUBS 0.014819f
C141 VDD1.n112 VSUBS 0.035027f
C142 VDD1.n113 VSUBS 0.015691f
C143 VDD1.n114 VSUBS 0.027578f
C144 VDD1.n115 VSUBS 0.014819f
C145 VDD1.n116 VSUBS 0.035027f
C146 VDD1.n117 VSUBS 0.015691f
C147 VDD1.n118 VSUBS 0.027578f
C148 VDD1.n119 VSUBS 0.014819f
C149 VDD1.n120 VSUBS 0.035027f
C150 VDD1.n121 VSUBS 0.015691f
C151 VDD1.n122 VSUBS 0.027578f
C152 VDD1.n123 VSUBS 0.014819f
C153 VDD1.n124 VSUBS 0.035027f
C154 VDD1.n125 VSUBS 0.015691f
C155 VDD1.n126 VSUBS 0.027578f
C156 VDD1.n127 VSUBS 0.014819f
C157 VDD1.n128 VSUBS 0.035027f
C158 VDD1.n129 VSUBS 0.015691f
C159 VDD1.n130 VSUBS 0.027578f
C160 VDD1.n131 VSUBS 0.014819f
C161 VDD1.n132 VSUBS 0.035027f
C162 VDD1.n133 VSUBS 0.015691f
C163 VDD1.n134 VSUBS 0.027578f
C164 VDD1.n135 VSUBS 0.014819f
C165 VDD1.n136 VSUBS 0.035027f
C166 VDD1.n137 VSUBS 0.015691f
C167 VDD1.n138 VSUBS 0.311333f
C168 VDD1.t0 VSUBS 0.076182f
C169 VDD1.n139 VSUBS 0.02627f
C170 VDD1.n140 VSUBS 0.026349f
C171 VDD1.n141 VSUBS 0.014819f
C172 VDD1.n142 VSUBS 2.26727f
C173 VDD1.n143 VSUBS 0.027578f
C174 VDD1.n144 VSUBS 0.014819f
C175 VDD1.n145 VSUBS 0.015691f
C176 VDD1.n146 VSUBS 0.035027f
C177 VDD1.n147 VSUBS 0.035027f
C178 VDD1.n148 VSUBS 0.015691f
C179 VDD1.n149 VSUBS 0.014819f
C180 VDD1.n150 VSUBS 0.027578f
C181 VDD1.n151 VSUBS 0.027578f
C182 VDD1.n152 VSUBS 0.014819f
C183 VDD1.n153 VSUBS 0.015691f
C184 VDD1.n154 VSUBS 0.035027f
C185 VDD1.n155 VSUBS 0.035027f
C186 VDD1.n156 VSUBS 0.035027f
C187 VDD1.n157 VSUBS 0.015691f
C188 VDD1.n158 VSUBS 0.014819f
C189 VDD1.n159 VSUBS 0.027578f
C190 VDD1.n160 VSUBS 0.027578f
C191 VDD1.n161 VSUBS 0.014819f
C192 VDD1.n162 VSUBS 0.015255f
C193 VDD1.n163 VSUBS 0.015255f
C194 VDD1.n164 VSUBS 0.035027f
C195 VDD1.n165 VSUBS 0.035027f
C196 VDD1.n166 VSUBS 0.015691f
C197 VDD1.n167 VSUBS 0.014819f
C198 VDD1.n168 VSUBS 0.027578f
C199 VDD1.n169 VSUBS 0.027578f
C200 VDD1.n170 VSUBS 0.014819f
C201 VDD1.n171 VSUBS 0.015691f
C202 VDD1.n172 VSUBS 0.035027f
C203 VDD1.n173 VSUBS 0.035027f
C204 VDD1.n174 VSUBS 0.015691f
C205 VDD1.n175 VSUBS 0.014819f
C206 VDD1.n176 VSUBS 0.027578f
C207 VDD1.n177 VSUBS 0.027578f
C208 VDD1.n178 VSUBS 0.014819f
C209 VDD1.n179 VSUBS 0.015691f
C210 VDD1.n180 VSUBS 0.035027f
C211 VDD1.n181 VSUBS 0.035027f
C212 VDD1.n182 VSUBS 0.015691f
C213 VDD1.n183 VSUBS 0.014819f
C214 VDD1.n184 VSUBS 0.027578f
C215 VDD1.n185 VSUBS 0.027578f
C216 VDD1.n186 VSUBS 0.014819f
C217 VDD1.n187 VSUBS 0.015691f
C218 VDD1.n188 VSUBS 0.035027f
C219 VDD1.n189 VSUBS 0.035027f
C220 VDD1.n190 VSUBS 0.015691f
C221 VDD1.n191 VSUBS 0.014819f
C222 VDD1.n192 VSUBS 0.027578f
C223 VDD1.n193 VSUBS 0.027578f
C224 VDD1.n194 VSUBS 0.014819f
C225 VDD1.n195 VSUBS 0.015691f
C226 VDD1.n196 VSUBS 0.035027f
C227 VDD1.n197 VSUBS 0.035027f
C228 VDD1.n198 VSUBS 0.015691f
C229 VDD1.n199 VSUBS 0.014819f
C230 VDD1.n200 VSUBS 0.027578f
C231 VDD1.n201 VSUBS 0.027578f
C232 VDD1.n202 VSUBS 0.014819f
C233 VDD1.n203 VSUBS 0.015691f
C234 VDD1.n204 VSUBS 0.035027f
C235 VDD1.n205 VSUBS 0.089044f
C236 VDD1.n206 VSUBS 0.015691f
C237 VDD1.n207 VSUBS 0.029101f
C238 VDD1.n208 VSUBS 0.072409f
C239 VDD1.n209 VSUBS 1.05525f
C240 VP.t0 VSUBS 4.43308f
C241 VP.t1 VSUBS 4.08429f
C242 VP.n0 VSUBS 7.23404f
C243 VDD2.n0 VSUBS 0.031029f
C244 VDD2.n1 VSUBS 0.027759f
C245 VDD2.n2 VSUBS 0.014916f
C246 VDD2.n3 VSUBS 0.035257f
C247 VDD2.n4 VSUBS 0.015794f
C248 VDD2.n5 VSUBS 0.027759f
C249 VDD2.n6 VSUBS 0.014916f
C250 VDD2.n7 VSUBS 0.035257f
C251 VDD2.n8 VSUBS 0.015794f
C252 VDD2.n9 VSUBS 0.027759f
C253 VDD2.n10 VSUBS 0.014916f
C254 VDD2.n11 VSUBS 0.035257f
C255 VDD2.n12 VSUBS 0.015794f
C256 VDD2.n13 VSUBS 0.027759f
C257 VDD2.n14 VSUBS 0.014916f
C258 VDD2.n15 VSUBS 0.035257f
C259 VDD2.n16 VSUBS 0.015794f
C260 VDD2.n17 VSUBS 0.027759f
C261 VDD2.n18 VSUBS 0.014916f
C262 VDD2.n19 VSUBS 0.035257f
C263 VDD2.n20 VSUBS 0.015794f
C264 VDD2.n21 VSUBS 0.027759f
C265 VDD2.n22 VSUBS 0.014916f
C266 VDD2.n23 VSUBS 0.035257f
C267 VDD2.n24 VSUBS 0.015794f
C268 VDD2.n25 VSUBS 0.027759f
C269 VDD2.n26 VSUBS 0.014916f
C270 VDD2.n27 VSUBS 0.035257f
C271 VDD2.n28 VSUBS 0.015794f
C272 VDD2.n29 VSUBS 0.027759f
C273 VDD2.n30 VSUBS 0.014916f
C274 VDD2.n31 VSUBS 0.035257f
C275 VDD2.n32 VSUBS 0.015794f
C276 VDD2.n33 VSUBS 0.313379f
C277 VDD2.t0 VSUBS 0.076683f
C278 VDD2.n34 VSUBS 0.026443f
C279 VDD2.n35 VSUBS 0.026522f
C280 VDD2.n36 VSUBS 0.014916f
C281 VDD2.n37 VSUBS 2.28217f
C282 VDD2.n38 VSUBS 0.027759f
C283 VDD2.n39 VSUBS 0.014916f
C284 VDD2.n40 VSUBS 0.015794f
C285 VDD2.n41 VSUBS 0.035257f
C286 VDD2.n42 VSUBS 0.035257f
C287 VDD2.n43 VSUBS 0.015794f
C288 VDD2.n44 VSUBS 0.014916f
C289 VDD2.n45 VSUBS 0.027759f
C290 VDD2.n46 VSUBS 0.027759f
C291 VDD2.n47 VSUBS 0.014916f
C292 VDD2.n48 VSUBS 0.015794f
C293 VDD2.n49 VSUBS 0.035257f
C294 VDD2.n50 VSUBS 0.035257f
C295 VDD2.n51 VSUBS 0.035257f
C296 VDD2.n52 VSUBS 0.015794f
C297 VDD2.n53 VSUBS 0.014916f
C298 VDD2.n54 VSUBS 0.027759f
C299 VDD2.n55 VSUBS 0.027759f
C300 VDD2.n56 VSUBS 0.014916f
C301 VDD2.n57 VSUBS 0.015355f
C302 VDD2.n58 VSUBS 0.015355f
C303 VDD2.n59 VSUBS 0.035257f
C304 VDD2.n60 VSUBS 0.035257f
C305 VDD2.n61 VSUBS 0.015794f
C306 VDD2.n62 VSUBS 0.014916f
C307 VDD2.n63 VSUBS 0.027759f
C308 VDD2.n64 VSUBS 0.027759f
C309 VDD2.n65 VSUBS 0.014916f
C310 VDD2.n66 VSUBS 0.015794f
C311 VDD2.n67 VSUBS 0.035257f
C312 VDD2.n68 VSUBS 0.035257f
C313 VDD2.n69 VSUBS 0.015794f
C314 VDD2.n70 VSUBS 0.014916f
C315 VDD2.n71 VSUBS 0.027759f
C316 VDD2.n72 VSUBS 0.027759f
C317 VDD2.n73 VSUBS 0.014916f
C318 VDD2.n74 VSUBS 0.015794f
C319 VDD2.n75 VSUBS 0.035257f
C320 VDD2.n76 VSUBS 0.035257f
C321 VDD2.n77 VSUBS 0.015794f
C322 VDD2.n78 VSUBS 0.014916f
C323 VDD2.n79 VSUBS 0.027759f
C324 VDD2.n80 VSUBS 0.027759f
C325 VDD2.n81 VSUBS 0.014916f
C326 VDD2.n82 VSUBS 0.015794f
C327 VDD2.n83 VSUBS 0.035257f
C328 VDD2.n84 VSUBS 0.035257f
C329 VDD2.n85 VSUBS 0.015794f
C330 VDD2.n86 VSUBS 0.014916f
C331 VDD2.n87 VSUBS 0.027759f
C332 VDD2.n88 VSUBS 0.027759f
C333 VDD2.n89 VSUBS 0.014916f
C334 VDD2.n90 VSUBS 0.015794f
C335 VDD2.n91 VSUBS 0.035257f
C336 VDD2.n92 VSUBS 0.035257f
C337 VDD2.n93 VSUBS 0.015794f
C338 VDD2.n94 VSUBS 0.014916f
C339 VDD2.n95 VSUBS 0.027759f
C340 VDD2.n96 VSUBS 0.027759f
C341 VDD2.n97 VSUBS 0.014916f
C342 VDD2.n98 VSUBS 0.015794f
C343 VDD2.n99 VSUBS 0.035257f
C344 VDD2.n100 VSUBS 0.08963f
C345 VDD2.n101 VSUBS 0.015794f
C346 VDD2.n102 VSUBS 0.029292f
C347 VDD2.n103 VSUBS 0.072885f
C348 VDD2.n104 VSUBS 1.01635f
C349 VDD2.n105 VSUBS 0.031029f
C350 VDD2.n106 VSUBS 0.027759f
C351 VDD2.n107 VSUBS 0.014916f
C352 VDD2.n108 VSUBS 0.035257f
C353 VDD2.n109 VSUBS 0.015794f
C354 VDD2.n110 VSUBS 0.027759f
C355 VDD2.n111 VSUBS 0.014916f
C356 VDD2.n112 VSUBS 0.035257f
C357 VDD2.n113 VSUBS 0.015794f
C358 VDD2.n114 VSUBS 0.027759f
C359 VDD2.n115 VSUBS 0.014916f
C360 VDD2.n116 VSUBS 0.035257f
C361 VDD2.n117 VSUBS 0.015794f
C362 VDD2.n118 VSUBS 0.027759f
C363 VDD2.n119 VSUBS 0.014916f
C364 VDD2.n120 VSUBS 0.035257f
C365 VDD2.n121 VSUBS 0.015794f
C366 VDD2.n122 VSUBS 0.027759f
C367 VDD2.n123 VSUBS 0.014916f
C368 VDD2.n124 VSUBS 0.035257f
C369 VDD2.n125 VSUBS 0.015794f
C370 VDD2.n126 VSUBS 0.027759f
C371 VDD2.n127 VSUBS 0.014916f
C372 VDD2.n128 VSUBS 0.035257f
C373 VDD2.n129 VSUBS 0.015794f
C374 VDD2.n130 VSUBS 0.027759f
C375 VDD2.n131 VSUBS 0.014916f
C376 VDD2.n132 VSUBS 0.035257f
C377 VDD2.n133 VSUBS 0.035257f
C378 VDD2.n134 VSUBS 0.015794f
C379 VDD2.n135 VSUBS 0.027759f
C380 VDD2.n136 VSUBS 0.014916f
C381 VDD2.n137 VSUBS 0.035257f
C382 VDD2.n138 VSUBS 0.015794f
C383 VDD2.n139 VSUBS 0.313379f
C384 VDD2.t1 VSUBS 0.076683f
C385 VDD2.n140 VSUBS 0.026443f
C386 VDD2.n141 VSUBS 0.026522f
C387 VDD2.n142 VSUBS 0.014916f
C388 VDD2.n143 VSUBS 2.28217f
C389 VDD2.n144 VSUBS 0.027759f
C390 VDD2.n145 VSUBS 0.014916f
C391 VDD2.n146 VSUBS 0.015794f
C392 VDD2.n147 VSUBS 0.035257f
C393 VDD2.n148 VSUBS 0.035257f
C394 VDD2.n149 VSUBS 0.015794f
C395 VDD2.n150 VSUBS 0.014916f
C396 VDD2.n151 VSUBS 0.027759f
C397 VDD2.n152 VSUBS 0.027759f
C398 VDD2.n153 VSUBS 0.014916f
C399 VDD2.n154 VSUBS 0.015794f
C400 VDD2.n155 VSUBS 0.035257f
C401 VDD2.n156 VSUBS 0.035257f
C402 VDD2.n157 VSUBS 0.015794f
C403 VDD2.n158 VSUBS 0.014916f
C404 VDD2.n159 VSUBS 0.027759f
C405 VDD2.n160 VSUBS 0.027759f
C406 VDD2.n161 VSUBS 0.014916f
C407 VDD2.n162 VSUBS 0.015355f
C408 VDD2.n163 VSUBS 0.015355f
C409 VDD2.n164 VSUBS 0.035257f
C410 VDD2.n165 VSUBS 0.035257f
C411 VDD2.n166 VSUBS 0.015794f
C412 VDD2.n167 VSUBS 0.014916f
C413 VDD2.n168 VSUBS 0.027759f
C414 VDD2.n169 VSUBS 0.027759f
C415 VDD2.n170 VSUBS 0.014916f
C416 VDD2.n171 VSUBS 0.015794f
C417 VDD2.n172 VSUBS 0.035257f
C418 VDD2.n173 VSUBS 0.035257f
C419 VDD2.n174 VSUBS 0.015794f
C420 VDD2.n175 VSUBS 0.014916f
C421 VDD2.n176 VSUBS 0.027759f
C422 VDD2.n177 VSUBS 0.027759f
C423 VDD2.n178 VSUBS 0.014916f
C424 VDD2.n179 VSUBS 0.015794f
C425 VDD2.n180 VSUBS 0.035257f
C426 VDD2.n181 VSUBS 0.035257f
C427 VDD2.n182 VSUBS 0.015794f
C428 VDD2.n183 VSUBS 0.014916f
C429 VDD2.n184 VSUBS 0.027759f
C430 VDD2.n185 VSUBS 0.027759f
C431 VDD2.n186 VSUBS 0.014916f
C432 VDD2.n187 VSUBS 0.015794f
C433 VDD2.n188 VSUBS 0.035257f
C434 VDD2.n189 VSUBS 0.035257f
C435 VDD2.n190 VSUBS 0.015794f
C436 VDD2.n191 VSUBS 0.014916f
C437 VDD2.n192 VSUBS 0.027759f
C438 VDD2.n193 VSUBS 0.027759f
C439 VDD2.n194 VSUBS 0.014916f
C440 VDD2.n195 VSUBS 0.015794f
C441 VDD2.n196 VSUBS 0.035257f
C442 VDD2.n197 VSUBS 0.035257f
C443 VDD2.n198 VSUBS 0.015794f
C444 VDD2.n199 VSUBS 0.014916f
C445 VDD2.n200 VSUBS 0.027759f
C446 VDD2.n201 VSUBS 0.027759f
C447 VDD2.n202 VSUBS 0.014916f
C448 VDD2.n203 VSUBS 0.015794f
C449 VDD2.n204 VSUBS 0.035257f
C450 VDD2.n205 VSUBS 0.08963f
C451 VDD2.n206 VSUBS 0.015794f
C452 VDD2.n207 VSUBS 0.029292f
C453 VDD2.n208 VSUBS 0.072885f
C454 VDD2.n209 VSUBS 0.08886f
C455 VDD2.n210 VSUBS 4.0236f
C456 VTAIL.n0 VSUBS 0.03086f
C457 VTAIL.n1 VSUBS 0.027608f
C458 VTAIL.n2 VSUBS 0.014835f
C459 VTAIL.n3 VSUBS 0.035065f
C460 VTAIL.n4 VSUBS 0.015708f
C461 VTAIL.n5 VSUBS 0.027608f
C462 VTAIL.n6 VSUBS 0.014835f
C463 VTAIL.n7 VSUBS 0.035065f
C464 VTAIL.n8 VSUBS 0.015708f
C465 VTAIL.n9 VSUBS 0.027608f
C466 VTAIL.n10 VSUBS 0.014835f
C467 VTAIL.n11 VSUBS 0.035065f
C468 VTAIL.n12 VSUBS 0.015708f
C469 VTAIL.n13 VSUBS 0.027608f
C470 VTAIL.n14 VSUBS 0.014835f
C471 VTAIL.n15 VSUBS 0.035065f
C472 VTAIL.n16 VSUBS 0.015708f
C473 VTAIL.n17 VSUBS 0.027608f
C474 VTAIL.n18 VSUBS 0.014835f
C475 VTAIL.n19 VSUBS 0.035065f
C476 VTAIL.n20 VSUBS 0.015708f
C477 VTAIL.n21 VSUBS 0.027608f
C478 VTAIL.n22 VSUBS 0.014835f
C479 VTAIL.n23 VSUBS 0.035065f
C480 VTAIL.n24 VSUBS 0.015708f
C481 VTAIL.n25 VSUBS 0.027608f
C482 VTAIL.n26 VSUBS 0.014835f
C483 VTAIL.n27 VSUBS 0.035065f
C484 VTAIL.n28 VSUBS 0.015708f
C485 VTAIL.n29 VSUBS 0.027608f
C486 VTAIL.n30 VSUBS 0.014835f
C487 VTAIL.n31 VSUBS 0.035065f
C488 VTAIL.n32 VSUBS 0.015708f
C489 VTAIL.n33 VSUBS 0.311677f
C490 VTAIL.t1 VSUBS 0.076266f
C491 VTAIL.n34 VSUBS 0.026299f
C492 VTAIL.n35 VSUBS 0.026378f
C493 VTAIL.n36 VSUBS 0.014835f
C494 VTAIL.n37 VSUBS 2.26977f
C495 VTAIL.n38 VSUBS 0.027608f
C496 VTAIL.n39 VSUBS 0.014835f
C497 VTAIL.n40 VSUBS 0.015708f
C498 VTAIL.n41 VSUBS 0.035065f
C499 VTAIL.n42 VSUBS 0.035065f
C500 VTAIL.n43 VSUBS 0.015708f
C501 VTAIL.n44 VSUBS 0.014835f
C502 VTAIL.n45 VSUBS 0.027608f
C503 VTAIL.n46 VSUBS 0.027608f
C504 VTAIL.n47 VSUBS 0.014835f
C505 VTAIL.n48 VSUBS 0.015708f
C506 VTAIL.n49 VSUBS 0.035065f
C507 VTAIL.n50 VSUBS 0.035065f
C508 VTAIL.n51 VSUBS 0.035065f
C509 VTAIL.n52 VSUBS 0.015708f
C510 VTAIL.n53 VSUBS 0.014835f
C511 VTAIL.n54 VSUBS 0.027608f
C512 VTAIL.n55 VSUBS 0.027608f
C513 VTAIL.n56 VSUBS 0.014835f
C514 VTAIL.n57 VSUBS 0.015272f
C515 VTAIL.n58 VSUBS 0.015272f
C516 VTAIL.n59 VSUBS 0.035065f
C517 VTAIL.n60 VSUBS 0.035065f
C518 VTAIL.n61 VSUBS 0.015708f
C519 VTAIL.n62 VSUBS 0.014835f
C520 VTAIL.n63 VSUBS 0.027608f
C521 VTAIL.n64 VSUBS 0.027608f
C522 VTAIL.n65 VSUBS 0.014835f
C523 VTAIL.n66 VSUBS 0.015708f
C524 VTAIL.n67 VSUBS 0.035065f
C525 VTAIL.n68 VSUBS 0.035065f
C526 VTAIL.n69 VSUBS 0.015708f
C527 VTAIL.n70 VSUBS 0.014835f
C528 VTAIL.n71 VSUBS 0.027608f
C529 VTAIL.n72 VSUBS 0.027608f
C530 VTAIL.n73 VSUBS 0.014835f
C531 VTAIL.n74 VSUBS 0.015708f
C532 VTAIL.n75 VSUBS 0.035065f
C533 VTAIL.n76 VSUBS 0.035065f
C534 VTAIL.n77 VSUBS 0.015708f
C535 VTAIL.n78 VSUBS 0.014835f
C536 VTAIL.n79 VSUBS 0.027608f
C537 VTAIL.n80 VSUBS 0.027608f
C538 VTAIL.n81 VSUBS 0.014835f
C539 VTAIL.n82 VSUBS 0.015708f
C540 VTAIL.n83 VSUBS 0.035065f
C541 VTAIL.n84 VSUBS 0.035065f
C542 VTAIL.n85 VSUBS 0.015708f
C543 VTAIL.n86 VSUBS 0.014835f
C544 VTAIL.n87 VSUBS 0.027608f
C545 VTAIL.n88 VSUBS 0.027608f
C546 VTAIL.n89 VSUBS 0.014835f
C547 VTAIL.n90 VSUBS 0.015708f
C548 VTAIL.n91 VSUBS 0.035065f
C549 VTAIL.n92 VSUBS 0.035065f
C550 VTAIL.n93 VSUBS 0.015708f
C551 VTAIL.n94 VSUBS 0.014835f
C552 VTAIL.n95 VSUBS 0.027608f
C553 VTAIL.n96 VSUBS 0.027608f
C554 VTAIL.n97 VSUBS 0.014835f
C555 VTAIL.n98 VSUBS 0.015708f
C556 VTAIL.n99 VSUBS 0.035065f
C557 VTAIL.n100 VSUBS 0.089143f
C558 VTAIL.n101 VSUBS 0.015708f
C559 VTAIL.n102 VSUBS 0.029133f
C560 VTAIL.n103 VSUBS 0.072489f
C561 VTAIL.n104 VSUBS 0.069374f
C562 VTAIL.n105 VSUBS 2.23618f
C563 VTAIL.n106 VSUBS 0.03086f
C564 VTAIL.n107 VSUBS 0.027608f
C565 VTAIL.n108 VSUBS 0.014835f
C566 VTAIL.n109 VSUBS 0.035065f
C567 VTAIL.n110 VSUBS 0.015708f
C568 VTAIL.n111 VSUBS 0.027608f
C569 VTAIL.n112 VSUBS 0.014835f
C570 VTAIL.n113 VSUBS 0.035065f
C571 VTAIL.n114 VSUBS 0.015708f
C572 VTAIL.n115 VSUBS 0.027608f
C573 VTAIL.n116 VSUBS 0.014835f
C574 VTAIL.n117 VSUBS 0.035065f
C575 VTAIL.n118 VSUBS 0.015708f
C576 VTAIL.n119 VSUBS 0.027608f
C577 VTAIL.n120 VSUBS 0.014835f
C578 VTAIL.n121 VSUBS 0.035065f
C579 VTAIL.n122 VSUBS 0.015708f
C580 VTAIL.n123 VSUBS 0.027608f
C581 VTAIL.n124 VSUBS 0.014835f
C582 VTAIL.n125 VSUBS 0.035065f
C583 VTAIL.n126 VSUBS 0.015708f
C584 VTAIL.n127 VSUBS 0.027608f
C585 VTAIL.n128 VSUBS 0.014835f
C586 VTAIL.n129 VSUBS 0.035065f
C587 VTAIL.n130 VSUBS 0.015708f
C588 VTAIL.n131 VSUBS 0.027608f
C589 VTAIL.n132 VSUBS 0.014835f
C590 VTAIL.n133 VSUBS 0.035065f
C591 VTAIL.n134 VSUBS 0.035065f
C592 VTAIL.n135 VSUBS 0.015708f
C593 VTAIL.n136 VSUBS 0.027608f
C594 VTAIL.n137 VSUBS 0.014835f
C595 VTAIL.n138 VSUBS 0.035065f
C596 VTAIL.n139 VSUBS 0.015708f
C597 VTAIL.n140 VSUBS 0.311677f
C598 VTAIL.t2 VSUBS 0.076266f
C599 VTAIL.n141 VSUBS 0.026299f
C600 VTAIL.n142 VSUBS 0.026378f
C601 VTAIL.n143 VSUBS 0.014835f
C602 VTAIL.n144 VSUBS 2.26977f
C603 VTAIL.n145 VSUBS 0.027608f
C604 VTAIL.n146 VSUBS 0.014835f
C605 VTAIL.n147 VSUBS 0.015708f
C606 VTAIL.n148 VSUBS 0.035065f
C607 VTAIL.n149 VSUBS 0.035065f
C608 VTAIL.n150 VSUBS 0.015708f
C609 VTAIL.n151 VSUBS 0.014835f
C610 VTAIL.n152 VSUBS 0.027608f
C611 VTAIL.n153 VSUBS 0.027608f
C612 VTAIL.n154 VSUBS 0.014835f
C613 VTAIL.n155 VSUBS 0.015708f
C614 VTAIL.n156 VSUBS 0.035065f
C615 VTAIL.n157 VSUBS 0.035065f
C616 VTAIL.n158 VSUBS 0.015708f
C617 VTAIL.n159 VSUBS 0.014835f
C618 VTAIL.n160 VSUBS 0.027608f
C619 VTAIL.n161 VSUBS 0.027608f
C620 VTAIL.n162 VSUBS 0.014835f
C621 VTAIL.n163 VSUBS 0.015272f
C622 VTAIL.n164 VSUBS 0.015272f
C623 VTAIL.n165 VSUBS 0.035065f
C624 VTAIL.n166 VSUBS 0.035065f
C625 VTAIL.n167 VSUBS 0.015708f
C626 VTAIL.n168 VSUBS 0.014835f
C627 VTAIL.n169 VSUBS 0.027608f
C628 VTAIL.n170 VSUBS 0.027608f
C629 VTAIL.n171 VSUBS 0.014835f
C630 VTAIL.n172 VSUBS 0.015708f
C631 VTAIL.n173 VSUBS 0.035065f
C632 VTAIL.n174 VSUBS 0.035065f
C633 VTAIL.n175 VSUBS 0.015708f
C634 VTAIL.n176 VSUBS 0.014835f
C635 VTAIL.n177 VSUBS 0.027608f
C636 VTAIL.n178 VSUBS 0.027608f
C637 VTAIL.n179 VSUBS 0.014835f
C638 VTAIL.n180 VSUBS 0.015708f
C639 VTAIL.n181 VSUBS 0.035065f
C640 VTAIL.n182 VSUBS 0.035065f
C641 VTAIL.n183 VSUBS 0.015708f
C642 VTAIL.n184 VSUBS 0.014835f
C643 VTAIL.n185 VSUBS 0.027608f
C644 VTAIL.n186 VSUBS 0.027608f
C645 VTAIL.n187 VSUBS 0.014835f
C646 VTAIL.n188 VSUBS 0.015708f
C647 VTAIL.n189 VSUBS 0.035065f
C648 VTAIL.n190 VSUBS 0.035065f
C649 VTAIL.n191 VSUBS 0.015708f
C650 VTAIL.n192 VSUBS 0.014835f
C651 VTAIL.n193 VSUBS 0.027608f
C652 VTAIL.n194 VSUBS 0.027608f
C653 VTAIL.n195 VSUBS 0.014835f
C654 VTAIL.n196 VSUBS 0.015708f
C655 VTAIL.n197 VSUBS 0.035065f
C656 VTAIL.n198 VSUBS 0.035065f
C657 VTAIL.n199 VSUBS 0.015708f
C658 VTAIL.n200 VSUBS 0.014835f
C659 VTAIL.n201 VSUBS 0.027608f
C660 VTAIL.n202 VSUBS 0.027608f
C661 VTAIL.n203 VSUBS 0.014835f
C662 VTAIL.n204 VSUBS 0.015708f
C663 VTAIL.n205 VSUBS 0.035065f
C664 VTAIL.n206 VSUBS 0.089143f
C665 VTAIL.n207 VSUBS 0.015708f
C666 VTAIL.n208 VSUBS 0.029133f
C667 VTAIL.n209 VSUBS 0.072489f
C668 VTAIL.n210 VSUBS 0.069374f
C669 VTAIL.n211 VSUBS 2.26283f
C670 VTAIL.n212 VSUBS 0.03086f
C671 VTAIL.n213 VSUBS 0.027608f
C672 VTAIL.n214 VSUBS 0.014835f
C673 VTAIL.n215 VSUBS 0.035065f
C674 VTAIL.n216 VSUBS 0.015708f
C675 VTAIL.n217 VSUBS 0.027608f
C676 VTAIL.n218 VSUBS 0.014835f
C677 VTAIL.n219 VSUBS 0.035065f
C678 VTAIL.n220 VSUBS 0.015708f
C679 VTAIL.n221 VSUBS 0.027608f
C680 VTAIL.n222 VSUBS 0.014835f
C681 VTAIL.n223 VSUBS 0.035065f
C682 VTAIL.n224 VSUBS 0.015708f
C683 VTAIL.n225 VSUBS 0.027608f
C684 VTAIL.n226 VSUBS 0.014835f
C685 VTAIL.n227 VSUBS 0.035065f
C686 VTAIL.n228 VSUBS 0.015708f
C687 VTAIL.n229 VSUBS 0.027608f
C688 VTAIL.n230 VSUBS 0.014835f
C689 VTAIL.n231 VSUBS 0.035065f
C690 VTAIL.n232 VSUBS 0.015708f
C691 VTAIL.n233 VSUBS 0.027608f
C692 VTAIL.n234 VSUBS 0.014835f
C693 VTAIL.n235 VSUBS 0.035065f
C694 VTAIL.n236 VSUBS 0.015708f
C695 VTAIL.n237 VSUBS 0.027608f
C696 VTAIL.n238 VSUBS 0.014835f
C697 VTAIL.n239 VSUBS 0.035065f
C698 VTAIL.n240 VSUBS 0.035065f
C699 VTAIL.n241 VSUBS 0.015708f
C700 VTAIL.n242 VSUBS 0.027608f
C701 VTAIL.n243 VSUBS 0.014835f
C702 VTAIL.n244 VSUBS 0.035065f
C703 VTAIL.n245 VSUBS 0.015708f
C704 VTAIL.n246 VSUBS 0.311677f
C705 VTAIL.t0 VSUBS 0.076266f
C706 VTAIL.n247 VSUBS 0.026299f
C707 VTAIL.n248 VSUBS 0.026378f
C708 VTAIL.n249 VSUBS 0.014835f
C709 VTAIL.n250 VSUBS 2.26977f
C710 VTAIL.n251 VSUBS 0.027608f
C711 VTAIL.n252 VSUBS 0.014835f
C712 VTAIL.n253 VSUBS 0.015708f
C713 VTAIL.n254 VSUBS 0.035065f
C714 VTAIL.n255 VSUBS 0.035065f
C715 VTAIL.n256 VSUBS 0.015708f
C716 VTAIL.n257 VSUBS 0.014835f
C717 VTAIL.n258 VSUBS 0.027608f
C718 VTAIL.n259 VSUBS 0.027608f
C719 VTAIL.n260 VSUBS 0.014835f
C720 VTAIL.n261 VSUBS 0.015708f
C721 VTAIL.n262 VSUBS 0.035065f
C722 VTAIL.n263 VSUBS 0.035065f
C723 VTAIL.n264 VSUBS 0.015708f
C724 VTAIL.n265 VSUBS 0.014835f
C725 VTAIL.n266 VSUBS 0.027608f
C726 VTAIL.n267 VSUBS 0.027608f
C727 VTAIL.n268 VSUBS 0.014835f
C728 VTAIL.n269 VSUBS 0.015272f
C729 VTAIL.n270 VSUBS 0.015272f
C730 VTAIL.n271 VSUBS 0.035065f
C731 VTAIL.n272 VSUBS 0.035065f
C732 VTAIL.n273 VSUBS 0.015708f
C733 VTAIL.n274 VSUBS 0.014835f
C734 VTAIL.n275 VSUBS 0.027608f
C735 VTAIL.n276 VSUBS 0.027608f
C736 VTAIL.n277 VSUBS 0.014835f
C737 VTAIL.n278 VSUBS 0.015708f
C738 VTAIL.n279 VSUBS 0.035065f
C739 VTAIL.n280 VSUBS 0.035065f
C740 VTAIL.n281 VSUBS 0.015708f
C741 VTAIL.n282 VSUBS 0.014835f
C742 VTAIL.n283 VSUBS 0.027608f
C743 VTAIL.n284 VSUBS 0.027608f
C744 VTAIL.n285 VSUBS 0.014835f
C745 VTAIL.n286 VSUBS 0.015708f
C746 VTAIL.n287 VSUBS 0.035065f
C747 VTAIL.n288 VSUBS 0.035065f
C748 VTAIL.n289 VSUBS 0.015708f
C749 VTAIL.n290 VSUBS 0.014835f
C750 VTAIL.n291 VSUBS 0.027608f
C751 VTAIL.n292 VSUBS 0.027608f
C752 VTAIL.n293 VSUBS 0.014835f
C753 VTAIL.n294 VSUBS 0.015708f
C754 VTAIL.n295 VSUBS 0.035065f
C755 VTAIL.n296 VSUBS 0.035065f
C756 VTAIL.n297 VSUBS 0.015708f
C757 VTAIL.n298 VSUBS 0.014835f
C758 VTAIL.n299 VSUBS 0.027608f
C759 VTAIL.n300 VSUBS 0.027608f
C760 VTAIL.n301 VSUBS 0.014835f
C761 VTAIL.n302 VSUBS 0.015708f
C762 VTAIL.n303 VSUBS 0.035065f
C763 VTAIL.n304 VSUBS 0.035065f
C764 VTAIL.n305 VSUBS 0.015708f
C765 VTAIL.n306 VSUBS 0.014835f
C766 VTAIL.n307 VSUBS 0.027608f
C767 VTAIL.n308 VSUBS 0.027608f
C768 VTAIL.n309 VSUBS 0.014835f
C769 VTAIL.n310 VSUBS 0.015708f
C770 VTAIL.n311 VSUBS 0.035065f
C771 VTAIL.n312 VSUBS 0.089143f
C772 VTAIL.n313 VSUBS 0.015708f
C773 VTAIL.n314 VSUBS 0.029133f
C774 VTAIL.n315 VSUBS 0.072489f
C775 VTAIL.n316 VSUBS 0.069374f
C776 VTAIL.n317 VSUBS 2.13553f
C777 VTAIL.n318 VSUBS 0.03086f
C778 VTAIL.n319 VSUBS 0.027608f
C779 VTAIL.n320 VSUBS 0.014835f
C780 VTAIL.n321 VSUBS 0.035065f
C781 VTAIL.n322 VSUBS 0.015708f
C782 VTAIL.n323 VSUBS 0.027608f
C783 VTAIL.n324 VSUBS 0.014835f
C784 VTAIL.n325 VSUBS 0.035065f
C785 VTAIL.n326 VSUBS 0.015708f
C786 VTAIL.n327 VSUBS 0.027608f
C787 VTAIL.n328 VSUBS 0.014835f
C788 VTAIL.n329 VSUBS 0.035065f
C789 VTAIL.n330 VSUBS 0.015708f
C790 VTAIL.n331 VSUBS 0.027608f
C791 VTAIL.n332 VSUBS 0.014835f
C792 VTAIL.n333 VSUBS 0.035065f
C793 VTAIL.n334 VSUBS 0.015708f
C794 VTAIL.n335 VSUBS 0.027608f
C795 VTAIL.n336 VSUBS 0.014835f
C796 VTAIL.n337 VSUBS 0.035065f
C797 VTAIL.n338 VSUBS 0.015708f
C798 VTAIL.n339 VSUBS 0.027608f
C799 VTAIL.n340 VSUBS 0.014835f
C800 VTAIL.n341 VSUBS 0.035065f
C801 VTAIL.n342 VSUBS 0.015708f
C802 VTAIL.n343 VSUBS 0.027608f
C803 VTAIL.n344 VSUBS 0.014835f
C804 VTAIL.n345 VSUBS 0.035065f
C805 VTAIL.n346 VSUBS 0.015708f
C806 VTAIL.n347 VSUBS 0.027608f
C807 VTAIL.n348 VSUBS 0.014835f
C808 VTAIL.n349 VSUBS 0.035065f
C809 VTAIL.n350 VSUBS 0.015708f
C810 VTAIL.n351 VSUBS 0.311677f
C811 VTAIL.t3 VSUBS 0.076266f
C812 VTAIL.n352 VSUBS 0.026299f
C813 VTAIL.n353 VSUBS 0.026378f
C814 VTAIL.n354 VSUBS 0.014835f
C815 VTAIL.n355 VSUBS 2.26977f
C816 VTAIL.n356 VSUBS 0.027608f
C817 VTAIL.n357 VSUBS 0.014835f
C818 VTAIL.n358 VSUBS 0.015708f
C819 VTAIL.n359 VSUBS 0.035065f
C820 VTAIL.n360 VSUBS 0.035065f
C821 VTAIL.n361 VSUBS 0.015708f
C822 VTAIL.n362 VSUBS 0.014835f
C823 VTAIL.n363 VSUBS 0.027608f
C824 VTAIL.n364 VSUBS 0.027608f
C825 VTAIL.n365 VSUBS 0.014835f
C826 VTAIL.n366 VSUBS 0.015708f
C827 VTAIL.n367 VSUBS 0.035065f
C828 VTAIL.n368 VSUBS 0.035065f
C829 VTAIL.n369 VSUBS 0.035065f
C830 VTAIL.n370 VSUBS 0.015708f
C831 VTAIL.n371 VSUBS 0.014835f
C832 VTAIL.n372 VSUBS 0.027608f
C833 VTAIL.n373 VSUBS 0.027608f
C834 VTAIL.n374 VSUBS 0.014835f
C835 VTAIL.n375 VSUBS 0.015272f
C836 VTAIL.n376 VSUBS 0.015272f
C837 VTAIL.n377 VSUBS 0.035065f
C838 VTAIL.n378 VSUBS 0.035065f
C839 VTAIL.n379 VSUBS 0.015708f
C840 VTAIL.n380 VSUBS 0.014835f
C841 VTAIL.n381 VSUBS 0.027608f
C842 VTAIL.n382 VSUBS 0.027608f
C843 VTAIL.n383 VSUBS 0.014835f
C844 VTAIL.n384 VSUBS 0.015708f
C845 VTAIL.n385 VSUBS 0.035065f
C846 VTAIL.n386 VSUBS 0.035065f
C847 VTAIL.n387 VSUBS 0.015708f
C848 VTAIL.n388 VSUBS 0.014835f
C849 VTAIL.n389 VSUBS 0.027608f
C850 VTAIL.n390 VSUBS 0.027608f
C851 VTAIL.n391 VSUBS 0.014835f
C852 VTAIL.n392 VSUBS 0.015708f
C853 VTAIL.n393 VSUBS 0.035065f
C854 VTAIL.n394 VSUBS 0.035065f
C855 VTAIL.n395 VSUBS 0.015708f
C856 VTAIL.n396 VSUBS 0.014835f
C857 VTAIL.n397 VSUBS 0.027608f
C858 VTAIL.n398 VSUBS 0.027608f
C859 VTAIL.n399 VSUBS 0.014835f
C860 VTAIL.n400 VSUBS 0.015708f
C861 VTAIL.n401 VSUBS 0.035065f
C862 VTAIL.n402 VSUBS 0.035065f
C863 VTAIL.n403 VSUBS 0.015708f
C864 VTAIL.n404 VSUBS 0.014835f
C865 VTAIL.n405 VSUBS 0.027608f
C866 VTAIL.n406 VSUBS 0.027608f
C867 VTAIL.n407 VSUBS 0.014835f
C868 VTAIL.n408 VSUBS 0.015708f
C869 VTAIL.n409 VSUBS 0.035065f
C870 VTAIL.n410 VSUBS 0.035065f
C871 VTAIL.n411 VSUBS 0.015708f
C872 VTAIL.n412 VSUBS 0.014835f
C873 VTAIL.n413 VSUBS 0.027608f
C874 VTAIL.n414 VSUBS 0.027608f
C875 VTAIL.n415 VSUBS 0.014835f
C876 VTAIL.n416 VSUBS 0.015708f
C877 VTAIL.n417 VSUBS 0.035065f
C878 VTAIL.n418 VSUBS 0.089143f
C879 VTAIL.n419 VSUBS 0.015708f
C880 VTAIL.n420 VSUBS 0.029133f
C881 VTAIL.n421 VSUBS 0.072489f
C882 VTAIL.n422 VSUBS 0.069374f
C883 VTAIL.n423 VSUBS 2.05673f
C884 VN.t1 VSUBS 3.98863f
C885 VN.t0 VSUBS 4.3333f
C886 B.n0 VSUBS 0.005031f
C887 B.n1 VSUBS 0.005031f
C888 B.n2 VSUBS 0.007957f
C889 B.n3 VSUBS 0.007957f
C890 B.n4 VSUBS 0.007957f
C891 B.n5 VSUBS 0.007957f
C892 B.n6 VSUBS 0.007957f
C893 B.n7 VSUBS 0.007957f
C894 B.n8 VSUBS 0.007957f
C895 B.n9 VSUBS 0.007957f
C896 B.n10 VSUBS 0.007957f
C897 B.n11 VSUBS 0.018754f
C898 B.n12 VSUBS 0.007957f
C899 B.n13 VSUBS 0.007957f
C900 B.n14 VSUBS 0.007957f
C901 B.n15 VSUBS 0.007957f
C902 B.n16 VSUBS 0.007957f
C903 B.n17 VSUBS 0.007957f
C904 B.n18 VSUBS 0.007957f
C905 B.n19 VSUBS 0.007957f
C906 B.n20 VSUBS 0.007957f
C907 B.n21 VSUBS 0.007957f
C908 B.n22 VSUBS 0.007957f
C909 B.n23 VSUBS 0.007957f
C910 B.n24 VSUBS 0.007957f
C911 B.n25 VSUBS 0.007957f
C912 B.n26 VSUBS 0.007957f
C913 B.n27 VSUBS 0.007957f
C914 B.n28 VSUBS 0.007957f
C915 B.n29 VSUBS 0.007957f
C916 B.n30 VSUBS 0.007957f
C917 B.n31 VSUBS 0.007957f
C918 B.n32 VSUBS 0.007957f
C919 B.n33 VSUBS 0.007957f
C920 B.n34 VSUBS 0.007957f
C921 B.n35 VSUBS 0.007957f
C922 B.n36 VSUBS 0.007957f
C923 B.n37 VSUBS 0.007957f
C924 B.n38 VSUBS 0.007957f
C925 B.n39 VSUBS 0.007957f
C926 B.n40 VSUBS 0.007957f
C927 B.n41 VSUBS 0.007957f
C928 B.n42 VSUBS 0.007957f
C929 B.n43 VSUBS 0.007957f
C930 B.t5 VSUBS 0.441938f
C931 B.t4 VSUBS 0.464264f
C932 B.t3 VSUBS 1.23853f
C933 B.n44 VSUBS 0.622209f
C934 B.n45 VSUBS 0.388466f
C935 B.n46 VSUBS 0.007957f
C936 B.n47 VSUBS 0.007957f
C937 B.n48 VSUBS 0.007957f
C938 B.n49 VSUBS 0.007957f
C939 B.t11 VSUBS 0.441942f
C940 B.t10 VSUBS 0.464268f
C941 B.t9 VSUBS 1.23853f
C942 B.n50 VSUBS 0.622206f
C943 B.n51 VSUBS 0.388461f
C944 B.n52 VSUBS 0.007957f
C945 B.n53 VSUBS 0.007957f
C946 B.n54 VSUBS 0.007957f
C947 B.n55 VSUBS 0.007957f
C948 B.n56 VSUBS 0.007957f
C949 B.n57 VSUBS 0.007957f
C950 B.n58 VSUBS 0.007957f
C951 B.n59 VSUBS 0.007957f
C952 B.n60 VSUBS 0.007957f
C953 B.n61 VSUBS 0.007957f
C954 B.n62 VSUBS 0.007957f
C955 B.n63 VSUBS 0.007957f
C956 B.n64 VSUBS 0.007957f
C957 B.n65 VSUBS 0.007957f
C958 B.n66 VSUBS 0.007957f
C959 B.n67 VSUBS 0.007957f
C960 B.n68 VSUBS 0.007957f
C961 B.n69 VSUBS 0.007957f
C962 B.n70 VSUBS 0.007957f
C963 B.n71 VSUBS 0.007957f
C964 B.n72 VSUBS 0.007957f
C965 B.n73 VSUBS 0.007957f
C966 B.n74 VSUBS 0.007957f
C967 B.n75 VSUBS 0.007957f
C968 B.n76 VSUBS 0.007957f
C969 B.n77 VSUBS 0.007957f
C970 B.n78 VSUBS 0.007957f
C971 B.n79 VSUBS 0.007957f
C972 B.n80 VSUBS 0.007957f
C973 B.n81 VSUBS 0.007957f
C974 B.n82 VSUBS 0.007957f
C975 B.n83 VSUBS 0.018754f
C976 B.n84 VSUBS 0.007957f
C977 B.n85 VSUBS 0.007957f
C978 B.n86 VSUBS 0.007957f
C979 B.n87 VSUBS 0.007957f
C980 B.n88 VSUBS 0.007957f
C981 B.n89 VSUBS 0.007957f
C982 B.n90 VSUBS 0.007957f
C983 B.n91 VSUBS 0.007957f
C984 B.n92 VSUBS 0.007957f
C985 B.n93 VSUBS 0.007957f
C986 B.n94 VSUBS 0.007957f
C987 B.n95 VSUBS 0.007957f
C988 B.n96 VSUBS 0.007957f
C989 B.n97 VSUBS 0.007957f
C990 B.n98 VSUBS 0.007957f
C991 B.n99 VSUBS 0.007957f
C992 B.n100 VSUBS 0.007957f
C993 B.n101 VSUBS 0.007957f
C994 B.n102 VSUBS 0.018754f
C995 B.n103 VSUBS 0.007957f
C996 B.n104 VSUBS 0.007957f
C997 B.n105 VSUBS 0.007957f
C998 B.n106 VSUBS 0.007957f
C999 B.n107 VSUBS 0.007957f
C1000 B.n108 VSUBS 0.007957f
C1001 B.n109 VSUBS 0.007957f
C1002 B.n110 VSUBS 0.007957f
C1003 B.n111 VSUBS 0.007957f
C1004 B.n112 VSUBS 0.007957f
C1005 B.n113 VSUBS 0.007957f
C1006 B.n114 VSUBS 0.007957f
C1007 B.n115 VSUBS 0.007957f
C1008 B.n116 VSUBS 0.007957f
C1009 B.n117 VSUBS 0.007957f
C1010 B.n118 VSUBS 0.007957f
C1011 B.n119 VSUBS 0.007957f
C1012 B.n120 VSUBS 0.007957f
C1013 B.n121 VSUBS 0.007957f
C1014 B.n122 VSUBS 0.007957f
C1015 B.n123 VSUBS 0.007957f
C1016 B.n124 VSUBS 0.007957f
C1017 B.n125 VSUBS 0.007957f
C1018 B.n126 VSUBS 0.007957f
C1019 B.n127 VSUBS 0.007957f
C1020 B.n128 VSUBS 0.007957f
C1021 B.n129 VSUBS 0.007957f
C1022 B.n130 VSUBS 0.007957f
C1023 B.n131 VSUBS 0.007957f
C1024 B.n132 VSUBS 0.007957f
C1025 B.n133 VSUBS 0.007957f
C1026 B.t1 VSUBS 0.441942f
C1027 B.t2 VSUBS 0.464268f
C1028 B.t0 VSUBS 1.23853f
C1029 B.n134 VSUBS 0.622206f
C1030 B.n135 VSUBS 0.388461f
C1031 B.n136 VSUBS 0.018435f
C1032 B.n137 VSUBS 0.007957f
C1033 B.n138 VSUBS 0.007957f
C1034 B.n139 VSUBS 0.007957f
C1035 B.n140 VSUBS 0.007957f
C1036 B.n141 VSUBS 0.007957f
C1037 B.t7 VSUBS 0.441938f
C1038 B.t8 VSUBS 0.464264f
C1039 B.t6 VSUBS 1.23853f
C1040 B.n142 VSUBS 0.622209f
C1041 B.n143 VSUBS 0.388466f
C1042 B.n144 VSUBS 0.007957f
C1043 B.n145 VSUBS 0.007957f
C1044 B.n146 VSUBS 0.007957f
C1045 B.n147 VSUBS 0.007957f
C1046 B.n148 VSUBS 0.007957f
C1047 B.n149 VSUBS 0.007957f
C1048 B.n150 VSUBS 0.007957f
C1049 B.n151 VSUBS 0.007957f
C1050 B.n152 VSUBS 0.007957f
C1051 B.n153 VSUBS 0.007957f
C1052 B.n154 VSUBS 0.007957f
C1053 B.n155 VSUBS 0.007957f
C1054 B.n156 VSUBS 0.007957f
C1055 B.n157 VSUBS 0.007957f
C1056 B.n158 VSUBS 0.007957f
C1057 B.n159 VSUBS 0.007957f
C1058 B.n160 VSUBS 0.007957f
C1059 B.n161 VSUBS 0.007957f
C1060 B.n162 VSUBS 0.007957f
C1061 B.n163 VSUBS 0.007957f
C1062 B.n164 VSUBS 0.007957f
C1063 B.n165 VSUBS 0.007957f
C1064 B.n166 VSUBS 0.007957f
C1065 B.n167 VSUBS 0.007957f
C1066 B.n168 VSUBS 0.007957f
C1067 B.n169 VSUBS 0.007957f
C1068 B.n170 VSUBS 0.007957f
C1069 B.n171 VSUBS 0.007957f
C1070 B.n172 VSUBS 0.007957f
C1071 B.n173 VSUBS 0.007957f
C1072 B.n174 VSUBS 0.007957f
C1073 B.n175 VSUBS 0.018221f
C1074 B.n176 VSUBS 0.007957f
C1075 B.n177 VSUBS 0.007957f
C1076 B.n178 VSUBS 0.007957f
C1077 B.n179 VSUBS 0.007957f
C1078 B.n180 VSUBS 0.007957f
C1079 B.n181 VSUBS 0.007957f
C1080 B.n182 VSUBS 0.007957f
C1081 B.n183 VSUBS 0.007957f
C1082 B.n184 VSUBS 0.007957f
C1083 B.n185 VSUBS 0.007957f
C1084 B.n186 VSUBS 0.007957f
C1085 B.n187 VSUBS 0.007957f
C1086 B.n188 VSUBS 0.007957f
C1087 B.n189 VSUBS 0.007957f
C1088 B.n190 VSUBS 0.007957f
C1089 B.n191 VSUBS 0.007957f
C1090 B.n192 VSUBS 0.007957f
C1091 B.n193 VSUBS 0.007957f
C1092 B.n194 VSUBS 0.007957f
C1093 B.n195 VSUBS 0.007957f
C1094 B.n196 VSUBS 0.007957f
C1095 B.n197 VSUBS 0.007957f
C1096 B.n198 VSUBS 0.007957f
C1097 B.n199 VSUBS 0.007957f
C1098 B.n200 VSUBS 0.007957f
C1099 B.n201 VSUBS 0.007957f
C1100 B.n202 VSUBS 0.007957f
C1101 B.n203 VSUBS 0.007957f
C1102 B.n204 VSUBS 0.007957f
C1103 B.n205 VSUBS 0.007957f
C1104 B.n206 VSUBS 0.007957f
C1105 B.n207 VSUBS 0.007957f
C1106 B.n208 VSUBS 0.018221f
C1107 B.n209 VSUBS 0.018754f
C1108 B.n210 VSUBS 0.018754f
C1109 B.n211 VSUBS 0.007957f
C1110 B.n212 VSUBS 0.007957f
C1111 B.n213 VSUBS 0.007957f
C1112 B.n214 VSUBS 0.007957f
C1113 B.n215 VSUBS 0.007957f
C1114 B.n216 VSUBS 0.007957f
C1115 B.n217 VSUBS 0.007957f
C1116 B.n218 VSUBS 0.007957f
C1117 B.n219 VSUBS 0.007957f
C1118 B.n220 VSUBS 0.007957f
C1119 B.n221 VSUBS 0.007957f
C1120 B.n222 VSUBS 0.007957f
C1121 B.n223 VSUBS 0.007957f
C1122 B.n224 VSUBS 0.007957f
C1123 B.n225 VSUBS 0.007957f
C1124 B.n226 VSUBS 0.007957f
C1125 B.n227 VSUBS 0.007957f
C1126 B.n228 VSUBS 0.007957f
C1127 B.n229 VSUBS 0.007957f
C1128 B.n230 VSUBS 0.007957f
C1129 B.n231 VSUBS 0.007957f
C1130 B.n232 VSUBS 0.007957f
C1131 B.n233 VSUBS 0.007957f
C1132 B.n234 VSUBS 0.007957f
C1133 B.n235 VSUBS 0.007957f
C1134 B.n236 VSUBS 0.007957f
C1135 B.n237 VSUBS 0.007957f
C1136 B.n238 VSUBS 0.007957f
C1137 B.n239 VSUBS 0.007957f
C1138 B.n240 VSUBS 0.007957f
C1139 B.n241 VSUBS 0.007957f
C1140 B.n242 VSUBS 0.007957f
C1141 B.n243 VSUBS 0.007957f
C1142 B.n244 VSUBS 0.007957f
C1143 B.n245 VSUBS 0.007957f
C1144 B.n246 VSUBS 0.007957f
C1145 B.n247 VSUBS 0.007957f
C1146 B.n248 VSUBS 0.007957f
C1147 B.n249 VSUBS 0.007957f
C1148 B.n250 VSUBS 0.007957f
C1149 B.n251 VSUBS 0.007957f
C1150 B.n252 VSUBS 0.007957f
C1151 B.n253 VSUBS 0.007957f
C1152 B.n254 VSUBS 0.007957f
C1153 B.n255 VSUBS 0.007957f
C1154 B.n256 VSUBS 0.007957f
C1155 B.n257 VSUBS 0.007957f
C1156 B.n258 VSUBS 0.007957f
C1157 B.n259 VSUBS 0.007957f
C1158 B.n260 VSUBS 0.007957f
C1159 B.n261 VSUBS 0.007957f
C1160 B.n262 VSUBS 0.007957f
C1161 B.n263 VSUBS 0.007957f
C1162 B.n264 VSUBS 0.007957f
C1163 B.n265 VSUBS 0.007957f
C1164 B.n266 VSUBS 0.007957f
C1165 B.n267 VSUBS 0.007957f
C1166 B.n268 VSUBS 0.007957f
C1167 B.n269 VSUBS 0.007957f
C1168 B.n270 VSUBS 0.007957f
C1169 B.n271 VSUBS 0.007957f
C1170 B.n272 VSUBS 0.007957f
C1171 B.n273 VSUBS 0.007957f
C1172 B.n274 VSUBS 0.007957f
C1173 B.n275 VSUBS 0.007957f
C1174 B.n276 VSUBS 0.007957f
C1175 B.n277 VSUBS 0.007957f
C1176 B.n278 VSUBS 0.007957f
C1177 B.n279 VSUBS 0.007957f
C1178 B.n280 VSUBS 0.007957f
C1179 B.n281 VSUBS 0.007957f
C1180 B.n282 VSUBS 0.007957f
C1181 B.n283 VSUBS 0.007957f
C1182 B.n284 VSUBS 0.007957f
C1183 B.n285 VSUBS 0.007957f
C1184 B.n286 VSUBS 0.007957f
C1185 B.n287 VSUBS 0.007957f
C1186 B.n288 VSUBS 0.007957f
C1187 B.n289 VSUBS 0.007957f
C1188 B.n290 VSUBS 0.007957f
C1189 B.n291 VSUBS 0.007957f
C1190 B.n292 VSUBS 0.007957f
C1191 B.n293 VSUBS 0.007957f
C1192 B.n294 VSUBS 0.007957f
C1193 B.n295 VSUBS 0.007957f
C1194 B.n296 VSUBS 0.007957f
C1195 B.n297 VSUBS 0.007957f
C1196 B.n298 VSUBS 0.007957f
C1197 B.n299 VSUBS 0.007957f
C1198 B.n300 VSUBS 0.007957f
C1199 B.n301 VSUBS 0.007957f
C1200 B.n302 VSUBS 0.007957f
C1201 B.n303 VSUBS 0.007957f
C1202 B.n304 VSUBS 0.005499f
C1203 B.n305 VSUBS 0.018435f
C1204 B.n306 VSUBS 0.006435f
C1205 B.n307 VSUBS 0.007957f
C1206 B.n308 VSUBS 0.007957f
C1207 B.n309 VSUBS 0.007957f
C1208 B.n310 VSUBS 0.007957f
C1209 B.n311 VSUBS 0.007957f
C1210 B.n312 VSUBS 0.007957f
C1211 B.n313 VSUBS 0.007957f
C1212 B.n314 VSUBS 0.007957f
C1213 B.n315 VSUBS 0.007957f
C1214 B.n316 VSUBS 0.007957f
C1215 B.n317 VSUBS 0.007957f
C1216 B.n318 VSUBS 0.006435f
C1217 B.n319 VSUBS 0.007957f
C1218 B.n320 VSUBS 0.007957f
C1219 B.n321 VSUBS 0.005499f
C1220 B.n322 VSUBS 0.007957f
C1221 B.n323 VSUBS 0.007957f
C1222 B.n324 VSUBS 0.007957f
C1223 B.n325 VSUBS 0.007957f
C1224 B.n326 VSUBS 0.007957f
C1225 B.n327 VSUBS 0.007957f
C1226 B.n328 VSUBS 0.007957f
C1227 B.n329 VSUBS 0.007957f
C1228 B.n330 VSUBS 0.007957f
C1229 B.n331 VSUBS 0.007957f
C1230 B.n332 VSUBS 0.007957f
C1231 B.n333 VSUBS 0.007957f
C1232 B.n334 VSUBS 0.007957f
C1233 B.n335 VSUBS 0.007957f
C1234 B.n336 VSUBS 0.007957f
C1235 B.n337 VSUBS 0.007957f
C1236 B.n338 VSUBS 0.007957f
C1237 B.n339 VSUBS 0.007957f
C1238 B.n340 VSUBS 0.007957f
C1239 B.n341 VSUBS 0.007957f
C1240 B.n342 VSUBS 0.007957f
C1241 B.n343 VSUBS 0.007957f
C1242 B.n344 VSUBS 0.007957f
C1243 B.n345 VSUBS 0.007957f
C1244 B.n346 VSUBS 0.007957f
C1245 B.n347 VSUBS 0.007957f
C1246 B.n348 VSUBS 0.007957f
C1247 B.n349 VSUBS 0.007957f
C1248 B.n350 VSUBS 0.007957f
C1249 B.n351 VSUBS 0.007957f
C1250 B.n352 VSUBS 0.007957f
C1251 B.n353 VSUBS 0.007957f
C1252 B.n354 VSUBS 0.007957f
C1253 B.n355 VSUBS 0.007957f
C1254 B.n356 VSUBS 0.007957f
C1255 B.n357 VSUBS 0.007957f
C1256 B.n358 VSUBS 0.007957f
C1257 B.n359 VSUBS 0.007957f
C1258 B.n360 VSUBS 0.007957f
C1259 B.n361 VSUBS 0.007957f
C1260 B.n362 VSUBS 0.007957f
C1261 B.n363 VSUBS 0.007957f
C1262 B.n364 VSUBS 0.007957f
C1263 B.n365 VSUBS 0.007957f
C1264 B.n366 VSUBS 0.007957f
C1265 B.n367 VSUBS 0.007957f
C1266 B.n368 VSUBS 0.007957f
C1267 B.n369 VSUBS 0.007957f
C1268 B.n370 VSUBS 0.007957f
C1269 B.n371 VSUBS 0.007957f
C1270 B.n372 VSUBS 0.007957f
C1271 B.n373 VSUBS 0.007957f
C1272 B.n374 VSUBS 0.007957f
C1273 B.n375 VSUBS 0.007957f
C1274 B.n376 VSUBS 0.007957f
C1275 B.n377 VSUBS 0.007957f
C1276 B.n378 VSUBS 0.007957f
C1277 B.n379 VSUBS 0.007957f
C1278 B.n380 VSUBS 0.007957f
C1279 B.n381 VSUBS 0.007957f
C1280 B.n382 VSUBS 0.007957f
C1281 B.n383 VSUBS 0.007957f
C1282 B.n384 VSUBS 0.007957f
C1283 B.n385 VSUBS 0.007957f
C1284 B.n386 VSUBS 0.007957f
C1285 B.n387 VSUBS 0.007957f
C1286 B.n388 VSUBS 0.007957f
C1287 B.n389 VSUBS 0.007957f
C1288 B.n390 VSUBS 0.007957f
C1289 B.n391 VSUBS 0.007957f
C1290 B.n392 VSUBS 0.007957f
C1291 B.n393 VSUBS 0.007957f
C1292 B.n394 VSUBS 0.007957f
C1293 B.n395 VSUBS 0.007957f
C1294 B.n396 VSUBS 0.007957f
C1295 B.n397 VSUBS 0.007957f
C1296 B.n398 VSUBS 0.007957f
C1297 B.n399 VSUBS 0.007957f
C1298 B.n400 VSUBS 0.007957f
C1299 B.n401 VSUBS 0.007957f
C1300 B.n402 VSUBS 0.007957f
C1301 B.n403 VSUBS 0.007957f
C1302 B.n404 VSUBS 0.007957f
C1303 B.n405 VSUBS 0.007957f
C1304 B.n406 VSUBS 0.007957f
C1305 B.n407 VSUBS 0.007957f
C1306 B.n408 VSUBS 0.007957f
C1307 B.n409 VSUBS 0.007957f
C1308 B.n410 VSUBS 0.007957f
C1309 B.n411 VSUBS 0.007957f
C1310 B.n412 VSUBS 0.007957f
C1311 B.n413 VSUBS 0.007957f
C1312 B.n414 VSUBS 0.007957f
C1313 B.n415 VSUBS 0.018754f
C1314 B.n416 VSUBS 0.018221f
C1315 B.n417 VSUBS 0.018221f
C1316 B.n418 VSUBS 0.007957f
C1317 B.n419 VSUBS 0.007957f
C1318 B.n420 VSUBS 0.007957f
C1319 B.n421 VSUBS 0.007957f
C1320 B.n422 VSUBS 0.007957f
C1321 B.n423 VSUBS 0.007957f
C1322 B.n424 VSUBS 0.007957f
C1323 B.n425 VSUBS 0.007957f
C1324 B.n426 VSUBS 0.007957f
C1325 B.n427 VSUBS 0.007957f
C1326 B.n428 VSUBS 0.007957f
C1327 B.n429 VSUBS 0.007957f
C1328 B.n430 VSUBS 0.007957f
C1329 B.n431 VSUBS 0.007957f
C1330 B.n432 VSUBS 0.007957f
C1331 B.n433 VSUBS 0.007957f
C1332 B.n434 VSUBS 0.007957f
C1333 B.n435 VSUBS 0.007957f
C1334 B.n436 VSUBS 0.007957f
C1335 B.n437 VSUBS 0.007957f
C1336 B.n438 VSUBS 0.007957f
C1337 B.n439 VSUBS 0.007957f
C1338 B.n440 VSUBS 0.007957f
C1339 B.n441 VSUBS 0.007957f
C1340 B.n442 VSUBS 0.007957f
C1341 B.n443 VSUBS 0.007957f
C1342 B.n444 VSUBS 0.007957f
C1343 B.n445 VSUBS 0.007957f
C1344 B.n446 VSUBS 0.007957f
C1345 B.n447 VSUBS 0.007957f
C1346 B.n448 VSUBS 0.007957f
C1347 B.n449 VSUBS 0.007957f
C1348 B.n450 VSUBS 0.007957f
C1349 B.n451 VSUBS 0.007957f
C1350 B.n452 VSUBS 0.007957f
C1351 B.n453 VSUBS 0.007957f
C1352 B.n454 VSUBS 0.007957f
C1353 B.n455 VSUBS 0.007957f
C1354 B.n456 VSUBS 0.007957f
C1355 B.n457 VSUBS 0.007957f
C1356 B.n458 VSUBS 0.007957f
C1357 B.n459 VSUBS 0.007957f
C1358 B.n460 VSUBS 0.007957f
C1359 B.n461 VSUBS 0.007957f
C1360 B.n462 VSUBS 0.007957f
C1361 B.n463 VSUBS 0.007957f
C1362 B.n464 VSUBS 0.007957f
C1363 B.n465 VSUBS 0.007957f
C1364 B.n466 VSUBS 0.007957f
C1365 B.n467 VSUBS 0.007957f
C1366 B.n468 VSUBS 0.007957f
C1367 B.n469 VSUBS 0.007957f
C1368 B.n470 VSUBS 0.018221f
C1369 B.n471 VSUBS 0.019171f
C1370 B.n472 VSUBS 0.017804f
C1371 B.n473 VSUBS 0.007957f
C1372 B.n474 VSUBS 0.007957f
C1373 B.n475 VSUBS 0.007957f
C1374 B.n476 VSUBS 0.007957f
C1375 B.n477 VSUBS 0.007957f
C1376 B.n478 VSUBS 0.007957f
C1377 B.n479 VSUBS 0.007957f
C1378 B.n480 VSUBS 0.007957f
C1379 B.n481 VSUBS 0.007957f
C1380 B.n482 VSUBS 0.007957f
C1381 B.n483 VSUBS 0.007957f
C1382 B.n484 VSUBS 0.007957f
C1383 B.n485 VSUBS 0.007957f
C1384 B.n486 VSUBS 0.007957f
C1385 B.n487 VSUBS 0.007957f
C1386 B.n488 VSUBS 0.007957f
C1387 B.n489 VSUBS 0.007957f
C1388 B.n490 VSUBS 0.007957f
C1389 B.n491 VSUBS 0.007957f
C1390 B.n492 VSUBS 0.007957f
C1391 B.n493 VSUBS 0.007957f
C1392 B.n494 VSUBS 0.007957f
C1393 B.n495 VSUBS 0.007957f
C1394 B.n496 VSUBS 0.007957f
C1395 B.n497 VSUBS 0.007957f
C1396 B.n498 VSUBS 0.007957f
C1397 B.n499 VSUBS 0.007957f
C1398 B.n500 VSUBS 0.007957f
C1399 B.n501 VSUBS 0.007957f
C1400 B.n502 VSUBS 0.007957f
C1401 B.n503 VSUBS 0.007957f
C1402 B.n504 VSUBS 0.007957f
C1403 B.n505 VSUBS 0.007957f
C1404 B.n506 VSUBS 0.007957f
C1405 B.n507 VSUBS 0.007957f
C1406 B.n508 VSUBS 0.007957f
C1407 B.n509 VSUBS 0.007957f
C1408 B.n510 VSUBS 0.007957f
C1409 B.n511 VSUBS 0.007957f
C1410 B.n512 VSUBS 0.007957f
C1411 B.n513 VSUBS 0.007957f
C1412 B.n514 VSUBS 0.007957f
C1413 B.n515 VSUBS 0.007957f
C1414 B.n516 VSUBS 0.007957f
C1415 B.n517 VSUBS 0.007957f
C1416 B.n518 VSUBS 0.007957f
C1417 B.n519 VSUBS 0.007957f
C1418 B.n520 VSUBS 0.007957f
C1419 B.n521 VSUBS 0.007957f
C1420 B.n522 VSUBS 0.007957f
C1421 B.n523 VSUBS 0.007957f
C1422 B.n524 VSUBS 0.007957f
C1423 B.n525 VSUBS 0.007957f
C1424 B.n526 VSUBS 0.007957f
C1425 B.n527 VSUBS 0.007957f
C1426 B.n528 VSUBS 0.007957f
C1427 B.n529 VSUBS 0.007957f
C1428 B.n530 VSUBS 0.007957f
C1429 B.n531 VSUBS 0.007957f
C1430 B.n532 VSUBS 0.007957f
C1431 B.n533 VSUBS 0.007957f
C1432 B.n534 VSUBS 0.007957f
C1433 B.n535 VSUBS 0.007957f
C1434 B.n536 VSUBS 0.007957f
C1435 B.n537 VSUBS 0.007957f
C1436 B.n538 VSUBS 0.007957f
C1437 B.n539 VSUBS 0.007957f
C1438 B.n540 VSUBS 0.007957f
C1439 B.n541 VSUBS 0.007957f
C1440 B.n542 VSUBS 0.007957f
C1441 B.n543 VSUBS 0.007957f
C1442 B.n544 VSUBS 0.007957f
C1443 B.n545 VSUBS 0.007957f
C1444 B.n546 VSUBS 0.007957f
C1445 B.n547 VSUBS 0.007957f
C1446 B.n548 VSUBS 0.007957f
C1447 B.n549 VSUBS 0.007957f
C1448 B.n550 VSUBS 0.007957f
C1449 B.n551 VSUBS 0.007957f
C1450 B.n552 VSUBS 0.007957f
C1451 B.n553 VSUBS 0.007957f
C1452 B.n554 VSUBS 0.007957f
C1453 B.n555 VSUBS 0.007957f
C1454 B.n556 VSUBS 0.007957f
C1455 B.n557 VSUBS 0.007957f
C1456 B.n558 VSUBS 0.007957f
C1457 B.n559 VSUBS 0.007957f
C1458 B.n560 VSUBS 0.007957f
C1459 B.n561 VSUBS 0.007957f
C1460 B.n562 VSUBS 0.007957f
C1461 B.n563 VSUBS 0.007957f
C1462 B.n564 VSUBS 0.007957f
C1463 B.n565 VSUBS 0.007957f
C1464 B.n566 VSUBS 0.007957f
C1465 B.n567 VSUBS 0.005499f
C1466 B.n568 VSUBS 0.018435f
C1467 B.n569 VSUBS 0.006435f
C1468 B.n570 VSUBS 0.007957f
C1469 B.n571 VSUBS 0.007957f
C1470 B.n572 VSUBS 0.007957f
C1471 B.n573 VSUBS 0.007957f
C1472 B.n574 VSUBS 0.007957f
C1473 B.n575 VSUBS 0.007957f
C1474 B.n576 VSUBS 0.007957f
C1475 B.n577 VSUBS 0.007957f
C1476 B.n578 VSUBS 0.007957f
C1477 B.n579 VSUBS 0.007957f
C1478 B.n580 VSUBS 0.007957f
C1479 B.n581 VSUBS 0.006435f
C1480 B.n582 VSUBS 0.018435f
C1481 B.n583 VSUBS 0.005499f
C1482 B.n584 VSUBS 0.007957f
C1483 B.n585 VSUBS 0.007957f
C1484 B.n586 VSUBS 0.007957f
C1485 B.n587 VSUBS 0.007957f
C1486 B.n588 VSUBS 0.007957f
C1487 B.n589 VSUBS 0.007957f
C1488 B.n590 VSUBS 0.007957f
C1489 B.n591 VSUBS 0.007957f
C1490 B.n592 VSUBS 0.007957f
C1491 B.n593 VSUBS 0.007957f
C1492 B.n594 VSUBS 0.007957f
C1493 B.n595 VSUBS 0.007957f
C1494 B.n596 VSUBS 0.007957f
C1495 B.n597 VSUBS 0.007957f
C1496 B.n598 VSUBS 0.007957f
C1497 B.n599 VSUBS 0.007957f
C1498 B.n600 VSUBS 0.007957f
C1499 B.n601 VSUBS 0.007957f
C1500 B.n602 VSUBS 0.007957f
C1501 B.n603 VSUBS 0.007957f
C1502 B.n604 VSUBS 0.007957f
C1503 B.n605 VSUBS 0.007957f
C1504 B.n606 VSUBS 0.007957f
C1505 B.n607 VSUBS 0.007957f
C1506 B.n608 VSUBS 0.007957f
C1507 B.n609 VSUBS 0.007957f
C1508 B.n610 VSUBS 0.007957f
C1509 B.n611 VSUBS 0.007957f
C1510 B.n612 VSUBS 0.007957f
C1511 B.n613 VSUBS 0.007957f
C1512 B.n614 VSUBS 0.007957f
C1513 B.n615 VSUBS 0.007957f
C1514 B.n616 VSUBS 0.007957f
C1515 B.n617 VSUBS 0.007957f
C1516 B.n618 VSUBS 0.007957f
C1517 B.n619 VSUBS 0.007957f
C1518 B.n620 VSUBS 0.007957f
C1519 B.n621 VSUBS 0.007957f
C1520 B.n622 VSUBS 0.007957f
C1521 B.n623 VSUBS 0.007957f
C1522 B.n624 VSUBS 0.007957f
C1523 B.n625 VSUBS 0.007957f
C1524 B.n626 VSUBS 0.007957f
C1525 B.n627 VSUBS 0.007957f
C1526 B.n628 VSUBS 0.007957f
C1527 B.n629 VSUBS 0.007957f
C1528 B.n630 VSUBS 0.007957f
C1529 B.n631 VSUBS 0.007957f
C1530 B.n632 VSUBS 0.007957f
C1531 B.n633 VSUBS 0.007957f
C1532 B.n634 VSUBS 0.007957f
C1533 B.n635 VSUBS 0.007957f
C1534 B.n636 VSUBS 0.007957f
C1535 B.n637 VSUBS 0.007957f
C1536 B.n638 VSUBS 0.007957f
C1537 B.n639 VSUBS 0.007957f
C1538 B.n640 VSUBS 0.007957f
C1539 B.n641 VSUBS 0.007957f
C1540 B.n642 VSUBS 0.007957f
C1541 B.n643 VSUBS 0.007957f
C1542 B.n644 VSUBS 0.007957f
C1543 B.n645 VSUBS 0.007957f
C1544 B.n646 VSUBS 0.007957f
C1545 B.n647 VSUBS 0.007957f
C1546 B.n648 VSUBS 0.007957f
C1547 B.n649 VSUBS 0.007957f
C1548 B.n650 VSUBS 0.007957f
C1549 B.n651 VSUBS 0.007957f
C1550 B.n652 VSUBS 0.007957f
C1551 B.n653 VSUBS 0.007957f
C1552 B.n654 VSUBS 0.007957f
C1553 B.n655 VSUBS 0.007957f
C1554 B.n656 VSUBS 0.007957f
C1555 B.n657 VSUBS 0.007957f
C1556 B.n658 VSUBS 0.007957f
C1557 B.n659 VSUBS 0.007957f
C1558 B.n660 VSUBS 0.007957f
C1559 B.n661 VSUBS 0.007957f
C1560 B.n662 VSUBS 0.007957f
C1561 B.n663 VSUBS 0.007957f
C1562 B.n664 VSUBS 0.007957f
C1563 B.n665 VSUBS 0.007957f
C1564 B.n666 VSUBS 0.007957f
C1565 B.n667 VSUBS 0.007957f
C1566 B.n668 VSUBS 0.007957f
C1567 B.n669 VSUBS 0.007957f
C1568 B.n670 VSUBS 0.007957f
C1569 B.n671 VSUBS 0.007957f
C1570 B.n672 VSUBS 0.007957f
C1571 B.n673 VSUBS 0.007957f
C1572 B.n674 VSUBS 0.007957f
C1573 B.n675 VSUBS 0.007957f
C1574 B.n676 VSUBS 0.007957f
C1575 B.n677 VSUBS 0.007957f
C1576 B.n678 VSUBS 0.018754f
C1577 B.n679 VSUBS 0.018221f
C1578 B.n680 VSUBS 0.018221f
C1579 B.n681 VSUBS 0.007957f
C1580 B.n682 VSUBS 0.007957f
C1581 B.n683 VSUBS 0.007957f
C1582 B.n684 VSUBS 0.007957f
C1583 B.n685 VSUBS 0.007957f
C1584 B.n686 VSUBS 0.007957f
C1585 B.n687 VSUBS 0.007957f
C1586 B.n688 VSUBS 0.007957f
C1587 B.n689 VSUBS 0.007957f
C1588 B.n690 VSUBS 0.007957f
C1589 B.n691 VSUBS 0.007957f
C1590 B.n692 VSUBS 0.007957f
C1591 B.n693 VSUBS 0.007957f
C1592 B.n694 VSUBS 0.007957f
C1593 B.n695 VSUBS 0.007957f
C1594 B.n696 VSUBS 0.007957f
C1595 B.n697 VSUBS 0.007957f
C1596 B.n698 VSUBS 0.007957f
C1597 B.n699 VSUBS 0.007957f
C1598 B.n700 VSUBS 0.007957f
C1599 B.n701 VSUBS 0.007957f
C1600 B.n702 VSUBS 0.007957f
C1601 B.n703 VSUBS 0.007957f
C1602 B.n704 VSUBS 0.007957f
C1603 B.n705 VSUBS 0.007957f
C1604 B.n706 VSUBS 0.007957f
C1605 B.n707 VSUBS 0.018017f
.ends

