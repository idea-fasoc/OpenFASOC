* NGSPICE file created from diff_pair_sample_1062.ext - technology: sky130A

.subckt diff_pair_sample_1062 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=5.9163 ps=31.12 w=15.17 l=0.79
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=0.79
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=0.79
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=5.9163 ps=31.12 w=15.17 l=0.79
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=0.79
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=5.9163 ps=31.12 w=15.17 l=0.79
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=5.9163 ps=31.12 w=15.17 l=0.79
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.9163 pd=31.12 as=0 ps=0 w=15.17 l=0.79
R0 VN VN.t0 716.765
R1 VN VN.t1 674.163
R2 VTAIL.n1 VTAIL.t2 48.8032
R3 VTAIL.n3 VTAIL.t3 48.803
R4 VTAIL.n0 VTAIL.t0 48.803
R5 VTAIL.n2 VTAIL.t1 48.803
R6 VTAIL.n1 VTAIL.n0 27.3927
R7 VTAIL.n3 VTAIL.n2 26.4272
R8 VTAIL.n2 VTAIL.n1 0.953086
R9 VTAIL VTAIL.n0 0.769897
R10 VTAIL VTAIL.n3 0.18369
R11 VDD2.n0 VDD2.t0 104.168
R12 VDD2.n0 VDD2.t1 65.4817
R13 VDD2 VDD2.n0 0.300069
R14 B.n58 B.t13 664.765
R15 B.n65 B.t6 664.765
R16 B.n151 B.t2 664.765
R17 B.n145 B.t10 664.765
R18 B.n466 B.n465 585
R19 B.n468 B.n91 585
R20 B.n471 B.n470 585
R21 B.n472 B.n90 585
R22 B.n474 B.n473 585
R23 B.n476 B.n89 585
R24 B.n479 B.n478 585
R25 B.n480 B.n88 585
R26 B.n482 B.n481 585
R27 B.n484 B.n87 585
R28 B.n487 B.n486 585
R29 B.n488 B.n86 585
R30 B.n490 B.n489 585
R31 B.n492 B.n85 585
R32 B.n495 B.n494 585
R33 B.n496 B.n84 585
R34 B.n498 B.n497 585
R35 B.n500 B.n83 585
R36 B.n503 B.n502 585
R37 B.n504 B.n82 585
R38 B.n506 B.n505 585
R39 B.n508 B.n81 585
R40 B.n511 B.n510 585
R41 B.n512 B.n80 585
R42 B.n514 B.n513 585
R43 B.n516 B.n79 585
R44 B.n519 B.n518 585
R45 B.n520 B.n78 585
R46 B.n522 B.n521 585
R47 B.n524 B.n77 585
R48 B.n527 B.n526 585
R49 B.n528 B.n76 585
R50 B.n530 B.n529 585
R51 B.n532 B.n75 585
R52 B.n535 B.n534 585
R53 B.n536 B.n74 585
R54 B.n538 B.n537 585
R55 B.n540 B.n73 585
R56 B.n543 B.n542 585
R57 B.n544 B.n72 585
R58 B.n546 B.n545 585
R59 B.n548 B.n71 585
R60 B.n551 B.n550 585
R61 B.n552 B.n70 585
R62 B.n554 B.n553 585
R63 B.n556 B.n69 585
R64 B.n559 B.n558 585
R65 B.n560 B.n68 585
R66 B.n562 B.n561 585
R67 B.n564 B.n67 585
R68 B.n567 B.n566 585
R69 B.n569 B.n64 585
R70 B.n571 B.n570 585
R71 B.n573 B.n63 585
R72 B.n576 B.n575 585
R73 B.n577 B.n62 585
R74 B.n579 B.n578 585
R75 B.n581 B.n61 585
R76 B.n584 B.n583 585
R77 B.n585 B.n57 585
R78 B.n587 B.n586 585
R79 B.n589 B.n56 585
R80 B.n592 B.n591 585
R81 B.n593 B.n55 585
R82 B.n595 B.n594 585
R83 B.n597 B.n54 585
R84 B.n600 B.n599 585
R85 B.n601 B.n53 585
R86 B.n603 B.n602 585
R87 B.n605 B.n52 585
R88 B.n608 B.n607 585
R89 B.n609 B.n51 585
R90 B.n611 B.n610 585
R91 B.n613 B.n50 585
R92 B.n616 B.n615 585
R93 B.n617 B.n49 585
R94 B.n619 B.n618 585
R95 B.n621 B.n48 585
R96 B.n624 B.n623 585
R97 B.n625 B.n47 585
R98 B.n627 B.n626 585
R99 B.n629 B.n46 585
R100 B.n632 B.n631 585
R101 B.n633 B.n45 585
R102 B.n635 B.n634 585
R103 B.n637 B.n44 585
R104 B.n640 B.n639 585
R105 B.n641 B.n43 585
R106 B.n643 B.n642 585
R107 B.n645 B.n42 585
R108 B.n648 B.n647 585
R109 B.n649 B.n41 585
R110 B.n651 B.n650 585
R111 B.n653 B.n40 585
R112 B.n656 B.n655 585
R113 B.n657 B.n39 585
R114 B.n659 B.n658 585
R115 B.n661 B.n38 585
R116 B.n664 B.n663 585
R117 B.n665 B.n37 585
R118 B.n667 B.n666 585
R119 B.n669 B.n36 585
R120 B.n672 B.n671 585
R121 B.n673 B.n35 585
R122 B.n675 B.n674 585
R123 B.n677 B.n34 585
R124 B.n680 B.n679 585
R125 B.n681 B.n33 585
R126 B.n683 B.n682 585
R127 B.n685 B.n32 585
R128 B.n688 B.n687 585
R129 B.n689 B.n31 585
R130 B.n464 B.n29 585
R131 B.n692 B.n29 585
R132 B.n463 B.n28 585
R133 B.n693 B.n28 585
R134 B.n462 B.n27 585
R135 B.n694 B.n27 585
R136 B.n461 B.n460 585
R137 B.n460 B.n23 585
R138 B.n459 B.n22 585
R139 B.n700 B.n22 585
R140 B.n458 B.n21 585
R141 B.n701 B.n21 585
R142 B.n457 B.n20 585
R143 B.n702 B.n20 585
R144 B.n456 B.n455 585
R145 B.n455 B.n16 585
R146 B.n454 B.n15 585
R147 B.n708 B.n15 585
R148 B.n453 B.n14 585
R149 B.n709 B.n14 585
R150 B.n452 B.n13 585
R151 B.n710 B.n13 585
R152 B.n451 B.n450 585
R153 B.n450 B.n12 585
R154 B.n449 B.n448 585
R155 B.n449 B.n8 585
R156 B.n447 B.n7 585
R157 B.n717 B.n7 585
R158 B.n446 B.n6 585
R159 B.n718 B.n6 585
R160 B.n445 B.n5 585
R161 B.n719 B.n5 585
R162 B.n444 B.n443 585
R163 B.n443 B.n4 585
R164 B.n442 B.n92 585
R165 B.n442 B.n441 585
R166 B.n431 B.n93 585
R167 B.n434 B.n93 585
R168 B.n433 B.n432 585
R169 B.n435 B.n433 585
R170 B.n430 B.n98 585
R171 B.n98 B.n97 585
R172 B.n429 B.n428 585
R173 B.n428 B.n427 585
R174 B.n100 B.n99 585
R175 B.n101 B.n100 585
R176 B.n420 B.n419 585
R177 B.n421 B.n420 585
R178 B.n418 B.n106 585
R179 B.n106 B.n105 585
R180 B.n417 B.n416 585
R181 B.n416 B.n415 585
R182 B.n108 B.n107 585
R183 B.n109 B.n108 585
R184 B.n408 B.n407 585
R185 B.n409 B.n408 585
R186 B.n406 B.n114 585
R187 B.n114 B.n113 585
R188 B.n405 B.n404 585
R189 B.n404 B.n403 585
R190 B.n400 B.n118 585
R191 B.n399 B.n398 585
R192 B.n396 B.n119 585
R193 B.n396 B.n117 585
R194 B.n395 B.n394 585
R195 B.n393 B.n392 585
R196 B.n391 B.n121 585
R197 B.n389 B.n388 585
R198 B.n387 B.n122 585
R199 B.n386 B.n385 585
R200 B.n383 B.n123 585
R201 B.n381 B.n380 585
R202 B.n379 B.n124 585
R203 B.n378 B.n377 585
R204 B.n375 B.n125 585
R205 B.n373 B.n372 585
R206 B.n371 B.n126 585
R207 B.n370 B.n369 585
R208 B.n367 B.n127 585
R209 B.n365 B.n364 585
R210 B.n363 B.n128 585
R211 B.n362 B.n361 585
R212 B.n359 B.n129 585
R213 B.n357 B.n356 585
R214 B.n355 B.n130 585
R215 B.n354 B.n353 585
R216 B.n351 B.n131 585
R217 B.n349 B.n348 585
R218 B.n347 B.n132 585
R219 B.n346 B.n345 585
R220 B.n343 B.n133 585
R221 B.n341 B.n340 585
R222 B.n339 B.n134 585
R223 B.n338 B.n337 585
R224 B.n335 B.n135 585
R225 B.n333 B.n332 585
R226 B.n331 B.n136 585
R227 B.n330 B.n329 585
R228 B.n327 B.n137 585
R229 B.n325 B.n324 585
R230 B.n323 B.n138 585
R231 B.n322 B.n321 585
R232 B.n319 B.n139 585
R233 B.n317 B.n316 585
R234 B.n315 B.n140 585
R235 B.n314 B.n313 585
R236 B.n311 B.n141 585
R237 B.n309 B.n308 585
R238 B.n307 B.n142 585
R239 B.n306 B.n305 585
R240 B.n303 B.n143 585
R241 B.n301 B.n300 585
R242 B.n298 B.n144 585
R243 B.n297 B.n296 585
R244 B.n294 B.n147 585
R245 B.n292 B.n291 585
R246 B.n290 B.n148 585
R247 B.n289 B.n288 585
R248 B.n286 B.n149 585
R249 B.n284 B.n283 585
R250 B.n282 B.n150 585
R251 B.n281 B.n280 585
R252 B.n278 B.n277 585
R253 B.n276 B.n275 585
R254 B.n274 B.n155 585
R255 B.n272 B.n271 585
R256 B.n270 B.n156 585
R257 B.n269 B.n268 585
R258 B.n266 B.n157 585
R259 B.n264 B.n263 585
R260 B.n262 B.n158 585
R261 B.n261 B.n260 585
R262 B.n258 B.n159 585
R263 B.n256 B.n255 585
R264 B.n254 B.n160 585
R265 B.n253 B.n252 585
R266 B.n250 B.n161 585
R267 B.n248 B.n247 585
R268 B.n246 B.n162 585
R269 B.n245 B.n244 585
R270 B.n242 B.n163 585
R271 B.n240 B.n239 585
R272 B.n238 B.n164 585
R273 B.n237 B.n236 585
R274 B.n234 B.n165 585
R275 B.n232 B.n231 585
R276 B.n230 B.n166 585
R277 B.n229 B.n228 585
R278 B.n226 B.n167 585
R279 B.n224 B.n223 585
R280 B.n222 B.n168 585
R281 B.n221 B.n220 585
R282 B.n218 B.n169 585
R283 B.n216 B.n215 585
R284 B.n214 B.n170 585
R285 B.n213 B.n212 585
R286 B.n210 B.n171 585
R287 B.n208 B.n207 585
R288 B.n206 B.n172 585
R289 B.n205 B.n204 585
R290 B.n202 B.n173 585
R291 B.n200 B.n199 585
R292 B.n198 B.n174 585
R293 B.n197 B.n196 585
R294 B.n194 B.n175 585
R295 B.n192 B.n191 585
R296 B.n190 B.n176 585
R297 B.n189 B.n188 585
R298 B.n186 B.n177 585
R299 B.n184 B.n183 585
R300 B.n182 B.n178 585
R301 B.n181 B.n180 585
R302 B.n116 B.n115 585
R303 B.n117 B.n116 585
R304 B.n402 B.n401 585
R305 B.n403 B.n402 585
R306 B.n112 B.n111 585
R307 B.n113 B.n112 585
R308 B.n411 B.n410 585
R309 B.n410 B.n409 585
R310 B.n412 B.n110 585
R311 B.n110 B.n109 585
R312 B.n414 B.n413 585
R313 B.n415 B.n414 585
R314 B.n104 B.n103 585
R315 B.n105 B.n104 585
R316 B.n423 B.n422 585
R317 B.n422 B.n421 585
R318 B.n424 B.n102 585
R319 B.n102 B.n101 585
R320 B.n426 B.n425 585
R321 B.n427 B.n426 585
R322 B.n96 B.n95 585
R323 B.n97 B.n96 585
R324 B.n437 B.n436 585
R325 B.n436 B.n435 585
R326 B.n438 B.n94 585
R327 B.n434 B.n94 585
R328 B.n440 B.n439 585
R329 B.n441 B.n440 585
R330 B.n3 B.n0 585
R331 B.n4 B.n3 585
R332 B.n716 B.n1 585
R333 B.n717 B.n716 585
R334 B.n715 B.n714 585
R335 B.n715 B.n8 585
R336 B.n713 B.n9 585
R337 B.n12 B.n9 585
R338 B.n712 B.n711 585
R339 B.n711 B.n710 585
R340 B.n11 B.n10 585
R341 B.n709 B.n11 585
R342 B.n707 B.n706 585
R343 B.n708 B.n707 585
R344 B.n705 B.n17 585
R345 B.n17 B.n16 585
R346 B.n704 B.n703 585
R347 B.n703 B.n702 585
R348 B.n19 B.n18 585
R349 B.n701 B.n19 585
R350 B.n699 B.n698 585
R351 B.n700 B.n699 585
R352 B.n697 B.n24 585
R353 B.n24 B.n23 585
R354 B.n696 B.n695 585
R355 B.n695 B.n694 585
R356 B.n26 B.n25 585
R357 B.n693 B.n26 585
R358 B.n691 B.n690 585
R359 B.n692 B.n691 585
R360 B.n720 B.n719 585
R361 B.n718 B.n2 585
R362 B.n691 B.n31 497.305
R363 B.n466 B.n29 497.305
R364 B.n404 B.n116 497.305
R365 B.n402 B.n118 497.305
R366 B.n467 B.n30 256.663
R367 B.n469 B.n30 256.663
R368 B.n475 B.n30 256.663
R369 B.n477 B.n30 256.663
R370 B.n483 B.n30 256.663
R371 B.n485 B.n30 256.663
R372 B.n491 B.n30 256.663
R373 B.n493 B.n30 256.663
R374 B.n499 B.n30 256.663
R375 B.n501 B.n30 256.663
R376 B.n507 B.n30 256.663
R377 B.n509 B.n30 256.663
R378 B.n515 B.n30 256.663
R379 B.n517 B.n30 256.663
R380 B.n523 B.n30 256.663
R381 B.n525 B.n30 256.663
R382 B.n531 B.n30 256.663
R383 B.n533 B.n30 256.663
R384 B.n539 B.n30 256.663
R385 B.n541 B.n30 256.663
R386 B.n547 B.n30 256.663
R387 B.n549 B.n30 256.663
R388 B.n555 B.n30 256.663
R389 B.n557 B.n30 256.663
R390 B.n563 B.n30 256.663
R391 B.n565 B.n30 256.663
R392 B.n572 B.n30 256.663
R393 B.n574 B.n30 256.663
R394 B.n580 B.n30 256.663
R395 B.n582 B.n30 256.663
R396 B.n588 B.n30 256.663
R397 B.n590 B.n30 256.663
R398 B.n596 B.n30 256.663
R399 B.n598 B.n30 256.663
R400 B.n604 B.n30 256.663
R401 B.n606 B.n30 256.663
R402 B.n612 B.n30 256.663
R403 B.n614 B.n30 256.663
R404 B.n620 B.n30 256.663
R405 B.n622 B.n30 256.663
R406 B.n628 B.n30 256.663
R407 B.n630 B.n30 256.663
R408 B.n636 B.n30 256.663
R409 B.n638 B.n30 256.663
R410 B.n644 B.n30 256.663
R411 B.n646 B.n30 256.663
R412 B.n652 B.n30 256.663
R413 B.n654 B.n30 256.663
R414 B.n660 B.n30 256.663
R415 B.n662 B.n30 256.663
R416 B.n668 B.n30 256.663
R417 B.n670 B.n30 256.663
R418 B.n676 B.n30 256.663
R419 B.n678 B.n30 256.663
R420 B.n684 B.n30 256.663
R421 B.n686 B.n30 256.663
R422 B.n397 B.n117 256.663
R423 B.n120 B.n117 256.663
R424 B.n390 B.n117 256.663
R425 B.n384 B.n117 256.663
R426 B.n382 B.n117 256.663
R427 B.n376 B.n117 256.663
R428 B.n374 B.n117 256.663
R429 B.n368 B.n117 256.663
R430 B.n366 B.n117 256.663
R431 B.n360 B.n117 256.663
R432 B.n358 B.n117 256.663
R433 B.n352 B.n117 256.663
R434 B.n350 B.n117 256.663
R435 B.n344 B.n117 256.663
R436 B.n342 B.n117 256.663
R437 B.n336 B.n117 256.663
R438 B.n334 B.n117 256.663
R439 B.n328 B.n117 256.663
R440 B.n326 B.n117 256.663
R441 B.n320 B.n117 256.663
R442 B.n318 B.n117 256.663
R443 B.n312 B.n117 256.663
R444 B.n310 B.n117 256.663
R445 B.n304 B.n117 256.663
R446 B.n302 B.n117 256.663
R447 B.n295 B.n117 256.663
R448 B.n293 B.n117 256.663
R449 B.n287 B.n117 256.663
R450 B.n285 B.n117 256.663
R451 B.n279 B.n117 256.663
R452 B.n154 B.n117 256.663
R453 B.n273 B.n117 256.663
R454 B.n267 B.n117 256.663
R455 B.n265 B.n117 256.663
R456 B.n259 B.n117 256.663
R457 B.n257 B.n117 256.663
R458 B.n251 B.n117 256.663
R459 B.n249 B.n117 256.663
R460 B.n243 B.n117 256.663
R461 B.n241 B.n117 256.663
R462 B.n235 B.n117 256.663
R463 B.n233 B.n117 256.663
R464 B.n227 B.n117 256.663
R465 B.n225 B.n117 256.663
R466 B.n219 B.n117 256.663
R467 B.n217 B.n117 256.663
R468 B.n211 B.n117 256.663
R469 B.n209 B.n117 256.663
R470 B.n203 B.n117 256.663
R471 B.n201 B.n117 256.663
R472 B.n195 B.n117 256.663
R473 B.n193 B.n117 256.663
R474 B.n187 B.n117 256.663
R475 B.n185 B.n117 256.663
R476 B.n179 B.n117 256.663
R477 B.n722 B.n721 256.663
R478 B.n687 B.n685 163.367
R479 B.n683 B.n33 163.367
R480 B.n679 B.n677 163.367
R481 B.n675 B.n35 163.367
R482 B.n671 B.n669 163.367
R483 B.n667 B.n37 163.367
R484 B.n663 B.n661 163.367
R485 B.n659 B.n39 163.367
R486 B.n655 B.n653 163.367
R487 B.n651 B.n41 163.367
R488 B.n647 B.n645 163.367
R489 B.n643 B.n43 163.367
R490 B.n639 B.n637 163.367
R491 B.n635 B.n45 163.367
R492 B.n631 B.n629 163.367
R493 B.n627 B.n47 163.367
R494 B.n623 B.n621 163.367
R495 B.n619 B.n49 163.367
R496 B.n615 B.n613 163.367
R497 B.n611 B.n51 163.367
R498 B.n607 B.n605 163.367
R499 B.n603 B.n53 163.367
R500 B.n599 B.n597 163.367
R501 B.n595 B.n55 163.367
R502 B.n591 B.n589 163.367
R503 B.n587 B.n57 163.367
R504 B.n583 B.n581 163.367
R505 B.n579 B.n62 163.367
R506 B.n575 B.n573 163.367
R507 B.n571 B.n64 163.367
R508 B.n566 B.n564 163.367
R509 B.n562 B.n68 163.367
R510 B.n558 B.n556 163.367
R511 B.n554 B.n70 163.367
R512 B.n550 B.n548 163.367
R513 B.n546 B.n72 163.367
R514 B.n542 B.n540 163.367
R515 B.n538 B.n74 163.367
R516 B.n534 B.n532 163.367
R517 B.n530 B.n76 163.367
R518 B.n526 B.n524 163.367
R519 B.n522 B.n78 163.367
R520 B.n518 B.n516 163.367
R521 B.n514 B.n80 163.367
R522 B.n510 B.n508 163.367
R523 B.n506 B.n82 163.367
R524 B.n502 B.n500 163.367
R525 B.n498 B.n84 163.367
R526 B.n494 B.n492 163.367
R527 B.n490 B.n86 163.367
R528 B.n486 B.n484 163.367
R529 B.n482 B.n88 163.367
R530 B.n478 B.n476 163.367
R531 B.n474 B.n90 163.367
R532 B.n470 B.n468 163.367
R533 B.n404 B.n114 163.367
R534 B.n408 B.n114 163.367
R535 B.n408 B.n108 163.367
R536 B.n416 B.n108 163.367
R537 B.n416 B.n106 163.367
R538 B.n420 B.n106 163.367
R539 B.n420 B.n100 163.367
R540 B.n428 B.n100 163.367
R541 B.n428 B.n98 163.367
R542 B.n433 B.n98 163.367
R543 B.n433 B.n93 163.367
R544 B.n442 B.n93 163.367
R545 B.n443 B.n442 163.367
R546 B.n443 B.n5 163.367
R547 B.n6 B.n5 163.367
R548 B.n7 B.n6 163.367
R549 B.n449 B.n7 163.367
R550 B.n450 B.n449 163.367
R551 B.n450 B.n13 163.367
R552 B.n14 B.n13 163.367
R553 B.n15 B.n14 163.367
R554 B.n455 B.n15 163.367
R555 B.n455 B.n20 163.367
R556 B.n21 B.n20 163.367
R557 B.n22 B.n21 163.367
R558 B.n460 B.n22 163.367
R559 B.n460 B.n27 163.367
R560 B.n28 B.n27 163.367
R561 B.n29 B.n28 163.367
R562 B.n398 B.n396 163.367
R563 B.n396 B.n395 163.367
R564 B.n392 B.n391 163.367
R565 B.n389 B.n122 163.367
R566 B.n385 B.n383 163.367
R567 B.n381 B.n124 163.367
R568 B.n377 B.n375 163.367
R569 B.n373 B.n126 163.367
R570 B.n369 B.n367 163.367
R571 B.n365 B.n128 163.367
R572 B.n361 B.n359 163.367
R573 B.n357 B.n130 163.367
R574 B.n353 B.n351 163.367
R575 B.n349 B.n132 163.367
R576 B.n345 B.n343 163.367
R577 B.n341 B.n134 163.367
R578 B.n337 B.n335 163.367
R579 B.n333 B.n136 163.367
R580 B.n329 B.n327 163.367
R581 B.n325 B.n138 163.367
R582 B.n321 B.n319 163.367
R583 B.n317 B.n140 163.367
R584 B.n313 B.n311 163.367
R585 B.n309 B.n142 163.367
R586 B.n305 B.n303 163.367
R587 B.n301 B.n144 163.367
R588 B.n296 B.n294 163.367
R589 B.n292 B.n148 163.367
R590 B.n288 B.n286 163.367
R591 B.n284 B.n150 163.367
R592 B.n280 B.n278 163.367
R593 B.n275 B.n274 163.367
R594 B.n272 B.n156 163.367
R595 B.n268 B.n266 163.367
R596 B.n264 B.n158 163.367
R597 B.n260 B.n258 163.367
R598 B.n256 B.n160 163.367
R599 B.n252 B.n250 163.367
R600 B.n248 B.n162 163.367
R601 B.n244 B.n242 163.367
R602 B.n240 B.n164 163.367
R603 B.n236 B.n234 163.367
R604 B.n232 B.n166 163.367
R605 B.n228 B.n226 163.367
R606 B.n224 B.n168 163.367
R607 B.n220 B.n218 163.367
R608 B.n216 B.n170 163.367
R609 B.n212 B.n210 163.367
R610 B.n208 B.n172 163.367
R611 B.n204 B.n202 163.367
R612 B.n200 B.n174 163.367
R613 B.n196 B.n194 163.367
R614 B.n192 B.n176 163.367
R615 B.n188 B.n186 163.367
R616 B.n184 B.n178 163.367
R617 B.n180 B.n116 163.367
R618 B.n402 B.n112 163.367
R619 B.n410 B.n112 163.367
R620 B.n410 B.n110 163.367
R621 B.n414 B.n110 163.367
R622 B.n414 B.n104 163.367
R623 B.n422 B.n104 163.367
R624 B.n422 B.n102 163.367
R625 B.n426 B.n102 163.367
R626 B.n426 B.n96 163.367
R627 B.n436 B.n96 163.367
R628 B.n436 B.n94 163.367
R629 B.n440 B.n94 163.367
R630 B.n440 B.n3 163.367
R631 B.n720 B.n3 163.367
R632 B.n716 B.n2 163.367
R633 B.n716 B.n715 163.367
R634 B.n715 B.n9 163.367
R635 B.n711 B.n9 163.367
R636 B.n711 B.n11 163.367
R637 B.n707 B.n11 163.367
R638 B.n707 B.n17 163.367
R639 B.n703 B.n17 163.367
R640 B.n703 B.n19 163.367
R641 B.n699 B.n19 163.367
R642 B.n699 B.n24 163.367
R643 B.n695 B.n24 163.367
R644 B.n695 B.n26 163.367
R645 B.n691 B.n26 163.367
R646 B.n65 B.t8 93.2435
R647 B.n151 B.t5 93.2435
R648 B.n58 B.t14 93.2238
R649 B.n145 B.t12 93.2238
R650 B.n403 B.n117 73.6384
R651 B.n692 B.n30 73.6384
R652 B.n686 B.n31 71.676
R653 B.n685 B.n684 71.676
R654 B.n678 B.n33 71.676
R655 B.n677 B.n676 71.676
R656 B.n670 B.n35 71.676
R657 B.n669 B.n668 71.676
R658 B.n662 B.n37 71.676
R659 B.n661 B.n660 71.676
R660 B.n654 B.n39 71.676
R661 B.n653 B.n652 71.676
R662 B.n646 B.n41 71.676
R663 B.n645 B.n644 71.676
R664 B.n638 B.n43 71.676
R665 B.n637 B.n636 71.676
R666 B.n630 B.n45 71.676
R667 B.n629 B.n628 71.676
R668 B.n622 B.n47 71.676
R669 B.n621 B.n620 71.676
R670 B.n614 B.n49 71.676
R671 B.n613 B.n612 71.676
R672 B.n606 B.n51 71.676
R673 B.n605 B.n604 71.676
R674 B.n598 B.n53 71.676
R675 B.n597 B.n596 71.676
R676 B.n590 B.n55 71.676
R677 B.n589 B.n588 71.676
R678 B.n582 B.n57 71.676
R679 B.n581 B.n580 71.676
R680 B.n574 B.n62 71.676
R681 B.n573 B.n572 71.676
R682 B.n565 B.n64 71.676
R683 B.n564 B.n563 71.676
R684 B.n557 B.n68 71.676
R685 B.n556 B.n555 71.676
R686 B.n549 B.n70 71.676
R687 B.n548 B.n547 71.676
R688 B.n541 B.n72 71.676
R689 B.n540 B.n539 71.676
R690 B.n533 B.n74 71.676
R691 B.n532 B.n531 71.676
R692 B.n525 B.n76 71.676
R693 B.n524 B.n523 71.676
R694 B.n517 B.n78 71.676
R695 B.n516 B.n515 71.676
R696 B.n509 B.n80 71.676
R697 B.n508 B.n507 71.676
R698 B.n501 B.n82 71.676
R699 B.n500 B.n499 71.676
R700 B.n493 B.n84 71.676
R701 B.n492 B.n491 71.676
R702 B.n485 B.n86 71.676
R703 B.n484 B.n483 71.676
R704 B.n477 B.n88 71.676
R705 B.n476 B.n475 71.676
R706 B.n469 B.n90 71.676
R707 B.n468 B.n467 71.676
R708 B.n467 B.n466 71.676
R709 B.n470 B.n469 71.676
R710 B.n475 B.n474 71.676
R711 B.n478 B.n477 71.676
R712 B.n483 B.n482 71.676
R713 B.n486 B.n485 71.676
R714 B.n491 B.n490 71.676
R715 B.n494 B.n493 71.676
R716 B.n499 B.n498 71.676
R717 B.n502 B.n501 71.676
R718 B.n507 B.n506 71.676
R719 B.n510 B.n509 71.676
R720 B.n515 B.n514 71.676
R721 B.n518 B.n517 71.676
R722 B.n523 B.n522 71.676
R723 B.n526 B.n525 71.676
R724 B.n531 B.n530 71.676
R725 B.n534 B.n533 71.676
R726 B.n539 B.n538 71.676
R727 B.n542 B.n541 71.676
R728 B.n547 B.n546 71.676
R729 B.n550 B.n549 71.676
R730 B.n555 B.n554 71.676
R731 B.n558 B.n557 71.676
R732 B.n563 B.n562 71.676
R733 B.n566 B.n565 71.676
R734 B.n572 B.n571 71.676
R735 B.n575 B.n574 71.676
R736 B.n580 B.n579 71.676
R737 B.n583 B.n582 71.676
R738 B.n588 B.n587 71.676
R739 B.n591 B.n590 71.676
R740 B.n596 B.n595 71.676
R741 B.n599 B.n598 71.676
R742 B.n604 B.n603 71.676
R743 B.n607 B.n606 71.676
R744 B.n612 B.n611 71.676
R745 B.n615 B.n614 71.676
R746 B.n620 B.n619 71.676
R747 B.n623 B.n622 71.676
R748 B.n628 B.n627 71.676
R749 B.n631 B.n630 71.676
R750 B.n636 B.n635 71.676
R751 B.n639 B.n638 71.676
R752 B.n644 B.n643 71.676
R753 B.n647 B.n646 71.676
R754 B.n652 B.n651 71.676
R755 B.n655 B.n654 71.676
R756 B.n660 B.n659 71.676
R757 B.n663 B.n662 71.676
R758 B.n668 B.n667 71.676
R759 B.n671 B.n670 71.676
R760 B.n676 B.n675 71.676
R761 B.n679 B.n678 71.676
R762 B.n684 B.n683 71.676
R763 B.n687 B.n686 71.676
R764 B.n397 B.n118 71.676
R765 B.n395 B.n120 71.676
R766 B.n391 B.n390 71.676
R767 B.n384 B.n122 71.676
R768 B.n383 B.n382 71.676
R769 B.n376 B.n124 71.676
R770 B.n375 B.n374 71.676
R771 B.n368 B.n126 71.676
R772 B.n367 B.n366 71.676
R773 B.n360 B.n128 71.676
R774 B.n359 B.n358 71.676
R775 B.n352 B.n130 71.676
R776 B.n351 B.n350 71.676
R777 B.n344 B.n132 71.676
R778 B.n343 B.n342 71.676
R779 B.n336 B.n134 71.676
R780 B.n335 B.n334 71.676
R781 B.n328 B.n136 71.676
R782 B.n327 B.n326 71.676
R783 B.n320 B.n138 71.676
R784 B.n319 B.n318 71.676
R785 B.n312 B.n140 71.676
R786 B.n311 B.n310 71.676
R787 B.n304 B.n142 71.676
R788 B.n303 B.n302 71.676
R789 B.n295 B.n144 71.676
R790 B.n294 B.n293 71.676
R791 B.n287 B.n148 71.676
R792 B.n286 B.n285 71.676
R793 B.n279 B.n150 71.676
R794 B.n278 B.n154 71.676
R795 B.n274 B.n273 71.676
R796 B.n267 B.n156 71.676
R797 B.n266 B.n265 71.676
R798 B.n259 B.n158 71.676
R799 B.n258 B.n257 71.676
R800 B.n251 B.n160 71.676
R801 B.n250 B.n249 71.676
R802 B.n243 B.n162 71.676
R803 B.n242 B.n241 71.676
R804 B.n235 B.n164 71.676
R805 B.n234 B.n233 71.676
R806 B.n227 B.n166 71.676
R807 B.n226 B.n225 71.676
R808 B.n219 B.n168 71.676
R809 B.n218 B.n217 71.676
R810 B.n211 B.n170 71.676
R811 B.n210 B.n209 71.676
R812 B.n203 B.n172 71.676
R813 B.n202 B.n201 71.676
R814 B.n195 B.n174 71.676
R815 B.n194 B.n193 71.676
R816 B.n187 B.n176 71.676
R817 B.n186 B.n185 71.676
R818 B.n179 B.n178 71.676
R819 B.n398 B.n397 71.676
R820 B.n392 B.n120 71.676
R821 B.n390 B.n389 71.676
R822 B.n385 B.n384 71.676
R823 B.n382 B.n381 71.676
R824 B.n377 B.n376 71.676
R825 B.n374 B.n373 71.676
R826 B.n369 B.n368 71.676
R827 B.n366 B.n365 71.676
R828 B.n361 B.n360 71.676
R829 B.n358 B.n357 71.676
R830 B.n353 B.n352 71.676
R831 B.n350 B.n349 71.676
R832 B.n345 B.n344 71.676
R833 B.n342 B.n341 71.676
R834 B.n337 B.n336 71.676
R835 B.n334 B.n333 71.676
R836 B.n329 B.n328 71.676
R837 B.n326 B.n325 71.676
R838 B.n321 B.n320 71.676
R839 B.n318 B.n317 71.676
R840 B.n313 B.n312 71.676
R841 B.n310 B.n309 71.676
R842 B.n305 B.n304 71.676
R843 B.n302 B.n301 71.676
R844 B.n296 B.n295 71.676
R845 B.n293 B.n292 71.676
R846 B.n288 B.n287 71.676
R847 B.n285 B.n284 71.676
R848 B.n280 B.n279 71.676
R849 B.n275 B.n154 71.676
R850 B.n273 B.n272 71.676
R851 B.n268 B.n267 71.676
R852 B.n265 B.n264 71.676
R853 B.n260 B.n259 71.676
R854 B.n257 B.n256 71.676
R855 B.n252 B.n251 71.676
R856 B.n249 B.n248 71.676
R857 B.n244 B.n243 71.676
R858 B.n241 B.n240 71.676
R859 B.n236 B.n235 71.676
R860 B.n233 B.n232 71.676
R861 B.n228 B.n227 71.676
R862 B.n225 B.n224 71.676
R863 B.n220 B.n219 71.676
R864 B.n217 B.n216 71.676
R865 B.n212 B.n211 71.676
R866 B.n209 B.n208 71.676
R867 B.n204 B.n203 71.676
R868 B.n201 B.n200 71.676
R869 B.n196 B.n195 71.676
R870 B.n193 B.n192 71.676
R871 B.n188 B.n187 71.676
R872 B.n185 B.n184 71.676
R873 B.n180 B.n179 71.676
R874 B.n721 B.n720 71.676
R875 B.n721 B.n2 71.676
R876 B.n66 B.t9 71.5223
R877 B.n152 B.t4 71.5223
R878 B.n59 B.t15 71.5026
R879 B.n146 B.t11 71.5026
R880 B.n60 B.n59 59.5399
R881 B.n568 B.n66 59.5399
R882 B.n153 B.n152 59.5399
R883 B.n299 B.n146 59.5399
R884 B.n403 B.n113 36.5507
R885 B.n409 B.n113 36.5507
R886 B.n409 B.n109 36.5507
R887 B.n415 B.n109 36.5507
R888 B.n421 B.n105 36.5507
R889 B.n421 B.n101 36.5507
R890 B.n427 B.n101 36.5507
R891 B.n427 B.n97 36.5507
R892 B.n435 B.n97 36.5507
R893 B.n435 B.n434 36.5507
R894 B.n441 B.n4 36.5507
R895 B.n719 B.n4 36.5507
R896 B.n719 B.n718 36.5507
R897 B.n718 B.n717 36.5507
R898 B.n717 B.n8 36.5507
R899 B.n710 B.n12 36.5507
R900 B.n710 B.n709 36.5507
R901 B.n709 B.n708 36.5507
R902 B.n708 B.n16 36.5507
R903 B.n702 B.n16 36.5507
R904 B.n702 B.n701 36.5507
R905 B.n700 B.n23 36.5507
R906 B.n694 B.n23 36.5507
R907 B.n694 B.n693 36.5507
R908 B.n693 B.n692 36.5507
R909 B.n401 B.n400 32.3127
R910 B.n405 B.n115 32.3127
R911 B.n465 B.n464 32.3127
R912 B.n690 B.n689 32.3127
R913 B.n415 B.t3 27.4132
R914 B.n441 B.t0 27.4132
R915 B.t1 B.n8 27.4132
R916 B.t7 B.n700 27.4132
R917 B.n59 B.n58 21.7217
R918 B.n66 B.n65 21.7217
R919 B.n152 B.n151 21.7217
R920 B.n146 B.n145 21.7217
R921 B B.n722 18.0485
R922 B.n401 B.n111 10.6151
R923 B.n411 B.n111 10.6151
R924 B.n412 B.n411 10.6151
R925 B.n413 B.n412 10.6151
R926 B.n413 B.n103 10.6151
R927 B.n423 B.n103 10.6151
R928 B.n424 B.n423 10.6151
R929 B.n425 B.n424 10.6151
R930 B.n425 B.n95 10.6151
R931 B.n437 B.n95 10.6151
R932 B.n438 B.n437 10.6151
R933 B.n439 B.n438 10.6151
R934 B.n439 B.n0 10.6151
R935 B.n400 B.n399 10.6151
R936 B.n399 B.n119 10.6151
R937 B.n394 B.n119 10.6151
R938 B.n394 B.n393 10.6151
R939 B.n393 B.n121 10.6151
R940 B.n388 B.n121 10.6151
R941 B.n388 B.n387 10.6151
R942 B.n387 B.n386 10.6151
R943 B.n386 B.n123 10.6151
R944 B.n380 B.n123 10.6151
R945 B.n380 B.n379 10.6151
R946 B.n379 B.n378 10.6151
R947 B.n378 B.n125 10.6151
R948 B.n372 B.n125 10.6151
R949 B.n372 B.n371 10.6151
R950 B.n371 B.n370 10.6151
R951 B.n370 B.n127 10.6151
R952 B.n364 B.n127 10.6151
R953 B.n364 B.n363 10.6151
R954 B.n363 B.n362 10.6151
R955 B.n362 B.n129 10.6151
R956 B.n356 B.n129 10.6151
R957 B.n356 B.n355 10.6151
R958 B.n355 B.n354 10.6151
R959 B.n354 B.n131 10.6151
R960 B.n348 B.n131 10.6151
R961 B.n348 B.n347 10.6151
R962 B.n347 B.n346 10.6151
R963 B.n346 B.n133 10.6151
R964 B.n340 B.n133 10.6151
R965 B.n340 B.n339 10.6151
R966 B.n339 B.n338 10.6151
R967 B.n338 B.n135 10.6151
R968 B.n332 B.n135 10.6151
R969 B.n332 B.n331 10.6151
R970 B.n331 B.n330 10.6151
R971 B.n330 B.n137 10.6151
R972 B.n324 B.n137 10.6151
R973 B.n324 B.n323 10.6151
R974 B.n323 B.n322 10.6151
R975 B.n322 B.n139 10.6151
R976 B.n316 B.n139 10.6151
R977 B.n316 B.n315 10.6151
R978 B.n315 B.n314 10.6151
R979 B.n314 B.n141 10.6151
R980 B.n308 B.n141 10.6151
R981 B.n308 B.n307 10.6151
R982 B.n307 B.n306 10.6151
R983 B.n306 B.n143 10.6151
R984 B.n300 B.n143 10.6151
R985 B.n298 B.n297 10.6151
R986 B.n297 B.n147 10.6151
R987 B.n291 B.n147 10.6151
R988 B.n291 B.n290 10.6151
R989 B.n290 B.n289 10.6151
R990 B.n289 B.n149 10.6151
R991 B.n283 B.n149 10.6151
R992 B.n283 B.n282 10.6151
R993 B.n282 B.n281 10.6151
R994 B.n277 B.n276 10.6151
R995 B.n276 B.n155 10.6151
R996 B.n271 B.n155 10.6151
R997 B.n271 B.n270 10.6151
R998 B.n270 B.n269 10.6151
R999 B.n269 B.n157 10.6151
R1000 B.n263 B.n157 10.6151
R1001 B.n263 B.n262 10.6151
R1002 B.n262 B.n261 10.6151
R1003 B.n261 B.n159 10.6151
R1004 B.n255 B.n159 10.6151
R1005 B.n255 B.n254 10.6151
R1006 B.n254 B.n253 10.6151
R1007 B.n253 B.n161 10.6151
R1008 B.n247 B.n161 10.6151
R1009 B.n247 B.n246 10.6151
R1010 B.n246 B.n245 10.6151
R1011 B.n245 B.n163 10.6151
R1012 B.n239 B.n163 10.6151
R1013 B.n239 B.n238 10.6151
R1014 B.n238 B.n237 10.6151
R1015 B.n237 B.n165 10.6151
R1016 B.n231 B.n165 10.6151
R1017 B.n231 B.n230 10.6151
R1018 B.n230 B.n229 10.6151
R1019 B.n229 B.n167 10.6151
R1020 B.n223 B.n167 10.6151
R1021 B.n223 B.n222 10.6151
R1022 B.n222 B.n221 10.6151
R1023 B.n221 B.n169 10.6151
R1024 B.n215 B.n169 10.6151
R1025 B.n215 B.n214 10.6151
R1026 B.n214 B.n213 10.6151
R1027 B.n213 B.n171 10.6151
R1028 B.n207 B.n171 10.6151
R1029 B.n207 B.n206 10.6151
R1030 B.n206 B.n205 10.6151
R1031 B.n205 B.n173 10.6151
R1032 B.n199 B.n173 10.6151
R1033 B.n199 B.n198 10.6151
R1034 B.n198 B.n197 10.6151
R1035 B.n197 B.n175 10.6151
R1036 B.n191 B.n175 10.6151
R1037 B.n191 B.n190 10.6151
R1038 B.n190 B.n189 10.6151
R1039 B.n189 B.n177 10.6151
R1040 B.n183 B.n177 10.6151
R1041 B.n183 B.n182 10.6151
R1042 B.n182 B.n181 10.6151
R1043 B.n181 B.n115 10.6151
R1044 B.n406 B.n405 10.6151
R1045 B.n407 B.n406 10.6151
R1046 B.n407 B.n107 10.6151
R1047 B.n417 B.n107 10.6151
R1048 B.n418 B.n417 10.6151
R1049 B.n419 B.n418 10.6151
R1050 B.n419 B.n99 10.6151
R1051 B.n429 B.n99 10.6151
R1052 B.n430 B.n429 10.6151
R1053 B.n432 B.n430 10.6151
R1054 B.n432 B.n431 10.6151
R1055 B.n431 B.n92 10.6151
R1056 B.n444 B.n92 10.6151
R1057 B.n445 B.n444 10.6151
R1058 B.n446 B.n445 10.6151
R1059 B.n447 B.n446 10.6151
R1060 B.n448 B.n447 10.6151
R1061 B.n451 B.n448 10.6151
R1062 B.n452 B.n451 10.6151
R1063 B.n453 B.n452 10.6151
R1064 B.n454 B.n453 10.6151
R1065 B.n456 B.n454 10.6151
R1066 B.n457 B.n456 10.6151
R1067 B.n458 B.n457 10.6151
R1068 B.n459 B.n458 10.6151
R1069 B.n461 B.n459 10.6151
R1070 B.n462 B.n461 10.6151
R1071 B.n463 B.n462 10.6151
R1072 B.n464 B.n463 10.6151
R1073 B.n714 B.n1 10.6151
R1074 B.n714 B.n713 10.6151
R1075 B.n713 B.n712 10.6151
R1076 B.n712 B.n10 10.6151
R1077 B.n706 B.n10 10.6151
R1078 B.n706 B.n705 10.6151
R1079 B.n705 B.n704 10.6151
R1080 B.n704 B.n18 10.6151
R1081 B.n698 B.n18 10.6151
R1082 B.n698 B.n697 10.6151
R1083 B.n697 B.n696 10.6151
R1084 B.n696 B.n25 10.6151
R1085 B.n690 B.n25 10.6151
R1086 B.n689 B.n688 10.6151
R1087 B.n688 B.n32 10.6151
R1088 B.n682 B.n32 10.6151
R1089 B.n682 B.n681 10.6151
R1090 B.n681 B.n680 10.6151
R1091 B.n680 B.n34 10.6151
R1092 B.n674 B.n34 10.6151
R1093 B.n674 B.n673 10.6151
R1094 B.n673 B.n672 10.6151
R1095 B.n672 B.n36 10.6151
R1096 B.n666 B.n36 10.6151
R1097 B.n666 B.n665 10.6151
R1098 B.n665 B.n664 10.6151
R1099 B.n664 B.n38 10.6151
R1100 B.n658 B.n38 10.6151
R1101 B.n658 B.n657 10.6151
R1102 B.n657 B.n656 10.6151
R1103 B.n656 B.n40 10.6151
R1104 B.n650 B.n40 10.6151
R1105 B.n650 B.n649 10.6151
R1106 B.n649 B.n648 10.6151
R1107 B.n648 B.n42 10.6151
R1108 B.n642 B.n42 10.6151
R1109 B.n642 B.n641 10.6151
R1110 B.n641 B.n640 10.6151
R1111 B.n640 B.n44 10.6151
R1112 B.n634 B.n44 10.6151
R1113 B.n634 B.n633 10.6151
R1114 B.n633 B.n632 10.6151
R1115 B.n632 B.n46 10.6151
R1116 B.n626 B.n46 10.6151
R1117 B.n626 B.n625 10.6151
R1118 B.n625 B.n624 10.6151
R1119 B.n624 B.n48 10.6151
R1120 B.n618 B.n48 10.6151
R1121 B.n618 B.n617 10.6151
R1122 B.n617 B.n616 10.6151
R1123 B.n616 B.n50 10.6151
R1124 B.n610 B.n50 10.6151
R1125 B.n610 B.n609 10.6151
R1126 B.n609 B.n608 10.6151
R1127 B.n608 B.n52 10.6151
R1128 B.n602 B.n52 10.6151
R1129 B.n602 B.n601 10.6151
R1130 B.n601 B.n600 10.6151
R1131 B.n600 B.n54 10.6151
R1132 B.n594 B.n54 10.6151
R1133 B.n594 B.n593 10.6151
R1134 B.n593 B.n592 10.6151
R1135 B.n592 B.n56 10.6151
R1136 B.n586 B.n585 10.6151
R1137 B.n585 B.n584 10.6151
R1138 B.n584 B.n61 10.6151
R1139 B.n578 B.n61 10.6151
R1140 B.n578 B.n577 10.6151
R1141 B.n577 B.n576 10.6151
R1142 B.n576 B.n63 10.6151
R1143 B.n570 B.n63 10.6151
R1144 B.n570 B.n569 10.6151
R1145 B.n567 B.n67 10.6151
R1146 B.n561 B.n67 10.6151
R1147 B.n561 B.n560 10.6151
R1148 B.n560 B.n559 10.6151
R1149 B.n559 B.n69 10.6151
R1150 B.n553 B.n69 10.6151
R1151 B.n553 B.n552 10.6151
R1152 B.n552 B.n551 10.6151
R1153 B.n551 B.n71 10.6151
R1154 B.n545 B.n71 10.6151
R1155 B.n545 B.n544 10.6151
R1156 B.n544 B.n543 10.6151
R1157 B.n543 B.n73 10.6151
R1158 B.n537 B.n73 10.6151
R1159 B.n537 B.n536 10.6151
R1160 B.n536 B.n535 10.6151
R1161 B.n535 B.n75 10.6151
R1162 B.n529 B.n75 10.6151
R1163 B.n529 B.n528 10.6151
R1164 B.n528 B.n527 10.6151
R1165 B.n527 B.n77 10.6151
R1166 B.n521 B.n77 10.6151
R1167 B.n521 B.n520 10.6151
R1168 B.n520 B.n519 10.6151
R1169 B.n519 B.n79 10.6151
R1170 B.n513 B.n79 10.6151
R1171 B.n513 B.n512 10.6151
R1172 B.n512 B.n511 10.6151
R1173 B.n511 B.n81 10.6151
R1174 B.n505 B.n81 10.6151
R1175 B.n505 B.n504 10.6151
R1176 B.n504 B.n503 10.6151
R1177 B.n503 B.n83 10.6151
R1178 B.n497 B.n83 10.6151
R1179 B.n497 B.n496 10.6151
R1180 B.n496 B.n495 10.6151
R1181 B.n495 B.n85 10.6151
R1182 B.n489 B.n85 10.6151
R1183 B.n489 B.n488 10.6151
R1184 B.n488 B.n487 10.6151
R1185 B.n487 B.n87 10.6151
R1186 B.n481 B.n87 10.6151
R1187 B.n481 B.n480 10.6151
R1188 B.n480 B.n479 10.6151
R1189 B.n479 B.n89 10.6151
R1190 B.n473 B.n89 10.6151
R1191 B.n473 B.n472 10.6151
R1192 B.n472 B.n471 10.6151
R1193 B.n471 B.n91 10.6151
R1194 B.n465 B.n91 10.6151
R1195 B.t3 B.n105 9.13805
R1196 B.n434 B.t0 9.13805
R1197 B.n12 B.t1 9.13805
R1198 B.n701 B.t7 9.13805
R1199 B.n300 B.n299 8.74196
R1200 B.n277 B.n153 8.74196
R1201 B.n60 B.n56 8.74196
R1202 B.n568 B.n567 8.74196
R1203 B.n722 B.n0 8.11757
R1204 B.n722 B.n1 8.11757
R1205 B.n299 B.n298 1.87367
R1206 B.n281 B.n153 1.87367
R1207 B.n586 B.n60 1.87367
R1208 B.n569 B.n568 1.87367
R1209 VP.n0 VP.t0 716.385
R1210 VP.n0 VP.t1 674.111
R1211 VP VP.n0 0.0516364
R1212 VDD1 VDD1.t0 104.933
R1213 VDD1 VDD1.t1 65.7813
C0 VP VDD2 0.259202f
C1 VP VTAIL 1.93853f
C2 VN VP 5.18947f
C3 VDD1 VP 2.66168f
C4 VDD2 VTAIL 6.67891f
C5 VN VDD2 2.55636f
C6 VN VTAIL 1.92383f
C7 VDD1 VDD2 0.471712f
C8 VDD1 VTAIL 6.6458f
C9 VDD1 VN 0.14863f
C10 VDD2 B 4.360122f
C11 VDD1 B 7.44312f
C12 VTAIL B 7.638114f
C13 VN B 8.87859f
C14 VP B 4.352852f
C15 VDD1.t1 B 2.86727f
C16 VDD1.t0 B 3.43075f
C17 VP.t0 B 1.77814f
C18 VP.t1 B 1.64314f
C19 VP.n0 B 4.46085f
C20 VDD2.t0 B 3.43249f
C21 VDD2.t1 B 2.88986f
C22 VDD2.n0 B 2.92454f
C23 VTAIL.t0 B 2.12436f
C24 VTAIL.n0 B 1.21581f
C25 VTAIL.t2 B 2.12437f
C26 VTAIL.n1 B 1.22509f
C27 VTAIL.t1 B 2.12436f
C28 VTAIL.n2 B 1.17618f
C29 VTAIL.t3 B 2.12436f
C30 VTAIL.n3 B 1.13719f
C31 VN.t1 B 1.60971f
C32 VN.t0 B 1.74474f
.ends

