* NGSPICE file created from diff_pair_sample_1621.ext - technology: sky130A

.subckt diff_pair_sample_1621 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=0 ps=0 w=6.5 l=3.58
X1 VDD1.t3 VP.t0 VTAIL.t4 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=1.0725 pd=6.83 as=2.535 ps=13.78 w=6.5 l=3.58
X2 VTAIL.t5 VP.t1 VDD1.t2 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=1.0725 ps=6.83 w=6.5 l=3.58
X3 B.t8 B.t6 B.t7 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=0 ps=0 w=6.5 l=3.58
X4 VTAIL.t6 VP.t2 VDD1.t1 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=1.0725 ps=6.83 w=6.5 l=3.58
X5 B.t5 B.t3 B.t4 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=0 ps=0 w=6.5 l=3.58
X6 VDD2.t3 VN.t0 VTAIL.t1 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=1.0725 pd=6.83 as=2.535 ps=13.78 w=6.5 l=3.58
X7 VDD1.t0 VP.t3 VTAIL.t7 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=1.0725 pd=6.83 as=2.535 ps=13.78 w=6.5 l=3.58
X8 VTAIL.t2 VN.t1 VDD2.t2 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=1.0725 ps=6.83 w=6.5 l=3.58
X9 B.t2 B.t0 B.t1 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=0 ps=0 w=6.5 l=3.58
X10 VDD2.t1 VN.t2 VTAIL.t3 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=1.0725 pd=6.83 as=2.535 ps=13.78 w=6.5 l=3.58
X11 VTAIL.t0 VN.t3 VDD2.t0 w_n3316_n2268# sky130_fd_pr__pfet_01v8 ad=2.535 pd=13.78 as=1.0725 ps=6.83 w=6.5 l=3.58
R0 B.n308 B.n101 585
R1 B.n307 B.n306 585
R2 B.n305 B.n102 585
R3 B.n304 B.n303 585
R4 B.n302 B.n103 585
R5 B.n301 B.n300 585
R6 B.n299 B.n104 585
R7 B.n298 B.n297 585
R8 B.n296 B.n105 585
R9 B.n295 B.n294 585
R10 B.n293 B.n106 585
R11 B.n292 B.n291 585
R12 B.n290 B.n107 585
R13 B.n289 B.n288 585
R14 B.n287 B.n108 585
R15 B.n286 B.n285 585
R16 B.n284 B.n109 585
R17 B.n283 B.n282 585
R18 B.n281 B.n110 585
R19 B.n280 B.n279 585
R20 B.n278 B.n111 585
R21 B.n277 B.n276 585
R22 B.n275 B.n112 585
R23 B.n274 B.n273 585
R24 B.n272 B.n113 585
R25 B.n271 B.n270 585
R26 B.n266 B.n114 585
R27 B.n265 B.n264 585
R28 B.n263 B.n115 585
R29 B.n262 B.n261 585
R30 B.n260 B.n116 585
R31 B.n259 B.n258 585
R32 B.n257 B.n117 585
R33 B.n256 B.n255 585
R34 B.n254 B.n118 585
R35 B.n252 B.n251 585
R36 B.n250 B.n121 585
R37 B.n249 B.n248 585
R38 B.n247 B.n122 585
R39 B.n246 B.n245 585
R40 B.n244 B.n123 585
R41 B.n243 B.n242 585
R42 B.n241 B.n124 585
R43 B.n240 B.n239 585
R44 B.n238 B.n125 585
R45 B.n237 B.n236 585
R46 B.n235 B.n126 585
R47 B.n234 B.n233 585
R48 B.n232 B.n127 585
R49 B.n231 B.n230 585
R50 B.n229 B.n128 585
R51 B.n228 B.n227 585
R52 B.n226 B.n129 585
R53 B.n225 B.n224 585
R54 B.n223 B.n130 585
R55 B.n222 B.n221 585
R56 B.n220 B.n131 585
R57 B.n219 B.n218 585
R58 B.n217 B.n132 585
R59 B.n216 B.n215 585
R60 B.n310 B.n309 585
R61 B.n311 B.n100 585
R62 B.n313 B.n312 585
R63 B.n314 B.n99 585
R64 B.n316 B.n315 585
R65 B.n317 B.n98 585
R66 B.n319 B.n318 585
R67 B.n320 B.n97 585
R68 B.n322 B.n321 585
R69 B.n323 B.n96 585
R70 B.n325 B.n324 585
R71 B.n326 B.n95 585
R72 B.n328 B.n327 585
R73 B.n329 B.n94 585
R74 B.n331 B.n330 585
R75 B.n332 B.n93 585
R76 B.n334 B.n333 585
R77 B.n335 B.n92 585
R78 B.n337 B.n336 585
R79 B.n338 B.n91 585
R80 B.n340 B.n339 585
R81 B.n341 B.n90 585
R82 B.n343 B.n342 585
R83 B.n344 B.n89 585
R84 B.n346 B.n345 585
R85 B.n347 B.n88 585
R86 B.n349 B.n348 585
R87 B.n350 B.n87 585
R88 B.n352 B.n351 585
R89 B.n353 B.n86 585
R90 B.n355 B.n354 585
R91 B.n356 B.n85 585
R92 B.n358 B.n357 585
R93 B.n359 B.n84 585
R94 B.n361 B.n360 585
R95 B.n362 B.n83 585
R96 B.n364 B.n363 585
R97 B.n365 B.n82 585
R98 B.n367 B.n366 585
R99 B.n368 B.n81 585
R100 B.n370 B.n369 585
R101 B.n371 B.n80 585
R102 B.n373 B.n372 585
R103 B.n374 B.n79 585
R104 B.n376 B.n375 585
R105 B.n377 B.n78 585
R106 B.n379 B.n378 585
R107 B.n380 B.n77 585
R108 B.n382 B.n381 585
R109 B.n383 B.n76 585
R110 B.n385 B.n384 585
R111 B.n386 B.n75 585
R112 B.n388 B.n387 585
R113 B.n389 B.n74 585
R114 B.n391 B.n390 585
R115 B.n392 B.n73 585
R116 B.n394 B.n393 585
R117 B.n395 B.n72 585
R118 B.n397 B.n396 585
R119 B.n398 B.n71 585
R120 B.n400 B.n399 585
R121 B.n401 B.n70 585
R122 B.n403 B.n402 585
R123 B.n404 B.n69 585
R124 B.n406 B.n405 585
R125 B.n407 B.n68 585
R126 B.n409 B.n408 585
R127 B.n410 B.n67 585
R128 B.n412 B.n411 585
R129 B.n413 B.n66 585
R130 B.n415 B.n414 585
R131 B.n416 B.n65 585
R132 B.n418 B.n417 585
R133 B.n419 B.n64 585
R134 B.n421 B.n420 585
R135 B.n422 B.n63 585
R136 B.n424 B.n423 585
R137 B.n425 B.n62 585
R138 B.n427 B.n426 585
R139 B.n428 B.n61 585
R140 B.n430 B.n429 585
R141 B.n431 B.n60 585
R142 B.n433 B.n432 585
R143 B.n434 B.n59 585
R144 B.n436 B.n435 585
R145 B.n437 B.n58 585
R146 B.n528 B.n23 585
R147 B.n527 B.n526 585
R148 B.n525 B.n24 585
R149 B.n524 B.n523 585
R150 B.n522 B.n25 585
R151 B.n521 B.n520 585
R152 B.n519 B.n26 585
R153 B.n518 B.n517 585
R154 B.n516 B.n27 585
R155 B.n515 B.n514 585
R156 B.n513 B.n28 585
R157 B.n512 B.n511 585
R158 B.n510 B.n29 585
R159 B.n509 B.n508 585
R160 B.n507 B.n30 585
R161 B.n506 B.n505 585
R162 B.n504 B.n31 585
R163 B.n503 B.n502 585
R164 B.n501 B.n32 585
R165 B.n500 B.n499 585
R166 B.n498 B.n33 585
R167 B.n497 B.n496 585
R168 B.n495 B.n34 585
R169 B.n494 B.n493 585
R170 B.n492 B.n35 585
R171 B.n490 B.n489 585
R172 B.n488 B.n38 585
R173 B.n487 B.n486 585
R174 B.n485 B.n39 585
R175 B.n484 B.n483 585
R176 B.n482 B.n40 585
R177 B.n481 B.n480 585
R178 B.n479 B.n41 585
R179 B.n478 B.n477 585
R180 B.n476 B.n42 585
R181 B.n475 B.n474 585
R182 B.n473 B.n43 585
R183 B.n472 B.n471 585
R184 B.n470 B.n47 585
R185 B.n469 B.n468 585
R186 B.n467 B.n48 585
R187 B.n466 B.n465 585
R188 B.n464 B.n49 585
R189 B.n463 B.n462 585
R190 B.n461 B.n50 585
R191 B.n460 B.n459 585
R192 B.n458 B.n51 585
R193 B.n457 B.n456 585
R194 B.n455 B.n52 585
R195 B.n454 B.n453 585
R196 B.n452 B.n53 585
R197 B.n451 B.n450 585
R198 B.n449 B.n54 585
R199 B.n448 B.n447 585
R200 B.n446 B.n55 585
R201 B.n445 B.n444 585
R202 B.n443 B.n56 585
R203 B.n442 B.n441 585
R204 B.n440 B.n57 585
R205 B.n439 B.n438 585
R206 B.n530 B.n529 585
R207 B.n531 B.n22 585
R208 B.n533 B.n532 585
R209 B.n534 B.n21 585
R210 B.n536 B.n535 585
R211 B.n537 B.n20 585
R212 B.n539 B.n538 585
R213 B.n540 B.n19 585
R214 B.n542 B.n541 585
R215 B.n543 B.n18 585
R216 B.n545 B.n544 585
R217 B.n546 B.n17 585
R218 B.n548 B.n547 585
R219 B.n549 B.n16 585
R220 B.n551 B.n550 585
R221 B.n552 B.n15 585
R222 B.n554 B.n553 585
R223 B.n555 B.n14 585
R224 B.n557 B.n556 585
R225 B.n558 B.n13 585
R226 B.n560 B.n559 585
R227 B.n561 B.n12 585
R228 B.n563 B.n562 585
R229 B.n564 B.n11 585
R230 B.n566 B.n565 585
R231 B.n567 B.n10 585
R232 B.n569 B.n568 585
R233 B.n570 B.n9 585
R234 B.n572 B.n571 585
R235 B.n573 B.n8 585
R236 B.n575 B.n574 585
R237 B.n576 B.n7 585
R238 B.n578 B.n577 585
R239 B.n579 B.n6 585
R240 B.n581 B.n580 585
R241 B.n582 B.n5 585
R242 B.n584 B.n583 585
R243 B.n585 B.n4 585
R244 B.n587 B.n586 585
R245 B.n588 B.n3 585
R246 B.n590 B.n589 585
R247 B.n591 B.n0 585
R248 B.n2 B.n1 585
R249 B.n154 B.n153 585
R250 B.n156 B.n155 585
R251 B.n157 B.n152 585
R252 B.n159 B.n158 585
R253 B.n160 B.n151 585
R254 B.n162 B.n161 585
R255 B.n163 B.n150 585
R256 B.n165 B.n164 585
R257 B.n166 B.n149 585
R258 B.n168 B.n167 585
R259 B.n169 B.n148 585
R260 B.n171 B.n170 585
R261 B.n172 B.n147 585
R262 B.n174 B.n173 585
R263 B.n175 B.n146 585
R264 B.n177 B.n176 585
R265 B.n178 B.n145 585
R266 B.n180 B.n179 585
R267 B.n181 B.n144 585
R268 B.n183 B.n182 585
R269 B.n184 B.n143 585
R270 B.n186 B.n185 585
R271 B.n187 B.n142 585
R272 B.n189 B.n188 585
R273 B.n190 B.n141 585
R274 B.n192 B.n191 585
R275 B.n193 B.n140 585
R276 B.n195 B.n194 585
R277 B.n196 B.n139 585
R278 B.n198 B.n197 585
R279 B.n199 B.n138 585
R280 B.n201 B.n200 585
R281 B.n202 B.n137 585
R282 B.n204 B.n203 585
R283 B.n205 B.n136 585
R284 B.n207 B.n206 585
R285 B.n208 B.n135 585
R286 B.n210 B.n209 585
R287 B.n211 B.n134 585
R288 B.n213 B.n212 585
R289 B.n214 B.n133 585
R290 B.n215 B.n214 554.963
R291 B.n309 B.n308 554.963
R292 B.n439 B.n58 554.963
R293 B.n530 B.n23 554.963
R294 B.n267 B.t1 352.526
R295 B.n44 B.t8 352.526
R296 B.n119 B.t4 352.526
R297 B.n36 B.t11 352.526
R298 B.n268 B.t2 276.695
R299 B.n45 B.t7 276.695
R300 B.n120 B.t5 276.695
R301 B.n37 B.t10 276.695
R302 B.n593 B.n592 256.663
R303 B.n119 B.t3 252.922
R304 B.n267 B.t0 252.922
R305 B.n44 B.t6 252.922
R306 B.n36 B.t9 252.922
R307 B.n592 B.n591 235.042
R308 B.n592 B.n2 235.042
R309 B.n215 B.n132 163.367
R310 B.n219 B.n132 163.367
R311 B.n220 B.n219 163.367
R312 B.n221 B.n220 163.367
R313 B.n221 B.n130 163.367
R314 B.n225 B.n130 163.367
R315 B.n226 B.n225 163.367
R316 B.n227 B.n226 163.367
R317 B.n227 B.n128 163.367
R318 B.n231 B.n128 163.367
R319 B.n232 B.n231 163.367
R320 B.n233 B.n232 163.367
R321 B.n233 B.n126 163.367
R322 B.n237 B.n126 163.367
R323 B.n238 B.n237 163.367
R324 B.n239 B.n238 163.367
R325 B.n239 B.n124 163.367
R326 B.n243 B.n124 163.367
R327 B.n244 B.n243 163.367
R328 B.n245 B.n244 163.367
R329 B.n245 B.n122 163.367
R330 B.n249 B.n122 163.367
R331 B.n250 B.n249 163.367
R332 B.n251 B.n250 163.367
R333 B.n251 B.n118 163.367
R334 B.n256 B.n118 163.367
R335 B.n257 B.n256 163.367
R336 B.n258 B.n257 163.367
R337 B.n258 B.n116 163.367
R338 B.n262 B.n116 163.367
R339 B.n263 B.n262 163.367
R340 B.n264 B.n263 163.367
R341 B.n264 B.n114 163.367
R342 B.n271 B.n114 163.367
R343 B.n272 B.n271 163.367
R344 B.n273 B.n272 163.367
R345 B.n273 B.n112 163.367
R346 B.n277 B.n112 163.367
R347 B.n278 B.n277 163.367
R348 B.n279 B.n278 163.367
R349 B.n279 B.n110 163.367
R350 B.n283 B.n110 163.367
R351 B.n284 B.n283 163.367
R352 B.n285 B.n284 163.367
R353 B.n285 B.n108 163.367
R354 B.n289 B.n108 163.367
R355 B.n290 B.n289 163.367
R356 B.n291 B.n290 163.367
R357 B.n291 B.n106 163.367
R358 B.n295 B.n106 163.367
R359 B.n296 B.n295 163.367
R360 B.n297 B.n296 163.367
R361 B.n297 B.n104 163.367
R362 B.n301 B.n104 163.367
R363 B.n302 B.n301 163.367
R364 B.n303 B.n302 163.367
R365 B.n303 B.n102 163.367
R366 B.n307 B.n102 163.367
R367 B.n308 B.n307 163.367
R368 B.n435 B.n58 163.367
R369 B.n435 B.n434 163.367
R370 B.n434 B.n433 163.367
R371 B.n433 B.n60 163.367
R372 B.n429 B.n60 163.367
R373 B.n429 B.n428 163.367
R374 B.n428 B.n427 163.367
R375 B.n427 B.n62 163.367
R376 B.n423 B.n62 163.367
R377 B.n423 B.n422 163.367
R378 B.n422 B.n421 163.367
R379 B.n421 B.n64 163.367
R380 B.n417 B.n64 163.367
R381 B.n417 B.n416 163.367
R382 B.n416 B.n415 163.367
R383 B.n415 B.n66 163.367
R384 B.n411 B.n66 163.367
R385 B.n411 B.n410 163.367
R386 B.n410 B.n409 163.367
R387 B.n409 B.n68 163.367
R388 B.n405 B.n68 163.367
R389 B.n405 B.n404 163.367
R390 B.n404 B.n403 163.367
R391 B.n403 B.n70 163.367
R392 B.n399 B.n70 163.367
R393 B.n399 B.n398 163.367
R394 B.n398 B.n397 163.367
R395 B.n397 B.n72 163.367
R396 B.n393 B.n72 163.367
R397 B.n393 B.n392 163.367
R398 B.n392 B.n391 163.367
R399 B.n391 B.n74 163.367
R400 B.n387 B.n74 163.367
R401 B.n387 B.n386 163.367
R402 B.n386 B.n385 163.367
R403 B.n385 B.n76 163.367
R404 B.n381 B.n76 163.367
R405 B.n381 B.n380 163.367
R406 B.n380 B.n379 163.367
R407 B.n379 B.n78 163.367
R408 B.n375 B.n78 163.367
R409 B.n375 B.n374 163.367
R410 B.n374 B.n373 163.367
R411 B.n373 B.n80 163.367
R412 B.n369 B.n80 163.367
R413 B.n369 B.n368 163.367
R414 B.n368 B.n367 163.367
R415 B.n367 B.n82 163.367
R416 B.n363 B.n82 163.367
R417 B.n363 B.n362 163.367
R418 B.n362 B.n361 163.367
R419 B.n361 B.n84 163.367
R420 B.n357 B.n84 163.367
R421 B.n357 B.n356 163.367
R422 B.n356 B.n355 163.367
R423 B.n355 B.n86 163.367
R424 B.n351 B.n86 163.367
R425 B.n351 B.n350 163.367
R426 B.n350 B.n349 163.367
R427 B.n349 B.n88 163.367
R428 B.n345 B.n88 163.367
R429 B.n345 B.n344 163.367
R430 B.n344 B.n343 163.367
R431 B.n343 B.n90 163.367
R432 B.n339 B.n90 163.367
R433 B.n339 B.n338 163.367
R434 B.n338 B.n337 163.367
R435 B.n337 B.n92 163.367
R436 B.n333 B.n92 163.367
R437 B.n333 B.n332 163.367
R438 B.n332 B.n331 163.367
R439 B.n331 B.n94 163.367
R440 B.n327 B.n94 163.367
R441 B.n327 B.n326 163.367
R442 B.n326 B.n325 163.367
R443 B.n325 B.n96 163.367
R444 B.n321 B.n96 163.367
R445 B.n321 B.n320 163.367
R446 B.n320 B.n319 163.367
R447 B.n319 B.n98 163.367
R448 B.n315 B.n98 163.367
R449 B.n315 B.n314 163.367
R450 B.n314 B.n313 163.367
R451 B.n313 B.n100 163.367
R452 B.n309 B.n100 163.367
R453 B.n526 B.n23 163.367
R454 B.n526 B.n525 163.367
R455 B.n525 B.n524 163.367
R456 B.n524 B.n25 163.367
R457 B.n520 B.n25 163.367
R458 B.n520 B.n519 163.367
R459 B.n519 B.n518 163.367
R460 B.n518 B.n27 163.367
R461 B.n514 B.n27 163.367
R462 B.n514 B.n513 163.367
R463 B.n513 B.n512 163.367
R464 B.n512 B.n29 163.367
R465 B.n508 B.n29 163.367
R466 B.n508 B.n507 163.367
R467 B.n507 B.n506 163.367
R468 B.n506 B.n31 163.367
R469 B.n502 B.n31 163.367
R470 B.n502 B.n501 163.367
R471 B.n501 B.n500 163.367
R472 B.n500 B.n33 163.367
R473 B.n496 B.n33 163.367
R474 B.n496 B.n495 163.367
R475 B.n495 B.n494 163.367
R476 B.n494 B.n35 163.367
R477 B.n489 B.n35 163.367
R478 B.n489 B.n488 163.367
R479 B.n488 B.n487 163.367
R480 B.n487 B.n39 163.367
R481 B.n483 B.n39 163.367
R482 B.n483 B.n482 163.367
R483 B.n482 B.n481 163.367
R484 B.n481 B.n41 163.367
R485 B.n477 B.n41 163.367
R486 B.n477 B.n476 163.367
R487 B.n476 B.n475 163.367
R488 B.n475 B.n43 163.367
R489 B.n471 B.n43 163.367
R490 B.n471 B.n470 163.367
R491 B.n470 B.n469 163.367
R492 B.n469 B.n48 163.367
R493 B.n465 B.n48 163.367
R494 B.n465 B.n464 163.367
R495 B.n464 B.n463 163.367
R496 B.n463 B.n50 163.367
R497 B.n459 B.n50 163.367
R498 B.n459 B.n458 163.367
R499 B.n458 B.n457 163.367
R500 B.n457 B.n52 163.367
R501 B.n453 B.n52 163.367
R502 B.n453 B.n452 163.367
R503 B.n452 B.n451 163.367
R504 B.n451 B.n54 163.367
R505 B.n447 B.n54 163.367
R506 B.n447 B.n446 163.367
R507 B.n446 B.n445 163.367
R508 B.n445 B.n56 163.367
R509 B.n441 B.n56 163.367
R510 B.n441 B.n440 163.367
R511 B.n440 B.n439 163.367
R512 B.n531 B.n530 163.367
R513 B.n532 B.n531 163.367
R514 B.n532 B.n21 163.367
R515 B.n536 B.n21 163.367
R516 B.n537 B.n536 163.367
R517 B.n538 B.n537 163.367
R518 B.n538 B.n19 163.367
R519 B.n542 B.n19 163.367
R520 B.n543 B.n542 163.367
R521 B.n544 B.n543 163.367
R522 B.n544 B.n17 163.367
R523 B.n548 B.n17 163.367
R524 B.n549 B.n548 163.367
R525 B.n550 B.n549 163.367
R526 B.n550 B.n15 163.367
R527 B.n554 B.n15 163.367
R528 B.n555 B.n554 163.367
R529 B.n556 B.n555 163.367
R530 B.n556 B.n13 163.367
R531 B.n560 B.n13 163.367
R532 B.n561 B.n560 163.367
R533 B.n562 B.n561 163.367
R534 B.n562 B.n11 163.367
R535 B.n566 B.n11 163.367
R536 B.n567 B.n566 163.367
R537 B.n568 B.n567 163.367
R538 B.n568 B.n9 163.367
R539 B.n572 B.n9 163.367
R540 B.n573 B.n572 163.367
R541 B.n574 B.n573 163.367
R542 B.n574 B.n7 163.367
R543 B.n578 B.n7 163.367
R544 B.n579 B.n578 163.367
R545 B.n580 B.n579 163.367
R546 B.n580 B.n5 163.367
R547 B.n584 B.n5 163.367
R548 B.n585 B.n584 163.367
R549 B.n586 B.n585 163.367
R550 B.n586 B.n3 163.367
R551 B.n590 B.n3 163.367
R552 B.n591 B.n590 163.367
R553 B.n154 B.n2 163.367
R554 B.n155 B.n154 163.367
R555 B.n155 B.n152 163.367
R556 B.n159 B.n152 163.367
R557 B.n160 B.n159 163.367
R558 B.n161 B.n160 163.367
R559 B.n161 B.n150 163.367
R560 B.n165 B.n150 163.367
R561 B.n166 B.n165 163.367
R562 B.n167 B.n166 163.367
R563 B.n167 B.n148 163.367
R564 B.n171 B.n148 163.367
R565 B.n172 B.n171 163.367
R566 B.n173 B.n172 163.367
R567 B.n173 B.n146 163.367
R568 B.n177 B.n146 163.367
R569 B.n178 B.n177 163.367
R570 B.n179 B.n178 163.367
R571 B.n179 B.n144 163.367
R572 B.n183 B.n144 163.367
R573 B.n184 B.n183 163.367
R574 B.n185 B.n184 163.367
R575 B.n185 B.n142 163.367
R576 B.n189 B.n142 163.367
R577 B.n190 B.n189 163.367
R578 B.n191 B.n190 163.367
R579 B.n191 B.n140 163.367
R580 B.n195 B.n140 163.367
R581 B.n196 B.n195 163.367
R582 B.n197 B.n196 163.367
R583 B.n197 B.n138 163.367
R584 B.n201 B.n138 163.367
R585 B.n202 B.n201 163.367
R586 B.n203 B.n202 163.367
R587 B.n203 B.n136 163.367
R588 B.n207 B.n136 163.367
R589 B.n208 B.n207 163.367
R590 B.n209 B.n208 163.367
R591 B.n209 B.n134 163.367
R592 B.n213 B.n134 163.367
R593 B.n214 B.n213 163.367
R594 B.n120 B.n119 75.8308
R595 B.n268 B.n267 75.8308
R596 B.n45 B.n44 75.8308
R597 B.n37 B.n36 75.8308
R598 B.n253 B.n120 59.5399
R599 B.n269 B.n268 59.5399
R600 B.n46 B.n45 59.5399
R601 B.n491 B.n37 59.5399
R602 B.n529 B.n528 36.059
R603 B.n438 B.n437 36.059
R604 B.n216 B.n133 36.059
R605 B.n310 B.n101 36.059
R606 B B.n593 18.0485
R607 B.n529 B.n22 10.6151
R608 B.n533 B.n22 10.6151
R609 B.n534 B.n533 10.6151
R610 B.n535 B.n534 10.6151
R611 B.n535 B.n20 10.6151
R612 B.n539 B.n20 10.6151
R613 B.n540 B.n539 10.6151
R614 B.n541 B.n540 10.6151
R615 B.n541 B.n18 10.6151
R616 B.n545 B.n18 10.6151
R617 B.n546 B.n545 10.6151
R618 B.n547 B.n546 10.6151
R619 B.n547 B.n16 10.6151
R620 B.n551 B.n16 10.6151
R621 B.n552 B.n551 10.6151
R622 B.n553 B.n552 10.6151
R623 B.n553 B.n14 10.6151
R624 B.n557 B.n14 10.6151
R625 B.n558 B.n557 10.6151
R626 B.n559 B.n558 10.6151
R627 B.n559 B.n12 10.6151
R628 B.n563 B.n12 10.6151
R629 B.n564 B.n563 10.6151
R630 B.n565 B.n564 10.6151
R631 B.n565 B.n10 10.6151
R632 B.n569 B.n10 10.6151
R633 B.n570 B.n569 10.6151
R634 B.n571 B.n570 10.6151
R635 B.n571 B.n8 10.6151
R636 B.n575 B.n8 10.6151
R637 B.n576 B.n575 10.6151
R638 B.n577 B.n576 10.6151
R639 B.n577 B.n6 10.6151
R640 B.n581 B.n6 10.6151
R641 B.n582 B.n581 10.6151
R642 B.n583 B.n582 10.6151
R643 B.n583 B.n4 10.6151
R644 B.n587 B.n4 10.6151
R645 B.n588 B.n587 10.6151
R646 B.n589 B.n588 10.6151
R647 B.n589 B.n0 10.6151
R648 B.n528 B.n527 10.6151
R649 B.n527 B.n24 10.6151
R650 B.n523 B.n24 10.6151
R651 B.n523 B.n522 10.6151
R652 B.n522 B.n521 10.6151
R653 B.n521 B.n26 10.6151
R654 B.n517 B.n26 10.6151
R655 B.n517 B.n516 10.6151
R656 B.n516 B.n515 10.6151
R657 B.n515 B.n28 10.6151
R658 B.n511 B.n28 10.6151
R659 B.n511 B.n510 10.6151
R660 B.n510 B.n509 10.6151
R661 B.n509 B.n30 10.6151
R662 B.n505 B.n30 10.6151
R663 B.n505 B.n504 10.6151
R664 B.n504 B.n503 10.6151
R665 B.n503 B.n32 10.6151
R666 B.n499 B.n32 10.6151
R667 B.n499 B.n498 10.6151
R668 B.n498 B.n497 10.6151
R669 B.n497 B.n34 10.6151
R670 B.n493 B.n34 10.6151
R671 B.n493 B.n492 10.6151
R672 B.n490 B.n38 10.6151
R673 B.n486 B.n38 10.6151
R674 B.n486 B.n485 10.6151
R675 B.n485 B.n484 10.6151
R676 B.n484 B.n40 10.6151
R677 B.n480 B.n40 10.6151
R678 B.n480 B.n479 10.6151
R679 B.n479 B.n478 10.6151
R680 B.n478 B.n42 10.6151
R681 B.n474 B.n473 10.6151
R682 B.n473 B.n472 10.6151
R683 B.n472 B.n47 10.6151
R684 B.n468 B.n47 10.6151
R685 B.n468 B.n467 10.6151
R686 B.n467 B.n466 10.6151
R687 B.n466 B.n49 10.6151
R688 B.n462 B.n49 10.6151
R689 B.n462 B.n461 10.6151
R690 B.n461 B.n460 10.6151
R691 B.n460 B.n51 10.6151
R692 B.n456 B.n51 10.6151
R693 B.n456 B.n455 10.6151
R694 B.n455 B.n454 10.6151
R695 B.n454 B.n53 10.6151
R696 B.n450 B.n53 10.6151
R697 B.n450 B.n449 10.6151
R698 B.n449 B.n448 10.6151
R699 B.n448 B.n55 10.6151
R700 B.n444 B.n55 10.6151
R701 B.n444 B.n443 10.6151
R702 B.n443 B.n442 10.6151
R703 B.n442 B.n57 10.6151
R704 B.n438 B.n57 10.6151
R705 B.n437 B.n436 10.6151
R706 B.n436 B.n59 10.6151
R707 B.n432 B.n59 10.6151
R708 B.n432 B.n431 10.6151
R709 B.n431 B.n430 10.6151
R710 B.n430 B.n61 10.6151
R711 B.n426 B.n61 10.6151
R712 B.n426 B.n425 10.6151
R713 B.n425 B.n424 10.6151
R714 B.n424 B.n63 10.6151
R715 B.n420 B.n63 10.6151
R716 B.n420 B.n419 10.6151
R717 B.n419 B.n418 10.6151
R718 B.n418 B.n65 10.6151
R719 B.n414 B.n65 10.6151
R720 B.n414 B.n413 10.6151
R721 B.n413 B.n412 10.6151
R722 B.n412 B.n67 10.6151
R723 B.n408 B.n67 10.6151
R724 B.n408 B.n407 10.6151
R725 B.n407 B.n406 10.6151
R726 B.n406 B.n69 10.6151
R727 B.n402 B.n69 10.6151
R728 B.n402 B.n401 10.6151
R729 B.n401 B.n400 10.6151
R730 B.n400 B.n71 10.6151
R731 B.n396 B.n71 10.6151
R732 B.n396 B.n395 10.6151
R733 B.n395 B.n394 10.6151
R734 B.n394 B.n73 10.6151
R735 B.n390 B.n73 10.6151
R736 B.n390 B.n389 10.6151
R737 B.n389 B.n388 10.6151
R738 B.n388 B.n75 10.6151
R739 B.n384 B.n75 10.6151
R740 B.n384 B.n383 10.6151
R741 B.n383 B.n382 10.6151
R742 B.n382 B.n77 10.6151
R743 B.n378 B.n77 10.6151
R744 B.n378 B.n377 10.6151
R745 B.n377 B.n376 10.6151
R746 B.n376 B.n79 10.6151
R747 B.n372 B.n79 10.6151
R748 B.n372 B.n371 10.6151
R749 B.n371 B.n370 10.6151
R750 B.n370 B.n81 10.6151
R751 B.n366 B.n81 10.6151
R752 B.n366 B.n365 10.6151
R753 B.n365 B.n364 10.6151
R754 B.n364 B.n83 10.6151
R755 B.n360 B.n83 10.6151
R756 B.n360 B.n359 10.6151
R757 B.n359 B.n358 10.6151
R758 B.n358 B.n85 10.6151
R759 B.n354 B.n85 10.6151
R760 B.n354 B.n353 10.6151
R761 B.n353 B.n352 10.6151
R762 B.n352 B.n87 10.6151
R763 B.n348 B.n87 10.6151
R764 B.n348 B.n347 10.6151
R765 B.n347 B.n346 10.6151
R766 B.n346 B.n89 10.6151
R767 B.n342 B.n89 10.6151
R768 B.n342 B.n341 10.6151
R769 B.n341 B.n340 10.6151
R770 B.n340 B.n91 10.6151
R771 B.n336 B.n91 10.6151
R772 B.n336 B.n335 10.6151
R773 B.n335 B.n334 10.6151
R774 B.n334 B.n93 10.6151
R775 B.n330 B.n93 10.6151
R776 B.n330 B.n329 10.6151
R777 B.n329 B.n328 10.6151
R778 B.n328 B.n95 10.6151
R779 B.n324 B.n95 10.6151
R780 B.n324 B.n323 10.6151
R781 B.n323 B.n322 10.6151
R782 B.n322 B.n97 10.6151
R783 B.n318 B.n97 10.6151
R784 B.n318 B.n317 10.6151
R785 B.n317 B.n316 10.6151
R786 B.n316 B.n99 10.6151
R787 B.n312 B.n99 10.6151
R788 B.n312 B.n311 10.6151
R789 B.n311 B.n310 10.6151
R790 B.n153 B.n1 10.6151
R791 B.n156 B.n153 10.6151
R792 B.n157 B.n156 10.6151
R793 B.n158 B.n157 10.6151
R794 B.n158 B.n151 10.6151
R795 B.n162 B.n151 10.6151
R796 B.n163 B.n162 10.6151
R797 B.n164 B.n163 10.6151
R798 B.n164 B.n149 10.6151
R799 B.n168 B.n149 10.6151
R800 B.n169 B.n168 10.6151
R801 B.n170 B.n169 10.6151
R802 B.n170 B.n147 10.6151
R803 B.n174 B.n147 10.6151
R804 B.n175 B.n174 10.6151
R805 B.n176 B.n175 10.6151
R806 B.n176 B.n145 10.6151
R807 B.n180 B.n145 10.6151
R808 B.n181 B.n180 10.6151
R809 B.n182 B.n181 10.6151
R810 B.n182 B.n143 10.6151
R811 B.n186 B.n143 10.6151
R812 B.n187 B.n186 10.6151
R813 B.n188 B.n187 10.6151
R814 B.n188 B.n141 10.6151
R815 B.n192 B.n141 10.6151
R816 B.n193 B.n192 10.6151
R817 B.n194 B.n193 10.6151
R818 B.n194 B.n139 10.6151
R819 B.n198 B.n139 10.6151
R820 B.n199 B.n198 10.6151
R821 B.n200 B.n199 10.6151
R822 B.n200 B.n137 10.6151
R823 B.n204 B.n137 10.6151
R824 B.n205 B.n204 10.6151
R825 B.n206 B.n205 10.6151
R826 B.n206 B.n135 10.6151
R827 B.n210 B.n135 10.6151
R828 B.n211 B.n210 10.6151
R829 B.n212 B.n211 10.6151
R830 B.n212 B.n133 10.6151
R831 B.n217 B.n216 10.6151
R832 B.n218 B.n217 10.6151
R833 B.n218 B.n131 10.6151
R834 B.n222 B.n131 10.6151
R835 B.n223 B.n222 10.6151
R836 B.n224 B.n223 10.6151
R837 B.n224 B.n129 10.6151
R838 B.n228 B.n129 10.6151
R839 B.n229 B.n228 10.6151
R840 B.n230 B.n229 10.6151
R841 B.n230 B.n127 10.6151
R842 B.n234 B.n127 10.6151
R843 B.n235 B.n234 10.6151
R844 B.n236 B.n235 10.6151
R845 B.n236 B.n125 10.6151
R846 B.n240 B.n125 10.6151
R847 B.n241 B.n240 10.6151
R848 B.n242 B.n241 10.6151
R849 B.n242 B.n123 10.6151
R850 B.n246 B.n123 10.6151
R851 B.n247 B.n246 10.6151
R852 B.n248 B.n247 10.6151
R853 B.n248 B.n121 10.6151
R854 B.n252 B.n121 10.6151
R855 B.n255 B.n254 10.6151
R856 B.n255 B.n117 10.6151
R857 B.n259 B.n117 10.6151
R858 B.n260 B.n259 10.6151
R859 B.n261 B.n260 10.6151
R860 B.n261 B.n115 10.6151
R861 B.n265 B.n115 10.6151
R862 B.n266 B.n265 10.6151
R863 B.n270 B.n266 10.6151
R864 B.n274 B.n113 10.6151
R865 B.n275 B.n274 10.6151
R866 B.n276 B.n275 10.6151
R867 B.n276 B.n111 10.6151
R868 B.n280 B.n111 10.6151
R869 B.n281 B.n280 10.6151
R870 B.n282 B.n281 10.6151
R871 B.n282 B.n109 10.6151
R872 B.n286 B.n109 10.6151
R873 B.n287 B.n286 10.6151
R874 B.n288 B.n287 10.6151
R875 B.n288 B.n107 10.6151
R876 B.n292 B.n107 10.6151
R877 B.n293 B.n292 10.6151
R878 B.n294 B.n293 10.6151
R879 B.n294 B.n105 10.6151
R880 B.n298 B.n105 10.6151
R881 B.n299 B.n298 10.6151
R882 B.n300 B.n299 10.6151
R883 B.n300 B.n103 10.6151
R884 B.n304 B.n103 10.6151
R885 B.n305 B.n304 10.6151
R886 B.n306 B.n305 10.6151
R887 B.n306 B.n101 10.6151
R888 B.n492 B.n491 9.36635
R889 B.n474 B.n46 9.36635
R890 B.n253 B.n252 9.36635
R891 B.n269 B.n113 9.36635
R892 B.n593 B.n0 8.11757
R893 B.n593 B.n1 8.11757
R894 B.n491 B.n490 1.24928
R895 B.n46 B.n42 1.24928
R896 B.n254 B.n253 1.24928
R897 B.n270 B.n269 1.24928
R898 VP.n19 VP.n18 161.3
R899 VP.n17 VP.n1 161.3
R900 VP.n16 VP.n15 161.3
R901 VP.n14 VP.n2 161.3
R902 VP.n13 VP.n12 161.3
R903 VP.n11 VP.n3 161.3
R904 VP.n10 VP.n9 161.3
R905 VP.n8 VP.n4 161.3
R906 VP.n7 VP.n6 80.1629
R907 VP.n20 VP.n0 80.1629
R908 VP.n5 VP.t1 78.629
R909 VP.n5 VP.t3 77.3889
R910 VP.n12 VP.n2 56.5617
R911 VP.n7 VP.n5 47.3439
R912 VP.n6 VP.t2 43.7575
R913 VP.n0 VP.t0 43.7575
R914 VP.n10 VP.n4 24.5923
R915 VP.n11 VP.n10 24.5923
R916 VP.n12 VP.n11 24.5923
R917 VP.n16 VP.n2 24.5923
R918 VP.n17 VP.n16 24.5923
R919 VP.n18 VP.n17 24.5923
R920 VP.n6 VP.n4 10.0832
R921 VP.n18 VP.n0 10.0832
R922 VP.n8 VP.n7 0.354861
R923 VP.n20 VP.n19 0.354861
R924 VP VP.n20 0.267071
R925 VP.n9 VP.n8 0.189894
R926 VP.n9 VP.n3 0.189894
R927 VP.n13 VP.n3 0.189894
R928 VP.n14 VP.n13 0.189894
R929 VP.n15 VP.n14 0.189894
R930 VP.n15 VP.n1 0.189894
R931 VP.n19 VP.n1 0.189894
R932 VTAIL.n270 VTAIL.n269 756.745
R933 VTAIL.n32 VTAIL.n31 756.745
R934 VTAIL.n66 VTAIL.n65 756.745
R935 VTAIL.n100 VTAIL.n99 756.745
R936 VTAIL.n236 VTAIL.n235 756.745
R937 VTAIL.n202 VTAIL.n201 756.745
R938 VTAIL.n168 VTAIL.n167 756.745
R939 VTAIL.n134 VTAIL.n133 756.745
R940 VTAIL.n248 VTAIL.n247 585
R941 VTAIL.n253 VTAIL.n252 585
R942 VTAIL.n255 VTAIL.n254 585
R943 VTAIL.n244 VTAIL.n243 585
R944 VTAIL.n261 VTAIL.n260 585
R945 VTAIL.n263 VTAIL.n262 585
R946 VTAIL.n240 VTAIL.n239 585
R947 VTAIL.n269 VTAIL.n268 585
R948 VTAIL.n10 VTAIL.n9 585
R949 VTAIL.n15 VTAIL.n14 585
R950 VTAIL.n17 VTAIL.n16 585
R951 VTAIL.n6 VTAIL.n5 585
R952 VTAIL.n23 VTAIL.n22 585
R953 VTAIL.n25 VTAIL.n24 585
R954 VTAIL.n2 VTAIL.n1 585
R955 VTAIL.n31 VTAIL.n30 585
R956 VTAIL.n44 VTAIL.n43 585
R957 VTAIL.n49 VTAIL.n48 585
R958 VTAIL.n51 VTAIL.n50 585
R959 VTAIL.n40 VTAIL.n39 585
R960 VTAIL.n57 VTAIL.n56 585
R961 VTAIL.n59 VTAIL.n58 585
R962 VTAIL.n36 VTAIL.n35 585
R963 VTAIL.n65 VTAIL.n64 585
R964 VTAIL.n78 VTAIL.n77 585
R965 VTAIL.n83 VTAIL.n82 585
R966 VTAIL.n85 VTAIL.n84 585
R967 VTAIL.n74 VTAIL.n73 585
R968 VTAIL.n91 VTAIL.n90 585
R969 VTAIL.n93 VTAIL.n92 585
R970 VTAIL.n70 VTAIL.n69 585
R971 VTAIL.n99 VTAIL.n98 585
R972 VTAIL.n235 VTAIL.n234 585
R973 VTAIL.n206 VTAIL.n205 585
R974 VTAIL.n229 VTAIL.n228 585
R975 VTAIL.n227 VTAIL.n226 585
R976 VTAIL.n210 VTAIL.n209 585
R977 VTAIL.n221 VTAIL.n220 585
R978 VTAIL.n219 VTAIL.n218 585
R979 VTAIL.n214 VTAIL.n213 585
R980 VTAIL.n201 VTAIL.n200 585
R981 VTAIL.n172 VTAIL.n171 585
R982 VTAIL.n195 VTAIL.n194 585
R983 VTAIL.n193 VTAIL.n192 585
R984 VTAIL.n176 VTAIL.n175 585
R985 VTAIL.n187 VTAIL.n186 585
R986 VTAIL.n185 VTAIL.n184 585
R987 VTAIL.n180 VTAIL.n179 585
R988 VTAIL.n167 VTAIL.n166 585
R989 VTAIL.n138 VTAIL.n137 585
R990 VTAIL.n161 VTAIL.n160 585
R991 VTAIL.n159 VTAIL.n158 585
R992 VTAIL.n142 VTAIL.n141 585
R993 VTAIL.n153 VTAIL.n152 585
R994 VTAIL.n151 VTAIL.n150 585
R995 VTAIL.n146 VTAIL.n145 585
R996 VTAIL.n133 VTAIL.n132 585
R997 VTAIL.n104 VTAIL.n103 585
R998 VTAIL.n127 VTAIL.n126 585
R999 VTAIL.n125 VTAIL.n124 585
R1000 VTAIL.n108 VTAIL.n107 585
R1001 VTAIL.n119 VTAIL.n118 585
R1002 VTAIL.n117 VTAIL.n116 585
R1003 VTAIL.n112 VTAIL.n111 585
R1004 VTAIL.n249 VTAIL.t3 329.084
R1005 VTAIL.n11 VTAIL.t2 329.084
R1006 VTAIL.n45 VTAIL.t4 329.084
R1007 VTAIL.n79 VTAIL.t6 329.084
R1008 VTAIL.n215 VTAIL.t7 329.084
R1009 VTAIL.n181 VTAIL.t5 329.084
R1010 VTAIL.n147 VTAIL.t1 329.084
R1011 VTAIL.n113 VTAIL.t0 329.084
R1012 VTAIL.n253 VTAIL.n247 171.744
R1013 VTAIL.n254 VTAIL.n253 171.744
R1014 VTAIL.n254 VTAIL.n243 171.744
R1015 VTAIL.n261 VTAIL.n243 171.744
R1016 VTAIL.n262 VTAIL.n261 171.744
R1017 VTAIL.n262 VTAIL.n239 171.744
R1018 VTAIL.n269 VTAIL.n239 171.744
R1019 VTAIL.n15 VTAIL.n9 171.744
R1020 VTAIL.n16 VTAIL.n15 171.744
R1021 VTAIL.n16 VTAIL.n5 171.744
R1022 VTAIL.n23 VTAIL.n5 171.744
R1023 VTAIL.n24 VTAIL.n23 171.744
R1024 VTAIL.n24 VTAIL.n1 171.744
R1025 VTAIL.n31 VTAIL.n1 171.744
R1026 VTAIL.n49 VTAIL.n43 171.744
R1027 VTAIL.n50 VTAIL.n49 171.744
R1028 VTAIL.n50 VTAIL.n39 171.744
R1029 VTAIL.n57 VTAIL.n39 171.744
R1030 VTAIL.n58 VTAIL.n57 171.744
R1031 VTAIL.n58 VTAIL.n35 171.744
R1032 VTAIL.n65 VTAIL.n35 171.744
R1033 VTAIL.n83 VTAIL.n77 171.744
R1034 VTAIL.n84 VTAIL.n83 171.744
R1035 VTAIL.n84 VTAIL.n73 171.744
R1036 VTAIL.n91 VTAIL.n73 171.744
R1037 VTAIL.n92 VTAIL.n91 171.744
R1038 VTAIL.n92 VTAIL.n69 171.744
R1039 VTAIL.n99 VTAIL.n69 171.744
R1040 VTAIL.n235 VTAIL.n205 171.744
R1041 VTAIL.n228 VTAIL.n205 171.744
R1042 VTAIL.n228 VTAIL.n227 171.744
R1043 VTAIL.n227 VTAIL.n209 171.744
R1044 VTAIL.n220 VTAIL.n209 171.744
R1045 VTAIL.n220 VTAIL.n219 171.744
R1046 VTAIL.n219 VTAIL.n213 171.744
R1047 VTAIL.n201 VTAIL.n171 171.744
R1048 VTAIL.n194 VTAIL.n171 171.744
R1049 VTAIL.n194 VTAIL.n193 171.744
R1050 VTAIL.n193 VTAIL.n175 171.744
R1051 VTAIL.n186 VTAIL.n175 171.744
R1052 VTAIL.n186 VTAIL.n185 171.744
R1053 VTAIL.n185 VTAIL.n179 171.744
R1054 VTAIL.n167 VTAIL.n137 171.744
R1055 VTAIL.n160 VTAIL.n137 171.744
R1056 VTAIL.n160 VTAIL.n159 171.744
R1057 VTAIL.n159 VTAIL.n141 171.744
R1058 VTAIL.n152 VTAIL.n141 171.744
R1059 VTAIL.n152 VTAIL.n151 171.744
R1060 VTAIL.n151 VTAIL.n145 171.744
R1061 VTAIL.n133 VTAIL.n103 171.744
R1062 VTAIL.n126 VTAIL.n103 171.744
R1063 VTAIL.n126 VTAIL.n125 171.744
R1064 VTAIL.n125 VTAIL.n107 171.744
R1065 VTAIL.n118 VTAIL.n107 171.744
R1066 VTAIL.n118 VTAIL.n117 171.744
R1067 VTAIL.n117 VTAIL.n111 171.744
R1068 VTAIL.t3 VTAIL.n247 85.8723
R1069 VTAIL.t2 VTAIL.n9 85.8723
R1070 VTAIL.t4 VTAIL.n43 85.8723
R1071 VTAIL.t6 VTAIL.n77 85.8723
R1072 VTAIL.t7 VTAIL.n213 85.8723
R1073 VTAIL.t5 VTAIL.n179 85.8723
R1074 VTAIL.t1 VTAIL.n145 85.8723
R1075 VTAIL.t0 VTAIL.n111 85.8723
R1076 VTAIL.n271 VTAIL.n270 34.5126
R1077 VTAIL.n33 VTAIL.n32 34.5126
R1078 VTAIL.n67 VTAIL.n66 34.5126
R1079 VTAIL.n101 VTAIL.n100 34.5126
R1080 VTAIL.n237 VTAIL.n236 34.5126
R1081 VTAIL.n203 VTAIL.n202 34.5126
R1082 VTAIL.n169 VTAIL.n168 34.5126
R1083 VTAIL.n135 VTAIL.n134 34.5126
R1084 VTAIL.n271 VTAIL.n237 21.341
R1085 VTAIL.n135 VTAIL.n101 21.341
R1086 VTAIL.n268 VTAIL.n238 12.8005
R1087 VTAIL.n30 VTAIL.n0 12.8005
R1088 VTAIL.n64 VTAIL.n34 12.8005
R1089 VTAIL.n98 VTAIL.n68 12.8005
R1090 VTAIL.n234 VTAIL.n204 12.8005
R1091 VTAIL.n200 VTAIL.n170 12.8005
R1092 VTAIL.n166 VTAIL.n136 12.8005
R1093 VTAIL.n132 VTAIL.n102 12.8005
R1094 VTAIL.n267 VTAIL.n240 12.0247
R1095 VTAIL.n29 VTAIL.n2 12.0247
R1096 VTAIL.n63 VTAIL.n36 12.0247
R1097 VTAIL.n97 VTAIL.n70 12.0247
R1098 VTAIL.n233 VTAIL.n206 12.0247
R1099 VTAIL.n199 VTAIL.n172 12.0247
R1100 VTAIL.n165 VTAIL.n138 12.0247
R1101 VTAIL.n131 VTAIL.n104 12.0247
R1102 VTAIL.n264 VTAIL.n263 11.249
R1103 VTAIL.n26 VTAIL.n25 11.249
R1104 VTAIL.n60 VTAIL.n59 11.249
R1105 VTAIL.n94 VTAIL.n93 11.249
R1106 VTAIL.n230 VTAIL.n229 11.249
R1107 VTAIL.n196 VTAIL.n195 11.249
R1108 VTAIL.n162 VTAIL.n161 11.249
R1109 VTAIL.n128 VTAIL.n127 11.249
R1110 VTAIL.n249 VTAIL.n248 10.7233
R1111 VTAIL.n11 VTAIL.n10 10.7233
R1112 VTAIL.n45 VTAIL.n44 10.7233
R1113 VTAIL.n79 VTAIL.n78 10.7233
R1114 VTAIL.n215 VTAIL.n214 10.7233
R1115 VTAIL.n181 VTAIL.n180 10.7233
R1116 VTAIL.n147 VTAIL.n146 10.7233
R1117 VTAIL.n113 VTAIL.n112 10.7233
R1118 VTAIL.n260 VTAIL.n242 10.4732
R1119 VTAIL.n22 VTAIL.n4 10.4732
R1120 VTAIL.n56 VTAIL.n38 10.4732
R1121 VTAIL.n90 VTAIL.n72 10.4732
R1122 VTAIL.n226 VTAIL.n208 10.4732
R1123 VTAIL.n192 VTAIL.n174 10.4732
R1124 VTAIL.n158 VTAIL.n140 10.4732
R1125 VTAIL.n124 VTAIL.n106 10.4732
R1126 VTAIL.n259 VTAIL.n244 9.69747
R1127 VTAIL.n21 VTAIL.n6 9.69747
R1128 VTAIL.n55 VTAIL.n40 9.69747
R1129 VTAIL.n89 VTAIL.n74 9.69747
R1130 VTAIL.n225 VTAIL.n210 9.69747
R1131 VTAIL.n191 VTAIL.n176 9.69747
R1132 VTAIL.n157 VTAIL.n142 9.69747
R1133 VTAIL.n123 VTAIL.n108 9.69747
R1134 VTAIL.n266 VTAIL.n238 9.45567
R1135 VTAIL.n28 VTAIL.n0 9.45567
R1136 VTAIL.n62 VTAIL.n34 9.45567
R1137 VTAIL.n96 VTAIL.n68 9.45567
R1138 VTAIL.n232 VTAIL.n204 9.45567
R1139 VTAIL.n198 VTAIL.n170 9.45567
R1140 VTAIL.n164 VTAIL.n136 9.45567
R1141 VTAIL.n130 VTAIL.n102 9.45567
R1142 VTAIL.n251 VTAIL.n250 9.3005
R1143 VTAIL.n246 VTAIL.n245 9.3005
R1144 VTAIL.n257 VTAIL.n256 9.3005
R1145 VTAIL.n259 VTAIL.n258 9.3005
R1146 VTAIL.n242 VTAIL.n241 9.3005
R1147 VTAIL.n265 VTAIL.n264 9.3005
R1148 VTAIL.n267 VTAIL.n266 9.3005
R1149 VTAIL.n13 VTAIL.n12 9.3005
R1150 VTAIL.n8 VTAIL.n7 9.3005
R1151 VTAIL.n19 VTAIL.n18 9.3005
R1152 VTAIL.n21 VTAIL.n20 9.3005
R1153 VTAIL.n4 VTAIL.n3 9.3005
R1154 VTAIL.n27 VTAIL.n26 9.3005
R1155 VTAIL.n29 VTAIL.n28 9.3005
R1156 VTAIL.n47 VTAIL.n46 9.3005
R1157 VTAIL.n42 VTAIL.n41 9.3005
R1158 VTAIL.n53 VTAIL.n52 9.3005
R1159 VTAIL.n55 VTAIL.n54 9.3005
R1160 VTAIL.n38 VTAIL.n37 9.3005
R1161 VTAIL.n61 VTAIL.n60 9.3005
R1162 VTAIL.n63 VTAIL.n62 9.3005
R1163 VTAIL.n81 VTAIL.n80 9.3005
R1164 VTAIL.n76 VTAIL.n75 9.3005
R1165 VTAIL.n87 VTAIL.n86 9.3005
R1166 VTAIL.n89 VTAIL.n88 9.3005
R1167 VTAIL.n72 VTAIL.n71 9.3005
R1168 VTAIL.n95 VTAIL.n94 9.3005
R1169 VTAIL.n97 VTAIL.n96 9.3005
R1170 VTAIL.n233 VTAIL.n232 9.3005
R1171 VTAIL.n231 VTAIL.n230 9.3005
R1172 VTAIL.n208 VTAIL.n207 9.3005
R1173 VTAIL.n225 VTAIL.n224 9.3005
R1174 VTAIL.n223 VTAIL.n222 9.3005
R1175 VTAIL.n212 VTAIL.n211 9.3005
R1176 VTAIL.n217 VTAIL.n216 9.3005
R1177 VTAIL.n178 VTAIL.n177 9.3005
R1178 VTAIL.n189 VTAIL.n188 9.3005
R1179 VTAIL.n191 VTAIL.n190 9.3005
R1180 VTAIL.n174 VTAIL.n173 9.3005
R1181 VTAIL.n197 VTAIL.n196 9.3005
R1182 VTAIL.n199 VTAIL.n198 9.3005
R1183 VTAIL.n183 VTAIL.n182 9.3005
R1184 VTAIL.n144 VTAIL.n143 9.3005
R1185 VTAIL.n155 VTAIL.n154 9.3005
R1186 VTAIL.n157 VTAIL.n156 9.3005
R1187 VTAIL.n140 VTAIL.n139 9.3005
R1188 VTAIL.n163 VTAIL.n162 9.3005
R1189 VTAIL.n165 VTAIL.n164 9.3005
R1190 VTAIL.n149 VTAIL.n148 9.3005
R1191 VTAIL.n110 VTAIL.n109 9.3005
R1192 VTAIL.n121 VTAIL.n120 9.3005
R1193 VTAIL.n123 VTAIL.n122 9.3005
R1194 VTAIL.n106 VTAIL.n105 9.3005
R1195 VTAIL.n129 VTAIL.n128 9.3005
R1196 VTAIL.n131 VTAIL.n130 9.3005
R1197 VTAIL.n115 VTAIL.n114 9.3005
R1198 VTAIL.n256 VTAIL.n255 8.92171
R1199 VTAIL.n18 VTAIL.n17 8.92171
R1200 VTAIL.n52 VTAIL.n51 8.92171
R1201 VTAIL.n86 VTAIL.n85 8.92171
R1202 VTAIL.n222 VTAIL.n221 8.92171
R1203 VTAIL.n188 VTAIL.n187 8.92171
R1204 VTAIL.n154 VTAIL.n153 8.92171
R1205 VTAIL.n120 VTAIL.n119 8.92171
R1206 VTAIL.n252 VTAIL.n246 8.14595
R1207 VTAIL.n14 VTAIL.n8 8.14595
R1208 VTAIL.n48 VTAIL.n42 8.14595
R1209 VTAIL.n82 VTAIL.n76 8.14595
R1210 VTAIL.n218 VTAIL.n212 8.14595
R1211 VTAIL.n184 VTAIL.n178 8.14595
R1212 VTAIL.n150 VTAIL.n144 8.14595
R1213 VTAIL.n116 VTAIL.n110 8.14595
R1214 VTAIL.n251 VTAIL.n248 7.3702
R1215 VTAIL.n13 VTAIL.n10 7.3702
R1216 VTAIL.n47 VTAIL.n44 7.3702
R1217 VTAIL.n81 VTAIL.n78 7.3702
R1218 VTAIL.n217 VTAIL.n214 7.3702
R1219 VTAIL.n183 VTAIL.n180 7.3702
R1220 VTAIL.n149 VTAIL.n146 7.3702
R1221 VTAIL.n115 VTAIL.n112 7.3702
R1222 VTAIL.n252 VTAIL.n251 5.81868
R1223 VTAIL.n14 VTAIL.n13 5.81868
R1224 VTAIL.n48 VTAIL.n47 5.81868
R1225 VTAIL.n82 VTAIL.n81 5.81868
R1226 VTAIL.n218 VTAIL.n217 5.81868
R1227 VTAIL.n184 VTAIL.n183 5.81868
R1228 VTAIL.n150 VTAIL.n149 5.81868
R1229 VTAIL.n116 VTAIL.n115 5.81868
R1230 VTAIL.n255 VTAIL.n246 5.04292
R1231 VTAIL.n17 VTAIL.n8 5.04292
R1232 VTAIL.n51 VTAIL.n42 5.04292
R1233 VTAIL.n85 VTAIL.n76 5.04292
R1234 VTAIL.n221 VTAIL.n212 5.04292
R1235 VTAIL.n187 VTAIL.n178 5.04292
R1236 VTAIL.n153 VTAIL.n144 5.04292
R1237 VTAIL.n119 VTAIL.n110 5.04292
R1238 VTAIL.n256 VTAIL.n244 4.26717
R1239 VTAIL.n18 VTAIL.n6 4.26717
R1240 VTAIL.n52 VTAIL.n40 4.26717
R1241 VTAIL.n86 VTAIL.n74 4.26717
R1242 VTAIL.n222 VTAIL.n210 4.26717
R1243 VTAIL.n188 VTAIL.n176 4.26717
R1244 VTAIL.n154 VTAIL.n142 4.26717
R1245 VTAIL.n120 VTAIL.n108 4.26717
R1246 VTAIL.n260 VTAIL.n259 3.49141
R1247 VTAIL.n22 VTAIL.n21 3.49141
R1248 VTAIL.n56 VTAIL.n55 3.49141
R1249 VTAIL.n90 VTAIL.n89 3.49141
R1250 VTAIL.n226 VTAIL.n225 3.49141
R1251 VTAIL.n192 VTAIL.n191 3.49141
R1252 VTAIL.n158 VTAIL.n157 3.49141
R1253 VTAIL.n124 VTAIL.n123 3.49141
R1254 VTAIL.n169 VTAIL.n135 3.37119
R1255 VTAIL.n237 VTAIL.n203 3.37119
R1256 VTAIL.n101 VTAIL.n67 3.37119
R1257 VTAIL.n263 VTAIL.n242 2.71565
R1258 VTAIL.n25 VTAIL.n4 2.71565
R1259 VTAIL.n59 VTAIL.n38 2.71565
R1260 VTAIL.n93 VTAIL.n72 2.71565
R1261 VTAIL.n229 VTAIL.n208 2.71565
R1262 VTAIL.n195 VTAIL.n174 2.71565
R1263 VTAIL.n161 VTAIL.n140 2.71565
R1264 VTAIL.n127 VTAIL.n106 2.71565
R1265 VTAIL.n182 VTAIL.n181 2.41347
R1266 VTAIL.n148 VTAIL.n147 2.41347
R1267 VTAIL.n114 VTAIL.n113 2.41347
R1268 VTAIL.n250 VTAIL.n249 2.41347
R1269 VTAIL.n12 VTAIL.n11 2.41347
R1270 VTAIL.n46 VTAIL.n45 2.41347
R1271 VTAIL.n80 VTAIL.n79 2.41347
R1272 VTAIL.n216 VTAIL.n215 2.41347
R1273 VTAIL.n264 VTAIL.n240 1.93989
R1274 VTAIL.n26 VTAIL.n2 1.93989
R1275 VTAIL.n60 VTAIL.n36 1.93989
R1276 VTAIL.n94 VTAIL.n70 1.93989
R1277 VTAIL.n230 VTAIL.n206 1.93989
R1278 VTAIL.n196 VTAIL.n172 1.93989
R1279 VTAIL.n162 VTAIL.n138 1.93989
R1280 VTAIL.n128 VTAIL.n104 1.93989
R1281 VTAIL VTAIL.n33 1.74403
R1282 VTAIL VTAIL.n271 1.62766
R1283 VTAIL.n268 VTAIL.n267 1.16414
R1284 VTAIL.n30 VTAIL.n29 1.16414
R1285 VTAIL.n64 VTAIL.n63 1.16414
R1286 VTAIL.n98 VTAIL.n97 1.16414
R1287 VTAIL.n234 VTAIL.n233 1.16414
R1288 VTAIL.n200 VTAIL.n199 1.16414
R1289 VTAIL.n166 VTAIL.n165 1.16414
R1290 VTAIL.n132 VTAIL.n131 1.16414
R1291 VTAIL.n203 VTAIL.n169 0.470328
R1292 VTAIL.n67 VTAIL.n33 0.470328
R1293 VTAIL.n270 VTAIL.n238 0.388379
R1294 VTAIL.n32 VTAIL.n0 0.388379
R1295 VTAIL.n66 VTAIL.n34 0.388379
R1296 VTAIL.n100 VTAIL.n68 0.388379
R1297 VTAIL.n236 VTAIL.n204 0.388379
R1298 VTAIL.n202 VTAIL.n170 0.388379
R1299 VTAIL.n168 VTAIL.n136 0.388379
R1300 VTAIL.n134 VTAIL.n102 0.388379
R1301 VTAIL.n250 VTAIL.n245 0.155672
R1302 VTAIL.n257 VTAIL.n245 0.155672
R1303 VTAIL.n258 VTAIL.n257 0.155672
R1304 VTAIL.n258 VTAIL.n241 0.155672
R1305 VTAIL.n265 VTAIL.n241 0.155672
R1306 VTAIL.n266 VTAIL.n265 0.155672
R1307 VTAIL.n12 VTAIL.n7 0.155672
R1308 VTAIL.n19 VTAIL.n7 0.155672
R1309 VTAIL.n20 VTAIL.n19 0.155672
R1310 VTAIL.n20 VTAIL.n3 0.155672
R1311 VTAIL.n27 VTAIL.n3 0.155672
R1312 VTAIL.n28 VTAIL.n27 0.155672
R1313 VTAIL.n46 VTAIL.n41 0.155672
R1314 VTAIL.n53 VTAIL.n41 0.155672
R1315 VTAIL.n54 VTAIL.n53 0.155672
R1316 VTAIL.n54 VTAIL.n37 0.155672
R1317 VTAIL.n61 VTAIL.n37 0.155672
R1318 VTAIL.n62 VTAIL.n61 0.155672
R1319 VTAIL.n80 VTAIL.n75 0.155672
R1320 VTAIL.n87 VTAIL.n75 0.155672
R1321 VTAIL.n88 VTAIL.n87 0.155672
R1322 VTAIL.n88 VTAIL.n71 0.155672
R1323 VTAIL.n95 VTAIL.n71 0.155672
R1324 VTAIL.n96 VTAIL.n95 0.155672
R1325 VTAIL.n232 VTAIL.n231 0.155672
R1326 VTAIL.n231 VTAIL.n207 0.155672
R1327 VTAIL.n224 VTAIL.n207 0.155672
R1328 VTAIL.n224 VTAIL.n223 0.155672
R1329 VTAIL.n223 VTAIL.n211 0.155672
R1330 VTAIL.n216 VTAIL.n211 0.155672
R1331 VTAIL.n198 VTAIL.n197 0.155672
R1332 VTAIL.n197 VTAIL.n173 0.155672
R1333 VTAIL.n190 VTAIL.n173 0.155672
R1334 VTAIL.n190 VTAIL.n189 0.155672
R1335 VTAIL.n189 VTAIL.n177 0.155672
R1336 VTAIL.n182 VTAIL.n177 0.155672
R1337 VTAIL.n164 VTAIL.n163 0.155672
R1338 VTAIL.n163 VTAIL.n139 0.155672
R1339 VTAIL.n156 VTAIL.n139 0.155672
R1340 VTAIL.n156 VTAIL.n155 0.155672
R1341 VTAIL.n155 VTAIL.n143 0.155672
R1342 VTAIL.n148 VTAIL.n143 0.155672
R1343 VTAIL.n130 VTAIL.n129 0.155672
R1344 VTAIL.n129 VTAIL.n105 0.155672
R1345 VTAIL.n122 VTAIL.n105 0.155672
R1346 VTAIL.n122 VTAIL.n121 0.155672
R1347 VTAIL.n121 VTAIL.n109 0.155672
R1348 VTAIL.n114 VTAIL.n109 0.155672
R1349 VDD1 VDD1.n1 130.525
R1350 VDD1 VDD1.n0 90.6284
R1351 VDD1.n0 VDD1.t2 5.00127
R1352 VDD1.n0 VDD1.t0 5.00127
R1353 VDD1.n1 VDD1.t1 5.00127
R1354 VDD1.n1 VDD1.t3 5.00127
R1355 VN.n1 VN.t0 78.6291
R1356 VN.n0 VN.t1 78.6291
R1357 VN.n0 VN.t2 77.3889
R1358 VN.n1 VN.t3 77.3889
R1359 VN VN.n1 47.5092
R1360 VN VN.n0 2.11145
R1361 VDD2.n2 VDD2.n0 130
R1362 VDD2.n2 VDD2.n1 90.5702
R1363 VDD2.n1 VDD2.t0 5.00127
R1364 VDD2.n1 VDD2.t3 5.00127
R1365 VDD2.n0 VDD2.t2 5.00127
R1366 VDD2.n0 VDD2.t1 5.00127
R1367 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 2.8547f
C1 VP w_n3316_n2268# 6.11351f
C2 VP B 1.94747f
C3 VDD2 VTAIL 4.56227f
C4 VN VTAIL 3.31615f
C5 VDD1 VP 3.16049f
C6 VDD2 w_n3316_n2268# 1.5693f
C7 VDD2 B 1.35573f
C8 VN B 1.2314f
C9 VN w_n3316_n2268# 5.68474f
C10 B VTAIL 3.44787f
C11 w_n3316_n2268# VTAIL 2.80399f
C12 VDD1 VDD2 1.26243f
C13 VDD1 VN 0.150371f
C14 VDD1 VTAIL 4.50149f
C15 B w_n3316_n2268# 8.91758f
C16 VDD2 VP 0.45715f
C17 VN VP 5.8733f
C18 VP VTAIL 3.33026f
C19 VDD1 w_n3316_n2268# 1.49157f
C20 VDD1 B 1.28736f
C21 VDD2 VSUBS 0.984277f
C22 VDD1 VSUBS 5.66774f
C23 VTAIL VSUBS 0.796395f
C24 VN VSUBS 5.89809f
C25 VP VSUBS 2.44998f
C26 B VSUBS 4.655326f
C27 w_n3316_n2268# VSUBS 93.710205f
C28 VDD2.t2 VSUBS 0.146223f
C29 VDD2.t1 VSUBS 0.146223f
C30 VDD2.n0 VSUBS 1.51774f
C31 VDD2.t0 VSUBS 0.146223f
C32 VDD2.t3 VSUBS 0.146223f
C33 VDD2.n1 VSUBS 1.00985f
C34 VDD2.n2 VSUBS 4.0722f
C35 VN.t2 VSUBS 2.61718f
C36 VN.t1 VSUBS 2.63337f
C37 VN.n0 VSUBS 1.53358f
C38 VN.t0 VSUBS 2.63337f
C39 VN.t3 VSUBS 2.61718f
C40 VN.n1 VSUBS 3.54219f
C41 VDD1.t2 VSUBS 0.148047f
C42 VDD1.t0 VSUBS 0.148047f
C43 VDD1.n0 VSUBS 1.02295f
C44 VDD1.t1 VSUBS 0.148047f
C45 VDD1.t3 VSUBS 0.148047f
C46 VDD1.n1 VSUBS 1.55899f
C47 VTAIL.n0 VSUBS 0.015883f
C48 VTAIL.n1 VSUBS 0.035868f
C49 VTAIL.n2 VSUBS 0.016068f
C50 VTAIL.n3 VSUBS 0.02824f
C51 VTAIL.n4 VSUBS 0.015175f
C52 VTAIL.n5 VSUBS 0.035868f
C53 VTAIL.n6 VSUBS 0.016068f
C54 VTAIL.n7 VSUBS 0.02824f
C55 VTAIL.n8 VSUBS 0.015175f
C56 VTAIL.n9 VSUBS 0.026901f
C57 VTAIL.n10 VSUBS 0.026978f
C58 VTAIL.t2 VSUBS 0.077089f
C59 VTAIL.n11 VSUBS 0.152438f
C60 VTAIL.n12 VSUBS 0.706389f
C61 VTAIL.n13 VSUBS 0.015175f
C62 VTAIL.n14 VSUBS 0.016068f
C63 VTAIL.n15 VSUBS 0.035868f
C64 VTAIL.n16 VSUBS 0.035868f
C65 VTAIL.n17 VSUBS 0.016068f
C66 VTAIL.n18 VSUBS 0.015175f
C67 VTAIL.n19 VSUBS 0.02824f
C68 VTAIL.n20 VSUBS 0.02824f
C69 VTAIL.n21 VSUBS 0.015175f
C70 VTAIL.n22 VSUBS 0.016068f
C71 VTAIL.n23 VSUBS 0.035868f
C72 VTAIL.n24 VSUBS 0.035868f
C73 VTAIL.n25 VSUBS 0.016068f
C74 VTAIL.n26 VSUBS 0.015175f
C75 VTAIL.n27 VSUBS 0.02824f
C76 VTAIL.n28 VSUBS 0.070676f
C77 VTAIL.n29 VSUBS 0.015175f
C78 VTAIL.n30 VSUBS 0.016068f
C79 VTAIL.n31 VSUBS 0.079091f
C80 VTAIL.n32 VSUBS 0.052009f
C81 VTAIL.n33 VSUBS 0.228143f
C82 VTAIL.n34 VSUBS 0.015883f
C83 VTAIL.n35 VSUBS 0.035868f
C84 VTAIL.n36 VSUBS 0.016068f
C85 VTAIL.n37 VSUBS 0.02824f
C86 VTAIL.n38 VSUBS 0.015175f
C87 VTAIL.n39 VSUBS 0.035868f
C88 VTAIL.n40 VSUBS 0.016068f
C89 VTAIL.n41 VSUBS 0.02824f
C90 VTAIL.n42 VSUBS 0.015175f
C91 VTAIL.n43 VSUBS 0.026901f
C92 VTAIL.n44 VSUBS 0.026978f
C93 VTAIL.t4 VSUBS 0.077089f
C94 VTAIL.n45 VSUBS 0.152438f
C95 VTAIL.n46 VSUBS 0.706389f
C96 VTAIL.n47 VSUBS 0.015175f
C97 VTAIL.n48 VSUBS 0.016068f
C98 VTAIL.n49 VSUBS 0.035868f
C99 VTAIL.n50 VSUBS 0.035868f
C100 VTAIL.n51 VSUBS 0.016068f
C101 VTAIL.n52 VSUBS 0.015175f
C102 VTAIL.n53 VSUBS 0.02824f
C103 VTAIL.n54 VSUBS 0.02824f
C104 VTAIL.n55 VSUBS 0.015175f
C105 VTAIL.n56 VSUBS 0.016068f
C106 VTAIL.n57 VSUBS 0.035868f
C107 VTAIL.n58 VSUBS 0.035868f
C108 VTAIL.n59 VSUBS 0.016068f
C109 VTAIL.n60 VSUBS 0.015175f
C110 VTAIL.n61 VSUBS 0.02824f
C111 VTAIL.n62 VSUBS 0.070676f
C112 VTAIL.n63 VSUBS 0.015175f
C113 VTAIL.n64 VSUBS 0.016068f
C114 VTAIL.n65 VSUBS 0.079091f
C115 VTAIL.n66 VSUBS 0.052009f
C116 VTAIL.n67 VSUBS 0.376207f
C117 VTAIL.n68 VSUBS 0.015883f
C118 VTAIL.n69 VSUBS 0.035868f
C119 VTAIL.n70 VSUBS 0.016068f
C120 VTAIL.n71 VSUBS 0.02824f
C121 VTAIL.n72 VSUBS 0.015175f
C122 VTAIL.n73 VSUBS 0.035868f
C123 VTAIL.n74 VSUBS 0.016068f
C124 VTAIL.n75 VSUBS 0.02824f
C125 VTAIL.n76 VSUBS 0.015175f
C126 VTAIL.n77 VSUBS 0.026901f
C127 VTAIL.n78 VSUBS 0.026978f
C128 VTAIL.t6 VSUBS 0.077089f
C129 VTAIL.n79 VSUBS 0.152438f
C130 VTAIL.n80 VSUBS 0.706389f
C131 VTAIL.n81 VSUBS 0.015175f
C132 VTAIL.n82 VSUBS 0.016068f
C133 VTAIL.n83 VSUBS 0.035868f
C134 VTAIL.n84 VSUBS 0.035868f
C135 VTAIL.n85 VSUBS 0.016068f
C136 VTAIL.n86 VSUBS 0.015175f
C137 VTAIL.n87 VSUBS 0.02824f
C138 VTAIL.n88 VSUBS 0.02824f
C139 VTAIL.n89 VSUBS 0.015175f
C140 VTAIL.n90 VSUBS 0.016068f
C141 VTAIL.n91 VSUBS 0.035868f
C142 VTAIL.n92 VSUBS 0.035868f
C143 VTAIL.n93 VSUBS 0.016068f
C144 VTAIL.n94 VSUBS 0.015175f
C145 VTAIL.n95 VSUBS 0.02824f
C146 VTAIL.n96 VSUBS 0.070676f
C147 VTAIL.n97 VSUBS 0.015175f
C148 VTAIL.n98 VSUBS 0.016068f
C149 VTAIL.n99 VSUBS 0.079091f
C150 VTAIL.n100 VSUBS 0.052009f
C151 VTAIL.n101 VSUBS 1.53367f
C152 VTAIL.n102 VSUBS 0.015883f
C153 VTAIL.n103 VSUBS 0.035868f
C154 VTAIL.n104 VSUBS 0.016068f
C155 VTAIL.n105 VSUBS 0.02824f
C156 VTAIL.n106 VSUBS 0.015175f
C157 VTAIL.n107 VSUBS 0.035868f
C158 VTAIL.n108 VSUBS 0.016068f
C159 VTAIL.n109 VSUBS 0.02824f
C160 VTAIL.n110 VSUBS 0.015175f
C161 VTAIL.n111 VSUBS 0.026901f
C162 VTAIL.n112 VSUBS 0.026978f
C163 VTAIL.t0 VSUBS 0.077089f
C164 VTAIL.n113 VSUBS 0.152438f
C165 VTAIL.n114 VSUBS 0.706389f
C166 VTAIL.n115 VSUBS 0.015175f
C167 VTAIL.n116 VSUBS 0.016068f
C168 VTAIL.n117 VSUBS 0.035868f
C169 VTAIL.n118 VSUBS 0.035868f
C170 VTAIL.n119 VSUBS 0.016068f
C171 VTAIL.n120 VSUBS 0.015175f
C172 VTAIL.n121 VSUBS 0.02824f
C173 VTAIL.n122 VSUBS 0.02824f
C174 VTAIL.n123 VSUBS 0.015175f
C175 VTAIL.n124 VSUBS 0.016068f
C176 VTAIL.n125 VSUBS 0.035868f
C177 VTAIL.n126 VSUBS 0.035868f
C178 VTAIL.n127 VSUBS 0.016068f
C179 VTAIL.n128 VSUBS 0.015175f
C180 VTAIL.n129 VSUBS 0.02824f
C181 VTAIL.n130 VSUBS 0.070676f
C182 VTAIL.n131 VSUBS 0.015175f
C183 VTAIL.n132 VSUBS 0.016068f
C184 VTAIL.n133 VSUBS 0.079091f
C185 VTAIL.n134 VSUBS 0.052009f
C186 VTAIL.n135 VSUBS 1.53367f
C187 VTAIL.n136 VSUBS 0.015883f
C188 VTAIL.n137 VSUBS 0.035868f
C189 VTAIL.n138 VSUBS 0.016068f
C190 VTAIL.n139 VSUBS 0.02824f
C191 VTAIL.n140 VSUBS 0.015175f
C192 VTAIL.n141 VSUBS 0.035868f
C193 VTAIL.n142 VSUBS 0.016068f
C194 VTAIL.n143 VSUBS 0.02824f
C195 VTAIL.n144 VSUBS 0.015175f
C196 VTAIL.n145 VSUBS 0.026901f
C197 VTAIL.n146 VSUBS 0.026978f
C198 VTAIL.t1 VSUBS 0.077089f
C199 VTAIL.n147 VSUBS 0.152438f
C200 VTAIL.n148 VSUBS 0.706389f
C201 VTAIL.n149 VSUBS 0.015175f
C202 VTAIL.n150 VSUBS 0.016068f
C203 VTAIL.n151 VSUBS 0.035868f
C204 VTAIL.n152 VSUBS 0.035868f
C205 VTAIL.n153 VSUBS 0.016068f
C206 VTAIL.n154 VSUBS 0.015175f
C207 VTAIL.n155 VSUBS 0.02824f
C208 VTAIL.n156 VSUBS 0.02824f
C209 VTAIL.n157 VSUBS 0.015175f
C210 VTAIL.n158 VSUBS 0.016068f
C211 VTAIL.n159 VSUBS 0.035868f
C212 VTAIL.n160 VSUBS 0.035868f
C213 VTAIL.n161 VSUBS 0.016068f
C214 VTAIL.n162 VSUBS 0.015175f
C215 VTAIL.n163 VSUBS 0.02824f
C216 VTAIL.n164 VSUBS 0.070676f
C217 VTAIL.n165 VSUBS 0.015175f
C218 VTAIL.n166 VSUBS 0.016068f
C219 VTAIL.n167 VSUBS 0.079091f
C220 VTAIL.n168 VSUBS 0.052009f
C221 VTAIL.n169 VSUBS 0.376207f
C222 VTAIL.n170 VSUBS 0.015883f
C223 VTAIL.n171 VSUBS 0.035868f
C224 VTAIL.n172 VSUBS 0.016068f
C225 VTAIL.n173 VSUBS 0.02824f
C226 VTAIL.n174 VSUBS 0.015175f
C227 VTAIL.n175 VSUBS 0.035868f
C228 VTAIL.n176 VSUBS 0.016068f
C229 VTAIL.n177 VSUBS 0.02824f
C230 VTAIL.n178 VSUBS 0.015175f
C231 VTAIL.n179 VSUBS 0.026901f
C232 VTAIL.n180 VSUBS 0.026978f
C233 VTAIL.t5 VSUBS 0.077089f
C234 VTAIL.n181 VSUBS 0.152438f
C235 VTAIL.n182 VSUBS 0.706389f
C236 VTAIL.n183 VSUBS 0.015175f
C237 VTAIL.n184 VSUBS 0.016068f
C238 VTAIL.n185 VSUBS 0.035868f
C239 VTAIL.n186 VSUBS 0.035868f
C240 VTAIL.n187 VSUBS 0.016068f
C241 VTAIL.n188 VSUBS 0.015175f
C242 VTAIL.n189 VSUBS 0.02824f
C243 VTAIL.n190 VSUBS 0.02824f
C244 VTAIL.n191 VSUBS 0.015175f
C245 VTAIL.n192 VSUBS 0.016068f
C246 VTAIL.n193 VSUBS 0.035868f
C247 VTAIL.n194 VSUBS 0.035868f
C248 VTAIL.n195 VSUBS 0.016068f
C249 VTAIL.n196 VSUBS 0.015175f
C250 VTAIL.n197 VSUBS 0.02824f
C251 VTAIL.n198 VSUBS 0.070676f
C252 VTAIL.n199 VSUBS 0.015175f
C253 VTAIL.n200 VSUBS 0.016068f
C254 VTAIL.n201 VSUBS 0.079091f
C255 VTAIL.n202 VSUBS 0.052009f
C256 VTAIL.n203 VSUBS 0.376207f
C257 VTAIL.n204 VSUBS 0.015883f
C258 VTAIL.n205 VSUBS 0.035868f
C259 VTAIL.n206 VSUBS 0.016068f
C260 VTAIL.n207 VSUBS 0.02824f
C261 VTAIL.n208 VSUBS 0.015175f
C262 VTAIL.n209 VSUBS 0.035868f
C263 VTAIL.n210 VSUBS 0.016068f
C264 VTAIL.n211 VSUBS 0.02824f
C265 VTAIL.n212 VSUBS 0.015175f
C266 VTAIL.n213 VSUBS 0.026901f
C267 VTAIL.n214 VSUBS 0.026978f
C268 VTAIL.t7 VSUBS 0.077089f
C269 VTAIL.n215 VSUBS 0.152438f
C270 VTAIL.n216 VSUBS 0.706389f
C271 VTAIL.n217 VSUBS 0.015175f
C272 VTAIL.n218 VSUBS 0.016068f
C273 VTAIL.n219 VSUBS 0.035868f
C274 VTAIL.n220 VSUBS 0.035868f
C275 VTAIL.n221 VSUBS 0.016068f
C276 VTAIL.n222 VSUBS 0.015175f
C277 VTAIL.n223 VSUBS 0.02824f
C278 VTAIL.n224 VSUBS 0.02824f
C279 VTAIL.n225 VSUBS 0.015175f
C280 VTAIL.n226 VSUBS 0.016068f
C281 VTAIL.n227 VSUBS 0.035868f
C282 VTAIL.n228 VSUBS 0.035868f
C283 VTAIL.n229 VSUBS 0.016068f
C284 VTAIL.n230 VSUBS 0.015175f
C285 VTAIL.n231 VSUBS 0.02824f
C286 VTAIL.n232 VSUBS 0.070676f
C287 VTAIL.n233 VSUBS 0.015175f
C288 VTAIL.n234 VSUBS 0.016068f
C289 VTAIL.n235 VSUBS 0.079091f
C290 VTAIL.n236 VSUBS 0.052009f
C291 VTAIL.n237 VSUBS 1.53367f
C292 VTAIL.n238 VSUBS 0.015883f
C293 VTAIL.n239 VSUBS 0.035868f
C294 VTAIL.n240 VSUBS 0.016068f
C295 VTAIL.n241 VSUBS 0.02824f
C296 VTAIL.n242 VSUBS 0.015175f
C297 VTAIL.n243 VSUBS 0.035868f
C298 VTAIL.n244 VSUBS 0.016068f
C299 VTAIL.n245 VSUBS 0.02824f
C300 VTAIL.n246 VSUBS 0.015175f
C301 VTAIL.n247 VSUBS 0.026901f
C302 VTAIL.n248 VSUBS 0.026978f
C303 VTAIL.t3 VSUBS 0.077089f
C304 VTAIL.n249 VSUBS 0.152438f
C305 VTAIL.n250 VSUBS 0.706389f
C306 VTAIL.n251 VSUBS 0.015175f
C307 VTAIL.n252 VSUBS 0.016068f
C308 VTAIL.n253 VSUBS 0.035868f
C309 VTAIL.n254 VSUBS 0.035868f
C310 VTAIL.n255 VSUBS 0.016068f
C311 VTAIL.n256 VSUBS 0.015175f
C312 VTAIL.n257 VSUBS 0.02824f
C313 VTAIL.n258 VSUBS 0.02824f
C314 VTAIL.n259 VSUBS 0.015175f
C315 VTAIL.n260 VSUBS 0.016068f
C316 VTAIL.n261 VSUBS 0.035868f
C317 VTAIL.n262 VSUBS 0.035868f
C318 VTAIL.n263 VSUBS 0.016068f
C319 VTAIL.n264 VSUBS 0.015175f
C320 VTAIL.n265 VSUBS 0.02824f
C321 VTAIL.n266 VSUBS 0.070676f
C322 VTAIL.n267 VSUBS 0.015175f
C323 VTAIL.n268 VSUBS 0.016068f
C324 VTAIL.n269 VSUBS 0.079091f
C325 VTAIL.n270 VSUBS 0.052009f
C326 VTAIL.n271 VSUBS 1.37502f
C327 VP.t0 VSUBS 2.2516f
C328 VP.n0 VSUBS 0.966905f
C329 VP.n1 VSUBS 0.036393f
C330 VP.n2 VSUBS 0.052903f
C331 VP.n3 VSUBS 0.036393f
C332 VP.n4 VSUBS 0.04783f
C333 VP.t1 VSUBS 2.74449f
C334 VP.t3 VSUBS 2.72763f
C335 VP.n5 VSUBS 3.67658f
C336 VP.t2 VSUBS 2.2516f
C337 VP.n6 VSUBS 0.966905f
C338 VP.n7 VSUBS 1.93025f
C339 VP.n8 VSUBS 0.058728f
C340 VP.n9 VSUBS 0.036393f
C341 VP.n10 VSUBS 0.067487f
C342 VP.n11 VSUBS 0.067487f
C343 VP.n12 VSUBS 0.052903f
C344 VP.n13 VSUBS 0.036393f
C345 VP.n14 VSUBS 0.036393f
C346 VP.n15 VSUBS 0.036393f
C347 VP.n16 VSUBS 0.067487f
C348 VP.n17 VSUBS 0.067487f
C349 VP.n18 VSUBS 0.04783f
C350 VP.n19 VSUBS 0.058728f
C351 VP.n20 VSUBS 0.098965f
C352 B.n0 VSUBS 0.006753f
C353 B.n1 VSUBS 0.006753f
C354 B.n2 VSUBS 0.009988f
C355 B.n3 VSUBS 0.007654f
C356 B.n4 VSUBS 0.007654f
C357 B.n5 VSUBS 0.007654f
C358 B.n6 VSUBS 0.007654f
C359 B.n7 VSUBS 0.007654f
C360 B.n8 VSUBS 0.007654f
C361 B.n9 VSUBS 0.007654f
C362 B.n10 VSUBS 0.007654f
C363 B.n11 VSUBS 0.007654f
C364 B.n12 VSUBS 0.007654f
C365 B.n13 VSUBS 0.007654f
C366 B.n14 VSUBS 0.007654f
C367 B.n15 VSUBS 0.007654f
C368 B.n16 VSUBS 0.007654f
C369 B.n17 VSUBS 0.007654f
C370 B.n18 VSUBS 0.007654f
C371 B.n19 VSUBS 0.007654f
C372 B.n20 VSUBS 0.007654f
C373 B.n21 VSUBS 0.007654f
C374 B.n22 VSUBS 0.007654f
C375 B.n23 VSUBS 0.019444f
C376 B.n24 VSUBS 0.007654f
C377 B.n25 VSUBS 0.007654f
C378 B.n26 VSUBS 0.007654f
C379 B.n27 VSUBS 0.007654f
C380 B.n28 VSUBS 0.007654f
C381 B.n29 VSUBS 0.007654f
C382 B.n30 VSUBS 0.007654f
C383 B.n31 VSUBS 0.007654f
C384 B.n32 VSUBS 0.007654f
C385 B.n33 VSUBS 0.007654f
C386 B.n34 VSUBS 0.007654f
C387 B.n35 VSUBS 0.007654f
C388 B.t10 VSUBS 0.107177f
C389 B.t11 VSUBS 0.144822f
C390 B.t9 VSUBS 1.21667f
C391 B.n36 VSUBS 0.23972f
C392 B.n37 VSUBS 0.185922f
C393 B.n38 VSUBS 0.007654f
C394 B.n39 VSUBS 0.007654f
C395 B.n40 VSUBS 0.007654f
C396 B.n41 VSUBS 0.007654f
C397 B.n42 VSUBS 0.004277f
C398 B.n43 VSUBS 0.007654f
C399 B.t7 VSUBS 0.107179f
C400 B.t8 VSUBS 0.144823f
C401 B.t6 VSUBS 1.21667f
C402 B.n44 VSUBS 0.239718f
C403 B.n45 VSUBS 0.18592f
C404 B.n46 VSUBS 0.017733f
C405 B.n47 VSUBS 0.007654f
C406 B.n48 VSUBS 0.007654f
C407 B.n49 VSUBS 0.007654f
C408 B.n50 VSUBS 0.007654f
C409 B.n51 VSUBS 0.007654f
C410 B.n52 VSUBS 0.007654f
C411 B.n53 VSUBS 0.007654f
C412 B.n54 VSUBS 0.007654f
C413 B.n55 VSUBS 0.007654f
C414 B.n56 VSUBS 0.007654f
C415 B.n57 VSUBS 0.007654f
C416 B.n58 VSUBS 0.018824f
C417 B.n59 VSUBS 0.007654f
C418 B.n60 VSUBS 0.007654f
C419 B.n61 VSUBS 0.007654f
C420 B.n62 VSUBS 0.007654f
C421 B.n63 VSUBS 0.007654f
C422 B.n64 VSUBS 0.007654f
C423 B.n65 VSUBS 0.007654f
C424 B.n66 VSUBS 0.007654f
C425 B.n67 VSUBS 0.007654f
C426 B.n68 VSUBS 0.007654f
C427 B.n69 VSUBS 0.007654f
C428 B.n70 VSUBS 0.007654f
C429 B.n71 VSUBS 0.007654f
C430 B.n72 VSUBS 0.007654f
C431 B.n73 VSUBS 0.007654f
C432 B.n74 VSUBS 0.007654f
C433 B.n75 VSUBS 0.007654f
C434 B.n76 VSUBS 0.007654f
C435 B.n77 VSUBS 0.007654f
C436 B.n78 VSUBS 0.007654f
C437 B.n79 VSUBS 0.007654f
C438 B.n80 VSUBS 0.007654f
C439 B.n81 VSUBS 0.007654f
C440 B.n82 VSUBS 0.007654f
C441 B.n83 VSUBS 0.007654f
C442 B.n84 VSUBS 0.007654f
C443 B.n85 VSUBS 0.007654f
C444 B.n86 VSUBS 0.007654f
C445 B.n87 VSUBS 0.007654f
C446 B.n88 VSUBS 0.007654f
C447 B.n89 VSUBS 0.007654f
C448 B.n90 VSUBS 0.007654f
C449 B.n91 VSUBS 0.007654f
C450 B.n92 VSUBS 0.007654f
C451 B.n93 VSUBS 0.007654f
C452 B.n94 VSUBS 0.007654f
C453 B.n95 VSUBS 0.007654f
C454 B.n96 VSUBS 0.007654f
C455 B.n97 VSUBS 0.007654f
C456 B.n98 VSUBS 0.007654f
C457 B.n99 VSUBS 0.007654f
C458 B.n100 VSUBS 0.007654f
C459 B.n101 VSUBS 0.018625f
C460 B.n102 VSUBS 0.007654f
C461 B.n103 VSUBS 0.007654f
C462 B.n104 VSUBS 0.007654f
C463 B.n105 VSUBS 0.007654f
C464 B.n106 VSUBS 0.007654f
C465 B.n107 VSUBS 0.007654f
C466 B.n108 VSUBS 0.007654f
C467 B.n109 VSUBS 0.007654f
C468 B.n110 VSUBS 0.007654f
C469 B.n111 VSUBS 0.007654f
C470 B.n112 VSUBS 0.007654f
C471 B.n113 VSUBS 0.007203f
C472 B.n114 VSUBS 0.007654f
C473 B.n115 VSUBS 0.007654f
C474 B.n116 VSUBS 0.007654f
C475 B.n117 VSUBS 0.007654f
C476 B.n118 VSUBS 0.007654f
C477 B.t5 VSUBS 0.107177f
C478 B.t4 VSUBS 0.144822f
C479 B.t3 VSUBS 1.21667f
C480 B.n119 VSUBS 0.23972f
C481 B.n120 VSUBS 0.185922f
C482 B.n121 VSUBS 0.007654f
C483 B.n122 VSUBS 0.007654f
C484 B.n123 VSUBS 0.007654f
C485 B.n124 VSUBS 0.007654f
C486 B.n125 VSUBS 0.007654f
C487 B.n126 VSUBS 0.007654f
C488 B.n127 VSUBS 0.007654f
C489 B.n128 VSUBS 0.007654f
C490 B.n129 VSUBS 0.007654f
C491 B.n130 VSUBS 0.007654f
C492 B.n131 VSUBS 0.007654f
C493 B.n132 VSUBS 0.007654f
C494 B.n133 VSUBS 0.018824f
C495 B.n134 VSUBS 0.007654f
C496 B.n135 VSUBS 0.007654f
C497 B.n136 VSUBS 0.007654f
C498 B.n137 VSUBS 0.007654f
C499 B.n138 VSUBS 0.007654f
C500 B.n139 VSUBS 0.007654f
C501 B.n140 VSUBS 0.007654f
C502 B.n141 VSUBS 0.007654f
C503 B.n142 VSUBS 0.007654f
C504 B.n143 VSUBS 0.007654f
C505 B.n144 VSUBS 0.007654f
C506 B.n145 VSUBS 0.007654f
C507 B.n146 VSUBS 0.007654f
C508 B.n147 VSUBS 0.007654f
C509 B.n148 VSUBS 0.007654f
C510 B.n149 VSUBS 0.007654f
C511 B.n150 VSUBS 0.007654f
C512 B.n151 VSUBS 0.007654f
C513 B.n152 VSUBS 0.007654f
C514 B.n153 VSUBS 0.007654f
C515 B.n154 VSUBS 0.007654f
C516 B.n155 VSUBS 0.007654f
C517 B.n156 VSUBS 0.007654f
C518 B.n157 VSUBS 0.007654f
C519 B.n158 VSUBS 0.007654f
C520 B.n159 VSUBS 0.007654f
C521 B.n160 VSUBS 0.007654f
C522 B.n161 VSUBS 0.007654f
C523 B.n162 VSUBS 0.007654f
C524 B.n163 VSUBS 0.007654f
C525 B.n164 VSUBS 0.007654f
C526 B.n165 VSUBS 0.007654f
C527 B.n166 VSUBS 0.007654f
C528 B.n167 VSUBS 0.007654f
C529 B.n168 VSUBS 0.007654f
C530 B.n169 VSUBS 0.007654f
C531 B.n170 VSUBS 0.007654f
C532 B.n171 VSUBS 0.007654f
C533 B.n172 VSUBS 0.007654f
C534 B.n173 VSUBS 0.007654f
C535 B.n174 VSUBS 0.007654f
C536 B.n175 VSUBS 0.007654f
C537 B.n176 VSUBS 0.007654f
C538 B.n177 VSUBS 0.007654f
C539 B.n178 VSUBS 0.007654f
C540 B.n179 VSUBS 0.007654f
C541 B.n180 VSUBS 0.007654f
C542 B.n181 VSUBS 0.007654f
C543 B.n182 VSUBS 0.007654f
C544 B.n183 VSUBS 0.007654f
C545 B.n184 VSUBS 0.007654f
C546 B.n185 VSUBS 0.007654f
C547 B.n186 VSUBS 0.007654f
C548 B.n187 VSUBS 0.007654f
C549 B.n188 VSUBS 0.007654f
C550 B.n189 VSUBS 0.007654f
C551 B.n190 VSUBS 0.007654f
C552 B.n191 VSUBS 0.007654f
C553 B.n192 VSUBS 0.007654f
C554 B.n193 VSUBS 0.007654f
C555 B.n194 VSUBS 0.007654f
C556 B.n195 VSUBS 0.007654f
C557 B.n196 VSUBS 0.007654f
C558 B.n197 VSUBS 0.007654f
C559 B.n198 VSUBS 0.007654f
C560 B.n199 VSUBS 0.007654f
C561 B.n200 VSUBS 0.007654f
C562 B.n201 VSUBS 0.007654f
C563 B.n202 VSUBS 0.007654f
C564 B.n203 VSUBS 0.007654f
C565 B.n204 VSUBS 0.007654f
C566 B.n205 VSUBS 0.007654f
C567 B.n206 VSUBS 0.007654f
C568 B.n207 VSUBS 0.007654f
C569 B.n208 VSUBS 0.007654f
C570 B.n209 VSUBS 0.007654f
C571 B.n210 VSUBS 0.007654f
C572 B.n211 VSUBS 0.007654f
C573 B.n212 VSUBS 0.007654f
C574 B.n213 VSUBS 0.007654f
C575 B.n214 VSUBS 0.018824f
C576 B.n215 VSUBS 0.019444f
C577 B.n216 VSUBS 0.019444f
C578 B.n217 VSUBS 0.007654f
C579 B.n218 VSUBS 0.007654f
C580 B.n219 VSUBS 0.007654f
C581 B.n220 VSUBS 0.007654f
C582 B.n221 VSUBS 0.007654f
C583 B.n222 VSUBS 0.007654f
C584 B.n223 VSUBS 0.007654f
C585 B.n224 VSUBS 0.007654f
C586 B.n225 VSUBS 0.007654f
C587 B.n226 VSUBS 0.007654f
C588 B.n227 VSUBS 0.007654f
C589 B.n228 VSUBS 0.007654f
C590 B.n229 VSUBS 0.007654f
C591 B.n230 VSUBS 0.007654f
C592 B.n231 VSUBS 0.007654f
C593 B.n232 VSUBS 0.007654f
C594 B.n233 VSUBS 0.007654f
C595 B.n234 VSUBS 0.007654f
C596 B.n235 VSUBS 0.007654f
C597 B.n236 VSUBS 0.007654f
C598 B.n237 VSUBS 0.007654f
C599 B.n238 VSUBS 0.007654f
C600 B.n239 VSUBS 0.007654f
C601 B.n240 VSUBS 0.007654f
C602 B.n241 VSUBS 0.007654f
C603 B.n242 VSUBS 0.007654f
C604 B.n243 VSUBS 0.007654f
C605 B.n244 VSUBS 0.007654f
C606 B.n245 VSUBS 0.007654f
C607 B.n246 VSUBS 0.007654f
C608 B.n247 VSUBS 0.007654f
C609 B.n248 VSUBS 0.007654f
C610 B.n249 VSUBS 0.007654f
C611 B.n250 VSUBS 0.007654f
C612 B.n251 VSUBS 0.007654f
C613 B.n252 VSUBS 0.007203f
C614 B.n253 VSUBS 0.017733f
C615 B.n254 VSUBS 0.004277f
C616 B.n255 VSUBS 0.007654f
C617 B.n256 VSUBS 0.007654f
C618 B.n257 VSUBS 0.007654f
C619 B.n258 VSUBS 0.007654f
C620 B.n259 VSUBS 0.007654f
C621 B.n260 VSUBS 0.007654f
C622 B.n261 VSUBS 0.007654f
C623 B.n262 VSUBS 0.007654f
C624 B.n263 VSUBS 0.007654f
C625 B.n264 VSUBS 0.007654f
C626 B.n265 VSUBS 0.007654f
C627 B.n266 VSUBS 0.007654f
C628 B.t2 VSUBS 0.107179f
C629 B.t1 VSUBS 0.144823f
C630 B.t0 VSUBS 1.21667f
C631 B.n267 VSUBS 0.239718f
C632 B.n268 VSUBS 0.18592f
C633 B.n269 VSUBS 0.017733f
C634 B.n270 VSUBS 0.004277f
C635 B.n271 VSUBS 0.007654f
C636 B.n272 VSUBS 0.007654f
C637 B.n273 VSUBS 0.007654f
C638 B.n274 VSUBS 0.007654f
C639 B.n275 VSUBS 0.007654f
C640 B.n276 VSUBS 0.007654f
C641 B.n277 VSUBS 0.007654f
C642 B.n278 VSUBS 0.007654f
C643 B.n279 VSUBS 0.007654f
C644 B.n280 VSUBS 0.007654f
C645 B.n281 VSUBS 0.007654f
C646 B.n282 VSUBS 0.007654f
C647 B.n283 VSUBS 0.007654f
C648 B.n284 VSUBS 0.007654f
C649 B.n285 VSUBS 0.007654f
C650 B.n286 VSUBS 0.007654f
C651 B.n287 VSUBS 0.007654f
C652 B.n288 VSUBS 0.007654f
C653 B.n289 VSUBS 0.007654f
C654 B.n290 VSUBS 0.007654f
C655 B.n291 VSUBS 0.007654f
C656 B.n292 VSUBS 0.007654f
C657 B.n293 VSUBS 0.007654f
C658 B.n294 VSUBS 0.007654f
C659 B.n295 VSUBS 0.007654f
C660 B.n296 VSUBS 0.007654f
C661 B.n297 VSUBS 0.007654f
C662 B.n298 VSUBS 0.007654f
C663 B.n299 VSUBS 0.007654f
C664 B.n300 VSUBS 0.007654f
C665 B.n301 VSUBS 0.007654f
C666 B.n302 VSUBS 0.007654f
C667 B.n303 VSUBS 0.007654f
C668 B.n304 VSUBS 0.007654f
C669 B.n305 VSUBS 0.007654f
C670 B.n306 VSUBS 0.007654f
C671 B.n307 VSUBS 0.007654f
C672 B.n308 VSUBS 0.019444f
C673 B.n309 VSUBS 0.018824f
C674 B.n310 VSUBS 0.019644f
C675 B.n311 VSUBS 0.007654f
C676 B.n312 VSUBS 0.007654f
C677 B.n313 VSUBS 0.007654f
C678 B.n314 VSUBS 0.007654f
C679 B.n315 VSUBS 0.007654f
C680 B.n316 VSUBS 0.007654f
C681 B.n317 VSUBS 0.007654f
C682 B.n318 VSUBS 0.007654f
C683 B.n319 VSUBS 0.007654f
C684 B.n320 VSUBS 0.007654f
C685 B.n321 VSUBS 0.007654f
C686 B.n322 VSUBS 0.007654f
C687 B.n323 VSUBS 0.007654f
C688 B.n324 VSUBS 0.007654f
C689 B.n325 VSUBS 0.007654f
C690 B.n326 VSUBS 0.007654f
C691 B.n327 VSUBS 0.007654f
C692 B.n328 VSUBS 0.007654f
C693 B.n329 VSUBS 0.007654f
C694 B.n330 VSUBS 0.007654f
C695 B.n331 VSUBS 0.007654f
C696 B.n332 VSUBS 0.007654f
C697 B.n333 VSUBS 0.007654f
C698 B.n334 VSUBS 0.007654f
C699 B.n335 VSUBS 0.007654f
C700 B.n336 VSUBS 0.007654f
C701 B.n337 VSUBS 0.007654f
C702 B.n338 VSUBS 0.007654f
C703 B.n339 VSUBS 0.007654f
C704 B.n340 VSUBS 0.007654f
C705 B.n341 VSUBS 0.007654f
C706 B.n342 VSUBS 0.007654f
C707 B.n343 VSUBS 0.007654f
C708 B.n344 VSUBS 0.007654f
C709 B.n345 VSUBS 0.007654f
C710 B.n346 VSUBS 0.007654f
C711 B.n347 VSUBS 0.007654f
C712 B.n348 VSUBS 0.007654f
C713 B.n349 VSUBS 0.007654f
C714 B.n350 VSUBS 0.007654f
C715 B.n351 VSUBS 0.007654f
C716 B.n352 VSUBS 0.007654f
C717 B.n353 VSUBS 0.007654f
C718 B.n354 VSUBS 0.007654f
C719 B.n355 VSUBS 0.007654f
C720 B.n356 VSUBS 0.007654f
C721 B.n357 VSUBS 0.007654f
C722 B.n358 VSUBS 0.007654f
C723 B.n359 VSUBS 0.007654f
C724 B.n360 VSUBS 0.007654f
C725 B.n361 VSUBS 0.007654f
C726 B.n362 VSUBS 0.007654f
C727 B.n363 VSUBS 0.007654f
C728 B.n364 VSUBS 0.007654f
C729 B.n365 VSUBS 0.007654f
C730 B.n366 VSUBS 0.007654f
C731 B.n367 VSUBS 0.007654f
C732 B.n368 VSUBS 0.007654f
C733 B.n369 VSUBS 0.007654f
C734 B.n370 VSUBS 0.007654f
C735 B.n371 VSUBS 0.007654f
C736 B.n372 VSUBS 0.007654f
C737 B.n373 VSUBS 0.007654f
C738 B.n374 VSUBS 0.007654f
C739 B.n375 VSUBS 0.007654f
C740 B.n376 VSUBS 0.007654f
C741 B.n377 VSUBS 0.007654f
C742 B.n378 VSUBS 0.007654f
C743 B.n379 VSUBS 0.007654f
C744 B.n380 VSUBS 0.007654f
C745 B.n381 VSUBS 0.007654f
C746 B.n382 VSUBS 0.007654f
C747 B.n383 VSUBS 0.007654f
C748 B.n384 VSUBS 0.007654f
C749 B.n385 VSUBS 0.007654f
C750 B.n386 VSUBS 0.007654f
C751 B.n387 VSUBS 0.007654f
C752 B.n388 VSUBS 0.007654f
C753 B.n389 VSUBS 0.007654f
C754 B.n390 VSUBS 0.007654f
C755 B.n391 VSUBS 0.007654f
C756 B.n392 VSUBS 0.007654f
C757 B.n393 VSUBS 0.007654f
C758 B.n394 VSUBS 0.007654f
C759 B.n395 VSUBS 0.007654f
C760 B.n396 VSUBS 0.007654f
C761 B.n397 VSUBS 0.007654f
C762 B.n398 VSUBS 0.007654f
C763 B.n399 VSUBS 0.007654f
C764 B.n400 VSUBS 0.007654f
C765 B.n401 VSUBS 0.007654f
C766 B.n402 VSUBS 0.007654f
C767 B.n403 VSUBS 0.007654f
C768 B.n404 VSUBS 0.007654f
C769 B.n405 VSUBS 0.007654f
C770 B.n406 VSUBS 0.007654f
C771 B.n407 VSUBS 0.007654f
C772 B.n408 VSUBS 0.007654f
C773 B.n409 VSUBS 0.007654f
C774 B.n410 VSUBS 0.007654f
C775 B.n411 VSUBS 0.007654f
C776 B.n412 VSUBS 0.007654f
C777 B.n413 VSUBS 0.007654f
C778 B.n414 VSUBS 0.007654f
C779 B.n415 VSUBS 0.007654f
C780 B.n416 VSUBS 0.007654f
C781 B.n417 VSUBS 0.007654f
C782 B.n418 VSUBS 0.007654f
C783 B.n419 VSUBS 0.007654f
C784 B.n420 VSUBS 0.007654f
C785 B.n421 VSUBS 0.007654f
C786 B.n422 VSUBS 0.007654f
C787 B.n423 VSUBS 0.007654f
C788 B.n424 VSUBS 0.007654f
C789 B.n425 VSUBS 0.007654f
C790 B.n426 VSUBS 0.007654f
C791 B.n427 VSUBS 0.007654f
C792 B.n428 VSUBS 0.007654f
C793 B.n429 VSUBS 0.007654f
C794 B.n430 VSUBS 0.007654f
C795 B.n431 VSUBS 0.007654f
C796 B.n432 VSUBS 0.007654f
C797 B.n433 VSUBS 0.007654f
C798 B.n434 VSUBS 0.007654f
C799 B.n435 VSUBS 0.007654f
C800 B.n436 VSUBS 0.007654f
C801 B.n437 VSUBS 0.018824f
C802 B.n438 VSUBS 0.019444f
C803 B.n439 VSUBS 0.019444f
C804 B.n440 VSUBS 0.007654f
C805 B.n441 VSUBS 0.007654f
C806 B.n442 VSUBS 0.007654f
C807 B.n443 VSUBS 0.007654f
C808 B.n444 VSUBS 0.007654f
C809 B.n445 VSUBS 0.007654f
C810 B.n446 VSUBS 0.007654f
C811 B.n447 VSUBS 0.007654f
C812 B.n448 VSUBS 0.007654f
C813 B.n449 VSUBS 0.007654f
C814 B.n450 VSUBS 0.007654f
C815 B.n451 VSUBS 0.007654f
C816 B.n452 VSUBS 0.007654f
C817 B.n453 VSUBS 0.007654f
C818 B.n454 VSUBS 0.007654f
C819 B.n455 VSUBS 0.007654f
C820 B.n456 VSUBS 0.007654f
C821 B.n457 VSUBS 0.007654f
C822 B.n458 VSUBS 0.007654f
C823 B.n459 VSUBS 0.007654f
C824 B.n460 VSUBS 0.007654f
C825 B.n461 VSUBS 0.007654f
C826 B.n462 VSUBS 0.007654f
C827 B.n463 VSUBS 0.007654f
C828 B.n464 VSUBS 0.007654f
C829 B.n465 VSUBS 0.007654f
C830 B.n466 VSUBS 0.007654f
C831 B.n467 VSUBS 0.007654f
C832 B.n468 VSUBS 0.007654f
C833 B.n469 VSUBS 0.007654f
C834 B.n470 VSUBS 0.007654f
C835 B.n471 VSUBS 0.007654f
C836 B.n472 VSUBS 0.007654f
C837 B.n473 VSUBS 0.007654f
C838 B.n474 VSUBS 0.007203f
C839 B.n475 VSUBS 0.007654f
C840 B.n476 VSUBS 0.007654f
C841 B.n477 VSUBS 0.007654f
C842 B.n478 VSUBS 0.007654f
C843 B.n479 VSUBS 0.007654f
C844 B.n480 VSUBS 0.007654f
C845 B.n481 VSUBS 0.007654f
C846 B.n482 VSUBS 0.007654f
C847 B.n483 VSUBS 0.007654f
C848 B.n484 VSUBS 0.007654f
C849 B.n485 VSUBS 0.007654f
C850 B.n486 VSUBS 0.007654f
C851 B.n487 VSUBS 0.007654f
C852 B.n488 VSUBS 0.007654f
C853 B.n489 VSUBS 0.007654f
C854 B.n490 VSUBS 0.004277f
C855 B.n491 VSUBS 0.017733f
C856 B.n492 VSUBS 0.007203f
C857 B.n493 VSUBS 0.007654f
C858 B.n494 VSUBS 0.007654f
C859 B.n495 VSUBS 0.007654f
C860 B.n496 VSUBS 0.007654f
C861 B.n497 VSUBS 0.007654f
C862 B.n498 VSUBS 0.007654f
C863 B.n499 VSUBS 0.007654f
C864 B.n500 VSUBS 0.007654f
C865 B.n501 VSUBS 0.007654f
C866 B.n502 VSUBS 0.007654f
C867 B.n503 VSUBS 0.007654f
C868 B.n504 VSUBS 0.007654f
C869 B.n505 VSUBS 0.007654f
C870 B.n506 VSUBS 0.007654f
C871 B.n507 VSUBS 0.007654f
C872 B.n508 VSUBS 0.007654f
C873 B.n509 VSUBS 0.007654f
C874 B.n510 VSUBS 0.007654f
C875 B.n511 VSUBS 0.007654f
C876 B.n512 VSUBS 0.007654f
C877 B.n513 VSUBS 0.007654f
C878 B.n514 VSUBS 0.007654f
C879 B.n515 VSUBS 0.007654f
C880 B.n516 VSUBS 0.007654f
C881 B.n517 VSUBS 0.007654f
C882 B.n518 VSUBS 0.007654f
C883 B.n519 VSUBS 0.007654f
C884 B.n520 VSUBS 0.007654f
C885 B.n521 VSUBS 0.007654f
C886 B.n522 VSUBS 0.007654f
C887 B.n523 VSUBS 0.007654f
C888 B.n524 VSUBS 0.007654f
C889 B.n525 VSUBS 0.007654f
C890 B.n526 VSUBS 0.007654f
C891 B.n527 VSUBS 0.007654f
C892 B.n528 VSUBS 0.019444f
C893 B.n529 VSUBS 0.018824f
C894 B.n530 VSUBS 0.018824f
C895 B.n531 VSUBS 0.007654f
C896 B.n532 VSUBS 0.007654f
C897 B.n533 VSUBS 0.007654f
C898 B.n534 VSUBS 0.007654f
C899 B.n535 VSUBS 0.007654f
C900 B.n536 VSUBS 0.007654f
C901 B.n537 VSUBS 0.007654f
C902 B.n538 VSUBS 0.007654f
C903 B.n539 VSUBS 0.007654f
C904 B.n540 VSUBS 0.007654f
C905 B.n541 VSUBS 0.007654f
C906 B.n542 VSUBS 0.007654f
C907 B.n543 VSUBS 0.007654f
C908 B.n544 VSUBS 0.007654f
C909 B.n545 VSUBS 0.007654f
C910 B.n546 VSUBS 0.007654f
C911 B.n547 VSUBS 0.007654f
C912 B.n548 VSUBS 0.007654f
C913 B.n549 VSUBS 0.007654f
C914 B.n550 VSUBS 0.007654f
C915 B.n551 VSUBS 0.007654f
C916 B.n552 VSUBS 0.007654f
C917 B.n553 VSUBS 0.007654f
C918 B.n554 VSUBS 0.007654f
C919 B.n555 VSUBS 0.007654f
C920 B.n556 VSUBS 0.007654f
C921 B.n557 VSUBS 0.007654f
C922 B.n558 VSUBS 0.007654f
C923 B.n559 VSUBS 0.007654f
C924 B.n560 VSUBS 0.007654f
C925 B.n561 VSUBS 0.007654f
C926 B.n562 VSUBS 0.007654f
C927 B.n563 VSUBS 0.007654f
C928 B.n564 VSUBS 0.007654f
C929 B.n565 VSUBS 0.007654f
C930 B.n566 VSUBS 0.007654f
C931 B.n567 VSUBS 0.007654f
C932 B.n568 VSUBS 0.007654f
C933 B.n569 VSUBS 0.007654f
C934 B.n570 VSUBS 0.007654f
C935 B.n571 VSUBS 0.007654f
C936 B.n572 VSUBS 0.007654f
C937 B.n573 VSUBS 0.007654f
C938 B.n574 VSUBS 0.007654f
C939 B.n575 VSUBS 0.007654f
C940 B.n576 VSUBS 0.007654f
C941 B.n577 VSUBS 0.007654f
C942 B.n578 VSUBS 0.007654f
C943 B.n579 VSUBS 0.007654f
C944 B.n580 VSUBS 0.007654f
C945 B.n581 VSUBS 0.007654f
C946 B.n582 VSUBS 0.007654f
C947 B.n583 VSUBS 0.007654f
C948 B.n584 VSUBS 0.007654f
C949 B.n585 VSUBS 0.007654f
C950 B.n586 VSUBS 0.007654f
C951 B.n587 VSUBS 0.007654f
C952 B.n588 VSUBS 0.007654f
C953 B.n589 VSUBS 0.007654f
C954 B.n590 VSUBS 0.007654f
C955 B.n591 VSUBS 0.009988f
C956 B.n592 VSUBS 0.010639f
C957 B.n593 VSUBS 0.021157f
.ends

