* NGSPICE file created from diff_pair_sample_0664.ext - technology: sky130A

.subckt diff_pair_sample_0664 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=0 ps=0 w=8.7 l=0.29
X1 VDD2.t9 VN.t0 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=1.4355 ps=9.03 w=8.7 l=0.29
X2 VTAIL.t6 VP.t0 VDD1.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X3 VDD2.t8 VN.t1 VTAIL.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X4 VDD1.t8 VP.t1 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=3.393 ps=18.18 w=8.7 l=0.29
X5 VDD2.t7 VN.t2 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=1.4355 ps=9.03 w=8.7 l=0.29
X6 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=0 ps=0 w=8.7 l=0.29
X7 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=0 ps=0 w=8.7 l=0.29
X8 VTAIL.t1 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X9 VTAIL.t11 VN.t3 VDD2.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X10 VTAIL.t12 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X11 VTAIL.t13 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X12 VDD1.t6 VP.t3 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=3.393 ps=18.18 w=8.7 l=0.29
X13 VDD1.t5 VP.t4 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=1.4355 ps=9.03 w=8.7 l=0.29
X14 VDD2.t3 VN.t6 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=3.393 ps=18.18 w=8.7 l=0.29
X15 VDD1.t4 VP.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=1.4355 ps=9.03 w=8.7 l=0.29
X16 VDD1.t3 VP.t6 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X17 VTAIL.t7 VN.t7 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X18 VDD2.t1 VN.t8 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X19 VDD1.t2 VP.t7 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X20 VTAIL.t18 VP.t8 VDD1.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X21 VTAIL.t19 VP.t9 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=1.4355 ps=9.03 w=8.7 l=0.29
X22 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.393 pd=18.18 as=0 ps=0 w=8.7 l=0.29
X23 VDD2.t0 VN.t9 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4355 pd=9.03 as=3.393 ps=18.18 w=8.7 l=0.29
R0 B.n294 B.t14 940.653
R1 B.n292 B.t10 940.653
R2 B.n78 B.t21 940.653
R3 B.n76 B.t17 940.653
R4 B.n528 B.n527 585
R5 B.n529 B.n528 585
R6 B.n220 B.n74 585
R7 B.n219 B.n218 585
R8 B.n217 B.n216 585
R9 B.n215 B.n214 585
R10 B.n213 B.n212 585
R11 B.n211 B.n210 585
R12 B.n209 B.n208 585
R13 B.n207 B.n206 585
R14 B.n205 B.n204 585
R15 B.n203 B.n202 585
R16 B.n201 B.n200 585
R17 B.n199 B.n198 585
R18 B.n197 B.n196 585
R19 B.n195 B.n194 585
R20 B.n193 B.n192 585
R21 B.n191 B.n190 585
R22 B.n189 B.n188 585
R23 B.n187 B.n186 585
R24 B.n185 B.n184 585
R25 B.n183 B.n182 585
R26 B.n181 B.n180 585
R27 B.n179 B.n178 585
R28 B.n177 B.n176 585
R29 B.n175 B.n174 585
R30 B.n173 B.n172 585
R31 B.n171 B.n170 585
R32 B.n169 B.n168 585
R33 B.n167 B.n166 585
R34 B.n165 B.n164 585
R35 B.n163 B.n162 585
R36 B.n161 B.n160 585
R37 B.n158 B.n157 585
R38 B.n156 B.n155 585
R39 B.n154 B.n153 585
R40 B.n152 B.n151 585
R41 B.n150 B.n149 585
R42 B.n148 B.n147 585
R43 B.n146 B.n145 585
R44 B.n144 B.n143 585
R45 B.n142 B.n141 585
R46 B.n140 B.n139 585
R47 B.n138 B.n137 585
R48 B.n136 B.n135 585
R49 B.n134 B.n133 585
R50 B.n132 B.n131 585
R51 B.n130 B.n129 585
R52 B.n128 B.n127 585
R53 B.n126 B.n125 585
R54 B.n124 B.n123 585
R55 B.n122 B.n121 585
R56 B.n120 B.n119 585
R57 B.n118 B.n117 585
R58 B.n116 B.n115 585
R59 B.n114 B.n113 585
R60 B.n112 B.n111 585
R61 B.n110 B.n109 585
R62 B.n108 B.n107 585
R63 B.n106 B.n105 585
R64 B.n104 B.n103 585
R65 B.n102 B.n101 585
R66 B.n100 B.n99 585
R67 B.n98 B.n97 585
R68 B.n96 B.n95 585
R69 B.n94 B.n93 585
R70 B.n92 B.n91 585
R71 B.n90 B.n89 585
R72 B.n88 B.n87 585
R73 B.n86 B.n85 585
R74 B.n84 B.n83 585
R75 B.n82 B.n81 585
R76 B.n38 B.n37 585
R77 B.n532 B.n531 585
R78 B.n526 B.n75 585
R79 B.n75 B.n35 585
R80 B.n525 B.n34 585
R81 B.n536 B.n34 585
R82 B.n524 B.n33 585
R83 B.n537 B.n33 585
R84 B.n523 B.n32 585
R85 B.n538 B.n32 585
R86 B.n522 B.n521 585
R87 B.n521 B.n31 585
R88 B.n520 B.n27 585
R89 B.n544 B.n27 585
R90 B.n519 B.n26 585
R91 B.n545 B.n26 585
R92 B.n518 B.n25 585
R93 B.n546 B.n25 585
R94 B.n517 B.n516 585
R95 B.n516 B.n21 585
R96 B.n515 B.n20 585
R97 B.n552 B.n20 585
R98 B.n514 B.n19 585
R99 B.n553 B.n19 585
R100 B.n513 B.n18 585
R101 B.n554 B.n18 585
R102 B.n512 B.n511 585
R103 B.n511 B.n510 585
R104 B.n509 B.n14 585
R105 B.n560 B.n14 585
R106 B.n508 B.n13 585
R107 B.n561 B.n13 585
R108 B.n507 B.n12 585
R109 B.n562 B.n12 585
R110 B.n506 B.n505 585
R111 B.n505 B.n11 585
R112 B.n504 B.n7 585
R113 B.n568 B.n7 585
R114 B.n503 B.n6 585
R115 B.n569 B.n6 585
R116 B.n502 B.n5 585
R117 B.n570 B.n5 585
R118 B.n501 B.n500 585
R119 B.n500 B.n4 585
R120 B.n499 B.n221 585
R121 B.n499 B.n498 585
R122 B.n488 B.n222 585
R123 B.n491 B.n222 585
R124 B.n490 B.n489 585
R125 B.n492 B.n490 585
R126 B.n487 B.n226 585
R127 B.n229 B.n226 585
R128 B.n486 B.n485 585
R129 B.n485 B.n484 585
R130 B.n228 B.n227 585
R131 B.n477 B.n228 585
R132 B.n476 B.n475 585
R133 B.n478 B.n476 585
R134 B.n474 B.n234 585
R135 B.n234 B.n233 585
R136 B.n473 B.n472 585
R137 B.n472 B.n471 585
R138 B.n236 B.n235 585
R139 B.n237 B.n236 585
R140 B.n464 B.n463 585
R141 B.n465 B.n464 585
R142 B.n462 B.n242 585
R143 B.n242 B.n241 585
R144 B.n461 B.n460 585
R145 B.n460 B.n459 585
R146 B.n244 B.n243 585
R147 B.n452 B.n244 585
R148 B.n451 B.n450 585
R149 B.n453 B.n451 585
R150 B.n449 B.n249 585
R151 B.n249 B.n248 585
R152 B.n448 B.n447 585
R153 B.n447 B.n446 585
R154 B.n251 B.n250 585
R155 B.n252 B.n251 585
R156 B.n442 B.n441 585
R157 B.n255 B.n254 585
R158 B.n438 B.n437 585
R159 B.n439 B.n438 585
R160 B.n436 B.n291 585
R161 B.n435 B.n434 585
R162 B.n433 B.n432 585
R163 B.n431 B.n430 585
R164 B.n429 B.n428 585
R165 B.n427 B.n426 585
R166 B.n425 B.n424 585
R167 B.n423 B.n422 585
R168 B.n421 B.n420 585
R169 B.n419 B.n418 585
R170 B.n417 B.n416 585
R171 B.n415 B.n414 585
R172 B.n413 B.n412 585
R173 B.n411 B.n410 585
R174 B.n409 B.n408 585
R175 B.n407 B.n406 585
R176 B.n405 B.n404 585
R177 B.n403 B.n402 585
R178 B.n401 B.n400 585
R179 B.n399 B.n398 585
R180 B.n397 B.n396 585
R181 B.n395 B.n394 585
R182 B.n393 B.n392 585
R183 B.n391 B.n390 585
R184 B.n389 B.n388 585
R185 B.n387 B.n386 585
R186 B.n385 B.n384 585
R187 B.n383 B.n382 585
R188 B.n381 B.n380 585
R189 B.n378 B.n377 585
R190 B.n376 B.n375 585
R191 B.n374 B.n373 585
R192 B.n372 B.n371 585
R193 B.n370 B.n369 585
R194 B.n368 B.n367 585
R195 B.n366 B.n365 585
R196 B.n364 B.n363 585
R197 B.n362 B.n361 585
R198 B.n360 B.n359 585
R199 B.n358 B.n357 585
R200 B.n356 B.n355 585
R201 B.n354 B.n353 585
R202 B.n352 B.n351 585
R203 B.n350 B.n349 585
R204 B.n348 B.n347 585
R205 B.n346 B.n345 585
R206 B.n344 B.n343 585
R207 B.n342 B.n341 585
R208 B.n340 B.n339 585
R209 B.n338 B.n337 585
R210 B.n336 B.n335 585
R211 B.n334 B.n333 585
R212 B.n332 B.n331 585
R213 B.n330 B.n329 585
R214 B.n328 B.n327 585
R215 B.n326 B.n325 585
R216 B.n324 B.n323 585
R217 B.n322 B.n321 585
R218 B.n320 B.n319 585
R219 B.n318 B.n317 585
R220 B.n316 B.n315 585
R221 B.n314 B.n313 585
R222 B.n312 B.n311 585
R223 B.n310 B.n309 585
R224 B.n308 B.n307 585
R225 B.n306 B.n305 585
R226 B.n304 B.n303 585
R227 B.n302 B.n301 585
R228 B.n300 B.n299 585
R229 B.n298 B.n297 585
R230 B.n443 B.n253 585
R231 B.n253 B.n252 585
R232 B.n445 B.n444 585
R233 B.n446 B.n445 585
R234 B.n247 B.n246 585
R235 B.n248 B.n247 585
R236 B.n455 B.n454 585
R237 B.n454 B.n453 585
R238 B.n456 B.n245 585
R239 B.n452 B.n245 585
R240 B.n458 B.n457 585
R241 B.n459 B.n458 585
R242 B.n240 B.n239 585
R243 B.n241 B.n240 585
R244 B.n467 B.n466 585
R245 B.n466 B.n465 585
R246 B.n468 B.n238 585
R247 B.n238 B.n237 585
R248 B.n470 B.n469 585
R249 B.n471 B.n470 585
R250 B.n232 B.n231 585
R251 B.n233 B.n232 585
R252 B.n480 B.n479 585
R253 B.n479 B.n478 585
R254 B.n481 B.n230 585
R255 B.n477 B.n230 585
R256 B.n483 B.n482 585
R257 B.n484 B.n483 585
R258 B.n225 B.n224 585
R259 B.n229 B.n225 585
R260 B.n494 B.n493 585
R261 B.n493 B.n492 585
R262 B.n495 B.n223 585
R263 B.n491 B.n223 585
R264 B.n497 B.n496 585
R265 B.n498 B.n497 585
R266 B.n2 B.n0 585
R267 B.n4 B.n2 585
R268 B.n3 B.n1 585
R269 B.n569 B.n3 585
R270 B.n567 B.n566 585
R271 B.n568 B.n567 585
R272 B.n565 B.n8 585
R273 B.n11 B.n8 585
R274 B.n564 B.n563 585
R275 B.n563 B.n562 585
R276 B.n10 B.n9 585
R277 B.n561 B.n10 585
R278 B.n559 B.n558 585
R279 B.n560 B.n559 585
R280 B.n557 B.n15 585
R281 B.n510 B.n15 585
R282 B.n556 B.n555 585
R283 B.n555 B.n554 585
R284 B.n17 B.n16 585
R285 B.n553 B.n17 585
R286 B.n551 B.n550 585
R287 B.n552 B.n551 585
R288 B.n549 B.n22 585
R289 B.n22 B.n21 585
R290 B.n548 B.n547 585
R291 B.n547 B.n546 585
R292 B.n24 B.n23 585
R293 B.n545 B.n24 585
R294 B.n543 B.n542 585
R295 B.n544 B.n543 585
R296 B.n541 B.n28 585
R297 B.n31 B.n28 585
R298 B.n540 B.n539 585
R299 B.n539 B.n538 585
R300 B.n30 B.n29 585
R301 B.n537 B.n30 585
R302 B.n535 B.n534 585
R303 B.n536 B.n535 585
R304 B.n533 B.n36 585
R305 B.n36 B.n35 585
R306 B.n572 B.n571 585
R307 B.n571 B.n570 585
R308 B.n441 B.n253 540.549
R309 B.n531 B.n36 540.549
R310 B.n297 B.n251 540.549
R311 B.n528 B.n75 540.549
R312 B.n529 B.n73 256.663
R313 B.n529 B.n72 256.663
R314 B.n529 B.n71 256.663
R315 B.n529 B.n70 256.663
R316 B.n529 B.n69 256.663
R317 B.n529 B.n68 256.663
R318 B.n529 B.n67 256.663
R319 B.n529 B.n66 256.663
R320 B.n529 B.n65 256.663
R321 B.n529 B.n64 256.663
R322 B.n529 B.n63 256.663
R323 B.n529 B.n62 256.663
R324 B.n529 B.n61 256.663
R325 B.n529 B.n60 256.663
R326 B.n529 B.n59 256.663
R327 B.n529 B.n58 256.663
R328 B.n529 B.n57 256.663
R329 B.n529 B.n56 256.663
R330 B.n529 B.n55 256.663
R331 B.n529 B.n54 256.663
R332 B.n529 B.n53 256.663
R333 B.n529 B.n52 256.663
R334 B.n529 B.n51 256.663
R335 B.n529 B.n50 256.663
R336 B.n529 B.n49 256.663
R337 B.n529 B.n48 256.663
R338 B.n529 B.n47 256.663
R339 B.n529 B.n46 256.663
R340 B.n529 B.n45 256.663
R341 B.n529 B.n44 256.663
R342 B.n529 B.n43 256.663
R343 B.n529 B.n42 256.663
R344 B.n529 B.n41 256.663
R345 B.n529 B.n40 256.663
R346 B.n529 B.n39 256.663
R347 B.n530 B.n529 256.663
R348 B.n440 B.n439 256.663
R349 B.n439 B.n256 256.663
R350 B.n439 B.n257 256.663
R351 B.n439 B.n258 256.663
R352 B.n439 B.n259 256.663
R353 B.n439 B.n260 256.663
R354 B.n439 B.n261 256.663
R355 B.n439 B.n262 256.663
R356 B.n439 B.n263 256.663
R357 B.n439 B.n264 256.663
R358 B.n439 B.n265 256.663
R359 B.n439 B.n266 256.663
R360 B.n439 B.n267 256.663
R361 B.n439 B.n268 256.663
R362 B.n439 B.n269 256.663
R363 B.n439 B.n270 256.663
R364 B.n439 B.n271 256.663
R365 B.n439 B.n272 256.663
R366 B.n439 B.n273 256.663
R367 B.n439 B.n274 256.663
R368 B.n439 B.n275 256.663
R369 B.n439 B.n276 256.663
R370 B.n439 B.n277 256.663
R371 B.n439 B.n278 256.663
R372 B.n439 B.n279 256.663
R373 B.n439 B.n280 256.663
R374 B.n439 B.n281 256.663
R375 B.n439 B.n282 256.663
R376 B.n439 B.n283 256.663
R377 B.n439 B.n284 256.663
R378 B.n439 B.n285 256.663
R379 B.n439 B.n286 256.663
R380 B.n439 B.n287 256.663
R381 B.n439 B.n288 256.663
R382 B.n439 B.n289 256.663
R383 B.n439 B.n290 256.663
R384 B.n294 B.t16 237.412
R385 B.n76 B.t19 237.412
R386 B.n292 B.t13 237.412
R387 B.n78 B.t22 237.412
R388 B.n295 B.t15 225.388
R389 B.n77 B.t20 225.388
R390 B.n293 B.t12 225.388
R391 B.n79 B.t23 225.388
R392 B.n445 B.n253 163.367
R393 B.n445 B.n247 163.367
R394 B.n454 B.n247 163.367
R395 B.n454 B.n245 163.367
R396 B.n458 B.n245 163.367
R397 B.n458 B.n240 163.367
R398 B.n466 B.n240 163.367
R399 B.n466 B.n238 163.367
R400 B.n470 B.n238 163.367
R401 B.n470 B.n232 163.367
R402 B.n479 B.n232 163.367
R403 B.n479 B.n230 163.367
R404 B.n483 B.n230 163.367
R405 B.n483 B.n225 163.367
R406 B.n493 B.n225 163.367
R407 B.n493 B.n223 163.367
R408 B.n497 B.n223 163.367
R409 B.n497 B.n2 163.367
R410 B.n571 B.n2 163.367
R411 B.n571 B.n3 163.367
R412 B.n567 B.n3 163.367
R413 B.n567 B.n8 163.367
R414 B.n563 B.n8 163.367
R415 B.n563 B.n10 163.367
R416 B.n559 B.n10 163.367
R417 B.n559 B.n15 163.367
R418 B.n555 B.n15 163.367
R419 B.n555 B.n17 163.367
R420 B.n551 B.n17 163.367
R421 B.n551 B.n22 163.367
R422 B.n547 B.n22 163.367
R423 B.n547 B.n24 163.367
R424 B.n543 B.n24 163.367
R425 B.n543 B.n28 163.367
R426 B.n539 B.n28 163.367
R427 B.n539 B.n30 163.367
R428 B.n535 B.n30 163.367
R429 B.n535 B.n36 163.367
R430 B.n438 B.n255 163.367
R431 B.n438 B.n291 163.367
R432 B.n434 B.n433 163.367
R433 B.n430 B.n429 163.367
R434 B.n426 B.n425 163.367
R435 B.n422 B.n421 163.367
R436 B.n418 B.n417 163.367
R437 B.n414 B.n413 163.367
R438 B.n410 B.n409 163.367
R439 B.n406 B.n405 163.367
R440 B.n402 B.n401 163.367
R441 B.n398 B.n397 163.367
R442 B.n394 B.n393 163.367
R443 B.n390 B.n389 163.367
R444 B.n386 B.n385 163.367
R445 B.n382 B.n381 163.367
R446 B.n377 B.n376 163.367
R447 B.n373 B.n372 163.367
R448 B.n369 B.n368 163.367
R449 B.n365 B.n364 163.367
R450 B.n361 B.n360 163.367
R451 B.n357 B.n356 163.367
R452 B.n353 B.n352 163.367
R453 B.n349 B.n348 163.367
R454 B.n345 B.n344 163.367
R455 B.n341 B.n340 163.367
R456 B.n337 B.n336 163.367
R457 B.n333 B.n332 163.367
R458 B.n329 B.n328 163.367
R459 B.n325 B.n324 163.367
R460 B.n321 B.n320 163.367
R461 B.n317 B.n316 163.367
R462 B.n313 B.n312 163.367
R463 B.n309 B.n308 163.367
R464 B.n305 B.n304 163.367
R465 B.n301 B.n300 163.367
R466 B.n447 B.n251 163.367
R467 B.n447 B.n249 163.367
R468 B.n451 B.n249 163.367
R469 B.n451 B.n244 163.367
R470 B.n460 B.n244 163.367
R471 B.n460 B.n242 163.367
R472 B.n464 B.n242 163.367
R473 B.n464 B.n236 163.367
R474 B.n472 B.n236 163.367
R475 B.n472 B.n234 163.367
R476 B.n476 B.n234 163.367
R477 B.n476 B.n228 163.367
R478 B.n485 B.n228 163.367
R479 B.n485 B.n226 163.367
R480 B.n490 B.n226 163.367
R481 B.n490 B.n222 163.367
R482 B.n499 B.n222 163.367
R483 B.n500 B.n499 163.367
R484 B.n500 B.n5 163.367
R485 B.n6 B.n5 163.367
R486 B.n7 B.n6 163.367
R487 B.n505 B.n7 163.367
R488 B.n505 B.n12 163.367
R489 B.n13 B.n12 163.367
R490 B.n14 B.n13 163.367
R491 B.n511 B.n14 163.367
R492 B.n511 B.n18 163.367
R493 B.n19 B.n18 163.367
R494 B.n20 B.n19 163.367
R495 B.n516 B.n20 163.367
R496 B.n516 B.n25 163.367
R497 B.n26 B.n25 163.367
R498 B.n27 B.n26 163.367
R499 B.n521 B.n27 163.367
R500 B.n521 B.n32 163.367
R501 B.n33 B.n32 163.367
R502 B.n34 B.n33 163.367
R503 B.n75 B.n34 163.367
R504 B.n81 B.n38 163.367
R505 B.n85 B.n84 163.367
R506 B.n89 B.n88 163.367
R507 B.n93 B.n92 163.367
R508 B.n97 B.n96 163.367
R509 B.n101 B.n100 163.367
R510 B.n105 B.n104 163.367
R511 B.n109 B.n108 163.367
R512 B.n113 B.n112 163.367
R513 B.n117 B.n116 163.367
R514 B.n121 B.n120 163.367
R515 B.n125 B.n124 163.367
R516 B.n129 B.n128 163.367
R517 B.n133 B.n132 163.367
R518 B.n137 B.n136 163.367
R519 B.n141 B.n140 163.367
R520 B.n145 B.n144 163.367
R521 B.n149 B.n148 163.367
R522 B.n153 B.n152 163.367
R523 B.n157 B.n156 163.367
R524 B.n162 B.n161 163.367
R525 B.n166 B.n165 163.367
R526 B.n170 B.n169 163.367
R527 B.n174 B.n173 163.367
R528 B.n178 B.n177 163.367
R529 B.n182 B.n181 163.367
R530 B.n186 B.n185 163.367
R531 B.n190 B.n189 163.367
R532 B.n194 B.n193 163.367
R533 B.n198 B.n197 163.367
R534 B.n202 B.n201 163.367
R535 B.n206 B.n205 163.367
R536 B.n210 B.n209 163.367
R537 B.n214 B.n213 163.367
R538 B.n218 B.n217 163.367
R539 B.n528 B.n74 163.367
R540 B.n439 B.n252 99.9647
R541 B.n529 B.n35 99.9647
R542 B.n441 B.n440 71.676
R543 B.n291 B.n256 71.676
R544 B.n433 B.n257 71.676
R545 B.n429 B.n258 71.676
R546 B.n425 B.n259 71.676
R547 B.n421 B.n260 71.676
R548 B.n417 B.n261 71.676
R549 B.n413 B.n262 71.676
R550 B.n409 B.n263 71.676
R551 B.n405 B.n264 71.676
R552 B.n401 B.n265 71.676
R553 B.n397 B.n266 71.676
R554 B.n393 B.n267 71.676
R555 B.n389 B.n268 71.676
R556 B.n385 B.n269 71.676
R557 B.n381 B.n270 71.676
R558 B.n376 B.n271 71.676
R559 B.n372 B.n272 71.676
R560 B.n368 B.n273 71.676
R561 B.n364 B.n274 71.676
R562 B.n360 B.n275 71.676
R563 B.n356 B.n276 71.676
R564 B.n352 B.n277 71.676
R565 B.n348 B.n278 71.676
R566 B.n344 B.n279 71.676
R567 B.n340 B.n280 71.676
R568 B.n336 B.n281 71.676
R569 B.n332 B.n282 71.676
R570 B.n328 B.n283 71.676
R571 B.n324 B.n284 71.676
R572 B.n320 B.n285 71.676
R573 B.n316 B.n286 71.676
R574 B.n312 B.n287 71.676
R575 B.n308 B.n288 71.676
R576 B.n304 B.n289 71.676
R577 B.n300 B.n290 71.676
R578 B.n531 B.n530 71.676
R579 B.n81 B.n39 71.676
R580 B.n85 B.n40 71.676
R581 B.n89 B.n41 71.676
R582 B.n93 B.n42 71.676
R583 B.n97 B.n43 71.676
R584 B.n101 B.n44 71.676
R585 B.n105 B.n45 71.676
R586 B.n109 B.n46 71.676
R587 B.n113 B.n47 71.676
R588 B.n117 B.n48 71.676
R589 B.n121 B.n49 71.676
R590 B.n125 B.n50 71.676
R591 B.n129 B.n51 71.676
R592 B.n133 B.n52 71.676
R593 B.n137 B.n53 71.676
R594 B.n141 B.n54 71.676
R595 B.n145 B.n55 71.676
R596 B.n149 B.n56 71.676
R597 B.n153 B.n57 71.676
R598 B.n157 B.n58 71.676
R599 B.n162 B.n59 71.676
R600 B.n166 B.n60 71.676
R601 B.n170 B.n61 71.676
R602 B.n174 B.n62 71.676
R603 B.n178 B.n63 71.676
R604 B.n182 B.n64 71.676
R605 B.n186 B.n65 71.676
R606 B.n190 B.n66 71.676
R607 B.n194 B.n67 71.676
R608 B.n198 B.n68 71.676
R609 B.n202 B.n69 71.676
R610 B.n206 B.n70 71.676
R611 B.n210 B.n71 71.676
R612 B.n214 B.n72 71.676
R613 B.n218 B.n73 71.676
R614 B.n74 B.n73 71.676
R615 B.n217 B.n72 71.676
R616 B.n213 B.n71 71.676
R617 B.n209 B.n70 71.676
R618 B.n205 B.n69 71.676
R619 B.n201 B.n68 71.676
R620 B.n197 B.n67 71.676
R621 B.n193 B.n66 71.676
R622 B.n189 B.n65 71.676
R623 B.n185 B.n64 71.676
R624 B.n181 B.n63 71.676
R625 B.n177 B.n62 71.676
R626 B.n173 B.n61 71.676
R627 B.n169 B.n60 71.676
R628 B.n165 B.n59 71.676
R629 B.n161 B.n58 71.676
R630 B.n156 B.n57 71.676
R631 B.n152 B.n56 71.676
R632 B.n148 B.n55 71.676
R633 B.n144 B.n54 71.676
R634 B.n140 B.n53 71.676
R635 B.n136 B.n52 71.676
R636 B.n132 B.n51 71.676
R637 B.n128 B.n50 71.676
R638 B.n124 B.n49 71.676
R639 B.n120 B.n48 71.676
R640 B.n116 B.n47 71.676
R641 B.n112 B.n46 71.676
R642 B.n108 B.n45 71.676
R643 B.n104 B.n44 71.676
R644 B.n100 B.n43 71.676
R645 B.n96 B.n42 71.676
R646 B.n92 B.n41 71.676
R647 B.n88 B.n40 71.676
R648 B.n84 B.n39 71.676
R649 B.n530 B.n38 71.676
R650 B.n440 B.n255 71.676
R651 B.n434 B.n256 71.676
R652 B.n430 B.n257 71.676
R653 B.n426 B.n258 71.676
R654 B.n422 B.n259 71.676
R655 B.n418 B.n260 71.676
R656 B.n414 B.n261 71.676
R657 B.n410 B.n262 71.676
R658 B.n406 B.n263 71.676
R659 B.n402 B.n264 71.676
R660 B.n398 B.n265 71.676
R661 B.n394 B.n266 71.676
R662 B.n390 B.n267 71.676
R663 B.n386 B.n268 71.676
R664 B.n382 B.n269 71.676
R665 B.n377 B.n270 71.676
R666 B.n373 B.n271 71.676
R667 B.n369 B.n272 71.676
R668 B.n365 B.n273 71.676
R669 B.n361 B.n274 71.676
R670 B.n357 B.n275 71.676
R671 B.n353 B.n276 71.676
R672 B.n349 B.n277 71.676
R673 B.n345 B.n278 71.676
R674 B.n341 B.n279 71.676
R675 B.n337 B.n280 71.676
R676 B.n333 B.n281 71.676
R677 B.n329 B.n282 71.676
R678 B.n325 B.n283 71.676
R679 B.n321 B.n284 71.676
R680 B.n317 B.n285 71.676
R681 B.n313 B.n286 71.676
R682 B.n309 B.n287 71.676
R683 B.n305 B.n288 71.676
R684 B.n301 B.n289 71.676
R685 B.n297 B.n290 71.676
R686 B.n296 B.n295 59.5399
R687 B.n379 B.n293 59.5399
R688 B.n80 B.n79 59.5399
R689 B.n159 B.n77 59.5399
R690 B.n446 B.n252 53.5246
R691 B.n446 B.n248 53.5246
R692 B.n453 B.n248 53.5246
R693 B.n453 B.n452 53.5246
R694 B.n459 B.n241 53.5246
R695 B.n465 B.n241 53.5246
R696 B.n465 B.n237 53.5246
R697 B.n471 B.n237 53.5246
R698 B.n478 B.n233 53.5246
R699 B.n484 B.n229 53.5246
R700 B.n492 B.n491 53.5246
R701 B.n498 B.n4 53.5246
R702 B.n570 B.n4 53.5246
R703 B.n570 B.n569 53.5246
R704 B.n569 B.n568 53.5246
R705 B.n562 B.n11 53.5246
R706 B.n561 B.n560 53.5246
R707 B.n554 B.n553 53.5246
R708 B.n552 B.n21 53.5246
R709 B.n546 B.n21 53.5246
R710 B.n546 B.n545 53.5246
R711 B.n545 B.n544 53.5246
R712 B.n538 B.n31 53.5246
R713 B.n538 B.n537 53.5246
R714 B.n537 B.n536 53.5246
R715 B.n536 B.n35 53.5246
R716 B.t4 B.n477 52.7375
R717 B.n510 B.t1 52.7375
R718 B.n459 B.t11 44.8663
R719 B.n477 B.t6 44.8663
R720 B.n510 B.t0 44.8663
R721 B.n544 B.t18 44.8663
R722 B.t7 B.n233 43.2921
R723 B.n553 B.t3 43.2921
R724 B.n229 B.t9 35.4209
R725 B.t8 B.n561 35.4209
R726 B.n533 B.n532 35.1225
R727 B.n527 B.n526 35.1225
R728 B.n298 B.n250 35.1225
R729 B.n443 B.n442 35.1225
R730 B.n498 B.t5 27.5497
R731 B.n568 B.t2 27.5497
R732 B.n491 B.t5 25.9755
R733 B.n11 B.t2 25.9755
R734 B.n492 B.t9 18.1043
R735 B.n562 B.t8 18.1043
R736 B B.n572 18.0485
R737 B.n295 B.n294 12.0247
R738 B.n293 B.n292 12.0247
R739 B.n79 B.n78 12.0247
R740 B.n77 B.n76 12.0247
R741 B.n532 B.n37 10.6151
R742 B.n82 B.n37 10.6151
R743 B.n83 B.n82 10.6151
R744 B.n86 B.n83 10.6151
R745 B.n87 B.n86 10.6151
R746 B.n90 B.n87 10.6151
R747 B.n91 B.n90 10.6151
R748 B.n94 B.n91 10.6151
R749 B.n95 B.n94 10.6151
R750 B.n98 B.n95 10.6151
R751 B.n99 B.n98 10.6151
R752 B.n102 B.n99 10.6151
R753 B.n103 B.n102 10.6151
R754 B.n106 B.n103 10.6151
R755 B.n107 B.n106 10.6151
R756 B.n110 B.n107 10.6151
R757 B.n111 B.n110 10.6151
R758 B.n114 B.n111 10.6151
R759 B.n115 B.n114 10.6151
R760 B.n118 B.n115 10.6151
R761 B.n119 B.n118 10.6151
R762 B.n122 B.n119 10.6151
R763 B.n123 B.n122 10.6151
R764 B.n126 B.n123 10.6151
R765 B.n127 B.n126 10.6151
R766 B.n130 B.n127 10.6151
R767 B.n131 B.n130 10.6151
R768 B.n134 B.n131 10.6151
R769 B.n135 B.n134 10.6151
R770 B.n138 B.n135 10.6151
R771 B.n139 B.n138 10.6151
R772 B.n143 B.n142 10.6151
R773 B.n146 B.n143 10.6151
R774 B.n147 B.n146 10.6151
R775 B.n150 B.n147 10.6151
R776 B.n151 B.n150 10.6151
R777 B.n154 B.n151 10.6151
R778 B.n155 B.n154 10.6151
R779 B.n158 B.n155 10.6151
R780 B.n163 B.n160 10.6151
R781 B.n164 B.n163 10.6151
R782 B.n167 B.n164 10.6151
R783 B.n168 B.n167 10.6151
R784 B.n171 B.n168 10.6151
R785 B.n172 B.n171 10.6151
R786 B.n175 B.n172 10.6151
R787 B.n176 B.n175 10.6151
R788 B.n179 B.n176 10.6151
R789 B.n180 B.n179 10.6151
R790 B.n183 B.n180 10.6151
R791 B.n184 B.n183 10.6151
R792 B.n187 B.n184 10.6151
R793 B.n188 B.n187 10.6151
R794 B.n191 B.n188 10.6151
R795 B.n192 B.n191 10.6151
R796 B.n195 B.n192 10.6151
R797 B.n196 B.n195 10.6151
R798 B.n199 B.n196 10.6151
R799 B.n200 B.n199 10.6151
R800 B.n203 B.n200 10.6151
R801 B.n204 B.n203 10.6151
R802 B.n207 B.n204 10.6151
R803 B.n208 B.n207 10.6151
R804 B.n211 B.n208 10.6151
R805 B.n212 B.n211 10.6151
R806 B.n215 B.n212 10.6151
R807 B.n216 B.n215 10.6151
R808 B.n219 B.n216 10.6151
R809 B.n220 B.n219 10.6151
R810 B.n527 B.n220 10.6151
R811 B.n448 B.n250 10.6151
R812 B.n449 B.n448 10.6151
R813 B.n450 B.n449 10.6151
R814 B.n450 B.n243 10.6151
R815 B.n461 B.n243 10.6151
R816 B.n462 B.n461 10.6151
R817 B.n463 B.n462 10.6151
R818 B.n463 B.n235 10.6151
R819 B.n473 B.n235 10.6151
R820 B.n474 B.n473 10.6151
R821 B.n475 B.n474 10.6151
R822 B.n475 B.n227 10.6151
R823 B.n486 B.n227 10.6151
R824 B.n487 B.n486 10.6151
R825 B.n489 B.n487 10.6151
R826 B.n489 B.n488 10.6151
R827 B.n488 B.n221 10.6151
R828 B.n501 B.n221 10.6151
R829 B.n502 B.n501 10.6151
R830 B.n503 B.n502 10.6151
R831 B.n504 B.n503 10.6151
R832 B.n506 B.n504 10.6151
R833 B.n507 B.n506 10.6151
R834 B.n508 B.n507 10.6151
R835 B.n509 B.n508 10.6151
R836 B.n512 B.n509 10.6151
R837 B.n513 B.n512 10.6151
R838 B.n514 B.n513 10.6151
R839 B.n515 B.n514 10.6151
R840 B.n517 B.n515 10.6151
R841 B.n518 B.n517 10.6151
R842 B.n519 B.n518 10.6151
R843 B.n520 B.n519 10.6151
R844 B.n522 B.n520 10.6151
R845 B.n523 B.n522 10.6151
R846 B.n524 B.n523 10.6151
R847 B.n525 B.n524 10.6151
R848 B.n526 B.n525 10.6151
R849 B.n442 B.n254 10.6151
R850 B.n437 B.n254 10.6151
R851 B.n437 B.n436 10.6151
R852 B.n436 B.n435 10.6151
R853 B.n435 B.n432 10.6151
R854 B.n432 B.n431 10.6151
R855 B.n431 B.n428 10.6151
R856 B.n428 B.n427 10.6151
R857 B.n427 B.n424 10.6151
R858 B.n424 B.n423 10.6151
R859 B.n423 B.n420 10.6151
R860 B.n420 B.n419 10.6151
R861 B.n419 B.n416 10.6151
R862 B.n416 B.n415 10.6151
R863 B.n415 B.n412 10.6151
R864 B.n412 B.n411 10.6151
R865 B.n411 B.n408 10.6151
R866 B.n408 B.n407 10.6151
R867 B.n407 B.n404 10.6151
R868 B.n404 B.n403 10.6151
R869 B.n403 B.n400 10.6151
R870 B.n400 B.n399 10.6151
R871 B.n399 B.n396 10.6151
R872 B.n396 B.n395 10.6151
R873 B.n395 B.n392 10.6151
R874 B.n392 B.n391 10.6151
R875 B.n391 B.n388 10.6151
R876 B.n388 B.n387 10.6151
R877 B.n387 B.n384 10.6151
R878 B.n384 B.n383 10.6151
R879 B.n383 B.n380 10.6151
R880 B.n378 B.n375 10.6151
R881 B.n375 B.n374 10.6151
R882 B.n374 B.n371 10.6151
R883 B.n371 B.n370 10.6151
R884 B.n370 B.n367 10.6151
R885 B.n367 B.n366 10.6151
R886 B.n366 B.n363 10.6151
R887 B.n363 B.n362 10.6151
R888 B.n359 B.n358 10.6151
R889 B.n358 B.n355 10.6151
R890 B.n355 B.n354 10.6151
R891 B.n354 B.n351 10.6151
R892 B.n351 B.n350 10.6151
R893 B.n350 B.n347 10.6151
R894 B.n347 B.n346 10.6151
R895 B.n346 B.n343 10.6151
R896 B.n343 B.n342 10.6151
R897 B.n342 B.n339 10.6151
R898 B.n339 B.n338 10.6151
R899 B.n338 B.n335 10.6151
R900 B.n335 B.n334 10.6151
R901 B.n334 B.n331 10.6151
R902 B.n331 B.n330 10.6151
R903 B.n330 B.n327 10.6151
R904 B.n327 B.n326 10.6151
R905 B.n326 B.n323 10.6151
R906 B.n323 B.n322 10.6151
R907 B.n322 B.n319 10.6151
R908 B.n319 B.n318 10.6151
R909 B.n318 B.n315 10.6151
R910 B.n315 B.n314 10.6151
R911 B.n314 B.n311 10.6151
R912 B.n311 B.n310 10.6151
R913 B.n310 B.n307 10.6151
R914 B.n307 B.n306 10.6151
R915 B.n306 B.n303 10.6151
R916 B.n303 B.n302 10.6151
R917 B.n302 B.n299 10.6151
R918 B.n299 B.n298 10.6151
R919 B.n444 B.n443 10.6151
R920 B.n444 B.n246 10.6151
R921 B.n455 B.n246 10.6151
R922 B.n456 B.n455 10.6151
R923 B.n457 B.n456 10.6151
R924 B.n457 B.n239 10.6151
R925 B.n467 B.n239 10.6151
R926 B.n468 B.n467 10.6151
R927 B.n469 B.n468 10.6151
R928 B.n469 B.n231 10.6151
R929 B.n480 B.n231 10.6151
R930 B.n481 B.n480 10.6151
R931 B.n482 B.n481 10.6151
R932 B.n482 B.n224 10.6151
R933 B.n494 B.n224 10.6151
R934 B.n495 B.n494 10.6151
R935 B.n496 B.n495 10.6151
R936 B.n496 B.n0 10.6151
R937 B.n566 B.n1 10.6151
R938 B.n566 B.n565 10.6151
R939 B.n565 B.n564 10.6151
R940 B.n564 B.n9 10.6151
R941 B.n558 B.n9 10.6151
R942 B.n558 B.n557 10.6151
R943 B.n557 B.n556 10.6151
R944 B.n556 B.n16 10.6151
R945 B.n550 B.n16 10.6151
R946 B.n550 B.n549 10.6151
R947 B.n549 B.n548 10.6151
R948 B.n548 B.n23 10.6151
R949 B.n542 B.n23 10.6151
R950 B.n542 B.n541 10.6151
R951 B.n541 B.n540 10.6151
R952 B.n540 B.n29 10.6151
R953 B.n534 B.n29 10.6151
R954 B.n534 B.n533 10.6151
R955 B.n471 B.t7 10.2331
R956 B.t3 B.n552 10.2331
R957 B.n452 B.t11 8.65882
R958 B.n484 B.t6 8.65882
R959 B.n560 B.t0 8.65882
R960 B.n31 B.t18 8.65882
R961 B.n142 B.n80 6.5566
R962 B.n159 B.n158 6.5566
R963 B.n379 B.n378 6.5566
R964 B.n362 B.n296 6.5566
R965 B.n139 B.n80 4.05904
R966 B.n160 B.n159 4.05904
R967 B.n380 B.n379 4.05904
R968 B.n359 B.n296 4.05904
R969 B.n572 B.n0 2.81026
R970 B.n572 B.n1 2.81026
R971 B.n478 B.t4 0.78762
R972 B.n554 B.t1 0.78762
R973 VN.n9 VN.t9 866.09
R974 VN.n3 VN.t0 866.09
R975 VN.n20 VN.t2 866.09
R976 VN.n14 VN.t6 866.09
R977 VN.n6 VN.t8 831.034
R978 VN.n8 VN.t7 831.034
R979 VN.n2 VN.t5 831.034
R980 VN.n17 VN.t1 831.034
R981 VN.n19 VN.t4 831.034
R982 VN.n13 VN.t3 831.034
R983 VN.n15 VN.n14 161.489
R984 VN.n4 VN.n3 161.489
R985 VN.n10 VN.n9 161.3
R986 VN.n21 VN.n20 161.3
R987 VN.n18 VN.n11 161.3
R988 VN.n17 VN.n16 161.3
R989 VN.n15 VN.n12 161.3
R990 VN.n7 VN.n0 161.3
R991 VN.n6 VN.n5 161.3
R992 VN.n4 VN.n1 161.3
R993 VN.n6 VN.n1 73.0308
R994 VN.n7 VN.n6 73.0308
R995 VN.n18 VN.n17 73.0308
R996 VN.n17 VN.n12 73.0308
R997 VN.n3 VN.n2 55.5035
R998 VN.n9 VN.n8 55.5035
R999 VN.n20 VN.n19 55.5035
R1000 VN.n14 VN.n13 55.5035
R1001 VN VN.n21 38.4721
R1002 VN.n2 VN.n1 17.5278
R1003 VN.n8 VN.n7 17.5278
R1004 VN.n19 VN.n18 17.5278
R1005 VN.n13 VN.n12 17.5278
R1006 VN.n21 VN.n11 0.189894
R1007 VN.n16 VN.n11 0.189894
R1008 VN.n16 VN.n15 0.189894
R1009 VN.n5 VN.n4 0.189894
R1010 VN.n5 VN.n0 0.189894
R1011 VN.n10 VN.n0 0.189894
R1012 VN VN.n10 0.0516364
R1013 VTAIL.n192 VTAIL.n152 289.615
R1014 VTAIL.n42 VTAIL.n2 289.615
R1015 VTAIL.n146 VTAIL.n106 289.615
R1016 VTAIL.n96 VTAIL.n56 289.615
R1017 VTAIL.n167 VTAIL.n166 185
R1018 VTAIL.n164 VTAIL.n163 185
R1019 VTAIL.n173 VTAIL.n172 185
R1020 VTAIL.n175 VTAIL.n174 185
R1021 VTAIL.n160 VTAIL.n159 185
R1022 VTAIL.n181 VTAIL.n180 185
R1023 VTAIL.n184 VTAIL.n183 185
R1024 VTAIL.n182 VTAIL.n156 185
R1025 VTAIL.n189 VTAIL.n155 185
R1026 VTAIL.n191 VTAIL.n190 185
R1027 VTAIL.n193 VTAIL.n192 185
R1028 VTAIL.n17 VTAIL.n16 185
R1029 VTAIL.n14 VTAIL.n13 185
R1030 VTAIL.n23 VTAIL.n22 185
R1031 VTAIL.n25 VTAIL.n24 185
R1032 VTAIL.n10 VTAIL.n9 185
R1033 VTAIL.n31 VTAIL.n30 185
R1034 VTAIL.n34 VTAIL.n33 185
R1035 VTAIL.n32 VTAIL.n6 185
R1036 VTAIL.n39 VTAIL.n5 185
R1037 VTAIL.n41 VTAIL.n40 185
R1038 VTAIL.n43 VTAIL.n42 185
R1039 VTAIL.n147 VTAIL.n146 185
R1040 VTAIL.n145 VTAIL.n144 185
R1041 VTAIL.n143 VTAIL.n109 185
R1042 VTAIL.n113 VTAIL.n110 185
R1043 VTAIL.n138 VTAIL.n137 185
R1044 VTAIL.n136 VTAIL.n135 185
R1045 VTAIL.n115 VTAIL.n114 185
R1046 VTAIL.n130 VTAIL.n129 185
R1047 VTAIL.n128 VTAIL.n127 185
R1048 VTAIL.n119 VTAIL.n118 185
R1049 VTAIL.n122 VTAIL.n121 185
R1050 VTAIL.n97 VTAIL.n96 185
R1051 VTAIL.n95 VTAIL.n94 185
R1052 VTAIL.n93 VTAIL.n59 185
R1053 VTAIL.n63 VTAIL.n60 185
R1054 VTAIL.n88 VTAIL.n87 185
R1055 VTAIL.n86 VTAIL.n85 185
R1056 VTAIL.n65 VTAIL.n64 185
R1057 VTAIL.n80 VTAIL.n79 185
R1058 VTAIL.n78 VTAIL.n77 185
R1059 VTAIL.n69 VTAIL.n68 185
R1060 VTAIL.n72 VTAIL.n71 185
R1061 VTAIL.t8 VTAIL.n165 149.524
R1062 VTAIL.t3 VTAIL.n15 149.524
R1063 VTAIL.t5 VTAIL.n120 149.524
R1064 VTAIL.t14 VTAIL.n70 149.524
R1065 VTAIL.n166 VTAIL.n163 104.615
R1066 VTAIL.n173 VTAIL.n163 104.615
R1067 VTAIL.n174 VTAIL.n173 104.615
R1068 VTAIL.n174 VTAIL.n159 104.615
R1069 VTAIL.n181 VTAIL.n159 104.615
R1070 VTAIL.n183 VTAIL.n181 104.615
R1071 VTAIL.n183 VTAIL.n182 104.615
R1072 VTAIL.n182 VTAIL.n155 104.615
R1073 VTAIL.n191 VTAIL.n155 104.615
R1074 VTAIL.n192 VTAIL.n191 104.615
R1075 VTAIL.n16 VTAIL.n13 104.615
R1076 VTAIL.n23 VTAIL.n13 104.615
R1077 VTAIL.n24 VTAIL.n23 104.615
R1078 VTAIL.n24 VTAIL.n9 104.615
R1079 VTAIL.n31 VTAIL.n9 104.615
R1080 VTAIL.n33 VTAIL.n31 104.615
R1081 VTAIL.n33 VTAIL.n32 104.615
R1082 VTAIL.n32 VTAIL.n5 104.615
R1083 VTAIL.n41 VTAIL.n5 104.615
R1084 VTAIL.n42 VTAIL.n41 104.615
R1085 VTAIL.n146 VTAIL.n145 104.615
R1086 VTAIL.n145 VTAIL.n109 104.615
R1087 VTAIL.n113 VTAIL.n109 104.615
R1088 VTAIL.n137 VTAIL.n113 104.615
R1089 VTAIL.n137 VTAIL.n136 104.615
R1090 VTAIL.n136 VTAIL.n114 104.615
R1091 VTAIL.n129 VTAIL.n114 104.615
R1092 VTAIL.n129 VTAIL.n128 104.615
R1093 VTAIL.n128 VTAIL.n118 104.615
R1094 VTAIL.n121 VTAIL.n118 104.615
R1095 VTAIL.n96 VTAIL.n95 104.615
R1096 VTAIL.n95 VTAIL.n59 104.615
R1097 VTAIL.n63 VTAIL.n59 104.615
R1098 VTAIL.n87 VTAIL.n63 104.615
R1099 VTAIL.n87 VTAIL.n86 104.615
R1100 VTAIL.n86 VTAIL.n64 104.615
R1101 VTAIL.n79 VTAIL.n64 104.615
R1102 VTAIL.n79 VTAIL.n78 104.615
R1103 VTAIL.n78 VTAIL.n68 104.615
R1104 VTAIL.n71 VTAIL.n68 104.615
R1105 VTAIL.n166 VTAIL.t8 52.3082
R1106 VTAIL.n16 VTAIL.t3 52.3082
R1107 VTAIL.n121 VTAIL.t5 52.3082
R1108 VTAIL.n71 VTAIL.t14 52.3082
R1109 VTAIL.n105 VTAIL.n104 50.2533
R1110 VTAIL.n103 VTAIL.n102 50.2533
R1111 VTAIL.n55 VTAIL.n54 50.2533
R1112 VTAIL.n53 VTAIL.n52 50.2533
R1113 VTAIL.n199 VTAIL.n198 50.2531
R1114 VTAIL.n1 VTAIL.n0 50.2531
R1115 VTAIL.n49 VTAIL.n48 50.2531
R1116 VTAIL.n51 VTAIL.n50 50.2531
R1117 VTAIL.n197 VTAIL.n196 35.6763
R1118 VTAIL.n47 VTAIL.n46 35.6763
R1119 VTAIL.n151 VTAIL.n150 35.6763
R1120 VTAIL.n101 VTAIL.n100 35.6763
R1121 VTAIL.n53 VTAIL.n51 20.9358
R1122 VTAIL.n197 VTAIL.n151 20.4014
R1123 VTAIL.n190 VTAIL.n189 13.1884
R1124 VTAIL.n40 VTAIL.n39 13.1884
R1125 VTAIL.n144 VTAIL.n143 13.1884
R1126 VTAIL.n94 VTAIL.n93 13.1884
R1127 VTAIL.n188 VTAIL.n156 12.8005
R1128 VTAIL.n193 VTAIL.n154 12.8005
R1129 VTAIL.n38 VTAIL.n6 12.8005
R1130 VTAIL.n43 VTAIL.n4 12.8005
R1131 VTAIL.n147 VTAIL.n108 12.8005
R1132 VTAIL.n142 VTAIL.n110 12.8005
R1133 VTAIL.n97 VTAIL.n58 12.8005
R1134 VTAIL.n92 VTAIL.n60 12.8005
R1135 VTAIL.n185 VTAIL.n184 12.0247
R1136 VTAIL.n194 VTAIL.n152 12.0247
R1137 VTAIL.n35 VTAIL.n34 12.0247
R1138 VTAIL.n44 VTAIL.n2 12.0247
R1139 VTAIL.n148 VTAIL.n106 12.0247
R1140 VTAIL.n139 VTAIL.n138 12.0247
R1141 VTAIL.n98 VTAIL.n56 12.0247
R1142 VTAIL.n89 VTAIL.n88 12.0247
R1143 VTAIL.n180 VTAIL.n158 11.249
R1144 VTAIL.n30 VTAIL.n8 11.249
R1145 VTAIL.n135 VTAIL.n112 11.249
R1146 VTAIL.n85 VTAIL.n62 11.249
R1147 VTAIL.n179 VTAIL.n160 10.4732
R1148 VTAIL.n29 VTAIL.n10 10.4732
R1149 VTAIL.n134 VTAIL.n115 10.4732
R1150 VTAIL.n84 VTAIL.n65 10.4732
R1151 VTAIL.n167 VTAIL.n165 10.2747
R1152 VTAIL.n17 VTAIL.n15 10.2747
R1153 VTAIL.n122 VTAIL.n120 10.2747
R1154 VTAIL.n72 VTAIL.n70 10.2747
R1155 VTAIL.n176 VTAIL.n175 9.69747
R1156 VTAIL.n26 VTAIL.n25 9.69747
R1157 VTAIL.n131 VTAIL.n130 9.69747
R1158 VTAIL.n81 VTAIL.n80 9.69747
R1159 VTAIL.n196 VTAIL.n195 9.45567
R1160 VTAIL.n46 VTAIL.n45 9.45567
R1161 VTAIL.n150 VTAIL.n149 9.45567
R1162 VTAIL.n100 VTAIL.n99 9.45567
R1163 VTAIL.n195 VTAIL.n194 9.3005
R1164 VTAIL.n154 VTAIL.n153 9.3005
R1165 VTAIL.n169 VTAIL.n168 9.3005
R1166 VTAIL.n171 VTAIL.n170 9.3005
R1167 VTAIL.n162 VTAIL.n161 9.3005
R1168 VTAIL.n177 VTAIL.n176 9.3005
R1169 VTAIL.n179 VTAIL.n178 9.3005
R1170 VTAIL.n158 VTAIL.n157 9.3005
R1171 VTAIL.n186 VTAIL.n185 9.3005
R1172 VTAIL.n188 VTAIL.n187 9.3005
R1173 VTAIL.n45 VTAIL.n44 9.3005
R1174 VTAIL.n4 VTAIL.n3 9.3005
R1175 VTAIL.n19 VTAIL.n18 9.3005
R1176 VTAIL.n21 VTAIL.n20 9.3005
R1177 VTAIL.n12 VTAIL.n11 9.3005
R1178 VTAIL.n27 VTAIL.n26 9.3005
R1179 VTAIL.n29 VTAIL.n28 9.3005
R1180 VTAIL.n8 VTAIL.n7 9.3005
R1181 VTAIL.n36 VTAIL.n35 9.3005
R1182 VTAIL.n38 VTAIL.n37 9.3005
R1183 VTAIL.n124 VTAIL.n123 9.3005
R1184 VTAIL.n126 VTAIL.n125 9.3005
R1185 VTAIL.n117 VTAIL.n116 9.3005
R1186 VTAIL.n132 VTAIL.n131 9.3005
R1187 VTAIL.n134 VTAIL.n133 9.3005
R1188 VTAIL.n112 VTAIL.n111 9.3005
R1189 VTAIL.n140 VTAIL.n139 9.3005
R1190 VTAIL.n142 VTAIL.n141 9.3005
R1191 VTAIL.n149 VTAIL.n148 9.3005
R1192 VTAIL.n108 VTAIL.n107 9.3005
R1193 VTAIL.n74 VTAIL.n73 9.3005
R1194 VTAIL.n76 VTAIL.n75 9.3005
R1195 VTAIL.n67 VTAIL.n66 9.3005
R1196 VTAIL.n82 VTAIL.n81 9.3005
R1197 VTAIL.n84 VTAIL.n83 9.3005
R1198 VTAIL.n62 VTAIL.n61 9.3005
R1199 VTAIL.n90 VTAIL.n89 9.3005
R1200 VTAIL.n92 VTAIL.n91 9.3005
R1201 VTAIL.n99 VTAIL.n98 9.3005
R1202 VTAIL.n58 VTAIL.n57 9.3005
R1203 VTAIL.n172 VTAIL.n162 8.92171
R1204 VTAIL.n22 VTAIL.n12 8.92171
R1205 VTAIL.n127 VTAIL.n117 8.92171
R1206 VTAIL.n77 VTAIL.n67 8.92171
R1207 VTAIL.n171 VTAIL.n164 8.14595
R1208 VTAIL.n21 VTAIL.n14 8.14595
R1209 VTAIL.n126 VTAIL.n119 8.14595
R1210 VTAIL.n76 VTAIL.n69 8.14595
R1211 VTAIL.n168 VTAIL.n167 7.3702
R1212 VTAIL.n18 VTAIL.n17 7.3702
R1213 VTAIL.n123 VTAIL.n122 7.3702
R1214 VTAIL.n73 VTAIL.n72 7.3702
R1215 VTAIL.n168 VTAIL.n164 5.81868
R1216 VTAIL.n18 VTAIL.n14 5.81868
R1217 VTAIL.n123 VTAIL.n119 5.81868
R1218 VTAIL.n73 VTAIL.n69 5.81868
R1219 VTAIL.n172 VTAIL.n171 5.04292
R1220 VTAIL.n22 VTAIL.n21 5.04292
R1221 VTAIL.n127 VTAIL.n126 5.04292
R1222 VTAIL.n77 VTAIL.n76 5.04292
R1223 VTAIL.n175 VTAIL.n162 4.26717
R1224 VTAIL.n25 VTAIL.n12 4.26717
R1225 VTAIL.n130 VTAIL.n117 4.26717
R1226 VTAIL.n80 VTAIL.n67 4.26717
R1227 VTAIL.n176 VTAIL.n160 3.49141
R1228 VTAIL.n26 VTAIL.n10 3.49141
R1229 VTAIL.n131 VTAIL.n115 3.49141
R1230 VTAIL.n81 VTAIL.n65 3.49141
R1231 VTAIL.n169 VTAIL.n165 2.84303
R1232 VTAIL.n19 VTAIL.n15 2.84303
R1233 VTAIL.n124 VTAIL.n120 2.84303
R1234 VTAIL.n74 VTAIL.n70 2.84303
R1235 VTAIL.n180 VTAIL.n179 2.71565
R1236 VTAIL.n30 VTAIL.n29 2.71565
R1237 VTAIL.n135 VTAIL.n134 2.71565
R1238 VTAIL.n85 VTAIL.n84 2.71565
R1239 VTAIL.n198 VTAIL.t10 2.27636
R1240 VTAIL.n198 VTAIL.t7 2.27636
R1241 VTAIL.n0 VTAIL.t15 2.27636
R1242 VTAIL.n0 VTAIL.t13 2.27636
R1243 VTAIL.n48 VTAIL.t17 2.27636
R1244 VTAIL.n48 VTAIL.t19 2.27636
R1245 VTAIL.n50 VTAIL.t4 2.27636
R1246 VTAIL.n50 VTAIL.t6 2.27636
R1247 VTAIL.n104 VTAIL.t2 2.27636
R1248 VTAIL.n104 VTAIL.t1 2.27636
R1249 VTAIL.n102 VTAIL.t0 2.27636
R1250 VTAIL.n102 VTAIL.t18 2.27636
R1251 VTAIL.n54 VTAIL.t9 2.27636
R1252 VTAIL.n54 VTAIL.t11 2.27636
R1253 VTAIL.n52 VTAIL.t16 2.27636
R1254 VTAIL.n52 VTAIL.t12 2.27636
R1255 VTAIL.n184 VTAIL.n158 1.93989
R1256 VTAIL.n196 VTAIL.n152 1.93989
R1257 VTAIL.n34 VTAIL.n8 1.93989
R1258 VTAIL.n46 VTAIL.n2 1.93989
R1259 VTAIL.n150 VTAIL.n106 1.93989
R1260 VTAIL.n138 VTAIL.n112 1.93989
R1261 VTAIL.n100 VTAIL.n56 1.93989
R1262 VTAIL.n88 VTAIL.n62 1.93989
R1263 VTAIL.n185 VTAIL.n156 1.16414
R1264 VTAIL.n194 VTAIL.n193 1.16414
R1265 VTAIL.n35 VTAIL.n6 1.16414
R1266 VTAIL.n44 VTAIL.n43 1.16414
R1267 VTAIL.n148 VTAIL.n147 1.16414
R1268 VTAIL.n139 VTAIL.n110 1.16414
R1269 VTAIL.n98 VTAIL.n97 1.16414
R1270 VTAIL.n89 VTAIL.n60 1.16414
R1271 VTAIL.n103 VTAIL.n101 0.737569
R1272 VTAIL.n47 VTAIL.n1 0.737569
R1273 VTAIL.n55 VTAIL.n53 0.534983
R1274 VTAIL.n101 VTAIL.n55 0.534983
R1275 VTAIL.n105 VTAIL.n103 0.534983
R1276 VTAIL.n151 VTAIL.n105 0.534983
R1277 VTAIL.n51 VTAIL.n49 0.534983
R1278 VTAIL.n49 VTAIL.n47 0.534983
R1279 VTAIL.n199 VTAIL.n197 0.534983
R1280 VTAIL VTAIL.n1 0.459552
R1281 VTAIL.n189 VTAIL.n188 0.388379
R1282 VTAIL.n190 VTAIL.n154 0.388379
R1283 VTAIL.n39 VTAIL.n38 0.388379
R1284 VTAIL.n40 VTAIL.n4 0.388379
R1285 VTAIL.n144 VTAIL.n108 0.388379
R1286 VTAIL.n143 VTAIL.n142 0.388379
R1287 VTAIL.n94 VTAIL.n58 0.388379
R1288 VTAIL.n93 VTAIL.n92 0.388379
R1289 VTAIL.n170 VTAIL.n169 0.155672
R1290 VTAIL.n170 VTAIL.n161 0.155672
R1291 VTAIL.n177 VTAIL.n161 0.155672
R1292 VTAIL.n178 VTAIL.n177 0.155672
R1293 VTAIL.n178 VTAIL.n157 0.155672
R1294 VTAIL.n186 VTAIL.n157 0.155672
R1295 VTAIL.n187 VTAIL.n186 0.155672
R1296 VTAIL.n187 VTAIL.n153 0.155672
R1297 VTAIL.n195 VTAIL.n153 0.155672
R1298 VTAIL.n20 VTAIL.n19 0.155672
R1299 VTAIL.n20 VTAIL.n11 0.155672
R1300 VTAIL.n27 VTAIL.n11 0.155672
R1301 VTAIL.n28 VTAIL.n27 0.155672
R1302 VTAIL.n28 VTAIL.n7 0.155672
R1303 VTAIL.n36 VTAIL.n7 0.155672
R1304 VTAIL.n37 VTAIL.n36 0.155672
R1305 VTAIL.n37 VTAIL.n3 0.155672
R1306 VTAIL.n45 VTAIL.n3 0.155672
R1307 VTAIL.n149 VTAIL.n107 0.155672
R1308 VTAIL.n141 VTAIL.n107 0.155672
R1309 VTAIL.n141 VTAIL.n140 0.155672
R1310 VTAIL.n140 VTAIL.n111 0.155672
R1311 VTAIL.n133 VTAIL.n111 0.155672
R1312 VTAIL.n133 VTAIL.n132 0.155672
R1313 VTAIL.n132 VTAIL.n116 0.155672
R1314 VTAIL.n125 VTAIL.n116 0.155672
R1315 VTAIL.n125 VTAIL.n124 0.155672
R1316 VTAIL.n99 VTAIL.n57 0.155672
R1317 VTAIL.n91 VTAIL.n57 0.155672
R1318 VTAIL.n91 VTAIL.n90 0.155672
R1319 VTAIL.n90 VTAIL.n61 0.155672
R1320 VTAIL.n83 VTAIL.n61 0.155672
R1321 VTAIL.n83 VTAIL.n82 0.155672
R1322 VTAIL.n82 VTAIL.n66 0.155672
R1323 VTAIL.n75 VTAIL.n66 0.155672
R1324 VTAIL.n75 VTAIL.n74 0.155672
R1325 VTAIL VTAIL.n199 0.075931
R1326 VDD2.n89 VDD2.n49 289.615
R1327 VDD2.n40 VDD2.n0 289.615
R1328 VDD2.n90 VDD2.n89 185
R1329 VDD2.n88 VDD2.n87 185
R1330 VDD2.n86 VDD2.n52 185
R1331 VDD2.n56 VDD2.n53 185
R1332 VDD2.n81 VDD2.n80 185
R1333 VDD2.n79 VDD2.n78 185
R1334 VDD2.n58 VDD2.n57 185
R1335 VDD2.n73 VDD2.n72 185
R1336 VDD2.n71 VDD2.n70 185
R1337 VDD2.n62 VDD2.n61 185
R1338 VDD2.n65 VDD2.n64 185
R1339 VDD2.n15 VDD2.n14 185
R1340 VDD2.n12 VDD2.n11 185
R1341 VDD2.n21 VDD2.n20 185
R1342 VDD2.n23 VDD2.n22 185
R1343 VDD2.n8 VDD2.n7 185
R1344 VDD2.n29 VDD2.n28 185
R1345 VDD2.n32 VDD2.n31 185
R1346 VDD2.n30 VDD2.n4 185
R1347 VDD2.n37 VDD2.n3 185
R1348 VDD2.n39 VDD2.n38 185
R1349 VDD2.n41 VDD2.n40 185
R1350 VDD2.t7 VDD2.n63 149.524
R1351 VDD2.t9 VDD2.n13 149.524
R1352 VDD2.n89 VDD2.n88 104.615
R1353 VDD2.n88 VDD2.n52 104.615
R1354 VDD2.n56 VDD2.n52 104.615
R1355 VDD2.n80 VDD2.n56 104.615
R1356 VDD2.n80 VDD2.n79 104.615
R1357 VDD2.n79 VDD2.n57 104.615
R1358 VDD2.n72 VDD2.n57 104.615
R1359 VDD2.n72 VDD2.n71 104.615
R1360 VDD2.n71 VDD2.n61 104.615
R1361 VDD2.n64 VDD2.n61 104.615
R1362 VDD2.n14 VDD2.n11 104.615
R1363 VDD2.n21 VDD2.n11 104.615
R1364 VDD2.n22 VDD2.n21 104.615
R1365 VDD2.n22 VDD2.n7 104.615
R1366 VDD2.n29 VDD2.n7 104.615
R1367 VDD2.n31 VDD2.n29 104.615
R1368 VDD2.n31 VDD2.n30 104.615
R1369 VDD2.n30 VDD2.n3 104.615
R1370 VDD2.n39 VDD2.n3 104.615
R1371 VDD2.n40 VDD2.n39 104.615
R1372 VDD2.n48 VDD2.n47 67.2774
R1373 VDD2 VDD2.n97 67.2746
R1374 VDD2.n96 VDD2.n95 66.9321
R1375 VDD2.n46 VDD2.n45 66.9319
R1376 VDD2.n46 VDD2.n44 52.8895
R1377 VDD2.n94 VDD2.n93 52.355
R1378 VDD2.n64 VDD2.t7 52.3082
R1379 VDD2.n14 VDD2.t9 52.3082
R1380 VDD2.n94 VDD2.n48 33.7541
R1381 VDD2.n87 VDD2.n86 13.1884
R1382 VDD2.n38 VDD2.n37 13.1884
R1383 VDD2.n90 VDD2.n51 12.8005
R1384 VDD2.n85 VDD2.n53 12.8005
R1385 VDD2.n36 VDD2.n4 12.8005
R1386 VDD2.n41 VDD2.n2 12.8005
R1387 VDD2.n91 VDD2.n49 12.0247
R1388 VDD2.n82 VDD2.n81 12.0247
R1389 VDD2.n33 VDD2.n32 12.0247
R1390 VDD2.n42 VDD2.n0 12.0247
R1391 VDD2.n78 VDD2.n55 11.249
R1392 VDD2.n28 VDD2.n6 11.249
R1393 VDD2.n77 VDD2.n58 10.4732
R1394 VDD2.n27 VDD2.n8 10.4732
R1395 VDD2.n65 VDD2.n63 10.2747
R1396 VDD2.n15 VDD2.n13 10.2747
R1397 VDD2.n74 VDD2.n73 9.69747
R1398 VDD2.n24 VDD2.n23 9.69747
R1399 VDD2.n93 VDD2.n92 9.45567
R1400 VDD2.n44 VDD2.n43 9.45567
R1401 VDD2.n67 VDD2.n66 9.3005
R1402 VDD2.n69 VDD2.n68 9.3005
R1403 VDD2.n60 VDD2.n59 9.3005
R1404 VDD2.n75 VDD2.n74 9.3005
R1405 VDD2.n77 VDD2.n76 9.3005
R1406 VDD2.n55 VDD2.n54 9.3005
R1407 VDD2.n83 VDD2.n82 9.3005
R1408 VDD2.n85 VDD2.n84 9.3005
R1409 VDD2.n92 VDD2.n91 9.3005
R1410 VDD2.n51 VDD2.n50 9.3005
R1411 VDD2.n43 VDD2.n42 9.3005
R1412 VDD2.n2 VDD2.n1 9.3005
R1413 VDD2.n17 VDD2.n16 9.3005
R1414 VDD2.n19 VDD2.n18 9.3005
R1415 VDD2.n10 VDD2.n9 9.3005
R1416 VDD2.n25 VDD2.n24 9.3005
R1417 VDD2.n27 VDD2.n26 9.3005
R1418 VDD2.n6 VDD2.n5 9.3005
R1419 VDD2.n34 VDD2.n33 9.3005
R1420 VDD2.n36 VDD2.n35 9.3005
R1421 VDD2.n70 VDD2.n60 8.92171
R1422 VDD2.n20 VDD2.n10 8.92171
R1423 VDD2.n69 VDD2.n62 8.14595
R1424 VDD2.n19 VDD2.n12 8.14595
R1425 VDD2.n66 VDD2.n65 7.3702
R1426 VDD2.n16 VDD2.n15 7.3702
R1427 VDD2.n66 VDD2.n62 5.81868
R1428 VDD2.n16 VDD2.n12 5.81868
R1429 VDD2.n70 VDD2.n69 5.04292
R1430 VDD2.n20 VDD2.n19 5.04292
R1431 VDD2.n73 VDD2.n60 4.26717
R1432 VDD2.n23 VDD2.n10 4.26717
R1433 VDD2.n74 VDD2.n58 3.49141
R1434 VDD2.n24 VDD2.n8 3.49141
R1435 VDD2.n17 VDD2.n13 2.84303
R1436 VDD2.n67 VDD2.n63 2.84303
R1437 VDD2.n78 VDD2.n77 2.71565
R1438 VDD2.n28 VDD2.n27 2.71565
R1439 VDD2.n97 VDD2.t6 2.27636
R1440 VDD2.n97 VDD2.t3 2.27636
R1441 VDD2.n95 VDD2.t5 2.27636
R1442 VDD2.n95 VDD2.t8 2.27636
R1443 VDD2.n47 VDD2.t2 2.27636
R1444 VDD2.n47 VDD2.t0 2.27636
R1445 VDD2.n45 VDD2.t4 2.27636
R1446 VDD2.n45 VDD2.t1 2.27636
R1447 VDD2.n93 VDD2.n49 1.93989
R1448 VDD2.n81 VDD2.n55 1.93989
R1449 VDD2.n32 VDD2.n6 1.93989
R1450 VDD2.n44 VDD2.n0 1.93989
R1451 VDD2.n91 VDD2.n90 1.16414
R1452 VDD2.n82 VDD2.n53 1.16414
R1453 VDD2.n33 VDD2.n4 1.16414
R1454 VDD2.n42 VDD2.n41 1.16414
R1455 VDD2.n96 VDD2.n94 0.534983
R1456 VDD2.n87 VDD2.n51 0.388379
R1457 VDD2.n86 VDD2.n85 0.388379
R1458 VDD2.n37 VDD2.n36 0.388379
R1459 VDD2.n38 VDD2.n2 0.388379
R1460 VDD2 VDD2.n96 0.19231
R1461 VDD2.n92 VDD2.n50 0.155672
R1462 VDD2.n84 VDD2.n50 0.155672
R1463 VDD2.n84 VDD2.n83 0.155672
R1464 VDD2.n83 VDD2.n54 0.155672
R1465 VDD2.n76 VDD2.n54 0.155672
R1466 VDD2.n76 VDD2.n75 0.155672
R1467 VDD2.n75 VDD2.n59 0.155672
R1468 VDD2.n68 VDD2.n59 0.155672
R1469 VDD2.n68 VDD2.n67 0.155672
R1470 VDD2.n18 VDD2.n17 0.155672
R1471 VDD2.n18 VDD2.n9 0.155672
R1472 VDD2.n25 VDD2.n9 0.155672
R1473 VDD2.n26 VDD2.n25 0.155672
R1474 VDD2.n26 VDD2.n5 0.155672
R1475 VDD2.n34 VDD2.n5 0.155672
R1476 VDD2.n35 VDD2.n34 0.155672
R1477 VDD2.n35 VDD2.n1 0.155672
R1478 VDD2.n43 VDD2.n1 0.155672
R1479 VDD2.n48 VDD2.n46 0.0787747
R1480 VP.n21 VP.t3 866.09
R1481 VP.n14 VP.t4 866.09
R1482 VP.n5 VP.t5 866.09
R1483 VP.n11 VP.t1 866.09
R1484 VP.n18 VP.t7 831.034
R1485 VP.n20 VP.t9 831.034
R1486 VP.n13 VP.t0 831.034
R1487 VP.n8 VP.t6 831.034
R1488 VP.n4 VP.t8 831.034
R1489 VP.n10 VP.t2 831.034
R1490 VP.n6 VP.n5 161.489
R1491 VP.n22 VP.n21 161.3
R1492 VP.n6 VP.n3 161.3
R1493 VP.n8 VP.n7 161.3
R1494 VP.n9 VP.n2 161.3
R1495 VP.n12 VP.n11 161.3
R1496 VP.n19 VP.n0 161.3
R1497 VP.n18 VP.n17 161.3
R1498 VP.n16 VP.n1 161.3
R1499 VP.n15 VP.n14 161.3
R1500 VP.n18 VP.n1 73.0308
R1501 VP.n19 VP.n18 73.0308
R1502 VP.n8 VP.n3 73.0308
R1503 VP.n9 VP.n8 73.0308
R1504 VP.n14 VP.n13 55.5035
R1505 VP.n21 VP.n20 55.5035
R1506 VP.n5 VP.n4 55.5035
R1507 VP.n11 VP.n10 55.5035
R1508 VP.n15 VP.n12 38.0914
R1509 VP.n13 VP.n1 17.5278
R1510 VP.n20 VP.n19 17.5278
R1511 VP.n4 VP.n3 17.5278
R1512 VP.n10 VP.n9 17.5278
R1513 VP.n7 VP.n6 0.189894
R1514 VP.n7 VP.n2 0.189894
R1515 VP.n12 VP.n2 0.189894
R1516 VP.n16 VP.n15 0.189894
R1517 VP.n17 VP.n16 0.189894
R1518 VP.n17 VP.n0 0.189894
R1519 VP.n22 VP.n0 0.189894
R1520 VP VP.n22 0.0516364
R1521 VDD1.n40 VDD1.n0 289.615
R1522 VDD1.n87 VDD1.n47 289.615
R1523 VDD1.n41 VDD1.n40 185
R1524 VDD1.n39 VDD1.n38 185
R1525 VDD1.n37 VDD1.n3 185
R1526 VDD1.n7 VDD1.n4 185
R1527 VDD1.n32 VDD1.n31 185
R1528 VDD1.n30 VDD1.n29 185
R1529 VDD1.n9 VDD1.n8 185
R1530 VDD1.n24 VDD1.n23 185
R1531 VDD1.n22 VDD1.n21 185
R1532 VDD1.n13 VDD1.n12 185
R1533 VDD1.n16 VDD1.n15 185
R1534 VDD1.n62 VDD1.n61 185
R1535 VDD1.n59 VDD1.n58 185
R1536 VDD1.n68 VDD1.n67 185
R1537 VDD1.n70 VDD1.n69 185
R1538 VDD1.n55 VDD1.n54 185
R1539 VDD1.n76 VDD1.n75 185
R1540 VDD1.n79 VDD1.n78 185
R1541 VDD1.n77 VDD1.n51 185
R1542 VDD1.n84 VDD1.n50 185
R1543 VDD1.n86 VDD1.n85 185
R1544 VDD1.n88 VDD1.n87 185
R1545 VDD1.t4 VDD1.n14 149.524
R1546 VDD1.t5 VDD1.n60 149.524
R1547 VDD1.n40 VDD1.n39 104.615
R1548 VDD1.n39 VDD1.n3 104.615
R1549 VDD1.n7 VDD1.n3 104.615
R1550 VDD1.n31 VDD1.n7 104.615
R1551 VDD1.n31 VDD1.n30 104.615
R1552 VDD1.n30 VDD1.n8 104.615
R1553 VDD1.n23 VDD1.n8 104.615
R1554 VDD1.n23 VDD1.n22 104.615
R1555 VDD1.n22 VDD1.n12 104.615
R1556 VDD1.n15 VDD1.n12 104.615
R1557 VDD1.n61 VDD1.n58 104.615
R1558 VDD1.n68 VDD1.n58 104.615
R1559 VDD1.n69 VDD1.n68 104.615
R1560 VDD1.n69 VDD1.n54 104.615
R1561 VDD1.n76 VDD1.n54 104.615
R1562 VDD1.n78 VDD1.n76 104.615
R1563 VDD1.n78 VDD1.n77 104.615
R1564 VDD1.n77 VDD1.n50 104.615
R1565 VDD1.n86 VDD1.n50 104.615
R1566 VDD1.n87 VDD1.n86 104.615
R1567 VDD1.n95 VDD1.n94 67.2774
R1568 VDD1.n46 VDD1.n45 66.9321
R1569 VDD1.n97 VDD1.n96 66.9319
R1570 VDD1.n93 VDD1.n92 66.9319
R1571 VDD1.n46 VDD1.n44 52.8895
R1572 VDD1.n93 VDD1.n91 52.8895
R1573 VDD1.n15 VDD1.t4 52.3082
R1574 VDD1.n61 VDD1.t5 52.3082
R1575 VDD1.n97 VDD1.n95 34.6043
R1576 VDD1.n38 VDD1.n37 13.1884
R1577 VDD1.n85 VDD1.n84 13.1884
R1578 VDD1.n41 VDD1.n2 12.8005
R1579 VDD1.n36 VDD1.n4 12.8005
R1580 VDD1.n83 VDD1.n51 12.8005
R1581 VDD1.n88 VDD1.n49 12.8005
R1582 VDD1.n42 VDD1.n0 12.0247
R1583 VDD1.n33 VDD1.n32 12.0247
R1584 VDD1.n80 VDD1.n79 12.0247
R1585 VDD1.n89 VDD1.n47 12.0247
R1586 VDD1.n29 VDD1.n6 11.249
R1587 VDD1.n75 VDD1.n53 11.249
R1588 VDD1.n28 VDD1.n9 10.4732
R1589 VDD1.n74 VDD1.n55 10.4732
R1590 VDD1.n16 VDD1.n14 10.2747
R1591 VDD1.n62 VDD1.n60 10.2747
R1592 VDD1.n25 VDD1.n24 9.69747
R1593 VDD1.n71 VDD1.n70 9.69747
R1594 VDD1.n44 VDD1.n43 9.45567
R1595 VDD1.n91 VDD1.n90 9.45567
R1596 VDD1.n18 VDD1.n17 9.3005
R1597 VDD1.n20 VDD1.n19 9.3005
R1598 VDD1.n11 VDD1.n10 9.3005
R1599 VDD1.n26 VDD1.n25 9.3005
R1600 VDD1.n28 VDD1.n27 9.3005
R1601 VDD1.n6 VDD1.n5 9.3005
R1602 VDD1.n34 VDD1.n33 9.3005
R1603 VDD1.n36 VDD1.n35 9.3005
R1604 VDD1.n43 VDD1.n42 9.3005
R1605 VDD1.n2 VDD1.n1 9.3005
R1606 VDD1.n90 VDD1.n89 9.3005
R1607 VDD1.n49 VDD1.n48 9.3005
R1608 VDD1.n64 VDD1.n63 9.3005
R1609 VDD1.n66 VDD1.n65 9.3005
R1610 VDD1.n57 VDD1.n56 9.3005
R1611 VDD1.n72 VDD1.n71 9.3005
R1612 VDD1.n74 VDD1.n73 9.3005
R1613 VDD1.n53 VDD1.n52 9.3005
R1614 VDD1.n81 VDD1.n80 9.3005
R1615 VDD1.n83 VDD1.n82 9.3005
R1616 VDD1.n21 VDD1.n11 8.92171
R1617 VDD1.n67 VDD1.n57 8.92171
R1618 VDD1.n20 VDD1.n13 8.14595
R1619 VDD1.n66 VDD1.n59 8.14595
R1620 VDD1.n17 VDD1.n16 7.3702
R1621 VDD1.n63 VDD1.n62 7.3702
R1622 VDD1.n17 VDD1.n13 5.81868
R1623 VDD1.n63 VDD1.n59 5.81868
R1624 VDD1.n21 VDD1.n20 5.04292
R1625 VDD1.n67 VDD1.n66 5.04292
R1626 VDD1.n24 VDD1.n11 4.26717
R1627 VDD1.n70 VDD1.n57 4.26717
R1628 VDD1.n25 VDD1.n9 3.49141
R1629 VDD1.n71 VDD1.n55 3.49141
R1630 VDD1.n64 VDD1.n60 2.84303
R1631 VDD1.n18 VDD1.n14 2.84303
R1632 VDD1.n29 VDD1.n28 2.71565
R1633 VDD1.n75 VDD1.n74 2.71565
R1634 VDD1.n96 VDD1.t7 2.27636
R1635 VDD1.n96 VDD1.t8 2.27636
R1636 VDD1.n45 VDD1.t1 2.27636
R1637 VDD1.n45 VDD1.t3 2.27636
R1638 VDD1.n94 VDD1.t0 2.27636
R1639 VDD1.n94 VDD1.t6 2.27636
R1640 VDD1.n92 VDD1.t9 2.27636
R1641 VDD1.n92 VDD1.t2 2.27636
R1642 VDD1.n44 VDD1.n0 1.93989
R1643 VDD1.n32 VDD1.n6 1.93989
R1644 VDD1.n79 VDD1.n53 1.93989
R1645 VDD1.n91 VDD1.n47 1.93989
R1646 VDD1.n42 VDD1.n41 1.16414
R1647 VDD1.n33 VDD1.n4 1.16414
R1648 VDD1.n80 VDD1.n51 1.16414
R1649 VDD1.n89 VDD1.n88 1.16414
R1650 VDD1.n38 VDD1.n2 0.388379
R1651 VDD1.n37 VDD1.n36 0.388379
R1652 VDD1.n84 VDD1.n83 0.388379
R1653 VDD1.n85 VDD1.n49 0.388379
R1654 VDD1 VDD1.n97 0.343172
R1655 VDD1 VDD1.n46 0.19231
R1656 VDD1.n43 VDD1.n1 0.155672
R1657 VDD1.n35 VDD1.n1 0.155672
R1658 VDD1.n35 VDD1.n34 0.155672
R1659 VDD1.n34 VDD1.n5 0.155672
R1660 VDD1.n27 VDD1.n5 0.155672
R1661 VDD1.n27 VDD1.n26 0.155672
R1662 VDD1.n26 VDD1.n10 0.155672
R1663 VDD1.n19 VDD1.n10 0.155672
R1664 VDD1.n19 VDD1.n18 0.155672
R1665 VDD1.n65 VDD1.n64 0.155672
R1666 VDD1.n65 VDD1.n56 0.155672
R1667 VDD1.n72 VDD1.n56 0.155672
R1668 VDD1.n73 VDD1.n72 0.155672
R1669 VDD1.n73 VDD1.n52 0.155672
R1670 VDD1.n81 VDD1.n52 0.155672
R1671 VDD1.n82 VDD1.n81 0.155672
R1672 VDD1.n82 VDD1.n48 0.155672
R1673 VDD1.n90 VDD1.n48 0.155672
R1674 VDD1.n95 VDD1.n93 0.0787747
C0 VDD2 VTAIL 15.9854f
C1 VDD2 VP 0.289192f
C2 VP VTAIL 2.68141f
C3 VDD1 VN 0.148358f
C4 VDD1 VDD2 0.718589f
C5 VDD2 VN 2.92739f
C6 VDD1 VTAIL 15.9534f
C7 VN VTAIL 2.66683f
C8 VDD1 VP 3.0644f
C9 VP VN 4.38034f
C10 VDD2 B 3.932622f
C11 VDD1 B 3.797672f
C12 VTAIL B 4.902755f
C13 VN B 7.3094f
C14 VP B 5.300401f
C15 VDD1.n0 B 0.041888f
C16 VDD1.n1 B 0.03009f
C17 VDD1.n2 B 0.016169f
C18 VDD1.n3 B 0.038218f
C19 VDD1.n4 B 0.01712f
C20 VDD1.n5 B 0.03009f
C21 VDD1.n6 B 0.016169f
C22 VDD1.n7 B 0.038218f
C23 VDD1.n8 B 0.038218f
C24 VDD1.n9 B 0.01712f
C25 VDD1.n10 B 0.03009f
C26 VDD1.n11 B 0.016169f
C27 VDD1.n12 B 0.038218f
C28 VDD1.n13 B 0.01712f
C29 VDD1.n14 B 0.178846f
C30 VDD1.t4 B 0.064025f
C31 VDD1.n15 B 0.028664f
C32 VDD1.n16 B 0.027017f
C33 VDD1.n17 B 0.016169f
C34 VDD1.n18 B 1.07631f
C35 VDD1.n19 B 0.03009f
C36 VDD1.n20 B 0.016169f
C37 VDD1.n21 B 0.01712f
C38 VDD1.n22 B 0.038218f
C39 VDD1.n23 B 0.038218f
C40 VDD1.n24 B 0.01712f
C41 VDD1.n25 B 0.016169f
C42 VDD1.n26 B 0.03009f
C43 VDD1.n27 B 0.03009f
C44 VDD1.n28 B 0.016169f
C45 VDD1.n29 B 0.01712f
C46 VDD1.n30 B 0.038218f
C47 VDD1.n31 B 0.038218f
C48 VDD1.n32 B 0.01712f
C49 VDD1.n33 B 0.016169f
C50 VDD1.n34 B 0.03009f
C51 VDD1.n35 B 0.03009f
C52 VDD1.n36 B 0.016169f
C53 VDD1.n37 B 0.016645f
C54 VDD1.n38 B 0.016645f
C55 VDD1.n39 B 0.038218f
C56 VDD1.n40 B 0.082018f
C57 VDD1.n41 B 0.01712f
C58 VDD1.n42 B 0.016169f
C59 VDD1.n43 B 0.076951f
C60 VDD1.n44 B 0.067913f
C61 VDD1.t1 B 0.206871f
C62 VDD1.t3 B 0.206871f
C63 VDD1.n45 B 1.80546f
C64 VDD1.n46 B 0.42278f
C65 VDD1.n47 B 0.041888f
C66 VDD1.n48 B 0.03009f
C67 VDD1.n49 B 0.016169f
C68 VDD1.n50 B 0.038218f
C69 VDD1.n51 B 0.01712f
C70 VDD1.n52 B 0.03009f
C71 VDD1.n53 B 0.016169f
C72 VDD1.n54 B 0.038218f
C73 VDD1.n55 B 0.01712f
C74 VDD1.n56 B 0.03009f
C75 VDD1.n57 B 0.016169f
C76 VDD1.n58 B 0.038218f
C77 VDD1.n59 B 0.01712f
C78 VDD1.n60 B 0.178846f
C79 VDD1.t5 B 0.064025f
C80 VDD1.n61 B 0.028664f
C81 VDD1.n62 B 0.027017f
C82 VDD1.n63 B 0.016169f
C83 VDD1.n64 B 1.07631f
C84 VDD1.n65 B 0.03009f
C85 VDD1.n66 B 0.016169f
C86 VDD1.n67 B 0.01712f
C87 VDD1.n68 B 0.038218f
C88 VDD1.n69 B 0.038218f
C89 VDD1.n70 B 0.01712f
C90 VDD1.n71 B 0.016169f
C91 VDD1.n72 B 0.03009f
C92 VDD1.n73 B 0.03009f
C93 VDD1.n74 B 0.016169f
C94 VDD1.n75 B 0.01712f
C95 VDD1.n76 B 0.038218f
C96 VDD1.n77 B 0.038218f
C97 VDD1.n78 B 0.038218f
C98 VDD1.n79 B 0.01712f
C99 VDD1.n80 B 0.016169f
C100 VDD1.n81 B 0.03009f
C101 VDD1.n82 B 0.03009f
C102 VDD1.n83 B 0.016169f
C103 VDD1.n84 B 0.016645f
C104 VDD1.n85 B 0.016645f
C105 VDD1.n86 B 0.038218f
C106 VDD1.n87 B 0.082018f
C107 VDD1.n88 B 0.01712f
C108 VDD1.n89 B 0.016169f
C109 VDD1.n90 B 0.076951f
C110 VDD1.n91 B 0.067913f
C111 VDD1.t9 B 0.206871f
C112 VDD1.t2 B 0.206871f
C113 VDD1.n92 B 1.80545f
C114 VDD1.n93 B 0.420691f
C115 VDD1.t0 B 0.206871f
C116 VDD1.t6 B 0.206871f
C117 VDD1.n94 B 1.80719f
C118 VDD1.n95 B 1.85824f
C119 VDD1.t7 B 0.206871f
C120 VDD1.t8 B 0.206871f
C121 VDD1.n96 B 1.80545f
C122 VDD1.n97 B 2.34743f
C123 VP.n0 B 0.055226f
C124 VP.t9 B 0.394974f
C125 VP.t7 B 0.394974f
C126 VP.n1 B 0.022406f
C127 VP.n2 B 0.055226f
C128 VP.t2 B 0.394974f
C129 VP.t6 B 0.394974f
C130 VP.n3 B 0.022406f
C131 VP.t5 B 0.40176f
C132 VP.t8 B 0.394974f
C133 VP.n4 B 0.166636f
C134 VP.n5 B 0.183354f
C135 VP.n6 B 0.119571f
C136 VP.n7 B 0.055226f
C137 VP.n8 B 0.184956f
C138 VP.n9 B 0.022406f
C139 VP.n10 B 0.166636f
C140 VP.t1 B 0.40176f
C141 VP.n11 B 0.183278f
C142 VP.n12 B 1.92573f
C143 VP.t4 B 0.40176f
C144 VP.t0 B 0.394974f
C145 VP.n13 B 0.166636f
C146 VP.n14 B 0.183278f
C147 VP.n15 B 1.978f
C148 VP.n16 B 0.055226f
C149 VP.n17 B 0.055226f
C150 VP.n18 B 0.184956f
C151 VP.n19 B 0.022406f
C152 VP.n20 B 0.166636f
C153 VP.t3 B 0.40176f
C154 VP.n21 B 0.183278f
C155 VP.n22 B 0.042798f
C156 VDD2.n0 B 0.041692f
C157 VDD2.n1 B 0.029949f
C158 VDD2.n2 B 0.016093f
C159 VDD2.n3 B 0.038039f
C160 VDD2.n4 B 0.01704f
C161 VDD2.n5 B 0.029949f
C162 VDD2.n6 B 0.016093f
C163 VDD2.n7 B 0.038039f
C164 VDD2.n8 B 0.01704f
C165 VDD2.n9 B 0.029949f
C166 VDD2.n10 B 0.016093f
C167 VDD2.n11 B 0.038039f
C168 VDD2.n12 B 0.01704f
C169 VDD2.n13 B 0.178009f
C170 VDD2.t9 B 0.063725f
C171 VDD2.n14 B 0.028529f
C172 VDD2.n15 B 0.026891f
C173 VDD2.n16 B 0.016093f
C174 VDD2.n17 B 1.07127f
C175 VDD2.n18 B 0.029949f
C176 VDD2.n19 B 0.016093f
C177 VDD2.n20 B 0.01704f
C178 VDD2.n21 B 0.038039f
C179 VDD2.n22 B 0.038039f
C180 VDD2.n23 B 0.01704f
C181 VDD2.n24 B 0.016093f
C182 VDD2.n25 B 0.029949f
C183 VDD2.n26 B 0.029949f
C184 VDD2.n27 B 0.016093f
C185 VDD2.n28 B 0.01704f
C186 VDD2.n29 B 0.038039f
C187 VDD2.n30 B 0.038039f
C188 VDD2.n31 B 0.038039f
C189 VDD2.n32 B 0.01704f
C190 VDD2.n33 B 0.016093f
C191 VDD2.n34 B 0.029949f
C192 VDD2.n35 B 0.029949f
C193 VDD2.n36 B 0.016093f
C194 VDD2.n37 B 0.016567f
C195 VDD2.n38 B 0.016567f
C196 VDD2.n39 B 0.038039f
C197 VDD2.n40 B 0.081634f
C198 VDD2.n41 B 0.01704f
C199 VDD2.n42 B 0.016093f
C200 VDD2.n43 B 0.076591f
C201 VDD2.n44 B 0.067595f
C202 VDD2.t4 B 0.205903f
C203 VDD2.t1 B 0.205903f
C204 VDD2.n45 B 1.797f
C205 VDD2.n46 B 0.418722f
C206 VDD2.t2 B 0.205903f
C207 VDD2.t0 B 0.205903f
C208 VDD2.n47 B 1.79874f
C209 VDD2.n48 B 1.76943f
C210 VDD2.n49 B 0.041692f
C211 VDD2.n50 B 0.029949f
C212 VDD2.n51 B 0.016093f
C213 VDD2.n52 B 0.038039f
C214 VDD2.n53 B 0.01704f
C215 VDD2.n54 B 0.029949f
C216 VDD2.n55 B 0.016093f
C217 VDD2.n56 B 0.038039f
C218 VDD2.n57 B 0.038039f
C219 VDD2.n58 B 0.01704f
C220 VDD2.n59 B 0.029949f
C221 VDD2.n60 B 0.016093f
C222 VDD2.n61 B 0.038039f
C223 VDD2.n62 B 0.01704f
C224 VDD2.n63 B 0.178009f
C225 VDD2.t7 B 0.063725f
C226 VDD2.n64 B 0.028529f
C227 VDD2.n65 B 0.026891f
C228 VDD2.n66 B 0.016093f
C229 VDD2.n67 B 1.07127f
C230 VDD2.n68 B 0.029949f
C231 VDD2.n69 B 0.016093f
C232 VDD2.n70 B 0.01704f
C233 VDD2.n71 B 0.038039f
C234 VDD2.n72 B 0.038039f
C235 VDD2.n73 B 0.01704f
C236 VDD2.n74 B 0.016093f
C237 VDD2.n75 B 0.029949f
C238 VDD2.n76 B 0.029949f
C239 VDD2.n77 B 0.016093f
C240 VDD2.n78 B 0.01704f
C241 VDD2.n79 B 0.038039f
C242 VDD2.n80 B 0.038039f
C243 VDD2.n81 B 0.01704f
C244 VDD2.n82 B 0.016093f
C245 VDD2.n83 B 0.029949f
C246 VDD2.n84 B 0.029949f
C247 VDD2.n85 B 0.016093f
C248 VDD2.n86 B 0.016567f
C249 VDD2.n87 B 0.016567f
C250 VDD2.n88 B 0.038039f
C251 VDD2.n89 B 0.081634f
C252 VDD2.n90 B 0.01704f
C253 VDD2.n91 B 0.016093f
C254 VDD2.n92 B 0.076591f
C255 VDD2.n93 B 0.066448f
C256 VDD2.n94 B 2.0843f
C257 VDD2.t5 B 0.205903f
C258 VDD2.t8 B 0.205903f
C259 VDD2.n95 B 1.79701f
C260 VDD2.n96 B 0.30848f
C261 VDD2.t6 B 0.205903f
C262 VDD2.t3 B 0.205903f
C263 VDD2.n97 B 1.79871f
C264 VTAIL.t15 B 0.217421f
C265 VTAIL.t13 B 0.217421f
C266 VTAIL.n0 B 1.81598f
C267 VTAIL.n1 B 0.412188f
C268 VTAIL.n2 B 0.044025f
C269 VTAIL.n3 B 0.031625f
C270 VTAIL.n4 B 0.016994f
C271 VTAIL.n5 B 0.040167f
C272 VTAIL.n6 B 0.017993f
C273 VTAIL.n7 B 0.031625f
C274 VTAIL.n8 B 0.016994f
C275 VTAIL.n9 B 0.040167f
C276 VTAIL.n10 B 0.017993f
C277 VTAIL.n11 B 0.031625f
C278 VTAIL.n12 B 0.016994f
C279 VTAIL.n13 B 0.040167f
C280 VTAIL.n14 B 0.017993f
C281 VTAIL.n15 B 0.187967f
C282 VTAIL.t3 B 0.06729f
C283 VTAIL.n16 B 0.030125f
C284 VTAIL.n17 B 0.028395f
C285 VTAIL.n18 B 0.016994f
C286 VTAIL.n19 B 1.1312f
C287 VTAIL.n20 B 0.031625f
C288 VTAIL.n21 B 0.016994f
C289 VTAIL.n22 B 0.017993f
C290 VTAIL.n23 B 0.040167f
C291 VTAIL.n24 B 0.040167f
C292 VTAIL.n25 B 0.017993f
C293 VTAIL.n26 B 0.016994f
C294 VTAIL.n27 B 0.031625f
C295 VTAIL.n28 B 0.031625f
C296 VTAIL.n29 B 0.016994f
C297 VTAIL.n30 B 0.017993f
C298 VTAIL.n31 B 0.040167f
C299 VTAIL.n32 B 0.040167f
C300 VTAIL.n33 B 0.040167f
C301 VTAIL.n34 B 0.017993f
C302 VTAIL.n35 B 0.016994f
C303 VTAIL.n36 B 0.031625f
C304 VTAIL.n37 B 0.031625f
C305 VTAIL.n38 B 0.016994f
C306 VTAIL.n39 B 0.017494f
C307 VTAIL.n40 B 0.017494f
C308 VTAIL.n41 B 0.040167f
C309 VTAIL.n42 B 0.0862f
C310 VTAIL.n43 B 0.017993f
C311 VTAIL.n44 B 0.016994f
C312 VTAIL.n45 B 0.080876f
C313 VTAIL.n46 B 0.048383f
C314 VTAIL.n47 B 0.160984f
C315 VTAIL.t17 B 0.217421f
C316 VTAIL.t19 B 0.217421f
C317 VTAIL.n48 B 1.81598f
C318 VTAIL.n49 B 0.399231f
C319 VTAIL.t4 B 0.217421f
C320 VTAIL.t6 B 0.217421f
C321 VTAIL.n50 B 1.81598f
C322 VTAIL.n51 B 1.64755f
C323 VTAIL.t16 B 0.217421f
C324 VTAIL.t12 B 0.217421f
C325 VTAIL.n52 B 1.81599f
C326 VTAIL.n53 B 1.64754f
C327 VTAIL.t9 B 0.217421f
C328 VTAIL.t11 B 0.217421f
C329 VTAIL.n54 B 1.81599f
C330 VTAIL.n55 B 0.39922f
C331 VTAIL.n56 B 0.044025f
C332 VTAIL.n57 B 0.031625f
C333 VTAIL.n58 B 0.016994f
C334 VTAIL.n59 B 0.040167f
C335 VTAIL.n60 B 0.017993f
C336 VTAIL.n61 B 0.031625f
C337 VTAIL.n62 B 0.016994f
C338 VTAIL.n63 B 0.040167f
C339 VTAIL.n64 B 0.040167f
C340 VTAIL.n65 B 0.017993f
C341 VTAIL.n66 B 0.031625f
C342 VTAIL.n67 B 0.016994f
C343 VTAIL.n68 B 0.040167f
C344 VTAIL.n69 B 0.017993f
C345 VTAIL.n70 B 0.187967f
C346 VTAIL.t14 B 0.06729f
C347 VTAIL.n71 B 0.030125f
C348 VTAIL.n72 B 0.028395f
C349 VTAIL.n73 B 0.016994f
C350 VTAIL.n74 B 1.1312f
C351 VTAIL.n75 B 0.031625f
C352 VTAIL.n76 B 0.016994f
C353 VTAIL.n77 B 0.017993f
C354 VTAIL.n78 B 0.040167f
C355 VTAIL.n79 B 0.040167f
C356 VTAIL.n80 B 0.017993f
C357 VTAIL.n81 B 0.016994f
C358 VTAIL.n82 B 0.031625f
C359 VTAIL.n83 B 0.031625f
C360 VTAIL.n84 B 0.016994f
C361 VTAIL.n85 B 0.017993f
C362 VTAIL.n86 B 0.040167f
C363 VTAIL.n87 B 0.040167f
C364 VTAIL.n88 B 0.017993f
C365 VTAIL.n89 B 0.016994f
C366 VTAIL.n90 B 0.031625f
C367 VTAIL.n91 B 0.031625f
C368 VTAIL.n92 B 0.016994f
C369 VTAIL.n93 B 0.017494f
C370 VTAIL.n94 B 0.017494f
C371 VTAIL.n95 B 0.040167f
C372 VTAIL.n96 B 0.0862f
C373 VTAIL.n97 B 0.017993f
C374 VTAIL.n98 B 0.016994f
C375 VTAIL.n99 B 0.080876f
C376 VTAIL.n100 B 0.048383f
C377 VTAIL.n101 B 0.160984f
C378 VTAIL.t0 B 0.217421f
C379 VTAIL.t18 B 0.217421f
C380 VTAIL.n102 B 1.81599f
C381 VTAIL.n103 B 0.419864f
C382 VTAIL.t2 B 0.217421f
C383 VTAIL.t1 B 0.217421f
C384 VTAIL.n104 B 1.81599f
C385 VTAIL.n105 B 0.39922f
C386 VTAIL.n106 B 0.044025f
C387 VTAIL.n107 B 0.031625f
C388 VTAIL.n108 B 0.016994f
C389 VTAIL.n109 B 0.040167f
C390 VTAIL.n110 B 0.017993f
C391 VTAIL.n111 B 0.031625f
C392 VTAIL.n112 B 0.016994f
C393 VTAIL.n113 B 0.040167f
C394 VTAIL.n114 B 0.040167f
C395 VTAIL.n115 B 0.017993f
C396 VTAIL.n116 B 0.031625f
C397 VTAIL.n117 B 0.016994f
C398 VTAIL.n118 B 0.040167f
C399 VTAIL.n119 B 0.017993f
C400 VTAIL.n120 B 0.187967f
C401 VTAIL.t5 B 0.06729f
C402 VTAIL.n121 B 0.030125f
C403 VTAIL.n122 B 0.028395f
C404 VTAIL.n123 B 0.016994f
C405 VTAIL.n124 B 1.1312f
C406 VTAIL.n125 B 0.031625f
C407 VTAIL.n126 B 0.016994f
C408 VTAIL.n127 B 0.017993f
C409 VTAIL.n128 B 0.040167f
C410 VTAIL.n129 B 0.040167f
C411 VTAIL.n130 B 0.017993f
C412 VTAIL.n131 B 0.016994f
C413 VTAIL.n132 B 0.031625f
C414 VTAIL.n133 B 0.031625f
C415 VTAIL.n134 B 0.016994f
C416 VTAIL.n135 B 0.017993f
C417 VTAIL.n136 B 0.040167f
C418 VTAIL.n137 B 0.040167f
C419 VTAIL.n138 B 0.017993f
C420 VTAIL.n139 B 0.016994f
C421 VTAIL.n140 B 0.031625f
C422 VTAIL.n141 B 0.031625f
C423 VTAIL.n142 B 0.016994f
C424 VTAIL.n143 B 0.017494f
C425 VTAIL.n144 B 0.017494f
C426 VTAIL.n145 B 0.040167f
C427 VTAIL.n146 B 0.0862f
C428 VTAIL.n147 B 0.017993f
C429 VTAIL.n148 B 0.016994f
C430 VTAIL.n149 B 0.080876f
C431 VTAIL.n150 B 0.048383f
C432 VTAIL.n151 B 1.33419f
C433 VTAIL.n152 B 0.044025f
C434 VTAIL.n153 B 0.031625f
C435 VTAIL.n154 B 0.016994f
C436 VTAIL.n155 B 0.040167f
C437 VTAIL.n156 B 0.017993f
C438 VTAIL.n157 B 0.031625f
C439 VTAIL.n158 B 0.016994f
C440 VTAIL.n159 B 0.040167f
C441 VTAIL.n160 B 0.017993f
C442 VTAIL.n161 B 0.031625f
C443 VTAIL.n162 B 0.016994f
C444 VTAIL.n163 B 0.040167f
C445 VTAIL.n164 B 0.017993f
C446 VTAIL.n165 B 0.187967f
C447 VTAIL.t8 B 0.06729f
C448 VTAIL.n166 B 0.030125f
C449 VTAIL.n167 B 0.028395f
C450 VTAIL.n168 B 0.016994f
C451 VTAIL.n169 B 1.1312f
C452 VTAIL.n170 B 0.031625f
C453 VTAIL.n171 B 0.016994f
C454 VTAIL.n172 B 0.017993f
C455 VTAIL.n173 B 0.040167f
C456 VTAIL.n174 B 0.040167f
C457 VTAIL.n175 B 0.017993f
C458 VTAIL.n176 B 0.016994f
C459 VTAIL.n177 B 0.031625f
C460 VTAIL.n178 B 0.031625f
C461 VTAIL.n179 B 0.016994f
C462 VTAIL.n180 B 0.017993f
C463 VTAIL.n181 B 0.040167f
C464 VTAIL.n182 B 0.040167f
C465 VTAIL.n183 B 0.040167f
C466 VTAIL.n184 B 0.017993f
C467 VTAIL.n185 B 0.016994f
C468 VTAIL.n186 B 0.031625f
C469 VTAIL.n187 B 0.031625f
C470 VTAIL.n188 B 0.016994f
C471 VTAIL.n189 B 0.017494f
C472 VTAIL.n190 B 0.017494f
C473 VTAIL.n191 B 0.040167f
C474 VTAIL.n192 B 0.0862f
C475 VTAIL.n193 B 0.017993f
C476 VTAIL.n194 B 0.016994f
C477 VTAIL.n195 B 0.080876f
C478 VTAIL.n196 B 0.048383f
C479 VTAIL.n197 B 1.33419f
C480 VTAIL.t10 B 0.217421f
C481 VTAIL.t7 B 0.217421f
C482 VTAIL.n198 B 1.81598f
C483 VTAIL.n199 B 0.352452f
C484 VN.n0 B 0.053734f
C485 VN.t7 B 0.384304f
C486 VN.t8 B 0.384304f
C487 VN.n1 B 0.021801f
C488 VN.t0 B 0.390907f
C489 VN.t5 B 0.384304f
C490 VN.n2 B 0.162135f
C491 VN.n3 B 0.178401f
C492 VN.n4 B 0.116341f
C493 VN.n5 B 0.053734f
C494 VN.n6 B 0.17996f
C495 VN.n7 B 0.021801f
C496 VN.n8 B 0.162135f
C497 VN.t9 B 0.390907f
C498 VN.n9 B 0.178327f
C499 VN.n10 B 0.041642f
C500 VN.n11 B 0.053734f
C501 VN.t2 B 0.390907f
C502 VN.t4 B 0.384304f
C503 VN.t1 B 0.384304f
C504 VN.n12 B 0.021801f
C505 VN.t3 B 0.384304f
C506 VN.n13 B 0.162135f
C507 VN.t6 B 0.390907f
C508 VN.n14 B 0.178401f
C509 VN.n15 B 0.116341f
C510 VN.n16 B 0.053734f
C511 VN.n17 B 0.17996f
C512 VN.n18 B 0.021801f
C513 VN.n19 B 0.162135f
C514 VN.n20 B 0.178327f
C515 VN.n21 B 1.90921f
.ends

