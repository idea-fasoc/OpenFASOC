* NGSPICE file created from diff_pair_sample_1752.ext - technology: sky130A

.subckt diff_pair_sample_1752 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X1 VTAIL.t3 VN.t0 VDD2.t9 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X2 VDD2.t8 VN.t1 VTAIL.t19 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X3 VDD1.t8 VP.t1 VTAIL.t13 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=1.0374 ps=6.1 w=2.66 l=3.36
X4 B.t11 B.t9 B.t10 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0 ps=0 w=2.66 l=3.36
X5 VDD1.t7 VP.t2 VTAIL.t9 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0.4389 ps=2.99 w=2.66 l=3.36
X6 VDD2.t7 VN.t2 VTAIL.t2 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=1.0374 ps=6.1 w=2.66 l=3.36
X7 VDD2.t6 VN.t3 VTAIL.t18 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0.4389 ps=2.99 w=2.66 l=3.36
X8 VDD2.t5 VN.t4 VTAIL.t17 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=1.0374 ps=6.1 w=2.66 l=3.36
X9 VTAIL.t4 VN.t5 VDD2.t4 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X10 B.t8 B.t6 B.t7 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0 ps=0 w=2.66 l=3.36
X11 VTAIL.t10 VP.t3 VDD1.t6 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X12 VDD1.t5 VP.t4 VTAIL.t8 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0.4389 ps=2.99 w=2.66 l=3.36
X13 VTAIL.t7 VP.t5 VDD1.t4 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X14 B.t5 B.t3 B.t4 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0 ps=0 w=2.66 l=3.36
X15 VTAIL.t12 VP.t6 VDD1.t3 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X16 VDD1.t2 VP.t7 VTAIL.t11 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X17 B.t2 B.t0 B.t1 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0 ps=0 w=2.66 l=3.36
X18 VTAIL.t15 VP.t8 VDD1.t1 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X19 VDD2.t3 VN.t6 VTAIL.t5 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=1.0374 pd=6.1 as=0.4389 ps=2.99 w=2.66 l=3.36
X20 VDD2.t2 VN.t7 VTAIL.t16 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X21 VTAIL.t0 VN.t8 VDD2.t1 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
X22 VDD1.t0 VP.t9 VTAIL.t6 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=1.0374 ps=6.1 w=2.66 l=3.36
X23 VTAIL.t1 VN.t9 VDD2.t0 w_n5398_n1500# sky130_fd_pr__pfet_01v8 ad=0.4389 pd=2.99 as=0.4389 ps=2.99 w=2.66 l=3.36
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n21 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n57 VP.n20 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n19 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n18 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n115 VP.n114 161.3
R23 VP.n113 VP.n1 161.3
R24 VP.n112 VP.n111 161.3
R25 VP.n110 VP.n2 161.3
R26 VP.n109 VP.n108 161.3
R27 VP.n107 VP.n3 161.3
R28 VP.n106 VP.n105 161.3
R29 VP.n104 VP.n4 161.3
R30 VP.n103 VP.n102 161.3
R31 VP.n100 VP.n5 161.3
R32 VP.n99 VP.n98 161.3
R33 VP.n97 VP.n6 161.3
R34 VP.n96 VP.n95 161.3
R35 VP.n94 VP.n7 161.3
R36 VP.n93 VP.n92 161.3
R37 VP.n91 VP.n90 161.3
R38 VP.n89 VP.n9 161.3
R39 VP.n88 VP.n87 161.3
R40 VP.n86 VP.n10 161.3
R41 VP.n85 VP.n84 161.3
R42 VP.n83 VP.n11 161.3
R43 VP.n82 VP.n81 161.3
R44 VP.n80 VP.n79 161.3
R45 VP.n78 VP.n13 161.3
R46 VP.n77 VP.n76 161.3
R47 VP.n75 VP.n14 161.3
R48 VP.n74 VP.n73 161.3
R49 VP.n72 VP.n15 161.3
R50 VP.n71 VP.n70 161.3
R51 VP.n69 VP.n16 161.3
R52 VP.n68 VP.n67 83.8517
R53 VP.n116 VP.n0 83.8517
R54 VP.n66 VP.n17 83.8517
R55 VP.n108 VP.n2 56.5617
R56 VP.n73 VP.n14 56.5617
R57 VP.n58 VP.n19 56.5617
R58 VP.n30 VP.n29 53.0779
R59 VP.n30 VP.t2 51.8941
R60 VP.n68 VP.n66 50.17
R61 VP.n84 VP.n10 49.7803
R62 VP.n99 VP.n6 49.7803
R63 VP.n49 VP.n23 49.7803
R64 VP.n34 VP.n27 49.7803
R65 VP.n88 VP.n10 31.3737
R66 VP.n95 VP.n6 31.3737
R67 VP.n45 VP.n23 31.3737
R68 VP.n38 VP.n27 31.3737
R69 VP.n71 VP.n16 24.5923
R70 VP.n72 VP.n71 24.5923
R71 VP.n73 VP.n72 24.5923
R72 VP.n77 VP.n14 24.5923
R73 VP.n78 VP.n77 24.5923
R74 VP.n79 VP.n78 24.5923
R75 VP.n83 VP.n82 24.5923
R76 VP.n84 VP.n83 24.5923
R77 VP.n89 VP.n88 24.5923
R78 VP.n90 VP.n89 24.5923
R79 VP.n94 VP.n93 24.5923
R80 VP.n95 VP.n94 24.5923
R81 VP.n100 VP.n99 24.5923
R82 VP.n102 VP.n100 24.5923
R83 VP.n106 VP.n4 24.5923
R84 VP.n107 VP.n106 24.5923
R85 VP.n108 VP.n107 24.5923
R86 VP.n112 VP.n2 24.5923
R87 VP.n113 VP.n112 24.5923
R88 VP.n114 VP.n113 24.5923
R89 VP.n62 VP.n19 24.5923
R90 VP.n63 VP.n62 24.5923
R91 VP.n64 VP.n63 24.5923
R92 VP.n50 VP.n49 24.5923
R93 VP.n52 VP.n50 24.5923
R94 VP.n56 VP.n21 24.5923
R95 VP.n57 VP.n56 24.5923
R96 VP.n58 VP.n57 24.5923
R97 VP.n39 VP.n38 24.5923
R98 VP.n40 VP.n39 24.5923
R99 VP.n44 VP.n43 24.5923
R100 VP.n45 VP.n44 24.5923
R101 VP.n33 VP.n32 24.5923
R102 VP.n34 VP.n33 24.5923
R103 VP.n82 VP.n12 21.6413
R104 VP.n102 VP.n101 21.6413
R105 VP.n52 VP.n51 21.6413
R106 VP.n32 VP.n29 21.6413
R107 VP.n67 VP.t4 19.0797
R108 VP.n12 VP.t5 19.0797
R109 VP.n8 VP.t7 19.0797
R110 VP.n101 VP.t3 19.0797
R111 VP.n0 VP.t9 19.0797
R112 VP.n17 VP.t1 19.0797
R113 VP.n51 VP.t6 19.0797
R114 VP.n25 VP.t0 19.0797
R115 VP.n29 VP.t8 19.0797
R116 VP.n90 VP.n8 12.2964
R117 VP.n93 VP.n8 12.2964
R118 VP.n40 VP.n25 12.2964
R119 VP.n43 VP.n25 12.2964
R120 VP.n67 VP.n16 6.39438
R121 VP.n114 VP.n0 6.39438
R122 VP.n64 VP.n17 6.39438
R123 VP.n31 VP.n30 3.26267
R124 VP.n79 VP.n12 2.95152
R125 VP.n101 VP.n4 2.95152
R126 VP.n51 VP.n21 2.95152
R127 VP.n66 VP.n65 0.354861
R128 VP.n69 VP.n68 0.354861
R129 VP.n116 VP.n115 0.354861
R130 VP VP.n116 0.267071
R131 VP.n31 VP.n28 0.189894
R132 VP.n35 VP.n28 0.189894
R133 VP.n36 VP.n35 0.189894
R134 VP.n37 VP.n36 0.189894
R135 VP.n37 VP.n26 0.189894
R136 VP.n41 VP.n26 0.189894
R137 VP.n42 VP.n41 0.189894
R138 VP.n42 VP.n24 0.189894
R139 VP.n46 VP.n24 0.189894
R140 VP.n47 VP.n46 0.189894
R141 VP.n48 VP.n47 0.189894
R142 VP.n48 VP.n22 0.189894
R143 VP.n53 VP.n22 0.189894
R144 VP.n54 VP.n53 0.189894
R145 VP.n55 VP.n54 0.189894
R146 VP.n55 VP.n20 0.189894
R147 VP.n59 VP.n20 0.189894
R148 VP.n60 VP.n59 0.189894
R149 VP.n61 VP.n60 0.189894
R150 VP.n61 VP.n18 0.189894
R151 VP.n65 VP.n18 0.189894
R152 VP.n70 VP.n69 0.189894
R153 VP.n70 VP.n15 0.189894
R154 VP.n74 VP.n15 0.189894
R155 VP.n75 VP.n74 0.189894
R156 VP.n76 VP.n75 0.189894
R157 VP.n76 VP.n13 0.189894
R158 VP.n80 VP.n13 0.189894
R159 VP.n81 VP.n80 0.189894
R160 VP.n81 VP.n11 0.189894
R161 VP.n85 VP.n11 0.189894
R162 VP.n86 VP.n85 0.189894
R163 VP.n87 VP.n86 0.189894
R164 VP.n87 VP.n9 0.189894
R165 VP.n91 VP.n9 0.189894
R166 VP.n92 VP.n91 0.189894
R167 VP.n92 VP.n7 0.189894
R168 VP.n96 VP.n7 0.189894
R169 VP.n97 VP.n96 0.189894
R170 VP.n98 VP.n97 0.189894
R171 VP.n98 VP.n5 0.189894
R172 VP.n103 VP.n5 0.189894
R173 VP.n104 VP.n103 0.189894
R174 VP.n105 VP.n104 0.189894
R175 VP.n105 VP.n3 0.189894
R176 VP.n109 VP.n3 0.189894
R177 VP.n110 VP.n109 0.189894
R178 VP.n111 VP.n110 0.189894
R179 VP.n111 VP.n1 0.189894
R180 VP.n115 VP.n1 0.189894
R181 VTAIL.n56 VTAIL.n50 756.745
R182 VTAIL.n8 VTAIL.n2 756.745
R183 VTAIL.n44 VTAIL.n38 756.745
R184 VTAIL.n28 VTAIL.n22 756.745
R185 VTAIL.n55 VTAIL.n54 585
R186 VTAIL.n57 VTAIL.n56 585
R187 VTAIL.n7 VTAIL.n6 585
R188 VTAIL.n9 VTAIL.n8 585
R189 VTAIL.n45 VTAIL.n44 585
R190 VTAIL.n43 VTAIL.n42 585
R191 VTAIL.n29 VTAIL.n28 585
R192 VTAIL.n27 VTAIL.n26 585
R193 VTAIL.n53 VTAIL.t17 357.269
R194 VTAIL.n5 VTAIL.t6 357.269
R195 VTAIL.n41 VTAIL.t13 357.269
R196 VTAIL.n25 VTAIL.t2 357.269
R197 VTAIL.n56 VTAIL.n55 171.744
R198 VTAIL.n8 VTAIL.n7 171.744
R199 VTAIL.n44 VTAIL.n43 171.744
R200 VTAIL.n28 VTAIL.n27 171.744
R201 VTAIL.n63 VTAIL.n62 134.511
R202 VTAIL.n1 VTAIL.n0 134.511
R203 VTAIL.n15 VTAIL.n14 134.511
R204 VTAIL.n17 VTAIL.n16 134.511
R205 VTAIL.n37 VTAIL.n36 134.511
R206 VTAIL.n35 VTAIL.n34 134.511
R207 VTAIL.n21 VTAIL.n20 134.511
R208 VTAIL.n19 VTAIL.n18 134.511
R209 VTAIL.n55 VTAIL.t17 85.8723
R210 VTAIL.n7 VTAIL.t6 85.8723
R211 VTAIL.n43 VTAIL.t13 85.8723
R212 VTAIL.n27 VTAIL.t2 85.8723
R213 VTAIL.n61 VTAIL.n60 30.246
R214 VTAIL.n13 VTAIL.n12 30.246
R215 VTAIL.n49 VTAIL.n48 30.246
R216 VTAIL.n33 VTAIL.n32 30.246
R217 VTAIL.n19 VTAIL.n17 21.0221
R218 VTAIL.n61 VTAIL.n49 17.841
R219 VTAIL.n62 VTAIL.t19 12.2204
R220 VTAIL.n62 VTAIL.t0 12.2204
R221 VTAIL.n0 VTAIL.t5 12.2204
R222 VTAIL.n0 VTAIL.t4 12.2204
R223 VTAIL.n14 VTAIL.t11 12.2204
R224 VTAIL.n14 VTAIL.t10 12.2204
R225 VTAIL.n16 VTAIL.t8 12.2204
R226 VTAIL.n16 VTAIL.t7 12.2204
R227 VTAIL.n36 VTAIL.t14 12.2204
R228 VTAIL.n36 VTAIL.t12 12.2204
R229 VTAIL.n34 VTAIL.t9 12.2204
R230 VTAIL.n34 VTAIL.t15 12.2204
R231 VTAIL.n20 VTAIL.t16 12.2204
R232 VTAIL.n20 VTAIL.t1 12.2204
R233 VTAIL.n18 VTAIL.t18 12.2204
R234 VTAIL.n18 VTAIL.t3 12.2204
R235 VTAIL.n54 VTAIL.n53 10.3978
R236 VTAIL.n6 VTAIL.n5 10.3978
R237 VTAIL.n42 VTAIL.n41 10.3978
R238 VTAIL.n26 VTAIL.n25 10.3978
R239 VTAIL.n60 VTAIL.n59 9.45567
R240 VTAIL.n12 VTAIL.n11 9.45567
R241 VTAIL.n48 VTAIL.n47 9.45567
R242 VTAIL.n32 VTAIL.n31 9.45567
R243 VTAIL.n52 VTAIL.n51 9.3005
R244 VTAIL.n59 VTAIL.n58 9.3005
R245 VTAIL.n4 VTAIL.n3 9.3005
R246 VTAIL.n11 VTAIL.n10 9.3005
R247 VTAIL.n40 VTAIL.n39 9.3005
R248 VTAIL.n47 VTAIL.n46 9.3005
R249 VTAIL.n31 VTAIL.n30 9.3005
R250 VTAIL.n24 VTAIL.n23 9.3005
R251 VTAIL.n60 VTAIL.n50 8.92171
R252 VTAIL.n12 VTAIL.n2 8.92171
R253 VTAIL.n48 VTAIL.n38 8.92171
R254 VTAIL.n32 VTAIL.n22 8.92171
R255 VTAIL.n58 VTAIL.n57 8.14595
R256 VTAIL.n10 VTAIL.n9 8.14595
R257 VTAIL.n46 VTAIL.n45 8.14595
R258 VTAIL.n30 VTAIL.n29 8.14595
R259 VTAIL.n54 VTAIL.n52 7.3702
R260 VTAIL.n6 VTAIL.n4 7.3702
R261 VTAIL.n42 VTAIL.n40 7.3702
R262 VTAIL.n26 VTAIL.n24 7.3702
R263 VTAIL.n57 VTAIL.n52 5.81868
R264 VTAIL.n9 VTAIL.n4 5.81868
R265 VTAIL.n45 VTAIL.n40 5.81868
R266 VTAIL.n29 VTAIL.n24 5.81868
R267 VTAIL.n58 VTAIL.n50 5.04292
R268 VTAIL.n10 VTAIL.n2 5.04292
R269 VTAIL.n46 VTAIL.n38 5.04292
R270 VTAIL.n30 VTAIL.n22 5.04292
R271 VTAIL.n21 VTAIL.n19 3.18153
R272 VTAIL.n33 VTAIL.n21 3.18153
R273 VTAIL.n37 VTAIL.n35 3.18153
R274 VTAIL.n49 VTAIL.n37 3.18153
R275 VTAIL.n17 VTAIL.n15 3.18153
R276 VTAIL.n15 VTAIL.n13 3.18153
R277 VTAIL.n63 VTAIL.n61 3.18153
R278 VTAIL.n53 VTAIL.n51 2.74506
R279 VTAIL.n5 VTAIL.n3 2.74506
R280 VTAIL.n41 VTAIL.n39 2.74506
R281 VTAIL.n25 VTAIL.n23 2.74506
R282 VTAIL VTAIL.n1 2.44447
R283 VTAIL.n35 VTAIL.n33 2.06084
R284 VTAIL.n13 VTAIL.n1 2.06084
R285 VTAIL VTAIL.n63 0.737569
R286 VTAIL.n59 VTAIL.n51 0.155672
R287 VTAIL.n11 VTAIL.n3 0.155672
R288 VTAIL.n47 VTAIL.n39 0.155672
R289 VTAIL.n31 VTAIL.n23 0.155672
R290 VDD1.n6 VDD1.n0 756.745
R291 VDD1.n19 VDD1.n13 756.745
R292 VDD1.n7 VDD1.n6 585
R293 VDD1.n5 VDD1.n4 585
R294 VDD1.n18 VDD1.n17 585
R295 VDD1.n20 VDD1.n19 585
R296 VDD1.n16 VDD1.t5 357.269
R297 VDD1.n3 VDD1.t7 357.269
R298 VDD1.n6 VDD1.n5 171.744
R299 VDD1.n19 VDD1.n18 171.744
R300 VDD1.n27 VDD1.n26 153.519
R301 VDD1.n29 VDD1.n28 151.19
R302 VDD1.n12 VDD1.n11 151.19
R303 VDD1.n25 VDD1.n24 151.19
R304 VDD1.n5 VDD1.t7 85.8723
R305 VDD1.n18 VDD1.t5 85.8723
R306 VDD1.n12 VDD1.n10 50.1058
R307 VDD1.n25 VDD1.n23 50.1058
R308 VDD1.n29 VDD1.n27 43.2918
R309 VDD1.n28 VDD1.t3 12.2204
R310 VDD1.n28 VDD1.t8 12.2204
R311 VDD1.n11 VDD1.t1 12.2204
R312 VDD1.n11 VDD1.t9 12.2204
R313 VDD1.n26 VDD1.t6 12.2204
R314 VDD1.n26 VDD1.t0 12.2204
R315 VDD1.n24 VDD1.t4 12.2204
R316 VDD1.n24 VDD1.t2 12.2204
R317 VDD1.n4 VDD1.n3 10.3978
R318 VDD1.n17 VDD1.n16 10.3978
R319 VDD1.n10 VDD1.n9 9.45567
R320 VDD1.n23 VDD1.n22 9.45567
R321 VDD1.n9 VDD1.n8 9.3005
R322 VDD1.n2 VDD1.n1 9.3005
R323 VDD1.n15 VDD1.n14 9.3005
R324 VDD1.n22 VDD1.n21 9.3005
R325 VDD1.n10 VDD1.n0 8.92171
R326 VDD1.n23 VDD1.n13 8.92171
R327 VDD1.n8 VDD1.n7 8.14595
R328 VDD1.n21 VDD1.n20 8.14595
R329 VDD1.n4 VDD1.n2 7.3702
R330 VDD1.n17 VDD1.n15 7.3702
R331 VDD1.n7 VDD1.n2 5.81868
R332 VDD1.n20 VDD1.n15 5.81868
R333 VDD1.n8 VDD1.n0 5.04292
R334 VDD1.n21 VDD1.n13 5.04292
R335 VDD1.n3 VDD1.n1 2.74506
R336 VDD1.n16 VDD1.n14 2.74506
R337 VDD1 VDD1.n29 2.32809
R338 VDD1 VDD1.n12 0.853948
R339 VDD1.n27 VDD1.n25 0.740413
R340 VDD1.n9 VDD1.n1 0.155672
R341 VDD1.n22 VDD1.n14 0.155672
R342 VN.n98 VN.n97 161.3
R343 VN.n96 VN.n51 161.3
R344 VN.n95 VN.n94 161.3
R345 VN.n93 VN.n52 161.3
R346 VN.n92 VN.n91 161.3
R347 VN.n90 VN.n53 161.3
R348 VN.n89 VN.n88 161.3
R349 VN.n87 VN.n54 161.3
R350 VN.n86 VN.n85 161.3
R351 VN.n84 VN.n55 161.3
R352 VN.n83 VN.n82 161.3
R353 VN.n81 VN.n57 161.3
R354 VN.n80 VN.n79 161.3
R355 VN.n78 VN.n58 161.3
R356 VN.n77 VN.n76 161.3
R357 VN.n75 VN.n74 161.3
R358 VN.n73 VN.n60 161.3
R359 VN.n72 VN.n71 161.3
R360 VN.n70 VN.n61 161.3
R361 VN.n69 VN.n68 161.3
R362 VN.n67 VN.n62 161.3
R363 VN.n66 VN.n65 161.3
R364 VN.n48 VN.n47 161.3
R365 VN.n46 VN.n1 161.3
R366 VN.n45 VN.n44 161.3
R367 VN.n43 VN.n2 161.3
R368 VN.n42 VN.n41 161.3
R369 VN.n40 VN.n3 161.3
R370 VN.n39 VN.n38 161.3
R371 VN.n37 VN.n4 161.3
R372 VN.n36 VN.n35 161.3
R373 VN.n33 VN.n5 161.3
R374 VN.n32 VN.n31 161.3
R375 VN.n30 VN.n6 161.3
R376 VN.n29 VN.n28 161.3
R377 VN.n27 VN.n7 161.3
R378 VN.n26 VN.n25 161.3
R379 VN.n24 VN.n23 161.3
R380 VN.n22 VN.n9 161.3
R381 VN.n21 VN.n20 161.3
R382 VN.n19 VN.n10 161.3
R383 VN.n18 VN.n17 161.3
R384 VN.n16 VN.n11 161.3
R385 VN.n15 VN.n14 161.3
R386 VN.n49 VN.n0 83.8517
R387 VN.n99 VN.n50 83.8517
R388 VN.n41 VN.n2 56.5617
R389 VN.n91 VN.n52 56.5617
R390 VN.n13 VN.n12 53.0779
R391 VN.n64 VN.n63 53.0779
R392 VN.n64 VN.t2 51.8942
R393 VN.n13 VN.t6 51.8942
R394 VN VN.n99 50.3353
R395 VN.n17 VN.n10 49.7803
R396 VN.n32 VN.n6 49.7803
R397 VN.n68 VN.n61 49.7803
R398 VN.n83 VN.n57 49.7803
R399 VN.n21 VN.n10 31.3737
R400 VN.n28 VN.n6 31.3737
R401 VN.n72 VN.n61 31.3737
R402 VN.n79 VN.n57 31.3737
R403 VN.n16 VN.n15 24.5923
R404 VN.n17 VN.n16 24.5923
R405 VN.n22 VN.n21 24.5923
R406 VN.n23 VN.n22 24.5923
R407 VN.n27 VN.n26 24.5923
R408 VN.n28 VN.n27 24.5923
R409 VN.n33 VN.n32 24.5923
R410 VN.n35 VN.n33 24.5923
R411 VN.n39 VN.n4 24.5923
R412 VN.n40 VN.n39 24.5923
R413 VN.n41 VN.n40 24.5923
R414 VN.n45 VN.n2 24.5923
R415 VN.n46 VN.n45 24.5923
R416 VN.n47 VN.n46 24.5923
R417 VN.n68 VN.n67 24.5923
R418 VN.n67 VN.n66 24.5923
R419 VN.n79 VN.n78 24.5923
R420 VN.n78 VN.n77 24.5923
R421 VN.n74 VN.n73 24.5923
R422 VN.n73 VN.n72 24.5923
R423 VN.n91 VN.n90 24.5923
R424 VN.n90 VN.n89 24.5923
R425 VN.n89 VN.n54 24.5923
R426 VN.n85 VN.n84 24.5923
R427 VN.n84 VN.n83 24.5923
R428 VN.n97 VN.n96 24.5923
R429 VN.n96 VN.n95 24.5923
R430 VN.n95 VN.n52 24.5923
R431 VN.n15 VN.n12 21.6413
R432 VN.n35 VN.n34 21.6413
R433 VN.n66 VN.n63 21.6413
R434 VN.n85 VN.n56 21.6413
R435 VN.n12 VN.t5 19.0797
R436 VN.n8 VN.t1 19.0797
R437 VN.n34 VN.t8 19.0797
R438 VN.n0 VN.t4 19.0797
R439 VN.n63 VN.t9 19.0797
R440 VN.n59 VN.t7 19.0797
R441 VN.n56 VN.t0 19.0797
R442 VN.n50 VN.t3 19.0797
R443 VN.n23 VN.n8 12.2964
R444 VN.n26 VN.n8 12.2964
R445 VN.n77 VN.n59 12.2964
R446 VN.n74 VN.n59 12.2964
R447 VN.n47 VN.n0 6.39438
R448 VN.n97 VN.n50 6.39438
R449 VN.n65 VN.n64 3.26269
R450 VN.n14 VN.n13 3.26269
R451 VN.n34 VN.n4 2.95152
R452 VN.n56 VN.n54 2.95152
R453 VN.n99 VN.n98 0.354861
R454 VN.n49 VN.n48 0.354861
R455 VN VN.n49 0.267071
R456 VN.n98 VN.n51 0.189894
R457 VN.n94 VN.n51 0.189894
R458 VN.n94 VN.n93 0.189894
R459 VN.n93 VN.n92 0.189894
R460 VN.n92 VN.n53 0.189894
R461 VN.n88 VN.n53 0.189894
R462 VN.n88 VN.n87 0.189894
R463 VN.n87 VN.n86 0.189894
R464 VN.n86 VN.n55 0.189894
R465 VN.n82 VN.n55 0.189894
R466 VN.n82 VN.n81 0.189894
R467 VN.n81 VN.n80 0.189894
R468 VN.n80 VN.n58 0.189894
R469 VN.n76 VN.n58 0.189894
R470 VN.n76 VN.n75 0.189894
R471 VN.n75 VN.n60 0.189894
R472 VN.n71 VN.n60 0.189894
R473 VN.n71 VN.n70 0.189894
R474 VN.n70 VN.n69 0.189894
R475 VN.n69 VN.n62 0.189894
R476 VN.n65 VN.n62 0.189894
R477 VN.n14 VN.n11 0.189894
R478 VN.n18 VN.n11 0.189894
R479 VN.n19 VN.n18 0.189894
R480 VN.n20 VN.n19 0.189894
R481 VN.n20 VN.n9 0.189894
R482 VN.n24 VN.n9 0.189894
R483 VN.n25 VN.n24 0.189894
R484 VN.n25 VN.n7 0.189894
R485 VN.n29 VN.n7 0.189894
R486 VN.n30 VN.n29 0.189894
R487 VN.n31 VN.n30 0.189894
R488 VN.n31 VN.n5 0.189894
R489 VN.n36 VN.n5 0.189894
R490 VN.n37 VN.n36 0.189894
R491 VN.n38 VN.n37 0.189894
R492 VN.n38 VN.n3 0.189894
R493 VN.n42 VN.n3 0.189894
R494 VN.n43 VN.n42 0.189894
R495 VN.n44 VN.n43 0.189894
R496 VN.n44 VN.n1 0.189894
R497 VN.n48 VN.n1 0.189894
R498 VDD2.n21 VDD2.n15 756.745
R499 VDD2.n6 VDD2.n0 756.745
R500 VDD2.n22 VDD2.n21 585
R501 VDD2.n20 VDD2.n19 585
R502 VDD2.n5 VDD2.n4 585
R503 VDD2.n7 VDD2.n6 585
R504 VDD2.n3 VDD2.t3 357.269
R505 VDD2.n18 VDD2.t6 357.269
R506 VDD2.n21 VDD2.n20 171.744
R507 VDD2.n6 VDD2.n5 171.744
R508 VDD2.n14 VDD2.n13 153.519
R509 VDD2 VDD2.n29 153.518
R510 VDD2.n28 VDD2.n27 151.19
R511 VDD2.n12 VDD2.n11 151.19
R512 VDD2.n20 VDD2.t6 85.8723
R513 VDD2.n5 VDD2.t3 85.8723
R514 VDD2.n12 VDD2.n10 50.1058
R515 VDD2.n26 VDD2.n25 46.9247
R516 VDD2.n26 VDD2.n14 41.1183
R517 VDD2.n29 VDD2.t0 12.2204
R518 VDD2.n29 VDD2.t7 12.2204
R519 VDD2.n27 VDD2.t9 12.2204
R520 VDD2.n27 VDD2.t2 12.2204
R521 VDD2.n13 VDD2.t1 12.2204
R522 VDD2.n13 VDD2.t5 12.2204
R523 VDD2.n11 VDD2.t4 12.2204
R524 VDD2.n11 VDD2.t8 12.2204
R525 VDD2.n19 VDD2.n18 10.3978
R526 VDD2.n4 VDD2.n3 10.3978
R527 VDD2.n25 VDD2.n24 9.45567
R528 VDD2.n10 VDD2.n9 9.45567
R529 VDD2.n24 VDD2.n23 9.3005
R530 VDD2.n17 VDD2.n16 9.3005
R531 VDD2.n2 VDD2.n1 9.3005
R532 VDD2.n9 VDD2.n8 9.3005
R533 VDD2.n25 VDD2.n15 8.92171
R534 VDD2.n10 VDD2.n0 8.92171
R535 VDD2.n23 VDD2.n22 8.14595
R536 VDD2.n8 VDD2.n7 8.14595
R537 VDD2.n19 VDD2.n17 7.3702
R538 VDD2.n4 VDD2.n2 7.3702
R539 VDD2.n22 VDD2.n17 5.81868
R540 VDD2.n7 VDD2.n2 5.81868
R541 VDD2.n23 VDD2.n15 5.04292
R542 VDD2.n8 VDD2.n0 5.04292
R543 VDD2.n28 VDD2.n26 3.18153
R544 VDD2.n18 VDD2.n16 2.74506
R545 VDD2.n3 VDD2.n1 2.74506
R546 VDD2 VDD2.n28 0.853948
R547 VDD2.n14 VDD2.n12 0.740413
R548 VDD2.n24 VDD2.n16 0.155672
R549 VDD2.n9 VDD2.n1 0.155672
R550 B.n583 B.n62 585
R551 B.n585 B.n584 585
R552 B.n586 B.n61 585
R553 B.n588 B.n587 585
R554 B.n589 B.n60 585
R555 B.n591 B.n590 585
R556 B.n592 B.n59 585
R557 B.n594 B.n593 585
R558 B.n595 B.n58 585
R559 B.n597 B.n596 585
R560 B.n598 B.n57 585
R561 B.n600 B.n599 585
R562 B.n601 B.n53 585
R563 B.n603 B.n602 585
R564 B.n604 B.n52 585
R565 B.n606 B.n605 585
R566 B.n607 B.n51 585
R567 B.n609 B.n608 585
R568 B.n610 B.n50 585
R569 B.n612 B.n611 585
R570 B.n613 B.n49 585
R571 B.n615 B.n614 585
R572 B.n616 B.n48 585
R573 B.n618 B.n617 585
R574 B.n620 B.n45 585
R575 B.n622 B.n621 585
R576 B.n623 B.n44 585
R577 B.n625 B.n624 585
R578 B.n626 B.n43 585
R579 B.n628 B.n627 585
R580 B.n629 B.n42 585
R581 B.n631 B.n630 585
R582 B.n632 B.n41 585
R583 B.n634 B.n633 585
R584 B.n635 B.n40 585
R585 B.n637 B.n636 585
R586 B.n638 B.n39 585
R587 B.n640 B.n639 585
R588 B.n582 B.n581 585
R589 B.n580 B.n63 585
R590 B.n579 B.n578 585
R591 B.n577 B.n64 585
R592 B.n576 B.n575 585
R593 B.n574 B.n65 585
R594 B.n573 B.n572 585
R595 B.n571 B.n66 585
R596 B.n570 B.n569 585
R597 B.n568 B.n67 585
R598 B.n567 B.n566 585
R599 B.n565 B.n68 585
R600 B.n564 B.n563 585
R601 B.n562 B.n69 585
R602 B.n561 B.n560 585
R603 B.n559 B.n70 585
R604 B.n558 B.n557 585
R605 B.n556 B.n71 585
R606 B.n555 B.n554 585
R607 B.n553 B.n72 585
R608 B.n552 B.n551 585
R609 B.n550 B.n73 585
R610 B.n549 B.n548 585
R611 B.n547 B.n74 585
R612 B.n546 B.n545 585
R613 B.n544 B.n75 585
R614 B.n543 B.n542 585
R615 B.n541 B.n76 585
R616 B.n540 B.n539 585
R617 B.n538 B.n77 585
R618 B.n537 B.n536 585
R619 B.n535 B.n78 585
R620 B.n534 B.n533 585
R621 B.n532 B.n79 585
R622 B.n531 B.n530 585
R623 B.n529 B.n80 585
R624 B.n528 B.n527 585
R625 B.n526 B.n81 585
R626 B.n525 B.n524 585
R627 B.n523 B.n82 585
R628 B.n522 B.n521 585
R629 B.n520 B.n83 585
R630 B.n519 B.n518 585
R631 B.n517 B.n84 585
R632 B.n516 B.n515 585
R633 B.n514 B.n85 585
R634 B.n513 B.n512 585
R635 B.n511 B.n86 585
R636 B.n510 B.n509 585
R637 B.n508 B.n87 585
R638 B.n507 B.n506 585
R639 B.n505 B.n88 585
R640 B.n504 B.n503 585
R641 B.n502 B.n89 585
R642 B.n501 B.n500 585
R643 B.n499 B.n90 585
R644 B.n498 B.n497 585
R645 B.n496 B.n91 585
R646 B.n495 B.n494 585
R647 B.n493 B.n92 585
R648 B.n492 B.n491 585
R649 B.n490 B.n93 585
R650 B.n489 B.n488 585
R651 B.n487 B.n94 585
R652 B.n486 B.n485 585
R653 B.n484 B.n95 585
R654 B.n483 B.n482 585
R655 B.n481 B.n96 585
R656 B.n480 B.n479 585
R657 B.n478 B.n97 585
R658 B.n477 B.n476 585
R659 B.n475 B.n98 585
R660 B.n474 B.n473 585
R661 B.n472 B.n99 585
R662 B.n471 B.n470 585
R663 B.n469 B.n100 585
R664 B.n468 B.n467 585
R665 B.n466 B.n101 585
R666 B.n465 B.n464 585
R667 B.n463 B.n102 585
R668 B.n462 B.n461 585
R669 B.n460 B.n103 585
R670 B.n459 B.n458 585
R671 B.n457 B.n104 585
R672 B.n456 B.n455 585
R673 B.n454 B.n105 585
R674 B.n453 B.n452 585
R675 B.n451 B.n106 585
R676 B.n450 B.n449 585
R677 B.n448 B.n107 585
R678 B.n447 B.n446 585
R679 B.n445 B.n108 585
R680 B.n444 B.n443 585
R681 B.n442 B.n109 585
R682 B.n441 B.n440 585
R683 B.n439 B.n110 585
R684 B.n438 B.n437 585
R685 B.n436 B.n111 585
R686 B.n435 B.n434 585
R687 B.n433 B.n112 585
R688 B.n432 B.n431 585
R689 B.n430 B.n113 585
R690 B.n429 B.n428 585
R691 B.n427 B.n114 585
R692 B.n426 B.n425 585
R693 B.n424 B.n115 585
R694 B.n423 B.n422 585
R695 B.n421 B.n116 585
R696 B.n420 B.n419 585
R697 B.n418 B.n117 585
R698 B.n417 B.n416 585
R699 B.n415 B.n118 585
R700 B.n414 B.n413 585
R701 B.n412 B.n119 585
R702 B.n411 B.n410 585
R703 B.n409 B.n120 585
R704 B.n408 B.n407 585
R705 B.n406 B.n121 585
R706 B.n405 B.n404 585
R707 B.n403 B.n122 585
R708 B.n402 B.n401 585
R709 B.n400 B.n123 585
R710 B.n399 B.n398 585
R711 B.n397 B.n124 585
R712 B.n396 B.n395 585
R713 B.n394 B.n125 585
R714 B.n393 B.n392 585
R715 B.n391 B.n126 585
R716 B.n390 B.n389 585
R717 B.n388 B.n127 585
R718 B.n387 B.n386 585
R719 B.n385 B.n128 585
R720 B.n384 B.n383 585
R721 B.n382 B.n129 585
R722 B.n381 B.n380 585
R723 B.n379 B.n130 585
R724 B.n378 B.n377 585
R725 B.n376 B.n131 585
R726 B.n375 B.n374 585
R727 B.n373 B.n132 585
R728 B.n372 B.n371 585
R729 B.n370 B.n133 585
R730 B.n369 B.n368 585
R731 B.n367 B.n134 585
R732 B.n366 B.n365 585
R733 B.n364 B.n135 585
R734 B.n363 B.n362 585
R735 B.n304 B.n159 585
R736 B.n306 B.n305 585
R737 B.n307 B.n158 585
R738 B.n309 B.n308 585
R739 B.n310 B.n157 585
R740 B.n312 B.n311 585
R741 B.n313 B.n156 585
R742 B.n315 B.n314 585
R743 B.n316 B.n155 585
R744 B.n318 B.n317 585
R745 B.n319 B.n154 585
R746 B.n321 B.n320 585
R747 B.n322 B.n153 585
R748 B.n324 B.n323 585
R749 B.n326 B.n150 585
R750 B.n328 B.n327 585
R751 B.n329 B.n149 585
R752 B.n331 B.n330 585
R753 B.n332 B.n148 585
R754 B.n334 B.n333 585
R755 B.n335 B.n147 585
R756 B.n337 B.n336 585
R757 B.n338 B.n146 585
R758 B.n340 B.n339 585
R759 B.n342 B.n341 585
R760 B.n343 B.n142 585
R761 B.n345 B.n344 585
R762 B.n346 B.n141 585
R763 B.n348 B.n347 585
R764 B.n349 B.n140 585
R765 B.n351 B.n350 585
R766 B.n352 B.n139 585
R767 B.n354 B.n353 585
R768 B.n355 B.n138 585
R769 B.n357 B.n356 585
R770 B.n358 B.n137 585
R771 B.n360 B.n359 585
R772 B.n361 B.n136 585
R773 B.n303 B.n302 585
R774 B.n301 B.n160 585
R775 B.n300 B.n299 585
R776 B.n298 B.n161 585
R777 B.n297 B.n296 585
R778 B.n295 B.n162 585
R779 B.n294 B.n293 585
R780 B.n292 B.n163 585
R781 B.n291 B.n290 585
R782 B.n289 B.n164 585
R783 B.n288 B.n287 585
R784 B.n286 B.n165 585
R785 B.n285 B.n284 585
R786 B.n283 B.n166 585
R787 B.n282 B.n281 585
R788 B.n280 B.n167 585
R789 B.n279 B.n278 585
R790 B.n277 B.n168 585
R791 B.n276 B.n275 585
R792 B.n274 B.n169 585
R793 B.n273 B.n272 585
R794 B.n271 B.n170 585
R795 B.n270 B.n269 585
R796 B.n268 B.n171 585
R797 B.n267 B.n266 585
R798 B.n265 B.n172 585
R799 B.n264 B.n263 585
R800 B.n262 B.n173 585
R801 B.n261 B.n260 585
R802 B.n259 B.n174 585
R803 B.n258 B.n257 585
R804 B.n256 B.n175 585
R805 B.n255 B.n254 585
R806 B.n253 B.n176 585
R807 B.n252 B.n251 585
R808 B.n250 B.n177 585
R809 B.n249 B.n248 585
R810 B.n247 B.n178 585
R811 B.n246 B.n245 585
R812 B.n244 B.n179 585
R813 B.n243 B.n242 585
R814 B.n241 B.n180 585
R815 B.n240 B.n239 585
R816 B.n238 B.n181 585
R817 B.n237 B.n236 585
R818 B.n235 B.n182 585
R819 B.n234 B.n233 585
R820 B.n232 B.n183 585
R821 B.n231 B.n230 585
R822 B.n229 B.n184 585
R823 B.n228 B.n227 585
R824 B.n226 B.n185 585
R825 B.n225 B.n224 585
R826 B.n223 B.n186 585
R827 B.n222 B.n221 585
R828 B.n220 B.n187 585
R829 B.n219 B.n218 585
R830 B.n217 B.n188 585
R831 B.n216 B.n215 585
R832 B.n214 B.n189 585
R833 B.n213 B.n212 585
R834 B.n211 B.n190 585
R835 B.n210 B.n209 585
R836 B.n208 B.n191 585
R837 B.n207 B.n206 585
R838 B.n205 B.n192 585
R839 B.n204 B.n203 585
R840 B.n202 B.n193 585
R841 B.n201 B.n200 585
R842 B.n199 B.n194 585
R843 B.n198 B.n197 585
R844 B.n196 B.n195 585
R845 B.n2 B.n0 585
R846 B.n749 B.n1 585
R847 B.n748 B.n747 585
R848 B.n746 B.n3 585
R849 B.n745 B.n744 585
R850 B.n743 B.n4 585
R851 B.n742 B.n741 585
R852 B.n740 B.n5 585
R853 B.n739 B.n738 585
R854 B.n737 B.n6 585
R855 B.n736 B.n735 585
R856 B.n734 B.n7 585
R857 B.n733 B.n732 585
R858 B.n731 B.n8 585
R859 B.n730 B.n729 585
R860 B.n728 B.n9 585
R861 B.n727 B.n726 585
R862 B.n725 B.n10 585
R863 B.n724 B.n723 585
R864 B.n722 B.n11 585
R865 B.n721 B.n720 585
R866 B.n719 B.n12 585
R867 B.n718 B.n717 585
R868 B.n716 B.n13 585
R869 B.n715 B.n714 585
R870 B.n713 B.n14 585
R871 B.n712 B.n711 585
R872 B.n710 B.n15 585
R873 B.n709 B.n708 585
R874 B.n707 B.n16 585
R875 B.n706 B.n705 585
R876 B.n704 B.n17 585
R877 B.n703 B.n702 585
R878 B.n701 B.n18 585
R879 B.n700 B.n699 585
R880 B.n698 B.n19 585
R881 B.n697 B.n696 585
R882 B.n695 B.n20 585
R883 B.n694 B.n693 585
R884 B.n692 B.n21 585
R885 B.n691 B.n690 585
R886 B.n689 B.n22 585
R887 B.n688 B.n687 585
R888 B.n686 B.n23 585
R889 B.n685 B.n684 585
R890 B.n683 B.n24 585
R891 B.n682 B.n681 585
R892 B.n680 B.n25 585
R893 B.n679 B.n678 585
R894 B.n677 B.n26 585
R895 B.n676 B.n675 585
R896 B.n674 B.n27 585
R897 B.n673 B.n672 585
R898 B.n671 B.n28 585
R899 B.n670 B.n669 585
R900 B.n668 B.n29 585
R901 B.n667 B.n666 585
R902 B.n665 B.n30 585
R903 B.n664 B.n663 585
R904 B.n662 B.n31 585
R905 B.n661 B.n660 585
R906 B.n659 B.n32 585
R907 B.n658 B.n657 585
R908 B.n656 B.n33 585
R909 B.n655 B.n654 585
R910 B.n653 B.n34 585
R911 B.n652 B.n651 585
R912 B.n650 B.n35 585
R913 B.n649 B.n648 585
R914 B.n647 B.n36 585
R915 B.n646 B.n645 585
R916 B.n644 B.n37 585
R917 B.n643 B.n642 585
R918 B.n641 B.n38 585
R919 B.n751 B.n750 585
R920 B.n304 B.n303 526.135
R921 B.n641 B.n640 526.135
R922 B.n363 B.n136 526.135
R923 B.n581 B.n62 526.135
R924 B.n143 B.t2 298.918
R925 B.n54 B.t4 298.918
R926 B.n151 B.t8 298.918
R927 B.n46 B.t10 298.918
R928 B.n143 B.t0 228.042
R929 B.n151 B.t6 228.042
R930 B.n46 B.t9 228.042
R931 B.n54 B.t3 228.042
R932 B.n144 B.t1 227.355
R933 B.n55 B.t5 227.355
R934 B.n152 B.t7 227.355
R935 B.n47 B.t11 227.355
R936 B.n303 B.n160 163.367
R937 B.n299 B.n160 163.367
R938 B.n299 B.n298 163.367
R939 B.n298 B.n297 163.367
R940 B.n297 B.n162 163.367
R941 B.n293 B.n162 163.367
R942 B.n293 B.n292 163.367
R943 B.n292 B.n291 163.367
R944 B.n291 B.n164 163.367
R945 B.n287 B.n164 163.367
R946 B.n287 B.n286 163.367
R947 B.n286 B.n285 163.367
R948 B.n285 B.n166 163.367
R949 B.n281 B.n166 163.367
R950 B.n281 B.n280 163.367
R951 B.n280 B.n279 163.367
R952 B.n279 B.n168 163.367
R953 B.n275 B.n168 163.367
R954 B.n275 B.n274 163.367
R955 B.n274 B.n273 163.367
R956 B.n273 B.n170 163.367
R957 B.n269 B.n170 163.367
R958 B.n269 B.n268 163.367
R959 B.n268 B.n267 163.367
R960 B.n267 B.n172 163.367
R961 B.n263 B.n172 163.367
R962 B.n263 B.n262 163.367
R963 B.n262 B.n261 163.367
R964 B.n261 B.n174 163.367
R965 B.n257 B.n174 163.367
R966 B.n257 B.n256 163.367
R967 B.n256 B.n255 163.367
R968 B.n255 B.n176 163.367
R969 B.n251 B.n176 163.367
R970 B.n251 B.n250 163.367
R971 B.n250 B.n249 163.367
R972 B.n249 B.n178 163.367
R973 B.n245 B.n178 163.367
R974 B.n245 B.n244 163.367
R975 B.n244 B.n243 163.367
R976 B.n243 B.n180 163.367
R977 B.n239 B.n180 163.367
R978 B.n239 B.n238 163.367
R979 B.n238 B.n237 163.367
R980 B.n237 B.n182 163.367
R981 B.n233 B.n182 163.367
R982 B.n233 B.n232 163.367
R983 B.n232 B.n231 163.367
R984 B.n231 B.n184 163.367
R985 B.n227 B.n184 163.367
R986 B.n227 B.n226 163.367
R987 B.n226 B.n225 163.367
R988 B.n225 B.n186 163.367
R989 B.n221 B.n186 163.367
R990 B.n221 B.n220 163.367
R991 B.n220 B.n219 163.367
R992 B.n219 B.n188 163.367
R993 B.n215 B.n188 163.367
R994 B.n215 B.n214 163.367
R995 B.n214 B.n213 163.367
R996 B.n213 B.n190 163.367
R997 B.n209 B.n190 163.367
R998 B.n209 B.n208 163.367
R999 B.n208 B.n207 163.367
R1000 B.n207 B.n192 163.367
R1001 B.n203 B.n192 163.367
R1002 B.n203 B.n202 163.367
R1003 B.n202 B.n201 163.367
R1004 B.n201 B.n194 163.367
R1005 B.n197 B.n194 163.367
R1006 B.n197 B.n196 163.367
R1007 B.n196 B.n2 163.367
R1008 B.n750 B.n2 163.367
R1009 B.n750 B.n749 163.367
R1010 B.n749 B.n748 163.367
R1011 B.n748 B.n3 163.367
R1012 B.n744 B.n3 163.367
R1013 B.n744 B.n743 163.367
R1014 B.n743 B.n742 163.367
R1015 B.n742 B.n5 163.367
R1016 B.n738 B.n5 163.367
R1017 B.n738 B.n737 163.367
R1018 B.n737 B.n736 163.367
R1019 B.n736 B.n7 163.367
R1020 B.n732 B.n7 163.367
R1021 B.n732 B.n731 163.367
R1022 B.n731 B.n730 163.367
R1023 B.n730 B.n9 163.367
R1024 B.n726 B.n9 163.367
R1025 B.n726 B.n725 163.367
R1026 B.n725 B.n724 163.367
R1027 B.n724 B.n11 163.367
R1028 B.n720 B.n11 163.367
R1029 B.n720 B.n719 163.367
R1030 B.n719 B.n718 163.367
R1031 B.n718 B.n13 163.367
R1032 B.n714 B.n13 163.367
R1033 B.n714 B.n713 163.367
R1034 B.n713 B.n712 163.367
R1035 B.n712 B.n15 163.367
R1036 B.n708 B.n15 163.367
R1037 B.n708 B.n707 163.367
R1038 B.n707 B.n706 163.367
R1039 B.n706 B.n17 163.367
R1040 B.n702 B.n17 163.367
R1041 B.n702 B.n701 163.367
R1042 B.n701 B.n700 163.367
R1043 B.n700 B.n19 163.367
R1044 B.n696 B.n19 163.367
R1045 B.n696 B.n695 163.367
R1046 B.n695 B.n694 163.367
R1047 B.n694 B.n21 163.367
R1048 B.n690 B.n21 163.367
R1049 B.n690 B.n689 163.367
R1050 B.n689 B.n688 163.367
R1051 B.n688 B.n23 163.367
R1052 B.n684 B.n23 163.367
R1053 B.n684 B.n683 163.367
R1054 B.n683 B.n682 163.367
R1055 B.n682 B.n25 163.367
R1056 B.n678 B.n25 163.367
R1057 B.n678 B.n677 163.367
R1058 B.n677 B.n676 163.367
R1059 B.n676 B.n27 163.367
R1060 B.n672 B.n27 163.367
R1061 B.n672 B.n671 163.367
R1062 B.n671 B.n670 163.367
R1063 B.n670 B.n29 163.367
R1064 B.n666 B.n29 163.367
R1065 B.n666 B.n665 163.367
R1066 B.n665 B.n664 163.367
R1067 B.n664 B.n31 163.367
R1068 B.n660 B.n31 163.367
R1069 B.n660 B.n659 163.367
R1070 B.n659 B.n658 163.367
R1071 B.n658 B.n33 163.367
R1072 B.n654 B.n33 163.367
R1073 B.n654 B.n653 163.367
R1074 B.n653 B.n652 163.367
R1075 B.n652 B.n35 163.367
R1076 B.n648 B.n35 163.367
R1077 B.n648 B.n647 163.367
R1078 B.n647 B.n646 163.367
R1079 B.n646 B.n37 163.367
R1080 B.n642 B.n37 163.367
R1081 B.n642 B.n641 163.367
R1082 B.n305 B.n304 163.367
R1083 B.n305 B.n158 163.367
R1084 B.n309 B.n158 163.367
R1085 B.n310 B.n309 163.367
R1086 B.n311 B.n310 163.367
R1087 B.n311 B.n156 163.367
R1088 B.n315 B.n156 163.367
R1089 B.n316 B.n315 163.367
R1090 B.n317 B.n316 163.367
R1091 B.n317 B.n154 163.367
R1092 B.n321 B.n154 163.367
R1093 B.n322 B.n321 163.367
R1094 B.n323 B.n322 163.367
R1095 B.n323 B.n150 163.367
R1096 B.n328 B.n150 163.367
R1097 B.n329 B.n328 163.367
R1098 B.n330 B.n329 163.367
R1099 B.n330 B.n148 163.367
R1100 B.n334 B.n148 163.367
R1101 B.n335 B.n334 163.367
R1102 B.n336 B.n335 163.367
R1103 B.n336 B.n146 163.367
R1104 B.n340 B.n146 163.367
R1105 B.n341 B.n340 163.367
R1106 B.n341 B.n142 163.367
R1107 B.n345 B.n142 163.367
R1108 B.n346 B.n345 163.367
R1109 B.n347 B.n346 163.367
R1110 B.n347 B.n140 163.367
R1111 B.n351 B.n140 163.367
R1112 B.n352 B.n351 163.367
R1113 B.n353 B.n352 163.367
R1114 B.n353 B.n138 163.367
R1115 B.n357 B.n138 163.367
R1116 B.n358 B.n357 163.367
R1117 B.n359 B.n358 163.367
R1118 B.n359 B.n136 163.367
R1119 B.n364 B.n363 163.367
R1120 B.n365 B.n364 163.367
R1121 B.n365 B.n134 163.367
R1122 B.n369 B.n134 163.367
R1123 B.n370 B.n369 163.367
R1124 B.n371 B.n370 163.367
R1125 B.n371 B.n132 163.367
R1126 B.n375 B.n132 163.367
R1127 B.n376 B.n375 163.367
R1128 B.n377 B.n376 163.367
R1129 B.n377 B.n130 163.367
R1130 B.n381 B.n130 163.367
R1131 B.n382 B.n381 163.367
R1132 B.n383 B.n382 163.367
R1133 B.n383 B.n128 163.367
R1134 B.n387 B.n128 163.367
R1135 B.n388 B.n387 163.367
R1136 B.n389 B.n388 163.367
R1137 B.n389 B.n126 163.367
R1138 B.n393 B.n126 163.367
R1139 B.n394 B.n393 163.367
R1140 B.n395 B.n394 163.367
R1141 B.n395 B.n124 163.367
R1142 B.n399 B.n124 163.367
R1143 B.n400 B.n399 163.367
R1144 B.n401 B.n400 163.367
R1145 B.n401 B.n122 163.367
R1146 B.n405 B.n122 163.367
R1147 B.n406 B.n405 163.367
R1148 B.n407 B.n406 163.367
R1149 B.n407 B.n120 163.367
R1150 B.n411 B.n120 163.367
R1151 B.n412 B.n411 163.367
R1152 B.n413 B.n412 163.367
R1153 B.n413 B.n118 163.367
R1154 B.n417 B.n118 163.367
R1155 B.n418 B.n417 163.367
R1156 B.n419 B.n418 163.367
R1157 B.n419 B.n116 163.367
R1158 B.n423 B.n116 163.367
R1159 B.n424 B.n423 163.367
R1160 B.n425 B.n424 163.367
R1161 B.n425 B.n114 163.367
R1162 B.n429 B.n114 163.367
R1163 B.n430 B.n429 163.367
R1164 B.n431 B.n430 163.367
R1165 B.n431 B.n112 163.367
R1166 B.n435 B.n112 163.367
R1167 B.n436 B.n435 163.367
R1168 B.n437 B.n436 163.367
R1169 B.n437 B.n110 163.367
R1170 B.n441 B.n110 163.367
R1171 B.n442 B.n441 163.367
R1172 B.n443 B.n442 163.367
R1173 B.n443 B.n108 163.367
R1174 B.n447 B.n108 163.367
R1175 B.n448 B.n447 163.367
R1176 B.n449 B.n448 163.367
R1177 B.n449 B.n106 163.367
R1178 B.n453 B.n106 163.367
R1179 B.n454 B.n453 163.367
R1180 B.n455 B.n454 163.367
R1181 B.n455 B.n104 163.367
R1182 B.n459 B.n104 163.367
R1183 B.n460 B.n459 163.367
R1184 B.n461 B.n460 163.367
R1185 B.n461 B.n102 163.367
R1186 B.n465 B.n102 163.367
R1187 B.n466 B.n465 163.367
R1188 B.n467 B.n466 163.367
R1189 B.n467 B.n100 163.367
R1190 B.n471 B.n100 163.367
R1191 B.n472 B.n471 163.367
R1192 B.n473 B.n472 163.367
R1193 B.n473 B.n98 163.367
R1194 B.n477 B.n98 163.367
R1195 B.n478 B.n477 163.367
R1196 B.n479 B.n478 163.367
R1197 B.n479 B.n96 163.367
R1198 B.n483 B.n96 163.367
R1199 B.n484 B.n483 163.367
R1200 B.n485 B.n484 163.367
R1201 B.n485 B.n94 163.367
R1202 B.n489 B.n94 163.367
R1203 B.n490 B.n489 163.367
R1204 B.n491 B.n490 163.367
R1205 B.n491 B.n92 163.367
R1206 B.n495 B.n92 163.367
R1207 B.n496 B.n495 163.367
R1208 B.n497 B.n496 163.367
R1209 B.n497 B.n90 163.367
R1210 B.n501 B.n90 163.367
R1211 B.n502 B.n501 163.367
R1212 B.n503 B.n502 163.367
R1213 B.n503 B.n88 163.367
R1214 B.n507 B.n88 163.367
R1215 B.n508 B.n507 163.367
R1216 B.n509 B.n508 163.367
R1217 B.n509 B.n86 163.367
R1218 B.n513 B.n86 163.367
R1219 B.n514 B.n513 163.367
R1220 B.n515 B.n514 163.367
R1221 B.n515 B.n84 163.367
R1222 B.n519 B.n84 163.367
R1223 B.n520 B.n519 163.367
R1224 B.n521 B.n520 163.367
R1225 B.n521 B.n82 163.367
R1226 B.n525 B.n82 163.367
R1227 B.n526 B.n525 163.367
R1228 B.n527 B.n526 163.367
R1229 B.n527 B.n80 163.367
R1230 B.n531 B.n80 163.367
R1231 B.n532 B.n531 163.367
R1232 B.n533 B.n532 163.367
R1233 B.n533 B.n78 163.367
R1234 B.n537 B.n78 163.367
R1235 B.n538 B.n537 163.367
R1236 B.n539 B.n538 163.367
R1237 B.n539 B.n76 163.367
R1238 B.n543 B.n76 163.367
R1239 B.n544 B.n543 163.367
R1240 B.n545 B.n544 163.367
R1241 B.n545 B.n74 163.367
R1242 B.n549 B.n74 163.367
R1243 B.n550 B.n549 163.367
R1244 B.n551 B.n550 163.367
R1245 B.n551 B.n72 163.367
R1246 B.n555 B.n72 163.367
R1247 B.n556 B.n555 163.367
R1248 B.n557 B.n556 163.367
R1249 B.n557 B.n70 163.367
R1250 B.n561 B.n70 163.367
R1251 B.n562 B.n561 163.367
R1252 B.n563 B.n562 163.367
R1253 B.n563 B.n68 163.367
R1254 B.n567 B.n68 163.367
R1255 B.n568 B.n567 163.367
R1256 B.n569 B.n568 163.367
R1257 B.n569 B.n66 163.367
R1258 B.n573 B.n66 163.367
R1259 B.n574 B.n573 163.367
R1260 B.n575 B.n574 163.367
R1261 B.n575 B.n64 163.367
R1262 B.n579 B.n64 163.367
R1263 B.n580 B.n579 163.367
R1264 B.n581 B.n580 163.367
R1265 B.n640 B.n39 163.367
R1266 B.n636 B.n39 163.367
R1267 B.n636 B.n635 163.367
R1268 B.n635 B.n634 163.367
R1269 B.n634 B.n41 163.367
R1270 B.n630 B.n41 163.367
R1271 B.n630 B.n629 163.367
R1272 B.n629 B.n628 163.367
R1273 B.n628 B.n43 163.367
R1274 B.n624 B.n43 163.367
R1275 B.n624 B.n623 163.367
R1276 B.n623 B.n622 163.367
R1277 B.n622 B.n45 163.367
R1278 B.n617 B.n45 163.367
R1279 B.n617 B.n616 163.367
R1280 B.n616 B.n615 163.367
R1281 B.n615 B.n49 163.367
R1282 B.n611 B.n49 163.367
R1283 B.n611 B.n610 163.367
R1284 B.n610 B.n609 163.367
R1285 B.n609 B.n51 163.367
R1286 B.n605 B.n51 163.367
R1287 B.n605 B.n604 163.367
R1288 B.n604 B.n603 163.367
R1289 B.n603 B.n53 163.367
R1290 B.n599 B.n53 163.367
R1291 B.n599 B.n598 163.367
R1292 B.n598 B.n597 163.367
R1293 B.n597 B.n58 163.367
R1294 B.n593 B.n58 163.367
R1295 B.n593 B.n592 163.367
R1296 B.n592 B.n591 163.367
R1297 B.n591 B.n60 163.367
R1298 B.n587 B.n60 163.367
R1299 B.n587 B.n586 163.367
R1300 B.n586 B.n585 163.367
R1301 B.n585 B.n62 163.367
R1302 B.n144 B.n143 71.5641
R1303 B.n152 B.n151 71.5641
R1304 B.n47 B.n46 71.5641
R1305 B.n55 B.n54 71.5641
R1306 B.n145 B.n144 59.5399
R1307 B.n325 B.n152 59.5399
R1308 B.n619 B.n47 59.5399
R1309 B.n56 B.n55 59.5399
R1310 B.n639 B.n38 34.1859
R1311 B.n583 B.n582 34.1859
R1312 B.n362 B.n361 34.1859
R1313 B.n302 B.n159 34.1859
R1314 B B.n751 18.0485
R1315 B.n639 B.n638 10.6151
R1316 B.n638 B.n637 10.6151
R1317 B.n637 B.n40 10.6151
R1318 B.n633 B.n40 10.6151
R1319 B.n633 B.n632 10.6151
R1320 B.n632 B.n631 10.6151
R1321 B.n631 B.n42 10.6151
R1322 B.n627 B.n42 10.6151
R1323 B.n627 B.n626 10.6151
R1324 B.n626 B.n625 10.6151
R1325 B.n625 B.n44 10.6151
R1326 B.n621 B.n44 10.6151
R1327 B.n621 B.n620 10.6151
R1328 B.n618 B.n48 10.6151
R1329 B.n614 B.n48 10.6151
R1330 B.n614 B.n613 10.6151
R1331 B.n613 B.n612 10.6151
R1332 B.n612 B.n50 10.6151
R1333 B.n608 B.n50 10.6151
R1334 B.n608 B.n607 10.6151
R1335 B.n607 B.n606 10.6151
R1336 B.n606 B.n52 10.6151
R1337 B.n602 B.n601 10.6151
R1338 B.n601 B.n600 10.6151
R1339 B.n600 B.n57 10.6151
R1340 B.n596 B.n57 10.6151
R1341 B.n596 B.n595 10.6151
R1342 B.n595 B.n594 10.6151
R1343 B.n594 B.n59 10.6151
R1344 B.n590 B.n59 10.6151
R1345 B.n590 B.n589 10.6151
R1346 B.n589 B.n588 10.6151
R1347 B.n588 B.n61 10.6151
R1348 B.n584 B.n61 10.6151
R1349 B.n584 B.n583 10.6151
R1350 B.n362 B.n135 10.6151
R1351 B.n366 B.n135 10.6151
R1352 B.n367 B.n366 10.6151
R1353 B.n368 B.n367 10.6151
R1354 B.n368 B.n133 10.6151
R1355 B.n372 B.n133 10.6151
R1356 B.n373 B.n372 10.6151
R1357 B.n374 B.n373 10.6151
R1358 B.n374 B.n131 10.6151
R1359 B.n378 B.n131 10.6151
R1360 B.n379 B.n378 10.6151
R1361 B.n380 B.n379 10.6151
R1362 B.n380 B.n129 10.6151
R1363 B.n384 B.n129 10.6151
R1364 B.n385 B.n384 10.6151
R1365 B.n386 B.n385 10.6151
R1366 B.n386 B.n127 10.6151
R1367 B.n390 B.n127 10.6151
R1368 B.n391 B.n390 10.6151
R1369 B.n392 B.n391 10.6151
R1370 B.n392 B.n125 10.6151
R1371 B.n396 B.n125 10.6151
R1372 B.n397 B.n396 10.6151
R1373 B.n398 B.n397 10.6151
R1374 B.n398 B.n123 10.6151
R1375 B.n402 B.n123 10.6151
R1376 B.n403 B.n402 10.6151
R1377 B.n404 B.n403 10.6151
R1378 B.n404 B.n121 10.6151
R1379 B.n408 B.n121 10.6151
R1380 B.n409 B.n408 10.6151
R1381 B.n410 B.n409 10.6151
R1382 B.n410 B.n119 10.6151
R1383 B.n414 B.n119 10.6151
R1384 B.n415 B.n414 10.6151
R1385 B.n416 B.n415 10.6151
R1386 B.n416 B.n117 10.6151
R1387 B.n420 B.n117 10.6151
R1388 B.n421 B.n420 10.6151
R1389 B.n422 B.n421 10.6151
R1390 B.n422 B.n115 10.6151
R1391 B.n426 B.n115 10.6151
R1392 B.n427 B.n426 10.6151
R1393 B.n428 B.n427 10.6151
R1394 B.n428 B.n113 10.6151
R1395 B.n432 B.n113 10.6151
R1396 B.n433 B.n432 10.6151
R1397 B.n434 B.n433 10.6151
R1398 B.n434 B.n111 10.6151
R1399 B.n438 B.n111 10.6151
R1400 B.n439 B.n438 10.6151
R1401 B.n440 B.n439 10.6151
R1402 B.n440 B.n109 10.6151
R1403 B.n444 B.n109 10.6151
R1404 B.n445 B.n444 10.6151
R1405 B.n446 B.n445 10.6151
R1406 B.n446 B.n107 10.6151
R1407 B.n450 B.n107 10.6151
R1408 B.n451 B.n450 10.6151
R1409 B.n452 B.n451 10.6151
R1410 B.n452 B.n105 10.6151
R1411 B.n456 B.n105 10.6151
R1412 B.n457 B.n456 10.6151
R1413 B.n458 B.n457 10.6151
R1414 B.n458 B.n103 10.6151
R1415 B.n462 B.n103 10.6151
R1416 B.n463 B.n462 10.6151
R1417 B.n464 B.n463 10.6151
R1418 B.n464 B.n101 10.6151
R1419 B.n468 B.n101 10.6151
R1420 B.n469 B.n468 10.6151
R1421 B.n470 B.n469 10.6151
R1422 B.n470 B.n99 10.6151
R1423 B.n474 B.n99 10.6151
R1424 B.n475 B.n474 10.6151
R1425 B.n476 B.n475 10.6151
R1426 B.n476 B.n97 10.6151
R1427 B.n480 B.n97 10.6151
R1428 B.n481 B.n480 10.6151
R1429 B.n482 B.n481 10.6151
R1430 B.n482 B.n95 10.6151
R1431 B.n486 B.n95 10.6151
R1432 B.n487 B.n486 10.6151
R1433 B.n488 B.n487 10.6151
R1434 B.n488 B.n93 10.6151
R1435 B.n492 B.n93 10.6151
R1436 B.n493 B.n492 10.6151
R1437 B.n494 B.n493 10.6151
R1438 B.n494 B.n91 10.6151
R1439 B.n498 B.n91 10.6151
R1440 B.n499 B.n498 10.6151
R1441 B.n500 B.n499 10.6151
R1442 B.n500 B.n89 10.6151
R1443 B.n504 B.n89 10.6151
R1444 B.n505 B.n504 10.6151
R1445 B.n506 B.n505 10.6151
R1446 B.n506 B.n87 10.6151
R1447 B.n510 B.n87 10.6151
R1448 B.n511 B.n510 10.6151
R1449 B.n512 B.n511 10.6151
R1450 B.n512 B.n85 10.6151
R1451 B.n516 B.n85 10.6151
R1452 B.n517 B.n516 10.6151
R1453 B.n518 B.n517 10.6151
R1454 B.n518 B.n83 10.6151
R1455 B.n522 B.n83 10.6151
R1456 B.n523 B.n522 10.6151
R1457 B.n524 B.n523 10.6151
R1458 B.n524 B.n81 10.6151
R1459 B.n528 B.n81 10.6151
R1460 B.n529 B.n528 10.6151
R1461 B.n530 B.n529 10.6151
R1462 B.n530 B.n79 10.6151
R1463 B.n534 B.n79 10.6151
R1464 B.n535 B.n534 10.6151
R1465 B.n536 B.n535 10.6151
R1466 B.n536 B.n77 10.6151
R1467 B.n540 B.n77 10.6151
R1468 B.n541 B.n540 10.6151
R1469 B.n542 B.n541 10.6151
R1470 B.n542 B.n75 10.6151
R1471 B.n546 B.n75 10.6151
R1472 B.n547 B.n546 10.6151
R1473 B.n548 B.n547 10.6151
R1474 B.n548 B.n73 10.6151
R1475 B.n552 B.n73 10.6151
R1476 B.n553 B.n552 10.6151
R1477 B.n554 B.n553 10.6151
R1478 B.n554 B.n71 10.6151
R1479 B.n558 B.n71 10.6151
R1480 B.n559 B.n558 10.6151
R1481 B.n560 B.n559 10.6151
R1482 B.n560 B.n69 10.6151
R1483 B.n564 B.n69 10.6151
R1484 B.n565 B.n564 10.6151
R1485 B.n566 B.n565 10.6151
R1486 B.n566 B.n67 10.6151
R1487 B.n570 B.n67 10.6151
R1488 B.n571 B.n570 10.6151
R1489 B.n572 B.n571 10.6151
R1490 B.n572 B.n65 10.6151
R1491 B.n576 B.n65 10.6151
R1492 B.n577 B.n576 10.6151
R1493 B.n578 B.n577 10.6151
R1494 B.n578 B.n63 10.6151
R1495 B.n582 B.n63 10.6151
R1496 B.n306 B.n159 10.6151
R1497 B.n307 B.n306 10.6151
R1498 B.n308 B.n307 10.6151
R1499 B.n308 B.n157 10.6151
R1500 B.n312 B.n157 10.6151
R1501 B.n313 B.n312 10.6151
R1502 B.n314 B.n313 10.6151
R1503 B.n314 B.n155 10.6151
R1504 B.n318 B.n155 10.6151
R1505 B.n319 B.n318 10.6151
R1506 B.n320 B.n319 10.6151
R1507 B.n320 B.n153 10.6151
R1508 B.n324 B.n153 10.6151
R1509 B.n327 B.n326 10.6151
R1510 B.n327 B.n149 10.6151
R1511 B.n331 B.n149 10.6151
R1512 B.n332 B.n331 10.6151
R1513 B.n333 B.n332 10.6151
R1514 B.n333 B.n147 10.6151
R1515 B.n337 B.n147 10.6151
R1516 B.n338 B.n337 10.6151
R1517 B.n339 B.n338 10.6151
R1518 B.n343 B.n342 10.6151
R1519 B.n344 B.n343 10.6151
R1520 B.n344 B.n141 10.6151
R1521 B.n348 B.n141 10.6151
R1522 B.n349 B.n348 10.6151
R1523 B.n350 B.n349 10.6151
R1524 B.n350 B.n139 10.6151
R1525 B.n354 B.n139 10.6151
R1526 B.n355 B.n354 10.6151
R1527 B.n356 B.n355 10.6151
R1528 B.n356 B.n137 10.6151
R1529 B.n360 B.n137 10.6151
R1530 B.n361 B.n360 10.6151
R1531 B.n302 B.n301 10.6151
R1532 B.n301 B.n300 10.6151
R1533 B.n300 B.n161 10.6151
R1534 B.n296 B.n161 10.6151
R1535 B.n296 B.n295 10.6151
R1536 B.n295 B.n294 10.6151
R1537 B.n294 B.n163 10.6151
R1538 B.n290 B.n163 10.6151
R1539 B.n290 B.n289 10.6151
R1540 B.n289 B.n288 10.6151
R1541 B.n288 B.n165 10.6151
R1542 B.n284 B.n165 10.6151
R1543 B.n284 B.n283 10.6151
R1544 B.n283 B.n282 10.6151
R1545 B.n282 B.n167 10.6151
R1546 B.n278 B.n167 10.6151
R1547 B.n278 B.n277 10.6151
R1548 B.n277 B.n276 10.6151
R1549 B.n276 B.n169 10.6151
R1550 B.n272 B.n169 10.6151
R1551 B.n272 B.n271 10.6151
R1552 B.n271 B.n270 10.6151
R1553 B.n270 B.n171 10.6151
R1554 B.n266 B.n171 10.6151
R1555 B.n266 B.n265 10.6151
R1556 B.n265 B.n264 10.6151
R1557 B.n264 B.n173 10.6151
R1558 B.n260 B.n173 10.6151
R1559 B.n260 B.n259 10.6151
R1560 B.n259 B.n258 10.6151
R1561 B.n258 B.n175 10.6151
R1562 B.n254 B.n175 10.6151
R1563 B.n254 B.n253 10.6151
R1564 B.n253 B.n252 10.6151
R1565 B.n252 B.n177 10.6151
R1566 B.n248 B.n177 10.6151
R1567 B.n248 B.n247 10.6151
R1568 B.n247 B.n246 10.6151
R1569 B.n246 B.n179 10.6151
R1570 B.n242 B.n179 10.6151
R1571 B.n242 B.n241 10.6151
R1572 B.n241 B.n240 10.6151
R1573 B.n240 B.n181 10.6151
R1574 B.n236 B.n181 10.6151
R1575 B.n236 B.n235 10.6151
R1576 B.n235 B.n234 10.6151
R1577 B.n234 B.n183 10.6151
R1578 B.n230 B.n183 10.6151
R1579 B.n230 B.n229 10.6151
R1580 B.n229 B.n228 10.6151
R1581 B.n228 B.n185 10.6151
R1582 B.n224 B.n185 10.6151
R1583 B.n224 B.n223 10.6151
R1584 B.n223 B.n222 10.6151
R1585 B.n222 B.n187 10.6151
R1586 B.n218 B.n187 10.6151
R1587 B.n218 B.n217 10.6151
R1588 B.n217 B.n216 10.6151
R1589 B.n216 B.n189 10.6151
R1590 B.n212 B.n189 10.6151
R1591 B.n212 B.n211 10.6151
R1592 B.n211 B.n210 10.6151
R1593 B.n210 B.n191 10.6151
R1594 B.n206 B.n191 10.6151
R1595 B.n206 B.n205 10.6151
R1596 B.n205 B.n204 10.6151
R1597 B.n204 B.n193 10.6151
R1598 B.n200 B.n193 10.6151
R1599 B.n200 B.n199 10.6151
R1600 B.n199 B.n198 10.6151
R1601 B.n198 B.n195 10.6151
R1602 B.n195 B.n0 10.6151
R1603 B.n747 B.n1 10.6151
R1604 B.n747 B.n746 10.6151
R1605 B.n746 B.n745 10.6151
R1606 B.n745 B.n4 10.6151
R1607 B.n741 B.n4 10.6151
R1608 B.n741 B.n740 10.6151
R1609 B.n740 B.n739 10.6151
R1610 B.n739 B.n6 10.6151
R1611 B.n735 B.n6 10.6151
R1612 B.n735 B.n734 10.6151
R1613 B.n734 B.n733 10.6151
R1614 B.n733 B.n8 10.6151
R1615 B.n729 B.n8 10.6151
R1616 B.n729 B.n728 10.6151
R1617 B.n728 B.n727 10.6151
R1618 B.n727 B.n10 10.6151
R1619 B.n723 B.n10 10.6151
R1620 B.n723 B.n722 10.6151
R1621 B.n722 B.n721 10.6151
R1622 B.n721 B.n12 10.6151
R1623 B.n717 B.n12 10.6151
R1624 B.n717 B.n716 10.6151
R1625 B.n716 B.n715 10.6151
R1626 B.n715 B.n14 10.6151
R1627 B.n711 B.n14 10.6151
R1628 B.n711 B.n710 10.6151
R1629 B.n710 B.n709 10.6151
R1630 B.n709 B.n16 10.6151
R1631 B.n705 B.n16 10.6151
R1632 B.n705 B.n704 10.6151
R1633 B.n704 B.n703 10.6151
R1634 B.n703 B.n18 10.6151
R1635 B.n699 B.n18 10.6151
R1636 B.n699 B.n698 10.6151
R1637 B.n698 B.n697 10.6151
R1638 B.n697 B.n20 10.6151
R1639 B.n693 B.n20 10.6151
R1640 B.n693 B.n692 10.6151
R1641 B.n692 B.n691 10.6151
R1642 B.n691 B.n22 10.6151
R1643 B.n687 B.n22 10.6151
R1644 B.n687 B.n686 10.6151
R1645 B.n686 B.n685 10.6151
R1646 B.n685 B.n24 10.6151
R1647 B.n681 B.n24 10.6151
R1648 B.n681 B.n680 10.6151
R1649 B.n680 B.n679 10.6151
R1650 B.n679 B.n26 10.6151
R1651 B.n675 B.n26 10.6151
R1652 B.n675 B.n674 10.6151
R1653 B.n674 B.n673 10.6151
R1654 B.n673 B.n28 10.6151
R1655 B.n669 B.n28 10.6151
R1656 B.n669 B.n668 10.6151
R1657 B.n668 B.n667 10.6151
R1658 B.n667 B.n30 10.6151
R1659 B.n663 B.n30 10.6151
R1660 B.n663 B.n662 10.6151
R1661 B.n662 B.n661 10.6151
R1662 B.n661 B.n32 10.6151
R1663 B.n657 B.n32 10.6151
R1664 B.n657 B.n656 10.6151
R1665 B.n656 B.n655 10.6151
R1666 B.n655 B.n34 10.6151
R1667 B.n651 B.n34 10.6151
R1668 B.n651 B.n650 10.6151
R1669 B.n650 B.n649 10.6151
R1670 B.n649 B.n36 10.6151
R1671 B.n645 B.n36 10.6151
R1672 B.n645 B.n644 10.6151
R1673 B.n644 B.n643 10.6151
R1674 B.n643 B.n38 10.6151
R1675 B.n620 B.n619 9.36635
R1676 B.n602 B.n56 9.36635
R1677 B.n325 B.n324 9.36635
R1678 B.n342 B.n145 9.36635
R1679 B.n751 B.n0 2.81026
R1680 B.n751 B.n1 2.81026
R1681 B.n619 B.n618 1.24928
R1682 B.n56 B.n52 1.24928
R1683 B.n326 B.n325 1.24928
R1684 B.n339 B.n145 1.24928
C0 VN w_n5398_n1500# 11.635099f
C1 VN VP 7.79359f
C2 VDD2 B 2.17395f
C3 VDD2 VDD1 2.6689f
C4 B VTAIL 1.75048f
C5 B w_n5398_n1500# 9.26553f
C6 VDD1 VTAIL 6.89695f
C7 VP B 2.59218f
C8 VDD1 w_n5398_n1500# 2.43279f
C9 VN B 1.40279f
C10 VP VDD1 3.42025f
C11 VDD2 VTAIL 6.95533f
C12 VN VDD1 0.161046f
C13 VDD2 w_n5398_n1500# 2.61525f
C14 VP VDD2 0.687102f
C15 VTAIL w_n5398_n1500# 2.01421f
C16 VN VDD2 2.89839f
C17 VP VTAIL 4.67357f
C18 VP w_n5398_n1500# 12.3373f
C19 VDD1 B 2.02613f
C20 VN VTAIL 4.65944f
C21 VDD2 VSUBS 2.409149f
C22 VDD1 VSUBS 2.096886f
C23 VTAIL VSUBS 0.687746f
C24 VN VSUBS 9.0365f
C25 VP VSUBS 4.502927f
C26 B VSUBS 5.167731f
C27 w_n5398_n1500# VSUBS 0.1028p
C28 B.n0 VSUBS 0.008558f
C29 B.n1 VSUBS 0.008558f
C30 B.n2 VSUBS 0.013533f
C31 B.n3 VSUBS 0.013533f
C32 B.n4 VSUBS 0.013533f
C33 B.n5 VSUBS 0.013533f
C34 B.n6 VSUBS 0.013533f
C35 B.n7 VSUBS 0.013533f
C36 B.n8 VSUBS 0.013533f
C37 B.n9 VSUBS 0.013533f
C38 B.n10 VSUBS 0.013533f
C39 B.n11 VSUBS 0.013533f
C40 B.n12 VSUBS 0.013533f
C41 B.n13 VSUBS 0.013533f
C42 B.n14 VSUBS 0.013533f
C43 B.n15 VSUBS 0.013533f
C44 B.n16 VSUBS 0.013533f
C45 B.n17 VSUBS 0.013533f
C46 B.n18 VSUBS 0.013533f
C47 B.n19 VSUBS 0.013533f
C48 B.n20 VSUBS 0.013533f
C49 B.n21 VSUBS 0.013533f
C50 B.n22 VSUBS 0.013533f
C51 B.n23 VSUBS 0.013533f
C52 B.n24 VSUBS 0.013533f
C53 B.n25 VSUBS 0.013533f
C54 B.n26 VSUBS 0.013533f
C55 B.n27 VSUBS 0.013533f
C56 B.n28 VSUBS 0.013533f
C57 B.n29 VSUBS 0.013533f
C58 B.n30 VSUBS 0.013533f
C59 B.n31 VSUBS 0.013533f
C60 B.n32 VSUBS 0.013533f
C61 B.n33 VSUBS 0.013533f
C62 B.n34 VSUBS 0.013533f
C63 B.n35 VSUBS 0.013533f
C64 B.n36 VSUBS 0.013533f
C65 B.n37 VSUBS 0.013533f
C66 B.n38 VSUBS 0.03154f
C67 B.n39 VSUBS 0.013533f
C68 B.n40 VSUBS 0.013533f
C69 B.n41 VSUBS 0.013533f
C70 B.n42 VSUBS 0.013533f
C71 B.n43 VSUBS 0.013533f
C72 B.n44 VSUBS 0.013533f
C73 B.n45 VSUBS 0.013533f
C74 B.t11 VSUBS 0.080166f
C75 B.t10 VSUBS 0.115746f
C76 B.t9 VSUBS 0.848322f
C77 B.n46 VSUBS 0.202087f
C78 B.n47 VSUBS 0.16792f
C79 B.n48 VSUBS 0.013533f
C80 B.n49 VSUBS 0.013533f
C81 B.n50 VSUBS 0.013533f
C82 B.n51 VSUBS 0.013533f
C83 B.n52 VSUBS 0.007563f
C84 B.n53 VSUBS 0.013533f
C85 B.t5 VSUBS 0.080166f
C86 B.t4 VSUBS 0.115747f
C87 B.t3 VSUBS 0.848322f
C88 B.n54 VSUBS 0.202086f
C89 B.n55 VSUBS 0.16792f
C90 B.n56 VSUBS 0.031355f
C91 B.n57 VSUBS 0.013533f
C92 B.n58 VSUBS 0.013533f
C93 B.n59 VSUBS 0.013533f
C94 B.n60 VSUBS 0.013533f
C95 B.n61 VSUBS 0.013533f
C96 B.n62 VSUBS 0.033739f
C97 B.n63 VSUBS 0.013533f
C98 B.n64 VSUBS 0.013533f
C99 B.n65 VSUBS 0.013533f
C100 B.n66 VSUBS 0.013533f
C101 B.n67 VSUBS 0.013533f
C102 B.n68 VSUBS 0.013533f
C103 B.n69 VSUBS 0.013533f
C104 B.n70 VSUBS 0.013533f
C105 B.n71 VSUBS 0.013533f
C106 B.n72 VSUBS 0.013533f
C107 B.n73 VSUBS 0.013533f
C108 B.n74 VSUBS 0.013533f
C109 B.n75 VSUBS 0.013533f
C110 B.n76 VSUBS 0.013533f
C111 B.n77 VSUBS 0.013533f
C112 B.n78 VSUBS 0.013533f
C113 B.n79 VSUBS 0.013533f
C114 B.n80 VSUBS 0.013533f
C115 B.n81 VSUBS 0.013533f
C116 B.n82 VSUBS 0.013533f
C117 B.n83 VSUBS 0.013533f
C118 B.n84 VSUBS 0.013533f
C119 B.n85 VSUBS 0.013533f
C120 B.n86 VSUBS 0.013533f
C121 B.n87 VSUBS 0.013533f
C122 B.n88 VSUBS 0.013533f
C123 B.n89 VSUBS 0.013533f
C124 B.n90 VSUBS 0.013533f
C125 B.n91 VSUBS 0.013533f
C126 B.n92 VSUBS 0.013533f
C127 B.n93 VSUBS 0.013533f
C128 B.n94 VSUBS 0.013533f
C129 B.n95 VSUBS 0.013533f
C130 B.n96 VSUBS 0.013533f
C131 B.n97 VSUBS 0.013533f
C132 B.n98 VSUBS 0.013533f
C133 B.n99 VSUBS 0.013533f
C134 B.n100 VSUBS 0.013533f
C135 B.n101 VSUBS 0.013533f
C136 B.n102 VSUBS 0.013533f
C137 B.n103 VSUBS 0.013533f
C138 B.n104 VSUBS 0.013533f
C139 B.n105 VSUBS 0.013533f
C140 B.n106 VSUBS 0.013533f
C141 B.n107 VSUBS 0.013533f
C142 B.n108 VSUBS 0.013533f
C143 B.n109 VSUBS 0.013533f
C144 B.n110 VSUBS 0.013533f
C145 B.n111 VSUBS 0.013533f
C146 B.n112 VSUBS 0.013533f
C147 B.n113 VSUBS 0.013533f
C148 B.n114 VSUBS 0.013533f
C149 B.n115 VSUBS 0.013533f
C150 B.n116 VSUBS 0.013533f
C151 B.n117 VSUBS 0.013533f
C152 B.n118 VSUBS 0.013533f
C153 B.n119 VSUBS 0.013533f
C154 B.n120 VSUBS 0.013533f
C155 B.n121 VSUBS 0.013533f
C156 B.n122 VSUBS 0.013533f
C157 B.n123 VSUBS 0.013533f
C158 B.n124 VSUBS 0.013533f
C159 B.n125 VSUBS 0.013533f
C160 B.n126 VSUBS 0.013533f
C161 B.n127 VSUBS 0.013533f
C162 B.n128 VSUBS 0.013533f
C163 B.n129 VSUBS 0.013533f
C164 B.n130 VSUBS 0.013533f
C165 B.n131 VSUBS 0.013533f
C166 B.n132 VSUBS 0.013533f
C167 B.n133 VSUBS 0.013533f
C168 B.n134 VSUBS 0.013533f
C169 B.n135 VSUBS 0.013533f
C170 B.n136 VSUBS 0.033739f
C171 B.n137 VSUBS 0.013533f
C172 B.n138 VSUBS 0.013533f
C173 B.n139 VSUBS 0.013533f
C174 B.n140 VSUBS 0.013533f
C175 B.n141 VSUBS 0.013533f
C176 B.n142 VSUBS 0.013533f
C177 B.t1 VSUBS 0.080166f
C178 B.t2 VSUBS 0.115747f
C179 B.t0 VSUBS 0.848322f
C180 B.n143 VSUBS 0.202086f
C181 B.n144 VSUBS 0.16792f
C182 B.n145 VSUBS 0.031355f
C183 B.n146 VSUBS 0.013533f
C184 B.n147 VSUBS 0.013533f
C185 B.n148 VSUBS 0.013533f
C186 B.n149 VSUBS 0.013533f
C187 B.n150 VSUBS 0.013533f
C188 B.t7 VSUBS 0.080166f
C189 B.t8 VSUBS 0.115746f
C190 B.t6 VSUBS 0.848322f
C191 B.n151 VSUBS 0.202087f
C192 B.n152 VSUBS 0.16792f
C193 B.n153 VSUBS 0.013533f
C194 B.n154 VSUBS 0.013533f
C195 B.n155 VSUBS 0.013533f
C196 B.n156 VSUBS 0.013533f
C197 B.n157 VSUBS 0.013533f
C198 B.n158 VSUBS 0.013533f
C199 B.n159 VSUBS 0.033739f
C200 B.n160 VSUBS 0.013533f
C201 B.n161 VSUBS 0.013533f
C202 B.n162 VSUBS 0.013533f
C203 B.n163 VSUBS 0.013533f
C204 B.n164 VSUBS 0.013533f
C205 B.n165 VSUBS 0.013533f
C206 B.n166 VSUBS 0.013533f
C207 B.n167 VSUBS 0.013533f
C208 B.n168 VSUBS 0.013533f
C209 B.n169 VSUBS 0.013533f
C210 B.n170 VSUBS 0.013533f
C211 B.n171 VSUBS 0.013533f
C212 B.n172 VSUBS 0.013533f
C213 B.n173 VSUBS 0.013533f
C214 B.n174 VSUBS 0.013533f
C215 B.n175 VSUBS 0.013533f
C216 B.n176 VSUBS 0.013533f
C217 B.n177 VSUBS 0.013533f
C218 B.n178 VSUBS 0.013533f
C219 B.n179 VSUBS 0.013533f
C220 B.n180 VSUBS 0.013533f
C221 B.n181 VSUBS 0.013533f
C222 B.n182 VSUBS 0.013533f
C223 B.n183 VSUBS 0.013533f
C224 B.n184 VSUBS 0.013533f
C225 B.n185 VSUBS 0.013533f
C226 B.n186 VSUBS 0.013533f
C227 B.n187 VSUBS 0.013533f
C228 B.n188 VSUBS 0.013533f
C229 B.n189 VSUBS 0.013533f
C230 B.n190 VSUBS 0.013533f
C231 B.n191 VSUBS 0.013533f
C232 B.n192 VSUBS 0.013533f
C233 B.n193 VSUBS 0.013533f
C234 B.n194 VSUBS 0.013533f
C235 B.n195 VSUBS 0.013533f
C236 B.n196 VSUBS 0.013533f
C237 B.n197 VSUBS 0.013533f
C238 B.n198 VSUBS 0.013533f
C239 B.n199 VSUBS 0.013533f
C240 B.n200 VSUBS 0.013533f
C241 B.n201 VSUBS 0.013533f
C242 B.n202 VSUBS 0.013533f
C243 B.n203 VSUBS 0.013533f
C244 B.n204 VSUBS 0.013533f
C245 B.n205 VSUBS 0.013533f
C246 B.n206 VSUBS 0.013533f
C247 B.n207 VSUBS 0.013533f
C248 B.n208 VSUBS 0.013533f
C249 B.n209 VSUBS 0.013533f
C250 B.n210 VSUBS 0.013533f
C251 B.n211 VSUBS 0.013533f
C252 B.n212 VSUBS 0.013533f
C253 B.n213 VSUBS 0.013533f
C254 B.n214 VSUBS 0.013533f
C255 B.n215 VSUBS 0.013533f
C256 B.n216 VSUBS 0.013533f
C257 B.n217 VSUBS 0.013533f
C258 B.n218 VSUBS 0.013533f
C259 B.n219 VSUBS 0.013533f
C260 B.n220 VSUBS 0.013533f
C261 B.n221 VSUBS 0.013533f
C262 B.n222 VSUBS 0.013533f
C263 B.n223 VSUBS 0.013533f
C264 B.n224 VSUBS 0.013533f
C265 B.n225 VSUBS 0.013533f
C266 B.n226 VSUBS 0.013533f
C267 B.n227 VSUBS 0.013533f
C268 B.n228 VSUBS 0.013533f
C269 B.n229 VSUBS 0.013533f
C270 B.n230 VSUBS 0.013533f
C271 B.n231 VSUBS 0.013533f
C272 B.n232 VSUBS 0.013533f
C273 B.n233 VSUBS 0.013533f
C274 B.n234 VSUBS 0.013533f
C275 B.n235 VSUBS 0.013533f
C276 B.n236 VSUBS 0.013533f
C277 B.n237 VSUBS 0.013533f
C278 B.n238 VSUBS 0.013533f
C279 B.n239 VSUBS 0.013533f
C280 B.n240 VSUBS 0.013533f
C281 B.n241 VSUBS 0.013533f
C282 B.n242 VSUBS 0.013533f
C283 B.n243 VSUBS 0.013533f
C284 B.n244 VSUBS 0.013533f
C285 B.n245 VSUBS 0.013533f
C286 B.n246 VSUBS 0.013533f
C287 B.n247 VSUBS 0.013533f
C288 B.n248 VSUBS 0.013533f
C289 B.n249 VSUBS 0.013533f
C290 B.n250 VSUBS 0.013533f
C291 B.n251 VSUBS 0.013533f
C292 B.n252 VSUBS 0.013533f
C293 B.n253 VSUBS 0.013533f
C294 B.n254 VSUBS 0.013533f
C295 B.n255 VSUBS 0.013533f
C296 B.n256 VSUBS 0.013533f
C297 B.n257 VSUBS 0.013533f
C298 B.n258 VSUBS 0.013533f
C299 B.n259 VSUBS 0.013533f
C300 B.n260 VSUBS 0.013533f
C301 B.n261 VSUBS 0.013533f
C302 B.n262 VSUBS 0.013533f
C303 B.n263 VSUBS 0.013533f
C304 B.n264 VSUBS 0.013533f
C305 B.n265 VSUBS 0.013533f
C306 B.n266 VSUBS 0.013533f
C307 B.n267 VSUBS 0.013533f
C308 B.n268 VSUBS 0.013533f
C309 B.n269 VSUBS 0.013533f
C310 B.n270 VSUBS 0.013533f
C311 B.n271 VSUBS 0.013533f
C312 B.n272 VSUBS 0.013533f
C313 B.n273 VSUBS 0.013533f
C314 B.n274 VSUBS 0.013533f
C315 B.n275 VSUBS 0.013533f
C316 B.n276 VSUBS 0.013533f
C317 B.n277 VSUBS 0.013533f
C318 B.n278 VSUBS 0.013533f
C319 B.n279 VSUBS 0.013533f
C320 B.n280 VSUBS 0.013533f
C321 B.n281 VSUBS 0.013533f
C322 B.n282 VSUBS 0.013533f
C323 B.n283 VSUBS 0.013533f
C324 B.n284 VSUBS 0.013533f
C325 B.n285 VSUBS 0.013533f
C326 B.n286 VSUBS 0.013533f
C327 B.n287 VSUBS 0.013533f
C328 B.n288 VSUBS 0.013533f
C329 B.n289 VSUBS 0.013533f
C330 B.n290 VSUBS 0.013533f
C331 B.n291 VSUBS 0.013533f
C332 B.n292 VSUBS 0.013533f
C333 B.n293 VSUBS 0.013533f
C334 B.n294 VSUBS 0.013533f
C335 B.n295 VSUBS 0.013533f
C336 B.n296 VSUBS 0.013533f
C337 B.n297 VSUBS 0.013533f
C338 B.n298 VSUBS 0.013533f
C339 B.n299 VSUBS 0.013533f
C340 B.n300 VSUBS 0.013533f
C341 B.n301 VSUBS 0.013533f
C342 B.n302 VSUBS 0.03154f
C343 B.n303 VSUBS 0.03154f
C344 B.n304 VSUBS 0.033739f
C345 B.n305 VSUBS 0.013533f
C346 B.n306 VSUBS 0.013533f
C347 B.n307 VSUBS 0.013533f
C348 B.n308 VSUBS 0.013533f
C349 B.n309 VSUBS 0.013533f
C350 B.n310 VSUBS 0.013533f
C351 B.n311 VSUBS 0.013533f
C352 B.n312 VSUBS 0.013533f
C353 B.n313 VSUBS 0.013533f
C354 B.n314 VSUBS 0.013533f
C355 B.n315 VSUBS 0.013533f
C356 B.n316 VSUBS 0.013533f
C357 B.n317 VSUBS 0.013533f
C358 B.n318 VSUBS 0.013533f
C359 B.n319 VSUBS 0.013533f
C360 B.n320 VSUBS 0.013533f
C361 B.n321 VSUBS 0.013533f
C362 B.n322 VSUBS 0.013533f
C363 B.n323 VSUBS 0.013533f
C364 B.n324 VSUBS 0.012737f
C365 B.n325 VSUBS 0.031355f
C366 B.n326 VSUBS 0.007563f
C367 B.n327 VSUBS 0.013533f
C368 B.n328 VSUBS 0.013533f
C369 B.n329 VSUBS 0.013533f
C370 B.n330 VSUBS 0.013533f
C371 B.n331 VSUBS 0.013533f
C372 B.n332 VSUBS 0.013533f
C373 B.n333 VSUBS 0.013533f
C374 B.n334 VSUBS 0.013533f
C375 B.n335 VSUBS 0.013533f
C376 B.n336 VSUBS 0.013533f
C377 B.n337 VSUBS 0.013533f
C378 B.n338 VSUBS 0.013533f
C379 B.n339 VSUBS 0.007563f
C380 B.n340 VSUBS 0.013533f
C381 B.n341 VSUBS 0.013533f
C382 B.n342 VSUBS 0.012737f
C383 B.n343 VSUBS 0.013533f
C384 B.n344 VSUBS 0.013533f
C385 B.n345 VSUBS 0.013533f
C386 B.n346 VSUBS 0.013533f
C387 B.n347 VSUBS 0.013533f
C388 B.n348 VSUBS 0.013533f
C389 B.n349 VSUBS 0.013533f
C390 B.n350 VSUBS 0.013533f
C391 B.n351 VSUBS 0.013533f
C392 B.n352 VSUBS 0.013533f
C393 B.n353 VSUBS 0.013533f
C394 B.n354 VSUBS 0.013533f
C395 B.n355 VSUBS 0.013533f
C396 B.n356 VSUBS 0.013533f
C397 B.n357 VSUBS 0.013533f
C398 B.n358 VSUBS 0.013533f
C399 B.n359 VSUBS 0.013533f
C400 B.n360 VSUBS 0.013533f
C401 B.n361 VSUBS 0.033739f
C402 B.n362 VSUBS 0.03154f
C403 B.n363 VSUBS 0.03154f
C404 B.n364 VSUBS 0.013533f
C405 B.n365 VSUBS 0.013533f
C406 B.n366 VSUBS 0.013533f
C407 B.n367 VSUBS 0.013533f
C408 B.n368 VSUBS 0.013533f
C409 B.n369 VSUBS 0.013533f
C410 B.n370 VSUBS 0.013533f
C411 B.n371 VSUBS 0.013533f
C412 B.n372 VSUBS 0.013533f
C413 B.n373 VSUBS 0.013533f
C414 B.n374 VSUBS 0.013533f
C415 B.n375 VSUBS 0.013533f
C416 B.n376 VSUBS 0.013533f
C417 B.n377 VSUBS 0.013533f
C418 B.n378 VSUBS 0.013533f
C419 B.n379 VSUBS 0.013533f
C420 B.n380 VSUBS 0.013533f
C421 B.n381 VSUBS 0.013533f
C422 B.n382 VSUBS 0.013533f
C423 B.n383 VSUBS 0.013533f
C424 B.n384 VSUBS 0.013533f
C425 B.n385 VSUBS 0.013533f
C426 B.n386 VSUBS 0.013533f
C427 B.n387 VSUBS 0.013533f
C428 B.n388 VSUBS 0.013533f
C429 B.n389 VSUBS 0.013533f
C430 B.n390 VSUBS 0.013533f
C431 B.n391 VSUBS 0.013533f
C432 B.n392 VSUBS 0.013533f
C433 B.n393 VSUBS 0.013533f
C434 B.n394 VSUBS 0.013533f
C435 B.n395 VSUBS 0.013533f
C436 B.n396 VSUBS 0.013533f
C437 B.n397 VSUBS 0.013533f
C438 B.n398 VSUBS 0.013533f
C439 B.n399 VSUBS 0.013533f
C440 B.n400 VSUBS 0.013533f
C441 B.n401 VSUBS 0.013533f
C442 B.n402 VSUBS 0.013533f
C443 B.n403 VSUBS 0.013533f
C444 B.n404 VSUBS 0.013533f
C445 B.n405 VSUBS 0.013533f
C446 B.n406 VSUBS 0.013533f
C447 B.n407 VSUBS 0.013533f
C448 B.n408 VSUBS 0.013533f
C449 B.n409 VSUBS 0.013533f
C450 B.n410 VSUBS 0.013533f
C451 B.n411 VSUBS 0.013533f
C452 B.n412 VSUBS 0.013533f
C453 B.n413 VSUBS 0.013533f
C454 B.n414 VSUBS 0.013533f
C455 B.n415 VSUBS 0.013533f
C456 B.n416 VSUBS 0.013533f
C457 B.n417 VSUBS 0.013533f
C458 B.n418 VSUBS 0.013533f
C459 B.n419 VSUBS 0.013533f
C460 B.n420 VSUBS 0.013533f
C461 B.n421 VSUBS 0.013533f
C462 B.n422 VSUBS 0.013533f
C463 B.n423 VSUBS 0.013533f
C464 B.n424 VSUBS 0.013533f
C465 B.n425 VSUBS 0.013533f
C466 B.n426 VSUBS 0.013533f
C467 B.n427 VSUBS 0.013533f
C468 B.n428 VSUBS 0.013533f
C469 B.n429 VSUBS 0.013533f
C470 B.n430 VSUBS 0.013533f
C471 B.n431 VSUBS 0.013533f
C472 B.n432 VSUBS 0.013533f
C473 B.n433 VSUBS 0.013533f
C474 B.n434 VSUBS 0.013533f
C475 B.n435 VSUBS 0.013533f
C476 B.n436 VSUBS 0.013533f
C477 B.n437 VSUBS 0.013533f
C478 B.n438 VSUBS 0.013533f
C479 B.n439 VSUBS 0.013533f
C480 B.n440 VSUBS 0.013533f
C481 B.n441 VSUBS 0.013533f
C482 B.n442 VSUBS 0.013533f
C483 B.n443 VSUBS 0.013533f
C484 B.n444 VSUBS 0.013533f
C485 B.n445 VSUBS 0.013533f
C486 B.n446 VSUBS 0.013533f
C487 B.n447 VSUBS 0.013533f
C488 B.n448 VSUBS 0.013533f
C489 B.n449 VSUBS 0.013533f
C490 B.n450 VSUBS 0.013533f
C491 B.n451 VSUBS 0.013533f
C492 B.n452 VSUBS 0.013533f
C493 B.n453 VSUBS 0.013533f
C494 B.n454 VSUBS 0.013533f
C495 B.n455 VSUBS 0.013533f
C496 B.n456 VSUBS 0.013533f
C497 B.n457 VSUBS 0.013533f
C498 B.n458 VSUBS 0.013533f
C499 B.n459 VSUBS 0.013533f
C500 B.n460 VSUBS 0.013533f
C501 B.n461 VSUBS 0.013533f
C502 B.n462 VSUBS 0.013533f
C503 B.n463 VSUBS 0.013533f
C504 B.n464 VSUBS 0.013533f
C505 B.n465 VSUBS 0.013533f
C506 B.n466 VSUBS 0.013533f
C507 B.n467 VSUBS 0.013533f
C508 B.n468 VSUBS 0.013533f
C509 B.n469 VSUBS 0.013533f
C510 B.n470 VSUBS 0.013533f
C511 B.n471 VSUBS 0.013533f
C512 B.n472 VSUBS 0.013533f
C513 B.n473 VSUBS 0.013533f
C514 B.n474 VSUBS 0.013533f
C515 B.n475 VSUBS 0.013533f
C516 B.n476 VSUBS 0.013533f
C517 B.n477 VSUBS 0.013533f
C518 B.n478 VSUBS 0.013533f
C519 B.n479 VSUBS 0.013533f
C520 B.n480 VSUBS 0.013533f
C521 B.n481 VSUBS 0.013533f
C522 B.n482 VSUBS 0.013533f
C523 B.n483 VSUBS 0.013533f
C524 B.n484 VSUBS 0.013533f
C525 B.n485 VSUBS 0.013533f
C526 B.n486 VSUBS 0.013533f
C527 B.n487 VSUBS 0.013533f
C528 B.n488 VSUBS 0.013533f
C529 B.n489 VSUBS 0.013533f
C530 B.n490 VSUBS 0.013533f
C531 B.n491 VSUBS 0.013533f
C532 B.n492 VSUBS 0.013533f
C533 B.n493 VSUBS 0.013533f
C534 B.n494 VSUBS 0.013533f
C535 B.n495 VSUBS 0.013533f
C536 B.n496 VSUBS 0.013533f
C537 B.n497 VSUBS 0.013533f
C538 B.n498 VSUBS 0.013533f
C539 B.n499 VSUBS 0.013533f
C540 B.n500 VSUBS 0.013533f
C541 B.n501 VSUBS 0.013533f
C542 B.n502 VSUBS 0.013533f
C543 B.n503 VSUBS 0.013533f
C544 B.n504 VSUBS 0.013533f
C545 B.n505 VSUBS 0.013533f
C546 B.n506 VSUBS 0.013533f
C547 B.n507 VSUBS 0.013533f
C548 B.n508 VSUBS 0.013533f
C549 B.n509 VSUBS 0.013533f
C550 B.n510 VSUBS 0.013533f
C551 B.n511 VSUBS 0.013533f
C552 B.n512 VSUBS 0.013533f
C553 B.n513 VSUBS 0.013533f
C554 B.n514 VSUBS 0.013533f
C555 B.n515 VSUBS 0.013533f
C556 B.n516 VSUBS 0.013533f
C557 B.n517 VSUBS 0.013533f
C558 B.n518 VSUBS 0.013533f
C559 B.n519 VSUBS 0.013533f
C560 B.n520 VSUBS 0.013533f
C561 B.n521 VSUBS 0.013533f
C562 B.n522 VSUBS 0.013533f
C563 B.n523 VSUBS 0.013533f
C564 B.n524 VSUBS 0.013533f
C565 B.n525 VSUBS 0.013533f
C566 B.n526 VSUBS 0.013533f
C567 B.n527 VSUBS 0.013533f
C568 B.n528 VSUBS 0.013533f
C569 B.n529 VSUBS 0.013533f
C570 B.n530 VSUBS 0.013533f
C571 B.n531 VSUBS 0.013533f
C572 B.n532 VSUBS 0.013533f
C573 B.n533 VSUBS 0.013533f
C574 B.n534 VSUBS 0.013533f
C575 B.n535 VSUBS 0.013533f
C576 B.n536 VSUBS 0.013533f
C577 B.n537 VSUBS 0.013533f
C578 B.n538 VSUBS 0.013533f
C579 B.n539 VSUBS 0.013533f
C580 B.n540 VSUBS 0.013533f
C581 B.n541 VSUBS 0.013533f
C582 B.n542 VSUBS 0.013533f
C583 B.n543 VSUBS 0.013533f
C584 B.n544 VSUBS 0.013533f
C585 B.n545 VSUBS 0.013533f
C586 B.n546 VSUBS 0.013533f
C587 B.n547 VSUBS 0.013533f
C588 B.n548 VSUBS 0.013533f
C589 B.n549 VSUBS 0.013533f
C590 B.n550 VSUBS 0.013533f
C591 B.n551 VSUBS 0.013533f
C592 B.n552 VSUBS 0.013533f
C593 B.n553 VSUBS 0.013533f
C594 B.n554 VSUBS 0.013533f
C595 B.n555 VSUBS 0.013533f
C596 B.n556 VSUBS 0.013533f
C597 B.n557 VSUBS 0.013533f
C598 B.n558 VSUBS 0.013533f
C599 B.n559 VSUBS 0.013533f
C600 B.n560 VSUBS 0.013533f
C601 B.n561 VSUBS 0.013533f
C602 B.n562 VSUBS 0.013533f
C603 B.n563 VSUBS 0.013533f
C604 B.n564 VSUBS 0.013533f
C605 B.n565 VSUBS 0.013533f
C606 B.n566 VSUBS 0.013533f
C607 B.n567 VSUBS 0.013533f
C608 B.n568 VSUBS 0.013533f
C609 B.n569 VSUBS 0.013533f
C610 B.n570 VSUBS 0.013533f
C611 B.n571 VSUBS 0.013533f
C612 B.n572 VSUBS 0.013533f
C613 B.n573 VSUBS 0.013533f
C614 B.n574 VSUBS 0.013533f
C615 B.n575 VSUBS 0.013533f
C616 B.n576 VSUBS 0.013533f
C617 B.n577 VSUBS 0.013533f
C618 B.n578 VSUBS 0.013533f
C619 B.n579 VSUBS 0.013533f
C620 B.n580 VSUBS 0.013533f
C621 B.n581 VSUBS 0.03154f
C622 B.n582 VSUBS 0.033068f
C623 B.n583 VSUBS 0.032211f
C624 B.n584 VSUBS 0.013533f
C625 B.n585 VSUBS 0.013533f
C626 B.n586 VSUBS 0.013533f
C627 B.n587 VSUBS 0.013533f
C628 B.n588 VSUBS 0.013533f
C629 B.n589 VSUBS 0.013533f
C630 B.n590 VSUBS 0.013533f
C631 B.n591 VSUBS 0.013533f
C632 B.n592 VSUBS 0.013533f
C633 B.n593 VSUBS 0.013533f
C634 B.n594 VSUBS 0.013533f
C635 B.n595 VSUBS 0.013533f
C636 B.n596 VSUBS 0.013533f
C637 B.n597 VSUBS 0.013533f
C638 B.n598 VSUBS 0.013533f
C639 B.n599 VSUBS 0.013533f
C640 B.n600 VSUBS 0.013533f
C641 B.n601 VSUBS 0.013533f
C642 B.n602 VSUBS 0.012737f
C643 B.n603 VSUBS 0.013533f
C644 B.n604 VSUBS 0.013533f
C645 B.n605 VSUBS 0.013533f
C646 B.n606 VSUBS 0.013533f
C647 B.n607 VSUBS 0.013533f
C648 B.n608 VSUBS 0.013533f
C649 B.n609 VSUBS 0.013533f
C650 B.n610 VSUBS 0.013533f
C651 B.n611 VSUBS 0.013533f
C652 B.n612 VSUBS 0.013533f
C653 B.n613 VSUBS 0.013533f
C654 B.n614 VSUBS 0.013533f
C655 B.n615 VSUBS 0.013533f
C656 B.n616 VSUBS 0.013533f
C657 B.n617 VSUBS 0.013533f
C658 B.n618 VSUBS 0.007563f
C659 B.n619 VSUBS 0.031355f
C660 B.n620 VSUBS 0.012737f
C661 B.n621 VSUBS 0.013533f
C662 B.n622 VSUBS 0.013533f
C663 B.n623 VSUBS 0.013533f
C664 B.n624 VSUBS 0.013533f
C665 B.n625 VSUBS 0.013533f
C666 B.n626 VSUBS 0.013533f
C667 B.n627 VSUBS 0.013533f
C668 B.n628 VSUBS 0.013533f
C669 B.n629 VSUBS 0.013533f
C670 B.n630 VSUBS 0.013533f
C671 B.n631 VSUBS 0.013533f
C672 B.n632 VSUBS 0.013533f
C673 B.n633 VSUBS 0.013533f
C674 B.n634 VSUBS 0.013533f
C675 B.n635 VSUBS 0.013533f
C676 B.n636 VSUBS 0.013533f
C677 B.n637 VSUBS 0.013533f
C678 B.n638 VSUBS 0.013533f
C679 B.n639 VSUBS 0.033739f
C680 B.n640 VSUBS 0.033739f
C681 B.n641 VSUBS 0.03154f
C682 B.n642 VSUBS 0.013533f
C683 B.n643 VSUBS 0.013533f
C684 B.n644 VSUBS 0.013533f
C685 B.n645 VSUBS 0.013533f
C686 B.n646 VSUBS 0.013533f
C687 B.n647 VSUBS 0.013533f
C688 B.n648 VSUBS 0.013533f
C689 B.n649 VSUBS 0.013533f
C690 B.n650 VSUBS 0.013533f
C691 B.n651 VSUBS 0.013533f
C692 B.n652 VSUBS 0.013533f
C693 B.n653 VSUBS 0.013533f
C694 B.n654 VSUBS 0.013533f
C695 B.n655 VSUBS 0.013533f
C696 B.n656 VSUBS 0.013533f
C697 B.n657 VSUBS 0.013533f
C698 B.n658 VSUBS 0.013533f
C699 B.n659 VSUBS 0.013533f
C700 B.n660 VSUBS 0.013533f
C701 B.n661 VSUBS 0.013533f
C702 B.n662 VSUBS 0.013533f
C703 B.n663 VSUBS 0.013533f
C704 B.n664 VSUBS 0.013533f
C705 B.n665 VSUBS 0.013533f
C706 B.n666 VSUBS 0.013533f
C707 B.n667 VSUBS 0.013533f
C708 B.n668 VSUBS 0.013533f
C709 B.n669 VSUBS 0.013533f
C710 B.n670 VSUBS 0.013533f
C711 B.n671 VSUBS 0.013533f
C712 B.n672 VSUBS 0.013533f
C713 B.n673 VSUBS 0.013533f
C714 B.n674 VSUBS 0.013533f
C715 B.n675 VSUBS 0.013533f
C716 B.n676 VSUBS 0.013533f
C717 B.n677 VSUBS 0.013533f
C718 B.n678 VSUBS 0.013533f
C719 B.n679 VSUBS 0.013533f
C720 B.n680 VSUBS 0.013533f
C721 B.n681 VSUBS 0.013533f
C722 B.n682 VSUBS 0.013533f
C723 B.n683 VSUBS 0.013533f
C724 B.n684 VSUBS 0.013533f
C725 B.n685 VSUBS 0.013533f
C726 B.n686 VSUBS 0.013533f
C727 B.n687 VSUBS 0.013533f
C728 B.n688 VSUBS 0.013533f
C729 B.n689 VSUBS 0.013533f
C730 B.n690 VSUBS 0.013533f
C731 B.n691 VSUBS 0.013533f
C732 B.n692 VSUBS 0.013533f
C733 B.n693 VSUBS 0.013533f
C734 B.n694 VSUBS 0.013533f
C735 B.n695 VSUBS 0.013533f
C736 B.n696 VSUBS 0.013533f
C737 B.n697 VSUBS 0.013533f
C738 B.n698 VSUBS 0.013533f
C739 B.n699 VSUBS 0.013533f
C740 B.n700 VSUBS 0.013533f
C741 B.n701 VSUBS 0.013533f
C742 B.n702 VSUBS 0.013533f
C743 B.n703 VSUBS 0.013533f
C744 B.n704 VSUBS 0.013533f
C745 B.n705 VSUBS 0.013533f
C746 B.n706 VSUBS 0.013533f
C747 B.n707 VSUBS 0.013533f
C748 B.n708 VSUBS 0.013533f
C749 B.n709 VSUBS 0.013533f
C750 B.n710 VSUBS 0.013533f
C751 B.n711 VSUBS 0.013533f
C752 B.n712 VSUBS 0.013533f
C753 B.n713 VSUBS 0.013533f
C754 B.n714 VSUBS 0.013533f
C755 B.n715 VSUBS 0.013533f
C756 B.n716 VSUBS 0.013533f
C757 B.n717 VSUBS 0.013533f
C758 B.n718 VSUBS 0.013533f
C759 B.n719 VSUBS 0.013533f
C760 B.n720 VSUBS 0.013533f
C761 B.n721 VSUBS 0.013533f
C762 B.n722 VSUBS 0.013533f
C763 B.n723 VSUBS 0.013533f
C764 B.n724 VSUBS 0.013533f
C765 B.n725 VSUBS 0.013533f
C766 B.n726 VSUBS 0.013533f
C767 B.n727 VSUBS 0.013533f
C768 B.n728 VSUBS 0.013533f
C769 B.n729 VSUBS 0.013533f
C770 B.n730 VSUBS 0.013533f
C771 B.n731 VSUBS 0.013533f
C772 B.n732 VSUBS 0.013533f
C773 B.n733 VSUBS 0.013533f
C774 B.n734 VSUBS 0.013533f
C775 B.n735 VSUBS 0.013533f
C776 B.n736 VSUBS 0.013533f
C777 B.n737 VSUBS 0.013533f
C778 B.n738 VSUBS 0.013533f
C779 B.n739 VSUBS 0.013533f
C780 B.n740 VSUBS 0.013533f
C781 B.n741 VSUBS 0.013533f
C782 B.n742 VSUBS 0.013533f
C783 B.n743 VSUBS 0.013533f
C784 B.n744 VSUBS 0.013533f
C785 B.n745 VSUBS 0.013533f
C786 B.n746 VSUBS 0.013533f
C787 B.n747 VSUBS 0.013533f
C788 B.n748 VSUBS 0.013533f
C789 B.n749 VSUBS 0.013533f
C790 B.n750 VSUBS 0.013533f
C791 B.n751 VSUBS 0.030644f
C792 VDD2.n0 VSUBS 0.045632f
C793 VDD2.n1 VSUBS 0.329762f
C794 VDD2.n2 VSUBS 0.021892f
C795 VDD2.t3 VSUBS 0.120706f
C796 VDD2.n3 VSUBS 0.145222f
C797 VDD2.n4 VSUBS 0.036696f
C798 VDD2.n5 VSUBS 0.03881f
C799 VDD2.n6 VSUBS 0.128221f
C800 VDD2.n7 VSUBS 0.02318f
C801 VDD2.n8 VSUBS 0.021892f
C802 VDD2.n9 VSUBS 0.088605f
C803 VDD2.n10 VSUBS 0.123905f
C804 VDD2.t4 VSUBS 0.085638f
C805 VDD2.t8 VSUBS 0.085638f
C806 VDD2.n11 VSUBS 0.409276f
C807 VDD2.n12 VSUBS 1.48683f
C808 VDD2.t1 VSUBS 0.085638f
C809 VDD2.t5 VSUBS 0.085638f
C810 VDD2.n13 VSUBS 0.428245f
C811 VDD2.n14 VSUBS 4.64773f
C812 VDD2.n15 VSUBS 0.045632f
C813 VDD2.n16 VSUBS 0.329762f
C814 VDD2.n17 VSUBS 0.021892f
C815 VDD2.t6 VSUBS 0.120706f
C816 VDD2.n18 VSUBS 0.145222f
C817 VDD2.n19 VSUBS 0.036696f
C818 VDD2.n20 VSUBS 0.03881f
C819 VDD2.n21 VSUBS 0.128221f
C820 VDD2.n22 VSUBS 0.02318f
C821 VDD2.n23 VSUBS 0.021892f
C822 VDD2.n24 VSUBS 0.088605f
C823 VDD2.n25 VSUBS 0.092614f
C824 VDD2.n26 VSUBS 4.0012f
C825 VDD2.t9 VSUBS 0.085638f
C826 VDD2.t2 VSUBS 0.085638f
C827 VDD2.n27 VSUBS 0.409277f
C828 VDD2.n28 VSUBS 1.03889f
C829 VDD2.t0 VSUBS 0.085638f
C830 VDD2.t7 VSUBS 0.085638f
C831 VDD2.n29 VSUBS 0.428212f
C832 VN.t4 VSUBS 0.968584f
C833 VN.n0 VSUBS 0.563985f
C834 VN.n1 VSUBS 0.04421f
C835 VN.n2 VSUBS 0.059985f
C836 VN.n3 VSUBS 0.04421f
C837 VN.n4 VSUBS 0.046367f
C838 VN.n5 VSUBS 0.04421f
C839 VN.n6 VSUBS 0.041069f
C840 VN.n7 VSUBS 0.04421f
C841 VN.t1 VSUBS 0.968584f
C842 VN.n8 VSUBS 0.40959f
C843 VN.n9 VSUBS 0.04421f
C844 VN.n10 VSUBS 0.041069f
C845 VN.n11 VSUBS 0.04421f
C846 VN.t5 VSUBS 0.968584f
C847 VN.n12 VSUBS 0.57535f
C848 VN.t6 VSUBS 1.42887f
C849 VN.n13 VSUBS 0.576688f
C850 VN.n14 VSUBS 0.540658f
C851 VN.n15 VSUBS 0.077127f
C852 VN.n16 VSUBS 0.081984f
C853 VN.n17 VSUBS 0.081165f
C854 VN.n18 VSUBS 0.04421f
C855 VN.n19 VSUBS 0.04421f
C856 VN.n20 VSUBS 0.04421f
C857 VN.n21 VSUBS 0.088283f
C858 VN.n22 VSUBS 0.081984f
C859 VN.n23 VSUBS 0.061747f
C860 VN.n24 VSUBS 0.04421f
C861 VN.n25 VSUBS 0.04421f
C862 VN.n26 VSUBS 0.061747f
C863 VN.n27 VSUBS 0.081984f
C864 VN.n28 VSUBS 0.088283f
C865 VN.n29 VSUBS 0.04421f
C866 VN.n30 VSUBS 0.04421f
C867 VN.n31 VSUBS 0.04421f
C868 VN.n32 VSUBS 0.081165f
C869 VN.n33 VSUBS 0.081984f
C870 VN.t8 VSUBS 0.968584f
C871 VN.n34 VSUBS 0.40959f
C872 VN.n35 VSUBS 0.077127f
C873 VN.n36 VSUBS 0.04421f
C874 VN.n37 VSUBS 0.04421f
C875 VN.n38 VSUBS 0.04421f
C876 VN.n39 VSUBS 0.081984f
C877 VN.n40 VSUBS 0.081984f
C878 VN.n41 VSUBS 0.068548f
C879 VN.n42 VSUBS 0.04421f
C880 VN.n43 VSUBS 0.04421f
C881 VN.n44 VSUBS 0.04421f
C882 VN.n45 VSUBS 0.081984f
C883 VN.n46 VSUBS 0.081984f
C884 VN.n47 VSUBS 0.052034f
C885 VN.n48 VSUBS 0.071343f
C886 VN.n49 VSUBS 0.120699f
C887 VN.t3 VSUBS 0.968584f
C888 VN.n50 VSUBS 0.563985f
C889 VN.n51 VSUBS 0.04421f
C890 VN.n52 VSUBS 0.059985f
C891 VN.n53 VSUBS 0.04421f
C892 VN.n54 VSUBS 0.046367f
C893 VN.n55 VSUBS 0.04421f
C894 VN.t0 VSUBS 0.968584f
C895 VN.n56 VSUBS 0.40959f
C896 VN.n57 VSUBS 0.041069f
C897 VN.n58 VSUBS 0.04421f
C898 VN.t7 VSUBS 0.968584f
C899 VN.n59 VSUBS 0.40959f
C900 VN.n60 VSUBS 0.04421f
C901 VN.n61 VSUBS 0.041069f
C902 VN.n62 VSUBS 0.04421f
C903 VN.t9 VSUBS 0.968584f
C904 VN.n63 VSUBS 0.57535f
C905 VN.t2 VSUBS 1.42887f
C906 VN.n64 VSUBS 0.576688f
C907 VN.n65 VSUBS 0.540658f
C908 VN.n66 VSUBS 0.077127f
C909 VN.n67 VSUBS 0.081984f
C910 VN.n68 VSUBS 0.081165f
C911 VN.n69 VSUBS 0.04421f
C912 VN.n70 VSUBS 0.04421f
C913 VN.n71 VSUBS 0.04421f
C914 VN.n72 VSUBS 0.088283f
C915 VN.n73 VSUBS 0.081984f
C916 VN.n74 VSUBS 0.061747f
C917 VN.n75 VSUBS 0.04421f
C918 VN.n76 VSUBS 0.04421f
C919 VN.n77 VSUBS 0.061747f
C920 VN.n78 VSUBS 0.081984f
C921 VN.n79 VSUBS 0.088283f
C922 VN.n80 VSUBS 0.04421f
C923 VN.n81 VSUBS 0.04421f
C924 VN.n82 VSUBS 0.04421f
C925 VN.n83 VSUBS 0.081165f
C926 VN.n84 VSUBS 0.081984f
C927 VN.n85 VSUBS 0.077127f
C928 VN.n86 VSUBS 0.04421f
C929 VN.n87 VSUBS 0.04421f
C930 VN.n88 VSUBS 0.04421f
C931 VN.n89 VSUBS 0.081984f
C932 VN.n90 VSUBS 0.081984f
C933 VN.n91 VSUBS 0.068548f
C934 VN.n92 VSUBS 0.04421f
C935 VN.n93 VSUBS 0.04421f
C936 VN.n94 VSUBS 0.04421f
C937 VN.n95 VSUBS 0.081984f
C938 VN.n96 VSUBS 0.081984f
C939 VN.n97 VSUBS 0.052034f
C940 VN.n98 VSUBS 0.071343f
C941 VN.n99 VSUBS 2.55492f
C942 VDD1.n0 VSUBS 0.04524f
C943 VDD1.n1 VSUBS 0.326935f
C944 VDD1.n2 VSUBS 0.021705f
C945 VDD1.t7 VSUBS 0.119671f
C946 VDD1.n3 VSUBS 0.143977f
C947 VDD1.n4 VSUBS 0.036381f
C948 VDD1.n5 VSUBS 0.038477f
C949 VDD1.n6 VSUBS 0.127121f
C950 VDD1.n7 VSUBS 0.022982f
C951 VDD1.n8 VSUBS 0.021705f
C952 VDD1.n9 VSUBS 0.087846f
C953 VDD1.n10 VSUBS 0.122842f
C954 VDD1.t1 VSUBS 0.084904f
C955 VDD1.t9 VSUBS 0.084904f
C956 VDD1.n11 VSUBS 0.405768f
C957 VDD1.n12 VSUBS 1.48759f
C958 VDD1.n13 VSUBS 0.04524f
C959 VDD1.n14 VSUBS 0.326935f
C960 VDD1.n15 VSUBS 0.021705f
C961 VDD1.t5 VSUBS 0.119671f
C962 VDD1.n16 VSUBS 0.143977f
C963 VDD1.n17 VSUBS 0.036381f
C964 VDD1.n18 VSUBS 0.038477f
C965 VDD1.n19 VSUBS 0.127121f
C966 VDD1.n20 VSUBS 0.022982f
C967 VDD1.n21 VSUBS 0.021705f
C968 VDD1.n22 VSUBS 0.087846f
C969 VDD1.n23 VSUBS 0.122842f
C970 VDD1.t4 VSUBS 0.084904f
C971 VDD1.t2 VSUBS 0.084904f
C972 VDD1.n24 VSUBS 0.405767f
C973 VDD1.n25 VSUBS 1.47408f
C974 VDD1.t6 VSUBS 0.084904f
C975 VDD1.t0 VSUBS 0.084904f
C976 VDD1.n26 VSUBS 0.424573f
C977 VDD1.n27 VSUBS 4.82869f
C978 VDD1.t3 VSUBS 0.084904f
C979 VDD1.t8 VSUBS 0.084904f
C980 VDD1.n28 VSUBS 0.405768f
C981 VDD1.n29 VSUBS 4.64474f
C982 VTAIL.t5 VSUBS 0.082229f
C983 VTAIL.t4 VSUBS 0.082229f
C984 VTAIL.n0 VSUBS 0.333272f
C985 VTAIL.n1 VSUBS 1.06328f
C986 VTAIL.n2 VSUBS 0.043815f
C987 VTAIL.n3 VSUBS 0.316632f
C988 VTAIL.n4 VSUBS 0.021021f
C989 VTAIL.t6 VSUBS 0.115899f
C990 VTAIL.n5 VSUBS 0.139439f
C991 VTAIL.n6 VSUBS 0.035235f
C992 VTAIL.n7 VSUBS 0.037264f
C993 VTAIL.n8 VSUBS 0.123115f
C994 VTAIL.n9 VSUBS 0.022257f
C995 VTAIL.n10 VSUBS 0.021021f
C996 VTAIL.n11 VSUBS 0.085078f
C997 VTAIL.n12 VSUBS 0.06187f
C998 VTAIL.n13 VSUBS 0.691075f
C999 VTAIL.t11 VSUBS 0.082229f
C1000 VTAIL.t10 VSUBS 0.082229f
C1001 VTAIL.n14 VSUBS 0.333272f
C1002 VTAIL.n15 VSUBS 1.29745f
C1003 VTAIL.t8 VSUBS 0.082229f
C1004 VTAIL.t7 VSUBS 0.082229f
C1005 VTAIL.n16 VSUBS 0.333272f
C1006 VTAIL.n17 VSUBS 2.51885f
C1007 VTAIL.t18 VSUBS 0.082229f
C1008 VTAIL.t3 VSUBS 0.082229f
C1009 VTAIL.n18 VSUBS 0.333274f
C1010 VTAIL.n19 VSUBS 2.51885f
C1011 VTAIL.t16 VSUBS 0.082229f
C1012 VTAIL.t1 VSUBS 0.082229f
C1013 VTAIL.n20 VSUBS 0.333274f
C1014 VTAIL.n21 VSUBS 1.29745f
C1015 VTAIL.n22 VSUBS 0.043815f
C1016 VTAIL.n23 VSUBS 0.316632f
C1017 VTAIL.n24 VSUBS 0.021021f
C1018 VTAIL.t2 VSUBS 0.115899f
C1019 VTAIL.n25 VSUBS 0.139439f
C1020 VTAIL.n26 VSUBS 0.035235f
C1021 VTAIL.n27 VSUBS 0.037264f
C1022 VTAIL.n28 VSUBS 0.123115f
C1023 VTAIL.n29 VSUBS 0.022257f
C1024 VTAIL.n30 VSUBS 0.021021f
C1025 VTAIL.n31 VSUBS 0.085078f
C1026 VTAIL.n32 VSUBS 0.06187f
C1027 VTAIL.n33 VSUBS 0.691075f
C1028 VTAIL.t9 VSUBS 0.082229f
C1029 VTAIL.t15 VSUBS 0.082229f
C1030 VTAIL.n34 VSUBS 0.333274f
C1031 VTAIL.n35 VSUBS 1.15619f
C1032 VTAIL.t14 VSUBS 0.082229f
C1033 VTAIL.t12 VSUBS 0.082229f
C1034 VTAIL.n36 VSUBS 0.333274f
C1035 VTAIL.n37 VSUBS 1.29745f
C1036 VTAIL.n38 VSUBS 0.043815f
C1037 VTAIL.n39 VSUBS 0.316632f
C1038 VTAIL.n40 VSUBS 0.021021f
C1039 VTAIL.t13 VSUBS 0.115899f
C1040 VTAIL.n41 VSUBS 0.139439f
C1041 VTAIL.n42 VSUBS 0.035235f
C1042 VTAIL.n43 VSUBS 0.037264f
C1043 VTAIL.n44 VSUBS 0.123115f
C1044 VTAIL.n45 VSUBS 0.022257f
C1045 VTAIL.n46 VSUBS 0.021021f
C1046 VTAIL.n47 VSUBS 0.085078f
C1047 VTAIL.n48 VSUBS 0.06187f
C1048 VTAIL.n49 VSUBS 1.65277f
C1049 VTAIL.n50 VSUBS 0.043815f
C1050 VTAIL.n51 VSUBS 0.316632f
C1051 VTAIL.n52 VSUBS 0.021021f
C1052 VTAIL.t17 VSUBS 0.115899f
C1053 VTAIL.n53 VSUBS 0.139439f
C1054 VTAIL.n54 VSUBS 0.035235f
C1055 VTAIL.n55 VSUBS 0.037264f
C1056 VTAIL.n56 VSUBS 0.123115f
C1057 VTAIL.n57 VSUBS 0.022257f
C1058 VTAIL.n58 VSUBS 0.021021f
C1059 VTAIL.n59 VSUBS 0.085078f
C1060 VTAIL.n60 VSUBS 0.06187f
C1061 VTAIL.n61 VSUBS 1.65277f
C1062 VTAIL.t19 VSUBS 0.082229f
C1063 VTAIL.t0 VSUBS 0.082229f
C1064 VTAIL.n62 VSUBS 0.333272f
C1065 VTAIL.n63 VSUBS 0.989391f
C1066 VP.t9 VSUBS 1.10745f
C1067 VP.n0 VSUBS 0.644845f
C1068 VP.n1 VSUBS 0.050549f
C1069 VP.n2 VSUBS 0.068586f
C1070 VP.n3 VSUBS 0.050549f
C1071 VP.n4 VSUBS 0.053015f
C1072 VP.n5 VSUBS 0.050549f
C1073 VP.n6 VSUBS 0.046958f
C1074 VP.n7 VSUBS 0.050549f
C1075 VP.t7 VSUBS 1.10745f
C1076 VP.n8 VSUBS 0.468314f
C1077 VP.n9 VSUBS 0.050549f
C1078 VP.n10 VSUBS 0.046958f
C1079 VP.n11 VSUBS 0.050549f
C1080 VP.t5 VSUBS 1.10745f
C1081 VP.n12 VSUBS 0.468314f
C1082 VP.n13 VSUBS 0.050549f
C1083 VP.n14 VSUBS 0.078375f
C1084 VP.n15 VSUBS 0.050549f
C1085 VP.n16 VSUBS 0.059494f
C1086 VP.t1 VSUBS 1.10745f
C1087 VP.n17 VSUBS 0.644845f
C1088 VP.n18 VSUBS 0.050549f
C1089 VP.n19 VSUBS 0.068586f
C1090 VP.n20 VSUBS 0.050549f
C1091 VP.n21 VSUBS 0.053015f
C1092 VP.n22 VSUBS 0.050549f
C1093 VP.n23 VSUBS 0.046958f
C1094 VP.n24 VSUBS 0.050549f
C1095 VP.t0 VSUBS 1.10745f
C1096 VP.n25 VSUBS 0.468314f
C1097 VP.n26 VSUBS 0.050549f
C1098 VP.n27 VSUBS 0.046958f
C1099 VP.n28 VSUBS 0.050549f
C1100 VP.t8 VSUBS 1.10745f
C1101 VP.n29 VSUBS 0.657839f
C1102 VP.t2 VSUBS 1.63373f
C1103 VP.n30 VSUBS 0.65937f
C1104 VP.n31 VSUBS 0.618174f
C1105 VP.n32 VSUBS 0.088185f
C1106 VP.n33 VSUBS 0.093738f
C1107 VP.n34 VSUBS 0.092801f
C1108 VP.n35 VSUBS 0.050549f
C1109 VP.n36 VSUBS 0.050549f
C1110 VP.n37 VSUBS 0.050549f
C1111 VP.n38 VSUBS 0.10094f
C1112 VP.n39 VSUBS 0.093738f
C1113 VP.n40 VSUBS 0.0706f
C1114 VP.n41 VSUBS 0.050549f
C1115 VP.n42 VSUBS 0.050549f
C1116 VP.n43 VSUBS 0.0706f
C1117 VP.n44 VSUBS 0.093738f
C1118 VP.n45 VSUBS 0.10094f
C1119 VP.n46 VSUBS 0.050549f
C1120 VP.n47 VSUBS 0.050549f
C1121 VP.n48 VSUBS 0.050549f
C1122 VP.n49 VSUBS 0.092801f
C1123 VP.n50 VSUBS 0.093738f
C1124 VP.t6 VSUBS 1.10745f
C1125 VP.n51 VSUBS 0.468314f
C1126 VP.n52 VSUBS 0.088185f
C1127 VP.n53 VSUBS 0.050549f
C1128 VP.n54 VSUBS 0.050549f
C1129 VP.n55 VSUBS 0.050549f
C1130 VP.n56 VSUBS 0.093738f
C1131 VP.n57 VSUBS 0.093738f
C1132 VP.n58 VSUBS 0.078375f
C1133 VP.n59 VSUBS 0.050549f
C1134 VP.n60 VSUBS 0.050549f
C1135 VP.n61 VSUBS 0.050549f
C1136 VP.n62 VSUBS 0.093738f
C1137 VP.n63 VSUBS 0.093738f
C1138 VP.n64 VSUBS 0.059494f
C1139 VP.n65 VSUBS 0.081572f
C1140 VP.n66 VSUBS 2.90055f
C1141 VP.t4 VSUBS 1.10745f
C1142 VP.n67 VSUBS 0.644845f
C1143 VP.n68 VSUBS 2.93688f
C1144 VP.n69 VSUBS 0.081572f
C1145 VP.n70 VSUBS 0.050549f
C1146 VP.n71 VSUBS 0.093738f
C1147 VP.n72 VSUBS 0.093738f
C1148 VP.n73 VSUBS 0.068586f
C1149 VP.n74 VSUBS 0.050549f
C1150 VP.n75 VSUBS 0.050549f
C1151 VP.n76 VSUBS 0.050549f
C1152 VP.n77 VSUBS 0.093738f
C1153 VP.n78 VSUBS 0.093738f
C1154 VP.n79 VSUBS 0.053015f
C1155 VP.n80 VSUBS 0.050549f
C1156 VP.n81 VSUBS 0.050549f
C1157 VP.n82 VSUBS 0.088185f
C1158 VP.n83 VSUBS 0.093738f
C1159 VP.n84 VSUBS 0.092801f
C1160 VP.n85 VSUBS 0.050549f
C1161 VP.n86 VSUBS 0.050549f
C1162 VP.n87 VSUBS 0.050549f
C1163 VP.n88 VSUBS 0.10094f
C1164 VP.n89 VSUBS 0.093738f
C1165 VP.n90 VSUBS 0.0706f
C1166 VP.n91 VSUBS 0.050549f
C1167 VP.n92 VSUBS 0.050549f
C1168 VP.n93 VSUBS 0.0706f
C1169 VP.n94 VSUBS 0.093738f
C1170 VP.n95 VSUBS 0.10094f
C1171 VP.n96 VSUBS 0.050549f
C1172 VP.n97 VSUBS 0.050549f
C1173 VP.n98 VSUBS 0.050549f
C1174 VP.n99 VSUBS 0.092801f
C1175 VP.n100 VSUBS 0.093738f
C1176 VP.t3 VSUBS 1.10745f
C1177 VP.n101 VSUBS 0.468314f
C1178 VP.n102 VSUBS 0.088185f
C1179 VP.n103 VSUBS 0.050549f
C1180 VP.n104 VSUBS 0.050549f
C1181 VP.n105 VSUBS 0.050549f
C1182 VP.n106 VSUBS 0.093738f
C1183 VP.n107 VSUBS 0.093738f
C1184 VP.n108 VSUBS 0.078375f
C1185 VP.n109 VSUBS 0.050549f
C1186 VP.n110 VSUBS 0.050549f
C1187 VP.n111 VSUBS 0.050549f
C1188 VP.n112 VSUBS 0.093738f
C1189 VP.n113 VSUBS 0.093738f
C1190 VP.n114 VSUBS 0.059494f
C1191 VP.n115 VSUBS 0.081572f
C1192 VP.n116 VSUBS 0.138004f
.ends

