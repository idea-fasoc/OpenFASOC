* NGSPICE file created from diff_pair_sample_0626.ext - technology: sky130A

.subckt diff_pair_sample_0626 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t4 VN.t0 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0.20295 ps=1.56 w=1.23 l=1.56
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0 ps=0 w=1.23 l=1.56
X2 VDD2.t1 VN.t1 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.20295 pd=1.56 as=0.4797 ps=3.24 w=1.23 l=1.56
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0 ps=0 w=1.23 l=1.56
X4 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.20295 pd=1.56 as=0.4797 ps=3.24 w=1.23 l=1.56
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0 ps=0 w=1.23 l=1.56
X6 VTAIL.t5 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0.20295 ps=1.56 w=1.23 l=1.56
X7 VTAIL.t2 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0.20295 ps=1.56 w=1.23 l=1.56
X8 VDD2.t0 VN.t3 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.20295 pd=1.56 as=0.4797 ps=3.24 w=1.23 l=1.56
X9 VDD1.t1 VP.t2 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.20295 pd=1.56 as=0.4797 ps=3.24 w=1.23 l=1.56
X10 VTAIL.t7 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0.20295 ps=1.56 w=1.23 l=1.56
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4797 pd=3.24 as=0 ps=0 w=1.23 l=1.56
R0 VN.n0 VN.t0 56.228
R1 VN.n1 VN.t3 56.228
R2 VN.n0 VN.t1 55.9065
R3 VN.n1 VN.t2 55.9065
R4 VN VN.n1 48.1218
R5 VN VN.n0 12.8529
R6 VDD2.n2 VDD2.n0 175.123
R7 VDD2.n2 VDD2.n1 145.459
R8 VDD2.n1 VDD2.t3 16.0981
R9 VDD2.n1 VDD2.t0 16.0981
R10 VDD2.n0 VDD2.t2 16.0981
R11 VDD2.n0 VDD2.t1 16.0981
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n7 VTAIL.t3 154.939
R14 VTAIL.n0 VTAIL.t4 154.939
R15 VTAIL.n1 VTAIL.t0 154.939
R16 VTAIL.n2 VTAIL.t5 154.939
R17 VTAIL.n6 VTAIL.t6 154.939
R18 VTAIL.n5 VTAIL.t7 154.939
R19 VTAIL.n4 VTAIL.t1 154.939
R20 VTAIL.n3 VTAIL.t2 154.939
R21 VTAIL.n7 VTAIL.n6 15.0565
R22 VTAIL.n3 VTAIL.n2 15.0565
R23 VTAIL.n4 VTAIL.n3 1.62981
R24 VTAIL.n6 VTAIL.n5 1.62981
R25 VTAIL.n2 VTAIL.n1 1.62981
R26 VTAIL VTAIL.n0 0.873345
R27 VTAIL VTAIL.n7 0.756965
R28 VTAIL.n5 VTAIL.n4 0.470328
R29 VTAIL.n1 VTAIL.n0 0.470328
R30 B.n353 B.n352 585
R31 B.n354 B.n353 585
R32 B.n121 B.n62 585
R33 B.n120 B.n119 585
R34 B.n118 B.n117 585
R35 B.n116 B.n115 585
R36 B.n114 B.n113 585
R37 B.n112 B.n111 585
R38 B.n110 B.n109 585
R39 B.n108 B.n107 585
R40 B.n106 B.n105 585
R41 B.n103 B.n102 585
R42 B.n101 B.n100 585
R43 B.n99 B.n98 585
R44 B.n97 B.n96 585
R45 B.n95 B.n94 585
R46 B.n93 B.n92 585
R47 B.n91 B.n90 585
R48 B.n89 B.n88 585
R49 B.n87 B.n86 585
R50 B.n85 B.n84 585
R51 B.n83 B.n82 585
R52 B.n81 B.n80 585
R53 B.n79 B.n78 585
R54 B.n77 B.n76 585
R55 B.n75 B.n74 585
R56 B.n73 B.n72 585
R57 B.n71 B.n70 585
R58 B.n69 B.n68 585
R59 B.n46 B.n45 585
R60 B.n351 B.n47 585
R61 B.n355 B.n47 585
R62 B.n350 B.n349 585
R63 B.n349 B.n43 585
R64 B.n348 B.n42 585
R65 B.n361 B.n42 585
R66 B.n347 B.n41 585
R67 B.n362 B.n41 585
R68 B.n346 B.n40 585
R69 B.n363 B.n40 585
R70 B.n345 B.n344 585
R71 B.n344 B.n39 585
R72 B.n343 B.n35 585
R73 B.n369 B.n35 585
R74 B.n342 B.n34 585
R75 B.n370 B.n34 585
R76 B.n341 B.n33 585
R77 B.n371 B.n33 585
R78 B.n340 B.n339 585
R79 B.n339 B.n29 585
R80 B.n338 B.n28 585
R81 B.n377 B.n28 585
R82 B.n337 B.n27 585
R83 B.n378 B.n27 585
R84 B.n336 B.n26 585
R85 B.n379 B.n26 585
R86 B.n335 B.n334 585
R87 B.n334 B.n22 585
R88 B.n333 B.n21 585
R89 B.n385 B.n21 585
R90 B.n332 B.n20 585
R91 B.n386 B.n20 585
R92 B.n331 B.n19 585
R93 B.n387 B.n19 585
R94 B.n330 B.n329 585
R95 B.n329 B.n15 585
R96 B.n328 B.n14 585
R97 B.n393 B.n14 585
R98 B.n327 B.n13 585
R99 B.n394 B.n13 585
R100 B.n326 B.n12 585
R101 B.n395 B.n12 585
R102 B.n325 B.n324 585
R103 B.n324 B.n323 585
R104 B.n322 B.n321 585
R105 B.n322 B.n8 585
R106 B.n320 B.n7 585
R107 B.n402 B.n7 585
R108 B.n319 B.n6 585
R109 B.n403 B.n6 585
R110 B.n318 B.n5 585
R111 B.n404 B.n5 585
R112 B.n317 B.n316 585
R113 B.n316 B.n4 585
R114 B.n315 B.n122 585
R115 B.n315 B.n314 585
R116 B.n305 B.n123 585
R117 B.n124 B.n123 585
R118 B.n307 B.n306 585
R119 B.n308 B.n307 585
R120 B.n304 B.n129 585
R121 B.n129 B.n128 585
R122 B.n303 B.n302 585
R123 B.n302 B.n301 585
R124 B.n131 B.n130 585
R125 B.n132 B.n131 585
R126 B.n294 B.n293 585
R127 B.n295 B.n294 585
R128 B.n292 B.n137 585
R129 B.n137 B.n136 585
R130 B.n291 B.n290 585
R131 B.n290 B.n289 585
R132 B.n139 B.n138 585
R133 B.n140 B.n139 585
R134 B.n282 B.n281 585
R135 B.n283 B.n282 585
R136 B.n280 B.n145 585
R137 B.n145 B.n144 585
R138 B.n279 B.n278 585
R139 B.n278 B.n277 585
R140 B.n147 B.n146 585
R141 B.n148 B.n147 585
R142 B.n270 B.n269 585
R143 B.n271 B.n270 585
R144 B.n268 B.n153 585
R145 B.n153 B.n152 585
R146 B.n267 B.n266 585
R147 B.n266 B.n265 585
R148 B.n155 B.n154 585
R149 B.n258 B.n155 585
R150 B.n257 B.n256 585
R151 B.n259 B.n257 585
R152 B.n255 B.n160 585
R153 B.n160 B.n159 585
R154 B.n254 B.n253 585
R155 B.n253 B.n252 585
R156 B.n162 B.n161 585
R157 B.n163 B.n162 585
R158 B.n245 B.n244 585
R159 B.n246 B.n245 585
R160 B.n166 B.n165 585
R161 B.n187 B.n185 585
R162 B.n188 B.n184 585
R163 B.n188 B.n167 585
R164 B.n191 B.n190 585
R165 B.n192 B.n183 585
R166 B.n194 B.n193 585
R167 B.n196 B.n182 585
R168 B.n199 B.n198 585
R169 B.n200 B.n181 585
R170 B.n205 B.n204 585
R171 B.n207 B.n180 585
R172 B.n210 B.n209 585
R173 B.n211 B.n179 585
R174 B.n213 B.n212 585
R175 B.n215 B.n178 585
R176 B.n218 B.n217 585
R177 B.n219 B.n177 585
R178 B.n221 B.n220 585
R179 B.n223 B.n176 585
R180 B.n226 B.n225 585
R181 B.n227 B.n172 585
R182 B.n229 B.n228 585
R183 B.n231 B.n171 585
R184 B.n234 B.n233 585
R185 B.n235 B.n170 585
R186 B.n237 B.n236 585
R187 B.n239 B.n169 585
R188 B.n242 B.n241 585
R189 B.n243 B.n168 585
R190 B.n248 B.n247 585
R191 B.n247 B.n246 585
R192 B.n249 B.n164 585
R193 B.n164 B.n163 585
R194 B.n251 B.n250 585
R195 B.n252 B.n251 585
R196 B.n158 B.n157 585
R197 B.n159 B.n158 585
R198 B.n261 B.n260 585
R199 B.n260 B.n259 585
R200 B.n262 B.n156 585
R201 B.n258 B.n156 585
R202 B.n264 B.n263 585
R203 B.n265 B.n264 585
R204 B.n151 B.n150 585
R205 B.n152 B.n151 585
R206 B.n273 B.n272 585
R207 B.n272 B.n271 585
R208 B.n274 B.n149 585
R209 B.n149 B.n148 585
R210 B.n276 B.n275 585
R211 B.n277 B.n276 585
R212 B.n143 B.n142 585
R213 B.n144 B.n143 585
R214 B.n285 B.n284 585
R215 B.n284 B.n283 585
R216 B.n286 B.n141 585
R217 B.n141 B.n140 585
R218 B.n288 B.n287 585
R219 B.n289 B.n288 585
R220 B.n135 B.n134 585
R221 B.n136 B.n135 585
R222 B.n297 B.n296 585
R223 B.n296 B.n295 585
R224 B.n298 B.n133 585
R225 B.n133 B.n132 585
R226 B.n300 B.n299 585
R227 B.n301 B.n300 585
R228 B.n127 B.n126 585
R229 B.n128 B.n127 585
R230 B.n310 B.n309 585
R231 B.n309 B.n308 585
R232 B.n311 B.n125 585
R233 B.n125 B.n124 585
R234 B.n313 B.n312 585
R235 B.n314 B.n313 585
R236 B.n3 B.n0 585
R237 B.n4 B.n3 585
R238 B.n401 B.n1 585
R239 B.n402 B.n401 585
R240 B.n400 B.n399 585
R241 B.n400 B.n8 585
R242 B.n398 B.n9 585
R243 B.n323 B.n9 585
R244 B.n397 B.n396 585
R245 B.n396 B.n395 585
R246 B.n11 B.n10 585
R247 B.n394 B.n11 585
R248 B.n392 B.n391 585
R249 B.n393 B.n392 585
R250 B.n390 B.n16 585
R251 B.n16 B.n15 585
R252 B.n389 B.n388 585
R253 B.n388 B.n387 585
R254 B.n18 B.n17 585
R255 B.n386 B.n18 585
R256 B.n384 B.n383 585
R257 B.n385 B.n384 585
R258 B.n382 B.n23 585
R259 B.n23 B.n22 585
R260 B.n381 B.n380 585
R261 B.n380 B.n379 585
R262 B.n25 B.n24 585
R263 B.n378 B.n25 585
R264 B.n376 B.n375 585
R265 B.n377 B.n376 585
R266 B.n374 B.n30 585
R267 B.n30 B.n29 585
R268 B.n373 B.n372 585
R269 B.n372 B.n371 585
R270 B.n32 B.n31 585
R271 B.n370 B.n32 585
R272 B.n368 B.n367 585
R273 B.n369 B.n368 585
R274 B.n366 B.n36 585
R275 B.n39 B.n36 585
R276 B.n365 B.n364 585
R277 B.n364 B.n363 585
R278 B.n38 B.n37 585
R279 B.n362 B.n38 585
R280 B.n360 B.n359 585
R281 B.n361 B.n360 585
R282 B.n358 B.n44 585
R283 B.n44 B.n43 585
R284 B.n357 B.n356 585
R285 B.n356 B.n355 585
R286 B.n405 B.n404 585
R287 B.n403 B.n2 585
R288 B.n356 B.n46 583.793
R289 B.n353 B.n47 583.793
R290 B.n245 B.n168 583.793
R291 B.n247 B.n166 583.793
R292 B.n354 B.n61 256.663
R293 B.n354 B.n60 256.663
R294 B.n354 B.n59 256.663
R295 B.n354 B.n58 256.663
R296 B.n354 B.n57 256.663
R297 B.n354 B.n56 256.663
R298 B.n354 B.n55 256.663
R299 B.n354 B.n54 256.663
R300 B.n354 B.n53 256.663
R301 B.n354 B.n52 256.663
R302 B.n354 B.n51 256.663
R303 B.n354 B.n50 256.663
R304 B.n354 B.n49 256.663
R305 B.n354 B.n48 256.663
R306 B.n186 B.n167 256.663
R307 B.n189 B.n167 256.663
R308 B.n195 B.n167 256.663
R309 B.n197 B.n167 256.663
R310 B.n206 B.n167 256.663
R311 B.n208 B.n167 256.663
R312 B.n214 B.n167 256.663
R313 B.n216 B.n167 256.663
R314 B.n222 B.n167 256.663
R315 B.n224 B.n167 256.663
R316 B.n230 B.n167 256.663
R317 B.n232 B.n167 256.663
R318 B.n238 B.n167 256.663
R319 B.n240 B.n167 256.663
R320 B.n407 B.n406 256.663
R321 B.n246 B.n167 241.815
R322 B.n355 B.n354 241.815
R323 B.n65 B.t15 224.659
R324 B.n63 B.t8 224.659
R325 B.n173 B.t4 224.659
R326 B.n201 B.t12 224.659
R327 B.n65 B.t16 185.476
R328 B.n63 B.t10 185.476
R329 B.n173 B.t7 185.476
R330 B.n201 B.t14 185.476
R331 B.n70 B.n69 163.367
R332 B.n74 B.n73 163.367
R333 B.n78 B.n77 163.367
R334 B.n82 B.n81 163.367
R335 B.n86 B.n85 163.367
R336 B.n90 B.n89 163.367
R337 B.n94 B.n93 163.367
R338 B.n98 B.n97 163.367
R339 B.n102 B.n101 163.367
R340 B.n107 B.n106 163.367
R341 B.n111 B.n110 163.367
R342 B.n115 B.n114 163.367
R343 B.n119 B.n118 163.367
R344 B.n353 B.n62 163.367
R345 B.n245 B.n162 163.367
R346 B.n253 B.n162 163.367
R347 B.n253 B.n160 163.367
R348 B.n257 B.n160 163.367
R349 B.n257 B.n155 163.367
R350 B.n266 B.n155 163.367
R351 B.n266 B.n153 163.367
R352 B.n270 B.n153 163.367
R353 B.n270 B.n147 163.367
R354 B.n278 B.n147 163.367
R355 B.n278 B.n145 163.367
R356 B.n282 B.n145 163.367
R357 B.n282 B.n139 163.367
R358 B.n290 B.n139 163.367
R359 B.n290 B.n137 163.367
R360 B.n294 B.n137 163.367
R361 B.n294 B.n131 163.367
R362 B.n302 B.n131 163.367
R363 B.n302 B.n129 163.367
R364 B.n307 B.n129 163.367
R365 B.n307 B.n123 163.367
R366 B.n315 B.n123 163.367
R367 B.n316 B.n315 163.367
R368 B.n316 B.n5 163.367
R369 B.n6 B.n5 163.367
R370 B.n7 B.n6 163.367
R371 B.n322 B.n7 163.367
R372 B.n324 B.n322 163.367
R373 B.n324 B.n12 163.367
R374 B.n13 B.n12 163.367
R375 B.n14 B.n13 163.367
R376 B.n329 B.n14 163.367
R377 B.n329 B.n19 163.367
R378 B.n20 B.n19 163.367
R379 B.n21 B.n20 163.367
R380 B.n334 B.n21 163.367
R381 B.n334 B.n26 163.367
R382 B.n27 B.n26 163.367
R383 B.n28 B.n27 163.367
R384 B.n339 B.n28 163.367
R385 B.n339 B.n33 163.367
R386 B.n34 B.n33 163.367
R387 B.n35 B.n34 163.367
R388 B.n344 B.n35 163.367
R389 B.n344 B.n40 163.367
R390 B.n41 B.n40 163.367
R391 B.n42 B.n41 163.367
R392 B.n349 B.n42 163.367
R393 B.n349 B.n47 163.367
R394 B.n188 B.n187 163.367
R395 B.n190 B.n188 163.367
R396 B.n194 B.n183 163.367
R397 B.n198 B.n196 163.367
R398 B.n205 B.n181 163.367
R399 B.n209 B.n207 163.367
R400 B.n213 B.n179 163.367
R401 B.n217 B.n215 163.367
R402 B.n221 B.n177 163.367
R403 B.n225 B.n223 163.367
R404 B.n229 B.n172 163.367
R405 B.n233 B.n231 163.367
R406 B.n237 B.n170 163.367
R407 B.n241 B.n239 163.367
R408 B.n247 B.n164 163.367
R409 B.n251 B.n164 163.367
R410 B.n251 B.n158 163.367
R411 B.n260 B.n158 163.367
R412 B.n260 B.n156 163.367
R413 B.n264 B.n156 163.367
R414 B.n264 B.n151 163.367
R415 B.n272 B.n151 163.367
R416 B.n272 B.n149 163.367
R417 B.n276 B.n149 163.367
R418 B.n276 B.n143 163.367
R419 B.n284 B.n143 163.367
R420 B.n284 B.n141 163.367
R421 B.n288 B.n141 163.367
R422 B.n288 B.n135 163.367
R423 B.n296 B.n135 163.367
R424 B.n296 B.n133 163.367
R425 B.n300 B.n133 163.367
R426 B.n300 B.n127 163.367
R427 B.n309 B.n127 163.367
R428 B.n309 B.n125 163.367
R429 B.n313 B.n125 163.367
R430 B.n313 B.n3 163.367
R431 B.n405 B.n3 163.367
R432 B.n401 B.n2 163.367
R433 B.n401 B.n400 163.367
R434 B.n400 B.n9 163.367
R435 B.n396 B.n9 163.367
R436 B.n396 B.n11 163.367
R437 B.n392 B.n11 163.367
R438 B.n392 B.n16 163.367
R439 B.n388 B.n16 163.367
R440 B.n388 B.n18 163.367
R441 B.n384 B.n18 163.367
R442 B.n384 B.n23 163.367
R443 B.n380 B.n23 163.367
R444 B.n380 B.n25 163.367
R445 B.n376 B.n25 163.367
R446 B.n376 B.n30 163.367
R447 B.n372 B.n30 163.367
R448 B.n372 B.n32 163.367
R449 B.n368 B.n32 163.367
R450 B.n368 B.n36 163.367
R451 B.n364 B.n36 163.367
R452 B.n364 B.n38 163.367
R453 B.n360 B.n38 163.367
R454 B.n360 B.n44 163.367
R455 B.n356 B.n44 163.367
R456 B.n66 B.t17 148.821
R457 B.n64 B.t11 148.821
R458 B.n174 B.t6 148.821
R459 B.n202 B.t13 148.821
R460 B.n246 B.n163 114.989
R461 B.n252 B.n163 114.989
R462 B.n252 B.n159 114.989
R463 B.n259 B.n159 114.989
R464 B.n259 B.n258 114.989
R465 B.n265 B.n152 114.989
R466 B.n271 B.n152 114.989
R467 B.n271 B.n148 114.989
R468 B.n277 B.n148 114.989
R469 B.n277 B.n144 114.989
R470 B.n283 B.n144 114.989
R471 B.n283 B.n140 114.989
R472 B.n289 B.n140 114.989
R473 B.n295 B.n136 114.989
R474 B.n295 B.n132 114.989
R475 B.n301 B.n132 114.989
R476 B.n301 B.n128 114.989
R477 B.n308 B.n128 114.989
R478 B.n314 B.n124 114.989
R479 B.n314 B.n4 114.989
R480 B.n404 B.n4 114.989
R481 B.n404 B.n403 114.989
R482 B.n403 B.n402 114.989
R483 B.n402 B.n8 114.989
R484 B.n323 B.n8 114.989
R485 B.n395 B.n394 114.989
R486 B.n394 B.n393 114.989
R487 B.n393 B.n15 114.989
R488 B.n387 B.n15 114.989
R489 B.n387 B.n386 114.989
R490 B.n385 B.n22 114.989
R491 B.n379 B.n22 114.989
R492 B.n379 B.n378 114.989
R493 B.n378 B.n377 114.989
R494 B.n377 B.n29 114.989
R495 B.n371 B.n29 114.989
R496 B.n371 B.n370 114.989
R497 B.n370 B.n369 114.989
R498 B.n363 B.n39 114.989
R499 B.n363 B.n362 114.989
R500 B.n362 B.n361 114.989
R501 B.n361 B.n43 114.989
R502 B.n355 B.n43 114.989
R503 B.t0 B.n124 101.46
R504 B.n323 B.t3 101.46
R505 B.n258 B.t5 91.3149
R506 B.n39 B.t9 91.3149
R507 B.n48 B.n46 71.676
R508 B.n70 B.n49 71.676
R509 B.n74 B.n50 71.676
R510 B.n78 B.n51 71.676
R511 B.n82 B.n52 71.676
R512 B.n86 B.n53 71.676
R513 B.n90 B.n54 71.676
R514 B.n94 B.n55 71.676
R515 B.n98 B.n56 71.676
R516 B.n102 B.n57 71.676
R517 B.n107 B.n58 71.676
R518 B.n111 B.n59 71.676
R519 B.n115 B.n60 71.676
R520 B.n119 B.n61 71.676
R521 B.n62 B.n61 71.676
R522 B.n118 B.n60 71.676
R523 B.n114 B.n59 71.676
R524 B.n110 B.n58 71.676
R525 B.n106 B.n57 71.676
R526 B.n101 B.n56 71.676
R527 B.n97 B.n55 71.676
R528 B.n93 B.n54 71.676
R529 B.n89 B.n53 71.676
R530 B.n85 B.n52 71.676
R531 B.n81 B.n51 71.676
R532 B.n77 B.n50 71.676
R533 B.n73 B.n49 71.676
R534 B.n69 B.n48 71.676
R535 B.n186 B.n166 71.676
R536 B.n190 B.n189 71.676
R537 B.n195 B.n194 71.676
R538 B.n198 B.n197 71.676
R539 B.n206 B.n205 71.676
R540 B.n209 B.n208 71.676
R541 B.n214 B.n213 71.676
R542 B.n217 B.n216 71.676
R543 B.n222 B.n221 71.676
R544 B.n225 B.n224 71.676
R545 B.n230 B.n229 71.676
R546 B.n233 B.n232 71.676
R547 B.n238 B.n237 71.676
R548 B.n241 B.n240 71.676
R549 B.n187 B.n186 71.676
R550 B.n189 B.n183 71.676
R551 B.n196 B.n195 71.676
R552 B.n197 B.n181 71.676
R553 B.n207 B.n206 71.676
R554 B.n208 B.n179 71.676
R555 B.n215 B.n214 71.676
R556 B.n216 B.n177 71.676
R557 B.n223 B.n222 71.676
R558 B.n224 B.n172 71.676
R559 B.n231 B.n230 71.676
R560 B.n232 B.n170 71.676
R561 B.n239 B.n238 71.676
R562 B.n240 B.n168 71.676
R563 B.n406 B.n405 71.676
R564 B.n406 B.n2 71.676
R565 B.n289 B.t1 64.2588
R566 B.t2 B.n385 64.2588
R567 B.n67 B.n66 59.5399
R568 B.n104 B.n64 59.5399
R569 B.n175 B.n174 59.5399
R570 B.n203 B.n202 59.5399
R571 B.t1 B.n136 50.7307
R572 B.n386 B.t2 50.7307
R573 B.n248 B.n165 37.9322
R574 B.n244 B.n243 37.9322
R575 B.n352 B.n351 37.9322
R576 B.n357 B.n45 37.9322
R577 B.n66 B.n65 36.655
R578 B.n64 B.n63 36.655
R579 B.n174 B.n173 36.655
R580 B.n202 B.n201 36.655
R581 B.n265 B.t5 23.6746
R582 B.n369 B.t9 23.6746
R583 B B.n407 18.0485
R584 B.n308 B.t0 13.5286
R585 B.n395 B.t3 13.5286
R586 B.n249 B.n248 10.6151
R587 B.n250 B.n249 10.6151
R588 B.n250 B.n157 10.6151
R589 B.n261 B.n157 10.6151
R590 B.n262 B.n261 10.6151
R591 B.n263 B.n262 10.6151
R592 B.n263 B.n150 10.6151
R593 B.n273 B.n150 10.6151
R594 B.n274 B.n273 10.6151
R595 B.n275 B.n274 10.6151
R596 B.n275 B.n142 10.6151
R597 B.n285 B.n142 10.6151
R598 B.n286 B.n285 10.6151
R599 B.n287 B.n286 10.6151
R600 B.n287 B.n134 10.6151
R601 B.n297 B.n134 10.6151
R602 B.n298 B.n297 10.6151
R603 B.n299 B.n298 10.6151
R604 B.n299 B.n126 10.6151
R605 B.n310 B.n126 10.6151
R606 B.n311 B.n310 10.6151
R607 B.n312 B.n311 10.6151
R608 B.n312 B.n0 10.6151
R609 B.n185 B.n165 10.6151
R610 B.n185 B.n184 10.6151
R611 B.n191 B.n184 10.6151
R612 B.n192 B.n191 10.6151
R613 B.n193 B.n192 10.6151
R614 B.n193 B.n182 10.6151
R615 B.n199 B.n182 10.6151
R616 B.n200 B.n199 10.6151
R617 B.n204 B.n200 10.6151
R618 B.n210 B.n180 10.6151
R619 B.n211 B.n210 10.6151
R620 B.n212 B.n211 10.6151
R621 B.n212 B.n178 10.6151
R622 B.n218 B.n178 10.6151
R623 B.n219 B.n218 10.6151
R624 B.n220 B.n219 10.6151
R625 B.n220 B.n176 10.6151
R626 B.n227 B.n226 10.6151
R627 B.n228 B.n227 10.6151
R628 B.n228 B.n171 10.6151
R629 B.n234 B.n171 10.6151
R630 B.n235 B.n234 10.6151
R631 B.n236 B.n235 10.6151
R632 B.n236 B.n169 10.6151
R633 B.n242 B.n169 10.6151
R634 B.n243 B.n242 10.6151
R635 B.n244 B.n161 10.6151
R636 B.n254 B.n161 10.6151
R637 B.n255 B.n254 10.6151
R638 B.n256 B.n255 10.6151
R639 B.n256 B.n154 10.6151
R640 B.n267 B.n154 10.6151
R641 B.n268 B.n267 10.6151
R642 B.n269 B.n268 10.6151
R643 B.n269 B.n146 10.6151
R644 B.n279 B.n146 10.6151
R645 B.n280 B.n279 10.6151
R646 B.n281 B.n280 10.6151
R647 B.n281 B.n138 10.6151
R648 B.n291 B.n138 10.6151
R649 B.n292 B.n291 10.6151
R650 B.n293 B.n292 10.6151
R651 B.n293 B.n130 10.6151
R652 B.n303 B.n130 10.6151
R653 B.n304 B.n303 10.6151
R654 B.n306 B.n304 10.6151
R655 B.n306 B.n305 10.6151
R656 B.n305 B.n122 10.6151
R657 B.n317 B.n122 10.6151
R658 B.n318 B.n317 10.6151
R659 B.n319 B.n318 10.6151
R660 B.n320 B.n319 10.6151
R661 B.n321 B.n320 10.6151
R662 B.n325 B.n321 10.6151
R663 B.n326 B.n325 10.6151
R664 B.n327 B.n326 10.6151
R665 B.n328 B.n327 10.6151
R666 B.n330 B.n328 10.6151
R667 B.n331 B.n330 10.6151
R668 B.n332 B.n331 10.6151
R669 B.n333 B.n332 10.6151
R670 B.n335 B.n333 10.6151
R671 B.n336 B.n335 10.6151
R672 B.n337 B.n336 10.6151
R673 B.n338 B.n337 10.6151
R674 B.n340 B.n338 10.6151
R675 B.n341 B.n340 10.6151
R676 B.n342 B.n341 10.6151
R677 B.n343 B.n342 10.6151
R678 B.n345 B.n343 10.6151
R679 B.n346 B.n345 10.6151
R680 B.n347 B.n346 10.6151
R681 B.n348 B.n347 10.6151
R682 B.n350 B.n348 10.6151
R683 B.n351 B.n350 10.6151
R684 B.n399 B.n1 10.6151
R685 B.n399 B.n398 10.6151
R686 B.n398 B.n397 10.6151
R687 B.n397 B.n10 10.6151
R688 B.n391 B.n10 10.6151
R689 B.n391 B.n390 10.6151
R690 B.n390 B.n389 10.6151
R691 B.n389 B.n17 10.6151
R692 B.n383 B.n17 10.6151
R693 B.n383 B.n382 10.6151
R694 B.n382 B.n381 10.6151
R695 B.n381 B.n24 10.6151
R696 B.n375 B.n24 10.6151
R697 B.n375 B.n374 10.6151
R698 B.n374 B.n373 10.6151
R699 B.n373 B.n31 10.6151
R700 B.n367 B.n31 10.6151
R701 B.n367 B.n366 10.6151
R702 B.n366 B.n365 10.6151
R703 B.n365 B.n37 10.6151
R704 B.n359 B.n37 10.6151
R705 B.n359 B.n358 10.6151
R706 B.n358 B.n357 10.6151
R707 B.n68 B.n45 10.6151
R708 B.n71 B.n68 10.6151
R709 B.n72 B.n71 10.6151
R710 B.n75 B.n72 10.6151
R711 B.n76 B.n75 10.6151
R712 B.n79 B.n76 10.6151
R713 B.n80 B.n79 10.6151
R714 B.n83 B.n80 10.6151
R715 B.n84 B.n83 10.6151
R716 B.n88 B.n87 10.6151
R717 B.n91 B.n88 10.6151
R718 B.n92 B.n91 10.6151
R719 B.n95 B.n92 10.6151
R720 B.n96 B.n95 10.6151
R721 B.n99 B.n96 10.6151
R722 B.n100 B.n99 10.6151
R723 B.n103 B.n100 10.6151
R724 B.n108 B.n105 10.6151
R725 B.n109 B.n108 10.6151
R726 B.n112 B.n109 10.6151
R727 B.n113 B.n112 10.6151
R728 B.n116 B.n113 10.6151
R729 B.n117 B.n116 10.6151
R730 B.n120 B.n117 10.6151
R731 B.n121 B.n120 10.6151
R732 B.n352 B.n121 10.6151
R733 B.n407 B.n0 8.11757
R734 B.n407 B.n1 8.11757
R735 B.n203 B.n180 6.5566
R736 B.n176 B.n175 6.5566
R737 B.n87 B.n67 6.5566
R738 B.n104 B.n103 6.5566
R739 B.n204 B.n203 4.05904
R740 B.n226 B.n175 4.05904
R741 B.n84 B.n67 4.05904
R742 B.n105 B.n104 4.05904
R743 VP.n4 VP.n3 176.226
R744 VP.n12 VP.n11 176.226
R745 VP.n10 VP.n0 161.3
R746 VP.n9 VP.n8 161.3
R747 VP.n7 VP.n1 161.3
R748 VP.n6 VP.n5 161.3
R749 VP.n9 VP.n1 56.5193
R750 VP.n2 VP.t3 56.228
R751 VP.n2 VP.t2 55.9065
R752 VP.n3 VP.n2 47.7412
R753 VP.n5 VP.n1 24.4675
R754 VP.n10 VP.n9 24.4675
R755 VP.n4 VP.t1 19.0024
R756 VP.n11 VP.t0 19.0024
R757 VP.n5 VP.n4 9.54263
R758 VP.n11 VP.n10 9.54263
R759 VP.n6 VP.n3 0.189894
R760 VP.n7 VP.n6 0.189894
R761 VP.n8 VP.n7 0.189894
R762 VP.n8 VP.n0 0.189894
R763 VP.n12 VP.n0 0.189894
R764 VP VP.n12 0.0516364
R765 VDD1 VDD1.n1 175.648
R766 VDD1 VDD1.n0 145.518
R767 VDD1.n0 VDD1.t0 16.0981
R768 VDD1.n0 VDD1.t1 16.0981
R769 VDD1.n1 VDD1.t2 16.0981
R770 VDD1.n1 VDD1.t3 16.0981
C0 VDD1 VP 0.889541f
C1 VTAIL VN 1.10349f
C2 VDD2 VTAIL 2.36286f
C3 VN VP 3.45468f
C4 VDD1 VN 0.154852f
C5 VDD2 VP 0.336017f
C6 VDD2 VDD1 0.774955f
C7 VTAIL VP 1.1176f
C8 VDD2 VN 0.710064f
C9 VDD1 VTAIL 2.31562f
C10 VDD2 B 2.30635f
C11 VDD1 B 4.31129f
C12 VTAIL B 2.765514f
C13 VN B 7.261f
C14 VP B 5.770038f
C15 VDD1.t0 B 0.019626f
C16 VDD1.t1 B 0.019626f
C17 VDD1.n0 B 0.098167f
C18 VDD1.t2 B 0.019626f
C19 VDD1.t3 B 0.019626f
C20 VDD1.n1 B 0.219395f
C21 VP.n0 B 0.029688f
C22 VP.t0 B 0.11638f
C23 VP.n1 B 0.043339f
C24 VP.t3 B 0.251867f
C25 VP.t2 B 0.25076f
C26 VP.n2 B 0.951387f
C27 VP.n3 B 1.19882f
C28 VP.t1 B 0.11638f
C29 VP.n4 B 0.143924f
C30 VP.n5 B 0.038666f
C31 VP.n6 B 0.029688f
C32 VP.n7 B 0.029688f
C33 VP.n8 B 0.029688f
C34 VP.n9 B 0.043339f
C35 VP.n10 B 0.038666f
C36 VP.n11 B 0.143924f
C37 VP.n12 B 0.028873f
C38 VTAIL.t4 B 0.109294f
C39 VTAIL.n0 B 0.229227f
C40 VTAIL.t0 B 0.109294f
C41 VTAIL.n1 B 0.276618f
C42 VTAIL.t5 B 0.109294f
C43 VTAIL.n2 B 0.679794f
C44 VTAIL.t2 B 0.109294f
C45 VTAIL.n3 B 0.679794f
C46 VTAIL.t1 B 0.109294f
C47 VTAIL.n4 B 0.276618f
C48 VTAIL.t7 B 0.109294f
C49 VTAIL.n5 B 0.276618f
C50 VTAIL.t6 B 0.109294f
C51 VTAIL.n6 B 0.679794f
C52 VTAIL.t3 B 0.109294f
C53 VTAIL.n7 B 0.625111f
C54 VDD2.t2 B 0.021166f
C55 VDD2.t1 B 0.021166f
C56 VDD2.n0 B 0.227148f
C57 VDD2.t3 B 0.021166f
C58 VDD2.t0 B 0.021166f
C59 VDD2.n1 B 0.105757f
C60 VDD2.n2 B 1.86342f
C61 VN.t0 B 0.248899f
C62 VN.t1 B 0.247805f
C63 VN.n0 B 0.183772f
C64 VN.t3 B 0.248899f
C65 VN.t2 B 0.247805f
C66 VN.n1 B 0.956686f
.ends

