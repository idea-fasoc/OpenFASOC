* NGSPICE file created from diff_pair_sample_1641.ext - technology: sky130A

.subckt diff_pair_sample_1641 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=1.95855 ps=12.2 w=11.87 l=2.95
X1 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=4.6293 ps=24.52 w=11.87 l=2.95
X2 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=1.95855 ps=12.2 w=11.87 l=2.95
X3 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=0 ps=0 w=11.87 l=2.95
X4 VDD1.t4 VP.t1 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=4.6293 ps=24.52 w=11.87 l=2.95
X5 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=0 ps=0 w=11.87 l=2.95
X6 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=4.6293 ps=24.52 w=11.87 l=2.95
X7 VTAIL.t4 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=1.95855 ps=12.2 w=11.87 l=2.95
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=0 ps=0 w=11.87 l=2.95
X9 VDD1.t3 VP.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=4.6293 ps=24.52 w=11.87 l=2.95
X10 VTAIL.t0 VN.t4 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=1.95855 ps=12.2 w=11.87 l=2.95
X11 VTAIL.t6 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=1.95855 ps=12.2 w=11.87 l=2.95
X12 VTAIL.t11 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.95855 pd=12.2 as=1.95855 ps=12.2 w=11.87 l=2.95
X13 VDD2.t0 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=1.95855 ps=12.2 w=11.87 l=2.95
X14 VDD1.t0 VP.t5 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=1.95855 ps=12.2 w=11.87 l=2.95
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.6293 pd=24.52 as=0 ps=0 w=11.87 l=2.95
R0 VP.n14 VP.n11 161.3
R1 VP.n16 VP.n15 161.3
R2 VP.n17 VP.n10 161.3
R3 VP.n19 VP.n18 161.3
R4 VP.n20 VP.n9 161.3
R5 VP.n22 VP.n21 161.3
R6 VP.n23 VP.n8 161.3
R7 VP.n48 VP.n0 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n45 VP.n1 161.3
R10 VP.n44 VP.n43 161.3
R11 VP.n42 VP.n2 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n39 VP.n3 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n35 VP.n4 161.3
R16 VP.n34 VP.n33 161.3
R17 VP.n32 VP.n5 161.3
R18 VP.n31 VP.n30 161.3
R19 VP.n29 VP.n6 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n13 VP.t5 129.436
R22 VP.n26 VP.n7 109.288
R23 VP.n50 VP.n49 109.288
R24 VP.n25 VP.n24 109.288
R25 VP.n7 VP.t0 96.9724
R26 VP.n36 VP.t4 96.9724
R27 VP.n49 VP.t1 96.9724
R28 VP.n24 VP.t2 96.9724
R29 VP.n12 VP.t3 96.9724
R30 VP.n13 VP.n12 61.6325
R31 VP.n34 VP.n5 51.1773
R32 VP.n43 VP.n42 51.1773
R33 VP.n18 VP.n17 51.1773
R34 VP.n26 VP.n25 49.9238
R35 VP.n30 VP.n5 29.8095
R36 VP.n43 VP.n1 29.8095
R37 VP.n18 VP.n9 29.8095
R38 VP.n29 VP.n28 24.4675
R39 VP.n30 VP.n29 24.4675
R40 VP.n35 VP.n34 24.4675
R41 VP.n37 VP.n35 24.4675
R42 VP.n41 VP.n3 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n1 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n22 VP.n9 24.4675
R47 VP.n23 VP.n22 24.4675
R48 VP.n16 VP.n11 24.4675
R49 VP.n17 VP.n16 24.4675
R50 VP.n37 VP.n36 12.234
R51 VP.n36 VP.n3 12.234
R52 VP.n12 VP.n11 12.234
R53 VP.n14 VP.n13 5.14959
R54 VP.n28 VP.n7 1.46852
R55 VP.n49 VP.n48 1.46852
R56 VP.n24 VP.n23 1.46852
R57 VP.n25 VP.n8 0.278367
R58 VP.n27 VP.n26 0.278367
R59 VP.n50 VP.n0 0.278367
R60 VP.n15 VP.n14 0.189894
R61 VP.n15 VP.n10 0.189894
R62 VP.n19 VP.n10 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n8 0.189894
R66 VP.n27 VP.n6 0.189894
R67 VP.n31 VP.n6 0.189894
R68 VP.n32 VP.n31 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n33 VP.n4 0.189894
R71 VP.n38 VP.n4 0.189894
R72 VP.n39 VP.n38 0.189894
R73 VP.n40 VP.n39 0.189894
R74 VP.n40 VP.n2 0.189894
R75 VP.n44 VP.n2 0.189894
R76 VP.n45 VP.n44 0.189894
R77 VP.n46 VP.n45 0.189894
R78 VP.n46 VP.n0 0.189894
R79 VP VP.n50 0.153454
R80 VTAIL.n7 VTAIL.t2 49.1026
R81 VTAIL.n11 VTAIL.t3 49.1024
R82 VTAIL.n2 VTAIL.t8 49.1024
R83 VTAIL.n10 VTAIL.t9 49.1024
R84 VTAIL.n9 VTAIL.n8 47.4346
R85 VTAIL.n6 VTAIL.n5 47.4346
R86 VTAIL.n1 VTAIL.n0 47.4343
R87 VTAIL.n4 VTAIL.n3 47.4343
R88 VTAIL.n6 VTAIL.n4 28.2548
R89 VTAIL.n11 VTAIL.n10 25.4272
R90 VTAIL.n7 VTAIL.n6 2.82809
R91 VTAIL.n10 VTAIL.n9 2.82809
R92 VTAIL.n4 VTAIL.n2 2.82809
R93 VTAIL VTAIL.n11 2.063
R94 VTAIL.n9 VTAIL.n7 1.88412
R95 VTAIL.n2 VTAIL.n1 1.88412
R96 VTAIL.n0 VTAIL.t1 1.66857
R97 VTAIL.n0 VTAIL.t0 1.66857
R98 VTAIL.n3 VTAIL.t10 1.66857
R99 VTAIL.n3 VTAIL.t11 1.66857
R100 VTAIL.n8 VTAIL.t7 1.66857
R101 VTAIL.n8 VTAIL.t6 1.66857
R102 VTAIL.n5 VTAIL.t5 1.66857
R103 VTAIL.n5 VTAIL.t4 1.66857
R104 VTAIL VTAIL.n1 0.765586
R105 VDD1 VDD1.t0 67.9603
R106 VDD1.n1 VDD1.t5 67.8465
R107 VDD1.n1 VDD1.n0 64.7647
R108 VDD1.n3 VDD1.n2 64.1132
R109 VDD1.n3 VDD1.n1 45.1345
R110 VDD1.n2 VDD1.t2 1.66857
R111 VDD1.n2 VDD1.t3 1.66857
R112 VDD1.n0 VDD1.t1 1.66857
R113 VDD1.n0 VDD1.t4 1.66857
R114 VDD1 VDD1.n3 0.649207
R115 B.n662 B.n661 585
R116 B.n664 B.n137 585
R117 B.n667 B.n666 585
R118 B.n668 B.n136 585
R119 B.n670 B.n669 585
R120 B.n672 B.n135 585
R121 B.n675 B.n674 585
R122 B.n676 B.n134 585
R123 B.n678 B.n677 585
R124 B.n680 B.n133 585
R125 B.n683 B.n682 585
R126 B.n684 B.n132 585
R127 B.n686 B.n685 585
R128 B.n688 B.n131 585
R129 B.n691 B.n690 585
R130 B.n692 B.n130 585
R131 B.n694 B.n693 585
R132 B.n696 B.n129 585
R133 B.n699 B.n698 585
R134 B.n700 B.n128 585
R135 B.n702 B.n701 585
R136 B.n704 B.n127 585
R137 B.n707 B.n706 585
R138 B.n708 B.n126 585
R139 B.n710 B.n709 585
R140 B.n712 B.n125 585
R141 B.n715 B.n714 585
R142 B.n716 B.n124 585
R143 B.n718 B.n717 585
R144 B.n720 B.n123 585
R145 B.n723 B.n722 585
R146 B.n724 B.n122 585
R147 B.n726 B.n725 585
R148 B.n728 B.n121 585
R149 B.n731 B.n730 585
R150 B.n732 B.n120 585
R151 B.n734 B.n733 585
R152 B.n736 B.n119 585
R153 B.n739 B.n738 585
R154 B.n740 B.n115 585
R155 B.n742 B.n741 585
R156 B.n744 B.n114 585
R157 B.n747 B.n746 585
R158 B.n748 B.n113 585
R159 B.n750 B.n749 585
R160 B.n752 B.n112 585
R161 B.n755 B.n754 585
R162 B.n756 B.n111 585
R163 B.n758 B.n757 585
R164 B.n760 B.n110 585
R165 B.n763 B.n762 585
R166 B.n765 B.n107 585
R167 B.n767 B.n766 585
R168 B.n769 B.n106 585
R169 B.n772 B.n771 585
R170 B.n773 B.n105 585
R171 B.n775 B.n774 585
R172 B.n777 B.n104 585
R173 B.n780 B.n779 585
R174 B.n781 B.n103 585
R175 B.n783 B.n782 585
R176 B.n785 B.n102 585
R177 B.n788 B.n787 585
R178 B.n789 B.n101 585
R179 B.n791 B.n790 585
R180 B.n793 B.n100 585
R181 B.n796 B.n795 585
R182 B.n797 B.n99 585
R183 B.n799 B.n798 585
R184 B.n801 B.n98 585
R185 B.n804 B.n803 585
R186 B.n805 B.n97 585
R187 B.n807 B.n806 585
R188 B.n809 B.n96 585
R189 B.n812 B.n811 585
R190 B.n813 B.n95 585
R191 B.n815 B.n814 585
R192 B.n817 B.n94 585
R193 B.n820 B.n819 585
R194 B.n821 B.n93 585
R195 B.n823 B.n822 585
R196 B.n825 B.n92 585
R197 B.n828 B.n827 585
R198 B.n829 B.n91 585
R199 B.n831 B.n830 585
R200 B.n833 B.n90 585
R201 B.n836 B.n835 585
R202 B.n837 B.n89 585
R203 B.n839 B.n838 585
R204 B.n841 B.n88 585
R205 B.n844 B.n843 585
R206 B.n845 B.n87 585
R207 B.n660 B.n85 585
R208 B.n848 B.n85 585
R209 B.n659 B.n84 585
R210 B.n849 B.n84 585
R211 B.n658 B.n83 585
R212 B.n850 B.n83 585
R213 B.n657 B.n656 585
R214 B.n656 B.n79 585
R215 B.n655 B.n78 585
R216 B.n856 B.n78 585
R217 B.n654 B.n77 585
R218 B.n857 B.n77 585
R219 B.n653 B.n76 585
R220 B.n858 B.n76 585
R221 B.n652 B.n651 585
R222 B.n651 B.n75 585
R223 B.n650 B.n71 585
R224 B.n864 B.n71 585
R225 B.n649 B.n70 585
R226 B.n865 B.n70 585
R227 B.n648 B.n69 585
R228 B.n866 B.n69 585
R229 B.n647 B.n646 585
R230 B.n646 B.n65 585
R231 B.n645 B.n64 585
R232 B.n872 B.n64 585
R233 B.n644 B.n63 585
R234 B.n873 B.n63 585
R235 B.n643 B.n62 585
R236 B.n874 B.n62 585
R237 B.n642 B.n641 585
R238 B.n641 B.n58 585
R239 B.n640 B.n57 585
R240 B.n880 B.n57 585
R241 B.n639 B.n56 585
R242 B.n881 B.n56 585
R243 B.n638 B.n55 585
R244 B.n882 B.n55 585
R245 B.n637 B.n636 585
R246 B.n636 B.n51 585
R247 B.n635 B.n50 585
R248 B.n888 B.n50 585
R249 B.n634 B.n49 585
R250 B.n889 B.n49 585
R251 B.n633 B.n48 585
R252 B.n890 B.n48 585
R253 B.n632 B.n631 585
R254 B.n631 B.n44 585
R255 B.n630 B.n43 585
R256 B.n896 B.n43 585
R257 B.n629 B.n42 585
R258 B.n897 B.n42 585
R259 B.n628 B.n41 585
R260 B.n898 B.n41 585
R261 B.n627 B.n626 585
R262 B.n626 B.n37 585
R263 B.n625 B.n36 585
R264 B.n904 B.n36 585
R265 B.n624 B.n35 585
R266 B.n905 B.n35 585
R267 B.n623 B.n34 585
R268 B.n906 B.n34 585
R269 B.n622 B.n621 585
R270 B.n621 B.n30 585
R271 B.n620 B.n29 585
R272 B.n912 B.n29 585
R273 B.n619 B.n28 585
R274 B.n913 B.n28 585
R275 B.n618 B.n27 585
R276 B.n914 B.n27 585
R277 B.n617 B.n616 585
R278 B.n616 B.n23 585
R279 B.n615 B.n22 585
R280 B.n920 B.n22 585
R281 B.n614 B.n21 585
R282 B.n921 B.n21 585
R283 B.n613 B.n20 585
R284 B.n922 B.n20 585
R285 B.n612 B.n611 585
R286 B.n611 B.n16 585
R287 B.n610 B.n15 585
R288 B.n928 B.n15 585
R289 B.n609 B.n14 585
R290 B.n929 B.n14 585
R291 B.n608 B.n13 585
R292 B.n930 B.n13 585
R293 B.n607 B.n606 585
R294 B.n606 B.n12 585
R295 B.n605 B.n604 585
R296 B.n605 B.n8 585
R297 B.n603 B.n7 585
R298 B.n937 B.n7 585
R299 B.n602 B.n6 585
R300 B.n938 B.n6 585
R301 B.n601 B.n5 585
R302 B.n939 B.n5 585
R303 B.n600 B.n599 585
R304 B.n599 B.n4 585
R305 B.n598 B.n138 585
R306 B.n598 B.n597 585
R307 B.n588 B.n139 585
R308 B.n140 B.n139 585
R309 B.n590 B.n589 585
R310 B.n591 B.n590 585
R311 B.n587 B.n145 585
R312 B.n145 B.n144 585
R313 B.n586 B.n585 585
R314 B.n585 B.n584 585
R315 B.n147 B.n146 585
R316 B.n148 B.n147 585
R317 B.n577 B.n576 585
R318 B.n578 B.n577 585
R319 B.n575 B.n153 585
R320 B.n153 B.n152 585
R321 B.n574 B.n573 585
R322 B.n573 B.n572 585
R323 B.n155 B.n154 585
R324 B.n156 B.n155 585
R325 B.n565 B.n564 585
R326 B.n566 B.n565 585
R327 B.n563 B.n161 585
R328 B.n161 B.n160 585
R329 B.n562 B.n561 585
R330 B.n561 B.n560 585
R331 B.n163 B.n162 585
R332 B.n164 B.n163 585
R333 B.n553 B.n552 585
R334 B.n554 B.n553 585
R335 B.n551 B.n169 585
R336 B.n169 B.n168 585
R337 B.n550 B.n549 585
R338 B.n549 B.n548 585
R339 B.n171 B.n170 585
R340 B.n172 B.n171 585
R341 B.n541 B.n540 585
R342 B.n542 B.n541 585
R343 B.n539 B.n177 585
R344 B.n177 B.n176 585
R345 B.n538 B.n537 585
R346 B.n537 B.n536 585
R347 B.n179 B.n178 585
R348 B.n180 B.n179 585
R349 B.n529 B.n528 585
R350 B.n530 B.n529 585
R351 B.n527 B.n185 585
R352 B.n185 B.n184 585
R353 B.n526 B.n525 585
R354 B.n525 B.n524 585
R355 B.n187 B.n186 585
R356 B.n188 B.n187 585
R357 B.n517 B.n516 585
R358 B.n518 B.n517 585
R359 B.n515 B.n193 585
R360 B.n193 B.n192 585
R361 B.n514 B.n513 585
R362 B.n513 B.n512 585
R363 B.n195 B.n194 585
R364 B.n196 B.n195 585
R365 B.n505 B.n504 585
R366 B.n506 B.n505 585
R367 B.n503 B.n201 585
R368 B.n201 B.n200 585
R369 B.n502 B.n501 585
R370 B.n501 B.n500 585
R371 B.n203 B.n202 585
R372 B.n204 B.n203 585
R373 B.n493 B.n492 585
R374 B.n494 B.n493 585
R375 B.n491 B.n209 585
R376 B.n209 B.n208 585
R377 B.n490 B.n489 585
R378 B.n489 B.n488 585
R379 B.n211 B.n210 585
R380 B.n481 B.n211 585
R381 B.n480 B.n479 585
R382 B.n482 B.n480 585
R383 B.n478 B.n216 585
R384 B.n216 B.n215 585
R385 B.n477 B.n476 585
R386 B.n476 B.n475 585
R387 B.n218 B.n217 585
R388 B.n219 B.n218 585
R389 B.n468 B.n467 585
R390 B.n469 B.n468 585
R391 B.n466 B.n224 585
R392 B.n224 B.n223 585
R393 B.n465 B.n464 585
R394 B.n464 B.n463 585
R395 B.n460 B.n228 585
R396 B.n459 B.n458 585
R397 B.n456 B.n229 585
R398 B.n456 B.n227 585
R399 B.n455 B.n454 585
R400 B.n453 B.n452 585
R401 B.n451 B.n231 585
R402 B.n449 B.n448 585
R403 B.n447 B.n232 585
R404 B.n446 B.n445 585
R405 B.n443 B.n233 585
R406 B.n441 B.n440 585
R407 B.n439 B.n234 585
R408 B.n438 B.n437 585
R409 B.n435 B.n235 585
R410 B.n433 B.n432 585
R411 B.n431 B.n236 585
R412 B.n430 B.n429 585
R413 B.n427 B.n237 585
R414 B.n425 B.n424 585
R415 B.n423 B.n238 585
R416 B.n422 B.n421 585
R417 B.n419 B.n239 585
R418 B.n417 B.n416 585
R419 B.n415 B.n240 585
R420 B.n414 B.n413 585
R421 B.n411 B.n241 585
R422 B.n409 B.n408 585
R423 B.n407 B.n242 585
R424 B.n406 B.n405 585
R425 B.n403 B.n243 585
R426 B.n401 B.n400 585
R427 B.n399 B.n244 585
R428 B.n398 B.n397 585
R429 B.n395 B.n245 585
R430 B.n393 B.n392 585
R431 B.n391 B.n246 585
R432 B.n390 B.n389 585
R433 B.n387 B.n247 585
R434 B.n385 B.n384 585
R435 B.n383 B.n248 585
R436 B.n382 B.n381 585
R437 B.n379 B.n378 585
R438 B.n377 B.n376 585
R439 B.n375 B.n253 585
R440 B.n373 B.n372 585
R441 B.n371 B.n254 585
R442 B.n370 B.n369 585
R443 B.n367 B.n255 585
R444 B.n365 B.n364 585
R445 B.n363 B.n256 585
R446 B.n362 B.n361 585
R447 B.n359 B.n358 585
R448 B.n357 B.n356 585
R449 B.n355 B.n261 585
R450 B.n353 B.n352 585
R451 B.n351 B.n262 585
R452 B.n350 B.n349 585
R453 B.n347 B.n263 585
R454 B.n345 B.n344 585
R455 B.n343 B.n264 585
R456 B.n342 B.n341 585
R457 B.n339 B.n265 585
R458 B.n337 B.n336 585
R459 B.n335 B.n266 585
R460 B.n334 B.n333 585
R461 B.n331 B.n267 585
R462 B.n329 B.n328 585
R463 B.n327 B.n268 585
R464 B.n326 B.n325 585
R465 B.n323 B.n269 585
R466 B.n321 B.n320 585
R467 B.n319 B.n270 585
R468 B.n318 B.n317 585
R469 B.n315 B.n271 585
R470 B.n313 B.n312 585
R471 B.n311 B.n272 585
R472 B.n310 B.n309 585
R473 B.n307 B.n273 585
R474 B.n305 B.n304 585
R475 B.n303 B.n274 585
R476 B.n302 B.n301 585
R477 B.n299 B.n275 585
R478 B.n297 B.n296 585
R479 B.n295 B.n276 585
R480 B.n294 B.n293 585
R481 B.n291 B.n277 585
R482 B.n289 B.n288 585
R483 B.n287 B.n278 585
R484 B.n286 B.n285 585
R485 B.n283 B.n279 585
R486 B.n281 B.n280 585
R487 B.n226 B.n225 585
R488 B.n227 B.n226 585
R489 B.n462 B.n461 585
R490 B.n463 B.n462 585
R491 B.n222 B.n221 585
R492 B.n223 B.n222 585
R493 B.n471 B.n470 585
R494 B.n470 B.n469 585
R495 B.n472 B.n220 585
R496 B.n220 B.n219 585
R497 B.n474 B.n473 585
R498 B.n475 B.n474 585
R499 B.n214 B.n213 585
R500 B.n215 B.n214 585
R501 B.n484 B.n483 585
R502 B.n483 B.n482 585
R503 B.n485 B.n212 585
R504 B.n481 B.n212 585
R505 B.n487 B.n486 585
R506 B.n488 B.n487 585
R507 B.n207 B.n206 585
R508 B.n208 B.n207 585
R509 B.n496 B.n495 585
R510 B.n495 B.n494 585
R511 B.n497 B.n205 585
R512 B.n205 B.n204 585
R513 B.n499 B.n498 585
R514 B.n500 B.n499 585
R515 B.n199 B.n198 585
R516 B.n200 B.n199 585
R517 B.n508 B.n507 585
R518 B.n507 B.n506 585
R519 B.n509 B.n197 585
R520 B.n197 B.n196 585
R521 B.n511 B.n510 585
R522 B.n512 B.n511 585
R523 B.n191 B.n190 585
R524 B.n192 B.n191 585
R525 B.n520 B.n519 585
R526 B.n519 B.n518 585
R527 B.n521 B.n189 585
R528 B.n189 B.n188 585
R529 B.n523 B.n522 585
R530 B.n524 B.n523 585
R531 B.n183 B.n182 585
R532 B.n184 B.n183 585
R533 B.n532 B.n531 585
R534 B.n531 B.n530 585
R535 B.n533 B.n181 585
R536 B.n181 B.n180 585
R537 B.n535 B.n534 585
R538 B.n536 B.n535 585
R539 B.n175 B.n174 585
R540 B.n176 B.n175 585
R541 B.n544 B.n543 585
R542 B.n543 B.n542 585
R543 B.n545 B.n173 585
R544 B.n173 B.n172 585
R545 B.n547 B.n546 585
R546 B.n548 B.n547 585
R547 B.n167 B.n166 585
R548 B.n168 B.n167 585
R549 B.n556 B.n555 585
R550 B.n555 B.n554 585
R551 B.n557 B.n165 585
R552 B.n165 B.n164 585
R553 B.n559 B.n558 585
R554 B.n560 B.n559 585
R555 B.n159 B.n158 585
R556 B.n160 B.n159 585
R557 B.n568 B.n567 585
R558 B.n567 B.n566 585
R559 B.n569 B.n157 585
R560 B.n157 B.n156 585
R561 B.n571 B.n570 585
R562 B.n572 B.n571 585
R563 B.n151 B.n150 585
R564 B.n152 B.n151 585
R565 B.n580 B.n579 585
R566 B.n579 B.n578 585
R567 B.n581 B.n149 585
R568 B.n149 B.n148 585
R569 B.n583 B.n582 585
R570 B.n584 B.n583 585
R571 B.n143 B.n142 585
R572 B.n144 B.n143 585
R573 B.n593 B.n592 585
R574 B.n592 B.n591 585
R575 B.n594 B.n141 585
R576 B.n141 B.n140 585
R577 B.n596 B.n595 585
R578 B.n597 B.n596 585
R579 B.n3 B.n0 585
R580 B.n4 B.n3 585
R581 B.n936 B.n1 585
R582 B.n937 B.n936 585
R583 B.n935 B.n934 585
R584 B.n935 B.n8 585
R585 B.n933 B.n9 585
R586 B.n12 B.n9 585
R587 B.n932 B.n931 585
R588 B.n931 B.n930 585
R589 B.n11 B.n10 585
R590 B.n929 B.n11 585
R591 B.n927 B.n926 585
R592 B.n928 B.n927 585
R593 B.n925 B.n17 585
R594 B.n17 B.n16 585
R595 B.n924 B.n923 585
R596 B.n923 B.n922 585
R597 B.n19 B.n18 585
R598 B.n921 B.n19 585
R599 B.n919 B.n918 585
R600 B.n920 B.n919 585
R601 B.n917 B.n24 585
R602 B.n24 B.n23 585
R603 B.n916 B.n915 585
R604 B.n915 B.n914 585
R605 B.n26 B.n25 585
R606 B.n913 B.n26 585
R607 B.n911 B.n910 585
R608 B.n912 B.n911 585
R609 B.n909 B.n31 585
R610 B.n31 B.n30 585
R611 B.n908 B.n907 585
R612 B.n907 B.n906 585
R613 B.n33 B.n32 585
R614 B.n905 B.n33 585
R615 B.n903 B.n902 585
R616 B.n904 B.n903 585
R617 B.n901 B.n38 585
R618 B.n38 B.n37 585
R619 B.n900 B.n899 585
R620 B.n899 B.n898 585
R621 B.n40 B.n39 585
R622 B.n897 B.n40 585
R623 B.n895 B.n894 585
R624 B.n896 B.n895 585
R625 B.n893 B.n45 585
R626 B.n45 B.n44 585
R627 B.n892 B.n891 585
R628 B.n891 B.n890 585
R629 B.n47 B.n46 585
R630 B.n889 B.n47 585
R631 B.n887 B.n886 585
R632 B.n888 B.n887 585
R633 B.n885 B.n52 585
R634 B.n52 B.n51 585
R635 B.n884 B.n883 585
R636 B.n883 B.n882 585
R637 B.n54 B.n53 585
R638 B.n881 B.n54 585
R639 B.n879 B.n878 585
R640 B.n880 B.n879 585
R641 B.n877 B.n59 585
R642 B.n59 B.n58 585
R643 B.n876 B.n875 585
R644 B.n875 B.n874 585
R645 B.n61 B.n60 585
R646 B.n873 B.n61 585
R647 B.n871 B.n870 585
R648 B.n872 B.n871 585
R649 B.n869 B.n66 585
R650 B.n66 B.n65 585
R651 B.n868 B.n867 585
R652 B.n867 B.n866 585
R653 B.n68 B.n67 585
R654 B.n865 B.n68 585
R655 B.n863 B.n862 585
R656 B.n864 B.n863 585
R657 B.n861 B.n72 585
R658 B.n75 B.n72 585
R659 B.n860 B.n859 585
R660 B.n859 B.n858 585
R661 B.n74 B.n73 585
R662 B.n857 B.n74 585
R663 B.n855 B.n854 585
R664 B.n856 B.n855 585
R665 B.n853 B.n80 585
R666 B.n80 B.n79 585
R667 B.n852 B.n851 585
R668 B.n851 B.n850 585
R669 B.n82 B.n81 585
R670 B.n849 B.n82 585
R671 B.n847 B.n846 585
R672 B.n848 B.n847 585
R673 B.n940 B.n939 585
R674 B.n938 B.n2 585
R675 B.n847 B.n87 535.745
R676 B.n662 B.n85 535.745
R677 B.n464 B.n226 535.745
R678 B.n462 B.n228 535.745
R679 B.n108 B.t14 305.493
R680 B.n116 B.t6 305.493
R681 B.n257 B.t10 305.493
R682 B.n249 B.t17 305.493
R683 B.n663 B.n86 256.663
R684 B.n665 B.n86 256.663
R685 B.n671 B.n86 256.663
R686 B.n673 B.n86 256.663
R687 B.n679 B.n86 256.663
R688 B.n681 B.n86 256.663
R689 B.n687 B.n86 256.663
R690 B.n689 B.n86 256.663
R691 B.n695 B.n86 256.663
R692 B.n697 B.n86 256.663
R693 B.n703 B.n86 256.663
R694 B.n705 B.n86 256.663
R695 B.n711 B.n86 256.663
R696 B.n713 B.n86 256.663
R697 B.n719 B.n86 256.663
R698 B.n721 B.n86 256.663
R699 B.n727 B.n86 256.663
R700 B.n729 B.n86 256.663
R701 B.n735 B.n86 256.663
R702 B.n737 B.n86 256.663
R703 B.n743 B.n86 256.663
R704 B.n745 B.n86 256.663
R705 B.n751 B.n86 256.663
R706 B.n753 B.n86 256.663
R707 B.n759 B.n86 256.663
R708 B.n761 B.n86 256.663
R709 B.n768 B.n86 256.663
R710 B.n770 B.n86 256.663
R711 B.n776 B.n86 256.663
R712 B.n778 B.n86 256.663
R713 B.n784 B.n86 256.663
R714 B.n786 B.n86 256.663
R715 B.n792 B.n86 256.663
R716 B.n794 B.n86 256.663
R717 B.n800 B.n86 256.663
R718 B.n802 B.n86 256.663
R719 B.n808 B.n86 256.663
R720 B.n810 B.n86 256.663
R721 B.n816 B.n86 256.663
R722 B.n818 B.n86 256.663
R723 B.n824 B.n86 256.663
R724 B.n826 B.n86 256.663
R725 B.n832 B.n86 256.663
R726 B.n834 B.n86 256.663
R727 B.n840 B.n86 256.663
R728 B.n842 B.n86 256.663
R729 B.n457 B.n227 256.663
R730 B.n230 B.n227 256.663
R731 B.n450 B.n227 256.663
R732 B.n444 B.n227 256.663
R733 B.n442 B.n227 256.663
R734 B.n436 B.n227 256.663
R735 B.n434 B.n227 256.663
R736 B.n428 B.n227 256.663
R737 B.n426 B.n227 256.663
R738 B.n420 B.n227 256.663
R739 B.n418 B.n227 256.663
R740 B.n412 B.n227 256.663
R741 B.n410 B.n227 256.663
R742 B.n404 B.n227 256.663
R743 B.n402 B.n227 256.663
R744 B.n396 B.n227 256.663
R745 B.n394 B.n227 256.663
R746 B.n388 B.n227 256.663
R747 B.n386 B.n227 256.663
R748 B.n380 B.n227 256.663
R749 B.n252 B.n227 256.663
R750 B.n374 B.n227 256.663
R751 B.n368 B.n227 256.663
R752 B.n366 B.n227 256.663
R753 B.n360 B.n227 256.663
R754 B.n260 B.n227 256.663
R755 B.n354 B.n227 256.663
R756 B.n348 B.n227 256.663
R757 B.n346 B.n227 256.663
R758 B.n340 B.n227 256.663
R759 B.n338 B.n227 256.663
R760 B.n332 B.n227 256.663
R761 B.n330 B.n227 256.663
R762 B.n324 B.n227 256.663
R763 B.n322 B.n227 256.663
R764 B.n316 B.n227 256.663
R765 B.n314 B.n227 256.663
R766 B.n308 B.n227 256.663
R767 B.n306 B.n227 256.663
R768 B.n300 B.n227 256.663
R769 B.n298 B.n227 256.663
R770 B.n292 B.n227 256.663
R771 B.n290 B.n227 256.663
R772 B.n284 B.n227 256.663
R773 B.n282 B.n227 256.663
R774 B.n942 B.n941 256.663
R775 B.n843 B.n841 163.367
R776 B.n839 B.n89 163.367
R777 B.n835 B.n833 163.367
R778 B.n831 B.n91 163.367
R779 B.n827 B.n825 163.367
R780 B.n823 B.n93 163.367
R781 B.n819 B.n817 163.367
R782 B.n815 B.n95 163.367
R783 B.n811 B.n809 163.367
R784 B.n807 B.n97 163.367
R785 B.n803 B.n801 163.367
R786 B.n799 B.n99 163.367
R787 B.n795 B.n793 163.367
R788 B.n791 B.n101 163.367
R789 B.n787 B.n785 163.367
R790 B.n783 B.n103 163.367
R791 B.n779 B.n777 163.367
R792 B.n775 B.n105 163.367
R793 B.n771 B.n769 163.367
R794 B.n767 B.n107 163.367
R795 B.n762 B.n760 163.367
R796 B.n758 B.n111 163.367
R797 B.n754 B.n752 163.367
R798 B.n750 B.n113 163.367
R799 B.n746 B.n744 163.367
R800 B.n742 B.n115 163.367
R801 B.n738 B.n736 163.367
R802 B.n734 B.n120 163.367
R803 B.n730 B.n728 163.367
R804 B.n726 B.n122 163.367
R805 B.n722 B.n720 163.367
R806 B.n718 B.n124 163.367
R807 B.n714 B.n712 163.367
R808 B.n710 B.n126 163.367
R809 B.n706 B.n704 163.367
R810 B.n702 B.n128 163.367
R811 B.n698 B.n696 163.367
R812 B.n694 B.n130 163.367
R813 B.n690 B.n688 163.367
R814 B.n686 B.n132 163.367
R815 B.n682 B.n680 163.367
R816 B.n678 B.n134 163.367
R817 B.n674 B.n672 163.367
R818 B.n670 B.n136 163.367
R819 B.n666 B.n664 163.367
R820 B.n464 B.n224 163.367
R821 B.n468 B.n224 163.367
R822 B.n468 B.n218 163.367
R823 B.n476 B.n218 163.367
R824 B.n476 B.n216 163.367
R825 B.n480 B.n216 163.367
R826 B.n480 B.n211 163.367
R827 B.n489 B.n211 163.367
R828 B.n489 B.n209 163.367
R829 B.n493 B.n209 163.367
R830 B.n493 B.n203 163.367
R831 B.n501 B.n203 163.367
R832 B.n501 B.n201 163.367
R833 B.n505 B.n201 163.367
R834 B.n505 B.n195 163.367
R835 B.n513 B.n195 163.367
R836 B.n513 B.n193 163.367
R837 B.n517 B.n193 163.367
R838 B.n517 B.n187 163.367
R839 B.n525 B.n187 163.367
R840 B.n525 B.n185 163.367
R841 B.n529 B.n185 163.367
R842 B.n529 B.n179 163.367
R843 B.n537 B.n179 163.367
R844 B.n537 B.n177 163.367
R845 B.n541 B.n177 163.367
R846 B.n541 B.n171 163.367
R847 B.n549 B.n171 163.367
R848 B.n549 B.n169 163.367
R849 B.n553 B.n169 163.367
R850 B.n553 B.n163 163.367
R851 B.n561 B.n163 163.367
R852 B.n561 B.n161 163.367
R853 B.n565 B.n161 163.367
R854 B.n565 B.n155 163.367
R855 B.n573 B.n155 163.367
R856 B.n573 B.n153 163.367
R857 B.n577 B.n153 163.367
R858 B.n577 B.n147 163.367
R859 B.n585 B.n147 163.367
R860 B.n585 B.n145 163.367
R861 B.n590 B.n145 163.367
R862 B.n590 B.n139 163.367
R863 B.n598 B.n139 163.367
R864 B.n599 B.n598 163.367
R865 B.n599 B.n5 163.367
R866 B.n6 B.n5 163.367
R867 B.n7 B.n6 163.367
R868 B.n605 B.n7 163.367
R869 B.n606 B.n605 163.367
R870 B.n606 B.n13 163.367
R871 B.n14 B.n13 163.367
R872 B.n15 B.n14 163.367
R873 B.n611 B.n15 163.367
R874 B.n611 B.n20 163.367
R875 B.n21 B.n20 163.367
R876 B.n22 B.n21 163.367
R877 B.n616 B.n22 163.367
R878 B.n616 B.n27 163.367
R879 B.n28 B.n27 163.367
R880 B.n29 B.n28 163.367
R881 B.n621 B.n29 163.367
R882 B.n621 B.n34 163.367
R883 B.n35 B.n34 163.367
R884 B.n36 B.n35 163.367
R885 B.n626 B.n36 163.367
R886 B.n626 B.n41 163.367
R887 B.n42 B.n41 163.367
R888 B.n43 B.n42 163.367
R889 B.n631 B.n43 163.367
R890 B.n631 B.n48 163.367
R891 B.n49 B.n48 163.367
R892 B.n50 B.n49 163.367
R893 B.n636 B.n50 163.367
R894 B.n636 B.n55 163.367
R895 B.n56 B.n55 163.367
R896 B.n57 B.n56 163.367
R897 B.n641 B.n57 163.367
R898 B.n641 B.n62 163.367
R899 B.n63 B.n62 163.367
R900 B.n64 B.n63 163.367
R901 B.n646 B.n64 163.367
R902 B.n646 B.n69 163.367
R903 B.n70 B.n69 163.367
R904 B.n71 B.n70 163.367
R905 B.n651 B.n71 163.367
R906 B.n651 B.n76 163.367
R907 B.n77 B.n76 163.367
R908 B.n78 B.n77 163.367
R909 B.n656 B.n78 163.367
R910 B.n656 B.n83 163.367
R911 B.n84 B.n83 163.367
R912 B.n85 B.n84 163.367
R913 B.n458 B.n456 163.367
R914 B.n456 B.n455 163.367
R915 B.n452 B.n451 163.367
R916 B.n449 B.n232 163.367
R917 B.n445 B.n443 163.367
R918 B.n441 B.n234 163.367
R919 B.n437 B.n435 163.367
R920 B.n433 B.n236 163.367
R921 B.n429 B.n427 163.367
R922 B.n425 B.n238 163.367
R923 B.n421 B.n419 163.367
R924 B.n417 B.n240 163.367
R925 B.n413 B.n411 163.367
R926 B.n409 B.n242 163.367
R927 B.n405 B.n403 163.367
R928 B.n401 B.n244 163.367
R929 B.n397 B.n395 163.367
R930 B.n393 B.n246 163.367
R931 B.n389 B.n387 163.367
R932 B.n385 B.n248 163.367
R933 B.n381 B.n379 163.367
R934 B.n376 B.n375 163.367
R935 B.n373 B.n254 163.367
R936 B.n369 B.n367 163.367
R937 B.n365 B.n256 163.367
R938 B.n361 B.n359 163.367
R939 B.n356 B.n355 163.367
R940 B.n353 B.n262 163.367
R941 B.n349 B.n347 163.367
R942 B.n345 B.n264 163.367
R943 B.n341 B.n339 163.367
R944 B.n337 B.n266 163.367
R945 B.n333 B.n331 163.367
R946 B.n329 B.n268 163.367
R947 B.n325 B.n323 163.367
R948 B.n321 B.n270 163.367
R949 B.n317 B.n315 163.367
R950 B.n313 B.n272 163.367
R951 B.n309 B.n307 163.367
R952 B.n305 B.n274 163.367
R953 B.n301 B.n299 163.367
R954 B.n297 B.n276 163.367
R955 B.n293 B.n291 163.367
R956 B.n289 B.n278 163.367
R957 B.n285 B.n283 163.367
R958 B.n281 B.n226 163.367
R959 B.n462 B.n222 163.367
R960 B.n470 B.n222 163.367
R961 B.n470 B.n220 163.367
R962 B.n474 B.n220 163.367
R963 B.n474 B.n214 163.367
R964 B.n483 B.n214 163.367
R965 B.n483 B.n212 163.367
R966 B.n487 B.n212 163.367
R967 B.n487 B.n207 163.367
R968 B.n495 B.n207 163.367
R969 B.n495 B.n205 163.367
R970 B.n499 B.n205 163.367
R971 B.n499 B.n199 163.367
R972 B.n507 B.n199 163.367
R973 B.n507 B.n197 163.367
R974 B.n511 B.n197 163.367
R975 B.n511 B.n191 163.367
R976 B.n519 B.n191 163.367
R977 B.n519 B.n189 163.367
R978 B.n523 B.n189 163.367
R979 B.n523 B.n183 163.367
R980 B.n531 B.n183 163.367
R981 B.n531 B.n181 163.367
R982 B.n535 B.n181 163.367
R983 B.n535 B.n175 163.367
R984 B.n543 B.n175 163.367
R985 B.n543 B.n173 163.367
R986 B.n547 B.n173 163.367
R987 B.n547 B.n167 163.367
R988 B.n555 B.n167 163.367
R989 B.n555 B.n165 163.367
R990 B.n559 B.n165 163.367
R991 B.n559 B.n159 163.367
R992 B.n567 B.n159 163.367
R993 B.n567 B.n157 163.367
R994 B.n571 B.n157 163.367
R995 B.n571 B.n151 163.367
R996 B.n579 B.n151 163.367
R997 B.n579 B.n149 163.367
R998 B.n583 B.n149 163.367
R999 B.n583 B.n143 163.367
R1000 B.n592 B.n143 163.367
R1001 B.n592 B.n141 163.367
R1002 B.n596 B.n141 163.367
R1003 B.n596 B.n3 163.367
R1004 B.n940 B.n3 163.367
R1005 B.n936 B.n2 163.367
R1006 B.n936 B.n935 163.367
R1007 B.n935 B.n9 163.367
R1008 B.n931 B.n9 163.367
R1009 B.n931 B.n11 163.367
R1010 B.n927 B.n11 163.367
R1011 B.n927 B.n17 163.367
R1012 B.n923 B.n17 163.367
R1013 B.n923 B.n19 163.367
R1014 B.n919 B.n19 163.367
R1015 B.n919 B.n24 163.367
R1016 B.n915 B.n24 163.367
R1017 B.n915 B.n26 163.367
R1018 B.n911 B.n26 163.367
R1019 B.n911 B.n31 163.367
R1020 B.n907 B.n31 163.367
R1021 B.n907 B.n33 163.367
R1022 B.n903 B.n33 163.367
R1023 B.n903 B.n38 163.367
R1024 B.n899 B.n38 163.367
R1025 B.n899 B.n40 163.367
R1026 B.n895 B.n40 163.367
R1027 B.n895 B.n45 163.367
R1028 B.n891 B.n45 163.367
R1029 B.n891 B.n47 163.367
R1030 B.n887 B.n47 163.367
R1031 B.n887 B.n52 163.367
R1032 B.n883 B.n52 163.367
R1033 B.n883 B.n54 163.367
R1034 B.n879 B.n54 163.367
R1035 B.n879 B.n59 163.367
R1036 B.n875 B.n59 163.367
R1037 B.n875 B.n61 163.367
R1038 B.n871 B.n61 163.367
R1039 B.n871 B.n66 163.367
R1040 B.n867 B.n66 163.367
R1041 B.n867 B.n68 163.367
R1042 B.n863 B.n68 163.367
R1043 B.n863 B.n72 163.367
R1044 B.n859 B.n72 163.367
R1045 B.n859 B.n74 163.367
R1046 B.n855 B.n74 163.367
R1047 B.n855 B.n80 163.367
R1048 B.n851 B.n80 163.367
R1049 B.n851 B.n82 163.367
R1050 B.n847 B.n82 163.367
R1051 B.n116 B.t8 137.431
R1052 B.n257 B.t13 137.431
R1053 B.n108 B.t15 137.417
R1054 B.n249 B.t19 137.417
R1055 B.n463 B.n227 87.8978
R1056 B.n848 B.n86 87.8978
R1057 B.n117 B.t9 73.8196
R1058 B.n258 B.t12 73.8196
R1059 B.n109 B.t16 73.8049
R1060 B.n250 B.t18 73.8049
R1061 B.n842 B.n87 71.676
R1062 B.n841 B.n840 71.676
R1063 B.n834 B.n89 71.676
R1064 B.n833 B.n832 71.676
R1065 B.n826 B.n91 71.676
R1066 B.n825 B.n824 71.676
R1067 B.n818 B.n93 71.676
R1068 B.n817 B.n816 71.676
R1069 B.n810 B.n95 71.676
R1070 B.n809 B.n808 71.676
R1071 B.n802 B.n97 71.676
R1072 B.n801 B.n800 71.676
R1073 B.n794 B.n99 71.676
R1074 B.n793 B.n792 71.676
R1075 B.n786 B.n101 71.676
R1076 B.n785 B.n784 71.676
R1077 B.n778 B.n103 71.676
R1078 B.n777 B.n776 71.676
R1079 B.n770 B.n105 71.676
R1080 B.n769 B.n768 71.676
R1081 B.n761 B.n107 71.676
R1082 B.n760 B.n759 71.676
R1083 B.n753 B.n111 71.676
R1084 B.n752 B.n751 71.676
R1085 B.n745 B.n113 71.676
R1086 B.n744 B.n743 71.676
R1087 B.n737 B.n115 71.676
R1088 B.n736 B.n735 71.676
R1089 B.n729 B.n120 71.676
R1090 B.n728 B.n727 71.676
R1091 B.n721 B.n122 71.676
R1092 B.n720 B.n719 71.676
R1093 B.n713 B.n124 71.676
R1094 B.n712 B.n711 71.676
R1095 B.n705 B.n126 71.676
R1096 B.n704 B.n703 71.676
R1097 B.n697 B.n128 71.676
R1098 B.n696 B.n695 71.676
R1099 B.n689 B.n130 71.676
R1100 B.n688 B.n687 71.676
R1101 B.n681 B.n132 71.676
R1102 B.n680 B.n679 71.676
R1103 B.n673 B.n134 71.676
R1104 B.n672 B.n671 71.676
R1105 B.n665 B.n136 71.676
R1106 B.n664 B.n663 71.676
R1107 B.n663 B.n662 71.676
R1108 B.n666 B.n665 71.676
R1109 B.n671 B.n670 71.676
R1110 B.n674 B.n673 71.676
R1111 B.n679 B.n678 71.676
R1112 B.n682 B.n681 71.676
R1113 B.n687 B.n686 71.676
R1114 B.n690 B.n689 71.676
R1115 B.n695 B.n694 71.676
R1116 B.n698 B.n697 71.676
R1117 B.n703 B.n702 71.676
R1118 B.n706 B.n705 71.676
R1119 B.n711 B.n710 71.676
R1120 B.n714 B.n713 71.676
R1121 B.n719 B.n718 71.676
R1122 B.n722 B.n721 71.676
R1123 B.n727 B.n726 71.676
R1124 B.n730 B.n729 71.676
R1125 B.n735 B.n734 71.676
R1126 B.n738 B.n737 71.676
R1127 B.n743 B.n742 71.676
R1128 B.n746 B.n745 71.676
R1129 B.n751 B.n750 71.676
R1130 B.n754 B.n753 71.676
R1131 B.n759 B.n758 71.676
R1132 B.n762 B.n761 71.676
R1133 B.n768 B.n767 71.676
R1134 B.n771 B.n770 71.676
R1135 B.n776 B.n775 71.676
R1136 B.n779 B.n778 71.676
R1137 B.n784 B.n783 71.676
R1138 B.n787 B.n786 71.676
R1139 B.n792 B.n791 71.676
R1140 B.n795 B.n794 71.676
R1141 B.n800 B.n799 71.676
R1142 B.n803 B.n802 71.676
R1143 B.n808 B.n807 71.676
R1144 B.n811 B.n810 71.676
R1145 B.n816 B.n815 71.676
R1146 B.n819 B.n818 71.676
R1147 B.n824 B.n823 71.676
R1148 B.n827 B.n826 71.676
R1149 B.n832 B.n831 71.676
R1150 B.n835 B.n834 71.676
R1151 B.n840 B.n839 71.676
R1152 B.n843 B.n842 71.676
R1153 B.n457 B.n228 71.676
R1154 B.n455 B.n230 71.676
R1155 B.n451 B.n450 71.676
R1156 B.n444 B.n232 71.676
R1157 B.n443 B.n442 71.676
R1158 B.n436 B.n234 71.676
R1159 B.n435 B.n434 71.676
R1160 B.n428 B.n236 71.676
R1161 B.n427 B.n426 71.676
R1162 B.n420 B.n238 71.676
R1163 B.n419 B.n418 71.676
R1164 B.n412 B.n240 71.676
R1165 B.n411 B.n410 71.676
R1166 B.n404 B.n242 71.676
R1167 B.n403 B.n402 71.676
R1168 B.n396 B.n244 71.676
R1169 B.n395 B.n394 71.676
R1170 B.n388 B.n246 71.676
R1171 B.n387 B.n386 71.676
R1172 B.n380 B.n248 71.676
R1173 B.n379 B.n252 71.676
R1174 B.n375 B.n374 71.676
R1175 B.n368 B.n254 71.676
R1176 B.n367 B.n366 71.676
R1177 B.n360 B.n256 71.676
R1178 B.n359 B.n260 71.676
R1179 B.n355 B.n354 71.676
R1180 B.n348 B.n262 71.676
R1181 B.n347 B.n346 71.676
R1182 B.n340 B.n264 71.676
R1183 B.n339 B.n338 71.676
R1184 B.n332 B.n266 71.676
R1185 B.n331 B.n330 71.676
R1186 B.n324 B.n268 71.676
R1187 B.n323 B.n322 71.676
R1188 B.n316 B.n270 71.676
R1189 B.n315 B.n314 71.676
R1190 B.n308 B.n272 71.676
R1191 B.n307 B.n306 71.676
R1192 B.n300 B.n274 71.676
R1193 B.n299 B.n298 71.676
R1194 B.n292 B.n276 71.676
R1195 B.n291 B.n290 71.676
R1196 B.n284 B.n278 71.676
R1197 B.n283 B.n282 71.676
R1198 B.n458 B.n457 71.676
R1199 B.n452 B.n230 71.676
R1200 B.n450 B.n449 71.676
R1201 B.n445 B.n444 71.676
R1202 B.n442 B.n441 71.676
R1203 B.n437 B.n436 71.676
R1204 B.n434 B.n433 71.676
R1205 B.n429 B.n428 71.676
R1206 B.n426 B.n425 71.676
R1207 B.n421 B.n420 71.676
R1208 B.n418 B.n417 71.676
R1209 B.n413 B.n412 71.676
R1210 B.n410 B.n409 71.676
R1211 B.n405 B.n404 71.676
R1212 B.n402 B.n401 71.676
R1213 B.n397 B.n396 71.676
R1214 B.n394 B.n393 71.676
R1215 B.n389 B.n388 71.676
R1216 B.n386 B.n385 71.676
R1217 B.n381 B.n380 71.676
R1218 B.n376 B.n252 71.676
R1219 B.n374 B.n373 71.676
R1220 B.n369 B.n368 71.676
R1221 B.n366 B.n365 71.676
R1222 B.n361 B.n360 71.676
R1223 B.n356 B.n260 71.676
R1224 B.n354 B.n353 71.676
R1225 B.n349 B.n348 71.676
R1226 B.n346 B.n345 71.676
R1227 B.n341 B.n340 71.676
R1228 B.n338 B.n337 71.676
R1229 B.n333 B.n332 71.676
R1230 B.n330 B.n329 71.676
R1231 B.n325 B.n324 71.676
R1232 B.n322 B.n321 71.676
R1233 B.n317 B.n316 71.676
R1234 B.n314 B.n313 71.676
R1235 B.n309 B.n308 71.676
R1236 B.n306 B.n305 71.676
R1237 B.n301 B.n300 71.676
R1238 B.n298 B.n297 71.676
R1239 B.n293 B.n292 71.676
R1240 B.n290 B.n289 71.676
R1241 B.n285 B.n284 71.676
R1242 B.n282 B.n281 71.676
R1243 B.n941 B.n940 71.676
R1244 B.n941 B.n2 71.676
R1245 B.n109 B.n108 63.6126
R1246 B.n117 B.n116 63.6126
R1247 B.n258 B.n257 63.6126
R1248 B.n250 B.n249 63.6126
R1249 B.n764 B.n109 59.5399
R1250 B.n118 B.n117 59.5399
R1251 B.n259 B.n258 59.5399
R1252 B.n251 B.n250 59.5399
R1253 B.n463 B.n223 43.6284
R1254 B.n469 B.n223 43.6284
R1255 B.n469 B.n219 43.6284
R1256 B.n475 B.n219 43.6284
R1257 B.n475 B.n215 43.6284
R1258 B.n482 B.n215 43.6284
R1259 B.n482 B.n481 43.6284
R1260 B.n488 B.n208 43.6284
R1261 B.n494 B.n208 43.6284
R1262 B.n494 B.n204 43.6284
R1263 B.n500 B.n204 43.6284
R1264 B.n500 B.n200 43.6284
R1265 B.n506 B.n200 43.6284
R1266 B.n506 B.n196 43.6284
R1267 B.n512 B.n196 43.6284
R1268 B.n512 B.n192 43.6284
R1269 B.n518 B.n192 43.6284
R1270 B.n518 B.n188 43.6284
R1271 B.n524 B.n188 43.6284
R1272 B.n530 B.n184 43.6284
R1273 B.n530 B.n180 43.6284
R1274 B.n536 B.n180 43.6284
R1275 B.n536 B.n176 43.6284
R1276 B.n542 B.n176 43.6284
R1277 B.n542 B.n172 43.6284
R1278 B.n548 B.n172 43.6284
R1279 B.n548 B.n168 43.6284
R1280 B.n554 B.n168 43.6284
R1281 B.n560 B.n164 43.6284
R1282 B.n560 B.n160 43.6284
R1283 B.n566 B.n160 43.6284
R1284 B.n566 B.n156 43.6284
R1285 B.n572 B.n156 43.6284
R1286 B.n572 B.n152 43.6284
R1287 B.n578 B.n152 43.6284
R1288 B.n578 B.n148 43.6284
R1289 B.n584 B.n148 43.6284
R1290 B.n591 B.n144 43.6284
R1291 B.n591 B.n140 43.6284
R1292 B.n597 B.n140 43.6284
R1293 B.n597 B.n4 43.6284
R1294 B.n939 B.n4 43.6284
R1295 B.n939 B.n938 43.6284
R1296 B.n938 B.n937 43.6284
R1297 B.n937 B.n8 43.6284
R1298 B.n12 B.n8 43.6284
R1299 B.n930 B.n12 43.6284
R1300 B.n930 B.n929 43.6284
R1301 B.n928 B.n16 43.6284
R1302 B.n922 B.n16 43.6284
R1303 B.n922 B.n921 43.6284
R1304 B.n921 B.n920 43.6284
R1305 B.n920 B.n23 43.6284
R1306 B.n914 B.n23 43.6284
R1307 B.n914 B.n913 43.6284
R1308 B.n913 B.n912 43.6284
R1309 B.n912 B.n30 43.6284
R1310 B.n906 B.n905 43.6284
R1311 B.n905 B.n904 43.6284
R1312 B.n904 B.n37 43.6284
R1313 B.n898 B.n37 43.6284
R1314 B.n898 B.n897 43.6284
R1315 B.n897 B.n896 43.6284
R1316 B.n896 B.n44 43.6284
R1317 B.n890 B.n44 43.6284
R1318 B.n890 B.n889 43.6284
R1319 B.n888 B.n51 43.6284
R1320 B.n882 B.n51 43.6284
R1321 B.n882 B.n881 43.6284
R1322 B.n881 B.n880 43.6284
R1323 B.n880 B.n58 43.6284
R1324 B.n874 B.n58 43.6284
R1325 B.n874 B.n873 43.6284
R1326 B.n873 B.n872 43.6284
R1327 B.n872 B.n65 43.6284
R1328 B.n866 B.n65 43.6284
R1329 B.n866 B.n865 43.6284
R1330 B.n865 B.n864 43.6284
R1331 B.n858 B.n75 43.6284
R1332 B.n858 B.n857 43.6284
R1333 B.n857 B.n856 43.6284
R1334 B.n856 B.n79 43.6284
R1335 B.n850 B.n79 43.6284
R1336 B.n850 B.n849 43.6284
R1337 B.n849 B.n848 43.6284
R1338 B.n481 B.t11 40.4204
R1339 B.t2 B.n144 40.4204
R1340 B.n929 B.t1 40.4204
R1341 B.n75 B.t7 40.4204
R1342 B.n461 B.n460 34.8103
R1343 B.n465 B.n225 34.8103
R1344 B.n661 B.n660 34.8103
R1345 B.n846 B.n845 34.8103
R1346 B.n524 B.t5 34.0046
R1347 B.t3 B.n888 34.0046
R1348 B.t4 B.n164 25.0224
R1349 B.t0 B.n30 25.0224
R1350 B.n554 B.t4 18.6065
R1351 B.n906 B.t0 18.6065
R1352 B B.n942 18.0485
R1353 B.n461 B.n221 10.6151
R1354 B.n471 B.n221 10.6151
R1355 B.n472 B.n471 10.6151
R1356 B.n473 B.n472 10.6151
R1357 B.n473 B.n213 10.6151
R1358 B.n484 B.n213 10.6151
R1359 B.n485 B.n484 10.6151
R1360 B.n486 B.n485 10.6151
R1361 B.n486 B.n206 10.6151
R1362 B.n496 B.n206 10.6151
R1363 B.n497 B.n496 10.6151
R1364 B.n498 B.n497 10.6151
R1365 B.n498 B.n198 10.6151
R1366 B.n508 B.n198 10.6151
R1367 B.n509 B.n508 10.6151
R1368 B.n510 B.n509 10.6151
R1369 B.n510 B.n190 10.6151
R1370 B.n520 B.n190 10.6151
R1371 B.n521 B.n520 10.6151
R1372 B.n522 B.n521 10.6151
R1373 B.n522 B.n182 10.6151
R1374 B.n532 B.n182 10.6151
R1375 B.n533 B.n532 10.6151
R1376 B.n534 B.n533 10.6151
R1377 B.n534 B.n174 10.6151
R1378 B.n544 B.n174 10.6151
R1379 B.n545 B.n544 10.6151
R1380 B.n546 B.n545 10.6151
R1381 B.n546 B.n166 10.6151
R1382 B.n556 B.n166 10.6151
R1383 B.n557 B.n556 10.6151
R1384 B.n558 B.n557 10.6151
R1385 B.n558 B.n158 10.6151
R1386 B.n568 B.n158 10.6151
R1387 B.n569 B.n568 10.6151
R1388 B.n570 B.n569 10.6151
R1389 B.n570 B.n150 10.6151
R1390 B.n580 B.n150 10.6151
R1391 B.n581 B.n580 10.6151
R1392 B.n582 B.n581 10.6151
R1393 B.n582 B.n142 10.6151
R1394 B.n593 B.n142 10.6151
R1395 B.n594 B.n593 10.6151
R1396 B.n595 B.n594 10.6151
R1397 B.n595 B.n0 10.6151
R1398 B.n460 B.n459 10.6151
R1399 B.n459 B.n229 10.6151
R1400 B.n454 B.n229 10.6151
R1401 B.n454 B.n453 10.6151
R1402 B.n453 B.n231 10.6151
R1403 B.n448 B.n231 10.6151
R1404 B.n448 B.n447 10.6151
R1405 B.n447 B.n446 10.6151
R1406 B.n446 B.n233 10.6151
R1407 B.n440 B.n233 10.6151
R1408 B.n440 B.n439 10.6151
R1409 B.n439 B.n438 10.6151
R1410 B.n438 B.n235 10.6151
R1411 B.n432 B.n235 10.6151
R1412 B.n432 B.n431 10.6151
R1413 B.n431 B.n430 10.6151
R1414 B.n430 B.n237 10.6151
R1415 B.n424 B.n237 10.6151
R1416 B.n424 B.n423 10.6151
R1417 B.n423 B.n422 10.6151
R1418 B.n422 B.n239 10.6151
R1419 B.n416 B.n239 10.6151
R1420 B.n416 B.n415 10.6151
R1421 B.n415 B.n414 10.6151
R1422 B.n414 B.n241 10.6151
R1423 B.n408 B.n241 10.6151
R1424 B.n408 B.n407 10.6151
R1425 B.n407 B.n406 10.6151
R1426 B.n406 B.n243 10.6151
R1427 B.n400 B.n243 10.6151
R1428 B.n400 B.n399 10.6151
R1429 B.n399 B.n398 10.6151
R1430 B.n398 B.n245 10.6151
R1431 B.n392 B.n245 10.6151
R1432 B.n392 B.n391 10.6151
R1433 B.n391 B.n390 10.6151
R1434 B.n390 B.n247 10.6151
R1435 B.n384 B.n247 10.6151
R1436 B.n384 B.n383 10.6151
R1437 B.n383 B.n382 10.6151
R1438 B.n378 B.n377 10.6151
R1439 B.n377 B.n253 10.6151
R1440 B.n372 B.n253 10.6151
R1441 B.n372 B.n371 10.6151
R1442 B.n371 B.n370 10.6151
R1443 B.n370 B.n255 10.6151
R1444 B.n364 B.n255 10.6151
R1445 B.n364 B.n363 10.6151
R1446 B.n363 B.n362 10.6151
R1447 B.n358 B.n357 10.6151
R1448 B.n357 B.n261 10.6151
R1449 B.n352 B.n261 10.6151
R1450 B.n352 B.n351 10.6151
R1451 B.n351 B.n350 10.6151
R1452 B.n350 B.n263 10.6151
R1453 B.n344 B.n263 10.6151
R1454 B.n344 B.n343 10.6151
R1455 B.n343 B.n342 10.6151
R1456 B.n342 B.n265 10.6151
R1457 B.n336 B.n265 10.6151
R1458 B.n336 B.n335 10.6151
R1459 B.n335 B.n334 10.6151
R1460 B.n334 B.n267 10.6151
R1461 B.n328 B.n267 10.6151
R1462 B.n328 B.n327 10.6151
R1463 B.n327 B.n326 10.6151
R1464 B.n326 B.n269 10.6151
R1465 B.n320 B.n269 10.6151
R1466 B.n320 B.n319 10.6151
R1467 B.n319 B.n318 10.6151
R1468 B.n318 B.n271 10.6151
R1469 B.n312 B.n271 10.6151
R1470 B.n312 B.n311 10.6151
R1471 B.n311 B.n310 10.6151
R1472 B.n310 B.n273 10.6151
R1473 B.n304 B.n273 10.6151
R1474 B.n304 B.n303 10.6151
R1475 B.n303 B.n302 10.6151
R1476 B.n302 B.n275 10.6151
R1477 B.n296 B.n275 10.6151
R1478 B.n296 B.n295 10.6151
R1479 B.n295 B.n294 10.6151
R1480 B.n294 B.n277 10.6151
R1481 B.n288 B.n277 10.6151
R1482 B.n288 B.n287 10.6151
R1483 B.n287 B.n286 10.6151
R1484 B.n286 B.n279 10.6151
R1485 B.n280 B.n279 10.6151
R1486 B.n280 B.n225 10.6151
R1487 B.n466 B.n465 10.6151
R1488 B.n467 B.n466 10.6151
R1489 B.n467 B.n217 10.6151
R1490 B.n477 B.n217 10.6151
R1491 B.n478 B.n477 10.6151
R1492 B.n479 B.n478 10.6151
R1493 B.n479 B.n210 10.6151
R1494 B.n490 B.n210 10.6151
R1495 B.n491 B.n490 10.6151
R1496 B.n492 B.n491 10.6151
R1497 B.n492 B.n202 10.6151
R1498 B.n502 B.n202 10.6151
R1499 B.n503 B.n502 10.6151
R1500 B.n504 B.n503 10.6151
R1501 B.n504 B.n194 10.6151
R1502 B.n514 B.n194 10.6151
R1503 B.n515 B.n514 10.6151
R1504 B.n516 B.n515 10.6151
R1505 B.n516 B.n186 10.6151
R1506 B.n526 B.n186 10.6151
R1507 B.n527 B.n526 10.6151
R1508 B.n528 B.n527 10.6151
R1509 B.n528 B.n178 10.6151
R1510 B.n538 B.n178 10.6151
R1511 B.n539 B.n538 10.6151
R1512 B.n540 B.n539 10.6151
R1513 B.n540 B.n170 10.6151
R1514 B.n550 B.n170 10.6151
R1515 B.n551 B.n550 10.6151
R1516 B.n552 B.n551 10.6151
R1517 B.n552 B.n162 10.6151
R1518 B.n562 B.n162 10.6151
R1519 B.n563 B.n562 10.6151
R1520 B.n564 B.n563 10.6151
R1521 B.n564 B.n154 10.6151
R1522 B.n574 B.n154 10.6151
R1523 B.n575 B.n574 10.6151
R1524 B.n576 B.n575 10.6151
R1525 B.n576 B.n146 10.6151
R1526 B.n586 B.n146 10.6151
R1527 B.n587 B.n586 10.6151
R1528 B.n589 B.n587 10.6151
R1529 B.n589 B.n588 10.6151
R1530 B.n588 B.n138 10.6151
R1531 B.n600 B.n138 10.6151
R1532 B.n601 B.n600 10.6151
R1533 B.n602 B.n601 10.6151
R1534 B.n603 B.n602 10.6151
R1535 B.n604 B.n603 10.6151
R1536 B.n607 B.n604 10.6151
R1537 B.n608 B.n607 10.6151
R1538 B.n609 B.n608 10.6151
R1539 B.n610 B.n609 10.6151
R1540 B.n612 B.n610 10.6151
R1541 B.n613 B.n612 10.6151
R1542 B.n614 B.n613 10.6151
R1543 B.n615 B.n614 10.6151
R1544 B.n617 B.n615 10.6151
R1545 B.n618 B.n617 10.6151
R1546 B.n619 B.n618 10.6151
R1547 B.n620 B.n619 10.6151
R1548 B.n622 B.n620 10.6151
R1549 B.n623 B.n622 10.6151
R1550 B.n624 B.n623 10.6151
R1551 B.n625 B.n624 10.6151
R1552 B.n627 B.n625 10.6151
R1553 B.n628 B.n627 10.6151
R1554 B.n629 B.n628 10.6151
R1555 B.n630 B.n629 10.6151
R1556 B.n632 B.n630 10.6151
R1557 B.n633 B.n632 10.6151
R1558 B.n634 B.n633 10.6151
R1559 B.n635 B.n634 10.6151
R1560 B.n637 B.n635 10.6151
R1561 B.n638 B.n637 10.6151
R1562 B.n639 B.n638 10.6151
R1563 B.n640 B.n639 10.6151
R1564 B.n642 B.n640 10.6151
R1565 B.n643 B.n642 10.6151
R1566 B.n644 B.n643 10.6151
R1567 B.n645 B.n644 10.6151
R1568 B.n647 B.n645 10.6151
R1569 B.n648 B.n647 10.6151
R1570 B.n649 B.n648 10.6151
R1571 B.n650 B.n649 10.6151
R1572 B.n652 B.n650 10.6151
R1573 B.n653 B.n652 10.6151
R1574 B.n654 B.n653 10.6151
R1575 B.n655 B.n654 10.6151
R1576 B.n657 B.n655 10.6151
R1577 B.n658 B.n657 10.6151
R1578 B.n659 B.n658 10.6151
R1579 B.n660 B.n659 10.6151
R1580 B.n934 B.n1 10.6151
R1581 B.n934 B.n933 10.6151
R1582 B.n933 B.n932 10.6151
R1583 B.n932 B.n10 10.6151
R1584 B.n926 B.n10 10.6151
R1585 B.n926 B.n925 10.6151
R1586 B.n925 B.n924 10.6151
R1587 B.n924 B.n18 10.6151
R1588 B.n918 B.n18 10.6151
R1589 B.n918 B.n917 10.6151
R1590 B.n917 B.n916 10.6151
R1591 B.n916 B.n25 10.6151
R1592 B.n910 B.n25 10.6151
R1593 B.n910 B.n909 10.6151
R1594 B.n909 B.n908 10.6151
R1595 B.n908 B.n32 10.6151
R1596 B.n902 B.n32 10.6151
R1597 B.n902 B.n901 10.6151
R1598 B.n901 B.n900 10.6151
R1599 B.n900 B.n39 10.6151
R1600 B.n894 B.n39 10.6151
R1601 B.n894 B.n893 10.6151
R1602 B.n893 B.n892 10.6151
R1603 B.n892 B.n46 10.6151
R1604 B.n886 B.n46 10.6151
R1605 B.n886 B.n885 10.6151
R1606 B.n885 B.n884 10.6151
R1607 B.n884 B.n53 10.6151
R1608 B.n878 B.n53 10.6151
R1609 B.n878 B.n877 10.6151
R1610 B.n877 B.n876 10.6151
R1611 B.n876 B.n60 10.6151
R1612 B.n870 B.n60 10.6151
R1613 B.n870 B.n869 10.6151
R1614 B.n869 B.n868 10.6151
R1615 B.n868 B.n67 10.6151
R1616 B.n862 B.n67 10.6151
R1617 B.n862 B.n861 10.6151
R1618 B.n861 B.n860 10.6151
R1619 B.n860 B.n73 10.6151
R1620 B.n854 B.n73 10.6151
R1621 B.n854 B.n853 10.6151
R1622 B.n853 B.n852 10.6151
R1623 B.n852 B.n81 10.6151
R1624 B.n846 B.n81 10.6151
R1625 B.n845 B.n844 10.6151
R1626 B.n844 B.n88 10.6151
R1627 B.n838 B.n88 10.6151
R1628 B.n838 B.n837 10.6151
R1629 B.n837 B.n836 10.6151
R1630 B.n836 B.n90 10.6151
R1631 B.n830 B.n90 10.6151
R1632 B.n830 B.n829 10.6151
R1633 B.n829 B.n828 10.6151
R1634 B.n828 B.n92 10.6151
R1635 B.n822 B.n92 10.6151
R1636 B.n822 B.n821 10.6151
R1637 B.n821 B.n820 10.6151
R1638 B.n820 B.n94 10.6151
R1639 B.n814 B.n94 10.6151
R1640 B.n814 B.n813 10.6151
R1641 B.n813 B.n812 10.6151
R1642 B.n812 B.n96 10.6151
R1643 B.n806 B.n96 10.6151
R1644 B.n806 B.n805 10.6151
R1645 B.n805 B.n804 10.6151
R1646 B.n804 B.n98 10.6151
R1647 B.n798 B.n98 10.6151
R1648 B.n798 B.n797 10.6151
R1649 B.n797 B.n796 10.6151
R1650 B.n796 B.n100 10.6151
R1651 B.n790 B.n100 10.6151
R1652 B.n790 B.n789 10.6151
R1653 B.n789 B.n788 10.6151
R1654 B.n788 B.n102 10.6151
R1655 B.n782 B.n102 10.6151
R1656 B.n782 B.n781 10.6151
R1657 B.n781 B.n780 10.6151
R1658 B.n780 B.n104 10.6151
R1659 B.n774 B.n104 10.6151
R1660 B.n774 B.n773 10.6151
R1661 B.n773 B.n772 10.6151
R1662 B.n772 B.n106 10.6151
R1663 B.n766 B.n106 10.6151
R1664 B.n766 B.n765 10.6151
R1665 B.n763 B.n110 10.6151
R1666 B.n757 B.n110 10.6151
R1667 B.n757 B.n756 10.6151
R1668 B.n756 B.n755 10.6151
R1669 B.n755 B.n112 10.6151
R1670 B.n749 B.n112 10.6151
R1671 B.n749 B.n748 10.6151
R1672 B.n748 B.n747 10.6151
R1673 B.n747 B.n114 10.6151
R1674 B.n741 B.n740 10.6151
R1675 B.n740 B.n739 10.6151
R1676 B.n739 B.n119 10.6151
R1677 B.n733 B.n119 10.6151
R1678 B.n733 B.n732 10.6151
R1679 B.n732 B.n731 10.6151
R1680 B.n731 B.n121 10.6151
R1681 B.n725 B.n121 10.6151
R1682 B.n725 B.n724 10.6151
R1683 B.n724 B.n723 10.6151
R1684 B.n723 B.n123 10.6151
R1685 B.n717 B.n123 10.6151
R1686 B.n717 B.n716 10.6151
R1687 B.n716 B.n715 10.6151
R1688 B.n715 B.n125 10.6151
R1689 B.n709 B.n125 10.6151
R1690 B.n709 B.n708 10.6151
R1691 B.n708 B.n707 10.6151
R1692 B.n707 B.n127 10.6151
R1693 B.n701 B.n127 10.6151
R1694 B.n701 B.n700 10.6151
R1695 B.n700 B.n699 10.6151
R1696 B.n699 B.n129 10.6151
R1697 B.n693 B.n129 10.6151
R1698 B.n693 B.n692 10.6151
R1699 B.n692 B.n691 10.6151
R1700 B.n691 B.n131 10.6151
R1701 B.n685 B.n131 10.6151
R1702 B.n685 B.n684 10.6151
R1703 B.n684 B.n683 10.6151
R1704 B.n683 B.n133 10.6151
R1705 B.n677 B.n133 10.6151
R1706 B.n677 B.n676 10.6151
R1707 B.n676 B.n675 10.6151
R1708 B.n675 B.n135 10.6151
R1709 B.n669 B.n135 10.6151
R1710 B.n669 B.n668 10.6151
R1711 B.n668 B.n667 10.6151
R1712 B.n667 B.n137 10.6151
R1713 B.n661 B.n137 10.6151
R1714 B.t5 B.n184 9.6243
R1715 B.n889 B.t3 9.6243
R1716 B.n382 B.n251 9.36635
R1717 B.n358 B.n259 9.36635
R1718 B.n765 B.n764 9.36635
R1719 B.n741 B.n118 9.36635
R1720 B.n942 B.n0 8.11757
R1721 B.n942 B.n1 8.11757
R1722 B.n488 B.t11 3.20843
R1723 B.n584 B.t2 3.20843
R1724 B.t1 B.n928 3.20843
R1725 B.n864 B.t7 3.20843
R1726 B.n378 B.n251 1.24928
R1727 B.n362 B.n259 1.24928
R1728 B.n764 B.n763 1.24928
R1729 B.n118 B.n114 1.24928
R1730 VN.n33 VN.n18 161.3
R1731 VN.n32 VN.n31 161.3
R1732 VN.n30 VN.n19 161.3
R1733 VN.n29 VN.n28 161.3
R1734 VN.n27 VN.n20 161.3
R1735 VN.n26 VN.n25 161.3
R1736 VN.n24 VN.n21 161.3
R1737 VN.n15 VN.n0 161.3
R1738 VN.n14 VN.n13 161.3
R1739 VN.n12 VN.n1 161.3
R1740 VN.n11 VN.n10 161.3
R1741 VN.n9 VN.n2 161.3
R1742 VN.n8 VN.n7 161.3
R1743 VN.n6 VN.n3 161.3
R1744 VN.n5 VN.t1 129.436
R1745 VN.n23 VN.t2 129.436
R1746 VN.n17 VN.n16 109.288
R1747 VN.n35 VN.n34 109.288
R1748 VN.n4 VN.t4 96.9724
R1749 VN.n16 VN.t0 96.9724
R1750 VN.n22 VN.t3 96.9724
R1751 VN.n34 VN.t5 96.9724
R1752 VN.n5 VN.n4 61.6325
R1753 VN.n23 VN.n22 61.6325
R1754 VN.n10 VN.n9 51.1773
R1755 VN.n28 VN.n27 51.1773
R1756 VN VN.n35 50.2027
R1757 VN.n10 VN.n1 29.8095
R1758 VN.n28 VN.n19 29.8095
R1759 VN.n8 VN.n3 24.4675
R1760 VN.n9 VN.n8 24.4675
R1761 VN.n14 VN.n1 24.4675
R1762 VN.n15 VN.n14 24.4675
R1763 VN.n27 VN.n26 24.4675
R1764 VN.n26 VN.n21 24.4675
R1765 VN.n33 VN.n32 24.4675
R1766 VN.n32 VN.n19 24.4675
R1767 VN.n4 VN.n3 12.234
R1768 VN.n22 VN.n21 12.234
R1769 VN.n24 VN.n23 5.14959
R1770 VN.n6 VN.n5 5.14959
R1771 VN.n16 VN.n15 1.46852
R1772 VN.n34 VN.n33 1.46852
R1773 VN.n35 VN.n18 0.278367
R1774 VN.n17 VN.n0 0.278367
R1775 VN.n31 VN.n18 0.189894
R1776 VN.n31 VN.n30 0.189894
R1777 VN.n30 VN.n29 0.189894
R1778 VN.n29 VN.n20 0.189894
R1779 VN.n25 VN.n20 0.189894
R1780 VN.n25 VN.n24 0.189894
R1781 VN.n7 VN.n6 0.189894
R1782 VN.n7 VN.n2 0.189894
R1783 VN.n11 VN.n2 0.189894
R1784 VN.n12 VN.n11 0.189894
R1785 VN.n13 VN.n12 0.189894
R1786 VN.n13 VN.n0 0.189894
R1787 VN VN.n17 0.153454
R1788 VDD2.n1 VDD2.t4 67.8465
R1789 VDD2.n2 VDD2.t0 65.7814
R1790 VDD2.n1 VDD2.n0 64.7647
R1791 VDD2 VDD2.n3 64.7619
R1792 VDD2.n2 VDD2.n1 43.1377
R1793 VDD2 VDD2.n2 2.17938
R1794 VDD2.n3 VDD2.t2 1.66857
R1795 VDD2.n3 VDD2.t3 1.66857
R1796 VDD2.n0 VDD2.t1 1.66857
R1797 VDD2.n0 VDD2.t5 1.66857
C0 VDD2 VP 0.487963f
C1 VDD1 VTAIL 7.76793f
C2 VN VP 7.24176f
C3 VDD1 VP 7.14175f
C4 VTAIL VP 7.073f
C5 VN VDD2 6.80808f
C6 VDD1 VDD2 1.5433f
C7 VDD1 VN 0.151198f
C8 VDD2 VTAIL 7.82148f
C9 VN VTAIL 7.05874f
C10 VDD2 B 6.228357f
C11 VDD1 B 6.568814f
C12 VTAIL B 7.99783f
C13 VN B 13.88596f
C14 VP B 12.553531f
C15 VDD2.t4 B 2.28618f
C16 VDD2.t1 B 0.200046f
C17 VDD2.t5 B 0.200046f
C18 VDD2.n0 B 1.78728f
C19 VDD2.n1 B 2.59794f
C20 VDD2.t0 B 2.27463f
C21 VDD2.n2 B 2.45425f
C22 VDD2.t2 B 0.200046f
C23 VDD2.t3 B 0.200046f
C24 VDD2.n3 B 1.78725f
C25 VN.n0 B 0.028365f
C26 VN.t0 B 2.05201f
C27 VN.n1 B 0.042864f
C28 VN.n2 B 0.021515f
C29 VN.n3 B 0.0302f
C30 VN.t1 B 2.27054f
C31 VN.t4 B 2.05201f
C32 VN.n4 B 0.791368f
C33 VN.n5 B 0.763719f
C34 VN.n6 B 0.229433f
C35 VN.n7 B 0.021515f
C36 VN.n8 B 0.040098f
C37 VN.n9 B 0.039063f
C38 VN.n10 B 0.020986f
C39 VN.n11 B 0.021515f
C40 VN.n12 B 0.021515f
C41 VN.n13 B 0.021515f
C42 VN.n14 B 0.040098f
C43 VN.n15 B 0.021489f
C44 VN.n16 B 0.79562f
C45 VN.n17 B 0.042099f
C46 VN.n18 B 0.028365f
C47 VN.t5 B 2.05201f
C48 VN.n19 B 0.042864f
C49 VN.n20 B 0.021515f
C50 VN.n21 B 0.0302f
C51 VN.t2 B 2.27054f
C52 VN.t3 B 2.05201f
C53 VN.n22 B 0.791368f
C54 VN.n23 B 0.763719f
C55 VN.n24 B 0.229433f
C56 VN.n25 B 0.021515f
C57 VN.n26 B 0.040098f
C58 VN.n27 B 0.039063f
C59 VN.n28 B 0.020986f
C60 VN.n29 B 0.021515f
C61 VN.n30 B 0.021515f
C62 VN.n31 B 0.021515f
C63 VN.n32 B 0.040098f
C64 VN.n33 B 0.021489f
C65 VN.n34 B 0.79562f
C66 VN.n35 B 1.21325f
C67 VDD1.t0 B 2.32151f
C68 VDD1.t5 B 2.32064f
C69 VDD1.t1 B 0.203061f
C70 VDD1.t4 B 0.203061f
C71 VDD1.n0 B 1.81422f
C72 VDD1.n1 B 2.75244f
C73 VDD1.t2 B 0.203061f
C74 VDD1.t3 B 0.203061f
C75 VDD1.n2 B 1.80989f
C76 VDD1.n3 B 2.49157f
C77 VTAIL.t1 B 0.225618f
C78 VTAIL.t0 B 0.225618f
C79 VTAIL.n0 B 1.94328f
C80 VTAIL.n1 B 0.437315f
C81 VTAIL.t8 B 2.47934f
C82 VTAIL.n2 B 0.676422f
C83 VTAIL.t10 B 0.225618f
C84 VTAIL.t11 B 0.225618f
C85 VTAIL.n3 B 1.94328f
C86 VTAIL.n4 B 2.00929f
C87 VTAIL.t5 B 0.225618f
C88 VTAIL.t4 B 0.225618f
C89 VTAIL.n5 B 1.94328f
C90 VTAIL.n6 B 2.00929f
C91 VTAIL.t2 B 2.47935f
C92 VTAIL.n7 B 0.676416f
C93 VTAIL.t7 B 0.225618f
C94 VTAIL.t6 B 0.225618f
C95 VTAIL.n8 B 1.94328f
C96 VTAIL.n9 B 0.597161f
C97 VTAIL.t9 B 2.47934f
C98 VTAIL.n10 B 1.8694f
C99 VTAIL.t3 B 2.47934f
C100 VTAIL.n11 B 1.8101f
C101 VP.n0 B 0.02881f
C102 VP.t1 B 2.08418f
C103 VP.n1 B 0.043536f
C104 VP.n2 B 0.021852f
C105 VP.n3 B 0.030673f
C106 VP.n4 B 0.021852f
C107 VP.n5 B 0.021315f
C108 VP.n6 B 0.021852f
C109 VP.t0 B 2.08418f
C110 VP.n7 B 0.80809f
C111 VP.n8 B 0.02881f
C112 VP.t2 B 2.08418f
C113 VP.n9 B 0.043536f
C114 VP.n10 B 0.021852f
C115 VP.n11 B 0.030673f
C116 VP.t5 B 2.30612f
C117 VP.t3 B 2.08418f
C118 VP.n12 B 0.803772f
C119 VP.n13 B 0.77569f
C120 VP.n14 B 0.23303f
C121 VP.n15 B 0.021852f
C122 VP.n16 B 0.040727f
C123 VP.n17 B 0.039675f
C124 VP.n18 B 0.021315f
C125 VP.n19 B 0.021852f
C126 VP.n20 B 0.021852f
C127 VP.n21 B 0.021852f
C128 VP.n22 B 0.040727f
C129 VP.n23 B 0.021826f
C130 VP.n24 B 0.80809f
C131 VP.n25 B 1.22053f
C132 VP.n26 B 1.23626f
C133 VP.n27 B 0.02881f
C134 VP.n28 B 0.021826f
C135 VP.n29 B 0.040727f
C136 VP.n30 B 0.043536f
C137 VP.n31 B 0.021852f
C138 VP.n32 B 0.021852f
C139 VP.n33 B 0.021852f
C140 VP.n34 B 0.039675f
C141 VP.n35 B 0.040727f
C142 VP.t4 B 2.08418f
C143 VP.n36 B 0.734906f
C144 VP.n37 B 0.030673f
C145 VP.n38 B 0.021852f
C146 VP.n39 B 0.021852f
C147 VP.n40 B 0.021852f
C148 VP.n41 B 0.040727f
C149 VP.n42 B 0.039675f
C150 VP.n43 B 0.021315f
C151 VP.n44 B 0.021852f
C152 VP.n45 B 0.021852f
C153 VP.n46 B 0.021852f
C154 VP.n47 B 0.040727f
C155 VP.n48 B 0.021826f
C156 VP.n49 B 0.80809f
C157 VP.n50 B 0.042759f
.ends

