* NGSPICE file created from diff_pair_sample_0053.ext - technology: sky130A

.subckt diff_pair_sample_0053 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=0 ps=0 w=8.65 l=0.93
X1 VDD1.t5 VP.t0 VTAIL.t9 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=1.42725 ps=8.98 w=8.65 l=0.93
X2 B.t8 B.t6 B.t7 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=0 ps=0 w=8.65 l=0.93
X3 VDD1.t4 VP.t1 VTAIL.t6 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=1.42725 ps=8.98 w=8.65 l=0.93
X4 VDD2.t5 VN.t0 VTAIL.t5 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=3.3735 ps=18.08 w=8.65 l=0.93
X5 VDD1.t3 VP.t2 VTAIL.t8 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=3.3735 ps=18.08 w=8.65 l=0.93
X6 VTAIL.t4 VN.t1 VDD2.t4 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=1.42725 ps=8.98 w=8.65 l=0.93
X7 VDD2.t3 VN.t2 VTAIL.t0 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=1.42725 ps=8.98 w=8.65 l=0.93
X8 VDD2.t2 VN.t3 VTAIL.t1 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=3.3735 ps=18.08 w=8.65 l=0.93
X9 VDD2.t1 VN.t4 VTAIL.t2 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=1.42725 ps=8.98 w=8.65 l=0.93
X10 B.t5 B.t3 B.t4 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=0 ps=0 w=8.65 l=0.93
X11 VDD1.t2 VP.t3 VTAIL.t7 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=3.3735 ps=18.08 w=8.65 l=0.93
X12 VTAIL.t11 VP.t4 VDD1.t1 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=1.42725 ps=8.98 w=8.65 l=0.93
X13 VTAIL.t10 VP.t5 VDD1.t0 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=1.42725 ps=8.98 w=8.65 l=0.93
X14 B.t2 B.t0 B.t1 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=3.3735 pd=18.08 as=0 ps=0 w=8.65 l=0.93
X15 VTAIL.t3 VN.t5 VDD2.t0 w_n1978_n2698# sky130_fd_pr__pfet_01v8 ad=1.42725 pd=8.98 as=1.42725 ps=8.98 w=8.65 l=0.93
R0 B.n345 B.n54 585
R1 B.n347 B.n346 585
R2 B.n348 B.n53 585
R3 B.n350 B.n349 585
R4 B.n351 B.n52 585
R5 B.n353 B.n352 585
R6 B.n354 B.n51 585
R7 B.n356 B.n355 585
R8 B.n357 B.n50 585
R9 B.n359 B.n358 585
R10 B.n360 B.n49 585
R11 B.n362 B.n361 585
R12 B.n363 B.n48 585
R13 B.n365 B.n364 585
R14 B.n366 B.n47 585
R15 B.n368 B.n367 585
R16 B.n369 B.n46 585
R17 B.n371 B.n370 585
R18 B.n372 B.n45 585
R19 B.n374 B.n373 585
R20 B.n375 B.n44 585
R21 B.n377 B.n376 585
R22 B.n378 B.n43 585
R23 B.n380 B.n379 585
R24 B.n381 B.n42 585
R25 B.n383 B.n382 585
R26 B.n384 B.n41 585
R27 B.n386 B.n385 585
R28 B.n387 B.n40 585
R29 B.n389 B.n388 585
R30 B.n390 B.n39 585
R31 B.n392 B.n391 585
R32 B.n394 B.n393 585
R33 B.n395 B.n35 585
R34 B.n397 B.n396 585
R35 B.n398 B.n34 585
R36 B.n400 B.n399 585
R37 B.n401 B.n33 585
R38 B.n403 B.n402 585
R39 B.n404 B.n32 585
R40 B.n406 B.n405 585
R41 B.n408 B.n29 585
R42 B.n410 B.n409 585
R43 B.n411 B.n28 585
R44 B.n413 B.n412 585
R45 B.n414 B.n27 585
R46 B.n416 B.n415 585
R47 B.n417 B.n26 585
R48 B.n419 B.n418 585
R49 B.n420 B.n25 585
R50 B.n422 B.n421 585
R51 B.n423 B.n24 585
R52 B.n425 B.n424 585
R53 B.n426 B.n23 585
R54 B.n428 B.n427 585
R55 B.n429 B.n22 585
R56 B.n431 B.n430 585
R57 B.n432 B.n21 585
R58 B.n434 B.n433 585
R59 B.n435 B.n20 585
R60 B.n437 B.n436 585
R61 B.n438 B.n19 585
R62 B.n440 B.n439 585
R63 B.n441 B.n18 585
R64 B.n443 B.n442 585
R65 B.n444 B.n17 585
R66 B.n446 B.n445 585
R67 B.n447 B.n16 585
R68 B.n449 B.n448 585
R69 B.n450 B.n15 585
R70 B.n452 B.n451 585
R71 B.n453 B.n14 585
R72 B.n455 B.n454 585
R73 B.n344 B.n343 585
R74 B.n342 B.n55 585
R75 B.n341 B.n340 585
R76 B.n339 B.n56 585
R77 B.n338 B.n337 585
R78 B.n336 B.n57 585
R79 B.n335 B.n334 585
R80 B.n333 B.n58 585
R81 B.n332 B.n331 585
R82 B.n330 B.n59 585
R83 B.n329 B.n328 585
R84 B.n327 B.n60 585
R85 B.n326 B.n325 585
R86 B.n324 B.n61 585
R87 B.n323 B.n322 585
R88 B.n321 B.n62 585
R89 B.n320 B.n319 585
R90 B.n318 B.n63 585
R91 B.n317 B.n316 585
R92 B.n315 B.n64 585
R93 B.n314 B.n313 585
R94 B.n312 B.n65 585
R95 B.n311 B.n310 585
R96 B.n309 B.n66 585
R97 B.n308 B.n307 585
R98 B.n306 B.n67 585
R99 B.n305 B.n304 585
R100 B.n303 B.n68 585
R101 B.n302 B.n301 585
R102 B.n300 B.n69 585
R103 B.n299 B.n298 585
R104 B.n297 B.n70 585
R105 B.n296 B.n295 585
R106 B.n294 B.n71 585
R107 B.n293 B.n292 585
R108 B.n291 B.n72 585
R109 B.n290 B.n289 585
R110 B.n288 B.n73 585
R111 B.n287 B.n286 585
R112 B.n285 B.n74 585
R113 B.n284 B.n283 585
R114 B.n282 B.n75 585
R115 B.n281 B.n280 585
R116 B.n279 B.n76 585
R117 B.n278 B.n277 585
R118 B.n276 B.n77 585
R119 B.n275 B.n274 585
R120 B.n164 B.n163 585
R121 B.n165 B.n118 585
R122 B.n167 B.n166 585
R123 B.n168 B.n117 585
R124 B.n170 B.n169 585
R125 B.n171 B.n116 585
R126 B.n173 B.n172 585
R127 B.n174 B.n115 585
R128 B.n176 B.n175 585
R129 B.n177 B.n114 585
R130 B.n179 B.n178 585
R131 B.n180 B.n113 585
R132 B.n182 B.n181 585
R133 B.n183 B.n112 585
R134 B.n185 B.n184 585
R135 B.n186 B.n111 585
R136 B.n188 B.n187 585
R137 B.n189 B.n110 585
R138 B.n191 B.n190 585
R139 B.n192 B.n109 585
R140 B.n194 B.n193 585
R141 B.n195 B.n108 585
R142 B.n197 B.n196 585
R143 B.n198 B.n107 585
R144 B.n200 B.n199 585
R145 B.n201 B.n106 585
R146 B.n203 B.n202 585
R147 B.n204 B.n105 585
R148 B.n206 B.n205 585
R149 B.n207 B.n104 585
R150 B.n209 B.n208 585
R151 B.n210 B.n101 585
R152 B.n213 B.n212 585
R153 B.n214 B.n100 585
R154 B.n216 B.n215 585
R155 B.n217 B.n99 585
R156 B.n219 B.n218 585
R157 B.n220 B.n98 585
R158 B.n222 B.n221 585
R159 B.n223 B.n97 585
R160 B.n225 B.n224 585
R161 B.n227 B.n226 585
R162 B.n228 B.n93 585
R163 B.n230 B.n229 585
R164 B.n231 B.n92 585
R165 B.n233 B.n232 585
R166 B.n234 B.n91 585
R167 B.n236 B.n235 585
R168 B.n237 B.n90 585
R169 B.n239 B.n238 585
R170 B.n240 B.n89 585
R171 B.n242 B.n241 585
R172 B.n243 B.n88 585
R173 B.n245 B.n244 585
R174 B.n246 B.n87 585
R175 B.n248 B.n247 585
R176 B.n249 B.n86 585
R177 B.n251 B.n250 585
R178 B.n252 B.n85 585
R179 B.n254 B.n253 585
R180 B.n255 B.n84 585
R181 B.n257 B.n256 585
R182 B.n258 B.n83 585
R183 B.n260 B.n259 585
R184 B.n261 B.n82 585
R185 B.n263 B.n262 585
R186 B.n264 B.n81 585
R187 B.n266 B.n265 585
R188 B.n267 B.n80 585
R189 B.n269 B.n268 585
R190 B.n270 B.n79 585
R191 B.n272 B.n271 585
R192 B.n273 B.n78 585
R193 B.n162 B.n119 585
R194 B.n161 B.n160 585
R195 B.n159 B.n120 585
R196 B.n158 B.n157 585
R197 B.n156 B.n121 585
R198 B.n155 B.n154 585
R199 B.n153 B.n122 585
R200 B.n152 B.n151 585
R201 B.n150 B.n123 585
R202 B.n149 B.n148 585
R203 B.n147 B.n124 585
R204 B.n146 B.n145 585
R205 B.n144 B.n125 585
R206 B.n143 B.n142 585
R207 B.n141 B.n126 585
R208 B.n140 B.n139 585
R209 B.n138 B.n127 585
R210 B.n137 B.n136 585
R211 B.n135 B.n128 585
R212 B.n134 B.n133 585
R213 B.n132 B.n129 585
R214 B.n131 B.n130 585
R215 B.n2 B.n0 585
R216 B.n489 B.n1 585
R217 B.n488 B.n487 585
R218 B.n486 B.n3 585
R219 B.n485 B.n484 585
R220 B.n483 B.n4 585
R221 B.n482 B.n481 585
R222 B.n480 B.n5 585
R223 B.n479 B.n478 585
R224 B.n477 B.n6 585
R225 B.n476 B.n475 585
R226 B.n474 B.n7 585
R227 B.n473 B.n472 585
R228 B.n471 B.n8 585
R229 B.n470 B.n469 585
R230 B.n468 B.n9 585
R231 B.n467 B.n466 585
R232 B.n465 B.n10 585
R233 B.n464 B.n463 585
R234 B.n462 B.n11 585
R235 B.n461 B.n460 585
R236 B.n459 B.n12 585
R237 B.n458 B.n457 585
R238 B.n456 B.n13 585
R239 B.n491 B.n490 585
R240 B.n164 B.n119 497.305
R241 B.n454 B.n13 497.305
R242 B.n274 B.n273 497.305
R243 B.n345 B.n344 497.305
R244 B.n94 B.t6 426.584
R245 B.n102 B.t9 426.584
R246 B.n30 B.t3 426.584
R247 B.n36 B.t0 426.584
R248 B.n94 B.t8 339.75
R249 B.n36 B.t1 339.75
R250 B.n102 B.t11 339.75
R251 B.n30 B.t4 339.75
R252 B.n95 B.t7 315.312
R253 B.n37 B.t2 315.312
R254 B.n103 B.t10 315.312
R255 B.n31 B.t5 315.312
R256 B.n160 B.n119 163.367
R257 B.n160 B.n159 163.367
R258 B.n159 B.n158 163.367
R259 B.n158 B.n121 163.367
R260 B.n154 B.n121 163.367
R261 B.n154 B.n153 163.367
R262 B.n153 B.n152 163.367
R263 B.n152 B.n123 163.367
R264 B.n148 B.n123 163.367
R265 B.n148 B.n147 163.367
R266 B.n147 B.n146 163.367
R267 B.n146 B.n125 163.367
R268 B.n142 B.n125 163.367
R269 B.n142 B.n141 163.367
R270 B.n141 B.n140 163.367
R271 B.n140 B.n127 163.367
R272 B.n136 B.n127 163.367
R273 B.n136 B.n135 163.367
R274 B.n135 B.n134 163.367
R275 B.n134 B.n129 163.367
R276 B.n130 B.n129 163.367
R277 B.n130 B.n2 163.367
R278 B.n490 B.n2 163.367
R279 B.n490 B.n489 163.367
R280 B.n489 B.n488 163.367
R281 B.n488 B.n3 163.367
R282 B.n484 B.n3 163.367
R283 B.n484 B.n483 163.367
R284 B.n483 B.n482 163.367
R285 B.n482 B.n5 163.367
R286 B.n478 B.n5 163.367
R287 B.n478 B.n477 163.367
R288 B.n477 B.n476 163.367
R289 B.n476 B.n7 163.367
R290 B.n472 B.n7 163.367
R291 B.n472 B.n471 163.367
R292 B.n471 B.n470 163.367
R293 B.n470 B.n9 163.367
R294 B.n466 B.n9 163.367
R295 B.n466 B.n465 163.367
R296 B.n465 B.n464 163.367
R297 B.n464 B.n11 163.367
R298 B.n460 B.n11 163.367
R299 B.n460 B.n459 163.367
R300 B.n459 B.n458 163.367
R301 B.n458 B.n13 163.367
R302 B.n165 B.n164 163.367
R303 B.n166 B.n165 163.367
R304 B.n166 B.n117 163.367
R305 B.n170 B.n117 163.367
R306 B.n171 B.n170 163.367
R307 B.n172 B.n171 163.367
R308 B.n172 B.n115 163.367
R309 B.n176 B.n115 163.367
R310 B.n177 B.n176 163.367
R311 B.n178 B.n177 163.367
R312 B.n178 B.n113 163.367
R313 B.n182 B.n113 163.367
R314 B.n183 B.n182 163.367
R315 B.n184 B.n183 163.367
R316 B.n184 B.n111 163.367
R317 B.n188 B.n111 163.367
R318 B.n189 B.n188 163.367
R319 B.n190 B.n189 163.367
R320 B.n190 B.n109 163.367
R321 B.n194 B.n109 163.367
R322 B.n195 B.n194 163.367
R323 B.n196 B.n195 163.367
R324 B.n196 B.n107 163.367
R325 B.n200 B.n107 163.367
R326 B.n201 B.n200 163.367
R327 B.n202 B.n201 163.367
R328 B.n202 B.n105 163.367
R329 B.n206 B.n105 163.367
R330 B.n207 B.n206 163.367
R331 B.n208 B.n207 163.367
R332 B.n208 B.n101 163.367
R333 B.n213 B.n101 163.367
R334 B.n214 B.n213 163.367
R335 B.n215 B.n214 163.367
R336 B.n215 B.n99 163.367
R337 B.n219 B.n99 163.367
R338 B.n220 B.n219 163.367
R339 B.n221 B.n220 163.367
R340 B.n221 B.n97 163.367
R341 B.n225 B.n97 163.367
R342 B.n226 B.n225 163.367
R343 B.n226 B.n93 163.367
R344 B.n230 B.n93 163.367
R345 B.n231 B.n230 163.367
R346 B.n232 B.n231 163.367
R347 B.n232 B.n91 163.367
R348 B.n236 B.n91 163.367
R349 B.n237 B.n236 163.367
R350 B.n238 B.n237 163.367
R351 B.n238 B.n89 163.367
R352 B.n242 B.n89 163.367
R353 B.n243 B.n242 163.367
R354 B.n244 B.n243 163.367
R355 B.n244 B.n87 163.367
R356 B.n248 B.n87 163.367
R357 B.n249 B.n248 163.367
R358 B.n250 B.n249 163.367
R359 B.n250 B.n85 163.367
R360 B.n254 B.n85 163.367
R361 B.n255 B.n254 163.367
R362 B.n256 B.n255 163.367
R363 B.n256 B.n83 163.367
R364 B.n260 B.n83 163.367
R365 B.n261 B.n260 163.367
R366 B.n262 B.n261 163.367
R367 B.n262 B.n81 163.367
R368 B.n266 B.n81 163.367
R369 B.n267 B.n266 163.367
R370 B.n268 B.n267 163.367
R371 B.n268 B.n79 163.367
R372 B.n272 B.n79 163.367
R373 B.n273 B.n272 163.367
R374 B.n274 B.n77 163.367
R375 B.n278 B.n77 163.367
R376 B.n279 B.n278 163.367
R377 B.n280 B.n279 163.367
R378 B.n280 B.n75 163.367
R379 B.n284 B.n75 163.367
R380 B.n285 B.n284 163.367
R381 B.n286 B.n285 163.367
R382 B.n286 B.n73 163.367
R383 B.n290 B.n73 163.367
R384 B.n291 B.n290 163.367
R385 B.n292 B.n291 163.367
R386 B.n292 B.n71 163.367
R387 B.n296 B.n71 163.367
R388 B.n297 B.n296 163.367
R389 B.n298 B.n297 163.367
R390 B.n298 B.n69 163.367
R391 B.n302 B.n69 163.367
R392 B.n303 B.n302 163.367
R393 B.n304 B.n303 163.367
R394 B.n304 B.n67 163.367
R395 B.n308 B.n67 163.367
R396 B.n309 B.n308 163.367
R397 B.n310 B.n309 163.367
R398 B.n310 B.n65 163.367
R399 B.n314 B.n65 163.367
R400 B.n315 B.n314 163.367
R401 B.n316 B.n315 163.367
R402 B.n316 B.n63 163.367
R403 B.n320 B.n63 163.367
R404 B.n321 B.n320 163.367
R405 B.n322 B.n321 163.367
R406 B.n322 B.n61 163.367
R407 B.n326 B.n61 163.367
R408 B.n327 B.n326 163.367
R409 B.n328 B.n327 163.367
R410 B.n328 B.n59 163.367
R411 B.n332 B.n59 163.367
R412 B.n333 B.n332 163.367
R413 B.n334 B.n333 163.367
R414 B.n334 B.n57 163.367
R415 B.n338 B.n57 163.367
R416 B.n339 B.n338 163.367
R417 B.n340 B.n339 163.367
R418 B.n340 B.n55 163.367
R419 B.n344 B.n55 163.367
R420 B.n454 B.n453 163.367
R421 B.n453 B.n452 163.367
R422 B.n452 B.n15 163.367
R423 B.n448 B.n15 163.367
R424 B.n448 B.n447 163.367
R425 B.n447 B.n446 163.367
R426 B.n446 B.n17 163.367
R427 B.n442 B.n17 163.367
R428 B.n442 B.n441 163.367
R429 B.n441 B.n440 163.367
R430 B.n440 B.n19 163.367
R431 B.n436 B.n19 163.367
R432 B.n436 B.n435 163.367
R433 B.n435 B.n434 163.367
R434 B.n434 B.n21 163.367
R435 B.n430 B.n21 163.367
R436 B.n430 B.n429 163.367
R437 B.n429 B.n428 163.367
R438 B.n428 B.n23 163.367
R439 B.n424 B.n23 163.367
R440 B.n424 B.n423 163.367
R441 B.n423 B.n422 163.367
R442 B.n422 B.n25 163.367
R443 B.n418 B.n25 163.367
R444 B.n418 B.n417 163.367
R445 B.n417 B.n416 163.367
R446 B.n416 B.n27 163.367
R447 B.n412 B.n27 163.367
R448 B.n412 B.n411 163.367
R449 B.n411 B.n410 163.367
R450 B.n410 B.n29 163.367
R451 B.n405 B.n29 163.367
R452 B.n405 B.n404 163.367
R453 B.n404 B.n403 163.367
R454 B.n403 B.n33 163.367
R455 B.n399 B.n33 163.367
R456 B.n399 B.n398 163.367
R457 B.n398 B.n397 163.367
R458 B.n397 B.n35 163.367
R459 B.n393 B.n35 163.367
R460 B.n393 B.n392 163.367
R461 B.n392 B.n39 163.367
R462 B.n388 B.n39 163.367
R463 B.n388 B.n387 163.367
R464 B.n387 B.n386 163.367
R465 B.n386 B.n41 163.367
R466 B.n382 B.n41 163.367
R467 B.n382 B.n381 163.367
R468 B.n381 B.n380 163.367
R469 B.n380 B.n43 163.367
R470 B.n376 B.n43 163.367
R471 B.n376 B.n375 163.367
R472 B.n375 B.n374 163.367
R473 B.n374 B.n45 163.367
R474 B.n370 B.n45 163.367
R475 B.n370 B.n369 163.367
R476 B.n369 B.n368 163.367
R477 B.n368 B.n47 163.367
R478 B.n364 B.n47 163.367
R479 B.n364 B.n363 163.367
R480 B.n363 B.n362 163.367
R481 B.n362 B.n49 163.367
R482 B.n358 B.n49 163.367
R483 B.n358 B.n357 163.367
R484 B.n357 B.n356 163.367
R485 B.n356 B.n51 163.367
R486 B.n352 B.n51 163.367
R487 B.n352 B.n351 163.367
R488 B.n351 B.n350 163.367
R489 B.n350 B.n53 163.367
R490 B.n346 B.n53 163.367
R491 B.n346 B.n345 163.367
R492 B.n96 B.n95 59.5399
R493 B.n211 B.n103 59.5399
R494 B.n407 B.n31 59.5399
R495 B.n38 B.n37 59.5399
R496 B.n456 B.n455 32.3127
R497 B.n343 B.n54 32.3127
R498 B.n275 B.n78 32.3127
R499 B.n163 B.n162 32.3127
R500 B.n95 B.n94 24.4369
R501 B.n103 B.n102 24.4369
R502 B.n31 B.n30 24.4369
R503 B.n37 B.n36 24.4369
R504 B B.n491 18.0485
R505 B.n455 B.n14 10.6151
R506 B.n451 B.n14 10.6151
R507 B.n451 B.n450 10.6151
R508 B.n450 B.n449 10.6151
R509 B.n449 B.n16 10.6151
R510 B.n445 B.n16 10.6151
R511 B.n445 B.n444 10.6151
R512 B.n444 B.n443 10.6151
R513 B.n443 B.n18 10.6151
R514 B.n439 B.n18 10.6151
R515 B.n439 B.n438 10.6151
R516 B.n438 B.n437 10.6151
R517 B.n437 B.n20 10.6151
R518 B.n433 B.n20 10.6151
R519 B.n433 B.n432 10.6151
R520 B.n432 B.n431 10.6151
R521 B.n431 B.n22 10.6151
R522 B.n427 B.n22 10.6151
R523 B.n427 B.n426 10.6151
R524 B.n426 B.n425 10.6151
R525 B.n425 B.n24 10.6151
R526 B.n421 B.n24 10.6151
R527 B.n421 B.n420 10.6151
R528 B.n420 B.n419 10.6151
R529 B.n419 B.n26 10.6151
R530 B.n415 B.n26 10.6151
R531 B.n415 B.n414 10.6151
R532 B.n414 B.n413 10.6151
R533 B.n413 B.n28 10.6151
R534 B.n409 B.n28 10.6151
R535 B.n409 B.n408 10.6151
R536 B.n406 B.n32 10.6151
R537 B.n402 B.n32 10.6151
R538 B.n402 B.n401 10.6151
R539 B.n401 B.n400 10.6151
R540 B.n400 B.n34 10.6151
R541 B.n396 B.n34 10.6151
R542 B.n396 B.n395 10.6151
R543 B.n395 B.n394 10.6151
R544 B.n391 B.n390 10.6151
R545 B.n390 B.n389 10.6151
R546 B.n389 B.n40 10.6151
R547 B.n385 B.n40 10.6151
R548 B.n385 B.n384 10.6151
R549 B.n384 B.n383 10.6151
R550 B.n383 B.n42 10.6151
R551 B.n379 B.n42 10.6151
R552 B.n379 B.n378 10.6151
R553 B.n378 B.n377 10.6151
R554 B.n377 B.n44 10.6151
R555 B.n373 B.n44 10.6151
R556 B.n373 B.n372 10.6151
R557 B.n372 B.n371 10.6151
R558 B.n371 B.n46 10.6151
R559 B.n367 B.n46 10.6151
R560 B.n367 B.n366 10.6151
R561 B.n366 B.n365 10.6151
R562 B.n365 B.n48 10.6151
R563 B.n361 B.n48 10.6151
R564 B.n361 B.n360 10.6151
R565 B.n360 B.n359 10.6151
R566 B.n359 B.n50 10.6151
R567 B.n355 B.n50 10.6151
R568 B.n355 B.n354 10.6151
R569 B.n354 B.n353 10.6151
R570 B.n353 B.n52 10.6151
R571 B.n349 B.n52 10.6151
R572 B.n349 B.n348 10.6151
R573 B.n348 B.n347 10.6151
R574 B.n347 B.n54 10.6151
R575 B.n276 B.n275 10.6151
R576 B.n277 B.n276 10.6151
R577 B.n277 B.n76 10.6151
R578 B.n281 B.n76 10.6151
R579 B.n282 B.n281 10.6151
R580 B.n283 B.n282 10.6151
R581 B.n283 B.n74 10.6151
R582 B.n287 B.n74 10.6151
R583 B.n288 B.n287 10.6151
R584 B.n289 B.n288 10.6151
R585 B.n289 B.n72 10.6151
R586 B.n293 B.n72 10.6151
R587 B.n294 B.n293 10.6151
R588 B.n295 B.n294 10.6151
R589 B.n295 B.n70 10.6151
R590 B.n299 B.n70 10.6151
R591 B.n300 B.n299 10.6151
R592 B.n301 B.n300 10.6151
R593 B.n301 B.n68 10.6151
R594 B.n305 B.n68 10.6151
R595 B.n306 B.n305 10.6151
R596 B.n307 B.n306 10.6151
R597 B.n307 B.n66 10.6151
R598 B.n311 B.n66 10.6151
R599 B.n312 B.n311 10.6151
R600 B.n313 B.n312 10.6151
R601 B.n313 B.n64 10.6151
R602 B.n317 B.n64 10.6151
R603 B.n318 B.n317 10.6151
R604 B.n319 B.n318 10.6151
R605 B.n319 B.n62 10.6151
R606 B.n323 B.n62 10.6151
R607 B.n324 B.n323 10.6151
R608 B.n325 B.n324 10.6151
R609 B.n325 B.n60 10.6151
R610 B.n329 B.n60 10.6151
R611 B.n330 B.n329 10.6151
R612 B.n331 B.n330 10.6151
R613 B.n331 B.n58 10.6151
R614 B.n335 B.n58 10.6151
R615 B.n336 B.n335 10.6151
R616 B.n337 B.n336 10.6151
R617 B.n337 B.n56 10.6151
R618 B.n341 B.n56 10.6151
R619 B.n342 B.n341 10.6151
R620 B.n343 B.n342 10.6151
R621 B.n163 B.n118 10.6151
R622 B.n167 B.n118 10.6151
R623 B.n168 B.n167 10.6151
R624 B.n169 B.n168 10.6151
R625 B.n169 B.n116 10.6151
R626 B.n173 B.n116 10.6151
R627 B.n174 B.n173 10.6151
R628 B.n175 B.n174 10.6151
R629 B.n175 B.n114 10.6151
R630 B.n179 B.n114 10.6151
R631 B.n180 B.n179 10.6151
R632 B.n181 B.n180 10.6151
R633 B.n181 B.n112 10.6151
R634 B.n185 B.n112 10.6151
R635 B.n186 B.n185 10.6151
R636 B.n187 B.n186 10.6151
R637 B.n187 B.n110 10.6151
R638 B.n191 B.n110 10.6151
R639 B.n192 B.n191 10.6151
R640 B.n193 B.n192 10.6151
R641 B.n193 B.n108 10.6151
R642 B.n197 B.n108 10.6151
R643 B.n198 B.n197 10.6151
R644 B.n199 B.n198 10.6151
R645 B.n199 B.n106 10.6151
R646 B.n203 B.n106 10.6151
R647 B.n204 B.n203 10.6151
R648 B.n205 B.n204 10.6151
R649 B.n205 B.n104 10.6151
R650 B.n209 B.n104 10.6151
R651 B.n210 B.n209 10.6151
R652 B.n212 B.n100 10.6151
R653 B.n216 B.n100 10.6151
R654 B.n217 B.n216 10.6151
R655 B.n218 B.n217 10.6151
R656 B.n218 B.n98 10.6151
R657 B.n222 B.n98 10.6151
R658 B.n223 B.n222 10.6151
R659 B.n224 B.n223 10.6151
R660 B.n228 B.n227 10.6151
R661 B.n229 B.n228 10.6151
R662 B.n229 B.n92 10.6151
R663 B.n233 B.n92 10.6151
R664 B.n234 B.n233 10.6151
R665 B.n235 B.n234 10.6151
R666 B.n235 B.n90 10.6151
R667 B.n239 B.n90 10.6151
R668 B.n240 B.n239 10.6151
R669 B.n241 B.n240 10.6151
R670 B.n241 B.n88 10.6151
R671 B.n245 B.n88 10.6151
R672 B.n246 B.n245 10.6151
R673 B.n247 B.n246 10.6151
R674 B.n247 B.n86 10.6151
R675 B.n251 B.n86 10.6151
R676 B.n252 B.n251 10.6151
R677 B.n253 B.n252 10.6151
R678 B.n253 B.n84 10.6151
R679 B.n257 B.n84 10.6151
R680 B.n258 B.n257 10.6151
R681 B.n259 B.n258 10.6151
R682 B.n259 B.n82 10.6151
R683 B.n263 B.n82 10.6151
R684 B.n264 B.n263 10.6151
R685 B.n265 B.n264 10.6151
R686 B.n265 B.n80 10.6151
R687 B.n269 B.n80 10.6151
R688 B.n270 B.n269 10.6151
R689 B.n271 B.n270 10.6151
R690 B.n271 B.n78 10.6151
R691 B.n162 B.n161 10.6151
R692 B.n161 B.n120 10.6151
R693 B.n157 B.n120 10.6151
R694 B.n157 B.n156 10.6151
R695 B.n156 B.n155 10.6151
R696 B.n155 B.n122 10.6151
R697 B.n151 B.n122 10.6151
R698 B.n151 B.n150 10.6151
R699 B.n150 B.n149 10.6151
R700 B.n149 B.n124 10.6151
R701 B.n145 B.n124 10.6151
R702 B.n145 B.n144 10.6151
R703 B.n144 B.n143 10.6151
R704 B.n143 B.n126 10.6151
R705 B.n139 B.n126 10.6151
R706 B.n139 B.n138 10.6151
R707 B.n138 B.n137 10.6151
R708 B.n137 B.n128 10.6151
R709 B.n133 B.n128 10.6151
R710 B.n133 B.n132 10.6151
R711 B.n132 B.n131 10.6151
R712 B.n131 B.n0 10.6151
R713 B.n487 B.n1 10.6151
R714 B.n487 B.n486 10.6151
R715 B.n486 B.n485 10.6151
R716 B.n485 B.n4 10.6151
R717 B.n481 B.n4 10.6151
R718 B.n481 B.n480 10.6151
R719 B.n480 B.n479 10.6151
R720 B.n479 B.n6 10.6151
R721 B.n475 B.n6 10.6151
R722 B.n475 B.n474 10.6151
R723 B.n474 B.n473 10.6151
R724 B.n473 B.n8 10.6151
R725 B.n469 B.n8 10.6151
R726 B.n469 B.n468 10.6151
R727 B.n468 B.n467 10.6151
R728 B.n467 B.n10 10.6151
R729 B.n463 B.n10 10.6151
R730 B.n463 B.n462 10.6151
R731 B.n462 B.n461 10.6151
R732 B.n461 B.n12 10.6151
R733 B.n457 B.n12 10.6151
R734 B.n457 B.n456 10.6151
R735 B.n407 B.n406 6.5566
R736 B.n394 B.n38 6.5566
R737 B.n212 B.n211 6.5566
R738 B.n224 B.n96 6.5566
R739 B.n408 B.n407 4.05904
R740 B.n391 B.n38 4.05904
R741 B.n211 B.n210 4.05904
R742 B.n227 B.n96 4.05904
R743 B.n491 B.n0 2.81026
R744 B.n491 B.n1 2.81026
R745 VP.n5 VP.t1 284.711
R746 VP.n12 VP.t0 266.656
R747 VP.n19 VP.t3 266.656
R748 VP.n9 VP.t2 266.656
R749 VP.n1 VP.t4 224.156
R750 VP.n4 VP.t5 224.156
R751 VP.n20 VP.n19 161.3
R752 VP.n7 VP.n6 161.3
R753 VP.n8 VP.n3 161.3
R754 VP.n10 VP.n9 161.3
R755 VP.n18 VP.n0 161.3
R756 VP.n17 VP.n16 161.3
R757 VP.n15 VP.n14 161.3
R758 VP.n13 VP.n2 161.3
R759 VP.n12 VP.n11 161.3
R760 VP.n14 VP.n13 52.1486
R761 VP.n18 VP.n17 52.1486
R762 VP.n8 VP.n7 52.1486
R763 VP.n6 VP.n5 43.399
R764 VP.n5 VP.n4 42.4117
R765 VP.n11 VP.n10 39.6066
R766 VP.n14 VP.n1 12.234
R767 VP.n17 VP.n1 12.234
R768 VP.n7 VP.n4 12.234
R769 VP.n13 VP.n12 6.57323
R770 VP.n19 VP.n18 6.57323
R771 VP.n9 VP.n8 6.57323
R772 VP.n6 VP.n3 0.189894
R773 VP.n10 VP.n3 0.189894
R774 VP.n11 VP.n2 0.189894
R775 VP.n15 VP.n2 0.189894
R776 VP.n16 VP.n15 0.189894
R777 VP.n16 VP.n0 0.189894
R778 VP.n20 VP.n0 0.189894
R779 VP VP.n20 0.0516364
R780 VTAIL.n186 VTAIL.n146 756.745
R781 VTAIL.n42 VTAIL.n2 756.745
R782 VTAIL.n140 VTAIL.n100 756.745
R783 VTAIL.n92 VTAIL.n52 756.745
R784 VTAIL.n161 VTAIL.n160 585
R785 VTAIL.n158 VTAIL.n157 585
R786 VTAIL.n167 VTAIL.n166 585
R787 VTAIL.n169 VTAIL.n168 585
R788 VTAIL.n154 VTAIL.n153 585
R789 VTAIL.n175 VTAIL.n174 585
R790 VTAIL.n178 VTAIL.n177 585
R791 VTAIL.n176 VTAIL.n150 585
R792 VTAIL.n183 VTAIL.n149 585
R793 VTAIL.n185 VTAIL.n184 585
R794 VTAIL.n187 VTAIL.n186 585
R795 VTAIL.n17 VTAIL.n16 585
R796 VTAIL.n14 VTAIL.n13 585
R797 VTAIL.n23 VTAIL.n22 585
R798 VTAIL.n25 VTAIL.n24 585
R799 VTAIL.n10 VTAIL.n9 585
R800 VTAIL.n31 VTAIL.n30 585
R801 VTAIL.n34 VTAIL.n33 585
R802 VTAIL.n32 VTAIL.n6 585
R803 VTAIL.n39 VTAIL.n5 585
R804 VTAIL.n41 VTAIL.n40 585
R805 VTAIL.n43 VTAIL.n42 585
R806 VTAIL.n141 VTAIL.n140 585
R807 VTAIL.n139 VTAIL.n138 585
R808 VTAIL.n137 VTAIL.n103 585
R809 VTAIL.n107 VTAIL.n104 585
R810 VTAIL.n132 VTAIL.n131 585
R811 VTAIL.n130 VTAIL.n129 585
R812 VTAIL.n109 VTAIL.n108 585
R813 VTAIL.n124 VTAIL.n123 585
R814 VTAIL.n122 VTAIL.n121 585
R815 VTAIL.n113 VTAIL.n112 585
R816 VTAIL.n116 VTAIL.n115 585
R817 VTAIL.n93 VTAIL.n92 585
R818 VTAIL.n91 VTAIL.n90 585
R819 VTAIL.n89 VTAIL.n55 585
R820 VTAIL.n59 VTAIL.n56 585
R821 VTAIL.n84 VTAIL.n83 585
R822 VTAIL.n82 VTAIL.n81 585
R823 VTAIL.n61 VTAIL.n60 585
R824 VTAIL.n76 VTAIL.n75 585
R825 VTAIL.n74 VTAIL.n73 585
R826 VTAIL.n65 VTAIL.n64 585
R827 VTAIL.n68 VTAIL.n67 585
R828 VTAIL.t8 VTAIL.n114 329.039
R829 VTAIL.t5 VTAIL.n66 329.039
R830 VTAIL.t1 VTAIL.n159 329.038
R831 VTAIL.t7 VTAIL.n15 329.038
R832 VTAIL.n160 VTAIL.n157 171.744
R833 VTAIL.n167 VTAIL.n157 171.744
R834 VTAIL.n168 VTAIL.n167 171.744
R835 VTAIL.n168 VTAIL.n153 171.744
R836 VTAIL.n175 VTAIL.n153 171.744
R837 VTAIL.n177 VTAIL.n175 171.744
R838 VTAIL.n177 VTAIL.n176 171.744
R839 VTAIL.n176 VTAIL.n149 171.744
R840 VTAIL.n185 VTAIL.n149 171.744
R841 VTAIL.n186 VTAIL.n185 171.744
R842 VTAIL.n16 VTAIL.n13 171.744
R843 VTAIL.n23 VTAIL.n13 171.744
R844 VTAIL.n24 VTAIL.n23 171.744
R845 VTAIL.n24 VTAIL.n9 171.744
R846 VTAIL.n31 VTAIL.n9 171.744
R847 VTAIL.n33 VTAIL.n31 171.744
R848 VTAIL.n33 VTAIL.n32 171.744
R849 VTAIL.n32 VTAIL.n5 171.744
R850 VTAIL.n41 VTAIL.n5 171.744
R851 VTAIL.n42 VTAIL.n41 171.744
R852 VTAIL.n140 VTAIL.n139 171.744
R853 VTAIL.n139 VTAIL.n103 171.744
R854 VTAIL.n107 VTAIL.n103 171.744
R855 VTAIL.n131 VTAIL.n107 171.744
R856 VTAIL.n131 VTAIL.n130 171.744
R857 VTAIL.n130 VTAIL.n108 171.744
R858 VTAIL.n123 VTAIL.n108 171.744
R859 VTAIL.n123 VTAIL.n122 171.744
R860 VTAIL.n122 VTAIL.n112 171.744
R861 VTAIL.n115 VTAIL.n112 171.744
R862 VTAIL.n92 VTAIL.n91 171.744
R863 VTAIL.n91 VTAIL.n55 171.744
R864 VTAIL.n59 VTAIL.n55 171.744
R865 VTAIL.n83 VTAIL.n59 171.744
R866 VTAIL.n83 VTAIL.n82 171.744
R867 VTAIL.n82 VTAIL.n60 171.744
R868 VTAIL.n75 VTAIL.n60 171.744
R869 VTAIL.n75 VTAIL.n74 171.744
R870 VTAIL.n74 VTAIL.n64 171.744
R871 VTAIL.n67 VTAIL.n64 171.744
R872 VTAIL.n160 VTAIL.t1 85.8723
R873 VTAIL.n16 VTAIL.t7 85.8723
R874 VTAIL.n115 VTAIL.t8 85.8723
R875 VTAIL.n67 VTAIL.t5 85.8723
R876 VTAIL.n99 VTAIL.n98 66.1467
R877 VTAIL.n51 VTAIL.n50 66.1467
R878 VTAIL.n1 VTAIL.n0 66.1465
R879 VTAIL.n49 VTAIL.n48 66.1465
R880 VTAIL.n191 VTAIL.n190 34.7066
R881 VTAIL.n47 VTAIL.n46 34.7066
R882 VTAIL.n145 VTAIL.n144 34.7066
R883 VTAIL.n97 VTAIL.n96 34.7066
R884 VTAIL.n51 VTAIL.n49 21.9962
R885 VTAIL.n191 VTAIL.n145 20.91
R886 VTAIL.n184 VTAIL.n183 13.1884
R887 VTAIL.n40 VTAIL.n39 13.1884
R888 VTAIL.n138 VTAIL.n137 13.1884
R889 VTAIL.n90 VTAIL.n89 13.1884
R890 VTAIL.n182 VTAIL.n150 12.8005
R891 VTAIL.n187 VTAIL.n148 12.8005
R892 VTAIL.n38 VTAIL.n6 12.8005
R893 VTAIL.n43 VTAIL.n4 12.8005
R894 VTAIL.n141 VTAIL.n102 12.8005
R895 VTAIL.n136 VTAIL.n104 12.8005
R896 VTAIL.n93 VTAIL.n54 12.8005
R897 VTAIL.n88 VTAIL.n56 12.8005
R898 VTAIL.n179 VTAIL.n178 12.0247
R899 VTAIL.n188 VTAIL.n146 12.0247
R900 VTAIL.n35 VTAIL.n34 12.0247
R901 VTAIL.n44 VTAIL.n2 12.0247
R902 VTAIL.n142 VTAIL.n100 12.0247
R903 VTAIL.n133 VTAIL.n132 12.0247
R904 VTAIL.n94 VTAIL.n52 12.0247
R905 VTAIL.n85 VTAIL.n84 12.0247
R906 VTAIL.n174 VTAIL.n152 11.249
R907 VTAIL.n30 VTAIL.n8 11.249
R908 VTAIL.n129 VTAIL.n106 11.249
R909 VTAIL.n81 VTAIL.n58 11.249
R910 VTAIL.n161 VTAIL.n159 10.7239
R911 VTAIL.n17 VTAIL.n15 10.7239
R912 VTAIL.n116 VTAIL.n114 10.7239
R913 VTAIL.n68 VTAIL.n66 10.7239
R914 VTAIL.n173 VTAIL.n154 10.4732
R915 VTAIL.n29 VTAIL.n10 10.4732
R916 VTAIL.n128 VTAIL.n109 10.4732
R917 VTAIL.n80 VTAIL.n61 10.4732
R918 VTAIL.n170 VTAIL.n169 9.69747
R919 VTAIL.n26 VTAIL.n25 9.69747
R920 VTAIL.n125 VTAIL.n124 9.69747
R921 VTAIL.n77 VTAIL.n76 9.69747
R922 VTAIL.n190 VTAIL.n189 9.45567
R923 VTAIL.n46 VTAIL.n45 9.45567
R924 VTAIL.n144 VTAIL.n143 9.45567
R925 VTAIL.n96 VTAIL.n95 9.45567
R926 VTAIL.n189 VTAIL.n188 9.3005
R927 VTAIL.n148 VTAIL.n147 9.3005
R928 VTAIL.n163 VTAIL.n162 9.3005
R929 VTAIL.n165 VTAIL.n164 9.3005
R930 VTAIL.n156 VTAIL.n155 9.3005
R931 VTAIL.n171 VTAIL.n170 9.3005
R932 VTAIL.n173 VTAIL.n172 9.3005
R933 VTAIL.n152 VTAIL.n151 9.3005
R934 VTAIL.n180 VTAIL.n179 9.3005
R935 VTAIL.n182 VTAIL.n181 9.3005
R936 VTAIL.n45 VTAIL.n44 9.3005
R937 VTAIL.n4 VTAIL.n3 9.3005
R938 VTAIL.n19 VTAIL.n18 9.3005
R939 VTAIL.n21 VTAIL.n20 9.3005
R940 VTAIL.n12 VTAIL.n11 9.3005
R941 VTAIL.n27 VTAIL.n26 9.3005
R942 VTAIL.n29 VTAIL.n28 9.3005
R943 VTAIL.n8 VTAIL.n7 9.3005
R944 VTAIL.n36 VTAIL.n35 9.3005
R945 VTAIL.n38 VTAIL.n37 9.3005
R946 VTAIL.n118 VTAIL.n117 9.3005
R947 VTAIL.n120 VTAIL.n119 9.3005
R948 VTAIL.n111 VTAIL.n110 9.3005
R949 VTAIL.n126 VTAIL.n125 9.3005
R950 VTAIL.n128 VTAIL.n127 9.3005
R951 VTAIL.n106 VTAIL.n105 9.3005
R952 VTAIL.n134 VTAIL.n133 9.3005
R953 VTAIL.n136 VTAIL.n135 9.3005
R954 VTAIL.n143 VTAIL.n142 9.3005
R955 VTAIL.n102 VTAIL.n101 9.3005
R956 VTAIL.n70 VTAIL.n69 9.3005
R957 VTAIL.n72 VTAIL.n71 9.3005
R958 VTAIL.n63 VTAIL.n62 9.3005
R959 VTAIL.n78 VTAIL.n77 9.3005
R960 VTAIL.n80 VTAIL.n79 9.3005
R961 VTAIL.n58 VTAIL.n57 9.3005
R962 VTAIL.n86 VTAIL.n85 9.3005
R963 VTAIL.n88 VTAIL.n87 9.3005
R964 VTAIL.n95 VTAIL.n94 9.3005
R965 VTAIL.n54 VTAIL.n53 9.3005
R966 VTAIL.n166 VTAIL.n156 8.92171
R967 VTAIL.n22 VTAIL.n12 8.92171
R968 VTAIL.n121 VTAIL.n111 8.92171
R969 VTAIL.n73 VTAIL.n63 8.92171
R970 VTAIL.n165 VTAIL.n158 8.14595
R971 VTAIL.n21 VTAIL.n14 8.14595
R972 VTAIL.n120 VTAIL.n113 8.14595
R973 VTAIL.n72 VTAIL.n65 8.14595
R974 VTAIL.n162 VTAIL.n161 7.3702
R975 VTAIL.n18 VTAIL.n17 7.3702
R976 VTAIL.n117 VTAIL.n116 7.3702
R977 VTAIL.n69 VTAIL.n68 7.3702
R978 VTAIL.n162 VTAIL.n158 5.81868
R979 VTAIL.n18 VTAIL.n14 5.81868
R980 VTAIL.n117 VTAIL.n113 5.81868
R981 VTAIL.n69 VTAIL.n65 5.81868
R982 VTAIL.n166 VTAIL.n165 5.04292
R983 VTAIL.n22 VTAIL.n21 5.04292
R984 VTAIL.n121 VTAIL.n120 5.04292
R985 VTAIL.n73 VTAIL.n72 5.04292
R986 VTAIL.n169 VTAIL.n156 4.26717
R987 VTAIL.n25 VTAIL.n12 4.26717
R988 VTAIL.n124 VTAIL.n111 4.26717
R989 VTAIL.n76 VTAIL.n63 4.26717
R990 VTAIL.n0 VTAIL.t0 3.7583
R991 VTAIL.n0 VTAIL.t4 3.7583
R992 VTAIL.n48 VTAIL.t9 3.7583
R993 VTAIL.n48 VTAIL.t11 3.7583
R994 VTAIL.n98 VTAIL.t6 3.7583
R995 VTAIL.n98 VTAIL.t10 3.7583
R996 VTAIL.n50 VTAIL.t2 3.7583
R997 VTAIL.n50 VTAIL.t3 3.7583
R998 VTAIL.n170 VTAIL.n154 3.49141
R999 VTAIL.n26 VTAIL.n10 3.49141
R1000 VTAIL.n125 VTAIL.n109 3.49141
R1001 VTAIL.n77 VTAIL.n61 3.49141
R1002 VTAIL.n174 VTAIL.n173 2.71565
R1003 VTAIL.n30 VTAIL.n29 2.71565
R1004 VTAIL.n129 VTAIL.n128 2.71565
R1005 VTAIL.n81 VTAIL.n80 2.71565
R1006 VTAIL.n163 VTAIL.n159 2.41285
R1007 VTAIL.n19 VTAIL.n15 2.41285
R1008 VTAIL.n118 VTAIL.n114 2.41285
R1009 VTAIL.n70 VTAIL.n66 2.41285
R1010 VTAIL.n178 VTAIL.n152 1.93989
R1011 VTAIL.n190 VTAIL.n146 1.93989
R1012 VTAIL.n34 VTAIL.n8 1.93989
R1013 VTAIL.n46 VTAIL.n2 1.93989
R1014 VTAIL.n144 VTAIL.n100 1.93989
R1015 VTAIL.n132 VTAIL.n106 1.93989
R1016 VTAIL.n96 VTAIL.n52 1.93989
R1017 VTAIL.n84 VTAIL.n58 1.93989
R1018 VTAIL.n179 VTAIL.n150 1.16414
R1019 VTAIL.n188 VTAIL.n187 1.16414
R1020 VTAIL.n35 VTAIL.n6 1.16414
R1021 VTAIL.n44 VTAIL.n43 1.16414
R1022 VTAIL.n142 VTAIL.n141 1.16414
R1023 VTAIL.n133 VTAIL.n104 1.16414
R1024 VTAIL.n94 VTAIL.n93 1.16414
R1025 VTAIL.n85 VTAIL.n56 1.16414
R1026 VTAIL.n97 VTAIL.n51 1.08671
R1027 VTAIL.n145 VTAIL.n99 1.08671
R1028 VTAIL.n49 VTAIL.n47 1.08671
R1029 VTAIL.n99 VTAIL.n97 1.01343
R1030 VTAIL.n47 VTAIL.n1 1.01343
R1031 VTAIL VTAIL.n191 0.756965
R1032 VTAIL.n183 VTAIL.n182 0.388379
R1033 VTAIL.n184 VTAIL.n148 0.388379
R1034 VTAIL.n39 VTAIL.n38 0.388379
R1035 VTAIL.n40 VTAIL.n4 0.388379
R1036 VTAIL.n138 VTAIL.n102 0.388379
R1037 VTAIL.n137 VTAIL.n136 0.388379
R1038 VTAIL.n90 VTAIL.n54 0.388379
R1039 VTAIL.n89 VTAIL.n88 0.388379
R1040 VTAIL VTAIL.n1 0.330241
R1041 VTAIL.n164 VTAIL.n163 0.155672
R1042 VTAIL.n164 VTAIL.n155 0.155672
R1043 VTAIL.n171 VTAIL.n155 0.155672
R1044 VTAIL.n172 VTAIL.n171 0.155672
R1045 VTAIL.n172 VTAIL.n151 0.155672
R1046 VTAIL.n180 VTAIL.n151 0.155672
R1047 VTAIL.n181 VTAIL.n180 0.155672
R1048 VTAIL.n181 VTAIL.n147 0.155672
R1049 VTAIL.n189 VTAIL.n147 0.155672
R1050 VTAIL.n20 VTAIL.n19 0.155672
R1051 VTAIL.n20 VTAIL.n11 0.155672
R1052 VTAIL.n27 VTAIL.n11 0.155672
R1053 VTAIL.n28 VTAIL.n27 0.155672
R1054 VTAIL.n28 VTAIL.n7 0.155672
R1055 VTAIL.n36 VTAIL.n7 0.155672
R1056 VTAIL.n37 VTAIL.n36 0.155672
R1057 VTAIL.n37 VTAIL.n3 0.155672
R1058 VTAIL.n45 VTAIL.n3 0.155672
R1059 VTAIL.n143 VTAIL.n101 0.155672
R1060 VTAIL.n135 VTAIL.n101 0.155672
R1061 VTAIL.n135 VTAIL.n134 0.155672
R1062 VTAIL.n134 VTAIL.n105 0.155672
R1063 VTAIL.n127 VTAIL.n105 0.155672
R1064 VTAIL.n127 VTAIL.n126 0.155672
R1065 VTAIL.n126 VTAIL.n110 0.155672
R1066 VTAIL.n119 VTAIL.n110 0.155672
R1067 VTAIL.n119 VTAIL.n118 0.155672
R1068 VTAIL.n95 VTAIL.n53 0.155672
R1069 VTAIL.n87 VTAIL.n53 0.155672
R1070 VTAIL.n87 VTAIL.n86 0.155672
R1071 VTAIL.n86 VTAIL.n57 0.155672
R1072 VTAIL.n79 VTAIL.n57 0.155672
R1073 VTAIL.n79 VTAIL.n78 0.155672
R1074 VTAIL.n78 VTAIL.n62 0.155672
R1075 VTAIL.n71 VTAIL.n62 0.155672
R1076 VTAIL.n71 VTAIL.n70 0.155672
R1077 VDD1.n40 VDD1.n0 756.745
R1078 VDD1.n85 VDD1.n45 756.745
R1079 VDD1.n41 VDD1.n40 585
R1080 VDD1.n39 VDD1.n38 585
R1081 VDD1.n37 VDD1.n3 585
R1082 VDD1.n7 VDD1.n4 585
R1083 VDD1.n32 VDD1.n31 585
R1084 VDD1.n30 VDD1.n29 585
R1085 VDD1.n9 VDD1.n8 585
R1086 VDD1.n24 VDD1.n23 585
R1087 VDD1.n22 VDD1.n21 585
R1088 VDD1.n13 VDD1.n12 585
R1089 VDD1.n16 VDD1.n15 585
R1090 VDD1.n60 VDD1.n59 585
R1091 VDD1.n57 VDD1.n56 585
R1092 VDD1.n66 VDD1.n65 585
R1093 VDD1.n68 VDD1.n67 585
R1094 VDD1.n53 VDD1.n52 585
R1095 VDD1.n74 VDD1.n73 585
R1096 VDD1.n77 VDD1.n76 585
R1097 VDD1.n75 VDD1.n49 585
R1098 VDD1.n82 VDD1.n48 585
R1099 VDD1.n84 VDD1.n83 585
R1100 VDD1.n86 VDD1.n85 585
R1101 VDD1.t4 VDD1.n14 329.039
R1102 VDD1.t5 VDD1.n58 329.038
R1103 VDD1.n40 VDD1.n39 171.744
R1104 VDD1.n39 VDD1.n3 171.744
R1105 VDD1.n7 VDD1.n3 171.744
R1106 VDD1.n31 VDD1.n7 171.744
R1107 VDD1.n31 VDD1.n30 171.744
R1108 VDD1.n30 VDD1.n8 171.744
R1109 VDD1.n23 VDD1.n8 171.744
R1110 VDD1.n23 VDD1.n22 171.744
R1111 VDD1.n22 VDD1.n12 171.744
R1112 VDD1.n15 VDD1.n12 171.744
R1113 VDD1.n59 VDD1.n56 171.744
R1114 VDD1.n66 VDD1.n56 171.744
R1115 VDD1.n67 VDD1.n66 171.744
R1116 VDD1.n67 VDD1.n52 171.744
R1117 VDD1.n74 VDD1.n52 171.744
R1118 VDD1.n76 VDD1.n74 171.744
R1119 VDD1.n76 VDD1.n75 171.744
R1120 VDD1.n75 VDD1.n48 171.744
R1121 VDD1.n84 VDD1.n48 171.744
R1122 VDD1.n85 VDD1.n84 171.744
R1123 VDD1.n15 VDD1.t4 85.8723
R1124 VDD1.n59 VDD1.t5 85.8723
R1125 VDD1.n91 VDD1.n90 83.0415
R1126 VDD1.n93 VDD1.n92 82.8253
R1127 VDD1 VDD1.n44 52.2582
R1128 VDD1.n91 VDD1.n89 52.1447
R1129 VDD1.n93 VDD1.n91 35.8285
R1130 VDD1.n38 VDD1.n37 13.1884
R1131 VDD1.n83 VDD1.n82 13.1884
R1132 VDD1.n41 VDD1.n2 12.8005
R1133 VDD1.n36 VDD1.n4 12.8005
R1134 VDD1.n81 VDD1.n49 12.8005
R1135 VDD1.n86 VDD1.n47 12.8005
R1136 VDD1.n42 VDD1.n0 12.0247
R1137 VDD1.n33 VDD1.n32 12.0247
R1138 VDD1.n78 VDD1.n77 12.0247
R1139 VDD1.n87 VDD1.n45 12.0247
R1140 VDD1.n29 VDD1.n6 11.249
R1141 VDD1.n73 VDD1.n51 11.249
R1142 VDD1.n16 VDD1.n14 10.7239
R1143 VDD1.n60 VDD1.n58 10.7239
R1144 VDD1.n28 VDD1.n9 10.4732
R1145 VDD1.n72 VDD1.n53 10.4732
R1146 VDD1.n25 VDD1.n24 9.69747
R1147 VDD1.n69 VDD1.n68 9.69747
R1148 VDD1.n44 VDD1.n43 9.45567
R1149 VDD1.n89 VDD1.n88 9.45567
R1150 VDD1.n18 VDD1.n17 9.3005
R1151 VDD1.n20 VDD1.n19 9.3005
R1152 VDD1.n11 VDD1.n10 9.3005
R1153 VDD1.n26 VDD1.n25 9.3005
R1154 VDD1.n28 VDD1.n27 9.3005
R1155 VDD1.n6 VDD1.n5 9.3005
R1156 VDD1.n34 VDD1.n33 9.3005
R1157 VDD1.n36 VDD1.n35 9.3005
R1158 VDD1.n43 VDD1.n42 9.3005
R1159 VDD1.n2 VDD1.n1 9.3005
R1160 VDD1.n88 VDD1.n87 9.3005
R1161 VDD1.n47 VDD1.n46 9.3005
R1162 VDD1.n62 VDD1.n61 9.3005
R1163 VDD1.n64 VDD1.n63 9.3005
R1164 VDD1.n55 VDD1.n54 9.3005
R1165 VDD1.n70 VDD1.n69 9.3005
R1166 VDD1.n72 VDD1.n71 9.3005
R1167 VDD1.n51 VDD1.n50 9.3005
R1168 VDD1.n79 VDD1.n78 9.3005
R1169 VDD1.n81 VDD1.n80 9.3005
R1170 VDD1.n21 VDD1.n11 8.92171
R1171 VDD1.n65 VDD1.n55 8.92171
R1172 VDD1.n20 VDD1.n13 8.14595
R1173 VDD1.n64 VDD1.n57 8.14595
R1174 VDD1.n17 VDD1.n16 7.3702
R1175 VDD1.n61 VDD1.n60 7.3702
R1176 VDD1.n17 VDD1.n13 5.81868
R1177 VDD1.n61 VDD1.n57 5.81868
R1178 VDD1.n21 VDD1.n20 5.04292
R1179 VDD1.n65 VDD1.n64 5.04292
R1180 VDD1.n24 VDD1.n11 4.26717
R1181 VDD1.n68 VDD1.n55 4.26717
R1182 VDD1.n92 VDD1.t0 3.7583
R1183 VDD1.n92 VDD1.t3 3.7583
R1184 VDD1.n90 VDD1.t1 3.7583
R1185 VDD1.n90 VDD1.t2 3.7583
R1186 VDD1.n25 VDD1.n9 3.49141
R1187 VDD1.n69 VDD1.n53 3.49141
R1188 VDD1.n29 VDD1.n28 2.71565
R1189 VDD1.n73 VDD1.n72 2.71565
R1190 VDD1.n18 VDD1.n14 2.41285
R1191 VDD1.n62 VDD1.n58 2.41285
R1192 VDD1.n44 VDD1.n0 1.93989
R1193 VDD1.n32 VDD1.n6 1.93989
R1194 VDD1.n77 VDD1.n51 1.93989
R1195 VDD1.n89 VDD1.n45 1.93989
R1196 VDD1.n42 VDD1.n41 1.16414
R1197 VDD1.n33 VDD1.n4 1.16414
R1198 VDD1.n78 VDD1.n49 1.16414
R1199 VDD1.n87 VDD1.n86 1.16414
R1200 VDD1.n38 VDD1.n2 0.388379
R1201 VDD1.n37 VDD1.n36 0.388379
R1202 VDD1.n82 VDD1.n81 0.388379
R1203 VDD1.n83 VDD1.n47 0.388379
R1204 VDD1 VDD1.n93 0.213862
R1205 VDD1.n43 VDD1.n1 0.155672
R1206 VDD1.n35 VDD1.n1 0.155672
R1207 VDD1.n35 VDD1.n34 0.155672
R1208 VDD1.n34 VDD1.n5 0.155672
R1209 VDD1.n27 VDD1.n5 0.155672
R1210 VDD1.n27 VDD1.n26 0.155672
R1211 VDD1.n26 VDD1.n10 0.155672
R1212 VDD1.n19 VDD1.n10 0.155672
R1213 VDD1.n19 VDD1.n18 0.155672
R1214 VDD1.n63 VDD1.n62 0.155672
R1215 VDD1.n63 VDD1.n54 0.155672
R1216 VDD1.n70 VDD1.n54 0.155672
R1217 VDD1.n71 VDD1.n70 0.155672
R1218 VDD1.n71 VDD1.n50 0.155672
R1219 VDD1.n79 VDD1.n50 0.155672
R1220 VDD1.n80 VDD1.n79 0.155672
R1221 VDD1.n80 VDD1.n46 0.155672
R1222 VDD1.n88 VDD1.n46 0.155672
R1223 VN.n2 VN.t2 284.711
R1224 VN.n10 VN.t0 284.711
R1225 VN.n6 VN.t3 266.656
R1226 VN.n14 VN.t4 266.656
R1227 VN.n1 VN.t1 224.156
R1228 VN.n9 VN.t5 224.156
R1229 VN.n7 VN.n6 161.3
R1230 VN.n15 VN.n14 161.3
R1231 VN.n13 VN.n8 161.3
R1232 VN.n12 VN.n11 161.3
R1233 VN.n5 VN.n0 161.3
R1234 VN.n4 VN.n3 161.3
R1235 VN.n5 VN.n4 52.1486
R1236 VN.n13 VN.n12 52.1486
R1237 VN.n11 VN.n10 43.399
R1238 VN.n3 VN.n2 43.399
R1239 VN.n2 VN.n1 42.4117
R1240 VN.n10 VN.n9 42.4117
R1241 VN VN.n15 39.9872
R1242 VN.n4 VN.n1 12.234
R1243 VN.n12 VN.n9 12.234
R1244 VN.n6 VN.n5 6.57323
R1245 VN.n14 VN.n13 6.57323
R1246 VN.n15 VN.n8 0.189894
R1247 VN.n11 VN.n8 0.189894
R1248 VN.n3 VN.n0 0.189894
R1249 VN.n7 VN.n0 0.189894
R1250 VN VN.n7 0.0516364
R1251 VDD2.n87 VDD2.n47 756.745
R1252 VDD2.n40 VDD2.n0 756.745
R1253 VDD2.n88 VDD2.n87 585
R1254 VDD2.n86 VDD2.n85 585
R1255 VDD2.n84 VDD2.n50 585
R1256 VDD2.n54 VDD2.n51 585
R1257 VDD2.n79 VDD2.n78 585
R1258 VDD2.n77 VDD2.n76 585
R1259 VDD2.n56 VDD2.n55 585
R1260 VDD2.n71 VDD2.n70 585
R1261 VDD2.n69 VDD2.n68 585
R1262 VDD2.n60 VDD2.n59 585
R1263 VDD2.n63 VDD2.n62 585
R1264 VDD2.n15 VDD2.n14 585
R1265 VDD2.n12 VDD2.n11 585
R1266 VDD2.n21 VDD2.n20 585
R1267 VDD2.n23 VDD2.n22 585
R1268 VDD2.n8 VDD2.n7 585
R1269 VDD2.n29 VDD2.n28 585
R1270 VDD2.n32 VDD2.n31 585
R1271 VDD2.n30 VDD2.n4 585
R1272 VDD2.n37 VDD2.n3 585
R1273 VDD2.n39 VDD2.n38 585
R1274 VDD2.n41 VDD2.n40 585
R1275 VDD2.t1 VDD2.n61 329.039
R1276 VDD2.t3 VDD2.n13 329.038
R1277 VDD2.n87 VDD2.n86 171.744
R1278 VDD2.n86 VDD2.n50 171.744
R1279 VDD2.n54 VDD2.n50 171.744
R1280 VDD2.n78 VDD2.n54 171.744
R1281 VDD2.n78 VDD2.n77 171.744
R1282 VDD2.n77 VDD2.n55 171.744
R1283 VDD2.n70 VDD2.n55 171.744
R1284 VDD2.n70 VDD2.n69 171.744
R1285 VDD2.n69 VDD2.n59 171.744
R1286 VDD2.n62 VDD2.n59 171.744
R1287 VDD2.n14 VDD2.n11 171.744
R1288 VDD2.n21 VDD2.n11 171.744
R1289 VDD2.n22 VDD2.n21 171.744
R1290 VDD2.n22 VDD2.n7 171.744
R1291 VDD2.n29 VDD2.n7 171.744
R1292 VDD2.n31 VDD2.n29 171.744
R1293 VDD2.n31 VDD2.n30 171.744
R1294 VDD2.n30 VDD2.n3 171.744
R1295 VDD2.n39 VDD2.n3 171.744
R1296 VDD2.n40 VDD2.n39 171.744
R1297 VDD2.n62 VDD2.t1 85.8723
R1298 VDD2.n14 VDD2.t3 85.8723
R1299 VDD2.n46 VDD2.n45 83.0415
R1300 VDD2 VDD2.n93 83.0387
R1301 VDD2.n46 VDD2.n44 52.1447
R1302 VDD2.n92 VDD2.n91 51.3853
R1303 VDD2.n92 VDD2.n46 34.7024
R1304 VDD2.n85 VDD2.n84 13.1884
R1305 VDD2.n38 VDD2.n37 13.1884
R1306 VDD2.n88 VDD2.n49 12.8005
R1307 VDD2.n83 VDD2.n51 12.8005
R1308 VDD2.n36 VDD2.n4 12.8005
R1309 VDD2.n41 VDD2.n2 12.8005
R1310 VDD2.n89 VDD2.n47 12.0247
R1311 VDD2.n80 VDD2.n79 12.0247
R1312 VDD2.n33 VDD2.n32 12.0247
R1313 VDD2.n42 VDD2.n0 12.0247
R1314 VDD2.n76 VDD2.n53 11.249
R1315 VDD2.n28 VDD2.n6 11.249
R1316 VDD2.n63 VDD2.n61 10.7239
R1317 VDD2.n15 VDD2.n13 10.7239
R1318 VDD2.n75 VDD2.n56 10.4732
R1319 VDD2.n27 VDD2.n8 10.4732
R1320 VDD2.n72 VDD2.n71 9.69747
R1321 VDD2.n24 VDD2.n23 9.69747
R1322 VDD2.n91 VDD2.n90 9.45567
R1323 VDD2.n44 VDD2.n43 9.45567
R1324 VDD2.n65 VDD2.n64 9.3005
R1325 VDD2.n67 VDD2.n66 9.3005
R1326 VDD2.n58 VDD2.n57 9.3005
R1327 VDD2.n73 VDD2.n72 9.3005
R1328 VDD2.n75 VDD2.n74 9.3005
R1329 VDD2.n53 VDD2.n52 9.3005
R1330 VDD2.n81 VDD2.n80 9.3005
R1331 VDD2.n83 VDD2.n82 9.3005
R1332 VDD2.n90 VDD2.n89 9.3005
R1333 VDD2.n49 VDD2.n48 9.3005
R1334 VDD2.n43 VDD2.n42 9.3005
R1335 VDD2.n2 VDD2.n1 9.3005
R1336 VDD2.n17 VDD2.n16 9.3005
R1337 VDD2.n19 VDD2.n18 9.3005
R1338 VDD2.n10 VDD2.n9 9.3005
R1339 VDD2.n25 VDD2.n24 9.3005
R1340 VDD2.n27 VDD2.n26 9.3005
R1341 VDD2.n6 VDD2.n5 9.3005
R1342 VDD2.n34 VDD2.n33 9.3005
R1343 VDD2.n36 VDD2.n35 9.3005
R1344 VDD2.n68 VDD2.n58 8.92171
R1345 VDD2.n20 VDD2.n10 8.92171
R1346 VDD2.n67 VDD2.n60 8.14595
R1347 VDD2.n19 VDD2.n12 8.14595
R1348 VDD2.n64 VDD2.n63 7.3702
R1349 VDD2.n16 VDD2.n15 7.3702
R1350 VDD2.n64 VDD2.n60 5.81868
R1351 VDD2.n16 VDD2.n12 5.81868
R1352 VDD2.n68 VDD2.n67 5.04292
R1353 VDD2.n20 VDD2.n19 5.04292
R1354 VDD2.n71 VDD2.n58 4.26717
R1355 VDD2.n23 VDD2.n10 4.26717
R1356 VDD2.n93 VDD2.t0 3.7583
R1357 VDD2.n93 VDD2.t5 3.7583
R1358 VDD2.n45 VDD2.t4 3.7583
R1359 VDD2.n45 VDD2.t2 3.7583
R1360 VDD2.n72 VDD2.n56 3.49141
R1361 VDD2.n24 VDD2.n8 3.49141
R1362 VDD2.n76 VDD2.n75 2.71565
R1363 VDD2.n28 VDD2.n27 2.71565
R1364 VDD2.n65 VDD2.n61 2.41285
R1365 VDD2.n17 VDD2.n13 2.41285
R1366 VDD2.n91 VDD2.n47 1.93989
R1367 VDD2.n79 VDD2.n53 1.93989
R1368 VDD2.n32 VDD2.n6 1.93989
R1369 VDD2.n44 VDD2.n0 1.93989
R1370 VDD2.n89 VDD2.n88 1.16414
R1371 VDD2.n80 VDD2.n51 1.16414
R1372 VDD2.n33 VDD2.n4 1.16414
R1373 VDD2.n42 VDD2.n41 1.16414
R1374 VDD2 VDD2.n92 0.873345
R1375 VDD2.n85 VDD2.n49 0.388379
R1376 VDD2.n84 VDD2.n83 0.388379
R1377 VDD2.n37 VDD2.n36 0.388379
R1378 VDD2.n38 VDD2.n2 0.388379
R1379 VDD2.n90 VDD2.n48 0.155672
R1380 VDD2.n82 VDD2.n48 0.155672
R1381 VDD2.n82 VDD2.n81 0.155672
R1382 VDD2.n81 VDD2.n52 0.155672
R1383 VDD2.n74 VDD2.n52 0.155672
R1384 VDD2.n74 VDD2.n73 0.155672
R1385 VDD2.n73 VDD2.n57 0.155672
R1386 VDD2.n66 VDD2.n57 0.155672
R1387 VDD2.n66 VDD2.n65 0.155672
R1388 VDD2.n18 VDD2.n17 0.155672
R1389 VDD2.n18 VDD2.n9 0.155672
R1390 VDD2.n25 VDD2.n9 0.155672
R1391 VDD2.n26 VDD2.n25 0.155672
R1392 VDD2.n26 VDD2.n5 0.155672
R1393 VDD2.n34 VDD2.n5 0.155672
R1394 VDD2.n35 VDD2.n34 0.155672
R1395 VDD2.n35 VDD2.n1 0.155672
R1396 VDD2.n43 VDD2.n1 0.155672
C0 VTAIL B 2.23389f
C1 VN w_n1978_n2698# 3.27683f
C2 VTAIL VDD1 7.06391f
C3 VN VDD2 3.6547f
C4 VP w_n1978_n2698# 3.5279f
C5 VP VDD2 0.316533f
C6 w_n1978_n2698# VDD2 1.65975f
C7 VN B 0.774094f
C8 VN VDD1 0.148427f
C9 VN VTAIL 3.53664f
C10 VP B 1.18488f
C11 VP VDD1 3.81962f
C12 w_n1978_n2698# B 6.43131f
C13 VP VTAIL 3.55106f
C14 VDD2 B 1.41614f
C15 w_n1978_n2698# VDD1 1.62829f
C16 VDD1 VDD2 0.7936f
C17 VTAIL w_n1978_n2698# 2.41261f
C18 VTAIL VDD2 7.10199f
C19 VN VP 4.68216f
C20 VDD1 B 1.38176f
C21 VDD2 VSUBS 1.201746f
C22 VDD1 VSUBS 1.09961f
C23 VTAIL VSUBS 0.714841f
C24 VN VSUBS 4.30936f
C25 VP VSUBS 1.521214f
C26 B VSUBS 2.696717f
C27 w_n1978_n2698# VSUBS 66.1048f
C28 VDD2.n0 VSUBS 0.02418f
C29 VDD2.n1 VSUBS 0.022706f
C30 VDD2.n2 VSUBS 0.012201f
C31 VDD2.n3 VSUBS 0.028839f
C32 VDD2.n4 VSUBS 0.012919f
C33 VDD2.n5 VSUBS 0.022706f
C34 VDD2.n6 VSUBS 0.012201f
C35 VDD2.n7 VSUBS 0.028839f
C36 VDD2.n8 VSUBS 0.012919f
C37 VDD2.n9 VSUBS 0.022706f
C38 VDD2.n10 VSUBS 0.012201f
C39 VDD2.n11 VSUBS 0.028839f
C40 VDD2.n12 VSUBS 0.012919f
C41 VDD2.n13 VSUBS 0.144481f
C42 VDD2.t3 VSUBS 0.061951f
C43 VDD2.n14 VSUBS 0.021629f
C44 VDD2.n15 VSUBS 0.021694f
C45 VDD2.n16 VSUBS 0.012201f
C46 VDD2.n17 VSUBS 0.782201f
C47 VDD2.n18 VSUBS 0.022706f
C48 VDD2.n19 VSUBS 0.012201f
C49 VDD2.n20 VSUBS 0.012919f
C50 VDD2.n21 VSUBS 0.028839f
C51 VDD2.n22 VSUBS 0.028839f
C52 VDD2.n23 VSUBS 0.012919f
C53 VDD2.n24 VSUBS 0.012201f
C54 VDD2.n25 VSUBS 0.022706f
C55 VDD2.n26 VSUBS 0.022706f
C56 VDD2.n27 VSUBS 0.012201f
C57 VDD2.n28 VSUBS 0.012919f
C58 VDD2.n29 VSUBS 0.028839f
C59 VDD2.n30 VSUBS 0.028839f
C60 VDD2.n31 VSUBS 0.028839f
C61 VDD2.n32 VSUBS 0.012919f
C62 VDD2.n33 VSUBS 0.012201f
C63 VDD2.n34 VSUBS 0.022706f
C64 VDD2.n35 VSUBS 0.022706f
C65 VDD2.n36 VSUBS 0.012201f
C66 VDD2.n37 VSUBS 0.01256f
C67 VDD2.n38 VSUBS 0.01256f
C68 VDD2.n39 VSUBS 0.028839f
C69 VDD2.n40 VSUBS 0.067197f
C70 VDD2.n41 VSUBS 0.012919f
C71 VDD2.n42 VSUBS 0.012201f
C72 VDD2.n43 VSUBS 0.056515f
C73 VDD2.n44 VSUBS 0.050934f
C74 VDD2.t4 VSUBS 0.155204f
C75 VDD2.t2 VSUBS 0.155204f
C76 VDD2.n45 VSUBS 1.14504f
C77 VDD2.n46 VSUBS 1.79649f
C78 VDD2.n47 VSUBS 0.02418f
C79 VDD2.n48 VSUBS 0.022706f
C80 VDD2.n49 VSUBS 0.012201f
C81 VDD2.n50 VSUBS 0.028839f
C82 VDD2.n51 VSUBS 0.012919f
C83 VDD2.n52 VSUBS 0.022706f
C84 VDD2.n53 VSUBS 0.012201f
C85 VDD2.n54 VSUBS 0.028839f
C86 VDD2.n55 VSUBS 0.028839f
C87 VDD2.n56 VSUBS 0.012919f
C88 VDD2.n57 VSUBS 0.022706f
C89 VDD2.n58 VSUBS 0.012201f
C90 VDD2.n59 VSUBS 0.028839f
C91 VDD2.n60 VSUBS 0.012919f
C92 VDD2.n61 VSUBS 0.144481f
C93 VDD2.t1 VSUBS 0.061951f
C94 VDD2.n62 VSUBS 0.021629f
C95 VDD2.n63 VSUBS 0.021694f
C96 VDD2.n64 VSUBS 0.012201f
C97 VDD2.n65 VSUBS 0.782201f
C98 VDD2.n66 VSUBS 0.022706f
C99 VDD2.n67 VSUBS 0.012201f
C100 VDD2.n68 VSUBS 0.012919f
C101 VDD2.n69 VSUBS 0.028839f
C102 VDD2.n70 VSUBS 0.028839f
C103 VDD2.n71 VSUBS 0.012919f
C104 VDD2.n72 VSUBS 0.012201f
C105 VDD2.n73 VSUBS 0.022706f
C106 VDD2.n74 VSUBS 0.022706f
C107 VDD2.n75 VSUBS 0.012201f
C108 VDD2.n76 VSUBS 0.012919f
C109 VDD2.n77 VSUBS 0.028839f
C110 VDD2.n78 VSUBS 0.028839f
C111 VDD2.n79 VSUBS 0.012919f
C112 VDD2.n80 VSUBS 0.012201f
C113 VDD2.n81 VSUBS 0.022706f
C114 VDD2.n82 VSUBS 0.022706f
C115 VDD2.n83 VSUBS 0.012201f
C116 VDD2.n84 VSUBS 0.01256f
C117 VDD2.n85 VSUBS 0.01256f
C118 VDD2.n86 VSUBS 0.028839f
C119 VDD2.n87 VSUBS 0.067197f
C120 VDD2.n88 VSUBS 0.012919f
C121 VDD2.n89 VSUBS 0.012201f
C122 VDD2.n90 VSUBS 0.056515f
C123 VDD2.n91 VSUBS 0.049445f
C124 VDD2.n92 VSUBS 1.67597f
C125 VDD2.t0 VSUBS 0.155204f
C126 VDD2.t5 VSUBS 0.155204f
C127 VDD2.n93 VSUBS 1.14501f
C128 VN.n0 VSUBS 0.053302f
C129 VN.t1 VSUBS 1.15535f
C130 VN.n1 VSUBS 0.500994f
C131 VN.t2 VSUBS 1.26454f
C132 VN.n2 VSUBS 0.515688f
C133 VN.n3 VSUBS 0.226865f
C134 VN.n4 VSUBS 0.071169f
C135 VN.n5 VSUBS 0.018239f
C136 VN.t3 VSUBS 1.2313f
C137 VN.n6 VSUBS 0.509789f
C138 VN.n7 VSUBS 0.041307f
C139 VN.n8 VSUBS 0.053302f
C140 VN.t5 VSUBS 1.15535f
C141 VN.n9 VSUBS 0.500994f
C142 VN.t0 VSUBS 1.26454f
C143 VN.n10 VSUBS 0.515688f
C144 VN.n11 VSUBS 0.226865f
C145 VN.n12 VSUBS 0.071169f
C146 VN.n13 VSUBS 0.018239f
C147 VN.t4 VSUBS 1.2313f
C148 VN.n14 VSUBS 0.509789f
C149 VN.n15 VSUBS 2.02623f
C150 VDD1.n0 VSUBS 0.024216f
C151 VDD1.n1 VSUBS 0.022739f
C152 VDD1.n2 VSUBS 0.012219f
C153 VDD1.n3 VSUBS 0.028882f
C154 VDD1.n4 VSUBS 0.012938f
C155 VDD1.n5 VSUBS 0.022739f
C156 VDD1.n6 VSUBS 0.012219f
C157 VDD1.n7 VSUBS 0.028882f
C158 VDD1.n8 VSUBS 0.028882f
C159 VDD1.n9 VSUBS 0.012938f
C160 VDD1.n10 VSUBS 0.022739f
C161 VDD1.n11 VSUBS 0.012219f
C162 VDD1.n12 VSUBS 0.028882f
C163 VDD1.n13 VSUBS 0.012938f
C164 VDD1.n14 VSUBS 0.144695f
C165 VDD1.t4 VSUBS 0.062042f
C166 VDD1.n15 VSUBS 0.021661f
C167 VDD1.n16 VSUBS 0.021726f
C168 VDD1.n17 VSUBS 0.012219f
C169 VDD1.n18 VSUBS 0.78336f
C170 VDD1.n19 VSUBS 0.022739f
C171 VDD1.n20 VSUBS 0.012219f
C172 VDD1.n21 VSUBS 0.012938f
C173 VDD1.n22 VSUBS 0.028882f
C174 VDD1.n23 VSUBS 0.028882f
C175 VDD1.n24 VSUBS 0.012938f
C176 VDD1.n25 VSUBS 0.012219f
C177 VDD1.n26 VSUBS 0.022739f
C178 VDD1.n27 VSUBS 0.022739f
C179 VDD1.n28 VSUBS 0.012219f
C180 VDD1.n29 VSUBS 0.012938f
C181 VDD1.n30 VSUBS 0.028882f
C182 VDD1.n31 VSUBS 0.028882f
C183 VDD1.n32 VSUBS 0.012938f
C184 VDD1.n33 VSUBS 0.012219f
C185 VDD1.n34 VSUBS 0.022739f
C186 VDD1.n35 VSUBS 0.022739f
C187 VDD1.n36 VSUBS 0.012219f
C188 VDD1.n37 VSUBS 0.012578f
C189 VDD1.n38 VSUBS 0.012578f
C190 VDD1.n39 VSUBS 0.028882f
C191 VDD1.n40 VSUBS 0.067297f
C192 VDD1.n41 VSUBS 0.012938f
C193 VDD1.n42 VSUBS 0.012219f
C194 VDD1.n43 VSUBS 0.056599f
C195 VDD1.n44 VSUBS 0.051356f
C196 VDD1.n45 VSUBS 0.024216f
C197 VDD1.n46 VSUBS 0.022739f
C198 VDD1.n47 VSUBS 0.012219f
C199 VDD1.n48 VSUBS 0.028882f
C200 VDD1.n49 VSUBS 0.012938f
C201 VDD1.n50 VSUBS 0.022739f
C202 VDD1.n51 VSUBS 0.012219f
C203 VDD1.n52 VSUBS 0.028882f
C204 VDD1.n53 VSUBS 0.012938f
C205 VDD1.n54 VSUBS 0.022739f
C206 VDD1.n55 VSUBS 0.012219f
C207 VDD1.n56 VSUBS 0.028882f
C208 VDD1.n57 VSUBS 0.012938f
C209 VDD1.n58 VSUBS 0.144695f
C210 VDD1.t5 VSUBS 0.062042f
C211 VDD1.n59 VSUBS 0.021661f
C212 VDD1.n60 VSUBS 0.021726f
C213 VDD1.n61 VSUBS 0.012219f
C214 VDD1.n62 VSUBS 0.78336f
C215 VDD1.n63 VSUBS 0.022739f
C216 VDD1.n64 VSUBS 0.012219f
C217 VDD1.n65 VSUBS 0.012938f
C218 VDD1.n66 VSUBS 0.028882f
C219 VDD1.n67 VSUBS 0.028882f
C220 VDD1.n68 VSUBS 0.012938f
C221 VDD1.n69 VSUBS 0.012219f
C222 VDD1.n70 VSUBS 0.022739f
C223 VDD1.n71 VSUBS 0.022739f
C224 VDD1.n72 VSUBS 0.012219f
C225 VDD1.n73 VSUBS 0.012938f
C226 VDD1.n74 VSUBS 0.028882f
C227 VDD1.n75 VSUBS 0.028882f
C228 VDD1.n76 VSUBS 0.028882f
C229 VDD1.n77 VSUBS 0.012938f
C230 VDD1.n78 VSUBS 0.012219f
C231 VDD1.n79 VSUBS 0.022739f
C232 VDD1.n80 VSUBS 0.022739f
C233 VDD1.n81 VSUBS 0.012219f
C234 VDD1.n82 VSUBS 0.012578f
C235 VDD1.n83 VSUBS 0.012578f
C236 VDD1.n84 VSUBS 0.028882f
C237 VDD1.n85 VSUBS 0.067297f
C238 VDD1.n86 VSUBS 0.012938f
C239 VDD1.n87 VSUBS 0.012219f
C240 VDD1.n88 VSUBS 0.056599f
C241 VDD1.n89 VSUBS 0.05101f
C242 VDD1.t1 VSUBS 0.155434f
C243 VDD1.t2 VSUBS 0.155434f
C244 VDD1.n90 VSUBS 1.14673f
C245 VDD1.n91 VSUBS 1.87282f
C246 VDD1.t0 VSUBS 0.155434f
C247 VDD1.t3 VSUBS 0.155434f
C248 VDD1.n92 VSUBS 1.14544f
C249 VDD1.n93 VSUBS 2.0745f
C250 VTAIL.t0 VSUBS 0.203128f
C251 VTAIL.t4 VSUBS 0.203128f
C252 VTAIL.n0 VSUBS 1.36936f
C253 VTAIL.n1 VSUBS 0.727231f
C254 VTAIL.n2 VSUBS 0.031646f
C255 VTAIL.n3 VSUBS 0.029717f
C256 VTAIL.n4 VSUBS 0.015968f
C257 VTAIL.n5 VSUBS 0.037744f
C258 VTAIL.n6 VSUBS 0.016908f
C259 VTAIL.n7 VSUBS 0.029717f
C260 VTAIL.n8 VSUBS 0.015968f
C261 VTAIL.n9 VSUBS 0.037744f
C262 VTAIL.n10 VSUBS 0.016908f
C263 VTAIL.n11 VSUBS 0.029717f
C264 VTAIL.n12 VSUBS 0.015968f
C265 VTAIL.n13 VSUBS 0.037744f
C266 VTAIL.n14 VSUBS 0.016908f
C267 VTAIL.n15 VSUBS 0.189094f
C268 VTAIL.t7 VSUBS 0.08108f
C269 VTAIL.n16 VSUBS 0.028308f
C270 VTAIL.n17 VSUBS 0.028393f
C271 VTAIL.n18 VSUBS 0.015968f
C272 VTAIL.n19 VSUBS 1.02373f
C273 VTAIL.n20 VSUBS 0.029717f
C274 VTAIL.n21 VSUBS 0.015968f
C275 VTAIL.n22 VSUBS 0.016908f
C276 VTAIL.n23 VSUBS 0.037744f
C277 VTAIL.n24 VSUBS 0.037744f
C278 VTAIL.n25 VSUBS 0.016908f
C279 VTAIL.n26 VSUBS 0.015968f
C280 VTAIL.n27 VSUBS 0.029717f
C281 VTAIL.n28 VSUBS 0.029717f
C282 VTAIL.n29 VSUBS 0.015968f
C283 VTAIL.n30 VSUBS 0.016908f
C284 VTAIL.n31 VSUBS 0.037744f
C285 VTAIL.n32 VSUBS 0.037744f
C286 VTAIL.n33 VSUBS 0.037744f
C287 VTAIL.n34 VSUBS 0.016908f
C288 VTAIL.n35 VSUBS 0.015968f
C289 VTAIL.n36 VSUBS 0.029717f
C290 VTAIL.n37 VSUBS 0.029717f
C291 VTAIL.n38 VSUBS 0.015968f
C292 VTAIL.n39 VSUBS 0.016438f
C293 VTAIL.n40 VSUBS 0.016438f
C294 VTAIL.n41 VSUBS 0.037744f
C295 VTAIL.n42 VSUBS 0.087947f
C296 VTAIL.n43 VSUBS 0.016908f
C297 VTAIL.n44 VSUBS 0.015968f
C298 VTAIL.n45 VSUBS 0.073966f
C299 VTAIL.n46 VSUBS 0.044232f
C300 VTAIL.n47 VSUBS 0.229365f
C301 VTAIL.t9 VSUBS 0.203128f
C302 VTAIL.t11 VSUBS 0.203128f
C303 VTAIL.n48 VSUBS 1.36936f
C304 VTAIL.n49 VSUBS 2.02838f
C305 VTAIL.t2 VSUBS 0.203128f
C306 VTAIL.t3 VSUBS 0.203128f
C307 VTAIL.n50 VSUBS 1.36937f
C308 VTAIL.n51 VSUBS 2.02837f
C309 VTAIL.n52 VSUBS 0.031646f
C310 VTAIL.n53 VSUBS 0.029717f
C311 VTAIL.n54 VSUBS 0.015968f
C312 VTAIL.n55 VSUBS 0.037744f
C313 VTAIL.n56 VSUBS 0.016908f
C314 VTAIL.n57 VSUBS 0.029717f
C315 VTAIL.n58 VSUBS 0.015968f
C316 VTAIL.n59 VSUBS 0.037744f
C317 VTAIL.n60 VSUBS 0.037744f
C318 VTAIL.n61 VSUBS 0.016908f
C319 VTAIL.n62 VSUBS 0.029717f
C320 VTAIL.n63 VSUBS 0.015968f
C321 VTAIL.n64 VSUBS 0.037744f
C322 VTAIL.n65 VSUBS 0.016908f
C323 VTAIL.n66 VSUBS 0.189094f
C324 VTAIL.t5 VSUBS 0.08108f
C325 VTAIL.n67 VSUBS 0.028308f
C326 VTAIL.n68 VSUBS 0.028393f
C327 VTAIL.n69 VSUBS 0.015968f
C328 VTAIL.n70 VSUBS 1.02373f
C329 VTAIL.n71 VSUBS 0.029717f
C330 VTAIL.n72 VSUBS 0.015968f
C331 VTAIL.n73 VSUBS 0.016908f
C332 VTAIL.n74 VSUBS 0.037744f
C333 VTAIL.n75 VSUBS 0.037744f
C334 VTAIL.n76 VSUBS 0.016908f
C335 VTAIL.n77 VSUBS 0.015968f
C336 VTAIL.n78 VSUBS 0.029717f
C337 VTAIL.n79 VSUBS 0.029717f
C338 VTAIL.n80 VSUBS 0.015968f
C339 VTAIL.n81 VSUBS 0.016908f
C340 VTAIL.n82 VSUBS 0.037744f
C341 VTAIL.n83 VSUBS 0.037744f
C342 VTAIL.n84 VSUBS 0.016908f
C343 VTAIL.n85 VSUBS 0.015968f
C344 VTAIL.n86 VSUBS 0.029717f
C345 VTAIL.n87 VSUBS 0.029717f
C346 VTAIL.n88 VSUBS 0.015968f
C347 VTAIL.n89 VSUBS 0.016438f
C348 VTAIL.n90 VSUBS 0.016438f
C349 VTAIL.n91 VSUBS 0.037744f
C350 VTAIL.n92 VSUBS 0.087947f
C351 VTAIL.n93 VSUBS 0.016908f
C352 VTAIL.n94 VSUBS 0.015968f
C353 VTAIL.n95 VSUBS 0.073966f
C354 VTAIL.n96 VSUBS 0.044232f
C355 VTAIL.n97 VSUBS 0.229365f
C356 VTAIL.t6 VSUBS 0.203128f
C357 VTAIL.t10 VSUBS 0.203128f
C358 VTAIL.n98 VSUBS 1.36937f
C359 VTAIL.n99 VSUBS 0.799657f
C360 VTAIL.n100 VSUBS 0.031646f
C361 VTAIL.n101 VSUBS 0.029717f
C362 VTAIL.n102 VSUBS 0.015968f
C363 VTAIL.n103 VSUBS 0.037744f
C364 VTAIL.n104 VSUBS 0.016908f
C365 VTAIL.n105 VSUBS 0.029717f
C366 VTAIL.n106 VSUBS 0.015968f
C367 VTAIL.n107 VSUBS 0.037744f
C368 VTAIL.n108 VSUBS 0.037744f
C369 VTAIL.n109 VSUBS 0.016908f
C370 VTAIL.n110 VSUBS 0.029717f
C371 VTAIL.n111 VSUBS 0.015968f
C372 VTAIL.n112 VSUBS 0.037744f
C373 VTAIL.n113 VSUBS 0.016908f
C374 VTAIL.n114 VSUBS 0.189094f
C375 VTAIL.t8 VSUBS 0.08108f
C376 VTAIL.n115 VSUBS 0.028308f
C377 VTAIL.n116 VSUBS 0.028393f
C378 VTAIL.n117 VSUBS 0.015968f
C379 VTAIL.n118 VSUBS 1.02373f
C380 VTAIL.n119 VSUBS 0.029717f
C381 VTAIL.n120 VSUBS 0.015968f
C382 VTAIL.n121 VSUBS 0.016908f
C383 VTAIL.n122 VSUBS 0.037744f
C384 VTAIL.n123 VSUBS 0.037744f
C385 VTAIL.n124 VSUBS 0.016908f
C386 VTAIL.n125 VSUBS 0.015968f
C387 VTAIL.n126 VSUBS 0.029717f
C388 VTAIL.n127 VSUBS 0.029717f
C389 VTAIL.n128 VSUBS 0.015968f
C390 VTAIL.n129 VSUBS 0.016908f
C391 VTAIL.n130 VSUBS 0.037744f
C392 VTAIL.n131 VSUBS 0.037744f
C393 VTAIL.n132 VSUBS 0.016908f
C394 VTAIL.n133 VSUBS 0.015968f
C395 VTAIL.n134 VSUBS 0.029717f
C396 VTAIL.n135 VSUBS 0.029717f
C397 VTAIL.n136 VSUBS 0.015968f
C398 VTAIL.n137 VSUBS 0.016438f
C399 VTAIL.n138 VSUBS 0.016438f
C400 VTAIL.n139 VSUBS 0.037744f
C401 VTAIL.n140 VSUBS 0.087947f
C402 VTAIL.n141 VSUBS 0.016908f
C403 VTAIL.n142 VSUBS 0.015968f
C404 VTAIL.n143 VSUBS 0.073966f
C405 VTAIL.n144 VSUBS 0.044232f
C406 VTAIL.n145 VSUBS 1.35407f
C407 VTAIL.n146 VSUBS 0.031646f
C408 VTAIL.n147 VSUBS 0.029717f
C409 VTAIL.n148 VSUBS 0.015968f
C410 VTAIL.n149 VSUBS 0.037744f
C411 VTAIL.n150 VSUBS 0.016908f
C412 VTAIL.n151 VSUBS 0.029717f
C413 VTAIL.n152 VSUBS 0.015968f
C414 VTAIL.n153 VSUBS 0.037744f
C415 VTAIL.n154 VSUBS 0.016908f
C416 VTAIL.n155 VSUBS 0.029717f
C417 VTAIL.n156 VSUBS 0.015968f
C418 VTAIL.n157 VSUBS 0.037744f
C419 VTAIL.n158 VSUBS 0.016908f
C420 VTAIL.n159 VSUBS 0.189094f
C421 VTAIL.t1 VSUBS 0.08108f
C422 VTAIL.n160 VSUBS 0.028308f
C423 VTAIL.n161 VSUBS 0.028393f
C424 VTAIL.n162 VSUBS 0.015968f
C425 VTAIL.n163 VSUBS 1.02373f
C426 VTAIL.n164 VSUBS 0.029717f
C427 VTAIL.n165 VSUBS 0.015968f
C428 VTAIL.n166 VSUBS 0.016908f
C429 VTAIL.n167 VSUBS 0.037744f
C430 VTAIL.n168 VSUBS 0.037744f
C431 VTAIL.n169 VSUBS 0.016908f
C432 VTAIL.n170 VSUBS 0.015968f
C433 VTAIL.n171 VSUBS 0.029717f
C434 VTAIL.n172 VSUBS 0.029717f
C435 VTAIL.n173 VSUBS 0.015968f
C436 VTAIL.n174 VSUBS 0.016908f
C437 VTAIL.n175 VSUBS 0.037744f
C438 VTAIL.n176 VSUBS 0.037744f
C439 VTAIL.n177 VSUBS 0.037744f
C440 VTAIL.n178 VSUBS 0.016908f
C441 VTAIL.n179 VSUBS 0.015968f
C442 VTAIL.n180 VSUBS 0.029717f
C443 VTAIL.n181 VSUBS 0.029717f
C444 VTAIL.n182 VSUBS 0.015968f
C445 VTAIL.n183 VSUBS 0.016438f
C446 VTAIL.n184 VSUBS 0.016438f
C447 VTAIL.n185 VSUBS 0.037744f
C448 VTAIL.n186 VSUBS 0.087947f
C449 VTAIL.n187 VSUBS 0.016908f
C450 VTAIL.n188 VSUBS 0.015968f
C451 VTAIL.n189 VSUBS 0.073966f
C452 VTAIL.n190 VSUBS 0.044232f
C453 VTAIL.n191 VSUBS 1.3225f
C454 VP.n0 VSUBS 0.054975f
C455 VP.t4 VSUBS 1.19163f
C456 VP.n1 VSUBS 0.463716f
C457 VP.n2 VSUBS 0.054975f
C458 VP.n3 VSUBS 0.054975f
C459 VP.t2 VSUBS 1.26996f
C460 VP.t5 VSUBS 1.19163f
C461 VP.n4 VSUBS 0.516725f
C462 VP.t1 VSUBS 1.30425f
C463 VP.n5 VSUBS 0.531881f
C464 VP.n6 VSUBS 0.233989f
C465 VP.n7 VSUBS 0.073404f
C466 VP.n8 VSUBS 0.018812f
C467 VP.n9 VSUBS 0.525796f
C468 VP.n10 VSUBS 2.05363f
C469 VP.n11 VSUBS 2.10352f
C470 VP.t0 VSUBS 1.26996f
C471 VP.n12 VSUBS 0.525796f
C472 VP.n13 VSUBS 0.018812f
C473 VP.n14 VSUBS 0.073404f
C474 VP.n15 VSUBS 0.054975f
C475 VP.n16 VSUBS 0.054975f
C476 VP.n17 VSUBS 0.073404f
C477 VP.n18 VSUBS 0.018812f
C478 VP.t3 VSUBS 1.26996f
C479 VP.n19 VSUBS 0.525796f
C480 VP.n20 VSUBS 0.042604f
C481 B.n0 VSUBS 0.004825f
C482 B.n1 VSUBS 0.004825f
C483 B.n2 VSUBS 0.00763f
C484 B.n3 VSUBS 0.00763f
C485 B.n4 VSUBS 0.00763f
C486 B.n5 VSUBS 0.00763f
C487 B.n6 VSUBS 0.00763f
C488 B.n7 VSUBS 0.00763f
C489 B.n8 VSUBS 0.00763f
C490 B.n9 VSUBS 0.00763f
C491 B.n10 VSUBS 0.00763f
C492 B.n11 VSUBS 0.00763f
C493 B.n12 VSUBS 0.00763f
C494 B.n13 VSUBS 0.017384f
C495 B.n14 VSUBS 0.00763f
C496 B.n15 VSUBS 0.00763f
C497 B.n16 VSUBS 0.00763f
C498 B.n17 VSUBS 0.00763f
C499 B.n18 VSUBS 0.00763f
C500 B.n19 VSUBS 0.00763f
C501 B.n20 VSUBS 0.00763f
C502 B.n21 VSUBS 0.00763f
C503 B.n22 VSUBS 0.00763f
C504 B.n23 VSUBS 0.00763f
C505 B.n24 VSUBS 0.00763f
C506 B.n25 VSUBS 0.00763f
C507 B.n26 VSUBS 0.00763f
C508 B.n27 VSUBS 0.00763f
C509 B.n28 VSUBS 0.00763f
C510 B.n29 VSUBS 0.00763f
C511 B.t5 VSUBS 0.152113f
C512 B.t4 VSUBS 0.16664f
C513 B.t3 VSUBS 0.377847f
C514 B.n30 VSUBS 0.267254f
C515 B.n31 VSUBS 0.212849f
C516 B.n32 VSUBS 0.00763f
C517 B.n33 VSUBS 0.00763f
C518 B.n34 VSUBS 0.00763f
C519 B.n35 VSUBS 0.00763f
C520 B.t2 VSUBS 0.152116f
C521 B.t1 VSUBS 0.166642f
C522 B.t0 VSUBS 0.377847f
C523 B.n36 VSUBS 0.267252f
C524 B.n37 VSUBS 0.212846f
C525 B.n38 VSUBS 0.017678f
C526 B.n39 VSUBS 0.00763f
C527 B.n40 VSUBS 0.00763f
C528 B.n41 VSUBS 0.00763f
C529 B.n42 VSUBS 0.00763f
C530 B.n43 VSUBS 0.00763f
C531 B.n44 VSUBS 0.00763f
C532 B.n45 VSUBS 0.00763f
C533 B.n46 VSUBS 0.00763f
C534 B.n47 VSUBS 0.00763f
C535 B.n48 VSUBS 0.00763f
C536 B.n49 VSUBS 0.00763f
C537 B.n50 VSUBS 0.00763f
C538 B.n51 VSUBS 0.00763f
C539 B.n52 VSUBS 0.00763f
C540 B.n53 VSUBS 0.00763f
C541 B.n54 VSUBS 0.017162f
C542 B.n55 VSUBS 0.00763f
C543 B.n56 VSUBS 0.00763f
C544 B.n57 VSUBS 0.00763f
C545 B.n58 VSUBS 0.00763f
C546 B.n59 VSUBS 0.00763f
C547 B.n60 VSUBS 0.00763f
C548 B.n61 VSUBS 0.00763f
C549 B.n62 VSUBS 0.00763f
C550 B.n63 VSUBS 0.00763f
C551 B.n64 VSUBS 0.00763f
C552 B.n65 VSUBS 0.00763f
C553 B.n66 VSUBS 0.00763f
C554 B.n67 VSUBS 0.00763f
C555 B.n68 VSUBS 0.00763f
C556 B.n69 VSUBS 0.00763f
C557 B.n70 VSUBS 0.00763f
C558 B.n71 VSUBS 0.00763f
C559 B.n72 VSUBS 0.00763f
C560 B.n73 VSUBS 0.00763f
C561 B.n74 VSUBS 0.00763f
C562 B.n75 VSUBS 0.00763f
C563 B.n76 VSUBS 0.00763f
C564 B.n77 VSUBS 0.00763f
C565 B.n78 VSUBS 0.018073f
C566 B.n79 VSUBS 0.00763f
C567 B.n80 VSUBS 0.00763f
C568 B.n81 VSUBS 0.00763f
C569 B.n82 VSUBS 0.00763f
C570 B.n83 VSUBS 0.00763f
C571 B.n84 VSUBS 0.00763f
C572 B.n85 VSUBS 0.00763f
C573 B.n86 VSUBS 0.00763f
C574 B.n87 VSUBS 0.00763f
C575 B.n88 VSUBS 0.00763f
C576 B.n89 VSUBS 0.00763f
C577 B.n90 VSUBS 0.00763f
C578 B.n91 VSUBS 0.00763f
C579 B.n92 VSUBS 0.00763f
C580 B.n93 VSUBS 0.00763f
C581 B.t7 VSUBS 0.152116f
C582 B.t8 VSUBS 0.166642f
C583 B.t6 VSUBS 0.377847f
C584 B.n94 VSUBS 0.267252f
C585 B.n95 VSUBS 0.212846f
C586 B.n96 VSUBS 0.017678f
C587 B.n97 VSUBS 0.00763f
C588 B.n98 VSUBS 0.00763f
C589 B.n99 VSUBS 0.00763f
C590 B.n100 VSUBS 0.00763f
C591 B.n101 VSUBS 0.00763f
C592 B.t10 VSUBS 0.152113f
C593 B.t11 VSUBS 0.16664f
C594 B.t9 VSUBS 0.377847f
C595 B.n102 VSUBS 0.267254f
C596 B.n103 VSUBS 0.212849f
C597 B.n104 VSUBS 0.00763f
C598 B.n105 VSUBS 0.00763f
C599 B.n106 VSUBS 0.00763f
C600 B.n107 VSUBS 0.00763f
C601 B.n108 VSUBS 0.00763f
C602 B.n109 VSUBS 0.00763f
C603 B.n110 VSUBS 0.00763f
C604 B.n111 VSUBS 0.00763f
C605 B.n112 VSUBS 0.00763f
C606 B.n113 VSUBS 0.00763f
C607 B.n114 VSUBS 0.00763f
C608 B.n115 VSUBS 0.00763f
C609 B.n116 VSUBS 0.00763f
C610 B.n117 VSUBS 0.00763f
C611 B.n118 VSUBS 0.00763f
C612 B.n119 VSUBS 0.017384f
C613 B.n120 VSUBS 0.00763f
C614 B.n121 VSUBS 0.00763f
C615 B.n122 VSUBS 0.00763f
C616 B.n123 VSUBS 0.00763f
C617 B.n124 VSUBS 0.00763f
C618 B.n125 VSUBS 0.00763f
C619 B.n126 VSUBS 0.00763f
C620 B.n127 VSUBS 0.00763f
C621 B.n128 VSUBS 0.00763f
C622 B.n129 VSUBS 0.00763f
C623 B.n130 VSUBS 0.00763f
C624 B.n131 VSUBS 0.00763f
C625 B.n132 VSUBS 0.00763f
C626 B.n133 VSUBS 0.00763f
C627 B.n134 VSUBS 0.00763f
C628 B.n135 VSUBS 0.00763f
C629 B.n136 VSUBS 0.00763f
C630 B.n137 VSUBS 0.00763f
C631 B.n138 VSUBS 0.00763f
C632 B.n139 VSUBS 0.00763f
C633 B.n140 VSUBS 0.00763f
C634 B.n141 VSUBS 0.00763f
C635 B.n142 VSUBS 0.00763f
C636 B.n143 VSUBS 0.00763f
C637 B.n144 VSUBS 0.00763f
C638 B.n145 VSUBS 0.00763f
C639 B.n146 VSUBS 0.00763f
C640 B.n147 VSUBS 0.00763f
C641 B.n148 VSUBS 0.00763f
C642 B.n149 VSUBS 0.00763f
C643 B.n150 VSUBS 0.00763f
C644 B.n151 VSUBS 0.00763f
C645 B.n152 VSUBS 0.00763f
C646 B.n153 VSUBS 0.00763f
C647 B.n154 VSUBS 0.00763f
C648 B.n155 VSUBS 0.00763f
C649 B.n156 VSUBS 0.00763f
C650 B.n157 VSUBS 0.00763f
C651 B.n158 VSUBS 0.00763f
C652 B.n159 VSUBS 0.00763f
C653 B.n160 VSUBS 0.00763f
C654 B.n161 VSUBS 0.00763f
C655 B.n162 VSUBS 0.017384f
C656 B.n163 VSUBS 0.018073f
C657 B.n164 VSUBS 0.018073f
C658 B.n165 VSUBS 0.00763f
C659 B.n166 VSUBS 0.00763f
C660 B.n167 VSUBS 0.00763f
C661 B.n168 VSUBS 0.00763f
C662 B.n169 VSUBS 0.00763f
C663 B.n170 VSUBS 0.00763f
C664 B.n171 VSUBS 0.00763f
C665 B.n172 VSUBS 0.00763f
C666 B.n173 VSUBS 0.00763f
C667 B.n174 VSUBS 0.00763f
C668 B.n175 VSUBS 0.00763f
C669 B.n176 VSUBS 0.00763f
C670 B.n177 VSUBS 0.00763f
C671 B.n178 VSUBS 0.00763f
C672 B.n179 VSUBS 0.00763f
C673 B.n180 VSUBS 0.00763f
C674 B.n181 VSUBS 0.00763f
C675 B.n182 VSUBS 0.00763f
C676 B.n183 VSUBS 0.00763f
C677 B.n184 VSUBS 0.00763f
C678 B.n185 VSUBS 0.00763f
C679 B.n186 VSUBS 0.00763f
C680 B.n187 VSUBS 0.00763f
C681 B.n188 VSUBS 0.00763f
C682 B.n189 VSUBS 0.00763f
C683 B.n190 VSUBS 0.00763f
C684 B.n191 VSUBS 0.00763f
C685 B.n192 VSUBS 0.00763f
C686 B.n193 VSUBS 0.00763f
C687 B.n194 VSUBS 0.00763f
C688 B.n195 VSUBS 0.00763f
C689 B.n196 VSUBS 0.00763f
C690 B.n197 VSUBS 0.00763f
C691 B.n198 VSUBS 0.00763f
C692 B.n199 VSUBS 0.00763f
C693 B.n200 VSUBS 0.00763f
C694 B.n201 VSUBS 0.00763f
C695 B.n202 VSUBS 0.00763f
C696 B.n203 VSUBS 0.00763f
C697 B.n204 VSUBS 0.00763f
C698 B.n205 VSUBS 0.00763f
C699 B.n206 VSUBS 0.00763f
C700 B.n207 VSUBS 0.00763f
C701 B.n208 VSUBS 0.00763f
C702 B.n209 VSUBS 0.00763f
C703 B.n210 VSUBS 0.005274f
C704 B.n211 VSUBS 0.017678f
C705 B.n212 VSUBS 0.006171f
C706 B.n213 VSUBS 0.00763f
C707 B.n214 VSUBS 0.00763f
C708 B.n215 VSUBS 0.00763f
C709 B.n216 VSUBS 0.00763f
C710 B.n217 VSUBS 0.00763f
C711 B.n218 VSUBS 0.00763f
C712 B.n219 VSUBS 0.00763f
C713 B.n220 VSUBS 0.00763f
C714 B.n221 VSUBS 0.00763f
C715 B.n222 VSUBS 0.00763f
C716 B.n223 VSUBS 0.00763f
C717 B.n224 VSUBS 0.006171f
C718 B.n225 VSUBS 0.00763f
C719 B.n226 VSUBS 0.00763f
C720 B.n227 VSUBS 0.005274f
C721 B.n228 VSUBS 0.00763f
C722 B.n229 VSUBS 0.00763f
C723 B.n230 VSUBS 0.00763f
C724 B.n231 VSUBS 0.00763f
C725 B.n232 VSUBS 0.00763f
C726 B.n233 VSUBS 0.00763f
C727 B.n234 VSUBS 0.00763f
C728 B.n235 VSUBS 0.00763f
C729 B.n236 VSUBS 0.00763f
C730 B.n237 VSUBS 0.00763f
C731 B.n238 VSUBS 0.00763f
C732 B.n239 VSUBS 0.00763f
C733 B.n240 VSUBS 0.00763f
C734 B.n241 VSUBS 0.00763f
C735 B.n242 VSUBS 0.00763f
C736 B.n243 VSUBS 0.00763f
C737 B.n244 VSUBS 0.00763f
C738 B.n245 VSUBS 0.00763f
C739 B.n246 VSUBS 0.00763f
C740 B.n247 VSUBS 0.00763f
C741 B.n248 VSUBS 0.00763f
C742 B.n249 VSUBS 0.00763f
C743 B.n250 VSUBS 0.00763f
C744 B.n251 VSUBS 0.00763f
C745 B.n252 VSUBS 0.00763f
C746 B.n253 VSUBS 0.00763f
C747 B.n254 VSUBS 0.00763f
C748 B.n255 VSUBS 0.00763f
C749 B.n256 VSUBS 0.00763f
C750 B.n257 VSUBS 0.00763f
C751 B.n258 VSUBS 0.00763f
C752 B.n259 VSUBS 0.00763f
C753 B.n260 VSUBS 0.00763f
C754 B.n261 VSUBS 0.00763f
C755 B.n262 VSUBS 0.00763f
C756 B.n263 VSUBS 0.00763f
C757 B.n264 VSUBS 0.00763f
C758 B.n265 VSUBS 0.00763f
C759 B.n266 VSUBS 0.00763f
C760 B.n267 VSUBS 0.00763f
C761 B.n268 VSUBS 0.00763f
C762 B.n269 VSUBS 0.00763f
C763 B.n270 VSUBS 0.00763f
C764 B.n271 VSUBS 0.00763f
C765 B.n272 VSUBS 0.00763f
C766 B.n273 VSUBS 0.018073f
C767 B.n274 VSUBS 0.017384f
C768 B.n275 VSUBS 0.017384f
C769 B.n276 VSUBS 0.00763f
C770 B.n277 VSUBS 0.00763f
C771 B.n278 VSUBS 0.00763f
C772 B.n279 VSUBS 0.00763f
C773 B.n280 VSUBS 0.00763f
C774 B.n281 VSUBS 0.00763f
C775 B.n282 VSUBS 0.00763f
C776 B.n283 VSUBS 0.00763f
C777 B.n284 VSUBS 0.00763f
C778 B.n285 VSUBS 0.00763f
C779 B.n286 VSUBS 0.00763f
C780 B.n287 VSUBS 0.00763f
C781 B.n288 VSUBS 0.00763f
C782 B.n289 VSUBS 0.00763f
C783 B.n290 VSUBS 0.00763f
C784 B.n291 VSUBS 0.00763f
C785 B.n292 VSUBS 0.00763f
C786 B.n293 VSUBS 0.00763f
C787 B.n294 VSUBS 0.00763f
C788 B.n295 VSUBS 0.00763f
C789 B.n296 VSUBS 0.00763f
C790 B.n297 VSUBS 0.00763f
C791 B.n298 VSUBS 0.00763f
C792 B.n299 VSUBS 0.00763f
C793 B.n300 VSUBS 0.00763f
C794 B.n301 VSUBS 0.00763f
C795 B.n302 VSUBS 0.00763f
C796 B.n303 VSUBS 0.00763f
C797 B.n304 VSUBS 0.00763f
C798 B.n305 VSUBS 0.00763f
C799 B.n306 VSUBS 0.00763f
C800 B.n307 VSUBS 0.00763f
C801 B.n308 VSUBS 0.00763f
C802 B.n309 VSUBS 0.00763f
C803 B.n310 VSUBS 0.00763f
C804 B.n311 VSUBS 0.00763f
C805 B.n312 VSUBS 0.00763f
C806 B.n313 VSUBS 0.00763f
C807 B.n314 VSUBS 0.00763f
C808 B.n315 VSUBS 0.00763f
C809 B.n316 VSUBS 0.00763f
C810 B.n317 VSUBS 0.00763f
C811 B.n318 VSUBS 0.00763f
C812 B.n319 VSUBS 0.00763f
C813 B.n320 VSUBS 0.00763f
C814 B.n321 VSUBS 0.00763f
C815 B.n322 VSUBS 0.00763f
C816 B.n323 VSUBS 0.00763f
C817 B.n324 VSUBS 0.00763f
C818 B.n325 VSUBS 0.00763f
C819 B.n326 VSUBS 0.00763f
C820 B.n327 VSUBS 0.00763f
C821 B.n328 VSUBS 0.00763f
C822 B.n329 VSUBS 0.00763f
C823 B.n330 VSUBS 0.00763f
C824 B.n331 VSUBS 0.00763f
C825 B.n332 VSUBS 0.00763f
C826 B.n333 VSUBS 0.00763f
C827 B.n334 VSUBS 0.00763f
C828 B.n335 VSUBS 0.00763f
C829 B.n336 VSUBS 0.00763f
C830 B.n337 VSUBS 0.00763f
C831 B.n338 VSUBS 0.00763f
C832 B.n339 VSUBS 0.00763f
C833 B.n340 VSUBS 0.00763f
C834 B.n341 VSUBS 0.00763f
C835 B.n342 VSUBS 0.00763f
C836 B.n343 VSUBS 0.018296f
C837 B.n344 VSUBS 0.017384f
C838 B.n345 VSUBS 0.018073f
C839 B.n346 VSUBS 0.00763f
C840 B.n347 VSUBS 0.00763f
C841 B.n348 VSUBS 0.00763f
C842 B.n349 VSUBS 0.00763f
C843 B.n350 VSUBS 0.00763f
C844 B.n351 VSUBS 0.00763f
C845 B.n352 VSUBS 0.00763f
C846 B.n353 VSUBS 0.00763f
C847 B.n354 VSUBS 0.00763f
C848 B.n355 VSUBS 0.00763f
C849 B.n356 VSUBS 0.00763f
C850 B.n357 VSUBS 0.00763f
C851 B.n358 VSUBS 0.00763f
C852 B.n359 VSUBS 0.00763f
C853 B.n360 VSUBS 0.00763f
C854 B.n361 VSUBS 0.00763f
C855 B.n362 VSUBS 0.00763f
C856 B.n363 VSUBS 0.00763f
C857 B.n364 VSUBS 0.00763f
C858 B.n365 VSUBS 0.00763f
C859 B.n366 VSUBS 0.00763f
C860 B.n367 VSUBS 0.00763f
C861 B.n368 VSUBS 0.00763f
C862 B.n369 VSUBS 0.00763f
C863 B.n370 VSUBS 0.00763f
C864 B.n371 VSUBS 0.00763f
C865 B.n372 VSUBS 0.00763f
C866 B.n373 VSUBS 0.00763f
C867 B.n374 VSUBS 0.00763f
C868 B.n375 VSUBS 0.00763f
C869 B.n376 VSUBS 0.00763f
C870 B.n377 VSUBS 0.00763f
C871 B.n378 VSUBS 0.00763f
C872 B.n379 VSUBS 0.00763f
C873 B.n380 VSUBS 0.00763f
C874 B.n381 VSUBS 0.00763f
C875 B.n382 VSUBS 0.00763f
C876 B.n383 VSUBS 0.00763f
C877 B.n384 VSUBS 0.00763f
C878 B.n385 VSUBS 0.00763f
C879 B.n386 VSUBS 0.00763f
C880 B.n387 VSUBS 0.00763f
C881 B.n388 VSUBS 0.00763f
C882 B.n389 VSUBS 0.00763f
C883 B.n390 VSUBS 0.00763f
C884 B.n391 VSUBS 0.005274f
C885 B.n392 VSUBS 0.00763f
C886 B.n393 VSUBS 0.00763f
C887 B.n394 VSUBS 0.006171f
C888 B.n395 VSUBS 0.00763f
C889 B.n396 VSUBS 0.00763f
C890 B.n397 VSUBS 0.00763f
C891 B.n398 VSUBS 0.00763f
C892 B.n399 VSUBS 0.00763f
C893 B.n400 VSUBS 0.00763f
C894 B.n401 VSUBS 0.00763f
C895 B.n402 VSUBS 0.00763f
C896 B.n403 VSUBS 0.00763f
C897 B.n404 VSUBS 0.00763f
C898 B.n405 VSUBS 0.00763f
C899 B.n406 VSUBS 0.006171f
C900 B.n407 VSUBS 0.017678f
C901 B.n408 VSUBS 0.005274f
C902 B.n409 VSUBS 0.00763f
C903 B.n410 VSUBS 0.00763f
C904 B.n411 VSUBS 0.00763f
C905 B.n412 VSUBS 0.00763f
C906 B.n413 VSUBS 0.00763f
C907 B.n414 VSUBS 0.00763f
C908 B.n415 VSUBS 0.00763f
C909 B.n416 VSUBS 0.00763f
C910 B.n417 VSUBS 0.00763f
C911 B.n418 VSUBS 0.00763f
C912 B.n419 VSUBS 0.00763f
C913 B.n420 VSUBS 0.00763f
C914 B.n421 VSUBS 0.00763f
C915 B.n422 VSUBS 0.00763f
C916 B.n423 VSUBS 0.00763f
C917 B.n424 VSUBS 0.00763f
C918 B.n425 VSUBS 0.00763f
C919 B.n426 VSUBS 0.00763f
C920 B.n427 VSUBS 0.00763f
C921 B.n428 VSUBS 0.00763f
C922 B.n429 VSUBS 0.00763f
C923 B.n430 VSUBS 0.00763f
C924 B.n431 VSUBS 0.00763f
C925 B.n432 VSUBS 0.00763f
C926 B.n433 VSUBS 0.00763f
C927 B.n434 VSUBS 0.00763f
C928 B.n435 VSUBS 0.00763f
C929 B.n436 VSUBS 0.00763f
C930 B.n437 VSUBS 0.00763f
C931 B.n438 VSUBS 0.00763f
C932 B.n439 VSUBS 0.00763f
C933 B.n440 VSUBS 0.00763f
C934 B.n441 VSUBS 0.00763f
C935 B.n442 VSUBS 0.00763f
C936 B.n443 VSUBS 0.00763f
C937 B.n444 VSUBS 0.00763f
C938 B.n445 VSUBS 0.00763f
C939 B.n446 VSUBS 0.00763f
C940 B.n447 VSUBS 0.00763f
C941 B.n448 VSUBS 0.00763f
C942 B.n449 VSUBS 0.00763f
C943 B.n450 VSUBS 0.00763f
C944 B.n451 VSUBS 0.00763f
C945 B.n452 VSUBS 0.00763f
C946 B.n453 VSUBS 0.00763f
C947 B.n454 VSUBS 0.018073f
C948 B.n455 VSUBS 0.018073f
C949 B.n456 VSUBS 0.017384f
C950 B.n457 VSUBS 0.00763f
C951 B.n458 VSUBS 0.00763f
C952 B.n459 VSUBS 0.00763f
C953 B.n460 VSUBS 0.00763f
C954 B.n461 VSUBS 0.00763f
C955 B.n462 VSUBS 0.00763f
C956 B.n463 VSUBS 0.00763f
C957 B.n464 VSUBS 0.00763f
C958 B.n465 VSUBS 0.00763f
C959 B.n466 VSUBS 0.00763f
C960 B.n467 VSUBS 0.00763f
C961 B.n468 VSUBS 0.00763f
C962 B.n469 VSUBS 0.00763f
C963 B.n470 VSUBS 0.00763f
C964 B.n471 VSUBS 0.00763f
C965 B.n472 VSUBS 0.00763f
C966 B.n473 VSUBS 0.00763f
C967 B.n474 VSUBS 0.00763f
C968 B.n475 VSUBS 0.00763f
C969 B.n476 VSUBS 0.00763f
C970 B.n477 VSUBS 0.00763f
C971 B.n478 VSUBS 0.00763f
C972 B.n479 VSUBS 0.00763f
C973 B.n480 VSUBS 0.00763f
C974 B.n481 VSUBS 0.00763f
C975 B.n482 VSUBS 0.00763f
C976 B.n483 VSUBS 0.00763f
C977 B.n484 VSUBS 0.00763f
C978 B.n485 VSUBS 0.00763f
C979 B.n486 VSUBS 0.00763f
C980 B.n487 VSUBS 0.00763f
C981 B.n488 VSUBS 0.00763f
C982 B.n489 VSUBS 0.00763f
C983 B.n490 VSUBS 0.00763f
C984 B.n491 VSUBS 0.017277f
.ends

