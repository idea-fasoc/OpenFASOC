* NGSPICE file created from diff_pair_sample_0692.ext - technology: sky130A

.subckt diff_pair_sample_0692 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=0 ps=0 w=10.77 l=0.45
X1 B.t8 B.t6 B.t7 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=0 ps=0 w=10.77 l=0.45
X2 VTAIL.t15 VP.t0 VDD1.t0 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=1.77705 ps=11.1 w=10.77 l=0.45
X3 VTAIL.t6 VN.t0 VDD2.t7 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=1.77705 ps=11.1 w=10.77 l=0.45
X4 VDD1.t2 VP.t1 VTAIL.t14 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X5 VTAIL.t13 VP.t2 VDD1.t6 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=1.77705 ps=11.1 w=10.77 l=0.45
X6 B.t5 B.t3 B.t4 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=0 ps=0 w=10.77 l=0.45
X7 VTAIL.t12 VP.t3 VDD1.t5 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X8 VDD2.t6 VN.t1 VTAIL.t3 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=4.2003 ps=22.32 w=10.77 l=0.45
X9 VTAIL.t11 VP.t4 VDD1.t4 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X10 VDD1.t1 VP.t5 VTAIL.t10 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=4.2003 ps=22.32 w=10.77 l=0.45
X11 B.t2 B.t0 B.t1 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=0 ps=0 w=10.77 l=0.45
X12 VDD2.t5 VN.t2 VTAIL.t5 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X13 VDD2.t4 VN.t3 VTAIL.t1 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=4.2003 ps=22.32 w=10.77 l=0.45
X14 VDD1.t7 VP.t6 VTAIL.t9 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X15 VTAIL.t2 VN.t4 VDD2.t3 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X16 VDD2.t2 VN.t5 VTAIL.t4 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X17 VTAIL.t7 VN.t6 VDD2.t1 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=1.77705 ps=11.1 w=10.77 l=0.45
X18 VTAIL.t0 VN.t7 VDD2.t0 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=4.2003 pd=22.32 as=1.77705 ps=11.1 w=10.77 l=0.45
X19 VDD1.t3 VP.t7 VTAIL.t8 w_n1750_n3122# sky130_fd_pr__pfet_01v8 ad=1.77705 pd=11.1 as=4.2003 ps=22.32 w=10.77 l=0.45
R0 B.n216 B.t9 784.54
R1 B.n99 B.t0 784.54
R2 B.n39 B.t6 784.54
R3 B.n32 B.t3 784.54
R4 B.n293 B.n292 585
R5 B.n291 B.n80 585
R6 B.n290 B.n289 585
R7 B.n288 B.n81 585
R8 B.n287 B.n286 585
R9 B.n285 B.n82 585
R10 B.n284 B.n283 585
R11 B.n282 B.n83 585
R12 B.n281 B.n280 585
R13 B.n279 B.n84 585
R14 B.n278 B.n277 585
R15 B.n276 B.n85 585
R16 B.n275 B.n274 585
R17 B.n273 B.n86 585
R18 B.n272 B.n271 585
R19 B.n270 B.n87 585
R20 B.n269 B.n268 585
R21 B.n267 B.n88 585
R22 B.n266 B.n265 585
R23 B.n264 B.n89 585
R24 B.n263 B.n262 585
R25 B.n261 B.n90 585
R26 B.n260 B.n259 585
R27 B.n258 B.n91 585
R28 B.n257 B.n256 585
R29 B.n255 B.n92 585
R30 B.n254 B.n253 585
R31 B.n252 B.n93 585
R32 B.n251 B.n250 585
R33 B.n249 B.n94 585
R34 B.n248 B.n247 585
R35 B.n246 B.n95 585
R36 B.n245 B.n244 585
R37 B.n243 B.n96 585
R38 B.n242 B.n241 585
R39 B.n240 B.n97 585
R40 B.n239 B.n238 585
R41 B.n237 B.n98 585
R42 B.n235 B.n234 585
R43 B.n233 B.n101 585
R44 B.n232 B.n231 585
R45 B.n230 B.n102 585
R46 B.n229 B.n228 585
R47 B.n227 B.n103 585
R48 B.n226 B.n225 585
R49 B.n224 B.n104 585
R50 B.n223 B.n222 585
R51 B.n221 B.n105 585
R52 B.n220 B.n219 585
R53 B.n215 B.n106 585
R54 B.n214 B.n213 585
R55 B.n212 B.n107 585
R56 B.n211 B.n210 585
R57 B.n209 B.n108 585
R58 B.n208 B.n207 585
R59 B.n206 B.n109 585
R60 B.n205 B.n204 585
R61 B.n203 B.n110 585
R62 B.n202 B.n201 585
R63 B.n200 B.n111 585
R64 B.n199 B.n198 585
R65 B.n197 B.n112 585
R66 B.n196 B.n195 585
R67 B.n194 B.n113 585
R68 B.n193 B.n192 585
R69 B.n191 B.n114 585
R70 B.n190 B.n189 585
R71 B.n188 B.n115 585
R72 B.n187 B.n186 585
R73 B.n185 B.n116 585
R74 B.n184 B.n183 585
R75 B.n182 B.n117 585
R76 B.n181 B.n180 585
R77 B.n179 B.n118 585
R78 B.n178 B.n177 585
R79 B.n176 B.n119 585
R80 B.n175 B.n174 585
R81 B.n173 B.n120 585
R82 B.n172 B.n171 585
R83 B.n170 B.n121 585
R84 B.n169 B.n168 585
R85 B.n167 B.n122 585
R86 B.n166 B.n165 585
R87 B.n164 B.n123 585
R88 B.n163 B.n162 585
R89 B.n161 B.n124 585
R90 B.n294 B.n79 585
R91 B.n296 B.n295 585
R92 B.n297 B.n78 585
R93 B.n299 B.n298 585
R94 B.n300 B.n77 585
R95 B.n302 B.n301 585
R96 B.n303 B.n76 585
R97 B.n305 B.n304 585
R98 B.n306 B.n75 585
R99 B.n308 B.n307 585
R100 B.n309 B.n74 585
R101 B.n311 B.n310 585
R102 B.n312 B.n73 585
R103 B.n314 B.n313 585
R104 B.n315 B.n72 585
R105 B.n317 B.n316 585
R106 B.n318 B.n71 585
R107 B.n320 B.n319 585
R108 B.n321 B.n70 585
R109 B.n323 B.n322 585
R110 B.n324 B.n69 585
R111 B.n326 B.n325 585
R112 B.n327 B.n68 585
R113 B.n329 B.n328 585
R114 B.n330 B.n67 585
R115 B.n332 B.n331 585
R116 B.n333 B.n66 585
R117 B.n335 B.n334 585
R118 B.n336 B.n65 585
R119 B.n338 B.n337 585
R120 B.n339 B.n64 585
R121 B.n341 B.n340 585
R122 B.n342 B.n63 585
R123 B.n344 B.n343 585
R124 B.n345 B.n62 585
R125 B.n347 B.n346 585
R126 B.n348 B.n61 585
R127 B.n350 B.n349 585
R128 B.n351 B.n60 585
R129 B.n353 B.n352 585
R130 B.n483 B.n482 585
R131 B.n481 B.n12 585
R132 B.n480 B.n479 585
R133 B.n478 B.n13 585
R134 B.n477 B.n476 585
R135 B.n475 B.n14 585
R136 B.n474 B.n473 585
R137 B.n472 B.n15 585
R138 B.n471 B.n470 585
R139 B.n469 B.n16 585
R140 B.n468 B.n467 585
R141 B.n466 B.n17 585
R142 B.n465 B.n464 585
R143 B.n463 B.n18 585
R144 B.n462 B.n461 585
R145 B.n460 B.n19 585
R146 B.n459 B.n458 585
R147 B.n457 B.n20 585
R148 B.n456 B.n455 585
R149 B.n454 B.n21 585
R150 B.n453 B.n452 585
R151 B.n451 B.n22 585
R152 B.n450 B.n449 585
R153 B.n448 B.n23 585
R154 B.n447 B.n446 585
R155 B.n445 B.n24 585
R156 B.n444 B.n443 585
R157 B.n442 B.n25 585
R158 B.n441 B.n440 585
R159 B.n439 B.n26 585
R160 B.n438 B.n437 585
R161 B.n436 B.n27 585
R162 B.n435 B.n434 585
R163 B.n433 B.n28 585
R164 B.n432 B.n431 585
R165 B.n430 B.n29 585
R166 B.n429 B.n428 585
R167 B.n427 B.n30 585
R168 B.n426 B.n425 585
R169 B.n424 B.n31 585
R170 B.n423 B.n422 585
R171 B.n421 B.n35 585
R172 B.n420 B.n419 585
R173 B.n418 B.n36 585
R174 B.n417 B.n416 585
R175 B.n415 B.n37 585
R176 B.n414 B.n413 585
R177 B.n412 B.n38 585
R178 B.n410 B.n409 585
R179 B.n408 B.n41 585
R180 B.n407 B.n406 585
R181 B.n405 B.n42 585
R182 B.n404 B.n403 585
R183 B.n402 B.n43 585
R184 B.n401 B.n400 585
R185 B.n399 B.n44 585
R186 B.n398 B.n397 585
R187 B.n396 B.n45 585
R188 B.n395 B.n394 585
R189 B.n393 B.n46 585
R190 B.n392 B.n391 585
R191 B.n390 B.n47 585
R192 B.n389 B.n388 585
R193 B.n387 B.n48 585
R194 B.n386 B.n385 585
R195 B.n384 B.n49 585
R196 B.n383 B.n382 585
R197 B.n381 B.n50 585
R198 B.n380 B.n379 585
R199 B.n378 B.n51 585
R200 B.n377 B.n376 585
R201 B.n375 B.n52 585
R202 B.n374 B.n373 585
R203 B.n372 B.n53 585
R204 B.n371 B.n370 585
R205 B.n369 B.n54 585
R206 B.n368 B.n367 585
R207 B.n366 B.n55 585
R208 B.n365 B.n364 585
R209 B.n363 B.n56 585
R210 B.n362 B.n361 585
R211 B.n360 B.n57 585
R212 B.n359 B.n358 585
R213 B.n357 B.n58 585
R214 B.n356 B.n355 585
R215 B.n354 B.n59 585
R216 B.n484 B.n11 585
R217 B.n486 B.n485 585
R218 B.n487 B.n10 585
R219 B.n489 B.n488 585
R220 B.n490 B.n9 585
R221 B.n492 B.n491 585
R222 B.n493 B.n8 585
R223 B.n495 B.n494 585
R224 B.n496 B.n7 585
R225 B.n498 B.n497 585
R226 B.n499 B.n6 585
R227 B.n501 B.n500 585
R228 B.n502 B.n5 585
R229 B.n504 B.n503 585
R230 B.n505 B.n4 585
R231 B.n507 B.n506 585
R232 B.n508 B.n3 585
R233 B.n510 B.n509 585
R234 B.n511 B.n0 585
R235 B.n2 B.n1 585
R236 B.n134 B.n133 585
R237 B.n136 B.n135 585
R238 B.n137 B.n132 585
R239 B.n139 B.n138 585
R240 B.n140 B.n131 585
R241 B.n142 B.n141 585
R242 B.n143 B.n130 585
R243 B.n145 B.n144 585
R244 B.n146 B.n129 585
R245 B.n148 B.n147 585
R246 B.n149 B.n128 585
R247 B.n151 B.n150 585
R248 B.n152 B.n127 585
R249 B.n154 B.n153 585
R250 B.n155 B.n126 585
R251 B.n157 B.n156 585
R252 B.n158 B.n125 585
R253 B.n160 B.n159 585
R254 B.n159 B.n124 478.086
R255 B.n294 B.n293 478.086
R256 B.n354 B.n353 478.086
R257 B.n482 B.n11 478.086
R258 B.n99 B.t1 368.69
R259 B.n39 B.t8 368.69
R260 B.n216 B.t10 368.69
R261 B.n32 B.t5 368.69
R262 B.n100 B.t2 353.562
R263 B.n40 B.t7 353.562
R264 B.n217 B.t11 353.562
R265 B.n33 B.t4 353.562
R266 B.n513 B.n512 256.663
R267 B.n512 B.n511 235.042
R268 B.n512 B.n2 235.042
R269 B.n163 B.n124 163.367
R270 B.n164 B.n163 163.367
R271 B.n165 B.n164 163.367
R272 B.n165 B.n122 163.367
R273 B.n169 B.n122 163.367
R274 B.n170 B.n169 163.367
R275 B.n171 B.n170 163.367
R276 B.n171 B.n120 163.367
R277 B.n175 B.n120 163.367
R278 B.n176 B.n175 163.367
R279 B.n177 B.n176 163.367
R280 B.n177 B.n118 163.367
R281 B.n181 B.n118 163.367
R282 B.n182 B.n181 163.367
R283 B.n183 B.n182 163.367
R284 B.n183 B.n116 163.367
R285 B.n187 B.n116 163.367
R286 B.n188 B.n187 163.367
R287 B.n189 B.n188 163.367
R288 B.n189 B.n114 163.367
R289 B.n193 B.n114 163.367
R290 B.n194 B.n193 163.367
R291 B.n195 B.n194 163.367
R292 B.n195 B.n112 163.367
R293 B.n199 B.n112 163.367
R294 B.n200 B.n199 163.367
R295 B.n201 B.n200 163.367
R296 B.n201 B.n110 163.367
R297 B.n205 B.n110 163.367
R298 B.n206 B.n205 163.367
R299 B.n207 B.n206 163.367
R300 B.n207 B.n108 163.367
R301 B.n211 B.n108 163.367
R302 B.n212 B.n211 163.367
R303 B.n213 B.n212 163.367
R304 B.n213 B.n106 163.367
R305 B.n220 B.n106 163.367
R306 B.n221 B.n220 163.367
R307 B.n222 B.n221 163.367
R308 B.n222 B.n104 163.367
R309 B.n226 B.n104 163.367
R310 B.n227 B.n226 163.367
R311 B.n228 B.n227 163.367
R312 B.n228 B.n102 163.367
R313 B.n232 B.n102 163.367
R314 B.n233 B.n232 163.367
R315 B.n234 B.n233 163.367
R316 B.n234 B.n98 163.367
R317 B.n239 B.n98 163.367
R318 B.n240 B.n239 163.367
R319 B.n241 B.n240 163.367
R320 B.n241 B.n96 163.367
R321 B.n245 B.n96 163.367
R322 B.n246 B.n245 163.367
R323 B.n247 B.n246 163.367
R324 B.n247 B.n94 163.367
R325 B.n251 B.n94 163.367
R326 B.n252 B.n251 163.367
R327 B.n253 B.n252 163.367
R328 B.n253 B.n92 163.367
R329 B.n257 B.n92 163.367
R330 B.n258 B.n257 163.367
R331 B.n259 B.n258 163.367
R332 B.n259 B.n90 163.367
R333 B.n263 B.n90 163.367
R334 B.n264 B.n263 163.367
R335 B.n265 B.n264 163.367
R336 B.n265 B.n88 163.367
R337 B.n269 B.n88 163.367
R338 B.n270 B.n269 163.367
R339 B.n271 B.n270 163.367
R340 B.n271 B.n86 163.367
R341 B.n275 B.n86 163.367
R342 B.n276 B.n275 163.367
R343 B.n277 B.n276 163.367
R344 B.n277 B.n84 163.367
R345 B.n281 B.n84 163.367
R346 B.n282 B.n281 163.367
R347 B.n283 B.n282 163.367
R348 B.n283 B.n82 163.367
R349 B.n287 B.n82 163.367
R350 B.n288 B.n287 163.367
R351 B.n289 B.n288 163.367
R352 B.n289 B.n80 163.367
R353 B.n293 B.n80 163.367
R354 B.n353 B.n60 163.367
R355 B.n349 B.n60 163.367
R356 B.n349 B.n348 163.367
R357 B.n348 B.n347 163.367
R358 B.n347 B.n62 163.367
R359 B.n343 B.n62 163.367
R360 B.n343 B.n342 163.367
R361 B.n342 B.n341 163.367
R362 B.n341 B.n64 163.367
R363 B.n337 B.n64 163.367
R364 B.n337 B.n336 163.367
R365 B.n336 B.n335 163.367
R366 B.n335 B.n66 163.367
R367 B.n331 B.n66 163.367
R368 B.n331 B.n330 163.367
R369 B.n330 B.n329 163.367
R370 B.n329 B.n68 163.367
R371 B.n325 B.n68 163.367
R372 B.n325 B.n324 163.367
R373 B.n324 B.n323 163.367
R374 B.n323 B.n70 163.367
R375 B.n319 B.n70 163.367
R376 B.n319 B.n318 163.367
R377 B.n318 B.n317 163.367
R378 B.n317 B.n72 163.367
R379 B.n313 B.n72 163.367
R380 B.n313 B.n312 163.367
R381 B.n312 B.n311 163.367
R382 B.n311 B.n74 163.367
R383 B.n307 B.n74 163.367
R384 B.n307 B.n306 163.367
R385 B.n306 B.n305 163.367
R386 B.n305 B.n76 163.367
R387 B.n301 B.n76 163.367
R388 B.n301 B.n300 163.367
R389 B.n300 B.n299 163.367
R390 B.n299 B.n78 163.367
R391 B.n295 B.n78 163.367
R392 B.n295 B.n294 163.367
R393 B.n482 B.n481 163.367
R394 B.n481 B.n480 163.367
R395 B.n480 B.n13 163.367
R396 B.n476 B.n13 163.367
R397 B.n476 B.n475 163.367
R398 B.n475 B.n474 163.367
R399 B.n474 B.n15 163.367
R400 B.n470 B.n15 163.367
R401 B.n470 B.n469 163.367
R402 B.n469 B.n468 163.367
R403 B.n468 B.n17 163.367
R404 B.n464 B.n17 163.367
R405 B.n464 B.n463 163.367
R406 B.n463 B.n462 163.367
R407 B.n462 B.n19 163.367
R408 B.n458 B.n19 163.367
R409 B.n458 B.n457 163.367
R410 B.n457 B.n456 163.367
R411 B.n456 B.n21 163.367
R412 B.n452 B.n21 163.367
R413 B.n452 B.n451 163.367
R414 B.n451 B.n450 163.367
R415 B.n450 B.n23 163.367
R416 B.n446 B.n23 163.367
R417 B.n446 B.n445 163.367
R418 B.n445 B.n444 163.367
R419 B.n444 B.n25 163.367
R420 B.n440 B.n25 163.367
R421 B.n440 B.n439 163.367
R422 B.n439 B.n438 163.367
R423 B.n438 B.n27 163.367
R424 B.n434 B.n27 163.367
R425 B.n434 B.n433 163.367
R426 B.n433 B.n432 163.367
R427 B.n432 B.n29 163.367
R428 B.n428 B.n29 163.367
R429 B.n428 B.n427 163.367
R430 B.n427 B.n426 163.367
R431 B.n426 B.n31 163.367
R432 B.n422 B.n31 163.367
R433 B.n422 B.n421 163.367
R434 B.n421 B.n420 163.367
R435 B.n420 B.n36 163.367
R436 B.n416 B.n36 163.367
R437 B.n416 B.n415 163.367
R438 B.n415 B.n414 163.367
R439 B.n414 B.n38 163.367
R440 B.n409 B.n38 163.367
R441 B.n409 B.n408 163.367
R442 B.n408 B.n407 163.367
R443 B.n407 B.n42 163.367
R444 B.n403 B.n42 163.367
R445 B.n403 B.n402 163.367
R446 B.n402 B.n401 163.367
R447 B.n401 B.n44 163.367
R448 B.n397 B.n44 163.367
R449 B.n397 B.n396 163.367
R450 B.n396 B.n395 163.367
R451 B.n395 B.n46 163.367
R452 B.n391 B.n46 163.367
R453 B.n391 B.n390 163.367
R454 B.n390 B.n389 163.367
R455 B.n389 B.n48 163.367
R456 B.n385 B.n48 163.367
R457 B.n385 B.n384 163.367
R458 B.n384 B.n383 163.367
R459 B.n383 B.n50 163.367
R460 B.n379 B.n50 163.367
R461 B.n379 B.n378 163.367
R462 B.n378 B.n377 163.367
R463 B.n377 B.n52 163.367
R464 B.n373 B.n52 163.367
R465 B.n373 B.n372 163.367
R466 B.n372 B.n371 163.367
R467 B.n371 B.n54 163.367
R468 B.n367 B.n54 163.367
R469 B.n367 B.n366 163.367
R470 B.n366 B.n365 163.367
R471 B.n365 B.n56 163.367
R472 B.n361 B.n56 163.367
R473 B.n361 B.n360 163.367
R474 B.n360 B.n359 163.367
R475 B.n359 B.n58 163.367
R476 B.n355 B.n58 163.367
R477 B.n355 B.n354 163.367
R478 B.n486 B.n11 163.367
R479 B.n487 B.n486 163.367
R480 B.n488 B.n487 163.367
R481 B.n488 B.n9 163.367
R482 B.n492 B.n9 163.367
R483 B.n493 B.n492 163.367
R484 B.n494 B.n493 163.367
R485 B.n494 B.n7 163.367
R486 B.n498 B.n7 163.367
R487 B.n499 B.n498 163.367
R488 B.n500 B.n499 163.367
R489 B.n500 B.n5 163.367
R490 B.n504 B.n5 163.367
R491 B.n505 B.n504 163.367
R492 B.n506 B.n505 163.367
R493 B.n506 B.n3 163.367
R494 B.n510 B.n3 163.367
R495 B.n511 B.n510 163.367
R496 B.n134 B.n2 163.367
R497 B.n135 B.n134 163.367
R498 B.n135 B.n132 163.367
R499 B.n139 B.n132 163.367
R500 B.n140 B.n139 163.367
R501 B.n141 B.n140 163.367
R502 B.n141 B.n130 163.367
R503 B.n145 B.n130 163.367
R504 B.n146 B.n145 163.367
R505 B.n147 B.n146 163.367
R506 B.n147 B.n128 163.367
R507 B.n151 B.n128 163.367
R508 B.n152 B.n151 163.367
R509 B.n153 B.n152 163.367
R510 B.n153 B.n126 163.367
R511 B.n157 B.n126 163.367
R512 B.n158 B.n157 163.367
R513 B.n159 B.n158 163.367
R514 B.n218 B.n217 59.5399
R515 B.n236 B.n100 59.5399
R516 B.n411 B.n40 59.5399
R517 B.n34 B.n33 59.5399
R518 B.n484 B.n483 31.0639
R519 B.n352 B.n59 31.0639
R520 B.n292 B.n79 31.0639
R521 B.n161 B.n160 31.0639
R522 B B.n513 18.0485
R523 B.n217 B.n216 15.1278
R524 B.n100 B.n99 15.1278
R525 B.n40 B.n39 15.1278
R526 B.n33 B.n32 15.1278
R527 B.n485 B.n484 10.6151
R528 B.n485 B.n10 10.6151
R529 B.n489 B.n10 10.6151
R530 B.n490 B.n489 10.6151
R531 B.n491 B.n490 10.6151
R532 B.n491 B.n8 10.6151
R533 B.n495 B.n8 10.6151
R534 B.n496 B.n495 10.6151
R535 B.n497 B.n496 10.6151
R536 B.n497 B.n6 10.6151
R537 B.n501 B.n6 10.6151
R538 B.n502 B.n501 10.6151
R539 B.n503 B.n502 10.6151
R540 B.n503 B.n4 10.6151
R541 B.n507 B.n4 10.6151
R542 B.n508 B.n507 10.6151
R543 B.n509 B.n508 10.6151
R544 B.n509 B.n0 10.6151
R545 B.n483 B.n12 10.6151
R546 B.n479 B.n12 10.6151
R547 B.n479 B.n478 10.6151
R548 B.n478 B.n477 10.6151
R549 B.n477 B.n14 10.6151
R550 B.n473 B.n14 10.6151
R551 B.n473 B.n472 10.6151
R552 B.n472 B.n471 10.6151
R553 B.n471 B.n16 10.6151
R554 B.n467 B.n16 10.6151
R555 B.n467 B.n466 10.6151
R556 B.n466 B.n465 10.6151
R557 B.n465 B.n18 10.6151
R558 B.n461 B.n18 10.6151
R559 B.n461 B.n460 10.6151
R560 B.n460 B.n459 10.6151
R561 B.n459 B.n20 10.6151
R562 B.n455 B.n20 10.6151
R563 B.n455 B.n454 10.6151
R564 B.n454 B.n453 10.6151
R565 B.n453 B.n22 10.6151
R566 B.n449 B.n22 10.6151
R567 B.n449 B.n448 10.6151
R568 B.n448 B.n447 10.6151
R569 B.n447 B.n24 10.6151
R570 B.n443 B.n24 10.6151
R571 B.n443 B.n442 10.6151
R572 B.n442 B.n441 10.6151
R573 B.n441 B.n26 10.6151
R574 B.n437 B.n26 10.6151
R575 B.n437 B.n436 10.6151
R576 B.n436 B.n435 10.6151
R577 B.n435 B.n28 10.6151
R578 B.n431 B.n28 10.6151
R579 B.n431 B.n430 10.6151
R580 B.n430 B.n429 10.6151
R581 B.n429 B.n30 10.6151
R582 B.n425 B.n424 10.6151
R583 B.n424 B.n423 10.6151
R584 B.n423 B.n35 10.6151
R585 B.n419 B.n35 10.6151
R586 B.n419 B.n418 10.6151
R587 B.n418 B.n417 10.6151
R588 B.n417 B.n37 10.6151
R589 B.n413 B.n37 10.6151
R590 B.n413 B.n412 10.6151
R591 B.n410 B.n41 10.6151
R592 B.n406 B.n41 10.6151
R593 B.n406 B.n405 10.6151
R594 B.n405 B.n404 10.6151
R595 B.n404 B.n43 10.6151
R596 B.n400 B.n43 10.6151
R597 B.n400 B.n399 10.6151
R598 B.n399 B.n398 10.6151
R599 B.n398 B.n45 10.6151
R600 B.n394 B.n45 10.6151
R601 B.n394 B.n393 10.6151
R602 B.n393 B.n392 10.6151
R603 B.n392 B.n47 10.6151
R604 B.n388 B.n47 10.6151
R605 B.n388 B.n387 10.6151
R606 B.n387 B.n386 10.6151
R607 B.n386 B.n49 10.6151
R608 B.n382 B.n49 10.6151
R609 B.n382 B.n381 10.6151
R610 B.n381 B.n380 10.6151
R611 B.n380 B.n51 10.6151
R612 B.n376 B.n51 10.6151
R613 B.n376 B.n375 10.6151
R614 B.n375 B.n374 10.6151
R615 B.n374 B.n53 10.6151
R616 B.n370 B.n53 10.6151
R617 B.n370 B.n369 10.6151
R618 B.n369 B.n368 10.6151
R619 B.n368 B.n55 10.6151
R620 B.n364 B.n55 10.6151
R621 B.n364 B.n363 10.6151
R622 B.n363 B.n362 10.6151
R623 B.n362 B.n57 10.6151
R624 B.n358 B.n57 10.6151
R625 B.n358 B.n357 10.6151
R626 B.n357 B.n356 10.6151
R627 B.n356 B.n59 10.6151
R628 B.n352 B.n351 10.6151
R629 B.n351 B.n350 10.6151
R630 B.n350 B.n61 10.6151
R631 B.n346 B.n61 10.6151
R632 B.n346 B.n345 10.6151
R633 B.n345 B.n344 10.6151
R634 B.n344 B.n63 10.6151
R635 B.n340 B.n63 10.6151
R636 B.n340 B.n339 10.6151
R637 B.n339 B.n338 10.6151
R638 B.n338 B.n65 10.6151
R639 B.n334 B.n65 10.6151
R640 B.n334 B.n333 10.6151
R641 B.n333 B.n332 10.6151
R642 B.n332 B.n67 10.6151
R643 B.n328 B.n67 10.6151
R644 B.n328 B.n327 10.6151
R645 B.n327 B.n326 10.6151
R646 B.n326 B.n69 10.6151
R647 B.n322 B.n69 10.6151
R648 B.n322 B.n321 10.6151
R649 B.n321 B.n320 10.6151
R650 B.n320 B.n71 10.6151
R651 B.n316 B.n71 10.6151
R652 B.n316 B.n315 10.6151
R653 B.n315 B.n314 10.6151
R654 B.n314 B.n73 10.6151
R655 B.n310 B.n73 10.6151
R656 B.n310 B.n309 10.6151
R657 B.n309 B.n308 10.6151
R658 B.n308 B.n75 10.6151
R659 B.n304 B.n75 10.6151
R660 B.n304 B.n303 10.6151
R661 B.n303 B.n302 10.6151
R662 B.n302 B.n77 10.6151
R663 B.n298 B.n77 10.6151
R664 B.n298 B.n297 10.6151
R665 B.n297 B.n296 10.6151
R666 B.n296 B.n79 10.6151
R667 B.n133 B.n1 10.6151
R668 B.n136 B.n133 10.6151
R669 B.n137 B.n136 10.6151
R670 B.n138 B.n137 10.6151
R671 B.n138 B.n131 10.6151
R672 B.n142 B.n131 10.6151
R673 B.n143 B.n142 10.6151
R674 B.n144 B.n143 10.6151
R675 B.n144 B.n129 10.6151
R676 B.n148 B.n129 10.6151
R677 B.n149 B.n148 10.6151
R678 B.n150 B.n149 10.6151
R679 B.n150 B.n127 10.6151
R680 B.n154 B.n127 10.6151
R681 B.n155 B.n154 10.6151
R682 B.n156 B.n155 10.6151
R683 B.n156 B.n125 10.6151
R684 B.n160 B.n125 10.6151
R685 B.n162 B.n161 10.6151
R686 B.n162 B.n123 10.6151
R687 B.n166 B.n123 10.6151
R688 B.n167 B.n166 10.6151
R689 B.n168 B.n167 10.6151
R690 B.n168 B.n121 10.6151
R691 B.n172 B.n121 10.6151
R692 B.n173 B.n172 10.6151
R693 B.n174 B.n173 10.6151
R694 B.n174 B.n119 10.6151
R695 B.n178 B.n119 10.6151
R696 B.n179 B.n178 10.6151
R697 B.n180 B.n179 10.6151
R698 B.n180 B.n117 10.6151
R699 B.n184 B.n117 10.6151
R700 B.n185 B.n184 10.6151
R701 B.n186 B.n185 10.6151
R702 B.n186 B.n115 10.6151
R703 B.n190 B.n115 10.6151
R704 B.n191 B.n190 10.6151
R705 B.n192 B.n191 10.6151
R706 B.n192 B.n113 10.6151
R707 B.n196 B.n113 10.6151
R708 B.n197 B.n196 10.6151
R709 B.n198 B.n197 10.6151
R710 B.n198 B.n111 10.6151
R711 B.n202 B.n111 10.6151
R712 B.n203 B.n202 10.6151
R713 B.n204 B.n203 10.6151
R714 B.n204 B.n109 10.6151
R715 B.n208 B.n109 10.6151
R716 B.n209 B.n208 10.6151
R717 B.n210 B.n209 10.6151
R718 B.n210 B.n107 10.6151
R719 B.n214 B.n107 10.6151
R720 B.n215 B.n214 10.6151
R721 B.n219 B.n215 10.6151
R722 B.n223 B.n105 10.6151
R723 B.n224 B.n223 10.6151
R724 B.n225 B.n224 10.6151
R725 B.n225 B.n103 10.6151
R726 B.n229 B.n103 10.6151
R727 B.n230 B.n229 10.6151
R728 B.n231 B.n230 10.6151
R729 B.n231 B.n101 10.6151
R730 B.n235 B.n101 10.6151
R731 B.n238 B.n237 10.6151
R732 B.n238 B.n97 10.6151
R733 B.n242 B.n97 10.6151
R734 B.n243 B.n242 10.6151
R735 B.n244 B.n243 10.6151
R736 B.n244 B.n95 10.6151
R737 B.n248 B.n95 10.6151
R738 B.n249 B.n248 10.6151
R739 B.n250 B.n249 10.6151
R740 B.n250 B.n93 10.6151
R741 B.n254 B.n93 10.6151
R742 B.n255 B.n254 10.6151
R743 B.n256 B.n255 10.6151
R744 B.n256 B.n91 10.6151
R745 B.n260 B.n91 10.6151
R746 B.n261 B.n260 10.6151
R747 B.n262 B.n261 10.6151
R748 B.n262 B.n89 10.6151
R749 B.n266 B.n89 10.6151
R750 B.n267 B.n266 10.6151
R751 B.n268 B.n267 10.6151
R752 B.n268 B.n87 10.6151
R753 B.n272 B.n87 10.6151
R754 B.n273 B.n272 10.6151
R755 B.n274 B.n273 10.6151
R756 B.n274 B.n85 10.6151
R757 B.n278 B.n85 10.6151
R758 B.n279 B.n278 10.6151
R759 B.n280 B.n279 10.6151
R760 B.n280 B.n83 10.6151
R761 B.n284 B.n83 10.6151
R762 B.n285 B.n284 10.6151
R763 B.n286 B.n285 10.6151
R764 B.n286 B.n81 10.6151
R765 B.n290 B.n81 10.6151
R766 B.n291 B.n290 10.6151
R767 B.n292 B.n291 10.6151
R768 B.n34 B.n30 9.36635
R769 B.n411 B.n410 9.36635
R770 B.n219 B.n218 9.36635
R771 B.n237 B.n236 9.36635
R772 B.n513 B.n0 8.11757
R773 B.n513 B.n1 8.11757
R774 B.n425 B.n34 1.24928
R775 B.n412 B.n411 1.24928
R776 B.n218 B.n105 1.24928
R777 B.n236 B.n235 1.24928
R778 VP.n4 VP.t0 685.606
R779 VP.n10 VP.t2 664.625
R780 VP.n1 VP.t1 664.625
R781 VP.n15 VP.t3 664.625
R782 VP.n16 VP.t5 664.625
R783 VP.n8 VP.t7 664.625
R784 VP.n7 VP.t4 664.625
R785 VP.n3 VP.t6 664.625
R786 VP.n17 VP.n16 161.3
R787 VP.n6 VP.n5 161.3
R788 VP.n7 VP.n2 161.3
R789 VP.n9 VP.n8 161.3
R790 VP.n15 VP.n0 161.3
R791 VP.n14 VP.n13 161.3
R792 VP.n12 VP.n1 161.3
R793 VP.n11 VP.n10 161.3
R794 VP.n5 VP.n4 70.4033
R795 VP.n10 VP.n1 48.2005
R796 VP.n16 VP.n15 48.2005
R797 VP.n8 VP.n7 48.2005
R798 VP.n11 VP.n9 39.9247
R799 VP.n14 VP.n1 24.1005
R800 VP.n15 VP.n14 24.1005
R801 VP.n6 VP.n3 24.1005
R802 VP.n7 VP.n6 24.1005
R803 VP.n4 VP.n3 20.9576
R804 VP.n5 VP.n2 0.189894
R805 VP.n9 VP.n2 0.189894
R806 VP.n12 VP.n11 0.189894
R807 VP.n13 VP.n12 0.189894
R808 VP.n13 VP.n0 0.189894
R809 VP.n17 VP.n0 0.189894
R810 VP VP.n17 0.0516364
R811 VDD1 VDD1.n0 78.006
R812 VDD1.n3 VDD1.n2 77.8923
R813 VDD1.n3 VDD1.n1 77.8923
R814 VDD1.n5 VDD1.n4 77.6114
R815 VDD1.n5 VDD1.n3 36.6086
R816 VDD1.n4 VDD1.t4 3.01861
R817 VDD1.n4 VDD1.t3 3.01861
R818 VDD1.n0 VDD1.t0 3.01861
R819 VDD1.n0 VDD1.t7 3.01861
R820 VDD1.n2 VDD1.t5 3.01861
R821 VDD1.n2 VDD1.t1 3.01861
R822 VDD1.n1 VDD1.t6 3.01861
R823 VDD1.n1 VDD1.t2 3.01861
R824 VDD1 VDD1.n5 0.278517
R825 VTAIL.n466 VTAIL.n414 756.745
R826 VTAIL.n54 VTAIL.n2 756.745
R827 VTAIL.n112 VTAIL.n60 756.745
R828 VTAIL.n172 VTAIL.n120 756.745
R829 VTAIL.n408 VTAIL.n356 756.745
R830 VTAIL.n348 VTAIL.n296 756.745
R831 VTAIL.n290 VTAIL.n238 756.745
R832 VTAIL.n230 VTAIL.n178 756.745
R833 VTAIL.n433 VTAIL.n432 585
R834 VTAIL.n430 VTAIL.n429 585
R835 VTAIL.n439 VTAIL.n438 585
R836 VTAIL.n441 VTAIL.n440 585
R837 VTAIL.n426 VTAIL.n425 585
R838 VTAIL.n447 VTAIL.n446 585
R839 VTAIL.n450 VTAIL.n449 585
R840 VTAIL.n448 VTAIL.n422 585
R841 VTAIL.n455 VTAIL.n421 585
R842 VTAIL.n457 VTAIL.n456 585
R843 VTAIL.n459 VTAIL.n458 585
R844 VTAIL.n418 VTAIL.n417 585
R845 VTAIL.n465 VTAIL.n464 585
R846 VTAIL.n467 VTAIL.n466 585
R847 VTAIL.n21 VTAIL.n20 585
R848 VTAIL.n18 VTAIL.n17 585
R849 VTAIL.n27 VTAIL.n26 585
R850 VTAIL.n29 VTAIL.n28 585
R851 VTAIL.n14 VTAIL.n13 585
R852 VTAIL.n35 VTAIL.n34 585
R853 VTAIL.n38 VTAIL.n37 585
R854 VTAIL.n36 VTAIL.n10 585
R855 VTAIL.n43 VTAIL.n9 585
R856 VTAIL.n45 VTAIL.n44 585
R857 VTAIL.n47 VTAIL.n46 585
R858 VTAIL.n6 VTAIL.n5 585
R859 VTAIL.n53 VTAIL.n52 585
R860 VTAIL.n55 VTAIL.n54 585
R861 VTAIL.n79 VTAIL.n78 585
R862 VTAIL.n76 VTAIL.n75 585
R863 VTAIL.n85 VTAIL.n84 585
R864 VTAIL.n87 VTAIL.n86 585
R865 VTAIL.n72 VTAIL.n71 585
R866 VTAIL.n93 VTAIL.n92 585
R867 VTAIL.n96 VTAIL.n95 585
R868 VTAIL.n94 VTAIL.n68 585
R869 VTAIL.n101 VTAIL.n67 585
R870 VTAIL.n103 VTAIL.n102 585
R871 VTAIL.n105 VTAIL.n104 585
R872 VTAIL.n64 VTAIL.n63 585
R873 VTAIL.n111 VTAIL.n110 585
R874 VTAIL.n113 VTAIL.n112 585
R875 VTAIL.n139 VTAIL.n138 585
R876 VTAIL.n136 VTAIL.n135 585
R877 VTAIL.n145 VTAIL.n144 585
R878 VTAIL.n147 VTAIL.n146 585
R879 VTAIL.n132 VTAIL.n131 585
R880 VTAIL.n153 VTAIL.n152 585
R881 VTAIL.n156 VTAIL.n155 585
R882 VTAIL.n154 VTAIL.n128 585
R883 VTAIL.n161 VTAIL.n127 585
R884 VTAIL.n163 VTAIL.n162 585
R885 VTAIL.n165 VTAIL.n164 585
R886 VTAIL.n124 VTAIL.n123 585
R887 VTAIL.n171 VTAIL.n170 585
R888 VTAIL.n173 VTAIL.n172 585
R889 VTAIL.n409 VTAIL.n408 585
R890 VTAIL.n407 VTAIL.n406 585
R891 VTAIL.n360 VTAIL.n359 585
R892 VTAIL.n401 VTAIL.n400 585
R893 VTAIL.n399 VTAIL.n398 585
R894 VTAIL.n397 VTAIL.n363 585
R895 VTAIL.n367 VTAIL.n364 585
R896 VTAIL.n392 VTAIL.n391 585
R897 VTAIL.n390 VTAIL.n389 585
R898 VTAIL.n369 VTAIL.n368 585
R899 VTAIL.n384 VTAIL.n383 585
R900 VTAIL.n382 VTAIL.n381 585
R901 VTAIL.n373 VTAIL.n372 585
R902 VTAIL.n376 VTAIL.n375 585
R903 VTAIL.n349 VTAIL.n348 585
R904 VTAIL.n347 VTAIL.n346 585
R905 VTAIL.n300 VTAIL.n299 585
R906 VTAIL.n341 VTAIL.n340 585
R907 VTAIL.n339 VTAIL.n338 585
R908 VTAIL.n337 VTAIL.n303 585
R909 VTAIL.n307 VTAIL.n304 585
R910 VTAIL.n332 VTAIL.n331 585
R911 VTAIL.n330 VTAIL.n329 585
R912 VTAIL.n309 VTAIL.n308 585
R913 VTAIL.n324 VTAIL.n323 585
R914 VTAIL.n322 VTAIL.n321 585
R915 VTAIL.n313 VTAIL.n312 585
R916 VTAIL.n316 VTAIL.n315 585
R917 VTAIL.n291 VTAIL.n290 585
R918 VTAIL.n289 VTAIL.n288 585
R919 VTAIL.n242 VTAIL.n241 585
R920 VTAIL.n283 VTAIL.n282 585
R921 VTAIL.n281 VTAIL.n280 585
R922 VTAIL.n279 VTAIL.n245 585
R923 VTAIL.n249 VTAIL.n246 585
R924 VTAIL.n274 VTAIL.n273 585
R925 VTAIL.n272 VTAIL.n271 585
R926 VTAIL.n251 VTAIL.n250 585
R927 VTAIL.n266 VTAIL.n265 585
R928 VTAIL.n264 VTAIL.n263 585
R929 VTAIL.n255 VTAIL.n254 585
R930 VTAIL.n258 VTAIL.n257 585
R931 VTAIL.n231 VTAIL.n230 585
R932 VTAIL.n229 VTAIL.n228 585
R933 VTAIL.n182 VTAIL.n181 585
R934 VTAIL.n223 VTAIL.n222 585
R935 VTAIL.n221 VTAIL.n220 585
R936 VTAIL.n219 VTAIL.n185 585
R937 VTAIL.n189 VTAIL.n186 585
R938 VTAIL.n214 VTAIL.n213 585
R939 VTAIL.n212 VTAIL.n211 585
R940 VTAIL.n191 VTAIL.n190 585
R941 VTAIL.n206 VTAIL.n205 585
R942 VTAIL.n204 VTAIL.n203 585
R943 VTAIL.n195 VTAIL.n194 585
R944 VTAIL.n198 VTAIL.n197 585
R945 VTAIL.t8 VTAIL.n374 329.038
R946 VTAIL.t15 VTAIL.n314 329.038
R947 VTAIL.t3 VTAIL.n256 329.038
R948 VTAIL.t6 VTAIL.n196 329.038
R949 VTAIL.t1 VTAIL.n431 329.038
R950 VTAIL.t0 VTAIL.n19 329.038
R951 VTAIL.t10 VTAIL.n77 329.038
R952 VTAIL.t13 VTAIL.n137 329.038
R953 VTAIL.n432 VTAIL.n429 171.744
R954 VTAIL.n439 VTAIL.n429 171.744
R955 VTAIL.n440 VTAIL.n439 171.744
R956 VTAIL.n440 VTAIL.n425 171.744
R957 VTAIL.n447 VTAIL.n425 171.744
R958 VTAIL.n449 VTAIL.n447 171.744
R959 VTAIL.n449 VTAIL.n448 171.744
R960 VTAIL.n448 VTAIL.n421 171.744
R961 VTAIL.n457 VTAIL.n421 171.744
R962 VTAIL.n458 VTAIL.n457 171.744
R963 VTAIL.n458 VTAIL.n417 171.744
R964 VTAIL.n465 VTAIL.n417 171.744
R965 VTAIL.n466 VTAIL.n465 171.744
R966 VTAIL.n20 VTAIL.n17 171.744
R967 VTAIL.n27 VTAIL.n17 171.744
R968 VTAIL.n28 VTAIL.n27 171.744
R969 VTAIL.n28 VTAIL.n13 171.744
R970 VTAIL.n35 VTAIL.n13 171.744
R971 VTAIL.n37 VTAIL.n35 171.744
R972 VTAIL.n37 VTAIL.n36 171.744
R973 VTAIL.n36 VTAIL.n9 171.744
R974 VTAIL.n45 VTAIL.n9 171.744
R975 VTAIL.n46 VTAIL.n45 171.744
R976 VTAIL.n46 VTAIL.n5 171.744
R977 VTAIL.n53 VTAIL.n5 171.744
R978 VTAIL.n54 VTAIL.n53 171.744
R979 VTAIL.n78 VTAIL.n75 171.744
R980 VTAIL.n85 VTAIL.n75 171.744
R981 VTAIL.n86 VTAIL.n85 171.744
R982 VTAIL.n86 VTAIL.n71 171.744
R983 VTAIL.n93 VTAIL.n71 171.744
R984 VTAIL.n95 VTAIL.n93 171.744
R985 VTAIL.n95 VTAIL.n94 171.744
R986 VTAIL.n94 VTAIL.n67 171.744
R987 VTAIL.n103 VTAIL.n67 171.744
R988 VTAIL.n104 VTAIL.n103 171.744
R989 VTAIL.n104 VTAIL.n63 171.744
R990 VTAIL.n111 VTAIL.n63 171.744
R991 VTAIL.n112 VTAIL.n111 171.744
R992 VTAIL.n138 VTAIL.n135 171.744
R993 VTAIL.n145 VTAIL.n135 171.744
R994 VTAIL.n146 VTAIL.n145 171.744
R995 VTAIL.n146 VTAIL.n131 171.744
R996 VTAIL.n153 VTAIL.n131 171.744
R997 VTAIL.n155 VTAIL.n153 171.744
R998 VTAIL.n155 VTAIL.n154 171.744
R999 VTAIL.n154 VTAIL.n127 171.744
R1000 VTAIL.n163 VTAIL.n127 171.744
R1001 VTAIL.n164 VTAIL.n163 171.744
R1002 VTAIL.n164 VTAIL.n123 171.744
R1003 VTAIL.n171 VTAIL.n123 171.744
R1004 VTAIL.n172 VTAIL.n171 171.744
R1005 VTAIL.n408 VTAIL.n407 171.744
R1006 VTAIL.n407 VTAIL.n359 171.744
R1007 VTAIL.n400 VTAIL.n359 171.744
R1008 VTAIL.n400 VTAIL.n399 171.744
R1009 VTAIL.n399 VTAIL.n363 171.744
R1010 VTAIL.n367 VTAIL.n363 171.744
R1011 VTAIL.n391 VTAIL.n367 171.744
R1012 VTAIL.n391 VTAIL.n390 171.744
R1013 VTAIL.n390 VTAIL.n368 171.744
R1014 VTAIL.n383 VTAIL.n368 171.744
R1015 VTAIL.n383 VTAIL.n382 171.744
R1016 VTAIL.n382 VTAIL.n372 171.744
R1017 VTAIL.n375 VTAIL.n372 171.744
R1018 VTAIL.n348 VTAIL.n347 171.744
R1019 VTAIL.n347 VTAIL.n299 171.744
R1020 VTAIL.n340 VTAIL.n299 171.744
R1021 VTAIL.n340 VTAIL.n339 171.744
R1022 VTAIL.n339 VTAIL.n303 171.744
R1023 VTAIL.n307 VTAIL.n303 171.744
R1024 VTAIL.n331 VTAIL.n307 171.744
R1025 VTAIL.n331 VTAIL.n330 171.744
R1026 VTAIL.n330 VTAIL.n308 171.744
R1027 VTAIL.n323 VTAIL.n308 171.744
R1028 VTAIL.n323 VTAIL.n322 171.744
R1029 VTAIL.n322 VTAIL.n312 171.744
R1030 VTAIL.n315 VTAIL.n312 171.744
R1031 VTAIL.n290 VTAIL.n289 171.744
R1032 VTAIL.n289 VTAIL.n241 171.744
R1033 VTAIL.n282 VTAIL.n241 171.744
R1034 VTAIL.n282 VTAIL.n281 171.744
R1035 VTAIL.n281 VTAIL.n245 171.744
R1036 VTAIL.n249 VTAIL.n245 171.744
R1037 VTAIL.n273 VTAIL.n249 171.744
R1038 VTAIL.n273 VTAIL.n272 171.744
R1039 VTAIL.n272 VTAIL.n250 171.744
R1040 VTAIL.n265 VTAIL.n250 171.744
R1041 VTAIL.n265 VTAIL.n264 171.744
R1042 VTAIL.n264 VTAIL.n254 171.744
R1043 VTAIL.n257 VTAIL.n254 171.744
R1044 VTAIL.n230 VTAIL.n229 171.744
R1045 VTAIL.n229 VTAIL.n181 171.744
R1046 VTAIL.n222 VTAIL.n181 171.744
R1047 VTAIL.n222 VTAIL.n221 171.744
R1048 VTAIL.n221 VTAIL.n185 171.744
R1049 VTAIL.n189 VTAIL.n185 171.744
R1050 VTAIL.n213 VTAIL.n189 171.744
R1051 VTAIL.n213 VTAIL.n212 171.744
R1052 VTAIL.n212 VTAIL.n190 171.744
R1053 VTAIL.n205 VTAIL.n190 171.744
R1054 VTAIL.n205 VTAIL.n204 171.744
R1055 VTAIL.n204 VTAIL.n194 171.744
R1056 VTAIL.n197 VTAIL.n194 171.744
R1057 VTAIL.n432 VTAIL.t1 85.8723
R1058 VTAIL.n20 VTAIL.t0 85.8723
R1059 VTAIL.n78 VTAIL.t10 85.8723
R1060 VTAIL.n138 VTAIL.t13 85.8723
R1061 VTAIL.n375 VTAIL.t8 85.8723
R1062 VTAIL.n315 VTAIL.t15 85.8723
R1063 VTAIL.n257 VTAIL.t3 85.8723
R1064 VTAIL.n197 VTAIL.t6 85.8723
R1065 VTAIL.n355 VTAIL.n354 60.9328
R1066 VTAIL.n237 VTAIL.n236 60.9328
R1067 VTAIL.n1 VTAIL.n0 60.9326
R1068 VTAIL.n119 VTAIL.n118 60.9326
R1069 VTAIL.n471 VTAIL.n470 33.9308
R1070 VTAIL.n59 VTAIL.n58 33.9308
R1071 VTAIL.n117 VTAIL.n116 33.9308
R1072 VTAIL.n177 VTAIL.n176 33.9308
R1073 VTAIL.n413 VTAIL.n412 33.9308
R1074 VTAIL.n353 VTAIL.n352 33.9308
R1075 VTAIL.n295 VTAIL.n294 33.9308
R1076 VTAIL.n235 VTAIL.n234 33.9308
R1077 VTAIL.n471 VTAIL.n413 22.3238
R1078 VTAIL.n235 VTAIL.n177 22.3238
R1079 VTAIL.n456 VTAIL.n455 13.1884
R1080 VTAIL.n44 VTAIL.n43 13.1884
R1081 VTAIL.n102 VTAIL.n101 13.1884
R1082 VTAIL.n162 VTAIL.n161 13.1884
R1083 VTAIL.n398 VTAIL.n397 13.1884
R1084 VTAIL.n338 VTAIL.n337 13.1884
R1085 VTAIL.n280 VTAIL.n279 13.1884
R1086 VTAIL.n220 VTAIL.n219 13.1884
R1087 VTAIL.n454 VTAIL.n422 12.8005
R1088 VTAIL.n459 VTAIL.n420 12.8005
R1089 VTAIL.n42 VTAIL.n10 12.8005
R1090 VTAIL.n47 VTAIL.n8 12.8005
R1091 VTAIL.n100 VTAIL.n68 12.8005
R1092 VTAIL.n105 VTAIL.n66 12.8005
R1093 VTAIL.n160 VTAIL.n128 12.8005
R1094 VTAIL.n165 VTAIL.n126 12.8005
R1095 VTAIL.n401 VTAIL.n362 12.8005
R1096 VTAIL.n396 VTAIL.n364 12.8005
R1097 VTAIL.n341 VTAIL.n302 12.8005
R1098 VTAIL.n336 VTAIL.n304 12.8005
R1099 VTAIL.n283 VTAIL.n244 12.8005
R1100 VTAIL.n278 VTAIL.n246 12.8005
R1101 VTAIL.n223 VTAIL.n184 12.8005
R1102 VTAIL.n218 VTAIL.n186 12.8005
R1103 VTAIL.n451 VTAIL.n450 12.0247
R1104 VTAIL.n460 VTAIL.n418 12.0247
R1105 VTAIL.n39 VTAIL.n38 12.0247
R1106 VTAIL.n48 VTAIL.n6 12.0247
R1107 VTAIL.n97 VTAIL.n96 12.0247
R1108 VTAIL.n106 VTAIL.n64 12.0247
R1109 VTAIL.n157 VTAIL.n156 12.0247
R1110 VTAIL.n166 VTAIL.n124 12.0247
R1111 VTAIL.n402 VTAIL.n360 12.0247
R1112 VTAIL.n393 VTAIL.n392 12.0247
R1113 VTAIL.n342 VTAIL.n300 12.0247
R1114 VTAIL.n333 VTAIL.n332 12.0247
R1115 VTAIL.n284 VTAIL.n242 12.0247
R1116 VTAIL.n275 VTAIL.n274 12.0247
R1117 VTAIL.n224 VTAIL.n182 12.0247
R1118 VTAIL.n215 VTAIL.n214 12.0247
R1119 VTAIL.n446 VTAIL.n424 11.249
R1120 VTAIL.n464 VTAIL.n463 11.249
R1121 VTAIL.n34 VTAIL.n12 11.249
R1122 VTAIL.n52 VTAIL.n51 11.249
R1123 VTAIL.n92 VTAIL.n70 11.249
R1124 VTAIL.n110 VTAIL.n109 11.249
R1125 VTAIL.n152 VTAIL.n130 11.249
R1126 VTAIL.n170 VTAIL.n169 11.249
R1127 VTAIL.n406 VTAIL.n405 11.249
R1128 VTAIL.n389 VTAIL.n366 11.249
R1129 VTAIL.n346 VTAIL.n345 11.249
R1130 VTAIL.n329 VTAIL.n306 11.249
R1131 VTAIL.n288 VTAIL.n287 11.249
R1132 VTAIL.n271 VTAIL.n248 11.249
R1133 VTAIL.n228 VTAIL.n227 11.249
R1134 VTAIL.n211 VTAIL.n188 11.249
R1135 VTAIL.n433 VTAIL.n431 10.7239
R1136 VTAIL.n21 VTAIL.n19 10.7239
R1137 VTAIL.n79 VTAIL.n77 10.7239
R1138 VTAIL.n139 VTAIL.n137 10.7239
R1139 VTAIL.n376 VTAIL.n374 10.7239
R1140 VTAIL.n316 VTAIL.n314 10.7239
R1141 VTAIL.n258 VTAIL.n256 10.7239
R1142 VTAIL.n198 VTAIL.n196 10.7239
R1143 VTAIL.n445 VTAIL.n426 10.4732
R1144 VTAIL.n467 VTAIL.n416 10.4732
R1145 VTAIL.n33 VTAIL.n14 10.4732
R1146 VTAIL.n55 VTAIL.n4 10.4732
R1147 VTAIL.n91 VTAIL.n72 10.4732
R1148 VTAIL.n113 VTAIL.n62 10.4732
R1149 VTAIL.n151 VTAIL.n132 10.4732
R1150 VTAIL.n173 VTAIL.n122 10.4732
R1151 VTAIL.n409 VTAIL.n358 10.4732
R1152 VTAIL.n388 VTAIL.n369 10.4732
R1153 VTAIL.n349 VTAIL.n298 10.4732
R1154 VTAIL.n328 VTAIL.n309 10.4732
R1155 VTAIL.n291 VTAIL.n240 10.4732
R1156 VTAIL.n270 VTAIL.n251 10.4732
R1157 VTAIL.n231 VTAIL.n180 10.4732
R1158 VTAIL.n210 VTAIL.n191 10.4732
R1159 VTAIL.n442 VTAIL.n441 9.69747
R1160 VTAIL.n468 VTAIL.n414 9.69747
R1161 VTAIL.n30 VTAIL.n29 9.69747
R1162 VTAIL.n56 VTAIL.n2 9.69747
R1163 VTAIL.n88 VTAIL.n87 9.69747
R1164 VTAIL.n114 VTAIL.n60 9.69747
R1165 VTAIL.n148 VTAIL.n147 9.69747
R1166 VTAIL.n174 VTAIL.n120 9.69747
R1167 VTAIL.n410 VTAIL.n356 9.69747
R1168 VTAIL.n385 VTAIL.n384 9.69747
R1169 VTAIL.n350 VTAIL.n296 9.69747
R1170 VTAIL.n325 VTAIL.n324 9.69747
R1171 VTAIL.n292 VTAIL.n238 9.69747
R1172 VTAIL.n267 VTAIL.n266 9.69747
R1173 VTAIL.n232 VTAIL.n178 9.69747
R1174 VTAIL.n207 VTAIL.n206 9.69747
R1175 VTAIL.n470 VTAIL.n469 9.45567
R1176 VTAIL.n58 VTAIL.n57 9.45567
R1177 VTAIL.n116 VTAIL.n115 9.45567
R1178 VTAIL.n176 VTAIL.n175 9.45567
R1179 VTAIL.n412 VTAIL.n411 9.45567
R1180 VTAIL.n352 VTAIL.n351 9.45567
R1181 VTAIL.n294 VTAIL.n293 9.45567
R1182 VTAIL.n234 VTAIL.n233 9.45567
R1183 VTAIL.n469 VTAIL.n468 9.3005
R1184 VTAIL.n416 VTAIL.n415 9.3005
R1185 VTAIL.n463 VTAIL.n462 9.3005
R1186 VTAIL.n461 VTAIL.n460 9.3005
R1187 VTAIL.n420 VTAIL.n419 9.3005
R1188 VTAIL.n435 VTAIL.n434 9.3005
R1189 VTAIL.n437 VTAIL.n436 9.3005
R1190 VTAIL.n428 VTAIL.n427 9.3005
R1191 VTAIL.n443 VTAIL.n442 9.3005
R1192 VTAIL.n445 VTAIL.n444 9.3005
R1193 VTAIL.n424 VTAIL.n423 9.3005
R1194 VTAIL.n452 VTAIL.n451 9.3005
R1195 VTAIL.n454 VTAIL.n453 9.3005
R1196 VTAIL.n57 VTAIL.n56 9.3005
R1197 VTAIL.n4 VTAIL.n3 9.3005
R1198 VTAIL.n51 VTAIL.n50 9.3005
R1199 VTAIL.n49 VTAIL.n48 9.3005
R1200 VTAIL.n8 VTAIL.n7 9.3005
R1201 VTAIL.n23 VTAIL.n22 9.3005
R1202 VTAIL.n25 VTAIL.n24 9.3005
R1203 VTAIL.n16 VTAIL.n15 9.3005
R1204 VTAIL.n31 VTAIL.n30 9.3005
R1205 VTAIL.n33 VTAIL.n32 9.3005
R1206 VTAIL.n12 VTAIL.n11 9.3005
R1207 VTAIL.n40 VTAIL.n39 9.3005
R1208 VTAIL.n42 VTAIL.n41 9.3005
R1209 VTAIL.n115 VTAIL.n114 9.3005
R1210 VTAIL.n62 VTAIL.n61 9.3005
R1211 VTAIL.n109 VTAIL.n108 9.3005
R1212 VTAIL.n107 VTAIL.n106 9.3005
R1213 VTAIL.n66 VTAIL.n65 9.3005
R1214 VTAIL.n81 VTAIL.n80 9.3005
R1215 VTAIL.n83 VTAIL.n82 9.3005
R1216 VTAIL.n74 VTAIL.n73 9.3005
R1217 VTAIL.n89 VTAIL.n88 9.3005
R1218 VTAIL.n91 VTAIL.n90 9.3005
R1219 VTAIL.n70 VTAIL.n69 9.3005
R1220 VTAIL.n98 VTAIL.n97 9.3005
R1221 VTAIL.n100 VTAIL.n99 9.3005
R1222 VTAIL.n175 VTAIL.n174 9.3005
R1223 VTAIL.n122 VTAIL.n121 9.3005
R1224 VTAIL.n169 VTAIL.n168 9.3005
R1225 VTAIL.n167 VTAIL.n166 9.3005
R1226 VTAIL.n126 VTAIL.n125 9.3005
R1227 VTAIL.n141 VTAIL.n140 9.3005
R1228 VTAIL.n143 VTAIL.n142 9.3005
R1229 VTAIL.n134 VTAIL.n133 9.3005
R1230 VTAIL.n149 VTAIL.n148 9.3005
R1231 VTAIL.n151 VTAIL.n150 9.3005
R1232 VTAIL.n130 VTAIL.n129 9.3005
R1233 VTAIL.n158 VTAIL.n157 9.3005
R1234 VTAIL.n160 VTAIL.n159 9.3005
R1235 VTAIL.n378 VTAIL.n377 9.3005
R1236 VTAIL.n380 VTAIL.n379 9.3005
R1237 VTAIL.n371 VTAIL.n370 9.3005
R1238 VTAIL.n386 VTAIL.n385 9.3005
R1239 VTAIL.n388 VTAIL.n387 9.3005
R1240 VTAIL.n366 VTAIL.n365 9.3005
R1241 VTAIL.n394 VTAIL.n393 9.3005
R1242 VTAIL.n396 VTAIL.n395 9.3005
R1243 VTAIL.n411 VTAIL.n410 9.3005
R1244 VTAIL.n358 VTAIL.n357 9.3005
R1245 VTAIL.n405 VTAIL.n404 9.3005
R1246 VTAIL.n403 VTAIL.n402 9.3005
R1247 VTAIL.n362 VTAIL.n361 9.3005
R1248 VTAIL.n318 VTAIL.n317 9.3005
R1249 VTAIL.n320 VTAIL.n319 9.3005
R1250 VTAIL.n311 VTAIL.n310 9.3005
R1251 VTAIL.n326 VTAIL.n325 9.3005
R1252 VTAIL.n328 VTAIL.n327 9.3005
R1253 VTAIL.n306 VTAIL.n305 9.3005
R1254 VTAIL.n334 VTAIL.n333 9.3005
R1255 VTAIL.n336 VTAIL.n335 9.3005
R1256 VTAIL.n351 VTAIL.n350 9.3005
R1257 VTAIL.n298 VTAIL.n297 9.3005
R1258 VTAIL.n345 VTAIL.n344 9.3005
R1259 VTAIL.n343 VTAIL.n342 9.3005
R1260 VTAIL.n302 VTAIL.n301 9.3005
R1261 VTAIL.n260 VTAIL.n259 9.3005
R1262 VTAIL.n262 VTAIL.n261 9.3005
R1263 VTAIL.n253 VTAIL.n252 9.3005
R1264 VTAIL.n268 VTAIL.n267 9.3005
R1265 VTAIL.n270 VTAIL.n269 9.3005
R1266 VTAIL.n248 VTAIL.n247 9.3005
R1267 VTAIL.n276 VTAIL.n275 9.3005
R1268 VTAIL.n278 VTAIL.n277 9.3005
R1269 VTAIL.n293 VTAIL.n292 9.3005
R1270 VTAIL.n240 VTAIL.n239 9.3005
R1271 VTAIL.n287 VTAIL.n286 9.3005
R1272 VTAIL.n285 VTAIL.n284 9.3005
R1273 VTAIL.n244 VTAIL.n243 9.3005
R1274 VTAIL.n200 VTAIL.n199 9.3005
R1275 VTAIL.n202 VTAIL.n201 9.3005
R1276 VTAIL.n193 VTAIL.n192 9.3005
R1277 VTAIL.n208 VTAIL.n207 9.3005
R1278 VTAIL.n210 VTAIL.n209 9.3005
R1279 VTAIL.n188 VTAIL.n187 9.3005
R1280 VTAIL.n216 VTAIL.n215 9.3005
R1281 VTAIL.n218 VTAIL.n217 9.3005
R1282 VTAIL.n233 VTAIL.n232 9.3005
R1283 VTAIL.n180 VTAIL.n179 9.3005
R1284 VTAIL.n227 VTAIL.n226 9.3005
R1285 VTAIL.n225 VTAIL.n224 9.3005
R1286 VTAIL.n184 VTAIL.n183 9.3005
R1287 VTAIL.n438 VTAIL.n428 8.92171
R1288 VTAIL.n26 VTAIL.n16 8.92171
R1289 VTAIL.n84 VTAIL.n74 8.92171
R1290 VTAIL.n144 VTAIL.n134 8.92171
R1291 VTAIL.n381 VTAIL.n371 8.92171
R1292 VTAIL.n321 VTAIL.n311 8.92171
R1293 VTAIL.n263 VTAIL.n253 8.92171
R1294 VTAIL.n203 VTAIL.n193 8.92171
R1295 VTAIL.n437 VTAIL.n430 8.14595
R1296 VTAIL.n25 VTAIL.n18 8.14595
R1297 VTAIL.n83 VTAIL.n76 8.14595
R1298 VTAIL.n143 VTAIL.n136 8.14595
R1299 VTAIL.n380 VTAIL.n373 8.14595
R1300 VTAIL.n320 VTAIL.n313 8.14595
R1301 VTAIL.n262 VTAIL.n255 8.14595
R1302 VTAIL.n202 VTAIL.n195 8.14595
R1303 VTAIL.n434 VTAIL.n433 7.3702
R1304 VTAIL.n22 VTAIL.n21 7.3702
R1305 VTAIL.n80 VTAIL.n79 7.3702
R1306 VTAIL.n140 VTAIL.n139 7.3702
R1307 VTAIL.n377 VTAIL.n376 7.3702
R1308 VTAIL.n317 VTAIL.n316 7.3702
R1309 VTAIL.n259 VTAIL.n258 7.3702
R1310 VTAIL.n199 VTAIL.n198 7.3702
R1311 VTAIL.n434 VTAIL.n430 5.81868
R1312 VTAIL.n22 VTAIL.n18 5.81868
R1313 VTAIL.n80 VTAIL.n76 5.81868
R1314 VTAIL.n140 VTAIL.n136 5.81868
R1315 VTAIL.n377 VTAIL.n373 5.81868
R1316 VTAIL.n317 VTAIL.n313 5.81868
R1317 VTAIL.n259 VTAIL.n255 5.81868
R1318 VTAIL.n199 VTAIL.n195 5.81868
R1319 VTAIL.n438 VTAIL.n437 5.04292
R1320 VTAIL.n26 VTAIL.n25 5.04292
R1321 VTAIL.n84 VTAIL.n83 5.04292
R1322 VTAIL.n144 VTAIL.n143 5.04292
R1323 VTAIL.n381 VTAIL.n380 5.04292
R1324 VTAIL.n321 VTAIL.n320 5.04292
R1325 VTAIL.n263 VTAIL.n262 5.04292
R1326 VTAIL.n203 VTAIL.n202 5.04292
R1327 VTAIL.n441 VTAIL.n428 4.26717
R1328 VTAIL.n470 VTAIL.n414 4.26717
R1329 VTAIL.n29 VTAIL.n16 4.26717
R1330 VTAIL.n58 VTAIL.n2 4.26717
R1331 VTAIL.n87 VTAIL.n74 4.26717
R1332 VTAIL.n116 VTAIL.n60 4.26717
R1333 VTAIL.n147 VTAIL.n134 4.26717
R1334 VTAIL.n176 VTAIL.n120 4.26717
R1335 VTAIL.n412 VTAIL.n356 4.26717
R1336 VTAIL.n384 VTAIL.n371 4.26717
R1337 VTAIL.n352 VTAIL.n296 4.26717
R1338 VTAIL.n324 VTAIL.n311 4.26717
R1339 VTAIL.n294 VTAIL.n238 4.26717
R1340 VTAIL.n266 VTAIL.n253 4.26717
R1341 VTAIL.n234 VTAIL.n178 4.26717
R1342 VTAIL.n206 VTAIL.n193 4.26717
R1343 VTAIL.n442 VTAIL.n426 3.49141
R1344 VTAIL.n468 VTAIL.n467 3.49141
R1345 VTAIL.n30 VTAIL.n14 3.49141
R1346 VTAIL.n56 VTAIL.n55 3.49141
R1347 VTAIL.n88 VTAIL.n72 3.49141
R1348 VTAIL.n114 VTAIL.n113 3.49141
R1349 VTAIL.n148 VTAIL.n132 3.49141
R1350 VTAIL.n174 VTAIL.n173 3.49141
R1351 VTAIL.n410 VTAIL.n409 3.49141
R1352 VTAIL.n385 VTAIL.n369 3.49141
R1353 VTAIL.n350 VTAIL.n349 3.49141
R1354 VTAIL.n325 VTAIL.n309 3.49141
R1355 VTAIL.n292 VTAIL.n291 3.49141
R1356 VTAIL.n267 VTAIL.n251 3.49141
R1357 VTAIL.n232 VTAIL.n231 3.49141
R1358 VTAIL.n207 VTAIL.n191 3.49141
R1359 VTAIL.n0 VTAIL.t4 3.01861
R1360 VTAIL.n0 VTAIL.t2 3.01861
R1361 VTAIL.n118 VTAIL.t14 3.01861
R1362 VTAIL.n118 VTAIL.t12 3.01861
R1363 VTAIL.n354 VTAIL.t9 3.01861
R1364 VTAIL.n354 VTAIL.t11 3.01861
R1365 VTAIL.n236 VTAIL.t5 3.01861
R1366 VTAIL.n236 VTAIL.t7 3.01861
R1367 VTAIL.n446 VTAIL.n445 2.71565
R1368 VTAIL.n464 VTAIL.n416 2.71565
R1369 VTAIL.n34 VTAIL.n33 2.71565
R1370 VTAIL.n52 VTAIL.n4 2.71565
R1371 VTAIL.n92 VTAIL.n91 2.71565
R1372 VTAIL.n110 VTAIL.n62 2.71565
R1373 VTAIL.n152 VTAIL.n151 2.71565
R1374 VTAIL.n170 VTAIL.n122 2.71565
R1375 VTAIL.n406 VTAIL.n358 2.71565
R1376 VTAIL.n389 VTAIL.n388 2.71565
R1377 VTAIL.n346 VTAIL.n298 2.71565
R1378 VTAIL.n329 VTAIL.n328 2.71565
R1379 VTAIL.n288 VTAIL.n240 2.71565
R1380 VTAIL.n271 VTAIL.n270 2.71565
R1381 VTAIL.n228 VTAIL.n180 2.71565
R1382 VTAIL.n211 VTAIL.n210 2.71565
R1383 VTAIL.n435 VTAIL.n431 2.41282
R1384 VTAIL.n23 VTAIL.n19 2.41282
R1385 VTAIL.n81 VTAIL.n77 2.41282
R1386 VTAIL.n141 VTAIL.n137 2.41282
R1387 VTAIL.n378 VTAIL.n374 2.41282
R1388 VTAIL.n318 VTAIL.n314 2.41282
R1389 VTAIL.n260 VTAIL.n256 2.41282
R1390 VTAIL.n200 VTAIL.n196 2.41282
R1391 VTAIL.n450 VTAIL.n424 1.93989
R1392 VTAIL.n463 VTAIL.n418 1.93989
R1393 VTAIL.n38 VTAIL.n12 1.93989
R1394 VTAIL.n51 VTAIL.n6 1.93989
R1395 VTAIL.n96 VTAIL.n70 1.93989
R1396 VTAIL.n109 VTAIL.n64 1.93989
R1397 VTAIL.n156 VTAIL.n130 1.93989
R1398 VTAIL.n169 VTAIL.n124 1.93989
R1399 VTAIL.n405 VTAIL.n360 1.93989
R1400 VTAIL.n392 VTAIL.n366 1.93989
R1401 VTAIL.n345 VTAIL.n300 1.93989
R1402 VTAIL.n332 VTAIL.n306 1.93989
R1403 VTAIL.n287 VTAIL.n242 1.93989
R1404 VTAIL.n274 VTAIL.n248 1.93989
R1405 VTAIL.n227 VTAIL.n182 1.93989
R1406 VTAIL.n214 VTAIL.n188 1.93989
R1407 VTAIL.n451 VTAIL.n422 1.16414
R1408 VTAIL.n460 VTAIL.n459 1.16414
R1409 VTAIL.n39 VTAIL.n10 1.16414
R1410 VTAIL.n48 VTAIL.n47 1.16414
R1411 VTAIL.n97 VTAIL.n68 1.16414
R1412 VTAIL.n106 VTAIL.n105 1.16414
R1413 VTAIL.n157 VTAIL.n128 1.16414
R1414 VTAIL.n166 VTAIL.n165 1.16414
R1415 VTAIL.n402 VTAIL.n401 1.16414
R1416 VTAIL.n393 VTAIL.n364 1.16414
R1417 VTAIL.n342 VTAIL.n341 1.16414
R1418 VTAIL.n333 VTAIL.n304 1.16414
R1419 VTAIL.n284 VTAIL.n283 1.16414
R1420 VTAIL.n275 VTAIL.n246 1.16414
R1421 VTAIL.n224 VTAIL.n223 1.16414
R1422 VTAIL.n215 VTAIL.n186 1.16414
R1423 VTAIL.n237 VTAIL.n235 0.672914
R1424 VTAIL.n295 VTAIL.n237 0.672914
R1425 VTAIL.n355 VTAIL.n353 0.672914
R1426 VTAIL.n413 VTAIL.n355 0.672914
R1427 VTAIL.n177 VTAIL.n119 0.672914
R1428 VTAIL.n119 VTAIL.n117 0.672914
R1429 VTAIL.n59 VTAIL.n1 0.672914
R1430 VTAIL VTAIL.n471 0.614724
R1431 VTAIL.n353 VTAIL.n295 0.470328
R1432 VTAIL.n117 VTAIL.n59 0.470328
R1433 VTAIL.n455 VTAIL.n454 0.388379
R1434 VTAIL.n456 VTAIL.n420 0.388379
R1435 VTAIL.n43 VTAIL.n42 0.388379
R1436 VTAIL.n44 VTAIL.n8 0.388379
R1437 VTAIL.n101 VTAIL.n100 0.388379
R1438 VTAIL.n102 VTAIL.n66 0.388379
R1439 VTAIL.n161 VTAIL.n160 0.388379
R1440 VTAIL.n162 VTAIL.n126 0.388379
R1441 VTAIL.n398 VTAIL.n362 0.388379
R1442 VTAIL.n397 VTAIL.n396 0.388379
R1443 VTAIL.n338 VTAIL.n302 0.388379
R1444 VTAIL.n337 VTAIL.n336 0.388379
R1445 VTAIL.n280 VTAIL.n244 0.388379
R1446 VTAIL.n279 VTAIL.n278 0.388379
R1447 VTAIL.n220 VTAIL.n184 0.388379
R1448 VTAIL.n219 VTAIL.n218 0.388379
R1449 VTAIL.n436 VTAIL.n435 0.155672
R1450 VTAIL.n436 VTAIL.n427 0.155672
R1451 VTAIL.n443 VTAIL.n427 0.155672
R1452 VTAIL.n444 VTAIL.n443 0.155672
R1453 VTAIL.n444 VTAIL.n423 0.155672
R1454 VTAIL.n452 VTAIL.n423 0.155672
R1455 VTAIL.n453 VTAIL.n452 0.155672
R1456 VTAIL.n453 VTAIL.n419 0.155672
R1457 VTAIL.n461 VTAIL.n419 0.155672
R1458 VTAIL.n462 VTAIL.n461 0.155672
R1459 VTAIL.n462 VTAIL.n415 0.155672
R1460 VTAIL.n469 VTAIL.n415 0.155672
R1461 VTAIL.n24 VTAIL.n23 0.155672
R1462 VTAIL.n24 VTAIL.n15 0.155672
R1463 VTAIL.n31 VTAIL.n15 0.155672
R1464 VTAIL.n32 VTAIL.n31 0.155672
R1465 VTAIL.n32 VTAIL.n11 0.155672
R1466 VTAIL.n40 VTAIL.n11 0.155672
R1467 VTAIL.n41 VTAIL.n40 0.155672
R1468 VTAIL.n41 VTAIL.n7 0.155672
R1469 VTAIL.n49 VTAIL.n7 0.155672
R1470 VTAIL.n50 VTAIL.n49 0.155672
R1471 VTAIL.n50 VTAIL.n3 0.155672
R1472 VTAIL.n57 VTAIL.n3 0.155672
R1473 VTAIL.n82 VTAIL.n81 0.155672
R1474 VTAIL.n82 VTAIL.n73 0.155672
R1475 VTAIL.n89 VTAIL.n73 0.155672
R1476 VTAIL.n90 VTAIL.n89 0.155672
R1477 VTAIL.n90 VTAIL.n69 0.155672
R1478 VTAIL.n98 VTAIL.n69 0.155672
R1479 VTAIL.n99 VTAIL.n98 0.155672
R1480 VTAIL.n99 VTAIL.n65 0.155672
R1481 VTAIL.n107 VTAIL.n65 0.155672
R1482 VTAIL.n108 VTAIL.n107 0.155672
R1483 VTAIL.n108 VTAIL.n61 0.155672
R1484 VTAIL.n115 VTAIL.n61 0.155672
R1485 VTAIL.n142 VTAIL.n141 0.155672
R1486 VTAIL.n142 VTAIL.n133 0.155672
R1487 VTAIL.n149 VTAIL.n133 0.155672
R1488 VTAIL.n150 VTAIL.n149 0.155672
R1489 VTAIL.n150 VTAIL.n129 0.155672
R1490 VTAIL.n158 VTAIL.n129 0.155672
R1491 VTAIL.n159 VTAIL.n158 0.155672
R1492 VTAIL.n159 VTAIL.n125 0.155672
R1493 VTAIL.n167 VTAIL.n125 0.155672
R1494 VTAIL.n168 VTAIL.n167 0.155672
R1495 VTAIL.n168 VTAIL.n121 0.155672
R1496 VTAIL.n175 VTAIL.n121 0.155672
R1497 VTAIL.n411 VTAIL.n357 0.155672
R1498 VTAIL.n404 VTAIL.n357 0.155672
R1499 VTAIL.n404 VTAIL.n403 0.155672
R1500 VTAIL.n403 VTAIL.n361 0.155672
R1501 VTAIL.n395 VTAIL.n361 0.155672
R1502 VTAIL.n395 VTAIL.n394 0.155672
R1503 VTAIL.n394 VTAIL.n365 0.155672
R1504 VTAIL.n387 VTAIL.n365 0.155672
R1505 VTAIL.n387 VTAIL.n386 0.155672
R1506 VTAIL.n386 VTAIL.n370 0.155672
R1507 VTAIL.n379 VTAIL.n370 0.155672
R1508 VTAIL.n379 VTAIL.n378 0.155672
R1509 VTAIL.n351 VTAIL.n297 0.155672
R1510 VTAIL.n344 VTAIL.n297 0.155672
R1511 VTAIL.n344 VTAIL.n343 0.155672
R1512 VTAIL.n343 VTAIL.n301 0.155672
R1513 VTAIL.n335 VTAIL.n301 0.155672
R1514 VTAIL.n335 VTAIL.n334 0.155672
R1515 VTAIL.n334 VTAIL.n305 0.155672
R1516 VTAIL.n327 VTAIL.n305 0.155672
R1517 VTAIL.n327 VTAIL.n326 0.155672
R1518 VTAIL.n326 VTAIL.n310 0.155672
R1519 VTAIL.n319 VTAIL.n310 0.155672
R1520 VTAIL.n319 VTAIL.n318 0.155672
R1521 VTAIL.n293 VTAIL.n239 0.155672
R1522 VTAIL.n286 VTAIL.n239 0.155672
R1523 VTAIL.n286 VTAIL.n285 0.155672
R1524 VTAIL.n285 VTAIL.n243 0.155672
R1525 VTAIL.n277 VTAIL.n243 0.155672
R1526 VTAIL.n277 VTAIL.n276 0.155672
R1527 VTAIL.n276 VTAIL.n247 0.155672
R1528 VTAIL.n269 VTAIL.n247 0.155672
R1529 VTAIL.n269 VTAIL.n268 0.155672
R1530 VTAIL.n268 VTAIL.n252 0.155672
R1531 VTAIL.n261 VTAIL.n252 0.155672
R1532 VTAIL.n261 VTAIL.n260 0.155672
R1533 VTAIL.n233 VTAIL.n179 0.155672
R1534 VTAIL.n226 VTAIL.n179 0.155672
R1535 VTAIL.n226 VTAIL.n225 0.155672
R1536 VTAIL.n225 VTAIL.n183 0.155672
R1537 VTAIL.n217 VTAIL.n183 0.155672
R1538 VTAIL.n217 VTAIL.n216 0.155672
R1539 VTAIL.n216 VTAIL.n187 0.155672
R1540 VTAIL.n209 VTAIL.n187 0.155672
R1541 VTAIL.n209 VTAIL.n208 0.155672
R1542 VTAIL.n208 VTAIL.n192 0.155672
R1543 VTAIL.n201 VTAIL.n192 0.155672
R1544 VTAIL.n201 VTAIL.n200 0.155672
R1545 VTAIL VTAIL.n1 0.0586897
R1546 VN.n2 VN.t7 685.606
R1547 VN.n10 VN.t1 685.606
R1548 VN.n1 VN.t5 664.625
R1549 VN.n5 VN.t4 664.625
R1550 VN.n6 VN.t3 664.625
R1551 VN.n9 VN.t6 664.625
R1552 VN.n13 VN.t2 664.625
R1553 VN.n14 VN.t0 664.625
R1554 VN.n7 VN.n6 161.3
R1555 VN.n15 VN.n14 161.3
R1556 VN.n13 VN.n8 161.3
R1557 VN.n12 VN.n11 161.3
R1558 VN.n5 VN.n0 161.3
R1559 VN.n4 VN.n3 161.3
R1560 VN.n11 VN.n10 70.4033
R1561 VN.n3 VN.n2 70.4033
R1562 VN.n6 VN.n5 48.2005
R1563 VN.n14 VN.n13 48.2005
R1564 VN VN.n15 40.3054
R1565 VN.n4 VN.n1 24.1005
R1566 VN.n5 VN.n4 24.1005
R1567 VN.n13 VN.n12 24.1005
R1568 VN.n12 VN.n9 24.1005
R1569 VN.n10 VN.n9 20.9576
R1570 VN.n2 VN.n1 20.9576
R1571 VN.n15 VN.n8 0.189894
R1572 VN.n11 VN.n8 0.189894
R1573 VN.n3 VN.n0 0.189894
R1574 VN.n7 VN.n0 0.189894
R1575 VN VN.n7 0.0516364
R1576 VDD2.n2 VDD2.n1 77.8923
R1577 VDD2.n2 VDD2.n0 77.8923
R1578 VDD2 VDD2.n5 77.8894
R1579 VDD2.n4 VDD2.n3 77.6116
R1580 VDD2.n4 VDD2.n2 36.0256
R1581 VDD2.n5 VDD2.t1 3.01861
R1582 VDD2.n5 VDD2.t6 3.01861
R1583 VDD2.n3 VDD2.t7 3.01861
R1584 VDD2.n3 VDD2.t5 3.01861
R1585 VDD2.n1 VDD2.t3 3.01861
R1586 VDD2.n1 VDD2.t4 3.01861
R1587 VDD2.n0 VDD2.t0 3.01861
R1588 VDD2.n0 VDD2.t2 3.01861
R1589 VDD2 VDD2.n4 0.394897
C0 VDD1 VP 4.03212f
C1 B w_n1750_n3122# 6.48214f
C2 VTAIL B 3.3119f
C3 VDD2 w_n1750_n3122# 1.19282f
C4 VDD2 VTAIL 12.4381f
C5 VDD1 w_n1750_n3122# 1.16834f
C6 VTAIL VDD1 12.3981f
C7 VP w_n1750_n3122# 3.16087f
C8 VTAIL VP 3.61326f
C9 VTAIL w_n1750_n3122# 3.92178f
C10 VN B 0.707475f
C11 VDD2 VN 3.88939f
C12 VDD1 VN 0.147876f
C13 VDD2 B 0.98949f
C14 VN VP 4.80635f
C15 VDD1 B 0.96054f
C16 VDD2 VDD1 0.704224f
C17 VN w_n1750_n3122# 2.94002f
C18 VP B 1.06623f
C19 VTAIL VN 3.59916f
C20 VDD2 VP 0.290923f
C21 VDD2 VSUBS 1.285159f
C22 VDD1 VSUBS 1.547103f
C23 VTAIL VSUBS 0.761351f
C24 VN VSUBS 4.42573f
C25 VP VSUBS 1.348084f
C26 B VSUBS 2.497035f
C27 w_n1750_n3122# VSUBS 67.389f
C28 VDD2.t0 VSUBS 0.254277f
C29 VDD2.t2 VSUBS 0.254277f
C30 VDD2.n0 VSUBS 1.95526f
C31 VDD2.t3 VSUBS 0.254277f
C32 VDD2.t4 VSUBS 0.254277f
C33 VDD2.n1 VSUBS 1.95526f
C34 VDD2.n2 VSUBS 2.9235f
C35 VDD2.t7 VSUBS 0.254277f
C36 VDD2.t5 VSUBS 0.254277f
C37 VDD2.n3 VSUBS 1.95293f
C38 VDD2.n4 VSUBS 2.81506f
C39 VDD2.t1 VSUBS 0.254277f
C40 VDD2.t6 VSUBS 0.254277f
C41 VDD2.n5 VSUBS 1.95523f
C42 VN.n0 VSUBS 0.062332f
C43 VN.t5 VSUBS 0.863368f
C44 VN.n1 VSUBS 0.36295f
C45 VN.t7 VSUBS 0.874284f
C46 VN.n2 VSUBS 0.346145f
C47 VN.n3 VSUBS 0.197688f
C48 VN.n4 VSUBS 0.014144f
C49 VN.t4 VSUBS 0.863368f
C50 VN.n5 VSUBS 0.36295f
C51 VN.t3 VSUBS 0.863368f
C52 VN.n6 VSUBS 0.356609f
C53 VN.n7 VSUBS 0.048305f
C54 VN.n8 VSUBS 0.062332f
C55 VN.t6 VSUBS 0.863368f
C56 VN.n9 VSUBS 0.36295f
C57 VN.t1 VSUBS 0.874284f
C58 VN.n10 VSUBS 0.346145f
C59 VN.n11 VSUBS 0.197688f
C60 VN.n12 VSUBS 0.014144f
C61 VN.t2 VSUBS 0.863368f
C62 VN.n13 VSUBS 0.36295f
C63 VN.t0 VSUBS 0.863368f
C64 VN.n14 VSUBS 0.356609f
C65 VN.n15 VSUBS 2.40197f
C66 VTAIL.t4 VSUBS 0.228014f
C67 VTAIL.t2 VSUBS 0.228014f
C68 VTAIL.n0 VSUBS 1.61943f
C69 VTAIL.n1 VSUBS 0.644986f
C70 VTAIL.n2 VSUBS 0.029439f
C71 VTAIL.n3 VSUBS 0.026791f
C72 VTAIL.n4 VSUBS 0.014396f
C73 VTAIL.n5 VSUBS 0.034028f
C74 VTAIL.n6 VSUBS 0.015243f
C75 VTAIL.n7 VSUBS 0.026791f
C76 VTAIL.n8 VSUBS 0.014396f
C77 VTAIL.n9 VSUBS 0.034028f
C78 VTAIL.n10 VSUBS 0.015243f
C79 VTAIL.n11 VSUBS 0.026791f
C80 VTAIL.n12 VSUBS 0.014396f
C81 VTAIL.n13 VSUBS 0.034028f
C82 VTAIL.n14 VSUBS 0.015243f
C83 VTAIL.n15 VSUBS 0.026791f
C84 VTAIL.n16 VSUBS 0.014396f
C85 VTAIL.n17 VSUBS 0.034028f
C86 VTAIL.n18 VSUBS 0.015243f
C87 VTAIL.n19 VSUBS 0.196107f
C88 VTAIL.t0 VSUBS 0.073227f
C89 VTAIL.n20 VSUBS 0.025521f
C90 VTAIL.n21 VSUBS 0.025598f
C91 VTAIL.n22 VSUBS 0.014396f
C92 VTAIL.n23 VSUBS 1.17193f
C93 VTAIL.n24 VSUBS 0.026791f
C94 VTAIL.n25 VSUBS 0.014396f
C95 VTAIL.n26 VSUBS 0.015243f
C96 VTAIL.n27 VSUBS 0.034028f
C97 VTAIL.n28 VSUBS 0.034028f
C98 VTAIL.n29 VSUBS 0.015243f
C99 VTAIL.n30 VSUBS 0.014396f
C100 VTAIL.n31 VSUBS 0.026791f
C101 VTAIL.n32 VSUBS 0.026791f
C102 VTAIL.n33 VSUBS 0.014396f
C103 VTAIL.n34 VSUBS 0.015243f
C104 VTAIL.n35 VSUBS 0.034028f
C105 VTAIL.n36 VSUBS 0.034028f
C106 VTAIL.n37 VSUBS 0.034028f
C107 VTAIL.n38 VSUBS 0.015243f
C108 VTAIL.n39 VSUBS 0.014396f
C109 VTAIL.n40 VSUBS 0.026791f
C110 VTAIL.n41 VSUBS 0.026791f
C111 VTAIL.n42 VSUBS 0.014396f
C112 VTAIL.n43 VSUBS 0.01482f
C113 VTAIL.n44 VSUBS 0.01482f
C114 VTAIL.n45 VSUBS 0.034028f
C115 VTAIL.n46 VSUBS 0.034028f
C116 VTAIL.n47 VSUBS 0.015243f
C117 VTAIL.n48 VSUBS 0.014396f
C118 VTAIL.n49 VSUBS 0.026791f
C119 VTAIL.n50 VSUBS 0.026791f
C120 VTAIL.n51 VSUBS 0.014396f
C121 VTAIL.n52 VSUBS 0.015243f
C122 VTAIL.n53 VSUBS 0.034028f
C123 VTAIL.n54 VSUBS 0.082383f
C124 VTAIL.n55 VSUBS 0.015243f
C125 VTAIL.n56 VSUBS 0.014396f
C126 VTAIL.n57 VSUBS 0.06522f
C127 VTAIL.n58 VSUBS 0.041529f
C128 VTAIL.n59 VSUBS 0.12335f
C129 VTAIL.n60 VSUBS 0.029439f
C130 VTAIL.n61 VSUBS 0.026791f
C131 VTAIL.n62 VSUBS 0.014396f
C132 VTAIL.n63 VSUBS 0.034028f
C133 VTAIL.n64 VSUBS 0.015243f
C134 VTAIL.n65 VSUBS 0.026791f
C135 VTAIL.n66 VSUBS 0.014396f
C136 VTAIL.n67 VSUBS 0.034028f
C137 VTAIL.n68 VSUBS 0.015243f
C138 VTAIL.n69 VSUBS 0.026791f
C139 VTAIL.n70 VSUBS 0.014396f
C140 VTAIL.n71 VSUBS 0.034028f
C141 VTAIL.n72 VSUBS 0.015243f
C142 VTAIL.n73 VSUBS 0.026791f
C143 VTAIL.n74 VSUBS 0.014396f
C144 VTAIL.n75 VSUBS 0.034028f
C145 VTAIL.n76 VSUBS 0.015243f
C146 VTAIL.n77 VSUBS 0.196107f
C147 VTAIL.t10 VSUBS 0.073227f
C148 VTAIL.n78 VSUBS 0.025521f
C149 VTAIL.n79 VSUBS 0.025598f
C150 VTAIL.n80 VSUBS 0.014396f
C151 VTAIL.n81 VSUBS 1.17193f
C152 VTAIL.n82 VSUBS 0.026791f
C153 VTAIL.n83 VSUBS 0.014396f
C154 VTAIL.n84 VSUBS 0.015243f
C155 VTAIL.n85 VSUBS 0.034028f
C156 VTAIL.n86 VSUBS 0.034028f
C157 VTAIL.n87 VSUBS 0.015243f
C158 VTAIL.n88 VSUBS 0.014396f
C159 VTAIL.n89 VSUBS 0.026791f
C160 VTAIL.n90 VSUBS 0.026791f
C161 VTAIL.n91 VSUBS 0.014396f
C162 VTAIL.n92 VSUBS 0.015243f
C163 VTAIL.n93 VSUBS 0.034028f
C164 VTAIL.n94 VSUBS 0.034028f
C165 VTAIL.n95 VSUBS 0.034028f
C166 VTAIL.n96 VSUBS 0.015243f
C167 VTAIL.n97 VSUBS 0.014396f
C168 VTAIL.n98 VSUBS 0.026791f
C169 VTAIL.n99 VSUBS 0.026791f
C170 VTAIL.n100 VSUBS 0.014396f
C171 VTAIL.n101 VSUBS 0.01482f
C172 VTAIL.n102 VSUBS 0.01482f
C173 VTAIL.n103 VSUBS 0.034028f
C174 VTAIL.n104 VSUBS 0.034028f
C175 VTAIL.n105 VSUBS 0.015243f
C176 VTAIL.n106 VSUBS 0.014396f
C177 VTAIL.n107 VSUBS 0.026791f
C178 VTAIL.n108 VSUBS 0.026791f
C179 VTAIL.n109 VSUBS 0.014396f
C180 VTAIL.n110 VSUBS 0.015243f
C181 VTAIL.n111 VSUBS 0.034028f
C182 VTAIL.n112 VSUBS 0.082383f
C183 VTAIL.n113 VSUBS 0.015243f
C184 VTAIL.n114 VSUBS 0.014396f
C185 VTAIL.n115 VSUBS 0.06522f
C186 VTAIL.n116 VSUBS 0.041529f
C187 VTAIL.n117 VSUBS 0.12335f
C188 VTAIL.t14 VSUBS 0.228014f
C189 VTAIL.t12 VSUBS 0.228014f
C190 VTAIL.n118 VSUBS 1.61943f
C191 VTAIL.n119 VSUBS 0.69801f
C192 VTAIL.n120 VSUBS 0.029439f
C193 VTAIL.n121 VSUBS 0.026791f
C194 VTAIL.n122 VSUBS 0.014396f
C195 VTAIL.n123 VSUBS 0.034028f
C196 VTAIL.n124 VSUBS 0.015243f
C197 VTAIL.n125 VSUBS 0.026791f
C198 VTAIL.n126 VSUBS 0.014396f
C199 VTAIL.n127 VSUBS 0.034028f
C200 VTAIL.n128 VSUBS 0.015243f
C201 VTAIL.n129 VSUBS 0.026791f
C202 VTAIL.n130 VSUBS 0.014396f
C203 VTAIL.n131 VSUBS 0.034028f
C204 VTAIL.n132 VSUBS 0.015243f
C205 VTAIL.n133 VSUBS 0.026791f
C206 VTAIL.n134 VSUBS 0.014396f
C207 VTAIL.n135 VSUBS 0.034028f
C208 VTAIL.n136 VSUBS 0.015243f
C209 VTAIL.n137 VSUBS 0.196107f
C210 VTAIL.t13 VSUBS 0.073227f
C211 VTAIL.n138 VSUBS 0.025521f
C212 VTAIL.n139 VSUBS 0.025598f
C213 VTAIL.n140 VSUBS 0.014396f
C214 VTAIL.n141 VSUBS 1.17193f
C215 VTAIL.n142 VSUBS 0.026791f
C216 VTAIL.n143 VSUBS 0.014396f
C217 VTAIL.n144 VSUBS 0.015243f
C218 VTAIL.n145 VSUBS 0.034028f
C219 VTAIL.n146 VSUBS 0.034028f
C220 VTAIL.n147 VSUBS 0.015243f
C221 VTAIL.n148 VSUBS 0.014396f
C222 VTAIL.n149 VSUBS 0.026791f
C223 VTAIL.n150 VSUBS 0.026791f
C224 VTAIL.n151 VSUBS 0.014396f
C225 VTAIL.n152 VSUBS 0.015243f
C226 VTAIL.n153 VSUBS 0.034028f
C227 VTAIL.n154 VSUBS 0.034028f
C228 VTAIL.n155 VSUBS 0.034028f
C229 VTAIL.n156 VSUBS 0.015243f
C230 VTAIL.n157 VSUBS 0.014396f
C231 VTAIL.n158 VSUBS 0.026791f
C232 VTAIL.n159 VSUBS 0.026791f
C233 VTAIL.n160 VSUBS 0.014396f
C234 VTAIL.n161 VSUBS 0.01482f
C235 VTAIL.n162 VSUBS 0.01482f
C236 VTAIL.n163 VSUBS 0.034028f
C237 VTAIL.n164 VSUBS 0.034028f
C238 VTAIL.n165 VSUBS 0.015243f
C239 VTAIL.n166 VSUBS 0.014396f
C240 VTAIL.n167 VSUBS 0.026791f
C241 VTAIL.n168 VSUBS 0.026791f
C242 VTAIL.n169 VSUBS 0.014396f
C243 VTAIL.n170 VSUBS 0.015243f
C244 VTAIL.n171 VSUBS 0.034028f
C245 VTAIL.n172 VSUBS 0.082383f
C246 VTAIL.n173 VSUBS 0.015243f
C247 VTAIL.n174 VSUBS 0.014396f
C248 VTAIL.n175 VSUBS 0.06522f
C249 VTAIL.n176 VSUBS 0.041529f
C250 VTAIL.n177 VSUBS 1.30627f
C251 VTAIL.n178 VSUBS 0.029439f
C252 VTAIL.n179 VSUBS 0.026791f
C253 VTAIL.n180 VSUBS 0.014396f
C254 VTAIL.n181 VSUBS 0.034028f
C255 VTAIL.n182 VSUBS 0.015243f
C256 VTAIL.n183 VSUBS 0.026791f
C257 VTAIL.n184 VSUBS 0.014396f
C258 VTAIL.n185 VSUBS 0.034028f
C259 VTAIL.n186 VSUBS 0.015243f
C260 VTAIL.n187 VSUBS 0.026791f
C261 VTAIL.n188 VSUBS 0.014396f
C262 VTAIL.n189 VSUBS 0.034028f
C263 VTAIL.n190 VSUBS 0.034028f
C264 VTAIL.n191 VSUBS 0.015243f
C265 VTAIL.n192 VSUBS 0.026791f
C266 VTAIL.n193 VSUBS 0.014396f
C267 VTAIL.n194 VSUBS 0.034028f
C268 VTAIL.n195 VSUBS 0.015243f
C269 VTAIL.n196 VSUBS 0.196107f
C270 VTAIL.t6 VSUBS 0.073227f
C271 VTAIL.n197 VSUBS 0.025521f
C272 VTAIL.n198 VSUBS 0.025598f
C273 VTAIL.n199 VSUBS 0.014396f
C274 VTAIL.n200 VSUBS 1.17193f
C275 VTAIL.n201 VSUBS 0.026791f
C276 VTAIL.n202 VSUBS 0.014396f
C277 VTAIL.n203 VSUBS 0.015243f
C278 VTAIL.n204 VSUBS 0.034028f
C279 VTAIL.n205 VSUBS 0.034028f
C280 VTAIL.n206 VSUBS 0.015243f
C281 VTAIL.n207 VSUBS 0.014396f
C282 VTAIL.n208 VSUBS 0.026791f
C283 VTAIL.n209 VSUBS 0.026791f
C284 VTAIL.n210 VSUBS 0.014396f
C285 VTAIL.n211 VSUBS 0.015243f
C286 VTAIL.n212 VSUBS 0.034028f
C287 VTAIL.n213 VSUBS 0.034028f
C288 VTAIL.n214 VSUBS 0.015243f
C289 VTAIL.n215 VSUBS 0.014396f
C290 VTAIL.n216 VSUBS 0.026791f
C291 VTAIL.n217 VSUBS 0.026791f
C292 VTAIL.n218 VSUBS 0.014396f
C293 VTAIL.n219 VSUBS 0.01482f
C294 VTAIL.n220 VSUBS 0.01482f
C295 VTAIL.n221 VSUBS 0.034028f
C296 VTAIL.n222 VSUBS 0.034028f
C297 VTAIL.n223 VSUBS 0.015243f
C298 VTAIL.n224 VSUBS 0.014396f
C299 VTAIL.n225 VSUBS 0.026791f
C300 VTAIL.n226 VSUBS 0.026791f
C301 VTAIL.n227 VSUBS 0.014396f
C302 VTAIL.n228 VSUBS 0.015243f
C303 VTAIL.n229 VSUBS 0.034028f
C304 VTAIL.n230 VSUBS 0.082383f
C305 VTAIL.n231 VSUBS 0.015243f
C306 VTAIL.n232 VSUBS 0.014396f
C307 VTAIL.n233 VSUBS 0.06522f
C308 VTAIL.n234 VSUBS 0.041529f
C309 VTAIL.n235 VSUBS 1.30627f
C310 VTAIL.t5 VSUBS 0.228014f
C311 VTAIL.t7 VSUBS 0.228014f
C312 VTAIL.n236 VSUBS 1.61944f
C313 VTAIL.n237 VSUBS 0.697999f
C314 VTAIL.n238 VSUBS 0.029439f
C315 VTAIL.n239 VSUBS 0.026791f
C316 VTAIL.n240 VSUBS 0.014396f
C317 VTAIL.n241 VSUBS 0.034028f
C318 VTAIL.n242 VSUBS 0.015243f
C319 VTAIL.n243 VSUBS 0.026791f
C320 VTAIL.n244 VSUBS 0.014396f
C321 VTAIL.n245 VSUBS 0.034028f
C322 VTAIL.n246 VSUBS 0.015243f
C323 VTAIL.n247 VSUBS 0.026791f
C324 VTAIL.n248 VSUBS 0.014396f
C325 VTAIL.n249 VSUBS 0.034028f
C326 VTAIL.n250 VSUBS 0.034028f
C327 VTAIL.n251 VSUBS 0.015243f
C328 VTAIL.n252 VSUBS 0.026791f
C329 VTAIL.n253 VSUBS 0.014396f
C330 VTAIL.n254 VSUBS 0.034028f
C331 VTAIL.n255 VSUBS 0.015243f
C332 VTAIL.n256 VSUBS 0.196107f
C333 VTAIL.t3 VSUBS 0.073227f
C334 VTAIL.n257 VSUBS 0.025521f
C335 VTAIL.n258 VSUBS 0.025598f
C336 VTAIL.n259 VSUBS 0.014396f
C337 VTAIL.n260 VSUBS 1.17193f
C338 VTAIL.n261 VSUBS 0.026791f
C339 VTAIL.n262 VSUBS 0.014396f
C340 VTAIL.n263 VSUBS 0.015243f
C341 VTAIL.n264 VSUBS 0.034028f
C342 VTAIL.n265 VSUBS 0.034028f
C343 VTAIL.n266 VSUBS 0.015243f
C344 VTAIL.n267 VSUBS 0.014396f
C345 VTAIL.n268 VSUBS 0.026791f
C346 VTAIL.n269 VSUBS 0.026791f
C347 VTAIL.n270 VSUBS 0.014396f
C348 VTAIL.n271 VSUBS 0.015243f
C349 VTAIL.n272 VSUBS 0.034028f
C350 VTAIL.n273 VSUBS 0.034028f
C351 VTAIL.n274 VSUBS 0.015243f
C352 VTAIL.n275 VSUBS 0.014396f
C353 VTAIL.n276 VSUBS 0.026791f
C354 VTAIL.n277 VSUBS 0.026791f
C355 VTAIL.n278 VSUBS 0.014396f
C356 VTAIL.n279 VSUBS 0.01482f
C357 VTAIL.n280 VSUBS 0.01482f
C358 VTAIL.n281 VSUBS 0.034028f
C359 VTAIL.n282 VSUBS 0.034028f
C360 VTAIL.n283 VSUBS 0.015243f
C361 VTAIL.n284 VSUBS 0.014396f
C362 VTAIL.n285 VSUBS 0.026791f
C363 VTAIL.n286 VSUBS 0.026791f
C364 VTAIL.n287 VSUBS 0.014396f
C365 VTAIL.n288 VSUBS 0.015243f
C366 VTAIL.n289 VSUBS 0.034028f
C367 VTAIL.n290 VSUBS 0.082383f
C368 VTAIL.n291 VSUBS 0.015243f
C369 VTAIL.n292 VSUBS 0.014396f
C370 VTAIL.n293 VSUBS 0.06522f
C371 VTAIL.n294 VSUBS 0.041529f
C372 VTAIL.n295 VSUBS 0.12335f
C373 VTAIL.n296 VSUBS 0.029439f
C374 VTAIL.n297 VSUBS 0.026791f
C375 VTAIL.n298 VSUBS 0.014396f
C376 VTAIL.n299 VSUBS 0.034028f
C377 VTAIL.n300 VSUBS 0.015243f
C378 VTAIL.n301 VSUBS 0.026791f
C379 VTAIL.n302 VSUBS 0.014396f
C380 VTAIL.n303 VSUBS 0.034028f
C381 VTAIL.n304 VSUBS 0.015243f
C382 VTAIL.n305 VSUBS 0.026791f
C383 VTAIL.n306 VSUBS 0.014396f
C384 VTAIL.n307 VSUBS 0.034028f
C385 VTAIL.n308 VSUBS 0.034028f
C386 VTAIL.n309 VSUBS 0.015243f
C387 VTAIL.n310 VSUBS 0.026791f
C388 VTAIL.n311 VSUBS 0.014396f
C389 VTAIL.n312 VSUBS 0.034028f
C390 VTAIL.n313 VSUBS 0.015243f
C391 VTAIL.n314 VSUBS 0.196107f
C392 VTAIL.t15 VSUBS 0.073227f
C393 VTAIL.n315 VSUBS 0.025521f
C394 VTAIL.n316 VSUBS 0.025598f
C395 VTAIL.n317 VSUBS 0.014396f
C396 VTAIL.n318 VSUBS 1.17193f
C397 VTAIL.n319 VSUBS 0.026791f
C398 VTAIL.n320 VSUBS 0.014396f
C399 VTAIL.n321 VSUBS 0.015243f
C400 VTAIL.n322 VSUBS 0.034028f
C401 VTAIL.n323 VSUBS 0.034028f
C402 VTAIL.n324 VSUBS 0.015243f
C403 VTAIL.n325 VSUBS 0.014396f
C404 VTAIL.n326 VSUBS 0.026791f
C405 VTAIL.n327 VSUBS 0.026791f
C406 VTAIL.n328 VSUBS 0.014396f
C407 VTAIL.n329 VSUBS 0.015243f
C408 VTAIL.n330 VSUBS 0.034028f
C409 VTAIL.n331 VSUBS 0.034028f
C410 VTAIL.n332 VSUBS 0.015243f
C411 VTAIL.n333 VSUBS 0.014396f
C412 VTAIL.n334 VSUBS 0.026791f
C413 VTAIL.n335 VSUBS 0.026791f
C414 VTAIL.n336 VSUBS 0.014396f
C415 VTAIL.n337 VSUBS 0.01482f
C416 VTAIL.n338 VSUBS 0.01482f
C417 VTAIL.n339 VSUBS 0.034028f
C418 VTAIL.n340 VSUBS 0.034028f
C419 VTAIL.n341 VSUBS 0.015243f
C420 VTAIL.n342 VSUBS 0.014396f
C421 VTAIL.n343 VSUBS 0.026791f
C422 VTAIL.n344 VSUBS 0.026791f
C423 VTAIL.n345 VSUBS 0.014396f
C424 VTAIL.n346 VSUBS 0.015243f
C425 VTAIL.n347 VSUBS 0.034028f
C426 VTAIL.n348 VSUBS 0.082383f
C427 VTAIL.n349 VSUBS 0.015243f
C428 VTAIL.n350 VSUBS 0.014396f
C429 VTAIL.n351 VSUBS 0.06522f
C430 VTAIL.n352 VSUBS 0.041529f
C431 VTAIL.n353 VSUBS 0.12335f
C432 VTAIL.t9 VSUBS 0.228014f
C433 VTAIL.t11 VSUBS 0.228014f
C434 VTAIL.n354 VSUBS 1.61944f
C435 VTAIL.n355 VSUBS 0.697999f
C436 VTAIL.n356 VSUBS 0.029439f
C437 VTAIL.n357 VSUBS 0.026791f
C438 VTAIL.n358 VSUBS 0.014396f
C439 VTAIL.n359 VSUBS 0.034028f
C440 VTAIL.n360 VSUBS 0.015243f
C441 VTAIL.n361 VSUBS 0.026791f
C442 VTAIL.n362 VSUBS 0.014396f
C443 VTAIL.n363 VSUBS 0.034028f
C444 VTAIL.n364 VSUBS 0.015243f
C445 VTAIL.n365 VSUBS 0.026791f
C446 VTAIL.n366 VSUBS 0.014396f
C447 VTAIL.n367 VSUBS 0.034028f
C448 VTAIL.n368 VSUBS 0.034028f
C449 VTAIL.n369 VSUBS 0.015243f
C450 VTAIL.n370 VSUBS 0.026791f
C451 VTAIL.n371 VSUBS 0.014396f
C452 VTAIL.n372 VSUBS 0.034028f
C453 VTAIL.n373 VSUBS 0.015243f
C454 VTAIL.n374 VSUBS 0.196107f
C455 VTAIL.t8 VSUBS 0.073227f
C456 VTAIL.n375 VSUBS 0.025521f
C457 VTAIL.n376 VSUBS 0.025598f
C458 VTAIL.n377 VSUBS 0.014396f
C459 VTAIL.n378 VSUBS 1.17193f
C460 VTAIL.n379 VSUBS 0.026791f
C461 VTAIL.n380 VSUBS 0.014396f
C462 VTAIL.n381 VSUBS 0.015243f
C463 VTAIL.n382 VSUBS 0.034028f
C464 VTAIL.n383 VSUBS 0.034028f
C465 VTAIL.n384 VSUBS 0.015243f
C466 VTAIL.n385 VSUBS 0.014396f
C467 VTAIL.n386 VSUBS 0.026791f
C468 VTAIL.n387 VSUBS 0.026791f
C469 VTAIL.n388 VSUBS 0.014396f
C470 VTAIL.n389 VSUBS 0.015243f
C471 VTAIL.n390 VSUBS 0.034028f
C472 VTAIL.n391 VSUBS 0.034028f
C473 VTAIL.n392 VSUBS 0.015243f
C474 VTAIL.n393 VSUBS 0.014396f
C475 VTAIL.n394 VSUBS 0.026791f
C476 VTAIL.n395 VSUBS 0.026791f
C477 VTAIL.n396 VSUBS 0.014396f
C478 VTAIL.n397 VSUBS 0.01482f
C479 VTAIL.n398 VSUBS 0.01482f
C480 VTAIL.n399 VSUBS 0.034028f
C481 VTAIL.n400 VSUBS 0.034028f
C482 VTAIL.n401 VSUBS 0.015243f
C483 VTAIL.n402 VSUBS 0.014396f
C484 VTAIL.n403 VSUBS 0.026791f
C485 VTAIL.n404 VSUBS 0.026791f
C486 VTAIL.n405 VSUBS 0.014396f
C487 VTAIL.n406 VSUBS 0.015243f
C488 VTAIL.n407 VSUBS 0.034028f
C489 VTAIL.n408 VSUBS 0.082383f
C490 VTAIL.n409 VSUBS 0.015243f
C491 VTAIL.n410 VSUBS 0.014396f
C492 VTAIL.n411 VSUBS 0.06522f
C493 VTAIL.n412 VSUBS 0.041529f
C494 VTAIL.n413 VSUBS 1.30627f
C495 VTAIL.n414 VSUBS 0.029439f
C496 VTAIL.n415 VSUBS 0.026791f
C497 VTAIL.n416 VSUBS 0.014396f
C498 VTAIL.n417 VSUBS 0.034028f
C499 VTAIL.n418 VSUBS 0.015243f
C500 VTAIL.n419 VSUBS 0.026791f
C501 VTAIL.n420 VSUBS 0.014396f
C502 VTAIL.n421 VSUBS 0.034028f
C503 VTAIL.n422 VSUBS 0.015243f
C504 VTAIL.n423 VSUBS 0.026791f
C505 VTAIL.n424 VSUBS 0.014396f
C506 VTAIL.n425 VSUBS 0.034028f
C507 VTAIL.n426 VSUBS 0.015243f
C508 VTAIL.n427 VSUBS 0.026791f
C509 VTAIL.n428 VSUBS 0.014396f
C510 VTAIL.n429 VSUBS 0.034028f
C511 VTAIL.n430 VSUBS 0.015243f
C512 VTAIL.n431 VSUBS 0.196107f
C513 VTAIL.t1 VSUBS 0.073227f
C514 VTAIL.n432 VSUBS 0.025521f
C515 VTAIL.n433 VSUBS 0.025598f
C516 VTAIL.n434 VSUBS 0.014396f
C517 VTAIL.n435 VSUBS 1.17193f
C518 VTAIL.n436 VSUBS 0.026791f
C519 VTAIL.n437 VSUBS 0.014396f
C520 VTAIL.n438 VSUBS 0.015243f
C521 VTAIL.n439 VSUBS 0.034028f
C522 VTAIL.n440 VSUBS 0.034028f
C523 VTAIL.n441 VSUBS 0.015243f
C524 VTAIL.n442 VSUBS 0.014396f
C525 VTAIL.n443 VSUBS 0.026791f
C526 VTAIL.n444 VSUBS 0.026791f
C527 VTAIL.n445 VSUBS 0.014396f
C528 VTAIL.n446 VSUBS 0.015243f
C529 VTAIL.n447 VSUBS 0.034028f
C530 VTAIL.n448 VSUBS 0.034028f
C531 VTAIL.n449 VSUBS 0.034028f
C532 VTAIL.n450 VSUBS 0.015243f
C533 VTAIL.n451 VSUBS 0.014396f
C534 VTAIL.n452 VSUBS 0.026791f
C535 VTAIL.n453 VSUBS 0.026791f
C536 VTAIL.n454 VSUBS 0.014396f
C537 VTAIL.n455 VSUBS 0.01482f
C538 VTAIL.n456 VSUBS 0.01482f
C539 VTAIL.n457 VSUBS 0.034028f
C540 VTAIL.n458 VSUBS 0.034028f
C541 VTAIL.n459 VSUBS 0.015243f
C542 VTAIL.n460 VSUBS 0.014396f
C543 VTAIL.n461 VSUBS 0.026791f
C544 VTAIL.n462 VSUBS 0.026791f
C545 VTAIL.n463 VSUBS 0.014396f
C546 VTAIL.n464 VSUBS 0.015243f
C547 VTAIL.n465 VSUBS 0.034028f
C548 VTAIL.n466 VSUBS 0.082383f
C549 VTAIL.n467 VSUBS 0.015243f
C550 VTAIL.n468 VSUBS 0.014396f
C551 VTAIL.n469 VSUBS 0.06522f
C552 VTAIL.n470 VSUBS 0.041529f
C553 VTAIL.n471 VSUBS 1.30125f
C554 VDD1.t0 VSUBS 0.254117f
C555 VDD1.t7 VSUBS 0.254117f
C556 VDD1.n0 VSUBS 1.95502f
C557 VDD1.t6 VSUBS 0.254117f
C558 VDD1.t2 VSUBS 0.254117f
C559 VDD1.n1 VSUBS 1.95403f
C560 VDD1.t5 VSUBS 0.254117f
C561 VDD1.t1 VSUBS 0.254117f
C562 VDD1.n2 VSUBS 1.95403f
C563 VDD1.n3 VSUBS 2.98569f
C564 VDD1.t4 VSUBS 0.254117f
C565 VDD1.t3 VSUBS 0.254117f
C566 VDD1.n4 VSUBS 1.95169f
C567 VDD1.n5 VSUBS 2.84834f
C568 VP.n0 VSUBS 0.064343f
C569 VP.t1 VSUBS 0.891225f
C570 VP.n1 VSUBS 0.374661f
C571 VP.n2 VSUBS 0.064343f
C572 VP.t7 VSUBS 0.891225f
C573 VP.t4 VSUBS 0.891225f
C574 VP.t6 VSUBS 0.891225f
C575 VP.n3 VSUBS 0.374661f
C576 VP.t0 VSUBS 0.902494f
C577 VP.n4 VSUBS 0.357313f
C578 VP.n5 VSUBS 0.204067f
C579 VP.n6 VSUBS 0.014601f
C580 VP.n7 VSUBS 0.374661f
C581 VP.n8 VSUBS 0.368116f
C582 VP.n9 VSUBS 2.4371f
C583 VP.t2 VSUBS 0.891225f
C584 VP.n10 VSUBS 0.368116f
C585 VP.n11 VSUBS 2.49503f
C586 VP.n12 VSUBS 0.064343f
C587 VP.n13 VSUBS 0.064343f
C588 VP.n14 VSUBS 0.014601f
C589 VP.t3 VSUBS 0.891225f
C590 VP.n15 VSUBS 0.374661f
C591 VP.t5 VSUBS 0.891225f
C592 VP.n16 VSUBS 0.368116f
C593 VP.n17 VSUBS 0.049863f
C594 B.n0 VSUBS 0.007575f
C595 B.n1 VSUBS 0.007575f
C596 B.n2 VSUBS 0.011204f
C597 B.n3 VSUBS 0.008586f
C598 B.n4 VSUBS 0.008586f
C599 B.n5 VSUBS 0.008586f
C600 B.n6 VSUBS 0.008586f
C601 B.n7 VSUBS 0.008586f
C602 B.n8 VSUBS 0.008586f
C603 B.n9 VSUBS 0.008586f
C604 B.n10 VSUBS 0.008586f
C605 B.n11 VSUBS 0.018676f
C606 B.n12 VSUBS 0.008586f
C607 B.n13 VSUBS 0.008586f
C608 B.n14 VSUBS 0.008586f
C609 B.n15 VSUBS 0.008586f
C610 B.n16 VSUBS 0.008586f
C611 B.n17 VSUBS 0.008586f
C612 B.n18 VSUBS 0.008586f
C613 B.n19 VSUBS 0.008586f
C614 B.n20 VSUBS 0.008586f
C615 B.n21 VSUBS 0.008586f
C616 B.n22 VSUBS 0.008586f
C617 B.n23 VSUBS 0.008586f
C618 B.n24 VSUBS 0.008586f
C619 B.n25 VSUBS 0.008586f
C620 B.n26 VSUBS 0.008586f
C621 B.n27 VSUBS 0.008586f
C622 B.n28 VSUBS 0.008586f
C623 B.n29 VSUBS 0.008586f
C624 B.n30 VSUBS 0.008081f
C625 B.n31 VSUBS 0.008586f
C626 B.t4 VSUBS 0.225818f
C627 B.t5 VSUBS 0.236656f
C628 B.t3 VSUBS 0.239768f
C629 B.n32 VSUBS 0.326687f
C630 B.n33 VSUBS 0.276413f
C631 B.n34 VSUBS 0.019892f
C632 B.n35 VSUBS 0.008586f
C633 B.n36 VSUBS 0.008586f
C634 B.n37 VSUBS 0.008586f
C635 B.n38 VSUBS 0.008586f
C636 B.t7 VSUBS 0.225821f
C637 B.t8 VSUBS 0.23666f
C638 B.t6 VSUBS 0.239768f
C639 B.n39 VSUBS 0.326683f
C640 B.n40 VSUBS 0.27641f
C641 B.n41 VSUBS 0.008586f
C642 B.n42 VSUBS 0.008586f
C643 B.n43 VSUBS 0.008586f
C644 B.n44 VSUBS 0.008586f
C645 B.n45 VSUBS 0.008586f
C646 B.n46 VSUBS 0.008586f
C647 B.n47 VSUBS 0.008586f
C648 B.n48 VSUBS 0.008586f
C649 B.n49 VSUBS 0.008586f
C650 B.n50 VSUBS 0.008586f
C651 B.n51 VSUBS 0.008586f
C652 B.n52 VSUBS 0.008586f
C653 B.n53 VSUBS 0.008586f
C654 B.n54 VSUBS 0.008586f
C655 B.n55 VSUBS 0.008586f
C656 B.n56 VSUBS 0.008586f
C657 B.n57 VSUBS 0.008586f
C658 B.n58 VSUBS 0.008586f
C659 B.n59 VSUBS 0.020211f
C660 B.n60 VSUBS 0.008586f
C661 B.n61 VSUBS 0.008586f
C662 B.n62 VSUBS 0.008586f
C663 B.n63 VSUBS 0.008586f
C664 B.n64 VSUBS 0.008586f
C665 B.n65 VSUBS 0.008586f
C666 B.n66 VSUBS 0.008586f
C667 B.n67 VSUBS 0.008586f
C668 B.n68 VSUBS 0.008586f
C669 B.n69 VSUBS 0.008586f
C670 B.n70 VSUBS 0.008586f
C671 B.n71 VSUBS 0.008586f
C672 B.n72 VSUBS 0.008586f
C673 B.n73 VSUBS 0.008586f
C674 B.n74 VSUBS 0.008586f
C675 B.n75 VSUBS 0.008586f
C676 B.n76 VSUBS 0.008586f
C677 B.n77 VSUBS 0.008586f
C678 B.n78 VSUBS 0.008586f
C679 B.n79 VSUBS 0.019743f
C680 B.n80 VSUBS 0.008586f
C681 B.n81 VSUBS 0.008586f
C682 B.n82 VSUBS 0.008586f
C683 B.n83 VSUBS 0.008586f
C684 B.n84 VSUBS 0.008586f
C685 B.n85 VSUBS 0.008586f
C686 B.n86 VSUBS 0.008586f
C687 B.n87 VSUBS 0.008586f
C688 B.n88 VSUBS 0.008586f
C689 B.n89 VSUBS 0.008586f
C690 B.n90 VSUBS 0.008586f
C691 B.n91 VSUBS 0.008586f
C692 B.n92 VSUBS 0.008586f
C693 B.n93 VSUBS 0.008586f
C694 B.n94 VSUBS 0.008586f
C695 B.n95 VSUBS 0.008586f
C696 B.n96 VSUBS 0.008586f
C697 B.n97 VSUBS 0.008586f
C698 B.n98 VSUBS 0.008586f
C699 B.t2 VSUBS 0.225821f
C700 B.t1 VSUBS 0.23666f
C701 B.t0 VSUBS 0.239768f
C702 B.n99 VSUBS 0.326683f
C703 B.n100 VSUBS 0.27641f
C704 B.n101 VSUBS 0.008586f
C705 B.n102 VSUBS 0.008586f
C706 B.n103 VSUBS 0.008586f
C707 B.n104 VSUBS 0.008586f
C708 B.n105 VSUBS 0.004798f
C709 B.n106 VSUBS 0.008586f
C710 B.n107 VSUBS 0.008586f
C711 B.n108 VSUBS 0.008586f
C712 B.n109 VSUBS 0.008586f
C713 B.n110 VSUBS 0.008586f
C714 B.n111 VSUBS 0.008586f
C715 B.n112 VSUBS 0.008586f
C716 B.n113 VSUBS 0.008586f
C717 B.n114 VSUBS 0.008586f
C718 B.n115 VSUBS 0.008586f
C719 B.n116 VSUBS 0.008586f
C720 B.n117 VSUBS 0.008586f
C721 B.n118 VSUBS 0.008586f
C722 B.n119 VSUBS 0.008586f
C723 B.n120 VSUBS 0.008586f
C724 B.n121 VSUBS 0.008586f
C725 B.n122 VSUBS 0.008586f
C726 B.n123 VSUBS 0.008586f
C727 B.n124 VSUBS 0.020211f
C728 B.n125 VSUBS 0.008586f
C729 B.n126 VSUBS 0.008586f
C730 B.n127 VSUBS 0.008586f
C731 B.n128 VSUBS 0.008586f
C732 B.n129 VSUBS 0.008586f
C733 B.n130 VSUBS 0.008586f
C734 B.n131 VSUBS 0.008586f
C735 B.n132 VSUBS 0.008586f
C736 B.n133 VSUBS 0.008586f
C737 B.n134 VSUBS 0.008586f
C738 B.n135 VSUBS 0.008586f
C739 B.n136 VSUBS 0.008586f
C740 B.n137 VSUBS 0.008586f
C741 B.n138 VSUBS 0.008586f
C742 B.n139 VSUBS 0.008586f
C743 B.n140 VSUBS 0.008586f
C744 B.n141 VSUBS 0.008586f
C745 B.n142 VSUBS 0.008586f
C746 B.n143 VSUBS 0.008586f
C747 B.n144 VSUBS 0.008586f
C748 B.n145 VSUBS 0.008586f
C749 B.n146 VSUBS 0.008586f
C750 B.n147 VSUBS 0.008586f
C751 B.n148 VSUBS 0.008586f
C752 B.n149 VSUBS 0.008586f
C753 B.n150 VSUBS 0.008586f
C754 B.n151 VSUBS 0.008586f
C755 B.n152 VSUBS 0.008586f
C756 B.n153 VSUBS 0.008586f
C757 B.n154 VSUBS 0.008586f
C758 B.n155 VSUBS 0.008586f
C759 B.n156 VSUBS 0.008586f
C760 B.n157 VSUBS 0.008586f
C761 B.n158 VSUBS 0.008586f
C762 B.n159 VSUBS 0.018676f
C763 B.n160 VSUBS 0.018676f
C764 B.n161 VSUBS 0.020211f
C765 B.n162 VSUBS 0.008586f
C766 B.n163 VSUBS 0.008586f
C767 B.n164 VSUBS 0.008586f
C768 B.n165 VSUBS 0.008586f
C769 B.n166 VSUBS 0.008586f
C770 B.n167 VSUBS 0.008586f
C771 B.n168 VSUBS 0.008586f
C772 B.n169 VSUBS 0.008586f
C773 B.n170 VSUBS 0.008586f
C774 B.n171 VSUBS 0.008586f
C775 B.n172 VSUBS 0.008586f
C776 B.n173 VSUBS 0.008586f
C777 B.n174 VSUBS 0.008586f
C778 B.n175 VSUBS 0.008586f
C779 B.n176 VSUBS 0.008586f
C780 B.n177 VSUBS 0.008586f
C781 B.n178 VSUBS 0.008586f
C782 B.n179 VSUBS 0.008586f
C783 B.n180 VSUBS 0.008586f
C784 B.n181 VSUBS 0.008586f
C785 B.n182 VSUBS 0.008586f
C786 B.n183 VSUBS 0.008586f
C787 B.n184 VSUBS 0.008586f
C788 B.n185 VSUBS 0.008586f
C789 B.n186 VSUBS 0.008586f
C790 B.n187 VSUBS 0.008586f
C791 B.n188 VSUBS 0.008586f
C792 B.n189 VSUBS 0.008586f
C793 B.n190 VSUBS 0.008586f
C794 B.n191 VSUBS 0.008586f
C795 B.n192 VSUBS 0.008586f
C796 B.n193 VSUBS 0.008586f
C797 B.n194 VSUBS 0.008586f
C798 B.n195 VSUBS 0.008586f
C799 B.n196 VSUBS 0.008586f
C800 B.n197 VSUBS 0.008586f
C801 B.n198 VSUBS 0.008586f
C802 B.n199 VSUBS 0.008586f
C803 B.n200 VSUBS 0.008586f
C804 B.n201 VSUBS 0.008586f
C805 B.n202 VSUBS 0.008586f
C806 B.n203 VSUBS 0.008586f
C807 B.n204 VSUBS 0.008586f
C808 B.n205 VSUBS 0.008586f
C809 B.n206 VSUBS 0.008586f
C810 B.n207 VSUBS 0.008586f
C811 B.n208 VSUBS 0.008586f
C812 B.n209 VSUBS 0.008586f
C813 B.n210 VSUBS 0.008586f
C814 B.n211 VSUBS 0.008586f
C815 B.n212 VSUBS 0.008586f
C816 B.n213 VSUBS 0.008586f
C817 B.n214 VSUBS 0.008586f
C818 B.n215 VSUBS 0.008586f
C819 B.t11 VSUBS 0.225818f
C820 B.t10 VSUBS 0.236656f
C821 B.t9 VSUBS 0.239768f
C822 B.n216 VSUBS 0.326687f
C823 B.n217 VSUBS 0.276413f
C824 B.n218 VSUBS 0.019892f
C825 B.n219 VSUBS 0.008081f
C826 B.n220 VSUBS 0.008586f
C827 B.n221 VSUBS 0.008586f
C828 B.n222 VSUBS 0.008586f
C829 B.n223 VSUBS 0.008586f
C830 B.n224 VSUBS 0.008586f
C831 B.n225 VSUBS 0.008586f
C832 B.n226 VSUBS 0.008586f
C833 B.n227 VSUBS 0.008586f
C834 B.n228 VSUBS 0.008586f
C835 B.n229 VSUBS 0.008586f
C836 B.n230 VSUBS 0.008586f
C837 B.n231 VSUBS 0.008586f
C838 B.n232 VSUBS 0.008586f
C839 B.n233 VSUBS 0.008586f
C840 B.n234 VSUBS 0.008586f
C841 B.n235 VSUBS 0.004798f
C842 B.n236 VSUBS 0.019892f
C843 B.n237 VSUBS 0.008081f
C844 B.n238 VSUBS 0.008586f
C845 B.n239 VSUBS 0.008586f
C846 B.n240 VSUBS 0.008586f
C847 B.n241 VSUBS 0.008586f
C848 B.n242 VSUBS 0.008586f
C849 B.n243 VSUBS 0.008586f
C850 B.n244 VSUBS 0.008586f
C851 B.n245 VSUBS 0.008586f
C852 B.n246 VSUBS 0.008586f
C853 B.n247 VSUBS 0.008586f
C854 B.n248 VSUBS 0.008586f
C855 B.n249 VSUBS 0.008586f
C856 B.n250 VSUBS 0.008586f
C857 B.n251 VSUBS 0.008586f
C858 B.n252 VSUBS 0.008586f
C859 B.n253 VSUBS 0.008586f
C860 B.n254 VSUBS 0.008586f
C861 B.n255 VSUBS 0.008586f
C862 B.n256 VSUBS 0.008586f
C863 B.n257 VSUBS 0.008586f
C864 B.n258 VSUBS 0.008586f
C865 B.n259 VSUBS 0.008586f
C866 B.n260 VSUBS 0.008586f
C867 B.n261 VSUBS 0.008586f
C868 B.n262 VSUBS 0.008586f
C869 B.n263 VSUBS 0.008586f
C870 B.n264 VSUBS 0.008586f
C871 B.n265 VSUBS 0.008586f
C872 B.n266 VSUBS 0.008586f
C873 B.n267 VSUBS 0.008586f
C874 B.n268 VSUBS 0.008586f
C875 B.n269 VSUBS 0.008586f
C876 B.n270 VSUBS 0.008586f
C877 B.n271 VSUBS 0.008586f
C878 B.n272 VSUBS 0.008586f
C879 B.n273 VSUBS 0.008586f
C880 B.n274 VSUBS 0.008586f
C881 B.n275 VSUBS 0.008586f
C882 B.n276 VSUBS 0.008586f
C883 B.n277 VSUBS 0.008586f
C884 B.n278 VSUBS 0.008586f
C885 B.n279 VSUBS 0.008586f
C886 B.n280 VSUBS 0.008586f
C887 B.n281 VSUBS 0.008586f
C888 B.n282 VSUBS 0.008586f
C889 B.n283 VSUBS 0.008586f
C890 B.n284 VSUBS 0.008586f
C891 B.n285 VSUBS 0.008586f
C892 B.n286 VSUBS 0.008586f
C893 B.n287 VSUBS 0.008586f
C894 B.n288 VSUBS 0.008586f
C895 B.n289 VSUBS 0.008586f
C896 B.n290 VSUBS 0.008586f
C897 B.n291 VSUBS 0.008586f
C898 B.n292 VSUBS 0.019145f
C899 B.n293 VSUBS 0.020211f
C900 B.n294 VSUBS 0.018676f
C901 B.n295 VSUBS 0.008586f
C902 B.n296 VSUBS 0.008586f
C903 B.n297 VSUBS 0.008586f
C904 B.n298 VSUBS 0.008586f
C905 B.n299 VSUBS 0.008586f
C906 B.n300 VSUBS 0.008586f
C907 B.n301 VSUBS 0.008586f
C908 B.n302 VSUBS 0.008586f
C909 B.n303 VSUBS 0.008586f
C910 B.n304 VSUBS 0.008586f
C911 B.n305 VSUBS 0.008586f
C912 B.n306 VSUBS 0.008586f
C913 B.n307 VSUBS 0.008586f
C914 B.n308 VSUBS 0.008586f
C915 B.n309 VSUBS 0.008586f
C916 B.n310 VSUBS 0.008586f
C917 B.n311 VSUBS 0.008586f
C918 B.n312 VSUBS 0.008586f
C919 B.n313 VSUBS 0.008586f
C920 B.n314 VSUBS 0.008586f
C921 B.n315 VSUBS 0.008586f
C922 B.n316 VSUBS 0.008586f
C923 B.n317 VSUBS 0.008586f
C924 B.n318 VSUBS 0.008586f
C925 B.n319 VSUBS 0.008586f
C926 B.n320 VSUBS 0.008586f
C927 B.n321 VSUBS 0.008586f
C928 B.n322 VSUBS 0.008586f
C929 B.n323 VSUBS 0.008586f
C930 B.n324 VSUBS 0.008586f
C931 B.n325 VSUBS 0.008586f
C932 B.n326 VSUBS 0.008586f
C933 B.n327 VSUBS 0.008586f
C934 B.n328 VSUBS 0.008586f
C935 B.n329 VSUBS 0.008586f
C936 B.n330 VSUBS 0.008586f
C937 B.n331 VSUBS 0.008586f
C938 B.n332 VSUBS 0.008586f
C939 B.n333 VSUBS 0.008586f
C940 B.n334 VSUBS 0.008586f
C941 B.n335 VSUBS 0.008586f
C942 B.n336 VSUBS 0.008586f
C943 B.n337 VSUBS 0.008586f
C944 B.n338 VSUBS 0.008586f
C945 B.n339 VSUBS 0.008586f
C946 B.n340 VSUBS 0.008586f
C947 B.n341 VSUBS 0.008586f
C948 B.n342 VSUBS 0.008586f
C949 B.n343 VSUBS 0.008586f
C950 B.n344 VSUBS 0.008586f
C951 B.n345 VSUBS 0.008586f
C952 B.n346 VSUBS 0.008586f
C953 B.n347 VSUBS 0.008586f
C954 B.n348 VSUBS 0.008586f
C955 B.n349 VSUBS 0.008586f
C956 B.n350 VSUBS 0.008586f
C957 B.n351 VSUBS 0.008586f
C958 B.n352 VSUBS 0.018676f
C959 B.n353 VSUBS 0.018676f
C960 B.n354 VSUBS 0.020211f
C961 B.n355 VSUBS 0.008586f
C962 B.n356 VSUBS 0.008586f
C963 B.n357 VSUBS 0.008586f
C964 B.n358 VSUBS 0.008586f
C965 B.n359 VSUBS 0.008586f
C966 B.n360 VSUBS 0.008586f
C967 B.n361 VSUBS 0.008586f
C968 B.n362 VSUBS 0.008586f
C969 B.n363 VSUBS 0.008586f
C970 B.n364 VSUBS 0.008586f
C971 B.n365 VSUBS 0.008586f
C972 B.n366 VSUBS 0.008586f
C973 B.n367 VSUBS 0.008586f
C974 B.n368 VSUBS 0.008586f
C975 B.n369 VSUBS 0.008586f
C976 B.n370 VSUBS 0.008586f
C977 B.n371 VSUBS 0.008586f
C978 B.n372 VSUBS 0.008586f
C979 B.n373 VSUBS 0.008586f
C980 B.n374 VSUBS 0.008586f
C981 B.n375 VSUBS 0.008586f
C982 B.n376 VSUBS 0.008586f
C983 B.n377 VSUBS 0.008586f
C984 B.n378 VSUBS 0.008586f
C985 B.n379 VSUBS 0.008586f
C986 B.n380 VSUBS 0.008586f
C987 B.n381 VSUBS 0.008586f
C988 B.n382 VSUBS 0.008586f
C989 B.n383 VSUBS 0.008586f
C990 B.n384 VSUBS 0.008586f
C991 B.n385 VSUBS 0.008586f
C992 B.n386 VSUBS 0.008586f
C993 B.n387 VSUBS 0.008586f
C994 B.n388 VSUBS 0.008586f
C995 B.n389 VSUBS 0.008586f
C996 B.n390 VSUBS 0.008586f
C997 B.n391 VSUBS 0.008586f
C998 B.n392 VSUBS 0.008586f
C999 B.n393 VSUBS 0.008586f
C1000 B.n394 VSUBS 0.008586f
C1001 B.n395 VSUBS 0.008586f
C1002 B.n396 VSUBS 0.008586f
C1003 B.n397 VSUBS 0.008586f
C1004 B.n398 VSUBS 0.008586f
C1005 B.n399 VSUBS 0.008586f
C1006 B.n400 VSUBS 0.008586f
C1007 B.n401 VSUBS 0.008586f
C1008 B.n402 VSUBS 0.008586f
C1009 B.n403 VSUBS 0.008586f
C1010 B.n404 VSUBS 0.008586f
C1011 B.n405 VSUBS 0.008586f
C1012 B.n406 VSUBS 0.008586f
C1013 B.n407 VSUBS 0.008586f
C1014 B.n408 VSUBS 0.008586f
C1015 B.n409 VSUBS 0.008586f
C1016 B.n410 VSUBS 0.008081f
C1017 B.n411 VSUBS 0.019892f
C1018 B.n412 VSUBS 0.004798f
C1019 B.n413 VSUBS 0.008586f
C1020 B.n414 VSUBS 0.008586f
C1021 B.n415 VSUBS 0.008586f
C1022 B.n416 VSUBS 0.008586f
C1023 B.n417 VSUBS 0.008586f
C1024 B.n418 VSUBS 0.008586f
C1025 B.n419 VSUBS 0.008586f
C1026 B.n420 VSUBS 0.008586f
C1027 B.n421 VSUBS 0.008586f
C1028 B.n422 VSUBS 0.008586f
C1029 B.n423 VSUBS 0.008586f
C1030 B.n424 VSUBS 0.008586f
C1031 B.n425 VSUBS 0.004798f
C1032 B.n426 VSUBS 0.008586f
C1033 B.n427 VSUBS 0.008586f
C1034 B.n428 VSUBS 0.008586f
C1035 B.n429 VSUBS 0.008586f
C1036 B.n430 VSUBS 0.008586f
C1037 B.n431 VSUBS 0.008586f
C1038 B.n432 VSUBS 0.008586f
C1039 B.n433 VSUBS 0.008586f
C1040 B.n434 VSUBS 0.008586f
C1041 B.n435 VSUBS 0.008586f
C1042 B.n436 VSUBS 0.008586f
C1043 B.n437 VSUBS 0.008586f
C1044 B.n438 VSUBS 0.008586f
C1045 B.n439 VSUBS 0.008586f
C1046 B.n440 VSUBS 0.008586f
C1047 B.n441 VSUBS 0.008586f
C1048 B.n442 VSUBS 0.008586f
C1049 B.n443 VSUBS 0.008586f
C1050 B.n444 VSUBS 0.008586f
C1051 B.n445 VSUBS 0.008586f
C1052 B.n446 VSUBS 0.008586f
C1053 B.n447 VSUBS 0.008586f
C1054 B.n448 VSUBS 0.008586f
C1055 B.n449 VSUBS 0.008586f
C1056 B.n450 VSUBS 0.008586f
C1057 B.n451 VSUBS 0.008586f
C1058 B.n452 VSUBS 0.008586f
C1059 B.n453 VSUBS 0.008586f
C1060 B.n454 VSUBS 0.008586f
C1061 B.n455 VSUBS 0.008586f
C1062 B.n456 VSUBS 0.008586f
C1063 B.n457 VSUBS 0.008586f
C1064 B.n458 VSUBS 0.008586f
C1065 B.n459 VSUBS 0.008586f
C1066 B.n460 VSUBS 0.008586f
C1067 B.n461 VSUBS 0.008586f
C1068 B.n462 VSUBS 0.008586f
C1069 B.n463 VSUBS 0.008586f
C1070 B.n464 VSUBS 0.008586f
C1071 B.n465 VSUBS 0.008586f
C1072 B.n466 VSUBS 0.008586f
C1073 B.n467 VSUBS 0.008586f
C1074 B.n468 VSUBS 0.008586f
C1075 B.n469 VSUBS 0.008586f
C1076 B.n470 VSUBS 0.008586f
C1077 B.n471 VSUBS 0.008586f
C1078 B.n472 VSUBS 0.008586f
C1079 B.n473 VSUBS 0.008586f
C1080 B.n474 VSUBS 0.008586f
C1081 B.n475 VSUBS 0.008586f
C1082 B.n476 VSUBS 0.008586f
C1083 B.n477 VSUBS 0.008586f
C1084 B.n478 VSUBS 0.008586f
C1085 B.n479 VSUBS 0.008586f
C1086 B.n480 VSUBS 0.008586f
C1087 B.n481 VSUBS 0.008586f
C1088 B.n482 VSUBS 0.020211f
C1089 B.n483 VSUBS 0.020211f
C1090 B.n484 VSUBS 0.018676f
C1091 B.n485 VSUBS 0.008586f
C1092 B.n486 VSUBS 0.008586f
C1093 B.n487 VSUBS 0.008586f
C1094 B.n488 VSUBS 0.008586f
C1095 B.n489 VSUBS 0.008586f
C1096 B.n490 VSUBS 0.008586f
C1097 B.n491 VSUBS 0.008586f
C1098 B.n492 VSUBS 0.008586f
C1099 B.n493 VSUBS 0.008586f
C1100 B.n494 VSUBS 0.008586f
C1101 B.n495 VSUBS 0.008586f
C1102 B.n496 VSUBS 0.008586f
C1103 B.n497 VSUBS 0.008586f
C1104 B.n498 VSUBS 0.008586f
C1105 B.n499 VSUBS 0.008586f
C1106 B.n500 VSUBS 0.008586f
C1107 B.n501 VSUBS 0.008586f
C1108 B.n502 VSUBS 0.008586f
C1109 B.n503 VSUBS 0.008586f
C1110 B.n504 VSUBS 0.008586f
C1111 B.n505 VSUBS 0.008586f
C1112 B.n506 VSUBS 0.008586f
C1113 B.n507 VSUBS 0.008586f
C1114 B.n508 VSUBS 0.008586f
C1115 B.n509 VSUBS 0.008586f
C1116 B.n510 VSUBS 0.008586f
C1117 B.n511 VSUBS 0.011204f
C1118 B.n512 VSUBS 0.011935f
C1119 B.n513 VSUBS 0.023733f
.ends

