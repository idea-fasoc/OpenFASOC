* NGSPICE file created from diff_pair_sample_0651.ext - technology: sky130A

.subckt diff_pair_sample_0651 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=2.8509 ps=15.4 w=7.31 l=0.28
X1 B.t11 B.t9 B.t10 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=0.28
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=2.8509 ps=15.4 w=7.31 l=0.28
X3 B.t8 B.t6 B.t7 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=0.28
X4 B.t5 B.t3 B.t4 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=0.28
X5 VDD2.t0 VN.t1 VTAIL.t3 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=2.8509 ps=15.4 w=7.31 l=0.28
X6 B.t2 B.t0 B.t1 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=0 ps=0 w=7.31 l=0.28
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1214_n2434# sky130_fd_pr__pfet_01v8 ad=2.8509 pd=15.4 as=2.8509 ps=15.4 w=7.31 l=0.28
R0 VN VN.t1 962.683
R1 VN VN.t0 927.388
R2 VTAIL.n121 VTAIL.n120 585
R3 VTAIL.n123 VTAIL.n122 585
R4 VTAIL.n116 VTAIL.n115 585
R5 VTAIL.n129 VTAIL.n128 585
R6 VTAIL.n131 VTAIL.n130 585
R7 VTAIL.n112 VTAIL.n111 585
R8 VTAIL.n137 VTAIL.n136 585
R9 VTAIL.n139 VTAIL.n138 585
R10 VTAIL.n13 VTAIL.n12 585
R11 VTAIL.n15 VTAIL.n14 585
R12 VTAIL.n8 VTAIL.n7 585
R13 VTAIL.n21 VTAIL.n20 585
R14 VTAIL.n23 VTAIL.n22 585
R15 VTAIL.n4 VTAIL.n3 585
R16 VTAIL.n29 VTAIL.n28 585
R17 VTAIL.n31 VTAIL.n30 585
R18 VTAIL.n103 VTAIL.n102 585
R19 VTAIL.n101 VTAIL.n100 585
R20 VTAIL.n76 VTAIL.n75 585
R21 VTAIL.n95 VTAIL.n94 585
R22 VTAIL.n93 VTAIL.n92 585
R23 VTAIL.n80 VTAIL.n79 585
R24 VTAIL.n87 VTAIL.n86 585
R25 VTAIL.n85 VTAIL.n84 585
R26 VTAIL.n67 VTAIL.n66 585
R27 VTAIL.n65 VTAIL.n64 585
R28 VTAIL.n40 VTAIL.n39 585
R29 VTAIL.n59 VTAIL.n58 585
R30 VTAIL.n57 VTAIL.n56 585
R31 VTAIL.n44 VTAIL.n43 585
R32 VTAIL.n51 VTAIL.n50 585
R33 VTAIL.n49 VTAIL.n48 585
R34 VTAIL.n138 VTAIL.n108 498.474
R35 VTAIL.n30 VTAIL.n0 498.474
R36 VTAIL.n102 VTAIL.n72 498.474
R37 VTAIL.n66 VTAIL.n36 498.474
R38 VTAIL.n119 VTAIL.t2 329.053
R39 VTAIL.n11 VTAIL.t0 329.053
R40 VTAIL.n83 VTAIL.t1 329.053
R41 VTAIL.n47 VTAIL.t3 329.053
R42 VTAIL.n122 VTAIL.n121 171.744
R43 VTAIL.n122 VTAIL.n115 171.744
R44 VTAIL.n129 VTAIL.n115 171.744
R45 VTAIL.n130 VTAIL.n129 171.744
R46 VTAIL.n130 VTAIL.n111 171.744
R47 VTAIL.n137 VTAIL.n111 171.744
R48 VTAIL.n138 VTAIL.n137 171.744
R49 VTAIL.n14 VTAIL.n13 171.744
R50 VTAIL.n14 VTAIL.n7 171.744
R51 VTAIL.n21 VTAIL.n7 171.744
R52 VTAIL.n22 VTAIL.n21 171.744
R53 VTAIL.n22 VTAIL.n3 171.744
R54 VTAIL.n29 VTAIL.n3 171.744
R55 VTAIL.n30 VTAIL.n29 171.744
R56 VTAIL.n102 VTAIL.n101 171.744
R57 VTAIL.n101 VTAIL.n75 171.744
R58 VTAIL.n94 VTAIL.n75 171.744
R59 VTAIL.n94 VTAIL.n93 171.744
R60 VTAIL.n93 VTAIL.n79 171.744
R61 VTAIL.n86 VTAIL.n79 171.744
R62 VTAIL.n86 VTAIL.n85 171.744
R63 VTAIL.n66 VTAIL.n65 171.744
R64 VTAIL.n65 VTAIL.n39 171.744
R65 VTAIL.n58 VTAIL.n39 171.744
R66 VTAIL.n58 VTAIL.n57 171.744
R67 VTAIL.n57 VTAIL.n43 171.744
R68 VTAIL.n50 VTAIL.n43 171.744
R69 VTAIL.n50 VTAIL.n49 171.744
R70 VTAIL.n121 VTAIL.t2 85.8723
R71 VTAIL.n13 VTAIL.t0 85.8723
R72 VTAIL.n85 VTAIL.t1 85.8723
R73 VTAIL.n49 VTAIL.t3 85.8723
R74 VTAIL.n143 VTAIL.n142 36.646
R75 VTAIL.n35 VTAIL.n34 36.646
R76 VTAIL.n107 VTAIL.n106 36.646
R77 VTAIL.n71 VTAIL.n70 36.646
R78 VTAIL.n71 VTAIL.n35 19.7376
R79 VTAIL.n143 VTAIL.n107 19.2117
R80 VTAIL.n140 VTAIL.n139 12.8005
R81 VTAIL.n32 VTAIL.n31 12.8005
R82 VTAIL.n104 VTAIL.n103 12.8005
R83 VTAIL.n68 VTAIL.n67 12.8005
R84 VTAIL.n136 VTAIL.n110 12.0247
R85 VTAIL.n28 VTAIL.n2 12.0247
R86 VTAIL.n100 VTAIL.n74 12.0247
R87 VTAIL.n64 VTAIL.n38 12.0247
R88 VTAIL.n135 VTAIL.n112 11.249
R89 VTAIL.n27 VTAIL.n4 11.249
R90 VTAIL.n99 VTAIL.n76 11.249
R91 VTAIL.n63 VTAIL.n40 11.249
R92 VTAIL.n120 VTAIL.n119 10.7237
R93 VTAIL.n12 VTAIL.n11 10.7237
R94 VTAIL.n84 VTAIL.n83 10.7237
R95 VTAIL.n48 VTAIL.n47 10.7237
R96 VTAIL.n132 VTAIL.n131 10.4732
R97 VTAIL.n24 VTAIL.n23 10.4732
R98 VTAIL.n96 VTAIL.n95 10.4732
R99 VTAIL.n60 VTAIL.n59 10.4732
R100 VTAIL.n128 VTAIL.n114 9.69747
R101 VTAIL.n20 VTAIL.n6 9.69747
R102 VTAIL.n92 VTAIL.n78 9.69747
R103 VTAIL.n56 VTAIL.n42 9.69747
R104 VTAIL.n142 VTAIL.n141 9.45567
R105 VTAIL.n34 VTAIL.n33 9.45567
R106 VTAIL.n106 VTAIL.n105 9.45567
R107 VTAIL.n70 VTAIL.n69 9.45567
R108 VTAIL.n118 VTAIL.n117 9.3005
R109 VTAIL.n125 VTAIL.n124 9.3005
R110 VTAIL.n127 VTAIL.n126 9.3005
R111 VTAIL.n114 VTAIL.n113 9.3005
R112 VTAIL.n133 VTAIL.n132 9.3005
R113 VTAIL.n135 VTAIL.n134 9.3005
R114 VTAIL.n110 VTAIL.n109 9.3005
R115 VTAIL.n141 VTAIL.n140 9.3005
R116 VTAIL.n10 VTAIL.n9 9.3005
R117 VTAIL.n17 VTAIL.n16 9.3005
R118 VTAIL.n19 VTAIL.n18 9.3005
R119 VTAIL.n6 VTAIL.n5 9.3005
R120 VTAIL.n25 VTAIL.n24 9.3005
R121 VTAIL.n27 VTAIL.n26 9.3005
R122 VTAIL.n2 VTAIL.n1 9.3005
R123 VTAIL.n33 VTAIL.n32 9.3005
R124 VTAIL.n82 VTAIL.n81 9.3005
R125 VTAIL.n89 VTAIL.n88 9.3005
R126 VTAIL.n91 VTAIL.n90 9.3005
R127 VTAIL.n78 VTAIL.n77 9.3005
R128 VTAIL.n97 VTAIL.n96 9.3005
R129 VTAIL.n99 VTAIL.n98 9.3005
R130 VTAIL.n74 VTAIL.n73 9.3005
R131 VTAIL.n105 VTAIL.n104 9.3005
R132 VTAIL.n46 VTAIL.n45 9.3005
R133 VTAIL.n53 VTAIL.n52 9.3005
R134 VTAIL.n55 VTAIL.n54 9.3005
R135 VTAIL.n42 VTAIL.n41 9.3005
R136 VTAIL.n61 VTAIL.n60 9.3005
R137 VTAIL.n63 VTAIL.n62 9.3005
R138 VTAIL.n38 VTAIL.n37 9.3005
R139 VTAIL.n69 VTAIL.n68 9.3005
R140 VTAIL.n127 VTAIL.n116 8.92171
R141 VTAIL.n19 VTAIL.n8 8.92171
R142 VTAIL.n91 VTAIL.n80 8.92171
R143 VTAIL.n55 VTAIL.n44 8.92171
R144 VTAIL.n124 VTAIL.n123 8.14595
R145 VTAIL.n16 VTAIL.n15 8.14595
R146 VTAIL.n88 VTAIL.n87 8.14595
R147 VTAIL.n52 VTAIL.n51 8.14595
R148 VTAIL.n142 VTAIL.n108 7.75445
R149 VTAIL.n34 VTAIL.n0 7.75445
R150 VTAIL.n106 VTAIL.n72 7.75445
R151 VTAIL.n70 VTAIL.n36 7.75445
R152 VTAIL.n120 VTAIL.n118 7.3702
R153 VTAIL.n12 VTAIL.n10 7.3702
R154 VTAIL.n84 VTAIL.n82 7.3702
R155 VTAIL.n48 VTAIL.n46 7.3702
R156 VTAIL.n140 VTAIL.n108 6.08283
R157 VTAIL.n32 VTAIL.n0 6.08283
R158 VTAIL.n104 VTAIL.n72 6.08283
R159 VTAIL.n68 VTAIL.n36 6.08283
R160 VTAIL.n123 VTAIL.n118 5.81868
R161 VTAIL.n15 VTAIL.n10 5.81868
R162 VTAIL.n87 VTAIL.n82 5.81868
R163 VTAIL.n51 VTAIL.n46 5.81868
R164 VTAIL.n124 VTAIL.n116 5.04292
R165 VTAIL.n16 VTAIL.n8 5.04292
R166 VTAIL.n88 VTAIL.n80 5.04292
R167 VTAIL.n52 VTAIL.n44 5.04292
R168 VTAIL.n128 VTAIL.n127 4.26717
R169 VTAIL.n20 VTAIL.n19 4.26717
R170 VTAIL.n92 VTAIL.n91 4.26717
R171 VTAIL.n56 VTAIL.n55 4.26717
R172 VTAIL.n131 VTAIL.n114 3.49141
R173 VTAIL.n23 VTAIL.n6 3.49141
R174 VTAIL.n95 VTAIL.n78 3.49141
R175 VTAIL.n59 VTAIL.n42 3.49141
R176 VTAIL.n132 VTAIL.n112 2.71565
R177 VTAIL.n24 VTAIL.n4 2.71565
R178 VTAIL.n96 VTAIL.n76 2.71565
R179 VTAIL.n60 VTAIL.n40 2.71565
R180 VTAIL.n119 VTAIL.n117 2.41305
R181 VTAIL.n11 VTAIL.n9 2.41305
R182 VTAIL.n83 VTAIL.n81 2.41305
R183 VTAIL.n47 VTAIL.n45 2.41305
R184 VTAIL.n136 VTAIL.n135 1.93989
R185 VTAIL.n28 VTAIL.n27 1.93989
R186 VTAIL.n100 VTAIL.n99 1.93989
R187 VTAIL.n64 VTAIL.n63 1.93989
R188 VTAIL.n139 VTAIL.n110 1.16414
R189 VTAIL.n31 VTAIL.n2 1.16414
R190 VTAIL.n103 VTAIL.n74 1.16414
R191 VTAIL.n67 VTAIL.n38 1.16414
R192 VTAIL.n107 VTAIL.n71 0.733259
R193 VTAIL VTAIL.n35 0.659983
R194 VTAIL.n125 VTAIL.n117 0.155672
R195 VTAIL.n126 VTAIL.n125 0.155672
R196 VTAIL.n126 VTAIL.n113 0.155672
R197 VTAIL.n133 VTAIL.n113 0.155672
R198 VTAIL.n134 VTAIL.n133 0.155672
R199 VTAIL.n134 VTAIL.n109 0.155672
R200 VTAIL.n141 VTAIL.n109 0.155672
R201 VTAIL.n17 VTAIL.n9 0.155672
R202 VTAIL.n18 VTAIL.n17 0.155672
R203 VTAIL.n18 VTAIL.n5 0.155672
R204 VTAIL.n25 VTAIL.n5 0.155672
R205 VTAIL.n26 VTAIL.n25 0.155672
R206 VTAIL.n26 VTAIL.n1 0.155672
R207 VTAIL.n33 VTAIL.n1 0.155672
R208 VTAIL.n105 VTAIL.n73 0.155672
R209 VTAIL.n98 VTAIL.n73 0.155672
R210 VTAIL.n98 VTAIL.n97 0.155672
R211 VTAIL.n97 VTAIL.n77 0.155672
R212 VTAIL.n90 VTAIL.n77 0.155672
R213 VTAIL.n90 VTAIL.n89 0.155672
R214 VTAIL.n89 VTAIL.n81 0.155672
R215 VTAIL.n69 VTAIL.n37 0.155672
R216 VTAIL.n62 VTAIL.n37 0.155672
R217 VTAIL.n62 VTAIL.n61 0.155672
R218 VTAIL.n61 VTAIL.n41 0.155672
R219 VTAIL.n54 VTAIL.n41 0.155672
R220 VTAIL.n54 VTAIL.n53 0.155672
R221 VTAIL.n53 VTAIL.n45 0.155672
R222 VTAIL VTAIL.n143 0.0737759
R223 VDD2.n66 VDD2.n65 585
R224 VDD2.n64 VDD2.n63 585
R225 VDD2.n39 VDD2.n38 585
R226 VDD2.n58 VDD2.n57 585
R227 VDD2.n56 VDD2.n55 585
R228 VDD2.n43 VDD2.n42 585
R229 VDD2.n50 VDD2.n49 585
R230 VDD2.n48 VDD2.n47 585
R231 VDD2.n13 VDD2.n12 585
R232 VDD2.n15 VDD2.n14 585
R233 VDD2.n8 VDD2.n7 585
R234 VDD2.n21 VDD2.n20 585
R235 VDD2.n23 VDD2.n22 585
R236 VDD2.n4 VDD2.n3 585
R237 VDD2.n29 VDD2.n28 585
R238 VDD2.n31 VDD2.n30 585
R239 VDD2.n65 VDD2.n35 498.474
R240 VDD2.n30 VDD2.n0 498.474
R241 VDD2.n46 VDD2.t0 329.053
R242 VDD2.n11 VDD2.t1 329.053
R243 VDD2.n65 VDD2.n64 171.744
R244 VDD2.n64 VDD2.n38 171.744
R245 VDD2.n57 VDD2.n38 171.744
R246 VDD2.n57 VDD2.n56 171.744
R247 VDD2.n56 VDD2.n42 171.744
R248 VDD2.n49 VDD2.n42 171.744
R249 VDD2.n49 VDD2.n48 171.744
R250 VDD2.n14 VDD2.n13 171.744
R251 VDD2.n14 VDD2.n7 171.744
R252 VDD2.n21 VDD2.n7 171.744
R253 VDD2.n22 VDD2.n21 171.744
R254 VDD2.n22 VDD2.n3 171.744
R255 VDD2.n29 VDD2.n3 171.744
R256 VDD2.n30 VDD2.n29 171.744
R257 VDD2.n48 VDD2.t0 85.8723
R258 VDD2.n13 VDD2.t1 85.8723
R259 VDD2.n70 VDD2.n34 84.3549
R260 VDD2.n70 VDD2.n69 53.3247
R261 VDD2.n67 VDD2.n66 12.8005
R262 VDD2.n32 VDD2.n31 12.8005
R263 VDD2.n63 VDD2.n37 12.0247
R264 VDD2.n28 VDD2.n2 12.0247
R265 VDD2.n62 VDD2.n39 11.249
R266 VDD2.n27 VDD2.n4 11.249
R267 VDD2.n47 VDD2.n46 10.7237
R268 VDD2.n12 VDD2.n11 10.7237
R269 VDD2.n59 VDD2.n58 10.4732
R270 VDD2.n24 VDD2.n23 10.4732
R271 VDD2.n55 VDD2.n41 9.69747
R272 VDD2.n20 VDD2.n6 9.69747
R273 VDD2.n69 VDD2.n68 9.45567
R274 VDD2.n34 VDD2.n33 9.45567
R275 VDD2.n45 VDD2.n44 9.3005
R276 VDD2.n52 VDD2.n51 9.3005
R277 VDD2.n54 VDD2.n53 9.3005
R278 VDD2.n41 VDD2.n40 9.3005
R279 VDD2.n60 VDD2.n59 9.3005
R280 VDD2.n62 VDD2.n61 9.3005
R281 VDD2.n37 VDD2.n36 9.3005
R282 VDD2.n68 VDD2.n67 9.3005
R283 VDD2.n10 VDD2.n9 9.3005
R284 VDD2.n17 VDD2.n16 9.3005
R285 VDD2.n19 VDD2.n18 9.3005
R286 VDD2.n6 VDD2.n5 9.3005
R287 VDD2.n25 VDD2.n24 9.3005
R288 VDD2.n27 VDD2.n26 9.3005
R289 VDD2.n2 VDD2.n1 9.3005
R290 VDD2.n33 VDD2.n32 9.3005
R291 VDD2.n54 VDD2.n43 8.92171
R292 VDD2.n19 VDD2.n8 8.92171
R293 VDD2.n51 VDD2.n50 8.14595
R294 VDD2.n16 VDD2.n15 8.14595
R295 VDD2.n69 VDD2.n35 7.75445
R296 VDD2.n34 VDD2.n0 7.75445
R297 VDD2.n47 VDD2.n45 7.3702
R298 VDD2.n12 VDD2.n10 7.3702
R299 VDD2.n67 VDD2.n35 6.08283
R300 VDD2.n32 VDD2.n0 6.08283
R301 VDD2.n50 VDD2.n45 5.81868
R302 VDD2.n15 VDD2.n10 5.81868
R303 VDD2.n51 VDD2.n43 5.04292
R304 VDD2.n16 VDD2.n8 5.04292
R305 VDD2.n55 VDD2.n54 4.26717
R306 VDD2.n20 VDD2.n19 4.26717
R307 VDD2.n58 VDD2.n41 3.49141
R308 VDD2.n23 VDD2.n6 3.49141
R309 VDD2.n59 VDD2.n39 2.71565
R310 VDD2.n24 VDD2.n4 2.71565
R311 VDD2.n46 VDD2.n44 2.41305
R312 VDD2.n11 VDD2.n9 2.41305
R313 VDD2.n63 VDD2.n62 1.93989
R314 VDD2.n28 VDD2.n27 1.93989
R315 VDD2.n66 VDD2.n37 1.16414
R316 VDD2.n31 VDD2.n2 1.16414
R317 VDD2 VDD2.n70 0.190155
R318 VDD2.n68 VDD2.n36 0.155672
R319 VDD2.n61 VDD2.n36 0.155672
R320 VDD2.n61 VDD2.n60 0.155672
R321 VDD2.n60 VDD2.n40 0.155672
R322 VDD2.n53 VDD2.n40 0.155672
R323 VDD2.n53 VDD2.n52 0.155672
R324 VDD2.n52 VDD2.n44 0.155672
R325 VDD2.n17 VDD2.n9 0.155672
R326 VDD2.n18 VDD2.n17 0.155672
R327 VDD2.n18 VDD2.n5 0.155672
R328 VDD2.n25 VDD2.n5 0.155672
R329 VDD2.n26 VDD2.n25 0.155672
R330 VDD2.n26 VDD2.n1 0.155672
R331 VDD2.n33 VDD2.n1 0.155672
R332 B.n76 B.t3 848.318
R333 B.n166 B.t9 848.318
R334 B.n28 B.t6 848.318
R335 B.n22 B.t0 848.318
R336 B.n212 B.n211 585
R337 B.n210 B.n57 585
R338 B.n209 B.n208 585
R339 B.n207 B.n58 585
R340 B.n206 B.n205 585
R341 B.n204 B.n59 585
R342 B.n203 B.n202 585
R343 B.n201 B.n60 585
R344 B.n200 B.n199 585
R345 B.n198 B.n61 585
R346 B.n197 B.n196 585
R347 B.n195 B.n62 585
R348 B.n194 B.n193 585
R349 B.n192 B.n63 585
R350 B.n191 B.n190 585
R351 B.n189 B.n64 585
R352 B.n188 B.n187 585
R353 B.n186 B.n65 585
R354 B.n185 B.n184 585
R355 B.n183 B.n66 585
R356 B.n182 B.n181 585
R357 B.n180 B.n67 585
R358 B.n179 B.n178 585
R359 B.n177 B.n68 585
R360 B.n176 B.n175 585
R361 B.n174 B.n69 585
R362 B.n173 B.n172 585
R363 B.n171 B.n70 585
R364 B.n170 B.n169 585
R365 B.n165 B.n71 585
R366 B.n164 B.n163 585
R367 B.n162 B.n72 585
R368 B.n161 B.n160 585
R369 B.n159 B.n73 585
R370 B.n158 B.n157 585
R371 B.n156 B.n74 585
R372 B.n155 B.n154 585
R373 B.n152 B.n75 585
R374 B.n151 B.n150 585
R375 B.n149 B.n78 585
R376 B.n148 B.n147 585
R377 B.n146 B.n79 585
R378 B.n145 B.n144 585
R379 B.n143 B.n80 585
R380 B.n142 B.n141 585
R381 B.n140 B.n81 585
R382 B.n139 B.n138 585
R383 B.n137 B.n82 585
R384 B.n136 B.n135 585
R385 B.n134 B.n83 585
R386 B.n133 B.n132 585
R387 B.n131 B.n84 585
R388 B.n130 B.n129 585
R389 B.n128 B.n85 585
R390 B.n127 B.n126 585
R391 B.n125 B.n86 585
R392 B.n124 B.n123 585
R393 B.n122 B.n87 585
R394 B.n121 B.n120 585
R395 B.n119 B.n88 585
R396 B.n118 B.n117 585
R397 B.n116 B.n89 585
R398 B.n115 B.n114 585
R399 B.n113 B.n90 585
R400 B.n112 B.n111 585
R401 B.n213 B.n56 585
R402 B.n215 B.n214 585
R403 B.n216 B.n55 585
R404 B.n218 B.n217 585
R405 B.n219 B.n54 585
R406 B.n221 B.n220 585
R407 B.n222 B.n53 585
R408 B.n224 B.n223 585
R409 B.n225 B.n52 585
R410 B.n227 B.n226 585
R411 B.n228 B.n51 585
R412 B.n230 B.n229 585
R413 B.n231 B.n50 585
R414 B.n233 B.n232 585
R415 B.n234 B.n49 585
R416 B.n236 B.n235 585
R417 B.n237 B.n48 585
R418 B.n239 B.n238 585
R419 B.n240 B.n47 585
R420 B.n242 B.n241 585
R421 B.n243 B.n46 585
R422 B.n245 B.n244 585
R423 B.n246 B.n45 585
R424 B.n248 B.n247 585
R425 B.n347 B.n346 585
R426 B.n345 B.n8 585
R427 B.n344 B.n343 585
R428 B.n342 B.n9 585
R429 B.n341 B.n340 585
R430 B.n339 B.n10 585
R431 B.n338 B.n337 585
R432 B.n336 B.n11 585
R433 B.n335 B.n334 585
R434 B.n333 B.n12 585
R435 B.n332 B.n331 585
R436 B.n330 B.n13 585
R437 B.n329 B.n328 585
R438 B.n327 B.n14 585
R439 B.n326 B.n325 585
R440 B.n324 B.n15 585
R441 B.n323 B.n322 585
R442 B.n321 B.n16 585
R443 B.n320 B.n319 585
R444 B.n318 B.n17 585
R445 B.n317 B.n316 585
R446 B.n315 B.n18 585
R447 B.n314 B.n313 585
R448 B.n312 B.n19 585
R449 B.n311 B.n310 585
R450 B.n309 B.n20 585
R451 B.n308 B.n307 585
R452 B.n306 B.n21 585
R453 B.n304 B.n303 585
R454 B.n302 B.n24 585
R455 B.n301 B.n300 585
R456 B.n299 B.n25 585
R457 B.n298 B.n297 585
R458 B.n296 B.n26 585
R459 B.n295 B.n294 585
R460 B.n293 B.n27 585
R461 B.n292 B.n291 585
R462 B.n290 B.n289 585
R463 B.n288 B.n31 585
R464 B.n287 B.n286 585
R465 B.n285 B.n32 585
R466 B.n284 B.n283 585
R467 B.n282 B.n33 585
R468 B.n281 B.n280 585
R469 B.n279 B.n34 585
R470 B.n278 B.n277 585
R471 B.n276 B.n35 585
R472 B.n275 B.n274 585
R473 B.n273 B.n36 585
R474 B.n272 B.n271 585
R475 B.n270 B.n37 585
R476 B.n269 B.n268 585
R477 B.n267 B.n38 585
R478 B.n266 B.n265 585
R479 B.n264 B.n39 585
R480 B.n263 B.n262 585
R481 B.n261 B.n40 585
R482 B.n260 B.n259 585
R483 B.n258 B.n41 585
R484 B.n257 B.n256 585
R485 B.n255 B.n42 585
R486 B.n254 B.n253 585
R487 B.n252 B.n43 585
R488 B.n251 B.n250 585
R489 B.n249 B.n44 585
R490 B.n348 B.n7 585
R491 B.n350 B.n349 585
R492 B.n351 B.n6 585
R493 B.n353 B.n352 585
R494 B.n354 B.n5 585
R495 B.n356 B.n355 585
R496 B.n357 B.n4 585
R497 B.n359 B.n358 585
R498 B.n360 B.n3 585
R499 B.n362 B.n361 585
R500 B.n363 B.n0 585
R501 B.n2 B.n1 585
R502 B.n97 B.n96 585
R503 B.n98 B.n95 585
R504 B.n100 B.n99 585
R505 B.n101 B.n94 585
R506 B.n103 B.n102 585
R507 B.n104 B.n93 585
R508 B.n106 B.n105 585
R509 B.n107 B.n92 585
R510 B.n109 B.n108 585
R511 B.n110 B.n91 585
R512 B.n112 B.n91 559.769
R513 B.n213 B.n212 559.769
R514 B.n249 B.n248 559.769
R515 B.n346 B.n7 559.769
R516 B.n166 B.t10 303.156
R517 B.n28 B.t8 303.156
R518 B.n76 B.t4 303.156
R519 B.n22 B.t2 303.156
R520 B.n167 B.t11 291.325
R521 B.n29 B.t7 291.325
R522 B.n77 B.t5 291.325
R523 B.n23 B.t1 291.325
R524 B.n365 B.n364 256.663
R525 B.n364 B.n363 235.042
R526 B.n364 B.n2 235.042
R527 B.n113 B.n112 163.367
R528 B.n114 B.n113 163.367
R529 B.n114 B.n89 163.367
R530 B.n118 B.n89 163.367
R531 B.n119 B.n118 163.367
R532 B.n120 B.n119 163.367
R533 B.n120 B.n87 163.367
R534 B.n124 B.n87 163.367
R535 B.n125 B.n124 163.367
R536 B.n126 B.n125 163.367
R537 B.n126 B.n85 163.367
R538 B.n130 B.n85 163.367
R539 B.n131 B.n130 163.367
R540 B.n132 B.n131 163.367
R541 B.n132 B.n83 163.367
R542 B.n136 B.n83 163.367
R543 B.n137 B.n136 163.367
R544 B.n138 B.n137 163.367
R545 B.n138 B.n81 163.367
R546 B.n142 B.n81 163.367
R547 B.n143 B.n142 163.367
R548 B.n144 B.n143 163.367
R549 B.n144 B.n79 163.367
R550 B.n148 B.n79 163.367
R551 B.n149 B.n148 163.367
R552 B.n150 B.n149 163.367
R553 B.n150 B.n75 163.367
R554 B.n155 B.n75 163.367
R555 B.n156 B.n155 163.367
R556 B.n157 B.n156 163.367
R557 B.n157 B.n73 163.367
R558 B.n161 B.n73 163.367
R559 B.n162 B.n161 163.367
R560 B.n163 B.n162 163.367
R561 B.n163 B.n71 163.367
R562 B.n170 B.n71 163.367
R563 B.n171 B.n170 163.367
R564 B.n172 B.n171 163.367
R565 B.n172 B.n69 163.367
R566 B.n176 B.n69 163.367
R567 B.n177 B.n176 163.367
R568 B.n178 B.n177 163.367
R569 B.n178 B.n67 163.367
R570 B.n182 B.n67 163.367
R571 B.n183 B.n182 163.367
R572 B.n184 B.n183 163.367
R573 B.n184 B.n65 163.367
R574 B.n188 B.n65 163.367
R575 B.n189 B.n188 163.367
R576 B.n190 B.n189 163.367
R577 B.n190 B.n63 163.367
R578 B.n194 B.n63 163.367
R579 B.n195 B.n194 163.367
R580 B.n196 B.n195 163.367
R581 B.n196 B.n61 163.367
R582 B.n200 B.n61 163.367
R583 B.n201 B.n200 163.367
R584 B.n202 B.n201 163.367
R585 B.n202 B.n59 163.367
R586 B.n206 B.n59 163.367
R587 B.n207 B.n206 163.367
R588 B.n208 B.n207 163.367
R589 B.n208 B.n57 163.367
R590 B.n212 B.n57 163.367
R591 B.n248 B.n45 163.367
R592 B.n244 B.n45 163.367
R593 B.n244 B.n243 163.367
R594 B.n243 B.n242 163.367
R595 B.n242 B.n47 163.367
R596 B.n238 B.n47 163.367
R597 B.n238 B.n237 163.367
R598 B.n237 B.n236 163.367
R599 B.n236 B.n49 163.367
R600 B.n232 B.n49 163.367
R601 B.n232 B.n231 163.367
R602 B.n231 B.n230 163.367
R603 B.n230 B.n51 163.367
R604 B.n226 B.n51 163.367
R605 B.n226 B.n225 163.367
R606 B.n225 B.n224 163.367
R607 B.n224 B.n53 163.367
R608 B.n220 B.n53 163.367
R609 B.n220 B.n219 163.367
R610 B.n219 B.n218 163.367
R611 B.n218 B.n55 163.367
R612 B.n214 B.n55 163.367
R613 B.n214 B.n213 163.367
R614 B.n346 B.n345 163.367
R615 B.n345 B.n344 163.367
R616 B.n344 B.n9 163.367
R617 B.n340 B.n9 163.367
R618 B.n340 B.n339 163.367
R619 B.n339 B.n338 163.367
R620 B.n338 B.n11 163.367
R621 B.n334 B.n11 163.367
R622 B.n334 B.n333 163.367
R623 B.n333 B.n332 163.367
R624 B.n332 B.n13 163.367
R625 B.n328 B.n13 163.367
R626 B.n328 B.n327 163.367
R627 B.n327 B.n326 163.367
R628 B.n326 B.n15 163.367
R629 B.n322 B.n15 163.367
R630 B.n322 B.n321 163.367
R631 B.n321 B.n320 163.367
R632 B.n320 B.n17 163.367
R633 B.n316 B.n17 163.367
R634 B.n316 B.n315 163.367
R635 B.n315 B.n314 163.367
R636 B.n314 B.n19 163.367
R637 B.n310 B.n19 163.367
R638 B.n310 B.n309 163.367
R639 B.n309 B.n308 163.367
R640 B.n308 B.n21 163.367
R641 B.n303 B.n21 163.367
R642 B.n303 B.n302 163.367
R643 B.n302 B.n301 163.367
R644 B.n301 B.n25 163.367
R645 B.n297 B.n25 163.367
R646 B.n297 B.n296 163.367
R647 B.n296 B.n295 163.367
R648 B.n295 B.n27 163.367
R649 B.n291 B.n27 163.367
R650 B.n291 B.n290 163.367
R651 B.n290 B.n31 163.367
R652 B.n286 B.n31 163.367
R653 B.n286 B.n285 163.367
R654 B.n285 B.n284 163.367
R655 B.n284 B.n33 163.367
R656 B.n280 B.n33 163.367
R657 B.n280 B.n279 163.367
R658 B.n279 B.n278 163.367
R659 B.n278 B.n35 163.367
R660 B.n274 B.n35 163.367
R661 B.n274 B.n273 163.367
R662 B.n273 B.n272 163.367
R663 B.n272 B.n37 163.367
R664 B.n268 B.n37 163.367
R665 B.n268 B.n267 163.367
R666 B.n267 B.n266 163.367
R667 B.n266 B.n39 163.367
R668 B.n262 B.n39 163.367
R669 B.n262 B.n261 163.367
R670 B.n261 B.n260 163.367
R671 B.n260 B.n41 163.367
R672 B.n256 B.n41 163.367
R673 B.n256 B.n255 163.367
R674 B.n255 B.n254 163.367
R675 B.n254 B.n43 163.367
R676 B.n250 B.n43 163.367
R677 B.n250 B.n249 163.367
R678 B.n350 B.n7 163.367
R679 B.n351 B.n350 163.367
R680 B.n352 B.n351 163.367
R681 B.n352 B.n5 163.367
R682 B.n356 B.n5 163.367
R683 B.n357 B.n356 163.367
R684 B.n358 B.n357 163.367
R685 B.n358 B.n3 163.367
R686 B.n362 B.n3 163.367
R687 B.n363 B.n362 163.367
R688 B.n96 B.n2 163.367
R689 B.n96 B.n95 163.367
R690 B.n100 B.n95 163.367
R691 B.n101 B.n100 163.367
R692 B.n102 B.n101 163.367
R693 B.n102 B.n93 163.367
R694 B.n106 B.n93 163.367
R695 B.n107 B.n106 163.367
R696 B.n108 B.n107 163.367
R697 B.n108 B.n91 163.367
R698 B.n153 B.n77 59.5399
R699 B.n168 B.n167 59.5399
R700 B.n30 B.n29 59.5399
R701 B.n305 B.n23 59.5399
R702 B.n348 B.n347 36.3712
R703 B.n247 B.n44 36.3712
R704 B.n211 B.n56 36.3712
R705 B.n111 B.n110 36.3712
R706 B B.n365 18.0485
R707 B.n77 B.n76 11.8308
R708 B.n167 B.n166 11.8308
R709 B.n29 B.n28 11.8308
R710 B.n23 B.n22 11.8308
R711 B.n349 B.n348 10.6151
R712 B.n349 B.n6 10.6151
R713 B.n353 B.n6 10.6151
R714 B.n354 B.n353 10.6151
R715 B.n355 B.n354 10.6151
R716 B.n355 B.n4 10.6151
R717 B.n359 B.n4 10.6151
R718 B.n360 B.n359 10.6151
R719 B.n361 B.n360 10.6151
R720 B.n361 B.n0 10.6151
R721 B.n347 B.n8 10.6151
R722 B.n343 B.n8 10.6151
R723 B.n343 B.n342 10.6151
R724 B.n342 B.n341 10.6151
R725 B.n341 B.n10 10.6151
R726 B.n337 B.n10 10.6151
R727 B.n337 B.n336 10.6151
R728 B.n336 B.n335 10.6151
R729 B.n335 B.n12 10.6151
R730 B.n331 B.n12 10.6151
R731 B.n331 B.n330 10.6151
R732 B.n330 B.n329 10.6151
R733 B.n329 B.n14 10.6151
R734 B.n325 B.n14 10.6151
R735 B.n325 B.n324 10.6151
R736 B.n324 B.n323 10.6151
R737 B.n323 B.n16 10.6151
R738 B.n319 B.n16 10.6151
R739 B.n319 B.n318 10.6151
R740 B.n318 B.n317 10.6151
R741 B.n317 B.n18 10.6151
R742 B.n313 B.n18 10.6151
R743 B.n313 B.n312 10.6151
R744 B.n312 B.n311 10.6151
R745 B.n311 B.n20 10.6151
R746 B.n307 B.n20 10.6151
R747 B.n307 B.n306 10.6151
R748 B.n304 B.n24 10.6151
R749 B.n300 B.n24 10.6151
R750 B.n300 B.n299 10.6151
R751 B.n299 B.n298 10.6151
R752 B.n298 B.n26 10.6151
R753 B.n294 B.n26 10.6151
R754 B.n294 B.n293 10.6151
R755 B.n293 B.n292 10.6151
R756 B.n289 B.n288 10.6151
R757 B.n288 B.n287 10.6151
R758 B.n287 B.n32 10.6151
R759 B.n283 B.n32 10.6151
R760 B.n283 B.n282 10.6151
R761 B.n282 B.n281 10.6151
R762 B.n281 B.n34 10.6151
R763 B.n277 B.n34 10.6151
R764 B.n277 B.n276 10.6151
R765 B.n276 B.n275 10.6151
R766 B.n275 B.n36 10.6151
R767 B.n271 B.n36 10.6151
R768 B.n271 B.n270 10.6151
R769 B.n270 B.n269 10.6151
R770 B.n269 B.n38 10.6151
R771 B.n265 B.n38 10.6151
R772 B.n265 B.n264 10.6151
R773 B.n264 B.n263 10.6151
R774 B.n263 B.n40 10.6151
R775 B.n259 B.n40 10.6151
R776 B.n259 B.n258 10.6151
R777 B.n258 B.n257 10.6151
R778 B.n257 B.n42 10.6151
R779 B.n253 B.n42 10.6151
R780 B.n253 B.n252 10.6151
R781 B.n252 B.n251 10.6151
R782 B.n251 B.n44 10.6151
R783 B.n247 B.n246 10.6151
R784 B.n246 B.n245 10.6151
R785 B.n245 B.n46 10.6151
R786 B.n241 B.n46 10.6151
R787 B.n241 B.n240 10.6151
R788 B.n240 B.n239 10.6151
R789 B.n239 B.n48 10.6151
R790 B.n235 B.n48 10.6151
R791 B.n235 B.n234 10.6151
R792 B.n234 B.n233 10.6151
R793 B.n233 B.n50 10.6151
R794 B.n229 B.n50 10.6151
R795 B.n229 B.n228 10.6151
R796 B.n228 B.n227 10.6151
R797 B.n227 B.n52 10.6151
R798 B.n223 B.n52 10.6151
R799 B.n223 B.n222 10.6151
R800 B.n222 B.n221 10.6151
R801 B.n221 B.n54 10.6151
R802 B.n217 B.n54 10.6151
R803 B.n217 B.n216 10.6151
R804 B.n216 B.n215 10.6151
R805 B.n215 B.n56 10.6151
R806 B.n97 B.n1 10.6151
R807 B.n98 B.n97 10.6151
R808 B.n99 B.n98 10.6151
R809 B.n99 B.n94 10.6151
R810 B.n103 B.n94 10.6151
R811 B.n104 B.n103 10.6151
R812 B.n105 B.n104 10.6151
R813 B.n105 B.n92 10.6151
R814 B.n109 B.n92 10.6151
R815 B.n110 B.n109 10.6151
R816 B.n111 B.n90 10.6151
R817 B.n115 B.n90 10.6151
R818 B.n116 B.n115 10.6151
R819 B.n117 B.n116 10.6151
R820 B.n117 B.n88 10.6151
R821 B.n121 B.n88 10.6151
R822 B.n122 B.n121 10.6151
R823 B.n123 B.n122 10.6151
R824 B.n123 B.n86 10.6151
R825 B.n127 B.n86 10.6151
R826 B.n128 B.n127 10.6151
R827 B.n129 B.n128 10.6151
R828 B.n129 B.n84 10.6151
R829 B.n133 B.n84 10.6151
R830 B.n134 B.n133 10.6151
R831 B.n135 B.n134 10.6151
R832 B.n135 B.n82 10.6151
R833 B.n139 B.n82 10.6151
R834 B.n140 B.n139 10.6151
R835 B.n141 B.n140 10.6151
R836 B.n141 B.n80 10.6151
R837 B.n145 B.n80 10.6151
R838 B.n146 B.n145 10.6151
R839 B.n147 B.n146 10.6151
R840 B.n147 B.n78 10.6151
R841 B.n151 B.n78 10.6151
R842 B.n152 B.n151 10.6151
R843 B.n154 B.n74 10.6151
R844 B.n158 B.n74 10.6151
R845 B.n159 B.n158 10.6151
R846 B.n160 B.n159 10.6151
R847 B.n160 B.n72 10.6151
R848 B.n164 B.n72 10.6151
R849 B.n165 B.n164 10.6151
R850 B.n169 B.n165 10.6151
R851 B.n173 B.n70 10.6151
R852 B.n174 B.n173 10.6151
R853 B.n175 B.n174 10.6151
R854 B.n175 B.n68 10.6151
R855 B.n179 B.n68 10.6151
R856 B.n180 B.n179 10.6151
R857 B.n181 B.n180 10.6151
R858 B.n181 B.n66 10.6151
R859 B.n185 B.n66 10.6151
R860 B.n186 B.n185 10.6151
R861 B.n187 B.n186 10.6151
R862 B.n187 B.n64 10.6151
R863 B.n191 B.n64 10.6151
R864 B.n192 B.n191 10.6151
R865 B.n193 B.n192 10.6151
R866 B.n193 B.n62 10.6151
R867 B.n197 B.n62 10.6151
R868 B.n198 B.n197 10.6151
R869 B.n199 B.n198 10.6151
R870 B.n199 B.n60 10.6151
R871 B.n203 B.n60 10.6151
R872 B.n204 B.n203 10.6151
R873 B.n205 B.n204 10.6151
R874 B.n205 B.n58 10.6151
R875 B.n209 B.n58 10.6151
R876 B.n210 B.n209 10.6151
R877 B.n211 B.n210 10.6151
R878 B.n365 B.n0 8.11757
R879 B.n365 B.n1 8.11757
R880 B.n305 B.n304 7.18099
R881 B.n292 B.n30 7.18099
R882 B.n154 B.n153 7.18099
R883 B.n169 B.n168 7.18099
R884 B.n306 B.n305 3.43465
R885 B.n289 B.n30 3.43465
R886 B.n153 B.n152 3.43465
R887 B.n168 B.n70 3.43465
R888 VP.n0 VP.t0 962.303
R889 VP.n0 VP.t1 927.337
R890 VP VP.n0 0.0516364
R891 VDD1.n31 VDD1.n30 585
R892 VDD1.n29 VDD1.n28 585
R893 VDD1.n4 VDD1.n3 585
R894 VDD1.n23 VDD1.n22 585
R895 VDD1.n21 VDD1.n20 585
R896 VDD1.n8 VDD1.n7 585
R897 VDD1.n15 VDD1.n14 585
R898 VDD1.n13 VDD1.n12 585
R899 VDD1.n48 VDD1.n47 585
R900 VDD1.n50 VDD1.n49 585
R901 VDD1.n43 VDD1.n42 585
R902 VDD1.n56 VDD1.n55 585
R903 VDD1.n58 VDD1.n57 585
R904 VDD1.n39 VDD1.n38 585
R905 VDD1.n64 VDD1.n63 585
R906 VDD1.n66 VDD1.n65 585
R907 VDD1.n30 VDD1.n0 498.474
R908 VDD1.n65 VDD1.n35 498.474
R909 VDD1.n11 VDD1.t1 329.053
R910 VDD1.n46 VDD1.t0 329.053
R911 VDD1.n30 VDD1.n29 171.744
R912 VDD1.n29 VDD1.n3 171.744
R913 VDD1.n22 VDD1.n3 171.744
R914 VDD1.n22 VDD1.n21 171.744
R915 VDD1.n21 VDD1.n7 171.744
R916 VDD1.n14 VDD1.n7 171.744
R917 VDD1.n14 VDD1.n13 171.744
R918 VDD1.n49 VDD1.n48 171.744
R919 VDD1.n49 VDD1.n42 171.744
R920 VDD1.n56 VDD1.n42 171.744
R921 VDD1.n57 VDD1.n56 171.744
R922 VDD1.n57 VDD1.n38 171.744
R923 VDD1.n64 VDD1.n38 171.744
R924 VDD1.n65 VDD1.n64 171.744
R925 VDD1.n13 VDD1.t1 85.8723
R926 VDD1.n48 VDD1.t0 85.8723
R927 VDD1 VDD1.n69 85.0112
R928 VDD1 VDD1.n34 53.5144
R929 VDD1.n32 VDD1.n31 12.8005
R930 VDD1.n67 VDD1.n66 12.8005
R931 VDD1.n28 VDD1.n2 12.0247
R932 VDD1.n63 VDD1.n37 12.0247
R933 VDD1.n27 VDD1.n4 11.249
R934 VDD1.n62 VDD1.n39 11.249
R935 VDD1.n12 VDD1.n11 10.7237
R936 VDD1.n47 VDD1.n46 10.7237
R937 VDD1.n24 VDD1.n23 10.4732
R938 VDD1.n59 VDD1.n58 10.4732
R939 VDD1.n20 VDD1.n6 9.69747
R940 VDD1.n55 VDD1.n41 9.69747
R941 VDD1.n34 VDD1.n33 9.45567
R942 VDD1.n69 VDD1.n68 9.45567
R943 VDD1.n10 VDD1.n9 9.3005
R944 VDD1.n17 VDD1.n16 9.3005
R945 VDD1.n19 VDD1.n18 9.3005
R946 VDD1.n6 VDD1.n5 9.3005
R947 VDD1.n25 VDD1.n24 9.3005
R948 VDD1.n27 VDD1.n26 9.3005
R949 VDD1.n2 VDD1.n1 9.3005
R950 VDD1.n33 VDD1.n32 9.3005
R951 VDD1.n45 VDD1.n44 9.3005
R952 VDD1.n52 VDD1.n51 9.3005
R953 VDD1.n54 VDD1.n53 9.3005
R954 VDD1.n41 VDD1.n40 9.3005
R955 VDD1.n60 VDD1.n59 9.3005
R956 VDD1.n62 VDD1.n61 9.3005
R957 VDD1.n37 VDD1.n36 9.3005
R958 VDD1.n68 VDD1.n67 9.3005
R959 VDD1.n19 VDD1.n8 8.92171
R960 VDD1.n54 VDD1.n43 8.92171
R961 VDD1.n16 VDD1.n15 8.14595
R962 VDD1.n51 VDD1.n50 8.14595
R963 VDD1.n34 VDD1.n0 7.75445
R964 VDD1.n69 VDD1.n35 7.75445
R965 VDD1.n12 VDD1.n10 7.3702
R966 VDD1.n47 VDD1.n45 7.3702
R967 VDD1.n32 VDD1.n0 6.08283
R968 VDD1.n67 VDD1.n35 6.08283
R969 VDD1.n15 VDD1.n10 5.81868
R970 VDD1.n50 VDD1.n45 5.81868
R971 VDD1.n16 VDD1.n8 5.04292
R972 VDD1.n51 VDD1.n43 5.04292
R973 VDD1.n20 VDD1.n19 4.26717
R974 VDD1.n55 VDD1.n54 4.26717
R975 VDD1.n23 VDD1.n6 3.49141
R976 VDD1.n58 VDD1.n41 3.49141
R977 VDD1.n24 VDD1.n4 2.71565
R978 VDD1.n59 VDD1.n39 2.71565
R979 VDD1.n11 VDD1.n9 2.41305
R980 VDD1.n46 VDD1.n44 2.41305
R981 VDD1.n28 VDD1.n27 1.93989
R982 VDD1.n63 VDD1.n62 1.93989
R983 VDD1.n31 VDD1.n2 1.16414
R984 VDD1.n66 VDD1.n37 1.16414
R985 VDD1.n33 VDD1.n1 0.155672
R986 VDD1.n26 VDD1.n1 0.155672
R987 VDD1.n26 VDD1.n25 0.155672
R988 VDD1.n25 VDD1.n5 0.155672
R989 VDD1.n18 VDD1.n5 0.155672
R990 VDD1.n18 VDD1.n17 0.155672
R991 VDD1.n17 VDD1.n9 0.155672
R992 VDD1.n52 VDD1.n44 0.155672
R993 VDD1.n53 VDD1.n52 0.155672
R994 VDD1.n53 VDD1.n40 0.155672
R995 VDD1.n60 VDD1.n40 0.155672
R996 VDD1.n61 VDD1.n60 0.155672
R997 VDD1.n61 VDD1.n36 0.155672
R998 VDD1.n68 VDD1.n36 0.155672
C0 VN B 0.599354f
C1 B VDD1 1.0063f
C2 VTAIL VP 0.602263f
C3 VN VP 3.50601f
C4 w_n1214_n2434# VTAIL 2.18676f
C5 VP VDD1 1.03096f
C6 VDD2 VTAIL 4.780221f
C7 VN w_n1214_n2434# 1.41962f
C8 w_n1214_n2434# VDD1 1.17299f
C9 VDD2 VN 0.945712f
C10 VDD2 VDD1 0.42332f
C11 VN VTAIL 0.587752f
C12 VTAIL VDD1 4.74771f
C13 VP B 0.836058f
C14 VN VDD1 0.14839f
C15 w_n1214_n2434# B 5.01138f
C16 VDD2 B 1.01809f
C17 w_n1214_n2434# VP 1.56925f
C18 VDD2 VP 0.236748f
C19 VTAIL B 1.66836f
C20 VDD2 w_n1214_n2434# 1.1735f
C21 VDD2 VSUBS 0.557513f
C22 VDD1 VSUBS 2.344347f
C23 VTAIL VSUBS 0.205364f
C24 VN VSUBS 4.16496f
C25 VP VSUBS 0.809692f
C26 B VSUBS 1.791293f
C27 w_n1214_n2434# VSUBS 36.7259f
C28 VDD1.n0 VSUBS 0.021198f
C29 VDD1.n1 VSUBS 0.018964f
C30 VDD1.n2 VSUBS 0.01019f
C31 VDD1.n3 VSUBS 0.024087f
C32 VDD1.n4 VSUBS 0.01079f
C33 VDD1.n5 VSUBS 0.018964f
C34 VDD1.n6 VSUBS 0.01019f
C35 VDD1.n7 VSUBS 0.024087f
C36 VDD1.n8 VSUBS 0.01079f
C37 VDD1.n9 VSUBS 0.541745f
C38 VDD1.n10 VSUBS 0.01019f
C39 VDD1.t1 VSUBS 0.051775f
C40 VDD1.n11 VSUBS 0.10928f
C41 VDD1.n12 VSUBS 0.018118f
C42 VDD1.n13 VSUBS 0.018065f
C43 VDD1.n14 VSUBS 0.024087f
C44 VDD1.n15 VSUBS 0.01079f
C45 VDD1.n16 VSUBS 0.01019f
C46 VDD1.n17 VSUBS 0.018964f
C47 VDD1.n18 VSUBS 0.018964f
C48 VDD1.n19 VSUBS 0.01019f
C49 VDD1.n20 VSUBS 0.01079f
C50 VDD1.n21 VSUBS 0.024087f
C51 VDD1.n22 VSUBS 0.024087f
C52 VDD1.n23 VSUBS 0.01079f
C53 VDD1.n24 VSUBS 0.01019f
C54 VDD1.n25 VSUBS 0.018964f
C55 VDD1.n26 VSUBS 0.018964f
C56 VDD1.n27 VSUBS 0.01019f
C57 VDD1.n28 VSUBS 0.01079f
C58 VDD1.n29 VSUBS 0.024087f
C59 VDD1.n30 VSUBS 0.061233f
C60 VDD1.n31 VSUBS 0.01079f
C61 VDD1.n32 VSUBS 0.020012f
C62 VDD1.n33 VSUBS 0.049793f
C63 VDD1.n34 VSUBS 0.06089f
C64 VDD1.n35 VSUBS 0.021198f
C65 VDD1.n36 VSUBS 0.018964f
C66 VDD1.n37 VSUBS 0.01019f
C67 VDD1.n38 VSUBS 0.024087f
C68 VDD1.n39 VSUBS 0.01079f
C69 VDD1.n40 VSUBS 0.018964f
C70 VDD1.n41 VSUBS 0.01019f
C71 VDD1.n42 VSUBS 0.024087f
C72 VDD1.n43 VSUBS 0.01079f
C73 VDD1.n44 VSUBS 0.541745f
C74 VDD1.n45 VSUBS 0.01019f
C75 VDD1.t0 VSUBS 0.051775f
C76 VDD1.n46 VSUBS 0.10928f
C77 VDD1.n47 VSUBS 0.018118f
C78 VDD1.n48 VSUBS 0.018065f
C79 VDD1.n49 VSUBS 0.024087f
C80 VDD1.n50 VSUBS 0.01079f
C81 VDD1.n51 VSUBS 0.01019f
C82 VDD1.n52 VSUBS 0.018964f
C83 VDD1.n53 VSUBS 0.018964f
C84 VDD1.n54 VSUBS 0.01019f
C85 VDD1.n55 VSUBS 0.01079f
C86 VDD1.n56 VSUBS 0.024087f
C87 VDD1.n57 VSUBS 0.024087f
C88 VDD1.n58 VSUBS 0.01079f
C89 VDD1.n59 VSUBS 0.01019f
C90 VDD1.n60 VSUBS 0.018964f
C91 VDD1.n61 VSUBS 0.018964f
C92 VDD1.n62 VSUBS 0.01019f
C93 VDD1.n63 VSUBS 0.01079f
C94 VDD1.n64 VSUBS 0.024087f
C95 VDD1.n65 VSUBS 0.061233f
C96 VDD1.n66 VSUBS 0.01079f
C97 VDD1.n67 VSUBS 0.020012f
C98 VDD1.n68 VSUBS 0.049793f
C99 VDD1.n69 VSUBS 0.360093f
C100 VP.t0 VSUBS 0.339575f
C101 VP.t1 VSUBS 0.287281f
C102 VP.n0 VSUBS 2.8677f
C103 B.n0 VSUBS 0.005711f
C104 B.n1 VSUBS 0.005711f
C105 B.n2 VSUBS 0.008446f
C106 B.n3 VSUBS 0.006472f
C107 B.n4 VSUBS 0.006472f
C108 B.n5 VSUBS 0.006472f
C109 B.n6 VSUBS 0.006472f
C110 B.n7 VSUBS 0.015932f
C111 B.n8 VSUBS 0.006472f
C112 B.n9 VSUBS 0.006472f
C113 B.n10 VSUBS 0.006472f
C114 B.n11 VSUBS 0.006472f
C115 B.n12 VSUBS 0.006472f
C116 B.n13 VSUBS 0.006472f
C117 B.n14 VSUBS 0.006472f
C118 B.n15 VSUBS 0.006472f
C119 B.n16 VSUBS 0.006472f
C120 B.n17 VSUBS 0.006472f
C121 B.n18 VSUBS 0.006472f
C122 B.n19 VSUBS 0.006472f
C123 B.n20 VSUBS 0.006472f
C124 B.n21 VSUBS 0.006472f
C125 B.t1 VSUBS 0.104747f
C126 B.t2 VSUBS 0.110535f
C127 B.t0 VSUBS 0.075858f
C128 B.n22 VSUBS 0.171423f
C129 B.n23 VSUBS 0.157542f
C130 B.n24 VSUBS 0.006472f
C131 B.n25 VSUBS 0.006472f
C132 B.n26 VSUBS 0.006472f
C133 B.n27 VSUBS 0.006472f
C134 B.t7 VSUBS 0.104749f
C135 B.t8 VSUBS 0.110537f
C136 B.t6 VSUBS 0.075858f
C137 B.n28 VSUBS 0.171421f
C138 B.n29 VSUBS 0.15754f
C139 B.n30 VSUBS 0.014995f
C140 B.n31 VSUBS 0.006472f
C141 B.n32 VSUBS 0.006472f
C142 B.n33 VSUBS 0.006472f
C143 B.n34 VSUBS 0.006472f
C144 B.n35 VSUBS 0.006472f
C145 B.n36 VSUBS 0.006472f
C146 B.n37 VSUBS 0.006472f
C147 B.n38 VSUBS 0.006472f
C148 B.n39 VSUBS 0.006472f
C149 B.n40 VSUBS 0.006472f
C150 B.n41 VSUBS 0.006472f
C151 B.n42 VSUBS 0.006472f
C152 B.n43 VSUBS 0.006472f
C153 B.n44 VSUBS 0.016619f
C154 B.n45 VSUBS 0.006472f
C155 B.n46 VSUBS 0.006472f
C156 B.n47 VSUBS 0.006472f
C157 B.n48 VSUBS 0.006472f
C158 B.n49 VSUBS 0.006472f
C159 B.n50 VSUBS 0.006472f
C160 B.n51 VSUBS 0.006472f
C161 B.n52 VSUBS 0.006472f
C162 B.n53 VSUBS 0.006472f
C163 B.n54 VSUBS 0.006472f
C164 B.n55 VSUBS 0.006472f
C165 B.n56 VSUBS 0.016619f
C166 B.n57 VSUBS 0.006472f
C167 B.n58 VSUBS 0.006472f
C168 B.n59 VSUBS 0.006472f
C169 B.n60 VSUBS 0.006472f
C170 B.n61 VSUBS 0.006472f
C171 B.n62 VSUBS 0.006472f
C172 B.n63 VSUBS 0.006472f
C173 B.n64 VSUBS 0.006472f
C174 B.n65 VSUBS 0.006472f
C175 B.n66 VSUBS 0.006472f
C176 B.n67 VSUBS 0.006472f
C177 B.n68 VSUBS 0.006472f
C178 B.n69 VSUBS 0.006472f
C179 B.n70 VSUBS 0.004283f
C180 B.n71 VSUBS 0.006472f
C181 B.n72 VSUBS 0.006472f
C182 B.n73 VSUBS 0.006472f
C183 B.n74 VSUBS 0.006472f
C184 B.n75 VSUBS 0.006472f
C185 B.t5 VSUBS 0.104747f
C186 B.t4 VSUBS 0.110535f
C187 B.t3 VSUBS 0.075858f
C188 B.n76 VSUBS 0.171423f
C189 B.n77 VSUBS 0.157542f
C190 B.n78 VSUBS 0.006472f
C191 B.n79 VSUBS 0.006472f
C192 B.n80 VSUBS 0.006472f
C193 B.n81 VSUBS 0.006472f
C194 B.n82 VSUBS 0.006472f
C195 B.n83 VSUBS 0.006472f
C196 B.n84 VSUBS 0.006472f
C197 B.n85 VSUBS 0.006472f
C198 B.n86 VSUBS 0.006472f
C199 B.n87 VSUBS 0.006472f
C200 B.n88 VSUBS 0.006472f
C201 B.n89 VSUBS 0.006472f
C202 B.n90 VSUBS 0.006472f
C203 B.n91 VSUBS 0.015932f
C204 B.n92 VSUBS 0.006472f
C205 B.n93 VSUBS 0.006472f
C206 B.n94 VSUBS 0.006472f
C207 B.n95 VSUBS 0.006472f
C208 B.n96 VSUBS 0.006472f
C209 B.n97 VSUBS 0.006472f
C210 B.n98 VSUBS 0.006472f
C211 B.n99 VSUBS 0.006472f
C212 B.n100 VSUBS 0.006472f
C213 B.n101 VSUBS 0.006472f
C214 B.n102 VSUBS 0.006472f
C215 B.n103 VSUBS 0.006472f
C216 B.n104 VSUBS 0.006472f
C217 B.n105 VSUBS 0.006472f
C218 B.n106 VSUBS 0.006472f
C219 B.n107 VSUBS 0.006472f
C220 B.n108 VSUBS 0.006472f
C221 B.n109 VSUBS 0.006472f
C222 B.n110 VSUBS 0.015932f
C223 B.n111 VSUBS 0.016619f
C224 B.n112 VSUBS 0.016619f
C225 B.n113 VSUBS 0.006472f
C226 B.n114 VSUBS 0.006472f
C227 B.n115 VSUBS 0.006472f
C228 B.n116 VSUBS 0.006472f
C229 B.n117 VSUBS 0.006472f
C230 B.n118 VSUBS 0.006472f
C231 B.n119 VSUBS 0.006472f
C232 B.n120 VSUBS 0.006472f
C233 B.n121 VSUBS 0.006472f
C234 B.n122 VSUBS 0.006472f
C235 B.n123 VSUBS 0.006472f
C236 B.n124 VSUBS 0.006472f
C237 B.n125 VSUBS 0.006472f
C238 B.n126 VSUBS 0.006472f
C239 B.n127 VSUBS 0.006472f
C240 B.n128 VSUBS 0.006472f
C241 B.n129 VSUBS 0.006472f
C242 B.n130 VSUBS 0.006472f
C243 B.n131 VSUBS 0.006472f
C244 B.n132 VSUBS 0.006472f
C245 B.n133 VSUBS 0.006472f
C246 B.n134 VSUBS 0.006472f
C247 B.n135 VSUBS 0.006472f
C248 B.n136 VSUBS 0.006472f
C249 B.n137 VSUBS 0.006472f
C250 B.n138 VSUBS 0.006472f
C251 B.n139 VSUBS 0.006472f
C252 B.n140 VSUBS 0.006472f
C253 B.n141 VSUBS 0.006472f
C254 B.n142 VSUBS 0.006472f
C255 B.n143 VSUBS 0.006472f
C256 B.n144 VSUBS 0.006472f
C257 B.n145 VSUBS 0.006472f
C258 B.n146 VSUBS 0.006472f
C259 B.n147 VSUBS 0.006472f
C260 B.n148 VSUBS 0.006472f
C261 B.n149 VSUBS 0.006472f
C262 B.n150 VSUBS 0.006472f
C263 B.n151 VSUBS 0.006472f
C264 B.n152 VSUBS 0.004283f
C265 B.n153 VSUBS 0.014995f
C266 B.n154 VSUBS 0.005425f
C267 B.n155 VSUBS 0.006472f
C268 B.n156 VSUBS 0.006472f
C269 B.n157 VSUBS 0.006472f
C270 B.n158 VSUBS 0.006472f
C271 B.n159 VSUBS 0.006472f
C272 B.n160 VSUBS 0.006472f
C273 B.n161 VSUBS 0.006472f
C274 B.n162 VSUBS 0.006472f
C275 B.n163 VSUBS 0.006472f
C276 B.n164 VSUBS 0.006472f
C277 B.n165 VSUBS 0.006472f
C278 B.t11 VSUBS 0.104749f
C279 B.t10 VSUBS 0.110537f
C280 B.t9 VSUBS 0.075858f
C281 B.n166 VSUBS 0.171421f
C282 B.n167 VSUBS 0.15754f
C283 B.n168 VSUBS 0.014995f
C284 B.n169 VSUBS 0.005425f
C285 B.n170 VSUBS 0.006472f
C286 B.n171 VSUBS 0.006472f
C287 B.n172 VSUBS 0.006472f
C288 B.n173 VSUBS 0.006472f
C289 B.n174 VSUBS 0.006472f
C290 B.n175 VSUBS 0.006472f
C291 B.n176 VSUBS 0.006472f
C292 B.n177 VSUBS 0.006472f
C293 B.n178 VSUBS 0.006472f
C294 B.n179 VSUBS 0.006472f
C295 B.n180 VSUBS 0.006472f
C296 B.n181 VSUBS 0.006472f
C297 B.n182 VSUBS 0.006472f
C298 B.n183 VSUBS 0.006472f
C299 B.n184 VSUBS 0.006472f
C300 B.n185 VSUBS 0.006472f
C301 B.n186 VSUBS 0.006472f
C302 B.n187 VSUBS 0.006472f
C303 B.n188 VSUBS 0.006472f
C304 B.n189 VSUBS 0.006472f
C305 B.n190 VSUBS 0.006472f
C306 B.n191 VSUBS 0.006472f
C307 B.n192 VSUBS 0.006472f
C308 B.n193 VSUBS 0.006472f
C309 B.n194 VSUBS 0.006472f
C310 B.n195 VSUBS 0.006472f
C311 B.n196 VSUBS 0.006472f
C312 B.n197 VSUBS 0.006472f
C313 B.n198 VSUBS 0.006472f
C314 B.n199 VSUBS 0.006472f
C315 B.n200 VSUBS 0.006472f
C316 B.n201 VSUBS 0.006472f
C317 B.n202 VSUBS 0.006472f
C318 B.n203 VSUBS 0.006472f
C319 B.n204 VSUBS 0.006472f
C320 B.n205 VSUBS 0.006472f
C321 B.n206 VSUBS 0.006472f
C322 B.n207 VSUBS 0.006472f
C323 B.n208 VSUBS 0.006472f
C324 B.n209 VSUBS 0.006472f
C325 B.n210 VSUBS 0.006472f
C326 B.n211 VSUBS 0.015932f
C327 B.n212 VSUBS 0.016619f
C328 B.n213 VSUBS 0.015932f
C329 B.n214 VSUBS 0.006472f
C330 B.n215 VSUBS 0.006472f
C331 B.n216 VSUBS 0.006472f
C332 B.n217 VSUBS 0.006472f
C333 B.n218 VSUBS 0.006472f
C334 B.n219 VSUBS 0.006472f
C335 B.n220 VSUBS 0.006472f
C336 B.n221 VSUBS 0.006472f
C337 B.n222 VSUBS 0.006472f
C338 B.n223 VSUBS 0.006472f
C339 B.n224 VSUBS 0.006472f
C340 B.n225 VSUBS 0.006472f
C341 B.n226 VSUBS 0.006472f
C342 B.n227 VSUBS 0.006472f
C343 B.n228 VSUBS 0.006472f
C344 B.n229 VSUBS 0.006472f
C345 B.n230 VSUBS 0.006472f
C346 B.n231 VSUBS 0.006472f
C347 B.n232 VSUBS 0.006472f
C348 B.n233 VSUBS 0.006472f
C349 B.n234 VSUBS 0.006472f
C350 B.n235 VSUBS 0.006472f
C351 B.n236 VSUBS 0.006472f
C352 B.n237 VSUBS 0.006472f
C353 B.n238 VSUBS 0.006472f
C354 B.n239 VSUBS 0.006472f
C355 B.n240 VSUBS 0.006472f
C356 B.n241 VSUBS 0.006472f
C357 B.n242 VSUBS 0.006472f
C358 B.n243 VSUBS 0.006472f
C359 B.n244 VSUBS 0.006472f
C360 B.n245 VSUBS 0.006472f
C361 B.n246 VSUBS 0.006472f
C362 B.n247 VSUBS 0.015932f
C363 B.n248 VSUBS 0.015932f
C364 B.n249 VSUBS 0.016619f
C365 B.n250 VSUBS 0.006472f
C366 B.n251 VSUBS 0.006472f
C367 B.n252 VSUBS 0.006472f
C368 B.n253 VSUBS 0.006472f
C369 B.n254 VSUBS 0.006472f
C370 B.n255 VSUBS 0.006472f
C371 B.n256 VSUBS 0.006472f
C372 B.n257 VSUBS 0.006472f
C373 B.n258 VSUBS 0.006472f
C374 B.n259 VSUBS 0.006472f
C375 B.n260 VSUBS 0.006472f
C376 B.n261 VSUBS 0.006472f
C377 B.n262 VSUBS 0.006472f
C378 B.n263 VSUBS 0.006472f
C379 B.n264 VSUBS 0.006472f
C380 B.n265 VSUBS 0.006472f
C381 B.n266 VSUBS 0.006472f
C382 B.n267 VSUBS 0.006472f
C383 B.n268 VSUBS 0.006472f
C384 B.n269 VSUBS 0.006472f
C385 B.n270 VSUBS 0.006472f
C386 B.n271 VSUBS 0.006472f
C387 B.n272 VSUBS 0.006472f
C388 B.n273 VSUBS 0.006472f
C389 B.n274 VSUBS 0.006472f
C390 B.n275 VSUBS 0.006472f
C391 B.n276 VSUBS 0.006472f
C392 B.n277 VSUBS 0.006472f
C393 B.n278 VSUBS 0.006472f
C394 B.n279 VSUBS 0.006472f
C395 B.n280 VSUBS 0.006472f
C396 B.n281 VSUBS 0.006472f
C397 B.n282 VSUBS 0.006472f
C398 B.n283 VSUBS 0.006472f
C399 B.n284 VSUBS 0.006472f
C400 B.n285 VSUBS 0.006472f
C401 B.n286 VSUBS 0.006472f
C402 B.n287 VSUBS 0.006472f
C403 B.n288 VSUBS 0.006472f
C404 B.n289 VSUBS 0.004283f
C405 B.n290 VSUBS 0.006472f
C406 B.n291 VSUBS 0.006472f
C407 B.n292 VSUBS 0.005425f
C408 B.n293 VSUBS 0.006472f
C409 B.n294 VSUBS 0.006472f
C410 B.n295 VSUBS 0.006472f
C411 B.n296 VSUBS 0.006472f
C412 B.n297 VSUBS 0.006472f
C413 B.n298 VSUBS 0.006472f
C414 B.n299 VSUBS 0.006472f
C415 B.n300 VSUBS 0.006472f
C416 B.n301 VSUBS 0.006472f
C417 B.n302 VSUBS 0.006472f
C418 B.n303 VSUBS 0.006472f
C419 B.n304 VSUBS 0.005425f
C420 B.n305 VSUBS 0.014995f
C421 B.n306 VSUBS 0.004283f
C422 B.n307 VSUBS 0.006472f
C423 B.n308 VSUBS 0.006472f
C424 B.n309 VSUBS 0.006472f
C425 B.n310 VSUBS 0.006472f
C426 B.n311 VSUBS 0.006472f
C427 B.n312 VSUBS 0.006472f
C428 B.n313 VSUBS 0.006472f
C429 B.n314 VSUBS 0.006472f
C430 B.n315 VSUBS 0.006472f
C431 B.n316 VSUBS 0.006472f
C432 B.n317 VSUBS 0.006472f
C433 B.n318 VSUBS 0.006472f
C434 B.n319 VSUBS 0.006472f
C435 B.n320 VSUBS 0.006472f
C436 B.n321 VSUBS 0.006472f
C437 B.n322 VSUBS 0.006472f
C438 B.n323 VSUBS 0.006472f
C439 B.n324 VSUBS 0.006472f
C440 B.n325 VSUBS 0.006472f
C441 B.n326 VSUBS 0.006472f
C442 B.n327 VSUBS 0.006472f
C443 B.n328 VSUBS 0.006472f
C444 B.n329 VSUBS 0.006472f
C445 B.n330 VSUBS 0.006472f
C446 B.n331 VSUBS 0.006472f
C447 B.n332 VSUBS 0.006472f
C448 B.n333 VSUBS 0.006472f
C449 B.n334 VSUBS 0.006472f
C450 B.n335 VSUBS 0.006472f
C451 B.n336 VSUBS 0.006472f
C452 B.n337 VSUBS 0.006472f
C453 B.n338 VSUBS 0.006472f
C454 B.n339 VSUBS 0.006472f
C455 B.n340 VSUBS 0.006472f
C456 B.n341 VSUBS 0.006472f
C457 B.n342 VSUBS 0.006472f
C458 B.n343 VSUBS 0.006472f
C459 B.n344 VSUBS 0.006472f
C460 B.n345 VSUBS 0.006472f
C461 B.n346 VSUBS 0.016619f
C462 B.n347 VSUBS 0.016619f
C463 B.n348 VSUBS 0.015932f
C464 B.n349 VSUBS 0.006472f
C465 B.n350 VSUBS 0.006472f
C466 B.n351 VSUBS 0.006472f
C467 B.n352 VSUBS 0.006472f
C468 B.n353 VSUBS 0.006472f
C469 B.n354 VSUBS 0.006472f
C470 B.n355 VSUBS 0.006472f
C471 B.n356 VSUBS 0.006472f
C472 B.n357 VSUBS 0.006472f
C473 B.n358 VSUBS 0.006472f
C474 B.n359 VSUBS 0.006472f
C475 B.n360 VSUBS 0.006472f
C476 B.n361 VSUBS 0.006472f
C477 B.n362 VSUBS 0.006472f
C478 B.n363 VSUBS 0.008446f
C479 B.n364 VSUBS 0.008997f
C480 B.n365 VSUBS 0.017891f
C481 VDD2.n0 VSUBS 0.021976f
C482 VDD2.n1 VSUBS 0.019661f
C483 VDD2.n2 VSUBS 0.010565f
C484 VDD2.n3 VSUBS 0.024971f
C485 VDD2.n4 VSUBS 0.011186f
C486 VDD2.n5 VSUBS 0.019661f
C487 VDD2.n6 VSUBS 0.010565f
C488 VDD2.n7 VSUBS 0.024971f
C489 VDD2.n8 VSUBS 0.011186f
C490 VDD2.n9 VSUBS 0.561641f
C491 VDD2.n10 VSUBS 0.010565f
C492 VDD2.t1 VSUBS 0.053676f
C493 VDD2.n11 VSUBS 0.113294f
C494 VDD2.n12 VSUBS 0.018784f
C495 VDD2.n13 VSUBS 0.018728f
C496 VDD2.n14 VSUBS 0.024971f
C497 VDD2.n15 VSUBS 0.011186f
C498 VDD2.n16 VSUBS 0.010565f
C499 VDD2.n17 VSUBS 0.019661f
C500 VDD2.n18 VSUBS 0.019661f
C501 VDD2.n19 VSUBS 0.010565f
C502 VDD2.n20 VSUBS 0.011186f
C503 VDD2.n21 VSUBS 0.024971f
C504 VDD2.n22 VSUBS 0.024971f
C505 VDD2.n23 VSUBS 0.011186f
C506 VDD2.n24 VSUBS 0.010565f
C507 VDD2.n25 VSUBS 0.019661f
C508 VDD2.n26 VSUBS 0.019661f
C509 VDD2.n27 VSUBS 0.010565f
C510 VDD2.n28 VSUBS 0.011186f
C511 VDD2.n29 VSUBS 0.024971f
C512 VDD2.n30 VSUBS 0.063482f
C513 VDD2.n31 VSUBS 0.011186f
C514 VDD2.n32 VSUBS 0.020747f
C515 VDD2.n33 VSUBS 0.051622f
C516 VDD2.n34 VSUBS 0.352582f
C517 VDD2.n35 VSUBS 0.021976f
C518 VDD2.n36 VSUBS 0.019661f
C519 VDD2.n37 VSUBS 0.010565f
C520 VDD2.n38 VSUBS 0.024971f
C521 VDD2.n39 VSUBS 0.011186f
C522 VDD2.n40 VSUBS 0.019661f
C523 VDD2.n41 VSUBS 0.010565f
C524 VDD2.n42 VSUBS 0.024971f
C525 VDD2.n43 VSUBS 0.011186f
C526 VDD2.n44 VSUBS 0.561641f
C527 VDD2.n45 VSUBS 0.010565f
C528 VDD2.t0 VSUBS 0.053676f
C529 VDD2.n46 VSUBS 0.113294f
C530 VDD2.n47 VSUBS 0.018784f
C531 VDD2.n48 VSUBS 0.018728f
C532 VDD2.n49 VSUBS 0.024971f
C533 VDD2.n50 VSUBS 0.011186f
C534 VDD2.n51 VSUBS 0.010565f
C535 VDD2.n52 VSUBS 0.019661f
C536 VDD2.n53 VSUBS 0.019661f
C537 VDD2.n54 VSUBS 0.010565f
C538 VDD2.n55 VSUBS 0.011186f
C539 VDD2.n56 VSUBS 0.024971f
C540 VDD2.n57 VSUBS 0.024971f
C541 VDD2.n58 VSUBS 0.011186f
C542 VDD2.n59 VSUBS 0.010565f
C543 VDD2.n60 VSUBS 0.019661f
C544 VDD2.n61 VSUBS 0.019661f
C545 VDD2.n62 VSUBS 0.010565f
C546 VDD2.n63 VSUBS 0.011186f
C547 VDD2.n64 VSUBS 0.024971f
C548 VDD2.n65 VSUBS 0.063482f
C549 VDD2.n66 VSUBS 0.011186f
C550 VDD2.n67 VSUBS 0.020747f
C551 VDD2.n68 VSUBS 0.051622f
C552 VDD2.n69 VSUBS 0.062937f
C553 VDD2.n70 VSUBS 1.66727f
C554 VTAIL.n0 VSUBS 0.029521f
C555 VTAIL.n1 VSUBS 0.02641f
C556 VTAIL.n2 VSUBS 0.014192f
C557 VTAIL.n3 VSUBS 0.033544f
C558 VTAIL.n4 VSUBS 0.015027f
C559 VTAIL.n5 VSUBS 0.02641f
C560 VTAIL.n6 VSUBS 0.014192f
C561 VTAIL.n7 VSUBS 0.033544f
C562 VTAIL.n8 VSUBS 0.015027f
C563 VTAIL.n9 VSUBS 0.754458f
C564 VTAIL.n10 VSUBS 0.014192f
C565 VTAIL.t0 VSUBS 0.072104f
C566 VTAIL.n11 VSUBS 0.152188f
C567 VTAIL.n12 VSUBS 0.025232f
C568 VTAIL.n13 VSUBS 0.025158f
C569 VTAIL.n14 VSUBS 0.033544f
C570 VTAIL.n15 VSUBS 0.015027f
C571 VTAIL.n16 VSUBS 0.014192f
C572 VTAIL.n17 VSUBS 0.02641f
C573 VTAIL.n18 VSUBS 0.02641f
C574 VTAIL.n19 VSUBS 0.014192f
C575 VTAIL.n20 VSUBS 0.015027f
C576 VTAIL.n21 VSUBS 0.033544f
C577 VTAIL.n22 VSUBS 0.033544f
C578 VTAIL.n23 VSUBS 0.015027f
C579 VTAIL.n24 VSUBS 0.014192f
C580 VTAIL.n25 VSUBS 0.02641f
C581 VTAIL.n26 VSUBS 0.02641f
C582 VTAIL.n27 VSUBS 0.014192f
C583 VTAIL.n28 VSUBS 0.015027f
C584 VTAIL.n29 VSUBS 0.033544f
C585 VTAIL.n30 VSUBS 0.085275f
C586 VTAIL.n31 VSUBS 0.015027f
C587 VTAIL.n32 VSUBS 0.027869f
C588 VTAIL.n33 VSUBS 0.069344f
C589 VTAIL.n34 VSUBS 0.066364f
C590 VTAIL.n35 VSUBS 1.06937f
C591 VTAIL.n36 VSUBS 0.029521f
C592 VTAIL.n37 VSUBS 0.02641f
C593 VTAIL.n38 VSUBS 0.014192f
C594 VTAIL.n39 VSUBS 0.033544f
C595 VTAIL.n40 VSUBS 0.015027f
C596 VTAIL.n41 VSUBS 0.02641f
C597 VTAIL.n42 VSUBS 0.014192f
C598 VTAIL.n43 VSUBS 0.033544f
C599 VTAIL.n44 VSUBS 0.015027f
C600 VTAIL.n45 VSUBS 0.754458f
C601 VTAIL.n46 VSUBS 0.014192f
C602 VTAIL.t3 VSUBS 0.072104f
C603 VTAIL.n47 VSUBS 0.152188f
C604 VTAIL.n48 VSUBS 0.025232f
C605 VTAIL.n49 VSUBS 0.025158f
C606 VTAIL.n50 VSUBS 0.033544f
C607 VTAIL.n51 VSUBS 0.015027f
C608 VTAIL.n52 VSUBS 0.014192f
C609 VTAIL.n53 VSUBS 0.02641f
C610 VTAIL.n54 VSUBS 0.02641f
C611 VTAIL.n55 VSUBS 0.014192f
C612 VTAIL.n56 VSUBS 0.015027f
C613 VTAIL.n57 VSUBS 0.033544f
C614 VTAIL.n58 VSUBS 0.033544f
C615 VTAIL.n59 VSUBS 0.015027f
C616 VTAIL.n60 VSUBS 0.014192f
C617 VTAIL.n61 VSUBS 0.02641f
C618 VTAIL.n62 VSUBS 0.02641f
C619 VTAIL.n63 VSUBS 0.014192f
C620 VTAIL.n64 VSUBS 0.015027f
C621 VTAIL.n65 VSUBS 0.033544f
C622 VTAIL.n66 VSUBS 0.085275f
C623 VTAIL.n67 VSUBS 0.015027f
C624 VTAIL.n68 VSUBS 0.027869f
C625 VTAIL.n69 VSUBS 0.069344f
C626 VTAIL.n70 VSUBS 0.066364f
C627 VTAIL.n71 VSUBS 1.07561f
C628 VTAIL.n72 VSUBS 0.029521f
C629 VTAIL.n73 VSUBS 0.02641f
C630 VTAIL.n74 VSUBS 0.014192f
C631 VTAIL.n75 VSUBS 0.033544f
C632 VTAIL.n76 VSUBS 0.015027f
C633 VTAIL.n77 VSUBS 0.02641f
C634 VTAIL.n78 VSUBS 0.014192f
C635 VTAIL.n79 VSUBS 0.033544f
C636 VTAIL.n80 VSUBS 0.015027f
C637 VTAIL.n81 VSUBS 0.754458f
C638 VTAIL.n82 VSUBS 0.014192f
C639 VTAIL.t1 VSUBS 0.072104f
C640 VTAIL.n83 VSUBS 0.152188f
C641 VTAIL.n84 VSUBS 0.025232f
C642 VTAIL.n85 VSUBS 0.025158f
C643 VTAIL.n86 VSUBS 0.033544f
C644 VTAIL.n87 VSUBS 0.015027f
C645 VTAIL.n88 VSUBS 0.014192f
C646 VTAIL.n89 VSUBS 0.02641f
C647 VTAIL.n90 VSUBS 0.02641f
C648 VTAIL.n91 VSUBS 0.014192f
C649 VTAIL.n92 VSUBS 0.015027f
C650 VTAIL.n93 VSUBS 0.033544f
C651 VTAIL.n94 VSUBS 0.033544f
C652 VTAIL.n95 VSUBS 0.015027f
C653 VTAIL.n96 VSUBS 0.014192f
C654 VTAIL.n97 VSUBS 0.02641f
C655 VTAIL.n98 VSUBS 0.02641f
C656 VTAIL.n99 VSUBS 0.014192f
C657 VTAIL.n100 VSUBS 0.015027f
C658 VTAIL.n101 VSUBS 0.033544f
C659 VTAIL.n102 VSUBS 0.085275f
C660 VTAIL.n103 VSUBS 0.015027f
C661 VTAIL.n104 VSUBS 0.027869f
C662 VTAIL.n105 VSUBS 0.069344f
C663 VTAIL.n106 VSUBS 0.066364f
C664 VTAIL.n107 VSUBS 1.03086f
C665 VTAIL.n108 VSUBS 0.029521f
C666 VTAIL.n109 VSUBS 0.02641f
C667 VTAIL.n110 VSUBS 0.014192f
C668 VTAIL.n111 VSUBS 0.033544f
C669 VTAIL.n112 VSUBS 0.015027f
C670 VTAIL.n113 VSUBS 0.02641f
C671 VTAIL.n114 VSUBS 0.014192f
C672 VTAIL.n115 VSUBS 0.033544f
C673 VTAIL.n116 VSUBS 0.015027f
C674 VTAIL.n117 VSUBS 0.754458f
C675 VTAIL.n118 VSUBS 0.014192f
C676 VTAIL.t2 VSUBS 0.072104f
C677 VTAIL.n119 VSUBS 0.152188f
C678 VTAIL.n120 VSUBS 0.025232f
C679 VTAIL.n121 VSUBS 0.025158f
C680 VTAIL.n122 VSUBS 0.033544f
C681 VTAIL.n123 VSUBS 0.015027f
C682 VTAIL.n124 VSUBS 0.014192f
C683 VTAIL.n125 VSUBS 0.02641f
C684 VTAIL.n126 VSUBS 0.02641f
C685 VTAIL.n127 VSUBS 0.014192f
C686 VTAIL.n128 VSUBS 0.015027f
C687 VTAIL.n129 VSUBS 0.033544f
C688 VTAIL.n130 VSUBS 0.033544f
C689 VTAIL.n131 VSUBS 0.015027f
C690 VTAIL.n132 VSUBS 0.014192f
C691 VTAIL.n133 VSUBS 0.02641f
C692 VTAIL.n134 VSUBS 0.02641f
C693 VTAIL.n135 VSUBS 0.014192f
C694 VTAIL.n136 VSUBS 0.015027f
C695 VTAIL.n137 VSUBS 0.033544f
C696 VTAIL.n138 VSUBS 0.085275f
C697 VTAIL.n139 VSUBS 0.015027f
C698 VTAIL.n140 VSUBS 0.027869f
C699 VTAIL.n141 VSUBS 0.069344f
C700 VTAIL.n142 VSUBS 0.066364f
C701 VTAIL.n143 VSUBS 0.974735f
C702 VN.t0 VSUBS 0.282158f
C703 VN.t1 VSUBS 0.335135f
.ends

