* NGSPICE file created from diff_pair_sample_1159.ext - technology: sky130A

.subckt diff_pair_sample_1159 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=1.06
X1 VDD2.t9 VN.t0 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=1.06
X2 VTAIL.t11 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X3 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=1.06
X4 VTAIL.t0 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X5 VTAIL.t9 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X6 VDD1.t6 VP.t3 VTAIL.t14 B.t8 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X7 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=1.06
X8 VTAIL.t7 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X9 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=1.06
X10 VTAIL.t10 VP.t4 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X11 VDD2.t5 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=1.06
X12 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=1.06
X13 VTAIL.t18 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X14 VDD1.t3 VP.t6 VTAIL.t17 B.t5 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X15 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=1.06
X16 VDD1.t2 VP.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=1.06
X17 VDD1.t1 VP.t8 VTAIL.t15 B.t1 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=1.06
X18 VDD1.t0 VP.t9 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=1.06
X19 VTAIL.t4 VN.t6 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X20 VTAIL.t2 VN.t7 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X21 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=1.06
X22 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
X23 VDD2.t0 VN.t9 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=1.06
R0 VP.n10 VP.t0 294.608
R1 VP.n5 VP.t7 274.423
R2 VP.n41 VP.t8 274.423
R3 VP.n23 VP.t9 274.423
R4 VP.n34 VP.t3 237.136
R5 VP.n29 VP.t1 237.136
R6 VP.n1 VP.t5 237.136
R7 VP.n16 VP.t6 237.136
R8 VP.n7 VP.t4 237.136
R9 VP.n11 VP.t2 237.136
R10 VP.n13 VP.n12 161.3
R11 VP.n14 VP.n9 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n8 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n22 VP.n6 161.3
R17 VP.n40 VP.n0 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n2 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n3 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n28 VP.n4 161.3
R25 VP.n27 VP.n26 161.3
R26 VP.n24 VP.n23 80.6037
R27 VP.n42 VP.n41 80.6037
R28 VP.n25 VP.n5 80.6037
R29 VP.n30 VP.n3 56.5193
R30 VP.n36 VP.n35 56.5193
R31 VP.n18 VP.n17 56.5193
R32 VP.n12 VP.n9 56.5193
R33 VP.n25 VP.n24 43.6188
R34 VP.n11 VP.n10 38.2823
R35 VP.n27 VP.n5 36.5157
R36 VP.n41 VP.n40 36.5157
R37 VP.n23 VP.n22 36.5157
R38 VP.n28 VP.n27 32.2376
R39 VP.n40 VP.n39 32.2376
R40 VP.n22 VP.n21 32.2376
R41 VP.n13 VP.n10 29.1642
R42 VP.n34 VP.n3 24.4675
R43 VP.n35 VP.n34 24.4675
R44 VP.n16 VP.n9 24.4675
R45 VP.n17 VP.n16 24.4675
R46 VP.n30 VP.n29 19.0848
R47 VP.n36 VP.n1 19.0848
R48 VP.n18 VP.n7 19.0848
R49 VP.n12 VP.n11 19.0848
R50 VP.n29 VP.n28 5.38324
R51 VP.n39 VP.n1 5.38324
R52 VP.n21 VP.n7 5.38324
R53 VP.n24 VP.n6 0.285035
R54 VP.n26 VP.n25 0.285035
R55 VP.n42 VP.n0 0.285035
R56 VP.n14 VP.n13 0.189894
R57 VP.n15 VP.n14 0.189894
R58 VP.n15 VP.n8 0.189894
R59 VP.n19 VP.n8 0.189894
R60 VP.n20 VP.n19 0.189894
R61 VP.n20 VP.n6 0.189894
R62 VP.n26 VP.n4 0.189894
R63 VP.n31 VP.n4 0.189894
R64 VP.n32 VP.n31 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n33 VP.n2 0.189894
R67 VP.n37 VP.n2 0.189894
R68 VP.n38 VP.n37 0.189894
R69 VP.n38 VP.n0 0.189894
R70 VP VP.n42 0.146778
R71 VTAIL.n11 VTAIL.t1 49.8359
R72 VTAIL.n17 VTAIL.t6 49.8357
R73 VTAIL.n2 VTAIL.t15 49.8357
R74 VTAIL.n16 VTAIL.t12 49.8357
R75 VTAIL.n15 VTAIL.n14 47.9375
R76 VTAIL.n13 VTAIL.n12 47.9375
R77 VTAIL.n10 VTAIL.n9 47.9375
R78 VTAIL.n8 VTAIL.n7 47.9375
R79 VTAIL.n19 VTAIL.n18 47.9373
R80 VTAIL.n1 VTAIL.n0 47.9373
R81 VTAIL.n4 VTAIL.n3 47.9373
R82 VTAIL.n6 VTAIL.n5 47.9373
R83 VTAIL.n8 VTAIL.n6 23.7548
R84 VTAIL.n17 VTAIL.n16 22.5565
R85 VTAIL.n18 VTAIL.t5 1.89887
R86 VTAIL.n18 VTAIL.t7 1.89887
R87 VTAIL.n0 VTAIL.t19 1.89887
R88 VTAIL.n0 VTAIL.t4 1.89887
R89 VTAIL.n3 VTAIL.t14 1.89887
R90 VTAIL.n3 VTAIL.t18 1.89887
R91 VTAIL.n5 VTAIL.t13 1.89887
R92 VTAIL.n5 VTAIL.t11 1.89887
R93 VTAIL.n14 VTAIL.t17 1.89887
R94 VTAIL.n14 VTAIL.t10 1.89887
R95 VTAIL.n12 VTAIL.t16 1.89887
R96 VTAIL.n12 VTAIL.t9 1.89887
R97 VTAIL.n9 VTAIL.t8 1.89887
R98 VTAIL.n9 VTAIL.t2 1.89887
R99 VTAIL.n7 VTAIL.t3 1.89887
R100 VTAIL.n7 VTAIL.t0 1.89887
R101 VTAIL.n10 VTAIL.n8 1.19878
R102 VTAIL.n11 VTAIL.n10 1.19878
R103 VTAIL.n15 VTAIL.n13 1.19878
R104 VTAIL.n16 VTAIL.n15 1.19878
R105 VTAIL.n6 VTAIL.n4 1.19878
R106 VTAIL.n4 VTAIL.n2 1.19878
R107 VTAIL.n19 VTAIL.n17 1.19878
R108 VTAIL.n13 VTAIL.n11 1.06947
R109 VTAIL.n2 VTAIL.n1 1.06947
R110 VTAIL VTAIL.n1 0.957397
R111 VTAIL VTAIL.n19 0.241879
R112 VDD1.n1 VDD1.t9 67.713
R113 VDD1.n3 VDD1.t2 67.7127
R114 VDD1.n5 VDD1.n4 65.4594
R115 VDD1.n1 VDD1.n0 64.6163
R116 VDD1.n7 VDD1.n6 64.6162
R117 VDD1.n3 VDD1.n2 64.6161
R118 VDD1.n7 VDD1.n5 39.5806
R119 VDD1.n6 VDD1.t5 1.89887
R120 VDD1.n6 VDD1.t0 1.89887
R121 VDD1.n0 VDD1.t7 1.89887
R122 VDD1.n0 VDD1.t3 1.89887
R123 VDD1.n4 VDD1.t4 1.89887
R124 VDD1.n4 VDD1.t1 1.89887
R125 VDD1.n2 VDD1.t8 1.89887
R126 VDD1.n2 VDD1.t6 1.89887
R127 VDD1 VDD1.n7 0.841017
R128 VDD1 VDD1.n1 0.358259
R129 VDD1.n5 VDD1.n3 0.244723
R130 B.n691 B.n690 585
R131 B.n272 B.n103 585
R132 B.n271 B.n270 585
R133 B.n269 B.n268 585
R134 B.n267 B.n266 585
R135 B.n265 B.n264 585
R136 B.n263 B.n262 585
R137 B.n261 B.n260 585
R138 B.n259 B.n258 585
R139 B.n257 B.n256 585
R140 B.n255 B.n254 585
R141 B.n253 B.n252 585
R142 B.n251 B.n250 585
R143 B.n249 B.n248 585
R144 B.n247 B.n246 585
R145 B.n245 B.n244 585
R146 B.n243 B.n242 585
R147 B.n241 B.n240 585
R148 B.n239 B.n238 585
R149 B.n237 B.n236 585
R150 B.n235 B.n234 585
R151 B.n233 B.n232 585
R152 B.n231 B.n230 585
R153 B.n229 B.n228 585
R154 B.n227 B.n226 585
R155 B.n225 B.n224 585
R156 B.n223 B.n222 585
R157 B.n221 B.n220 585
R158 B.n219 B.n218 585
R159 B.n217 B.n216 585
R160 B.n215 B.n214 585
R161 B.n213 B.n212 585
R162 B.n211 B.n210 585
R163 B.n209 B.n208 585
R164 B.n207 B.n206 585
R165 B.n205 B.n204 585
R166 B.n203 B.n202 585
R167 B.n200 B.n199 585
R168 B.n198 B.n197 585
R169 B.n196 B.n195 585
R170 B.n194 B.n193 585
R171 B.n192 B.n191 585
R172 B.n190 B.n189 585
R173 B.n188 B.n187 585
R174 B.n186 B.n185 585
R175 B.n184 B.n183 585
R176 B.n182 B.n181 585
R177 B.n179 B.n178 585
R178 B.n177 B.n176 585
R179 B.n175 B.n174 585
R180 B.n173 B.n172 585
R181 B.n171 B.n170 585
R182 B.n169 B.n168 585
R183 B.n167 B.n166 585
R184 B.n165 B.n164 585
R185 B.n163 B.n162 585
R186 B.n161 B.n160 585
R187 B.n159 B.n158 585
R188 B.n157 B.n156 585
R189 B.n155 B.n154 585
R190 B.n153 B.n152 585
R191 B.n151 B.n150 585
R192 B.n149 B.n148 585
R193 B.n147 B.n146 585
R194 B.n145 B.n144 585
R195 B.n143 B.n142 585
R196 B.n141 B.n140 585
R197 B.n139 B.n138 585
R198 B.n137 B.n136 585
R199 B.n135 B.n134 585
R200 B.n133 B.n132 585
R201 B.n131 B.n130 585
R202 B.n129 B.n128 585
R203 B.n127 B.n126 585
R204 B.n125 B.n124 585
R205 B.n123 B.n122 585
R206 B.n121 B.n120 585
R207 B.n119 B.n118 585
R208 B.n117 B.n116 585
R209 B.n115 B.n114 585
R210 B.n113 B.n112 585
R211 B.n111 B.n110 585
R212 B.n109 B.n108 585
R213 B.n60 B.n59 585
R214 B.n689 B.n61 585
R215 B.n694 B.n61 585
R216 B.n688 B.n687 585
R217 B.n687 B.n57 585
R218 B.n686 B.n56 585
R219 B.n700 B.n56 585
R220 B.n685 B.n55 585
R221 B.n701 B.n55 585
R222 B.n684 B.n54 585
R223 B.n702 B.n54 585
R224 B.n683 B.n682 585
R225 B.n682 B.n53 585
R226 B.n681 B.n49 585
R227 B.n708 B.n49 585
R228 B.n680 B.n48 585
R229 B.n709 B.n48 585
R230 B.n679 B.n47 585
R231 B.n710 B.n47 585
R232 B.n678 B.n677 585
R233 B.n677 B.n43 585
R234 B.n676 B.n42 585
R235 B.n716 B.n42 585
R236 B.n675 B.n41 585
R237 B.n717 B.n41 585
R238 B.n674 B.n40 585
R239 B.n718 B.n40 585
R240 B.n673 B.n672 585
R241 B.n672 B.n36 585
R242 B.n671 B.n35 585
R243 B.n724 B.n35 585
R244 B.n670 B.n34 585
R245 B.n725 B.n34 585
R246 B.n669 B.n33 585
R247 B.n726 B.n33 585
R248 B.n668 B.n667 585
R249 B.n667 B.n29 585
R250 B.n666 B.n28 585
R251 B.n732 B.n28 585
R252 B.n665 B.n27 585
R253 B.n733 B.n27 585
R254 B.n664 B.n26 585
R255 B.n734 B.n26 585
R256 B.n663 B.n662 585
R257 B.n662 B.n22 585
R258 B.n661 B.n21 585
R259 B.n740 B.n21 585
R260 B.n660 B.n20 585
R261 B.n741 B.n20 585
R262 B.n659 B.n19 585
R263 B.n742 B.n19 585
R264 B.n658 B.n657 585
R265 B.n657 B.n15 585
R266 B.n656 B.n14 585
R267 B.n748 B.n14 585
R268 B.n655 B.n13 585
R269 B.n749 B.n13 585
R270 B.n654 B.n12 585
R271 B.n750 B.n12 585
R272 B.n653 B.n652 585
R273 B.n652 B.n651 585
R274 B.n650 B.n649 585
R275 B.n650 B.n8 585
R276 B.n648 B.n7 585
R277 B.n757 B.n7 585
R278 B.n647 B.n6 585
R279 B.n758 B.n6 585
R280 B.n646 B.n5 585
R281 B.n759 B.n5 585
R282 B.n645 B.n644 585
R283 B.n644 B.n4 585
R284 B.n643 B.n273 585
R285 B.n643 B.n642 585
R286 B.n633 B.n274 585
R287 B.n275 B.n274 585
R288 B.n635 B.n634 585
R289 B.n636 B.n635 585
R290 B.n632 B.n280 585
R291 B.n280 B.n279 585
R292 B.n631 B.n630 585
R293 B.n630 B.n629 585
R294 B.n282 B.n281 585
R295 B.n283 B.n282 585
R296 B.n622 B.n621 585
R297 B.n623 B.n622 585
R298 B.n620 B.n288 585
R299 B.n288 B.n287 585
R300 B.n619 B.n618 585
R301 B.n618 B.n617 585
R302 B.n290 B.n289 585
R303 B.n291 B.n290 585
R304 B.n610 B.n609 585
R305 B.n611 B.n610 585
R306 B.n608 B.n296 585
R307 B.n296 B.n295 585
R308 B.n607 B.n606 585
R309 B.n606 B.n605 585
R310 B.n298 B.n297 585
R311 B.n299 B.n298 585
R312 B.n598 B.n597 585
R313 B.n599 B.n598 585
R314 B.n596 B.n304 585
R315 B.n304 B.n303 585
R316 B.n595 B.n594 585
R317 B.n594 B.n593 585
R318 B.n306 B.n305 585
R319 B.n307 B.n306 585
R320 B.n586 B.n585 585
R321 B.n587 B.n586 585
R322 B.n584 B.n312 585
R323 B.n312 B.n311 585
R324 B.n583 B.n582 585
R325 B.n582 B.n581 585
R326 B.n314 B.n313 585
R327 B.n315 B.n314 585
R328 B.n574 B.n573 585
R329 B.n575 B.n574 585
R330 B.n572 B.n320 585
R331 B.n320 B.n319 585
R332 B.n571 B.n570 585
R333 B.n570 B.n569 585
R334 B.n322 B.n321 585
R335 B.n562 B.n322 585
R336 B.n561 B.n560 585
R337 B.n563 B.n561 585
R338 B.n559 B.n327 585
R339 B.n327 B.n326 585
R340 B.n558 B.n557 585
R341 B.n557 B.n556 585
R342 B.n329 B.n328 585
R343 B.n330 B.n329 585
R344 B.n549 B.n548 585
R345 B.n550 B.n549 585
R346 B.n333 B.n332 585
R347 B.n384 B.n383 585
R348 B.n385 B.n381 585
R349 B.n381 B.n334 585
R350 B.n387 B.n386 585
R351 B.n389 B.n380 585
R352 B.n392 B.n391 585
R353 B.n393 B.n379 585
R354 B.n395 B.n394 585
R355 B.n397 B.n378 585
R356 B.n400 B.n399 585
R357 B.n401 B.n377 585
R358 B.n403 B.n402 585
R359 B.n405 B.n376 585
R360 B.n408 B.n407 585
R361 B.n409 B.n375 585
R362 B.n411 B.n410 585
R363 B.n413 B.n374 585
R364 B.n416 B.n415 585
R365 B.n417 B.n373 585
R366 B.n419 B.n418 585
R367 B.n421 B.n372 585
R368 B.n424 B.n423 585
R369 B.n425 B.n371 585
R370 B.n427 B.n426 585
R371 B.n429 B.n370 585
R372 B.n432 B.n431 585
R373 B.n433 B.n369 585
R374 B.n435 B.n434 585
R375 B.n437 B.n368 585
R376 B.n440 B.n439 585
R377 B.n441 B.n367 585
R378 B.n443 B.n442 585
R379 B.n445 B.n366 585
R380 B.n448 B.n447 585
R381 B.n449 B.n365 585
R382 B.n451 B.n450 585
R383 B.n453 B.n364 585
R384 B.n456 B.n455 585
R385 B.n457 B.n360 585
R386 B.n459 B.n458 585
R387 B.n461 B.n359 585
R388 B.n464 B.n463 585
R389 B.n465 B.n358 585
R390 B.n467 B.n466 585
R391 B.n469 B.n357 585
R392 B.n472 B.n471 585
R393 B.n473 B.n354 585
R394 B.n476 B.n475 585
R395 B.n478 B.n353 585
R396 B.n481 B.n480 585
R397 B.n482 B.n352 585
R398 B.n484 B.n483 585
R399 B.n486 B.n351 585
R400 B.n489 B.n488 585
R401 B.n490 B.n350 585
R402 B.n492 B.n491 585
R403 B.n494 B.n349 585
R404 B.n497 B.n496 585
R405 B.n498 B.n348 585
R406 B.n500 B.n499 585
R407 B.n502 B.n347 585
R408 B.n505 B.n504 585
R409 B.n506 B.n346 585
R410 B.n508 B.n507 585
R411 B.n510 B.n345 585
R412 B.n513 B.n512 585
R413 B.n514 B.n344 585
R414 B.n516 B.n515 585
R415 B.n518 B.n343 585
R416 B.n521 B.n520 585
R417 B.n522 B.n342 585
R418 B.n524 B.n523 585
R419 B.n526 B.n341 585
R420 B.n529 B.n528 585
R421 B.n530 B.n340 585
R422 B.n532 B.n531 585
R423 B.n534 B.n339 585
R424 B.n537 B.n536 585
R425 B.n538 B.n338 585
R426 B.n540 B.n539 585
R427 B.n542 B.n337 585
R428 B.n543 B.n336 585
R429 B.n546 B.n545 585
R430 B.n547 B.n335 585
R431 B.n335 B.n334 585
R432 B.n552 B.n551 585
R433 B.n551 B.n550 585
R434 B.n553 B.n331 585
R435 B.n331 B.n330 585
R436 B.n555 B.n554 585
R437 B.n556 B.n555 585
R438 B.n325 B.n324 585
R439 B.n326 B.n325 585
R440 B.n565 B.n564 585
R441 B.n564 B.n563 585
R442 B.n566 B.n323 585
R443 B.n562 B.n323 585
R444 B.n568 B.n567 585
R445 B.n569 B.n568 585
R446 B.n318 B.n317 585
R447 B.n319 B.n318 585
R448 B.n577 B.n576 585
R449 B.n576 B.n575 585
R450 B.n578 B.n316 585
R451 B.n316 B.n315 585
R452 B.n580 B.n579 585
R453 B.n581 B.n580 585
R454 B.n310 B.n309 585
R455 B.n311 B.n310 585
R456 B.n589 B.n588 585
R457 B.n588 B.n587 585
R458 B.n590 B.n308 585
R459 B.n308 B.n307 585
R460 B.n592 B.n591 585
R461 B.n593 B.n592 585
R462 B.n302 B.n301 585
R463 B.n303 B.n302 585
R464 B.n601 B.n600 585
R465 B.n600 B.n599 585
R466 B.n602 B.n300 585
R467 B.n300 B.n299 585
R468 B.n604 B.n603 585
R469 B.n605 B.n604 585
R470 B.n294 B.n293 585
R471 B.n295 B.n294 585
R472 B.n613 B.n612 585
R473 B.n612 B.n611 585
R474 B.n614 B.n292 585
R475 B.n292 B.n291 585
R476 B.n616 B.n615 585
R477 B.n617 B.n616 585
R478 B.n286 B.n285 585
R479 B.n287 B.n286 585
R480 B.n625 B.n624 585
R481 B.n624 B.n623 585
R482 B.n626 B.n284 585
R483 B.n284 B.n283 585
R484 B.n628 B.n627 585
R485 B.n629 B.n628 585
R486 B.n278 B.n277 585
R487 B.n279 B.n278 585
R488 B.n638 B.n637 585
R489 B.n637 B.n636 585
R490 B.n639 B.n276 585
R491 B.n276 B.n275 585
R492 B.n641 B.n640 585
R493 B.n642 B.n641 585
R494 B.n3 B.n0 585
R495 B.n4 B.n3 585
R496 B.n756 B.n1 585
R497 B.n757 B.n756 585
R498 B.n755 B.n754 585
R499 B.n755 B.n8 585
R500 B.n753 B.n9 585
R501 B.n651 B.n9 585
R502 B.n752 B.n751 585
R503 B.n751 B.n750 585
R504 B.n11 B.n10 585
R505 B.n749 B.n11 585
R506 B.n747 B.n746 585
R507 B.n748 B.n747 585
R508 B.n745 B.n16 585
R509 B.n16 B.n15 585
R510 B.n744 B.n743 585
R511 B.n743 B.n742 585
R512 B.n18 B.n17 585
R513 B.n741 B.n18 585
R514 B.n739 B.n738 585
R515 B.n740 B.n739 585
R516 B.n737 B.n23 585
R517 B.n23 B.n22 585
R518 B.n736 B.n735 585
R519 B.n735 B.n734 585
R520 B.n25 B.n24 585
R521 B.n733 B.n25 585
R522 B.n731 B.n730 585
R523 B.n732 B.n731 585
R524 B.n729 B.n30 585
R525 B.n30 B.n29 585
R526 B.n728 B.n727 585
R527 B.n727 B.n726 585
R528 B.n32 B.n31 585
R529 B.n725 B.n32 585
R530 B.n723 B.n722 585
R531 B.n724 B.n723 585
R532 B.n721 B.n37 585
R533 B.n37 B.n36 585
R534 B.n720 B.n719 585
R535 B.n719 B.n718 585
R536 B.n39 B.n38 585
R537 B.n717 B.n39 585
R538 B.n715 B.n714 585
R539 B.n716 B.n715 585
R540 B.n713 B.n44 585
R541 B.n44 B.n43 585
R542 B.n712 B.n711 585
R543 B.n711 B.n710 585
R544 B.n46 B.n45 585
R545 B.n709 B.n46 585
R546 B.n707 B.n706 585
R547 B.n708 B.n707 585
R548 B.n705 B.n50 585
R549 B.n53 B.n50 585
R550 B.n704 B.n703 585
R551 B.n703 B.n702 585
R552 B.n52 B.n51 585
R553 B.n701 B.n52 585
R554 B.n699 B.n698 585
R555 B.n700 B.n699 585
R556 B.n697 B.n58 585
R557 B.n58 B.n57 585
R558 B.n696 B.n695 585
R559 B.n695 B.n694 585
R560 B.n760 B.n759 585
R561 B.n758 B.n2 585
R562 B.n695 B.n60 487.695
R563 B.n691 B.n61 487.695
R564 B.n549 B.n335 487.695
R565 B.n551 B.n333 487.695
R566 B.n106 B.t14 440.452
R567 B.n104 B.t10 440.452
R568 B.n355 B.t17 440.452
R569 B.n361 B.t21 440.452
R570 B.n693 B.n692 256.663
R571 B.n693 B.n102 256.663
R572 B.n693 B.n101 256.663
R573 B.n693 B.n100 256.663
R574 B.n693 B.n99 256.663
R575 B.n693 B.n98 256.663
R576 B.n693 B.n97 256.663
R577 B.n693 B.n96 256.663
R578 B.n693 B.n95 256.663
R579 B.n693 B.n94 256.663
R580 B.n693 B.n93 256.663
R581 B.n693 B.n92 256.663
R582 B.n693 B.n91 256.663
R583 B.n693 B.n90 256.663
R584 B.n693 B.n89 256.663
R585 B.n693 B.n88 256.663
R586 B.n693 B.n87 256.663
R587 B.n693 B.n86 256.663
R588 B.n693 B.n85 256.663
R589 B.n693 B.n84 256.663
R590 B.n693 B.n83 256.663
R591 B.n693 B.n82 256.663
R592 B.n693 B.n81 256.663
R593 B.n693 B.n80 256.663
R594 B.n693 B.n79 256.663
R595 B.n693 B.n78 256.663
R596 B.n693 B.n77 256.663
R597 B.n693 B.n76 256.663
R598 B.n693 B.n75 256.663
R599 B.n693 B.n74 256.663
R600 B.n693 B.n73 256.663
R601 B.n693 B.n72 256.663
R602 B.n693 B.n71 256.663
R603 B.n693 B.n70 256.663
R604 B.n693 B.n69 256.663
R605 B.n693 B.n68 256.663
R606 B.n693 B.n67 256.663
R607 B.n693 B.n66 256.663
R608 B.n693 B.n65 256.663
R609 B.n693 B.n64 256.663
R610 B.n693 B.n63 256.663
R611 B.n693 B.n62 256.663
R612 B.n382 B.n334 256.663
R613 B.n388 B.n334 256.663
R614 B.n390 B.n334 256.663
R615 B.n396 B.n334 256.663
R616 B.n398 B.n334 256.663
R617 B.n404 B.n334 256.663
R618 B.n406 B.n334 256.663
R619 B.n412 B.n334 256.663
R620 B.n414 B.n334 256.663
R621 B.n420 B.n334 256.663
R622 B.n422 B.n334 256.663
R623 B.n428 B.n334 256.663
R624 B.n430 B.n334 256.663
R625 B.n436 B.n334 256.663
R626 B.n438 B.n334 256.663
R627 B.n444 B.n334 256.663
R628 B.n446 B.n334 256.663
R629 B.n452 B.n334 256.663
R630 B.n454 B.n334 256.663
R631 B.n460 B.n334 256.663
R632 B.n462 B.n334 256.663
R633 B.n468 B.n334 256.663
R634 B.n470 B.n334 256.663
R635 B.n477 B.n334 256.663
R636 B.n479 B.n334 256.663
R637 B.n485 B.n334 256.663
R638 B.n487 B.n334 256.663
R639 B.n493 B.n334 256.663
R640 B.n495 B.n334 256.663
R641 B.n501 B.n334 256.663
R642 B.n503 B.n334 256.663
R643 B.n509 B.n334 256.663
R644 B.n511 B.n334 256.663
R645 B.n517 B.n334 256.663
R646 B.n519 B.n334 256.663
R647 B.n525 B.n334 256.663
R648 B.n527 B.n334 256.663
R649 B.n533 B.n334 256.663
R650 B.n535 B.n334 256.663
R651 B.n541 B.n334 256.663
R652 B.n544 B.n334 256.663
R653 B.n762 B.n761 256.663
R654 B.n110 B.n109 163.367
R655 B.n114 B.n113 163.367
R656 B.n118 B.n117 163.367
R657 B.n122 B.n121 163.367
R658 B.n126 B.n125 163.367
R659 B.n130 B.n129 163.367
R660 B.n134 B.n133 163.367
R661 B.n138 B.n137 163.367
R662 B.n142 B.n141 163.367
R663 B.n146 B.n145 163.367
R664 B.n150 B.n149 163.367
R665 B.n154 B.n153 163.367
R666 B.n158 B.n157 163.367
R667 B.n162 B.n161 163.367
R668 B.n166 B.n165 163.367
R669 B.n170 B.n169 163.367
R670 B.n174 B.n173 163.367
R671 B.n178 B.n177 163.367
R672 B.n183 B.n182 163.367
R673 B.n187 B.n186 163.367
R674 B.n191 B.n190 163.367
R675 B.n195 B.n194 163.367
R676 B.n199 B.n198 163.367
R677 B.n204 B.n203 163.367
R678 B.n208 B.n207 163.367
R679 B.n212 B.n211 163.367
R680 B.n216 B.n215 163.367
R681 B.n220 B.n219 163.367
R682 B.n224 B.n223 163.367
R683 B.n228 B.n227 163.367
R684 B.n232 B.n231 163.367
R685 B.n236 B.n235 163.367
R686 B.n240 B.n239 163.367
R687 B.n244 B.n243 163.367
R688 B.n248 B.n247 163.367
R689 B.n252 B.n251 163.367
R690 B.n256 B.n255 163.367
R691 B.n260 B.n259 163.367
R692 B.n264 B.n263 163.367
R693 B.n268 B.n267 163.367
R694 B.n270 B.n103 163.367
R695 B.n549 B.n329 163.367
R696 B.n557 B.n329 163.367
R697 B.n557 B.n327 163.367
R698 B.n561 B.n327 163.367
R699 B.n561 B.n322 163.367
R700 B.n570 B.n322 163.367
R701 B.n570 B.n320 163.367
R702 B.n574 B.n320 163.367
R703 B.n574 B.n314 163.367
R704 B.n582 B.n314 163.367
R705 B.n582 B.n312 163.367
R706 B.n586 B.n312 163.367
R707 B.n586 B.n306 163.367
R708 B.n594 B.n306 163.367
R709 B.n594 B.n304 163.367
R710 B.n598 B.n304 163.367
R711 B.n598 B.n298 163.367
R712 B.n606 B.n298 163.367
R713 B.n606 B.n296 163.367
R714 B.n610 B.n296 163.367
R715 B.n610 B.n290 163.367
R716 B.n618 B.n290 163.367
R717 B.n618 B.n288 163.367
R718 B.n622 B.n288 163.367
R719 B.n622 B.n282 163.367
R720 B.n630 B.n282 163.367
R721 B.n630 B.n280 163.367
R722 B.n635 B.n280 163.367
R723 B.n635 B.n274 163.367
R724 B.n643 B.n274 163.367
R725 B.n644 B.n643 163.367
R726 B.n644 B.n5 163.367
R727 B.n6 B.n5 163.367
R728 B.n7 B.n6 163.367
R729 B.n650 B.n7 163.367
R730 B.n652 B.n650 163.367
R731 B.n652 B.n12 163.367
R732 B.n13 B.n12 163.367
R733 B.n14 B.n13 163.367
R734 B.n657 B.n14 163.367
R735 B.n657 B.n19 163.367
R736 B.n20 B.n19 163.367
R737 B.n21 B.n20 163.367
R738 B.n662 B.n21 163.367
R739 B.n662 B.n26 163.367
R740 B.n27 B.n26 163.367
R741 B.n28 B.n27 163.367
R742 B.n667 B.n28 163.367
R743 B.n667 B.n33 163.367
R744 B.n34 B.n33 163.367
R745 B.n35 B.n34 163.367
R746 B.n672 B.n35 163.367
R747 B.n672 B.n40 163.367
R748 B.n41 B.n40 163.367
R749 B.n42 B.n41 163.367
R750 B.n677 B.n42 163.367
R751 B.n677 B.n47 163.367
R752 B.n48 B.n47 163.367
R753 B.n49 B.n48 163.367
R754 B.n682 B.n49 163.367
R755 B.n682 B.n54 163.367
R756 B.n55 B.n54 163.367
R757 B.n56 B.n55 163.367
R758 B.n687 B.n56 163.367
R759 B.n687 B.n61 163.367
R760 B.n383 B.n381 163.367
R761 B.n387 B.n381 163.367
R762 B.n391 B.n389 163.367
R763 B.n395 B.n379 163.367
R764 B.n399 B.n397 163.367
R765 B.n403 B.n377 163.367
R766 B.n407 B.n405 163.367
R767 B.n411 B.n375 163.367
R768 B.n415 B.n413 163.367
R769 B.n419 B.n373 163.367
R770 B.n423 B.n421 163.367
R771 B.n427 B.n371 163.367
R772 B.n431 B.n429 163.367
R773 B.n435 B.n369 163.367
R774 B.n439 B.n437 163.367
R775 B.n443 B.n367 163.367
R776 B.n447 B.n445 163.367
R777 B.n451 B.n365 163.367
R778 B.n455 B.n453 163.367
R779 B.n459 B.n360 163.367
R780 B.n463 B.n461 163.367
R781 B.n467 B.n358 163.367
R782 B.n471 B.n469 163.367
R783 B.n476 B.n354 163.367
R784 B.n480 B.n478 163.367
R785 B.n484 B.n352 163.367
R786 B.n488 B.n486 163.367
R787 B.n492 B.n350 163.367
R788 B.n496 B.n494 163.367
R789 B.n500 B.n348 163.367
R790 B.n504 B.n502 163.367
R791 B.n508 B.n346 163.367
R792 B.n512 B.n510 163.367
R793 B.n516 B.n344 163.367
R794 B.n520 B.n518 163.367
R795 B.n524 B.n342 163.367
R796 B.n528 B.n526 163.367
R797 B.n532 B.n340 163.367
R798 B.n536 B.n534 163.367
R799 B.n540 B.n338 163.367
R800 B.n543 B.n542 163.367
R801 B.n545 B.n335 163.367
R802 B.n551 B.n331 163.367
R803 B.n555 B.n331 163.367
R804 B.n555 B.n325 163.367
R805 B.n564 B.n325 163.367
R806 B.n564 B.n323 163.367
R807 B.n568 B.n323 163.367
R808 B.n568 B.n318 163.367
R809 B.n576 B.n318 163.367
R810 B.n576 B.n316 163.367
R811 B.n580 B.n316 163.367
R812 B.n580 B.n310 163.367
R813 B.n588 B.n310 163.367
R814 B.n588 B.n308 163.367
R815 B.n592 B.n308 163.367
R816 B.n592 B.n302 163.367
R817 B.n600 B.n302 163.367
R818 B.n600 B.n300 163.367
R819 B.n604 B.n300 163.367
R820 B.n604 B.n294 163.367
R821 B.n612 B.n294 163.367
R822 B.n612 B.n292 163.367
R823 B.n616 B.n292 163.367
R824 B.n616 B.n286 163.367
R825 B.n624 B.n286 163.367
R826 B.n624 B.n284 163.367
R827 B.n628 B.n284 163.367
R828 B.n628 B.n278 163.367
R829 B.n637 B.n278 163.367
R830 B.n637 B.n276 163.367
R831 B.n641 B.n276 163.367
R832 B.n641 B.n3 163.367
R833 B.n760 B.n3 163.367
R834 B.n756 B.n2 163.367
R835 B.n756 B.n755 163.367
R836 B.n755 B.n9 163.367
R837 B.n751 B.n9 163.367
R838 B.n751 B.n11 163.367
R839 B.n747 B.n11 163.367
R840 B.n747 B.n16 163.367
R841 B.n743 B.n16 163.367
R842 B.n743 B.n18 163.367
R843 B.n739 B.n18 163.367
R844 B.n739 B.n23 163.367
R845 B.n735 B.n23 163.367
R846 B.n735 B.n25 163.367
R847 B.n731 B.n25 163.367
R848 B.n731 B.n30 163.367
R849 B.n727 B.n30 163.367
R850 B.n727 B.n32 163.367
R851 B.n723 B.n32 163.367
R852 B.n723 B.n37 163.367
R853 B.n719 B.n37 163.367
R854 B.n719 B.n39 163.367
R855 B.n715 B.n39 163.367
R856 B.n715 B.n44 163.367
R857 B.n711 B.n44 163.367
R858 B.n711 B.n46 163.367
R859 B.n707 B.n46 163.367
R860 B.n707 B.n50 163.367
R861 B.n703 B.n50 163.367
R862 B.n703 B.n52 163.367
R863 B.n699 B.n52 163.367
R864 B.n699 B.n58 163.367
R865 B.n695 B.n58 163.367
R866 B.n104 B.t12 99.454
R867 B.n355 B.t20 99.454
R868 B.n106 B.t15 99.4412
R869 B.n361 B.t23 99.4412
R870 B.n550 B.n334 93.1555
R871 B.n694 B.n693 93.1555
R872 B.n105 B.t13 72.4964
R873 B.n356 B.t19 72.4964
R874 B.n107 B.t16 72.4837
R875 B.n362 B.t22 72.4837
R876 B.n62 B.n60 71.676
R877 B.n110 B.n63 71.676
R878 B.n114 B.n64 71.676
R879 B.n118 B.n65 71.676
R880 B.n122 B.n66 71.676
R881 B.n126 B.n67 71.676
R882 B.n130 B.n68 71.676
R883 B.n134 B.n69 71.676
R884 B.n138 B.n70 71.676
R885 B.n142 B.n71 71.676
R886 B.n146 B.n72 71.676
R887 B.n150 B.n73 71.676
R888 B.n154 B.n74 71.676
R889 B.n158 B.n75 71.676
R890 B.n162 B.n76 71.676
R891 B.n166 B.n77 71.676
R892 B.n170 B.n78 71.676
R893 B.n174 B.n79 71.676
R894 B.n178 B.n80 71.676
R895 B.n183 B.n81 71.676
R896 B.n187 B.n82 71.676
R897 B.n191 B.n83 71.676
R898 B.n195 B.n84 71.676
R899 B.n199 B.n85 71.676
R900 B.n204 B.n86 71.676
R901 B.n208 B.n87 71.676
R902 B.n212 B.n88 71.676
R903 B.n216 B.n89 71.676
R904 B.n220 B.n90 71.676
R905 B.n224 B.n91 71.676
R906 B.n228 B.n92 71.676
R907 B.n232 B.n93 71.676
R908 B.n236 B.n94 71.676
R909 B.n240 B.n95 71.676
R910 B.n244 B.n96 71.676
R911 B.n248 B.n97 71.676
R912 B.n252 B.n98 71.676
R913 B.n256 B.n99 71.676
R914 B.n260 B.n100 71.676
R915 B.n264 B.n101 71.676
R916 B.n268 B.n102 71.676
R917 B.n692 B.n103 71.676
R918 B.n692 B.n691 71.676
R919 B.n270 B.n102 71.676
R920 B.n267 B.n101 71.676
R921 B.n263 B.n100 71.676
R922 B.n259 B.n99 71.676
R923 B.n255 B.n98 71.676
R924 B.n251 B.n97 71.676
R925 B.n247 B.n96 71.676
R926 B.n243 B.n95 71.676
R927 B.n239 B.n94 71.676
R928 B.n235 B.n93 71.676
R929 B.n231 B.n92 71.676
R930 B.n227 B.n91 71.676
R931 B.n223 B.n90 71.676
R932 B.n219 B.n89 71.676
R933 B.n215 B.n88 71.676
R934 B.n211 B.n87 71.676
R935 B.n207 B.n86 71.676
R936 B.n203 B.n85 71.676
R937 B.n198 B.n84 71.676
R938 B.n194 B.n83 71.676
R939 B.n190 B.n82 71.676
R940 B.n186 B.n81 71.676
R941 B.n182 B.n80 71.676
R942 B.n177 B.n79 71.676
R943 B.n173 B.n78 71.676
R944 B.n169 B.n77 71.676
R945 B.n165 B.n76 71.676
R946 B.n161 B.n75 71.676
R947 B.n157 B.n74 71.676
R948 B.n153 B.n73 71.676
R949 B.n149 B.n72 71.676
R950 B.n145 B.n71 71.676
R951 B.n141 B.n70 71.676
R952 B.n137 B.n69 71.676
R953 B.n133 B.n68 71.676
R954 B.n129 B.n67 71.676
R955 B.n125 B.n66 71.676
R956 B.n121 B.n65 71.676
R957 B.n117 B.n64 71.676
R958 B.n113 B.n63 71.676
R959 B.n109 B.n62 71.676
R960 B.n382 B.n333 71.676
R961 B.n388 B.n387 71.676
R962 B.n391 B.n390 71.676
R963 B.n396 B.n395 71.676
R964 B.n399 B.n398 71.676
R965 B.n404 B.n403 71.676
R966 B.n407 B.n406 71.676
R967 B.n412 B.n411 71.676
R968 B.n415 B.n414 71.676
R969 B.n420 B.n419 71.676
R970 B.n423 B.n422 71.676
R971 B.n428 B.n427 71.676
R972 B.n431 B.n430 71.676
R973 B.n436 B.n435 71.676
R974 B.n439 B.n438 71.676
R975 B.n444 B.n443 71.676
R976 B.n447 B.n446 71.676
R977 B.n452 B.n451 71.676
R978 B.n455 B.n454 71.676
R979 B.n460 B.n459 71.676
R980 B.n463 B.n462 71.676
R981 B.n468 B.n467 71.676
R982 B.n471 B.n470 71.676
R983 B.n477 B.n476 71.676
R984 B.n480 B.n479 71.676
R985 B.n485 B.n484 71.676
R986 B.n488 B.n487 71.676
R987 B.n493 B.n492 71.676
R988 B.n496 B.n495 71.676
R989 B.n501 B.n500 71.676
R990 B.n504 B.n503 71.676
R991 B.n509 B.n508 71.676
R992 B.n512 B.n511 71.676
R993 B.n517 B.n516 71.676
R994 B.n520 B.n519 71.676
R995 B.n525 B.n524 71.676
R996 B.n528 B.n527 71.676
R997 B.n533 B.n532 71.676
R998 B.n536 B.n535 71.676
R999 B.n541 B.n540 71.676
R1000 B.n544 B.n543 71.676
R1001 B.n383 B.n382 71.676
R1002 B.n389 B.n388 71.676
R1003 B.n390 B.n379 71.676
R1004 B.n397 B.n396 71.676
R1005 B.n398 B.n377 71.676
R1006 B.n405 B.n404 71.676
R1007 B.n406 B.n375 71.676
R1008 B.n413 B.n412 71.676
R1009 B.n414 B.n373 71.676
R1010 B.n421 B.n420 71.676
R1011 B.n422 B.n371 71.676
R1012 B.n429 B.n428 71.676
R1013 B.n430 B.n369 71.676
R1014 B.n437 B.n436 71.676
R1015 B.n438 B.n367 71.676
R1016 B.n445 B.n444 71.676
R1017 B.n446 B.n365 71.676
R1018 B.n453 B.n452 71.676
R1019 B.n454 B.n360 71.676
R1020 B.n461 B.n460 71.676
R1021 B.n462 B.n358 71.676
R1022 B.n469 B.n468 71.676
R1023 B.n470 B.n354 71.676
R1024 B.n478 B.n477 71.676
R1025 B.n479 B.n352 71.676
R1026 B.n486 B.n485 71.676
R1027 B.n487 B.n350 71.676
R1028 B.n494 B.n493 71.676
R1029 B.n495 B.n348 71.676
R1030 B.n502 B.n501 71.676
R1031 B.n503 B.n346 71.676
R1032 B.n510 B.n509 71.676
R1033 B.n511 B.n344 71.676
R1034 B.n518 B.n517 71.676
R1035 B.n519 B.n342 71.676
R1036 B.n526 B.n525 71.676
R1037 B.n527 B.n340 71.676
R1038 B.n534 B.n533 71.676
R1039 B.n535 B.n338 71.676
R1040 B.n542 B.n541 71.676
R1041 B.n545 B.n544 71.676
R1042 B.n761 B.n760 71.676
R1043 B.n761 B.n2 71.676
R1044 B.n180 B.n107 59.5399
R1045 B.n201 B.n105 59.5399
R1046 B.n474 B.n356 59.5399
R1047 B.n363 B.n362 59.5399
R1048 B.n550 B.n330 47.6286
R1049 B.n556 B.n330 47.6286
R1050 B.n556 B.n326 47.6286
R1051 B.n563 B.n326 47.6286
R1052 B.n563 B.n562 47.6286
R1053 B.n569 B.n319 47.6286
R1054 B.n575 B.n319 47.6286
R1055 B.n575 B.n315 47.6286
R1056 B.n581 B.n315 47.6286
R1057 B.n581 B.n311 47.6286
R1058 B.n587 B.n311 47.6286
R1059 B.n593 B.n307 47.6286
R1060 B.n593 B.n303 47.6286
R1061 B.n599 B.n303 47.6286
R1062 B.n605 B.n299 47.6286
R1063 B.n605 B.n295 47.6286
R1064 B.n611 B.n295 47.6286
R1065 B.n617 B.n291 47.6286
R1066 B.n617 B.n287 47.6286
R1067 B.n623 B.n287 47.6286
R1068 B.n629 B.n283 47.6286
R1069 B.n629 B.n279 47.6286
R1070 B.n636 B.n279 47.6286
R1071 B.n642 B.n275 47.6286
R1072 B.n642 B.n4 47.6286
R1073 B.n759 B.n4 47.6286
R1074 B.n759 B.n758 47.6286
R1075 B.n758 B.n757 47.6286
R1076 B.n757 B.n8 47.6286
R1077 B.n651 B.n8 47.6286
R1078 B.n750 B.n749 47.6286
R1079 B.n749 B.n748 47.6286
R1080 B.n748 B.n15 47.6286
R1081 B.n742 B.n741 47.6286
R1082 B.n741 B.n740 47.6286
R1083 B.n740 B.n22 47.6286
R1084 B.n734 B.n733 47.6286
R1085 B.n733 B.n732 47.6286
R1086 B.n732 B.n29 47.6286
R1087 B.n726 B.n725 47.6286
R1088 B.n725 B.n724 47.6286
R1089 B.n724 B.n36 47.6286
R1090 B.n718 B.n717 47.6286
R1091 B.n717 B.n716 47.6286
R1092 B.n716 B.n43 47.6286
R1093 B.n710 B.n43 47.6286
R1094 B.n710 B.n709 47.6286
R1095 B.n709 B.n708 47.6286
R1096 B.n702 B.n53 47.6286
R1097 B.n702 B.n701 47.6286
R1098 B.n701 B.n700 47.6286
R1099 B.n700 B.n57 47.6286
R1100 B.n694 B.n57 47.6286
R1101 B.n636 B.t1 40.6245
R1102 B.n750 B.t9 40.6245
R1103 B.n569 B.t18 37.8228
R1104 B.n708 B.t11 37.8228
R1105 B.n623 B.t2 36.422
R1106 B.n742 B.t4 36.422
R1107 B.n611 B.t8 32.2195
R1108 B.n734 B.t5 32.2195
R1109 B.n552 B.n332 31.6883
R1110 B.n548 B.n547 31.6883
R1111 B.n690 B.n689 31.6883
R1112 B.n696 B.n59 31.6883
R1113 B.n599 B.t0 28.0171
R1114 B.n726 B.t7 28.0171
R1115 B.n107 B.n106 26.9581
R1116 B.n105 B.n104 26.9581
R1117 B.n356 B.n355 26.9581
R1118 B.n362 B.n361 26.9581
R1119 B.n587 B.t3 23.8146
R1120 B.t3 B.n307 23.8146
R1121 B.t6 B.n36 23.8146
R1122 B.n718 B.t6 23.8146
R1123 B.t0 B.n299 19.6121
R1124 B.t7 B.n29 19.6121
R1125 B B.n762 18.0485
R1126 B.t8 B.n291 15.4096
R1127 B.t5 B.n22 15.4096
R1128 B.t2 B.n283 11.2071
R1129 B.t4 B.n15 11.2071
R1130 B.n553 B.n552 10.6151
R1131 B.n554 B.n553 10.6151
R1132 B.n554 B.n324 10.6151
R1133 B.n565 B.n324 10.6151
R1134 B.n566 B.n565 10.6151
R1135 B.n567 B.n566 10.6151
R1136 B.n567 B.n317 10.6151
R1137 B.n577 B.n317 10.6151
R1138 B.n578 B.n577 10.6151
R1139 B.n579 B.n578 10.6151
R1140 B.n579 B.n309 10.6151
R1141 B.n589 B.n309 10.6151
R1142 B.n590 B.n589 10.6151
R1143 B.n591 B.n590 10.6151
R1144 B.n591 B.n301 10.6151
R1145 B.n601 B.n301 10.6151
R1146 B.n602 B.n601 10.6151
R1147 B.n603 B.n602 10.6151
R1148 B.n603 B.n293 10.6151
R1149 B.n613 B.n293 10.6151
R1150 B.n614 B.n613 10.6151
R1151 B.n615 B.n614 10.6151
R1152 B.n615 B.n285 10.6151
R1153 B.n625 B.n285 10.6151
R1154 B.n626 B.n625 10.6151
R1155 B.n627 B.n626 10.6151
R1156 B.n627 B.n277 10.6151
R1157 B.n638 B.n277 10.6151
R1158 B.n639 B.n638 10.6151
R1159 B.n640 B.n639 10.6151
R1160 B.n640 B.n0 10.6151
R1161 B.n384 B.n332 10.6151
R1162 B.n385 B.n384 10.6151
R1163 B.n386 B.n385 10.6151
R1164 B.n386 B.n380 10.6151
R1165 B.n392 B.n380 10.6151
R1166 B.n393 B.n392 10.6151
R1167 B.n394 B.n393 10.6151
R1168 B.n394 B.n378 10.6151
R1169 B.n400 B.n378 10.6151
R1170 B.n401 B.n400 10.6151
R1171 B.n402 B.n401 10.6151
R1172 B.n402 B.n376 10.6151
R1173 B.n408 B.n376 10.6151
R1174 B.n409 B.n408 10.6151
R1175 B.n410 B.n409 10.6151
R1176 B.n410 B.n374 10.6151
R1177 B.n416 B.n374 10.6151
R1178 B.n417 B.n416 10.6151
R1179 B.n418 B.n417 10.6151
R1180 B.n418 B.n372 10.6151
R1181 B.n424 B.n372 10.6151
R1182 B.n425 B.n424 10.6151
R1183 B.n426 B.n425 10.6151
R1184 B.n426 B.n370 10.6151
R1185 B.n432 B.n370 10.6151
R1186 B.n433 B.n432 10.6151
R1187 B.n434 B.n433 10.6151
R1188 B.n434 B.n368 10.6151
R1189 B.n440 B.n368 10.6151
R1190 B.n441 B.n440 10.6151
R1191 B.n442 B.n441 10.6151
R1192 B.n442 B.n366 10.6151
R1193 B.n448 B.n366 10.6151
R1194 B.n449 B.n448 10.6151
R1195 B.n450 B.n449 10.6151
R1196 B.n450 B.n364 10.6151
R1197 B.n457 B.n456 10.6151
R1198 B.n458 B.n457 10.6151
R1199 B.n458 B.n359 10.6151
R1200 B.n464 B.n359 10.6151
R1201 B.n465 B.n464 10.6151
R1202 B.n466 B.n465 10.6151
R1203 B.n466 B.n357 10.6151
R1204 B.n472 B.n357 10.6151
R1205 B.n473 B.n472 10.6151
R1206 B.n475 B.n353 10.6151
R1207 B.n481 B.n353 10.6151
R1208 B.n482 B.n481 10.6151
R1209 B.n483 B.n482 10.6151
R1210 B.n483 B.n351 10.6151
R1211 B.n489 B.n351 10.6151
R1212 B.n490 B.n489 10.6151
R1213 B.n491 B.n490 10.6151
R1214 B.n491 B.n349 10.6151
R1215 B.n497 B.n349 10.6151
R1216 B.n498 B.n497 10.6151
R1217 B.n499 B.n498 10.6151
R1218 B.n499 B.n347 10.6151
R1219 B.n505 B.n347 10.6151
R1220 B.n506 B.n505 10.6151
R1221 B.n507 B.n506 10.6151
R1222 B.n507 B.n345 10.6151
R1223 B.n513 B.n345 10.6151
R1224 B.n514 B.n513 10.6151
R1225 B.n515 B.n514 10.6151
R1226 B.n515 B.n343 10.6151
R1227 B.n521 B.n343 10.6151
R1228 B.n522 B.n521 10.6151
R1229 B.n523 B.n522 10.6151
R1230 B.n523 B.n341 10.6151
R1231 B.n529 B.n341 10.6151
R1232 B.n530 B.n529 10.6151
R1233 B.n531 B.n530 10.6151
R1234 B.n531 B.n339 10.6151
R1235 B.n537 B.n339 10.6151
R1236 B.n538 B.n537 10.6151
R1237 B.n539 B.n538 10.6151
R1238 B.n539 B.n337 10.6151
R1239 B.n337 B.n336 10.6151
R1240 B.n546 B.n336 10.6151
R1241 B.n547 B.n546 10.6151
R1242 B.n548 B.n328 10.6151
R1243 B.n558 B.n328 10.6151
R1244 B.n559 B.n558 10.6151
R1245 B.n560 B.n559 10.6151
R1246 B.n560 B.n321 10.6151
R1247 B.n571 B.n321 10.6151
R1248 B.n572 B.n571 10.6151
R1249 B.n573 B.n572 10.6151
R1250 B.n573 B.n313 10.6151
R1251 B.n583 B.n313 10.6151
R1252 B.n584 B.n583 10.6151
R1253 B.n585 B.n584 10.6151
R1254 B.n585 B.n305 10.6151
R1255 B.n595 B.n305 10.6151
R1256 B.n596 B.n595 10.6151
R1257 B.n597 B.n596 10.6151
R1258 B.n597 B.n297 10.6151
R1259 B.n607 B.n297 10.6151
R1260 B.n608 B.n607 10.6151
R1261 B.n609 B.n608 10.6151
R1262 B.n609 B.n289 10.6151
R1263 B.n619 B.n289 10.6151
R1264 B.n620 B.n619 10.6151
R1265 B.n621 B.n620 10.6151
R1266 B.n621 B.n281 10.6151
R1267 B.n631 B.n281 10.6151
R1268 B.n632 B.n631 10.6151
R1269 B.n634 B.n632 10.6151
R1270 B.n634 B.n633 10.6151
R1271 B.n633 B.n273 10.6151
R1272 B.n645 B.n273 10.6151
R1273 B.n646 B.n645 10.6151
R1274 B.n647 B.n646 10.6151
R1275 B.n648 B.n647 10.6151
R1276 B.n649 B.n648 10.6151
R1277 B.n653 B.n649 10.6151
R1278 B.n654 B.n653 10.6151
R1279 B.n655 B.n654 10.6151
R1280 B.n656 B.n655 10.6151
R1281 B.n658 B.n656 10.6151
R1282 B.n659 B.n658 10.6151
R1283 B.n660 B.n659 10.6151
R1284 B.n661 B.n660 10.6151
R1285 B.n663 B.n661 10.6151
R1286 B.n664 B.n663 10.6151
R1287 B.n665 B.n664 10.6151
R1288 B.n666 B.n665 10.6151
R1289 B.n668 B.n666 10.6151
R1290 B.n669 B.n668 10.6151
R1291 B.n670 B.n669 10.6151
R1292 B.n671 B.n670 10.6151
R1293 B.n673 B.n671 10.6151
R1294 B.n674 B.n673 10.6151
R1295 B.n675 B.n674 10.6151
R1296 B.n676 B.n675 10.6151
R1297 B.n678 B.n676 10.6151
R1298 B.n679 B.n678 10.6151
R1299 B.n680 B.n679 10.6151
R1300 B.n681 B.n680 10.6151
R1301 B.n683 B.n681 10.6151
R1302 B.n684 B.n683 10.6151
R1303 B.n685 B.n684 10.6151
R1304 B.n686 B.n685 10.6151
R1305 B.n688 B.n686 10.6151
R1306 B.n689 B.n688 10.6151
R1307 B.n754 B.n1 10.6151
R1308 B.n754 B.n753 10.6151
R1309 B.n753 B.n752 10.6151
R1310 B.n752 B.n10 10.6151
R1311 B.n746 B.n10 10.6151
R1312 B.n746 B.n745 10.6151
R1313 B.n745 B.n744 10.6151
R1314 B.n744 B.n17 10.6151
R1315 B.n738 B.n17 10.6151
R1316 B.n738 B.n737 10.6151
R1317 B.n737 B.n736 10.6151
R1318 B.n736 B.n24 10.6151
R1319 B.n730 B.n24 10.6151
R1320 B.n730 B.n729 10.6151
R1321 B.n729 B.n728 10.6151
R1322 B.n728 B.n31 10.6151
R1323 B.n722 B.n31 10.6151
R1324 B.n722 B.n721 10.6151
R1325 B.n721 B.n720 10.6151
R1326 B.n720 B.n38 10.6151
R1327 B.n714 B.n38 10.6151
R1328 B.n714 B.n713 10.6151
R1329 B.n713 B.n712 10.6151
R1330 B.n712 B.n45 10.6151
R1331 B.n706 B.n45 10.6151
R1332 B.n706 B.n705 10.6151
R1333 B.n705 B.n704 10.6151
R1334 B.n704 B.n51 10.6151
R1335 B.n698 B.n51 10.6151
R1336 B.n698 B.n697 10.6151
R1337 B.n697 B.n696 10.6151
R1338 B.n108 B.n59 10.6151
R1339 B.n111 B.n108 10.6151
R1340 B.n112 B.n111 10.6151
R1341 B.n115 B.n112 10.6151
R1342 B.n116 B.n115 10.6151
R1343 B.n119 B.n116 10.6151
R1344 B.n120 B.n119 10.6151
R1345 B.n123 B.n120 10.6151
R1346 B.n124 B.n123 10.6151
R1347 B.n127 B.n124 10.6151
R1348 B.n128 B.n127 10.6151
R1349 B.n131 B.n128 10.6151
R1350 B.n132 B.n131 10.6151
R1351 B.n135 B.n132 10.6151
R1352 B.n136 B.n135 10.6151
R1353 B.n139 B.n136 10.6151
R1354 B.n140 B.n139 10.6151
R1355 B.n143 B.n140 10.6151
R1356 B.n144 B.n143 10.6151
R1357 B.n147 B.n144 10.6151
R1358 B.n148 B.n147 10.6151
R1359 B.n151 B.n148 10.6151
R1360 B.n152 B.n151 10.6151
R1361 B.n155 B.n152 10.6151
R1362 B.n156 B.n155 10.6151
R1363 B.n159 B.n156 10.6151
R1364 B.n160 B.n159 10.6151
R1365 B.n163 B.n160 10.6151
R1366 B.n164 B.n163 10.6151
R1367 B.n167 B.n164 10.6151
R1368 B.n168 B.n167 10.6151
R1369 B.n171 B.n168 10.6151
R1370 B.n172 B.n171 10.6151
R1371 B.n175 B.n172 10.6151
R1372 B.n176 B.n175 10.6151
R1373 B.n179 B.n176 10.6151
R1374 B.n184 B.n181 10.6151
R1375 B.n185 B.n184 10.6151
R1376 B.n188 B.n185 10.6151
R1377 B.n189 B.n188 10.6151
R1378 B.n192 B.n189 10.6151
R1379 B.n193 B.n192 10.6151
R1380 B.n196 B.n193 10.6151
R1381 B.n197 B.n196 10.6151
R1382 B.n200 B.n197 10.6151
R1383 B.n205 B.n202 10.6151
R1384 B.n206 B.n205 10.6151
R1385 B.n209 B.n206 10.6151
R1386 B.n210 B.n209 10.6151
R1387 B.n213 B.n210 10.6151
R1388 B.n214 B.n213 10.6151
R1389 B.n217 B.n214 10.6151
R1390 B.n218 B.n217 10.6151
R1391 B.n221 B.n218 10.6151
R1392 B.n222 B.n221 10.6151
R1393 B.n225 B.n222 10.6151
R1394 B.n226 B.n225 10.6151
R1395 B.n229 B.n226 10.6151
R1396 B.n230 B.n229 10.6151
R1397 B.n233 B.n230 10.6151
R1398 B.n234 B.n233 10.6151
R1399 B.n237 B.n234 10.6151
R1400 B.n238 B.n237 10.6151
R1401 B.n241 B.n238 10.6151
R1402 B.n242 B.n241 10.6151
R1403 B.n245 B.n242 10.6151
R1404 B.n246 B.n245 10.6151
R1405 B.n249 B.n246 10.6151
R1406 B.n250 B.n249 10.6151
R1407 B.n253 B.n250 10.6151
R1408 B.n254 B.n253 10.6151
R1409 B.n257 B.n254 10.6151
R1410 B.n258 B.n257 10.6151
R1411 B.n261 B.n258 10.6151
R1412 B.n262 B.n261 10.6151
R1413 B.n265 B.n262 10.6151
R1414 B.n266 B.n265 10.6151
R1415 B.n269 B.n266 10.6151
R1416 B.n271 B.n269 10.6151
R1417 B.n272 B.n271 10.6151
R1418 B.n690 B.n272 10.6151
R1419 B.n562 B.t18 9.80629
R1420 B.n53 B.t11 9.80629
R1421 B.n364 B.n363 9.36635
R1422 B.n475 B.n474 9.36635
R1423 B.n180 B.n179 9.36635
R1424 B.n202 B.n201 9.36635
R1425 B.n762 B.n0 8.11757
R1426 B.n762 B.n1 8.11757
R1427 B.t1 B.n275 7.00464
R1428 B.n651 B.t9 7.00464
R1429 B.n456 B.n363 1.24928
R1430 B.n474 B.n473 1.24928
R1431 B.n181 B.n180 1.24928
R1432 B.n201 B.n200 1.24928
R1433 VN.n4 VN.t0 294.608
R1434 VN.n23 VN.t5 294.608
R1435 VN.n17 VN.t1 274.423
R1436 VN.n36 VN.t4 274.423
R1437 VN.n10 VN.t8 237.136
R1438 VN.n5 VN.t6 237.136
R1439 VN.n1 VN.t3 237.136
R1440 VN.n29 VN.t9 237.136
R1441 VN.n24 VN.t7 237.136
R1442 VN.n20 VN.t2 237.136
R1443 VN.n35 VN.n19 161.3
R1444 VN.n34 VN.n33 161.3
R1445 VN.n32 VN.n31 161.3
R1446 VN.n30 VN.n21 161.3
R1447 VN.n29 VN.n28 161.3
R1448 VN.n27 VN.n22 161.3
R1449 VN.n26 VN.n25 161.3
R1450 VN.n16 VN.n0 161.3
R1451 VN.n15 VN.n14 161.3
R1452 VN.n13 VN.n12 161.3
R1453 VN.n11 VN.n2 161.3
R1454 VN.n10 VN.n9 161.3
R1455 VN.n8 VN.n3 161.3
R1456 VN.n7 VN.n6 161.3
R1457 VN.n37 VN.n36 80.6037
R1458 VN.n18 VN.n17 80.6037
R1459 VN.n6 VN.n3 56.5193
R1460 VN.n12 VN.n11 56.5193
R1461 VN.n25 VN.n22 56.5193
R1462 VN.n31 VN.n30 56.5193
R1463 VN VN.n37 43.9044
R1464 VN.n5 VN.n4 38.2823
R1465 VN.n24 VN.n23 38.2823
R1466 VN.n17 VN.n16 36.5157
R1467 VN.n36 VN.n35 36.5157
R1468 VN.n16 VN.n15 32.2376
R1469 VN.n35 VN.n34 32.2376
R1470 VN.n26 VN.n23 29.1642
R1471 VN.n7 VN.n4 29.1642
R1472 VN.n10 VN.n3 24.4675
R1473 VN.n11 VN.n10 24.4675
R1474 VN.n30 VN.n29 24.4675
R1475 VN.n29 VN.n22 24.4675
R1476 VN.n6 VN.n5 19.0848
R1477 VN.n12 VN.n1 19.0848
R1478 VN.n25 VN.n24 19.0848
R1479 VN.n31 VN.n20 19.0848
R1480 VN.n15 VN.n1 5.38324
R1481 VN.n34 VN.n20 5.38324
R1482 VN.n37 VN.n19 0.285035
R1483 VN.n18 VN.n0 0.285035
R1484 VN.n33 VN.n19 0.189894
R1485 VN.n33 VN.n32 0.189894
R1486 VN.n32 VN.n21 0.189894
R1487 VN.n28 VN.n21 0.189894
R1488 VN.n28 VN.n27 0.189894
R1489 VN.n27 VN.n26 0.189894
R1490 VN.n8 VN.n7 0.189894
R1491 VN.n9 VN.n8 0.189894
R1492 VN.n9 VN.n2 0.189894
R1493 VN.n13 VN.n2 0.189894
R1494 VN.n14 VN.n13 0.189894
R1495 VN.n14 VN.n0 0.189894
R1496 VN VN.n18 0.146778
R1497 VDD2.n1 VDD2.t9 67.7127
R1498 VDD2.n4 VDD2.t5 66.5147
R1499 VDD2.n3 VDD2.n2 65.4594
R1500 VDD2 VDD2.n7 65.4567
R1501 VDD2.n6 VDD2.n5 64.6163
R1502 VDD2.n1 VDD2.n0 64.6161
R1503 VDD2.n4 VDD2.n3 38.3985
R1504 VDD2.n7 VDD2.t2 1.89887
R1505 VDD2.n7 VDD2.t4 1.89887
R1506 VDD2.n5 VDD2.t7 1.89887
R1507 VDD2.n5 VDD2.t0 1.89887
R1508 VDD2.n2 VDD2.t6 1.89887
R1509 VDD2.n2 VDD2.t8 1.89887
R1510 VDD2.n0 VDD2.t3 1.89887
R1511 VDD2.n0 VDD2.t1 1.89887
R1512 VDD2.n6 VDD2.n4 1.19878
R1513 VDD2 VDD2.n6 0.358259
R1514 VDD2.n3 VDD2.n1 0.244723
C0 VP VDD1 7.36902f
C1 VP VDD2 0.387133f
C2 VDD1 VDD2 1.19887f
C3 VN VTAIL 7.195741f
C4 VP VTAIL 7.21019f
C5 VTAIL VDD1 10.871599f
C6 VTAIL VDD2 10.910099f
C7 VN VP 5.84154f
C8 VN VDD1 0.149823f
C9 VN VDD2 7.135601f
C10 VDD2 B 5.10667f
C11 VDD1 B 5.060066f
C12 VTAIL B 6.302358f
C13 VN B 10.875731f
C14 VP B 9.151324f
C15 VDD2.t9 B 2.15202f
C16 VDD2.t3 B 0.190489f
C17 VDD2.t1 B 0.190489f
C18 VDD2.n0 B 1.68388f
C19 VDD2.n1 B 0.634469f
C20 VDD2.t6 B 0.190489f
C21 VDD2.t8 B 0.190489f
C22 VDD2.n2 B 1.68838f
C23 VDD2.n3 B 1.84606f
C24 VDD2.t5 B 2.14595f
C25 VDD2.n4 B 2.2164f
C26 VDD2.t7 B 0.190489f
C27 VDD2.t0 B 0.190489f
C28 VDD2.n5 B 1.68388f
C29 VDD2.n6 B 0.303343f
C30 VDD2.t2 B 0.190489f
C31 VDD2.t4 B 0.190489f
C32 VDD2.n7 B 1.68835f
C33 VN.n0 B 0.04792f
C34 VN.t3 B 1.07711f
C35 VN.n1 B 0.403935f
C36 VN.n2 B 0.035912f
C37 VN.t8 B 1.07711f
C38 VN.n3 B 0.046924f
C39 VN.t0 B 1.1675f
C40 VN.n4 B 0.453782f
C41 VN.t6 B 1.07711f
C42 VN.n5 B 0.453138f
C43 VN.n6 B 0.050662f
C44 VN.n7 B 0.180606f
C45 VN.n8 B 0.035912f
C46 VN.n9 B 0.035912f
C47 VN.n10 B 0.437822f
C48 VN.n11 B 0.046924f
C49 VN.n12 B 0.050662f
C50 VN.n13 B 0.035912f
C51 VN.n14 B 0.035912f
C52 VN.n15 B 0.046572f
C53 VN.n16 B 0.026974f
C54 VN.t1 B 1.13543f
C55 VN.n17 B 0.4599f
C56 VN.n18 B 0.033633f
C57 VN.n19 B 0.04792f
C58 VN.t2 B 1.07711f
C59 VN.n20 B 0.403935f
C60 VN.n21 B 0.035912f
C61 VN.t9 B 1.07711f
C62 VN.n22 B 0.046924f
C63 VN.t5 B 1.1675f
C64 VN.n23 B 0.453782f
C65 VN.t7 B 1.07711f
C66 VN.n24 B 0.453138f
C67 VN.n25 B 0.050662f
C68 VN.n26 B 0.180606f
C69 VN.n27 B 0.035912f
C70 VN.n28 B 0.035912f
C71 VN.n29 B 0.437822f
C72 VN.n30 B 0.046924f
C73 VN.n31 B 0.050662f
C74 VN.n32 B 0.035912f
C75 VN.n33 B 0.035912f
C76 VN.n34 B 0.046572f
C77 VN.n35 B 0.026974f
C78 VN.t4 B 1.13543f
C79 VN.n36 B 0.4599f
C80 VN.n37 B 1.61032f
C81 VDD1.t9 B 2.17756f
C82 VDD1.t7 B 0.19275f
C83 VDD1.t3 B 0.19275f
C84 VDD1.n0 B 1.70386f
C85 VDD1.n1 B 0.648327f
C86 VDD1.t2 B 2.17756f
C87 VDD1.t8 B 0.19275f
C88 VDD1.t6 B 0.19275f
C89 VDD1.n2 B 1.70386f
C90 VDD1.n3 B 0.641999f
C91 VDD1.t4 B 0.19275f
C92 VDD1.t1 B 0.19275f
C93 VDD1.n4 B 1.70842f
C94 VDD1.n5 B 1.94739f
C95 VDD1.t5 B 0.19275f
C96 VDD1.t0 B 0.19275f
C97 VDD1.n6 B 1.70386f
C98 VDD1.n7 B 2.25487f
C99 VTAIL.t19 B 0.206329f
C100 VTAIL.t4 B 0.206329f
C101 VTAIL.n0 B 1.75491f
C102 VTAIL.n1 B 0.401435f
C103 VTAIL.t15 B 2.2372f
C104 VTAIL.n2 B 0.501331f
C105 VTAIL.t14 B 0.206329f
C106 VTAIL.t18 B 0.206329f
C107 VTAIL.n3 B 1.75491f
C108 VTAIL.n4 B 0.431336f
C109 VTAIL.t13 B 0.206329f
C110 VTAIL.t11 B 0.206329f
C111 VTAIL.n5 B 1.75491f
C112 VTAIL.n6 B 1.59332f
C113 VTAIL.t3 B 0.206329f
C114 VTAIL.t0 B 0.206329f
C115 VTAIL.n7 B 1.75491f
C116 VTAIL.n8 B 1.59332f
C117 VTAIL.t8 B 0.206329f
C118 VTAIL.t2 B 0.206329f
C119 VTAIL.n9 B 1.75491f
C120 VTAIL.n10 B 0.431331f
C121 VTAIL.t1 B 2.23721f
C122 VTAIL.n11 B 0.501325f
C123 VTAIL.t16 B 0.206329f
C124 VTAIL.t9 B 0.206329f
C125 VTAIL.n12 B 1.75491f
C126 VTAIL.n13 B 0.4209f
C127 VTAIL.t17 B 0.206329f
C128 VTAIL.t10 B 0.206329f
C129 VTAIL.n14 B 1.75491f
C130 VTAIL.n15 B 0.431331f
C131 VTAIL.t12 B 2.2372f
C132 VTAIL.n16 B 1.57709f
C133 VTAIL.t6 B 2.2372f
C134 VTAIL.n17 B 1.57709f
C135 VTAIL.t5 B 0.206329f
C136 VTAIL.t7 B 0.206329f
C137 VTAIL.n18 B 1.75491f
C138 VTAIL.n19 B 0.354149f
C139 VP.n0 B 0.048757f
C140 VP.t5 B 1.09594f
C141 VP.n1 B 0.410996f
C142 VP.n2 B 0.03654f
C143 VP.t3 B 1.09594f
C144 VP.n3 B 0.047745f
C145 VP.n4 B 0.03654f
C146 VP.t1 B 1.09594f
C147 VP.t7 B 1.15528f
C148 VP.n5 B 0.467939f
C149 VP.n6 B 0.048757f
C150 VP.t9 B 1.15528f
C151 VP.t4 B 1.09594f
C152 VP.n7 B 0.410996f
C153 VP.n8 B 0.03654f
C154 VP.t6 B 1.09594f
C155 VP.n9 B 0.047744f
C156 VP.t0 B 1.18791f
C157 VP.n10 B 0.461714f
C158 VP.t2 B 1.09594f
C159 VP.n11 B 0.46106f
C160 VP.n12 B 0.051548f
C161 VP.n13 B 0.183764f
C162 VP.n14 B 0.03654f
C163 VP.n15 B 0.03654f
C164 VP.n16 B 0.445475f
C165 VP.n17 B 0.047745f
C166 VP.n18 B 0.051548f
C167 VP.n19 B 0.03654f
C168 VP.n20 B 0.03654f
C169 VP.n21 B 0.047386f
C170 VP.n22 B 0.027446f
C171 VP.n23 B 0.467939f
C172 VP.n24 B 1.6181f
C173 VP.n25 B 1.64822f
C174 VP.n26 B 0.048757f
C175 VP.n27 B 0.027446f
C176 VP.n28 B 0.047386f
C177 VP.n29 B 0.410996f
C178 VP.n30 B 0.051548f
C179 VP.n31 B 0.03654f
C180 VP.n32 B 0.03654f
C181 VP.n33 B 0.03654f
C182 VP.n34 B 0.445475f
C183 VP.n35 B 0.047744f
C184 VP.n36 B 0.051548f
C185 VP.n37 B 0.03654f
C186 VP.n38 B 0.03654f
C187 VP.n39 B 0.047386f
C188 VP.n40 B 0.027446f
C189 VP.t8 B 1.15528f
C190 VP.n41 B 0.467939f
C191 VP.n42 B 0.034221f
.ends

