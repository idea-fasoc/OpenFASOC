* NGSPICE file created from diff_pair_sample_1358.ext - technology: sky130A

.subckt diff_pair_sample_1358 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VP.t0 VDD1.t2 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=1.70445 ps=10.66 w=10.33 l=3.94
X1 B.t11 B.t9 B.t10 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=0 ps=0 w=10.33 l=3.94
X2 VDD1.t1 VP.t1 VTAIL.t5 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=1.70445 pd=10.66 as=4.0287 ps=21.44 w=10.33 l=3.94
X3 B.t8 B.t6 B.t7 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=0 ps=0 w=10.33 l=3.94
X4 VDD2.t3 VN.t0 VTAIL.t1 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=1.70445 pd=10.66 as=4.0287 ps=21.44 w=10.33 l=3.94
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=1.70445 pd=10.66 as=4.0287 ps=21.44 w=10.33 l=3.94
X6 B.t5 B.t3 B.t4 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=0 ps=0 w=10.33 l=3.94
X7 VTAIL.t2 VN.t2 VDD2.t1 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=1.70445 ps=10.66 w=10.33 l=3.94
X8 VDD1.t0 VP.t2 VTAIL.t4 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=1.70445 pd=10.66 as=4.0287 ps=21.44 w=10.33 l=3.94
X9 VTAIL.t7 VN.t3 VDD2.t0 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=1.70445 ps=10.66 w=10.33 l=3.94
X10 VTAIL.t3 VP.t3 VDD1.t3 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=1.70445 ps=10.66 w=10.33 l=3.94
X11 B.t2 B.t0 B.t1 w_n3532_n3034# sky130_fd_pr__pfet_01v8 ad=4.0287 pd=21.44 as=0 ps=0 w=10.33 l=3.94
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t3 97.0083
R9 VP.n4 VP.t2 95.5786
R10 VP.n6 VP.n5 63.3422
R11 VP.n20 VP.n19 63.3422
R12 VP.n6 VP.t0 63.1865
R13 VP.n19 VP.t1 63.1865
R14 VP.n13 VP.n12 56.5193
R15 VP.n5 VP.n4 51.0231
R16 VP.n7 VP.n3 24.4675
R17 VP.n11 VP.n3 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n13 VP.n1 24.4675
R20 VP.n17 VP.n1 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n7 VP.n6 18.8401
R23 VP.n19 VP.n18 18.8401
R24 VP.n8 VP.n5 0.417535
R25 VP.n20 VP.n0 0.417535
R26 VP VP.n20 0.394291
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VDD1 VDD1.n1 120.85
R35 VDD1 VDD1.n0 76.7206
R36 VDD1.n0 VDD1.t3 3.14716
R37 VDD1.n0 VDD1.t0 3.14716
R38 VDD1.n1 VDD1.t2 3.14716
R39 VDD1.n1 VDD1.t1 3.14716
R40 VTAIL.n5 VTAIL.t3 63.1305
R41 VTAIL.n4 VTAIL.t0 63.1305
R42 VTAIL.n3 VTAIL.t2 63.1305
R43 VTAIL.n6 VTAIL.t4 63.1303
R44 VTAIL.n7 VTAIL.t1 63.1303
R45 VTAIL.n0 VTAIL.t7 63.1303
R46 VTAIL.n1 VTAIL.t5 63.1303
R47 VTAIL.n2 VTAIL.t6 63.1303
R48 VTAIL.n7 VTAIL.n6 24.9531
R49 VTAIL.n3 VTAIL.n2 24.9531
R50 VTAIL.n4 VTAIL.n3 3.68153
R51 VTAIL.n6 VTAIL.n5 3.68153
R52 VTAIL.n2 VTAIL.n1 3.68153
R53 VTAIL VTAIL.n0 1.89921
R54 VTAIL VTAIL.n7 1.78283
R55 VTAIL.n5 VTAIL.n4 0.470328
R56 VTAIL.n1 VTAIL.n0 0.470328
R57 B.n520 B.n519 585
R58 B.n521 B.n70 585
R59 B.n523 B.n522 585
R60 B.n524 B.n69 585
R61 B.n526 B.n525 585
R62 B.n527 B.n68 585
R63 B.n529 B.n528 585
R64 B.n530 B.n67 585
R65 B.n532 B.n531 585
R66 B.n533 B.n66 585
R67 B.n535 B.n534 585
R68 B.n536 B.n65 585
R69 B.n538 B.n537 585
R70 B.n539 B.n64 585
R71 B.n541 B.n540 585
R72 B.n542 B.n63 585
R73 B.n544 B.n543 585
R74 B.n545 B.n62 585
R75 B.n547 B.n546 585
R76 B.n548 B.n61 585
R77 B.n550 B.n549 585
R78 B.n551 B.n60 585
R79 B.n553 B.n552 585
R80 B.n554 B.n59 585
R81 B.n556 B.n555 585
R82 B.n557 B.n58 585
R83 B.n559 B.n558 585
R84 B.n560 B.n57 585
R85 B.n562 B.n561 585
R86 B.n563 B.n56 585
R87 B.n565 B.n564 585
R88 B.n566 B.n55 585
R89 B.n568 B.n567 585
R90 B.n569 B.n54 585
R91 B.n571 B.n570 585
R92 B.n572 B.n53 585
R93 B.n574 B.n573 585
R94 B.n576 B.n575 585
R95 B.n577 B.n49 585
R96 B.n579 B.n578 585
R97 B.n580 B.n48 585
R98 B.n582 B.n581 585
R99 B.n583 B.n47 585
R100 B.n585 B.n584 585
R101 B.n586 B.n46 585
R102 B.n588 B.n587 585
R103 B.n590 B.n43 585
R104 B.n592 B.n591 585
R105 B.n593 B.n42 585
R106 B.n595 B.n594 585
R107 B.n596 B.n41 585
R108 B.n598 B.n597 585
R109 B.n599 B.n40 585
R110 B.n601 B.n600 585
R111 B.n602 B.n39 585
R112 B.n604 B.n603 585
R113 B.n605 B.n38 585
R114 B.n607 B.n606 585
R115 B.n608 B.n37 585
R116 B.n610 B.n609 585
R117 B.n611 B.n36 585
R118 B.n613 B.n612 585
R119 B.n614 B.n35 585
R120 B.n616 B.n615 585
R121 B.n617 B.n34 585
R122 B.n619 B.n618 585
R123 B.n620 B.n33 585
R124 B.n622 B.n621 585
R125 B.n623 B.n32 585
R126 B.n625 B.n624 585
R127 B.n626 B.n31 585
R128 B.n628 B.n627 585
R129 B.n629 B.n30 585
R130 B.n631 B.n630 585
R131 B.n632 B.n29 585
R132 B.n634 B.n633 585
R133 B.n635 B.n28 585
R134 B.n637 B.n636 585
R135 B.n638 B.n27 585
R136 B.n640 B.n639 585
R137 B.n641 B.n26 585
R138 B.n643 B.n642 585
R139 B.n644 B.n25 585
R140 B.n518 B.n71 585
R141 B.n517 B.n516 585
R142 B.n515 B.n72 585
R143 B.n514 B.n513 585
R144 B.n512 B.n73 585
R145 B.n511 B.n510 585
R146 B.n509 B.n74 585
R147 B.n508 B.n507 585
R148 B.n506 B.n75 585
R149 B.n505 B.n504 585
R150 B.n503 B.n76 585
R151 B.n502 B.n501 585
R152 B.n500 B.n77 585
R153 B.n499 B.n498 585
R154 B.n497 B.n78 585
R155 B.n496 B.n495 585
R156 B.n494 B.n79 585
R157 B.n493 B.n492 585
R158 B.n491 B.n80 585
R159 B.n490 B.n489 585
R160 B.n488 B.n81 585
R161 B.n487 B.n486 585
R162 B.n485 B.n82 585
R163 B.n484 B.n483 585
R164 B.n482 B.n83 585
R165 B.n481 B.n480 585
R166 B.n479 B.n84 585
R167 B.n478 B.n477 585
R168 B.n476 B.n85 585
R169 B.n475 B.n474 585
R170 B.n473 B.n86 585
R171 B.n472 B.n471 585
R172 B.n470 B.n87 585
R173 B.n469 B.n468 585
R174 B.n467 B.n88 585
R175 B.n466 B.n465 585
R176 B.n464 B.n89 585
R177 B.n463 B.n462 585
R178 B.n461 B.n90 585
R179 B.n460 B.n459 585
R180 B.n458 B.n91 585
R181 B.n457 B.n456 585
R182 B.n455 B.n92 585
R183 B.n454 B.n453 585
R184 B.n452 B.n93 585
R185 B.n451 B.n450 585
R186 B.n449 B.n94 585
R187 B.n448 B.n447 585
R188 B.n446 B.n95 585
R189 B.n445 B.n444 585
R190 B.n443 B.n96 585
R191 B.n442 B.n441 585
R192 B.n440 B.n97 585
R193 B.n439 B.n438 585
R194 B.n437 B.n98 585
R195 B.n436 B.n435 585
R196 B.n434 B.n99 585
R197 B.n433 B.n432 585
R198 B.n431 B.n100 585
R199 B.n430 B.n429 585
R200 B.n428 B.n101 585
R201 B.n427 B.n426 585
R202 B.n425 B.n102 585
R203 B.n424 B.n423 585
R204 B.n422 B.n103 585
R205 B.n421 B.n420 585
R206 B.n419 B.n104 585
R207 B.n418 B.n417 585
R208 B.n416 B.n105 585
R209 B.n415 B.n414 585
R210 B.n413 B.n106 585
R211 B.n412 B.n411 585
R212 B.n410 B.n107 585
R213 B.n409 B.n408 585
R214 B.n407 B.n108 585
R215 B.n406 B.n405 585
R216 B.n404 B.n109 585
R217 B.n403 B.n402 585
R218 B.n401 B.n110 585
R219 B.n400 B.n399 585
R220 B.n398 B.n111 585
R221 B.n397 B.n396 585
R222 B.n395 B.n112 585
R223 B.n394 B.n393 585
R224 B.n392 B.n113 585
R225 B.n391 B.n390 585
R226 B.n389 B.n114 585
R227 B.n388 B.n387 585
R228 B.n386 B.n115 585
R229 B.n385 B.n384 585
R230 B.n383 B.n116 585
R231 B.n382 B.n381 585
R232 B.n380 B.n117 585
R233 B.n254 B.n163 585
R234 B.n256 B.n255 585
R235 B.n257 B.n162 585
R236 B.n259 B.n258 585
R237 B.n260 B.n161 585
R238 B.n262 B.n261 585
R239 B.n263 B.n160 585
R240 B.n265 B.n264 585
R241 B.n266 B.n159 585
R242 B.n268 B.n267 585
R243 B.n269 B.n158 585
R244 B.n271 B.n270 585
R245 B.n272 B.n157 585
R246 B.n274 B.n273 585
R247 B.n275 B.n156 585
R248 B.n277 B.n276 585
R249 B.n278 B.n155 585
R250 B.n280 B.n279 585
R251 B.n281 B.n154 585
R252 B.n283 B.n282 585
R253 B.n284 B.n153 585
R254 B.n286 B.n285 585
R255 B.n287 B.n152 585
R256 B.n289 B.n288 585
R257 B.n290 B.n151 585
R258 B.n292 B.n291 585
R259 B.n293 B.n150 585
R260 B.n295 B.n294 585
R261 B.n296 B.n149 585
R262 B.n298 B.n297 585
R263 B.n299 B.n148 585
R264 B.n301 B.n300 585
R265 B.n302 B.n147 585
R266 B.n304 B.n303 585
R267 B.n305 B.n146 585
R268 B.n307 B.n306 585
R269 B.n308 B.n143 585
R270 B.n311 B.n310 585
R271 B.n312 B.n142 585
R272 B.n314 B.n313 585
R273 B.n315 B.n141 585
R274 B.n317 B.n316 585
R275 B.n318 B.n140 585
R276 B.n320 B.n319 585
R277 B.n321 B.n139 585
R278 B.n323 B.n322 585
R279 B.n325 B.n324 585
R280 B.n326 B.n135 585
R281 B.n328 B.n327 585
R282 B.n329 B.n134 585
R283 B.n331 B.n330 585
R284 B.n332 B.n133 585
R285 B.n334 B.n333 585
R286 B.n335 B.n132 585
R287 B.n337 B.n336 585
R288 B.n338 B.n131 585
R289 B.n340 B.n339 585
R290 B.n341 B.n130 585
R291 B.n343 B.n342 585
R292 B.n344 B.n129 585
R293 B.n346 B.n345 585
R294 B.n347 B.n128 585
R295 B.n349 B.n348 585
R296 B.n350 B.n127 585
R297 B.n352 B.n351 585
R298 B.n353 B.n126 585
R299 B.n355 B.n354 585
R300 B.n356 B.n125 585
R301 B.n358 B.n357 585
R302 B.n359 B.n124 585
R303 B.n361 B.n360 585
R304 B.n362 B.n123 585
R305 B.n364 B.n363 585
R306 B.n365 B.n122 585
R307 B.n367 B.n366 585
R308 B.n368 B.n121 585
R309 B.n370 B.n369 585
R310 B.n371 B.n120 585
R311 B.n373 B.n372 585
R312 B.n374 B.n119 585
R313 B.n376 B.n375 585
R314 B.n377 B.n118 585
R315 B.n379 B.n378 585
R316 B.n253 B.n252 585
R317 B.n251 B.n164 585
R318 B.n250 B.n249 585
R319 B.n248 B.n165 585
R320 B.n247 B.n246 585
R321 B.n245 B.n166 585
R322 B.n244 B.n243 585
R323 B.n242 B.n167 585
R324 B.n241 B.n240 585
R325 B.n239 B.n168 585
R326 B.n238 B.n237 585
R327 B.n236 B.n169 585
R328 B.n235 B.n234 585
R329 B.n233 B.n170 585
R330 B.n232 B.n231 585
R331 B.n230 B.n171 585
R332 B.n229 B.n228 585
R333 B.n227 B.n172 585
R334 B.n226 B.n225 585
R335 B.n224 B.n173 585
R336 B.n223 B.n222 585
R337 B.n221 B.n174 585
R338 B.n220 B.n219 585
R339 B.n218 B.n175 585
R340 B.n217 B.n216 585
R341 B.n215 B.n176 585
R342 B.n214 B.n213 585
R343 B.n212 B.n177 585
R344 B.n211 B.n210 585
R345 B.n209 B.n178 585
R346 B.n208 B.n207 585
R347 B.n206 B.n179 585
R348 B.n205 B.n204 585
R349 B.n203 B.n180 585
R350 B.n202 B.n201 585
R351 B.n200 B.n181 585
R352 B.n199 B.n198 585
R353 B.n197 B.n182 585
R354 B.n196 B.n195 585
R355 B.n194 B.n183 585
R356 B.n193 B.n192 585
R357 B.n191 B.n184 585
R358 B.n190 B.n189 585
R359 B.n188 B.n185 585
R360 B.n187 B.n186 585
R361 B.n2 B.n0 585
R362 B.n713 B.n1 585
R363 B.n712 B.n711 585
R364 B.n710 B.n3 585
R365 B.n709 B.n708 585
R366 B.n707 B.n4 585
R367 B.n706 B.n705 585
R368 B.n704 B.n5 585
R369 B.n703 B.n702 585
R370 B.n701 B.n6 585
R371 B.n700 B.n699 585
R372 B.n698 B.n7 585
R373 B.n697 B.n696 585
R374 B.n695 B.n8 585
R375 B.n694 B.n693 585
R376 B.n692 B.n9 585
R377 B.n691 B.n690 585
R378 B.n689 B.n10 585
R379 B.n688 B.n687 585
R380 B.n686 B.n11 585
R381 B.n685 B.n684 585
R382 B.n683 B.n12 585
R383 B.n682 B.n681 585
R384 B.n680 B.n13 585
R385 B.n679 B.n678 585
R386 B.n677 B.n14 585
R387 B.n676 B.n675 585
R388 B.n674 B.n15 585
R389 B.n673 B.n672 585
R390 B.n671 B.n16 585
R391 B.n670 B.n669 585
R392 B.n668 B.n17 585
R393 B.n667 B.n666 585
R394 B.n665 B.n18 585
R395 B.n664 B.n663 585
R396 B.n662 B.n19 585
R397 B.n661 B.n660 585
R398 B.n659 B.n20 585
R399 B.n658 B.n657 585
R400 B.n656 B.n21 585
R401 B.n655 B.n654 585
R402 B.n653 B.n22 585
R403 B.n652 B.n651 585
R404 B.n650 B.n23 585
R405 B.n649 B.n648 585
R406 B.n647 B.n24 585
R407 B.n646 B.n645 585
R408 B.n715 B.n714 585
R409 B.n252 B.n163 463.671
R410 B.n646 B.n25 463.671
R411 B.n378 B.n117 463.671
R412 B.n520 B.n71 463.671
R413 B.n136 B.t0 272.635
R414 B.n144 B.t9 272.635
R415 B.n44 B.t6 272.635
R416 B.n50 B.t3 272.635
R417 B.n136 B.t2 192.897
R418 B.n50 B.t4 192.897
R419 B.n144 B.t11 192.885
R420 B.n44 B.t7 192.885
R421 B.n252 B.n251 163.367
R422 B.n251 B.n250 163.367
R423 B.n250 B.n165 163.367
R424 B.n246 B.n165 163.367
R425 B.n246 B.n245 163.367
R426 B.n245 B.n244 163.367
R427 B.n244 B.n167 163.367
R428 B.n240 B.n167 163.367
R429 B.n240 B.n239 163.367
R430 B.n239 B.n238 163.367
R431 B.n238 B.n169 163.367
R432 B.n234 B.n169 163.367
R433 B.n234 B.n233 163.367
R434 B.n233 B.n232 163.367
R435 B.n232 B.n171 163.367
R436 B.n228 B.n171 163.367
R437 B.n228 B.n227 163.367
R438 B.n227 B.n226 163.367
R439 B.n226 B.n173 163.367
R440 B.n222 B.n173 163.367
R441 B.n222 B.n221 163.367
R442 B.n221 B.n220 163.367
R443 B.n220 B.n175 163.367
R444 B.n216 B.n175 163.367
R445 B.n216 B.n215 163.367
R446 B.n215 B.n214 163.367
R447 B.n214 B.n177 163.367
R448 B.n210 B.n177 163.367
R449 B.n210 B.n209 163.367
R450 B.n209 B.n208 163.367
R451 B.n208 B.n179 163.367
R452 B.n204 B.n179 163.367
R453 B.n204 B.n203 163.367
R454 B.n203 B.n202 163.367
R455 B.n202 B.n181 163.367
R456 B.n198 B.n181 163.367
R457 B.n198 B.n197 163.367
R458 B.n197 B.n196 163.367
R459 B.n196 B.n183 163.367
R460 B.n192 B.n183 163.367
R461 B.n192 B.n191 163.367
R462 B.n191 B.n190 163.367
R463 B.n190 B.n185 163.367
R464 B.n186 B.n185 163.367
R465 B.n186 B.n2 163.367
R466 B.n714 B.n2 163.367
R467 B.n714 B.n713 163.367
R468 B.n713 B.n712 163.367
R469 B.n712 B.n3 163.367
R470 B.n708 B.n3 163.367
R471 B.n708 B.n707 163.367
R472 B.n707 B.n706 163.367
R473 B.n706 B.n5 163.367
R474 B.n702 B.n5 163.367
R475 B.n702 B.n701 163.367
R476 B.n701 B.n700 163.367
R477 B.n700 B.n7 163.367
R478 B.n696 B.n7 163.367
R479 B.n696 B.n695 163.367
R480 B.n695 B.n694 163.367
R481 B.n694 B.n9 163.367
R482 B.n690 B.n9 163.367
R483 B.n690 B.n689 163.367
R484 B.n689 B.n688 163.367
R485 B.n688 B.n11 163.367
R486 B.n684 B.n11 163.367
R487 B.n684 B.n683 163.367
R488 B.n683 B.n682 163.367
R489 B.n682 B.n13 163.367
R490 B.n678 B.n13 163.367
R491 B.n678 B.n677 163.367
R492 B.n677 B.n676 163.367
R493 B.n676 B.n15 163.367
R494 B.n672 B.n15 163.367
R495 B.n672 B.n671 163.367
R496 B.n671 B.n670 163.367
R497 B.n670 B.n17 163.367
R498 B.n666 B.n17 163.367
R499 B.n666 B.n665 163.367
R500 B.n665 B.n664 163.367
R501 B.n664 B.n19 163.367
R502 B.n660 B.n19 163.367
R503 B.n660 B.n659 163.367
R504 B.n659 B.n658 163.367
R505 B.n658 B.n21 163.367
R506 B.n654 B.n21 163.367
R507 B.n654 B.n653 163.367
R508 B.n653 B.n652 163.367
R509 B.n652 B.n23 163.367
R510 B.n648 B.n23 163.367
R511 B.n648 B.n647 163.367
R512 B.n647 B.n646 163.367
R513 B.n256 B.n163 163.367
R514 B.n257 B.n256 163.367
R515 B.n258 B.n257 163.367
R516 B.n258 B.n161 163.367
R517 B.n262 B.n161 163.367
R518 B.n263 B.n262 163.367
R519 B.n264 B.n263 163.367
R520 B.n264 B.n159 163.367
R521 B.n268 B.n159 163.367
R522 B.n269 B.n268 163.367
R523 B.n270 B.n269 163.367
R524 B.n270 B.n157 163.367
R525 B.n274 B.n157 163.367
R526 B.n275 B.n274 163.367
R527 B.n276 B.n275 163.367
R528 B.n276 B.n155 163.367
R529 B.n280 B.n155 163.367
R530 B.n281 B.n280 163.367
R531 B.n282 B.n281 163.367
R532 B.n282 B.n153 163.367
R533 B.n286 B.n153 163.367
R534 B.n287 B.n286 163.367
R535 B.n288 B.n287 163.367
R536 B.n288 B.n151 163.367
R537 B.n292 B.n151 163.367
R538 B.n293 B.n292 163.367
R539 B.n294 B.n293 163.367
R540 B.n294 B.n149 163.367
R541 B.n298 B.n149 163.367
R542 B.n299 B.n298 163.367
R543 B.n300 B.n299 163.367
R544 B.n300 B.n147 163.367
R545 B.n304 B.n147 163.367
R546 B.n305 B.n304 163.367
R547 B.n306 B.n305 163.367
R548 B.n306 B.n143 163.367
R549 B.n311 B.n143 163.367
R550 B.n312 B.n311 163.367
R551 B.n313 B.n312 163.367
R552 B.n313 B.n141 163.367
R553 B.n317 B.n141 163.367
R554 B.n318 B.n317 163.367
R555 B.n319 B.n318 163.367
R556 B.n319 B.n139 163.367
R557 B.n323 B.n139 163.367
R558 B.n324 B.n323 163.367
R559 B.n324 B.n135 163.367
R560 B.n328 B.n135 163.367
R561 B.n329 B.n328 163.367
R562 B.n330 B.n329 163.367
R563 B.n330 B.n133 163.367
R564 B.n334 B.n133 163.367
R565 B.n335 B.n334 163.367
R566 B.n336 B.n335 163.367
R567 B.n336 B.n131 163.367
R568 B.n340 B.n131 163.367
R569 B.n341 B.n340 163.367
R570 B.n342 B.n341 163.367
R571 B.n342 B.n129 163.367
R572 B.n346 B.n129 163.367
R573 B.n347 B.n346 163.367
R574 B.n348 B.n347 163.367
R575 B.n348 B.n127 163.367
R576 B.n352 B.n127 163.367
R577 B.n353 B.n352 163.367
R578 B.n354 B.n353 163.367
R579 B.n354 B.n125 163.367
R580 B.n358 B.n125 163.367
R581 B.n359 B.n358 163.367
R582 B.n360 B.n359 163.367
R583 B.n360 B.n123 163.367
R584 B.n364 B.n123 163.367
R585 B.n365 B.n364 163.367
R586 B.n366 B.n365 163.367
R587 B.n366 B.n121 163.367
R588 B.n370 B.n121 163.367
R589 B.n371 B.n370 163.367
R590 B.n372 B.n371 163.367
R591 B.n372 B.n119 163.367
R592 B.n376 B.n119 163.367
R593 B.n377 B.n376 163.367
R594 B.n378 B.n377 163.367
R595 B.n382 B.n117 163.367
R596 B.n383 B.n382 163.367
R597 B.n384 B.n383 163.367
R598 B.n384 B.n115 163.367
R599 B.n388 B.n115 163.367
R600 B.n389 B.n388 163.367
R601 B.n390 B.n389 163.367
R602 B.n390 B.n113 163.367
R603 B.n394 B.n113 163.367
R604 B.n395 B.n394 163.367
R605 B.n396 B.n395 163.367
R606 B.n396 B.n111 163.367
R607 B.n400 B.n111 163.367
R608 B.n401 B.n400 163.367
R609 B.n402 B.n401 163.367
R610 B.n402 B.n109 163.367
R611 B.n406 B.n109 163.367
R612 B.n407 B.n406 163.367
R613 B.n408 B.n407 163.367
R614 B.n408 B.n107 163.367
R615 B.n412 B.n107 163.367
R616 B.n413 B.n412 163.367
R617 B.n414 B.n413 163.367
R618 B.n414 B.n105 163.367
R619 B.n418 B.n105 163.367
R620 B.n419 B.n418 163.367
R621 B.n420 B.n419 163.367
R622 B.n420 B.n103 163.367
R623 B.n424 B.n103 163.367
R624 B.n425 B.n424 163.367
R625 B.n426 B.n425 163.367
R626 B.n426 B.n101 163.367
R627 B.n430 B.n101 163.367
R628 B.n431 B.n430 163.367
R629 B.n432 B.n431 163.367
R630 B.n432 B.n99 163.367
R631 B.n436 B.n99 163.367
R632 B.n437 B.n436 163.367
R633 B.n438 B.n437 163.367
R634 B.n438 B.n97 163.367
R635 B.n442 B.n97 163.367
R636 B.n443 B.n442 163.367
R637 B.n444 B.n443 163.367
R638 B.n444 B.n95 163.367
R639 B.n448 B.n95 163.367
R640 B.n449 B.n448 163.367
R641 B.n450 B.n449 163.367
R642 B.n450 B.n93 163.367
R643 B.n454 B.n93 163.367
R644 B.n455 B.n454 163.367
R645 B.n456 B.n455 163.367
R646 B.n456 B.n91 163.367
R647 B.n460 B.n91 163.367
R648 B.n461 B.n460 163.367
R649 B.n462 B.n461 163.367
R650 B.n462 B.n89 163.367
R651 B.n466 B.n89 163.367
R652 B.n467 B.n466 163.367
R653 B.n468 B.n467 163.367
R654 B.n468 B.n87 163.367
R655 B.n472 B.n87 163.367
R656 B.n473 B.n472 163.367
R657 B.n474 B.n473 163.367
R658 B.n474 B.n85 163.367
R659 B.n478 B.n85 163.367
R660 B.n479 B.n478 163.367
R661 B.n480 B.n479 163.367
R662 B.n480 B.n83 163.367
R663 B.n484 B.n83 163.367
R664 B.n485 B.n484 163.367
R665 B.n486 B.n485 163.367
R666 B.n486 B.n81 163.367
R667 B.n490 B.n81 163.367
R668 B.n491 B.n490 163.367
R669 B.n492 B.n491 163.367
R670 B.n492 B.n79 163.367
R671 B.n496 B.n79 163.367
R672 B.n497 B.n496 163.367
R673 B.n498 B.n497 163.367
R674 B.n498 B.n77 163.367
R675 B.n502 B.n77 163.367
R676 B.n503 B.n502 163.367
R677 B.n504 B.n503 163.367
R678 B.n504 B.n75 163.367
R679 B.n508 B.n75 163.367
R680 B.n509 B.n508 163.367
R681 B.n510 B.n509 163.367
R682 B.n510 B.n73 163.367
R683 B.n514 B.n73 163.367
R684 B.n515 B.n514 163.367
R685 B.n516 B.n515 163.367
R686 B.n516 B.n71 163.367
R687 B.n642 B.n25 163.367
R688 B.n642 B.n641 163.367
R689 B.n641 B.n640 163.367
R690 B.n640 B.n27 163.367
R691 B.n636 B.n27 163.367
R692 B.n636 B.n635 163.367
R693 B.n635 B.n634 163.367
R694 B.n634 B.n29 163.367
R695 B.n630 B.n29 163.367
R696 B.n630 B.n629 163.367
R697 B.n629 B.n628 163.367
R698 B.n628 B.n31 163.367
R699 B.n624 B.n31 163.367
R700 B.n624 B.n623 163.367
R701 B.n623 B.n622 163.367
R702 B.n622 B.n33 163.367
R703 B.n618 B.n33 163.367
R704 B.n618 B.n617 163.367
R705 B.n617 B.n616 163.367
R706 B.n616 B.n35 163.367
R707 B.n612 B.n35 163.367
R708 B.n612 B.n611 163.367
R709 B.n611 B.n610 163.367
R710 B.n610 B.n37 163.367
R711 B.n606 B.n37 163.367
R712 B.n606 B.n605 163.367
R713 B.n605 B.n604 163.367
R714 B.n604 B.n39 163.367
R715 B.n600 B.n39 163.367
R716 B.n600 B.n599 163.367
R717 B.n599 B.n598 163.367
R718 B.n598 B.n41 163.367
R719 B.n594 B.n41 163.367
R720 B.n594 B.n593 163.367
R721 B.n593 B.n592 163.367
R722 B.n592 B.n43 163.367
R723 B.n587 B.n43 163.367
R724 B.n587 B.n586 163.367
R725 B.n586 B.n585 163.367
R726 B.n585 B.n47 163.367
R727 B.n581 B.n47 163.367
R728 B.n581 B.n580 163.367
R729 B.n580 B.n579 163.367
R730 B.n579 B.n49 163.367
R731 B.n575 B.n49 163.367
R732 B.n575 B.n574 163.367
R733 B.n574 B.n53 163.367
R734 B.n570 B.n53 163.367
R735 B.n570 B.n569 163.367
R736 B.n569 B.n568 163.367
R737 B.n568 B.n55 163.367
R738 B.n564 B.n55 163.367
R739 B.n564 B.n563 163.367
R740 B.n563 B.n562 163.367
R741 B.n562 B.n57 163.367
R742 B.n558 B.n57 163.367
R743 B.n558 B.n557 163.367
R744 B.n557 B.n556 163.367
R745 B.n556 B.n59 163.367
R746 B.n552 B.n59 163.367
R747 B.n552 B.n551 163.367
R748 B.n551 B.n550 163.367
R749 B.n550 B.n61 163.367
R750 B.n546 B.n61 163.367
R751 B.n546 B.n545 163.367
R752 B.n545 B.n544 163.367
R753 B.n544 B.n63 163.367
R754 B.n540 B.n63 163.367
R755 B.n540 B.n539 163.367
R756 B.n539 B.n538 163.367
R757 B.n538 B.n65 163.367
R758 B.n534 B.n65 163.367
R759 B.n534 B.n533 163.367
R760 B.n533 B.n532 163.367
R761 B.n532 B.n67 163.367
R762 B.n528 B.n67 163.367
R763 B.n528 B.n527 163.367
R764 B.n527 B.n526 163.367
R765 B.n526 B.n69 163.367
R766 B.n522 B.n69 163.367
R767 B.n522 B.n521 163.367
R768 B.n521 B.n520 163.367
R769 B.n137 B.t1 110.085
R770 B.n51 B.t5 110.085
R771 B.n145 B.t10 110.073
R772 B.n45 B.t8 110.073
R773 B.n137 B.n136 82.8126
R774 B.n145 B.n144 82.8126
R775 B.n45 B.n44 82.8126
R776 B.n51 B.n50 82.8126
R777 B.n138 B.n137 59.5399
R778 B.n309 B.n145 59.5399
R779 B.n589 B.n45 59.5399
R780 B.n52 B.n51 59.5399
R781 B.n645 B.n644 30.1273
R782 B.n380 B.n379 30.1273
R783 B.n254 B.n253 30.1273
R784 B.n519 B.n518 30.1273
R785 B B.n715 18.0485
R786 B.n644 B.n643 10.6151
R787 B.n643 B.n26 10.6151
R788 B.n639 B.n26 10.6151
R789 B.n639 B.n638 10.6151
R790 B.n638 B.n637 10.6151
R791 B.n637 B.n28 10.6151
R792 B.n633 B.n28 10.6151
R793 B.n633 B.n632 10.6151
R794 B.n632 B.n631 10.6151
R795 B.n631 B.n30 10.6151
R796 B.n627 B.n30 10.6151
R797 B.n627 B.n626 10.6151
R798 B.n626 B.n625 10.6151
R799 B.n625 B.n32 10.6151
R800 B.n621 B.n32 10.6151
R801 B.n621 B.n620 10.6151
R802 B.n620 B.n619 10.6151
R803 B.n619 B.n34 10.6151
R804 B.n615 B.n34 10.6151
R805 B.n615 B.n614 10.6151
R806 B.n614 B.n613 10.6151
R807 B.n613 B.n36 10.6151
R808 B.n609 B.n36 10.6151
R809 B.n609 B.n608 10.6151
R810 B.n608 B.n607 10.6151
R811 B.n607 B.n38 10.6151
R812 B.n603 B.n38 10.6151
R813 B.n603 B.n602 10.6151
R814 B.n602 B.n601 10.6151
R815 B.n601 B.n40 10.6151
R816 B.n597 B.n40 10.6151
R817 B.n597 B.n596 10.6151
R818 B.n596 B.n595 10.6151
R819 B.n595 B.n42 10.6151
R820 B.n591 B.n42 10.6151
R821 B.n591 B.n590 10.6151
R822 B.n588 B.n46 10.6151
R823 B.n584 B.n46 10.6151
R824 B.n584 B.n583 10.6151
R825 B.n583 B.n582 10.6151
R826 B.n582 B.n48 10.6151
R827 B.n578 B.n48 10.6151
R828 B.n578 B.n577 10.6151
R829 B.n577 B.n576 10.6151
R830 B.n573 B.n572 10.6151
R831 B.n572 B.n571 10.6151
R832 B.n571 B.n54 10.6151
R833 B.n567 B.n54 10.6151
R834 B.n567 B.n566 10.6151
R835 B.n566 B.n565 10.6151
R836 B.n565 B.n56 10.6151
R837 B.n561 B.n56 10.6151
R838 B.n561 B.n560 10.6151
R839 B.n560 B.n559 10.6151
R840 B.n559 B.n58 10.6151
R841 B.n555 B.n58 10.6151
R842 B.n555 B.n554 10.6151
R843 B.n554 B.n553 10.6151
R844 B.n553 B.n60 10.6151
R845 B.n549 B.n60 10.6151
R846 B.n549 B.n548 10.6151
R847 B.n548 B.n547 10.6151
R848 B.n547 B.n62 10.6151
R849 B.n543 B.n62 10.6151
R850 B.n543 B.n542 10.6151
R851 B.n542 B.n541 10.6151
R852 B.n541 B.n64 10.6151
R853 B.n537 B.n64 10.6151
R854 B.n537 B.n536 10.6151
R855 B.n536 B.n535 10.6151
R856 B.n535 B.n66 10.6151
R857 B.n531 B.n66 10.6151
R858 B.n531 B.n530 10.6151
R859 B.n530 B.n529 10.6151
R860 B.n529 B.n68 10.6151
R861 B.n525 B.n68 10.6151
R862 B.n525 B.n524 10.6151
R863 B.n524 B.n523 10.6151
R864 B.n523 B.n70 10.6151
R865 B.n519 B.n70 10.6151
R866 B.n381 B.n380 10.6151
R867 B.n381 B.n116 10.6151
R868 B.n385 B.n116 10.6151
R869 B.n386 B.n385 10.6151
R870 B.n387 B.n386 10.6151
R871 B.n387 B.n114 10.6151
R872 B.n391 B.n114 10.6151
R873 B.n392 B.n391 10.6151
R874 B.n393 B.n392 10.6151
R875 B.n393 B.n112 10.6151
R876 B.n397 B.n112 10.6151
R877 B.n398 B.n397 10.6151
R878 B.n399 B.n398 10.6151
R879 B.n399 B.n110 10.6151
R880 B.n403 B.n110 10.6151
R881 B.n404 B.n403 10.6151
R882 B.n405 B.n404 10.6151
R883 B.n405 B.n108 10.6151
R884 B.n409 B.n108 10.6151
R885 B.n410 B.n409 10.6151
R886 B.n411 B.n410 10.6151
R887 B.n411 B.n106 10.6151
R888 B.n415 B.n106 10.6151
R889 B.n416 B.n415 10.6151
R890 B.n417 B.n416 10.6151
R891 B.n417 B.n104 10.6151
R892 B.n421 B.n104 10.6151
R893 B.n422 B.n421 10.6151
R894 B.n423 B.n422 10.6151
R895 B.n423 B.n102 10.6151
R896 B.n427 B.n102 10.6151
R897 B.n428 B.n427 10.6151
R898 B.n429 B.n428 10.6151
R899 B.n429 B.n100 10.6151
R900 B.n433 B.n100 10.6151
R901 B.n434 B.n433 10.6151
R902 B.n435 B.n434 10.6151
R903 B.n435 B.n98 10.6151
R904 B.n439 B.n98 10.6151
R905 B.n440 B.n439 10.6151
R906 B.n441 B.n440 10.6151
R907 B.n441 B.n96 10.6151
R908 B.n445 B.n96 10.6151
R909 B.n446 B.n445 10.6151
R910 B.n447 B.n446 10.6151
R911 B.n447 B.n94 10.6151
R912 B.n451 B.n94 10.6151
R913 B.n452 B.n451 10.6151
R914 B.n453 B.n452 10.6151
R915 B.n453 B.n92 10.6151
R916 B.n457 B.n92 10.6151
R917 B.n458 B.n457 10.6151
R918 B.n459 B.n458 10.6151
R919 B.n459 B.n90 10.6151
R920 B.n463 B.n90 10.6151
R921 B.n464 B.n463 10.6151
R922 B.n465 B.n464 10.6151
R923 B.n465 B.n88 10.6151
R924 B.n469 B.n88 10.6151
R925 B.n470 B.n469 10.6151
R926 B.n471 B.n470 10.6151
R927 B.n471 B.n86 10.6151
R928 B.n475 B.n86 10.6151
R929 B.n476 B.n475 10.6151
R930 B.n477 B.n476 10.6151
R931 B.n477 B.n84 10.6151
R932 B.n481 B.n84 10.6151
R933 B.n482 B.n481 10.6151
R934 B.n483 B.n482 10.6151
R935 B.n483 B.n82 10.6151
R936 B.n487 B.n82 10.6151
R937 B.n488 B.n487 10.6151
R938 B.n489 B.n488 10.6151
R939 B.n489 B.n80 10.6151
R940 B.n493 B.n80 10.6151
R941 B.n494 B.n493 10.6151
R942 B.n495 B.n494 10.6151
R943 B.n495 B.n78 10.6151
R944 B.n499 B.n78 10.6151
R945 B.n500 B.n499 10.6151
R946 B.n501 B.n500 10.6151
R947 B.n501 B.n76 10.6151
R948 B.n505 B.n76 10.6151
R949 B.n506 B.n505 10.6151
R950 B.n507 B.n506 10.6151
R951 B.n507 B.n74 10.6151
R952 B.n511 B.n74 10.6151
R953 B.n512 B.n511 10.6151
R954 B.n513 B.n512 10.6151
R955 B.n513 B.n72 10.6151
R956 B.n517 B.n72 10.6151
R957 B.n518 B.n517 10.6151
R958 B.n255 B.n254 10.6151
R959 B.n255 B.n162 10.6151
R960 B.n259 B.n162 10.6151
R961 B.n260 B.n259 10.6151
R962 B.n261 B.n260 10.6151
R963 B.n261 B.n160 10.6151
R964 B.n265 B.n160 10.6151
R965 B.n266 B.n265 10.6151
R966 B.n267 B.n266 10.6151
R967 B.n267 B.n158 10.6151
R968 B.n271 B.n158 10.6151
R969 B.n272 B.n271 10.6151
R970 B.n273 B.n272 10.6151
R971 B.n273 B.n156 10.6151
R972 B.n277 B.n156 10.6151
R973 B.n278 B.n277 10.6151
R974 B.n279 B.n278 10.6151
R975 B.n279 B.n154 10.6151
R976 B.n283 B.n154 10.6151
R977 B.n284 B.n283 10.6151
R978 B.n285 B.n284 10.6151
R979 B.n285 B.n152 10.6151
R980 B.n289 B.n152 10.6151
R981 B.n290 B.n289 10.6151
R982 B.n291 B.n290 10.6151
R983 B.n291 B.n150 10.6151
R984 B.n295 B.n150 10.6151
R985 B.n296 B.n295 10.6151
R986 B.n297 B.n296 10.6151
R987 B.n297 B.n148 10.6151
R988 B.n301 B.n148 10.6151
R989 B.n302 B.n301 10.6151
R990 B.n303 B.n302 10.6151
R991 B.n303 B.n146 10.6151
R992 B.n307 B.n146 10.6151
R993 B.n308 B.n307 10.6151
R994 B.n310 B.n142 10.6151
R995 B.n314 B.n142 10.6151
R996 B.n315 B.n314 10.6151
R997 B.n316 B.n315 10.6151
R998 B.n316 B.n140 10.6151
R999 B.n320 B.n140 10.6151
R1000 B.n321 B.n320 10.6151
R1001 B.n322 B.n321 10.6151
R1002 B.n326 B.n325 10.6151
R1003 B.n327 B.n326 10.6151
R1004 B.n327 B.n134 10.6151
R1005 B.n331 B.n134 10.6151
R1006 B.n332 B.n331 10.6151
R1007 B.n333 B.n332 10.6151
R1008 B.n333 B.n132 10.6151
R1009 B.n337 B.n132 10.6151
R1010 B.n338 B.n337 10.6151
R1011 B.n339 B.n338 10.6151
R1012 B.n339 B.n130 10.6151
R1013 B.n343 B.n130 10.6151
R1014 B.n344 B.n343 10.6151
R1015 B.n345 B.n344 10.6151
R1016 B.n345 B.n128 10.6151
R1017 B.n349 B.n128 10.6151
R1018 B.n350 B.n349 10.6151
R1019 B.n351 B.n350 10.6151
R1020 B.n351 B.n126 10.6151
R1021 B.n355 B.n126 10.6151
R1022 B.n356 B.n355 10.6151
R1023 B.n357 B.n356 10.6151
R1024 B.n357 B.n124 10.6151
R1025 B.n361 B.n124 10.6151
R1026 B.n362 B.n361 10.6151
R1027 B.n363 B.n362 10.6151
R1028 B.n363 B.n122 10.6151
R1029 B.n367 B.n122 10.6151
R1030 B.n368 B.n367 10.6151
R1031 B.n369 B.n368 10.6151
R1032 B.n369 B.n120 10.6151
R1033 B.n373 B.n120 10.6151
R1034 B.n374 B.n373 10.6151
R1035 B.n375 B.n374 10.6151
R1036 B.n375 B.n118 10.6151
R1037 B.n379 B.n118 10.6151
R1038 B.n253 B.n164 10.6151
R1039 B.n249 B.n164 10.6151
R1040 B.n249 B.n248 10.6151
R1041 B.n248 B.n247 10.6151
R1042 B.n247 B.n166 10.6151
R1043 B.n243 B.n166 10.6151
R1044 B.n243 B.n242 10.6151
R1045 B.n242 B.n241 10.6151
R1046 B.n241 B.n168 10.6151
R1047 B.n237 B.n168 10.6151
R1048 B.n237 B.n236 10.6151
R1049 B.n236 B.n235 10.6151
R1050 B.n235 B.n170 10.6151
R1051 B.n231 B.n170 10.6151
R1052 B.n231 B.n230 10.6151
R1053 B.n230 B.n229 10.6151
R1054 B.n229 B.n172 10.6151
R1055 B.n225 B.n172 10.6151
R1056 B.n225 B.n224 10.6151
R1057 B.n224 B.n223 10.6151
R1058 B.n223 B.n174 10.6151
R1059 B.n219 B.n174 10.6151
R1060 B.n219 B.n218 10.6151
R1061 B.n218 B.n217 10.6151
R1062 B.n217 B.n176 10.6151
R1063 B.n213 B.n176 10.6151
R1064 B.n213 B.n212 10.6151
R1065 B.n212 B.n211 10.6151
R1066 B.n211 B.n178 10.6151
R1067 B.n207 B.n178 10.6151
R1068 B.n207 B.n206 10.6151
R1069 B.n206 B.n205 10.6151
R1070 B.n205 B.n180 10.6151
R1071 B.n201 B.n180 10.6151
R1072 B.n201 B.n200 10.6151
R1073 B.n200 B.n199 10.6151
R1074 B.n199 B.n182 10.6151
R1075 B.n195 B.n182 10.6151
R1076 B.n195 B.n194 10.6151
R1077 B.n194 B.n193 10.6151
R1078 B.n193 B.n184 10.6151
R1079 B.n189 B.n184 10.6151
R1080 B.n189 B.n188 10.6151
R1081 B.n188 B.n187 10.6151
R1082 B.n187 B.n0 10.6151
R1083 B.n711 B.n1 10.6151
R1084 B.n711 B.n710 10.6151
R1085 B.n710 B.n709 10.6151
R1086 B.n709 B.n4 10.6151
R1087 B.n705 B.n4 10.6151
R1088 B.n705 B.n704 10.6151
R1089 B.n704 B.n703 10.6151
R1090 B.n703 B.n6 10.6151
R1091 B.n699 B.n6 10.6151
R1092 B.n699 B.n698 10.6151
R1093 B.n698 B.n697 10.6151
R1094 B.n697 B.n8 10.6151
R1095 B.n693 B.n8 10.6151
R1096 B.n693 B.n692 10.6151
R1097 B.n692 B.n691 10.6151
R1098 B.n691 B.n10 10.6151
R1099 B.n687 B.n10 10.6151
R1100 B.n687 B.n686 10.6151
R1101 B.n686 B.n685 10.6151
R1102 B.n685 B.n12 10.6151
R1103 B.n681 B.n12 10.6151
R1104 B.n681 B.n680 10.6151
R1105 B.n680 B.n679 10.6151
R1106 B.n679 B.n14 10.6151
R1107 B.n675 B.n14 10.6151
R1108 B.n675 B.n674 10.6151
R1109 B.n674 B.n673 10.6151
R1110 B.n673 B.n16 10.6151
R1111 B.n669 B.n16 10.6151
R1112 B.n669 B.n668 10.6151
R1113 B.n668 B.n667 10.6151
R1114 B.n667 B.n18 10.6151
R1115 B.n663 B.n18 10.6151
R1116 B.n663 B.n662 10.6151
R1117 B.n662 B.n661 10.6151
R1118 B.n661 B.n20 10.6151
R1119 B.n657 B.n20 10.6151
R1120 B.n657 B.n656 10.6151
R1121 B.n656 B.n655 10.6151
R1122 B.n655 B.n22 10.6151
R1123 B.n651 B.n22 10.6151
R1124 B.n651 B.n650 10.6151
R1125 B.n650 B.n649 10.6151
R1126 B.n649 B.n24 10.6151
R1127 B.n645 B.n24 10.6151
R1128 B.n589 B.n588 6.5566
R1129 B.n576 B.n52 6.5566
R1130 B.n310 B.n309 6.5566
R1131 B.n322 B.n138 6.5566
R1132 B.n590 B.n589 4.05904
R1133 B.n573 B.n52 4.05904
R1134 B.n309 B.n308 4.05904
R1135 B.n325 B.n138 4.05904
R1136 B.n715 B.n0 2.81026
R1137 B.n715 B.n1 2.81026
R1138 VN.n0 VN.t3 97.0087
R1139 VN.n1 VN.t1 97.0087
R1140 VN.n0 VN.t0 95.5786
R1141 VN.n1 VN.t2 95.5786
R1142 VN VN.n1 51.0612
R1143 VN VN.n0 1.77706
R1144 VDD2.n2 VDD2.n0 120.326
R1145 VDD2.n2 VDD2.n1 76.6625
R1146 VDD2.n1 VDD2.t1 3.14716
R1147 VDD2.n1 VDD2.t2 3.14716
R1148 VDD2.n0 VDD2.t0 3.14716
R1149 VDD2.n0 VDD2.t3 3.14716
R1150 VDD2 VDD2.n2 0.0586897
C0 VDD1 B 1.45442f
C1 VDD2 B 1.52874f
C2 VP w_n3532_n3034# 6.66321f
C3 VTAIL w_n3532_n3034# 3.65539f
C4 VN w_n3532_n3034# 6.20576f
C5 VDD1 w_n3532_n3034# 1.66046f
C6 VP VTAIL 4.60171f
C7 VDD2 w_n3532_n3034# 1.7461f
C8 VP VN 6.85163f
C9 VP VDD1 4.72256f
C10 B w_n3532_n3034# 10.4255f
C11 VN VTAIL 4.5876f
C12 VDD2 VP 0.47973f
C13 VDD1 VTAIL 5.45802f
C14 VDD2 VTAIL 5.52121f
C15 VDD1 VN 0.150369f
C16 VP B 2.10855f
C17 VDD2 VN 4.39428f
C18 VTAIL B 4.89575f
C19 VDD2 VDD1 1.35628f
C20 VN B 1.34321f
C21 VDD2 VSUBS 1.12168f
C22 VDD1 VSUBS 6.338389f
C23 VTAIL VSUBS 1.328008f
C24 VN VSUBS 6.21381f
C25 VP VSUBS 2.956659f
C26 B VSUBS 5.288486f
C27 w_n3532_n3034# VSUBS 0.13228p
C28 VDD2.t0 VSUBS 0.224835f
C29 VDD2.t3 VSUBS 0.224835f
C30 VDD2.n0 VSUBS 2.42261f
C31 VDD2.t1 VSUBS 0.224835f
C32 VDD2.t2 VSUBS 0.224835f
C33 VDD2.n1 VSUBS 1.70852f
C34 VDD2.n2 VSUBS 4.53692f
C35 VN.t3 VSUBS 3.54433f
C36 VN.t0 VSUBS 3.52572f
C37 VN.n0 VSUBS 2.09486f
C38 VN.t1 VSUBS 3.54433f
C39 VN.t2 VSUBS 3.52572f
C40 VN.n1 VSUBS 3.90453f
C41 B.n0 VSUBS 0.004615f
C42 B.n1 VSUBS 0.004615f
C43 B.n2 VSUBS 0.007297f
C44 B.n3 VSUBS 0.007297f
C45 B.n4 VSUBS 0.007297f
C46 B.n5 VSUBS 0.007297f
C47 B.n6 VSUBS 0.007297f
C48 B.n7 VSUBS 0.007297f
C49 B.n8 VSUBS 0.007297f
C50 B.n9 VSUBS 0.007297f
C51 B.n10 VSUBS 0.007297f
C52 B.n11 VSUBS 0.007297f
C53 B.n12 VSUBS 0.007297f
C54 B.n13 VSUBS 0.007297f
C55 B.n14 VSUBS 0.007297f
C56 B.n15 VSUBS 0.007297f
C57 B.n16 VSUBS 0.007297f
C58 B.n17 VSUBS 0.007297f
C59 B.n18 VSUBS 0.007297f
C60 B.n19 VSUBS 0.007297f
C61 B.n20 VSUBS 0.007297f
C62 B.n21 VSUBS 0.007297f
C63 B.n22 VSUBS 0.007297f
C64 B.n23 VSUBS 0.007297f
C65 B.n24 VSUBS 0.007297f
C66 B.n25 VSUBS 0.01649f
C67 B.n26 VSUBS 0.007297f
C68 B.n27 VSUBS 0.007297f
C69 B.n28 VSUBS 0.007297f
C70 B.n29 VSUBS 0.007297f
C71 B.n30 VSUBS 0.007297f
C72 B.n31 VSUBS 0.007297f
C73 B.n32 VSUBS 0.007297f
C74 B.n33 VSUBS 0.007297f
C75 B.n34 VSUBS 0.007297f
C76 B.n35 VSUBS 0.007297f
C77 B.n36 VSUBS 0.007297f
C78 B.n37 VSUBS 0.007297f
C79 B.n38 VSUBS 0.007297f
C80 B.n39 VSUBS 0.007297f
C81 B.n40 VSUBS 0.007297f
C82 B.n41 VSUBS 0.007297f
C83 B.n42 VSUBS 0.007297f
C84 B.n43 VSUBS 0.007297f
C85 B.t8 VSUBS 0.344877f
C86 B.t7 VSUBS 0.374965f
C87 B.t6 VSUBS 1.9976f
C88 B.n44 VSUBS 0.215574f
C89 B.n45 VSUBS 0.080489f
C90 B.n46 VSUBS 0.007297f
C91 B.n47 VSUBS 0.007297f
C92 B.n48 VSUBS 0.007297f
C93 B.n49 VSUBS 0.007297f
C94 B.t5 VSUBS 0.344872f
C95 B.t4 VSUBS 0.37496f
C96 B.t3 VSUBS 1.9976f
C97 B.n50 VSUBS 0.215579f
C98 B.n51 VSUBS 0.080494f
C99 B.n52 VSUBS 0.016907f
C100 B.n53 VSUBS 0.007297f
C101 B.n54 VSUBS 0.007297f
C102 B.n55 VSUBS 0.007297f
C103 B.n56 VSUBS 0.007297f
C104 B.n57 VSUBS 0.007297f
C105 B.n58 VSUBS 0.007297f
C106 B.n59 VSUBS 0.007297f
C107 B.n60 VSUBS 0.007297f
C108 B.n61 VSUBS 0.007297f
C109 B.n62 VSUBS 0.007297f
C110 B.n63 VSUBS 0.007297f
C111 B.n64 VSUBS 0.007297f
C112 B.n65 VSUBS 0.007297f
C113 B.n66 VSUBS 0.007297f
C114 B.n67 VSUBS 0.007297f
C115 B.n68 VSUBS 0.007297f
C116 B.n69 VSUBS 0.007297f
C117 B.n70 VSUBS 0.007297f
C118 B.n71 VSUBS 0.01592f
C119 B.n72 VSUBS 0.007297f
C120 B.n73 VSUBS 0.007297f
C121 B.n74 VSUBS 0.007297f
C122 B.n75 VSUBS 0.007297f
C123 B.n76 VSUBS 0.007297f
C124 B.n77 VSUBS 0.007297f
C125 B.n78 VSUBS 0.007297f
C126 B.n79 VSUBS 0.007297f
C127 B.n80 VSUBS 0.007297f
C128 B.n81 VSUBS 0.007297f
C129 B.n82 VSUBS 0.007297f
C130 B.n83 VSUBS 0.007297f
C131 B.n84 VSUBS 0.007297f
C132 B.n85 VSUBS 0.007297f
C133 B.n86 VSUBS 0.007297f
C134 B.n87 VSUBS 0.007297f
C135 B.n88 VSUBS 0.007297f
C136 B.n89 VSUBS 0.007297f
C137 B.n90 VSUBS 0.007297f
C138 B.n91 VSUBS 0.007297f
C139 B.n92 VSUBS 0.007297f
C140 B.n93 VSUBS 0.007297f
C141 B.n94 VSUBS 0.007297f
C142 B.n95 VSUBS 0.007297f
C143 B.n96 VSUBS 0.007297f
C144 B.n97 VSUBS 0.007297f
C145 B.n98 VSUBS 0.007297f
C146 B.n99 VSUBS 0.007297f
C147 B.n100 VSUBS 0.007297f
C148 B.n101 VSUBS 0.007297f
C149 B.n102 VSUBS 0.007297f
C150 B.n103 VSUBS 0.007297f
C151 B.n104 VSUBS 0.007297f
C152 B.n105 VSUBS 0.007297f
C153 B.n106 VSUBS 0.007297f
C154 B.n107 VSUBS 0.007297f
C155 B.n108 VSUBS 0.007297f
C156 B.n109 VSUBS 0.007297f
C157 B.n110 VSUBS 0.007297f
C158 B.n111 VSUBS 0.007297f
C159 B.n112 VSUBS 0.007297f
C160 B.n113 VSUBS 0.007297f
C161 B.n114 VSUBS 0.007297f
C162 B.n115 VSUBS 0.007297f
C163 B.n116 VSUBS 0.007297f
C164 B.n117 VSUBS 0.01592f
C165 B.n118 VSUBS 0.007297f
C166 B.n119 VSUBS 0.007297f
C167 B.n120 VSUBS 0.007297f
C168 B.n121 VSUBS 0.007297f
C169 B.n122 VSUBS 0.007297f
C170 B.n123 VSUBS 0.007297f
C171 B.n124 VSUBS 0.007297f
C172 B.n125 VSUBS 0.007297f
C173 B.n126 VSUBS 0.007297f
C174 B.n127 VSUBS 0.007297f
C175 B.n128 VSUBS 0.007297f
C176 B.n129 VSUBS 0.007297f
C177 B.n130 VSUBS 0.007297f
C178 B.n131 VSUBS 0.007297f
C179 B.n132 VSUBS 0.007297f
C180 B.n133 VSUBS 0.007297f
C181 B.n134 VSUBS 0.007297f
C182 B.n135 VSUBS 0.007297f
C183 B.t1 VSUBS 0.344872f
C184 B.t2 VSUBS 0.37496f
C185 B.t0 VSUBS 1.9976f
C186 B.n136 VSUBS 0.215579f
C187 B.n137 VSUBS 0.080494f
C188 B.n138 VSUBS 0.016907f
C189 B.n139 VSUBS 0.007297f
C190 B.n140 VSUBS 0.007297f
C191 B.n141 VSUBS 0.007297f
C192 B.n142 VSUBS 0.007297f
C193 B.n143 VSUBS 0.007297f
C194 B.t10 VSUBS 0.344877f
C195 B.t11 VSUBS 0.374965f
C196 B.t9 VSUBS 1.9976f
C197 B.n144 VSUBS 0.215574f
C198 B.n145 VSUBS 0.080489f
C199 B.n146 VSUBS 0.007297f
C200 B.n147 VSUBS 0.007297f
C201 B.n148 VSUBS 0.007297f
C202 B.n149 VSUBS 0.007297f
C203 B.n150 VSUBS 0.007297f
C204 B.n151 VSUBS 0.007297f
C205 B.n152 VSUBS 0.007297f
C206 B.n153 VSUBS 0.007297f
C207 B.n154 VSUBS 0.007297f
C208 B.n155 VSUBS 0.007297f
C209 B.n156 VSUBS 0.007297f
C210 B.n157 VSUBS 0.007297f
C211 B.n158 VSUBS 0.007297f
C212 B.n159 VSUBS 0.007297f
C213 B.n160 VSUBS 0.007297f
C214 B.n161 VSUBS 0.007297f
C215 B.n162 VSUBS 0.007297f
C216 B.n163 VSUBS 0.01649f
C217 B.n164 VSUBS 0.007297f
C218 B.n165 VSUBS 0.007297f
C219 B.n166 VSUBS 0.007297f
C220 B.n167 VSUBS 0.007297f
C221 B.n168 VSUBS 0.007297f
C222 B.n169 VSUBS 0.007297f
C223 B.n170 VSUBS 0.007297f
C224 B.n171 VSUBS 0.007297f
C225 B.n172 VSUBS 0.007297f
C226 B.n173 VSUBS 0.007297f
C227 B.n174 VSUBS 0.007297f
C228 B.n175 VSUBS 0.007297f
C229 B.n176 VSUBS 0.007297f
C230 B.n177 VSUBS 0.007297f
C231 B.n178 VSUBS 0.007297f
C232 B.n179 VSUBS 0.007297f
C233 B.n180 VSUBS 0.007297f
C234 B.n181 VSUBS 0.007297f
C235 B.n182 VSUBS 0.007297f
C236 B.n183 VSUBS 0.007297f
C237 B.n184 VSUBS 0.007297f
C238 B.n185 VSUBS 0.007297f
C239 B.n186 VSUBS 0.007297f
C240 B.n187 VSUBS 0.007297f
C241 B.n188 VSUBS 0.007297f
C242 B.n189 VSUBS 0.007297f
C243 B.n190 VSUBS 0.007297f
C244 B.n191 VSUBS 0.007297f
C245 B.n192 VSUBS 0.007297f
C246 B.n193 VSUBS 0.007297f
C247 B.n194 VSUBS 0.007297f
C248 B.n195 VSUBS 0.007297f
C249 B.n196 VSUBS 0.007297f
C250 B.n197 VSUBS 0.007297f
C251 B.n198 VSUBS 0.007297f
C252 B.n199 VSUBS 0.007297f
C253 B.n200 VSUBS 0.007297f
C254 B.n201 VSUBS 0.007297f
C255 B.n202 VSUBS 0.007297f
C256 B.n203 VSUBS 0.007297f
C257 B.n204 VSUBS 0.007297f
C258 B.n205 VSUBS 0.007297f
C259 B.n206 VSUBS 0.007297f
C260 B.n207 VSUBS 0.007297f
C261 B.n208 VSUBS 0.007297f
C262 B.n209 VSUBS 0.007297f
C263 B.n210 VSUBS 0.007297f
C264 B.n211 VSUBS 0.007297f
C265 B.n212 VSUBS 0.007297f
C266 B.n213 VSUBS 0.007297f
C267 B.n214 VSUBS 0.007297f
C268 B.n215 VSUBS 0.007297f
C269 B.n216 VSUBS 0.007297f
C270 B.n217 VSUBS 0.007297f
C271 B.n218 VSUBS 0.007297f
C272 B.n219 VSUBS 0.007297f
C273 B.n220 VSUBS 0.007297f
C274 B.n221 VSUBS 0.007297f
C275 B.n222 VSUBS 0.007297f
C276 B.n223 VSUBS 0.007297f
C277 B.n224 VSUBS 0.007297f
C278 B.n225 VSUBS 0.007297f
C279 B.n226 VSUBS 0.007297f
C280 B.n227 VSUBS 0.007297f
C281 B.n228 VSUBS 0.007297f
C282 B.n229 VSUBS 0.007297f
C283 B.n230 VSUBS 0.007297f
C284 B.n231 VSUBS 0.007297f
C285 B.n232 VSUBS 0.007297f
C286 B.n233 VSUBS 0.007297f
C287 B.n234 VSUBS 0.007297f
C288 B.n235 VSUBS 0.007297f
C289 B.n236 VSUBS 0.007297f
C290 B.n237 VSUBS 0.007297f
C291 B.n238 VSUBS 0.007297f
C292 B.n239 VSUBS 0.007297f
C293 B.n240 VSUBS 0.007297f
C294 B.n241 VSUBS 0.007297f
C295 B.n242 VSUBS 0.007297f
C296 B.n243 VSUBS 0.007297f
C297 B.n244 VSUBS 0.007297f
C298 B.n245 VSUBS 0.007297f
C299 B.n246 VSUBS 0.007297f
C300 B.n247 VSUBS 0.007297f
C301 B.n248 VSUBS 0.007297f
C302 B.n249 VSUBS 0.007297f
C303 B.n250 VSUBS 0.007297f
C304 B.n251 VSUBS 0.007297f
C305 B.n252 VSUBS 0.01592f
C306 B.n253 VSUBS 0.01592f
C307 B.n254 VSUBS 0.01649f
C308 B.n255 VSUBS 0.007297f
C309 B.n256 VSUBS 0.007297f
C310 B.n257 VSUBS 0.007297f
C311 B.n258 VSUBS 0.007297f
C312 B.n259 VSUBS 0.007297f
C313 B.n260 VSUBS 0.007297f
C314 B.n261 VSUBS 0.007297f
C315 B.n262 VSUBS 0.007297f
C316 B.n263 VSUBS 0.007297f
C317 B.n264 VSUBS 0.007297f
C318 B.n265 VSUBS 0.007297f
C319 B.n266 VSUBS 0.007297f
C320 B.n267 VSUBS 0.007297f
C321 B.n268 VSUBS 0.007297f
C322 B.n269 VSUBS 0.007297f
C323 B.n270 VSUBS 0.007297f
C324 B.n271 VSUBS 0.007297f
C325 B.n272 VSUBS 0.007297f
C326 B.n273 VSUBS 0.007297f
C327 B.n274 VSUBS 0.007297f
C328 B.n275 VSUBS 0.007297f
C329 B.n276 VSUBS 0.007297f
C330 B.n277 VSUBS 0.007297f
C331 B.n278 VSUBS 0.007297f
C332 B.n279 VSUBS 0.007297f
C333 B.n280 VSUBS 0.007297f
C334 B.n281 VSUBS 0.007297f
C335 B.n282 VSUBS 0.007297f
C336 B.n283 VSUBS 0.007297f
C337 B.n284 VSUBS 0.007297f
C338 B.n285 VSUBS 0.007297f
C339 B.n286 VSUBS 0.007297f
C340 B.n287 VSUBS 0.007297f
C341 B.n288 VSUBS 0.007297f
C342 B.n289 VSUBS 0.007297f
C343 B.n290 VSUBS 0.007297f
C344 B.n291 VSUBS 0.007297f
C345 B.n292 VSUBS 0.007297f
C346 B.n293 VSUBS 0.007297f
C347 B.n294 VSUBS 0.007297f
C348 B.n295 VSUBS 0.007297f
C349 B.n296 VSUBS 0.007297f
C350 B.n297 VSUBS 0.007297f
C351 B.n298 VSUBS 0.007297f
C352 B.n299 VSUBS 0.007297f
C353 B.n300 VSUBS 0.007297f
C354 B.n301 VSUBS 0.007297f
C355 B.n302 VSUBS 0.007297f
C356 B.n303 VSUBS 0.007297f
C357 B.n304 VSUBS 0.007297f
C358 B.n305 VSUBS 0.007297f
C359 B.n306 VSUBS 0.007297f
C360 B.n307 VSUBS 0.007297f
C361 B.n308 VSUBS 0.005044f
C362 B.n309 VSUBS 0.016907f
C363 B.n310 VSUBS 0.005902f
C364 B.n311 VSUBS 0.007297f
C365 B.n312 VSUBS 0.007297f
C366 B.n313 VSUBS 0.007297f
C367 B.n314 VSUBS 0.007297f
C368 B.n315 VSUBS 0.007297f
C369 B.n316 VSUBS 0.007297f
C370 B.n317 VSUBS 0.007297f
C371 B.n318 VSUBS 0.007297f
C372 B.n319 VSUBS 0.007297f
C373 B.n320 VSUBS 0.007297f
C374 B.n321 VSUBS 0.007297f
C375 B.n322 VSUBS 0.005902f
C376 B.n323 VSUBS 0.007297f
C377 B.n324 VSUBS 0.007297f
C378 B.n325 VSUBS 0.005044f
C379 B.n326 VSUBS 0.007297f
C380 B.n327 VSUBS 0.007297f
C381 B.n328 VSUBS 0.007297f
C382 B.n329 VSUBS 0.007297f
C383 B.n330 VSUBS 0.007297f
C384 B.n331 VSUBS 0.007297f
C385 B.n332 VSUBS 0.007297f
C386 B.n333 VSUBS 0.007297f
C387 B.n334 VSUBS 0.007297f
C388 B.n335 VSUBS 0.007297f
C389 B.n336 VSUBS 0.007297f
C390 B.n337 VSUBS 0.007297f
C391 B.n338 VSUBS 0.007297f
C392 B.n339 VSUBS 0.007297f
C393 B.n340 VSUBS 0.007297f
C394 B.n341 VSUBS 0.007297f
C395 B.n342 VSUBS 0.007297f
C396 B.n343 VSUBS 0.007297f
C397 B.n344 VSUBS 0.007297f
C398 B.n345 VSUBS 0.007297f
C399 B.n346 VSUBS 0.007297f
C400 B.n347 VSUBS 0.007297f
C401 B.n348 VSUBS 0.007297f
C402 B.n349 VSUBS 0.007297f
C403 B.n350 VSUBS 0.007297f
C404 B.n351 VSUBS 0.007297f
C405 B.n352 VSUBS 0.007297f
C406 B.n353 VSUBS 0.007297f
C407 B.n354 VSUBS 0.007297f
C408 B.n355 VSUBS 0.007297f
C409 B.n356 VSUBS 0.007297f
C410 B.n357 VSUBS 0.007297f
C411 B.n358 VSUBS 0.007297f
C412 B.n359 VSUBS 0.007297f
C413 B.n360 VSUBS 0.007297f
C414 B.n361 VSUBS 0.007297f
C415 B.n362 VSUBS 0.007297f
C416 B.n363 VSUBS 0.007297f
C417 B.n364 VSUBS 0.007297f
C418 B.n365 VSUBS 0.007297f
C419 B.n366 VSUBS 0.007297f
C420 B.n367 VSUBS 0.007297f
C421 B.n368 VSUBS 0.007297f
C422 B.n369 VSUBS 0.007297f
C423 B.n370 VSUBS 0.007297f
C424 B.n371 VSUBS 0.007297f
C425 B.n372 VSUBS 0.007297f
C426 B.n373 VSUBS 0.007297f
C427 B.n374 VSUBS 0.007297f
C428 B.n375 VSUBS 0.007297f
C429 B.n376 VSUBS 0.007297f
C430 B.n377 VSUBS 0.007297f
C431 B.n378 VSUBS 0.01649f
C432 B.n379 VSUBS 0.01649f
C433 B.n380 VSUBS 0.01592f
C434 B.n381 VSUBS 0.007297f
C435 B.n382 VSUBS 0.007297f
C436 B.n383 VSUBS 0.007297f
C437 B.n384 VSUBS 0.007297f
C438 B.n385 VSUBS 0.007297f
C439 B.n386 VSUBS 0.007297f
C440 B.n387 VSUBS 0.007297f
C441 B.n388 VSUBS 0.007297f
C442 B.n389 VSUBS 0.007297f
C443 B.n390 VSUBS 0.007297f
C444 B.n391 VSUBS 0.007297f
C445 B.n392 VSUBS 0.007297f
C446 B.n393 VSUBS 0.007297f
C447 B.n394 VSUBS 0.007297f
C448 B.n395 VSUBS 0.007297f
C449 B.n396 VSUBS 0.007297f
C450 B.n397 VSUBS 0.007297f
C451 B.n398 VSUBS 0.007297f
C452 B.n399 VSUBS 0.007297f
C453 B.n400 VSUBS 0.007297f
C454 B.n401 VSUBS 0.007297f
C455 B.n402 VSUBS 0.007297f
C456 B.n403 VSUBS 0.007297f
C457 B.n404 VSUBS 0.007297f
C458 B.n405 VSUBS 0.007297f
C459 B.n406 VSUBS 0.007297f
C460 B.n407 VSUBS 0.007297f
C461 B.n408 VSUBS 0.007297f
C462 B.n409 VSUBS 0.007297f
C463 B.n410 VSUBS 0.007297f
C464 B.n411 VSUBS 0.007297f
C465 B.n412 VSUBS 0.007297f
C466 B.n413 VSUBS 0.007297f
C467 B.n414 VSUBS 0.007297f
C468 B.n415 VSUBS 0.007297f
C469 B.n416 VSUBS 0.007297f
C470 B.n417 VSUBS 0.007297f
C471 B.n418 VSUBS 0.007297f
C472 B.n419 VSUBS 0.007297f
C473 B.n420 VSUBS 0.007297f
C474 B.n421 VSUBS 0.007297f
C475 B.n422 VSUBS 0.007297f
C476 B.n423 VSUBS 0.007297f
C477 B.n424 VSUBS 0.007297f
C478 B.n425 VSUBS 0.007297f
C479 B.n426 VSUBS 0.007297f
C480 B.n427 VSUBS 0.007297f
C481 B.n428 VSUBS 0.007297f
C482 B.n429 VSUBS 0.007297f
C483 B.n430 VSUBS 0.007297f
C484 B.n431 VSUBS 0.007297f
C485 B.n432 VSUBS 0.007297f
C486 B.n433 VSUBS 0.007297f
C487 B.n434 VSUBS 0.007297f
C488 B.n435 VSUBS 0.007297f
C489 B.n436 VSUBS 0.007297f
C490 B.n437 VSUBS 0.007297f
C491 B.n438 VSUBS 0.007297f
C492 B.n439 VSUBS 0.007297f
C493 B.n440 VSUBS 0.007297f
C494 B.n441 VSUBS 0.007297f
C495 B.n442 VSUBS 0.007297f
C496 B.n443 VSUBS 0.007297f
C497 B.n444 VSUBS 0.007297f
C498 B.n445 VSUBS 0.007297f
C499 B.n446 VSUBS 0.007297f
C500 B.n447 VSUBS 0.007297f
C501 B.n448 VSUBS 0.007297f
C502 B.n449 VSUBS 0.007297f
C503 B.n450 VSUBS 0.007297f
C504 B.n451 VSUBS 0.007297f
C505 B.n452 VSUBS 0.007297f
C506 B.n453 VSUBS 0.007297f
C507 B.n454 VSUBS 0.007297f
C508 B.n455 VSUBS 0.007297f
C509 B.n456 VSUBS 0.007297f
C510 B.n457 VSUBS 0.007297f
C511 B.n458 VSUBS 0.007297f
C512 B.n459 VSUBS 0.007297f
C513 B.n460 VSUBS 0.007297f
C514 B.n461 VSUBS 0.007297f
C515 B.n462 VSUBS 0.007297f
C516 B.n463 VSUBS 0.007297f
C517 B.n464 VSUBS 0.007297f
C518 B.n465 VSUBS 0.007297f
C519 B.n466 VSUBS 0.007297f
C520 B.n467 VSUBS 0.007297f
C521 B.n468 VSUBS 0.007297f
C522 B.n469 VSUBS 0.007297f
C523 B.n470 VSUBS 0.007297f
C524 B.n471 VSUBS 0.007297f
C525 B.n472 VSUBS 0.007297f
C526 B.n473 VSUBS 0.007297f
C527 B.n474 VSUBS 0.007297f
C528 B.n475 VSUBS 0.007297f
C529 B.n476 VSUBS 0.007297f
C530 B.n477 VSUBS 0.007297f
C531 B.n478 VSUBS 0.007297f
C532 B.n479 VSUBS 0.007297f
C533 B.n480 VSUBS 0.007297f
C534 B.n481 VSUBS 0.007297f
C535 B.n482 VSUBS 0.007297f
C536 B.n483 VSUBS 0.007297f
C537 B.n484 VSUBS 0.007297f
C538 B.n485 VSUBS 0.007297f
C539 B.n486 VSUBS 0.007297f
C540 B.n487 VSUBS 0.007297f
C541 B.n488 VSUBS 0.007297f
C542 B.n489 VSUBS 0.007297f
C543 B.n490 VSUBS 0.007297f
C544 B.n491 VSUBS 0.007297f
C545 B.n492 VSUBS 0.007297f
C546 B.n493 VSUBS 0.007297f
C547 B.n494 VSUBS 0.007297f
C548 B.n495 VSUBS 0.007297f
C549 B.n496 VSUBS 0.007297f
C550 B.n497 VSUBS 0.007297f
C551 B.n498 VSUBS 0.007297f
C552 B.n499 VSUBS 0.007297f
C553 B.n500 VSUBS 0.007297f
C554 B.n501 VSUBS 0.007297f
C555 B.n502 VSUBS 0.007297f
C556 B.n503 VSUBS 0.007297f
C557 B.n504 VSUBS 0.007297f
C558 B.n505 VSUBS 0.007297f
C559 B.n506 VSUBS 0.007297f
C560 B.n507 VSUBS 0.007297f
C561 B.n508 VSUBS 0.007297f
C562 B.n509 VSUBS 0.007297f
C563 B.n510 VSUBS 0.007297f
C564 B.n511 VSUBS 0.007297f
C565 B.n512 VSUBS 0.007297f
C566 B.n513 VSUBS 0.007297f
C567 B.n514 VSUBS 0.007297f
C568 B.n515 VSUBS 0.007297f
C569 B.n516 VSUBS 0.007297f
C570 B.n517 VSUBS 0.007297f
C571 B.n518 VSUBS 0.016854f
C572 B.n519 VSUBS 0.015555f
C573 B.n520 VSUBS 0.01649f
C574 B.n521 VSUBS 0.007297f
C575 B.n522 VSUBS 0.007297f
C576 B.n523 VSUBS 0.007297f
C577 B.n524 VSUBS 0.007297f
C578 B.n525 VSUBS 0.007297f
C579 B.n526 VSUBS 0.007297f
C580 B.n527 VSUBS 0.007297f
C581 B.n528 VSUBS 0.007297f
C582 B.n529 VSUBS 0.007297f
C583 B.n530 VSUBS 0.007297f
C584 B.n531 VSUBS 0.007297f
C585 B.n532 VSUBS 0.007297f
C586 B.n533 VSUBS 0.007297f
C587 B.n534 VSUBS 0.007297f
C588 B.n535 VSUBS 0.007297f
C589 B.n536 VSUBS 0.007297f
C590 B.n537 VSUBS 0.007297f
C591 B.n538 VSUBS 0.007297f
C592 B.n539 VSUBS 0.007297f
C593 B.n540 VSUBS 0.007297f
C594 B.n541 VSUBS 0.007297f
C595 B.n542 VSUBS 0.007297f
C596 B.n543 VSUBS 0.007297f
C597 B.n544 VSUBS 0.007297f
C598 B.n545 VSUBS 0.007297f
C599 B.n546 VSUBS 0.007297f
C600 B.n547 VSUBS 0.007297f
C601 B.n548 VSUBS 0.007297f
C602 B.n549 VSUBS 0.007297f
C603 B.n550 VSUBS 0.007297f
C604 B.n551 VSUBS 0.007297f
C605 B.n552 VSUBS 0.007297f
C606 B.n553 VSUBS 0.007297f
C607 B.n554 VSUBS 0.007297f
C608 B.n555 VSUBS 0.007297f
C609 B.n556 VSUBS 0.007297f
C610 B.n557 VSUBS 0.007297f
C611 B.n558 VSUBS 0.007297f
C612 B.n559 VSUBS 0.007297f
C613 B.n560 VSUBS 0.007297f
C614 B.n561 VSUBS 0.007297f
C615 B.n562 VSUBS 0.007297f
C616 B.n563 VSUBS 0.007297f
C617 B.n564 VSUBS 0.007297f
C618 B.n565 VSUBS 0.007297f
C619 B.n566 VSUBS 0.007297f
C620 B.n567 VSUBS 0.007297f
C621 B.n568 VSUBS 0.007297f
C622 B.n569 VSUBS 0.007297f
C623 B.n570 VSUBS 0.007297f
C624 B.n571 VSUBS 0.007297f
C625 B.n572 VSUBS 0.007297f
C626 B.n573 VSUBS 0.005044f
C627 B.n574 VSUBS 0.007297f
C628 B.n575 VSUBS 0.007297f
C629 B.n576 VSUBS 0.005902f
C630 B.n577 VSUBS 0.007297f
C631 B.n578 VSUBS 0.007297f
C632 B.n579 VSUBS 0.007297f
C633 B.n580 VSUBS 0.007297f
C634 B.n581 VSUBS 0.007297f
C635 B.n582 VSUBS 0.007297f
C636 B.n583 VSUBS 0.007297f
C637 B.n584 VSUBS 0.007297f
C638 B.n585 VSUBS 0.007297f
C639 B.n586 VSUBS 0.007297f
C640 B.n587 VSUBS 0.007297f
C641 B.n588 VSUBS 0.005902f
C642 B.n589 VSUBS 0.016907f
C643 B.n590 VSUBS 0.005044f
C644 B.n591 VSUBS 0.007297f
C645 B.n592 VSUBS 0.007297f
C646 B.n593 VSUBS 0.007297f
C647 B.n594 VSUBS 0.007297f
C648 B.n595 VSUBS 0.007297f
C649 B.n596 VSUBS 0.007297f
C650 B.n597 VSUBS 0.007297f
C651 B.n598 VSUBS 0.007297f
C652 B.n599 VSUBS 0.007297f
C653 B.n600 VSUBS 0.007297f
C654 B.n601 VSUBS 0.007297f
C655 B.n602 VSUBS 0.007297f
C656 B.n603 VSUBS 0.007297f
C657 B.n604 VSUBS 0.007297f
C658 B.n605 VSUBS 0.007297f
C659 B.n606 VSUBS 0.007297f
C660 B.n607 VSUBS 0.007297f
C661 B.n608 VSUBS 0.007297f
C662 B.n609 VSUBS 0.007297f
C663 B.n610 VSUBS 0.007297f
C664 B.n611 VSUBS 0.007297f
C665 B.n612 VSUBS 0.007297f
C666 B.n613 VSUBS 0.007297f
C667 B.n614 VSUBS 0.007297f
C668 B.n615 VSUBS 0.007297f
C669 B.n616 VSUBS 0.007297f
C670 B.n617 VSUBS 0.007297f
C671 B.n618 VSUBS 0.007297f
C672 B.n619 VSUBS 0.007297f
C673 B.n620 VSUBS 0.007297f
C674 B.n621 VSUBS 0.007297f
C675 B.n622 VSUBS 0.007297f
C676 B.n623 VSUBS 0.007297f
C677 B.n624 VSUBS 0.007297f
C678 B.n625 VSUBS 0.007297f
C679 B.n626 VSUBS 0.007297f
C680 B.n627 VSUBS 0.007297f
C681 B.n628 VSUBS 0.007297f
C682 B.n629 VSUBS 0.007297f
C683 B.n630 VSUBS 0.007297f
C684 B.n631 VSUBS 0.007297f
C685 B.n632 VSUBS 0.007297f
C686 B.n633 VSUBS 0.007297f
C687 B.n634 VSUBS 0.007297f
C688 B.n635 VSUBS 0.007297f
C689 B.n636 VSUBS 0.007297f
C690 B.n637 VSUBS 0.007297f
C691 B.n638 VSUBS 0.007297f
C692 B.n639 VSUBS 0.007297f
C693 B.n640 VSUBS 0.007297f
C694 B.n641 VSUBS 0.007297f
C695 B.n642 VSUBS 0.007297f
C696 B.n643 VSUBS 0.007297f
C697 B.n644 VSUBS 0.01649f
C698 B.n645 VSUBS 0.01592f
C699 B.n646 VSUBS 0.01592f
C700 B.n647 VSUBS 0.007297f
C701 B.n648 VSUBS 0.007297f
C702 B.n649 VSUBS 0.007297f
C703 B.n650 VSUBS 0.007297f
C704 B.n651 VSUBS 0.007297f
C705 B.n652 VSUBS 0.007297f
C706 B.n653 VSUBS 0.007297f
C707 B.n654 VSUBS 0.007297f
C708 B.n655 VSUBS 0.007297f
C709 B.n656 VSUBS 0.007297f
C710 B.n657 VSUBS 0.007297f
C711 B.n658 VSUBS 0.007297f
C712 B.n659 VSUBS 0.007297f
C713 B.n660 VSUBS 0.007297f
C714 B.n661 VSUBS 0.007297f
C715 B.n662 VSUBS 0.007297f
C716 B.n663 VSUBS 0.007297f
C717 B.n664 VSUBS 0.007297f
C718 B.n665 VSUBS 0.007297f
C719 B.n666 VSUBS 0.007297f
C720 B.n667 VSUBS 0.007297f
C721 B.n668 VSUBS 0.007297f
C722 B.n669 VSUBS 0.007297f
C723 B.n670 VSUBS 0.007297f
C724 B.n671 VSUBS 0.007297f
C725 B.n672 VSUBS 0.007297f
C726 B.n673 VSUBS 0.007297f
C727 B.n674 VSUBS 0.007297f
C728 B.n675 VSUBS 0.007297f
C729 B.n676 VSUBS 0.007297f
C730 B.n677 VSUBS 0.007297f
C731 B.n678 VSUBS 0.007297f
C732 B.n679 VSUBS 0.007297f
C733 B.n680 VSUBS 0.007297f
C734 B.n681 VSUBS 0.007297f
C735 B.n682 VSUBS 0.007297f
C736 B.n683 VSUBS 0.007297f
C737 B.n684 VSUBS 0.007297f
C738 B.n685 VSUBS 0.007297f
C739 B.n686 VSUBS 0.007297f
C740 B.n687 VSUBS 0.007297f
C741 B.n688 VSUBS 0.007297f
C742 B.n689 VSUBS 0.007297f
C743 B.n690 VSUBS 0.007297f
C744 B.n691 VSUBS 0.007297f
C745 B.n692 VSUBS 0.007297f
C746 B.n693 VSUBS 0.007297f
C747 B.n694 VSUBS 0.007297f
C748 B.n695 VSUBS 0.007297f
C749 B.n696 VSUBS 0.007297f
C750 B.n697 VSUBS 0.007297f
C751 B.n698 VSUBS 0.007297f
C752 B.n699 VSUBS 0.007297f
C753 B.n700 VSUBS 0.007297f
C754 B.n701 VSUBS 0.007297f
C755 B.n702 VSUBS 0.007297f
C756 B.n703 VSUBS 0.007297f
C757 B.n704 VSUBS 0.007297f
C758 B.n705 VSUBS 0.007297f
C759 B.n706 VSUBS 0.007297f
C760 B.n707 VSUBS 0.007297f
C761 B.n708 VSUBS 0.007297f
C762 B.n709 VSUBS 0.007297f
C763 B.n710 VSUBS 0.007297f
C764 B.n711 VSUBS 0.007297f
C765 B.n712 VSUBS 0.007297f
C766 B.n713 VSUBS 0.007297f
C767 B.n714 VSUBS 0.007297f
C768 B.n715 VSUBS 0.016524f
C769 VTAIL.t7 VSUBS 1.93654f
C770 VTAIL.n0 VSUBS 0.843909f
C771 VTAIL.t5 VSUBS 1.93654f
C772 VTAIL.n1 VSUBS 0.990739f
C773 VTAIL.t6 VSUBS 1.93654f
C774 VTAIL.n2 VSUBS 2.33619f
C775 VTAIL.t2 VSUBS 1.93654f
C776 VTAIL.n3 VSUBS 2.33619f
C777 VTAIL.t0 VSUBS 1.93654f
C778 VTAIL.n4 VSUBS 0.990733f
C779 VTAIL.t3 VSUBS 1.93654f
C780 VTAIL.n5 VSUBS 0.990733f
C781 VTAIL.t4 VSUBS 1.93653f
C782 VTAIL.n6 VSUBS 2.33619f
C783 VTAIL.t1 VSUBS 1.93654f
C784 VTAIL.n7 VSUBS 2.17977f
C785 VDD1.t3 VSUBS 0.229292f
C786 VDD1.t0 VSUBS 0.229292f
C787 VDD1.n0 VSUBS 1.74304f
C788 VDD1.t2 VSUBS 0.229292f
C789 VDD1.t1 VSUBS 0.229292f
C790 VDD1.n1 VSUBS 2.49644f
C791 VP.n0 VSUBS 0.059564f
C792 VP.t1 VSUBS 3.49534f
C793 VP.n1 VSUBS 0.059018f
C794 VP.n2 VSUBS 0.031666f
C795 VP.n3 VSUBS 0.059018f
C796 VP.t2 VSUBS 3.99547f
C797 VP.t3 VSUBS 4.01656f
C798 VP.n4 VSUBS 4.4166f
C799 VP.n5 VSUBS 1.90847f
C800 VP.t0 VSUBS 3.49534f
C801 VP.n6 VSUBS 1.3681f
C802 VP.n7 VSUBS 0.052315f
C803 VP.n8 VSUBS 0.059564f
C804 VP.n9 VSUBS 0.031666f
C805 VP.n10 VSUBS 0.031666f
C806 VP.n11 VSUBS 0.059018f
C807 VP.n12 VSUBS 0.046227f
C808 VP.n13 VSUBS 0.046227f
C809 VP.n14 VSUBS 0.031666f
C810 VP.n15 VSUBS 0.031666f
C811 VP.n16 VSUBS 0.031666f
C812 VP.n17 VSUBS 0.059018f
C813 VP.n18 VSUBS 0.052315f
C814 VP.n19 VSUBS 1.3681f
C815 VP.n20 VSUBS 0.10279f
.ends

