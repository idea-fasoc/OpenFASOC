* NGSPICE file created from diff_pair_sample_1545.ext - technology: sky130A

.subckt diff_pair_sample_1545 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VN.t0 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X1 VTAIL.t11 VN.t1 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=0.87
X2 VDD2.t0 VN.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X3 VTAIL.t13 VP.t0 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X4 VDD1.t6 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=0.87
X5 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=0.87
X6 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=0.87
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=0.87
X8 VTAIL.t9 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X9 VTAIL.t14 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=0.87
X10 VDD2.t1 VN.t4 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=0.87
X11 VTAIL.t1 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X12 VDD1.t3 VP.t4 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0 ps=0 w=2.74 l=0.87
X14 VDD2.t5 VN.t5 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=0.87
X15 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X16 VTAIL.t5 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=0.87
X17 VDD1.t2 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=1.0686 ps=6.26 w=2.74 l=0.87
X18 VDD1.t1 VP.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4521 pd=3.07 as=0.4521 ps=3.07 w=2.74 l=0.87
X19 VTAIL.t2 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0686 pd=6.26 as=0.4521 ps=3.07 w=2.74 l=0.87
R0 VN.n12 VN.n11 161.3
R1 VN.n25 VN.n24 161.3
R2 VN.n23 VN.n13 161.3
R3 VN.n22 VN.n21 161.3
R4 VN.n20 VN.n19 161.3
R5 VN.n18 VN.n15 161.3
R6 VN.n10 VN.n0 161.3
R7 VN.n9 VN.n8 161.3
R8 VN.n7 VN.n6 161.3
R9 VN.n5 VN.n2 161.3
R10 VN.n3 VN.t7 143.125
R11 VN.n16 VN.t5 143.125
R12 VN.n11 VN.t4 121.055
R13 VN.n24 VN.t1 121.055
R14 VN.n4 VN.t2 75.9016
R15 VN.n1 VN.t3 75.9016
R16 VN.n17 VN.t0 75.9016
R17 VN.n14 VN.t6 75.9016
R18 VN.n6 VN.n5 56.5617
R19 VN.n19 VN.n18 56.5617
R20 VN.n10 VN.n9 45.4209
R21 VN.n23 VN.n22 45.4209
R22 VN.n16 VN.n15 42.7264
R23 VN.n3 VN.n2 42.7264
R24 VN.n4 VN.n3 36.9171
R25 VN.n17 VN.n16 36.9171
R26 VN VN.n25 36.1994
R27 VN.n5 VN.n4 17.2148
R28 VN.n6 VN.n1 17.2148
R29 VN.n18 VN.n17 17.2148
R30 VN.n19 VN.n14 17.2148
R31 VN.n11 VN.n10 16.7975
R32 VN.n24 VN.n23 16.7975
R33 VN.n9 VN.n1 7.37805
R34 VN.n22 VN.n14 7.37805
R35 VN.n25 VN.n13 0.189894
R36 VN.n21 VN.n13 0.189894
R37 VN.n21 VN.n20 0.189894
R38 VN.n20 VN.n15 0.189894
R39 VN.n7 VN.n2 0.189894
R40 VN.n8 VN.n7 0.189894
R41 VN.n8 VN.n0 0.189894
R42 VN.n12 VN.n0 0.189894
R43 VN VN.n12 0.0516364
R44 VDD2.n2 VDD2.n1 80.9024
R45 VDD2.n2 VDD2.n0 80.9024
R46 VDD2 VDD2.n5 80.8996
R47 VDD2.n4 VDD2.n3 80.4407
R48 VDD2.n4 VDD2.n2 30.7325
R49 VDD2.n5 VDD2.t6 7.22678
R50 VDD2.n5 VDD2.t5 7.22678
R51 VDD2.n3 VDD2.t7 7.22678
R52 VDD2.n3 VDD2.t3 7.22678
R53 VDD2.n1 VDD2.t4 7.22678
R54 VDD2.n1 VDD2.t1 7.22678
R55 VDD2.n0 VDD2.t2 7.22678
R56 VDD2.n0 VDD2.t0 7.22678
R57 VDD2 VDD2.n4 0.575931
R58 VTAIL.n11 VTAIL.t14 70.9882
R59 VTAIL.n10 VTAIL.t7 70.9882
R60 VTAIL.n7 VTAIL.t11 70.9882
R61 VTAIL.n15 VTAIL.t8 70.9879
R62 VTAIL.n2 VTAIL.t5 70.9879
R63 VTAIL.n3 VTAIL.t4 70.9879
R64 VTAIL.n6 VTAIL.t2 70.9879
R65 VTAIL.n14 VTAIL.t0 70.9879
R66 VTAIL.n13 VTAIL.n12 63.7619
R67 VTAIL.n9 VTAIL.n8 63.7619
R68 VTAIL.n1 VTAIL.n0 63.7617
R69 VTAIL.n5 VTAIL.n4 63.7617
R70 VTAIL.n15 VTAIL.n14 15.7634
R71 VTAIL.n7 VTAIL.n6 15.7634
R72 VTAIL.n0 VTAIL.t10 7.22678
R73 VTAIL.n0 VTAIL.t9 7.22678
R74 VTAIL.n4 VTAIL.t15 7.22678
R75 VTAIL.n4 VTAIL.t1 7.22678
R76 VTAIL.n12 VTAIL.t3 7.22678
R77 VTAIL.n12 VTAIL.t13 7.22678
R78 VTAIL.n8 VTAIL.t6 7.22678
R79 VTAIL.n8 VTAIL.t12 7.22678
R80 VTAIL.n9 VTAIL.n7 1.03498
R81 VTAIL.n10 VTAIL.n9 1.03498
R82 VTAIL.n13 VTAIL.n11 1.03498
R83 VTAIL.n14 VTAIL.n13 1.03498
R84 VTAIL.n6 VTAIL.n5 1.03498
R85 VTAIL.n5 VTAIL.n3 1.03498
R86 VTAIL.n2 VTAIL.n1 1.03498
R87 VTAIL VTAIL.n15 0.976793
R88 VTAIL.n11 VTAIL.n10 0.470328
R89 VTAIL.n3 VTAIL.n2 0.470328
R90 VTAIL VTAIL.n1 0.0586897
R91 B.n406 B.n405 585
R92 B.n147 B.n68 585
R93 B.n146 B.n145 585
R94 B.n144 B.n143 585
R95 B.n142 B.n141 585
R96 B.n140 B.n139 585
R97 B.n138 B.n137 585
R98 B.n136 B.n135 585
R99 B.n134 B.n133 585
R100 B.n132 B.n131 585
R101 B.n130 B.n129 585
R102 B.n128 B.n127 585
R103 B.n126 B.n125 585
R104 B.n124 B.n123 585
R105 B.n122 B.n121 585
R106 B.n120 B.n119 585
R107 B.n118 B.n117 585
R108 B.n116 B.n115 585
R109 B.n114 B.n113 585
R110 B.n112 B.n111 585
R111 B.n110 B.n109 585
R112 B.n108 B.n107 585
R113 B.n106 B.n105 585
R114 B.n104 B.n103 585
R115 B.n102 B.n101 585
R116 B.n100 B.n99 585
R117 B.n98 B.n97 585
R118 B.n96 B.n95 585
R119 B.n94 B.n93 585
R120 B.n92 B.n91 585
R121 B.n90 B.n89 585
R122 B.n88 B.n87 585
R123 B.n86 B.n85 585
R124 B.n84 B.n83 585
R125 B.n82 B.n81 585
R126 B.n80 B.n79 585
R127 B.n78 B.n77 585
R128 B.n76 B.n75 585
R129 B.n404 B.n49 585
R130 B.n409 B.n49 585
R131 B.n403 B.n48 585
R132 B.n410 B.n48 585
R133 B.n402 B.n401 585
R134 B.n401 B.n44 585
R135 B.n400 B.n43 585
R136 B.n416 B.n43 585
R137 B.n399 B.n42 585
R138 B.n417 B.n42 585
R139 B.n398 B.n41 585
R140 B.n418 B.n41 585
R141 B.n397 B.n396 585
R142 B.n396 B.n37 585
R143 B.n395 B.n36 585
R144 B.n424 B.n36 585
R145 B.n394 B.n35 585
R146 B.n425 B.n35 585
R147 B.n393 B.n34 585
R148 B.n426 B.n34 585
R149 B.n392 B.n391 585
R150 B.n391 B.n30 585
R151 B.n390 B.n29 585
R152 B.n432 B.n29 585
R153 B.n389 B.n28 585
R154 B.n433 B.n28 585
R155 B.n388 B.n27 585
R156 B.n434 B.n27 585
R157 B.n387 B.n386 585
R158 B.n386 B.n23 585
R159 B.n385 B.n22 585
R160 B.n440 B.n22 585
R161 B.n384 B.n21 585
R162 B.n441 B.n21 585
R163 B.n383 B.n20 585
R164 B.n442 B.n20 585
R165 B.n382 B.n381 585
R166 B.n381 B.n19 585
R167 B.n380 B.n15 585
R168 B.n448 B.n15 585
R169 B.n379 B.n14 585
R170 B.n449 B.n14 585
R171 B.n378 B.n13 585
R172 B.n450 B.n13 585
R173 B.n377 B.n376 585
R174 B.n376 B.n12 585
R175 B.n375 B.n374 585
R176 B.n375 B.n8 585
R177 B.n373 B.n7 585
R178 B.n457 B.n7 585
R179 B.n372 B.n6 585
R180 B.n458 B.n6 585
R181 B.n371 B.n5 585
R182 B.n459 B.n5 585
R183 B.n370 B.n369 585
R184 B.n369 B.n4 585
R185 B.n368 B.n148 585
R186 B.n368 B.n367 585
R187 B.n357 B.n149 585
R188 B.n360 B.n149 585
R189 B.n359 B.n358 585
R190 B.n361 B.n359 585
R191 B.n356 B.n154 585
R192 B.n154 B.n153 585
R193 B.n355 B.n354 585
R194 B.n354 B.n353 585
R195 B.n156 B.n155 585
R196 B.n346 B.n156 585
R197 B.n345 B.n344 585
R198 B.n347 B.n345 585
R199 B.n343 B.n161 585
R200 B.n161 B.n160 585
R201 B.n342 B.n341 585
R202 B.n341 B.n340 585
R203 B.n163 B.n162 585
R204 B.n164 B.n163 585
R205 B.n333 B.n332 585
R206 B.n334 B.n333 585
R207 B.n331 B.n169 585
R208 B.n169 B.n168 585
R209 B.n330 B.n329 585
R210 B.n329 B.n328 585
R211 B.n171 B.n170 585
R212 B.n172 B.n171 585
R213 B.n321 B.n320 585
R214 B.n322 B.n321 585
R215 B.n319 B.n177 585
R216 B.n177 B.n176 585
R217 B.n318 B.n317 585
R218 B.n317 B.n316 585
R219 B.n179 B.n178 585
R220 B.n180 B.n179 585
R221 B.n309 B.n308 585
R222 B.n310 B.n309 585
R223 B.n307 B.n184 585
R224 B.n188 B.n184 585
R225 B.n306 B.n305 585
R226 B.n305 B.n304 585
R227 B.n186 B.n185 585
R228 B.n187 B.n186 585
R229 B.n297 B.n296 585
R230 B.n298 B.n297 585
R231 B.n295 B.n193 585
R232 B.n193 B.n192 585
R233 B.n290 B.n289 585
R234 B.n288 B.n214 585
R235 B.n287 B.n213 585
R236 B.n292 B.n213 585
R237 B.n286 B.n285 585
R238 B.n284 B.n283 585
R239 B.n282 B.n281 585
R240 B.n280 B.n279 585
R241 B.n278 B.n277 585
R242 B.n276 B.n275 585
R243 B.n274 B.n273 585
R244 B.n272 B.n271 585
R245 B.n270 B.n269 585
R246 B.n268 B.n267 585
R247 B.n266 B.n265 585
R248 B.n263 B.n262 585
R249 B.n261 B.n260 585
R250 B.n259 B.n258 585
R251 B.n257 B.n256 585
R252 B.n255 B.n254 585
R253 B.n253 B.n252 585
R254 B.n251 B.n250 585
R255 B.n249 B.n248 585
R256 B.n247 B.n246 585
R257 B.n245 B.n244 585
R258 B.n242 B.n241 585
R259 B.n240 B.n239 585
R260 B.n238 B.n237 585
R261 B.n236 B.n235 585
R262 B.n234 B.n233 585
R263 B.n232 B.n231 585
R264 B.n230 B.n229 585
R265 B.n228 B.n227 585
R266 B.n226 B.n225 585
R267 B.n224 B.n223 585
R268 B.n222 B.n221 585
R269 B.n220 B.n219 585
R270 B.n195 B.n194 585
R271 B.n294 B.n293 585
R272 B.n293 B.n292 585
R273 B.n191 B.n190 585
R274 B.n192 B.n191 585
R275 B.n300 B.n299 585
R276 B.n299 B.n298 585
R277 B.n301 B.n189 585
R278 B.n189 B.n187 585
R279 B.n303 B.n302 585
R280 B.n304 B.n303 585
R281 B.n183 B.n182 585
R282 B.n188 B.n183 585
R283 B.n312 B.n311 585
R284 B.n311 B.n310 585
R285 B.n313 B.n181 585
R286 B.n181 B.n180 585
R287 B.n315 B.n314 585
R288 B.n316 B.n315 585
R289 B.n175 B.n174 585
R290 B.n176 B.n175 585
R291 B.n324 B.n323 585
R292 B.n323 B.n322 585
R293 B.n325 B.n173 585
R294 B.n173 B.n172 585
R295 B.n327 B.n326 585
R296 B.n328 B.n327 585
R297 B.n167 B.n166 585
R298 B.n168 B.n167 585
R299 B.n336 B.n335 585
R300 B.n335 B.n334 585
R301 B.n337 B.n165 585
R302 B.n165 B.n164 585
R303 B.n339 B.n338 585
R304 B.n340 B.n339 585
R305 B.n159 B.n158 585
R306 B.n160 B.n159 585
R307 B.n349 B.n348 585
R308 B.n348 B.n347 585
R309 B.n350 B.n157 585
R310 B.n346 B.n157 585
R311 B.n352 B.n351 585
R312 B.n353 B.n352 585
R313 B.n152 B.n151 585
R314 B.n153 B.n152 585
R315 B.n363 B.n362 585
R316 B.n362 B.n361 585
R317 B.n364 B.n150 585
R318 B.n360 B.n150 585
R319 B.n366 B.n365 585
R320 B.n367 B.n366 585
R321 B.n3 B.n0 585
R322 B.n4 B.n3 585
R323 B.n456 B.n1 585
R324 B.n457 B.n456 585
R325 B.n455 B.n454 585
R326 B.n455 B.n8 585
R327 B.n453 B.n9 585
R328 B.n12 B.n9 585
R329 B.n452 B.n451 585
R330 B.n451 B.n450 585
R331 B.n11 B.n10 585
R332 B.n449 B.n11 585
R333 B.n447 B.n446 585
R334 B.n448 B.n447 585
R335 B.n445 B.n16 585
R336 B.n19 B.n16 585
R337 B.n444 B.n443 585
R338 B.n443 B.n442 585
R339 B.n18 B.n17 585
R340 B.n441 B.n18 585
R341 B.n439 B.n438 585
R342 B.n440 B.n439 585
R343 B.n437 B.n24 585
R344 B.n24 B.n23 585
R345 B.n436 B.n435 585
R346 B.n435 B.n434 585
R347 B.n26 B.n25 585
R348 B.n433 B.n26 585
R349 B.n431 B.n430 585
R350 B.n432 B.n431 585
R351 B.n429 B.n31 585
R352 B.n31 B.n30 585
R353 B.n428 B.n427 585
R354 B.n427 B.n426 585
R355 B.n33 B.n32 585
R356 B.n425 B.n33 585
R357 B.n423 B.n422 585
R358 B.n424 B.n423 585
R359 B.n421 B.n38 585
R360 B.n38 B.n37 585
R361 B.n420 B.n419 585
R362 B.n419 B.n418 585
R363 B.n40 B.n39 585
R364 B.n417 B.n40 585
R365 B.n415 B.n414 585
R366 B.n416 B.n415 585
R367 B.n413 B.n45 585
R368 B.n45 B.n44 585
R369 B.n412 B.n411 585
R370 B.n411 B.n410 585
R371 B.n47 B.n46 585
R372 B.n409 B.n47 585
R373 B.n460 B.n459 585
R374 B.n458 B.n2 585
R375 B.n75 B.n47 569.379
R376 B.n406 B.n49 569.379
R377 B.n293 B.n193 569.379
R378 B.n290 B.n191 569.379
R379 B.n72 B.t8 277.858
R380 B.n69 B.t19 277.858
R381 B.n217 B.t12 277.858
R382 B.n215 B.t16 277.858
R383 B.n408 B.n407 256.663
R384 B.n408 B.n67 256.663
R385 B.n408 B.n66 256.663
R386 B.n408 B.n65 256.663
R387 B.n408 B.n64 256.663
R388 B.n408 B.n63 256.663
R389 B.n408 B.n62 256.663
R390 B.n408 B.n61 256.663
R391 B.n408 B.n60 256.663
R392 B.n408 B.n59 256.663
R393 B.n408 B.n58 256.663
R394 B.n408 B.n57 256.663
R395 B.n408 B.n56 256.663
R396 B.n408 B.n55 256.663
R397 B.n408 B.n54 256.663
R398 B.n408 B.n53 256.663
R399 B.n408 B.n52 256.663
R400 B.n408 B.n51 256.663
R401 B.n408 B.n50 256.663
R402 B.n292 B.n291 256.663
R403 B.n292 B.n196 256.663
R404 B.n292 B.n197 256.663
R405 B.n292 B.n198 256.663
R406 B.n292 B.n199 256.663
R407 B.n292 B.n200 256.663
R408 B.n292 B.n201 256.663
R409 B.n292 B.n202 256.663
R410 B.n292 B.n203 256.663
R411 B.n292 B.n204 256.663
R412 B.n292 B.n205 256.663
R413 B.n292 B.n206 256.663
R414 B.n292 B.n207 256.663
R415 B.n292 B.n208 256.663
R416 B.n292 B.n209 256.663
R417 B.n292 B.n210 256.663
R418 B.n292 B.n211 256.663
R419 B.n292 B.n212 256.663
R420 B.n462 B.n461 256.663
R421 B.n292 B.n192 193.512
R422 B.n409 B.n408 193.512
R423 B.n79 B.n78 163.367
R424 B.n83 B.n82 163.367
R425 B.n87 B.n86 163.367
R426 B.n91 B.n90 163.367
R427 B.n95 B.n94 163.367
R428 B.n99 B.n98 163.367
R429 B.n103 B.n102 163.367
R430 B.n107 B.n106 163.367
R431 B.n111 B.n110 163.367
R432 B.n115 B.n114 163.367
R433 B.n119 B.n118 163.367
R434 B.n123 B.n122 163.367
R435 B.n127 B.n126 163.367
R436 B.n131 B.n130 163.367
R437 B.n135 B.n134 163.367
R438 B.n139 B.n138 163.367
R439 B.n143 B.n142 163.367
R440 B.n145 B.n68 163.367
R441 B.n297 B.n193 163.367
R442 B.n297 B.n186 163.367
R443 B.n305 B.n186 163.367
R444 B.n305 B.n184 163.367
R445 B.n309 B.n184 163.367
R446 B.n309 B.n179 163.367
R447 B.n317 B.n179 163.367
R448 B.n317 B.n177 163.367
R449 B.n321 B.n177 163.367
R450 B.n321 B.n171 163.367
R451 B.n329 B.n171 163.367
R452 B.n329 B.n169 163.367
R453 B.n333 B.n169 163.367
R454 B.n333 B.n163 163.367
R455 B.n341 B.n163 163.367
R456 B.n341 B.n161 163.367
R457 B.n345 B.n161 163.367
R458 B.n345 B.n156 163.367
R459 B.n354 B.n156 163.367
R460 B.n354 B.n154 163.367
R461 B.n359 B.n154 163.367
R462 B.n359 B.n149 163.367
R463 B.n368 B.n149 163.367
R464 B.n369 B.n368 163.367
R465 B.n369 B.n5 163.367
R466 B.n6 B.n5 163.367
R467 B.n7 B.n6 163.367
R468 B.n375 B.n7 163.367
R469 B.n376 B.n375 163.367
R470 B.n376 B.n13 163.367
R471 B.n14 B.n13 163.367
R472 B.n15 B.n14 163.367
R473 B.n381 B.n15 163.367
R474 B.n381 B.n20 163.367
R475 B.n21 B.n20 163.367
R476 B.n22 B.n21 163.367
R477 B.n386 B.n22 163.367
R478 B.n386 B.n27 163.367
R479 B.n28 B.n27 163.367
R480 B.n29 B.n28 163.367
R481 B.n391 B.n29 163.367
R482 B.n391 B.n34 163.367
R483 B.n35 B.n34 163.367
R484 B.n36 B.n35 163.367
R485 B.n396 B.n36 163.367
R486 B.n396 B.n41 163.367
R487 B.n42 B.n41 163.367
R488 B.n43 B.n42 163.367
R489 B.n401 B.n43 163.367
R490 B.n401 B.n48 163.367
R491 B.n49 B.n48 163.367
R492 B.n214 B.n213 163.367
R493 B.n285 B.n213 163.367
R494 B.n283 B.n282 163.367
R495 B.n279 B.n278 163.367
R496 B.n275 B.n274 163.367
R497 B.n271 B.n270 163.367
R498 B.n267 B.n266 163.367
R499 B.n262 B.n261 163.367
R500 B.n258 B.n257 163.367
R501 B.n254 B.n253 163.367
R502 B.n250 B.n249 163.367
R503 B.n246 B.n245 163.367
R504 B.n241 B.n240 163.367
R505 B.n237 B.n236 163.367
R506 B.n233 B.n232 163.367
R507 B.n229 B.n228 163.367
R508 B.n225 B.n224 163.367
R509 B.n221 B.n220 163.367
R510 B.n293 B.n195 163.367
R511 B.n299 B.n191 163.367
R512 B.n299 B.n189 163.367
R513 B.n303 B.n189 163.367
R514 B.n303 B.n183 163.367
R515 B.n311 B.n183 163.367
R516 B.n311 B.n181 163.367
R517 B.n315 B.n181 163.367
R518 B.n315 B.n175 163.367
R519 B.n323 B.n175 163.367
R520 B.n323 B.n173 163.367
R521 B.n327 B.n173 163.367
R522 B.n327 B.n167 163.367
R523 B.n335 B.n167 163.367
R524 B.n335 B.n165 163.367
R525 B.n339 B.n165 163.367
R526 B.n339 B.n159 163.367
R527 B.n348 B.n159 163.367
R528 B.n348 B.n157 163.367
R529 B.n352 B.n157 163.367
R530 B.n352 B.n152 163.367
R531 B.n362 B.n152 163.367
R532 B.n362 B.n150 163.367
R533 B.n366 B.n150 163.367
R534 B.n366 B.n3 163.367
R535 B.n460 B.n3 163.367
R536 B.n456 B.n2 163.367
R537 B.n456 B.n455 163.367
R538 B.n455 B.n9 163.367
R539 B.n451 B.n9 163.367
R540 B.n451 B.n11 163.367
R541 B.n447 B.n11 163.367
R542 B.n447 B.n16 163.367
R543 B.n443 B.n16 163.367
R544 B.n443 B.n18 163.367
R545 B.n439 B.n18 163.367
R546 B.n439 B.n24 163.367
R547 B.n435 B.n24 163.367
R548 B.n435 B.n26 163.367
R549 B.n431 B.n26 163.367
R550 B.n431 B.n31 163.367
R551 B.n427 B.n31 163.367
R552 B.n427 B.n33 163.367
R553 B.n423 B.n33 163.367
R554 B.n423 B.n38 163.367
R555 B.n419 B.n38 163.367
R556 B.n419 B.n40 163.367
R557 B.n415 B.n40 163.367
R558 B.n415 B.n45 163.367
R559 B.n411 B.n45 163.367
R560 B.n411 B.n47 163.367
R561 B.n69 B.t20 99.4714
R562 B.n217 B.t15 99.4714
R563 B.n72 B.t10 99.4696
R564 B.n215 B.t18 99.4696
R565 B.n298 B.n192 93.3255
R566 B.n298 B.n187 93.3255
R567 B.n304 B.n187 93.3255
R568 B.n304 B.n188 93.3255
R569 B.n310 B.n180 93.3255
R570 B.n316 B.n180 93.3255
R571 B.n316 B.n176 93.3255
R572 B.n322 B.n176 93.3255
R573 B.n322 B.n172 93.3255
R574 B.n328 B.n172 93.3255
R575 B.n334 B.n168 93.3255
R576 B.n334 B.n164 93.3255
R577 B.n340 B.n164 93.3255
R578 B.n347 B.n160 93.3255
R579 B.n347 B.n346 93.3255
R580 B.n353 B.n153 93.3255
R581 B.n361 B.n153 93.3255
R582 B.n361 B.n360 93.3255
R583 B.n367 B.n4 93.3255
R584 B.n459 B.n4 93.3255
R585 B.n459 B.n458 93.3255
R586 B.n458 B.n457 93.3255
R587 B.n457 B.n8 93.3255
R588 B.n450 B.n12 93.3255
R589 B.n450 B.n449 93.3255
R590 B.n449 B.n448 93.3255
R591 B.n442 B.n19 93.3255
R592 B.n442 B.n441 93.3255
R593 B.n440 B.n23 93.3255
R594 B.n434 B.n23 93.3255
R595 B.n434 B.n433 93.3255
R596 B.n432 B.n30 93.3255
R597 B.n426 B.n30 93.3255
R598 B.n426 B.n425 93.3255
R599 B.n425 B.n424 93.3255
R600 B.n424 B.n37 93.3255
R601 B.n418 B.n37 93.3255
R602 B.n417 B.n416 93.3255
R603 B.n416 B.n44 93.3255
R604 B.n410 B.n44 93.3255
R605 B.n410 B.n409 93.3255
R606 B.t6 B.n160 86.4634
R607 B.n441 B.t7 86.4634
R608 B.n367 B.t4 80.9737
R609 B.t5 B.n8 80.9737
R610 B.n70 B.t21 76.1987
R611 B.n218 B.t14 76.1987
R612 B.n73 B.t11 76.1968
R613 B.n216 B.t17 76.1968
R614 B.n188 B.t13 75.484
R615 B.t9 B.n417 75.484
R616 B.n75 B.n50 71.676
R617 B.n79 B.n51 71.676
R618 B.n83 B.n52 71.676
R619 B.n87 B.n53 71.676
R620 B.n91 B.n54 71.676
R621 B.n95 B.n55 71.676
R622 B.n99 B.n56 71.676
R623 B.n103 B.n57 71.676
R624 B.n107 B.n58 71.676
R625 B.n111 B.n59 71.676
R626 B.n115 B.n60 71.676
R627 B.n119 B.n61 71.676
R628 B.n123 B.n62 71.676
R629 B.n127 B.n63 71.676
R630 B.n131 B.n64 71.676
R631 B.n135 B.n65 71.676
R632 B.n139 B.n66 71.676
R633 B.n143 B.n67 71.676
R634 B.n407 B.n68 71.676
R635 B.n407 B.n406 71.676
R636 B.n145 B.n67 71.676
R637 B.n142 B.n66 71.676
R638 B.n138 B.n65 71.676
R639 B.n134 B.n64 71.676
R640 B.n130 B.n63 71.676
R641 B.n126 B.n62 71.676
R642 B.n122 B.n61 71.676
R643 B.n118 B.n60 71.676
R644 B.n114 B.n59 71.676
R645 B.n110 B.n58 71.676
R646 B.n106 B.n57 71.676
R647 B.n102 B.n56 71.676
R648 B.n98 B.n55 71.676
R649 B.n94 B.n54 71.676
R650 B.n90 B.n53 71.676
R651 B.n86 B.n52 71.676
R652 B.n82 B.n51 71.676
R653 B.n78 B.n50 71.676
R654 B.n291 B.n290 71.676
R655 B.n285 B.n196 71.676
R656 B.n282 B.n197 71.676
R657 B.n278 B.n198 71.676
R658 B.n274 B.n199 71.676
R659 B.n270 B.n200 71.676
R660 B.n266 B.n201 71.676
R661 B.n261 B.n202 71.676
R662 B.n257 B.n203 71.676
R663 B.n253 B.n204 71.676
R664 B.n249 B.n205 71.676
R665 B.n245 B.n206 71.676
R666 B.n240 B.n207 71.676
R667 B.n236 B.n208 71.676
R668 B.n232 B.n209 71.676
R669 B.n228 B.n210 71.676
R670 B.n224 B.n211 71.676
R671 B.n220 B.n212 71.676
R672 B.n291 B.n214 71.676
R673 B.n283 B.n196 71.676
R674 B.n279 B.n197 71.676
R675 B.n275 B.n198 71.676
R676 B.n271 B.n199 71.676
R677 B.n267 B.n200 71.676
R678 B.n262 B.n201 71.676
R679 B.n258 B.n202 71.676
R680 B.n254 B.n203 71.676
R681 B.n250 B.n204 71.676
R682 B.n246 B.n205 71.676
R683 B.n241 B.n206 71.676
R684 B.n237 B.n207 71.676
R685 B.n233 B.n208 71.676
R686 B.n229 B.n209 71.676
R687 B.n225 B.n210 71.676
R688 B.n221 B.n211 71.676
R689 B.n212 B.n195 71.676
R690 B.n461 B.n460 71.676
R691 B.n461 B.n2 71.676
R692 B.n74 B.n73 59.5399
R693 B.n71 B.n70 59.5399
R694 B.n243 B.n218 59.5399
R695 B.n264 B.n216 59.5399
R696 B.n346 B.t1 56.27
R697 B.n19 B.t3 56.27
R698 B.n328 B.t2 50.7803
R699 B.t0 B.n432 50.7803
R700 B.t2 B.n168 42.5457
R701 B.n433 B.t0 42.5457
R702 B.n353 B.t1 37.056
R703 B.n448 B.t3 37.056
R704 B.n289 B.n190 36.9956
R705 B.n295 B.n294 36.9956
R706 B.n405 B.n404 36.9956
R707 B.n76 B.n46 36.9956
R708 B.n73 B.n72 23.2732
R709 B.n70 B.n69 23.2732
R710 B.n218 B.n217 23.2732
R711 B.n216 B.n215 23.2732
R712 B B.n462 18.0485
R713 B.n310 B.t13 17.842
R714 B.n418 B.t9 17.842
R715 B.n360 B.t4 12.3523
R716 B.n12 B.t5 12.3523
R717 B.n300 B.n190 10.6151
R718 B.n301 B.n300 10.6151
R719 B.n302 B.n301 10.6151
R720 B.n302 B.n182 10.6151
R721 B.n312 B.n182 10.6151
R722 B.n313 B.n312 10.6151
R723 B.n314 B.n313 10.6151
R724 B.n314 B.n174 10.6151
R725 B.n324 B.n174 10.6151
R726 B.n325 B.n324 10.6151
R727 B.n326 B.n325 10.6151
R728 B.n326 B.n166 10.6151
R729 B.n336 B.n166 10.6151
R730 B.n337 B.n336 10.6151
R731 B.n338 B.n337 10.6151
R732 B.n338 B.n158 10.6151
R733 B.n349 B.n158 10.6151
R734 B.n350 B.n349 10.6151
R735 B.n351 B.n350 10.6151
R736 B.n351 B.n151 10.6151
R737 B.n363 B.n151 10.6151
R738 B.n364 B.n363 10.6151
R739 B.n365 B.n364 10.6151
R740 B.n365 B.n0 10.6151
R741 B.n289 B.n288 10.6151
R742 B.n288 B.n287 10.6151
R743 B.n287 B.n286 10.6151
R744 B.n286 B.n284 10.6151
R745 B.n284 B.n281 10.6151
R746 B.n281 B.n280 10.6151
R747 B.n280 B.n277 10.6151
R748 B.n277 B.n276 10.6151
R749 B.n276 B.n273 10.6151
R750 B.n273 B.n272 10.6151
R751 B.n272 B.n269 10.6151
R752 B.n269 B.n268 10.6151
R753 B.n268 B.n265 10.6151
R754 B.n263 B.n260 10.6151
R755 B.n260 B.n259 10.6151
R756 B.n259 B.n256 10.6151
R757 B.n256 B.n255 10.6151
R758 B.n255 B.n252 10.6151
R759 B.n252 B.n251 10.6151
R760 B.n251 B.n248 10.6151
R761 B.n248 B.n247 10.6151
R762 B.n247 B.n244 10.6151
R763 B.n242 B.n239 10.6151
R764 B.n239 B.n238 10.6151
R765 B.n238 B.n235 10.6151
R766 B.n235 B.n234 10.6151
R767 B.n234 B.n231 10.6151
R768 B.n231 B.n230 10.6151
R769 B.n230 B.n227 10.6151
R770 B.n227 B.n226 10.6151
R771 B.n226 B.n223 10.6151
R772 B.n223 B.n222 10.6151
R773 B.n222 B.n219 10.6151
R774 B.n219 B.n194 10.6151
R775 B.n294 B.n194 10.6151
R776 B.n296 B.n295 10.6151
R777 B.n296 B.n185 10.6151
R778 B.n306 B.n185 10.6151
R779 B.n307 B.n306 10.6151
R780 B.n308 B.n307 10.6151
R781 B.n308 B.n178 10.6151
R782 B.n318 B.n178 10.6151
R783 B.n319 B.n318 10.6151
R784 B.n320 B.n319 10.6151
R785 B.n320 B.n170 10.6151
R786 B.n330 B.n170 10.6151
R787 B.n331 B.n330 10.6151
R788 B.n332 B.n331 10.6151
R789 B.n332 B.n162 10.6151
R790 B.n342 B.n162 10.6151
R791 B.n343 B.n342 10.6151
R792 B.n344 B.n343 10.6151
R793 B.n344 B.n155 10.6151
R794 B.n355 B.n155 10.6151
R795 B.n356 B.n355 10.6151
R796 B.n358 B.n356 10.6151
R797 B.n358 B.n357 10.6151
R798 B.n357 B.n148 10.6151
R799 B.n370 B.n148 10.6151
R800 B.n371 B.n370 10.6151
R801 B.n372 B.n371 10.6151
R802 B.n373 B.n372 10.6151
R803 B.n374 B.n373 10.6151
R804 B.n377 B.n374 10.6151
R805 B.n378 B.n377 10.6151
R806 B.n379 B.n378 10.6151
R807 B.n380 B.n379 10.6151
R808 B.n382 B.n380 10.6151
R809 B.n383 B.n382 10.6151
R810 B.n384 B.n383 10.6151
R811 B.n385 B.n384 10.6151
R812 B.n387 B.n385 10.6151
R813 B.n388 B.n387 10.6151
R814 B.n389 B.n388 10.6151
R815 B.n390 B.n389 10.6151
R816 B.n392 B.n390 10.6151
R817 B.n393 B.n392 10.6151
R818 B.n394 B.n393 10.6151
R819 B.n395 B.n394 10.6151
R820 B.n397 B.n395 10.6151
R821 B.n398 B.n397 10.6151
R822 B.n399 B.n398 10.6151
R823 B.n400 B.n399 10.6151
R824 B.n402 B.n400 10.6151
R825 B.n403 B.n402 10.6151
R826 B.n404 B.n403 10.6151
R827 B.n454 B.n1 10.6151
R828 B.n454 B.n453 10.6151
R829 B.n453 B.n452 10.6151
R830 B.n452 B.n10 10.6151
R831 B.n446 B.n10 10.6151
R832 B.n446 B.n445 10.6151
R833 B.n445 B.n444 10.6151
R834 B.n444 B.n17 10.6151
R835 B.n438 B.n17 10.6151
R836 B.n438 B.n437 10.6151
R837 B.n437 B.n436 10.6151
R838 B.n436 B.n25 10.6151
R839 B.n430 B.n25 10.6151
R840 B.n430 B.n429 10.6151
R841 B.n429 B.n428 10.6151
R842 B.n428 B.n32 10.6151
R843 B.n422 B.n32 10.6151
R844 B.n422 B.n421 10.6151
R845 B.n421 B.n420 10.6151
R846 B.n420 B.n39 10.6151
R847 B.n414 B.n39 10.6151
R848 B.n414 B.n413 10.6151
R849 B.n413 B.n412 10.6151
R850 B.n412 B.n46 10.6151
R851 B.n77 B.n76 10.6151
R852 B.n80 B.n77 10.6151
R853 B.n81 B.n80 10.6151
R854 B.n84 B.n81 10.6151
R855 B.n85 B.n84 10.6151
R856 B.n88 B.n85 10.6151
R857 B.n89 B.n88 10.6151
R858 B.n92 B.n89 10.6151
R859 B.n93 B.n92 10.6151
R860 B.n96 B.n93 10.6151
R861 B.n97 B.n96 10.6151
R862 B.n100 B.n97 10.6151
R863 B.n101 B.n100 10.6151
R864 B.n105 B.n104 10.6151
R865 B.n108 B.n105 10.6151
R866 B.n109 B.n108 10.6151
R867 B.n112 B.n109 10.6151
R868 B.n113 B.n112 10.6151
R869 B.n116 B.n113 10.6151
R870 B.n117 B.n116 10.6151
R871 B.n120 B.n117 10.6151
R872 B.n121 B.n120 10.6151
R873 B.n125 B.n124 10.6151
R874 B.n128 B.n125 10.6151
R875 B.n129 B.n128 10.6151
R876 B.n132 B.n129 10.6151
R877 B.n133 B.n132 10.6151
R878 B.n136 B.n133 10.6151
R879 B.n137 B.n136 10.6151
R880 B.n140 B.n137 10.6151
R881 B.n141 B.n140 10.6151
R882 B.n144 B.n141 10.6151
R883 B.n146 B.n144 10.6151
R884 B.n147 B.n146 10.6151
R885 B.n405 B.n147 10.6151
R886 B.n265 B.n264 9.36635
R887 B.n243 B.n242 9.36635
R888 B.n101 B.n74 9.36635
R889 B.n124 B.n71 9.36635
R890 B.n462 B.n0 8.11757
R891 B.n462 B.n1 8.11757
R892 B.n340 B.t6 6.86263
R893 B.t7 B.n440 6.86263
R894 B.n264 B.n263 1.24928
R895 B.n244 B.n243 1.24928
R896 B.n104 B.n74 1.24928
R897 B.n121 B.n71 1.24928
R898 VP.n30 VP.n29 161.3
R899 VP.n9 VP.n6 161.3
R900 VP.n11 VP.n10 161.3
R901 VP.n13 VP.n12 161.3
R902 VP.n14 VP.n4 161.3
R903 VP.n16 VP.n15 161.3
R904 VP.n28 VP.n0 161.3
R905 VP.n27 VP.n26 161.3
R906 VP.n25 VP.n24 161.3
R907 VP.n23 VP.n2 161.3
R908 VP.n21 VP.n20 161.3
R909 VP.n19 VP.n3 161.3
R910 VP.n18 VP.n17 161.3
R911 VP.n7 VP.t2 143.125
R912 VP.n17 VP.t7 121.055
R913 VP.n29 VP.t1 121.055
R914 VP.n15 VP.t5 121.055
R915 VP.n22 VP.t4 75.9016
R916 VP.n1 VP.t3 75.9016
R917 VP.n5 VP.t0 75.9016
R918 VP.n8 VP.t6 75.9016
R919 VP.n24 VP.n23 56.5617
R920 VP.n10 VP.n9 56.5617
R921 VP.n21 VP.n3 45.4209
R922 VP.n28 VP.n27 45.4209
R923 VP.n14 VP.n13 45.4209
R924 VP.n7 VP.n6 42.7264
R925 VP.n8 VP.n7 36.9171
R926 VP.n18 VP.n16 35.8187
R927 VP.n23 VP.n22 17.2148
R928 VP.n24 VP.n1 17.2148
R929 VP.n10 VP.n5 17.2148
R930 VP.n9 VP.n8 17.2148
R931 VP.n17 VP.n3 16.7975
R932 VP.n29 VP.n28 16.7975
R933 VP.n15 VP.n14 16.7975
R934 VP.n22 VP.n21 7.37805
R935 VP.n27 VP.n1 7.37805
R936 VP.n13 VP.n5 7.37805
R937 VP.n11 VP.n6 0.189894
R938 VP.n12 VP.n11 0.189894
R939 VP.n12 VP.n4 0.189894
R940 VP.n16 VP.n4 0.189894
R941 VP.n19 VP.n18 0.189894
R942 VP.n20 VP.n19 0.189894
R943 VP.n20 VP.n2 0.189894
R944 VP.n25 VP.n2 0.189894
R945 VP.n26 VP.n25 0.189894
R946 VP.n26 VP.n0 0.189894
R947 VP.n30 VP.n0 0.189894
R948 VP VP.n30 0.0516364
R949 VDD1 VDD1.n0 81.0161
R950 VDD1.n3 VDD1.n2 80.9024
R951 VDD1.n3 VDD1.n1 80.9024
R952 VDD1.n5 VDD1.n4 80.4406
R953 VDD1.n5 VDD1.n3 31.3155
R954 VDD1.n4 VDD1.t7 7.22678
R955 VDD1.n4 VDD1.t2 7.22678
R956 VDD1.n0 VDD1.t5 7.22678
R957 VDD1.n0 VDD1.t1 7.22678
R958 VDD1.n2 VDD1.t4 7.22678
R959 VDD1.n2 VDD1.t6 7.22678
R960 VDD1.n1 VDD1.t0 7.22678
R961 VDD1.n1 VDD1.t3 7.22678
R962 VDD1 VDD1.n5 0.459552
C0 VN VTAIL 1.99952f
C1 VN VDD1 0.153711f
C2 VN VDD2 1.7105f
C3 VTAIL VDD1 4.06931f
C4 VTAIL VDD2 4.11212f
C5 VN VP 3.83366f
C6 VP VTAIL 2.01362f
C7 VDD2 VDD1 0.908091f
C8 VP VDD1 1.8969f
C9 VP VDD2 0.341283f
C10 VDD2 B 2.766656f
C11 VDD1 B 3.010755f
C12 VTAIL B 3.611238f
C13 VN B 7.343754f
C14 VP B 6.515849f
C15 VDD1.t5 B 0.038424f
C16 VDD1.t1 B 0.038424f
C17 VDD1.n0 B 0.2822f
C18 VDD1.t0 B 0.038424f
C19 VDD1.t3 B 0.038424f
C20 VDD1.n1 B 0.281848f
C21 VDD1.t4 B 0.038424f
C22 VDD1.t6 B 0.038424f
C23 VDD1.n2 B 0.281848f
C24 VDD1.n3 B 1.23026f
C25 VDD1.t7 B 0.038424f
C26 VDD1.t2 B 0.038424f
C27 VDD1.n4 B 0.280569f
C28 VDD1.n5 B 1.14895f
C29 VP.n0 B 0.033932f
C30 VP.t3 B 0.199109f
C31 VP.n1 B 0.106626f
C32 VP.n2 B 0.033932f
C33 VP.t4 B 0.199109f
C34 VP.n3 B 0.014553f
C35 VP.n4 B 0.033932f
C36 VP.t5 B 0.24406f
C37 VP.t0 B 0.199109f
C38 VP.n5 B 0.106626f
C39 VP.n6 B 0.144826f
C40 VP.t6 B 0.199109f
C41 VP.t2 B 0.267189f
C42 VP.n7 B 0.140965f
C43 VP.n8 B 0.142912f
C44 VP.n9 B 0.040007f
C45 VP.n10 B 0.040007f
C46 VP.n11 B 0.033932f
C47 VP.n12 B 0.033932f
C48 VP.n13 B 0.043174f
C49 VP.n14 B 0.014553f
C50 VP.n15 B 0.141917f
C51 VP.n16 B 1.05667f
C52 VP.t7 B 0.24406f
C53 VP.n17 B 0.141917f
C54 VP.n18 B 1.09082f
C55 VP.n19 B 0.033932f
C56 VP.n20 B 0.033932f
C57 VP.n21 B 0.043174f
C58 VP.n22 B 0.106626f
C59 VP.n23 B 0.040007f
C60 VP.n24 B 0.040007f
C61 VP.n25 B 0.033932f
C62 VP.n26 B 0.033932f
C63 VP.n27 B 0.043174f
C64 VP.n28 B 0.014553f
C65 VP.t1 B 0.24406f
C66 VP.n29 B 0.141917f
C67 VP.n30 B 0.026296f
C68 VTAIL.t10 B 0.045676f
C69 VTAIL.t9 B 0.045676f
C70 VTAIL.n0 B 0.29409f
C71 VTAIL.n1 B 0.239805f
C72 VTAIL.t5 B 0.380693f
C73 VTAIL.n2 B 0.305754f
C74 VTAIL.t4 B 0.380693f
C75 VTAIL.n3 B 0.305754f
C76 VTAIL.t15 B 0.045676f
C77 VTAIL.t1 B 0.045676f
C78 VTAIL.n4 B 0.29409f
C79 VTAIL.n5 B 0.306167f
C80 VTAIL.t2 B 0.380693f
C81 VTAIL.n6 B 0.79125f
C82 VTAIL.t11 B 0.380694f
C83 VTAIL.n7 B 0.791249f
C84 VTAIL.t6 B 0.045676f
C85 VTAIL.t12 B 0.045676f
C86 VTAIL.n8 B 0.294091f
C87 VTAIL.n9 B 0.306166f
C88 VTAIL.t7 B 0.380694f
C89 VTAIL.n10 B 0.305753f
C90 VTAIL.t14 B 0.380694f
C91 VTAIL.n11 B 0.305753f
C92 VTAIL.t3 B 0.045676f
C93 VTAIL.t13 B 0.045676f
C94 VTAIL.n12 B 0.294091f
C95 VTAIL.n13 B 0.306166f
C96 VTAIL.t0 B 0.380693f
C97 VTAIL.n14 B 0.79125f
C98 VTAIL.t8 B 0.380693f
C99 VTAIL.n15 B 0.787295f
C100 VDD2.t2 B 0.039048f
C101 VDD2.t0 B 0.039048f
C102 VDD2.n0 B 0.286427f
C103 VDD2.t4 B 0.039048f
C104 VDD2.t1 B 0.039048f
C105 VDD2.n1 B 0.286427f
C106 VDD2.n2 B 1.2117f
C107 VDD2.t7 B 0.039048f
C108 VDD2.t3 B 0.039048f
C109 VDD2.n3 B 0.285129f
C110 VDD2.n4 B 1.14633f
C111 VDD2.t6 B 0.039048f
C112 VDD2.t5 B 0.039048f
C113 VDD2.n5 B 0.286412f
C114 VN.n0 B 0.02205f
C115 VN.t3 B 0.129387f
C116 VN.n1 B 0.069289f
C117 VN.n2 B 0.094112f
C118 VN.t2 B 0.129387f
C119 VN.t7 B 0.173627f
C120 VN.n3 B 0.091603f
C121 VN.n4 B 0.092868f
C122 VN.n5 B 0.025997f
C123 VN.n6 B 0.025997f
C124 VN.n7 B 0.02205f
C125 VN.n8 B 0.02205f
C126 VN.n9 B 0.028056f
C127 VN.n10 B 0.009457f
C128 VN.t4 B 0.158597f
C129 VN.n11 B 0.092221f
C130 VN.n12 B 0.017088f
C131 VN.n13 B 0.02205f
C132 VN.t6 B 0.129387f
C133 VN.n14 B 0.069289f
C134 VN.n15 B 0.094112f
C135 VN.t0 B 0.129387f
C136 VN.t5 B 0.173627f
C137 VN.n16 B 0.091603f
C138 VN.n17 B 0.092868f
C139 VN.n18 B 0.025997f
C140 VN.n19 B 0.025997f
C141 VN.n20 B 0.02205f
C142 VN.n21 B 0.02205f
C143 VN.n22 B 0.028056f
C144 VN.n23 B 0.009457f
C145 VN.t1 B 0.158597f
C146 VN.n24 B 0.092221f
C147 VN.n25 B 0.701287f
.ends

