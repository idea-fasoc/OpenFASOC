* NGSPICE file created from diff_pair_sample_1738.ext - technology: sky130A

.subckt diff_pair_sample_1738 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=4.3914 ps=23.3 w=11.26 l=3
X1 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=4.3914 ps=23.3 w=11.26 l=3
X2 VTAIL.t3 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X3 VTAIL.t12 VN.t1 VDD2.t6 B.t21 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=1.8579 ps=11.59 w=11.26 l=3
X4 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=0 ps=0 w=11.26 l=3
X5 VTAIL.t10 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=1.8579 ps=11.59 w=11.26 l=3
X6 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=0 ps=0 w=11.26 l=3
X7 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=0 ps=0 w=11.26 l=3
X8 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=0 ps=0 w=11.26 l=3
X9 VDD1.t5 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=4.3914 ps=23.3 w=11.26 l=3
X10 VDD2.t4 VN.t3 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X11 VTAIL.t8 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X12 VDD1.t4 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X13 VDD2.t2 VN.t5 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=4.3914 ps=23.3 w=11.26 l=3
X14 VTAIL.t14 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X15 VDD2.t0 VN.t7 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X16 VDD1.t3 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
X17 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=1.8579 ps=11.59 w=11.26 l=3
X18 VTAIL.t15 VP.t6 VDD1.t1 B.t21 sky130_fd_pr__nfet_01v8 ad=4.3914 pd=23.3 as=1.8579 ps=11.59 w=11.26 l=3
X19 VTAIL.t0 VP.t7 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8579 pd=11.59 as=1.8579 ps=11.59 w=11.26 l=3
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n50 VN.n49 161.3
R7 VN.n48 VN.n35 161.3
R8 VN.n47 VN.n46 161.3
R9 VN.n45 VN.n36 161.3
R10 VN.n44 VN.n43 161.3
R11 VN.n42 VN.n37 161.3
R12 VN.n41 VN.n40 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n19 VN.n18 161.3
R20 VN.n17 VN.n4 161.3
R21 VN.n16 VN.n15 161.3
R22 VN.n14 VN.n5 161.3
R23 VN.n13 VN.n12 161.3
R24 VN.n11 VN.n6 161.3
R25 VN.n10 VN.n9 161.3
R26 VN.n38 VN.t5 122.287
R27 VN.n7 VN.t2 122.287
R28 VN.n8 VN.t7 90.4558
R29 VN.n20 VN.t4 90.4558
R30 VN.n0 VN.t0 90.4558
R31 VN.n39 VN.t6 90.4558
R32 VN.n51 VN.t3 90.4558
R33 VN.n31 VN.t1 90.4558
R34 VN.n8 VN.n7 66.0722
R35 VN.n39 VN.n38 66.0722
R36 VN.n30 VN.n0 65.8996
R37 VN.n61 VN.n31 65.8996
R38 VN.n26 VN.n2 56.5617
R39 VN.n57 VN.n33 56.5617
R40 VN VN.n61 52.5587
R41 VN.n14 VN.n13 40.577
R42 VN.n15 VN.n14 40.577
R43 VN.n45 VN.n44 40.577
R44 VN.n46 VN.n45 40.577
R45 VN.n9 VN.n6 24.5923
R46 VN.n13 VN.n6 24.5923
R47 VN.n15 VN.n4 24.5923
R48 VN.n19 VN.n4 24.5923
R49 VN.n22 VN.n21 24.5923
R50 VN.n22 VN.n2 24.5923
R51 VN.n27 VN.n26 24.5923
R52 VN.n28 VN.n27 24.5923
R53 VN.n44 VN.n37 24.5923
R54 VN.n40 VN.n37 24.5923
R55 VN.n53 VN.n33 24.5923
R56 VN.n53 VN.n52 24.5923
R57 VN.n50 VN.n35 24.5923
R58 VN.n46 VN.n35 24.5923
R59 VN.n59 VN.n58 24.5923
R60 VN.n58 VN.n57 24.5923
R61 VN.n28 VN.n0 24.3464
R62 VN.n59 VN.n31 24.3464
R63 VN.n21 VN.n20 16.477
R64 VN.n52 VN.n51 16.477
R65 VN.n9 VN.n8 8.11581
R66 VN.n20 VN.n19 8.11581
R67 VN.n40 VN.n39 8.11581
R68 VN.n51 VN.n50 8.11581
R69 VN.n41 VN.n38 5.23312
R70 VN.n10 VN.n7 5.23312
R71 VN.n61 VN.n60 0.354861
R72 VN.n30 VN.n29 0.354861
R73 VN VN.n30 0.267071
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n49 VN.n34 0.189894
R80 VN.n49 VN.n48 0.189894
R81 VN.n48 VN.n47 0.189894
R82 VN.n47 VN.n36 0.189894
R83 VN.n43 VN.n36 0.189894
R84 VN.n43 VN.n42 0.189894
R85 VN.n42 VN.n41 0.189894
R86 VN.n11 VN.n10 0.189894
R87 VN.n12 VN.n11 0.189894
R88 VN.n12 VN.n5 0.189894
R89 VN.n16 VN.n5 0.189894
R90 VN.n17 VN.n16 0.189894
R91 VN.n18 VN.n17 0.189894
R92 VN.n18 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VTAIL.n502 VTAIL.n501 289.615
R99 VTAIL.n62 VTAIL.n61 289.615
R100 VTAIL.n124 VTAIL.n123 289.615
R101 VTAIL.n188 VTAIL.n187 289.615
R102 VTAIL.n440 VTAIL.n439 289.615
R103 VTAIL.n376 VTAIL.n375 289.615
R104 VTAIL.n314 VTAIL.n313 289.615
R105 VTAIL.n250 VTAIL.n249 289.615
R106 VTAIL.n463 VTAIL.n462 185
R107 VTAIL.n460 VTAIL.n459 185
R108 VTAIL.n469 VTAIL.n468 185
R109 VTAIL.n471 VTAIL.n470 185
R110 VTAIL.n456 VTAIL.n455 185
R111 VTAIL.n477 VTAIL.n476 185
R112 VTAIL.n479 VTAIL.n478 185
R113 VTAIL.n452 VTAIL.n451 185
R114 VTAIL.n485 VTAIL.n484 185
R115 VTAIL.n487 VTAIL.n486 185
R116 VTAIL.n448 VTAIL.n447 185
R117 VTAIL.n493 VTAIL.n492 185
R118 VTAIL.n495 VTAIL.n494 185
R119 VTAIL.n444 VTAIL.n443 185
R120 VTAIL.n501 VTAIL.n500 185
R121 VTAIL.n23 VTAIL.n22 185
R122 VTAIL.n20 VTAIL.n19 185
R123 VTAIL.n29 VTAIL.n28 185
R124 VTAIL.n31 VTAIL.n30 185
R125 VTAIL.n16 VTAIL.n15 185
R126 VTAIL.n37 VTAIL.n36 185
R127 VTAIL.n39 VTAIL.n38 185
R128 VTAIL.n12 VTAIL.n11 185
R129 VTAIL.n45 VTAIL.n44 185
R130 VTAIL.n47 VTAIL.n46 185
R131 VTAIL.n8 VTAIL.n7 185
R132 VTAIL.n53 VTAIL.n52 185
R133 VTAIL.n55 VTAIL.n54 185
R134 VTAIL.n4 VTAIL.n3 185
R135 VTAIL.n61 VTAIL.n60 185
R136 VTAIL.n85 VTAIL.n84 185
R137 VTAIL.n82 VTAIL.n81 185
R138 VTAIL.n91 VTAIL.n90 185
R139 VTAIL.n93 VTAIL.n92 185
R140 VTAIL.n78 VTAIL.n77 185
R141 VTAIL.n99 VTAIL.n98 185
R142 VTAIL.n101 VTAIL.n100 185
R143 VTAIL.n74 VTAIL.n73 185
R144 VTAIL.n107 VTAIL.n106 185
R145 VTAIL.n109 VTAIL.n108 185
R146 VTAIL.n70 VTAIL.n69 185
R147 VTAIL.n115 VTAIL.n114 185
R148 VTAIL.n117 VTAIL.n116 185
R149 VTAIL.n66 VTAIL.n65 185
R150 VTAIL.n123 VTAIL.n122 185
R151 VTAIL.n149 VTAIL.n148 185
R152 VTAIL.n146 VTAIL.n145 185
R153 VTAIL.n155 VTAIL.n154 185
R154 VTAIL.n157 VTAIL.n156 185
R155 VTAIL.n142 VTAIL.n141 185
R156 VTAIL.n163 VTAIL.n162 185
R157 VTAIL.n165 VTAIL.n164 185
R158 VTAIL.n138 VTAIL.n137 185
R159 VTAIL.n171 VTAIL.n170 185
R160 VTAIL.n173 VTAIL.n172 185
R161 VTAIL.n134 VTAIL.n133 185
R162 VTAIL.n179 VTAIL.n178 185
R163 VTAIL.n181 VTAIL.n180 185
R164 VTAIL.n130 VTAIL.n129 185
R165 VTAIL.n187 VTAIL.n186 185
R166 VTAIL.n439 VTAIL.n438 185
R167 VTAIL.n382 VTAIL.n381 185
R168 VTAIL.n433 VTAIL.n432 185
R169 VTAIL.n431 VTAIL.n430 185
R170 VTAIL.n386 VTAIL.n385 185
R171 VTAIL.n425 VTAIL.n424 185
R172 VTAIL.n423 VTAIL.n422 185
R173 VTAIL.n390 VTAIL.n389 185
R174 VTAIL.n417 VTAIL.n416 185
R175 VTAIL.n415 VTAIL.n414 185
R176 VTAIL.n394 VTAIL.n393 185
R177 VTAIL.n409 VTAIL.n408 185
R178 VTAIL.n407 VTAIL.n406 185
R179 VTAIL.n398 VTAIL.n397 185
R180 VTAIL.n401 VTAIL.n400 185
R181 VTAIL.n375 VTAIL.n374 185
R182 VTAIL.n318 VTAIL.n317 185
R183 VTAIL.n369 VTAIL.n368 185
R184 VTAIL.n367 VTAIL.n366 185
R185 VTAIL.n322 VTAIL.n321 185
R186 VTAIL.n361 VTAIL.n360 185
R187 VTAIL.n359 VTAIL.n358 185
R188 VTAIL.n326 VTAIL.n325 185
R189 VTAIL.n353 VTAIL.n352 185
R190 VTAIL.n351 VTAIL.n350 185
R191 VTAIL.n330 VTAIL.n329 185
R192 VTAIL.n345 VTAIL.n344 185
R193 VTAIL.n343 VTAIL.n342 185
R194 VTAIL.n334 VTAIL.n333 185
R195 VTAIL.n337 VTAIL.n336 185
R196 VTAIL.n313 VTAIL.n312 185
R197 VTAIL.n256 VTAIL.n255 185
R198 VTAIL.n307 VTAIL.n306 185
R199 VTAIL.n305 VTAIL.n304 185
R200 VTAIL.n260 VTAIL.n259 185
R201 VTAIL.n299 VTAIL.n298 185
R202 VTAIL.n297 VTAIL.n296 185
R203 VTAIL.n264 VTAIL.n263 185
R204 VTAIL.n291 VTAIL.n290 185
R205 VTAIL.n289 VTAIL.n288 185
R206 VTAIL.n268 VTAIL.n267 185
R207 VTAIL.n283 VTAIL.n282 185
R208 VTAIL.n281 VTAIL.n280 185
R209 VTAIL.n272 VTAIL.n271 185
R210 VTAIL.n275 VTAIL.n274 185
R211 VTAIL.n249 VTAIL.n248 185
R212 VTAIL.n192 VTAIL.n191 185
R213 VTAIL.n243 VTAIL.n242 185
R214 VTAIL.n241 VTAIL.n240 185
R215 VTAIL.n196 VTAIL.n195 185
R216 VTAIL.n235 VTAIL.n234 185
R217 VTAIL.n233 VTAIL.n232 185
R218 VTAIL.n200 VTAIL.n199 185
R219 VTAIL.n227 VTAIL.n226 185
R220 VTAIL.n225 VTAIL.n224 185
R221 VTAIL.n204 VTAIL.n203 185
R222 VTAIL.n219 VTAIL.n218 185
R223 VTAIL.n217 VTAIL.n216 185
R224 VTAIL.n208 VTAIL.n207 185
R225 VTAIL.n211 VTAIL.n210 185
R226 VTAIL.t9 VTAIL.n461 147.659
R227 VTAIL.t10 VTAIL.n21 147.659
R228 VTAIL.t6 VTAIL.n83 147.659
R229 VTAIL.t15 VTAIL.n147 147.659
R230 VTAIL.t1 VTAIL.n399 147.659
R231 VTAIL.t4 VTAIL.n335 147.659
R232 VTAIL.t11 VTAIL.n273 147.659
R233 VTAIL.t12 VTAIL.n209 147.659
R234 VTAIL.n462 VTAIL.n459 104.615
R235 VTAIL.n469 VTAIL.n459 104.615
R236 VTAIL.n470 VTAIL.n469 104.615
R237 VTAIL.n470 VTAIL.n455 104.615
R238 VTAIL.n477 VTAIL.n455 104.615
R239 VTAIL.n478 VTAIL.n477 104.615
R240 VTAIL.n478 VTAIL.n451 104.615
R241 VTAIL.n485 VTAIL.n451 104.615
R242 VTAIL.n486 VTAIL.n485 104.615
R243 VTAIL.n486 VTAIL.n447 104.615
R244 VTAIL.n493 VTAIL.n447 104.615
R245 VTAIL.n494 VTAIL.n493 104.615
R246 VTAIL.n494 VTAIL.n443 104.615
R247 VTAIL.n501 VTAIL.n443 104.615
R248 VTAIL.n22 VTAIL.n19 104.615
R249 VTAIL.n29 VTAIL.n19 104.615
R250 VTAIL.n30 VTAIL.n29 104.615
R251 VTAIL.n30 VTAIL.n15 104.615
R252 VTAIL.n37 VTAIL.n15 104.615
R253 VTAIL.n38 VTAIL.n37 104.615
R254 VTAIL.n38 VTAIL.n11 104.615
R255 VTAIL.n45 VTAIL.n11 104.615
R256 VTAIL.n46 VTAIL.n45 104.615
R257 VTAIL.n46 VTAIL.n7 104.615
R258 VTAIL.n53 VTAIL.n7 104.615
R259 VTAIL.n54 VTAIL.n53 104.615
R260 VTAIL.n54 VTAIL.n3 104.615
R261 VTAIL.n61 VTAIL.n3 104.615
R262 VTAIL.n84 VTAIL.n81 104.615
R263 VTAIL.n91 VTAIL.n81 104.615
R264 VTAIL.n92 VTAIL.n91 104.615
R265 VTAIL.n92 VTAIL.n77 104.615
R266 VTAIL.n99 VTAIL.n77 104.615
R267 VTAIL.n100 VTAIL.n99 104.615
R268 VTAIL.n100 VTAIL.n73 104.615
R269 VTAIL.n107 VTAIL.n73 104.615
R270 VTAIL.n108 VTAIL.n107 104.615
R271 VTAIL.n108 VTAIL.n69 104.615
R272 VTAIL.n115 VTAIL.n69 104.615
R273 VTAIL.n116 VTAIL.n115 104.615
R274 VTAIL.n116 VTAIL.n65 104.615
R275 VTAIL.n123 VTAIL.n65 104.615
R276 VTAIL.n148 VTAIL.n145 104.615
R277 VTAIL.n155 VTAIL.n145 104.615
R278 VTAIL.n156 VTAIL.n155 104.615
R279 VTAIL.n156 VTAIL.n141 104.615
R280 VTAIL.n163 VTAIL.n141 104.615
R281 VTAIL.n164 VTAIL.n163 104.615
R282 VTAIL.n164 VTAIL.n137 104.615
R283 VTAIL.n171 VTAIL.n137 104.615
R284 VTAIL.n172 VTAIL.n171 104.615
R285 VTAIL.n172 VTAIL.n133 104.615
R286 VTAIL.n179 VTAIL.n133 104.615
R287 VTAIL.n180 VTAIL.n179 104.615
R288 VTAIL.n180 VTAIL.n129 104.615
R289 VTAIL.n187 VTAIL.n129 104.615
R290 VTAIL.n439 VTAIL.n381 104.615
R291 VTAIL.n432 VTAIL.n381 104.615
R292 VTAIL.n432 VTAIL.n431 104.615
R293 VTAIL.n431 VTAIL.n385 104.615
R294 VTAIL.n424 VTAIL.n385 104.615
R295 VTAIL.n424 VTAIL.n423 104.615
R296 VTAIL.n423 VTAIL.n389 104.615
R297 VTAIL.n416 VTAIL.n389 104.615
R298 VTAIL.n416 VTAIL.n415 104.615
R299 VTAIL.n415 VTAIL.n393 104.615
R300 VTAIL.n408 VTAIL.n393 104.615
R301 VTAIL.n408 VTAIL.n407 104.615
R302 VTAIL.n407 VTAIL.n397 104.615
R303 VTAIL.n400 VTAIL.n397 104.615
R304 VTAIL.n375 VTAIL.n317 104.615
R305 VTAIL.n368 VTAIL.n317 104.615
R306 VTAIL.n368 VTAIL.n367 104.615
R307 VTAIL.n367 VTAIL.n321 104.615
R308 VTAIL.n360 VTAIL.n321 104.615
R309 VTAIL.n360 VTAIL.n359 104.615
R310 VTAIL.n359 VTAIL.n325 104.615
R311 VTAIL.n352 VTAIL.n325 104.615
R312 VTAIL.n352 VTAIL.n351 104.615
R313 VTAIL.n351 VTAIL.n329 104.615
R314 VTAIL.n344 VTAIL.n329 104.615
R315 VTAIL.n344 VTAIL.n343 104.615
R316 VTAIL.n343 VTAIL.n333 104.615
R317 VTAIL.n336 VTAIL.n333 104.615
R318 VTAIL.n313 VTAIL.n255 104.615
R319 VTAIL.n306 VTAIL.n255 104.615
R320 VTAIL.n306 VTAIL.n305 104.615
R321 VTAIL.n305 VTAIL.n259 104.615
R322 VTAIL.n298 VTAIL.n259 104.615
R323 VTAIL.n298 VTAIL.n297 104.615
R324 VTAIL.n297 VTAIL.n263 104.615
R325 VTAIL.n290 VTAIL.n263 104.615
R326 VTAIL.n290 VTAIL.n289 104.615
R327 VTAIL.n289 VTAIL.n267 104.615
R328 VTAIL.n282 VTAIL.n267 104.615
R329 VTAIL.n282 VTAIL.n281 104.615
R330 VTAIL.n281 VTAIL.n271 104.615
R331 VTAIL.n274 VTAIL.n271 104.615
R332 VTAIL.n249 VTAIL.n191 104.615
R333 VTAIL.n242 VTAIL.n191 104.615
R334 VTAIL.n242 VTAIL.n241 104.615
R335 VTAIL.n241 VTAIL.n195 104.615
R336 VTAIL.n234 VTAIL.n195 104.615
R337 VTAIL.n234 VTAIL.n233 104.615
R338 VTAIL.n233 VTAIL.n199 104.615
R339 VTAIL.n226 VTAIL.n199 104.615
R340 VTAIL.n226 VTAIL.n225 104.615
R341 VTAIL.n225 VTAIL.n203 104.615
R342 VTAIL.n218 VTAIL.n203 104.615
R343 VTAIL.n218 VTAIL.n217 104.615
R344 VTAIL.n217 VTAIL.n207 104.615
R345 VTAIL.n210 VTAIL.n207 104.615
R346 VTAIL.n462 VTAIL.t9 52.3082
R347 VTAIL.n22 VTAIL.t10 52.3082
R348 VTAIL.n84 VTAIL.t6 52.3082
R349 VTAIL.n148 VTAIL.t15 52.3082
R350 VTAIL.n400 VTAIL.t1 52.3082
R351 VTAIL.n336 VTAIL.t4 52.3082
R352 VTAIL.n274 VTAIL.t11 52.3082
R353 VTAIL.n210 VTAIL.t12 52.3082
R354 VTAIL.n379 VTAIL.n378 48.9724
R355 VTAIL.n253 VTAIL.n252 48.9724
R356 VTAIL.n1 VTAIL.n0 48.9723
R357 VTAIL.n127 VTAIL.n126 48.9723
R358 VTAIL.n503 VTAIL.n502 34.5126
R359 VTAIL.n63 VTAIL.n62 34.5126
R360 VTAIL.n125 VTAIL.n124 34.5126
R361 VTAIL.n189 VTAIL.n188 34.5126
R362 VTAIL.n441 VTAIL.n440 34.5126
R363 VTAIL.n377 VTAIL.n376 34.5126
R364 VTAIL.n315 VTAIL.n314 34.5126
R365 VTAIL.n251 VTAIL.n250 34.5126
R366 VTAIL.n503 VTAIL.n441 24.9445
R367 VTAIL.n251 VTAIL.n189 24.9445
R368 VTAIL.n463 VTAIL.n461 15.6677
R369 VTAIL.n23 VTAIL.n21 15.6677
R370 VTAIL.n85 VTAIL.n83 15.6677
R371 VTAIL.n149 VTAIL.n147 15.6677
R372 VTAIL.n401 VTAIL.n399 15.6677
R373 VTAIL.n337 VTAIL.n335 15.6677
R374 VTAIL.n275 VTAIL.n273 15.6677
R375 VTAIL.n211 VTAIL.n209 15.6677
R376 VTAIL.n464 VTAIL.n460 12.8005
R377 VTAIL.n24 VTAIL.n20 12.8005
R378 VTAIL.n86 VTAIL.n82 12.8005
R379 VTAIL.n150 VTAIL.n146 12.8005
R380 VTAIL.n402 VTAIL.n398 12.8005
R381 VTAIL.n338 VTAIL.n334 12.8005
R382 VTAIL.n276 VTAIL.n272 12.8005
R383 VTAIL.n212 VTAIL.n208 12.8005
R384 VTAIL.n468 VTAIL.n467 12.0247
R385 VTAIL.n28 VTAIL.n27 12.0247
R386 VTAIL.n90 VTAIL.n89 12.0247
R387 VTAIL.n154 VTAIL.n153 12.0247
R388 VTAIL.n406 VTAIL.n405 12.0247
R389 VTAIL.n342 VTAIL.n341 12.0247
R390 VTAIL.n280 VTAIL.n279 12.0247
R391 VTAIL.n216 VTAIL.n215 12.0247
R392 VTAIL.n471 VTAIL.n458 11.249
R393 VTAIL.n500 VTAIL.n442 11.249
R394 VTAIL.n31 VTAIL.n18 11.249
R395 VTAIL.n60 VTAIL.n2 11.249
R396 VTAIL.n93 VTAIL.n80 11.249
R397 VTAIL.n122 VTAIL.n64 11.249
R398 VTAIL.n157 VTAIL.n144 11.249
R399 VTAIL.n186 VTAIL.n128 11.249
R400 VTAIL.n438 VTAIL.n380 11.249
R401 VTAIL.n409 VTAIL.n396 11.249
R402 VTAIL.n374 VTAIL.n316 11.249
R403 VTAIL.n345 VTAIL.n332 11.249
R404 VTAIL.n312 VTAIL.n254 11.249
R405 VTAIL.n283 VTAIL.n270 11.249
R406 VTAIL.n248 VTAIL.n190 11.249
R407 VTAIL.n219 VTAIL.n206 11.249
R408 VTAIL.n472 VTAIL.n456 10.4732
R409 VTAIL.n499 VTAIL.n444 10.4732
R410 VTAIL.n32 VTAIL.n16 10.4732
R411 VTAIL.n59 VTAIL.n4 10.4732
R412 VTAIL.n94 VTAIL.n78 10.4732
R413 VTAIL.n121 VTAIL.n66 10.4732
R414 VTAIL.n158 VTAIL.n142 10.4732
R415 VTAIL.n185 VTAIL.n130 10.4732
R416 VTAIL.n437 VTAIL.n382 10.4732
R417 VTAIL.n410 VTAIL.n394 10.4732
R418 VTAIL.n373 VTAIL.n318 10.4732
R419 VTAIL.n346 VTAIL.n330 10.4732
R420 VTAIL.n311 VTAIL.n256 10.4732
R421 VTAIL.n284 VTAIL.n268 10.4732
R422 VTAIL.n247 VTAIL.n192 10.4732
R423 VTAIL.n220 VTAIL.n204 10.4732
R424 VTAIL.n476 VTAIL.n475 9.69747
R425 VTAIL.n496 VTAIL.n495 9.69747
R426 VTAIL.n36 VTAIL.n35 9.69747
R427 VTAIL.n56 VTAIL.n55 9.69747
R428 VTAIL.n98 VTAIL.n97 9.69747
R429 VTAIL.n118 VTAIL.n117 9.69747
R430 VTAIL.n162 VTAIL.n161 9.69747
R431 VTAIL.n182 VTAIL.n181 9.69747
R432 VTAIL.n434 VTAIL.n433 9.69747
R433 VTAIL.n414 VTAIL.n413 9.69747
R434 VTAIL.n370 VTAIL.n369 9.69747
R435 VTAIL.n350 VTAIL.n349 9.69747
R436 VTAIL.n308 VTAIL.n307 9.69747
R437 VTAIL.n288 VTAIL.n287 9.69747
R438 VTAIL.n244 VTAIL.n243 9.69747
R439 VTAIL.n224 VTAIL.n223 9.69747
R440 VTAIL.n498 VTAIL.n442 9.45567
R441 VTAIL.n58 VTAIL.n2 9.45567
R442 VTAIL.n120 VTAIL.n64 9.45567
R443 VTAIL.n184 VTAIL.n128 9.45567
R444 VTAIL.n436 VTAIL.n380 9.45567
R445 VTAIL.n372 VTAIL.n316 9.45567
R446 VTAIL.n310 VTAIL.n254 9.45567
R447 VTAIL.n246 VTAIL.n190 9.45567
R448 VTAIL.n450 VTAIL.n449 9.3005
R449 VTAIL.n489 VTAIL.n488 9.3005
R450 VTAIL.n491 VTAIL.n490 9.3005
R451 VTAIL.n446 VTAIL.n445 9.3005
R452 VTAIL.n497 VTAIL.n496 9.3005
R453 VTAIL.n499 VTAIL.n498 9.3005
R454 VTAIL.n481 VTAIL.n480 9.3005
R455 VTAIL.n454 VTAIL.n453 9.3005
R456 VTAIL.n475 VTAIL.n474 9.3005
R457 VTAIL.n473 VTAIL.n472 9.3005
R458 VTAIL.n458 VTAIL.n457 9.3005
R459 VTAIL.n467 VTAIL.n466 9.3005
R460 VTAIL.n465 VTAIL.n464 9.3005
R461 VTAIL.n483 VTAIL.n482 9.3005
R462 VTAIL.n10 VTAIL.n9 9.3005
R463 VTAIL.n49 VTAIL.n48 9.3005
R464 VTAIL.n51 VTAIL.n50 9.3005
R465 VTAIL.n6 VTAIL.n5 9.3005
R466 VTAIL.n57 VTAIL.n56 9.3005
R467 VTAIL.n59 VTAIL.n58 9.3005
R468 VTAIL.n41 VTAIL.n40 9.3005
R469 VTAIL.n14 VTAIL.n13 9.3005
R470 VTAIL.n35 VTAIL.n34 9.3005
R471 VTAIL.n33 VTAIL.n32 9.3005
R472 VTAIL.n18 VTAIL.n17 9.3005
R473 VTAIL.n27 VTAIL.n26 9.3005
R474 VTAIL.n25 VTAIL.n24 9.3005
R475 VTAIL.n43 VTAIL.n42 9.3005
R476 VTAIL.n72 VTAIL.n71 9.3005
R477 VTAIL.n111 VTAIL.n110 9.3005
R478 VTAIL.n113 VTAIL.n112 9.3005
R479 VTAIL.n68 VTAIL.n67 9.3005
R480 VTAIL.n119 VTAIL.n118 9.3005
R481 VTAIL.n121 VTAIL.n120 9.3005
R482 VTAIL.n103 VTAIL.n102 9.3005
R483 VTAIL.n76 VTAIL.n75 9.3005
R484 VTAIL.n97 VTAIL.n96 9.3005
R485 VTAIL.n95 VTAIL.n94 9.3005
R486 VTAIL.n80 VTAIL.n79 9.3005
R487 VTAIL.n89 VTAIL.n88 9.3005
R488 VTAIL.n87 VTAIL.n86 9.3005
R489 VTAIL.n105 VTAIL.n104 9.3005
R490 VTAIL.n136 VTAIL.n135 9.3005
R491 VTAIL.n175 VTAIL.n174 9.3005
R492 VTAIL.n177 VTAIL.n176 9.3005
R493 VTAIL.n132 VTAIL.n131 9.3005
R494 VTAIL.n183 VTAIL.n182 9.3005
R495 VTAIL.n185 VTAIL.n184 9.3005
R496 VTAIL.n167 VTAIL.n166 9.3005
R497 VTAIL.n140 VTAIL.n139 9.3005
R498 VTAIL.n161 VTAIL.n160 9.3005
R499 VTAIL.n159 VTAIL.n158 9.3005
R500 VTAIL.n144 VTAIL.n143 9.3005
R501 VTAIL.n153 VTAIL.n152 9.3005
R502 VTAIL.n151 VTAIL.n150 9.3005
R503 VTAIL.n169 VTAIL.n168 9.3005
R504 VTAIL.n437 VTAIL.n436 9.3005
R505 VTAIL.n435 VTAIL.n434 9.3005
R506 VTAIL.n384 VTAIL.n383 9.3005
R507 VTAIL.n429 VTAIL.n428 9.3005
R508 VTAIL.n427 VTAIL.n426 9.3005
R509 VTAIL.n388 VTAIL.n387 9.3005
R510 VTAIL.n421 VTAIL.n420 9.3005
R511 VTAIL.n419 VTAIL.n418 9.3005
R512 VTAIL.n392 VTAIL.n391 9.3005
R513 VTAIL.n413 VTAIL.n412 9.3005
R514 VTAIL.n411 VTAIL.n410 9.3005
R515 VTAIL.n396 VTAIL.n395 9.3005
R516 VTAIL.n405 VTAIL.n404 9.3005
R517 VTAIL.n403 VTAIL.n402 9.3005
R518 VTAIL.n363 VTAIL.n362 9.3005
R519 VTAIL.n365 VTAIL.n364 9.3005
R520 VTAIL.n320 VTAIL.n319 9.3005
R521 VTAIL.n371 VTAIL.n370 9.3005
R522 VTAIL.n373 VTAIL.n372 9.3005
R523 VTAIL.n324 VTAIL.n323 9.3005
R524 VTAIL.n357 VTAIL.n356 9.3005
R525 VTAIL.n355 VTAIL.n354 9.3005
R526 VTAIL.n328 VTAIL.n327 9.3005
R527 VTAIL.n349 VTAIL.n348 9.3005
R528 VTAIL.n347 VTAIL.n346 9.3005
R529 VTAIL.n332 VTAIL.n331 9.3005
R530 VTAIL.n341 VTAIL.n340 9.3005
R531 VTAIL.n339 VTAIL.n338 9.3005
R532 VTAIL.n301 VTAIL.n300 9.3005
R533 VTAIL.n303 VTAIL.n302 9.3005
R534 VTAIL.n258 VTAIL.n257 9.3005
R535 VTAIL.n309 VTAIL.n308 9.3005
R536 VTAIL.n311 VTAIL.n310 9.3005
R537 VTAIL.n262 VTAIL.n261 9.3005
R538 VTAIL.n295 VTAIL.n294 9.3005
R539 VTAIL.n293 VTAIL.n292 9.3005
R540 VTAIL.n266 VTAIL.n265 9.3005
R541 VTAIL.n287 VTAIL.n286 9.3005
R542 VTAIL.n285 VTAIL.n284 9.3005
R543 VTAIL.n270 VTAIL.n269 9.3005
R544 VTAIL.n279 VTAIL.n278 9.3005
R545 VTAIL.n277 VTAIL.n276 9.3005
R546 VTAIL.n237 VTAIL.n236 9.3005
R547 VTAIL.n239 VTAIL.n238 9.3005
R548 VTAIL.n194 VTAIL.n193 9.3005
R549 VTAIL.n245 VTAIL.n244 9.3005
R550 VTAIL.n247 VTAIL.n246 9.3005
R551 VTAIL.n198 VTAIL.n197 9.3005
R552 VTAIL.n231 VTAIL.n230 9.3005
R553 VTAIL.n229 VTAIL.n228 9.3005
R554 VTAIL.n202 VTAIL.n201 9.3005
R555 VTAIL.n223 VTAIL.n222 9.3005
R556 VTAIL.n221 VTAIL.n220 9.3005
R557 VTAIL.n206 VTAIL.n205 9.3005
R558 VTAIL.n215 VTAIL.n214 9.3005
R559 VTAIL.n213 VTAIL.n212 9.3005
R560 VTAIL.n479 VTAIL.n454 8.92171
R561 VTAIL.n492 VTAIL.n446 8.92171
R562 VTAIL.n39 VTAIL.n14 8.92171
R563 VTAIL.n52 VTAIL.n6 8.92171
R564 VTAIL.n101 VTAIL.n76 8.92171
R565 VTAIL.n114 VTAIL.n68 8.92171
R566 VTAIL.n165 VTAIL.n140 8.92171
R567 VTAIL.n178 VTAIL.n132 8.92171
R568 VTAIL.n430 VTAIL.n384 8.92171
R569 VTAIL.n417 VTAIL.n392 8.92171
R570 VTAIL.n366 VTAIL.n320 8.92171
R571 VTAIL.n353 VTAIL.n328 8.92171
R572 VTAIL.n304 VTAIL.n258 8.92171
R573 VTAIL.n291 VTAIL.n266 8.92171
R574 VTAIL.n240 VTAIL.n194 8.92171
R575 VTAIL.n227 VTAIL.n202 8.92171
R576 VTAIL.n480 VTAIL.n452 8.14595
R577 VTAIL.n491 VTAIL.n448 8.14595
R578 VTAIL.n40 VTAIL.n12 8.14595
R579 VTAIL.n51 VTAIL.n8 8.14595
R580 VTAIL.n102 VTAIL.n74 8.14595
R581 VTAIL.n113 VTAIL.n70 8.14595
R582 VTAIL.n166 VTAIL.n138 8.14595
R583 VTAIL.n177 VTAIL.n134 8.14595
R584 VTAIL.n429 VTAIL.n386 8.14595
R585 VTAIL.n418 VTAIL.n390 8.14595
R586 VTAIL.n365 VTAIL.n322 8.14595
R587 VTAIL.n354 VTAIL.n326 8.14595
R588 VTAIL.n303 VTAIL.n260 8.14595
R589 VTAIL.n292 VTAIL.n264 8.14595
R590 VTAIL.n239 VTAIL.n196 8.14595
R591 VTAIL.n228 VTAIL.n200 8.14595
R592 VTAIL.n484 VTAIL.n483 7.3702
R593 VTAIL.n488 VTAIL.n487 7.3702
R594 VTAIL.n44 VTAIL.n43 7.3702
R595 VTAIL.n48 VTAIL.n47 7.3702
R596 VTAIL.n106 VTAIL.n105 7.3702
R597 VTAIL.n110 VTAIL.n109 7.3702
R598 VTAIL.n170 VTAIL.n169 7.3702
R599 VTAIL.n174 VTAIL.n173 7.3702
R600 VTAIL.n426 VTAIL.n425 7.3702
R601 VTAIL.n422 VTAIL.n421 7.3702
R602 VTAIL.n362 VTAIL.n361 7.3702
R603 VTAIL.n358 VTAIL.n357 7.3702
R604 VTAIL.n300 VTAIL.n299 7.3702
R605 VTAIL.n296 VTAIL.n295 7.3702
R606 VTAIL.n236 VTAIL.n235 7.3702
R607 VTAIL.n232 VTAIL.n231 7.3702
R608 VTAIL.n484 VTAIL.n450 6.59444
R609 VTAIL.n487 VTAIL.n450 6.59444
R610 VTAIL.n44 VTAIL.n10 6.59444
R611 VTAIL.n47 VTAIL.n10 6.59444
R612 VTAIL.n106 VTAIL.n72 6.59444
R613 VTAIL.n109 VTAIL.n72 6.59444
R614 VTAIL.n170 VTAIL.n136 6.59444
R615 VTAIL.n173 VTAIL.n136 6.59444
R616 VTAIL.n425 VTAIL.n388 6.59444
R617 VTAIL.n422 VTAIL.n388 6.59444
R618 VTAIL.n361 VTAIL.n324 6.59444
R619 VTAIL.n358 VTAIL.n324 6.59444
R620 VTAIL.n299 VTAIL.n262 6.59444
R621 VTAIL.n296 VTAIL.n262 6.59444
R622 VTAIL.n235 VTAIL.n198 6.59444
R623 VTAIL.n232 VTAIL.n198 6.59444
R624 VTAIL.n483 VTAIL.n452 5.81868
R625 VTAIL.n488 VTAIL.n448 5.81868
R626 VTAIL.n43 VTAIL.n12 5.81868
R627 VTAIL.n48 VTAIL.n8 5.81868
R628 VTAIL.n105 VTAIL.n74 5.81868
R629 VTAIL.n110 VTAIL.n70 5.81868
R630 VTAIL.n169 VTAIL.n138 5.81868
R631 VTAIL.n174 VTAIL.n134 5.81868
R632 VTAIL.n426 VTAIL.n386 5.81868
R633 VTAIL.n421 VTAIL.n390 5.81868
R634 VTAIL.n362 VTAIL.n322 5.81868
R635 VTAIL.n357 VTAIL.n326 5.81868
R636 VTAIL.n300 VTAIL.n260 5.81868
R637 VTAIL.n295 VTAIL.n264 5.81868
R638 VTAIL.n236 VTAIL.n196 5.81868
R639 VTAIL.n231 VTAIL.n200 5.81868
R640 VTAIL.n480 VTAIL.n479 5.04292
R641 VTAIL.n492 VTAIL.n491 5.04292
R642 VTAIL.n40 VTAIL.n39 5.04292
R643 VTAIL.n52 VTAIL.n51 5.04292
R644 VTAIL.n102 VTAIL.n101 5.04292
R645 VTAIL.n114 VTAIL.n113 5.04292
R646 VTAIL.n166 VTAIL.n165 5.04292
R647 VTAIL.n178 VTAIL.n177 5.04292
R648 VTAIL.n430 VTAIL.n429 5.04292
R649 VTAIL.n418 VTAIL.n417 5.04292
R650 VTAIL.n366 VTAIL.n365 5.04292
R651 VTAIL.n354 VTAIL.n353 5.04292
R652 VTAIL.n304 VTAIL.n303 5.04292
R653 VTAIL.n292 VTAIL.n291 5.04292
R654 VTAIL.n240 VTAIL.n239 5.04292
R655 VTAIL.n228 VTAIL.n227 5.04292
R656 VTAIL.n465 VTAIL.n461 4.38563
R657 VTAIL.n25 VTAIL.n21 4.38563
R658 VTAIL.n87 VTAIL.n83 4.38563
R659 VTAIL.n151 VTAIL.n147 4.38563
R660 VTAIL.n403 VTAIL.n399 4.38563
R661 VTAIL.n339 VTAIL.n335 4.38563
R662 VTAIL.n277 VTAIL.n273 4.38563
R663 VTAIL.n213 VTAIL.n209 4.38563
R664 VTAIL.n476 VTAIL.n454 4.26717
R665 VTAIL.n495 VTAIL.n446 4.26717
R666 VTAIL.n36 VTAIL.n14 4.26717
R667 VTAIL.n55 VTAIL.n6 4.26717
R668 VTAIL.n98 VTAIL.n76 4.26717
R669 VTAIL.n117 VTAIL.n68 4.26717
R670 VTAIL.n162 VTAIL.n140 4.26717
R671 VTAIL.n181 VTAIL.n132 4.26717
R672 VTAIL.n433 VTAIL.n384 4.26717
R673 VTAIL.n414 VTAIL.n392 4.26717
R674 VTAIL.n369 VTAIL.n320 4.26717
R675 VTAIL.n350 VTAIL.n328 4.26717
R676 VTAIL.n307 VTAIL.n258 4.26717
R677 VTAIL.n288 VTAIL.n266 4.26717
R678 VTAIL.n243 VTAIL.n194 4.26717
R679 VTAIL.n224 VTAIL.n202 4.26717
R680 VTAIL.n475 VTAIL.n456 3.49141
R681 VTAIL.n496 VTAIL.n444 3.49141
R682 VTAIL.n35 VTAIL.n16 3.49141
R683 VTAIL.n56 VTAIL.n4 3.49141
R684 VTAIL.n97 VTAIL.n78 3.49141
R685 VTAIL.n118 VTAIL.n66 3.49141
R686 VTAIL.n161 VTAIL.n142 3.49141
R687 VTAIL.n182 VTAIL.n130 3.49141
R688 VTAIL.n434 VTAIL.n382 3.49141
R689 VTAIL.n413 VTAIL.n394 3.49141
R690 VTAIL.n370 VTAIL.n318 3.49141
R691 VTAIL.n349 VTAIL.n330 3.49141
R692 VTAIL.n308 VTAIL.n256 3.49141
R693 VTAIL.n287 VTAIL.n268 3.49141
R694 VTAIL.n244 VTAIL.n192 3.49141
R695 VTAIL.n223 VTAIL.n204 3.49141
R696 VTAIL.n253 VTAIL.n251 2.87119
R697 VTAIL.n315 VTAIL.n253 2.87119
R698 VTAIL.n379 VTAIL.n377 2.87119
R699 VTAIL.n441 VTAIL.n379 2.87119
R700 VTAIL.n189 VTAIL.n127 2.87119
R701 VTAIL.n127 VTAIL.n125 2.87119
R702 VTAIL.n63 VTAIL.n1 2.87119
R703 VTAIL VTAIL.n503 2.813
R704 VTAIL.n472 VTAIL.n471 2.71565
R705 VTAIL.n500 VTAIL.n499 2.71565
R706 VTAIL.n32 VTAIL.n31 2.71565
R707 VTAIL.n60 VTAIL.n59 2.71565
R708 VTAIL.n94 VTAIL.n93 2.71565
R709 VTAIL.n122 VTAIL.n121 2.71565
R710 VTAIL.n158 VTAIL.n157 2.71565
R711 VTAIL.n186 VTAIL.n185 2.71565
R712 VTAIL.n438 VTAIL.n437 2.71565
R713 VTAIL.n410 VTAIL.n409 2.71565
R714 VTAIL.n374 VTAIL.n373 2.71565
R715 VTAIL.n346 VTAIL.n345 2.71565
R716 VTAIL.n312 VTAIL.n311 2.71565
R717 VTAIL.n284 VTAIL.n283 2.71565
R718 VTAIL.n248 VTAIL.n247 2.71565
R719 VTAIL.n220 VTAIL.n219 2.71565
R720 VTAIL.n468 VTAIL.n458 1.93989
R721 VTAIL.n502 VTAIL.n442 1.93989
R722 VTAIL.n28 VTAIL.n18 1.93989
R723 VTAIL.n62 VTAIL.n2 1.93989
R724 VTAIL.n90 VTAIL.n80 1.93989
R725 VTAIL.n124 VTAIL.n64 1.93989
R726 VTAIL.n154 VTAIL.n144 1.93989
R727 VTAIL.n188 VTAIL.n128 1.93989
R728 VTAIL.n440 VTAIL.n380 1.93989
R729 VTAIL.n406 VTAIL.n396 1.93989
R730 VTAIL.n376 VTAIL.n316 1.93989
R731 VTAIL.n342 VTAIL.n332 1.93989
R732 VTAIL.n314 VTAIL.n254 1.93989
R733 VTAIL.n280 VTAIL.n270 1.93989
R734 VTAIL.n250 VTAIL.n190 1.93989
R735 VTAIL.n216 VTAIL.n206 1.93989
R736 VTAIL.n0 VTAIL.t13 1.75894
R737 VTAIL.n0 VTAIL.t8 1.75894
R738 VTAIL.n126 VTAIL.t5 1.75894
R739 VTAIL.n126 VTAIL.t0 1.75894
R740 VTAIL.n378 VTAIL.t2 1.75894
R741 VTAIL.n378 VTAIL.t3 1.75894
R742 VTAIL.n252 VTAIL.t7 1.75894
R743 VTAIL.n252 VTAIL.t14 1.75894
R744 VTAIL.n467 VTAIL.n460 1.16414
R745 VTAIL.n27 VTAIL.n20 1.16414
R746 VTAIL.n89 VTAIL.n82 1.16414
R747 VTAIL.n153 VTAIL.n146 1.16414
R748 VTAIL.n405 VTAIL.n398 1.16414
R749 VTAIL.n341 VTAIL.n334 1.16414
R750 VTAIL.n279 VTAIL.n272 1.16414
R751 VTAIL.n215 VTAIL.n208 1.16414
R752 VTAIL.n377 VTAIL.n315 0.470328
R753 VTAIL.n125 VTAIL.n63 0.470328
R754 VTAIL.n464 VTAIL.n463 0.388379
R755 VTAIL.n24 VTAIL.n23 0.388379
R756 VTAIL.n86 VTAIL.n85 0.388379
R757 VTAIL.n150 VTAIL.n149 0.388379
R758 VTAIL.n402 VTAIL.n401 0.388379
R759 VTAIL.n338 VTAIL.n337 0.388379
R760 VTAIL.n276 VTAIL.n275 0.388379
R761 VTAIL.n212 VTAIL.n211 0.388379
R762 VTAIL.n466 VTAIL.n465 0.155672
R763 VTAIL.n466 VTAIL.n457 0.155672
R764 VTAIL.n473 VTAIL.n457 0.155672
R765 VTAIL.n474 VTAIL.n473 0.155672
R766 VTAIL.n474 VTAIL.n453 0.155672
R767 VTAIL.n481 VTAIL.n453 0.155672
R768 VTAIL.n482 VTAIL.n481 0.155672
R769 VTAIL.n482 VTAIL.n449 0.155672
R770 VTAIL.n489 VTAIL.n449 0.155672
R771 VTAIL.n490 VTAIL.n489 0.155672
R772 VTAIL.n490 VTAIL.n445 0.155672
R773 VTAIL.n497 VTAIL.n445 0.155672
R774 VTAIL.n498 VTAIL.n497 0.155672
R775 VTAIL.n26 VTAIL.n25 0.155672
R776 VTAIL.n26 VTAIL.n17 0.155672
R777 VTAIL.n33 VTAIL.n17 0.155672
R778 VTAIL.n34 VTAIL.n33 0.155672
R779 VTAIL.n34 VTAIL.n13 0.155672
R780 VTAIL.n41 VTAIL.n13 0.155672
R781 VTAIL.n42 VTAIL.n41 0.155672
R782 VTAIL.n42 VTAIL.n9 0.155672
R783 VTAIL.n49 VTAIL.n9 0.155672
R784 VTAIL.n50 VTAIL.n49 0.155672
R785 VTAIL.n50 VTAIL.n5 0.155672
R786 VTAIL.n57 VTAIL.n5 0.155672
R787 VTAIL.n58 VTAIL.n57 0.155672
R788 VTAIL.n88 VTAIL.n87 0.155672
R789 VTAIL.n88 VTAIL.n79 0.155672
R790 VTAIL.n95 VTAIL.n79 0.155672
R791 VTAIL.n96 VTAIL.n95 0.155672
R792 VTAIL.n96 VTAIL.n75 0.155672
R793 VTAIL.n103 VTAIL.n75 0.155672
R794 VTAIL.n104 VTAIL.n103 0.155672
R795 VTAIL.n104 VTAIL.n71 0.155672
R796 VTAIL.n111 VTAIL.n71 0.155672
R797 VTAIL.n112 VTAIL.n111 0.155672
R798 VTAIL.n112 VTAIL.n67 0.155672
R799 VTAIL.n119 VTAIL.n67 0.155672
R800 VTAIL.n120 VTAIL.n119 0.155672
R801 VTAIL.n152 VTAIL.n151 0.155672
R802 VTAIL.n152 VTAIL.n143 0.155672
R803 VTAIL.n159 VTAIL.n143 0.155672
R804 VTAIL.n160 VTAIL.n159 0.155672
R805 VTAIL.n160 VTAIL.n139 0.155672
R806 VTAIL.n167 VTAIL.n139 0.155672
R807 VTAIL.n168 VTAIL.n167 0.155672
R808 VTAIL.n168 VTAIL.n135 0.155672
R809 VTAIL.n175 VTAIL.n135 0.155672
R810 VTAIL.n176 VTAIL.n175 0.155672
R811 VTAIL.n176 VTAIL.n131 0.155672
R812 VTAIL.n183 VTAIL.n131 0.155672
R813 VTAIL.n184 VTAIL.n183 0.155672
R814 VTAIL.n436 VTAIL.n435 0.155672
R815 VTAIL.n435 VTAIL.n383 0.155672
R816 VTAIL.n428 VTAIL.n383 0.155672
R817 VTAIL.n428 VTAIL.n427 0.155672
R818 VTAIL.n427 VTAIL.n387 0.155672
R819 VTAIL.n420 VTAIL.n387 0.155672
R820 VTAIL.n420 VTAIL.n419 0.155672
R821 VTAIL.n419 VTAIL.n391 0.155672
R822 VTAIL.n412 VTAIL.n391 0.155672
R823 VTAIL.n412 VTAIL.n411 0.155672
R824 VTAIL.n411 VTAIL.n395 0.155672
R825 VTAIL.n404 VTAIL.n395 0.155672
R826 VTAIL.n404 VTAIL.n403 0.155672
R827 VTAIL.n372 VTAIL.n371 0.155672
R828 VTAIL.n371 VTAIL.n319 0.155672
R829 VTAIL.n364 VTAIL.n319 0.155672
R830 VTAIL.n364 VTAIL.n363 0.155672
R831 VTAIL.n363 VTAIL.n323 0.155672
R832 VTAIL.n356 VTAIL.n323 0.155672
R833 VTAIL.n356 VTAIL.n355 0.155672
R834 VTAIL.n355 VTAIL.n327 0.155672
R835 VTAIL.n348 VTAIL.n327 0.155672
R836 VTAIL.n348 VTAIL.n347 0.155672
R837 VTAIL.n347 VTAIL.n331 0.155672
R838 VTAIL.n340 VTAIL.n331 0.155672
R839 VTAIL.n340 VTAIL.n339 0.155672
R840 VTAIL.n310 VTAIL.n309 0.155672
R841 VTAIL.n309 VTAIL.n257 0.155672
R842 VTAIL.n302 VTAIL.n257 0.155672
R843 VTAIL.n302 VTAIL.n301 0.155672
R844 VTAIL.n301 VTAIL.n261 0.155672
R845 VTAIL.n294 VTAIL.n261 0.155672
R846 VTAIL.n294 VTAIL.n293 0.155672
R847 VTAIL.n293 VTAIL.n265 0.155672
R848 VTAIL.n286 VTAIL.n265 0.155672
R849 VTAIL.n286 VTAIL.n285 0.155672
R850 VTAIL.n285 VTAIL.n269 0.155672
R851 VTAIL.n278 VTAIL.n269 0.155672
R852 VTAIL.n278 VTAIL.n277 0.155672
R853 VTAIL.n246 VTAIL.n245 0.155672
R854 VTAIL.n245 VTAIL.n193 0.155672
R855 VTAIL.n238 VTAIL.n193 0.155672
R856 VTAIL.n238 VTAIL.n237 0.155672
R857 VTAIL.n237 VTAIL.n197 0.155672
R858 VTAIL.n230 VTAIL.n197 0.155672
R859 VTAIL.n230 VTAIL.n229 0.155672
R860 VTAIL.n229 VTAIL.n201 0.155672
R861 VTAIL.n222 VTAIL.n201 0.155672
R862 VTAIL.n222 VTAIL.n221 0.155672
R863 VTAIL.n221 VTAIL.n205 0.155672
R864 VTAIL.n214 VTAIL.n205 0.155672
R865 VTAIL.n214 VTAIL.n213 0.155672
R866 VTAIL VTAIL.n1 0.0586897
R867 VDD2.n2 VDD2.n1 67.0311
R868 VDD2.n2 VDD2.n0 67.0311
R869 VDD2 VDD2.n5 67.0274
R870 VDD2.n4 VDD2.n3 65.6512
R871 VDD2.n4 VDD2.n2 46.3403
R872 VDD2.n5 VDD2.t1 1.75894
R873 VDD2.n5 VDD2.t2 1.75894
R874 VDD2.n3 VDD2.t6 1.75894
R875 VDD2.n3 VDD2.t4 1.75894
R876 VDD2.n1 VDD2.t3 1.75894
R877 VDD2.n1 VDD2.t7 1.75894
R878 VDD2.n0 VDD2.t5 1.75894
R879 VDD2.n0 VDD2.t0 1.75894
R880 VDD2 VDD2.n4 1.49403
R881 B.n909 B.n908 585
R882 B.n327 B.n148 585
R883 B.n326 B.n325 585
R884 B.n324 B.n323 585
R885 B.n322 B.n321 585
R886 B.n320 B.n319 585
R887 B.n318 B.n317 585
R888 B.n316 B.n315 585
R889 B.n314 B.n313 585
R890 B.n312 B.n311 585
R891 B.n310 B.n309 585
R892 B.n308 B.n307 585
R893 B.n306 B.n305 585
R894 B.n304 B.n303 585
R895 B.n302 B.n301 585
R896 B.n300 B.n299 585
R897 B.n298 B.n297 585
R898 B.n296 B.n295 585
R899 B.n294 B.n293 585
R900 B.n292 B.n291 585
R901 B.n290 B.n289 585
R902 B.n288 B.n287 585
R903 B.n286 B.n285 585
R904 B.n284 B.n283 585
R905 B.n282 B.n281 585
R906 B.n280 B.n279 585
R907 B.n278 B.n277 585
R908 B.n276 B.n275 585
R909 B.n274 B.n273 585
R910 B.n272 B.n271 585
R911 B.n270 B.n269 585
R912 B.n268 B.n267 585
R913 B.n266 B.n265 585
R914 B.n264 B.n263 585
R915 B.n262 B.n261 585
R916 B.n260 B.n259 585
R917 B.n258 B.n257 585
R918 B.n256 B.n255 585
R919 B.n254 B.n253 585
R920 B.n251 B.n250 585
R921 B.n249 B.n248 585
R922 B.n247 B.n246 585
R923 B.n245 B.n244 585
R924 B.n243 B.n242 585
R925 B.n241 B.n240 585
R926 B.n239 B.n238 585
R927 B.n237 B.n236 585
R928 B.n235 B.n234 585
R929 B.n233 B.n232 585
R930 B.n230 B.n229 585
R931 B.n228 B.n227 585
R932 B.n226 B.n225 585
R933 B.n224 B.n223 585
R934 B.n222 B.n221 585
R935 B.n220 B.n219 585
R936 B.n218 B.n217 585
R937 B.n216 B.n215 585
R938 B.n214 B.n213 585
R939 B.n212 B.n211 585
R940 B.n210 B.n209 585
R941 B.n208 B.n207 585
R942 B.n206 B.n205 585
R943 B.n204 B.n203 585
R944 B.n202 B.n201 585
R945 B.n200 B.n199 585
R946 B.n198 B.n197 585
R947 B.n196 B.n195 585
R948 B.n194 B.n193 585
R949 B.n192 B.n191 585
R950 B.n190 B.n189 585
R951 B.n188 B.n187 585
R952 B.n186 B.n185 585
R953 B.n184 B.n183 585
R954 B.n182 B.n181 585
R955 B.n180 B.n179 585
R956 B.n178 B.n177 585
R957 B.n176 B.n175 585
R958 B.n174 B.n173 585
R959 B.n172 B.n171 585
R960 B.n170 B.n169 585
R961 B.n168 B.n167 585
R962 B.n166 B.n165 585
R963 B.n164 B.n163 585
R964 B.n162 B.n161 585
R965 B.n160 B.n159 585
R966 B.n158 B.n157 585
R967 B.n156 B.n155 585
R968 B.n154 B.n153 585
R969 B.n907 B.n104 585
R970 B.n912 B.n104 585
R971 B.n906 B.n103 585
R972 B.n913 B.n103 585
R973 B.n905 B.n904 585
R974 B.n904 B.n99 585
R975 B.n903 B.n98 585
R976 B.n919 B.n98 585
R977 B.n902 B.n97 585
R978 B.n920 B.n97 585
R979 B.n901 B.n96 585
R980 B.n921 B.n96 585
R981 B.n900 B.n899 585
R982 B.n899 B.n92 585
R983 B.n898 B.n91 585
R984 B.n927 B.n91 585
R985 B.n897 B.n90 585
R986 B.n928 B.n90 585
R987 B.n896 B.n89 585
R988 B.n929 B.n89 585
R989 B.n895 B.n894 585
R990 B.n894 B.n85 585
R991 B.n893 B.n84 585
R992 B.n935 B.n84 585
R993 B.n892 B.n83 585
R994 B.n936 B.n83 585
R995 B.n891 B.n82 585
R996 B.n937 B.n82 585
R997 B.n890 B.n889 585
R998 B.n889 B.n78 585
R999 B.n888 B.n77 585
R1000 B.n943 B.n77 585
R1001 B.n887 B.n76 585
R1002 B.n944 B.n76 585
R1003 B.n886 B.n75 585
R1004 B.n945 B.n75 585
R1005 B.n885 B.n884 585
R1006 B.n884 B.n71 585
R1007 B.n883 B.n70 585
R1008 B.n951 B.n70 585
R1009 B.n882 B.n69 585
R1010 B.n952 B.n69 585
R1011 B.n881 B.n68 585
R1012 B.n953 B.n68 585
R1013 B.n880 B.n879 585
R1014 B.n879 B.n64 585
R1015 B.n878 B.n63 585
R1016 B.n959 B.n63 585
R1017 B.n877 B.n62 585
R1018 B.n960 B.n62 585
R1019 B.n876 B.n61 585
R1020 B.n961 B.n61 585
R1021 B.n875 B.n874 585
R1022 B.n874 B.n57 585
R1023 B.n873 B.n56 585
R1024 B.n967 B.n56 585
R1025 B.n872 B.n55 585
R1026 B.n968 B.n55 585
R1027 B.n871 B.n54 585
R1028 B.n969 B.n54 585
R1029 B.n870 B.n869 585
R1030 B.n869 B.n53 585
R1031 B.n868 B.n49 585
R1032 B.n975 B.n49 585
R1033 B.n867 B.n48 585
R1034 B.n976 B.n48 585
R1035 B.n866 B.n47 585
R1036 B.n977 B.n47 585
R1037 B.n865 B.n864 585
R1038 B.n864 B.n43 585
R1039 B.n863 B.n42 585
R1040 B.n983 B.n42 585
R1041 B.n862 B.n41 585
R1042 B.n984 B.n41 585
R1043 B.n861 B.n40 585
R1044 B.n985 B.n40 585
R1045 B.n860 B.n859 585
R1046 B.n859 B.n36 585
R1047 B.n858 B.n35 585
R1048 B.n991 B.n35 585
R1049 B.n857 B.n34 585
R1050 B.n992 B.n34 585
R1051 B.n856 B.n33 585
R1052 B.n993 B.n33 585
R1053 B.n855 B.n854 585
R1054 B.n854 B.n29 585
R1055 B.n853 B.n28 585
R1056 B.n999 B.n28 585
R1057 B.n852 B.n27 585
R1058 B.n1000 B.n27 585
R1059 B.n851 B.n26 585
R1060 B.n1001 B.n26 585
R1061 B.n850 B.n849 585
R1062 B.n849 B.n22 585
R1063 B.n848 B.n21 585
R1064 B.n1007 B.n21 585
R1065 B.n847 B.n20 585
R1066 B.n1008 B.n20 585
R1067 B.n846 B.n19 585
R1068 B.n1009 B.n19 585
R1069 B.n845 B.n844 585
R1070 B.n844 B.n18 585
R1071 B.n843 B.n14 585
R1072 B.n1015 B.n14 585
R1073 B.n842 B.n13 585
R1074 B.n1016 B.n13 585
R1075 B.n841 B.n12 585
R1076 B.n1017 B.n12 585
R1077 B.n840 B.n839 585
R1078 B.n839 B.n8 585
R1079 B.n838 B.n7 585
R1080 B.n1023 B.n7 585
R1081 B.n837 B.n6 585
R1082 B.n1024 B.n6 585
R1083 B.n836 B.n5 585
R1084 B.n1025 B.n5 585
R1085 B.n835 B.n834 585
R1086 B.n834 B.n4 585
R1087 B.n833 B.n328 585
R1088 B.n833 B.n832 585
R1089 B.n823 B.n329 585
R1090 B.n330 B.n329 585
R1091 B.n825 B.n824 585
R1092 B.n826 B.n825 585
R1093 B.n822 B.n335 585
R1094 B.n335 B.n334 585
R1095 B.n821 B.n820 585
R1096 B.n820 B.n819 585
R1097 B.n337 B.n336 585
R1098 B.n812 B.n337 585
R1099 B.n811 B.n810 585
R1100 B.n813 B.n811 585
R1101 B.n809 B.n342 585
R1102 B.n342 B.n341 585
R1103 B.n808 B.n807 585
R1104 B.n807 B.n806 585
R1105 B.n344 B.n343 585
R1106 B.n345 B.n344 585
R1107 B.n799 B.n798 585
R1108 B.n800 B.n799 585
R1109 B.n797 B.n350 585
R1110 B.n350 B.n349 585
R1111 B.n796 B.n795 585
R1112 B.n795 B.n794 585
R1113 B.n352 B.n351 585
R1114 B.n353 B.n352 585
R1115 B.n787 B.n786 585
R1116 B.n788 B.n787 585
R1117 B.n785 B.n357 585
R1118 B.n361 B.n357 585
R1119 B.n784 B.n783 585
R1120 B.n783 B.n782 585
R1121 B.n359 B.n358 585
R1122 B.n360 B.n359 585
R1123 B.n775 B.n774 585
R1124 B.n776 B.n775 585
R1125 B.n773 B.n366 585
R1126 B.n366 B.n365 585
R1127 B.n772 B.n771 585
R1128 B.n771 B.n770 585
R1129 B.n368 B.n367 585
R1130 B.n369 B.n368 585
R1131 B.n763 B.n762 585
R1132 B.n764 B.n763 585
R1133 B.n761 B.n374 585
R1134 B.n374 B.n373 585
R1135 B.n760 B.n759 585
R1136 B.n759 B.n758 585
R1137 B.n376 B.n375 585
R1138 B.n751 B.n376 585
R1139 B.n750 B.n749 585
R1140 B.n752 B.n750 585
R1141 B.n748 B.n381 585
R1142 B.n381 B.n380 585
R1143 B.n747 B.n746 585
R1144 B.n746 B.n745 585
R1145 B.n383 B.n382 585
R1146 B.n384 B.n383 585
R1147 B.n738 B.n737 585
R1148 B.n739 B.n738 585
R1149 B.n736 B.n389 585
R1150 B.n389 B.n388 585
R1151 B.n735 B.n734 585
R1152 B.n734 B.n733 585
R1153 B.n391 B.n390 585
R1154 B.n392 B.n391 585
R1155 B.n726 B.n725 585
R1156 B.n727 B.n726 585
R1157 B.n724 B.n397 585
R1158 B.n397 B.n396 585
R1159 B.n723 B.n722 585
R1160 B.n722 B.n721 585
R1161 B.n399 B.n398 585
R1162 B.n400 B.n399 585
R1163 B.n714 B.n713 585
R1164 B.n715 B.n714 585
R1165 B.n712 B.n405 585
R1166 B.n405 B.n404 585
R1167 B.n711 B.n710 585
R1168 B.n710 B.n709 585
R1169 B.n407 B.n406 585
R1170 B.n408 B.n407 585
R1171 B.n702 B.n701 585
R1172 B.n703 B.n702 585
R1173 B.n700 B.n413 585
R1174 B.n413 B.n412 585
R1175 B.n699 B.n698 585
R1176 B.n698 B.n697 585
R1177 B.n415 B.n414 585
R1178 B.n416 B.n415 585
R1179 B.n690 B.n689 585
R1180 B.n691 B.n690 585
R1181 B.n688 B.n420 585
R1182 B.n424 B.n420 585
R1183 B.n687 B.n686 585
R1184 B.n686 B.n685 585
R1185 B.n422 B.n421 585
R1186 B.n423 B.n422 585
R1187 B.n678 B.n677 585
R1188 B.n679 B.n678 585
R1189 B.n676 B.n429 585
R1190 B.n429 B.n428 585
R1191 B.n675 B.n674 585
R1192 B.n674 B.n673 585
R1193 B.n431 B.n430 585
R1194 B.n432 B.n431 585
R1195 B.n666 B.n665 585
R1196 B.n667 B.n666 585
R1197 B.n664 B.n437 585
R1198 B.n437 B.n436 585
R1199 B.n659 B.n658 585
R1200 B.n657 B.n483 585
R1201 B.n656 B.n482 585
R1202 B.n661 B.n482 585
R1203 B.n655 B.n654 585
R1204 B.n653 B.n652 585
R1205 B.n651 B.n650 585
R1206 B.n649 B.n648 585
R1207 B.n647 B.n646 585
R1208 B.n645 B.n644 585
R1209 B.n643 B.n642 585
R1210 B.n641 B.n640 585
R1211 B.n639 B.n638 585
R1212 B.n637 B.n636 585
R1213 B.n635 B.n634 585
R1214 B.n633 B.n632 585
R1215 B.n631 B.n630 585
R1216 B.n629 B.n628 585
R1217 B.n627 B.n626 585
R1218 B.n625 B.n624 585
R1219 B.n623 B.n622 585
R1220 B.n621 B.n620 585
R1221 B.n619 B.n618 585
R1222 B.n617 B.n616 585
R1223 B.n615 B.n614 585
R1224 B.n613 B.n612 585
R1225 B.n611 B.n610 585
R1226 B.n609 B.n608 585
R1227 B.n607 B.n606 585
R1228 B.n605 B.n604 585
R1229 B.n603 B.n602 585
R1230 B.n601 B.n600 585
R1231 B.n599 B.n598 585
R1232 B.n597 B.n596 585
R1233 B.n595 B.n594 585
R1234 B.n593 B.n592 585
R1235 B.n591 B.n590 585
R1236 B.n589 B.n588 585
R1237 B.n587 B.n586 585
R1238 B.n585 B.n584 585
R1239 B.n583 B.n582 585
R1240 B.n581 B.n580 585
R1241 B.n579 B.n578 585
R1242 B.n577 B.n576 585
R1243 B.n575 B.n574 585
R1244 B.n573 B.n572 585
R1245 B.n571 B.n570 585
R1246 B.n569 B.n568 585
R1247 B.n567 B.n566 585
R1248 B.n565 B.n564 585
R1249 B.n563 B.n562 585
R1250 B.n561 B.n560 585
R1251 B.n559 B.n558 585
R1252 B.n557 B.n556 585
R1253 B.n555 B.n554 585
R1254 B.n553 B.n552 585
R1255 B.n551 B.n550 585
R1256 B.n549 B.n548 585
R1257 B.n547 B.n546 585
R1258 B.n545 B.n544 585
R1259 B.n543 B.n542 585
R1260 B.n541 B.n540 585
R1261 B.n539 B.n538 585
R1262 B.n537 B.n536 585
R1263 B.n535 B.n534 585
R1264 B.n533 B.n532 585
R1265 B.n531 B.n530 585
R1266 B.n529 B.n528 585
R1267 B.n527 B.n526 585
R1268 B.n525 B.n524 585
R1269 B.n523 B.n522 585
R1270 B.n521 B.n520 585
R1271 B.n519 B.n518 585
R1272 B.n517 B.n516 585
R1273 B.n515 B.n514 585
R1274 B.n513 B.n512 585
R1275 B.n511 B.n510 585
R1276 B.n509 B.n508 585
R1277 B.n507 B.n506 585
R1278 B.n505 B.n504 585
R1279 B.n503 B.n502 585
R1280 B.n501 B.n500 585
R1281 B.n499 B.n498 585
R1282 B.n497 B.n496 585
R1283 B.n495 B.n494 585
R1284 B.n493 B.n492 585
R1285 B.n491 B.n490 585
R1286 B.n439 B.n438 585
R1287 B.n663 B.n662 585
R1288 B.n662 B.n661 585
R1289 B.n435 B.n434 585
R1290 B.n436 B.n435 585
R1291 B.n669 B.n668 585
R1292 B.n668 B.n667 585
R1293 B.n670 B.n433 585
R1294 B.n433 B.n432 585
R1295 B.n672 B.n671 585
R1296 B.n673 B.n672 585
R1297 B.n427 B.n426 585
R1298 B.n428 B.n427 585
R1299 B.n681 B.n680 585
R1300 B.n680 B.n679 585
R1301 B.n682 B.n425 585
R1302 B.n425 B.n423 585
R1303 B.n684 B.n683 585
R1304 B.n685 B.n684 585
R1305 B.n419 B.n418 585
R1306 B.n424 B.n419 585
R1307 B.n693 B.n692 585
R1308 B.n692 B.n691 585
R1309 B.n694 B.n417 585
R1310 B.n417 B.n416 585
R1311 B.n696 B.n695 585
R1312 B.n697 B.n696 585
R1313 B.n411 B.n410 585
R1314 B.n412 B.n411 585
R1315 B.n705 B.n704 585
R1316 B.n704 B.n703 585
R1317 B.n706 B.n409 585
R1318 B.n409 B.n408 585
R1319 B.n708 B.n707 585
R1320 B.n709 B.n708 585
R1321 B.n403 B.n402 585
R1322 B.n404 B.n403 585
R1323 B.n717 B.n716 585
R1324 B.n716 B.n715 585
R1325 B.n718 B.n401 585
R1326 B.n401 B.n400 585
R1327 B.n720 B.n719 585
R1328 B.n721 B.n720 585
R1329 B.n395 B.n394 585
R1330 B.n396 B.n395 585
R1331 B.n729 B.n728 585
R1332 B.n728 B.n727 585
R1333 B.n730 B.n393 585
R1334 B.n393 B.n392 585
R1335 B.n732 B.n731 585
R1336 B.n733 B.n732 585
R1337 B.n387 B.n386 585
R1338 B.n388 B.n387 585
R1339 B.n741 B.n740 585
R1340 B.n740 B.n739 585
R1341 B.n742 B.n385 585
R1342 B.n385 B.n384 585
R1343 B.n744 B.n743 585
R1344 B.n745 B.n744 585
R1345 B.n379 B.n378 585
R1346 B.n380 B.n379 585
R1347 B.n754 B.n753 585
R1348 B.n753 B.n752 585
R1349 B.n755 B.n377 585
R1350 B.n751 B.n377 585
R1351 B.n757 B.n756 585
R1352 B.n758 B.n757 585
R1353 B.n372 B.n371 585
R1354 B.n373 B.n372 585
R1355 B.n766 B.n765 585
R1356 B.n765 B.n764 585
R1357 B.n767 B.n370 585
R1358 B.n370 B.n369 585
R1359 B.n769 B.n768 585
R1360 B.n770 B.n769 585
R1361 B.n364 B.n363 585
R1362 B.n365 B.n364 585
R1363 B.n778 B.n777 585
R1364 B.n777 B.n776 585
R1365 B.n779 B.n362 585
R1366 B.n362 B.n360 585
R1367 B.n781 B.n780 585
R1368 B.n782 B.n781 585
R1369 B.n356 B.n355 585
R1370 B.n361 B.n356 585
R1371 B.n790 B.n789 585
R1372 B.n789 B.n788 585
R1373 B.n791 B.n354 585
R1374 B.n354 B.n353 585
R1375 B.n793 B.n792 585
R1376 B.n794 B.n793 585
R1377 B.n348 B.n347 585
R1378 B.n349 B.n348 585
R1379 B.n802 B.n801 585
R1380 B.n801 B.n800 585
R1381 B.n803 B.n346 585
R1382 B.n346 B.n345 585
R1383 B.n805 B.n804 585
R1384 B.n806 B.n805 585
R1385 B.n340 B.n339 585
R1386 B.n341 B.n340 585
R1387 B.n815 B.n814 585
R1388 B.n814 B.n813 585
R1389 B.n816 B.n338 585
R1390 B.n812 B.n338 585
R1391 B.n818 B.n817 585
R1392 B.n819 B.n818 585
R1393 B.n333 B.n332 585
R1394 B.n334 B.n333 585
R1395 B.n828 B.n827 585
R1396 B.n827 B.n826 585
R1397 B.n829 B.n331 585
R1398 B.n331 B.n330 585
R1399 B.n831 B.n830 585
R1400 B.n832 B.n831 585
R1401 B.n2 B.n0 585
R1402 B.n4 B.n2 585
R1403 B.n3 B.n1 585
R1404 B.n1024 B.n3 585
R1405 B.n1022 B.n1021 585
R1406 B.n1023 B.n1022 585
R1407 B.n1020 B.n9 585
R1408 B.n9 B.n8 585
R1409 B.n1019 B.n1018 585
R1410 B.n1018 B.n1017 585
R1411 B.n11 B.n10 585
R1412 B.n1016 B.n11 585
R1413 B.n1014 B.n1013 585
R1414 B.n1015 B.n1014 585
R1415 B.n1012 B.n15 585
R1416 B.n18 B.n15 585
R1417 B.n1011 B.n1010 585
R1418 B.n1010 B.n1009 585
R1419 B.n17 B.n16 585
R1420 B.n1008 B.n17 585
R1421 B.n1006 B.n1005 585
R1422 B.n1007 B.n1006 585
R1423 B.n1004 B.n23 585
R1424 B.n23 B.n22 585
R1425 B.n1003 B.n1002 585
R1426 B.n1002 B.n1001 585
R1427 B.n25 B.n24 585
R1428 B.n1000 B.n25 585
R1429 B.n998 B.n997 585
R1430 B.n999 B.n998 585
R1431 B.n996 B.n30 585
R1432 B.n30 B.n29 585
R1433 B.n995 B.n994 585
R1434 B.n994 B.n993 585
R1435 B.n32 B.n31 585
R1436 B.n992 B.n32 585
R1437 B.n990 B.n989 585
R1438 B.n991 B.n990 585
R1439 B.n988 B.n37 585
R1440 B.n37 B.n36 585
R1441 B.n987 B.n986 585
R1442 B.n986 B.n985 585
R1443 B.n39 B.n38 585
R1444 B.n984 B.n39 585
R1445 B.n982 B.n981 585
R1446 B.n983 B.n982 585
R1447 B.n980 B.n44 585
R1448 B.n44 B.n43 585
R1449 B.n979 B.n978 585
R1450 B.n978 B.n977 585
R1451 B.n46 B.n45 585
R1452 B.n976 B.n46 585
R1453 B.n974 B.n973 585
R1454 B.n975 B.n974 585
R1455 B.n972 B.n50 585
R1456 B.n53 B.n50 585
R1457 B.n971 B.n970 585
R1458 B.n970 B.n969 585
R1459 B.n52 B.n51 585
R1460 B.n968 B.n52 585
R1461 B.n966 B.n965 585
R1462 B.n967 B.n966 585
R1463 B.n964 B.n58 585
R1464 B.n58 B.n57 585
R1465 B.n963 B.n962 585
R1466 B.n962 B.n961 585
R1467 B.n60 B.n59 585
R1468 B.n960 B.n60 585
R1469 B.n958 B.n957 585
R1470 B.n959 B.n958 585
R1471 B.n956 B.n65 585
R1472 B.n65 B.n64 585
R1473 B.n955 B.n954 585
R1474 B.n954 B.n953 585
R1475 B.n67 B.n66 585
R1476 B.n952 B.n67 585
R1477 B.n950 B.n949 585
R1478 B.n951 B.n950 585
R1479 B.n948 B.n72 585
R1480 B.n72 B.n71 585
R1481 B.n947 B.n946 585
R1482 B.n946 B.n945 585
R1483 B.n74 B.n73 585
R1484 B.n944 B.n74 585
R1485 B.n942 B.n941 585
R1486 B.n943 B.n942 585
R1487 B.n940 B.n79 585
R1488 B.n79 B.n78 585
R1489 B.n939 B.n938 585
R1490 B.n938 B.n937 585
R1491 B.n81 B.n80 585
R1492 B.n936 B.n81 585
R1493 B.n934 B.n933 585
R1494 B.n935 B.n934 585
R1495 B.n932 B.n86 585
R1496 B.n86 B.n85 585
R1497 B.n931 B.n930 585
R1498 B.n930 B.n929 585
R1499 B.n88 B.n87 585
R1500 B.n928 B.n88 585
R1501 B.n926 B.n925 585
R1502 B.n927 B.n926 585
R1503 B.n924 B.n93 585
R1504 B.n93 B.n92 585
R1505 B.n923 B.n922 585
R1506 B.n922 B.n921 585
R1507 B.n95 B.n94 585
R1508 B.n920 B.n95 585
R1509 B.n918 B.n917 585
R1510 B.n919 B.n918 585
R1511 B.n916 B.n100 585
R1512 B.n100 B.n99 585
R1513 B.n915 B.n914 585
R1514 B.n914 B.n913 585
R1515 B.n102 B.n101 585
R1516 B.n912 B.n102 585
R1517 B.n1027 B.n1026 585
R1518 B.n1026 B.n1025 585
R1519 B.n659 B.n435 550.159
R1520 B.n153 B.n102 550.159
R1521 B.n662 B.n437 550.159
R1522 B.n909 B.n104 550.159
R1523 B.n487 B.t17 333.714
R1524 B.n149 B.t19 333.714
R1525 B.n484 B.t10 333.714
R1526 B.n151 B.t13 333.714
R1527 B.n487 B.t15 299.036
R1528 B.n484 B.t7 299.036
R1529 B.n151 B.t11 299.036
R1530 B.n149 B.t18 299.036
R1531 B.n488 B.t16 269.132
R1532 B.n150 B.t20 269.132
R1533 B.n485 B.t9 269.132
R1534 B.n152 B.t14 269.132
R1535 B.n911 B.n910 256.663
R1536 B.n911 B.n147 256.663
R1537 B.n911 B.n146 256.663
R1538 B.n911 B.n145 256.663
R1539 B.n911 B.n144 256.663
R1540 B.n911 B.n143 256.663
R1541 B.n911 B.n142 256.663
R1542 B.n911 B.n141 256.663
R1543 B.n911 B.n140 256.663
R1544 B.n911 B.n139 256.663
R1545 B.n911 B.n138 256.663
R1546 B.n911 B.n137 256.663
R1547 B.n911 B.n136 256.663
R1548 B.n911 B.n135 256.663
R1549 B.n911 B.n134 256.663
R1550 B.n911 B.n133 256.663
R1551 B.n911 B.n132 256.663
R1552 B.n911 B.n131 256.663
R1553 B.n911 B.n130 256.663
R1554 B.n911 B.n129 256.663
R1555 B.n911 B.n128 256.663
R1556 B.n911 B.n127 256.663
R1557 B.n911 B.n126 256.663
R1558 B.n911 B.n125 256.663
R1559 B.n911 B.n124 256.663
R1560 B.n911 B.n123 256.663
R1561 B.n911 B.n122 256.663
R1562 B.n911 B.n121 256.663
R1563 B.n911 B.n120 256.663
R1564 B.n911 B.n119 256.663
R1565 B.n911 B.n118 256.663
R1566 B.n911 B.n117 256.663
R1567 B.n911 B.n116 256.663
R1568 B.n911 B.n115 256.663
R1569 B.n911 B.n114 256.663
R1570 B.n911 B.n113 256.663
R1571 B.n911 B.n112 256.663
R1572 B.n911 B.n111 256.663
R1573 B.n911 B.n110 256.663
R1574 B.n911 B.n109 256.663
R1575 B.n911 B.n108 256.663
R1576 B.n911 B.n107 256.663
R1577 B.n911 B.n106 256.663
R1578 B.n911 B.n105 256.663
R1579 B.n661 B.n660 256.663
R1580 B.n661 B.n440 256.663
R1581 B.n661 B.n441 256.663
R1582 B.n661 B.n442 256.663
R1583 B.n661 B.n443 256.663
R1584 B.n661 B.n444 256.663
R1585 B.n661 B.n445 256.663
R1586 B.n661 B.n446 256.663
R1587 B.n661 B.n447 256.663
R1588 B.n661 B.n448 256.663
R1589 B.n661 B.n449 256.663
R1590 B.n661 B.n450 256.663
R1591 B.n661 B.n451 256.663
R1592 B.n661 B.n452 256.663
R1593 B.n661 B.n453 256.663
R1594 B.n661 B.n454 256.663
R1595 B.n661 B.n455 256.663
R1596 B.n661 B.n456 256.663
R1597 B.n661 B.n457 256.663
R1598 B.n661 B.n458 256.663
R1599 B.n661 B.n459 256.663
R1600 B.n661 B.n460 256.663
R1601 B.n661 B.n461 256.663
R1602 B.n661 B.n462 256.663
R1603 B.n661 B.n463 256.663
R1604 B.n661 B.n464 256.663
R1605 B.n661 B.n465 256.663
R1606 B.n661 B.n466 256.663
R1607 B.n661 B.n467 256.663
R1608 B.n661 B.n468 256.663
R1609 B.n661 B.n469 256.663
R1610 B.n661 B.n470 256.663
R1611 B.n661 B.n471 256.663
R1612 B.n661 B.n472 256.663
R1613 B.n661 B.n473 256.663
R1614 B.n661 B.n474 256.663
R1615 B.n661 B.n475 256.663
R1616 B.n661 B.n476 256.663
R1617 B.n661 B.n477 256.663
R1618 B.n661 B.n478 256.663
R1619 B.n661 B.n479 256.663
R1620 B.n661 B.n480 256.663
R1621 B.n661 B.n481 256.663
R1622 B.n668 B.n435 163.367
R1623 B.n668 B.n433 163.367
R1624 B.n672 B.n433 163.367
R1625 B.n672 B.n427 163.367
R1626 B.n680 B.n427 163.367
R1627 B.n680 B.n425 163.367
R1628 B.n684 B.n425 163.367
R1629 B.n684 B.n419 163.367
R1630 B.n692 B.n419 163.367
R1631 B.n692 B.n417 163.367
R1632 B.n696 B.n417 163.367
R1633 B.n696 B.n411 163.367
R1634 B.n704 B.n411 163.367
R1635 B.n704 B.n409 163.367
R1636 B.n708 B.n409 163.367
R1637 B.n708 B.n403 163.367
R1638 B.n716 B.n403 163.367
R1639 B.n716 B.n401 163.367
R1640 B.n720 B.n401 163.367
R1641 B.n720 B.n395 163.367
R1642 B.n728 B.n395 163.367
R1643 B.n728 B.n393 163.367
R1644 B.n732 B.n393 163.367
R1645 B.n732 B.n387 163.367
R1646 B.n740 B.n387 163.367
R1647 B.n740 B.n385 163.367
R1648 B.n744 B.n385 163.367
R1649 B.n744 B.n379 163.367
R1650 B.n753 B.n379 163.367
R1651 B.n753 B.n377 163.367
R1652 B.n757 B.n377 163.367
R1653 B.n757 B.n372 163.367
R1654 B.n765 B.n372 163.367
R1655 B.n765 B.n370 163.367
R1656 B.n769 B.n370 163.367
R1657 B.n769 B.n364 163.367
R1658 B.n777 B.n364 163.367
R1659 B.n777 B.n362 163.367
R1660 B.n781 B.n362 163.367
R1661 B.n781 B.n356 163.367
R1662 B.n789 B.n356 163.367
R1663 B.n789 B.n354 163.367
R1664 B.n793 B.n354 163.367
R1665 B.n793 B.n348 163.367
R1666 B.n801 B.n348 163.367
R1667 B.n801 B.n346 163.367
R1668 B.n805 B.n346 163.367
R1669 B.n805 B.n340 163.367
R1670 B.n814 B.n340 163.367
R1671 B.n814 B.n338 163.367
R1672 B.n818 B.n338 163.367
R1673 B.n818 B.n333 163.367
R1674 B.n827 B.n333 163.367
R1675 B.n827 B.n331 163.367
R1676 B.n831 B.n331 163.367
R1677 B.n831 B.n2 163.367
R1678 B.n1026 B.n2 163.367
R1679 B.n1026 B.n3 163.367
R1680 B.n1022 B.n3 163.367
R1681 B.n1022 B.n9 163.367
R1682 B.n1018 B.n9 163.367
R1683 B.n1018 B.n11 163.367
R1684 B.n1014 B.n11 163.367
R1685 B.n1014 B.n15 163.367
R1686 B.n1010 B.n15 163.367
R1687 B.n1010 B.n17 163.367
R1688 B.n1006 B.n17 163.367
R1689 B.n1006 B.n23 163.367
R1690 B.n1002 B.n23 163.367
R1691 B.n1002 B.n25 163.367
R1692 B.n998 B.n25 163.367
R1693 B.n998 B.n30 163.367
R1694 B.n994 B.n30 163.367
R1695 B.n994 B.n32 163.367
R1696 B.n990 B.n32 163.367
R1697 B.n990 B.n37 163.367
R1698 B.n986 B.n37 163.367
R1699 B.n986 B.n39 163.367
R1700 B.n982 B.n39 163.367
R1701 B.n982 B.n44 163.367
R1702 B.n978 B.n44 163.367
R1703 B.n978 B.n46 163.367
R1704 B.n974 B.n46 163.367
R1705 B.n974 B.n50 163.367
R1706 B.n970 B.n50 163.367
R1707 B.n970 B.n52 163.367
R1708 B.n966 B.n52 163.367
R1709 B.n966 B.n58 163.367
R1710 B.n962 B.n58 163.367
R1711 B.n962 B.n60 163.367
R1712 B.n958 B.n60 163.367
R1713 B.n958 B.n65 163.367
R1714 B.n954 B.n65 163.367
R1715 B.n954 B.n67 163.367
R1716 B.n950 B.n67 163.367
R1717 B.n950 B.n72 163.367
R1718 B.n946 B.n72 163.367
R1719 B.n946 B.n74 163.367
R1720 B.n942 B.n74 163.367
R1721 B.n942 B.n79 163.367
R1722 B.n938 B.n79 163.367
R1723 B.n938 B.n81 163.367
R1724 B.n934 B.n81 163.367
R1725 B.n934 B.n86 163.367
R1726 B.n930 B.n86 163.367
R1727 B.n930 B.n88 163.367
R1728 B.n926 B.n88 163.367
R1729 B.n926 B.n93 163.367
R1730 B.n922 B.n93 163.367
R1731 B.n922 B.n95 163.367
R1732 B.n918 B.n95 163.367
R1733 B.n918 B.n100 163.367
R1734 B.n914 B.n100 163.367
R1735 B.n914 B.n102 163.367
R1736 B.n483 B.n482 163.367
R1737 B.n654 B.n482 163.367
R1738 B.n652 B.n651 163.367
R1739 B.n648 B.n647 163.367
R1740 B.n644 B.n643 163.367
R1741 B.n640 B.n639 163.367
R1742 B.n636 B.n635 163.367
R1743 B.n632 B.n631 163.367
R1744 B.n628 B.n627 163.367
R1745 B.n624 B.n623 163.367
R1746 B.n620 B.n619 163.367
R1747 B.n616 B.n615 163.367
R1748 B.n612 B.n611 163.367
R1749 B.n608 B.n607 163.367
R1750 B.n604 B.n603 163.367
R1751 B.n600 B.n599 163.367
R1752 B.n596 B.n595 163.367
R1753 B.n592 B.n591 163.367
R1754 B.n588 B.n587 163.367
R1755 B.n584 B.n583 163.367
R1756 B.n580 B.n579 163.367
R1757 B.n576 B.n575 163.367
R1758 B.n572 B.n571 163.367
R1759 B.n568 B.n567 163.367
R1760 B.n564 B.n563 163.367
R1761 B.n560 B.n559 163.367
R1762 B.n556 B.n555 163.367
R1763 B.n552 B.n551 163.367
R1764 B.n548 B.n547 163.367
R1765 B.n544 B.n543 163.367
R1766 B.n540 B.n539 163.367
R1767 B.n536 B.n535 163.367
R1768 B.n532 B.n531 163.367
R1769 B.n528 B.n527 163.367
R1770 B.n524 B.n523 163.367
R1771 B.n520 B.n519 163.367
R1772 B.n516 B.n515 163.367
R1773 B.n512 B.n511 163.367
R1774 B.n508 B.n507 163.367
R1775 B.n504 B.n503 163.367
R1776 B.n500 B.n499 163.367
R1777 B.n496 B.n495 163.367
R1778 B.n492 B.n491 163.367
R1779 B.n662 B.n439 163.367
R1780 B.n666 B.n437 163.367
R1781 B.n666 B.n431 163.367
R1782 B.n674 B.n431 163.367
R1783 B.n674 B.n429 163.367
R1784 B.n678 B.n429 163.367
R1785 B.n678 B.n422 163.367
R1786 B.n686 B.n422 163.367
R1787 B.n686 B.n420 163.367
R1788 B.n690 B.n420 163.367
R1789 B.n690 B.n415 163.367
R1790 B.n698 B.n415 163.367
R1791 B.n698 B.n413 163.367
R1792 B.n702 B.n413 163.367
R1793 B.n702 B.n407 163.367
R1794 B.n710 B.n407 163.367
R1795 B.n710 B.n405 163.367
R1796 B.n714 B.n405 163.367
R1797 B.n714 B.n399 163.367
R1798 B.n722 B.n399 163.367
R1799 B.n722 B.n397 163.367
R1800 B.n726 B.n397 163.367
R1801 B.n726 B.n391 163.367
R1802 B.n734 B.n391 163.367
R1803 B.n734 B.n389 163.367
R1804 B.n738 B.n389 163.367
R1805 B.n738 B.n383 163.367
R1806 B.n746 B.n383 163.367
R1807 B.n746 B.n381 163.367
R1808 B.n750 B.n381 163.367
R1809 B.n750 B.n376 163.367
R1810 B.n759 B.n376 163.367
R1811 B.n759 B.n374 163.367
R1812 B.n763 B.n374 163.367
R1813 B.n763 B.n368 163.367
R1814 B.n771 B.n368 163.367
R1815 B.n771 B.n366 163.367
R1816 B.n775 B.n366 163.367
R1817 B.n775 B.n359 163.367
R1818 B.n783 B.n359 163.367
R1819 B.n783 B.n357 163.367
R1820 B.n787 B.n357 163.367
R1821 B.n787 B.n352 163.367
R1822 B.n795 B.n352 163.367
R1823 B.n795 B.n350 163.367
R1824 B.n799 B.n350 163.367
R1825 B.n799 B.n344 163.367
R1826 B.n807 B.n344 163.367
R1827 B.n807 B.n342 163.367
R1828 B.n811 B.n342 163.367
R1829 B.n811 B.n337 163.367
R1830 B.n820 B.n337 163.367
R1831 B.n820 B.n335 163.367
R1832 B.n825 B.n335 163.367
R1833 B.n825 B.n329 163.367
R1834 B.n833 B.n329 163.367
R1835 B.n834 B.n833 163.367
R1836 B.n834 B.n5 163.367
R1837 B.n6 B.n5 163.367
R1838 B.n7 B.n6 163.367
R1839 B.n839 B.n7 163.367
R1840 B.n839 B.n12 163.367
R1841 B.n13 B.n12 163.367
R1842 B.n14 B.n13 163.367
R1843 B.n844 B.n14 163.367
R1844 B.n844 B.n19 163.367
R1845 B.n20 B.n19 163.367
R1846 B.n21 B.n20 163.367
R1847 B.n849 B.n21 163.367
R1848 B.n849 B.n26 163.367
R1849 B.n27 B.n26 163.367
R1850 B.n28 B.n27 163.367
R1851 B.n854 B.n28 163.367
R1852 B.n854 B.n33 163.367
R1853 B.n34 B.n33 163.367
R1854 B.n35 B.n34 163.367
R1855 B.n859 B.n35 163.367
R1856 B.n859 B.n40 163.367
R1857 B.n41 B.n40 163.367
R1858 B.n42 B.n41 163.367
R1859 B.n864 B.n42 163.367
R1860 B.n864 B.n47 163.367
R1861 B.n48 B.n47 163.367
R1862 B.n49 B.n48 163.367
R1863 B.n869 B.n49 163.367
R1864 B.n869 B.n54 163.367
R1865 B.n55 B.n54 163.367
R1866 B.n56 B.n55 163.367
R1867 B.n874 B.n56 163.367
R1868 B.n874 B.n61 163.367
R1869 B.n62 B.n61 163.367
R1870 B.n63 B.n62 163.367
R1871 B.n879 B.n63 163.367
R1872 B.n879 B.n68 163.367
R1873 B.n69 B.n68 163.367
R1874 B.n70 B.n69 163.367
R1875 B.n884 B.n70 163.367
R1876 B.n884 B.n75 163.367
R1877 B.n76 B.n75 163.367
R1878 B.n77 B.n76 163.367
R1879 B.n889 B.n77 163.367
R1880 B.n889 B.n82 163.367
R1881 B.n83 B.n82 163.367
R1882 B.n84 B.n83 163.367
R1883 B.n894 B.n84 163.367
R1884 B.n894 B.n89 163.367
R1885 B.n90 B.n89 163.367
R1886 B.n91 B.n90 163.367
R1887 B.n899 B.n91 163.367
R1888 B.n899 B.n96 163.367
R1889 B.n97 B.n96 163.367
R1890 B.n98 B.n97 163.367
R1891 B.n904 B.n98 163.367
R1892 B.n904 B.n103 163.367
R1893 B.n104 B.n103 163.367
R1894 B.n157 B.n156 163.367
R1895 B.n161 B.n160 163.367
R1896 B.n165 B.n164 163.367
R1897 B.n169 B.n168 163.367
R1898 B.n173 B.n172 163.367
R1899 B.n177 B.n176 163.367
R1900 B.n181 B.n180 163.367
R1901 B.n185 B.n184 163.367
R1902 B.n189 B.n188 163.367
R1903 B.n193 B.n192 163.367
R1904 B.n197 B.n196 163.367
R1905 B.n201 B.n200 163.367
R1906 B.n205 B.n204 163.367
R1907 B.n209 B.n208 163.367
R1908 B.n213 B.n212 163.367
R1909 B.n217 B.n216 163.367
R1910 B.n221 B.n220 163.367
R1911 B.n225 B.n224 163.367
R1912 B.n229 B.n228 163.367
R1913 B.n234 B.n233 163.367
R1914 B.n238 B.n237 163.367
R1915 B.n242 B.n241 163.367
R1916 B.n246 B.n245 163.367
R1917 B.n250 B.n249 163.367
R1918 B.n255 B.n254 163.367
R1919 B.n259 B.n258 163.367
R1920 B.n263 B.n262 163.367
R1921 B.n267 B.n266 163.367
R1922 B.n271 B.n270 163.367
R1923 B.n275 B.n274 163.367
R1924 B.n279 B.n278 163.367
R1925 B.n283 B.n282 163.367
R1926 B.n287 B.n286 163.367
R1927 B.n291 B.n290 163.367
R1928 B.n295 B.n294 163.367
R1929 B.n299 B.n298 163.367
R1930 B.n303 B.n302 163.367
R1931 B.n307 B.n306 163.367
R1932 B.n311 B.n310 163.367
R1933 B.n315 B.n314 163.367
R1934 B.n319 B.n318 163.367
R1935 B.n323 B.n322 163.367
R1936 B.n325 B.n148 163.367
R1937 B.n661 B.n436 85.8185
R1938 B.n912 B.n911 85.8185
R1939 B.n660 B.n659 71.676
R1940 B.n654 B.n440 71.676
R1941 B.n651 B.n441 71.676
R1942 B.n647 B.n442 71.676
R1943 B.n643 B.n443 71.676
R1944 B.n639 B.n444 71.676
R1945 B.n635 B.n445 71.676
R1946 B.n631 B.n446 71.676
R1947 B.n627 B.n447 71.676
R1948 B.n623 B.n448 71.676
R1949 B.n619 B.n449 71.676
R1950 B.n615 B.n450 71.676
R1951 B.n611 B.n451 71.676
R1952 B.n607 B.n452 71.676
R1953 B.n603 B.n453 71.676
R1954 B.n599 B.n454 71.676
R1955 B.n595 B.n455 71.676
R1956 B.n591 B.n456 71.676
R1957 B.n587 B.n457 71.676
R1958 B.n583 B.n458 71.676
R1959 B.n579 B.n459 71.676
R1960 B.n575 B.n460 71.676
R1961 B.n571 B.n461 71.676
R1962 B.n567 B.n462 71.676
R1963 B.n563 B.n463 71.676
R1964 B.n559 B.n464 71.676
R1965 B.n555 B.n465 71.676
R1966 B.n551 B.n466 71.676
R1967 B.n547 B.n467 71.676
R1968 B.n543 B.n468 71.676
R1969 B.n539 B.n469 71.676
R1970 B.n535 B.n470 71.676
R1971 B.n531 B.n471 71.676
R1972 B.n527 B.n472 71.676
R1973 B.n523 B.n473 71.676
R1974 B.n519 B.n474 71.676
R1975 B.n515 B.n475 71.676
R1976 B.n511 B.n476 71.676
R1977 B.n507 B.n477 71.676
R1978 B.n503 B.n478 71.676
R1979 B.n499 B.n479 71.676
R1980 B.n495 B.n480 71.676
R1981 B.n491 B.n481 71.676
R1982 B.n153 B.n105 71.676
R1983 B.n157 B.n106 71.676
R1984 B.n161 B.n107 71.676
R1985 B.n165 B.n108 71.676
R1986 B.n169 B.n109 71.676
R1987 B.n173 B.n110 71.676
R1988 B.n177 B.n111 71.676
R1989 B.n181 B.n112 71.676
R1990 B.n185 B.n113 71.676
R1991 B.n189 B.n114 71.676
R1992 B.n193 B.n115 71.676
R1993 B.n197 B.n116 71.676
R1994 B.n201 B.n117 71.676
R1995 B.n205 B.n118 71.676
R1996 B.n209 B.n119 71.676
R1997 B.n213 B.n120 71.676
R1998 B.n217 B.n121 71.676
R1999 B.n221 B.n122 71.676
R2000 B.n225 B.n123 71.676
R2001 B.n229 B.n124 71.676
R2002 B.n234 B.n125 71.676
R2003 B.n238 B.n126 71.676
R2004 B.n242 B.n127 71.676
R2005 B.n246 B.n128 71.676
R2006 B.n250 B.n129 71.676
R2007 B.n255 B.n130 71.676
R2008 B.n259 B.n131 71.676
R2009 B.n263 B.n132 71.676
R2010 B.n267 B.n133 71.676
R2011 B.n271 B.n134 71.676
R2012 B.n275 B.n135 71.676
R2013 B.n279 B.n136 71.676
R2014 B.n283 B.n137 71.676
R2015 B.n287 B.n138 71.676
R2016 B.n291 B.n139 71.676
R2017 B.n295 B.n140 71.676
R2018 B.n299 B.n141 71.676
R2019 B.n303 B.n142 71.676
R2020 B.n307 B.n143 71.676
R2021 B.n311 B.n144 71.676
R2022 B.n315 B.n145 71.676
R2023 B.n319 B.n146 71.676
R2024 B.n323 B.n147 71.676
R2025 B.n910 B.n148 71.676
R2026 B.n910 B.n909 71.676
R2027 B.n325 B.n147 71.676
R2028 B.n322 B.n146 71.676
R2029 B.n318 B.n145 71.676
R2030 B.n314 B.n144 71.676
R2031 B.n310 B.n143 71.676
R2032 B.n306 B.n142 71.676
R2033 B.n302 B.n141 71.676
R2034 B.n298 B.n140 71.676
R2035 B.n294 B.n139 71.676
R2036 B.n290 B.n138 71.676
R2037 B.n286 B.n137 71.676
R2038 B.n282 B.n136 71.676
R2039 B.n278 B.n135 71.676
R2040 B.n274 B.n134 71.676
R2041 B.n270 B.n133 71.676
R2042 B.n266 B.n132 71.676
R2043 B.n262 B.n131 71.676
R2044 B.n258 B.n130 71.676
R2045 B.n254 B.n129 71.676
R2046 B.n249 B.n128 71.676
R2047 B.n245 B.n127 71.676
R2048 B.n241 B.n126 71.676
R2049 B.n237 B.n125 71.676
R2050 B.n233 B.n124 71.676
R2051 B.n228 B.n123 71.676
R2052 B.n224 B.n122 71.676
R2053 B.n220 B.n121 71.676
R2054 B.n216 B.n120 71.676
R2055 B.n212 B.n119 71.676
R2056 B.n208 B.n118 71.676
R2057 B.n204 B.n117 71.676
R2058 B.n200 B.n116 71.676
R2059 B.n196 B.n115 71.676
R2060 B.n192 B.n114 71.676
R2061 B.n188 B.n113 71.676
R2062 B.n184 B.n112 71.676
R2063 B.n180 B.n111 71.676
R2064 B.n176 B.n110 71.676
R2065 B.n172 B.n109 71.676
R2066 B.n168 B.n108 71.676
R2067 B.n164 B.n107 71.676
R2068 B.n160 B.n106 71.676
R2069 B.n156 B.n105 71.676
R2070 B.n660 B.n483 71.676
R2071 B.n652 B.n440 71.676
R2072 B.n648 B.n441 71.676
R2073 B.n644 B.n442 71.676
R2074 B.n640 B.n443 71.676
R2075 B.n636 B.n444 71.676
R2076 B.n632 B.n445 71.676
R2077 B.n628 B.n446 71.676
R2078 B.n624 B.n447 71.676
R2079 B.n620 B.n448 71.676
R2080 B.n616 B.n449 71.676
R2081 B.n612 B.n450 71.676
R2082 B.n608 B.n451 71.676
R2083 B.n604 B.n452 71.676
R2084 B.n600 B.n453 71.676
R2085 B.n596 B.n454 71.676
R2086 B.n592 B.n455 71.676
R2087 B.n588 B.n456 71.676
R2088 B.n584 B.n457 71.676
R2089 B.n580 B.n458 71.676
R2090 B.n576 B.n459 71.676
R2091 B.n572 B.n460 71.676
R2092 B.n568 B.n461 71.676
R2093 B.n564 B.n462 71.676
R2094 B.n560 B.n463 71.676
R2095 B.n556 B.n464 71.676
R2096 B.n552 B.n465 71.676
R2097 B.n548 B.n466 71.676
R2098 B.n544 B.n467 71.676
R2099 B.n540 B.n468 71.676
R2100 B.n536 B.n469 71.676
R2101 B.n532 B.n470 71.676
R2102 B.n528 B.n471 71.676
R2103 B.n524 B.n472 71.676
R2104 B.n520 B.n473 71.676
R2105 B.n516 B.n474 71.676
R2106 B.n512 B.n475 71.676
R2107 B.n508 B.n476 71.676
R2108 B.n504 B.n477 71.676
R2109 B.n500 B.n478 71.676
R2110 B.n496 B.n479 71.676
R2111 B.n492 B.n480 71.676
R2112 B.n481 B.n439 71.676
R2113 B.n488 B.n487 64.5823
R2114 B.n485 B.n484 64.5823
R2115 B.n152 B.n151 64.5823
R2116 B.n150 B.n149 64.5823
R2117 B.n489 B.n488 59.5399
R2118 B.n486 B.n485 59.5399
R2119 B.n231 B.n152 59.5399
R2120 B.n252 B.n150 59.5399
R2121 B.n667 B.n436 45.2379
R2122 B.n667 B.n432 45.2379
R2123 B.n673 B.n432 45.2379
R2124 B.n673 B.n428 45.2379
R2125 B.n679 B.n428 45.2379
R2126 B.n679 B.n423 45.2379
R2127 B.n685 B.n423 45.2379
R2128 B.n685 B.n424 45.2379
R2129 B.n691 B.n416 45.2379
R2130 B.n697 B.n416 45.2379
R2131 B.n697 B.n412 45.2379
R2132 B.n703 B.n412 45.2379
R2133 B.n703 B.n408 45.2379
R2134 B.n709 B.n408 45.2379
R2135 B.n709 B.n404 45.2379
R2136 B.n715 B.n404 45.2379
R2137 B.n715 B.n400 45.2379
R2138 B.n721 B.n400 45.2379
R2139 B.n721 B.n396 45.2379
R2140 B.n727 B.n396 45.2379
R2141 B.n733 B.n392 45.2379
R2142 B.n733 B.n388 45.2379
R2143 B.n739 B.n388 45.2379
R2144 B.n739 B.n384 45.2379
R2145 B.n745 B.n384 45.2379
R2146 B.n745 B.n380 45.2379
R2147 B.n752 B.n380 45.2379
R2148 B.n752 B.n751 45.2379
R2149 B.n758 B.n373 45.2379
R2150 B.n764 B.n373 45.2379
R2151 B.n764 B.n369 45.2379
R2152 B.n770 B.n369 45.2379
R2153 B.n770 B.n365 45.2379
R2154 B.n776 B.n365 45.2379
R2155 B.n776 B.n360 45.2379
R2156 B.n782 B.n360 45.2379
R2157 B.n782 B.n361 45.2379
R2158 B.n788 B.n353 45.2379
R2159 B.n794 B.n353 45.2379
R2160 B.n794 B.n349 45.2379
R2161 B.n800 B.n349 45.2379
R2162 B.n800 B.n345 45.2379
R2163 B.n806 B.n345 45.2379
R2164 B.n806 B.n341 45.2379
R2165 B.n813 B.n341 45.2379
R2166 B.n813 B.n812 45.2379
R2167 B.n819 B.n334 45.2379
R2168 B.n826 B.n334 45.2379
R2169 B.n826 B.n330 45.2379
R2170 B.n832 B.n330 45.2379
R2171 B.n832 B.n4 45.2379
R2172 B.n1025 B.n4 45.2379
R2173 B.n1025 B.n1024 45.2379
R2174 B.n1024 B.n1023 45.2379
R2175 B.n1023 B.n8 45.2379
R2176 B.n1017 B.n8 45.2379
R2177 B.n1017 B.n1016 45.2379
R2178 B.n1016 B.n1015 45.2379
R2179 B.n1009 B.n18 45.2379
R2180 B.n1009 B.n1008 45.2379
R2181 B.n1008 B.n1007 45.2379
R2182 B.n1007 B.n22 45.2379
R2183 B.n1001 B.n22 45.2379
R2184 B.n1001 B.n1000 45.2379
R2185 B.n1000 B.n999 45.2379
R2186 B.n999 B.n29 45.2379
R2187 B.n993 B.n29 45.2379
R2188 B.n992 B.n991 45.2379
R2189 B.n991 B.n36 45.2379
R2190 B.n985 B.n36 45.2379
R2191 B.n985 B.n984 45.2379
R2192 B.n984 B.n983 45.2379
R2193 B.n983 B.n43 45.2379
R2194 B.n977 B.n43 45.2379
R2195 B.n977 B.n976 45.2379
R2196 B.n976 B.n975 45.2379
R2197 B.n969 B.n53 45.2379
R2198 B.n969 B.n968 45.2379
R2199 B.n968 B.n967 45.2379
R2200 B.n967 B.n57 45.2379
R2201 B.n961 B.n57 45.2379
R2202 B.n961 B.n960 45.2379
R2203 B.n960 B.n959 45.2379
R2204 B.n959 B.n64 45.2379
R2205 B.n953 B.n952 45.2379
R2206 B.n952 B.n951 45.2379
R2207 B.n951 B.n71 45.2379
R2208 B.n945 B.n71 45.2379
R2209 B.n945 B.n944 45.2379
R2210 B.n944 B.n943 45.2379
R2211 B.n943 B.n78 45.2379
R2212 B.n937 B.n78 45.2379
R2213 B.n937 B.n936 45.2379
R2214 B.n936 B.n935 45.2379
R2215 B.n935 B.n85 45.2379
R2216 B.n929 B.n85 45.2379
R2217 B.n928 B.n927 45.2379
R2218 B.n927 B.n92 45.2379
R2219 B.n921 B.n92 45.2379
R2220 B.n921 B.n920 45.2379
R2221 B.n920 B.n919 45.2379
R2222 B.n919 B.n99 45.2379
R2223 B.n913 B.n99 45.2379
R2224 B.n913 B.n912 45.2379
R2225 B.n751 B.t5 41.2463
R2226 B.n53 B.t3 41.2463
R2227 B.n691 B.t8 39.9158
R2228 B.t21 B.n392 39.9158
R2229 B.t1 B.n64 39.9158
R2230 B.n929 B.t12 39.9158
R2231 B.n154 B.n101 35.7468
R2232 B.n664 B.n663 35.7468
R2233 B.n658 B.n434 35.7468
R2234 B.n908 B.n907 35.7468
R2235 B.n361 B.t0 31.9328
R2236 B.t2 B.n992 31.9328
R2237 B.n812 B.t6 22.6192
R2238 B.n819 B.t6 22.6192
R2239 B.n1015 B.t4 22.6192
R2240 B.n18 B.t4 22.6192
R2241 B B.n1027 18.0485
R2242 B.n788 B.t0 13.3056
R2243 B.n993 B.t2 13.3056
R2244 B.n155 B.n154 10.6151
R2245 B.n158 B.n155 10.6151
R2246 B.n159 B.n158 10.6151
R2247 B.n162 B.n159 10.6151
R2248 B.n163 B.n162 10.6151
R2249 B.n166 B.n163 10.6151
R2250 B.n167 B.n166 10.6151
R2251 B.n170 B.n167 10.6151
R2252 B.n171 B.n170 10.6151
R2253 B.n174 B.n171 10.6151
R2254 B.n175 B.n174 10.6151
R2255 B.n178 B.n175 10.6151
R2256 B.n179 B.n178 10.6151
R2257 B.n182 B.n179 10.6151
R2258 B.n183 B.n182 10.6151
R2259 B.n186 B.n183 10.6151
R2260 B.n187 B.n186 10.6151
R2261 B.n190 B.n187 10.6151
R2262 B.n191 B.n190 10.6151
R2263 B.n194 B.n191 10.6151
R2264 B.n195 B.n194 10.6151
R2265 B.n198 B.n195 10.6151
R2266 B.n199 B.n198 10.6151
R2267 B.n202 B.n199 10.6151
R2268 B.n203 B.n202 10.6151
R2269 B.n206 B.n203 10.6151
R2270 B.n207 B.n206 10.6151
R2271 B.n210 B.n207 10.6151
R2272 B.n211 B.n210 10.6151
R2273 B.n214 B.n211 10.6151
R2274 B.n215 B.n214 10.6151
R2275 B.n218 B.n215 10.6151
R2276 B.n219 B.n218 10.6151
R2277 B.n222 B.n219 10.6151
R2278 B.n223 B.n222 10.6151
R2279 B.n226 B.n223 10.6151
R2280 B.n227 B.n226 10.6151
R2281 B.n230 B.n227 10.6151
R2282 B.n235 B.n232 10.6151
R2283 B.n236 B.n235 10.6151
R2284 B.n239 B.n236 10.6151
R2285 B.n240 B.n239 10.6151
R2286 B.n243 B.n240 10.6151
R2287 B.n244 B.n243 10.6151
R2288 B.n247 B.n244 10.6151
R2289 B.n248 B.n247 10.6151
R2290 B.n251 B.n248 10.6151
R2291 B.n256 B.n253 10.6151
R2292 B.n257 B.n256 10.6151
R2293 B.n260 B.n257 10.6151
R2294 B.n261 B.n260 10.6151
R2295 B.n264 B.n261 10.6151
R2296 B.n265 B.n264 10.6151
R2297 B.n268 B.n265 10.6151
R2298 B.n269 B.n268 10.6151
R2299 B.n272 B.n269 10.6151
R2300 B.n273 B.n272 10.6151
R2301 B.n276 B.n273 10.6151
R2302 B.n277 B.n276 10.6151
R2303 B.n280 B.n277 10.6151
R2304 B.n281 B.n280 10.6151
R2305 B.n284 B.n281 10.6151
R2306 B.n285 B.n284 10.6151
R2307 B.n288 B.n285 10.6151
R2308 B.n289 B.n288 10.6151
R2309 B.n292 B.n289 10.6151
R2310 B.n293 B.n292 10.6151
R2311 B.n296 B.n293 10.6151
R2312 B.n297 B.n296 10.6151
R2313 B.n300 B.n297 10.6151
R2314 B.n301 B.n300 10.6151
R2315 B.n304 B.n301 10.6151
R2316 B.n305 B.n304 10.6151
R2317 B.n308 B.n305 10.6151
R2318 B.n309 B.n308 10.6151
R2319 B.n312 B.n309 10.6151
R2320 B.n313 B.n312 10.6151
R2321 B.n316 B.n313 10.6151
R2322 B.n317 B.n316 10.6151
R2323 B.n320 B.n317 10.6151
R2324 B.n321 B.n320 10.6151
R2325 B.n324 B.n321 10.6151
R2326 B.n326 B.n324 10.6151
R2327 B.n327 B.n326 10.6151
R2328 B.n908 B.n327 10.6151
R2329 B.n665 B.n664 10.6151
R2330 B.n665 B.n430 10.6151
R2331 B.n675 B.n430 10.6151
R2332 B.n676 B.n675 10.6151
R2333 B.n677 B.n676 10.6151
R2334 B.n677 B.n421 10.6151
R2335 B.n687 B.n421 10.6151
R2336 B.n688 B.n687 10.6151
R2337 B.n689 B.n688 10.6151
R2338 B.n689 B.n414 10.6151
R2339 B.n699 B.n414 10.6151
R2340 B.n700 B.n699 10.6151
R2341 B.n701 B.n700 10.6151
R2342 B.n701 B.n406 10.6151
R2343 B.n711 B.n406 10.6151
R2344 B.n712 B.n711 10.6151
R2345 B.n713 B.n712 10.6151
R2346 B.n713 B.n398 10.6151
R2347 B.n723 B.n398 10.6151
R2348 B.n724 B.n723 10.6151
R2349 B.n725 B.n724 10.6151
R2350 B.n725 B.n390 10.6151
R2351 B.n735 B.n390 10.6151
R2352 B.n736 B.n735 10.6151
R2353 B.n737 B.n736 10.6151
R2354 B.n737 B.n382 10.6151
R2355 B.n747 B.n382 10.6151
R2356 B.n748 B.n747 10.6151
R2357 B.n749 B.n748 10.6151
R2358 B.n749 B.n375 10.6151
R2359 B.n760 B.n375 10.6151
R2360 B.n761 B.n760 10.6151
R2361 B.n762 B.n761 10.6151
R2362 B.n762 B.n367 10.6151
R2363 B.n772 B.n367 10.6151
R2364 B.n773 B.n772 10.6151
R2365 B.n774 B.n773 10.6151
R2366 B.n774 B.n358 10.6151
R2367 B.n784 B.n358 10.6151
R2368 B.n785 B.n784 10.6151
R2369 B.n786 B.n785 10.6151
R2370 B.n786 B.n351 10.6151
R2371 B.n796 B.n351 10.6151
R2372 B.n797 B.n796 10.6151
R2373 B.n798 B.n797 10.6151
R2374 B.n798 B.n343 10.6151
R2375 B.n808 B.n343 10.6151
R2376 B.n809 B.n808 10.6151
R2377 B.n810 B.n809 10.6151
R2378 B.n810 B.n336 10.6151
R2379 B.n821 B.n336 10.6151
R2380 B.n822 B.n821 10.6151
R2381 B.n824 B.n822 10.6151
R2382 B.n824 B.n823 10.6151
R2383 B.n823 B.n328 10.6151
R2384 B.n835 B.n328 10.6151
R2385 B.n836 B.n835 10.6151
R2386 B.n837 B.n836 10.6151
R2387 B.n838 B.n837 10.6151
R2388 B.n840 B.n838 10.6151
R2389 B.n841 B.n840 10.6151
R2390 B.n842 B.n841 10.6151
R2391 B.n843 B.n842 10.6151
R2392 B.n845 B.n843 10.6151
R2393 B.n846 B.n845 10.6151
R2394 B.n847 B.n846 10.6151
R2395 B.n848 B.n847 10.6151
R2396 B.n850 B.n848 10.6151
R2397 B.n851 B.n850 10.6151
R2398 B.n852 B.n851 10.6151
R2399 B.n853 B.n852 10.6151
R2400 B.n855 B.n853 10.6151
R2401 B.n856 B.n855 10.6151
R2402 B.n857 B.n856 10.6151
R2403 B.n858 B.n857 10.6151
R2404 B.n860 B.n858 10.6151
R2405 B.n861 B.n860 10.6151
R2406 B.n862 B.n861 10.6151
R2407 B.n863 B.n862 10.6151
R2408 B.n865 B.n863 10.6151
R2409 B.n866 B.n865 10.6151
R2410 B.n867 B.n866 10.6151
R2411 B.n868 B.n867 10.6151
R2412 B.n870 B.n868 10.6151
R2413 B.n871 B.n870 10.6151
R2414 B.n872 B.n871 10.6151
R2415 B.n873 B.n872 10.6151
R2416 B.n875 B.n873 10.6151
R2417 B.n876 B.n875 10.6151
R2418 B.n877 B.n876 10.6151
R2419 B.n878 B.n877 10.6151
R2420 B.n880 B.n878 10.6151
R2421 B.n881 B.n880 10.6151
R2422 B.n882 B.n881 10.6151
R2423 B.n883 B.n882 10.6151
R2424 B.n885 B.n883 10.6151
R2425 B.n886 B.n885 10.6151
R2426 B.n887 B.n886 10.6151
R2427 B.n888 B.n887 10.6151
R2428 B.n890 B.n888 10.6151
R2429 B.n891 B.n890 10.6151
R2430 B.n892 B.n891 10.6151
R2431 B.n893 B.n892 10.6151
R2432 B.n895 B.n893 10.6151
R2433 B.n896 B.n895 10.6151
R2434 B.n897 B.n896 10.6151
R2435 B.n898 B.n897 10.6151
R2436 B.n900 B.n898 10.6151
R2437 B.n901 B.n900 10.6151
R2438 B.n902 B.n901 10.6151
R2439 B.n903 B.n902 10.6151
R2440 B.n905 B.n903 10.6151
R2441 B.n906 B.n905 10.6151
R2442 B.n907 B.n906 10.6151
R2443 B.n658 B.n657 10.6151
R2444 B.n657 B.n656 10.6151
R2445 B.n656 B.n655 10.6151
R2446 B.n655 B.n653 10.6151
R2447 B.n653 B.n650 10.6151
R2448 B.n650 B.n649 10.6151
R2449 B.n649 B.n646 10.6151
R2450 B.n646 B.n645 10.6151
R2451 B.n645 B.n642 10.6151
R2452 B.n642 B.n641 10.6151
R2453 B.n641 B.n638 10.6151
R2454 B.n638 B.n637 10.6151
R2455 B.n637 B.n634 10.6151
R2456 B.n634 B.n633 10.6151
R2457 B.n633 B.n630 10.6151
R2458 B.n630 B.n629 10.6151
R2459 B.n629 B.n626 10.6151
R2460 B.n626 B.n625 10.6151
R2461 B.n625 B.n622 10.6151
R2462 B.n622 B.n621 10.6151
R2463 B.n621 B.n618 10.6151
R2464 B.n618 B.n617 10.6151
R2465 B.n617 B.n614 10.6151
R2466 B.n614 B.n613 10.6151
R2467 B.n613 B.n610 10.6151
R2468 B.n610 B.n609 10.6151
R2469 B.n609 B.n606 10.6151
R2470 B.n606 B.n605 10.6151
R2471 B.n605 B.n602 10.6151
R2472 B.n602 B.n601 10.6151
R2473 B.n601 B.n598 10.6151
R2474 B.n598 B.n597 10.6151
R2475 B.n597 B.n594 10.6151
R2476 B.n594 B.n593 10.6151
R2477 B.n593 B.n590 10.6151
R2478 B.n590 B.n589 10.6151
R2479 B.n589 B.n586 10.6151
R2480 B.n586 B.n585 10.6151
R2481 B.n582 B.n581 10.6151
R2482 B.n581 B.n578 10.6151
R2483 B.n578 B.n577 10.6151
R2484 B.n577 B.n574 10.6151
R2485 B.n574 B.n573 10.6151
R2486 B.n573 B.n570 10.6151
R2487 B.n570 B.n569 10.6151
R2488 B.n569 B.n566 10.6151
R2489 B.n566 B.n565 10.6151
R2490 B.n562 B.n561 10.6151
R2491 B.n561 B.n558 10.6151
R2492 B.n558 B.n557 10.6151
R2493 B.n557 B.n554 10.6151
R2494 B.n554 B.n553 10.6151
R2495 B.n553 B.n550 10.6151
R2496 B.n550 B.n549 10.6151
R2497 B.n549 B.n546 10.6151
R2498 B.n546 B.n545 10.6151
R2499 B.n545 B.n542 10.6151
R2500 B.n542 B.n541 10.6151
R2501 B.n541 B.n538 10.6151
R2502 B.n538 B.n537 10.6151
R2503 B.n537 B.n534 10.6151
R2504 B.n534 B.n533 10.6151
R2505 B.n533 B.n530 10.6151
R2506 B.n530 B.n529 10.6151
R2507 B.n529 B.n526 10.6151
R2508 B.n526 B.n525 10.6151
R2509 B.n525 B.n522 10.6151
R2510 B.n522 B.n521 10.6151
R2511 B.n521 B.n518 10.6151
R2512 B.n518 B.n517 10.6151
R2513 B.n517 B.n514 10.6151
R2514 B.n514 B.n513 10.6151
R2515 B.n513 B.n510 10.6151
R2516 B.n510 B.n509 10.6151
R2517 B.n509 B.n506 10.6151
R2518 B.n506 B.n505 10.6151
R2519 B.n505 B.n502 10.6151
R2520 B.n502 B.n501 10.6151
R2521 B.n501 B.n498 10.6151
R2522 B.n498 B.n497 10.6151
R2523 B.n497 B.n494 10.6151
R2524 B.n494 B.n493 10.6151
R2525 B.n493 B.n490 10.6151
R2526 B.n490 B.n438 10.6151
R2527 B.n663 B.n438 10.6151
R2528 B.n669 B.n434 10.6151
R2529 B.n670 B.n669 10.6151
R2530 B.n671 B.n670 10.6151
R2531 B.n671 B.n426 10.6151
R2532 B.n681 B.n426 10.6151
R2533 B.n682 B.n681 10.6151
R2534 B.n683 B.n682 10.6151
R2535 B.n683 B.n418 10.6151
R2536 B.n693 B.n418 10.6151
R2537 B.n694 B.n693 10.6151
R2538 B.n695 B.n694 10.6151
R2539 B.n695 B.n410 10.6151
R2540 B.n705 B.n410 10.6151
R2541 B.n706 B.n705 10.6151
R2542 B.n707 B.n706 10.6151
R2543 B.n707 B.n402 10.6151
R2544 B.n717 B.n402 10.6151
R2545 B.n718 B.n717 10.6151
R2546 B.n719 B.n718 10.6151
R2547 B.n719 B.n394 10.6151
R2548 B.n729 B.n394 10.6151
R2549 B.n730 B.n729 10.6151
R2550 B.n731 B.n730 10.6151
R2551 B.n731 B.n386 10.6151
R2552 B.n741 B.n386 10.6151
R2553 B.n742 B.n741 10.6151
R2554 B.n743 B.n742 10.6151
R2555 B.n743 B.n378 10.6151
R2556 B.n754 B.n378 10.6151
R2557 B.n755 B.n754 10.6151
R2558 B.n756 B.n755 10.6151
R2559 B.n756 B.n371 10.6151
R2560 B.n766 B.n371 10.6151
R2561 B.n767 B.n766 10.6151
R2562 B.n768 B.n767 10.6151
R2563 B.n768 B.n363 10.6151
R2564 B.n778 B.n363 10.6151
R2565 B.n779 B.n778 10.6151
R2566 B.n780 B.n779 10.6151
R2567 B.n780 B.n355 10.6151
R2568 B.n790 B.n355 10.6151
R2569 B.n791 B.n790 10.6151
R2570 B.n792 B.n791 10.6151
R2571 B.n792 B.n347 10.6151
R2572 B.n802 B.n347 10.6151
R2573 B.n803 B.n802 10.6151
R2574 B.n804 B.n803 10.6151
R2575 B.n804 B.n339 10.6151
R2576 B.n815 B.n339 10.6151
R2577 B.n816 B.n815 10.6151
R2578 B.n817 B.n816 10.6151
R2579 B.n817 B.n332 10.6151
R2580 B.n828 B.n332 10.6151
R2581 B.n829 B.n828 10.6151
R2582 B.n830 B.n829 10.6151
R2583 B.n830 B.n0 10.6151
R2584 B.n1021 B.n1 10.6151
R2585 B.n1021 B.n1020 10.6151
R2586 B.n1020 B.n1019 10.6151
R2587 B.n1019 B.n10 10.6151
R2588 B.n1013 B.n10 10.6151
R2589 B.n1013 B.n1012 10.6151
R2590 B.n1012 B.n1011 10.6151
R2591 B.n1011 B.n16 10.6151
R2592 B.n1005 B.n16 10.6151
R2593 B.n1005 B.n1004 10.6151
R2594 B.n1004 B.n1003 10.6151
R2595 B.n1003 B.n24 10.6151
R2596 B.n997 B.n24 10.6151
R2597 B.n997 B.n996 10.6151
R2598 B.n996 B.n995 10.6151
R2599 B.n995 B.n31 10.6151
R2600 B.n989 B.n31 10.6151
R2601 B.n989 B.n988 10.6151
R2602 B.n988 B.n987 10.6151
R2603 B.n987 B.n38 10.6151
R2604 B.n981 B.n38 10.6151
R2605 B.n981 B.n980 10.6151
R2606 B.n980 B.n979 10.6151
R2607 B.n979 B.n45 10.6151
R2608 B.n973 B.n45 10.6151
R2609 B.n973 B.n972 10.6151
R2610 B.n972 B.n971 10.6151
R2611 B.n971 B.n51 10.6151
R2612 B.n965 B.n51 10.6151
R2613 B.n965 B.n964 10.6151
R2614 B.n964 B.n963 10.6151
R2615 B.n963 B.n59 10.6151
R2616 B.n957 B.n59 10.6151
R2617 B.n957 B.n956 10.6151
R2618 B.n956 B.n955 10.6151
R2619 B.n955 B.n66 10.6151
R2620 B.n949 B.n66 10.6151
R2621 B.n949 B.n948 10.6151
R2622 B.n948 B.n947 10.6151
R2623 B.n947 B.n73 10.6151
R2624 B.n941 B.n73 10.6151
R2625 B.n941 B.n940 10.6151
R2626 B.n940 B.n939 10.6151
R2627 B.n939 B.n80 10.6151
R2628 B.n933 B.n80 10.6151
R2629 B.n933 B.n932 10.6151
R2630 B.n932 B.n931 10.6151
R2631 B.n931 B.n87 10.6151
R2632 B.n925 B.n87 10.6151
R2633 B.n925 B.n924 10.6151
R2634 B.n924 B.n923 10.6151
R2635 B.n923 B.n94 10.6151
R2636 B.n917 B.n94 10.6151
R2637 B.n917 B.n916 10.6151
R2638 B.n916 B.n915 10.6151
R2639 B.n915 B.n101 10.6151
R2640 B.n231 B.n230 9.36635
R2641 B.n253 B.n252 9.36635
R2642 B.n585 B.n486 9.36635
R2643 B.n562 B.n489 9.36635
R2644 B.n424 B.t8 5.32254
R2645 B.n727 B.t21 5.32254
R2646 B.n953 B.t1 5.32254
R2647 B.t12 B.n928 5.32254
R2648 B.n758 B.t5 3.99203
R2649 B.n975 B.t3 3.99203
R2650 B.n1027 B.n0 2.81026
R2651 B.n1027 B.n1 2.81026
R2652 B.n232 B.n231 1.24928
R2653 B.n252 B.n251 1.24928
R2654 B.n582 B.n486 1.24928
R2655 B.n565 B.n489 1.24928
R2656 VP.n21 VP.n20 161.3
R2657 VP.n22 VP.n17 161.3
R2658 VP.n24 VP.n23 161.3
R2659 VP.n25 VP.n16 161.3
R2660 VP.n27 VP.n26 161.3
R2661 VP.n28 VP.n15 161.3
R2662 VP.n30 VP.n29 161.3
R2663 VP.n32 VP.n14 161.3
R2664 VP.n34 VP.n33 161.3
R2665 VP.n35 VP.n13 161.3
R2666 VP.n37 VP.n36 161.3
R2667 VP.n38 VP.n12 161.3
R2668 VP.n40 VP.n39 161.3
R2669 VP.n73 VP.n72 161.3
R2670 VP.n71 VP.n1 161.3
R2671 VP.n70 VP.n69 161.3
R2672 VP.n68 VP.n2 161.3
R2673 VP.n67 VP.n66 161.3
R2674 VP.n65 VP.n3 161.3
R2675 VP.n63 VP.n62 161.3
R2676 VP.n61 VP.n4 161.3
R2677 VP.n60 VP.n59 161.3
R2678 VP.n58 VP.n5 161.3
R2679 VP.n57 VP.n56 161.3
R2680 VP.n55 VP.n6 161.3
R2681 VP.n54 VP.n53 161.3
R2682 VP.n51 VP.n7 161.3
R2683 VP.n50 VP.n49 161.3
R2684 VP.n48 VP.n8 161.3
R2685 VP.n47 VP.n46 161.3
R2686 VP.n45 VP.n9 161.3
R2687 VP.n44 VP.n43 161.3
R2688 VP.n18 VP.t5 122.287
R2689 VP.n10 VP.t6 90.4558
R2690 VP.n52 VP.t4 90.4558
R2691 VP.n64 VP.t7 90.4558
R2692 VP.n0 VP.t2 90.4558
R2693 VP.n11 VP.t0 90.4558
R2694 VP.n31 VP.t1 90.4558
R2695 VP.n19 VP.t3 90.4558
R2696 VP.n19 VP.n18 66.0722
R2697 VP.n42 VP.n10 65.8996
R2698 VP.n74 VP.n0 65.8996
R2699 VP.n41 VP.n11 65.8996
R2700 VP.n46 VP.n8 56.5617
R2701 VP.n70 VP.n2 56.5617
R2702 VP.n37 VP.n13 56.5617
R2703 VP.n42 VP.n41 52.3935
R2704 VP.n58 VP.n57 40.577
R2705 VP.n59 VP.n58 40.577
R2706 VP.n26 VP.n25 40.577
R2707 VP.n25 VP.n24 40.577
R2708 VP.n45 VP.n44 24.5923
R2709 VP.n46 VP.n45 24.5923
R2710 VP.n50 VP.n8 24.5923
R2711 VP.n51 VP.n50 24.5923
R2712 VP.n53 VP.n6 24.5923
R2713 VP.n57 VP.n6 24.5923
R2714 VP.n59 VP.n4 24.5923
R2715 VP.n63 VP.n4 24.5923
R2716 VP.n66 VP.n65 24.5923
R2717 VP.n66 VP.n2 24.5923
R2718 VP.n71 VP.n70 24.5923
R2719 VP.n72 VP.n71 24.5923
R2720 VP.n38 VP.n37 24.5923
R2721 VP.n39 VP.n38 24.5923
R2722 VP.n26 VP.n15 24.5923
R2723 VP.n30 VP.n15 24.5923
R2724 VP.n33 VP.n32 24.5923
R2725 VP.n33 VP.n13 24.5923
R2726 VP.n20 VP.n17 24.5923
R2727 VP.n24 VP.n17 24.5923
R2728 VP.n44 VP.n10 24.3464
R2729 VP.n72 VP.n0 24.3464
R2730 VP.n39 VP.n11 24.3464
R2731 VP.n52 VP.n51 16.477
R2732 VP.n65 VP.n64 16.477
R2733 VP.n32 VP.n31 16.477
R2734 VP.n53 VP.n52 8.11581
R2735 VP.n64 VP.n63 8.11581
R2736 VP.n31 VP.n30 8.11581
R2737 VP.n20 VP.n19 8.11581
R2738 VP.n21 VP.n18 5.23308
R2739 VP.n41 VP.n40 0.354861
R2740 VP.n43 VP.n42 0.354861
R2741 VP.n74 VP.n73 0.354861
R2742 VP VP.n74 0.267071
R2743 VP.n22 VP.n21 0.189894
R2744 VP.n23 VP.n22 0.189894
R2745 VP.n23 VP.n16 0.189894
R2746 VP.n27 VP.n16 0.189894
R2747 VP.n28 VP.n27 0.189894
R2748 VP.n29 VP.n28 0.189894
R2749 VP.n29 VP.n14 0.189894
R2750 VP.n34 VP.n14 0.189894
R2751 VP.n35 VP.n34 0.189894
R2752 VP.n36 VP.n35 0.189894
R2753 VP.n36 VP.n12 0.189894
R2754 VP.n40 VP.n12 0.189894
R2755 VP.n43 VP.n9 0.189894
R2756 VP.n47 VP.n9 0.189894
R2757 VP.n48 VP.n47 0.189894
R2758 VP.n49 VP.n48 0.189894
R2759 VP.n49 VP.n7 0.189894
R2760 VP.n54 VP.n7 0.189894
R2761 VP.n55 VP.n54 0.189894
R2762 VP.n56 VP.n55 0.189894
R2763 VP.n56 VP.n5 0.189894
R2764 VP.n60 VP.n5 0.189894
R2765 VP.n61 VP.n60 0.189894
R2766 VP.n62 VP.n61 0.189894
R2767 VP.n62 VP.n3 0.189894
R2768 VP.n67 VP.n3 0.189894
R2769 VP.n68 VP.n67 0.189894
R2770 VP.n69 VP.n68 0.189894
R2771 VP.n69 VP.n1 0.189894
R2772 VP.n73 VP.n1 0.189894
R2773 VDD1 VDD1.n0 67.1447
R2774 VDD1.n3 VDD1.n2 67.0311
R2775 VDD1.n3 VDD1.n1 67.0311
R2776 VDD1.n5 VDD1.n4 65.6502
R2777 VDD1.n5 VDD1.n3 46.9233
R2778 VDD1.n4 VDD1.t6 1.75894
R2779 VDD1.n4 VDD1.t7 1.75894
R2780 VDD1.n0 VDD1.t2 1.75894
R2781 VDD1.n0 VDD1.t4 1.75894
R2782 VDD1.n2 VDD1.t0 1.75894
R2783 VDD1.n2 VDD1.t5 1.75894
R2784 VDD1.n1 VDD1.t1 1.75894
R2785 VDD1.n1 VDD1.t3 1.75894
R2786 VDD1 VDD1.n5 1.37766
C0 VP VDD2 0.562687f
C1 VN VP 8.00764f
C2 VP VDD1 8.80651f
C3 VTAIL VP 8.98732f
C4 VN VDD2 8.39832f
C5 VDD1 VDD2 1.98659f
C6 VTAIL VDD2 8.01935f
C7 VN VDD1 0.152903f
C8 VN VTAIL 8.973209f
C9 VTAIL VDD1 7.96226f
C10 VDD2 B 5.660152f
C11 VDD1 B 6.143567f
C12 VTAIL B 10.309671f
C13 VN B 16.98502f
C14 VP B 15.613184f
C15 VDD1.t2 B 0.218818f
C16 VDD1.t4 B 0.218818f
C17 VDD1.n0 B 1.96504f
C18 VDD1.t1 B 0.218818f
C19 VDD1.t3 B 0.218818f
C20 VDD1.n1 B 1.96395f
C21 VDD1.t0 B 0.218818f
C22 VDD1.t5 B 0.218818f
C23 VDD1.n2 B 1.96395f
C24 VDD1.n3 B 3.43788f
C25 VDD1.t6 B 0.218818f
C26 VDD1.t7 B 0.218818f
C27 VDD1.n4 B 1.95286f
C28 VDD1.n5 B 3.00296f
C29 VP.t2 B 1.90629f
C30 VP.n0 B 0.761664f
C31 VP.n1 B 0.020751f
C32 VP.n2 B 0.034758f
C33 VP.n3 B 0.020751f
C34 VP.t7 B 1.90629f
C35 VP.n4 B 0.038481f
C36 VP.n5 B 0.020751f
C37 VP.n6 B 0.038481f
C38 VP.n7 B 0.020751f
C39 VP.t4 B 1.90629f
C40 VP.n8 B 0.034758f
C41 VP.n9 B 0.020751f
C42 VP.t6 B 1.90629f
C43 VP.n10 B 0.761664f
C44 VP.t0 B 1.90629f
C45 VP.n11 B 0.761664f
C46 VP.n12 B 0.020751f
C47 VP.n13 B 0.034758f
C48 VP.n14 B 0.020751f
C49 VP.t1 B 1.90629f
C50 VP.n15 B 0.038481f
C51 VP.n16 B 0.020751f
C52 VP.n17 B 0.038481f
C53 VP.t5 B 2.11871f
C54 VP.n18 B 0.713095f
C55 VP.t3 B 1.90629f
C56 VP.n19 B 0.736418f
C57 VP.n20 B 0.025753f
C58 VP.n21 B 0.222516f
C59 VP.n22 B 0.020751f
C60 VP.n23 B 0.020751f
C61 VP.n24 B 0.041025f
C62 VP.n25 B 0.01676f
C63 VP.n26 B 0.041025f
C64 VP.n27 B 0.020751f
C65 VP.n28 B 0.020751f
C66 VP.n29 B 0.020751f
C67 VP.n30 B 0.025753f
C68 VP.n31 B 0.673812f
C69 VP.n32 B 0.032212f
C70 VP.n33 B 0.038481f
C71 VP.n34 B 0.020751f
C72 VP.n35 B 0.020751f
C73 VP.n36 B 0.020751f
C74 VP.n37 B 0.025572f
C75 VP.n38 B 0.038481f
C76 VP.n39 B 0.038291f
C77 VP.n40 B 0.033486f
C78 VP.n41 B 1.25094f
C79 VP.n42 B 1.26522f
C80 VP.n43 B 0.033486f
C81 VP.n44 B 0.038291f
C82 VP.n45 B 0.038481f
C83 VP.n46 B 0.025572f
C84 VP.n47 B 0.020751f
C85 VP.n48 B 0.020751f
C86 VP.n49 B 0.020751f
C87 VP.n50 B 0.038481f
C88 VP.n51 B 0.032212f
C89 VP.n52 B 0.673812f
C90 VP.n53 B 0.025753f
C91 VP.n54 B 0.020751f
C92 VP.n55 B 0.020751f
C93 VP.n56 B 0.020751f
C94 VP.n57 B 0.041025f
C95 VP.n58 B 0.01676f
C96 VP.n59 B 0.041025f
C97 VP.n60 B 0.020751f
C98 VP.n61 B 0.020751f
C99 VP.n62 B 0.020751f
C100 VP.n63 B 0.025753f
C101 VP.n64 B 0.673812f
C102 VP.n65 B 0.032212f
C103 VP.n66 B 0.038481f
C104 VP.n67 B 0.020751f
C105 VP.n68 B 0.020751f
C106 VP.n69 B 0.020751f
C107 VP.n70 B 0.025572f
C108 VP.n71 B 0.038481f
C109 VP.n72 B 0.038291f
C110 VP.n73 B 0.033486f
C111 VP.n74 B 0.038804f
C112 VDD2.t5 B 0.214769f
C113 VDD2.t0 B 0.214769f
C114 VDD2.n0 B 1.92761f
C115 VDD2.t3 B 0.214769f
C116 VDD2.t7 B 0.214769f
C117 VDD2.n1 B 1.92761f
C118 VDD2.n2 B 3.32418f
C119 VDD2.t6 B 0.214769f
C120 VDD2.t4 B 0.214769f
C121 VDD2.n3 B 1.91672f
C122 VDD2.n4 B 2.91738f
C123 VDD2.t1 B 0.214769f
C124 VDD2.t2 B 0.214769f
C125 VDD2.n5 B 1.92758f
C126 VTAIL.t13 B 0.181588f
C127 VTAIL.t8 B 0.181588f
C128 VTAIL.n0 B 1.5677f
C129 VTAIL.n1 B 0.376921f
C130 VTAIL.n2 B 0.011515f
C131 VTAIL.n3 B 0.02592f
C132 VTAIL.n4 B 0.011611f
C133 VTAIL.n5 B 0.020408f
C134 VTAIL.n6 B 0.010966f
C135 VTAIL.n7 B 0.02592f
C136 VTAIL.n8 B 0.011611f
C137 VTAIL.n9 B 0.020408f
C138 VTAIL.n10 B 0.010966f
C139 VTAIL.n11 B 0.02592f
C140 VTAIL.n12 B 0.011611f
C141 VTAIL.n13 B 0.020408f
C142 VTAIL.n14 B 0.010966f
C143 VTAIL.n15 B 0.02592f
C144 VTAIL.n16 B 0.011611f
C145 VTAIL.n17 B 0.020408f
C146 VTAIL.n18 B 0.010966f
C147 VTAIL.n19 B 0.02592f
C148 VTAIL.n20 B 0.011611f
C149 VTAIL.n21 B 0.113968f
C150 VTAIL.t10 B 0.042478f
C151 VTAIL.n22 B 0.01944f
C152 VTAIL.n23 B 0.015312f
C153 VTAIL.n24 B 0.010966f
C154 VTAIL.n25 B 0.977956f
C155 VTAIL.n26 B 0.020408f
C156 VTAIL.n27 B 0.010966f
C157 VTAIL.n28 B 0.011611f
C158 VTAIL.n29 B 0.02592f
C159 VTAIL.n30 B 0.02592f
C160 VTAIL.n31 B 0.011611f
C161 VTAIL.n32 B 0.010966f
C162 VTAIL.n33 B 0.020408f
C163 VTAIL.n34 B 0.020408f
C164 VTAIL.n35 B 0.010966f
C165 VTAIL.n36 B 0.011611f
C166 VTAIL.n37 B 0.02592f
C167 VTAIL.n38 B 0.02592f
C168 VTAIL.n39 B 0.011611f
C169 VTAIL.n40 B 0.010966f
C170 VTAIL.n41 B 0.020408f
C171 VTAIL.n42 B 0.020408f
C172 VTAIL.n43 B 0.010966f
C173 VTAIL.n44 B 0.011611f
C174 VTAIL.n45 B 0.02592f
C175 VTAIL.n46 B 0.02592f
C176 VTAIL.n47 B 0.011611f
C177 VTAIL.n48 B 0.010966f
C178 VTAIL.n49 B 0.020408f
C179 VTAIL.n50 B 0.020408f
C180 VTAIL.n51 B 0.010966f
C181 VTAIL.n52 B 0.011611f
C182 VTAIL.n53 B 0.02592f
C183 VTAIL.n54 B 0.02592f
C184 VTAIL.n55 B 0.011611f
C185 VTAIL.n56 B 0.010966f
C186 VTAIL.n57 B 0.020408f
C187 VTAIL.n58 B 0.053305f
C188 VTAIL.n59 B 0.010966f
C189 VTAIL.n60 B 0.011611f
C190 VTAIL.n61 B 0.05173f
C191 VTAIL.n62 B 0.0443f
C192 VTAIL.n63 B 0.238987f
C193 VTAIL.n64 B 0.011515f
C194 VTAIL.n65 B 0.02592f
C195 VTAIL.n66 B 0.011611f
C196 VTAIL.n67 B 0.020408f
C197 VTAIL.n68 B 0.010966f
C198 VTAIL.n69 B 0.02592f
C199 VTAIL.n70 B 0.011611f
C200 VTAIL.n71 B 0.020408f
C201 VTAIL.n72 B 0.010966f
C202 VTAIL.n73 B 0.02592f
C203 VTAIL.n74 B 0.011611f
C204 VTAIL.n75 B 0.020408f
C205 VTAIL.n76 B 0.010966f
C206 VTAIL.n77 B 0.02592f
C207 VTAIL.n78 B 0.011611f
C208 VTAIL.n79 B 0.020408f
C209 VTAIL.n80 B 0.010966f
C210 VTAIL.n81 B 0.02592f
C211 VTAIL.n82 B 0.011611f
C212 VTAIL.n83 B 0.113968f
C213 VTAIL.t6 B 0.042478f
C214 VTAIL.n84 B 0.01944f
C215 VTAIL.n85 B 0.015312f
C216 VTAIL.n86 B 0.010966f
C217 VTAIL.n87 B 0.977956f
C218 VTAIL.n88 B 0.020408f
C219 VTAIL.n89 B 0.010966f
C220 VTAIL.n90 B 0.011611f
C221 VTAIL.n91 B 0.02592f
C222 VTAIL.n92 B 0.02592f
C223 VTAIL.n93 B 0.011611f
C224 VTAIL.n94 B 0.010966f
C225 VTAIL.n95 B 0.020408f
C226 VTAIL.n96 B 0.020408f
C227 VTAIL.n97 B 0.010966f
C228 VTAIL.n98 B 0.011611f
C229 VTAIL.n99 B 0.02592f
C230 VTAIL.n100 B 0.02592f
C231 VTAIL.n101 B 0.011611f
C232 VTAIL.n102 B 0.010966f
C233 VTAIL.n103 B 0.020408f
C234 VTAIL.n104 B 0.020408f
C235 VTAIL.n105 B 0.010966f
C236 VTAIL.n106 B 0.011611f
C237 VTAIL.n107 B 0.02592f
C238 VTAIL.n108 B 0.02592f
C239 VTAIL.n109 B 0.011611f
C240 VTAIL.n110 B 0.010966f
C241 VTAIL.n111 B 0.020408f
C242 VTAIL.n112 B 0.020408f
C243 VTAIL.n113 B 0.010966f
C244 VTAIL.n114 B 0.011611f
C245 VTAIL.n115 B 0.02592f
C246 VTAIL.n116 B 0.02592f
C247 VTAIL.n117 B 0.011611f
C248 VTAIL.n118 B 0.010966f
C249 VTAIL.n119 B 0.020408f
C250 VTAIL.n120 B 0.053305f
C251 VTAIL.n121 B 0.010966f
C252 VTAIL.n122 B 0.011611f
C253 VTAIL.n123 B 0.05173f
C254 VTAIL.n124 B 0.0443f
C255 VTAIL.n125 B 0.238987f
C256 VTAIL.t5 B 0.181588f
C257 VTAIL.t0 B 0.181588f
C258 VTAIL.n126 B 1.5677f
C259 VTAIL.n127 B 0.561866f
C260 VTAIL.n128 B 0.011515f
C261 VTAIL.n129 B 0.02592f
C262 VTAIL.n130 B 0.011611f
C263 VTAIL.n131 B 0.020408f
C264 VTAIL.n132 B 0.010966f
C265 VTAIL.n133 B 0.02592f
C266 VTAIL.n134 B 0.011611f
C267 VTAIL.n135 B 0.020408f
C268 VTAIL.n136 B 0.010966f
C269 VTAIL.n137 B 0.02592f
C270 VTAIL.n138 B 0.011611f
C271 VTAIL.n139 B 0.020408f
C272 VTAIL.n140 B 0.010966f
C273 VTAIL.n141 B 0.02592f
C274 VTAIL.n142 B 0.011611f
C275 VTAIL.n143 B 0.020408f
C276 VTAIL.n144 B 0.010966f
C277 VTAIL.n145 B 0.02592f
C278 VTAIL.n146 B 0.011611f
C279 VTAIL.n147 B 0.113968f
C280 VTAIL.t15 B 0.042478f
C281 VTAIL.n148 B 0.01944f
C282 VTAIL.n149 B 0.015312f
C283 VTAIL.n150 B 0.010966f
C284 VTAIL.n151 B 0.977956f
C285 VTAIL.n152 B 0.020408f
C286 VTAIL.n153 B 0.010966f
C287 VTAIL.n154 B 0.011611f
C288 VTAIL.n155 B 0.02592f
C289 VTAIL.n156 B 0.02592f
C290 VTAIL.n157 B 0.011611f
C291 VTAIL.n158 B 0.010966f
C292 VTAIL.n159 B 0.020408f
C293 VTAIL.n160 B 0.020408f
C294 VTAIL.n161 B 0.010966f
C295 VTAIL.n162 B 0.011611f
C296 VTAIL.n163 B 0.02592f
C297 VTAIL.n164 B 0.02592f
C298 VTAIL.n165 B 0.011611f
C299 VTAIL.n166 B 0.010966f
C300 VTAIL.n167 B 0.020408f
C301 VTAIL.n168 B 0.020408f
C302 VTAIL.n169 B 0.010966f
C303 VTAIL.n170 B 0.011611f
C304 VTAIL.n171 B 0.02592f
C305 VTAIL.n172 B 0.02592f
C306 VTAIL.n173 B 0.011611f
C307 VTAIL.n174 B 0.010966f
C308 VTAIL.n175 B 0.020408f
C309 VTAIL.n176 B 0.020408f
C310 VTAIL.n177 B 0.010966f
C311 VTAIL.n178 B 0.011611f
C312 VTAIL.n179 B 0.02592f
C313 VTAIL.n180 B 0.02592f
C314 VTAIL.n181 B 0.011611f
C315 VTAIL.n182 B 0.010966f
C316 VTAIL.n183 B 0.020408f
C317 VTAIL.n184 B 0.053305f
C318 VTAIL.n185 B 0.010966f
C319 VTAIL.n186 B 0.011611f
C320 VTAIL.n187 B 0.05173f
C321 VTAIL.n188 B 0.0443f
C322 VTAIL.n189 B 1.31239f
C323 VTAIL.n190 B 0.011515f
C324 VTAIL.n191 B 0.02592f
C325 VTAIL.n192 B 0.011611f
C326 VTAIL.n193 B 0.020408f
C327 VTAIL.n194 B 0.010966f
C328 VTAIL.n195 B 0.02592f
C329 VTAIL.n196 B 0.011611f
C330 VTAIL.n197 B 0.020408f
C331 VTAIL.n198 B 0.010966f
C332 VTAIL.n199 B 0.02592f
C333 VTAIL.n200 B 0.011611f
C334 VTAIL.n201 B 0.020408f
C335 VTAIL.n202 B 0.010966f
C336 VTAIL.n203 B 0.02592f
C337 VTAIL.n204 B 0.011611f
C338 VTAIL.n205 B 0.020408f
C339 VTAIL.n206 B 0.010966f
C340 VTAIL.n207 B 0.02592f
C341 VTAIL.n208 B 0.011611f
C342 VTAIL.n209 B 0.113968f
C343 VTAIL.t12 B 0.042478f
C344 VTAIL.n210 B 0.01944f
C345 VTAIL.n211 B 0.015312f
C346 VTAIL.n212 B 0.010966f
C347 VTAIL.n213 B 0.977956f
C348 VTAIL.n214 B 0.020408f
C349 VTAIL.n215 B 0.010966f
C350 VTAIL.n216 B 0.011611f
C351 VTAIL.n217 B 0.02592f
C352 VTAIL.n218 B 0.02592f
C353 VTAIL.n219 B 0.011611f
C354 VTAIL.n220 B 0.010966f
C355 VTAIL.n221 B 0.020408f
C356 VTAIL.n222 B 0.020408f
C357 VTAIL.n223 B 0.010966f
C358 VTAIL.n224 B 0.011611f
C359 VTAIL.n225 B 0.02592f
C360 VTAIL.n226 B 0.02592f
C361 VTAIL.n227 B 0.011611f
C362 VTAIL.n228 B 0.010966f
C363 VTAIL.n229 B 0.020408f
C364 VTAIL.n230 B 0.020408f
C365 VTAIL.n231 B 0.010966f
C366 VTAIL.n232 B 0.011611f
C367 VTAIL.n233 B 0.02592f
C368 VTAIL.n234 B 0.02592f
C369 VTAIL.n235 B 0.011611f
C370 VTAIL.n236 B 0.010966f
C371 VTAIL.n237 B 0.020408f
C372 VTAIL.n238 B 0.020408f
C373 VTAIL.n239 B 0.010966f
C374 VTAIL.n240 B 0.011611f
C375 VTAIL.n241 B 0.02592f
C376 VTAIL.n242 B 0.02592f
C377 VTAIL.n243 B 0.011611f
C378 VTAIL.n244 B 0.010966f
C379 VTAIL.n245 B 0.020408f
C380 VTAIL.n246 B 0.053305f
C381 VTAIL.n247 B 0.010966f
C382 VTAIL.n248 B 0.011611f
C383 VTAIL.n249 B 0.05173f
C384 VTAIL.n250 B 0.0443f
C385 VTAIL.n251 B 1.31239f
C386 VTAIL.t7 B 0.181588f
C387 VTAIL.t14 B 0.181588f
C388 VTAIL.n252 B 1.56771f
C389 VTAIL.n253 B 0.561861f
C390 VTAIL.n254 B 0.011515f
C391 VTAIL.n255 B 0.02592f
C392 VTAIL.n256 B 0.011611f
C393 VTAIL.n257 B 0.020408f
C394 VTAIL.n258 B 0.010966f
C395 VTAIL.n259 B 0.02592f
C396 VTAIL.n260 B 0.011611f
C397 VTAIL.n261 B 0.020408f
C398 VTAIL.n262 B 0.010966f
C399 VTAIL.n263 B 0.02592f
C400 VTAIL.n264 B 0.011611f
C401 VTAIL.n265 B 0.020408f
C402 VTAIL.n266 B 0.010966f
C403 VTAIL.n267 B 0.02592f
C404 VTAIL.n268 B 0.011611f
C405 VTAIL.n269 B 0.020408f
C406 VTAIL.n270 B 0.010966f
C407 VTAIL.n271 B 0.02592f
C408 VTAIL.n272 B 0.011611f
C409 VTAIL.n273 B 0.113968f
C410 VTAIL.t11 B 0.042478f
C411 VTAIL.n274 B 0.01944f
C412 VTAIL.n275 B 0.015312f
C413 VTAIL.n276 B 0.010966f
C414 VTAIL.n277 B 0.977956f
C415 VTAIL.n278 B 0.020408f
C416 VTAIL.n279 B 0.010966f
C417 VTAIL.n280 B 0.011611f
C418 VTAIL.n281 B 0.02592f
C419 VTAIL.n282 B 0.02592f
C420 VTAIL.n283 B 0.011611f
C421 VTAIL.n284 B 0.010966f
C422 VTAIL.n285 B 0.020408f
C423 VTAIL.n286 B 0.020408f
C424 VTAIL.n287 B 0.010966f
C425 VTAIL.n288 B 0.011611f
C426 VTAIL.n289 B 0.02592f
C427 VTAIL.n290 B 0.02592f
C428 VTAIL.n291 B 0.011611f
C429 VTAIL.n292 B 0.010966f
C430 VTAIL.n293 B 0.020408f
C431 VTAIL.n294 B 0.020408f
C432 VTAIL.n295 B 0.010966f
C433 VTAIL.n296 B 0.011611f
C434 VTAIL.n297 B 0.02592f
C435 VTAIL.n298 B 0.02592f
C436 VTAIL.n299 B 0.011611f
C437 VTAIL.n300 B 0.010966f
C438 VTAIL.n301 B 0.020408f
C439 VTAIL.n302 B 0.020408f
C440 VTAIL.n303 B 0.010966f
C441 VTAIL.n304 B 0.011611f
C442 VTAIL.n305 B 0.02592f
C443 VTAIL.n306 B 0.02592f
C444 VTAIL.n307 B 0.011611f
C445 VTAIL.n308 B 0.010966f
C446 VTAIL.n309 B 0.020408f
C447 VTAIL.n310 B 0.053305f
C448 VTAIL.n311 B 0.010966f
C449 VTAIL.n312 B 0.011611f
C450 VTAIL.n313 B 0.05173f
C451 VTAIL.n314 B 0.0443f
C452 VTAIL.n315 B 0.238987f
C453 VTAIL.n316 B 0.011515f
C454 VTAIL.n317 B 0.02592f
C455 VTAIL.n318 B 0.011611f
C456 VTAIL.n319 B 0.020408f
C457 VTAIL.n320 B 0.010966f
C458 VTAIL.n321 B 0.02592f
C459 VTAIL.n322 B 0.011611f
C460 VTAIL.n323 B 0.020408f
C461 VTAIL.n324 B 0.010966f
C462 VTAIL.n325 B 0.02592f
C463 VTAIL.n326 B 0.011611f
C464 VTAIL.n327 B 0.020408f
C465 VTAIL.n328 B 0.010966f
C466 VTAIL.n329 B 0.02592f
C467 VTAIL.n330 B 0.011611f
C468 VTAIL.n331 B 0.020408f
C469 VTAIL.n332 B 0.010966f
C470 VTAIL.n333 B 0.02592f
C471 VTAIL.n334 B 0.011611f
C472 VTAIL.n335 B 0.113968f
C473 VTAIL.t4 B 0.042478f
C474 VTAIL.n336 B 0.01944f
C475 VTAIL.n337 B 0.015312f
C476 VTAIL.n338 B 0.010966f
C477 VTAIL.n339 B 0.977956f
C478 VTAIL.n340 B 0.020408f
C479 VTAIL.n341 B 0.010966f
C480 VTAIL.n342 B 0.011611f
C481 VTAIL.n343 B 0.02592f
C482 VTAIL.n344 B 0.02592f
C483 VTAIL.n345 B 0.011611f
C484 VTAIL.n346 B 0.010966f
C485 VTAIL.n347 B 0.020408f
C486 VTAIL.n348 B 0.020408f
C487 VTAIL.n349 B 0.010966f
C488 VTAIL.n350 B 0.011611f
C489 VTAIL.n351 B 0.02592f
C490 VTAIL.n352 B 0.02592f
C491 VTAIL.n353 B 0.011611f
C492 VTAIL.n354 B 0.010966f
C493 VTAIL.n355 B 0.020408f
C494 VTAIL.n356 B 0.020408f
C495 VTAIL.n357 B 0.010966f
C496 VTAIL.n358 B 0.011611f
C497 VTAIL.n359 B 0.02592f
C498 VTAIL.n360 B 0.02592f
C499 VTAIL.n361 B 0.011611f
C500 VTAIL.n362 B 0.010966f
C501 VTAIL.n363 B 0.020408f
C502 VTAIL.n364 B 0.020408f
C503 VTAIL.n365 B 0.010966f
C504 VTAIL.n366 B 0.011611f
C505 VTAIL.n367 B 0.02592f
C506 VTAIL.n368 B 0.02592f
C507 VTAIL.n369 B 0.011611f
C508 VTAIL.n370 B 0.010966f
C509 VTAIL.n371 B 0.020408f
C510 VTAIL.n372 B 0.053305f
C511 VTAIL.n373 B 0.010966f
C512 VTAIL.n374 B 0.011611f
C513 VTAIL.n375 B 0.05173f
C514 VTAIL.n376 B 0.0443f
C515 VTAIL.n377 B 0.238987f
C516 VTAIL.t2 B 0.181588f
C517 VTAIL.t3 B 0.181588f
C518 VTAIL.n378 B 1.56771f
C519 VTAIL.n379 B 0.561861f
C520 VTAIL.n380 B 0.011515f
C521 VTAIL.n381 B 0.02592f
C522 VTAIL.n382 B 0.011611f
C523 VTAIL.n383 B 0.020408f
C524 VTAIL.n384 B 0.010966f
C525 VTAIL.n385 B 0.02592f
C526 VTAIL.n386 B 0.011611f
C527 VTAIL.n387 B 0.020408f
C528 VTAIL.n388 B 0.010966f
C529 VTAIL.n389 B 0.02592f
C530 VTAIL.n390 B 0.011611f
C531 VTAIL.n391 B 0.020408f
C532 VTAIL.n392 B 0.010966f
C533 VTAIL.n393 B 0.02592f
C534 VTAIL.n394 B 0.011611f
C535 VTAIL.n395 B 0.020408f
C536 VTAIL.n396 B 0.010966f
C537 VTAIL.n397 B 0.02592f
C538 VTAIL.n398 B 0.011611f
C539 VTAIL.n399 B 0.113968f
C540 VTAIL.t1 B 0.042478f
C541 VTAIL.n400 B 0.01944f
C542 VTAIL.n401 B 0.015312f
C543 VTAIL.n402 B 0.010966f
C544 VTAIL.n403 B 0.977956f
C545 VTAIL.n404 B 0.020408f
C546 VTAIL.n405 B 0.010966f
C547 VTAIL.n406 B 0.011611f
C548 VTAIL.n407 B 0.02592f
C549 VTAIL.n408 B 0.02592f
C550 VTAIL.n409 B 0.011611f
C551 VTAIL.n410 B 0.010966f
C552 VTAIL.n411 B 0.020408f
C553 VTAIL.n412 B 0.020408f
C554 VTAIL.n413 B 0.010966f
C555 VTAIL.n414 B 0.011611f
C556 VTAIL.n415 B 0.02592f
C557 VTAIL.n416 B 0.02592f
C558 VTAIL.n417 B 0.011611f
C559 VTAIL.n418 B 0.010966f
C560 VTAIL.n419 B 0.020408f
C561 VTAIL.n420 B 0.020408f
C562 VTAIL.n421 B 0.010966f
C563 VTAIL.n422 B 0.011611f
C564 VTAIL.n423 B 0.02592f
C565 VTAIL.n424 B 0.02592f
C566 VTAIL.n425 B 0.011611f
C567 VTAIL.n426 B 0.010966f
C568 VTAIL.n427 B 0.020408f
C569 VTAIL.n428 B 0.020408f
C570 VTAIL.n429 B 0.010966f
C571 VTAIL.n430 B 0.011611f
C572 VTAIL.n431 B 0.02592f
C573 VTAIL.n432 B 0.02592f
C574 VTAIL.n433 B 0.011611f
C575 VTAIL.n434 B 0.010966f
C576 VTAIL.n435 B 0.020408f
C577 VTAIL.n436 B 0.053305f
C578 VTAIL.n437 B 0.010966f
C579 VTAIL.n438 B 0.011611f
C580 VTAIL.n439 B 0.05173f
C581 VTAIL.n440 B 0.0443f
C582 VTAIL.n441 B 1.31239f
C583 VTAIL.n442 B 0.011515f
C584 VTAIL.n443 B 0.02592f
C585 VTAIL.n444 B 0.011611f
C586 VTAIL.n445 B 0.020408f
C587 VTAIL.n446 B 0.010966f
C588 VTAIL.n447 B 0.02592f
C589 VTAIL.n448 B 0.011611f
C590 VTAIL.n449 B 0.020408f
C591 VTAIL.n450 B 0.010966f
C592 VTAIL.n451 B 0.02592f
C593 VTAIL.n452 B 0.011611f
C594 VTAIL.n453 B 0.020408f
C595 VTAIL.n454 B 0.010966f
C596 VTAIL.n455 B 0.02592f
C597 VTAIL.n456 B 0.011611f
C598 VTAIL.n457 B 0.020408f
C599 VTAIL.n458 B 0.010966f
C600 VTAIL.n459 B 0.02592f
C601 VTAIL.n460 B 0.011611f
C602 VTAIL.n461 B 0.113968f
C603 VTAIL.t9 B 0.042478f
C604 VTAIL.n462 B 0.01944f
C605 VTAIL.n463 B 0.015312f
C606 VTAIL.n464 B 0.010966f
C607 VTAIL.n465 B 0.977956f
C608 VTAIL.n466 B 0.020408f
C609 VTAIL.n467 B 0.010966f
C610 VTAIL.n468 B 0.011611f
C611 VTAIL.n469 B 0.02592f
C612 VTAIL.n470 B 0.02592f
C613 VTAIL.n471 B 0.011611f
C614 VTAIL.n472 B 0.010966f
C615 VTAIL.n473 B 0.020408f
C616 VTAIL.n474 B 0.020408f
C617 VTAIL.n475 B 0.010966f
C618 VTAIL.n476 B 0.011611f
C619 VTAIL.n477 B 0.02592f
C620 VTAIL.n478 B 0.02592f
C621 VTAIL.n479 B 0.011611f
C622 VTAIL.n480 B 0.010966f
C623 VTAIL.n481 B 0.020408f
C624 VTAIL.n482 B 0.020408f
C625 VTAIL.n483 B 0.010966f
C626 VTAIL.n484 B 0.011611f
C627 VTAIL.n485 B 0.02592f
C628 VTAIL.n486 B 0.02592f
C629 VTAIL.n487 B 0.011611f
C630 VTAIL.n488 B 0.010966f
C631 VTAIL.n489 B 0.020408f
C632 VTAIL.n490 B 0.020408f
C633 VTAIL.n491 B 0.010966f
C634 VTAIL.n492 B 0.011611f
C635 VTAIL.n493 B 0.02592f
C636 VTAIL.n494 B 0.02592f
C637 VTAIL.n495 B 0.011611f
C638 VTAIL.n496 B 0.010966f
C639 VTAIL.n497 B 0.020408f
C640 VTAIL.n498 B 0.053305f
C641 VTAIL.n499 B 0.010966f
C642 VTAIL.n500 B 0.011611f
C643 VTAIL.n501 B 0.05173f
C644 VTAIL.n502 B 0.0443f
C645 VTAIL.n503 B 1.30856f
C646 VN.t0 B 1.87462f
C647 VN.n0 B 0.749009f
C648 VN.n1 B 0.020406f
C649 VN.n2 B 0.03418f
C650 VN.n3 B 0.020406f
C651 VN.t4 B 1.87462f
C652 VN.n4 B 0.037841f
C653 VN.n5 B 0.020406f
C654 VN.n6 B 0.037841f
C655 VN.t2 B 2.08351f
C656 VN.n7 B 0.701246f
C657 VN.t7 B 1.87462f
C658 VN.n8 B 0.724182f
C659 VN.n9 B 0.025325f
C660 VN.n10 B 0.218819f
C661 VN.n11 B 0.020406f
C662 VN.n12 B 0.020406f
C663 VN.n13 B 0.040344f
C664 VN.n14 B 0.016481f
C665 VN.n15 B 0.040344f
C666 VN.n16 B 0.020406f
C667 VN.n17 B 0.020406f
C668 VN.n18 B 0.020406f
C669 VN.n19 B 0.025325f
C670 VN.n20 B 0.662617f
C671 VN.n21 B 0.031677f
C672 VN.n22 B 0.037841f
C673 VN.n23 B 0.020406f
C674 VN.n24 B 0.020406f
C675 VN.n25 B 0.020406f
C676 VN.n26 B 0.025147f
C677 VN.n27 B 0.037841f
C678 VN.n28 B 0.037655f
C679 VN.n29 B 0.03293f
C680 VN.n30 B 0.038159f
C681 VN.t1 B 1.87462f
C682 VN.n31 B 0.749009f
C683 VN.n32 B 0.020406f
C684 VN.n33 B 0.03418f
C685 VN.n34 B 0.020406f
C686 VN.t3 B 1.87462f
C687 VN.n35 B 0.037841f
C688 VN.n36 B 0.020406f
C689 VN.n37 B 0.037841f
C690 VN.t5 B 2.08351f
C691 VN.n38 B 0.701246f
C692 VN.t6 B 1.87462f
C693 VN.n39 B 0.724182f
C694 VN.n40 B 0.025325f
C695 VN.n41 B 0.218819f
C696 VN.n42 B 0.020406f
C697 VN.n43 B 0.020406f
C698 VN.n44 B 0.040344f
C699 VN.n45 B 0.016481f
C700 VN.n46 B 0.040344f
C701 VN.n47 B 0.020406f
C702 VN.n48 B 0.020406f
C703 VN.n49 B 0.020406f
C704 VN.n50 B 0.025325f
C705 VN.n51 B 0.662617f
C706 VN.n52 B 0.031677f
C707 VN.n53 B 0.037841f
C708 VN.n54 B 0.020406f
C709 VN.n55 B 0.020406f
C710 VN.n56 B 0.020406f
C711 VN.n57 B 0.025147f
C712 VN.n58 B 0.037841f
C713 VN.n59 B 0.037655f
C714 VN.n60 B 0.03293f
C715 VN.n61 B 1.23837f
.ends

