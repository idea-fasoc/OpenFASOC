* NGSPICE file created from diff_pair_sample_0713.ext - technology: sky130A

.subckt diff_pair_sample_0713 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0 ps=0 w=1.15 l=2.41
X1 B.t8 B.t6 B.t7 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0 ps=0 w=1.15 l=2.41
X2 VDD1.t1 VP.t0 VTAIL.t2 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0.4485 ps=3.08 w=1.15 l=2.41
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0.4485 ps=3.08 w=1.15 l=2.41
X4 B.t5 B.t3 B.t4 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0 ps=0 w=1.15 l=2.41
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0.4485 ps=3.08 w=1.15 l=2.41
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0.4485 ps=3.08 w=1.15 l=2.41
X7 B.t2 B.t0 B.t1 w_n2066_n1198# sky130_fd_pr__pfet_01v8 ad=0.4485 pd=3.08 as=0 ps=0 w=1.15 l=2.41
R0 B.n241 B.n32 585
R1 B.n243 B.n242 585
R2 B.n244 B.n31 585
R3 B.n246 B.n245 585
R4 B.n247 B.n30 585
R5 B.n249 B.n248 585
R6 B.n250 B.n29 585
R7 B.n252 B.n251 585
R8 B.n253 B.n28 585
R9 B.n255 B.n254 585
R10 B.n257 B.n25 585
R11 B.n259 B.n258 585
R12 B.n260 B.n24 585
R13 B.n262 B.n261 585
R14 B.n263 B.n23 585
R15 B.n265 B.n264 585
R16 B.n266 B.n22 585
R17 B.n268 B.n267 585
R18 B.n269 B.n19 585
R19 B.n272 B.n271 585
R20 B.n273 B.n18 585
R21 B.n275 B.n274 585
R22 B.n276 B.n17 585
R23 B.n278 B.n277 585
R24 B.n279 B.n16 585
R25 B.n281 B.n280 585
R26 B.n282 B.n15 585
R27 B.n284 B.n283 585
R28 B.n285 B.n14 585
R29 B.n240 B.n239 585
R30 B.n238 B.n33 585
R31 B.n237 B.n236 585
R32 B.n235 B.n34 585
R33 B.n234 B.n233 585
R34 B.n232 B.n35 585
R35 B.n231 B.n230 585
R36 B.n229 B.n36 585
R37 B.n228 B.n227 585
R38 B.n226 B.n37 585
R39 B.n225 B.n224 585
R40 B.n223 B.n38 585
R41 B.n222 B.n221 585
R42 B.n220 B.n39 585
R43 B.n219 B.n218 585
R44 B.n217 B.n40 585
R45 B.n216 B.n215 585
R46 B.n214 B.n41 585
R47 B.n213 B.n212 585
R48 B.n211 B.n42 585
R49 B.n210 B.n209 585
R50 B.n208 B.n43 585
R51 B.n207 B.n206 585
R52 B.n205 B.n44 585
R53 B.n204 B.n203 585
R54 B.n202 B.n45 585
R55 B.n201 B.n200 585
R56 B.n199 B.n46 585
R57 B.n198 B.n197 585
R58 B.n196 B.n47 585
R59 B.n195 B.n194 585
R60 B.n193 B.n48 585
R61 B.n192 B.n191 585
R62 B.n190 B.n49 585
R63 B.n189 B.n188 585
R64 B.n187 B.n50 585
R65 B.n186 B.n185 585
R66 B.n184 B.n51 585
R67 B.n183 B.n182 585
R68 B.n181 B.n52 585
R69 B.n180 B.n179 585
R70 B.n178 B.n53 585
R71 B.n177 B.n176 585
R72 B.n175 B.n54 585
R73 B.n174 B.n173 585
R74 B.n172 B.n55 585
R75 B.n171 B.n170 585
R76 B.n169 B.n56 585
R77 B.n168 B.n167 585
R78 B.n123 B.n122 585
R79 B.n124 B.n75 585
R80 B.n126 B.n125 585
R81 B.n127 B.n74 585
R82 B.n129 B.n128 585
R83 B.n130 B.n73 585
R84 B.n132 B.n131 585
R85 B.n133 B.n72 585
R86 B.n135 B.n134 585
R87 B.n136 B.n69 585
R88 B.n139 B.n138 585
R89 B.n140 B.n68 585
R90 B.n142 B.n141 585
R91 B.n143 B.n67 585
R92 B.n145 B.n144 585
R93 B.n146 B.n66 585
R94 B.n148 B.n147 585
R95 B.n149 B.n65 585
R96 B.n151 B.n150 585
R97 B.n153 B.n152 585
R98 B.n154 B.n61 585
R99 B.n156 B.n155 585
R100 B.n157 B.n60 585
R101 B.n159 B.n158 585
R102 B.n160 B.n59 585
R103 B.n162 B.n161 585
R104 B.n163 B.n58 585
R105 B.n165 B.n164 585
R106 B.n166 B.n57 585
R107 B.n121 B.n76 585
R108 B.n120 B.n119 585
R109 B.n118 B.n77 585
R110 B.n117 B.n116 585
R111 B.n115 B.n78 585
R112 B.n114 B.n113 585
R113 B.n112 B.n79 585
R114 B.n111 B.n110 585
R115 B.n109 B.n80 585
R116 B.n108 B.n107 585
R117 B.n106 B.n81 585
R118 B.n105 B.n104 585
R119 B.n103 B.n82 585
R120 B.n102 B.n101 585
R121 B.n100 B.n83 585
R122 B.n99 B.n98 585
R123 B.n97 B.n84 585
R124 B.n96 B.n95 585
R125 B.n94 B.n85 585
R126 B.n93 B.n92 585
R127 B.n91 B.n86 585
R128 B.n90 B.n89 585
R129 B.n88 B.n87 585
R130 B.n2 B.n0 585
R131 B.n321 B.n1 585
R132 B.n320 B.n319 585
R133 B.n318 B.n3 585
R134 B.n317 B.n316 585
R135 B.n315 B.n4 585
R136 B.n314 B.n313 585
R137 B.n312 B.n5 585
R138 B.n311 B.n310 585
R139 B.n309 B.n6 585
R140 B.n308 B.n307 585
R141 B.n306 B.n7 585
R142 B.n305 B.n304 585
R143 B.n303 B.n8 585
R144 B.n302 B.n301 585
R145 B.n300 B.n9 585
R146 B.n299 B.n298 585
R147 B.n297 B.n10 585
R148 B.n296 B.n295 585
R149 B.n294 B.n11 585
R150 B.n293 B.n292 585
R151 B.n291 B.n12 585
R152 B.n290 B.n289 585
R153 B.n288 B.n13 585
R154 B.n287 B.n286 585
R155 B.n323 B.n322 585
R156 B.n122 B.n121 535.745
R157 B.n286 B.n285 535.745
R158 B.n168 B.n57 535.745
R159 B.n241 B.n240 535.745
R160 B.n62 B.t2 417.248
R161 B.n70 B.t8 417.248
R162 B.n20 B.t10 417.248
R163 B.n26 B.t4 417.248
R164 B.n63 B.t1 364.108
R165 B.n71 B.t7 364.108
R166 B.n21 B.t11 364.108
R167 B.n27 B.t5 364.108
R168 B.n62 B.t0 208.587
R169 B.n70 B.t6 208.587
R170 B.n20 B.t9 208.587
R171 B.n26 B.t3 208.587
R172 B.n121 B.n120 163.367
R173 B.n120 B.n77 163.367
R174 B.n116 B.n77 163.367
R175 B.n116 B.n115 163.367
R176 B.n115 B.n114 163.367
R177 B.n114 B.n79 163.367
R178 B.n110 B.n79 163.367
R179 B.n110 B.n109 163.367
R180 B.n109 B.n108 163.367
R181 B.n108 B.n81 163.367
R182 B.n104 B.n81 163.367
R183 B.n104 B.n103 163.367
R184 B.n103 B.n102 163.367
R185 B.n102 B.n83 163.367
R186 B.n98 B.n83 163.367
R187 B.n98 B.n97 163.367
R188 B.n97 B.n96 163.367
R189 B.n96 B.n85 163.367
R190 B.n92 B.n85 163.367
R191 B.n92 B.n91 163.367
R192 B.n91 B.n90 163.367
R193 B.n90 B.n87 163.367
R194 B.n87 B.n2 163.367
R195 B.n322 B.n2 163.367
R196 B.n322 B.n321 163.367
R197 B.n321 B.n320 163.367
R198 B.n320 B.n3 163.367
R199 B.n316 B.n3 163.367
R200 B.n316 B.n315 163.367
R201 B.n315 B.n314 163.367
R202 B.n314 B.n5 163.367
R203 B.n310 B.n5 163.367
R204 B.n310 B.n309 163.367
R205 B.n309 B.n308 163.367
R206 B.n308 B.n7 163.367
R207 B.n304 B.n7 163.367
R208 B.n304 B.n303 163.367
R209 B.n303 B.n302 163.367
R210 B.n302 B.n9 163.367
R211 B.n298 B.n9 163.367
R212 B.n298 B.n297 163.367
R213 B.n297 B.n296 163.367
R214 B.n296 B.n11 163.367
R215 B.n292 B.n11 163.367
R216 B.n292 B.n291 163.367
R217 B.n291 B.n290 163.367
R218 B.n290 B.n13 163.367
R219 B.n286 B.n13 163.367
R220 B.n122 B.n75 163.367
R221 B.n126 B.n75 163.367
R222 B.n127 B.n126 163.367
R223 B.n128 B.n127 163.367
R224 B.n128 B.n73 163.367
R225 B.n132 B.n73 163.367
R226 B.n133 B.n132 163.367
R227 B.n134 B.n133 163.367
R228 B.n134 B.n69 163.367
R229 B.n139 B.n69 163.367
R230 B.n140 B.n139 163.367
R231 B.n141 B.n140 163.367
R232 B.n141 B.n67 163.367
R233 B.n145 B.n67 163.367
R234 B.n146 B.n145 163.367
R235 B.n147 B.n146 163.367
R236 B.n147 B.n65 163.367
R237 B.n151 B.n65 163.367
R238 B.n152 B.n151 163.367
R239 B.n152 B.n61 163.367
R240 B.n156 B.n61 163.367
R241 B.n157 B.n156 163.367
R242 B.n158 B.n157 163.367
R243 B.n158 B.n59 163.367
R244 B.n162 B.n59 163.367
R245 B.n163 B.n162 163.367
R246 B.n164 B.n163 163.367
R247 B.n164 B.n57 163.367
R248 B.n169 B.n168 163.367
R249 B.n170 B.n169 163.367
R250 B.n170 B.n55 163.367
R251 B.n174 B.n55 163.367
R252 B.n175 B.n174 163.367
R253 B.n176 B.n175 163.367
R254 B.n176 B.n53 163.367
R255 B.n180 B.n53 163.367
R256 B.n181 B.n180 163.367
R257 B.n182 B.n181 163.367
R258 B.n182 B.n51 163.367
R259 B.n186 B.n51 163.367
R260 B.n187 B.n186 163.367
R261 B.n188 B.n187 163.367
R262 B.n188 B.n49 163.367
R263 B.n192 B.n49 163.367
R264 B.n193 B.n192 163.367
R265 B.n194 B.n193 163.367
R266 B.n194 B.n47 163.367
R267 B.n198 B.n47 163.367
R268 B.n199 B.n198 163.367
R269 B.n200 B.n199 163.367
R270 B.n200 B.n45 163.367
R271 B.n204 B.n45 163.367
R272 B.n205 B.n204 163.367
R273 B.n206 B.n205 163.367
R274 B.n206 B.n43 163.367
R275 B.n210 B.n43 163.367
R276 B.n211 B.n210 163.367
R277 B.n212 B.n211 163.367
R278 B.n212 B.n41 163.367
R279 B.n216 B.n41 163.367
R280 B.n217 B.n216 163.367
R281 B.n218 B.n217 163.367
R282 B.n218 B.n39 163.367
R283 B.n222 B.n39 163.367
R284 B.n223 B.n222 163.367
R285 B.n224 B.n223 163.367
R286 B.n224 B.n37 163.367
R287 B.n228 B.n37 163.367
R288 B.n229 B.n228 163.367
R289 B.n230 B.n229 163.367
R290 B.n230 B.n35 163.367
R291 B.n234 B.n35 163.367
R292 B.n235 B.n234 163.367
R293 B.n236 B.n235 163.367
R294 B.n236 B.n33 163.367
R295 B.n240 B.n33 163.367
R296 B.n285 B.n284 163.367
R297 B.n284 B.n15 163.367
R298 B.n280 B.n15 163.367
R299 B.n280 B.n279 163.367
R300 B.n279 B.n278 163.367
R301 B.n278 B.n17 163.367
R302 B.n274 B.n17 163.367
R303 B.n274 B.n273 163.367
R304 B.n273 B.n272 163.367
R305 B.n272 B.n19 163.367
R306 B.n267 B.n19 163.367
R307 B.n267 B.n266 163.367
R308 B.n266 B.n265 163.367
R309 B.n265 B.n23 163.367
R310 B.n261 B.n23 163.367
R311 B.n261 B.n260 163.367
R312 B.n260 B.n259 163.367
R313 B.n259 B.n25 163.367
R314 B.n254 B.n25 163.367
R315 B.n254 B.n253 163.367
R316 B.n253 B.n252 163.367
R317 B.n252 B.n29 163.367
R318 B.n248 B.n29 163.367
R319 B.n248 B.n247 163.367
R320 B.n247 B.n246 163.367
R321 B.n246 B.n31 163.367
R322 B.n242 B.n31 163.367
R323 B.n242 B.n241 163.367
R324 B.n64 B.n63 59.5399
R325 B.n137 B.n71 59.5399
R326 B.n270 B.n21 59.5399
R327 B.n256 B.n27 59.5399
R328 B.n63 B.n62 53.1399
R329 B.n71 B.n70 53.1399
R330 B.n21 B.n20 53.1399
R331 B.n27 B.n26 53.1399
R332 B.n287 B.n14 34.8103
R333 B.n239 B.n32 34.8103
R334 B.n167 B.n166 34.8103
R335 B.n123 B.n76 34.8103
R336 B B.n323 18.0485
R337 B.n283 B.n14 10.6151
R338 B.n283 B.n282 10.6151
R339 B.n282 B.n281 10.6151
R340 B.n281 B.n16 10.6151
R341 B.n277 B.n16 10.6151
R342 B.n277 B.n276 10.6151
R343 B.n276 B.n275 10.6151
R344 B.n275 B.n18 10.6151
R345 B.n271 B.n18 10.6151
R346 B.n269 B.n268 10.6151
R347 B.n268 B.n22 10.6151
R348 B.n264 B.n22 10.6151
R349 B.n264 B.n263 10.6151
R350 B.n263 B.n262 10.6151
R351 B.n262 B.n24 10.6151
R352 B.n258 B.n24 10.6151
R353 B.n258 B.n257 10.6151
R354 B.n255 B.n28 10.6151
R355 B.n251 B.n28 10.6151
R356 B.n251 B.n250 10.6151
R357 B.n250 B.n249 10.6151
R358 B.n249 B.n30 10.6151
R359 B.n245 B.n30 10.6151
R360 B.n245 B.n244 10.6151
R361 B.n244 B.n243 10.6151
R362 B.n243 B.n32 10.6151
R363 B.n167 B.n56 10.6151
R364 B.n171 B.n56 10.6151
R365 B.n172 B.n171 10.6151
R366 B.n173 B.n172 10.6151
R367 B.n173 B.n54 10.6151
R368 B.n177 B.n54 10.6151
R369 B.n178 B.n177 10.6151
R370 B.n179 B.n178 10.6151
R371 B.n179 B.n52 10.6151
R372 B.n183 B.n52 10.6151
R373 B.n184 B.n183 10.6151
R374 B.n185 B.n184 10.6151
R375 B.n185 B.n50 10.6151
R376 B.n189 B.n50 10.6151
R377 B.n190 B.n189 10.6151
R378 B.n191 B.n190 10.6151
R379 B.n191 B.n48 10.6151
R380 B.n195 B.n48 10.6151
R381 B.n196 B.n195 10.6151
R382 B.n197 B.n196 10.6151
R383 B.n197 B.n46 10.6151
R384 B.n201 B.n46 10.6151
R385 B.n202 B.n201 10.6151
R386 B.n203 B.n202 10.6151
R387 B.n203 B.n44 10.6151
R388 B.n207 B.n44 10.6151
R389 B.n208 B.n207 10.6151
R390 B.n209 B.n208 10.6151
R391 B.n209 B.n42 10.6151
R392 B.n213 B.n42 10.6151
R393 B.n214 B.n213 10.6151
R394 B.n215 B.n214 10.6151
R395 B.n215 B.n40 10.6151
R396 B.n219 B.n40 10.6151
R397 B.n220 B.n219 10.6151
R398 B.n221 B.n220 10.6151
R399 B.n221 B.n38 10.6151
R400 B.n225 B.n38 10.6151
R401 B.n226 B.n225 10.6151
R402 B.n227 B.n226 10.6151
R403 B.n227 B.n36 10.6151
R404 B.n231 B.n36 10.6151
R405 B.n232 B.n231 10.6151
R406 B.n233 B.n232 10.6151
R407 B.n233 B.n34 10.6151
R408 B.n237 B.n34 10.6151
R409 B.n238 B.n237 10.6151
R410 B.n239 B.n238 10.6151
R411 B.n124 B.n123 10.6151
R412 B.n125 B.n124 10.6151
R413 B.n125 B.n74 10.6151
R414 B.n129 B.n74 10.6151
R415 B.n130 B.n129 10.6151
R416 B.n131 B.n130 10.6151
R417 B.n131 B.n72 10.6151
R418 B.n135 B.n72 10.6151
R419 B.n136 B.n135 10.6151
R420 B.n138 B.n68 10.6151
R421 B.n142 B.n68 10.6151
R422 B.n143 B.n142 10.6151
R423 B.n144 B.n143 10.6151
R424 B.n144 B.n66 10.6151
R425 B.n148 B.n66 10.6151
R426 B.n149 B.n148 10.6151
R427 B.n150 B.n149 10.6151
R428 B.n154 B.n153 10.6151
R429 B.n155 B.n154 10.6151
R430 B.n155 B.n60 10.6151
R431 B.n159 B.n60 10.6151
R432 B.n160 B.n159 10.6151
R433 B.n161 B.n160 10.6151
R434 B.n161 B.n58 10.6151
R435 B.n165 B.n58 10.6151
R436 B.n166 B.n165 10.6151
R437 B.n119 B.n76 10.6151
R438 B.n119 B.n118 10.6151
R439 B.n118 B.n117 10.6151
R440 B.n117 B.n78 10.6151
R441 B.n113 B.n78 10.6151
R442 B.n113 B.n112 10.6151
R443 B.n112 B.n111 10.6151
R444 B.n111 B.n80 10.6151
R445 B.n107 B.n80 10.6151
R446 B.n107 B.n106 10.6151
R447 B.n106 B.n105 10.6151
R448 B.n105 B.n82 10.6151
R449 B.n101 B.n82 10.6151
R450 B.n101 B.n100 10.6151
R451 B.n100 B.n99 10.6151
R452 B.n99 B.n84 10.6151
R453 B.n95 B.n84 10.6151
R454 B.n95 B.n94 10.6151
R455 B.n94 B.n93 10.6151
R456 B.n93 B.n86 10.6151
R457 B.n89 B.n86 10.6151
R458 B.n89 B.n88 10.6151
R459 B.n88 B.n0 10.6151
R460 B.n319 B.n1 10.6151
R461 B.n319 B.n318 10.6151
R462 B.n318 B.n317 10.6151
R463 B.n317 B.n4 10.6151
R464 B.n313 B.n4 10.6151
R465 B.n313 B.n312 10.6151
R466 B.n312 B.n311 10.6151
R467 B.n311 B.n6 10.6151
R468 B.n307 B.n6 10.6151
R469 B.n307 B.n306 10.6151
R470 B.n306 B.n305 10.6151
R471 B.n305 B.n8 10.6151
R472 B.n301 B.n8 10.6151
R473 B.n301 B.n300 10.6151
R474 B.n300 B.n299 10.6151
R475 B.n299 B.n10 10.6151
R476 B.n295 B.n10 10.6151
R477 B.n295 B.n294 10.6151
R478 B.n294 B.n293 10.6151
R479 B.n293 B.n12 10.6151
R480 B.n289 B.n12 10.6151
R481 B.n289 B.n288 10.6151
R482 B.n288 B.n287 10.6151
R483 B.n270 B.n269 6.5566
R484 B.n257 B.n256 6.5566
R485 B.n138 B.n137 6.5566
R486 B.n150 B.n64 6.5566
R487 B.n271 B.n270 4.05904
R488 B.n256 B.n255 4.05904
R489 B.n137 B.n136 4.05904
R490 B.n153 B.n64 4.05904
R491 B.n323 B.n0 2.81026
R492 B.n323 B.n1 2.81026
R493 VP.n0 VP.t1 96.6037
R494 VP.n0 VP.t0 60.6708
R495 VP VP.n0 0.336784
R496 VTAIL.n3 VTAIL.t1 373.493
R497 VTAIL.n0 VTAIL.t2 373.493
R498 VTAIL.n2 VTAIL.t3 373.493
R499 VTAIL.n1 VTAIL.t0 373.493
R500 VTAIL.n1 VTAIL.n0 18.0824
R501 VTAIL.n3 VTAIL.n2 15.7203
R502 VTAIL.n2 VTAIL.n1 1.65136
R503 VTAIL VTAIL.n0 1.11903
R504 VTAIL VTAIL.n3 0.532828
R505 VDD1 VDD1.t1 420.661
R506 VDD1 VDD1.t0 390.82
R507 VN VN.t1 96.7003
R508 VN VN.t0 61.0071
R509 VDD2.n0 VDD2.t1 419.546
R510 VDD2.n0 VDD2.t0 390.171
R511 VDD2 VDD2.n0 0.649207
C0 VN B 0.830406f
C1 VTAIL VP 0.865834f
C2 VN w_n2066_n1198# 2.59327f
C3 VDD2 VP 0.332781f
C4 VN VDD1 0.15556f
C5 VTAIL VDD2 2.18588f
C6 B VP 1.26048f
C7 VTAIL B 1.04056f
C8 VP w_n2066_n1198# 2.8488f
C9 B VDD2 0.854978f
C10 VTAIL w_n2066_n1198# 1.14237f
C11 VDD1 VP 0.669984f
C12 VTAIL VDD1 2.13404f
C13 VDD2 w_n2066_n1198# 1.01653f
C14 VDD1 VDD2 0.650557f
C15 B w_n2066_n1198# 5.60181f
C16 VDD1 B 0.826043f
C17 VDD1 w_n2066_n1198# 0.993923f
C18 VN VP 3.36541f
C19 VTAIL VN 0.851709f
C20 VN VDD2 0.494569f
C21 VDD2 VSUBS 0.513073f
C22 VDD1 VSUBS 2.52186f
C23 VTAIL VSUBS 0.328758f
C24 VN VSUBS 5.45144f
C25 VP VSUBS 1.140724f
C26 B VSUBS 2.69943f
C27 w_n2066_n1198# VSUBS 31.857698f
C28 VDD2.t1 VSUBS 0.148626f
C29 VDD2.t0 VSUBS 0.093179f
C30 VDD2.n0 VSUBS 1.84705f
C31 VN.t0 VSUBS 0.786375f
C32 VN.t1 VSUBS 1.59272f
C33 VDD1.t0 VSUBS 0.08655f
C34 VDD1.t1 VSUBS 0.143152f
C35 VTAIL.t2 VSUBS 0.107575f
C36 VTAIL.n0 VSUBS 1.01646f
C37 VTAIL.t0 VSUBS 0.107575f
C38 VTAIL.n1 VSUBS 1.0567f
C39 VTAIL.t3 VSUBS 0.107575f
C40 VTAIL.n2 VSUBS 0.878152f
C41 VTAIL.t1 VSUBS 0.107575f
C42 VTAIL.n3 VSUBS 0.793603f
C43 VP.t1 VSUBS 1.65798f
C44 VP.t0 VSUBS 0.821811f
C45 VP.n0 VSUBS 3.58578f
C46 B.n0 VSUBS 0.006892f
C47 B.n1 VSUBS 0.006892f
C48 B.n2 VSUBS 0.010899f
C49 B.n3 VSUBS 0.010899f
C50 B.n4 VSUBS 0.010899f
C51 B.n5 VSUBS 0.010899f
C52 B.n6 VSUBS 0.010899f
C53 B.n7 VSUBS 0.010899f
C54 B.n8 VSUBS 0.010899f
C55 B.n9 VSUBS 0.010899f
C56 B.n10 VSUBS 0.010899f
C57 B.n11 VSUBS 0.010899f
C58 B.n12 VSUBS 0.010899f
C59 B.n13 VSUBS 0.010899f
C60 B.n14 VSUBS 0.027417f
C61 B.n15 VSUBS 0.010899f
C62 B.n16 VSUBS 0.010899f
C63 B.n17 VSUBS 0.010899f
C64 B.n18 VSUBS 0.010899f
C65 B.n19 VSUBS 0.010899f
C66 B.t11 VSUBS 0.03374f
C67 B.t10 VSUBS 0.041302f
C68 B.t9 VSUBS 0.219162f
C69 B.n20 VSUBS 0.093213f
C70 B.n21 VSUBS 0.074926f
C71 B.n22 VSUBS 0.010899f
C72 B.n23 VSUBS 0.010899f
C73 B.n24 VSUBS 0.010899f
C74 B.n25 VSUBS 0.010899f
C75 B.t5 VSUBS 0.03374f
C76 B.t4 VSUBS 0.041302f
C77 B.t3 VSUBS 0.219162f
C78 B.n26 VSUBS 0.093213f
C79 B.n27 VSUBS 0.074926f
C80 B.n28 VSUBS 0.010899f
C81 B.n29 VSUBS 0.010899f
C82 B.n30 VSUBS 0.010899f
C83 B.n31 VSUBS 0.010899f
C84 B.n32 VSUBS 0.026209f
C85 B.n33 VSUBS 0.010899f
C86 B.n34 VSUBS 0.010899f
C87 B.n35 VSUBS 0.010899f
C88 B.n36 VSUBS 0.010899f
C89 B.n37 VSUBS 0.010899f
C90 B.n38 VSUBS 0.010899f
C91 B.n39 VSUBS 0.010899f
C92 B.n40 VSUBS 0.010899f
C93 B.n41 VSUBS 0.010899f
C94 B.n42 VSUBS 0.010899f
C95 B.n43 VSUBS 0.010899f
C96 B.n44 VSUBS 0.010899f
C97 B.n45 VSUBS 0.010899f
C98 B.n46 VSUBS 0.010899f
C99 B.n47 VSUBS 0.010899f
C100 B.n48 VSUBS 0.010899f
C101 B.n49 VSUBS 0.010899f
C102 B.n50 VSUBS 0.010899f
C103 B.n51 VSUBS 0.010899f
C104 B.n52 VSUBS 0.010899f
C105 B.n53 VSUBS 0.010899f
C106 B.n54 VSUBS 0.010899f
C107 B.n55 VSUBS 0.010899f
C108 B.n56 VSUBS 0.010899f
C109 B.n57 VSUBS 0.027417f
C110 B.n58 VSUBS 0.010899f
C111 B.n59 VSUBS 0.010899f
C112 B.n60 VSUBS 0.010899f
C113 B.n61 VSUBS 0.010899f
C114 B.t1 VSUBS 0.03374f
C115 B.t2 VSUBS 0.041302f
C116 B.t0 VSUBS 0.219162f
C117 B.n62 VSUBS 0.093213f
C118 B.n63 VSUBS 0.074926f
C119 B.n64 VSUBS 0.025252f
C120 B.n65 VSUBS 0.010899f
C121 B.n66 VSUBS 0.010899f
C122 B.n67 VSUBS 0.010899f
C123 B.n68 VSUBS 0.010899f
C124 B.n69 VSUBS 0.010899f
C125 B.t7 VSUBS 0.03374f
C126 B.t8 VSUBS 0.041302f
C127 B.t6 VSUBS 0.219162f
C128 B.n70 VSUBS 0.093213f
C129 B.n71 VSUBS 0.074926f
C130 B.n72 VSUBS 0.010899f
C131 B.n73 VSUBS 0.010899f
C132 B.n74 VSUBS 0.010899f
C133 B.n75 VSUBS 0.010899f
C134 B.n76 VSUBS 0.025796f
C135 B.n77 VSUBS 0.010899f
C136 B.n78 VSUBS 0.010899f
C137 B.n79 VSUBS 0.010899f
C138 B.n80 VSUBS 0.010899f
C139 B.n81 VSUBS 0.010899f
C140 B.n82 VSUBS 0.010899f
C141 B.n83 VSUBS 0.010899f
C142 B.n84 VSUBS 0.010899f
C143 B.n85 VSUBS 0.010899f
C144 B.n86 VSUBS 0.010899f
C145 B.n87 VSUBS 0.010899f
C146 B.n88 VSUBS 0.010899f
C147 B.n89 VSUBS 0.010899f
C148 B.n90 VSUBS 0.010899f
C149 B.n91 VSUBS 0.010899f
C150 B.n92 VSUBS 0.010899f
C151 B.n93 VSUBS 0.010899f
C152 B.n94 VSUBS 0.010899f
C153 B.n95 VSUBS 0.010899f
C154 B.n96 VSUBS 0.010899f
C155 B.n97 VSUBS 0.010899f
C156 B.n98 VSUBS 0.010899f
C157 B.n99 VSUBS 0.010899f
C158 B.n100 VSUBS 0.010899f
C159 B.n101 VSUBS 0.010899f
C160 B.n102 VSUBS 0.010899f
C161 B.n103 VSUBS 0.010899f
C162 B.n104 VSUBS 0.010899f
C163 B.n105 VSUBS 0.010899f
C164 B.n106 VSUBS 0.010899f
C165 B.n107 VSUBS 0.010899f
C166 B.n108 VSUBS 0.010899f
C167 B.n109 VSUBS 0.010899f
C168 B.n110 VSUBS 0.010899f
C169 B.n111 VSUBS 0.010899f
C170 B.n112 VSUBS 0.010899f
C171 B.n113 VSUBS 0.010899f
C172 B.n114 VSUBS 0.010899f
C173 B.n115 VSUBS 0.010899f
C174 B.n116 VSUBS 0.010899f
C175 B.n117 VSUBS 0.010899f
C176 B.n118 VSUBS 0.010899f
C177 B.n119 VSUBS 0.010899f
C178 B.n120 VSUBS 0.010899f
C179 B.n121 VSUBS 0.025796f
C180 B.n122 VSUBS 0.027417f
C181 B.n123 VSUBS 0.027417f
C182 B.n124 VSUBS 0.010899f
C183 B.n125 VSUBS 0.010899f
C184 B.n126 VSUBS 0.010899f
C185 B.n127 VSUBS 0.010899f
C186 B.n128 VSUBS 0.010899f
C187 B.n129 VSUBS 0.010899f
C188 B.n130 VSUBS 0.010899f
C189 B.n131 VSUBS 0.010899f
C190 B.n132 VSUBS 0.010899f
C191 B.n133 VSUBS 0.010899f
C192 B.n134 VSUBS 0.010899f
C193 B.n135 VSUBS 0.010899f
C194 B.n136 VSUBS 0.007533f
C195 B.n137 VSUBS 0.025252f
C196 B.n138 VSUBS 0.008816f
C197 B.n139 VSUBS 0.010899f
C198 B.n140 VSUBS 0.010899f
C199 B.n141 VSUBS 0.010899f
C200 B.n142 VSUBS 0.010899f
C201 B.n143 VSUBS 0.010899f
C202 B.n144 VSUBS 0.010899f
C203 B.n145 VSUBS 0.010899f
C204 B.n146 VSUBS 0.010899f
C205 B.n147 VSUBS 0.010899f
C206 B.n148 VSUBS 0.010899f
C207 B.n149 VSUBS 0.010899f
C208 B.n150 VSUBS 0.008816f
C209 B.n151 VSUBS 0.010899f
C210 B.n152 VSUBS 0.010899f
C211 B.n153 VSUBS 0.007533f
C212 B.n154 VSUBS 0.010899f
C213 B.n155 VSUBS 0.010899f
C214 B.n156 VSUBS 0.010899f
C215 B.n157 VSUBS 0.010899f
C216 B.n158 VSUBS 0.010899f
C217 B.n159 VSUBS 0.010899f
C218 B.n160 VSUBS 0.010899f
C219 B.n161 VSUBS 0.010899f
C220 B.n162 VSUBS 0.010899f
C221 B.n163 VSUBS 0.010899f
C222 B.n164 VSUBS 0.010899f
C223 B.n165 VSUBS 0.010899f
C224 B.n166 VSUBS 0.027417f
C225 B.n167 VSUBS 0.025796f
C226 B.n168 VSUBS 0.025796f
C227 B.n169 VSUBS 0.010899f
C228 B.n170 VSUBS 0.010899f
C229 B.n171 VSUBS 0.010899f
C230 B.n172 VSUBS 0.010899f
C231 B.n173 VSUBS 0.010899f
C232 B.n174 VSUBS 0.010899f
C233 B.n175 VSUBS 0.010899f
C234 B.n176 VSUBS 0.010899f
C235 B.n177 VSUBS 0.010899f
C236 B.n178 VSUBS 0.010899f
C237 B.n179 VSUBS 0.010899f
C238 B.n180 VSUBS 0.010899f
C239 B.n181 VSUBS 0.010899f
C240 B.n182 VSUBS 0.010899f
C241 B.n183 VSUBS 0.010899f
C242 B.n184 VSUBS 0.010899f
C243 B.n185 VSUBS 0.010899f
C244 B.n186 VSUBS 0.010899f
C245 B.n187 VSUBS 0.010899f
C246 B.n188 VSUBS 0.010899f
C247 B.n189 VSUBS 0.010899f
C248 B.n190 VSUBS 0.010899f
C249 B.n191 VSUBS 0.010899f
C250 B.n192 VSUBS 0.010899f
C251 B.n193 VSUBS 0.010899f
C252 B.n194 VSUBS 0.010899f
C253 B.n195 VSUBS 0.010899f
C254 B.n196 VSUBS 0.010899f
C255 B.n197 VSUBS 0.010899f
C256 B.n198 VSUBS 0.010899f
C257 B.n199 VSUBS 0.010899f
C258 B.n200 VSUBS 0.010899f
C259 B.n201 VSUBS 0.010899f
C260 B.n202 VSUBS 0.010899f
C261 B.n203 VSUBS 0.010899f
C262 B.n204 VSUBS 0.010899f
C263 B.n205 VSUBS 0.010899f
C264 B.n206 VSUBS 0.010899f
C265 B.n207 VSUBS 0.010899f
C266 B.n208 VSUBS 0.010899f
C267 B.n209 VSUBS 0.010899f
C268 B.n210 VSUBS 0.010899f
C269 B.n211 VSUBS 0.010899f
C270 B.n212 VSUBS 0.010899f
C271 B.n213 VSUBS 0.010899f
C272 B.n214 VSUBS 0.010899f
C273 B.n215 VSUBS 0.010899f
C274 B.n216 VSUBS 0.010899f
C275 B.n217 VSUBS 0.010899f
C276 B.n218 VSUBS 0.010899f
C277 B.n219 VSUBS 0.010899f
C278 B.n220 VSUBS 0.010899f
C279 B.n221 VSUBS 0.010899f
C280 B.n222 VSUBS 0.010899f
C281 B.n223 VSUBS 0.010899f
C282 B.n224 VSUBS 0.010899f
C283 B.n225 VSUBS 0.010899f
C284 B.n226 VSUBS 0.010899f
C285 B.n227 VSUBS 0.010899f
C286 B.n228 VSUBS 0.010899f
C287 B.n229 VSUBS 0.010899f
C288 B.n230 VSUBS 0.010899f
C289 B.n231 VSUBS 0.010899f
C290 B.n232 VSUBS 0.010899f
C291 B.n233 VSUBS 0.010899f
C292 B.n234 VSUBS 0.010899f
C293 B.n235 VSUBS 0.010899f
C294 B.n236 VSUBS 0.010899f
C295 B.n237 VSUBS 0.010899f
C296 B.n238 VSUBS 0.010899f
C297 B.n239 VSUBS 0.027005f
C298 B.n240 VSUBS 0.025796f
C299 B.n241 VSUBS 0.027417f
C300 B.n242 VSUBS 0.010899f
C301 B.n243 VSUBS 0.010899f
C302 B.n244 VSUBS 0.010899f
C303 B.n245 VSUBS 0.010899f
C304 B.n246 VSUBS 0.010899f
C305 B.n247 VSUBS 0.010899f
C306 B.n248 VSUBS 0.010899f
C307 B.n249 VSUBS 0.010899f
C308 B.n250 VSUBS 0.010899f
C309 B.n251 VSUBS 0.010899f
C310 B.n252 VSUBS 0.010899f
C311 B.n253 VSUBS 0.010899f
C312 B.n254 VSUBS 0.010899f
C313 B.n255 VSUBS 0.007533f
C314 B.n256 VSUBS 0.025252f
C315 B.n257 VSUBS 0.008816f
C316 B.n258 VSUBS 0.010899f
C317 B.n259 VSUBS 0.010899f
C318 B.n260 VSUBS 0.010899f
C319 B.n261 VSUBS 0.010899f
C320 B.n262 VSUBS 0.010899f
C321 B.n263 VSUBS 0.010899f
C322 B.n264 VSUBS 0.010899f
C323 B.n265 VSUBS 0.010899f
C324 B.n266 VSUBS 0.010899f
C325 B.n267 VSUBS 0.010899f
C326 B.n268 VSUBS 0.010899f
C327 B.n269 VSUBS 0.008816f
C328 B.n270 VSUBS 0.025252f
C329 B.n271 VSUBS 0.007533f
C330 B.n272 VSUBS 0.010899f
C331 B.n273 VSUBS 0.010899f
C332 B.n274 VSUBS 0.010899f
C333 B.n275 VSUBS 0.010899f
C334 B.n276 VSUBS 0.010899f
C335 B.n277 VSUBS 0.010899f
C336 B.n278 VSUBS 0.010899f
C337 B.n279 VSUBS 0.010899f
C338 B.n280 VSUBS 0.010899f
C339 B.n281 VSUBS 0.010899f
C340 B.n282 VSUBS 0.010899f
C341 B.n283 VSUBS 0.010899f
C342 B.n284 VSUBS 0.010899f
C343 B.n285 VSUBS 0.027417f
C344 B.n286 VSUBS 0.025796f
C345 B.n287 VSUBS 0.025796f
C346 B.n288 VSUBS 0.010899f
C347 B.n289 VSUBS 0.010899f
C348 B.n290 VSUBS 0.010899f
C349 B.n291 VSUBS 0.010899f
C350 B.n292 VSUBS 0.010899f
C351 B.n293 VSUBS 0.010899f
C352 B.n294 VSUBS 0.010899f
C353 B.n295 VSUBS 0.010899f
C354 B.n296 VSUBS 0.010899f
C355 B.n297 VSUBS 0.010899f
C356 B.n298 VSUBS 0.010899f
C357 B.n299 VSUBS 0.010899f
C358 B.n300 VSUBS 0.010899f
C359 B.n301 VSUBS 0.010899f
C360 B.n302 VSUBS 0.010899f
C361 B.n303 VSUBS 0.010899f
C362 B.n304 VSUBS 0.010899f
C363 B.n305 VSUBS 0.010899f
C364 B.n306 VSUBS 0.010899f
C365 B.n307 VSUBS 0.010899f
C366 B.n308 VSUBS 0.010899f
C367 B.n309 VSUBS 0.010899f
C368 B.n310 VSUBS 0.010899f
C369 B.n311 VSUBS 0.010899f
C370 B.n312 VSUBS 0.010899f
C371 B.n313 VSUBS 0.010899f
C372 B.n314 VSUBS 0.010899f
C373 B.n315 VSUBS 0.010899f
C374 B.n316 VSUBS 0.010899f
C375 B.n317 VSUBS 0.010899f
C376 B.n318 VSUBS 0.010899f
C377 B.n319 VSUBS 0.010899f
C378 B.n320 VSUBS 0.010899f
C379 B.n321 VSUBS 0.010899f
C380 B.n322 VSUBS 0.010899f
C381 B.n323 VSUBS 0.02468f
.ends

