* NGSPICE file created from diff_pair_sample_0251.ext - technology: sky130A

.subckt diff_pair_sample_0251 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t12 VP.t0 VDD1.t7 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X1 VTAIL.t15 VN.t0 VDD2.t7 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0.1254 ps=1.09 w=0.76 l=3.35
X2 B.t11 B.t9 B.t10 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0 ps=0 w=0.76 l=3.35
X3 VDD1.t2 VP.t1 VTAIL.t11 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X4 VDD2.t6 VN.t1 VTAIL.t4 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X5 VDD1.t0 VP.t2 VTAIL.t10 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.2964 ps=2.3 w=0.76 l=3.35
X6 VDD2.t5 VN.t2 VTAIL.t14 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.2964 ps=2.3 w=0.76 l=3.35
X7 VDD1.t4 VP.t3 VTAIL.t9 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X8 VTAIL.t1 VN.t3 VDD2.t4 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X9 VDD2.t3 VN.t4 VTAIL.t2 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.2964 ps=2.3 w=0.76 l=3.35
X10 VTAIL.t8 VP.t4 VDD1.t3 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X11 VDD1.t1 VP.t5 VTAIL.t7 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.2964 ps=2.3 w=0.76 l=3.35
X12 VTAIL.t3 VN.t5 VDD2.t2 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X13 VTAIL.t6 VP.t6 VDD1.t6 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0.1254 ps=1.09 w=0.76 l=3.35
X14 B.t8 B.t6 B.t7 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0 ps=0 w=0.76 l=3.35
X15 B.t5 B.t3 B.t4 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0 ps=0 w=0.76 l=3.35
X16 VDD2.t1 VN.t6 VTAIL.t13 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.1254 pd=1.09 as=0.1254 ps=1.09 w=0.76 l=3.35
X17 VTAIL.t0 VN.t7 VDD2.t0 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0.1254 ps=1.09 w=0.76 l=3.35
X18 B.t2 B.t0 B.t1 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0 ps=0 w=0.76 l=3.35
X19 VTAIL.t5 VP.t7 VDD1.t5 w_n4650_n1120# sky130_fd_pr__pfet_01v8 ad=0.2964 pd=2.3 as=0.1254 ps=1.09 w=0.76 l=3.35
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n48 VP.n12 76.966
R38 VP.n84 VP.n0 76.966
R39 VP.n47 VP.n13 76.966
R40 VP.n23 VP.n22 70.385
R41 VP.n65 VP.n6 56.5617
R42 VP.n28 VP.n19 56.5617
R43 VP.n56 VP.n10 47.3584
R44 VP.n76 VP.n2 47.3584
R45 VP.n39 VP.n15 47.3584
R46 VP.n48 VP.n47 45.992
R47 VP.n23 VP.t7 38.2121
R48 VP.n52 VP.n10 33.7956
R49 VP.n80 VP.n2 33.7956
R50 VP.n43 VP.n15 33.7956
R51 VP.n51 VP.n50 24.5923
R52 VP.n52 VP.n51 24.5923
R53 VP.n57 VP.n56 24.5923
R54 VP.n59 VP.n57 24.5923
R55 VP.n63 VP.n8 24.5923
R56 VP.n64 VP.n63 24.5923
R57 VP.n65 VP.n64 24.5923
R58 VP.n69 VP.n6 24.5923
R59 VP.n70 VP.n69 24.5923
R60 VP.n71 VP.n70 24.5923
R61 VP.n75 VP.n74 24.5923
R62 VP.n76 VP.n75 24.5923
R63 VP.n81 VP.n80 24.5923
R64 VP.n82 VP.n81 24.5923
R65 VP.n44 VP.n43 24.5923
R66 VP.n45 VP.n44 24.5923
R67 VP.n32 VP.n19 24.5923
R68 VP.n33 VP.n32 24.5923
R69 VP.n34 VP.n33 24.5923
R70 VP.n38 VP.n37 24.5923
R71 VP.n39 VP.n38 24.5923
R72 VP.n26 VP.n21 24.5923
R73 VP.n27 VP.n26 24.5923
R74 VP.n28 VP.n27 24.5923
R75 VP.n59 VP.n58 20.1658
R76 VP.n74 VP.n4 20.1658
R77 VP.n37 VP.n17 20.1658
R78 VP.n50 VP.n12 13.2801
R79 VP.n82 VP.n0 13.2801
R80 VP.n45 VP.n13 13.2801
R81 VP.n12 VP.t6 5.46796
R82 VP.n58 VP.t3 5.46796
R83 VP.n4 VP.t4 5.46796
R84 VP.n0 VP.t5 5.46796
R85 VP.n13 VP.t2 5.46796
R86 VP.n17 VP.t0 5.46796
R87 VP.n22 VP.t1 5.46796
R88 VP.n58 VP.n8 4.42703
R89 VP.n71 VP.n4 4.42703
R90 VP.n34 VP.n17 4.42703
R91 VP.n22 VP.n21 4.42703
R92 VP.n24 VP.n23 4.22517
R93 VP.n47 VP.n46 0.354861
R94 VP.n49 VP.n48 0.354861
R95 VP.n84 VP.n83 0.354861
R96 VP VP.n84 0.267071
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VDD1 VDD1.n0 638.611
R133 VDD1.n3 VDD1.n2 638.497
R134 VDD1.n3 VDD1.n1 638.497
R135 VDD1.n5 VDD1.n4 636.967
R136 VDD1.n4 VDD1.t7 42.7702
R137 VDD1.n4 VDD1.t0 42.7702
R138 VDD1.n0 VDD1.t5 42.7702
R139 VDD1.n0 VDD1.t2 42.7702
R140 VDD1.n2 VDD1.t3 42.7702
R141 VDD1.n2 VDD1.t1 42.7702
R142 VDD1.n1 VDD1.t6 42.7702
R143 VDD1.n1 VDD1.t4 42.7702
R144 VDD1.n5 VDD1.n3 39.2293
R145 VDD1 VDD1.n5 1.52852
R146 VTAIL.n15 VTAIL.t14 663.058
R147 VTAIL.n2 VTAIL.t0 663.058
R148 VTAIL.n3 VTAIL.t7 663.058
R149 VTAIL.n6 VTAIL.t6 663.058
R150 VTAIL.n14 VTAIL.t10 663.058
R151 VTAIL.n11 VTAIL.t5 663.058
R152 VTAIL.n10 VTAIL.t2 663.058
R153 VTAIL.n7 VTAIL.t15 663.058
R154 VTAIL.n1 VTAIL.n0 620.288
R155 VTAIL.n5 VTAIL.n4 620.288
R156 VTAIL.n13 VTAIL.n12 620.288
R157 VTAIL.n9 VTAIL.n8 620.288
R158 VTAIL.n0 VTAIL.t13 42.7702
R159 VTAIL.n0 VTAIL.t1 42.7702
R160 VTAIL.n4 VTAIL.t9 42.7702
R161 VTAIL.n4 VTAIL.t8 42.7702
R162 VTAIL.n12 VTAIL.t11 42.7702
R163 VTAIL.n12 VTAIL.t12 42.7702
R164 VTAIL.n8 VTAIL.t4 42.7702
R165 VTAIL.n8 VTAIL.t3 42.7702
R166 VTAIL.n15 VTAIL.n14 16.1945
R167 VTAIL.n7 VTAIL.n6 16.1945
R168 VTAIL.n9 VTAIL.n7 3.17291
R169 VTAIL.n10 VTAIL.n9 3.17291
R170 VTAIL.n13 VTAIL.n11 3.17291
R171 VTAIL.n14 VTAIL.n13 3.17291
R172 VTAIL.n6 VTAIL.n5 3.17291
R173 VTAIL.n5 VTAIL.n3 3.17291
R174 VTAIL.n2 VTAIL.n1 3.17291
R175 VTAIL VTAIL.n15 3.11472
R176 VTAIL.n11 VTAIL.n10 0.470328
R177 VTAIL.n3 VTAIL.n2 0.470328
R178 VTAIL VTAIL.n1 0.0586897
R179 VN.n68 VN.n67 161.3
R180 VN.n66 VN.n36 161.3
R181 VN.n65 VN.n64 161.3
R182 VN.n63 VN.n37 161.3
R183 VN.n62 VN.n61 161.3
R184 VN.n60 VN.n38 161.3
R185 VN.n59 VN.n58 161.3
R186 VN.n57 VN.n56 161.3
R187 VN.n55 VN.n40 161.3
R188 VN.n54 VN.n53 161.3
R189 VN.n52 VN.n41 161.3
R190 VN.n51 VN.n50 161.3
R191 VN.n49 VN.n42 161.3
R192 VN.n48 VN.n47 161.3
R193 VN.n46 VN.n43 161.3
R194 VN.n33 VN.n32 161.3
R195 VN.n31 VN.n1 161.3
R196 VN.n30 VN.n29 161.3
R197 VN.n28 VN.n2 161.3
R198 VN.n27 VN.n26 161.3
R199 VN.n25 VN.n3 161.3
R200 VN.n24 VN.n23 161.3
R201 VN.n22 VN.n21 161.3
R202 VN.n20 VN.n5 161.3
R203 VN.n19 VN.n18 161.3
R204 VN.n17 VN.n6 161.3
R205 VN.n16 VN.n15 161.3
R206 VN.n14 VN.n7 161.3
R207 VN.n13 VN.n12 161.3
R208 VN.n11 VN.n8 161.3
R209 VN.n34 VN.n0 76.966
R210 VN.n69 VN.n35 76.966
R211 VN.n10 VN.n9 70.385
R212 VN.n45 VN.n44 70.385
R213 VN.n15 VN.n6 56.5617
R214 VN.n50 VN.n41 56.5617
R215 VN.n26 VN.n2 47.3584
R216 VN.n61 VN.n37 47.3584
R217 VN VN.n69 46.1572
R218 VN.n45 VN.t4 38.2123
R219 VN.n10 VN.t7 38.2123
R220 VN.n30 VN.n2 33.7956
R221 VN.n65 VN.n37 33.7956
R222 VN.n13 VN.n8 24.5923
R223 VN.n14 VN.n13 24.5923
R224 VN.n15 VN.n14 24.5923
R225 VN.n19 VN.n6 24.5923
R226 VN.n20 VN.n19 24.5923
R227 VN.n21 VN.n20 24.5923
R228 VN.n25 VN.n24 24.5923
R229 VN.n26 VN.n25 24.5923
R230 VN.n31 VN.n30 24.5923
R231 VN.n32 VN.n31 24.5923
R232 VN.n50 VN.n49 24.5923
R233 VN.n49 VN.n48 24.5923
R234 VN.n48 VN.n43 24.5923
R235 VN.n61 VN.n60 24.5923
R236 VN.n60 VN.n59 24.5923
R237 VN.n56 VN.n55 24.5923
R238 VN.n55 VN.n54 24.5923
R239 VN.n54 VN.n41 24.5923
R240 VN.n67 VN.n66 24.5923
R241 VN.n66 VN.n65 24.5923
R242 VN.n24 VN.n4 20.1658
R243 VN.n59 VN.n39 20.1658
R244 VN.n32 VN.n0 13.2801
R245 VN.n67 VN.n35 13.2801
R246 VN.n9 VN.t6 5.46796
R247 VN.n4 VN.t3 5.46796
R248 VN.n0 VN.t2 5.46796
R249 VN.n44 VN.t5 5.46796
R250 VN.n39 VN.t1 5.46796
R251 VN.n35 VN.t0 5.46796
R252 VN.n9 VN.n8 4.42703
R253 VN.n21 VN.n4 4.42703
R254 VN.n44 VN.n43 4.42703
R255 VN.n56 VN.n39 4.42703
R256 VN.n46 VN.n45 4.22519
R257 VN.n11 VN.n10 4.22519
R258 VN.n69 VN.n68 0.354861
R259 VN.n34 VN.n33 0.354861
R260 VN VN.n34 0.267071
R261 VN.n68 VN.n36 0.189894
R262 VN.n64 VN.n36 0.189894
R263 VN.n64 VN.n63 0.189894
R264 VN.n63 VN.n62 0.189894
R265 VN.n62 VN.n38 0.189894
R266 VN.n58 VN.n38 0.189894
R267 VN.n58 VN.n57 0.189894
R268 VN.n57 VN.n40 0.189894
R269 VN.n53 VN.n40 0.189894
R270 VN.n53 VN.n52 0.189894
R271 VN.n52 VN.n51 0.189894
R272 VN.n51 VN.n42 0.189894
R273 VN.n47 VN.n42 0.189894
R274 VN.n47 VN.n46 0.189894
R275 VN.n12 VN.n11 0.189894
R276 VN.n12 VN.n7 0.189894
R277 VN.n16 VN.n7 0.189894
R278 VN.n17 VN.n16 0.189894
R279 VN.n18 VN.n17 0.189894
R280 VN.n18 VN.n5 0.189894
R281 VN.n22 VN.n5 0.189894
R282 VN.n23 VN.n22 0.189894
R283 VN.n23 VN.n3 0.189894
R284 VN.n27 VN.n3 0.189894
R285 VN.n28 VN.n27 0.189894
R286 VN.n29 VN.n28 0.189894
R287 VN.n29 VN.n1 0.189894
R288 VN.n33 VN.n1 0.189894
R289 VDD2.n2 VDD2.n1 638.497
R290 VDD2.n2 VDD2.n0 638.497
R291 VDD2 VDD2.n5 638.495
R292 VDD2.n4 VDD2.n3 636.967
R293 VDD2.n5 VDD2.t2 42.7702
R294 VDD2.n5 VDD2.t3 42.7702
R295 VDD2.n3 VDD2.t7 42.7702
R296 VDD2.n3 VDD2.t6 42.7702
R297 VDD2.n1 VDD2.t4 42.7702
R298 VDD2.n1 VDD2.t5 42.7702
R299 VDD2.n0 VDD2.t0 42.7702
R300 VDD2.n0 VDD2.t1 42.7702
R301 VDD2.n4 VDD2.n2 38.6463
R302 VDD2 VDD2.n4 1.6449
R303 B.n118 B.t11 723.577
R304 B.n126 B.t5 723.577
R305 B.n38 B.t1 723.577
R306 B.n44 B.t7 723.577
R307 B.n119 B.t10 652.207
R308 B.n127 B.t4 652.207
R309 B.n39 B.t2 652.207
R310 B.n45 B.t8 652.207
R311 B.n484 B.n483 585
R312 B.n485 B.n50 585
R313 B.n487 B.n486 585
R314 B.n488 B.n49 585
R315 B.n490 B.n489 585
R316 B.n491 B.n48 585
R317 B.n493 B.n492 585
R318 B.n494 B.n47 585
R319 B.n496 B.n495 585
R320 B.n498 B.n497 585
R321 B.n499 B.n43 585
R322 B.n501 B.n500 585
R323 B.n502 B.n42 585
R324 B.n504 B.n503 585
R325 B.n505 B.n41 585
R326 B.n507 B.n506 585
R327 B.n508 B.n40 585
R328 B.n510 B.n509 585
R329 B.n512 B.n37 585
R330 B.n514 B.n513 585
R331 B.n515 B.n36 585
R332 B.n517 B.n516 585
R333 B.n518 B.n35 585
R334 B.n520 B.n519 585
R335 B.n521 B.n34 585
R336 B.n523 B.n522 585
R337 B.n524 B.n33 585
R338 B.n482 B.n51 585
R339 B.n481 B.n480 585
R340 B.n479 B.n52 585
R341 B.n478 B.n477 585
R342 B.n476 B.n53 585
R343 B.n475 B.n474 585
R344 B.n473 B.n54 585
R345 B.n472 B.n471 585
R346 B.n470 B.n55 585
R347 B.n469 B.n468 585
R348 B.n467 B.n56 585
R349 B.n466 B.n465 585
R350 B.n464 B.n57 585
R351 B.n463 B.n462 585
R352 B.n461 B.n58 585
R353 B.n460 B.n459 585
R354 B.n458 B.n59 585
R355 B.n457 B.n456 585
R356 B.n455 B.n60 585
R357 B.n454 B.n453 585
R358 B.n452 B.n61 585
R359 B.n451 B.n450 585
R360 B.n449 B.n62 585
R361 B.n448 B.n447 585
R362 B.n446 B.n63 585
R363 B.n445 B.n444 585
R364 B.n443 B.n64 585
R365 B.n442 B.n441 585
R366 B.n440 B.n65 585
R367 B.n439 B.n438 585
R368 B.n437 B.n66 585
R369 B.n436 B.n435 585
R370 B.n434 B.n67 585
R371 B.n433 B.n432 585
R372 B.n431 B.n68 585
R373 B.n430 B.n429 585
R374 B.n428 B.n69 585
R375 B.n427 B.n426 585
R376 B.n425 B.n70 585
R377 B.n424 B.n423 585
R378 B.n422 B.n71 585
R379 B.n421 B.n420 585
R380 B.n419 B.n72 585
R381 B.n418 B.n417 585
R382 B.n416 B.n73 585
R383 B.n415 B.n414 585
R384 B.n413 B.n74 585
R385 B.n412 B.n411 585
R386 B.n410 B.n75 585
R387 B.n409 B.n408 585
R388 B.n407 B.n76 585
R389 B.n406 B.n405 585
R390 B.n404 B.n77 585
R391 B.n403 B.n402 585
R392 B.n401 B.n78 585
R393 B.n400 B.n399 585
R394 B.n398 B.n79 585
R395 B.n397 B.n396 585
R396 B.n395 B.n80 585
R397 B.n394 B.n393 585
R398 B.n392 B.n81 585
R399 B.n391 B.n390 585
R400 B.n389 B.n82 585
R401 B.n388 B.n387 585
R402 B.n386 B.n83 585
R403 B.n385 B.n384 585
R404 B.n383 B.n84 585
R405 B.n382 B.n381 585
R406 B.n380 B.n85 585
R407 B.n379 B.n378 585
R408 B.n377 B.n86 585
R409 B.n376 B.n375 585
R410 B.n374 B.n87 585
R411 B.n373 B.n372 585
R412 B.n371 B.n88 585
R413 B.n370 B.n369 585
R414 B.n368 B.n89 585
R415 B.n367 B.n366 585
R416 B.n365 B.n90 585
R417 B.n364 B.n363 585
R418 B.n362 B.n91 585
R419 B.n361 B.n360 585
R420 B.n359 B.n92 585
R421 B.n358 B.n357 585
R422 B.n356 B.n93 585
R423 B.n355 B.n354 585
R424 B.n353 B.n94 585
R425 B.n352 B.n351 585
R426 B.n350 B.n95 585
R427 B.n349 B.n348 585
R428 B.n347 B.n96 585
R429 B.n346 B.n345 585
R430 B.n344 B.n97 585
R431 B.n343 B.n342 585
R432 B.n341 B.n98 585
R433 B.n340 B.n339 585
R434 B.n338 B.n99 585
R435 B.n337 B.n336 585
R436 B.n335 B.n100 585
R437 B.n334 B.n333 585
R438 B.n332 B.n101 585
R439 B.n331 B.n330 585
R440 B.n329 B.n102 585
R441 B.n328 B.n327 585
R442 B.n326 B.n103 585
R443 B.n325 B.n324 585
R444 B.n323 B.n104 585
R445 B.n322 B.n321 585
R446 B.n320 B.n105 585
R447 B.n319 B.n318 585
R448 B.n317 B.n106 585
R449 B.n316 B.n315 585
R450 B.n314 B.n107 585
R451 B.n313 B.n312 585
R452 B.n311 B.n108 585
R453 B.n310 B.n309 585
R454 B.n308 B.n109 585
R455 B.n307 B.n306 585
R456 B.n305 B.n110 585
R457 B.n304 B.n303 585
R458 B.n302 B.n111 585
R459 B.n301 B.n300 585
R460 B.n299 B.n112 585
R461 B.n298 B.n297 585
R462 B.n296 B.n113 585
R463 B.n254 B.n131 585
R464 B.n256 B.n255 585
R465 B.n257 B.n130 585
R466 B.n259 B.n258 585
R467 B.n260 B.n129 585
R468 B.n262 B.n261 585
R469 B.n263 B.n128 585
R470 B.n265 B.n264 585
R471 B.n266 B.n125 585
R472 B.n269 B.n268 585
R473 B.n270 B.n124 585
R474 B.n272 B.n271 585
R475 B.n273 B.n123 585
R476 B.n275 B.n274 585
R477 B.n276 B.n122 585
R478 B.n278 B.n277 585
R479 B.n279 B.n121 585
R480 B.n281 B.n280 585
R481 B.n283 B.n282 585
R482 B.n284 B.n117 585
R483 B.n286 B.n285 585
R484 B.n287 B.n116 585
R485 B.n289 B.n288 585
R486 B.n290 B.n115 585
R487 B.n292 B.n291 585
R488 B.n293 B.n114 585
R489 B.n295 B.n294 585
R490 B.n253 B.n252 585
R491 B.n251 B.n132 585
R492 B.n250 B.n249 585
R493 B.n248 B.n133 585
R494 B.n247 B.n246 585
R495 B.n245 B.n134 585
R496 B.n244 B.n243 585
R497 B.n242 B.n135 585
R498 B.n241 B.n240 585
R499 B.n239 B.n136 585
R500 B.n238 B.n237 585
R501 B.n236 B.n137 585
R502 B.n235 B.n234 585
R503 B.n233 B.n138 585
R504 B.n232 B.n231 585
R505 B.n230 B.n139 585
R506 B.n229 B.n228 585
R507 B.n227 B.n140 585
R508 B.n226 B.n225 585
R509 B.n224 B.n141 585
R510 B.n223 B.n222 585
R511 B.n221 B.n142 585
R512 B.n220 B.n219 585
R513 B.n218 B.n143 585
R514 B.n217 B.n216 585
R515 B.n215 B.n144 585
R516 B.n214 B.n213 585
R517 B.n212 B.n145 585
R518 B.n211 B.n210 585
R519 B.n209 B.n146 585
R520 B.n208 B.n207 585
R521 B.n206 B.n147 585
R522 B.n205 B.n204 585
R523 B.n203 B.n148 585
R524 B.n202 B.n201 585
R525 B.n200 B.n149 585
R526 B.n199 B.n198 585
R527 B.n197 B.n150 585
R528 B.n196 B.n195 585
R529 B.n194 B.n151 585
R530 B.n193 B.n192 585
R531 B.n191 B.n152 585
R532 B.n190 B.n189 585
R533 B.n188 B.n153 585
R534 B.n187 B.n186 585
R535 B.n185 B.n154 585
R536 B.n184 B.n183 585
R537 B.n182 B.n155 585
R538 B.n181 B.n180 585
R539 B.n179 B.n156 585
R540 B.n178 B.n177 585
R541 B.n176 B.n157 585
R542 B.n175 B.n174 585
R543 B.n173 B.n158 585
R544 B.n172 B.n171 585
R545 B.n170 B.n159 585
R546 B.n169 B.n168 585
R547 B.n167 B.n160 585
R548 B.n166 B.n165 585
R549 B.n164 B.n161 585
R550 B.n163 B.n162 585
R551 B.n2 B.n0 585
R552 B.n617 B.n1 585
R553 B.n616 B.n615 585
R554 B.n614 B.n3 585
R555 B.n613 B.n612 585
R556 B.n611 B.n4 585
R557 B.n610 B.n609 585
R558 B.n608 B.n5 585
R559 B.n607 B.n606 585
R560 B.n605 B.n6 585
R561 B.n604 B.n603 585
R562 B.n602 B.n7 585
R563 B.n601 B.n600 585
R564 B.n599 B.n8 585
R565 B.n598 B.n597 585
R566 B.n596 B.n9 585
R567 B.n595 B.n594 585
R568 B.n593 B.n10 585
R569 B.n592 B.n591 585
R570 B.n590 B.n11 585
R571 B.n589 B.n588 585
R572 B.n587 B.n12 585
R573 B.n586 B.n585 585
R574 B.n584 B.n13 585
R575 B.n583 B.n582 585
R576 B.n581 B.n14 585
R577 B.n580 B.n579 585
R578 B.n578 B.n15 585
R579 B.n577 B.n576 585
R580 B.n575 B.n16 585
R581 B.n574 B.n573 585
R582 B.n572 B.n17 585
R583 B.n571 B.n570 585
R584 B.n569 B.n18 585
R585 B.n568 B.n567 585
R586 B.n566 B.n19 585
R587 B.n565 B.n564 585
R588 B.n563 B.n20 585
R589 B.n562 B.n561 585
R590 B.n560 B.n21 585
R591 B.n559 B.n558 585
R592 B.n557 B.n22 585
R593 B.n556 B.n555 585
R594 B.n554 B.n23 585
R595 B.n553 B.n552 585
R596 B.n551 B.n24 585
R597 B.n550 B.n549 585
R598 B.n548 B.n25 585
R599 B.n547 B.n546 585
R600 B.n545 B.n26 585
R601 B.n544 B.n543 585
R602 B.n542 B.n27 585
R603 B.n541 B.n540 585
R604 B.n539 B.n28 585
R605 B.n538 B.n537 585
R606 B.n536 B.n29 585
R607 B.n535 B.n534 585
R608 B.n533 B.n30 585
R609 B.n532 B.n531 585
R610 B.n530 B.n31 585
R611 B.n529 B.n528 585
R612 B.n527 B.n32 585
R613 B.n526 B.n525 585
R614 B.n619 B.n618 585
R615 B.n252 B.n131 511.721
R616 B.n526 B.n33 511.721
R617 B.n294 B.n113 511.721
R618 B.n484 B.n51 511.721
R619 B.n118 B.t9 209.843
R620 B.n126 B.t3 209.843
R621 B.n38 B.t0 209.843
R622 B.n44 B.t6 209.843
R623 B.n252 B.n251 163.367
R624 B.n251 B.n250 163.367
R625 B.n250 B.n133 163.367
R626 B.n246 B.n133 163.367
R627 B.n246 B.n245 163.367
R628 B.n245 B.n244 163.367
R629 B.n244 B.n135 163.367
R630 B.n240 B.n135 163.367
R631 B.n240 B.n239 163.367
R632 B.n239 B.n238 163.367
R633 B.n238 B.n137 163.367
R634 B.n234 B.n137 163.367
R635 B.n234 B.n233 163.367
R636 B.n233 B.n232 163.367
R637 B.n232 B.n139 163.367
R638 B.n228 B.n139 163.367
R639 B.n228 B.n227 163.367
R640 B.n227 B.n226 163.367
R641 B.n226 B.n141 163.367
R642 B.n222 B.n141 163.367
R643 B.n222 B.n221 163.367
R644 B.n221 B.n220 163.367
R645 B.n220 B.n143 163.367
R646 B.n216 B.n143 163.367
R647 B.n216 B.n215 163.367
R648 B.n215 B.n214 163.367
R649 B.n214 B.n145 163.367
R650 B.n210 B.n145 163.367
R651 B.n210 B.n209 163.367
R652 B.n209 B.n208 163.367
R653 B.n208 B.n147 163.367
R654 B.n204 B.n147 163.367
R655 B.n204 B.n203 163.367
R656 B.n203 B.n202 163.367
R657 B.n202 B.n149 163.367
R658 B.n198 B.n149 163.367
R659 B.n198 B.n197 163.367
R660 B.n197 B.n196 163.367
R661 B.n196 B.n151 163.367
R662 B.n192 B.n151 163.367
R663 B.n192 B.n191 163.367
R664 B.n191 B.n190 163.367
R665 B.n190 B.n153 163.367
R666 B.n186 B.n153 163.367
R667 B.n186 B.n185 163.367
R668 B.n185 B.n184 163.367
R669 B.n184 B.n155 163.367
R670 B.n180 B.n155 163.367
R671 B.n180 B.n179 163.367
R672 B.n179 B.n178 163.367
R673 B.n178 B.n157 163.367
R674 B.n174 B.n157 163.367
R675 B.n174 B.n173 163.367
R676 B.n173 B.n172 163.367
R677 B.n172 B.n159 163.367
R678 B.n168 B.n159 163.367
R679 B.n168 B.n167 163.367
R680 B.n167 B.n166 163.367
R681 B.n166 B.n161 163.367
R682 B.n162 B.n161 163.367
R683 B.n162 B.n2 163.367
R684 B.n618 B.n2 163.367
R685 B.n618 B.n617 163.367
R686 B.n617 B.n616 163.367
R687 B.n616 B.n3 163.367
R688 B.n612 B.n3 163.367
R689 B.n612 B.n611 163.367
R690 B.n611 B.n610 163.367
R691 B.n610 B.n5 163.367
R692 B.n606 B.n5 163.367
R693 B.n606 B.n605 163.367
R694 B.n605 B.n604 163.367
R695 B.n604 B.n7 163.367
R696 B.n600 B.n7 163.367
R697 B.n600 B.n599 163.367
R698 B.n599 B.n598 163.367
R699 B.n598 B.n9 163.367
R700 B.n594 B.n9 163.367
R701 B.n594 B.n593 163.367
R702 B.n593 B.n592 163.367
R703 B.n592 B.n11 163.367
R704 B.n588 B.n11 163.367
R705 B.n588 B.n587 163.367
R706 B.n587 B.n586 163.367
R707 B.n586 B.n13 163.367
R708 B.n582 B.n13 163.367
R709 B.n582 B.n581 163.367
R710 B.n581 B.n580 163.367
R711 B.n580 B.n15 163.367
R712 B.n576 B.n15 163.367
R713 B.n576 B.n575 163.367
R714 B.n575 B.n574 163.367
R715 B.n574 B.n17 163.367
R716 B.n570 B.n17 163.367
R717 B.n570 B.n569 163.367
R718 B.n569 B.n568 163.367
R719 B.n568 B.n19 163.367
R720 B.n564 B.n19 163.367
R721 B.n564 B.n563 163.367
R722 B.n563 B.n562 163.367
R723 B.n562 B.n21 163.367
R724 B.n558 B.n21 163.367
R725 B.n558 B.n557 163.367
R726 B.n557 B.n556 163.367
R727 B.n556 B.n23 163.367
R728 B.n552 B.n23 163.367
R729 B.n552 B.n551 163.367
R730 B.n551 B.n550 163.367
R731 B.n550 B.n25 163.367
R732 B.n546 B.n25 163.367
R733 B.n546 B.n545 163.367
R734 B.n545 B.n544 163.367
R735 B.n544 B.n27 163.367
R736 B.n540 B.n27 163.367
R737 B.n540 B.n539 163.367
R738 B.n539 B.n538 163.367
R739 B.n538 B.n29 163.367
R740 B.n534 B.n29 163.367
R741 B.n534 B.n533 163.367
R742 B.n533 B.n532 163.367
R743 B.n532 B.n31 163.367
R744 B.n528 B.n31 163.367
R745 B.n528 B.n527 163.367
R746 B.n527 B.n526 163.367
R747 B.n256 B.n131 163.367
R748 B.n257 B.n256 163.367
R749 B.n258 B.n257 163.367
R750 B.n258 B.n129 163.367
R751 B.n262 B.n129 163.367
R752 B.n263 B.n262 163.367
R753 B.n264 B.n263 163.367
R754 B.n264 B.n125 163.367
R755 B.n269 B.n125 163.367
R756 B.n270 B.n269 163.367
R757 B.n271 B.n270 163.367
R758 B.n271 B.n123 163.367
R759 B.n275 B.n123 163.367
R760 B.n276 B.n275 163.367
R761 B.n277 B.n276 163.367
R762 B.n277 B.n121 163.367
R763 B.n281 B.n121 163.367
R764 B.n282 B.n281 163.367
R765 B.n282 B.n117 163.367
R766 B.n286 B.n117 163.367
R767 B.n287 B.n286 163.367
R768 B.n288 B.n287 163.367
R769 B.n288 B.n115 163.367
R770 B.n292 B.n115 163.367
R771 B.n293 B.n292 163.367
R772 B.n294 B.n293 163.367
R773 B.n298 B.n113 163.367
R774 B.n299 B.n298 163.367
R775 B.n300 B.n299 163.367
R776 B.n300 B.n111 163.367
R777 B.n304 B.n111 163.367
R778 B.n305 B.n304 163.367
R779 B.n306 B.n305 163.367
R780 B.n306 B.n109 163.367
R781 B.n310 B.n109 163.367
R782 B.n311 B.n310 163.367
R783 B.n312 B.n311 163.367
R784 B.n312 B.n107 163.367
R785 B.n316 B.n107 163.367
R786 B.n317 B.n316 163.367
R787 B.n318 B.n317 163.367
R788 B.n318 B.n105 163.367
R789 B.n322 B.n105 163.367
R790 B.n323 B.n322 163.367
R791 B.n324 B.n323 163.367
R792 B.n324 B.n103 163.367
R793 B.n328 B.n103 163.367
R794 B.n329 B.n328 163.367
R795 B.n330 B.n329 163.367
R796 B.n330 B.n101 163.367
R797 B.n334 B.n101 163.367
R798 B.n335 B.n334 163.367
R799 B.n336 B.n335 163.367
R800 B.n336 B.n99 163.367
R801 B.n340 B.n99 163.367
R802 B.n341 B.n340 163.367
R803 B.n342 B.n341 163.367
R804 B.n342 B.n97 163.367
R805 B.n346 B.n97 163.367
R806 B.n347 B.n346 163.367
R807 B.n348 B.n347 163.367
R808 B.n348 B.n95 163.367
R809 B.n352 B.n95 163.367
R810 B.n353 B.n352 163.367
R811 B.n354 B.n353 163.367
R812 B.n354 B.n93 163.367
R813 B.n358 B.n93 163.367
R814 B.n359 B.n358 163.367
R815 B.n360 B.n359 163.367
R816 B.n360 B.n91 163.367
R817 B.n364 B.n91 163.367
R818 B.n365 B.n364 163.367
R819 B.n366 B.n365 163.367
R820 B.n366 B.n89 163.367
R821 B.n370 B.n89 163.367
R822 B.n371 B.n370 163.367
R823 B.n372 B.n371 163.367
R824 B.n372 B.n87 163.367
R825 B.n376 B.n87 163.367
R826 B.n377 B.n376 163.367
R827 B.n378 B.n377 163.367
R828 B.n378 B.n85 163.367
R829 B.n382 B.n85 163.367
R830 B.n383 B.n382 163.367
R831 B.n384 B.n383 163.367
R832 B.n384 B.n83 163.367
R833 B.n388 B.n83 163.367
R834 B.n389 B.n388 163.367
R835 B.n390 B.n389 163.367
R836 B.n390 B.n81 163.367
R837 B.n394 B.n81 163.367
R838 B.n395 B.n394 163.367
R839 B.n396 B.n395 163.367
R840 B.n396 B.n79 163.367
R841 B.n400 B.n79 163.367
R842 B.n401 B.n400 163.367
R843 B.n402 B.n401 163.367
R844 B.n402 B.n77 163.367
R845 B.n406 B.n77 163.367
R846 B.n407 B.n406 163.367
R847 B.n408 B.n407 163.367
R848 B.n408 B.n75 163.367
R849 B.n412 B.n75 163.367
R850 B.n413 B.n412 163.367
R851 B.n414 B.n413 163.367
R852 B.n414 B.n73 163.367
R853 B.n418 B.n73 163.367
R854 B.n419 B.n418 163.367
R855 B.n420 B.n419 163.367
R856 B.n420 B.n71 163.367
R857 B.n424 B.n71 163.367
R858 B.n425 B.n424 163.367
R859 B.n426 B.n425 163.367
R860 B.n426 B.n69 163.367
R861 B.n430 B.n69 163.367
R862 B.n431 B.n430 163.367
R863 B.n432 B.n431 163.367
R864 B.n432 B.n67 163.367
R865 B.n436 B.n67 163.367
R866 B.n437 B.n436 163.367
R867 B.n438 B.n437 163.367
R868 B.n438 B.n65 163.367
R869 B.n442 B.n65 163.367
R870 B.n443 B.n442 163.367
R871 B.n444 B.n443 163.367
R872 B.n444 B.n63 163.367
R873 B.n448 B.n63 163.367
R874 B.n449 B.n448 163.367
R875 B.n450 B.n449 163.367
R876 B.n450 B.n61 163.367
R877 B.n454 B.n61 163.367
R878 B.n455 B.n454 163.367
R879 B.n456 B.n455 163.367
R880 B.n456 B.n59 163.367
R881 B.n460 B.n59 163.367
R882 B.n461 B.n460 163.367
R883 B.n462 B.n461 163.367
R884 B.n462 B.n57 163.367
R885 B.n466 B.n57 163.367
R886 B.n467 B.n466 163.367
R887 B.n468 B.n467 163.367
R888 B.n468 B.n55 163.367
R889 B.n472 B.n55 163.367
R890 B.n473 B.n472 163.367
R891 B.n474 B.n473 163.367
R892 B.n474 B.n53 163.367
R893 B.n478 B.n53 163.367
R894 B.n479 B.n478 163.367
R895 B.n480 B.n479 163.367
R896 B.n480 B.n51 163.367
R897 B.n522 B.n33 163.367
R898 B.n522 B.n521 163.367
R899 B.n521 B.n520 163.367
R900 B.n520 B.n35 163.367
R901 B.n516 B.n35 163.367
R902 B.n516 B.n515 163.367
R903 B.n515 B.n514 163.367
R904 B.n514 B.n37 163.367
R905 B.n509 B.n37 163.367
R906 B.n509 B.n508 163.367
R907 B.n508 B.n507 163.367
R908 B.n507 B.n41 163.367
R909 B.n503 B.n41 163.367
R910 B.n503 B.n502 163.367
R911 B.n502 B.n501 163.367
R912 B.n501 B.n43 163.367
R913 B.n497 B.n43 163.367
R914 B.n497 B.n496 163.367
R915 B.n496 B.n47 163.367
R916 B.n492 B.n47 163.367
R917 B.n492 B.n491 163.367
R918 B.n491 B.n490 163.367
R919 B.n490 B.n49 163.367
R920 B.n486 B.n49 163.367
R921 B.n486 B.n485 163.367
R922 B.n485 B.n484 163.367
R923 B.n119 B.n118 71.3702
R924 B.n127 B.n126 71.3702
R925 B.n39 B.n38 71.3702
R926 B.n45 B.n44 71.3702
R927 B.n120 B.n119 59.5399
R928 B.n267 B.n127 59.5399
R929 B.n511 B.n39 59.5399
R930 B.n46 B.n45 59.5399
R931 B.n525 B.n524 33.2493
R932 B.n483 B.n482 33.2493
R933 B.n296 B.n295 33.2493
R934 B.n254 B.n253 33.2493
R935 B B.n619 18.0485
R936 B.n524 B.n523 10.6151
R937 B.n523 B.n34 10.6151
R938 B.n519 B.n34 10.6151
R939 B.n519 B.n518 10.6151
R940 B.n518 B.n517 10.6151
R941 B.n517 B.n36 10.6151
R942 B.n513 B.n36 10.6151
R943 B.n513 B.n512 10.6151
R944 B.n510 B.n40 10.6151
R945 B.n506 B.n40 10.6151
R946 B.n506 B.n505 10.6151
R947 B.n505 B.n504 10.6151
R948 B.n504 B.n42 10.6151
R949 B.n500 B.n42 10.6151
R950 B.n500 B.n499 10.6151
R951 B.n499 B.n498 10.6151
R952 B.n495 B.n494 10.6151
R953 B.n494 B.n493 10.6151
R954 B.n493 B.n48 10.6151
R955 B.n489 B.n48 10.6151
R956 B.n489 B.n488 10.6151
R957 B.n488 B.n487 10.6151
R958 B.n487 B.n50 10.6151
R959 B.n483 B.n50 10.6151
R960 B.n297 B.n296 10.6151
R961 B.n297 B.n112 10.6151
R962 B.n301 B.n112 10.6151
R963 B.n302 B.n301 10.6151
R964 B.n303 B.n302 10.6151
R965 B.n303 B.n110 10.6151
R966 B.n307 B.n110 10.6151
R967 B.n308 B.n307 10.6151
R968 B.n309 B.n308 10.6151
R969 B.n309 B.n108 10.6151
R970 B.n313 B.n108 10.6151
R971 B.n314 B.n313 10.6151
R972 B.n315 B.n314 10.6151
R973 B.n315 B.n106 10.6151
R974 B.n319 B.n106 10.6151
R975 B.n320 B.n319 10.6151
R976 B.n321 B.n320 10.6151
R977 B.n321 B.n104 10.6151
R978 B.n325 B.n104 10.6151
R979 B.n326 B.n325 10.6151
R980 B.n327 B.n326 10.6151
R981 B.n327 B.n102 10.6151
R982 B.n331 B.n102 10.6151
R983 B.n332 B.n331 10.6151
R984 B.n333 B.n332 10.6151
R985 B.n333 B.n100 10.6151
R986 B.n337 B.n100 10.6151
R987 B.n338 B.n337 10.6151
R988 B.n339 B.n338 10.6151
R989 B.n339 B.n98 10.6151
R990 B.n343 B.n98 10.6151
R991 B.n344 B.n343 10.6151
R992 B.n345 B.n344 10.6151
R993 B.n345 B.n96 10.6151
R994 B.n349 B.n96 10.6151
R995 B.n350 B.n349 10.6151
R996 B.n351 B.n350 10.6151
R997 B.n351 B.n94 10.6151
R998 B.n355 B.n94 10.6151
R999 B.n356 B.n355 10.6151
R1000 B.n357 B.n356 10.6151
R1001 B.n357 B.n92 10.6151
R1002 B.n361 B.n92 10.6151
R1003 B.n362 B.n361 10.6151
R1004 B.n363 B.n362 10.6151
R1005 B.n363 B.n90 10.6151
R1006 B.n367 B.n90 10.6151
R1007 B.n368 B.n367 10.6151
R1008 B.n369 B.n368 10.6151
R1009 B.n369 B.n88 10.6151
R1010 B.n373 B.n88 10.6151
R1011 B.n374 B.n373 10.6151
R1012 B.n375 B.n374 10.6151
R1013 B.n375 B.n86 10.6151
R1014 B.n379 B.n86 10.6151
R1015 B.n380 B.n379 10.6151
R1016 B.n381 B.n380 10.6151
R1017 B.n381 B.n84 10.6151
R1018 B.n385 B.n84 10.6151
R1019 B.n386 B.n385 10.6151
R1020 B.n387 B.n386 10.6151
R1021 B.n387 B.n82 10.6151
R1022 B.n391 B.n82 10.6151
R1023 B.n392 B.n391 10.6151
R1024 B.n393 B.n392 10.6151
R1025 B.n393 B.n80 10.6151
R1026 B.n397 B.n80 10.6151
R1027 B.n398 B.n397 10.6151
R1028 B.n399 B.n398 10.6151
R1029 B.n399 B.n78 10.6151
R1030 B.n403 B.n78 10.6151
R1031 B.n404 B.n403 10.6151
R1032 B.n405 B.n404 10.6151
R1033 B.n405 B.n76 10.6151
R1034 B.n409 B.n76 10.6151
R1035 B.n410 B.n409 10.6151
R1036 B.n411 B.n410 10.6151
R1037 B.n411 B.n74 10.6151
R1038 B.n415 B.n74 10.6151
R1039 B.n416 B.n415 10.6151
R1040 B.n417 B.n416 10.6151
R1041 B.n417 B.n72 10.6151
R1042 B.n421 B.n72 10.6151
R1043 B.n422 B.n421 10.6151
R1044 B.n423 B.n422 10.6151
R1045 B.n423 B.n70 10.6151
R1046 B.n427 B.n70 10.6151
R1047 B.n428 B.n427 10.6151
R1048 B.n429 B.n428 10.6151
R1049 B.n429 B.n68 10.6151
R1050 B.n433 B.n68 10.6151
R1051 B.n434 B.n433 10.6151
R1052 B.n435 B.n434 10.6151
R1053 B.n435 B.n66 10.6151
R1054 B.n439 B.n66 10.6151
R1055 B.n440 B.n439 10.6151
R1056 B.n441 B.n440 10.6151
R1057 B.n441 B.n64 10.6151
R1058 B.n445 B.n64 10.6151
R1059 B.n446 B.n445 10.6151
R1060 B.n447 B.n446 10.6151
R1061 B.n447 B.n62 10.6151
R1062 B.n451 B.n62 10.6151
R1063 B.n452 B.n451 10.6151
R1064 B.n453 B.n452 10.6151
R1065 B.n453 B.n60 10.6151
R1066 B.n457 B.n60 10.6151
R1067 B.n458 B.n457 10.6151
R1068 B.n459 B.n458 10.6151
R1069 B.n459 B.n58 10.6151
R1070 B.n463 B.n58 10.6151
R1071 B.n464 B.n463 10.6151
R1072 B.n465 B.n464 10.6151
R1073 B.n465 B.n56 10.6151
R1074 B.n469 B.n56 10.6151
R1075 B.n470 B.n469 10.6151
R1076 B.n471 B.n470 10.6151
R1077 B.n471 B.n54 10.6151
R1078 B.n475 B.n54 10.6151
R1079 B.n476 B.n475 10.6151
R1080 B.n477 B.n476 10.6151
R1081 B.n477 B.n52 10.6151
R1082 B.n481 B.n52 10.6151
R1083 B.n482 B.n481 10.6151
R1084 B.n255 B.n254 10.6151
R1085 B.n255 B.n130 10.6151
R1086 B.n259 B.n130 10.6151
R1087 B.n260 B.n259 10.6151
R1088 B.n261 B.n260 10.6151
R1089 B.n261 B.n128 10.6151
R1090 B.n265 B.n128 10.6151
R1091 B.n266 B.n265 10.6151
R1092 B.n268 B.n124 10.6151
R1093 B.n272 B.n124 10.6151
R1094 B.n273 B.n272 10.6151
R1095 B.n274 B.n273 10.6151
R1096 B.n274 B.n122 10.6151
R1097 B.n278 B.n122 10.6151
R1098 B.n279 B.n278 10.6151
R1099 B.n280 B.n279 10.6151
R1100 B.n284 B.n283 10.6151
R1101 B.n285 B.n284 10.6151
R1102 B.n285 B.n116 10.6151
R1103 B.n289 B.n116 10.6151
R1104 B.n290 B.n289 10.6151
R1105 B.n291 B.n290 10.6151
R1106 B.n291 B.n114 10.6151
R1107 B.n295 B.n114 10.6151
R1108 B.n253 B.n132 10.6151
R1109 B.n249 B.n132 10.6151
R1110 B.n249 B.n248 10.6151
R1111 B.n248 B.n247 10.6151
R1112 B.n247 B.n134 10.6151
R1113 B.n243 B.n134 10.6151
R1114 B.n243 B.n242 10.6151
R1115 B.n242 B.n241 10.6151
R1116 B.n241 B.n136 10.6151
R1117 B.n237 B.n136 10.6151
R1118 B.n237 B.n236 10.6151
R1119 B.n236 B.n235 10.6151
R1120 B.n235 B.n138 10.6151
R1121 B.n231 B.n138 10.6151
R1122 B.n231 B.n230 10.6151
R1123 B.n230 B.n229 10.6151
R1124 B.n229 B.n140 10.6151
R1125 B.n225 B.n140 10.6151
R1126 B.n225 B.n224 10.6151
R1127 B.n224 B.n223 10.6151
R1128 B.n223 B.n142 10.6151
R1129 B.n219 B.n142 10.6151
R1130 B.n219 B.n218 10.6151
R1131 B.n218 B.n217 10.6151
R1132 B.n217 B.n144 10.6151
R1133 B.n213 B.n144 10.6151
R1134 B.n213 B.n212 10.6151
R1135 B.n212 B.n211 10.6151
R1136 B.n211 B.n146 10.6151
R1137 B.n207 B.n146 10.6151
R1138 B.n207 B.n206 10.6151
R1139 B.n206 B.n205 10.6151
R1140 B.n205 B.n148 10.6151
R1141 B.n201 B.n148 10.6151
R1142 B.n201 B.n200 10.6151
R1143 B.n200 B.n199 10.6151
R1144 B.n199 B.n150 10.6151
R1145 B.n195 B.n150 10.6151
R1146 B.n195 B.n194 10.6151
R1147 B.n194 B.n193 10.6151
R1148 B.n193 B.n152 10.6151
R1149 B.n189 B.n152 10.6151
R1150 B.n189 B.n188 10.6151
R1151 B.n188 B.n187 10.6151
R1152 B.n187 B.n154 10.6151
R1153 B.n183 B.n154 10.6151
R1154 B.n183 B.n182 10.6151
R1155 B.n182 B.n181 10.6151
R1156 B.n181 B.n156 10.6151
R1157 B.n177 B.n156 10.6151
R1158 B.n177 B.n176 10.6151
R1159 B.n176 B.n175 10.6151
R1160 B.n175 B.n158 10.6151
R1161 B.n171 B.n158 10.6151
R1162 B.n171 B.n170 10.6151
R1163 B.n170 B.n169 10.6151
R1164 B.n169 B.n160 10.6151
R1165 B.n165 B.n160 10.6151
R1166 B.n165 B.n164 10.6151
R1167 B.n164 B.n163 10.6151
R1168 B.n163 B.n0 10.6151
R1169 B.n615 B.n1 10.6151
R1170 B.n615 B.n614 10.6151
R1171 B.n614 B.n613 10.6151
R1172 B.n613 B.n4 10.6151
R1173 B.n609 B.n4 10.6151
R1174 B.n609 B.n608 10.6151
R1175 B.n608 B.n607 10.6151
R1176 B.n607 B.n6 10.6151
R1177 B.n603 B.n6 10.6151
R1178 B.n603 B.n602 10.6151
R1179 B.n602 B.n601 10.6151
R1180 B.n601 B.n8 10.6151
R1181 B.n597 B.n8 10.6151
R1182 B.n597 B.n596 10.6151
R1183 B.n596 B.n595 10.6151
R1184 B.n595 B.n10 10.6151
R1185 B.n591 B.n10 10.6151
R1186 B.n591 B.n590 10.6151
R1187 B.n590 B.n589 10.6151
R1188 B.n589 B.n12 10.6151
R1189 B.n585 B.n12 10.6151
R1190 B.n585 B.n584 10.6151
R1191 B.n584 B.n583 10.6151
R1192 B.n583 B.n14 10.6151
R1193 B.n579 B.n14 10.6151
R1194 B.n579 B.n578 10.6151
R1195 B.n578 B.n577 10.6151
R1196 B.n577 B.n16 10.6151
R1197 B.n573 B.n16 10.6151
R1198 B.n573 B.n572 10.6151
R1199 B.n572 B.n571 10.6151
R1200 B.n571 B.n18 10.6151
R1201 B.n567 B.n18 10.6151
R1202 B.n567 B.n566 10.6151
R1203 B.n566 B.n565 10.6151
R1204 B.n565 B.n20 10.6151
R1205 B.n561 B.n20 10.6151
R1206 B.n561 B.n560 10.6151
R1207 B.n560 B.n559 10.6151
R1208 B.n559 B.n22 10.6151
R1209 B.n555 B.n22 10.6151
R1210 B.n555 B.n554 10.6151
R1211 B.n554 B.n553 10.6151
R1212 B.n553 B.n24 10.6151
R1213 B.n549 B.n24 10.6151
R1214 B.n549 B.n548 10.6151
R1215 B.n548 B.n547 10.6151
R1216 B.n547 B.n26 10.6151
R1217 B.n543 B.n26 10.6151
R1218 B.n543 B.n542 10.6151
R1219 B.n542 B.n541 10.6151
R1220 B.n541 B.n28 10.6151
R1221 B.n537 B.n28 10.6151
R1222 B.n537 B.n536 10.6151
R1223 B.n536 B.n535 10.6151
R1224 B.n535 B.n30 10.6151
R1225 B.n531 B.n30 10.6151
R1226 B.n531 B.n530 10.6151
R1227 B.n530 B.n529 10.6151
R1228 B.n529 B.n32 10.6151
R1229 B.n525 B.n32 10.6151
R1230 B.n511 B.n510 6.5566
R1231 B.n498 B.n46 6.5566
R1232 B.n268 B.n267 6.5566
R1233 B.n280 B.n120 6.5566
R1234 B.n512 B.n511 4.05904
R1235 B.n495 B.n46 4.05904
R1236 B.n267 B.n266 4.05904
R1237 B.n283 B.n120 4.05904
R1238 B.n619 B.n0 2.81026
R1239 B.n619 B.n1 2.81026
C0 VTAIL VP 2.74681f
C1 VTAIL VDD1 5.03296f
C2 B VDD2 1.69625f
C3 w_n4650_n1120# VDD2 2.02671f
C4 VN VDD2 1.03373f
C5 VP VDD2 0.609601f
C6 w_n4650_n1120# B 8.2524f
C7 VN B 1.21827f
C8 w_n4650_n1120# VN 9.51439f
C9 VDD1 VDD2 2.16401f
C10 B VP 2.23652f
C11 w_n4650_n1120# VP 10.1116f
C12 VN VP 6.50228f
C13 B VDD1 1.57574f
C14 VTAIL VDD2 5.0924f
C15 w_n4650_n1120# VDD1 1.88176f
C16 VN VDD1 0.160728f
C17 VDD1 VP 1.47765f
C18 VTAIL B 1.24732f
C19 VTAIL w_n4650_n1120# 1.72149f
C20 VTAIL VN 2.7327f
C21 VDD2 VSUBS 1.757041f
C22 VDD1 VSUBS 2.268828f
C23 VTAIL VSUBS 0.705189f
C24 VN VSUBS 8.44728f
C25 VP VSUBS 3.696873f
C26 B VSUBS 4.58358f
C27 w_n4650_n1120# VSUBS 67.3506f
C28 B.n0 VSUBS 0.008352f
C29 B.n1 VSUBS 0.008352f
C30 B.n2 VSUBS 0.013209f
C31 B.n3 VSUBS 0.013209f
C32 B.n4 VSUBS 0.013209f
C33 B.n5 VSUBS 0.013209f
C34 B.n6 VSUBS 0.013209f
C35 B.n7 VSUBS 0.013209f
C36 B.n8 VSUBS 0.013209f
C37 B.n9 VSUBS 0.013209f
C38 B.n10 VSUBS 0.013209f
C39 B.n11 VSUBS 0.013209f
C40 B.n12 VSUBS 0.013209f
C41 B.n13 VSUBS 0.013209f
C42 B.n14 VSUBS 0.013209f
C43 B.n15 VSUBS 0.013209f
C44 B.n16 VSUBS 0.013209f
C45 B.n17 VSUBS 0.013209f
C46 B.n18 VSUBS 0.013209f
C47 B.n19 VSUBS 0.013209f
C48 B.n20 VSUBS 0.013209f
C49 B.n21 VSUBS 0.013209f
C50 B.n22 VSUBS 0.013209f
C51 B.n23 VSUBS 0.013209f
C52 B.n24 VSUBS 0.013209f
C53 B.n25 VSUBS 0.013209f
C54 B.n26 VSUBS 0.013209f
C55 B.n27 VSUBS 0.013209f
C56 B.n28 VSUBS 0.013209f
C57 B.n29 VSUBS 0.013209f
C58 B.n30 VSUBS 0.013209f
C59 B.n31 VSUBS 0.013209f
C60 B.n32 VSUBS 0.013209f
C61 B.n33 VSUBS 0.032488f
C62 B.n34 VSUBS 0.013209f
C63 B.n35 VSUBS 0.013209f
C64 B.n36 VSUBS 0.013209f
C65 B.n37 VSUBS 0.013209f
C66 B.t2 VSUBS 0.027447f
C67 B.t1 VSUBS 0.033971f
C68 B.t0 VSUBS 0.242262f
C69 B.n38 VSUBS 0.126453f
C70 B.n39 VSUBS 0.084985f
C71 B.n40 VSUBS 0.013209f
C72 B.n41 VSUBS 0.013209f
C73 B.n42 VSUBS 0.013209f
C74 B.n43 VSUBS 0.013209f
C75 B.t8 VSUBS 0.027447f
C76 B.t7 VSUBS 0.033971f
C77 B.t6 VSUBS 0.242262f
C78 B.n44 VSUBS 0.126453f
C79 B.n45 VSUBS 0.084985f
C80 B.n46 VSUBS 0.030603f
C81 B.n47 VSUBS 0.013209f
C82 B.n48 VSUBS 0.013209f
C83 B.n49 VSUBS 0.013209f
C84 B.n50 VSUBS 0.013209f
C85 B.n51 VSUBS 0.030058f
C86 B.n52 VSUBS 0.013209f
C87 B.n53 VSUBS 0.013209f
C88 B.n54 VSUBS 0.013209f
C89 B.n55 VSUBS 0.013209f
C90 B.n56 VSUBS 0.013209f
C91 B.n57 VSUBS 0.013209f
C92 B.n58 VSUBS 0.013209f
C93 B.n59 VSUBS 0.013209f
C94 B.n60 VSUBS 0.013209f
C95 B.n61 VSUBS 0.013209f
C96 B.n62 VSUBS 0.013209f
C97 B.n63 VSUBS 0.013209f
C98 B.n64 VSUBS 0.013209f
C99 B.n65 VSUBS 0.013209f
C100 B.n66 VSUBS 0.013209f
C101 B.n67 VSUBS 0.013209f
C102 B.n68 VSUBS 0.013209f
C103 B.n69 VSUBS 0.013209f
C104 B.n70 VSUBS 0.013209f
C105 B.n71 VSUBS 0.013209f
C106 B.n72 VSUBS 0.013209f
C107 B.n73 VSUBS 0.013209f
C108 B.n74 VSUBS 0.013209f
C109 B.n75 VSUBS 0.013209f
C110 B.n76 VSUBS 0.013209f
C111 B.n77 VSUBS 0.013209f
C112 B.n78 VSUBS 0.013209f
C113 B.n79 VSUBS 0.013209f
C114 B.n80 VSUBS 0.013209f
C115 B.n81 VSUBS 0.013209f
C116 B.n82 VSUBS 0.013209f
C117 B.n83 VSUBS 0.013209f
C118 B.n84 VSUBS 0.013209f
C119 B.n85 VSUBS 0.013209f
C120 B.n86 VSUBS 0.013209f
C121 B.n87 VSUBS 0.013209f
C122 B.n88 VSUBS 0.013209f
C123 B.n89 VSUBS 0.013209f
C124 B.n90 VSUBS 0.013209f
C125 B.n91 VSUBS 0.013209f
C126 B.n92 VSUBS 0.013209f
C127 B.n93 VSUBS 0.013209f
C128 B.n94 VSUBS 0.013209f
C129 B.n95 VSUBS 0.013209f
C130 B.n96 VSUBS 0.013209f
C131 B.n97 VSUBS 0.013209f
C132 B.n98 VSUBS 0.013209f
C133 B.n99 VSUBS 0.013209f
C134 B.n100 VSUBS 0.013209f
C135 B.n101 VSUBS 0.013209f
C136 B.n102 VSUBS 0.013209f
C137 B.n103 VSUBS 0.013209f
C138 B.n104 VSUBS 0.013209f
C139 B.n105 VSUBS 0.013209f
C140 B.n106 VSUBS 0.013209f
C141 B.n107 VSUBS 0.013209f
C142 B.n108 VSUBS 0.013209f
C143 B.n109 VSUBS 0.013209f
C144 B.n110 VSUBS 0.013209f
C145 B.n111 VSUBS 0.013209f
C146 B.n112 VSUBS 0.013209f
C147 B.n113 VSUBS 0.030058f
C148 B.n114 VSUBS 0.013209f
C149 B.n115 VSUBS 0.013209f
C150 B.n116 VSUBS 0.013209f
C151 B.n117 VSUBS 0.013209f
C152 B.t10 VSUBS 0.027447f
C153 B.t11 VSUBS 0.033971f
C154 B.t9 VSUBS 0.242262f
C155 B.n118 VSUBS 0.126453f
C156 B.n119 VSUBS 0.084985f
C157 B.n120 VSUBS 0.030603f
C158 B.n121 VSUBS 0.013209f
C159 B.n122 VSUBS 0.013209f
C160 B.n123 VSUBS 0.013209f
C161 B.n124 VSUBS 0.013209f
C162 B.n125 VSUBS 0.013209f
C163 B.t4 VSUBS 0.027447f
C164 B.t5 VSUBS 0.033971f
C165 B.t3 VSUBS 0.242262f
C166 B.n126 VSUBS 0.126453f
C167 B.n127 VSUBS 0.084985f
C168 B.n128 VSUBS 0.013209f
C169 B.n129 VSUBS 0.013209f
C170 B.n130 VSUBS 0.013209f
C171 B.n131 VSUBS 0.032488f
C172 B.n132 VSUBS 0.013209f
C173 B.n133 VSUBS 0.013209f
C174 B.n134 VSUBS 0.013209f
C175 B.n135 VSUBS 0.013209f
C176 B.n136 VSUBS 0.013209f
C177 B.n137 VSUBS 0.013209f
C178 B.n138 VSUBS 0.013209f
C179 B.n139 VSUBS 0.013209f
C180 B.n140 VSUBS 0.013209f
C181 B.n141 VSUBS 0.013209f
C182 B.n142 VSUBS 0.013209f
C183 B.n143 VSUBS 0.013209f
C184 B.n144 VSUBS 0.013209f
C185 B.n145 VSUBS 0.013209f
C186 B.n146 VSUBS 0.013209f
C187 B.n147 VSUBS 0.013209f
C188 B.n148 VSUBS 0.013209f
C189 B.n149 VSUBS 0.013209f
C190 B.n150 VSUBS 0.013209f
C191 B.n151 VSUBS 0.013209f
C192 B.n152 VSUBS 0.013209f
C193 B.n153 VSUBS 0.013209f
C194 B.n154 VSUBS 0.013209f
C195 B.n155 VSUBS 0.013209f
C196 B.n156 VSUBS 0.013209f
C197 B.n157 VSUBS 0.013209f
C198 B.n158 VSUBS 0.013209f
C199 B.n159 VSUBS 0.013209f
C200 B.n160 VSUBS 0.013209f
C201 B.n161 VSUBS 0.013209f
C202 B.n162 VSUBS 0.013209f
C203 B.n163 VSUBS 0.013209f
C204 B.n164 VSUBS 0.013209f
C205 B.n165 VSUBS 0.013209f
C206 B.n166 VSUBS 0.013209f
C207 B.n167 VSUBS 0.013209f
C208 B.n168 VSUBS 0.013209f
C209 B.n169 VSUBS 0.013209f
C210 B.n170 VSUBS 0.013209f
C211 B.n171 VSUBS 0.013209f
C212 B.n172 VSUBS 0.013209f
C213 B.n173 VSUBS 0.013209f
C214 B.n174 VSUBS 0.013209f
C215 B.n175 VSUBS 0.013209f
C216 B.n176 VSUBS 0.013209f
C217 B.n177 VSUBS 0.013209f
C218 B.n178 VSUBS 0.013209f
C219 B.n179 VSUBS 0.013209f
C220 B.n180 VSUBS 0.013209f
C221 B.n181 VSUBS 0.013209f
C222 B.n182 VSUBS 0.013209f
C223 B.n183 VSUBS 0.013209f
C224 B.n184 VSUBS 0.013209f
C225 B.n185 VSUBS 0.013209f
C226 B.n186 VSUBS 0.013209f
C227 B.n187 VSUBS 0.013209f
C228 B.n188 VSUBS 0.013209f
C229 B.n189 VSUBS 0.013209f
C230 B.n190 VSUBS 0.013209f
C231 B.n191 VSUBS 0.013209f
C232 B.n192 VSUBS 0.013209f
C233 B.n193 VSUBS 0.013209f
C234 B.n194 VSUBS 0.013209f
C235 B.n195 VSUBS 0.013209f
C236 B.n196 VSUBS 0.013209f
C237 B.n197 VSUBS 0.013209f
C238 B.n198 VSUBS 0.013209f
C239 B.n199 VSUBS 0.013209f
C240 B.n200 VSUBS 0.013209f
C241 B.n201 VSUBS 0.013209f
C242 B.n202 VSUBS 0.013209f
C243 B.n203 VSUBS 0.013209f
C244 B.n204 VSUBS 0.013209f
C245 B.n205 VSUBS 0.013209f
C246 B.n206 VSUBS 0.013209f
C247 B.n207 VSUBS 0.013209f
C248 B.n208 VSUBS 0.013209f
C249 B.n209 VSUBS 0.013209f
C250 B.n210 VSUBS 0.013209f
C251 B.n211 VSUBS 0.013209f
C252 B.n212 VSUBS 0.013209f
C253 B.n213 VSUBS 0.013209f
C254 B.n214 VSUBS 0.013209f
C255 B.n215 VSUBS 0.013209f
C256 B.n216 VSUBS 0.013209f
C257 B.n217 VSUBS 0.013209f
C258 B.n218 VSUBS 0.013209f
C259 B.n219 VSUBS 0.013209f
C260 B.n220 VSUBS 0.013209f
C261 B.n221 VSUBS 0.013209f
C262 B.n222 VSUBS 0.013209f
C263 B.n223 VSUBS 0.013209f
C264 B.n224 VSUBS 0.013209f
C265 B.n225 VSUBS 0.013209f
C266 B.n226 VSUBS 0.013209f
C267 B.n227 VSUBS 0.013209f
C268 B.n228 VSUBS 0.013209f
C269 B.n229 VSUBS 0.013209f
C270 B.n230 VSUBS 0.013209f
C271 B.n231 VSUBS 0.013209f
C272 B.n232 VSUBS 0.013209f
C273 B.n233 VSUBS 0.013209f
C274 B.n234 VSUBS 0.013209f
C275 B.n235 VSUBS 0.013209f
C276 B.n236 VSUBS 0.013209f
C277 B.n237 VSUBS 0.013209f
C278 B.n238 VSUBS 0.013209f
C279 B.n239 VSUBS 0.013209f
C280 B.n240 VSUBS 0.013209f
C281 B.n241 VSUBS 0.013209f
C282 B.n242 VSUBS 0.013209f
C283 B.n243 VSUBS 0.013209f
C284 B.n244 VSUBS 0.013209f
C285 B.n245 VSUBS 0.013209f
C286 B.n246 VSUBS 0.013209f
C287 B.n247 VSUBS 0.013209f
C288 B.n248 VSUBS 0.013209f
C289 B.n249 VSUBS 0.013209f
C290 B.n250 VSUBS 0.013209f
C291 B.n251 VSUBS 0.013209f
C292 B.n252 VSUBS 0.030058f
C293 B.n253 VSUBS 0.030058f
C294 B.n254 VSUBS 0.032488f
C295 B.n255 VSUBS 0.013209f
C296 B.n256 VSUBS 0.013209f
C297 B.n257 VSUBS 0.013209f
C298 B.n258 VSUBS 0.013209f
C299 B.n259 VSUBS 0.013209f
C300 B.n260 VSUBS 0.013209f
C301 B.n261 VSUBS 0.013209f
C302 B.n262 VSUBS 0.013209f
C303 B.n263 VSUBS 0.013209f
C304 B.n264 VSUBS 0.013209f
C305 B.n265 VSUBS 0.013209f
C306 B.n266 VSUBS 0.009129f
C307 B.n267 VSUBS 0.030603f
C308 B.n268 VSUBS 0.010683f
C309 B.n269 VSUBS 0.013209f
C310 B.n270 VSUBS 0.013209f
C311 B.n271 VSUBS 0.013209f
C312 B.n272 VSUBS 0.013209f
C313 B.n273 VSUBS 0.013209f
C314 B.n274 VSUBS 0.013209f
C315 B.n275 VSUBS 0.013209f
C316 B.n276 VSUBS 0.013209f
C317 B.n277 VSUBS 0.013209f
C318 B.n278 VSUBS 0.013209f
C319 B.n279 VSUBS 0.013209f
C320 B.n280 VSUBS 0.010683f
C321 B.n281 VSUBS 0.013209f
C322 B.n282 VSUBS 0.013209f
C323 B.n283 VSUBS 0.009129f
C324 B.n284 VSUBS 0.013209f
C325 B.n285 VSUBS 0.013209f
C326 B.n286 VSUBS 0.013209f
C327 B.n287 VSUBS 0.013209f
C328 B.n288 VSUBS 0.013209f
C329 B.n289 VSUBS 0.013209f
C330 B.n290 VSUBS 0.013209f
C331 B.n291 VSUBS 0.013209f
C332 B.n292 VSUBS 0.013209f
C333 B.n293 VSUBS 0.013209f
C334 B.n294 VSUBS 0.032488f
C335 B.n295 VSUBS 0.032488f
C336 B.n296 VSUBS 0.030058f
C337 B.n297 VSUBS 0.013209f
C338 B.n298 VSUBS 0.013209f
C339 B.n299 VSUBS 0.013209f
C340 B.n300 VSUBS 0.013209f
C341 B.n301 VSUBS 0.013209f
C342 B.n302 VSUBS 0.013209f
C343 B.n303 VSUBS 0.013209f
C344 B.n304 VSUBS 0.013209f
C345 B.n305 VSUBS 0.013209f
C346 B.n306 VSUBS 0.013209f
C347 B.n307 VSUBS 0.013209f
C348 B.n308 VSUBS 0.013209f
C349 B.n309 VSUBS 0.013209f
C350 B.n310 VSUBS 0.013209f
C351 B.n311 VSUBS 0.013209f
C352 B.n312 VSUBS 0.013209f
C353 B.n313 VSUBS 0.013209f
C354 B.n314 VSUBS 0.013209f
C355 B.n315 VSUBS 0.013209f
C356 B.n316 VSUBS 0.013209f
C357 B.n317 VSUBS 0.013209f
C358 B.n318 VSUBS 0.013209f
C359 B.n319 VSUBS 0.013209f
C360 B.n320 VSUBS 0.013209f
C361 B.n321 VSUBS 0.013209f
C362 B.n322 VSUBS 0.013209f
C363 B.n323 VSUBS 0.013209f
C364 B.n324 VSUBS 0.013209f
C365 B.n325 VSUBS 0.013209f
C366 B.n326 VSUBS 0.013209f
C367 B.n327 VSUBS 0.013209f
C368 B.n328 VSUBS 0.013209f
C369 B.n329 VSUBS 0.013209f
C370 B.n330 VSUBS 0.013209f
C371 B.n331 VSUBS 0.013209f
C372 B.n332 VSUBS 0.013209f
C373 B.n333 VSUBS 0.013209f
C374 B.n334 VSUBS 0.013209f
C375 B.n335 VSUBS 0.013209f
C376 B.n336 VSUBS 0.013209f
C377 B.n337 VSUBS 0.013209f
C378 B.n338 VSUBS 0.013209f
C379 B.n339 VSUBS 0.013209f
C380 B.n340 VSUBS 0.013209f
C381 B.n341 VSUBS 0.013209f
C382 B.n342 VSUBS 0.013209f
C383 B.n343 VSUBS 0.013209f
C384 B.n344 VSUBS 0.013209f
C385 B.n345 VSUBS 0.013209f
C386 B.n346 VSUBS 0.013209f
C387 B.n347 VSUBS 0.013209f
C388 B.n348 VSUBS 0.013209f
C389 B.n349 VSUBS 0.013209f
C390 B.n350 VSUBS 0.013209f
C391 B.n351 VSUBS 0.013209f
C392 B.n352 VSUBS 0.013209f
C393 B.n353 VSUBS 0.013209f
C394 B.n354 VSUBS 0.013209f
C395 B.n355 VSUBS 0.013209f
C396 B.n356 VSUBS 0.013209f
C397 B.n357 VSUBS 0.013209f
C398 B.n358 VSUBS 0.013209f
C399 B.n359 VSUBS 0.013209f
C400 B.n360 VSUBS 0.013209f
C401 B.n361 VSUBS 0.013209f
C402 B.n362 VSUBS 0.013209f
C403 B.n363 VSUBS 0.013209f
C404 B.n364 VSUBS 0.013209f
C405 B.n365 VSUBS 0.013209f
C406 B.n366 VSUBS 0.013209f
C407 B.n367 VSUBS 0.013209f
C408 B.n368 VSUBS 0.013209f
C409 B.n369 VSUBS 0.013209f
C410 B.n370 VSUBS 0.013209f
C411 B.n371 VSUBS 0.013209f
C412 B.n372 VSUBS 0.013209f
C413 B.n373 VSUBS 0.013209f
C414 B.n374 VSUBS 0.013209f
C415 B.n375 VSUBS 0.013209f
C416 B.n376 VSUBS 0.013209f
C417 B.n377 VSUBS 0.013209f
C418 B.n378 VSUBS 0.013209f
C419 B.n379 VSUBS 0.013209f
C420 B.n380 VSUBS 0.013209f
C421 B.n381 VSUBS 0.013209f
C422 B.n382 VSUBS 0.013209f
C423 B.n383 VSUBS 0.013209f
C424 B.n384 VSUBS 0.013209f
C425 B.n385 VSUBS 0.013209f
C426 B.n386 VSUBS 0.013209f
C427 B.n387 VSUBS 0.013209f
C428 B.n388 VSUBS 0.013209f
C429 B.n389 VSUBS 0.013209f
C430 B.n390 VSUBS 0.013209f
C431 B.n391 VSUBS 0.013209f
C432 B.n392 VSUBS 0.013209f
C433 B.n393 VSUBS 0.013209f
C434 B.n394 VSUBS 0.013209f
C435 B.n395 VSUBS 0.013209f
C436 B.n396 VSUBS 0.013209f
C437 B.n397 VSUBS 0.013209f
C438 B.n398 VSUBS 0.013209f
C439 B.n399 VSUBS 0.013209f
C440 B.n400 VSUBS 0.013209f
C441 B.n401 VSUBS 0.013209f
C442 B.n402 VSUBS 0.013209f
C443 B.n403 VSUBS 0.013209f
C444 B.n404 VSUBS 0.013209f
C445 B.n405 VSUBS 0.013209f
C446 B.n406 VSUBS 0.013209f
C447 B.n407 VSUBS 0.013209f
C448 B.n408 VSUBS 0.013209f
C449 B.n409 VSUBS 0.013209f
C450 B.n410 VSUBS 0.013209f
C451 B.n411 VSUBS 0.013209f
C452 B.n412 VSUBS 0.013209f
C453 B.n413 VSUBS 0.013209f
C454 B.n414 VSUBS 0.013209f
C455 B.n415 VSUBS 0.013209f
C456 B.n416 VSUBS 0.013209f
C457 B.n417 VSUBS 0.013209f
C458 B.n418 VSUBS 0.013209f
C459 B.n419 VSUBS 0.013209f
C460 B.n420 VSUBS 0.013209f
C461 B.n421 VSUBS 0.013209f
C462 B.n422 VSUBS 0.013209f
C463 B.n423 VSUBS 0.013209f
C464 B.n424 VSUBS 0.013209f
C465 B.n425 VSUBS 0.013209f
C466 B.n426 VSUBS 0.013209f
C467 B.n427 VSUBS 0.013209f
C468 B.n428 VSUBS 0.013209f
C469 B.n429 VSUBS 0.013209f
C470 B.n430 VSUBS 0.013209f
C471 B.n431 VSUBS 0.013209f
C472 B.n432 VSUBS 0.013209f
C473 B.n433 VSUBS 0.013209f
C474 B.n434 VSUBS 0.013209f
C475 B.n435 VSUBS 0.013209f
C476 B.n436 VSUBS 0.013209f
C477 B.n437 VSUBS 0.013209f
C478 B.n438 VSUBS 0.013209f
C479 B.n439 VSUBS 0.013209f
C480 B.n440 VSUBS 0.013209f
C481 B.n441 VSUBS 0.013209f
C482 B.n442 VSUBS 0.013209f
C483 B.n443 VSUBS 0.013209f
C484 B.n444 VSUBS 0.013209f
C485 B.n445 VSUBS 0.013209f
C486 B.n446 VSUBS 0.013209f
C487 B.n447 VSUBS 0.013209f
C488 B.n448 VSUBS 0.013209f
C489 B.n449 VSUBS 0.013209f
C490 B.n450 VSUBS 0.013209f
C491 B.n451 VSUBS 0.013209f
C492 B.n452 VSUBS 0.013209f
C493 B.n453 VSUBS 0.013209f
C494 B.n454 VSUBS 0.013209f
C495 B.n455 VSUBS 0.013209f
C496 B.n456 VSUBS 0.013209f
C497 B.n457 VSUBS 0.013209f
C498 B.n458 VSUBS 0.013209f
C499 B.n459 VSUBS 0.013209f
C500 B.n460 VSUBS 0.013209f
C501 B.n461 VSUBS 0.013209f
C502 B.n462 VSUBS 0.013209f
C503 B.n463 VSUBS 0.013209f
C504 B.n464 VSUBS 0.013209f
C505 B.n465 VSUBS 0.013209f
C506 B.n466 VSUBS 0.013209f
C507 B.n467 VSUBS 0.013209f
C508 B.n468 VSUBS 0.013209f
C509 B.n469 VSUBS 0.013209f
C510 B.n470 VSUBS 0.013209f
C511 B.n471 VSUBS 0.013209f
C512 B.n472 VSUBS 0.013209f
C513 B.n473 VSUBS 0.013209f
C514 B.n474 VSUBS 0.013209f
C515 B.n475 VSUBS 0.013209f
C516 B.n476 VSUBS 0.013209f
C517 B.n477 VSUBS 0.013209f
C518 B.n478 VSUBS 0.013209f
C519 B.n479 VSUBS 0.013209f
C520 B.n480 VSUBS 0.013209f
C521 B.n481 VSUBS 0.013209f
C522 B.n482 VSUBS 0.031591f
C523 B.n483 VSUBS 0.030955f
C524 B.n484 VSUBS 0.032488f
C525 B.n485 VSUBS 0.013209f
C526 B.n486 VSUBS 0.013209f
C527 B.n487 VSUBS 0.013209f
C528 B.n488 VSUBS 0.013209f
C529 B.n489 VSUBS 0.013209f
C530 B.n490 VSUBS 0.013209f
C531 B.n491 VSUBS 0.013209f
C532 B.n492 VSUBS 0.013209f
C533 B.n493 VSUBS 0.013209f
C534 B.n494 VSUBS 0.013209f
C535 B.n495 VSUBS 0.009129f
C536 B.n496 VSUBS 0.013209f
C537 B.n497 VSUBS 0.013209f
C538 B.n498 VSUBS 0.010683f
C539 B.n499 VSUBS 0.013209f
C540 B.n500 VSUBS 0.013209f
C541 B.n501 VSUBS 0.013209f
C542 B.n502 VSUBS 0.013209f
C543 B.n503 VSUBS 0.013209f
C544 B.n504 VSUBS 0.013209f
C545 B.n505 VSUBS 0.013209f
C546 B.n506 VSUBS 0.013209f
C547 B.n507 VSUBS 0.013209f
C548 B.n508 VSUBS 0.013209f
C549 B.n509 VSUBS 0.013209f
C550 B.n510 VSUBS 0.010683f
C551 B.n511 VSUBS 0.030603f
C552 B.n512 VSUBS 0.009129f
C553 B.n513 VSUBS 0.013209f
C554 B.n514 VSUBS 0.013209f
C555 B.n515 VSUBS 0.013209f
C556 B.n516 VSUBS 0.013209f
C557 B.n517 VSUBS 0.013209f
C558 B.n518 VSUBS 0.013209f
C559 B.n519 VSUBS 0.013209f
C560 B.n520 VSUBS 0.013209f
C561 B.n521 VSUBS 0.013209f
C562 B.n522 VSUBS 0.013209f
C563 B.n523 VSUBS 0.013209f
C564 B.n524 VSUBS 0.032488f
C565 B.n525 VSUBS 0.030058f
C566 B.n526 VSUBS 0.030058f
C567 B.n527 VSUBS 0.013209f
C568 B.n528 VSUBS 0.013209f
C569 B.n529 VSUBS 0.013209f
C570 B.n530 VSUBS 0.013209f
C571 B.n531 VSUBS 0.013209f
C572 B.n532 VSUBS 0.013209f
C573 B.n533 VSUBS 0.013209f
C574 B.n534 VSUBS 0.013209f
C575 B.n535 VSUBS 0.013209f
C576 B.n536 VSUBS 0.013209f
C577 B.n537 VSUBS 0.013209f
C578 B.n538 VSUBS 0.013209f
C579 B.n539 VSUBS 0.013209f
C580 B.n540 VSUBS 0.013209f
C581 B.n541 VSUBS 0.013209f
C582 B.n542 VSUBS 0.013209f
C583 B.n543 VSUBS 0.013209f
C584 B.n544 VSUBS 0.013209f
C585 B.n545 VSUBS 0.013209f
C586 B.n546 VSUBS 0.013209f
C587 B.n547 VSUBS 0.013209f
C588 B.n548 VSUBS 0.013209f
C589 B.n549 VSUBS 0.013209f
C590 B.n550 VSUBS 0.013209f
C591 B.n551 VSUBS 0.013209f
C592 B.n552 VSUBS 0.013209f
C593 B.n553 VSUBS 0.013209f
C594 B.n554 VSUBS 0.013209f
C595 B.n555 VSUBS 0.013209f
C596 B.n556 VSUBS 0.013209f
C597 B.n557 VSUBS 0.013209f
C598 B.n558 VSUBS 0.013209f
C599 B.n559 VSUBS 0.013209f
C600 B.n560 VSUBS 0.013209f
C601 B.n561 VSUBS 0.013209f
C602 B.n562 VSUBS 0.013209f
C603 B.n563 VSUBS 0.013209f
C604 B.n564 VSUBS 0.013209f
C605 B.n565 VSUBS 0.013209f
C606 B.n566 VSUBS 0.013209f
C607 B.n567 VSUBS 0.013209f
C608 B.n568 VSUBS 0.013209f
C609 B.n569 VSUBS 0.013209f
C610 B.n570 VSUBS 0.013209f
C611 B.n571 VSUBS 0.013209f
C612 B.n572 VSUBS 0.013209f
C613 B.n573 VSUBS 0.013209f
C614 B.n574 VSUBS 0.013209f
C615 B.n575 VSUBS 0.013209f
C616 B.n576 VSUBS 0.013209f
C617 B.n577 VSUBS 0.013209f
C618 B.n578 VSUBS 0.013209f
C619 B.n579 VSUBS 0.013209f
C620 B.n580 VSUBS 0.013209f
C621 B.n581 VSUBS 0.013209f
C622 B.n582 VSUBS 0.013209f
C623 B.n583 VSUBS 0.013209f
C624 B.n584 VSUBS 0.013209f
C625 B.n585 VSUBS 0.013209f
C626 B.n586 VSUBS 0.013209f
C627 B.n587 VSUBS 0.013209f
C628 B.n588 VSUBS 0.013209f
C629 B.n589 VSUBS 0.013209f
C630 B.n590 VSUBS 0.013209f
C631 B.n591 VSUBS 0.013209f
C632 B.n592 VSUBS 0.013209f
C633 B.n593 VSUBS 0.013209f
C634 B.n594 VSUBS 0.013209f
C635 B.n595 VSUBS 0.013209f
C636 B.n596 VSUBS 0.013209f
C637 B.n597 VSUBS 0.013209f
C638 B.n598 VSUBS 0.013209f
C639 B.n599 VSUBS 0.013209f
C640 B.n600 VSUBS 0.013209f
C641 B.n601 VSUBS 0.013209f
C642 B.n602 VSUBS 0.013209f
C643 B.n603 VSUBS 0.013209f
C644 B.n604 VSUBS 0.013209f
C645 B.n605 VSUBS 0.013209f
C646 B.n606 VSUBS 0.013209f
C647 B.n607 VSUBS 0.013209f
C648 B.n608 VSUBS 0.013209f
C649 B.n609 VSUBS 0.013209f
C650 B.n610 VSUBS 0.013209f
C651 B.n611 VSUBS 0.013209f
C652 B.n612 VSUBS 0.013209f
C653 B.n613 VSUBS 0.013209f
C654 B.n614 VSUBS 0.013209f
C655 B.n615 VSUBS 0.013209f
C656 B.n616 VSUBS 0.013209f
C657 B.n617 VSUBS 0.013209f
C658 B.n618 VSUBS 0.013209f
C659 B.n619 VSUBS 0.029909f
C660 VDD2.t0 VSUBS 0.023506f
C661 VDD2.t1 VSUBS 0.023506f
C662 VDD2.n0 VSUBS 0.052524f
C663 VDD2.t4 VSUBS 0.023506f
C664 VDD2.t5 VSUBS 0.023506f
C665 VDD2.n1 VSUBS 0.052524f
C666 VDD2.n2 VSUBS 4.3434f
C667 VDD2.t7 VSUBS 0.023506f
C668 VDD2.t6 VSUBS 0.023506f
C669 VDD2.n3 VSUBS 0.050806f
C670 VDD2.n4 VSUBS 3.44603f
C671 VDD2.t2 VSUBS 0.023506f
C672 VDD2.t3 VSUBS 0.023506f
C673 VDD2.n5 VSUBS 0.052519f
C674 VN.t2 VSUBS 0.246518f
C675 VN.n0 VSUBS 0.440931f
C676 VN.n1 VSUBS 0.061542f
C677 VN.n2 VSUBS 0.05366f
C678 VN.n3 VSUBS 0.061542f
C679 VN.t3 VSUBS 0.246518f
C680 VN.n4 VSUBS 0.202711f
C681 VN.n5 VSUBS 0.061542f
C682 VN.n6 VSUBS 0.089462f
C683 VN.n7 VSUBS 0.061542f
C684 VN.n8 VSUBS 0.067926f
C685 VN.t6 VSUBS 0.246518f
C686 VN.n9 VSUBS 0.392708f
C687 VN.t7 VSUBS 0.795051f
C688 VN.n10 VSUBS 0.496899f
C689 VN.n11 VSUBS 0.728431f
C690 VN.n12 VSUBS 0.061542f
C691 VN.n13 VSUBS 0.114125f
C692 VN.n14 VSUBS 0.114125f
C693 VN.n15 VSUBS 0.089462f
C694 VN.n16 VSUBS 0.061542f
C695 VN.n17 VSUBS 0.061542f
C696 VN.n18 VSUBS 0.061542f
C697 VN.n19 VSUBS 0.114125f
C698 VN.n20 VSUBS 0.114125f
C699 VN.n21 VSUBS 0.067926f
C700 VN.n22 VSUBS 0.061542f
C701 VN.n23 VSUBS 0.061542f
C702 VN.n24 VSUBS 0.103983f
C703 VN.n25 VSUBS 0.114125f
C704 VN.n26 VSUBS 0.11575f
C705 VN.n27 VSUBS 0.061542f
C706 VN.n28 VSUBS 0.061542f
C707 VN.n29 VSUBS 0.061542f
C708 VN.n30 VSUBS 0.123637f
C709 VN.n31 VSUBS 0.114125f
C710 VN.n32 VSUBS 0.088208f
C711 VN.n33 VSUBS 0.099312f
C712 VN.n34 VSUBS 0.153622f
C713 VN.t0 VSUBS 0.246518f
C714 VN.n35 VSUBS 0.440931f
C715 VN.n36 VSUBS 0.061542f
C716 VN.n37 VSUBS 0.05366f
C717 VN.n38 VSUBS 0.061542f
C718 VN.t1 VSUBS 0.246518f
C719 VN.n39 VSUBS 0.202711f
C720 VN.n40 VSUBS 0.061542f
C721 VN.n41 VSUBS 0.089462f
C722 VN.n42 VSUBS 0.061542f
C723 VN.n43 VSUBS 0.067926f
C724 VN.t4 VSUBS 0.795051f
C725 VN.t5 VSUBS 0.246518f
C726 VN.n44 VSUBS 0.392708f
C727 VN.n45 VSUBS 0.4969f
C728 VN.n46 VSUBS 0.728431f
C729 VN.n47 VSUBS 0.061542f
C730 VN.n48 VSUBS 0.114125f
C731 VN.n49 VSUBS 0.114125f
C732 VN.n50 VSUBS 0.089462f
C733 VN.n51 VSUBS 0.061542f
C734 VN.n52 VSUBS 0.061542f
C735 VN.n53 VSUBS 0.061542f
C736 VN.n54 VSUBS 0.114125f
C737 VN.n55 VSUBS 0.114125f
C738 VN.n56 VSUBS 0.067926f
C739 VN.n57 VSUBS 0.061542f
C740 VN.n58 VSUBS 0.061542f
C741 VN.n59 VSUBS 0.103983f
C742 VN.n60 VSUBS 0.114125f
C743 VN.n61 VSUBS 0.11575f
C744 VN.n62 VSUBS 0.061542f
C745 VN.n63 VSUBS 0.061542f
C746 VN.n64 VSUBS 0.061542f
C747 VN.n65 VSUBS 0.123637f
C748 VN.n66 VSUBS 0.114125f
C749 VN.n67 VSUBS 0.088208f
C750 VN.n68 VSUBS 0.099312f
C751 VN.n69 VSUBS 3.12813f
C752 VTAIL.t13 VSUBS 0.028792f
C753 VTAIL.t1 VSUBS 0.028792f
C754 VTAIL.n0 VSUBS 0.058944f
C755 VTAIL.n1 VSUBS 0.568468f
C756 VTAIL.t0 VSUBS 0.130456f
C757 VTAIL.n2 VSUBS 0.639065f
C758 VTAIL.t7 VSUBS 0.130456f
C759 VTAIL.n3 VSUBS 0.639065f
C760 VTAIL.t9 VSUBS 0.028792f
C761 VTAIL.t8 VSUBS 0.028792f
C762 VTAIL.n4 VSUBS 0.058944f
C763 VTAIL.n5 VSUBS 1.04953f
C764 VTAIL.t6 VSUBS 0.130456f
C765 VTAIL.n6 VSUBS 1.80896f
C766 VTAIL.t15 VSUBS 0.130456f
C767 VTAIL.n7 VSUBS 1.80896f
C768 VTAIL.t4 VSUBS 0.028792f
C769 VTAIL.t3 VSUBS 0.028792f
C770 VTAIL.n8 VSUBS 0.058944f
C771 VTAIL.n9 VSUBS 1.04953f
C772 VTAIL.t2 VSUBS 0.130456f
C773 VTAIL.n10 VSUBS 0.639065f
C774 VTAIL.t5 VSUBS 0.130456f
C775 VTAIL.n11 VSUBS 0.639065f
C776 VTAIL.t11 VSUBS 0.028792f
C777 VTAIL.t12 VSUBS 0.028792f
C778 VTAIL.n12 VSUBS 0.058944f
C779 VTAIL.n13 VSUBS 1.04953f
C780 VTAIL.t10 VSUBS 0.130456f
C781 VTAIL.n14 VSUBS 1.80896f
C782 VTAIL.t14 VSUBS 0.130456f
C783 VTAIL.n15 VSUBS 1.79997f
C784 VDD1.t5 VSUBS 0.01792f
C785 VDD1.t2 VSUBS 0.01792f
C786 VDD1.n0 VSUBS 0.040165f
C787 VDD1.t6 VSUBS 0.01792f
C788 VDD1.t4 VSUBS 0.01792f
C789 VDD1.n1 VSUBS 0.040041f
C790 VDD1.t3 VSUBS 0.01792f
C791 VDD1.t1 VSUBS 0.01792f
C792 VDD1.n2 VSUBS 0.040041f
C793 VDD1.n3 VSUBS 3.37307f
C794 VDD1.t7 VSUBS 0.01792f
C795 VDD1.t0 VSUBS 0.01792f
C796 VDD1.n4 VSUBS 0.038731f
C797 VDD1.n5 VSUBS 2.66416f
C798 VP.t5 VSUBS 0.284747f
C799 VP.n0 VSUBS 0.50931f
C800 VP.n1 VSUBS 0.071086f
C801 VP.n2 VSUBS 0.061982f
C802 VP.n3 VSUBS 0.071086f
C803 VP.t4 VSUBS 0.284747f
C804 VP.n4 VSUBS 0.234146f
C805 VP.n5 VSUBS 0.071086f
C806 VP.n6 VSUBS 0.103335f
C807 VP.n7 VSUBS 0.071086f
C808 VP.n8 VSUBS 0.078459f
C809 VP.n9 VSUBS 0.071086f
C810 VP.n10 VSUBS 0.061982f
C811 VP.n11 VSUBS 0.071086f
C812 VP.t6 VSUBS 0.284747f
C813 VP.n12 VSUBS 0.50931f
C814 VP.t2 VSUBS 0.284747f
C815 VP.n13 VSUBS 0.50931f
C816 VP.n14 VSUBS 0.071086f
C817 VP.n15 VSUBS 0.061982f
C818 VP.n16 VSUBS 0.071086f
C819 VP.t0 VSUBS 0.284747f
C820 VP.n17 VSUBS 0.234146f
C821 VP.n18 VSUBS 0.071086f
C822 VP.n19 VSUBS 0.103335f
C823 VP.n20 VSUBS 0.071086f
C824 VP.n21 VSUBS 0.078459f
C825 VP.t7 VSUBS 0.918343f
C826 VP.t1 VSUBS 0.284747f
C827 VP.n22 VSUBS 0.453608f
C828 VP.n23 VSUBS 0.573958f
C829 VP.n24 VSUBS 0.841395f
C830 VP.n25 VSUBS 0.071086f
C831 VP.n26 VSUBS 0.131823f
C832 VP.n27 VSUBS 0.131823f
C833 VP.n28 VSUBS 0.103335f
C834 VP.n29 VSUBS 0.071086f
C835 VP.n30 VSUBS 0.071086f
C836 VP.n31 VSUBS 0.071086f
C837 VP.n32 VSUBS 0.131823f
C838 VP.n33 VSUBS 0.131823f
C839 VP.n34 VSUBS 0.078459f
C840 VP.n35 VSUBS 0.071086f
C841 VP.n36 VSUBS 0.071086f
C842 VP.n37 VSUBS 0.120109f
C843 VP.n38 VSUBS 0.131823f
C844 VP.n39 VSUBS 0.1337f
C845 VP.n40 VSUBS 0.071086f
C846 VP.n41 VSUBS 0.071086f
C847 VP.n42 VSUBS 0.071086f
C848 VP.n43 VSUBS 0.142811f
C849 VP.n44 VSUBS 0.131823f
C850 VP.n45 VSUBS 0.101887f
C851 VP.n46 VSUBS 0.114714f
C852 VP.n47 VSUBS 3.58329f
C853 VP.n48 VSUBS 3.63901f
C854 VP.n49 VSUBS 0.114714f
C855 VP.n50 VSUBS 0.101887f
C856 VP.n51 VSUBS 0.131823f
C857 VP.n52 VSUBS 0.142811f
C858 VP.n53 VSUBS 0.071086f
C859 VP.n54 VSUBS 0.071086f
C860 VP.n55 VSUBS 0.071086f
C861 VP.n56 VSUBS 0.1337f
C862 VP.n57 VSUBS 0.131823f
C863 VP.t3 VSUBS 0.284747f
C864 VP.n58 VSUBS 0.234146f
C865 VP.n59 VSUBS 0.120109f
C866 VP.n60 VSUBS 0.071086f
C867 VP.n61 VSUBS 0.071086f
C868 VP.n62 VSUBS 0.071086f
C869 VP.n63 VSUBS 0.131823f
C870 VP.n64 VSUBS 0.131823f
C871 VP.n65 VSUBS 0.103335f
C872 VP.n66 VSUBS 0.071086f
C873 VP.n67 VSUBS 0.071086f
C874 VP.n68 VSUBS 0.071086f
C875 VP.n69 VSUBS 0.131823f
C876 VP.n70 VSUBS 0.131823f
C877 VP.n71 VSUBS 0.078459f
C878 VP.n72 VSUBS 0.071086f
C879 VP.n73 VSUBS 0.071086f
C880 VP.n74 VSUBS 0.120109f
C881 VP.n75 VSUBS 0.131823f
C882 VP.n76 VSUBS 0.1337f
C883 VP.n77 VSUBS 0.071086f
C884 VP.n78 VSUBS 0.071086f
C885 VP.n79 VSUBS 0.071086f
C886 VP.n80 VSUBS 0.142811f
C887 VP.n81 VSUBS 0.131823f
C888 VP.n82 VSUBS 0.101887f
C889 VP.n83 VSUBS 0.114714f
C890 VP.n84 VSUBS 0.177445f
.ends

