* NGSPICE file created from diff_pair_sample_1242.ext - technology: sky130A

.subckt diff_pair_sample_1242 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X1 VDD1.t4 VP.t1 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X2 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=0 ps=0 w=15.74 l=1.76
X3 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=0 ps=0 w=15.74 l=1.76
X4 VDD1.t3 VP.t2 VTAIL.t12 B.t23 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=6.1386 ps=32.26 w=15.74 l=1.76
X5 VTAIL.t4 VN.t0 VDD2.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X6 VDD1.t1 VP.t3 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=6.1386 ps=32.26 w=15.74 l=1.76
X7 VDD2.t8 VN.t1 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=2.5971 ps=16.07 w=15.74 l=1.76
X8 VDD2.t7 VN.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X9 VTAIL.t0 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X10 VTAIL.t2 VN.t4 VDD2.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X11 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X12 VTAIL.t16 VN.t6 VDD2.t3 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X13 VTAIL.t10 VP.t4 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X14 VDD2.t2 VN.t7 VTAIL.t18 B.t23 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=6.1386 ps=32.26 w=15.74 l=1.76
X15 VDD1.t9 VP.t5 VTAIL.t9 B.t21 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=2.5971 ps=16.07 w=15.74 l=1.76
X16 VDD1.t8 VP.t6 VTAIL.t8 B.t20 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=2.5971 ps=16.07 w=15.74 l=1.76
X17 VTAIL.t7 VP.t7 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X18 VDD2.t1 VN.t8 VTAIL.t17 B.t20 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=2.5971 ps=16.07 w=15.74 l=1.76
X19 VDD1.t5 VP.t8 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X20 VTAIL.t5 VP.t9 VDD1.t2 B.t19 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=2.5971 ps=16.07 w=15.74 l=1.76
X21 VDD2.t0 VN.t9 VTAIL.t19 B.t22 sky130_fd_pr__nfet_01v8 ad=2.5971 pd=16.07 as=6.1386 ps=32.26 w=15.74 l=1.76
X22 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=0 ps=0 w=15.74 l=1.76
X23 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=6.1386 pd=32.26 as=0 ps=0 w=15.74 l=1.76
R0 VP.n14 VP.t5 246.417
R1 VP.n39 VP.t6 215.531
R2 VP.n46 VP.t4 215.531
R3 VP.n53 VP.t1 215.531
R4 VP.n60 VP.t0 215.531
R5 VP.n67 VP.t2 215.531
R6 VP.n36 VP.t3 215.531
R7 VP.n29 VP.t7 215.531
R8 VP.n22 VP.t8 215.531
R9 VP.n15 VP.t9 215.531
R10 VP.n17 VP.n16 161.3
R11 VP.n18 VP.n13 161.3
R12 VP.n20 VP.n19 161.3
R13 VP.n21 VP.n12 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n25 VP.n11 161.3
R16 VP.n27 VP.n26 161.3
R17 VP.n28 VP.n10 161.3
R18 VP.n31 VP.n30 161.3
R19 VP.n32 VP.n9 161.3
R20 VP.n34 VP.n33 161.3
R21 VP.n35 VP.n8 161.3
R22 VP.n66 VP.n0 161.3
R23 VP.n65 VP.n64 161.3
R24 VP.n63 VP.n1 161.3
R25 VP.n62 VP.n61 161.3
R26 VP.n59 VP.n2 161.3
R27 VP.n58 VP.n57 161.3
R28 VP.n56 VP.n3 161.3
R29 VP.n55 VP.n54 161.3
R30 VP.n52 VP.n4 161.3
R31 VP.n51 VP.n50 161.3
R32 VP.n49 VP.n5 161.3
R33 VP.n48 VP.n47 161.3
R34 VP.n45 VP.n6 161.3
R35 VP.n44 VP.n43 161.3
R36 VP.n42 VP.n7 161.3
R37 VP.n41 VP.n40 161.3
R38 VP.n39 VP.n38 89.6708
R39 VP.n68 VP.n67 89.6708
R40 VP.n37 VP.n36 89.6708
R41 VP.n51 VP.n5 56.4773
R42 VP.n58 VP.n3 56.4773
R43 VP.n27 VP.n11 56.4773
R44 VP.n20 VP.n13 56.4773
R45 VP.n15 VP.n14 52.8339
R46 VP.n44 VP.n7 51.6086
R47 VP.n65 VP.n1 51.6086
R48 VP.n34 VP.n9 51.6086
R49 VP.n38 VP.n37 51.3669
R50 VP.n40 VP.n7 29.2126
R51 VP.n66 VP.n65 29.2126
R52 VP.n35 VP.n34 29.2126
R53 VP.n45 VP.n44 24.3439
R54 VP.n47 VP.n5 24.3439
R55 VP.n52 VP.n51 24.3439
R56 VP.n54 VP.n3 24.3439
R57 VP.n59 VP.n58 24.3439
R58 VP.n61 VP.n1 24.3439
R59 VP.n28 VP.n27 24.3439
R60 VP.n30 VP.n9 24.3439
R61 VP.n21 VP.n20 24.3439
R62 VP.n23 VP.n11 24.3439
R63 VP.n16 VP.n13 24.3439
R64 VP.n40 VP.n39 20.9359
R65 VP.n67 VP.n66 20.9359
R66 VP.n36 VP.n35 20.9359
R67 VP.n47 VP.n46 16.554
R68 VP.n60 VP.n59 16.554
R69 VP.n29 VP.n28 16.554
R70 VP.n16 VP.n15 16.554
R71 VP.n17 VP.n14 13.1234
R72 VP.n53 VP.n52 12.1722
R73 VP.n54 VP.n53 12.1722
R74 VP.n22 VP.n21 12.1722
R75 VP.n23 VP.n22 12.1722
R76 VP.n46 VP.n45 7.7904
R77 VP.n61 VP.n60 7.7904
R78 VP.n30 VP.n29 7.7904
R79 VP.n37 VP.n8 0.278398
R80 VP.n41 VP.n38 0.278398
R81 VP.n68 VP.n0 0.278398
R82 VP.n18 VP.n17 0.189894
R83 VP.n19 VP.n18 0.189894
R84 VP.n19 VP.n12 0.189894
R85 VP.n24 VP.n12 0.189894
R86 VP.n25 VP.n24 0.189894
R87 VP.n26 VP.n25 0.189894
R88 VP.n26 VP.n10 0.189894
R89 VP.n31 VP.n10 0.189894
R90 VP.n32 VP.n31 0.189894
R91 VP.n33 VP.n32 0.189894
R92 VP.n33 VP.n8 0.189894
R93 VP.n42 VP.n41 0.189894
R94 VP.n43 VP.n42 0.189894
R95 VP.n43 VP.n6 0.189894
R96 VP.n48 VP.n6 0.189894
R97 VP.n49 VP.n48 0.189894
R98 VP.n50 VP.n49 0.189894
R99 VP.n50 VP.n4 0.189894
R100 VP.n55 VP.n4 0.189894
R101 VP.n56 VP.n55 0.189894
R102 VP.n57 VP.n56 0.189894
R103 VP.n57 VP.n2 0.189894
R104 VP.n62 VP.n2 0.189894
R105 VP.n63 VP.n62 0.189894
R106 VP.n64 VP.n63 0.189894
R107 VP.n64 VP.n0 0.189894
R108 VP VP.n68 0.153422
R109 VDD1.n1 VDD1.t9 64.2558
R110 VDD1.n3 VDD1.t8 64.2557
R111 VDD1.n5 VDD1.n4 62.4919
R112 VDD1.n1 VDD1.n0 61.1962
R113 VDD1.n7 VDD1.n6 61.196
R114 VDD1.n3 VDD1.n2 61.1959
R115 VDD1.n7 VDD1.n5 47.3263
R116 VDD1 VDD1.n7 1.2936
R117 VDD1.n6 VDD1.t6 1.25844
R118 VDD1.n6 VDD1.t1 1.25844
R119 VDD1.n0 VDD1.t2 1.25844
R120 VDD1.n0 VDD1.t5 1.25844
R121 VDD1.n4 VDD1.t7 1.25844
R122 VDD1.n4 VDD1.t3 1.25844
R123 VDD1.n2 VDD1.t0 1.25844
R124 VDD1.n2 VDD1.t4 1.25844
R125 VDD1 VDD1.n1 0.509121
R126 VDD1.n5 VDD1.n3 0.395585
R127 VTAIL.n11 VTAIL.t18 45.7753
R128 VTAIL.n17 VTAIL.t19 45.7752
R129 VTAIL.n2 VTAIL.t12 45.7752
R130 VTAIL.n16 VTAIL.t11 45.7752
R131 VTAIL.n15 VTAIL.n14 44.5174
R132 VTAIL.n13 VTAIL.n12 44.5174
R133 VTAIL.n10 VTAIL.n9 44.5174
R134 VTAIL.n8 VTAIL.n7 44.5174
R135 VTAIL.n19 VTAIL.n18 44.5171
R136 VTAIL.n1 VTAIL.n0 44.5171
R137 VTAIL.n4 VTAIL.n3 44.5171
R138 VTAIL.n6 VTAIL.n5 44.5171
R139 VTAIL.n8 VTAIL.n6 29.5393
R140 VTAIL.n17 VTAIL.n16 27.7376
R141 VTAIL.n10 VTAIL.n8 1.80222
R142 VTAIL.n11 VTAIL.n10 1.80222
R143 VTAIL.n15 VTAIL.n13 1.80222
R144 VTAIL.n16 VTAIL.n15 1.80222
R145 VTAIL.n6 VTAIL.n4 1.80222
R146 VTAIL.n4 VTAIL.n2 1.80222
R147 VTAIL.n19 VTAIL.n17 1.80222
R148 VTAIL VTAIL.n1 1.40998
R149 VTAIL.n13 VTAIL.n11 1.37119
R150 VTAIL.n2 VTAIL.n1 1.37119
R151 VTAIL.n18 VTAIL.t1 1.25844
R152 VTAIL.n18 VTAIL.t4 1.25844
R153 VTAIL.n0 VTAIL.t15 1.25844
R154 VTAIL.n0 VTAIL.t16 1.25844
R155 VTAIL.n3 VTAIL.t13 1.25844
R156 VTAIL.n3 VTAIL.t14 1.25844
R157 VTAIL.n5 VTAIL.t8 1.25844
R158 VTAIL.n5 VTAIL.t10 1.25844
R159 VTAIL.n14 VTAIL.t6 1.25844
R160 VTAIL.n14 VTAIL.t7 1.25844
R161 VTAIL.n12 VTAIL.t9 1.25844
R162 VTAIL.n12 VTAIL.t5 1.25844
R163 VTAIL.n9 VTAIL.t3 1.25844
R164 VTAIL.n9 VTAIL.t2 1.25844
R165 VTAIL.n7 VTAIL.t17 1.25844
R166 VTAIL.n7 VTAIL.t0 1.25844
R167 VTAIL VTAIL.n19 0.392741
R168 B.n949 B.n948 585
R169 B.n950 B.n949 585
R170 B.n374 B.n141 585
R171 B.n373 B.n372 585
R172 B.n371 B.n370 585
R173 B.n369 B.n368 585
R174 B.n367 B.n366 585
R175 B.n365 B.n364 585
R176 B.n363 B.n362 585
R177 B.n361 B.n360 585
R178 B.n359 B.n358 585
R179 B.n357 B.n356 585
R180 B.n355 B.n354 585
R181 B.n353 B.n352 585
R182 B.n351 B.n350 585
R183 B.n349 B.n348 585
R184 B.n347 B.n346 585
R185 B.n345 B.n344 585
R186 B.n343 B.n342 585
R187 B.n341 B.n340 585
R188 B.n339 B.n338 585
R189 B.n337 B.n336 585
R190 B.n335 B.n334 585
R191 B.n333 B.n332 585
R192 B.n331 B.n330 585
R193 B.n329 B.n328 585
R194 B.n327 B.n326 585
R195 B.n325 B.n324 585
R196 B.n323 B.n322 585
R197 B.n321 B.n320 585
R198 B.n319 B.n318 585
R199 B.n317 B.n316 585
R200 B.n315 B.n314 585
R201 B.n313 B.n312 585
R202 B.n311 B.n310 585
R203 B.n309 B.n308 585
R204 B.n307 B.n306 585
R205 B.n305 B.n304 585
R206 B.n303 B.n302 585
R207 B.n301 B.n300 585
R208 B.n299 B.n298 585
R209 B.n297 B.n296 585
R210 B.n295 B.n294 585
R211 B.n293 B.n292 585
R212 B.n291 B.n290 585
R213 B.n289 B.n288 585
R214 B.n287 B.n286 585
R215 B.n285 B.n284 585
R216 B.n283 B.n282 585
R217 B.n281 B.n280 585
R218 B.n279 B.n278 585
R219 B.n277 B.n276 585
R220 B.n275 B.n274 585
R221 B.n273 B.n272 585
R222 B.n271 B.n270 585
R223 B.n269 B.n268 585
R224 B.n267 B.n266 585
R225 B.n265 B.n264 585
R226 B.n263 B.n262 585
R227 B.n261 B.n260 585
R228 B.n259 B.n258 585
R229 B.n257 B.n256 585
R230 B.n255 B.n254 585
R231 B.n252 B.n251 585
R232 B.n250 B.n249 585
R233 B.n248 B.n247 585
R234 B.n246 B.n245 585
R235 B.n244 B.n243 585
R236 B.n242 B.n241 585
R237 B.n240 B.n239 585
R238 B.n238 B.n237 585
R239 B.n236 B.n235 585
R240 B.n234 B.n233 585
R241 B.n232 B.n231 585
R242 B.n230 B.n229 585
R243 B.n228 B.n227 585
R244 B.n226 B.n225 585
R245 B.n224 B.n223 585
R246 B.n222 B.n221 585
R247 B.n220 B.n219 585
R248 B.n218 B.n217 585
R249 B.n216 B.n215 585
R250 B.n214 B.n213 585
R251 B.n212 B.n211 585
R252 B.n210 B.n209 585
R253 B.n208 B.n207 585
R254 B.n206 B.n205 585
R255 B.n204 B.n203 585
R256 B.n202 B.n201 585
R257 B.n200 B.n199 585
R258 B.n198 B.n197 585
R259 B.n196 B.n195 585
R260 B.n194 B.n193 585
R261 B.n192 B.n191 585
R262 B.n190 B.n189 585
R263 B.n188 B.n187 585
R264 B.n186 B.n185 585
R265 B.n184 B.n183 585
R266 B.n182 B.n181 585
R267 B.n180 B.n179 585
R268 B.n178 B.n177 585
R269 B.n176 B.n175 585
R270 B.n174 B.n173 585
R271 B.n172 B.n171 585
R272 B.n170 B.n169 585
R273 B.n168 B.n167 585
R274 B.n166 B.n165 585
R275 B.n164 B.n163 585
R276 B.n162 B.n161 585
R277 B.n160 B.n159 585
R278 B.n158 B.n157 585
R279 B.n156 B.n155 585
R280 B.n154 B.n153 585
R281 B.n152 B.n151 585
R282 B.n150 B.n149 585
R283 B.n148 B.n147 585
R284 B.n947 B.n83 585
R285 B.n951 B.n83 585
R286 B.n946 B.n82 585
R287 B.n952 B.n82 585
R288 B.n945 B.n944 585
R289 B.n944 B.n78 585
R290 B.n943 B.n77 585
R291 B.n958 B.n77 585
R292 B.n942 B.n76 585
R293 B.n959 B.n76 585
R294 B.n941 B.n75 585
R295 B.n960 B.n75 585
R296 B.n940 B.n939 585
R297 B.n939 B.n74 585
R298 B.n938 B.n70 585
R299 B.n966 B.n70 585
R300 B.n937 B.n69 585
R301 B.n967 B.n69 585
R302 B.n936 B.n68 585
R303 B.n968 B.n68 585
R304 B.n935 B.n934 585
R305 B.n934 B.n64 585
R306 B.n933 B.n63 585
R307 B.n974 B.n63 585
R308 B.n932 B.n62 585
R309 B.n975 B.n62 585
R310 B.n931 B.n61 585
R311 B.n976 B.n61 585
R312 B.n930 B.n929 585
R313 B.n929 B.n57 585
R314 B.n928 B.n56 585
R315 B.n982 B.n56 585
R316 B.n927 B.n55 585
R317 B.n983 B.n55 585
R318 B.n926 B.n54 585
R319 B.n984 B.n54 585
R320 B.n925 B.n924 585
R321 B.n924 B.n50 585
R322 B.n923 B.n49 585
R323 B.n990 B.n49 585
R324 B.n922 B.n48 585
R325 B.n991 B.n48 585
R326 B.n921 B.n47 585
R327 B.n992 B.n47 585
R328 B.n920 B.n919 585
R329 B.n919 B.n43 585
R330 B.n918 B.n42 585
R331 B.n998 B.n42 585
R332 B.n917 B.n41 585
R333 B.n999 B.n41 585
R334 B.n916 B.n40 585
R335 B.n1000 B.n40 585
R336 B.n915 B.n914 585
R337 B.n914 B.n36 585
R338 B.n913 B.n35 585
R339 B.n1006 B.n35 585
R340 B.n912 B.n34 585
R341 B.n1007 B.n34 585
R342 B.n911 B.n33 585
R343 B.n1008 B.n33 585
R344 B.n910 B.n909 585
R345 B.n909 B.n29 585
R346 B.n908 B.n28 585
R347 B.n1014 B.n28 585
R348 B.n907 B.n27 585
R349 B.n1015 B.n27 585
R350 B.n906 B.n26 585
R351 B.n1016 B.n26 585
R352 B.n905 B.n904 585
R353 B.n904 B.n25 585
R354 B.n903 B.n21 585
R355 B.n1022 B.n21 585
R356 B.n902 B.n20 585
R357 B.n1023 B.n20 585
R358 B.n901 B.n19 585
R359 B.n1024 B.n19 585
R360 B.n900 B.n899 585
R361 B.n899 B.n15 585
R362 B.n898 B.n14 585
R363 B.n1030 B.n14 585
R364 B.n897 B.n13 585
R365 B.n1031 B.n13 585
R366 B.n896 B.n12 585
R367 B.n1032 B.n12 585
R368 B.n895 B.n894 585
R369 B.n894 B.n8 585
R370 B.n893 B.n7 585
R371 B.n1038 B.n7 585
R372 B.n892 B.n6 585
R373 B.n1039 B.n6 585
R374 B.n891 B.n5 585
R375 B.n1040 B.n5 585
R376 B.n890 B.n889 585
R377 B.n889 B.n4 585
R378 B.n888 B.n375 585
R379 B.n888 B.n887 585
R380 B.n878 B.n376 585
R381 B.n377 B.n376 585
R382 B.n880 B.n879 585
R383 B.n881 B.n880 585
R384 B.n877 B.n381 585
R385 B.n385 B.n381 585
R386 B.n876 B.n875 585
R387 B.n875 B.n874 585
R388 B.n383 B.n382 585
R389 B.n384 B.n383 585
R390 B.n867 B.n866 585
R391 B.n868 B.n867 585
R392 B.n865 B.n390 585
R393 B.n390 B.n389 585
R394 B.n864 B.n863 585
R395 B.n863 B.n862 585
R396 B.n392 B.n391 585
R397 B.n855 B.n392 585
R398 B.n854 B.n853 585
R399 B.n856 B.n854 585
R400 B.n852 B.n397 585
R401 B.n397 B.n396 585
R402 B.n851 B.n850 585
R403 B.n850 B.n849 585
R404 B.n399 B.n398 585
R405 B.n400 B.n399 585
R406 B.n842 B.n841 585
R407 B.n843 B.n842 585
R408 B.n840 B.n404 585
R409 B.n408 B.n404 585
R410 B.n839 B.n838 585
R411 B.n838 B.n837 585
R412 B.n406 B.n405 585
R413 B.n407 B.n406 585
R414 B.n830 B.n829 585
R415 B.n831 B.n830 585
R416 B.n828 B.n413 585
R417 B.n413 B.n412 585
R418 B.n827 B.n826 585
R419 B.n826 B.n825 585
R420 B.n415 B.n414 585
R421 B.n416 B.n415 585
R422 B.n818 B.n817 585
R423 B.n819 B.n818 585
R424 B.n816 B.n421 585
R425 B.n421 B.n420 585
R426 B.n815 B.n814 585
R427 B.n814 B.n813 585
R428 B.n423 B.n422 585
R429 B.n424 B.n423 585
R430 B.n806 B.n805 585
R431 B.n807 B.n806 585
R432 B.n804 B.n429 585
R433 B.n429 B.n428 585
R434 B.n803 B.n802 585
R435 B.n802 B.n801 585
R436 B.n431 B.n430 585
R437 B.n432 B.n431 585
R438 B.n794 B.n793 585
R439 B.n795 B.n794 585
R440 B.n792 B.n437 585
R441 B.n437 B.n436 585
R442 B.n791 B.n790 585
R443 B.n790 B.n789 585
R444 B.n439 B.n438 585
R445 B.n440 B.n439 585
R446 B.n782 B.n781 585
R447 B.n783 B.n782 585
R448 B.n780 B.n445 585
R449 B.n445 B.n444 585
R450 B.n779 B.n778 585
R451 B.n778 B.n777 585
R452 B.n447 B.n446 585
R453 B.n770 B.n447 585
R454 B.n769 B.n768 585
R455 B.n771 B.n769 585
R456 B.n767 B.n452 585
R457 B.n452 B.n451 585
R458 B.n766 B.n765 585
R459 B.n765 B.n764 585
R460 B.n454 B.n453 585
R461 B.n455 B.n454 585
R462 B.n757 B.n756 585
R463 B.n758 B.n757 585
R464 B.n755 B.n460 585
R465 B.n460 B.n459 585
R466 B.n749 B.n748 585
R467 B.n747 B.n519 585
R468 B.n746 B.n518 585
R469 B.n751 B.n518 585
R470 B.n745 B.n744 585
R471 B.n743 B.n742 585
R472 B.n741 B.n740 585
R473 B.n739 B.n738 585
R474 B.n737 B.n736 585
R475 B.n735 B.n734 585
R476 B.n733 B.n732 585
R477 B.n731 B.n730 585
R478 B.n729 B.n728 585
R479 B.n727 B.n726 585
R480 B.n725 B.n724 585
R481 B.n723 B.n722 585
R482 B.n721 B.n720 585
R483 B.n719 B.n718 585
R484 B.n717 B.n716 585
R485 B.n715 B.n714 585
R486 B.n713 B.n712 585
R487 B.n711 B.n710 585
R488 B.n709 B.n708 585
R489 B.n707 B.n706 585
R490 B.n705 B.n704 585
R491 B.n703 B.n702 585
R492 B.n701 B.n700 585
R493 B.n699 B.n698 585
R494 B.n697 B.n696 585
R495 B.n695 B.n694 585
R496 B.n693 B.n692 585
R497 B.n691 B.n690 585
R498 B.n689 B.n688 585
R499 B.n687 B.n686 585
R500 B.n685 B.n684 585
R501 B.n683 B.n682 585
R502 B.n681 B.n680 585
R503 B.n679 B.n678 585
R504 B.n677 B.n676 585
R505 B.n675 B.n674 585
R506 B.n673 B.n672 585
R507 B.n671 B.n670 585
R508 B.n669 B.n668 585
R509 B.n667 B.n666 585
R510 B.n665 B.n664 585
R511 B.n663 B.n662 585
R512 B.n661 B.n660 585
R513 B.n659 B.n658 585
R514 B.n657 B.n656 585
R515 B.n655 B.n654 585
R516 B.n653 B.n652 585
R517 B.n651 B.n650 585
R518 B.n649 B.n648 585
R519 B.n647 B.n646 585
R520 B.n645 B.n644 585
R521 B.n643 B.n642 585
R522 B.n641 B.n640 585
R523 B.n639 B.n638 585
R524 B.n637 B.n636 585
R525 B.n635 B.n634 585
R526 B.n633 B.n632 585
R527 B.n631 B.n630 585
R528 B.n629 B.n628 585
R529 B.n626 B.n625 585
R530 B.n624 B.n623 585
R531 B.n622 B.n621 585
R532 B.n620 B.n619 585
R533 B.n618 B.n617 585
R534 B.n616 B.n615 585
R535 B.n614 B.n613 585
R536 B.n612 B.n611 585
R537 B.n610 B.n609 585
R538 B.n608 B.n607 585
R539 B.n606 B.n605 585
R540 B.n604 B.n603 585
R541 B.n602 B.n601 585
R542 B.n600 B.n599 585
R543 B.n598 B.n597 585
R544 B.n596 B.n595 585
R545 B.n594 B.n593 585
R546 B.n592 B.n591 585
R547 B.n590 B.n589 585
R548 B.n588 B.n587 585
R549 B.n586 B.n585 585
R550 B.n584 B.n583 585
R551 B.n582 B.n581 585
R552 B.n580 B.n579 585
R553 B.n578 B.n577 585
R554 B.n576 B.n575 585
R555 B.n574 B.n573 585
R556 B.n572 B.n571 585
R557 B.n570 B.n569 585
R558 B.n568 B.n567 585
R559 B.n566 B.n565 585
R560 B.n564 B.n563 585
R561 B.n562 B.n561 585
R562 B.n560 B.n559 585
R563 B.n558 B.n557 585
R564 B.n556 B.n555 585
R565 B.n554 B.n553 585
R566 B.n552 B.n551 585
R567 B.n550 B.n549 585
R568 B.n548 B.n547 585
R569 B.n546 B.n545 585
R570 B.n544 B.n543 585
R571 B.n542 B.n541 585
R572 B.n540 B.n539 585
R573 B.n538 B.n537 585
R574 B.n536 B.n535 585
R575 B.n534 B.n533 585
R576 B.n532 B.n531 585
R577 B.n530 B.n529 585
R578 B.n528 B.n527 585
R579 B.n526 B.n525 585
R580 B.n462 B.n461 585
R581 B.n754 B.n753 585
R582 B.n458 B.n457 585
R583 B.n459 B.n458 585
R584 B.n760 B.n759 585
R585 B.n759 B.n758 585
R586 B.n761 B.n456 585
R587 B.n456 B.n455 585
R588 B.n763 B.n762 585
R589 B.n764 B.n763 585
R590 B.n450 B.n449 585
R591 B.n451 B.n450 585
R592 B.n773 B.n772 585
R593 B.n772 B.n771 585
R594 B.n774 B.n448 585
R595 B.n770 B.n448 585
R596 B.n776 B.n775 585
R597 B.n777 B.n776 585
R598 B.n443 B.n442 585
R599 B.n444 B.n443 585
R600 B.n785 B.n784 585
R601 B.n784 B.n783 585
R602 B.n786 B.n441 585
R603 B.n441 B.n440 585
R604 B.n788 B.n787 585
R605 B.n789 B.n788 585
R606 B.n435 B.n434 585
R607 B.n436 B.n435 585
R608 B.n797 B.n796 585
R609 B.n796 B.n795 585
R610 B.n798 B.n433 585
R611 B.n433 B.n432 585
R612 B.n800 B.n799 585
R613 B.n801 B.n800 585
R614 B.n427 B.n426 585
R615 B.n428 B.n427 585
R616 B.n809 B.n808 585
R617 B.n808 B.n807 585
R618 B.n810 B.n425 585
R619 B.n425 B.n424 585
R620 B.n812 B.n811 585
R621 B.n813 B.n812 585
R622 B.n419 B.n418 585
R623 B.n420 B.n419 585
R624 B.n821 B.n820 585
R625 B.n820 B.n819 585
R626 B.n822 B.n417 585
R627 B.n417 B.n416 585
R628 B.n824 B.n823 585
R629 B.n825 B.n824 585
R630 B.n411 B.n410 585
R631 B.n412 B.n411 585
R632 B.n833 B.n832 585
R633 B.n832 B.n831 585
R634 B.n834 B.n409 585
R635 B.n409 B.n407 585
R636 B.n836 B.n835 585
R637 B.n837 B.n836 585
R638 B.n403 B.n402 585
R639 B.n408 B.n403 585
R640 B.n845 B.n844 585
R641 B.n844 B.n843 585
R642 B.n846 B.n401 585
R643 B.n401 B.n400 585
R644 B.n848 B.n847 585
R645 B.n849 B.n848 585
R646 B.n395 B.n394 585
R647 B.n396 B.n395 585
R648 B.n858 B.n857 585
R649 B.n857 B.n856 585
R650 B.n859 B.n393 585
R651 B.n855 B.n393 585
R652 B.n861 B.n860 585
R653 B.n862 B.n861 585
R654 B.n388 B.n387 585
R655 B.n389 B.n388 585
R656 B.n870 B.n869 585
R657 B.n869 B.n868 585
R658 B.n871 B.n386 585
R659 B.n386 B.n384 585
R660 B.n873 B.n872 585
R661 B.n874 B.n873 585
R662 B.n380 B.n379 585
R663 B.n385 B.n380 585
R664 B.n883 B.n882 585
R665 B.n882 B.n881 585
R666 B.n884 B.n378 585
R667 B.n378 B.n377 585
R668 B.n886 B.n885 585
R669 B.n887 B.n886 585
R670 B.n2 B.n0 585
R671 B.n4 B.n2 585
R672 B.n3 B.n1 585
R673 B.n1039 B.n3 585
R674 B.n1037 B.n1036 585
R675 B.n1038 B.n1037 585
R676 B.n1035 B.n9 585
R677 B.n9 B.n8 585
R678 B.n1034 B.n1033 585
R679 B.n1033 B.n1032 585
R680 B.n11 B.n10 585
R681 B.n1031 B.n11 585
R682 B.n1029 B.n1028 585
R683 B.n1030 B.n1029 585
R684 B.n1027 B.n16 585
R685 B.n16 B.n15 585
R686 B.n1026 B.n1025 585
R687 B.n1025 B.n1024 585
R688 B.n18 B.n17 585
R689 B.n1023 B.n18 585
R690 B.n1021 B.n1020 585
R691 B.n1022 B.n1021 585
R692 B.n1019 B.n22 585
R693 B.n25 B.n22 585
R694 B.n1018 B.n1017 585
R695 B.n1017 B.n1016 585
R696 B.n24 B.n23 585
R697 B.n1015 B.n24 585
R698 B.n1013 B.n1012 585
R699 B.n1014 B.n1013 585
R700 B.n1011 B.n30 585
R701 B.n30 B.n29 585
R702 B.n1010 B.n1009 585
R703 B.n1009 B.n1008 585
R704 B.n32 B.n31 585
R705 B.n1007 B.n32 585
R706 B.n1005 B.n1004 585
R707 B.n1006 B.n1005 585
R708 B.n1003 B.n37 585
R709 B.n37 B.n36 585
R710 B.n1002 B.n1001 585
R711 B.n1001 B.n1000 585
R712 B.n39 B.n38 585
R713 B.n999 B.n39 585
R714 B.n997 B.n996 585
R715 B.n998 B.n997 585
R716 B.n995 B.n44 585
R717 B.n44 B.n43 585
R718 B.n994 B.n993 585
R719 B.n993 B.n992 585
R720 B.n46 B.n45 585
R721 B.n991 B.n46 585
R722 B.n989 B.n988 585
R723 B.n990 B.n989 585
R724 B.n987 B.n51 585
R725 B.n51 B.n50 585
R726 B.n986 B.n985 585
R727 B.n985 B.n984 585
R728 B.n53 B.n52 585
R729 B.n983 B.n53 585
R730 B.n981 B.n980 585
R731 B.n982 B.n981 585
R732 B.n979 B.n58 585
R733 B.n58 B.n57 585
R734 B.n978 B.n977 585
R735 B.n977 B.n976 585
R736 B.n60 B.n59 585
R737 B.n975 B.n60 585
R738 B.n973 B.n972 585
R739 B.n974 B.n973 585
R740 B.n971 B.n65 585
R741 B.n65 B.n64 585
R742 B.n970 B.n969 585
R743 B.n969 B.n968 585
R744 B.n67 B.n66 585
R745 B.n967 B.n67 585
R746 B.n965 B.n964 585
R747 B.n966 B.n965 585
R748 B.n963 B.n71 585
R749 B.n74 B.n71 585
R750 B.n962 B.n961 585
R751 B.n961 B.n960 585
R752 B.n73 B.n72 585
R753 B.n959 B.n73 585
R754 B.n957 B.n956 585
R755 B.n958 B.n957 585
R756 B.n955 B.n79 585
R757 B.n79 B.n78 585
R758 B.n954 B.n953 585
R759 B.n953 B.n952 585
R760 B.n81 B.n80 585
R761 B.n951 B.n81 585
R762 B.n1042 B.n1041 585
R763 B.n1041 B.n1040 585
R764 B.n749 B.n458 482.89
R765 B.n147 B.n81 482.89
R766 B.n753 B.n460 482.89
R767 B.n949 B.n83 482.89
R768 B.n523 B.t13 422.471
R769 B.n142 B.t5 422.471
R770 B.n520 B.t9 422.045
R771 B.n145 B.t16 422.045
R772 B.n950 B.n140 256.663
R773 B.n950 B.n139 256.663
R774 B.n950 B.n138 256.663
R775 B.n950 B.n137 256.663
R776 B.n950 B.n136 256.663
R777 B.n950 B.n135 256.663
R778 B.n950 B.n134 256.663
R779 B.n950 B.n133 256.663
R780 B.n950 B.n132 256.663
R781 B.n950 B.n131 256.663
R782 B.n950 B.n130 256.663
R783 B.n950 B.n129 256.663
R784 B.n950 B.n128 256.663
R785 B.n950 B.n127 256.663
R786 B.n950 B.n126 256.663
R787 B.n950 B.n125 256.663
R788 B.n950 B.n124 256.663
R789 B.n950 B.n123 256.663
R790 B.n950 B.n122 256.663
R791 B.n950 B.n121 256.663
R792 B.n950 B.n120 256.663
R793 B.n950 B.n119 256.663
R794 B.n950 B.n118 256.663
R795 B.n950 B.n117 256.663
R796 B.n950 B.n116 256.663
R797 B.n950 B.n115 256.663
R798 B.n950 B.n114 256.663
R799 B.n950 B.n113 256.663
R800 B.n950 B.n112 256.663
R801 B.n950 B.n111 256.663
R802 B.n950 B.n110 256.663
R803 B.n950 B.n109 256.663
R804 B.n950 B.n108 256.663
R805 B.n950 B.n107 256.663
R806 B.n950 B.n106 256.663
R807 B.n950 B.n105 256.663
R808 B.n950 B.n104 256.663
R809 B.n950 B.n103 256.663
R810 B.n950 B.n102 256.663
R811 B.n950 B.n101 256.663
R812 B.n950 B.n100 256.663
R813 B.n950 B.n99 256.663
R814 B.n950 B.n98 256.663
R815 B.n950 B.n97 256.663
R816 B.n950 B.n96 256.663
R817 B.n950 B.n95 256.663
R818 B.n950 B.n94 256.663
R819 B.n950 B.n93 256.663
R820 B.n950 B.n92 256.663
R821 B.n950 B.n91 256.663
R822 B.n950 B.n90 256.663
R823 B.n950 B.n89 256.663
R824 B.n950 B.n88 256.663
R825 B.n950 B.n87 256.663
R826 B.n950 B.n86 256.663
R827 B.n950 B.n85 256.663
R828 B.n950 B.n84 256.663
R829 B.n751 B.n750 256.663
R830 B.n751 B.n463 256.663
R831 B.n751 B.n464 256.663
R832 B.n751 B.n465 256.663
R833 B.n751 B.n466 256.663
R834 B.n751 B.n467 256.663
R835 B.n751 B.n468 256.663
R836 B.n751 B.n469 256.663
R837 B.n751 B.n470 256.663
R838 B.n751 B.n471 256.663
R839 B.n751 B.n472 256.663
R840 B.n751 B.n473 256.663
R841 B.n751 B.n474 256.663
R842 B.n751 B.n475 256.663
R843 B.n751 B.n476 256.663
R844 B.n751 B.n477 256.663
R845 B.n751 B.n478 256.663
R846 B.n751 B.n479 256.663
R847 B.n751 B.n480 256.663
R848 B.n751 B.n481 256.663
R849 B.n751 B.n482 256.663
R850 B.n751 B.n483 256.663
R851 B.n751 B.n484 256.663
R852 B.n751 B.n485 256.663
R853 B.n751 B.n486 256.663
R854 B.n751 B.n487 256.663
R855 B.n751 B.n488 256.663
R856 B.n751 B.n489 256.663
R857 B.n751 B.n490 256.663
R858 B.n751 B.n491 256.663
R859 B.n751 B.n492 256.663
R860 B.n751 B.n493 256.663
R861 B.n751 B.n494 256.663
R862 B.n751 B.n495 256.663
R863 B.n751 B.n496 256.663
R864 B.n751 B.n497 256.663
R865 B.n751 B.n498 256.663
R866 B.n751 B.n499 256.663
R867 B.n751 B.n500 256.663
R868 B.n751 B.n501 256.663
R869 B.n751 B.n502 256.663
R870 B.n751 B.n503 256.663
R871 B.n751 B.n504 256.663
R872 B.n751 B.n505 256.663
R873 B.n751 B.n506 256.663
R874 B.n751 B.n507 256.663
R875 B.n751 B.n508 256.663
R876 B.n751 B.n509 256.663
R877 B.n751 B.n510 256.663
R878 B.n751 B.n511 256.663
R879 B.n751 B.n512 256.663
R880 B.n751 B.n513 256.663
R881 B.n751 B.n514 256.663
R882 B.n751 B.n515 256.663
R883 B.n751 B.n516 256.663
R884 B.n751 B.n517 256.663
R885 B.n752 B.n751 256.663
R886 B.n759 B.n458 163.367
R887 B.n759 B.n456 163.367
R888 B.n763 B.n456 163.367
R889 B.n763 B.n450 163.367
R890 B.n772 B.n450 163.367
R891 B.n772 B.n448 163.367
R892 B.n776 B.n448 163.367
R893 B.n776 B.n443 163.367
R894 B.n784 B.n443 163.367
R895 B.n784 B.n441 163.367
R896 B.n788 B.n441 163.367
R897 B.n788 B.n435 163.367
R898 B.n796 B.n435 163.367
R899 B.n796 B.n433 163.367
R900 B.n800 B.n433 163.367
R901 B.n800 B.n427 163.367
R902 B.n808 B.n427 163.367
R903 B.n808 B.n425 163.367
R904 B.n812 B.n425 163.367
R905 B.n812 B.n419 163.367
R906 B.n820 B.n419 163.367
R907 B.n820 B.n417 163.367
R908 B.n824 B.n417 163.367
R909 B.n824 B.n411 163.367
R910 B.n832 B.n411 163.367
R911 B.n832 B.n409 163.367
R912 B.n836 B.n409 163.367
R913 B.n836 B.n403 163.367
R914 B.n844 B.n403 163.367
R915 B.n844 B.n401 163.367
R916 B.n848 B.n401 163.367
R917 B.n848 B.n395 163.367
R918 B.n857 B.n395 163.367
R919 B.n857 B.n393 163.367
R920 B.n861 B.n393 163.367
R921 B.n861 B.n388 163.367
R922 B.n869 B.n388 163.367
R923 B.n869 B.n386 163.367
R924 B.n873 B.n386 163.367
R925 B.n873 B.n380 163.367
R926 B.n882 B.n380 163.367
R927 B.n882 B.n378 163.367
R928 B.n886 B.n378 163.367
R929 B.n886 B.n2 163.367
R930 B.n1041 B.n2 163.367
R931 B.n1041 B.n3 163.367
R932 B.n1037 B.n3 163.367
R933 B.n1037 B.n9 163.367
R934 B.n1033 B.n9 163.367
R935 B.n1033 B.n11 163.367
R936 B.n1029 B.n11 163.367
R937 B.n1029 B.n16 163.367
R938 B.n1025 B.n16 163.367
R939 B.n1025 B.n18 163.367
R940 B.n1021 B.n18 163.367
R941 B.n1021 B.n22 163.367
R942 B.n1017 B.n22 163.367
R943 B.n1017 B.n24 163.367
R944 B.n1013 B.n24 163.367
R945 B.n1013 B.n30 163.367
R946 B.n1009 B.n30 163.367
R947 B.n1009 B.n32 163.367
R948 B.n1005 B.n32 163.367
R949 B.n1005 B.n37 163.367
R950 B.n1001 B.n37 163.367
R951 B.n1001 B.n39 163.367
R952 B.n997 B.n39 163.367
R953 B.n997 B.n44 163.367
R954 B.n993 B.n44 163.367
R955 B.n993 B.n46 163.367
R956 B.n989 B.n46 163.367
R957 B.n989 B.n51 163.367
R958 B.n985 B.n51 163.367
R959 B.n985 B.n53 163.367
R960 B.n981 B.n53 163.367
R961 B.n981 B.n58 163.367
R962 B.n977 B.n58 163.367
R963 B.n977 B.n60 163.367
R964 B.n973 B.n60 163.367
R965 B.n973 B.n65 163.367
R966 B.n969 B.n65 163.367
R967 B.n969 B.n67 163.367
R968 B.n965 B.n67 163.367
R969 B.n965 B.n71 163.367
R970 B.n961 B.n71 163.367
R971 B.n961 B.n73 163.367
R972 B.n957 B.n73 163.367
R973 B.n957 B.n79 163.367
R974 B.n953 B.n79 163.367
R975 B.n953 B.n81 163.367
R976 B.n519 B.n518 163.367
R977 B.n744 B.n518 163.367
R978 B.n742 B.n741 163.367
R979 B.n738 B.n737 163.367
R980 B.n734 B.n733 163.367
R981 B.n730 B.n729 163.367
R982 B.n726 B.n725 163.367
R983 B.n722 B.n721 163.367
R984 B.n718 B.n717 163.367
R985 B.n714 B.n713 163.367
R986 B.n710 B.n709 163.367
R987 B.n706 B.n705 163.367
R988 B.n702 B.n701 163.367
R989 B.n698 B.n697 163.367
R990 B.n694 B.n693 163.367
R991 B.n690 B.n689 163.367
R992 B.n686 B.n685 163.367
R993 B.n682 B.n681 163.367
R994 B.n678 B.n677 163.367
R995 B.n674 B.n673 163.367
R996 B.n670 B.n669 163.367
R997 B.n666 B.n665 163.367
R998 B.n662 B.n661 163.367
R999 B.n658 B.n657 163.367
R1000 B.n654 B.n653 163.367
R1001 B.n650 B.n649 163.367
R1002 B.n646 B.n645 163.367
R1003 B.n642 B.n641 163.367
R1004 B.n638 B.n637 163.367
R1005 B.n634 B.n633 163.367
R1006 B.n630 B.n629 163.367
R1007 B.n625 B.n624 163.367
R1008 B.n621 B.n620 163.367
R1009 B.n617 B.n616 163.367
R1010 B.n613 B.n612 163.367
R1011 B.n609 B.n608 163.367
R1012 B.n605 B.n604 163.367
R1013 B.n601 B.n600 163.367
R1014 B.n597 B.n596 163.367
R1015 B.n593 B.n592 163.367
R1016 B.n589 B.n588 163.367
R1017 B.n585 B.n584 163.367
R1018 B.n581 B.n580 163.367
R1019 B.n577 B.n576 163.367
R1020 B.n573 B.n572 163.367
R1021 B.n569 B.n568 163.367
R1022 B.n565 B.n564 163.367
R1023 B.n561 B.n560 163.367
R1024 B.n557 B.n556 163.367
R1025 B.n553 B.n552 163.367
R1026 B.n549 B.n548 163.367
R1027 B.n545 B.n544 163.367
R1028 B.n541 B.n540 163.367
R1029 B.n537 B.n536 163.367
R1030 B.n533 B.n532 163.367
R1031 B.n529 B.n528 163.367
R1032 B.n525 B.n462 163.367
R1033 B.n757 B.n460 163.367
R1034 B.n757 B.n454 163.367
R1035 B.n765 B.n454 163.367
R1036 B.n765 B.n452 163.367
R1037 B.n769 B.n452 163.367
R1038 B.n769 B.n447 163.367
R1039 B.n778 B.n447 163.367
R1040 B.n778 B.n445 163.367
R1041 B.n782 B.n445 163.367
R1042 B.n782 B.n439 163.367
R1043 B.n790 B.n439 163.367
R1044 B.n790 B.n437 163.367
R1045 B.n794 B.n437 163.367
R1046 B.n794 B.n431 163.367
R1047 B.n802 B.n431 163.367
R1048 B.n802 B.n429 163.367
R1049 B.n806 B.n429 163.367
R1050 B.n806 B.n423 163.367
R1051 B.n814 B.n423 163.367
R1052 B.n814 B.n421 163.367
R1053 B.n818 B.n421 163.367
R1054 B.n818 B.n415 163.367
R1055 B.n826 B.n415 163.367
R1056 B.n826 B.n413 163.367
R1057 B.n830 B.n413 163.367
R1058 B.n830 B.n406 163.367
R1059 B.n838 B.n406 163.367
R1060 B.n838 B.n404 163.367
R1061 B.n842 B.n404 163.367
R1062 B.n842 B.n399 163.367
R1063 B.n850 B.n399 163.367
R1064 B.n850 B.n397 163.367
R1065 B.n854 B.n397 163.367
R1066 B.n854 B.n392 163.367
R1067 B.n863 B.n392 163.367
R1068 B.n863 B.n390 163.367
R1069 B.n867 B.n390 163.367
R1070 B.n867 B.n383 163.367
R1071 B.n875 B.n383 163.367
R1072 B.n875 B.n381 163.367
R1073 B.n880 B.n381 163.367
R1074 B.n880 B.n376 163.367
R1075 B.n888 B.n376 163.367
R1076 B.n889 B.n888 163.367
R1077 B.n889 B.n5 163.367
R1078 B.n6 B.n5 163.367
R1079 B.n7 B.n6 163.367
R1080 B.n894 B.n7 163.367
R1081 B.n894 B.n12 163.367
R1082 B.n13 B.n12 163.367
R1083 B.n14 B.n13 163.367
R1084 B.n899 B.n14 163.367
R1085 B.n899 B.n19 163.367
R1086 B.n20 B.n19 163.367
R1087 B.n21 B.n20 163.367
R1088 B.n904 B.n21 163.367
R1089 B.n904 B.n26 163.367
R1090 B.n27 B.n26 163.367
R1091 B.n28 B.n27 163.367
R1092 B.n909 B.n28 163.367
R1093 B.n909 B.n33 163.367
R1094 B.n34 B.n33 163.367
R1095 B.n35 B.n34 163.367
R1096 B.n914 B.n35 163.367
R1097 B.n914 B.n40 163.367
R1098 B.n41 B.n40 163.367
R1099 B.n42 B.n41 163.367
R1100 B.n919 B.n42 163.367
R1101 B.n919 B.n47 163.367
R1102 B.n48 B.n47 163.367
R1103 B.n49 B.n48 163.367
R1104 B.n924 B.n49 163.367
R1105 B.n924 B.n54 163.367
R1106 B.n55 B.n54 163.367
R1107 B.n56 B.n55 163.367
R1108 B.n929 B.n56 163.367
R1109 B.n929 B.n61 163.367
R1110 B.n62 B.n61 163.367
R1111 B.n63 B.n62 163.367
R1112 B.n934 B.n63 163.367
R1113 B.n934 B.n68 163.367
R1114 B.n69 B.n68 163.367
R1115 B.n70 B.n69 163.367
R1116 B.n939 B.n70 163.367
R1117 B.n939 B.n75 163.367
R1118 B.n76 B.n75 163.367
R1119 B.n77 B.n76 163.367
R1120 B.n944 B.n77 163.367
R1121 B.n944 B.n82 163.367
R1122 B.n83 B.n82 163.367
R1123 B.n151 B.n150 163.367
R1124 B.n155 B.n154 163.367
R1125 B.n159 B.n158 163.367
R1126 B.n163 B.n162 163.367
R1127 B.n167 B.n166 163.367
R1128 B.n171 B.n170 163.367
R1129 B.n175 B.n174 163.367
R1130 B.n179 B.n178 163.367
R1131 B.n183 B.n182 163.367
R1132 B.n187 B.n186 163.367
R1133 B.n191 B.n190 163.367
R1134 B.n195 B.n194 163.367
R1135 B.n199 B.n198 163.367
R1136 B.n203 B.n202 163.367
R1137 B.n207 B.n206 163.367
R1138 B.n211 B.n210 163.367
R1139 B.n215 B.n214 163.367
R1140 B.n219 B.n218 163.367
R1141 B.n223 B.n222 163.367
R1142 B.n227 B.n226 163.367
R1143 B.n231 B.n230 163.367
R1144 B.n235 B.n234 163.367
R1145 B.n239 B.n238 163.367
R1146 B.n243 B.n242 163.367
R1147 B.n247 B.n246 163.367
R1148 B.n251 B.n250 163.367
R1149 B.n256 B.n255 163.367
R1150 B.n260 B.n259 163.367
R1151 B.n264 B.n263 163.367
R1152 B.n268 B.n267 163.367
R1153 B.n272 B.n271 163.367
R1154 B.n276 B.n275 163.367
R1155 B.n280 B.n279 163.367
R1156 B.n284 B.n283 163.367
R1157 B.n288 B.n287 163.367
R1158 B.n292 B.n291 163.367
R1159 B.n296 B.n295 163.367
R1160 B.n300 B.n299 163.367
R1161 B.n304 B.n303 163.367
R1162 B.n308 B.n307 163.367
R1163 B.n312 B.n311 163.367
R1164 B.n316 B.n315 163.367
R1165 B.n320 B.n319 163.367
R1166 B.n324 B.n323 163.367
R1167 B.n328 B.n327 163.367
R1168 B.n332 B.n331 163.367
R1169 B.n336 B.n335 163.367
R1170 B.n340 B.n339 163.367
R1171 B.n344 B.n343 163.367
R1172 B.n348 B.n347 163.367
R1173 B.n352 B.n351 163.367
R1174 B.n356 B.n355 163.367
R1175 B.n360 B.n359 163.367
R1176 B.n364 B.n363 163.367
R1177 B.n368 B.n367 163.367
R1178 B.n372 B.n371 163.367
R1179 B.n949 B.n141 163.367
R1180 B.n523 B.t15 110.07
R1181 B.n142 B.t7 110.07
R1182 B.n520 B.t12 110.049
R1183 B.n145 B.t17 110.049
R1184 B.n750 B.n749 71.676
R1185 B.n744 B.n463 71.676
R1186 B.n741 B.n464 71.676
R1187 B.n737 B.n465 71.676
R1188 B.n733 B.n466 71.676
R1189 B.n729 B.n467 71.676
R1190 B.n725 B.n468 71.676
R1191 B.n721 B.n469 71.676
R1192 B.n717 B.n470 71.676
R1193 B.n713 B.n471 71.676
R1194 B.n709 B.n472 71.676
R1195 B.n705 B.n473 71.676
R1196 B.n701 B.n474 71.676
R1197 B.n697 B.n475 71.676
R1198 B.n693 B.n476 71.676
R1199 B.n689 B.n477 71.676
R1200 B.n685 B.n478 71.676
R1201 B.n681 B.n479 71.676
R1202 B.n677 B.n480 71.676
R1203 B.n673 B.n481 71.676
R1204 B.n669 B.n482 71.676
R1205 B.n665 B.n483 71.676
R1206 B.n661 B.n484 71.676
R1207 B.n657 B.n485 71.676
R1208 B.n653 B.n486 71.676
R1209 B.n649 B.n487 71.676
R1210 B.n645 B.n488 71.676
R1211 B.n641 B.n489 71.676
R1212 B.n637 B.n490 71.676
R1213 B.n633 B.n491 71.676
R1214 B.n629 B.n492 71.676
R1215 B.n624 B.n493 71.676
R1216 B.n620 B.n494 71.676
R1217 B.n616 B.n495 71.676
R1218 B.n612 B.n496 71.676
R1219 B.n608 B.n497 71.676
R1220 B.n604 B.n498 71.676
R1221 B.n600 B.n499 71.676
R1222 B.n596 B.n500 71.676
R1223 B.n592 B.n501 71.676
R1224 B.n588 B.n502 71.676
R1225 B.n584 B.n503 71.676
R1226 B.n580 B.n504 71.676
R1227 B.n576 B.n505 71.676
R1228 B.n572 B.n506 71.676
R1229 B.n568 B.n507 71.676
R1230 B.n564 B.n508 71.676
R1231 B.n560 B.n509 71.676
R1232 B.n556 B.n510 71.676
R1233 B.n552 B.n511 71.676
R1234 B.n548 B.n512 71.676
R1235 B.n544 B.n513 71.676
R1236 B.n540 B.n514 71.676
R1237 B.n536 B.n515 71.676
R1238 B.n532 B.n516 71.676
R1239 B.n528 B.n517 71.676
R1240 B.n752 B.n462 71.676
R1241 B.n147 B.n84 71.676
R1242 B.n151 B.n85 71.676
R1243 B.n155 B.n86 71.676
R1244 B.n159 B.n87 71.676
R1245 B.n163 B.n88 71.676
R1246 B.n167 B.n89 71.676
R1247 B.n171 B.n90 71.676
R1248 B.n175 B.n91 71.676
R1249 B.n179 B.n92 71.676
R1250 B.n183 B.n93 71.676
R1251 B.n187 B.n94 71.676
R1252 B.n191 B.n95 71.676
R1253 B.n195 B.n96 71.676
R1254 B.n199 B.n97 71.676
R1255 B.n203 B.n98 71.676
R1256 B.n207 B.n99 71.676
R1257 B.n211 B.n100 71.676
R1258 B.n215 B.n101 71.676
R1259 B.n219 B.n102 71.676
R1260 B.n223 B.n103 71.676
R1261 B.n227 B.n104 71.676
R1262 B.n231 B.n105 71.676
R1263 B.n235 B.n106 71.676
R1264 B.n239 B.n107 71.676
R1265 B.n243 B.n108 71.676
R1266 B.n247 B.n109 71.676
R1267 B.n251 B.n110 71.676
R1268 B.n256 B.n111 71.676
R1269 B.n260 B.n112 71.676
R1270 B.n264 B.n113 71.676
R1271 B.n268 B.n114 71.676
R1272 B.n272 B.n115 71.676
R1273 B.n276 B.n116 71.676
R1274 B.n280 B.n117 71.676
R1275 B.n284 B.n118 71.676
R1276 B.n288 B.n119 71.676
R1277 B.n292 B.n120 71.676
R1278 B.n296 B.n121 71.676
R1279 B.n300 B.n122 71.676
R1280 B.n304 B.n123 71.676
R1281 B.n308 B.n124 71.676
R1282 B.n312 B.n125 71.676
R1283 B.n316 B.n126 71.676
R1284 B.n320 B.n127 71.676
R1285 B.n324 B.n128 71.676
R1286 B.n328 B.n129 71.676
R1287 B.n332 B.n130 71.676
R1288 B.n336 B.n131 71.676
R1289 B.n340 B.n132 71.676
R1290 B.n344 B.n133 71.676
R1291 B.n348 B.n134 71.676
R1292 B.n352 B.n135 71.676
R1293 B.n356 B.n136 71.676
R1294 B.n360 B.n137 71.676
R1295 B.n364 B.n138 71.676
R1296 B.n368 B.n139 71.676
R1297 B.n372 B.n140 71.676
R1298 B.n141 B.n140 71.676
R1299 B.n371 B.n139 71.676
R1300 B.n367 B.n138 71.676
R1301 B.n363 B.n137 71.676
R1302 B.n359 B.n136 71.676
R1303 B.n355 B.n135 71.676
R1304 B.n351 B.n134 71.676
R1305 B.n347 B.n133 71.676
R1306 B.n343 B.n132 71.676
R1307 B.n339 B.n131 71.676
R1308 B.n335 B.n130 71.676
R1309 B.n331 B.n129 71.676
R1310 B.n327 B.n128 71.676
R1311 B.n323 B.n127 71.676
R1312 B.n319 B.n126 71.676
R1313 B.n315 B.n125 71.676
R1314 B.n311 B.n124 71.676
R1315 B.n307 B.n123 71.676
R1316 B.n303 B.n122 71.676
R1317 B.n299 B.n121 71.676
R1318 B.n295 B.n120 71.676
R1319 B.n291 B.n119 71.676
R1320 B.n287 B.n118 71.676
R1321 B.n283 B.n117 71.676
R1322 B.n279 B.n116 71.676
R1323 B.n275 B.n115 71.676
R1324 B.n271 B.n114 71.676
R1325 B.n267 B.n113 71.676
R1326 B.n263 B.n112 71.676
R1327 B.n259 B.n111 71.676
R1328 B.n255 B.n110 71.676
R1329 B.n250 B.n109 71.676
R1330 B.n246 B.n108 71.676
R1331 B.n242 B.n107 71.676
R1332 B.n238 B.n106 71.676
R1333 B.n234 B.n105 71.676
R1334 B.n230 B.n104 71.676
R1335 B.n226 B.n103 71.676
R1336 B.n222 B.n102 71.676
R1337 B.n218 B.n101 71.676
R1338 B.n214 B.n100 71.676
R1339 B.n210 B.n99 71.676
R1340 B.n206 B.n98 71.676
R1341 B.n202 B.n97 71.676
R1342 B.n198 B.n96 71.676
R1343 B.n194 B.n95 71.676
R1344 B.n190 B.n94 71.676
R1345 B.n186 B.n93 71.676
R1346 B.n182 B.n92 71.676
R1347 B.n178 B.n91 71.676
R1348 B.n174 B.n90 71.676
R1349 B.n170 B.n89 71.676
R1350 B.n166 B.n88 71.676
R1351 B.n162 B.n87 71.676
R1352 B.n158 B.n86 71.676
R1353 B.n154 B.n85 71.676
R1354 B.n150 B.n84 71.676
R1355 B.n750 B.n519 71.676
R1356 B.n742 B.n463 71.676
R1357 B.n738 B.n464 71.676
R1358 B.n734 B.n465 71.676
R1359 B.n730 B.n466 71.676
R1360 B.n726 B.n467 71.676
R1361 B.n722 B.n468 71.676
R1362 B.n718 B.n469 71.676
R1363 B.n714 B.n470 71.676
R1364 B.n710 B.n471 71.676
R1365 B.n706 B.n472 71.676
R1366 B.n702 B.n473 71.676
R1367 B.n698 B.n474 71.676
R1368 B.n694 B.n475 71.676
R1369 B.n690 B.n476 71.676
R1370 B.n686 B.n477 71.676
R1371 B.n682 B.n478 71.676
R1372 B.n678 B.n479 71.676
R1373 B.n674 B.n480 71.676
R1374 B.n670 B.n481 71.676
R1375 B.n666 B.n482 71.676
R1376 B.n662 B.n483 71.676
R1377 B.n658 B.n484 71.676
R1378 B.n654 B.n485 71.676
R1379 B.n650 B.n486 71.676
R1380 B.n646 B.n487 71.676
R1381 B.n642 B.n488 71.676
R1382 B.n638 B.n489 71.676
R1383 B.n634 B.n490 71.676
R1384 B.n630 B.n491 71.676
R1385 B.n625 B.n492 71.676
R1386 B.n621 B.n493 71.676
R1387 B.n617 B.n494 71.676
R1388 B.n613 B.n495 71.676
R1389 B.n609 B.n496 71.676
R1390 B.n605 B.n497 71.676
R1391 B.n601 B.n498 71.676
R1392 B.n597 B.n499 71.676
R1393 B.n593 B.n500 71.676
R1394 B.n589 B.n501 71.676
R1395 B.n585 B.n502 71.676
R1396 B.n581 B.n503 71.676
R1397 B.n577 B.n504 71.676
R1398 B.n573 B.n505 71.676
R1399 B.n569 B.n506 71.676
R1400 B.n565 B.n507 71.676
R1401 B.n561 B.n508 71.676
R1402 B.n557 B.n509 71.676
R1403 B.n553 B.n510 71.676
R1404 B.n549 B.n511 71.676
R1405 B.n545 B.n512 71.676
R1406 B.n541 B.n513 71.676
R1407 B.n537 B.n514 71.676
R1408 B.n533 B.n515 71.676
R1409 B.n529 B.n516 71.676
R1410 B.n525 B.n517 71.676
R1411 B.n753 B.n752 71.676
R1412 B.n524 B.t14 69.5367
R1413 B.n143 B.t8 69.5367
R1414 B.n521 B.t11 69.5159
R1415 B.n146 B.t18 69.5159
R1416 B.n751 B.n459 64.3831
R1417 B.n951 B.n950 64.3831
R1418 B.n627 B.n524 59.5399
R1419 B.n522 B.n521 59.5399
R1420 B.n253 B.n146 59.5399
R1421 B.n144 B.n143 59.5399
R1422 B.n524 B.n523 40.5338
R1423 B.n521 B.n520 40.5338
R1424 B.n146 B.n145 40.5338
R1425 B.n143 B.n142 40.5338
R1426 B.n758 B.n459 35.5941
R1427 B.n758 B.n455 35.5941
R1428 B.n764 B.n455 35.5941
R1429 B.n764 B.n451 35.5941
R1430 B.n771 B.n451 35.5941
R1431 B.n771 B.n770 35.5941
R1432 B.n777 B.n444 35.5941
R1433 B.n783 B.n444 35.5941
R1434 B.n783 B.n440 35.5941
R1435 B.n789 B.n440 35.5941
R1436 B.n789 B.n436 35.5941
R1437 B.n795 B.n436 35.5941
R1438 B.n795 B.n432 35.5941
R1439 B.n801 B.n432 35.5941
R1440 B.n807 B.n428 35.5941
R1441 B.n807 B.n424 35.5941
R1442 B.n813 B.n424 35.5941
R1443 B.n813 B.n420 35.5941
R1444 B.n819 B.n420 35.5941
R1445 B.n825 B.n416 35.5941
R1446 B.n825 B.n412 35.5941
R1447 B.n831 B.n412 35.5941
R1448 B.n831 B.n407 35.5941
R1449 B.n837 B.n407 35.5941
R1450 B.n837 B.n408 35.5941
R1451 B.n843 B.n400 35.5941
R1452 B.n849 B.n400 35.5941
R1453 B.n849 B.n396 35.5941
R1454 B.n856 B.n396 35.5941
R1455 B.n856 B.n855 35.5941
R1456 B.n862 B.n389 35.5941
R1457 B.n868 B.n389 35.5941
R1458 B.n868 B.n384 35.5941
R1459 B.n874 B.n384 35.5941
R1460 B.n874 B.n385 35.5941
R1461 B.n881 B.n377 35.5941
R1462 B.n887 B.n377 35.5941
R1463 B.n887 B.n4 35.5941
R1464 B.n1040 B.n4 35.5941
R1465 B.n1040 B.n1039 35.5941
R1466 B.n1039 B.n1038 35.5941
R1467 B.n1038 B.n8 35.5941
R1468 B.n1032 B.n8 35.5941
R1469 B.n1031 B.n1030 35.5941
R1470 B.n1030 B.n15 35.5941
R1471 B.n1024 B.n15 35.5941
R1472 B.n1024 B.n1023 35.5941
R1473 B.n1023 B.n1022 35.5941
R1474 B.n1016 B.n25 35.5941
R1475 B.n1016 B.n1015 35.5941
R1476 B.n1015 B.n1014 35.5941
R1477 B.n1014 B.n29 35.5941
R1478 B.n1008 B.n29 35.5941
R1479 B.n1007 B.n1006 35.5941
R1480 B.n1006 B.n36 35.5941
R1481 B.n1000 B.n36 35.5941
R1482 B.n1000 B.n999 35.5941
R1483 B.n999 B.n998 35.5941
R1484 B.n998 B.n43 35.5941
R1485 B.n992 B.n991 35.5941
R1486 B.n991 B.n990 35.5941
R1487 B.n990 B.n50 35.5941
R1488 B.n984 B.n50 35.5941
R1489 B.n984 B.n983 35.5941
R1490 B.n982 B.n57 35.5941
R1491 B.n976 B.n57 35.5941
R1492 B.n976 B.n975 35.5941
R1493 B.n975 B.n974 35.5941
R1494 B.n974 B.n64 35.5941
R1495 B.n968 B.n64 35.5941
R1496 B.n968 B.n967 35.5941
R1497 B.n967 B.n966 35.5941
R1498 B.n960 B.n74 35.5941
R1499 B.n960 B.n959 35.5941
R1500 B.n959 B.n958 35.5941
R1501 B.n958 B.n78 35.5941
R1502 B.n952 B.n78 35.5941
R1503 B.n952 B.n951 35.5941
R1504 B.n843 B.t3 34.5473
R1505 B.n1008 B.t1 34.5473
R1506 B.n819 B.t0 31.4066
R1507 B.n992 B.t4 31.4066
R1508 B.n148 B.n80 31.3761
R1509 B.n948 B.n947 31.3761
R1510 B.n755 B.n754 31.3761
R1511 B.n748 B.n457 31.3761
R1512 B.n862 B.t2 29.3129
R1513 B.n1022 B.t19 29.3129
R1514 B.n801 B.t20 26.1723
R1515 B.t22 B.n982 26.1723
R1516 B.n881 B.t23 24.0785
R1517 B.n1032 B.t21 24.0785
R1518 B.n777 B.t10 21.9848
R1519 B.n966 B.t6 21.9848
R1520 B B.n1042 18.0485
R1521 B.n770 B.t10 13.6098
R1522 B.n74 B.t6 13.6098
R1523 B.n385 B.t23 11.5161
R1524 B.t21 B.n1031 11.5161
R1525 B.n149 B.n148 10.6151
R1526 B.n152 B.n149 10.6151
R1527 B.n153 B.n152 10.6151
R1528 B.n156 B.n153 10.6151
R1529 B.n157 B.n156 10.6151
R1530 B.n160 B.n157 10.6151
R1531 B.n161 B.n160 10.6151
R1532 B.n164 B.n161 10.6151
R1533 B.n165 B.n164 10.6151
R1534 B.n168 B.n165 10.6151
R1535 B.n169 B.n168 10.6151
R1536 B.n172 B.n169 10.6151
R1537 B.n173 B.n172 10.6151
R1538 B.n176 B.n173 10.6151
R1539 B.n177 B.n176 10.6151
R1540 B.n180 B.n177 10.6151
R1541 B.n181 B.n180 10.6151
R1542 B.n184 B.n181 10.6151
R1543 B.n185 B.n184 10.6151
R1544 B.n188 B.n185 10.6151
R1545 B.n189 B.n188 10.6151
R1546 B.n192 B.n189 10.6151
R1547 B.n193 B.n192 10.6151
R1548 B.n196 B.n193 10.6151
R1549 B.n197 B.n196 10.6151
R1550 B.n200 B.n197 10.6151
R1551 B.n201 B.n200 10.6151
R1552 B.n204 B.n201 10.6151
R1553 B.n205 B.n204 10.6151
R1554 B.n208 B.n205 10.6151
R1555 B.n209 B.n208 10.6151
R1556 B.n212 B.n209 10.6151
R1557 B.n213 B.n212 10.6151
R1558 B.n216 B.n213 10.6151
R1559 B.n217 B.n216 10.6151
R1560 B.n220 B.n217 10.6151
R1561 B.n221 B.n220 10.6151
R1562 B.n224 B.n221 10.6151
R1563 B.n225 B.n224 10.6151
R1564 B.n228 B.n225 10.6151
R1565 B.n229 B.n228 10.6151
R1566 B.n232 B.n229 10.6151
R1567 B.n233 B.n232 10.6151
R1568 B.n236 B.n233 10.6151
R1569 B.n237 B.n236 10.6151
R1570 B.n240 B.n237 10.6151
R1571 B.n241 B.n240 10.6151
R1572 B.n244 B.n241 10.6151
R1573 B.n245 B.n244 10.6151
R1574 B.n248 B.n245 10.6151
R1575 B.n249 B.n248 10.6151
R1576 B.n252 B.n249 10.6151
R1577 B.n257 B.n254 10.6151
R1578 B.n258 B.n257 10.6151
R1579 B.n261 B.n258 10.6151
R1580 B.n262 B.n261 10.6151
R1581 B.n265 B.n262 10.6151
R1582 B.n266 B.n265 10.6151
R1583 B.n269 B.n266 10.6151
R1584 B.n270 B.n269 10.6151
R1585 B.n274 B.n273 10.6151
R1586 B.n277 B.n274 10.6151
R1587 B.n278 B.n277 10.6151
R1588 B.n281 B.n278 10.6151
R1589 B.n282 B.n281 10.6151
R1590 B.n285 B.n282 10.6151
R1591 B.n286 B.n285 10.6151
R1592 B.n289 B.n286 10.6151
R1593 B.n290 B.n289 10.6151
R1594 B.n293 B.n290 10.6151
R1595 B.n294 B.n293 10.6151
R1596 B.n297 B.n294 10.6151
R1597 B.n298 B.n297 10.6151
R1598 B.n301 B.n298 10.6151
R1599 B.n302 B.n301 10.6151
R1600 B.n305 B.n302 10.6151
R1601 B.n306 B.n305 10.6151
R1602 B.n309 B.n306 10.6151
R1603 B.n310 B.n309 10.6151
R1604 B.n313 B.n310 10.6151
R1605 B.n314 B.n313 10.6151
R1606 B.n317 B.n314 10.6151
R1607 B.n318 B.n317 10.6151
R1608 B.n321 B.n318 10.6151
R1609 B.n322 B.n321 10.6151
R1610 B.n325 B.n322 10.6151
R1611 B.n326 B.n325 10.6151
R1612 B.n329 B.n326 10.6151
R1613 B.n330 B.n329 10.6151
R1614 B.n333 B.n330 10.6151
R1615 B.n334 B.n333 10.6151
R1616 B.n337 B.n334 10.6151
R1617 B.n338 B.n337 10.6151
R1618 B.n341 B.n338 10.6151
R1619 B.n342 B.n341 10.6151
R1620 B.n345 B.n342 10.6151
R1621 B.n346 B.n345 10.6151
R1622 B.n349 B.n346 10.6151
R1623 B.n350 B.n349 10.6151
R1624 B.n353 B.n350 10.6151
R1625 B.n354 B.n353 10.6151
R1626 B.n357 B.n354 10.6151
R1627 B.n358 B.n357 10.6151
R1628 B.n361 B.n358 10.6151
R1629 B.n362 B.n361 10.6151
R1630 B.n365 B.n362 10.6151
R1631 B.n366 B.n365 10.6151
R1632 B.n369 B.n366 10.6151
R1633 B.n370 B.n369 10.6151
R1634 B.n373 B.n370 10.6151
R1635 B.n374 B.n373 10.6151
R1636 B.n948 B.n374 10.6151
R1637 B.n756 B.n755 10.6151
R1638 B.n756 B.n453 10.6151
R1639 B.n766 B.n453 10.6151
R1640 B.n767 B.n766 10.6151
R1641 B.n768 B.n767 10.6151
R1642 B.n768 B.n446 10.6151
R1643 B.n779 B.n446 10.6151
R1644 B.n780 B.n779 10.6151
R1645 B.n781 B.n780 10.6151
R1646 B.n781 B.n438 10.6151
R1647 B.n791 B.n438 10.6151
R1648 B.n792 B.n791 10.6151
R1649 B.n793 B.n792 10.6151
R1650 B.n793 B.n430 10.6151
R1651 B.n803 B.n430 10.6151
R1652 B.n804 B.n803 10.6151
R1653 B.n805 B.n804 10.6151
R1654 B.n805 B.n422 10.6151
R1655 B.n815 B.n422 10.6151
R1656 B.n816 B.n815 10.6151
R1657 B.n817 B.n816 10.6151
R1658 B.n817 B.n414 10.6151
R1659 B.n827 B.n414 10.6151
R1660 B.n828 B.n827 10.6151
R1661 B.n829 B.n828 10.6151
R1662 B.n829 B.n405 10.6151
R1663 B.n839 B.n405 10.6151
R1664 B.n840 B.n839 10.6151
R1665 B.n841 B.n840 10.6151
R1666 B.n841 B.n398 10.6151
R1667 B.n851 B.n398 10.6151
R1668 B.n852 B.n851 10.6151
R1669 B.n853 B.n852 10.6151
R1670 B.n853 B.n391 10.6151
R1671 B.n864 B.n391 10.6151
R1672 B.n865 B.n864 10.6151
R1673 B.n866 B.n865 10.6151
R1674 B.n866 B.n382 10.6151
R1675 B.n876 B.n382 10.6151
R1676 B.n877 B.n876 10.6151
R1677 B.n879 B.n877 10.6151
R1678 B.n879 B.n878 10.6151
R1679 B.n878 B.n375 10.6151
R1680 B.n890 B.n375 10.6151
R1681 B.n891 B.n890 10.6151
R1682 B.n892 B.n891 10.6151
R1683 B.n893 B.n892 10.6151
R1684 B.n895 B.n893 10.6151
R1685 B.n896 B.n895 10.6151
R1686 B.n897 B.n896 10.6151
R1687 B.n898 B.n897 10.6151
R1688 B.n900 B.n898 10.6151
R1689 B.n901 B.n900 10.6151
R1690 B.n902 B.n901 10.6151
R1691 B.n903 B.n902 10.6151
R1692 B.n905 B.n903 10.6151
R1693 B.n906 B.n905 10.6151
R1694 B.n907 B.n906 10.6151
R1695 B.n908 B.n907 10.6151
R1696 B.n910 B.n908 10.6151
R1697 B.n911 B.n910 10.6151
R1698 B.n912 B.n911 10.6151
R1699 B.n913 B.n912 10.6151
R1700 B.n915 B.n913 10.6151
R1701 B.n916 B.n915 10.6151
R1702 B.n917 B.n916 10.6151
R1703 B.n918 B.n917 10.6151
R1704 B.n920 B.n918 10.6151
R1705 B.n921 B.n920 10.6151
R1706 B.n922 B.n921 10.6151
R1707 B.n923 B.n922 10.6151
R1708 B.n925 B.n923 10.6151
R1709 B.n926 B.n925 10.6151
R1710 B.n927 B.n926 10.6151
R1711 B.n928 B.n927 10.6151
R1712 B.n930 B.n928 10.6151
R1713 B.n931 B.n930 10.6151
R1714 B.n932 B.n931 10.6151
R1715 B.n933 B.n932 10.6151
R1716 B.n935 B.n933 10.6151
R1717 B.n936 B.n935 10.6151
R1718 B.n937 B.n936 10.6151
R1719 B.n938 B.n937 10.6151
R1720 B.n940 B.n938 10.6151
R1721 B.n941 B.n940 10.6151
R1722 B.n942 B.n941 10.6151
R1723 B.n943 B.n942 10.6151
R1724 B.n945 B.n943 10.6151
R1725 B.n946 B.n945 10.6151
R1726 B.n947 B.n946 10.6151
R1727 B.n748 B.n747 10.6151
R1728 B.n747 B.n746 10.6151
R1729 B.n746 B.n745 10.6151
R1730 B.n745 B.n743 10.6151
R1731 B.n743 B.n740 10.6151
R1732 B.n740 B.n739 10.6151
R1733 B.n739 B.n736 10.6151
R1734 B.n736 B.n735 10.6151
R1735 B.n735 B.n732 10.6151
R1736 B.n732 B.n731 10.6151
R1737 B.n731 B.n728 10.6151
R1738 B.n728 B.n727 10.6151
R1739 B.n727 B.n724 10.6151
R1740 B.n724 B.n723 10.6151
R1741 B.n723 B.n720 10.6151
R1742 B.n720 B.n719 10.6151
R1743 B.n719 B.n716 10.6151
R1744 B.n716 B.n715 10.6151
R1745 B.n715 B.n712 10.6151
R1746 B.n712 B.n711 10.6151
R1747 B.n711 B.n708 10.6151
R1748 B.n708 B.n707 10.6151
R1749 B.n707 B.n704 10.6151
R1750 B.n704 B.n703 10.6151
R1751 B.n703 B.n700 10.6151
R1752 B.n700 B.n699 10.6151
R1753 B.n699 B.n696 10.6151
R1754 B.n696 B.n695 10.6151
R1755 B.n695 B.n692 10.6151
R1756 B.n692 B.n691 10.6151
R1757 B.n691 B.n688 10.6151
R1758 B.n688 B.n687 10.6151
R1759 B.n687 B.n684 10.6151
R1760 B.n684 B.n683 10.6151
R1761 B.n683 B.n680 10.6151
R1762 B.n680 B.n679 10.6151
R1763 B.n679 B.n676 10.6151
R1764 B.n676 B.n675 10.6151
R1765 B.n675 B.n672 10.6151
R1766 B.n672 B.n671 10.6151
R1767 B.n671 B.n668 10.6151
R1768 B.n668 B.n667 10.6151
R1769 B.n667 B.n664 10.6151
R1770 B.n664 B.n663 10.6151
R1771 B.n663 B.n660 10.6151
R1772 B.n660 B.n659 10.6151
R1773 B.n659 B.n656 10.6151
R1774 B.n656 B.n655 10.6151
R1775 B.n655 B.n652 10.6151
R1776 B.n652 B.n651 10.6151
R1777 B.n651 B.n648 10.6151
R1778 B.n648 B.n647 10.6151
R1779 B.n644 B.n643 10.6151
R1780 B.n643 B.n640 10.6151
R1781 B.n640 B.n639 10.6151
R1782 B.n639 B.n636 10.6151
R1783 B.n636 B.n635 10.6151
R1784 B.n635 B.n632 10.6151
R1785 B.n632 B.n631 10.6151
R1786 B.n631 B.n628 10.6151
R1787 B.n626 B.n623 10.6151
R1788 B.n623 B.n622 10.6151
R1789 B.n622 B.n619 10.6151
R1790 B.n619 B.n618 10.6151
R1791 B.n618 B.n615 10.6151
R1792 B.n615 B.n614 10.6151
R1793 B.n614 B.n611 10.6151
R1794 B.n611 B.n610 10.6151
R1795 B.n610 B.n607 10.6151
R1796 B.n607 B.n606 10.6151
R1797 B.n606 B.n603 10.6151
R1798 B.n603 B.n602 10.6151
R1799 B.n602 B.n599 10.6151
R1800 B.n599 B.n598 10.6151
R1801 B.n598 B.n595 10.6151
R1802 B.n595 B.n594 10.6151
R1803 B.n594 B.n591 10.6151
R1804 B.n591 B.n590 10.6151
R1805 B.n590 B.n587 10.6151
R1806 B.n587 B.n586 10.6151
R1807 B.n586 B.n583 10.6151
R1808 B.n583 B.n582 10.6151
R1809 B.n582 B.n579 10.6151
R1810 B.n579 B.n578 10.6151
R1811 B.n578 B.n575 10.6151
R1812 B.n575 B.n574 10.6151
R1813 B.n574 B.n571 10.6151
R1814 B.n571 B.n570 10.6151
R1815 B.n570 B.n567 10.6151
R1816 B.n567 B.n566 10.6151
R1817 B.n566 B.n563 10.6151
R1818 B.n563 B.n562 10.6151
R1819 B.n562 B.n559 10.6151
R1820 B.n559 B.n558 10.6151
R1821 B.n558 B.n555 10.6151
R1822 B.n555 B.n554 10.6151
R1823 B.n554 B.n551 10.6151
R1824 B.n551 B.n550 10.6151
R1825 B.n550 B.n547 10.6151
R1826 B.n547 B.n546 10.6151
R1827 B.n546 B.n543 10.6151
R1828 B.n543 B.n542 10.6151
R1829 B.n542 B.n539 10.6151
R1830 B.n539 B.n538 10.6151
R1831 B.n538 B.n535 10.6151
R1832 B.n535 B.n534 10.6151
R1833 B.n534 B.n531 10.6151
R1834 B.n531 B.n530 10.6151
R1835 B.n530 B.n527 10.6151
R1836 B.n527 B.n526 10.6151
R1837 B.n526 B.n461 10.6151
R1838 B.n754 B.n461 10.6151
R1839 B.n760 B.n457 10.6151
R1840 B.n761 B.n760 10.6151
R1841 B.n762 B.n761 10.6151
R1842 B.n762 B.n449 10.6151
R1843 B.n773 B.n449 10.6151
R1844 B.n774 B.n773 10.6151
R1845 B.n775 B.n774 10.6151
R1846 B.n775 B.n442 10.6151
R1847 B.n785 B.n442 10.6151
R1848 B.n786 B.n785 10.6151
R1849 B.n787 B.n786 10.6151
R1850 B.n787 B.n434 10.6151
R1851 B.n797 B.n434 10.6151
R1852 B.n798 B.n797 10.6151
R1853 B.n799 B.n798 10.6151
R1854 B.n799 B.n426 10.6151
R1855 B.n809 B.n426 10.6151
R1856 B.n810 B.n809 10.6151
R1857 B.n811 B.n810 10.6151
R1858 B.n811 B.n418 10.6151
R1859 B.n821 B.n418 10.6151
R1860 B.n822 B.n821 10.6151
R1861 B.n823 B.n822 10.6151
R1862 B.n823 B.n410 10.6151
R1863 B.n833 B.n410 10.6151
R1864 B.n834 B.n833 10.6151
R1865 B.n835 B.n834 10.6151
R1866 B.n835 B.n402 10.6151
R1867 B.n845 B.n402 10.6151
R1868 B.n846 B.n845 10.6151
R1869 B.n847 B.n846 10.6151
R1870 B.n847 B.n394 10.6151
R1871 B.n858 B.n394 10.6151
R1872 B.n859 B.n858 10.6151
R1873 B.n860 B.n859 10.6151
R1874 B.n860 B.n387 10.6151
R1875 B.n870 B.n387 10.6151
R1876 B.n871 B.n870 10.6151
R1877 B.n872 B.n871 10.6151
R1878 B.n872 B.n379 10.6151
R1879 B.n883 B.n379 10.6151
R1880 B.n884 B.n883 10.6151
R1881 B.n885 B.n884 10.6151
R1882 B.n885 B.n0 10.6151
R1883 B.n1036 B.n1 10.6151
R1884 B.n1036 B.n1035 10.6151
R1885 B.n1035 B.n1034 10.6151
R1886 B.n1034 B.n10 10.6151
R1887 B.n1028 B.n10 10.6151
R1888 B.n1028 B.n1027 10.6151
R1889 B.n1027 B.n1026 10.6151
R1890 B.n1026 B.n17 10.6151
R1891 B.n1020 B.n17 10.6151
R1892 B.n1020 B.n1019 10.6151
R1893 B.n1019 B.n1018 10.6151
R1894 B.n1018 B.n23 10.6151
R1895 B.n1012 B.n23 10.6151
R1896 B.n1012 B.n1011 10.6151
R1897 B.n1011 B.n1010 10.6151
R1898 B.n1010 B.n31 10.6151
R1899 B.n1004 B.n31 10.6151
R1900 B.n1004 B.n1003 10.6151
R1901 B.n1003 B.n1002 10.6151
R1902 B.n1002 B.n38 10.6151
R1903 B.n996 B.n38 10.6151
R1904 B.n996 B.n995 10.6151
R1905 B.n995 B.n994 10.6151
R1906 B.n994 B.n45 10.6151
R1907 B.n988 B.n45 10.6151
R1908 B.n988 B.n987 10.6151
R1909 B.n987 B.n986 10.6151
R1910 B.n986 B.n52 10.6151
R1911 B.n980 B.n52 10.6151
R1912 B.n980 B.n979 10.6151
R1913 B.n979 B.n978 10.6151
R1914 B.n978 B.n59 10.6151
R1915 B.n972 B.n59 10.6151
R1916 B.n972 B.n971 10.6151
R1917 B.n971 B.n970 10.6151
R1918 B.n970 B.n66 10.6151
R1919 B.n964 B.n66 10.6151
R1920 B.n964 B.n963 10.6151
R1921 B.n963 B.n962 10.6151
R1922 B.n962 B.n72 10.6151
R1923 B.n956 B.n72 10.6151
R1924 B.n956 B.n955 10.6151
R1925 B.n955 B.n954 10.6151
R1926 B.n954 B.n80 10.6151
R1927 B.t20 B.n428 9.42234
R1928 B.n983 B.t22 9.42234
R1929 B.n254 B.n253 6.4005
R1930 B.n270 B.n144 6.4005
R1931 B.n644 B.n522 6.4005
R1932 B.n628 B.n627 6.4005
R1933 B.n855 B.t2 6.28173
R1934 B.n25 B.t19 6.28173
R1935 B.n253 B.n252 4.21513
R1936 B.n273 B.n144 4.21513
R1937 B.n647 B.n522 4.21513
R1938 B.n627 B.n626 4.21513
R1939 B.t0 B.n416 4.18799
R1940 B.t4 B.n43 4.18799
R1941 B.n1042 B.n0 2.81026
R1942 B.n1042 B.n1 2.81026
R1943 B.n408 B.t3 1.04737
R1944 B.t1 B.n1007 1.04737
R1945 VN.n6 VN.t1 246.417
R1946 VN.n36 VN.t7 246.417
R1947 VN.n7 VN.t6 215.531
R1948 VN.n14 VN.t5 215.531
R1949 VN.n21 VN.t0 215.531
R1950 VN.n28 VN.t9 215.531
R1951 VN.n37 VN.t4 215.531
R1952 VN.n44 VN.t2 215.531
R1953 VN.n51 VN.t3 215.531
R1954 VN.n58 VN.t8 215.531
R1955 VN.n57 VN.n30 161.3
R1956 VN.n56 VN.n55 161.3
R1957 VN.n54 VN.n31 161.3
R1958 VN.n53 VN.n52 161.3
R1959 VN.n50 VN.n32 161.3
R1960 VN.n49 VN.n48 161.3
R1961 VN.n47 VN.n33 161.3
R1962 VN.n46 VN.n45 161.3
R1963 VN.n43 VN.n34 161.3
R1964 VN.n42 VN.n41 161.3
R1965 VN.n40 VN.n35 161.3
R1966 VN.n39 VN.n38 161.3
R1967 VN.n27 VN.n0 161.3
R1968 VN.n26 VN.n25 161.3
R1969 VN.n24 VN.n1 161.3
R1970 VN.n23 VN.n22 161.3
R1971 VN.n20 VN.n2 161.3
R1972 VN.n19 VN.n18 161.3
R1973 VN.n17 VN.n3 161.3
R1974 VN.n16 VN.n15 161.3
R1975 VN.n13 VN.n4 161.3
R1976 VN.n12 VN.n11 161.3
R1977 VN.n10 VN.n5 161.3
R1978 VN.n9 VN.n8 161.3
R1979 VN.n29 VN.n28 89.6708
R1980 VN.n59 VN.n58 89.6708
R1981 VN.n12 VN.n5 56.4773
R1982 VN.n19 VN.n3 56.4773
R1983 VN.n42 VN.n35 56.4773
R1984 VN.n49 VN.n33 56.4773
R1985 VN.n7 VN.n6 52.8339
R1986 VN.n37 VN.n36 52.8339
R1987 VN VN.n59 51.6458
R1988 VN.n26 VN.n1 51.6086
R1989 VN.n56 VN.n31 51.6086
R1990 VN.n27 VN.n26 29.2126
R1991 VN.n57 VN.n56 29.2126
R1992 VN.n8 VN.n5 24.3439
R1993 VN.n13 VN.n12 24.3439
R1994 VN.n15 VN.n3 24.3439
R1995 VN.n20 VN.n19 24.3439
R1996 VN.n22 VN.n1 24.3439
R1997 VN.n38 VN.n35 24.3439
R1998 VN.n45 VN.n33 24.3439
R1999 VN.n43 VN.n42 24.3439
R2000 VN.n52 VN.n31 24.3439
R2001 VN.n50 VN.n49 24.3439
R2002 VN.n28 VN.n27 20.9359
R2003 VN.n58 VN.n57 20.9359
R2004 VN.n8 VN.n7 16.554
R2005 VN.n21 VN.n20 16.554
R2006 VN.n38 VN.n37 16.554
R2007 VN.n51 VN.n50 16.554
R2008 VN.n39 VN.n36 13.1234
R2009 VN.n9 VN.n6 13.1234
R2010 VN.n14 VN.n13 12.1722
R2011 VN.n15 VN.n14 12.1722
R2012 VN.n45 VN.n44 12.1722
R2013 VN.n44 VN.n43 12.1722
R2014 VN.n22 VN.n21 7.7904
R2015 VN.n52 VN.n51 7.7904
R2016 VN.n59 VN.n30 0.278398
R2017 VN.n29 VN.n0 0.278398
R2018 VN.n55 VN.n30 0.189894
R2019 VN.n55 VN.n54 0.189894
R2020 VN.n54 VN.n53 0.189894
R2021 VN.n53 VN.n32 0.189894
R2022 VN.n48 VN.n32 0.189894
R2023 VN.n48 VN.n47 0.189894
R2024 VN.n47 VN.n46 0.189894
R2025 VN.n46 VN.n34 0.189894
R2026 VN.n41 VN.n34 0.189894
R2027 VN.n41 VN.n40 0.189894
R2028 VN.n40 VN.n39 0.189894
R2029 VN.n10 VN.n9 0.189894
R2030 VN.n11 VN.n10 0.189894
R2031 VN.n11 VN.n4 0.189894
R2032 VN.n16 VN.n4 0.189894
R2033 VN.n17 VN.n16 0.189894
R2034 VN.n18 VN.n17 0.189894
R2035 VN.n18 VN.n2 0.189894
R2036 VN.n23 VN.n2 0.189894
R2037 VN.n24 VN.n23 0.189894
R2038 VN.n25 VN.n24 0.189894
R2039 VN.n25 VN.n0 0.189894
R2040 VN VN.n29 0.153422
R2041 VDD2.n1 VDD2.t8 64.2557
R2042 VDD2.n3 VDD2.n2 62.4919
R2043 VDD2 VDD2.n7 62.4891
R2044 VDD2.n4 VDD2.t1 62.4541
R2045 VDD2.n6 VDD2.n5 61.1962
R2046 VDD2.n1 VDD2.n0 61.1959
R2047 VDD2.n4 VDD2.n3 45.8425
R2048 VDD2.n6 VDD2.n4 1.80222
R2049 VDD2.n7 VDD2.t5 1.25844
R2050 VDD2.n7 VDD2.t2 1.25844
R2051 VDD2.n5 VDD2.t6 1.25844
R2052 VDD2.n5 VDD2.t7 1.25844
R2053 VDD2.n2 VDD2.t9 1.25844
R2054 VDD2.n2 VDD2.t0 1.25844
R2055 VDD2.n0 VDD2.t3 1.25844
R2056 VDD2.n0 VDD2.t4 1.25844
R2057 VDD2 VDD2.n6 0.509121
R2058 VDD2.n3 VDD2.n1 0.395585
C0 VDD1 VDD2 1.62902f
C1 VP VTAIL 12.7463f
C2 VN VDD2 12.5925f
C3 VDD1 VP 12.913099f
C4 VDD1 VTAIL 12.7231f
C5 VN VP 7.862871f
C6 VN VTAIL 12.7318f
C7 VDD1 VN 0.151176f
C8 VP VDD2 0.476619f
C9 VDD2 VTAIL 12.766001f
C10 VDD2 B 6.876759f
C11 VDD1 B 6.858693f
C12 VTAIL B 8.972833f
C13 VN B 14.587881f
C14 VP B 12.905174f
C15 VDD2.t8 B 3.21074f
C16 VDD2.t3 B 0.276584f
C17 VDD2.t4 B 0.276584f
C18 VDD2.n0 B 2.50585f
C19 VDD2.n1 B 0.711134f
C20 VDD2.t9 B 0.276584f
C21 VDD2.t0 B 0.276584f
C22 VDD2.n2 B 2.51443f
C23 VDD2.n3 B 2.39807f
C24 VDD2.t1 B 3.20008f
C25 VDD2.n4 B 2.74503f
C26 VDD2.t6 B 0.276584f
C27 VDD2.t7 B 0.276584f
C28 VDD2.n5 B 2.50585f
C29 VDD2.n6 B 0.348009f
C30 VDD2.t5 B 0.276584f
C31 VDD2.t2 B 0.276584f
C32 VDD2.n7 B 2.51439f
C33 VN.n0 B 0.035288f
C34 VN.t9 B 2.03296f
C35 VN.n1 B 0.048563f
C36 VN.n2 B 0.026764f
C37 VN.t0 B 2.03296f
C38 VN.n3 B 0.042621f
C39 VN.n4 B 0.026764f
C40 VN.t5 B 2.03296f
C41 VN.n5 B 0.035861f
C42 VN.t1 B 2.13798f
C43 VN.n6 B 0.787162f
C44 VN.t6 B 2.03296f
C45 VN.n7 B 0.780616f
C46 VN.n8 B 0.042211f
C47 VN.n9 B 0.194644f
C48 VN.n10 B 0.026764f
C49 VN.n11 B 0.026764f
C50 VN.n12 B 0.042621f
C51 VN.n13 B 0.037756f
C52 VN.n14 B 0.717368f
C53 VN.n15 B 0.037756f
C54 VN.n16 B 0.026764f
C55 VN.n17 B 0.026764f
C56 VN.n18 B 0.026764f
C57 VN.n19 B 0.035861f
C58 VN.n20 B 0.042211f
C59 VN.n21 B 0.717368f
C60 VN.n22 B 0.033301f
C61 VN.n23 B 0.026764f
C62 VN.n24 B 0.026764f
C63 VN.n25 B 0.026764f
C64 VN.n26 B 0.026619f
C65 VN.n27 B 0.049967f
C66 VN.n28 B 0.791985f
C67 VN.n29 B 0.030583f
C68 VN.n30 B 0.035288f
C69 VN.t8 B 2.03296f
C70 VN.n31 B 0.048563f
C71 VN.n32 B 0.026764f
C72 VN.t3 B 2.03296f
C73 VN.n33 B 0.042621f
C74 VN.n34 B 0.026764f
C75 VN.t2 B 2.03296f
C76 VN.n35 B 0.035861f
C77 VN.t7 B 2.13798f
C78 VN.n36 B 0.787162f
C79 VN.t4 B 2.03296f
C80 VN.n37 B 0.780616f
C81 VN.n38 B 0.042211f
C82 VN.n39 B 0.194644f
C83 VN.n40 B 0.026764f
C84 VN.n41 B 0.026764f
C85 VN.n42 B 0.042621f
C86 VN.n43 B 0.037756f
C87 VN.n44 B 0.717368f
C88 VN.n45 B 0.037756f
C89 VN.n46 B 0.026764f
C90 VN.n47 B 0.026764f
C91 VN.n48 B 0.026764f
C92 VN.n49 B 0.035861f
C93 VN.n50 B 0.042211f
C94 VN.n51 B 0.717368f
C95 VN.n52 B 0.033301f
C96 VN.n53 B 0.026764f
C97 VN.n54 B 0.026764f
C98 VN.n55 B 0.026764f
C99 VN.n56 B 0.026619f
C100 VN.n57 B 0.049967f
C101 VN.n58 B 0.791985f
C102 VN.n59 B 1.54892f
C103 VTAIL.t15 B 0.295325f
C104 VTAIL.t16 B 0.295325f
C105 VTAIL.n0 B 2.60434f
C106 VTAIL.n1 B 0.446569f
C107 VTAIL.t12 B 3.32417f
C108 VTAIL.n2 B 0.562176f
C109 VTAIL.t13 B 0.295325f
C110 VTAIL.t14 B 0.295325f
C111 VTAIL.n3 B 2.60434f
C112 VTAIL.n4 B 0.509555f
C113 VTAIL.t8 B 0.295325f
C114 VTAIL.t10 B 0.295325f
C115 VTAIL.n5 B 2.60434f
C116 VTAIL.n6 B 2.00804f
C117 VTAIL.t17 B 0.295325f
C118 VTAIL.t0 B 0.295325f
C119 VTAIL.n7 B 2.60434f
C120 VTAIL.n8 B 2.00803f
C121 VTAIL.t3 B 0.295325f
C122 VTAIL.t2 B 0.295325f
C123 VTAIL.n9 B 2.60434f
C124 VTAIL.n10 B 0.509552f
C125 VTAIL.t18 B 3.3242f
C126 VTAIL.n11 B 0.562154f
C127 VTAIL.t9 B 0.295325f
C128 VTAIL.t5 B 0.295325f
C129 VTAIL.n12 B 2.60434f
C130 VTAIL.n13 B 0.476575f
C131 VTAIL.t6 B 0.295325f
C132 VTAIL.t7 B 0.295325f
C133 VTAIL.n14 B 2.60434f
C134 VTAIL.n15 B 0.509552f
C135 VTAIL.t11 B 3.32417f
C136 VTAIL.n16 B 1.95579f
C137 VTAIL.t19 B 3.32417f
C138 VTAIL.n17 B 1.95579f
C139 VTAIL.t1 B 0.295325f
C140 VTAIL.t4 B 0.295325f
C141 VTAIL.n18 B 2.60434f
C142 VTAIL.n19 B 0.401721f
C143 VDD1.t9 B 3.22561f
C144 VDD1.t2 B 0.277863f
C145 VDD1.t5 B 0.277863f
C146 VDD1.n0 B 2.51744f
C147 VDD1.n1 B 0.721269f
C148 VDD1.t8 B 3.22559f
C149 VDD1.t0 B 0.277863f
C150 VDD1.t4 B 0.277863f
C151 VDD1.n2 B 2.51744f
C152 VDD1.n3 B 0.714424f
C153 VDD1.t7 B 0.277863f
C154 VDD1.t3 B 0.277863f
C155 VDD1.n4 B 2.52606f
C156 VDD1.n5 B 2.50292f
C157 VDD1.t6 B 0.277863f
C158 VDD1.t1 B 0.277863f
C159 VDD1.n6 B 2.51743f
C160 VDD1.n7 B 2.77921f
C161 VP.n0 B 0.035647f
C162 VP.t2 B 2.05366f
C163 VP.n1 B 0.049057f
C164 VP.n2 B 0.027037f
C165 VP.t0 B 2.05366f
C166 VP.n3 B 0.043055f
C167 VP.n4 B 0.027037f
C168 VP.t1 B 2.05366f
C169 VP.n5 B 0.036226f
C170 VP.n6 B 0.027037f
C171 VP.t4 B 2.05366f
C172 VP.n7 B 0.02689f
C173 VP.n8 B 0.035647f
C174 VP.t3 B 2.05366f
C175 VP.n9 B 0.049057f
C176 VP.n10 B 0.027037f
C177 VP.t7 B 2.05366f
C178 VP.n11 B 0.043055f
C179 VP.n12 B 0.027037f
C180 VP.t8 B 2.05366f
C181 VP.n13 B 0.036226f
C182 VP.t5 B 2.15974f
C183 VP.n14 B 0.795176f
C184 VP.t9 B 2.05366f
C185 VP.n15 B 0.788564f
C186 VP.n16 B 0.042641f
C187 VP.n17 B 0.196626f
C188 VP.n18 B 0.027037f
C189 VP.n19 B 0.027037f
C190 VP.n20 B 0.043055f
C191 VP.n21 B 0.03814f
C192 VP.n22 B 0.724672f
C193 VP.n23 B 0.03814f
C194 VP.n24 B 0.027037f
C195 VP.n25 B 0.027037f
C196 VP.n26 B 0.027037f
C197 VP.n27 B 0.036226f
C198 VP.n28 B 0.042641f
C199 VP.n29 B 0.724672f
C200 VP.n30 B 0.03364f
C201 VP.n31 B 0.027037f
C202 VP.n32 B 0.027037f
C203 VP.n33 B 0.027037f
C204 VP.n34 B 0.02689f
C205 VP.n35 B 0.050476f
C206 VP.n36 B 0.800048f
C207 VP.n37 B 1.55022f
C208 VP.n38 B 1.56908f
C209 VP.t6 B 2.05366f
C210 VP.n39 B 0.800048f
C211 VP.n40 B 0.050476f
C212 VP.n41 B 0.035647f
C213 VP.n42 B 0.027037f
C214 VP.n43 B 0.027037f
C215 VP.n44 B 0.049057f
C216 VP.n45 B 0.03364f
C217 VP.n46 B 0.724672f
C218 VP.n47 B 0.042641f
C219 VP.n48 B 0.027037f
C220 VP.n49 B 0.027037f
C221 VP.n50 B 0.027037f
C222 VP.n51 B 0.043055f
C223 VP.n52 B 0.03814f
C224 VP.n53 B 0.724672f
C225 VP.n54 B 0.03814f
C226 VP.n55 B 0.027037f
C227 VP.n56 B 0.027037f
C228 VP.n57 B 0.027037f
C229 VP.n58 B 0.036226f
C230 VP.n59 B 0.042641f
C231 VP.n60 B 0.724672f
C232 VP.n61 B 0.03364f
C233 VP.n62 B 0.027037f
C234 VP.n63 B 0.027037f
C235 VP.n64 B 0.027037f
C236 VP.n65 B 0.02689f
C237 VP.n66 B 0.050476f
C238 VP.n67 B 0.800048f
C239 VP.n68 B 0.030894f
.ends

