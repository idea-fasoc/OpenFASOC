* NGSPICE file created from diff_pair_sample_1110.ext - technology: sky130A

.subckt diff_pair_sample_1110 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=4.5357 ps=24.04 w=11.63 l=1.9
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=0 ps=0 w=11.63 l=1.9
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=0 ps=0 w=11.63 l=1.9
X3 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=4.5357 ps=24.04 w=11.63 l=1.9
X4 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=4.5357 ps=24.04 w=11.63 l=1.9
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=0 ps=0 w=11.63 l=1.9
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=4.5357 ps=24.04 w=11.63 l=1.9
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5357 pd=24.04 as=0 ps=0 w=11.63 l=1.9
R0 VN VN.t1 249.089
R1 VN VN.t0 206.619
R2 VTAIL.n1 VTAIL.t1 50.8153
R3 VTAIL.n3 VTAIL.t2 50.8144
R4 VTAIL.n0 VTAIL.t3 50.8144
R5 VTAIL.n2 VTAIL.t0 50.8142
R6 VTAIL.n1 VTAIL.n0 26.2376
R7 VTAIL.n3 VTAIL.n2 24.3152
R8 VTAIL.n2 VTAIL.n1 1.43153
R9 VTAIL VTAIL.n0 1.00912
R10 VTAIL VTAIL.n3 0.422914
R11 VDD2.n0 VDD2.t1 105.023
R12 VDD2.n0 VDD2.t0 67.493
R13 VDD2 VDD2.n0 0.539293
R14 B.n637 B.n636 585
R15 B.n638 B.n637 585
R16 B.n272 B.n87 585
R17 B.n271 B.n270 585
R18 B.n269 B.n268 585
R19 B.n267 B.n266 585
R20 B.n265 B.n264 585
R21 B.n263 B.n262 585
R22 B.n261 B.n260 585
R23 B.n259 B.n258 585
R24 B.n257 B.n256 585
R25 B.n255 B.n254 585
R26 B.n253 B.n252 585
R27 B.n251 B.n250 585
R28 B.n249 B.n248 585
R29 B.n247 B.n246 585
R30 B.n245 B.n244 585
R31 B.n243 B.n242 585
R32 B.n241 B.n240 585
R33 B.n239 B.n238 585
R34 B.n237 B.n236 585
R35 B.n235 B.n234 585
R36 B.n233 B.n232 585
R37 B.n231 B.n230 585
R38 B.n229 B.n228 585
R39 B.n227 B.n226 585
R40 B.n225 B.n224 585
R41 B.n223 B.n222 585
R42 B.n221 B.n220 585
R43 B.n219 B.n218 585
R44 B.n217 B.n216 585
R45 B.n215 B.n214 585
R46 B.n213 B.n212 585
R47 B.n211 B.n210 585
R48 B.n209 B.n208 585
R49 B.n207 B.n206 585
R50 B.n205 B.n204 585
R51 B.n203 B.n202 585
R52 B.n201 B.n200 585
R53 B.n199 B.n198 585
R54 B.n197 B.n196 585
R55 B.n195 B.n194 585
R56 B.n193 B.n192 585
R57 B.n191 B.n190 585
R58 B.n189 B.n188 585
R59 B.n187 B.n186 585
R60 B.n185 B.n184 585
R61 B.n183 B.n182 585
R62 B.n181 B.n180 585
R63 B.n179 B.n178 585
R64 B.n177 B.n176 585
R65 B.n174 B.n173 585
R66 B.n172 B.n171 585
R67 B.n170 B.n169 585
R68 B.n168 B.n167 585
R69 B.n166 B.n165 585
R70 B.n164 B.n163 585
R71 B.n162 B.n161 585
R72 B.n160 B.n159 585
R73 B.n158 B.n157 585
R74 B.n156 B.n155 585
R75 B.n154 B.n153 585
R76 B.n152 B.n151 585
R77 B.n150 B.n149 585
R78 B.n148 B.n147 585
R79 B.n146 B.n145 585
R80 B.n144 B.n143 585
R81 B.n142 B.n141 585
R82 B.n140 B.n139 585
R83 B.n138 B.n137 585
R84 B.n136 B.n135 585
R85 B.n134 B.n133 585
R86 B.n132 B.n131 585
R87 B.n130 B.n129 585
R88 B.n128 B.n127 585
R89 B.n126 B.n125 585
R90 B.n124 B.n123 585
R91 B.n122 B.n121 585
R92 B.n120 B.n119 585
R93 B.n118 B.n117 585
R94 B.n116 B.n115 585
R95 B.n114 B.n113 585
R96 B.n112 B.n111 585
R97 B.n110 B.n109 585
R98 B.n108 B.n107 585
R99 B.n106 B.n105 585
R100 B.n104 B.n103 585
R101 B.n102 B.n101 585
R102 B.n100 B.n99 585
R103 B.n98 B.n97 585
R104 B.n96 B.n95 585
R105 B.n94 B.n93 585
R106 B.n635 B.n41 585
R107 B.n639 B.n41 585
R108 B.n634 B.n40 585
R109 B.n640 B.n40 585
R110 B.n633 B.n632 585
R111 B.n632 B.n36 585
R112 B.n631 B.n35 585
R113 B.n646 B.n35 585
R114 B.n630 B.n34 585
R115 B.n647 B.n34 585
R116 B.n629 B.n33 585
R117 B.n648 B.n33 585
R118 B.n628 B.n627 585
R119 B.n627 B.n32 585
R120 B.n626 B.n28 585
R121 B.n654 B.n28 585
R122 B.n625 B.n27 585
R123 B.n655 B.n27 585
R124 B.n624 B.n26 585
R125 B.n656 B.n26 585
R126 B.n623 B.n622 585
R127 B.n622 B.n22 585
R128 B.n621 B.n21 585
R129 B.n662 B.n21 585
R130 B.n620 B.n20 585
R131 B.n663 B.n20 585
R132 B.n619 B.n19 585
R133 B.n664 B.n19 585
R134 B.n618 B.n617 585
R135 B.n617 B.n15 585
R136 B.n616 B.n14 585
R137 B.n670 B.n14 585
R138 B.n615 B.n13 585
R139 B.n671 B.n13 585
R140 B.n614 B.n12 585
R141 B.n672 B.n12 585
R142 B.n613 B.n612 585
R143 B.n612 B.n8 585
R144 B.n611 B.n7 585
R145 B.n678 B.n7 585
R146 B.n610 B.n6 585
R147 B.n679 B.n6 585
R148 B.n609 B.n5 585
R149 B.n680 B.n5 585
R150 B.n608 B.n607 585
R151 B.n607 B.n4 585
R152 B.n606 B.n273 585
R153 B.n606 B.n605 585
R154 B.n596 B.n274 585
R155 B.n275 B.n274 585
R156 B.n598 B.n597 585
R157 B.n599 B.n598 585
R158 B.n595 B.n279 585
R159 B.n283 B.n279 585
R160 B.n594 B.n593 585
R161 B.n593 B.n592 585
R162 B.n281 B.n280 585
R163 B.n282 B.n281 585
R164 B.n585 B.n584 585
R165 B.n586 B.n585 585
R166 B.n583 B.n288 585
R167 B.n288 B.n287 585
R168 B.n582 B.n581 585
R169 B.n581 B.n580 585
R170 B.n290 B.n289 585
R171 B.n291 B.n290 585
R172 B.n573 B.n572 585
R173 B.n574 B.n573 585
R174 B.n571 B.n296 585
R175 B.n296 B.n295 585
R176 B.n570 B.n569 585
R177 B.n569 B.n568 585
R178 B.n298 B.n297 585
R179 B.n561 B.n298 585
R180 B.n560 B.n559 585
R181 B.n562 B.n560 585
R182 B.n558 B.n303 585
R183 B.n303 B.n302 585
R184 B.n557 B.n556 585
R185 B.n556 B.n555 585
R186 B.n305 B.n304 585
R187 B.n306 B.n305 585
R188 B.n548 B.n547 585
R189 B.n549 B.n548 585
R190 B.n546 B.n311 585
R191 B.n311 B.n310 585
R192 B.n540 B.n539 585
R193 B.n538 B.n358 585
R194 B.n537 B.n357 585
R195 B.n542 B.n357 585
R196 B.n536 B.n535 585
R197 B.n534 B.n533 585
R198 B.n532 B.n531 585
R199 B.n530 B.n529 585
R200 B.n528 B.n527 585
R201 B.n526 B.n525 585
R202 B.n524 B.n523 585
R203 B.n522 B.n521 585
R204 B.n520 B.n519 585
R205 B.n518 B.n517 585
R206 B.n516 B.n515 585
R207 B.n514 B.n513 585
R208 B.n512 B.n511 585
R209 B.n510 B.n509 585
R210 B.n508 B.n507 585
R211 B.n506 B.n505 585
R212 B.n504 B.n503 585
R213 B.n502 B.n501 585
R214 B.n500 B.n499 585
R215 B.n498 B.n497 585
R216 B.n496 B.n495 585
R217 B.n494 B.n493 585
R218 B.n492 B.n491 585
R219 B.n490 B.n489 585
R220 B.n488 B.n487 585
R221 B.n486 B.n485 585
R222 B.n484 B.n483 585
R223 B.n482 B.n481 585
R224 B.n480 B.n479 585
R225 B.n478 B.n477 585
R226 B.n476 B.n475 585
R227 B.n474 B.n473 585
R228 B.n472 B.n471 585
R229 B.n470 B.n469 585
R230 B.n468 B.n467 585
R231 B.n466 B.n465 585
R232 B.n464 B.n463 585
R233 B.n462 B.n461 585
R234 B.n460 B.n459 585
R235 B.n458 B.n457 585
R236 B.n456 B.n455 585
R237 B.n454 B.n453 585
R238 B.n452 B.n451 585
R239 B.n450 B.n449 585
R240 B.n448 B.n447 585
R241 B.n446 B.n445 585
R242 B.n444 B.n443 585
R243 B.n441 B.n440 585
R244 B.n439 B.n438 585
R245 B.n437 B.n436 585
R246 B.n435 B.n434 585
R247 B.n433 B.n432 585
R248 B.n431 B.n430 585
R249 B.n429 B.n428 585
R250 B.n427 B.n426 585
R251 B.n425 B.n424 585
R252 B.n423 B.n422 585
R253 B.n421 B.n420 585
R254 B.n419 B.n418 585
R255 B.n417 B.n416 585
R256 B.n415 B.n414 585
R257 B.n413 B.n412 585
R258 B.n411 B.n410 585
R259 B.n409 B.n408 585
R260 B.n407 B.n406 585
R261 B.n405 B.n404 585
R262 B.n403 B.n402 585
R263 B.n401 B.n400 585
R264 B.n399 B.n398 585
R265 B.n397 B.n396 585
R266 B.n395 B.n394 585
R267 B.n393 B.n392 585
R268 B.n391 B.n390 585
R269 B.n389 B.n388 585
R270 B.n387 B.n386 585
R271 B.n385 B.n384 585
R272 B.n383 B.n382 585
R273 B.n381 B.n380 585
R274 B.n379 B.n378 585
R275 B.n377 B.n376 585
R276 B.n375 B.n374 585
R277 B.n373 B.n372 585
R278 B.n371 B.n370 585
R279 B.n369 B.n368 585
R280 B.n367 B.n366 585
R281 B.n365 B.n364 585
R282 B.n313 B.n312 585
R283 B.n545 B.n544 585
R284 B.n309 B.n308 585
R285 B.n310 B.n309 585
R286 B.n551 B.n550 585
R287 B.n550 B.n549 585
R288 B.n552 B.n307 585
R289 B.n307 B.n306 585
R290 B.n554 B.n553 585
R291 B.n555 B.n554 585
R292 B.n301 B.n300 585
R293 B.n302 B.n301 585
R294 B.n564 B.n563 585
R295 B.n563 B.n562 585
R296 B.n565 B.n299 585
R297 B.n561 B.n299 585
R298 B.n567 B.n566 585
R299 B.n568 B.n567 585
R300 B.n294 B.n293 585
R301 B.n295 B.n294 585
R302 B.n576 B.n575 585
R303 B.n575 B.n574 585
R304 B.n577 B.n292 585
R305 B.n292 B.n291 585
R306 B.n579 B.n578 585
R307 B.n580 B.n579 585
R308 B.n286 B.n285 585
R309 B.n287 B.n286 585
R310 B.n588 B.n587 585
R311 B.n587 B.n586 585
R312 B.n589 B.n284 585
R313 B.n284 B.n282 585
R314 B.n591 B.n590 585
R315 B.n592 B.n591 585
R316 B.n278 B.n277 585
R317 B.n283 B.n278 585
R318 B.n601 B.n600 585
R319 B.n600 B.n599 585
R320 B.n602 B.n276 585
R321 B.n276 B.n275 585
R322 B.n604 B.n603 585
R323 B.n605 B.n604 585
R324 B.n2 B.n0 585
R325 B.n4 B.n2 585
R326 B.n3 B.n1 585
R327 B.n679 B.n3 585
R328 B.n677 B.n676 585
R329 B.n678 B.n677 585
R330 B.n675 B.n9 585
R331 B.n9 B.n8 585
R332 B.n674 B.n673 585
R333 B.n673 B.n672 585
R334 B.n11 B.n10 585
R335 B.n671 B.n11 585
R336 B.n669 B.n668 585
R337 B.n670 B.n669 585
R338 B.n667 B.n16 585
R339 B.n16 B.n15 585
R340 B.n666 B.n665 585
R341 B.n665 B.n664 585
R342 B.n18 B.n17 585
R343 B.n663 B.n18 585
R344 B.n661 B.n660 585
R345 B.n662 B.n661 585
R346 B.n659 B.n23 585
R347 B.n23 B.n22 585
R348 B.n658 B.n657 585
R349 B.n657 B.n656 585
R350 B.n25 B.n24 585
R351 B.n655 B.n25 585
R352 B.n653 B.n652 585
R353 B.n654 B.n653 585
R354 B.n651 B.n29 585
R355 B.n32 B.n29 585
R356 B.n650 B.n649 585
R357 B.n649 B.n648 585
R358 B.n31 B.n30 585
R359 B.n647 B.n31 585
R360 B.n645 B.n644 585
R361 B.n646 B.n645 585
R362 B.n643 B.n37 585
R363 B.n37 B.n36 585
R364 B.n642 B.n641 585
R365 B.n641 B.n640 585
R366 B.n39 B.n38 585
R367 B.n639 B.n39 585
R368 B.n682 B.n681 585
R369 B.n681 B.n680 585
R370 B.n540 B.n309 506.916
R371 B.n93 B.n39 506.916
R372 B.n544 B.n311 506.916
R373 B.n637 B.n41 506.916
R374 B.n362 B.t6 354.19
R375 B.n359 B.t10 354.19
R376 B.n91 B.t13 354.19
R377 B.n88 B.t2 354.19
R378 B.n638 B.n86 256.663
R379 B.n638 B.n85 256.663
R380 B.n638 B.n84 256.663
R381 B.n638 B.n83 256.663
R382 B.n638 B.n82 256.663
R383 B.n638 B.n81 256.663
R384 B.n638 B.n80 256.663
R385 B.n638 B.n79 256.663
R386 B.n638 B.n78 256.663
R387 B.n638 B.n77 256.663
R388 B.n638 B.n76 256.663
R389 B.n638 B.n75 256.663
R390 B.n638 B.n74 256.663
R391 B.n638 B.n73 256.663
R392 B.n638 B.n72 256.663
R393 B.n638 B.n71 256.663
R394 B.n638 B.n70 256.663
R395 B.n638 B.n69 256.663
R396 B.n638 B.n68 256.663
R397 B.n638 B.n67 256.663
R398 B.n638 B.n66 256.663
R399 B.n638 B.n65 256.663
R400 B.n638 B.n64 256.663
R401 B.n638 B.n63 256.663
R402 B.n638 B.n62 256.663
R403 B.n638 B.n61 256.663
R404 B.n638 B.n60 256.663
R405 B.n638 B.n59 256.663
R406 B.n638 B.n58 256.663
R407 B.n638 B.n57 256.663
R408 B.n638 B.n56 256.663
R409 B.n638 B.n55 256.663
R410 B.n638 B.n54 256.663
R411 B.n638 B.n53 256.663
R412 B.n638 B.n52 256.663
R413 B.n638 B.n51 256.663
R414 B.n638 B.n50 256.663
R415 B.n638 B.n49 256.663
R416 B.n638 B.n48 256.663
R417 B.n638 B.n47 256.663
R418 B.n638 B.n46 256.663
R419 B.n638 B.n45 256.663
R420 B.n638 B.n44 256.663
R421 B.n638 B.n43 256.663
R422 B.n638 B.n42 256.663
R423 B.n542 B.n541 256.663
R424 B.n542 B.n314 256.663
R425 B.n542 B.n315 256.663
R426 B.n542 B.n316 256.663
R427 B.n542 B.n317 256.663
R428 B.n542 B.n318 256.663
R429 B.n542 B.n319 256.663
R430 B.n542 B.n320 256.663
R431 B.n542 B.n321 256.663
R432 B.n542 B.n322 256.663
R433 B.n542 B.n323 256.663
R434 B.n542 B.n324 256.663
R435 B.n542 B.n325 256.663
R436 B.n542 B.n326 256.663
R437 B.n542 B.n327 256.663
R438 B.n542 B.n328 256.663
R439 B.n542 B.n329 256.663
R440 B.n542 B.n330 256.663
R441 B.n542 B.n331 256.663
R442 B.n542 B.n332 256.663
R443 B.n542 B.n333 256.663
R444 B.n542 B.n334 256.663
R445 B.n542 B.n335 256.663
R446 B.n542 B.n336 256.663
R447 B.n542 B.n337 256.663
R448 B.n542 B.n338 256.663
R449 B.n542 B.n339 256.663
R450 B.n542 B.n340 256.663
R451 B.n542 B.n341 256.663
R452 B.n542 B.n342 256.663
R453 B.n542 B.n343 256.663
R454 B.n542 B.n344 256.663
R455 B.n542 B.n345 256.663
R456 B.n542 B.n346 256.663
R457 B.n542 B.n347 256.663
R458 B.n542 B.n348 256.663
R459 B.n542 B.n349 256.663
R460 B.n542 B.n350 256.663
R461 B.n542 B.n351 256.663
R462 B.n542 B.n352 256.663
R463 B.n542 B.n353 256.663
R464 B.n542 B.n354 256.663
R465 B.n542 B.n355 256.663
R466 B.n542 B.n356 256.663
R467 B.n543 B.n542 256.663
R468 B.n550 B.n309 163.367
R469 B.n550 B.n307 163.367
R470 B.n554 B.n307 163.367
R471 B.n554 B.n301 163.367
R472 B.n563 B.n301 163.367
R473 B.n563 B.n299 163.367
R474 B.n567 B.n299 163.367
R475 B.n567 B.n294 163.367
R476 B.n575 B.n294 163.367
R477 B.n575 B.n292 163.367
R478 B.n579 B.n292 163.367
R479 B.n579 B.n286 163.367
R480 B.n587 B.n286 163.367
R481 B.n587 B.n284 163.367
R482 B.n591 B.n284 163.367
R483 B.n591 B.n278 163.367
R484 B.n600 B.n278 163.367
R485 B.n600 B.n276 163.367
R486 B.n604 B.n276 163.367
R487 B.n604 B.n2 163.367
R488 B.n681 B.n2 163.367
R489 B.n681 B.n3 163.367
R490 B.n677 B.n3 163.367
R491 B.n677 B.n9 163.367
R492 B.n673 B.n9 163.367
R493 B.n673 B.n11 163.367
R494 B.n669 B.n11 163.367
R495 B.n669 B.n16 163.367
R496 B.n665 B.n16 163.367
R497 B.n665 B.n18 163.367
R498 B.n661 B.n18 163.367
R499 B.n661 B.n23 163.367
R500 B.n657 B.n23 163.367
R501 B.n657 B.n25 163.367
R502 B.n653 B.n25 163.367
R503 B.n653 B.n29 163.367
R504 B.n649 B.n29 163.367
R505 B.n649 B.n31 163.367
R506 B.n645 B.n31 163.367
R507 B.n645 B.n37 163.367
R508 B.n641 B.n37 163.367
R509 B.n641 B.n39 163.367
R510 B.n358 B.n357 163.367
R511 B.n535 B.n357 163.367
R512 B.n533 B.n532 163.367
R513 B.n529 B.n528 163.367
R514 B.n525 B.n524 163.367
R515 B.n521 B.n520 163.367
R516 B.n517 B.n516 163.367
R517 B.n513 B.n512 163.367
R518 B.n509 B.n508 163.367
R519 B.n505 B.n504 163.367
R520 B.n501 B.n500 163.367
R521 B.n497 B.n496 163.367
R522 B.n493 B.n492 163.367
R523 B.n489 B.n488 163.367
R524 B.n485 B.n484 163.367
R525 B.n481 B.n480 163.367
R526 B.n477 B.n476 163.367
R527 B.n473 B.n472 163.367
R528 B.n469 B.n468 163.367
R529 B.n465 B.n464 163.367
R530 B.n461 B.n460 163.367
R531 B.n457 B.n456 163.367
R532 B.n453 B.n452 163.367
R533 B.n449 B.n448 163.367
R534 B.n445 B.n444 163.367
R535 B.n440 B.n439 163.367
R536 B.n436 B.n435 163.367
R537 B.n432 B.n431 163.367
R538 B.n428 B.n427 163.367
R539 B.n424 B.n423 163.367
R540 B.n420 B.n419 163.367
R541 B.n416 B.n415 163.367
R542 B.n412 B.n411 163.367
R543 B.n408 B.n407 163.367
R544 B.n404 B.n403 163.367
R545 B.n400 B.n399 163.367
R546 B.n396 B.n395 163.367
R547 B.n392 B.n391 163.367
R548 B.n388 B.n387 163.367
R549 B.n384 B.n383 163.367
R550 B.n380 B.n379 163.367
R551 B.n376 B.n375 163.367
R552 B.n372 B.n371 163.367
R553 B.n368 B.n367 163.367
R554 B.n364 B.n313 163.367
R555 B.n548 B.n311 163.367
R556 B.n548 B.n305 163.367
R557 B.n556 B.n305 163.367
R558 B.n556 B.n303 163.367
R559 B.n560 B.n303 163.367
R560 B.n560 B.n298 163.367
R561 B.n569 B.n298 163.367
R562 B.n569 B.n296 163.367
R563 B.n573 B.n296 163.367
R564 B.n573 B.n290 163.367
R565 B.n581 B.n290 163.367
R566 B.n581 B.n288 163.367
R567 B.n585 B.n288 163.367
R568 B.n585 B.n281 163.367
R569 B.n593 B.n281 163.367
R570 B.n593 B.n279 163.367
R571 B.n598 B.n279 163.367
R572 B.n598 B.n274 163.367
R573 B.n606 B.n274 163.367
R574 B.n607 B.n606 163.367
R575 B.n607 B.n5 163.367
R576 B.n6 B.n5 163.367
R577 B.n7 B.n6 163.367
R578 B.n612 B.n7 163.367
R579 B.n612 B.n12 163.367
R580 B.n13 B.n12 163.367
R581 B.n14 B.n13 163.367
R582 B.n617 B.n14 163.367
R583 B.n617 B.n19 163.367
R584 B.n20 B.n19 163.367
R585 B.n21 B.n20 163.367
R586 B.n622 B.n21 163.367
R587 B.n622 B.n26 163.367
R588 B.n27 B.n26 163.367
R589 B.n28 B.n27 163.367
R590 B.n627 B.n28 163.367
R591 B.n627 B.n33 163.367
R592 B.n34 B.n33 163.367
R593 B.n35 B.n34 163.367
R594 B.n632 B.n35 163.367
R595 B.n632 B.n40 163.367
R596 B.n41 B.n40 163.367
R597 B.n97 B.n96 163.367
R598 B.n101 B.n100 163.367
R599 B.n105 B.n104 163.367
R600 B.n109 B.n108 163.367
R601 B.n113 B.n112 163.367
R602 B.n117 B.n116 163.367
R603 B.n121 B.n120 163.367
R604 B.n125 B.n124 163.367
R605 B.n129 B.n128 163.367
R606 B.n133 B.n132 163.367
R607 B.n137 B.n136 163.367
R608 B.n141 B.n140 163.367
R609 B.n145 B.n144 163.367
R610 B.n149 B.n148 163.367
R611 B.n153 B.n152 163.367
R612 B.n157 B.n156 163.367
R613 B.n161 B.n160 163.367
R614 B.n165 B.n164 163.367
R615 B.n169 B.n168 163.367
R616 B.n173 B.n172 163.367
R617 B.n178 B.n177 163.367
R618 B.n182 B.n181 163.367
R619 B.n186 B.n185 163.367
R620 B.n190 B.n189 163.367
R621 B.n194 B.n193 163.367
R622 B.n198 B.n197 163.367
R623 B.n202 B.n201 163.367
R624 B.n206 B.n205 163.367
R625 B.n210 B.n209 163.367
R626 B.n214 B.n213 163.367
R627 B.n218 B.n217 163.367
R628 B.n222 B.n221 163.367
R629 B.n226 B.n225 163.367
R630 B.n230 B.n229 163.367
R631 B.n234 B.n233 163.367
R632 B.n238 B.n237 163.367
R633 B.n242 B.n241 163.367
R634 B.n246 B.n245 163.367
R635 B.n250 B.n249 163.367
R636 B.n254 B.n253 163.367
R637 B.n258 B.n257 163.367
R638 B.n262 B.n261 163.367
R639 B.n266 B.n265 163.367
R640 B.n270 B.n269 163.367
R641 B.n637 B.n87 163.367
R642 B.n362 B.t9 112.448
R643 B.n88 B.t4 112.448
R644 B.n359 B.t12 112.433
R645 B.n91 B.t14 112.433
R646 B.n542 B.n310 90.4471
R647 B.n639 B.n638 90.4471
R648 B.n541 B.n540 71.676
R649 B.n535 B.n314 71.676
R650 B.n532 B.n315 71.676
R651 B.n528 B.n316 71.676
R652 B.n524 B.n317 71.676
R653 B.n520 B.n318 71.676
R654 B.n516 B.n319 71.676
R655 B.n512 B.n320 71.676
R656 B.n508 B.n321 71.676
R657 B.n504 B.n322 71.676
R658 B.n500 B.n323 71.676
R659 B.n496 B.n324 71.676
R660 B.n492 B.n325 71.676
R661 B.n488 B.n326 71.676
R662 B.n484 B.n327 71.676
R663 B.n480 B.n328 71.676
R664 B.n476 B.n329 71.676
R665 B.n472 B.n330 71.676
R666 B.n468 B.n331 71.676
R667 B.n464 B.n332 71.676
R668 B.n460 B.n333 71.676
R669 B.n456 B.n334 71.676
R670 B.n452 B.n335 71.676
R671 B.n448 B.n336 71.676
R672 B.n444 B.n337 71.676
R673 B.n439 B.n338 71.676
R674 B.n435 B.n339 71.676
R675 B.n431 B.n340 71.676
R676 B.n427 B.n341 71.676
R677 B.n423 B.n342 71.676
R678 B.n419 B.n343 71.676
R679 B.n415 B.n344 71.676
R680 B.n411 B.n345 71.676
R681 B.n407 B.n346 71.676
R682 B.n403 B.n347 71.676
R683 B.n399 B.n348 71.676
R684 B.n395 B.n349 71.676
R685 B.n391 B.n350 71.676
R686 B.n387 B.n351 71.676
R687 B.n383 B.n352 71.676
R688 B.n379 B.n353 71.676
R689 B.n375 B.n354 71.676
R690 B.n371 B.n355 71.676
R691 B.n367 B.n356 71.676
R692 B.n543 B.n313 71.676
R693 B.n93 B.n42 71.676
R694 B.n97 B.n43 71.676
R695 B.n101 B.n44 71.676
R696 B.n105 B.n45 71.676
R697 B.n109 B.n46 71.676
R698 B.n113 B.n47 71.676
R699 B.n117 B.n48 71.676
R700 B.n121 B.n49 71.676
R701 B.n125 B.n50 71.676
R702 B.n129 B.n51 71.676
R703 B.n133 B.n52 71.676
R704 B.n137 B.n53 71.676
R705 B.n141 B.n54 71.676
R706 B.n145 B.n55 71.676
R707 B.n149 B.n56 71.676
R708 B.n153 B.n57 71.676
R709 B.n157 B.n58 71.676
R710 B.n161 B.n59 71.676
R711 B.n165 B.n60 71.676
R712 B.n169 B.n61 71.676
R713 B.n173 B.n62 71.676
R714 B.n178 B.n63 71.676
R715 B.n182 B.n64 71.676
R716 B.n186 B.n65 71.676
R717 B.n190 B.n66 71.676
R718 B.n194 B.n67 71.676
R719 B.n198 B.n68 71.676
R720 B.n202 B.n69 71.676
R721 B.n206 B.n70 71.676
R722 B.n210 B.n71 71.676
R723 B.n214 B.n72 71.676
R724 B.n218 B.n73 71.676
R725 B.n222 B.n74 71.676
R726 B.n226 B.n75 71.676
R727 B.n230 B.n76 71.676
R728 B.n234 B.n77 71.676
R729 B.n238 B.n78 71.676
R730 B.n242 B.n79 71.676
R731 B.n246 B.n80 71.676
R732 B.n250 B.n81 71.676
R733 B.n254 B.n82 71.676
R734 B.n258 B.n83 71.676
R735 B.n262 B.n84 71.676
R736 B.n266 B.n85 71.676
R737 B.n270 B.n86 71.676
R738 B.n87 B.n86 71.676
R739 B.n269 B.n85 71.676
R740 B.n265 B.n84 71.676
R741 B.n261 B.n83 71.676
R742 B.n257 B.n82 71.676
R743 B.n253 B.n81 71.676
R744 B.n249 B.n80 71.676
R745 B.n245 B.n79 71.676
R746 B.n241 B.n78 71.676
R747 B.n237 B.n77 71.676
R748 B.n233 B.n76 71.676
R749 B.n229 B.n75 71.676
R750 B.n225 B.n74 71.676
R751 B.n221 B.n73 71.676
R752 B.n217 B.n72 71.676
R753 B.n213 B.n71 71.676
R754 B.n209 B.n70 71.676
R755 B.n205 B.n69 71.676
R756 B.n201 B.n68 71.676
R757 B.n197 B.n67 71.676
R758 B.n193 B.n66 71.676
R759 B.n189 B.n65 71.676
R760 B.n185 B.n64 71.676
R761 B.n181 B.n63 71.676
R762 B.n177 B.n62 71.676
R763 B.n172 B.n61 71.676
R764 B.n168 B.n60 71.676
R765 B.n164 B.n59 71.676
R766 B.n160 B.n58 71.676
R767 B.n156 B.n57 71.676
R768 B.n152 B.n56 71.676
R769 B.n148 B.n55 71.676
R770 B.n144 B.n54 71.676
R771 B.n140 B.n53 71.676
R772 B.n136 B.n52 71.676
R773 B.n132 B.n51 71.676
R774 B.n128 B.n50 71.676
R775 B.n124 B.n49 71.676
R776 B.n120 B.n48 71.676
R777 B.n116 B.n47 71.676
R778 B.n112 B.n46 71.676
R779 B.n108 B.n45 71.676
R780 B.n104 B.n44 71.676
R781 B.n100 B.n43 71.676
R782 B.n96 B.n42 71.676
R783 B.n541 B.n358 71.676
R784 B.n533 B.n314 71.676
R785 B.n529 B.n315 71.676
R786 B.n525 B.n316 71.676
R787 B.n521 B.n317 71.676
R788 B.n517 B.n318 71.676
R789 B.n513 B.n319 71.676
R790 B.n509 B.n320 71.676
R791 B.n505 B.n321 71.676
R792 B.n501 B.n322 71.676
R793 B.n497 B.n323 71.676
R794 B.n493 B.n324 71.676
R795 B.n489 B.n325 71.676
R796 B.n485 B.n326 71.676
R797 B.n481 B.n327 71.676
R798 B.n477 B.n328 71.676
R799 B.n473 B.n329 71.676
R800 B.n469 B.n330 71.676
R801 B.n465 B.n331 71.676
R802 B.n461 B.n332 71.676
R803 B.n457 B.n333 71.676
R804 B.n453 B.n334 71.676
R805 B.n449 B.n335 71.676
R806 B.n445 B.n336 71.676
R807 B.n440 B.n337 71.676
R808 B.n436 B.n338 71.676
R809 B.n432 B.n339 71.676
R810 B.n428 B.n340 71.676
R811 B.n424 B.n341 71.676
R812 B.n420 B.n342 71.676
R813 B.n416 B.n343 71.676
R814 B.n412 B.n344 71.676
R815 B.n408 B.n345 71.676
R816 B.n404 B.n346 71.676
R817 B.n400 B.n347 71.676
R818 B.n396 B.n348 71.676
R819 B.n392 B.n349 71.676
R820 B.n388 B.n350 71.676
R821 B.n384 B.n351 71.676
R822 B.n380 B.n352 71.676
R823 B.n376 B.n353 71.676
R824 B.n372 B.n354 71.676
R825 B.n368 B.n355 71.676
R826 B.n364 B.n356 71.676
R827 B.n544 B.n543 71.676
R828 B.n363 B.t8 69.1995
R829 B.n89 B.t5 69.1995
R830 B.n360 B.t11 69.1847
R831 B.n92 B.t15 69.1847
R832 B.n442 B.n363 59.5399
R833 B.n361 B.n360 59.5399
R834 B.n175 B.n92 59.5399
R835 B.n90 B.n89 59.5399
R836 B.n549 B.n310 44.2478
R837 B.n549 B.n306 44.2478
R838 B.n555 B.n306 44.2478
R839 B.n555 B.n302 44.2478
R840 B.n562 B.n302 44.2478
R841 B.n562 B.n561 44.2478
R842 B.n568 B.n295 44.2478
R843 B.n574 B.n295 44.2478
R844 B.n574 B.n291 44.2478
R845 B.n580 B.n291 44.2478
R846 B.n580 B.n287 44.2478
R847 B.n586 B.n287 44.2478
R848 B.n586 B.n282 44.2478
R849 B.n592 B.n282 44.2478
R850 B.n592 B.n283 44.2478
R851 B.n599 B.n275 44.2478
R852 B.n605 B.n275 44.2478
R853 B.n605 B.n4 44.2478
R854 B.n680 B.n4 44.2478
R855 B.n680 B.n679 44.2478
R856 B.n679 B.n678 44.2478
R857 B.n678 B.n8 44.2478
R858 B.n672 B.n8 44.2478
R859 B.n671 B.n670 44.2478
R860 B.n670 B.n15 44.2478
R861 B.n664 B.n15 44.2478
R862 B.n664 B.n663 44.2478
R863 B.n663 B.n662 44.2478
R864 B.n662 B.n22 44.2478
R865 B.n656 B.n22 44.2478
R866 B.n656 B.n655 44.2478
R867 B.n655 B.n654 44.2478
R868 B.n648 B.n32 44.2478
R869 B.n648 B.n647 44.2478
R870 B.n647 B.n646 44.2478
R871 B.n646 B.n36 44.2478
R872 B.n640 B.n36 44.2478
R873 B.n640 B.n639 44.2478
R874 B.n363 B.n362 43.249
R875 B.n360 B.n359 43.249
R876 B.n92 B.n91 43.249
R877 B.n89 B.n88 43.249
R878 B.n599 B.t1 39.0422
R879 B.n672 B.t0 39.0422
R880 B.n94 B.n38 32.9371
R881 B.n636 B.n635 32.9371
R882 B.n546 B.n545 32.9371
R883 B.n539 B.n308 32.9371
R884 B.n568 B.t7 28.6311
R885 B.n654 B.t3 28.6311
R886 B B.n682 18.0485
R887 B.n561 B.t7 15.6172
R888 B.n32 B.t3 15.6172
R889 B.n95 B.n94 10.6151
R890 B.n98 B.n95 10.6151
R891 B.n99 B.n98 10.6151
R892 B.n102 B.n99 10.6151
R893 B.n103 B.n102 10.6151
R894 B.n106 B.n103 10.6151
R895 B.n107 B.n106 10.6151
R896 B.n110 B.n107 10.6151
R897 B.n111 B.n110 10.6151
R898 B.n114 B.n111 10.6151
R899 B.n115 B.n114 10.6151
R900 B.n118 B.n115 10.6151
R901 B.n119 B.n118 10.6151
R902 B.n122 B.n119 10.6151
R903 B.n123 B.n122 10.6151
R904 B.n126 B.n123 10.6151
R905 B.n127 B.n126 10.6151
R906 B.n130 B.n127 10.6151
R907 B.n131 B.n130 10.6151
R908 B.n134 B.n131 10.6151
R909 B.n135 B.n134 10.6151
R910 B.n138 B.n135 10.6151
R911 B.n139 B.n138 10.6151
R912 B.n142 B.n139 10.6151
R913 B.n143 B.n142 10.6151
R914 B.n146 B.n143 10.6151
R915 B.n147 B.n146 10.6151
R916 B.n150 B.n147 10.6151
R917 B.n151 B.n150 10.6151
R918 B.n154 B.n151 10.6151
R919 B.n155 B.n154 10.6151
R920 B.n158 B.n155 10.6151
R921 B.n159 B.n158 10.6151
R922 B.n162 B.n159 10.6151
R923 B.n163 B.n162 10.6151
R924 B.n166 B.n163 10.6151
R925 B.n167 B.n166 10.6151
R926 B.n170 B.n167 10.6151
R927 B.n171 B.n170 10.6151
R928 B.n174 B.n171 10.6151
R929 B.n179 B.n176 10.6151
R930 B.n180 B.n179 10.6151
R931 B.n183 B.n180 10.6151
R932 B.n184 B.n183 10.6151
R933 B.n187 B.n184 10.6151
R934 B.n188 B.n187 10.6151
R935 B.n191 B.n188 10.6151
R936 B.n192 B.n191 10.6151
R937 B.n196 B.n195 10.6151
R938 B.n199 B.n196 10.6151
R939 B.n200 B.n199 10.6151
R940 B.n203 B.n200 10.6151
R941 B.n204 B.n203 10.6151
R942 B.n207 B.n204 10.6151
R943 B.n208 B.n207 10.6151
R944 B.n211 B.n208 10.6151
R945 B.n212 B.n211 10.6151
R946 B.n215 B.n212 10.6151
R947 B.n216 B.n215 10.6151
R948 B.n219 B.n216 10.6151
R949 B.n220 B.n219 10.6151
R950 B.n223 B.n220 10.6151
R951 B.n224 B.n223 10.6151
R952 B.n227 B.n224 10.6151
R953 B.n228 B.n227 10.6151
R954 B.n231 B.n228 10.6151
R955 B.n232 B.n231 10.6151
R956 B.n235 B.n232 10.6151
R957 B.n236 B.n235 10.6151
R958 B.n239 B.n236 10.6151
R959 B.n240 B.n239 10.6151
R960 B.n243 B.n240 10.6151
R961 B.n244 B.n243 10.6151
R962 B.n247 B.n244 10.6151
R963 B.n248 B.n247 10.6151
R964 B.n251 B.n248 10.6151
R965 B.n252 B.n251 10.6151
R966 B.n255 B.n252 10.6151
R967 B.n256 B.n255 10.6151
R968 B.n259 B.n256 10.6151
R969 B.n260 B.n259 10.6151
R970 B.n263 B.n260 10.6151
R971 B.n264 B.n263 10.6151
R972 B.n267 B.n264 10.6151
R973 B.n268 B.n267 10.6151
R974 B.n271 B.n268 10.6151
R975 B.n272 B.n271 10.6151
R976 B.n636 B.n272 10.6151
R977 B.n547 B.n546 10.6151
R978 B.n547 B.n304 10.6151
R979 B.n557 B.n304 10.6151
R980 B.n558 B.n557 10.6151
R981 B.n559 B.n558 10.6151
R982 B.n559 B.n297 10.6151
R983 B.n570 B.n297 10.6151
R984 B.n571 B.n570 10.6151
R985 B.n572 B.n571 10.6151
R986 B.n572 B.n289 10.6151
R987 B.n582 B.n289 10.6151
R988 B.n583 B.n582 10.6151
R989 B.n584 B.n583 10.6151
R990 B.n584 B.n280 10.6151
R991 B.n594 B.n280 10.6151
R992 B.n595 B.n594 10.6151
R993 B.n597 B.n595 10.6151
R994 B.n597 B.n596 10.6151
R995 B.n596 B.n273 10.6151
R996 B.n608 B.n273 10.6151
R997 B.n609 B.n608 10.6151
R998 B.n610 B.n609 10.6151
R999 B.n611 B.n610 10.6151
R1000 B.n613 B.n611 10.6151
R1001 B.n614 B.n613 10.6151
R1002 B.n615 B.n614 10.6151
R1003 B.n616 B.n615 10.6151
R1004 B.n618 B.n616 10.6151
R1005 B.n619 B.n618 10.6151
R1006 B.n620 B.n619 10.6151
R1007 B.n621 B.n620 10.6151
R1008 B.n623 B.n621 10.6151
R1009 B.n624 B.n623 10.6151
R1010 B.n625 B.n624 10.6151
R1011 B.n626 B.n625 10.6151
R1012 B.n628 B.n626 10.6151
R1013 B.n629 B.n628 10.6151
R1014 B.n630 B.n629 10.6151
R1015 B.n631 B.n630 10.6151
R1016 B.n633 B.n631 10.6151
R1017 B.n634 B.n633 10.6151
R1018 B.n635 B.n634 10.6151
R1019 B.n539 B.n538 10.6151
R1020 B.n538 B.n537 10.6151
R1021 B.n537 B.n536 10.6151
R1022 B.n536 B.n534 10.6151
R1023 B.n534 B.n531 10.6151
R1024 B.n531 B.n530 10.6151
R1025 B.n530 B.n527 10.6151
R1026 B.n527 B.n526 10.6151
R1027 B.n526 B.n523 10.6151
R1028 B.n523 B.n522 10.6151
R1029 B.n522 B.n519 10.6151
R1030 B.n519 B.n518 10.6151
R1031 B.n518 B.n515 10.6151
R1032 B.n515 B.n514 10.6151
R1033 B.n514 B.n511 10.6151
R1034 B.n511 B.n510 10.6151
R1035 B.n510 B.n507 10.6151
R1036 B.n507 B.n506 10.6151
R1037 B.n506 B.n503 10.6151
R1038 B.n503 B.n502 10.6151
R1039 B.n502 B.n499 10.6151
R1040 B.n499 B.n498 10.6151
R1041 B.n498 B.n495 10.6151
R1042 B.n495 B.n494 10.6151
R1043 B.n494 B.n491 10.6151
R1044 B.n491 B.n490 10.6151
R1045 B.n490 B.n487 10.6151
R1046 B.n487 B.n486 10.6151
R1047 B.n486 B.n483 10.6151
R1048 B.n483 B.n482 10.6151
R1049 B.n482 B.n479 10.6151
R1050 B.n479 B.n478 10.6151
R1051 B.n478 B.n475 10.6151
R1052 B.n475 B.n474 10.6151
R1053 B.n474 B.n471 10.6151
R1054 B.n471 B.n470 10.6151
R1055 B.n470 B.n467 10.6151
R1056 B.n467 B.n466 10.6151
R1057 B.n466 B.n463 10.6151
R1058 B.n463 B.n462 10.6151
R1059 B.n459 B.n458 10.6151
R1060 B.n458 B.n455 10.6151
R1061 B.n455 B.n454 10.6151
R1062 B.n454 B.n451 10.6151
R1063 B.n451 B.n450 10.6151
R1064 B.n450 B.n447 10.6151
R1065 B.n447 B.n446 10.6151
R1066 B.n446 B.n443 10.6151
R1067 B.n441 B.n438 10.6151
R1068 B.n438 B.n437 10.6151
R1069 B.n437 B.n434 10.6151
R1070 B.n434 B.n433 10.6151
R1071 B.n433 B.n430 10.6151
R1072 B.n430 B.n429 10.6151
R1073 B.n429 B.n426 10.6151
R1074 B.n426 B.n425 10.6151
R1075 B.n425 B.n422 10.6151
R1076 B.n422 B.n421 10.6151
R1077 B.n421 B.n418 10.6151
R1078 B.n418 B.n417 10.6151
R1079 B.n417 B.n414 10.6151
R1080 B.n414 B.n413 10.6151
R1081 B.n413 B.n410 10.6151
R1082 B.n410 B.n409 10.6151
R1083 B.n409 B.n406 10.6151
R1084 B.n406 B.n405 10.6151
R1085 B.n405 B.n402 10.6151
R1086 B.n402 B.n401 10.6151
R1087 B.n401 B.n398 10.6151
R1088 B.n398 B.n397 10.6151
R1089 B.n397 B.n394 10.6151
R1090 B.n394 B.n393 10.6151
R1091 B.n393 B.n390 10.6151
R1092 B.n390 B.n389 10.6151
R1093 B.n389 B.n386 10.6151
R1094 B.n386 B.n385 10.6151
R1095 B.n385 B.n382 10.6151
R1096 B.n382 B.n381 10.6151
R1097 B.n381 B.n378 10.6151
R1098 B.n378 B.n377 10.6151
R1099 B.n377 B.n374 10.6151
R1100 B.n374 B.n373 10.6151
R1101 B.n373 B.n370 10.6151
R1102 B.n370 B.n369 10.6151
R1103 B.n369 B.n366 10.6151
R1104 B.n366 B.n365 10.6151
R1105 B.n365 B.n312 10.6151
R1106 B.n545 B.n312 10.6151
R1107 B.n551 B.n308 10.6151
R1108 B.n552 B.n551 10.6151
R1109 B.n553 B.n552 10.6151
R1110 B.n553 B.n300 10.6151
R1111 B.n564 B.n300 10.6151
R1112 B.n565 B.n564 10.6151
R1113 B.n566 B.n565 10.6151
R1114 B.n566 B.n293 10.6151
R1115 B.n576 B.n293 10.6151
R1116 B.n577 B.n576 10.6151
R1117 B.n578 B.n577 10.6151
R1118 B.n578 B.n285 10.6151
R1119 B.n588 B.n285 10.6151
R1120 B.n589 B.n588 10.6151
R1121 B.n590 B.n589 10.6151
R1122 B.n590 B.n277 10.6151
R1123 B.n601 B.n277 10.6151
R1124 B.n602 B.n601 10.6151
R1125 B.n603 B.n602 10.6151
R1126 B.n603 B.n0 10.6151
R1127 B.n676 B.n1 10.6151
R1128 B.n676 B.n675 10.6151
R1129 B.n675 B.n674 10.6151
R1130 B.n674 B.n10 10.6151
R1131 B.n668 B.n10 10.6151
R1132 B.n668 B.n667 10.6151
R1133 B.n667 B.n666 10.6151
R1134 B.n666 B.n17 10.6151
R1135 B.n660 B.n17 10.6151
R1136 B.n660 B.n659 10.6151
R1137 B.n659 B.n658 10.6151
R1138 B.n658 B.n24 10.6151
R1139 B.n652 B.n24 10.6151
R1140 B.n652 B.n651 10.6151
R1141 B.n651 B.n650 10.6151
R1142 B.n650 B.n30 10.6151
R1143 B.n644 B.n30 10.6151
R1144 B.n644 B.n643 10.6151
R1145 B.n643 B.n642 10.6151
R1146 B.n642 B.n38 10.6151
R1147 B.n176 B.n175 6.5566
R1148 B.n192 B.n90 6.5566
R1149 B.n459 B.n361 6.5566
R1150 B.n443 B.n442 6.5566
R1151 B.n283 B.t1 5.20606
R1152 B.t0 B.n671 5.20606
R1153 B.n175 B.n174 4.05904
R1154 B.n195 B.n90 4.05904
R1155 B.n462 B.n361 4.05904
R1156 B.n442 B.n441 4.05904
R1157 B.n682 B.n0 2.81026
R1158 B.n682 B.n1 2.81026
R1159 VP.n0 VP.t1 248.899
R1160 VP.n0 VP.t0 206.379
R1161 VP VP.n0 0.241678
R1162 VDD1 VDD1.t1 106.028
R1163 VDD1 VDD1.t0 68.0318
C0 VN VP 5.05806f
C1 VP VTAIL 2.20186f
C2 VDD1 VP 2.71026f
C3 VN VTAIL 2.18751f
C4 VN VDD1 0.147801f
C5 VDD2 VP 0.303684f
C6 VDD1 VTAIL 4.91582f
C7 VDD2 VN 2.55727f
C8 VDD2 VTAIL 4.96092f
C9 VDD2 VDD1 0.591683f
C10 VDD2 B 4.119998f
C11 VDD1 B 7.05448f
C12 VTAIL B 6.868188f
C13 VN B 9.98105f
C14 VP B 5.502343f
C15 VDD1.t0 B 2.12201f
C16 VDD1.t1 B 2.62745f
C17 VP.t1 B 2.9821f
C18 VP.t0 B 2.56965f
C19 VP.n0 B 4.38755f
C20 VDD2.t1 B 2.62279f
C21 VDD2.t0 B 2.14108f
C22 VDD2.n0 B 2.73678f
C23 VTAIL.t3 B 2.09046f
C24 VTAIL.n0 B 1.52032f
C25 VTAIL.t1 B 2.09046f
C26 VTAIL.n1 B 1.54837f
C27 VTAIL.t0 B 2.09045f
C28 VTAIL.n2 B 1.42073f
C29 VTAIL.t2 B 2.09046f
C30 VTAIL.n3 B 1.35375f
C31 VN.t0 B 2.53143f
C32 VN.t1 B 2.94111f
.ends

