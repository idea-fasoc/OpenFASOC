* NGSPICE file created from diff_pair_sample_0362.ext - technology: sky130A

.subckt diff_pair_sample_0362 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=7.3164 ps=38.3 w=18.76 l=2.46
X1 B.t11 B.t9 B.t10 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=2.46
X2 VDD2.t0 VN.t1 VTAIL.t2 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=7.3164 ps=38.3 w=18.76 l=2.46
X3 VDD1.t1 VP.t0 VTAIL.t1 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=7.3164 ps=38.3 w=18.76 l=2.46
X4 VDD1.t0 VP.t1 VTAIL.t0 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=7.3164 ps=38.3 w=18.76 l=2.46
X5 B.t8 B.t6 B.t7 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=2.46
X6 B.t5 B.t3 B.t4 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=2.46
X7 B.t2 B.t0 B.t1 w_n2086_n4720# sky130_fd_pr__pfet_01v8 ad=7.3164 pd=38.3 as=0 ps=0 w=18.76 l=2.46
R0 VN VN.t1 282.416
R1 VN VN.t0 233.25
R2 VTAIL.n414 VTAIL.n413 756.745
R3 VTAIL.n102 VTAIL.n101 756.745
R4 VTAIL.n310 VTAIL.n309 756.745
R5 VTAIL.n206 VTAIL.n205 756.745
R6 VTAIL.n347 VTAIL.n346 585
R7 VTAIL.n349 VTAIL.n348 585
R8 VTAIL.n342 VTAIL.n341 585
R9 VTAIL.n355 VTAIL.n354 585
R10 VTAIL.n357 VTAIL.n356 585
R11 VTAIL.n338 VTAIL.n337 585
R12 VTAIL.n364 VTAIL.n363 585
R13 VTAIL.n365 VTAIL.n336 585
R14 VTAIL.n367 VTAIL.n366 585
R15 VTAIL.n334 VTAIL.n333 585
R16 VTAIL.n373 VTAIL.n372 585
R17 VTAIL.n375 VTAIL.n374 585
R18 VTAIL.n330 VTAIL.n329 585
R19 VTAIL.n381 VTAIL.n380 585
R20 VTAIL.n383 VTAIL.n382 585
R21 VTAIL.n326 VTAIL.n325 585
R22 VTAIL.n389 VTAIL.n388 585
R23 VTAIL.n391 VTAIL.n390 585
R24 VTAIL.n322 VTAIL.n321 585
R25 VTAIL.n397 VTAIL.n396 585
R26 VTAIL.n399 VTAIL.n398 585
R27 VTAIL.n318 VTAIL.n317 585
R28 VTAIL.n405 VTAIL.n404 585
R29 VTAIL.n407 VTAIL.n406 585
R30 VTAIL.n314 VTAIL.n313 585
R31 VTAIL.n413 VTAIL.n412 585
R32 VTAIL.n35 VTAIL.n34 585
R33 VTAIL.n37 VTAIL.n36 585
R34 VTAIL.n30 VTAIL.n29 585
R35 VTAIL.n43 VTAIL.n42 585
R36 VTAIL.n45 VTAIL.n44 585
R37 VTAIL.n26 VTAIL.n25 585
R38 VTAIL.n52 VTAIL.n51 585
R39 VTAIL.n53 VTAIL.n24 585
R40 VTAIL.n55 VTAIL.n54 585
R41 VTAIL.n22 VTAIL.n21 585
R42 VTAIL.n61 VTAIL.n60 585
R43 VTAIL.n63 VTAIL.n62 585
R44 VTAIL.n18 VTAIL.n17 585
R45 VTAIL.n69 VTAIL.n68 585
R46 VTAIL.n71 VTAIL.n70 585
R47 VTAIL.n14 VTAIL.n13 585
R48 VTAIL.n77 VTAIL.n76 585
R49 VTAIL.n79 VTAIL.n78 585
R50 VTAIL.n10 VTAIL.n9 585
R51 VTAIL.n85 VTAIL.n84 585
R52 VTAIL.n87 VTAIL.n86 585
R53 VTAIL.n6 VTAIL.n5 585
R54 VTAIL.n93 VTAIL.n92 585
R55 VTAIL.n95 VTAIL.n94 585
R56 VTAIL.n2 VTAIL.n1 585
R57 VTAIL.n101 VTAIL.n100 585
R58 VTAIL.n309 VTAIL.n308 585
R59 VTAIL.n210 VTAIL.n209 585
R60 VTAIL.n303 VTAIL.n302 585
R61 VTAIL.n301 VTAIL.n300 585
R62 VTAIL.n214 VTAIL.n213 585
R63 VTAIL.n295 VTAIL.n294 585
R64 VTAIL.n293 VTAIL.n292 585
R65 VTAIL.n218 VTAIL.n217 585
R66 VTAIL.n287 VTAIL.n286 585
R67 VTAIL.n285 VTAIL.n284 585
R68 VTAIL.n222 VTAIL.n221 585
R69 VTAIL.n279 VTAIL.n278 585
R70 VTAIL.n277 VTAIL.n276 585
R71 VTAIL.n226 VTAIL.n225 585
R72 VTAIL.n271 VTAIL.n270 585
R73 VTAIL.n269 VTAIL.n268 585
R74 VTAIL.n230 VTAIL.n229 585
R75 VTAIL.n234 VTAIL.n232 585
R76 VTAIL.n263 VTAIL.n262 585
R77 VTAIL.n261 VTAIL.n260 585
R78 VTAIL.n236 VTAIL.n235 585
R79 VTAIL.n255 VTAIL.n254 585
R80 VTAIL.n253 VTAIL.n252 585
R81 VTAIL.n240 VTAIL.n239 585
R82 VTAIL.n247 VTAIL.n246 585
R83 VTAIL.n245 VTAIL.n244 585
R84 VTAIL.n205 VTAIL.n204 585
R85 VTAIL.n106 VTAIL.n105 585
R86 VTAIL.n199 VTAIL.n198 585
R87 VTAIL.n197 VTAIL.n196 585
R88 VTAIL.n110 VTAIL.n109 585
R89 VTAIL.n191 VTAIL.n190 585
R90 VTAIL.n189 VTAIL.n188 585
R91 VTAIL.n114 VTAIL.n113 585
R92 VTAIL.n183 VTAIL.n182 585
R93 VTAIL.n181 VTAIL.n180 585
R94 VTAIL.n118 VTAIL.n117 585
R95 VTAIL.n175 VTAIL.n174 585
R96 VTAIL.n173 VTAIL.n172 585
R97 VTAIL.n122 VTAIL.n121 585
R98 VTAIL.n167 VTAIL.n166 585
R99 VTAIL.n165 VTAIL.n164 585
R100 VTAIL.n126 VTAIL.n125 585
R101 VTAIL.n130 VTAIL.n128 585
R102 VTAIL.n159 VTAIL.n158 585
R103 VTAIL.n157 VTAIL.n156 585
R104 VTAIL.n132 VTAIL.n131 585
R105 VTAIL.n151 VTAIL.n150 585
R106 VTAIL.n149 VTAIL.n148 585
R107 VTAIL.n136 VTAIL.n135 585
R108 VTAIL.n143 VTAIL.n142 585
R109 VTAIL.n141 VTAIL.n140 585
R110 VTAIL.n345 VTAIL.t3 329.036
R111 VTAIL.n33 VTAIL.t0 329.036
R112 VTAIL.n243 VTAIL.t1 329.036
R113 VTAIL.n139 VTAIL.t2 329.036
R114 VTAIL.n348 VTAIL.n347 171.744
R115 VTAIL.n348 VTAIL.n341 171.744
R116 VTAIL.n355 VTAIL.n341 171.744
R117 VTAIL.n356 VTAIL.n355 171.744
R118 VTAIL.n356 VTAIL.n337 171.744
R119 VTAIL.n364 VTAIL.n337 171.744
R120 VTAIL.n365 VTAIL.n364 171.744
R121 VTAIL.n366 VTAIL.n365 171.744
R122 VTAIL.n366 VTAIL.n333 171.744
R123 VTAIL.n373 VTAIL.n333 171.744
R124 VTAIL.n374 VTAIL.n373 171.744
R125 VTAIL.n374 VTAIL.n329 171.744
R126 VTAIL.n381 VTAIL.n329 171.744
R127 VTAIL.n382 VTAIL.n381 171.744
R128 VTAIL.n382 VTAIL.n325 171.744
R129 VTAIL.n389 VTAIL.n325 171.744
R130 VTAIL.n390 VTAIL.n389 171.744
R131 VTAIL.n390 VTAIL.n321 171.744
R132 VTAIL.n397 VTAIL.n321 171.744
R133 VTAIL.n398 VTAIL.n397 171.744
R134 VTAIL.n398 VTAIL.n317 171.744
R135 VTAIL.n405 VTAIL.n317 171.744
R136 VTAIL.n406 VTAIL.n405 171.744
R137 VTAIL.n406 VTAIL.n313 171.744
R138 VTAIL.n413 VTAIL.n313 171.744
R139 VTAIL.n36 VTAIL.n35 171.744
R140 VTAIL.n36 VTAIL.n29 171.744
R141 VTAIL.n43 VTAIL.n29 171.744
R142 VTAIL.n44 VTAIL.n43 171.744
R143 VTAIL.n44 VTAIL.n25 171.744
R144 VTAIL.n52 VTAIL.n25 171.744
R145 VTAIL.n53 VTAIL.n52 171.744
R146 VTAIL.n54 VTAIL.n53 171.744
R147 VTAIL.n54 VTAIL.n21 171.744
R148 VTAIL.n61 VTAIL.n21 171.744
R149 VTAIL.n62 VTAIL.n61 171.744
R150 VTAIL.n62 VTAIL.n17 171.744
R151 VTAIL.n69 VTAIL.n17 171.744
R152 VTAIL.n70 VTAIL.n69 171.744
R153 VTAIL.n70 VTAIL.n13 171.744
R154 VTAIL.n77 VTAIL.n13 171.744
R155 VTAIL.n78 VTAIL.n77 171.744
R156 VTAIL.n78 VTAIL.n9 171.744
R157 VTAIL.n85 VTAIL.n9 171.744
R158 VTAIL.n86 VTAIL.n85 171.744
R159 VTAIL.n86 VTAIL.n5 171.744
R160 VTAIL.n93 VTAIL.n5 171.744
R161 VTAIL.n94 VTAIL.n93 171.744
R162 VTAIL.n94 VTAIL.n1 171.744
R163 VTAIL.n101 VTAIL.n1 171.744
R164 VTAIL.n309 VTAIL.n209 171.744
R165 VTAIL.n302 VTAIL.n209 171.744
R166 VTAIL.n302 VTAIL.n301 171.744
R167 VTAIL.n301 VTAIL.n213 171.744
R168 VTAIL.n294 VTAIL.n213 171.744
R169 VTAIL.n294 VTAIL.n293 171.744
R170 VTAIL.n293 VTAIL.n217 171.744
R171 VTAIL.n286 VTAIL.n217 171.744
R172 VTAIL.n286 VTAIL.n285 171.744
R173 VTAIL.n285 VTAIL.n221 171.744
R174 VTAIL.n278 VTAIL.n221 171.744
R175 VTAIL.n278 VTAIL.n277 171.744
R176 VTAIL.n277 VTAIL.n225 171.744
R177 VTAIL.n270 VTAIL.n225 171.744
R178 VTAIL.n270 VTAIL.n269 171.744
R179 VTAIL.n269 VTAIL.n229 171.744
R180 VTAIL.n234 VTAIL.n229 171.744
R181 VTAIL.n262 VTAIL.n234 171.744
R182 VTAIL.n262 VTAIL.n261 171.744
R183 VTAIL.n261 VTAIL.n235 171.744
R184 VTAIL.n254 VTAIL.n235 171.744
R185 VTAIL.n254 VTAIL.n253 171.744
R186 VTAIL.n253 VTAIL.n239 171.744
R187 VTAIL.n246 VTAIL.n239 171.744
R188 VTAIL.n246 VTAIL.n245 171.744
R189 VTAIL.n205 VTAIL.n105 171.744
R190 VTAIL.n198 VTAIL.n105 171.744
R191 VTAIL.n198 VTAIL.n197 171.744
R192 VTAIL.n197 VTAIL.n109 171.744
R193 VTAIL.n190 VTAIL.n109 171.744
R194 VTAIL.n190 VTAIL.n189 171.744
R195 VTAIL.n189 VTAIL.n113 171.744
R196 VTAIL.n182 VTAIL.n113 171.744
R197 VTAIL.n182 VTAIL.n181 171.744
R198 VTAIL.n181 VTAIL.n117 171.744
R199 VTAIL.n174 VTAIL.n117 171.744
R200 VTAIL.n174 VTAIL.n173 171.744
R201 VTAIL.n173 VTAIL.n121 171.744
R202 VTAIL.n166 VTAIL.n121 171.744
R203 VTAIL.n166 VTAIL.n165 171.744
R204 VTAIL.n165 VTAIL.n125 171.744
R205 VTAIL.n130 VTAIL.n125 171.744
R206 VTAIL.n158 VTAIL.n130 171.744
R207 VTAIL.n158 VTAIL.n157 171.744
R208 VTAIL.n157 VTAIL.n131 171.744
R209 VTAIL.n150 VTAIL.n131 171.744
R210 VTAIL.n150 VTAIL.n149 171.744
R211 VTAIL.n149 VTAIL.n135 171.744
R212 VTAIL.n142 VTAIL.n135 171.744
R213 VTAIL.n142 VTAIL.n141 171.744
R214 VTAIL.n347 VTAIL.t3 85.8723
R215 VTAIL.n35 VTAIL.t0 85.8723
R216 VTAIL.n245 VTAIL.t1 85.8723
R217 VTAIL.n141 VTAIL.t2 85.8723
R218 VTAIL.n415 VTAIL.n414 34.9005
R219 VTAIL.n103 VTAIL.n102 34.9005
R220 VTAIL.n311 VTAIL.n310 34.9005
R221 VTAIL.n207 VTAIL.n206 34.9005
R222 VTAIL.n207 VTAIL.n103 33.3496
R223 VTAIL.n415 VTAIL.n311 30.9445
R224 VTAIL.n367 VTAIL.n334 13.1884
R225 VTAIL.n55 VTAIL.n22 13.1884
R226 VTAIL.n232 VTAIL.n230 13.1884
R227 VTAIL.n128 VTAIL.n126 13.1884
R228 VTAIL.n368 VTAIL.n336 12.8005
R229 VTAIL.n372 VTAIL.n371 12.8005
R230 VTAIL.n412 VTAIL.n312 12.8005
R231 VTAIL.n56 VTAIL.n24 12.8005
R232 VTAIL.n60 VTAIL.n59 12.8005
R233 VTAIL.n100 VTAIL.n0 12.8005
R234 VTAIL.n308 VTAIL.n208 12.8005
R235 VTAIL.n268 VTAIL.n267 12.8005
R236 VTAIL.n264 VTAIL.n263 12.8005
R237 VTAIL.n204 VTAIL.n104 12.8005
R238 VTAIL.n164 VTAIL.n163 12.8005
R239 VTAIL.n160 VTAIL.n159 12.8005
R240 VTAIL.n363 VTAIL.n362 12.0247
R241 VTAIL.n375 VTAIL.n332 12.0247
R242 VTAIL.n411 VTAIL.n314 12.0247
R243 VTAIL.n51 VTAIL.n50 12.0247
R244 VTAIL.n63 VTAIL.n20 12.0247
R245 VTAIL.n99 VTAIL.n2 12.0247
R246 VTAIL.n307 VTAIL.n210 12.0247
R247 VTAIL.n271 VTAIL.n228 12.0247
R248 VTAIL.n260 VTAIL.n233 12.0247
R249 VTAIL.n203 VTAIL.n106 12.0247
R250 VTAIL.n167 VTAIL.n124 12.0247
R251 VTAIL.n156 VTAIL.n129 12.0247
R252 VTAIL.n361 VTAIL.n338 11.249
R253 VTAIL.n376 VTAIL.n330 11.249
R254 VTAIL.n408 VTAIL.n407 11.249
R255 VTAIL.n49 VTAIL.n26 11.249
R256 VTAIL.n64 VTAIL.n18 11.249
R257 VTAIL.n96 VTAIL.n95 11.249
R258 VTAIL.n304 VTAIL.n303 11.249
R259 VTAIL.n272 VTAIL.n226 11.249
R260 VTAIL.n259 VTAIL.n236 11.249
R261 VTAIL.n200 VTAIL.n199 11.249
R262 VTAIL.n168 VTAIL.n122 11.249
R263 VTAIL.n155 VTAIL.n132 11.249
R264 VTAIL.n346 VTAIL.n345 10.7239
R265 VTAIL.n34 VTAIL.n33 10.7239
R266 VTAIL.n244 VTAIL.n243 10.7239
R267 VTAIL.n140 VTAIL.n139 10.7239
R268 VTAIL.n358 VTAIL.n357 10.4732
R269 VTAIL.n380 VTAIL.n379 10.4732
R270 VTAIL.n404 VTAIL.n316 10.4732
R271 VTAIL.n46 VTAIL.n45 10.4732
R272 VTAIL.n68 VTAIL.n67 10.4732
R273 VTAIL.n92 VTAIL.n4 10.4732
R274 VTAIL.n300 VTAIL.n212 10.4732
R275 VTAIL.n276 VTAIL.n275 10.4732
R276 VTAIL.n256 VTAIL.n255 10.4732
R277 VTAIL.n196 VTAIL.n108 10.4732
R278 VTAIL.n172 VTAIL.n171 10.4732
R279 VTAIL.n152 VTAIL.n151 10.4732
R280 VTAIL.n354 VTAIL.n340 9.69747
R281 VTAIL.n383 VTAIL.n328 9.69747
R282 VTAIL.n403 VTAIL.n318 9.69747
R283 VTAIL.n42 VTAIL.n28 9.69747
R284 VTAIL.n71 VTAIL.n16 9.69747
R285 VTAIL.n91 VTAIL.n6 9.69747
R286 VTAIL.n299 VTAIL.n214 9.69747
R287 VTAIL.n279 VTAIL.n224 9.69747
R288 VTAIL.n252 VTAIL.n238 9.69747
R289 VTAIL.n195 VTAIL.n110 9.69747
R290 VTAIL.n175 VTAIL.n120 9.69747
R291 VTAIL.n148 VTAIL.n134 9.69747
R292 VTAIL.n410 VTAIL.n312 9.45567
R293 VTAIL.n98 VTAIL.n0 9.45567
R294 VTAIL.n306 VTAIL.n208 9.45567
R295 VTAIL.n202 VTAIL.n104 9.45567
R296 VTAIL.n393 VTAIL.n392 9.3005
R297 VTAIL.n395 VTAIL.n394 9.3005
R298 VTAIL.n320 VTAIL.n319 9.3005
R299 VTAIL.n401 VTAIL.n400 9.3005
R300 VTAIL.n403 VTAIL.n402 9.3005
R301 VTAIL.n316 VTAIL.n315 9.3005
R302 VTAIL.n409 VTAIL.n408 9.3005
R303 VTAIL.n411 VTAIL.n410 9.3005
R304 VTAIL.n387 VTAIL.n386 9.3005
R305 VTAIL.n385 VTAIL.n384 9.3005
R306 VTAIL.n328 VTAIL.n327 9.3005
R307 VTAIL.n379 VTAIL.n378 9.3005
R308 VTAIL.n377 VTAIL.n376 9.3005
R309 VTAIL.n332 VTAIL.n331 9.3005
R310 VTAIL.n371 VTAIL.n370 9.3005
R311 VTAIL.n344 VTAIL.n343 9.3005
R312 VTAIL.n351 VTAIL.n350 9.3005
R313 VTAIL.n353 VTAIL.n352 9.3005
R314 VTAIL.n340 VTAIL.n339 9.3005
R315 VTAIL.n359 VTAIL.n358 9.3005
R316 VTAIL.n361 VTAIL.n360 9.3005
R317 VTAIL.n362 VTAIL.n335 9.3005
R318 VTAIL.n369 VTAIL.n368 9.3005
R319 VTAIL.n324 VTAIL.n323 9.3005
R320 VTAIL.n81 VTAIL.n80 9.3005
R321 VTAIL.n83 VTAIL.n82 9.3005
R322 VTAIL.n8 VTAIL.n7 9.3005
R323 VTAIL.n89 VTAIL.n88 9.3005
R324 VTAIL.n91 VTAIL.n90 9.3005
R325 VTAIL.n4 VTAIL.n3 9.3005
R326 VTAIL.n97 VTAIL.n96 9.3005
R327 VTAIL.n99 VTAIL.n98 9.3005
R328 VTAIL.n75 VTAIL.n74 9.3005
R329 VTAIL.n73 VTAIL.n72 9.3005
R330 VTAIL.n16 VTAIL.n15 9.3005
R331 VTAIL.n67 VTAIL.n66 9.3005
R332 VTAIL.n65 VTAIL.n64 9.3005
R333 VTAIL.n20 VTAIL.n19 9.3005
R334 VTAIL.n59 VTAIL.n58 9.3005
R335 VTAIL.n32 VTAIL.n31 9.3005
R336 VTAIL.n39 VTAIL.n38 9.3005
R337 VTAIL.n41 VTAIL.n40 9.3005
R338 VTAIL.n28 VTAIL.n27 9.3005
R339 VTAIL.n47 VTAIL.n46 9.3005
R340 VTAIL.n49 VTAIL.n48 9.3005
R341 VTAIL.n50 VTAIL.n23 9.3005
R342 VTAIL.n57 VTAIL.n56 9.3005
R343 VTAIL.n12 VTAIL.n11 9.3005
R344 VTAIL.n307 VTAIL.n306 9.3005
R345 VTAIL.n305 VTAIL.n304 9.3005
R346 VTAIL.n212 VTAIL.n211 9.3005
R347 VTAIL.n299 VTAIL.n298 9.3005
R348 VTAIL.n297 VTAIL.n296 9.3005
R349 VTAIL.n216 VTAIL.n215 9.3005
R350 VTAIL.n291 VTAIL.n290 9.3005
R351 VTAIL.n289 VTAIL.n288 9.3005
R352 VTAIL.n220 VTAIL.n219 9.3005
R353 VTAIL.n283 VTAIL.n282 9.3005
R354 VTAIL.n281 VTAIL.n280 9.3005
R355 VTAIL.n224 VTAIL.n223 9.3005
R356 VTAIL.n275 VTAIL.n274 9.3005
R357 VTAIL.n273 VTAIL.n272 9.3005
R358 VTAIL.n228 VTAIL.n227 9.3005
R359 VTAIL.n267 VTAIL.n266 9.3005
R360 VTAIL.n265 VTAIL.n264 9.3005
R361 VTAIL.n233 VTAIL.n231 9.3005
R362 VTAIL.n259 VTAIL.n258 9.3005
R363 VTAIL.n257 VTAIL.n256 9.3005
R364 VTAIL.n238 VTAIL.n237 9.3005
R365 VTAIL.n251 VTAIL.n250 9.3005
R366 VTAIL.n249 VTAIL.n248 9.3005
R367 VTAIL.n242 VTAIL.n241 9.3005
R368 VTAIL.n138 VTAIL.n137 9.3005
R369 VTAIL.n145 VTAIL.n144 9.3005
R370 VTAIL.n147 VTAIL.n146 9.3005
R371 VTAIL.n134 VTAIL.n133 9.3005
R372 VTAIL.n153 VTAIL.n152 9.3005
R373 VTAIL.n155 VTAIL.n154 9.3005
R374 VTAIL.n129 VTAIL.n127 9.3005
R375 VTAIL.n161 VTAIL.n160 9.3005
R376 VTAIL.n187 VTAIL.n186 9.3005
R377 VTAIL.n112 VTAIL.n111 9.3005
R378 VTAIL.n193 VTAIL.n192 9.3005
R379 VTAIL.n195 VTAIL.n194 9.3005
R380 VTAIL.n108 VTAIL.n107 9.3005
R381 VTAIL.n201 VTAIL.n200 9.3005
R382 VTAIL.n203 VTAIL.n202 9.3005
R383 VTAIL.n185 VTAIL.n184 9.3005
R384 VTAIL.n116 VTAIL.n115 9.3005
R385 VTAIL.n179 VTAIL.n178 9.3005
R386 VTAIL.n177 VTAIL.n176 9.3005
R387 VTAIL.n120 VTAIL.n119 9.3005
R388 VTAIL.n171 VTAIL.n170 9.3005
R389 VTAIL.n169 VTAIL.n168 9.3005
R390 VTAIL.n124 VTAIL.n123 9.3005
R391 VTAIL.n163 VTAIL.n162 9.3005
R392 VTAIL.n353 VTAIL.n342 8.92171
R393 VTAIL.n384 VTAIL.n326 8.92171
R394 VTAIL.n400 VTAIL.n399 8.92171
R395 VTAIL.n41 VTAIL.n30 8.92171
R396 VTAIL.n72 VTAIL.n14 8.92171
R397 VTAIL.n88 VTAIL.n87 8.92171
R398 VTAIL.n296 VTAIL.n295 8.92171
R399 VTAIL.n280 VTAIL.n222 8.92171
R400 VTAIL.n251 VTAIL.n240 8.92171
R401 VTAIL.n192 VTAIL.n191 8.92171
R402 VTAIL.n176 VTAIL.n118 8.92171
R403 VTAIL.n147 VTAIL.n136 8.92171
R404 VTAIL.n350 VTAIL.n349 8.14595
R405 VTAIL.n388 VTAIL.n387 8.14595
R406 VTAIL.n396 VTAIL.n320 8.14595
R407 VTAIL.n38 VTAIL.n37 8.14595
R408 VTAIL.n76 VTAIL.n75 8.14595
R409 VTAIL.n84 VTAIL.n8 8.14595
R410 VTAIL.n292 VTAIL.n216 8.14595
R411 VTAIL.n284 VTAIL.n283 8.14595
R412 VTAIL.n248 VTAIL.n247 8.14595
R413 VTAIL.n188 VTAIL.n112 8.14595
R414 VTAIL.n180 VTAIL.n179 8.14595
R415 VTAIL.n144 VTAIL.n143 8.14595
R416 VTAIL.n346 VTAIL.n344 7.3702
R417 VTAIL.n391 VTAIL.n324 7.3702
R418 VTAIL.n395 VTAIL.n322 7.3702
R419 VTAIL.n34 VTAIL.n32 7.3702
R420 VTAIL.n79 VTAIL.n12 7.3702
R421 VTAIL.n83 VTAIL.n10 7.3702
R422 VTAIL.n291 VTAIL.n218 7.3702
R423 VTAIL.n287 VTAIL.n220 7.3702
R424 VTAIL.n244 VTAIL.n242 7.3702
R425 VTAIL.n187 VTAIL.n114 7.3702
R426 VTAIL.n183 VTAIL.n116 7.3702
R427 VTAIL.n140 VTAIL.n138 7.3702
R428 VTAIL.n392 VTAIL.n391 6.59444
R429 VTAIL.n392 VTAIL.n322 6.59444
R430 VTAIL.n80 VTAIL.n79 6.59444
R431 VTAIL.n80 VTAIL.n10 6.59444
R432 VTAIL.n288 VTAIL.n218 6.59444
R433 VTAIL.n288 VTAIL.n287 6.59444
R434 VTAIL.n184 VTAIL.n114 6.59444
R435 VTAIL.n184 VTAIL.n183 6.59444
R436 VTAIL.n349 VTAIL.n344 5.81868
R437 VTAIL.n388 VTAIL.n324 5.81868
R438 VTAIL.n396 VTAIL.n395 5.81868
R439 VTAIL.n37 VTAIL.n32 5.81868
R440 VTAIL.n76 VTAIL.n12 5.81868
R441 VTAIL.n84 VTAIL.n83 5.81868
R442 VTAIL.n292 VTAIL.n291 5.81868
R443 VTAIL.n284 VTAIL.n220 5.81868
R444 VTAIL.n247 VTAIL.n242 5.81868
R445 VTAIL.n188 VTAIL.n187 5.81868
R446 VTAIL.n180 VTAIL.n116 5.81868
R447 VTAIL.n143 VTAIL.n138 5.81868
R448 VTAIL.n350 VTAIL.n342 5.04292
R449 VTAIL.n387 VTAIL.n326 5.04292
R450 VTAIL.n399 VTAIL.n320 5.04292
R451 VTAIL.n38 VTAIL.n30 5.04292
R452 VTAIL.n75 VTAIL.n14 5.04292
R453 VTAIL.n87 VTAIL.n8 5.04292
R454 VTAIL.n295 VTAIL.n216 5.04292
R455 VTAIL.n283 VTAIL.n222 5.04292
R456 VTAIL.n248 VTAIL.n240 5.04292
R457 VTAIL.n191 VTAIL.n112 5.04292
R458 VTAIL.n179 VTAIL.n118 5.04292
R459 VTAIL.n144 VTAIL.n136 5.04292
R460 VTAIL.n354 VTAIL.n353 4.26717
R461 VTAIL.n384 VTAIL.n383 4.26717
R462 VTAIL.n400 VTAIL.n318 4.26717
R463 VTAIL.n42 VTAIL.n41 4.26717
R464 VTAIL.n72 VTAIL.n71 4.26717
R465 VTAIL.n88 VTAIL.n6 4.26717
R466 VTAIL.n296 VTAIL.n214 4.26717
R467 VTAIL.n280 VTAIL.n279 4.26717
R468 VTAIL.n252 VTAIL.n251 4.26717
R469 VTAIL.n192 VTAIL.n110 4.26717
R470 VTAIL.n176 VTAIL.n175 4.26717
R471 VTAIL.n148 VTAIL.n147 4.26717
R472 VTAIL.n357 VTAIL.n340 3.49141
R473 VTAIL.n380 VTAIL.n328 3.49141
R474 VTAIL.n404 VTAIL.n403 3.49141
R475 VTAIL.n45 VTAIL.n28 3.49141
R476 VTAIL.n68 VTAIL.n16 3.49141
R477 VTAIL.n92 VTAIL.n91 3.49141
R478 VTAIL.n300 VTAIL.n299 3.49141
R479 VTAIL.n276 VTAIL.n224 3.49141
R480 VTAIL.n255 VTAIL.n238 3.49141
R481 VTAIL.n196 VTAIL.n195 3.49141
R482 VTAIL.n172 VTAIL.n120 3.49141
R483 VTAIL.n151 VTAIL.n134 3.49141
R484 VTAIL.n358 VTAIL.n338 2.71565
R485 VTAIL.n379 VTAIL.n330 2.71565
R486 VTAIL.n407 VTAIL.n316 2.71565
R487 VTAIL.n46 VTAIL.n26 2.71565
R488 VTAIL.n67 VTAIL.n18 2.71565
R489 VTAIL.n95 VTAIL.n4 2.71565
R490 VTAIL.n303 VTAIL.n212 2.71565
R491 VTAIL.n275 VTAIL.n226 2.71565
R492 VTAIL.n256 VTAIL.n236 2.71565
R493 VTAIL.n199 VTAIL.n108 2.71565
R494 VTAIL.n171 VTAIL.n122 2.71565
R495 VTAIL.n152 VTAIL.n132 2.71565
R496 VTAIL.n243 VTAIL.n241 2.41282
R497 VTAIL.n139 VTAIL.n137 2.41282
R498 VTAIL.n345 VTAIL.n343 2.41282
R499 VTAIL.n33 VTAIL.n31 2.41282
R500 VTAIL.n363 VTAIL.n361 1.93989
R501 VTAIL.n376 VTAIL.n375 1.93989
R502 VTAIL.n408 VTAIL.n314 1.93989
R503 VTAIL.n51 VTAIL.n49 1.93989
R504 VTAIL.n64 VTAIL.n63 1.93989
R505 VTAIL.n96 VTAIL.n2 1.93989
R506 VTAIL.n304 VTAIL.n210 1.93989
R507 VTAIL.n272 VTAIL.n271 1.93989
R508 VTAIL.n260 VTAIL.n259 1.93989
R509 VTAIL.n200 VTAIL.n106 1.93989
R510 VTAIL.n168 VTAIL.n167 1.93989
R511 VTAIL.n156 VTAIL.n155 1.93989
R512 VTAIL.n311 VTAIL.n207 1.67291
R513 VTAIL.n362 VTAIL.n336 1.16414
R514 VTAIL.n372 VTAIL.n332 1.16414
R515 VTAIL.n412 VTAIL.n411 1.16414
R516 VTAIL.n50 VTAIL.n24 1.16414
R517 VTAIL.n60 VTAIL.n20 1.16414
R518 VTAIL.n100 VTAIL.n99 1.16414
R519 VTAIL.n308 VTAIL.n307 1.16414
R520 VTAIL.n268 VTAIL.n228 1.16414
R521 VTAIL.n263 VTAIL.n233 1.16414
R522 VTAIL.n204 VTAIL.n203 1.16414
R523 VTAIL.n164 VTAIL.n124 1.16414
R524 VTAIL.n159 VTAIL.n129 1.16414
R525 VTAIL VTAIL.n103 1.12981
R526 VTAIL VTAIL.n415 0.543603
R527 VTAIL.n368 VTAIL.n367 0.388379
R528 VTAIL.n371 VTAIL.n334 0.388379
R529 VTAIL.n414 VTAIL.n312 0.388379
R530 VTAIL.n56 VTAIL.n55 0.388379
R531 VTAIL.n59 VTAIL.n22 0.388379
R532 VTAIL.n102 VTAIL.n0 0.388379
R533 VTAIL.n310 VTAIL.n208 0.388379
R534 VTAIL.n267 VTAIL.n230 0.388379
R535 VTAIL.n264 VTAIL.n232 0.388379
R536 VTAIL.n206 VTAIL.n104 0.388379
R537 VTAIL.n163 VTAIL.n126 0.388379
R538 VTAIL.n160 VTAIL.n128 0.388379
R539 VTAIL.n351 VTAIL.n343 0.155672
R540 VTAIL.n352 VTAIL.n351 0.155672
R541 VTAIL.n352 VTAIL.n339 0.155672
R542 VTAIL.n359 VTAIL.n339 0.155672
R543 VTAIL.n360 VTAIL.n359 0.155672
R544 VTAIL.n360 VTAIL.n335 0.155672
R545 VTAIL.n369 VTAIL.n335 0.155672
R546 VTAIL.n370 VTAIL.n369 0.155672
R547 VTAIL.n370 VTAIL.n331 0.155672
R548 VTAIL.n377 VTAIL.n331 0.155672
R549 VTAIL.n378 VTAIL.n377 0.155672
R550 VTAIL.n378 VTAIL.n327 0.155672
R551 VTAIL.n385 VTAIL.n327 0.155672
R552 VTAIL.n386 VTAIL.n385 0.155672
R553 VTAIL.n386 VTAIL.n323 0.155672
R554 VTAIL.n393 VTAIL.n323 0.155672
R555 VTAIL.n394 VTAIL.n393 0.155672
R556 VTAIL.n394 VTAIL.n319 0.155672
R557 VTAIL.n401 VTAIL.n319 0.155672
R558 VTAIL.n402 VTAIL.n401 0.155672
R559 VTAIL.n402 VTAIL.n315 0.155672
R560 VTAIL.n409 VTAIL.n315 0.155672
R561 VTAIL.n410 VTAIL.n409 0.155672
R562 VTAIL.n39 VTAIL.n31 0.155672
R563 VTAIL.n40 VTAIL.n39 0.155672
R564 VTAIL.n40 VTAIL.n27 0.155672
R565 VTAIL.n47 VTAIL.n27 0.155672
R566 VTAIL.n48 VTAIL.n47 0.155672
R567 VTAIL.n48 VTAIL.n23 0.155672
R568 VTAIL.n57 VTAIL.n23 0.155672
R569 VTAIL.n58 VTAIL.n57 0.155672
R570 VTAIL.n58 VTAIL.n19 0.155672
R571 VTAIL.n65 VTAIL.n19 0.155672
R572 VTAIL.n66 VTAIL.n65 0.155672
R573 VTAIL.n66 VTAIL.n15 0.155672
R574 VTAIL.n73 VTAIL.n15 0.155672
R575 VTAIL.n74 VTAIL.n73 0.155672
R576 VTAIL.n74 VTAIL.n11 0.155672
R577 VTAIL.n81 VTAIL.n11 0.155672
R578 VTAIL.n82 VTAIL.n81 0.155672
R579 VTAIL.n82 VTAIL.n7 0.155672
R580 VTAIL.n89 VTAIL.n7 0.155672
R581 VTAIL.n90 VTAIL.n89 0.155672
R582 VTAIL.n90 VTAIL.n3 0.155672
R583 VTAIL.n97 VTAIL.n3 0.155672
R584 VTAIL.n98 VTAIL.n97 0.155672
R585 VTAIL.n306 VTAIL.n305 0.155672
R586 VTAIL.n305 VTAIL.n211 0.155672
R587 VTAIL.n298 VTAIL.n211 0.155672
R588 VTAIL.n298 VTAIL.n297 0.155672
R589 VTAIL.n297 VTAIL.n215 0.155672
R590 VTAIL.n290 VTAIL.n215 0.155672
R591 VTAIL.n290 VTAIL.n289 0.155672
R592 VTAIL.n289 VTAIL.n219 0.155672
R593 VTAIL.n282 VTAIL.n219 0.155672
R594 VTAIL.n282 VTAIL.n281 0.155672
R595 VTAIL.n281 VTAIL.n223 0.155672
R596 VTAIL.n274 VTAIL.n223 0.155672
R597 VTAIL.n274 VTAIL.n273 0.155672
R598 VTAIL.n273 VTAIL.n227 0.155672
R599 VTAIL.n266 VTAIL.n227 0.155672
R600 VTAIL.n266 VTAIL.n265 0.155672
R601 VTAIL.n265 VTAIL.n231 0.155672
R602 VTAIL.n258 VTAIL.n231 0.155672
R603 VTAIL.n258 VTAIL.n257 0.155672
R604 VTAIL.n257 VTAIL.n237 0.155672
R605 VTAIL.n250 VTAIL.n237 0.155672
R606 VTAIL.n250 VTAIL.n249 0.155672
R607 VTAIL.n249 VTAIL.n241 0.155672
R608 VTAIL.n202 VTAIL.n201 0.155672
R609 VTAIL.n201 VTAIL.n107 0.155672
R610 VTAIL.n194 VTAIL.n107 0.155672
R611 VTAIL.n194 VTAIL.n193 0.155672
R612 VTAIL.n193 VTAIL.n111 0.155672
R613 VTAIL.n186 VTAIL.n111 0.155672
R614 VTAIL.n186 VTAIL.n185 0.155672
R615 VTAIL.n185 VTAIL.n115 0.155672
R616 VTAIL.n178 VTAIL.n115 0.155672
R617 VTAIL.n178 VTAIL.n177 0.155672
R618 VTAIL.n177 VTAIL.n119 0.155672
R619 VTAIL.n170 VTAIL.n119 0.155672
R620 VTAIL.n170 VTAIL.n169 0.155672
R621 VTAIL.n169 VTAIL.n123 0.155672
R622 VTAIL.n162 VTAIL.n123 0.155672
R623 VTAIL.n162 VTAIL.n161 0.155672
R624 VTAIL.n161 VTAIL.n127 0.155672
R625 VTAIL.n154 VTAIL.n127 0.155672
R626 VTAIL.n154 VTAIL.n153 0.155672
R627 VTAIL.n153 VTAIL.n133 0.155672
R628 VTAIL.n146 VTAIL.n133 0.155672
R629 VTAIL.n146 VTAIL.n145 0.155672
R630 VTAIL.n145 VTAIL.n137 0.155672
R631 VDD2.n205 VDD2.n204 756.745
R632 VDD2.n102 VDD2.n101 756.745
R633 VDD2.n204 VDD2.n203 585
R634 VDD2.n105 VDD2.n104 585
R635 VDD2.n198 VDD2.n197 585
R636 VDD2.n196 VDD2.n195 585
R637 VDD2.n109 VDD2.n108 585
R638 VDD2.n190 VDD2.n189 585
R639 VDD2.n188 VDD2.n187 585
R640 VDD2.n113 VDD2.n112 585
R641 VDD2.n182 VDD2.n181 585
R642 VDD2.n180 VDD2.n179 585
R643 VDD2.n117 VDD2.n116 585
R644 VDD2.n174 VDD2.n173 585
R645 VDD2.n172 VDD2.n171 585
R646 VDD2.n121 VDD2.n120 585
R647 VDD2.n166 VDD2.n165 585
R648 VDD2.n164 VDD2.n163 585
R649 VDD2.n125 VDD2.n124 585
R650 VDD2.n129 VDD2.n127 585
R651 VDD2.n158 VDD2.n157 585
R652 VDD2.n156 VDD2.n155 585
R653 VDD2.n131 VDD2.n130 585
R654 VDD2.n150 VDD2.n149 585
R655 VDD2.n148 VDD2.n147 585
R656 VDD2.n135 VDD2.n134 585
R657 VDD2.n142 VDD2.n141 585
R658 VDD2.n140 VDD2.n139 585
R659 VDD2.n35 VDD2.n34 585
R660 VDD2.n37 VDD2.n36 585
R661 VDD2.n30 VDD2.n29 585
R662 VDD2.n43 VDD2.n42 585
R663 VDD2.n45 VDD2.n44 585
R664 VDD2.n26 VDD2.n25 585
R665 VDD2.n52 VDD2.n51 585
R666 VDD2.n53 VDD2.n24 585
R667 VDD2.n55 VDD2.n54 585
R668 VDD2.n22 VDD2.n21 585
R669 VDD2.n61 VDD2.n60 585
R670 VDD2.n63 VDD2.n62 585
R671 VDD2.n18 VDD2.n17 585
R672 VDD2.n69 VDD2.n68 585
R673 VDD2.n71 VDD2.n70 585
R674 VDD2.n14 VDD2.n13 585
R675 VDD2.n77 VDD2.n76 585
R676 VDD2.n79 VDD2.n78 585
R677 VDD2.n10 VDD2.n9 585
R678 VDD2.n85 VDD2.n84 585
R679 VDD2.n87 VDD2.n86 585
R680 VDD2.n6 VDD2.n5 585
R681 VDD2.n93 VDD2.n92 585
R682 VDD2.n95 VDD2.n94 585
R683 VDD2.n2 VDD2.n1 585
R684 VDD2.n101 VDD2.n100 585
R685 VDD2.n138 VDD2.t0 329.036
R686 VDD2.n33 VDD2.t1 329.036
R687 VDD2.n204 VDD2.n104 171.744
R688 VDD2.n197 VDD2.n104 171.744
R689 VDD2.n197 VDD2.n196 171.744
R690 VDD2.n196 VDD2.n108 171.744
R691 VDD2.n189 VDD2.n108 171.744
R692 VDD2.n189 VDD2.n188 171.744
R693 VDD2.n188 VDD2.n112 171.744
R694 VDD2.n181 VDD2.n112 171.744
R695 VDD2.n181 VDD2.n180 171.744
R696 VDD2.n180 VDD2.n116 171.744
R697 VDD2.n173 VDD2.n116 171.744
R698 VDD2.n173 VDD2.n172 171.744
R699 VDD2.n172 VDD2.n120 171.744
R700 VDD2.n165 VDD2.n120 171.744
R701 VDD2.n165 VDD2.n164 171.744
R702 VDD2.n164 VDD2.n124 171.744
R703 VDD2.n129 VDD2.n124 171.744
R704 VDD2.n157 VDD2.n129 171.744
R705 VDD2.n157 VDD2.n156 171.744
R706 VDD2.n156 VDD2.n130 171.744
R707 VDD2.n149 VDD2.n130 171.744
R708 VDD2.n149 VDD2.n148 171.744
R709 VDD2.n148 VDD2.n134 171.744
R710 VDD2.n141 VDD2.n134 171.744
R711 VDD2.n141 VDD2.n140 171.744
R712 VDD2.n36 VDD2.n35 171.744
R713 VDD2.n36 VDD2.n29 171.744
R714 VDD2.n43 VDD2.n29 171.744
R715 VDD2.n44 VDD2.n43 171.744
R716 VDD2.n44 VDD2.n25 171.744
R717 VDD2.n52 VDD2.n25 171.744
R718 VDD2.n53 VDD2.n52 171.744
R719 VDD2.n54 VDD2.n53 171.744
R720 VDD2.n54 VDD2.n21 171.744
R721 VDD2.n61 VDD2.n21 171.744
R722 VDD2.n62 VDD2.n61 171.744
R723 VDD2.n62 VDD2.n17 171.744
R724 VDD2.n69 VDD2.n17 171.744
R725 VDD2.n70 VDD2.n69 171.744
R726 VDD2.n70 VDD2.n13 171.744
R727 VDD2.n77 VDD2.n13 171.744
R728 VDD2.n78 VDD2.n77 171.744
R729 VDD2.n78 VDD2.n9 171.744
R730 VDD2.n85 VDD2.n9 171.744
R731 VDD2.n86 VDD2.n85 171.744
R732 VDD2.n86 VDD2.n5 171.744
R733 VDD2.n93 VDD2.n5 171.744
R734 VDD2.n94 VDD2.n93 171.744
R735 VDD2.n94 VDD2.n1 171.744
R736 VDD2.n101 VDD2.n1 171.744
R737 VDD2.n206 VDD2.n102 96.2215
R738 VDD2.n140 VDD2.t0 85.8723
R739 VDD2.n35 VDD2.t1 85.8723
R740 VDD2.n206 VDD2.n205 51.5793
R741 VDD2.n127 VDD2.n125 13.1884
R742 VDD2.n55 VDD2.n22 13.1884
R743 VDD2.n203 VDD2.n103 12.8005
R744 VDD2.n163 VDD2.n162 12.8005
R745 VDD2.n159 VDD2.n158 12.8005
R746 VDD2.n56 VDD2.n24 12.8005
R747 VDD2.n60 VDD2.n59 12.8005
R748 VDD2.n100 VDD2.n0 12.8005
R749 VDD2.n202 VDD2.n105 12.0247
R750 VDD2.n166 VDD2.n123 12.0247
R751 VDD2.n155 VDD2.n128 12.0247
R752 VDD2.n51 VDD2.n50 12.0247
R753 VDD2.n63 VDD2.n20 12.0247
R754 VDD2.n99 VDD2.n2 12.0247
R755 VDD2.n199 VDD2.n198 11.249
R756 VDD2.n167 VDD2.n121 11.249
R757 VDD2.n154 VDD2.n131 11.249
R758 VDD2.n49 VDD2.n26 11.249
R759 VDD2.n64 VDD2.n18 11.249
R760 VDD2.n96 VDD2.n95 11.249
R761 VDD2.n139 VDD2.n138 10.7239
R762 VDD2.n34 VDD2.n33 10.7239
R763 VDD2.n195 VDD2.n107 10.4732
R764 VDD2.n171 VDD2.n170 10.4732
R765 VDD2.n151 VDD2.n150 10.4732
R766 VDD2.n46 VDD2.n45 10.4732
R767 VDD2.n68 VDD2.n67 10.4732
R768 VDD2.n92 VDD2.n4 10.4732
R769 VDD2.n194 VDD2.n109 9.69747
R770 VDD2.n174 VDD2.n119 9.69747
R771 VDD2.n147 VDD2.n133 9.69747
R772 VDD2.n42 VDD2.n28 9.69747
R773 VDD2.n71 VDD2.n16 9.69747
R774 VDD2.n91 VDD2.n6 9.69747
R775 VDD2.n201 VDD2.n103 9.45567
R776 VDD2.n98 VDD2.n0 9.45567
R777 VDD2.n202 VDD2.n201 9.3005
R778 VDD2.n200 VDD2.n199 9.3005
R779 VDD2.n107 VDD2.n106 9.3005
R780 VDD2.n194 VDD2.n193 9.3005
R781 VDD2.n192 VDD2.n191 9.3005
R782 VDD2.n111 VDD2.n110 9.3005
R783 VDD2.n186 VDD2.n185 9.3005
R784 VDD2.n184 VDD2.n183 9.3005
R785 VDD2.n115 VDD2.n114 9.3005
R786 VDD2.n178 VDD2.n177 9.3005
R787 VDD2.n176 VDD2.n175 9.3005
R788 VDD2.n119 VDD2.n118 9.3005
R789 VDD2.n170 VDD2.n169 9.3005
R790 VDD2.n168 VDD2.n167 9.3005
R791 VDD2.n123 VDD2.n122 9.3005
R792 VDD2.n162 VDD2.n161 9.3005
R793 VDD2.n160 VDD2.n159 9.3005
R794 VDD2.n128 VDD2.n126 9.3005
R795 VDD2.n154 VDD2.n153 9.3005
R796 VDD2.n152 VDD2.n151 9.3005
R797 VDD2.n133 VDD2.n132 9.3005
R798 VDD2.n146 VDD2.n145 9.3005
R799 VDD2.n144 VDD2.n143 9.3005
R800 VDD2.n137 VDD2.n136 9.3005
R801 VDD2.n81 VDD2.n80 9.3005
R802 VDD2.n83 VDD2.n82 9.3005
R803 VDD2.n8 VDD2.n7 9.3005
R804 VDD2.n89 VDD2.n88 9.3005
R805 VDD2.n91 VDD2.n90 9.3005
R806 VDD2.n4 VDD2.n3 9.3005
R807 VDD2.n97 VDD2.n96 9.3005
R808 VDD2.n99 VDD2.n98 9.3005
R809 VDD2.n75 VDD2.n74 9.3005
R810 VDD2.n73 VDD2.n72 9.3005
R811 VDD2.n16 VDD2.n15 9.3005
R812 VDD2.n67 VDD2.n66 9.3005
R813 VDD2.n65 VDD2.n64 9.3005
R814 VDD2.n20 VDD2.n19 9.3005
R815 VDD2.n59 VDD2.n58 9.3005
R816 VDD2.n32 VDD2.n31 9.3005
R817 VDD2.n39 VDD2.n38 9.3005
R818 VDD2.n41 VDD2.n40 9.3005
R819 VDD2.n28 VDD2.n27 9.3005
R820 VDD2.n47 VDD2.n46 9.3005
R821 VDD2.n49 VDD2.n48 9.3005
R822 VDD2.n50 VDD2.n23 9.3005
R823 VDD2.n57 VDD2.n56 9.3005
R824 VDD2.n12 VDD2.n11 9.3005
R825 VDD2.n191 VDD2.n190 8.92171
R826 VDD2.n175 VDD2.n117 8.92171
R827 VDD2.n146 VDD2.n135 8.92171
R828 VDD2.n41 VDD2.n30 8.92171
R829 VDD2.n72 VDD2.n14 8.92171
R830 VDD2.n88 VDD2.n87 8.92171
R831 VDD2.n187 VDD2.n111 8.14595
R832 VDD2.n179 VDD2.n178 8.14595
R833 VDD2.n143 VDD2.n142 8.14595
R834 VDD2.n38 VDD2.n37 8.14595
R835 VDD2.n76 VDD2.n75 8.14595
R836 VDD2.n84 VDD2.n8 8.14595
R837 VDD2.n186 VDD2.n113 7.3702
R838 VDD2.n182 VDD2.n115 7.3702
R839 VDD2.n139 VDD2.n137 7.3702
R840 VDD2.n34 VDD2.n32 7.3702
R841 VDD2.n79 VDD2.n12 7.3702
R842 VDD2.n83 VDD2.n10 7.3702
R843 VDD2.n183 VDD2.n113 6.59444
R844 VDD2.n183 VDD2.n182 6.59444
R845 VDD2.n80 VDD2.n79 6.59444
R846 VDD2.n80 VDD2.n10 6.59444
R847 VDD2.n187 VDD2.n186 5.81868
R848 VDD2.n179 VDD2.n115 5.81868
R849 VDD2.n142 VDD2.n137 5.81868
R850 VDD2.n37 VDD2.n32 5.81868
R851 VDD2.n76 VDD2.n12 5.81868
R852 VDD2.n84 VDD2.n83 5.81868
R853 VDD2.n190 VDD2.n111 5.04292
R854 VDD2.n178 VDD2.n117 5.04292
R855 VDD2.n143 VDD2.n135 5.04292
R856 VDD2.n38 VDD2.n30 5.04292
R857 VDD2.n75 VDD2.n14 5.04292
R858 VDD2.n87 VDD2.n8 5.04292
R859 VDD2.n191 VDD2.n109 4.26717
R860 VDD2.n175 VDD2.n174 4.26717
R861 VDD2.n147 VDD2.n146 4.26717
R862 VDD2.n42 VDD2.n41 4.26717
R863 VDD2.n72 VDD2.n71 4.26717
R864 VDD2.n88 VDD2.n6 4.26717
R865 VDD2.n195 VDD2.n194 3.49141
R866 VDD2.n171 VDD2.n119 3.49141
R867 VDD2.n150 VDD2.n133 3.49141
R868 VDD2.n45 VDD2.n28 3.49141
R869 VDD2.n68 VDD2.n16 3.49141
R870 VDD2.n92 VDD2.n91 3.49141
R871 VDD2.n198 VDD2.n107 2.71565
R872 VDD2.n170 VDD2.n121 2.71565
R873 VDD2.n151 VDD2.n131 2.71565
R874 VDD2.n46 VDD2.n26 2.71565
R875 VDD2.n67 VDD2.n18 2.71565
R876 VDD2.n95 VDD2.n4 2.71565
R877 VDD2.n138 VDD2.n136 2.41282
R878 VDD2.n33 VDD2.n31 2.41282
R879 VDD2.n199 VDD2.n105 1.93989
R880 VDD2.n167 VDD2.n166 1.93989
R881 VDD2.n155 VDD2.n154 1.93989
R882 VDD2.n51 VDD2.n49 1.93989
R883 VDD2.n64 VDD2.n63 1.93989
R884 VDD2.n96 VDD2.n2 1.93989
R885 VDD2.n203 VDD2.n202 1.16414
R886 VDD2.n163 VDD2.n123 1.16414
R887 VDD2.n158 VDD2.n128 1.16414
R888 VDD2.n50 VDD2.n24 1.16414
R889 VDD2.n60 VDD2.n20 1.16414
R890 VDD2.n100 VDD2.n99 1.16414
R891 VDD2 VDD2.n206 0.659983
R892 VDD2.n205 VDD2.n103 0.388379
R893 VDD2.n162 VDD2.n125 0.388379
R894 VDD2.n159 VDD2.n127 0.388379
R895 VDD2.n56 VDD2.n55 0.388379
R896 VDD2.n59 VDD2.n22 0.388379
R897 VDD2.n102 VDD2.n0 0.388379
R898 VDD2.n201 VDD2.n200 0.155672
R899 VDD2.n200 VDD2.n106 0.155672
R900 VDD2.n193 VDD2.n106 0.155672
R901 VDD2.n193 VDD2.n192 0.155672
R902 VDD2.n192 VDD2.n110 0.155672
R903 VDD2.n185 VDD2.n110 0.155672
R904 VDD2.n185 VDD2.n184 0.155672
R905 VDD2.n184 VDD2.n114 0.155672
R906 VDD2.n177 VDD2.n114 0.155672
R907 VDD2.n177 VDD2.n176 0.155672
R908 VDD2.n176 VDD2.n118 0.155672
R909 VDD2.n169 VDD2.n118 0.155672
R910 VDD2.n169 VDD2.n168 0.155672
R911 VDD2.n168 VDD2.n122 0.155672
R912 VDD2.n161 VDD2.n122 0.155672
R913 VDD2.n161 VDD2.n160 0.155672
R914 VDD2.n160 VDD2.n126 0.155672
R915 VDD2.n153 VDD2.n126 0.155672
R916 VDD2.n153 VDD2.n152 0.155672
R917 VDD2.n152 VDD2.n132 0.155672
R918 VDD2.n145 VDD2.n132 0.155672
R919 VDD2.n145 VDD2.n144 0.155672
R920 VDD2.n144 VDD2.n136 0.155672
R921 VDD2.n39 VDD2.n31 0.155672
R922 VDD2.n40 VDD2.n39 0.155672
R923 VDD2.n40 VDD2.n27 0.155672
R924 VDD2.n47 VDD2.n27 0.155672
R925 VDD2.n48 VDD2.n47 0.155672
R926 VDD2.n48 VDD2.n23 0.155672
R927 VDD2.n57 VDD2.n23 0.155672
R928 VDD2.n58 VDD2.n57 0.155672
R929 VDD2.n58 VDD2.n19 0.155672
R930 VDD2.n65 VDD2.n19 0.155672
R931 VDD2.n66 VDD2.n65 0.155672
R932 VDD2.n66 VDD2.n15 0.155672
R933 VDD2.n73 VDD2.n15 0.155672
R934 VDD2.n74 VDD2.n73 0.155672
R935 VDD2.n74 VDD2.n11 0.155672
R936 VDD2.n81 VDD2.n11 0.155672
R937 VDD2.n82 VDD2.n81 0.155672
R938 VDD2.n82 VDD2.n7 0.155672
R939 VDD2.n89 VDD2.n7 0.155672
R940 VDD2.n90 VDD2.n89 0.155672
R941 VDD2.n90 VDD2.n3 0.155672
R942 VDD2.n97 VDD2.n3 0.155672
R943 VDD2.n98 VDD2.n97 0.155672
R944 B.n427 B.n426 585
R945 B.n425 B.n110 585
R946 B.n424 B.n423 585
R947 B.n422 B.n111 585
R948 B.n421 B.n420 585
R949 B.n419 B.n112 585
R950 B.n418 B.n417 585
R951 B.n416 B.n113 585
R952 B.n415 B.n414 585
R953 B.n413 B.n114 585
R954 B.n412 B.n411 585
R955 B.n410 B.n115 585
R956 B.n409 B.n408 585
R957 B.n407 B.n116 585
R958 B.n406 B.n405 585
R959 B.n404 B.n117 585
R960 B.n403 B.n402 585
R961 B.n401 B.n118 585
R962 B.n400 B.n399 585
R963 B.n398 B.n119 585
R964 B.n397 B.n396 585
R965 B.n395 B.n120 585
R966 B.n394 B.n393 585
R967 B.n392 B.n121 585
R968 B.n391 B.n390 585
R969 B.n389 B.n122 585
R970 B.n388 B.n387 585
R971 B.n386 B.n123 585
R972 B.n385 B.n384 585
R973 B.n383 B.n124 585
R974 B.n382 B.n381 585
R975 B.n380 B.n125 585
R976 B.n379 B.n378 585
R977 B.n377 B.n126 585
R978 B.n376 B.n375 585
R979 B.n374 B.n127 585
R980 B.n373 B.n372 585
R981 B.n371 B.n128 585
R982 B.n370 B.n369 585
R983 B.n368 B.n129 585
R984 B.n367 B.n366 585
R985 B.n365 B.n130 585
R986 B.n364 B.n363 585
R987 B.n362 B.n131 585
R988 B.n361 B.n360 585
R989 B.n359 B.n132 585
R990 B.n358 B.n357 585
R991 B.n356 B.n133 585
R992 B.n355 B.n354 585
R993 B.n353 B.n134 585
R994 B.n352 B.n351 585
R995 B.n350 B.n135 585
R996 B.n349 B.n348 585
R997 B.n347 B.n136 585
R998 B.n346 B.n345 585
R999 B.n344 B.n137 585
R1000 B.n343 B.n342 585
R1001 B.n341 B.n138 585
R1002 B.n340 B.n339 585
R1003 B.n338 B.n139 585
R1004 B.n337 B.n336 585
R1005 B.n335 B.n140 585
R1006 B.n334 B.n333 585
R1007 B.n329 B.n141 585
R1008 B.n328 B.n327 585
R1009 B.n326 B.n142 585
R1010 B.n325 B.n324 585
R1011 B.n323 B.n143 585
R1012 B.n322 B.n321 585
R1013 B.n320 B.n144 585
R1014 B.n319 B.n318 585
R1015 B.n316 B.n145 585
R1016 B.n315 B.n314 585
R1017 B.n313 B.n148 585
R1018 B.n312 B.n311 585
R1019 B.n310 B.n149 585
R1020 B.n309 B.n308 585
R1021 B.n307 B.n150 585
R1022 B.n306 B.n305 585
R1023 B.n304 B.n151 585
R1024 B.n303 B.n302 585
R1025 B.n301 B.n152 585
R1026 B.n300 B.n299 585
R1027 B.n298 B.n153 585
R1028 B.n297 B.n296 585
R1029 B.n295 B.n154 585
R1030 B.n294 B.n293 585
R1031 B.n292 B.n155 585
R1032 B.n291 B.n290 585
R1033 B.n289 B.n156 585
R1034 B.n288 B.n287 585
R1035 B.n286 B.n157 585
R1036 B.n285 B.n284 585
R1037 B.n283 B.n158 585
R1038 B.n282 B.n281 585
R1039 B.n280 B.n159 585
R1040 B.n279 B.n278 585
R1041 B.n277 B.n160 585
R1042 B.n276 B.n275 585
R1043 B.n274 B.n161 585
R1044 B.n273 B.n272 585
R1045 B.n271 B.n162 585
R1046 B.n270 B.n269 585
R1047 B.n268 B.n163 585
R1048 B.n267 B.n266 585
R1049 B.n265 B.n164 585
R1050 B.n264 B.n263 585
R1051 B.n262 B.n165 585
R1052 B.n261 B.n260 585
R1053 B.n259 B.n166 585
R1054 B.n258 B.n257 585
R1055 B.n256 B.n167 585
R1056 B.n255 B.n254 585
R1057 B.n253 B.n168 585
R1058 B.n252 B.n251 585
R1059 B.n250 B.n169 585
R1060 B.n249 B.n248 585
R1061 B.n247 B.n170 585
R1062 B.n246 B.n245 585
R1063 B.n244 B.n171 585
R1064 B.n243 B.n242 585
R1065 B.n241 B.n172 585
R1066 B.n240 B.n239 585
R1067 B.n238 B.n173 585
R1068 B.n237 B.n236 585
R1069 B.n235 B.n174 585
R1070 B.n234 B.n233 585
R1071 B.n232 B.n175 585
R1072 B.n231 B.n230 585
R1073 B.n229 B.n176 585
R1074 B.n228 B.n227 585
R1075 B.n226 B.n177 585
R1076 B.n225 B.n224 585
R1077 B.n428 B.n109 585
R1078 B.n430 B.n429 585
R1079 B.n431 B.n108 585
R1080 B.n433 B.n432 585
R1081 B.n434 B.n107 585
R1082 B.n436 B.n435 585
R1083 B.n437 B.n106 585
R1084 B.n439 B.n438 585
R1085 B.n440 B.n105 585
R1086 B.n442 B.n441 585
R1087 B.n443 B.n104 585
R1088 B.n445 B.n444 585
R1089 B.n446 B.n103 585
R1090 B.n448 B.n447 585
R1091 B.n449 B.n102 585
R1092 B.n451 B.n450 585
R1093 B.n452 B.n101 585
R1094 B.n454 B.n453 585
R1095 B.n455 B.n100 585
R1096 B.n457 B.n456 585
R1097 B.n458 B.n99 585
R1098 B.n460 B.n459 585
R1099 B.n461 B.n98 585
R1100 B.n463 B.n462 585
R1101 B.n464 B.n97 585
R1102 B.n466 B.n465 585
R1103 B.n467 B.n96 585
R1104 B.n469 B.n468 585
R1105 B.n470 B.n95 585
R1106 B.n472 B.n471 585
R1107 B.n473 B.n94 585
R1108 B.n475 B.n474 585
R1109 B.n476 B.n93 585
R1110 B.n478 B.n477 585
R1111 B.n479 B.n92 585
R1112 B.n481 B.n480 585
R1113 B.n482 B.n91 585
R1114 B.n484 B.n483 585
R1115 B.n485 B.n90 585
R1116 B.n487 B.n486 585
R1117 B.n488 B.n89 585
R1118 B.n490 B.n489 585
R1119 B.n491 B.n88 585
R1120 B.n493 B.n492 585
R1121 B.n494 B.n87 585
R1122 B.n496 B.n495 585
R1123 B.n497 B.n86 585
R1124 B.n499 B.n498 585
R1125 B.n500 B.n85 585
R1126 B.n502 B.n501 585
R1127 B.n703 B.n14 585
R1128 B.n702 B.n701 585
R1129 B.n700 B.n15 585
R1130 B.n699 B.n698 585
R1131 B.n697 B.n16 585
R1132 B.n696 B.n695 585
R1133 B.n694 B.n17 585
R1134 B.n693 B.n692 585
R1135 B.n691 B.n18 585
R1136 B.n690 B.n689 585
R1137 B.n688 B.n19 585
R1138 B.n687 B.n686 585
R1139 B.n685 B.n20 585
R1140 B.n684 B.n683 585
R1141 B.n682 B.n21 585
R1142 B.n681 B.n680 585
R1143 B.n679 B.n22 585
R1144 B.n678 B.n677 585
R1145 B.n676 B.n23 585
R1146 B.n675 B.n674 585
R1147 B.n673 B.n24 585
R1148 B.n672 B.n671 585
R1149 B.n670 B.n25 585
R1150 B.n669 B.n668 585
R1151 B.n667 B.n26 585
R1152 B.n666 B.n665 585
R1153 B.n664 B.n27 585
R1154 B.n663 B.n662 585
R1155 B.n661 B.n28 585
R1156 B.n660 B.n659 585
R1157 B.n658 B.n29 585
R1158 B.n657 B.n656 585
R1159 B.n655 B.n30 585
R1160 B.n654 B.n653 585
R1161 B.n652 B.n31 585
R1162 B.n651 B.n650 585
R1163 B.n649 B.n32 585
R1164 B.n648 B.n647 585
R1165 B.n646 B.n33 585
R1166 B.n645 B.n644 585
R1167 B.n643 B.n34 585
R1168 B.n642 B.n641 585
R1169 B.n640 B.n35 585
R1170 B.n639 B.n638 585
R1171 B.n637 B.n36 585
R1172 B.n636 B.n635 585
R1173 B.n634 B.n37 585
R1174 B.n633 B.n632 585
R1175 B.n631 B.n38 585
R1176 B.n630 B.n629 585
R1177 B.n628 B.n39 585
R1178 B.n627 B.n626 585
R1179 B.n625 B.n40 585
R1180 B.n624 B.n623 585
R1181 B.n622 B.n41 585
R1182 B.n621 B.n620 585
R1183 B.n619 B.n42 585
R1184 B.n618 B.n617 585
R1185 B.n616 B.n43 585
R1186 B.n615 B.n614 585
R1187 B.n613 B.n44 585
R1188 B.n612 B.n611 585
R1189 B.n609 B.n45 585
R1190 B.n608 B.n607 585
R1191 B.n606 B.n48 585
R1192 B.n605 B.n604 585
R1193 B.n603 B.n49 585
R1194 B.n602 B.n601 585
R1195 B.n600 B.n50 585
R1196 B.n599 B.n598 585
R1197 B.n597 B.n51 585
R1198 B.n595 B.n594 585
R1199 B.n593 B.n54 585
R1200 B.n592 B.n591 585
R1201 B.n590 B.n55 585
R1202 B.n589 B.n588 585
R1203 B.n587 B.n56 585
R1204 B.n586 B.n585 585
R1205 B.n584 B.n57 585
R1206 B.n583 B.n582 585
R1207 B.n581 B.n58 585
R1208 B.n580 B.n579 585
R1209 B.n578 B.n59 585
R1210 B.n577 B.n576 585
R1211 B.n575 B.n60 585
R1212 B.n574 B.n573 585
R1213 B.n572 B.n61 585
R1214 B.n571 B.n570 585
R1215 B.n569 B.n62 585
R1216 B.n568 B.n567 585
R1217 B.n566 B.n63 585
R1218 B.n565 B.n564 585
R1219 B.n563 B.n64 585
R1220 B.n562 B.n561 585
R1221 B.n560 B.n65 585
R1222 B.n559 B.n558 585
R1223 B.n557 B.n66 585
R1224 B.n556 B.n555 585
R1225 B.n554 B.n67 585
R1226 B.n553 B.n552 585
R1227 B.n551 B.n68 585
R1228 B.n550 B.n549 585
R1229 B.n548 B.n69 585
R1230 B.n547 B.n546 585
R1231 B.n545 B.n70 585
R1232 B.n544 B.n543 585
R1233 B.n542 B.n71 585
R1234 B.n541 B.n540 585
R1235 B.n539 B.n72 585
R1236 B.n538 B.n537 585
R1237 B.n536 B.n73 585
R1238 B.n535 B.n534 585
R1239 B.n533 B.n74 585
R1240 B.n532 B.n531 585
R1241 B.n530 B.n75 585
R1242 B.n529 B.n528 585
R1243 B.n527 B.n76 585
R1244 B.n526 B.n525 585
R1245 B.n524 B.n77 585
R1246 B.n523 B.n522 585
R1247 B.n521 B.n78 585
R1248 B.n520 B.n519 585
R1249 B.n518 B.n79 585
R1250 B.n517 B.n516 585
R1251 B.n515 B.n80 585
R1252 B.n514 B.n513 585
R1253 B.n512 B.n81 585
R1254 B.n511 B.n510 585
R1255 B.n509 B.n82 585
R1256 B.n508 B.n507 585
R1257 B.n506 B.n83 585
R1258 B.n505 B.n504 585
R1259 B.n503 B.n84 585
R1260 B.n705 B.n704 585
R1261 B.n706 B.n13 585
R1262 B.n708 B.n707 585
R1263 B.n709 B.n12 585
R1264 B.n711 B.n710 585
R1265 B.n712 B.n11 585
R1266 B.n714 B.n713 585
R1267 B.n715 B.n10 585
R1268 B.n717 B.n716 585
R1269 B.n718 B.n9 585
R1270 B.n720 B.n719 585
R1271 B.n721 B.n8 585
R1272 B.n723 B.n722 585
R1273 B.n724 B.n7 585
R1274 B.n726 B.n725 585
R1275 B.n727 B.n6 585
R1276 B.n729 B.n728 585
R1277 B.n730 B.n5 585
R1278 B.n732 B.n731 585
R1279 B.n733 B.n4 585
R1280 B.n735 B.n734 585
R1281 B.n736 B.n3 585
R1282 B.n738 B.n737 585
R1283 B.n739 B.n0 585
R1284 B.n2 B.n1 585
R1285 B.n190 B.n189 585
R1286 B.n192 B.n191 585
R1287 B.n193 B.n188 585
R1288 B.n195 B.n194 585
R1289 B.n196 B.n187 585
R1290 B.n198 B.n197 585
R1291 B.n199 B.n186 585
R1292 B.n201 B.n200 585
R1293 B.n202 B.n185 585
R1294 B.n204 B.n203 585
R1295 B.n205 B.n184 585
R1296 B.n207 B.n206 585
R1297 B.n208 B.n183 585
R1298 B.n210 B.n209 585
R1299 B.n211 B.n182 585
R1300 B.n213 B.n212 585
R1301 B.n214 B.n181 585
R1302 B.n216 B.n215 585
R1303 B.n217 B.n180 585
R1304 B.n219 B.n218 585
R1305 B.n220 B.n179 585
R1306 B.n222 B.n221 585
R1307 B.n223 B.n178 585
R1308 B.n330 B.t10 551.343
R1309 B.n52 B.t5 551.343
R1310 B.n146 B.t7 551.343
R1311 B.n46 B.t2 551.343
R1312 B.n331 B.t11 497.235
R1313 B.n53 B.t4 497.235
R1314 B.n147 B.t8 497.235
R1315 B.n47 B.t1 497.235
R1316 B.n224 B.n223 468.476
R1317 B.n426 B.n109 468.476
R1318 B.n503 B.n502 468.476
R1319 B.n704 B.n703 468.476
R1320 B.n146 B.t6 391.613
R1321 B.n330 B.t9 391.613
R1322 B.n52 B.t3 391.613
R1323 B.n46 B.t0 391.613
R1324 B.n741 B.n740 256.663
R1325 B.n740 B.n739 235.042
R1326 B.n740 B.n2 235.042
R1327 B.n224 B.n177 163.367
R1328 B.n228 B.n177 163.367
R1329 B.n229 B.n228 163.367
R1330 B.n230 B.n229 163.367
R1331 B.n230 B.n175 163.367
R1332 B.n234 B.n175 163.367
R1333 B.n235 B.n234 163.367
R1334 B.n236 B.n235 163.367
R1335 B.n236 B.n173 163.367
R1336 B.n240 B.n173 163.367
R1337 B.n241 B.n240 163.367
R1338 B.n242 B.n241 163.367
R1339 B.n242 B.n171 163.367
R1340 B.n246 B.n171 163.367
R1341 B.n247 B.n246 163.367
R1342 B.n248 B.n247 163.367
R1343 B.n248 B.n169 163.367
R1344 B.n252 B.n169 163.367
R1345 B.n253 B.n252 163.367
R1346 B.n254 B.n253 163.367
R1347 B.n254 B.n167 163.367
R1348 B.n258 B.n167 163.367
R1349 B.n259 B.n258 163.367
R1350 B.n260 B.n259 163.367
R1351 B.n260 B.n165 163.367
R1352 B.n264 B.n165 163.367
R1353 B.n265 B.n264 163.367
R1354 B.n266 B.n265 163.367
R1355 B.n266 B.n163 163.367
R1356 B.n270 B.n163 163.367
R1357 B.n271 B.n270 163.367
R1358 B.n272 B.n271 163.367
R1359 B.n272 B.n161 163.367
R1360 B.n276 B.n161 163.367
R1361 B.n277 B.n276 163.367
R1362 B.n278 B.n277 163.367
R1363 B.n278 B.n159 163.367
R1364 B.n282 B.n159 163.367
R1365 B.n283 B.n282 163.367
R1366 B.n284 B.n283 163.367
R1367 B.n284 B.n157 163.367
R1368 B.n288 B.n157 163.367
R1369 B.n289 B.n288 163.367
R1370 B.n290 B.n289 163.367
R1371 B.n290 B.n155 163.367
R1372 B.n294 B.n155 163.367
R1373 B.n295 B.n294 163.367
R1374 B.n296 B.n295 163.367
R1375 B.n296 B.n153 163.367
R1376 B.n300 B.n153 163.367
R1377 B.n301 B.n300 163.367
R1378 B.n302 B.n301 163.367
R1379 B.n302 B.n151 163.367
R1380 B.n306 B.n151 163.367
R1381 B.n307 B.n306 163.367
R1382 B.n308 B.n307 163.367
R1383 B.n308 B.n149 163.367
R1384 B.n312 B.n149 163.367
R1385 B.n313 B.n312 163.367
R1386 B.n314 B.n313 163.367
R1387 B.n314 B.n145 163.367
R1388 B.n319 B.n145 163.367
R1389 B.n320 B.n319 163.367
R1390 B.n321 B.n320 163.367
R1391 B.n321 B.n143 163.367
R1392 B.n325 B.n143 163.367
R1393 B.n326 B.n325 163.367
R1394 B.n327 B.n326 163.367
R1395 B.n327 B.n141 163.367
R1396 B.n334 B.n141 163.367
R1397 B.n335 B.n334 163.367
R1398 B.n336 B.n335 163.367
R1399 B.n336 B.n139 163.367
R1400 B.n340 B.n139 163.367
R1401 B.n341 B.n340 163.367
R1402 B.n342 B.n341 163.367
R1403 B.n342 B.n137 163.367
R1404 B.n346 B.n137 163.367
R1405 B.n347 B.n346 163.367
R1406 B.n348 B.n347 163.367
R1407 B.n348 B.n135 163.367
R1408 B.n352 B.n135 163.367
R1409 B.n353 B.n352 163.367
R1410 B.n354 B.n353 163.367
R1411 B.n354 B.n133 163.367
R1412 B.n358 B.n133 163.367
R1413 B.n359 B.n358 163.367
R1414 B.n360 B.n359 163.367
R1415 B.n360 B.n131 163.367
R1416 B.n364 B.n131 163.367
R1417 B.n365 B.n364 163.367
R1418 B.n366 B.n365 163.367
R1419 B.n366 B.n129 163.367
R1420 B.n370 B.n129 163.367
R1421 B.n371 B.n370 163.367
R1422 B.n372 B.n371 163.367
R1423 B.n372 B.n127 163.367
R1424 B.n376 B.n127 163.367
R1425 B.n377 B.n376 163.367
R1426 B.n378 B.n377 163.367
R1427 B.n378 B.n125 163.367
R1428 B.n382 B.n125 163.367
R1429 B.n383 B.n382 163.367
R1430 B.n384 B.n383 163.367
R1431 B.n384 B.n123 163.367
R1432 B.n388 B.n123 163.367
R1433 B.n389 B.n388 163.367
R1434 B.n390 B.n389 163.367
R1435 B.n390 B.n121 163.367
R1436 B.n394 B.n121 163.367
R1437 B.n395 B.n394 163.367
R1438 B.n396 B.n395 163.367
R1439 B.n396 B.n119 163.367
R1440 B.n400 B.n119 163.367
R1441 B.n401 B.n400 163.367
R1442 B.n402 B.n401 163.367
R1443 B.n402 B.n117 163.367
R1444 B.n406 B.n117 163.367
R1445 B.n407 B.n406 163.367
R1446 B.n408 B.n407 163.367
R1447 B.n408 B.n115 163.367
R1448 B.n412 B.n115 163.367
R1449 B.n413 B.n412 163.367
R1450 B.n414 B.n413 163.367
R1451 B.n414 B.n113 163.367
R1452 B.n418 B.n113 163.367
R1453 B.n419 B.n418 163.367
R1454 B.n420 B.n419 163.367
R1455 B.n420 B.n111 163.367
R1456 B.n424 B.n111 163.367
R1457 B.n425 B.n424 163.367
R1458 B.n426 B.n425 163.367
R1459 B.n502 B.n85 163.367
R1460 B.n498 B.n85 163.367
R1461 B.n498 B.n497 163.367
R1462 B.n497 B.n496 163.367
R1463 B.n496 B.n87 163.367
R1464 B.n492 B.n87 163.367
R1465 B.n492 B.n491 163.367
R1466 B.n491 B.n490 163.367
R1467 B.n490 B.n89 163.367
R1468 B.n486 B.n89 163.367
R1469 B.n486 B.n485 163.367
R1470 B.n485 B.n484 163.367
R1471 B.n484 B.n91 163.367
R1472 B.n480 B.n91 163.367
R1473 B.n480 B.n479 163.367
R1474 B.n479 B.n478 163.367
R1475 B.n478 B.n93 163.367
R1476 B.n474 B.n93 163.367
R1477 B.n474 B.n473 163.367
R1478 B.n473 B.n472 163.367
R1479 B.n472 B.n95 163.367
R1480 B.n468 B.n95 163.367
R1481 B.n468 B.n467 163.367
R1482 B.n467 B.n466 163.367
R1483 B.n466 B.n97 163.367
R1484 B.n462 B.n97 163.367
R1485 B.n462 B.n461 163.367
R1486 B.n461 B.n460 163.367
R1487 B.n460 B.n99 163.367
R1488 B.n456 B.n99 163.367
R1489 B.n456 B.n455 163.367
R1490 B.n455 B.n454 163.367
R1491 B.n454 B.n101 163.367
R1492 B.n450 B.n101 163.367
R1493 B.n450 B.n449 163.367
R1494 B.n449 B.n448 163.367
R1495 B.n448 B.n103 163.367
R1496 B.n444 B.n103 163.367
R1497 B.n444 B.n443 163.367
R1498 B.n443 B.n442 163.367
R1499 B.n442 B.n105 163.367
R1500 B.n438 B.n105 163.367
R1501 B.n438 B.n437 163.367
R1502 B.n437 B.n436 163.367
R1503 B.n436 B.n107 163.367
R1504 B.n432 B.n107 163.367
R1505 B.n432 B.n431 163.367
R1506 B.n431 B.n430 163.367
R1507 B.n430 B.n109 163.367
R1508 B.n703 B.n702 163.367
R1509 B.n702 B.n15 163.367
R1510 B.n698 B.n15 163.367
R1511 B.n698 B.n697 163.367
R1512 B.n697 B.n696 163.367
R1513 B.n696 B.n17 163.367
R1514 B.n692 B.n17 163.367
R1515 B.n692 B.n691 163.367
R1516 B.n691 B.n690 163.367
R1517 B.n690 B.n19 163.367
R1518 B.n686 B.n19 163.367
R1519 B.n686 B.n685 163.367
R1520 B.n685 B.n684 163.367
R1521 B.n684 B.n21 163.367
R1522 B.n680 B.n21 163.367
R1523 B.n680 B.n679 163.367
R1524 B.n679 B.n678 163.367
R1525 B.n678 B.n23 163.367
R1526 B.n674 B.n23 163.367
R1527 B.n674 B.n673 163.367
R1528 B.n673 B.n672 163.367
R1529 B.n672 B.n25 163.367
R1530 B.n668 B.n25 163.367
R1531 B.n668 B.n667 163.367
R1532 B.n667 B.n666 163.367
R1533 B.n666 B.n27 163.367
R1534 B.n662 B.n27 163.367
R1535 B.n662 B.n661 163.367
R1536 B.n661 B.n660 163.367
R1537 B.n660 B.n29 163.367
R1538 B.n656 B.n29 163.367
R1539 B.n656 B.n655 163.367
R1540 B.n655 B.n654 163.367
R1541 B.n654 B.n31 163.367
R1542 B.n650 B.n31 163.367
R1543 B.n650 B.n649 163.367
R1544 B.n649 B.n648 163.367
R1545 B.n648 B.n33 163.367
R1546 B.n644 B.n33 163.367
R1547 B.n644 B.n643 163.367
R1548 B.n643 B.n642 163.367
R1549 B.n642 B.n35 163.367
R1550 B.n638 B.n35 163.367
R1551 B.n638 B.n637 163.367
R1552 B.n637 B.n636 163.367
R1553 B.n636 B.n37 163.367
R1554 B.n632 B.n37 163.367
R1555 B.n632 B.n631 163.367
R1556 B.n631 B.n630 163.367
R1557 B.n630 B.n39 163.367
R1558 B.n626 B.n39 163.367
R1559 B.n626 B.n625 163.367
R1560 B.n625 B.n624 163.367
R1561 B.n624 B.n41 163.367
R1562 B.n620 B.n41 163.367
R1563 B.n620 B.n619 163.367
R1564 B.n619 B.n618 163.367
R1565 B.n618 B.n43 163.367
R1566 B.n614 B.n43 163.367
R1567 B.n614 B.n613 163.367
R1568 B.n613 B.n612 163.367
R1569 B.n612 B.n45 163.367
R1570 B.n607 B.n45 163.367
R1571 B.n607 B.n606 163.367
R1572 B.n606 B.n605 163.367
R1573 B.n605 B.n49 163.367
R1574 B.n601 B.n49 163.367
R1575 B.n601 B.n600 163.367
R1576 B.n600 B.n599 163.367
R1577 B.n599 B.n51 163.367
R1578 B.n594 B.n51 163.367
R1579 B.n594 B.n593 163.367
R1580 B.n593 B.n592 163.367
R1581 B.n592 B.n55 163.367
R1582 B.n588 B.n55 163.367
R1583 B.n588 B.n587 163.367
R1584 B.n587 B.n586 163.367
R1585 B.n586 B.n57 163.367
R1586 B.n582 B.n57 163.367
R1587 B.n582 B.n581 163.367
R1588 B.n581 B.n580 163.367
R1589 B.n580 B.n59 163.367
R1590 B.n576 B.n59 163.367
R1591 B.n576 B.n575 163.367
R1592 B.n575 B.n574 163.367
R1593 B.n574 B.n61 163.367
R1594 B.n570 B.n61 163.367
R1595 B.n570 B.n569 163.367
R1596 B.n569 B.n568 163.367
R1597 B.n568 B.n63 163.367
R1598 B.n564 B.n63 163.367
R1599 B.n564 B.n563 163.367
R1600 B.n563 B.n562 163.367
R1601 B.n562 B.n65 163.367
R1602 B.n558 B.n65 163.367
R1603 B.n558 B.n557 163.367
R1604 B.n557 B.n556 163.367
R1605 B.n556 B.n67 163.367
R1606 B.n552 B.n67 163.367
R1607 B.n552 B.n551 163.367
R1608 B.n551 B.n550 163.367
R1609 B.n550 B.n69 163.367
R1610 B.n546 B.n69 163.367
R1611 B.n546 B.n545 163.367
R1612 B.n545 B.n544 163.367
R1613 B.n544 B.n71 163.367
R1614 B.n540 B.n71 163.367
R1615 B.n540 B.n539 163.367
R1616 B.n539 B.n538 163.367
R1617 B.n538 B.n73 163.367
R1618 B.n534 B.n73 163.367
R1619 B.n534 B.n533 163.367
R1620 B.n533 B.n532 163.367
R1621 B.n532 B.n75 163.367
R1622 B.n528 B.n75 163.367
R1623 B.n528 B.n527 163.367
R1624 B.n527 B.n526 163.367
R1625 B.n526 B.n77 163.367
R1626 B.n522 B.n77 163.367
R1627 B.n522 B.n521 163.367
R1628 B.n521 B.n520 163.367
R1629 B.n520 B.n79 163.367
R1630 B.n516 B.n79 163.367
R1631 B.n516 B.n515 163.367
R1632 B.n515 B.n514 163.367
R1633 B.n514 B.n81 163.367
R1634 B.n510 B.n81 163.367
R1635 B.n510 B.n509 163.367
R1636 B.n509 B.n508 163.367
R1637 B.n508 B.n83 163.367
R1638 B.n504 B.n83 163.367
R1639 B.n504 B.n503 163.367
R1640 B.n704 B.n13 163.367
R1641 B.n708 B.n13 163.367
R1642 B.n709 B.n708 163.367
R1643 B.n710 B.n709 163.367
R1644 B.n710 B.n11 163.367
R1645 B.n714 B.n11 163.367
R1646 B.n715 B.n714 163.367
R1647 B.n716 B.n715 163.367
R1648 B.n716 B.n9 163.367
R1649 B.n720 B.n9 163.367
R1650 B.n721 B.n720 163.367
R1651 B.n722 B.n721 163.367
R1652 B.n722 B.n7 163.367
R1653 B.n726 B.n7 163.367
R1654 B.n727 B.n726 163.367
R1655 B.n728 B.n727 163.367
R1656 B.n728 B.n5 163.367
R1657 B.n732 B.n5 163.367
R1658 B.n733 B.n732 163.367
R1659 B.n734 B.n733 163.367
R1660 B.n734 B.n3 163.367
R1661 B.n738 B.n3 163.367
R1662 B.n739 B.n738 163.367
R1663 B.n189 B.n2 163.367
R1664 B.n192 B.n189 163.367
R1665 B.n193 B.n192 163.367
R1666 B.n194 B.n193 163.367
R1667 B.n194 B.n187 163.367
R1668 B.n198 B.n187 163.367
R1669 B.n199 B.n198 163.367
R1670 B.n200 B.n199 163.367
R1671 B.n200 B.n185 163.367
R1672 B.n204 B.n185 163.367
R1673 B.n205 B.n204 163.367
R1674 B.n206 B.n205 163.367
R1675 B.n206 B.n183 163.367
R1676 B.n210 B.n183 163.367
R1677 B.n211 B.n210 163.367
R1678 B.n212 B.n211 163.367
R1679 B.n212 B.n181 163.367
R1680 B.n216 B.n181 163.367
R1681 B.n217 B.n216 163.367
R1682 B.n218 B.n217 163.367
R1683 B.n218 B.n179 163.367
R1684 B.n222 B.n179 163.367
R1685 B.n223 B.n222 163.367
R1686 B.n317 B.n147 59.5399
R1687 B.n332 B.n331 59.5399
R1688 B.n596 B.n53 59.5399
R1689 B.n610 B.n47 59.5399
R1690 B.n147 B.n146 54.1096
R1691 B.n331 B.n330 54.1096
R1692 B.n53 B.n52 54.1096
R1693 B.n47 B.n46 54.1096
R1694 B.n428 B.n427 30.4395
R1695 B.n705 B.n14 30.4395
R1696 B.n501 B.n84 30.4395
R1697 B.n225 B.n178 30.4395
R1698 B B.n741 18.0485
R1699 B.n706 B.n705 10.6151
R1700 B.n707 B.n706 10.6151
R1701 B.n707 B.n12 10.6151
R1702 B.n711 B.n12 10.6151
R1703 B.n712 B.n711 10.6151
R1704 B.n713 B.n712 10.6151
R1705 B.n713 B.n10 10.6151
R1706 B.n717 B.n10 10.6151
R1707 B.n718 B.n717 10.6151
R1708 B.n719 B.n718 10.6151
R1709 B.n719 B.n8 10.6151
R1710 B.n723 B.n8 10.6151
R1711 B.n724 B.n723 10.6151
R1712 B.n725 B.n724 10.6151
R1713 B.n725 B.n6 10.6151
R1714 B.n729 B.n6 10.6151
R1715 B.n730 B.n729 10.6151
R1716 B.n731 B.n730 10.6151
R1717 B.n731 B.n4 10.6151
R1718 B.n735 B.n4 10.6151
R1719 B.n736 B.n735 10.6151
R1720 B.n737 B.n736 10.6151
R1721 B.n737 B.n0 10.6151
R1722 B.n701 B.n14 10.6151
R1723 B.n701 B.n700 10.6151
R1724 B.n700 B.n699 10.6151
R1725 B.n699 B.n16 10.6151
R1726 B.n695 B.n16 10.6151
R1727 B.n695 B.n694 10.6151
R1728 B.n694 B.n693 10.6151
R1729 B.n693 B.n18 10.6151
R1730 B.n689 B.n18 10.6151
R1731 B.n689 B.n688 10.6151
R1732 B.n688 B.n687 10.6151
R1733 B.n687 B.n20 10.6151
R1734 B.n683 B.n20 10.6151
R1735 B.n683 B.n682 10.6151
R1736 B.n682 B.n681 10.6151
R1737 B.n681 B.n22 10.6151
R1738 B.n677 B.n22 10.6151
R1739 B.n677 B.n676 10.6151
R1740 B.n676 B.n675 10.6151
R1741 B.n675 B.n24 10.6151
R1742 B.n671 B.n24 10.6151
R1743 B.n671 B.n670 10.6151
R1744 B.n670 B.n669 10.6151
R1745 B.n669 B.n26 10.6151
R1746 B.n665 B.n26 10.6151
R1747 B.n665 B.n664 10.6151
R1748 B.n664 B.n663 10.6151
R1749 B.n663 B.n28 10.6151
R1750 B.n659 B.n28 10.6151
R1751 B.n659 B.n658 10.6151
R1752 B.n658 B.n657 10.6151
R1753 B.n657 B.n30 10.6151
R1754 B.n653 B.n30 10.6151
R1755 B.n653 B.n652 10.6151
R1756 B.n652 B.n651 10.6151
R1757 B.n651 B.n32 10.6151
R1758 B.n647 B.n32 10.6151
R1759 B.n647 B.n646 10.6151
R1760 B.n646 B.n645 10.6151
R1761 B.n645 B.n34 10.6151
R1762 B.n641 B.n34 10.6151
R1763 B.n641 B.n640 10.6151
R1764 B.n640 B.n639 10.6151
R1765 B.n639 B.n36 10.6151
R1766 B.n635 B.n36 10.6151
R1767 B.n635 B.n634 10.6151
R1768 B.n634 B.n633 10.6151
R1769 B.n633 B.n38 10.6151
R1770 B.n629 B.n38 10.6151
R1771 B.n629 B.n628 10.6151
R1772 B.n628 B.n627 10.6151
R1773 B.n627 B.n40 10.6151
R1774 B.n623 B.n40 10.6151
R1775 B.n623 B.n622 10.6151
R1776 B.n622 B.n621 10.6151
R1777 B.n621 B.n42 10.6151
R1778 B.n617 B.n42 10.6151
R1779 B.n617 B.n616 10.6151
R1780 B.n616 B.n615 10.6151
R1781 B.n615 B.n44 10.6151
R1782 B.n611 B.n44 10.6151
R1783 B.n609 B.n608 10.6151
R1784 B.n608 B.n48 10.6151
R1785 B.n604 B.n48 10.6151
R1786 B.n604 B.n603 10.6151
R1787 B.n603 B.n602 10.6151
R1788 B.n602 B.n50 10.6151
R1789 B.n598 B.n50 10.6151
R1790 B.n598 B.n597 10.6151
R1791 B.n595 B.n54 10.6151
R1792 B.n591 B.n54 10.6151
R1793 B.n591 B.n590 10.6151
R1794 B.n590 B.n589 10.6151
R1795 B.n589 B.n56 10.6151
R1796 B.n585 B.n56 10.6151
R1797 B.n585 B.n584 10.6151
R1798 B.n584 B.n583 10.6151
R1799 B.n583 B.n58 10.6151
R1800 B.n579 B.n58 10.6151
R1801 B.n579 B.n578 10.6151
R1802 B.n578 B.n577 10.6151
R1803 B.n577 B.n60 10.6151
R1804 B.n573 B.n60 10.6151
R1805 B.n573 B.n572 10.6151
R1806 B.n572 B.n571 10.6151
R1807 B.n571 B.n62 10.6151
R1808 B.n567 B.n62 10.6151
R1809 B.n567 B.n566 10.6151
R1810 B.n566 B.n565 10.6151
R1811 B.n565 B.n64 10.6151
R1812 B.n561 B.n64 10.6151
R1813 B.n561 B.n560 10.6151
R1814 B.n560 B.n559 10.6151
R1815 B.n559 B.n66 10.6151
R1816 B.n555 B.n66 10.6151
R1817 B.n555 B.n554 10.6151
R1818 B.n554 B.n553 10.6151
R1819 B.n553 B.n68 10.6151
R1820 B.n549 B.n68 10.6151
R1821 B.n549 B.n548 10.6151
R1822 B.n548 B.n547 10.6151
R1823 B.n547 B.n70 10.6151
R1824 B.n543 B.n70 10.6151
R1825 B.n543 B.n542 10.6151
R1826 B.n542 B.n541 10.6151
R1827 B.n541 B.n72 10.6151
R1828 B.n537 B.n72 10.6151
R1829 B.n537 B.n536 10.6151
R1830 B.n536 B.n535 10.6151
R1831 B.n535 B.n74 10.6151
R1832 B.n531 B.n74 10.6151
R1833 B.n531 B.n530 10.6151
R1834 B.n530 B.n529 10.6151
R1835 B.n529 B.n76 10.6151
R1836 B.n525 B.n76 10.6151
R1837 B.n525 B.n524 10.6151
R1838 B.n524 B.n523 10.6151
R1839 B.n523 B.n78 10.6151
R1840 B.n519 B.n78 10.6151
R1841 B.n519 B.n518 10.6151
R1842 B.n518 B.n517 10.6151
R1843 B.n517 B.n80 10.6151
R1844 B.n513 B.n80 10.6151
R1845 B.n513 B.n512 10.6151
R1846 B.n512 B.n511 10.6151
R1847 B.n511 B.n82 10.6151
R1848 B.n507 B.n82 10.6151
R1849 B.n507 B.n506 10.6151
R1850 B.n506 B.n505 10.6151
R1851 B.n505 B.n84 10.6151
R1852 B.n501 B.n500 10.6151
R1853 B.n500 B.n499 10.6151
R1854 B.n499 B.n86 10.6151
R1855 B.n495 B.n86 10.6151
R1856 B.n495 B.n494 10.6151
R1857 B.n494 B.n493 10.6151
R1858 B.n493 B.n88 10.6151
R1859 B.n489 B.n88 10.6151
R1860 B.n489 B.n488 10.6151
R1861 B.n488 B.n487 10.6151
R1862 B.n487 B.n90 10.6151
R1863 B.n483 B.n90 10.6151
R1864 B.n483 B.n482 10.6151
R1865 B.n482 B.n481 10.6151
R1866 B.n481 B.n92 10.6151
R1867 B.n477 B.n92 10.6151
R1868 B.n477 B.n476 10.6151
R1869 B.n476 B.n475 10.6151
R1870 B.n475 B.n94 10.6151
R1871 B.n471 B.n94 10.6151
R1872 B.n471 B.n470 10.6151
R1873 B.n470 B.n469 10.6151
R1874 B.n469 B.n96 10.6151
R1875 B.n465 B.n96 10.6151
R1876 B.n465 B.n464 10.6151
R1877 B.n464 B.n463 10.6151
R1878 B.n463 B.n98 10.6151
R1879 B.n459 B.n98 10.6151
R1880 B.n459 B.n458 10.6151
R1881 B.n458 B.n457 10.6151
R1882 B.n457 B.n100 10.6151
R1883 B.n453 B.n100 10.6151
R1884 B.n453 B.n452 10.6151
R1885 B.n452 B.n451 10.6151
R1886 B.n451 B.n102 10.6151
R1887 B.n447 B.n102 10.6151
R1888 B.n447 B.n446 10.6151
R1889 B.n446 B.n445 10.6151
R1890 B.n445 B.n104 10.6151
R1891 B.n441 B.n104 10.6151
R1892 B.n441 B.n440 10.6151
R1893 B.n440 B.n439 10.6151
R1894 B.n439 B.n106 10.6151
R1895 B.n435 B.n106 10.6151
R1896 B.n435 B.n434 10.6151
R1897 B.n434 B.n433 10.6151
R1898 B.n433 B.n108 10.6151
R1899 B.n429 B.n108 10.6151
R1900 B.n429 B.n428 10.6151
R1901 B.n190 B.n1 10.6151
R1902 B.n191 B.n190 10.6151
R1903 B.n191 B.n188 10.6151
R1904 B.n195 B.n188 10.6151
R1905 B.n196 B.n195 10.6151
R1906 B.n197 B.n196 10.6151
R1907 B.n197 B.n186 10.6151
R1908 B.n201 B.n186 10.6151
R1909 B.n202 B.n201 10.6151
R1910 B.n203 B.n202 10.6151
R1911 B.n203 B.n184 10.6151
R1912 B.n207 B.n184 10.6151
R1913 B.n208 B.n207 10.6151
R1914 B.n209 B.n208 10.6151
R1915 B.n209 B.n182 10.6151
R1916 B.n213 B.n182 10.6151
R1917 B.n214 B.n213 10.6151
R1918 B.n215 B.n214 10.6151
R1919 B.n215 B.n180 10.6151
R1920 B.n219 B.n180 10.6151
R1921 B.n220 B.n219 10.6151
R1922 B.n221 B.n220 10.6151
R1923 B.n221 B.n178 10.6151
R1924 B.n226 B.n225 10.6151
R1925 B.n227 B.n226 10.6151
R1926 B.n227 B.n176 10.6151
R1927 B.n231 B.n176 10.6151
R1928 B.n232 B.n231 10.6151
R1929 B.n233 B.n232 10.6151
R1930 B.n233 B.n174 10.6151
R1931 B.n237 B.n174 10.6151
R1932 B.n238 B.n237 10.6151
R1933 B.n239 B.n238 10.6151
R1934 B.n239 B.n172 10.6151
R1935 B.n243 B.n172 10.6151
R1936 B.n244 B.n243 10.6151
R1937 B.n245 B.n244 10.6151
R1938 B.n245 B.n170 10.6151
R1939 B.n249 B.n170 10.6151
R1940 B.n250 B.n249 10.6151
R1941 B.n251 B.n250 10.6151
R1942 B.n251 B.n168 10.6151
R1943 B.n255 B.n168 10.6151
R1944 B.n256 B.n255 10.6151
R1945 B.n257 B.n256 10.6151
R1946 B.n257 B.n166 10.6151
R1947 B.n261 B.n166 10.6151
R1948 B.n262 B.n261 10.6151
R1949 B.n263 B.n262 10.6151
R1950 B.n263 B.n164 10.6151
R1951 B.n267 B.n164 10.6151
R1952 B.n268 B.n267 10.6151
R1953 B.n269 B.n268 10.6151
R1954 B.n269 B.n162 10.6151
R1955 B.n273 B.n162 10.6151
R1956 B.n274 B.n273 10.6151
R1957 B.n275 B.n274 10.6151
R1958 B.n275 B.n160 10.6151
R1959 B.n279 B.n160 10.6151
R1960 B.n280 B.n279 10.6151
R1961 B.n281 B.n280 10.6151
R1962 B.n281 B.n158 10.6151
R1963 B.n285 B.n158 10.6151
R1964 B.n286 B.n285 10.6151
R1965 B.n287 B.n286 10.6151
R1966 B.n287 B.n156 10.6151
R1967 B.n291 B.n156 10.6151
R1968 B.n292 B.n291 10.6151
R1969 B.n293 B.n292 10.6151
R1970 B.n293 B.n154 10.6151
R1971 B.n297 B.n154 10.6151
R1972 B.n298 B.n297 10.6151
R1973 B.n299 B.n298 10.6151
R1974 B.n299 B.n152 10.6151
R1975 B.n303 B.n152 10.6151
R1976 B.n304 B.n303 10.6151
R1977 B.n305 B.n304 10.6151
R1978 B.n305 B.n150 10.6151
R1979 B.n309 B.n150 10.6151
R1980 B.n310 B.n309 10.6151
R1981 B.n311 B.n310 10.6151
R1982 B.n311 B.n148 10.6151
R1983 B.n315 B.n148 10.6151
R1984 B.n316 B.n315 10.6151
R1985 B.n318 B.n144 10.6151
R1986 B.n322 B.n144 10.6151
R1987 B.n323 B.n322 10.6151
R1988 B.n324 B.n323 10.6151
R1989 B.n324 B.n142 10.6151
R1990 B.n328 B.n142 10.6151
R1991 B.n329 B.n328 10.6151
R1992 B.n333 B.n329 10.6151
R1993 B.n337 B.n140 10.6151
R1994 B.n338 B.n337 10.6151
R1995 B.n339 B.n338 10.6151
R1996 B.n339 B.n138 10.6151
R1997 B.n343 B.n138 10.6151
R1998 B.n344 B.n343 10.6151
R1999 B.n345 B.n344 10.6151
R2000 B.n345 B.n136 10.6151
R2001 B.n349 B.n136 10.6151
R2002 B.n350 B.n349 10.6151
R2003 B.n351 B.n350 10.6151
R2004 B.n351 B.n134 10.6151
R2005 B.n355 B.n134 10.6151
R2006 B.n356 B.n355 10.6151
R2007 B.n357 B.n356 10.6151
R2008 B.n357 B.n132 10.6151
R2009 B.n361 B.n132 10.6151
R2010 B.n362 B.n361 10.6151
R2011 B.n363 B.n362 10.6151
R2012 B.n363 B.n130 10.6151
R2013 B.n367 B.n130 10.6151
R2014 B.n368 B.n367 10.6151
R2015 B.n369 B.n368 10.6151
R2016 B.n369 B.n128 10.6151
R2017 B.n373 B.n128 10.6151
R2018 B.n374 B.n373 10.6151
R2019 B.n375 B.n374 10.6151
R2020 B.n375 B.n126 10.6151
R2021 B.n379 B.n126 10.6151
R2022 B.n380 B.n379 10.6151
R2023 B.n381 B.n380 10.6151
R2024 B.n381 B.n124 10.6151
R2025 B.n385 B.n124 10.6151
R2026 B.n386 B.n385 10.6151
R2027 B.n387 B.n386 10.6151
R2028 B.n387 B.n122 10.6151
R2029 B.n391 B.n122 10.6151
R2030 B.n392 B.n391 10.6151
R2031 B.n393 B.n392 10.6151
R2032 B.n393 B.n120 10.6151
R2033 B.n397 B.n120 10.6151
R2034 B.n398 B.n397 10.6151
R2035 B.n399 B.n398 10.6151
R2036 B.n399 B.n118 10.6151
R2037 B.n403 B.n118 10.6151
R2038 B.n404 B.n403 10.6151
R2039 B.n405 B.n404 10.6151
R2040 B.n405 B.n116 10.6151
R2041 B.n409 B.n116 10.6151
R2042 B.n410 B.n409 10.6151
R2043 B.n411 B.n410 10.6151
R2044 B.n411 B.n114 10.6151
R2045 B.n415 B.n114 10.6151
R2046 B.n416 B.n415 10.6151
R2047 B.n417 B.n416 10.6151
R2048 B.n417 B.n112 10.6151
R2049 B.n421 B.n112 10.6151
R2050 B.n422 B.n421 10.6151
R2051 B.n423 B.n422 10.6151
R2052 B.n423 B.n110 10.6151
R2053 B.n427 B.n110 10.6151
R2054 B.n741 B.n0 8.11757
R2055 B.n741 B.n1 8.11757
R2056 B.n610 B.n609 6.5566
R2057 B.n597 B.n596 6.5566
R2058 B.n318 B.n317 6.5566
R2059 B.n333 B.n332 6.5566
R2060 B.n611 B.n610 4.05904
R2061 B.n596 B.n595 4.05904
R2062 B.n317 B.n316 4.05904
R2063 B.n332 B.n140 4.05904
R2064 VP.n0 VP.t0 282.32
R2065 VP.n0 VP.t1 232.913
R2066 VP VP.n0 0.336784
R2067 VDD1.n102 VDD1.n101 756.745
R2068 VDD1.n205 VDD1.n204 756.745
R2069 VDD1.n101 VDD1.n100 585
R2070 VDD1.n2 VDD1.n1 585
R2071 VDD1.n95 VDD1.n94 585
R2072 VDD1.n93 VDD1.n92 585
R2073 VDD1.n6 VDD1.n5 585
R2074 VDD1.n87 VDD1.n86 585
R2075 VDD1.n85 VDD1.n84 585
R2076 VDD1.n10 VDD1.n9 585
R2077 VDD1.n79 VDD1.n78 585
R2078 VDD1.n77 VDD1.n76 585
R2079 VDD1.n14 VDD1.n13 585
R2080 VDD1.n71 VDD1.n70 585
R2081 VDD1.n69 VDD1.n68 585
R2082 VDD1.n18 VDD1.n17 585
R2083 VDD1.n63 VDD1.n62 585
R2084 VDD1.n61 VDD1.n60 585
R2085 VDD1.n22 VDD1.n21 585
R2086 VDD1.n26 VDD1.n24 585
R2087 VDD1.n55 VDD1.n54 585
R2088 VDD1.n53 VDD1.n52 585
R2089 VDD1.n28 VDD1.n27 585
R2090 VDD1.n47 VDD1.n46 585
R2091 VDD1.n45 VDD1.n44 585
R2092 VDD1.n32 VDD1.n31 585
R2093 VDD1.n39 VDD1.n38 585
R2094 VDD1.n37 VDD1.n36 585
R2095 VDD1.n138 VDD1.n137 585
R2096 VDD1.n140 VDD1.n139 585
R2097 VDD1.n133 VDD1.n132 585
R2098 VDD1.n146 VDD1.n145 585
R2099 VDD1.n148 VDD1.n147 585
R2100 VDD1.n129 VDD1.n128 585
R2101 VDD1.n155 VDD1.n154 585
R2102 VDD1.n156 VDD1.n127 585
R2103 VDD1.n158 VDD1.n157 585
R2104 VDD1.n125 VDD1.n124 585
R2105 VDD1.n164 VDD1.n163 585
R2106 VDD1.n166 VDD1.n165 585
R2107 VDD1.n121 VDD1.n120 585
R2108 VDD1.n172 VDD1.n171 585
R2109 VDD1.n174 VDD1.n173 585
R2110 VDD1.n117 VDD1.n116 585
R2111 VDD1.n180 VDD1.n179 585
R2112 VDD1.n182 VDD1.n181 585
R2113 VDD1.n113 VDD1.n112 585
R2114 VDD1.n188 VDD1.n187 585
R2115 VDD1.n190 VDD1.n189 585
R2116 VDD1.n109 VDD1.n108 585
R2117 VDD1.n196 VDD1.n195 585
R2118 VDD1.n198 VDD1.n197 585
R2119 VDD1.n105 VDD1.n104 585
R2120 VDD1.n204 VDD1.n203 585
R2121 VDD1.n35 VDD1.t1 329.036
R2122 VDD1.n136 VDD1.t0 329.036
R2123 VDD1.n101 VDD1.n1 171.744
R2124 VDD1.n94 VDD1.n1 171.744
R2125 VDD1.n94 VDD1.n93 171.744
R2126 VDD1.n93 VDD1.n5 171.744
R2127 VDD1.n86 VDD1.n5 171.744
R2128 VDD1.n86 VDD1.n85 171.744
R2129 VDD1.n85 VDD1.n9 171.744
R2130 VDD1.n78 VDD1.n9 171.744
R2131 VDD1.n78 VDD1.n77 171.744
R2132 VDD1.n77 VDD1.n13 171.744
R2133 VDD1.n70 VDD1.n13 171.744
R2134 VDD1.n70 VDD1.n69 171.744
R2135 VDD1.n69 VDD1.n17 171.744
R2136 VDD1.n62 VDD1.n17 171.744
R2137 VDD1.n62 VDD1.n61 171.744
R2138 VDD1.n61 VDD1.n21 171.744
R2139 VDD1.n26 VDD1.n21 171.744
R2140 VDD1.n54 VDD1.n26 171.744
R2141 VDD1.n54 VDD1.n53 171.744
R2142 VDD1.n53 VDD1.n27 171.744
R2143 VDD1.n46 VDD1.n27 171.744
R2144 VDD1.n46 VDD1.n45 171.744
R2145 VDD1.n45 VDD1.n31 171.744
R2146 VDD1.n38 VDD1.n31 171.744
R2147 VDD1.n38 VDD1.n37 171.744
R2148 VDD1.n139 VDD1.n138 171.744
R2149 VDD1.n139 VDD1.n132 171.744
R2150 VDD1.n146 VDD1.n132 171.744
R2151 VDD1.n147 VDD1.n146 171.744
R2152 VDD1.n147 VDD1.n128 171.744
R2153 VDD1.n155 VDD1.n128 171.744
R2154 VDD1.n156 VDD1.n155 171.744
R2155 VDD1.n157 VDD1.n156 171.744
R2156 VDD1.n157 VDD1.n124 171.744
R2157 VDD1.n164 VDD1.n124 171.744
R2158 VDD1.n165 VDD1.n164 171.744
R2159 VDD1.n165 VDD1.n120 171.744
R2160 VDD1.n172 VDD1.n120 171.744
R2161 VDD1.n173 VDD1.n172 171.744
R2162 VDD1.n173 VDD1.n116 171.744
R2163 VDD1.n180 VDD1.n116 171.744
R2164 VDD1.n181 VDD1.n180 171.744
R2165 VDD1.n181 VDD1.n112 171.744
R2166 VDD1.n188 VDD1.n112 171.744
R2167 VDD1.n189 VDD1.n188 171.744
R2168 VDD1.n189 VDD1.n108 171.744
R2169 VDD1.n196 VDD1.n108 171.744
R2170 VDD1.n197 VDD1.n196 171.744
R2171 VDD1.n197 VDD1.n104 171.744
R2172 VDD1.n204 VDD1.n104 171.744
R2173 VDD1 VDD1.n205 97.3476
R2174 VDD1.n37 VDD1.t1 85.8723
R2175 VDD1.n138 VDD1.t0 85.8723
R2176 VDD1 VDD1.n102 52.2388
R2177 VDD1.n24 VDD1.n22 13.1884
R2178 VDD1.n158 VDD1.n125 13.1884
R2179 VDD1.n100 VDD1.n0 12.8005
R2180 VDD1.n60 VDD1.n59 12.8005
R2181 VDD1.n56 VDD1.n55 12.8005
R2182 VDD1.n159 VDD1.n127 12.8005
R2183 VDD1.n163 VDD1.n162 12.8005
R2184 VDD1.n203 VDD1.n103 12.8005
R2185 VDD1.n99 VDD1.n2 12.0247
R2186 VDD1.n63 VDD1.n20 12.0247
R2187 VDD1.n52 VDD1.n25 12.0247
R2188 VDD1.n154 VDD1.n153 12.0247
R2189 VDD1.n166 VDD1.n123 12.0247
R2190 VDD1.n202 VDD1.n105 12.0247
R2191 VDD1.n96 VDD1.n95 11.249
R2192 VDD1.n64 VDD1.n18 11.249
R2193 VDD1.n51 VDD1.n28 11.249
R2194 VDD1.n152 VDD1.n129 11.249
R2195 VDD1.n167 VDD1.n121 11.249
R2196 VDD1.n199 VDD1.n198 11.249
R2197 VDD1.n36 VDD1.n35 10.7239
R2198 VDD1.n137 VDD1.n136 10.7239
R2199 VDD1.n92 VDD1.n4 10.4732
R2200 VDD1.n68 VDD1.n67 10.4732
R2201 VDD1.n48 VDD1.n47 10.4732
R2202 VDD1.n149 VDD1.n148 10.4732
R2203 VDD1.n171 VDD1.n170 10.4732
R2204 VDD1.n195 VDD1.n107 10.4732
R2205 VDD1.n91 VDD1.n6 9.69747
R2206 VDD1.n71 VDD1.n16 9.69747
R2207 VDD1.n44 VDD1.n30 9.69747
R2208 VDD1.n145 VDD1.n131 9.69747
R2209 VDD1.n174 VDD1.n119 9.69747
R2210 VDD1.n194 VDD1.n109 9.69747
R2211 VDD1.n98 VDD1.n0 9.45567
R2212 VDD1.n201 VDD1.n103 9.45567
R2213 VDD1.n99 VDD1.n98 9.3005
R2214 VDD1.n97 VDD1.n96 9.3005
R2215 VDD1.n4 VDD1.n3 9.3005
R2216 VDD1.n91 VDD1.n90 9.3005
R2217 VDD1.n89 VDD1.n88 9.3005
R2218 VDD1.n8 VDD1.n7 9.3005
R2219 VDD1.n83 VDD1.n82 9.3005
R2220 VDD1.n81 VDD1.n80 9.3005
R2221 VDD1.n12 VDD1.n11 9.3005
R2222 VDD1.n75 VDD1.n74 9.3005
R2223 VDD1.n73 VDD1.n72 9.3005
R2224 VDD1.n16 VDD1.n15 9.3005
R2225 VDD1.n67 VDD1.n66 9.3005
R2226 VDD1.n65 VDD1.n64 9.3005
R2227 VDD1.n20 VDD1.n19 9.3005
R2228 VDD1.n59 VDD1.n58 9.3005
R2229 VDD1.n57 VDD1.n56 9.3005
R2230 VDD1.n25 VDD1.n23 9.3005
R2231 VDD1.n51 VDD1.n50 9.3005
R2232 VDD1.n49 VDD1.n48 9.3005
R2233 VDD1.n30 VDD1.n29 9.3005
R2234 VDD1.n43 VDD1.n42 9.3005
R2235 VDD1.n41 VDD1.n40 9.3005
R2236 VDD1.n34 VDD1.n33 9.3005
R2237 VDD1.n184 VDD1.n183 9.3005
R2238 VDD1.n186 VDD1.n185 9.3005
R2239 VDD1.n111 VDD1.n110 9.3005
R2240 VDD1.n192 VDD1.n191 9.3005
R2241 VDD1.n194 VDD1.n193 9.3005
R2242 VDD1.n107 VDD1.n106 9.3005
R2243 VDD1.n200 VDD1.n199 9.3005
R2244 VDD1.n202 VDD1.n201 9.3005
R2245 VDD1.n178 VDD1.n177 9.3005
R2246 VDD1.n176 VDD1.n175 9.3005
R2247 VDD1.n119 VDD1.n118 9.3005
R2248 VDD1.n170 VDD1.n169 9.3005
R2249 VDD1.n168 VDD1.n167 9.3005
R2250 VDD1.n123 VDD1.n122 9.3005
R2251 VDD1.n162 VDD1.n161 9.3005
R2252 VDD1.n135 VDD1.n134 9.3005
R2253 VDD1.n142 VDD1.n141 9.3005
R2254 VDD1.n144 VDD1.n143 9.3005
R2255 VDD1.n131 VDD1.n130 9.3005
R2256 VDD1.n150 VDD1.n149 9.3005
R2257 VDD1.n152 VDD1.n151 9.3005
R2258 VDD1.n153 VDD1.n126 9.3005
R2259 VDD1.n160 VDD1.n159 9.3005
R2260 VDD1.n115 VDD1.n114 9.3005
R2261 VDD1.n88 VDD1.n87 8.92171
R2262 VDD1.n72 VDD1.n14 8.92171
R2263 VDD1.n43 VDD1.n32 8.92171
R2264 VDD1.n144 VDD1.n133 8.92171
R2265 VDD1.n175 VDD1.n117 8.92171
R2266 VDD1.n191 VDD1.n190 8.92171
R2267 VDD1.n84 VDD1.n8 8.14595
R2268 VDD1.n76 VDD1.n75 8.14595
R2269 VDD1.n40 VDD1.n39 8.14595
R2270 VDD1.n141 VDD1.n140 8.14595
R2271 VDD1.n179 VDD1.n178 8.14595
R2272 VDD1.n187 VDD1.n111 8.14595
R2273 VDD1.n83 VDD1.n10 7.3702
R2274 VDD1.n79 VDD1.n12 7.3702
R2275 VDD1.n36 VDD1.n34 7.3702
R2276 VDD1.n137 VDD1.n135 7.3702
R2277 VDD1.n182 VDD1.n115 7.3702
R2278 VDD1.n186 VDD1.n113 7.3702
R2279 VDD1.n80 VDD1.n10 6.59444
R2280 VDD1.n80 VDD1.n79 6.59444
R2281 VDD1.n183 VDD1.n182 6.59444
R2282 VDD1.n183 VDD1.n113 6.59444
R2283 VDD1.n84 VDD1.n83 5.81868
R2284 VDD1.n76 VDD1.n12 5.81868
R2285 VDD1.n39 VDD1.n34 5.81868
R2286 VDD1.n140 VDD1.n135 5.81868
R2287 VDD1.n179 VDD1.n115 5.81868
R2288 VDD1.n187 VDD1.n186 5.81868
R2289 VDD1.n87 VDD1.n8 5.04292
R2290 VDD1.n75 VDD1.n14 5.04292
R2291 VDD1.n40 VDD1.n32 5.04292
R2292 VDD1.n141 VDD1.n133 5.04292
R2293 VDD1.n178 VDD1.n117 5.04292
R2294 VDD1.n190 VDD1.n111 5.04292
R2295 VDD1.n88 VDD1.n6 4.26717
R2296 VDD1.n72 VDD1.n71 4.26717
R2297 VDD1.n44 VDD1.n43 4.26717
R2298 VDD1.n145 VDD1.n144 4.26717
R2299 VDD1.n175 VDD1.n174 4.26717
R2300 VDD1.n191 VDD1.n109 4.26717
R2301 VDD1.n92 VDD1.n91 3.49141
R2302 VDD1.n68 VDD1.n16 3.49141
R2303 VDD1.n47 VDD1.n30 3.49141
R2304 VDD1.n148 VDD1.n131 3.49141
R2305 VDD1.n171 VDD1.n119 3.49141
R2306 VDD1.n195 VDD1.n194 3.49141
R2307 VDD1.n95 VDD1.n4 2.71565
R2308 VDD1.n67 VDD1.n18 2.71565
R2309 VDD1.n48 VDD1.n28 2.71565
R2310 VDD1.n149 VDD1.n129 2.71565
R2311 VDD1.n170 VDD1.n121 2.71565
R2312 VDD1.n198 VDD1.n107 2.71565
R2313 VDD1.n35 VDD1.n33 2.41282
R2314 VDD1.n136 VDD1.n134 2.41282
R2315 VDD1.n96 VDD1.n2 1.93989
R2316 VDD1.n64 VDD1.n63 1.93989
R2317 VDD1.n52 VDD1.n51 1.93989
R2318 VDD1.n154 VDD1.n152 1.93989
R2319 VDD1.n167 VDD1.n166 1.93989
R2320 VDD1.n199 VDD1.n105 1.93989
R2321 VDD1.n100 VDD1.n99 1.16414
R2322 VDD1.n60 VDD1.n20 1.16414
R2323 VDD1.n55 VDD1.n25 1.16414
R2324 VDD1.n153 VDD1.n127 1.16414
R2325 VDD1.n163 VDD1.n123 1.16414
R2326 VDD1.n203 VDD1.n202 1.16414
R2327 VDD1.n102 VDD1.n0 0.388379
R2328 VDD1.n59 VDD1.n22 0.388379
R2329 VDD1.n56 VDD1.n24 0.388379
R2330 VDD1.n159 VDD1.n158 0.388379
R2331 VDD1.n162 VDD1.n125 0.388379
R2332 VDD1.n205 VDD1.n103 0.388379
R2333 VDD1.n98 VDD1.n97 0.155672
R2334 VDD1.n97 VDD1.n3 0.155672
R2335 VDD1.n90 VDD1.n3 0.155672
R2336 VDD1.n90 VDD1.n89 0.155672
R2337 VDD1.n89 VDD1.n7 0.155672
R2338 VDD1.n82 VDD1.n7 0.155672
R2339 VDD1.n82 VDD1.n81 0.155672
R2340 VDD1.n81 VDD1.n11 0.155672
R2341 VDD1.n74 VDD1.n11 0.155672
R2342 VDD1.n74 VDD1.n73 0.155672
R2343 VDD1.n73 VDD1.n15 0.155672
R2344 VDD1.n66 VDD1.n15 0.155672
R2345 VDD1.n66 VDD1.n65 0.155672
R2346 VDD1.n65 VDD1.n19 0.155672
R2347 VDD1.n58 VDD1.n19 0.155672
R2348 VDD1.n58 VDD1.n57 0.155672
R2349 VDD1.n57 VDD1.n23 0.155672
R2350 VDD1.n50 VDD1.n23 0.155672
R2351 VDD1.n50 VDD1.n49 0.155672
R2352 VDD1.n49 VDD1.n29 0.155672
R2353 VDD1.n42 VDD1.n29 0.155672
R2354 VDD1.n42 VDD1.n41 0.155672
R2355 VDD1.n41 VDD1.n33 0.155672
R2356 VDD1.n142 VDD1.n134 0.155672
R2357 VDD1.n143 VDD1.n142 0.155672
R2358 VDD1.n143 VDD1.n130 0.155672
R2359 VDD1.n150 VDD1.n130 0.155672
R2360 VDD1.n151 VDD1.n150 0.155672
R2361 VDD1.n151 VDD1.n126 0.155672
R2362 VDD1.n160 VDD1.n126 0.155672
R2363 VDD1.n161 VDD1.n160 0.155672
R2364 VDD1.n161 VDD1.n122 0.155672
R2365 VDD1.n168 VDD1.n122 0.155672
R2366 VDD1.n169 VDD1.n168 0.155672
R2367 VDD1.n169 VDD1.n118 0.155672
R2368 VDD1.n176 VDD1.n118 0.155672
R2369 VDD1.n177 VDD1.n176 0.155672
R2370 VDD1.n177 VDD1.n114 0.155672
R2371 VDD1.n184 VDD1.n114 0.155672
R2372 VDD1.n185 VDD1.n184 0.155672
R2373 VDD1.n185 VDD1.n110 0.155672
R2374 VDD1.n192 VDD1.n110 0.155672
R2375 VDD1.n193 VDD1.n192 0.155672
R2376 VDD1.n193 VDD1.n106 0.155672
R2377 VDD1.n200 VDD1.n106 0.155672
R2378 VDD1.n201 VDD1.n200 0.155672
C0 VN VDD2 4.16931f
C1 w_n2086_n4720# VDD2 2.26034f
C2 VN VP 6.6436f
C3 w_n2086_n4720# VP 3.26372f
C4 VTAIL VDD1 6.85241f
C5 VTAIL VDD2 6.90027f
C6 VTAIL VP 3.53201f
C7 VN B 1.10199f
C8 w_n2086_n4720# B 10.5533f
C9 VDD1 VDD2 0.658665f
C10 VP VDD1 4.34517f
C11 VTAIL B 5.09995f
C12 VP VDD2 0.32742f
C13 VN w_n2086_n4720# 2.99831f
C14 B VDD1 2.21857f
C15 B VDD2 2.24741f
C16 VN VTAIL 3.5176f
C17 VTAIL w_n2086_n4720# 3.72431f
C18 B VP 1.53778f
C19 VN VDD1 0.147724f
C20 w_n2086_n4720# VDD1 2.23613f
C21 VDD2 VSUBS 1.136696f
C22 VDD1 VSUBS 5.59969f
C23 VTAIL VSUBS 1.256024f
C24 VN VSUBS 9.20466f
C25 VP VSUBS 1.888048f
C26 B VSUBS 4.379263f
C27 w_n2086_n4720# VSUBS 0.120329p
C28 VDD1.n0 VSUBS 0.015677f
C29 VDD1.n1 VSUBS 0.035374f
C30 VDD1.n2 VSUBS 0.015846f
C31 VDD1.n3 VSUBS 0.027851f
C32 VDD1.n4 VSUBS 0.014966f
C33 VDD1.n5 VSUBS 0.035374f
C34 VDD1.n6 VSUBS 0.015846f
C35 VDD1.n7 VSUBS 0.027851f
C36 VDD1.n8 VSUBS 0.014966f
C37 VDD1.n9 VSUBS 0.035374f
C38 VDD1.n10 VSUBS 0.015846f
C39 VDD1.n11 VSUBS 0.027851f
C40 VDD1.n12 VSUBS 0.014966f
C41 VDD1.n13 VSUBS 0.035374f
C42 VDD1.n14 VSUBS 0.015846f
C43 VDD1.n15 VSUBS 0.027851f
C44 VDD1.n16 VSUBS 0.014966f
C45 VDD1.n17 VSUBS 0.035374f
C46 VDD1.n18 VSUBS 0.015846f
C47 VDD1.n19 VSUBS 0.027851f
C48 VDD1.n20 VSUBS 0.014966f
C49 VDD1.n21 VSUBS 0.035374f
C50 VDD1.n22 VSUBS 0.015406f
C51 VDD1.n23 VSUBS 0.027851f
C52 VDD1.n24 VSUBS 0.015406f
C53 VDD1.n25 VSUBS 0.014966f
C54 VDD1.n26 VSUBS 0.035374f
C55 VDD1.n27 VSUBS 0.035374f
C56 VDD1.n28 VSUBS 0.015846f
C57 VDD1.n29 VSUBS 0.027851f
C58 VDD1.n30 VSUBS 0.014966f
C59 VDD1.n31 VSUBS 0.035374f
C60 VDD1.n32 VSUBS 0.015846f
C61 VDD1.n33 VSUBS 2.19333f
C62 VDD1.n34 VSUBS 0.014966f
C63 VDD1.t1 VSUBS 0.076862f
C64 VDD1.n35 VSUBS 0.304468f
C65 VDD1.n36 VSUBS 0.02661f
C66 VDD1.n37 VSUBS 0.02653f
C67 VDD1.n38 VSUBS 0.035374f
C68 VDD1.n39 VSUBS 0.015846f
C69 VDD1.n40 VSUBS 0.014966f
C70 VDD1.n41 VSUBS 0.027851f
C71 VDD1.n42 VSUBS 0.027851f
C72 VDD1.n43 VSUBS 0.014966f
C73 VDD1.n44 VSUBS 0.015846f
C74 VDD1.n45 VSUBS 0.035374f
C75 VDD1.n46 VSUBS 0.035374f
C76 VDD1.n47 VSUBS 0.015846f
C77 VDD1.n48 VSUBS 0.014966f
C78 VDD1.n49 VSUBS 0.027851f
C79 VDD1.n50 VSUBS 0.027851f
C80 VDD1.n51 VSUBS 0.014966f
C81 VDD1.n52 VSUBS 0.015846f
C82 VDD1.n53 VSUBS 0.035374f
C83 VDD1.n54 VSUBS 0.035374f
C84 VDD1.n55 VSUBS 0.015846f
C85 VDD1.n56 VSUBS 0.014966f
C86 VDD1.n57 VSUBS 0.027851f
C87 VDD1.n58 VSUBS 0.027851f
C88 VDD1.n59 VSUBS 0.014966f
C89 VDD1.n60 VSUBS 0.015846f
C90 VDD1.n61 VSUBS 0.035374f
C91 VDD1.n62 VSUBS 0.035374f
C92 VDD1.n63 VSUBS 0.015846f
C93 VDD1.n64 VSUBS 0.014966f
C94 VDD1.n65 VSUBS 0.027851f
C95 VDD1.n66 VSUBS 0.027851f
C96 VDD1.n67 VSUBS 0.014966f
C97 VDD1.n68 VSUBS 0.015846f
C98 VDD1.n69 VSUBS 0.035374f
C99 VDD1.n70 VSUBS 0.035374f
C100 VDD1.n71 VSUBS 0.015846f
C101 VDD1.n72 VSUBS 0.014966f
C102 VDD1.n73 VSUBS 0.027851f
C103 VDD1.n74 VSUBS 0.027851f
C104 VDD1.n75 VSUBS 0.014966f
C105 VDD1.n76 VSUBS 0.015846f
C106 VDD1.n77 VSUBS 0.035374f
C107 VDD1.n78 VSUBS 0.035374f
C108 VDD1.n79 VSUBS 0.015846f
C109 VDD1.n80 VSUBS 0.014966f
C110 VDD1.n81 VSUBS 0.027851f
C111 VDD1.n82 VSUBS 0.027851f
C112 VDD1.n83 VSUBS 0.014966f
C113 VDD1.n84 VSUBS 0.015846f
C114 VDD1.n85 VSUBS 0.035374f
C115 VDD1.n86 VSUBS 0.035374f
C116 VDD1.n87 VSUBS 0.015846f
C117 VDD1.n88 VSUBS 0.014966f
C118 VDD1.n89 VSUBS 0.027851f
C119 VDD1.n90 VSUBS 0.027851f
C120 VDD1.n91 VSUBS 0.014966f
C121 VDD1.n92 VSUBS 0.015846f
C122 VDD1.n93 VSUBS 0.035374f
C123 VDD1.n94 VSUBS 0.035374f
C124 VDD1.n95 VSUBS 0.015846f
C125 VDD1.n96 VSUBS 0.014966f
C126 VDD1.n97 VSUBS 0.027851f
C127 VDD1.n98 VSUBS 0.070463f
C128 VDD1.n99 VSUBS 0.014966f
C129 VDD1.n100 VSUBS 0.015846f
C130 VDD1.n101 VSUBS 0.078805f
C131 VDD1.n102 VSUBS 0.072632f
C132 VDD1.n103 VSUBS 0.015677f
C133 VDD1.n104 VSUBS 0.035374f
C134 VDD1.n105 VSUBS 0.015846f
C135 VDD1.n106 VSUBS 0.027851f
C136 VDD1.n107 VSUBS 0.014966f
C137 VDD1.n108 VSUBS 0.035374f
C138 VDD1.n109 VSUBS 0.015846f
C139 VDD1.n110 VSUBS 0.027851f
C140 VDD1.n111 VSUBS 0.014966f
C141 VDD1.n112 VSUBS 0.035374f
C142 VDD1.n113 VSUBS 0.015846f
C143 VDD1.n114 VSUBS 0.027851f
C144 VDD1.n115 VSUBS 0.014966f
C145 VDD1.n116 VSUBS 0.035374f
C146 VDD1.n117 VSUBS 0.015846f
C147 VDD1.n118 VSUBS 0.027851f
C148 VDD1.n119 VSUBS 0.014966f
C149 VDD1.n120 VSUBS 0.035374f
C150 VDD1.n121 VSUBS 0.015846f
C151 VDD1.n122 VSUBS 0.027851f
C152 VDD1.n123 VSUBS 0.014966f
C153 VDD1.n124 VSUBS 0.035374f
C154 VDD1.n125 VSUBS 0.015406f
C155 VDD1.n126 VSUBS 0.027851f
C156 VDD1.n127 VSUBS 0.015846f
C157 VDD1.n128 VSUBS 0.035374f
C158 VDD1.n129 VSUBS 0.015846f
C159 VDD1.n130 VSUBS 0.027851f
C160 VDD1.n131 VSUBS 0.014966f
C161 VDD1.n132 VSUBS 0.035374f
C162 VDD1.n133 VSUBS 0.015846f
C163 VDD1.n134 VSUBS 2.19333f
C164 VDD1.n135 VSUBS 0.014966f
C165 VDD1.t0 VSUBS 0.076862f
C166 VDD1.n136 VSUBS 0.304468f
C167 VDD1.n137 VSUBS 0.02661f
C168 VDD1.n138 VSUBS 0.02653f
C169 VDD1.n139 VSUBS 0.035374f
C170 VDD1.n140 VSUBS 0.015846f
C171 VDD1.n141 VSUBS 0.014966f
C172 VDD1.n142 VSUBS 0.027851f
C173 VDD1.n143 VSUBS 0.027851f
C174 VDD1.n144 VSUBS 0.014966f
C175 VDD1.n145 VSUBS 0.015846f
C176 VDD1.n146 VSUBS 0.035374f
C177 VDD1.n147 VSUBS 0.035374f
C178 VDD1.n148 VSUBS 0.015846f
C179 VDD1.n149 VSUBS 0.014966f
C180 VDD1.n150 VSUBS 0.027851f
C181 VDD1.n151 VSUBS 0.027851f
C182 VDD1.n152 VSUBS 0.014966f
C183 VDD1.n153 VSUBS 0.014966f
C184 VDD1.n154 VSUBS 0.015846f
C185 VDD1.n155 VSUBS 0.035374f
C186 VDD1.n156 VSUBS 0.035374f
C187 VDD1.n157 VSUBS 0.035374f
C188 VDD1.n158 VSUBS 0.015406f
C189 VDD1.n159 VSUBS 0.014966f
C190 VDD1.n160 VSUBS 0.027851f
C191 VDD1.n161 VSUBS 0.027851f
C192 VDD1.n162 VSUBS 0.014966f
C193 VDD1.n163 VSUBS 0.015846f
C194 VDD1.n164 VSUBS 0.035374f
C195 VDD1.n165 VSUBS 0.035374f
C196 VDD1.n166 VSUBS 0.015846f
C197 VDD1.n167 VSUBS 0.014966f
C198 VDD1.n168 VSUBS 0.027851f
C199 VDD1.n169 VSUBS 0.027851f
C200 VDD1.n170 VSUBS 0.014966f
C201 VDD1.n171 VSUBS 0.015846f
C202 VDD1.n172 VSUBS 0.035374f
C203 VDD1.n173 VSUBS 0.035374f
C204 VDD1.n174 VSUBS 0.015846f
C205 VDD1.n175 VSUBS 0.014966f
C206 VDD1.n176 VSUBS 0.027851f
C207 VDD1.n177 VSUBS 0.027851f
C208 VDD1.n178 VSUBS 0.014966f
C209 VDD1.n179 VSUBS 0.015846f
C210 VDD1.n180 VSUBS 0.035374f
C211 VDD1.n181 VSUBS 0.035374f
C212 VDD1.n182 VSUBS 0.015846f
C213 VDD1.n183 VSUBS 0.014966f
C214 VDD1.n184 VSUBS 0.027851f
C215 VDD1.n185 VSUBS 0.027851f
C216 VDD1.n186 VSUBS 0.014966f
C217 VDD1.n187 VSUBS 0.015846f
C218 VDD1.n188 VSUBS 0.035374f
C219 VDD1.n189 VSUBS 0.035374f
C220 VDD1.n190 VSUBS 0.015846f
C221 VDD1.n191 VSUBS 0.014966f
C222 VDD1.n192 VSUBS 0.027851f
C223 VDD1.n193 VSUBS 0.027851f
C224 VDD1.n194 VSUBS 0.014966f
C225 VDD1.n195 VSUBS 0.015846f
C226 VDD1.n196 VSUBS 0.035374f
C227 VDD1.n197 VSUBS 0.035374f
C228 VDD1.n198 VSUBS 0.015846f
C229 VDD1.n199 VSUBS 0.014966f
C230 VDD1.n200 VSUBS 0.027851f
C231 VDD1.n201 VSUBS 0.070463f
C232 VDD1.n202 VSUBS 0.014966f
C233 VDD1.n203 VSUBS 0.015846f
C234 VDD1.n204 VSUBS 0.078805f
C235 VDD1.n205 VSUBS 1.12975f
C236 VP.t0 VSUBS 5.81688f
C237 VP.t1 VSUBS 5.17637f
C238 VP.n0 VSUBS 6.62148f
C239 B.n0 VSUBS 0.006109f
C240 B.n1 VSUBS 0.006109f
C241 B.n2 VSUBS 0.009034f
C242 B.n3 VSUBS 0.006923f
C243 B.n4 VSUBS 0.006923f
C244 B.n5 VSUBS 0.006923f
C245 B.n6 VSUBS 0.006923f
C246 B.n7 VSUBS 0.006923f
C247 B.n8 VSUBS 0.006923f
C248 B.n9 VSUBS 0.006923f
C249 B.n10 VSUBS 0.006923f
C250 B.n11 VSUBS 0.006923f
C251 B.n12 VSUBS 0.006923f
C252 B.n13 VSUBS 0.006923f
C253 B.n14 VSUBS 0.016064f
C254 B.n15 VSUBS 0.006923f
C255 B.n16 VSUBS 0.006923f
C256 B.n17 VSUBS 0.006923f
C257 B.n18 VSUBS 0.006923f
C258 B.n19 VSUBS 0.006923f
C259 B.n20 VSUBS 0.006923f
C260 B.n21 VSUBS 0.006923f
C261 B.n22 VSUBS 0.006923f
C262 B.n23 VSUBS 0.006923f
C263 B.n24 VSUBS 0.006923f
C264 B.n25 VSUBS 0.006923f
C265 B.n26 VSUBS 0.006923f
C266 B.n27 VSUBS 0.006923f
C267 B.n28 VSUBS 0.006923f
C268 B.n29 VSUBS 0.006923f
C269 B.n30 VSUBS 0.006923f
C270 B.n31 VSUBS 0.006923f
C271 B.n32 VSUBS 0.006923f
C272 B.n33 VSUBS 0.006923f
C273 B.n34 VSUBS 0.006923f
C274 B.n35 VSUBS 0.006923f
C275 B.n36 VSUBS 0.006923f
C276 B.n37 VSUBS 0.006923f
C277 B.n38 VSUBS 0.006923f
C278 B.n39 VSUBS 0.006923f
C279 B.n40 VSUBS 0.006923f
C280 B.n41 VSUBS 0.006923f
C281 B.n42 VSUBS 0.006923f
C282 B.n43 VSUBS 0.006923f
C283 B.n44 VSUBS 0.006923f
C284 B.n45 VSUBS 0.006923f
C285 B.t1 VSUBS 0.365297f
C286 B.t2 VSUBS 0.39707f
C287 B.t0 VSUBS 2.01051f
C288 B.n46 VSUBS 0.601688f
C289 B.n47 VSUBS 0.333624f
C290 B.n48 VSUBS 0.006923f
C291 B.n49 VSUBS 0.006923f
C292 B.n50 VSUBS 0.006923f
C293 B.n51 VSUBS 0.006923f
C294 B.t4 VSUBS 0.3653f
C295 B.t5 VSUBS 0.397073f
C296 B.t3 VSUBS 2.01051f
C297 B.n52 VSUBS 0.601685f
C298 B.n53 VSUBS 0.33362f
C299 B.n54 VSUBS 0.006923f
C300 B.n55 VSUBS 0.006923f
C301 B.n56 VSUBS 0.006923f
C302 B.n57 VSUBS 0.006923f
C303 B.n58 VSUBS 0.006923f
C304 B.n59 VSUBS 0.006923f
C305 B.n60 VSUBS 0.006923f
C306 B.n61 VSUBS 0.006923f
C307 B.n62 VSUBS 0.006923f
C308 B.n63 VSUBS 0.006923f
C309 B.n64 VSUBS 0.006923f
C310 B.n65 VSUBS 0.006923f
C311 B.n66 VSUBS 0.006923f
C312 B.n67 VSUBS 0.006923f
C313 B.n68 VSUBS 0.006923f
C314 B.n69 VSUBS 0.006923f
C315 B.n70 VSUBS 0.006923f
C316 B.n71 VSUBS 0.006923f
C317 B.n72 VSUBS 0.006923f
C318 B.n73 VSUBS 0.006923f
C319 B.n74 VSUBS 0.006923f
C320 B.n75 VSUBS 0.006923f
C321 B.n76 VSUBS 0.006923f
C322 B.n77 VSUBS 0.006923f
C323 B.n78 VSUBS 0.006923f
C324 B.n79 VSUBS 0.006923f
C325 B.n80 VSUBS 0.006923f
C326 B.n81 VSUBS 0.006923f
C327 B.n82 VSUBS 0.006923f
C328 B.n83 VSUBS 0.006923f
C329 B.n84 VSUBS 0.016064f
C330 B.n85 VSUBS 0.006923f
C331 B.n86 VSUBS 0.006923f
C332 B.n87 VSUBS 0.006923f
C333 B.n88 VSUBS 0.006923f
C334 B.n89 VSUBS 0.006923f
C335 B.n90 VSUBS 0.006923f
C336 B.n91 VSUBS 0.006923f
C337 B.n92 VSUBS 0.006923f
C338 B.n93 VSUBS 0.006923f
C339 B.n94 VSUBS 0.006923f
C340 B.n95 VSUBS 0.006923f
C341 B.n96 VSUBS 0.006923f
C342 B.n97 VSUBS 0.006923f
C343 B.n98 VSUBS 0.006923f
C344 B.n99 VSUBS 0.006923f
C345 B.n100 VSUBS 0.006923f
C346 B.n101 VSUBS 0.006923f
C347 B.n102 VSUBS 0.006923f
C348 B.n103 VSUBS 0.006923f
C349 B.n104 VSUBS 0.006923f
C350 B.n105 VSUBS 0.006923f
C351 B.n106 VSUBS 0.006923f
C352 B.n107 VSUBS 0.006923f
C353 B.n108 VSUBS 0.006923f
C354 B.n109 VSUBS 0.014886f
C355 B.n110 VSUBS 0.006923f
C356 B.n111 VSUBS 0.006923f
C357 B.n112 VSUBS 0.006923f
C358 B.n113 VSUBS 0.006923f
C359 B.n114 VSUBS 0.006923f
C360 B.n115 VSUBS 0.006923f
C361 B.n116 VSUBS 0.006923f
C362 B.n117 VSUBS 0.006923f
C363 B.n118 VSUBS 0.006923f
C364 B.n119 VSUBS 0.006923f
C365 B.n120 VSUBS 0.006923f
C366 B.n121 VSUBS 0.006923f
C367 B.n122 VSUBS 0.006923f
C368 B.n123 VSUBS 0.006923f
C369 B.n124 VSUBS 0.006923f
C370 B.n125 VSUBS 0.006923f
C371 B.n126 VSUBS 0.006923f
C372 B.n127 VSUBS 0.006923f
C373 B.n128 VSUBS 0.006923f
C374 B.n129 VSUBS 0.006923f
C375 B.n130 VSUBS 0.006923f
C376 B.n131 VSUBS 0.006923f
C377 B.n132 VSUBS 0.006923f
C378 B.n133 VSUBS 0.006923f
C379 B.n134 VSUBS 0.006923f
C380 B.n135 VSUBS 0.006923f
C381 B.n136 VSUBS 0.006923f
C382 B.n137 VSUBS 0.006923f
C383 B.n138 VSUBS 0.006923f
C384 B.n139 VSUBS 0.006923f
C385 B.n140 VSUBS 0.004785f
C386 B.n141 VSUBS 0.006923f
C387 B.n142 VSUBS 0.006923f
C388 B.n143 VSUBS 0.006923f
C389 B.n144 VSUBS 0.006923f
C390 B.n145 VSUBS 0.006923f
C391 B.t8 VSUBS 0.365297f
C392 B.t7 VSUBS 0.39707f
C393 B.t6 VSUBS 2.01051f
C394 B.n146 VSUBS 0.601688f
C395 B.n147 VSUBS 0.333624f
C396 B.n148 VSUBS 0.006923f
C397 B.n149 VSUBS 0.006923f
C398 B.n150 VSUBS 0.006923f
C399 B.n151 VSUBS 0.006923f
C400 B.n152 VSUBS 0.006923f
C401 B.n153 VSUBS 0.006923f
C402 B.n154 VSUBS 0.006923f
C403 B.n155 VSUBS 0.006923f
C404 B.n156 VSUBS 0.006923f
C405 B.n157 VSUBS 0.006923f
C406 B.n158 VSUBS 0.006923f
C407 B.n159 VSUBS 0.006923f
C408 B.n160 VSUBS 0.006923f
C409 B.n161 VSUBS 0.006923f
C410 B.n162 VSUBS 0.006923f
C411 B.n163 VSUBS 0.006923f
C412 B.n164 VSUBS 0.006923f
C413 B.n165 VSUBS 0.006923f
C414 B.n166 VSUBS 0.006923f
C415 B.n167 VSUBS 0.006923f
C416 B.n168 VSUBS 0.006923f
C417 B.n169 VSUBS 0.006923f
C418 B.n170 VSUBS 0.006923f
C419 B.n171 VSUBS 0.006923f
C420 B.n172 VSUBS 0.006923f
C421 B.n173 VSUBS 0.006923f
C422 B.n174 VSUBS 0.006923f
C423 B.n175 VSUBS 0.006923f
C424 B.n176 VSUBS 0.006923f
C425 B.n177 VSUBS 0.006923f
C426 B.n178 VSUBS 0.014886f
C427 B.n179 VSUBS 0.006923f
C428 B.n180 VSUBS 0.006923f
C429 B.n181 VSUBS 0.006923f
C430 B.n182 VSUBS 0.006923f
C431 B.n183 VSUBS 0.006923f
C432 B.n184 VSUBS 0.006923f
C433 B.n185 VSUBS 0.006923f
C434 B.n186 VSUBS 0.006923f
C435 B.n187 VSUBS 0.006923f
C436 B.n188 VSUBS 0.006923f
C437 B.n189 VSUBS 0.006923f
C438 B.n190 VSUBS 0.006923f
C439 B.n191 VSUBS 0.006923f
C440 B.n192 VSUBS 0.006923f
C441 B.n193 VSUBS 0.006923f
C442 B.n194 VSUBS 0.006923f
C443 B.n195 VSUBS 0.006923f
C444 B.n196 VSUBS 0.006923f
C445 B.n197 VSUBS 0.006923f
C446 B.n198 VSUBS 0.006923f
C447 B.n199 VSUBS 0.006923f
C448 B.n200 VSUBS 0.006923f
C449 B.n201 VSUBS 0.006923f
C450 B.n202 VSUBS 0.006923f
C451 B.n203 VSUBS 0.006923f
C452 B.n204 VSUBS 0.006923f
C453 B.n205 VSUBS 0.006923f
C454 B.n206 VSUBS 0.006923f
C455 B.n207 VSUBS 0.006923f
C456 B.n208 VSUBS 0.006923f
C457 B.n209 VSUBS 0.006923f
C458 B.n210 VSUBS 0.006923f
C459 B.n211 VSUBS 0.006923f
C460 B.n212 VSUBS 0.006923f
C461 B.n213 VSUBS 0.006923f
C462 B.n214 VSUBS 0.006923f
C463 B.n215 VSUBS 0.006923f
C464 B.n216 VSUBS 0.006923f
C465 B.n217 VSUBS 0.006923f
C466 B.n218 VSUBS 0.006923f
C467 B.n219 VSUBS 0.006923f
C468 B.n220 VSUBS 0.006923f
C469 B.n221 VSUBS 0.006923f
C470 B.n222 VSUBS 0.006923f
C471 B.n223 VSUBS 0.014886f
C472 B.n224 VSUBS 0.016064f
C473 B.n225 VSUBS 0.016064f
C474 B.n226 VSUBS 0.006923f
C475 B.n227 VSUBS 0.006923f
C476 B.n228 VSUBS 0.006923f
C477 B.n229 VSUBS 0.006923f
C478 B.n230 VSUBS 0.006923f
C479 B.n231 VSUBS 0.006923f
C480 B.n232 VSUBS 0.006923f
C481 B.n233 VSUBS 0.006923f
C482 B.n234 VSUBS 0.006923f
C483 B.n235 VSUBS 0.006923f
C484 B.n236 VSUBS 0.006923f
C485 B.n237 VSUBS 0.006923f
C486 B.n238 VSUBS 0.006923f
C487 B.n239 VSUBS 0.006923f
C488 B.n240 VSUBS 0.006923f
C489 B.n241 VSUBS 0.006923f
C490 B.n242 VSUBS 0.006923f
C491 B.n243 VSUBS 0.006923f
C492 B.n244 VSUBS 0.006923f
C493 B.n245 VSUBS 0.006923f
C494 B.n246 VSUBS 0.006923f
C495 B.n247 VSUBS 0.006923f
C496 B.n248 VSUBS 0.006923f
C497 B.n249 VSUBS 0.006923f
C498 B.n250 VSUBS 0.006923f
C499 B.n251 VSUBS 0.006923f
C500 B.n252 VSUBS 0.006923f
C501 B.n253 VSUBS 0.006923f
C502 B.n254 VSUBS 0.006923f
C503 B.n255 VSUBS 0.006923f
C504 B.n256 VSUBS 0.006923f
C505 B.n257 VSUBS 0.006923f
C506 B.n258 VSUBS 0.006923f
C507 B.n259 VSUBS 0.006923f
C508 B.n260 VSUBS 0.006923f
C509 B.n261 VSUBS 0.006923f
C510 B.n262 VSUBS 0.006923f
C511 B.n263 VSUBS 0.006923f
C512 B.n264 VSUBS 0.006923f
C513 B.n265 VSUBS 0.006923f
C514 B.n266 VSUBS 0.006923f
C515 B.n267 VSUBS 0.006923f
C516 B.n268 VSUBS 0.006923f
C517 B.n269 VSUBS 0.006923f
C518 B.n270 VSUBS 0.006923f
C519 B.n271 VSUBS 0.006923f
C520 B.n272 VSUBS 0.006923f
C521 B.n273 VSUBS 0.006923f
C522 B.n274 VSUBS 0.006923f
C523 B.n275 VSUBS 0.006923f
C524 B.n276 VSUBS 0.006923f
C525 B.n277 VSUBS 0.006923f
C526 B.n278 VSUBS 0.006923f
C527 B.n279 VSUBS 0.006923f
C528 B.n280 VSUBS 0.006923f
C529 B.n281 VSUBS 0.006923f
C530 B.n282 VSUBS 0.006923f
C531 B.n283 VSUBS 0.006923f
C532 B.n284 VSUBS 0.006923f
C533 B.n285 VSUBS 0.006923f
C534 B.n286 VSUBS 0.006923f
C535 B.n287 VSUBS 0.006923f
C536 B.n288 VSUBS 0.006923f
C537 B.n289 VSUBS 0.006923f
C538 B.n290 VSUBS 0.006923f
C539 B.n291 VSUBS 0.006923f
C540 B.n292 VSUBS 0.006923f
C541 B.n293 VSUBS 0.006923f
C542 B.n294 VSUBS 0.006923f
C543 B.n295 VSUBS 0.006923f
C544 B.n296 VSUBS 0.006923f
C545 B.n297 VSUBS 0.006923f
C546 B.n298 VSUBS 0.006923f
C547 B.n299 VSUBS 0.006923f
C548 B.n300 VSUBS 0.006923f
C549 B.n301 VSUBS 0.006923f
C550 B.n302 VSUBS 0.006923f
C551 B.n303 VSUBS 0.006923f
C552 B.n304 VSUBS 0.006923f
C553 B.n305 VSUBS 0.006923f
C554 B.n306 VSUBS 0.006923f
C555 B.n307 VSUBS 0.006923f
C556 B.n308 VSUBS 0.006923f
C557 B.n309 VSUBS 0.006923f
C558 B.n310 VSUBS 0.006923f
C559 B.n311 VSUBS 0.006923f
C560 B.n312 VSUBS 0.006923f
C561 B.n313 VSUBS 0.006923f
C562 B.n314 VSUBS 0.006923f
C563 B.n315 VSUBS 0.006923f
C564 B.n316 VSUBS 0.004785f
C565 B.n317 VSUBS 0.01604f
C566 B.n318 VSUBS 0.0056f
C567 B.n319 VSUBS 0.006923f
C568 B.n320 VSUBS 0.006923f
C569 B.n321 VSUBS 0.006923f
C570 B.n322 VSUBS 0.006923f
C571 B.n323 VSUBS 0.006923f
C572 B.n324 VSUBS 0.006923f
C573 B.n325 VSUBS 0.006923f
C574 B.n326 VSUBS 0.006923f
C575 B.n327 VSUBS 0.006923f
C576 B.n328 VSUBS 0.006923f
C577 B.n329 VSUBS 0.006923f
C578 B.t11 VSUBS 0.3653f
C579 B.t10 VSUBS 0.397073f
C580 B.t9 VSUBS 2.01051f
C581 B.n330 VSUBS 0.601685f
C582 B.n331 VSUBS 0.33362f
C583 B.n332 VSUBS 0.01604f
C584 B.n333 VSUBS 0.0056f
C585 B.n334 VSUBS 0.006923f
C586 B.n335 VSUBS 0.006923f
C587 B.n336 VSUBS 0.006923f
C588 B.n337 VSUBS 0.006923f
C589 B.n338 VSUBS 0.006923f
C590 B.n339 VSUBS 0.006923f
C591 B.n340 VSUBS 0.006923f
C592 B.n341 VSUBS 0.006923f
C593 B.n342 VSUBS 0.006923f
C594 B.n343 VSUBS 0.006923f
C595 B.n344 VSUBS 0.006923f
C596 B.n345 VSUBS 0.006923f
C597 B.n346 VSUBS 0.006923f
C598 B.n347 VSUBS 0.006923f
C599 B.n348 VSUBS 0.006923f
C600 B.n349 VSUBS 0.006923f
C601 B.n350 VSUBS 0.006923f
C602 B.n351 VSUBS 0.006923f
C603 B.n352 VSUBS 0.006923f
C604 B.n353 VSUBS 0.006923f
C605 B.n354 VSUBS 0.006923f
C606 B.n355 VSUBS 0.006923f
C607 B.n356 VSUBS 0.006923f
C608 B.n357 VSUBS 0.006923f
C609 B.n358 VSUBS 0.006923f
C610 B.n359 VSUBS 0.006923f
C611 B.n360 VSUBS 0.006923f
C612 B.n361 VSUBS 0.006923f
C613 B.n362 VSUBS 0.006923f
C614 B.n363 VSUBS 0.006923f
C615 B.n364 VSUBS 0.006923f
C616 B.n365 VSUBS 0.006923f
C617 B.n366 VSUBS 0.006923f
C618 B.n367 VSUBS 0.006923f
C619 B.n368 VSUBS 0.006923f
C620 B.n369 VSUBS 0.006923f
C621 B.n370 VSUBS 0.006923f
C622 B.n371 VSUBS 0.006923f
C623 B.n372 VSUBS 0.006923f
C624 B.n373 VSUBS 0.006923f
C625 B.n374 VSUBS 0.006923f
C626 B.n375 VSUBS 0.006923f
C627 B.n376 VSUBS 0.006923f
C628 B.n377 VSUBS 0.006923f
C629 B.n378 VSUBS 0.006923f
C630 B.n379 VSUBS 0.006923f
C631 B.n380 VSUBS 0.006923f
C632 B.n381 VSUBS 0.006923f
C633 B.n382 VSUBS 0.006923f
C634 B.n383 VSUBS 0.006923f
C635 B.n384 VSUBS 0.006923f
C636 B.n385 VSUBS 0.006923f
C637 B.n386 VSUBS 0.006923f
C638 B.n387 VSUBS 0.006923f
C639 B.n388 VSUBS 0.006923f
C640 B.n389 VSUBS 0.006923f
C641 B.n390 VSUBS 0.006923f
C642 B.n391 VSUBS 0.006923f
C643 B.n392 VSUBS 0.006923f
C644 B.n393 VSUBS 0.006923f
C645 B.n394 VSUBS 0.006923f
C646 B.n395 VSUBS 0.006923f
C647 B.n396 VSUBS 0.006923f
C648 B.n397 VSUBS 0.006923f
C649 B.n398 VSUBS 0.006923f
C650 B.n399 VSUBS 0.006923f
C651 B.n400 VSUBS 0.006923f
C652 B.n401 VSUBS 0.006923f
C653 B.n402 VSUBS 0.006923f
C654 B.n403 VSUBS 0.006923f
C655 B.n404 VSUBS 0.006923f
C656 B.n405 VSUBS 0.006923f
C657 B.n406 VSUBS 0.006923f
C658 B.n407 VSUBS 0.006923f
C659 B.n408 VSUBS 0.006923f
C660 B.n409 VSUBS 0.006923f
C661 B.n410 VSUBS 0.006923f
C662 B.n411 VSUBS 0.006923f
C663 B.n412 VSUBS 0.006923f
C664 B.n413 VSUBS 0.006923f
C665 B.n414 VSUBS 0.006923f
C666 B.n415 VSUBS 0.006923f
C667 B.n416 VSUBS 0.006923f
C668 B.n417 VSUBS 0.006923f
C669 B.n418 VSUBS 0.006923f
C670 B.n419 VSUBS 0.006923f
C671 B.n420 VSUBS 0.006923f
C672 B.n421 VSUBS 0.006923f
C673 B.n422 VSUBS 0.006923f
C674 B.n423 VSUBS 0.006923f
C675 B.n424 VSUBS 0.006923f
C676 B.n425 VSUBS 0.006923f
C677 B.n426 VSUBS 0.016064f
C678 B.n427 VSUBS 0.015186f
C679 B.n428 VSUBS 0.015764f
C680 B.n429 VSUBS 0.006923f
C681 B.n430 VSUBS 0.006923f
C682 B.n431 VSUBS 0.006923f
C683 B.n432 VSUBS 0.006923f
C684 B.n433 VSUBS 0.006923f
C685 B.n434 VSUBS 0.006923f
C686 B.n435 VSUBS 0.006923f
C687 B.n436 VSUBS 0.006923f
C688 B.n437 VSUBS 0.006923f
C689 B.n438 VSUBS 0.006923f
C690 B.n439 VSUBS 0.006923f
C691 B.n440 VSUBS 0.006923f
C692 B.n441 VSUBS 0.006923f
C693 B.n442 VSUBS 0.006923f
C694 B.n443 VSUBS 0.006923f
C695 B.n444 VSUBS 0.006923f
C696 B.n445 VSUBS 0.006923f
C697 B.n446 VSUBS 0.006923f
C698 B.n447 VSUBS 0.006923f
C699 B.n448 VSUBS 0.006923f
C700 B.n449 VSUBS 0.006923f
C701 B.n450 VSUBS 0.006923f
C702 B.n451 VSUBS 0.006923f
C703 B.n452 VSUBS 0.006923f
C704 B.n453 VSUBS 0.006923f
C705 B.n454 VSUBS 0.006923f
C706 B.n455 VSUBS 0.006923f
C707 B.n456 VSUBS 0.006923f
C708 B.n457 VSUBS 0.006923f
C709 B.n458 VSUBS 0.006923f
C710 B.n459 VSUBS 0.006923f
C711 B.n460 VSUBS 0.006923f
C712 B.n461 VSUBS 0.006923f
C713 B.n462 VSUBS 0.006923f
C714 B.n463 VSUBS 0.006923f
C715 B.n464 VSUBS 0.006923f
C716 B.n465 VSUBS 0.006923f
C717 B.n466 VSUBS 0.006923f
C718 B.n467 VSUBS 0.006923f
C719 B.n468 VSUBS 0.006923f
C720 B.n469 VSUBS 0.006923f
C721 B.n470 VSUBS 0.006923f
C722 B.n471 VSUBS 0.006923f
C723 B.n472 VSUBS 0.006923f
C724 B.n473 VSUBS 0.006923f
C725 B.n474 VSUBS 0.006923f
C726 B.n475 VSUBS 0.006923f
C727 B.n476 VSUBS 0.006923f
C728 B.n477 VSUBS 0.006923f
C729 B.n478 VSUBS 0.006923f
C730 B.n479 VSUBS 0.006923f
C731 B.n480 VSUBS 0.006923f
C732 B.n481 VSUBS 0.006923f
C733 B.n482 VSUBS 0.006923f
C734 B.n483 VSUBS 0.006923f
C735 B.n484 VSUBS 0.006923f
C736 B.n485 VSUBS 0.006923f
C737 B.n486 VSUBS 0.006923f
C738 B.n487 VSUBS 0.006923f
C739 B.n488 VSUBS 0.006923f
C740 B.n489 VSUBS 0.006923f
C741 B.n490 VSUBS 0.006923f
C742 B.n491 VSUBS 0.006923f
C743 B.n492 VSUBS 0.006923f
C744 B.n493 VSUBS 0.006923f
C745 B.n494 VSUBS 0.006923f
C746 B.n495 VSUBS 0.006923f
C747 B.n496 VSUBS 0.006923f
C748 B.n497 VSUBS 0.006923f
C749 B.n498 VSUBS 0.006923f
C750 B.n499 VSUBS 0.006923f
C751 B.n500 VSUBS 0.006923f
C752 B.n501 VSUBS 0.014886f
C753 B.n502 VSUBS 0.014886f
C754 B.n503 VSUBS 0.016064f
C755 B.n504 VSUBS 0.006923f
C756 B.n505 VSUBS 0.006923f
C757 B.n506 VSUBS 0.006923f
C758 B.n507 VSUBS 0.006923f
C759 B.n508 VSUBS 0.006923f
C760 B.n509 VSUBS 0.006923f
C761 B.n510 VSUBS 0.006923f
C762 B.n511 VSUBS 0.006923f
C763 B.n512 VSUBS 0.006923f
C764 B.n513 VSUBS 0.006923f
C765 B.n514 VSUBS 0.006923f
C766 B.n515 VSUBS 0.006923f
C767 B.n516 VSUBS 0.006923f
C768 B.n517 VSUBS 0.006923f
C769 B.n518 VSUBS 0.006923f
C770 B.n519 VSUBS 0.006923f
C771 B.n520 VSUBS 0.006923f
C772 B.n521 VSUBS 0.006923f
C773 B.n522 VSUBS 0.006923f
C774 B.n523 VSUBS 0.006923f
C775 B.n524 VSUBS 0.006923f
C776 B.n525 VSUBS 0.006923f
C777 B.n526 VSUBS 0.006923f
C778 B.n527 VSUBS 0.006923f
C779 B.n528 VSUBS 0.006923f
C780 B.n529 VSUBS 0.006923f
C781 B.n530 VSUBS 0.006923f
C782 B.n531 VSUBS 0.006923f
C783 B.n532 VSUBS 0.006923f
C784 B.n533 VSUBS 0.006923f
C785 B.n534 VSUBS 0.006923f
C786 B.n535 VSUBS 0.006923f
C787 B.n536 VSUBS 0.006923f
C788 B.n537 VSUBS 0.006923f
C789 B.n538 VSUBS 0.006923f
C790 B.n539 VSUBS 0.006923f
C791 B.n540 VSUBS 0.006923f
C792 B.n541 VSUBS 0.006923f
C793 B.n542 VSUBS 0.006923f
C794 B.n543 VSUBS 0.006923f
C795 B.n544 VSUBS 0.006923f
C796 B.n545 VSUBS 0.006923f
C797 B.n546 VSUBS 0.006923f
C798 B.n547 VSUBS 0.006923f
C799 B.n548 VSUBS 0.006923f
C800 B.n549 VSUBS 0.006923f
C801 B.n550 VSUBS 0.006923f
C802 B.n551 VSUBS 0.006923f
C803 B.n552 VSUBS 0.006923f
C804 B.n553 VSUBS 0.006923f
C805 B.n554 VSUBS 0.006923f
C806 B.n555 VSUBS 0.006923f
C807 B.n556 VSUBS 0.006923f
C808 B.n557 VSUBS 0.006923f
C809 B.n558 VSUBS 0.006923f
C810 B.n559 VSUBS 0.006923f
C811 B.n560 VSUBS 0.006923f
C812 B.n561 VSUBS 0.006923f
C813 B.n562 VSUBS 0.006923f
C814 B.n563 VSUBS 0.006923f
C815 B.n564 VSUBS 0.006923f
C816 B.n565 VSUBS 0.006923f
C817 B.n566 VSUBS 0.006923f
C818 B.n567 VSUBS 0.006923f
C819 B.n568 VSUBS 0.006923f
C820 B.n569 VSUBS 0.006923f
C821 B.n570 VSUBS 0.006923f
C822 B.n571 VSUBS 0.006923f
C823 B.n572 VSUBS 0.006923f
C824 B.n573 VSUBS 0.006923f
C825 B.n574 VSUBS 0.006923f
C826 B.n575 VSUBS 0.006923f
C827 B.n576 VSUBS 0.006923f
C828 B.n577 VSUBS 0.006923f
C829 B.n578 VSUBS 0.006923f
C830 B.n579 VSUBS 0.006923f
C831 B.n580 VSUBS 0.006923f
C832 B.n581 VSUBS 0.006923f
C833 B.n582 VSUBS 0.006923f
C834 B.n583 VSUBS 0.006923f
C835 B.n584 VSUBS 0.006923f
C836 B.n585 VSUBS 0.006923f
C837 B.n586 VSUBS 0.006923f
C838 B.n587 VSUBS 0.006923f
C839 B.n588 VSUBS 0.006923f
C840 B.n589 VSUBS 0.006923f
C841 B.n590 VSUBS 0.006923f
C842 B.n591 VSUBS 0.006923f
C843 B.n592 VSUBS 0.006923f
C844 B.n593 VSUBS 0.006923f
C845 B.n594 VSUBS 0.006923f
C846 B.n595 VSUBS 0.004785f
C847 B.n596 VSUBS 0.01604f
C848 B.n597 VSUBS 0.0056f
C849 B.n598 VSUBS 0.006923f
C850 B.n599 VSUBS 0.006923f
C851 B.n600 VSUBS 0.006923f
C852 B.n601 VSUBS 0.006923f
C853 B.n602 VSUBS 0.006923f
C854 B.n603 VSUBS 0.006923f
C855 B.n604 VSUBS 0.006923f
C856 B.n605 VSUBS 0.006923f
C857 B.n606 VSUBS 0.006923f
C858 B.n607 VSUBS 0.006923f
C859 B.n608 VSUBS 0.006923f
C860 B.n609 VSUBS 0.0056f
C861 B.n610 VSUBS 0.01604f
C862 B.n611 VSUBS 0.004785f
C863 B.n612 VSUBS 0.006923f
C864 B.n613 VSUBS 0.006923f
C865 B.n614 VSUBS 0.006923f
C866 B.n615 VSUBS 0.006923f
C867 B.n616 VSUBS 0.006923f
C868 B.n617 VSUBS 0.006923f
C869 B.n618 VSUBS 0.006923f
C870 B.n619 VSUBS 0.006923f
C871 B.n620 VSUBS 0.006923f
C872 B.n621 VSUBS 0.006923f
C873 B.n622 VSUBS 0.006923f
C874 B.n623 VSUBS 0.006923f
C875 B.n624 VSUBS 0.006923f
C876 B.n625 VSUBS 0.006923f
C877 B.n626 VSUBS 0.006923f
C878 B.n627 VSUBS 0.006923f
C879 B.n628 VSUBS 0.006923f
C880 B.n629 VSUBS 0.006923f
C881 B.n630 VSUBS 0.006923f
C882 B.n631 VSUBS 0.006923f
C883 B.n632 VSUBS 0.006923f
C884 B.n633 VSUBS 0.006923f
C885 B.n634 VSUBS 0.006923f
C886 B.n635 VSUBS 0.006923f
C887 B.n636 VSUBS 0.006923f
C888 B.n637 VSUBS 0.006923f
C889 B.n638 VSUBS 0.006923f
C890 B.n639 VSUBS 0.006923f
C891 B.n640 VSUBS 0.006923f
C892 B.n641 VSUBS 0.006923f
C893 B.n642 VSUBS 0.006923f
C894 B.n643 VSUBS 0.006923f
C895 B.n644 VSUBS 0.006923f
C896 B.n645 VSUBS 0.006923f
C897 B.n646 VSUBS 0.006923f
C898 B.n647 VSUBS 0.006923f
C899 B.n648 VSUBS 0.006923f
C900 B.n649 VSUBS 0.006923f
C901 B.n650 VSUBS 0.006923f
C902 B.n651 VSUBS 0.006923f
C903 B.n652 VSUBS 0.006923f
C904 B.n653 VSUBS 0.006923f
C905 B.n654 VSUBS 0.006923f
C906 B.n655 VSUBS 0.006923f
C907 B.n656 VSUBS 0.006923f
C908 B.n657 VSUBS 0.006923f
C909 B.n658 VSUBS 0.006923f
C910 B.n659 VSUBS 0.006923f
C911 B.n660 VSUBS 0.006923f
C912 B.n661 VSUBS 0.006923f
C913 B.n662 VSUBS 0.006923f
C914 B.n663 VSUBS 0.006923f
C915 B.n664 VSUBS 0.006923f
C916 B.n665 VSUBS 0.006923f
C917 B.n666 VSUBS 0.006923f
C918 B.n667 VSUBS 0.006923f
C919 B.n668 VSUBS 0.006923f
C920 B.n669 VSUBS 0.006923f
C921 B.n670 VSUBS 0.006923f
C922 B.n671 VSUBS 0.006923f
C923 B.n672 VSUBS 0.006923f
C924 B.n673 VSUBS 0.006923f
C925 B.n674 VSUBS 0.006923f
C926 B.n675 VSUBS 0.006923f
C927 B.n676 VSUBS 0.006923f
C928 B.n677 VSUBS 0.006923f
C929 B.n678 VSUBS 0.006923f
C930 B.n679 VSUBS 0.006923f
C931 B.n680 VSUBS 0.006923f
C932 B.n681 VSUBS 0.006923f
C933 B.n682 VSUBS 0.006923f
C934 B.n683 VSUBS 0.006923f
C935 B.n684 VSUBS 0.006923f
C936 B.n685 VSUBS 0.006923f
C937 B.n686 VSUBS 0.006923f
C938 B.n687 VSUBS 0.006923f
C939 B.n688 VSUBS 0.006923f
C940 B.n689 VSUBS 0.006923f
C941 B.n690 VSUBS 0.006923f
C942 B.n691 VSUBS 0.006923f
C943 B.n692 VSUBS 0.006923f
C944 B.n693 VSUBS 0.006923f
C945 B.n694 VSUBS 0.006923f
C946 B.n695 VSUBS 0.006923f
C947 B.n696 VSUBS 0.006923f
C948 B.n697 VSUBS 0.006923f
C949 B.n698 VSUBS 0.006923f
C950 B.n699 VSUBS 0.006923f
C951 B.n700 VSUBS 0.006923f
C952 B.n701 VSUBS 0.006923f
C953 B.n702 VSUBS 0.006923f
C954 B.n703 VSUBS 0.016064f
C955 B.n704 VSUBS 0.014886f
C956 B.n705 VSUBS 0.014886f
C957 B.n706 VSUBS 0.006923f
C958 B.n707 VSUBS 0.006923f
C959 B.n708 VSUBS 0.006923f
C960 B.n709 VSUBS 0.006923f
C961 B.n710 VSUBS 0.006923f
C962 B.n711 VSUBS 0.006923f
C963 B.n712 VSUBS 0.006923f
C964 B.n713 VSUBS 0.006923f
C965 B.n714 VSUBS 0.006923f
C966 B.n715 VSUBS 0.006923f
C967 B.n716 VSUBS 0.006923f
C968 B.n717 VSUBS 0.006923f
C969 B.n718 VSUBS 0.006923f
C970 B.n719 VSUBS 0.006923f
C971 B.n720 VSUBS 0.006923f
C972 B.n721 VSUBS 0.006923f
C973 B.n722 VSUBS 0.006923f
C974 B.n723 VSUBS 0.006923f
C975 B.n724 VSUBS 0.006923f
C976 B.n725 VSUBS 0.006923f
C977 B.n726 VSUBS 0.006923f
C978 B.n727 VSUBS 0.006923f
C979 B.n728 VSUBS 0.006923f
C980 B.n729 VSUBS 0.006923f
C981 B.n730 VSUBS 0.006923f
C982 B.n731 VSUBS 0.006923f
C983 B.n732 VSUBS 0.006923f
C984 B.n733 VSUBS 0.006923f
C985 B.n734 VSUBS 0.006923f
C986 B.n735 VSUBS 0.006923f
C987 B.n736 VSUBS 0.006923f
C988 B.n737 VSUBS 0.006923f
C989 B.n738 VSUBS 0.006923f
C990 B.n739 VSUBS 0.009034f
C991 B.n740 VSUBS 0.009624f
C992 B.n741 VSUBS 0.019138f
C993 VDD2.n0 VSUBS 0.015781f
C994 VDD2.n1 VSUBS 0.035608f
C995 VDD2.n2 VSUBS 0.015951f
C996 VDD2.n3 VSUBS 0.028036f
C997 VDD2.n4 VSUBS 0.015065f
C998 VDD2.n5 VSUBS 0.035608f
C999 VDD2.n6 VSUBS 0.015951f
C1000 VDD2.n7 VSUBS 0.028036f
C1001 VDD2.n8 VSUBS 0.015065f
C1002 VDD2.n9 VSUBS 0.035608f
C1003 VDD2.n10 VSUBS 0.015951f
C1004 VDD2.n11 VSUBS 0.028036f
C1005 VDD2.n12 VSUBS 0.015065f
C1006 VDD2.n13 VSUBS 0.035608f
C1007 VDD2.n14 VSUBS 0.015951f
C1008 VDD2.n15 VSUBS 0.028036f
C1009 VDD2.n16 VSUBS 0.015065f
C1010 VDD2.n17 VSUBS 0.035608f
C1011 VDD2.n18 VSUBS 0.015951f
C1012 VDD2.n19 VSUBS 0.028036f
C1013 VDD2.n20 VSUBS 0.015065f
C1014 VDD2.n21 VSUBS 0.035608f
C1015 VDD2.n22 VSUBS 0.015508f
C1016 VDD2.n23 VSUBS 0.028036f
C1017 VDD2.n24 VSUBS 0.015951f
C1018 VDD2.n25 VSUBS 0.035608f
C1019 VDD2.n26 VSUBS 0.015951f
C1020 VDD2.n27 VSUBS 0.028036f
C1021 VDD2.n28 VSUBS 0.015065f
C1022 VDD2.n29 VSUBS 0.035608f
C1023 VDD2.n30 VSUBS 0.015951f
C1024 VDD2.n31 VSUBS 2.20789f
C1025 VDD2.n32 VSUBS 0.015065f
C1026 VDD2.t1 VSUBS 0.077372f
C1027 VDD2.n33 VSUBS 0.306489f
C1028 VDD2.n34 VSUBS 0.026787f
C1029 VDD2.n35 VSUBS 0.026706f
C1030 VDD2.n36 VSUBS 0.035608f
C1031 VDD2.n37 VSUBS 0.015951f
C1032 VDD2.n38 VSUBS 0.015065f
C1033 VDD2.n39 VSUBS 0.028036f
C1034 VDD2.n40 VSUBS 0.028036f
C1035 VDD2.n41 VSUBS 0.015065f
C1036 VDD2.n42 VSUBS 0.015951f
C1037 VDD2.n43 VSUBS 0.035608f
C1038 VDD2.n44 VSUBS 0.035608f
C1039 VDD2.n45 VSUBS 0.015951f
C1040 VDD2.n46 VSUBS 0.015065f
C1041 VDD2.n47 VSUBS 0.028036f
C1042 VDD2.n48 VSUBS 0.028036f
C1043 VDD2.n49 VSUBS 0.015065f
C1044 VDD2.n50 VSUBS 0.015065f
C1045 VDD2.n51 VSUBS 0.015951f
C1046 VDD2.n52 VSUBS 0.035608f
C1047 VDD2.n53 VSUBS 0.035608f
C1048 VDD2.n54 VSUBS 0.035608f
C1049 VDD2.n55 VSUBS 0.015508f
C1050 VDD2.n56 VSUBS 0.015065f
C1051 VDD2.n57 VSUBS 0.028036f
C1052 VDD2.n58 VSUBS 0.028036f
C1053 VDD2.n59 VSUBS 0.015065f
C1054 VDD2.n60 VSUBS 0.015951f
C1055 VDD2.n61 VSUBS 0.035608f
C1056 VDD2.n62 VSUBS 0.035608f
C1057 VDD2.n63 VSUBS 0.015951f
C1058 VDD2.n64 VSUBS 0.015065f
C1059 VDD2.n65 VSUBS 0.028036f
C1060 VDD2.n66 VSUBS 0.028036f
C1061 VDD2.n67 VSUBS 0.015065f
C1062 VDD2.n68 VSUBS 0.015951f
C1063 VDD2.n69 VSUBS 0.035608f
C1064 VDD2.n70 VSUBS 0.035608f
C1065 VDD2.n71 VSUBS 0.015951f
C1066 VDD2.n72 VSUBS 0.015065f
C1067 VDD2.n73 VSUBS 0.028036f
C1068 VDD2.n74 VSUBS 0.028036f
C1069 VDD2.n75 VSUBS 0.015065f
C1070 VDD2.n76 VSUBS 0.015951f
C1071 VDD2.n77 VSUBS 0.035608f
C1072 VDD2.n78 VSUBS 0.035608f
C1073 VDD2.n79 VSUBS 0.015951f
C1074 VDD2.n80 VSUBS 0.015065f
C1075 VDD2.n81 VSUBS 0.028036f
C1076 VDD2.n82 VSUBS 0.028036f
C1077 VDD2.n83 VSUBS 0.015065f
C1078 VDD2.n84 VSUBS 0.015951f
C1079 VDD2.n85 VSUBS 0.035608f
C1080 VDD2.n86 VSUBS 0.035608f
C1081 VDD2.n87 VSUBS 0.015951f
C1082 VDD2.n88 VSUBS 0.015065f
C1083 VDD2.n89 VSUBS 0.028036f
C1084 VDD2.n90 VSUBS 0.028036f
C1085 VDD2.n91 VSUBS 0.015065f
C1086 VDD2.n92 VSUBS 0.015951f
C1087 VDD2.n93 VSUBS 0.035608f
C1088 VDD2.n94 VSUBS 0.035608f
C1089 VDD2.n95 VSUBS 0.015951f
C1090 VDD2.n96 VSUBS 0.015065f
C1091 VDD2.n97 VSUBS 0.028036f
C1092 VDD2.n98 VSUBS 0.070931f
C1093 VDD2.n99 VSUBS 0.015065f
C1094 VDD2.n100 VSUBS 0.015951f
C1095 VDD2.n101 VSUBS 0.079328f
C1096 VDD2.n102 VSUBS 1.07917f
C1097 VDD2.n103 VSUBS 0.015781f
C1098 VDD2.n104 VSUBS 0.035608f
C1099 VDD2.n105 VSUBS 0.015951f
C1100 VDD2.n106 VSUBS 0.028036f
C1101 VDD2.n107 VSUBS 0.015065f
C1102 VDD2.n108 VSUBS 0.035608f
C1103 VDD2.n109 VSUBS 0.015951f
C1104 VDD2.n110 VSUBS 0.028036f
C1105 VDD2.n111 VSUBS 0.015065f
C1106 VDD2.n112 VSUBS 0.035608f
C1107 VDD2.n113 VSUBS 0.015951f
C1108 VDD2.n114 VSUBS 0.028036f
C1109 VDD2.n115 VSUBS 0.015065f
C1110 VDD2.n116 VSUBS 0.035608f
C1111 VDD2.n117 VSUBS 0.015951f
C1112 VDD2.n118 VSUBS 0.028036f
C1113 VDD2.n119 VSUBS 0.015065f
C1114 VDD2.n120 VSUBS 0.035608f
C1115 VDD2.n121 VSUBS 0.015951f
C1116 VDD2.n122 VSUBS 0.028036f
C1117 VDD2.n123 VSUBS 0.015065f
C1118 VDD2.n124 VSUBS 0.035608f
C1119 VDD2.n125 VSUBS 0.015508f
C1120 VDD2.n126 VSUBS 0.028036f
C1121 VDD2.n127 VSUBS 0.015508f
C1122 VDD2.n128 VSUBS 0.015065f
C1123 VDD2.n129 VSUBS 0.035608f
C1124 VDD2.n130 VSUBS 0.035608f
C1125 VDD2.n131 VSUBS 0.015951f
C1126 VDD2.n132 VSUBS 0.028036f
C1127 VDD2.n133 VSUBS 0.015065f
C1128 VDD2.n134 VSUBS 0.035608f
C1129 VDD2.n135 VSUBS 0.015951f
C1130 VDD2.n136 VSUBS 2.20789f
C1131 VDD2.n137 VSUBS 0.015065f
C1132 VDD2.t0 VSUBS 0.077372f
C1133 VDD2.n138 VSUBS 0.306489f
C1134 VDD2.n139 VSUBS 0.026787f
C1135 VDD2.n140 VSUBS 0.026706f
C1136 VDD2.n141 VSUBS 0.035608f
C1137 VDD2.n142 VSUBS 0.015951f
C1138 VDD2.n143 VSUBS 0.015065f
C1139 VDD2.n144 VSUBS 0.028036f
C1140 VDD2.n145 VSUBS 0.028036f
C1141 VDD2.n146 VSUBS 0.015065f
C1142 VDD2.n147 VSUBS 0.015951f
C1143 VDD2.n148 VSUBS 0.035608f
C1144 VDD2.n149 VSUBS 0.035608f
C1145 VDD2.n150 VSUBS 0.015951f
C1146 VDD2.n151 VSUBS 0.015065f
C1147 VDD2.n152 VSUBS 0.028036f
C1148 VDD2.n153 VSUBS 0.028036f
C1149 VDD2.n154 VSUBS 0.015065f
C1150 VDD2.n155 VSUBS 0.015951f
C1151 VDD2.n156 VSUBS 0.035608f
C1152 VDD2.n157 VSUBS 0.035608f
C1153 VDD2.n158 VSUBS 0.015951f
C1154 VDD2.n159 VSUBS 0.015065f
C1155 VDD2.n160 VSUBS 0.028036f
C1156 VDD2.n161 VSUBS 0.028036f
C1157 VDD2.n162 VSUBS 0.015065f
C1158 VDD2.n163 VSUBS 0.015951f
C1159 VDD2.n164 VSUBS 0.035608f
C1160 VDD2.n165 VSUBS 0.035608f
C1161 VDD2.n166 VSUBS 0.015951f
C1162 VDD2.n167 VSUBS 0.015065f
C1163 VDD2.n168 VSUBS 0.028036f
C1164 VDD2.n169 VSUBS 0.028036f
C1165 VDD2.n170 VSUBS 0.015065f
C1166 VDD2.n171 VSUBS 0.015951f
C1167 VDD2.n172 VSUBS 0.035608f
C1168 VDD2.n173 VSUBS 0.035608f
C1169 VDD2.n174 VSUBS 0.015951f
C1170 VDD2.n175 VSUBS 0.015065f
C1171 VDD2.n176 VSUBS 0.028036f
C1172 VDD2.n177 VSUBS 0.028036f
C1173 VDD2.n178 VSUBS 0.015065f
C1174 VDD2.n179 VSUBS 0.015951f
C1175 VDD2.n180 VSUBS 0.035608f
C1176 VDD2.n181 VSUBS 0.035608f
C1177 VDD2.n182 VSUBS 0.015951f
C1178 VDD2.n183 VSUBS 0.015065f
C1179 VDD2.n184 VSUBS 0.028036f
C1180 VDD2.n185 VSUBS 0.028036f
C1181 VDD2.n186 VSUBS 0.015065f
C1182 VDD2.n187 VSUBS 0.015951f
C1183 VDD2.n188 VSUBS 0.035608f
C1184 VDD2.n189 VSUBS 0.035608f
C1185 VDD2.n190 VSUBS 0.015951f
C1186 VDD2.n191 VSUBS 0.015065f
C1187 VDD2.n192 VSUBS 0.028036f
C1188 VDD2.n193 VSUBS 0.028036f
C1189 VDD2.n194 VSUBS 0.015065f
C1190 VDD2.n195 VSUBS 0.015951f
C1191 VDD2.n196 VSUBS 0.035608f
C1192 VDD2.n197 VSUBS 0.035608f
C1193 VDD2.n198 VSUBS 0.015951f
C1194 VDD2.n199 VSUBS 0.015065f
C1195 VDD2.n200 VSUBS 0.028036f
C1196 VDD2.n201 VSUBS 0.070931f
C1197 VDD2.n202 VSUBS 0.015065f
C1198 VDD2.n203 VSUBS 0.015951f
C1199 VDD2.n204 VSUBS 0.079328f
C1200 VDD2.n205 VSUBS 0.071642f
C1201 VDD2.n206 VSUBS 4.19595f
C1202 VTAIL.n0 VSUBS 0.015696f
C1203 VTAIL.n1 VSUBS 0.035416f
C1204 VTAIL.n2 VSUBS 0.015865f
C1205 VTAIL.n3 VSUBS 0.027884f
C1206 VTAIL.n4 VSUBS 0.014984f
C1207 VTAIL.n5 VSUBS 0.035416f
C1208 VTAIL.n6 VSUBS 0.015865f
C1209 VTAIL.n7 VSUBS 0.027884f
C1210 VTAIL.n8 VSUBS 0.014984f
C1211 VTAIL.n9 VSUBS 0.035416f
C1212 VTAIL.n10 VSUBS 0.015865f
C1213 VTAIL.n11 VSUBS 0.027884f
C1214 VTAIL.n12 VSUBS 0.014984f
C1215 VTAIL.n13 VSUBS 0.035416f
C1216 VTAIL.n14 VSUBS 0.015865f
C1217 VTAIL.n15 VSUBS 0.027884f
C1218 VTAIL.n16 VSUBS 0.014984f
C1219 VTAIL.n17 VSUBS 0.035416f
C1220 VTAIL.n18 VSUBS 0.015865f
C1221 VTAIL.n19 VSUBS 0.027884f
C1222 VTAIL.n20 VSUBS 0.014984f
C1223 VTAIL.n21 VSUBS 0.035416f
C1224 VTAIL.n22 VSUBS 0.015424f
C1225 VTAIL.n23 VSUBS 0.027884f
C1226 VTAIL.n24 VSUBS 0.015865f
C1227 VTAIL.n25 VSUBS 0.035416f
C1228 VTAIL.n26 VSUBS 0.015865f
C1229 VTAIL.n27 VSUBS 0.027884f
C1230 VTAIL.n28 VSUBS 0.014984f
C1231 VTAIL.n29 VSUBS 0.035416f
C1232 VTAIL.n30 VSUBS 0.015865f
C1233 VTAIL.n31 VSUBS 2.19595f
C1234 VTAIL.n32 VSUBS 0.014984f
C1235 VTAIL.t0 VSUBS 0.076954f
C1236 VTAIL.n33 VSUBS 0.304833f
C1237 VTAIL.n34 VSUBS 0.026642f
C1238 VTAIL.n35 VSUBS 0.026562f
C1239 VTAIL.n36 VSUBS 0.035416f
C1240 VTAIL.n37 VSUBS 0.015865f
C1241 VTAIL.n38 VSUBS 0.014984f
C1242 VTAIL.n39 VSUBS 0.027884f
C1243 VTAIL.n40 VSUBS 0.027884f
C1244 VTAIL.n41 VSUBS 0.014984f
C1245 VTAIL.n42 VSUBS 0.015865f
C1246 VTAIL.n43 VSUBS 0.035416f
C1247 VTAIL.n44 VSUBS 0.035416f
C1248 VTAIL.n45 VSUBS 0.015865f
C1249 VTAIL.n46 VSUBS 0.014984f
C1250 VTAIL.n47 VSUBS 0.027884f
C1251 VTAIL.n48 VSUBS 0.027884f
C1252 VTAIL.n49 VSUBS 0.014984f
C1253 VTAIL.n50 VSUBS 0.014984f
C1254 VTAIL.n51 VSUBS 0.015865f
C1255 VTAIL.n52 VSUBS 0.035416f
C1256 VTAIL.n53 VSUBS 0.035416f
C1257 VTAIL.n54 VSUBS 0.035416f
C1258 VTAIL.n55 VSUBS 0.015424f
C1259 VTAIL.n56 VSUBS 0.014984f
C1260 VTAIL.n57 VSUBS 0.027884f
C1261 VTAIL.n58 VSUBS 0.027884f
C1262 VTAIL.n59 VSUBS 0.014984f
C1263 VTAIL.n60 VSUBS 0.015865f
C1264 VTAIL.n61 VSUBS 0.035416f
C1265 VTAIL.n62 VSUBS 0.035416f
C1266 VTAIL.n63 VSUBS 0.015865f
C1267 VTAIL.n64 VSUBS 0.014984f
C1268 VTAIL.n65 VSUBS 0.027884f
C1269 VTAIL.n66 VSUBS 0.027884f
C1270 VTAIL.n67 VSUBS 0.014984f
C1271 VTAIL.n68 VSUBS 0.015865f
C1272 VTAIL.n69 VSUBS 0.035416f
C1273 VTAIL.n70 VSUBS 0.035416f
C1274 VTAIL.n71 VSUBS 0.015865f
C1275 VTAIL.n72 VSUBS 0.014984f
C1276 VTAIL.n73 VSUBS 0.027884f
C1277 VTAIL.n74 VSUBS 0.027884f
C1278 VTAIL.n75 VSUBS 0.014984f
C1279 VTAIL.n76 VSUBS 0.015865f
C1280 VTAIL.n77 VSUBS 0.035416f
C1281 VTAIL.n78 VSUBS 0.035416f
C1282 VTAIL.n79 VSUBS 0.015865f
C1283 VTAIL.n80 VSUBS 0.014984f
C1284 VTAIL.n81 VSUBS 0.027884f
C1285 VTAIL.n82 VSUBS 0.027884f
C1286 VTAIL.n83 VSUBS 0.014984f
C1287 VTAIL.n84 VSUBS 0.015865f
C1288 VTAIL.n85 VSUBS 0.035416f
C1289 VTAIL.n86 VSUBS 0.035416f
C1290 VTAIL.n87 VSUBS 0.015865f
C1291 VTAIL.n88 VSUBS 0.014984f
C1292 VTAIL.n89 VSUBS 0.027884f
C1293 VTAIL.n90 VSUBS 0.027884f
C1294 VTAIL.n91 VSUBS 0.014984f
C1295 VTAIL.n92 VSUBS 0.015865f
C1296 VTAIL.n93 VSUBS 0.035416f
C1297 VTAIL.n94 VSUBS 0.035416f
C1298 VTAIL.n95 VSUBS 0.015865f
C1299 VTAIL.n96 VSUBS 0.014984f
C1300 VTAIL.n97 VSUBS 0.027884f
C1301 VTAIL.n98 VSUBS 0.070547f
C1302 VTAIL.n99 VSUBS 0.014984f
C1303 VTAIL.n100 VSUBS 0.015865f
C1304 VTAIL.n101 VSUBS 0.078899f
C1305 VTAIL.n102 VSUBS 0.05204f
C1306 VTAIL.n103 VSUBS 2.39234f
C1307 VTAIL.n104 VSUBS 0.015696f
C1308 VTAIL.n105 VSUBS 0.035416f
C1309 VTAIL.n106 VSUBS 0.015865f
C1310 VTAIL.n107 VSUBS 0.027884f
C1311 VTAIL.n108 VSUBS 0.014984f
C1312 VTAIL.n109 VSUBS 0.035416f
C1313 VTAIL.n110 VSUBS 0.015865f
C1314 VTAIL.n111 VSUBS 0.027884f
C1315 VTAIL.n112 VSUBS 0.014984f
C1316 VTAIL.n113 VSUBS 0.035416f
C1317 VTAIL.n114 VSUBS 0.015865f
C1318 VTAIL.n115 VSUBS 0.027884f
C1319 VTAIL.n116 VSUBS 0.014984f
C1320 VTAIL.n117 VSUBS 0.035416f
C1321 VTAIL.n118 VSUBS 0.015865f
C1322 VTAIL.n119 VSUBS 0.027884f
C1323 VTAIL.n120 VSUBS 0.014984f
C1324 VTAIL.n121 VSUBS 0.035416f
C1325 VTAIL.n122 VSUBS 0.015865f
C1326 VTAIL.n123 VSUBS 0.027884f
C1327 VTAIL.n124 VSUBS 0.014984f
C1328 VTAIL.n125 VSUBS 0.035416f
C1329 VTAIL.n126 VSUBS 0.015424f
C1330 VTAIL.n127 VSUBS 0.027884f
C1331 VTAIL.n128 VSUBS 0.015424f
C1332 VTAIL.n129 VSUBS 0.014984f
C1333 VTAIL.n130 VSUBS 0.035416f
C1334 VTAIL.n131 VSUBS 0.035416f
C1335 VTAIL.n132 VSUBS 0.015865f
C1336 VTAIL.n133 VSUBS 0.027884f
C1337 VTAIL.n134 VSUBS 0.014984f
C1338 VTAIL.n135 VSUBS 0.035416f
C1339 VTAIL.n136 VSUBS 0.015865f
C1340 VTAIL.n137 VSUBS 2.19595f
C1341 VTAIL.n138 VSUBS 0.014984f
C1342 VTAIL.t2 VSUBS 0.076954f
C1343 VTAIL.n139 VSUBS 0.304833f
C1344 VTAIL.n140 VSUBS 0.026642f
C1345 VTAIL.n141 VSUBS 0.026562f
C1346 VTAIL.n142 VSUBS 0.035416f
C1347 VTAIL.n143 VSUBS 0.015865f
C1348 VTAIL.n144 VSUBS 0.014984f
C1349 VTAIL.n145 VSUBS 0.027884f
C1350 VTAIL.n146 VSUBS 0.027884f
C1351 VTAIL.n147 VSUBS 0.014984f
C1352 VTAIL.n148 VSUBS 0.015865f
C1353 VTAIL.n149 VSUBS 0.035416f
C1354 VTAIL.n150 VSUBS 0.035416f
C1355 VTAIL.n151 VSUBS 0.015865f
C1356 VTAIL.n152 VSUBS 0.014984f
C1357 VTAIL.n153 VSUBS 0.027884f
C1358 VTAIL.n154 VSUBS 0.027884f
C1359 VTAIL.n155 VSUBS 0.014984f
C1360 VTAIL.n156 VSUBS 0.015865f
C1361 VTAIL.n157 VSUBS 0.035416f
C1362 VTAIL.n158 VSUBS 0.035416f
C1363 VTAIL.n159 VSUBS 0.015865f
C1364 VTAIL.n160 VSUBS 0.014984f
C1365 VTAIL.n161 VSUBS 0.027884f
C1366 VTAIL.n162 VSUBS 0.027884f
C1367 VTAIL.n163 VSUBS 0.014984f
C1368 VTAIL.n164 VSUBS 0.015865f
C1369 VTAIL.n165 VSUBS 0.035416f
C1370 VTAIL.n166 VSUBS 0.035416f
C1371 VTAIL.n167 VSUBS 0.015865f
C1372 VTAIL.n168 VSUBS 0.014984f
C1373 VTAIL.n169 VSUBS 0.027884f
C1374 VTAIL.n170 VSUBS 0.027884f
C1375 VTAIL.n171 VSUBS 0.014984f
C1376 VTAIL.n172 VSUBS 0.015865f
C1377 VTAIL.n173 VSUBS 0.035416f
C1378 VTAIL.n174 VSUBS 0.035416f
C1379 VTAIL.n175 VSUBS 0.015865f
C1380 VTAIL.n176 VSUBS 0.014984f
C1381 VTAIL.n177 VSUBS 0.027884f
C1382 VTAIL.n178 VSUBS 0.027884f
C1383 VTAIL.n179 VSUBS 0.014984f
C1384 VTAIL.n180 VSUBS 0.015865f
C1385 VTAIL.n181 VSUBS 0.035416f
C1386 VTAIL.n182 VSUBS 0.035416f
C1387 VTAIL.n183 VSUBS 0.015865f
C1388 VTAIL.n184 VSUBS 0.014984f
C1389 VTAIL.n185 VSUBS 0.027884f
C1390 VTAIL.n186 VSUBS 0.027884f
C1391 VTAIL.n187 VSUBS 0.014984f
C1392 VTAIL.n188 VSUBS 0.015865f
C1393 VTAIL.n189 VSUBS 0.035416f
C1394 VTAIL.n190 VSUBS 0.035416f
C1395 VTAIL.n191 VSUBS 0.015865f
C1396 VTAIL.n192 VSUBS 0.014984f
C1397 VTAIL.n193 VSUBS 0.027884f
C1398 VTAIL.n194 VSUBS 0.027884f
C1399 VTAIL.n195 VSUBS 0.014984f
C1400 VTAIL.n196 VSUBS 0.015865f
C1401 VTAIL.n197 VSUBS 0.035416f
C1402 VTAIL.n198 VSUBS 0.035416f
C1403 VTAIL.n199 VSUBS 0.015865f
C1404 VTAIL.n200 VSUBS 0.014984f
C1405 VTAIL.n201 VSUBS 0.027884f
C1406 VTAIL.n202 VSUBS 0.070547f
C1407 VTAIL.n203 VSUBS 0.014984f
C1408 VTAIL.n204 VSUBS 0.015865f
C1409 VTAIL.n205 VSUBS 0.078899f
C1410 VTAIL.n206 VSUBS 0.05204f
C1411 VTAIL.n207 VSUBS 2.44114f
C1412 VTAIL.n208 VSUBS 0.015696f
C1413 VTAIL.n209 VSUBS 0.035416f
C1414 VTAIL.n210 VSUBS 0.015865f
C1415 VTAIL.n211 VSUBS 0.027884f
C1416 VTAIL.n212 VSUBS 0.014984f
C1417 VTAIL.n213 VSUBS 0.035416f
C1418 VTAIL.n214 VSUBS 0.015865f
C1419 VTAIL.n215 VSUBS 0.027884f
C1420 VTAIL.n216 VSUBS 0.014984f
C1421 VTAIL.n217 VSUBS 0.035416f
C1422 VTAIL.n218 VSUBS 0.015865f
C1423 VTAIL.n219 VSUBS 0.027884f
C1424 VTAIL.n220 VSUBS 0.014984f
C1425 VTAIL.n221 VSUBS 0.035416f
C1426 VTAIL.n222 VSUBS 0.015865f
C1427 VTAIL.n223 VSUBS 0.027884f
C1428 VTAIL.n224 VSUBS 0.014984f
C1429 VTAIL.n225 VSUBS 0.035416f
C1430 VTAIL.n226 VSUBS 0.015865f
C1431 VTAIL.n227 VSUBS 0.027884f
C1432 VTAIL.n228 VSUBS 0.014984f
C1433 VTAIL.n229 VSUBS 0.035416f
C1434 VTAIL.n230 VSUBS 0.015424f
C1435 VTAIL.n231 VSUBS 0.027884f
C1436 VTAIL.n232 VSUBS 0.015424f
C1437 VTAIL.n233 VSUBS 0.014984f
C1438 VTAIL.n234 VSUBS 0.035416f
C1439 VTAIL.n235 VSUBS 0.035416f
C1440 VTAIL.n236 VSUBS 0.015865f
C1441 VTAIL.n237 VSUBS 0.027884f
C1442 VTAIL.n238 VSUBS 0.014984f
C1443 VTAIL.n239 VSUBS 0.035416f
C1444 VTAIL.n240 VSUBS 0.015865f
C1445 VTAIL.n241 VSUBS 2.19595f
C1446 VTAIL.n242 VSUBS 0.014984f
C1447 VTAIL.t1 VSUBS 0.076954f
C1448 VTAIL.n243 VSUBS 0.304832f
C1449 VTAIL.n244 VSUBS 0.026642f
C1450 VTAIL.n245 VSUBS 0.026562f
C1451 VTAIL.n246 VSUBS 0.035416f
C1452 VTAIL.n247 VSUBS 0.015865f
C1453 VTAIL.n248 VSUBS 0.014984f
C1454 VTAIL.n249 VSUBS 0.027884f
C1455 VTAIL.n250 VSUBS 0.027884f
C1456 VTAIL.n251 VSUBS 0.014984f
C1457 VTAIL.n252 VSUBS 0.015865f
C1458 VTAIL.n253 VSUBS 0.035416f
C1459 VTAIL.n254 VSUBS 0.035416f
C1460 VTAIL.n255 VSUBS 0.015865f
C1461 VTAIL.n256 VSUBS 0.014984f
C1462 VTAIL.n257 VSUBS 0.027884f
C1463 VTAIL.n258 VSUBS 0.027884f
C1464 VTAIL.n259 VSUBS 0.014984f
C1465 VTAIL.n260 VSUBS 0.015865f
C1466 VTAIL.n261 VSUBS 0.035416f
C1467 VTAIL.n262 VSUBS 0.035416f
C1468 VTAIL.n263 VSUBS 0.015865f
C1469 VTAIL.n264 VSUBS 0.014984f
C1470 VTAIL.n265 VSUBS 0.027884f
C1471 VTAIL.n266 VSUBS 0.027884f
C1472 VTAIL.n267 VSUBS 0.014984f
C1473 VTAIL.n268 VSUBS 0.015865f
C1474 VTAIL.n269 VSUBS 0.035416f
C1475 VTAIL.n270 VSUBS 0.035416f
C1476 VTAIL.n271 VSUBS 0.015865f
C1477 VTAIL.n272 VSUBS 0.014984f
C1478 VTAIL.n273 VSUBS 0.027884f
C1479 VTAIL.n274 VSUBS 0.027884f
C1480 VTAIL.n275 VSUBS 0.014984f
C1481 VTAIL.n276 VSUBS 0.015865f
C1482 VTAIL.n277 VSUBS 0.035416f
C1483 VTAIL.n278 VSUBS 0.035416f
C1484 VTAIL.n279 VSUBS 0.015865f
C1485 VTAIL.n280 VSUBS 0.014984f
C1486 VTAIL.n281 VSUBS 0.027884f
C1487 VTAIL.n282 VSUBS 0.027884f
C1488 VTAIL.n283 VSUBS 0.014984f
C1489 VTAIL.n284 VSUBS 0.015865f
C1490 VTAIL.n285 VSUBS 0.035416f
C1491 VTAIL.n286 VSUBS 0.035416f
C1492 VTAIL.n287 VSUBS 0.015865f
C1493 VTAIL.n288 VSUBS 0.014984f
C1494 VTAIL.n289 VSUBS 0.027884f
C1495 VTAIL.n290 VSUBS 0.027884f
C1496 VTAIL.n291 VSUBS 0.014984f
C1497 VTAIL.n292 VSUBS 0.015865f
C1498 VTAIL.n293 VSUBS 0.035416f
C1499 VTAIL.n294 VSUBS 0.035416f
C1500 VTAIL.n295 VSUBS 0.015865f
C1501 VTAIL.n296 VSUBS 0.014984f
C1502 VTAIL.n297 VSUBS 0.027884f
C1503 VTAIL.n298 VSUBS 0.027884f
C1504 VTAIL.n299 VSUBS 0.014984f
C1505 VTAIL.n300 VSUBS 0.015865f
C1506 VTAIL.n301 VSUBS 0.035416f
C1507 VTAIL.n302 VSUBS 0.035416f
C1508 VTAIL.n303 VSUBS 0.015865f
C1509 VTAIL.n304 VSUBS 0.014984f
C1510 VTAIL.n305 VSUBS 0.027884f
C1511 VTAIL.n306 VSUBS 0.070547f
C1512 VTAIL.n307 VSUBS 0.014984f
C1513 VTAIL.n308 VSUBS 0.015865f
C1514 VTAIL.n309 VSUBS 0.078899f
C1515 VTAIL.n310 VSUBS 0.05204f
C1516 VTAIL.n311 VSUBS 2.22504f
C1517 VTAIL.n312 VSUBS 0.015696f
C1518 VTAIL.n313 VSUBS 0.035416f
C1519 VTAIL.n314 VSUBS 0.015865f
C1520 VTAIL.n315 VSUBS 0.027884f
C1521 VTAIL.n316 VSUBS 0.014984f
C1522 VTAIL.n317 VSUBS 0.035416f
C1523 VTAIL.n318 VSUBS 0.015865f
C1524 VTAIL.n319 VSUBS 0.027884f
C1525 VTAIL.n320 VSUBS 0.014984f
C1526 VTAIL.n321 VSUBS 0.035416f
C1527 VTAIL.n322 VSUBS 0.015865f
C1528 VTAIL.n323 VSUBS 0.027884f
C1529 VTAIL.n324 VSUBS 0.014984f
C1530 VTAIL.n325 VSUBS 0.035416f
C1531 VTAIL.n326 VSUBS 0.015865f
C1532 VTAIL.n327 VSUBS 0.027884f
C1533 VTAIL.n328 VSUBS 0.014984f
C1534 VTAIL.n329 VSUBS 0.035416f
C1535 VTAIL.n330 VSUBS 0.015865f
C1536 VTAIL.n331 VSUBS 0.027884f
C1537 VTAIL.n332 VSUBS 0.014984f
C1538 VTAIL.n333 VSUBS 0.035416f
C1539 VTAIL.n334 VSUBS 0.015424f
C1540 VTAIL.n335 VSUBS 0.027884f
C1541 VTAIL.n336 VSUBS 0.015865f
C1542 VTAIL.n337 VSUBS 0.035416f
C1543 VTAIL.n338 VSUBS 0.015865f
C1544 VTAIL.n339 VSUBS 0.027884f
C1545 VTAIL.n340 VSUBS 0.014984f
C1546 VTAIL.n341 VSUBS 0.035416f
C1547 VTAIL.n342 VSUBS 0.015865f
C1548 VTAIL.n343 VSUBS 2.19595f
C1549 VTAIL.n344 VSUBS 0.014984f
C1550 VTAIL.t3 VSUBS 0.076954f
C1551 VTAIL.n345 VSUBS 0.304833f
C1552 VTAIL.n346 VSUBS 0.026642f
C1553 VTAIL.n347 VSUBS 0.026562f
C1554 VTAIL.n348 VSUBS 0.035416f
C1555 VTAIL.n349 VSUBS 0.015865f
C1556 VTAIL.n350 VSUBS 0.014984f
C1557 VTAIL.n351 VSUBS 0.027884f
C1558 VTAIL.n352 VSUBS 0.027884f
C1559 VTAIL.n353 VSUBS 0.014984f
C1560 VTAIL.n354 VSUBS 0.015865f
C1561 VTAIL.n355 VSUBS 0.035416f
C1562 VTAIL.n356 VSUBS 0.035416f
C1563 VTAIL.n357 VSUBS 0.015865f
C1564 VTAIL.n358 VSUBS 0.014984f
C1565 VTAIL.n359 VSUBS 0.027884f
C1566 VTAIL.n360 VSUBS 0.027884f
C1567 VTAIL.n361 VSUBS 0.014984f
C1568 VTAIL.n362 VSUBS 0.014984f
C1569 VTAIL.n363 VSUBS 0.015865f
C1570 VTAIL.n364 VSUBS 0.035416f
C1571 VTAIL.n365 VSUBS 0.035416f
C1572 VTAIL.n366 VSUBS 0.035416f
C1573 VTAIL.n367 VSUBS 0.015424f
C1574 VTAIL.n368 VSUBS 0.014984f
C1575 VTAIL.n369 VSUBS 0.027884f
C1576 VTAIL.n370 VSUBS 0.027884f
C1577 VTAIL.n371 VSUBS 0.014984f
C1578 VTAIL.n372 VSUBS 0.015865f
C1579 VTAIL.n373 VSUBS 0.035416f
C1580 VTAIL.n374 VSUBS 0.035416f
C1581 VTAIL.n375 VSUBS 0.015865f
C1582 VTAIL.n376 VSUBS 0.014984f
C1583 VTAIL.n377 VSUBS 0.027884f
C1584 VTAIL.n378 VSUBS 0.027884f
C1585 VTAIL.n379 VSUBS 0.014984f
C1586 VTAIL.n380 VSUBS 0.015865f
C1587 VTAIL.n381 VSUBS 0.035416f
C1588 VTAIL.n382 VSUBS 0.035416f
C1589 VTAIL.n383 VSUBS 0.015865f
C1590 VTAIL.n384 VSUBS 0.014984f
C1591 VTAIL.n385 VSUBS 0.027884f
C1592 VTAIL.n386 VSUBS 0.027884f
C1593 VTAIL.n387 VSUBS 0.014984f
C1594 VTAIL.n388 VSUBS 0.015865f
C1595 VTAIL.n389 VSUBS 0.035416f
C1596 VTAIL.n390 VSUBS 0.035416f
C1597 VTAIL.n391 VSUBS 0.015865f
C1598 VTAIL.n392 VSUBS 0.014984f
C1599 VTAIL.n393 VSUBS 0.027884f
C1600 VTAIL.n394 VSUBS 0.027884f
C1601 VTAIL.n395 VSUBS 0.014984f
C1602 VTAIL.n396 VSUBS 0.015865f
C1603 VTAIL.n397 VSUBS 0.035416f
C1604 VTAIL.n398 VSUBS 0.035416f
C1605 VTAIL.n399 VSUBS 0.015865f
C1606 VTAIL.n400 VSUBS 0.014984f
C1607 VTAIL.n401 VSUBS 0.027884f
C1608 VTAIL.n402 VSUBS 0.027884f
C1609 VTAIL.n403 VSUBS 0.014984f
C1610 VTAIL.n404 VSUBS 0.015865f
C1611 VTAIL.n405 VSUBS 0.035416f
C1612 VTAIL.n406 VSUBS 0.035416f
C1613 VTAIL.n407 VSUBS 0.015865f
C1614 VTAIL.n408 VSUBS 0.014984f
C1615 VTAIL.n409 VSUBS 0.027884f
C1616 VTAIL.n410 VSUBS 0.070547f
C1617 VTAIL.n411 VSUBS 0.014984f
C1618 VTAIL.n412 VSUBS 0.015865f
C1619 VTAIL.n413 VSUBS 0.078899f
C1620 VTAIL.n414 VSUBS 0.05204f
C1621 VTAIL.n415 VSUBS 2.12357f
C1622 VN.t0 VSUBS 5.04665f
C1623 VN.t1 VSUBS 5.67164f
.ends

