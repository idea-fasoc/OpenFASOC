* NGSPICE file created from diff_pair_sample_1126.ext - technology: sky130A

.subckt diff_pair_sample_1126 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=0 ps=0 w=11.56 l=1.59
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=0 ps=0 w=11.56 l=1.59
X2 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=0 ps=0 w=11.56 l=1.59
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=0 ps=0 w=11.56 l=1.59
X4 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=4.5084 ps=23.9 w=11.56 l=1.59
X5 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=4.5084 ps=23.9 w=11.56 l=1.59
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=4.5084 ps=23.9 w=11.56 l=1.59
X7 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5084 pd=23.9 as=4.5084 ps=23.9 w=11.56 l=1.59
R0 B.n615 B.n614 585
R1 B.n263 B.n83 585
R2 B.n262 B.n261 585
R3 B.n260 B.n259 585
R4 B.n258 B.n257 585
R5 B.n256 B.n255 585
R6 B.n254 B.n253 585
R7 B.n252 B.n251 585
R8 B.n250 B.n249 585
R9 B.n248 B.n247 585
R10 B.n246 B.n245 585
R11 B.n244 B.n243 585
R12 B.n242 B.n241 585
R13 B.n240 B.n239 585
R14 B.n238 B.n237 585
R15 B.n236 B.n235 585
R16 B.n234 B.n233 585
R17 B.n232 B.n231 585
R18 B.n230 B.n229 585
R19 B.n228 B.n227 585
R20 B.n226 B.n225 585
R21 B.n224 B.n223 585
R22 B.n222 B.n221 585
R23 B.n220 B.n219 585
R24 B.n218 B.n217 585
R25 B.n216 B.n215 585
R26 B.n214 B.n213 585
R27 B.n212 B.n211 585
R28 B.n210 B.n209 585
R29 B.n208 B.n207 585
R30 B.n206 B.n205 585
R31 B.n204 B.n203 585
R32 B.n202 B.n201 585
R33 B.n200 B.n199 585
R34 B.n198 B.n197 585
R35 B.n196 B.n195 585
R36 B.n194 B.n193 585
R37 B.n192 B.n191 585
R38 B.n190 B.n189 585
R39 B.n188 B.n187 585
R40 B.n186 B.n185 585
R41 B.n184 B.n183 585
R42 B.n182 B.n181 585
R43 B.n180 B.n179 585
R44 B.n178 B.n177 585
R45 B.n176 B.n175 585
R46 B.n174 B.n173 585
R47 B.n172 B.n171 585
R48 B.n170 B.n169 585
R49 B.n168 B.n167 585
R50 B.n166 B.n165 585
R51 B.n164 B.n163 585
R52 B.n162 B.n161 585
R53 B.n160 B.n159 585
R54 B.n158 B.n157 585
R55 B.n156 B.n155 585
R56 B.n154 B.n153 585
R57 B.n152 B.n151 585
R58 B.n150 B.n149 585
R59 B.n148 B.n147 585
R60 B.n146 B.n145 585
R61 B.n144 B.n143 585
R62 B.n142 B.n141 585
R63 B.n140 B.n139 585
R64 B.n138 B.n137 585
R65 B.n136 B.n135 585
R66 B.n134 B.n133 585
R67 B.n132 B.n131 585
R68 B.n130 B.n129 585
R69 B.n128 B.n127 585
R70 B.n126 B.n125 585
R71 B.n124 B.n123 585
R72 B.n122 B.n121 585
R73 B.n120 B.n119 585
R74 B.n118 B.n117 585
R75 B.n116 B.n115 585
R76 B.n114 B.n113 585
R77 B.n112 B.n111 585
R78 B.n110 B.n109 585
R79 B.n108 B.n107 585
R80 B.n106 B.n105 585
R81 B.n104 B.n103 585
R82 B.n102 B.n101 585
R83 B.n100 B.n99 585
R84 B.n98 B.n97 585
R85 B.n96 B.n95 585
R86 B.n94 B.n93 585
R87 B.n92 B.n91 585
R88 B.n39 B.n38 585
R89 B.n620 B.n619 585
R90 B.n613 B.n84 585
R91 B.n84 B.n36 585
R92 B.n612 B.n35 585
R93 B.n624 B.n35 585
R94 B.n611 B.n34 585
R95 B.n625 B.n34 585
R96 B.n610 B.n33 585
R97 B.n626 B.n33 585
R98 B.n609 B.n608 585
R99 B.n608 B.n29 585
R100 B.n607 B.n28 585
R101 B.n632 B.n28 585
R102 B.n606 B.n27 585
R103 B.n633 B.n27 585
R104 B.n605 B.n26 585
R105 B.n634 B.n26 585
R106 B.n604 B.n603 585
R107 B.n603 B.n22 585
R108 B.n602 B.n21 585
R109 B.n640 B.n21 585
R110 B.n601 B.n20 585
R111 B.n641 B.n20 585
R112 B.n600 B.n19 585
R113 B.n642 B.n19 585
R114 B.n599 B.n598 585
R115 B.n598 B.n15 585
R116 B.n597 B.n14 585
R117 B.n648 B.n14 585
R118 B.n596 B.n13 585
R119 B.n649 B.n13 585
R120 B.n595 B.n12 585
R121 B.n650 B.n12 585
R122 B.n594 B.n593 585
R123 B.n593 B.n592 585
R124 B.n591 B.n590 585
R125 B.n591 B.n8 585
R126 B.n589 B.n7 585
R127 B.n657 B.n7 585
R128 B.n588 B.n6 585
R129 B.n658 B.n6 585
R130 B.n587 B.n5 585
R131 B.n659 B.n5 585
R132 B.n586 B.n585 585
R133 B.n585 B.n4 585
R134 B.n584 B.n264 585
R135 B.n584 B.n583 585
R136 B.n574 B.n265 585
R137 B.n266 B.n265 585
R138 B.n576 B.n575 585
R139 B.n577 B.n576 585
R140 B.n573 B.n271 585
R141 B.n271 B.n270 585
R142 B.n572 B.n571 585
R143 B.n571 B.n570 585
R144 B.n273 B.n272 585
R145 B.n274 B.n273 585
R146 B.n563 B.n562 585
R147 B.n564 B.n563 585
R148 B.n561 B.n279 585
R149 B.n279 B.n278 585
R150 B.n560 B.n559 585
R151 B.n559 B.n558 585
R152 B.n281 B.n280 585
R153 B.n282 B.n281 585
R154 B.n551 B.n550 585
R155 B.n552 B.n551 585
R156 B.n549 B.n286 585
R157 B.n290 B.n286 585
R158 B.n548 B.n547 585
R159 B.n547 B.n546 585
R160 B.n288 B.n287 585
R161 B.n289 B.n288 585
R162 B.n539 B.n538 585
R163 B.n540 B.n539 585
R164 B.n537 B.n295 585
R165 B.n295 B.n294 585
R166 B.n536 B.n535 585
R167 B.n535 B.n534 585
R168 B.n297 B.n296 585
R169 B.n298 B.n297 585
R170 B.n530 B.n529 585
R171 B.n301 B.n300 585
R172 B.n526 B.n525 585
R173 B.n527 B.n526 585
R174 B.n524 B.n346 585
R175 B.n523 B.n522 585
R176 B.n521 B.n520 585
R177 B.n519 B.n518 585
R178 B.n517 B.n516 585
R179 B.n515 B.n514 585
R180 B.n513 B.n512 585
R181 B.n511 B.n510 585
R182 B.n509 B.n508 585
R183 B.n507 B.n506 585
R184 B.n505 B.n504 585
R185 B.n503 B.n502 585
R186 B.n501 B.n500 585
R187 B.n499 B.n498 585
R188 B.n497 B.n496 585
R189 B.n495 B.n494 585
R190 B.n493 B.n492 585
R191 B.n491 B.n490 585
R192 B.n489 B.n488 585
R193 B.n487 B.n486 585
R194 B.n485 B.n484 585
R195 B.n483 B.n482 585
R196 B.n481 B.n480 585
R197 B.n479 B.n478 585
R198 B.n477 B.n476 585
R199 B.n475 B.n474 585
R200 B.n473 B.n472 585
R201 B.n471 B.n470 585
R202 B.n469 B.n468 585
R203 B.n467 B.n466 585
R204 B.n465 B.n464 585
R205 B.n463 B.n462 585
R206 B.n461 B.n460 585
R207 B.n459 B.n458 585
R208 B.n457 B.n456 585
R209 B.n455 B.n454 585
R210 B.n453 B.n452 585
R211 B.n450 B.n449 585
R212 B.n448 B.n447 585
R213 B.n446 B.n445 585
R214 B.n444 B.n443 585
R215 B.n442 B.n441 585
R216 B.n440 B.n439 585
R217 B.n438 B.n437 585
R218 B.n436 B.n435 585
R219 B.n434 B.n433 585
R220 B.n432 B.n431 585
R221 B.n429 B.n428 585
R222 B.n427 B.n426 585
R223 B.n425 B.n424 585
R224 B.n423 B.n422 585
R225 B.n421 B.n420 585
R226 B.n419 B.n418 585
R227 B.n417 B.n416 585
R228 B.n415 B.n414 585
R229 B.n413 B.n412 585
R230 B.n411 B.n410 585
R231 B.n409 B.n408 585
R232 B.n407 B.n406 585
R233 B.n405 B.n404 585
R234 B.n403 B.n402 585
R235 B.n401 B.n400 585
R236 B.n399 B.n398 585
R237 B.n397 B.n396 585
R238 B.n395 B.n394 585
R239 B.n393 B.n392 585
R240 B.n391 B.n390 585
R241 B.n389 B.n388 585
R242 B.n387 B.n386 585
R243 B.n385 B.n384 585
R244 B.n383 B.n382 585
R245 B.n381 B.n380 585
R246 B.n379 B.n378 585
R247 B.n377 B.n376 585
R248 B.n375 B.n374 585
R249 B.n373 B.n372 585
R250 B.n371 B.n370 585
R251 B.n369 B.n368 585
R252 B.n367 B.n366 585
R253 B.n365 B.n364 585
R254 B.n363 B.n362 585
R255 B.n361 B.n360 585
R256 B.n359 B.n358 585
R257 B.n357 B.n356 585
R258 B.n355 B.n354 585
R259 B.n353 B.n352 585
R260 B.n351 B.n345 585
R261 B.n527 B.n345 585
R262 B.n531 B.n299 585
R263 B.n299 B.n298 585
R264 B.n533 B.n532 585
R265 B.n534 B.n533 585
R266 B.n293 B.n292 585
R267 B.n294 B.n293 585
R268 B.n542 B.n541 585
R269 B.n541 B.n540 585
R270 B.n543 B.n291 585
R271 B.n291 B.n289 585
R272 B.n545 B.n544 585
R273 B.n546 B.n545 585
R274 B.n285 B.n284 585
R275 B.n290 B.n285 585
R276 B.n554 B.n553 585
R277 B.n553 B.n552 585
R278 B.n555 B.n283 585
R279 B.n283 B.n282 585
R280 B.n557 B.n556 585
R281 B.n558 B.n557 585
R282 B.n277 B.n276 585
R283 B.n278 B.n277 585
R284 B.n566 B.n565 585
R285 B.n565 B.n564 585
R286 B.n567 B.n275 585
R287 B.n275 B.n274 585
R288 B.n569 B.n568 585
R289 B.n570 B.n569 585
R290 B.n269 B.n268 585
R291 B.n270 B.n269 585
R292 B.n579 B.n578 585
R293 B.n578 B.n577 585
R294 B.n580 B.n267 585
R295 B.n267 B.n266 585
R296 B.n582 B.n581 585
R297 B.n583 B.n582 585
R298 B.n3 B.n0 585
R299 B.n4 B.n3 585
R300 B.n656 B.n1 585
R301 B.n657 B.n656 585
R302 B.n655 B.n654 585
R303 B.n655 B.n8 585
R304 B.n653 B.n9 585
R305 B.n592 B.n9 585
R306 B.n652 B.n651 585
R307 B.n651 B.n650 585
R308 B.n11 B.n10 585
R309 B.n649 B.n11 585
R310 B.n647 B.n646 585
R311 B.n648 B.n647 585
R312 B.n645 B.n16 585
R313 B.n16 B.n15 585
R314 B.n644 B.n643 585
R315 B.n643 B.n642 585
R316 B.n18 B.n17 585
R317 B.n641 B.n18 585
R318 B.n639 B.n638 585
R319 B.n640 B.n639 585
R320 B.n637 B.n23 585
R321 B.n23 B.n22 585
R322 B.n636 B.n635 585
R323 B.n635 B.n634 585
R324 B.n25 B.n24 585
R325 B.n633 B.n25 585
R326 B.n631 B.n630 585
R327 B.n632 B.n631 585
R328 B.n629 B.n30 585
R329 B.n30 B.n29 585
R330 B.n628 B.n627 585
R331 B.n627 B.n626 585
R332 B.n32 B.n31 585
R333 B.n625 B.n32 585
R334 B.n623 B.n622 585
R335 B.n624 B.n623 585
R336 B.n621 B.n37 585
R337 B.n37 B.n36 585
R338 B.n660 B.n659 585
R339 B.n658 B.n2 585
R340 B.n619 B.n37 502.111
R341 B.n615 B.n84 502.111
R342 B.n345 B.n297 502.111
R343 B.n529 B.n299 502.111
R344 B.n88 B.t6 380.978
R345 B.n85 B.t2 380.978
R346 B.n349 B.t13 380.978
R347 B.n347 B.t9 380.978
R348 B.n617 B.n616 256.663
R349 B.n617 B.n82 256.663
R350 B.n617 B.n81 256.663
R351 B.n617 B.n80 256.663
R352 B.n617 B.n79 256.663
R353 B.n617 B.n78 256.663
R354 B.n617 B.n77 256.663
R355 B.n617 B.n76 256.663
R356 B.n617 B.n75 256.663
R357 B.n617 B.n74 256.663
R358 B.n617 B.n73 256.663
R359 B.n617 B.n72 256.663
R360 B.n617 B.n71 256.663
R361 B.n617 B.n70 256.663
R362 B.n617 B.n69 256.663
R363 B.n617 B.n68 256.663
R364 B.n617 B.n67 256.663
R365 B.n617 B.n66 256.663
R366 B.n617 B.n65 256.663
R367 B.n617 B.n64 256.663
R368 B.n617 B.n63 256.663
R369 B.n617 B.n62 256.663
R370 B.n617 B.n61 256.663
R371 B.n617 B.n60 256.663
R372 B.n617 B.n59 256.663
R373 B.n617 B.n58 256.663
R374 B.n617 B.n57 256.663
R375 B.n617 B.n56 256.663
R376 B.n617 B.n55 256.663
R377 B.n617 B.n54 256.663
R378 B.n617 B.n53 256.663
R379 B.n617 B.n52 256.663
R380 B.n617 B.n51 256.663
R381 B.n617 B.n50 256.663
R382 B.n617 B.n49 256.663
R383 B.n617 B.n48 256.663
R384 B.n617 B.n47 256.663
R385 B.n617 B.n46 256.663
R386 B.n617 B.n45 256.663
R387 B.n617 B.n44 256.663
R388 B.n617 B.n43 256.663
R389 B.n617 B.n42 256.663
R390 B.n617 B.n41 256.663
R391 B.n617 B.n40 256.663
R392 B.n618 B.n617 256.663
R393 B.n528 B.n527 256.663
R394 B.n527 B.n302 256.663
R395 B.n527 B.n303 256.663
R396 B.n527 B.n304 256.663
R397 B.n527 B.n305 256.663
R398 B.n527 B.n306 256.663
R399 B.n527 B.n307 256.663
R400 B.n527 B.n308 256.663
R401 B.n527 B.n309 256.663
R402 B.n527 B.n310 256.663
R403 B.n527 B.n311 256.663
R404 B.n527 B.n312 256.663
R405 B.n527 B.n313 256.663
R406 B.n527 B.n314 256.663
R407 B.n527 B.n315 256.663
R408 B.n527 B.n316 256.663
R409 B.n527 B.n317 256.663
R410 B.n527 B.n318 256.663
R411 B.n527 B.n319 256.663
R412 B.n527 B.n320 256.663
R413 B.n527 B.n321 256.663
R414 B.n527 B.n322 256.663
R415 B.n527 B.n323 256.663
R416 B.n527 B.n324 256.663
R417 B.n527 B.n325 256.663
R418 B.n527 B.n326 256.663
R419 B.n527 B.n327 256.663
R420 B.n527 B.n328 256.663
R421 B.n527 B.n329 256.663
R422 B.n527 B.n330 256.663
R423 B.n527 B.n331 256.663
R424 B.n527 B.n332 256.663
R425 B.n527 B.n333 256.663
R426 B.n527 B.n334 256.663
R427 B.n527 B.n335 256.663
R428 B.n527 B.n336 256.663
R429 B.n527 B.n337 256.663
R430 B.n527 B.n338 256.663
R431 B.n527 B.n339 256.663
R432 B.n527 B.n340 256.663
R433 B.n527 B.n341 256.663
R434 B.n527 B.n342 256.663
R435 B.n527 B.n343 256.663
R436 B.n527 B.n344 256.663
R437 B.n662 B.n661 256.663
R438 B.n91 B.n39 163.367
R439 B.n95 B.n94 163.367
R440 B.n99 B.n98 163.367
R441 B.n103 B.n102 163.367
R442 B.n107 B.n106 163.367
R443 B.n111 B.n110 163.367
R444 B.n115 B.n114 163.367
R445 B.n119 B.n118 163.367
R446 B.n123 B.n122 163.367
R447 B.n127 B.n126 163.367
R448 B.n131 B.n130 163.367
R449 B.n135 B.n134 163.367
R450 B.n139 B.n138 163.367
R451 B.n143 B.n142 163.367
R452 B.n147 B.n146 163.367
R453 B.n151 B.n150 163.367
R454 B.n155 B.n154 163.367
R455 B.n159 B.n158 163.367
R456 B.n163 B.n162 163.367
R457 B.n167 B.n166 163.367
R458 B.n171 B.n170 163.367
R459 B.n175 B.n174 163.367
R460 B.n179 B.n178 163.367
R461 B.n183 B.n182 163.367
R462 B.n187 B.n186 163.367
R463 B.n191 B.n190 163.367
R464 B.n195 B.n194 163.367
R465 B.n199 B.n198 163.367
R466 B.n203 B.n202 163.367
R467 B.n207 B.n206 163.367
R468 B.n211 B.n210 163.367
R469 B.n215 B.n214 163.367
R470 B.n219 B.n218 163.367
R471 B.n223 B.n222 163.367
R472 B.n227 B.n226 163.367
R473 B.n231 B.n230 163.367
R474 B.n235 B.n234 163.367
R475 B.n239 B.n238 163.367
R476 B.n243 B.n242 163.367
R477 B.n247 B.n246 163.367
R478 B.n251 B.n250 163.367
R479 B.n255 B.n254 163.367
R480 B.n259 B.n258 163.367
R481 B.n261 B.n83 163.367
R482 B.n535 B.n297 163.367
R483 B.n535 B.n295 163.367
R484 B.n539 B.n295 163.367
R485 B.n539 B.n288 163.367
R486 B.n547 B.n288 163.367
R487 B.n547 B.n286 163.367
R488 B.n551 B.n286 163.367
R489 B.n551 B.n281 163.367
R490 B.n559 B.n281 163.367
R491 B.n559 B.n279 163.367
R492 B.n563 B.n279 163.367
R493 B.n563 B.n273 163.367
R494 B.n571 B.n273 163.367
R495 B.n571 B.n271 163.367
R496 B.n576 B.n271 163.367
R497 B.n576 B.n265 163.367
R498 B.n584 B.n265 163.367
R499 B.n585 B.n584 163.367
R500 B.n585 B.n5 163.367
R501 B.n6 B.n5 163.367
R502 B.n7 B.n6 163.367
R503 B.n591 B.n7 163.367
R504 B.n593 B.n591 163.367
R505 B.n593 B.n12 163.367
R506 B.n13 B.n12 163.367
R507 B.n14 B.n13 163.367
R508 B.n598 B.n14 163.367
R509 B.n598 B.n19 163.367
R510 B.n20 B.n19 163.367
R511 B.n21 B.n20 163.367
R512 B.n603 B.n21 163.367
R513 B.n603 B.n26 163.367
R514 B.n27 B.n26 163.367
R515 B.n28 B.n27 163.367
R516 B.n608 B.n28 163.367
R517 B.n608 B.n33 163.367
R518 B.n34 B.n33 163.367
R519 B.n35 B.n34 163.367
R520 B.n84 B.n35 163.367
R521 B.n526 B.n301 163.367
R522 B.n526 B.n346 163.367
R523 B.n522 B.n521 163.367
R524 B.n518 B.n517 163.367
R525 B.n514 B.n513 163.367
R526 B.n510 B.n509 163.367
R527 B.n506 B.n505 163.367
R528 B.n502 B.n501 163.367
R529 B.n498 B.n497 163.367
R530 B.n494 B.n493 163.367
R531 B.n490 B.n489 163.367
R532 B.n486 B.n485 163.367
R533 B.n482 B.n481 163.367
R534 B.n478 B.n477 163.367
R535 B.n474 B.n473 163.367
R536 B.n470 B.n469 163.367
R537 B.n466 B.n465 163.367
R538 B.n462 B.n461 163.367
R539 B.n458 B.n457 163.367
R540 B.n454 B.n453 163.367
R541 B.n449 B.n448 163.367
R542 B.n445 B.n444 163.367
R543 B.n441 B.n440 163.367
R544 B.n437 B.n436 163.367
R545 B.n433 B.n432 163.367
R546 B.n428 B.n427 163.367
R547 B.n424 B.n423 163.367
R548 B.n420 B.n419 163.367
R549 B.n416 B.n415 163.367
R550 B.n412 B.n411 163.367
R551 B.n408 B.n407 163.367
R552 B.n404 B.n403 163.367
R553 B.n400 B.n399 163.367
R554 B.n396 B.n395 163.367
R555 B.n392 B.n391 163.367
R556 B.n388 B.n387 163.367
R557 B.n384 B.n383 163.367
R558 B.n380 B.n379 163.367
R559 B.n376 B.n375 163.367
R560 B.n372 B.n371 163.367
R561 B.n368 B.n367 163.367
R562 B.n364 B.n363 163.367
R563 B.n360 B.n359 163.367
R564 B.n356 B.n355 163.367
R565 B.n352 B.n345 163.367
R566 B.n533 B.n299 163.367
R567 B.n533 B.n293 163.367
R568 B.n541 B.n293 163.367
R569 B.n541 B.n291 163.367
R570 B.n545 B.n291 163.367
R571 B.n545 B.n285 163.367
R572 B.n553 B.n285 163.367
R573 B.n553 B.n283 163.367
R574 B.n557 B.n283 163.367
R575 B.n557 B.n277 163.367
R576 B.n565 B.n277 163.367
R577 B.n565 B.n275 163.367
R578 B.n569 B.n275 163.367
R579 B.n569 B.n269 163.367
R580 B.n578 B.n269 163.367
R581 B.n578 B.n267 163.367
R582 B.n582 B.n267 163.367
R583 B.n582 B.n3 163.367
R584 B.n660 B.n3 163.367
R585 B.n656 B.n2 163.367
R586 B.n656 B.n655 163.367
R587 B.n655 B.n9 163.367
R588 B.n651 B.n9 163.367
R589 B.n651 B.n11 163.367
R590 B.n647 B.n11 163.367
R591 B.n647 B.n16 163.367
R592 B.n643 B.n16 163.367
R593 B.n643 B.n18 163.367
R594 B.n639 B.n18 163.367
R595 B.n639 B.n23 163.367
R596 B.n635 B.n23 163.367
R597 B.n635 B.n25 163.367
R598 B.n631 B.n25 163.367
R599 B.n631 B.n30 163.367
R600 B.n627 B.n30 163.367
R601 B.n627 B.n32 163.367
R602 B.n623 B.n32 163.367
R603 B.n623 B.n37 163.367
R604 B.n85 B.t4 105.088
R605 B.n349 B.t15 105.088
R606 B.n88 B.t7 105.073
R607 B.n347 B.t12 105.073
R608 B.n527 B.n298 76.4484
R609 B.n617 B.n36 76.4484
R610 B.n619 B.n618 71.676
R611 B.n91 B.n40 71.676
R612 B.n95 B.n41 71.676
R613 B.n99 B.n42 71.676
R614 B.n103 B.n43 71.676
R615 B.n107 B.n44 71.676
R616 B.n111 B.n45 71.676
R617 B.n115 B.n46 71.676
R618 B.n119 B.n47 71.676
R619 B.n123 B.n48 71.676
R620 B.n127 B.n49 71.676
R621 B.n131 B.n50 71.676
R622 B.n135 B.n51 71.676
R623 B.n139 B.n52 71.676
R624 B.n143 B.n53 71.676
R625 B.n147 B.n54 71.676
R626 B.n151 B.n55 71.676
R627 B.n155 B.n56 71.676
R628 B.n159 B.n57 71.676
R629 B.n163 B.n58 71.676
R630 B.n167 B.n59 71.676
R631 B.n171 B.n60 71.676
R632 B.n175 B.n61 71.676
R633 B.n179 B.n62 71.676
R634 B.n183 B.n63 71.676
R635 B.n187 B.n64 71.676
R636 B.n191 B.n65 71.676
R637 B.n195 B.n66 71.676
R638 B.n199 B.n67 71.676
R639 B.n203 B.n68 71.676
R640 B.n207 B.n69 71.676
R641 B.n211 B.n70 71.676
R642 B.n215 B.n71 71.676
R643 B.n219 B.n72 71.676
R644 B.n223 B.n73 71.676
R645 B.n227 B.n74 71.676
R646 B.n231 B.n75 71.676
R647 B.n235 B.n76 71.676
R648 B.n239 B.n77 71.676
R649 B.n243 B.n78 71.676
R650 B.n247 B.n79 71.676
R651 B.n251 B.n80 71.676
R652 B.n255 B.n81 71.676
R653 B.n259 B.n82 71.676
R654 B.n616 B.n83 71.676
R655 B.n616 B.n615 71.676
R656 B.n261 B.n82 71.676
R657 B.n258 B.n81 71.676
R658 B.n254 B.n80 71.676
R659 B.n250 B.n79 71.676
R660 B.n246 B.n78 71.676
R661 B.n242 B.n77 71.676
R662 B.n238 B.n76 71.676
R663 B.n234 B.n75 71.676
R664 B.n230 B.n74 71.676
R665 B.n226 B.n73 71.676
R666 B.n222 B.n72 71.676
R667 B.n218 B.n71 71.676
R668 B.n214 B.n70 71.676
R669 B.n210 B.n69 71.676
R670 B.n206 B.n68 71.676
R671 B.n202 B.n67 71.676
R672 B.n198 B.n66 71.676
R673 B.n194 B.n65 71.676
R674 B.n190 B.n64 71.676
R675 B.n186 B.n63 71.676
R676 B.n182 B.n62 71.676
R677 B.n178 B.n61 71.676
R678 B.n174 B.n60 71.676
R679 B.n170 B.n59 71.676
R680 B.n166 B.n58 71.676
R681 B.n162 B.n57 71.676
R682 B.n158 B.n56 71.676
R683 B.n154 B.n55 71.676
R684 B.n150 B.n54 71.676
R685 B.n146 B.n53 71.676
R686 B.n142 B.n52 71.676
R687 B.n138 B.n51 71.676
R688 B.n134 B.n50 71.676
R689 B.n130 B.n49 71.676
R690 B.n126 B.n48 71.676
R691 B.n122 B.n47 71.676
R692 B.n118 B.n46 71.676
R693 B.n114 B.n45 71.676
R694 B.n110 B.n44 71.676
R695 B.n106 B.n43 71.676
R696 B.n102 B.n42 71.676
R697 B.n98 B.n41 71.676
R698 B.n94 B.n40 71.676
R699 B.n618 B.n39 71.676
R700 B.n529 B.n528 71.676
R701 B.n346 B.n302 71.676
R702 B.n521 B.n303 71.676
R703 B.n517 B.n304 71.676
R704 B.n513 B.n305 71.676
R705 B.n509 B.n306 71.676
R706 B.n505 B.n307 71.676
R707 B.n501 B.n308 71.676
R708 B.n497 B.n309 71.676
R709 B.n493 B.n310 71.676
R710 B.n489 B.n311 71.676
R711 B.n485 B.n312 71.676
R712 B.n481 B.n313 71.676
R713 B.n477 B.n314 71.676
R714 B.n473 B.n315 71.676
R715 B.n469 B.n316 71.676
R716 B.n465 B.n317 71.676
R717 B.n461 B.n318 71.676
R718 B.n457 B.n319 71.676
R719 B.n453 B.n320 71.676
R720 B.n448 B.n321 71.676
R721 B.n444 B.n322 71.676
R722 B.n440 B.n323 71.676
R723 B.n436 B.n324 71.676
R724 B.n432 B.n325 71.676
R725 B.n427 B.n326 71.676
R726 B.n423 B.n327 71.676
R727 B.n419 B.n328 71.676
R728 B.n415 B.n329 71.676
R729 B.n411 B.n330 71.676
R730 B.n407 B.n331 71.676
R731 B.n403 B.n332 71.676
R732 B.n399 B.n333 71.676
R733 B.n395 B.n334 71.676
R734 B.n391 B.n335 71.676
R735 B.n387 B.n336 71.676
R736 B.n383 B.n337 71.676
R737 B.n379 B.n338 71.676
R738 B.n375 B.n339 71.676
R739 B.n371 B.n340 71.676
R740 B.n367 B.n341 71.676
R741 B.n363 B.n342 71.676
R742 B.n359 B.n343 71.676
R743 B.n355 B.n344 71.676
R744 B.n528 B.n301 71.676
R745 B.n522 B.n302 71.676
R746 B.n518 B.n303 71.676
R747 B.n514 B.n304 71.676
R748 B.n510 B.n305 71.676
R749 B.n506 B.n306 71.676
R750 B.n502 B.n307 71.676
R751 B.n498 B.n308 71.676
R752 B.n494 B.n309 71.676
R753 B.n490 B.n310 71.676
R754 B.n486 B.n311 71.676
R755 B.n482 B.n312 71.676
R756 B.n478 B.n313 71.676
R757 B.n474 B.n314 71.676
R758 B.n470 B.n315 71.676
R759 B.n466 B.n316 71.676
R760 B.n462 B.n317 71.676
R761 B.n458 B.n318 71.676
R762 B.n454 B.n319 71.676
R763 B.n449 B.n320 71.676
R764 B.n445 B.n321 71.676
R765 B.n441 B.n322 71.676
R766 B.n437 B.n323 71.676
R767 B.n433 B.n324 71.676
R768 B.n428 B.n325 71.676
R769 B.n424 B.n326 71.676
R770 B.n420 B.n327 71.676
R771 B.n416 B.n328 71.676
R772 B.n412 B.n329 71.676
R773 B.n408 B.n330 71.676
R774 B.n404 B.n331 71.676
R775 B.n400 B.n332 71.676
R776 B.n396 B.n333 71.676
R777 B.n392 B.n334 71.676
R778 B.n388 B.n335 71.676
R779 B.n384 B.n336 71.676
R780 B.n380 B.n337 71.676
R781 B.n376 B.n338 71.676
R782 B.n372 B.n339 71.676
R783 B.n368 B.n340 71.676
R784 B.n364 B.n341 71.676
R785 B.n360 B.n342 71.676
R786 B.n356 B.n343 71.676
R787 B.n352 B.n344 71.676
R788 B.n661 B.n660 71.676
R789 B.n661 B.n2 71.676
R790 B.n86 B.t5 67.8522
R791 B.n350 B.t14 67.8522
R792 B.n89 B.t8 67.8375
R793 B.n348 B.t11 67.8375
R794 B.n90 B.n89 59.5399
R795 B.n87 B.n86 59.5399
R796 B.n430 B.n350 59.5399
R797 B.n451 B.n348 59.5399
R798 B.n534 B.n298 44.4317
R799 B.n534 B.n294 44.4317
R800 B.n540 B.n294 44.4317
R801 B.n540 B.n289 44.4317
R802 B.n546 B.n289 44.4317
R803 B.n546 B.n290 44.4317
R804 B.n552 B.n282 44.4317
R805 B.n558 B.n282 44.4317
R806 B.n558 B.n278 44.4317
R807 B.n564 B.n278 44.4317
R808 B.n564 B.n274 44.4317
R809 B.n570 B.n274 44.4317
R810 B.n570 B.n270 44.4317
R811 B.n577 B.n270 44.4317
R812 B.n583 B.n266 44.4317
R813 B.n583 B.n4 44.4317
R814 B.n659 B.n4 44.4317
R815 B.n659 B.n658 44.4317
R816 B.n658 B.n657 44.4317
R817 B.n657 B.n8 44.4317
R818 B.n592 B.n8 44.4317
R819 B.n650 B.n649 44.4317
R820 B.n649 B.n648 44.4317
R821 B.n648 B.n15 44.4317
R822 B.n642 B.n15 44.4317
R823 B.n642 B.n641 44.4317
R824 B.n641 B.n640 44.4317
R825 B.n640 B.n22 44.4317
R826 B.n634 B.n22 44.4317
R827 B.n633 B.n632 44.4317
R828 B.n632 B.n29 44.4317
R829 B.n626 B.n29 44.4317
R830 B.n626 B.n625 44.4317
R831 B.n625 B.n624 44.4317
R832 B.n624 B.n36 44.4317
R833 B.t0 B.n266 41.1647
R834 B.n592 B.t1 41.1647
R835 B.n89 B.n88 37.2369
R836 B.n86 B.n85 37.2369
R837 B.n350 B.n349 37.2369
R838 B.n348 B.n347 37.2369
R839 B.n552 B.t10 34.6307
R840 B.n634 B.t3 34.6307
R841 B.n531 B.n530 32.6249
R842 B.n351 B.n296 32.6249
R843 B.n614 B.n613 32.6249
R844 B.n621 B.n620 32.6249
R845 B B.n662 18.0485
R846 B.n532 B.n531 10.6151
R847 B.n532 B.n292 10.6151
R848 B.n542 B.n292 10.6151
R849 B.n543 B.n542 10.6151
R850 B.n544 B.n543 10.6151
R851 B.n544 B.n284 10.6151
R852 B.n554 B.n284 10.6151
R853 B.n555 B.n554 10.6151
R854 B.n556 B.n555 10.6151
R855 B.n556 B.n276 10.6151
R856 B.n566 B.n276 10.6151
R857 B.n567 B.n566 10.6151
R858 B.n568 B.n567 10.6151
R859 B.n568 B.n268 10.6151
R860 B.n579 B.n268 10.6151
R861 B.n580 B.n579 10.6151
R862 B.n581 B.n580 10.6151
R863 B.n581 B.n0 10.6151
R864 B.n530 B.n300 10.6151
R865 B.n525 B.n300 10.6151
R866 B.n525 B.n524 10.6151
R867 B.n524 B.n523 10.6151
R868 B.n523 B.n520 10.6151
R869 B.n520 B.n519 10.6151
R870 B.n519 B.n516 10.6151
R871 B.n516 B.n515 10.6151
R872 B.n515 B.n512 10.6151
R873 B.n512 B.n511 10.6151
R874 B.n511 B.n508 10.6151
R875 B.n508 B.n507 10.6151
R876 B.n507 B.n504 10.6151
R877 B.n504 B.n503 10.6151
R878 B.n503 B.n500 10.6151
R879 B.n500 B.n499 10.6151
R880 B.n499 B.n496 10.6151
R881 B.n496 B.n495 10.6151
R882 B.n495 B.n492 10.6151
R883 B.n492 B.n491 10.6151
R884 B.n491 B.n488 10.6151
R885 B.n488 B.n487 10.6151
R886 B.n487 B.n484 10.6151
R887 B.n484 B.n483 10.6151
R888 B.n483 B.n480 10.6151
R889 B.n480 B.n479 10.6151
R890 B.n479 B.n476 10.6151
R891 B.n476 B.n475 10.6151
R892 B.n475 B.n472 10.6151
R893 B.n472 B.n471 10.6151
R894 B.n471 B.n468 10.6151
R895 B.n468 B.n467 10.6151
R896 B.n467 B.n464 10.6151
R897 B.n464 B.n463 10.6151
R898 B.n463 B.n460 10.6151
R899 B.n460 B.n459 10.6151
R900 B.n459 B.n456 10.6151
R901 B.n456 B.n455 10.6151
R902 B.n455 B.n452 10.6151
R903 B.n450 B.n447 10.6151
R904 B.n447 B.n446 10.6151
R905 B.n446 B.n443 10.6151
R906 B.n443 B.n442 10.6151
R907 B.n442 B.n439 10.6151
R908 B.n439 B.n438 10.6151
R909 B.n438 B.n435 10.6151
R910 B.n435 B.n434 10.6151
R911 B.n434 B.n431 10.6151
R912 B.n429 B.n426 10.6151
R913 B.n426 B.n425 10.6151
R914 B.n425 B.n422 10.6151
R915 B.n422 B.n421 10.6151
R916 B.n421 B.n418 10.6151
R917 B.n418 B.n417 10.6151
R918 B.n417 B.n414 10.6151
R919 B.n414 B.n413 10.6151
R920 B.n413 B.n410 10.6151
R921 B.n410 B.n409 10.6151
R922 B.n409 B.n406 10.6151
R923 B.n406 B.n405 10.6151
R924 B.n405 B.n402 10.6151
R925 B.n402 B.n401 10.6151
R926 B.n401 B.n398 10.6151
R927 B.n398 B.n397 10.6151
R928 B.n397 B.n394 10.6151
R929 B.n394 B.n393 10.6151
R930 B.n393 B.n390 10.6151
R931 B.n390 B.n389 10.6151
R932 B.n389 B.n386 10.6151
R933 B.n386 B.n385 10.6151
R934 B.n385 B.n382 10.6151
R935 B.n382 B.n381 10.6151
R936 B.n381 B.n378 10.6151
R937 B.n378 B.n377 10.6151
R938 B.n377 B.n374 10.6151
R939 B.n374 B.n373 10.6151
R940 B.n373 B.n370 10.6151
R941 B.n370 B.n369 10.6151
R942 B.n369 B.n366 10.6151
R943 B.n366 B.n365 10.6151
R944 B.n365 B.n362 10.6151
R945 B.n362 B.n361 10.6151
R946 B.n361 B.n358 10.6151
R947 B.n358 B.n357 10.6151
R948 B.n357 B.n354 10.6151
R949 B.n354 B.n353 10.6151
R950 B.n353 B.n351 10.6151
R951 B.n536 B.n296 10.6151
R952 B.n537 B.n536 10.6151
R953 B.n538 B.n537 10.6151
R954 B.n538 B.n287 10.6151
R955 B.n548 B.n287 10.6151
R956 B.n549 B.n548 10.6151
R957 B.n550 B.n549 10.6151
R958 B.n550 B.n280 10.6151
R959 B.n560 B.n280 10.6151
R960 B.n561 B.n560 10.6151
R961 B.n562 B.n561 10.6151
R962 B.n562 B.n272 10.6151
R963 B.n572 B.n272 10.6151
R964 B.n573 B.n572 10.6151
R965 B.n575 B.n573 10.6151
R966 B.n575 B.n574 10.6151
R967 B.n574 B.n264 10.6151
R968 B.n586 B.n264 10.6151
R969 B.n587 B.n586 10.6151
R970 B.n588 B.n587 10.6151
R971 B.n589 B.n588 10.6151
R972 B.n590 B.n589 10.6151
R973 B.n594 B.n590 10.6151
R974 B.n595 B.n594 10.6151
R975 B.n596 B.n595 10.6151
R976 B.n597 B.n596 10.6151
R977 B.n599 B.n597 10.6151
R978 B.n600 B.n599 10.6151
R979 B.n601 B.n600 10.6151
R980 B.n602 B.n601 10.6151
R981 B.n604 B.n602 10.6151
R982 B.n605 B.n604 10.6151
R983 B.n606 B.n605 10.6151
R984 B.n607 B.n606 10.6151
R985 B.n609 B.n607 10.6151
R986 B.n610 B.n609 10.6151
R987 B.n611 B.n610 10.6151
R988 B.n612 B.n611 10.6151
R989 B.n613 B.n612 10.6151
R990 B.n654 B.n1 10.6151
R991 B.n654 B.n653 10.6151
R992 B.n653 B.n652 10.6151
R993 B.n652 B.n10 10.6151
R994 B.n646 B.n10 10.6151
R995 B.n646 B.n645 10.6151
R996 B.n645 B.n644 10.6151
R997 B.n644 B.n17 10.6151
R998 B.n638 B.n17 10.6151
R999 B.n638 B.n637 10.6151
R1000 B.n637 B.n636 10.6151
R1001 B.n636 B.n24 10.6151
R1002 B.n630 B.n24 10.6151
R1003 B.n630 B.n629 10.6151
R1004 B.n629 B.n628 10.6151
R1005 B.n628 B.n31 10.6151
R1006 B.n622 B.n31 10.6151
R1007 B.n622 B.n621 10.6151
R1008 B.n620 B.n38 10.6151
R1009 B.n92 B.n38 10.6151
R1010 B.n93 B.n92 10.6151
R1011 B.n96 B.n93 10.6151
R1012 B.n97 B.n96 10.6151
R1013 B.n100 B.n97 10.6151
R1014 B.n101 B.n100 10.6151
R1015 B.n104 B.n101 10.6151
R1016 B.n105 B.n104 10.6151
R1017 B.n108 B.n105 10.6151
R1018 B.n109 B.n108 10.6151
R1019 B.n112 B.n109 10.6151
R1020 B.n113 B.n112 10.6151
R1021 B.n116 B.n113 10.6151
R1022 B.n117 B.n116 10.6151
R1023 B.n120 B.n117 10.6151
R1024 B.n121 B.n120 10.6151
R1025 B.n124 B.n121 10.6151
R1026 B.n125 B.n124 10.6151
R1027 B.n128 B.n125 10.6151
R1028 B.n129 B.n128 10.6151
R1029 B.n132 B.n129 10.6151
R1030 B.n133 B.n132 10.6151
R1031 B.n136 B.n133 10.6151
R1032 B.n137 B.n136 10.6151
R1033 B.n140 B.n137 10.6151
R1034 B.n141 B.n140 10.6151
R1035 B.n144 B.n141 10.6151
R1036 B.n145 B.n144 10.6151
R1037 B.n148 B.n145 10.6151
R1038 B.n149 B.n148 10.6151
R1039 B.n152 B.n149 10.6151
R1040 B.n153 B.n152 10.6151
R1041 B.n156 B.n153 10.6151
R1042 B.n157 B.n156 10.6151
R1043 B.n160 B.n157 10.6151
R1044 B.n161 B.n160 10.6151
R1045 B.n164 B.n161 10.6151
R1046 B.n165 B.n164 10.6151
R1047 B.n169 B.n168 10.6151
R1048 B.n172 B.n169 10.6151
R1049 B.n173 B.n172 10.6151
R1050 B.n176 B.n173 10.6151
R1051 B.n177 B.n176 10.6151
R1052 B.n180 B.n177 10.6151
R1053 B.n181 B.n180 10.6151
R1054 B.n184 B.n181 10.6151
R1055 B.n185 B.n184 10.6151
R1056 B.n189 B.n188 10.6151
R1057 B.n192 B.n189 10.6151
R1058 B.n193 B.n192 10.6151
R1059 B.n196 B.n193 10.6151
R1060 B.n197 B.n196 10.6151
R1061 B.n200 B.n197 10.6151
R1062 B.n201 B.n200 10.6151
R1063 B.n204 B.n201 10.6151
R1064 B.n205 B.n204 10.6151
R1065 B.n208 B.n205 10.6151
R1066 B.n209 B.n208 10.6151
R1067 B.n212 B.n209 10.6151
R1068 B.n213 B.n212 10.6151
R1069 B.n216 B.n213 10.6151
R1070 B.n217 B.n216 10.6151
R1071 B.n220 B.n217 10.6151
R1072 B.n221 B.n220 10.6151
R1073 B.n224 B.n221 10.6151
R1074 B.n225 B.n224 10.6151
R1075 B.n228 B.n225 10.6151
R1076 B.n229 B.n228 10.6151
R1077 B.n232 B.n229 10.6151
R1078 B.n233 B.n232 10.6151
R1079 B.n236 B.n233 10.6151
R1080 B.n237 B.n236 10.6151
R1081 B.n240 B.n237 10.6151
R1082 B.n241 B.n240 10.6151
R1083 B.n244 B.n241 10.6151
R1084 B.n245 B.n244 10.6151
R1085 B.n248 B.n245 10.6151
R1086 B.n249 B.n248 10.6151
R1087 B.n252 B.n249 10.6151
R1088 B.n253 B.n252 10.6151
R1089 B.n256 B.n253 10.6151
R1090 B.n257 B.n256 10.6151
R1091 B.n260 B.n257 10.6151
R1092 B.n262 B.n260 10.6151
R1093 B.n263 B.n262 10.6151
R1094 B.n614 B.n263 10.6151
R1095 B.n290 B.t10 9.80151
R1096 B.t3 B.n633 9.80151
R1097 B.n452 B.n451 9.36635
R1098 B.n430 B.n429 9.36635
R1099 B.n165 B.n90 9.36635
R1100 B.n188 B.n87 9.36635
R1101 B.n662 B.n0 8.11757
R1102 B.n662 B.n1 8.11757
R1103 B.n577 B.t0 3.2675
R1104 B.n650 B.t1 3.2675
R1105 B.n451 B.n450 1.24928
R1106 B.n431 B.n430 1.24928
R1107 B.n168 B.n90 1.24928
R1108 B.n185 B.n87 1.24928
R1109 VP.n0 VP.t1 322.476
R1110 VP.n0 VP.t0 280.83
R1111 VP VP.n0 0.146778
R1112 VTAIL.n1 VTAIL.t0 49.4681
R1113 VTAIL.n3 VTAIL.t1 49.4671
R1114 VTAIL.n0 VTAIL.t3 49.4671
R1115 VTAIL.n2 VTAIL.t2 49.467
R1116 VTAIL.n1 VTAIL.n0 25.6427
R1117 VTAIL.n3 VTAIL.n2 23.9876
R1118 VTAIL.n2 VTAIL.n1 1.29791
R1119 VTAIL VTAIL.n0 0.94231
R1120 VTAIL VTAIL.n3 0.356103
R1121 VDD1 VDD1.t1 104.019
R1122 VDD1 VDD1.t0 66.6177
R1123 VN VN.t0 322.762
R1124 VN VN.t1 280.978
R1125 VDD2.n0 VDD2.t0 103.082
R1126 VDD2.n0 VDD2.t1 66.1458
R1127 VDD2 VDD2.n0 0.472483
C0 VP VTAIL 2.08058f
C1 VN VDD2 2.44857f
C2 VDD2 VDD1 0.556215f
C3 VP VDD2 0.29037f
C4 VN VDD1 0.147325f
C5 VN VP 4.8988f
C6 VP VDD1 2.58849f
C7 VDD2 VTAIL 4.96179f
C8 VN VTAIL 2.06619f
C9 VTAIL VDD1 4.91929f
C10 VDD2 B 3.996558f
C11 VDD1 B 6.86986f
C12 VTAIL B 6.673841f
C13 VN B 9.523129f
C14 VP B 5.093344f
C15 VDD2.t0 B 2.56832f
C16 VDD2.t1 B 2.10129f
C17 VDD2.n0 B 2.64522f
C18 VN.t1 B 2.36647f
C19 VN.t0 B 2.66632f
C20 VDD1.t0 B 2.11019f
C21 VDD1.t1 B 2.60595f
C22 VTAIL.t3 B 2.0743f
C23 VTAIL.n0 B 1.48207f
C24 VTAIL.t0 B 2.0743f
C25 VTAIL.n1 B 1.5057f
C26 VTAIL.t2 B 2.07429f
C27 VTAIL.n2 B 1.3957f
C28 VTAIL.t1 B 2.0743f
C29 VTAIL.n3 B 1.3331f
C30 VP.t1 B 2.7348f
C31 VP.t0 B 2.4312f
C32 VP.n0 B 4.38851f
.ends

