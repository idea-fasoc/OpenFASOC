* NGSPICE file created from diff_pair_sample_0528.ext - technology: sky130A

.subckt diff_pair_sample_0528 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=3.6192 ps=19.34 w=9.28 l=2.56
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=3.6192 ps=19.34 w=9.28 l=2.56
X2 B.t11 B.t9 B.t10 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=0 ps=0 w=9.28 l=2.56
X3 VDD2.t0 VN.t1 VTAIL.t2 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=3.6192 ps=19.34 w=9.28 l=2.56
X4 B.t8 B.t6 B.t7 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=0 ps=0 w=9.28 l=2.56
X5 B.t5 B.t3 B.t4 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=0 ps=0 w=9.28 l=2.56
X6 B.t2 B.t0 B.t1 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=0 ps=0 w=9.28 l=2.56
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n2126_n2824# sky130_fd_pr__pfet_01v8 ad=3.6192 pd=19.34 as=3.6192 ps=19.34 w=9.28 l=2.56
R0 VN VN.t1 179.165
R1 VN VN.t0 136.915
R2 VTAIL.n194 VTAIL.n150 756.745
R3 VTAIL.n44 VTAIL.n0 756.745
R4 VTAIL.n144 VTAIL.n100 756.745
R5 VTAIL.n94 VTAIL.n50 756.745
R6 VTAIL.n167 VTAIL.n166 585
R7 VTAIL.n169 VTAIL.n168 585
R8 VTAIL.n162 VTAIL.n161 585
R9 VTAIL.n175 VTAIL.n174 585
R10 VTAIL.n177 VTAIL.n176 585
R11 VTAIL.n158 VTAIL.n157 585
R12 VTAIL.n184 VTAIL.n183 585
R13 VTAIL.n185 VTAIL.n156 585
R14 VTAIL.n187 VTAIL.n186 585
R15 VTAIL.n154 VTAIL.n153 585
R16 VTAIL.n193 VTAIL.n192 585
R17 VTAIL.n195 VTAIL.n194 585
R18 VTAIL.n17 VTAIL.n16 585
R19 VTAIL.n19 VTAIL.n18 585
R20 VTAIL.n12 VTAIL.n11 585
R21 VTAIL.n25 VTAIL.n24 585
R22 VTAIL.n27 VTAIL.n26 585
R23 VTAIL.n8 VTAIL.n7 585
R24 VTAIL.n34 VTAIL.n33 585
R25 VTAIL.n35 VTAIL.n6 585
R26 VTAIL.n37 VTAIL.n36 585
R27 VTAIL.n4 VTAIL.n3 585
R28 VTAIL.n43 VTAIL.n42 585
R29 VTAIL.n45 VTAIL.n44 585
R30 VTAIL.n145 VTAIL.n144 585
R31 VTAIL.n143 VTAIL.n142 585
R32 VTAIL.n104 VTAIL.n103 585
R33 VTAIL.n108 VTAIL.n106 585
R34 VTAIL.n137 VTAIL.n136 585
R35 VTAIL.n135 VTAIL.n134 585
R36 VTAIL.n110 VTAIL.n109 585
R37 VTAIL.n129 VTAIL.n128 585
R38 VTAIL.n127 VTAIL.n126 585
R39 VTAIL.n114 VTAIL.n113 585
R40 VTAIL.n121 VTAIL.n120 585
R41 VTAIL.n119 VTAIL.n118 585
R42 VTAIL.n95 VTAIL.n94 585
R43 VTAIL.n93 VTAIL.n92 585
R44 VTAIL.n54 VTAIL.n53 585
R45 VTAIL.n58 VTAIL.n56 585
R46 VTAIL.n87 VTAIL.n86 585
R47 VTAIL.n85 VTAIL.n84 585
R48 VTAIL.n60 VTAIL.n59 585
R49 VTAIL.n79 VTAIL.n78 585
R50 VTAIL.n77 VTAIL.n76 585
R51 VTAIL.n64 VTAIL.n63 585
R52 VTAIL.n71 VTAIL.n70 585
R53 VTAIL.n69 VTAIL.n68 585
R54 VTAIL.n165 VTAIL.t3 329.038
R55 VTAIL.n15 VTAIL.t1 329.038
R56 VTAIL.n117 VTAIL.t0 329.038
R57 VTAIL.n67 VTAIL.t2 329.038
R58 VTAIL.n168 VTAIL.n167 171.744
R59 VTAIL.n168 VTAIL.n161 171.744
R60 VTAIL.n175 VTAIL.n161 171.744
R61 VTAIL.n176 VTAIL.n175 171.744
R62 VTAIL.n176 VTAIL.n157 171.744
R63 VTAIL.n184 VTAIL.n157 171.744
R64 VTAIL.n185 VTAIL.n184 171.744
R65 VTAIL.n186 VTAIL.n185 171.744
R66 VTAIL.n186 VTAIL.n153 171.744
R67 VTAIL.n193 VTAIL.n153 171.744
R68 VTAIL.n194 VTAIL.n193 171.744
R69 VTAIL.n18 VTAIL.n17 171.744
R70 VTAIL.n18 VTAIL.n11 171.744
R71 VTAIL.n25 VTAIL.n11 171.744
R72 VTAIL.n26 VTAIL.n25 171.744
R73 VTAIL.n26 VTAIL.n7 171.744
R74 VTAIL.n34 VTAIL.n7 171.744
R75 VTAIL.n35 VTAIL.n34 171.744
R76 VTAIL.n36 VTAIL.n35 171.744
R77 VTAIL.n36 VTAIL.n3 171.744
R78 VTAIL.n43 VTAIL.n3 171.744
R79 VTAIL.n44 VTAIL.n43 171.744
R80 VTAIL.n144 VTAIL.n143 171.744
R81 VTAIL.n143 VTAIL.n103 171.744
R82 VTAIL.n108 VTAIL.n103 171.744
R83 VTAIL.n136 VTAIL.n108 171.744
R84 VTAIL.n136 VTAIL.n135 171.744
R85 VTAIL.n135 VTAIL.n109 171.744
R86 VTAIL.n128 VTAIL.n109 171.744
R87 VTAIL.n128 VTAIL.n127 171.744
R88 VTAIL.n127 VTAIL.n113 171.744
R89 VTAIL.n120 VTAIL.n113 171.744
R90 VTAIL.n120 VTAIL.n119 171.744
R91 VTAIL.n94 VTAIL.n93 171.744
R92 VTAIL.n93 VTAIL.n53 171.744
R93 VTAIL.n58 VTAIL.n53 171.744
R94 VTAIL.n86 VTAIL.n58 171.744
R95 VTAIL.n86 VTAIL.n85 171.744
R96 VTAIL.n85 VTAIL.n59 171.744
R97 VTAIL.n78 VTAIL.n59 171.744
R98 VTAIL.n78 VTAIL.n77 171.744
R99 VTAIL.n77 VTAIL.n63 171.744
R100 VTAIL.n70 VTAIL.n63 171.744
R101 VTAIL.n70 VTAIL.n69 171.744
R102 VTAIL.n167 VTAIL.t3 85.8723
R103 VTAIL.n17 VTAIL.t1 85.8723
R104 VTAIL.n119 VTAIL.t0 85.8723
R105 VTAIL.n69 VTAIL.t2 85.8723
R106 VTAIL.n199 VTAIL.n198 32.9611
R107 VTAIL.n49 VTAIL.n48 32.9611
R108 VTAIL.n149 VTAIL.n148 32.9611
R109 VTAIL.n99 VTAIL.n98 32.9611
R110 VTAIL.n99 VTAIL.n49 25.3496
R111 VTAIL.n199 VTAIL.n149 22.8583
R112 VTAIL.n187 VTAIL.n154 13.1884
R113 VTAIL.n37 VTAIL.n4 13.1884
R114 VTAIL.n106 VTAIL.n104 13.1884
R115 VTAIL.n56 VTAIL.n54 13.1884
R116 VTAIL.n188 VTAIL.n156 12.8005
R117 VTAIL.n192 VTAIL.n191 12.8005
R118 VTAIL.n38 VTAIL.n6 12.8005
R119 VTAIL.n42 VTAIL.n41 12.8005
R120 VTAIL.n142 VTAIL.n141 12.8005
R121 VTAIL.n138 VTAIL.n137 12.8005
R122 VTAIL.n92 VTAIL.n91 12.8005
R123 VTAIL.n88 VTAIL.n87 12.8005
R124 VTAIL.n183 VTAIL.n182 12.0247
R125 VTAIL.n195 VTAIL.n152 12.0247
R126 VTAIL.n33 VTAIL.n32 12.0247
R127 VTAIL.n45 VTAIL.n2 12.0247
R128 VTAIL.n145 VTAIL.n102 12.0247
R129 VTAIL.n134 VTAIL.n107 12.0247
R130 VTAIL.n95 VTAIL.n52 12.0247
R131 VTAIL.n84 VTAIL.n57 12.0247
R132 VTAIL.n181 VTAIL.n158 11.249
R133 VTAIL.n196 VTAIL.n150 11.249
R134 VTAIL.n31 VTAIL.n8 11.249
R135 VTAIL.n46 VTAIL.n0 11.249
R136 VTAIL.n146 VTAIL.n100 11.249
R137 VTAIL.n133 VTAIL.n110 11.249
R138 VTAIL.n96 VTAIL.n50 11.249
R139 VTAIL.n83 VTAIL.n60 11.249
R140 VTAIL.n166 VTAIL.n165 10.7239
R141 VTAIL.n16 VTAIL.n15 10.7239
R142 VTAIL.n118 VTAIL.n117 10.7239
R143 VTAIL.n68 VTAIL.n67 10.7239
R144 VTAIL.n178 VTAIL.n177 10.4732
R145 VTAIL.n28 VTAIL.n27 10.4732
R146 VTAIL.n130 VTAIL.n129 10.4732
R147 VTAIL.n80 VTAIL.n79 10.4732
R148 VTAIL.n174 VTAIL.n160 9.69747
R149 VTAIL.n24 VTAIL.n10 9.69747
R150 VTAIL.n126 VTAIL.n112 9.69747
R151 VTAIL.n76 VTAIL.n62 9.69747
R152 VTAIL.n198 VTAIL.n197 9.45567
R153 VTAIL.n48 VTAIL.n47 9.45567
R154 VTAIL.n148 VTAIL.n147 9.45567
R155 VTAIL.n98 VTAIL.n97 9.45567
R156 VTAIL.n197 VTAIL.n196 9.3005
R157 VTAIL.n152 VTAIL.n151 9.3005
R158 VTAIL.n191 VTAIL.n190 9.3005
R159 VTAIL.n164 VTAIL.n163 9.3005
R160 VTAIL.n171 VTAIL.n170 9.3005
R161 VTAIL.n173 VTAIL.n172 9.3005
R162 VTAIL.n160 VTAIL.n159 9.3005
R163 VTAIL.n179 VTAIL.n178 9.3005
R164 VTAIL.n181 VTAIL.n180 9.3005
R165 VTAIL.n182 VTAIL.n155 9.3005
R166 VTAIL.n189 VTAIL.n188 9.3005
R167 VTAIL.n47 VTAIL.n46 9.3005
R168 VTAIL.n2 VTAIL.n1 9.3005
R169 VTAIL.n41 VTAIL.n40 9.3005
R170 VTAIL.n14 VTAIL.n13 9.3005
R171 VTAIL.n21 VTAIL.n20 9.3005
R172 VTAIL.n23 VTAIL.n22 9.3005
R173 VTAIL.n10 VTAIL.n9 9.3005
R174 VTAIL.n29 VTAIL.n28 9.3005
R175 VTAIL.n31 VTAIL.n30 9.3005
R176 VTAIL.n32 VTAIL.n5 9.3005
R177 VTAIL.n39 VTAIL.n38 9.3005
R178 VTAIL.n116 VTAIL.n115 9.3005
R179 VTAIL.n123 VTAIL.n122 9.3005
R180 VTAIL.n125 VTAIL.n124 9.3005
R181 VTAIL.n112 VTAIL.n111 9.3005
R182 VTAIL.n131 VTAIL.n130 9.3005
R183 VTAIL.n133 VTAIL.n132 9.3005
R184 VTAIL.n107 VTAIL.n105 9.3005
R185 VTAIL.n139 VTAIL.n138 9.3005
R186 VTAIL.n147 VTAIL.n146 9.3005
R187 VTAIL.n102 VTAIL.n101 9.3005
R188 VTAIL.n141 VTAIL.n140 9.3005
R189 VTAIL.n66 VTAIL.n65 9.3005
R190 VTAIL.n73 VTAIL.n72 9.3005
R191 VTAIL.n75 VTAIL.n74 9.3005
R192 VTAIL.n62 VTAIL.n61 9.3005
R193 VTAIL.n81 VTAIL.n80 9.3005
R194 VTAIL.n83 VTAIL.n82 9.3005
R195 VTAIL.n57 VTAIL.n55 9.3005
R196 VTAIL.n89 VTAIL.n88 9.3005
R197 VTAIL.n97 VTAIL.n96 9.3005
R198 VTAIL.n52 VTAIL.n51 9.3005
R199 VTAIL.n91 VTAIL.n90 9.3005
R200 VTAIL.n173 VTAIL.n162 8.92171
R201 VTAIL.n23 VTAIL.n12 8.92171
R202 VTAIL.n125 VTAIL.n114 8.92171
R203 VTAIL.n75 VTAIL.n64 8.92171
R204 VTAIL.n170 VTAIL.n169 8.14595
R205 VTAIL.n20 VTAIL.n19 8.14595
R206 VTAIL.n122 VTAIL.n121 8.14595
R207 VTAIL.n72 VTAIL.n71 8.14595
R208 VTAIL.n166 VTAIL.n164 7.3702
R209 VTAIL.n16 VTAIL.n14 7.3702
R210 VTAIL.n118 VTAIL.n116 7.3702
R211 VTAIL.n68 VTAIL.n66 7.3702
R212 VTAIL.n169 VTAIL.n164 5.81868
R213 VTAIL.n19 VTAIL.n14 5.81868
R214 VTAIL.n121 VTAIL.n116 5.81868
R215 VTAIL.n71 VTAIL.n66 5.81868
R216 VTAIL.n170 VTAIL.n162 5.04292
R217 VTAIL.n20 VTAIL.n12 5.04292
R218 VTAIL.n122 VTAIL.n114 5.04292
R219 VTAIL.n72 VTAIL.n64 5.04292
R220 VTAIL.n174 VTAIL.n173 4.26717
R221 VTAIL.n24 VTAIL.n23 4.26717
R222 VTAIL.n126 VTAIL.n125 4.26717
R223 VTAIL.n76 VTAIL.n75 4.26717
R224 VTAIL.n177 VTAIL.n160 3.49141
R225 VTAIL.n27 VTAIL.n10 3.49141
R226 VTAIL.n129 VTAIL.n112 3.49141
R227 VTAIL.n79 VTAIL.n62 3.49141
R228 VTAIL.n178 VTAIL.n158 2.71565
R229 VTAIL.n198 VTAIL.n150 2.71565
R230 VTAIL.n28 VTAIL.n8 2.71565
R231 VTAIL.n48 VTAIL.n0 2.71565
R232 VTAIL.n148 VTAIL.n100 2.71565
R233 VTAIL.n130 VTAIL.n110 2.71565
R234 VTAIL.n98 VTAIL.n50 2.71565
R235 VTAIL.n80 VTAIL.n60 2.71565
R236 VTAIL.n165 VTAIL.n163 2.41283
R237 VTAIL.n15 VTAIL.n13 2.41283
R238 VTAIL.n117 VTAIL.n115 2.41283
R239 VTAIL.n67 VTAIL.n65 2.41283
R240 VTAIL.n183 VTAIL.n181 1.93989
R241 VTAIL.n196 VTAIL.n195 1.93989
R242 VTAIL.n33 VTAIL.n31 1.93989
R243 VTAIL.n46 VTAIL.n45 1.93989
R244 VTAIL.n146 VTAIL.n145 1.93989
R245 VTAIL.n134 VTAIL.n133 1.93989
R246 VTAIL.n96 VTAIL.n95 1.93989
R247 VTAIL.n84 VTAIL.n83 1.93989
R248 VTAIL.n149 VTAIL.n99 1.71602
R249 VTAIL.n182 VTAIL.n156 1.16414
R250 VTAIL.n192 VTAIL.n152 1.16414
R251 VTAIL.n32 VTAIL.n6 1.16414
R252 VTAIL.n42 VTAIL.n2 1.16414
R253 VTAIL.n142 VTAIL.n102 1.16414
R254 VTAIL.n137 VTAIL.n107 1.16414
R255 VTAIL.n92 VTAIL.n52 1.16414
R256 VTAIL.n87 VTAIL.n57 1.16414
R257 VTAIL VTAIL.n49 1.15136
R258 VTAIL VTAIL.n199 0.565155
R259 VTAIL.n188 VTAIL.n187 0.388379
R260 VTAIL.n191 VTAIL.n154 0.388379
R261 VTAIL.n38 VTAIL.n37 0.388379
R262 VTAIL.n41 VTAIL.n4 0.388379
R263 VTAIL.n141 VTAIL.n104 0.388379
R264 VTAIL.n138 VTAIL.n106 0.388379
R265 VTAIL.n91 VTAIL.n54 0.388379
R266 VTAIL.n88 VTAIL.n56 0.388379
R267 VTAIL.n171 VTAIL.n163 0.155672
R268 VTAIL.n172 VTAIL.n171 0.155672
R269 VTAIL.n172 VTAIL.n159 0.155672
R270 VTAIL.n179 VTAIL.n159 0.155672
R271 VTAIL.n180 VTAIL.n179 0.155672
R272 VTAIL.n180 VTAIL.n155 0.155672
R273 VTAIL.n189 VTAIL.n155 0.155672
R274 VTAIL.n190 VTAIL.n189 0.155672
R275 VTAIL.n190 VTAIL.n151 0.155672
R276 VTAIL.n197 VTAIL.n151 0.155672
R277 VTAIL.n21 VTAIL.n13 0.155672
R278 VTAIL.n22 VTAIL.n21 0.155672
R279 VTAIL.n22 VTAIL.n9 0.155672
R280 VTAIL.n29 VTAIL.n9 0.155672
R281 VTAIL.n30 VTAIL.n29 0.155672
R282 VTAIL.n30 VTAIL.n5 0.155672
R283 VTAIL.n39 VTAIL.n5 0.155672
R284 VTAIL.n40 VTAIL.n39 0.155672
R285 VTAIL.n40 VTAIL.n1 0.155672
R286 VTAIL.n47 VTAIL.n1 0.155672
R287 VTAIL.n147 VTAIL.n101 0.155672
R288 VTAIL.n140 VTAIL.n101 0.155672
R289 VTAIL.n140 VTAIL.n139 0.155672
R290 VTAIL.n139 VTAIL.n105 0.155672
R291 VTAIL.n132 VTAIL.n105 0.155672
R292 VTAIL.n132 VTAIL.n131 0.155672
R293 VTAIL.n131 VTAIL.n111 0.155672
R294 VTAIL.n124 VTAIL.n111 0.155672
R295 VTAIL.n124 VTAIL.n123 0.155672
R296 VTAIL.n123 VTAIL.n115 0.155672
R297 VTAIL.n97 VTAIL.n51 0.155672
R298 VTAIL.n90 VTAIL.n51 0.155672
R299 VTAIL.n90 VTAIL.n89 0.155672
R300 VTAIL.n89 VTAIL.n55 0.155672
R301 VTAIL.n82 VTAIL.n55 0.155672
R302 VTAIL.n82 VTAIL.n81 0.155672
R303 VTAIL.n81 VTAIL.n61 0.155672
R304 VTAIL.n74 VTAIL.n61 0.155672
R305 VTAIL.n74 VTAIL.n73 0.155672
R306 VTAIL.n73 VTAIL.n65 0.155672
R307 VDD2.n93 VDD2.n49 756.745
R308 VDD2.n44 VDD2.n0 756.745
R309 VDD2.n94 VDD2.n93 585
R310 VDD2.n92 VDD2.n91 585
R311 VDD2.n53 VDD2.n52 585
R312 VDD2.n57 VDD2.n55 585
R313 VDD2.n86 VDD2.n85 585
R314 VDD2.n84 VDD2.n83 585
R315 VDD2.n59 VDD2.n58 585
R316 VDD2.n78 VDD2.n77 585
R317 VDD2.n76 VDD2.n75 585
R318 VDD2.n63 VDD2.n62 585
R319 VDD2.n70 VDD2.n69 585
R320 VDD2.n68 VDD2.n67 585
R321 VDD2.n17 VDD2.n16 585
R322 VDD2.n19 VDD2.n18 585
R323 VDD2.n12 VDD2.n11 585
R324 VDD2.n25 VDD2.n24 585
R325 VDD2.n27 VDD2.n26 585
R326 VDD2.n8 VDD2.n7 585
R327 VDD2.n34 VDD2.n33 585
R328 VDD2.n35 VDD2.n6 585
R329 VDD2.n37 VDD2.n36 585
R330 VDD2.n4 VDD2.n3 585
R331 VDD2.n43 VDD2.n42 585
R332 VDD2.n45 VDD2.n44 585
R333 VDD2.n66 VDD2.t0 329.038
R334 VDD2.n15 VDD2.t1 329.038
R335 VDD2.n93 VDD2.n92 171.744
R336 VDD2.n92 VDD2.n52 171.744
R337 VDD2.n57 VDD2.n52 171.744
R338 VDD2.n85 VDD2.n57 171.744
R339 VDD2.n85 VDD2.n84 171.744
R340 VDD2.n84 VDD2.n58 171.744
R341 VDD2.n77 VDD2.n58 171.744
R342 VDD2.n77 VDD2.n76 171.744
R343 VDD2.n76 VDD2.n62 171.744
R344 VDD2.n69 VDD2.n62 171.744
R345 VDD2.n69 VDD2.n68 171.744
R346 VDD2.n18 VDD2.n17 171.744
R347 VDD2.n18 VDD2.n11 171.744
R348 VDD2.n25 VDD2.n11 171.744
R349 VDD2.n26 VDD2.n25 171.744
R350 VDD2.n26 VDD2.n7 171.744
R351 VDD2.n34 VDD2.n7 171.744
R352 VDD2.n35 VDD2.n34 171.744
R353 VDD2.n36 VDD2.n35 171.744
R354 VDD2.n36 VDD2.n3 171.744
R355 VDD2.n43 VDD2.n3 171.744
R356 VDD2.n44 VDD2.n43 171.744
R357 VDD2.n98 VDD2.n48 86.2821
R358 VDD2.n68 VDD2.t0 85.8723
R359 VDD2.n17 VDD2.t1 85.8723
R360 VDD2.n98 VDD2.n97 49.6399
R361 VDD2.n55 VDD2.n53 13.1884
R362 VDD2.n37 VDD2.n4 13.1884
R363 VDD2.n91 VDD2.n90 12.8005
R364 VDD2.n87 VDD2.n86 12.8005
R365 VDD2.n38 VDD2.n6 12.8005
R366 VDD2.n42 VDD2.n41 12.8005
R367 VDD2.n94 VDD2.n51 12.0247
R368 VDD2.n83 VDD2.n56 12.0247
R369 VDD2.n33 VDD2.n32 12.0247
R370 VDD2.n45 VDD2.n2 12.0247
R371 VDD2.n95 VDD2.n49 11.249
R372 VDD2.n82 VDD2.n59 11.249
R373 VDD2.n31 VDD2.n8 11.249
R374 VDD2.n46 VDD2.n0 11.249
R375 VDD2.n67 VDD2.n66 10.7239
R376 VDD2.n16 VDD2.n15 10.7239
R377 VDD2.n79 VDD2.n78 10.4732
R378 VDD2.n28 VDD2.n27 10.4732
R379 VDD2.n75 VDD2.n61 9.69747
R380 VDD2.n24 VDD2.n10 9.69747
R381 VDD2.n97 VDD2.n96 9.45567
R382 VDD2.n48 VDD2.n47 9.45567
R383 VDD2.n65 VDD2.n64 9.3005
R384 VDD2.n72 VDD2.n71 9.3005
R385 VDD2.n74 VDD2.n73 9.3005
R386 VDD2.n61 VDD2.n60 9.3005
R387 VDD2.n80 VDD2.n79 9.3005
R388 VDD2.n82 VDD2.n81 9.3005
R389 VDD2.n56 VDD2.n54 9.3005
R390 VDD2.n88 VDD2.n87 9.3005
R391 VDD2.n96 VDD2.n95 9.3005
R392 VDD2.n51 VDD2.n50 9.3005
R393 VDD2.n90 VDD2.n89 9.3005
R394 VDD2.n47 VDD2.n46 9.3005
R395 VDD2.n2 VDD2.n1 9.3005
R396 VDD2.n41 VDD2.n40 9.3005
R397 VDD2.n14 VDD2.n13 9.3005
R398 VDD2.n21 VDD2.n20 9.3005
R399 VDD2.n23 VDD2.n22 9.3005
R400 VDD2.n10 VDD2.n9 9.3005
R401 VDD2.n29 VDD2.n28 9.3005
R402 VDD2.n31 VDD2.n30 9.3005
R403 VDD2.n32 VDD2.n5 9.3005
R404 VDD2.n39 VDD2.n38 9.3005
R405 VDD2.n74 VDD2.n63 8.92171
R406 VDD2.n23 VDD2.n12 8.92171
R407 VDD2.n71 VDD2.n70 8.14595
R408 VDD2.n20 VDD2.n19 8.14595
R409 VDD2.n67 VDD2.n65 7.3702
R410 VDD2.n16 VDD2.n14 7.3702
R411 VDD2.n70 VDD2.n65 5.81868
R412 VDD2.n19 VDD2.n14 5.81868
R413 VDD2.n71 VDD2.n63 5.04292
R414 VDD2.n20 VDD2.n12 5.04292
R415 VDD2.n75 VDD2.n74 4.26717
R416 VDD2.n24 VDD2.n23 4.26717
R417 VDD2.n78 VDD2.n61 3.49141
R418 VDD2.n27 VDD2.n10 3.49141
R419 VDD2.n97 VDD2.n49 2.71565
R420 VDD2.n79 VDD2.n59 2.71565
R421 VDD2.n28 VDD2.n8 2.71565
R422 VDD2.n48 VDD2.n0 2.71565
R423 VDD2.n66 VDD2.n64 2.41283
R424 VDD2.n15 VDD2.n13 2.41283
R425 VDD2.n95 VDD2.n94 1.93989
R426 VDD2.n83 VDD2.n82 1.93989
R427 VDD2.n33 VDD2.n31 1.93989
R428 VDD2.n46 VDD2.n45 1.93989
R429 VDD2.n91 VDD2.n51 1.16414
R430 VDD2.n86 VDD2.n56 1.16414
R431 VDD2.n32 VDD2.n6 1.16414
R432 VDD2.n42 VDD2.n2 1.16414
R433 VDD2 VDD2.n98 0.681535
R434 VDD2.n90 VDD2.n53 0.388379
R435 VDD2.n87 VDD2.n55 0.388379
R436 VDD2.n38 VDD2.n37 0.388379
R437 VDD2.n41 VDD2.n4 0.388379
R438 VDD2.n96 VDD2.n50 0.155672
R439 VDD2.n89 VDD2.n50 0.155672
R440 VDD2.n89 VDD2.n88 0.155672
R441 VDD2.n88 VDD2.n54 0.155672
R442 VDD2.n81 VDD2.n54 0.155672
R443 VDD2.n81 VDD2.n80 0.155672
R444 VDD2.n80 VDD2.n60 0.155672
R445 VDD2.n73 VDD2.n60 0.155672
R446 VDD2.n73 VDD2.n72 0.155672
R447 VDD2.n72 VDD2.n64 0.155672
R448 VDD2.n21 VDD2.n13 0.155672
R449 VDD2.n22 VDD2.n21 0.155672
R450 VDD2.n22 VDD2.n9 0.155672
R451 VDD2.n29 VDD2.n9 0.155672
R452 VDD2.n30 VDD2.n29 0.155672
R453 VDD2.n30 VDD2.n5 0.155672
R454 VDD2.n39 VDD2.n5 0.155672
R455 VDD2.n40 VDD2.n39 0.155672
R456 VDD2.n40 VDD2.n1 0.155672
R457 VDD2.n47 VDD2.n1 0.155672
R458 VP.n0 VP.t1 179.067
R459 VP.n0 VP.t0 136.578
R460 VP VP.n0 0.336784
R461 VDD1.n44 VDD1.n0 756.745
R462 VDD1.n93 VDD1.n49 756.745
R463 VDD1.n45 VDD1.n44 585
R464 VDD1.n43 VDD1.n42 585
R465 VDD1.n4 VDD1.n3 585
R466 VDD1.n8 VDD1.n6 585
R467 VDD1.n37 VDD1.n36 585
R468 VDD1.n35 VDD1.n34 585
R469 VDD1.n10 VDD1.n9 585
R470 VDD1.n29 VDD1.n28 585
R471 VDD1.n27 VDD1.n26 585
R472 VDD1.n14 VDD1.n13 585
R473 VDD1.n21 VDD1.n20 585
R474 VDD1.n19 VDD1.n18 585
R475 VDD1.n66 VDD1.n65 585
R476 VDD1.n68 VDD1.n67 585
R477 VDD1.n61 VDD1.n60 585
R478 VDD1.n74 VDD1.n73 585
R479 VDD1.n76 VDD1.n75 585
R480 VDD1.n57 VDD1.n56 585
R481 VDD1.n83 VDD1.n82 585
R482 VDD1.n84 VDD1.n55 585
R483 VDD1.n86 VDD1.n85 585
R484 VDD1.n53 VDD1.n52 585
R485 VDD1.n92 VDD1.n91 585
R486 VDD1.n94 VDD1.n93 585
R487 VDD1.n17 VDD1.t0 329.038
R488 VDD1.n64 VDD1.t1 329.038
R489 VDD1.n44 VDD1.n43 171.744
R490 VDD1.n43 VDD1.n3 171.744
R491 VDD1.n8 VDD1.n3 171.744
R492 VDD1.n36 VDD1.n8 171.744
R493 VDD1.n36 VDD1.n35 171.744
R494 VDD1.n35 VDD1.n9 171.744
R495 VDD1.n28 VDD1.n9 171.744
R496 VDD1.n28 VDD1.n27 171.744
R497 VDD1.n27 VDD1.n13 171.744
R498 VDD1.n20 VDD1.n13 171.744
R499 VDD1.n20 VDD1.n19 171.744
R500 VDD1.n67 VDD1.n66 171.744
R501 VDD1.n67 VDD1.n60 171.744
R502 VDD1.n74 VDD1.n60 171.744
R503 VDD1.n75 VDD1.n74 171.744
R504 VDD1.n75 VDD1.n56 171.744
R505 VDD1.n83 VDD1.n56 171.744
R506 VDD1.n84 VDD1.n83 171.744
R507 VDD1.n85 VDD1.n84 171.744
R508 VDD1.n85 VDD1.n52 171.744
R509 VDD1.n92 VDD1.n52 171.744
R510 VDD1.n93 VDD1.n92 171.744
R511 VDD1 VDD1.n97 87.4298
R512 VDD1.n19 VDD1.t0 85.8723
R513 VDD1.n66 VDD1.t1 85.8723
R514 VDD1 VDD1.n48 50.3209
R515 VDD1.n6 VDD1.n4 13.1884
R516 VDD1.n86 VDD1.n53 13.1884
R517 VDD1.n42 VDD1.n41 12.8005
R518 VDD1.n38 VDD1.n37 12.8005
R519 VDD1.n87 VDD1.n55 12.8005
R520 VDD1.n91 VDD1.n90 12.8005
R521 VDD1.n45 VDD1.n2 12.0247
R522 VDD1.n34 VDD1.n7 12.0247
R523 VDD1.n82 VDD1.n81 12.0247
R524 VDD1.n94 VDD1.n51 12.0247
R525 VDD1.n46 VDD1.n0 11.249
R526 VDD1.n33 VDD1.n10 11.249
R527 VDD1.n80 VDD1.n57 11.249
R528 VDD1.n95 VDD1.n49 11.249
R529 VDD1.n18 VDD1.n17 10.7239
R530 VDD1.n65 VDD1.n64 10.7239
R531 VDD1.n30 VDD1.n29 10.4732
R532 VDD1.n77 VDD1.n76 10.4732
R533 VDD1.n26 VDD1.n12 9.69747
R534 VDD1.n73 VDD1.n59 9.69747
R535 VDD1.n48 VDD1.n47 9.45567
R536 VDD1.n97 VDD1.n96 9.45567
R537 VDD1.n16 VDD1.n15 9.3005
R538 VDD1.n23 VDD1.n22 9.3005
R539 VDD1.n25 VDD1.n24 9.3005
R540 VDD1.n12 VDD1.n11 9.3005
R541 VDD1.n31 VDD1.n30 9.3005
R542 VDD1.n33 VDD1.n32 9.3005
R543 VDD1.n7 VDD1.n5 9.3005
R544 VDD1.n39 VDD1.n38 9.3005
R545 VDD1.n47 VDD1.n46 9.3005
R546 VDD1.n2 VDD1.n1 9.3005
R547 VDD1.n41 VDD1.n40 9.3005
R548 VDD1.n96 VDD1.n95 9.3005
R549 VDD1.n51 VDD1.n50 9.3005
R550 VDD1.n90 VDD1.n89 9.3005
R551 VDD1.n63 VDD1.n62 9.3005
R552 VDD1.n70 VDD1.n69 9.3005
R553 VDD1.n72 VDD1.n71 9.3005
R554 VDD1.n59 VDD1.n58 9.3005
R555 VDD1.n78 VDD1.n77 9.3005
R556 VDD1.n80 VDD1.n79 9.3005
R557 VDD1.n81 VDD1.n54 9.3005
R558 VDD1.n88 VDD1.n87 9.3005
R559 VDD1.n25 VDD1.n14 8.92171
R560 VDD1.n72 VDD1.n61 8.92171
R561 VDD1.n22 VDD1.n21 8.14595
R562 VDD1.n69 VDD1.n68 8.14595
R563 VDD1.n18 VDD1.n16 7.3702
R564 VDD1.n65 VDD1.n63 7.3702
R565 VDD1.n21 VDD1.n16 5.81868
R566 VDD1.n68 VDD1.n63 5.81868
R567 VDD1.n22 VDD1.n14 5.04292
R568 VDD1.n69 VDD1.n61 5.04292
R569 VDD1.n26 VDD1.n25 4.26717
R570 VDD1.n73 VDD1.n72 4.26717
R571 VDD1.n29 VDD1.n12 3.49141
R572 VDD1.n76 VDD1.n59 3.49141
R573 VDD1.n48 VDD1.n0 2.71565
R574 VDD1.n30 VDD1.n10 2.71565
R575 VDD1.n77 VDD1.n57 2.71565
R576 VDD1.n97 VDD1.n49 2.71565
R577 VDD1.n17 VDD1.n15 2.41283
R578 VDD1.n64 VDD1.n62 2.41283
R579 VDD1.n46 VDD1.n45 1.93989
R580 VDD1.n34 VDD1.n33 1.93989
R581 VDD1.n82 VDD1.n80 1.93989
R582 VDD1.n95 VDD1.n94 1.93989
R583 VDD1.n42 VDD1.n2 1.16414
R584 VDD1.n37 VDD1.n7 1.16414
R585 VDD1.n81 VDD1.n55 1.16414
R586 VDD1.n91 VDD1.n51 1.16414
R587 VDD1.n41 VDD1.n4 0.388379
R588 VDD1.n38 VDD1.n6 0.388379
R589 VDD1.n87 VDD1.n86 0.388379
R590 VDD1.n90 VDD1.n53 0.388379
R591 VDD1.n47 VDD1.n1 0.155672
R592 VDD1.n40 VDD1.n1 0.155672
R593 VDD1.n40 VDD1.n39 0.155672
R594 VDD1.n39 VDD1.n5 0.155672
R595 VDD1.n32 VDD1.n5 0.155672
R596 VDD1.n32 VDD1.n31 0.155672
R597 VDD1.n31 VDD1.n11 0.155672
R598 VDD1.n24 VDD1.n11 0.155672
R599 VDD1.n24 VDD1.n23 0.155672
R600 VDD1.n23 VDD1.n15 0.155672
R601 VDD1.n70 VDD1.n62 0.155672
R602 VDD1.n71 VDD1.n70 0.155672
R603 VDD1.n71 VDD1.n58 0.155672
R604 VDD1.n78 VDD1.n58 0.155672
R605 VDD1.n79 VDD1.n78 0.155672
R606 VDD1.n79 VDD1.n54 0.155672
R607 VDD1.n88 VDD1.n54 0.155672
R608 VDD1.n89 VDD1.n88 0.155672
R609 VDD1.n89 VDD1.n50 0.155672
R610 VDD1.n96 VDD1.n50 0.155672
R611 B.n368 B.n57 585
R612 B.n370 B.n369 585
R613 B.n371 B.n56 585
R614 B.n373 B.n372 585
R615 B.n374 B.n55 585
R616 B.n376 B.n375 585
R617 B.n377 B.n54 585
R618 B.n379 B.n378 585
R619 B.n380 B.n53 585
R620 B.n382 B.n381 585
R621 B.n383 B.n52 585
R622 B.n385 B.n384 585
R623 B.n386 B.n51 585
R624 B.n388 B.n387 585
R625 B.n389 B.n50 585
R626 B.n391 B.n390 585
R627 B.n392 B.n49 585
R628 B.n394 B.n393 585
R629 B.n395 B.n48 585
R630 B.n397 B.n396 585
R631 B.n398 B.n47 585
R632 B.n400 B.n399 585
R633 B.n401 B.n46 585
R634 B.n403 B.n402 585
R635 B.n404 B.n45 585
R636 B.n406 B.n405 585
R637 B.n407 B.n44 585
R638 B.n409 B.n408 585
R639 B.n410 B.n43 585
R640 B.n412 B.n411 585
R641 B.n413 B.n42 585
R642 B.n415 B.n414 585
R643 B.n416 B.n41 585
R644 B.n418 B.n417 585
R645 B.n420 B.n419 585
R646 B.n421 B.n37 585
R647 B.n423 B.n422 585
R648 B.n424 B.n36 585
R649 B.n426 B.n425 585
R650 B.n427 B.n35 585
R651 B.n429 B.n428 585
R652 B.n430 B.n34 585
R653 B.n432 B.n431 585
R654 B.n434 B.n31 585
R655 B.n436 B.n435 585
R656 B.n437 B.n30 585
R657 B.n439 B.n438 585
R658 B.n440 B.n29 585
R659 B.n442 B.n441 585
R660 B.n443 B.n28 585
R661 B.n445 B.n444 585
R662 B.n446 B.n27 585
R663 B.n448 B.n447 585
R664 B.n449 B.n26 585
R665 B.n451 B.n450 585
R666 B.n452 B.n25 585
R667 B.n454 B.n453 585
R668 B.n455 B.n24 585
R669 B.n457 B.n456 585
R670 B.n458 B.n23 585
R671 B.n460 B.n459 585
R672 B.n461 B.n22 585
R673 B.n463 B.n462 585
R674 B.n464 B.n21 585
R675 B.n466 B.n465 585
R676 B.n467 B.n20 585
R677 B.n469 B.n468 585
R678 B.n470 B.n19 585
R679 B.n472 B.n471 585
R680 B.n473 B.n18 585
R681 B.n475 B.n474 585
R682 B.n476 B.n17 585
R683 B.n478 B.n477 585
R684 B.n479 B.n16 585
R685 B.n481 B.n480 585
R686 B.n482 B.n15 585
R687 B.n484 B.n483 585
R688 B.n367 B.n366 585
R689 B.n365 B.n58 585
R690 B.n364 B.n363 585
R691 B.n362 B.n59 585
R692 B.n361 B.n360 585
R693 B.n359 B.n60 585
R694 B.n358 B.n357 585
R695 B.n356 B.n61 585
R696 B.n355 B.n354 585
R697 B.n353 B.n62 585
R698 B.n352 B.n351 585
R699 B.n350 B.n63 585
R700 B.n349 B.n348 585
R701 B.n347 B.n64 585
R702 B.n346 B.n345 585
R703 B.n344 B.n65 585
R704 B.n343 B.n342 585
R705 B.n341 B.n66 585
R706 B.n340 B.n339 585
R707 B.n338 B.n67 585
R708 B.n337 B.n336 585
R709 B.n335 B.n68 585
R710 B.n334 B.n333 585
R711 B.n332 B.n69 585
R712 B.n331 B.n330 585
R713 B.n329 B.n70 585
R714 B.n328 B.n327 585
R715 B.n326 B.n71 585
R716 B.n325 B.n324 585
R717 B.n323 B.n72 585
R718 B.n322 B.n321 585
R719 B.n320 B.n73 585
R720 B.n319 B.n318 585
R721 B.n317 B.n74 585
R722 B.n316 B.n315 585
R723 B.n314 B.n75 585
R724 B.n313 B.n312 585
R725 B.n311 B.n76 585
R726 B.n310 B.n309 585
R727 B.n308 B.n77 585
R728 B.n307 B.n306 585
R729 B.n305 B.n78 585
R730 B.n304 B.n303 585
R731 B.n302 B.n79 585
R732 B.n301 B.n300 585
R733 B.n299 B.n80 585
R734 B.n298 B.n297 585
R735 B.n296 B.n81 585
R736 B.n295 B.n294 585
R737 B.n293 B.n82 585
R738 B.n292 B.n291 585
R739 B.n175 B.n174 585
R740 B.n176 B.n125 585
R741 B.n178 B.n177 585
R742 B.n179 B.n124 585
R743 B.n181 B.n180 585
R744 B.n182 B.n123 585
R745 B.n184 B.n183 585
R746 B.n185 B.n122 585
R747 B.n187 B.n186 585
R748 B.n188 B.n121 585
R749 B.n190 B.n189 585
R750 B.n191 B.n120 585
R751 B.n193 B.n192 585
R752 B.n194 B.n119 585
R753 B.n196 B.n195 585
R754 B.n197 B.n118 585
R755 B.n199 B.n198 585
R756 B.n200 B.n117 585
R757 B.n202 B.n201 585
R758 B.n203 B.n116 585
R759 B.n205 B.n204 585
R760 B.n206 B.n115 585
R761 B.n208 B.n207 585
R762 B.n209 B.n114 585
R763 B.n211 B.n210 585
R764 B.n212 B.n113 585
R765 B.n214 B.n213 585
R766 B.n215 B.n112 585
R767 B.n217 B.n216 585
R768 B.n218 B.n111 585
R769 B.n220 B.n219 585
R770 B.n221 B.n110 585
R771 B.n223 B.n222 585
R772 B.n224 B.n107 585
R773 B.n227 B.n226 585
R774 B.n228 B.n106 585
R775 B.n230 B.n229 585
R776 B.n231 B.n105 585
R777 B.n233 B.n232 585
R778 B.n234 B.n104 585
R779 B.n236 B.n235 585
R780 B.n237 B.n103 585
R781 B.n239 B.n238 585
R782 B.n241 B.n240 585
R783 B.n242 B.n99 585
R784 B.n244 B.n243 585
R785 B.n245 B.n98 585
R786 B.n247 B.n246 585
R787 B.n248 B.n97 585
R788 B.n250 B.n249 585
R789 B.n251 B.n96 585
R790 B.n253 B.n252 585
R791 B.n254 B.n95 585
R792 B.n256 B.n255 585
R793 B.n257 B.n94 585
R794 B.n259 B.n258 585
R795 B.n260 B.n93 585
R796 B.n262 B.n261 585
R797 B.n263 B.n92 585
R798 B.n265 B.n264 585
R799 B.n266 B.n91 585
R800 B.n268 B.n267 585
R801 B.n269 B.n90 585
R802 B.n271 B.n270 585
R803 B.n272 B.n89 585
R804 B.n274 B.n273 585
R805 B.n275 B.n88 585
R806 B.n277 B.n276 585
R807 B.n278 B.n87 585
R808 B.n280 B.n279 585
R809 B.n281 B.n86 585
R810 B.n283 B.n282 585
R811 B.n284 B.n85 585
R812 B.n286 B.n285 585
R813 B.n287 B.n84 585
R814 B.n289 B.n288 585
R815 B.n290 B.n83 585
R816 B.n173 B.n126 585
R817 B.n172 B.n171 585
R818 B.n170 B.n127 585
R819 B.n169 B.n168 585
R820 B.n167 B.n128 585
R821 B.n166 B.n165 585
R822 B.n164 B.n129 585
R823 B.n163 B.n162 585
R824 B.n161 B.n130 585
R825 B.n160 B.n159 585
R826 B.n158 B.n131 585
R827 B.n157 B.n156 585
R828 B.n155 B.n132 585
R829 B.n154 B.n153 585
R830 B.n152 B.n133 585
R831 B.n151 B.n150 585
R832 B.n149 B.n134 585
R833 B.n148 B.n147 585
R834 B.n146 B.n135 585
R835 B.n145 B.n144 585
R836 B.n143 B.n136 585
R837 B.n142 B.n141 585
R838 B.n140 B.n137 585
R839 B.n139 B.n138 585
R840 B.n2 B.n0 585
R841 B.n521 B.n1 585
R842 B.n520 B.n519 585
R843 B.n518 B.n3 585
R844 B.n517 B.n516 585
R845 B.n515 B.n4 585
R846 B.n514 B.n513 585
R847 B.n512 B.n5 585
R848 B.n511 B.n510 585
R849 B.n509 B.n6 585
R850 B.n508 B.n507 585
R851 B.n506 B.n7 585
R852 B.n505 B.n504 585
R853 B.n503 B.n8 585
R854 B.n502 B.n501 585
R855 B.n500 B.n9 585
R856 B.n499 B.n498 585
R857 B.n497 B.n10 585
R858 B.n496 B.n495 585
R859 B.n494 B.n11 585
R860 B.n493 B.n492 585
R861 B.n491 B.n12 585
R862 B.n490 B.n489 585
R863 B.n488 B.n13 585
R864 B.n487 B.n486 585
R865 B.n485 B.n14 585
R866 B.n523 B.n522 585
R867 B.n174 B.n173 502.111
R868 B.n485 B.n484 502.111
R869 B.n292 B.n83 502.111
R870 B.n366 B.n57 502.111
R871 B.n100 B.t2 382.615
R872 B.n38 B.t7 382.615
R873 B.n108 B.t11 382.615
R874 B.n32 B.t4 382.615
R875 B.n101 B.t1 326.567
R876 B.n39 B.t8 326.567
R877 B.n109 B.t10 326.567
R878 B.n33 B.t5 326.567
R879 B.n100 B.t0 295.349
R880 B.n108 B.t9 295.349
R881 B.n32 B.t3 295.349
R882 B.n38 B.t6 295.349
R883 B.n173 B.n172 163.367
R884 B.n172 B.n127 163.367
R885 B.n168 B.n127 163.367
R886 B.n168 B.n167 163.367
R887 B.n167 B.n166 163.367
R888 B.n166 B.n129 163.367
R889 B.n162 B.n129 163.367
R890 B.n162 B.n161 163.367
R891 B.n161 B.n160 163.367
R892 B.n160 B.n131 163.367
R893 B.n156 B.n131 163.367
R894 B.n156 B.n155 163.367
R895 B.n155 B.n154 163.367
R896 B.n154 B.n133 163.367
R897 B.n150 B.n133 163.367
R898 B.n150 B.n149 163.367
R899 B.n149 B.n148 163.367
R900 B.n148 B.n135 163.367
R901 B.n144 B.n135 163.367
R902 B.n144 B.n143 163.367
R903 B.n143 B.n142 163.367
R904 B.n142 B.n137 163.367
R905 B.n138 B.n137 163.367
R906 B.n138 B.n2 163.367
R907 B.n522 B.n2 163.367
R908 B.n522 B.n521 163.367
R909 B.n521 B.n520 163.367
R910 B.n520 B.n3 163.367
R911 B.n516 B.n3 163.367
R912 B.n516 B.n515 163.367
R913 B.n515 B.n514 163.367
R914 B.n514 B.n5 163.367
R915 B.n510 B.n5 163.367
R916 B.n510 B.n509 163.367
R917 B.n509 B.n508 163.367
R918 B.n508 B.n7 163.367
R919 B.n504 B.n7 163.367
R920 B.n504 B.n503 163.367
R921 B.n503 B.n502 163.367
R922 B.n502 B.n9 163.367
R923 B.n498 B.n9 163.367
R924 B.n498 B.n497 163.367
R925 B.n497 B.n496 163.367
R926 B.n496 B.n11 163.367
R927 B.n492 B.n11 163.367
R928 B.n492 B.n491 163.367
R929 B.n491 B.n490 163.367
R930 B.n490 B.n13 163.367
R931 B.n486 B.n13 163.367
R932 B.n486 B.n485 163.367
R933 B.n174 B.n125 163.367
R934 B.n178 B.n125 163.367
R935 B.n179 B.n178 163.367
R936 B.n180 B.n179 163.367
R937 B.n180 B.n123 163.367
R938 B.n184 B.n123 163.367
R939 B.n185 B.n184 163.367
R940 B.n186 B.n185 163.367
R941 B.n186 B.n121 163.367
R942 B.n190 B.n121 163.367
R943 B.n191 B.n190 163.367
R944 B.n192 B.n191 163.367
R945 B.n192 B.n119 163.367
R946 B.n196 B.n119 163.367
R947 B.n197 B.n196 163.367
R948 B.n198 B.n197 163.367
R949 B.n198 B.n117 163.367
R950 B.n202 B.n117 163.367
R951 B.n203 B.n202 163.367
R952 B.n204 B.n203 163.367
R953 B.n204 B.n115 163.367
R954 B.n208 B.n115 163.367
R955 B.n209 B.n208 163.367
R956 B.n210 B.n209 163.367
R957 B.n210 B.n113 163.367
R958 B.n214 B.n113 163.367
R959 B.n215 B.n214 163.367
R960 B.n216 B.n215 163.367
R961 B.n216 B.n111 163.367
R962 B.n220 B.n111 163.367
R963 B.n221 B.n220 163.367
R964 B.n222 B.n221 163.367
R965 B.n222 B.n107 163.367
R966 B.n227 B.n107 163.367
R967 B.n228 B.n227 163.367
R968 B.n229 B.n228 163.367
R969 B.n229 B.n105 163.367
R970 B.n233 B.n105 163.367
R971 B.n234 B.n233 163.367
R972 B.n235 B.n234 163.367
R973 B.n235 B.n103 163.367
R974 B.n239 B.n103 163.367
R975 B.n240 B.n239 163.367
R976 B.n240 B.n99 163.367
R977 B.n244 B.n99 163.367
R978 B.n245 B.n244 163.367
R979 B.n246 B.n245 163.367
R980 B.n246 B.n97 163.367
R981 B.n250 B.n97 163.367
R982 B.n251 B.n250 163.367
R983 B.n252 B.n251 163.367
R984 B.n252 B.n95 163.367
R985 B.n256 B.n95 163.367
R986 B.n257 B.n256 163.367
R987 B.n258 B.n257 163.367
R988 B.n258 B.n93 163.367
R989 B.n262 B.n93 163.367
R990 B.n263 B.n262 163.367
R991 B.n264 B.n263 163.367
R992 B.n264 B.n91 163.367
R993 B.n268 B.n91 163.367
R994 B.n269 B.n268 163.367
R995 B.n270 B.n269 163.367
R996 B.n270 B.n89 163.367
R997 B.n274 B.n89 163.367
R998 B.n275 B.n274 163.367
R999 B.n276 B.n275 163.367
R1000 B.n276 B.n87 163.367
R1001 B.n280 B.n87 163.367
R1002 B.n281 B.n280 163.367
R1003 B.n282 B.n281 163.367
R1004 B.n282 B.n85 163.367
R1005 B.n286 B.n85 163.367
R1006 B.n287 B.n286 163.367
R1007 B.n288 B.n287 163.367
R1008 B.n288 B.n83 163.367
R1009 B.n293 B.n292 163.367
R1010 B.n294 B.n293 163.367
R1011 B.n294 B.n81 163.367
R1012 B.n298 B.n81 163.367
R1013 B.n299 B.n298 163.367
R1014 B.n300 B.n299 163.367
R1015 B.n300 B.n79 163.367
R1016 B.n304 B.n79 163.367
R1017 B.n305 B.n304 163.367
R1018 B.n306 B.n305 163.367
R1019 B.n306 B.n77 163.367
R1020 B.n310 B.n77 163.367
R1021 B.n311 B.n310 163.367
R1022 B.n312 B.n311 163.367
R1023 B.n312 B.n75 163.367
R1024 B.n316 B.n75 163.367
R1025 B.n317 B.n316 163.367
R1026 B.n318 B.n317 163.367
R1027 B.n318 B.n73 163.367
R1028 B.n322 B.n73 163.367
R1029 B.n323 B.n322 163.367
R1030 B.n324 B.n323 163.367
R1031 B.n324 B.n71 163.367
R1032 B.n328 B.n71 163.367
R1033 B.n329 B.n328 163.367
R1034 B.n330 B.n329 163.367
R1035 B.n330 B.n69 163.367
R1036 B.n334 B.n69 163.367
R1037 B.n335 B.n334 163.367
R1038 B.n336 B.n335 163.367
R1039 B.n336 B.n67 163.367
R1040 B.n340 B.n67 163.367
R1041 B.n341 B.n340 163.367
R1042 B.n342 B.n341 163.367
R1043 B.n342 B.n65 163.367
R1044 B.n346 B.n65 163.367
R1045 B.n347 B.n346 163.367
R1046 B.n348 B.n347 163.367
R1047 B.n348 B.n63 163.367
R1048 B.n352 B.n63 163.367
R1049 B.n353 B.n352 163.367
R1050 B.n354 B.n353 163.367
R1051 B.n354 B.n61 163.367
R1052 B.n358 B.n61 163.367
R1053 B.n359 B.n358 163.367
R1054 B.n360 B.n359 163.367
R1055 B.n360 B.n59 163.367
R1056 B.n364 B.n59 163.367
R1057 B.n365 B.n364 163.367
R1058 B.n366 B.n365 163.367
R1059 B.n484 B.n15 163.367
R1060 B.n480 B.n15 163.367
R1061 B.n480 B.n479 163.367
R1062 B.n479 B.n478 163.367
R1063 B.n478 B.n17 163.367
R1064 B.n474 B.n17 163.367
R1065 B.n474 B.n473 163.367
R1066 B.n473 B.n472 163.367
R1067 B.n472 B.n19 163.367
R1068 B.n468 B.n19 163.367
R1069 B.n468 B.n467 163.367
R1070 B.n467 B.n466 163.367
R1071 B.n466 B.n21 163.367
R1072 B.n462 B.n21 163.367
R1073 B.n462 B.n461 163.367
R1074 B.n461 B.n460 163.367
R1075 B.n460 B.n23 163.367
R1076 B.n456 B.n23 163.367
R1077 B.n456 B.n455 163.367
R1078 B.n455 B.n454 163.367
R1079 B.n454 B.n25 163.367
R1080 B.n450 B.n25 163.367
R1081 B.n450 B.n449 163.367
R1082 B.n449 B.n448 163.367
R1083 B.n448 B.n27 163.367
R1084 B.n444 B.n27 163.367
R1085 B.n444 B.n443 163.367
R1086 B.n443 B.n442 163.367
R1087 B.n442 B.n29 163.367
R1088 B.n438 B.n29 163.367
R1089 B.n438 B.n437 163.367
R1090 B.n437 B.n436 163.367
R1091 B.n436 B.n31 163.367
R1092 B.n431 B.n31 163.367
R1093 B.n431 B.n430 163.367
R1094 B.n430 B.n429 163.367
R1095 B.n429 B.n35 163.367
R1096 B.n425 B.n35 163.367
R1097 B.n425 B.n424 163.367
R1098 B.n424 B.n423 163.367
R1099 B.n423 B.n37 163.367
R1100 B.n419 B.n37 163.367
R1101 B.n419 B.n418 163.367
R1102 B.n418 B.n41 163.367
R1103 B.n414 B.n41 163.367
R1104 B.n414 B.n413 163.367
R1105 B.n413 B.n412 163.367
R1106 B.n412 B.n43 163.367
R1107 B.n408 B.n43 163.367
R1108 B.n408 B.n407 163.367
R1109 B.n407 B.n406 163.367
R1110 B.n406 B.n45 163.367
R1111 B.n402 B.n45 163.367
R1112 B.n402 B.n401 163.367
R1113 B.n401 B.n400 163.367
R1114 B.n400 B.n47 163.367
R1115 B.n396 B.n47 163.367
R1116 B.n396 B.n395 163.367
R1117 B.n395 B.n394 163.367
R1118 B.n394 B.n49 163.367
R1119 B.n390 B.n49 163.367
R1120 B.n390 B.n389 163.367
R1121 B.n389 B.n388 163.367
R1122 B.n388 B.n51 163.367
R1123 B.n384 B.n51 163.367
R1124 B.n384 B.n383 163.367
R1125 B.n383 B.n382 163.367
R1126 B.n382 B.n53 163.367
R1127 B.n378 B.n53 163.367
R1128 B.n378 B.n377 163.367
R1129 B.n377 B.n376 163.367
R1130 B.n376 B.n55 163.367
R1131 B.n372 B.n55 163.367
R1132 B.n372 B.n371 163.367
R1133 B.n371 B.n370 163.367
R1134 B.n370 B.n57 163.367
R1135 B.n102 B.n101 59.5399
R1136 B.n225 B.n109 59.5399
R1137 B.n433 B.n33 59.5399
R1138 B.n40 B.n39 59.5399
R1139 B.n101 B.n100 56.049
R1140 B.n109 B.n108 56.049
R1141 B.n33 B.n32 56.049
R1142 B.n39 B.n38 56.049
R1143 B.n483 B.n14 32.6249
R1144 B.n368 B.n367 32.6249
R1145 B.n291 B.n290 32.6249
R1146 B.n175 B.n126 32.6249
R1147 B B.n523 18.0485
R1148 B.n483 B.n482 10.6151
R1149 B.n482 B.n481 10.6151
R1150 B.n481 B.n16 10.6151
R1151 B.n477 B.n16 10.6151
R1152 B.n477 B.n476 10.6151
R1153 B.n476 B.n475 10.6151
R1154 B.n475 B.n18 10.6151
R1155 B.n471 B.n18 10.6151
R1156 B.n471 B.n470 10.6151
R1157 B.n470 B.n469 10.6151
R1158 B.n469 B.n20 10.6151
R1159 B.n465 B.n20 10.6151
R1160 B.n465 B.n464 10.6151
R1161 B.n464 B.n463 10.6151
R1162 B.n463 B.n22 10.6151
R1163 B.n459 B.n22 10.6151
R1164 B.n459 B.n458 10.6151
R1165 B.n458 B.n457 10.6151
R1166 B.n457 B.n24 10.6151
R1167 B.n453 B.n24 10.6151
R1168 B.n453 B.n452 10.6151
R1169 B.n452 B.n451 10.6151
R1170 B.n451 B.n26 10.6151
R1171 B.n447 B.n26 10.6151
R1172 B.n447 B.n446 10.6151
R1173 B.n446 B.n445 10.6151
R1174 B.n445 B.n28 10.6151
R1175 B.n441 B.n28 10.6151
R1176 B.n441 B.n440 10.6151
R1177 B.n440 B.n439 10.6151
R1178 B.n439 B.n30 10.6151
R1179 B.n435 B.n30 10.6151
R1180 B.n435 B.n434 10.6151
R1181 B.n432 B.n34 10.6151
R1182 B.n428 B.n34 10.6151
R1183 B.n428 B.n427 10.6151
R1184 B.n427 B.n426 10.6151
R1185 B.n426 B.n36 10.6151
R1186 B.n422 B.n36 10.6151
R1187 B.n422 B.n421 10.6151
R1188 B.n421 B.n420 10.6151
R1189 B.n417 B.n416 10.6151
R1190 B.n416 B.n415 10.6151
R1191 B.n415 B.n42 10.6151
R1192 B.n411 B.n42 10.6151
R1193 B.n411 B.n410 10.6151
R1194 B.n410 B.n409 10.6151
R1195 B.n409 B.n44 10.6151
R1196 B.n405 B.n44 10.6151
R1197 B.n405 B.n404 10.6151
R1198 B.n404 B.n403 10.6151
R1199 B.n403 B.n46 10.6151
R1200 B.n399 B.n46 10.6151
R1201 B.n399 B.n398 10.6151
R1202 B.n398 B.n397 10.6151
R1203 B.n397 B.n48 10.6151
R1204 B.n393 B.n48 10.6151
R1205 B.n393 B.n392 10.6151
R1206 B.n392 B.n391 10.6151
R1207 B.n391 B.n50 10.6151
R1208 B.n387 B.n50 10.6151
R1209 B.n387 B.n386 10.6151
R1210 B.n386 B.n385 10.6151
R1211 B.n385 B.n52 10.6151
R1212 B.n381 B.n52 10.6151
R1213 B.n381 B.n380 10.6151
R1214 B.n380 B.n379 10.6151
R1215 B.n379 B.n54 10.6151
R1216 B.n375 B.n54 10.6151
R1217 B.n375 B.n374 10.6151
R1218 B.n374 B.n373 10.6151
R1219 B.n373 B.n56 10.6151
R1220 B.n369 B.n56 10.6151
R1221 B.n369 B.n368 10.6151
R1222 B.n291 B.n82 10.6151
R1223 B.n295 B.n82 10.6151
R1224 B.n296 B.n295 10.6151
R1225 B.n297 B.n296 10.6151
R1226 B.n297 B.n80 10.6151
R1227 B.n301 B.n80 10.6151
R1228 B.n302 B.n301 10.6151
R1229 B.n303 B.n302 10.6151
R1230 B.n303 B.n78 10.6151
R1231 B.n307 B.n78 10.6151
R1232 B.n308 B.n307 10.6151
R1233 B.n309 B.n308 10.6151
R1234 B.n309 B.n76 10.6151
R1235 B.n313 B.n76 10.6151
R1236 B.n314 B.n313 10.6151
R1237 B.n315 B.n314 10.6151
R1238 B.n315 B.n74 10.6151
R1239 B.n319 B.n74 10.6151
R1240 B.n320 B.n319 10.6151
R1241 B.n321 B.n320 10.6151
R1242 B.n321 B.n72 10.6151
R1243 B.n325 B.n72 10.6151
R1244 B.n326 B.n325 10.6151
R1245 B.n327 B.n326 10.6151
R1246 B.n327 B.n70 10.6151
R1247 B.n331 B.n70 10.6151
R1248 B.n332 B.n331 10.6151
R1249 B.n333 B.n332 10.6151
R1250 B.n333 B.n68 10.6151
R1251 B.n337 B.n68 10.6151
R1252 B.n338 B.n337 10.6151
R1253 B.n339 B.n338 10.6151
R1254 B.n339 B.n66 10.6151
R1255 B.n343 B.n66 10.6151
R1256 B.n344 B.n343 10.6151
R1257 B.n345 B.n344 10.6151
R1258 B.n345 B.n64 10.6151
R1259 B.n349 B.n64 10.6151
R1260 B.n350 B.n349 10.6151
R1261 B.n351 B.n350 10.6151
R1262 B.n351 B.n62 10.6151
R1263 B.n355 B.n62 10.6151
R1264 B.n356 B.n355 10.6151
R1265 B.n357 B.n356 10.6151
R1266 B.n357 B.n60 10.6151
R1267 B.n361 B.n60 10.6151
R1268 B.n362 B.n361 10.6151
R1269 B.n363 B.n362 10.6151
R1270 B.n363 B.n58 10.6151
R1271 B.n367 B.n58 10.6151
R1272 B.n176 B.n175 10.6151
R1273 B.n177 B.n176 10.6151
R1274 B.n177 B.n124 10.6151
R1275 B.n181 B.n124 10.6151
R1276 B.n182 B.n181 10.6151
R1277 B.n183 B.n182 10.6151
R1278 B.n183 B.n122 10.6151
R1279 B.n187 B.n122 10.6151
R1280 B.n188 B.n187 10.6151
R1281 B.n189 B.n188 10.6151
R1282 B.n189 B.n120 10.6151
R1283 B.n193 B.n120 10.6151
R1284 B.n194 B.n193 10.6151
R1285 B.n195 B.n194 10.6151
R1286 B.n195 B.n118 10.6151
R1287 B.n199 B.n118 10.6151
R1288 B.n200 B.n199 10.6151
R1289 B.n201 B.n200 10.6151
R1290 B.n201 B.n116 10.6151
R1291 B.n205 B.n116 10.6151
R1292 B.n206 B.n205 10.6151
R1293 B.n207 B.n206 10.6151
R1294 B.n207 B.n114 10.6151
R1295 B.n211 B.n114 10.6151
R1296 B.n212 B.n211 10.6151
R1297 B.n213 B.n212 10.6151
R1298 B.n213 B.n112 10.6151
R1299 B.n217 B.n112 10.6151
R1300 B.n218 B.n217 10.6151
R1301 B.n219 B.n218 10.6151
R1302 B.n219 B.n110 10.6151
R1303 B.n223 B.n110 10.6151
R1304 B.n224 B.n223 10.6151
R1305 B.n226 B.n106 10.6151
R1306 B.n230 B.n106 10.6151
R1307 B.n231 B.n230 10.6151
R1308 B.n232 B.n231 10.6151
R1309 B.n232 B.n104 10.6151
R1310 B.n236 B.n104 10.6151
R1311 B.n237 B.n236 10.6151
R1312 B.n238 B.n237 10.6151
R1313 B.n242 B.n241 10.6151
R1314 B.n243 B.n242 10.6151
R1315 B.n243 B.n98 10.6151
R1316 B.n247 B.n98 10.6151
R1317 B.n248 B.n247 10.6151
R1318 B.n249 B.n248 10.6151
R1319 B.n249 B.n96 10.6151
R1320 B.n253 B.n96 10.6151
R1321 B.n254 B.n253 10.6151
R1322 B.n255 B.n254 10.6151
R1323 B.n255 B.n94 10.6151
R1324 B.n259 B.n94 10.6151
R1325 B.n260 B.n259 10.6151
R1326 B.n261 B.n260 10.6151
R1327 B.n261 B.n92 10.6151
R1328 B.n265 B.n92 10.6151
R1329 B.n266 B.n265 10.6151
R1330 B.n267 B.n266 10.6151
R1331 B.n267 B.n90 10.6151
R1332 B.n271 B.n90 10.6151
R1333 B.n272 B.n271 10.6151
R1334 B.n273 B.n272 10.6151
R1335 B.n273 B.n88 10.6151
R1336 B.n277 B.n88 10.6151
R1337 B.n278 B.n277 10.6151
R1338 B.n279 B.n278 10.6151
R1339 B.n279 B.n86 10.6151
R1340 B.n283 B.n86 10.6151
R1341 B.n284 B.n283 10.6151
R1342 B.n285 B.n284 10.6151
R1343 B.n285 B.n84 10.6151
R1344 B.n289 B.n84 10.6151
R1345 B.n290 B.n289 10.6151
R1346 B.n171 B.n126 10.6151
R1347 B.n171 B.n170 10.6151
R1348 B.n170 B.n169 10.6151
R1349 B.n169 B.n128 10.6151
R1350 B.n165 B.n128 10.6151
R1351 B.n165 B.n164 10.6151
R1352 B.n164 B.n163 10.6151
R1353 B.n163 B.n130 10.6151
R1354 B.n159 B.n130 10.6151
R1355 B.n159 B.n158 10.6151
R1356 B.n158 B.n157 10.6151
R1357 B.n157 B.n132 10.6151
R1358 B.n153 B.n132 10.6151
R1359 B.n153 B.n152 10.6151
R1360 B.n152 B.n151 10.6151
R1361 B.n151 B.n134 10.6151
R1362 B.n147 B.n134 10.6151
R1363 B.n147 B.n146 10.6151
R1364 B.n146 B.n145 10.6151
R1365 B.n145 B.n136 10.6151
R1366 B.n141 B.n136 10.6151
R1367 B.n141 B.n140 10.6151
R1368 B.n140 B.n139 10.6151
R1369 B.n139 B.n0 10.6151
R1370 B.n519 B.n1 10.6151
R1371 B.n519 B.n518 10.6151
R1372 B.n518 B.n517 10.6151
R1373 B.n517 B.n4 10.6151
R1374 B.n513 B.n4 10.6151
R1375 B.n513 B.n512 10.6151
R1376 B.n512 B.n511 10.6151
R1377 B.n511 B.n6 10.6151
R1378 B.n507 B.n6 10.6151
R1379 B.n507 B.n506 10.6151
R1380 B.n506 B.n505 10.6151
R1381 B.n505 B.n8 10.6151
R1382 B.n501 B.n8 10.6151
R1383 B.n501 B.n500 10.6151
R1384 B.n500 B.n499 10.6151
R1385 B.n499 B.n10 10.6151
R1386 B.n495 B.n10 10.6151
R1387 B.n495 B.n494 10.6151
R1388 B.n494 B.n493 10.6151
R1389 B.n493 B.n12 10.6151
R1390 B.n489 B.n12 10.6151
R1391 B.n489 B.n488 10.6151
R1392 B.n488 B.n487 10.6151
R1393 B.n487 B.n14 10.6151
R1394 B.n433 B.n432 6.5566
R1395 B.n420 B.n40 6.5566
R1396 B.n226 B.n225 6.5566
R1397 B.n238 B.n102 6.5566
R1398 B.n434 B.n433 4.05904
R1399 B.n417 B.n40 4.05904
R1400 B.n225 B.n224 4.05904
R1401 B.n241 B.n102 4.05904
R1402 B.n523 B.n0 2.81026
R1403 B.n523 B.n1 2.81026
C0 w_n2126_n2824# B 8.00332f
C1 VDD1 VN 0.148438f
C2 VP VTAIL 1.99996f
C3 VDD1 w_n2126_n2824# 1.58759f
C4 VDD2 VTAIL 4.39175f
C5 VP B 1.45989f
C6 B VDD2 1.51502f
C7 VP VDD1 2.38165f
C8 VDD1 VDD2 0.669474f
C9 w_n2126_n2824# VN 2.8761f
C10 B VTAIL 3.03369f
C11 VP VN 4.92734f
C12 VN VDD2 2.20066f
C13 VDD1 VTAIL 4.34081f
C14 VP w_n2126_n2824# 3.14683f
C15 w_n2126_n2824# VDD2 1.61298f
C16 VDD1 B 1.48529f
C17 VP VDD2 0.331502f
C18 VN VTAIL 1.98571f
C19 w_n2126_n2824# VTAIL 2.3715f
C20 VN B 1.01497f
C21 VDD2 VSUBS 0.801683f
C22 VDD1 VSUBS 3.376427f
C23 VTAIL VSUBS 0.858134f
C24 VN VSUBS 6.45706f
C25 VP VSUBS 1.561969f
C26 B VSUBS 3.64996f
C27 w_n2126_n2824# VSUBS 74.265396f
C28 B.n0 VSUBS 0.004211f
C29 B.n1 VSUBS 0.004211f
C30 B.n2 VSUBS 0.00666f
C31 B.n3 VSUBS 0.00666f
C32 B.n4 VSUBS 0.00666f
C33 B.n5 VSUBS 0.00666f
C34 B.n6 VSUBS 0.00666f
C35 B.n7 VSUBS 0.00666f
C36 B.n8 VSUBS 0.00666f
C37 B.n9 VSUBS 0.00666f
C38 B.n10 VSUBS 0.00666f
C39 B.n11 VSUBS 0.00666f
C40 B.n12 VSUBS 0.00666f
C41 B.n13 VSUBS 0.00666f
C42 B.n14 VSUBS 0.015063f
C43 B.n15 VSUBS 0.00666f
C44 B.n16 VSUBS 0.00666f
C45 B.n17 VSUBS 0.00666f
C46 B.n18 VSUBS 0.00666f
C47 B.n19 VSUBS 0.00666f
C48 B.n20 VSUBS 0.00666f
C49 B.n21 VSUBS 0.00666f
C50 B.n22 VSUBS 0.00666f
C51 B.n23 VSUBS 0.00666f
C52 B.n24 VSUBS 0.00666f
C53 B.n25 VSUBS 0.00666f
C54 B.n26 VSUBS 0.00666f
C55 B.n27 VSUBS 0.00666f
C56 B.n28 VSUBS 0.00666f
C57 B.n29 VSUBS 0.00666f
C58 B.n30 VSUBS 0.00666f
C59 B.n31 VSUBS 0.00666f
C60 B.t5 VSUBS 0.14495f
C61 B.t4 VSUBS 0.173105f
C62 B.t3 VSUBS 1.0443f
C63 B.n32 VSUBS 0.282729f
C64 B.n33 VSUBS 0.201702f
C65 B.n34 VSUBS 0.00666f
C66 B.n35 VSUBS 0.00666f
C67 B.n36 VSUBS 0.00666f
C68 B.n37 VSUBS 0.00666f
C69 B.t8 VSUBS 0.144952f
C70 B.t7 VSUBS 0.173107f
C71 B.t6 VSUBS 1.0443f
C72 B.n38 VSUBS 0.282727f
C73 B.n39 VSUBS 0.2017f
C74 B.n40 VSUBS 0.01543f
C75 B.n41 VSUBS 0.00666f
C76 B.n42 VSUBS 0.00666f
C77 B.n43 VSUBS 0.00666f
C78 B.n44 VSUBS 0.00666f
C79 B.n45 VSUBS 0.00666f
C80 B.n46 VSUBS 0.00666f
C81 B.n47 VSUBS 0.00666f
C82 B.n48 VSUBS 0.00666f
C83 B.n49 VSUBS 0.00666f
C84 B.n50 VSUBS 0.00666f
C85 B.n51 VSUBS 0.00666f
C86 B.n52 VSUBS 0.00666f
C87 B.n53 VSUBS 0.00666f
C88 B.n54 VSUBS 0.00666f
C89 B.n55 VSUBS 0.00666f
C90 B.n56 VSUBS 0.00666f
C91 B.n57 VSUBS 0.016082f
C92 B.n58 VSUBS 0.00666f
C93 B.n59 VSUBS 0.00666f
C94 B.n60 VSUBS 0.00666f
C95 B.n61 VSUBS 0.00666f
C96 B.n62 VSUBS 0.00666f
C97 B.n63 VSUBS 0.00666f
C98 B.n64 VSUBS 0.00666f
C99 B.n65 VSUBS 0.00666f
C100 B.n66 VSUBS 0.00666f
C101 B.n67 VSUBS 0.00666f
C102 B.n68 VSUBS 0.00666f
C103 B.n69 VSUBS 0.00666f
C104 B.n70 VSUBS 0.00666f
C105 B.n71 VSUBS 0.00666f
C106 B.n72 VSUBS 0.00666f
C107 B.n73 VSUBS 0.00666f
C108 B.n74 VSUBS 0.00666f
C109 B.n75 VSUBS 0.00666f
C110 B.n76 VSUBS 0.00666f
C111 B.n77 VSUBS 0.00666f
C112 B.n78 VSUBS 0.00666f
C113 B.n79 VSUBS 0.00666f
C114 B.n80 VSUBS 0.00666f
C115 B.n81 VSUBS 0.00666f
C116 B.n82 VSUBS 0.00666f
C117 B.n83 VSUBS 0.016082f
C118 B.n84 VSUBS 0.00666f
C119 B.n85 VSUBS 0.00666f
C120 B.n86 VSUBS 0.00666f
C121 B.n87 VSUBS 0.00666f
C122 B.n88 VSUBS 0.00666f
C123 B.n89 VSUBS 0.00666f
C124 B.n90 VSUBS 0.00666f
C125 B.n91 VSUBS 0.00666f
C126 B.n92 VSUBS 0.00666f
C127 B.n93 VSUBS 0.00666f
C128 B.n94 VSUBS 0.00666f
C129 B.n95 VSUBS 0.00666f
C130 B.n96 VSUBS 0.00666f
C131 B.n97 VSUBS 0.00666f
C132 B.n98 VSUBS 0.00666f
C133 B.n99 VSUBS 0.00666f
C134 B.t1 VSUBS 0.144952f
C135 B.t2 VSUBS 0.173107f
C136 B.t0 VSUBS 1.0443f
C137 B.n100 VSUBS 0.282727f
C138 B.n101 VSUBS 0.2017f
C139 B.n102 VSUBS 0.01543f
C140 B.n103 VSUBS 0.00666f
C141 B.n104 VSUBS 0.00666f
C142 B.n105 VSUBS 0.00666f
C143 B.n106 VSUBS 0.00666f
C144 B.n107 VSUBS 0.00666f
C145 B.t10 VSUBS 0.14495f
C146 B.t11 VSUBS 0.173105f
C147 B.t9 VSUBS 1.0443f
C148 B.n108 VSUBS 0.282729f
C149 B.n109 VSUBS 0.201702f
C150 B.n110 VSUBS 0.00666f
C151 B.n111 VSUBS 0.00666f
C152 B.n112 VSUBS 0.00666f
C153 B.n113 VSUBS 0.00666f
C154 B.n114 VSUBS 0.00666f
C155 B.n115 VSUBS 0.00666f
C156 B.n116 VSUBS 0.00666f
C157 B.n117 VSUBS 0.00666f
C158 B.n118 VSUBS 0.00666f
C159 B.n119 VSUBS 0.00666f
C160 B.n120 VSUBS 0.00666f
C161 B.n121 VSUBS 0.00666f
C162 B.n122 VSUBS 0.00666f
C163 B.n123 VSUBS 0.00666f
C164 B.n124 VSUBS 0.00666f
C165 B.n125 VSUBS 0.00666f
C166 B.n126 VSUBS 0.015063f
C167 B.n127 VSUBS 0.00666f
C168 B.n128 VSUBS 0.00666f
C169 B.n129 VSUBS 0.00666f
C170 B.n130 VSUBS 0.00666f
C171 B.n131 VSUBS 0.00666f
C172 B.n132 VSUBS 0.00666f
C173 B.n133 VSUBS 0.00666f
C174 B.n134 VSUBS 0.00666f
C175 B.n135 VSUBS 0.00666f
C176 B.n136 VSUBS 0.00666f
C177 B.n137 VSUBS 0.00666f
C178 B.n138 VSUBS 0.00666f
C179 B.n139 VSUBS 0.00666f
C180 B.n140 VSUBS 0.00666f
C181 B.n141 VSUBS 0.00666f
C182 B.n142 VSUBS 0.00666f
C183 B.n143 VSUBS 0.00666f
C184 B.n144 VSUBS 0.00666f
C185 B.n145 VSUBS 0.00666f
C186 B.n146 VSUBS 0.00666f
C187 B.n147 VSUBS 0.00666f
C188 B.n148 VSUBS 0.00666f
C189 B.n149 VSUBS 0.00666f
C190 B.n150 VSUBS 0.00666f
C191 B.n151 VSUBS 0.00666f
C192 B.n152 VSUBS 0.00666f
C193 B.n153 VSUBS 0.00666f
C194 B.n154 VSUBS 0.00666f
C195 B.n155 VSUBS 0.00666f
C196 B.n156 VSUBS 0.00666f
C197 B.n157 VSUBS 0.00666f
C198 B.n158 VSUBS 0.00666f
C199 B.n159 VSUBS 0.00666f
C200 B.n160 VSUBS 0.00666f
C201 B.n161 VSUBS 0.00666f
C202 B.n162 VSUBS 0.00666f
C203 B.n163 VSUBS 0.00666f
C204 B.n164 VSUBS 0.00666f
C205 B.n165 VSUBS 0.00666f
C206 B.n166 VSUBS 0.00666f
C207 B.n167 VSUBS 0.00666f
C208 B.n168 VSUBS 0.00666f
C209 B.n169 VSUBS 0.00666f
C210 B.n170 VSUBS 0.00666f
C211 B.n171 VSUBS 0.00666f
C212 B.n172 VSUBS 0.00666f
C213 B.n173 VSUBS 0.015063f
C214 B.n174 VSUBS 0.016082f
C215 B.n175 VSUBS 0.016082f
C216 B.n176 VSUBS 0.00666f
C217 B.n177 VSUBS 0.00666f
C218 B.n178 VSUBS 0.00666f
C219 B.n179 VSUBS 0.00666f
C220 B.n180 VSUBS 0.00666f
C221 B.n181 VSUBS 0.00666f
C222 B.n182 VSUBS 0.00666f
C223 B.n183 VSUBS 0.00666f
C224 B.n184 VSUBS 0.00666f
C225 B.n185 VSUBS 0.00666f
C226 B.n186 VSUBS 0.00666f
C227 B.n187 VSUBS 0.00666f
C228 B.n188 VSUBS 0.00666f
C229 B.n189 VSUBS 0.00666f
C230 B.n190 VSUBS 0.00666f
C231 B.n191 VSUBS 0.00666f
C232 B.n192 VSUBS 0.00666f
C233 B.n193 VSUBS 0.00666f
C234 B.n194 VSUBS 0.00666f
C235 B.n195 VSUBS 0.00666f
C236 B.n196 VSUBS 0.00666f
C237 B.n197 VSUBS 0.00666f
C238 B.n198 VSUBS 0.00666f
C239 B.n199 VSUBS 0.00666f
C240 B.n200 VSUBS 0.00666f
C241 B.n201 VSUBS 0.00666f
C242 B.n202 VSUBS 0.00666f
C243 B.n203 VSUBS 0.00666f
C244 B.n204 VSUBS 0.00666f
C245 B.n205 VSUBS 0.00666f
C246 B.n206 VSUBS 0.00666f
C247 B.n207 VSUBS 0.00666f
C248 B.n208 VSUBS 0.00666f
C249 B.n209 VSUBS 0.00666f
C250 B.n210 VSUBS 0.00666f
C251 B.n211 VSUBS 0.00666f
C252 B.n212 VSUBS 0.00666f
C253 B.n213 VSUBS 0.00666f
C254 B.n214 VSUBS 0.00666f
C255 B.n215 VSUBS 0.00666f
C256 B.n216 VSUBS 0.00666f
C257 B.n217 VSUBS 0.00666f
C258 B.n218 VSUBS 0.00666f
C259 B.n219 VSUBS 0.00666f
C260 B.n220 VSUBS 0.00666f
C261 B.n221 VSUBS 0.00666f
C262 B.n222 VSUBS 0.00666f
C263 B.n223 VSUBS 0.00666f
C264 B.n224 VSUBS 0.004603f
C265 B.n225 VSUBS 0.01543f
C266 B.n226 VSUBS 0.005387f
C267 B.n227 VSUBS 0.00666f
C268 B.n228 VSUBS 0.00666f
C269 B.n229 VSUBS 0.00666f
C270 B.n230 VSUBS 0.00666f
C271 B.n231 VSUBS 0.00666f
C272 B.n232 VSUBS 0.00666f
C273 B.n233 VSUBS 0.00666f
C274 B.n234 VSUBS 0.00666f
C275 B.n235 VSUBS 0.00666f
C276 B.n236 VSUBS 0.00666f
C277 B.n237 VSUBS 0.00666f
C278 B.n238 VSUBS 0.005387f
C279 B.n239 VSUBS 0.00666f
C280 B.n240 VSUBS 0.00666f
C281 B.n241 VSUBS 0.004603f
C282 B.n242 VSUBS 0.00666f
C283 B.n243 VSUBS 0.00666f
C284 B.n244 VSUBS 0.00666f
C285 B.n245 VSUBS 0.00666f
C286 B.n246 VSUBS 0.00666f
C287 B.n247 VSUBS 0.00666f
C288 B.n248 VSUBS 0.00666f
C289 B.n249 VSUBS 0.00666f
C290 B.n250 VSUBS 0.00666f
C291 B.n251 VSUBS 0.00666f
C292 B.n252 VSUBS 0.00666f
C293 B.n253 VSUBS 0.00666f
C294 B.n254 VSUBS 0.00666f
C295 B.n255 VSUBS 0.00666f
C296 B.n256 VSUBS 0.00666f
C297 B.n257 VSUBS 0.00666f
C298 B.n258 VSUBS 0.00666f
C299 B.n259 VSUBS 0.00666f
C300 B.n260 VSUBS 0.00666f
C301 B.n261 VSUBS 0.00666f
C302 B.n262 VSUBS 0.00666f
C303 B.n263 VSUBS 0.00666f
C304 B.n264 VSUBS 0.00666f
C305 B.n265 VSUBS 0.00666f
C306 B.n266 VSUBS 0.00666f
C307 B.n267 VSUBS 0.00666f
C308 B.n268 VSUBS 0.00666f
C309 B.n269 VSUBS 0.00666f
C310 B.n270 VSUBS 0.00666f
C311 B.n271 VSUBS 0.00666f
C312 B.n272 VSUBS 0.00666f
C313 B.n273 VSUBS 0.00666f
C314 B.n274 VSUBS 0.00666f
C315 B.n275 VSUBS 0.00666f
C316 B.n276 VSUBS 0.00666f
C317 B.n277 VSUBS 0.00666f
C318 B.n278 VSUBS 0.00666f
C319 B.n279 VSUBS 0.00666f
C320 B.n280 VSUBS 0.00666f
C321 B.n281 VSUBS 0.00666f
C322 B.n282 VSUBS 0.00666f
C323 B.n283 VSUBS 0.00666f
C324 B.n284 VSUBS 0.00666f
C325 B.n285 VSUBS 0.00666f
C326 B.n286 VSUBS 0.00666f
C327 B.n287 VSUBS 0.00666f
C328 B.n288 VSUBS 0.00666f
C329 B.n289 VSUBS 0.00666f
C330 B.n290 VSUBS 0.016082f
C331 B.n291 VSUBS 0.015063f
C332 B.n292 VSUBS 0.015063f
C333 B.n293 VSUBS 0.00666f
C334 B.n294 VSUBS 0.00666f
C335 B.n295 VSUBS 0.00666f
C336 B.n296 VSUBS 0.00666f
C337 B.n297 VSUBS 0.00666f
C338 B.n298 VSUBS 0.00666f
C339 B.n299 VSUBS 0.00666f
C340 B.n300 VSUBS 0.00666f
C341 B.n301 VSUBS 0.00666f
C342 B.n302 VSUBS 0.00666f
C343 B.n303 VSUBS 0.00666f
C344 B.n304 VSUBS 0.00666f
C345 B.n305 VSUBS 0.00666f
C346 B.n306 VSUBS 0.00666f
C347 B.n307 VSUBS 0.00666f
C348 B.n308 VSUBS 0.00666f
C349 B.n309 VSUBS 0.00666f
C350 B.n310 VSUBS 0.00666f
C351 B.n311 VSUBS 0.00666f
C352 B.n312 VSUBS 0.00666f
C353 B.n313 VSUBS 0.00666f
C354 B.n314 VSUBS 0.00666f
C355 B.n315 VSUBS 0.00666f
C356 B.n316 VSUBS 0.00666f
C357 B.n317 VSUBS 0.00666f
C358 B.n318 VSUBS 0.00666f
C359 B.n319 VSUBS 0.00666f
C360 B.n320 VSUBS 0.00666f
C361 B.n321 VSUBS 0.00666f
C362 B.n322 VSUBS 0.00666f
C363 B.n323 VSUBS 0.00666f
C364 B.n324 VSUBS 0.00666f
C365 B.n325 VSUBS 0.00666f
C366 B.n326 VSUBS 0.00666f
C367 B.n327 VSUBS 0.00666f
C368 B.n328 VSUBS 0.00666f
C369 B.n329 VSUBS 0.00666f
C370 B.n330 VSUBS 0.00666f
C371 B.n331 VSUBS 0.00666f
C372 B.n332 VSUBS 0.00666f
C373 B.n333 VSUBS 0.00666f
C374 B.n334 VSUBS 0.00666f
C375 B.n335 VSUBS 0.00666f
C376 B.n336 VSUBS 0.00666f
C377 B.n337 VSUBS 0.00666f
C378 B.n338 VSUBS 0.00666f
C379 B.n339 VSUBS 0.00666f
C380 B.n340 VSUBS 0.00666f
C381 B.n341 VSUBS 0.00666f
C382 B.n342 VSUBS 0.00666f
C383 B.n343 VSUBS 0.00666f
C384 B.n344 VSUBS 0.00666f
C385 B.n345 VSUBS 0.00666f
C386 B.n346 VSUBS 0.00666f
C387 B.n347 VSUBS 0.00666f
C388 B.n348 VSUBS 0.00666f
C389 B.n349 VSUBS 0.00666f
C390 B.n350 VSUBS 0.00666f
C391 B.n351 VSUBS 0.00666f
C392 B.n352 VSUBS 0.00666f
C393 B.n353 VSUBS 0.00666f
C394 B.n354 VSUBS 0.00666f
C395 B.n355 VSUBS 0.00666f
C396 B.n356 VSUBS 0.00666f
C397 B.n357 VSUBS 0.00666f
C398 B.n358 VSUBS 0.00666f
C399 B.n359 VSUBS 0.00666f
C400 B.n360 VSUBS 0.00666f
C401 B.n361 VSUBS 0.00666f
C402 B.n362 VSUBS 0.00666f
C403 B.n363 VSUBS 0.00666f
C404 B.n364 VSUBS 0.00666f
C405 B.n365 VSUBS 0.00666f
C406 B.n366 VSUBS 0.015063f
C407 B.n367 VSUBS 0.015851f
C408 B.n368 VSUBS 0.015294f
C409 B.n369 VSUBS 0.00666f
C410 B.n370 VSUBS 0.00666f
C411 B.n371 VSUBS 0.00666f
C412 B.n372 VSUBS 0.00666f
C413 B.n373 VSUBS 0.00666f
C414 B.n374 VSUBS 0.00666f
C415 B.n375 VSUBS 0.00666f
C416 B.n376 VSUBS 0.00666f
C417 B.n377 VSUBS 0.00666f
C418 B.n378 VSUBS 0.00666f
C419 B.n379 VSUBS 0.00666f
C420 B.n380 VSUBS 0.00666f
C421 B.n381 VSUBS 0.00666f
C422 B.n382 VSUBS 0.00666f
C423 B.n383 VSUBS 0.00666f
C424 B.n384 VSUBS 0.00666f
C425 B.n385 VSUBS 0.00666f
C426 B.n386 VSUBS 0.00666f
C427 B.n387 VSUBS 0.00666f
C428 B.n388 VSUBS 0.00666f
C429 B.n389 VSUBS 0.00666f
C430 B.n390 VSUBS 0.00666f
C431 B.n391 VSUBS 0.00666f
C432 B.n392 VSUBS 0.00666f
C433 B.n393 VSUBS 0.00666f
C434 B.n394 VSUBS 0.00666f
C435 B.n395 VSUBS 0.00666f
C436 B.n396 VSUBS 0.00666f
C437 B.n397 VSUBS 0.00666f
C438 B.n398 VSUBS 0.00666f
C439 B.n399 VSUBS 0.00666f
C440 B.n400 VSUBS 0.00666f
C441 B.n401 VSUBS 0.00666f
C442 B.n402 VSUBS 0.00666f
C443 B.n403 VSUBS 0.00666f
C444 B.n404 VSUBS 0.00666f
C445 B.n405 VSUBS 0.00666f
C446 B.n406 VSUBS 0.00666f
C447 B.n407 VSUBS 0.00666f
C448 B.n408 VSUBS 0.00666f
C449 B.n409 VSUBS 0.00666f
C450 B.n410 VSUBS 0.00666f
C451 B.n411 VSUBS 0.00666f
C452 B.n412 VSUBS 0.00666f
C453 B.n413 VSUBS 0.00666f
C454 B.n414 VSUBS 0.00666f
C455 B.n415 VSUBS 0.00666f
C456 B.n416 VSUBS 0.00666f
C457 B.n417 VSUBS 0.004603f
C458 B.n418 VSUBS 0.00666f
C459 B.n419 VSUBS 0.00666f
C460 B.n420 VSUBS 0.005387f
C461 B.n421 VSUBS 0.00666f
C462 B.n422 VSUBS 0.00666f
C463 B.n423 VSUBS 0.00666f
C464 B.n424 VSUBS 0.00666f
C465 B.n425 VSUBS 0.00666f
C466 B.n426 VSUBS 0.00666f
C467 B.n427 VSUBS 0.00666f
C468 B.n428 VSUBS 0.00666f
C469 B.n429 VSUBS 0.00666f
C470 B.n430 VSUBS 0.00666f
C471 B.n431 VSUBS 0.00666f
C472 B.n432 VSUBS 0.005387f
C473 B.n433 VSUBS 0.01543f
C474 B.n434 VSUBS 0.004603f
C475 B.n435 VSUBS 0.00666f
C476 B.n436 VSUBS 0.00666f
C477 B.n437 VSUBS 0.00666f
C478 B.n438 VSUBS 0.00666f
C479 B.n439 VSUBS 0.00666f
C480 B.n440 VSUBS 0.00666f
C481 B.n441 VSUBS 0.00666f
C482 B.n442 VSUBS 0.00666f
C483 B.n443 VSUBS 0.00666f
C484 B.n444 VSUBS 0.00666f
C485 B.n445 VSUBS 0.00666f
C486 B.n446 VSUBS 0.00666f
C487 B.n447 VSUBS 0.00666f
C488 B.n448 VSUBS 0.00666f
C489 B.n449 VSUBS 0.00666f
C490 B.n450 VSUBS 0.00666f
C491 B.n451 VSUBS 0.00666f
C492 B.n452 VSUBS 0.00666f
C493 B.n453 VSUBS 0.00666f
C494 B.n454 VSUBS 0.00666f
C495 B.n455 VSUBS 0.00666f
C496 B.n456 VSUBS 0.00666f
C497 B.n457 VSUBS 0.00666f
C498 B.n458 VSUBS 0.00666f
C499 B.n459 VSUBS 0.00666f
C500 B.n460 VSUBS 0.00666f
C501 B.n461 VSUBS 0.00666f
C502 B.n462 VSUBS 0.00666f
C503 B.n463 VSUBS 0.00666f
C504 B.n464 VSUBS 0.00666f
C505 B.n465 VSUBS 0.00666f
C506 B.n466 VSUBS 0.00666f
C507 B.n467 VSUBS 0.00666f
C508 B.n468 VSUBS 0.00666f
C509 B.n469 VSUBS 0.00666f
C510 B.n470 VSUBS 0.00666f
C511 B.n471 VSUBS 0.00666f
C512 B.n472 VSUBS 0.00666f
C513 B.n473 VSUBS 0.00666f
C514 B.n474 VSUBS 0.00666f
C515 B.n475 VSUBS 0.00666f
C516 B.n476 VSUBS 0.00666f
C517 B.n477 VSUBS 0.00666f
C518 B.n478 VSUBS 0.00666f
C519 B.n479 VSUBS 0.00666f
C520 B.n480 VSUBS 0.00666f
C521 B.n481 VSUBS 0.00666f
C522 B.n482 VSUBS 0.00666f
C523 B.n483 VSUBS 0.016082f
C524 B.n484 VSUBS 0.016082f
C525 B.n485 VSUBS 0.015063f
C526 B.n486 VSUBS 0.00666f
C527 B.n487 VSUBS 0.00666f
C528 B.n488 VSUBS 0.00666f
C529 B.n489 VSUBS 0.00666f
C530 B.n490 VSUBS 0.00666f
C531 B.n491 VSUBS 0.00666f
C532 B.n492 VSUBS 0.00666f
C533 B.n493 VSUBS 0.00666f
C534 B.n494 VSUBS 0.00666f
C535 B.n495 VSUBS 0.00666f
C536 B.n496 VSUBS 0.00666f
C537 B.n497 VSUBS 0.00666f
C538 B.n498 VSUBS 0.00666f
C539 B.n499 VSUBS 0.00666f
C540 B.n500 VSUBS 0.00666f
C541 B.n501 VSUBS 0.00666f
C542 B.n502 VSUBS 0.00666f
C543 B.n503 VSUBS 0.00666f
C544 B.n504 VSUBS 0.00666f
C545 B.n505 VSUBS 0.00666f
C546 B.n506 VSUBS 0.00666f
C547 B.n507 VSUBS 0.00666f
C548 B.n508 VSUBS 0.00666f
C549 B.n509 VSUBS 0.00666f
C550 B.n510 VSUBS 0.00666f
C551 B.n511 VSUBS 0.00666f
C552 B.n512 VSUBS 0.00666f
C553 B.n513 VSUBS 0.00666f
C554 B.n514 VSUBS 0.00666f
C555 B.n515 VSUBS 0.00666f
C556 B.n516 VSUBS 0.00666f
C557 B.n517 VSUBS 0.00666f
C558 B.n518 VSUBS 0.00666f
C559 B.n519 VSUBS 0.00666f
C560 B.n520 VSUBS 0.00666f
C561 B.n521 VSUBS 0.00666f
C562 B.n522 VSUBS 0.00666f
C563 B.n523 VSUBS 0.01508f
C564 VDD1.n0 VSUBS 0.021498f
C565 VDD1.n1 VSUBS 0.020597f
C566 VDD1.n2 VSUBS 0.011068f
C567 VDD1.n3 VSUBS 0.026161f
C568 VDD1.n4 VSUBS 0.011394f
C569 VDD1.n5 VSUBS 0.020597f
C570 VDD1.n6 VSUBS 0.011394f
C571 VDD1.n7 VSUBS 0.011068f
C572 VDD1.n8 VSUBS 0.026161f
C573 VDD1.n9 VSUBS 0.026161f
C574 VDD1.n10 VSUBS 0.011719f
C575 VDD1.n11 VSUBS 0.020597f
C576 VDD1.n12 VSUBS 0.011068f
C577 VDD1.n13 VSUBS 0.026161f
C578 VDD1.n14 VSUBS 0.011719f
C579 VDD1.n15 VSUBS 0.766478f
C580 VDD1.n16 VSUBS 0.011068f
C581 VDD1.t0 VSUBS 0.056211f
C582 VDD1.n17 VSUBS 0.136906f
C583 VDD1.n18 VSUBS 0.019679f
C584 VDD1.n19 VSUBS 0.019621f
C585 VDD1.n20 VSUBS 0.026161f
C586 VDD1.n21 VSUBS 0.011719f
C587 VDD1.n22 VSUBS 0.011068f
C588 VDD1.n23 VSUBS 0.020597f
C589 VDD1.n24 VSUBS 0.020597f
C590 VDD1.n25 VSUBS 0.011068f
C591 VDD1.n26 VSUBS 0.011719f
C592 VDD1.n27 VSUBS 0.026161f
C593 VDD1.n28 VSUBS 0.026161f
C594 VDD1.n29 VSUBS 0.011719f
C595 VDD1.n30 VSUBS 0.011068f
C596 VDD1.n31 VSUBS 0.020597f
C597 VDD1.n32 VSUBS 0.020597f
C598 VDD1.n33 VSUBS 0.011068f
C599 VDD1.n34 VSUBS 0.011719f
C600 VDD1.n35 VSUBS 0.026161f
C601 VDD1.n36 VSUBS 0.026161f
C602 VDD1.n37 VSUBS 0.011719f
C603 VDD1.n38 VSUBS 0.011068f
C604 VDD1.n39 VSUBS 0.020597f
C605 VDD1.n40 VSUBS 0.020597f
C606 VDD1.n41 VSUBS 0.011068f
C607 VDD1.n42 VSUBS 0.011719f
C608 VDD1.n43 VSUBS 0.026161f
C609 VDD1.n44 VSUBS 0.05947f
C610 VDD1.n45 VSUBS 0.011719f
C611 VDD1.n46 VSUBS 0.011068f
C612 VDD1.n47 VSUBS 0.048735f
C613 VDD1.n48 VSUBS 0.04514f
C614 VDD1.n49 VSUBS 0.021498f
C615 VDD1.n50 VSUBS 0.020597f
C616 VDD1.n51 VSUBS 0.011068f
C617 VDD1.n52 VSUBS 0.026161f
C618 VDD1.n53 VSUBS 0.011394f
C619 VDD1.n54 VSUBS 0.020597f
C620 VDD1.n55 VSUBS 0.011719f
C621 VDD1.n56 VSUBS 0.026161f
C622 VDD1.n57 VSUBS 0.011719f
C623 VDD1.n58 VSUBS 0.020597f
C624 VDD1.n59 VSUBS 0.011068f
C625 VDD1.n60 VSUBS 0.026161f
C626 VDD1.n61 VSUBS 0.011719f
C627 VDD1.n62 VSUBS 0.766478f
C628 VDD1.n63 VSUBS 0.011068f
C629 VDD1.t1 VSUBS 0.056211f
C630 VDD1.n64 VSUBS 0.136906f
C631 VDD1.n65 VSUBS 0.019679f
C632 VDD1.n66 VSUBS 0.019621f
C633 VDD1.n67 VSUBS 0.026161f
C634 VDD1.n68 VSUBS 0.011719f
C635 VDD1.n69 VSUBS 0.011068f
C636 VDD1.n70 VSUBS 0.020597f
C637 VDD1.n71 VSUBS 0.020597f
C638 VDD1.n72 VSUBS 0.011068f
C639 VDD1.n73 VSUBS 0.011719f
C640 VDD1.n74 VSUBS 0.026161f
C641 VDD1.n75 VSUBS 0.026161f
C642 VDD1.n76 VSUBS 0.011719f
C643 VDD1.n77 VSUBS 0.011068f
C644 VDD1.n78 VSUBS 0.020597f
C645 VDD1.n79 VSUBS 0.020597f
C646 VDD1.n80 VSUBS 0.011068f
C647 VDD1.n81 VSUBS 0.011068f
C648 VDD1.n82 VSUBS 0.011719f
C649 VDD1.n83 VSUBS 0.026161f
C650 VDD1.n84 VSUBS 0.026161f
C651 VDD1.n85 VSUBS 0.026161f
C652 VDD1.n86 VSUBS 0.011394f
C653 VDD1.n87 VSUBS 0.011068f
C654 VDD1.n88 VSUBS 0.020597f
C655 VDD1.n89 VSUBS 0.020597f
C656 VDD1.n90 VSUBS 0.011068f
C657 VDD1.n91 VSUBS 0.011719f
C658 VDD1.n92 VSUBS 0.026161f
C659 VDD1.n93 VSUBS 0.05947f
C660 VDD1.n94 VSUBS 0.011719f
C661 VDD1.n95 VSUBS 0.011068f
C662 VDD1.n96 VSUBS 0.048735f
C663 VDD1.n97 VSUBS 0.558074f
C664 VP.t1 VSUBS 3.34244f
C665 VP.t0 VSUBS 2.76941f
C666 VP.n0 VSUBS 4.20095f
C667 VDD2.n0 VSUBS 0.02142f
C668 VDD2.n1 VSUBS 0.020523f
C669 VDD2.n2 VSUBS 0.011028f
C670 VDD2.n3 VSUBS 0.026066f
C671 VDD2.n4 VSUBS 0.011352f
C672 VDD2.n5 VSUBS 0.020523f
C673 VDD2.n6 VSUBS 0.011677f
C674 VDD2.n7 VSUBS 0.026066f
C675 VDD2.n8 VSUBS 0.011677f
C676 VDD2.n9 VSUBS 0.020523f
C677 VDD2.n10 VSUBS 0.011028f
C678 VDD2.n11 VSUBS 0.026066f
C679 VDD2.n12 VSUBS 0.011677f
C680 VDD2.n13 VSUBS 0.763709f
C681 VDD2.n14 VSUBS 0.011028f
C682 VDD2.t1 VSUBS 0.056008f
C683 VDD2.n15 VSUBS 0.136412f
C684 VDD2.n16 VSUBS 0.019608f
C685 VDD2.n17 VSUBS 0.01955f
C686 VDD2.n18 VSUBS 0.026066f
C687 VDD2.n19 VSUBS 0.011677f
C688 VDD2.n20 VSUBS 0.011028f
C689 VDD2.n21 VSUBS 0.020523f
C690 VDD2.n22 VSUBS 0.020523f
C691 VDD2.n23 VSUBS 0.011028f
C692 VDD2.n24 VSUBS 0.011677f
C693 VDD2.n25 VSUBS 0.026066f
C694 VDD2.n26 VSUBS 0.026066f
C695 VDD2.n27 VSUBS 0.011677f
C696 VDD2.n28 VSUBS 0.011028f
C697 VDD2.n29 VSUBS 0.020523f
C698 VDD2.n30 VSUBS 0.020523f
C699 VDD2.n31 VSUBS 0.011028f
C700 VDD2.n32 VSUBS 0.011028f
C701 VDD2.n33 VSUBS 0.011677f
C702 VDD2.n34 VSUBS 0.026066f
C703 VDD2.n35 VSUBS 0.026066f
C704 VDD2.n36 VSUBS 0.026066f
C705 VDD2.n37 VSUBS 0.011352f
C706 VDD2.n38 VSUBS 0.011028f
C707 VDD2.n39 VSUBS 0.020523f
C708 VDD2.n40 VSUBS 0.020523f
C709 VDD2.n41 VSUBS 0.011028f
C710 VDD2.n42 VSUBS 0.011677f
C711 VDD2.n43 VSUBS 0.026066f
C712 VDD2.n44 VSUBS 0.059255f
C713 VDD2.n45 VSUBS 0.011677f
C714 VDD2.n46 VSUBS 0.011028f
C715 VDD2.n47 VSUBS 0.048559f
C716 VDD2.n48 VSUBS 0.51832f
C717 VDD2.n49 VSUBS 0.02142f
C718 VDD2.n50 VSUBS 0.020523f
C719 VDD2.n51 VSUBS 0.011028f
C720 VDD2.n52 VSUBS 0.026066f
C721 VDD2.n53 VSUBS 0.011352f
C722 VDD2.n54 VSUBS 0.020523f
C723 VDD2.n55 VSUBS 0.011352f
C724 VDD2.n56 VSUBS 0.011028f
C725 VDD2.n57 VSUBS 0.026066f
C726 VDD2.n58 VSUBS 0.026066f
C727 VDD2.n59 VSUBS 0.011677f
C728 VDD2.n60 VSUBS 0.020523f
C729 VDD2.n61 VSUBS 0.011028f
C730 VDD2.n62 VSUBS 0.026066f
C731 VDD2.n63 VSUBS 0.011677f
C732 VDD2.n64 VSUBS 0.763709f
C733 VDD2.n65 VSUBS 0.011028f
C734 VDD2.t0 VSUBS 0.056008f
C735 VDD2.n66 VSUBS 0.136412f
C736 VDD2.n67 VSUBS 0.019608f
C737 VDD2.n68 VSUBS 0.01955f
C738 VDD2.n69 VSUBS 0.026066f
C739 VDD2.n70 VSUBS 0.011677f
C740 VDD2.n71 VSUBS 0.011028f
C741 VDD2.n72 VSUBS 0.020523f
C742 VDD2.n73 VSUBS 0.020523f
C743 VDD2.n74 VSUBS 0.011028f
C744 VDD2.n75 VSUBS 0.011677f
C745 VDD2.n76 VSUBS 0.026066f
C746 VDD2.n77 VSUBS 0.026066f
C747 VDD2.n78 VSUBS 0.011677f
C748 VDD2.n79 VSUBS 0.011028f
C749 VDD2.n80 VSUBS 0.020523f
C750 VDD2.n81 VSUBS 0.020523f
C751 VDD2.n82 VSUBS 0.011028f
C752 VDD2.n83 VSUBS 0.011677f
C753 VDD2.n84 VSUBS 0.026066f
C754 VDD2.n85 VSUBS 0.026066f
C755 VDD2.n86 VSUBS 0.011677f
C756 VDD2.n87 VSUBS 0.011028f
C757 VDD2.n88 VSUBS 0.020523f
C758 VDD2.n89 VSUBS 0.020523f
C759 VDD2.n90 VSUBS 0.011028f
C760 VDD2.n91 VSUBS 0.011677f
C761 VDD2.n92 VSUBS 0.026066f
C762 VDD2.n93 VSUBS 0.059255f
C763 VDD2.n94 VSUBS 0.011677f
C764 VDD2.n95 VSUBS 0.011028f
C765 VDD2.n96 VSUBS 0.048559f
C766 VDD2.n97 VSUBS 0.043824f
C767 VDD2.n98 VSUBS 2.27188f
C768 VTAIL.n0 VSUBS 0.024877f
C769 VTAIL.n1 VSUBS 0.023835f
C770 VTAIL.n2 VSUBS 0.012808f
C771 VTAIL.n3 VSUBS 0.030273f
C772 VTAIL.n4 VSUBS 0.013184f
C773 VTAIL.n5 VSUBS 0.023835f
C774 VTAIL.n6 VSUBS 0.013561f
C775 VTAIL.n7 VSUBS 0.030273f
C776 VTAIL.n8 VSUBS 0.013561f
C777 VTAIL.n9 VSUBS 0.023835f
C778 VTAIL.n10 VSUBS 0.012808f
C779 VTAIL.n11 VSUBS 0.030273f
C780 VTAIL.n12 VSUBS 0.013561f
C781 VTAIL.n13 VSUBS 0.88695f
C782 VTAIL.n14 VSUBS 0.012808f
C783 VTAIL.t1 VSUBS 0.065047f
C784 VTAIL.n15 VSUBS 0.158425f
C785 VTAIL.n16 VSUBS 0.022773f
C786 VTAIL.n17 VSUBS 0.022705f
C787 VTAIL.n18 VSUBS 0.030273f
C788 VTAIL.n19 VSUBS 0.013561f
C789 VTAIL.n20 VSUBS 0.012808f
C790 VTAIL.n21 VSUBS 0.023835f
C791 VTAIL.n22 VSUBS 0.023835f
C792 VTAIL.n23 VSUBS 0.012808f
C793 VTAIL.n24 VSUBS 0.013561f
C794 VTAIL.n25 VSUBS 0.030273f
C795 VTAIL.n26 VSUBS 0.030273f
C796 VTAIL.n27 VSUBS 0.013561f
C797 VTAIL.n28 VSUBS 0.012808f
C798 VTAIL.n29 VSUBS 0.023835f
C799 VTAIL.n30 VSUBS 0.023835f
C800 VTAIL.n31 VSUBS 0.012808f
C801 VTAIL.n32 VSUBS 0.012808f
C802 VTAIL.n33 VSUBS 0.013561f
C803 VTAIL.n34 VSUBS 0.030273f
C804 VTAIL.n35 VSUBS 0.030273f
C805 VTAIL.n36 VSUBS 0.030273f
C806 VTAIL.n37 VSUBS 0.013184f
C807 VTAIL.n38 VSUBS 0.012808f
C808 VTAIL.n39 VSUBS 0.023835f
C809 VTAIL.n40 VSUBS 0.023835f
C810 VTAIL.n41 VSUBS 0.012808f
C811 VTAIL.n42 VSUBS 0.013561f
C812 VTAIL.n43 VSUBS 0.030273f
C813 VTAIL.n44 VSUBS 0.068818f
C814 VTAIL.n45 VSUBS 0.013561f
C815 VTAIL.n46 VSUBS 0.012808f
C816 VTAIL.n47 VSUBS 0.056395f
C817 VTAIL.n48 VSUBS 0.034449f
C818 VTAIL.n49 VSUBS 1.43032f
C819 VTAIL.n50 VSUBS 0.024877f
C820 VTAIL.n51 VSUBS 0.023835f
C821 VTAIL.n52 VSUBS 0.012808f
C822 VTAIL.n53 VSUBS 0.030273f
C823 VTAIL.n54 VSUBS 0.013184f
C824 VTAIL.n55 VSUBS 0.023835f
C825 VTAIL.n56 VSUBS 0.013184f
C826 VTAIL.n57 VSUBS 0.012808f
C827 VTAIL.n58 VSUBS 0.030273f
C828 VTAIL.n59 VSUBS 0.030273f
C829 VTAIL.n60 VSUBS 0.013561f
C830 VTAIL.n61 VSUBS 0.023835f
C831 VTAIL.n62 VSUBS 0.012808f
C832 VTAIL.n63 VSUBS 0.030273f
C833 VTAIL.n64 VSUBS 0.013561f
C834 VTAIL.n65 VSUBS 0.88695f
C835 VTAIL.n66 VSUBS 0.012808f
C836 VTAIL.t2 VSUBS 0.065047f
C837 VTAIL.n67 VSUBS 0.158425f
C838 VTAIL.n68 VSUBS 0.022773f
C839 VTAIL.n69 VSUBS 0.022705f
C840 VTAIL.n70 VSUBS 0.030273f
C841 VTAIL.n71 VSUBS 0.013561f
C842 VTAIL.n72 VSUBS 0.012808f
C843 VTAIL.n73 VSUBS 0.023835f
C844 VTAIL.n74 VSUBS 0.023835f
C845 VTAIL.n75 VSUBS 0.012808f
C846 VTAIL.n76 VSUBS 0.013561f
C847 VTAIL.n77 VSUBS 0.030273f
C848 VTAIL.n78 VSUBS 0.030273f
C849 VTAIL.n79 VSUBS 0.013561f
C850 VTAIL.n80 VSUBS 0.012808f
C851 VTAIL.n81 VSUBS 0.023835f
C852 VTAIL.n82 VSUBS 0.023835f
C853 VTAIL.n83 VSUBS 0.012808f
C854 VTAIL.n84 VSUBS 0.013561f
C855 VTAIL.n85 VSUBS 0.030273f
C856 VTAIL.n86 VSUBS 0.030273f
C857 VTAIL.n87 VSUBS 0.013561f
C858 VTAIL.n88 VSUBS 0.012808f
C859 VTAIL.n89 VSUBS 0.023835f
C860 VTAIL.n90 VSUBS 0.023835f
C861 VTAIL.n91 VSUBS 0.012808f
C862 VTAIL.n92 VSUBS 0.013561f
C863 VTAIL.n93 VSUBS 0.030273f
C864 VTAIL.n94 VSUBS 0.068818f
C865 VTAIL.n95 VSUBS 0.013561f
C866 VTAIL.n96 VSUBS 0.012808f
C867 VTAIL.n97 VSUBS 0.056395f
C868 VTAIL.n98 VSUBS 0.034449f
C869 VTAIL.n99 VSUBS 1.47369f
C870 VTAIL.n100 VSUBS 0.024877f
C871 VTAIL.n101 VSUBS 0.023835f
C872 VTAIL.n102 VSUBS 0.012808f
C873 VTAIL.n103 VSUBS 0.030273f
C874 VTAIL.n104 VSUBS 0.013184f
C875 VTAIL.n105 VSUBS 0.023835f
C876 VTAIL.n106 VSUBS 0.013184f
C877 VTAIL.n107 VSUBS 0.012808f
C878 VTAIL.n108 VSUBS 0.030273f
C879 VTAIL.n109 VSUBS 0.030273f
C880 VTAIL.n110 VSUBS 0.013561f
C881 VTAIL.n111 VSUBS 0.023835f
C882 VTAIL.n112 VSUBS 0.012808f
C883 VTAIL.n113 VSUBS 0.030273f
C884 VTAIL.n114 VSUBS 0.013561f
C885 VTAIL.n115 VSUBS 0.88695f
C886 VTAIL.n116 VSUBS 0.012808f
C887 VTAIL.t0 VSUBS 0.065047f
C888 VTAIL.n117 VSUBS 0.158425f
C889 VTAIL.n118 VSUBS 0.022773f
C890 VTAIL.n119 VSUBS 0.022705f
C891 VTAIL.n120 VSUBS 0.030273f
C892 VTAIL.n121 VSUBS 0.013561f
C893 VTAIL.n122 VSUBS 0.012808f
C894 VTAIL.n123 VSUBS 0.023835f
C895 VTAIL.n124 VSUBS 0.023835f
C896 VTAIL.n125 VSUBS 0.012808f
C897 VTAIL.n126 VSUBS 0.013561f
C898 VTAIL.n127 VSUBS 0.030273f
C899 VTAIL.n128 VSUBS 0.030273f
C900 VTAIL.n129 VSUBS 0.013561f
C901 VTAIL.n130 VSUBS 0.012808f
C902 VTAIL.n131 VSUBS 0.023835f
C903 VTAIL.n132 VSUBS 0.023835f
C904 VTAIL.n133 VSUBS 0.012808f
C905 VTAIL.n134 VSUBS 0.013561f
C906 VTAIL.n135 VSUBS 0.030273f
C907 VTAIL.n136 VSUBS 0.030273f
C908 VTAIL.n137 VSUBS 0.013561f
C909 VTAIL.n138 VSUBS 0.012808f
C910 VTAIL.n139 VSUBS 0.023835f
C911 VTAIL.n140 VSUBS 0.023835f
C912 VTAIL.n141 VSUBS 0.012808f
C913 VTAIL.n142 VSUBS 0.013561f
C914 VTAIL.n143 VSUBS 0.030273f
C915 VTAIL.n144 VSUBS 0.068818f
C916 VTAIL.n145 VSUBS 0.013561f
C917 VTAIL.n146 VSUBS 0.012808f
C918 VTAIL.n147 VSUBS 0.056395f
C919 VTAIL.n148 VSUBS 0.034449f
C920 VTAIL.n149 VSUBS 1.28235f
C921 VTAIL.n150 VSUBS 0.024877f
C922 VTAIL.n151 VSUBS 0.023835f
C923 VTAIL.n152 VSUBS 0.012808f
C924 VTAIL.n153 VSUBS 0.030273f
C925 VTAIL.n154 VSUBS 0.013184f
C926 VTAIL.n155 VSUBS 0.023835f
C927 VTAIL.n156 VSUBS 0.013561f
C928 VTAIL.n157 VSUBS 0.030273f
C929 VTAIL.n158 VSUBS 0.013561f
C930 VTAIL.n159 VSUBS 0.023835f
C931 VTAIL.n160 VSUBS 0.012808f
C932 VTAIL.n161 VSUBS 0.030273f
C933 VTAIL.n162 VSUBS 0.013561f
C934 VTAIL.n163 VSUBS 0.88695f
C935 VTAIL.n164 VSUBS 0.012808f
C936 VTAIL.t3 VSUBS 0.065047f
C937 VTAIL.n165 VSUBS 0.158425f
C938 VTAIL.n166 VSUBS 0.022773f
C939 VTAIL.n167 VSUBS 0.022705f
C940 VTAIL.n168 VSUBS 0.030273f
C941 VTAIL.n169 VSUBS 0.013561f
C942 VTAIL.n170 VSUBS 0.012808f
C943 VTAIL.n171 VSUBS 0.023835f
C944 VTAIL.n172 VSUBS 0.023835f
C945 VTAIL.n173 VSUBS 0.012808f
C946 VTAIL.n174 VSUBS 0.013561f
C947 VTAIL.n175 VSUBS 0.030273f
C948 VTAIL.n176 VSUBS 0.030273f
C949 VTAIL.n177 VSUBS 0.013561f
C950 VTAIL.n178 VSUBS 0.012808f
C951 VTAIL.n179 VSUBS 0.023835f
C952 VTAIL.n180 VSUBS 0.023835f
C953 VTAIL.n181 VSUBS 0.012808f
C954 VTAIL.n182 VSUBS 0.012808f
C955 VTAIL.n183 VSUBS 0.013561f
C956 VTAIL.n184 VSUBS 0.030273f
C957 VTAIL.n185 VSUBS 0.030273f
C958 VTAIL.n186 VSUBS 0.030273f
C959 VTAIL.n187 VSUBS 0.013184f
C960 VTAIL.n188 VSUBS 0.012808f
C961 VTAIL.n189 VSUBS 0.023835f
C962 VTAIL.n190 VSUBS 0.023835f
C963 VTAIL.n191 VSUBS 0.012808f
C964 VTAIL.n192 VSUBS 0.013561f
C965 VTAIL.n193 VSUBS 0.030273f
C966 VTAIL.n194 VSUBS 0.068818f
C967 VTAIL.n195 VSUBS 0.013561f
C968 VTAIL.n196 VSUBS 0.012808f
C969 VTAIL.n197 VSUBS 0.056395f
C970 VTAIL.n198 VSUBS 0.034449f
C971 VTAIL.n199 VSUBS 1.19396f
C972 VN.t0 VSUBS 2.65168f
C973 VN.t1 VSUBS 3.2019f
.ends

