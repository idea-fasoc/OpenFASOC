* NGSPICE file created from diff_pair_sample_0178.ext - technology: sky130A

.subckt diff_pair_sample_0178 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t2 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=1.4388 ps=9.05 w=8.72 l=1.27
X1 VTAIL.t2 VN.t0 VDD2.t5 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=1.4388 ps=9.05 w=8.72 l=1.27
X2 VDD1.t1 VP.t1 VTAIL.t8 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=3.4008 ps=18.22 w=8.72 l=1.27
X3 B.t11 B.t9 B.t10 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=0 ps=0 w=8.72 l=1.27
X4 VDD1.t0 VP.t2 VTAIL.t7 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=1.4388 ps=9.05 w=8.72 l=1.27
X5 VTAIL.t6 VP.t3 VDD1.t5 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=1.4388 ps=9.05 w=8.72 l=1.27
X6 VTAIL.t10 VN.t1 VDD2.t4 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=1.4388 ps=9.05 w=8.72 l=1.27
X7 VDD2.t3 VN.t2 VTAIL.t11 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=3.4008 ps=18.22 w=8.72 l=1.27
X8 VDD1.t4 VP.t4 VTAIL.t5 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=3.4008 ps=18.22 w=8.72 l=1.27
X9 VDD2.t2 VN.t3 VTAIL.t0 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=1.4388 pd=9.05 as=3.4008 ps=18.22 w=8.72 l=1.27
X10 VDD1.t3 VP.t5 VTAIL.t4 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=1.4388 ps=9.05 w=8.72 l=1.27
X11 VDD2.t1 VN.t4 VTAIL.t1 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=1.4388 ps=9.05 w=8.72 l=1.27
X12 B.t8 B.t6 B.t7 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=0 ps=0 w=8.72 l=1.27
X13 B.t5 B.t3 B.t4 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=0 ps=0 w=8.72 l=1.27
X14 VDD2.t0 VN.t5 VTAIL.t3 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=1.4388 ps=9.05 w=8.72 l=1.27
X15 B.t2 B.t0 B.t1 w_n2250_n2712# sky130_fd_pr__pfet_01v8 ad=3.4008 pd=18.22 as=0 ps=0 w=8.72 l=1.27
R0 VP.n5 VP.t2 215.903
R1 VP.n12 VP.t5 196.786
R2 VP.n19 VP.t1 196.786
R3 VP.n9 VP.t4 196.786
R4 VP.n1 VP.t3 165.475
R5 VP.n4 VP.t0 165.475
R6 VP.n7 VP.n6 161.3
R7 VP.n8 VP.n3 161.3
R8 VP.n18 VP.n0 161.3
R9 VP.n17 VP.n16 161.3
R10 VP.n15 VP.n14 161.3
R11 VP.n13 VP.n2 161.3
R12 VP.n10 VP.n9 80.6037
R13 VP.n20 VP.n19 80.6037
R14 VP.n12 VP.n11 80.6037
R15 VP.n5 VP.n4 45.2962
R16 VP.n11 VP.n10 41.1453
R17 VP.n14 VP.n13 35.5419
R18 VP.n18 VP.n17 35.5419
R19 VP.n8 VP.n7 35.5419
R20 VP.n13 VP.n12 31.4035
R21 VP.n19 VP.n18 31.4035
R22 VP.n9 VP.n8 31.4035
R23 VP.n6 VP.n5 29.5285
R24 VP.n14 VP.n1 12.1722
R25 VP.n17 VP.n1 12.1722
R26 VP.n7 VP.n4 12.1722
R27 VP.n10 VP.n3 0.285035
R28 VP.n11 VP.n2 0.285035
R29 VP.n20 VP.n0 0.285035
R30 VP.n6 VP.n3 0.189894
R31 VP.n15 VP.n2 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VP VP.n20 0.146778
R35 VDD1.n40 VDD1.n0 756.745
R36 VDD1.n85 VDD1.n45 756.745
R37 VDD1.n41 VDD1.n40 585
R38 VDD1.n39 VDD1.n38 585
R39 VDD1.n37 VDD1.n3 585
R40 VDD1.n7 VDD1.n4 585
R41 VDD1.n32 VDD1.n31 585
R42 VDD1.n30 VDD1.n29 585
R43 VDD1.n9 VDD1.n8 585
R44 VDD1.n24 VDD1.n23 585
R45 VDD1.n22 VDD1.n21 585
R46 VDD1.n13 VDD1.n12 585
R47 VDD1.n16 VDD1.n15 585
R48 VDD1.n60 VDD1.n59 585
R49 VDD1.n57 VDD1.n56 585
R50 VDD1.n66 VDD1.n65 585
R51 VDD1.n68 VDD1.n67 585
R52 VDD1.n53 VDD1.n52 585
R53 VDD1.n74 VDD1.n73 585
R54 VDD1.n77 VDD1.n76 585
R55 VDD1.n75 VDD1.n49 585
R56 VDD1.n82 VDD1.n48 585
R57 VDD1.n84 VDD1.n83 585
R58 VDD1.n86 VDD1.n85 585
R59 VDD1.t0 VDD1.n14 329.039
R60 VDD1.t3 VDD1.n58 329.038
R61 VDD1.n40 VDD1.n39 171.744
R62 VDD1.n39 VDD1.n3 171.744
R63 VDD1.n7 VDD1.n3 171.744
R64 VDD1.n31 VDD1.n7 171.744
R65 VDD1.n31 VDD1.n30 171.744
R66 VDD1.n30 VDD1.n8 171.744
R67 VDD1.n23 VDD1.n8 171.744
R68 VDD1.n23 VDD1.n22 171.744
R69 VDD1.n22 VDD1.n12 171.744
R70 VDD1.n15 VDD1.n12 171.744
R71 VDD1.n59 VDD1.n56 171.744
R72 VDD1.n66 VDD1.n56 171.744
R73 VDD1.n67 VDD1.n66 171.744
R74 VDD1.n67 VDD1.n52 171.744
R75 VDD1.n74 VDD1.n52 171.744
R76 VDD1.n76 VDD1.n74 171.744
R77 VDD1.n76 VDD1.n75 171.744
R78 VDD1.n75 VDD1.n48 171.744
R79 VDD1.n84 VDD1.n48 171.744
R80 VDD1.n85 VDD1.n84 171.744
R81 VDD1.n15 VDD1.t0 85.8723
R82 VDD1.n59 VDD1.t3 85.8723
R83 VDD1.n91 VDD1.n90 84.4724
R84 VDD1.n93 VDD1.n92 84.1829
R85 VDD1 VDD1.n44 53.8356
R86 VDD1.n91 VDD1.n89 53.7221
R87 VDD1.n93 VDD1.n91 36.988
R88 VDD1.n38 VDD1.n37 13.1884
R89 VDD1.n83 VDD1.n82 13.1884
R90 VDD1.n41 VDD1.n2 12.8005
R91 VDD1.n36 VDD1.n4 12.8005
R92 VDD1.n81 VDD1.n49 12.8005
R93 VDD1.n86 VDD1.n47 12.8005
R94 VDD1.n42 VDD1.n0 12.0247
R95 VDD1.n33 VDD1.n32 12.0247
R96 VDD1.n78 VDD1.n77 12.0247
R97 VDD1.n87 VDD1.n45 12.0247
R98 VDD1.n29 VDD1.n6 11.249
R99 VDD1.n73 VDD1.n51 11.249
R100 VDD1.n16 VDD1.n14 10.7239
R101 VDD1.n60 VDD1.n58 10.7239
R102 VDD1.n28 VDD1.n9 10.4732
R103 VDD1.n72 VDD1.n53 10.4732
R104 VDD1.n25 VDD1.n24 9.69747
R105 VDD1.n69 VDD1.n68 9.69747
R106 VDD1.n44 VDD1.n43 9.45567
R107 VDD1.n89 VDD1.n88 9.45567
R108 VDD1.n18 VDD1.n17 9.3005
R109 VDD1.n20 VDD1.n19 9.3005
R110 VDD1.n11 VDD1.n10 9.3005
R111 VDD1.n26 VDD1.n25 9.3005
R112 VDD1.n28 VDD1.n27 9.3005
R113 VDD1.n6 VDD1.n5 9.3005
R114 VDD1.n34 VDD1.n33 9.3005
R115 VDD1.n36 VDD1.n35 9.3005
R116 VDD1.n43 VDD1.n42 9.3005
R117 VDD1.n2 VDD1.n1 9.3005
R118 VDD1.n88 VDD1.n87 9.3005
R119 VDD1.n47 VDD1.n46 9.3005
R120 VDD1.n62 VDD1.n61 9.3005
R121 VDD1.n64 VDD1.n63 9.3005
R122 VDD1.n55 VDD1.n54 9.3005
R123 VDD1.n70 VDD1.n69 9.3005
R124 VDD1.n72 VDD1.n71 9.3005
R125 VDD1.n51 VDD1.n50 9.3005
R126 VDD1.n79 VDD1.n78 9.3005
R127 VDD1.n81 VDD1.n80 9.3005
R128 VDD1.n21 VDD1.n11 8.92171
R129 VDD1.n65 VDD1.n55 8.92171
R130 VDD1.n20 VDD1.n13 8.14595
R131 VDD1.n64 VDD1.n57 8.14595
R132 VDD1.n17 VDD1.n16 7.3702
R133 VDD1.n61 VDD1.n60 7.3702
R134 VDD1.n17 VDD1.n13 5.81868
R135 VDD1.n61 VDD1.n57 5.81868
R136 VDD1.n21 VDD1.n20 5.04292
R137 VDD1.n65 VDD1.n64 5.04292
R138 VDD1.n24 VDD1.n11 4.26717
R139 VDD1.n68 VDD1.n55 4.26717
R140 VDD1.n92 VDD1.t2 3.72814
R141 VDD1.n92 VDD1.t4 3.72814
R142 VDD1.n90 VDD1.t5 3.72814
R143 VDD1.n90 VDD1.t1 3.72814
R144 VDD1.n25 VDD1.n9 3.49141
R145 VDD1.n69 VDD1.n53 3.49141
R146 VDD1.n29 VDD1.n28 2.71565
R147 VDD1.n73 VDD1.n72 2.71565
R148 VDD1.n18 VDD1.n14 2.41285
R149 VDD1.n62 VDD1.n58 2.41285
R150 VDD1.n44 VDD1.n0 1.93989
R151 VDD1.n32 VDD1.n6 1.93989
R152 VDD1.n77 VDD1.n51 1.93989
R153 VDD1.n89 VDD1.n45 1.93989
R154 VDD1.n42 VDD1.n41 1.16414
R155 VDD1.n33 VDD1.n4 1.16414
R156 VDD1.n78 VDD1.n49 1.16414
R157 VDD1.n87 VDD1.n86 1.16414
R158 VDD1.n38 VDD1.n2 0.388379
R159 VDD1.n37 VDD1.n36 0.388379
R160 VDD1.n82 VDD1.n81 0.388379
R161 VDD1.n83 VDD1.n47 0.388379
R162 VDD1 VDD1.n93 0.287138
R163 VDD1.n43 VDD1.n1 0.155672
R164 VDD1.n35 VDD1.n1 0.155672
R165 VDD1.n35 VDD1.n34 0.155672
R166 VDD1.n34 VDD1.n5 0.155672
R167 VDD1.n27 VDD1.n5 0.155672
R168 VDD1.n27 VDD1.n26 0.155672
R169 VDD1.n26 VDD1.n10 0.155672
R170 VDD1.n19 VDD1.n10 0.155672
R171 VDD1.n19 VDD1.n18 0.155672
R172 VDD1.n63 VDD1.n62 0.155672
R173 VDD1.n63 VDD1.n54 0.155672
R174 VDD1.n70 VDD1.n54 0.155672
R175 VDD1.n71 VDD1.n70 0.155672
R176 VDD1.n71 VDD1.n50 0.155672
R177 VDD1.n79 VDD1.n50 0.155672
R178 VDD1.n80 VDD1.n79 0.155672
R179 VDD1.n80 VDD1.n46 0.155672
R180 VDD1.n88 VDD1.n46 0.155672
R181 VTAIL.n186 VTAIL.n146 756.745
R182 VTAIL.n42 VTAIL.n2 756.745
R183 VTAIL.n140 VTAIL.n100 756.745
R184 VTAIL.n92 VTAIL.n52 756.745
R185 VTAIL.n161 VTAIL.n160 585
R186 VTAIL.n158 VTAIL.n157 585
R187 VTAIL.n167 VTAIL.n166 585
R188 VTAIL.n169 VTAIL.n168 585
R189 VTAIL.n154 VTAIL.n153 585
R190 VTAIL.n175 VTAIL.n174 585
R191 VTAIL.n178 VTAIL.n177 585
R192 VTAIL.n176 VTAIL.n150 585
R193 VTAIL.n183 VTAIL.n149 585
R194 VTAIL.n185 VTAIL.n184 585
R195 VTAIL.n187 VTAIL.n186 585
R196 VTAIL.n17 VTAIL.n16 585
R197 VTAIL.n14 VTAIL.n13 585
R198 VTAIL.n23 VTAIL.n22 585
R199 VTAIL.n25 VTAIL.n24 585
R200 VTAIL.n10 VTAIL.n9 585
R201 VTAIL.n31 VTAIL.n30 585
R202 VTAIL.n34 VTAIL.n33 585
R203 VTAIL.n32 VTAIL.n6 585
R204 VTAIL.n39 VTAIL.n5 585
R205 VTAIL.n41 VTAIL.n40 585
R206 VTAIL.n43 VTAIL.n42 585
R207 VTAIL.n141 VTAIL.n140 585
R208 VTAIL.n139 VTAIL.n138 585
R209 VTAIL.n137 VTAIL.n103 585
R210 VTAIL.n107 VTAIL.n104 585
R211 VTAIL.n132 VTAIL.n131 585
R212 VTAIL.n130 VTAIL.n129 585
R213 VTAIL.n109 VTAIL.n108 585
R214 VTAIL.n124 VTAIL.n123 585
R215 VTAIL.n122 VTAIL.n121 585
R216 VTAIL.n113 VTAIL.n112 585
R217 VTAIL.n116 VTAIL.n115 585
R218 VTAIL.n93 VTAIL.n92 585
R219 VTAIL.n91 VTAIL.n90 585
R220 VTAIL.n89 VTAIL.n55 585
R221 VTAIL.n59 VTAIL.n56 585
R222 VTAIL.n84 VTAIL.n83 585
R223 VTAIL.n82 VTAIL.n81 585
R224 VTAIL.n61 VTAIL.n60 585
R225 VTAIL.n76 VTAIL.n75 585
R226 VTAIL.n74 VTAIL.n73 585
R227 VTAIL.n65 VTAIL.n64 585
R228 VTAIL.n68 VTAIL.n67 585
R229 VTAIL.t5 VTAIL.n114 329.039
R230 VTAIL.t11 VTAIL.n66 329.039
R231 VTAIL.t0 VTAIL.n159 329.038
R232 VTAIL.t8 VTAIL.n15 329.038
R233 VTAIL.n160 VTAIL.n157 171.744
R234 VTAIL.n167 VTAIL.n157 171.744
R235 VTAIL.n168 VTAIL.n167 171.744
R236 VTAIL.n168 VTAIL.n153 171.744
R237 VTAIL.n175 VTAIL.n153 171.744
R238 VTAIL.n177 VTAIL.n175 171.744
R239 VTAIL.n177 VTAIL.n176 171.744
R240 VTAIL.n176 VTAIL.n149 171.744
R241 VTAIL.n185 VTAIL.n149 171.744
R242 VTAIL.n186 VTAIL.n185 171.744
R243 VTAIL.n16 VTAIL.n13 171.744
R244 VTAIL.n23 VTAIL.n13 171.744
R245 VTAIL.n24 VTAIL.n23 171.744
R246 VTAIL.n24 VTAIL.n9 171.744
R247 VTAIL.n31 VTAIL.n9 171.744
R248 VTAIL.n33 VTAIL.n31 171.744
R249 VTAIL.n33 VTAIL.n32 171.744
R250 VTAIL.n32 VTAIL.n5 171.744
R251 VTAIL.n41 VTAIL.n5 171.744
R252 VTAIL.n42 VTAIL.n41 171.744
R253 VTAIL.n140 VTAIL.n139 171.744
R254 VTAIL.n139 VTAIL.n103 171.744
R255 VTAIL.n107 VTAIL.n103 171.744
R256 VTAIL.n131 VTAIL.n107 171.744
R257 VTAIL.n131 VTAIL.n130 171.744
R258 VTAIL.n130 VTAIL.n108 171.744
R259 VTAIL.n123 VTAIL.n108 171.744
R260 VTAIL.n123 VTAIL.n122 171.744
R261 VTAIL.n122 VTAIL.n112 171.744
R262 VTAIL.n115 VTAIL.n112 171.744
R263 VTAIL.n92 VTAIL.n91 171.744
R264 VTAIL.n91 VTAIL.n55 171.744
R265 VTAIL.n59 VTAIL.n55 171.744
R266 VTAIL.n83 VTAIL.n59 171.744
R267 VTAIL.n83 VTAIL.n82 171.744
R268 VTAIL.n82 VTAIL.n60 171.744
R269 VTAIL.n75 VTAIL.n60 171.744
R270 VTAIL.n75 VTAIL.n74 171.744
R271 VTAIL.n74 VTAIL.n64 171.744
R272 VTAIL.n67 VTAIL.n64 171.744
R273 VTAIL.n160 VTAIL.t0 85.8723
R274 VTAIL.n16 VTAIL.t8 85.8723
R275 VTAIL.n115 VTAIL.t5 85.8723
R276 VTAIL.n67 VTAIL.t11 85.8723
R277 VTAIL.n99 VTAIL.n98 67.5043
R278 VTAIL.n51 VTAIL.n50 67.5043
R279 VTAIL.n1 VTAIL.n0 67.5041
R280 VTAIL.n49 VTAIL.n48 67.5041
R281 VTAIL.n191 VTAIL.n190 36.0641
R282 VTAIL.n47 VTAIL.n46 36.0641
R283 VTAIL.n145 VTAIL.n144 36.0641
R284 VTAIL.n97 VTAIL.n96 36.0641
R285 VTAIL.n51 VTAIL.n49 22.6427
R286 VTAIL.n191 VTAIL.n145 21.2634
R287 VTAIL.n184 VTAIL.n183 13.1884
R288 VTAIL.n40 VTAIL.n39 13.1884
R289 VTAIL.n138 VTAIL.n137 13.1884
R290 VTAIL.n90 VTAIL.n89 13.1884
R291 VTAIL.n182 VTAIL.n150 12.8005
R292 VTAIL.n187 VTAIL.n148 12.8005
R293 VTAIL.n38 VTAIL.n6 12.8005
R294 VTAIL.n43 VTAIL.n4 12.8005
R295 VTAIL.n141 VTAIL.n102 12.8005
R296 VTAIL.n136 VTAIL.n104 12.8005
R297 VTAIL.n93 VTAIL.n54 12.8005
R298 VTAIL.n88 VTAIL.n56 12.8005
R299 VTAIL.n179 VTAIL.n178 12.0247
R300 VTAIL.n188 VTAIL.n146 12.0247
R301 VTAIL.n35 VTAIL.n34 12.0247
R302 VTAIL.n44 VTAIL.n2 12.0247
R303 VTAIL.n142 VTAIL.n100 12.0247
R304 VTAIL.n133 VTAIL.n132 12.0247
R305 VTAIL.n94 VTAIL.n52 12.0247
R306 VTAIL.n85 VTAIL.n84 12.0247
R307 VTAIL.n174 VTAIL.n152 11.249
R308 VTAIL.n30 VTAIL.n8 11.249
R309 VTAIL.n129 VTAIL.n106 11.249
R310 VTAIL.n81 VTAIL.n58 11.249
R311 VTAIL.n161 VTAIL.n159 10.7239
R312 VTAIL.n17 VTAIL.n15 10.7239
R313 VTAIL.n116 VTAIL.n114 10.7239
R314 VTAIL.n68 VTAIL.n66 10.7239
R315 VTAIL.n173 VTAIL.n154 10.4732
R316 VTAIL.n29 VTAIL.n10 10.4732
R317 VTAIL.n128 VTAIL.n109 10.4732
R318 VTAIL.n80 VTAIL.n61 10.4732
R319 VTAIL.n170 VTAIL.n169 9.69747
R320 VTAIL.n26 VTAIL.n25 9.69747
R321 VTAIL.n125 VTAIL.n124 9.69747
R322 VTAIL.n77 VTAIL.n76 9.69747
R323 VTAIL.n190 VTAIL.n189 9.45567
R324 VTAIL.n46 VTAIL.n45 9.45567
R325 VTAIL.n144 VTAIL.n143 9.45567
R326 VTAIL.n96 VTAIL.n95 9.45567
R327 VTAIL.n189 VTAIL.n188 9.3005
R328 VTAIL.n148 VTAIL.n147 9.3005
R329 VTAIL.n163 VTAIL.n162 9.3005
R330 VTAIL.n165 VTAIL.n164 9.3005
R331 VTAIL.n156 VTAIL.n155 9.3005
R332 VTAIL.n171 VTAIL.n170 9.3005
R333 VTAIL.n173 VTAIL.n172 9.3005
R334 VTAIL.n152 VTAIL.n151 9.3005
R335 VTAIL.n180 VTAIL.n179 9.3005
R336 VTAIL.n182 VTAIL.n181 9.3005
R337 VTAIL.n45 VTAIL.n44 9.3005
R338 VTAIL.n4 VTAIL.n3 9.3005
R339 VTAIL.n19 VTAIL.n18 9.3005
R340 VTAIL.n21 VTAIL.n20 9.3005
R341 VTAIL.n12 VTAIL.n11 9.3005
R342 VTAIL.n27 VTAIL.n26 9.3005
R343 VTAIL.n29 VTAIL.n28 9.3005
R344 VTAIL.n8 VTAIL.n7 9.3005
R345 VTAIL.n36 VTAIL.n35 9.3005
R346 VTAIL.n38 VTAIL.n37 9.3005
R347 VTAIL.n118 VTAIL.n117 9.3005
R348 VTAIL.n120 VTAIL.n119 9.3005
R349 VTAIL.n111 VTAIL.n110 9.3005
R350 VTAIL.n126 VTAIL.n125 9.3005
R351 VTAIL.n128 VTAIL.n127 9.3005
R352 VTAIL.n106 VTAIL.n105 9.3005
R353 VTAIL.n134 VTAIL.n133 9.3005
R354 VTAIL.n136 VTAIL.n135 9.3005
R355 VTAIL.n143 VTAIL.n142 9.3005
R356 VTAIL.n102 VTAIL.n101 9.3005
R357 VTAIL.n70 VTAIL.n69 9.3005
R358 VTAIL.n72 VTAIL.n71 9.3005
R359 VTAIL.n63 VTAIL.n62 9.3005
R360 VTAIL.n78 VTAIL.n77 9.3005
R361 VTAIL.n80 VTAIL.n79 9.3005
R362 VTAIL.n58 VTAIL.n57 9.3005
R363 VTAIL.n86 VTAIL.n85 9.3005
R364 VTAIL.n88 VTAIL.n87 9.3005
R365 VTAIL.n95 VTAIL.n94 9.3005
R366 VTAIL.n54 VTAIL.n53 9.3005
R367 VTAIL.n166 VTAIL.n156 8.92171
R368 VTAIL.n22 VTAIL.n12 8.92171
R369 VTAIL.n121 VTAIL.n111 8.92171
R370 VTAIL.n73 VTAIL.n63 8.92171
R371 VTAIL.n165 VTAIL.n158 8.14595
R372 VTAIL.n21 VTAIL.n14 8.14595
R373 VTAIL.n120 VTAIL.n113 8.14595
R374 VTAIL.n72 VTAIL.n65 8.14595
R375 VTAIL.n162 VTAIL.n161 7.3702
R376 VTAIL.n18 VTAIL.n17 7.3702
R377 VTAIL.n117 VTAIL.n116 7.3702
R378 VTAIL.n69 VTAIL.n68 7.3702
R379 VTAIL.n162 VTAIL.n158 5.81868
R380 VTAIL.n18 VTAIL.n14 5.81868
R381 VTAIL.n117 VTAIL.n113 5.81868
R382 VTAIL.n69 VTAIL.n65 5.81868
R383 VTAIL.n166 VTAIL.n165 5.04292
R384 VTAIL.n22 VTAIL.n21 5.04292
R385 VTAIL.n121 VTAIL.n120 5.04292
R386 VTAIL.n73 VTAIL.n72 5.04292
R387 VTAIL.n169 VTAIL.n156 4.26717
R388 VTAIL.n25 VTAIL.n12 4.26717
R389 VTAIL.n124 VTAIL.n111 4.26717
R390 VTAIL.n76 VTAIL.n63 4.26717
R391 VTAIL.n0 VTAIL.t3 3.72814
R392 VTAIL.n0 VTAIL.t10 3.72814
R393 VTAIL.n48 VTAIL.t4 3.72814
R394 VTAIL.n48 VTAIL.t6 3.72814
R395 VTAIL.n98 VTAIL.t7 3.72814
R396 VTAIL.n98 VTAIL.t9 3.72814
R397 VTAIL.n50 VTAIL.t1 3.72814
R398 VTAIL.n50 VTAIL.t2 3.72814
R399 VTAIL.n170 VTAIL.n154 3.49141
R400 VTAIL.n26 VTAIL.n10 3.49141
R401 VTAIL.n125 VTAIL.n109 3.49141
R402 VTAIL.n77 VTAIL.n61 3.49141
R403 VTAIL.n174 VTAIL.n173 2.71565
R404 VTAIL.n30 VTAIL.n29 2.71565
R405 VTAIL.n129 VTAIL.n128 2.71565
R406 VTAIL.n81 VTAIL.n80 2.71565
R407 VTAIL.n163 VTAIL.n159 2.41285
R408 VTAIL.n19 VTAIL.n15 2.41285
R409 VTAIL.n118 VTAIL.n114 2.41285
R410 VTAIL.n70 VTAIL.n66 2.41285
R411 VTAIL.n178 VTAIL.n152 1.93989
R412 VTAIL.n190 VTAIL.n146 1.93989
R413 VTAIL.n34 VTAIL.n8 1.93989
R414 VTAIL.n46 VTAIL.n2 1.93989
R415 VTAIL.n144 VTAIL.n100 1.93989
R416 VTAIL.n132 VTAIL.n106 1.93989
R417 VTAIL.n96 VTAIL.n52 1.93989
R418 VTAIL.n84 VTAIL.n58 1.93989
R419 VTAIL.n97 VTAIL.n51 1.37981
R420 VTAIL.n145 VTAIL.n99 1.37981
R421 VTAIL.n49 VTAIL.n47 1.37981
R422 VTAIL.n179 VTAIL.n150 1.16414
R423 VTAIL.n188 VTAIL.n187 1.16414
R424 VTAIL.n35 VTAIL.n6 1.16414
R425 VTAIL.n44 VTAIL.n43 1.16414
R426 VTAIL.n142 VTAIL.n141 1.16414
R427 VTAIL.n133 VTAIL.n104 1.16414
R428 VTAIL.n94 VTAIL.n93 1.16414
R429 VTAIL.n85 VTAIL.n56 1.16414
R430 VTAIL.n99 VTAIL.n97 1.15998
R431 VTAIL.n47 VTAIL.n1 1.15998
R432 VTAIL VTAIL.n191 0.976793
R433 VTAIL VTAIL.n1 0.403517
R434 VTAIL.n183 VTAIL.n182 0.388379
R435 VTAIL.n184 VTAIL.n148 0.388379
R436 VTAIL.n39 VTAIL.n38 0.388379
R437 VTAIL.n40 VTAIL.n4 0.388379
R438 VTAIL.n138 VTAIL.n102 0.388379
R439 VTAIL.n137 VTAIL.n136 0.388379
R440 VTAIL.n90 VTAIL.n54 0.388379
R441 VTAIL.n89 VTAIL.n88 0.388379
R442 VTAIL.n164 VTAIL.n163 0.155672
R443 VTAIL.n164 VTAIL.n155 0.155672
R444 VTAIL.n171 VTAIL.n155 0.155672
R445 VTAIL.n172 VTAIL.n171 0.155672
R446 VTAIL.n172 VTAIL.n151 0.155672
R447 VTAIL.n180 VTAIL.n151 0.155672
R448 VTAIL.n181 VTAIL.n180 0.155672
R449 VTAIL.n181 VTAIL.n147 0.155672
R450 VTAIL.n189 VTAIL.n147 0.155672
R451 VTAIL.n20 VTAIL.n19 0.155672
R452 VTAIL.n20 VTAIL.n11 0.155672
R453 VTAIL.n27 VTAIL.n11 0.155672
R454 VTAIL.n28 VTAIL.n27 0.155672
R455 VTAIL.n28 VTAIL.n7 0.155672
R456 VTAIL.n36 VTAIL.n7 0.155672
R457 VTAIL.n37 VTAIL.n36 0.155672
R458 VTAIL.n37 VTAIL.n3 0.155672
R459 VTAIL.n45 VTAIL.n3 0.155672
R460 VTAIL.n143 VTAIL.n101 0.155672
R461 VTAIL.n135 VTAIL.n101 0.155672
R462 VTAIL.n135 VTAIL.n134 0.155672
R463 VTAIL.n134 VTAIL.n105 0.155672
R464 VTAIL.n127 VTAIL.n105 0.155672
R465 VTAIL.n127 VTAIL.n126 0.155672
R466 VTAIL.n126 VTAIL.n110 0.155672
R467 VTAIL.n119 VTAIL.n110 0.155672
R468 VTAIL.n119 VTAIL.n118 0.155672
R469 VTAIL.n95 VTAIL.n53 0.155672
R470 VTAIL.n87 VTAIL.n53 0.155672
R471 VTAIL.n87 VTAIL.n86 0.155672
R472 VTAIL.n86 VTAIL.n57 0.155672
R473 VTAIL.n79 VTAIL.n57 0.155672
R474 VTAIL.n79 VTAIL.n78 0.155672
R475 VTAIL.n78 VTAIL.n62 0.155672
R476 VTAIL.n71 VTAIL.n62 0.155672
R477 VTAIL.n71 VTAIL.n70 0.155672
R478 VN.n2 VN.t5 215.903
R479 VN.n10 VN.t2 215.903
R480 VN.n6 VN.t3 196.786
R481 VN.n14 VN.t4 196.786
R482 VN.n1 VN.t1 165.475
R483 VN.n9 VN.t0 165.475
R484 VN.n13 VN.n8 161.3
R485 VN.n12 VN.n11 161.3
R486 VN.n5 VN.n0 161.3
R487 VN.n4 VN.n3 161.3
R488 VN.n15 VN.n14 80.6037
R489 VN.n7 VN.n6 80.6037
R490 VN.n2 VN.n1 45.2962
R491 VN.n10 VN.n9 45.2962
R492 VN VN.n15 41.4309
R493 VN.n5 VN.n4 35.5419
R494 VN.n13 VN.n12 35.5419
R495 VN.n6 VN.n5 31.4035
R496 VN.n14 VN.n13 31.4035
R497 VN.n11 VN.n10 29.5285
R498 VN.n3 VN.n2 29.5285
R499 VN.n4 VN.n1 12.1722
R500 VN.n12 VN.n9 12.1722
R501 VN.n15 VN.n8 0.285035
R502 VN.n7 VN.n0 0.285035
R503 VN.n11 VN.n8 0.189894
R504 VN.n3 VN.n0 0.189894
R505 VN VN.n7 0.146778
R506 VDD2.n87 VDD2.n47 756.745
R507 VDD2.n40 VDD2.n0 756.745
R508 VDD2.n88 VDD2.n87 585
R509 VDD2.n86 VDD2.n85 585
R510 VDD2.n84 VDD2.n50 585
R511 VDD2.n54 VDD2.n51 585
R512 VDD2.n79 VDD2.n78 585
R513 VDD2.n77 VDD2.n76 585
R514 VDD2.n56 VDD2.n55 585
R515 VDD2.n71 VDD2.n70 585
R516 VDD2.n69 VDD2.n68 585
R517 VDD2.n60 VDD2.n59 585
R518 VDD2.n63 VDD2.n62 585
R519 VDD2.n15 VDD2.n14 585
R520 VDD2.n12 VDD2.n11 585
R521 VDD2.n21 VDD2.n20 585
R522 VDD2.n23 VDD2.n22 585
R523 VDD2.n8 VDD2.n7 585
R524 VDD2.n29 VDD2.n28 585
R525 VDD2.n32 VDD2.n31 585
R526 VDD2.n30 VDD2.n4 585
R527 VDD2.n37 VDD2.n3 585
R528 VDD2.n39 VDD2.n38 585
R529 VDD2.n41 VDD2.n40 585
R530 VDD2.t1 VDD2.n61 329.039
R531 VDD2.t0 VDD2.n13 329.038
R532 VDD2.n87 VDD2.n86 171.744
R533 VDD2.n86 VDD2.n50 171.744
R534 VDD2.n54 VDD2.n50 171.744
R535 VDD2.n78 VDD2.n54 171.744
R536 VDD2.n78 VDD2.n77 171.744
R537 VDD2.n77 VDD2.n55 171.744
R538 VDD2.n70 VDD2.n55 171.744
R539 VDD2.n70 VDD2.n69 171.744
R540 VDD2.n69 VDD2.n59 171.744
R541 VDD2.n62 VDD2.n59 171.744
R542 VDD2.n14 VDD2.n11 171.744
R543 VDD2.n21 VDD2.n11 171.744
R544 VDD2.n22 VDD2.n21 171.744
R545 VDD2.n22 VDD2.n7 171.744
R546 VDD2.n29 VDD2.n7 171.744
R547 VDD2.n31 VDD2.n29 171.744
R548 VDD2.n31 VDD2.n30 171.744
R549 VDD2.n30 VDD2.n3 171.744
R550 VDD2.n39 VDD2.n3 171.744
R551 VDD2.n40 VDD2.n39 171.744
R552 VDD2.n62 VDD2.t1 85.8723
R553 VDD2.n14 VDD2.t0 85.8723
R554 VDD2.n46 VDD2.n45 84.4724
R555 VDD2 VDD2.n93 84.4695
R556 VDD2.n46 VDD2.n44 53.7221
R557 VDD2.n92 VDD2.n91 52.7429
R558 VDD2.n92 VDD2.n46 35.7153
R559 VDD2.n85 VDD2.n84 13.1884
R560 VDD2.n38 VDD2.n37 13.1884
R561 VDD2.n88 VDD2.n49 12.8005
R562 VDD2.n83 VDD2.n51 12.8005
R563 VDD2.n36 VDD2.n4 12.8005
R564 VDD2.n41 VDD2.n2 12.8005
R565 VDD2.n89 VDD2.n47 12.0247
R566 VDD2.n80 VDD2.n79 12.0247
R567 VDD2.n33 VDD2.n32 12.0247
R568 VDD2.n42 VDD2.n0 12.0247
R569 VDD2.n76 VDD2.n53 11.249
R570 VDD2.n28 VDD2.n6 11.249
R571 VDD2.n63 VDD2.n61 10.7239
R572 VDD2.n15 VDD2.n13 10.7239
R573 VDD2.n75 VDD2.n56 10.4732
R574 VDD2.n27 VDD2.n8 10.4732
R575 VDD2.n72 VDD2.n71 9.69747
R576 VDD2.n24 VDD2.n23 9.69747
R577 VDD2.n91 VDD2.n90 9.45567
R578 VDD2.n44 VDD2.n43 9.45567
R579 VDD2.n65 VDD2.n64 9.3005
R580 VDD2.n67 VDD2.n66 9.3005
R581 VDD2.n58 VDD2.n57 9.3005
R582 VDD2.n73 VDD2.n72 9.3005
R583 VDD2.n75 VDD2.n74 9.3005
R584 VDD2.n53 VDD2.n52 9.3005
R585 VDD2.n81 VDD2.n80 9.3005
R586 VDD2.n83 VDD2.n82 9.3005
R587 VDD2.n90 VDD2.n89 9.3005
R588 VDD2.n49 VDD2.n48 9.3005
R589 VDD2.n43 VDD2.n42 9.3005
R590 VDD2.n2 VDD2.n1 9.3005
R591 VDD2.n17 VDD2.n16 9.3005
R592 VDD2.n19 VDD2.n18 9.3005
R593 VDD2.n10 VDD2.n9 9.3005
R594 VDD2.n25 VDD2.n24 9.3005
R595 VDD2.n27 VDD2.n26 9.3005
R596 VDD2.n6 VDD2.n5 9.3005
R597 VDD2.n34 VDD2.n33 9.3005
R598 VDD2.n36 VDD2.n35 9.3005
R599 VDD2.n68 VDD2.n58 8.92171
R600 VDD2.n20 VDD2.n10 8.92171
R601 VDD2.n67 VDD2.n60 8.14595
R602 VDD2.n19 VDD2.n12 8.14595
R603 VDD2.n64 VDD2.n63 7.3702
R604 VDD2.n16 VDD2.n15 7.3702
R605 VDD2.n64 VDD2.n60 5.81868
R606 VDD2.n16 VDD2.n12 5.81868
R607 VDD2.n68 VDD2.n67 5.04292
R608 VDD2.n20 VDD2.n19 5.04292
R609 VDD2.n71 VDD2.n58 4.26717
R610 VDD2.n23 VDD2.n10 4.26717
R611 VDD2.n93 VDD2.t5 3.72814
R612 VDD2.n93 VDD2.t3 3.72814
R613 VDD2.n45 VDD2.t4 3.72814
R614 VDD2.n45 VDD2.t2 3.72814
R615 VDD2.n72 VDD2.n56 3.49141
R616 VDD2.n24 VDD2.n8 3.49141
R617 VDD2.n76 VDD2.n75 2.71565
R618 VDD2.n28 VDD2.n27 2.71565
R619 VDD2.n65 VDD2.n61 2.41285
R620 VDD2.n17 VDD2.n13 2.41285
R621 VDD2.n91 VDD2.n47 1.93989
R622 VDD2.n79 VDD2.n53 1.93989
R623 VDD2.n32 VDD2.n6 1.93989
R624 VDD2.n44 VDD2.n0 1.93989
R625 VDD2.n89 VDD2.n88 1.16414
R626 VDD2.n80 VDD2.n51 1.16414
R627 VDD2.n33 VDD2.n4 1.16414
R628 VDD2.n42 VDD2.n41 1.16414
R629 VDD2 VDD2.n92 1.09317
R630 VDD2.n85 VDD2.n49 0.388379
R631 VDD2.n84 VDD2.n83 0.388379
R632 VDD2.n37 VDD2.n36 0.388379
R633 VDD2.n38 VDD2.n2 0.388379
R634 VDD2.n90 VDD2.n48 0.155672
R635 VDD2.n82 VDD2.n48 0.155672
R636 VDD2.n82 VDD2.n81 0.155672
R637 VDD2.n81 VDD2.n52 0.155672
R638 VDD2.n74 VDD2.n52 0.155672
R639 VDD2.n74 VDD2.n73 0.155672
R640 VDD2.n73 VDD2.n57 0.155672
R641 VDD2.n66 VDD2.n57 0.155672
R642 VDD2.n66 VDD2.n65 0.155672
R643 VDD2.n18 VDD2.n17 0.155672
R644 VDD2.n18 VDD2.n9 0.155672
R645 VDD2.n25 VDD2.n9 0.155672
R646 VDD2.n26 VDD2.n25 0.155672
R647 VDD2.n26 VDD2.n5 0.155672
R648 VDD2.n34 VDD2.n5 0.155672
R649 VDD2.n35 VDD2.n34 0.155672
R650 VDD2.n35 VDD2.n1 0.155672
R651 VDD2.n43 VDD2.n1 0.155672
R652 B.n374 B.n57 585
R653 B.n376 B.n375 585
R654 B.n377 B.n56 585
R655 B.n379 B.n378 585
R656 B.n380 B.n55 585
R657 B.n382 B.n381 585
R658 B.n383 B.n54 585
R659 B.n385 B.n384 585
R660 B.n386 B.n53 585
R661 B.n388 B.n387 585
R662 B.n389 B.n52 585
R663 B.n391 B.n390 585
R664 B.n392 B.n51 585
R665 B.n394 B.n393 585
R666 B.n395 B.n50 585
R667 B.n397 B.n396 585
R668 B.n398 B.n49 585
R669 B.n400 B.n399 585
R670 B.n401 B.n48 585
R671 B.n403 B.n402 585
R672 B.n404 B.n47 585
R673 B.n406 B.n405 585
R674 B.n407 B.n46 585
R675 B.n409 B.n408 585
R676 B.n410 B.n45 585
R677 B.n412 B.n411 585
R678 B.n413 B.n44 585
R679 B.n415 B.n414 585
R680 B.n416 B.n43 585
R681 B.n418 B.n417 585
R682 B.n419 B.n39 585
R683 B.n421 B.n420 585
R684 B.n422 B.n38 585
R685 B.n424 B.n423 585
R686 B.n425 B.n37 585
R687 B.n427 B.n426 585
R688 B.n428 B.n36 585
R689 B.n430 B.n429 585
R690 B.n431 B.n35 585
R691 B.n433 B.n432 585
R692 B.n434 B.n34 585
R693 B.n436 B.n435 585
R694 B.n438 B.n31 585
R695 B.n440 B.n439 585
R696 B.n441 B.n30 585
R697 B.n443 B.n442 585
R698 B.n444 B.n29 585
R699 B.n446 B.n445 585
R700 B.n447 B.n28 585
R701 B.n449 B.n448 585
R702 B.n450 B.n27 585
R703 B.n452 B.n451 585
R704 B.n453 B.n26 585
R705 B.n455 B.n454 585
R706 B.n456 B.n25 585
R707 B.n458 B.n457 585
R708 B.n459 B.n24 585
R709 B.n461 B.n460 585
R710 B.n462 B.n23 585
R711 B.n464 B.n463 585
R712 B.n465 B.n22 585
R713 B.n467 B.n466 585
R714 B.n468 B.n21 585
R715 B.n470 B.n469 585
R716 B.n471 B.n20 585
R717 B.n473 B.n472 585
R718 B.n474 B.n19 585
R719 B.n476 B.n475 585
R720 B.n477 B.n18 585
R721 B.n479 B.n478 585
R722 B.n480 B.n17 585
R723 B.n482 B.n481 585
R724 B.n483 B.n16 585
R725 B.n485 B.n484 585
R726 B.n373 B.n372 585
R727 B.n371 B.n58 585
R728 B.n370 B.n369 585
R729 B.n368 B.n59 585
R730 B.n367 B.n366 585
R731 B.n365 B.n60 585
R732 B.n364 B.n363 585
R733 B.n362 B.n61 585
R734 B.n361 B.n360 585
R735 B.n359 B.n62 585
R736 B.n358 B.n357 585
R737 B.n356 B.n63 585
R738 B.n355 B.n354 585
R739 B.n353 B.n64 585
R740 B.n352 B.n351 585
R741 B.n350 B.n65 585
R742 B.n349 B.n348 585
R743 B.n347 B.n66 585
R744 B.n346 B.n345 585
R745 B.n344 B.n67 585
R746 B.n343 B.n342 585
R747 B.n341 B.n68 585
R748 B.n340 B.n339 585
R749 B.n338 B.n69 585
R750 B.n337 B.n336 585
R751 B.n335 B.n70 585
R752 B.n334 B.n333 585
R753 B.n332 B.n71 585
R754 B.n331 B.n330 585
R755 B.n329 B.n72 585
R756 B.n328 B.n327 585
R757 B.n326 B.n73 585
R758 B.n325 B.n324 585
R759 B.n323 B.n74 585
R760 B.n322 B.n321 585
R761 B.n320 B.n75 585
R762 B.n319 B.n318 585
R763 B.n317 B.n76 585
R764 B.n316 B.n315 585
R765 B.n314 B.n77 585
R766 B.n313 B.n312 585
R767 B.n311 B.n78 585
R768 B.n310 B.n309 585
R769 B.n308 B.n79 585
R770 B.n307 B.n306 585
R771 B.n305 B.n80 585
R772 B.n304 B.n303 585
R773 B.n302 B.n81 585
R774 B.n301 B.n300 585
R775 B.n299 B.n82 585
R776 B.n298 B.n297 585
R777 B.n296 B.n83 585
R778 B.n295 B.n294 585
R779 B.n293 B.n84 585
R780 B.n292 B.n291 585
R781 B.n179 B.n126 585
R782 B.n181 B.n180 585
R783 B.n182 B.n125 585
R784 B.n184 B.n183 585
R785 B.n185 B.n124 585
R786 B.n187 B.n186 585
R787 B.n188 B.n123 585
R788 B.n190 B.n189 585
R789 B.n191 B.n122 585
R790 B.n193 B.n192 585
R791 B.n194 B.n121 585
R792 B.n196 B.n195 585
R793 B.n197 B.n120 585
R794 B.n199 B.n198 585
R795 B.n200 B.n119 585
R796 B.n202 B.n201 585
R797 B.n203 B.n118 585
R798 B.n205 B.n204 585
R799 B.n206 B.n117 585
R800 B.n208 B.n207 585
R801 B.n209 B.n116 585
R802 B.n211 B.n210 585
R803 B.n212 B.n115 585
R804 B.n214 B.n213 585
R805 B.n215 B.n114 585
R806 B.n217 B.n216 585
R807 B.n218 B.n113 585
R808 B.n220 B.n219 585
R809 B.n221 B.n112 585
R810 B.n223 B.n222 585
R811 B.n224 B.n111 585
R812 B.n226 B.n225 585
R813 B.n228 B.n108 585
R814 B.n230 B.n229 585
R815 B.n231 B.n107 585
R816 B.n233 B.n232 585
R817 B.n234 B.n106 585
R818 B.n236 B.n235 585
R819 B.n237 B.n105 585
R820 B.n239 B.n238 585
R821 B.n240 B.n104 585
R822 B.n242 B.n241 585
R823 B.n244 B.n243 585
R824 B.n245 B.n100 585
R825 B.n247 B.n246 585
R826 B.n248 B.n99 585
R827 B.n250 B.n249 585
R828 B.n251 B.n98 585
R829 B.n253 B.n252 585
R830 B.n254 B.n97 585
R831 B.n256 B.n255 585
R832 B.n257 B.n96 585
R833 B.n259 B.n258 585
R834 B.n260 B.n95 585
R835 B.n262 B.n261 585
R836 B.n263 B.n94 585
R837 B.n265 B.n264 585
R838 B.n266 B.n93 585
R839 B.n268 B.n267 585
R840 B.n269 B.n92 585
R841 B.n271 B.n270 585
R842 B.n272 B.n91 585
R843 B.n274 B.n273 585
R844 B.n275 B.n90 585
R845 B.n277 B.n276 585
R846 B.n278 B.n89 585
R847 B.n280 B.n279 585
R848 B.n281 B.n88 585
R849 B.n283 B.n282 585
R850 B.n284 B.n87 585
R851 B.n286 B.n285 585
R852 B.n287 B.n86 585
R853 B.n289 B.n288 585
R854 B.n290 B.n85 585
R855 B.n178 B.n177 585
R856 B.n176 B.n127 585
R857 B.n175 B.n174 585
R858 B.n173 B.n128 585
R859 B.n172 B.n171 585
R860 B.n170 B.n129 585
R861 B.n169 B.n168 585
R862 B.n167 B.n130 585
R863 B.n166 B.n165 585
R864 B.n164 B.n131 585
R865 B.n163 B.n162 585
R866 B.n161 B.n132 585
R867 B.n160 B.n159 585
R868 B.n158 B.n133 585
R869 B.n157 B.n156 585
R870 B.n155 B.n134 585
R871 B.n154 B.n153 585
R872 B.n152 B.n135 585
R873 B.n151 B.n150 585
R874 B.n149 B.n136 585
R875 B.n148 B.n147 585
R876 B.n146 B.n137 585
R877 B.n145 B.n144 585
R878 B.n143 B.n138 585
R879 B.n142 B.n141 585
R880 B.n140 B.n139 585
R881 B.n2 B.n0 585
R882 B.n525 B.n1 585
R883 B.n524 B.n523 585
R884 B.n522 B.n3 585
R885 B.n521 B.n520 585
R886 B.n519 B.n4 585
R887 B.n518 B.n517 585
R888 B.n516 B.n5 585
R889 B.n515 B.n514 585
R890 B.n513 B.n6 585
R891 B.n512 B.n511 585
R892 B.n510 B.n7 585
R893 B.n509 B.n508 585
R894 B.n507 B.n8 585
R895 B.n506 B.n505 585
R896 B.n504 B.n9 585
R897 B.n503 B.n502 585
R898 B.n501 B.n10 585
R899 B.n500 B.n499 585
R900 B.n498 B.n11 585
R901 B.n497 B.n496 585
R902 B.n495 B.n12 585
R903 B.n494 B.n493 585
R904 B.n492 B.n13 585
R905 B.n491 B.n490 585
R906 B.n489 B.n14 585
R907 B.n488 B.n487 585
R908 B.n486 B.n15 585
R909 B.n527 B.n526 585
R910 B.n177 B.n126 449.257
R911 B.n484 B.n15 449.257
R912 B.n291 B.n290 449.257
R913 B.n374 B.n373 449.257
R914 B.n101 B.t0 369.942
R915 B.n109 B.t9 369.942
R916 B.n32 B.t6 369.942
R917 B.n40 B.t3 369.942
R918 B.n101 B.t2 347.7
R919 B.n40 B.t4 347.7
R920 B.n109 B.t11 347.7
R921 B.n32 B.t7 347.7
R922 B.n102 B.t1 316.671
R923 B.n41 B.t5 316.671
R924 B.n110 B.t10 316.671
R925 B.n33 B.t8 316.671
R926 B.n177 B.n176 163.367
R927 B.n176 B.n175 163.367
R928 B.n175 B.n128 163.367
R929 B.n171 B.n128 163.367
R930 B.n171 B.n170 163.367
R931 B.n170 B.n169 163.367
R932 B.n169 B.n130 163.367
R933 B.n165 B.n130 163.367
R934 B.n165 B.n164 163.367
R935 B.n164 B.n163 163.367
R936 B.n163 B.n132 163.367
R937 B.n159 B.n132 163.367
R938 B.n159 B.n158 163.367
R939 B.n158 B.n157 163.367
R940 B.n157 B.n134 163.367
R941 B.n153 B.n134 163.367
R942 B.n153 B.n152 163.367
R943 B.n152 B.n151 163.367
R944 B.n151 B.n136 163.367
R945 B.n147 B.n136 163.367
R946 B.n147 B.n146 163.367
R947 B.n146 B.n145 163.367
R948 B.n145 B.n138 163.367
R949 B.n141 B.n138 163.367
R950 B.n141 B.n140 163.367
R951 B.n140 B.n2 163.367
R952 B.n526 B.n2 163.367
R953 B.n526 B.n525 163.367
R954 B.n525 B.n524 163.367
R955 B.n524 B.n3 163.367
R956 B.n520 B.n3 163.367
R957 B.n520 B.n519 163.367
R958 B.n519 B.n518 163.367
R959 B.n518 B.n5 163.367
R960 B.n514 B.n5 163.367
R961 B.n514 B.n513 163.367
R962 B.n513 B.n512 163.367
R963 B.n512 B.n7 163.367
R964 B.n508 B.n7 163.367
R965 B.n508 B.n507 163.367
R966 B.n507 B.n506 163.367
R967 B.n506 B.n9 163.367
R968 B.n502 B.n9 163.367
R969 B.n502 B.n501 163.367
R970 B.n501 B.n500 163.367
R971 B.n500 B.n11 163.367
R972 B.n496 B.n11 163.367
R973 B.n496 B.n495 163.367
R974 B.n495 B.n494 163.367
R975 B.n494 B.n13 163.367
R976 B.n490 B.n13 163.367
R977 B.n490 B.n489 163.367
R978 B.n489 B.n488 163.367
R979 B.n488 B.n15 163.367
R980 B.n181 B.n126 163.367
R981 B.n182 B.n181 163.367
R982 B.n183 B.n182 163.367
R983 B.n183 B.n124 163.367
R984 B.n187 B.n124 163.367
R985 B.n188 B.n187 163.367
R986 B.n189 B.n188 163.367
R987 B.n189 B.n122 163.367
R988 B.n193 B.n122 163.367
R989 B.n194 B.n193 163.367
R990 B.n195 B.n194 163.367
R991 B.n195 B.n120 163.367
R992 B.n199 B.n120 163.367
R993 B.n200 B.n199 163.367
R994 B.n201 B.n200 163.367
R995 B.n201 B.n118 163.367
R996 B.n205 B.n118 163.367
R997 B.n206 B.n205 163.367
R998 B.n207 B.n206 163.367
R999 B.n207 B.n116 163.367
R1000 B.n211 B.n116 163.367
R1001 B.n212 B.n211 163.367
R1002 B.n213 B.n212 163.367
R1003 B.n213 B.n114 163.367
R1004 B.n217 B.n114 163.367
R1005 B.n218 B.n217 163.367
R1006 B.n219 B.n218 163.367
R1007 B.n219 B.n112 163.367
R1008 B.n223 B.n112 163.367
R1009 B.n224 B.n223 163.367
R1010 B.n225 B.n224 163.367
R1011 B.n225 B.n108 163.367
R1012 B.n230 B.n108 163.367
R1013 B.n231 B.n230 163.367
R1014 B.n232 B.n231 163.367
R1015 B.n232 B.n106 163.367
R1016 B.n236 B.n106 163.367
R1017 B.n237 B.n236 163.367
R1018 B.n238 B.n237 163.367
R1019 B.n238 B.n104 163.367
R1020 B.n242 B.n104 163.367
R1021 B.n243 B.n242 163.367
R1022 B.n243 B.n100 163.367
R1023 B.n247 B.n100 163.367
R1024 B.n248 B.n247 163.367
R1025 B.n249 B.n248 163.367
R1026 B.n249 B.n98 163.367
R1027 B.n253 B.n98 163.367
R1028 B.n254 B.n253 163.367
R1029 B.n255 B.n254 163.367
R1030 B.n255 B.n96 163.367
R1031 B.n259 B.n96 163.367
R1032 B.n260 B.n259 163.367
R1033 B.n261 B.n260 163.367
R1034 B.n261 B.n94 163.367
R1035 B.n265 B.n94 163.367
R1036 B.n266 B.n265 163.367
R1037 B.n267 B.n266 163.367
R1038 B.n267 B.n92 163.367
R1039 B.n271 B.n92 163.367
R1040 B.n272 B.n271 163.367
R1041 B.n273 B.n272 163.367
R1042 B.n273 B.n90 163.367
R1043 B.n277 B.n90 163.367
R1044 B.n278 B.n277 163.367
R1045 B.n279 B.n278 163.367
R1046 B.n279 B.n88 163.367
R1047 B.n283 B.n88 163.367
R1048 B.n284 B.n283 163.367
R1049 B.n285 B.n284 163.367
R1050 B.n285 B.n86 163.367
R1051 B.n289 B.n86 163.367
R1052 B.n290 B.n289 163.367
R1053 B.n291 B.n84 163.367
R1054 B.n295 B.n84 163.367
R1055 B.n296 B.n295 163.367
R1056 B.n297 B.n296 163.367
R1057 B.n297 B.n82 163.367
R1058 B.n301 B.n82 163.367
R1059 B.n302 B.n301 163.367
R1060 B.n303 B.n302 163.367
R1061 B.n303 B.n80 163.367
R1062 B.n307 B.n80 163.367
R1063 B.n308 B.n307 163.367
R1064 B.n309 B.n308 163.367
R1065 B.n309 B.n78 163.367
R1066 B.n313 B.n78 163.367
R1067 B.n314 B.n313 163.367
R1068 B.n315 B.n314 163.367
R1069 B.n315 B.n76 163.367
R1070 B.n319 B.n76 163.367
R1071 B.n320 B.n319 163.367
R1072 B.n321 B.n320 163.367
R1073 B.n321 B.n74 163.367
R1074 B.n325 B.n74 163.367
R1075 B.n326 B.n325 163.367
R1076 B.n327 B.n326 163.367
R1077 B.n327 B.n72 163.367
R1078 B.n331 B.n72 163.367
R1079 B.n332 B.n331 163.367
R1080 B.n333 B.n332 163.367
R1081 B.n333 B.n70 163.367
R1082 B.n337 B.n70 163.367
R1083 B.n338 B.n337 163.367
R1084 B.n339 B.n338 163.367
R1085 B.n339 B.n68 163.367
R1086 B.n343 B.n68 163.367
R1087 B.n344 B.n343 163.367
R1088 B.n345 B.n344 163.367
R1089 B.n345 B.n66 163.367
R1090 B.n349 B.n66 163.367
R1091 B.n350 B.n349 163.367
R1092 B.n351 B.n350 163.367
R1093 B.n351 B.n64 163.367
R1094 B.n355 B.n64 163.367
R1095 B.n356 B.n355 163.367
R1096 B.n357 B.n356 163.367
R1097 B.n357 B.n62 163.367
R1098 B.n361 B.n62 163.367
R1099 B.n362 B.n361 163.367
R1100 B.n363 B.n362 163.367
R1101 B.n363 B.n60 163.367
R1102 B.n367 B.n60 163.367
R1103 B.n368 B.n367 163.367
R1104 B.n369 B.n368 163.367
R1105 B.n369 B.n58 163.367
R1106 B.n373 B.n58 163.367
R1107 B.n484 B.n483 163.367
R1108 B.n483 B.n482 163.367
R1109 B.n482 B.n17 163.367
R1110 B.n478 B.n17 163.367
R1111 B.n478 B.n477 163.367
R1112 B.n477 B.n476 163.367
R1113 B.n476 B.n19 163.367
R1114 B.n472 B.n19 163.367
R1115 B.n472 B.n471 163.367
R1116 B.n471 B.n470 163.367
R1117 B.n470 B.n21 163.367
R1118 B.n466 B.n21 163.367
R1119 B.n466 B.n465 163.367
R1120 B.n465 B.n464 163.367
R1121 B.n464 B.n23 163.367
R1122 B.n460 B.n23 163.367
R1123 B.n460 B.n459 163.367
R1124 B.n459 B.n458 163.367
R1125 B.n458 B.n25 163.367
R1126 B.n454 B.n25 163.367
R1127 B.n454 B.n453 163.367
R1128 B.n453 B.n452 163.367
R1129 B.n452 B.n27 163.367
R1130 B.n448 B.n27 163.367
R1131 B.n448 B.n447 163.367
R1132 B.n447 B.n446 163.367
R1133 B.n446 B.n29 163.367
R1134 B.n442 B.n29 163.367
R1135 B.n442 B.n441 163.367
R1136 B.n441 B.n440 163.367
R1137 B.n440 B.n31 163.367
R1138 B.n435 B.n31 163.367
R1139 B.n435 B.n434 163.367
R1140 B.n434 B.n433 163.367
R1141 B.n433 B.n35 163.367
R1142 B.n429 B.n35 163.367
R1143 B.n429 B.n428 163.367
R1144 B.n428 B.n427 163.367
R1145 B.n427 B.n37 163.367
R1146 B.n423 B.n37 163.367
R1147 B.n423 B.n422 163.367
R1148 B.n422 B.n421 163.367
R1149 B.n421 B.n39 163.367
R1150 B.n417 B.n39 163.367
R1151 B.n417 B.n416 163.367
R1152 B.n416 B.n415 163.367
R1153 B.n415 B.n44 163.367
R1154 B.n411 B.n44 163.367
R1155 B.n411 B.n410 163.367
R1156 B.n410 B.n409 163.367
R1157 B.n409 B.n46 163.367
R1158 B.n405 B.n46 163.367
R1159 B.n405 B.n404 163.367
R1160 B.n404 B.n403 163.367
R1161 B.n403 B.n48 163.367
R1162 B.n399 B.n48 163.367
R1163 B.n399 B.n398 163.367
R1164 B.n398 B.n397 163.367
R1165 B.n397 B.n50 163.367
R1166 B.n393 B.n50 163.367
R1167 B.n393 B.n392 163.367
R1168 B.n392 B.n391 163.367
R1169 B.n391 B.n52 163.367
R1170 B.n387 B.n52 163.367
R1171 B.n387 B.n386 163.367
R1172 B.n386 B.n385 163.367
R1173 B.n385 B.n54 163.367
R1174 B.n381 B.n54 163.367
R1175 B.n381 B.n380 163.367
R1176 B.n380 B.n379 163.367
R1177 B.n379 B.n56 163.367
R1178 B.n375 B.n56 163.367
R1179 B.n375 B.n374 163.367
R1180 B.n103 B.n102 59.5399
R1181 B.n227 B.n110 59.5399
R1182 B.n437 B.n33 59.5399
R1183 B.n42 B.n41 59.5399
R1184 B.n102 B.n101 31.0308
R1185 B.n110 B.n109 31.0308
R1186 B.n33 B.n32 31.0308
R1187 B.n41 B.n40 31.0308
R1188 B.n372 B.n57 29.1907
R1189 B.n486 B.n485 29.1907
R1190 B.n292 B.n85 29.1907
R1191 B.n179 B.n178 29.1907
R1192 B B.n527 18.0485
R1193 B.n485 B.n16 10.6151
R1194 B.n481 B.n16 10.6151
R1195 B.n481 B.n480 10.6151
R1196 B.n480 B.n479 10.6151
R1197 B.n479 B.n18 10.6151
R1198 B.n475 B.n18 10.6151
R1199 B.n475 B.n474 10.6151
R1200 B.n474 B.n473 10.6151
R1201 B.n473 B.n20 10.6151
R1202 B.n469 B.n20 10.6151
R1203 B.n469 B.n468 10.6151
R1204 B.n468 B.n467 10.6151
R1205 B.n467 B.n22 10.6151
R1206 B.n463 B.n22 10.6151
R1207 B.n463 B.n462 10.6151
R1208 B.n462 B.n461 10.6151
R1209 B.n461 B.n24 10.6151
R1210 B.n457 B.n24 10.6151
R1211 B.n457 B.n456 10.6151
R1212 B.n456 B.n455 10.6151
R1213 B.n455 B.n26 10.6151
R1214 B.n451 B.n26 10.6151
R1215 B.n451 B.n450 10.6151
R1216 B.n450 B.n449 10.6151
R1217 B.n449 B.n28 10.6151
R1218 B.n445 B.n28 10.6151
R1219 B.n445 B.n444 10.6151
R1220 B.n444 B.n443 10.6151
R1221 B.n443 B.n30 10.6151
R1222 B.n439 B.n30 10.6151
R1223 B.n439 B.n438 10.6151
R1224 B.n436 B.n34 10.6151
R1225 B.n432 B.n34 10.6151
R1226 B.n432 B.n431 10.6151
R1227 B.n431 B.n430 10.6151
R1228 B.n430 B.n36 10.6151
R1229 B.n426 B.n36 10.6151
R1230 B.n426 B.n425 10.6151
R1231 B.n425 B.n424 10.6151
R1232 B.n424 B.n38 10.6151
R1233 B.n420 B.n419 10.6151
R1234 B.n419 B.n418 10.6151
R1235 B.n418 B.n43 10.6151
R1236 B.n414 B.n43 10.6151
R1237 B.n414 B.n413 10.6151
R1238 B.n413 B.n412 10.6151
R1239 B.n412 B.n45 10.6151
R1240 B.n408 B.n45 10.6151
R1241 B.n408 B.n407 10.6151
R1242 B.n407 B.n406 10.6151
R1243 B.n406 B.n47 10.6151
R1244 B.n402 B.n47 10.6151
R1245 B.n402 B.n401 10.6151
R1246 B.n401 B.n400 10.6151
R1247 B.n400 B.n49 10.6151
R1248 B.n396 B.n49 10.6151
R1249 B.n396 B.n395 10.6151
R1250 B.n395 B.n394 10.6151
R1251 B.n394 B.n51 10.6151
R1252 B.n390 B.n51 10.6151
R1253 B.n390 B.n389 10.6151
R1254 B.n389 B.n388 10.6151
R1255 B.n388 B.n53 10.6151
R1256 B.n384 B.n53 10.6151
R1257 B.n384 B.n383 10.6151
R1258 B.n383 B.n382 10.6151
R1259 B.n382 B.n55 10.6151
R1260 B.n378 B.n55 10.6151
R1261 B.n378 B.n377 10.6151
R1262 B.n377 B.n376 10.6151
R1263 B.n376 B.n57 10.6151
R1264 B.n293 B.n292 10.6151
R1265 B.n294 B.n293 10.6151
R1266 B.n294 B.n83 10.6151
R1267 B.n298 B.n83 10.6151
R1268 B.n299 B.n298 10.6151
R1269 B.n300 B.n299 10.6151
R1270 B.n300 B.n81 10.6151
R1271 B.n304 B.n81 10.6151
R1272 B.n305 B.n304 10.6151
R1273 B.n306 B.n305 10.6151
R1274 B.n306 B.n79 10.6151
R1275 B.n310 B.n79 10.6151
R1276 B.n311 B.n310 10.6151
R1277 B.n312 B.n311 10.6151
R1278 B.n312 B.n77 10.6151
R1279 B.n316 B.n77 10.6151
R1280 B.n317 B.n316 10.6151
R1281 B.n318 B.n317 10.6151
R1282 B.n318 B.n75 10.6151
R1283 B.n322 B.n75 10.6151
R1284 B.n323 B.n322 10.6151
R1285 B.n324 B.n323 10.6151
R1286 B.n324 B.n73 10.6151
R1287 B.n328 B.n73 10.6151
R1288 B.n329 B.n328 10.6151
R1289 B.n330 B.n329 10.6151
R1290 B.n330 B.n71 10.6151
R1291 B.n334 B.n71 10.6151
R1292 B.n335 B.n334 10.6151
R1293 B.n336 B.n335 10.6151
R1294 B.n336 B.n69 10.6151
R1295 B.n340 B.n69 10.6151
R1296 B.n341 B.n340 10.6151
R1297 B.n342 B.n341 10.6151
R1298 B.n342 B.n67 10.6151
R1299 B.n346 B.n67 10.6151
R1300 B.n347 B.n346 10.6151
R1301 B.n348 B.n347 10.6151
R1302 B.n348 B.n65 10.6151
R1303 B.n352 B.n65 10.6151
R1304 B.n353 B.n352 10.6151
R1305 B.n354 B.n353 10.6151
R1306 B.n354 B.n63 10.6151
R1307 B.n358 B.n63 10.6151
R1308 B.n359 B.n358 10.6151
R1309 B.n360 B.n359 10.6151
R1310 B.n360 B.n61 10.6151
R1311 B.n364 B.n61 10.6151
R1312 B.n365 B.n364 10.6151
R1313 B.n366 B.n365 10.6151
R1314 B.n366 B.n59 10.6151
R1315 B.n370 B.n59 10.6151
R1316 B.n371 B.n370 10.6151
R1317 B.n372 B.n371 10.6151
R1318 B.n180 B.n179 10.6151
R1319 B.n180 B.n125 10.6151
R1320 B.n184 B.n125 10.6151
R1321 B.n185 B.n184 10.6151
R1322 B.n186 B.n185 10.6151
R1323 B.n186 B.n123 10.6151
R1324 B.n190 B.n123 10.6151
R1325 B.n191 B.n190 10.6151
R1326 B.n192 B.n191 10.6151
R1327 B.n192 B.n121 10.6151
R1328 B.n196 B.n121 10.6151
R1329 B.n197 B.n196 10.6151
R1330 B.n198 B.n197 10.6151
R1331 B.n198 B.n119 10.6151
R1332 B.n202 B.n119 10.6151
R1333 B.n203 B.n202 10.6151
R1334 B.n204 B.n203 10.6151
R1335 B.n204 B.n117 10.6151
R1336 B.n208 B.n117 10.6151
R1337 B.n209 B.n208 10.6151
R1338 B.n210 B.n209 10.6151
R1339 B.n210 B.n115 10.6151
R1340 B.n214 B.n115 10.6151
R1341 B.n215 B.n214 10.6151
R1342 B.n216 B.n215 10.6151
R1343 B.n216 B.n113 10.6151
R1344 B.n220 B.n113 10.6151
R1345 B.n221 B.n220 10.6151
R1346 B.n222 B.n221 10.6151
R1347 B.n222 B.n111 10.6151
R1348 B.n226 B.n111 10.6151
R1349 B.n229 B.n228 10.6151
R1350 B.n229 B.n107 10.6151
R1351 B.n233 B.n107 10.6151
R1352 B.n234 B.n233 10.6151
R1353 B.n235 B.n234 10.6151
R1354 B.n235 B.n105 10.6151
R1355 B.n239 B.n105 10.6151
R1356 B.n240 B.n239 10.6151
R1357 B.n241 B.n240 10.6151
R1358 B.n245 B.n244 10.6151
R1359 B.n246 B.n245 10.6151
R1360 B.n246 B.n99 10.6151
R1361 B.n250 B.n99 10.6151
R1362 B.n251 B.n250 10.6151
R1363 B.n252 B.n251 10.6151
R1364 B.n252 B.n97 10.6151
R1365 B.n256 B.n97 10.6151
R1366 B.n257 B.n256 10.6151
R1367 B.n258 B.n257 10.6151
R1368 B.n258 B.n95 10.6151
R1369 B.n262 B.n95 10.6151
R1370 B.n263 B.n262 10.6151
R1371 B.n264 B.n263 10.6151
R1372 B.n264 B.n93 10.6151
R1373 B.n268 B.n93 10.6151
R1374 B.n269 B.n268 10.6151
R1375 B.n270 B.n269 10.6151
R1376 B.n270 B.n91 10.6151
R1377 B.n274 B.n91 10.6151
R1378 B.n275 B.n274 10.6151
R1379 B.n276 B.n275 10.6151
R1380 B.n276 B.n89 10.6151
R1381 B.n280 B.n89 10.6151
R1382 B.n281 B.n280 10.6151
R1383 B.n282 B.n281 10.6151
R1384 B.n282 B.n87 10.6151
R1385 B.n286 B.n87 10.6151
R1386 B.n287 B.n286 10.6151
R1387 B.n288 B.n287 10.6151
R1388 B.n288 B.n85 10.6151
R1389 B.n178 B.n127 10.6151
R1390 B.n174 B.n127 10.6151
R1391 B.n174 B.n173 10.6151
R1392 B.n173 B.n172 10.6151
R1393 B.n172 B.n129 10.6151
R1394 B.n168 B.n129 10.6151
R1395 B.n168 B.n167 10.6151
R1396 B.n167 B.n166 10.6151
R1397 B.n166 B.n131 10.6151
R1398 B.n162 B.n131 10.6151
R1399 B.n162 B.n161 10.6151
R1400 B.n161 B.n160 10.6151
R1401 B.n160 B.n133 10.6151
R1402 B.n156 B.n133 10.6151
R1403 B.n156 B.n155 10.6151
R1404 B.n155 B.n154 10.6151
R1405 B.n154 B.n135 10.6151
R1406 B.n150 B.n135 10.6151
R1407 B.n150 B.n149 10.6151
R1408 B.n149 B.n148 10.6151
R1409 B.n148 B.n137 10.6151
R1410 B.n144 B.n137 10.6151
R1411 B.n144 B.n143 10.6151
R1412 B.n143 B.n142 10.6151
R1413 B.n142 B.n139 10.6151
R1414 B.n139 B.n0 10.6151
R1415 B.n523 B.n1 10.6151
R1416 B.n523 B.n522 10.6151
R1417 B.n522 B.n521 10.6151
R1418 B.n521 B.n4 10.6151
R1419 B.n517 B.n4 10.6151
R1420 B.n517 B.n516 10.6151
R1421 B.n516 B.n515 10.6151
R1422 B.n515 B.n6 10.6151
R1423 B.n511 B.n6 10.6151
R1424 B.n511 B.n510 10.6151
R1425 B.n510 B.n509 10.6151
R1426 B.n509 B.n8 10.6151
R1427 B.n505 B.n8 10.6151
R1428 B.n505 B.n504 10.6151
R1429 B.n504 B.n503 10.6151
R1430 B.n503 B.n10 10.6151
R1431 B.n499 B.n10 10.6151
R1432 B.n499 B.n498 10.6151
R1433 B.n498 B.n497 10.6151
R1434 B.n497 B.n12 10.6151
R1435 B.n493 B.n12 10.6151
R1436 B.n493 B.n492 10.6151
R1437 B.n492 B.n491 10.6151
R1438 B.n491 B.n14 10.6151
R1439 B.n487 B.n14 10.6151
R1440 B.n487 B.n486 10.6151
R1441 B.n438 B.n437 9.36635
R1442 B.n420 B.n42 9.36635
R1443 B.n227 B.n226 9.36635
R1444 B.n244 B.n103 9.36635
R1445 B.n527 B.n0 2.81026
R1446 B.n527 B.n1 2.81026
R1447 B.n437 B.n436 1.24928
R1448 B.n42 B.n38 1.24928
R1449 B.n228 B.n227 1.24928
R1450 B.n241 B.n103 1.24928
C0 VTAIL VDD1 6.63866f
C1 VP w_n2250_n2712# 4.17045f
C2 VN B 0.844579f
C3 VDD2 w_n2250_n2712# 1.76574f
C4 VN VDD1 0.148439f
C5 VTAIL w_n2250_n2712# 2.40687f
C6 B VDD1 1.48193f
C7 VP VDD2 0.344857f
C8 VP VTAIL 4.14033f
C9 VTAIL VDD2 6.67971f
C10 VN w_n2250_n2712# 3.88326f
C11 B w_n2250_n2712# 6.91975f
C12 VDD1 w_n2250_n2712# 1.72358f
C13 VN VP 5.02887f
C14 VP B 1.31737f
C15 VN VDD2 4.14452f
C16 VP VDD1 4.33795f
C17 VN VTAIL 4.12597f
C18 B VDD2 1.52432f
C19 B VTAIL 2.41557f
C20 VDD1 VDD2 0.919051f
C21 VDD2 VSUBS 1.253017f
C22 VDD1 VSUBS 1.200491f
C23 VTAIL VSUBS 0.80727f
C24 VN VSUBS 4.54747f
C25 VP VSUBS 1.802902f
C26 B VSUBS 3.046108f
C27 w_n2250_n2712# VSUBS 75.573f
C28 B.n0 VSUBS 0.00469f
C29 B.n1 VSUBS 0.00469f
C30 B.n2 VSUBS 0.007417f
C31 B.n3 VSUBS 0.007417f
C32 B.n4 VSUBS 0.007417f
C33 B.n5 VSUBS 0.007417f
C34 B.n6 VSUBS 0.007417f
C35 B.n7 VSUBS 0.007417f
C36 B.n8 VSUBS 0.007417f
C37 B.n9 VSUBS 0.007417f
C38 B.n10 VSUBS 0.007417f
C39 B.n11 VSUBS 0.007417f
C40 B.n12 VSUBS 0.007417f
C41 B.n13 VSUBS 0.007417f
C42 B.n14 VSUBS 0.007417f
C43 B.n15 VSUBS 0.015534f
C44 B.n16 VSUBS 0.007417f
C45 B.n17 VSUBS 0.007417f
C46 B.n18 VSUBS 0.007417f
C47 B.n19 VSUBS 0.007417f
C48 B.n20 VSUBS 0.007417f
C49 B.n21 VSUBS 0.007417f
C50 B.n22 VSUBS 0.007417f
C51 B.n23 VSUBS 0.007417f
C52 B.n24 VSUBS 0.007417f
C53 B.n25 VSUBS 0.007417f
C54 B.n26 VSUBS 0.007417f
C55 B.n27 VSUBS 0.007417f
C56 B.n28 VSUBS 0.007417f
C57 B.n29 VSUBS 0.007417f
C58 B.n30 VSUBS 0.007417f
C59 B.n31 VSUBS 0.007417f
C60 B.t8 VSUBS 0.1495f
C61 B.t7 VSUBS 0.167249f
C62 B.t6 VSUBS 0.518058f
C63 B.n32 VSUBS 0.272179f
C64 B.n33 VSUBS 0.20946f
C65 B.n34 VSUBS 0.007417f
C66 B.n35 VSUBS 0.007417f
C67 B.n36 VSUBS 0.007417f
C68 B.n37 VSUBS 0.007417f
C69 B.n38 VSUBS 0.004145f
C70 B.n39 VSUBS 0.007417f
C71 B.t5 VSUBS 0.149503f
C72 B.t4 VSUBS 0.167252f
C73 B.t3 VSUBS 0.518058f
C74 B.n40 VSUBS 0.272176f
C75 B.n41 VSUBS 0.209458f
C76 B.n42 VSUBS 0.017185f
C77 B.n43 VSUBS 0.007417f
C78 B.n44 VSUBS 0.007417f
C79 B.n45 VSUBS 0.007417f
C80 B.n46 VSUBS 0.007417f
C81 B.n47 VSUBS 0.007417f
C82 B.n48 VSUBS 0.007417f
C83 B.n49 VSUBS 0.007417f
C84 B.n50 VSUBS 0.007417f
C85 B.n51 VSUBS 0.007417f
C86 B.n52 VSUBS 0.007417f
C87 B.n53 VSUBS 0.007417f
C88 B.n54 VSUBS 0.007417f
C89 B.n55 VSUBS 0.007417f
C90 B.n56 VSUBS 0.007417f
C91 B.n57 VSUBS 0.015773f
C92 B.n58 VSUBS 0.007417f
C93 B.n59 VSUBS 0.007417f
C94 B.n60 VSUBS 0.007417f
C95 B.n61 VSUBS 0.007417f
C96 B.n62 VSUBS 0.007417f
C97 B.n63 VSUBS 0.007417f
C98 B.n64 VSUBS 0.007417f
C99 B.n65 VSUBS 0.007417f
C100 B.n66 VSUBS 0.007417f
C101 B.n67 VSUBS 0.007417f
C102 B.n68 VSUBS 0.007417f
C103 B.n69 VSUBS 0.007417f
C104 B.n70 VSUBS 0.007417f
C105 B.n71 VSUBS 0.007417f
C106 B.n72 VSUBS 0.007417f
C107 B.n73 VSUBS 0.007417f
C108 B.n74 VSUBS 0.007417f
C109 B.n75 VSUBS 0.007417f
C110 B.n76 VSUBS 0.007417f
C111 B.n77 VSUBS 0.007417f
C112 B.n78 VSUBS 0.007417f
C113 B.n79 VSUBS 0.007417f
C114 B.n80 VSUBS 0.007417f
C115 B.n81 VSUBS 0.007417f
C116 B.n82 VSUBS 0.007417f
C117 B.n83 VSUBS 0.007417f
C118 B.n84 VSUBS 0.007417f
C119 B.n85 VSUBS 0.016754f
C120 B.n86 VSUBS 0.007417f
C121 B.n87 VSUBS 0.007417f
C122 B.n88 VSUBS 0.007417f
C123 B.n89 VSUBS 0.007417f
C124 B.n90 VSUBS 0.007417f
C125 B.n91 VSUBS 0.007417f
C126 B.n92 VSUBS 0.007417f
C127 B.n93 VSUBS 0.007417f
C128 B.n94 VSUBS 0.007417f
C129 B.n95 VSUBS 0.007417f
C130 B.n96 VSUBS 0.007417f
C131 B.n97 VSUBS 0.007417f
C132 B.n98 VSUBS 0.007417f
C133 B.n99 VSUBS 0.007417f
C134 B.n100 VSUBS 0.007417f
C135 B.t1 VSUBS 0.149503f
C136 B.t2 VSUBS 0.167252f
C137 B.t0 VSUBS 0.518058f
C138 B.n101 VSUBS 0.272176f
C139 B.n102 VSUBS 0.209458f
C140 B.n103 VSUBS 0.017185f
C141 B.n104 VSUBS 0.007417f
C142 B.n105 VSUBS 0.007417f
C143 B.n106 VSUBS 0.007417f
C144 B.n107 VSUBS 0.007417f
C145 B.n108 VSUBS 0.007417f
C146 B.t10 VSUBS 0.1495f
C147 B.t11 VSUBS 0.167249f
C148 B.t9 VSUBS 0.518058f
C149 B.n109 VSUBS 0.272179f
C150 B.n110 VSUBS 0.20946f
C151 B.n111 VSUBS 0.007417f
C152 B.n112 VSUBS 0.007417f
C153 B.n113 VSUBS 0.007417f
C154 B.n114 VSUBS 0.007417f
C155 B.n115 VSUBS 0.007417f
C156 B.n116 VSUBS 0.007417f
C157 B.n117 VSUBS 0.007417f
C158 B.n118 VSUBS 0.007417f
C159 B.n119 VSUBS 0.007417f
C160 B.n120 VSUBS 0.007417f
C161 B.n121 VSUBS 0.007417f
C162 B.n122 VSUBS 0.007417f
C163 B.n123 VSUBS 0.007417f
C164 B.n124 VSUBS 0.007417f
C165 B.n125 VSUBS 0.007417f
C166 B.n126 VSUBS 0.016754f
C167 B.n127 VSUBS 0.007417f
C168 B.n128 VSUBS 0.007417f
C169 B.n129 VSUBS 0.007417f
C170 B.n130 VSUBS 0.007417f
C171 B.n131 VSUBS 0.007417f
C172 B.n132 VSUBS 0.007417f
C173 B.n133 VSUBS 0.007417f
C174 B.n134 VSUBS 0.007417f
C175 B.n135 VSUBS 0.007417f
C176 B.n136 VSUBS 0.007417f
C177 B.n137 VSUBS 0.007417f
C178 B.n138 VSUBS 0.007417f
C179 B.n139 VSUBS 0.007417f
C180 B.n140 VSUBS 0.007417f
C181 B.n141 VSUBS 0.007417f
C182 B.n142 VSUBS 0.007417f
C183 B.n143 VSUBS 0.007417f
C184 B.n144 VSUBS 0.007417f
C185 B.n145 VSUBS 0.007417f
C186 B.n146 VSUBS 0.007417f
C187 B.n147 VSUBS 0.007417f
C188 B.n148 VSUBS 0.007417f
C189 B.n149 VSUBS 0.007417f
C190 B.n150 VSUBS 0.007417f
C191 B.n151 VSUBS 0.007417f
C192 B.n152 VSUBS 0.007417f
C193 B.n153 VSUBS 0.007417f
C194 B.n154 VSUBS 0.007417f
C195 B.n155 VSUBS 0.007417f
C196 B.n156 VSUBS 0.007417f
C197 B.n157 VSUBS 0.007417f
C198 B.n158 VSUBS 0.007417f
C199 B.n159 VSUBS 0.007417f
C200 B.n160 VSUBS 0.007417f
C201 B.n161 VSUBS 0.007417f
C202 B.n162 VSUBS 0.007417f
C203 B.n163 VSUBS 0.007417f
C204 B.n164 VSUBS 0.007417f
C205 B.n165 VSUBS 0.007417f
C206 B.n166 VSUBS 0.007417f
C207 B.n167 VSUBS 0.007417f
C208 B.n168 VSUBS 0.007417f
C209 B.n169 VSUBS 0.007417f
C210 B.n170 VSUBS 0.007417f
C211 B.n171 VSUBS 0.007417f
C212 B.n172 VSUBS 0.007417f
C213 B.n173 VSUBS 0.007417f
C214 B.n174 VSUBS 0.007417f
C215 B.n175 VSUBS 0.007417f
C216 B.n176 VSUBS 0.007417f
C217 B.n177 VSUBS 0.015534f
C218 B.n178 VSUBS 0.015534f
C219 B.n179 VSUBS 0.016754f
C220 B.n180 VSUBS 0.007417f
C221 B.n181 VSUBS 0.007417f
C222 B.n182 VSUBS 0.007417f
C223 B.n183 VSUBS 0.007417f
C224 B.n184 VSUBS 0.007417f
C225 B.n185 VSUBS 0.007417f
C226 B.n186 VSUBS 0.007417f
C227 B.n187 VSUBS 0.007417f
C228 B.n188 VSUBS 0.007417f
C229 B.n189 VSUBS 0.007417f
C230 B.n190 VSUBS 0.007417f
C231 B.n191 VSUBS 0.007417f
C232 B.n192 VSUBS 0.007417f
C233 B.n193 VSUBS 0.007417f
C234 B.n194 VSUBS 0.007417f
C235 B.n195 VSUBS 0.007417f
C236 B.n196 VSUBS 0.007417f
C237 B.n197 VSUBS 0.007417f
C238 B.n198 VSUBS 0.007417f
C239 B.n199 VSUBS 0.007417f
C240 B.n200 VSUBS 0.007417f
C241 B.n201 VSUBS 0.007417f
C242 B.n202 VSUBS 0.007417f
C243 B.n203 VSUBS 0.007417f
C244 B.n204 VSUBS 0.007417f
C245 B.n205 VSUBS 0.007417f
C246 B.n206 VSUBS 0.007417f
C247 B.n207 VSUBS 0.007417f
C248 B.n208 VSUBS 0.007417f
C249 B.n209 VSUBS 0.007417f
C250 B.n210 VSUBS 0.007417f
C251 B.n211 VSUBS 0.007417f
C252 B.n212 VSUBS 0.007417f
C253 B.n213 VSUBS 0.007417f
C254 B.n214 VSUBS 0.007417f
C255 B.n215 VSUBS 0.007417f
C256 B.n216 VSUBS 0.007417f
C257 B.n217 VSUBS 0.007417f
C258 B.n218 VSUBS 0.007417f
C259 B.n219 VSUBS 0.007417f
C260 B.n220 VSUBS 0.007417f
C261 B.n221 VSUBS 0.007417f
C262 B.n222 VSUBS 0.007417f
C263 B.n223 VSUBS 0.007417f
C264 B.n224 VSUBS 0.007417f
C265 B.n225 VSUBS 0.007417f
C266 B.n226 VSUBS 0.006981f
C267 B.n227 VSUBS 0.017185f
C268 B.n228 VSUBS 0.004145f
C269 B.n229 VSUBS 0.007417f
C270 B.n230 VSUBS 0.007417f
C271 B.n231 VSUBS 0.007417f
C272 B.n232 VSUBS 0.007417f
C273 B.n233 VSUBS 0.007417f
C274 B.n234 VSUBS 0.007417f
C275 B.n235 VSUBS 0.007417f
C276 B.n236 VSUBS 0.007417f
C277 B.n237 VSUBS 0.007417f
C278 B.n238 VSUBS 0.007417f
C279 B.n239 VSUBS 0.007417f
C280 B.n240 VSUBS 0.007417f
C281 B.n241 VSUBS 0.004145f
C282 B.n242 VSUBS 0.007417f
C283 B.n243 VSUBS 0.007417f
C284 B.n244 VSUBS 0.006981f
C285 B.n245 VSUBS 0.007417f
C286 B.n246 VSUBS 0.007417f
C287 B.n247 VSUBS 0.007417f
C288 B.n248 VSUBS 0.007417f
C289 B.n249 VSUBS 0.007417f
C290 B.n250 VSUBS 0.007417f
C291 B.n251 VSUBS 0.007417f
C292 B.n252 VSUBS 0.007417f
C293 B.n253 VSUBS 0.007417f
C294 B.n254 VSUBS 0.007417f
C295 B.n255 VSUBS 0.007417f
C296 B.n256 VSUBS 0.007417f
C297 B.n257 VSUBS 0.007417f
C298 B.n258 VSUBS 0.007417f
C299 B.n259 VSUBS 0.007417f
C300 B.n260 VSUBS 0.007417f
C301 B.n261 VSUBS 0.007417f
C302 B.n262 VSUBS 0.007417f
C303 B.n263 VSUBS 0.007417f
C304 B.n264 VSUBS 0.007417f
C305 B.n265 VSUBS 0.007417f
C306 B.n266 VSUBS 0.007417f
C307 B.n267 VSUBS 0.007417f
C308 B.n268 VSUBS 0.007417f
C309 B.n269 VSUBS 0.007417f
C310 B.n270 VSUBS 0.007417f
C311 B.n271 VSUBS 0.007417f
C312 B.n272 VSUBS 0.007417f
C313 B.n273 VSUBS 0.007417f
C314 B.n274 VSUBS 0.007417f
C315 B.n275 VSUBS 0.007417f
C316 B.n276 VSUBS 0.007417f
C317 B.n277 VSUBS 0.007417f
C318 B.n278 VSUBS 0.007417f
C319 B.n279 VSUBS 0.007417f
C320 B.n280 VSUBS 0.007417f
C321 B.n281 VSUBS 0.007417f
C322 B.n282 VSUBS 0.007417f
C323 B.n283 VSUBS 0.007417f
C324 B.n284 VSUBS 0.007417f
C325 B.n285 VSUBS 0.007417f
C326 B.n286 VSUBS 0.007417f
C327 B.n287 VSUBS 0.007417f
C328 B.n288 VSUBS 0.007417f
C329 B.n289 VSUBS 0.007417f
C330 B.n290 VSUBS 0.016754f
C331 B.n291 VSUBS 0.015534f
C332 B.n292 VSUBS 0.015534f
C333 B.n293 VSUBS 0.007417f
C334 B.n294 VSUBS 0.007417f
C335 B.n295 VSUBS 0.007417f
C336 B.n296 VSUBS 0.007417f
C337 B.n297 VSUBS 0.007417f
C338 B.n298 VSUBS 0.007417f
C339 B.n299 VSUBS 0.007417f
C340 B.n300 VSUBS 0.007417f
C341 B.n301 VSUBS 0.007417f
C342 B.n302 VSUBS 0.007417f
C343 B.n303 VSUBS 0.007417f
C344 B.n304 VSUBS 0.007417f
C345 B.n305 VSUBS 0.007417f
C346 B.n306 VSUBS 0.007417f
C347 B.n307 VSUBS 0.007417f
C348 B.n308 VSUBS 0.007417f
C349 B.n309 VSUBS 0.007417f
C350 B.n310 VSUBS 0.007417f
C351 B.n311 VSUBS 0.007417f
C352 B.n312 VSUBS 0.007417f
C353 B.n313 VSUBS 0.007417f
C354 B.n314 VSUBS 0.007417f
C355 B.n315 VSUBS 0.007417f
C356 B.n316 VSUBS 0.007417f
C357 B.n317 VSUBS 0.007417f
C358 B.n318 VSUBS 0.007417f
C359 B.n319 VSUBS 0.007417f
C360 B.n320 VSUBS 0.007417f
C361 B.n321 VSUBS 0.007417f
C362 B.n322 VSUBS 0.007417f
C363 B.n323 VSUBS 0.007417f
C364 B.n324 VSUBS 0.007417f
C365 B.n325 VSUBS 0.007417f
C366 B.n326 VSUBS 0.007417f
C367 B.n327 VSUBS 0.007417f
C368 B.n328 VSUBS 0.007417f
C369 B.n329 VSUBS 0.007417f
C370 B.n330 VSUBS 0.007417f
C371 B.n331 VSUBS 0.007417f
C372 B.n332 VSUBS 0.007417f
C373 B.n333 VSUBS 0.007417f
C374 B.n334 VSUBS 0.007417f
C375 B.n335 VSUBS 0.007417f
C376 B.n336 VSUBS 0.007417f
C377 B.n337 VSUBS 0.007417f
C378 B.n338 VSUBS 0.007417f
C379 B.n339 VSUBS 0.007417f
C380 B.n340 VSUBS 0.007417f
C381 B.n341 VSUBS 0.007417f
C382 B.n342 VSUBS 0.007417f
C383 B.n343 VSUBS 0.007417f
C384 B.n344 VSUBS 0.007417f
C385 B.n345 VSUBS 0.007417f
C386 B.n346 VSUBS 0.007417f
C387 B.n347 VSUBS 0.007417f
C388 B.n348 VSUBS 0.007417f
C389 B.n349 VSUBS 0.007417f
C390 B.n350 VSUBS 0.007417f
C391 B.n351 VSUBS 0.007417f
C392 B.n352 VSUBS 0.007417f
C393 B.n353 VSUBS 0.007417f
C394 B.n354 VSUBS 0.007417f
C395 B.n355 VSUBS 0.007417f
C396 B.n356 VSUBS 0.007417f
C397 B.n357 VSUBS 0.007417f
C398 B.n358 VSUBS 0.007417f
C399 B.n359 VSUBS 0.007417f
C400 B.n360 VSUBS 0.007417f
C401 B.n361 VSUBS 0.007417f
C402 B.n362 VSUBS 0.007417f
C403 B.n363 VSUBS 0.007417f
C404 B.n364 VSUBS 0.007417f
C405 B.n365 VSUBS 0.007417f
C406 B.n366 VSUBS 0.007417f
C407 B.n367 VSUBS 0.007417f
C408 B.n368 VSUBS 0.007417f
C409 B.n369 VSUBS 0.007417f
C410 B.n370 VSUBS 0.007417f
C411 B.n371 VSUBS 0.007417f
C412 B.n372 VSUBS 0.016515f
C413 B.n373 VSUBS 0.015534f
C414 B.n374 VSUBS 0.016754f
C415 B.n375 VSUBS 0.007417f
C416 B.n376 VSUBS 0.007417f
C417 B.n377 VSUBS 0.007417f
C418 B.n378 VSUBS 0.007417f
C419 B.n379 VSUBS 0.007417f
C420 B.n380 VSUBS 0.007417f
C421 B.n381 VSUBS 0.007417f
C422 B.n382 VSUBS 0.007417f
C423 B.n383 VSUBS 0.007417f
C424 B.n384 VSUBS 0.007417f
C425 B.n385 VSUBS 0.007417f
C426 B.n386 VSUBS 0.007417f
C427 B.n387 VSUBS 0.007417f
C428 B.n388 VSUBS 0.007417f
C429 B.n389 VSUBS 0.007417f
C430 B.n390 VSUBS 0.007417f
C431 B.n391 VSUBS 0.007417f
C432 B.n392 VSUBS 0.007417f
C433 B.n393 VSUBS 0.007417f
C434 B.n394 VSUBS 0.007417f
C435 B.n395 VSUBS 0.007417f
C436 B.n396 VSUBS 0.007417f
C437 B.n397 VSUBS 0.007417f
C438 B.n398 VSUBS 0.007417f
C439 B.n399 VSUBS 0.007417f
C440 B.n400 VSUBS 0.007417f
C441 B.n401 VSUBS 0.007417f
C442 B.n402 VSUBS 0.007417f
C443 B.n403 VSUBS 0.007417f
C444 B.n404 VSUBS 0.007417f
C445 B.n405 VSUBS 0.007417f
C446 B.n406 VSUBS 0.007417f
C447 B.n407 VSUBS 0.007417f
C448 B.n408 VSUBS 0.007417f
C449 B.n409 VSUBS 0.007417f
C450 B.n410 VSUBS 0.007417f
C451 B.n411 VSUBS 0.007417f
C452 B.n412 VSUBS 0.007417f
C453 B.n413 VSUBS 0.007417f
C454 B.n414 VSUBS 0.007417f
C455 B.n415 VSUBS 0.007417f
C456 B.n416 VSUBS 0.007417f
C457 B.n417 VSUBS 0.007417f
C458 B.n418 VSUBS 0.007417f
C459 B.n419 VSUBS 0.007417f
C460 B.n420 VSUBS 0.006981f
C461 B.n421 VSUBS 0.007417f
C462 B.n422 VSUBS 0.007417f
C463 B.n423 VSUBS 0.007417f
C464 B.n424 VSUBS 0.007417f
C465 B.n425 VSUBS 0.007417f
C466 B.n426 VSUBS 0.007417f
C467 B.n427 VSUBS 0.007417f
C468 B.n428 VSUBS 0.007417f
C469 B.n429 VSUBS 0.007417f
C470 B.n430 VSUBS 0.007417f
C471 B.n431 VSUBS 0.007417f
C472 B.n432 VSUBS 0.007417f
C473 B.n433 VSUBS 0.007417f
C474 B.n434 VSUBS 0.007417f
C475 B.n435 VSUBS 0.007417f
C476 B.n436 VSUBS 0.004145f
C477 B.n437 VSUBS 0.017185f
C478 B.n438 VSUBS 0.006981f
C479 B.n439 VSUBS 0.007417f
C480 B.n440 VSUBS 0.007417f
C481 B.n441 VSUBS 0.007417f
C482 B.n442 VSUBS 0.007417f
C483 B.n443 VSUBS 0.007417f
C484 B.n444 VSUBS 0.007417f
C485 B.n445 VSUBS 0.007417f
C486 B.n446 VSUBS 0.007417f
C487 B.n447 VSUBS 0.007417f
C488 B.n448 VSUBS 0.007417f
C489 B.n449 VSUBS 0.007417f
C490 B.n450 VSUBS 0.007417f
C491 B.n451 VSUBS 0.007417f
C492 B.n452 VSUBS 0.007417f
C493 B.n453 VSUBS 0.007417f
C494 B.n454 VSUBS 0.007417f
C495 B.n455 VSUBS 0.007417f
C496 B.n456 VSUBS 0.007417f
C497 B.n457 VSUBS 0.007417f
C498 B.n458 VSUBS 0.007417f
C499 B.n459 VSUBS 0.007417f
C500 B.n460 VSUBS 0.007417f
C501 B.n461 VSUBS 0.007417f
C502 B.n462 VSUBS 0.007417f
C503 B.n463 VSUBS 0.007417f
C504 B.n464 VSUBS 0.007417f
C505 B.n465 VSUBS 0.007417f
C506 B.n466 VSUBS 0.007417f
C507 B.n467 VSUBS 0.007417f
C508 B.n468 VSUBS 0.007417f
C509 B.n469 VSUBS 0.007417f
C510 B.n470 VSUBS 0.007417f
C511 B.n471 VSUBS 0.007417f
C512 B.n472 VSUBS 0.007417f
C513 B.n473 VSUBS 0.007417f
C514 B.n474 VSUBS 0.007417f
C515 B.n475 VSUBS 0.007417f
C516 B.n476 VSUBS 0.007417f
C517 B.n477 VSUBS 0.007417f
C518 B.n478 VSUBS 0.007417f
C519 B.n479 VSUBS 0.007417f
C520 B.n480 VSUBS 0.007417f
C521 B.n481 VSUBS 0.007417f
C522 B.n482 VSUBS 0.007417f
C523 B.n483 VSUBS 0.007417f
C524 B.n484 VSUBS 0.016754f
C525 B.n485 VSUBS 0.016754f
C526 B.n486 VSUBS 0.015534f
C527 B.n487 VSUBS 0.007417f
C528 B.n488 VSUBS 0.007417f
C529 B.n489 VSUBS 0.007417f
C530 B.n490 VSUBS 0.007417f
C531 B.n491 VSUBS 0.007417f
C532 B.n492 VSUBS 0.007417f
C533 B.n493 VSUBS 0.007417f
C534 B.n494 VSUBS 0.007417f
C535 B.n495 VSUBS 0.007417f
C536 B.n496 VSUBS 0.007417f
C537 B.n497 VSUBS 0.007417f
C538 B.n498 VSUBS 0.007417f
C539 B.n499 VSUBS 0.007417f
C540 B.n500 VSUBS 0.007417f
C541 B.n501 VSUBS 0.007417f
C542 B.n502 VSUBS 0.007417f
C543 B.n503 VSUBS 0.007417f
C544 B.n504 VSUBS 0.007417f
C545 B.n505 VSUBS 0.007417f
C546 B.n506 VSUBS 0.007417f
C547 B.n507 VSUBS 0.007417f
C548 B.n508 VSUBS 0.007417f
C549 B.n509 VSUBS 0.007417f
C550 B.n510 VSUBS 0.007417f
C551 B.n511 VSUBS 0.007417f
C552 B.n512 VSUBS 0.007417f
C553 B.n513 VSUBS 0.007417f
C554 B.n514 VSUBS 0.007417f
C555 B.n515 VSUBS 0.007417f
C556 B.n516 VSUBS 0.007417f
C557 B.n517 VSUBS 0.007417f
C558 B.n518 VSUBS 0.007417f
C559 B.n519 VSUBS 0.007417f
C560 B.n520 VSUBS 0.007417f
C561 B.n521 VSUBS 0.007417f
C562 B.n522 VSUBS 0.007417f
C563 B.n523 VSUBS 0.007417f
C564 B.n524 VSUBS 0.007417f
C565 B.n525 VSUBS 0.007417f
C566 B.n526 VSUBS 0.007417f
C567 B.n527 VSUBS 0.016796f
C568 VDD2.n0 VSUBS 0.024103f
C569 VDD2.n1 VSUBS 0.022019f
C570 VDD2.n2 VSUBS 0.011832f
C571 VDD2.n3 VSUBS 0.027967f
C572 VDD2.n4 VSUBS 0.012528f
C573 VDD2.n5 VSUBS 0.022019f
C574 VDD2.n6 VSUBS 0.011832f
C575 VDD2.n7 VSUBS 0.027967f
C576 VDD2.n8 VSUBS 0.012528f
C577 VDD2.n9 VSUBS 0.022019f
C578 VDD2.n10 VSUBS 0.011832f
C579 VDD2.n11 VSUBS 0.027967f
C580 VDD2.n12 VSUBS 0.012528f
C581 VDD2.n13 VSUBS 0.14082f
C582 VDD2.t0 VSUBS 0.060094f
C583 VDD2.n14 VSUBS 0.020975f
C584 VDD2.n15 VSUBS 0.021038f
C585 VDD2.n16 VSUBS 0.011832f
C586 VDD2.n17 VSUBS 0.765296f
C587 VDD2.n18 VSUBS 0.022019f
C588 VDD2.n19 VSUBS 0.011832f
C589 VDD2.n20 VSUBS 0.012528f
C590 VDD2.n21 VSUBS 0.027967f
C591 VDD2.n22 VSUBS 0.027967f
C592 VDD2.n23 VSUBS 0.012528f
C593 VDD2.n24 VSUBS 0.011832f
C594 VDD2.n25 VSUBS 0.022019f
C595 VDD2.n26 VSUBS 0.022019f
C596 VDD2.n27 VSUBS 0.011832f
C597 VDD2.n28 VSUBS 0.012528f
C598 VDD2.n29 VSUBS 0.027967f
C599 VDD2.n30 VSUBS 0.027967f
C600 VDD2.n31 VSUBS 0.027967f
C601 VDD2.n32 VSUBS 0.012528f
C602 VDD2.n33 VSUBS 0.011832f
C603 VDD2.n34 VSUBS 0.022019f
C604 VDD2.n35 VSUBS 0.022019f
C605 VDD2.n36 VSUBS 0.011832f
C606 VDD2.n37 VSUBS 0.01218f
C607 VDD2.n38 VSUBS 0.01218f
C608 VDD2.n39 VSUBS 0.027967f
C609 VDD2.n40 VSUBS 0.067392f
C610 VDD2.n41 VSUBS 0.012528f
C611 VDD2.n42 VSUBS 0.011832f
C612 VDD2.n43 VSUBS 0.056913f
C613 VDD2.n44 VSUBS 0.051327f
C614 VDD2.t4 VSUBS 0.151732f
C615 VDD2.t2 VSUBS 0.151732f
C616 VDD2.n45 VSUBS 1.12443f
C617 VDD2.n46 VSUBS 1.87516f
C618 VDD2.n47 VSUBS 0.024103f
C619 VDD2.n48 VSUBS 0.022019f
C620 VDD2.n49 VSUBS 0.011832f
C621 VDD2.n50 VSUBS 0.027967f
C622 VDD2.n51 VSUBS 0.012528f
C623 VDD2.n52 VSUBS 0.022019f
C624 VDD2.n53 VSUBS 0.011832f
C625 VDD2.n54 VSUBS 0.027967f
C626 VDD2.n55 VSUBS 0.027967f
C627 VDD2.n56 VSUBS 0.012528f
C628 VDD2.n57 VSUBS 0.022019f
C629 VDD2.n58 VSUBS 0.011832f
C630 VDD2.n59 VSUBS 0.027967f
C631 VDD2.n60 VSUBS 0.012528f
C632 VDD2.n61 VSUBS 0.14082f
C633 VDD2.t1 VSUBS 0.060094f
C634 VDD2.n62 VSUBS 0.020975f
C635 VDD2.n63 VSUBS 0.021038f
C636 VDD2.n64 VSUBS 0.011832f
C637 VDD2.n65 VSUBS 0.765296f
C638 VDD2.n66 VSUBS 0.022019f
C639 VDD2.n67 VSUBS 0.011832f
C640 VDD2.n68 VSUBS 0.012528f
C641 VDD2.n69 VSUBS 0.027967f
C642 VDD2.n70 VSUBS 0.027967f
C643 VDD2.n71 VSUBS 0.012528f
C644 VDD2.n72 VSUBS 0.011832f
C645 VDD2.n73 VSUBS 0.022019f
C646 VDD2.n74 VSUBS 0.022019f
C647 VDD2.n75 VSUBS 0.011832f
C648 VDD2.n76 VSUBS 0.012528f
C649 VDD2.n77 VSUBS 0.027967f
C650 VDD2.n78 VSUBS 0.027967f
C651 VDD2.n79 VSUBS 0.012528f
C652 VDD2.n80 VSUBS 0.011832f
C653 VDD2.n81 VSUBS 0.022019f
C654 VDD2.n82 VSUBS 0.022019f
C655 VDD2.n83 VSUBS 0.011832f
C656 VDD2.n84 VSUBS 0.01218f
C657 VDD2.n85 VSUBS 0.01218f
C658 VDD2.n86 VSUBS 0.027967f
C659 VDD2.n87 VSUBS 0.067392f
C660 VDD2.n88 VSUBS 0.012528f
C661 VDD2.n89 VSUBS 0.011832f
C662 VDD2.n90 VSUBS 0.056913f
C663 VDD2.n91 VSUBS 0.049215f
C664 VDD2.n92 VSUBS 1.71342f
C665 VDD2.t5 VSUBS 0.151732f
C666 VDD2.t3 VSUBS 0.151732f
C667 VDD2.n93 VSUBS 1.1244f
C668 VN.n0 VSUBS 0.062114f
C669 VN.t1 VSUBS 1.38947f
C670 VN.n1 VSUBS 0.585451f
C671 VN.t5 VSUBS 1.53621f
C672 VN.n2 VSUBS 0.606003f
C673 VN.n3 VSUBS 0.244036f
C674 VN.n4 VSUBS 0.072991f
C675 VN.n5 VSUBS 0.029786f
C676 VN.t3 VSUBS 1.48059f
C677 VN.n6 VSUBS 0.617489f
C678 VN.n7 VSUBS 0.043595f
C679 VN.n8 VSUBS 0.062114f
C680 VN.t0 VSUBS 1.38947f
C681 VN.n9 VSUBS 0.585451f
C682 VN.t2 VSUBS 1.53621f
C683 VN.n10 VSUBS 0.606003f
C684 VN.n11 VSUBS 0.244036f
C685 VN.n12 VSUBS 0.072991f
C686 VN.n13 VSUBS 0.029786f
C687 VN.t4 VSUBS 1.48059f
C688 VN.n14 VSUBS 0.617489f
C689 VN.n15 VSUBS 1.89908f
C690 VTAIL.t3 VSUBS 0.203009f
C691 VTAIL.t10 VSUBS 0.203009f
C692 VTAIL.n0 VSUBS 1.37883f
C693 VTAIL.n1 VSUBS 0.73608f
C694 VTAIL.n2 VSUBS 0.032248f
C695 VTAIL.n3 VSUBS 0.029461f
C696 VTAIL.n4 VSUBS 0.015831f
C697 VTAIL.n5 VSUBS 0.037419f
C698 VTAIL.n6 VSUBS 0.016762f
C699 VTAIL.n7 VSUBS 0.029461f
C700 VTAIL.n8 VSUBS 0.015831f
C701 VTAIL.n9 VSUBS 0.037419f
C702 VTAIL.n10 VSUBS 0.016762f
C703 VTAIL.n11 VSUBS 0.029461f
C704 VTAIL.n12 VSUBS 0.015831f
C705 VTAIL.n13 VSUBS 0.037419f
C706 VTAIL.n14 VSUBS 0.016762f
C707 VTAIL.n15 VSUBS 0.18841f
C708 VTAIL.t8 VSUBS 0.080402f
C709 VTAIL.n16 VSUBS 0.028064f
C710 VTAIL.n17 VSUBS 0.028148f
C711 VTAIL.n18 VSUBS 0.015831f
C712 VTAIL.n19 VSUBS 1.02393f
C713 VTAIL.n20 VSUBS 0.029461f
C714 VTAIL.n21 VSUBS 0.015831f
C715 VTAIL.n22 VSUBS 0.016762f
C716 VTAIL.n23 VSUBS 0.037419f
C717 VTAIL.n24 VSUBS 0.037419f
C718 VTAIL.n25 VSUBS 0.016762f
C719 VTAIL.n26 VSUBS 0.015831f
C720 VTAIL.n27 VSUBS 0.029461f
C721 VTAIL.n28 VSUBS 0.029461f
C722 VTAIL.n29 VSUBS 0.015831f
C723 VTAIL.n30 VSUBS 0.016762f
C724 VTAIL.n31 VSUBS 0.037419f
C725 VTAIL.n32 VSUBS 0.037419f
C726 VTAIL.n33 VSUBS 0.037419f
C727 VTAIL.n34 VSUBS 0.016762f
C728 VTAIL.n35 VSUBS 0.015831f
C729 VTAIL.n36 VSUBS 0.029461f
C730 VTAIL.n37 VSUBS 0.029461f
C731 VTAIL.n38 VSUBS 0.015831f
C732 VTAIL.n39 VSUBS 0.016297f
C733 VTAIL.n40 VSUBS 0.016297f
C734 VTAIL.n41 VSUBS 0.037419f
C735 VTAIL.n42 VSUBS 0.090167f
C736 VTAIL.n43 VSUBS 0.016762f
C737 VTAIL.n44 VSUBS 0.015831f
C738 VTAIL.n45 VSUBS 0.076147f
C739 VTAIL.n46 VSUBS 0.045561f
C740 VTAIL.n47 VSUBS 0.270723f
C741 VTAIL.t4 VSUBS 0.203009f
C742 VTAIL.t6 VSUBS 0.203009f
C743 VTAIL.n48 VSUBS 1.37883f
C744 VTAIL.n49 VSUBS 2.09436f
C745 VTAIL.t1 VSUBS 0.203009f
C746 VTAIL.t2 VSUBS 0.203009f
C747 VTAIL.n50 VSUBS 1.37884f
C748 VTAIL.n51 VSUBS 2.09435f
C749 VTAIL.n52 VSUBS 0.032248f
C750 VTAIL.n53 VSUBS 0.029461f
C751 VTAIL.n54 VSUBS 0.015831f
C752 VTAIL.n55 VSUBS 0.037419f
C753 VTAIL.n56 VSUBS 0.016762f
C754 VTAIL.n57 VSUBS 0.029461f
C755 VTAIL.n58 VSUBS 0.015831f
C756 VTAIL.n59 VSUBS 0.037419f
C757 VTAIL.n60 VSUBS 0.037419f
C758 VTAIL.n61 VSUBS 0.016762f
C759 VTAIL.n62 VSUBS 0.029461f
C760 VTAIL.n63 VSUBS 0.015831f
C761 VTAIL.n64 VSUBS 0.037419f
C762 VTAIL.n65 VSUBS 0.016762f
C763 VTAIL.n66 VSUBS 0.18841f
C764 VTAIL.t11 VSUBS 0.080402f
C765 VTAIL.n67 VSUBS 0.028064f
C766 VTAIL.n68 VSUBS 0.028148f
C767 VTAIL.n69 VSUBS 0.015831f
C768 VTAIL.n70 VSUBS 1.02393f
C769 VTAIL.n71 VSUBS 0.029461f
C770 VTAIL.n72 VSUBS 0.015831f
C771 VTAIL.n73 VSUBS 0.016762f
C772 VTAIL.n74 VSUBS 0.037419f
C773 VTAIL.n75 VSUBS 0.037419f
C774 VTAIL.n76 VSUBS 0.016762f
C775 VTAIL.n77 VSUBS 0.015831f
C776 VTAIL.n78 VSUBS 0.029461f
C777 VTAIL.n79 VSUBS 0.029461f
C778 VTAIL.n80 VSUBS 0.015831f
C779 VTAIL.n81 VSUBS 0.016762f
C780 VTAIL.n82 VSUBS 0.037419f
C781 VTAIL.n83 VSUBS 0.037419f
C782 VTAIL.n84 VSUBS 0.016762f
C783 VTAIL.n85 VSUBS 0.015831f
C784 VTAIL.n86 VSUBS 0.029461f
C785 VTAIL.n87 VSUBS 0.029461f
C786 VTAIL.n88 VSUBS 0.015831f
C787 VTAIL.n89 VSUBS 0.016297f
C788 VTAIL.n90 VSUBS 0.016297f
C789 VTAIL.n91 VSUBS 0.037419f
C790 VTAIL.n92 VSUBS 0.090167f
C791 VTAIL.n93 VSUBS 0.016762f
C792 VTAIL.n94 VSUBS 0.015831f
C793 VTAIL.n95 VSUBS 0.076147f
C794 VTAIL.n96 VSUBS 0.045561f
C795 VTAIL.n97 VSUBS 0.270723f
C796 VTAIL.t7 VSUBS 0.203009f
C797 VTAIL.t9 VSUBS 0.203009f
C798 VTAIL.n98 VSUBS 1.37884f
C799 VTAIL.n99 VSUBS 0.82875f
C800 VTAIL.n100 VSUBS 0.032248f
C801 VTAIL.n101 VSUBS 0.029461f
C802 VTAIL.n102 VSUBS 0.015831f
C803 VTAIL.n103 VSUBS 0.037419f
C804 VTAIL.n104 VSUBS 0.016762f
C805 VTAIL.n105 VSUBS 0.029461f
C806 VTAIL.n106 VSUBS 0.015831f
C807 VTAIL.n107 VSUBS 0.037419f
C808 VTAIL.n108 VSUBS 0.037419f
C809 VTAIL.n109 VSUBS 0.016762f
C810 VTAIL.n110 VSUBS 0.029461f
C811 VTAIL.n111 VSUBS 0.015831f
C812 VTAIL.n112 VSUBS 0.037419f
C813 VTAIL.n113 VSUBS 0.016762f
C814 VTAIL.n114 VSUBS 0.18841f
C815 VTAIL.t5 VSUBS 0.080402f
C816 VTAIL.n115 VSUBS 0.028064f
C817 VTAIL.n116 VSUBS 0.028148f
C818 VTAIL.n117 VSUBS 0.015831f
C819 VTAIL.n118 VSUBS 1.02393f
C820 VTAIL.n119 VSUBS 0.029461f
C821 VTAIL.n120 VSUBS 0.015831f
C822 VTAIL.n121 VSUBS 0.016762f
C823 VTAIL.n122 VSUBS 0.037419f
C824 VTAIL.n123 VSUBS 0.037419f
C825 VTAIL.n124 VSUBS 0.016762f
C826 VTAIL.n125 VSUBS 0.015831f
C827 VTAIL.n126 VSUBS 0.029461f
C828 VTAIL.n127 VSUBS 0.029461f
C829 VTAIL.n128 VSUBS 0.015831f
C830 VTAIL.n129 VSUBS 0.016762f
C831 VTAIL.n130 VSUBS 0.037419f
C832 VTAIL.n131 VSUBS 0.037419f
C833 VTAIL.n132 VSUBS 0.016762f
C834 VTAIL.n133 VSUBS 0.015831f
C835 VTAIL.n134 VSUBS 0.029461f
C836 VTAIL.n135 VSUBS 0.029461f
C837 VTAIL.n136 VSUBS 0.015831f
C838 VTAIL.n137 VSUBS 0.016297f
C839 VTAIL.n138 VSUBS 0.016297f
C840 VTAIL.n139 VSUBS 0.037419f
C841 VTAIL.n140 VSUBS 0.090167f
C842 VTAIL.n141 VSUBS 0.016762f
C843 VTAIL.n142 VSUBS 0.015831f
C844 VTAIL.n143 VSUBS 0.076147f
C845 VTAIL.n144 VSUBS 0.045561f
C846 VTAIL.n145 VSUBS 1.40539f
C847 VTAIL.n146 VSUBS 0.032248f
C848 VTAIL.n147 VSUBS 0.029461f
C849 VTAIL.n148 VSUBS 0.015831f
C850 VTAIL.n149 VSUBS 0.037419f
C851 VTAIL.n150 VSUBS 0.016762f
C852 VTAIL.n151 VSUBS 0.029461f
C853 VTAIL.n152 VSUBS 0.015831f
C854 VTAIL.n153 VSUBS 0.037419f
C855 VTAIL.n154 VSUBS 0.016762f
C856 VTAIL.n155 VSUBS 0.029461f
C857 VTAIL.n156 VSUBS 0.015831f
C858 VTAIL.n157 VSUBS 0.037419f
C859 VTAIL.n158 VSUBS 0.016762f
C860 VTAIL.n159 VSUBS 0.18841f
C861 VTAIL.t0 VSUBS 0.080402f
C862 VTAIL.n160 VSUBS 0.028064f
C863 VTAIL.n161 VSUBS 0.028148f
C864 VTAIL.n162 VSUBS 0.015831f
C865 VTAIL.n163 VSUBS 1.02393f
C866 VTAIL.n164 VSUBS 0.029461f
C867 VTAIL.n165 VSUBS 0.015831f
C868 VTAIL.n166 VSUBS 0.016762f
C869 VTAIL.n167 VSUBS 0.037419f
C870 VTAIL.n168 VSUBS 0.037419f
C871 VTAIL.n169 VSUBS 0.016762f
C872 VTAIL.n170 VSUBS 0.015831f
C873 VTAIL.n171 VSUBS 0.029461f
C874 VTAIL.n172 VSUBS 0.029461f
C875 VTAIL.n173 VSUBS 0.015831f
C876 VTAIL.n174 VSUBS 0.016762f
C877 VTAIL.n175 VSUBS 0.037419f
C878 VTAIL.n176 VSUBS 0.037419f
C879 VTAIL.n177 VSUBS 0.037419f
C880 VTAIL.n178 VSUBS 0.016762f
C881 VTAIL.n179 VSUBS 0.015831f
C882 VTAIL.n180 VSUBS 0.029461f
C883 VTAIL.n181 VSUBS 0.029461f
C884 VTAIL.n182 VSUBS 0.015831f
C885 VTAIL.n183 VSUBS 0.016297f
C886 VTAIL.n184 VSUBS 0.016297f
C887 VTAIL.n185 VSUBS 0.037419f
C888 VTAIL.n186 VSUBS 0.090167f
C889 VTAIL.n187 VSUBS 0.016762f
C890 VTAIL.n188 VSUBS 0.015831f
C891 VTAIL.n189 VSUBS 0.076147f
C892 VTAIL.n190 VSUBS 0.045561f
C893 VTAIL.n191 VSUBS 1.36713f
C894 VDD1.n0 VSUBS 0.024144f
C895 VDD1.n1 VSUBS 0.022057f
C896 VDD1.n2 VSUBS 0.011853f
C897 VDD1.n3 VSUBS 0.028015f
C898 VDD1.n4 VSUBS 0.01255f
C899 VDD1.n5 VSUBS 0.022057f
C900 VDD1.n6 VSUBS 0.011853f
C901 VDD1.n7 VSUBS 0.028015f
C902 VDD1.n8 VSUBS 0.028015f
C903 VDD1.n9 VSUBS 0.01255f
C904 VDD1.n10 VSUBS 0.022057f
C905 VDD1.n11 VSUBS 0.011853f
C906 VDD1.n12 VSUBS 0.028015f
C907 VDD1.n13 VSUBS 0.01255f
C908 VDD1.n14 VSUBS 0.141062f
C909 VDD1.t0 VSUBS 0.060197f
C910 VDD1.n15 VSUBS 0.021011f
C911 VDD1.n16 VSUBS 0.021074f
C912 VDD1.n17 VSUBS 0.011853f
C913 VDD1.n18 VSUBS 0.76661f
C914 VDD1.n19 VSUBS 0.022057f
C915 VDD1.n20 VSUBS 0.011853f
C916 VDD1.n21 VSUBS 0.01255f
C917 VDD1.n22 VSUBS 0.028015f
C918 VDD1.n23 VSUBS 0.028015f
C919 VDD1.n24 VSUBS 0.01255f
C920 VDD1.n25 VSUBS 0.011853f
C921 VDD1.n26 VSUBS 0.022057f
C922 VDD1.n27 VSUBS 0.022057f
C923 VDD1.n28 VSUBS 0.011853f
C924 VDD1.n29 VSUBS 0.01255f
C925 VDD1.n30 VSUBS 0.028015f
C926 VDD1.n31 VSUBS 0.028015f
C927 VDD1.n32 VSUBS 0.01255f
C928 VDD1.n33 VSUBS 0.011853f
C929 VDD1.n34 VSUBS 0.022057f
C930 VDD1.n35 VSUBS 0.022057f
C931 VDD1.n36 VSUBS 0.011853f
C932 VDD1.n37 VSUBS 0.012201f
C933 VDD1.n38 VSUBS 0.012201f
C934 VDD1.n39 VSUBS 0.028015f
C935 VDD1.n40 VSUBS 0.067508f
C936 VDD1.n41 VSUBS 0.01255f
C937 VDD1.n42 VSUBS 0.011853f
C938 VDD1.n43 VSUBS 0.057011f
C939 VDD1.n44 VSUBS 0.051808f
C940 VDD1.n45 VSUBS 0.024144f
C941 VDD1.n46 VSUBS 0.022057f
C942 VDD1.n47 VSUBS 0.011853f
C943 VDD1.n48 VSUBS 0.028015f
C944 VDD1.n49 VSUBS 0.01255f
C945 VDD1.n50 VSUBS 0.022057f
C946 VDD1.n51 VSUBS 0.011853f
C947 VDD1.n52 VSUBS 0.028015f
C948 VDD1.n53 VSUBS 0.01255f
C949 VDD1.n54 VSUBS 0.022057f
C950 VDD1.n55 VSUBS 0.011853f
C951 VDD1.n56 VSUBS 0.028015f
C952 VDD1.n57 VSUBS 0.01255f
C953 VDD1.n58 VSUBS 0.141062f
C954 VDD1.t3 VSUBS 0.060197f
C955 VDD1.n59 VSUBS 0.021011f
C956 VDD1.n60 VSUBS 0.021074f
C957 VDD1.n61 VSUBS 0.011853f
C958 VDD1.n62 VSUBS 0.76661f
C959 VDD1.n63 VSUBS 0.022057f
C960 VDD1.n64 VSUBS 0.011853f
C961 VDD1.n65 VSUBS 0.01255f
C962 VDD1.n66 VSUBS 0.028015f
C963 VDD1.n67 VSUBS 0.028015f
C964 VDD1.n68 VSUBS 0.01255f
C965 VDD1.n69 VSUBS 0.011853f
C966 VDD1.n70 VSUBS 0.022057f
C967 VDD1.n71 VSUBS 0.022057f
C968 VDD1.n72 VSUBS 0.011853f
C969 VDD1.n73 VSUBS 0.01255f
C970 VDD1.n74 VSUBS 0.028015f
C971 VDD1.n75 VSUBS 0.028015f
C972 VDD1.n76 VSUBS 0.028015f
C973 VDD1.n77 VSUBS 0.01255f
C974 VDD1.n78 VSUBS 0.011853f
C975 VDD1.n79 VSUBS 0.022057f
C976 VDD1.n80 VSUBS 0.022057f
C977 VDD1.n81 VSUBS 0.011853f
C978 VDD1.n82 VSUBS 0.012201f
C979 VDD1.n83 VSUBS 0.012201f
C980 VDD1.n84 VSUBS 0.028015f
C981 VDD1.n85 VSUBS 0.067508f
C982 VDD1.n86 VSUBS 0.01255f
C983 VDD1.n87 VSUBS 0.011853f
C984 VDD1.n88 VSUBS 0.057011f
C985 VDD1.n89 VSUBS 0.051415f
C986 VDD1.t5 VSUBS 0.151992f
C987 VDD1.t1 VSUBS 0.151992f
C988 VDD1.n90 VSUBS 1.12636f
C989 VDD1.n91 VSUBS 1.95675f
C990 VDD1.t2 VSUBS 0.151992f
C991 VDD1.t4 VSUBS 0.151992f
C992 VDD1.n92 VSUBS 1.12462f
C993 VDD1.n93 VSUBS 2.10089f
C994 VP.n0 VSUBS 0.064176f
C995 VP.t3 VSUBS 1.43559f
C996 VP.n1 VSUBS 0.542027f
C997 VP.n2 VSUBS 0.064176f
C998 VP.n3 VSUBS 0.064176f
C999 VP.t4 VSUBS 1.52973f
C1000 VP.t0 VSUBS 1.43559f
C1001 VP.n4 VSUBS 0.604884f
C1002 VP.t2 VSUBS 1.5872f
C1003 VP.n5 VSUBS 0.626118f
C1004 VP.n6 VSUBS 0.252137f
C1005 VP.n7 VSUBS 0.075414f
C1006 VP.n8 VSUBS 0.030775f
C1007 VP.n9 VSUBS 0.637985f
C1008 VP.n10 VSUBS 1.93504f
C1009 VP.n11 VSUBS 1.97694f
C1010 VP.t5 VSUBS 1.52973f
C1011 VP.n12 VSUBS 0.637985f
C1012 VP.n13 VSUBS 0.030775f
C1013 VP.n14 VSUBS 0.075414f
C1014 VP.n15 VSUBS 0.048094f
C1015 VP.n16 VSUBS 0.048094f
C1016 VP.n17 VSUBS 0.075414f
C1017 VP.n18 VSUBS 0.030775f
C1018 VP.t1 VSUBS 1.52973f
C1019 VP.n19 VSUBS 0.637985f
C1020 VP.n20 VSUBS 0.045042f
.ends

