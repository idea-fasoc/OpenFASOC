* NGSPICE file created from diff_pair_sample_1090.ext - technology: sky130A

.subckt diff_pair_sample_1090 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=0 ps=0 w=7.18 l=3.48
X1 B.t8 B.t6 B.t7 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=0 ps=0 w=7.18 l=3.48
X2 B.t5 B.t3 B.t4 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=0 ps=0 w=7.18 l=3.48
X3 VTAIL.t11 VP.t0 VDD1.t1 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=1.1847 ps=7.51 w=7.18 l=3.48
X4 VDD2.t5 VN.t0 VTAIL.t2 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=1.1847 ps=7.51 w=7.18 l=3.48
X5 VTAIL.t3 VN.t1 VDD2.t4 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=1.1847 ps=7.51 w=7.18 l=3.48
X6 VDD2.t3 VN.t2 VTAIL.t0 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=2.8002 ps=15.14 w=7.18 l=3.48
X7 VTAIL.t5 VN.t3 VDD2.t2 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=1.1847 ps=7.51 w=7.18 l=3.48
X8 B.t2 B.t0 B.t1 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=0 ps=0 w=7.18 l=3.48
X9 VTAIL.t10 VP.t1 VDD1.t0 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=1.1847 ps=7.51 w=7.18 l=3.48
X10 VDD1.t5 VP.t2 VTAIL.t9 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=1.1847 ps=7.51 w=7.18 l=3.48
X11 VDD2.t1 VN.t4 VTAIL.t4 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=2.8002 ps=15.14 w=7.18 l=3.48
X12 VDD1.t4 VP.t3 VTAIL.t8 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=1.1847 ps=7.51 w=7.18 l=3.48
X13 VDD1.t3 VP.t4 VTAIL.t7 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=2.8002 ps=15.14 w=7.18 l=3.48
X14 VDD1.t2 VP.t5 VTAIL.t6 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=1.1847 pd=7.51 as=2.8002 ps=15.14 w=7.18 l=3.48
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n4018_n2404# sky130_fd_pr__pfet_01v8 ad=2.8002 pd=15.14 as=1.1847 ps=7.51 w=7.18 l=3.48
R0 B.n518 B.n517 585
R1 B.n519 B.n64 585
R2 B.n521 B.n520 585
R3 B.n522 B.n63 585
R4 B.n524 B.n523 585
R5 B.n525 B.n62 585
R6 B.n527 B.n526 585
R7 B.n528 B.n61 585
R8 B.n530 B.n529 585
R9 B.n531 B.n60 585
R10 B.n533 B.n532 585
R11 B.n534 B.n59 585
R12 B.n536 B.n535 585
R13 B.n537 B.n58 585
R14 B.n539 B.n538 585
R15 B.n540 B.n57 585
R16 B.n542 B.n541 585
R17 B.n543 B.n56 585
R18 B.n545 B.n544 585
R19 B.n546 B.n55 585
R20 B.n548 B.n547 585
R21 B.n549 B.n54 585
R22 B.n551 B.n550 585
R23 B.n552 B.n53 585
R24 B.n554 B.n553 585
R25 B.n555 B.n52 585
R26 B.n557 B.n556 585
R27 B.n559 B.n49 585
R28 B.n561 B.n560 585
R29 B.n562 B.n48 585
R30 B.n564 B.n563 585
R31 B.n565 B.n47 585
R32 B.n567 B.n566 585
R33 B.n568 B.n46 585
R34 B.n570 B.n569 585
R35 B.n571 B.n45 585
R36 B.n573 B.n572 585
R37 B.n575 B.n574 585
R38 B.n576 B.n41 585
R39 B.n578 B.n577 585
R40 B.n579 B.n40 585
R41 B.n581 B.n580 585
R42 B.n582 B.n39 585
R43 B.n584 B.n583 585
R44 B.n585 B.n38 585
R45 B.n587 B.n586 585
R46 B.n588 B.n37 585
R47 B.n590 B.n589 585
R48 B.n591 B.n36 585
R49 B.n593 B.n592 585
R50 B.n594 B.n35 585
R51 B.n596 B.n595 585
R52 B.n597 B.n34 585
R53 B.n599 B.n598 585
R54 B.n600 B.n33 585
R55 B.n602 B.n601 585
R56 B.n603 B.n32 585
R57 B.n605 B.n604 585
R58 B.n606 B.n31 585
R59 B.n608 B.n607 585
R60 B.n609 B.n30 585
R61 B.n611 B.n610 585
R62 B.n612 B.n29 585
R63 B.n614 B.n613 585
R64 B.n516 B.n65 585
R65 B.n515 B.n514 585
R66 B.n513 B.n66 585
R67 B.n512 B.n511 585
R68 B.n510 B.n67 585
R69 B.n509 B.n508 585
R70 B.n507 B.n68 585
R71 B.n506 B.n505 585
R72 B.n504 B.n69 585
R73 B.n503 B.n502 585
R74 B.n501 B.n70 585
R75 B.n500 B.n499 585
R76 B.n498 B.n71 585
R77 B.n497 B.n496 585
R78 B.n495 B.n72 585
R79 B.n494 B.n493 585
R80 B.n492 B.n73 585
R81 B.n491 B.n490 585
R82 B.n489 B.n74 585
R83 B.n488 B.n487 585
R84 B.n486 B.n75 585
R85 B.n485 B.n484 585
R86 B.n483 B.n76 585
R87 B.n482 B.n481 585
R88 B.n480 B.n77 585
R89 B.n479 B.n478 585
R90 B.n477 B.n78 585
R91 B.n476 B.n475 585
R92 B.n474 B.n79 585
R93 B.n473 B.n472 585
R94 B.n471 B.n80 585
R95 B.n470 B.n469 585
R96 B.n468 B.n81 585
R97 B.n467 B.n466 585
R98 B.n465 B.n82 585
R99 B.n464 B.n463 585
R100 B.n462 B.n83 585
R101 B.n461 B.n460 585
R102 B.n459 B.n84 585
R103 B.n458 B.n457 585
R104 B.n456 B.n85 585
R105 B.n455 B.n454 585
R106 B.n453 B.n86 585
R107 B.n452 B.n451 585
R108 B.n450 B.n87 585
R109 B.n449 B.n448 585
R110 B.n447 B.n88 585
R111 B.n446 B.n445 585
R112 B.n444 B.n89 585
R113 B.n443 B.n442 585
R114 B.n441 B.n90 585
R115 B.n440 B.n439 585
R116 B.n438 B.n91 585
R117 B.n437 B.n436 585
R118 B.n435 B.n92 585
R119 B.n434 B.n433 585
R120 B.n432 B.n93 585
R121 B.n431 B.n430 585
R122 B.n429 B.n94 585
R123 B.n428 B.n427 585
R124 B.n426 B.n95 585
R125 B.n425 B.n424 585
R126 B.n423 B.n96 585
R127 B.n422 B.n421 585
R128 B.n420 B.n97 585
R129 B.n419 B.n418 585
R130 B.n417 B.n98 585
R131 B.n416 B.n415 585
R132 B.n414 B.n99 585
R133 B.n413 B.n412 585
R134 B.n411 B.n100 585
R135 B.n410 B.n409 585
R136 B.n408 B.n101 585
R137 B.n407 B.n406 585
R138 B.n405 B.n102 585
R139 B.n404 B.n403 585
R140 B.n402 B.n103 585
R141 B.n401 B.n400 585
R142 B.n399 B.n104 585
R143 B.n398 B.n397 585
R144 B.n396 B.n105 585
R145 B.n395 B.n394 585
R146 B.n393 B.n106 585
R147 B.n392 B.n391 585
R148 B.n390 B.n107 585
R149 B.n389 B.n388 585
R150 B.n387 B.n108 585
R151 B.n386 B.n385 585
R152 B.n384 B.n109 585
R153 B.n383 B.n382 585
R154 B.n381 B.n110 585
R155 B.n380 B.n379 585
R156 B.n378 B.n111 585
R157 B.n377 B.n376 585
R158 B.n375 B.n112 585
R159 B.n374 B.n373 585
R160 B.n372 B.n113 585
R161 B.n371 B.n370 585
R162 B.n369 B.n114 585
R163 B.n368 B.n367 585
R164 B.n366 B.n115 585
R165 B.n365 B.n364 585
R166 B.n363 B.n116 585
R167 B.n362 B.n361 585
R168 B.n360 B.n117 585
R169 B.n359 B.n358 585
R170 B.n357 B.n118 585
R171 B.n260 B.n259 585
R172 B.n261 B.n154 585
R173 B.n263 B.n262 585
R174 B.n264 B.n153 585
R175 B.n266 B.n265 585
R176 B.n267 B.n152 585
R177 B.n269 B.n268 585
R178 B.n270 B.n151 585
R179 B.n272 B.n271 585
R180 B.n273 B.n150 585
R181 B.n275 B.n274 585
R182 B.n276 B.n149 585
R183 B.n278 B.n277 585
R184 B.n279 B.n148 585
R185 B.n281 B.n280 585
R186 B.n282 B.n147 585
R187 B.n284 B.n283 585
R188 B.n285 B.n146 585
R189 B.n287 B.n286 585
R190 B.n288 B.n145 585
R191 B.n290 B.n289 585
R192 B.n291 B.n144 585
R193 B.n293 B.n292 585
R194 B.n294 B.n143 585
R195 B.n296 B.n295 585
R196 B.n297 B.n142 585
R197 B.n299 B.n298 585
R198 B.n301 B.n139 585
R199 B.n303 B.n302 585
R200 B.n304 B.n138 585
R201 B.n306 B.n305 585
R202 B.n307 B.n137 585
R203 B.n309 B.n308 585
R204 B.n310 B.n136 585
R205 B.n312 B.n311 585
R206 B.n313 B.n135 585
R207 B.n315 B.n314 585
R208 B.n317 B.n316 585
R209 B.n318 B.n131 585
R210 B.n320 B.n319 585
R211 B.n321 B.n130 585
R212 B.n323 B.n322 585
R213 B.n324 B.n129 585
R214 B.n326 B.n325 585
R215 B.n327 B.n128 585
R216 B.n329 B.n328 585
R217 B.n330 B.n127 585
R218 B.n332 B.n331 585
R219 B.n333 B.n126 585
R220 B.n335 B.n334 585
R221 B.n336 B.n125 585
R222 B.n338 B.n337 585
R223 B.n339 B.n124 585
R224 B.n341 B.n340 585
R225 B.n342 B.n123 585
R226 B.n344 B.n343 585
R227 B.n345 B.n122 585
R228 B.n347 B.n346 585
R229 B.n348 B.n121 585
R230 B.n350 B.n349 585
R231 B.n351 B.n120 585
R232 B.n353 B.n352 585
R233 B.n354 B.n119 585
R234 B.n356 B.n355 585
R235 B.n258 B.n155 585
R236 B.n257 B.n256 585
R237 B.n255 B.n156 585
R238 B.n254 B.n253 585
R239 B.n252 B.n157 585
R240 B.n251 B.n250 585
R241 B.n249 B.n158 585
R242 B.n248 B.n247 585
R243 B.n246 B.n159 585
R244 B.n245 B.n244 585
R245 B.n243 B.n160 585
R246 B.n242 B.n241 585
R247 B.n240 B.n161 585
R248 B.n239 B.n238 585
R249 B.n237 B.n162 585
R250 B.n236 B.n235 585
R251 B.n234 B.n163 585
R252 B.n233 B.n232 585
R253 B.n231 B.n164 585
R254 B.n230 B.n229 585
R255 B.n228 B.n165 585
R256 B.n227 B.n226 585
R257 B.n225 B.n166 585
R258 B.n224 B.n223 585
R259 B.n222 B.n167 585
R260 B.n221 B.n220 585
R261 B.n219 B.n168 585
R262 B.n218 B.n217 585
R263 B.n216 B.n169 585
R264 B.n215 B.n214 585
R265 B.n213 B.n170 585
R266 B.n212 B.n211 585
R267 B.n210 B.n171 585
R268 B.n209 B.n208 585
R269 B.n207 B.n172 585
R270 B.n206 B.n205 585
R271 B.n204 B.n173 585
R272 B.n203 B.n202 585
R273 B.n201 B.n174 585
R274 B.n200 B.n199 585
R275 B.n198 B.n175 585
R276 B.n197 B.n196 585
R277 B.n195 B.n176 585
R278 B.n194 B.n193 585
R279 B.n192 B.n177 585
R280 B.n191 B.n190 585
R281 B.n189 B.n178 585
R282 B.n188 B.n187 585
R283 B.n186 B.n179 585
R284 B.n185 B.n184 585
R285 B.n183 B.n180 585
R286 B.n182 B.n181 585
R287 B.n2 B.n0 585
R288 B.n693 B.n1 585
R289 B.n692 B.n691 585
R290 B.n690 B.n3 585
R291 B.n689 B.n688 585
R292 B.n687 B.n4 585
R293 B.n686 B.n685 585
R294 B.n684 B.n5 585
R295 B.n683 B.n682 585
R296 B.n681 B.n6 585
R297 B.n680 B.n679 585
R298 B.n678 B.n7 585
R299 B.n677 B.n676 585
R300 B.n675 B.n8 585
R301 B.n674 B.n673 585
R302 B.n672 B.n9 585
R303 B.n671 B.n670 585
R304 B.n669 B.n10 585
R305 B.n668 B.n667 585
R306 B.n666 B.n11 585
R307 B.n665 B.n664 585
R308 B.n663 B.n12 585
R309 B.n662 B.n661 585
R310 B.n660 B.n13 585
R311 B.n659 B.n658 585
R312 B.n657 B.n14 585
R313 B.n656 B.n655 585
R314 B.n654 B.n15 585
R315 B.n653 B.n652 585
R316 B.n651 B.n16 585
R317 B.n650 B.n649 585
R318 B.n648 B.n17 585
R319 B.n647 B.n646 585
R320 B.n645 B.n18 585
R321 B.n644 B.n643 585
R322 B.n642 B.n19 585
R323 B.n641 B.n640 585
R324 B.n639 B.n20 585
R325 B.n638 B.n637 585
R326 B.n636 B.n21 585
R327 B.n635 B.n634 585
R328 B.n633 B.n22 585
R329 B.n632 B.n631 585
R330 B.n630 B.n23 585
R331 B.n629 B.n628 585
R332 B.n627 B.n24 585
R333 B.n626 B.n625 585
R334 B.n624 B.n25 585
R335 B.n623 B.n622 585
R336 B.n621 B.n26 585
R337 B.n620 B.n619 585
R338 B.n618 B.n27 585
R339 B.n617 B.n616 585
R340 B.n615 B.n28 585
R341 B.n695 B.n694 585
R342 B.n260 B.n155 526.135
R343 B.n615 B.n614 526.135
R344 B.n357 B.n356 526.135
R345 B.n518 B.n65 526.135
R346 B.n132 B.t8 362.695
R347 B.n50 B.t10 362.695
R348 B.n140 B.t2 362.695
R349 B.n42 B.t4 362.695
R350 B.n133 B.t7 288.805
R351 B.n51 B.t11 288.805
R352 B.n141 B.t1 288.805
R353 B.n43 B.t5 288.805
R354 B.n132 B.t6 258.8
R355 B.n140 B.t0 258.8
R356 B.n42 B.t3 258.8
R357 B.n50 B.t9 258.8
R358 B.n256 B.n155 163.367
R359 B.n256 B.n255 163.367
R360 B.n255 B.n254 163.367
R361 B.n254 B.n157 163.367
R362 B.n250 B.n157 163.367
R363 B.n250 B.n249 163.367
R364 B.n249 B.n248 163.367
R365 B.n248 B.n159 163.367
R366 B.n244 B.n159 163.367
R367 B.n244 B.n243 163.367
R368 B.n243 B.n242 163.367
R369 B.n242 B.n161 163.367
R370 B.n238 B.n161 163.367
R371 B.n238 B.n237 163.367
R372 B.n237 B.n236 163.367
R373 B.n236 B.n163 163.367
R374 B.n232 B.n163 163.367
R375 B.n232 B.n231 163.367
R376 B.n231 B.n230 163.367
R377 B.n230 B.n165 163.367
R378 B.n226 B.n165 163.367
R379 B.n226 B.n225 163.367
R380 B.n225 B.n224 163.367
R381 B.n224 B.n167 163.367
R382 B.n220 B.n167 163.367
R383 B.n220 B.n219 163.367
R384 B.n219 B.n218 163.367
R385 B.n218 B.n169 163.367
R386 B.n214 B.n169 163.367
R387 B.n214 B.n213 163.367
R388 B.n213 B.n212 163.367
R389 B.n212 B.n171 163.367
R390 B.n208 B.n171 163.367
R391 B.n208 B.n207 163.367
R392 B.n207 B.n206 163.367
R393 B.n206 B.n173 163.367
R394 B.n202 B.n173 163.367
R395 B.n202 B.n201 163.367
R396 B.n201 B.n200 163.367
R397 B.n200 B.n175 163.367
R398 B.n196 B.n175 163.367
R399 B.n196 B.n195 163.367
R400 B.n195 B.n194 163.367
R401 B.n194 B.n177 163.367
R402 B.n190 B.n177 163.367
R403 B.n190 B.n189 163.367
R404 B.n189 B.n188 163.367
R405 B.n188 B.n179 163.367
R406 B.n184 B.n179 163.367
R407 B.n184 B.n183 163.367
R408 B.n183 B.n182 163.367
R409 B.n182 B.n2 163.367
R410 B.n694 B.n2 163.367
R411 B.n694 B.n693 163.367
R412 B.n693 B.n692 163.367
R413 B.n692 B.n3 163.367
R414 B.n688 B.n3 163.367
R415 B.n688 B.n687 163.367
R416 B.n687 B.n686 163.367
R417 B.n686 B.n5 163.367
R418 B.n682 B.n5 163.367
R419 B.n682 B.n681 163.367
R420 B.n681 B.n680 163.367
R421 B.n680 B.n7 163.367
R422 B.n676 B.n7 163.367
R423 B.n676 B.n675 163.367
R424 B.n675 B.n674 163.367
R425 B.n674 B.n9 163.367
R426 B.n670 B.n9 163.367
R427 B.n670 B.n669 163.367
R428 B.n669 B.n668 163.367
R429 B.n668 B.n11 163.367
R430 B.n664 B.n11 163.367
R431 B.n664 B.n663 163.367
R432 B.n663 B.n662 163.367
R433 B.n662 B.n13 163.367
R434 B.n658 B.n13 163.367
R435 B.n658 B.n657 163.367
R436 B.n657 B.n656 163.367
R437 B.n656 B.n15 163.367
R438 B.n652 B.n15 163.367
R439 B.n652 B.n651 163.367
R440 B.n651 B.n650 163.367
R441 B.n650 B.n17 163.367
R442 B.n646 B.n17 163.367
R443 B.n646 B.n645 163.367
R444 B.n645 B.n644 163.367
R445 B.n644 B.n19 163.367
R446 B.n640 B.n19 163.367
R447 B.n640 B.n639 163.367
R448 B.n639 B.n638 163.367
R449 B.n638 B.n21 163.367
R450 B.n634 B.n21 163.367
R451 B.n634 B.n633 163.367
R452 B.n633 B.n632 163.367
R453 B.n632 B.n23 163.367
R454 B.n628 B.n23 163.367
R455 B.n628 B.n627 163.367
R456 B.n627 B.n626 163.367
R457 B.n626 B.n25 163.367
R458 B.n622 B.n25 163.367
R459 B.n622 B.n621 163.367
R460 B.n621 B.n620 163.367
R461 B.n620 B.n27 163.367
R462 B.n616 B.n27 163.367
R463 B.n616 B.n615 163.367
R464 B.n261 B.n260 163.367
R465 B.n262 B.n261 163.367
R466 B.n262 B.n153 163.367
R467 B.n266 B.n153 163.367
R468 B.n267 B.n266 163.367
R469 B.n268 B.n267 163.367
R470 B.n268 B.n151 163.367
R471 B.n272 B.n151 163.367
R472 B.n273 B.n272 163.367
R473 B.n274 B.n273 163.367
R474 B.n274 B.n149 163.367
R475 B.n278 B.n149 163.367
R476 B.n279 B.n278 163.367
R477 B.n280 B.n279 163.367
R478 B.n280 B.n147 163.367
R479 B.n284 B.n147 163.367
R480 B.n285 B.n284 163.367
R481 B.n286 B.n285 163.367
R482 B.n286 B.n145 163.367
R483 B.n290 B.n145 163.367
R484 B.n291 B.n290 163.367
R485 B.n292 B.n291 163.367
R486 B.n292 B.n143 163.367
R487 B.n296 B.n143 163.367
R488 B.n297 B.n296 163.367
R489 B.n298 B.n297 163.367
R490 B.n298 B.n139 163.367
R491 B.n303 B.n139 163.367
R492 B.n304 B.n303 163.367
R493 B.n305 B.n304 163.367
R494 B.n305 B.n137 163.367
R495 B.n309 B.n137 163.367
R496 B.n310 B.n309 163.367
R497 B.n311 B.n310 163.367
R498 B.n311 B.n135 163.367
R499 B.n315 B.n135 163.367
R500 B.n316 B.n315 163.367
R501 B.n316 B.n131 163.367
R502 B.n320 B.n131 163.367
R503 B.n321 B.n320 163.367
R504 B.n322 B.n321 163.367
R505 B.n322 B.n129 163.367
R506 B.n326 B.n129 163.367
R507 B.n327 B.n326 163.367
R508 B.n328 B.n327 163.367
R509 B.n328 B.n127 163.367
R510 B.n332 B.n127 163.367
R511 B.n333 B.n332 163.367
R512 B.n334 B.n333 163.367
R513 B.n334 B.n125 163.367
R514 B.n338 B.n125 163.367
R515 B.n339 B.n338 163.367
R516 B.n340 B.n339 163.367
R517 B.n340 B.n123 163.367
R518 B.n344 B.n123 163.367
R519 B.n345 B.n344 163.367
R520 B.n346 B.n345 163.367
R521 B.n346 B.n121 163.367
R522 B.n350 B.n121 163.367
R523 B.n351 B.n350 163.367
R524 B.n352 B.n351 163.367
R525 B.n352 B.n119 163.367
R526 B.n356 B.n119 163.367
R527 B.n358 B.n357 163.367
R528 B.n358 B.n117 163.367
R529 B.n362 B.n117 163.367
R530 B.n363 B.n362 163.367
R531 B.n364 B.n363 163.367
R532 B.n364 B.n115 163.367
R533 B.n368 B.n115 163.367
R534 B.n369 B.n368 163.367
R535 B.n370 B.n369 163.367
R536 B.n370 B.n113 163.367
R537 B.n374 B.n113 163.367
R538 B.n375 B.n374 163.367
R539 B.n376 B.n375 163.367
R540 B.n376 B.n111 163.367
R541 B.n380 B.n111 163.367
R542 B.n381 B.n380 163.367
R543 B.n382 B.n381 163.367
R544 B.n382 B.n109 163.367
R545 B.n386 B.n109 163.367
R546 B.n387 B.n386 163.367
R547 B.n388 B.n387 163.367
R548 B.n388 B.n107 163.367
R549 B.n392 B.n107 163.367
R550 B.n393 B.n392 163.367
R551 B.n394 B.n393 163.367
R552 B.n394 B.n105 163.367
R553 B.n398 B.n105 163.367
R554 B.n399 B.n398 163.367
R555 B.n400 B.n399 163.367
R556 B.n400 B.n103 163.367
R557 B.n404 B.n103 163.367
R558 B.n405 B.n404 163.367
R559 B.n406 B.n405 163.367
R560 B.n406 B.n101 163.367
R561 B.n410 B.n101 163.367
R562 B.n411 B.n410 163.367
R563 B.n412 B.n411 163.367
R564 B.n412 B.n99 163.367
R565 B.n416 B.n99 163.367
R566 B.n417 B.n416 163.367
R567 B.n418 B.n417 163.367
R568 B.n418 B.n97 163.367
R569 B.n422 B.n97 163.367
R570 B.n423 B.n422 163.367
R571 B.n424 B.n423 163.367
R572 B.n424 B.n95 163.367
R573 B.n428 B.n95 163.367
R574 B.n429 B.n428 163.367
R575 B.n430 B.n429 163.367
R576 B.n430 B.n93 163.367
R577 B.n434 B.n93 163.367
R578 B.n435 B.n434 163.367
R579 B.n436 B.n435 163.367
R580 B.n436 B.n91 163.367
R581 B.n440 B.n91 163.367
R582 B.n441 B.n440 163.367
R583 B.n442 B.n441 163.367
R584 B.n442 B.n89 163.367
R585 B.n446 B.n89 163.367
R586 B.n447 B.n446 163.367
R587 B.n448 B.n447 163.367
R588 B.n448 B.n87 163.367
R589 B.n452 B.n87 163.367
R590 B.n453 B.n452 163.367
R591 B.n454 B.n453 163.367
R592 B.n454 B.n85 163.367
R593 B.n458 B.n85 163.367
R594 B.n459 B.n458 163.367
R595 B.n460 B.n459 163.367
R596 B.n460 B.n83 163.367
R597 B.n464 B.n83 163.367
R598 B.n465 B.n464 163.367
R599 B.n466 B.n465 163.367
R600 B.n466 B.n81 163.367
R601 B.n470 B.n81 163.367
R602 B.n471 B.n470 163.367
R603 B.n472 B.n471 163.367
R604 B.n472 B.n79 163.367
R605 B.n476 B.n79 163.367
R606 B.n477 B.n476 163.367
R607 B.n478 B.n477 163.367
R608 B.n478 B.n77 163.367
R609 B.n482 B.n77 163.367
R610 B.n483 B.n482 163.367
R611 B.n484 B.n483 163.367
R612 B.n484 B.n75 163.367
R613 B.n488 B.n75 163.367
R614 B.n489 B.n488 163.367
R615 B.n490 B.n489 163.367
R616 B.n490 B.n73 163.367
R617 B.n494 B.n73 163.367
R618 B.n495 B.n494 163.367
R619 B.n496 B.n495 163.367
R620 B.n496 B.n71 163.367
R621 B.n500 B.n71 163.367
R622 B.n501 B.n500 163.367
R623 B.n502 B.n501 163.367
R624 B.n502 B.n69 163.367
R625 B.n506 B.n69 163.367
R626 B.n507 B.n506 163.367
R627 B.n508 B.n507 163.367
R628 B.n508 B.n67 163.367
R629 B.n512 B.n67 163.367
R630 B.n513 B.n512 163.367
R631 B.n514 B.n513 163.367
R632 B.n514 B.n65 163.367
R633 B.n614 B.n29 163.367
R634 B.n610 B.n29 163.367
R635 B.n610 B.n609 163.367
R636 B.n609 B.n608 163.367
R637 B.n608 B.n31 163.367
R638 B.n604 B.n31 163.367
R639 B.n604 B.n603 163.367
R640 B.n603 B.n602 163.367
R641 B.n602 B.n33 163.367
R642 B.n598 B.n33 163.367
R643 B.n598 B.n597 163.367
R644 B.n597 B.n596 163.367
R645 B.n596 B.n35 163.367
R646 B.n592 B.n35 163.367
R647 B.n592 B.n591 163.367
R648 B.n591 B.n590 163.367
R649 B.n590 B.n37 163.367
R650 B.n586 B.n37 163.367
R651 B.n586 B.n585 163.367
R652 B.n585 B.n584 163.367
R653 B.n584 B.n39 163.367
R654 B.n580 B.n39 163.367
R655 B.n580 B.n579 163.367
R656 B.n579 B.n578 163.367
R657 B.n578 B.n41 163.367
R658 B.n574 B.n41 163.367
R659 B.n574 B.n573 163.367
R660 B.n573 B.n45 163.367
R661 B.n569 B.n45 163.367
R662 B.n569 B.n568 163.367
R663 B.n568 B.n567 163.367
R664 B.n567 B.n47 163.367
R665 B.n563 B.n47 163.367
R666 B.n563 B.n562 163.367
R667 B.n562 B.n561 163.367
R668 B.n561 B.n49 163.367
R669 B.n556 B.n49 163.367
R670 B.n556 B.n555 163.367
R671 B.n555 B.n554 163.367
R672 B.n554 B.n53 163.367
R673 B.n550 B.n53 163.367
R674 B.n550 B.n549 163.367
R675 B.n549 B.n548 163.367
R676 B.n548 B.n55 163.367
R677 B.n544 B.n55 163.367
R678 B.n544 B.n543 163.367
R679 B.n543 B.n542 163.367
R680 B.n542 B.n57 163.367
R681 B.n538 B.n57 163.367
R682 B.n538 B.n537 163.367
R683 B.n537 B.n536 163.367
R684 B.n536 B.n59 163.367
R685 B.n532 B.n59 163.367
R686 B.n532 B.n531 163.367
R687 B.n531 B.n530 163.367
R688 B.n530 B.n61 163.367
R689 B.n526 B.n61 163.367
R690 B.n526 B.n525 163.367
R691 B.n525 B.n524 163.367
R692 B.n524 B.n63 163.367
R693 B.n520 B.n63 163.367
R694 B.n520 B.n519 163.367
R695 B.n519 B.n518 163.367
R696 B.n133 B.n132 73.8914
R697 B.n141 B.n140 73.8914
R698 B.n43 B.n42 73.8914
R699 B.n51 B.n50 73.8914
R700 B.n134 B.n133 59.5399
R701 B.n300 B.n141 59.5399
R702 B.n44 B.n43 59.5399
R703 B.n558 B.n51 59.5399
R704 B.n613 B.n28 34.1859
R705 B.n517 B.n516 34.1859
R706 B.n355 B.n118 34.1859
R707 B.n259 B.n258 34.1859
R708 B B.n695 18.0485
R709 B.n613 B.n612 10.6151
R710 B.n612 B.n611 10.6151
R711 B.n611 B.n30 10.6151
R712 B.n607 B.n30 10.6151
R713 B.n607 B.n606 10.6151
R714 B.n606 B.n605 10.6151
R715 B.n605 B.n32 10.6151
R716 B.n601 B.n32 10.6151
R717 B.n601 B.n600 10.6151
R718 B.n600 B.n599 10.6151
R719 B.n599 B.n34 10.6151
R720 B.n595 B.n34 10.6151
R721 B.n595 B.n594 10.6151
R722 B.n594 B.n593 10.6151
R723 B.n593 B.n36 10.6151
R724 B.n589 B.n36 10.6151
R725 B.n589 B.n588 10.6151
R726 B.n588 B.n587 10.6151
R727 B.n587 B.n38 10.6151
R728 B.n583 B.n38 10.6151
R729 B.n583 B.n582 10.6151
R730 B.n582 B.n581 10.6151
R731 B.n581 B.n40 10.6151
R732 B.n577 B.n40 10.6151
R733 B.n577 B.n576 10.6151
R734 B.n576 B.n575 10.6151
R735 B.n572 B.n571 10.6151
R736 B.n571 B.n570 10.6151
R737 B.n570 B.n46 10.6151
R738 B.n566 B.n46 10.6151
R739 B.n566 B.n565 10.6151
R740 B.n565 B.n564 10.6151
R741 B.n564 B.n48 10.6151
R742 B.n560 B.n48 10.6151
R743 B.n560 B.n559 10.6151
R744 B.n557 B.n52 10.6151
R745 B.n553 B.n52 10.6151
R746 B.n553 B.n552 10.6151
R747 B.n552 B.n551 10.6151
R748 B.n551 B.n54 10.6151
R749 B.n547 B.n54 10.6151
R750 B.n547 B.n546 10.6151
R751 B.n546 B.n545 10.6151
R752 B.n545 B.n56 10.6151
R753 B.n541 B.n56 10.6151
R754 B.n541 B.n540 10.6151
R755 B.n540 B.n539 10.6151
R756 B.n539 B.n58 10.6151
R757 B.n535 B.n58 10.6151
R758 B.n535 B.n534 10.6151
R759 B.n534 B.n533 10.6151
R760 B.n533 B.n60 10.6151
R761 B.n529 B.n60 10.6151
R762 B.n529 B.n528 10.6151
R763 B.n528 B.n527 10.6151
R764 B.n527 B.n62 10.6151
R765 B.n523 B.n62 10.6151
R766 B.n523 B.n522 10.6151
R767 B.n522 B.n521 10.6151
R768 B.n521 B.n64 10.6151
R769 B.n517 B.n64 10.6151
R770 B.n359 B.n118 10.6151
R771 B.n360 B.n359 10.6151
R772 B.n361 B.n360 10.6151
R773 B.n361 B.n116 10.6151
R774 B.n365 B.n116 10.6151
R775 B.n366 B.n365 10.6151
R776 B.n367 B.n366 10.6151
R777 B.n367 B.n114 10.6151
R778 B.n371 B.n114 10.6151
R779 B.n372 B.n371 10.6151
R780 B.n373 B.n372 10.6151
R781 B.n373 B.n112 10.6151
R782 B.n377 B.n112 10.6151
R783 B.n378 B.n377 10.6151
R784 B.n379 B.n378 10.6151
R785 B.n379 B.n110 10.6151
R786 B.n383 B.n110 10.6151
R787 B.n384 B.n383 10.6151
R788 B.n385 B.n384 10.6151
R789 B.n385 B.n108 10.6151
R790 B.n389 B.n108 10.6151
R791 B.n390 B.n389 10.6151
R792 B.n391 B.n390 10.6151
R793 B.n391 B.n106 10.6151
R794 B.n395 B.n106 10.6151
R795 B.n396 B.n395 10.6151
R796 B.n397 B.n396 10.6151
R797 B.n397 B.n104 10.6151
R798 B.n401 B.n104 10.6151
R799 B.n402 B.n401 10.6151
R800 B.n403 B.n402 10.6151
R801 B.n403 B.n102 10.6151
R802 B.n407 B.n102 10.6151
R803 B.n408 B.n407 10.6151
R804 B.n409 B.n408 10.6151
R805 B.n409 B.n100 10.6151
R806 B.n413 B.n100 10.6151
R807 B.n414 B.n413 10.6151
R808 B.n415 B.n414 10.6151
R809 B.n415 B.n98 10.6151
R810 B.n419 B.n98 10.6151
R811 B.n420 B.n419 10.6151
R812 B.n421 B.n420 10.6151
R813 B.n421 B.n96 10.6151
R814 B.n425 B.n96 10.6151
R815 B.n426 B.n425 10.6151
R816 B.n427 B.n426 10.6151
R817 B.n427 B.n94 10.6151
R818 B.n431 B.n94 10.6151
R819 B.n432 B.n431 10.6151
R820 B.n433 B.n432 10.6151
R821 B.n433 B.n92 10.6151
R822 B.n437 B.n92 10.6151
R823 B.n438 B.n437 10.6151
R824 B.n439 B.n438 10.6151
R825 B.n439 B.n90 10.6151
R826 B.n443 B.n90 10.6151
R827 B.n444 B.n443 10.6151
R828 B.n445 B.n444 10.6151
R829 B.n445 B.n88 10.6151
R830 B.n449 B.n88 10.6151
R831 B.n450 B.n449 10.6151
R832 B.n451 B.n450 10.6151
R833 B.n451 B.n86 10.6151
R834 B.n455 B.n86 10.6151
R835 B.n456 B.n455 10.6151
R836 B.n457 B.n456 10.6151
R837 B.n457 B.n84 10.6151
R838 B.n461 B.n84 10.6151
R839 B.n462 B.n461 10.6151
R840 B.n463 B.n462 10.6151
R841 B.n463 B.n82 10.6151
R842 B.n467 B.n82 10.6151
R843 B.n468 B.n467 10.6151
R844 B.n469 B.n468 10.6151
R845 B.n469 B.n80 10.6151
R846 B.n473 B.n80 10.6151
R847 B.n474 B.n473 10.6151
R848 B.n475 B.n474 10.6151
R849 B.n475 B.n78 10.6151
R850 B.n479 B.n78 10.6151
R851 B.n480 B.n479 10.6151
R852 B.n481 B.n480 10.6151
R853 B.n481 B.n76 10.6151
R854 B.n485 B.n76 10.6151
R855 B.n486 B.n485 10.6151
R856 B.n487 B.n486 10.6151
R857 B.n487 B.n74 10.6151
R858 B.n491 B.n74 10.6151
R859 B.n492 B.n491 10.6151
R860 B.n493 B.n492 10.6151
R861 B.n493 B.n72 10.6151
R862 B.n497 B.n72 10.6151
R863 B.n498 B.n497 10.6151
R864 B.n499 B.n498 10.6151
R865 B.n499 B.n70 10.6151
R866 B.n503 B.n70 10.6151
R867 B.n504 B.n503 10.6151
R868 B.n505 B.n504 10.6151
R869 B.n505 B.n68 10.6151
R870 B.n509 B.n68 10.6151
R871 B.n510 B.n509 10.6151
R872 B.n511 B.n510 10.6151
R873 B.n511 B.n66 10.6151
R874 B.n515 B.n66 10.6151
R875 B.n516 B.n515 10.6151
R876 B.n259 B.n154 10.6151
R877 B.n263 B.n154 10.6151
R878 B.n264 B.n263 10.6151
R879 B.n265 B.n264 10.6151
R880 B.n265 B.n152 10.6151
R881 B.n269 B.n152 10.6151
R882 B.n270 B.n269 10.6151
R883 B.n271 B.n270 10.6151
R884 B.n271 B.n150 10.6151
R885 B.n275 B.n150 10.6151
R886 B.n276 B.n275 10.6151
R887 B.n277 B.n276 10.6151
R888 B.n277 B.n148 10.6151
R889 B.n281 B.n148 10.6151
R890 B.n282 B.n281 10.6151
R891 B.n283 B.n282 10.6151
R892 B.n283 B.n146 10.6151
R893 B.n287 B.n146 10.6151
R894 B.n288 B.n287 10.6151
R895 B.n289 B.n288 10.6151
R896 B.n289 B.n144 10.6151
R897 B.n293 B.n144 10.6151
R898 B.n294 B.n293 10.6151
R899 B.n295 B.n294 10.6151
R900 B.n295 B.n142 10.6151
R901 B.n299 B.n142 10.6151
R902 B.n302 B.n301 10.6151
R903 B.n302 B.n138 10.6151
R904 B.n306 B.n138 10.6151
R905 B.n307 B.n306 10.6151
R906 B.n308 B.n307 10.6151
R907 B.n308 B.n136 10.6151
R908 B.n312 B.n136 10.6151
R909 B.n313 B.n312 10.6151
R910 B.n314 B.n313 10.6151
R911 B.n318 B.n317 10.6151
R912 B.n319 B.n318 10.6151
R913 B.n319 B.n130 10.6151
R914 B.n323 B.n130 10.6151
R915 B.n324 B.n323 10.6151
R916 B.n325 B.n324 10.6151
R917 B.n325 B.n128 10.6151
R918 B.n329 B.n128 10.6151
R919 B.n330 B.n329 10.6151
R920 B.n331 B.n330 10.6151
R921 B.n331 B.n126 10.6151
R922 B.n335 B.n126 10.6151
R923 B.n336 B.n335 10.6151
R924 B.n337 B.n336 10.6151
R925 B.n337 B.n124 10.6151
R926 B.n341 B.n124 10.6151
R927 B.n342 B.n341 10.6151
R928 B.n343 B.n342 10.6151
R929 B.n343 B.n122 10.6151
R930 B.n347 B.n122 10.6151
R931 B.n348 B.n347 10.6151
R932 B.n349 B.n348 10.6151
R933 B.n349 B.n120 10.6151
R934 B.n353 B.n120 10.6151
R935 B.n354 B.n353 10.6151
R936 B.n355 B.n354 10.6151
R937 B.n258 B.n257 10.6151
R938 B.n257 B.n156 10.6151
R939 B.n253 B.n156 10.6151
R940 B.n253 B.n252 10.6151
R941 B.n252 B.n251 10.6151
R942 B.n251 B.n158 10.6151
R943 B.n247 B.n158 10.6151
R944 B.n247 B.n246 10.6151
R945 B.n246 B.n245 10.6151
R946 B.n245 B.n160 10.6151
R947 B.n241 B.n160 10.6151
R948 B.n241 B.n240 10.6151
R949 B.n240 B.n239 10.6151
R950 B.n239 B.n162 10.6151
R951 B.n235 B.n162 10.6151
R952 B.n235 B.n234 10.6151
R953 B.n234 B.n233 10.6151
R954 B.n233 B.n164 10.6151
R955 B.n229 B.n164 10.6151
R956 B.n229 B.n228 10.6151
R957 B.n228 B.n227 10.6151
R958 B.n227 B.n166 10.6151
R959 B.n223 B.n166 10.6151
R960 B.n223 B.n222 10.6151
R961 B.n222 B.n221 10.6151
R962 B.n221 B.n168 10.6151
R963 B.n217 B.n168 10.6151
R964 B.n217 B.n216 10.6151
R965 B.n216 B.n215 10.6151
R966 B.n215 B.n170 10.6151
R967 B.n211 B.n170 10.6151
R968 B.n211 B.n210 10.6151
R969 B.n210 B.n209 10.6151
R970 B.n209 B.n172 10.6151
R971 B.n205 B.n172 10.6151
R972 B.n205 B.n204 10.6151
R973 B.n204 B.n203 10.6151
R974 B.n203 B.n174 10.6151
R975 B.n199 B.n174 10.6151
R976 B.n199 B.n198 10.6151
R977 B.n198 B.n197 10.6151
R978 B.n197 B.n176 10.6151
R979 B.n193 B.n176 10.6151
R980 B.n193 B.n192 10.6151
R981 B.n192 B.n191 10.6151
R982 B.n191 B.n178 10.6151
R983 B.n187 B.n178 10.6151
R984 B.n187 B.n186 10.6151
R985 B.n186 B.n185 10.6151
R986 B.n185 B.n180 10.6151
R987 B.n181 B.n180 10.6151
R988 B.n181 B.n0 10.6151
R989 B.n691 B.n1 10.6151
R990 B.n691 B.n690 10.6151
R991 B.n690 B.n689 10.6151
R992 B.n689 B.n4 10.6151
R993 B.n685 B.n4 10.6151
R994 B.n685 B.n684 10.6151
R995 B.n684 B.n683 10.6151
R996 B.n683 B.n6 10.6151
R997 B.n679 B.n6 10.6151
R998 B.n679 B.n678 10.6151
R999 B.n678 B.n677 10.6151
R1000 B.n677 B.n8 10.6151
R1001 B.n673 B.n8 10.6151
R1002 B.n673 B.n672 10.6151
R1003 B.n672 B.n671 10.6151
R1004 B.n671 B.n10 10.6151
R1005 B.n667 B.n10 10.6151
R1006 B.n667 B.n666 10.6151
R1007 B.n666 B.n665 10.6151
R1008 B.n665 B.n12 10.6151
R1009 B.n661 B.n12 10.6151
R1010 B.n661 B.n660 10.6151
R1011 B.n660 B.n659 10.6151
R1012 B.n659 B.n14 10.6151
R1013 B.n655 B.n14 10.6151
R1014 B.n655 B.n654 10.6151
R1015 B.n654 B.n653 10.6151
R1016 B.n653 B.n16 10.6151
R1017 B.n649 B.n16 10.6151
R1018 B.n649 B.n648 10.6151
R1019 B.n648 B.n647 10.6151
R1020 B.n647 B.n18 10.6151
R1021 B.n643 B.n18 10.6151
R1022 B.n643 B.n642 10.6151
R1023 B.n642 B.n641 10.6151
R1024 B.n641 B.n20 10.6151
R1025 B.n637 B.n20 10.6151
R1026 B.n637 B.n636 10.6151
R1027 B.n636 B.n635 10.6151
R1028 B.n635 B.n22 10.6151
R1029 B.n631 B.n22 10.6151
R1030 B.n631 B.n630 10.6151
R1031 B.n630 B.n629 10.6151
R1032 B.n629 B.n24 10.6151
R1033 B.n625 B.n24 10.6151
R1034 B.n625 B.n624 10.6151
R1035 B.n624 B.n623 10.6151
R1036 B.n623 B.n26 10.6151
R1037 B.n619 B.n26 10.6151
R1038 B.n619 B.n618 10.6151
R1039 B.n618 B.n617 10.6151
R1040 B.n617 B.n28 10.6151
R1041 B.n575 B.n44 9.36635
R1042 B.n558 B.n557 9.36635
R1043 B.n300 B.n299 9.36635
R1044 B.n317 B.n134 9.36635
R1045 B.n695 B.n0 2.81026
R1046 B.n695 B.n1 2.81026
R1047 B.n572 B.n44 1.24928
R1048 B.n559 B.n558 1.24928
R1049 B.n301 B.n300 1.24928
R1050 B.n314 B.n134 1.24928
R1051 VP.n16 VP.n15 161.3
R1052 VP.n17 VP.n12 161.3
R1053 VP.n19 VP.n18 161.3
R1054 VP.n20 VP.n11 161.3
R1055 VP.n22 VP.n21 161.3
R1056 VP.n23 VP.n10 161.3
R1057 VP.n25 VP.n24 161.3
R1058 VP.n50 VP.n49 161.3
R1059 VP.n48 VP.n1 161.3
R1060 VP.n47 VP.n46 161.3
R1061 VP.n45 VP.n2 161.3
R1062 VP.n44 VP.n43 161.3
R1063 VP.n42 VP.n3 161.3
R1064 VP.n41 VP.n40 161.3
R1065 VP.n39 VP.n4 161.3
R1066 VP.n38 VP.n37 161.3
R1067 VP.n36 VP.n5 161.3
R1068 VP.n35 VP.n34 161.3
R1069 VP.n33 VP.n6 161.3
R1070 VP.n32 VP.n31 161.3
R1071 VP.n30 VP.n7 161.3
R1072 VP.n29 VP.n28 161.3
R1073 VP.n14 VP.t2 83.9337
R1074 VP.n27 VP.n8 74.9986
R1075 VP.n51 VP.n0 74.9986
R1076 VP.n26 VP.n9 74.9986
R1077 VP.n14 VP.n13 50.3132
R1078 VP.n35 VP.n6 49.7803
R1079 VP.n43 VP.n2 49.7803
R1080 VP.n18 VP.n11 49.7803
R1081 VP.n4 VP.t1 49.7241
R1082 VP.n8 VP.t3 49.7241
R1083 VP.n0 VP.t5 49.7241
R1084 VP.n13 VP.t0 49.7241
R1085 VP.n9 VP.t4 49.7241
R1086 VP.n27 VP.n26 48.6397
R1087 VP.n31 VP.n6 31.3737
R1088 VP.n47 VP.n2 31.3737
R1089 VP.n22 VP.n11 31.3737
R1090 VP.n30 VP.n29 24.5923
R1091 VP.n31 VP.n30 24.5923
R1092 VP.n36 VP.n35 24.5923
R1093 VP.n37 VP.n36 24.5923
R1094 VP.n37 VP.n4 24.5923
R1095 VP.n41 VP.n4 24.5923
R1096 VP.n42 VP.n41 24.5923
R1097 VP.n43 VP.n42 24.5923
R1098 VP.n48 VP.n47 24.5923
R1099 VP.n49 VP.n48 24.5923
R1100 VP.n23 VP.n22 24.5923
R1101 VP.n24 VP.n23 24.5923
R1102 VP.n16 VP.n13 24.5923
R1103 VP.n17 VP.n16 24.5923
R1104 VP.n18 VP.n17 24.5923
R1105 VP.n29 VP.n8 15.2474
R1106 VP.n49 VP.n0 15.2474
R1107 VP.n24 VP.n9 15.2474
R1108 VP.n15 VP.n14 2.96487
R1109 VP.n26 VP.n25 0.354861
R1110 VP.n28 VP.n27 0.354861
R1111 VP.n51 VP.n50 0.354861
R1112 VP VP.n51 0.267071
R1113 VP.n15 VP.n12 0.189894
R1114 VP.n19 VP.n12 0.189894
R1115 VP.n20 VP.n19 0.189894
R1116 VP.n21 VP.n20 0.189894
R1117 VP.n21 VP.n10 0.189894
R1118 VP.n25 VP.n10 0.189894
R1119 VP.n28 VP.n7 0.189894
R1120 VP.n32 VP.n7 0.189894
R1121 VP.n33 VP.n32 0.189894
R1122 VP.n34 VP.n33 0.189894
R1123 VP.n34 VP.n5 0.189894
R1124 VP.n38 VP.n5 0.189894
R1125 VP.n39 VP.n38 0.189894
R1126 VP.n40 VP.n39 0.189894
R1127 VP.n40 VP.n3 0.189894
R1128 VP.n44 VP.n3 0.189894
R1129 VP.n45 VP.n44 0.189894
R1130 VP.n46 VP.n45 0.189894
R1131 VP.n46 VP.n1 0.189894
R1132 VP.n50 VP.n1 0.189894
R1133 VDD1.n31 VDD1.n30 585
R1134 VDD1.n29 VDD1.n28 585
R1135 VDD1.n4 VDD1.n3 585
R1136 VDD1.n23 VDD1.n22 585
R1137 VDD1.n21 VDD1.n20 585
R1138 VDD1.n8 VDD1.n7 585
R1139 VDD1.n15 VDD1.n14 585
R1140 VDD1.n13 VDD1.n12 585
R1141 VDD1.n48 VDD1.n47 585
R1142 VDD1.n50 VDD1.n49 585
R1143 VDD1.n43 VDD1.n42 585
R1144 VDD1.n56 VDD1.n55 585
R1145 VDD1.n58 VDD1.n57 585
R1146 VDD1.n39 VDD1.n38 585
R1147 VDD1.n64 VDD1.n63 585
R1148 VDD1.n66 VDD1.n65 585
R1149 VDD1.n30 VDD1.n0 498.474
R1150 VDD1.n65 VDD1.n35 498.474
R1151 VDD1.n11 VDD1.t5 329.053
R1152 VDD1.n46 VDD1.t4 329.053
R1153 VDD1.n30 VDD1.n29 171.744
R1154 VDD1.n29 VDD1.n3 171.744
R1155 VDD1.n22 VDD1.n3 171.744
R1156 VDD1.n22 VDD1.n21 171.744
R1157 VDD1.n21 VDD1.n7 171.744
R1158 VDD1.n14 VDD1.n7 171.744
R1159 VDD1.n14 VDD1.n13 171.744
R1160 VDD1.n49 VDD1.n48 171.744
R1161 VDD1.n49 VDD1.n42 171.744
R1162 VDD1.n56 VDD1.n42 171.744
R1163 VDD1.n57 VDD1.n56 171.744
R1164 VDD1.n57 VDD1.n38 171.744
R1165 VDD1.n64 VDD1.n38 171.744
R1166 VDD1.n65 VDD1.n64 171.744
R1167 VDD1.n71 VDD1.n70 87.5439
R1168 VDD1.n73 VDD1.n72 86.7781
R1169 VDD1.n13 VDD1.t5 85.8723
R1170 VDD1.n48 VDD1.t4 85.8723
R1171 VDD1 VDD1.n34 53.3251
R1172 VDD1.n71 VDD1.n69 53.2115
R1173 VDD1.n73 VDD1.n71 42.8048
R1174 VDD1.n32 VDD1.n31 12.8005
R1175 VDD1.n67 VDD1.n66 12.8005
R1176 VDD1.n28 VDD1.n2 12.0247
R1177 VDD1.n63 VDD1.n37 12.0247
R1178 VDD1.n27 VDD1.n4 11.249
R1179 VDD1.n62 VDD1.n39 11.249
R1180 VDD1.n12 VDD1.n11 10.7237
R1181 VDD1.n47 VDD1.n46 10.7237
R1182 VDD1.n24 VDD1.n23 10.4732
R1183 VDD1.n59 VDD1.n58 10.4732
R1184 VDD1.n20 VDD1.n6 9.69747
R1185 VDD1.n55 VDD1.n41 9.69747
R1186 VDD1.n34 VDD1.n33 9.45567
R1187 VDD1.n69 VDD1.n68 9.45567
R1188 VDD1.n10 VDD1.n9 9.3005
R1189 VDD1.n17 VDD1.n16 9.3005
R1190 VDD1.n19 VDD1.n18 9.3005
R1191 VDD1.n6 VDD1.n5 9.3005
R1192 VDD1.n25 VDD1.n24 9.3005
R1193 VDD1.n27 VDD1.n26 9.3005
R1194 VDD1.n2 VDD1.n1 9.3005
R1195 VDD1.n33 VDD1.n32 9.3005
R1196 VDD1.n45 VDD1.n44 9.3005
R1197 VDD1.n52 VDD1.n51 9.3005
R1198 VDD1.n54 VDD1.n53 9.3005
R1199 VDD1.n41 VDD1.n40 9.3005
R1200 VDD1.n60 VDD1.n59 9.3005
R1201 VDD1.n62 VDD1.n61 9.3005
R1202 VDD1.n37 VDD1.n36 9.3005
R1203 VDD1.n68 VDD1.n67 9.3005
R1204 VDD1.n19 VDD1.n8 8.92171
R1205 VDD1.n54 VDD1.n43 8.92171
R1206 VDD1.n16 VDD1.n15 8.14595
R1207 VDD1.n51 VDD1.n50 8.14595
R1208 VDD1.n34 VDD1.n0 7.75445
R1209 VDD1.n69 VDD1.n35 7.75445
R1210 VDD1.n12 VDD1.n10 7.3702
R1211 VDD1.n47 VDD1.n45 7.3702
R1212 VDD1.n32 VDD1.n0 6.08283
R1213 VDD1.n67 VDD1.n35 6.08283
R1214 VDD1.n15 VDD1.n10 5.81868
R1215 VDD1.n50 VDD1.n45 5.81868
R1216 VDD1.n16 VDD1.n8 5.04292
R1217 VDD1.n51 VDD1.n43 5.04292
R1218 VDD1.n72 VDD1.t1 4.52766
R1219 VDD1.n72 VDD1.t3 4.52766
R1220 VDD1.n70 VDD1.t0 4.52766
R1221 VDD1.n70 VDD1.t2 4.52766
R1222 VDD1.n20 VDD1.n19 4.26717
R1223 VDD1.n55 VDD1.n54 4.26717
R1224 VDD1.n23 VDD1.n6 3.49141
R1225 VDD1.n58 VDD1.n41 3.49141
R1226 VDD1.n24 VDD1.n4 2.71565
R1227 VDD1.n59 VDD1.n39 2.71565
R1228 VDD1.n11 VDD1.n9 2.41305
R1229 VDD1.n46 VDD1.n44 2.41305
R1230 VDD1.n28 VDD1.n27 1.93989
R1231 VDD1.n63 VDD1.n62 1.93989
R1232 VDD1.n31 VDD1.n2 1.16414
R1233 VDD1.n66 VDD1.n37 1.16414
R1234 VDD1 VDD1.n73 0.763431
R1235 VDD1.n33 VDD1.n1 0.155672
R1236 VDD1.n26 VDD1.n1 0.155672
R1237 VDD1.n26 VDD1.n25 0.155672
R1238 VDD1.n25 VDD1.n5 0.155672
R1239 VDD1.n18 VDD1.n5 0.155672
R1240 VDD1.n18 VDD1.n17 0.155672
R1241 VDD1.n17 VDD1.n9 0.155672
R1242 VDD1.n52 VDD1.n44 0.155672
R1243 VDD1.n53 VDD1.n52 0.155672
R1244 VDD1.n53 VDD1.n40 0.155672
R1245 VDD1.n60 VDD1.n40 0.155672
R1246 VDD1.n61 VDD1.n60 0.155672
R1247 VDD1.n61 VDD1.n36 0.155672
R1248 VDD1.n68 VDD1.n36 0.155672
R1249 VTAIL.n129 VTAIL.n128 585
R1250 VTAIL.n131 VTAIL.n130 585
R1251 VTAIL.n124 VTAIL.n123 585
R1252 VTAIL.n137 VTAIL.n136 585
R1253 VTAIL.n139 VTAIL.n138 585
R1254 VTAIL.n120 VTAIL.n119 585
R1255 VTAIL.n145 VTAIL.n144 585
R1256 VTAIL.n147 VTAIL.n146 585
R1257 VTAIL.n15 VTAIL.n14 585
R1258 VTAIL.n17 VTAIL.n16 585
R1259 VTAIL.n10 VTAIL.n9 585
R1260 VTAIL.n23 VTAIL.n22 585
R1261 VTAIL.n25 VTAIL.n24 585
R1262 VTAIL.n6 VTAIL.n5 585
R1263 VTAIL.n31 VTAIL.n30 585
R1264 VTAIL.n33 VTAIL.n32 585
R1265 VTAIL.n111 VTAIL.n110 585
R1266 VTAIL.n109 VTAIL.n108 585
R1267 VTAIL.n84 VTAIL.n83 585
R1268 VTAIL.n103 VTAIL.n102 585
R1269 VTAIL.n101 VTAIL.n100 585
R1270 VTAIL.n88 VTAIL.n87 585
R1271 VTAIL.n95 VTAIL.n94 585
R1272 VTAIL.n93 VTAIL.n92 585
R1273 VTAIL.n73 VTAIL.n72 585
R1274 VTAIL.n71 VTAIL.n70 585
R1275 VTAIL.n46 VTAIL.n45 585
R1276 VTAIL.n65 VTAIL.n64 585
R1277 VTAIL.n63 VTAIL.n62 585
R1278 VTAIL.n50 VTAIL.n49 585
R1279 VTAIL.n57 VTAIL.n56 585
R1280 VTAIL.n55 VTAIL.n54 585
R1281 VTAIL.n146 VTAIL.n116 498.474
R1282 VTAIL.n32 VTAIL.n2 498.474
R1283 VTAIL.n110 VTAIL.n80 498.474
R1284 VTAIL.n72 VTAIL.n42 498.474
R1285 VTAIL.n127 VTAIL.t4 329.053
R1286 VTAIL.n13 VTAIL.t6 329.053
R1287 VTAIL.n91 VTAIL.t7 329.053
R1288 VTAIL.n53 VTAIL.t0 329.053
R1289 VTAIL.n130 VTAIL.n129 171.744
R1290 VTAIL.n130 VTAIL.n123 171.744
R1291 VTAIL.n137 VTAIL.n123 171.744
R1292 VTAIL.n138 VTAIL.n137 171.744
R1293 VTAIL.n138 VTAIL.n119 171.744
R1294 VTAIL.n145 VTAIL.n119 171.744
R1295 VTAIL.n146 VTAIL.n145 171.744
R1296 VTAIL.n16 VTAIL.n15 171.744
R1297 VTAIL.n16 VTAIL.n9 171.744
R1298 VTAIL.n23 VTAIL.n9 171.744
R1299 VTAIL.n24 VTAIL.n23 171.744
R1300 VTAIL.n24 VTAIL.n5 171.744
R1301 VTAIL.n31 VTAIL.n5 171.744
R1302 VTAIL.n32 VTAIL.n31 171.744
R1303 VTAIL.n110 VTAIL.n109 171.744
R1304 VTAIL.n109 VTAIL.n83 171.744
R1305 VTAIL.n102 VTAIL.n83 171.744
R1306 VTAIL.n102 VTAIL.n101 171.744
R1307 VTAIL.n101 VTAIL.n87 171.744
R1308 VTAIL.n94 VTAIL.n87 171.744
R1309 VTAIL.n94 VTAIL.n93 171.744
R1310 VTAIL.n72 VTAIL.n71 171.744
R1311 VTAIL.n71 VTAIL.n45 171.744
R1312 VTAIL.n64 VTAIL.n45 171.744
R1313 VTAIL.n64 VTAIL.n63 171.744
R1314 VTAIL.n63 VTAIL.n49 171.744
R1315 VTAIL.n56 VTAIL.n49 171.744
R1316 VTAIL.n56 VTAIL.n55 171.744
R1317 VTAIL.n129 VTAIL.t4 85.8723
R1318 VTAIL.n15 VTAIL.t6 85.8723
R1319 VTAIL.n93 VTAIL.t7 85.8723
R1320 VTAIL.n55 VTAIL.t0 85.8723
R1321 VTAIL.n79 VTAIL.n78 70.0994
R1322 VTAIL.n41 VTAIL.n40 70.0994
R1323 VTAIL.n1 VTAIL.n0 70.0993
R1324 VTAIL.n39 VTAIL.n38 70.0993
R1325 VTAIL.n151 VTAIL.n150 34.1247
R1326 VTAIL.n37 VTAIL.n36 34.1247
R1327 VTAIL.n115 VTAIL.n114 34.1247
R1328 VTAIL.n77 VTAIL.n76 34.1247
R1329 VTAIL.n41 VTAIL.n39 25.1255
R1330 VTAIL.n151 VTAIL.n115 21.841
R1331 VTAIL.n148 VTAIL.n147 12.8005
R1332 VTAIL.n34 VTAIL.n33 12.8005
R1333 VTAIL.n112 VTAIL.n111 12.8005
R1334 VTAIL.n74 VTAIL.n73 12.8005
R1335 VTAIL.n144 VTAIL.n118 12.0247
R1336 VTAIL.n30 VTAIL.n4 12.0247
R1337 VTAIL.n108 VTAIL.n82 12.0247
R1338 VTAIL.n70 VTAIL.n44 12.0247
R1339 VTAIL.n143 VTAIL.n120 11.249
R1340 VTAIL.n29 VTAIL.n6 11.249
R1341 VTAIL.n107 VTAIL.n84 11.249
R1342 VTAIL.n69 VTAIL.n46 11.249
R1343 VTAIL.n128 VTAIL.n127 10.7237
R1344 VTAIL.n14 VTAIL.n13 10.7237
R1345 VTAIL.n92 VTAIL.n91 10.7237
R1346 VTAIL.n54 VTAIL.n53 10.7237
R1347 VTAIL.n140 VTAIL.n139 10.4732
R1348 VTAIL.n26 VTAIL.n25 10.4732
R1349 VTAIL.n104 VTAIL.n103 10.4732
R1350 VTAIL.n66 VTAIL.n65 10.4732
R1351 VTAIL.n136 VTAIL.n122 9.69747
R1352 VTAIL.n22 VTAIL.n8 9.69747
R1353 VTAIL.n100 VTAIL.n86 9.69747
R1354 VTAIL.n62 VTAIL.n48 9.69747
R1355 VTAIL.n150 VTAIL.n149 9.45567
R1356 VTAIL.n36 VTAIL.n35 9.45567
R1357 VTAIL.n114 VTAIL.n113 9.45567
R1358 VTAIL.n76 VTAIL.n75 9.45567
R1359 VTAIL.n126 VTAIL.n125 9.3005
R1360 VTAIL.n133 VTAIL.n132 9.3005
R1361 VTAIL.n135 VTAIL.n134 9.3005
R1362 VTAIL.n122 VTAIL.n121 9.3005
R1363 VTAIL.n141 VTAIL.n140 9.3005
R1364 VTAIL.n143 VTAIL.n142 9.3005
R1365 VTAIL.n118 VTAIL.n117 9.3005
R1366 VTAIL.n149 VTAIL.n148 9.3005
R1367 VTAIL.n12 VTAIL.n11 9.3005
R1368 VTAIL.n19 VTAIL.n18 9.3005
R1369 VTAIL.n21 VTAIL.n20 9.3005
R1370 VTAIL.n8 VTAIL.n7 9.3005
R1371 VTAIL.n27 VTAIL.n26 9.3005
R1372 VTAIL.n29 VTAIL.n28 9.3005
R1373 VTAIL.n4 VTAIL.n3 9.3005
R1374 VTAIL.n35 VTAIL.n34 9.3005
R1375 VTAIL.n90 VTAIL.n89 9.3005
R1376 VTAIL.n97 VTAIL.n96 9.3005
R1377 VTAIL.n99 VTAIL.n98 9.3005
R1378 VTAIL.n86 VTAIL.n85 9.3005
R1379 VTAIL.n105 VTAIL.n104 9.3005
R1380 VTAIL.n107 VTAIL.n106 9.3005
R1381 VTAIL.n82 VTAIL.n81 9.3005
R1382 VTAIL.n113 VTAIL.n112 9.3005
R1383 VTAIL.n52 VTAIL.n51 9.3005
R1384 VTAIL.n59 VTAIL.n58 9.3005
R1385 VTAIL.n61 VTAIL.n60 9.3005
R1386 VTAIL.n48 VTAIL.n47 9.3005
R1387 VTAIL.n67 VTAIL.n66 9.3005
R1388 VTAIL.n69 VTAIL.n68 9.3005
R1389 VTAIL.n44 VTAIL.n43 9.3005
R1390 VTAIL.n75 VTAIL.n74 9.3005
R1391 VTAIL.n135 VTAIL.n124 8.92171
R1392 VTAIL.n21 VTAIL.n10 8.92171
R1393 VTAIL.n99 VTAIL.n88 8.92171
R1394 VTAIL.n61 VTAIL.n50 8.92171
R1395 VTAIL.n132 VTAIL.n131 8.14595
R1396 VTAIL.n18 VTAIL.n17 8.14595
R1397 VTAIL.n96 VTAIL.n95 8.14595
R1398 VTAIL.n58 VTAIL.n57 8.14595
R1399 VTAIL.n150 VTAIL.n116 7.75445
R1400 VTAIL.n36 VTAIL.n2 7.75445
R1401 VTAIL.n114 VTAIL.n80 7.75445
R1402 VTAIL.n76 VTAIL.n42 7.75445
R1403 VTAIL.n128 VTAIL.n126 7.3702
R1404 VTAIL.n14 VTAIL.n12 7.3702
R1405 VTAIL.n92 VTAIL.n90 7.3702
R1406 VTAIL.n54 VTAIL.n52 7.3702
R1407 VTAIL.n148 VTAIL.n116 6.08283
R1408 VTAIL.n34 VTAIL.n2 6.08283
R1409 VTAIL.n112 VTAIL.n80 6.08283
R1410 VTAIL.n74 VTAIL.n42 6.08283
R1411 VTAIL.n131 VTAIL.n126 5.81868
R1412 VTAIL.n17 VTAIL.n12 5.81868
R1413 VTAIL.n95 VTAIL.n90 5.81868
R1414 VTAIL.n57 VTAIL.n52 5.81868
R1415 VTAIL.n132 VTAIL.n124 5.04292
R1416 VTAIL.n18 VTAIL.n10 5.04292
R1417 VTAIL.n96 VTAIL.n88 5.04292
R1418 VTAIL.n58 VTAIL.n50 5.04292
R1419 VTAIL.n0 VTAIL.t1 4.52766
R1420 VTAIL.n0 VTAIL.t3 4.52766
R1421 VTAIL.n38 VTAIL.t8 4.52766
R1422 VTAIL.n38 VTAIL.t10 4.52766
R1423 VTAIL.n78 VTAIL.t9 4.52766
R1424 VTAIL.n78 VTAIL.t11 4.52766
R1425 VTAIL.n40 VTAIL.t2 4.52766
R1426 VTAIL.n40 VTAIL.t5 4.52766
R1427 VTAIL.n136 VTAIL.n135 4.26717
R1428 VTAIL.n22 VTAIL.n21 4.26717
R1429 VTAIL.n100 VTAIL.n99 4.26717
R1430 VTAIL.n62 VTAIL.n61 4.26717
R1431 VTAIL.n139 VTAIL.n122 3.49141
R1432 VTAIL.n25 VTAIL.n8 3.49141
R1433 VTAIL.n103 VTAIL.n86 3.49141
R1434 VTAIL.n65 VTAIL.n48 3.49141
R1435 VTAIL.n77 VTAIL.n41 3.28498
R1436 VTAIL.n115 VTAIL.n79 3.28498
R1437 VTAIL.n39 VTAIL.n37 3.28498
R1438 VTAIL.n140 VTAIL.n120 2.71565
R1439 VTAIL.n26 VTAIL.n6 2.71565
R1440 VTAIL.n104 VTAIL.n84 2.71565
R1441 VTAIL.n66 VTAIL.n46 2.71565
R1442 VTAIL.n127 VTAIL.n125 2.41305
R1443 VTAIL.n13 VTAIL.n11 2.41305
R1444 VTAIL.n91 VTAIL.n89 2.41305
R1445 VTAIL.n53 VTAIL.n51 2.41305
R1446 VTAIL VTAIL.n151 2.40567
R1447 VTAIL.n79 VTAIL.n77 2.11257
R1448 VTAIL.n37 VTAIL.n1 2.11257
R1449 VTAIL.n144 VTAIL.n143 1.93989
R1450 VTAIL.n30 VTAIL.n29 1.93989
R1451 VTAIL.n108 VTAIL.n107 1.93989
R1452 VTAIL.n70 VTAIL.n69 1.93989
R1453 VTAIL.n147 VTAIL.n118 1.16414
R1454 VTAIL.n33 VTAIL.n4 1.16414
R1455 VTAIL.n111 VTAIL.n82 1.16414
R1456 VTAIL.n73 VTAIL.n44 1.16414
R1457 VTAIL VTAIL.n1 0.87981
R1458 VTAIL.n133 VTAIL.n125 0.155672
R1459 VTAIL.n134 VTAIL.n133 0.155672
R1460 VTAIL.n134 VTAIL.n121 0.155672
R1461 VTAIL.n141 VTAIL.n121 0.155672
R1462 VTAIL.n142 VTAIL.n141 0.155672
R1463 VTAIL.n142 VTAIL.n117 0.155672
R1464 VTAIL.n149 VTAIL.n117 0.155672
R1465 VTAIL.n19 VTAIL.n11 0.155672
R1466 VTAIL.n20 VTAIL.n19 0.155672
R1467 VTAIL.n20 VTAIL.n7 0.155672
R1468 VTAIL.n27 VTAIL.n7 0.155672
R1469 VTAIL.n28 VTAIL.n27 0.155672
R1470 VTAIL.n28 VTAIL.n3 0.155672
R1471 VTAIL.n35 VTAIL.n3 0.155672
R1472 VTAIL.n113 VTAIL.n81 0.155672
R1473 VTAIL.n106 VTAIL.n81 0.155672
R1474 VTAIL.n106 VTAIL.n105 0.155672
R1475 VTAIL.n105 VTAIL.n85 0.155672
R1476 VTAIL.n98 VTAIL.n85 0.155672
R1477 VTAIL.n98 VTAIL.n97 0.155672
R1478 VTAIL.n97 VTAIL.n89 0.155672
R1479 VTAIL.n75 VTAIL.n43 0.155672
R1480 VTAIL.n68 VTAIL.n43 0.155672
R1481 VTAIL.n68 VTAIL.n67 0.155672
R1482 VTAIL.n67 VTAIL.n47 0.155672
R1483 VTAIL.n60 VTAIL.n47 0.155672
R1484 VTAIL.n60 VTAIL.n59 0.155672
R1485 VTAIL.n59 VTAIL.n51 0.155672
R1486 VN.n34 VN.n33 161.3
R1487 VN.n32 VN.n19 161.3
R1488 VN.n31 VN.n30 161.3
R1489 VN.n29 VN.n20 161.3
R1490 VN.n28 VN.n27 161.3
R1491 VN.n26 VN.n21 161.3
R1492 VN.n25 VN.n24 161.3
R1493 VN.n16 VN.n15 161.3
R1494 VN.n14 VN.n1 161.3
R1495 VN.n13 VN.n12 161.3
R1496 VN.n11 VN.n2 161.3
R1497 VN.n10 VN.n9 161.3
R1498 VN.n8 VN.n3 161.3
R1499 VN.n7 VN.n6 161.3
R1500 VN.n23 VN.t2 83.9339
R1501 VN.n5 VN.t5 83.9339
R1502 VN.n17 VN.n0 74.9986
R1503 VN.n35 VN.n18 74.9986
R1504 VN.n5 VN.n4 50.3132
R1505 VN.n23 VN.n22 50.3132
R1506 VN.n9 VN.n2 49.7803
R1507 VN.n27 VN.n20 49.7803
R1508 VN.n4 VN.t1 49.7241
R1509 VN.n0 VN.t4 49.7241
R1510 VN.n22 VN.t3 49.7241
R1511 VN.n18 VN.t0 49.7241
R1512 VN VN.n35 48.805
R1513 VN.n13 VN.n2 31.3737
R1514 VN.n31 VN.n20 31.3737
R1515 VN.n7 VN.n4 24.5923
R1516 VN.n8 VN.n7 24.5923
R1517 VN.n9 VN.n8 24.5923
R1518 VN.n14 VN.n13 24.5923
R1519 VN.n15 VN.n14 24.5923
R1520 VN.n27 VN.n26 24.5923
R1521 VN.n26 VN.n25 24.5923
R1522 VN.n25 VN.n22 24.5923
R1523 VN.n33 VN.n32 24.5923
R1524 VN.n32 VN.n31 24.5923
R1525 VN.n15 VN.n0 15.2474
R1526 VN.n33 VN.n18 15.2474
R1527 VN.n24 VN.n23 2.96489
R1528 VN.n6 VN.n5 2.96489
R1529 VN.n35 VN.n34 0.354861
R1530 VN.n17 VN.n16 0.354861
R1531 VN VN.n17 0.267071
R1532 VN.n34 VN.n19 0.189894
R1533 VN.n30 VN.n19 0.189894
R1534 VN.n30 VN.n29 0.189894
R1535 VN.n29 VN.n28 0.189894
R1536 VN.n28 VN.n21 0.189894
R1537 VN.n24 VN.n21 0.189894
R1538 VN.n6 VN.n3 0.189894
R1539 VN.n10 VN.n3 0.189894
R1540 VN.n11 VN.n10 0.189894
R1541 VN.n12 VN.n11 0.189894
R1542 VN.n12 VN.n1 0.189894
R1543 VN.n16 VN.n1 0.189894
R1544 VDD2.n68 VDD2.n67 585
R1545 VDD2.n66 VDD2.n65 585
R1546 VDD2.n41 VDD2.n40 585
R1547 VDD2.n60 VDD2.n59 585
R1548 VDD2.n58 VDD2.n57 585
R1549 VDD2.n45 VDD2.n44 585
R1550 VDD2.n52 VDD2.n51 585
R1551 VDD2.n50 VDD2.n49 585
R1552 VDD2.n13 VDD2.n12 585
R1553 VDD2.n15 VDD2.n14 585
R1554 VDD2.n8 VDD2.n7 585
R1555 VDD2.n21 VDD2.n20 585
R1556 VDD2.n23 VDD2.n22 585
R1557 VDD2.n4 VDD2.n3 585
R1558 VDD2.n29 VDD2.n28 585
R1559 VDD2.n31 VDD2.n30 585
R1560 VDD2.n67 VDD2.n37 498.474
R1561 VDD2.n30 VDD2.n0 498.474
R1562 VDD2.n48 VDD2.t5 329.053
R1563 VDD2.n11 VDD2.t0 329.053
R1564 VDD2.n67 VDD2.n66 171.744
R1565 VDD2.n66 VDD2.n40 171.744
R1566 VDD2.n59 VDD2.n40 171.744
R1567 VDD2.n59 VDD2.n58 171.744
R1568 VDD2.n58 VDD2.n44 171.744
R1569 VDD2.n51 VDD2.n44 171.744
R1570 VDD2.n51 VDD2.n50 171.744
R1571 VDD2.n14 VDD2.n13 171.744
R1572 VDD2.n14 VDD2.n7 171.744
R1573 VDD2.n21 VDD2.n7 171.744
R1574 VDD2.n22 VDD2.n21 171.744
R1575 VDD2.n22 VDD2.n3 171.744
R1576 VDD2.n29 VDD2.n3 171.744
R1577 VDD2.n30 VDD2.n29 171.744
R1578 VDD2.n36 VDD2.n35 87.5439
R1579 VDD2 VDD2.n73 87.541
R1580 VDD2.n50 VDD2.t5 85.8723
R1581 VDD2.n13 VDD2.t0 85.8723
R1582 VDD2.n36 VDD2.n34 53.2115
R1583 VDD2.n72 VDD2.n71 50.8035
R1584 VDD2.n72 VDD2.n36 40.5795
R1585 VDD2.n69 VDD2.n68 12.8005
R1586 VDD2.n32 VDD2.n31 12.8005
R1587 VDD2.n65 VDD2.n39 12.0247
R1588 VDD2.n28 VDD2.n2 12.0247
R1589 VDD2.n64 VDD2.n41 11.249
R1590 VDD2.n27 VDD2.n4 11.249
R1591 VDD2.n49 VDD2.n48 10.7237
R1592 VDD2.n12 VDD2.n11 10.7237
R1593 VDD2.n61 VDD2.n60 10.4732
R1594 VDD2.n24 VDD2.n23 10.4732
R1595 VDD2.n57 VDD2.n43 9.69747
R1596 VDD2.n20 VDD2.n6 9.69747
R1597 VDD2.n71 VDD2.n70 9.45567
R1598 VDD2.n34 VDD2.n33 9.45567
R1599 VDD2.n47 VDD2.n46 9.3005
R1600 VDD2.n54 VDD2.n53 9.3005
R1601 VDD2.n56 VDD2.n55 9.3005
R1602 VDD2.n43 VDD2.n42 9.3005
R1603 VDD2.n62 VDD2.n61 9.3005
R1604 VDD2.n64 VDD2.n63 9.3005
R1605 VDD2.n39 VDD2.n38 9.3005
R1606 VDD2.n70 VDD2.n69 9.3005
R1607 VDD2.n10 VDD2.n9 9.3005
R1608 VDD2.n17 VDD2.n16 9.3005
R1609 VDD2.n19 VDD2.n18 9.3005
R1610 VDD2.n6 VDD2.n5 9.3005
R1611 VDD2.n25 VDD2.n24 9.3005
R1612 VDD2.n27 VDD2.n26 9.3005
R1613 VDD2.n2 VDD2.n1 9.3005
R1614 VDD2.n33 VDD2.n32 9.3005
R1615 VDD2.n56 VDD2.n45 8.92171
R1616 VDD2.n19 VDD2.n8 8.92171
R1617 VDD2.n53 VDD2.n52 8.14595
R1618 VDD2.n16 VDD2.n15 8.14595
R1619 VDD2.n71 VDD2.n37 7.75445
R1620 VDD2.n34 VDD2.n0 7.75445
R1621 VDD2.n49 VDD2.n47 7.3702
R1622 VDD2.n12 VDD2.n10 7.3702
R1623 VDD2.n69 VDD2.n37 6.08283
R1624 VDD2.n32 VDD2.n0 6.08283
R1625 VDD2.n52 VDD2.n47 5.81868
R1626 VDD2.n15 VDD2.n10 5.81868
R1627 VDD2.n53 VDD2.n45 5.04292
R1628 VDD2.n16 VDD2.n8 5.04292
R1629 VDD2.n73 VDD2.t2 4.52766
R1630 VDD2.n73 VDD2.t3 4.52766
R1631 VDD2.n35 VDD2.t4 4.52766
R1632 VDD2.n35 VDD2.t1 4.52766
R1633 VDD2.n57 VDD2.n56 4.26717
R1634 VDD2.n20 VDD2.n19 4.26717
R1635 VDD2.n60 VDD2.n43 3.49141
R1636 VDD2.n23 VDD2.n6 3.49141
R1637 VDD2.n61 VDD2.n41 2.71565
R1638 VDD2.n24 VDD2.n4 2.71565
R1639 VDD2 VDD2.n72 2.52205
R1640 VDD2.n48 VDD2.n46 2.41305
R1641 VDD2.n11 VDD2.n9 2.41305
R1642 VDD2.n65 VDD2.n64 1.93989
R1643 VDD2.n28 VDD2.n27 1.93989
R1644 VDD2.n68 VDD2.n39 1.16414
R1645 VDD2.n31 VDD2.n2 1.16414
R1646 VDD2.n70 VDD2.n38 0.155672
R1647 VDD2.n63 VDD2.n38 0.155672
R1648 VDD2.n63 VDD2.n62 0.155672
R1649 VDD2.n62 VDD2.n42 0.155672
R1650 VDD2.n55 VDD2.n42 0.155672
R1651 VDD2.n55 VDD2.n54 0.155672
R1652 VDD2.n54 VDD2.n46 0.155672
R1653 VDD2.n17 VDD2.n9 0.155672
R1654 VDD2.n18 VDD2.n17 0.155672
R1655 VDD2.n18 VDD2.n5 0.155672
R1656 VDD2.n25 VDD2.n5 0.155672
R1657 VDD2.n26 VDD2.n25 0.155672
R1658 VDD2.n26 VDD2.n1 0.155672
R1659 VDD2.n33 VDD2.n1 0.155672
C0 VDD2 VTAIL 6.49388f
C1 VP VDD2 0.532937f
C2 B VTAIL 2.89004f
C3 VP B 2.17648f
C4 VN VTAIL 5.15567f
C5 VDD1 VTAIL 6.43556f
C6 VP VN 6.88112f
C7 VP VDD1 4.76214f
C8 VDD2 w_n4018_n2404# 2.28742f
C9 w_n4018_n2404# B 9.54269f
C10 w_n4018_n2404# VN 7.71874f
C11 w_n4018_n2404# VDD1 2.17422f
C12 VP VTAIL 5.16985f
C13 w_n4018_n2404# VTAIL 2.39684f
C14 VP w_n4018_n2404# 8.24067f
C15 VDD2 B 2.02998f
C16 VDD2 VN 4.38384f
C17 VDD2 VDD1 1.74962f
C18 B VN 1.30065f
C19 B VDD1 1.93478f
C20 VN VDD1 0.152237f
C21 VDD2 VSUBS 2.014889f
C22 VDD1 VSUBS 1.956715f
C23 VTAIL VSUBS 0.808794f
C24 VN VSUBS 6.46888f
C25 VP VSUBS 3.262168f
C26 B VSUBS 5.100217f
C27 w_n4018_n2404# VSUBS 0.120106p
C28 VDD2.n0 VSUBS 0.031878f
C29 VDD2.n1 VSUBS 0.03035f
C30 VDD2.n2 VSUBS 0.016309f
C31 VDD2.n3 VSUBS 0.038547f
C32 VDD2.n4 VSUBS 0.017268f
C33 VDD2.n5 VSUBS 0.03035f
C34 VDD2.n6 VSUBS 0.016309f
C35 VDD2.n7 VSUBS 0.038547f
C36 VDD2.n8 VSUBS 0.017268f
C37 VDD2.n9 VSUBS 0.84984f
C38 VDD2.n10 VSUBS 0.016309f
C39 VDD2.t0 VSUBS 0.082771f
C40 VDD2.n11 VSUBS 0.17304f
C41 VDD2.n12 VSUBS 0.028996f
C42 VDD2.n13 VSUBS 0.02891f
C43 VDD2.n14 VSUBS 0.038547f
C44 VDD2.n15 VSUBS 0.017268f
C45 VDD2.n16 VSUBS 0.016309f
C46 VDD2.n17 VSUBS 0.03035f
C47 VDD2.n18 VSUBS 0.03035f
C48 VDD2.n19 VSUBS 0.016309f
C49 VDD2.n20 VSUBS 0.017268f
C50 VDD2.n21 VSUBS 0.038547f
C51 VDD2.n22 VSUBS 0.038547f
C52 VDD2.n23 VSUBS 0.017268f
C53 VDD2.n24 VSUBS 0.016309f
C54 VDD2.n25 VSUBS 0.03035f
C55 VDD2.n26 VSUBS 0.03035f
C56 VDD2.n27 VSUBS 0.016309f
C57 VDD2.n28 VSUBS 0.017268f
C58 VDD2.n29 VSUBS 0.038547f
C59 VDD2.n30 VSUBS 0.094261f
C60 VDD2.n31 VSUBS 0.017268f
C61 VDD2.n32 VSUBS 0.032026f
C62 VDD2.n33 VSUBS 0.074297f
C63 VDD2.n34 VSUBS 0.10575f
C64 VDD2.t4 VSUBS 0.172199f
C65 VDD2.t1 VSUBS 0.172199f
C66 VDD2.n35 VSUBS 1.22438f
C67 VDD2.n36 VSUBS 3.60552f
C68 VDD2.n37 VSUBS 0.031878f
C69 VDD2.n38 VSUBS 0.03035f
C70 VDD2.n39 VSUBS 0.016309f
C71 VDD2.n40 VSUBS 0.038547f
C72 VDD2.n41 VSUBS 0.017268f
C73 VDD2.n42 VSUBS 0.03035f
C74 VDD2.n43 VSUBS 0.016309f
C75 VDD2.n44 VSUBS 0.038547f
C76 VDD2.n45 VSUBS 0.017268f
C77 VDD2.n46 VSUBS 0.84984f
C78 VDD2.n47 VSUBS 0.016309f
C79 VDD2.t5 VSUBS 0.082771f
C80 VDD2.n48 VSUBS 0.17304f
C81 VDD2.n49 VSUBS 0.028996f
C82 VDD2.n50 VSUBS 0.02891f
C83 VDD2.n51 VSUBS 0.038547f
C84 VDD2.n52 VSUBS 0.017268f
C85 VDD2.n53 VSUBS 0.016309f
C86 VDD2.n54 VSUBS 0.03035f
C87 VDD2.n55 VSUBS 0.03035f
C88 VDD2.n56 VSUBS 0.016309f
C89 VDD2.n57 VSUBS 0.017268f
C90 VDD2.n58 VSUBS 0.038547f
C91 VDD2.n59 VSUBS 0.038547f
C92 VDD2.n60 VSUBS 0.017268f
C93 VDD2.n61 VSUBS 0.016309f
C94 VDD2.n62 VSUBS 0.03035f
C95 VDD2.n63 VSUBS 0.03035f
C96 VDD2.n64 VSUBS 0.016309f
C97 VDD2.n65 VSUBS 0.017268f
C98 VDD2.n66 VSUBS 0.038547f
C99 VDD2.n67 VSUBS 0.094261f
C100 VDD2.n68 VSUBS 0.017268f
C101 VDD2.n69 VSUBS 0.032026f
C102 VDD2.n70 VSUBS 0.074297f
C103 VDD2.n71 VSUBS 0.092328f
C104 VDD2.n72 VSUBS 2.94941f
C105 VDD2.t2 VSUBS 0.172199f
C106 VDD2.t3 VSUBS 0.172199f
C107 VDD2.n73 VSUBS 1.22434f
C108 VN.t4 VSUBS 2.11084f
C109 VN.n0 VSUBS 0.897545f
C110 VN.n1 VSUBS 0.031612f
C111 VN.n2 VSUBS 0.029367f
C112 VN.n3 VSUBS 0.031612f
C113 VN.t1 VSUBS 2.11084f
C114 VN.n4 VSUBS 0.891973f
C115 VN.t5 VSUBS 2.52136f
C116 VN.n5 VSUBS 0.8329f
C117 VN.n6 VSUBS 0.385625f
C118 VN.n7 VSUBS 0.058622f
C119 VN.n8 VSUBS 0.058622f
C120 VN.n9 VSUBS 0.058036f
C121 VN.n10 VSUBS 0.031612f
C122 VN.n11 VSUBS 0.031612f
C123 VN.n12 VSUBS 0.031612f
C124 VN.n13 VSUBS 0.063126f
C125 VN.n14 VSUBS 0.058622f
C126 VN.n15 VSUBS 0.047625f
C127 VN.n16 VSUBS 0.051014f
C128 VN.n17 VSUBS 0.078086f
C129 VN.t0 VSUBS 2.11084f
C130 VN.n18 VSUBS 0.897545f
C131 VN.n19 VSUBS 0.031612f
C132 VN.n20 VSUBS 0.029367f
C133 VN.n21 VSUBS 0.031612f
C134 VN.t3 VSUBS 2.11084f
C135 VN.n22 VSUBS 0.891973f
C136 VN.t2 VSUBS 2.52136f
C137 VN.n23 VSUBS 0.8329f
C138 VN.n24 VSUBS 0.385625f
C139 VN.n25 VSUBS 0.058622f
C140 VN.n26 VSUBS 0.058622f
C141 VN.n27 VSUBS 0.058036f
C142 VN.n28 VSUBS 0.031612f
C143 VN.n29 VSUBS 0.031612f
C144 VN.n30 VSUBS 0.031612f
C145 VN.n31 VSUBS 0.063126f
C146 VN.n32 VSUBS 0.058622f
C147 VN.n33 VSUBS 0.047625f
C148 VN.n34 VSUBS 0.051014f
C149 VN.n35 VSUBS 1.74493f
C150 VTAIL.t1 VSUBS 0.18909f
C151 VTAIL.t3 VSUBS 0.18909f
C152 VTAIL.n0 VSUBS 1.20682f
C153 VTAIL.n1 VSUBS 0.953142f
C154 VTAIL.n2 VSUBS 0.035005f
C155 VTAIL.n3 VSUBS 0.033327f
C156 VTAIL.n4 VSUBS 0.017908f
C157 VTAIL.n5 VSUBS 0.042329f
C158 VTAIL.n6 VSUBS 0.018962f
C159 VTAIL.n7 VSUBS 0.033327f
C160 VTAIL.n8 VSUBS 0.017908f
C161 VTAIL.n9 VSUBS 0.042329f
C162 VTAIL.n10 VSUBS 0.018962f
C163 VTAIL.n11 VSUBS 0.933205f
C164 VTAIL.n12 VSUBS 0.017908f
C165 VTAIL.t6 VSUBS 0.09089f
C166 VTAIL.n13 VSUBS 0.190014f
C167 VTAIL.n14 VSUBS 0.03184f
C168 VTAIL.n15 VSUBS 0.031746f
C169 VTAIL.n16 VSUBS 0.042329f
C170 VTAIL.n17 VSUBS 0.018962f
C171 VTAIL.n18 VSUBS 0.017908f
C172 VTAIL.n19 VSUBS 0.033327f
C173 VTAIL.n20 VSUBS 0.033327f
C174 VTAIL.n21 VSUBS 0.017908f
C175 VTAIL.n22 VSUBS 0.018962f
C176 VTAIL.n23 VSUBS 0.042329f
C177 VTAIL.n24 VSUBS 0.042329f
C178 VTAIL.n25 VSUBS 0.018962f
C179 VTAIL.n26 VSUBS 0.017908f
C180 VTAIL.n27 VSUBS 0.033327f
C181 VTAIL.n28 VSUBS 0.033327f
C182 VTAIL.n29 VSUBS 0.017908f
C183 VTAIL.n30 VSUBS 0.018962f
C184 VTAIL.n31 VSUBS 0.042329f
C185 VTAIL.n32 VSUBS 0.103507f
C186 VTAIL.n33 VSUBS 0.018962f
C187 VTAIL.n34 VSUBS 0.035168f
C188 VTAIL.n35 VSUBS 0.081586f
C189 VTAIL.n36 VSUBS 0.078408f
C190 VTAIL.n37 VSUBS 0.61055f
C191 VTAIL.t8 VSUBS 0.18909f
C192 VTAIL.t10 VSUBS 0.18909f
C193 VTAIL.n38 VSUBS 1.20682f
C194 VTAIL.n39 VSUBS 2.80741f
C195 VTAIL.t2 VSUBS 0.18909f
C196 VTAIL.t5 VSUBS 0.18909f
C197 VTAIL.n40 VSUBS 1.20683f
C198 VTAIL.n41 VSUBS 2.80741f
C199 VTAIL.n42 VSUBS 0.035005f
C200 VTAIL.n43 VSUBS 0.033327f
C201 VTAIL.n44 VSUBS 0.017908f
C202 VTAIL.n45 VSUBS 0.042329f
C203 VTAIL.n46 VSUBS 0.018962f
C204 VTAIL.n47 VSUBS 0.033327f
C205 VTAIL.n48 VSUBS 0.017908f
C206 VTAIL.n49 VSUBS 0.042329f
C207 VTAIL.n50 VSUBS 0.018962f
C208 VTAIL.n51 VSUBS 0.933206f
C209 VTAIL.n52 VSUBS 0.017908f
C210 VTAIL.t0 VSUBS 0.09089f
C211 VTAIL.n53 VSUBS 0.190014f
C212 VTAIL.n54 VSUBS 0.03184f
C213 VTAIL.n55 VSUBS 0.031746f
C214 VTAIL.n56 VSUBS 0.042329f
C215 VTAIL.n57 VSUBS 0.018962f
C216 VTAIL.n58 VSUBS 0.017908f
C217 VTAIL.n59 VSUBS 0.033327f
C218 VTAIL.n60 VSUBS 0.033327f
C219 VTAIL.n61 VSUBS 0.017908f
C220 VTAIL.n62 VSUBS 0.018962f
C221 VTAIL.n63 VSUBS 0.042329f
C222 VTAIL.n64 VSUBS 0.042329f
C223 VTAIL.n65 VSUBS 0.018962f
C224 VTAIL.n66 VSUBS 0.017908f
C225 VTAIL.n67 VSUBS 0.033327f
C226 VTAIL.n68 VSUBS 0.033327f
C227 VTAIL.n69 VSUBS 0.017908f
C228 VTAIL.n70 VSUBS 0.018962f
C229 VTAIL.n71 VSUBS 0.042329f
C230 VTAIL.n72 VSUBS 0.103507f
C231 VTAIL.n73 VSUBS 0.018962f
C232 VTAIL.n74 VSUBS 0.035168f
C233 VTAIL.n75 VSUBS 0.081586f
C234 VTAIL.n76 VSUBS 0.078408f
C235 VTAIL.n77 VSUBS 0.61055f
C236 VTAIL.t9 VSUBS 0.18909f
C237 VTAIL.t11 VSUBS 0.18909f
C238 VTAIL.n78 VSUBS 1.20683f
C239 VTAIL.n79 VSUBS 1.21141f
C240 VTAIL.n80 VSUBS 0.035005f
C241 VTAIL.n81 VSUBS 0.033327f
C242 VTAIL.n82 VSUBS 0.017908f
C243 VTAIL.n83 VSUBS 0.042329f
C244 VTAIL.n84 VSUBS 0.018962f
C245 VTAIL.n85 VSUBS 0.033327f
C246 VTAIL.n86 VSUBS 0.017908f
C247 VTAIL.n87 VSUBS 0.042329f
C248 VTAIL.n88 VSUBS 0.018962f
C249 VTAIL.n89 VSUBS 0.933206f
C250 VTAIL.n90 VSUBS 0.017908f
C251 VTAIL.t7 VSUBS 0.09089f
C252 VTAIL.n91 VSUBS 0.190014f
C253 VTAIL.n92 VSUBS 0.03184f
C254 VTAIL.n93 VSUBS 0.031746f
C255 VTAIL.n94 VSUBS 0.042329f
C256 VTAIL.n95 VSUBS 0.018962f
C257 VTAIL.n96 VSUBS 0.017908f
C258 VTAIL.n97 VSUBS 0.033327f
C259 VTAIL.n98 VSUBS 0.033327f
C260 VTAIL.n99 VSUBS 0.017908f
C261 VTAIL.n100 VSUBS 0.018962f
C262 VTAIL.n101 VSUBS 0.042329f
C263 VTAIL.n102 VSUBS 0.042329f
C264 VTAIL.n103 VSUBS 0.018962f
C265 VTAIL.n104 VSUBS 0.017908f
C266 VTAIL.n105 VSUBS 0.033327f
C267 VTAIL.n106 VSUBS 0.033327f
C268 VTAIL.n107 VSUBS 0.017908f
C269 VTAIL.n108 VSUBS 0.018962f
C270 VTAIL.n109 VSUBS 0.042329f
C271 VTAIL.n110 VSUBS 0.103507f
C272 VTAIL.n111 VSUBS 0.018962f
C273 VTAIL.n112 VSUBS 0.035168f
C274 VTAIL.n113 VSUBS 0.081586f
C275 VTAIL.n114 VSUBS 0.078408f
C276 VTAIL.n115 VSUBS 1.85383f
C277 VTAIL.n116 VSUBS 0.035005f
C278 VTAIL.n117 VSUBS 0.033327f
C279 VTAIL.n118 VSUBS 0.017908f
C280 VTAIL.n119 VSUBS 0.042329f
C281 VTAIL.n120 VSUBS 0.018962f
C282 VTAIL.n121 VSUBS 0.033327f
C283 VTAIL.n122 VSUBS 0.017908f
C284 VTAIL.n123 VSUBS 0.042329f
C285 VTAIL.n124 VSUBS 0.018962f
C286 VTAIL.n125 VSUBS 0.933205f
C287 VTAIL.n126 VSUBS 0.017908f
C288 VTAIL.t4 VSUBS 0.09089f
C289 VTAIL.n127 VSUBS 0.190014f
C290 VTAIL.n128 VSUBS 0.03184f
C291 VTAIL.n129 VSUBS 0.031746f
C292 VTAIL.n130 VSUBS 0.042329f
C293 VTAIL.n131 VSUBS 0.018962f
C294 VTAIL.n132 VSUBS 0.017908f
C295 VTAIL.n133 VSUBS 0.033327f
C296 VTAIL.n134 VSUBS 0.033327f
C297 VTAIL.n135 VSUBS 0.017908f
C298 VTAIL.n136 VSUBS 0.018962f
C299 VTAIL.n137 VSUBS 0.042329f
C300 VTAIL.n138 VSUBS 0.042329f
C301 VTAIL.n139 VSUBS 0.018962f
C302 VTAIL.n140 VSUBS 0.017908f
C303 VTAIL.n141 VSUBS 0.033327f
C304 VTAIL.n142 VSUBS 0.033327f
C305 VTAIL.n143 VSUBS 0.017908f
C306 VTAIL.n144 VSUBS 0.018962f
C307 VTAIL.n145 VSUBS 0.042329f
C308 VTAIL.n146 VSUBS 0.103507f
C309 VTAIL.n147 VSUBS 0.018962f
C310 VTAIL.n148 VSUBS 0.035168f
C311 VTAIL.n149 VSUBS 0.081586f
C312 VTAIL.n150 VSUBS 0.078408f
C313 VTAIL.n151 VSUBS 1.75941f
C314 VDD1.n0 VSUBS 0.027897f
C315 VDD1.n1 VSUBS 0.02656f
C316 VDD1.n2 VSUBS 0.014272f
C317 VDD1.n3 VSUBS 0.033734f
C318 VDD1.n4 VSUBS 0.015111f
C319 VDD1.n5 VSUBS 0.02656f
C320 VDD1.n6 VSUBS 0.014272f
C321 VDD1.n7 VSUBS 0.033734f
C322 VDD1.n8 VSUBS 0.015111f
C323 VDD1.n9 VSUBS 0.743717f
C324 VDD1.n10 VSUBS 0.014272f
C325 VDD1.t5 VSUBS 0.072435f
C326 VDD1.n11 VSUBS 0.151432f
C327 VDD1.n12 VSUBS 0.025375f
C328 VDD1.n13 VSUBS 0.0253f
C329 VDD1.n14 VSUBS 0.033734f
C330 VDD1.n15 VSUBS 0.015111f
C331 VDD1.n16 VSUBS 0.014272f
C332 VDD1.n17 VSUBS 0.02656f
C333 VDD1.n18 VSUBS 0.02656f
C334 VDD1.n19 VSUBS 0.014272f
C335 VDD1.n20 VSUBS 0.015111f
C336 VDD1.n21 VSUBS 0.033734f
C337 VDD1.n22 VSUBS 0.033734f
C338 VDD1.n23 VSUBS 0.015111f
C339 VDD1.n24 VSUBS 0.014272f
C340 VDD1.n25 VSUBS 0.02656f
C341 VDD1.n26 VSUBS 0.02656f
C342 VDD1.n27 VSUBS 0.014272f
C343 VDD1.n28 VSUBS 0.015111f
C344 VDD1.n29 VSUBS 0.033734f
C345 VDD1.n30 VSUBS 0.08249f
C346 VDD1.n31 VSUBS 0.015111f
C347 VDD1.n32 VSUBS 0.028027f
C348 VDD1.n33 VSUBS 0.06502f
C349 VDD1.n34 VSUBS 0.09352f
C350 VDD1.n35 VSUBS 0.027897f
C351 VDD1.n36 VSUBS 0.02656f
C352 VDD1.n37 VSUBS 0.014272f
C353 VDD1.n38 VSUBS 0.033734f
C354 VDD1.n39 VSUBS 0.015111f
C355 VDD1.n40 VSUBS 0.02656f
C356 VDD1.n41 VSUBS 0.014272f
C357 VDD1.n42 VSUBS 0.033734f
C358 VDD1.n43 VSUBS 0.015111f
C359 VDD1.n44 VSUBS 0.743717f
C360 VDD1.n45 VSUBS 0.014272f
C361 VDD1.t4 VSUBS 0.072435f
C362 VDD1.n46 VSUBS 0.151432f
C363 VDD1.n47 VSUBS 0.025375f
C364 VDD1.n48 VSUBS 0.0253f
C365 VDD1.n49 VSUBS 0.033734f
C366 VDD1.n50 VSUBS 0.015111f
C367 VDD1.n51 VSUBS 0.014272f
C368 VDD1.n52 VSUBS 0.02656f
C369 VDD1.n53 VSUBS 0.02656f
C370 VDD1.n54 VSUBS 0.014272f
C371 VDD1.n55 VSUBS 0.015111f
C372 VDD1.n56 VSUBS 0.033734f
C373 VDD1.n57 VSUBS 0.033734f
C374 VDD1.n58 VSUBS 0.015111f
C375 VDD1.n59 VSUBS 0.014272f
C376 VDD1.n60 VSUBS 0.02656f
C377 VDD1.n61 VSUBS 0.02656f
C378 VDD1.n62 VSUBS 0.014272f
C379 VDD1.n63 VSUBS 0.015111f
C380 VDD1.n64 VSUBS 0.033734f
C381 VDD1.n65 VSUBS 0.08249f
C382 VDD1.n66 VSUBS 0.015111f
C383 VDD1.n67 VSUBS 0.028027f
C384 VDD1.n68 VSUBS 0.06502f
C385 VDD1.n69 VSUBS 0.092545f
C386 VDD1.t0 VSUBS 0.150695f
C387 VDD1.t2 VSUBS 0.150695f
C388 VDD1.n70 VSUBS 1.07148f
C389 VDD1.n71 VSUBS 3.30667f
C390 VDD1.t1 VSUBS 0.150695f
C391 VDD1.t3 VSUBS 0.150695f
C392 VDD1.n72 VSUBS 1.06453f
C393 VDD1.n73 VSUBS 3.05281f
C394 VP.t5 VSUBS 2.38562f
C395 VP.n0 VSUBS 1.01438f
C396 VP.n1 VSUBS 0.035727f
C397 VP.n2 VSUBS 0.033189f
C398 VP.n3 VSUBS 0.035727f
C399 VP.t1 VSUBS 2.38562f
C400 VP.n4 VSUBS 0.900175f
C401 VP.n5 VSUBS 0.035727f
C402 VP.n6 VSUBS 0.033189f
C403 VP.n7 VSUBS 0.035727f
C404 VP.t3 VSUBS 2.38562f
C405 VP.n8 VSUBS 1.01438f
C406 VP.t4 VSUBS 2.38562f
C407 VP.n9 VSUBS 1.01438f
C408 VP.n10 VSUBS 0.035727f
C409 VP.n11 VSUBS 0.033189f
C410 VP.n12 VSUBS 0.035727f
C411 VP.t0 VSUBS 2.38562f
C412 VP.n13 VSUBS 1.00809f
C413 VP.t2 VSUBS 2.84957f
C414 VP.n14 VSUBS 0.941325f
C415 VP.n15 VSUBS 0.435824f
C416 VP.n16 VSUBS 0.066253f
C417 VP.n17 VSUBS 0.066253f
C418 VP.n18 VSUBS 0.065591f
C419 VP.n19 VSUBS 0.035727f
C420 VP.n20 VSUBS 0.035727f
C421 VP.n21 VSUBS 0.035727f
C422 VP.n22 VSUBS 0.071344f
C423 VP.n23 VSUBS 0.066253f
C424 VP.n24 VSUBS 0.053824f
C425 VP.n25 VSUBS 0.057654f
C426 VP.n26 VSUBS 1.95733f
C427 VP.n27 VSUBS 1.98381f
C428 VP.n28 VSUBS 0.057654f
C429 VP.n29 VSUBS 0.053824f
C430 VP.n30 VSUBS 0.066253f
C431 VP.n31 VSUBS 0.071344f
C432 VP.n32 VSUBS 0.035727f
C433 VP.n33 VSUBS 0.035727f
C434 VP.n34 VSUBS 0.035727f
C435 VP.n35 VSUBS 0.065591f
C436 VP.n36 VSUBS 0.066253f
C437 VP.n37 VSUBS 0.066253f
C438 VP.n38 VSUBS 0.035727f
C439 VP.n39 VSUBS 0.035727f
C440 VP.n40 VSUBS 0.035727f
C441 VP.n41 VSUBS 0.066253f
C442 VP.n42 VSUBS 0.066253f
C443 VP.n43 VSUBS 0.065591f
C444 VP.n44 VSUBS 0.035727f
C445 VP.n45 VSUBS 0.035727f
C446 VP.n46 VSUBS 0.035727f
C447 VP.n47 VSUBS 0.071344f
C448 VP.n48 VSUBS 0.066253f
C449 VP.n49 VSUBS 0.053824f
C450 VP.n50 VSUBS 0.057654f
C451 VP.n51 VSUBS 0.08825f
C452 B.n0 VSUBS 0.00589f
C453 B.n1 VSUBS 0.00589f
C454 B.n2 VSUBS 0.009315f
C455 B.n3 VSUBS 0.009315f
C456 B.n4 VSUBS 0.009315f
C457 B.n5 VSUBS 0.009315f
C458 B.n6 VSUBS 0.009315f
C459 B.n7 VSUBS 0.009315f
C460 B.n8 VSUBS 0.009315f
C461 B.n9 VSUBS 0.009315f
C462 B.n10 VSUBS 0.009315f
C463 B.n11 VSUBS 0.009315f
C464 B.n12 VSUBS 0.009315f
C465 B.n13 VSUBS 0.009315f
C466 B.n14 VSUBS 0.009315f
C467 B.n15 VSUBS 0.009315f
C468 B.n16 VSUBS 0.009315f
C469 B.n17 VSUBS 0.009315f
C470 B.n18 VSUBS 0.009315f
C471 B.n19 VSUBS 0.009315f
C472 B.n20 VSUBS 0.009315f
C473 B.n21 VSUBS 0.009315f
C474 B.n22 VSUBS 0.009315f
C475 B.n23 VSUBS 0.009315f
C476 B.n24 VSUBS 0.009315f
C477 B.n25 VSUBS 0.009315f
C478 B.n26 VSUBS 0.009315f
C479 B.n27 VSUBS 0.009315f
C480 B.n28 VSUBS 0.022222f
C481 B.n29 VSUBS 0.009315f
C482 B.n30 VSUBS 0.009315f
C483 B.n31 VSUBS 0.009315f
C484 B.n32 VSUBS 0.009315f
C485 B.n33 VSUBS 0.009315f
C486 B.n34 VSUBS 0.009315f
C487 B.n35 VSUBS 0.009315f
C488 B.n36 VSUBS 0.009315f
C489 B.n37 VSUBS 0.009315f
C490 B.n38 VSUBS 0.009315f
C491 B.n39 VSUBS 0.009315f
C492 B.n40 VSUBS 0.009315f
C493 B.n41 VSUBS 0.009315f
C494 B.t5 VSUBS 0.147174f
C495 B.t4 VSUBS 0.193711f
C496 B.t3 VSUBS 1.58165f
C497 B.n42 VSUBS 0.31918f
C498 B.n43 VSUBS 0.241712f
C499 B.n44 VSUBS 0.021582f
C500 B.n45 VSUBS 0.009315f
C501 B.n46 VSUBS 0.009315f
C502 B.n47 VSUBS 0.009315f
C503 B.n48 VSUBS 0.009315f
C504 B.n49 VSUBS 0.009315f
C505 B.t11 VSUBS 0.147177f
C506 B.t10 VSUBS 0.193713f
C507 B.t9 VSUBS 1.58165f
C508 B.n50 VSUBS 0.319177f
C509 B.n51 VSUBS 0.241709f
C510 B.n52 VSUBS 0.009315f
C511 B.n53 VSUBS 0.009315f
C512 B.n54 VSUBS 0.009315f
C513 B.n55 VSUBS 0.009315f
C514 B.n56 VSUBS 0.009315f
C515 B.n57 VSUBS 0.009315f
C516 B.n58 VSUBS 0.009315f
C517 B.n59 VSUBS 0.009315f
C518 B.n60 VSUBS 0.009315f
C519 B.n61 VSUBS 0.009315f
C520 B.n62 VSUBS 0.009315f
C521 B.n63 VSUBS 0.009315f
C522 B.n64 VSUBS 0.009315f
C523 B.n65 VSUBS 0.022222f
C524 B.n66 VSUBS 0.009315f
C525 B.n67 VSUBS 0.009315f
C526 B.n68 VSUBS 0.009315f
C527 B.n69 VSUBS 0.009315f
C528 B.n70 VSUBS 0.009315f
C529 B.n71 VSUBS 0.009315f
C530 B.n72 VSUBS 0.009315f
C531 B.n73 VSUBS 0.009315f
C532 B.n74 VSUBS 0.009315f
C533 B.n75 VSUBS 0.009315f
C534 B.n76 VSUBS 0.009315f
C535 B.n77 VSUBS 0.009315f
C536 B.n78 VSUBS 0.009315f
C537 B.n79 VSUBS 0.009315f
C538 B.n80 VSUBS 0.009315f
C539 B.n81 VSUBS 0.009315f
C540 B.n82 VSUBS 0.009315f
C541 B.n83 VSUBS 0.009315f
C542 B.n84 VSUBS 0.009315f
C543 B.n85 VSUBS 0.009315f
C544 B.n86 VSUBS 0.009315f
C545 B.n87 VSUBS 0.009315f
C546 B.n88 VSUBS 0.009315f
C547 B.n89 VSUBS 0.009315f
C548 B.n90 VSUBS 0.009315f
C549 B.n91 VSUBS 0.009315f
C550 B.n92 VSUBS 0.009315f
C551 B.n93 VSUBS 0.009315f
C552 B.n94 VSUBS 0.009315f
C553 B.n95 VSUBS 0.009315f
C554 B.n96 VSUBS 0.009315f
C555 B.n97 VSUBS 0.009315f
C556 B.n98 VSUBS 0.009315f
C557 B.n99 VSUBS 0.009315f
C558 B.n100 VSUBS 0.009315f
C559 B.n101 VSUBS 0.009315f
C560 B.n102 VSUBS 0.009315f
C561 B.n103 VSUBS 0.009315f
C562 B.n104 VSUBS 0.009315f
C563 B.n105 VSUBS 0.009315f
C564 B.n106 VSUBS 0.009315f
C565 B.n107 VSUBS 0.009315f
C566 B.n108 VSUBS 0.009315f
C567 B.n109 VSUBS 0.009315f
C568 B.n110 VSUBS 0.009315f
C569 B.n111 VSUBS 0.009315f
C570 B.n112 VSUBS 0.009315f
C571 B.n113 VSUBS 0.009315f
C572 B.n114 VSUBS 0.009315f
C573 B.n115 VSUBS 0.009315f
C574 B.n116 VSUBS 0.009315f
C575 B.n117 VSUBS 0.009315f
C576 B.n118 VSUBS 0.022222f
C577 B.n119 VSUBS 0.009315f
C578 B.n120 VSUBS 0.009315f
C579 B.n121 VSUBS 0.009315f
C580 B.n122 VSUBS 0.009315f
C581 B.n123 VSUBS 0.009315f
C582 B.n124 VSUBS 0.009315f
C583 B.n125 VSUBS 0.009315f
C584 B.n126 VSUBS 0.009315f
C585 B.n127 VSUBS 0.009315f
C586 B.n128 VSUBS 0.009315f
C587 B.n129 VSUBS 0.009315f
C588 B.n130 VSUBS 0.009315f
C589 B.n131 VSUBS 0.009315f
C590 B.t7 VSUBS 0.147177f
C591 B.t8 VSUBS 0.193713f
C592 B.t6 VSUBS 1.58165f
C593 B.n132 VSUBS 0.319177f
C594 B.n133 VSUBS 0.241709f
C595 B.n134 VSUBS 0.021582f
C596 B.n135 VSUBS 0.009315f
C597 B.n136 VSUBS 0.009315f
C598 B.n137 VSUBS 0.009315f
C599 B.n138 VSUBS 0.009315f
C600 B.n139 VSUBS 0.009315f
C601 B.t1 VSUBS 0.147174f
C602 B.t2 VSUBS 0.193711f
C603 B.t0 VSUBS 1.58165f
C604 B.n140 VSUBS 0.31918f
C605 B.n141 VSUBS 0.241712f
C606 B.n142 VSUBS 0.009315f
C607 B.n143 VSUBS 0.009315f
C608 B.n144 VSUBS 0.009315f
C609 B.n145 VSUBS 0.009315f
C610 B.n146 VSUBS 0.009315f
C611 B.n147 VSUBS 0.009315f
C612 B.n148 VSUBS 0.009315f
C613 B.n149 VSUBS 0.009315f
C614 B.n150 VSUBS 0.009315f
C615 B.n151 VSUBS 0.009315f
C616 B.n152 VSUBS 0.009315f
C617 B.n153 VSUBS 0.009315f
C618 B.n154 VSUBS 0.009315f
C619 B.n155 VSUBS 0.022222f
C620 B.n156 VSUBS 0.009315f
C621 B.n157 VSUBS 0.009315f
C622 B.n158 VSUBS 0.009315f
C623 B.n159 VSUBS 0.009315f
C624 B.n160 VSUBS 0.009315f
C625 B.n161 VSUBS 0.009315f
C626 B.n162 VSUBS 0.009315f
C627 B.n163 VSUBS 0.009315f
C628 B.n164 VSUBS 0.009315f
C629 B.n165 VSUBS 0.009315f
C630 B.n166 VSUBS 0.009315f
C631 B.n167 VSUBS 0.009315f
C632 B.n168 VSUBS 0.009315f
C633 B.n169 VSUBS 0.009315f
C634 B.n170 VSUBS 0.009315f
C635 B.n171 VSUBS 0.009315f
C636 B.n172 VSUBS 0.009315f
C637 B.n173 VSUBS 0.009315f
C638 B.n174 VSUBS 0.009315f
C639 B.n175 VSUBS 0.009315f
C640 B.n176 VSUBS 0.009315f
C641 B.n177 VSUBS 0.009315f
C642 B.n178 VSUBS 0.009315f
C643 B.n179 VSUBS 0.009315f
C644 B.n180 VSUBS 0.009315f
C645 B.n181 VSUBS 0.009315f
C646 B.n182 VSUBS 0.009315f
C647 B.n183 VSUBS 0.009315f
C648 B.n184 VSUBS 0.009315f
C649 B.n185 VSUBS 0.009315f
C650 B.n186 VSUBS 0.009315f
C651 B.n187 VSUBS 0.009315f
C652 B.n188 VSUBS 0.009315f
C653 B.n189 VSUBS 0.009315f
C654 B.n190 VSUBS 0.009315f
C655 B.n191 VSUBS 0.009315f
C656 B.n192 VSUBS 0.009315f
C657 B.n193 VSUBS 0.009315f
C658 B.n194 VSUBS 0.009315f
C659 B.n195 VSUBS 0.009315f
C660 B.n196 VSUBS 0.009315f
C661 B.n197 VSUBS 0.009315f
C662 B.n198 VSUBS 0.009315f
C663 B.n199 VSUBS 0.009315f
C664 B.n200 VSUBS 0.009315f
C665 B.n201 VSUBS 0.009315f
C666 B.n202 VSUBS 0.009315f
C667 B.n203 VSUBS 0.009315f
C668 B.n204 VSUBS 0.009315f
C669 B.n205 VSUBS 0.009315f
C670 B.n206 VSUBS 0.009315f
C671 B.n207 VSUBS 0.009315f
C672 B.n208 VSUBS 0.009315f
C673 B.n209 VSUBS 0.009315f
C674 B.n210 VSUBS 0.009315f
C675 B.n211 VSUBS 0.009315f
C676 B.n212 VSUBS 0.009315f
C677 B.n213 VSUBS 0.009315f
C678 B.n214 VSUBS 0.009315f
C679 B.n215 VSUBS 0.009315f
C680 B.n216 VSUBS 0.009315f
C681 B.n217 VSUBS 0.009315f
C682 B.n218 VSUBS 0.009315f
C683 B.n219 VSUBS 0.009315f
C684 B.n220 VSUBS 0.009315f
C685 B.n221 VSUBS 0.009315f
C686 B.n222 VSUBS 0.009315f
C687 B.n223 VSUBS 0.009315f
C688 B.n224 VSUBS 0.009315f
C689 B.n225 VSUBS 0.009315f
C690 B.n226 VSUBS 0.009315f
C691 B.n227 VSUBS 0.009315f
C692 B.n228 VSUBS 0.009315f
C693 B.n229 VSUBS 0.009315f
C694 B.n230 VSUBS 0.009315f
C695 B.n231 VSUBS 0.009315f
C696 B.n232 VSUBS 0.009315f
C697 B.n233 VSUBS 0.009315f
C698 B.n234 VSUBS 0.009315f
C699 B.n235 VSUBS 0.009315f
C700 B.n236 VSUBS 0.009315f
C701 B.n237 VSUBS 0.009315f
C702 B.n238 VSUBS 0.009315f
C703 B.n239 VSUBS 0.009315f
C704 B.n240 VSUBS 0.009315f
C705 B.n241 VSUBS 0.009315f
C706 B.n242 VSUBS 0.009315f
C707 B.n243 VSUBS 0.009315f
C708 B.n244 VSUBS 0.009315f
C709 B.n245 VSUBS 0.009315f
C710 B.n246 VSUBS 0.009315f
C711 B.n247 VSUBS 0.009315f
C712 B.n248 VSUBS 0.009315f
C713 B.n249 VSUBS 0.009315f
C714 B.n250 VSUBS 0.009315f
C715 B.n251 VSUBS 0.009315f
C716 B.n252 VSUBS 0.009315f
C717 B.n253 VSUBS 0.009315f
C718 B.n254 VSUBS 0.009315f
C719 B.n255 VSUBS 0.009315f
C720 B.n256 VSUBS 0.009315f
C721 B.n257 VSUBS 0.009315f
C722 B.n258 VSUBS 0.022222f
C723 B.n259 VSUBS 0.022709f
C724 B.n260 VSUBS 0.022709f
C725 B.n261 VSUBS 0.009315f
C726 B.n262 VSUBS 0.009315f
C727 B.n263 VSUBS 0.009315f
C728 B.n264 VSUBS 0.009315f
C729 B.n265 VSUBS 0.009315f
C730 B.n266 VSUBS 0.009315f
C731 B.n267 VSUBS 0.009315f
C732 B.n268 VSUBS 0.009315f
C733 B.n269 VSUBS 0.009315f
C734 B.n270 VSUBS 0.009315f
C735 B.n271 VSUBS 0.009315f
C736 B.n272 VSUBS 0.009315f
C737 B.n273 VSUBS 0.009315f
C738 B.n274 VSUBS 0.009315f
C739 B.n275 VSUBS 0.009315f
C740 B.n276 VSUBS 0.009315f
C741 B.n277 VSUBS 0.009315f
C742 B.n278 VSUBS 0.009315f
C743 B.n279 VSUBS 0.009315f
C744 B.n280 VSUBS 0.009315f
C745 B.n281 VSUBS 0.009315f
C746 B.n282 VSUBS 0.009315f
C747 B.n283 VSUBS 0.009315f
C748 B.n284 VSUBS 0.009315f
C749 B.n285 VSUBS 0.009315f
C750 B.n286 VSUBS 0.009315f
C751 B.n287 VSUBS 0.009315f
C752 B.n288 VSUBS 0.009315f
C753 B.n289 VSUBS 0.009315f
C754 B.n290 VSUBS 0.009315f
C755 B.n291 VSUBS 0.009315f
C756 B.n292 VSUBS 0.009315f
C757 B.n293 VSUBS 0.009315f
C758 B.n294 VSUBS 0.009315f
C759 B.n295 VSUBS 0.009315f
C760 B.n296 VSUBS 0.009315f
C761 B.n297 VSUBS 0.009315f
C762 B.n298 VSUBS 0.009315f
C763 B.n299 VSUBS 0.008767f
C764 B.n300 VSUBS 0.021582f
C765 B.n301 VSUBS 0.005205f
C766 B.n302 VSUBS 0.009315f
C767 B.n303 VSUBS 0.009315f
C768 B.n304 VSUBS 0.009315f
C769 B.n305 VSUBS 0.009315f
C770 B.n306 VSUBS 0.009315f
C771 B.n307 VSUBS 0.009315f
C772 B.n308 VSUBS 0.009315f
C773 B.n309 VSUBS 0.009315f
C774 B.n310 VSUBS 0.009315f
C775 B.n311 VSUBS 0.009315f
C776 B.n312 VSUBS 0.009315f
C777 B.n313 VSUBS 0.009315f
C778 B.n314 VSUBS 0.005205f
C779 B.n315 VSUBS 0.009315f
C780 B.n316 VSUBS 0.009315f
C781 B.n317 VSUBS 0.008767f
C782 B.n318 VSUBS 0.009315f
C783 B.n319 VSUBS 0.009315f
C784 B.n320 VSUBS 0.009315f
C785 B.n321 VSUBS 0.009315f
C786 B.n322 VSUBS 0.009315f
C787 B.n323 VSUBS 0.009315f
C788 B.n324 VSUBS 0.009315f
C789 B.n325 VSUBS 0.009315f
C790 B.n326 VSUBS 0.009315f
C791 B.n327 VSUBS 0.009315f
C792 B.n328 VSUBS 0.009315f
C793 B.n329 VSUBS 0.009315f
C794 B.n330 VSUBS 0.009315f
C795 B.n331 VSUBS 0.009315f
C796 B.n332 VSUBS 0.009315f
C797 B.n333 VSUBS 0.009315f
C798 B.n334 VSUBS 0.009315f
C799 B.n335 VSUBS 0.009315f
C800 B.n336 VSUBS 0.009315f
C801 B.n337 VSUBS 0.009315f
C802 B.n338 VSUBS 0.009315f
C803 B.n339 VSUBS 0.009315f
C804 B.n340 VSUBS 0.009315f
C805 B.n341 VSUBS 0.009315f
C806 B.n342 VSUBS 0.009315f
C807 B.n343 VSUBS 0.009315f
C808 B.n344 VSUBS 0.009315f
C809 B.n345 VSUBS 0.009315f
C810 B.n346 VSUBS 0.009315f
C811 B.n347 VSUBS 0.009315f
C812 B.n348 VSUBS 0.009315f
C813 B.n349 VSUBS 0.009315f
C814 B.n350 VSUBS 0.009315f
C815 B.n351 VSUBS 0.009315f
C816 B.n352 VSUBS 0.009315f
C817 B.n353 VSUBS 0.009315f
C818 B.n354 VSUBS 0.009315f
C819 B.n355 VSUBS 0.022709f
C820 B.n356 VSUBS 0.022709f
C821 B.n357 VSUBS 0.022222f
C822 B.n358 VSUBS 0.009315f
C823 B.n359 VSUBS 0.009315f
C824 B.n360 VSUBS 0.009315f
C825 B.n361 VSUBS 0.009315f
C826 B.n362 VSUBS 0.009315f
C827 B.n363 VSUBS 0.009315f
C828 B.n364 VSUBS 0.009315f
C829 B.n365 VSUBS 0.009315f
C830 B.n366 VSUBS 0.009315f
C831 B.n367 VSUBS 0.009315f
C832 B.n368 VSUBS 0.009315f
C833 B.n369 VSUBS 0.009315f
C834 B.n370 VSUBS 0.009315f
C835 B.n371 VSUBS 0.009315f
C836 B.n372 VSUBS 0.009315f
C837 B.n373 VSUBS 0.009315f
C838 B.n374 VSUBS 0.009315f
C839 B.n375 VSUBS 0.009315f
C840 B.n376 VSUBS 0.009315f
C841 B.n377 VSUBS 0.009315f
C842 B.n378 VSUBS 0.009315f
C843 B.n379 VSUBS 0.009315f
C844 B.n380 VSUBS 0.009315f
C845 B.n381 VSUBS 0.009315f
C846 B.n382 VSUBS 0.009315f
C847 B.n383 VSUBS 0.009315f
C848 B.n384 VSUBS 0.009315f
C849 B.n385 VSUBS 0.009315f
C850 B.n386 VSUBS 0.009315f
C851 B.n387 VSUBS 0.009315f
C852 B.n388 VSUBS 0.009315f
C853 B.n389 VSUBS 0.009315f
C854 B.n390 VSUBS 0.009315f
C855 B.n391 VSUBS 0.009315f
C856 B.n392 VSUBS 0.009315f
C857 B.n393 VSUBS 0.009315f
C858 B.n394 VSUBS 0.009315f
C859 B.n395 VSUBS 0.009315f
C860 B.n396 VSUBS 0.009315f
C861 B.n397 VSUBS 0.009315f
C862 B.n398 VSUBS 0.009315f
C863 B.n399 VSUBS 0.009315f
C864 B.n400 VSUBS 0.009315f
C865 B.n401 VSUBS 0.009315f
C866 B.n402 VSUBS 0.009315f
C867 B.n403 VSUBS 0.009315f
C868 B.n404 VSUBS 0.009315f
C869 B.n405 VSUBS 0.009315f
C870 B.n406 VSUBS 0.009315f
C871 B.n407 VSUBS 0.009315f
C872 B.n408 VSUBS 0.009315f
C873 B.n409 VSUBS 0.009315f
C874 B.n410 VSUBS 0.009315f
C875 B.n411 VSUBS 0.009315f
C876 B.n412 VSUBS 0.009315f
C877 B.n413 VSUBS 0.009315f
C878 B.n414 VSUBS 0.009315f
C879 B.n415 VSUBS 0.009315f
C880 B.n416 VSUBS 0.009315f
C881 B.n417 VSUBS 0.009315f
C882 B.n418 VSUBS 0.009315f
C883 B.n419 VSUBS 0.009315f
C884 B.n420 VSUBS 0.009315f
C885 B.n421 VSUBS 0.009315f
C886 B.n422 VSUBS 0.009315f
C887 B.n423 VSUBS 0.009315f
C888 B.n424 VSUBS 0.009315f
C889 B.n425 VSUBS 0.009315f
C890 B.n426 VSUBS 0.009315f
C891 B.n427 VSUBS 0.009315f
C892 B.n428 VSUBS 0.009315f
C893 B.n429 VSUBS 0.009315f
C894 B.n430 VSUBS 0.009315f
C895 B.n431 VSUBS 0.009315f
C896 B.n432 VSUBS 0.009315f
C897 B.n433 VSUBS 0.009315f
C898 B.n434 VSUBS 0.009315f
C899 B.n435 VSUBS 0.009315f
C900 B.n436 VSUBS 0.009315f
C901 B.n437 VSUBS 0.009315f
C902 B.n438 VSUBS 0.009315f
C903 B.n439 VSUBS 0.009315f
C904 B.n440 VSUBS 0.009315f
C905 B.n441 VSUBS 0.009315f
C906 B.n442 VSUBS 0.009315f
C907 B.n443 VSUBS 0.009315f
C908 B.n444 VSUBS 0.009315f
C909 B.n445 VSUBS 0.009315f
C910 B.n446 VSUBS 0.009315f
C911 B.n447 VSUBS 0.009315f
C912 B.n448 VSUBS 0.009315f
C913 B.n449 VSUBS 0.009315f
C914 B.n450 VSUBS 0.009315f
C915 B.n451 VSUBS 0.009315f
C916 B.n452 VSUBS 0.009315f
C917 B.n453 VSUBS 0.009315f
C918 B.n454 VSUBS 0.009315f
C919 B.n455 VSUBS 0.009315f
C920 B.n456 VSUBS 0.009315f
C921 B.n457 VSUBS 0.009315f
C922 B.n458 VSUBS 0.009315f
C923 B.n459 VSUBS 0.009315f
C924 B.n460 VSUBS 0.009315f
C925 B.n461 VSUBS 0.009315f
C926 B.n462 VSUBS 0.009315f
C927 B.n463 VSUBS 0.009315f
C928 B.n464 VSUBS 0.009315f
C929 B.n465 VSUBS 0.009315f
C930 B.n466 VSUBS 0.009315f
C931 B.n467 VSUBS 0.009315f
C932 B.n468 VSUBS 0.009315f
C933 B.n469 VSUBS 0.009315f
C934 B.n470 VSUBS 0.009315f
C935 B.n471 VSUBS 0.009315f
C936 B.n472 VSUBS 0.009315f
C937 B.n473 VSUBS 0.009315f
C938 B.n474 VSUBS 0.009315f
C939 B.n475 VSUBS 0.009315f
C940 B.n476 VSUBS 0.009315f
C941 B.n477 VSUBS 0.009315f
C942 B.n478 VSUBS 0.009315f
C943 B.n479 VSUBS 0.009315f
C944 B.n480 VSUBS 0.009315f
C945 B.n481 VSUBS 0.009315f
C946 B.n482 VSUBS 0.009315f
C947 B.n483 VSUBS 0.009315f
C948 B.n484 VSUBS 0.009315f
C949 B.n485 VSUBS 0.009315f
C950 B.n486 VSUBS 0.009315f
C951 B.n487 VSUBS 0.009315f
C952 B.n488 VSUBS 0.009315f
C953 B.n489 VSUBS 0.009315f
C954 B.n490 VSUBS 0.009315f
C955 B.n491 VSUBS 0.009315f
C956 B.n492 VSUBS 0.009315f
C957 B.n493 VSUBS 0.009315f
C958 B.n494 VSUBS 0.009315f
C959 B.n495 VSUBS 0.009315f
C960 B.n496 VSUBS 0.009315f
C961 B.n497 VSUBS 0.009315f
C962 B.n498 VSUBS 0.009315f
C963 B.n499 VSUBS 0.009315f
C964 B.n500 VSUBS 0.009315f
C965 B.n501 VSUBS 0.009315f
C966 B.n502 VSUBS 0.009315f
C967 B.n503 VSUBS 0.009315f
C968 B.n504 VSUBS 0.009315f
C969 B.n505 VSUBS 0.009315f
C970 B.n506 VSUBS 0.009315f
C971 B.n507 VSUBS 0.009315f
C972 B.n508 VSUBS 0.009315f
C973 B.n509 VSUBS 0.009315f
C974 B.n510 VSUBS 0.009315f
C975 B.n511 VSUBS 0.009315f
C976 B.n512 VSUBS 0.009315f
C977 B.n513 VSUBS 0.009315f
C978 B.n514 VSUBS 0.009315f
C979 B.n515 VSUBS 0.009315f
C980 B.n516 VSUBS 0.023274f
C981 B.n517 VSUBS 0.021658f
C982 B.n518 VSUBS 0.022709f
C983 B.n519 VSUBS 0.009315f
C984 B.n520 VSUBS 0.009315f
C985 B.n521 VSUBS 0.009315f
C986 B.n522 VSUBS 0.009315f
C987 B.n523 VSUBS 0.009315f
C988 B.n524 VSUBS 0.009315f
C989 B.n525 VSUBS 0.009315f
C990 B.n526 VSUBS 0.009315f
C991 B.n527 VSUBS 0.009315f
C992 B.n528 VSUBS 0.009315f
C993 B.n529 VSUBS 0.009315f
C994 B.n530 VSUBS 0.009315f
C995 B.n531 VSUBS 0.009315f
C996 B.n532 VSUBS 0.009315f
C997 B.n533 VSUBS 0.009315f
C998 B.n534 VSUBS 0.009315f
C999 B.n535 VSUBS 0.009315f
C1000 B.n536 VSUBS 0.009315f
C1001 B.n537 VSUBS 0.009315f
C1002 B.n538 VSUBS 0.009315f
C1003 B.n539 VSUBS 0.009315f
C1004 B.n540 VSUBS 0.009315f
C1005 B.n541 VSUBS 0.009315f
C1006 B.n542 VSUBS 0.009315f
C1007 B.n543 VSUBS 0.009315f
C1008 B.n544 VSUBS 0.009315f
C1009 B.n545 VSUBS 0.009315f
C1010 B.n546 VSUBS 0.009315f
C1011 B.n547 VSUBS 0.009315f
C1012 B.n548 VSUBS 0.009315f
C1013 B.n549 VSUBS 0.009315f
C1014 B.n550 VSUBS 0.009315f
C1015 B.n551 VSUBS 0.009315f
C1016 B.n552 VSUBS 0.009315f
C1017 B.n553 VSUBS 0.009315f
C1018 B.n554 VSUBS 0.009315f
C1019 B.n555 VSUBS 0.009315f
C1020 B.n556 VSUBS 0.009315f
C1021 B.n557 VSUBS 0.008767f
C1022 B.n558 VSUBS 0.021582f
C1023 B.n559 VSUBS 0.005205f
C1024 B.n560 VSUBS 0.009315f
C1025 B.n561 VSUBS 0.009315f
C1026 B.n562 VSUBS 0.009315f
C1027 B.n563 VSUBS 0.009315f
C1028 B.n564 VSUBS 0.009315f
C1029 B.n565 VSUBS 0.009315f
C1030 B.n566 VSUBS 0.009315f
C1031 B.n567 VSUBS 0.009315f
C1032 B.n568 VSUBS 0.009315f
C1033 B.n569 VSUBS 0.009315f
C1034 B.n570 VSUBS 0.009315f
C1035 B.n571 VSUBS 0.009315f
C1036 B.n572 VSUBS 0.005205f
C1037 B.n573 VSUBS 0.009315f
C1038 B.n574 VSUBS 0.009315f
C1039 B.n575 VSUBS 0.008767f
C1040 B.n576 VSUBS 0.009315f
C1041 B.n577 VSUBS 0.009315f
C1042 B.n578 VSUBS 0.009315f
C1043 B.n579 VSUBS 0.009315f
C1044 B.n580 VSUBS 0.009315f
C1045 B.n581 VSUBS 0.009315f
C1046 B.n582 VSUBS 0.009315f
C1047 B.n583 VSUBS 0.009315f
C1048 B.n584 VSUBS 0.009315f
C1049 B.n585 VSUBS 0.009315f
C1050 B.n586 VSUBS 0.009315f
C1051 B.n587 VSUBS 0.009315f
C1052 B.n588 VSUBS 0.009315f
C1053 B.n589 VSUBS 0.009315f
C1054 B.n590 VSUBS 0.009315f
C1055 B.n591 VSUBS 0.009315f
C1056 B.n592 VSUBS 0.009315f
C1057 B.n593 VSUBS 0.009315f
C1058 B.n594 VSUBS 0.009315f
C1059 B.n595 VSUBS 0.009315f
C1060 B.n596 VSUBS 0.009315f
C1061 B.n597 VSUBS 0.009315f
C1062 B.n598 VSUBS 0.009315f
C1063 B.n599 VSUBS 0.009315f
C1064 B.n600 VSUBS 0.009315f
C1065 B.n601 VSUBS 0.009315f
C1066 B.n602 VSUBS 0.009315f
C1067 B.n603 VSUBS 0.009315f
C1068 B.n604 VSUBS 0.009315f
C1069 B.n605 VSUBS 0.009315f
C1070 B.n606 VSUBS 0.009315f
C1071 B.n607 VSUBS 0.009315f
C1072 B.n608 VSUBS 0.009315f
C1073 B.n609 VSUBS 0.009315f
C1074 B.n610 VSUBS 0.009315f
C1075 B.n611 VSUBS 0.009315f
C1076 B.n612 VSUBS 0.009315f
C1077 B.n613 VSUBS 0.022709f
C1078 B.n614 VSUBS 0.022709f
C1079 B.n615 VSUBS 0.022222f
C1080 B.n616 VSUBS 0.009315f
C1081 B.n617 VSUBS 0.009315f
C1082 B.n618 VSUBS 0.009315f
C1083 B.n619 VSUBS 0.009315f
C1084 B.n620 VSUBS 0.009315f
C1085 B.n621 VSUBS 0.009315f
C1086 B.n622 VSUBS 0.009315f
C1087 B.n623 VSUBS 0.009315f
C1088 B.n624 VSUBS 0.009315f
C1089 B.n625 VSUBS 0.009315f
C1090 B.n626 VSUBS 0.009315f
C1091 B.n627 VSUBS 0.009315f
C1092 B.n628 VSUBS 0.009315f
C1093 B.n629 VSUBS 0.009315f
C1094 B.n630 VSUBS 0.009315f
C1095 B.n631 VSUBS 0.009315f
C1096 B.n632 VSUBS 0.009315f
C1097 B.n633 VSUBS 0.009315f
C1098 B.n634 VSUBS 0.009315f
C1099 B.n635 VSUBS 0.009315f
C1100 B.n636 VSUBS 0.009315f
C1101 B.n637 VSUBS 0.009315f
C1102 B.n638 VSUBS 0.009315f
C1103 B.n639 VSUBS 0.009315f
C1104 B.n640 VSUBS 0.009315f
C1105 B.n641 VSUBS 0.009315f
C1106 B.n642 VSUBS 0.009315f
C1107 B.n643 VSUBS 0.009315f
C1108 B.n644 VSUBS 0.009315f
C1109 B.n645 VSUBS 0.009315f
C1110 B.n646 VSUBS 0.009315f
C1111 B.n647 VSUBS 0.009315f
C1112 B.n648 VSUBS 0.009315f
C1113 B.n649 VSUBS 0.009315f
C1114 B.n650 VSUBS 0.009315f
C1115 B.n651 VSUBS 0.009315f
C1116 B.n652 VSUBS 0.009315f
C1117 B.n653 VSUBS 0.009315f
C1118 B.n654 VSUBS 0.009315f
C1119 B.n655 VSUBS 0.009315f
C1120 B.n656 VSUBS 0.009315f
C1121 B.n657 VSUBS 0.009315f
C1122 B.n658 VSUBS 0.009315f
C1123 B.n659 VSUBS 0.009315f
C1124 B.n660 VSUBS 0.009315f
C1125 B.n661 VSUBS 0.009315f
C1126 B.n662 VSUBS 0.009315f
C1127 B.n663 VSUBS 0.009315f
C1128 B.n664 VSUBS 0.009315f
C1129 B.n665 VSUBS 0.009315f
C1130 B.n666 VSUBS 0.009315f
C1131 B.n667 VSUBS 0.009315f
C1132 B.n668 VSUBS 0.009315f
C1133 B.n669 VSUBS 0.009315f
C1134 B.n670 VSUBS 0.009315f
C1135 B.n671 VSUBS 0.009315f
C1136 B.n672 VSUBS 0.009315f
C1137 B.n673 VSUBS 0.009315f
C1138 B.n674 VSUBS 0.009315f
C1139 B.n675 VSUBS 0.009315f
C1140 B.n676 VSUBS 0.009315f
C1141 B.n677 VSUBS 0.009315f
C1142 B.n678 VSUBS 0.009315f
C1143 B.n679 VSUBS 0.009315f
C1144 B.n680 VSUBS 0.009315f
C1145 B.n681 VSUBS 0.009315f
C1146 B.n682 VSUBS 0.009315f
C1147 B.n683 VSUBS 0.009315f
C1148 B.n684 VSUBS 0.009315f
C1149 B.n685 VSUBS 0.009315f
C1150 B.n686 VSUBS 0.009315f
C1151 B.n687 VSUBS 0.009315f
C1152 B.n688 VSUBS 0.009315f
C1153 B.n689 VSUBS 0.009315f
C1154 B.n690 VSUBS 0.009315f
C1155 B.n691 VSUBS 0.009315f
C1156 B.n692 VSUBS 0.009315f
C1157 B.n693 VSUBS 0.009315f
C1158 B.n694 VSUBS 0.009315f
C1159 B.n695 VSUBS 0.021093f
.ends

