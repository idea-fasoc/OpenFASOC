* NGSPICE file created from diff_pair_sample_1599.ext - technology: sky130A

.subckt diff_pair_sample_1599 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=0 ps=0 w=15.86 l=2.62
X1 VDD1.t9 VP.t0 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=6.1854 ps=32.5 w=15.86 l=2.62
X2 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=0 ps=0 w=15.86 l=2.62
X3 VDD1.t8 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X4 VTAIL.t7 VN.t0 VDD2.t9 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X5 VTAIL.t6 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X6 VTAIL.t5 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X7 VDD2.t6 VN.t3 VTAIL.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=2.6169 ps=16.19 w=15.86 l=2.62
X8 VDD1.t7 VP.t2 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=2.6169 ps=16.19 w=15.86 l=2.62
X9 VTAIL.t19 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X10 VDD1.t5 VP.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X11 VDD2.t5 VN.t4 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=2.6169 ps=16.19 w=15.86 l=2.62
X12 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=0 ps=0 w=15.86 l=2.62
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=0 ps=0 w=15.86 l=2.62
X14 VDD1.t4 VP.t5 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=6.1854 ps=32.5 w=15.86 l=2.62
X15 VDD1.t3 VP.t6 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=6.1854 pd=32.5 as=2.6169 ps=16.19 w=15.86 l=2.62
X16 VDD2.t4 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X17 VTAIL.t18 VP.t7 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X18 VDD2.t3 VN.t6 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=6.1854 ps=32.5 w=15.86 l=2.62
X19 VDD2.t2 VN.t7 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X20 VDD2.t1 VN.t8 VTAIL.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=6.1854 ps=32.5 w=15.86 l=2.62
X21 VTAIL.t10 VP.t8 VDD1.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X22 VTAIL.t0 VN.t9 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
X23 VTAIL.t15 VP.t9 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6169 pd=16.19 as=2.6169 ps=16.19 w=15.86 l=2.62
R0 B.n1072 B.n1071 585
R1 B.n401 B.n168 585
R2 B.n400 B.n399 585
R3 B.n398 B.n397 585
R4 B.n396 B.n395 585
R5 B.n394 B.n393 585
R6 B.n392 B.n391 585
R7 B.n390 B.n389 585
R8 B.n388 B.n387 585
R9 B.n386 B.n385 585
R10 B.n384 B.n383 585
R11 B.n382 B.n381 585
R12 B.n380 B.n379 585
R13 B.n378 B.n377 585
R14 B.n376 B.n375 585
R15 B.n374 B.n373 585
R16 B.n372 B.n371 585
R17 B.n370 B.n369 585
R18 B.n368 B.n367 585
R19 B.n366 B.n365 585
R20 B.n364 B.n363 585
R21 B.n362 B.n361 585
R22 B.n360 B.n359 585
R23 B.n358 B.n357 585
R24 B.n356 B.n355 585
R25 B.n354 B.n353 585
R26 B.n352 B.n351 585
R27 B.n350 B.n349 585
R28 B.n348 B.n347 585
R29 B.n346 B.n345 585
R30 B.n344 B.n343 585
R31 B.n342 B.n341 585
R32 B.n340 B.n339 585
R33 B.n338 B.n337 585
R34 B.n336 B.n335 585
R35 B.n334 B.n333 585
R36 B.n332 B.n331 585
R37 B.n330 B.n329 585
R38 B.n328 B.n327 585
R39 B.n326 B.n325 585
R40 B.n324 B.n323 585
R41 B.n322 B.n321 585
R42 B.n320 B.n319 585
R43 B.n318 B.n317 585
R44 B.n316 B.n315 585
R45 B.n314 B.n313 585
R46 B.n312 B.n311 585
R47 B.n310 B.n309 585
R48 B.n308 B.n307 585
R49 B.n306 B.n305 585
R50 B.n304 B.n303 585
R51 B.n302 B.n301 585
R52 B.n300 B.n299 585
R53 B.n297 B.n296 585
R54 B.n295 B.n294 585
R55 B.n293 B.n292 585
R56 B.n291 B.n290 585
R57 B.n289 B.n288 585
R58 B.n287 B.n286 585
R59 B.n285 B.n284 585
R60 B.n283 B.n282 585
R61 B.n281 B.n280 585
R62 B.n279 B.n278 585
R63 B.n276 B.n275 585
R64 B.n274 B.n273 585
R65 B.n272 B.n271 585
R66 B.n270 B.n269 585
R67 B.n268 B.n267 585
R68 B.n266 B.n265 585
R69 B.n264 B.n263 585
R70 B.n262 B.n261 585
R71 B.n260 B.n259 585
R72 B.n258 B.n257 585
R73 B.n256 B.n255 585
R74 B.n254 B.n253 585
R75 B.n252 B.n251 585
R76 B.n250 B.n249 585
R77 B.n248 B.n247 585
R78 B.n246 B.n245 585
R79 B.n244 B.n243 585
R80 B.n242 B.n241 585
R81 B.n240 B.n239 585
R82 B.n238 B.n237 585
R83 B.n236 B.n235 585
R84 B.n234 B.n233 585
R85 B.n232 B.n231 585
R86 B.n230 B.n229 585
R87 B.n228 B.n227 585
R88 B.n226 B.n225 585
R89 B.n224 B.n223 585
R90 B.n222 B.n221 585
R91 B.n220 B.n219 585
R92 B.n218 B.n217 585
R93 B.n216 B.n215 585
R94 B.n214 B.n213 585
R95 B.n212 B.n211 585
R96 B.n210 B.n209 585
R97 B.n208 B.n207 585
R98 B.n206 B.n205 585
R99 B.n204 B.n203 585
R100 B.n202 B.n201 585
R101 B.n200 B.n199 585
R102 B.n198 B.n197 585
R103 B.n196 B.n195 585
R104 B.n194 B.n193 585
R105 B.n192 B.n191 585
R106 B.n190 B.n189 585
R107 B.n188 B.n187 585
R108 B.n186 B.n185 585
R109 B.n184 B.n183 585
R110 B.n182 B.n181 585
R111 B.n180 B.n179 585
R112 B.n178 B.n177 585
R113 B.n176 B.n175 585
R114 B.n174 B.n173 585
R115 B.n109 B.n108 585
R116 B.n1070 B.n110 585
R117 B.n1075 B.n110 585
R118 B.n1069 B.n1068 585
R119 B.n1068 B.n106 585
R120 B.n1067 B.n105 585
R121 B.n1081 B.n105 585
R122 B.n1066 B.n104 585
R123 B.n1082 B.n104 585
R124 B.n1065 B.n103 585
R125 B.n1083 B.n103 585
R126 B.n1064 B.n1063 585
R127 B.n1063 B.n99 585
R128 B.n1062 B.n98 585
R129 B.n1089 B.n98 585
R130 B.n1061 B.n97 585
R131 B.n1090 B.n97 585
R132 B.n1060 B.n96 585
R133 B.n1091 B.n96 585
R134 B.n1059 B.n1058 585
R135 B.n1058 B.n92 585
R136 B.n1057 B.n91 585
R137 B.n1097 B.n91 585
R138 B.n1056 B.n90 585
R139 B.n1098 B.n90 585
R140 B.n1055 B.n89 585
R141 B.n1099 B.n89 585
R142 B.n1054 B.n1053 585
R143 B.n1053 B.n85 585
R144 B.n1052 B.n84 585
R145 B.n1105 B.n84 585
R146 B.n1051 B.n83 585
R147 B.n1106 B.n83 585
R148 B.n1050 B.n82 585
R149 B.n1107 B.n82 585
R150 B.n1049 B.n1048 585
R151 B.n1048 B.n78 585
R152 B.n1047 B.n77 585
R153 B.n1113 B.n77 585
R154 B.n1046 B.n76 585
R155 B.n1114 B.n76 585
R156 B.n1045 B.n75 585
R157 B.n1115 B.n75 585
R158 B.n1044 B.n1043 585
R159 B.n1043 B.n71 585
R160 B.n1042 B.n70 585
R161 B.n1121 B.n70 585
R162 B.n1041 B.n69 585
R163 B.n1122 B.n69 585
R164 B.n1040 B.n68 585
R165 B.n1123 B.n68 585
R166 B.n1039 B.n1038 585
R167 B.n1038 B.n64 585
R168 B.n1037 B.n63 585
R169 B.n1129 B.n63 585
R170 B.n1036 B.n62 585
R171 B.n1130 B.n62 585
R172 B.n1035 B.n61 585
R173 B.n1131 B.n61 585
R174 B.n1034 B.n1033 585
R175 B.n1033 B.n57 585
R176 B.n1032 B.n56 585
R177 B.n1137 B.n56 585
R178 B.n1031 B.n55 585
R179 B.n1138 B.n55 585
R180 B.n1030 B.n54 585
R181 B.n1139 B.n54 585
R182 B.n1029 B.n1028 585
R183 B.n1028 B.n50 585
R184 B.n1027 B.n49 585
R185 B.n1145 B.n49 585
R186 B.n1026 B.n48 585
R187 B.n1146 B.n48 585
R188 B.n1025 B.n47 585
R189 B.n1147 B.n47 585
R190 B.n1024 B.n1023 585
R191 B.n1023 B.n43 585
R192 B.n1022 B.n42 585
R193 B.n1153 B.n42 585
R194 B.n1021 B.n41 585
R195 B.n1154 B.n41 585
R196 B.n1020 B.n40 585
R197 B.n1155 B.n40 585
R198 B.n1019 B.n1018 585
R199 B.n1018 B.n36 585
R200 B.n1017 B.n35 585
R201 B.n1161 B.n35 585
R202 B.n1016 B.n34 585
R203 B.n1162 B.n34 585
R204 B.n1015 B.n33 585
R205 B.n1163 B.n33 585
R206 B.n1014 B.n1013 585
R207 B.n1013 B.n32 585
R208 B.n1012 B.n28 585
R209 B.n1169 B.n28 585
R210 B.n1011 B.n27 585
R211 B.n1170 B.n27 585
R212 B.n1010 B.n26 585
R213 B.n1171 B.n26 585
R214 B.n1009 B.n1008 585
R215 B.n1008 B.n22 585
R216 B.n1007 B.n21 585
R217 B.n1177 B.n21 585
R218 B.n1006 B.n20 585
R219 B.n1178 B.n20 585
R220 B.n1005 B.n19 585
R221 B.n1179 B.n19 585
R222 B.n1004 B.n1003 585
R223 B.n1003 B.n15 585
R224 B.n1002 B.n14 585
R225 B.n1185 B.n14 585
R226 B.n1001 B.n13 585
R227 B.n1186 B.n13 585
R228 B.n1000 B.n12 585
R229 B.n1187 B.n12 585
R230 B.n999 B.n998 585
R231 B.n998 B.n8 585
R232 B.n997 B.n7 585
R233 B.n1193 B.n7 585
R234 B.n996 B.n6 585
R235 B.n1194 B.n6 585
R236 B.n995 B.n5 585
R237 B.n1195 B.n5 585
R238 B.n994 B.n993 585
R239 B.n993 B.n4 585
R240 B.n992 B.n402 585
R241 B.n992 B.n991 585
R242 B.n982 B.n403 585
R243 B.n404 B.n403 585
R244 B.n984 B.n983 585
R245 B.n985 B.n984 585
R246 B.n981 B.n409 585
R247 B.n409 B.n408 585
R248 B.n980 B.n979 585
R249 B.n979 B.n978 585
R250 B.n411 B.n410 585
R251 B.n412 B.n411 585
R252 B.n971 B.n970 585
R253 B.n972 B.n971 585
R254 B.n969 B.n417 585
R255 B.n417 B.n416 585
R256 B.n968 B.n967 585
R257 B.n967 B.n966 585
R258 B.n419 B.n418 585
R259 B.n420 B.n419 585
R260 B.n959 B.n958 585
R261 B.n960 B.n959 585
R262 B.n957 B.n425 585
R263 B.n425 B.n424 585
R264 B.n956 B.n955 585
R265 B.n955 B.n954 585
R266 B.n427 B.n426 585
R267 B.n947 B.n427 585
R268 B.n946 B.n945 585
R269 B.n948 B.n946 585
R270 B.n944 B.n432 585
R271 B.n432 B.n431 585
R272 B.n943 B.n942 585
R273 B.n942 B.n941 585
R274 B.n434 B.n433 585
R275 B.n435 B.n434 585
R276 B.n934 B.n933 585
R277 B.n935 B.n934 585
R278 B.n932 B.n440 585
R279 B.n440 B.n439 585
R280 B.n931 B.n930 585
R281 B.n930 B.n929 585
R282 B.n442 B.n441 585
R283 B.n443 B.n442 585
R284 B.n922 B.n921 585
R285 B.n923 B.n922 585
R286 B.n920 B.n448 585
R287 B.n448 B.n447 585
R288 B.n919 B.n918 585
R289 B.n918 B.n917 585
R290 B.n450 B.n449 585
R291 B.n451 B.n450 585
R292 B.n910 B.n909 585
R293 B.n911 B.n910 585
R294 B.n908 B.n456 585
R295 B.n456 B.n455 585
R296 B.n907 B.n906 585
R297 B.n906 B.n905 585
R298 B.n458 B.n457 585
R299 B.n459 B.n458 585
R300 B.n898 B.n897 585
R301 B.n899 B.n898 585
R302 B.n896 B.n464 585
R303 B.n464 B.n463 585
R304 B.n895 B.n894 585
R305 B.n894 B.n893 585
R306 B.n466 B.n465 585
R307 B.n467 B.n466 585
R308 B.n886 B.n885 585
R309 B.n887 B.n886 585
R310 B.n884 B.n472 585
R311 B.n472 B.n471 585
R312 B.n883 B.n882 585
R313 B.n882 B.n881 585
R314 B.n474 B.n473 585
R315 B.n475 B.n474 585
R316 B.n874 B.n873 585
R317 B.n875 B.n874 585
R318 B.n872 B.n479 585
R319 B.n483 B.n479 585
R320 B.n871 B.n870 585
R321 B.n870 B.n869 585
R322 B.n481 B.n480 585
R323 B.n482 B.n481 585
R324 B.n862 B.n861 585
R325 B.n863 B.n862 585
R326 B.n860 B.n488 585
R327 B.n488 B.n487 585
R328 B.n859 B.n858 585
R329 B.n858 B.n857 585
R330 B.n490 B.n489 585
R331 B.n491 B.n490 585
R332 B.n850 B.n849 585
R333 B.n851 B.n850 585
R334 B.n848 B.n496 585
R335 B.n496 B.n495 585
R336 B.n847 B.n846 585
R337 B.n846 B.n845 585
R338 B.n498 B.n497 585
R339 B.n499 B.n498 585
R340 B.n838 B.n837 585
R341 B.n839 B.n838 585
R342 B.n836 B.n503 585
R343 B.n507 B.n503 585
R344 B.n835 B.n834 585
R345 B.n834 B.n833 585
R346 B.n505 B.n504 585
R347 B.n506 B.n505 585
R348 B.n826 B.n825 585
R349 B.n827 B.n826 585
R350 B.n824 B.n512 585
R351 B.n512 B.n511 585
R352 B.n823 B.n822 585
R353 B.n822 B.n821 585
R354 B.n514 B.n513 585
R355 B.n515 B.n514 585
R356 B.n814 B.n813 585
R357 B.n815 B.n814 585
R358 B.n518 B.n517 585
R359 B.n585 B.n584 585
R360 B.n586 B.n582 585
R361 B.n582 B.n519 585
R362 B.n588 B.n587 585
R363 B.n590 B.n581 585
R364 B.n593 B.n592 585
R365 B.n594 B.n580 585
R366 B.n596 B.n595 585
R367 B.n598 B.n579 585
R368 B.n601 B.n600 585
R369 B.n602 B.n578 585
R370 B.n604 B.n603 585
R371 B.n606 B.n577 585
R372 B.n609 B.n608 585
R373 B.n610 B.n576 585
R374 B.n612 B.n611 585
R375 B.n614 B.n575 585
R376 B.n617 B.n616 585
R377 B.n618 B.n574 585
R378 B.n620 B.n619 585
R379 B.n622 B.n573 585
R380 B.n625 B.n624 585
R381 B.n626 B.n572 585
R382 B.n628 B.n627 585
R383 B.n630 B.n571 585
R384 B.n633 B.n632 585
R385 B.n634 B.n570 585
R386 B.n636 B.n635 585
R387 B.n638 B.n569 585
R388 B.n641 B.n640 585
R389 B.n642 B.n568 585
R390 B.n644 B.n643 585
R391 B.n646 B.n567 585
R392 B.n649 B.n648 585
R393 B.n650 B.n566 585
R394 B.n652 B.n651 585
R395 B.n654 B.n565 585
R396 B.n657 B.n656 585
R397 B.n658 B.n564 585
R398 B.n660 B.n659 585
R399 B.n662 B.n563 585
R400 B.n665 B.n664 585
R401 B.n666 B.n562 585
R402 B.n668 B.n667 585
R403 B.n670 B.n561 585
R404 B.n673 B.n672 585
R405 B.n674 B.n560 585
R406 B.n676 B.n675 585
R407 B.n678 B.n559 585
R408 B.n681 B.n680 585
R409 B.n682 B.n558 585
R410 B.n684 B.n683 585
R411 B.n686 B.n557 585
R412 B.n689 B.n688 585
R413 B.n690 B.n553 585
R414 B.n692 B.n691 585
R415 B.n694 B.n552 585
R416 B.n697 B.n696 585
R417 B.n698 B.n551 585
R418 B.n700 B.n699 585
R419 B.n702 B.n550 585
R420 B.n705 B.n704 585
R421 B.n706 B.n547 585
R422 B.n709 B.n708 585
R423 B.n711 B.n546 585
R424 B.n714 B.n713 585
R425 B.n715 B.n545 585
R426 B.n717 B.n716 585
R427 B.n719 B.n544 585
R428 B.n722 B.n721 585
R429 B.n723 B.n543 585
R430 B.n725 B.n724 585
R431 B.n727 B.n542 585
R432 B.n730 B.n729 585
R433 B.n731 B.n541 585
R434 B.n733 B.n732 585
R435 B.n735 B.n540 585
R436 B.n738 B.n737 585
R437 B.n739 B.n539 585
R438 B.n741 B.n740 585
R439 B.n743 B.n538 585
R440 B.n746 B.n745 585
R441 B.n747 B.n537 585
R442 B.n749 B.n748 585
R443 B.n751 B.n536 585
R444 B.n754 B.n753 585
R445 B.n755 B.n535 585
R446 B.n757 B.n756 585
R447 B.n759 B.n534 585
R448 B.n762 B.n761 585
R449 B.n763 B.n533 585
R450 B.n765 B.n764 585
R451 B.n767 B.n532 585
R452 B.n770 B.n769 585
R453 B.n771 B.n531 585
R454 B.n773 B.n772 585
R455 B.n775 B.n530 585
R456 B.n778 B.n777 585
R457 B.n779 B.n529 585
R458 B.n781 B.n780 585
R459 B.n783 B.n528 585
R460 B.n786 B.n785 585
R461 B.n787 B.n527 585
R462 B.n789 B.n788 585
R463 B.n791 B.n526 585
R464 B.n794 B.n793 585
R465 B.n795 B.n525 585
R466 B.n797 B.n796 585
R467 B.n799 B.n524 585
R468 B.n802 B.n801 585
R469 B.n803 B.n523 585
R470 B.n805 B.n804 585
R471 B.n807 B.n522 585
R472 B.n808 B.n521 585
R473 B.n811 B.n810 585
R474 B.n812 B.n520 585
R475 B.n520 B.n519 585
R476 B.n817 B.n816 585
R477 B.n816 B.n815 585
R478 B.n818 B.n516 585
R479 B.n516 B.n515 585
R480 B.n820 B.n819 585
R481 B.n821 B.n820 585
R482 B.n510 B.n509 585
R483 B.n511 B.n510 585
R484 B.n829 B.n828 585
R485 B.n828 B.n827 585
R486 B.n830 B.n508 585
R487 B.n508 B.n506 585
R488 B.n832 B.n831 585
R489 B.n833 B.n832 585
R490 B.n502 B.n501 585
R491 B.n507 B.n502 585
R492 B.n841 B.n840 585
R493 B.n840 B.n839 585
R494 B.n842 B.n500 585
R495 B.n500 B.n499 585
R496 B.n844 B.n843 585
R497 B.n845 B.n844 585
R498 B.n494 B.n493 585
R499 B.n495 B.n494 585
R500 B.n853 B.n852 585
R501 B.n852 B.n851 585
R502 B.n854 B.n492 585
R503 B.n492 B.n491 585
R504 B.n856 B.n855 585
R505 B.n857 B.n856 585
R506 B.n486 B.n485 585
R507 B.n487 B.n486 585
R508 B.n865 B.n864 585
R509 B.n864 B.n863 585
R510 B.n866 B.n484 585
R511 B.n484 B.n482 585
R512 B.n868 B.n867 585
R513 B.n869 B.n868 585
R514 B.n478 B.n477 585
R515 B.n483 B.n478 585
R516 B.n877 B.n876 585
R517 B.n876 B.n875 585
R518 B.n878 B.n476 585
R519 B.n476 B.n475 585
R520 B.n880 B.n879 585
R521 B.n881 B.n880 585
R522 B.n470 B.n469 585
R523 B.n471 B.n470 585
R524 B.n889 B.n888 585
R525 B.n888 B.n887 585
R526 B.n890 B.n468 585
R527 B.n468 B.n467 585
R528 B.n892 B.n891 585
R529 B.n893 B.n892 585
R530 B.n462 B.n461 585
R531 B.n463 B.n462 585
R532 B.n901 B.n900 585
R533 B.n900 B.n899 585
R534 B.n902 B.n460 585
R535 B.n460 B.n459 585
R536 B.n904 B.n903 585
R537 B.n905 B.n904 585
R538 B.n454 B.n453 585
R539 B.n455 B.n454 585
R540 B.n913 B.n912 585
R541 B.n912 B.n911 585
R542 B.n914 B.n452 585
R543 B.n452 B.n451 585
R544 B.n916 B.n915 585
R545 B.n917 B.n916 585
R546 B.n446 B.n445 585
R547 B.n447 B.n446 585
R548 B.n925 B.n924 585
R549 B.n924 B.n923 585
R550 B.n926 B.n444 585
R551 B.n444 B.n443 585
R552 B.n928 B.n927 585
R553 B.n929 B.n928 585
R554 B.n438 B.n437 585
R555 B.n439 B.n438 585
R556 B.n937 B.n936 585
R557 B.n936 B.n935 585
R558 B.n938 B.n436 585
R559 B.n436 B.n435 585
R560 B.n940 B.n939 585
R561 B.n941 B.n940 585
R562 B.n430 B.n429 585
R563 B.n431 B.n430 585
R564 B.n950 B.n949 585
R565 B.n949 B.n948 585
R566 B.n951 B.n428 585
R567 B.n947 B.n428 585
R568 B.n953 B.n952 585
R569 B.n954 B.n953 585
R570 B.n423 B.n422 585
R571 B.n424 B.n423 585
R572 B.n962 B.n961 585
R573 B.n961 B.n960 585
R574 B.n963 B.n421 585
R575 B.n421 B.n420 585
R576 B.n965 B.n964 585
R577 B.n966 B.n965 585
R578 B.n415 B.n414 585
R579 B.n416 B.n415 585
R580 B.n974 B.n973 585
R581 B.n973 B.n972 585
R582 B.n975 B.n413 585
R583 B.n413 B.n412 585
R584 B.n977 B.n976 585
R585 B.n978 B.n977 585
R586 B.n407 B.n406 585
R587 B.n408 B.n407 585
R588 B.n987 B.n986 585
R589 B.n986 B.n985 585
R590 B.n988 B.n405 585
R591 B.n405 B.n404 585
R592 B.n990 B.n989 585
R593 B.n991 B.n990 585
R594 B.n2 B.n0 585
R595 B.n4 B.n2 585
R596 B.n3 B.n1 585
R597 B.n1194 B.n3 585
R598 B.n1192 B.n1191 585
R599 B.n1193 B.n1192 585
R600 B.n1190 B.n9 585
R601 B.n9 B.n8 585
R602 B.n1189 B.n1188 585
R603 B.n1188 B.n1187 585
R604 B.n11 B.n10 585
R605 B.n1186 B.n11 585
R606 B.n1184 B.n1183 585
R607 B.n1185 B.n1184 585
R608 B.n1182 B.n16 585
R609 B.n16 B.n15 585
R610 B.n1181 B.n1180 585
R611 B.n1180 B.n1179 585
R612 B.n18 B.n17 585
R613 B.n1178 B.n18 585
R614 B.n1176 B.n1175 585
R615 B.n1177 B.n1176 585
R616 B.n1174 B.n23 585
R617 B.n23 B.n22 585
R618 B.n1173 B.n1172 585
R619 B.n1172 B.n1171 585
R620 B.n25 B.n24 585
R621 B.n1170 B.n25 585
R622 B.n1168 B.n1167 585
R623 B.n1169 B.n1168 585
R624 B.n1166 B.n29 585
R625 B.n32 B.n29 585
R626 B.n1165 B.n1164 585
R627 B.n1164 B.n1163 585
R628 B.n31 B.n30 585
R629 B.n1162 B.n31 585
R630 B.n1160 B.n1159 585
R631 B.n1161 B.n1160 585
R632 B.n1158 B.n37 585
R633 B.n37 B.n36 585
R634 B.n1157 B.n1156 585
R635 B.n1156 B.n1155 585
R636 B.n39 B.n38 585
R637 B.n1154 B.n39 585
R638 B.n1152 B.n1151 585
R639 B.n1153 B.n1152 585
R640 B.n1150 B.n44 585
R641 B.n44 B.n43 585
R642 B.n1149 B.n1148 585
R643 B.n1148 B.n1147 585
R644 B.n46 B.n45 585
R645 B.n1146 B.n46 585
R646 B.n1144 B.n1143 585
R647 B.n1145 B.n1144 585
R648 B.n1142 B.n51 585
R649 B.n51 B.n50 585
R650 B.n1141 B.n1140 585
R651 B.n1140 B.n1139 585
R652 B.n53 B.n52 585
R653 B.n1138 B.n53 585
R654 B.n1136 B.n1135 585
R655 B.n1137 B.n1136 585
R656 B.n1134 B.n58 585
R657 B.n58 B.n57 585
R658 B.n1133 B.n1132 585
R659 B.n1132 B.n1131 585
R660 B.n60 B.n59 585
R661 B.n1130 B.n60 585
R662 B.n1128 B.n1127 585
R663 B.n1129 B.n1128 585
R664 B.n1126 B.n65 585
R665 B.n65 B.n64 585
R666 B.n1125 B.n1124 585
R667 B.n1124 B.n1123 585
R668 B.n67 B.n66 585
R669 B.n1122 B.n67 585
R670 B.n1120 B.n1119 585
R671 B.n1121 B.n1120 585
R672 B.n1118 B.n72 585
R673 B.n72 B.n71 585
R674 B.n1117 B.n1116 585
R675 B.n1116 B.n1115 585
R676 B.n74 B.n73 585
R677 B.n1114 B.n74 585
R678 B.n1112 B.n1111 585
R679 B.n1113 B.n1112 585
R680 B.n1110 B.n79 585
R681 B.n79 B.n78 585
R682 B.n1109 B.n1108 585
R683 B.n1108 B.n1107 585
R684 B.n81 B.n80 585
R685 B.n1106 B.n81 585
R686 B.n1104 B.n1103 585
R687 B.n1105 B.n1104 585
R688 B.n1102 B.n86 585
R689 B.n86 B.n85 585
R690 B.n1101 B.n1100 585
R691 B.n1100 B.n1099 585
R692 B.n88 B.n87 585
R693 B.n1098 B.n88 585
R694 B.n1096 B.n1095 585
R695 B.n1097 B.n1096 585
R696 B.n1094 B.n93 585
R697 B.n93 B.n92 585
R698 B.n1093 B.n1092 585
R699 B.n1092 B.n1091 585
R700 B.n95 B.n94 585
R701 B.n1090 B.n95 585
R702 B.n1088 B.n1087 585
R703 B.n1089 B.n1088 585
R704 B.n1086 B.n100 585
R705 B.n100 B.n99 585
R706 B.n1085 B.n1084 585
R707 B.n1084 B.n1083 585
R708 B.n102 B.n101 585
R709 B.n1082 B.n102 585
R710 B.n1080 B.n1079 585
R711 B.n1081 B.n1080 585
R712 B.n1078 B.n107 585
R713 B.n107 B.n106 585
R714 B.n1077 B.n1076 585
R715 B.n1076 B.n1075 585
R716 B.n1197 B.n1196 585
R717 B.n1196 B.n1195 585
R718 B.n816 B.n518 487.695
R719 B.n1076 B.n109 487.695
R720 B.n814 B.n520 487.695
R721 B.n1072 B.n110 487.695
R722 B.n548 B.t17 353.964
R723 B.n554 B.t21 353.964
R724 B.n171 B.t10 353.964
R725 B.n169 B.t14 353.964
R726 B.n1074 B.n1073 256.663
R727 B.n1074 B.n167 256.663
R728 B.n1074 B.n166 256.663
R729 B.n1074 B.n165 256.663
R730 B.n1074 B.n164 256.663
R731 B.n1074 B.n163 256.663
R732 B.n1074 B.n162 256.663
R733 B.n1074 B.n161 256.663
R734 B.n1074 B.n160 256.663
R735 B.n1074 B.n159 256.663
R736 B.n1074 B.n158 256.663
R737 B.n1074 B.n157 256.663
R738 B.n1074 B.n156 256.663
R739 B.n1074 B.n155 256.663
R740 B.n1074 B.n154 256.663
R741 B.n1074 B.n153 256.663
R742 B.n1074 B.n152 256.663
R743 B.n1074 B.n151 256.663
R744 B.n1074 B.n150 256.663
R745 B.n1074 B.n149 256.663
R746 B.n1074 B.n148 256.663
R747 B.n1074 B.n147 256.663
R748 B.n1074 B.n146 256.663
R749 B.n1074 B.n145 256.663
R750 B.n1074 B.n144 256.663
R751 B.n1074 B.n143 256.663
R752 B.n1074 B.n142 256.663
R753 B.n1074 B.n141 256.663
R754 B.n1074 B.n140 256.663
R755 B.n1074 B.n139 256.663
R756 B.n1074 B.n138 256.663
R757 B.n1074 B.n137 256.663
R758 B.n1074 B.n136 256.663
R759 B.n1074 B.n135 256.663
R760 B.n1074 B.n134 256.663
R761 B.n1074 B.n133 256.663
R762 B.n1074 B.n132 256.663
R763 B.n1074 B.n131 256.663
R764 B.n1074 B.n130 256.663
R765 B.n1074 B.n129 256.663
R766 B.n1074 B.n128 256.663
R767 B.n1074 B.n127 256.663
R768 B.n1074 B.n126 256.663
R769 B.n1074 B.n125 256.663
R770 B.n1074 B.n124 256.663
R771 B.n1074 B.n123 256.663
R772 B.n1074 B.n122 256.663
R773 B.n1074 B.n121 256.663
R774 B.n1074 B.n120 256.663
R775 B.n1074 B.n119 256.663
R776 B.n1074 B.n118 256.663
R777 B.n1074 B.n117 256.663
R778 B.n1074 B.n116 256.663
R779 B.n1074 B.n115 256.663
R780 B.n1074 B.n114 256.663
R781 B.n1074 B.n113 256.663
R782 B.n1074 B.n112 256.663
R783 B.n1074 B.n111 256.663
R784 B.n583 B.n519 256.663
R785 B.n589 B.n519 256.663
R786 B.n591 B.n519 256.663
R787 B.n597 B.n519 256.663
R788 B.n599 B.n519 256.663
R789 B.n605 B.n519 256.663
R790 B.n607 B.n519 256.663
R791 B.n613 B.n519 256.663
R792 B.n615 B.n519 256.663
R793 B.n621 B.n519 256.663
R794 B.n623 B.n519 256.663
R795 B.n629 B.n519 256.663
R796 B.n631 B.n519 256.663
R797 B.n637 B.n519 256.663
R798 B.n639 B.n519 256.663
R799 B.n645 B.n519 256.663
R800 B.n647 B.n519 256.663
R801 B.n653 B.n519 256.663
R802 B.n655 B.n519 256.663
R803 B.n661 B.n519 256.663
R804 B.n663 B.n519 256.663
R805 B.n669 B.n519 256.663
R806 B.n671 B.n519 256.663
R807 B.n677 B.n519 256.663
R808 B.n679 B.n519 256.663
R809 B.n685 B.n519 256.663
R810 B.n687 B.n519 256.663
R811 B.n693 B.n519 256.663
R812 B.n695 B.n519 256.663
R813 B.n701 B.n519 256.663
R814 B.n703 B.n519 256.663
R815 B.n710 B.n519 256.663
R816 B.n712 B.n519 256.663
R817 B.n718 B.n519 256.663
R818 B.n720 B.n519 256.663
R819 B.n726 B.n519 256.663
R820 B.n728 B.n519 256.663
R821 B.n734 B.n519 256.663
R822 B.n736 B.n519 256.663
R823 B.n742 B.n519 256.663
R824 B.n744 B.n519 256.663
R825 B.n750 B.n519 256.663
R826 B.n752 B.n519 256.663
R827 B.n758 B.n519 256.663
R828 B.n760 B.n519 256.663
R829 B.n766 B.n519 256.663
R830 B.n768 B.n519 256.663
R831 B.n774 B.n519 256.663
R832 B.n776 B.n519 256.663
R833 B.n782 B.n519 256.663
R834 B.n784 B.n519 256.663
R835 B.n790 B.n519 256.663
R836 B.n792 B.n519 256.663
R837 B.n798 B.n519 256.663
R838 B.n800 B.n519 256.663
R839 B.n806 B.n519 256.663
R840 B.n809 B.n519 256.663
R841 B.n816 B.n516 163.367
R842 B.n820 B.n516 163.367
R843 B.n820 B.n510 163.367
R844 B.n828 B.n510 163.367
R845 B.n828 B.n508 163.367
R846 B.n832 B.n508 163.367
R847 B.n832 B.n502 163.367
R848 B.n840 B.n502 163.367
R849 B.n840 B.n500 163.367
R850 B.n844 B.n500 163.367
R851 B.n844 B.n494 163.367
R852 B.n852 B.n494 163.367
R853 B.n852 B.n492 163.367
R854 B.n856 B.n492 163.367
R855 B.n856 B.n486 163.367
R856 B.n864 B.n486 163.367
R857 B.n864 B.n484 163.367
R858 B.n868 B.n484 163.367
R859 B.n868 B.n478 163.367
R860 B.n876 B.n478 163.367
R861 B.n876 B.n476 163.367
R862 B.n880 B.n476 163.367
R863 B.n880 B.n470 163.367
R864 B.n888 B.n470 163.367
R865 B.n888 B.n468 163.367
R866 B.n892 B.n468 163.367
R867 B.n892 B.n462 163.367
R868 B.n900 B.n462 163.367
R869 B.n900 B.n460 163.367
R870 B.n904 B.n460 163.367
R871 B.n904 B.n454 163.367
R872 B.n912 B.n454 163.367
R873 B.n912 B.n452 163.367
R874 B.n916 B.n452 163.367
R875 B.n916 B.n446 163.367
R876 B.n924 B.n446 163.367
R877 B.n924 B.n444 163.367
R878 B.n928 B.n444 163.367
R879 B.n928 B.n438 163.367
R880 B.n936 B.n438 163.367
R881 B.n936 B.n436 163.367
R882 B.n940 B.n436 163.367
R883 B.n940 B.n430 163.367
R884 B.n949 B.n430 163.367
R885 B.n949 B.n428 163.367
R886 B.n953 B.n428 163.367
R887 B.n953 B.n423 163.367
R888 B.n961 B.n423 163.367
R889 B.n961 B.n421 163.367
R890 B.n965 B.n421 163.367
R891 B.n965 B.n415 163.367
R892 B.n973 B.n415 163.367
R893 B.n973 B.n413 163.367
R894 B.n977 B.n413 163.367
R895 B.n977 B.n407 163.367
R896 B.n986 B.n407 163.367
R897 B.n986 B.n405 163.367
R898 B.n990 B.n405 163.367
R899 B.n990 B.n2 163.367
R900 B.n1196 B.n2 163.367
R901 B.n1196 B.n3 163.367
R902 B.n1192 B.n3 163.367
R903 B.n1192 B.n9 163.367
R904 B.n1188 B.n9 163.367
R905 B.n1188 B.n11 163.367
R906 B.n1184 B.n11 163.367
R907 B.n1184 B.n16 163.367
R908 B.n1180 B.n16 163.367
R909 B.n1180 B.n18 163.367
R910 B.n1176 B.n18 163.367
R911 B.n1176 B.n23 163.367
R912 B.n1172 B.n23 163.367
R913 B.n1172 B.n25 163.367
R914 B.n1168 B.n25 163.367
R915 B.n1168 B.n29 163.367
R916 B.n1164 B.n29 163.367
R917 B.n1164 B.n31 163.367
R918 B.n1160 B.n31 163.367
R919 B.n1160 B.n37 163.367
R920 B.n1156 B.n37 163.367
R921 B.n1156 B.n39 163.367
R922 B.n1152 B.n39 163.367
R923 B.n1152 B.n44 163.367
R924 B.n1148 B.n44 163.367
R925 B.n1148 B.n46 163.367
R926 B.n1144 B.n46 163.367
R927 B.n1144 B.n51 163.367
R928 B.n1140 B.n51 163.367
R929 B.n1140 B.n53 163.367
R930 B.n1136 B.n53 163.367
R931 B.n1136 B.n58 163.367
R932 B.n1132 B.n58 163.367
R933 B.n1132 B.n60 163.367
R934 B.n1128 B.n60 163.367
R935 B.n1128 B.n65 163.367
R936 B.n1124 B.n65 163.367
R937 B.n1124 B.n67 163.367
R938 B.n1120 B.n67 163.367
R939 B.n1120 B.n72 163.367
R940 B.n1116 B.n72 163.367
R941 B.n1116 B.n74 163.367
R942 B.n1112 B.n74 163.367
R943 B.n1112 B.n79 163.367
R944 B.n1108 B.n79 163.367
R945 B.n1108 B.n81 163.367
R946 B.n1104 B.n81 163.367
R947 B.n1104 B.n86 163.367
R948 B.n1100 B.n86 163.367
R949 B.n1100 B.n88 163.367
R950 B.n1096 B.n88 163.367
R951 B.n1096 B.n93 163.367
R952 B.n1092 B.n93 163.367
R953 B.n1092 B.n95 163.367
R954 B.n1088 B.n95 163.367
R955 B.n1088 B.n100 163.367
R956 B.n1084 B.n100 163.367
R957 B.n1084 B.n102 163.367
R958 B.n1080 B.n102 163.367
R959 B.n1080 B.n107 163.367
R960 B.n1076 B.n107 163.367
R961 B.n584 B.n582 163.367
R962 B.n588 B.n582 163.367
R963 B.n592 B.n590 163.367
R964 B.n596 B.n580 163.367
R965 B.n600 B.n598 163.367
R966 B.n604 B.n578 163.367
R967 B.n608 B.n606 163.367
R968 B.n612 B.n576 163.367
R969 B.n616 B.n614 163.367
R970 B.n620 B.n574 163.367
R971 B.n624 B.n622 163.367
R972 B.n628 B.n572 163.367
R973 B.n632 B.n630 163.367
R974 B.n636 B.n570 163.367
R975 B.n640 B.n638 163.367
R976 B.n644 B.n568 163.367
R977 B.n648 B.n646 163.367
R978 B.n652 B.n566 163.367
R979 B.n656 B.n654 163.367
R980 B.n660 B.n564 163.367
R981 B.n664 B.n662 163.367
R982 B.n668 B.n562 163.367
R983 B.n672 B.n670 163.367
R984 B.n676 B.n560 163.367
R985 B.n680 B.n678 163.367
R986 B.n684 B.n558 163.367
R987 B.n688 B.n686 163.367
R988 B.n692 B.n553 163.367
R989 B.n696 B.n694 163.367
R990 B.n700 B.n551 163.367
R991 B.n704 B.n702 163.367
R992 B.n709 B.n547 163.367
R993 B.n713 B.n711 163.367
R994 B.n717 B.n545 163.367
R995 B.n721 B.n719 163.367
R996 B.n725 B.n543 163.367
R997 B.n729 B.n727 163.367
R998 B.n733 B.n541 163.367
R999 B.n737 B.n735 163.367
R1000 B.n741 B.n539 163.367
R1001 B.n745 B.n743 163.367
R1002 B.n749 B.n537 163.367
R1003 B.n753 B.n751 163.367
R1004 B.n757 B.n535 163.367
R1005 B.n761 B.n759 163.367
R1006 B.n765 B.n533 163.367
R1007 B.n769 B.n767 163.367
R1008 B.n773 B.n531 163.367
R1009 B.n777 B.n775 163.367
R1010 B.n781 B.n529 163.367
R1011 B.n785 B.n783 163.367
R1012 B.n789 B.n527 163.367
R1013 B.n793 B.n791 163.367
R1014 B.n797 B.n525 163.367
R1015 B.n801 B.n799 163.367
R1016 B.n805 B.n523 163.367
R1017 B.n808 B.n807 163.367
R1018 B.n810 B.n520 163.367
R1019 B.n814 B.n514 163.367
R1020 B.n822 B.n514 163.367
R1021 B.n822 B.n512 163.367
R1022 B.n826 B.n512 163.367
R1023 B.n826 B.n505 163.367
R1024 B.n834 B.n505 163.367
R1025 B.n834 B.n503 163.367
R1026 B.n838 B.n503 163.367
R1027 B.n838 B.n498 163.367
R1028 B.n846 B.n498 163.367
R1029 B.n846 B.n496 163.367
R1030 B.n850 B.n496 163.367
R1031 B.n850 B.n490 163.367
R1032 B.n858 B.n490 163.367
R1033 B.n858 B.n488 163.367
R1034 B.n862 B.n488 163.367
R1035 B.n862 B.n481 163.367
R1036 B.n870 B.n481 163.367
R1037 B.n870 B.n479 163.367
R1038 B.n874 B.n479 163.367
R1039 B.n874 B.n474 163.367
R1040 B.n882 B.n474 163.367
R1041 B.n882 B.n472 163.367
R1042 B.n886 B.n472 163.367
R1043 B.n886 B.n466 163.367
R1044 B.n894 B.n466 163.367
R1045 B.n894 B.n464 163.367
R1046 B.n898 B.n464 163.367
R1047 B.n898 B.n458 163.367
R1048 B.n906 B.n458 163.367
R1049 B.n906 B.n456 163.367
R1050 B.n910 B.n456 163.367
R1051 B.n910 B.n450 163.367
R1052 B.n918 B.n450 163.367
R1053 B.n918 B.n448 163.367
R1054 B.n922 B.n448 163.367
R1055 B.n922 B.n442 163.367
R1056 B.n930 B.n442 163.367
R1057 B.n930 B.n440 163.367
R1058 B.n934 B.n440 163.367
R1059 B.n934 B.n434 163.367
R1060 B.n942 B.n434 163.367
R1061 B.n942 B.n432 163.367
R1062 B.n946 B.n432 163.367
R1063 B.n946 B.n427 163.367
R1064 B.n955 B.n427 163.367
R1065 B.n955 B.n425 163.367
R1066 B.n959 B.n425 163.367
R1067 B.n959 B.n419 163.367
R1068 B.n967 B.n419 163.367
R1069 B.n967 B.n417 163.367
R1070 B.n971 B.n417 163.367
R1071 B.n971 B.n411 163.367
R1072 B.n979 B.n411 163.367
R1073 B.n979 B.n409 163.367
R1074 B.n984 B.n409 163.367
R1075 B.n984 B.n403 163.367
R1076 B.n992 B.n403 163.367
R1077 B.n993 B.n992 163.367
R1078 B.n993 B.n5 163.367
R1079 B.n6 B.n5 163.367
R1080 B.n7 B.n6 163.367
R1081 B.n998 B.n7 163.367
R1082 B.n998 B.n12 163.367
R1083 B.n13 B.n12 163.367
R1084 B.n14 B.n13 163.367
R1085 B.n1003 B.n14 163.367
R1086 B.n1003 B.n19 163.367
R1087 B.n20 B.n19 163.367
R1088 B.n21 B.n20 163.367
R1089 B.n1008 B.n21 163.367
R1090 B.n1008 B.n26 163.367
R1091 B.n27 B.n26 163.367
R1092 B.n28 B.n27 163.367
R1093 B.n1013 B.n28 163.367
R1094 B.n1013 B.n33 163.367
R1095 B.n34 B.n33 163.367
R1096 B.n35 B.n34 163.367
R1097 B.n1018 B.n35 163.367
R1098 B.n1018 B.n40 163.367
R1099 B.n41 B.n40 163.367
R1100 B.n42 B.n41 163.367
R1101 B.n1023 B.n42 163.367
R1102 B.n1023 B.n47 163.367
R1103 B.n48 B.n47 163.367
R1104 B.n49 B.n48 163.367
R1105 B.n1028 B.n49 163.367
R1106 B.n1028 B.n54 163.367
R1107 B.n55 B.n54 163.367
R1108 B.n56 B.n55 163.367
R1109 B.n1033 B.n56 163.367
R1110 B.n1033 B.n61 163.367
R1111 B.n62 B.n61 163.367
R1112 B.n63 B.n62 163.367
R1113 B.n1038 B.n63 163.367
R1114 B.n1038 B.n68 163.367
R1115 B.n69 B.n68 163.367
R1116 B.n70 B.n69 163.367
R1117 B.n1043 B.n70 163.367
R1118 B.n1043 B.n75 163.367
R1119 B.n76 B.n75 163.367
R1120 B.n77 B.n76 163.367
R1121 B.n1048 B.n77 163.367
R1122 B.n1048 B.n82 163.367
R1123 B.n83 B.n82 163.367
R1124 B.n84 B.n83 163.367
R1125 B.n1053 B.n84 163.367
R1126 B.n1053 B.n89 163.367
R1127 B.n90 B.n89 163.367
R1128 B.n91 B.n90 163.367
R1129 B.n1058 B.n91 163.367
R1130 B.n1058 B.n96 163.367
R1131 B.n97 B.n96 163.367
R1132 B.n98 B.n97 163.367
R1133 B.n1063 B.n98 163.367
R1134 B.n1063 B.n103 163.367
R1135 B.n104 B.n103 163.367
R1136 B.n105 B.n104 163.367
R1137 B.n1068 B.n105 163.367
R1138 B.n1068 B.n110 163.367
R1139 B.n175 B.n174 163.367
R1140 B.n179 B.n178 163.367
R1141 B.n183 B.n182 163.367
R1142 B.n187 B.n186 163.367
R1143 B.n191 B.n190 163.367
R1144 B.n195 B.n194 163.367
R1145 B.n199 B.n198 163.367
R1146 B.n203 B.n202 163.367
R1147 B.n207 B.n206 163.367
R1148 B.n211 B.n210 163.367
R1149 B.n215 B.n214 163.367
R1150 B.n219 B.n218 163.367
R1151 B.n223 B.n222 163.367
R1152 B.n227 B.n226 163.367
R1153 B.n231 B.n230 163.367
R1154 B.n235 B.n234 163.367
R1155 B.n239 B.n238 163.367
R1156 B.n243 B.n242 163.367
R1157 B.n247 B.n246 163.367
R1158 B.n251 B.n250 163.367
R1159 B.n255 B.n254 163.367
R1160 B.n259 B.n258 163.367
R1161 B.n263 B.n262 163.367
R1162 B.n267 B.n266 163.367
R1163 B.n271 B.n270 163.367
R1164 B.n275 B.n274 163.367
R1165 B.n280 B.n279 163.367
R1166 B.n284 B.n283 163.367
R1167 B.n288 B.n287 163.367
R1168 B.n292 B.n291 163.367
R1169 B.n296 B.n295 163.367
R1170 B.n301 B.n300 163.367
R1171 B.n305 B.n304 163.367
R1172 B.n309 B.n308 163.367
R1173 B.n313 B.n312 163.367
R1174 B.n317 B.n316 163.367
R1175 B.n321 B.n320 163.367
R1176 B.n325 B.n324 163.367
R1177 B.n329 B.n328 163.367
R1178 B.n333 B.n332 163.367
R1179 B.n337 B.n336 163.367
R1180 B.n341 B.n340 163.367
R1181 B.n345 B.n344 163.367
R1182 B.n349 B.n348 163.367
R1183 B.n353 B.n352 163.367
R1184 B.n357 B.n356 163.367
R1185 B.n361 B.n360 163.367
R1186 B.n365 B.n364 163.367
R1187 B.n369 B.n368 163.367
R1188 B.n373 B.n372 163.367
R1189 B.n377 B.n376 163.367
R1190 B.n381 B.n380 163.367
R1191 B.n385 B.n384 163.367
R1192 B.n389 B.n388 163.367
R1193 B.n393 B.n392 163.367
R1194 B.n397 B.n396 163.367
R1195 B.n399 B.n168 163.367
R1196 B.n548 B.t20 128.873
R1197 B.n169 B.t15 128.873
R1198 B.n554 B.t23 128.851
R1199 B.n171 B.t12 128.851
R1200 B.n583 B.n518 71.676
R1201 B.n589 B.n588 71.676
R1202 B.n592 B.n591 71.676
R1203 B.n597 B.n596 71.676
R1204 B.n600 B.n599 71.676
R1205 B.n605 B.n604 71.676
R1206 B.n608 B.n607 71.676
R1207 B.n613 B.n612 71.676
R1208 B.n616 B.n615 71.676
R1209 B.n621 B.n620 71.676
R1210 B.n624 B.n623 71.676
R1211 B.n629 B.n628 71.676
R1212 B.n632 B.n631 71.676
R1213 B.n637 B.n636 71.676
R1214 B.n640 B.n639 71.676
R1215 B.n645 B.n644 71.676
R1216 B.n648 B.n647 71.676
R1217 B.n653 B.n652 71.676
R1218 B.n656 B.n655 71.676
R1219 B.n661 B.n660 71.676
R1220 B.n664 B.n663 71.676
R1221 B.n669 B.n668 71.676
R1222 B.n672 B.n671 71.676
R1223 B.n677 B.n676 71.676
R1224 B.n680 B.n679 71.676
R1225 B.n685 B.n684 71.676
R1226 B.n688 B.n687 71.676
R1227 B.n693 B.n692 71.676
R1228 B.n696 B.n695 71.676
R1229 B.n701 B.n700 71.676
R1230 B.n704 B.n703 71.676
R1231 B.n710 B.n709 71.676
R1232 B.n713 B.n712 71.676
R1233 B.n718 B.n717 71.676
R1234 B.n721 B.n720 71.676
R1235 B.n726 B.n725 71.676
R1236 B.n729 B.n728 71.676
R1237 B.n734 B.n733 71.676
R1238 B.n737 B.n736 71.676
R1239 B.n742 B.n741 71.676
R1240 B.n745 B.n744 71.676
R1241 B.n750 B.n749 71.676
R1242 B.n753 B.n752 71.676
R1243 B.n758 B.n757 71.676
R1244 B.n761 B.n760 71.676
R1245 B.n766 B.n765 71.676
R1246 B.n769 B.n768 71.676
R1247 B.n774 B.n773 71.676
R1248 B.n777 B.n776 71.676
R1249 B.n782 B.n781 71.676
R1250 B.n785 B.n784 71.676
R1251 B.n790 B.n789 71.676
R1252 B.n793 B.n792 71.676
R1253 B.n798 B.n797 71.676
R1254 B.n801 B.n800 71.676
R1255 B.n806 B.n805 71.676
R1256 B.n809 B.n808 71.676
R1257 B.n111 B.n109 71.676
R1258 B.n175 B.n112 71.676
R1259 B.n179 B.n113 71.676
R1260 B.n183 B.n114 71.676
R1261 B.n187 B.n115 71.676
R1262 B.n191 B.n116 71.676
R1263 B.n195 B.n117 71.676
R1264 B.n199 B.n118 71.676
R1265 B.n203 B.n119 71.676
R1266 B.n207 B.n120 71.676
R1267 B.n211 B.n121 71.676
R1268 B.n215 B.n122 71.676
R1269 B.n219 B.n123 71.676
R1270 B.n223 B.n124 71.676
R1271 B.n227 B.n125 71.676
R1272 B.n231 B.n126 71.676
R1273 B.n235 B.n127 71.676
R1274 B.n239 B.n128 71.676
R1275 B.n243 B.n129 71.676
R1276 B.n247 B.n130 71.676
R1277 B.n251 B.n131 71.676
R1278 B.n255 B.n132 71.676
R1279 B.n259 B.n133 71.676
R1280 B.n263 B.n134 71.676
R1281 B.n267 B.n135 71.676
R1282 B.n271 B.n136 71.676
R1283 B.n275 B.n137 71.676
R1284 B.n280 B.n138 71.676
R1285 B.n284 B.n139 71.676
R1286 B.n288 B.n140 71.676
R1287 B.n292 B.n141 71.676
R1288 B.n296 B.n142 71.676
R1289 B.n301 B.n143 71.676
R1290 B.n305 B.n144 71.676
R1291 B.n309 B.n145 71.676
R1292 B.n313 B.n146 71.676
R1293 B.n317 B.n147 71.676
R1294 B.n321 B.n148 71.676
R1295 B.n325 B.n149 71.676
R1296 B.n329 B.n150 71.676
R1297 B.n333 B.n151 71.676
R1298 B.n337 B.n152 71.676
R1299 B.n341 B.n153 71.676
R1300 B.n345 B.n154 71.676
R1301 B.n349 B.n155 71.676
R1302 B.n353 B.n156 71.676
R1303 B.n357 B.n157 71.676
R1304 B.n361 B.n158 71.676
R1305 B.n365 B.n159 71.676
R1306 B.n369 B.n160 71.676
R1307 B.n373 B.n161 71.676
R1308 B.n377 B.n162 71.676
R1309 B.n381 B.n163 71.676
R1310 B.n385 B.n164 71.676
R1311 B.n389 B.n165 71.676
R1312 B.n393 B.n166 71.676
R1313 B.n397 B.n167 71.676
R1314 B.n1073 B.n168 71.676
R1315 B.n1073 B.n1072 71.676
R1316 B.n399 B.n167 71.676
R1317 B.n396 B.n166 71.676
R1318 B.n392 B.n165 71.676
R1319 B.n388 B.n164 71.676
R1320 B.n384 B.n163 71.676
R1321 B.n380 B.n162 71.676
R1322 B.n376 B.n161 71.676
R1323 B.n372 B.n160 71.676
R1324 B.n368 B.n159 71.676
R1325 B.n364 B.n158 71.676
R1326 B.n360 B.n157 71.676
R1327 B.n356 B.n156 71.676
R1328 B.n352 B.n155 71.676
R1329 B.n348 B.n154 71.676
R1330 B.n344 B.n153 71.676
R1331 B.n340 B.n152 71.676
R1332 B.n336 B.n151 71.676
R1333 B.n332 B.n150 71.676
R1334 B.n328 B.n149 71.676
R1335 B.n324 B.n148 71.676
R1336 B.n320 B.n147 71.676
R1337 B.n316 B.n146 71.676
R1338 B.n312 B.n145 71.676
R1339 B.n308 B.n144 71.676
R1340 B.n304 B.n143 71.676
R1341 B.n300 B.n142 71.676
R1342 B.n295 B.n141 71.676
R1343 B.n291 B.n140 71.676
R1344 B.n287 B.n139 71.676
R1345 B.n283 B.n138 71.676
R1346 B.n279 B.n137 71.676
R1347 B.n274 B.n136 71.676
R1348 B.n270 B.n135 71.676
R1349 B.n266 B.n134 71.676
R1350 B.n262 B.n133 71.676
R1351 B.n258 B.n132 71.676
R1352 B.n254 B.n131 71.676
R1353 B.n250 B.n130 71.676
R1354 B.n246 B.n129 71.676
R1355 B.n242 B.n128 71.676
R1356 B.n238 B.n127 71.676
R1357 B.n234 B.n126 71.676
R1358 B.n230 B.n125 71.676
R1359 B.n226 B.n124 71.676
R1360 B.n222 B.n123 71.676
R1361 B.n218 B.n122 71.676
R1362 B.n214 B.n121 71.676
R1363 B.n210 B.n120 71.676
R1364 B.n206 B.n119 71.676
R1365 B.n202 B.n118 71.676
R1366 B.n198 B.n117 71.676
R1367 B.n194 B.n116 71.676
R1368 B.n190 B.n115 71.676
R1369 B.n186 B.n114 71.676
R1370 B.n182 B.n113 71.676
R1371 B.n178 B.n112 71.676
R1372 B.n174 B.n111 71.676
R1373 B.n584 B.n583 71.676
R1374 B.n590 B.n589 71.676
R1375 B.n591 B.n580 71.676
R1376 B.n598 B.n597 71.676
R1377 B.n599 B.n578 71.676
R1378 B.n606 B.n605 71.676
R1379 B.n607 B.n576 71.676
R1380 B.n614 B.n613 71.676
R1381 B.n615 B.n574 71.676
R1382 B.n622 B.n621 71.676
R1383 B.n623 B.n572 71.676
R1384 B.n630 B.n629 71.676
R1385 B.n631 B.n570 71.676
R1386 B.n638 B.n637 71.676
R1387 B.n639 B.n568 71.676
R1388 B.n646 B.n645 71.676
R1389 B.n647 B.n566 71.676
R1390 B.n654 B.n653 71.676
R1391 B.n655 B.n564 71.676
R1392 B.n662 B.n661 71.676
R1393 B.n663 B.n562 71.676
R1394 B.n670 B.n669 71.676
R1395 B.n671 B.n560 71.676
R1396 B.n678 B.n677 71.676
R1397 B.n679 B.n558 71.676
R1398 B.n686 B.n685 71.676
R1399 B.n687 B.n553 71.676
R1400 B.n694 B.n693 71.676
R1401 B.n695 B.n551 71.676
R1402 B.n702 B.n701 71.676
R1403 B.n703 B.n547 71.676
R1404 B.n711 B.n710 71.676
R1405 B.n712 B.n545 71.676
R1406 B.n719 B.n718 71.676
R1407 B.n720 B.n543 71.676
R1408 B.n727 B.n726 71.676
R1409 B.n728 B.n541 71.676
R1410 B.n735 B.n734 71.676
R1411 B.n736 B.n539 71.676
R1412 B.n743 B.n742 71.676
R1413 B.n744 B.n537 71.676
R1414 B.n751 B.n750 71.676
R1415 B.n752 B.n535 71.676
R1416 B.n759 B.n758 71.676
R1417 B.n760 B.n533 71.676
R1418 B.n767 B.n766 71.676
R1419 B.n768 B.n531 71.676
R1420 B.n775 B.n774 71.676
R1421 B.n776 B.n529 71.676
R1422 B.n783 B.n782 71.676
R1423 B.n784 B.n527 71.676
R1424 B.n791 B.n790 71.676
R1425 B.n792 B.n525 71.676
R1426 B.n799 B.n798 71.676
R1427 B.n800 B.n523 71.676
R1428 B.n807 B.n806 71.676
R1429 B.n810 B.n809 71.676
R1430 B.n549 B.t19 71.6605
R1431 B.n170 B.t16 71.6605
R1432 B.n555 B.t22 71.6398
R1433 B.n172 B.t13 71.6398
R1434 B.n815 B.n519 70.2631
R1435 B.n1075 B.n1074 70.2631
R1436 B.n707 B.n549 59.5399
R1437 B.n556 B.n555 59.5399
R1438 B.n277 B.n172 59.5399
R1439 B.n298 B.n170 59.5399
R1440 B.n549 B.n548 57.2126
R1441 B.n555 B.n554 57.2126
R1442 B.n172 B.n171 57.2126
R1443 B.n170 B.n169 57.2126
R1444 B.n815 B.n515 35.392
R1445 B.n821 B.n515 35.392
R1446 B.n821 B.n511 35.392
R1447 B.n827 B.n511 35.392
R1448 B.n827 B.n506 35.392
R1449 B.n833 B.n506 35.392
R1450 B.n833 B.n507 35.392
R1451 B.n839 B.n499 35.392
R1452 B.n845 B.n499 35.392
R1453 B.n845 B.n495 35.392
R1454 B.n851 B.n495 35.392
R1455 B.n851 B.n491 35.392
R1456 B.n857 B.n491 35.392
R1457 B.n857 B.n487 35.392
R1458 B.n863 B.n487 35.392
R1459 B.n863 B.n482 35.392
R1460 B.n869 B.n482 35.392
R1461 B.n869 B.n483 35.392
R1462 B.n875 B.n475 35.392
R1463 B.n881 B.n475 35.392
R1464 B.n881 B.n471 35.392
R1465 B.n887 B.n471 35.392
R1466 B.n887 B.n467 35.392
R1467 B.n893 B.n467 35.392
R1468 B.n893 B.n463 35.392
R1469 B.n899 B.n463 35.392
R1470 B.n905 B.n459 35.392
R1471 B.n905 B.n455 35.392
R1472 B.n911 B.n455 35.392
R1473 B.n911 B.n451 35.392
R1474 B.n917 B.n451 35.392
R1475 B.n917 B.n447 35.392
R1476 B.n923 B.n447 35.392
R1477 B.n929 B.n443 35.392
R1478 B.n929 B.n439 35.392
R1479 B.n935 B.n439 35.392
R1480 B.n935 B.n435 35.392
R1481 B.n941 B.n435 35.392
R1482 B.n941 B.n431 35.392
R1483 B.n948 B.n431 35.392
R1484 B.n948 B.n947 35.392
R1485 B.n954 B.n424 35.392
R1486 B.n960 B.n424 35.392
R1487 B.n960 B.n420 35.392
R1488 B.n966 B.n420 35.392
R1489 B.n966 B.n416 35.392
R1490 B.n972 B.n416 35.392
R1491 B.n972 B.n412 35.392
R1492 B.n978 B.n412 35.392
R1493 B.n985 B.n408 35.392
R1494 B.n985 B.n404 35.392
R1495 B.n991 B.n404 35.392
R1496 B.n991 B.n4 35.392
R1497 B.n1195 B.n4 35.392
R1498 B.n1195 B.n1194 35.392
R1499 B.n1194 B.n1193 35.392
R1500 B.n1193 B.n8 35.392
R1501 B.n1187 B.n8 35.392
R1502 B.n1187 B.n1186 35.392
R1503 B.n1185 B.n15 35.392
R1504 B.n1179 B.n15 35.392
R1505 B.n1179 B.n1178 35.392
R1506 B.n1178 B.n1177 35.392
R1507 B.n1177 B.n22 35.392
R1508 B.n1171 B.n22 35.392
R1509 B.n1171 B.n1170 35.392
R1510 B.n1170 B.n1169 35.392
R1511 B.n1163 B.n32 35.392
R1512 B.n1163 B.n1162 35.392
R1513 B.n1162 B.n1161 35.392
R1514 B.n1161 B.n36 35.392
R1515 B.n1155 B.n36 35.392
R1516 B.n1155 B.n1154 35.392
R1517 B.n1154 B.n1153 35.392
R1518 B.n1153 B.n43 35.392
R1519 B.n1147 B.n1146 35.392
R1520 B.n1146 B.n1145 35.392
R1521 B.n1145 B.n50 35.392
R1522 B.n1139 B.n50 35.392
R1523 B.n1139 B.n1138 35.392
R1524 B.n1138 B.n1137 35.392
R1525 B.n1137 B.n57 35.392
R1526 B.n1131 B.n1130 35.392
R1527 B.n1130 B.n1129 35.392
R1528 B.n1129 B.n64 35.392
R1529 B.n1123 B.n64 35.392
R1530 B.n1123 B.n1122 35.392
R1531 B.n1122 B.n1121 35.392
R1532 B.n1121 B.n71 35.392
R1533 B.n1115 B.n71 35.392
R1534 B.n1114 B.n1113 35.392
R1535 B.n1113 B.n78 35.392
R1536 B.n1107 B.n78 35.392
R1537 B.n1107 B.n1106 35.392
R1538 B.n1106 B.n1105 35.392
R1539 B.n1105 B.n85 35.392
R1540 B.n1099 B.n85 35.392
R1541 B.n1099 B.n1098 35.392
R1542 B.n1098 B.n1097 35.392
R1543 B.n1097 B.n92 35.392
R1544 B.n1091 B.n92 35.392
R1545 B.n1090 B.n1089 35.392
R1546 B.n1089 B.n99 35.392
R1547 B.n1083 B.n99 35.392
R1548 B.n1083 B.n1082 35.392
R1549 B.n1082 B.n1081 35.392
R1550 B.n1081 B.n106 35.392
R1551 B.n1075 B.n106 35.392
R1552 B.t3 B.n459 34.3511
R1553 B.t9 B.n57 34.3511
R1554 B.t2 B.n408 33.3102
R1555 B.n1186 B.t8 33.3102
R1556 B.n1077 B.n108 31.6883
R1557 B.n1071 B.n1070 31.6883
R1558 B.n813 B.n812 31.6883
R1559 B.n817 B.n517 31.6883
R1560 B.n923 B.t5 24.9828
R1561 B.n1147 B.t1 24.9828
R1562 B.n875 B.t7 22.9009
R1563 B.n1115 B.t4 22.9009
R1564 B.n954 B.t6 21.86
R1565 B.n1169 B.t0 21.86
R1566 B.n839 B.t18 18.7372
R1567 B.n1091 B.t11 18.7372
R1568 B B.n1197 18.0485
R1569 B.n507 B.t18 16.6553
R1570 B.t11 B.n1090 16.6553
R1571 B.n947 B.t6 13.5326
R1572 B.n32 B.t0 13.5326
R1573 B.n483 B.t7 12.4916
R1574 B.t4 B.n1114 12.4916
R1575 B.n173 B.n108 10.6151
R1576 B.n176 B.n173 10.6151
R1577 B.n177 B.n176 10.6151
R1578 B.n180 B.n177 10.6151
R1579 B.n181 B.n180 10.6151
R1580 B.n184 B.n181 10.6151
R1581 B.n185 B.n184 10.6151
R1582 B.n188 B.n185 10.6151
R1583 B.n189 B.n188 10.6151
R1584 B.n192 B.n189 10.6151
R1585 B.n193 B.n192 10.6151
R1586 B.n196 B.n193 10.6151
R1587 B.n197 B.n196 10.6151
R1588 B.n200 B.n197 10.6151
R1589 B.n201 B.n200 10.6151
R1590 B.n204 B.n201 10.6151
R1591 B.n205 B.n204 10.6151
R1592 B.n208 B.n205 10.6151
R1593 B.n209 B.n208 10.6151
R1594 B.n212 B.n209 10.6151
R1595 B.n213 B.n212 10.6151
R1596 B.n216 B.n213 10.6151
R1597 B.n217 B.n216 10.6151
R1598 B.n220 B.n217 10.6151
R1599 B.n221 B.n220 10.6151
R1600 B.n224 B.n221 10.6151
R1601 B.n225 B.n224 10.6151
R1602 B.n228 B.n225 10.6151
R1603 B.n229 B.n228 10.6151
R1604 B.n232 B.n229 10.6151
R1605 B.n233 B.n232 10.6151
R1606 B.n236 B.n233 10.6151
R1607 B.n237 B.n236 10.6151
R1608 B.n240 B.n237 10.6151
R1609 B.n241 B.n240 10.6151
R1610 B.n244 B.n241 10.6151
R1611 B.n245 B.n244 10.6151
R1612 B.n248 B.n245 10.6151
R1613 B.n249 B.n248 10.6151
R1614 B.n252 B.n249 10.6151
R1615 B.n253 B.n252 10.6151
R1616 B.n256 B.n253 10.6151
R1617 B.n257 B.n256 10.6151
R1618 B.n260 B.n257 10.6151
R1619 B.n261 B.n260 10.6151
R1620 B.n264 B.n261 10.6151
R1621 B.n265 B.n264 10.6151
R1622 B.n268 B.n265 10.6151
R1623 B.n269 B.n268 10.6151
R1624 B.n272 B.n269 10.6151
R1625 B.n273 B.n272 10.6151
R1626 B.n276 B.n273 10.6151
R1627 B.n281 B.n278 10.6151
R1628 B.n282 B.n281 10.6151
R1629 B.n285 B.n282 10.6151
R1630 B.n286 B.n285 10.6151
R1631 B.n289 B.n286 10.6151
R1632 B.n290 B.n289 10.6151
R1633 B.n293 B.n290 10.6151
R1634 B.n294 B.n293 10.6151
R1635 B.n297 B.n294 10.6151
R1636 B.n302 B.n299 10.6151
R1637 B.n303 B.n302 10.6151
R1638 B.n306 B.n303 10.6151
R1639 B.n307 B.n306 10.6151
R1640 B.n310 B.n307 10.6151
R1641 B.n311 B.n310 10.6151
R1642 B.n314 B.n311 10.6151
R1643 B.n315 B.n314 10.6151
R1644 B.n318 B.n315 10.6151
R1645 B.n319 B.n318 10.6151
R1646 B.n322 B.n319 10.6151
R1647 B.n323 B.n322 10.6151
R1648 B.n326 B.n323 10.6151
R1649 B.n327 B.n326 10.6151
R1650 B.n330 B.n327 10.6151
R1651 B.n331 B.n330 10.6151
R1652 B.n334 B.n331 10.6151
R1653 B.n335 B.n334 10.6151
R1654 B.n338 B.n335 10.6151
R1655 B.n339 B.n338 10.6151
R1656 B.n342 B.n339 10.6151
R1657 B.n343 B.n342 10.6151
R1658 B.n346 B.n343 10.6151
R1659 B.n347 B.n346 10.6151
R1660 B.n350 B.n347 10.6151
R1661 B.n351 B.n350 10.6151
R1662 B.n354 B.n351 10.6151
R1663 B.n355 B.n354 10.6151
R1664 B.n358 B.n355 10.6151
R1665 B.n359 B.n358 10.6151
R1666 B.n362 B.n359 10.6151
R1667 B.n363 B.n362 10.6151
R1668 B.n366 B.n363 10.6151
R1669 B.n367 B.n366 10.6151
R1670 B.n370 B.n367 10.6151
R1671 B.n371 B.n370 10.6151
R1672 B.n374 B.n371 10.6151
R1673 B.n375 B.n374 10.6151
R1674 B.n378 B.n375 10.6151
R1675 B.n379 B.n378 10.6151
R1676 B.n382 B.n379 10.6151
R1677 B.n383 B.n382 10.6151
R1678 B.n386 B.n383 10.6151
R1679 B.n387 B.n386 10.6151
R1680 B.n390 B.n387 10.6151
R1681 B.n391 B.n390 10.6151
R1682 B.n394 B.n391 10.6151
R1683 B.n395 B.n394 10.6151
R1684 B.n398 B.n395 10.6151
R1685 B.n400 B.n398 10.6151
R1686 B.n401 B.n400 10.6151
R1687 B.n1071 B.n401 10.6151
R1688 B.n813 B.n513 10.6151
R1689 B.n823 B.n513 10.6151
R1690 B.n824 B.n823 10.6151
R1691 B.n825 B.n824 10.6151
R1692 B.n825 B.n504 10.6151
R1693 B.n835 B.n504 10.6151
R1694 B.n836 B.n835 10.6151
R1695 B.n837 B.n836 10.6151
R1696 B.n837 B.n497 10.6151
R1697 B.n847 B.n497 10.6151
R1698 B.n848 B.n847 10.6151
R1699 B.n849 B.n848 10.6151
R1700 B.n849 B.n489 10.6151
R1701 B.n859 B.n489 10.6151
R1702 B.n860 B.n859 10.6151
R1703 B.n861 B.n860 10.6151
R1704 B.n861 B.n480 10.6151
R1705 B.n871 B.n480 10.6151
R1706 B.n872 B.n871 10.6151
R1707 B.n873 B.n872 10.6151
R1708 B.n873 B.n473 10.6151
R1709 B.n883 B.n473 10.6151
R1710 B.n884 B.n883 10.6151
R1711 B.n885 B.n884 10.6151
R1712 B.n885 B.n465 10.6151
R1713 B.n895 B.n465 10.6151
R1714 B.n896 B.n895 10.6151
R1715 B.n897 B.n896 10.6151
R1716 B.n897 B.n457 10.6151
R1717 B.n907 B.n457 10.6151
R1718 B.n908 B.n907 10.6151
R1719 B.n909 B.n908 10.6151
R1720 B.n909 B.n449 10.6151
R1721 B.n919 B.n449 10.6151
R1722 B.n920 B.n919 10.6151
R1723 B.n921 B.n920 10.6151
R1724 B.n921 B.n441 10.6151
R1725 B.n931 B.n441 10.6151
R1726 B.n932 B.n931 10.6151
R1727 B.n933 B.n932 10.6151
R1728 B.n933 B.n433 10.6151
R1729 B.n943 B.n433 10.6151
R1730 B.n944 B.n943 10.6151
R1731 B.n945 B.n944 10.6151
R1732 B.n945 B.n426 10.6151
R1733 B.n956 B.n426 10.6151
R1734 B.n957 B.n956 10.6151
R1735 B.n958 B.n957 10.6151
R1736 B.n958 B.n418 10.6151
R1737 B.n968 B.n418 10.6151
R1738 B.n969 B.n968 10.6151
R1739 B.n970 B.n969 10.6151
R1740 B.n970 B.n410 10.6151
R1741 B.n980 B.n410 10.6151
R1742 B.n981 B.n980 10.6151
R1743 B.n983 B.n981 10.6151
R1744 B.n983 B.n982 10.6151
R1745 B.n982 B.n402 10.6151
R1746 B.n994 B.n402 10.6151
R1747 B.n995 B.n994 10.6151
R1748 B.n996 B.n995 10.6151
R1749 B.n997 B.n996 10.6151
R1750 B.n999 B.n997 10.6151
R1751 B.n1000 B.n999 10.6151
R1752 B.n1001 B.n1000 10.6151
R1753 B.n1002 B.n1001 10.6151
R1754 B.n1004 B.n1002 10.6151
R1755 B.n1005 B.n1004 10.6151
R1756 B.n1006 B.n1005 10.6151
R1757 B.n1007 B.n1006 10.6151
R1758 B.n1009 B.n1007 10.6151
R1759 B.n1010 B.n1009 10.6151
R1760 B.n1011 B.n1010 10.6151
R1761 B.n1012 B.n1011 10.6151
R1762 B.n1014 B.n1012 10.6151
R1763 B.n1015 B.n1014 10.6151
R1764 B.n1016 B.n1015 10.6151
R1765 B.n1017 B.n1016 10.6151
R1766 B.n1019 B.n1017 10.6151
R1767 B.n1020 B.n1019 10.6151
R1768 B.n1021 B.n1020 10.6151
R1769 B.n1022 B.n1021 10.6151
R1770 B.n1024 B.n1022 10.6151
R1771 B.n1025 B.n1024 10.6151
R1772 B.n1026 B.n1025 10.6151
R1773 B.n1027 B.n1026 10.6151
R1774 B.n1029 B.n1027 10.6151
R1775 B.n1030 B.n1029 10.6151
R1776 B.n1031 B.n1030 10.6151
R1777 B.n1032 B.n1031 10.6151
R1778 B.n1034 B.n1032 10.6151
R1779 B.n1035 B.n1034 10.6151
R1780 B.n1036 B.n1035 10.6151
R1781 B.n1037 B.n1036 10.6151
R1782 B.n1039 B.n1037 10.6151
R1783 B.n1040 B.n1039 10.6151
R1784 B.n1041 B.n1040 10.6151
R1785 B.n1042 B.n1041 10.6151
R1786 B.n1044 B.n1042 10.6151
R1787 B.n1045 B.n1044 10.6151
R1788 B.n1046 B.n1045 10.6151
R1789 B.n1047 B.n1046 10.6151
R1790 B.n1049 B.n1047 10.6151
R1791 B.n1050 B.n1049 10.6151
R1792 B.n1051 B.n1050 10.6151
R1793 B.n1052 B.n1051 10.6151
R1794 B.n1054 B.n1052 10.6151
R1795 B.n1055 B.n1054 10.6151
R1796 B.n1056 B.n1055 10.6151
R1797 B.n1057 B.n1056 10.6151
R1798 B.n1059 B.n1057 10.6151
R1799 B.n1060 B.n1059 10.6151
R1800 B.n1061 B.n1060 10.6151
R1801 B.n1062 B.n1061 10.6151
R1802 B.n1064 B.n1062 10.6151
R1803 B.n1065 B.n1064 10.6151
R1804 B.n1066 B.n1065 10.6151
R1805 B.n1067 B.n1066 10.6151
R1806 B.n1069 B.n1067 10.6151
R1807 B.n1070 B.n1069 10.6151
R1808 B.n585 B.n517 10.6151
R1809 B.n586 B.n585 10.6151
R1810 B.n587 B.n586 10.6151
R1811 B.n587 B.n581 10.6151
R1812 B.n593 B.n581 10.6151
R1813 B.n594 B.n593 10.6151
R1814 B.n595 B.n594 10.6151
R1815 B.n595 B.n579 10.6151
R1816 B.n601 B.n579 10.6151
R1817 B.n602 B.n601 10.6151
R1818 B.n603 B.n602 10.6151
R1819 B.n603 B.n577 10.6151
R1820 B.n609 B.n577 10.6151
R1821 B.n610 B.n609 10.6151
R1822 B.n611 B.n610 10.6151
R1823 B.n611 B.n575 10.6151
R1824 B.n617 B.n575 10.6151
R1825 B.n618 B.n617 10.6151
R1826 B.n619 B.n618 10.6151
R1827 B.n619 B.n573 10.6151
R1828 B.n625 B.n573 10.6151
R1829 B.n626 B.n625 10.6151
R1830 B.n627 B.n626 10.6151
R1831 B.n627 B.n571 10.6151
R1832 B.n633 B.n571 10.6151
R1833 B.n634 B.n633 10.6151
R1834 B.n635 B.n634 10.6151
R1835 B.n635 B.n569 10.6151
R1836 B.n641 B.n569 10.6151
R1837 B.n642 B.n641 10.6151
R1838 B.n643 B.n642 10.6151
R1839 B.n643 B.n567 10.6151
R1840 B.n649 B.n567 10.6151
R1841 B.n650 B.n649 10.6151
R1842 B.n651 B.n650 10.6151
R1843 B.n651 B.n565 10.6151
R1844 B.n657 B.n565 10.6151
R1845 B.n658 B.n657 10.6151
R1846 B.n659 B.n658 10.6151
R1847 B.n659 B.n563 10.6151
R1848 B.n665 B.n563 10.6151
R1849 B.n666 B.n665 10.6151
R1850 B.n667 B.n666 10.6151
R1851 B.n667 B.n561 10.6151
R1852 B.n673 B.n561 10.6151
R1853 B.n674 B.n673 10.6151
R1854 B.n675 B.n674 10.6151
R1855 B.n675 B.n559 10.6151
R1856 B.n681 B.n559 10.6151
R1857 B.n682 B.n681 10.6151
R1858 B.n683 B.n682 10.6151
R1859 B.n683 B.n557 10.6151
R1860 B.n690 B.n689 10.6151
R1861 B.n691 B.n690 10.6151
R1862 B.n691 B.n552 10.6151
R1863 B.n697 B.n552 10.6151
R1864 B.n698 B.n697 10.6151
R1865 B.n699 B.n698 10.6151
R1866 B.n699 B.n550 10.6151
R1867 B.n705 B.n550 10.6151
R1868 B.n706 B.n705 10.6151
R1869 B.n708 B.n546 10.6151
R1870 B.n714 B.n546 10.6151
R1871 B.n715 B.n714 10.6151
R1872 B.n716 B.n715 10.6151
R1873 B.n716 B.n544 10.6151
R1874 B.n722 B.n544 10.6151
R1875 B.n723 B.n722 10.6151
R1876 B.n724 B.n723 10.6151
R1877 B.n724 B.n542 10.6151
R1878 B.n730 B.n542 10.6151
R1879 B.n731 B.n730 10.6151
R1880 B.n732 B.n731 10.6151
R1881 B.n732 B.n540 10.6151
R1882 B.n738 B.n540 10.6151
R1883 B.n739 B.n738 10.6151
R1884 B.n740 B.n739 10.6151
R1885 B.n740 B.n538 10.6151
R1886 B.n746 B.n538 10.6151
R1887 B.n747 B.n746 10.6151
R1888 B.n748 B.n747 10.6151
R1889 B.n748 B.n536 10.6151
R1890 B.n754 B.n536 10.6151
R1891 B.n755 B.n754 10.6151
R1892 B.n756 B.n755 10.6151
R1893 B.n756 B.n534 10.6151
R1894 B.n762 B.n534 10.6151
R1895 B.n763 B.n762 10.6151
R1896 B.n764 B.n763 10.6151
R1897 B.n764 B.n532 10.6151
R1898 B.n770 B.n532 10.6151
R1899 B.n771 B.n770 10.6151
R1900 B.n772 B.n771 10.6151
R1901 B.n772 B.n530 10.6151
R1902 B.n778 B.n530 10.6151
R1903 B.n779 B.n778 10.6151
R1904 B.n780 B.n779 10.6151
R1905 B.n780 B.n528 10.6151
R1906 B.n786 B.n528 10.6151
R1907 B.n787 B.n786 10.6151
R1908 B.n788 B.n787 10.6151
R1909 B.n788 B.n526 10.6151
R1910 B.n794 B.n526 10.6151
R1911 B.n795 B.n794 10.6151
R1912 B.n796 B.n795 10.6151
R1913 B.n796 B.n524 10.6151
R1914 B.n802 B.n524 10.6151
R1915 B.n803 B.n802 10.6151
R1916 B.n804 B.n803 10.6151
R1917 B.n804 B.n522 10.6151
R1918 B.n522 B.n521 10.6151
R1919 B.n811 B.n521 10.6151
R1920 B.n812 B.n811 10.6151
R1921 B.n818 B.n817 10.6151
R1922 B.n819 B.n818 10.6151
R1923 B.n819 B.n509 10.6151
R1924 B.n829 B.n509 10.6151
R1925 B.n830 B.n829 10.6151
R1926 B.n831 B.n830 10.6151
R1927 B.n831 B.n501 10.6151
R1928 B.n841 B.n501 10.6151
R1929 B.n842 B.n841 10.6151
R1930 B.n843 B.n842 10.6151
R1931 B.n843 B.n493 10.6151
R1932 B.n853 B.n493 10.6151
R1933 B.n854 B.n853 10.6151
R1934 B.n855 B.n854 10.6151
R1935 B.n855 B.n485 10.6151
R1936 B.n865 B.n485 10.6151
R1937 B.n866 B.n865 10.6151
R1938 B.n867 B.n866 10.6151
R1939 B.n867 B.n477 10.6151
R1940 B.n877 B.n477 10.6151
R1941 B.n878 B.n877 10.6151
R1942 B.n879 B.n878 10.6151
R1943 B.n879 B.n469 10.6151
R1944 B.n889 B.n469 10.6151
R1945 B.n890 B.n889 10.6151
R1946 B.n891 B.n890 10.6151
R1947 B.n891 B.n461 10.6151
R1948 B.n901 B.n461 10.6151
R1949 B.n902 B.n901 10.6151
R1950 B.n903 B.n902 10.6151
R1951 B.n903 B.n453 10.6151
R1952 B.n913 B.n453 10.6151
R1953 B.n914 B.n913 10.6151
R1954 B.n915 B.n914 10.6151
R1955 B.n915 B.n445 10.6151
R1956 B.n925 B.n445 10.6151
R1957 B.n926 B.n925 10.6151
R1958 B.n927 B.n926 10.6151
R1959 B.n927 B.n437 10.6151
R1960 B.n937 B.n437 10.6151
R1961 B.n938 B.n937 10.6151
R1962 B.n939 B.n938 10.6151
R1963 B.n939 B.n429 10.6151
R1964 B.n950 B.n429 10.6151
R1965 B.n951 B.n950 10.6151
R1966 B.n952 B.n951 10.6151
R1967 B.n952 B.n422 10.6151
R1968 B.n962 B.n422 10.6151
R1969 B.n963 B.n962 10.6151
R1970 B.n964 B.n963 10.6151
R1971 B.n964 B.n414 10.6151
R1972 B.n974 B.n414 10.6151
R1973 B.n975 B.n974 10.6151
R1974 B.n976 B.n975 10.6151
R1975 B.n976 B.n406 10.6151
R1976 B.n987 B.n406 10.6151
R1977 B.n988 B.n987 10.6151
R1978 B.n989 B.n988 10.6151
R1979 B.n989 B.n0 10.6151
R1980 B.n1191 B.n1 10.6151
R1981 B.n1191 B.n1190 10.6151
R1982 B.n1190 B.n1189 10.6151
R1983 B.n1189 B.n10 10.6151
R1984 B.n1183 B.n10 10.6151
R1985 B.n1183 B.n1182 10.6151
R1986 B.n1182 B.n1181 10.6151
R1987 B.n1181 B.n17 10.6151
R1988 B.n1175 B.n17 10.6151
R1989 B.n1175 B.n1174 10.6151
R1990 B.n1174 B.n1173 10.6151
R1991 B.n1173 B.n24 10.6151
R1992 B.n1167 B.n24 10.6151
R1993 B.n1167 B.n1166 10.6151
R1994 B.n1166 B.n1165 10.6151
R1995 B.n1165 B.n30 10.6151
R1996 B.n1159 B.n30 10.6151
R1997 B.n1159 B.n1158 10.6151
R1998 B.n1158 B.n1157 10.6151
R1999 B.n1157 B.n38 10.6151
R2000 B.n1151 B.n38 10.6151
R2001 B.n1151 B.n1150 10.6151
R2002 B.n1150 B.n1149 10.6151
R2003 B.n1149 B.n45 10.6151
R2004 B.n1143 B.n45 10.6151
R2005 B.n1143 B.n1142 10.6151
R2006 B.n1142 B.n1141 10.6151
R2007 B.n1141 B.n52 10.6151
R2008 B.n1135 B.n52 10.6151
R2009 B.n1135 B.n1134 10.6151
R2010 B.n1134 B.n1133 10.6151
R2011 B.n1133 B.n59 10.6151
R2012 B.n1127 B.n59 10.6151
R2013 B.n1127 B.n1126 10.6151
R2014 B.n1126 B.n1125 10.6151
R2015 B.n1125 B.n66 10.6151
R2016 B.n1119 B.n66 10.6151
R2017 B.n1119 B.n1118 10.6151
R2018 B.n1118 B.n1117 10.6151
R2019 B.n1117 B.n73 10.6151
R2020 B.n1111 B.n73 10.6151
R2021 B.n1111 B.n1110 10.6151
R2022 B.n1110 B.n1109 10.6151
R2023 B.n1109 B.n80 10.6151
R2024 B.n1103 B.n80 10.6151
R2025 B.n1103 B.n1102 10.6151
R2026 B.n1102 B.n1101 10.6151
R2027 B.n1101 B.n87 10.6151
R2028 B.n1095 B.n87 10.6151
R2029 B.n1095 B.n1094 10.6151
R2030 B.n1094 B.n1093 10.6151
R2031 B.n1093 B.n94 10.6151
R2032 B.n1087 B.n94 10.6151
R2033 B.n1087 B.n1086 10.6151
R2034 B.n1086 B.n1085 10.6151
R2035 B.n1085 B.n101 10.6151
R2036 B.n1079 B.n101 10.6151
R2037 B.n1079 B.n1078 10.6151
R2038 B.n1078 B.n1077 10.6151
R2039 B.t5 B.n443 10.4098
R2040 B.t1 B.n43 10.4098
R2041 B.n277 B.n276 9.36635
R2042 B.n299 B.n298 9.36635
R2043 B.n557 B.n556 9.36635
R2044 B.n708 B.n707 9.36635
R2045 B.n1197 B.n0 2.81026
R2046 B.n1197 B.n1 2.81026
R2047 B.n978 B.t2 2.08235
R2048 B.t8 B.n1185 2.08235
R2049 B.n278 B.n277 1.24928
R2050 B.n298 B.n297 1.24928
R2051 B.n689 B.n556 1.24928
R2052 B.n707 B.n706 1.24928
R2053 B.n899 B.t3 1.04143
R2054 B.n1131 B.t9 1.04143
R2055 VP.n24 VP.t2 178.786
R2056 VP.n25 VP.n22 161.3
R2057 VP.n27 VP.n26 161.3
R2058 VP.n28 VP.n21 161.3
R2059 VP.n30 VP.n29 161.3
R2060 VP.n31 VP.n20 161.3
R2061 VP.n33 VP.n32 161.3
R2062 VP.n35 VP.n19 161.3
R2063 VP.n37 VP.n36 161.3
R2064 VP.n38 VP.n18 161.3
R2065 VP.n40 VP.n39 161.3
R2066 VP.n41 VP.n17 161.3
R2067 VP.n43 VP.n42 161.3
R2068 VP.n45 VP.n44 161.3
R2069 VP.n46 VP.n15 161.3
R2070 VP.n48 VP.n47 161.3
R2071 VP.n49 VP.n14 161.3
R2072 VP.n51 VP.n50 161.3
R2073 VP.n52 VP.n13 161.3
R2074 VP.n94 VP.n0 161.3
R2075 VP.n93 VP.n92 161.3
R2076 VP.n91 VP.n1 161.3
R2077 VP.n90 VP.n89 161.3
R2078 VP.n88 VP.n2 161.3
R2079 VP.n87 VP.n86 161.3
R2080 VP.n85 VP.n84 161.3
R2081 VP.n83 VP.n4 161.3
R2082 VP.n82 VP.n81 161.3
R2083 VP.n80 VP.n5 161.3
R2084 VP.n79 VP.n78 161.3
R2085 VP.n77 VP.n6 161.3
R2086 VP.n75 VP.n74 161.3
R2087 VP.n73 VP.n7 161.3
R2088 VP.n72 VP.n71 161.3
R2089 VP.n70 VP.n8 161.3
R2090 VP.n69 VP.n68 161.3
R2091 VP.n67 VP.n9 161.3
R2092 VP.n66 VP.n65 161.3
R2093 VP.n63 VP.n10 161.3
R2094 VP.n62 VP.n61 161.3
R2095 VP.n60 VP.n11 161.3
R2096 VP.n59 VP.n58 161.3
R2097 VP.n57 VP.n12 161.3
R2098 VP.n56 VP.t6 145.888
R2099 VP.n64 VP.t9 145.888
R2100 VP.n76 VP.t4 145.888
R2101 VP.n3 VP.t8 145.888
R2102 VP.n95 VP.t0 145.888
R2103 VP.n53 VP.t5 145.888
R2104 VP.n16 VP.t3 145.888
R2105 VP.n34 VP.t1 145.888
R2106 VP.n23 VP.t7 145.888
R2107 VP.n56 VP.n55 103.531
R2108 VP.n96 VP.n95 103.531
R2109 VP.n54 VP.n53 103.531
R2110 VP.n24 VP.n23 62.6783
R2111 VP.n62 VP.n11 56.5617
R2112 VP.n71 VP.n70 56.5617
R2113 VP.n82 VP.n5 56.5617
R2114 VP.n89 VP.n1 56.5617
R2115 VP.n47 VP.n14 56.5617
R2116 VP.n40 VP.n18 56.5617
R2117 VP.n29 VP.n28 56.5617
R2118 VP.n55 VP.n54 56.1322
R2119 VP.n58 VP.n57 24.5923
R2120 VP.n58 VP.n11 24.5923
R2121 VP.n63 VP.n62 24.5923
R2122 VP.n65 VP.n63 24.5923
R2123 VP.n69 VP.n9 24.5923
R2124 VP.n70 VP.n69 24.5923
R2125 VP.n71 VP.n7 24.5923
R2126 VP.n75 VP.n7 24.5923
R2127 VP.n78 VP.n77 24.5923
R2128 VP.n78 VP.n5 24.5923
R2129 VP.n83 VP.n82 24.5923
R2130 VP.n84 VP.n83 24.5923
R2131 VP.n88 VP.n87 24.5923
R2132 VP.n89 VP.n88 24.5923
R2133 VP.n93 VP.n1 24.5923
R2134 VP.n94 VP.n93 24.5923
R2135 VP.n51 VP.n14 24.5923
R2136 VP.n52 VP.n51 24.5923
R2137 VP.n41 VP.n40 24.5923
R2138 VP.n42 VP.n41 24.5923
R2139 VP.n46 VP.n45 24.5923
R2140 VP.n47 VP.n46 24.5923
R2141 VP.n29 VP.n20 24.5923
R2142 VP.n33 VP.n20 24.5923
R2143 VP.n36 VP.n35 24.5923
R2144 VP.n36 VP.n18 24.5923
R2145 VP.n27 VP.n22 24.5923
R2146 VP.n28 VP.n27 24.5923
R2147 VP.n65 VP.n64 14.7556
R2148 VP.n87 VP.n3 14.7556
R2149 VP.n45 VP.n16 14.7556
R2150 VP.n76 VP.n75 12.2964
R2151 VP.n77 VP.n76 12.2964
R2152 VP.n34 VP.n33 12.2964
R2153 VP.n35 VP.n34 12.2964
R2154 VP.n64 VP.n9 9.83723
R2155 VP.n84 VP.n3 9.83723
R2156 VP.n42 VP.n16 9.83723
R2157 VP.n23 VP.n22 9.83723
R2158 VP.n57 VP.n56 7.37805
R2159 VP.n95 VP.n94 7.37805
R2160 VP.n53 VP.n52 7.37805
R2161 VP.n25 VP.n24 6.9978
R2162 VP.n54 VP.n13 0.278335
R2163 VP.n55 VP.n12 0.278335
R2164 VP.n96 VP.n0 0.278335
R2165 VP.n26 VP.n25 0.189894
R2166 VP.n26 VP.n21 0.189894
R2167 VP.n30 VP.n21 0.189894
R2168 VP.n31 VP.n30 0.189894
R2169 VP.n32 VP.n31 0.189894
R2170 VP.n32 VP.n19 0.189894
R2171 VP.n37 VP.n19 0.189894
R2172 VP.n38 VP.n37 0.189894
R2173 VP.n39 VP.n38 0.189894
R2174 VP.n39 VP.n17 0.189894
R2175 VP.n43 VP.n17 0.189894
R2176 VP.n44 VP.n43 0.189894
R2177 VP.n44 VP.n15 0.189894
R2178 VP.n48 VP.n15 0.189894
R2179 VP.n49 VP.n48 0.189894
R2180 VP.n50 VP.n49 0.189894
R2181 VP.n50 VP.n13 0.189894
R2182 VP.n59 VP.n12 0.189894
R2183 VP.n60 VP.n59 0.189894
R2184 VP.n61 VP.n60 0.189894
R2185 VP.n61 VP.n10 0.189894
R2186 VP.n66 VP.n10 0.189894
R2187 VP.n67 VP.n66 0.189894
R2188 VP.n68 VP.n67 0.189894
R2189 VP.n68 VP.n8 0.189894
R2190 VP.n72 VP.n8 0.189894
R2191 VP.n73 VP.n72 0.189894
R2192 VP.n74 VP.n73 0.189894
R2193 VP.n74 VP.n6 0.189894
R2194 VP.n79 VP.n6 0.189894
R2195 VP.n80 VP.n79 0.189894
R2196 VP.n81 VP.n80 0.189894
R2197 VP.n81 VP.n4 0.189894
R2198 VP.n85 VP.n4 0.189894
R2199 VP.n86 VP.n85 0.189894
R2200 VP.n86 VP.n2 0.189894
R2201 VP.n90 VP.n2 0.189894
R2202 VP.n91 VP.n90 0.189894
R2203 VP.n92 VP.n91 0.189894
R2204 VP.n92 VP.n0 0.189894
R2205 VP VP.n96 0.153485
R2206 VTAIL.n11 VTAIL.t8 48.093
R2207 VTAIL.n17 VTAIL.t2 48.0929
R2208 VTAIL.n2 VTAIL.t16 48.0929
R2209 VTAIL.n16 VTAIL.t12 48.0929
R2210 VTAIL.n15 VTAIL.n14 46.8447
R2211 VTAIL.n13 VTAIL.n12 46.8447
R2212 VTAIL.n10 VTAIL.n9 46.8447
R2213 VTAIL.n8 VTAIL.n7 46.8447
R2214 VTAIL.n19 VTAIL.n18 46.8444
R2215 VTAIL.n1 VTAIL.n0 46.8444
R2216 VTAIL.n4 VTAIL.n3 46.8444
R2217 VTAIL.n6 VTAIL.n5 46.8444
R2218 VTAIL.n8 VTAIL.n6 31.1255
R2219 VTAIL.n17 VTAIL.n16 28.5824
R2220 VTAIL.n10 VTAIL.n8 2.5436
R2221 VTAIL.n11 VTAIL.n10 2.5436
R2222 VTAIL.n15 VTAIL.n13 2.5436
R2223 VTAIL.n16 VTAIL.n15 2.5436
R2224 VTAIL.n6 VTAIL.n4 2.5436
R2225 VTAIL.n4 VTAIL.n2 2.5436
R2226 VTAIL.n19 VTAIL.n17 2.5436
R2227 VTAIL VTAIL.n1 1.96602
R2228 VTAIL.n13 VTAIL.n11 1.74188
R2229 VTAIL.n2 VTAIL.n1 1.74188
R2230 VTAIL.n18 VTAIL.t1 1.24892
R2231 VTAIL.n18 VTAIL.t5 1.24892
R2232 VTAIL.n0 VTAIL.t4 1.24892
R2233 VTAIL.n0 VTAIL.t0 1.24892
R2234 VTAIL.n3 VTAIL.t11 1.24892
R2235 VTAIL.n3 VTAIL.t10 1.24892
R2236 VTAIL.n5 VTAIL.t17 1.24892
R2237 VTAIL.n5 VTAIL.t15 1.24892
R2238 VTAIL.n14 VTAIL.t14 1.24892
R2239 VTAIL.n14 VTAIL.t19 1.24892
R2240 VTAIL.n12 VTAIL.t13 1.24892
R2241 VTAIL.n12 VTAIL.t18 1.24892
R2242 VTAIL.n9 VTAIL.t3 1.24892
R2243 VTAIL.n9 VTAIL.t7 1.24892
R2244 VTAIL.n7 VTAIL.t9 1.24892
R2245 VTAIL.n7 VTAIL.t6 1.24892
R2246 VTAIL VTAIL.n19 0.578086
R2247 VDD1.n1 VDD1.t7 67.3149
R2248 VDD1.n3 VDD1.t3 67.3148
R2249 VDD1.n5 VDD1.n4 65.3752
R2250 VDD1.n1 VDD1.n0 63.5234
R2251 VDD1.n7 VDD1.n6 63.5233
R2252 VDD1.n3 VDD1.n2 63.5232
R2253 VDD1.n7 VDD1.n5 51.322
R2254 VDD1 VDD1.n7 1.84964
R2255 VDD1.n6 VDD1.t6 1.24892
R2256 VDD1.n6 VDD1.t4 1.24892
R2257 VDD1.n0 VDD1.t2 1.24892
R2258 VDD1.n0 VDD1.t8 1.24892
R2259 VDD1.n4 VDD1.t1 1.24892
R2260 VDD1.n4 VDD1.t9 1.24892
R2261 VDD1.n2 VDD1.t0 1.24892
R2262 VDD1.n2 VDD1.t5 1.24892
R2263 VDD1 VDD1.n1 0.694465
R2264 VDD1.n5 VDD1.n3 0.58093
R2265 VN.n11 VN.t3 178.786
R2266 VN.n53 VN.t6 178.786
R2267 VN.n81 VN.n42 161.3
R2268 VN.n80 VN.n79 161.3
R2269 VN.n78 VN.n43 161.3
R2270 VN.n77 VN.n76 161.3
R2271 VN.n75 VN.n44 161.3
R2272 VN.n74 VN.n73 161.3
R2273 VN.n72 VN.n71 161.3
R2274 VN.n70 VN.n46 161.3
R2275 VN.n69 VN.n68 161.3
R2276 VN.n67 VN.n47 161.3
R2277 VN.n66 VN.n65 161.3
R2278 VN.n64 VN.n48 161.3
R2279 VN.n62 VN.n61 161.3
R2280 VN.n60 VN.n49 161.3
R2281 VN.n59 VN.n58 161.3
R2282 VN.n57 VN.n50 161.3
R2283 VN.n56 VN.n55 161.3
R2284 VN.n54 VN.n51 161.3
R2285 VN.n39 VN.n0 161.3
R2286 VN.n38 VN.n37 161.3
R2287 VN.n36 VN.n1 161.3
R2288 VN.n35 VN.n34 161.3
R2289 VN.n33 VN.n2 161.3
R2290 VN.n32 VN.n31 161.3
R2291 VN.n30 VN.n29 161.3
R2292 VN.n28 VN.n4 161.3
R2293 VN.n27 VN.n26 161.3
R2294 VN.n25 VN.n5 161.3
R2295 VN.n24 VN.n23 161.3
R2296 VN.n22 VN.n6 161.3
R2297 VN.n20 VN.n19 161.3
R2298 VN.n18 VN.n7 161.3
R2299 VN.n17 VN.n16 161.3
R2300 VN.n15 VN.n8 161.3
R2301 VN.n14 VN.n13 161.3
R2302 VN.n12 VN.n9 161.3
R2303 VN.n10 VN.t9 145.888
R2304 VN.n21 VN.t5 145.888
R2305 VN.n3 VN.t2 145.888
R2306 VN.n40 VN.t8 145.888
R2307 VN.n52 VN.t0 145.888
R2308 VN.n63 VN.t7 145.888
R2309 VN.n45 VN.t1 145.888
R2310 VN.n82 VN.t4 145.888
R2311 VN.n41 VN.n40 103.531
R2312 VN.n83 VN.n82 103.531
R2313 VN.n11 VN.n10 62.6783
R2314 VN.n53 VN.n52 62.6783
R2315 VN.n16 VN.n15 56.5617
R2316 VN.n27 VN.n5 56.5617
R2317 VN.n34 VN.n1 56.5617
R2318 VN.n58 VN.n57 56.5617
R2319 VN.n69 VN.n47 56.5617
R2320 VN.n76 VN.n43 56.5617
R2321 VN VN.n83 56.4111
R2322 VN.n14 VN.n9 24.5923
R2323 VN.n15 VN.n14 24.5923
R2324 VN.n16 VN.n7 24.5923
R2325 VN.n20 VN.n7 24.5923
R2326 VN.n23 VN.n22 24.5923
R2327 VN.n23 VN.n5 24.5923
R2328 VN.n28 VN.n27 24.5923
R2329 VN.n29 VN.n28 24.5923
R2330 VN.n33 VN.n32 24.5923
R2331 VN.n34 VN.n33 24.5923
R2332 VN.n38 VN.n1 24.5923
R2333 VN.n39 VN.n38 24.5923
R2334 VN.n57 VN.n56 24.5923
R2335 VN.n56 VN.n51 24.5923
R2336 VN.n65 VN.n47 24.5923
R2337 VN.n65 VN.n64 24.5923
R2338 VN.n62 VN.n49 24.5923
R2339 VN.n58 VN.n49 24.5923
R2340 VN.n76 VN.n75 24.5923
R2341 VN.n75 VN.n74 24.5923
R2342 VN.n71 VN.n70 24.5923
R2343 VN.n70 VN.n69 24.5923
R2344 VN.n81 VN.n80 24.5923
R2345 VN.n80 VN.n43 24.5923
R2346 VN.n32 VN.n3 14.7556
R2347 VN.n74 VN.n45 14.7556
R2348 VN.n21 VN.n20 12.2964
R2349 VN.n22 VN.n21 12.2964
R2350 VN.n64 VN.n63 12.2964
R2351 VN.n63 VN.n62 12.2964
R2352 VN.n10 VN.n9 9.83723
R2353 VN.n29 VN.n3 9.83723
R2354 VN.n52 VN.n51 9.83723
R2355 VN.n71 VN.n45 9.83723
R2356 VN.n40 VN.n39 7.37805
R2357 VN.n82 VN.n81 7.37805
R2358 VN.n54 VN.n53 6.9978
R2359 VN.n12 VN.n11 6.9978
R2360 VN.n83 VN.n42 0.278335
R2361 VN.n41 VN.n0 0.278335
R2362 VN.n79 VN.n42 0.189894
R2363 VN.n79 VN.n78 0.189894
R2364 VN.n78 VN.n77 0.189894
R2365 VN.n77 VN.n44 0.189894
R2366 VN.n73 VN.n44 0.189894
R2367 VN.n73 VN.n72 0.189894
R2368 VN.n72 VN.n46 0.189894
R2369 VN.n68 VN.n46 0.189894
R2370 VN.n68 VN.n67 0.189894
R2371 VN.n67 VN.n66 0.189894
R2372 VN.n66 VN.n48 0.189894
R2373 VN.n61 VN.n48 0.189894
R2374 VN.n61 VN.n60 0.189894
R2375 VN.n60 VN.n59 0.189894
R2376 VN.n59 VN.n50 0.189894
R2377 VN.n55 VN.n50 0.189894
R2378 VN.n55 VN.n54 0.189894
R2379 VN.n13 VN.n12 0.189894
R2380 VN.n13 VN.n8 0.189894
R2381 VN.n17 VN.n8 0.189894
R2382 VN.n18 VN.n17 0.189894
R2383 VN.n19 VN.n18 0.189894
R2384 VN.n19 VN.n6 0.189894
R2385 VN.n24 VN.n6 0.189894
R2386 VN.n25 VN.n24 0.189894
R2387 VN.n26 VN.n25 0.189894
R2388 VN.n26 VN.n4 0.189894
R2389 VN.n30 VN.n4 0.189894
R2390 VN.n31 VN.n30 0.189894
R2391 VN.n31 VN.n2 0.189894
R2392 VN.n35 VN.n2 0.189894
R2393 VN.n36 VN.n35 0.189894
R2394 VN.n37 VN.n36 0.189894
R2395 VN.n37 VN.n0 0.189894
R2396 VN VN.n41 0.153485
R2397 VDD2.n1 VDD2.t6 67.3148
R2398 VDD2.n3 VDD2.n2 65.3752
R2399 VDD2 VDD2.n7 65.3724
R2400 VDD2.n4 VDD2.t5 64.7718
R2401 VDD2.n6 VDD2.n5 63.5234
R2402 VDD2.n1 VDD2.n0 63.5232
R2403 VDD2.n4 VDD2.n3 49.4674
R2404 VDD2.n6 VDD2.n4 2.5436
R2405 VDD2.n7 VDD2.t9 1.24892
R2406 VDD2.n7 VDD2.t3 1.24892
R2407 VDD2.n5 VDD2.t8 1.24892
R2408 VDD2.n5 VDD2.t2 1.24892
R2409 VDD2.n2 VDD2.t7 1.24892
R2410 VDD2.n2 VDD2.t1 1.24892
R2411 VDD2.n0 VDD2.t0 1.24892
R2412 VDD2.n0 VDD2.t4 1.24892
R2413 VDD2 VDD2.n6 0.694465
R2414 VDD2.n3 VDD2.n1 0.58093
C0 VDD2 VP 0.586928f
C1 VDD1 VDD2 2.18898f
C2 VDD1 VP 14.379801f
C3 VDD2 VN 13.9512f
C4 VP VN 9.13617f
C5 VDD2 VTAIL 12.2207f
C6 VDD1 VN 0.153897f
C7 VP VTAIL 14.442599f
C8 VDD1 VTAIL 12.170401f
C9 VN VTAIL 14.4283f
C10 VDD2 B 7.916133f
C11 VDD1 B 7.891484f
C12 VTAIL B 9.763324f
C13 VN B 18.539072f
C14 VP B 17.012846f
C15 VDD2.t6 B 3.46614f
C16 VDD2.t0 B 0.297558f
C17 VDD2.t4 B 0.297558f
C18 VDD2.n0 B 2.69923f
C19 VDD2.n1 B 0.87361f
C20 VDD2.t7 B 0.297558f
C21 VDD2.t1 B 0.297558f
C22 VDD2.n2 B 2.71449f
C23 VDD2.n3 B 2.99515f
C24 VDD2.t5 B 3.44883f
C25 VDD2.n4 B 3.25087f
C26 VDD2.t8 B 0.297558f
C27 VDD2.t2 B 0.297558f
C28 VDD2.n5 B 2.69924f
C29 VDD2.n6 B 0.440127f
C30 VDD2.t9 B 0.297558f
C31 VDD2.t3 B 0.297558f
C32 VDD2.n7 B 2.71445f
C33 VN.n0 B 0.027262f
C34 VN.t8 B 2.35754f
C35 VN.n1 B 0.034352f
C36 VN.n2 B 0.020679f
C37 VN.t2 B 2.35754f
C38 VN.n3 B 0.821647f
C39 VN.n4 B 0.020679f
C40 VN.n5 B 0.02863f
C41 VN.n6 B 0.020679f
C42 VN.t5 B 2.35754f
C43 VN.n7 B 0.038348f
C44 VN.n8 B 0.020679f
C45 VN.n9 B 0.026989f
C46 VN.t3 B 2.53212f
C47 VN.t9 B 2.35754f
C48 VN.n10 B 0.879272f
C49 VN.n11 B 0.860316f
C50 VN.n12 B 0.200201f
C51 VN.n13 B 0.020679f
C52 VN.n14 B 0.038348f
C53 VN.n15 B 0.031491f
C54 VN.n16 B 0.02863f
C55 VN.n17 B 0.020679f
C56 VN.n18 B 0.020679f
C57 VN.n19 B 0.020679f
C58 VN.n20 B 0.028882f
C59 VN.n21 B 0.821647f
C60 VN.n22 B 0.028882f
C61 VN.n23 B 0.038348f
C62 VN.n24 B 0.020679f
C63 VN.n25 B 0.020679f
C64 VN.n26 B 0.020679f
C65 VN.n27 B 0.031491f
C66 VN.n28 B 0.038348f
C67 VN.n29 B 0.026989f
C68 VN.n30 B 0.020679f
C69 VN.n31 B 0.020679f
C70 VN.n32 B 0.030776f
C71 VN.n33 B 0.038348f
C72 VN.n34 B 0.02577f
C73 VN.n35 B 0.020679f
C74 VN.n36 B 0.020679f
C75 VN.n37 B 0.020679f
C76 VN.n38 B 0.038348f
C77 VN.n39 B 0.025096f
C78 VN.n40 B 0.888131f
C79 VN.n41 B 0.035111f
C80 VN.n42 B 0.027262f
C81 VN.t4 B 2.35754f
C82 VN.n43 B 0.034352f
C83 VN.n44 B 0.020679f
C84 VN.t1 B 2.35754f
C85 VN.n45 B 0.821647f
C86 VN.n46 B 0.020679f
C87 VN.n47 B 0.02863f
C88 VN.n48 B 0.020679f
C89 VN.t7 B 2.35754f
C90 VN.n49 B 0.038348f
C91 VN.n50 B 0.020679f
C92 VN.n51 B 0.026989f
C93 VN.t6 B 2.53212f
C94 VN.t0 B 2.35754f
C95 VN.n52 B 0.879272f
C96 VN.n53 B 0.860316f
C97 VN.n54 B 0.200201f
C98 VN.n55 B 0.020679f
C99 VN.n56 B 0.038348f
C100 VN.n57 B 0.031491f
C101 VN.n58 B 0.02863f
C102 VN.n59 B 0.020679f
C103 VN.n60 B 0.020679f
C104 VN.n61 B 0.020679f
C105 VN.n62 B 0.028882f
C106 VN.n63 B 0.821647f
C107 VN.n64 B 0.028882f
C108 VN.n65 B 0.038348f
C109 VN.n66 B 0.020679f
C110 VN.n67 B 0.020679f
C111 VN.n68 B 0.020679f
C112 VN.n69 B 0.031491f
C113 VN.n70 B 0.038348f
C114 VN.n71 B 0.026989f
C115 VN.n72 B 0.020679f
C116 VN.n73 B 0.020679f
C117 VN.n74 B 0.030776f
C118 VN.n75 B 0.038348f
C119 VN.n76 B 0.02577f
C120 VN.n77 B 0.020679f
C121 VN.n78 B 0.020679f
C122 VN.n79 B 0.020679f
C123 VN.n80 B 0.038348f
C124 VN.n81 B 0.025096f
C125 VN.n82 B 0.888131f
C126 VN.n83 B 1.37007f
C127 VDD1.t7 B 3.50415f
C128 VDD1.t2 B 0.30082f
C129 VDD1.t8 B 0.30082f
C130 VDD1.n0 B 2.72883f
C131 VDD1.n1 B 0.890993f
C132 VDD1.t3 B 3.50414f
C133 VDD1.t0 B 0.30082f
C134 VDD1.t5 B 0.30082f
C135 VDD1.n2 B 2.72882f
C136 VDD1.n3 B 0.883188f
C137 VDD1.t1 B 0.30082f
C138 VDD1.t9 B 0.30082f
C139 VDD1.n4 B 2.74425f
C140 VDD1.n5 B 3.1509f
C141 VDD1.t6 B 0.30082f
C142 VDD1.t4 B 0.30082f
C143 VDD1.n6 B 2.72882f
C144 VDD1.n7 B 3.33266f
C145 VTAIL.t4 B 0.30091f
C146 VTAIL.t0 B 0.30091f
C147 VTAIL.n0 B 2.66196f
C148 VTAIL.n1 B 0.516482f
C149 VTAIL.t16 B 3.40002f
C150 VTAIL.n2 B 0.643769f
C151 VTAIL.t11 B 0.30091f
C152 VTAIL.t10 B 0.30091f
C153 VTAIL.n3 B 2.66196f
C154 VTAIL.n4 B 0.623191f
C155 VTAIL.t17 B 0.30091f
C156 VTAIL.t15 B 0.30091f
C157 VTAIL.n5 B 2.66196f
C158 VTAIL.n6 B 2.20382f
C159 VTAIL.t9 B 0.30091f
C160 VTAIL.t6 B 0.30091f
C161 VTAIL.n7 B 2.66197f
C162 VTAIL.n8 B 2.20381f
C163 VTAIL.t3 B 0.30091f
C164 VTAIL.t7 B 0.30091f
C165 VTAIL.n9 B 2.66197f
C166 VTAIL.n10 B 0.623187f
C167 VTAIL.t8 B 3.40005f
C168 VTAIL.n11 B 0.643748f
C169 VTAIL.t13 B 0.30091f
C170 VTAIL.t18 B 0.30091f
C171 VTAIL.n12 B 2.66197f
C172 VTAIL.n13 B 0.561163f
C173 VTAIL.t14 B 0.30091f
C174 VTAIL.t19 B 0.30091f
C175 VTAIL.n14 B 2.66197f
C176 VTAIL.n15 B 0.623187f
C177 VTAIL.t12 B 3.40002f
C178 VTAIL.n16 B 2.08968f
C179 VTAIL.t2 B 3.40002f
C180 VTAIL.n17 B 2.08968f
C181 VTAIL.t1 B 0.30091f
C182 VTAIL.t5 B 0.30091f
C183 VTAIL.n18 B 2.66196f
C184 VTAIL.n19 B 0.471131f
C185 VP.n0 B 0.027574f
C186 VP.t0 B 2.38453f
C187 VP.n1 B 0.034745f
C188 VP.n2 B 0.020916f
C189 VP.t8 B 2.38453f
C190 VP.n3 B 0.831056f
C191 VP.n4 B 0.020916f
C192 VP.n5 B 0.028958f
C193 VP.n6 B 0.020916f
C194 VP.t4 B 2.38453f
C195 VP.n7 B 0.038787f
C196 VP.n8 B 0.020916f
C197 VP.n9 B 0.027298f
C198 VP.n10 B 0.020916f
C199 VP.n11 B 0.034745f
C200 VP.n12 B 0.027574f
C201 VP.t6 B 2.38453f
C202 VP.n13 B 0.027574f
C203 VP.t5 B 2.38453f
C204 VP.n14 B 0.034745f
C205 VP.n15 B 0.020916f
C206 VP.t3 B 2.38453f
C207 VP.n16 B 0.831056f
C208 VP.n17 B 0.020916f
C209 VP.n18 B 0.028958f
C210 VP.n19 B 0.020916f
C211 VP.t1 B 2.38453f
C212 VP.n20 B 0.038787f
C213 VP.n21 B 0.020916f
C214 VP.n22 B 0.027298f
C215 VP.t2 B 2.56111f
C216 VP.t7 B 2.38453f
C217 VP.n23 B 0.88934f
C218 VP.n24 B 0.870167f
C219 VP.n25 B 0.202494f
C220 VP.n26 B 0.020916f
C221 VP.n27 B 0.038787f
C222 VP.n28 B 0.031852f
C223 VP.n29 B 0.028958f
C224 VP.n30 B 0.020916f
C225 VP.n31 B 0.020916f
C226 VP.n32 B 0.020916f
C227 VP.n33 B 0.029213f
C228 VP.n34 B 0.831056f
C229 VP.n35 B 0.029213f
C230 VP.n36 B 0.038787f
C231 VP.n37 B 0.020916f
C232 VP.n38 B 0.020916f
C233 VP.n39 B 0.020916f
C234 VP.n40 B 0.031852f
C235 VP.n41 B 0.038787f
C236 VP.n42 B 0.027298f
C237 VP.n43 B 0.020916f
C238 VP.n44 B 0.020916f
C239 VP.n45 B 0.031128f
C240 VP.n46 B 0.038787f
C241 VP.n47 B 0.026065f
C242 VP.n48 B 0.020916f
C243 VP.n49 B 0.020916f
C244 VP.n50 B 0.020916f
C245 VP.n51 B 0.038787f
C246 VP.n52 B 0.025383f
C247 VP.n53 B 0.8983f
C248 VP.n54 B 1.37471f
C249 VP.n55 B 1.38814f
C250 VP.n56 B 0.8983f
C251 VP.n57 B 0.025383f
C252 VP.n58 B 0.038787f
C253 VP.n59 B 0.020916f
C254 VP.n60 B 0.020916f
C255 VP.n61 B 0.020916f
C256 VP.n62 B 0.026065f
C257 VP.n63 B 0.038787f
C258 VP.t9 B 2.38453f
C259 VP.n64 B 0.831056f
C260 VP.n65 B 0.031128f
C261 VP.n66 B 0.020916f
C262 VP.n67 B 0.020916f
C263 VP.n68 B 0.020916f
C264 VP.n69 B 0.038787f
C265 VP.n70 B 0.031852f
C266 VP.n71 B 0.028958f
C267 VP.n72 B 0.020916f
C268 VP.n73 B 0.020916f
C269 VP.n74 B 0.020916f
C270 VP.n75 B 0.029213f
C271 VP.n76 B 0.831056f
C272 VP.n77 B 0.029213f
C273 VP.n78 B 0.038787f
C274 VP.n79 B 0.020916f
C275 VP.n80 B 0.020916f
C276 VP.n81 B 0.020916f
C277 VP.n82 B 0.031852f
C278 VP.n83 B 0.038787f
C279 VP.n84 B 0.027298f
C280 VP.n85 B 0.020916f
C281 VP.n86 B 0.020916f
C282 VP.n87 B 0.031128f
C283 VP.n88 B 0.038787f
C284 VP.n89 B 0.026065f
C285 VP.n90 B 0.020916f
C286 VP.n91 B 0.020916f
C287 VP.n92 B 0.020916f
C288 VP.n93 B 0.038787f
C289 VP.n94 B 0.025383f
C290 VP.n95 B 0.8983f
C291 VP.n96 B 0.035513f
.ends

