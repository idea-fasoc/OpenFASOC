* NGSPICE file created from diff_pair_sample_1202.ext - technology: sky130A

.subckt diff_pair_sample_1202 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=7.7259 ps=40.4 w=19.81 l=2.48
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=7.7259 ps=40.4 w=19.81 l=2.48
X2 B.t11 B.t9 B.t10 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=2.48
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=7.7259 ps=40.4 w=19.81 l=2.48
X4 B.t8 B.t6 B.t7 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=2.48
X5 B.t5 B.t3 B.t4 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=2.48
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=7.7259 ps=40.4 w=19.81 l=2.48
X7 B.t2 B.t0 B.t1 w_n2094_n4930# sky130_fd_pr__pfet_01v8 ad=7.7259 pd=40.4 as=0 ps=0 w=19.81 l=2.48
R0 VN VN.t1 292.031
R1 VN VN.t0 242.016
R2 VTAIL.n1 VTAIL.t1 55.2055
R3 VTAIL.n3 VTAIL.t2 55.2053
R4 VTAIL.n0 VTAIL.t3 55.2053
R5 VTAIL.n2 VTAIL.t0 55.2053
R6 VTAIL.n1 VTAIL.n0 34.2893
R7 VTAIL.n3 VTAIL.n2 31.8669
R8 VTAIL.n2 VTAIL.n1 1.68153
R9 VTAIL VTAIL.n0 1.13412
R10 VTAIL VTAIL.n3 0.547914
R11 VDD2.n0 VDD2.t1 117.466
R12 VDD2.n0 VDD2.t0 71.884
R13 VDD2 VDD2.n0 0.664293
R14 VP.n0 VP.t0 291.935
R15 VP.n0 VP.t1 241.679
R16 VP VP.n0 0.336784
R17 VDD1 VDD1.t0 118.597
R18 VDD1 VDD1.t1 72.5478
R19 B.n443 B.n442 585
R20 B.n441 B.n114 585
R21 B.n440 B.n439 585
R22 B.n438 B.n115 585
R23 B.n437 B.n436 585
R24 B.n435 B.n116 585
R25 B.n434 B.n433 585
R26 B.n432 B.n117 585
R27 B.n431 B.n430 585
R28 B.n429 B.n118 585
R29 B.n428 B.n427 585
R30 B.n426 B.n119 585
R31 B.n425 B.n424 585
R32 B.n423 B.n120 585
R33 B.n422 B.n421 585
R34 B.n420 B.n121 585
R35 B.n419 B.n418 585
R36 B.n417 B.n122 585
R37 B.n416 B.n415 585
R38 B.n414 B.n123 585
R39 B.n413 B.n412 585
R40 B.n411 B.n124 585
R41 B.n410 B.n409 585
R42 B.n408 B.n125 585
R43 B.n407 B.n406 585
R44 B.n405 B.n126 585
R45 B.n404 B.n403 585
R46 B.n402 B.n127 585
R47 B.n401 B.n400 585
R48 B.n399 B.n128 585
R49 B.n398 B.n397 585
R50 B.n396 B.n129 585
R51 B.n395 B.n394 585
R52 B.n393 B.n130 585
R53 B.n392 B.n391 585
R54 B.n390 B.n131 585
R55 B.n389 B.n388 585
R56 B.n387 B.n132 585
R57 B.n386 B.n385 585
R58 B.n384 B.n133 585
R59 B.n383 B.n382 585
R60 B.n381 B.n134 585
R61 B.n380 B.n379 585
R62 B.n378 B.n135 585
R63 B.n377 B.n376 585
R64 B.n375 B.n136 585
R65 B.n374 B.n373 585
R66 B.n372 B.n137 585
R67 B.n371 B.n370 585
R68 B.n369 B.n138 585
R69 B.n368 B.n367 585
R70 B.n366 B.n139 585
R71 B.n365 B.n364 585
R72 B.n363 B.n140 585
R73 B.n362 B.n361 585
R74 B.n360 B.n141 585
R75 B.n359 B.n358 585
R76 B.n357 B.n142 585
R77 B.n356 B.n355 585
R78 B.n354 B.n143 585
R79 B.n353 B.n352 585
R80 B.n351 B.n144 585
R81 B.n350 B.n349 585
R82 B.n348 B.n145 585
R83 B.n347 B.n346 585
R84 B.n344 B.n146 585
R85 B.n343 B.n342 585
R86 B.n341 B.n149 585
R87 B.n340 B.n339 585
R88 B.n338 B.n150 585
R89 B.n337 B.n336 585
R90 B.n335 B.n151 585
R91 B.n334 B.n333 585
R92 B.n332 B.n152 585
R93 B.n330 B.n329 585
R94 B.n328 B.n155 585
R95 B.n327 B.n326 585
R96 B.n325 B.n156 585
R97 B.n324 B.n323 585
R98 B.n322 B.n157 585
R99 B.n321 B.n320 585
R100 B.n319 B.n158 585
R101 B.n318 B.n317 585
R102 B.n316 B.n159 585
R103 B.n315 B.n314 585
R104 B.n313 B.n160 585
R105 B.n312 B.n311 585
R106 B.n310 B.n161 585
R107 B.n309 B.n308 585
R108 B.n307 B.n162 585
R109 B.n306 B.n305 585
R110 B.n304 B.n163 585
R111 B.n303 B.n302 585
R112 B.n301 B.n164 585
R113 B.n300 B.n299 585
R114 B.n298 B.n165 585
R115 B.n297 B.n296 585
R116 B.n295 B.n166 585
R117 B.n294 B.n293 585
R118 B.n292 B.n167 585
R119 B.n291 B.n290 585
R120 B.n289 B.n168 585
R121 B.n288 B.n287 585
R122 B.n286 B.n169 585
R123 B.n285 B.n284 585
R124 B.n283 B.n170 585
R125 B.n282 B.n281 585
R126 B.n280 B.n171 585
R127 B.n279 B.n278 585
R128 B.n277 B.n172 585
R129 B.n276 B.n275 585
R130 B.n274 B.n173 585
R131 B.n273 B.n272 585
R132 B.n271 B.n174 585
R133 B.n270 B.n269 585
R134 B.n268 B.n175 585
R135 B.n267 B.n266 585
R136 B.n265 B.n176 585
R137 B.n264 B.n263 585
R138 B.n262 B.n177 585
R139 B.n261 B.n260 585
R140 B.n259 B.n178 585
R141 B.n258 B.n257 585
R142 B.n256 B.n179 585
R143 B.n255 B.n254 585
R144 B.n253 B.n180 585
R145 B.n252 B.n251 585
R146 B.n250 B.n181 585
R147 B.n249 B.n248 585
R148 B.n247 B.n182 585
R149 B.n246 B.n245 585
R150 B.n244 B.n183 585
R151 B.n243 B.n242 585
R152 B.n241 B.n184 585
R153 B.n240 B.n239 585
R154 B.n238 B.n185 585
R155 B.n237 B.n236 585
R156 B.n235 B.n186 585
R157 B.n234 B.n233 585
R158 B.n444 B.n113 585
R159 B.n446 B.n445 585
R160 B.n447 B.n112 585
R161 B.n449 B.n448 585
R162 B.n450 B.n111 585
R163 B.n452 B.n451 585
R164 B.n453 B.n110 585
R165 B.n455 B.n454 585
R166 B.n456 B.n109 585
R167 B.n458 B.n457 585
R168 B.n459 B.n108 585
R169 B.n461 B.n460 585
R170 B.n462 B.n107 585
R171 B.n464 B.n463 585
R172 B.n465 B.n106 585
R173 B.n467 B.n466 585
R174 B.n468 B.n105 585
R175 B.n470 B.n469 585
R176 B.n471 B.n104 585
R177 B.n473 B.n472 585
R178 B.n474 B.n103 585
R179 B.n476 B.n475 585
R180 B.n477 B.n102 585
R181 B.n479 B.n478 585
R182 B.n480 B.n101 585
R183 B.n482 B.n481 585
R184 B.n483 B.n100 585
R185 B.n485 B.n484 585
R186 B.n486 B.n99 585
R187 B.n488 B.n487 585
R188 B.n489 B.n98 585
R189 B.n491 B.n490 585
R190 B.n492 B.n97 585
R191 B.n494 B.n493 585
R192 B.n495 B.n96 585
R193 B.n497 B.n496 585
R194 B.n498 B.n95 585
R195 B.n500 B.n499 585
R196 B.n501 B.n94 585
R197 B.n503 B.n502 585
R198 B.n504 B.n93 585
R199 B.n506 B.n505 585
R200 B.n507 B.n92 585
R201 B.n509 B.n508 585
R202 B.n510 B.n91 585
R203 B.n512 B.n511 585
R204 B.n513 B.n90 585
R205 B.n515 B.n514 585
R206 B.n516 B.n89 585
R207 B.n518 B.n517 585
R208 B.n727 B.n14 585
R209 B.n726 B.n725 585
R210 B.n724 B.n15 585
R211 B.n723 B.n722 585
R212 B.n721 B.n16 585
R213 B.n720 B.n719 585
R214 B.n718 B.n17 585
R215 B.n717 B.n716 585
R216 B.n715 B.n18 585
R217 B.n714 B.n713 585
R218 B.n712 B.n19 585
R219 B.n711 B.n710 585
R220 B.n709 B.n20 585
R221 B.n708 B.n707 585
R222 B.n706 B.n21 585
R223 B.n705 B.n704 585
R224 B.n703 B.n22 585
R225 B.n702 B.n701 585
R226 B.n700 B.n23 585
R227 B.n699 B.n698 585
R228 B.n697 B.n24 585
R229 B.n696 B.n695 585
R230 B.n694 B.n25 585
R231 B.n693 B.n692 585
R232 B.n691 B.n26 585
R233 B.n690 B.n689 585
R234 B.n688 B.n27 585
R235 B.n687 B.n686 585
R236 B.n685 B.n28 585
R237 B.n684 B.n683 585
R238 B.n682 B.n29 585
R239 B.n681 B.n680 585
R240 B.n679 B.n30 585
R241 B.n678 B.n677 585
R242 B.n676 B.n31 585
R243 B.n675 B.n674 585
R244 B.n673 B.n32 585
R245 B.n672 B.n671 585
R246 B.n670 B.n33 585
R247 B.n669 B.n668 585
R248 B.n667 B.n34 585
R249 B.n666 B.n665 585
R250 B.n664 B.n35 585
R251 B.n663 B.n662 585
R252 B.n661 B.n36 585
R253 B.n660 B.n659 585
R254 B.n658 B.n37 585
R255 B.n657 B.n656 585
R256 B.n655 B.n38 585
R257 B.n654 B.n653 585
R258 B.n652 B.n39 585
R259 B.n651 B.n650 585
R260 B.n649 B.n40 585
R261 B.n648 B.n647 585
R262 B.n646 B.n41 585
R263 B.n645 B.n644 585
R264 B.n643 B.n42 585
R265 B.n642 B.n641 585
R266 B.n640 B.n43 585
R267 B.n639 B.n638 585
R268 B.n637 B.n44 585
R269 B.n636 B.n635 585
R270 B.n634 B.n45 585
R271 B.n633 B.n632 585
R272 B.n631 B.n46 585
R273 B.n630 B.n629 585
R274 B.n628 B.n47 585
R275 B.n627 B.n626 585
R276 B.n625 B.n51 585
R277 B.n624 B.n623 585
R278 B.n622 B.n52 585
R279 B.n621 B.n620 585
R280 B.n619 B.n53 585
R281 B.n618 B.n617 585
R282 B.n615 B.n54 585
R283 B.n614 B.n613 585
R284 B.n612 B.n57 585
R285 B.n611 B.n610 585
R286 B.n609 B.n58 585
R287 B.n608 B.n607 585
R288 B.n606 B.n59 585
R289 B.n605 B.n604 585
R290 B.n603 B.n60 585
R291 B.n602 B.n601 585
R292 B.n600 B.n61 585
R293 B.n599 B.n598 585
R294 B.n597 B.n62 585
R295 B.n596 B.n595 585
R296 B.n594 B.n63 585
R297 B.n593 B.n592 585
R298 B.n591 B.n64 585
R299 B.n590 B.n589 585
R300 B.n588 B.n65 585
R301 B.n587 B.n586 585
R302 B.n585 B.n66 585
R303 B.n584 B.n583 585
R304 B.n582 B.n67 585
R305 B.n581 B.n580 585
R306 B.n579 B.n68 585
R307 B.n578 B.n577 585
R308 B.n576 B.n69 585
R309 B.n575 B.n574 585
R310 B.n573 B.n70 585
R311 B.n572 B.n571 585
R312 B.n570 B.n71 585
R313 B.n569 B.n568 585
R314 B.n567 B.n72 585
R315 B.n566 B.n565 585
R316 B.n564 B.n73 585
R317 B.n563 B.n562 585
R318 B.n561 B.n74 585
R319 B.n560 B.n559 585
R320 B.n558 B.n75 585
R321 B.n557 B.n556 585
R322 B.n555 B.n76 585
R323 B.n554 B.n553 585
R324 B.n552 B.n77 585
R325 B.n551 B.n550 585
R326 B.n549 B.n78 585
R327 B.n548 B.n547 585
R328 B.n546 B.n79 585
R329 B.n545 B.n544 585
R330 B.n543 B.n80 585
R331 B.n542 B.n541 585
R332 B.n540 B.n81 585
R333 B.n539 B.n538 585
R334 B.n537 B.n82 585
R335 B.n536 B.n535 585
R336 B.n534 B.n83 585
R337 B.n533 B.n532 585
R338 B.n531 B.n84 585
R339 B.n530 B.n529 585
R340 B.n528 B.n85 585
R341 B.n527 B.n526 585
R342 B.n525 B.n86 585
R343 B.n524 B.n523 585
R344 B.n522 B.n87 585
R345 B.n521 B.n520 585
R346 B.n519 B.n88 585
R347 B.n729 B.n728 585
R348 B.n730 B.n13 585
R349 B.n732 B.n731 585
R350 B.n733 B.n12 585
R351 B.n735 B.n734 585
R352 B.n736 B.n11 585
R353 B.n738 B.n737 585
R354 B.n739 B.n10 585
R355 B.n741 B.n740 585
R356 B.n742 B.n9 585
R357 B.n744 B.n743 585
R358 B.n745 B.n8 585
R359 B.n747 B.n746 585
R360 B.n748 B.n7 585
R361 B.n750 B.n749 585
R362 B.n751 B.n6 585
R363 B.n753 B.n752 585
R364 B.n754 B.n5 585
R365 B.n756 B.n755 585
R366 B.n757 B.n4 585
R367 B.n759 B.n758 585
R368 B.n760 B.n3 585
R369 B.n762 B.n761 585
R370 B.n763 B.n0 585
R371 B.n2 B.n1 585
R372 B.n199 B.n198 585
R373 B.n201 B.n200 585
R374 B.n202 B.n197 585
R375 B.n204 B.n203 585
R376 B.n205 B.n196 585
R377 B.n207 B.n206 585
R378 B.n208 B.n195 585
R379 B.n210 B.n209 585
R380 B.n211 B.n194 585
R381 B.n213 B.n212 585
R382 B.n214 B.n193 585
R383 B.n216 B.n215 585
R384 B.n217 B.n192 585
R385 B.n219 B.n218 585
R386 B.n220 B.n191 585
R387 B.n222 B.n221 585
R388 B.n223 B.n190 585
R389 B.n225 B.n224 585
R390 B.n226 B.n189 585
R391 B.n228 B.n227 585
R392 B.n229 B.n188 585
R393 B.n231 B.n230 585
R394 B.n232 B.n187 585
R395 B.n233 B.n232 502.111
R396 B.n444 B.n443 502.111
R397 B.n517 B.n88 502.111
R398 B.n728 B.n727 502.111
R399 B.n153 B.t9 400.366
R400 B.n147 B.t0 400.366
R401 B.n55 B.t6 400.366
R402 B.n48 B.t3 400.366
R403 B.n765 B.n764 256.663
R404 B.n764 B.n763 235.042
R405 B.n764 B.n2 235.042
R406 B.n233 B.n186 163.367
R407 B.n237 B.n186 163.367
R408 B.n238 B.n237 163.367
R409 B.n239 B.n238 163.367
R410 B.n239 B.n184 163.367
R411 B.n243 B.n184 163.367
R412 B.n244 B.n243 163.367
R413 B.n245 B.n244 163.367
R414 B.n245 B.n182 163.367
R415 B.n249 B.n182 163.367
R416 B.n250 B.n249 163.367
R417 B.n251 B.n250 163.367
R418 B.n251 B.n180 163.367
R419 B.n255 B.n180 163.367
R420 B.n256 B.n255 163.367
R421 B.n257 B.n256 163.367
R422 B.n257 B.n178 163.367
R423 B.n261 B.n178 163.367
R424 B.n262 B.n261 163.367
R425 B.n263 B.n262 163.367
R426 B.n263 B.n176 163.367
R427 B.n267 B.n176 163.367
R428 B.n268 B.n267 163.367
R429 B.n269 B.n268 163.367
R430 B.n269 B.n174 163.367
R431 B.n273 B.n174 163.367
R432 B.n274 B.n273 163.367
R433 B.n275 B.n274 163.367
R434 B.n275 B.n172 163.367
R435 B.n279 B.n172 163.367
R436 B.n280 B.n279 163.367
R437 B.n281 B.n280 163.367
R438 B.n281 B.n170 163.367
R439 B.n285 B.n170 163.367
R440 B.n286 B.n285 163.367
R441 B.n287 B.n286 163.367
R442 B.n287 B.n168 163.367
R443 B.n291 B.n168 163.367
R444 B.n292 B.n291 163.367
R445 B.n293 B.n292 163.367
R446 B.n293 B.n166 163.367
R447 B.n297 B.n166 163.367
R448 B.n298 B.n297 163.367
R449 B.n299 B.n298 163.367
R450 B.n299 B.n164 163.367
R451 B.n303 B.n164 163.367
R452 B.n304 B.n303 163.367
R453 B.n305 B.n304 163.367
R454 B.n305 B.n162 163.367
R455 B.n309 B.n162 163.367
R456 B.n310 B.n309 163.367
R457 B.n311 B.n310 163.367
R458 B.n311 B.n160 163.367
R459 B.n315 B.n160 163.367
R460 B.n316 B.n315 163.367
R461 B.n317 B.n316 163.367
R462 B.n317 B.n158 163.367
R463 B.n321 B.n158 163.367
R464 B.n322 B.n321 163.367
R465 B.n323 B.n322 163.367
R466 B.n323 B.n156 163.367
R467 B.n327 B.n156 163.367
R468 B.n328 B.n327 163.367
R469 B.n329 B.n328 163.367
R470 B.n329 B.n152 163.367
R471 B.n334 B.n152 163.367
R472 B.n335 B.n334 163.367
R473 B.n336 B.n335 163.367
R474 B.n336 B.n150 163.367
R475 B.n340 B.n150 163.367
R476 B.n341 B.n340 163.367
R477 B.n342 B.n341 163.367
R478 B.n342 B.n146 163.367
R479 B.n347 B.n146 163.367
R480 B.n348 B.n347 163.367
R481 B.n349 B.n348 163.367
R482 B.n349 B.n144 163.367
R483 B.n353 B.n144 163.367
R484 B.n354 B.n353 163.367
R485 B.n355 B.n354 163.367
R486 B.n355 B.n142 163.367
R487 B.n359 B.n142 163.367
R488 B.n360 B.n359 163.367
R489 B.n361 B.n360 163.367
R490 B.n361 B.n140 163.367
R491 B.n365 B.n140 163.367
R492 B.n366 B.n365 163.367
R493 B.n367 B.n366 163.367
R494 B.n367 B.n138 163.367
R495 B.n371 B.n138 163.367
R496 B.n372 B.n371 163.367
R497 B.n373 B.n372 163.367
R498 B.n373 B.n136 163.367
R499 B.n377 B.n136 163.367
R500 B.n378 B.n377 163.367
R501 B.n379 B.n378 163.367
R502 B.n379 B.n134 163.367
R503 B.n383 B.n134 163.367
R504 B.n384 B.n383 163.367
R505 B.n385 B.n384 163.367
R506 B.n385 B.n132 163.367
R507 B.n389 B.n132 163.367
R508 B.n390 B.n389 163.367
R509 B.n391 B.n390 163.367
R510 B.n391 B.n130 163.367
R511 B.n395 B.n130 163.367
R512 B.n396 B.n395 163.367
R513 B.n397 B.n396 163.367
R514 B.n397 B.n128 163.367
R515 B.n401 B.n128 163.367
R516 B.n402 B.n401 163.367
R517 B.n403 B.n402 163.367
R518 B.n403 B.n126 163.367
R519 B.n407 B.n126 163.367
R520 B.n408 B.n407 163.367
R521 B.n409 B.n408 163.367
R522 B.n409 B.n124 163.367
R523 B.n413 B.n124 163.367
R524 B.n414 B.n413 163.367
R525 B.n415 B.n414 163.367
R526 B.n415 B.n122 163.367
R527 B.n419 B.n122 163.367
R528 B.n420 B.n419 163.367
R529 B.n421 B.n420 163.367
R530 B.n421 B.n120 163.367
R531 B.n425 B.n120 163.367
R532 B.n426 B.n425 163.367
R533 B.n427 B.n426 163.367
R534 B.n427 B.n118 163.367
R535 B.n431 B.n118 163.367
R536 B.n432 B.n431 163.367
R537 B.n433 B.n432 163.367
R538 B.n433 B.n116 163.367
R539 B.n437 B.n116 163.367
R540 B.n438 B.n437 163.367
R541 B.n439 B.n438 163.367
R542 B.n439 B.n114 163.367
R543 B.n443 B.n114 163.367
R544 B.n517 B.n516 163.367
R545 B.n516 B.n515 163.367
R546 B.n515 B.n90 163.367
R547 B.n511 B.n90 163.367
R548 B.n511 B.n510 163.367
R549 B.n510 B.n509 163.367
R550 B.n509 B.n92 163.367
R551 B.n505 B.n92 163.367
R552 B.n505 B.n504 163.367
R553 B.n504 B.n503 163.367
R554 B.n503 B.n94 163.367
R555 B.n499 B.n94 163.367
R556 B.n499 B.n498 163.367
R557 B.n498 B.n497 163.367
R558 B.n497 B.n96 163.367
R559 B.n493 B.n96 163.367
R560 B.n493 B.n492 163.367
R561 B.n492 B.n491 163.367
R562 B.n491 B.n98 163.367
R563 B.n487 B.n98 163.367
R564 B.n487 B.n486 163.367
R565 B.n486 B.n485 163.367
R566 B.n485 B.n100 163.367
R567 B.n481 B.n100 163.367
R568 B.n481 B.n480 163.367
R569 B.n480 B.n479 163.367
R570 B.n479 B.n102 163.367
R571 B.n475 B.n102 163.367
R572 B.n475 B.n474 163.367
R573 B.n474 B.n473 163.367
R574 B.n473 B.n104 163.367
R575 B.n469 B.n104 163.367
R576 B.n469 B.n468 163.367
R577 B.n468 B.n467 163.367
R578 B.n467 B.n106 163.367
R579 B.n463 B.n106 163.367
R580 B.n463 B.n462 163.367
R581 B.n462 B.n461 163.367
R582 B.n461 B.n108 163.367
R583 B.n457 B.n108 163.367
R584 B.n457 B.n456 163.367
R585 B.n456 B.n455 163.367
R586 B.n455 B.n110 163.367
R587 B.n451 B.n110 163.367
R588 B.n451 B.n450 163.367
R589 B.n450 B.n449 163.367
R590 B.n449 B.n112 163.367
R591 B.n445 B.n112 163.367
R592 B.n445 B.n444 163.367
R593 B.n727 B.n726 163.367
R594 B.n726 B.n15 163.367
R595 B.n722 B.n15 163.367
R596 B.n722 B.n721 163.367
R597 B.n721 B.n720 163.367
R598 B.n720 B.n17 163.367
R599 B.n716 B.n17 163.367
R600 B.n716 B.n715 163.367
R601 B.n715 B.n714 163.367
R602 B.n714 B.n19 163.367
R603 B.n710 B.n19 163.367
R604 B.n710 B.n709 163.367
R605 B.n709 B.n708 163.367
R606 B.n708 B.n21 163.367
R607 B.n704 B.n21 163.367
R608 B.n704 B.n703 163.367
R609 B.n703 B.n702 163.367
R610 B.n702 B.n23 163.367
R611 B.n698 B.n23 163.367
R612 B.n698 B.n697 163.367
R613 B.n697 B.n696 163.367
R614 B.n696 B.n25 163.367
R615 B.n692 B.n25 163.367
R616 B.n692 B.n691 163.367
R617 B.n691 B.n690 163.367
R618 B.n690 B.n27 163.367
R619 B.n686 B.n27 163.367
R620 B.n686 B.n685 163.367
R621 B.n685 B.n684 163.367
R622 B.n684 B.n29 163.367
R623 B.n680 B.n29 163.367
R624 B.n680 B.n679 163.367
R625 B.n679 B.n678 163.367
R626 B.n678 B.n31 163.367
R627 B.n674 B.n31 163.367
R628 B.n674 B.n673 163.367
R629 B.n673 B.n672 163.367
R630 B.n672 B.n33 163.367
R631 B.n668 B.n33 163.367
R632 B.n668 B.n667 163.367
R633 B.n667 B.n666 163.367
R634 B.n666 B.n35 163.367
R635 B.n662 B.n35 163.367
R636 B.n662 B.n661 163.367
R637 B.n661 B.n660 163.367
R638 B.n660 B.n37 163.367
R639 B.n656 B.n37 163.367
R640 B.n656 B.n655 163.367
R641 B.n655 B.n654 163.367
R642 B.n654 B.n39 163.367
R643 B.n650 B.n39 163.367
R644 B.n650 B.n649 163.367
R645 B.n649 B.n648 163.367
R646 B.n648 B.n41 163.367
R647 B.n644 B.n41 163.367
R648 B.n644 B.n643 163.367
R649 B.n643 B.n642 163.367
R650 B.n642 B.n43 163.367
R651 B.n638 B.n43 163.367
R652 B.n638 B.n637 163.367
R653 B.n637 B.n636 163.367
R654 B.n636 B.n45 163.367
R655 B.n632 B.n45 163.367
R656 B.n632 B.n631 163.367
R657 B.n631 B.n630 163.367
R658 B.n630 B.n47 163.367
R659 B.n626 B.n47 163.367
R660 B.n626 B.n625 163.367
R661 B.n625 B.n624 163.367
R662 B.n624 B.n52 163.367
R663 B.n620 B.n52 163.367
R664 B.n620 B.n619 163.367
R665 B.n619 B.n618 163.367
R666 B.n618 B.n54 163.367
R667 B.n613 B.n54 163.367
R668 B.n613 B.n612 163.367
R669 B.n612 B.n611 163.367
R670 B.n611 B.n58 163.367
R671 B.n607 B.n58 163.367
R672 B.n607 B.n606 163.367
R673 B.n606 B.n605 163.367
R674 B.n605 B.n60 163.367
R675 B.n601 B.n60 163.367
R676 B.n601 B.n600 163.367
R677 B.n600 B.n599 163.367
R678 B.n599 B.n62 163.367
R679 B.n595 B.n62 163.367
R680 B.n595 B.n594 163.367
R681 B.n594 B.n593 163.367
R682 B.n593 B.n64 163.367
R683 B.n589 B.n64 163.367
R684 B.n589 B.n588 163.367
R685 B.n588 B.n587 163.367
R686 B.n587 B.n66 163.367
R687 B.n583 B.n66 163.367
R688 B.n583 B.n582 163.367
R689 B.n582 B.n581 163.367
R690 B.n581 B.n68 163.367
R691 B.n577 B.n68 163.367
R692 B.n577 B.n576 163.367
R693 B.n576 B.n575 163.367
R694 B.n575 B.n70 163.367
R695 B.n571 B.n70 163.367
R696 B.n571 B.n570 163.367
R697 B.n570 B.n569 163.367
R698 B.n569 B.n72 163.367
R699 B.n565 B.n72 163.367
R700 B.n565 B.n564 163.367
R701 B.n564 B.n563 163.367
R702 B.n563 B.n74 163.367
R703 B.n559 B.n74 163.367
R704 B.n559 B.n558 163.367
R705 B.n558 B.n557 163.367
R706 B.n557 B.n76 163.367
R707 B.n553 B.n76 163.367
R708 B.n553 B.n552 163.367
R709 B.n552 B.n551 163.367
R710 B.n551 B.n78 163.367
R711 B.n547 B.n78 163.367
R712 B.n547 B.n546 163.367
R713 B.n546 B.n545 163.367
R714 B.n545 B.n80 163.367
R715 B.n541 B.n80 163.367
R716 B.n541 B.n540 163.367
R717 B.n540 B.n539 163.367
R718 B.n539 B.n82 163.367
R719 B.n535 B.n82 163.367
R720 B.n535 B.n534 163.367
R721 B.n534 B.n533 163.367
R722 B.n533 B.n84 163.367
R723 B.n529 B.n84 163.367
R724 B.n529 B.n528 163.367
R725 B.n528 B.n527 163.367
R726 B.n527 B.n86 163.367
R727 B.n523 B.n86 163.367
R728 B.n523 B.n522 163.367
R729 B.n522 B.n521 163.367
R730 B.n521 B.n88 163.367
R731 B.n728 B.n13 163.367
R732 B.n732 B.n13 163.367
R733 B.n733 B.n732 163.367
R734 B.n734 B.n733 163.367
R735 B.n734 B.n11 163.367
R736 B.n738 B.n11 163.367
R737 B.n739 B.n738 163.367
R738 B.n740 B.n739 163.367
R739 B.n740 B.n9 163.367
R740 B.n744 B.n9 163.367
R741 B.n745 B.n744 163.367
R742 B.n746 B.n745 163.367
R743 B.n746 B.n7 163.367
R744 B.n750 B.n7 163.367
R745 B.n751 B.n750 163.367
R746 B.n752 B.n751 163.367
R747 B.n752 B.n5 163.367
R748 B.n756 B.n5 163.367
R749 B.n757 B.n756 163.367
R750 B.n758 B.n757 163.367
R751 B.n758 B.n3 163.367
R752 B.n762 B.n3 163.367
R753 B.n763 B.n762 163.367
R754 B.n198 B.n2 163.367
R755 B.n201 B.n198 163.367
R756 B.n202 B.n201 163.367
R757 B.n203 B.n202 163.367
R758 B.n203 B.n196 163.367
R759 B.n207 B.n196 163.367
R760 B.n208 B.n207 163.367
R761 B.n209 B.n208 163.367
R762 B.n209 B.n194 163.367
R763 B.n213 B.n194 163.367
R764 B.n214 B.n213 163.367
R765 B.n215 B.n214 163.367
R766 B.n215 B.n192 163.367
R767 B.n219 B.n192 163.367
R768 B.n220 B.n219 163.367
R769 B.n221 B.n220 163.367
R770 B.n221 B.n190 163.367
R771 B.n225 B.n190 163.367
R772 B.n226 B.n225 163.367
R773 B.n227 B.n226 163.367
R774 B.n227 B.n188 163.367
R775 B.n231 B.n188 163.367
R776 B.n232 B.n231 163.367
R777 B.n147 B.t1 162.285
R778 B.n55 B.t8 162.285
R779 B.n153 B.t10 162.258
R780 B.n48 B.t5 162.258
R781 B.n148 B.t2 107.787
R782 B.n56 B.t7 107.787
R783 B.n154 B.t11 107.761
R784 B.n49 B.t4 107.761
R785 B.n331 B.n154 59.5399
R786 B.n345 B.n148 59.5399
R787 B.n616 B.n56 59.5399
R788 B.n50 B.n49 59.5399
R789 B.n154 B.n153 54.4975
R790 B.n148 B.n147 54.4975
R791 B.n56 B.n55 54.4975
R792 B.n49 B.n48 54.4975
R793 B.n729 B.n14 32.6249
R794 B.n519 B.n518 32.6249
R795 B.n442 B.n113 32.6249
R796 B.n234 B.n187 32.6249
R797 B B.n765 18.0485
R798 B.n730 B.n729 10.6151
R799 B.n731 B.n730 10.6151
R800 B.n731 B.n12 10.6151
R801 B.n735 B.n12 10.6151
R802 B.n736 B.n735 10.6151
R803 B.n737 B.n736 10.6151
R804 B.n737 B.n10 10.6151
R805 B.n741 B.n10 10.6151
R806 B.n742 B.n741 10.6151
R807 B.n743 B.n742 10.6151
R808 B.n743 B.n8 10.6151
R809 B.n747 B.n8 10.6151
R810 B.n748 B.n747 10.6151
R811 B.n749 B.n748 10.6151
R812 B.n749 B.n6 10.6151
R813 B.n753 B.n6 10.6151
R814 B.n754 B.n753 10.6151
R815 B.n755 B.n754 10.6151
R816 B.n755 B.n4 10.6151
R817 B.n759 B.n4 10.6151
R818 B.n760 B.n759 10.6151
R819 B.n761 B.n760 10.6151
R820 B.n761 B.n0 10.6151
R821 B.n725 B.n14 10.6151
R822 B.n725 B.n724 10.6151
R823 B.n724 B.n723 10.6151
R824 B.n723 B.n16 10.6151
R825 B.n719 B.n16 10.6151
R826 B.n719 B.n718 10.6151
R827 B.n718 B.n717 10.6151
R828 B.n717 B.n18 10.6151
R829 B.n713 B.n18 10.6151
R830 B.n713 B.n712 10.6151
R831 B.n712 B.n711 10.6151
R832 B.n711 B.n20 10.6151
R833 B.n707 B.n20 10.6151
R834 B.n707 B.n706 10.6151
R835 B.n706 B.n705 10.6151
R836 B.n705 B.n22 10.6151
R837 B.n701 B.n22 10.6151
R838 B.n701 B.n700 10.6151
R839 B.n700 B.n699 10.6151
R840 B.n699 B.n24 10.6151
R841 B.n695 B.n24 10.6151
R842 B.n695 B.n694 10.6151
R843 B.n694 B.n693 10.6151
R844 B.n693 B.n26 10.6151
R845 B.n689 B.n26 10.6151
R846 B.n689 B.n688 10.6151
R847 B.n688 B.n687 10.6151
R848 B.n687 B.n28 10.6151
R849 B.n683 B.n28 10.6151
R850 B.n683 B.n682 10.6151
R851 B.n682 B.n681 10.6151
R852 B.n681 B.n30 10.6151
R853 B.n677 B.n30 10.6151
R854 B.n677 B.n676 10.6151
R855 B.n676 B.n675 10.6151
R856 B.n675 B.n32 10.6151
R857 B.n671 B.n32 10.6151
R858 B.n671 B.n670 10.6151
R859 B.n670 B.n669 10.6151
R860 B.n669 B.n34 10.6151
R861 B.n665 B.n34 10.6151
R862 B.n665 B.n664 10.6151
R863 B.n664 B.n663 10.6151
R864 B.n663 B.n36 10.6151
R865 B.n659 B.n36 10.6151
R866 B.n659 B.n658 10.6151
R867 B.n658 B.n657 10.6151
R868 B.n657 B.n38 10.6151
R869 B.n653 B.n38 10.6151
R870 B.n653 B.n652 10.6151
R871 B.n652 B.n651 10.6151
R872 B.n651 B.n40 10.6151
R873 B.n647 B.n40 10.6151
R874 B.n647 B.n646 10.6151
R875 B.n646 B.n645 10.6151
R876 B.n645 B.n42 10.6151
R877 B.n641 B.n42 10.6151
R878 B.n641 B.n640 10.6151
R879 B.n640 B.n639 10.6151
R880 B.n639 B.n44 10.6151
R881 B.n635 B.n44 10.6151
R882 B.n635 B.n634 10.6151
R883 B.n634 B.n633 10.6151
R884 B.n633 B.n46 10.6151
R885 B.n629 B.n628 10.6151
R886 B.n628 B.n627 10.6151
R887 B.n627 B.n51 10.6151
R888 B.n623 B.n51 10.6151
R889 B.n623 B.n622 10.6151
R890 B.n622 B.n621 10.6151
R891 B.n621 B.n53 10.6151
R892 B.n617 B.n53 10.6151
R893 B.n615 B.n614 10.6151
R894 B.n614 B.n57 10.6151
R895 B.n610 B.n57 10.6151
R896 B.n610 B.n609 10.6151
R897 B.n609 B.n608 10.6151
R898 B.n608 B.n59 10.6151
R899 B.n604 B.n59 10.6151
R900 B.n604 B.n603 10.6151
R901 B.n603 B.n602 10.6151
R902 B.n602 B.n61 10.6151
R903 B.n598 B.n61 10.6151
R904 B.n598 B.n597 10.6151
R905 B.n597 B.n596 10.6151
R906 B.n596 B.n63 10.6151
R907 B.n592 B.n63 10.6151
R908 B.n592 B.n591 10.6151
R909 B.n591 B.n590 10.6151
R910 B.n590 B.n65 10.6151
R911 B.n586 B.n65 10.6151
R912 B.n586 B.n585 10.6151
R913 B.n585 B.n584 10.6151
R914 B.n584 B.n67 10.6151
R915 B.n580 B.n67 10.6151
R916 B.n580 B.n579 10.6151
R917 B.n579 B.n578 10.6151
R918 B.n578 B.n69 10.6151
R919 B.n574 B.n69 10.6151
R920 B.n574 B.n573 10.6151
R921 B.n573 B.n572 10.6151
R922 B.n572 B.n71 10.6151
R923 B.n568 B.n71 10.6151
R924 B.n568 B.n567 10.6151
R925 B.n567 B.n566 10.6151
R926 B.n566 B.n73 10.6151
R927 B.n562 B.n73 10.6151
R928 B.n562 B.n561 10.6151
R929 B.n561 B.n560 10.6151
R930 B.n560 B.n75 10.6151
R931 B.n556 B.n75 10.6151
R932 B.n556 B.n555 10.6151
R933 B.n555 B.n554 10.6151
R934 B.n554 B.n77 10.6151
R935 B.n550 B.n77 10.6151
R936 B.n550 B.n549 10.6151
R937 B.n549 B.n548 10.6151
R938 B.n548 B.n79 10.6151
R939 B.n544 B.n79 10.6151
R940 B.n544 B.n543 10.6151
R941 B.n543 B.n542 10.6151
R942 B.n542 B.n81 10.6151
R943 B.n538 B.n81 10.6151
R944 B.n538 B.n537 10.6151
R945 B.n537 B.n536 10.6151
R946 B.n536 B.n83 10.6151
R947 B.n532 B.n83 10.6151
R948 B.n532 B.n531 10.6151
R949 B.n531 B.n530 10.6151
R950 B.n530 B.n85 10.6151
R951 B.n526 B.n85 10.6151
R952 B.n526 B.n525 10.6151
R953 B.n525 B.n524 10.6151
R954 B.n524 B.n87 10.6151
R955 B.n520 B.n87 10.6151
R956 B.n520 B.n519 10.6151
R957 B.n518 B.n89 10.6151
R958 B.n514 B.n89 10.6151
R959 B.n514 B.n513 10.6151
R960 B.n513 B.n512 10.6151
R961 B.n512 B.n91 10.6151
R962 B.n508 B.n91 10.6151
R963 B.n508 B.n507 10.6151
R964 B.n507 B.n506 10.6151
R965 B.n506 B.n93 10.6151
R966 B.n502 B.n93 10.6151
R967 B.n502 B.n501 10.6151
R968 B.n501 B.n500 10.6151
R969 B.n500 B.n95 10.6151
R970 B.n496 B.n95 10.6151
R971 B.n496 B.n495 10.6151
R972 B.n495 B.n494 10.6151
R973 B.n494 B.n97 10.6151
R974 B.n490 B.n97 10.6151
R975 B.n490 B.n489 10.6151
R976 B.n489 B.n488 10.6151
R977 B.n488 B.n99 10.6151
R978 B.n484 B.n99 10.6151
R979 B.n484 B.n483 10.6151
R980 B.n483 B.n482 10.6151
R981 B.n482 B.n101 10.6151
R982 B.n478 B.n101 10.6151
R983 B.n478 B.n477 10.6151
R984 B.n477 B.n476 10.6151
R985 B.n476 B.n103 10.6151
R986 B.n472 B.n103 10.6151
R987 B.n472 B.n471 10.6151
R988 B.n471 B.n470 10.6151
R989 B.n470 B.n105 10.6151
R990 B.n466 B.n105 10.6151
R991 B.n466 B.n465 10.6151
R992 B.n465 B.n464 10.6151
R993 B.n464 B.n107 10.6151
R994 B.n460 B.n107 10.6151
R995 B.n460 B.n459 10.6151
R996 B.n459 B.n458 10.6151
R997 B.n458 B.n109 10.6151
R998 B.n454 B.n109 10.6151
R999 B.n454 B.n453 10.6151
R1000 B.n453 B.n452 10.6151
R1001 B.n452 B.n111 10.6151
R1002 B.n448 B.n111 10.6151
R1003 B.n448 B.n447 10.6151
R1004 B.n447 B.n446 10.6151
R1005 B.n446 B.n113 10.6151
R1006 B.n199 B.n1 10.6151
R1007 B.n200 B.n199 10.6151
R1008 B.n200 B.n197 10.6151
R1009 B.n204 B.n197 10.6151
R1010 B.n205 B.n204 10.6151
R1011 B.n206 B.n205 10.6151
R1012 B.n206 B.n195 10.6151
R1013 B.n210 B.n195 10.6151
R1014 B.n211 B.n210 10.6151
R1015 B.n212 B.n211 10.6151
R1016 B.n212 B.n193 10.6151
R1017 B.n216 B.n193 10.6151
R1018 B.n217 B.n216 10.6151
R1019 B.n218 B.n217 10.6151
R1020 B.n218 B.n191 10.6151
R1021 B.n222 B.n191 10.6151
R1022 B.n223 B.n222 10.6151
R1023 B.n224 B.n223 10.6151
R1024 B.n224 B.n189 10.6151
R1025 B.n228 B.n189 10.6151
R1026 B.n229 B.n228 10.6151
R1027 B.n230 B.n229 10.6151
R1028 B.n230 B.n187 10.6151
R1029 B.n235 B.n234 10.6151
R1030 B.n236 B.n235 10.6151
R1031 B.n236 B.n185 10.6151
R1032 B.n240 B.n185 10.6151
R1033 B.n241 B.n240 10.6151
R1034 B.n242 B.n241 10.6151
R1035 B.n242 B.n183 10.6151
R1036 B.n246 B.n183 10.6151
R1037 B.n247 B.n246 10.6151
R1038 B.n248 B.n247 10.6151
R1039 B.n248 B.n181 10.6151
R1040 B.n252 B.n181 10.6151
R1041 B.n253 B.n252 10.6151
R1042 B.n254 B.n253 10.6151
R1043 B.n254 B.n179 10.6151
R1044 B.n258 B.n179 10.6151
R1045 B.n259 B.n258 10.6151
R1046 B.n260 B.n259 10.6151
R1047 B.n260 B.n177 10.6151
R1048 B.n264 B.n177 10.6151
R1049 B.n265 B.n264 10.6151
R1050 B.n266 B.n265 10.6151
R1051 B.n266 B.n175 10.6151
R1052 B.n270 B.n175 10.6151
R1053 B.n271 B.n270 10.6151
R1054 B.n272 B.n271 10.6151
R1055 B.n272 B.n173 10.6151
R1056 B.n276 B.n173 10.6151
R1057 B.n277 B.n276 10.6151
R1058 B.n278 B.n277 10.6151
R1059 B.n278 B.n171 10.6151
R1060 B.n282 B.n171 10.6151
R1061 B.n283 B.n282 10.6151
R1062 B.n284 B.n283 10.6151
R1063 B.n284 B.n169 10.6151
R1064 B.n288 B.n169 10.6151
R1065 B.n289 B.n288 10.6151
R1066 B.n290 B.n289 10.6151
R1067 B.n290 B.n167 10.6151
R1068 B.n294 B.n167 10.6151
R1069 B.n295 B.n294 10.6151
R1070 B.n296 B.n295 10.6151
R1071 B.n296 B.n165 10.6151
R1072 B.n300 B.n165 10.6151
R1073 B.n301 B.n300 10.6151
R1074 B.n302 B.n301 10.6151
R1075 B.n302 B.n163 10.6151
R1076 B.n306 B.n163 10.6151
R1077 B.n307 B.n306 10.6151
R1078 B.n308 B.n307 10.6151
R1079 B.n308 B.n161 10.6151
R1080 B.n312 B.n161 10.6151
R1081 B.n313 B.n312 10.6151
R1082 B.n314 B.n313 10.6151
R1083 B.n314 B.n159 10.6151
R1084 B.n318 B.n159 10.6151
R1085 B.n319 B.n318 10.6151
R1086 B.n320 B.n319 10.6151
R1087 B.n320 B.n157 10.6151
R1088 B.n324 B.n157 10.6151
R1089 B.n325 B.n324 10.6151
R1090 B.n326 B.n325 10.6151
R1091 B.n326 B.n155 10.6151
R1092 B.n330 B.n155 10.6151
R1093 B.n333 B.n332 10.6151
R1094 B.n333 B.n151 10.6151
R1095 B.n337 B.n151 10.6151
R1096 B.n338 B.n337 10.6151
R1097 B.n339 B.n338 10.6151
R1098 B.n339 B.n149 10.6151
R1099 B.n343 B.n149 10.6151
R1100 B.n344 B.n343 10.6151
R1101 B.n346 B.n145 10.6151
R1102 B.n350 B.n145 10.6151
R1103 B.n351 B.n350 10.6151
R1104 B.n352 B.n351 10.6151
R1105 B.n352 B.n143 10.6151
R1106 B.n356 B.n143 10.6151
R1107 B.n357 B.n356 10.6151
R1108 B.n358 B.n357 10.6151
R1109 B.n358 B.n141 10.6151
R1110 B.n362 B.n141 10.6151
R1111 B.n363 B.n362 10.6151
R1112 B.n364 B.n363 10.6151
R1113 B.n364 B.n139 10.6151
R1114 B.n368 B.n139 10.6151
R1115 B.n369 B.n368 10.6151
R1116 B.n370 B.n369 10.6151
R1117 B.n370 B.n137 10.6151
R1118 B.n374 B.n137 10.6151
R1119 B.n375 B.n374 10.6151
R1120 B.n376 B.n375 10.6151
R1121 B.n376 B.n135 10.6151
R1122 B.n380 B.n135 10.6151
R1123 B.n381 B.n380 10.6151
R1124 B.n382 B.n381 10.6151
R1125 B.n382 B.n133 10.6151
R1126 B.n386 B.n133 10.6151
R1127 B.n387 B.n386 10.6151
R1128 B.n388 B.n387 10.6151
R1129 B.n388 B.n131 10.6151
R1130 B.n392 B.n131 10.6151
R1131 B.n393 B.n392 10.6151
R1132 B.n394 B.n393 10.6151
R1133 B.n394 B.n129 10.6151
R1134 B.n398 B.n129 10.6151
R1135 B.n399 B.n398 10.6151
R1136 B.n400 B.n399 10.6151
R1137 B.n400 B.n127 10.6151
R1138 B.n404 B.n127 10.6151
R1139 B.n405 B.n404 10.6151
R1140 B.n406 B.n405 10.6151
R1141 B.n406 B.n125 10.6151
R1142 B.n410 B.n125 10.6151
R1143 B.n411 B.n410 10.6151
R1144 B.n412 B.n411 10.6151
R1145 B.n412 B.n123 10.6151
R1146 B.n416 B.n123 10.6151
R1147 B.n417 B.n416 10.6151
R1148 B.n418 B.n417 10.6151
R1149 B.n418 B.n121 10.6151
R1150 B.n422 B.n121 10.6151
R1151 B.n423 B.n422 10.6151
R1152 B.n424 B.n423 10.6151
R1153 B.n424 B.n119 10.6151
R1154 B.n428 B.n119 10.6151
R1155 B.n429 B.n428 10.6151
R1156 B.n430 B.n429 10.6151
R1157 B.n430 B.n117 10.6151
R1158 B.n434 B.n117 10.6151
R1159 B.n435 B.n434 10.6151
R1160 B.n436 B.n435 10.6151
R1161 B.n436 B.n115 10.6151
R1162 B.n440 B.n115 10.6151
R1163 B.n441 B.n440 10.6151
R1164 B.n442 B.n441 10.6151
R1165 B.n765 B.n0 8.11757
R1166 B.n765 B.n1 8.11757
R1167 B.n629 B.n50 6.5566
R1168 B.n617 B.n616 6.5566
R1169 B.n332 B.n331 6.5566
R1170 B.n345 B.n344 6.5566
R1171 B.n50 B.n46 4.05904
R1172 B.n616 B.n615 4.05904
R1173 B.n331 B.n330 4.05904
R1174 B.n346 B.n345 4.05904
C0 VN w_n2094_n4930# 3.02735f
C1 VDD1 VP 4.5711f
C2 VDD1 VDD2 0.661173f
C3 w_n2094_n4930# B 10.8693f
C4 w_n2094_n4930# VTAIL 3.86957f
C5 VN B 1.12137f
C6 VN VTAIL 3.69748f
C7 VDD2 VP 0.328676f
C8 VDD1 w_n2094_n4930# 2.31126f
C9 VTAIL B 5.34364f
C10 VN VDD1 0.148067f
C11 VDD1 B 2.30433f
C12 w_n2094_n4930# VP 3.29382f
C13 w_n2094_n4930# VDD2 2.3357f
C14 VDD1 VTAIL 7.13192f
C15 VN VP 6.84411f
C16 VN VDD2 4.3945f
C17 VP B 1.55899f
C18 VDD2 B 2.33334f
C19 VTAIL VP 3.7119f
C20 VTAIL VDD2 7.17969f
C21 VDD2 VSUBS 1.169801f
C22 VDD1 VSUBS 6.87782f
C23 VTAIL VSUBS 1.299369f
C24 VN VSUBS 9.41134f
C25 VP VSUBS 1.932106f
C26 B VSUBS 4.48264f
C27 w_n2094_n4930# VSUBS 0.126067p
C28 B.n0 VSUBS 0.006002f
C29 B.n1 VSUBS 0.006002f
C30 B.n2 VSUBS 0.008876f
C31 B.n3 VSUBS 0.006802f
C32 B.n4 VSUBS 0.006802f
C33 B.n5 VSUBS 0.006802f
C34 B.n6 VSUBS 0.006802f
C35 B.n7 VSUBS 0.006802f
C36 B.n8 VSUBS 0.006802f
C37 B.n9 VSUBS 0.006802f
C38 B.n10 VSUBS 0.006802f
C39 B.n11 VSUBS 0.006802f
C40 B.n12 VSUBS 0.006802f
C41 B.n13 VSUBS 0.006802f
C42 B.n14 VSUBS 0.016463f
C43 B.n15 VSUBS 0.006802f
C44 B.n16 VSUBS 0.006802f
C45 B.n17 VSUBS 0.006802f
C46 B.n18 VSUBS 0.006802f
C47 B.n19 VSUBS 0.006802f
C48 B.n20 VSUBS 0.006802f
C49 B.n21 VSUBS 0.006802f
C50 B.n22 VSUBS 0.006802f
C51 B.n23 VSUBS 0.006802f
C52 B.n24 VSUBS 0.006802f
C53 B.n25 VSUBS 0.006802f
C54 B.n26 VSUBS 0.006802f
C55 B.n27 VSUBS 0.006802f
C56 B.n28 VSUBS 0.006802f
C57 B.n29 VSUBS 0.006802f
C58 B.n30 VSUBS 0.006802f
C59 B.n31 VSUBS 0.006802f
C60 B.n32 VSUBS 0.006802f
C61 B.n33 VSUBS 0.006802f
C62 B.n34 VSUBS 0.006802f
C63 B.n35 VSUBS 0.006802f
C64 B.n36 VSUBS 0.006802f
C65 B.n37 VSUBS 0.006802f
C66 B.n38 VSUBS 0.006802f
C67 B.n39 VSUBS 0.006802f
C68 B.n40 VSUBS 0.006802f
C69 B.n41 VSUBS 0.006802f
C70 B.n42 VSUBS 0.006802f
C71 B.n43 VSUBS 0.006802f
C72 B.n44 VSUBS 0.006802f
C73 B.n45 VSUBS 0.006802f
C74 B.n46 VSUBS 0.004701f
C75 B.n47 VSUBS 0.006802f
C76 B.t4 VSUBS 0.653974f
C77 B.t5 VSUBS 0.674114f
C78 B.t3 VSUBS 2.09617f
C79 B.n48 VSUBS 0.368732f
C80 B.n49 VSUBS 0.069665f
C81 B.n50 VSUBS 0.015759f
C82 B.n51 VSUBS 0.006802f
C83 B.n52 VSUBS 0.006802f
C84 B.n53 VSUBS 0.006802f
C85 B.n54 VSUBS 0.006802f
C86 B.t7 VSUBS 0.653946f
C87 B.t8 VSUBS 0.674092f
C88 B.t6 VSUBS 2.09617f
C89 B.n55 VSUBS 0.368754f
C90 B.n56 VSUBS 0.069693f
C91 B.n57 VSUBS 0.006802f
C92 B.n58 VSUBS 0.006802f
C93 B.n59 VSUBS 0.006802f
C94 B.n60 VSUBS 0.006802f
C95 B.n61 VSUBS 0.006802f
C96 B.n62 VSUBS 0.006802f
C97 B.n63 VSUBS 0.006802f
C98 B.n64 VSUBS 0.006802f
C99 B.n65 VSUBS 0.006802f
C100 B.n66 VSUBS 0.006802f
C101 B.n67 VSUBS 0.006802f
C102 B.n68 VSUBS 0.006802f
C103 B.n69 VSUBS 0.006802f
C104 B.n70 VSUBS 0.006802f
C105 B.n71 VSUBS 0.006802f
C106 B.n72 VSUBS 0.006802f
C107 B.n73 VSUBS 0.006802f
C108 B.n74 VSUBS 0.006802f
C109 B.n75 VSUBS 0.006802f
C110 B.n76 VSUBS 0.006802f
C111 B.n77 VSUBS 0.006802f
C112 B.n78 VSUBS 0.006802f
C113 B.n79 VSUBS 0.006802f
C114 B.n80 VSUBS 0.006802f
C115 B.n81 VSUBS 0.006802f
C116 B.n82 VSUBS 0.006802f
C117 B.n83 VSUBS 0.006802f
C118 B.n84 VSUBS 0.006802f
C119 B.n85 VSUBS 0.006802f
C120 B.n86 VSUBS 0.006802f
C121 B.n87 VSUBS 0.006802f
C122 B.n88 VSUBS 0.016463f
C123 B.n89 VSUBS 0.006802f
C124 B.n90 VSUBS 0.006802f
C125 B.n91 VSUBS 0.006802f
C126 B.n92 VSUBS 0.006802f
C127 B.n93 VSUBS 0.006802f
C128 B.n94 VSUBS 0.006802f
C129 B.n95 VSUBS 0.006802f
C130 B.n96 VSUBS 0.006802f
C131 B.n97 VSUBS 0.006802f
C132 B.n98 VSUBS 0.006802f
C133 B.n99 VSUBS 0.006802f
C134 B.n100 VSUBS 0.006802f
C135 B.n101 VSUBS 0.006802f
C136 B.n102 VSUBS 0.006802f
C137 B.n103 VSUBS 0.006802f
C138 B.n104 VSUBS 0.006802f
C139 B.n105 VSUBS 0.006802f
C140 B.n106 VSUBS 0.006802f
C141 B.n107 VSUBS 0.006802f
C142 B.n108 VSUBS 0.006802f
C143 B.n109 VSUBS 0.006802f
C144 B.n110 VSUBS 0.006802f
C145 B.n111 VSUBS 0.006802f
C146 B.n112 VSUBS 0.006802f
C147 B.n113 VSUBS 0.016149f
C148 B.n114 VSUBS 0.006802f
C149 B.n115 VSUBS 0.006802f
C150 B.n116 VSUBS 0.006802f
C151 B.n117 VSUBS 0.006802f
C152 B.n118 VSUBS 0.006802f
C153 B.n119 VSUBS 0.006802f
C154 B.n120 VSUBS 0.006802f
C155 B.n121 VSUBS 0.006802f
C156 B.n122 VSUBS 0.006802f
C157 B.n123 VSUBS 0.006802f
C158 B.n124 VSUBS 0.006802f
C159 B.n125 VSUBS 0.006802f
C160 B.n126 VSUBS 0.006802f
C161 B.n127 VSUBS 0.006802f
C162 B.n128 VSUBS 0.006802f
C163 B.n129 VSUBS 0.006802f
C164 B.n130 VSUBS 0.006802f
C165 B.n131 VSUBS 0.006802f
C166 B.n132 VSUBS 0.006802f
C167 B.n133 VSUBS 0.006802f
C168 B.n134 VSUBS 0.006802f
C169 B.n135 VSUBS 0.006802f
C170 B.n136 VSUBS 0.006802f
C171 B.n137 VSUBS 0.006802f
C172 B.n138 VSUBS 0.006802f
C173 B.n139 VSUBS 0.006802f
C174 B.n140 VSUBS 0.006802f
C175 B.n141 VSUBS 0.006802f
C176 B.n142 VSUBS 0.006802f
C177 B.n143 VSUBS 0.006802f
C178 B.n144 VSUBS 0.006802f
C179 B.n145 VSUBS 0.006802f
C180 B.n146 VSUBS 0.006802f
C181 B.t2 VSUBS 0.653946f
C182 B.t1 VSUBS 0.674092f
C183 B.t0 VSUBS 2.09617f
C184 B.n147 VSUBS 0.368754f
C185 B.n148 VSUBS 0.069693f
C186 B.n149 VSUBS 0.006802f
C187 B.n150 VSUBS 0.006802f
C188 B.n151 VSUBS 0.006802f
C189 B.n152 VSUBS 0.006802f
C190 B.t11 VSUBS 0.653974f
C191 B.t10 VSUBS 0.674114f
C192 B.t9 VSUBS 2.09617f
C193 B.n153 VSUBS 0.368732f
C194 B.n154 VSUBS 0.069665f
C195 B.n155 VSUBS 0.006802f
C196 B.n156 VSUBS 0.006802f
C197 B.n157 VSUBS 0.006802f
C198 B.n158 VSUBS 0.006802f
C199 B.n159 VSUBS 0.006802f
C200 B.n160 VSUBS 0.006802f
C201 B.n161 VSUBS 0.006802f
C202 B.n162 VSUBS 0.006802f
C203 B.n163 VSUBS 0.006802f
C204 B.n164 VSUBS 0.006802f
C205 B.n165 VSUBS 0.006802f
C206 B.n166 VSUBS 0.006802f
C207 B.n167 VSUBS 0.006802f
C208 B.n168 VSUBS 0.006802f
C209 B.n169 VSUBS 0.006802f
C210 B.n170 VSUBS 0.006802f
C211 B.n171 VSUBS 0.006802f
C212 B.n172 VSUBS 0.006802f
C213 B.n173 VSUBS 0.006802f
C214 B.n174 VSUBS 0.006802f
C215 B.n175 VSUBS 0.006802f
C216 B.n176 VSUBS 0.006802f
C217 B.n177 VSUBS 0.006802f
C218 B.n178 VSUBS 0.006802f
C219 B.n179 VSUBS 0.006802f
C220 B.n180 VSUBS 0.006802f
C221 B.n181 VSUBS 0.006802f
C222 B.n182 VSUBS 0.006802f
C223 B.n183 VSUBS 0.006802f
C224 B.n184 VSUBS 0.006802f
C225 B.n185 VSUBS 0.006802f
C226 B.n186 VSUBS 0.006802f
C227 B.n187 VSUBS 0.015345f
C228 B.n188 VSUBS 0.006802f
C229 B.n189 VSUBS 0.006802f
C230 B.n190 VSUBS 0.006802f
C231 B.n191 VSUBS 0.006802f
C232 B.n192 VSUBS 0.006802f
C233 B.n193 VSUBS 0.006802f
C234 B.n194 VSUBS 0.006802f
C235 B.n195 VSUBS 0.006802f
C236 B.n196 VSUBS 0.006802f
C237 B.n197 VSUBS 0.006802f
C238 B.n198 VSUBS 0.006802f
C239 B.n199 VSUBS 0.006802f
C240 B.n200 VSUBS 0.006802f
C241 B.n201 VSUBS 0.006802f
C242 B.n202 VSUBS 0.006802f
C243 B.n203 VSUBS 0.006802f
C244 B.n204 VSUBS 0.006802f
C245 B.n205 VSUBS 0.006802f
C246 B.n206 VSUBS 0.006802f
C247 B.n207 VSUBS 0.006802f
C248 B.n208 VSUBS 0.006802f
C249 B.n209 VSUBS 0.006802f
C250 B.n210 VSUBS 0.006802f
C251 B.n211 VSUBS 0.006802f
C252 B.n212 VSUBS 0.006802f
C253 B.n213 VSUBS 0.006802f
C254 B.n214 VSUBS 0.006802f
C255 B.n215 VSUBS 0.006802f
C256 B.n216 VSUBS 0.006802f
C257 B.n217 VSUBS 0.006802f
C258 B.n218 VSUBS 0.006802f
C259 B.n219 VSUBS 0.006802f
C260 B.n220 VSUBS 0.006802f
C261 B.n221 VSUBS 0.006802f
C262 B.n222 VSUBS 0.006802f
C263 B.n223 VSUBS 0.006802f
C264 B.n224 VSUBS 0.006802f
C265 B.n225 VSUBS 0.006802f
C266 B.n226 VSUBS 0.006802f
C267 B.n227 VSUBS 0.006802f
C268 B.n228 VSUBS 0.006802f
C269 B.n229 VSUBS 0.006802f
C270 B.n230 VSUBS 0.006802f
C271 B.n231 VSUBS 0.006802f
C272 B.n232 VSUBS 0.015345f
C273 B.n233 VSUBS 0.016463f
C274 B.n234 VSUBS 0.016463f
C275 B.n235 VSUBS 0.006802f
C276 B.n236 VSUBS 0.006802f
C277 B.n237 VSUBS 0.006802f
C278 B.n238 VSUBS 0.006802f
C279 B.n239 VSUBS 0.006802f
C280 B.n240 VSUBS 0.006802f
C281 B.n241 VSUBS 0.006802f
C282 B.n242 VSUBS 0.006802f
C283 B.n243 VSUBS 0.006802f
C284 B.n244 VSUBS 0.006802f
C285 B.n245 VSUBS 0.006802f
C286 B.n246 VSUBS 0.006802f
C287 B.n247 VSUBS 0.006802f
C288 B.n248 VSUBS 0.006802f
C289 B.n249 VSUBS 0.006802f
C290 B.n250 VSUBS 0.006802f
C291 B.n251 VSUBS 0.006802f
C292 B.n252 VSUBS 0.006802f
C293 B.n253 VSUBS 0.006802f
C294 B.n254 VSUBS 0.006802f
C295 B.n255 VSUBS 0.006802f
C296 B.n256 VSUBS 0.006802f
C297 B.n257 VSUBS 0.006802f
C298 B.n258 VSUBS 0.006802f
C299 B.n259 VSUBS 0.006802f
C300 B.n260 VSUBS 0.006802f
C301 B.n261 VSUBS 0.006802f
C302 B.n262 VSUBS 0.006802f
C303 B.n263 VSUBS 0.006802f
C304 B.n264 VSUBS 0.006802f
C305 B.n265 VSUBS 0.006802f
C306 B.n266 VSUBS 0.006802f
C307 B.n267 VSUBS 0.006802f
C308 B.n268 VSUBS 0.006802f
C309 B.n269 VSUBS 0.006802f
C310 B.n270 VSUBS 0.006802f
C311 B.n271 VSUBS 0.006802f
C312 B.n272 VSUBS 0.006802f
C313 B.n273 VSUBS 0.006802f
C314 B.n274 VSUBS 0.006802f
C315 B.n275 VSUBS 0.006802f
C316 B.n276 VSUBS 0.006802f
C317 B.n277 VSUBS 0.006802f
C318 B.n278 VSUBS 0.006802f
C319 B.n279 VSUBS 0.006802f
C320 B.n280 VSUBS 0.006802f
C321 B.n281 VSUBS 0.006802f
C322 B.n282 VSUBS 0.006802f
C323 B.n283 VSUBS 0.006802f
C324 B.n284 VSUBS 0.006802f
C325 B.n285 VSUBS 0.006802f
C326 B.n286 VSUBS 0.006802f
C327 B.n287 VSUBS 0.006802f
C328 B.n288 VSUBS 0.006802f
C329 B.n289 VSUBS 0.006802f
C330 B.n290 VSUBS 0.006802f
C331 B.n291 VSUBS 0.006802f
C332 B.n292 VSUBS 0.006802f
C333 B.n293 VSUBS 0.006802f
C334 B.n294 VSUBS 0.006802f
C335 B.n295 VSUBS 0.006802f
C336 B.n296 VSUBS 0.006802f
C337 B.n297 VSUBS 0.006802f
C338 B.n298 VSUBS 0.006802f
C339 B.n299 VSUBS 0.006802f
C340 B.n300 VSUBS 0.006802f
C341 B.n301 VSUBS 0.006802f
C342 B.n302 VSUBS 0.006802f
C343 B.n303 VSUBS 0.006802f
C344 B.n304 VSUBS 0.006802f
C345 B.n305 VSUBS 0.006802f
C346 B.n306 VSUBS 0.006802f
C347 B.n307 VSUBS 0.006802f
C348 B.n308 VSUBS 0.006802f
C349 B.n309 VSUBS 0.006802f
C350 B.n310 VSUBS 0.006802f
C351 B.n311 VSUBS 0.006802f
C352 B.n312 VSUBS 0.006802f
C353 B.n313 VSUBS 0.006802f
C354 B.n314 VSUBS 0.006802f
C355 B.n315 VSUBS 0.006802f
C356 B.n316 VSUBS 0.006802f
C357 B.n317 VSUBS 0.006802f
C358 B.n318 VSUBS 0.006802f
C359 B.n319 VSUBS 0.006802f
C360 B.n320 VSUBS 0.006802f
C361 B.n321 VSUBS 0.006802f
C362 B.n322 VSUBS 0.006802f
C363 B.n323 VSUBS 0.006802f
C364 B.n324 VSUBS 0.006802f
C365 B.n325 VSUBS 0.006802f
C366 B.n326 VSUBS 0.006802f
C367 B.n327 VSUBS 0.006802f
C368 B.n328 VSUBS 0.006802f
C369 B.n329 VSUBS 0.006802f
C370 B.n330 VSUBS 0.004701f
C371 B.n331 VSUBS 0.015759f
C372 B.n332 VSUBS 0.005501f
C373 B.n333 VSUBS 0.006802f
C374 B.n334 VSUBS 0.006802f
C375 B.n335 VSUBS 0.006802f
C376 B.n336 VSUBS 0.006802f
C377 B.n337 VSUBS 0.006802f
C378 B.n338 VSUBS 0.006802f
C379 B.n339 VSUBS 0.006802f
C380 B.n340 VSUBS 0.006802f
C381 B.n341 VSUBS 0.006802f
C382 B.n342 VSUBS 0.006802f
C383 B.n343 VSUBS 0.006802f
C384 B.n344 VSUBS 0.005501f
C385 B.n345 VSUBS 0.015759f
C386 B.n346 VSUBS 0.004701f
C387 B.n347 VSUBS 0.006802f
C388 B.n348 VSUBS 0.006802f
C389 B.n349 VSUBS 0.006802f
C390 B.n350 VSUBS 0.006802f
C391 B.n351 VSUBS 0.006802f
C392 B.n352 VSUBS 0.006802f
C393 B.n353 VSUBS 0.006802f
C394 B.n354 VSUBS 0.006802f
C395 B.n355 VSUBS 0.006802f
C396 B.n356 VSUBS 0.006802f
C397 B.n357 VSUBS 0.006802f
C398 B.n358 VSUBS 0.006802f
C399 B.n359 VSUBS 0.006802f
C400 B.n360 VSUBS 0.006802f
C401 B.n361 VSUBS 0.006802f
C402 B.n362 VSUBS 0.006802f
C403 B.n363 VSUBS 0.006802f
C404 B.n364 VSUBS 0.006802f
C405 B.n365 VSUBS 0.006802f
C406 B.n366 VSUBS 0.006802f
C407 B.n367 VSUBS 0.006802f
C408 B.n368 VSUBS 0.006802f
C409 B.n369 VSUBS 0.006802f
C410 B.n370 VSUBS 0.006802f
C411 B.n371 VSUBS 0.006802f
C412 B.n372 VSUBS 0.006802f
C413 B.n373 VSUBS 0.006802f
C414 B.n374 VSUBS 0.006802f
C415 B.n375 VSUBS 0.006802f
C416 B.n376 VSUBS 0.006802f
C417 B.n377 VSUBS 0.006802f
C418 B.n378 VSUBS 0.006802f
C419 B.n379 VSUBS 0.006802f
C420 B.n380 VSUBS 0.006802f
C421 B.n381 VSUBS 0.006802f
C422 B.n382 VSUBS 0.006802f
C423 B.n383 VSUBS 0.006802f
C424 B.n384 VSUBS 0.006802f
C425 B.n385 VSUBS 0.006802f
C426 B.n386 VSUBS 0.006802f
C427 B.n387 VSUBS 0.006802f
C428 B.n388 VSUBS 0.006802f
C429 B.n389 VSUBS 0.006802f
C430 B.n390 VSUBS 0.006802f
C431 B.n391 VSUBS 0.006802f
C432 B.n392 VSUBS 0.006802f
C433 B.n393 VSUBS 0.006802f
C434 B.n394 VSUBS 0.006802f
C435 B.n395 VSUBS 0.006802f
C436 B.n396 VSUBS 0.006802f
C437 B.n397 VSUBS 0.006802f
C438 B.n398 VSUBS 0.006802f
C439 B.n399 VSUBS 0.006802f
C440 B.n400 VSUBS 0.006802f
C441 B.n401 VSUBS 0.006802f
C442 B.n402 VSUBS 0.006802f
C443 B.n403 VSUBS 0.006802f
C444 B.n404 VSUBS 0.006802f
C445 B.n405 VSUBS 0.006802f
C446 B.n406 VSUBS 0.006802f
C447 B.n407 VSUBS 0.006802f
C448 B.n408 VSUBS 0.006802f
C449 B.n409 VSUBS 0.006802f
C450 B.n410 VSUBS 0.006802f
C451 B.n411 VSUBS 0.006802f
C452 B.n412 VSUBS 0.006802f
C453 B.n413 VSUBS 0.006802f
C454 B.n414 VSUBS 0.006802f
C455 B.n415 VSUBS 0.006802f
C456 B.n416 VSUBS 0.006802f
C457 B.n417 VSUBS 0.006802f
C458 B.n418 VSUBS 0.006802f
C459 B.n419 VSUBS 0.006802f
C460 B.n420 VSUBS 0.006802f
C461 B.n421 VSUBS 0.006802f
C462 B.n422 VSUBS 0.006802f
C463 B.n423 VSUBS 0.006802f
C464 B.n424 VSUBS 0.006802f
C465 B.n425 VSUBS 0.006802f
C466 B.n426 VSUBS 0.006802f
C467 B.n427 VSUBS 0.006802f
C468 B.n428 VSUBS 0.006802f
C469 B.n429 VSUBS 0.006802f
C470 B.n430 VSUBS 0.006802f
C471 B.n431 VSUBS 0.006802f
C472 B.n432 VSUBS 0.006802f
C473 B.n433 VSUBS 0.006802f
C474 B.n434 VSUBS 0.006802f
C475 B.n435 VSUBS 0.006802f
C476 B.n436 VSUBS 0.006802f
C477 B.n437 VSUBS 0.006802f
C478 B.n438 VSUBS 0.006802f
C479 B.n439 VSUBS 0.006802f
C480 B.n440 VSUBS 0.006802f
C481 B.n441 VSUBS 0.006802f
C482 B.n442 VSUBS 0.015659f
C483 B.n443 VSUBS 0.016463f
C484 B.n444 VSUBS 0.015345f
C485 B.n445 VSUBS 0.006802f
C486 B.n446 VSUBS 0.006802f
C487 B.n447 VSUBS 0.006802f
C488 B.n448 VSUBS 0.006802f
C489 B.n449 VSUBS 0.006802f
C490 B.n450 VSUBS 0.006802f
C491 B.n451 VSUBS 0.006802f
C492 B.n452 VSUBS 0.006802f
C493 B.n453 VSUBS 0.006802f
C494 B.n454 VSUBS 0.006802f
C495 B.n455 VSUBS 0.006802f
C496 B.n456 VSUBS 0.006802f
C497 B.n457 VSUBS 0.006802f
C498 B.n458 VSUBS 0.006802f
C499 B.n459 VSUBS 0.006802f
C500 B.n460 VSUBS 0.006802f
C501 B.n461 VSUBS 0.006802f
C502 B.n462 VSUBS 0.006802f
C503 B.n463 VSUBS 0.006802f
C504 B.n464 VSUBS 0.006802f
C505 B.n465 VSUBS 0.006802f
C506 B.n466 VSUBS 0.006802f
C507 B.n467 VSUBS 0.006802f
C508 B.n468 VSUBS 0.006802f
C509 B.n469 VSUBS 0.006802f
C510 B.n470 VSUBS 0.006802f
C511 B.n471 VSUBS 0.006802f
C512 B.n472 VSUBS 0.006802f
C513 B.n473 VSUBS 0.006802f
C514 B.n474 VSUBS 0.006802f
C515 B.n475 VSUBS 0.006802f
C516 B.n476 VSUBS 0.006802f
C517 B.n477 VSUBS 0.006802f
C518 B.n478 VSUBS 0.006802f
C519 B.n479 VSUBS 0.006802f
C520 B.n480 VSUBS 0.006802f
C521 B.n481 VSUBS 0.006802f
C522 B.n482 VSUBS 0.006802f
C523 B.n483 VSUBS 0.006802f
C524 B.n484 VSUBS 0.006802f
C525 B.n485 VSUBS 0.006802f
C526 B.n486 VSUBS 0.006802f
C527 B.n487 VSUBS 0.006802f
C528 B.n488 VSUBS 0.006802f
C529 B.n489 VSUBS 0.006802f
C530 B.n490 VSUBS 0.006802f
C531 B.n491 VSUBS 0.006802f
C532 B.n492 VSUBS 0.006802f
C533 B.n493 VSUBS 0.006802f
C534 B.n494 VSUBS 0.006802f
C535 B.n495 VSUBS 0.006802f
C536 B.n496 VSUBS 0.006802f
C537 B.n497 VSUBS 0.006802f
C538 B.n498 VSUBS 0.006802f
C539 B.n499 VSUBS 0.006802f
C540 B.n500 VSUBS 0.006802f
C541 B.n501 VSUBS 0.006802f
C542 B.n502 VSUBS 0.006802f
C543 B.n503 VSUBS 0.006802f
C544 B.n504 VSUBS 0.006802f
C545 B.n505 VSUBS 0.006802f
C546 B.n506 VSUBS 0.006802f
C547 B.n507 VSUBS 0.006802f
C548 B.n508 VSUBS 0.006802f
C549 B.n509 VSUBS 0.006802f
C550 B.n510 VSUBS 0.006802f
C551 B.n511 VSUBS 0.006802f
C552 B.n512 VSUBS 0.006802f
C553 B.n513 VSUBS 0.006802f
C554 B.n514 VSUBS 0.006802f
C555 B.n515 VSUBS 0.006802f
C556 B.n516 VSUBS 0.006802f
C557 B.n517 VSUBS 0.015345f
C558 B.n518 VSUBS 0.015345f
C559 B.n519 VSUBS 0.016463f
C560 B.n520 VSUBS 0.006802f
C561 B.n521 VSUBS 0.006802f
C562 B.n522 VSUBS 0.006802f
C563 B.n523 VSUBS 0.006802f
C564 B.n524 VSUBS 0.006802f
C565 B.n525 VSUBS 0.006802f
C566 B.n526 VSUBS 0.006802f
C567 B.n527 VSUBS 0.006802f
C568 B.n528 VSUBS 0.006802f
C569 B.n529 VSUBS 0.006802f
C570 B.n530 VSUBS 0.006802f
C571 B.n531 VSUBS 0.006802f
C572 B.n532 VSUBS 0.006802f
C573 B.n533 VSUBS 0.006802f
C574 B.n534 VSUBS 0.006802f
C575 B.n535 VSUBS 0.006802f
C576 B.n536 VSUBS 0.006802f
C577 B.n537 VSUBS 0.006802f
C578 B.n538 VSUBS 0.006802f
C579 B.n539 VSUBS 0.006802f
C580 B.n540 VSUBS 0.006802f
C581 B.n541 VSUBS 0.006802f
C582 B.n542 VSUBS 0.006802f
C583 B.n543 VSUBS 0.006802f
C584 B.n544 VSUBS 0.006802f
C585 B.n545 VSUBS 0.006802f
C586 B.n546 VSUBS 0.006802f
C587 B.n547 VSUBS 0.006802f
C588 B.n548 VSUBS 0.006802f
C589 B.n549 VSUBS 0.006802f
C590 B.n550 VSUBS 0.006802f
C591 B.n551 VSUBS 0.006802f
C592 B.n552 VSUBS 0.006802f
C593 B.n553 VSUBS 0.006802f
C594 B.n554 VSUBS 0.006802f
C595 B.n555 VSUBS 0.006802f
C596 B.n556 VSUBS 0.006802f
C597 B.n557 VSUBS 0.006802f
C598 B.n558 VSUBS 0.006802f
C599 B.n559 VSUBS 0.006802f
C600 B.n560 VSUBS 0.006802f
C601 B.n561 VSUBS 0.006802f
C602 B.n562 VSUBS 0.006802f
C603 B.n563 VSUBS 0.006802f
C604 B.n564 VSUBS 0.006802f
C605 B.n565 VSUBS 0.006802f
C606 B.n566 VSUBS 0.006802f
C607 B.n567 VSUBS 0.006802f
C608 B.n568 VSUBS 0.006802f
C609 B.n569 VSUBS 0.006802f
C610 B.n570 VSUBS 0.006802f
C611 B.n571 VSUBS 0.006802f
C612 B.n572 VSUBS 0.006802f
C613 B.n573 VSUBS 0.006802f
C614 B.n574 VSUBS 0.006802f
C615 B.n575 VSUBS 0.006802f
C616 B.n576 VSUBS 0.006802f
C617 B.n577 VSUBS 0.006802f
C618 B.n578 VSUBS 0.006802f
C619 B.n579 VSUBS 0.006802f
C620 B.n580 VSUBS 0.006802f
C621 B.n581 VSUBS 0.006802f
C622 B.n582 VSUBS 0.006802f
C623 B.n583 VSUBS 0.006802f
C624 B.n584 VSUBS 0.006802f
C625 B.n585 VSUBS 0.006802f
C626 B.n586 VSUBS 0.006802f
C627 B.n587 VSUBS 0.006802f
C628 B.n588 VSUBS 0.006802f
C629 B.n589 VSUBS 0.006802f
C630 B.n590 VSUBS 0.006802f
C631 B.n591 VSUBS 0.006802f
C632 B.n592 VSUBS 0.006802f
C633 B.n593 VSUBS 0.006802f
C634 B.n594 VSUBS 0.006802f
C635 B.n595 VSUBS 0.006802f
C636 B.n596 VSUBS 0.006802f
C637 B.n597 VSUBS 0.006802f
C638 B.n598 VSUBS 0.006802f
C639 B.n599 VSUBS 0.006802f
C640 B.n600 VSUBS 0.006802f
C641 B.n601 VSUBS 0.006802f
C642 B.n602 VSUBS 0.006802f
C643 B.n603 VSUBS 0.006802f
C644 B.n604 VSUBS 0.006802f
C645 B.n605 VSUBS 0.006802f
C646 B.n606 VSUBS 0.006802f
C647 B.n607 VSUBS 0.006802f
C648 B.n608 VSUBS 0.006802f
C649 B.n609 VSUBS 0.006802f
C650 B.n610 VSUBS 0.006802f
C651 B.n611 VSUBS 0.006802f
C652 B.n612 VSUBS 0.006802f
C653 B.n613 VSUBS 0.006802f
C654 B.n614 VSUBS 0.006802f
C655 B.n615 VSUBS 0.004701f
C656 B.n616 VSUBS 0.015759f
C657 B.n617 VSUBS 0.005501f
C658 B.n618 VSUBS 0.006802f
C659 B.n619 VSUBS 0.006802f
C660 B.n620 VSUBS 0.006802f
C661 B.n621 VSUBS 0.006802f
C662 B.n622 VSUBS 0.006802f
C663 B.n623 VSUBS 0.006802f
C664 B.n624 VSUBS 0.006802f
C665 B.n625 VSUBS 0.006802f
C666 B.n626 VSUBS 0.006802f
C667 B.n627 VSUBS 0.006802f
C668 B.n628 VSUBS 0.006802f
C669 B.n629 VSUBS 0.005501f
C670 B.n630 VSUBS 0.006802f
C671 B.n631 VSUBS 0.006802f
C672 B.n632 VSUBS 0.006802f
C673 B.n633 VSUBS 0.006802f
C674 B.n634 VSUBS 0.006802f
C675 B.n635 VSUBS 0.006802f
C676 B.n636 VSUBS 0.006802f
C677 B.n637 VSUBS 0.006802f
C678 B.n638 VSUBS 0.006802f
C679 B.n639 VSUBS 0.006802f
C680 B.n640 VSUBS 0.006802f
C681 B.n641 VSUBS 0.006802f
C682 B.n642 VSUBS 0.006802f
C683 B.n643 VSUBS 0.006802f
C684 B.n644 VSUBS 0.006802f
C685 B.n645 VSUBS 0.006802f
C686 B.n646 VSUBS 0.006802f
C687 B.n647 VSUBS 0.006802f
C688 B.n648 VSUBS 0.006802f
C689 B.n649 VSUBS 0.006802f
C690 B.n650 VSUBS 0.006802f
C691 B.n651 VSUBS 0.006802f
C692 B.n652 VSUBS 0.006802f
C693 B.n653 VSUBS 0.006802f
C694 B.n654 VSUBS 0.006802f
C695 B.n655 VSUBS 0.006802f
C696 B.n656 VSUBS 0.006802f
C697 B.n657 VSUBS 0.006802f
C698 B.n658 VSUBS 0.006802f
C699 B.n659 VSUBS 0.006802f
C700 B.n660 VSUBS 0.006802f
C701 B.n661 VSUBS 0.006802f
C702 B.n662 VSUBS 0.006802f
C703 B.n663 VSUBS 0.006802f
C704 B.n664 VSUBS 0.006802f
C705 B.n665 VSUBS 0.006802f
C706 B.n666 VSUBS 0.006802f
C707 B.n667 VSUBS 0.006802f
C708 B.n668 VSUBS 0.006802f
C709 B.n669 VSUBS 0.006802f
C710 B.n670 VSUBS 0.006802f
C711 B.n671 VSUBS 0.006802f
C712 B.n672 VSUBS 0.006802f
C713 B.n673 VSUBS 0.006802f
C714 B.n674 VSUBS 0.006802f
C715 B.n675 VSUBS 0.006802f
C716 B.n676 VSUBS 0.006802f
C717 B.n677 VSUBS 0.006802f
C718 B.n678 VSUBS 0.006802f
C719 B.n679 VSUBS 0.006802f
C720 B.n680 VSUBS 0.006802f
C721 B.n681 VSUBS 0.006802f
C722 B.n682 VSUBS 0.006802f
C723 B.n683 VSUBS 0.006802f
C724 B.n684 VSUBS 0.006802f
C725 B.n685 VSUBS 0.006802f
C726 B.n686 VSUBS 0.006802f
C727 B.n687 VSUBS 0.006802f
C728 B.n688 VSUBS 0.006802f
C729 B.n689 VSUBS 0.006802f
C730 B.n690 VSUBS 0.006802f
C731 B.n691 VSUBS 0.006802f
C732 B.n692 VSUBS 0.006802f
C733 B.n693 VSUBS 0.006802f
C734 B.n694 VSUBS 0.006802f
C735 B.n695 VSUBS 0.006802f
C736 B.n696 VSUBS 0.006802f
C737 B.n697 VSUBS 0.006802f
C738 B.n698 VSUBS 0.006802f
C739 B.n699 VSUBS 0.006802f
C740 B.n700 VSUBS 0.006802f
C741 B.n701 VSUBS 0.006802f
C742 B.n702 VSUBS 0.006802f
C743 B.n703 VSUBS 0.006802f
C744 B.n704 VSUBS 0.006802f
C745 B.n705 VSUBS 0.006802f
C746 B.n706 VSUBS 0.006802f
C747 B.n707 VSUBS 0.006802f
C748 B.n708 VSUBS 0.006802f
C749 B.n709 VSUBS 0.006802f
C750 B.n710 VSUBS 0.006802f
C751 B.n711 VSUBS 0.006802f
C752 B.n712 VSUBS 0.006802f
C753 B.n713 VSUBS 0.006802f
C754 B.n714 VSUBS 0.006802f
C755 B.n715 VSUBS 0.006802f
C756 B.n716 VSUBS 0.006802f
C757 B.n717 VSUBS 0.006802f
C758 B.n718 VSUBS 0.006802f
C759 B.n719 VSUBS 0.006802f
C760 B.n720 VSUBS 0.006802f
C761 B.n721 VSUBS 0.006802f
C762 B.n722 VSUBS 0.006802f
C763 B.n723 VSUBS 0.006802f
C764 B.n724 VSUBS 0.006802f
C765 B.n725 VSUBS 0.006802f
C766 B.n726 VSUBS 0.006802f
C767 B.n727 VSUBS 0.016463f
C768 B.n728 VSUBS 0.015345f
C769 B.n729 VSUBS 0.015345f
C770 B.n730 VSUBS 0.006802f
C771 B.n731 VSUBS 0.006802f
C772 B.n732 VSUBS 0.006802f
C773 B.n733 VSUBS 0.006802f
C774 B.n734 VSUBS 0.006802f
C775 B.n735 VSUBS 0.006802f
C776 B.n736 VSUBS 0.006802f
C777 B.n737 VSUBS 0.006802f
C778 B.n738 VSUBS 0.006802f
C779 B.n739 VSUBS 0.006802f
C780 B.n740 VSUBS 0.006802f
C781 B.n741 VSUBS 0.006802f
C782 B.n742 VSUBS 0.006802f
C783 B.n743 VSUBS 0.006802f
C784 B.n744 VSUBS 0.006802f
C785 B.n745 VSUBS 0.006802f
C786 B.n746 VSUBS 0.006802f
C787 B.n747 VSUBS 0.006802f
C788 B.n748 VSUBS 0.006802f
C789 B.n749 VSUBS 0.006802f
C790 B.n750 VSUBS 0.006802f
C791 B.n751 VSUBS 0.006802f
C792 B.n752 VSUBS 0.006802f
C793 B.n753 VSUBS 0.006802f
C794 B.n754 VSUBS 0.006802f
C795 B.n755 VSUBS 0.006802f
C796 B.n756 VSUBS 0.006802f
C797 B.n757 VSUBS 0.006802f
C798 B.n758 VSUBS 0.006802f
C799 B.n759 VSUBS 0.006802f
C800 B.n760 VSUBS 0.006802f
C801 B.n761 VSUBS 0.006802f
C802 B.n762 VSUBS 0.006802f
C803 B.n763 VSUBS 0.008876f
C804 B.n764 VSUBS 0.009455f
C805 B.n765 VSUBS 0.018802f
C806 VDD1.t1 VSUBS 4.7676f
C807 VDD1.t0 VSUBS 5.9088f
C808 VP.t0 VSUBS 6.07274f
C809 VP.t1 VSUBS 5.4252f
C810 VP.n0 VSUBS 6.81723f
C811 VDD2.t1 VSUBS 5.85604f
C812 VDD2.t0 VSUBS 4.76192f
C813 VDD2.n0 VSUBS 5.41334f
C814 VTAIL.t3 VSUBS 4.56087f
C815 VTAIL.n0 VSUBS 3.22344f
C816 VTAIL.t1 VSUBS 4.56087f
C817 VTAIL.n1 VSUBS 3.27236f
C818 VTAIL.t0 VSUBS 4.56087f
C819 VTAIL.n2 VSUBS 3.0559f
C820 VTAIL.t2 VSUBS 4.56087f
C821 VTAIL.n3 VSUBS 2.95461f
C822 VN.t0 VSUBS 5.26519f
C823 VN.t1 VSUBS 5.89406f
.ends

