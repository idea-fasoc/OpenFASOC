* NGSPICE file created from diff_pair_sample_0299.ext - technology: sky130A

.subckt diff_pair_sample_0299 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0.49005 ps=3.3 w=2.97 l=2.27
X1 VDD2.t9 VN.t0 VTAIL.t19 B.t6 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0 ps=0 w=2.97 l=2.27
X3 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0 ps=0 w=2.97 l=2.27
X4 VDD1.t8 VP.t1 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=1.1583 ps=6.72 w=2.97 l=2.27
X5 VTAIL.t8 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X6 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0 ps=0 w=2.97 l=2.27
X7 VTAIL.t12 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X8 VTAIL.t1 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X9 VDD1.t5 VP.t4 VTAIL.t10 B.t8 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X10 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=1.1583 ps=6.72 w=2.97 l=2.27
X11 VTAIL.t18 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X12 VDD1.t4 VP.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=1.1583 ps=6.72 w=2.97 l=2.27
X13 VTAIL.t14 VP.t6 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X14 VDD2.t5 VN.t4 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X15 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0.49005 ps=3.3 w=2.97 l=2.27
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0 ps=0 w=2.97 l=2.27
X17 VDD1.t2 VP.t7 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0.49005 ps=3.3 w=2.97 l=2.27
X18 VDD2.t3 VN.t6 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=1.1583 ps=6.72 w=2.97 l=2.27
X19 VDD1.t1 VP.t8 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X20 VTAIL.t7 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X21 VTAIL.t17 VN.t7 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X22 VTAIL.t15 VN.t8 VDD2.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.49005 pd=3.3 as=0.49005 ps=3.3 w=2.97 l=2.27
X23 VDD2.t0 VN.t9 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1583 pd=6.72 as=0.49005 ps=3.3 w=2.97 l=2.27
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n16 161.3
R6 VP.n31 VP.n30 161.3
R7 VP.n32 VP.n15 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n14 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n39 VP.n13 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n42 VP.n12 161.3
R14 VP.n44 VP.n43 161.3
R15 VP.n45 VP.n11 161.3
R16 VP.n82 VP.n0 161.3
R17 VP.n81 VP.n80 161.3
R18 VP.n79 VP.n1 161.3
R19 VP.n78 VP.n77 161.3
R20 VP.n76 VP.n2 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n3 161.3
R23 VP.n71 VP.n70 161.3
R24 VP.n69 VP.n4 161.3
R25 VP.n68 VP.n67 161.3
R26 VP.n66 VP.n5 161.3
R27 VP.n65 VP.n64 161.3
R28 VP.n63 VP.n6 161.3
R29 VP.n62 VP.n61 161.3
R30 VP.n60 VP.n7 161.3
R31 VP.n59 VP.n58 161.3
R32 VP.n56 VP.n8 161.3
R33 VP.n55 VP.n54 161.3
R34 VP.n53 VP.n9 161.3
R35 VP.n52 VP.n51 161.3
R36 VP.n50 VP.n10 161.3
R37 VP.n49 VP.n48 100.969
R38 VP.n84 VP.n83 100.969
R39 VP.n47 VP.n46 100.969
R40 VP.n20 VP.n19 67.1934
R41 VP.n19 VP.t7 62.4054
R42 VP.n63 VP.n62 56.5193
R43 VP.n70 VP.n69 56.5193
R44 VP.n33 VP.n32 56.5193
R45 VP.n26 VP.n25 56.5193
R46 VP.n55 VP.n9 50.2061
R47 VP.n77 VP.n1 50.2061
R48 VP.n40 VP.n12 50.2061
R49 VP.n48 VP.n47 44.4163
R50 VP.n5 VP.t4 31.5322
R51 VP.n49 VP.t0 31.5322
R52 VP.n57 VP.t3 31.5322
R53 VP.n75 VP.t2 31.5322
R54 VP.n83 VP.t1 31.5322
R55 VP.n16 VP.t8 31.5322
R56 VP.n46 VP.t5 31.5322
R57 VP.n38 VP.t6 31.5322
R58 VP.n20 VP.t9 31.5322
R59 VP.n51 VP.n9 30.7807
R60 VP.n81 VP.n1 30.7807
R61 VP.n44 VP.n12 30.7807
R62 VP.n51 VP.n50 24.4675
R63 VP.n56 VP.n55 24.4675
R64 VP.n58 VP.n7 24.4675
R65 VP.n62 VP.n7 24.4675
R66 VP.n64 VP.n63 24.4675
R67 VP.n64 VP.n5 24.4675
R68 VP.n68 VP.n5 24.4675
R69 VP.n69 VP.n68 24.4675
R70 VP.n70 VP.n3 24.4675
R71 VP.n74 VP.n3 24.4675
R72 VP.n77 VP.n76 24.4675
R73 VP.n82 VP.n81 24.4675
R74 VP.n45 VP.n44 24.4675
R75 VP.n33 VP.n14 24.4675
R76 VP.n37 VP.n14 24.4675
R77 VP.n40 VP.n39 24.4675
R78 VP.n27 VP.n26 24.4675
R79 VP.n27 VP.n16 24.4675
R80 VP.n31 VP.n16 24.4675
R81 VP.n32 VP.n31 24.4675
R82 VP.n21 VP.n18 24.4675
R83 VP.n25 VP.n18 24.4675
R84 VP.n57 VP.n56 19.5741
R85 VP.n76 VP.n75 19.5741
R86 VP.n39 VP.n38 19.5741
R87 VP.n22 VP.n19 10.026
R88 VP.n50 VP.n49 9.7873
R89 VP.n83 VP.n82 9.7873
R90 VP.n46 VP.n45 9.7873
R91 VP.n58 VP.n57 4.8939
R92 VP.n75 VP.n74 4.8939
R93 VP.n38 VP.n37 4.8939
R94 VP.n21 VP.n20 4.8939
R95 VP.n47 VP.n11 0.278367
R96 VP.n48 VP.n10 0.278367
R97 VP.n84 VP.n0 0.278367
R98 VP.n23 VP.n22 0.189894
R99 VP.n24 VP.n23 0.189894
R100 VP.n24 VP.n17 0.189894
R101 VP.n28 VP.n17 0.189894
R102 VP.n29 VP.n28 0.189894
R103 VP.n30 VP.n29 0.189894
R104 VP.n30 VP.n15 0.189894
R105 VP.n34 VP.n15 0.189894
R106 VP.n35 VP.n34 0.189894
R107 VP.n36 VP.n35 0.189894
R108 VP.n36 VP.n13 0.189894
R109 VP.n41 VP.n13 0.189894
R110 VP.n42 VP.n41 0.189894
R111 VP.n43 VP.n42 0.189894
R112 VP.n43 VP.n11 0.189894
R113 VP.n52 VP.n10 0.189894
R114 VP.n53 VP.n52 0.189894
R115 VP.n54 VP.n53 0.189894
R116 VP.n54 VP.n8 0.189894
R117 VP.n59 VP.n8 0.189894
R118 VP.n60 VP.n59 0.189894
R119 VP.n61 VP.n60 0.189894
R120 VP.n61 VP.n6 0.189894
R121 VP.n65 VP.n6 0.189894
R122 VP.n66 VP.n65 0.189894
R123 VP.n67 VP.n66 0.189894
R124 VP.n67 VP.n4 0.189894
R125 VP.n71 VP.n4 0.189894
R126 VP.n72 VP.n71 0.189894
R127 VP.n73 VP.n72 0.189894
R128 VP.n73 VP.n2 0.189894
R129 VP.n78 VP.n2 0.189894
R130 VP.n79 VP.n78 0.189894
R131 VP.n80 VP.n79 0.189894
R132 VP.n80 VP.n0 0.189894
R133 VP VP.n84 0.153454
R134 VTAIL.n11 VTAIL.t4 74.8892
R135 VTAIL.n17 VTAIL.t3 74.889
R136 VTAIL.n2 VTAIL.t9 74.889
R137 VTAIL.n16 VTAIL.t6 74.889
R138 VTAIL.n15 VTAIL.n14 68.2225
R139 VTAIL.n13 VTAIL.n12 68.2225
R140 VTAIL.n10 VTAIL.n9 68.2225
R141 VTAIL.n8 VTAIL.n7 68.2225
R142 VTAIL.n19 VTAIL.n18 68.2223
R143 VTAIL.n1 VTAIL.n0 68.2223
R144 VTAIL.n4 VTAIL.n3 68.2223
R145 VTAIL.n6 VTAIL.n5 68.2223
R146 VTAIL.n8 VTAIL.n6 19.41
R147 VTAIL.n17 VTAIL.n16 17.1686
R148 VTAIL.n18 VTAIL.t19 6.66717
R149 VTAIL.n18 VTAIL.t18 6.66717
R150 VTAIL.n0 VTAIL.t2 6.66717
R151 VTAIL.n0 VTAIL.t17 6.66717
R152 VTAIL.n3 VTAIL.t10 6.66717
R153 VTAIL.n3 VTAIL.t8 6.66717
R154 VTAIL.n5 VTAIL.t13 6.66717
R155 VTAIL.n5 VTAIL.t12 6.66717
R156 VTAIL.n14 VTAIL.t11 6.66717
R157 VTAIL.n14 VTAIL.t14 6.66717
R158 VTAIL.n12 VTAIL.t5 6.66717
R159 VTAIL.n12 VTAIL.t7 6.66717
R160 VTAIL.n9 VTAIL.t16 6.66717
R161 VTAIL.n9 VTAIL.t1 6.66717
R162 VTAIL.n7 VTAIL.t0 6.66717
R163 VTAIL.n7 VTAIL.t15 6.66717
R164 VTAIL.n10 VTAIL.n8 2.24188
R165 VTAIL.n11 VTAIL.n10 2.24188
R166 VTAIL.n15 VTAIL.n13 2.24188
R167 VTAIL.n16 VTAIL.n15 2.24188
R168 VTAIL.n6 VTAIL.n4 2.24188
R169 VTAIL.n4 VTAIL.n2 2.24188
R170 VTAIL.n19 VTAIL.n17 2.24188
R171 VTAIL VTAIL.n1 1.73972
R172 VTAIL.n13 VTAIL.n11 1.59102
R173 VTAIL.n2 VTAIL.n1 1.59102
R174 VTAIL VTAIL.n19 0.502655
R175 VDD1.n1 VDD1.t2 93.8094
R176 VDD1.n3 VDD1.t9 93.8091
R177 VDD1.n5 VDD1.n4 86.5268
R178 VDD1.n1 VDD1.n0 84.9013
R179 VDD1.n7 VDD1.n6 84.9012
R180 VDD1.n3 VDD1.n2 84.9011
R181 VDD1.n7 VDD1.n5 38.6259
R182 VDD1.n6 VDD1.t3 6.66717
R183 VDD1.n6 VDD1.t4 6.66717
R184 VDD1.n0 VDD1.t0 6.66717
R185 VDD1.n0 VDD1.t1 6.66717
R186 VDD1.n4 VDD1.t7 6.66717
R187 VDD1.n4 VDD1.t8 6.66717
R188 VDD1.n2 VDD1.t6 6.66717
R189 VDD1.n2 VDD1.t5 6.66717
R190 VDD1 VDD1.n7 1.62334
R191 VDD1 VDD1.n1 0.619035
R192 VDD1.n5 VDD1.n3 0.505499
R193 B.n567 B.n566 585
R194 B.n569 B.n124 585
R195 B.n572 B.n571 585
R196 B.n573 B.n123 585
R197 B.n575 B.n574 585
R198 B.n577 B.n122 585
R199 B.n580 B.n579 585
R200 B.n581 B.n121 585
R201 B.n583 B.n582 585
R202 B.n585 B.n120 585
R203 B.n588 B.n587 585
R204 B.n589 B.n119 585
R205 B.n591 B.n590 585
R206 B.n593 B.n118 585
R207 B.n596 B.n595 585
R208 B.n598 B.n115 585
R209 B.n600 B.n599 585
R210 B.n602 B.n114 585
R211 B.n605 B.n604 585
R212 B.n606 B.n113 585
R213 B.n608 B.n607 585
R214 B.n610 B.n112 585
R215 B.n613 B.n612 585
R216 B.n614 B.n108 585
R217 B.n616 B.n615 585
R218 B.n618 B.n107 585
R219 B.n621 B.n620 585
R220 B.n622 B.n106 585
R221 B.n624 B.n623 585
R222 B.n626 B.n105 585
R223 B.n629 B.n628 585
R224 B.n630 B.n104 585
R225 B.n632 B.n631 585
R226 B.n634 B.n103 585
R227 B.n637 B.n636 585
R228 B.n638 B.n102 585
R229 B.n640 B.n639 585
R230 B.n642 B.n101 585
R231 B.n645 B.n644 585
R232 B.n646 B.n100 585
R233 B.n565 B.n98 585
R234 B.n649 B.n98 585
R235 B.n564 B.n97 585
R236 B.n650 B.n97 585
R237 B.n563 B.n96 585
R238 B.n651 B.n96 585
R239 B.n562 B.n561 585
R240 B.n561 B.n92 585
R241 B.n560 B.n91 585
R242 B.n657 B.n91 585
R243 B.n559 B.n90 585
R244 B.n658 B.n90 585
R245 B.n558 B.n89 585
R246 B.n659 B.n89 585
R247 B.n557 B.n556 585
R248 B.n556 B.n88 585
R249 B.n555 B.n84 585
R250 B.n665 B.n84 585
R251 B.n554 B.n83 585
R252 B.n666 B.n83 585
R253 B.n553 B.n82 585
R254 B.n667 B.n82 585
R255 B.n552 B.n551 585
R256 B.n551 B.n78 585
R257 B.n550 B.n77 585
R258 B.n673 B.n77 585
R259 B.n549 B.n76 585
R260 B.n674 B.n76 585
R261 B.n548 B.n75 585
R262 B.n675 B.n75 585
R263 B.n547 B.n546 585
R264 B.n546 B.n71 585
R265 B.n545 B.n70 585
R266 B.n681 B.n70 585
R267 B.n544 B.n69 585
R268 B.n682 B.n69 585
R269 B.n543 B.n68 585
R270 B.n683 B.n68 585
R271 B.n542 B.n541 585
R272 B.n541 B.n64 585
R273 B.n540 B.n63 585
R274 B.n689 B.n63 585
R275 B.n539 B.n62 585
R276 B.n690 B.n62 585
R277 B.n538 B.n61 585
R278 B.n691 B.n61 585
R279 B.n537 B.n536 585
R280 B.n536 B.n57 585
R281 B.n535 B.n56 585
R282 B.n697 B.n56 585
R283 B.n534 B.n55 585
R284 B.n698 B.n55 585
R285 B.n533 B.n54 585
R286 B.n699 B.n54 585
R287 B.n532 B.n531 585
R288 B.n531 B.n50 585
R289 B.n530 B.n49 585
R290 B.n705 B.n49 585
R291 B.n529 B.n48 585
R292 B.n706 B.n48 585
R293 B.n528 B.n47 585
R294 B.n707 B.n47 585
R295 B.n527 B.n526 585
R296 B.n526 B.n43 585
R297 B.n525 B.n42 585
R298 B.n713 B.n42 585
R299 B.n524 B.n41 585
R300 B.n714 B.n41 585
R301 B.n523 B.n40 585
R302 B.n715 B.n40 585
R303 B.n522 B.n521 585
R304 B.n521 B.n36 585
R305 B.n520 B.n35 585
R306 B.n721 B.n35 585
R307 B.n519 B.n34 585
R308 B.n722 B.n34 585
R309 B.n518 B.n33 585
R310 B.n723 B.n33 585
R311 B.n517 B.n516 585
R312 B.n516 B.n29 585
R313 B.n515 B.n28 585
R314 B.n729 B.n28 585
R315 B.n514 B.n27 585
R316 B.n730 B.n27 585
R317 B.n513 B.n26 585
R318 B.n731 B.n26 585
R319 B.n512 B.n511 585
R320 B.n511 B.n22 585
R321 B.n510 B.n21 585
R322 B.n737 B.n21 585
R323 B.n509 B.n20 585
R324 B.n738 B.n20 585
R325 B.n508 B.n19 585
R326 B.n739 B.n19 585
R327 B.n507 B.n506 585
R328 B.n506 B.n15 585
R329 B.n505 B.n14 585
R330 B.n745 B.n14 585
R331 B.n504 B.n13 585
R332 B.n746 B.n13 585
R333 B.n503 B.n12 585
R334 B.n747 B.n12 585
R335 B.n502 B.n501 585
R336 B.n501 B.n8 585
R337 B.n500 B.n7 585
R338 B.n753 B.n7 585
R339 B.n499 B.n6 585
R340 B.n754 B.n6 585
R341 B.n498 B.n5 585
R342 B.n755 B.n5 585
R343 B.n497 B.n496 585
R344 B.n496 B.n4 585
R345 B.n495 B.n125 585
R346 B.n495 B.n494 585
R347 B.n485 B.n126 585
R348 B.n127 B.n126 585
R349 B.n487 B.n486 585
R350 B.n488 B.n487 585
R351 B.n484 B.n132 585
R352 B.n132 B.n131 585
R353 B.n483 B.n482 585
R354 B.n482 B.n481 585
R355 B.n134 B.n133 585
R356 B.n135 B.n134 585
R357 B.n474 B.n473 585
R358 B.n475 B.n474 585
R359 B.n472 B.n140 585
R360 B.n140 B.n139 585
R361 B.n471 B.n470 585
R362 B.n470 B.n469 585
R363 B.n142 B.n141 585
R364 B.n143 B.n142 585
R365 B.n462 B.n461 585
R366 B.n463 B.n462 585
R367 B.n460 B.n148 585
R368 B.n148 B.n147 585
R369 B.n459 B.n458 585
R370 B.n458 B.n457 585
R371 B.n150 B.n149 585
R372 B.n151 B.n150 585
R373 B.n450 B.n449 585
R374 B.n451 B.n450 585
R375 B.n448 B.n156 585
R376 B.n156 B.n155 585
R377 B.n447 B.n446 585
R378 B.n446 B.n445 585
R379 B.n158 B.n157 585
R380 B.n159 B.n158 585
R381 B.n438 B.n437 585
R382 B.n439 B.n438 585
R383 B.n436 B.n163 585
R384 B.n167 B.n163 585
R385 B.n435 B.n434 585
R386 B.n434 B.n433 585
R387 B.n165 B.n164 585
R388 B.n166 B.n165 585
R389 B.n426 B.n425 585
R390 B.n427 B.n426 585
R391 B.n424 B.n172 585
R392 B.n172 B.n171 585
R393 B.n423 B.n422 585
R394 B.n422 B.n421 585
R395 B.n174 B.n173 585
R396 B.n175 B.n174 585
R397 B.n414 B.n413 585
R398 B.n415 B.n414 585
R399 B.n412 B.n179 585
R400 B.n183 B.n179 585
R401 B.n411 B.n410 585
R402 B.n410 B.n409 585
R403 B.n181 B.n180 585
R404 B.n182 B.n181 585
R405 B.n402 B.n401 585
R406 B.n403 B.n402 585
R407 B.n400 B.n188 585
R408 B.n188 B.n187 585
R409 B.n399 B.n398 585
R410 B.n398 B.n397 585
R411 B.n190 B.n189 585
R412 B.n191 B.n190 585
R413 B.n390 B.n389 585
R414 B.n391 B.n390 585
R415 B.n388 B.n195 585
R416 B.n199 B.n195 585
R417 B.n387 B.n386 585
R418 B.n386 B.n385 585
R419 B.n197 B.n196 585
R420 B.n198 B.n197 585
R421 B.n378 B.n377 585
R422 B.n379 B.n378 585
R423 B.n376 B.n204 585
R424 B.n204 B.n203 585
R425 B.n375 B.n374 585
R426 B.n374 B.n373 585
R427 B.n206 B.n205 585
R428 B.n207 B.n206 585
R429 B.n366 B.n365 585
R430 B.n367 B.n366 585
R431 B.n364 B.n212 585
R432 B.n212 B.n211 585
R433 B.n363 B.n362 585
R434 B.n362 B.n361 585
R435 B.n214 B.n213 585
R436 B.n354 B.n214 585
R437 B.n353 B.n352 585
R438 B.n355 B.n353 585
R439 B.n351 B.n219 585
R440 B.n219 B.n218 585
R441 B.n350 B.n349 585
R442 B.n349 B.n348 585
R443 B.n221 B.n220 585
R444 B.n222 B.n221 585
R445 B.n341 B.n340 585
R446 B.n342 B.n341 585
R447 B.n339 B.n227 585
R448 B.n227 B.n226 585
R449 B.n338 B.n337 585
R450 B.n337 B.n336 585
R451 B.n333 B.n231 585
R452 B.n332 B.n331 585
R453 B.n329 B.n232 585
R454 B.n329 B.n230 585
R455 B.n328 B.n327 585
R456 B.n326 B.n325 585
R457 B.n324 B.n234 585
R458 B.n322 B.n321 585
R459 B.n320 B.n235 585
R460 B.n319 B.n318 585
R461 B.n316 B.n236 585
R462 B.n314 B.n313 585
R463 B.n312 B.n237 585
R464 B.n311 B.n310 585
R465 B.n308 B.n238 585
R466 B.n306 B.n305 585
R467 B.n303 B.n239 585
R468 B.n302 B.n301 585
R469 B.n299 B.n242 585
R470 B.n297 B.n296 585
R471 B.n295 B.n243 585
R472 B.n294 B.n293 585
R473 B.n291 B.n244 585
R474 B.n289 B.n288 585
R475 B.n287 B.n245 585
R476 B.n286 B.n285 585
R477 B.n283 B.n282 585
R478 B.n281 B.n280 585
R479 B.n279 B.n250 585
R480 B.n277 B.n276 585
R481 B.n275 B.n251 585
R482 B.n274 B.n273 585
R483 B.n271 B.n252 585
R484 B.n269 B.n268 585
R485 B.n267 B.n253 585
R486 B.n266 B.n265 585
R487 B.n263 B.n254 585
R488 B.n261 B.n260 585
R489 B.n259 B.n255 585
R490 B.n258 B.n257 585
R491 B.n229 B.n228 585
R492 B.n230 B.n229 585
R493 B.n335 B.n334 585
R494 B.n336 B.n335 585
R495 B.n225 B.n224 585
R496 B.n226 B.n225 585
R497 B.n344 B.n343 585
R498 B.n343 B.n342 585
R499 B.n345 B.n223 585
R500 B.n223 B.n222 585
R501 B.n347 B.n346 585
R502 B.n348 B.n347 585
R503 B.n217 B.n216 585
R504 B.n218 B.n217 585
R505 B.n357 B.n356 585
R506 B.n356 B.n355 585
R507 B.n358 B.n215 585
R508 B.n354 B.n215 585
R509 B.n360 B.n359 585
R510 B.n361 B.n360 585
R511 B.n210 B.n209 585
R512 B.n211 B.n210 585
R513 B.n369 B.n368 585
R514 B.n368 B.n367 585
R515 B.n370 B.n208 585
R516 B.n208 B.n207 585
R517 B.n372 B.n371 585
R518 B.n373 B.n372 585
R519 B.n202 B.n201 585
R520 B.n203 B.n202 585
R521 B.n381 B.n380 585
R522 B.n380 B.n379 585
R523 B.n382 B.n200 585
R524 B.n200 B.n198 585
R525 B.n384 B.n383 585
R526 B.n385 B.n384 585
R527 B.n194 B.n193 585
R528 B.n199 B.n194 585
R529 B.n393 B.n392 585
R530 B.n392 B.n391 585
R531 B.n394 B.n192 585
R532 B.n192 B.n191 585
R533 B.n396 B.n395 585
R534 B.n397 B.n396 585
R535 B.n186 B.n185 585
R536 B.n187 B.n186 585
R537 B.n405 B.n404 585
R538 B.n404 B.n403 585
R539 B.n406 B.n184 585
R540 B.n184 B.n182 585
R541 B.n408 B.n407 585
R542 B.n409 B.n408 585
R543 B.n178 B.n177 585
R544 B.n183 B.n178 585
R545 B.n417 B.n416 585
R546 B.n416 B.n415 585
R547 B.n418 B.n176 585
R548 B.n176 B.n175 585
R549 B.n420 B.n419 585
R550 B.n421 B.n420 585
R551 B.n170 B.n169 585
R552 B.n171 B.n170 585
R553 B.n429 B.n428 585
R554 B.n428 B.n427 585
R555 B.n430 B.n168 585
R556 B.n168 B.n166 585
R557 B.n432 B.n431 585
R558 B.n433 B.n432 585
R559 B.n162 B.n161 585
R560 B.n167 B.n162 585
R561 B.n441 B.n440 585
R562 B.n440 B.n439 585
R563 B.n442 B.n160 585
R564 B.n160 B.n159 585
R565 B.n444 B.n443 585
R566 B.n445 B.n444 585
R567 B.n154 B.n153 585
R568 B.n155 B.n154 585
R569 B.n453 B.n452 585
R570 B.n452 B.n451 585
R571 B.n454 B.n152 585
R572 B.n152 B.n151 585
R573 B.n456 B.n455 585
R574 B.n457 B.n456 585
R575 B.n146 B.n145 585
R576 B.n147 B.n146 585
R577 B.n465 B.n464 585
R578 B.n464 B.n463 585
R579 B.n466 B.n144 585
R580 B.n144 B.n143 585
R581 B.n468 B.n467 585
R582 B.n469 B.n468 585
R583 B.n138 B.n137 585
R584 B.n139 B.n138 585
R585 B.n477 B.n476 585
R586 B.n476 B.n475 585
R587 B.n478 B.n136 585
R588 B.n136 B.n135 585
R589 B.n480 B.n479 585
R590 B.n481 B.n480 585
R591 B.n130 B.n129 585
R592 B.n131 B.n130 585
R593 B.n490 B.n489 585
R594 B.n489 B.n488 585
R595 B.n491 B.n128 585
R596 B.n128 B.n127 585
R597 B.n493 B.n492 585
R598 B.n494 B.n493 585
R599 B.n2 B.n0 585
R600 B.n4 B.n2 585
R601 B.n3 B.n1 585
R602 B.n754 B.n3 585
R603 B.n752 B.n751 585
R604 B.n753 B.n752 585
R605 B.n750 B.n9 585
R606 B.n9 B.n8 585
R607 B.n749 B.n748 585
R608 B.n748 B.n747 585
R609 B.n11 B.n10 585
R610 B.n746 B.n11 585
R611 B.n744 B.n743 585
R612 B.n745 B.n744 585
R613 B.n742 B.n16 585
R614 B.n16 B.n15 585
R615 B.n741 B.n740 585
R616 B.n740 B.n739 585
R617 B.n18 B.n17 585
R618 B.n738 B.n18 585
R619 B.n736 B.n735 585
R620 B.n737 B.n736 585
R621 B.n734 B.n23 585
R622 B.n23 B.n22 585
R623 B.n733 B.n732 585
R624 B.n732 B.n731 585
R625 B.n25 B.n24 585
R626 B.n730 B.n25 585
R627 B.n728 B.n727 585
R628 B.n729 B.n728 585
R629 B.n726 B.n30 585
R630 B.n30 B.n29 585
R631 B.n725 B.n724 585
R632 B.n724 B.n723 585
R633 B.n32 B.n31 585
R634 B.n722 B.n32 585
R635 B.n720 B.n719 585
R636 B.n721 B.n720 585
R637 B.n718 B.n37 585
R638 B.n37 B.n36 585
R639 B.n717 B.n716 585
R640 B.n716 B.n715 585
R641 B.n39 B.n38 585
R642 B.n714 B.n39 585
R643 B.n712 B.n711 585
R644 B.n713 B.n712 585
R645 B.n710 B.n44 585
R646 B.n44 B.n43 585
R647 B.n709 B.n708 585
R648 B.n708 B.n707 585
R649 B.n46 B.n45 585
R650 B.n706 B.n46 585
R651 B.n704 B.n703 585
R652 B.n705 B.n704 585
R653 B.n702 B.n51 585
R654 B.n51 B.n50 585
R655 B.n701 B.n700 585
R656 B.n700 B.n699 585
R657 B.n53 B.n52 585
R658 B.n698 B.n53 585
R659 B.n696 B.n695 585
R660 B.n697 B.n696 585
R661 B.n694 B.n58 585
R662 B.n58 B.n57 585
R663 B.n693 B.n692 585
R664 B.n692 B.n691 585
R665 B.n60 B.n59 585
R666 B.n690 B.n60 585
R667 B.n688 B.n687 585
R668 B.n689 B.n688 585
R669 B.n686 B.n65 585
R670 B.n65 B.n64 585
R671 B.n685 B.n684 585
R672 B.n684 B.n683 585
R673 B.n67 B.n66 585
R674 B.n682 B.n67 585
R675 B.n680 B.n679 585
R676 B.n681 B.n680 585
R677 B.n678 B.n72 585
R678 B.n72 B.n71 585
R679 B.n677 B.n676 585
R680 B.n676 B.n675 585
R681 B.n74 B.n73 585
R682 B.n674 B.n74 585
R683 B.n672 B.n671 585
R684 B.n673 B.n672 585
R685 B.n670 B.n79 585
R686 B.n79 B.n78 585
R687 B.n669 B.n668 585
R688 B.n668 B.n667 585
R689 B.n81 B.n80 585
R690 B.n666 B.n81 585
R691 B.n664 B.n663 585
R692 B.n665 B.n664 585
R693 B.n662 B.n85 585
R694 B.n88 B.n85 585
R695 B.n661 B.n660 585
R696 B.n660 B.n659 585
R697 B.n87 B.n86 585
R698 B.n658 B.n87 585
R699 B.n656 B.n655 585
R700 B.n657 B.n656 585
R701 B.n654 B.n93 585
R702 B.n93 B.n92 585
R703 B.n653 B.n652 585
R704 B.n652 B.n651 585
R705 B.n95 B.n94 585
R706 B.n650 B.n95 585
R707 B.n648 B.n647 585
R708 B.n649 B.n648 585
R709 B.n757 B.n756 585
R710 B.n756 B.n755 585
R711 B.n335 B.n231 473.281
R712 B.n648 B.n100 473.281
R713 B.n337 B.n229 473.281
R714 B.n567 B.n98 473.281
R715 B.n568 B.n99 256.663
R716 B.n570 B.n99 256.663
R717 B.n576 B.n99 256.663
R718 B.n578 B.n99 256.663
R719 B.n584 B.n99 256.663
R720 B.n586 B.n99 256.663
R721 B.n592 B.n99 256.663
R722 B.n594 B.n99 256.663
R723 B.n601 B.n99 256.663
R724 B.n603 B.n99 256.663
R725 B.n609 B.n99 256.663
R726 B.n611 B.n99 256.663
R727 B.n617 B.n99 256.663
R728 B.n619 B.n99 256.663
R729 B.n625 B.n99 256.663
R730 B.n627 B.n99 256.663
R731 B.n633 B.n99 256.663
R732 B.n635 B.n99 256.663
R733 B.n641 B.n99 256.663
R734 B.n643 B.n99 256.663
R735 B.n330 B.n230 256.663
R736 B.n233 B.n230 256.663
R737 B.n323 B.n230 256.663
R738 B.n317 B.n230 256.663
R739 B.n315 B.n230 256.663
R740 B.n309 B.n230 256.663
R741 B.n307 B.n230 256.663
R742 B.n300 B.n230 256.663
R743 B.n298 B.n230 256.663
R744 B.n292 B.n230 256.663
R745 B.n290 B.n230 256.663
R746 B.n284 B.n230 256.663
R747 B.n249 B.n230 256.663
R748 B.n278 B.n230 256.663
R749 B.n272 B.n230 256.663
R750 B.n270 B.n230 256.663
R751 B.n264 B.n230 256.663
R752 B.n262 B.n230 256.663
R753 B.n256 B.n230 256.663
R754 B.n246 B.t10 239.02
R755 B.n240 B.t18 239.02
R756 B.n109 B.t21 239.02
R757 B.n116 B.t14 239.02
R758 B.n336 B.n230 164.1
R759 B.n649 B.n99 164.1
R760 B.n335 B.n225 163.367
R761 B.n343 B.n225 163.367
R762 B.n343 B.n223 163.367
R763 B.n347 B.n223 163.367
R764 B.n347 B.n217 163.367
R765 B.n356 B.n217 163.367
R766 B.n356 B.n215 163.367
R767 B.n360 B.n215 163.367
R768 B.n360 B.n210 163.367
R769 B.n368 B.n210 163.367
R770 B.n368 B.n208 163.367
R771 B.n372 B.n208 163.367
R772 B.n372 B.n202 163.367
R773 B.n380 B.n202 163.367
R774 B.n380 B.n200 163.367
R775 B.n384 B.n200 163.367
R776 B.n384 B.n194 163.367
R777 B.n392 B.n194 163.367
R778 B.n392 B.n192 163.367
R779 B.n396 B.n192 163.367
R780 B.n396 B.n186 163.367
R781 B.n404 B.n186 163.367
R782 B.n404 B.n184 163.367
R783 B.n408 B.n184 163.367
R784 B.n408 B.n178 163.367
R785 B.n416 B.n178 163.367
R786 B.n416 B.n176 163.367
R787 B.n420 B.n176 163.367
R788 B.n420 B.n170 163.367
R789 B.n428 B.n170 163.367
R790 B.n428 B.n168 163.367
R791 B.n432 B.n168 163.367
R792 B.n432 B.n162 163.367
R793 B.n440 B.n162 163.367
R794 B.n440 B.n160 163.367
R795 B.n444 B.n160 163.367
R796 B.n444 B.n154 163.367
R797 B.n452 B.n154 163.367
R798 B.n452 B.n152 163.367
R799 B.n456 B.n152 163.367
R800 B.n456 B.n146 163.367
R801 B.n464 B.n146 163.367
R802 B.n464 B.n144 163.367
R803 B.n468 B.n144 163.367
R804 B.n468 B.n138 163.367
R805 B.n476 B.n138 163.367
R806 B.n476 B.n136 163.367
R807 B.n480 B.n136 163.367
R808 B.n480 B.n130 163.367
R809 B.n489 B.n130 163.367
R810 B.n489 B.n128 163.367
R811 B.n493 B.n128 163.367
R812 B.n493 B.n2 163.367
R813 B.n756 B.n2 163.367
R814 B.n756 B.n3 163.367
R815 B.n752 B.n3 163.367
R816 B.n752 B.n9 163.367
R817 B.n748 B.n9 163.367
R818 B.n748 B.n11 163.367
R819 B.n744 B.n11 163.367
R820 B.n744 B.n16 163.367
R821 B.n740 B.n16 163.367
R822 B.n740 B.n18 163.367
R823 B.n736 B.n18 163.367
R824 B.n736 B.n23 163.367
R825 B.n732 B.n23 163.367
R826 B.n732 B.n25 163.367
R827 B.n728 B.n25 163.367
R828 B.n728 B.n30 163.367
R829 B.n724 B.n30 163.367
R830 B.n724 B.n32 163.367
R831 B.n720 B.n32 163.367
R832 B.n720 B.n37 163.367
R833 B.n716 B.n37 163.367
R834 B.n716 B.n39 163.367
R835 B.n712 B.n39 163.367
R836 B.n712 B.n44 163.367
R837 B.n708 B.n44 163.367
R838 B.n708 B.n46 163.367
R839 B.n704 B.n46 163.367
R840 B.n704 B.n51 163.367
R841 B.n700 B.n51 163.367
R842 B.n700 B.n53 163.367
R843 B.n696 B.n53 163.367
R844 B.n696 B.n58 163.367
R845 B.n692 B.n58 163.367
R846 B.n692 B.n60 163.367
R847 B.n688 B.n60 163.367
R848 B.n688 B.n65 163.367
R849 B.n684 B.n65 163.367
R850 B.n684 B.n67 163.367
R851 B.n680 B.n67 163.367
R852 B.n680 B.n72 163.367
R853 B.n676 B.n72 163.367
R854 B.n676 B.n74 163.367
R855 B.n672 B.n74 163.367
R856 B.n672 B.n79 163.367
R857 B.n668 B.n79 163.367
R858 B.n668 B.n81 163.367
R859 B.n664 B.n81 163.367
R860 B.n664 B.n85 163.367
R861 B.n660 B.n85 163.367
R862 B.n660 B.n87 163.367
R863 B.n656 B.n87 163.367
R864 B.n656 B.n93 163.367
R865 B.n652 B.n93 163.367
R866 B.n652 B.n95 163.367
R867 B.n648 B.n95 163.367
R868 B.n331 B.n329 163.367
R869 B.n329 B.n328 163.367
R870 B.n325 B.n324 163.367
R871 B.n322 B.n235 163.367
R872 B.n318 B.n316 163.367
R873 B.n314 B.n237 163.367
R874 B.n310 B.n308 163.367
R875 B.n306 B.n239 163.367
R876 B.n301 B.n299 163.367
R877 B.n297 B.n243 163.367
R878 B.n293 B.n291 163.367
R879 B.n289 B.n245 163.367
R880 B.n285 B.n283 163.367
R881 B.n280 B.n279 163.367
R882 B.n277 B.n251 163.367
R883 B.n273 B.n271 163.367
R884 B.n269 B.n253 163.367
R885 B.n265 B.n263 163.367
R886 B.n261 B.n255 163.367
R887 B.n257 B.n229 163.367
R888 B.n337 B.n227 163.367
R889 B.n341 B.n227 163.367
R890 B.n341 B.n221 163.367
R891 B.n349 B.n221 163.367
R892 B.n349 B.n219 163.367
R893 B.n353 B.n219 163.367
R894 B.n353 B.n214 163.367
R895 B.n362 B.n214 163.367
R896 B.n362 B.n212 163.367
R897 B.n366 B.n212 163.367
R898 B.n366 B.n206 163.367
R899 B.n374 B.n206 163.367
R900 B.n374 B.n204 163.367
R901 B.n378 B.n204 163.367
R902 B.n378 B.n197 163.367
R903 B.n386 B.n197 163.367
R904 B.n386 B.n195 163.367
R905 B.n390 B.n195 163.367
R906 B.n390 B.n190 163.367
R907 B.n398 B.n190 163.367
R908 B.n398 B.n188 163.367
R909 B.n402 B.n188 163.367
R910 B.n402 B.n181 163.367
R911 B.n410 B.n181 163.367
R912 B.n410 B.n179 163.367
R913 B.n414 B.n179 163.367
R914 B.n414 B.n174 163.367
R915 B.n422 B.n174 163.367
R916 B.n422 B.n172 163.367
R917 B.n426 B.n172 163.367
R918 B.n426 B.n165 163.367
R919 B.n434 B.n165 163.367
R920 B.n434 B.n163 163.367
R921 B.n438 B.n163 163.367
R922 B.n438 B.n158 163.367
R923 B.n446 B.n158 163.367
R924 B.n446 B.n156 163.367
R925 B.n450 B.n156 163.367
R926 B.n450 B.n150 163.367
R927 B.n458 B.n150 163.367
R928 B.n458 B.n148 163.367
R929 B.n462 B.n148 163.367
R930 B.n462 B.n142 163.367
R931 B.n470 B.n142 163.367
R932 B.n470 B.n140 163.367
R933 B.n474 B.n140 163.367
R934 B.n474 B.n134 163.367
R935 B.n482 B.n134 163.367
R936 B.n482 B.n132 163.367
R937 B.n487 B.n132 163.367
R938 B.n487 B.n126 163.367
R939 B.n495 B.n126 163.367
R940 B.n496 B.n495 163.367
R941 B.n496 B.n5 163.367
R942 B.n6 B.n5 163.367
R943 B.n7 B.n6 163.367
R944 B.n501 B.n7 163.367
R945 B.n501 B.n12 163.367
R946 B.n13 B.n12 163.367
R947 B.n14 B.n13 163.367
R948 B.n506 B.n14 163.367
R949 B.n506 B.n19 163.367
R950 B.n20 B.n19 163.367
R951 B.n21 B.n20 163.367
R952 B.n511 B.n21 163.367
R953 B.n511 B.n26 163.367
R954 B.n27 B.n26 163.367
R955 B.n28 B.n27 163.367
R956 B.n516 B.n28 163.367
R957 B.n516 B.n33 163.367
R958 B.n34 B.n33 163.367
R959 B.n35 B.n34 163.367
R960 B.n521 B.n35 163.367
R961 B.n521 B.n40 163.367
R962 B.n41 B.n40 163.367
R963 B.n42 B.n41 163.367
R964 B.n526 B.n42 163.367
R965 B.n526 B.n47 163.367
R966 B.n48 B.n47 163.367
R967 B.n49 B.n48 163.367
R968 B.n531 B.n49 163.367
R969 B.n531 B.n54 163.367
R970 B.n55 B.n54 163.367
R971 B.n56 B.n55 163.367
R972 B.n536 B.n56 163.367
R973 B.n536 B.n61 163.367
R974 B.n62 B.n61 163.367
R975 B.n63 B.n62 163.367
R976 B.n541 B.n63 163.367
R977 B.n541 B.n68 163.367
R978 B.n69 B.n68 163.367
R979 B.n70 B.n69 163.367
R980 B.n546 B.n70 163.367
R981 B.n546 B.n75 163.367
R982 B.n76 B.n75 163.367
R983 B.n77 B.n76 163.367
R984 B.n551 B.n77 163.367
R985 B.n551 B.n82 163.367
R986 B.n83 B.n82 163.367
R987 B.n84 B.n83 163.367
R988 B.n556 B.n84 163.367
R989 B.n556 B.n89 163.367
R990 B.n90 B.n89 163.367
R991 B.n91 B.n90 163.367
R992 B.n561 B.n91 163.367
R993 B.n561 B.n96 163.367
R994 B.n97 B.n96 163.367
R995 B.n98 B.n97 163.367
R996 B.n644 B.n642 163.367
R997 B.n640 B.n102 163.367
R998 B.n636 B.n634 163.367
R999 B.n632 B.n104 163.367
R1000 B.n628 B.n626 163.367
R1001 B.n624 B.n106 163.367
R1002 B.n620 B.n618 163.367
R1003 B.n616 B.n108 163.367
R1004 B.n612 B.n610 163.367
R1005 B.n608 B.n113 163.367
R1006 B.n604 B.n602 163.367
R1007 B.n600 B.n115 163.367
R1008 B.n595 B.n593 163.367
R1009 B.n591 B.n119 163.367
R1010 B.n587 B.n585 163.367
R1011 B.n583 B.n121 163.367
R1012 B.n579 B.n577 163.367
R1013 B.n575 B.n123 163.367
R1014 B.n571 B.n569 163.367
R1015 B.n246 B.t13 130.524
R1016 B.n116 B.t16 130.524
R1017 B.n240 B.t20 130.523
R1018 B.n109 B.t22 130.523
R1019 B.n336 B.n226 90.7221
R1020 B.n342 B.n226 90.7221
R1021 B.n342 B.n222 90.7221
R1022 B.n348 B.n222 90.7221
R1023 B.n348 B.n218 90.7221
R1024 B.n355 B.n218 90.7221
R1025 B.n355 B.n354 90.7221
R1026 B.n361 B.n211 90.7221
R1027 B.n367 B.n211 90.7221
R1028 B.n367 B.n207 90.7221
R1029 B.n373 B.n207 90.7221
R1030 B.n373 B.n203 90.7221
R1031 B.n379 B.n203 90.7221
R1032 B.n379 B.n198 90.7221
R1033 B.n385 B.n198 90.7221
R1034 B.n385 B.n199 90.7221
R1035 B.n391 B.n191 90.7221
R1036 B.n397 B.n191 90.7221
R1037 B.n397 B.n187 90.7221
R1038 B.n403 B.n187 90.7221
R1039 B.n403 B.n182 90.7221
R1040 B.n409 B.n182 90.7221
R1041 B.n409 B.n183 90.7221
R1042 B.n415 B.n175 90.7221
R1043 B.n421 B.n175 90.7221
R1044 B.n421 B.n171 90.7221
R1045 B.n427 B.n171 90.7221
R1046 B.n427 B.n166 90.7221
R1047 B.n433 B.n166 90.7221
R1048 B.n433 B.n167 90.7221
R1049 B.n439 B.n159 90.7221
R1050 B.n445 B.n159 90.7221
R1051 B.n445 B.n155 90.7221
R1052 B.n451 B.n155 90.7221
R1053 B.n451 B.n151 90.7221
R1054 B.n457 B.n151 90.7221
R1055 B.n463 B.n147 90.7221
R1056 B.n463 B.n143 90.7221
R1057 B.n469 B.n143 90.7221
R1058 B.n469 B.n139 90.7221
R1059 B.n475 B.n139 90.7221
R1060 B.n475 B.n135 90.7221
R1061 B.n481 B.n135 90.7221
R1062 B.n488 B.n131 90.7221
R1063 B.n488 B.n127 90.7221
R1064 B.n494 B.n127 90.7221
R1065 B.n494 B.n4 90.7221
R1066 B.n755 B.n4 90.7221
R1067 B.n755 B.n754 90.7221
R1068 B.n754 B.n753 90.7221
R1069 B.n753 B.n8 90.7221
R1070 B.n747 B.n8 90.7221
R1071 B.n747 B.n746 90.7221
R1072 B.n745 B.n15 90.7221
R1073 B.n739 B.n15 90.7221
R1074 B.n739 B.n738 90.7221
R1075 B.n738 B.n737 90.7221
R1076 B.n737 B.n22 90.7221
R1077 B.n731 B.n22 90.7221
R1078 B.n731 B.n730 90.7221
R1079 B.n729 B.n29 90.7221
R1080 B.n723 B.n29 90.7221
R1081 B.n723 B.n722 90.7221
R1082 B.n722 B.n721 90.7221
R1083 B.n721 B.n36 90.7221
R1084 B.n715 B.n36 90.7221
R1085 B.n714 B.n713 90.7221
R1086 B.n713 B.n43 90.7221
R1087 B.n707 B.n43 90.7221
R1088 B.n707 B.n706 90.7221
R1089 B.n706 B.n705 90.7221
R1090 B.n705 B.n50 90.7221
R1091 B.n699 B.n50 90.7221
R1092 B.n698 B.n697 90.7221
R1093 B.n697 B.n57 90.7221
R1094 B.n691 B.n57 90.7221
R1095 B.n691 B.n690 90.7221
R1096 B.n690 B.n689 90.7221
R1097 B.n689 B.n64 90.7221
R1098 B.n683 B.n64 90.7221
R1099 B.n682 B.n681 90.7221
R1100 B.n681 B.n71 90.7221
R1101 B.n675 B.n71 90.7221
R1102 B.n675 B.n674 90.7221
R1103 B.n674 B.n673 90.7221
R1104 B.n673 B.n78 90.7221
R1105 B.n667 B.n78 90.7221
R1106 B.n667 B.n666 90.7221
R1107 B.n666 B.n665 90.7221
R1108 B.n659 B.n88 90.7221
R1109 B.n659 B.n658 90.7221
R1110 B.n658 B.n657 90.7221
R1111 B.n657 B.n92 90.7221
R1112 B.n651 B.n92 90.7221
R1113 B.n651 B.n650 90.7221
R1114 B.n650 B.n649 90.7221
R1115 B.n199 B.t0 89.388
R1116 B.t3 B.n682 89.388
R1117 B.n457 B.t1 84.0514
R1118 B.t5 B.n729 84.0514
R1119 B.n247 B.t12 80.0997
R1120 B.n117 B.t17 80.0997
R1121 B.n241 B.t19 80.0978
R1122 B.n110 B.t23 80.0978
R1123 B.n361 B.t11 78.7149
R1124 B.n665 B.t15 78.7149
R1125 B.n330 B.n231 71.676
R1126 B.n328 B.n233 71.676
R1127 B.n324 B.n323 71.676
R1128 B.n317 B.n235 71.676
R1129 B.n316 B.n315 71.676
R1130 B.n309 B.n237 71.676
R1131 B.n308 B.n307 71.676
R1132 B.n300 B.n239 71.676
R1133 B.n299 B.n298 71.676
R1134 B.n292 B.n243 71.676
R1135 B.n291 B.n290 71.676
R1136 B.n284 B.n245 71.676
R1137 B.n283 B.n249 71.676
R1138 B.n279 B.n278 71.676
R1139 B.n272 B.n251 71.676
R1140 B.n271 B.n270 71.676
R1141 B.n264 B.n253 71.676
R1142 B.n263 B.n262 71.676
R1143 B.n256 B.n255 71.676
R1144 B.n643 B.n100 71.676
R1145 B.n642 B.n641 71.676
R1146 B.n635 B.n102 71.676
R1147 B.n634 B.n633 71.676
R1148 B.n627 B.n104 71.676
R1149 B.n626 B.n625 71.676
R1150 B.n619 B.n106 71.676
R1151 B.n618 B.n617 71.676
R1152 B.n611 B.n108 71.676
R1153 B.n610 B.n609 71.676
R1154 B.n603 B.n113 71.676
R1155 B.n602 B.n601 71.676
R1156 B.n594 B.n115 71.676
R1157 B.n593 B.n592 71.676
R1158 B.n586 B.n119 71.676
R1159 B.n585 B.n584 71.676
R1160 B.n578 B.n121 71.676
R1161 B.n577 B.n576 71.676
R1162 B.n570 B.n123 71.676
R1163 B.n569 B.n568 71.676
R1164 B.n568 B.n567 71.676
R1165 B.n571 B.n570 71.676
R1166 B.n576 B.n575 71.676
R1167 B.n579 B.n578 71.676
R1168 B.n584 B.n583 71.676
R1169 B.n587 B.n586 71.676
R1170 B.n592 B.n591 71.676
R1171 B.n595 B.n594 71.676
R1172 B.n601 B.n600 71.676
R1173 B.n604 B.n603 71.676
R1174 B.n609 B.n608 71.676
R1175 B.n612 B.n611 71.676
R1176 B.n617 B.n616 71.676
R1177 B.n620 B.n619 71.676
R1178 B.n625 B.n624 71.676
R1179 B.n628 B.n627 71.676
R1180 B.n633 B.n632 71.676
R1181 B.n636 B.n635 71.676
R1182 B.n641 B.n640 71.676
R1183 B.n644 B.n643 71.676
R1184 B.n331 B.n330 71.676
R1185 B.n325 B.n233 71.676
R1186 B.n323 B.n322 71.676
R1187 B.n318 B.n317 71.676
R1188 B.n315 B.n314 71.676
R1189 B.n310 B.n309 71.676
R1190 B.n307 B.n306 71.676
R1191 B.n301 B.n300 71.676
R1192 B.n298 B.n297 71.676
R1193 B.n293 B.n292 71.676
R1194 B.n290 B.n289 71.676
R1195 B.n285 B.n284 71.676
R1196 B.n280 B.n249 71.676
R1197 B.n278 B.n277 71.676
R1198 B.n273 B.n272 71.676
R1199 B.n270 B.n269 71.676
R1200 B.n265 B.n264 71.676
R1201 B.n262 B.n261 71.676
R1202 B.n257 B.n256 71.676
R1203 B.n439 B.t8 65.3735
R1204 B.n715 B.t6 65.3735
R1205 B.n248 B.n247 59.5399
R1206 B.n304 B.n241 59.5399
R1207 B.n111 B.n110 59.5399
R1208 B.n597 B.n117 59.5399
R1209 B.n183 B.t9 57.3686
R1210 B.t7 B.n698 57.3686
R1211 B.n481 B.t4 52.032
R1212 B.t2 B.n745 52.032
R1213 B.n247 B.n246 50.4247
R1214 B.n241 B.n240 50.4247
R1215 B.n110 B.n109 50.4247
R1216 B.n117 B.n116 50.4247
R1217 B.t4 B.n131 38.6906
R1218 B.n746 B.t2 38.6906
R1219 B.n415 B.t9 33.354
R1220 B.n699 B.t7 33.354
R1221 B.n647 B.n646 30.7517
R1222 B.n566 B.n565 30.7517
R1223 B.n338 B.n228 30.7517
R1224 B.n334 B.n333 30.7517
R1225 B.n167 B.t8 25.3492
R1226 B.t6 B.n714 25.3492
R1227 B B.n757 18.0485
R1228 B.n354 B.t11 12.0078
R1229 B.n88 B.t15 12.0078
R1230 B.n646 B.n645 10.6151
R1231 B.n645 B.n101 10.6151
R1232 B.n639 B.n101 10.6151
R1233 B.n639 B.n638 10.6151
R1234 B.n638 B.n637 10.6151
R1235 B.n637 B.n103 10.6151
R1236 B.n631 B.n103 10.6151
R1237 B.n631 B.n630 10.6151
R1238 B.n630 B.n629 10.6151
R1239 B.n629 B.n105 10.6151
R1240 B.n623 B.n105 10.6151
R1241 B.n623 B.n622 10.6151
R1242 B.n622 B.n621 10.6151
R1243 B.n621 B.n107 10.6151
R1244 B.n615 B.n614 10.6151
R1245 B.n614 B.n613 10.6151
R1246 B.n613 B.n112 10.6151
R1247 B.n607 B.n112 10.6151
R1248 B.n607 B.n606 10.6151
R1249 B.n606 B.n605 10.6151
R1250 B.n605 B.n114 10.6151
R1251 B.n599 B.n114 10.6151
R1252 B.n599 B.n598 10.6151
R1253 B.n596 B.n118 10.6151
R1254 B.n590 B.n118 10.6151
R1255 B.n590 B.n589 10.6151
R1256 B.n589 B.n588 10.6151
R1257 B.n588 B.n120 10.6151
R1258 B.n582 B.n120 10.6151
R1259 B.n582 B.n581 10.6151
R1260 B.n581 B.n580 10.6151
R1261 B.n580 B.n122 10.6151
R1262 B.n574 B.n122 10.6151
R1263 B.n574 B.n573 10.6151
R1264 B.n573 B.n572 10.6151
R1265 B.n572 B.n124 10.6151
R1266 B.n566 B.n124 10.6151
R1267 B.n339 B.n338 10.6151
R1268 B.n340 B.n339 10.6151
R1269 B.n340 B.n220 10.6151
R1270 B.n350 B.n220 10.6151
R1271 B.n351 B.n350 10.6151
R1272 B.n352 B.n351 10.6151
R1273 B.n352 B.n213 10.6151
R1274 B.n363 B.n213 10.6151
R1275 B.n364 B.n363 10.6151
R1276 B.n365 B.n364 10.6151
R1277 B.n365 B.n205 10.6151
R1278 B.n375 B.n205 10.6151
R1279 B.n376 B.n375 10.6151
R1280 B.n377 B.n376 10.6151
R1281 B.n377 B.n196 10.6151
R1282 B.n387 B.n196 10.6151
R1283 B.n388 B.n387 10.6151
R1284 B.n389 B.n388 10.6151
R1285 B.n389 B.n189 10.6151
R1286 B.n399 B.n189 10.6151
R1287 B.n400 B.n399 10.6151
R1288 B.n401 B.n400 10.6151
R1289 B.n401 B.n180 10.6151
R1290 B.n411 B.n180 10.6151
R1291 B.n412 B.n411 10.6151
R1292 B.n413 B.n412 10.6151
R1293 B.n413 B.n173 10.6151
R1294 B.n423 B.n173 10.6151
R1295 B.n424 B.n423 10.6151
R1296 B.n425 B.n424 10.6151
R1297 B.n425 B.n164 10.6151
R1298 B.n435 B.n164 10.6151
R1299 B.n436 B.n435 10.6151
R1300 B.n437 B.n436 10.6151
R1301 B.n437 B.n157 10.6151
R1302 B.n447 B.n157 10.6151
R1303 B.n448 B.n447 10.6151
R1304 B.n449 B.n448 10.6151
R1305 B.n449 B.n149 10.6151
R1306 B.n459 B.n149 10.6151
R1307 B.n460 B.n459 10.6151
R1308 B.n461 B.n460 10.6151
R1309 B.n461 B.n141 10.6151
R1310 B.n471 B.n141 10.6151
R1311 B.n472 B.n471 10.6151
R1312 B.n473 B.n472 10.6151
R1313 B.n473 B.n133 10.6151
R1314 B.n483 B.n133 10.6151
R1315 B.n484 B.n483 10.6151
R1316 B.n486 B.n484 10.6151
R1317 B.n486 B.n485 10.6151
R1318 B.n485 B.n125 10.6151
R1319 B.n497 B.n125 10.6151
R1320 B.n498 B.n497 10.6151
R1321 B.n499 B.n498 10.6151
R1322 B.n500 B.n499 10.6151
R1323 B.n502 B.n500 10.6151
R1324 B.n503 B.n502 10.6151
R1325 B.n504 B.n503 10.6151
R1326 B.n505 B.n504 10.6151
R1327 B.n507 B.n505 10.6151
R1328 B.n508 B.n507 10.6151
R1329 B.n509 B.n508 10.6151
R1330 B.n510 B.n509 10.6151
R1331 B.n512 B.n510 10.6151
R1332 B.n513 B.n512 10.6151
R1333 B.n514 B.n513 10.6151
R1334 B.n515 B.n514 10.6151
R1335 B.n517 B.n515 10.6151
R1336 B.n518 B.n517 10.6151
R1337 B.n519 B.n518 10.6151
R1338 B.n520 B.n519 10.6151
R1339 B.n522 B.n520 10.6151
R1340 B.n523 B.n522 10.6151
R1341 B.n524 B.n523 10.6151
R1342 B.n525 B.n524 10.6151
R1343 B.n527 B.n525 10.6151
R1344 B.n528 B.n527 10.6151
R1345 B.n529 B.n528 10.6151
R1346 B.n530 B.n529 10.6151
R1347 B.n532 B.n530 10.6151
R1348 B.n533 B.n532 10.6151
R1349 B.n534 B.n533 10.6151
R1350 B.n535 B.n534 10.6151
R1351 B.n537 B.n535 10.6151
R1352 B.n538 B.n537 10.6151
R1353 B.n539 B.n538 10.6151
R1354 B.n540 B.n539 10.6151
R1355 B.n542 B.n540 10.6151
R1356 B.n543 B.n542 10.6151
R1357 B.n544 B.n543 10.6151
R1358 B.n545 B.n544 10.6151
R1359 B.n547 B.n545 10.6151
R1360 B.n548 B.n547 10.6151
R1361 B.n549 B.n548 10.6151
R1362 B.n550 B.n549 10.6151
R1363 B.n552 B.n550 10.6151
R1364 B.n553 B.n552 10.6151
R1365 B.n554 B.n553 10.6151
R1366 B.n555 B.n554 10.6151
R1367 B.n557 B.n555 10.6151
R1368 B.n558 B.n557 10.6151
R1369 B.n559 B.n558 10.6151
R1370 B.n560 B.n559 10.6151
R1371 B.n562 B.n560 10.6151
R1372 B.n563 B.n562 10.6151
R1373 B.n564 B.n563 10.6151
R1374 B.n565 B.n564 10.6151
R1375 B.n333 B.n332 10.6151
R1376 B.n332 B.n232 10.6151
R1377 B.n327 B.n232 10.6151
R1378 B.n327 B.n326 10.6151
R1379 B.n326 B.n234 10.6151
R1380 B.n321 B.n234 10.6151
R1381 B.n321 B.n320 10.6151
R1382 B.n320 B.n319 10.6151
R1383 B.n319 B.n236 10.6151
R1384 B.n313 B.n236 10.6151
R1385 B.n313 B.n312 10.6151
R1386 B.n312 B.n311 10.6151
R1387 B.n311 B.n238 10.6151
R1388 B.n305 B.n238 10.6151
R1389 B.n303 B.n302 10.6151
R1390 B.n302 B.n242 10.6151
R1391 B.n296 B.n242 10.6151
R1392 B.n296 B.n295 10.6151
R1393 B.n295 B.n294 10.6151
R1394 B.n294 B.n244 10.6151
R1395 B.n288 B.n244 10.6151
R1396 B.n288 B.n287 10.6151
R1397 B.n287 B.n286 10.6151
R1398 B.n282 B.n281 10.6151
R1399 B.n281 B.n250 10.6151
R1400 B.n276 B.n250 10.6151
R1401 B.n276 B.n275 10.6151
R1402 B.n275 B.n274 10.6151
R1403 B.n274 B.n252 10.6151
R1404 B.n268 B.n252 10.6151
R1405 B.n268 B.n267 10.6151
R1406 B.n267 B.n266 10.6151
R1407 B.n266 B.n254 10.6151
R1408 B.n260 B.n254 10.6151
R1409 B.n260 B.n259 10.6151
R1410 B.n259 B.n258 10.6151
R1411 B.n258 B.n228 10.6151
R1412 B.n334 B.n224 10.6151
R1413 B.n344 B.n224 10.6151
R1414 B.n345 B.n344 10.6151
R1415 B.n346 B.n345 10.6151
R1416 B.n346 B.n216 10.6151
R1417 B.n357 B.n216 10.6151
R1418 B.n358 B.n357 10.6151
R1419 B.n359 B.n358 10.6151
R1420 B.n359 B.n209 10.6151
R1421 B.n369 B.n209 10.6151
R1422 B.n370 B.n369 10.6151
R1423 B.n371 B.n370 10.6151
R1424 B.n371 B.n201 10.6151
R1425 B.n381 B.n201 10.6151
R1426 B.n382 B.n381 10.6151
R1427 B.n383 B.n382 10.6151
R1428 B.n383 B.n193 10.6151
R1429 B.n393 B.n193 10.6151
R1430 B.n394 B.n393 10.6151
R1431 B.n395 B.n394 10.6151
R1432 B.n395 B.n185 10.6151
R1433 B.n405 B.n185 10.6151
R1434 B.n406 B.n405 10.6151
R1435 B.n407 B.n406 10.6151
R1436 B.n407 B.n177 10.6151
R1437 B.n417 B.n177 10.6151
R1438 B.n418 B.n417 10.6151
R1439 B.n419 B.n418 10.6151
R1440 B.n419 B.n169 10.6151
R1441 B.n429 B.n169 10.6151
R1442 B.n430 B.n429 10.6151
R1443 B.n431 B.n430 10.6151
R1444 B.n431 B.n161 10.6151
R1445 B.n441 B.n161 10.6151
R1446 B.n442 B.n441 10.6151
R1447 B.n443 B.n442 10.6151
R1448 B.n443 B.n153 10.6151
R1449 B.n453 B.n153 10.6151
R1450 B.n454 B.n453 10.6151
R1451 B.n455 B.n454 10.6151
R1452 B.n455 B.n145 10.6151
R1453 B.n465 B.n145 10.6151
R1454 B.n466 B.n465 10.6151
R1455 B.n467 B.n466 10.6151
R1456 B.n467 B.n137 10.6151
R1457 B.n477 B.n137 10.6151
R1458 B.n478 B.n477 10.6151
R1459 B.n479 B.n478 10.6151
R1460 B.n479 B.n129 10.6151
R1461 B.n490 B.n129 10.6151
R1462 B.n491 B.n490 10.6151
R1463 B.n492 B.n491 10.6151
R1464 B.n492 B.n0 10.6151
R1465 B.n751 B.n1 10.6151
R1466 B.n751 B.n750 10.6151
R1467 B.n750 B.n749 10.6151
R1468 B.n749 B.n10 10.6151
R1469 B.n743 B.n10 10.6151
R1470 B.n743 B.n742 10.6151
R1471 B.n742 B.n741 10.6151
R1472 B.n741 B.n17 10.6151
R1473 B.n735 B.n17 10.6151
R1474 B.n735 B.n734 10.6151
R1475 B.n734 B.n733 10.6151
R1476 B.n733 B.n24 10.6151
R1477 B.n727 B.n24 10.6151
R1478 B.n727 B.n726 10.6151
R1479 B.n726 B.n725 10.6151
R1480 B.n725 B.n31 10.6151
R1481 B.n719 B.n31 10.6151
R1482 B.n719 B.n718 10.6151
R1483 B.n718 B.n717 10.6151
R1484 B.n717 B.n38 10.6151
R1485 B.n711 B.n38 10.6151
R1486 B.n711 B.n710 10.6151
R1487 B.n710 B.n709 10.6151
R1488 B.n709 B.n45 10.6151
R1489 B.n703 B.n45 10.6151
R1490 B.n703 B.n702 10.6151
R1491 B.n702 B.n701 10.6151
R1492 B.n701 B.n52 10.6151
R1493 B.n695 B.n52 10.6151
R1494 B.n695 B.n694 10.6151
R1495 B.n694 B.n693 10.6151
R1496 B.n693 B.n59 10.6151
R1497 B.n687 B.n59 10.6151
R1498 B.n687 B.n686 10.6151
R1499 B.n686 B.n685 10.6151
R1500 B.n685 B.n66 10.6151
R1501 B.n679 B.n66 10.6151
R1502 B.n679 B.n678 10.6151
R1503 B.n678 B.n677 10.6151
R1504 B.n677 B.n73 10.6151
R1505 B.n671 B.n73 10.6151
R1506 B.n671 B.n670 10.6151
R1507 B.n670 B.n669 10.6151
R1508 B.n669 B.n80 10.6151
R1509 B.n663 B.n80 10.6151
R1510 B.n663 B.n662 10.6151
R1511 B.n662 B.n661 10.6151
R1512 B.n661 B.n86 10.6151
R1513 B.n655 B.n86 10.6151
R1514 B.n655 B.n654 10.6151
R1515 B.n654 B.n653 10.6151
R1516 B.n653 B.n94 10.6151
R1517 B.n647 B.n94 10.6151
R1518 B.n111 B.n107 9.36635
R1519 B.n597 B.n596 9.36635
R1520 B.n305 B.n304 9.36635
R1521 B.n282 B.n248 9.36635
R1522 B.t1 B.n147 6.67121
R1523 B.n730 B.t5 6.67121
R1524 B.n757 B.n0 2.81026
R1525 B.n757 B.n1 2.81026
R1526 B.n391 B.t0 1.33464
R1527 B.n683 B.t3 1.33464
R1528 B.n615 B.n111 1.24928
R1529 B.n598 B.n597 1.24928
R1530 B.n304 B.n303 1.24928
R1531 B.n286 B.n248 1.24928
R1532 VN.n71 VN.n37 161.3
R1533 VN.n70 VN.n69 161.3
R1534 VN.n68 VN.n38 161.3
R1535 VN.n67 VN.n66 161.3
R1536 VN.n65 VN.n39 161.3
R1537 VN.n63 VN.n62 161.3
R1538 VN.n61 VN.n40 161.3
R1539 VN.n60 VN.n59 161.3
R1540 VN.n58 VN.n41 161.3
R1541 VN.n57 VN.n56 161.3
R1542 VN.n55 VN.n42 161.3
R1543 VN.n54 VN.n53 161.3
R1544 VN.n52 VN.n43 161.3
R1545 VN.n51 VN.n50 161.3
R1546 VN.n49 VN.n44 161.3
R1547 VN.n48 VN.n47 161.3
R1548 VN.n34 VN.n0 161.3
R1549 VN.n33 VN.n32 161.3
R1550 VN.n31 VN.n1 161.3
R1551 VN.n30 VN.n29 161.3
R1552 VN.n28 VN.n2 161.3
R1553 VN.n26 VN.n25 161.3
R1554 VN.n24 VN.n3 161.3
R1555 VN.n23 VN.n22 161.3
R1556 VN.n21 VN.n4 161.3
R1557 VN.n20 VN.n19 161.3
R1558 VN.n18 VN.n5 161.3
R1559 VN.n17 VN.n16 161.3
R1560 VN.n15 VN.n6 161.3
R1561 VN.n14 VN.n13 161.3
R1562 VN.n12 VN.n7 161.3
R1563 VN.n11 VN.n10 161.3
R1564 VN.n36 VN.n35 100.969
R1565 VN.n73 VN.n72 100.969
R1566 VN.n9 VN.n8 67.1934
R1567 VN.n46 VN.n45 67.1934
R1568 VN.n8 VN.t9 62.4054
R1569 VN.n45 VN.t2 62.4054
R1570 VN.n15 VN.n14 56.5193
R1571 VN.n22 VN.n21 56.5193
R1572 VN.n52 VN.n51 56.5193
R1573 VN.n59 VN.n58 56.5193
R1574 VN.n29 VN.n1 50.2061
R1575 VN.n66 VN.n38 50.2061
R1576 VN VN.n73 44.6951
R1577 VN.n5 VN.t0 31.5322
R1578 VN.n9 VN.t7 31.5322
R1579 VN.n27 VN.t3 31.5322
R1580 VN.n35 VN.t6 31.5322
R1581 VN.n42 VN.t4 31.5322
R1582 VN.n46 VN.t1 31.5322
R1583 VN.n64 VN.t8 31.5322
R1584 VN.n72 VN.t5 31.5322
R1585 VN.n33 VN.n1 30.7807
R1586 VN.n70 VN.n38 30.7807
R1587 VN.n10 VN.n7 24.4675
R1588 VN.n14 VN.n7 24.4675
R1589 VN.n16 VN.n15 24.4675
R1590 VN.n16 VN.n5 24.4675
R1591 VN.n20 VN.n5 24.4675
R1592 VN.n21 VN.n20 24.4675
R1593 VN.n22 VN.n3 24.4675
R1594 VN.n26 VN.n3 24.4675
R1595 VN.n29 VN.n28 24.4675
R1596 VN.n34 VN.n33 24.4675
R1597 VN.n51 VN.n44 24.4675
R1598 VN.n47 VN.n44 24.4675
R1599 VN.n58 VN.n57 24.4675
R1600 VN.n57 VN.n42 24.4675
R1601 VN.n53 VN.n42 24.4675
R1602 VN.n53 VN.n52 24.4675
R1603 VN.n66 VN.n65 24.4675
R1604 VN.n63 VN.n40 24.4675
R1605 VN.n59 VN.n40 24.4675
R1606 VN.n71 VN.n70 24.4675
R1607 VN.n28 VN.n27 19.5741
R1608 VN.n65 VN.n64 19.5741
R1609 VN.n48 VN.n45 10.026
R1610 VN.n11 VN.n8 10.026
R1611 VN.n35 VN.n34 9.7873
R1612 VN.n72 VN.n71 9.7873
R1613 VN.n10 VN.n9 4.8939
R1614 VN.n27 VN.n26 4.8939
R1615 VN.n47 VN.n46 4.8939
R1616 VN.n64 VN.n63 4.8939
R1617 VN.n73 VN.n37 0.278367
R1618 VN.n36 VN.n0 0.278367
R1619 VN.n69 VN.n37 0.189894
R1620 VN.n69 VN.n68 0.189894
R1621 VN.n68 VN.n67 0.189894
R1622 VN.n67 VN.n39 0.189894
R1623 VN.n62 VN.n39 0.189894
R1624 VN.n62 VN.n61 0.189894
R1625 VN.n61 VN.n60 0.189894
R1626 VN.n60 VN.n41 0.189894
R1627 VN.n56 VN.n41 0.189894
R1628 VN.n56 VN.n55 0.189894
R1629 VN.n55 VN.n54 0.189894
R1630 VN.n54 VN.n43 0.189894
R1631 VN.n50 VN.n43 0.189894
R1632 VN.n50 VN.n49 0.189894
R1633 VN.n49 VN.n48 0.189894
R1634 VN.n12 VN.n11 0.189894
R1635 VN.n13 VN.n12 0.189894
R1636 VN.n13 VN.n6 0.189894
R1637 VN.n17 VN.n6 0.189894
R1638 VN.n18 VN.n17 0.189894
R1639 VN.n19 VN.n18 0.189894
R1640 VN.n19 VN.n4 0.189894
R1641 VN.n23 VN.n4 0.189894
R1642 VN.n24 VN.n23 0.189894
R1643 VN.n25 VN.n24 0.189894
R1644 VN.n25 VN.n2 0.189894
R1645 VN.n30 VN.n2 0.189894
R1646 VN.n31 VN.n30 0.189894
R1647 VN.n32 VN.n31 0.189894
R1648 VN.n32 VN.n0 0.189894
R1649 VN VN.n36 0.153454
R1650 VDD2.n1 VDD2.t0 93.8091
R1651 VDD2.n4 VDD2.t4 91.568
R1652 VDD2.n3 VDD2.n2 86.5268
R1653 VDD2 VDD2.n7 86.524
R1654 VDD2.n6 VDD2.n5 84.9013
R1655 VDD2.n1 VDD2.n0 84.9011
R1656 VDD2.n4 VDD2.n3 36.9222
R1657 VDD2.n7 VDD2.t8 6.66717
R1658 VDD2.n7 VDD2.t7 6.66717
R1659 VDD2.n5 VDD2.t1 6.66717
R1660 VDD2.n5 VDD2.t5 6.66717
R1661 VDD2.n2 VDD2.t6 6.66717
R1662 VDD2.n2 VDD2.t3 6.66717
R1663 VDD2.n0 VDD2.t2 6.66717
R1664 VDD2.n0 VDD2.t9 6.66717
R1665 VDD2.n6 VDD2.n4 2.24188
R1666 VDD2 VDD2.n6 0.619035
R1667 VDD2.n3 VDD2.n1 0.505499
C0 VP VTAIL 4.10096f
C1 VP VN 6.25049f
C2 VTAIL VN 4.0868f
C3 VDD1 VP 3.33303f
C4 VDD1 VTAIL 5.91218f
C5 VDD1 VN 0.157862f
C6 VP VDD2 0.546826f
C7 VDD2 VTAIL 5.9629f
C8 VDD2 VN 2.94726f
C9 VDD1 VDD2 1.95869f
C10 VDD2 B 5.182257f
C11 VDD1 B 5.176446f
C12 VTAIL B 3.956847f
C13 VN B 15.741529f
C14 VP B 14.22704f
C15 VDD2.t0 B 0.518165f
C16 VDD2.t2 B 0.053968f
C17 VDD2.t9 B 0.053968f
C18 VDD2.n0 B 0.397494f
C19 VDD2.n1 B 0.755446f
C20 VDD2.t6 B 0.053968f
C21 VDD2.t3 B 0.053968f
C22 VDD2.n2 B 0.406337f
C23 VDD2.n3 B 2.00334f
C24 VDD2.t4 B 0.508953f
C25 VDD2.n4 B 2.06093f
C26 VDD2.t1 B 0.053968f
C27 VDD2.t5 B 0.053968f
C28 VDD2.n5 B 0.397495f
C29 VDD2.n6 B 0.386427f
C30 VDD2.t8 B 0.053968f
C31 VDD2.t7 B 0.053968f
C32 VDD2.n7 B 0.406311f
C33 VN.n0 B 0.038209f
C34 VN.t6 B 0.486114f
C35 VN.n1 B 0.027378f
C36 VN.n2 B 0.028981f
C37 VN.t3 B 0.486114f
C38 VN.n3 B 0.054014f
C39 VN.n4 B 0.028981f
C40 VN.t0 B 0.486114f
C41 VN.n5 B 0.236537f
C42 VN.n6 B 0.028981f
C43 VN.n7 B 0.054014f
C44 VN.t9 B 0.666291f
C45 VN.n8 B 0.277868f
C46 VN.t7 B 0.486114f
C47 VN.n9 B 0.278697f
C48 VN.n10 B 0.03268f
C49 VN.n11 B 0.248276f
C50 VN.n12 B 0.028981f
C51 VN.n13 B 0.028981f
C52 VN.n14 B 0.038269f
C53 VN.n15 B 0.046345f
C54 VN.n16 B 0.054014f
C55 VN.n17 B 0.028981f
C56 VN.n18 B 0.028981f
C57 VN.n19 B 0.028981f
C58 VN.n20 B 0.054014f
C59 VN.n21 B 0.046345f
C60 VN.n22 B 0.038269f
C61 VN.n23 B 0.028981f
C62 VN.n24 B 0.028981f
C63 VN.n25 B 0.028981f
C64 VN.n26 B 0.03268f
C65 VN.n27 B 0.20919f
C66 VN.n28 B 0.04868f
C67 VN.n29 B 0.053191f
C68 VN.n30 B 0.028981f
C69 VN.n31 B 0.028981f
C70 VN.n32 B 0.028981f
C71 VN.n33 B 0.058059f
C72 VN.n34 B 0.038014f
C73 VN.n35 B 0.293044f
C74 VN.n36 B 0.044306f
C75 VN.n37 B 0.038209f
C76 VN.t5 B 0.486114f
C77 VN.n38 B 0.027378f
C78 VN.n39 B 0.028981f
C79 VN.t8 B 0.486114f
C80 VN.n40 B 0.054014f
C81 VN.n41 B 0.028981f
C82 VN.t4 B 0.486114f
C83 VN.n42 B 0.236537f
C84 VN.n43 B 0.028981f
C85 VN.n44 B 0.054014f
C86 VN.t2 B 0.666291f
C87 VN.n45 B 0.277868f
C88 VN.t1 B 0.486114f
C89 VN.n46 B 0.278697f
C90 VN.n47 B 0.03268f
C91 VN.n48 B 0.248276f
C92 VN.n49 B 0.028981f
C93 VN.n50 B 0.028981f
C94 VN.n51 B 0.038269f
C95 VN.n52 B 0.046345f
C96 VN.n53 B 0.054014f
C97 VN.n54 B 0.028981f
C98 VN.n55 B 0.028981f
C99 VN.n56 B 0.028981f
C100 VN.n57 B 0.054014f
C101 VN.n58 B 0.046345f
C102 VN.n59 B 0.038269f
C103 VN.n60 B 0.028981f
C104 VN.n61 B 0.028981f
C105 VN.n62 B 0.028981f
C106 VN.n63 B 0.03268f
C107 VN.n64 B 0.20919f
C108 VN.n65 B 0.04868f
C109 VN.n66 B 0.053191f
C110 VN.n67 B 0.028981f
C111 VN.n68 B 0.028981f
C112 VN.n69 B 0.028981f
C113 VN.n70 B 0.058059f
C114 VN.n71 B 0.038014f
C115 VN.n72 B 0.293044f
C116 VN.n73 B 1.35952f
C117 VDD1.t2 B 0.530569f
C118 VDD1.t0 B 0.055259f
C119 VDD1.t1 B 0.055259f
C120 VDD1.n0 B 0.40701f
C121 VDD1.n1 B 0.781059f
C122 VDD1.t9 B 0.530568f
C123 VDD1.t6 B 0.055259f
C124 VDD1.t5 B 0.055259f
C125 VDD1.n2 B 0.407009f
C126 VDD1.n3 B 0.773529f
C127 VDD1.t7 B 0.055259f
C128 VDD1.t8 B 0.055259f
C129 VDD1.n4 B 0.416063f
C130 VDD1.n5 B 2.15362f
C131 VDD1.t3 B 0.055259f
C132 VDD1.t4 B 0.055259f
C133 VDD1.n6 B 0.407009f
C134 VDD1.n7 B 2.18144f
C135 VTAIL.t2 B 0.077071f
C136 VTAIL.t17 B 0.077071f
C137 VTAIL.n0 B 0.508257f
C138 VTAIL.n1 B 0.616344f
C139 VTAIL.t9 B 0.661355f
C140 VTAIL.n2 B 0.726575f
C141 VTAIL.t10 B 0.077071f
C142 VTAIL.t8 B 0.077071f
C143 VTAIL.n3 B 0.508257f
C144 VTAIL.n4 B 0.738349f
C145 VTAIL.t13 B 0.077071f
C146 VTAIL.t12 B 0.077071f
C147 VTAIL.n5 B 0.508257f
C148 VTAIL.n6 B 1.69251f
C149 VTAIL.t0 B 0.077071f
C150 VTAIL.t15 B 0.077071f
C151 VTAIL.n7 B 0.508259f
C152 VTAIL.n8 B 1.6925f
C153 VTAIL.t16 B 0.077071f
C154 VTAIL.t1 B 0.077071f
C155 VTAIL.n9 B 0.508259f
C156 VTAIL.n10 B 0.738346f
C157 VTAIL.t4 B 0.661357f
C158 VTAIL.n11 B 0.726573f
C159 VTAIL.t5 B 0.077071f
C160 VTAIL.t7 B 0.077071f
C161 VTAIL.n12 B 0.508259f
C162 VTAIL.n13 B 0.669477f
C163 VTAIL.t11 B 0.077071f
C164 VTAIL.t14 B 0.077071f
C165 VTAIL.n14 B 0.508259f
C166 VTAIL.n15 B 0.738346f
C167 VTAIL.t6 B 0.661355f
C168 VTAIL.n16 B 1.51243f
C169 VTAIL.t3 B 0.661355f
C170 VTAIL.n17 B 1.51243f
C171 VTAIL.t19 B 0.077071f
C172 VTAIL.t18 B 0.077071f
C173 VTAIL.n18 B 0.508257f
C174 VTAIL.n19 B 0.554316f
C175 VP.n0 B 0.039479f
C176 VP.t1 B 0.502273f
C177 VP.n1 B 0.028288f
C178 VP.n2 B 0.029945f
C179 VP.t2 B 0.502273f
C180 VP.n3 B 0.055809f
C181 VP.n4 B 0.029945f
C182 VP.t4 B 0.502273f
C183 VP.n5 B 0.2444f
C184 VP.n6 B 0.029945f
C185 VP.n7 B 0.055809f
C186 VP.n8 B 0.029945f
C187 VP.t3 B 0.502273f
C188 VP.n9 B 0.028288f
C189 VP.n10 B 0.039479f
C190 VP.t0 B 0.502273f
C191 VP.n11 B 0.039479f
C192 VP.t5 B 0.502273f
C193 VP.n12 B 0.028288f
C194 VP.n13 B 0.029945f
C195 VP.t6 B 0.502273f
C196 VP.n14 B 0.055809f
C197 VP.n15 B 0.029945f
C198 VP.t8 B 0.502273f
C199 VP.n16 B 0.2444f
C200 VP.n17 B 0.029945f
C201 VP.n18 B 0.055809f
C202 VP.t7 B 0.688439f
C203 VP.n19 B 0.287104f
C204 VP.t9 B 0.502273f
C205 VP.n20 B 0.287961f
C206 VP.n21 B 0.033766f
C207 VP.n22 B 0.256529f
C208 VP.n23 B 0.029945f
C209 VP.n24 B 0.029945f
C210 VP.n25 B 0.039542f
C211 VP.n26 B 0.047886f
C212 VP.n27 B 0.055809f
C213 VP.n28 B 0.029945f
C214 VP.n29 B 0.029945f
C215 VP.n30 B 0.029945f
C216 VP.n31 B 0.055809f
C217 VP.n32 B 0.047886f
C218 VP.n33 B 0.039542f
C219 VP.n34 B 0.029945f
C220 VP.n35 B 0.029945f
C221 VP.n36 B 0.029945f
C222 VP.n37 B 0.033766f
C223 VP.n38 B 0.216144f
C224 VP.n39 B 0.050299f
C225 VP.n40 B 0.054959f
C226 VP.n41 B 0.029945f
C227 VP.n42 B 0.029945f
C228 VP.n43 B 0.029945f
C229 VP.n44 B 0.059989f
C230 VP.n45 B 0.039277f
C231 VP.n46 B 0.302784f
C232 VP.n47 B 1.38829f
C233 VP.n48 B 1.41253f
C234 VP.n49 B 0.302784f
C235 VP.n50 B 0.039277f
C236 VP.n51 B 0.059989f
C237 VP.n52 B 0.029945f
C238 VP.n53 B 0.029945f
C239 VP.n54 B 0.029945f
C240 VP.n55 B 0.054959f
C241 VP.n56 B 0.050299f
C242 VP.n57 B 0.216144f
C243 VP.n58 B 0.033766f
C244 VP.n59 B 0.029945f
C245 VP.n60 B 0.029945f
C246 VP.n61 B 0.029945f
C247 VP.n62 B 0.039542f
C248 VP.n63 B 0.047886f
C249 VP.n64 B 0.055809f
C250 VP.n65 B 0.029945f
C251 VP.n66 B 0.029945f
C252 VP.n67 B 0.029945f
C253 VP.n68 B 0.055809f
C254 VP.n69 B 0.047886f
C255 VP.n70 B 0.039542f
C256 VP.n71 B 0.029945f
C257 VP.n72 B 0.029945f
C258 VP.n73 B 0.029945f
C259 VP.n74 B 0.033766f
C260 VP.n75 B 0.216144f
C261 VP.n76 B 0.050299f
C262 VP.n77 B 0.054959f
C263 VP.n78 B 0.029945f
C264 VP.n79 B 0.029945f
C265 VP.n80 B 0.029945f
C266 VP.n81 B 0.059989f
C267 VP.n82 B 0.039277f
C268 VP.n83 B 0.302784f
C269 VP.n84 B 0.045779f
.ends

