* NGSPICE file created from diff_pair_sample_1012.ext - technology: sky130A

.subckt diff_pair_sample_1012 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X1 B.t11 B.t9 B.t10 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=0 ps=0 w=13.62 l=2.47
X2 B.t8 B.t6 B.t7 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=0 ps=0 w=13.62 l=2.47
X3 VDD2.t7 VN.t0 VTAIL.t3 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=5.3118 ps=28.02 w=13.62 l=2.47
X4 VTAIL.t14 VP.t1 VDD1.t6 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=2.2473 ps=13.95 w=13.62 l=2.47
X5 VDD2.t6 VN.t1 VTAIL.t6 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=5.3118 ps=28.02 w=13.62 l=2.47
X6 B.t5 B.t3 B.t4 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=0 ps=0 w=13.62 l=2.47
X7 VTAIL.t7 VN.t2 VDD2.t5 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=2.2473 ps=13.95 w=13.62 l=2.47
X8 VDD2.t4 VN.t3 VTAIL.t5 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X9 B.t2 B.t0 B.t1 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=0 ps=0 w=13.62 l=2.47
X10 VDD1.t5 VP.t2 VTAIL.t13 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=5.3118 ps=28.02 w=13.62 l=2.47
X11 VTAIL.t2 VN.t4 VDD2.t3 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X12 VDD1.t4 VP.t3 VTAIL.t12 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X13 VDD2.t2 VN.t5 VTAIL.t4 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X14 VTAIL.t11 VP.t4 VDD1.t1 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=2.2473 ps=13.95 w=13.62 l=2.47
X15 VDD1.t0 VP.t5 VTAIL.t10 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=5.3118 ps=28.02 w=13.62 l=2.47
X16 VTAIL.t9 VP.t6 VDD1.t7 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X17 VDD1.t2 VP.t7 VTAIL.t8 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
X18 VTAIL.t1 VN.t6 VDD2.t1 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=5.3118 pd=28.02 as=2.2473 ps=13.95 w=13.62 l=2.47
X19 VTAIL.t0 VN.t7 VDD2.t0 w_n3770_n3692# sky130_fd_pr__pfet_01v8 ad=2.2473 pd=13.95 as=2.2473 ps=13.95 w=13.62 l=2.47
R0 VP.n16 VP.t4 166.523
R1 VP.n19 VP.n18 161.3
R2 VP.n20 VP.n15 161.3
R3 VP.n22 VP.n21 161.3
R4 VP.n23 VP.n14 161.3
R5 VP.n25 VP.n24 161.3
R6 VP.n27 VP.n26 161.3
R7 VP.n28 VP.n12 161.3
R8 VP.n30 VP.n29 161.3
R9 VP.n31 VP.n11 161.3
R10 VP.n33 VP.n32 161.3
R11 VP.n34 VP.n10 161.3
R12 VP.n64 VP.n0 161.3
R13 VP.n63 VP.n62 161.3
R14 VP.n61 VP.n1 161.3
R15 VP.n60 VP.n59 161.3
R16 VP.n58 VP.n2 161.3
R17 VP.n57 VP.n56 161.3
R18 VP.n55 VP.n54 161.3
R19 VP.n53 VP.n4 161.3
R20 VP.n52 VP.n51 161.3
R21 VP.n50 VP.n5 161.3
R22 VP.n49 VP.n48 161.3
R23 VP.n46 VP.n6 161.3
R24 VP.n45 VP.n44 161.3
R25 VP.n43 VP.n7 161.3
R26 VP.n42 VP.n41 161.3
R27 VP.n40 VP.n8 161.3
R28 VP.n39 VP.n38 161.3
R29 VP.n9 VP.t1 132.892
R30 VP.n47 VP.t7 132.892
R31 VP.n3 VP.t0 132.892
R32 VP.n65 VP.t2 132.892
R33 VP.n35 VP.t5 132.892
R34 VP.n13 VP.t6 132.892
R35 VP.n17 VP.t3 132.892
R36 VP.n37 VP.n9 101.072
R37 VP.n66 VP.n65 101.072
R38 VP.n36 VP.n35 101.072
R39 VP.n41 VP.n7 56.5617
R40 VP.n59 VP.n1 56.5617
R41 VP.n29 VP.n11 56.5617
R42 VP.n17 VP.n16 52.9956
R43 VP.n37 VP.n36 51.4997
R44 VP.n52 VP.n5 40.577
R45 VP.n53 VP.n52 40.577
R46 VP.n23 VP.n22 40.577
R47 VP.n22 VP.n15 40.577
R48 VP.n40 VP.n39 24.5923
R49 VP.n41 VP.n40 24.5923
R50 VP.n45 VP.n7 24.5923
R51 VP.n46 VP.n45 24.5923
R52 VP.n48 VP.n5 24.5923
R53 VP.n54 VP.n53 24.5923
R54 VP.n58 VP.n57 24.5923
R55 VP.n59 VP.n58 24.5923
R56 VP.n63 VP.n1 24.5923
R57 VP.n64 VP.n63 24.5923
R58 VP.n33 VP.n11 24.5923
R59 VP.n34 VP.n33 24.5923
R60 VP.n24 VP.n23 24.5923
R61 VP.n28 VP.n27 24.5923
R62 VP.n29 VP.n28 24.5923
R63 VP.n18 VP.n15 24.5923
R64 VP.n48 VP.n47 19.674
R65 VP.n54 VP.n3 19.674
R66 VP.n24 VP.n13 19.674
R67 VP.n18 VP.n17 19.674
R68 VP.n39 VP.n9 9.83723
R69 VP.n65 VP.n64 9.83723
R70 VP.n35 VP.n34 9.83723
R71 VP.n19 VP.n16 6.84375
R72 VP.n47 VP.n46 4.91887
R73 VP.n57 VP.n3 4.91887
R74 VP.n27 VP.n13 4.91887
R75 VP.n36 VP.n10 0.278335
R76 VP.n38 VP.n37 0.278335
R77 VP.n66 VP.n0 0.278335
R78 VP.n20 VP.n19 0.189894
R79 VP.n21 VP.n20 0.189894
R80 VP.n21 VP.n14 0.189894
R81 VP.n25 VP.n14 0.189894
R82 VP.n26 VP.n25 0.189894
R83 VP.n26 VP.n12 0.189894
R84 VP.n30 VP.n12 0.189894
R85 VP.n31 VP.n30 0.189894
R86 VP.n32 VP.n31 0.189894
R87 VP.n32 VP.n10 0.189894
R88 VP.n38 VP.n8 0.189894
R89 VP.n42 VP.n8 0.189894
R90 VP.n43 VP.n42 0.189894
R91 VP.n44 VP.n43 0.189894
R92 VP.n44 VP.n6 0.189894
R93 VP.n49 VP.n6 0.189894
R94 VP.n50 VP.n49 0.189894
R95 VP.n51 VP.n50 0.189894
R96 VP.n51 VP.n4 0.189894
R97 VP.n55 VP.n4 0.189894
R98 VP.n56 VP.n55 0.189894
R99 VP.n56 VP.n2 0.189894
R100 VP.n60 VP.n2 0.189894
R101 VP.n61 VP.n60 0.189894
R102 VP.n62 VP.n61 0.189894
R103 VP.n62 VP.n0 0.189894
R104 VP VP.n66 0.153485
R105 VDD1 VDD1.n0 74.0718
R106 VDD1.n3 VDD1.n2 73.958
R107 VDD1.n3 VDD1.n1 73.958
R108 VDD1.n5 VDD1.n4 72.8065
R109 VDD1.n5 VDD1.n3 46.9018
R110 VDD1.n4 VDD1.t7 2.38706
R111 VDD1.n4 VDD1.t0 2.38706
R112 VDD1.n0 VDD1.t1 2.38706
R113 VDD1.n0 VDD1.t4 2.38706
R114 VDD1.n2 VDD1.t3 2.38706
R115 VDD1.n2 VDD1.t5 2.38706
R116 VDD1.n1 VDD1.t6 2.38706
R117 VDD1.n1 VDD1.t2 2.38706
R118 VDD1 VDD1.n5 1.14921
R119 VTAIL.n11 VTAIL.t11 58.5144
R120 VTAIL.n10 VTAIL.t6 58.5144
R121 VTAIL.n7 VTAIL.t1 58.5144
R122 VTAIL.n15 VTAIL.t3 58.5142
R123 VTAIL.n2 VTAIL.t7 58.5142
R124 VTAIL.n3 VTAIL.t13 58.5142
R125 VTAIL.n6 VTAIL.t14 58.5142
R126 VTAIL.n14 VTAIL.t10 58.5142
R127 VTAIL.n13 VTAIL.n12 56.1279
R128 VTAIL.n9 VTAIL.n8 56.1279
R129 VTAIL.n1 VTAIL.n0 56.1277
R130 VTAIL.n5 VTAIL.n4 56.1277
R131 VTAIL.n15 VTAIL.n14 26.5221
R132 VTAIL.n7 VTAIL.n6 26.5221
R133 VTAIL.n9 VTAIL.n7 2.41429
R134 VTAIL.n10 VTAIL.n9 2.41429
R135 VTAIL.n13 VTAIL.n11 2.41429
R136 VTAIL.n14 VTAIL.n13 2.41429
R137 VTAIL.n6 VTAIL.n5 2.41429
R138 VTAIL.n5 VTAIL.n3 2.41429
R139 VTAIL.n2 VTAIL.n1 2.41429
R140 VTAIL.n0 VTAIL.t5 2.38706
R141 VTAIL.n0 VTAIL.t0 2.38706
R142 VTAIL.n4 VTAIL.t8 2.38706
R143 VTAIL.n4 VTAIL.t15 2.38706
R144 VTAIL.n12 VTAIL.t12 2.38706
R145 VTAIL.n12 VTAIL.t9 2.38706
R146 VTAIL.n8 VTAIL.t4 2.38706
R147 VTAIL.n8 VTAIL.t2 2.38706
R148 VTAIL VTAIL.n15 2.3561
R149 VTAIL.n11 VTAIL.n10 0.470328
R150 VTAIL.n3 VTAIL.n2 0.470328
R151 VTAIL VTAIL.n1 0.0586897
R152 B.n438 B.n437 585
R153 B.n436 B.n133 585
R154 B.n435 B.n434 585
R155 B.n433 B.n134 585
R156 B.n432 B.n431 585
R157 B.n430 B.n135 585
R158 B.n429 B.n428 585
R159 B.n427 B.n136 585
R160 B.n426 B.n425 585
R161 B.n424 B.n137 585
R162 B.n423 B.n422 585
R163 B.n421 B.n138 585
R164 B.n420 B.n419 585
R165 B.n418 B.n139 585
R166 B.n417 B.n416 585
R167 B.n415 B.n140 585
R168 B.n414 B.n413 585
R169 B.n412 B.n141 585
R170 B.n411 B.n410 585
R171 B.n409 B.n142 585
R172 B.n408 B.n407 585
R173 B.n406 B.n143 585
R174 B.n405 B.n404 585
R175 B.n403 B.n144 585
R176 B.n402 B.n401 585
R177 B.n400 B.n145 585
R178 B.n399 B.n398 585
R179 B.n397 B.n146 585
R180 B.n396 B.n395 585
R181 B.n394 B.n147 585
R182 B.n393 B.n392 585
R183 B.n391 B.n148 585
R184 B.n390 B.n389 585
R185 B.n388 B.n149 585
R186 B.n387 B.n386 585
R187 B.n385 B.n150 585
R188 B.n384 B.n383 585
R189 B.n382 B.n151 585
R190 B.n381 B.n380 585
R191 B.n379 B.n152 585
R192 B.n378 B.n377 585
R193 B.n376 B.n153 585
R194 B.n375 B.n374 585
R195 B.n373 B.n154 585
R196 B.n372 B.n371 585
R197 B.n370 B.n155 585
R198 B.n369 B.n368 585
R199 B.n364 B.n156 585
R200 B.n363 B.n362 585
R201 B.n361 B.n157 585
R202 B.n360 B.n359 585
R203 B.n358 B.n158 585
R204 B.n357 B.n356 585
R205 B.n355 B.n159 585
R206 B.n354 B.n353 585
R207 B.n352 B.n160 585
R208 B.n350 B.n349 585
R209 B.n348 B.n163 585
R210 B.n347 B.n346 585
R211 B.n345 B.n164 585
R212 B.n344 B.n343 585
R213 B.n342 B.n165 585
R214 B.n341 B.n340 585
R215 B.n339 B.n166 585
R216 B.n338 B.n337 585
R217 B.n336 B.n167 585
R218 B.n335 B.n334 585
R219 B.n333 B.n168 585
R220 B.n332 B.n331 585
R221 B.n330 B.n169 585
R222 B.n329 B.n328 585
R223 B.n327 B.n170 585
R224 B.n326 B.n325 585
R225 B.n324 B.n171 585
R226 B.n323 B.n322 585
R227 B.n321 B.n172 585
R228 B.n320 B.n319 585
R229 B.n318 B.n173 585
R230 B.n317 B.n316 585
R231 B.n315 B.n174 585
R232 B.n314 B.n313 585
R233 B.n312 B.n175 585
R234 B.n311 B.n310 585
R235 B.n309 B.n176 585
R236 B.n308 B.n307 585
R237 B.n306 B.n177 585
R238 B.n305 B.n304 585
R239 B.n303 B.n178 585
R240 B.n302 B.n301 585
R241 B.n300 B.n179 585
R242 B.n299 B.n298 585
R243 B.n297 B.n180 585
R244 B.n296 B.n295 585
R245 B.n294 B.n181 585
R246 B.n293 B.n292 585
R247 B.n291 B.n182 585
R248 B.n290 B.n289 585
R249 B.n288 B.n183 585
R250 B.n287 B.n286 585
R251 B.n285 B.n184 585
R252 B.n284 B.n283 585
R253 B.n282 B.n185 585
R254 B.n439 B.n132 585
R255 B.n441 B.n440 585
R256 B.n442 B.n131 585
R257 B.n444 B.n443 585
R258 B.n445 B.n130 585
R259 B.n447 B.n446 585
R260 B.n448 B.n129 585
R261 B.n450 B.n449 585
R262 B.n451 B.n128 585
R263 B.n453 B.n452 585
R264 B.n454 B.n127 585
R265 B.n456 B.n455 585
R266 B.n457 B.n126 585
R267 B.n459 B.n458 585
R268 B.n460 B.n125 585
R269 B.n462 B.n461 585
R270 B.n463 B.n124 585
R271 B.n465 B.n464 585
R272 B.n466 B.n123 585
R273 B.n468 B.n467 585
R274 B.n469 B.n122 585
R275 B.n471 B.n470 585
R276 B.n472 B.n121 585
R277 B.n474 B.n473 585
R278 B.n475 B.n120 585
R279 B.n477 B.n476 585
R280 B.n478 B.n119 585
R281 B.n480 B.n479 585
R282 B.n481 B.n118 585
R283 B.n483 B.n482 585
R284 B.n484 B.n117 585
R285 B.n486 B.n485 585
R286 B.n487 B.n116 585
R287 B.n489 B.n488 585
R288 B.n490 B.n115 585
R289 B.n492 B.n491 585
R290 B.n493 B.n114 585
R291 B.n495 B.n494 585
R292 B.n496 B.n113 585
R293 B.n498 B.n497 585
R294 B.n499 B.n112 585
R295 B.n501 B.n500 585
R296 B.n502 B.n111 585
R297 B.n504 B.n503 585
R298 B.n505 B.n110 585
R299 B.n507 B.n506 585
R300 B.n508 B.n109 585
R301 B.n510 B.n509 585
R302 B.n511 B.n108 585
R303 B.n513 B.n512 585
R304 B.n514 B.n107 585
R305 B.n516 B.n515 585
R306 B.n517 B.n106 585
R307 B.n519 B.n518 585
R308 B.n520 B.n105 585
R309 B.n522 B.n521 585
R310 B.n523 B.n104 585
R311 B.n525 B.n524 585
R312 B.n526 B.n103 585
R313 B.n528 B.n527 585
R314 B.n529 B.n102 585
R315 B.n531 B.n530 585
R316 B.n532 B.n101 585
R317 B.n534 B.n533 585
R318 B.n535 B.n100 585
R319 B.n537 B.n536 585
R320 B.n538 B.n99 585
R321 B.n540 B.n539 585
R322 B.n541 B.n98 585
R323 B.n543 B.n542 585
R324 B.n544 B.n97 585
R325 B.n546 B.n545 585
R326 B.n547 B.n96 585
R327 B.n549 B.n548 585
R328 B.n550 B.n95 585
R329 B.n552 B.n551 585
R330 B.n553 B.n94 585
R331 B.n555 B.n554 585
R332 B.n556 B.n93 585
R333 B.n558 B.n557 585
R334 B.n559 B.n92 585
R335 B.n561 B.n560 585
R336 B.n562 B.n91 585
R337 B.n564 B.n563 585
R338 B.n565 B.n90 585
R339 B.n567 B.n566 585
R340 B.n568 B.n89 585
R341 B.n570 B.n569 585
R342 B.n571 B.n88 585
R343 B.n573 B.n572 585
R344 B.n574 B.n87 585
R345 B.n576 B.n575 585
R346 B.n577 B.n86 585
R347 B.n579 B.n578 585
R348 B.n580 B.n85 585
R349 B.n582 B.n581 585
R350 B.n583 B.n84 585
R351 B.n585 B.n584 585
R352 B.n586 B.n83 585
R353 B.n588 B.n587 585
R354 B.n742 B.n741 585
R355 B.n740 B.n27 585
R356 B.n739 B.n738 585
R357 B.n737 B.n28 585
R358 B.n736 B.n735 585
R359 B.n734 B.n29 585
R360 B.n733 B.n732 585
R361 B.n731 B.n30 585
R362 B.n730 B.n729 585
R363 B.n728 B.n31 585
R364 B.n727 B.n726 585
R365 B.n725 B.n32 585
R366 B.n724 B.n723 585
R367 B.n722 B.n33 585
R368 B.n721 B.n720 585
R369 B.n719 B.n34 585
R370 B.n718 B.n717 585
R371 B.n716 B.n35 585
R372 B.n715 B.n714 585
R373 B.n713 B.n36 585
R374 B.n712 B.n711 585
R375 B.n710 B.n37 585
R376 B.n709 B.n708 585
R377 B.n707 B.n38 585
R378 B.n706 B.n705 585
R379 B.n704 B.n39 585
R380 B.n703 B.n702 585
R381 B.n701 B.n40 585
R382 B.n700 B.n699 585
R383 B.n698 B.n41 585
R384 B.n697 B.n696 585
R385 B.n695 B.n42 585
R386 B.n694 B.n693 585
R387 B.n692 B.n43 585
R388 B.n691 B.n690 585
R389 B.n689 B.n44 585
R390 B.n688 B.n687 585
R391 B.n686 B.n45 585
R392 B.n685 B.n684 585
R393 B.n683 B.n46 585
R394 B.n682 B.n681 585
R395 B.n680 B.n47 585
R396 B.n679 B.n678 585
R397 B.n677 B.n48 585
R398 B.n676 B.n675 585
R399 B.n674 B.n49 585
R400 B.n672 B.n671 585
R401 B.n670 B.n52 585
R402 B.n669 B.n668 585
R403 B.n667 B.n53 585
R404 B.n666 B.n665 585
R405 B.n664 B.n54 585
R406 B.n663 B.n662 585
R407 B.n661 B.n55 585
R408 B.n660 B.n659 585
R409 B.n658 B.n56 585
R410 B.n657 B.n656 585
R411 B.n655 B.n57 585
R412 B.n654 B.n653 585
R413 B.n652 B.n61 585
R414 B.n651 B.n650 585
R415 B.n649 B.n62 585
R416 B.n648 B.n647 585
R417 B.n646 B.n63 585
R418 B.n645 B.n644 585
R419 B.n643 B.n64 585
R420 B.n642 B.n641 585
R421 B.n640 B.n65 585
R422 B.n639 B.n638 585
R423 B.n637 B.n66 585
R424 B.n636 B.n635 585
R425 B.n634 B.n67 585
R426 B.n633 B.n632 585
R427 B.n631 B.n68 585
R428 B.n630 B.n629 585
R429 B.n628 B.n69 585
R430 B.n627 B.n626 585
R431 B.n625 B.n70 585
R432 B.n624 B.n623 585
R433 B.n622 B.n71 585
R434 B.n621 B.n620 585
R435 B.n619 B.n72 585
R436 B.n618 B.n617 585
R437 B.n616 B.n73 585
R438 B.n615 B.n614 585
R439 B.n613 B.n74 585
R440 B.n612 B.n611 585
R441 B.n610 B.n75 585
R442 B.n609 B.n608 585
R443 B.n607 B.n76 585
R444 B.n606 B.n605 585
R445 B.n604 B.n77 585
R446 B.n603 B.n602 585
R447 B.n601 B.n78 585
R448 B.n600 B.n599 585
R449 B.n598 B.n79 585
R450 B.n597 B.n596 585
R451 B.n595 B.n80 585
R452 B.n594 B.n593 585
R453 B.n592 B.n81 585
R454 B.n591 B.n590 585
R455 B.n589 B.n82 585
R456 B.n743 B.n26 585
R457 B.n745 B.n744 585
R458 B.n746 B.n25 585
R459 B.n748 B.n747 585
R460 B.n749 B.n24 585
R461 B.n751 B.n750 585
R462 B.n752 B.n23 585
R463 B.n754 B.n753 585
R464 B.n755 B.n22 585
R465 B.n757 B.n756 585
R466 B.n758 B.n21 585
R467 B.n760 B.n759 585
R468 B.n761 B.n20 585
R469 B.n763 B.n762 585
R470 B.n764 B.n19 585
R471 B.n766 B.n765 585
R472 B.n767 B.n18 585
R473 B.n769 B.n768 585
R474 B.n770 B.n17 585
R475 B.n772 B.n771 585
R476 B.n773 B.n16 585
R477 B.n775 B.n774 585
R478 B.n776 B.n15 585
R479 B.n778 B.n777 585
R480 B.n779 B.n14 585
R481 B.n781 B.n780 585
R482 B.n782 B.n13 585
R483 B.n784 B.n783 585
R484 B.n785 B.n12 585
R485 B.n787 B.n786 585
R486 B.n788 B.n11 585
R487 B.n790 B.n789 585
R488 B.n791 B.n10 585
R489 B.n793 B.n792 585
R490 B.n794 B.n9 585
R491 B.n796 B.n795 585
R492 B.n797 B.n8 585
R493 B.n799 B.n798 585
R494 B.n800 B.n7 585
R495 B.n802 B.n801 585
R496 B.n803 B.n6 585
R497 B.n805 B.n804 585
R498 B.n806 B.n5 585
R499 B.n808 B.n807 585
R500 B.n809 B.n4 585
R501 B.n811 B.n810 585
R502 B.n812 B.n3 585
R503 B.n814 B.n813 585
R504 B.n815 B.n0 585
R505 B.n2 B.n1 585
R506 B.n210 B.n209 585
R507 B.n212 B.n211 585
R508 B.n213 B.n208 585
R509 B.n215 B.n214 585
R510 B.n216 B.n207 585
R511 B.n218 B.n217 585
R512 B.n219 B.n206 585
R513 B.n221 B.n220 585
R514 B.n222 B.n205 585
R515 B.n224 B.n223 585
R516 B.n225 B.n204 585
R517 B.n227 B.n226 585
R518 B.n228 B.n203 585
R519 B.n230 B.n229 585
R520 B.n231 B.n202 585
R521 B.n233 B.n232 585
R522 B.n234 B.n201 585
R523 B.n236 B.n235 585
R524 B.n237 B.n200 585
R525 B.n239 B.n238 585
R526 B.n240 B.n199 585
R527 B.n242 B.n241 585
R528 B.n243 B.n198 585
R529 B.n245 B.n244 585
R530 B.n246 B.n197 585
R531 B.n248 B.n247 585
R532 B.n249 B.n196 585
R533 B.n251 B.n250 585
R534 B.n252 B.n195 585
R535 B.n254 B.n253 585
R536 B.n255 B.n194 585
R537 B.n257 B.n256 585
R538 B.n258 B.n193 585
R539 B.n260 B.n259 585
R540 B.n261 B.n192 585
R541 B.n263 B.n262 585
R542 B.n264 B.n191 585
R543 B.n266 B.n265 585
R544 B.n267 B.n190 585
R545 B.n269 B.n268 585
R546 B.n270 B.n189 585
R547 B.n272 B.n271 585
R548 B.n273 B.n188 585
R549 B.n275 B.n274 585
R550 B.n276 B.n187 585
R551 B.n278 B.n277 585
R552 B.n279 B.n186 585
R553 B.n281 B.n280 585
R554 B.n282 B.n281 492.5
R555 B.n437 B.n132 492.5
R556 B.n587 B.n82 492.5
R557 B.n743 B.n742 492.5
R558 B.n161 B.t9 340.733
R559 B.n365 B.t6 340.733
R560 B.n58 B.t0 340.733
R561 B.n50 B.t3 340.733
R562 B.n817 B.n816 256.663
R563 B.n816 B.n815 235.042
R564 B.n816 B.n2 235.042
R565 B.n283 B.n282 163.367
R566 B.n283 B.n184 163.367
R567 B.n287 B.n184 163.367
R568 B.n288 B.n287 163.367
R569 B.n289 B.n288 163.367
R570 B.n289 B.n182 163.367
R571 B.n293 B.n182 163.367
R572 B.n294 B.n293 163.367
R573 B.n295 B.n294 163.367
R574 B.n295 B.n180 163.367
R575 B.n299 B.n180 163.367
R576 B.n300 B.n299 163.367
R577 B.n301 B.n300 163.367
R578 B.n301 B.n178 163.367
R579 B.n305 B.n178 163.367
R580 B.n306 B.n305 163.367
R581 B.n307 B.n306 163.367
R582 B.n307 B.n176 163.367
R583 B.n311 B.n176 163.367
R584 B.n312 B.n311 163.367
R585 B.n313 B.n312 163.367
R586 B.n313 B.n174 163.367
R587 B.n317 B.n174 163.367
R588 B.n318 B.n317 163.367
R589 B.n319 B.n318 163.367
R590 B.n319 B.n172 163.367
R591 B.n323 B.n172 163.367
R592 B.n324 B.n323 163.367
R593 B.n325 B.n324 163.367
R594 B.n325 B.n170 163.367
R595 B.n329 B.n170 163.367
R596 B.n330 B.n329 163.367
R597 B.n331 B.n330 163.367
R598 B.n331 B.n168 163.367
R599 B.n335 B.n168 163.367
R600 B.n336 B.n335 163.367
R601 B.n337 B.n336 163.367
R602 B.n337 B.n166 163.367
R603 B.n341 B.n166 163.367
R604 B.n342 B.n341 163.367
R605 B.n343 B.n342 163.367
R606 B.n343 B.n164 163.367
R607 B.n347 B.n164 163.367
R608 B.n348 B.n347 163.367
R609 B.n349 B.n348 163.367
R610 B.n349 B.n160 163.367
R611 B.n354 B.n160 163.367
R612 B.n355 B.n354 163.367
R613 B.n356 B.n355 163.367
R614 B.n356 B.n158 163.367
R615 B.n360 B.n158 163.367
R616 B.n361 B.n360 163.367
R617 B.n362 B.n361 163.367
R618 B.n362 B.n156 163.367
R619 B.n369 B.n156 163.367
R620 B.n370 B.n369 163.367
R621 B.n371 B.n370 163.367
R622 B.n371 B.n154 163.367
R623 B.n375 B.n154 163.367
R624 B.n376 B.n375 163.367
R625 B.n377 B.n376 163.367
R626 B.n377 B.n152 163.367
R627 B.n381 B.n152 163.367
R628 B.n382 B.n381 163.367
R629 B.n383 B.n382 163.367
R630 B.n383 B.n150 163.367
R631 B.n387 B.n150 163.367
R632 B.n388 B.n387 163.367
R633 B.n389 B.n388 163.367
R634 B.n389 B.n148 163.367
R635 B.n393 B.n148 163.367
R636 B.n394 B.n393 163.367
R637 B.n395 B.n394 163.367
R638 B.n395 B.n146 163.367
R639 B.n399 B.n146 163.367
R640 B.n400 B.n399 163.367
R641 B.n401 B.n400 163.367
R642 B.n401 B.n144 163.367
R643 B.n405 B.n144 163.367
R644 B.n406 B.n405 163.367
R645 B.n407 B.n406 163.367
R646 B.n407 B.n142 163.367
R647 B.n411 B.n142 163.367
R648 B.n412 B.n411 163.367
R649 B.n413 B.n412 163.367
R650 B.n413 B.n140 163.367
R651 B.n417 B.n140 163.367
R652 B.n418 B.n417 163.367
R653 B.n419 B.n418 163.367
R654 B.n419 B.n138 163.367
R655 B.n423 B.n138 163.367
R656 B.n424 B.n423 163.367
R657 B.n425 B.n424 163.367
R658 B.n425 B.n136 163.367
R659 B.n429 B.n136 163.367
R660 B.n430 B.n429 163.367
R661 B.n431 B.n430 163.367
R662 B.n431 B.n134 163.367
R663 B.n435 B.n134 163.367
R664 B.n436 B.n435 163.367
R665 B.n437 B.n436 163.367
R666 B.n587 B.n586 163.367
R667 B.n586 B.n585 163.367
R668 B.n585 B.n84 163.367
R669 B.n581 B.n84 163.367
R670 B.n581 B.n580 163.367
R671 B.n580 B.n579 163.367
R672 B.n579 B.n86 163.367
R673 B.n575 B.n86 163.367
R674 B.n575 B.n574 163.367
R675 B.n574 B.n573 163.367
R676 B.n573 B.n88 163.367
R677 B.n569 B.n88 163.367
R678 B.n569 B.n568 163.367
R679 B.n568 B.n567 163.367
R680 B.n567 B.n90 163.367
R681 B.n563 B.n90 163.367
R682 B.n563 B.n562 163.367
R683 B.n562 B.n561 163.367
R684 B.n561 B.n92 163.367
R685 B.n557 B.n92 163.367
R686 B.n557 B.n556 163.367
R687 B.n556 B.n555 163.367
R688 B.n555 B.n94 163.367
R689 B.n551 B.n94 163.367
R690 B.n551 B.n550 163.367
R691 B.n550 B.n549 163.367
R692 B.n549 B.n96 163.367
R693 B.n545 B.n96 163.367
R694 B.n545 B.n544 163.367
R695 B.n544 B.n543 163.367
R696 B.n543 B.n98 163.367
R697 B.n539 B.n98 163.367
R698 B.n539 B.n538 163.367
R699 B.n538 B.n537 163.367
R700 B.n537 B.n100 163.367
R701 B.n533 B.n100 163.367
R702 B.n533 B.n532 163.367
R703 B.n532 B.n531 163.367
R704 B.n531 B.n102 163.367
R705 B.n527 B.n102 163.367
R706 B.n527 B.n526 163.367
R707 B.n526 B.n525 163.367
R708 B.n525 B.n104 163.367
R709 B.n521 B.n104 163.367
R710 B.n521 B.n520 163.367
R711 B.n520 B.n519 163.367
R712 B.n519 B.n106 163.367
R713 B.n515 B.n106 163.367
R714 B.n515 B.n514 163.367
R715 B.n514 B.n513 163.367
R716 B.n513 B.n108 163.367
R717 B.n509 B.n108 163.367
R718 B.n509 B.n508 163.367
R719 B.n508 B.n507 163.367
R720 B.n507 B.n110 163.367
R721 B.n503 B.n110 163.367
R722 B.n503 B.n502 163.367
R723 B.n502 B.n501 163.367
R724 B.n501 B.n112 163.367
R725 B.n497 B.n112 163.367
R726 B.n497 B.n496 163.367
R727 B.n496 B.n495 163.367
R728 B.n495 B.n114 163.367
R729 B.n491 B.n114 163.367
R730 B.n491 B.n490 163.367
R731 B.n490 B.n489 163.367
R732 B.n489 B.n116 163.367
R733 B.n485 B.n116 163.367
R734 B.n485 B.n484 163.367
R735 B.n484 B.n483 163.367
R736 B.n483 B.n118 163.367
R737 B.n479 B.n118 163.367
R738 B.n479 B.n478 163.367
R739 B.n478 B.n477 163.367
R740 B.n477 B.n120 163.367
R741 B.n473 B.n120 163.367
R742 B.n473 B.n472 163.367
R743 B.n472 B.n471 163.367
R744 B.n471 B.n122 163.367
R745 B.n467 B.n122 163.367
R746 B.n467 B.n466 163.367
R747 B.n466 B.n465 163.367
R748 B.n465 B.n124 163.367
R749 B.n461 B.n124 163.367
R750 B.n461 B.n460 163.367
R751 B.n460 B.n459 163.367
R752 B.n459 B.n126 163.367
R753 B.n455 B.n126 163.367
R754 B.n455 B.n454 163.367
R755 B.n454 B.n453 163.367
R756 B.n453 B.n128 163.367
R757 B.n449 B.n128 163.367
R758 B.n449 B.n448 163.367
R759 B.n448 B.n447 163.367
R760 B.n447 B.n130 163.367
R761 B.n443 B.n130 163.367
R762 B.n443 B.n442 163.367
R763 B.n442 B.n441 163.367
R764 B.n441 B.n132 163.367
R765 B.n742 B.n27 163.367
R766 B.n738 B.n27 163.367
R767 B.n738 B.n737 163.367
R768 B.n737 B.n736 163.367
R769 B.n736 B.n29 163.367
R770 B.n732 B.n29 163.367
R771 B.n732 B.n731 163.367
R772 B.n731 B.n730 163.367
R773 B.n730 B.n31 163.367
R774 B.n726 B.n31 163.367
R775 B.n726 B.n725 163.367
R776 B.n725 B.n724 163.367
R777 B.n724 B.n33 163.367
R778 B.n720 B.n33 163.367
R779 B.n720 B.n719 163.367
R780 B.n719 B.n718 163.367
R781 B.n718 B.n35 163.367
R782 B.n714 B.n35 163.367
R783 B.n714 B.n713 163.367
R784 B.n713 B.n712 163.367
R785 B.n712 B.n37 163.367
R786 B.n708 B.n37 163.367
R787 B.n708 B.n707 163.367
R788 B.n707 B.n706 163.367
R789 B.n706 B.n39 163.367
R790 B.n702 B.n39 163.367
R791 B.n702 B.n701 163.367
R792 B.n701 B.n700 163.367
R793 B.n700 B.n41 163.367
R794 B.n696 B.n41 163.367
R795 B.n696 B.n695 163.367
R796 B.n695 B.n694 163.367
R797 B.n694 B.n43 163.367
R798 B.n690 B.n43 163.367
R799 B.n690 B.n689 163.367
R800 B.n689 B.n688 163.367
R801 B.n688 B.n45 163.367
R802 B.n684 B.n45 163.367
R803 B.n684 B.n683 163.367
R804 B.n683 B.n682 163.367
R805 B.n682 B.n47 163.367
R806 B.n678 B.n47 163.367
R807 B.n678 B.n677 163.367
R808 B.n677 B.n676 163.367
R809 B.n676 B.n49 163.367
R810 B.n671 B.n49 163.367
R811 B.n671 B.n670 163.367
R812 B.n670 B.n669 163.367
R813 B.n669 B.n53 163.367
R814 B.n665 B.n53 163.367
R815 B.n665 B.n664 163.367
R816 B.n664 B.n663 163.367
R817 B.n663 B.n55 163.367
R818 B.n659 B.n55 163.367
R819 B.n659 B.n658 163.367
R820 B.n658 B.n657 163.367
R821 B.n657 B.n57 163.367
R822 B.n653 B.n57 163.367
R823 B.n653 B.n652 163.367
R824 B.n652 B.n651 163.367
R825 B.n651 B.n62 163.367
R826 B.n647 B.n62 163.367
R827 B.n647 B.n646 163.367
R828 B.n646 B.n645 163.367
R829 B.n645 B.n64 163.367
R830 B.n641 B.n64 163.367
R831 B.n641 B.n640 163.367
R832 B.n640 B.n639 163.367
R833 B.n639 B.n66 163.367
R834 B.n635 B.n66 163.367
R835 B.n635 B.n634 163.367
R836 B.n634 B.n633 163.367
R837 B.n633 B.n68 163.367
R838 B.n629 B.n68 163.367
R839 B.n629 B.n628 163.367
R840 B.n628 B.n627 163.367
R841 B.n627 B.n70 163.367
R842 B.n623 B.n70 163.367
R843 B.n623 B.n622 163.367
R844 B.n622 B.n621 163.367
R845 B.n621 B.n72 163.367
R846 B.n617 B.n72 163.367
R847 B.n617 B.n616 163.367
R848 B.n616 B.n615 163.367
R849 B.n615 B.n74 163.367
R850 B.n611 B.n74 163.367
R851 B.n611 B.n610 163.367
R852 B.n610 B.n609 163.367
R853 B.n609 B.n76 163.367
R854 B.n605 B.n76 163.367
R855 B.n605 B.n604 163.367
R856 B.n604 B.n603 163.367
R857 B.n603 B.n78 163.367
R858 B.n599 B.n78 163.367
R859 B.n599 B.n598 163.367
R860 B.n598 B.n597 163.367
R861 B.n597 B.n80 163.367
R862 B.n593 B.n80 163.367
R863 B.n593 B.n592 163.367
R864 B.n592 B.n591 163.367
R865 B.n591 B.n82 163.367
R866 B.n744 B.n743 163.367
R867 B.n744 B.n25 163.367
R868 B.n748 B.n25 163.367
R869 B.n749 B.n748 163.367
R870 B.n750 B.n749 163.367
R871 B.n750 B.n23 163.367
R872 B.n754 B.n23 163.367
R873 B.n755 B.n754 163.367
R874 B.n756 B.n755 163.367
R875 B.n756 B.n21 163.367
R876 B.n760 B.n21 163.367
R877 B.n761 B.n760 163.367
R878 B.n762 B.n761 163.367
R879 B.n762 B.n19 163.367
R880 B.n766 B.n19 163.367
R881 B.n767 B.n766 163.367
R882 B.n768 B.n767 163.367
R883 B.n768 B.n17 163.367
R884 B.n772 B.n17 163.367
R885 B.n773 B.n772 163.367
R886 B.n774 B.n773 163.367
R887 B.n774 B.n15 163.367
R888 B.n778 B.n15 163.367
R889 B.n779 B.n778 163.367
R890 B.n780 B.n779 163.367
R891 B.n780 B.n13 163.367
R892 B.n784 B.n13 163.367
R893 B.n785 B.n784 163.367
R894 B.n786 B.n785 163.367
R895 B.n786 B.n11 163.367
R896 B.n790 B.n11 163.367
R897 B.n791 B.n790 163.367
R898 B.n792 B.n791 163.367
R899 B.n792 B.n9 163.367
R900 B.n796 B.n9 163.367
R901 B.n797 B.n796 163.367
R902 B.n798 B.n797 163.367
R903 B.n798 B.n7 163.367
R904 B.n802 B.n7 163.367
R905 B.n803 B.n802 163.367
R906 B.n804 B.n803 163.367
R907 B.n804 B.n5 163.367
R908 B.n808 B.n5 163.367
R909 B.n809 B.n808 163.367
R910 B.n810 B.n809 163.367
R911 B.n810 B.n3 163.367
R912 B.n814 B.n3 163.367
R913 B.n815 B.n814 163.367
R914 B.n210 B.n2 163.367
R915 B.n211 B.n210 163.367
R916 B.n211 B.n208 163.367
R917 B.n215 B.n208 163.367
R918 B.n216 B.n215 163.367
R919 B.n217 B.n216 163.367
R920 B.n217 B.n206 163.367
R921 B.n221 B.n206 163.367
R922 B.n222 B.n221 163.367
R923 B.n223 B.n222 163.367
R924 B.n223 B.n204 163.367
R925 B.n227 B.n204 163.367
R926 B.n228 B.n227 163.367
R927 B.n229 B.n228 163.367
R928 B.n229 B.n202 163.367
R929 B.n233 B.n202 163.367
R930 B.n234 B.n233 163.367
R931 B.n235 B.n234 163.367
R932 B.n235 B.n200 163.367
R933 B.n239 B.n200 163.367
R934 B.n240 B.n239 163.367
R935 B.n241 B.n240 163.367
R936 B.n241 B.n198 163.367
R937 B.n245 B.n198 163.367
R938 B.n246 B.n245 163.367
R939 B.n247 B.n246 163.367
R940 B.n247 B.n196 163.367
R941 B.n251 B.n196 163.367
R942 B.n252 B.n251 163.367
R943 B.n253 B.n252 163.367
R944 B.n253 B.n194 163.367
R945 B.n257 B.n194 163.367
R946 B.n258 B.n257 163.367
R947 B.n259 B.n258 163.367
R948 B.n259 B.n192 163.367
R949 B.n263 B.n192 163.367
R950 B.n264 B.n263 163.367
R951 B.n265 B.n264 163.367
R952 B.n265 B.n190 163.367
R953 B.n269 B.n190 163.367
R954 B.n270 B.n269 163.367
R955 B.n271 B.n270 163.367
R956 B.n271 B.n188 163.367
R957 B.n275 B.n188 163.367
R958 B.n276 B.n275 163.367
R959 B.n277 B.n276 163.367
R960 B.n277 B.n186 163.367
R961 B.n281 B.n186 163.367
R962 B.n365 B.t7 161.47
R963 B.n58 B.t2 161.47
R964 B.n161 B.t10 161.453
R965 B.n50 B.t5 161.453
R966 B.n366 B.t8 107.168
R967 B.n59 B.t1 107.168
R968 B.n162 B.t11 107.15
R969 B.n51 B.t4 107.15
R970 B.n351 B.n162 59.5399
R971 B.n367 B.n366 59.5399
R972 B.n60 B.n59 59.5399
R973 B.n673 B.n51 59.5399
R974 B.n162 B.n161 54.3035
R975 B.n366 B.n365 54.3035
R976 B.n59 B.n58 54.3035
R977 B.n51 B.n50 54.3035
R978 B.n741 B.n26 32.0005
R979 B.n589 B.n588 32.0005
R980 B.n439 B.n438 32.0005
R981 B.n280 B.n185 32.0005
R982 B B.n817 18.0485
R983 B.n745 B.n26 10.6151
R984 B.n746 B.n745 10.6151
R985 B.n747 B.n746 10.6151
R986 B.n747 B.n24 10.6151
R987 B.n751 B.n24 10.6151
R988 B.n752 B.n751 10.6151
R989 B.n753 B.n752 10.6151
R990 B.n753 B.n22 10.6151
R991 B.n757 B.n22 10.6151
R992 B.n758 B.n757 10.6151
R993 B.n759 B.n758 10.6151
R994 B.n759 B.n20 10.6151
R995 B.n763 B.n20 10.6151
R996 B.n764 B.n763 10.6151
R997 B.n765 B.n764 10.6151
R998 B.n765 B.n18 10.6151
R999 B.n769 B.n18 10.6151
R1000 B.n770 B.n769 10.6151
R1001 B.n771 B.n770 10.6151
R1002 B.n771 B.n16 10.6151
R1003 B.n775 B.n16 10.6151
R1004 B.n776 B.n775 10.6151
R1005 B.n777 B.n776 10.6151
R1006 B.n777 B.n14 10.6151
R1007 B.n781 B.n14 10.6151
R1008 B.n782 B.n781 10.6151
R1009 B.n783 B.n782 10.6151
R1010 B.n783 B.n12 10.6151
R1011 B.n787 B.n12 10.6151
R1012 B.n788 B.n787 10.6151
R1013 B.n789 B.n788 10.6151
R1014 B.n789 B.n10 10.6151
R1015 B.n793 B.n10 10.6151
R1016 B.n794 B.n793 10.6151
R1017 B.n795 B.n794 10.6151
R1018 B.n795 B.n8 10.6151
R1019 B.n799 B.n8 10.6151
R1020 B.n800 B.n799 10.6151
R1021 B.n801 B.n800 10.6151
R1022 B.n801 B.n6 10.6151
R1023 B.n805 B.n6 10.6151
R1024 B.n806 B.n805 10.6151
R1025 B.n807 B.n806 10.6151
R1026 B.n807 B.n4 10.6151
R1027 B.n811 B.n4 10.6151
R1028 B.n812 B.n811 10.6151
R1029 B.n813 B.n812 10.6151
R1030 B.n813 B.n0 10.6151
R1031 B.n741 B.n740 10.6151
R1032 B.n740 B.n739 10.6151
R1033 B.n739 B.n28 10.6151
R1034 B.n735 B.n28 10.6151
R1035 B.n735 B.n734 10.6151
R1036 B.n734 B.n733 10.6151
R1037 B.n733 B.n30 10.6151
R1038 B.n729 B.n30 10.6151
R1039 B.n729 B.n728 10.6151
R1040 B.n728 B.n727 10.6151
R1041 B.n727 B.n32 10.6151
R1042 B.n723 B.n32 10.6151
R1043 B.n723 B.n722 10.6151
R1044 B.n722 B.n721 10.6151
R1045 B.n721 B.n34 10.6151
R1046 B.n717 B.n34 10.6151
R1047 B.n717 B.n716 10.6151
R1048 B.n716 B.n715 10.6151
R1049 B.n715 B.n36 10.6151
R1050 B.n711 B.n36 10.6151
R1051 B.n711 B.n710 10.6151
R1052 B.n710 B.n709 10.6151
R1053 B.n709 B.n38 10.6151
R1054 B.n705 B.n38 10.6151
R1055 B.n705 B.n704 10.6151
R1056 B.n704 B.n703 10.6151
R1057 B.n703 B.n40 10.6151
R1058 B.n699 B.n40 10.6151
R1059 B.n699 B.n698 10.6151
R1060 B.n698 B.n697 10.6151
R1061 B.n697 B.n42 10.6151
R1062 B.n693 B.n42 10.6151
R1063 B.n693 B.n692 10.6151
R1064 B.n692 B.n691 10.6151
R1065 B.n691 B.n44 10.6151
R1066 B.n687 B.n44 10.6151
R1067 B.n687 B.n686 10.6151
R1068 B.n686 B.n685 10.6151
R1069 B.n685 B.n46 10.6151
R1070 B.n681 B.n46 10.6151
R1071 B.n681 B.n680 10.6151
R1072 B.n680 B.n679 10.6151
R1073 B.n679 B.n48 10.6151
R1074 B.n675 B.n48 10.6151
R1075 B.n675 B.n674 10.6151
R1076 B.n672 B.n52 10.6151
R1077 B.n668 B.n52 10.6151
R1078 B.n668 B.n667 10.6151
R1079 B.n667 B.n666 10.6151
R1080 B.n666 B.n54 10.6151
R1081 B.n662 B.n54 10.6151
R1082 B.n662 B.n661 10.6151
R1083 B.n661 B.n660 10.6151
R1084 B.n660 B.n56 10.6151
R1085 B.n656 B.n655 10.6151
R1086 B.n655 B.n654 10.6151
R1087 B.n654 B.n61 10.6151
R1088 B.n650 B.n61 10.6151
R1089 B.n650 B.n649 10.6151
R1090 B.n649 B.n648 10.6151
R1091 B.n648 B.n63 10.6151
R1092 B.n644 B.n63 10.6151
R1093 B.n644 B.n643 10.6151
R1094 B.n643 B.n642 10.6151
R1095 B.n642 B.n65 10.6151
R1096 B.n638 B.n65 10.6151
R1097 B.n638 B.n637 10.6151
R1098 B.n637 B.n636 10.6151
R1099 B.n636 B.n67 10.6151
R1100 B.n632 B.n67 10.6151
R1101 B.n632 B.n631 10.6151
R1102 B.n631 B.n630 10.6151
R1103 B.n630 B.n69 10.6151
R1104 B.n626 B.n69 10.6151
R1105 B.n626 B.n625 10.6151
R1106 B.n625 B.n624 10.6151
R1107 B.n624 B.n71 10.6151
R1108 B.n620 B.n71 10.6151
R1109 B.n620 B.n619 10.6151
R1110 B.n619 B.n618 10.6151
R1111 B.n618 B.n73 10.6151
R1112 B.n614 B.n73 10.6151
R1113 B.n614 B.n613 10.6151
R1114 B.n613 B.n612 10.6151
R1115 B.n612 B.n75 10.6151
R1116 B.n608 B.n75 10.6151
R1117 B.n608 B.n607 10.6151
R1118 B.n607 B.n606 10.6151
R1119 B.n606 B.n77 10.6151
R1120 B.n602 B.n77 10.6151
R1121 B.n602 B.n601 10.6151
R1122 B.n601 B.n600 10.6151
R1123 B.n600 B.n79 10.6151
R1124 B.n596 B.n79 10.6151
R1125 B.n596 B.n595 10.6151
R1126 B.n595 B.n594 10.6151
R1127 B.n594 B.n81 10.6151
R1128 B.n590 B.n81 10.6151
R1129 B.n590 B.n589 10.6151
R1130 B.n588 B.n83 10.6151
R1131 B.n584 B.n83 10.6151
R1132 B.n584 B.n583 10.6151
R1133 B.n583 B.n582 10.6151
R1134 B.n582 B.n85 10.6151
R1135 B.n578 B.n85 10.6151
R1136 B.n578 B.n577 10.6151
R1137 B.n577 B.n576 10.6151
R1138 B.n576 B.n87 10.6151
R1139 B.n572 B.n87 10.6151
R1140 B.n572 B.n571 10.6151
R1141 B.n571 B.n570 10.6151
R1142 B.n570 B.n89 10.6151
R1143 B.n566 B.n89 10.6151
R1144 B.n566 B.n565 10.6151
R1145 B.n565 B.n564 10.6151
R1146 B.n564 B.n91 10.6151
R1147 B.n560 B.n91 10.6151
R1148 B.n560 B.n559 10.6151
R1149 B.n559 B.n558 10.6151
R1150 B.n558 B.n93 10.6151
R1151 B.n554 B.n93 10.6151
R1152 B.n554 B.n553 10.6151
R1153 B.n553 B.n552 10.6151
R1154 B.n552 B.n95 10.6151
R1155 B.n548 B.n95 10.6151
R1156 B.n548 B.n547 10.6151
R1157 B.n547 B.n546 10.6151
R1158 B.n546 B.n97 10.6151
R1159 B.n542 B.n97 10.6151
R1160 B.n542 B.n541 10.6151
R1161 B.n541 B.n540 10.6151
R1162 B.n540 B.n99 10.6151
R1163 B.n536 B.n99 10.6151
R1164 B.n536 B.n535 10.6151
R1165 B.n535 B.n534 10.6151
R1166 B.n534 B.n101 10.6151
R1167 B.n530 B.n101 10.6151
R1168 B.n530 B.n529 10.6151
R1169 B.n529 B.n528 10.6151
R1170 B.n528 B.n103 10.6151
R1171 B.n524 B.n103 10.6151
R1172 B.n524 B.n523 10.6151
R1173 B.n523 B.n522 10.6151
R1174 B.n522 B.n105 10.6151
R1175 B.n518 B.n105 10.6151
R1176 B.n518 B.n517 10.6151
R1177 B.n517 B.n516 10.6151
R1178 B.n516 B.n107 10.6151
R1179 B.n512 B.n107 10.6151
R1180 B.n512 B.n511 10.6151
R1181 B.n511 B.n510 10.6151
R1182 B.n510 B.n109 10.6151
R1183 B.n506 B.n109 10.6151
R1184 B.n506 B.n505 10.6151
R1185 B.n505 B.n504 10.6151
R1186 B.n504 B.n111 10.6151
R1187 B.n500 B.n111 10.6151
R1188 B.n500 B.n499 10.6151
R1189 B.n499 B.n498 10.6151
R1190 B.n498 B.n113 10.6151
R1191 B.n494 B.n113 10.6151
R1192 B.n494 B.n493 10.6151
R1193 B.n493 B.n492 10.6151
R1194 B.n492 B.n115 10.6151
R1195 B.n488 B.n115 10.6151
R1196 B.n488 B.n487 10.6151
R1197 B.n487 B.n486 10.6151
R1198 B.n486 B.n117 10.6151
R1199 B.n482 B.n117 10.6151
R1200 B.n482 B.n481 10.6151
R1201 B.n481 B.n480 10.6151
R1202 B.n480 B.n119 10.6151
R1203 B.n476 B.n119 10.6151
R1204 B.n476 B.n475 10.6151
R1205 B.n475 B.n474 10.6151
R1206 B.n474 B.n121 10.6151
R1207 B.n470 B.n121 10.6151
R1208 B.n470 B.n469 10.6151
R1209 B.n469 B.n468 10.6151
R1210 B.n468 B.n123 10.6151
R1211 B.n464 B.n123 10.6151
R1212 B.n464 B.n463 10.6151
R1213 B.n463 B.n462 10.6151
R1214 B.n462 B.n125 10.6151
R1215 B.n458 B.n125 10.6151
R1216 B.n458 B.n457 10.6151
R1217 B.n457 B.n456 10.6151
R1218 B.n456 B.n127 10.6151
R1219 B.n452 B.n127 10.6151
R1220 B.n452 B.n451 10.6151
R1221 B.n451 B.n450 10.6151
R1222 B.n450 B.n129 10.6151
R1223 B.n446 B.n129 10.6151
R1224 B.n446 B.n445 10.6151
R1225 B.n445 B.n444 10.6151
R1226 B.n444 B.n131 10.6151
R1227 B.n440 B.n131 10.6151
R1228 B.n440 B.n439 10.6151
R1229 B.n209 B.n1 10.6151
R1230 B.n212 B.n209 10.6151
R1231 B.n213 B.n212 10.6151
R1232 B.n214 B.n213 10.6151
R1233 B.n214 B.n207 10.6151
R1234 B.n218 B.n207 10.6151
R1235 B.n219 B.n218 10.6151
R1236 B.n220 B.n219 10.6151
R1237 B.n220 B.n205 10.6151
R1238 B.n224 B.n205 10.6151
R1239 B.n225 B.n224 10.6151
R1240 B.n226 B.n225 10.6151
R1241 B.n226 B.n203 10.6151
R1242 B.n230 B.n203 10.6151
R1243 B.n231 B.n230 10.6151
R1244 B.n232 B.n231 10.6151
R1245 B.n232 B.n201 10.6151
R1246 B.n236 B.n201 10.6151
R1247 B.n237 B.n236 10.6151
R1248 B.n238 B.n237 10.6151
R1249 B.n238 B.n199 10.6151
R1250 B.n242 B.n199 10.6151
R1251 B.n243 B.n242 10.6151
R1252 B.n244 B.n243 10.6151
R1253 B.n244 B.n197 10.6151
R1254 B.n248 B.n197 10.6151
R1255 B.n249 B.n248 10.6151
R1256 B.n250 B.n249 10.6151
R1257 B.n250 B.n195 10.6151
R1258 B.n254 B.n195 10.6151
R1259 B.n255 B.n254 10.6151
R1260 B.n256 B.n255 10.6151
R1261 B.n256 B.n193 10.6151
R1262 B.n260 B.n193 10.6151
R1263 B.n261 B.n260 10.6151
R1264 B.n262 B.n261 10.6151
R1265 B.n262 B.n191 10.6151
R1266 B.n266 B.n191 10.6151
R1267 B.n267 B.n266 10.6151
R1268 B.n268 B.n267 10.6151
R1269 B.n268 B.n189 10.6151
R1270 B.n272 B.n189 10.6151
R1271 B.n273 B.n272 10.6151
R1272 B.n274 B.n273 10.6151
R1273 B.n274 B.n187 10.6151
R1274 B.n278 B.n187 10.6151
R1275 B.n279 B.n278 10.6151
R1276 B.n280 B.n279 10.6151
R1277 B.n284 B.n185 10.6151
R1278 B.n285 B.n284 10.6151
R1279 B.n286 B.n285 10.6151
R1280 B.n286 B.n183 10.6151
R1281 B.n290 B.n183 10.6151
R1282 B.n291 B.n290 10.6151
R1283 B.n292 B.n291 10.6151
R1284 B.n292 B.n181 10.6151
R1285 B.n296 B.n181 10.6151
R1286 B.n297 B.n296 10.6151
R1287 B.n298 B.n297 10.6151
R1288 B.n298 B.n179 10.6151
R1289 B.n302 B.n179 10.6151
R1290 B.n303 B.n302 10.6151
R1291 B.n304 B.n303 10.6151
R1292 B.n304 B.n177 10.6151
R1293 B.n308 B.n177 10.6151
R1294 B.n309 B.n308 10.6151
R1295 B.n310 B.n309 10.6151
R1296 B.n310 B.n175 10.6151
R1297 B.n314 B.n175 10.6151
R1298 B.n315 B.n314 10.6151
R1299 B.n316 B.n315 10.6151
R1300 B.n316 B.n173 10.6151
R1301 B.n320 B.n173 10.6151
R1302 B.n321 B.n320 10.6151
R1303 B.n322 B.n321 10.6151
R1304 B.n322 B.n171 10.6151
R1305 B.n326 B.n171 10.6151
R1306 B.n327 B.n326 10.6151
R1307 B.n328 B.n327 10.6151
R1308 B.n328 B.n169 10.6151
R1309 B.n332 B.n169 10.6151
R1310 B.n333 B.n332 10.6151
R1311 B.n334 B.n333 10.6151
R1312 B.n334 B.n167 10.6151
R1313 B.n338 B.n167 10.6151
R1314 B.n339 B.n338 10.6151
R1315 B.n340 B.n339 10.6151
R1316 B.n340 B.n165 10.6151
R1317 B.n344 B.n165 10.6151
R1318 B.n345 B.n344 10.6151
R1319 B.n346 B.n345 10.6151
R1320 B.n346 B.n163 10.6151
R1321 B.n350 B.n163 10.6151
R1322 B.n353 B.n352 10.6151
R1323 B.n353 B.n159 10.6151
R1324 B.n357 B.n159 10.6151
R1325 B.n358 B.n357 10.6151
R1326 B.n359 B.n358 10.6151
R1327 B.n359 B.n157 10.6151
R1328 B.n363 B.n157 10.6151
R1329 B.n364 B.n363 10.6151
R1330 B.n368 B.n364 10.6151
R1331 B.n372 B.n155 10.6151
R1332 B.n373 B.n372 10.6151
R1333 B.n374 B.n373 10.6151
R1334 B.n374 B.n153 10.6151
R1335 B.n378 B.n153 10.6151
R1336 B.n379 B.n378 10.6151
R1337 B.n380 B.n379 10.6151
R1338 B.n380 B.n151 10.6151
R1339 B.n384 B.n151 10.6151
R1340 B.n385 B.n384 10.6151
R1341 B.n386 B.n385 10.6151
R1342 B.n386 B.n149 10.6151
R1343 B.n390 B.n149 10.6151
R1344 B.n391 B.n390 10.6151
R1345 B.n392 B.n391 10.6151
R1346 B.n392 B.n147 10.6151
R1347 B.n396 B.n147 10.6151
R1348 B.n397 B.n396 10.6151
R1349 B.n398 B.n397 10.6151
R1350 B.n398 B.n145 10.6151
R1351 B.n402 B.n145 10.6151
R1352 B.n403 B.n402 10.6151
R1353 B.n404 B.n403 10.6151
R1354 B.n404 B.n143 10.6151
R1355 B.n408 B.n143 10.6151
R1356 B.n409 B.n408 10.6151
R1357 B.n410 B.n409 10.6151
R1358 B.n410 B.n141 10.6151
R1359 B.n414 B.n141 10.6151
R1360 B.n415 B.n414 10.6151
R1361 B.n416 B.n415 10.6151
R1362 B.n416 B.n139 10.6151
R1363 B.n420 B.n139 10.6151
R1364 B.n421 B.n420 10.6151
R1365 B.n422 B.n421 10.6151
R1366 B.n422 B.n137 10.6151
R1367 B.n426 B.n137 10.6151
R1368 B.n427 B.n426 10.6151
R1369 B.n428 B.n427 10.6151
R1370 B.n428 B.n135 10.6151
R1371 B.n432 B.n135 10.6151
R1372 B.n433 B.n432 10.6151
R1373 B.n434 B.n433 10.6151
R1374 B.n434 B.n133 10.6151
R1375 B.n438 B.n133 10.6151
R1376 B.n674 B.n673 9.36635
R1377 B.n656 B.n60 9.36635
R1378 B.n351 B.n350 9.36635
R1379 B.n367 B.n155 9.36635
R1380 B.n817 B.n0 8.11757
R1381 B.n817 B.n1 8.11757
R1382 B.n673 B.n672 1.24928
R1383 B.n60 B.n56 1.24928
R1384 B.n352 B.n351 1.24928
R1385 B.n368 B.n367 1.24928
R1386 VN.n6 VN.t2 166.523
R1387 VN.n33 VN.t1 166.523
R1388 VN.n51 VN.n27 161.3
R1389 VN.n50 VN.n49 161.3
R1390 VN.n48 VN.n28 161.3
R1391 VN.n47 VN.n46 161.3
R1392 VN.n45 VN.n29 161.3
R1393 VN.n44 VN.n43 161.3
R1394 VN.n42 VN.n41 161.3
R1395 VN.n40 VN.n31 161.3
R1396 VN.n39 VN.n38 161.3
R1397 VN.n37 VN.n32 161.3
R1398 VN.n36 VN.n35 161.3
R1399 VN.n24 VN.n0 161.3
R1400 VN.n23 VN.n22 161.3
R1401 VN.n21 VN.n1 161.3
R1402 VN.n20 VN.n19 161.3
R1403 VN.n18 VN.n2 161.3
R1404 VN.n17 VN.n16 161.3
R1405 VN.n15 VN.n14 161.3
R1406 VN.n13 VN.n4 161.3
R1407 VN.n12 VN.n11 161.3
R1408 VN.n10 VN.n5 161.3
R1409 VN.n9 VN.n8 161.3
R1410 VN.n7 VN.t3 132.892
R1411 VN.n3 VN.t7 132.892
R1412 VN.n25 VN.t0 132.892
R1413 VN.n34 VN.t4 132.892
R1414 VN.n30 VN.t5 132.892
R1415 VN.n52 VN.t6 132.892
R1416 VN.n26 VN.n25 101.072
R1417 VN.n53 VN.n52 101.072
R1418 VN.n19 VN.n1 56.5617
R1419 VN.n46 VN.n28 56.5617
R1420 VN.n7 VN.n6 52.9956
R1421 VN.n34 VN.n33 52.9956
R1422 VN VN.n53 51.7785
R1423 VN.n12 VN.n5 40.577
R1424 VN.n13 VN.n12 40.577
R1425 VN.n39 VN.n32 40.577
R1426 VN.n40 VN.n39 40.577
R1427 VN.n8 VN.n5 24.5923
R1428 VN.n14 VN.n13 24.5923
R1429 VN.n18 VN.n17 24.5923
R1430 VN.n19 VN.n18 24.5923
R1431 VN.n23 VN.n1 24.5923
R1432 VN.n24 VN.n23 24.5923
R1433 VN.n35 VN.n32 24.5923
R1434 VN.n46 VN.n45 24.5923
R1435 VN.n45 VN.n44 24.5923
R1436 VN.n41 VN.n40 24.5923
R1437 VN.n51 VN.n50 24.5923
R1438 VN.n50 VN.n28 24.5923
R1439 VN.n8 VN.n7 19.674
R1440 VN.n14 VN.n3 19.674
R1441 VN.n35 VN.n34 19.674
R1442 VN.n41 VN.n30 19.674
R1443 VN.n25 VN.n24 9.83723
R1444 VN.n52 VN.n51 9.83723
R1445 VN.n36 VN.n33 6.84375
R1446 VN.n9 VN.n6 6.84375
R1447 VN.n17 VN.n3 4.91887
R1448 VN.n44 VN.n30 4.91887
R1449 VN.n53 VN.n27 0.278335
R1450 VN.n26 VN.n0 0.278335
R1451 VN.n49 VN.n27 0.189894
R1452 VN.n49 VN.n48 0.189894
R1453 VN.n48 VN.n47 0.189894
R1454 VN.n47 VN.n29 0.189894
R1455 VN.n43 VN.n29 0.189894
R1456 VN.n43 VN.n42 0.189894
R1457 VN.n42 VN.n31 0.189894
R1458 VN.n38 VN.n31 0.189894
R1459 VN.n38 VN.n37 0.189894
R1460 VN.n37 VN.n36 0.189894
R1461 VN.n10 VN.n9 0.189894
R1462 VN.n11 VN.n10 0.189894
R1463 VN.n11 VN.n4 0.189894
R1464 VN.n15 VN.n4 0.189894
R1465 VN.n16 VN.n15 0.189894
R1466 VN.n16 VN.n2 0.189894
R1467 VN.n20 VN.n2 0.189894
R1468 VN.n21 VN.n20 0.189894
R1469 VN.n22 VN.n21 0.189894
R1470 VN.n22 VN.n0 0.189894
R1471 VN VN.n26 0.153485
R1472 VDD2.n2 VDD2.n1 73.958
R1473 VDD2.n2 VDD2.n0 73.958
R1474 VDD2 VDD2.n5 73.9552
R1475 VDD2.n4 VDD2.n3 72.8067
R1476 VDD2.n4 VDD2.n2 46.3187
R1477 VDD2.n5 VDD2.t3 2.38706
R1478 VDD2.n5 VDD2.t6 2.38706
R1479 VDD2.n3 VDD2.t1 2.38706
R1480 VDD2.n3 VDD2.t2 2.38706
R1481 VDD2.n1 VDD2.t0 2.38706
R1482 VDD2.n1 VDD2.t7 2.38706
R1483 VDD2.n0 VDD2.t5 2.38706
R1484 VDD2.n0 VDD2.t4 2.38706
R1485 VDD2 VDD2.n4 1.26559
C0 w_n3770_n3692# VP 8.1476f
C1 VDD2 VTAIL 8.67311f
C2 VDD2 B 1.74398f
C3 VDD2 VN 9.70143f
C4 w_n3770_n3692# VDD2 2.06779f
C5 VDD2 VP 0.506271f
C6 VDD1 VTAIL 8.61957f
C7 VDD1 B 1.65205f
C8 VDD1 VN 0.151927f
C9 w_n3770_n3692# VDD1 1.95853f
C10 VTAIL B 5.45065f
C11 VN VTAIL 9.99226f
C12 VDD1 VP 10.0544f
C13 VN B 1.21769f
C14 w_n3770_n3692# VTAIL 4.56033f
C15 w_n3770_n3692# B 10.371099f
C16 w_n3770_n3692# VN 7.65856f
C17 VDD1 VDD2 1.71044f
C18 VP VTAIL 10.0064f
C19 VP B 2.0368f
C20 VP VN 7.79889f
C21 VDD2 VSUBS 1.8947f
C22 VDD1 VSUBS 2.41572f
C23 VTAIL VSUBS 1.387234f
C24 VN VSUBS 6.63048f
C25 VP VSUBS 3.510638f
C26 B VSUBS 4.998524f
C27 w_n3770_n3692# VSUBS 0.170962p
C28 VDD2.t5 VSUBS 0.292271f
C29 VDD2.t4 VSUBS 0.292271f
C30 VDD2.n0 VSUBS 2.35607f
C31 VDD2.t0 VSUBS 0.292271f
C32 VDD2.t7 VSUBS 0.292271f
C33 VDD2.n1 VSUBS 2.35607f
C34 VDD2.n2 VSUBS 4.14967f
C35 VDD2.t1 VSUBS 0.292271f
C36 VDD2.t2 VSUBS 0.292271f
C37 VDD2.n3 VSUBS 2.34314f
C38 VDD2.n4 VSUBS 3.57292f
C39 VDD2.t3 VSUBS 0.292271f
C40 VDD2.t6 VSUBS 0.292271f
C41 VDD2.n5 VSUBS 2.35602f
C42 VN.n0 VSUBS 0.038084f
C43 VN.t0 VSUBS 2.65687f
C44 VN.n1 VSUBS 0.037997f
C45 VN.n2 VSUBS 0.028888f
C46 VN.t7 VSUBS 2.65687f
C47 VN.n3 VSUBS 0.934287f
C48 VN.n4 VSUBS 0.028888f
C49 VN.n5 VSUBS 0.057112f
C50 VN.t2 VSUBS 2.88021f
C51 VN.n6 VSUBS 0.990414f
C52 VN.t3 VSUBS 2.65687f
C53 VN.n7 VSUBS 1.02338f
C54 VN.n8 VSUBS 0.048281f
C55 VN.n9 VSUBS 0.275395f
C56 VN.n10 VSUBS 0.028888f
C57 VN.n11 VSUBS 0.028888f
C58 VN.n12 VSUBS 0.023332f
C59 VN.n13 VSUBS 0.057112f
C60 VN.n14 VSUBS 0.048281f
C61 VN.n15 VSUBS 0.028888f
C62 VN.n16 VSUBS 0.028888f
C63 VN.n17 VSUBS 0.032413f
C64 VN.n18 VSUBS 0.05357f
C65 VN.n19 VSUBS 0.045989f
C66 VN.n20 VSUBS 0.028888f
C67 VN.n21 VSUBS 0.028888f
C68 VN.n22 VSUBS 0.028888f
C69 VN.n23 VSUBS 0.05357f
C70 VN.n24 VSUBS 0.037702f
C71 VN.n25 VSUBS 1.0252f
C72 VN.n26 VSUBS 0.045951f
C73 VN.n27 VSUBS 0.038084f
C74 VN.t6 VSUBS 2.65687f
C75 VN.n28 VSUBS 0.037997f
C76 VN.n29 VSUBS 0.028888f
C77 VN.t5 VSUBS 2.65687f
C78 VN.n30 VSUBS 0.934287f
C79 VN.n31 VSUBS 0.028888f
C80 VN.n32 VSUBS 0.057112f
C81 VN.t1 VSUBS 2.88021f
C82 VN.n33 VSUBS 0.990414f
C83 VN.t4 VSUBS 2.65687f
C84 VN.n34 VSUBS 1.02338f
C85 VN.n35 VSUBS 0.048281f
C86 VN.n36 VSUBS 0.275395f
C87 VN.n37 VSUBS 0.028888f
C88 VN.n38 VSUBS 0.028888f
C89 VN.n39 VSUBS 0.023332f
C90 VN.n40 VSUBS 0.057112f
C91 VN.n41 VSUBS 0.048281f
C92 VN.n42 VSUBS 0.028888f
C93 VN.n43 VSUBS 0.028888f
C94 VN.n44 VSUBS 0.032413f
C95 VN.n45 VSUBS 0.05357f
C96 VN.n46 VSUBS 0.045989f
C97 VN.n47 VSUBS 0.028888f
C98 VN.n48 VSUBS 0.028888f
C99 VN.n49 VSUBS 0.028888f
C100 VN.n50 VSUBS 0.05357f
C101 VN.n51 VSUBS 0.037702f
C102 VN.n52 VSUBS 1.0252f
C103 VN.n53 VSUBS 1.69211f
C104 B.n0 VSUBS 0.006555f
C105 B.n1 VSUBS 0.006555f
C106 B.n2 VSUBS 0.009695f
C107 B.n3 VSUBS 0.00743f
C108 B.n4 VSUBS 0.00743f
C109 B.n5 VSUBS 0.00743f
C110 B.n6 VSUBS 0.00743f
C111 B.n7 VSUBS 0.00743f
C112 B.n8 VSUBS 0.00743f
C113 B.n9 VSUBS 0.00743f
C114 B.n10 VSUBS 0.00743f
C115 B.n11 VSUBS 0.00743f
C116 B.n12 VSUBS 0.00743f
C117 B.n13 VSUBS 0.00743f
C118 B.n14 VSUBS 0.00743f
C119 B.n15 VSUBS 0.00743f
C120 B.n16 VSUBS 0.00743f
C121 B.n17 VSUBS 0.00743f
C122 B.n18 VSUBS 0.00743f
C123 B.n19 VSUBS 0.00743f
C124 B.n20 VSUBS 0.00743f
C125 B.n21 VSUBS 0.00743f
C126 B.n22 VSUBS 0.00743f
C127 B.n23 VSUBS 0.00743f
C128 B.n24 VSUBS 0.00743f
C129 B.n25 VSUBS 0.00743f
C130 B.n26 VSUBS 0.017011f
C131 B.n27 VSUBS 0.00743f
C132 B.n28 VSUBS 0.00743f
C133 B.n29 VSUBS 0.00743f
C134 B.n30 VSUBS 0.00743f
C135 B.n31 VSUBS 0.00743f
C136 B.n32 VSUBS 0.00743f
C137 B.n33 VSUBS 0.00743f
C138 B.n34 VSUBS 0.00743f
C139 B.n35 VSUBS 0.00743f
C140 B.n36 VSUBS 0.00743f
C141 B.n37 VSUBS 0.00743f
C142 B.n38 VSUBS 0.00743f
C143 B.n39 VSUBS 0.00743f
C144 B.n40 VSUBS 0.00743f
C145 B.n41 VSUBS 0.00743f
C146 B.n42 VSUBS 0.00743f
C147 B.n43 VSUBS 0.00743f
C148 B.n44 VSUBS 0.00743f
C149 B.n45 VSUBS 0.00743f
C150 B.n46 VSUBS 0.00743f
C151 B.n47 VSUBS 0.00743f
C152 B.n48 VSUBS 0.00743f
C153 B.n49 VSUBS 0.00743f
C154 B.t4 VSUBS 0.477079f
C155 B.t5 VSUBS 0.499001f
C156 B.t3 VSUBS 1.60753f
C157 B.n50 VSUBS 0.259121f
C158 B.n51 VSUBS 0.075776f
C159 B.n52 VSUBS 0.00743f
C160 B.n53 VSUBS 0.00743f
C161 B.n54 VSUBS 0.00743f
C162 B.n55 VSUBS 0.00743f
C163 B.n56 VSUBS 0.004152f
C164 B.n57 VSUBS 0.00743f
C165 B.t1 VSUBS 0.477066f
C166 B.t2 VSUBS 0.49899f
C167 B.t0 VSUBS 1.60753f
C168 B.n58 VSUBS 0.259131f
C169 B.n59 VSUBS 0.075788f
C170 B.n60 VSUBS 0.017213f
C171 B.n61 VSUBS 0.00743f
C172 B.n62 VSUBS 0.00743f
C173 B.n63 VSUBS 0.00743f
C174 B.n64 VSUBS 0.00743f
C175 B.n65 VSUBS 0.00743f
C176 B.n66 VSUBS 0.00743f
C177 B.n67 VSUBS 0.00743f
C178 B.n68 VSUBS 0.00743f
C179 B.n69 VSUBS 0.00743f
C180 B.n70 VSUBS 0.00743f
C181 B.n71 VSUBS 0.00743f
C182 B.n72 VSUBS 0.00743f
C183 B.n73 VSUBS 0.00743f
C184 B.n74 VSUBS 0.00743f
C185 B.n75 VSUBS 0.00743f
C186 B.n76 VSUBS 0.00743f
C187 B.n77 VSUBS 0.00743f
C188 B.n78 VSUBS 0.00743f
C189 B.n79 VSUBS 0.00743f
C190 B.n80 VSUBS 0.00743f
C191 B.n81 VSUBS 0.00743f
C192 B.n82 VSUBS 0.017296f
C193 B.n83 VSUBS 0.00743f
C194 B.n84 VSUBS 0.00743f
C195 B.n85 VSUBS 0.00743f
C196 B.n86 VSUBS 0.00743f
C197 B.n87 VSUBS 0.00743f
C198 B.n88 VSUBS 0.00743f
C199 B.n89 VSUBS 0.00743f
C200 B.n90 VSUBS 0.00743f
C201 B.n91 VSUBS 0.00743f
C202 B.n92 VSUBS 0.00743f
C203 B.n93 VSUBS 0.00743f
C204 B.n94 VSUBS 0.00743f
C205 B.n95 VSUBS 0.00743f
C206 B.n96 VSUBS 0.00743f
C207 B.n97 VSUBS 0.00743f
C208 B.n98 VSUBS 0.00743f
C209 B.n99 VSUBS 0.00743f
C210 B.n100 VSUBS 0.00743f
C211 B.n101 VSUBS 0.00743f
C212 B.n102 VSUBS 0.00743f
C213 B.n103 VSUBS 0.00743f
C214 B.n104 VSUBS 0.00743f
C215 B.n105 VSUBS 0.00743f
C216 B.n106 VSUBS 0.00743f
C217 B.n107 VSUBS 0.00743f
C218 B.n108 VSUBS 0.00743f
C219 B.n109 VSUBS 0.00743f
C220 B.n110 VSUBS 0.00743f
C221 B.n111 VSUBS 0.00743f
C222 B.n112 VSUBS 0.00743f
C223 B.n113 VSUBS 0.00743f
C224 B.n114 VSUBS 0.00743f
C225 B.n115 VSUBS 0.00743f
C226 B.n116 VSUBS 0.00743f
C227 B.n117 VSUBS 0.00743f
C228 B.n118 VSUBS 0.00743f
C229 B.n119 VSUBS 0.00743f
C230 B.n120 VSUBS 0.00743f
C231 B.n121 VSUBS 0.00743f
C232 B.n122 VSUBS 0.00743f
C233 B.n123 VSUBS 0.00743f
C234 B.n124 VSUBS 0.00743f
C235 B.n125 VSUBS 0.00743f
C236 B.n126 VSUBS 0.00743f
C237 B.n127 VSUBS 0.00743f
C238 B.n128 VSUBS 0.00743f
C239 B.n129 VSUBS 0.00743f
C240 B.n130 VSUBS 0.00743f
C241 B.n131 VSUBS 0.00743f
C242 B.n132 VSUBS 0.017011f
C243 B.n133 VSUBS 0.00743f
C244 B.n134 VSUBS 0.00743f
C245 B.n135 VSUBS 0.00743f
C246 B.n136 VSUBS 0.00743f
C247 B.n137 VSUBS 0.00743f
C248 B.n138 VSUBS 0.00743f
C249 B.n139 VSUBS 0.00743f
C250 B.n140 VSUBS 0.00743f
C251 B.n141 VSUBS 0.00743f
C252 B.n142 VSUBS 0.00743f
C253 B.n143 VSUBS 0.00743f
C254 B.n144 VSUBS 0.00743f
C255 B.n145 VSUBS 0.00743f
C256 B.n146 VSUBS 0.00743f
C257 B.n147 VSUBS 0.00743f
C258 B.n148 VSUBS 0.00743f
C259 B.n149 VSUBS 0.00743f
C260 B.n150 VSUBS 0.00743f
C261 B.n151 VSUBS 0.00743f
C262 B.n152 VSUBS 0.00743f
C263 B.n153 VSUBS 0.00743f
C264 B.n154 VSUBS 0.00743f
C265 B.n155 VSUBS 0.006993f
C266 B.n156 VSUBS 0.00743f
C267 B.n157 VSUBS 0.00743f
C268 B.n158 VSUBS 0.00743f
C269 B.n159 VSUBS 0.00743f
C270 B.n160 VSUBS 0.00743f
C271 B.t11 VSUBS 0.477079f
C272 B.t10 VSUBS 0.499001f
C273 B.t9 VSUBS 1.60753f
C274 B.n161 VSUBS 0.259121f
C275 B.n162 VSUBS 0.075776f
C276 B.n163 VSUBS 0.00743f
C277 B.n164 VSUBS 0.00743f
C278 B.n165 VSUBS 0.00743f
C279 B.n166 VSUBS 0.00743f
C280 B.n167 VSUBS 0.00743f
C281 B.n168 VSUBS 0.00743f
C282 B.n169 VSUBS 0.00743f
C283 B.n170 VSUBS 0.00743f
C284 B.n171 VSUBS 0.00743f
C285 B.n172 VSUBS 0.00743f
C286 B.n173 VSUBS 0.00743f
C287 B.n174 VSUBS 0.00743f
C288 B.n175 VSUBS 0.00743f
C289 B.n176 VSUBS 0.00743f
C290 B.n177 VSUBS 0.00743f
C291 B.n178 VSUBS 0.00743f
C292 B.n179 VSUBS 0.00743f
C293 B.n180 VSUBS 0.00743f
C294 B.n181 VSUBS 0.00743f
C295 B.n182 VSUBS 0.00743f
C296 B.n183 VSUBS 0.00743f
C297 B.n184 VSUBS 0.00743f
C298 B.n185 VSUBS 0.017296f
C299 B.n186 VSUBS 0.00743f
C300 B.n187 VSUBS 0.00743f
C301 B.n188 VSUBS 0.00743f
C302 B.n189 VSUBS 0.00743f
C303 B.n190 VSUBS 0.00743f
C304 B.n191 VSUBS 0.00743f
C305 B.n192 VSUBS 0.00743f
C306 B.n193 VSUBS 0.00743f
C307 B.n194 VSUBS 0.00743f
C308 B.n195 VSUBS 0.00743f
C309 B.n196 VSUBS 0.00743f
C310 B.n197 VSUBS 0.00743f
C311 B.n198 VSUBS 0.00743f
C312 B.n199 VSUBS 0.00743f
C313 B.n200 VSUBS 0.00743f
C314 B.n201 VSUBS 0.00743f
C315 B.n202 VSUBS 0.00743f
C316 B.n203 VSUBS 0.00743f
C317 B.n204 VSUBS 0.00743f
C318 B.n205 VSUBS 0.00743f
C319 B.n206 VSUBS 0.00743f
C320 B.n207 VSUBS 0.00743f
C321 B.n208 VSUBS 0.00743f
C322 B.n209 VSUBS 0.00743f
C323 B.n210 VSUBS 0.00743f
C324 B.n211 VSUBS 0.00743f
C325 B.n212 VSUBS 0.00743f
C326 B.n213 VSUBS 0.00743f
C327 B.n214 VSUBS 0.00743f
C328 B.n215 VSUBS 0.00743f
C329 B.n216 VSUBS 0.00743f
C330 B.n217 VSUBS 0.00743f
C331 B.n218 VSUBS 0.00743f
C332 B.n219 VSUBS 0.00743f
C333 B.n220 VSUBS 0.00743f
C334 B.n221 VSUBS 0.00743f
C335 B.n222 VSUBS 0.00743f
C336 B.n223 VSUBS 0.00743f
C337 B.n224 VSUBS 0.00743f
C338 B.n225 VSUBS 0.00743f
C339 B.n226 VSUBS 0.00743f
C340 B.n227 VSUBS 0.00743f
C341 B.n228 VSUBS 0.00743f
C342 B.n229 VSUBS 0.00743f
C343 B.n230 VSUBS 0.00743f
C344 B.n231 VSUBS 0.00743f
C345 B.n232 VSUBS 0.00743f
C346 B.n233 VSUBS 0.00743f
C347 B.n234 VSUBS 0.00743f
C348 B.n235 VSUBS 0.00743f
C349 B.n236 VSUBS 0.00743f
C350 B.n237 VSUBS 0.00743f
C351 B.n238 VSUBS 0.00743f
C352 B.n239 VSUBS 0.00743f
C353 B.n240 VSUBS 0.00743f
C354 B.n241 VSUBS 0.00743f
C355 B.n242 VSUBS 0.00743f
C356 B.n243 VSUBS 0.00743f
C357 B.n244 VSUBS 0.00743f
C358 B.n245 VSUBS 0.00743f
C359 B.n246 VSUBS 0.00743f
C360 B.n247 VSUBS 0.00743f
C361 B.n248 VSUBS 0.00743f
C362 B.n249 VSUBS 0.00743f
C363 B.n250 VSUBS 0.00743f
C364 B.n251 VSUBS 0.00743f
C365 B.n252 VSUBS 0.00743f
C366 B.n253 VSUBS 0.00743f
C367 B.n254 VSUBS 0.00743f
C368 B.n255 VSUBS 0.00743f
C369 B.n256 VSUBS 0.00743f
C370 B.n257 VSUBS 0.00743f
C371 B.n258 VSUBS 0.00743f
C372 B.n259 VSUBS 0.00743f
C373 B.n260 VSUBS 0.00743f
C374 B.n261 VSUBS 0.00743f
C375 B.n262 VSUBS 0.00743f
C376 B.n263 VSUBS 0.00743f
C377 B.n264 VSUBS 0.00743f
C378 B.n265 VSUBS 0.00743f
C379 B.n266 VSUBS 0.00743f
C380 B.n267 VSUBS 0.00743f
C381 B.n268 VSUBS 0.00743f
C382 B.n269 VSUBS 0.00743f
C383 B.n270 VSUBS 0.00743f
C384 B.n271 VSUBS 0.00743f
C385 B.n272 VSUBS 0.00743f
C386 B.n273 VSUBS 0.00743f
C387 B.n274 VSUBS 0.00743f
C388 B.n275 VSUBS 0.00743f
C389 B.n276 VSUBS 0.00743f
C390 B.n277 VSUBS 0.00743f
C391 B.n278 VSUBS 0.00743f
C392 B.n279 VSUBS 0.00743f
C393 B.n280 VSUBS 0.017011f
C394 B.n281 VSUBS 0.017011f
C395 B.n282 VSUBS 0.017296f
C396 B.n283 VSUBS 0.00743f
C397 B.n284 VSUBS 0.00743f
C398 B.n285 VSUBS 0.00743f
C399 B.n286 VSUBS 0.00743f
C400 B.n287 VSUBS 0.00743f
C401 B.n288 VSUBS 0.00743f
C402 B.n289 VSUBS 0.00743f
C403 B.n290 VSUBS 0.00743f
C404 B.n291 VSUBS 0.00743f
C405 B.n292 VSUBS 0.00743f
C406 B.n293 VSUBS 0.00743f
C407 B.n294 VSUBS 0.00743f
C408 B.n295 VSUBS 0.00743f
C409 B.n296 VSUBS 0.00743f
C410 B.n297 VSUBS 0.00743f
C411 B.n298 VSUBS 0.00743f
C412 B.n299 VSUBS 0.00743f
C413 B.n300 VSUBS 0.00743f
C414 B.n301 VSUBS 0.00743f
C415 B.n302 VSUBS 0.00743f
C416 B.n303 VSUBS 0.00743f
C417 B.n304 VSUBS 0.00743f
C418 B.n305 VSUBS 0.00743f
C419 B.n306 VSUBS 0.00743f
C420 B.n307 VSUBS 0.00743f
C421 B.n308 VSUBS 0.00743f
C422 B.n309 VSUBS 0.00743f
C423 B.n310 VSUBS 0.00743f
C424 B.n311 VSUBS 0.00743f
C425 B.n312 VSUBS 0.00743f
C426 B.n313 VSUBS 0.00743f
C427 B.n314 VSUBS 0.00743f
C428 B.n315 VSUBS 0.00743f
C429 B.n316 VSUBS 0.00743f
C430 B.n317 VSUBS 0.00743f
C431 B.n318 VSUBS 0.00743f
C432 B.n319 VSUBS 0.00743f
C433 B.n320 VSUBS 0.00743f
C434 B.n321 VSUBS 0.00743f
C435 B.n322 VSUBS 0.00743f
C436 B.n323 VSUBS 0.00743f
C437 B.n324 VSUBS 0.00743f
C438 B.n325 VSUBS 0.00743f
C439 B.n326 VSUBS 0.00743f
C440 B.n327 VSUBS 0.00743f
C441 B.n328 VSUBS 0.00743f
C442 B.n329 VSUBS 0.00743f
C443 B.n330 VSUBS 0.00743f
C444 B.n331 VSUBS 0.00743f
C445 B.n332 VSUBS 0.00743f
C446 B.n333 VSUBS 0.00743f
C447 B.n334 VSUBS 0.00743f
C448 B.n335 VSUBS 0.00743f
C449 B.n336 VSUBS 0.00743f
C450 B.n337 VSUBS 0.00743f
C451 B.n338 VSUBS 0.00743f
C452 B.n339 VSUBS 0.00743f
C453 B.n340 VSUBS 0.00743f
C454 B.n341 VSUBS 0.00743f
C455 B.n342 VSUBS 0.00743f
C456 B.n343 VSUBS 0.00743f
C457 B.n344 VSUBS 0.00743f
C458 B.n345 VSUBS 0.00743f
C459 B.n346 VSUBS 0.00743f
C460 B.n347 VSUBS 0.00743f
C461 B.n348 VSUBS 0.00743f
C462 B.n349 VSUBS 0.00743f
C463 B.n350 VSUBS 0.006993f
C464 B.n351 VSUBS 0.017213f
C465 B.n352 VSUBS 0.004152f
C466 B.n353 VSUBS 0.00743f
C467 B.n354 VSUBS 0.00743f
C468 B.n355 VSUBS 0.00743f
C469 B.n356 VSUBS 0.00743f
C470 B.n357 VSUBS 0.00743f
C471 B.n358 VSUBS 0.00743f
C472 B.n359 VSUBS 0.00743f
C473 B.n360 VSUBS 0.00743f
C474 B.n361 VSUBS 0.00743f
C475 B.n362 VSUBS 0.00743f
C476 B.n363 VSUBS 0.00743f
C477 B.n364 VSUBS 0.00743f
C478 B.t8 VSUBS 0.477066f
C479 B.t7 VSUBS 0.49899f
C480 B.t6 VSUBS 1.60753f
C481 B.n365 VSUBS 0.259131f
C482 B.n366 VSUBS 0.075788f
C483 B.n367 VSUBS 0.017213f
C484 B.n368 VSUBS 0.004152f
C485 B.n369 VSUBS 0.00743f
C486 B.n370 VSUBS 0.00743f
C487 B.n371 VSUBS 0.00743f
C488 B.n372 VSUBS 0.00743f
C489 B.n373 VSUBS 0.00743f
C490 B.n374 VSUBS 0.00743f
C491 B.n375 VSUBS 0.00743f
C492 B.n376 VSUBS 0.00743f
C493 B.n377 VSUBS 0.00743f
C494 B.n378 VSUBS 0.00743f
C495 B.n379 VSUBS 0.00743f
C496 B.n380 VSUBS 0.00743f
C497 B.n381 VSUBS 0.00743f
C498 B.n382 VSUBS 0.00743f
C499 B.n383 VSUBS 0.00743f
C500 B.n384 VSUBS 0.00743f
C501 B.n385 VSUBS 0.00743f
C502 B.n386 VSUBS 0.00743f
C503 B.n387 VSUBS 0.00743f
C504 B.n388 VSUBS 0.00743f
C505 B.n389 VSUBS 0.00743f
C506 B.n390 VSUBS 0.00743f
C507 B.n391 VSUBS 0.00743f
C508 B.n392 VSUBS 0.00743f
C509 B.n393 VSUBS 0.00743f
C510 B.n394 VSUBS 0.00743f
C511 B.n395 VSUBS 0.00743f
C512 B.n396 VSUBS 0.00743f
C513 B.n397 VSUBS 0.00743f
C514 B.n398 VSUBS 0.00743f
C515 B.n399 VSUBS 0.00743f
C516 B.n400 VSUBS 0.00743f
C517 B.n401 VSUBS 0.00743f
C518 B.n402 VSUBS 0.00743f
C519 B.n403 VSUBS 0.00743f
C520 B.n404 VSUBS 0.00743f
C521 B.n405 VSUBS 0.00743f
C522 B.n406 VSUBS 0.00743f
C523 B.n407 VSUBS 0.00743f
C524 B.n408 VSUBS 0.00743f
C525 B.n409 VSUBS 0.00743f
C526 B.n410 VSUBS 0.00743f
C527 B.n411 VSUBS 0.00743f
C528 B.n412 VSUBS 0.00743f
C529 B.n413 VSUBS 0.00743f
C530 B.n414 VSUBS 0.00743f
C531 B.n415 VSUBS 0.00743f
C532 B.n416 VSUBS 0.00743f
C533 B.n417 VSUBS 0.00743f
C534 B.n418 VSUBS 0.00743f
C535 B.n419 VSUBS 0.00743f
C536 B.n420 VSUBS 0.00743f
C537 B.n421 VSUBS 0.00743f
C538 B.n422 VSUBS 0.00743f
C539 B.n423 VSUBS 0.00743f
C540 B.n424 VSUBS 0.00743f
C541 B.n425 VSUBS 0.00743f
C542 B.n426 VSUBS 0.00743f
C543 B.n427 VSUBS 0.00743f
C544 B.n428 VSUBS 0.00743f
C545 B.n429 VSUBS 0.00743f
C546 B.n430 VSUBS 0.00743f
C547 B.n431 VSUBS 0.00743f
C548 B.n432 VSUBS 0.00743f
C549 B.n433 VSUBS 0.00743f
C550 B.n434 VSUBS 0.00743f
C551 B.n435 VSUBS 0.00743f
C552 B.n436 VSUBS 0.00743f
C553 B.n437 VSUBS 0.017296f
C554 B.n438 VSUBS 0.0164f
C555 B.n439 VSUBS 0.017907f
C556 B.n440 VSUBS 0.00743f
C557 B.n441 VSUBS 0.00743f
C558 B.n442 VSUBS 0.00743f
C559 B.n443 VSUBS 0.00743f
C560 B.n444 VSUBS 0.00743f
C561 B.n445 VSUBS 0.00743f
C562 B.n446 VSUBS 0.00743f
C563 B.n447 VSUBS 0.00743f
C564 B.n448 VSUBS 0.00743f
C565 B.n449 VSUBS 0.00743f
C566 B.n450 VSUBS 0.00743f
C567 B.n451 VSUBS 0.00743f
C568 B.n452 VSUBS 0.00743f
C569 B.n453 VSUBS 0.00743f
C570 B.n454 VSUBS 0.00743f
C571 B.n455 VSUBS 0.00743f
C572 B.n456 VSUBS 0.00743f
C573 B.n457 VSUBS 0.00743f
C574 B.n458 VSUBS 0.00743f
C575 B.n459 VSUBS 0.00743f
C576 B.n460 VSUBS 0.00743f
C577 B.n461 VSUBS 0.00743f
C578 B.n462 VSUBS 0.00743f
C579 B.n463 VSUBS 0.00743f
C580 B.n464 VSUBS 0.00743f
C581 B.n465 VSUBS 0.00743f
C582 B.n466 VSUBS 0.00743f
C583 B.n467 VSUBS 0.00743f
C584 B.n468 VSUBS 0.00743f
C585 B.n469 VSUBS 0.00743f
C586 B.n470 VSUBS 0.00743f
C587 B.n471 VSUBS 0.00743f
C588 B.n472 VSUBS 0.00743f
C589 B.n473 VSUBS 0.00743f
C590 B.n474 VSUBS 0.00743f
C591 B.n475 VSUBS 0.00743f
C592 B.n476 VSUBS 0.00743f
C593 B.n477 VSUBS 0.00743f
C594 B.n478 VSUBS 0.00743f
C595 B.n479 VSUBS 0.00743f
C596 B.n480 VSUBS 0.00743f
C597 B.n481 VSUBS 0.00743f
C598 B.n482 VSUBS 0.00743f
C599 B.n483 VSUBS 0.00743f
C600 B.n484 VSUBS 0.00743f
C601 B.n485 VSUBS 0.00743f
C602 B.n486 VSUBS 0.00743f
C603 B.n487 VSUBS 0.00743f
C604 B.n488 VSUBS 0.00743f
C605 B.n489 VSUBS 0.00743f
C606 B.n490 VSUBS 0.00743f
C607 B.n491 VSUBS 0.00743f
C608 B.n492 VSUBS 0.00743f
C609 B.n493 VSUBS 0.00743f
C610 B.n494 VSUBS 0.00743f
C611 B.n495 VSUBS 0.00743f
C612 B.n496 VSUBS 0.00743f
C613 B.n497 VSUBS 0.00743f
C614 B.n498 VSUBS 0.00743f
C615 B.n499 VSUBS 0.00743f
C616 B.n500 VSUBS 0.00743f
C617 B.n501 VSUBS 0.00743f
C618 B.n502 VSUBS 0.00743f
C619 B.n503 VSUBS 0.00743f
C620 B.n504 VSUBS 0.00743f
C621 B.n505 VSUBS 0.00743f
C622 B.n506 VSUBS 0.00743f
C623 B.n507 VSUBS 0.00743f
C624 B.n508 VSUBS 0.00743f
C625 B.n509 VSUBS 0.00743f
C626 B.n510 VSUBS 0.00743f
C627 B.n511 VSUBS 0.00743f
C628 B.n512 VSUBS 0.00743f
C629 B.n513 VSUBS 0.00743f
C630 B.n514 VSUBS 0.00743f
C631 B.n515 VSUBS 0.00743f
C632 B.n516 VSUBS 0.00743f
C633 B.n517 VSUBS 0.00743f
C634 B.n518 VSUBS 0.00743f
C635 B.n519 VSUBS 0.00743f
C636 B.n520 VSUBS 0.00743f
C637 B.n521 VSUBS 0.00743f
C638 B.n522 VSUBS 0.00743f
C639 B.n523 VSUBS 0.00743f
C640 B.n524 VSUBS 0.00743f
C641 B.n525 VSUBS 0.00743f
C642 B.n526 VSUBS 0.00743f
C643 B.n527 VSUBS 0.00743f
C644 B.n528 VSUBS 0.00743f
C645 B.n529 VSUBS 0.00743f
C646 B.n530 VSUBS 0.00743f
C647 B.n531 VSUBS 0.00743f
C648 B.n532 VSUBS 0.00743f
C649 B.n533 VSUBS 0.00743f
C650 B.n534 VSUBS 0.00743f
C651 B.n535 VSUBS 0.00743f
C652 B.n536 VSUBS 0.00743f
C653 B.n537 VSUBS 0.00743f
C654 B.n538 VSUBS 0.00743f
C655 B.n539 VSUBS 0.00743f
C656 B.n540 VSUBS 0.00743f
C657 B.n541 VSUBS 0.00743f
C658 B.n542 VSUBS 0.00743f
C659 B.n543 VSUBS 0.00743f
C660 B.n544 VSUBS 0.00743f
C661 B.n545 VSUBS 0.00743f
C662 B.n546 VSUBS 0.00743f
C663 B.n547 VSUBS 0.00743f
C664 B.n548 VSUBS 0.00743f
C665 B.n549 VSUBS 0.00743f
C666 B.n550 VSUBS 0.00743f
C667 B.n551 VSUBS 0.00743f
C668 B.n552 VSUBS 0.00743f
C669 B.n553 VSUBS 0.00743f
C670 B.n554 VSUBS 0.00743f
C671 B.n555 VSUBS 0.00743f
C672 B.n556 VSUBS 0.00743f
C673 B.n557 VSUBS 0.00743f
C674 B.n558 VSUBS 0.00743f
C675 B.n559 VSUBS 0.00743f
C676 B.n560 VSUBS 0.00743f
C677 B.n561 VSUBS 0.00743f
C678 B.n562 VSUBS 0.00743f
C679 B.n563 VSUBS 0.00743f
C680 B.n564 VSUBS 0.00743f
C681 B.n565 VSUBS 0.00743f
C682 B.n566 VSUBS 0.00743f
C683 B.n567 VSUBS 0.00743f
C684 B.n568 VSUBS 0.00743f
C685 B.n569 VSUBS 0.00743f
C686 B.n570 VSUBS 0.00743f
C687 B.n571 VSUBS 0.00743f
C688 B.n572 VSUBS 0.00743f
C689 B.n573 VSUBS 0.00743f
C690 B.n574 VSUBS 0.00743f
C691 B.n575 VSUBS 0.00743f
C692 B.n576 VSUBS 0.00743f
C693 B.n577 VSUBS 0.00743f
C694 B.n578 VSUBS 0.00743f
C695 B.n579 VSUBS 0.00743f
C696 B.n580 VSUBS 0.00743f
C697 B.n581 VSUBS 0.00743f
C698 B.n582 VSUBS 0.00743f
C699 B.n583 VSUBS 0.00743f
C700 B.n584 VSUBS 0.00743f
C701 B.n585 VSUBS 0.00743f
C702 B.n586 VSUBS 0.00743f
C703 B.n587 VSUBS 0.017011f
C704 B.n588 VSUBS 0.017011f
C705 B.n589 VSUBS 0.017296f
C706 B.n590 VSUBS 0.00743f
C707 B.n591 VSUBS 0.00743f
C708 B.n592 VSUBS 0.00743f
C709 B.n593 VSUBS 0.00743f
C710 B.n594 VSUBS 0.00743f
C711 B.n595 VSUBS 0.00743f
C712 B.n596 VSUBS 0.00743f
C713 B.n597 VSUBS 0.00743f
C714 B.n598 VSUBS 0.00743f
C715 B.n599 VSUBS 0.00743f
C716 B.n600 VSUBS 0.00743f
C717 B.n601 VSUBS 0.00743f
C718 B.n602 VSUBS 0.00743f
C719 B.n603 VSUBS 0.00743f
C720 B.n604 VSUBS 0.00743f
C721 B.n605 VSUBS 0.00743f
C722 B.n606 VSUBS 0.00743f
C723 B.n607 VSUBS 0.00743f
C724 B.n608 VSUBS 0.00743f
C725 B.n609 VSUBS 0.00743f
C726 B.n610 VSUBS 0.00743f
C727 B.n611 VSUBS 0.00743f
C728 B.n612 VSUBS 0.00743f
C729 B.n613 VSUBS 0.00743f
C730 B.n614 VSUBS 0.00743f
C731 B.n615 VSUBS 0.00743f
C732 B.n616 VSUBS 0.00743f
C733 B.n617 VSUBS 0.00743f
C734 B.n618 VSUBS 0.00743f
C735 B.n619 VSUBS 0.00743f
C736 B.n620 VSUBS 0.00743f
C737 B.n621 VSUBS 0.00743f
C738 B.n622 VSUBS 0.00743f
C739 B.n623 VSUBS 0.00743f
C740 B.n624 VSUBS 0.00743f
C741 B.n625 VSUBS 0.00743f
C742 B.n626 VSUBS 0.00743f
C743 B.n627 VSUBS 0.00743f
C744 B.n628 VSUBS 0.00743f
C745 B.n629 VSUBS 0.00743f
C746 B.n630 VSUBS 0.00743f
C747 B.n631 VSUBS 0.00743f
C748 B.n632 VSUBS 0.00743f
C749 B.n633 VSUBS 0.00743f
C750 B.n634 VSUBS 0.00743f
C751 B.n635 VSUBS 0.00743f
C752 B.n636 VSUBS 0.00743f
C753 B.n637 VSUBS 0.00743f
C754 B.n638 VSUBS 0.00743f
C755 B.n639 VSUBS 0.00743f
C756 B.n640 VSUBS 0.00743f
C757 B.n641 VSUBS 0.00743f
C758 B.n642 VSUBS 0.00743f
C759 B.n643 VSUBS 0.00743f
C760 B.n644 VSUBS 0.00743f
C761 B.n645 VSUBS 0.00743f
C762 B.n646 VSUBS 0.00743f
C763 B.n647 VSUBS 0.00743f
C764 B.n648 VSUBS 0.00743f
C765 B.n649 VSUBS 0.00743f
C766 B.n650 VSUBS 0.00743f
C767 B.n651 VSUBS 0.00743f
C768 B.n652 VSUBS 0.00743f
C769 B.n653 VSUBS 0.00743f
C770 B.n654 VSUBS 0.00743f
C771 B.n655 VSUBS 0.00743f
C772 B.n656 VSUBS 0.006993f
C773 B.n657 VSUBS 0.00743f
C774 B.n658 VSUBS 0.00743f
C775 B.n659 VSUBS 0.00743f
C776 B.n660 VSUBS 0.00743f
C777 B.n661 VSUBS 0.00743f
C778 B.n662 VSUBS 0.00743f
C779 B.n663 VSUBS 0.00743f
C780 B.n664 VSUBS 0.00743f
C781 B.n665 VSUBS 0.00743f
C782 B.n666 VSUBS 0.00743f
C783 B.n667 VSUBS 0.00743f
C784 B.n668 VSUBS 0.00743f
C785 B.n669 VSUBS 0.00743f
C786 B.n670 VSUBS 0.00743f
C787 B.n671 VSUBS 0.00743f
C788 B.n672 VSUBS 0.004152f
C789 B.n673 VSUBS 0.017213f
C790 B.n674 VSUBS 0.006993f
C791 B.n675 VSUBS 0.00743f
C792 B.n676 VSUBS 0.00743f
C793 B.n677 VSUBS 0.00743f
C794 B.n678 VSUBS 0.00743f
C795 B.n679 VSUBS 0.00743f
C796 B.n680 VSUBS 0.00743f
C797 B.n681 VSUBS 0.00743f
C798 B.n682 VSUBS 0.00743f
C799 B.n683 VSUBS 0.00743f
C800 B.n684 VSUBS 0.00743f
C801 B.n685 VSUBS 0.00743f
C802 B.n686 VSUBS 0.00743f
C803 B.n687 VSUBS 0.00743f
C804 B.n688 VSUBS 0.00743f
C805 B.n689 VSUBS 0.00743f
C806 B.n690 VSUBS 0.00743f
C807 B.n691 VSUBS 0.00743f
C808 B.n692 VSUBS 0.00743f
C809 B.n693 VSUBS 0.00743f
C810 B.n694 VSUBS 0.00743f
C811 B.n695 VSUBS 0.00743f
C812 B.n696 VSUBS 0.00743f
C813 B.n697 VSUBS 0.00743f
C814 B.n698 VSUBS 0.00743f
C815 B.n699 VSUBS 0.00743f
C816 B.n700 VSUBS 0.00743f
C817 B.n701 VSUBS 0.00743f
C818 B.n702 VSUBS 0.00743f
C819 B.n703 VSUBS 0.00743f
C820 B.n704 VSUBS 0.00743f
C821 B.n705 VSUBS 0.00743f
C822 B.n706 VSUBS 0.00743f
C823 B.n707 VSUBS 0.00743f
C824 B.n708 VSUBS 0.00743f
C825 B.n709 VSUBS 0.00743f
C826 B.n710 VSUBS 0.00743f
C827 B.n711 VSUBS 0.00743f
C828 B.n712 VSUBS 0.00743f
C829 B.n713 VSUBS 0.00743f
C830 B.n714 VSUBS 0.00743f
C831 B.n715 VSUBS 0.00743f
C832 B.n716 VSUBS 0.00743f
C833 B.n717 VSUBS 0.00743f
C834 B.n718 VSUBS 0.00743f
C835 B.n719 VSUBS 0.00743f
C836 B.n720 VSUBS 0.00743f
C837 B.n721 VSUBS 0.00743f
C838 B.n722 VSUBS 0.00743f
C839 B.n723 VSUBS 0.00743f
C840 B.n724 VSUBS 0.00743f
C841 B.n725 VSUBS 0.00743f
C842 B.n726 VSUBS 0.00743f
C843 B.n727 VSUBS 0.00743f
C844 B.n728 VSUBS 0.00743f
C845 B.n729 VSUBS 0.00743f
C846 B.n730 VSUBS 0.00743f
C847 B.n731 VSUBS 0.00743f
C848 B.n732 VSUBS 0.00743f
C849 B.n733 VSUBS 0.00743f
C850 B.n734 VSUBS 0.00743f
C851 B.n735 VSUBS 0.00743f
C852 B.n736 VSUBS 0.00743f
C853 B.n737 VSUBS 0.00743f
C854 B.n738 VSUBS 0.00743f
C855 B.n739 VSUBS 0.00743f
C856 B.n740 VSUBS 0.00743f
C857 B.n741 VSUBS 0.017296f
C858 B.n742 VSUBS 0.017296f
C859 B.n743 VSUBS 0.017011f
C860 B.n744 VSUBS 0.00743f
C861 B.n745 VSUBS 0.00743f
C862 B.n746 VSUBS 0.00743f
C863 B.n747 VSUBS 0.00743f
C864 B.n748 VSUBS 0.00743f
C865 B.n749 VSUBS 0.00743f
C866 B.n750 VSUBS 0.00743f
C867 B.n751 VSUBS 0.00743f
C868 B.n752 VSUBS 0.00743f
C869 B.n753 VSUBS 0.00743f
C870 B.n754 VSUBS 0.00743f
C871 B.n755 VSUBS 0.00743f
C872 B.n756 VSUBS 0.00743f
C873 B.n757 VSUBS 0.00743f
C874 B.n758 VSUBS 0.00743f
C875 B.n759 VSUBS 0.00743f
C876 B.n760 VSUBS 0.00743f
C877 B.n761 VSUBS 0.00743f
C878 B.n762 VSUBS 0.00743f
C879 B.n763 VSUBS 0.00743f
C880 B.n764 VSUBS 0.00743f
C881 B.n765 VSUBS 0.00743f
C882 B.n766 VSUBS 0.00743f
C883 B.n767 VSUBS 0.00743f
C884 B.n768 VSUBS 0.00743f
C885 B.n769 VSUBS 0.00743f
C886 B.n770 VSUBS 0.00743f
C887 B.n771 VSUBS 0.00743f
C888 B.n772 VSUBS 0.00743f
C889 B.n773 VSUBS 0.00743f
C890 B.n774 VSUBS 0.00743f
C891 B.n775 VSUBS 0.00743f
C892 B.n776 VSUBS 0.00743f
C893 B.n777 VSUBS 0.00743f
C894 B.n778 VSUBS 0.00743f
C895 B.n779 VSUBS 0.00743f
C896 B.n780 VSUBS 0.00743f
C897 B.n781 VSUBS 0.00743f
C898 B.n782 VSUBS 0.00743f
C899 B.n783 VSUBS 0.00743f
C900 B.n784 VSUBS 0.00743f
C901 B.n785 VSUBS 0.00743f
C902 B.n786 VSUBS 0.00743f
C903 B.n787 VSUBS 0.00743f
C904 B.n788 VSUBS 0.00743f
C905 B.n789 VSUBS 0.00743f
C906 B.n790 VSUBS 0.00743f
C907 B.n791 VSUBS 0.00743f
C908 B.n792 VSUBS 0.00743f
C909 B.n793 VSUBS 0.00743f
C910 B.n794 VSUBS 0.00743f
C911 B.n795 VSUBS 0.00743f
C912 B.n796 VSUBS 0.00743f
C913 B.n797 VSUBS 0.00743f
C914 B.n798 VSUBS 0.00743f
C915 B.n799 VSUBS 0.00743f
C916 B.n800 VSUBS 0.00743f
C917 B.n801 VSUBS 0.00743f
C918 B.n802 VSUBS 0.00743f
C919 B.n803 VSUBS 0.00743f
C920 B.n804 VSUBS 0.00743f
C921 B.n805 VSUBS 0.00743f
C922 B.n806 VSUBS 0.00743f
C923 B.n807 VSUBS 0.00743f
C924 B.n808 VSUBS 0.00743f
C925 B.n809 VSUBS 0.00743f
C926 B.n810 VSUBS 0.00743f
C927 B.n811 VSUBS 0.00743f
C928 B.n812 VSUBS 0.00743f
C929 B.n813 VSUBS 0.00743f
C930 B.n814 VSUBS 0.00743f
C931 B.n815 VSUBS 0.009695f
C932 B.n816 VSUBS 0.010328f
C933 B.n817 VSUBS 0.020538f
C934 VTAIL.t5 VSUBS 0.264146f
C935 VTAIL.t0 VSUBS 0.264146f
C936 VTAIL.n0 VSUBS 1.98289f
C937 VTAIL.n1 VSUBS 0.755073f
C938 VTAIL.t7 VSUBS 2.60381f
C939 VTAIL.n2 VSUBS 0.887109f
C940 VTAIL.t13 VSUBS 2.60381f
C941 VTAIL.n3 VSUBS 0.887109f
C942 VTAIL.t8 VSUBS 0.264146f
C943 VTAIL.t15 VSUBS 0.264146f
C944 VTAIL.n4 VSUBS 1.98289f
C945 VTAIL.n5 VSUBS 0.941355f
C946 VTAIL.t14 VSUBS 2.60381f
C947 VTAIL.n6 VSUBS 2.30273f
C948 VTAIL.t1 VSUBS 2.60381f
C949 VTAIL.n7 VSUBS 2.30273f
C950 VTAIL.t4 VSUBS 0.264146f
C951 VTAIL.t2 VSUBS 0.264146f
C952 VTAIL.n8 VSUBS 1.9829f
C953 VTAIL.n9 VSUBS 0.941351f
C954 VTAIL.t6 VSUBS 2.60381f
C955 VTAIL.n10 VSUBS 0.887105f
C956 VTAIL.t11 VSUBS 2.60381f
C957 VTAIL.n11 VSUBS 0.887105f
C958 VTAIL.t12 VSUBS 0.264146f
C959 VTAIL.t9 VSUBS 0.264146f
C960 VTAIL.n12 VSUBS 1.9829f
C961 VTAIL.n13 VSUBS 0.941351f
C962 VTAIL.t10 VSUBS 2.60381f
C963 VTAIL.n14 VSUBS 2.30273f
C964 VTAIL.t3 VSUBS 2.60381f
C965 VTAIL.n15 VSUBS 2.29813f
C966 VDD1.t1 VSUBS 0.26531f
C967 VDD1.t4 VSUBS 0.26531f
C968 VDD1.n0 VSUBS 2.14001f
C969 VDD1.t6 VSUBS 0.26531f
C970 VDD1.t2 VSUBS 0.26531f
C971 VDD1.n1 VSUBS 2.13873f
C972 VDD1.t3 VSUBS 0.26531f
C973 VDD1.t5 VSUBS 0.26531f
C974 VDD1.n2 VSUBS 2.13873f
C975 VDD1.n3 VSUBS 3.81823f
C976 VDD1.t7 VSUBS 0.26531f
C977 VDD1.t0 VSUBS 0.26531f
C978 VDD1.n4 VSUBS 2.12699f
C979 VDD1.n5 VSUBS 3.27378f
C980 VP.n0 VSUBS 0.041161f
C981 VP.t2 VSUBS 2.87152f
C982 VP.n1 VSUBS 0.041067f
C983 VP.n2 VSUBS 0.031222f
C984 VP.t0 VSUBS 2.87152f
C985 VP.n3 VSUBS 1.00977f
C986 VP.n4 VSUBS 0.031222f
C987 VP.n5 VSUBS 0.061726f
C988 VP.n6 VSUBS 0.031222f
C989 VP.t7 VSUBS 2.87152f
C990 VP.n7 VSUBS 0.049705f
C991 VP.n8 VSUBS 0.031222f
C992 VP.t1 VSUBS 2.87152f
C993 VP.n9 VSUBS 1.10803f
C994 VP.n10 VSUBS 0.041161f
C995 VP.t5 VSUBS 2.87152f
C996 VP.n11 VSUBS 0.041067f
C997 VP.n12 VSUBS 0.031222f
C998 VP.t6 VSUBS 2.87152f
C999 VP.n13 VSUBS 1.00977f
C1000 VP.n14 VSUBS 0.031222f
C1001 VP.n15 VSUBS 0.061726f
C1002 VP.t4 VSUBS 3.11291f
C1003 VP.n16 VSUBS 1.07043f
C1004 VP.t3 VSUBS 2.87152f
C1005 VP.n17 VSUBS 1.10606f
C1006 VP.n18 VSUBS 0.052182f
C1007 VP.n19 VSUBS 0.297645f
C1008 VP.n20 VSUBS 0.031222f
C1009 VP.n21 VSUBS 0.031222f
C1010 VP.n22 VSUBS 0.025217f
C1011 VP.n23 VSUBS 0.061726f
C1012 VP.n24 VSUBS 0.052182f
C1013 VP.n25 VSUBS 0.031222f
C1014 VP.n26 VSUBS 0.031222f
C1015 VP.n27 VSUBS 0.035032f
C1016 VP.n28 VSUBS 0.057898f
C1017 VP.n29 VSUBS 0.049705f
C1018 VP.n30 VSUBS 0.031222f
C1019 VP.n31 VSUBS 0.031222f
C1020 VP.n32 VSUBS 0.031222f
C1021 VP.n33 VSUBS 0.057898f
C1022 VP.n34 VSUBS 0.040748f
C1023 VP.n35 VSUBS 1.10803f
C1024 VP.n36 VSUBS 1.81212f
C1025 VP.n37 VSUBS 1.83398f
C1026 VP.n38 VSUBS 0.041161f
C1027 VP.n39 VSUBS 0.040748f
C1028 VP.n40 VSUBS 0.057898f
C1029 VP.n41 VSUBS 0.041067f
C1030 VP.n42 VSUBS 0.031222f
C1031 VP.n43 VSUBS 0.031222f
C1032 VP.n44 VSUBS 0.031222f
C1033 VP.n45 VSUBS 0.057898f
C1034 VP.n46 VSUBS 0.035032f
C1035 VP.n47 VSUBS 1.00977f
C1036 VP.n48 VSUBS 0.052182f
C1037 VP.n49 VSUBS 0.031222f
C1038 VP.n50 VSUBS 0.031222f
C1039 VP.n51 VSUBS 0.031222f
C1040 VP.n52 VSUBS 0.025217f
C1041 VP.n53 VSUBS 0.061726f
C1042 VP.n54 VSUBS 0.052182f
C1043 VP.n55 VSUBS 0.031222f
C1044 VP.n56 VSUBS 0.031222f
C1045 VP.n57 VSUBS 0.035032f
C1046 VP.n58 VSUBS 0.057898f
C1047 VP.n59 VSUBS 0.049705f
C1048 VP.n60 VSUBS 0.031222f
C1049 VP.n61 VSUBS 0.031222f
C1050 VP.n62 VSUBS 0.031222f
C1051 VP.n63 VSUBS 0.057898f
C1052 VP.n64 VSUBS 0.040748f
C1053 VP.n65 VSUBS 1.10803f
C1054 VP.n66 VSUBS 0.049663f
.ends

