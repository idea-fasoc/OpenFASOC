* NGSPICE file created from diff_pair_sample_1128.ext - technology: sky130A

.subckt diff_pair_sample_1128 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=5.5224 ps=29.1 w=14.16 l=1.44
X1 VDD2.t1 VN.t0 VTAIL.t1 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=5.5224 ps=29.1 w=14.16 l=1.44
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=5.5224 ps=29.1 w=14.16 l=1.44
X3 VDD2.t0 VN.t1 VTAIL.t0 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=5.5224 ps=29.1 w=14.16 l=1.44
X4 B.t11 B.t9 B.t10 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=0 ps=0 w=14.16 l=1.44
X5 B.t8 B.t6 B.t7 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=0 ps=0 w=14.16 l=1.44
X6 B.t5 B.t3 B.t4 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=0 ps=0 w=14.16 l=1.44
X7 B.t2 B.t0 B.t1 w_n1678_n3800# sky130_fd_pr__pfet_01v8 ad=5.5224 pd=29.1 as=0 ps=0 w=14.16 l=1.44
R0 VP.n0 VP.t1 388.084
R1 VP.n0 VP.t0 344.866
R2 VP VP.n0 0.146778
R3 VTAIL.n306 VTAIL.n234 756.745
R4 VTAIL.n72 VTAIL.n0 756.745
R5 VTAIL.n228 VTAIL.n156 756.745
R6 VTAIL.n150 VTAIL.n78 756.745
R7 VTAIL.n258 VTAIL.n257 585
R8 VTAIL.n263 VTAIL.n262 585
R9 VTAIL.n265 VTAIL.n264 585
R10 VTAIL.n254 VTAIL.n253 585
R11 VTAIL.n271 VTAIL.n270 585
R12 VTAIL.n273 VTAIL.n272 585
R13 VTAIL.n250 VTAIL.n249 585
R14 VTAIL.n280 VTAIL.n279 585
R15 VTAIL.n281 VTAIL.n248 585
R16 VTAIL.n283 VTAIL.n282 585
R17 VTAIL.n246 VTAIL.n245 585
R18 VTAIL.n289 VTAIL.n288 585
R19 VTAIL.n291 VTAIL.n290 585
R20 VTAIL.n242 VTAIL.n241 585
R21 VTAIL.n297 VTAIL.n296 585
R22 VTAIL.n299 VTAIL.n298 585
R23 VTAIL.n238 VTAIL.n237 585
R24 VTAIL.n305 VTAIL.n304 585
R25 VTAIL.n307 VTAIL.n306 585
R26 VTAIL.n24 VTAIL.n23 585
R27 VTAIL.n29 VTAIL.n28 585
R28 VTAIL.n31 VTAIL.n30 585
R29 VTAIL.n20 VTAIL.n19 585
R30 VTAIL.n37 VTAIL.n36 585
R31 VTAIL.n39 VTAIL.n38 585
R32 VTAIL.n16 VTAIL.n15 585
R33 VTAIL.n46 VTAIL.n45 585
R34 VTAIL.n47 VTAIL.n14 585
R35 VTAIL.n49 VTAIL.n48 585
R36 VTAIL.n12 VTAIL.n11 585
R37 VTAIL.n55 VTAIL.n54 585
R38 VTAIL.n57 VTAIL.n56 585
R39 VTAIL.n8 VTAIL.n7 585
R40 VTAIL.n63 VTAIL.n62 585
R41 VTAIL.n65 VTAIL.n64 585
R42 VTAIL.n4 VTAIL.n3 585
R43 VTAIL.n71 VTAIL.n70 585
R44 VTAIL.n73 VTAIL.n72 585
R45 VTAIL.n229 VTAIL.n228 585
R46 VTAIL.n227 VTAIL.n226 585
R47 VTAIL.n160 VTAIL.n159 585
R48 VTAIL.n221 VTAIL.n220 585
R49 VTAIL.n219 VTAIL.n218 585
R50 VTAIL.n164 VTAIL.n163 585
R51 VTAIL.n213 VTAIL.n212 585
R52 VTAIL.n211 VTAIL.n210 585
R53 VTAIL.n168 VTAIL.n167 585
R54 VTAIL.n205 VTAIL.n204 585
R55 VTAIL.n203 VTAIL.n170 585
R56 VTAIL.n202 VTAIL.n201 585
R57 VTAIL.n173 VTAIL.n171 585
R58 VTAIL.n196 VTAIL.n195 585
R59 VTAIL.n194 VTAIL.n193 585
R60 VTAIL.n177 VTAIL.n176 585
R61 VTAIL.n188 VTAIL.n187 585
R62 VTAIL.n186 VTAIL.n185 585
R63 VTAIL.n181 VTAIL.n180 585
R64 VTAIL.n151 VTAIL.n150 585
R65 VTAIL.n149 VTAIL.n148 585
R66 VTAIL.n82 VTAIL.n81 585
R67 VTAIL.n143 VTAIL.n142 585
R68 VTAIL.n141 VTAIL.n140 585
R69 VTAIL.n86 VTAIL.n85 585
R70 VTAIL.n135 VTAIL.n134 585
R71 VTAIL.n133 VTAIL.n132 585
R72 VTAIL.n90 VTAIL.n89 585
R73 VTAIL.n127 VTAIL.n126 585
R74 VTAIL.n125 VTAIL.n92 585
R75 VTAIL.n124 VTAIL.n123 585
R76 VTAIL.n95 VTAIL.n93 585
R77 VTAIL.n118 VTAIL.n117 585
R78 VTAIL.n116 VTAIL.n115 585
R79 VTAIL.n99 VTAIL.n98 585
R80 VTAIL.n110 VTAIL.n109 585
R81 VTAIL.n108 VTAIL.n107 585
R82 VTAIL.n103 VTAIL.n102 585
R83 VTAIL.n259 VTAIL.t1 329.036
R84 VTAIL.n25 VTAIL.t2 329.036
R85 VTAIL.n104 VTAIL.t0 329.036
R86 VTAIL.n182 VTAIL.t3 329.036
R87 VTAIL.n263 VTAIL.n257 171.744
R88 VTAIL.n264 VTAIL.n263 171.744
R89 VTAIL.n264 VTAIL.n253 171.744
R90 VTAIL.n271 VTAIL.n253 171.744
R91 VTAIL.n272 VTAIL.n271 171.744
R92 VTAIL.n272 VTAIL.n249 171.744
R93 VTAIL.n280 VTAIL.n249 171.744
R94 VTAIL.n281 VTAIL.n280 171.744
R95 VTAIL.n282 VTAIL.n281 171.744
R96 VTAIL.n282 VTAIL.n245 171.744
R97 VTAIL.n289 VTAIL.n245 171.744
R98 VTAIL.n290 VTAIL.n289 171.744
R99 VTAIL.n290 VTAIL.n241 171.744
R100 VTAIL.n297 VTAIL.n241 171.744
R101 VTAIL.n298 VTAIL.n297 171.744
R102 VTAIL.n298 VTAIL.n237 171.744
R103 VTAIL.n305 VTAIL.n237 171.744
R104 VTAIL.n306 VTAIL.n305 171.744
R105 VTAIL.n29 VTAIL.n23 171.744
R106 VTAIL.n30 VTAIL.n29 171.744
R107 VTAIL.n30 VTAIL.n19 171.744
R108 VTAIL.n37 VTAIL.n19 171.744
R109 VTAIL.n38 VTAIL.n37 171.744
R110 VTAIL.n38 VTAIL.n15 171.744
R111 VTAIL.n46 VTAIL.n15 171.744
R112 VTAIL.n47 VTAIL.n46 171.744
R113 VTAIL.n48 VTAIL.n47 171.744
R114 VTAIL.n48 VTAIL.n11 171.744
R115 VTAIL.n55 VTAIL.n11 171.744
R116 VTAIL.n56 VTAIL.n55 171.744
R117 VTAIL.n56 VTAIL.n7 171.744
R118 VTAIL.n63 VTAIL.n7 171.744
R119 VTAIL.n64 VTAIL.n63 171.744
R120 VTAIL.n64 VTAIL.n3 171.744
R121 VTAIL.n71 VTAIL.n3 171.744
R122 VTAIL.n72 VTAIL.n71 171.744
R123 VTAIL.n228 VTAIL.n227 171.744
R124 VTAIL.n227 VTAIL.n159 171.744
R125 VTAIL.n220 VTAIL.n159 171.744
R126 VTAIL.n220 VTAIL.n219 171.744
R127 VTAIL.n219 VTAIL.n163 171.744
R128 VTAIL.n212 VTAIL.n163 171.744
R129 VTAIL.n212 VTAIL.n211 171.744
R130 VTAIL.n211 VTAIL.n167 171.744
R131 VTAIL.n204 VTAIL.n167 171.744
R132 VTAIL.n204 VTAIL.n203 171.744
R133 VTAIL.n203 VTAIL.n202 171.744
R134 VTAIL.n202 VTAIL.n171 171.744
R135 VTAIL.n195 VTAIL.n171 171.744
R136 VTAIL.n195 VTAIL.n194 171.744
R137 VTAIL.n194 VTAIL.n176 171.744
R138 VTAIL.n187 VTAIL.n176 171.744
R139 VTAIL.n187 VTAIL.n186 171.744
R140 VTAIL.n186 VTAIL.n180 171.744
R141 VTAIL.n150 VTAIL.n149 171.744
R142 VTAIL.n149 VTAIL.n81 171.744
R143 VTAIL.n142 VTAIL.n81 171.744
R144 VTAIL.n142 VTAIL.n141 171.744
R145 VTAIL.n141 VTAIL.n85 171.744
R146 VTAIL.n134 VTAIL.n85 171.744
R147 VTAIL.n134 VTAIL.n133 171.744
R148 VTAIL.n133 VTAIL.n89 171.744
R149 VTAIL.n126 VTAIL.n89 171.744
R150 VTAIL.n126 VTAIL.n125 171.744
R151 VTAIL.n125 VTAIL.n124 171.744
R152 VTAIL.n124 VTAIL.n93 171.744
R153 VTAIL.n117 VTAIL.n93 171.744
R154 VTAIL.n117 VTAIL.n116 171.744
R155 VTAIL.n116 VTAIL.n98 171.744
R156 VTAIL.n109 VTAIL.n98 171.744
R157 VTAIL.n109 VTAIL.n108 171.744
R158 VTAIL.n108 VTAIL.n102 171.744
R159 VTAIL.t1 VTAIL.n257 85.8723
R160 VTAIL.t2 VTAIL.n23 85.8723
R161 VTAIL.t3 VTAIL.n180 85.8723
R162 VTAIL.t0 VTAIL.n102 85.8723
R163 VTAIL.n311 VTAIL.n310 29.8581
R164 VTAIL.n77 VTAIL.n76 29.8581
R165 VTAIL.n233 VTAIL.n232 29.8581
R166 VTAIL.n155 VTAIL.n154 29.8581
R167 VTAIL.n155 VTAIL.n77 27.6255
R168 VTAIL.n311 VTAIL.n233 26.0996
R169 VTAIL.n283 VTAIL.n248 13.1884
R170 VTAIL.n49 VTAIL.n14 13.1884
R171 VTAIL.n205 VTAIL.n170 13.1884
R172 VTAIL.n127 VTAIL.n92 13.1884
R173 VTAIL.n279 VTAIL.n278 12.8005
R174 VTAIL.n284 VTAIL.n246 12.8005
R175 VTAIL.n45 VTAIL.n44 12.8005
R176 VTAIL.n50 VTAIL.n12 12.8005
R177 VTAIL.n206 VTAIL.n168 12.8005
R178 VTAIL.n201 VTAIL.n172 12.8005
R179 VTAIL.n128 VTAIL.n90 12.8005
R180 VTAIL.n123 VTAIL.n94 12.8005
R181 VTAIL.n277 VTAIL.n250 12.0247
R182 VTAIL.n288 VTAIL.n287 12.0247
R183 VTAIL.n43 VTAIL.n16 12.0247
R184 VTAIL.n54 VTAIL.n53 12.0247
R185 VTAIL.n210 VTAIL.n209 12.0247
R186 VTAIL.n200 VTAIL.n173 12.0247
R187 VTAIL.n132 VTAIL.n131 12.0247
R188 VTAIL.n122 VTAIL.n95 12.0247
R189 VTAIL.n274 VTAIL.n273 11.249
R190 VTAIL.n291 VTAIL.n244 11.249
R191 VTAIL.n40 VTAIL.n39 11.249
R192 VTAIL.n57 VTAIL.n10 11.249
R193 VTAIL.n213 VTAIL.n166 11.249
R194 VTAIL.n197 VTAIL.n196 11.249
R195 VTAIL.n135 VTAIL.n88 11.249
R196 VTAIL.n119 VTAIL.n118 11.249
R197 VTAIL.n259 VTAIL.n258 10.7239
R198 VTAIL.n25 VTAIL.n24 10.7239
R199 VTAIL.n182 VTAIL.n181 10.7239
R200 VTAIL.n104 VTAIL.n103 10.7239
R201 VTAIL.n270 VTAIL.n252 10.4732
R202 VTAIL.n292 VTAIL.n242 10.4732
R203 VTAIL.n36 VTAIL.n18 10.4732
R204 VTAIL.n58 VTAIL.n8 10.4732
R205 VTAIL.n214 VTAIL.n164 10.4732
R206 VTAIL.n193 VTAIL.n175 10.4732
R207 VTAIL.n136 VTAIL.n86 10.4732
R208 VTAIL.n115 VTAIL.n97 10.4732
R209 VTAIL.n269 VTAIL.n254 9.69747
R210 VTAIL.n296 VTAIL.n295 9.69747
R211 VTAIL.n35 VTAIL.n20 9.69747
R212 VTAIL.n62 VTAIL.n61 9.69747
R213 VTAIL.n218 VTAIL.n217 9.69747
R214 VTAIL.n192 VTAIL.n177 9.69747
R215 VTAIL.n140 VTAIL.n139 9.69747
R216 VTAIL.n114 VTAIL.n99 9.69747
R217 VTAIL.n310 VTAIL.n309 9.45567
R218 VTAIL.n76 VTAIL.n75 9.45567
R219 VTAIL.n232 VTAIL.n231 9.45567
R220 VTAIL.n154 VTAIL.n153 9.45567
R221 VTAIL.n236 VTAIL.n235 9.3005
R222 VTAIL.n309 VTAIL.n308 9.3005
R223 VTAIL.n301 VTAIL.n300 9.3005
R224 VTAIL.n240 VTAIL.n239 9.3005
R225 VTAIL.n295 VTAIL.n294 9.3005
R226 VTAIL.n293 VTAIL.n292 9.3005
R227 VTAIL.n244 VTAIL.n243 9.3005
R228 VTAIL.n287 VTAIL.n286 9.3005
R229 VTAIL.n285 VTAIL.n284 9.3005
R230 VTAIL.n261 VTAIL.n260 9.3005
R231 VTAIL.n256 VTAIL.n255 9.3005
R232 VTAIL.n267 VTAIL.n266 9.3005
R233 VTAIL.n269 VTAIL.n268 9.3005
R234 VTAIL.n252 VTAIL.n251 9.3005
R235 VTAIL.n275 VTAIL.n274 9.3005
R236 VTAIL.n277 VTAIL.n276 9.3005
R237 VTAIL.n278 VTAIL.n247 9.3005
R238 VTAIL.n303 VTAIL.n302 9.3005
R239 VTAIL.n2 VTAIL.n1 9.3005
R240 VTAIL.n75 VTAIL.n74 9.3005
R241 VTAIL.n67 VTAIL.n66 9.3005
R242 VTAIL.n6 VTAIL.n5 9.3005
R243 VTAIL.n61 VTAIL.n60 9.3005
R244 VTAIL.n59 VTAIL.n58 9.3005
R245 VTAIL.n10 VTAIL.n9 9.3005
R246 VTAIL.n53 VTAIL.n52 9.3005
R247 VTAIL.n51 VTAIL.n50 9.3005
R248 VTAIL.n27 VTAIL.n26 9.3005
R249 VTAIL.n22 VTAIL.n21 9.3005
R250 VTAIL.n33 VTAIL.n32 9.3005
R251 VTAIL.n35 VTAIL.n34 9.3005
R252 VTAIL.n18 VTAIL.n17 9.3005
R253 VTAIL.n41 VTAIL.n40 9.3005
R254 VTAIL.n43 VTAIL.n42 9.3005
R255 VTAIL.n44 VTAIL.n13 9.3005
R256 VTAIL.n69 VTAIL.n68 9.3005
R257 VTAIL.n158 VTAIL.n157 9.3005
R258 VTAIL.n225 VTAIL.n224 9.3005
R259 VTAIL.n223 VTAIL.n222 9.3005
R260 VTAIL.n162 VTAIL.n161 9.3005
R261 VTAIL.n217 VTAIL.n216 9.3005
R262 VTAIL.n215 VTAIL.n214 9.3005
R263 VTAIL.n166 VTAIL.n165 9.3005
R264 VTAIL.n209 VTAIL.n208 9.3005
R265 VTAIL.n207 VTAIL.n206 9.3005
R266 VTAIL.n172 VTAIL.n169 9.3005
R267 VTAIL.n200 VTAIL.n199 9.3005
R268 VTAIL.n198 VTAIL.n197 9.3005
R269 VTAIL.n175 VTAIL.n174 9.3005
R270 VTAIL.n192 VTAIL.n191 9.3005
R271 VTAIL.n190 VTAIL.n189 9.3005
R272 VTAIL.n179 VTAIL.n178 9.3005
R273 VTAIL.n184 VTAIL.n183 9.3005
R274 VTAIL.n231 VTAIL.n230 9.3005
R275 VTAIL.n106 VTAIL.n105 9.3005
R276 VTAIL.n101 VTAIL.n100 9.3005
R277 VTAIL.n112 VTAIL.n111 9.3005
R278 VTAIL.n114 VTAIL.n113 9.3005
R279 VTAIL.n97 VTAIL.n96 9.3005
R280 VTAIL.n120 VTAIL.n119 9.3005
R281 VTAIL.n122 VTAIL.n121 9.3005
R282 VTAIL.n94 VTAIL.n91 9.3005
R283 VTAIL.n153 VTAIL.n152 9.3005
R284 VTAIL.n80 VTAIL.n79 9.3005
R285 VTAIL.n147 VTAIL.n146 9.3005
R286 VTAIL.n145 VTAIL.n144 9.3005
R287 VTAIL.n84 VTAIL.n83 9.3005
R288 VTAIL.n139 VTAIL.n138 9.3005
R289 VTAIL.n137 VTAIL.n136 9.3005
R290 VTAIL.n88 VTAIL.n87 9.3005
R291 VTAIL.n131 VTAIL.n130 9.3005
R292 VTAIL.n129 VTAIL.n128 9.3005
R293 VTAIL.n266 VTAIL.n265 8.92171
R294 VTAIL.n299 VTAIL.n240 8.92171
R295 VTAIL.n32 VTAIL.n31 8.92171
R296 VTAIL.n65 VTAIL.n6 8.92171
R297 VTAIL.n221 VTAIL.n162 8.92171
R298 VTAIL.n189 VTAIL.n188 8.92171
R299 VTAIL.n143 VTAIL.n84 8.92171
R300 VTAIL.n111 VTAIL.n110 8.92171
R301 VTAIL.n262 VTAIL.n256 8.14595
R302 VTAIL.n300 VTAIL.n238 8.14595
R303 VTAIL.n310 VTAIL.n234 8.14595
R304 VTAIL.n28 VTAIL.n22 8.14595
R305 VTAIL.n66 VTAIL.n4 8.14595
R306 VTAIL.n76 VTAIL.n0 8.14595
R307 VTAIL.n232 VTAIL.n156 8.14595
R308 VTAIL.n222 VTAIL.n160 8.14595
R309 VTAIL.n185 VTAIL.n179 8.14595
R310 VTAIL.n154 VTAIL.n78 8.14595
R311 VTAIL.n144 VTAIL.n82 8.14595
R312 VTAIL.n107 VTAIL.n101 8.14595
R313 VTAIL.n261 VTAIL.n258 7.3702
R314 VTAIL.n304 VTAIL.n303 7.3702
R315 VTAIL.n308 VTAIL.n307 7.3702
R316 VTAIL.n27 VTAIL.n24 7.3702
R317 VTAIL.n70 VTAIL.n69 7.3702
R318 VTAIL.n74 VTAIL.n73 7.3702
R319 VTAIL.n230 VTAIL.n229 7.3702
R320 VTAIL.n226 VTAIL.n225 7.3702
R321 VTAIL.n184 VTAIL.n181 7.3702
R322 VTAIL.n152 VTAIL.n151 7.3702
R323 VTAIL.n148 VTAIL.n147 7.3702
R324 VTAIL.n106 VTAIL.n103 7.3702
R325 VTAIL.n304 VTAIL.n236 6.59444
R326 VTAIL.n307 VTAIL.n236 6.59444
R327 VTAIL.n70 VTAIL.n2 6.59444
R328 VTAIL.n73 VTAIL.n2 6.59444
R329 VTAIL.n229 VTAIL.n158 6.59444
R330 VTAIL.n226 VTAIL.n158 6.59444
R331 VTAIL.n151 VTAIL.n80 6.59444
R332 VTAIL.n148 VTAIL.n80 6.59444
R333 VTAIL.n262 VTAIL.n261 5.81868
R334 VTAIL.n303 VTAIL.n238 5.81868
R335 VTAIL.n308 VTAIL.n234 5.81868
R336 VTAIL.n28 VTAIL.n27 5.81868
R337 VTAIL.n69 VTAIL.n4 5.81868
R338 VTAIL.n74 VTAIL.n0 5.81868
R339 VTAIL.n230 VTAIL.n156 5.81868
R340 VTAIL.n225 VTAIL.n160 5.81868
R341 VTAIL.n185 VTAIL.n184 5.81868
R342 VTAIL.n152 VTAIL.n78 5.81868
R343 VTAIL.n147 VTAIL.n82 5.81868
R344 VTAIL.n107 VTAIL.n106 5.81868
R345 VTAIL.n265 VTAIL.n256 5.04292
R346 VTAIL.n300 VTAIL.n299 5.04292
R347 VTAIL.n31 VTAIL.n22 5.04292
R348 VTAIL.n66 VTAIL.n65 5.04292
R349 VTAIL.n222 VTAIL.n221 5.04292
R350 VTAIL.n188 VTAIL.n179 5.04292
R351 VTAIL.n144 VTAIL.n143 5.04292
R352 VTAIL.n110 VTAIL.n101 5.04292
R353 VTAIL.n266 VTAIL.n254 4.26717
R354 VTAIL.n296 VTAIL.n240 4.26717
R355 VTAIL.n32 VTAIL.n20 4.26717
R356 VTAIL.n62 VTAIL.n6 4.26717
R357 VTAIL.n218 VTAIL.n162 4.26717
R358 VTAIL.n189 VTAIL.n177 4.26717
R359 VTAIL.n140 VTAIL.n84 4.26717
R360 VTAIL.n111 VTAIL.n99 4.26717
R361 VTAIL.n270 VTAIL.n269 3.49141
R362 VTAIL.n295 VTAIL.n242 3.49141
R363 VTAIL.n36 VTAIL.n35 3.49141
R364 VTAIL.n61 VTAIL.n8 3.49141
R365 VTAIL.n217 VTAIL.n164 3.49141
R366 VTAIL.n193 VTAIL.n192 3.49141
R367 VTAIL.n139 VTAIL.n86 3.49141
R368 VTAIL.n115 VTAIL.n114 3.49141
R369 VTAIL.n273 VTAIL.n252 2.71565
R370 VTAIL.n292 VTAIL.n291 2.71565
R371 VTAIL.n39 VTAIL.n18 2.71565
R372 VTAIL.n58 VTAIL.n57 2.71565
R373 VTAIL.n214 VTAIL.n213 2.71565
R374 VTAIL.n196 VTAIL.n175 2.71565
R375 VTAIL.n136 VTAIL.n135 2.71565
R376 VTAIL.n118 VTAIL.n97 2.71565
R377 VTAIL.n183 VTAIL.n182 2.41282
R378 VTAIL.n105 VTAIL.n104 2.41282
R379 VTAIL.n260 VTAIL.n259 2.41282
R380 VTAIL.n26 VTAIL.n25 2.41282
R381 VTAIL.n274 VTAIL.n250 1.93989
R382 VTAIL.n288 VTAIL.n244 1.93989
R383 VTAIL.n40 VTAIL.n16 1.93989
R384 VTAIL.n54 VTAIL.n10 1.93989
R385 VTAIL.n210 VTAIL.n166 1.93989
R386 VTAIL.n197 VTAIL.n173 1.93989
R387 VTAIL.n132 VTAIL.n88 1.93989
R388 VTAIL.n119 VTAIL.n95 1.93989
R389 VTAIL.n233 VTAIL.n155 1.23326
R390 VTAIL.n279 VTAIL.n277 1.16414
R391 VTAIL.n287 VTAIL.n246 1.16414
R392 VTAIL.n45 VTAIL.n43 1.16414
R393 VTAIL.n53 VTAIL.n12 1.16414
R394 VTAIL.n209 VTAIL.n168 1.16414
R395 VTAIL.n201 VTAIL.n200 1.16414
R396 VTAIL.n131 VTAIL.n90 1.16414
R397 VTAIL.n123 VTAIL.n122 1.16414
R398 VTAIL VTAIL.n77 0.909983
R399 VTAIL.n278 VTAIL.n248 0.388379
R400 VTAIL.n284 VTAIL.n283 0.388379
R401 VTAIL.n44 VTAIL.n14 0.388379
R402 VTAIL.n50 VTAIL.n49 0.388379
R403 VTAIL.n206 VTAIL.n205 0.388379
R404 VTAIL.n172 VTAIL.n170 0.388379
R405 VTAIL.n128 VTAIL.n127 0.388379
R406 VTAIL.n94 VTAIL.n92 0.388379
R407 VTAIL VTAIL.n311 0.323776
R408 VTAIL.n260 VTAIL.n255 0.155672
R409 VTAIL.n267 VTAIL.n255 0.155672
R410 VTAIL.n268 VTAIL.n267 0.155672
R411 VTAIL.n268 VTAIL.n251 0.155672
R412 VTAIL.n275 VTAIL.n251 0.155672
R413 VTAIL.n276 VTAIL.n275 0.155672
R414 VTAIL.n276 VTAIL.n247 0.155672
R415 VTAIL.n285 VTAIL.n247 0.155672
R416 VTAIL.n286 VTAIL.n285 0.155672
R417 VTAIL.n286 VTAIL.n243 0.155672
R418 VTAIL.n293 VTAIL.n243 0.155672
R419 VTAIL.n294 VTAIL.n293 0.155672
R420 VTAIL.n294 VTAIL.n239 0.155672
R421 VTAIL.n301 VTAIL.n239 0.155672
R422 VTAIL.n302 VTAIL.n301 0.155672
R423 VTAIL.n302 VTAIL.n235 0.155672
R424 VTAIL.n309 VTAIL.n235 0.155672
R425 VTAIL.n26 VTAIL.n21 0.155672
R426 VTAIL.n33 VTAIL.n21 0.155672
R427 VTAIL.n34 VTAIL.n33 0.155672
R428 VTAIL.n34 VTAIL.n17 0.155672
R429 VTAIL.n41 VTAIL.n17 0.155672
R430 VTAIL.n42 VTAIL.n41 0.155672
R431 VTAIL.n42 VTAIL.n13 0.155672
R432 VTAIL.n51 VTAIL.n13 0.155672
R433 VTAIL.n52 VTAIL.n51 0.155672
R434 VTAIL.n52 VTAIL.n9 0.155672
R435 VTAIL.n59 VTAIL.n9 0.155672
R436 VTAIL.n60 VTAIL.n59 0.155672
R437 VTAIL.n60 VTAIL.n5 0.155672
R438 VTAIL.n67 VTAIL.n5 0.155672
R439 VTAIL.n68 VTAIL.n67 0.155672
R440 VTAIL.n68 VTAIL.n1 0.155672
R441 VTAIL.n75 VTAIL.n1 0.155672
R442 VTAIL.n231 VTAIL.n157 0.155672
R443 VTAIL.n224 VTAIL.n157 0.155672
R444 VTAIL.n224 VTAIL.n223 0.155672
R445 VTAIL.n223 VTAIL.n161 0.155672
R446 VTAIL.n216 VTAIL.n161 0.155672
R447 VTAIL.n216 VTAIL.n215 0.155672
R448 VTAIL.n215 VTAIL.n165 0.155672
R449 VTAIL.n208 VTAIL.n165 0.155672
R450 VTAIL.n208 VTAIL.n207 0.155672
R451 VTAIL.n207 VTAIL.n169 0.155672
R452 VTAIL.n199 VTAIL.n169 0.155672
R453 VTAIL.n199 VTAIL.n198 0.155672
R454 VTAIL.n198 VTAIL.n174 0.155672
R455 VTAIL.n191 VTAIL.n174 0.155672
R456 VTAIL.n191 VTAIL.n190 0.155672
R457 VTAIL.n190 VTAIL.n178 0.155672
R458 VTAIL.n183 VTAIL.n178 0.155672
R459 VTAIL.n153 VTAIL.n79 0.155672
R460 VTAIL.n146 VTAIL.n79 0.155672
R461 VTAIL.n146 VTAIL.n145 0.155672
R462 VTAIL.n145 VTAIL.n83 0.155672
R463 VTAIL.n138 VTAIL.n83 0.155672
R464 VTAIL.n138 VTAIL.n137 0.155672
R465 VTAIL.n137 VTAIL.n87 0.155672
R466 VTAIL.n130 VTAIL.n87 0.155672
R467 VTAIL.n130 VTAIL.n129 0.155672
R468 VTAIL.n129 VTAIL.n91 0.155672
R469 VTAIL.n121 VTAIL.n91 0.155672
R470 VTAIL.n121 VTAIL.n120 0.155672
R471 VTAIL.n120 VTAIL.n96 0.155672
R472 VTAIL.n113 VTAIL.n96 0.155672
R473 VTAIL.n113 VTAIL.n112 0.155672
R474 VTAIL.n112 VTAIL.n100 0.155672
R475 VTAIL.n105 VTAIL.n100 0.155672
R476 VDD1.n72 VDD1.n0 756.745
R477 VDD1.n149 VDD1.n77 756.745
R478 VDD1.n73 VDD1.n72 585
R479 VDD1.n71 VDD1.n70 585
R480 VDD1.n4 VDD1.n3 585
R481 VDD1.n65 VDD1.n64 585
R482 VDD1.n63 VDD1.n62 585
R483 VDD1.n8 VDD1.n7 585
R484 VDD1.n57 VDD1.n56 585
R485 VDD1.n55 VDD1.n54 585
R486 VDD1.n12 VDD1.n11 585
R487 VDD1.n49 VDD1.n48 585
R488 VDD1.n47 VDD1.n14 585
R489 VDD1.n46 VDD1.n45 585
R490 VDD1.n17 VDD1.n15 585
R491 VDD1.n40 VDD1.n39 585
R492 VDD1.n38 VDD1.n37 585
R493 VDD1.n21 VDD1.n20 585
R494 VDD1.n32 VDD1.n31 585
R495 VDD1.n30 VDD1.n29 585
R496 VDD1.n25 VDD1.n24 585
R497 VDD1.n101 VDD1.n100 585
R498 VDD1.n106 VDD1.n105 585
R499 VDD1.n108 VDD1.n107 585
R500 VDD1.n97 VDD1.n96 585
R501 VDD1.n114 VDD1.n113 585
R502 VDD1.n116 VDD1.n115 585
R503 VDD1.n93 VDD1.n92 585
R504 VDD1.n123 VDD1.n122 585
R505 VDD1.n124 VDD1.n91 585
R506 VDD1.n126 VDD1.n125 585
R507 VDD1.n89 VDD1.n88 585
R508 VDD1.n132 VDD1.n131 585
R509 VDD1.n134 VDD1.n133 585
R510 VDD1.n85 VDD1.n84 585
R511 VDD1.n140 VDD1.n139 585
R512 VDD1.n142 VDD1.n141 585
R513 VDD1.n81 VDD1.n80 585
R514 VDD1.n148 VDD1.n147 585
R515 VDD1.n150 VDD1.n149 585
R516 VDD1.n102 VDD1.t1 329.036
R517 VDD1.n26 VDD1.t0 329.036
R518 VDD1.n72 VDD1.n71 171.744
R519 VDD1.n71 VDD1.n3 171.744
R520 VDD1.n64 VDD1.n3 171.744
R521 VDD1.n64 VDD1.n63 171.744
R522 VDD1.n63 VDD1.n7 171.744
R523 VDD1.n56 VDD1.n7 171.744
R524 VDD1.n56 VDD1.n55 171.744
R525 VDD1.n55 VDD1.n11 171.744
R526 VDD1.n48 VDD1.n11 171.744
R527 VDD1.n48 VDD1.n47 171.744
R528 VDD1.n47 VDD1.n46 171.744
R529 VDD1.n46 VDD1.n15 171.744
R530 VDD1.n39 VDD1.n15 171.744
R531 VDD1.n39 VDD1.n38 171.744
R532 VDD1.n38 VDD1.n20 171.744
R533 VDD1.n31 VDD1.n20 171.744
R534 VDD1.n31 VDD1.n30 171.744
R535 VDD1.n30 VDD1.n24 171.744
R536 VDD1.n106 VDD1.n100 171.744
R537 VDD1.n107 VDD1.n106 171.744
R538 VDD1.n107 VDD1.n96 171.744
R539 VDD1.n114 VDD1.n96 171.744
R540 VDD1.n115 VDD1.n114 171.744
R541 VDD1.n115 VDD1.n92 171.744
R542 VDD1.n123 VDD1.n92 171.744
R543 VDD1.n124 VDD1.n123 171.744
R544 VDD1.n125 VDD1.n124 171.744
R545 VDD1.n125 VDD1.n88 171.744
R546 VDD1.n132 VDD1.n88 171.744
R547 VDD1.n133 VDD1.n132 171.744
R548 VDD1.n133 VDD1.n84 171.744
R549 VDD1.n140 VDD1.n84 171.744
R550 VDD1.n141 VDD1.n140 171.744
R551 VDD1.n141 VDD1.n80 171.744
R552 VDD1.n148 VDD1.n80 171.744
R553 VDD1.n149 VDD1.n148 171.744
R554 VDD1 VDD1.n153 86.3612
R555 VDD1.t0 VDD1.n24 85.8723
R556 VDD1.t1 VDD1.n100 85.8723
R557 VDD1 VDD1.n76 46.9765
R558 VDD1.n49 VDD1.n14 13.1884
R559 VDD1.n126 VDD1.n91 13.1884
R560 VDD1.n50 VDD1.n12 12.8005
R561 VDD1.n45 VDD1.n16 12.8005
R562 VDD1.n122 VDD1.n121 12.8005
R563 VDD1.n127 VDD1.n89 12.8005
R564 VDD1.n54 VDD1.n53 12.0247
R565 VDD1.n44 VDD1.n17 12.0247
R566 VDD1.n120 VDD1.n93 12.0247
R567 VDD1.n131 VDD1.n130 12.0247
R568 VDD1.n57 VDD1.n10 11.249
R569 VDD1.n41 VDD1.n40 11.249
R570 VDD1.n117 VDD1.n116 11.249
R571 VDD1.n134 VDD1.n87 11.249
R572 VDD1.n26 VDD1.n25 10.7239
R573 VDD1.n102 VDD1.n101 10.7239
R574 VDD1.n58 VDD1.n8 10.4732
R575 VDD1.n37 VDD1.n19 10.4732
R576 VDD1.n113 VDD1.n95 10.4732
R577 VDD1.n135 VDD1.n85 10.4732
R578 VDD1.n62 VDD1.n61 9.69747
R579 VDD1.n36 VDD1.n21 9.69747
R580 VDD1.n112 VDD1.n97 9.69747
R581 VDD1.n139 VDD1.n138 9.69747
R582 VDD1.n76 VDD1.n75 9.45567
R583 VDD1.n153 VDD1.n152 9.45567
R584 VDD1.n2 VDD1.n1 9.3005
R585 VDD1.n69 VDD1.n68 9.3005
R586 VDD1.n67 VDD1.n66 9.3005
R587 VDD1.n6 VDD1.n5 9.3005
R588 VDD1.n61 VDD1.n60 9.3005
R589 VDD1.n59 VDD1.n58 9.3005
R590 VDD1.n10 VDD1.n9 9.3005
R591 VDD1.n53 VDD1.n52 9.3005
R592 VDD1.n51 VDD1.n50 9.3005
R593 VDD1.n16 VDD1.n13 9.3005
R594 VDD1.n44 VDD1.n43 9.3005
R595 VDD1.n42 VDD1.n41 9.3005
R596 VDD1.n19 VDD1.n18 9.3005
R597 VDD1.n36 VDD1.n35 9.3005
R598 VDD1.n34 VDD1.n33 9.3005
R599 VDD1.n23 VDD1.n22 9.3005
R600 VDD1.n28 VDD1.n27 9.3005
R601 VDD1.n75 VDD1.n74 9.3005
R602 VDD1.n79 VDD1.n78 9.3005
R603 VDD1.n152 VDD1.n151 9.3005
R604 VDD1.n144 VDD1.n143 9.3005
R605 VDD1.n83 VDD1.n82 9.3005
R606 VDD1.n138 VDD1.n137 9.3005
R607 VDD1.n136 VDD1.n135 9.3005
R608 VDD1.n87 VDD1.n86 9.3005
R609 VDD1.n130 VDD1.n129 9.3005
R610 VDD1.n128 VDD1.n127 9.3005
R611 VDD1.n104 VDD1.n103 9.3005
R612 VDD1.n99 VDD1.n98 9.3005
R613 VDD1.n110 VDD1.n109 9.3005
R614 VDD1.n112 VDD1.n111 9.3005
R615 VDD1.n95 VDD1.n94 9.3005
R616 VDD1.n118 VDD1.n117 9.3005
R617 VDD1.n120 VDD1.n119 9.3005
R618 VDD1.n121 VDD1.n90 9.3005
R619 VDD1.n146 VDD1.n145 9.3005
R620 VDD1.n65 VDD1.n6 8.92171
R621 VDD1.n33 VDD1.n32 8.92171
R622 VDD1.n109 VDD1.n108 8.92171
R623 VDD1.n142 VDD1.n83 8.92171
R624 VDD1.n76 VDD1.n0 8.14595
R625 VDD1.n66 VDD1.n4 8.14595
R626 VDD1.n29 VDD1.n23 8.14595
R627 VDD1.n105 VDD1.n99 8.14595
R628 VDD1.n143 VDD1.n81 8.14595
R629 VDD1.n153 VDD1.n77 8.14595
R630 VDD1.n74 VDD1.n73 7.3702
R631 VDD1.n70 VDD1.n69 7.3702
R632 VDD1.n28 VDD1.n25 7.3702
R633 VDD1.n104 VDD1.n101 7.3702
R634 VDD1.n147 VDD1.n146 7.3702
R635 VDD1.n151 VDD1.n150 7.3702
R636 VDD1.n73 VDD1.n2 6.59444
R637 VDD1.n70 VDD1.n2 6.59444
R638 VDD1.n147 VDD1.n79 6.59444
R639 VDD1.n150 VDD1.n79 6.59444
R640 VDD1.n74 VDD1.n0 5.81868
R641 VDD1.n69 VDD1.n4 5.81868
R642 VDD1.n29 VDD1.n28 5.81868
R643 VDD1.n105 VDD1.n104 5.81868
R644 VDD1.n146 VDD1.n81 5.81868
R645 VDD1.n151 VDD1.n77 5.81868
R646 VDD1.n66 VDD1.n65 5.04292
R647 VDD1.n32 VDD1.n23 5.04292
R648 VDD1.n108 VDD1.n99 5.04292
R649 VDD1.n143 VDD1.n142 5.04292
R650 VDD1.n62 VDD1.n6 4.26717
R651 VDD1.n33 VDD1.n21 4.26717
R652 VDD1.n109 VDD1.n97 4.26717
R653 VDD1.n139 VDD1.n83 4.26717
R654 VDD1.n61 VDD1.n8 3.49141
R655 VDD1.n37 VDD1.n36 3.49141
R656 VDD1.n113 VDD1.n112 3.49141
R657 VDD1.n138 VDD1.n85 3.49141
R658 VDD1.n58 VDD1.n57 2.71565
R659 VDD1.n40 VDD1.n19 2.71565
R660 VDD1.n116 VDD1.n95 2.71565
R661 VDD1.n135 VDD1.n134 2.71565
R662 VDD1.n27 VDD1.n26 2.41282
R663 VDD1.n103 VDD1.n102 2.41282
R664 VDD1.n54 VDD1.n10 1.93989
R665 VDD1.n41 VDD1.n17 1.93989
R666 VDD1.n117 VDD1.n93 1.93989
R667 VDD1.n131 VDD1.n87 1.93989
R668 VDD1.n53 VDD1.n12 1.16414
R669 VDD1.n45 VDD1.n44 1.16414
R670 VDD1.n122 VDD1.n120 1.16414
R671 VDD1.n130 VDD1.n89 1.16414
R672 VDD1.n50 VDD1.n49 0.388379
R673 VDD1.n16 VDD1.n14 0.388379
R674 VDD1.n121 VDD1.n91 0.388379
R675 VDD1.n127 VDD1.n126 0.388379
R676 VDD1.n75 VDD1.n1 0.155672
R677 VDD1.n68 VDD1.n1 0.155672
R678 VDD1.n68 VDD1.n67 0.155672
R679 VDD1.n67 VDD1.n5 0.155672
R680 VDD1.n60 VDD1.n5 0.155672
R681 VDD1.n60 VDD1.n59 0.155672
R682 VDD1.n59 VDD1.n9 0.155672
R683 VDD1.n52 VDD1.n9 0.155672
R684 VDD1.n52 VDD1.n51 0.155672
R685 VDD1.n51 VDD1.n13 0.155672
R686 VDD1.n43 VDD1.n13 0.155672
R687 VDD1.n43 VDD1.n42 0.155672
R688 VDD1.n42 VDD1.n18 0.155672
R689 VDD1.n35 VDD1.n18 0.155672
R690 VDD1.n35 VDD1.n34 0.155672
R691 VDD1.n34 VDD1.n22 0.155672
R692 VDD1.n27 VDD1.n22 0.155672
R693 VDD1.n103 VDD1.n98 0.155672
R694 VDD1.n110 VDD1.n98 0.155672
R695 VDD1.n111 VDD1.n110 0.155672
R696 VDD1.n111 VDD1.n94 0.155672
R697 VDD1.n118 VDD1.n94 0.155672
R698 VDD1.n119 VDD1.n118 0.155672
R699 VDD1.n119 VDD1.n90 0.155672
R700 VDD1.n128 VDD1.n90 0.155672
R701 VDD1.n129 VDD1.n128 0.155672
R702 VDD1.n129 VDD1.n86 0.155672
R703 VDD1.n136 VDD1.n86 0.155672
R704 VDD1.n137 VDD1.n136 0.155672
R705 VDD1.n137 VDD1.n82 0.155672
R706 VDD1.n144 VDD1.n82 0.155672
R707 VDD1.n145 VDD1.n144 0.155672
R708 VDD1.n145 VDD1.n78 0.155672
R709 VDD1.n152 VDD1.n78 0.155672
R710 VN VN.t1 388.37
R711 VN VN.t0 345.014
R712 VDD2.n149 VDD2.n77 756.745
R713 VDD2.n72 VDD2.n0 756.745
R714 VDD2.n150 VDD2.n149 585
R715 VDD2.n148 VDD2.n147 585
R716 VDD2.n81 VDD2.n80 585
R717 VDD2.n142 VDD2.n141 585
R718 VDD2.n140 VDD2.n139 585
R719 VDD2.n85 VDD2.n84 585
R720 VDD2.n134 VDD2.n133 585
R721 VDD2.n132 VDD2.n131 585
R722 VDD2.n89 VDD2.n88 585
R723 VDD2.n126 VDD2.n125 585
R724 VDD2.n124 VDD2.n91 585
R725 VDD2.n123 VDD2.n122 585
R726 VDD2.n94 VDD2.n92 585
R727 VDD2.n117 VDD2.n116 585
R728 VDD2.n115 VDD2.n114 585
R729 VDD2.n98 VDD2.n97 585
R730 VDD2.n109 VDD2.n108 585
R731 VDD2.n107 VDD2.n106 585
R732 VDD2.n102 VDD2.n101 585
R733 VDD2.n24 VDD2.n23 585
R734 VDD2.n29 VDD2.n28 585
R735 VDD2.n31 VDD2.n30 585
R736 VDD2.n20 VDD2.n19 585
R737 VDD2.n37 VDD2.n36 585
R738 VDD2.n39 VDD2.n38 585
R739 VDD2.n16 VDD2.n15 585
R740 VDD2.n46 VDD2.n45 585
R741 VDD2.n47 VDD2.n14 585
R742 VDD2.n49 VDD2.n48 585
R743 VDD2.n12 VDD2.n11 585
R744 VDD2.n55 VDD2.n54 585
R745 VDD2.n57 VDD2.n56 585
R746 VDD2.n8 VDD2.n7 585
R747 VDD2.n63 VDD2.n62 585
R748 VDD2.n65 VDD2.n64 585
R749 VDD2.n4 VDD2.n3 585
R750 VDD2.n71 VDD2.n70 585
R751 VDD2.n73 VDD2.n72 585
R752 VDD2.n25 VDD2.t1 329.036
R753 VDD2.n103 VDD2.t0 329.036
R754 VDD2.n149 VDD2.n148 171.744
R755 VDD2.n148 VDD2.n80 171.744
R756 VDD2.n141 VDD2.n80 171.744
R757 VDD2.n141 VDD2.n140 171.744
R758 VDD2.n140 VDD2.n84 171.744
R759 VDD2.n133 VDD2.n84 171.744
R760 VDD2.n133 VDD2.n132 171.744
R761 VDD2.n132 VDD2.n88 171.744
R762 VDD2.n125 VDD2.n88 171.744
R763 VDD2.n125 VDD2.n124 171.744
R764 VDD2.n124 VDD2.n123 171.744
R765 VDD2.n123 VDD2.n92 171.744
R766 VDD2.n116 VDD2.n92 171.744
R767 VDD2.n116 VDD2.n115 171.744
R768 VDD2.n115 VDD2.n97 171.744
R769 VDD2.n108 VDD2.n97 171.744
R770 VDD2.n108 VDD2.n107 171.744
R771 VDD2.n107 VDD2.n101 171.744
R772 VDD2.n29 VDD2.n23 171.744
R773 VDD2.n30 VDD2.n29 171.744
R774 VDD2.n30 VDD2.n19 171.744
R775 VDD2.n37 VDD2.n19 171.744
R776 VDD2.n38 VDD2.n37 171.744
R777 VDD2.n38 VDD2.n15 171.744
R778 VDD2.n46 VDD2.n15 171.744
R779 VDD2.n47 VDD2.n46 171.744
R780 VDD2.n48 VDD2.n47 171.744
R781 VDD2.n48 VDD2.n11 171.744
R782 VDD2.n55 VDD2.n11 171.744
R783 VDD2.n56 VDD2.n55 171.744
R784 VDD2.n56 VDD2.n7 171.744
R785 VDD2.n63 VDD2.n7 171.744
R786 VDD2.n64 VDD2.n63 171.744
R787 VDD2.n64 VDD2.n3 171.744
R788 VDD2.n71 VDD2.n3 171.744
R789 VDD2.n72 VDD2.n71 171.744
R790 VDD2.t0 VDD2.n101 85.8723
R791 VDD2.t1 VDD2.n23 85.8723
R792 VDD2.n154 VDD2.n76 85.4549
R793 VDD2.n154 VDD2.n153 46.5369
R794 VDD2.n126 VDD2.n91 13.1884
R795 VDD2.n49 VDD2.n14 13.1884
R796 VDD2.n127 VDD2.n89 12.8005
R797 VDD2.n122 VDD2.n93 12.8005
R798 VDD2.n45 VDD2.n44 12.8005
R799 VDD2.n50 VDD2.n12 12.8005
R800 VDD2.n131 VDD2.n130 12.0247
R801 VDD2.n121 VDD2.n94 12.0247
R802 VDD2.n43 VDD2.n16 12.0247
R803 VDD2.n54 VDD2.n53 12.0247
R804 VDD2.n134 VDD2.n87 11.249
R805 VDD2.n118 VDD2.n117 11.249
R806 VDD2.n40 VDD2.n39 11.249
R807 VDD2.n57 VDD2.n10 11.249
R808 VDD2.n103 VDD2.n102 10.7239
R809 VDD2.n25 VDD2.n24 10.7239
R810 VDD2.n135 VDD2.n85 10.4732
R811 VDD2.n114 VDD2.n96 10.4732
R812 VDD2.n36 VDD2.n18 10.4732
R813 VDD2.n58 VDD2.n8 10.4732
R814 VDD2.n139 VDD2.n138 9.69747
R815 VDD2.n113 VDD2.n98 9.69747
R816 VDD2.n35 VDD2.n20 9.69747
R817 VDD2.n62 VDD2.n61 9.69747
R818 VDD2.n153 VDD2.n152 9.45567
R819 VDD2.n76 VDD2.n75 9.45567
R820 VDD2.n79 VDD2.n78 9.3005
R821 VDD2.n146 VDD2.n145 9.3005
R822 VDD2.n144 VDD2.n143 9.3005
R823 VDD2.n83 VDD2.n82 9.3005
R824 VDD2.n138 VDD2.n137 9.3005
R825 VDD2.n136 VDD2.n135 9.3005
R826 VDD2.n87 VDD2.n86 9.3005
R827 VDD2.n130 VDD2.n129 9.3005
R828 VDD2.n128 VDD2.n127 9.3005
R829 VDD2.n93 VDD2.n90 9.3005
R830 VDD2.n121 VDD2.n120 9.3005
R831 VDD2.n119 VDD2.n118 9.3005
R832 VDD2.n96 VDD2.n95 9.3005
R833 VDD2.n113 VDD2.n112 9.3005
R834 VDD2.n111 VDD2.n110 9.3005
R835 VDD2.n100 VDD2.n99 9.3005
R836 VDD2.n105 VDD2.n104 9.3005
R837 VDD2.n152 VDD2.n151 9.3005
R838 VDD2.n2 VDD2.n1 9.3005
R839 VDD2.n75 VDD2.n74 9.3005
R840 VDD2.n67 VDD2.n66 9.3005
R841 VDD2.n6 VDD2.n5 9.3005
R842 VDD2.n61 VDD2.n60 9.3005
R843 VDD2.n59 VDD2.n58 9.3005
R844 VDD2.n10 VDD2.n9 9.3005
R845 VDD2.n53 VDD2.n52 9.3005
R846 VDD2.n51 VDD2.n50 9.3005
R847 VDD2.n27 VDD2.n26 9.3005
R848 VDD2.n22 VDD2.n21 9.3005
R849 VDD2.n33 VDD2.n32 9.3005
R850 VDD2.n35 VDD2.n34 9.3005
R851 VDD2.n18 VDD2.n17 9.3005
R852 VDD2.n41 VDD2.n40 9.3005
R853 VDD2.n43 VDD2.n42 9.3005
R854 VDD2.n44 VDD2.n13 9.3005
R855 VDD2.n69 VDD2.n68 9.3005
R856 VDD2.n142 VDD2.n83 8.92171
R857 VDD2.n110 VDD2.n109 8.92171
R858 VDD2.n32 VDD2.n31 8.92171
R859 VDD2.n65 VDD2.n6 8.92171
R860 VDD2.n153 VDD2.n77 8.14595
R861 VDD2.n143 VDD2.n81 8.14595
R862 VDD2.n106 VDD2.n100 8.14595
R863 VDD2.n28 VDD2.n22 8.14595
R864 VDD2.n66 VDD2.n4 8.14595
R865 VDD2.n76 VDD2.n0 8.14595
R866 VDD2.n151 VDD2.n150 7.3702
R867 VDD2.n147 VDD2.n146 7.3702
R868 VDD2.n105 VDD2.n102 7.3702
R869 VDD2.n27 VDD2.n24 7.3702
R870 VDD2.n70 VDD2.n69 7.3702
R871 VDD2.n74 VDD2.n73 7.3702
R872 VDD2.n150 VDD2.n79 6.59444
R873 VDD2.n147 VDD2.n79 6.59444
R874 VDD2.n70 VDD2.n2 6.59444
R875 VDD2.n73 VDD2.n2 6.59444
R876 VDD2.n151 VDD2.n77 5.81868
R877 VDD2.n146 VDD2.n81 5.81868
R878 VDD2.n106 VDD2.n105 5.81868
R879 VDD2.n28 VDD2.n27 5.81868
R880 VDD2.n69 VDD2.n4 5.81868
R881 VDD2.n74 VDD2.n0 5.81868
R882 VDD2.n143 VDD2.n142 5.04292
R883 VDD2.n109 VDD2.n100 5.04292
R884 VDD2.n31 VDD2.n22 5.04292
R885 VDD2.n66 VDD2.n65 5.04292
R886 VDD2.n139 VDD2.n83 4.26717
R887 VDD2.n110 VDD2.n98 4.26717
R888 VDD2.n32 VDD2.n20 4.26717
R889 VDD2.n62 VDD2.n6 4.26717
R890 VDD2.n138 VDD2.n85 3.49141
R891 VDD2.n114 VDD2.n113 3.49141
R892 VDD2.n36 VDD2.n35 3.49141
R893 VDD2.n61 VDD2.n8 3.49141
R894 VDD2.n135 VDD2.n134 2.71565
R895 VDD2.n117 VDD2.n96 2.71565
R896 VDD2.n39 VDD2.n18 2.71565
R897 VDD2.n58 VDD2.n57 2.71565
R898 VDD2.n104 VDD2.n103 2.41282
R899 VDD2.n26 VDD2.n25 2.41282
R900 VDD2.n131 VDD2.n87 1.93989
R901 VDD2.n118 VDD2.n94 1.93989
R902 VDD2.n40 VDD2.n16 1.93989
R903 VDD2.n54 VDD2.n10 1.93989
R904 VDD2.n130 VDD2.n89 1.16414
R905 VDD2.n122 VDD2.n121 1.16414
R906 VDD2.n45 VDD2.n43 1.16414
R907 VDD2.n53 VDD2.n12 1.16414
R908 VDD2 VDD2.n154 0.440155
R909 VDD2.n127 VDD2.n126 0.388379
R910 VDD2.n93 VDD2.n91 0.388379
R911 VDD2.n44 VDD2.n14 0.388379
R912 VDD2.n50 VDD2.n49 0.388379
R913 VDD2.n152 VDD2.n78 0.155672
R914 VDD2.n145 VDD2.n78 0.155672
R915 VDD2.n145 VDD2.n144 0.155672
R916 VDD2.n144 VDD2.n82 0.155672
R917 VDD2.n137 VDD2.n82 0.155672
R918 VDD2.n137 VDD2.n136 0.155672
R919 VDD2.n136 VDD2.n86 0.155672
R920 VDD2.n129 VDD2.n86 0.155672
R921 VDD2.n129 VDD2.n128 0.155672
R922 VDD2.n128 VDD2.n90 0.155672
R923 VDD2.n120 VDD2.n90 0.155672
R924 VDD2.n120 VDD2.n119 0.155672
R925 VDD2.n119 VDD2.n95 0.155672
R926 VDD2.n112 VDD2.n95 0.155672
R927 VDD2.n112 VDD2.n111 0.155672
R928 VDD2.n111 VDD2.n99 0.155672
R929 VDD2.n104 VDD2.n99 0.155672
R930 VDD2.n26 VDD2.n21 0.155672
R931 VDD2.n33 VDD2.n21 0.155672
R932 VDD2.n34 VDD2.n33 0.155672
R933 VDD2.n34 VDD2.n17 0.155672
R934 VDD2.n41 VDD2.n17 0.155672
R935 VDD2.n42 VDD2.n41 0.155672
R936 VDD2.n42 VDD2.n13 0.155672
R937 VDD2.n51 VDD2.n13 0.155672
R938 VDD2.n52 VDD2.n51 0.155672
R939 VDD2.n52 VDD2.n9 0.155672
R940 VDD2.n59 VDD2.n9 0.155672
R941 VDD2.n60 VDD2.n59 0.155672
R942 VDD2.n60 VDD2.n5 0.155672
R943 VDD2.n67 VDD2.n5 0.155672
R944 VDD2.n68 VDD2.n67 0.155672
R945 VDD2.n68 VDD2.n1 0.155672
R946 VDD2.n75 VDD2.n1 0.155672
R947 B.n339 B.n338 585
R948 B.n337 B.n88 585
R949 B.n336 B.n335 585
R950 B.n334 B.n89 585
R951 B.n333 B.n332 585
R952 B.n331 B.n90 585
R953 B.n330 B.n329 585
R954 B.n328 B.n91 585
R955 B.n327 B.n326 585
R956 B.n325 B.n92 585
R957 B.n324 B.n323 585
R958 B.n322 B.n93 585
R959 B.n321 B.n320 585
R960 B.n319 B.n94 585
R961 B.n318 B.n317 585
R962 B.n316 B.n95 585
R963 B.n315 B.n314 585
R964 B.n313 B.n96 585
R965 B.n312 B.n311 585
R966 B.n310 B.n97 585
R967 B.n309 B.n308 585
R968 B.n307 B.n98 585
R969 B.n306 B.n305 585
R970 B.n304 B.n99 585
R971 B.n303 B.n302 585
R972 B.n301 B.n100 585
R973 B.n300 B.n299 585
R974 B.n298 B.n101 585
R975 B.n297 B.n296 585
R976 B.n295 B.n102 585
R977 B.n294 B.n293 585
R978 B.n292 B.n103 585
R979 B.n291 B.n290 585
R980 B.n289 B.n104 585
R981 B.n288 B.n287 585
R982 B.n286 B.n105 585
R983 B.n285 B.n284 585
R984 B.n283 B.n106 585
R985 B.n282 B.n281 585
R986 B.n280 B.n107 585
R987 B.n279 B.n278 585
R988 B.n277 B.n108 585
R989 B.n276 B.n275 585
R990 B.n274 B.n109 585
R991 B.n273 B.n272 585
R992 B.n271 B.n110 585
R993 B.n270 B.n269 585
R994 B.n268 B.n111 585
R995 B.n266 B.n265 585
R996 B.n264 B.n114 585
R997 B.n263 B.n262 585
R998 B.n261 B.n115 585
R999 B.n260 B.n259 585
R1000 B.n258 B.n116 585
R1001 B.n257 B.n256 585
R1002 B.n255 B.n117 585
R1003 B.n254 B.n253 585
R1004 B.n252 B.n118 585
R1005 B.n251 B.n250 585
R1006 B.n246 B.n119 585
R1007 B.n245 B.n244 585
R1008 B.n243 B.n120 585
R1009 B.n242 B.n241 585
R1010 B.n240 B.n121 585
R1011 B.n239 B.n238 585
R1012 B.n237 B.n122 585
R1013 B.n236 B.n235 585
R1014 B.n234 B.n123 585
R1015 B.n233 B.n232 585
R1016 B.n231 B.n124 585
R1017 B.n230 B.n229 585
R1018 B.n228 B.n125 585
R1019 B.n227 B.n226 585
R1020 B.n225 B.n126 585
R1021 B.n224 B.n223 585
R1022 B.n222 B.n127 585
R1023 B.n221 B.n220 585
R1024 B.n219 B.n128 585
R1025 B.n218 B.n217 585
R1026 B.n216 B.n129 585
R1027 B.n215 B.n214 585
R1028 B.n213 B.n130 585
R1029 B.n212 B.n211 585
R1030 B.n210 B.n131 585
R1031 B.n209 B.n208 585
R1032 B.n207 B.n132 585
R1033 B.n206 B.n205 585
R1034 B.n204 B.n133 585
R1035 B.n203 B.n202 585
R1036 B.n201 B.n134 585
R1037 B.n200 B.n199 585
R1038 B.n198 B.n135 585
R1039 B.n197 B.n196 585
R1040 B.n195 B.n136 585
R1041 B.n194 B.n193 585
R1042 B.n192 B.n137 585
R1043 B.n191 B.n190 585
R1044 B.n189 B.n138 585
R1045 B.n188 B.n187 585
R1046 B.n186 B.n139 585
R1047 B.n185 B.n184 585
R1048 B.n183 B.n140 585
R1049 B.n182 B.n181 585
R1050 B.n180 B.n141 585
R1051 B.n179 B.n178 585
R1052 B.n177 B.n142 585
R1053 B.n340 B.n87 585
R1054 B.n342 B.n341 585
R1055 B.n343 B.n86 585
R1056 B.n345 B.n344 585
R1057 B.n346 B.n85 585
R1058 B.n348 B.n347 585
R1059 B.n349 B.n84 585
R1060 B.n351 B.n350 585
R1061 B.n352 B.n83 585
R1062 B.n354 B.n353 585
R1063 B.n355 B.n82 585
R1064 B.n357 B.n356 585
R1065 B.n358 B.n81 585
R1066 B.n360 B.n359 585
R1067 B.n361 B.n80 585
R1068 B.n363 B.n362 585
R1069 B.n364 B.n79 585
R1070 B.n366 B.n365 585
R1071 B.n367 B.n78 585
R1072 B.n369 B.n368 585
R1073 B.n370 B.n77 585
R1074 B.n372 B.n371 585
R1075 B.n373 B.n76 585
R1076 B.n375 B.n374 585
R1077 B.n376 B.n75 585
R1078 B.n378 B.n377 585
R1079 B.n379 B.n74 585
R1080 B.n381 B.n380 585
R1081 B.n382 B.n73 585
R1082 B.n384 B.n383 585
R1083 B.n385 B.n72 585
R1084 B.n387 B.n386 585
R1085 B.n388 B.n71 585
R1086 B.n390 B.n389 585
R1087 B.n391 B.n70 585
R1088 B.n393 B.n392 585
R1089 B.n394 B.n69 585
R1090 B.n396 B.n395 585
R1091 B.n556 B.n11 585
R1092 B.n555 B.n554 585
R1093 B.n553 B.n12 585
R1094 B.n552 B.n551 585
R1095 B.n550 B.n13 585
R1096 B.n549 B.n548 585
R1097 B.n547 B.n14 585
R1098 B.n546 B.n545 585
R1099 B.n544 B.n15 585
R1100 B.n543 B.n542 585
R1101 B.n541 B.n16 585
R1102 B.n540 B.n539 585
R1103 B.n538 B.n17 585
R1104 B.n537 B.n536 585
R1105 B.n535 B.n18 585
R1106 B.n534 B.n533 585
R1107 B.n532 B.n19 585
R1108 B.n531 B.n530 585
R1109 B.n529 B.n20 585
R1110 B.n528 B.n527 585
R1111 B.n526 B.n21 585
R1112 B.n525 B.n524 585
R1113 B.n523 B.n22 585
R1114 B.n522 B.n521 585
R1115 B.n520 B.n23 585
R1116 B.n519 B.n518 585
R1117 B.n517 B.n24 585
R1118 B.n516 B.n515 585
R1119 B.n514 B.n25 585
R1120 B.n513 B.n512 585
R1121 B.n511 B.n26 585
R1122 B.n510 B.n509 585
R1123 B.n508 B.n27 585
R1124 B.n507 B.n506 585
R1125 B.n505 B.n28 585
R1126 B.n504 B.n503 585
R1127 B.n502 B.n29 585
R1128 B.n501 B.n500 585
R1129 B.n499 B.n30 585
R1130 B.n498 B.n497 585
R1131 B.n496 B.n31 585
R1132 B.n495 B.n494 585
R1133 B.n493 B.n32 585
R1134 B.n492 B.n491 585
R1135 B.n490 B.n33 585
R1136 B.n489 B.n488 585
R1137 B.n487 B.n34 585
R1138 B.n486 B.n485 585
R1139 B.n483 B.n35 585
R1140 B.n482 B.n481 585
R1141 B.n480 B.n38 585
R1142 B.n479 B.n478 585
R1143 B.n477 B.n39 585
R1144 B.n476 B.n475 585
R1145 B.n474 B.n40 585
R1146 B.n473 B.n472 585
R1147 B.n471 B.n41 585
R1148 B.n470 B.n469 585
R1149 B.n468 B.n467 585
R1150 B.n466 B.n45 585
R1151 B.n465 B.n464 585
R1152 B.n463 B.n46 585
R1153 B.n462 B.n461 585
R1154 B.n460 B.n47 585
R1155 B.n459 B.n458 585
R1156 B.n457 B.n48 585
R1157 B.n456 B.n455 585
R1158 B.n454 B.n49 585
R1159 B.n453 B.n452 585
R1160 B.n451 B.n50 585
R1161 B.n450 B.n449 585
R1162 B.n448 B.n51 585
R1163 B.n447 B.n446 585
R1164 B.n445 B.n52 585
R1165 B.n444 B.n443 585
R1166 B.n442 B.n53 585
R1167 B.n441 B.n440 585
R1168 B.n439 B.n54 585
R1169 B.n438 B.n437 585
R1170 B.n436 B.n55 585
R1171 B.n435 B.n434 585
R1172 B.n433 B.n56 585
R1173 B.n432 B.n431 585
R1174 B.n430 B.n57 585
R1175 B.n429 B.n428 585
R1176 B.n427 B.n58 585
R1177 B.n426 B.n425 585
R1178 B.n424 B.n59 585
R1179 B.n423 B.n422 585
R1180 B.n421 B.n60 585
R1181 B.n420 B.n419 585
R1182 B.n418 B.n61 585
R1183 B.n417 B.n416 585
R1184 B.n415 B.n62 585
R1185 B.n414 B.n413 585
R1186 B.n412 B.n63 585
R1187 B.n411 B.n410 585
R1188 B.n409 B.n64 585
R1189 B.n408 B.n407 585
R1190 B.n406 B.n65 585
R1191 B.n405 B.n404 585
R1192 B.n403 B.n66 585
R1193 B.n402 B.n401 585
R1194 B.n400 B.n67 585
R1195 B.n399 B.n398 585
R1196 B.n397 B.n68 585
R1197 B.n558 B.n557 585
R1198 B.n559 B.n10 585
R1199 B.n561 B.n560 585
R1200 B.n562 B.n9 585
R1201 B.n564 B.n563 585
R1202 B.n565 B.n8 585
R1203 B.n567 B.n566 585
R1204 B.n568 B.n7 585
R1205 B.n570 B.n569 585
R1206 B.n571 B.n6 585
R1207 B.n573 B.n572 585
R1208 B.n574 B.n5 585
R1209 B.n576 B.n575 585
R1210 B.n577 B.n4 585
R1211 B.n579 B.n578 585
R1212 B.n580 B.n3 585
R1213 B.n582 B.n581 585
R1214 B.n583 B.n0 585
R1215 B.n2 B.n1 585
R1216 B.n152 B.n151 585
R1217 B.n153 B.n150 585
R1218 B.n155 B.n154 585
R1219 B.n156 B.n149 585
R1220 B.n158 B.n157 585
R1221 B.n159 B.n148 585
R1222 B.n161 B.n160 585
R1223 B.n162 B.n147 585
R1224 B.n164 B.n163 585
R1225 B.n165 B.n146 585
R1226 B.n167 B.n166 585
R1227 B.n168 B.n145 585
R1228 B.n170 B.n169 585
R1229 B.n171 B.n144 585
R1230 B.n173 B.n172 585
R1231 B.n174 B.n143 585
R1232 B.n176 B.n175 585
R1233 B.n177 B.n176 463.671
R1234 B.n338 B.n87 463.671
R1235 B.n397 B.n396 463.671
R1236 B.n558 B.n11 463.671
R1237 B.n112 B.t10 448.926
R1238 B.n42 B.t5 448.926
R1239 B.n247 B.t7 448.926
R1240 B.n36 B.t2 448.926
R1241 B.n247 B.t6 442.192
R1242 B.n112 B.t9 442.192
R1243 B.n42 B.t3 442.192
R1244 B.n36 B.t0 442.192
R1245 B.n113 B.t11 414.599
R1246 B.n43 B.t4 414.599
R1247 B.n248 B.t8 414.599
R1248 B.n37 B.t1 414.599
R1249 B.n585 B.n584 256.663
R1250 B.n584 B.n583 235.042
R1251 B.n584 B.n2 235.042
R1252 B.n178 B.n177 163.367
R1253 B.n178 B.n141 163.367
R1254 B.n182 B.n141 163.367
R1255 B.n183 B.n182 163.367
R1256 B.n184 B.n183 163.367
R1257 B.n184 B.n139 163.367
R1258 B.n188 B.n139 163.367
R1259 B.n189 B.n188 163.367
R1260 B.n190 B.n189 163.367
R1261 B.n190 B.n137 163.367
R1262 B.n194 B.n137 163.367
R1263 B.n195 B.n194 163.367
R1264 B.n196 B.n195 163.367
R1265 B.n196 B.n135 163.367
R1266 B.n200 B.n135 163.367
R1267 B.n201 B.n200 163.367
R1268 B.n202 B.n201 163.367
R1269 B.n202 B.n133 163.367
R1270 B.n206 B.n133 163.367
R1271 B.n207 B.n206 163.367
R1272 B.n208 B.n207 163.367
R1273 B.n208 B.n131 163.367
R1274 B.n212 B.n131 163.367
R1275 B.n213 B.n212 163.367
R1276 B.n214 B.n213 163.367
R1277 B.n214 B.n129 163.367
R1278 B.n218 B.n129 163.367
R1279 B.n219 B.n218 163.367
R1280 B.n220 B.n219 163.367
R1281 B.n220 B.n127 163.367
R1282 B.n224 B.n127 163.367
R1283 B.n225 B.n224 163.367
R1284 B.n226 B.n225 163.367
R1285 B.n226 B.n125 163.367
R1286 B.n230 B.n125 163.367
R1287 B.n231 B.n230 163.367
R1288 B.n232 B.n231 163.367
R1289 B.n232 B.n123 163.367
R1290 B.n236 B.n123 163.367
R1291 B.n237 B.n236 163.367
R1292 B.n238 B.n237 163.367
R1293 B.n238 B.n121 163.367
R1294 B.n242 B.n121 163.367
R1295 B.n243 B.n242 163.367
R1296 B.n244 B.n243 163.367
R1297 B.n244 B.n119 163.367
R1298 B.n251 B.n119 163.367
R1299 B.n252 B.n251 163.367
R1300 B.n253 B.n252 163.367
R1301 B.n253 B.n117 163.367
R1302 B.n257 B.n117 163.367
R1303 B.n258 B.n257 163.367
R1304 B.n259 B.n258 163.367
R1305 B.n259 B.n115 163.367
R1306 B.n263 B.n115 163.367
R1307 B.n264 B.n263 163.367
R1308 B.n265 B.n264 163.367
R1309 B.n265 B.n111 163.367
R1310 B.n270 B.n111 163.367
R1311 B.n271 B.n270 163.367
R1312 B.n272 B.n271 163.367
R1313 B.n272 B.n109 163.367
R1314 B.n276 B.n109 163.367
R1315 B.n277 B.n276 163.367
R1316 B.n278 B.n277 163.367
R1317 B.n278 B.n107 163.367
R1318 B.n282 B.n107 163.367
R1319 B.n283 B.n282 163.367
R1320 B.n284 B.n283 163.367
R1321 B.n284 B.n105 163.367
R1322 B.n288 B.n105 163.367
R1323 B.n289 B.n288 163.367
R1324 B.n290 B.n289 163.367
R1325 B.n290 B.n103 163.367
R1326 B.n294 B.n103 163.367
R1327 B.n295 B.n294 163.367
R1328 B.n296 B.n295 163.367
R1329 B.n296 B.n101 163.367
R1330 B.n300 B.n101 163.367
R1331 B.n301 B.n300 163.367
R1332 B.n302 B.n301 163.367
R1333 B.n302 B.n99 163.367
R1334 B.n306 B.n99 163.367
R1335 B.n307 B.n306 163.367
R1336 B.n308 B.n307 163.367
R1337 B.n308 B.n97 163.367
R1338 B.n312 B.n97 163.367
R1339 B.n313 B.n312 163.367
R1340 B.n314 B.n313 163.367
R1341 B.n314 B.n95 163.367
R1342 B.n318 B.n95 163.367
R1343 B.n319 B.n318 163.367
R1344 B.n320 B.n319 163.367
R1345 B.n320 B.n93 163.367
R1346 B.n324 B.n93 163.367
R1347 B.n325 B.n324 163.367
R1348 B.n326 B.n325 163.367
R1349 B.n326 B.n91 163.367
R1350 B.n330 B.n91 163.367
R1351 B.n331 B.n330 163.367
R1352 B.n332 B.n331 163.367
R1353 B.n332 B.n89 163.367
R1354 B.n336 B.n89 163.367
R1355 B.n337 B.n336 163.367
R1356 B.n338 B.n337 163.367
R1357 B.n396 B.n69 163.367
R1358 B.n392 B.n69 163.367
R1359 B.n392 B.n391 163.367
R1360 B.n391 B.n390 163.367
R1361 B.n390 B.n71 163.367
R1362 B.n386 B.n71 163.367
R1363 B.n386 B.n385 163.367
R1364 B.n385 B.n384 163.367
R1365 B.n384 B.n73 163.367
R1366 B.n380 B.n73 163.367
R1367 B.n380 B.n379 163.367
R1368 B.n379 B.n378 163.367
R1369 B.n378 B.n75 163.367
R1370 B.n374 B.n75 163.367
R1371 B.n374 B.n373 163.367
R1372 B.n373 B.n372 163.367
R1373 B.n372 B.n77 163.367
R1374 B.n368 B.n77 163.367
R1375 B.n368 B.n367 163.367
R1376 B.n367 B.n366 163.367
R1377 B.n366 B.n79 163.367
R1378 B.n362 B.n79 163.367
R1379 B.n362 B.n361 163.367
R1380 B.n361 B.n360 163.367
R1381 B.n360 B.n81 163.367
R1382 B.n356 B.n81 163.367
R1383 B.n356 B.n355 163.367
R1384 B.n355 B.n354 163.367
R1385 B.n354 B.n83 163.367
R1386 B.n350 B.n83 163.367
R1387 B.n350 B.n349 163.367
R1388 B.n349 B.n348 163.367
R1389 B.n348 B.n85 163.367
R1390 B.n344 B.n85 163.367
R1391 B.n344 B.n343 163.367
R1392 B.n343 B.n342 163.367
R1393 B.n342 B.n87 163.367
R1394 B.n554 B.n11 163.367
R1395 B.n554 B.n553 163.367
R1396 B.n553 B.n552 163.367
R1397 B.n552 B.n13 163.367
R1398 B.n548 B.n13 163.367
R1399 B.n548 B.n547 163.367
R1400 B.n547 B.n546 163.367
R1401 B.n546 B.n15 163.367
R1402 B.n542 B.n15 163.367
R1403 B.n542 B.n541 163.367
R1404 B.n541 B.n540 163.367
R1405 B.n540 B.n17 163.367
R1406 B.n536 B.n17 163.367
R1407 B.n536 B.n535 163.367
R1408 B.n535 B.n534 163.367
R1409 B.n534 B.n19 163.367
R1410 B.n530 B.n19 163.367
R1411 B.n530 B.n529 163.367
R1412 B.n529 B.n528 163.367
R1413 B.n528 B.n21 163.367
R1414 B.n524 B.n21 163.367
R1415 B.n524 B.n523 163.367
R1416 B.n523 B.n522 163.367
R1417 B.n522 B.n23 163.367
R1418 B.n518 B.n23 163.367
R1419 B.n518 B.n517 163.367
R1420 B.n517 B.n516 163.367
R1421 B.n516 B.n25 163.367
R1422 B.n512 B.n25 163.367
R1423 B.n512 B.n511 163.367
R1424 B.n511 B.n510 163.367
R1425 B.n510 B.n27 163.367
R1426 B.n506 B.n27 163.367
R1427 B.n506 B.n505 163.367
R1428 B.n505 B.n504 163.367
R1429 B.n504 B.n29 163.367
R1430 B.n500 B.n29 163.367
R1431 B.n500 B.n499 163.367
R1432 B.n499 B.n498 163.367
R1433 B.n498 B.n31 163.367
R1434 B.n494 B.n31 163.367
R1435 B.n494 B.n493 163.367
R1436 B.n493 B.n492 163.367
R1437 B.n492 B.n33 163.367
R1438 B.n488 B.n33 163.367
R1439 B.n488 B.n487 163.367
R1440 B.n487 B.n486 163.367
R1441 B.n486 B.n35 163.367
R1442 B.n481 B.n35 163.367
R1443 B.n481 B.n480 163.367
R1444 B.n480 B.n479 163.367
R1445 B.n479 B.n39 163.367
R1446 B.n475 B.n39 163.367
R1447 B.n475 B.n474 163.367
R1448 B.n474 B.n473 163.367
R1449 B.n473 B.n41 163.367
R1450 B.n469 B.n41 163.367
R1451 B.n469 B.n468 163.367
R1452 B.n468 B.n45 163.367
R1453 B.n464 B.n45 163.367
R1454 B.n464 B.n463 163.367
R1455 B.n463 B.n462 163.367
R1456 B.n462 B.n47 163.367
R1457 B.n458 B.n47 163.367
R1458 B.n458 B.n457 163.367
R1459 B.n457 B.n456 163.367
R1460 B.n456 B.n49 163.367
R1461 B.n452 B.n49 163.367
R1462 B.n452 B.n451 163.367
R1463 B.n451 B.n450 163.367
R1464 B.n450 B.n51 163.367
R1465 B.n446 B.n51 163.367
R1466 B.n446 B.n445 163.367
R1467 B.n445 B.n444 163.367
R1468 B.n444 B.n53 163.367
R1469 B.n440 B.n53 163.367
R1470 B.n440 B.n439 163.367
R1471 B.n439 B.n438 163.367
R1472 B.n438 B.n55 163.367
R1473 B.n434 B.n55 163.367
R1474 B.n434 B.n433 163.367
R1475 B.n433 B.n432 163.367
R1476 B.n432 B.n57 163.367
R1477 B.n428 B.n57 163.367
R1478 B.n428 B.n427 163.367
R1479 B.n427 B.n426 163.367
R1480 B.n426 B.n59 163.367
R1481 B.n422 B.n59 163.367
R1482 B.n422 B.n421 163.367
R1483 B.n421 B.n420 163.367
R1484 B.n420 B.n61 163.367
R1485 B.n416 B.n61 163.367
R1486 B.n416 B.n415 163.367
R1487 B.n415 B.n414 163.367
R1488 B.n414 B.n63 163.367
R1489 B.n410 B.n63 163.367
R1490 B.n410 B.n409 163.367
R1491 B.n409 B.n408 163.367
R1492 B.n408 B.n65 163.367
R1493 B.n404 B.n65 163.367
R1494 B.n404 B.n403 163.367
R1495 B.n403 B.n402 163.367
R1496 B.n402 B.n67 163.367
R1497 B.n398 B.n67 163.367
R1498 B.n398 B.n397 163.367
R1499 B.n559 B.n558 163.367
R1500 B.n560 B.n559 163.367
R1501 B.n560 B.n9 163.367
R1502 B.n564 B.n9 163.367
R1503 B.n565 B.n564 163.367
R1504 B.n566 B.n565 163.367
R1505 B.n566 B.n7 163.367
R1506 B.n570 B.n7 163.367
R1507 B.n571 B.n570 163.367
R1508 B.n572 B.n571 163.367
R1509 B.n572 B.n5 163.367
R1510 B.n576 B.n5 163.367
R1511 B.n577 B.n576 163.367
R1512 B.n578 B.n577 163.367
R1513 B.n578 B.n3 163.367
R1514 B.n582 B.n3 163.367
R1515 B.n583 B.n582 163.367
R1516 B.n152 B.n2 163.367
R1517 B.n153 B.n152 163.367
R1518 B.n154 B.n153 163.367
R1519 B.n154 B.n149 163.367
R1520 B.n158 B.n149 163.367
R1521 B.n159 B.n158 163.367
R1522 B.n160 B.n159 163.367
R1523 B.n160 B.n147 163.367
R1524 B.n164 B.n147 163.367
R1525 B.n165 B.n164 163.367
R1526 B.n166 B.n165 163.367
R1527 B.n166 B.n145 163.367
R1528 B.n170 B.n145 163.367
R1529 B.n171 B.n170 163.367
R1530 B.n172 B.n171 163.367
R1531 B.n172 B.n143 163.367
R1532 B.n176 B.n143 163.367
R1533 B.n249 B.n248 59.5399
R1534 B.n267 B.n113 59.5399
R1535 B.n44 B.n43 59.5399
R1536 B.n484 B.n37 59.5399
R1537 B.n248 B.n247 34.3278
R1538 B.n113 B.n112 34.3278
R1539 B.n43 B.n42 34.3278
R1540 B.n37 B.n36 34.3278
R1541 B.n340 B.n339 30.1273
R1542 B.n557 B.n556 30.1273
R1543 B.n395 B.n68 30.1273
R1544 B.n175 B.n142 30.1273
R1545 B B.n585 18.0485
R1546 B.n557 B.n10 10.6151
R1547 B.n561 B.n10 10.6151
R1548 B.n562 B.n561 10.6151
R1549 B.n563 B.n562 10.6151
R1550 B.n563 B.n8 10.6151
R1551 B.n567 B.n8 10.6151
R1552 B.n568 B.n567 10.6151
R1553 B.n569 B.n568 10.6151
R1554 B.n569 B.n6 10.6151
R1555 B.n573 B.n6 10.6151
R1556 B.n574 B.n573 10.6151
R1557 B.n575 B.n574 10.6151
R1558 B.n575 B.n4 10.6151
R1559 B.n579 B.n4 10.6151
R1560 B.n580 B.n579 10.6151
R1561 B.n581 B.n580 10.6151
R1562 B.n581 B.n0 10.6151
R1563 B.n556 B.n555 10.6151
R1564 B.n555 B.n12 10.6151
R1565 B.n551 B.n12 10.6151
R1566 B.n551 B.n550 10.6151
R1567 B.n550 B.n549 10.6151
R1568 B.n549 B.n14 10.6151
R1569 B.n545 B.n14 10.6151
R1570 B.n545 B.n544 10.6151
R1571 B.n544 B.n543 10.6151
R1572 B.n543 B.n16 10.6151
R1573 B.n539 B.n16 10.6151
R1574 B.n539 B.n538 10.6151
R1575 B.n538 B.n537 10.6151
R1576 B.n537 B.n18 10.6151
R1577 B.n533 B.n18 10.6151
R1578 B.n533 B.n532 10.6151
R1579 B.n532 B.n531 10.6151
R1580 B.n531 B.n20 10.6151
R1581 B.n527 B.n20 10.6151
R1582 B.n527 B.n526 10.6151
R1583 B.n526 B.n525 10.6151
R1584 B.n525 B.n22 10.6151
R1585 B.n521 B.n22 10.6151
R1586 B.n521 B.n520 10.6151
R1587 B.n520 B.n519 10.6151
R1588 B.n519 B.n24 10.6151
R1589 B.n515 B.n24 10.6151
R1590 B.n515 B.n514 10.6151
R1591 B.n514 B.n513 10.6151
R1592 B.n513 B.n26 10.6151
R1593 B.n509 B.n26 10.6151
R1594 B.n509 B.n508 10.6151
R1595 B.n508 B.n507 10.6151
R1596 B.n507 B.n28 10.6151
R1597 B.n503 B.n28 10.6151
R1598 B.n503 B.n502 10.6151
R1599 B.n502 B.n501 10.6151
R1600 B.n501 B.n30 10.6151
R1601 B.n497 B.n30 10.6151
R1602 B.n497 B.n496 10.6151
R1603 B.n496 B.n495 10.6151
R1604 B.n495 B.n32 10.6151
R1605 B.n491 B.n32 10.6151
R1606 B.n491 B.n490 10.6151
R1607 B.n490 B.n489 10.6151
R1608 B.n489 B.n34 10.6151
R1609 B.n485 B.n34 10.6151
R1610 B.n483 B.n482 10.6151
R1611 B.n482 B.n38 10.6151
R1612 B.n478 B.n38 10.6151
R1613 B.n478 B.n477 10.6151
R1614 B.n477 B.n476 10.6151
R1615 B.n476 B.n40 10.6151
R1616 B.n472 B.n40 10.6151
R1617 B.n472 B.n471 10.6151
R1618 B.n471 B.n470 10.6151
R1619 B.n467 B.n466 10.6151
R1620 B.n466 B.n465 10.6151
R1621 B.n465 B.n46 10.6151
R1622 B.n461 B.n46 10.6151
R1623 B.n461 B.n460 10.6151
R1624 B.n460 B.n459 10.6151
R1625 B.n459 B.n48 10.6151
R1626 B.n455 B.n48 10.6151
R1627 B.n455 B.n454 10.6151
R1628 B.n454 B.n453 10.6151
R1629 B.n453 B.n50 10.6151
R1630 B.n449 B.n50 10.6151
R1631 B.n449 B.n448 10.6151
R1632 B.n448 B.n447 10.6151
R1633 B.n447 B.n52 10.6151
R1634 B.n443 B.n52 10.6151
R1635 B.n443 B.n442 10.6151
R1636 B.n442 B.n441 10.6151
R1637 B.n441 B.n54 10.6151
R1638 B.n437 B.n54 10.6151
R1639 B.n437 B.n436 10.6151
R1640 B.n436 B.n435 10.6151
R1641 B.n435 B.n56 10.6151
R1642 B.n431 B.n56 10.6151
R1643 B.n431 B.n430 10.6151
R1644 B.n430 B.n429 10.6151
R1645 B.n429 B.n58 10.6151
R1646 B.n425 B.n58 10.6151
R1647 B.n425 B.n424 10.6151
R1648 B.n424 B.n423 10.6151
R1649 B.n423 B.n60 10.6151
R1650 B.n419 B.n60 10.6151
R1651 B.n419 B.n418 10.6151
R1652 B.n418 B.n417 10.6151
R1653 B.n417 B.n62 10.6151
R1654 B.n413 B.n62 10.6151
R1655 B.n413 B.n412 10.6151
R1656 B.n412 B.n411 10.6151
R1657 B.n411 B.n64 10.6151
R1658 B.n407 B.n64 10.6151
R1659 B.n407 B.n406 10.6151
R1660 B.n406 B.n405 10.6151
R1661 B.n405 B.n66 10.6151
R1662 B.n401 B.n66 10.6151
R1663 B.n401 B.n400 10.6151
R1664 B.n400 B.n399 10.6151
R1665 B.n399 B.n68 10.6151
R1666 B.n395 B.n394 10.6151
R1667 B.n394 B.n393 10.6151
R1668 B.n393 B.n70 10.6151
R1669 B.n389 B.n70 10.6151
R1670 B.n389 B.n388 10.6151
R1671 B.n388 B.n387 10.6151
R1672 B.n387 B.n72 10.6151
R1673 B.n383 B.n72 10.6151
R1674 B.n383 B.n382 10.6151
R1675 B.n382 B.n381 10.6151
R1676 B.n381 B.n74 10.6151
R1677 B.n377 B.n74 10.6151
R1678 B.n377 B.n376 10.6151
R1679 B.n376 B.n375 10.6151
R1680 B.n375 B.n76 10.6151
R1681 B.n371 B.n76 10.6151
R1682 B.n371 B.n370 10.6151
R1683 B.n370 B.n369 10.6151
R1684 B.n369 B.n78 10.6151
R1685 B.n365 B.n78 10.6151
R1686 B.n365 B.n364 10.6151
R1687 B.n364 B.n363 10.6151
R1688 B.n363 B.n80 10.6151
R1689 B.n359 B.n80 10.6151
R1690 B.n359 B.n358 10.6151
R1691 B.n358 B.n357 10.6151
R1692 B.n357 B.n82 10.6151
R1693 B.n353 B.n82 10.6151
R1694 B.n353 B.n352 10.6151
R1695 B.n352 B.n351 10.6151
R1696 B.n351 B.n84 10.6151
R1697 B.n347 B.n84 10.6151
R1698 B.n347 B.n346 10.6151
R1699 B.n346 B.n345 10.6151
R1700 B.n345 B.n86 10.6151
R1701 B.n341 B.n86 10.6151
R1702 B.n341 B.n340 10.6151
R1703 B.n151 B.n1 10.6151
R1704 B.n151 B.n150 10.6151
R1705 B.n155 B.n150 10.6151
R1706 B.n156 B.n155 10.6151
R1707 B.n157 B.n156 10.6151
R1708 B.n157 B.n148 10.6151
R1709 B.n161 B.n148 10.6151
R1710 B.n162 B.n161 10.6151
R1711 B.n163 B.n162 10.6151
R1712 B.n163 B.n146 10.6151
R1713 B.n167 B.n146 10.6151
R1714 B.n168 B.n167 10.6151
R1715 B.n169 B.n168 10.6151
R1716 B.n169 B.n144 10.6151
R1717 B.n173 B.n144 10.6151
R1718 B.n174 B.n173 10.6151
R1719 B.n175 B.n174 10.6151
R1720 B.n179 B.n142 10.6151
R1721 B.n180 B.n179 10.6151
R1722 B.n181 B.n180 10.6151
R1723 B.n181 B.n140 10.6151
R1724 B.n185 B.n140 10.6151
R1725 B.n186 B.n185 10.6151
R1726 B.n187 B.n186 10.6151
R1727 B.n187 B.n138 10.6151
R1728 B.n191 B.n138 10.6151
R1729 B.n192 B.n191 10.6151
R1730 B.n193 B.n192 10.6151
R1731 B.n193 B.n136 10.6151
R1732 B.n197 B.n136 10.6151
R1733 B.n198 B.n197 10.6151
R1734 B.n199 B.n198 10.6151
R1735 B.n199 B.n134 10.6151
R1736 B.n203 B.n134 10.6151
R1737 B.n204 B.n203 10.6151
R1738 B.n205 B.n204 10.6151
R1739 B.n205 B.n132 10.6151
R1740 B.n209 B.n132 10.6151
R1741 B.n210 B.n209 10.6151
R1742 B.n211 B.n210 10.6151
R1743 B.n211 B.n130 10.6151
R1744 B.n215 B.n130 10.6151
R1745 B.n216 B.n215 10.6151
R1746 B.n217 B.n216 10.6151
R1747 B.n217 B.n128 10.6151
R1748 B.n221 B.n128 10.6151
R1749 B.n222 B.n221 10.6151
R1750 B.n223 B.n222 10.6151
R1751 B.n223 B.n126 10.6151
R1752 B.n227 B.n126 10.6151
R1753 B.n228 B.n227 10.6151
R1754 B.n229 B.n228 10.6151
R1755 B.n229 B.n124 10.6151
R1756 B.n233 B.n124 10.6151
R1757 B.n234 B.n233 10.6151
R1758 B.n235 B.n234 10.6151
R1759 B.n235 B.n122 10.6151
R1760 B.n239 B.n122 10.6151
R1761 B.n240 B.n239 10.6151
R1762 B.n241 B.n240 10.6151
R1763 B.n241 B.n120 10.6151
R1764 B.n245 B.n120 10.6151
R1765 B.n246 B.n245 10.6151
R1766 B.n250 B.n246 10.6151
R1767 B.n254 B.n118 10.6151
R1768 B.n255 B.n254 10.6151
R1769 B.n256 B.n255 10.6151
R1770 B.n256 B.n116 10.6151
R1771 B.n260 B.n116 10.6151
R1772 B.n261 B.n260 10.6151
R1773 B.n262 B.n261 10.6151
R1774 B.n262 B.n114 10.6151
R1775 B.n266 B.n114 10.6151
R1776 B.n269 B.n268 10.6151
R1777 B.n269 B.n110 10.6151
R1778 B.n273 B.n110 10.6151
R1779 B.n274 B.n273 10.6151
R1780 B.n275 B.n274 10.6151
R1781 B.n275 B.n108 10.6151
R1782 B.n279 B.n108 10.6151
R1783 B.n280 B.n279 10.6151
R1784 B.n281 B.n280 10.6151
R1785 B.n281 B.n106 10.6151
R1786 B.n285 B.n106 10.6151
R1787 B.n286 B.n285 10.6151
R1788 B.n287 B.n286 10.6151
R1789 B.n287 B.n104 10.6151
R1790 B.n291 B.n104 10.6151
R1791 B.n292 B.n291 10.6151
R1792 B.n293 B.n292 10.6151
R1793 B.n293 B.n102 10.6151
R1794 B.n297 B.n102 10.6151
R1795 B.n298 B.n297 10.6151
R1796 B.n299 B.n298 10.6151
R1797 B.n299 B.n100 10.6151
R1798 B.n303 B.n100 10.6151
R1799 B.n304 B.n303 10.6151
R1800 B.n305 B.n304 10.6151
R1801 B.n305 B.n98 10.6151
R1802 B.n309 B.n98 10.6151
R1803 B.n310 B.n309 10.6151
R1804 B.n311 B.n310 10.6151
R1805 B.n311 B.n96 10.6151
R1806 B.n315 B.n96 10.6151
R1807 B.n316 B.n315 10.6151
R1808 B.n317 B.n316 10.6151
R1809 B.n317 B.n94 10.6151
R1810 B.n321 B.n94 10.6151
R1811 B.n322 B.n321 10.6151
R1812 B.n323 B.n322 10.6151
R1813 B.n323 B.n92 10.6151
R1814 B.n327 B.n92 10.6151
R1815 B.n328 B.n327 10.6151
R1816 B.n329 B.n328 10.6151
R1817 B.n329 B.n90 10.6151
R1818 B.n333 B.n90 10.6151
R1819 B.n334 B.n333 10.6151
R1820 B.n335 B.n334 10.6151
R1821 B.n335 B.n88 10.6151
R1822 B.n339 B.n88 10.6151
R1823 B.n485 B.n484 9.36635
R1824 B.n467 B.n44 9.36635
R1825 B.n250 B.n249 9.36635
R1826 B.n268 B.n267 9.36635
R1827 B.n585 B.n0 8.11757
R1828 B.n585 B.n1 8.11757
R1829 B.n484 B.n483 1.24928
R1830 B.n470 B.n44 1.24928
R1831 B.n249 B.n118 1.24928
R1832 B.n267 B.n266 1.24928
C0 VN VDD2 2.87549f
C1 VDD1 VP 3.00869f
C2 VTAIL VDD1 5.72778f
C3 w_n1678_n3800# VP 2.46163f
C4 VDD1 B 1.70333f
C5 VN VDD1 0.147924f
C6 VTAIL w_n1678_n3800# 3.12256f
C7 w_n1678_n3800# B 8.16034f
C8 VTAIL VP 2.38872f
C9 VDD1 VDD2 0.53991f
C10 VN w_n1678_n3800# 2.25038f
C11 VP B 1.22455f
C12 VN VP 5.30728f
C13 w_n1678_n3800# VDD2 1.81852f
C14 VTAIL B 3.55781f
C15 VN VTAIL 2.37423f
C16 VP VDD2 0.285067f
C17 VN B 0.881914f
C18 VTAIL VDD2 5.76798f
C19 B VDD2 1.72328f
C20 VDD1 w_n1678_n3800# 1.80634f
C21 VDD2 VSUBS 0.869464f
C22 VDD1 VSUBS 3.53013f
C23 VTAIL VSUBS 0.954075f
C24 VN VSUBS 8.07545f
C25 VP VSUBS 1.416988f
C26 B VSUBS 3.219021f
C27 w_n1678_n3800# VSUBS 78.2686f
C28 B.n0 VSUBS 0.005758f
C29 B.n1 VSUBS 0.005758f
C30 B.n2 VSUBS 0.008516f
C31 B.n3 VSUBS 0.006526f
C32 B.n4 VSUBS 0.006526f
C33 B.n5 VSUBS 0.006526f
C34 B.n6 VSUBS 0.006526f
C35 B.n7 VSUBS 0.006526f
C36 B.n8 VSUBS 0.006526f
C37 B.n9 VSUBS 0.006526f
C38 B.n10 VSUBS 0.006526f
C39 B.n11 VSUBS 0.015072f
C40 B.n12 VSUBS 0.006526f
C41 B.n13 VSUBS 0.006526f
C42 B.n14 VSUBS 0.006526f
C43 B.n15 VSUBS 0.006526f
C44 B.n16 VSUBS 0.006526f
C45 B.n17 VSUBS 0.006526f
C46 B.n18 VSUBS 0.006526f
C47 B.n19 VSUBS 0.006526f
C48 B.n20 VSUBS 0.006526f
C49 B.n21 VSUBS 0.006526f
C50 B.n22 VSUBS 0.006526f
C51 B.n23 VSUBS 0.006526f
C52 B.n24 VSUBS 0.006526f
C53 B.n25 VSUBS 0.006526f
C54 B.n26 VSUBS 0.006526f
C55 B.n27 VSUBS 0.006526f
C56 B.n28 VSUBS 0.006526f
C57 B.n29 VSUBS 0.006526f
C58 B.n30 VSUBS 0.006526f
C59 B.n31 VSUBS 0.006526f
C60 B.n32 VSUBS 0.006526f
C61 B.n33 VSUBS 0.006526f
C62 B.n34 VSUBS 0.006526f
C63 B.n35 VSUBS 0.006526f
C64 B.t1 VSUBS 0.242527f
C65 B.t2 VSUBS 0.26149f
C66 B.t0 VSUBS 0.819247f
C67 B.n36 VSUBS 0.383088f
C68 B.n37 VSUBS 0.257297f
C69 B.n38 VSUBS 0.006526f
C70 B.n39 VSUBS 0.006526f
C71 B.n40 VSUBS 0.006526f
C72 B.n41 VSUBS 0.006526f
C73 B.t4 VSUBS 0.24253f
C74 B.t5 VSUBS 0.261492f
C75 B.t3 VSUBS 0.819247f
C76 B.n42 VSUBS 0.383085f
C77 B.n43 VSUBS 0.257294f
C78 B.n44 VSUBS 0.01512f
C79 B.n45 VSUBS 0.006526f
C80 B.n46 VSUBS 0.006526f
C81 B.n47 VSUBS 0.006526f
C82 B.n48 VSUBS 0.006526f
C83 B.n49 VSUBS 0.006526f
C84 B.n50 VSUBS 0.006526f
C85 B.n51 VSUBS 0.006526f
C86 B.n52 VSUBS 0.006526f
C87 B.n53 VSUBS 0.006526f
C88 B.n54 VSUBS 0.006526f
C89 B.n55 VSUBS 0.006526f
C90 B.n56 VSUBS 0.006526f
C91 B.n57 VSUBS 0.006526f
C92 B.n58 VSUBS 0.006526f
C93 B.n59 VSUBS 0.006526f
C94 B.n60 VSUBS 0.006526f
C95 B.n61 VSUBS 0.006526f
C96 B.n62 VSUBS 0.006526f
C97 B.n63 VSUBS 0.006526f
C98 B.n64 VSUBS 0.006526f
C99 B.n65 VSUBS 0.006526f
C100 B.n66 VSUBS 0.006526f
C101 B.n67 VSUBS 0.006526f
C102 B.n68 VSUBS 0.015072f
C103 B.n69 VSUBS 0.006526f
C104 B.n70 VSUBS 0.006526f
C105 B.n71 VSUBS 0.006526f
C106 B.n72 VSUBS 0.006526f
C107 B.n73 VSUBS 0.006526f
C108 B.n74 VSUBS 0.006526f
C109 B.n75 VSUBS 0.006526f
C110 B.n76 VSUBS 0.006526f
C111 B.n77 VSUBS 0.006526f
C112 B.n78 VSUBS 0.006526f
C113 B.n79 VSUBS 0.006526f
C114 B.n80 VSUBS 0.006526f
C115 B.n81 VSUBS 0.006526f
C116 B.n82 VSUBS 0.006526f
C117 B.n83 VSUBS 0.006526f
C118 B.n84 VSUBS 0.006526f
C119 B.n85 VSUBS 0.006526f
C120 B.n86 VSUBS 0.006526f
C121 B.n87 VSUBS 0.01391f
C122 B.n88 VSUBS 0.006526f
C123 B.n89 VSUBS 0.006526f
C124 B.n90 VSUBS 0.006526f
C125 B.n91 VSUBS 0.006526f
C126 B.n92 VSUBS 0.006526f
C127 B.n93 VSUBS 0.006526f
C128 B.n94 VSUBS 0.006526f
C129 B.n95 VSUBS 0.006526f
C130 B.n96 VSUBS 0.006526f
C131 B.n97 VSUBS 0.006526f
C132 B.n98 VSUBS 0.006526f
C133 B.n99 VSUBS 0.006526f
C134 B.n100 VSUBS 0.006526f
C135 B.n101 VSUBS 0.006526f
C136 B.n102 VSUBS 0.006526f
C137 B.n103 VSUBS 0.006526f
C138 B.n104 VSUBS 0.006526f
C139 B.n105 VSUBS 0.006526f
C140 B.n106 VSUBS 0.006526f
C141 B.n107 VSUBS 0.006526f
C142 B.n108 VSUBS 0.006526f
C143 B.n109 VSUBS 0.006526f
C144 B.n110 VSUBS 0.006526f
C145 B.n111 VSUBS 0.006526f
C146 B.t11 VSUBS 0.24253f
C147 B.t10 VSUBS 0.261492f
C148 B.t9 VSUBS 0.819247f
C149 B.n112 VSUBS 0.383085f
C150 B.n113 VSUBS 0.257294f
C151 B.n114 VSUBS 0.006526f
C152 B.n115 VSUBS 0.006526f
C153 B.n116 VSUBS 0.006526f
C154 B.n117 VSUBS 0.006526f
C155 B.n118 VSUBS 0.003647f
C156 B.n119 VSUBS 0.006526f
C157 B.n120 VSUBS 0.006526f
C158 B.n121 VSUBS 0.006526f
C159 B.n122 VSUBS 0.006526f
C160 B.n123 VSUBS 0.006526f
C161 B.n124 VSUBS 0.006526f
C162 B.n125 VSUBS 0.006526f
C163 B.n126 VSUBS 0.006526f
C164 B.n127 VSUBS 0.006526f
C165 B.n128 VSUBS 0.006526f
C166 B.n129 VSUBS 0.006526f
C167 B.n130 VSUBS 0.006526f
C168 B.n131 VSUBS 0.006526f
C169 B.n132 VSUBS 0.006526f
C170 B.n133 VSUBS 0.006526f
C171 B.n134 VSUBS 0.006526f
C172 B.n135 VSUBS 0.006526f
C173 B.n136 VSUBS 0.006526f
C174 B.n137 VSUBS 0.006526f
C175 B.n138 VSUBS 0.006526f
C176 B.n139 VSUBS 0.006526f
C177 B.n140 VSUBS 0.006526f
C178 B.n141 VSUBS 0.006526f
C179 B.n142 VSUBS 0.015072f
C180 B.n143 VSUBS 0.006526f
C181 B.n144 VSUBS 0.006526f
C182 B.n145 VSUBS 0.006526f
C183 B.n146 VSUBS 0.006526f
C184 B.n147 VSUBS 0.006526f
C185 B.n148 VSUBS 0.006526f
C186 B.n149 VSUBS 0.006526f
C187 B.n150 VSUBS 0.006526f
C188 B.n151 VSUBS 0.006526f
C189 B.n152 VSUBS 0.006526f
C190 B.n153 VSUBS 0.006526f
C191 B.n154 VSUBS 0.006526f
C192 B.n155 VSUBS 0.006526f
C193 B.n156 VSUBS 0.006526f
C194 B.n157 VSUBS 0.006526f
C195 B.n158 VSUBS 0.006526f
C196 B.n159 VSUBS 0.006526f
C197 B.n160 VSUBS 0.006526f
C198 B.n161 VSUBS 0.006526f
C199 B.n162 VSUBS 0.006526f
C200 B.n163 VSUBS 0.006526f
C201 B.n164 VSUBS 0.006526f
C202 B.n165 VSUBS 0.006526f
C203 B.n166 VSUBS 0.006526f
C204 B.n167 VSUBS 0.006526f
C205 B.n168 VSUBS 0.006526f
C206 B.n169 VSUBS 0.006526f
C207 B.n170 VSUBS 0.006526f
C208 B.n171 VSUBS 0.006526f
C209 B.n172 VSUBS 0.006526f
C210 B.n173 VSUBS 0.006526f
C211 B.n174 VSUBS 0.006526f
C212 B.n175 VSUBS 0.01391f
C213 B.n176 VSUBS 0.01391f
C214 B.n177 VSUBS 0.015072f
C215 B.n178 VSUBS 0.006526f
C216 B.n179 VSUBS 0.006526f
C217 B.n180 VSUBS 0.006526f
C218 B.n181 VSUBS 0.006526f
C219 B.n182 VSUBS 0.006526f
C220 B.n183 VSUBS 0.006526f
C221 B.n184 VSUBS 0.006526f
C222 B.n185 VSUBS 0.006526f
C223 B.n186 VSUBS 0.006526f
C224 B.n187 VSUBS 0.006526f
C225 B.n188 VSUBS 0.006526f
C226 B.n189 VSUBS 0.006526f
C227 B.n190 VSUBS 0.006526f
C228 B.n191 VSUBS 0.006526f
C229 B.n192 VSUBS 0.006526f
C230 B.n193 VSUBS 0.006526f
C231 B.n194 VSUBS 0.006526f
C232 B.n195 VSUBS 0.006526f
C233 B.n196 VSUBS 0.006526f
C234 B.n197 VSUBS 0.006526f
C235 B.n198 VSUBS 0.006526f
C236 B.n199 VSUBS 0.006526f
C237 B.n200 VSUBS 0.006526f
C238 B.n201 VSUBS 0.006526f
C239 B.n202 VSUBS 0.006526f
C240 B.n203 VSUBS 0.006526f
C241 B.n204 VSUBS 0.006526f
C242 B.n205 VSUBS 0.006526f
C243 B.n206 VSUBS 0.006526f
C244 B.n207 VSUBS 0.006526f
C245 B.n208 VSUBS 0.006526f
C246 B.n209 VSUBS 0.006526f
C247 B.n210 VSUBS 0.006526f
C248 B.n211 VSUBS 0.006526f
C249 B.n212 VSUBS 0.006526f
C250 B.n213 VSUBS 0.006526f
C251 B.n214 VSUBS 0.006526f
C252 B.n215 VSUBS 0.006526f
C253 B.n216 VSUBS 0.006526f
C254 B.n217 VSUBS 0.006526f
C255 B.n218 VSUBS 0.006526f
C256 B.n219 VSUBS 0.006526f
C257 B.n220 VSUBS 0.006526f
C258 B.n221 VSUBS 0.006526f
C259 B.n222 VSUBS 0.006526f
C260 B.n223 VSUBS 0.006526f
C261 B.n224 VSUBS 0.006526f
C262 B.n225 VSUBS 0.006526f
C263 B.n226 VSUBS 0.006526f
C264 B.n227 VSUBS 0.006526f
C265 B.n228 VSUBS 0.006526f
C266 B.n229 VSUBS 0.006526f
C267 B.n230 VSUBS 0.006526f
C268 B.n231 VSUBS 0.006526f
C269 B.n232 VSUBS 0.006526f
C270 B.n233 VSUBS 0.006526f
C271 B.n234 VSUBS 0.006526f
C272 B.n235 VSUBS 0.006526f
C273 B.n236 VSUBS 0.006526f
C274 B.n237 VSUBS 0.006526f
C275 B.n238 VSUBS 0.006526f
C276 B.n239 VSUBS 0.006526f
C277 B.n240 VSUBS 0.006526f
C278 B.n241 VSUBS 0.006526f
C279 B.n242 VSUBS 0.006526f
C280 B.n243 VSUBS 0.006526f
C281 B.n244 VSUBS 0.006526f
C282 B.n245 VSUBS 0.006526f
C283 B.n246 VSUBS 0.006526f
C284 B.t8 VSUBS 0.242527f
C285 B.t7 VSUBS 0.26149f
C286 B.t6 VSUBS 0.819247f
C287 B.n247 VSUBS 0.383088f
C288 B.n248 VSUBS 0.257297f
C289 B.n249 VSUBS 0.01512f
C290 B.n250 VSUBS 0.006142f
C291 B.n251 VSUBS 0.006526f
C292 B.n252 VSUBS 0.006526f
C293 B.n253 VSUBS 0.006526f
C294 B.n254 VSUBS 0.006526f
C295 B.n255 VSUBS 0.006526f
C296 B.n256 VSUBS 0.006526f
C297 B.n257 VSUBS 0.006526f
C298 B.n258 VSUBS 0.006526f
C299 B.n259 VSUBS 0.006526f
C300 B.n260 VSUBS 0.006526f
C301 B.n261 VSUBS 0.006526f
C302 B.n262 VSUBS 0.006526f
C303 B.n263 VSUBS 0.006526f
C304 B.n264 VSUBS 0.006526f
C305 B.n265 VSUBS 0.006526f
C306 B.n266 VSUBS 0.003647f
C307 B.n267 VSUBS 0.01512f
C308 B.n268 VSUBS 0.006142f
C309 B.n269 VSUBS 0.006526f
C310 B.n270 VSUBS 0.006526f
C311 B.n271 VSUBS 0.006526f
C312 B.n272 VSUBS 0.006526f
C313 B.n273 VSUBS 0.006526f
C314 B.n274 VSUBS 0.006526f
C315 B.n275 VSUBS 0.006526f
C316 B.n276 VSUBS 0.006526f
C317 B.n277 VSUBS 0.006526f
C318 B.n278 VSUBS 0.006526f
C319 B.n279 VSUBS 0.006526f
C320 B.n280 VSUBS 0.006526f
C321 B.n281 VSUBS 0.006526f
C322 B.n282 VSUBS 0.006526f
C323 B.n283 VSUBS 0.006526f
C324 B.n284 VSUBS 0.006526f
C325 B.n285 VSUBS 0.006526f
C326 B.n286 VSUBS 0.006526f
C327 B.n287 VSUBS 0.006526f
C328 B.n288 VSUBS 0.006526f
C329 B.n289 VSUBS 0.006526f
C330 B.n290 VSUBS 0.006526f
C331 B.n291 VSUBS 0.006526f
C332 B.n292 VSUBS 0.006526f
C333 B.n293 VSUBS 0.006526f
C334 B.n294 VSUBS 0.006526f
C335 B.n295 VSUBS 0.006526f
C336 B.n296 VSUBS 0.006526f
C337 B.n297 VSUBS 0.006526f
C338 B.n298 VSUBS 0.006526f
C339 B.n299 VSUBS 0.006526f
C340 B.n300 VSUBS 0.006526f
C341 B.n301 VSUBS 0.006526f
C342 B.n302 VSUBS 0.006526f
C343 B.n303 VSUBS 0.006526f
C344 B.n304 VSUBS 0.006526f
C345 B.n305 VSUBS 0.006526f
C346 B.n306 VSUBS 0.006526f
C347 B.n307 VSUBS 0.006526f
C348 B.n308 VSUBS 0.006526f
C349 B.n309 VSUBS 0.006526f
C350 B.n310 VSUBS 0.006526f
C351 B.n311 VSUBS 0.006526f
C352 B.n312 VSUBS 0.006526f
C353 B.n313 VSUBS 0.006526f
C354 B.n314 VSUBS 0.006526f
C355 B.n315 VSUBS 0.006526f
C356 B.n316 VSUBS 0.006526f
C357 B.n317 VSUBS 0.006526f
C358 B.n318 VSUBS 0.006526f
C359 B.n319 VSUBS 0.006526f
C360 B.n320 VSUBS 0.006526f
C361 B.n321 VSUBS 0.006526f
C362 B.n322 VSUBS 0.006526f
C363 B.n323 VSUBS 0.006526f
C364 B.n324 VSUBS 0.006526f
C365 B.n325 VSUBS 0.006526f
C366 B.n326 VSUBS 0.006526f
C367 B.n327 VSUBS 0.006526f
C368 B.n328 VSUBS 0.006526f
C369 B.n329 VSUBS 0.006526f
C370 B.n330 VSUBS 0.006526f
C371 B.n331 VSUBS 0.006526f
C372 B.n332 VSUBS 0.006526f
C373 B.n333 VSUBS 0.006526f
C374 B.n334 VSUBS 0.006526f
C375 B.n335 VSUBS 0.006526f
C376 B.n336 VSUBS 0.006526f
C377 B.n337 VSUBS 0.006526f
C378 B.n338 VSUBS 0.015072f
C379 B.n339 VSUBS 0.014236f
C380 B.n340 VSUBS 0.014746f
C381 B.n341 VSUBS 0.006526f
C382 B.n342 VSUBS 0.006526f
C383 B.n343 VSUBS 0.006526f
C384 B.n344 VSUBS 0.006526f
C385 B.n345 VSUBS 0.006526f
C386 B.n346 VSUBS 0.006526f
C387 B.n347 VSUBS 0.006526f
C388 B.n348 VSUBS 0.006526f
C389 B.n349 VSUBS 0.006526f
C390 B.n350 VSUBS 0.006526f
C391 B.n351 VSUBS 0.006526f
C392 B.n352 VSUBS 0.006526f
C393 B.n353 VSUBS 0.006526f
C394 B.n354 VSUBS 0.006526f
C395 B.n355 VSUBS 0.006526f
C396 B.n356 VSUBS 0.006526f
C397 B.n357 VSUBS 0.006526f
C398 B.n358 VSUBS 0.006526f
C399 B.n359 VSUBS 0.006526f
C400 B.n360 VSUBS 0.006526f
C401 B.n361 VSUBS 0.006526f
C402 B.n362 VSUBS 0.006526f
C403 B.n363 VSUBS 0.006526f
C404 B.n364 VSUBS 0.006526f
C405 B.n365 VSUBS 0.006526f
C406 B.n366 VSUBS 0.006526f
C407 B.n367 VSUBS 0.006526f
C408 B.n368 VSUBS 0.006526f
C409 B.n369 VSUBS 0.006526f
C410 B.n370 VSUBS 0.006526f
C411 B.n371 VSUBS 0.006526f
C412 B.n372 VSUBS 0.006526f
C413 B.n373 VSUBS 0.006526f
C414 B.n374 VSUBS 0.006526f
C415 B.n375 VSUBS 0.006526f
C416 B.n376 VSUBS 0.006526f
C417 B.n377 VSUBS 0.006526f
C418 B.n378 VSUBS 0.006526f
C419 B.n379 VSUBS 0.006526f
C420 B.n380 VSUBS 0.006526f
C421 B.n381 VSUBS 0.006526f
C422 B.n382 VSUBS 0.006526f
C423 B.n383 VSUBS 0.006526f
C424 B.n384 VSUBS 0.006526f
C425 B.n385 VSUBS 0.006526f
C426 B.n386 VSUBS 0.006526f
C427 B.n387 VSUBS 0.006526f
C428 B.n388 VSUBS 0.006526f
C429 B.n389 VSUBS 0.006526f
C430 B.n390 VSUBS 0.006526f
C431 B.n391 VSUBS 0.006526f
C432 B.n392 VSUBS 0.006526f
C433 B.n393 VSUBS 0.006526f
C434 B.n394 VSUBS 0.006526f
C435 B.n395 VSUBS 0.01391f
C436 B.n396 VSUBS 0.01391f
C437 B.n397 VSUBS 0.015072f
C438 B.n398 VSUBS 0.006526f
C439 B.n399 VSUBS 0.006526f
C440 B.n400 VSUBS 0.006526f
C441 B.n401 VSUBS 0.006526f
C442 B.n402 VSUBS 0.006526f
C443 B.n403 VSUBS 0.006526f
C444 B.n404 VSUBS 0.006526f
C445 B.n405 VSUBS 0.006526f
C446 B.n406 VSUBS 0.006526f
C447 B.n407 VSUBS 0.006526f
C448 B.n408 VSUBS 0.006526f
C449 B.n409 VSUBS 0.006526f
C450 B.n410 VSUBS 0.006526f
C451 B.n411 VSUBS 0.006526f
C452 B.n412 VSUBS 0.006526f
C453 B.n413 VSUBS 0.006526f
C454 B.n414 VSUBS 0.006526f
C455 B.n415 VSUBS 0.006526f
C456 B.n416 VSUBS 0.006526f
C457 B.n417 VSUBS 0.006526f
C458 B.n418 VSUBS 0.006526f
C459 B.n419 VSUBS 0.006526f
C460 B.n420 VSUBS 0.006526f
C461 B.n421 VSUBS 0.006526f
C462 B.n422 VSUBS 0.006526f
C463 B.n423 VSUBS 0.006526f
C464 B.n424 VSUBS 0.006526f
C465 B.n425 VSUBS 0.006526f
C466 B.n426 VSUBS 0.006526f
C467 B.n427 VSUBS 0.006526f
C468 B.n428 VSUBS 0.006526f
C469 B.n429 VSUBS 0.006526f
C470 B.n430 VSUBS 0.006526f
C471 B.n431 VSUBS 0.006526f
C472 B.n432 VSUBS 0.006526f
C473 B.n433 VSUBS 0.006526f
C474 B.n434 VSUBS 0.006526f
C475 B.n435 VSUBS 0.006526f
C476 B.n436 VSUBS 0.006526f
C477 B.n437 VSUBS 0.006526f
C478 B.n438 VSUBS 0.006526f
C479 B.n439 VSUBS 0.006526f
C480 B.n440 VSUBS 0.006526f
C481 B.n441 VSUBS 0.006526f
C482 B.n442 VSUBS 0.006526f
C483 B.n443 VSUBS 0.006526f
C484 B.n444 VSUBS 0.006526f
C485 B.n445 VSUBS 0.006526f
C486 B.n446 VSUBS 0.006526f
C487 B.n447 VSUBS 0.006526f
C488 B.n448 VSUBS 0.006526f
C489 B.n449 VSUBS 0.006526f
C490 B.n450 VSUBS 0.006526f
C491 B.n451 VSUBS 0.006526f
C492 B.n452 VSUBS 0.006526f
C493 B.n453 VSUBS 0.006526f
C494 B.n454 VSUBS 0.006526f
C495 B.n455 VSUBS 0.006526f
C496 B.n456 VSUBS 0.006526f
C497 B.n457 VSUBS 0.006526f
C498 B.n458 VSUBS 0.006526f
C499 B.n459 VSUBS 0.006526f
C500 B.n460 VSUBS 0.006526f
C501 B.n461 VSUBS 0.006526f
C502 B.n462 VSUBS 0.006526f
C503 B.n463 VSUBS 0.006526f
C504 B.n464 VSUBS 0.006526f
C505 B.n465 VSUBS 0.006526f
C506 B.n466 VSUBS 0.006526f
C507 B.n467 VSUBS 0.006142f
C508 B.n468 VSUBS 0.006526f
C509 B.n469 VSUBS 0.006526f
C510 B.n470 VSUBS 0.003647f
C511 B.n471 VSUBS 0.006526f
C512 B.n472 VSUBS 0.006526f
C513 B.n473 VSUBS 0.006526f
C514 B.n474 VSUBS 0.006526f
C515 B.n475 VSUBS 0.006526f
C516 B.n476 VSUBS 0.006526f
C517 B.n477 VSUBS 0.006526f
C518 B.n478 VSUBS 0.006526f
C519 B.n479 VSUBS 0.006526f
C520 B.n480 VSUBS 0.006526f
C521 B.n481 VSUBS 0.006526f
C522 B.n482 VSUBS 0.006526f
C523 B.n483 VSUBS 0.003647f
C524 B.n484 VSUBS 0.01512f
C525 B.n485 VSUBS 0.006142f
C526 B.n486 VSUBS 0.006526f
C527 B.n487 VSUBS 0.006526f
C528 B.n488 VSUBS 0.006526f
C529 B.n489 VSUBS 0.006526f
C530 B.n490 VSUBS 0.006526f
C531 B.n491 VSUBS 0.006526f
C532 B.n492 VSUBS 0.006526f
C533 B.n493 VSUBS 0.006526f
C534 B.n494 VSUBS 0.006526f
C535 B.n495 VSUBS 0.006526f
C536 B.n496 VSUBS 0.006526f
C537 B.n497 VSUBS 0.006526f
C538 B.n498 VSUBS 0.006526f
C539 B.n499 VSUBS 0.006526f
C540 B.n500 VSUBS 0.006526f
C541 B.n501 VSUBS 0.006526f
C542 B.n502 VSUBS 0.006526f
C543 B.n503 VSUBS 0.006526f
C544 B.n504 VSUBS 0.006526f
C545 B.n505 VSUBS 0.006526f
C546 B.n506 VSUBS 0.006526f
C547 B.n507 VSUBS 0.006526f
C548 B.n508 VSUBS 0.006526f
C549 B.n509 VSUBS 0.006526f
C550 B.n510 VSUBS 0.006526f
C551 B.n511 VSUBS 0.006526f
C552 B.n512 VSUBS 0.006526f
C553 B.n513 VSUBS 0.006526f
C554 B.n514 VSUBS 0.006526f
C555 B.n515 VSUBS 0.006526f
C556 B.n516 VSUBS 0.006526f
C557 B.n517 VSUBS 0.006526f
C558 B.n518 VSUBS 0.006526f
C559 B.n519 VSUBS 0.006526f
C560 B.n520 VSUBS 0.006526f
C561 B.n521 VSUBS 0.006526f
C562 B.n522 VSUBS 0.006526f
C563 B.n523 VSUBS 0.006526f
C564 B.n524 VSUBS 0.006526f
C565 B.n525 VSUBS 0.006526f
C566 B.n526 VSUBS 0.006526f
C567 B.n527 VSUBS 0.006526f
C568 B.n528 VSUBS 0.006526f
C569 B.n529 VSUBS 0.006526f
C570 B.n530 VSUBS 0.006526f
C571 B.n531 VSUBS 0.006526f
C572 B.n532 VSUBS 0.006526f
C573 B.n533 VSUBS 0.006526f
C574 B.n534 VSUBS 0.006526f
C575 B.n535 VSUBS 0.006526f
C576 B.n536 VSUBS 0.006526f
C577 B.n537 VSUBS 0.006526f
C578 B.n538 VSUBS 0.006526f
C579 B.n539 VSUBS 0.006526f
C580 B.n540 VSUBS 0.006526f
C581 B.n541 VSUBS 0.006526f
C582 B.n542 VSUBS 0.006526f
C583 B.n543 VSUBS 0.006526f
C584 B.n544 VSUBS 0.006526f
C585 B.n545 VSUBS 0.006526f
C586 B.n546 VSUBS 0.006526f
C587 B.n547 VSUBS 0.006526f
C588 B.n548 VSUBS 0.006526f
C589 B.n549 VSUBS 0.006526f
C590 B.n550 VSUBS 0.006526f
C591 B.n551 VSUBS 0.006526f
C592 B.n552 VSUBS 0.006526f
C593 B.n553 VSUBS 0.006526f
C594 B.n554 VSUBS 0.006526f
C595 B.n555 VSUBS 0.006526f
C596 B.n556 VSUBS 0.015072f
C597 B.n557 VSUBS 0.01391f
C598 B.n558 VSUBS 0.01391f
C599 B.n559 VSUBS 0.006526f
C600 B.n560 VSUBS 0.006526f
C601 B.n561 VSUBS 0.006526f
C602 B.n562 VSUBS 0.006526f
C603 B.n563 VSUBS 0.006526f
C604 B.n564 VSUBS 0.006526f
C605 B.n565 VSUBS 0.006526f
C606 B.n566 VSUBS 0.006526f
C607 B.n567 VSUBS 0.006526f
C608 B.n568 VSUBS 0.006526f
C609 B.n569 VSUBS 0.006526f
C610 B.n570 VSUBS 0.006526f
C611 B.n571 VSUBS 0.006526f
C612 B.n572 VSUBS 0.006526f
C613 B.n573 VSUBS 0.006526f
C614 B.n574 VSUBS 0.006526f
C615 B.n575 VSUBS 0.006526f
C616 B.n576 VSUBS 0.006526f
C617 B.n577 VSUBS 0.006526f
C618 B.n578 VSUBS 0.006526f
C619 B.n579 VSUBS 0.006526f
C620 B.n580 VSUBS 0.006526f
C621 B.n581 VSUBS 0.006526f
C622 B.n582 VSUBS 0.006526f
C623 B.n583 VSUBS 0.008516f
C624 B.n584 VSUBS 0.009071f
C625 B.n585 VSUBS 0.018039f
C626 VDD2.n0 VSUBS 0.022192f
C627 VDD2.n1 VSUBS 0.020274f
C628 VDD2.n2 VSUBS 0.010894f
C629 VDD2.n3 VSUBS 0.02575f
C630 VDD2.n4 VSUBS 0.011535f
C631 VDD2.n5 VSUBS 0.020274f
C632 VDD2.n6 VSUBS 0.010894f
C633 VDD2.n7 VSUBS 0.02575f
C634 VDD2.n8 VSUBS 0.011535f
C635 VDD2.n9 VSUBS 0.020274f
C636 VDD2.n10 VSUBS 0.010894f
C637 VDD2.n11 VSUBS 0.02575f
C638 VDD2.n12 VSUBS 0.011535f
C639 VDD2.n13 VSUBS 0.020274f
C640 VDD2.n14 VSUBS 0.011215f
C641 VDD2.n15 VSUBS 0.02575f
C642 VDD2.n16 VSUBS 0.011535f
C643 VDD2.n17 VSUBS 0.020274f
C644 VDD2.n18 VSUBS 0.010894f
C645 VDD2.n19 VSUBS 0.02575f
C646 VDD2.n20 VSUBS 0.011535f
C647 VDD2.n21 VSUBS 0.020274f
C648 VDD2.n22 VSUBS 0.010894f
C649 VDD2.n23 VSUBS 0.019313f
C650 VDD2.n24 VSUBS 0.01937f
C651 VDD2.t1 VSUBS 0.055634f
C652 VDD2.n25 VSUBS 0.179466f
C653 VDD2.n26 VSUBS 1.188f
C654 VDD2.n27 VSUBS 0.010894f
C655 VDD2.n28 VSUBS 0.011535f
C656 VDD2.n29 VSUBS 0.02575f
C657 VDD2.n30 VSUBS 0.02575f
C658 VDD2.n31 VSUBS 0.011535f
C659 VDD2.n32 VSUBS 0.010894f
C660 VDD2.n33 VSUBS 0.020274f
C661 VDD2.n34 VSUBS 0.020274f
C662 VDD2.n35 VSUBS 0.010894f
C663 VDD2.n36 VSUBS 0.011535f
C664 VDD2.n37 VSUBS 0.02575f
C665 VDD2.n38 VSUBS 0.02575f
C666 VDD2.n39 VSUBS 0.011535f
C667 VDD2.n40 VSUBS 0.010894f
C668 VDD2.n41 VSUBS 0.020274f
C669 VDD2.n42 VSUBS 0.020274f
C670 VDD2.n43 VSUBS 0.010894f
C671 VDD2.n44 VSUBS 0.010894f
C672 VDD2.n45 VSUBS 0.011535f
C673 VDD2.n46 VSUBS 0.02575f
C674 VDD2.n47 VSUBS 0.02575f
C675 VDD2.n48 VSUBS 0.02575f
C676 VDD2.n49 VSUBS 0.011215f
C677 VDD2.n50 VSUBS 0.010894f
C678 VDD2.n51 VSUBS 0.020274f
C679 VDD2.n52 VSUBS 0.020274f
C680 VDD2.n53 VSUBS 0.010894f
C681 VDD2.n54 VSUBS 0.011535f
C682 VDD2.n55 VSUBS 0.02575f
C683 VDD2.n56 VSUBS 0.02575f
C684 VDD2.n57 VSUBS 0.011535f
C685 VDD2.n58 VSUBS 0.010894f
C686 VDD2.n59 VSUBS 0.020274f
C687 VDD2.n60 VSUBS 0.020274f
C688 VDD2.n61 VSUBS 0.010894f
C689 VDD2.n62 VSUBS 0.011535f
C690 VDD2.n63 VSUBS 0.02575f
C691 VDD2.n64 VSUBS 0.02575f
C692 VDD2.n65 VSUBS 0.011535f
C693 VDD2.n66 VSUBS 0.010894f
C694 VDD2.n67 VSUBS 0.020274f
C695 VDD2.n68 VSUBS 0.020274f
C696 VDD2.n69 VSUBS 0.010894f
C697 VDD2.n70 VSUBS 0.011535f
C698 VDD2.n71 VSUBS 0.02575f
C699 VDD2.n72 VSUBS 0.062049f
C700 VDD2.n73 VSUBS 0.011535f
C701 VDD2.n74 VSUBS 0.010894f
C702 VDD2.n75 VSUBS 0.043538f
C703 VDD2.n76 VSUBS 0.610654f
C704 VDD2.n77 VSUBS 0.022192f
C705 VDD2.n78 VSUBS 0.020274f
C706 VDD2.n79 VSUBS 0.010894f
C707 VDD2.n80 VSUBS 0.02575f
C708 VDD2.n81 VSUBS 0.011535f
C709 VDD2.n82 VSUBS 0.020274f
C710 VDD2.n83 VSUBS 0.010894f
C711 VDD2.n84 VSUBS 0.02575f
C712 VDD2.n85 VSUBS 0.011535f
C713 VDD2.n86 VSUBS 0.020274f
C714 VDD2.n87 VSUBS 0.010894f
C715 VDD2.n88 VSUBS 0.02575f
C716 VDD2.n89 VSUBS 0.011535f
C717 VDD2.n90 VSUBS 0.020274f
C718 VDD2.n91 VSUBS 0.011215f
C719 VDD2.n92 VSUBS 0.02575f
C720 VDD2.n93 VSUBS 0.010894f
C721 VDD2.n94 VSUBS 0.011535f
C722 VDD2.n95 VSUBS 0.020274f
C723 VDD2.n96 VSUBS 0.010894f
C724 VDD2.n97 VSUBS 0.02575f
C725 VDD2.n98 VSUBS 0.011535f
C726 VDD2.n99 VSUBS 0.020274f
C727 VDD2.n100 VSUBS 0.010894f
C728 VDD2.n101 VSUBS 0.019313f
C729 VDD2.n102 VSUBS 0.01937f
C730 VDD2.t0 VSUBS 0.055634f
C731 VDD2.n103 VSUBS 0.179466f
C732 VDD2.n104 VSUBS 1.188f
C733 VDD2.n105 VSUBS 0.010894f
C734 VDD2.n106 VSUBS 0.011535f
C735 VDD2.n107 VSUBS 0.02575f
C736 VDD2.n108 VSUBS 0.02575f
C737 VDD2.n109 VSUBS 0.011535f
C738 VDD2.n110 VSUBS 0.010894f
C739 VDD2.n111 VSUBS 0.020274f
C740 VDD2.n112 VSUBS 0.020274f
C741 VDD2.n113 VSUBS 0.010894f
C742 VDD2.n114 VSUBS 0.011535f
C743 VDD2.n115 VSUBS 0.02575f
C744 VDD2.n116 VSUBS 0.02575f
C745 VDD2.n117 VSUBS 0.011535f
C746 VDD2.n118 VSUBS 0.010894f
C747 VDD2.n119 VSUBS 0.020274f
C748 VDD2.n120 VSUBS 0.020274f
C749 VDD2.n121 VSUBS 0.010894f
C750 VDD2.n122 VSUBS 0.011535f
C751 VDD2.n123 VSUBS 0.02575f
C752 VDD2.n124 VSUBS 0.02575f
C753 VDD2.n125 VSUBS 0.02575f
C754 VDD2.n126 VSUBS 0.011215f
C755 VDD2.n127 VSUBS 0.010894f
C756 VDD2.n128 VSUBS 0.020274f
C757 VDD2.n129 VSUBS 0.020274f
C758 VDD2.n130 VSUBS 0.010894f
C759 VDD2.n131 VSUBS 0.011535f
C760 VDD2.n132 VSUBS 0.02575f
C761 VDD2.n133 VSUBS 0.02575f
C762 VDD2.n134 VSUBS 0.011535f
C763 VDD2.n135 VSUBS 0.010894f
C764 VDD2.n136 VSUBS 0.020274f
C765 VDD2.n137 VSUBS 0.020274f
C766 VDD2.n138 VSUBS 0.010894f
C767 VDD2.n139 VSUBS 0.011535f
C768 VDD2.n140 VSUBS 0.02575f
C769 VDD2.n141 VSUBS 0.02575f
C770 VDD2.n142 VSUBS 0.011535f
C771 VDD2.n143 VSUBS 0.010894f
C772 VDD2.n144 VSUBS 0.020274f
C773 VDD2.n145 VSUBS 0.020274f
C774 VDD2.n146 VSUBS 0.010894f
C775 VDD2.n147 VSUBS 0.011535f
C776 VDD2.n148 VSUBS 0.02575f
C777 VDD2.n149 VSUBS 0.062049f
C778 VDD2.n150 VSUBS 0.011535f
C779 VDD2.n151 VSUBS 0.010894f
C780 VDD2.n152 VSUBS 0.043538f
C781 VDD2.n153 VSUBS 0.045113f
C782 VDD2.n154 VSUBS 2.45556f
C783 VN.t0 VSUBS 3.24675f
C784 VN.t1 VSUBS 3.60196f
C785 VDD1.n0 VSUBS 0.022002f
C786 VDD1.n1 VSUBS 0.020101f
C787 VDD1.n2 VSUBS 0.010801f
C788 VDD1.n3 VSUBS 0.02553f
C789 VDD1.n4 VSUBS 0.011437f
C790 VDD1.n5 VSUBS 0.020101f
C791 VDD1.n6 VSUBS 0.010801f
C792 VDD1.n7 VSUBS 0.02553f
C793 VDD1.n8 VSUBS 0.011437f
C794 VDD1.n9 VSUBS 0.020101f
C795 VDD1.n10 VSUBS 0.010801f
C796 VDD1.n11 VSUBS 0.02553f
C797 VDD1.n12 VSUBS 0.011437f
C798 VDD1.n13 VSUBS 0.020101f
C799 VDD1.n14 VSUBS 0.011119f
C800 VDD1.n15 VSUBS 0.02553f
C801 VDD1.n16 VSUBS 0.010801f
C802 VDD1.n17 VSUBS 0.011437f
C803 VDD1.n18 VSUBS 0.020101f
C804 VDD1.n19 VSUBS 0.010801f
C805 VDD1.n20 VSUBS 0.02553f
C806 VDD1.n21 VSUBS 0.011437f
C807 VDD1.n22 VSUBS 0.020101f
C808 VDD1.n23 VSUBS 0.010801f
C809 VDD1.n24 VSUBS 0.019148f
C810 VDD1.n25 VSUBS 0.019205f
C811 VDD1.t0 VSUBS 0.055159f
C812 VDD1.n26 VSUBS 0.177935f
C813 VDD1.n27 VSUBS 1.17786f
C814 VDD1.n28 VSUBS 0.010801f
C815 VDD1.n29 VSUBS 0.011437f
C816 VDD1.n30 VSUBS 0.02553f
C817 VDD1.n31 VSUBS 0.02553f
C818 VDD1.n32 VSUBS 0.011437f
C819 VDD1.n33 VSUBS 0.010801f
C820 VDD1.n34 VSUBS 0.020101f
C821 VDD1.n35 VSUBS 0.020101f
C822 VDD1.n36 VSUBS 0.010801f
C823 VDD1.n37 VSUBS 0.011437f
C824 VDD1.n38 VSUBS 0.02553f
C825 VDD1.n39 VSUBS 0.02553f
C826 VDD1.n40 VSUBS 0.011437f
C827 VDD1.n41 VSUBS 0.010801f
C828 VDD1.n42 VSUBS 0.020101f
C829 VDD1.n43 VSUBS 0.020101f
C830 VDD1.n44 VSUBS 0.010801f
C831 VDD1.n45 VSUBS 0.011437f
C832 VDD1.n46 VSUBS 0.02553f
C833 VDD1.n47 VSUBS 0.02553f
C834 VDD1.n48 VSUBS 0.02553f
C835 VDD1.n49 VSUBS 0.011119f
C836 VDD1.n50 VSUBS 0.010801f
C837 VDD1.n51 VSUBS 0.020101f
C838 VDD1.n52 VSUBS 0.020101f
C839 VDD1.n53 VSUBS 0.010801f
C840 VDD1.n54 VSUBS 0.011437f
C841 VDD1.n55 VSUBS 0.02553f
C842 VDD1.n56 VSUBS 0.02553f
C843 VDD1.n57 VSUBS 0.011437f
C844 VDD1.n58 VSUBS 0.010801f
C845 VDD1.n59 VSUBS 0.020101f
C846 VDD1.n60 VSUBS 0.020101f
C847 VDD1.n61 VSUBS 0.010801f
C848 VDD1.n62 VSUBS 0.011437f
C849 VDD1.n63 VSUBS 0.02553f
C850 VDD1.n64 VSUBS 0.02553f
C851 VDD1.n65 VSUBS 0.011437f
C852 VDD1.n66 VSUBS 0.010801f
C853 VDD1.n67 VSUBS 0.020101f
C854 VDD1.n68 VSUBS 0.020101f
C855 VDD1.n69 VSUBS 0.010801f
C856 VDD1.n70 VSUBS 0.011437f
C857 VDD1.n71 VSUBS 0.02553f
C858 VDD1.n72 VSUBS 0.06152f
C859 VDD1.n73 VSUBS 0.011437f
C860 VDD1.n74 VSUBS 0.010801f
C861 VDD1.n75 VSUBS 0.043167f
C862 VDD1.n76 VSUBS 0.045339f
C863 VDD1.n77 VSUBS 0.022002f
C864 VDD1.n78 VSUBS 0.020101f
C865 VDD1.n79 VSUBS 0.010801f
C866 VDD1.n80 VSUBS 0.02553f
C867 VDD1.n81 VSUBS 0.011437f
C868 VDD1.n82 VSUBS 0.020101f
C869 VDD1.n83 VSUBS 0.010801f
C870 VDD1.n84 VSUBS 0.02553f
C871 VDD1.n85 VSUBS 0.011437f
C872 VDD1.n86 VSUBS 0.020101f
C873 VDD1.n87 VSUBS 0.010801f
C874 VDD1.n88 VSUBS 0.02553f
C875 VDD1.n89 VSUBS 0.011437f
C876 VDD1.n90 VSUBS 0.020101f
C877 VDD1.n91 VSUBS 0.011119f
C878 VDD1.n92 VSUBS 0.02553f
C879 VDD1.n93 VSUBS 0.011437f
C880 VDD1.n94 VSUBS 0.020101f
C881 VDD1.n95 VSUBS 0.010801f
C882 VDD1.n96 VSUBS 0.02553f
C883 VDD1.n97 VSUBS 0.011437f
C884 VDD1.n98 VSUBS 0.020101f
C885 VDD1.n99 VSUBS 0.010801f
C886 VDD1.n100 VSUBS 0.019148f
C887 VDD1.n101 VSUBS 0.019205f
C888 VDD1.t1 VSUBS 0.055159f
C889 VDD1.n102 VSUBS 0.177935f
C890 VDD1.n103 VSUBS 1.17786f
C891 VDD1.n104 VSUBS 0.010801f
C892 VDD1.n105 VSUBS 0.011437f
C893 VDD1.n106 VSUBS 0.02553f
C894 VDD1.n107 VSUBS 0.02553f
C895 VDD1.n108 VSUBS 0.011437f
C896 VDD1.n109 VSUBS 0.010801f
C897 VDD1.n110 VSUBS 0.020101f
C898 VDD1.n111 VSUBS 0.020101f
C899 VDD1.n112 VSUBS 0.010801f
C900 VDD1.n113 VSUBS 0.011437f
C901 VDD1.n114 VSUBS 0.02553f
C902 VDD1.n115 VSUBS 0.02553f
C903 VDD1.n116 VSUBS 0.011437f
C904 VDD1.n117 VSUBS 0.010801f
C905 VDD1.n118 VSUBS 0.020101f
C906 VDD1.n119 VSUBS 0.020101f
C907 VDD1.n120 VSUBS 0.010801f
C908 VDD1.n121 VSUBS 0.010801f
C909 VDD1.n122 VSUBS 0.011437f
C910 VDD1.n123 VSUBS 0.02553f
C911 VDD1.n124 VSUBS 0.02553f
C912 VDD1.n125 VSUBS 0.02553f
C913 VDD1.n126 VSUBS 0.011119f
C914 VDD1.n127 VSUBS 0.010801f
C915 VDD1.n128 VSUBS 0.020101f
C916 VDD1.n129 VSUBS 0.020101f
C917 VDD1.n130 VSUBS 0.010801f
C918 VDD1.n131 VSUBS 0.011437f
C919 VDD1.n132 VSUBS 0.02553f
C920 VDD1.n133 VSUBS 0.02553f
C921 VDD1.n134 VSUBS 0.011437f
C922 VDD1.n135 VSUBS 0.010801f
C923 VDD1.n136 VSUBS 0.020101f
C924 VDD1.n137 VSUBS 0.020101f
C925 VDD1.n138 VSUBS 0.010801f
C926 VDD1.n139 VSUBS 0.011437f
C927 VDD1.n140 VSUBS 0.02553f
C928 VDD1.n141 VSUBS 0.02553f
C929 VDD1.n142 VSUBS 0.011437f
C930 VDD1.n143 VSUBS 0.010801f
C931 VDD1.n144 VSUBS 0.020101f
C932 VDD1.n145 VSUBS 0.020101f
C933 VDD1.n146 VSUBS 0.010801f
C934 VDD1.n147 VSUBS 0.011437f
C935 VDD1.n148 VSUBS 0.02553f
C936 VDD1.n149 VSUBS 0.06152f
C937 VDD1.n150 VSUBS 0.011437f
C938 VDD1.n151 VSUBS 0.010801f
C939 VDD1.n152 VSUBS 0.043167f
C940 VDD1.n153 VSUBS 0.638836f
C941 VTAIL.n0 VSUBS 0.031091f
C942 VTAIL.n1 VSUBS 0.028404f
C943 VTAIL.n2 VSUBS 0.015263f
C944 VTAIL.n3 VSUBS 0.036076f
C945 VTAIL.n4 VSUBS 0.016161f
C946 VTAIL.n5 VSUBS 0.028404f
C947 VTAIL.n6 VSUBS 0.015263f
C948 VTAIL.n7 VSUBS 0.036076f
C949 VTAIL.n8 VSUBS 0.016161f
C950 VTAIL.n9 VSUBS 0.028404f
C951 VTAIL.n10 VSUBS 0.015263f
C952 VTAIL.n11 VSUBS 0.036076f
C953 VTAIL.n12 VSUBS 0.016161f
C954 VTAIL.n13 VSUBS 0.028404f
C955 VTAIL.n14 VSUBS 0.015712f
C956 VTAIL.n15 VSUBS 0.036076f
C957 VTAIL.n16 VSUBS 0.016161f
C958 VTAIL.n17 VSUBS 0.028404f
C959 VTAIL.n18 VSUBS 0.015263f
C960 VTAIL.n19 VSUBS 0.036076f
C961 VTAIL.n20 VSUBS 0.016161f
C962 VTAIL.n21 VSUBS 0.028404f
C963 VTAIL.n22 VSUBS 0.015263f
C964 VTAIL.n23 VSUBS 0.027057f
C965 VTAIL.n24 VSUBS 0.027138f
C966 VTAIL.t2 VSUBS 0.077944f
C967 VTAIL.n25 VSUBS 0.251434f
C968 VTAIL.n26 VSUBS 1.66439f
C969 VTAIL.n27 VSUBS 0.015263f
C970 VTAIL.n28 VSUBS 0.016161f
C971 VTAIL.n29 VSUBS 0.036076f
C972 VTAIL.n30 VSUBS 0.036076f
C973 VTAIL.n31 VSUBS 0.016161f
C974 VTAIL.n32 VSUBS 0.015263f
C975 VTAIL.n33 VSUBS 0.028404f
C976 VTAIL.n34 VSUBS 0.028404f
C977 VTAIL.n35 VSUBS 0.015263f
C978 VTAIL.n36 VSUBS 0.016161f
C979 VTAIL.n37 VSUBS 0.036076f
C980 VTAIL.n38 VSUBS 0.036076f
C981 VTAIL.n39 VSUBS 0.016161f
C982 VTAIL.n40 VSUBS 0.015263f
C983 VTAIL.n41 VSUBS 0.028404f
C984 VTAIL.n42 VSUBS 0.028404f
C985 VTAIL.n43 VSUBS 0.015263f
C986 VTAIL.n44 VSUBS 0.015263f
C987 VTAIL.n45 VSUBS 0.016161f
C988 VTAIL.n46 VSUBS 0.036076f
C989 VTAIL.n47 VSUBS 0.036076f
C990 VTAIL.n48 VSUBS 0.036076f
C991 VTAIL.n49 VSUBS 0.015712f
C992 VTAIL.n50 VSUBS 0.015263f
C993 VTAIL.n51 VSUBS 0.028404f
C994 VTAIL.n52 VSUBS 0.028404f
C995 VTAIL.n53 VSUBS 0.015263f
C996 VTAIL.n54 VSUBS 0.016161f
C997 VTAIL.n55 VSUBS 0.036076f
C998 VTAIL.n56 VSUBS 0.036076f
C999 VTAIL.n57 VSUBS 0.016161f
C1000 VTAIL.n58 VSUBS 0.015263f
C1001 VTAIL.n59 VSUBS 0.028404f
C1002 VTAIL.n60 VSUBS 0.028404f
C1003 VTAIL.n61 VSUBS 0.015263f
C1004 VTAIL.n62 VSUBS 0.016161f
C1005 VTAIL.n63 VSUBS 0.036076f
C1006 VTAIL.n64 VSUBS 0.036076f
C1007 VTAIL.n65 VSUBS 0.016161f
C1008 VTAIL.n66 VSUBS 0.015263f
C1009 VTAIL.n67 VSUBS 0.028404f
C1010 VTAIL.n68 VSUBS 0.028404f
C1011 VTAIL.n69 VSUBS 0.015263f
C1012 VTAIL.n70 VSUBS 0.016161f
C1013 VTAIL.n71 VSUBS 0.036076f
C1014 VTAIL.n72 VSUBS 0.086932f
C1015 VTAIL.n73 VSUBS 0.016161f
C1016 VTAIL.n74 VSUBS 0.015263f
C1017 VTAIL.n75 VSUBS 0.060998f
C1018 VTAIL.n76 VSUBS 0.043551f
C1019 VTAIL.n77 VSUBS 1.88722f
C1020 VTAIL.n78 VSUBS 0.031091f
C1021 VTAIL.n79 VSUBS 0.028404f
C1022 VTAIL.n80 VSUBS 0.015263f
C1023 VTAIL.n81 VSUBS 0.036076f
C1024 VTAIL.n82 VSUBS 0.016161f
C1025 VTAIL.n83 VSUBS 0.028404f
C1026 VTAIL.n84 VSUBS 0.015263f
C1027 VTAIL.n85 VSUBS 0.036076f
C1028 VTAIL.n86 VSUBS 0.016161f
C1029 VTAIL.n87 VSUBS 0.028404f
C1030 VTAIL.n88 VSUBS 0.015263f
C1031 VTAIL.n89 VSUBS 0.036076f
C1032 VTAIL.n90 VSUBS 0.016161f
C1033 VTAIL.n91 VSUBS 0.028404f
C1034 VTAIL.n92 VSUBS 0.015712f
C1035 VTAIL.n93 VSUBS 0.036076f
C1036 VTAIL.n94 VSUBS 0.015263f
C1037 VTAIL.n95 VSUBS 0.016161f
C1038 VTAIL.n96 VSUBS 0.028404f
C1039 VTAIL.n97 VSUBS 0.015263f
C1040 VTAIL.n98 VSUBS 0.036076f
C1041 VTAIL.n99 VSUBS 0.016161f
C1042 VTAIL.n100 VSUBS 0.028404f
C1043 VTAIL.n101 VSUBS 0.015263f
C1044 VTAIL.n102 VSUBS 0.027057f
C1045 VTAIL.n103 VSUBS 0.027138f
C1046 VTAIL.t0 VSUBS 0.077944f
C1047 VTAIL.n104 VSUBS 0.251434f
C1048 VTAIL.n105 VSUBS 1.66439f
C1049 VTAIL.n106 VSUBS 0.015263f
C1050 VTAIL.n107 VSUBS 0.016161f
C1051 VTAIL.n108 VSUBS 0.036076f
C1052 VTAIL.n109 VSUBS 0.036076f
C1053 VTAIL.n110 VSUBS 0.016161f
C1054 VTAIL.n111 VSUBS 0.015263f
C1055 VTAIL.n112 VSUBS 0.028404f
C1056 VTAIL.n113 VSUBS 0.028404f
C1057 VTAIL.n114 VSUBS 0.015263f
C1058 VTAIL.n115 VSUBS 0.016161f
C1059 VTAIL.n116 VSUBS 0.036076f
C1060 VTAIL.n117 VSUBS 0.036076f
C1061 VTAIL.n118 VSUBS 0.016161f
C1062 VTAIL.n119 VSUBS 0.015263f
C1063 VTAIL.n120 VSUBS 0.028404f
C1064 VTAIL.n121 VSUBS 0.028404f
C1065 VTAIL.n122 VSUBS 0.015263f
C1066 VTAIL.n123 VSUBS 0.016161f
C1067 VTAIL.n124 VSUBS 0.036076f
C1068 VTAIL.n125 VSUBS 0.036076f
C1069 VTAIL.n126 VSUBS 0.036076f
C1070 VTAIL.n127 VSUBS 0.015712f
C1071 VTAIL.n128 VSUBS 0.015263f
C1072 VTAIL.n129 VSUBS 0.028404f
C1073 VTAIL.n130 VSUBS 0.028404f
C1074 VTAIL.n131 VSUBS 0.015263f
C1075 VTAIL.n132 VSUBS 0.016161f
C1076 VTAIL.n133 VSUBS 0.036076f
C1077 VTAIL.n134 VSUBS 0.036076f
C1078 VTAIL.n135 VSUBS 0.016161f
C1079 VTAIL.n136 VSUBS 0.015263f
C1080 VTAIL.n137 VSUBS 0.028404f
C1081 VTAIL.n138 VSUBS 0.028404f
C1082 VTAIL.n139 VSUBS 0.015263f
C1083 VTAIL.n140 VSUBS 0.016161f
C1084 VTAIL.n141 VSUBS 0.036076f
C1085 VTAIL.n142 VSUBS 0.036076f
C1086 VTAIL.n143 VSUBS 0.016161f
C1087 VTAIL.n144 VSUBS 0.015263f
C1088 VTAIL.n145 VSUBS 0.028404f
C1089 VTAIL.n146 VSUBS 0.028404f
C1090 VTAIL.n147 VSUBS 0.015263f
C1091 VTAIL.n148 VSUBS 0.016161f
C1092 VTAIL.n149 VSUBS 0.036076f
C1093 VTAIL.n150 VSUBS 0.086932f
C1094 VTAIL.n151 VSUBS 0.016161f
C1095 VTAIL.n152 VSUBS 0.015263f
C1096 VTAIL.n153 VSUBS 0.060998f
C1097 VTAIL.n154 VSUBS 0.043551f
C1098 VTAIL.n155 VSUBS 1.91681f
C1099 VTAIL.n156 VSUBS 0.031091f
C1100 VTAIL.n157 VSUBS 0.028404f
C1101 VTAIL.n158 VSUBS 0.015263f
C1102 VTAIL.n159 VSUBS 0.036076f
C1103 VTAIL.n160 VSUBS 0.016161f
C1104 VTAIL.n161 VSUBS 0.028404f
C1105 VTAIL.n162 VSUBS 0.015263f
C1106 VTAIL.n163 VSUBS 0.036076f
C1107 VTAIL.n164 VSUBS 0.016161f
C1108 VTAIL.n165 VSUBS 0.028404f
C1109 VTAIL.n166 VSUBS 0.015263f
C1110 VTAIL.n167 VSUBS 0.036076f
C1111 VTAIL.n168 VSUBS 0.016161f
C1112 VTAIL.n169 VSUBS 0.028404f
C1113 VTAIL.n170 VSUBS 0.015712f
C1114 VTAIL.n171 VSUBS 0.036076f
C1115 VTAIL.n172 VSUBS 0.015263f
C1116 VTAIL.n173 VSUBS 0.016161f
C1117 VTAIL.n174 VSUBS 0.028404f
C1118 VTAIL.n175 VSUBS 0.015263f
C1119 VTAIL.n176 VSUBS 0.036076f
C1120 VTAIL.n177 VSUBS 0.016161f
C1121 VTAIL.n178 VSUBS 0.028404f
C1122 VTAIL.n179 VSUBS 0.015263f
C1123 VTAIL.n180 VSUBS 0.027057f
C1124 VTAIL.n181 VSUBS 0.027138f
C1125 VTAIL.t3 VSUBS 0.077944f
C1126 VTAIL.n182 VSUBS 0.251434f
C1127 VTAIL.n183 VSUBS 1.66439f
C1128 VTAIL.n184 VSUBS 0.015263f
C1129 VTAIL.n185 VSUBS 0.016161f
C1130 VTAIL.n186 VSUBS 0.036076f
C1131 VTAIL.n187 VSUBS 0.036076f
C1132 VTAIL.n188 VSUBS 0.016161f
C1133 VTAIL.n189 VSUBS 0.015263f
C1134 VTAIL.n190 VSUBS 0.028404f
C1135 VTAIL.n191 VSUBS 0.028404f
C1136 VTAIL.n192 VSUBS 0.015263f
C1137 VTAIL.n193 VSUBS 0.016161f
C1138 VTAIL.n194 VSUBS 0.036076f
C1139 VTAIL.n195 VSUBS 0.036076f
C1140 VTAIL.n196 VSUBS 0.016161f
C1141 VTAIL.n197 VSUBS 0.015263f
C1142 VTAIL.n198 VSUBS 0.028404f
C1143 VTAIL.n199 VSUBS 0.028404f
C1144 VTAIL.n200 VSUBS 0.015263f
C1145 VTAIL.n201 VSUBS 0.016161f
C1146 VTAIL.n202 VSUBS 0.036076f
C1147 VTAIL.n203 VSUBS 0.036076f
C1148 VTAIL.n204 VSUBS 0.036076f
C1149 VTAIL.n205 VSUBS 0.015712f
C1150 VTAIL.n206 VSUBS 0.015263f
C1151 VTAIL.n207 VSUBS 0.028404f
C1152 VTAIL.n208 VSUBS 0.028404f
C1153 VTAIL.n209 VSUBS 0.015263f
C1154 VTAIL.n210 VSUBS 0.016161f
C1155 VTAIL.n211 VSUBS 0.036076f
C1156 VTAIL.n212 VSUBS 0.036076f
C1157 VTAIL.n213 VSUBS 0.016161f
C1158 VTAIL.n214 VSUBS 0.015263f
C1159 VTAIL.n215 VSUBS 0.028404f
C1160 VTAIL.n216 VSUBS 0.028404f
C1161 VTAIL.n217 VSUBS 0.015263f
C1162 VTAIL.n218 VSUBS 0.016161f
C1163 VTAIL.n219 VSUBS 0.036076f
C1164 VTAIL.n220 VSUBS 0.036076f
C1165 VTAIL.n221 VSUBS 0.016161f
C1166 VTAIL.n222 VSUBS 0.015263f
C1167 VTAIL.n223 VSUBS 0.028404f
C1168 VTAIL.n224 VSUBS 0.028404f
C1169 VTAIL.n225 VSUBS 0.015263f
C1170 VTAIL.n226 VSUBS 0.016161f
C1171 VTAIL.n227 VSUBS 0.036076f
C1172 VTAIL.n228 VSUBS 0.086932f
C1173 VTAIL.n229 VSUBS 0.016161f
C1174 VTAIL.n230 VSUBS 0.015263f
C1175 VTAIL.n231 VSUBS 0.060998f
C1176 VTAIL.n232 VSUBS 0.043551f
C1177 VTAIL.n233 VSUBS 1.77716f
C1178 VTAIL.n234 VSUBS 0.031091f
C1179 VTAIL.n235 VSUBS 0.028404f
C1180 VTAIL.n236 VSUBS 0.015263f
C1181 VTAIL.n237 VSUBS 0.036076f
C1182 VTAIL.n238 VSUBS 0.016161f
C1183 VTAIL.n239 VSUBS 0.028404f
C1184 VTAIL.n240 VSUBS 0.015263f
C1185 VTAIL.n241 VSUBS 0.036076f
C1186 VTAIL.n242 VSUBS 0.016161f
C1187 VTAIL.n243 VSUBS 0.028404f
C1188 VTAIL.n244 VSUBS 0.015263f
C1189 VTAIL.n245 VSUBS 0.036076f
C1190 VTAIL.n246 VSUBS 0.016161f
C1191 VTAIL.n247 VSUBS 0.028404f
C1192 VTAIL.n248 VSUBS 0.015712f
C1193 VTAIL.n249 VSUBS 0.036076f
C1194 VTAIL.n250 VSUBS 0.016161f
C1195 VTAIL.n251 VSUBS 0.028404f
C1196 VTAIL.n252 VSUBS 0.015263f
C1197 VTAIL.n253 VSUBS 0.036076f
C1198 VTAIL.n254 VSUBS 0.016161f
C1199 VTAIL.n255 VSUBS 0.028404f
C1200 VTAIL.n256 VSUBS 0.015263f
C1201 VTAIL.n257 VSUBS 0.027057f
C1202 VTAIL.n258 VSUBS 0.027138f
C1203 VTAIL.t1 VSUBS 0.077944f
C1204 VTAIL.n259 VSUBS 0.251434f
C1205 VTAIL.n260 VSUBS 1.66439f
C1206 VTAIL.n261 VSUBS 0.015263f
C1207 VTAIL.n262 VSUBS 0.016161f
C1208 VTAIL.n263 VSUBS 0.036076f
C1209 VTAIL.n264 VSUBS 0.036076f
C1210 VTAIL.n265 VSUBS 0.016161f
C1211 VTAIL.n266 VSUBS 0.015263f
C1212 VTAIL.n267 VSUBS 0.028404f
C1213 VTAIL.n268 VSUBS 0.028404f
C1214 VTAIL.n269 VSUBS 0.015263f
C1215 VTAIL.n270 VSUBS 0.016161f
C1216 VTAIL.n271 VSUBS 0.036076f
C1217 VTAIL.n272 VSUBS 0.036076f
C1218 VTAIL.n273 VSUBS 0.016161f
C1219 VTAIL.n274 VSUBS 0.015263f
C1220 VTAIL.n275 VSUBS 0.028404f
C1221 VTAIL.n276 VSUBS 0.028404f
C1222 VTAIL.n277 VSUBS 0.015263f
C1223 VTAIL.n278 VSUBS 0.015263f
C1224 VTAIL.n279 VSUBS 0.016161f
C1225 VTAIL.n280 VSUBS 0.036076f
C1226 VTAIL.n281 VSUBS 0.036076f
C1227 VTAIL.n282 VSUBS 0.036076f
C1228 VTAIL.n283 VSUBS 0.015712f
C1229 VTAIL.n284 VSUBS 0.015263f
C1230 VTAIL.n285 VSUBS 0.028404f
C1231 VTAIL.n286 VSUBS 0.028404f
C1232 VTAIL.n287 VSUBS 0.015263f
C1233 VTAIL.n288 VSUBS 0.016161f
C1234 VTAIL.n289 VSUBS 0.036076f
C1235 VTAIL.n290 VSUBS 0.036076f
C1236 VTAIL.n291 VSUBS 0.016161f
C1237 VTAIL.n292 VSUBS 0.015263f
C1238 VTAIL.n293 VSUBS 0.028404f
C1239 VTAIL.n294 VSUBS 0.028404f
C1240 VTAIL.n295 VSUBS 0.015263f
C1241 VTAIL.n296 VSUBS 0.016161f
C1242 VTAIL.n297 VSUBS 0.036076f
C1243 VTAIL.n298 VSUBS 0.036076f
C1244 VTAIL.n299 VSUBS 0.016161f
C1245 VTAIL.n300 VSUBS 0.015263f
C1246 VTAIL.n301 VSUBS 0.028404f
C1247 VTAIL.n302 VSUBS 0.028404f
C1248 VTAIL.n303 VSUBS 0.015263f
C1249 VTAIL.n304 VSUBS 0.016161f
C1250 VTAIL.n305 VSUBS 0.036076f
C1251 VTAIL.n306 VSUBS 0.086932f
C1252 VTAIL.n307 VSUBS 0.016161f
C1253 VTAIL.n308 VSUBS 0.015263f
C1254 VTAIL.n309 VSUBS 0.060998f
C1255 VTAIL.n310 VSUBS 0.043551f
C1256 VTAIL.n311 VSUBS 1.69392f
C1257 VP.t1 VSUBS 3.70106f
C1258 VP.t0 VSUBS 3.34055f
C1259 VP.n0 VSUBS 6.10549f
.ends

