* NGSPICE file created from diff_pair_sample_1068.ext - technology: sky130A

.subckt diff_pair_sample_1068 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t8 VN.t0 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=0.70455 ps=4.6 w=4.27 l=3.97
X1 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0 ps=0 w=4.27 l=3.97
X2 VTAIL.t7 VN.t1 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=0.70455 ps=4.6 w=4.27 l=3.97
X3 VTAIL.t1 VP.t0 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=0.70455 ps=4.6 w=4.27 l=3.97
X4 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0.70455 ps=4.6 w=4.27 l=3.97
X5 VDD2.t4 VN.t2 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=1.6653 ps=9.32 w=4.27 l=3.97
X6 VDD2.t1 VN.t3 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0.70455 ps=4.6 w=4.27 l=3.97
X7 VDD1.t3 VP.t2 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=1.6653 ps=9.32 w=4.27 l=3.97
X8 VDD2.t0 VN.t4 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0.70455 ps=4.6 w=4.27 l=3.97
X9 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0 ps=0 w=4.27 l=3.97
X10 VDD1.t2 VP.t3 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0.70455 ps=4.6 w=4.27 l=3.97
X11 VTAIL.t10 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=0.70455 ps=4.6 w=4.27 l=3.97
X12 VDD2.t3 VN.t5 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=1.6653 ps=9.32 w=4.27 l=3.97
X13 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.70455 pd=4.6 as=1.6653 ps=9.32 w=4.27 l=3.97
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0 ps=0 w=4.27 l=3.97
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.6653 pd=9.32 as=0 ps=0 w=4.27 l=3.97
R0 VN.n42 VN.n41 161.3
R1 VN.n40 VN.n23 161.3
R2 VN.n39 VN.n38 161.3
R3 VN.n37 VN.n24 161.3
R4 VN.n36 VN.n35 161.3
R5 VN.n34 VN.n25 161.3
R6 VN.n33 VN.n32 161.3
R7 VN.n31 VN.n26 161.3
R8 VN.n30 VN.n29 161.3
R9 VN.n20 VN.n19 161.3
R10 VN.n18 VN.n1 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n2 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n12 VN.n3 161.3
R15 VN.n11 VN.n10 161.3
R16 VN.n9 VN.n4 161.3
R17 VN.n8 VN.n7 161.3
R18 VN.n21 VN.n0 87.6207
R19 VN.n43 VN.n22 87.6207
R20 VN.n28 VN.n27 62.9379
R21 VN.n6 VN.n5 62.9379
R22 VN.n27 VN.t5 58.6116
R23 VN.n5 VN.t4 58.6116
R24 VN.n13 VN.n12 50.2061
R25 VN.n35 VN.n34 50.2061
R26 VN VN.n43 48.445
R27 VN.n13 VN.n2 30.7807
R28 VN.n35 VN.n24 30.7807
R29 VN.n6 VN.t1 25.9217
R30 VN.n0 VN.t2 25.9217
R31 VN.n28 VN.t0 25.9217
R32 VN.n22 VN.t3 25.9217
R33 VN.n7 VN.n4 24.4675
R34 VN.n11 VN.n4 24.4675
R35 VN.n12 VN.n11 24.4675
R36 VN.n17 VN.n2 24.4675
R37 VN.n18 VN.n17 24.4675
R38 VN.n19 VN.n18 24.4675
R39 VN.n34 VN.n33 24.4675
R40 VN.n33 VN.n26 24.4675
R41 VN.n29 VN.n26 24.4675
R42 VN.n41 VN.n40 24.4675
R43 VN.n40 VN.n39 24.4675
R44 VN.n39 VN.n24 24.4675
R45 VN.n7 VN.n6 12.234
R46 VN.n29 VN.n28 12.234
R47 VN.n30 VN.n27 2.47757
R48 VN.n8 VN.n5 2.47757
R49 VN.n19 VN.n0 2.4472
R50 VN.n41 VN.n22 2.4472
R51 VN.n43 VN.n42 0.354971
R52 VN.n21 VN.n20 0.354971
R53 VN VN.n21 0.26696
R54 VN.n42 VN.n23 0.189894
R55 VN.n38 VN.n23 0.189894
R56 VN.n38 VN.n37 0.189894
R57 VN.n37 VN.n36 0.189894
R58 VN.n36 VN.n25 0.189894
R59 VN.n32 VN.n25 0.189894
R60 VN.n32 VN.n31 0.189894
R61 VN.n31 VN.n30 0.189894
R62 VN.n9 VN.n8 0.189894
R63 VN.n10 VN.n9 0.189894
R64 VN.n10 VN.n3 0.189894
R65 VN.n14 VN.n3 0.189894
R66 VN.n15 VN.n14 0.189894
R67 VN.n16 VN.n15 0.189894
R68 VN.n16 VN.n1 0.189894
R69 VN.n20 VN.n1 0.189894
R70 VDD2.n1 VDD2.t0 80.6376
R71 VDD2.n2 VDD2.t1 77.913
R72 VDD2.n1 VDD2.n0 74.1472
R73 VDD2 VDD2.n3 74.1444
R74 VDD2.n2 VDD2.n1 39.4437
R75 VDD2.n3 VDD2.t2 4.6375
R76 VDD2.n3 VDD2.t3 4.6375
R77 VDD2.n0 VDD2.t5 4.6375
R78 VDD2.n0 VDD2.t4 4.6375
R79 VDD2 VDD2.n2 2.83886
R80 VTAIL.n7 VTAIL.t3 61.2342
R81 VTAIL.n11 VTAIL.t6 61.234
R82 VTAIL.n2 VTAIL.t0 61.234
R83 VTAIL.n10 VTAIL.t9 61.234
R84 VTAIL.n9 VTAIL.n8 56.5972
R85 VTAIL.n6 VTAIL.n5 56.5972
R86 VTAIL.n1 VTAIL.n0 56.597
R87 VTAIL.n4 VTAIL.n3 56.597
R88 VTAIL.n6 VTAIL.n4 23.4617
R89 VTAIL.n11 VTAIL.n10 19.7548
R90 VTAIL.n0 VTAIL.t4 4.6375
R91 VTAIL.n0 VTAIL.t7 4.6375
R92 VTAIL.n3 VTAIL.t11 4.6375
R93 VTAIL.n3 VTAIL.t10 4.6375
R94 VTAIL.n8 VTAIL.t2 4.6375
R95 VTAIL.n8 VTAIL.t1 4.6375
R96 VTAIL.n5 VTAIL.t5 4.6375
R97 VTAIL.n5 VTAIL.t8 4.6375
R98 VTAIL.n7 VTAIL.n6 3.7074
R99 VTAIL.n10 VTAIL.n9 3.7074
R100 VTAIL.n4 VTAIL.n2 3.7074
R101 VTAIL VTAIL.n11 2.72248
R102 VTAIL.n9 VTAIL.n7 2.32378
R103 VTAIL.n2 VTAIL.n1 2.32378
R104 VTAIL VTAIL.n1 0.985414
R105 B.n623 B.n622 585
R106 B.n623 B.n107 585
R107 B.n626 B.n625 585
R108 B.n627 B.n135 585
R109 B.n629 B.n628 585
R110 B.n631 B.n134 585
R111 B.n634 B.n633 585
R112 B.n635 B.n133 585
R113 B.n637 B.n636 585
R114 B.n639 B.n132 585
R115 B.n642 B.n641 585
R116 B.n643 B.n131 585
R117 B.n645 B.n644 585
R118 B.n647 B.n130 585
R119 B.n650 B.n649 585
R120 B.n651 B.n129 585
R121 B.n653 B.n652 585
R122 B.n655 B.n128 585
R123 B.n658 B.n657 585
R124 B.n659 B.n125 585
R125 B.n662 B.n661 585
R126 B.n664 B.n124 585
R127 B.n667 B.n666 585
R128 B.n668 B.n123 585
R129 B.n670 B.n669 585
R130 B.n672 B.n122 585
R131 B.n675 B.n674 585
R132 B.n676 B.n118 585
R133 B.n678 B.n677 585
R134 B.n680 B.n117 585
R135 B.n683 B.n682 585
R136 B.n684 B.n116 585
R137 B.n686 B.n685 585
R138 B.n688 B.n115 585
R139 B.n691 B.n690 585
R140 B.n692 B.n114 585
R141 B.n694 B.n693 585
R142 B.n696 B.n113 585
R143 B.n699 B.n698 585
R144 B.n700 B.n112 585
R145 B.n702 B.n701 585
R146 B.n704 B.n111 585
R147 B.n707 B.n706 585
R148 B.n708 B.n110 585
R149 B.n710 B.n709 585
R150 B.n712 B.n109 585
R151 B.n715 B.n714 585
R152 B.n716 B.n108 585
R153 B.n621 B.n106 585
R154 B.n719 B.n106 585
R155 B.n620 B.n105 585
R156 B.n720 B.n105 585
R157 B.n619 B.n104 585
R158 B.n721 B.n104 585
R159 B.n618 B.n617 585
R160 B.n617 B.n100 585
R161 B.n616 B.n99 585
R162 B.n727 B.n99 585
R163 B.n615 B.n98 585
R164 B.n728 B.n98 585
R165 B.n614 B.n97 585
R166 B.n729 B.n97 585
R167 B.n613 B.n612 585
R168 B.n612 B.n93 585
R169 B.n611 B.n92 585
R170 B.n735 B.n92 585
R171 B.n610 B.n91 585
R172 B.n736 B.n91 585
R173 B.n609 B.n90 585
R174 B.n737 B.n90 585
R175 B.n608 B.n607 585
R176 B.n607 B.n86 585
R177 B.n606 B.n85 585
R178 B.n743 B.n85 585
R179 B.n605 B.n84 585
R180 B.n744 B.n84 585
R181 B.n604 B.n83 585
R182 B.n745 B.n83 585
R183 B.n603 B.n602 585
R184 B.n602 B.n79 585
R185 B.n601 B.n78 585
R186 B.n751 B.n78 585
R187 B.n600 B.n77 585
R188 B.n752 B.n77 585
R189 B.n599 B.n76 585
R190 B.n753 B.n76 585
R191 B.n598 B.n597 585
R192 B.n597 B.n72 585
R193 B.n596 B.n71 585
R194 B.n759 B.n71 585
R195 B.n595 B.n70 585
R196 B.n760 B.n70 585
R197 B.n594 B.n69 585
R198 B.n761 B.n69 585
R199 B.n593 B.n592 585
R200 B.n592 B.n65 585
R201 B.n591 B.n64 585
R202 B.n767 B.n64 585
R203 B.n590 B.n63 585
R204 B.n768 B.n63 585
R205 B.n589 B.n62 585
R206 B.n769 B.n62 585
R207 B.n588 B.n587 585
R208 B.n587 B.n58 585
R209 B.n586 B.n57 585
R210 B.n775 B.n57 585
R211 B.n585 B.n56 585
R212 B.n776 B.n56 585
R213 B.n584 B.n55 585
R214 B.n777 B.n55 585
R215 B.n583 B.n582 585
R216 B.n582 B.n51 585
R217 B.n581 B.n50 585
R218 B.n783 B.n50 585
R219 B.n580 B.n49 585
R220 B.n784 B.n49 585
R221 B.n579 B.n48 585
R222 B.n785 B.n48 585
R223 B.n578 B.n577 585
R224 B.n577 B.n44 585
R225 B.n576 B.n43 585
R226 B.n791 B.n43 585
R227 B.n575 B.n42 585
R228 B.n792 B.n42 585
R229 B.n574 B.n41 585
R230 B.n793 B.n41 585
R231 B.n573 B.n572 585
R232 B.n572 B.n37 585
R233 B.n571 B.n36 585
R234 B.n799 B.n36 585
R235 B.n570 B.n35 585
R236 B.n800 B.n35 585
R237 B.n569 B.n34 585
R238 B.n801 B.n34 585
R239 B.n568 B.n567 585
R240 B.n567 B.n30 585
R241 B.n566 B.n29 585
R242 B.n807 B.n29 585
R243 B.n565 B.n28 585
R244 B.n808 B.n28 585
R245 B.n564 B.n27 585
R246 B.n809 B.n27 585
R247 B.n563 B.n562 585
R248 B.n562 B.n23 585
R249 B.n561 B.n22 585
R250 B.n815 B.n22 585
R251 B.n560 B.n21 585
R252 B.n816 B.n21 585
R253 B.n559 B.n20 585
R254 B.n817 B.n20 585
R255 B.n558 B.n557 585
R256 B.n557 B.n16 585
R257 B.n556 B.n15 585
R258 B.n823 B.n15 585
R259 B.n555 B.n14 585
R260 B.n824 B.n14 585
R261 B.n554 B.n13 585
R262 B.n825 B.n13 585
R263 B.n553 B.n552 585
R264 B.n552 B.n12 585
R265 B.n551 B.n550 585
R266 B.n551 B.n8 585
R267 B.n549 B.n7 585
R268 B.n832 B.n7 585
R269 B.n548 B.n6 585
R270 B.n833 B.n6 585
R271 B.n547 B.n5 585
R272 B.n834 B.n5 585
R273 B.n546 B.n545 585
R274 B.n545 B.n4 585
R275 B.n544 B.n136 585
R276 B.n544 B.n543 585
R277 B.n534 B.n137 585
R278 B.n138 B.n137 585
R279 B.n536 B.n535 585
R280 B.n537 B.n536 585
R281 B.n533 B.n143 585
R282 B.n143 B.n142 585
R283 B.n532 B.n531 585
R284 B.n531 B.n530 585
R285 B.n145 B.n144 585
R286 B.n146 B.n145 585
R287 B.n523 B.n522 585
R288 B.n524 B.n523 585
R289 B.n521 B.n151 585
R290 B.n151 B.n150 585
R291 B.n520 B.n519 585
R292 B.n519 B.n518 585
R293 B.n153 B.n152 585
R294 B.n154 B.n153 585
R295 B.n511 B.n510 585
R296 B.n512 B.n511 585
R297 B.n509 B.n159 585
R298 B.n159 B.n158 585
R299 B.n508 B.n507 585
R300 B.n507 B.n506 585
R301 B.n161 B.n160 585
R302 B.n162 B.n161 585
R303 B.n499 B.n498 585
R304 B.n500 B.n499 585
R305 B.n497 B.n167 585
R306 B.n167 B.n166 585
R307 B.n496 B.n495 585
R308 B.n495 B.n494 585
R309 B.n169 B.n168 585
R310 B.n170 B.n169 585
R311 B.n487 B.n486 585
R312 B.n488 B.n487 585
R313 B.n485 B.n174 585
R314 B.n178 B.n174 585
R315 B.n484 B.n483 585
R316 B.n483 B.n482 585
R317 B.n176 B.n175 585
R318 B.n177 B.n176 585
R319 B.n475 B.n474 585
R320 B.n476 B.n475 585
R321 B.n473 B.n183 585
R322 B.n183 B.n182 585
R323 B.n472 B.n471 585
R324 B.n471 B.n470 585
R325 B.n185 B.n184 585
R326 B.n186 B.n185 585
R327 B.n463 B.n462 585
R328 B.n464 B.n463 585
R329 B.n461 B.n191 585
R330 B.n191 B.n190 585
R331 B.n460 B.n459 585
R332 B.n459 B.n458 585
R333 B.n193 B.n192 585
R334 B.n194 B.n193 585
R335 B.n451 B.n450 585
R336 B.n452 B.n451 585
R337 B.n449 B.n198 585
R338 B.n202 B.n198 585
R339 B.n448 B.n447 585
R340 B.n447 B.n446 585
R341 B.n200 B.n199 585
R342 B.n201 B.n200 585
R343 B.n439 B.n438 585
R344 B.n440 B.n439 585
R345 B.n437 B.n207 585
R346 B.n207 B.n206 585
R347 B.n436 B.n435 585
R348 B.n435 B.n434 585
R349 B.n209 B.n208 585
R350 B.n210 B.n209 585
R351 B.n427 B.n426 585
R352 B.n428 B.n427 585
R353 B.n425 B.n215 585
R354 B.n215 B.n214 585
R355 B.n424 B.n423 585
R356 B.n423 B.n422 585
R357 B.n217 B.n216 585
R358 B.n218 B.n217 585
R359 B.n415 B.n414 585
R360 B.n416 B.n415 585
R361 B.n413 B.n223 585
R362 B.n223 B.n222 585
R363 B.n412 B.n411 585
R364 B.n411 B.n410 585
R365 B.n225 B.n224 585
R366 B.n226 B.n225 585
R367 B.n403 B.n402 585
R368 B.n404 B.n403 585
R369 B.n401 B.n230 585
R370 B.n234 B.n230 585
R371 B.n400 B.n399 585
R372 B.n399 B.n398 585
R373 B.n232 B.n231 585
R374 B.n233 B.n232 585
R375 B.n391 B.n390 585
R376 B.n392 B.n391 585
R377 B.n389 B.n239 585
R378 B.n239 B.n238 585
R379 B.n388 B.n387 585
R380 B.n387 B.n386 585
R381 B.n241 B.n240 585
R382 B.n242 B.n241 585
R383 B.n379 B.n378 585
R384 B.n380 B.n379 585
R385 B.n377 B.n247 585
R386 B.n247 B.n246 585
R387 B.n376 B.n375 585
R388 B.n375 B.n374 585
R389 B.n371 B.n251 585
R390 B.n370 B.n369 585
R391 B.n367 B.n252 585
R392 B.n367 B.n250 585
R393 B.n366 B.n365 585
R394 B.n364 B.n363 585
R395 B.n362 B.n254 585
R396 B.n360 B.n359 585
R397 B.n358 B.n255 585
R398 B.n357 B.n356 585
R399 B.n354 B.n256 585
R400 B.n352 B.n351 585
R401 B.n350 B.n257 585
R402 B.n349 B.n348 585
R403 B.n346 B.n258 585
R404 B.n344 B.n343 585
R405 B.n342 B.n259 585
R406 B.n341 B.n340 585
R407 B.n338 B.n260 585
R408 B.n336 B.n335 585
R409 B.n333 B.n261 585
R410 B.n332 B.n331 585
R411 B.n329 B.n264 585
R412 B.n327 B.n326 585
R413 B.n325 B.n265 585
R414 B.n324 B.n323 585
R415 B.n321 B.n266 585
R416 B.n319 B.n318 585
R417 B.n317 B.n267 585
R418 B.n315 B.n314 585
R419 B.n312 B.n270 585
R420 B.n310 B.n309 585
R421 B.n308 B.n271 585
R422 B.n307 B.n306 585
R423 B.n304 B.n272 585
R424 B.n302 B.n301 585
R425 B.n300 B.n273 585
R426 B.n299 B.n298 585
R427 B.n296 B.n274 585
R428 B.n294 B.n293 585
R429 B.n292 B.n275 585
R430 B.n291 B.n290 585
R431 B.n288 B.n276 585
R432 B.n286 B.n285 585
R433 B.n284 B.n277 585
R434 B.n283 B.n282 585
R435 B.n280 B.n278 585
R436 B.n249 B.n248 585
R437 B.n373 B.n372 585
R438 B.n374 B.n373 585
R439 B.n245 B.n244 585
R440 B.n246 B.n245 585
R441 B.n382 B.n381 585
R442 B.n381 B.n380 585
R443 B.n383 B.n243 585
R444 B.n243 B.n242 585
R445 B.n385 B.n384 585
R446 B.n386 B.n385 585
R447 B.n237 B.n236 585
R448 B.n238 B.n237 585
R449 B.n394 B.n393 585
R450 B.n393 B.n392 585
R451 B.n395 B.n235 585
R452 B.n235 B.n233 585
R453 B.n397 B.n396 585
R454 B.n398 B.n397 585
R455 B.n229 B.n228 585
R456 B.n234 B.n229 585
R457 B.n406 B.n405 585
R458 B.n405 B.n404 585
R459 B.n407 B.n227 585
R460 B.n227 B.n226 585
R461 B.n409 B.n408 585
R462 B.n410 B.n409 585
R463 B.n221 B.n220 585
R464 B.n222 B.n221 585
R465 B.n418 B.n417 585
R466 B.n417 B.n416 585
R467 B.n419 B.n219 585
R468 B.n219 B.n218 585
R469 B.n421 B.n420 585
R470 B.n422 B.n421 585
R471 B.n213 B.n212 585
R472 B.n214 B.n213 585
R473 B.n430 B.n429 585
R474 B.n429 B.n428 585
R475 B.n431 B.n211 585
R476 B.n211 B.n210 585
R477 B.n433 B.n432 585
R478 B.n434 B.n433 585
R479 B.n205 B.n204 585
R480 B.n206 B.n205 585
R481 B.n442 B.n441 585
R482 B.n441 B.n440 585
R483 B.n443 B.n203 585
R484 B.n203 B.n201 585
R485 B.n445 B.n444 585
R486 B.n446 B.n445 585
R487 B.n197 B.n196 585
R488 B.n202 B.n197 585
R489 B.n454 B.n453 585
R490 B.n453 B.n452 585
R491 B.n455 B.n195 585
R492 B.n195 B.n194 585
R493 B.n457 B.n456 585
R494 B.n458 B.n457 585
R495 B.n189 B.n188 585
R496 B.n190 B.n189 585
R497 B.n466 B.n465 585
R498 B.n465 B.n464 585
R499 B.n467 B.n187 585
R500 B.n187 B.n186 585
R501 B.n469 B.n468 585
R502 B.n470 B.n469 585
R503 B.n181 B.n180 585
R504 B.n182 B.n181 585
R505 B.n478 B.n477 585
R506 B.n477 B.n476 585
R507 B.n479 B.n179 585
R508 B.n179 B.n177 585
R509 B.n481 B.n480 585
R510 B.n482 B.n481 585
R511 B.n173 B.n172 585
R512 B.n178 B.n173 585
R513 B.n490 B.n489 585
R514 B.n489 B.n488 585
R515 B.n491 B.n171 585
R516 B.n171 B.n170 585
R517 B.n493 B.n492 585
R518 B.n494 B.n493 585
R519 B.n165 B.n164 585
R520 B.n166 B.n165 585
R521 B.n502 B.n501 585
R522 B.n501 B.n500 585
R523 B.n503 B.n163 585
R524 B.n163 B.n162 585
R525 B.n505 B.n504 585
R526 B.n506 B.n505 585
R527 B.n157 B.n156 585
R528 B.n158 B.n157 585
R529 B.n514 B.n513 585
R530 B.n513 B.n512 585
R531 B.n515 B.n155 585
R532 B.n155 B.n154 585
R533 B.n517 B.n516 585
R534 B.n518 B.n517 585
R535 B.n149 B.n148 585
R536 B.n150 B.n149 585
R537 B.n526 B.n525 585
R538 B.n525 B.n524 585
R539 B.n527 B.n147 585
R540 B.n147 B.n146 585
R541 B.n529 B.n528 585
R542 B.n530 B.n529 585
R543 B.n141 B.n140 585
R544 B.n142 B.n141 585
R545 B.n539 B.n538 585
R546 B.n538 B.n537 585
R547 B.n540 B.n139 585
R548 B.n139 B.n138 585
R549 B.n542 B.n541 585
R550 B.n543 B.n542 585
R551 B.n3 B.n0 585
R552 B.n4 B.n3 585
R553 B.n831 B.n1 585
R554 B.n832 B.n831 585
R555 B.n830 B.n829 585
R556 B.n830 B.n8 585
R557 B.n828 B.n9 585
R558 B.n12 B.n9 585
R559 B.n827 B.n826 585
R560 B.n826 B.n825 585
R561 B.n11 B.n10 585
R562 B.n824 B.n11 585
R563 B.n822 B.n821 585
R564 B.n823 B.n822 585
R565 B.n820 B.n17 585
R566 B.n17 B.n16 585
R567 B.n819 B.n818 585
R568 B.n818 B.n817 585
R569 B.n19 B.n18 585
R570 B.n816 B.n19 585
R571 B.n814 B.n813 585
R572 B.n815 B.n814 585
R573 B.n812 B.n24 585
R574 B.n24 B.n23 585
R575 B.n811 B.n810 585
R576 B.n810 B.n809 585
R577 B.n26 B.n25 585
R578 B.n808 B.n26 585
R579 B.n806 B.n805 585
R580 B.n807 B.n806 585
R581 B.n804 B.n31 585
R582 B.n31 B.n30 585
R583 B.n803 B.n802 585
R584 B.n802 B.n801 585
R585 B.n33 B.n32 585
R586 B.n800 B.n33 585
R587 B.n798 B.n797 585
R588 B.n799 B.n798 585
R589 B.n796 B.n38 585
R590 B.n38 B.n37 585
R591 B.n795 B.n794 585
R592 B.n794 B.n793 585
R593 B.n40 B.n39 585
R594 B.n792 B.n40 585
R595 B.n790 B.n789 585
R596 B.n791 B.n790 585
R597 B.n788 B.n45 585
R598 B.n45 B.n44 585
R599 B.n787 B.n786 585
R600 B.n786 B.n785 585
R601 B.n47 B.n46 585
R602 B.n784 B.n47 585
R603 B.n782 B.n781 585
R604 B.n783 B.n782 585
R605 B.n780 B.n52 585
R606 B.n52 B.n51 585
R607 B.n779 B.n778 585
R608 B.n778 B.n777 585
R609 B.n54 B.n53 585
R610 B.n776 B.n54 585
R611 B.n774 B.n773 585
R612 B.n775 B.n774 585
R613 B.n772 B.n59 585
R614 B.n59 B.n58 585
R615 B.n771 B.n770 585
R616 B.n770 B.n769 585
R617 B.n61 B.n60 585
R618 B.n768 B.n61 585
R619 B.n766 B.n765 585
R620 B.n767 B.n766 585
R621 B.n764 B.n66 585
R622 B.n66 B.n65 585
R623 B.n763 B.n762 585
R624 B.n762 B.n761 585
R625 B.n68 B.n67 585
R626 B.n760 B.n68 585
R627 B.n758 B.n757 585
R628 B.n759 B.n758 585
R629 B.n756 B.n73 585
R630 B.n73 B.n72 585
R631 B.n755 B.n754 585
R632 B.n754 B.n753 585
R633 B.n75 B.n74 585
R634 B.n752 B.n75 585
R635 B.n750 B.n749 585
R636 B.n751 B.n750 585
R637 B.n748 B.n80 585
R638 B.n80 B.n79 585
R639 B.n747 B.n746 585
R640 B.n746 B.n745 585
R641 B.n82 B.n81 585
R642 B.n744 B.n82 585
R643 B.n742 B.n741 585
R644 B.n743 B.n742 585
R645 B.n740 B.n87 585
R646 B.n87 B.n86 585
R647 B.n739 B.n738 585
R648 B.n738 B.n737 585
R649 B.n89 B.n88 585
R650 B.n736 B.n89 585
R651 B.n734 B.n733 585
R652 B.n735 B.n734 585
R653 B.n732 B.n94 585
R654 B.n94 B.n93 585
R655 B.n731 B.n730 585
R656 B.n730 B.n729 585
R657 B.n96 B.n95 585
R658 B.n728 B.n96 585
R659 B.n726 B.n725 585
R660 B.n727 B.n726 585
R661 B.n724 B.n101 585
R662 B.n101 B.n100 585
R663 B.n723 B.n722 585
R664 B.n722 B.n721 585
R665 B.n103 B.n102 585
R666 B.n720 B.n103 585
R667 B.n718 B.n717 585
R668 B.n719 B.n718 585
R669 B.n835 B.n834 585
R670 B.n833 B.n2 585
R671 B.n718 B.n108 559.769
R672 B.n623 B.n106 559.769
R673 B.n375 B.n249 559.769
R674 B.n373 B.n251 559.769
R675 B.n624 B.n107 256.663
R676 B.n630 B.n107 256.663
R677 B.n632 B.n107 256.663
R678 B.n638 B.n107 256.663
R679 B.n640 B.n107 256.663
R680 B.n646 B.n107 256.663
R681 B.n648 B.n107 256.663
R682 B.n654 B.n107 256.663
R683 B.n656 B.n107 256.663
R684 B.n663 B.n107 256.663
R685 B.n665 B.n107 256.663
R686 B.n671 B.n107 256.663
R687 B.n673 B.n107 256.663
R688 B.n679 B.n107 256.663
R689 B.n681 B.n107 256.663
R690 B.n687 B.n107 256.663
R691 B.n689 B.n107 256.663
R692 B.n695 B.n107 256.663
R693 B.n697 B.n107 256.663
R694 B.n703 B.n107 256.663
R695 B.n705 B.n107 256.663
R696 B.n711 B.n107 256.663
R697 B.n713 B.n107 256.663
R698 B.n368 B.n250 256.663
R699 B.n253 B.n250 256.663
R700 B.n361 B.n250 256.663
R701 B.n355 B.n250 256.663
R702 B.n353 B.n250 256.663
R703 B.n347 B.n250 256.663
R704 B.n345 B.n250 256.663
R705 B.n339 B.n250 256.663
R706 B.n337 B.n250 256.663
R707 B.n330 B.n250 256.663
R708 B.n328 B.n250 256.663
R709 B.n322 B.n250 256.663
R710 B.n320 B.n250 256.663
R711 B.n313 B.n250 256.663
R712 B.n311 B.n250 256.663
R713 B.n305 B.n250 256.663
R714 B.n303 B.n250 256.663
R715 B.n297 B.n250 256.663
R716 B.n295 B.n250 256.663
R717 B.n289 B.n250 256.663
R718 B.n287 B.n250 256.663
R719 B.n281 B.n250 256.663
R720 B.n279 B.n250 256.663
R721 B.n837 B.n836 256.663
R722 B.n119 B.t6 235.392
R723 B.n126 B.t17 235.392
R724 B.n268 B.t14 235.392
R725 B.n262 B.t10 235.392
R726 B.n714 B.n712 163.367
R727 B.n710 B.n110 163.367
R728 B.n706 B.n704 163.367
R729 B.n702 B.n112 163.367
R730 B.n698 B.n696 163.367
R731 B.n694 B.n114 163.367
R732 B.n690 B.n688 163.367
R733 B.n686 B.n116 163.367
R734 B.n682 B.n680 163.367
R735 B.n678 B.n118 163.367
R736 B.n674 B.n672 163.367
R737 B.n670 B.n123 163.367
R738 B.n666 B.n664 163.367
R739 B.n662 B.n125 163.367
R740 B.n657 B.n655 163.367
R741 B.n653 B.n129 163.367
R742 B.n649 B.n647 163.367
R743 B.n645 B.n131 163.367
R744 B.n641 B.n639 163.367
R745 B.n637 B.n133 163.367
R746 B.n633 B.n631 163.367
R747 B.n629 B.n135 163.367
R748 B.n625 B.n623 163.367
R749 B.n375 B.n247 163.367
R750 B.n379 B.n247 163.367
R751 B.n379 B.n241 163.367
R752 B.n387 B.n241 163.367
R753 B.n387 B.n239 163.367
R754 B.n391 B.n239 163.367
R755 B.n391 B.n232 163.367
R756 B.n399 B.n232 163.367
R757 B.n399 B.n230 163.367
R758 B.n403 B.n230 163.367
R759 B.n403 B.n225 163.367
R760 B.n411 B.n225 163.367
R761 B.n411 B.n223 163.367
R762 B.n415 B.n223 163.367
R763 B.n415 B.n217 163.367
R764 B.n423 B.n217 163.367
R765 B.n423 B.n215 163.367
R766 B.n427 B.n215 163.367
R767 B.n427 B.n209 163.367
R768 B.n435 B.n209 163.367
R769 B.n435 B.n207 163.367
R770 B.n439 B.n207 163.367
R771 B.n439 B.n200 163.367
R772 B.n447 B.n200 163.367
R773 B.n447 B.n198 163.367
R774 B.n451 B.n198 163.367
R775 B.n451 B.n193 163.367
R776 B.n459 B.n193 163.367
R777 B.n459 B.n191 163.367
R778 B.n463 B.n191 163.367
R779 B.n463 B.n185 163.367
R780 B.n471 B.n185 163.367
R781 B.n471 B.n183 163.367
R782 B.n475 B.n183 163.367
R783 B.n475 B.n176 163.367
R784 B.n483 B.n176 163.367
R785 B.n483 B.n174 163.367
R786 B.n487 B.n174 163.367
R787 B.n487 B.n169 163.367
R788 B.n495 B.n169 163.367
R789 B.n495 B.n167 163.367
R790 B.n499 B.n167 163.367
R791 B.n499 B.n161 163.367
R792 B.n507 B.n161 163.367
R793 B.n507 B.n159 163.367
R794 B.n511 B.n159 163.367
R795 B.n511 B.n153 163.367
R796 B.n519 B.n153 163.367
R797 B.n519 B.n151 163.367
R798 B.n523 B.n151 163.367
R799 B.n523 B.n145 163.367
R800 B.n531 B.n145 163.367
R801 B.n531 B.n143 163.367
R802 B.n536 B.n143 163.367
R803 B.n536 B.n137 163.367
R804 B.n544 B.n137 163.367
R805 B.n545 B.n544 163.367
R806 B.n545 B.n5 163.367
R807 B.n6 B.n5 163.367
R808 B.n7 B.n6 163.367
R809 B.n551 B.n7 163.367
R810 B.n552 B.n551 163.367
R811 B.n552 B.n13 163.367
R812 B.n14 B.n13 163.367
R813 B.n15 B.n14 163.367
R814 B.n557 B.n15 163.367
R815 B.n557 B.n20 163.367
R816 B.n21 B.n20 163.367
R817 B.n22 B.n21 163.367
R818 B.n562 B.n22 163.367
R819 B.n562 B.n27 163.367
R820 B.n28 B.n27 163.367
R821 B.n29 B.n28 163.367
R822 B.n567 B.n29 163.367
R823 B.n567 B.n34 163.367
R824 B.n35 B.n34 163.367
R825 B.n36 B.n35 163.367
R826 B.n572 B.n36 163.367
R827 B.n572 B.n41 163.367
R828 B.n42 B.n41 163.367
R829 B.n43 B.n42 163.367
R830 B.n577 B.n43 163.367
R831 B.n577 B.n48 163.367
R832 B.n49 B.n48 163.367
R833 B.n50 B.n49 163.367
R834 B.n582 B.n50 163.367
R835 B.n582 B.n55 163.367
R836 B.n56 B.n55 163.367
R837 B.n57 B.n56 163.367
R838 B.n587 B.n57 163.367
R839 B.n587 B.n62 163.367
R840 B.n63 B.n62 163.367
R841 B.n64 B.n63 163.367
R842 B.n592 B.n64 163.367
R843 B.n592 B.n69 163.367
R844 B.n70 B.n69 163.367
R845 B.n71 B.n70 163.367
R846 B.n597 B.n71 163.367
R847 B.n597 B.n76 163.367
R848 B.n77 B.n76 163.367
R849 B.n78 B.n77 163.367
R850 B.n602 B.n78 163.367
R851 B.n602 B.n83 163.367
R852 B.n84 B.n83 163.367
R853 B.n85 B.n84 163.367
R854 B.n607 B.n85 163.367
R855 B.n607 B.n90 163.367
R856 B.n91 B.n90 163.367
R857 B.n92 B.n91 163.367
R858 B.n612 B.n92 163.367
R859 B.n612 B.n97 163.367
R860 B.n98 B.n97 163.367
R861 B.n99 B.n98 163.367
R862 B.n617 B.n99 163.367
R863 B.n617 B.n104 163.367
R864 B.n105 B.n104 163.367
R865 B.n106 B.n105 163.367
R866 B.n369 B.n367 163.367
R867 B.n367 B.n366 163.367
R868 B.n363 B.n362 163.367
R869 B.n360 B.n255 163.367
R870 B.n356 B.n354 163.367
R871 B.n352 B.n257 163.367
R872 B.n348 B.n346 163.367
R873 B.n344 B.n259 163.367
R874 B.n340 B.n338 163.367
R875 B.n336 B.n261 163.367
R876 B.n331 B.n329 163.367
R877 B.n327 B.n265 163.367
R878 B.n323 B.n321 163.367
R879 B.n319 B.n267 163.367
R880 B.n314 B.n312 163.367
R881 B.n310 B.n271 163.367
R882 B.n306 B.n304 163.367
R883 B.n302 B.n273 163.367
R884 B.n298 B.n296 163.367
R885 B.n294 B.n275 163.367
R886 B.n290 B.n288 163.367
R887 B.n286 B.n277 163.367
R888 B.n282 B.n280 163.367
R889 B.n373 B.n245 163.367
R890 B.n381 B.n245 163.367
R891 B.n381 B.n243 163.367
R892 B.n385 B.n243 163.367
R893 B.n385 B.n237 163.367
R894 B.n393 B.n237 163.367
R895 B.n393 B.n235 163.367
R896 B.n397 B.n235 163.367
R897 B.n397 B.n229 163.367
R898 B.n405 B.n229 163.367
R899 B.n405 B.n227 163.367
R900 B.n409 B.n227 163.367
R901 B.n409 B.n221 163.367
R902 B.n417 B.n221 163.367
R903 B.n417 B.n219 163.367
R904 B.n421 B.n219 163.367
R905 B.n421 B.n213 163.367
R906 B.n429 B.n213 163.367
R907 B.n429 B.n211 163.367
R908 B.n433 B.n211 163.367
R909 B.n433 B.n205 163.367
R910 B.n441 B.n205 163.367
R911 B.n441 B.n203 163.367
R912 B.n445 B.n203 163.367
R913 B.n445 B.n197 163.367
R914 B.n453 B.n197 163.367
R915 B.n453 B.n195 163.367
R916 B.n457 B.n195 163.367
R917 B.n457 B.n189 163.367
R918 B.n465 B.n189 163.367
R919 B.n465 B.n187 163.367
R920 B.n469 B.n187 163.367
R921 B.n469 B.n181 163.367
R922 B.n477 B.n181 163.367
R923 B.n477 B.n179 163.367
R924 B.n481 B.n179 163.367
R925 B.n481 B.n173 163.367
R926 B.n489 B.n173 163.367
R927 B.n489 B.n171 163.367
R928 B.n493 B.n171 163.367
R929 B.n493 B.n165 163.367
R930 B.n501 B.n165 163.367
R931 B.n501 B.n163 163.367
R932 B.n505 B.n163 163.367
R933 B.n505 B.n157 163.367
R934 B.n513 B.n157 163.367
R935 B.n513 B.n155 163.367
R936 B.n517 B.n155 163.367
R937 B.n517 B.n149 163.367
R938 B.n525 B.n149 163.367
R939 B.n525 B.n147 163.367
R940 B.n529 B.n147 163.367
R941 B.n529 B.n141 163.367
R942 B.n538 B.n141 163.367
R943 B.n538 B.n139 163.367
R944 B.n542 B.n139 163.367
R945 B.n542 B.n3 163.367
R946 B.n835 B.n3 163.367
R947 B.n831 B.n2 163.367
R948 B.n831 B.n830 163.367
R949 B.n830 B.n9 163.367
R950 B.n826 B.n9 163.367
R951 B.n826 B.n11 163.367
R952 B.n822 B.n11 163.367
R953 B.n822 B.n17 163.367
R954 B.n818 B.n17 163.367
R955 B.n818 B.n19 163.367
R956 B.n814 B.n19 163.367
R957 B.n814 B.n24 163.367
R958 B.n810 B.n24 163.367
R959 B.n810 B.n26 163.367
R960 B.n806 B.n26 163.367
R961 B.n806 B.n31 163.367
R962 B.n802 B.n31 163.367
R963 B.n802 B.n33 163.367
R964 B.n798 B.n33 163.367
R965 B.n798 B.n38 163.367
R966 B.n794 B.n38 163.367
R967 B.n794 B.n40 163.367
R968 B.n790 B.n40 163.367
R969 B.n790 B.n45 163.367
R970 B.n786 B.n45 163.367
R971 B.n786 B.n47 163.367
R972 B.n782 B.n47 163.367
R973 B.n782 B.n52 163.367
R974 B.n778 B.n52 163.367
R975 B.n778 B.n54 163.367
R976 B.n774 B.n54 163.367
R977 B.n774 B.n59 163.367
R978 B.n770 B.n59 163.367
R979 B.n770 B.n61 163.367
R980 B.n766 B.n61 163.367
R981 B.n766 B.n66 163.367
R982 B.n762 B.n66 163.367
R983 B.n762 B.n68 163.367
R984 B.n758 B.n68 163.367
R985 B.n758 B.n73 163.367
R986 B.n754 B.n73 163.367
R987 B.n754 B.n75 163.367
R988 B.n750 B.n75 163.367
R989 B.n750 B.n80 163.367
R990 B.n746 B.n80 163.367
R991 B.n746 B.n82 163.367
R992 B.n742 B.n82 163.367
R993 B.n742 B.n87 163.367
R994 B.n738 B.n87 163.367
R995 B.n738 B.n89 163.367
R996 B.n734 B.n89 163.367
R997 B.n734 B.n94 163.367
R998 B.n730 B.n94 163.367
R999 B.n730 B.n96 163.367
R1000 B.n726 B.n96 163.367
R1001 B.n726 B.n101 163.367
R1002 B.n722 B.n101 163.367
R1003 B.n722 B.n103 163.367
R1004 B.n718 B.n103 163.367
R1005 B.n126 B.t18 158.131
R1006 B.n268 B.t16 158.131
R1007 B.n119 B.t8 158.126
R1008 B.n262 B.t13 158.126
R1009 B.n374 B.n250 157.885
R1010 B.n719 B.n107 157.885
R1011 B.n120 B.n119 83.3944
R1012 B.n127 B.n126 83.3944
R1013 B.n269 B.n268 83.3944
R1014 B.n263 B.n262 83.3944
R1015 B.n374 B.n246 78.3661
R1016 B.n380 B.n246 78.3661
R1017 B.n380 B.n242 78.3661
R1018 B.n386 B.n242 78.3661
R1019 B.n386 B.n238 78.3661
R1020 B.n392 B.n238 78.3661
R1021 B.n392 B.n233 78.3661
R1022 B.n398 B.n233 78.3661
R1023 B.n398 B.n234 78.3661
R1024 B.n404 B.n226 78.3661
R1025 B.n410 B.n226 78.3661
R1026 B.n410 B.n222 78.3661
R1027 B.n416 B.n222 78.3661
R1028 B.n416 B.n218 78.3661
R1029 B.n422 B.n218 78.3661
R1030 B.n422 B.n214 78.3661
R1031 B.n428 B.n214 78.3661
R1032 B.n428 B.n210 78.3661
R1033 B.n434 B.n210 78.3661
R1034 B.n434 B.n206 78.3661
R1035 B.n440 B.n206 78.3661
R1036 B.n440 B.n201 78.3661
R1037 B.n446 B.n201 78.3661
R1038 B.n446 B.n202 78.3661
R1039 B.n452 B.n194 78.3661
R1040 B.n458 B.n194 78.3661
R1041 B.n458 B.n190 78.3661
R1042 B.n464 B.n190 78.3661
R1043 B.n464 B.n186 78.3661
R1044 B.n470 B.n186 78.3661
R1045 B.n470 B.n182 78.3661
R1046 B.n476 B.n182 78.3661
R1047 B.n476 B.n177 78.3661
R1048 B.n482 B.n177 78.3661
R1049 B.n482 B.n178 78.3661
R1050 B.n488 B.n170 78.3661
R1051 B.n494 B.n170 78.3661
R1052 B.n494 B.n166 78.3661
R1053 B.n500 B.n166 78.3661
R1054 B.n500 B.n162 78.3661
R1055 B.n506 B.n162 78.3661
R1056 B.n506 B.n158 78.3661
R1057 B.n512 B.n158 78.3661
R1058 B.n512 B.n154 78.3661
R1059 B.n518 B.n154 78.3661
R1060 B.n518 B.n150 78.3661
R1061 B.n524 B.n150 78.3661
R1062 B.n530 B.n146 78.3661
R1063 B.n530 B.n142 78.3661
R1064 B.n537 B.n142 78.3661
R1065 B.n537 B.n138 78.3661
R1066 B.n543 B.n138 78.3661
R1067 B.n543 B.n4 78.3661
R1068 B.n834 B.n4 78.3661
R1069 B.n834 B.n833 78.3661
R1070 B.n833 B.n832 78.3661
R1071 B.n832 B.n8 78.3661
R1072 B.n12 B.n8 78.3661
R1073 B.n825 B.n12 78.3661
R1074 B.n825 B.n824 78.3661
R1075 B.n824 B.n823 78.3661
R1076 B.n823 B.n16 78.3661
R1077 B.n817 B.n816 78.3661
R1078 B.n816 B.n815 78.3661
R1079 B.n815 B.n23 78.3661
R1080 B.n809 B.n23 78.3661
R1081 B.n809 B.n808 78.3661
R1082 B.n808 B.n807 78.3661
R1083 B.n807 B.n30 78.3661
R1084 B.n801 B.n30 78.3661
R1085 B.n801 B.n800 78.3661
R1086 B.n800 B.n799 78.3661
R1087 B.n799 B.n37 78.3661
R1088 B.n793 B.n37 78.3661
R1089 B.n792 B.n791 78.3661
R1090 B.n791 B.n44 78.3661
R1091 B.n785 B.n44 78.3661
R1092 B.n785 B.n784 78.3661
R1093 B.n784 B.n783 78.3661
R1094 B.n783 B.n51 78.3661
R1095 B.n777 B.n51 78.3661
R1096 B.n777 B.n776 78.3661
R1097 B.n776 B.n775 78.3661
R1098 B.n775 B.n58 78.3661
R1099 B.n769 B.n58 78.3661
R1100 B.n768 B.n767 78.3661
R1101 B.n767 B.n65 78.3661
R1102 B.n761 B.n65 78.3661
R1103 B.n761 B.n760 78.3661
R1104 B.n760 B.n759 78.3661
R1105 B.n759 B.n72 78.3661
R1106 B.n753 B.n72 78.3661
R1107 B.n753 B.n752 78.3661
R1108 B.n752 B.n751 78.3661
R1109 B.n751 B.n79 78.3661
R1110 B.n745 B.n79 78.3661
R1111 B.n745 B.n744 78.3661
R1112 B.n744 B.n743 78.3661
R1113 B.n743 B.n86 78.3661
R1114 B.n737 B.n86 78.3661
R1115 B.n736 B.n735 78.3661
R1116 B.n735 B.n93 78.3661
R1117 B.n729 B.n93 78.3661
R1118 B.n729 B.n728 78.3661
R1119 B.n728 B.n727 78.3661
R1120 B.n727 B.n100 78.3661
R1121 B.n721 B.n100 78.3661
R1122 B.n721 B.n720 78.3661
R1123 B.n720 B.n719 78.3661
R1124 B.n127 B.t19 74.7364
R1125 B.n269 B.t15 74.7364
R1126 B.n120 B.t9 74.7325
R1127 B.n263 B.t12 74.7325
R1128 B.n178 B.t5 72.604
R1129 B.t1 B.n792 72.604
R1130 B.n713 B.n108 71.676
R1131 B.n712 B.n711 71.676
R1132 B.n705 B.n110 71.676
R1133 B.n704 B.n703 71.676
R1134 B.n697 B.n112 71.676
R1135 B.n696 B.n695 71.676
R1136 B.n689 B.n114 71.676
R1137 B.n688 B.n687 71.676
R1138 B.n681 B.n116 71.676
R1139 B.n680 B.n679 71.676
R1140 B.n673 B.n118 71.676
R1141 B.n672 B.n671 71.676
R1142 B.n665 B.n123 71.676
R1143 B.n664 B.n663 71.676
R1144 B.n656 B.n125 71.676
R1145 B.n655 B.n654 71.676
R1146 B.n648 B.n129 71.676
R1147 B.n647 B.n646 71.676
R1148 B.n640 B.n131 71.676
R1149 B.n639 B.n638 71.676
R1150 B.n632 B.n133 71.676
R1151 B.n631 B.n630 71.676
R1152 B.n624 B.n135 71.676
R1153 B.n625 B.n624 71.676
R1154 B.n630 B.n629 71.676
R1155 B.n633 B.n632 71.676
R1156 B.n638 B.n637 71.676
R1157 B.n641 B.n640 71.676
R1158 B.n646 B.n645 71.676
R1159 B.n649 B.n648 71.676
R1160 B.n654 B.n653 71.676
R1161 B.n657 B.n656 71.676
R1162 B.n663 B.n662 71.676
R1163 B.n666 B.n665 71.676
R1164 B.n671 B.n670 71.676
R1165 B.n674 B.n673 71.676
R1166 B.n679 B.n678 71.676
R1167 B.n682 B.n681 71.676
R1168 B.n687 B.n686 71.676
R1169 B.n690 B.n689 71.676
R1170 B.n695 B.n694 71.676
R1171 B.n698 B.n697 71.676
R1172 B.n703 B.n702 71.676
R1173 B.n706 B.n705 71.676
R1174 B.n711 B.n710 71.676
R1175 B.n714 B.n713 71.676
R1176 B.n368 B.n251 71.676
R1177 B.n366 B.n253 71.676
R1178 B.n362 B.n361 71.676
R1179 B.n355 B.n255 71.676
R1180 B.n354 B.n353 71.676
R1181 B.n347 B.n257 71.676
R1182 B.n346 B.n345 71.676
R1183 B.n339 B.n259 71.676
R1184 B.n338 B.n337 71.676
R1185 B.n330 B.n261 71.676
R1186 B.n329 B.n328 71.676
R1187 B.n322 B.n265 71.676
R1188 B.n321 B.n320 71.676
R1189 B.n313 B.n267 71.676
R1190 B.n312 B.n311 71.676
R1191 B.n305 B.n271 71.676
R1192 B.n304 B.n303 71.676
R1193 B.n297 B.n273 71.676
R1194 B.n296 B.n295 71.676
R1195 B.n289 B.n275 71.676
R1196 B.n288 B.n287 71.676
R1197 B.n281 B.n277 71.676
R1198 B.n280 B.n279 71.676
R1199 B.n369 B.n368 71.676
R1200 B.n363 B.n253 71.676
R1201 B.n361 B.n360 71.676
R1202 B.n356 B.n355 71.676
R1203 B.n353 B.n352 71.676
R1204 B.n348 B.n347 71.676
R1205 B.n345 B.n344 71.676
R1206 B.n340 B.n339 71.676
R1207 B.n337 B.n336 71.676
R1208 B.n331 B.n330 71.676
R1209 B.n328 B.n327 71.676
R1210 B.n323 B.n322 71.676
R1211 B.n320 B.n319 71.676
R1212 B.n314 B.n313 71.676
R1213 B.n311 B.n310 71.676
R1214 B.n306 B.n305 71.676
R1215 B.n303 B.n302 71.676
R1216 B.n298 B.n297 71.676
R1217 B.n295 B.n294 71.676
R1218 B.n290 B.n289 71.676
R1219 B.n287 B.n286 71.676
R1220 B.n282 B.n281 71.676
R1221 B.n279 B.n249 71.676
R1222 B.n836 B.n835 71.676
R1223 B.n836 B.n2 71.676
R1224 B.n121 B.n120 59.5399
R1225 B.n660 B.n127 59.5399
R1226 B.n316 B.n269 59.5399
R1227 B.n334 B.n263 59.5399
R1228 B.n452 B.t3 56.4699
R1229 B.n769 B.t4 56.4699
R1230 B.n404 B.t11 44.9455
R1231 B.n524 B.t0 44.9455
R1232 B.n817 B.t2 44.9455
R1233 B.n737 B.t7 44.9455
R1234 B.n372 B.n371 36.3712
R1235 B.n376 B.n248 36.3712
R1236 B.n622 B.n621 36.3712
R1237 B.n717 B.n716 36.3712
R1238 B.n234 B.t11 33.4211
R1239 B.t0 B.n146 33.4211
R1240 B.t2 B.n16 33.4211
R1241 B.t7 B.n736 33.4211
R1242 B.n202 B.t3 21.8968
R1243 B.t4 B.n768 21.8968
R1244 B B.n837 18.0485
R1245 B.n372 B.n244 10.6151
R1246 B.n382 B.n244 10.6151
R1247 B.n383 B.n382 10.6151
R1248 B.n384 B.n383 10.6151
R1249 B.n384 B.n236 10.6151
R1250 B.n394 B.n236 10.6151
R1251 B.n395 B.n394 10.6151
R1252 B.n396 B.n395 10.6151
R1253 B.n396 B.n228 10.6151
R1254 B.n406 B.n228 10.6151
R1255 B.n407 B.n406 10.6151
R1256 B.n408 B.n407 10.6151
R1257 B.n408 B.n220 10.6151
R1258 B.n418 B.n220 10.6151
R1259 B.n419 B.n418 10.6151
R1260 B.n420 B.n419 10.6151
R1261 B.n420 B.n212 10.6151
R1262 B.n430 B.n212 10.6151
R1263 B.n431 B.n430 10.6151
R1264 B.n432 B.n431 10.6151
R1265 B.n432 B.n204 10.6151
R1266 B.n442 B.n204 10.6151
R1267 B.n443 B.n442 10.6151
R1268 B.n444 B.n443 10.6151
R1269 B.n444 B.n196 10.6151
R1270 B.n454 B.n196 10.6151
R1271 B.n455 B.n454 10.6151
R1272 B.n456 B.n455 10.6151
R1273 B.n456 B.n188 10.6151
R1274 B.n466 B.n188 10.6151
R1275 B.n467 B.n466 10.6151
R1276 B.n468 B.n467 10.6151
R1277 B.n468 B.n180 10.6151
R1278 B.n478 B.n180 10.6151
R1279 B.n479 B.n478 10.6151
R1280 B.n480 B.n479 10.6151
R1281 B.n480 B.n172 10.6151
R1282 B.n490 B.n172 10.6151
R1283 B.n491 B.n490 10.6151
R1284 B.n492 B.n491 10.6151
R1285 B.n492 B.n164 10.6151
R1286 B.n502 B.n164 10.6151
R1287 B.n503 B.n502 10.6151
R1288 B.n504 B.n503 10.6151
R1289 B.n504 B.n156 10.6151
R1290 B.n514 B.n156 10.6151
R1291 B.n515 B.n514 10.6151
R1292 B.n516 B.n515 10.6151
R1293 B.n516 B.n148 10.6151
R1294 B.n526 B.n148 10.6151
R1295 B.n527 B.n526 10.6151
R1296 B.n528 B.n527 10.6151
R1297 B.n528 B.n140 10.6151
R1298 B.n539 B.n140 10.6151
R1299 B.n540 B.n539 10.6151
R1300 B.n541 B.n540 10.6151
R1301 B.n541 B.n0 10.6151
R1302 B.n371 B.n370 10.6151
R1303 B.n370 B.n252 10.6151
R1304 B.n365 B.n252 10.6151
R1305 B.n365 B.n364 10.6151
R1306 B.n364 B.n254 10.6151
R1307 B.n359 B.n254 10.6151
R1308 B.n359 B.n358 10.6151
R1309 B.n358 B.n357 10.6151
R1310 B.n357 B.n256 10.6151
R1311 B.n351 B.n256 10.6151
R1312 B.n351 B.n350 10.6151
R1313 B.n350 B.n349 10.6151
R1314 B.n349 B.n258 10.6151
R1315 B.n343 B.n258 10.6151
R1316 B.n343 B.n342 10.6151
R1317 B.n342 B.n341 10.6151
R1318 B.n341 B.n260 10.6151
R1319 B.n335 B.n260 10.6151
R1320 B.n333 B.n332 10.6151
R1321 B.n332 B.n264 10.6151
R1322 B.n326 B.n264 10.6151
R1323 B.n326 B.n325 10.6151
R1324 B.n325 B.n324 10.6151
R1325 B.n324 B.n266 10.6151
R1326 B.n318 B.n266 10.6151
R1327 B.n318 B.n317 10.6151
R1328 B.n315 B.n270 10.6151
R1329 B.n309 B.n270 10.6151
R1330 B.n309 B.n308 10.6151
R1331 B.n308 B.n307 10.6151
R1332 B.n307 B.n272 10.6151
R1333 B.n301 B.n272 10.6151
R1334 B.n301 B.n300 10.6151
R1335 B.n300 B.n299 10.6151
R1336 B.n299 B.n274 10.6151
R1337 B.n293 B.n274 10.6151
R1338 B.n293 B.n292 10.6151
R1339 B.n292 B.n291 10.6151
R1340 B.n291 B.n276 10.6151
R1341 B.n285 B.n276 10.6151
R1342 B.n285 B.n284 10.6151
R1343 B.n284 B.n283 10.6151
R1344 B.n283 B.n278 10.6151
R1345 B.n278 B.n248 10.6151
R1346 B.n377 B.n376 10.6151
R1347 B.n378 B.n377 10.6151
R1348 B.n378 B.n240 10.6151
R1349 B.n388 B.n240 10.6151
R1350 B.n389 B.n388 10.6151
R1351 B.n390 B.n389 10.6151
R1352 B.n390 B.n231 10.6151
R1353 B.n400 B.n231 10.6151
R1354 B.n401 B.n400 10.6151
R1355 B.n402 B.n401 10.6151
R1356 B.n402 B.n224 10.6151
R1357 B.n412 B.n224 10.6151
R1358 B.n413 B.n412 10.6151
R1359 B.n414 B.n413 10.6151
R1360 B.n414 B.n216 10.6151
R1361 B.n424 B.n216 10.6151
R1362 B.n425 B.n424 10.6151
R1363 B.n426 B.n425 10.6151
R1364 B.n426 B.n208 10.6151
R1365 B.n436 B.n208 10.6151
R1366 B.n437 B.n436 10.6151
R1367 B.n438 B.n437 10.6151
R1368 B.n438 B.n199 10.6151
R1369 B.n448 B.n199 10.6151
R1370 B.n449 B.n448 10.6151
R1371 B.n450 B.n449 10.6151
R1372 B.n450 B.n192 10.6151
R1373 B.n460 B.n192 10.6151
R1374 B.n461 B.n460 10.6151
R1375 B.n462 B.n461 10.6151
R1376 B.n462 B.n184 10.6151
R1377 B.n472 B.n184 10.6151
R1378 B.n473 B.n472 10.6151
R1379 B.n474 B.n473 10.6151
R1380 B.n474 B.n175 10.6151
R1381 B.n484 B.n175 10.6151
R1382 B.n485 B.n484 10.6151
R1383 B.n486 B.n485 10.6151
R1384 B.n486 B.n168 10.6151
R1385 B.n496 B.n168 10.6151
R1386 B.n497 B.n496 10.6151
R1387 B.n498 B.n497 10.6151
R1388 B.n498 B.n160 10.6151
R1389 B.n508 B.n160 10.6151
R1390 B.n509 B.n508 10.6151
R1391 B.n510 B.n509 10.6151
R1392 B.n510 B.n152 10.6151
R1393 B.n520 B.n152 10.6151
R1394 B.n521 B.n520 10.6151
R1395 B.n522 B.n521 10.6151
R1396 B.n522 B.n144 10.6151
R1397 B.n532 B.n144 10.6151
R1398 B.n533 B.n532 10.6151
R1399 B.n535 B.n533 10.6151
R1400 B.n535 B.n534 10.6151
R1401 B.n534 B.n136 10.6151
R1402 B.n546 B.n136 10.6151
R1403 B.n547 B.n546 10.6151
R1404 B.n548 B.n547 10.6151
R1405 B.n549 B.n548 10.6151
R1406 B.n550 B.n549 10.6151
R1407 B.n553 B.n550 10.6151
R1408 B.n554 B.n553 10.6151
R1409 B.n555 B.n554 10.6151
R1410 B.n556 B.n555 10.6151
R1411 B.n558 B.n556 10.6151
R1412 B.n559 B.n558 10.6151
R1413 B.n560 B.n559 10.6151
R1414 B.n561 B.n560 10.6151
R1415 B.n563 B.n561 10.6151
R1416 B.n564 B.n563 10.6151
R1417 B.n565 B.n564 10.6151
R1418 B.n566 B.n565 10.6151
R1419 B.n568 B.n566 10.6151
R1420 B.n569 B.n568 10.6151
R1421 B.n570 B.n569 10.6151
R1422 B.n571 B.n570 10.6151
R1423 B.n573 B.n571 10.6151
R1424 B.n574 B.n573 10.6151
R1425 B.n575 B.n574 10.6151
R1426 B.n576 B.n575 10.6151
R1427 B.n578 B.n576 10.6151
R1428 B.n579 B.n578 10.6151
R1429 B.n580 B.n579 10.6151
R1430 B.n581 B.n580 10.6151
R1431 B.n583 B.n581 10.6151
R1432 B.n584 B.n583 10.6151
R1433 B.n585 B.n584 10.6151
R1434 B.n586 B.n585 10.6151
R1435 B.n588 B.n586 10.6151
R1436 B.n589 B.n588 10.6151
R1437 B.n590 B.n589 10.6151
R1438 B.n591 B.n590 10.6151
R1439 B.n593 B.n591 10.6151
R1440 B.n594 B.n593 10.6151
R1441 B.n595 B.n594 10.6151
R1442 B.n596 B.n595 10.6151
R1443 B.n598 B.n596 10.6151
R1444 B.n599 B.n598 10.6151
R1445 B.n600 B.n599 10.6151
R1446 B.n601 B.n600 10.6151
R1447 B.n603 B.n601 10.6151
R1448 B.n604 B.n603 10.6151
R1449 B.n605 B.n604 10.6151
R1450 B.n606 B.n605 10.6151
R1451 B.n608 B.n606 10.6151
R1452 B.n609 B.n608 10.6151
R1453 B.n610 B.n609 10.6151
R1454 B.n611 B.n610 10.6151
R1455 B.n613 B.n611 10.6151
R1456 B.n614 B.n613 10.6151
R1457 B.n615 B.n614 10.6151
R1458 B.n616 B.n615 10.6151
R1459 B.n618 B.n616 10.6151
R1460 B.n619 B.n618 10.6151
R1461 B.n620 B.n619 10.6151
R1462 B.n621 B.n620 10.6151
R1463 B.n829 B.n1 10.6151
R1464 B.n829 B.n828 10.6151
R1465 B.n828 B.n827 10.6151
R1466 B.n827 B.n10 10.6151
R1467 B.n821 B.n10 10.6151
R1468 B.n821 B.n820 10.6151
R1469 B.n820 B.n819 10.6151
R1470 B.n819 B.n18 10.6151
R1471 B.n813 B.n18 10.6151
R1472 B.n813 B.n812 10.6151
R1473 B.n812 B.n811 10.6151
R1474 B.n811 B.n25 10.6151
R1475 B.n805 B.n25 10.6151
R1476 B.n805 B.n804 10.6151
R1477 B.n804 B.n803 10.6151
R1478 B.n803 B.n32 10.6151
R1479 B.n797 B.n32 10.6151
R1480 B.n797 B.n796 10.6151
R1481 B.n796 B.n795 10.6151
R1482 B.n795 B.n39 10.6151
R1483 B.n789 B.n39 10.6151
R1484 B.n789 B.n788 10.6151
R1485 B.n788 B.n787 10.6151
R1486 B.n787 B.n46 10.6151
R1487 B.n781 B.n46 10.6151
R1488 B.n781 B.n780 10.6151
R1489 B.n780 B.n779 10.6151
R1490 B.n779 B.n53 10.6151
R1491 B.n773 B.n53 10.6151
R1492 B.n773 B.n772 10.6151
R1493 B.n772 B.n771 10.6151
R1494 B.n771 B.n60 10.6151
R1495 B.n765 B.n60 10.6151
R1496 B.n765 B.n764 10.6151
R1497 B.n764 B.n763 10.6151
R1498 B.n763 B.n67 10.6151
R1499 B.n757 B.n67 10.6151
R1500 B.n757 B.n756 10.6151
R1501 B.n756 B.n755 10.6151
R1502 B.n755 B.n74 10.6151
R1503 B.n749 B.n74 10.6151
R1504 B.n749 B.n748 10.6151
R1505 B.n748 B.n747 10.6151
R1506 B.n747 B.n81 10.6151
R1507 B.n741 B.n81 10.6151
R1508 B.n741 B.n740 10.6151
R1509 B.n740 B.n739 10.6151
R1510 B.n739 B.n88 10.6151
R1511 B.n733 B.n88 10.6151
R1512 B.n733 B.n732 10.6151
R1513 B.n732 B.n731 10.6151
R1514 B.n731 B.n95 10.6151
R1515 B.n725 B.n95 10.6151
R1516 B.n725 B.n724 10.6151
R1517 B.n724 B.n723 10.6151
R1518 B.n723 B.n102 10.6151
R1519 B.n717 B.n102 10.6151
R1520 B.n716 B.n715 10.6151
R1521 B.n715 B.n109 10.6151
R1522 B.n709 B.n109 10.6151
R1523 B.n709 B.n708 10.6151
R1524 B.n708 B.n707 10.6151
R1525 B.n707 B.n111 10.6151
R1526 B.n701 B.n111 10.6151
R1527 B.n701 B.n700 10.6151
R1528 B.n700 B.n699 10.6151
R1529 B.n699 B.n113 10.6151
R1530 B.n693 B.n113 10.6151
R1531 B.n693 B.n692 10.6151
R1532 B.n692 B.n691 10.6151
R1533 B.n691 B.n115 10.6151
R1534 B.n685 B.n115 10.6151
R1535 B.n685 B.n684 10.6151
R1536 B.n684 B.n683 10.6151
R1537 B.n683 B.n117 10.6151
R1538 B.n677 B.n676 10.6151
R1539 B.n676 B.n675 10.6151
R1540 B.n675 B.n122 10.6151
R1541 B.n669 B.n122 10.6151
R1542 B.n669 B.n668 10.6151
R1543 B.n668 B.n667 10.6151
R1544 B.n667 B.n124 10.6151
R1545 B.n661 B.n124 10.6151
R1546 B.n659 B.n658 10.6151
R1547 B.n658 B.n128 10.6151
R1548 B.n652 B.n128 10.6151
R1549 B.n652 B.n651 10.6151
R1550 B.n651 B.n650 10.6151
R1551 B.n650 B.n130 10.6151
R1552 B.n644 B.n130 10.6151
R1553 B.n644 B.n643 10.6151
R1554 B.n643 B.n642 10.6151
R1555 B.n642 B.n132 10.6151
R1556 B.n636 B.n132 10.6151
R1557 B.n636 B.n635 10.6151
R1558 B.n635 B.n634 10.6151
R1559 B.n634 B.n134 10.6151
R1560 B.n628 B.n134 10.6151
R1561 B.n628 B.n627 10.6151
R1562 B.n627 B.n626 10.6151
R1563 B.n626 B.n622 10.6151
R1564 B.n837 B.n0 8.11757
R1565 B.n837 B.n1 8.11757
R1566 B.n334 B.n333 6.5566
R1567 B.n317 B.n316 6.5566
R1568 B.n677 B.n121 6.5566
R1569 B.n661 B.n660 6.5566
R1570 B.n488 B.t5 5.76268
R1571 B.n793 B.t1 5.76268
R1572 B.n335 B.n334 4.05904
R1573 B.n316 B.n315 4.05904
R1574 B.n121 B.n117 4.05904
R1575 B.n660 B.n659 4.05904
R1576 VP.n18 VP.n17 161.3
R1577 VP.n19 VP.n14 161.3
R1578 VP.n21 VP.n20 161.3
R1579 VP.n22 VP.n13 161.3
R1580 VP.n24 VP.n23 161.3
R1581 VP.n25 VP.n12 161.3
R1582 VP.n27 VP.n26 161.3
R1583 VP.n28 VP.n11 161.3
R1584 VP.n30 VP.n29 161.3
R1585 VP.n61 VP.n60 161.3
R1586 VP.n59 VP.n1 161.3
R1587 VP.n58 VP.n57 161.3
R1588 VP.n56 VP.n2 161.3
R1589 VP.n55 VP.n54 161.3
R1590 VP.n53 VP.n3 161.3
R1591 VP.n52 VP.n51 161.3
R1592 VP.n50 VP.n4 161.3
R1593 VP.n49 VP.n48 161.3
R1594 VP.n46 VP.n5 161.3
R1595 VP.n45 VP.n44 161.3
R1596 VP.n43 VP.n6 161.3
R1597 VP.n42 VP.n41 161.3
R1598 VP.n40 VP.n7 161.3
R1599 VP.n39 VP.n38 161.3
R1600 VP.n37 VP.n8 161.3
R1601 VP.n36 VP.n35 161.3
R1602 VP.n34 VP.n9 161.3
R1603 VP.n33 VP.n32 87.6207
R1604 VP.n62 VP.n0 87.6207
R1605 VP.n31 VP.n10 87.6207
R1606 VP.n16 VP.n15 62.9379
R1607 VP.n15 VP.t1 58.6115
R1608 VP.n41 VP.n40 50.2061
R1609 VP.n54 VP.n53 50.2061
R1610 VP.n23 VP.n22 50.2061
R1611 VP.n32 VP.n31 48.2796
R1612 VP.n40 VP.n39 30.7807
R1613 VP.n54 VP.n2 30.7807
R1614 VP.n23 VP.n12 30.7807
R1615 VP.n33 VP.t3 25.9217
R1616 VP.n47 VP.t4 25.9217
R1617 VP.n0 VP.t5 25.9217
R1618 VP.n10 VP.t2 25.9217
R1619 VP.n16 VP.t0 25.9217
R1620 VP.n35 VP.n34 24.4675
R1621 VP.n35 VP.n8 24.4675
R1622 VP.n39 VP.n8 24.4675
R1623 VP.n41 VP.n6 24.4675
R1624 VP.n45 VP.n6 24.4675
R1625 VP.n46 VP.n45 24.4675
R1626 VP.n48 VP.n4 24.4675
R1627 VP.n52 VP.n4 24.4675
R1628 VP.n53 VP.n52 24.4675
R1629 VP.n58 VP.n2 24.4675
R1630 VP.n59 VP.n58 24.4675
R1631 VP.n60 VP.n59 24.4675
R1632 VP.n27 VP.n12 24.4675
R1633 VP.n28 VP.n27 24.4675
R1634 VP.n29 VP.n28 24.4675
R1635 VP.n17 VP.n14 24.4675
R1636 VP.n21 VP.n14 24.4675
R1637 VP.n22 VP.n21 24.4675
R1638 VP.n47 VP.n46 12.234
R1639 VP.n48 VP.n47 12.234
R1640 VP.n17 VP.n16 12.234
R1641 VP.n18 VP.n15 2.47756
R1642 VP.n34 VP.n33 2.4472
R1643 VP.n60 VP.n0 2.4472
R1644 VP.n29 VP.n10 2.4472
R1645 VP.n31 VP.n30 0.354971
R1646 VP.n32 VP.n9 0.354971
R1647 VP.n62 VP.n61 0.354971
R1648 VP VP.n62 0.26696
R1649 VP.n19 VP.n18 0.189894
R1650 VP.n20 VP.n19 0.189894
R1651 VP.n20 VP.n13 0.189894
R1652 VP.n24 VP.n13 0.189894
R1653 VP.n25 VP.n24 0.189894
R1654 VP.n26 VP.n25 0.189894
R1655 VP.n26 VP.n11 0.189894
R1656 VP.n30 VP.n11 0.189894
R1657 VP.n36 VP.n9 0.189894
R1658 VP.n37 VP.n36 0.189894
R1659 VP.n38 VP.n37 0.189894
R1660 VP.n38 VP.n7 0.189894
R1661 VP.n42 VP.n7 0.189894
R1662 VP.n43 VP.n42 0.189894
R1663 VP.n44 VP.n43 0.189894
R1664 VP.n44 VP.n5 0.189894
R1665 VP.n49 VP.n5 0.189894
R1666 VP.n50 VP.n49 0.189894
R1667 VP.n51 VP.n50 0.189894
R1668 VP.n51 VP.n3 0.189894
R1669 VP.n55 VP.n3 0.189894
R1670 VP.n56 VP.n55 0.189894
R1671 VP.n57 VP.n56 0.189894
R1672 VP.n57 VP.n1 0.189894
R1673 VP.n61 VP.n1 0.189894
R1674 VDD1 VDD1.t4 80.7514
R1675 VDD1.n1 VDD1.t2 80.6376
R1676 VDD1.n1 VDD1.n0 74.1472
R1677 VDD1.n3 VDD1.n2 73.2759
R1678 VDD1.n3 VDD1.n1 41.8802
R1679 VDD1.n2 VDD1.t5 4.6375
R1680 VDD1.n2 VDD1.t3 4.6375
R1681 VDD1.n0 VDD1.t1 4.6375
R1682 VDD1.n0 VDD1.t0 4.6375
R1683 VDD1 VDD1.n3 0.869035
C0 VDD1 VP 3.24349f
C1 VN VDD2 2.82428f
C2 VTAIL VP 3.94427f
C3 VTAIL VDD1 5.82151f
C4 VDD2 VP 0.578545f
C5 VDD1 VDD2 1.94096f
C6 VN VP 6.83061f
C7 VTAIL VDD2 5.88372f
C8 VN VDD1 0.156718f
C9 VTAIL VN 3.92989f
C10 VDD2 B 5.666094f
C11 VDD1 B 6.047897f
C12 VTAIL B 5.047755f
C13 VN B 16.22296f
C14 VP B 14.862272f
C15 VDD1.t4 B 0.789716f
C16 VDD1.t2 B 0.788843f
C17 VDD1.t1 B 0.076667f
C18 VDD1.t0 B 0.076667f
C19 VDD1.n0 B 0.615479f
C20 VDD1.n1 B 2.85747f
C21 VDD1.t5 B 0.076667f
C22 VDD1.t3 B 0.076667f
C23 VDD1.n2 B 0.609333f
C24 VDD1.n3 B 2.33746f
C25 VP.t5 B 1.01911f
C26 VP.n0 B 0.480363f
C27 VP.n1 B 0.023268f
C28 VP.n2 B 0.046614f
C29 VP.n3 B 0.023268f
C30 VP.n4 B 0.043366f
C31 VP.n5 B 0.023268f
C32 VP.t4 B 1.01911f
C33 VP.n6 B 0.043366f
C34 VP.n7 B 0.023268f
C35 VP.n8 B 0.043366f
C36 VP.n9 B 0.037554f
C37 VP.t3 B 1.01911f
C38 VP.t2 B 1.01911f
C39 VP.n10 B 0.480363f
C40 VP.n11 B 0.023268f
C41 VP.n12 B 0.046614f
C42 VP.n13 B 0.023268f
C43 VP.n14 B 0.043366f
C44 VP.t1 B 1.34233f
C45 VP.n15 B 0.481952f
C46 VP.t0 B 1.01911f
C47 VP.n16 B 0.474772f
C48 VP.n17 B 0.032661f
C49 VP.n18 B 0.304363f
C50 VP.n19 B 0.023268f
C51 VP.n20 B 0.023268f
C52 VP.n21 B 0.043366f
C53 VP.n22 B 0.042706f
C54 VP.n23 B 0.021981f
C55 VP.n24 B 0.023268f
C56 VP.n25 B 0.023268f
C57 VP.n26 B 0.023268f
C58 VP.n27 B 0.043366f
C59 VP.n28 B 0.043366f
C60 VP.n29 B 0.024097f
C61 VP.n30 B 0.037554f
C62 VP.n31 B 1.27738f
C63 VP.n32 B 1.29471f
C64 VP.n33 B 0.480363f
C65 VP.n34 B 0.024097f
C66 VP.n35 B 0.043366f
C67 VP.n36 B 0.023268f
C68 VP.n37 B 0.023268f
C69 VP.n38 B 0.023268f
C70 VP.n39 B 0.046614f
C71 VP.n40 B 0.021981f
C72 VP.n41 B 0.042706f
C73 VP.n42 B 0.023268f
C74 VP.n43 B 0.023268f
C75 VP.n44 B 0.023268f
C76 VP.n45 B 0.043366f
C77 VP.n46 B 0.032661f
C78 VP.n47 B 0.389878f
C79 VP.n48 B 0.032661f
C80 VP.n49 B 0.023268f
C81 VP.n50 B 0.023268f
C82 VP.n51 B 0.023268f
C83 VP.n52 B 0.043366f
C84 VP.n53 B 0.042706f
C85 VP.n54 B 0.021981f
C86 VP.n55 B 0.023268f
C87 VP.n56 B 0.023268f
C88 VP.n57 B 0.023268f
C89 VP.n58 B 0.043366f
C90 VP.n59 B 0.043366f
C91 VP.n60 B 0.024097f
C92 VP.n61 B 0.037554f
C93 VP.n62 B 0.074003f
C94 VTAIL.t4 B 0.104593f
C95 VTAIL.t7 B 0.104593f
C96 VTAIL.n0 B 0.761468f
C97 VTAIL.n1 B 0.600919f
C98 VTAIL.t0 B 0.975379f
C99 VTAIL.n2 B 0.944135f
C100 VTAIL.t11 B 0.104593f
C101 VTAIL.t10 B 0.104593f
C102 VTAIL.n3 B 0.761468f
C103 VTAIL.n4 B 2.16995f
C104 VTAIL.t5 B 0.104593f
C105 VTAIL.t8 B 0.104593f
C106 VTAIL.n5 B 0.761472f
C107 VTAIL.n6 B 2.16995f
C108 VTAIL.t3 B 0.975383f
C109 VTAIL.n7 B 0.944131f
C110 VTAIL.t2 B 0.104593f
C111 VTAIL.t1 B 0.104593f
C112 VTAIL.n8 B 0.761472f
C113 VTAIL.n9 B 0.872787f
C114 VTAIL.t9 B 0.975379f
C115 VTAIL.n10 B 1.87105f
C116 VTAIL.t6 B 0.975379f
C117 VTAIL.n11 B 1.77268f
C118 VDD2.t0 B 0.769725f
C119 VDD2.t5 B 0.074809f
C120 VDD2.t4 B 0.074809f
C121 VDD2.n0 B 0.600563f
C122 VDD2.n1 B 2.65373f
C123 VDD2.t1 B 0.755517f
C124 VDD2.n2 B 2.25239f
C125 VDD2.t2 B 0.074809f
C126 VDD2.t3 B 0.074809f
C127 VDD2.n3 B 0.600534f
C128 VN.t2 B 0.987461f
C129 VN.n0 B 0.465444f
C130 VN.n1 B 0.022545f
C131 VN.n2 B 0.045166f
C132 VN.n3 B 0.022545f
C133 VN.n4 B 0.042019f
C134 VN.t4 B 1.30064f
C135 VN.n5 B 0.466984f
C136 VN.t1 B 0.987461f
C137 VN.n6 B 0.460027f
C138 VN.n7 B 0.031647f
C139 VN.n8 B 0.29491f
C140 VN.n9 B 0.022545f
C141 VN.n10 B 0.022545f
C142 VN.n11 B 0.042019f
C143 VN.n12 B 0.041379f
C144 VN.n13 B 0.021298f
C145 VN.n14 B 0.022545f
C146 VN.n15 B 0.022545f
C147 VN.n16 B 0.022545f
C148 VN.n17 B 0.042019f
C149 VN.n18 B 0.042019f
C150 VN.n19 B 0.023349f
C151 VN.n20 B 0.036388f
C152 VN.n21 B 0.071704f
C153 VN.t3 B 0.987461f
C154 VN.n22 B 0.465444f
C155 VN.n23 B 0.022545f
C156 VN.n24 B 0.045166f
C157 VN.n25 B 0.022545f
C158 VN.n26 B 0.042019f
C159 VN.t5 B 1.30064f
C160 VN.n27 B 0.466984f
C161 VN.t0 B 0.987461f
C162 VN.n28 B 0.460027f
C163 VN.n29 B 0.031647f
C164 VN.n30 B 0.29491f
C165 VN.n31 B 0.022545f
C166 VN.n32 B 0.022545f
C167 VN.n33 B 0.042019f
C168 VN.n34 B 0.041379f
C169 VN.n35 B 0.021298f
C170 VN.n36 B 0.022545f
C171 VN.n37 B 0.022545f
C172 VN.n38 B 0.022545f
C173 VN.n39 B 0.042019f
C174 VN.n40 B 0.042019f
C175 VN.n41 B 0.023349f
C176 VN.n42 B 0.036388f
C177 VN.n43 B 1.24704f
.ends

