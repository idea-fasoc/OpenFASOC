* NGSPICE file created from diff_pair_sample_1416.ext - technology: sky130A

.subckt diff_pair_sample_1416 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0 ps=0 w=5.36 l=0.46
X1 VDD1.t9 VP.t0 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X2 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0 ps=0 w=5.36 l=0.46
X3 VDD2.t9 VN.t0 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0.8844 ps=5.69 w=5.36 l=0.46
X4 VTAIL.t18 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X5 VTAIL.t19 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X6 VDD2.t6 VN.t3 VTAIL.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=2.0904 ps=11.5 w=5.36 l=0.46
X7 VDD2.t5 VN.t4 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0.8844 ps=5.69 w=5.36 l=0.46
X8 VDD1.t8 VP.t1 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=2.0904 ps=11.5 w=5.36 l=0.46
X9 VTAIL.t14 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X10 VDD2.t4 VN.t5 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X11 VDD1.t6 VP.t3 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0.8844 ps=5.69 w=5.36 l=0.46
X12 VDD1.t5 VP.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=2.0904 ps=11.5 w=5.36 l=0.46
X13 VTAIL.t2 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X14 VTAIL.t12 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X15 VDD2.t2 VN.t7 VTAIL.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=2.0904 ps=11.5 w=5.36 l=0.46
X16 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0 ps=0 w=5.36 l=0.46
X17 VTAIL.t3 VN.t8 VDD2.t1 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0 ps=0 w=5.36 l=0.46
X19 VDD1.t3 VP.t6 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X20 VTAIL.t7 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X21 VDD1.t1 VP.t8 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.0904 pd=11.5 as=0.8844 ps=5.69 w=5.36 l=0.46
X22 VTAIL.t8 VP.t9 VDD1.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
X23 VDD2.t0 VN.t9 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8844 pd=5.69 as=0.8844 ps=5.69 w=5.36 l=0.46
R0 B.n355 B.n354 585
R1 B.n356 B.n76 585
R2 B.n358 B.n357 585
R3 B.n360 B.n75 585
R4 B.n363 B.n362 585
R5 B.n364 B.n74 585
R6 B.n366 B.n365 585
R7 B.n368 B.n73 585
R8 B.n371 B.n370 585
R9 B.n372 B.n72 585
R10 B.n374 B.n373 585
R11 B.n376 B.n71 585
R12 B.n379 B.n378 585
R13 B.n380 B.n70 585
R14 B.n382 B.n381 585
R15 B.n384 B.n69 585
R16 B.n387 B.n386 585
R17 B.n388 B.n68 585
R18 B.n390 B.n389 585
R19 B.n392 B.n67 585
R20 B.n394 B.n393 585
R21 B.n396 B.n395 585
R22 B.n399 B.n398 585
R23 B.n400 B.n62 585
R24 B.n402 B.n401 585
R25 B.n404 B.n61 585
R26 B.n407 B.n406 585
R27 B.n408 B.n60 585
R28 B.n410 B.n409 585
R29 B.n412 B.n59 585
R30 B.n414 B.n413 585
R31 B.n416 B.n415 585
R32 B.n419 B.n418 585
R33 B.n420 B.n54 585
R34 B.n422 B.n421 585
R35 B.n424 B.n53 585
R36 B.n427 B.n426 585
R37 B.n428 B.n52 585
R38 B.n430 B.n429 585
R39 B.n432 B.n51 585
R40 B.n435 B.n434 585
R41 B.n436 B.n50 585
R42 B.n438 B.n437 585
R43 B.n440 B.n49 585
R44 B.n443 B.n442 585
R45 B.n444 B.n48 585
R46 B.n446 B.n445 585
R47 B.n448 B.n47 585
R48 B.n451 B.n450 585
R49 B.n452 B.n46 585
R50 B.n454 B.n453 585
R51 B.n456 B.n45 585
R52 B.n459 B.n458 585
R53 B.n460 B.n44 585
R54 B.n352 B.n42 585
R55 B.n463 B.n42 585
R56 B.n351 B.n41 585
R57 B.n464 B.n41 585
R58 B.n350 B.n40 585
R59 B.n465 B.n40 585
R60 B.n349 B.n348 585
R61 B.n348 B.n36 585
R62 B.n347 B.n35 585
R63 B.n471 B.n35 585
R64 B.n346 B.n34 585
R65 B.n472 B.n34 585
R66 B.n345 B.n33 585
R67 B.n473 B.n33 585
R68 B.n344 B.n343 585
R69 B.n343 B.n29 585
R70 B.n342 B.n28 585
R71 B.n479 B.n28 585
R72 B.n341 B.n27 585
R73 B.n480 B.n27 585
R74 B.n340 B.n26 585
R75 B.n481 B.n26 585
R76 B.n339 B.n338 585
R77 B.n338 B.n22 585
R78 B.n337 B.n21 585
R79 B.n487 B.n21 585
R80 B.n336 B.n20 585
R81 B.n488 B.n20 585
R82 B.n335 B.n19 585
R83 B.n489 B.n19 585
R84 B.n334 B.n333 585
R85 B.n333 B.n15 585
R86 B.n332 B.n14 585
R87 B.n495 B.n14 585
R88 B.n331 B.n13 585
R89 B.n496 B.n13 585
R90 B.n330 B.n12 585
R91 B.n497 B.n12 585
R92 B.n329 B.n328 585
R93 B.n328 B.n11 585
R94 B.n327 B.n7 585
R95 B.n503 B.n7 585
R96 B.n326 B.n6 585
R97 B.n504 B.n6 585
R98 B.n325 B.n5 585
R99 B.n505 B.n5 585
R100 B.n324 B.n323 585
R101 B.n323 B.n4 585
R102 B.n322 B.n77 585
R103 B.n322 B.n321 585
R104 B.n311 B.n78 585
R105 B.n314 B.n78 585
R106 B.n313 B.n312 585
R107 B.n315 B.n313 585
R108 B.n310 B.n83 585
R109 B.n83 B.n82 585
R110 B.n309 B.n308 585
R111 B.n308 B.n307 585
R112 B.n85 B.n84 585
R113 B.n86 B.n85 585
R114 B.n300 B.n299 585
R115 B.n301 B.n300 585
R116 B.n298 B.n91 585
R117 B.n91 B.n90 585
R118 B.n297 B.n296 585
R119 B.n296 B.n295 585
R120 B.n93 B.n92 585
R121 B.n94 B.n93 585
R122 B.n288 B.n287 585
R123 B.n289 B.n288 585
R124 B.n286 B.n98 585
R125 B.n102 B.n98 585
R126 B.n285 B.n284 585
R127 B.n284 B.n283 585
R128 B.n100 B.n99 585
R129 B.n101 B.n100 585
R130 B.n276 B.n275 585
R131 B.n277 B.n276 585
R132 B.n274 B.n107 585
R133 B.n107 B.n106 585
R134 B.n273 B.n272 585
R135 B.n272 B.n271 585
R136 B.n109 B.n108 585
R137 B.n110 B.n109 585
R138 B.n264 B.n263 585
R139 B.n265 B.n264 585
R140 B.n262 B.n115 585
R141 B.n115 B.n114 585
R142 B.n261 B.n260 585
R143 B.n260 B.n259 585
R144 B.n256 B.n119 585
R145 B.n255 B.n254 585
R146 B.n252 B.n120 585
R147 B.n252 B.n118 585
R148 B.n251 B.n250 585
R149 B.n249 B.n248 585
R150 B.n247 B.n122 585
R151 B.n245 B.n244 585
R152 B.n243 B.n123 585
R153 B.n242 B.n241 585
R154 B.n239 B.n124 585
R155 B.n237 B.n236 585
R156 B.n235 B.n125 585
R157 B.n234 B.n233 585
R158 B.n231 B.n126 585
R159 B.n229 B.n228 585
R160 B.n227 B.n127 585
R161 B.n226 B.n225 585
R162 B.n223 B.n128 585
R163 B.n221 B.n220 585
R164 B.n219 B.n129 585
R165 B.n218 B.n217 585
R166 B.n215 B.n130 585
R167 B.n213 B.n212 585
R168 B.n211 B.n131 585
R169 B.n210 B.n209 585
R170 B.n207 B.n135 585
R171 B.n205 B.n204 585
R172 B.n203 B.n136 585
R173 B.n202 B.n201 585
R174 B.n199 B.n137 585
R175 B.n197 B.n196 585
R176 B.n195 B.n138 585
R177 B.n193 B.n192 585
R178 B.n190 B.n141 585
R179 B.n188 B.n187 585
R180 B.n186 B.n142 585
R181 B.n185 B.n184 585
R182 B.n182 B.n143 585
R183 B.n180 B.n179 585
R184 B.n178 B.n144 585
R185 B.n177 B.n176 585
R186 B.n174 B.n145 585
R187 B.n172 B.n171 585
R188 B.n170 B.n146 585
R189 B.n169 B.n168 585
R190 B.n166 B.n147 585
R191 B.n164 B.n163 585
R192 B.n162 B.n148 585
R193 B.n161 B.n160 585
R194 B.n158 B.n149 585
R195 B.n156 B.n155 585
R196 B.n154 B.n150 585
R197 B.n153 B.n152 585
R198 B.n117 B.n116 585
R199 B.n118 B.n117 585
R200 B.n258 B.n257 585
R201 B.n259 B.n258 585
R202 B.n113 B.n112 585
R203 B.n114 B.n113 585
R204 B.n267 B.n266 585
R205 B.n266 B.n265 585
R206 B.n268 B.n111 585
R207 B.n111 B.n110 585
R208 B.n270 B.n269 585
R209 B.n271 B.n270 585
R210 B.n105 B.n104 585
R211 B.n106 B.n105 585
R212 B.n279 B.n278 585
R213 B.n278 B.n277 585
R214 B.n280 B.n103 585
R215 B.n103 B.n101 585
R216 B.n282 B.n281 585
R217 B.n283 B.n282 585
R218 B.n97 B.n96 585
R219 B.n102 B.n97 585
R220 B.n291 B.n290 585
R221 B.n290 B.n289 585
R222 B.n292 B.n95 585
R223 B.n95 B.n94 585
R224 B.n294 B.n293 585
R225 B.n295 B.n294 585
R226 B.n89 B.n88 585
R227 B.n90 B.n89 585
R228 B.n303 B.n302 585
R229 B.n302 B.n301 585
R230 B.n304 B.n87 585
R231 B.n87 B.n86 585
R232 B.n306 B.n305 585
R233 B.n307 B.n306 585
R234 B.n81 B.n80 585
R235 B.n82 B.n81 585
R236 B.n317 B.n316 585
R237 B.n316 B.n315 585
R238 B.n318 B.n79 585
R239 B.n314 B.n79 585
R240 B.n320 B.n319 585
R241 B.n321 B.n320 585
R242 B.n2 B.n0 585
R243 B.n4 B.n2 585
R244 B.n3 B.n1 585
R245 B.n504 B.n3 585
R246 B.n502 B.n501 585
R247 B.n503 B.n502 585
R248 B.n500 B.n8 585
R249 B.n11 B.n8 585
R250 B.n499 B.n498 585
R251 B.n498 B.n497 585
R252 B.n10 B.n9 585
R253 B.n496 B.n10 585
R254 B.n494 B.n493 585
R255 B.n495 B.n494 585
R256 B.n492 B.n16 585
R257 B.n16 B.n15 585
R258 B.n491 B.n490 585
R259 B.n490 B.n489 585
R260 B.n18 B.n17 585
R261 B.n488 B.n18 585
R262 B.n486 B.n485 585
R263 B.n487 B.n486 585
R264 B.n484 B.n23 585
R265 B.n23 B.n22 585
R266 B.n483 B.n482 585
R267 B.n482 B.n481 585
R268 B.n25 B.n24 585
R269 B.n480 B.n25 585
R270 B.n478 B.n477 585
R271 B.n479 B.n478 585
R272 B.n476 B.n30 585
R273 B.n30 B.n29 585
R274 B.n475 B.n474 585
R275 B.n474 B.n473 585
R276 B.n32 B.n31 585
R277 B.n472 B.n32 585
R278 B.n470 B.n469 585
R279 B.n471 B.n470 585
R280 B.n468 B.n37 585
R281 B.n37 B.n36 585
R282 B.n467 B.n466 585
R283 B.n466 B.n465 585
R284 B.n39 B.n38 585
R285 B.n464 B.n39 585
R286 B.n462 B.n461 585
R287 B.n463 B.n462 585
R288 B.n507 B.n506 585
R289 B.n506 B.n505 585
R290 B.n139 B.t14 488.274
R291 B.n132 B.t21 488.274
R292 B.n55 B.t18 488.274
R293 B.n63 B.t10 488.274
R294 B.n258 B.n119 487.695
R295 B.n462 B.n44 487.695
R296 B.n260 B.n117 487.695
R297 B.n354 B.n42 487.695
R298 B.n353 B.n43 256.663
R299 B.n359 B.n43 256.663
R300 B.n361 B.n43 256.663
R301 B.n367 B.n43 256.663
R302 B.n369 B.n43 256.663
R303 B.n375 B.n43 256.663
R304 B.n377 B.n43 256.663
R305 B.n383 B.n43 256.663
R306 B.n385 B.n43 256.663
R307 B.n391 B.n43 256.663
R308 B.n66 B.n43 256.663
R309 B.n397 B.n43 256.663
R310 B.n403 B.n43 256.663
R311 B.n405 B.n43 256.663
R312 B.n411 B.n43 256.663
R313 B.n58 B.n43 256.663
R314 B.n417 B.n43 256.663
R315 B.n423 B.n43 256.663
R316 B.n425 B.n43 256.663
R317 B.n431 B.n43 256.663
R318 B.n433 B.n43 256.663
R319 B.n439 B.n43 256.663
R320 B.n441 B.n43 256.663
R321 B.n447 B.n43 256.663
R322 B.n449 B.n43 256.663
R323 B.n455 B.n43 256.663
R324 B.n457 B.n43 256.663
R325 B.n253 B.n118 256.663
R326 B.n121 B.n118 256.663
R327 B.n246 B.n118 256.663
R328 B.n240 B.n118 256.663
R329 B.n238 B.n118 256.663
R330 B.n232 B.n118 256.663
R331 B.n230 B.n118 256.663
R332 B.n224 B.n118 256.663
R333 B.n222 B.n118 256.663
R334 B.n216 B.n118 256.663
R335 B.n214 B.n118 256.663
R336 B.n208 B.n118 256.663
R337 B.n206 B.n118 256.663
R338 B.n200 B.n118 256.663
R339 B.n198 B.n118 256.663
R340 B.n191 B.n118 256.663
R341 B.n189 B.n118 256.663
R342 B.n183 B.n118 256.663
R343 B.n181 B.n118 256.663
R344 B.n175 B.n118 256.663
R345 B.n173 B.n118 256.663
R346 B.n167 B.n118 256.663
R347 B.n165 B.n118 256.663
R348 B.n159 B.n118 256.663
R349 B.n157 B.n118 256.663
R350 B.n151 B.n118 256.663
R351 B.n139 B.t17 183.446
R352 B.n63 B.t12 183.446
R353 B.n132 B.t23 183.446
R354 B.n55 B.t19 183.446
R355 B.n140 B.t16 168.125
R356 B.n64 B.t13 168.125
R357 B.n133 B.t22 168.125
R358 B.n56 B.t20 168.125
R359 B.n258 B.n113 163.367
R360 B.n266 B.n113 163.367
R361 B.n266 B.n111 163.367
R362 B.n270 B.n111 163.367
R363 B.n270 B.n105 163.367
R364 B.n278 B.n105 163.367
R365 B.n278 B.n103 163.367
R366 B.n282 B.n103 163.367
R367 B.n282 B.n97 163.367
R368 B.n290 B.n97 163.367
R369 B.n290 B.n95 163.367
R370 B.n294 B.n95 163.367
R371 B.n294 B.n89 163.367
R372 B.n302 B.n89 163.367
R373 B.n302 B.n87 163.367
R374 B.n306 B.n87 163.367
R375 B.n306 B.n81 163.367
R376 B.n316 B.n81 163.367
R377 B.n316 B.n79 163.367
R378 B.n320 B.n79 163.367
R379 B.n320 B.n2 163.367
R380 B.n506 B.n2 163.367
R381 B.n506 B.n3 163.367
R382 B.n502 B.n3 163.367
R383 B.n502 B.n8 163.367
R384 B.n498 B.n8 163.367
R385 B.n498 B.n10 163.367
R386 B.n494 B.n10 163.367
R387 B.n494 B.n16 163.367
R388 B.n490 B.n16 163.367
R389 B.n490 B.n18 163.367
R390 B.n486 B.n18 163.367
R391 B.n486 B.n23 163.367
R392 B.n482 B.n23 163.367
R393 B.n482 B.n25 163.367
R394 B.n478 B.n25 163.367
R395 B.n478 B.n30 163.367
R396 B.n474 B.n30 163.367
R397 B.n474 B.n32 163.367
R398 B.n470 B.n32 163.367
R399 B.n470 B.n37 163.367
R400 B.n466 B.n37 163.367
R401 B.n466 B.n39 163.367
R402 B.n462 B.n39 163.367
R403 B.n254 B.n252 163.367
R404 B.n252 B.n251 163.367
R405 B.n248 B.n247 163.367
R406 B.n245 B.n123 163.367
R407 B.n241 B.n239 163.367
R408 B.n237 B.n125 163.367
R409 B.n233 B.n231 163.367
R410 B.n229 B.n127 163.367
R411 B.n225 B.n223 163.367
R412 B.n221 B.n129 163.367
R413 B.n217 B.n215 163.367
R414 B.n213 B.n131 163.367
R415 B.n209 B.n207 163.367
R416 B.n205 B.n136 163.367
R417 B.n201 B.n199 163.367
R418 B.n197 B.n138 163.367
R419 B.n192 B.n190 163.367
R420 B.n188 B.n142 163.367
R421 B.n184 B.n182 163.367
R422 B.n180 B.n144 163.367
R423 B.n176 B.n174 163.367
R424 B.n172 B.n146 163.367
R425 B.n168 B.n166 163.367
R426 B.n164 B.n148 163.367
R427 B.n160 B.n158 163.367
R428 B.n156 B.n150 163.367
R429 B.n152 B.n117 163.367
R430 B.n260 B.n115 163.367
R431 B.n264 B.n115 163.367
R432 B.n264 B.n109 163.367
R433 B.n272 B.n109 163.367
R434 B.n272 B.n107 163.367
R435 B.n276 B.n107 163.367
R436 B.n276 B.n100 163.367
R437 B.n284 B.n100 163.367
R438 B.n284 B.n98 163.367
R439 B.n288 B.n98 163.367
R440 B.n288 B.n93 163.367
R441 B.n296 B.n93 163.367
R442 B.n296 B.n91 163.367
R443 B.n300 B.n91 163.367
R444 B.n300 B.n85 163.367
R445 B.n308 B.n85 163.367
R446 B.n308 B.n83 163.367
R447 B.n313 B.n83 163.367
R448 B.n313 B.n78 163.367
R449 B.n322 B.n78 163.367
R450 B.n323 B.n322 163.367
R451 B.n323 B.n5 163.367
R452 B.n6 B.n5 163.367
R453 B.n7 B.n6 163.367
R454 B.n328 B.n7 163.367
R455 B.n328 B.n12 163.367
R456 B.n13 B.n12 163.367
R457 B.n14 B.n13 163.367
R458 B.n333 B.n14 163.367
R459 B.n333 B.n19 163.367
R460 B.n20 B.n19 163.367
R461 B.n21 B.n20 163.367
R462 B.n338 B.n21 163.367
R463 B.n338 B.n26 163.367
R464 B.n27 B.n26 163.367
R465 B.n28 B.n27 163.367
R466 B.n343 B.n28 163.367
R467 B.n343 B.n33 163.367
R468 B.n34 B.n33 163.367
R469 B.n35 B.n34 163.367
R470 B.n348 B.n35 163.367
R471 B.n348 B.n40 163.367
R472 B.n41 B.n40 163.367
R473 B.n42 B.n41 163.367
R474 B.n458 B.n456 163.367
R475 B.n454 B.n46 163.367
R476 B.n450 B.n448 163.367
R477 B.n446 B.n48 163.367
R478 B.n442 B.n440 163.367
R479 B.n438 B.n50 163.367
R480 B.n434 B.n432 163.367
R481 B.n430 B.n52 163.367
R482 B.n426 B.n424 163.367
R483 B.n422 B.n54 163.367
R484 B.n418 B.n416 163.367
R485 B.n413 B.n412 163.367
R486 B.n410 B.n60 163.367
R487 B.n406 B.n404 163.367
R488 B.n402 B.n62 163.367
R489 B.n398 B.n396 163.367
R490 B.n393 B.n392 163.367
R491 B.n390 B.n68 163.367
R492 B.n386 B.n384 163.367
R493 B.n382 B.n70 163.367
R494 B.n378 B.n376 163.367
R495 B.n374 B.n72 163.367
R496 B.n370 B.n368 163.367
R497 B.n366 B.n74 163.367
R498 B.n362 B.n360 163.367
R499 B.n358 B.n76 163.367
R500 B.n259 B.n118 131.359
R501 B.n463 B.n43 131.359
R502 B.n253 B.n119 71.676
R503 B.n251 B.n121 71.676
R504 B.n247 B.n246 71.676
R505 B.n240 B.n123 71.676
R506 B.n239 B.n238 71.676
R507 B.n232 B.n125 71.676
R508 B.n231 B.n230 71.676
R509 B.n224 B.n127 71.676
R510 B.n223 B.n222 71.676
R511 B.n216 B.n129 71.676
R512 B.n215 B.n214 71.676
R513 B.n208 B.n131 71.676
R514 B.n207 B.n206 71.676
R515 B.n200 B.n136 71.676
R516 B.n199 B.n198 71.676
R517 B.n191 B.n138 71.676
R518 B.n190 B.n189 71.676
R519 B.n183 B.n142 71.676
R520 B.n182 B.n181 71.676
R521 B.n175 B.n144 71.676
R522 B.n174 B.n173 71.676
R523 B.n167 B.n146 71.676
R524 B.n166 B.n165 71.676
R525 B.n159 B.n148 71.676
R526 B.n158 B.n157 71.676
R527 B.n151 B.n150 71.676
R528 B.n457 B.n44 71.676
R529 B.n456 B.n455 71.676
R530 B.n449 B.n46 71.676
R531 B.n448 B.n447 71.676
R532 B.n441 B.n48 71.676
R533 B.n440 B.n439 71.676
R534 B.n433 B.n50 71.676
R535 B.n432 B.n431 71.676
R536 B.n425 B.n52 71.676
R537 B.n424 B.n423 71.676
R538 B.n417 B.n54 71.676
R539 B.n416 B.n58 71.676
R540 B.n412 B.n411 71.676
R541 B.n405 B.n60 71.676
R542 B.n404 B.n403 71.676
R543 B.n397 B.n62 71.676
R544 B.n396 B.n66 71.676
R545 B.n392 B.n391 71.676
R546 B.n385 B.n68 71.676
R547 B.n384 B.n383 71.676
R548 B.n377 B.n70 71.676
R549 B.n376 B.n375 71.676
R550 B.n369 B.n72 71.676
R551 B.n368 B.n367 71.676
R552 B.n361 B.n74 71.676
R553 B.n360 B.n359 71.676
R554 B.n353 B.n76 71.676
R555 B.n354 B.n353 71.676
R556 B.n359 B.n358 71.676
R557 B.n362 B.n361 71.676
R558 B.n367 B.n366 71.676
R559 B.n370 B.n369 71.676
R560 B.n375 B.n374 71.676
R561 B.n378 B.n377 71.676
R562 B.n383 B.n382 71.676
R563 B.n386 B.n385 71.676
R564 B.n391 B.n390 71.676
R565 B.n393 B.n66 71.676
R566 B.n398 B.n397 71.676
R567 B.n403 B.n402 71.676
R568 B.n406 B.n405 71.676
R569 B.n411 B.n410 71.676
R570 B.n413 B.n58 71.676
R571 B.n418 B.n417 71.676
R572 B.n423 B.n422 71.676
R573 B.n426 B.n425 71.676
R574 B.n431 B.n430 71.676
R575 B.n434 B.n433 71.676
R576 B.n439 B.n438 71.676
R577 B.n442 B.n441 71.676
R578 B.n447 B.n446 71.676
R579 B.n450 B.n449 71.676
R580 B.n455 B.n454 71.676
R581 B.n458 B.n457 71.676
R582 B.n254 B.n253 71.676
R583 B.n248 B.n121 71.676
R584 B.n246 B.n245 71.676
R585 B.n241 B.n240 71.676
R586 B.n238 B.n237 71.676
R587 B.n233 B.n232 71.676
R588 B.n230 B.n229 71.676
R589 B.n225 B.n224 71.676
R590 B.n222 B.n221 71.676
R591 B.n217 B.n216 71.676
R592 B.n214 B.n213 71.676
R593 B.n209 B.n208 71.676
R594 B.n206 B.n205 71.676
R595 B.n201 B.n200 71.676
R596 B.n198 B.n197 71.676
R597 B.n192 B.n191 71.676
R598 B.n189 B.n188 71.676
R599 B.n184 B.n183 71.676
R600 B.n181 B.n180 71.676
R601 B.n176 B.n175 71.676
R602 B.n173 B.n172 71.676
R603 B.n168 B.n167 71.676
R604 B.n165 B.n164 71.676
R605 B.n160 B.n159 71.676
R606 B.n157 B.n156 71.676
R607 B.n152 B.n151 71.676
R608 B.n259 B.n114 70.3343
R609 B.n265 B.n114 70.3343
R610 B.n265 B.n110 70.3343
R611 B.n271 B.n110 70.3343
R612 B.n277 B.n106 70.3343
R613 B.n277 B.n101 70.3343
R614 B.n283 B.n101 70.3343
R615 B.n283 B.n102 70.3343
R616 B.n289 B.n94 70.3343
R617 B.n295 B.n94 70.3343
R618 B.n301 B.n90 70.3343
R619 B.n307 B.n86 70.3343
R620 B.n315 B.n82 70.3343
R621 B.n315 B.n314 70.3343
R622 B.n321 B.n4 70.3343
R623 B.n505 B.n4 70.3343
R624 B.n505 B.n504 70.3343
R625 B.n504 B.n503 70.3343
R626 B.n497 B.n11 70.3343
R627 B.n497 B.n496 70.3343
R628 B.n495 B.n15 70.3343
R629 B.n489 B.n488 70.3343
R630 B.n487 B.n22 70.3343
R631 B.n481 B.n22 70.3343
R632 B.n480 B.n479 70.3343
R633 B.n479 B.n29 70.3343
R634 B.n473 B.n29 70.3343
R635 B.n473 B.n472 70.3343
R636 B.n471 B.n36 70.3343
R637 B.n465 B.n36 70.3343
R638 B.n465 B.n464 70.3343
R639 B.n464 B.n463 70.3343
R640 B.n102 B.t4 66.197
R641 B.t5 B.n480 66.197
R642 B.n307 B.t8 64.1284
R643 B.t3 B.n495 64.1284
R644 B.n194 B.n140 59.5399
R645 B.n134 B.n133 59.5399
R646 B.n57 B.n56 59.5399
R647 B.n65 B.n64 59.5399
R648 B.n321 B.t7 53.7852
R649 B.n503 B.t1 53.7852
R650 B.t2 B.n90 51.7165
R651 B.n488 B.t9 51.7165
R652 B.t15 B.n106 41.3733
R653 B.n301 B.t6 41.3733
R654 B.n489 B.t0 41.3733
R655 B.n472 B.t11 41.3733
R656 B.n461 B.n460 31.6883
R657 B.n355 B.n352 31.6883
R658 B.n261 B.n116 31.6883
R659 B.n257 B.n256 31.6883
R660 B.n271 B.t15 28.9615
R661 B.t6 B.n86 28.9615
R662 B.t0 B.n15 28.9615
R663 B.t11 B.n471 28.9615
R664 B.n295 B.t2 18.6183
R665 B.t9 B.n487 18.6183
R666 B B.n507 18.0485
R667 B.n314 B.t7 16.5496
R668 B.n11 B.t1 16.5496
R669 B.n140 B.n139 15.3217
R670 B.n133 B.n132 15.3217
R671 B.n56 B.n55 15.3217
R672 B.n64 B.n63 15.3217
R673 B.n460 B.n459 10.6151
R674 B.n459 B.n45 10.6151
R675 B.n453 B.n45 10.6151
R676 B.n453 B.n452 10.6151
R677 B.n452 B.n451 10.6151
R678 B.n451 B.n47 10.6151
R679 B.n445 B.n47 10.6151
R680 B.n445 B.n444 10.6151
R681 B.n444 B.n443 10.6151
R682 B.n443 B.n49 10.6151
R683 B.n437 B.n49 10.6151
R684 B.n437 B.n436 10.6151
R685 B.n436 B.n435 10.6151
R686 B.n435 B.n51 10.6151
R687 B.n429 B.n51 10.6151
R688 B.n429 B.n428 10.6151
R689 B.n428 B.n427 10.6151
R690 B.n427 B.n53 10.6151
R691 B.n421 B.n53 10.6151
R692 B.n421 B.n420 10.6151
R693 B.n420 B.n419 10.6151
R694 B.n415 B.n414 10.6151
R695 B.n414 B.n59 10.6151
R696 B.n409 B.n59 10.6151
R697 B.n409 B.n408 10.6151
R698 B.n408 B.n407 10.6151
R699 B.n407 B.n61 10.6151
R700 B.n401 B.n61 10.6151
R701 B.n401 B.n400 10.6151
R702 B.n400 B.n399 10.6151
R703 B.n395 B.n394 10.6151
R704 B.n394 B.n67 10.6151
R705 B.n389 B.n67 10.6151
R706 B.n389 B.n388 10.6151
R707 B.n388 B.n387 10.6151
R708 B.n387 B.n69 10.6151
R709 B.n381 B.n69 10.6151
R710 B.n381 B.n380 10.6151
R711 B.n380 B.n379 10.6151
R712 B.n379 B.n71 10.6151
R713 B.n373 B.n71 10.6151
R714 B.n373 B.n372 10.6151
R715 B.n372 B.n371 10.6151
R716 B.n371 B.n73 10.6151
R717 B.n365 B.n73 10.6151
R718 B.n365 B.n364 10.6151
R719 B.n364 B.n363 10.6151
R720 B.n363 B.n75 10.6151
R721 B.n357 B.n75 10.6151
R722 B.n357 B.n356 10.6151
R723 B.n356 B.n355 10.6151
R724 B.n262 B.n261 10.6151
R725 B.n263 B.n262 10.6151
R726 B.n263 B.n108 10.6151
R727 B.n273 B.n108 10.6151
R728 B.n274 B.n273 10.6151
R729 B.n275 B.n274 10.6151
R730 B.n275 B.n99 10.6151
R731 B.n285 B.n99 10.6151
R732 B.n286 B.n285 10.6151
R733 B.n287 B.n286 10.6151
R734 B.n287 B.n92 10.6151
R735 B.n297 B.n92 10.6151
R736 B.n298 B.n297 10.6151
R737 B.n299 B.n298 10.6151
R738 B.n299 B.n84 10.6151
R739 B.n309 B.n84 10.6151
R740 B.n310 B.n309 10.6151
R741 B.n312 B.n310 10.6151
R742 B.n312 B.n311 10.6151
R743 B.n311 B.n77 10.6151
R744 B.n324 B.n77 10.6151
R745 B.n325 B.n324 10.6151
R746 B.n326 B.n325 10.6151
R747 B.n327 B.n326 10.6151
R748 B.n329 B.n327 10.6151
R749 B.n330 B.n329 10.6151
R750 B.n331 B.n330 10.6151
R751 B.n332 B.n331 10.6151
R752 B.n334 B.n332 10.6151
R753 B.n335 B.n334 10.6151
R754 B.n336 B.n335 10.6151
R755 B.n337 B.n336 10.6151
R756 B.n339 B.n337 10.6151
R757 B.n340 B.n339 10.6151
R758 B.n341 B.n340 10.6151
R759 B.n342 B.n341 10.6151
R760 B.n344 B.n342 10.6151
R761 B.n345 B.n344 10.6151
R762 B.n346 B.n345 10.6151
R763 B.n347 B.n346 10.6151
R764 B.n349 B.n347 10.6151
R765 B.n350 B.n349 10.6151
R766 B.n351 B.n350 10.6151
R767 B.n352 B.n351 10.6151
R768 B.n256 B.n255 10.6151
R769 B.n255 B.n120 10.6151
R770 B.n250 B.n120 10.6151
R771 B.n250 B.n249 10.6151
R772 B.n249 B.n122 10.6151
R773 B.n244 B.n122 10.6151
R774 B.n244 B.n243 10.6151
R775 B.n243 B.n242 10.6151
R776 B.n242 B.n124 10.6151
R777 B.n236 B.n124 10.6151
R778 B.n236 B.n235 10.6151
R779 B.n235 B.n234 10.6151
R780 B.n234 B.n126 10.6151
R781 B.n228 B.n126 10.6151
R782 B.n228 B.n227 10.6151
R783 B.n227 B.n226 10.6151
R784 B.n226 B.n128 10.6151
R785 B.n220 B.n128 10.6151
R786 B.n220 B.n219 10.6151
R787 B.n219 B.n218 10.6151
R788 B.n218 B.n130 10.6151
R789 B.n212 B.n211 10.6151
R790 B.n211 B.n210 10.6151
R791 B.n210 B.n135 10.6151
R792 B.n204 B.n135 10.6151
R793 B.n204 B.n203 10.6151
R794 B.n203 B.n202 10.6151
R795 B.n202 B.n137 10.6151
R796 B.n196 B.n137 10.6151
R797 B.n196 B.n195 10.6151
R798 B.n193 B.n141 10.6151
R799 B.n187 B.n141 10.6151
R800 B.n187 B.n186 10.6151
R801 B.n186 B.n185 10.6151
R802 B.n185 B.n143 10.6151
R803 B.n179 B.n143 10.6151
R804 B.n179 B.n178 10.6151
R805 B.n178 B.n177 10.6151
R806 B.n177 B.n145 10.6151
R807 B.n171 B.n145 10.6151
R808 B.n171 B.n170 10.6151
R809 B.n170 B.n169 10.6151
R810 B.n169 B.n147 10.6151
R811 B.n163 B.n147 10.6151
R812 B.n163 B.n162 10.6151
R813 B.n162 B.n161 10.6151
R814 B.n161 B.n149 10.6151
R815 B.n155 B.n149 10.6151
R816 B.n155 B.n154 10.6151
R817 B.n154 B.n153 10.6151
R818 B.n153 B.n116 10.6151
R819 B.n257 B.n112 10.6151
R820 B.n267 B.n112 10.6151
R821 B.n268 B.n267 10.6151
R822 B.n269 B.n268 10.6151
R823 B.n269 B.n104 10.6151
R824 B.n279 B.n104 10.6151
R825 B.n280 B.n279 10.6151
R826 B.n281 B.n280 10.6151
R827 B.n281 B.n96 10.6151
R828 B.n291 B.n96 10.6151
R829 B.n292 B.n291 10.6151
R830 B.n293 B.n292 10.6151
R831 B.n293 B.n88 10.6151
R832 B.n303 B.n88 10.6151
R833 B.n304 B.n303 10.6151
R834 B.n305 B.n304 10.6151
R835 B.n305 B.n80 10.6151
R836 B.n317 B.n80 10.6151
R837 B.n318 B.n317 10.6151
R838 B.n319 B.n318 10.6151
R839 B.n319 B.n0 10.6151
R840 B.n501 B.n1 10.6151
R841 B.n501 B.n500 10.6151
R842 B.n500 B.n499 10.6151
R843 B.n499 B.n9 10.6151
R844 B.n493 B.n9 10.6151
R845 B.n493 B.n492 10.6151
R846 B.n492 B.n491 10.6151
R847 B.n491 B.n17 10.6151
R848 B.n485 B.n17 10.6151
R849 B.n485 B.n484 10.6151
R850 B.n484 B.n483 10.6151
R851 B.n483 B.n24 10.6151
R852 B.n477 B.n24 10.6151
R853 B.n477 B.n476 10.6151
R854 B.n476 B.n475 10.6151
R855 B.n475 B.n31 10.6151
R856 B.n469 B.n31 10.6151
R857 B.n469 B.n468 10.6151
R858 B.n468 B.n467 10.6151
R859 B.n467 B.n38 10.6151
R860 B.n461 B.n38 10.6151
R861 B.n419 B.n57 9.36635
R862 B.n395 B.n65 9.36635
R863 B.n134 B.n130 9.36635
R864 B.n194 B.n193 9.36635
R865 B.t8 B.n82 6.20642
R866 B.n496 B.t3 6.20642
R867 B.n289 B.t4 4.13778
R868 B.n481 B.t5 4.13778
R869 B.n507 B.n0 2.81026
R870 B.n507 B.n1 2.81026
R871 B.n415 B.n57 1.24928
R872 B.n399 B.n65 1.24928
R873 B.n212 B.n134 1.24928
R874 B.n195 B.n194 1.24928
R875 VP.n5 VP.t8 387.197
R876 VP.n16 VP.t3 366.216
R877 VP.n17 VP.t2 366.216
R878 VP.n1 VP.t0 366.216
R879 VP.n23 VP.t9 366.216
R880 VP.n24 VP.t1 366.216
R881 VP.n13 VP.t4 366.216
R882 VP.n12 VP.t7 366.216
R883 VP.n4 VP.t6 366.216
R884 VP.n6 VP.t5 366.216
R885 VP.n25 VP.n24 161.3
R886 VP.n8 VP.n7 161.3
R887 VP.n9 VP.n4 161.3
R888 VP.n11 VP.n10 161.3
R889 VP.n12 VP.n3 161.3
R890 VP.n14 VP.n13 161.3
R891 VP.n23 VP.n0 161.3
R892 VP.n22 VP.n21 161.3
R893 VP.n20 VP.n1 161.3
R894 VP.n19 VP.n18 161.3
R895 VP.n17 VP.n2 161.3
R896 VP.n16 VP.n15 161.3
R897 VP.n8 VP.n5 70.4033
R898 VP.n17 VP.n16 48.2005
R899 VP.n24 VP.n23 48.2005
R900 VP.n13 VP.n12 48.2005
R901 VP.n18 VP.n1 39.4369
R902 VP.n22 VP.n1 39.4369
R903 VP.n11 VP.n4 39.4369
R904 VP.n7 VP.n4 39.4369
R905 VP.n15 VP.n14 36.4058
R906 VP.n6 VP.n5 20.9576
R907 VP.n18 VP.n17 8.76414
R908 VP.n23 VP.n22 8.76414
R909 VP.n12 VP.n11 8.76414
R910 VP.n7 VP.n6 8.76414
R911 VP.n9 VP.n8 0.189894
R912 VP.n10 VP.n9 0.189894
R913 VP.n10 VP.n3 0.189894
R914 VP.n14 VP.n3 0.189894
R915 VP.n15 VP.n2 0.189894
R916 VP.n19 VP.n2 0.189894
R917 VP.n20 VP.n19 0.189894
R918 VP.n21 VP.n20 0.189894
R919 VP.n21 VP.n0 0.189894
R920 VP.n25 VP.n0 0.189894
R921 VP VP.n25 0.0516364
R922 VTAIL.n120 VTAIL.n98 289.615
R923 VTAIL.n24 VTAIL.n2 289.615
R924 VTAIL.n92 VTAIL.n70 289.615
R925 VTAIL.n60 VTAIL.n38 289.615
R926 VTAIL.n106 VTAIL.n105 185
R927 VTAIL.n111 VTAIL.n110 185
R928 VTAIL.n113 VTAIL.n112 185
R929 VTAIL.n102 VTAIL.n101 185
R930 VTAIL.n119 VTAIL.n118 185
R931 VTAIL.n121 VTAIL.n120 185
R932 VTAIL.n10 VTAIL.n9 185
R933 VTAIL.n15 VTAIL.n14 185
R934 VTAIL.n17 VTAIL.n16 185
R935 VTAIL.n6 VTAIL.n5 185
R936 VTAIL.n23 VTAIL.n22 185
R937 VTAIL.n25 VTAIL.n24 185
R938 VTAIL.n93 VTAIL.n92 185
R939 VTAIL.n91 VTAIL.n90 185
R940 VTAIL.n74 VTAIL.n73 185
R941 VTAIL.n85 VTAIL.n84 185
R942 VTAIL.n83 VTAIL.n82 185
R943 VTAIL.n78 VTAIL.n77 185
R944 VTAIL.n61 VTAIL.n60 185
R945 VTAIL.n59 VTAIL.n58 185
R946 VTAIL.n42 VTAIL.n41 185
R947 VTAIL.n53 VTAIL.n52 185
R948 VTAIL.n51 VTAIL.n50 185
R949 VTAIL.n46 VTAIL.n45 185
R950 VTAIL.n107 VTAIL.t1 147.672
R951 VTAIL.n11 VTAIL.t15 147.672
R952 VTAIL.n79 VTAIL.t11 147.672
R953 VTAIL.n47 VTAIL.t5 147.672
R954 VTAIL.n111 VTAIL.n105 104.615
R955 VTAIL.n112 VTAIL.n111 104.615
R956 VTAIL.n112 VTAIL.n101 104.615
R957 VTAIL.n119 VTAIL.n101 104.615
R958 VTAIL.n120 VTAIL.n119 104.615
R959 VTAIL.n15 VTAIL.n9 104.615
R960 VTAIL.n16 VTAIL.n15 104.615
R961 VTAIL.n16 VTAIL.n5 104.615
R962 VTAIL.n23 VTAIL.n5 104.615
R963 VTAIL.n24 VTAIL.n23 104.615
R964 VTAIL.n92 VTAIL.n91 104.615
R965 VTAIL.n91 VTAIL.n73 104.615
R966 VTAIL.n84 VTAIL.n73 104.615
R967 VTAIL.n84 VTAIL.n83 104.615
R968 VTAIL.n83 VTAIL.n77 104.615
R969 VTAIL.n60 VTAIL.n59 104.615
R970 VTAIL.n59 VTAIL.n41 104.615
R971 VTAIL.n52 VTAIL.n41 104.615
R972 VTAIL.n52 VTAIL.n51 104.615
R973 VTAIL.n51 VTAIL.n45 104.615
R974 VTAIL.n69 VTAIL.n68 53.528
R975 VTAIL.n67 VTAIL.n66 53.528
R976 VTAIL.n37 VTAIL.n36 53.528
R977 VTAIL.n35 VTAIL.n34 53.528
R978 VTAIL.n127 VTAIL.n126 53.5278
R979 VTAIL.n1 VTAIL.n0 53.5278
R980 VTAIL.n31 VTAIL.n30 53.5278
R981 VTAIL.n33 VTAIL.n32 53.5278
R982 VTAIL.t1 VTAIL.n105 52.3082
R983 VTAIL.t15 VTAIL.n9 52.3082
R984 VTAIL.t11 VTAIL.n77 52.3082
R985 VTAIL.t5 VTAIL.n45 52.3082
R986 VTAIL.n125 VTAIL.n124 33.7369
R987 VTAIL.n29 VTAIL.n28 33.7369
R988 VTAIL.n97 VTAIL.n96 33.7369
R989 VTAIL.n65 VTAIL.n64 33.7369
R990 VTAIL.n35 VTAIL.n33 18.3496
R991 VTAIL.n125 VTAIL.n97 17.6686
R992 VTAIL.n107 VTAIL.n106 15.6666
R993 VTAIL.n11 VTAIL.n10 15.6666
R994 VTAIL.n79 VTAIL.n78 15.6666
R995 VTAIL.n47 VTAIL.n46 15.6666
R996 VTAIL.n110 VTAIL.n109 12.8005
R997 VTAIL.n14 VTAIL.n13 12.8005
R998 VTAIL.n82 VTAIL.n81 12.8005
R999 VTAIL.n50 VTAIL.n49 12.8005
R1000 VTAIL.n113 VTAIL.n104 12.0247
R1001 VTAIL.n17 VTAIL.n8 12.0247
R1002 VTAIL.n85 VTAIL.n76 12.0247
R1003 VTAIL.n53 VTAIL.n44 12.0247
R1004 VTAIL.n114 VTAIL.n102 11.249
R1005 VTAIL.n18 VTAIL.n6 11.249
R1006 VTAIL.n86 VTAIL.n74 11.249
R1007 VTAIL.n54 VTAIL.n42 11.249
R1008 VTAIL.n118 VTAIL.n117 10.4732
R1009 VTAIL.n22 VTAIL.n21 10.4732
R1010 VTAIL.n90 VTAIL.n89 10.4732
R1011 VTAIL.n58 VTAIL.n57 10.4732
R1012 VTAIL.n121 VTAIL.n100 9.69747
R1013 VTAIL.n25 VTAIL.n4 9.69747
R1014 VTAIL.n93 VTAIL.n72 9.69747
R1015 VTAIL.n61 VTAIL.n40 9.69747
R1016 VTAIL.n124 VTAIL.n123 9.45567
R1017 VTAIL.n28 VTAIL.n27 9.45567
R1018 VTAIL.n96 VTAIL.n95 9.45567
R1019 VTAIL.n64 VTAIL.n63 9.45567
R1020 VTAIL.n123 VTAIL.n122 9.3005
R1021 VTAIL.n100 VTAIL.n99 9.3005
R1022 VTAIL.n117 VTAIL.n116 9.3005
R1023 VTAIL.n115 VTAIL.n114 9.3005
R1024 VTAIL.n104 VTAIL.n103 9.3005
R1025 VTAIL.n109 VTAIL.n108 9.3005
R1026 VTAIL.n27 VTAIL.n26 9.3005
R1027 VTAIL.n4 VTAIL.n3 9.3005
R1028 VTAIL.n21 VTAIL.n20 9.3005
R1029 VTAIL.n19 VTAIL.n18 9.3005
R1030 VTAIL.n8 VTAIL.n7 9.3005
R1031 VTAIL.n13 VTAIL.n12 9.3005
R1032 VTAIL.n95 VTAIL.n94 9.3005
R1033 VTAIL.n72 VTAIL.n71 9.3005
R1034 VTAIL.n89 VTAIL.n88 9.3005
R1035 VTAIL.n87 VTAIL.n86 9.3005
R1036 VTAIL.n76 VTAIL.n75 9.3005
R1037 VTAIL.n81 VTAIL.n80 9.3005
R1038 VTAIL.n63 VTAIL.n62 9.3005
R1039 VTAIL.n40 VTAIL.n39 9.3005
R1040 VTAIL.n57 VTAIL.n56 9.3005
R1041 VTAIL.n55 VTAIL.n54 9.3005
R1042 VTAIL.n44 VTAIL.n43 9.3005
R1043 VTAIL.n49 VTAIL.n48 9.3005
R1044 VTAIL.n122 VTAIL.n98 8.92171
R1045 VTAIL.n26 VTAIL.n2 8.92171
R1046 VTAIL.n94 VTAIL.n70 8.92171
R1047 VTAIL.n62 VTAIL.n38 8.92171
R1048 VTAIL.n124 VTAIL.n98 5.04292
R1049 VTAIL.n28 VTAIL.n2 5.04292
R1050 VTAIL.n96 VTAIL.n70 5.04292
R1051 VTAIL.n64 VTAIL.n38 5.04292
R1052 VTAIL.n108 VTAIL.n107 4.38687
R1053 VTAIL.n12 VTAIL.n11 4.38687
R1054 VTAIL.n80 VTAIL.n79 4.38687
R1055 VTAIL.n48 VTAIL.n47 4.38687
R1056 VTAIL.n122 VTAIL.n121 4.26717
R1057 VTAIL.n26 VTAIL.n25 4.26717
R1058 VTAIL.n94 VTAIL.n93 4.26717
R1059 VTAIL.n62 VTAIL.n61 4.26717
R1060 VTAIL.n126 VTAIL.t16 3.69453
R1061 VTAIL.n126 VTAIL.t19 3.69453
R1062 VTAIL.n0 VTAIL.t17 3.69453
R1063 VTAIL.n0 VTAIL.t18 3.69453
R1064 VTAIL.n30 VTAIL.t13 3.69453
R1065 VTAIL.n30 VTAIL.t8 3.69453
R1066 VTAIL.n32 VTAIL.t10 3.69453
R1067 VTAIL.n32 VTAIL.t14 3.69453
R1068 VTAIL.n68 VTAIL.t9 3.69453
R1069 VTAIL.n68 VTAIL.t7 3.69453
R1070 VTAIL.n66 VTAIL.t6 3.69453
R1071 VTAIL.n66 VTAIL.t12 3.69453
R1072 VTAIL.n36 VTAIL.t4 3.69453
R1073 VTAIL.n36 VTAIL.t3 3.69453
R1074 VTAIL.n34 VTAIL.t0 3.69453
R1075 VTAIL.n34 VTAIL.t2 3.69453
R1076 VTAIL.n118 VTAIL.n100 3.49141
R1077 VTAIL.n22 VTAIL.n4 3.49141
R1078 VTAIL.n90 VTAIL.n72 3.49141
R1079 VTAIL.n58 VTAIL.n40 3.49141
R1080 VTAIL.n117 VTAIL.n102 2.71565
R1081 VTAIL.n21 VTAIL.n6 2.71565
R1082 VTAIL.n89 VTAIL.n74 2.71565
R1083 VTAIL.n57 VTAIL.n42 2.71565
R1084 VTAIL.n114 VTAIL.n113 1.93989
R1085 VTAIL.n18 VTAIL.n17 1.93989
R1086 VTAIL.n86 VTAIL.n85 1.93989
R1087 VTAIL.n54 VTAIL.n53 1.93989
R1088 VTAIL.n110 VTAIL.n104 1.16414
R1089 VTAIL.n14 VTAIL.n8 1.16414
R1090 VTAIL.n82 VTAIL.n76 1.16414
R1091 VTAIL.n50 VTAIL.n44 1.16414
R1092 VTAIL.n67 VTAIL.n65 0.810845
R1093 VTAIL.n29 VTAIL.n1 0.810845
R1094 VTAIL.n37 VTAIL.n35 0.681535
R1095 VTAIL.n65 VTAIL.n37 0.681535
R1096 VTAIL.n69 VTAIL.n67 0.681535
R1097 VTAIL.n97 VTAIL.n69 0.681535
R1098 VTAIL.n33 VTAIL.n31 0.681535
R1099 VTAIL.n31 VTAIL.n29 0.681535
R1100 VTAIL.n127 VTAIL.n125 0.681535
R1101 VTAIL VTAIL.n1 0.569465
R1102 VTAIL.n109 VTAIL.n106 0.388379
R1103 VTAIL.n13 VTAIL.n10 0.388379
R1104 VTAIL.n81 VTAIL.n78 0.388379
R1105 VTAIL.n49 VTAIL.n46 0.388379
R1106 VTAIL.n108 VTAIL.n103 0.155672
R1107 VTAIL.n115 VTAIL.n103 0.155672
R1108 VTAIL.n116 VTAIL.n115 0.155672
R1109 VTAIL.n116 VTAIL.n99 0.155672
R1110 VTAIL.n123 VTAIL.n99 0.155672
R1111 VTAIL.n12 VTAIL.n7 0.155672
R1112 VTAIL.n19 VTAIL.n7 0.155672
R1113 VTAIL.n20 VTAIL.n19 0.155672
R1114 VTAIL.n20 VTAIL.n3 0.155672
R1115 VTAIL.n27 VTAIL.n3 0.155672
R1116 VTAIL.n95 VTAIL.n71 0.155672
R1117 VTAIL.n88 VTAIL.n71 0.155672
R1118 VTAIL.n88 VTAIL.n87 0.155672
R1119 VTAIL.n87 VTAIL.n75 0.155672
R1120 VTAIL.n80 VTAIL.n75 0.155672
R1121 VTAIL.n63 VTAIL.n39 0.155672
R1122 VTAIL.n56 VTAIL.n39 0.155672
R1123 VTAIL.n56 VTAIL.n55 0.155672
R1124 VTAIL.n55 VTAIL.n43 0.155672
R1125 VTAIL.n48 VTAIL.n43 0.155672
R1126 VTAIL VTAIL.n127 0.112569
R1127 VDD1.n22 VDD1.n0 289.615
R1128 VDD1.n51 VDD1.n29 289.615
R1129 VDD1.n23 VDD1.n22 185
R1130 VDD1.n21 VDD1.n20 185
R1131 VDD1.n4 VDD1.n3 185
R1132 VDD1.n15 VDD1.n14 185
R1133 VDD1.n13 VDD1.n12 185
R1134 VDD1.n8 VDD1.n7 185
R1135 VDD1.n37 VDD1.n36 185
R1136 VDD1.n42 VDD1.n41 185
R1137 VDD1.n44 VDD1.n43 185
R1138 VDD1.n33 VDD1.n32 185
R1139 VDD1.n50 VDD1.n49 185
R1140 VDD1.n52 VDD1.n51 185
R1141 VDD1.n9 VDD1.t1 147.672
R1142 VDD1.n38 VDD1.t6 147.672
R1143 VDD1.n22 VDD1.n21 104.615
R1144 VDD1.n21 VDD1.n3 104.615
R1145 VDD1.n14 VDD1.n3 104.615
R1146 VDD1.n14 VDD1.n13 104.615
R1147 VDD1.n13 VDD1.n7 104.615
R1148 VDD1.n42 VDD1.n36 104.615
R1149 VDD1.n43 VDD1.n42 104.615
R1150 VDD1.n43 VDD1.n32 104.615
R1151 VDD1.n50 VDD1.n32 104.615
R1152 VDD1.n51 VDD1.n50 104.615
R1153 VDD1.n59 VDD1.n58 70.6621
R1154 VDD1.n28 VDD1.n27 70.2068
R1155 VDD1.n61 VDD1.n60 70.2066
R1156 VDD1.n57 VDD1.n56 70.2066
R1157 VDD1.t1 VDD1.n7 52.3082
R1158 VDD1.t6 VDD1.n36 52.3082
R1159 VDD1.n28 VDD1.n26 51.0967
R1160 VDD1.n57 VDD1.n55 51.0967
R1161 VDD1.n61 VDD1.n59 32.4944
R1162 VDD1.n9 VDD1.n8 15.6666
R1163 VDD1.n38 VDD1.n37 15.6666
R1164 VDD1.n12 VDD1.n11 12.8005
R1165 VDD1.n41 VDD1.n40 12.8005
R1166 VDD1.n15 VDD1.n6 12.0247
R1167 VDD1.n44 VDD1.n35 12.0247
R1168 VDD1.n16 VDD1.n4 11.249
R1169 VDD1.n45 VDD1.n33 11.249
R1170 VDD1.n20 VDD1.n19 10.4732
R1171 VDD1.n49 VDD1.n48 10.4732
R1172 VDD1.n23 VDD1.n2 9.69747
R1173 VDD1.n52 VDD1.n31 9.69747
R1174 VDD1.n26 VDD1.n25 9.45567
R1175 VDD1.n55 VDD1.n54 9.45567
R1176 VDD1.n25 VDD1.n24 9.3005
R1177 VDD1.n2 VDD1.n1 9.3005
R1178 VDD1.n19 VDD1.n18 9.3005
R1179 VDD1.n17 VDD1.n16 9.3005
R1180 VDD1.n6 VDD1.n5 9.3005
R1181 VDD1.n11 VDD1.n10 9.3005
R1182 VDD1.n54 VDD1.n53 9.3005
R1183 VDD1.n31 VDD1.n30 9.3005
R1184 VDD1.n48 VDD1.n47 9.3005
R1185 VDD1.n46 VDD1.n45 9.3005
R1186 VDD1.n35 VDD1.n34 9.3005
R1187 VDD1.n40 VDD1.n39 9.3005
R1188 VDD1.n24 VDD1.n0 8.92171
R1189 VDD1.n53 VDD1.n29 8.92171
R1190 VDD1.n26 VDD1.n0 5.04292
R1191 VDD1.n55 VDD1.n29 5.04292
R1192 VDD1.n10 VDD1.n9 4.38687
R1193 VDD1.n39 VDD1.n38 4.38687
R1194 VDD1.n24 VDD1.n23 4.26717
R1195 VDD1.n53 VDD1.n52 4.26717
R1196 VDD1.n60 VDD1.t2 3.69453
R1197 VDD1.n60 VDD1.t5 3.69453
R1198 VDD1.n27 VDD1.t4 3.69453
R1199 VDD1.n27 VDD1.t3 3.69453
R1200 VDD1.n58 VDD1.t0 3.69453
R1201 VDD1.n58 VDD1.t8 3.69453
R1202 VDD1.n56 VDD1.t7 3.69453
R1203 VDD1.n56 VDD1.t9 3.69453
R1204 VDD1.n20 VDD1.n2 3.49141
R1205 VDD1.n49 VDD1.n31 3.49141
R1206 VDD1.n19 VDD1.n4 2.71565
R1207 VDD1.n48 VDD1.n33 2.71565
R1208 VDD1.n16 VDD1.n15 1.93989
R1209 VDD1.n45 VDD1.n44 1.93989
R1210 VDD1.n12 VDD1.n6 1.16414
R1211 VDD1.n41 VDD1.n35 1.16414
R1212 VDD1 VDD1.n61 0.453086
R1213 VDD1.n11 VDD1.n8 0.388379
R1214 VDD1.n40 VDD1.n37 0.388379
R1215 VDD1 VDD1.n28 0.228948
R1216 VDD1.n25 VDD1.n1 0.155672
R1217 VDD1.n18 VDD1.n1 0.155672
R1218 VDD1.n18 VDD1.n17 0.155672
R1219 VDD1.n17 VDD1.n5 0.155672
R1220 VDD1.n10 VDD1.n5 0.155672
R1221 VDD1.n39 VDD1.n34 0.155672
R1222 VDD1.n46 VDD1.n34 0.155672
R1223 VDD1.n47 VDD1.n46 0.155672
R1224 VDD1.n47 VDD1.n30 0.155672
R1225 VDD1.n54 VDD1.n30 0.155672
R1226 VDD1.n59 VDD1.n57 0.115413
R1227 VN.n2 VN.t0 387.197
R1228 VN.n14 VN.t7 387.197
R1229 VN.n3 VN.t1 366.216
R1230 VN.n1 VN.t9 366.216
R1231 VN.n9 VN.t2 366.216
R1232 VN.n10 VN.t3 366.216
R1233 VN.n15 VN.t8 366.216
R1234 VN.n13 VN.t5 366.216
R1235 VN.n21 VN.t6 366.216
R1236 VN.n22 VN.t4 366.216
R1237 VN.n11 VN.n10 161.3
R1238 VN.n23 VN.n22 161.3
R1239 VN.n21 VN.n12 161.3
R1240 VN.n20 VN.n19 161.3
R1241 VN.n18 VN.n13 161.3
R1242 VN.n17 VN.n16 161.3
R1243 VN.n9 VN.n0 161.3
R1244 VN.n8 VN.n7 161.3
R1245 VN.n6 VN.n1 161.3
R1246 VN.n5 VN.n4 161.3
R1247 VN.n17 VN.n14 70.4033
R1248 VN.n5 VN.n2 70.4033
R1249 VN.n10 VN.n9 48.2005
R1250 VN.n22 VN.n21 48.2005
R1251 VN.n4 VN.n1 39.4369
R1252 VN.n8 VN.n1 39.4369
R1253 VN.n16 VN.n13 39.4369
R1254 VN.n20 VN.n13 39.4369
R1255 VN VN.n23 36.7865
R1256 VN.n15 VN.n14 20.9576
R1257 VN.n3 VN.n2 20.9576
R1258 VN.n4 VN.n3 8.76414
R1259 VN.n9 VN.n8 8.76414
R1260 VN.n16 VN.n15 8.76414
R1261 VN.n21 VN.n20 8.76414
R1262 VN.n23 VN.n12 0.189894
R1263 VN.n19 VN.n12 0.189894
R1264 VN.n19 VN.n18 0.189894
R1265 VN.n18 VN.n17 0.189894
R1266 VN.n6 VN.n5 0.189894
R1267 VN.n7 VN.n6 0.189894
R1268 VN.n7 VN.n0 0.189894
R1269 VN.n11 VN.n0 0.189894
R1270 VN VN.n11 0.0516364
R1271 VDD2.n53 VDD2.n31 289.615
R1272 VDD2.n22 VDD2.n0 289.615
R1273 VDD2.n54 VDD2.n53 185
R1274 VDD2.n52 VDD2.n51 185
R1275 VDD2.n35 VDD2.n34 185
R1276 VDD2.n46 VDD2.n45 185
R1277 VDD2.n44 VDD2.n43 185
R1278 VDD2.n39 VDD2.n38 185
R1279 VDD2.n8 VDD2.n7 185
R1280 VDD2.n13 VDD2.n12 185
R1281 VDD2.n15 VDD2.n14 185
R1282 VDD2.n4 VDD2.n3 185
R1283 VDD2.n21 VDD2.n20 185
R1284 VDD2.n23 VDD2.n22 185
R1285 VDD2.n40 VDD2.t5 147.672
R1286 VDD2.n9 VDD2.t9 147.672
R1287 VDD2.n53 VDD2.n52 104.615
R1288 VDD2.n52 VDD2.n34 104.615
R1289 VDD2.n45 VDD2.n34 104.615
R1290 VDD2.n45 VDD2.n44 104.615
R1291 VDD2.n44 VDD2.n38 104.615
R1292 VDD2.n13 VDD2.n7 104.615
R1293 VDD2.n14 VDD2.n13 104.615
R1294 VDD2.n14 VDD2.n3 104.615
R1295 VDD2.n21 VDD2.n3 104.615
R1296 VDD2.n22 VDD2.n21 104.615
R1297 VDD2.n30 VDD2.n29 70.6621
R1298 VDD2 VDD2.n61 70.6592
R1299 VDD2.n60 VDD2.n59 70.2068
R1300 VDD2.n28 VDD2.n27 70.2066
R1301 VDD2.t5 VDD2.n38 52.3082
R1302 VDD2.t9 VDD2.n7 52.3082
R1303 VDD2.n28 VDD2.n26 51.0967
R1304 VDD2.n58 VDD2.n57 50.4157
R1305 VDD2.n58 VDD2.n30 31.5709
R1306 VDD2.n40 VDD2.n39 15.6666
R1307 VDD2.n9 VDD2.n8 15.6666
R1308 VDD2.n43 VDD2.n42 12.8005
R1309 VDD2.n12 VDD2.n11 12.8005
R1310 VDD2.n46 VDD2.n37 12.0247
R1311 VDD2.n15 VDD2.n6 12.0247
R1312 VDD2.n47 VDD2.n35 11.249
R1313 VDD2.n16 VDD2.n4 11.249
R1314 VDD2.n51 VDD2.n50 10.4732
R1315 VDD2.n20 VDD2.n19 10.4732
R1316 VDD2.n54 VDD2.n33 9.69747
R1317 VDD2.n23 VDD2.n2 9.69747
R1318 VDD2.n57 VDD2.n56 9.45567
R1319 VDD2.n26 VDD2.n25 9.45567
R1320 VDD2.n56 VDD2.n55 9.3005
R1321 VDD2.n33 VDD2.n32 9.3005
R1322 VDD2.n50 VDD2.n49 9.3005
R1323 VDD2.n48 VDD2.n47 9.3005
R1324 VDD2.n37 VDD2.n36 9.3005
R1325 VDD2.n42 VDD2.n41 9.3005
R1326 VDD2.n25 VDD2.n24 9.3005
R1327 VDD2.n2 VDD2.n1 9.3005
R1328 VDD2.n19 VDD2.n18 9.3005
R1329 VDD2.n17 VDD2.n16 9.3005
R1330 VDD2.n6 VDD2.n5 9.3005
R1331 VDD2.n11 VDD2.n10 9.3005
R1332 VDD2.n55 VDD2.n31 8.92171
R1333 VDD2.n24 VDD2.n0 8.92171
R1334 VDD2.n57 VDD2.n31 5.04292
R1335 VDD2.n26 VDD2.n0 5.04292
R1336 VDD2.n41 VDD2.n40 4.38687
R1337 VDD2.n10 VDD2.n9 4.38687
R1338 VDD2.n55 VDD2.n54 4.26717
R1339 VDD2.n24 VDD2.n23 4.26717
R1340 VDD2.n61 VDD2.t1 3.69453
R1341 VDD2.n61 VDD2.t2 3.69453
R1342 VDD2.n59 VDD2.t3 3.69453
R1343 VDD2.n59 VDD2.t4 3.69453
R1344 VDD2.n29 VDD2.t7 3.69453
R1345 VDD2.n29 VDD2.t6 3.69453
R1346 VDD2.n27 VDD2.t8 3.69453
R1347 VDD2.n27 VDD2.t0 3.69453
R1348 VDD2.n51 VDD2.n33 3.49141
R1349 VDD2.n20 VDD2.n2 3.49141
R1350 VDD2.n50 VDD2.n35 2.71565
R1351 VDD2.n19 VDD2.n4 2.71565
R1352 VDD2.n47 VDD2.n46 1.93989
R1353 VDD2.n16 VDD2.n15 1.93989
R1354 VDD2.n43 VDD2.n37 1.16414
R1355 VDD2.n12 VDD2.n6 1.16414
R1356 VDD2.n60 VDD2.n58 0.681535
R1357 VDD2.n42 VDD2.n39 0.388379
R1358 VDD2.n11 VDD2.n8 0.388379
R1359 VDD2 VDD2.n60 0.228948
R1360 VDD2.n56 VDD2.n32 0.155672
R1361 VDD2.n49 VDD2.n32 0.155672
R1362 VDD2.n49 VDD2.n48 0.155672
R1363 VDD2.n48 VDD2.n36 0.155672
R1364 VDD2.n41 VDD2.n36 0.155672
R1365 VDD2.n10 VDD2.n5 0.155672
R1366 VDD2.n17 VDD2.n5 0.155672
R1367 VDD2.n18 VDD2.n17 0.155672
R1368 VDD2.n18 VDD2.n1 0.155672
R1369 VDD2.n25 VDD2.n1 0.155672
R1370 VDD2.n30 VDD2.n28 0.115413
C0 VP VDD1 2.72939f
C1 VDD2 VDD1 0.821494f
C2 VP VDD2 0.314228f
C3 VDD1 VTAIL 8.927019f
C4 VP VTAIL 2.6154f
C5 VDD2 VTAIL 8.962799f
C6 VDD1 VN 0.14881f
C7 VP VN 4.01467f
C8 VDD2 VN 2.57037f
C9 VTAIL VN 2.60103f
C10 VDD2 B 3.510956f
C11 VDD1 B 3.415347f
C12 VTAIL B 3.776351f
C13 VN B 7.548049f
C14 VP B 5.817993f
C15 VDD2.n0 B 0.038156f
C16 VDD2.n1 B 0.026635f
C17 VDD2.n2 B 0.014312f
C18 VDD2.n3 B 0.033829f
C19 VDD2.n4 B 0.015154f
C20 VDD2.n5 B 0.026635f
C21 VDD2.n6 B 0.014312f
C22 VDD2.n7 B 0.025372f
C23 VDD2.n8 B 0.019979f
C24 VDD2.t9 B 0.055288f
C25 VDD2.n9 B 0.110111f
C26 VDD2.n10 B 0.555013f
C27 VDD2.n11 B 0.014312f
C28 VDD2.n12 B 0.015154f
C29 VDD2.n13 B 0.033829f
C30 VDD2.n14 B 0.033829f
C31 VDD2.n15 B 0.015154f
C32 VDD2.n16 B 0.014312f
C33 VDD2.n17 B 0.026635f
C34 VDD2.n18 B 0.026635f
C35 VDD2.n19 B 0.014312f
C36 VDD2.n20 B 0.015154f
C37 VDD2.n21 B 0.033829f
C38 VDD2.n22 B 0.074506f
C39 VDD2.n23 B 0.015154f
C40 VDD2.n24 B 0.014312f
C41 VDD2.n25 B 0.064476f
C42 VDD2.n26 B 0.061761f
C43 VDD2.t8 B 0.112815f
C44 VDD2.t0 B 0.112815f
C45 VDD2.n27 B 0.927719f
C46 VDD2.n28 B 0.39711f
C47 VDD2.t7 B 0.112815f
C48 VDD2.t6 B 0.112815f
C49 VDD2.n29 B 0.929801f
C50 VDD2.n30 B 1.46647f
C51 VDD2.n31 B 0.038156f
C52 VDD2.n32 B 0.026635f
C53 VDD2.n33 B 0.014312f
C54 VDD2.n34 B 0.033829f
C55 VDD2.n35 B 0.015154f
C56 VDD2.n36 B 0.026635f
C57 VDD2.n37 B 0.014312f
C58 VDD2.n38 B 0.025372f
C59 VDD2.n39 B 0.019979f
C60 VDD2.t5 B 0.055288f
C61 VDD2.n40 B 0.110111f
C62 VDD2.n41 B 0.555013f
C63 VDD2.n42 B 0.014312f
C64 VDD2.n43 B 0.015154f
C65 VDD2.n44 B 0.033829f
C66 VDD2.n45 B 0.033829f
C67 VDD2.n46 B 0.015154f
C68 VDD2.n47 B 0.014312f
C69 VDD2.n48 B 0.026635f
C70 VDD2.n49 B 0.026635f
C71 VDD2.n50 B 0.014312f
C72 VDD2.n51 B 0.015154f
C73 VDD2.n52 B 0.033829f
C74 VDD2.n53 B 0.074506f
C75 VDD2.n54 B 0.015154f
C76 VDD2.n55 B 0.014312f
C77 VDD2.n56 B 0.064476f
C78 VDD2.n57 B 0.060276f
C79 VDD2.n58 B 1.63456f
C80 VDD2.t3 B 0.112815f
C81 VDD2.t4 B 0.112815f
C82 VDD2.n59 B 0.927723f
C83 VDD2.n60 B 0.291558f
C84 VDD2.t1 B 0.112815f
C85 VDD2.t2 B 0.112815f
C86 VDD2.n61 B 0.929779f
C87 VN.n0 B 0.049194f
C88 VN.t9 B 0.353238f
C89 VN.n1 B 0.179248f
C90 VN.t0 B 0.36261f
C91 VN.n2 B 0.163844f
C92 VN.t1 B 0.353238f
C93 VN.n3 B 0.174699f
C94 VN.n4 B 0.011163f
C95 VN.n5 B 0.150886f
C96 VN.n6 B 0.049194f
C97 VN.n7 B 0.049194f
C98 VN.n8 B 0.011163f
C99 VN.t2 B 0.353238f
C100 VN.n9 B 0.174699f
C101 VN.t3 B 0.353238f
C102 VN.n10 B 0.172879f
C103 VN.n11 B 0.038124f
C104 VN.n12 B 0.049194f
C105 VN.t5 B 0.353238f
C106 VN.n13 B 0.179248f
C107 VN.t7 B 0.36261f
C108 VN.n14 B 0.163844f
C109 VN.t8 B 0.353238f
C110 VN.n15 B 0.174699f
C111 VN.n16 B 0.011163f
C112 VN.n17 B 0.150886f
C113 VN.n18 B 0.049194f
C114 VN.n19 B 0.049194f
C115 VN.n20 B 0.011163f
C116 VN.t6 B 0.353238f
C117 VN.n21 B 0.174699f
C118 VN.t4 B 0.353238f
C119 VN.n22 B 0.172879f
C120 VN.n23 B 1.61194f
C121 VDD1.n0 B 0.037836f
C122 VDD1.n1 B 0.026411f
C123 VDD1.n2 B 0.014192f
C124 VDD1.n3 B 0.033545f
C125 VDD1.n4 B 0.015027f
C126 VDD1.n5 B 0.026411f
C127 VDD1.n6 B 0.014192f
C128 VDD1.n7 B 0.025159f
C129 VDD1.n8 B 0.019811f
C130 VDD1.t1 B 0.054823f
C131 VDD1.n9 B 0.109185f
C132 VDD1.n10 B 0.550346f
C133 VDD1.n11 B 0.014192f
C134 VDD1.n12 B 0.015027f
C135 VDD1.n13 B 0.033545f
C136 VDD1.n14 B 0.033545f
C137 VDD1.n15 B 0.015027f
C138 VDD1.n16 B 0.014192f
C139 VDD1.n17 B 0.026411f
C140 VDD1.n18 B 0.026411f
C141 VDD1.n19 B 0.014192f
C142 VDD1.n20 B 0.015027f
C143 VDD1.n21 B 0.033545f
C144 VDD1.n22 B 0.073879f
C145 VDD1.n23 B 0.015027f
C146 VDD1.n24 B 0.014192f
C147 VDD1.n25 B 0.063934f
C148 VDD1.n26 B 0.061241f
C149 VDD1.t4 B 0.111866f
C150 VDD1.t3 B 0.111866f
C151 VDD1.n27 B 0.919922f
C152 VDD1.n28 B 0.3981f
C153 VDD1.n29 B 0.037836f
C154 VDD1.n30 B 0.026411f
C155 VDD1.n31 B 0.014192f
C156 VDD1.n32 B 0.033545f
C157 VDD1.n33 B 0.015027f
C158 VDD1.n34 B 0.026411f
C159 VDD1.n35 B 0.014192f
C160 VDD1.n36 B 0.025159f
C161 VDD1.n37 B 0.019811f
C162 VDD1.t6 B 0.054823f
C163 VDD1.n38 B 0.109185f
C164 VDD1.n39 B 0.550346f
C165 VDD1.n40 B 0.014192f
C166 VDD1.n41 B 0.015027f
C167 VDD1.n42 B 0.033545f
C168 VDD1.n43 B 0.033545f
C169 VDD1.n44 B 0.015027f
C170 VDD1.n45 B 0.014192f
C171 VDD1.n46 B 0.026411f
C172 VDD1.n47 B 0.026411f
C173 VDD1.n48 B 0.014192f
C174 VDD1.n49 B 0.015027f
C175 VDD1.n50 B 0.033545f
C176 VDD1.n51 B 0.073879f
C177 VDD1.n52 B 0.015027f
C178 VDD1.n53 B 0.014192f
C179 VDD1.n54 B 0.063934f
C180 VDD1.n55 B 0.061241f
C181 VDD1.t7 B 0.111866f
C182 VDD1.t9 B 0.111866f
C183 VDD1.n56 B 0.919917f
C184 VDD1.n57 B 0.39377f
C185 VDD1.t0 B 0.111866f
C186 VDD1.t8 B 0.111866f
C187 VDD1.n58 B 0.921982f
C188 VDD1.n59 B 1.5273f
C189 VDD1.t2 B 0.111866f
C190 VDD1.t5 B 0.111866f
C191 VDD1.n60 B 0.919917f
C192 VDD1.n61 B 1.85356f
C193 VTAIL.t17 B 0.124729f
C194 VTAIL.t18 B 0.124729f
C195 VTAIL.n0 B 0.953883f
C196 VTAIL.n1 B 0.398714f
C197 VTAIL.n2 B 0.042186f
C198 VTAIL.n3 B 0.029448f
C199 VTAIL.n4 B 0.015824f
C200 VTAIL.n5 B 0.037402f
C201 VTAIL.n6 B 0.016755f
C202 VTAIL.n7 B 0.029448f
C203 VTAIL.n8 B 0.015824f
C204 VTAIL.n9 B 0.028051f
C205 VTAIL.n10 B 0.022089f
C206 VTAIL.t15 B 0.061127f
C207 VTAIL.n11 B 0.121739f
C208 VTAIL.n12 B 0.613624f
C209 VTAIL.n13 B 0.015824f
C210 VTAIL.n14 B 0.016755f
C211 VTAIL.n15 B 0.037402f
C212 VTAIL.n16 B 0.037402f
C213 VTAIL.n17 B 0.016755f
C214 VTAIL.n18 B 0.015824f
C215 VTAIL.n19 B 0.029448f
C216 VTAIL.n20 B 0.029448f
C217 VTAIL.n21 B 0.015824f
C218 VTAIL.n22 B 0.016755f
C219 VTAIL.n23 B 0.037402f
C220 VTAIL.n24 B 0.082374f
C221 VTAIL.n25 B 0.016755f
C222 VTAIL.n26 B 0.015824f
C223 VTAIL.n27 B 0.071285f
C224 VTAIL.n28 B 0.046333f
C225 VTAIL.n29 B 0.16848f
C226 VTAIL.t13 B 0.124729f
C227 VTAIL.t8 B 0.124729f
C228 VTAIL.n30 B 0.953883f
C229 VTAIL.n31 B 0.397078f
C230 VTAIL.t10 B 0.124729f
C231 VTAIL.t14 B 0.124729f
C232 VTAIL.n32 B 0.953883f
C233 VTAIL.n33 B 1.30015f
C234 VTAIL.t0 B 0.124729f
C235 VTAIL.t2 B 0.124729f
C236 VTAIL.n34 B 0.95389f
C237 VTAIL.n35 B 1.30014f
C238 VTAIL.t4 B 0.124729f
C239 VTAIL.t3 B 0.124729f
C240 VTAIL.n36 B 0.95389f
C241 VTAIL.n37 B 0.397072f
C242 VTAIL.n38 B 0.042186f
C243 VTAIL.n39 B 0.029448f
C244 VTAIL.n40 B 0.015824f
C245 VTAIL.n41 B 0.037402f
C246 VTAIL.n42 B 0.016755f
C247 VTAIL.n43 B 0.029448f
C248 VTAIL.n44 B 0.015824f
C249 VTAIL.n45 B 0.028051f
C250 VTAIL.n46 B 0.022089f
C251 VTAIL.t5 B 0.061127f
C252 VTAIL.n47 B 0.121739f
C253 VTAIL.n48 B 0.613624f
C254 VTAIL.n49 B 0.015824f
C255 VTAIL.n50 B 0.016755f
C256 VTAIL.n51 B 0.037402f
C257 VTAIL.n52 B 0.037402f
C258 VTAIL.n53 B 0.016755f
C259 VTAIL.n54 B 0.015824f
C260 VTAIL.n55 B 0.029448f
C261 VTAIL.n56 B 0.029448f
C262 VTAIL.n57 B 0.015824f
C263 VTAIL.n58 B 0.016755f
C264 VTAIL.n59 B 0.037402f
C265 VTAIL.n60 B 0.082374f
C266 VTAIL.n61 B 0.016755f
C267 VTAIL.n62 B 0.015824f
C268 VTAIL.n63 B 0.071285f
C269 VTAIL.n64 B 0.046333f
C270 VTAIL.n65 B 0.16848f
C271 VTAIL.t6 B 0.124729f
C272 VTAIL.t12 B 0.124729f
C273 VTAIL.n66 B 0.95389f
C274 VTAIL.n67 B 0.409342f
C275 VTAIL.t9 B 0.124729f
C276 VTAIL.t7 B 0.124729f
C277 VTAIL.n68 B 0.95389f
C278 VTAIL.n69 B 0.397072f
C279 VTAIL.n70 B 0.042186f
C280 VTAIL.n71 B 0.029448f
C281 VTAIL.n72 B 0.015824f
C282 VTAIL.n73 B 0.037402f
C283 VTAIL.n74 B 0.016755f
C284 VTAIL.n75 B 0.029448f
C285 VTAIL.n76 B 0.015824f
C286 VTAIL.n77 B 0.028051f
C287 VTAIL.n78 B 0.022089f
C288 VTAIL.t11 B 0.061127f
C289 VTAIL.n79 B 0.121739f
C290 VTAIL.n80 B 0.613624f
C291 VTAIL.n81 B 0.015824f
C292 VTAIL.n82 B 0.016755f
C293 VTAIL.n83 B 0.037402f
C294 VTAIL.n84 B 0.037402f
C295 VTAIL.n85 B 0.016755f
C296 VTAIL.n86 B 0.015824f
C297 VTAIL.n87 B 0.029448f
C298 VTAIL.n88 B 0.029448f
C299 VTAIL.n89 B 0.015824f
C300 VTAIL.n90 B 0.016755f
C301 VTAIL.n91 B 0.037402f
C302 VTAIL.n92 B 0.082374f
C303 VTAIL.n93 B 0.016755f
C304 VTAIL.n94 B 0.015824f
C305 VTAIL.n95 B 0.071285f
C306 VTAIL.n96 B 0.046333f
C307 VTAIL.n97 B 0.994661f
C308 VTAIL.n98 B 0.042186f
C309 VTAIL.n99 B 0.029448f
C310 VTAIL.n100 B 0.015824f
C311 VTAIL.n101 B 0.037402f
C312 VTAIL.n102 B 0.016755f
C313 VTAIL.n103 B 0.029448f
C314 VTAIL.n104 B 0.015824f
C315 VTAIL.n105 B 0.028051f
C316 VTAIL.n106 B 0.022089f
C317 VTAIL.t1 B 0.061127f
C318 VTAIL.n107 B 0.121739f
C319 VTAIL.n108 B 0.613624f
C320 VTAIL.n109 B 0.015824f
C321 VTAIL.n110 B 0.016755f
C322 VTAIL.n111 B 0.037402f
C323 VTAIL.n112 B 0.037402f
C324 VTAIL.n113 B 0.016755f
C325 VTAIL.n114 B 0.015824f
C326 VTAIL.n115 B 0.029448f
C327 VTAIL.n116 B 0.029448f
C328 VTAIL.n117 B 0.015824f
C329 VTAIL.n118 B 0.016755f
C330 VTAIL.n119 B 0.037402f
C331 VTAIL.n120 B 0.082374f
C332 VTAIL.n121 B 0.016755f
C333 VTAIL.n122 B 0.015824f
C334 VTAIL.n123 B 0.071285f
C335 VTAIL.n124 B 0.046333f
C336 VTAIL.n125 B 0.994661f
C337 VTAIL.t16 B 0.124729f
C338 VTAIL.t19 B 0.124729f
C339 VTAIL.n126 B 0.953883f
C340 VTAIL.n127 B 0.343091f
C341 VP.n0 B 0.050106f
C342 VP.t0 B 0.359782f
C343 VP.n1 B 0.182569f
C344 VP.n2 B 0.050106f
C345 VP.n3 B 0.050106f
C346 VP.t4 B 0.359782f
C347 VP.t7 B 0.359782f
C348 VP.t6 B 0.359782f
C349 VP.n4 B 0.182569f
C350 VP.t8 B 0.369327f
C351 VP.n5 B 0.166879f
C352 VP.t5 B 0.359782f
C353 VP.n6 B 0.177935f
C354 VP.n7 B 0.01137f
C355 VP.n8 B 0.153681f
C356 VP.n9 B 0.050106f
C357 VP.n10 B 0.050106f
C358 VP.n11 B 0.01137f
C359 VP.n12 B 0.177935f
C360 VP.n13 B 0.176082f
C361 VP.n14 B 1.6086f
C362 VP.n15 B 1.65821f
C363 VP.t3 B 0.359782f
C364 VP.n16 B 0.176082f
C365 VP.t2 B 0.359782f
C366 VP.n17 B 0.177935f
C367 VP.n18 B 0.01137f
C368 VP.n19 B 0.050106f
C369 VP.n20 B 0.050106f
C370 VP.n21 B 0.050106f
C371 VP.n22 B 0.01137f
C372 VP.t9 B 0.359782f
C373 VP.n23 B 0.177935f
C374 VP.t1 B 0.359782f
C375 VP.n24 B 0.176082f
C376 VP.n25 B 0.03883f
.ends

