* NGSPICE file created from diff_pair_sample_0336.ext - technology: sky130A

.subckt diff_pair_sample_0336 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VN.t0 VDD2.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X1 VTAIL.t18 VP.t0 VDD1.t9 B.t21 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X2 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=0 ps=0 w=11.68 l=0.62
X3 VDD2.t5 VN.t1 VTAIL.t15 B.t23 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=4.5552 ps=24.14 w=11.68 l=0.62
X4 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=0 ps=0 w=11.68 l=0.62
X5 VDD2.t8 VN.t2 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=1.9272 ps=12.01 w=11.68 l=0.62
X6 VTAIL.t13 VN.t3 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X7 VDD1.t8 VP.t1 VTAIL.t19 B.t22 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=4.5552 ps=24.14 w=11.68 l=0.62
X8 VTAIL.t4 VP.t2 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X9 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=0 ps=0 w=11.68 l=0.62
X10 VDD1.t6 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=1.9272 ps=12.01 w=11.68 l=0.62
X11 VTAIL.t6 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X12 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X13 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=0 ps=0 w=11.68 l=0.62
X14 VTAIL.t2 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X15 VDD1.t2 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=1.9272 ps=12.01 w=11.68 l=0.62
X16 VTAIL.t12 VN.t4 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X17 VDD2.t6 VN.t5 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=4.5552 ps=24.14 w=11.68 l=0.62
X18 VDD1.t1 VP.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X19 VDD2.t3 VN.t6 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=4.5552 pd=24.14 as=1.9272 ps=12.01 w=11.68 l=0.62
X20 VTAIL.t9 VN.t7 VDD2.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X21 VDD2.t4 VN.t8 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
X22 VDD1.t0 VP.t9 VTAIL.t17 B.t23 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=4.5552 ps=24.14 w=11.68 l=0.62
X23 VDD2.t2 VN.t9 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9272 pd=12.01 as=1.9272 ps=12.01 w=11.68 l=0.62
R0 VN.n2 VN.t6 544.194
R1 VN.n10 VN.t5 544.194
R2 VN.n1 VN.t7 517.374
R3 VN.n4 VN.t9 517.374
R4 VN.n5 VN.t0 517.374
R5 VN.n6 VN.t1 517.374
R6 VN.n9 VN.t3 517.374
R7 VN.n12 VN.t8 517.374
R8 VN.n13 VN.t4 517.374
R9 VN.n14 VN.t2 517.374
R10 VN.n7 VN.n6 161.3
R11 VN.n15 VN.n14 161.3
R12 VN.n13 VN.n8 80.6037
R13 VN.n12 VN.n11 80.6037
R14 VN.n5 VN.n0 80.6037
R15 VN.n4 VN.n3 80.6037
R16 VN.n4 VN.n1 48.2005
R17 VN.n5 VN.n4 48.2005
R18 VN.n6 VN.n5 48.2005
R19 VN.n12 VN.n9 48.2005
R20 VN.n13 VN.n12 48.2005
R21 VN.n14 VN.n13 48.2005
R22 VN.n11 VN.n10 45.2318
R23 VN.n3 VN.n2 45.2318
R24 VN VN.n15 42.5365
R25 VN.n10 VN.n9 13.3799
R26 VN.n2 VN.n1 13.3799
R27 VN.n11 VN.n8 0.380177
R28 VN.n3 VN.n0 0.380177
R29 VN.n15 VN.n8 0.285035
R30 VN.n7 VN.n0 0.285035
R31 VN VN.n7 0.0516364
R32 VDD2.n1 VDD2.t3 62.9425
R33 VDD2.n4 VDD2.t8 62.1237
R34 VDD2.n3 VDD2.n2 60.9872
R35 VDD2 VDD2.n7 60.9844
R36 VDD2.n6 VDD2.n5 60.4285
R37 VDD2.n1 VDD2.n0 60.4283
R38 VDD2.n4 VDD2.n3 37.6743
R39 VDD2.n7 VDD2.t0 1.69571
R40 VDD2.n7 VDD2.t6 1.69571
R41 VDD2.n5 VDD2.t1 1.69571
R42 VDD2.n5 VDD2.t4 1.69571
R43 VDD2.n2 VDD2.t9 1.69571
R44 VDD2.n2 VDD2.t5 1.69571
R45 VDD2.n0 VDD2.t7 1.69571
R46 VDD2.n0 VDD2.t2 1.69571
R47 VDD2.n6 VDD2.n4 0.819465
R48 VDD2 VDD2.n6 0.263431
R49 VDD2.n3 VDD2.n1 0.149895
R50 VTAIL.n11 VTAIL.t11 45.4449
R51 VTAIL.n17 VTAIL.t15 45.4447
R52 VTAIL.n2 VTAIL.t19 45.4447
R53 VTAIL.n16 VTAIL.t17 45.4447
R54 VTAIL.n15 VTAIL.n14 43.7497
R55 VTAIL.n13 VTAIL.n12 43.7497
R56 VTAIL.n10 VTAIL.n9 43.7497
R57 VTAIL.n8 VTAIL.n7 43.7497
R58 VTAIL.n19 VTAIL.n18 43.7495
R59 VTAIL.n1 VTAIL.n0 43.7495
R60 VTAIL.n4 VTAIL.n3 43.7495
R61 VTAIL.n6 VTAIL.n5 43.7495
R62 VTAIL.n8 VTAIL.n6 24.0738
R63 VTAIL.n17 VTAIL.n16 23.2548
R64 VTAIL.n18 VTAIL.t7 1.69571
R65 VTAIL.n18 VTAIL.t16 1.69571
R66 VTAIL.n0 VTAIL.t10 1.69571
R67 VTAIL.n0 VTAIL.t9 1.69571
R68 VTAIL.n3 VTAIL.t1 1.69571
R69 VTAIL.n3 VTAIL.t6 1.69571
R70 VTAIL.n5 VTAIL.t5 1.69571
R71 VTAIL.n5 VTAIL.t2 1.69571
R72 VTAIL.n14 VTAIL.t0 1.69571
R73 VTAIL.n14 VTAIL.t4 1.69571
R74 VTAIL.n12 VTAIL.t3 1.69571
R75 VTAIL.n12 VTAIL.t18 1.69571
R76 VTAIL.n9 VTAIL.t8 1.69571
R77 VTAIL.n9 VTAIL.t13 1.69571
R78 VTAIL.n7 VTAIL.t14 1.69571
R79 VTAIL.n7 VTAIL.t12 1.69571
R80 VTAIL.n13 VTAIL.n11 0.87981
R81 VTAIL.n2 VTAIL.n1 0.87981
R82 VTAIL.n10 VTAIL.n8 0.819465
R83 VTAIL.n11 VTAIL.n10 0.819465
R84 VTAIL.n15 VTAIL.n13 0.819465
R85 VTAIL.n16 VTAIL.n15 0.819465
R86 VTAIL.n6 VTAIL.n4 0.819465
R87 VTAIL.n4 VTAIL.n2 0.819465
R88 VTAIL.n19 VTAIL.n17 0.819465
R89 VTAIL VTAIL.n1 0.672914
R90 VTAIL VTAIL.n19 0.147052
R91 B.n375 B.t11 658.088
R92 B.n372 B.t7 658.088
R93 B.n97 B.t14 658.088
R94 B.n94 B.t18 658.088
R95 B.n667 B.n666 585
R96 B.n668 B.n667 585
R97 B.n278 B.n93 585
R98 B.n277 B.n276 585
R99 B.n275 B.n274 585
R100 B.n273 B.n272 585
R101 B.n271 B.n270 585
R102 B.n269 B.n268 585
R103 B.n267 B.n266 585
R104 B.n265 B.n264 585
R105 B.n263 B.n262 585
R106 B.n261 B.n260 585
R107 B.n259 B.n258 585
R108 B.n257 B.n256 585
R109 B.n255 B.n254 585
R110 B.n253 B.n252 585
R111 B.n251 B.n250 585
R112 B.n249 B.n248 585
R113 B.n247 B.n246 585
R114 B.n245 B.n244 585
R115 B.n243 B.n242 585
R116 B.n241 B.n240 585
R117 B.n239 B.n238 585
R118 B.n237 B.n236 585
R119 B.n235 B.n234 585
R120 B.n233 B.n232 585
R121 B.n231 B.n230 585
R122 B.n229 B.n228 585
R123 B.n227 B.n226 585
R124 B.n225 B.n224 585
R125 B.n223 B.n222 585
R126 B.n221 B.n220 585
R127 B.n219 B.n218 585
R128 B.n217 B.n216 585
R129 B.n215 B.n214 585
R130 B.n213 B.n212 585
R131 B.n211 B.n210 585
R132 B.n209 B.n208 585
R133 B.n207 B.n206 585
R134 B.n205 B.n204 585
R135 B.n203 B.n202 585
R136 B.n201 B.n200 585
R137 B.n199 B.n198 585
R138 B.n197 B.n196 585
R139 B.n195 B.n194 585
R140 B.n193 B.n192 585
R141 B.n191 B.n190 585
R142 B.n189 B.n188 585
R143 B.n187 B.n186 585
R144 B.n185 B.n184 585
R145 B.n183 B.n182 585
R146 B.n180 B.n179 585
R147 B.n178 B.n177 585
R148 B.n176 B.n175 585
R149 B.n174 B.n173 585
R150 B.n172 B.n171 585
R151 B.n170 B.n169 585
R152 B.n168 B.n167 585
R153 B.n166 B.n165 585
R154 B.n164 B.n163 585
R155 B.n162 B.n161 585
R156 B.n160 B.n159 585
R157 B.n158 B.n157 585
R158 B.n156 B.n155 585
R159 B.n154 B.n153 585
R160 B.n152 B.n151 585
R161 B.n150 B.n149 585
R162 B.n148 B.n147 585
R163 B.n146 B.n145 585
R164 B.n144 B.n143 585
R165 B.n142 B.n141 585
R166 B.n140 B.n139 585
R167 B.n138 B.n137 585
R168 B.n136 B.n135 585
R169 B.n134 B.n133 585
R170 B.n132 B.n131 585
R171 B.n130 B.n129 585
R172 B.n128 B.n127 585
R173 B.n126 B.n125 585
R174 B.n124 B.n123 585
R175 B.n122 B.n121 585
R176 B.n120 B.n119 585
R177 B.n118 B.n117 585
R178 B.n116 B.n115 585
R179 B.n114 B.n113 585
R180 B.n112 B.n111 585
R181 B.n110 B.n109 585
R182 B.n108 B.n107 585
R183 B.n106 B.n105 585
R184 B.n104 B.n103 585
R185 B.n102 B.n101 585
R186 B.n100 B.n99 585
R187 B.n665 B.n47 585
R188 B.n669 B.n47 585
R189 B.n664 B.n46 585
R190 B.n670 B.n46 585
R191 B.n663 B.n662 585
R192 B.n662 B.n42 585
R193 B.n661 B.n41 585
R194 B.n676 B.n41 585
R195 B.n660 B.n40 585
R196 B.n677 B.n40 585
R197 B.n659 B.n39 585
R198 B.n678 B.n39 585
R199 B.n658 B.n657 585
R200 B.n657 B.n35 585
R201 B.n656 B.n34 585
R202 B.n684 B.n34 585
R203 B.n655 B.n33 585
R204 B.n685 B.n33 585
R205 B.n654 B.n32 585
R206 B.n686 B.n32 585
R207 B.n653 B.n652 585
R208 B.n652 B.n31 585
R209 B.n651 B.n27 585
R210 B.n692 B.n27 585
R211 B.n650 B.n26 585
R212 B.n693 B.n26 585
R213 B.n649 B.n25 585
R214 B.n694 B.n25 585
R215 B.n648 B.n647 585
R216 B.n647 B.n21 585
R217 B.n646 B.n20 585
R218 B.n700 B.n20 585
R219 B.n645 B.n19 585
R220 B.n701 B.n19 585
R221 B.n644 B.n18 585
R222 B.n702 B.n18 585
R223 B.n643 B.n642 585
R224 B.n642 B.n14 585
R225 B.n641 B.n13 585
R226 B.n708 B.n13 585
R227 B.n640 B.n12 585
R228 B.n709 B.n12 585
R229 B.n639 B.n11 585
R230 B.n710 B.n11 585
R231 B.n638 B.n637 585
R232 B.n637 B.t3 585
R233 B.n636 B.n7 585
R234 B.n716 B.n7 585
R235 B.n635 B.n6 585
R236 B.n717 B.n6 585
R237 B.n634 B.n5 585
R238 B.n718 B.n5 585
R239 B.n633 B.n632 585
R240 B.n632 B.n4 585
R241 B.n631 B.n279 585
R242 B.n631 B.n630 585
R243 B.n621 B.n280 585
R244 B.t22 B.n280 585
R245 B.n623 B.n622 585
R246 B.n624 B.n623 585
R247 B.n620 B.n285 585
R248 B.n285 B.n284 585
R249 B.n619 B.n618 585
R250 B.n618 B.n617 585
R251 B.n287 B.n286 585
R252 B.n288 B.n287 585
R253 B.n610 B.n609 585
R254 B.n611 B.n610 585
R255 B.n608 B.n292 585
R256 B.n296 B.n292 585
R257 B.n607 B.n606 585
R258 B.n606 B.n605 585
R259 B.n294 B.n293 585
R260 B.n295 B.n294 585
R261 B.n598 B.n597 585
R262 B.n599 B.n598 585
R263 B.n596 B.n301 585
R264 B.n301 B.n300 585
R265 B.n595 B.n594 585
R266 B.n594 B.n593 585
R267 B.n303 B.n302 585
R268 B.n586 B.n303 585
R269 B.n585 B.n584 585
R270 B.n587 B.n585 585
R271 B.n583 B.n308 585
R272 B.n308 B.n307 585
R273 B.n582 B.n581 585
R274 B.n581 B.n580 585
R275 B.n310 B.n309 585
R276 B.n311 B.n310 585
R277 B.n573 B.n572 585
R278 B.n574 B.n573 585
R279 B.n571 B.n315 585
R280 B.n319 B.n315 585
R281 B.n570 B.n569 585
R282 B.n569 B.n568 585
R283 B.n317 B.n316 585
R284 B.n318 B.n317 585
R285 B.n561 B.n560 585
R286 B.n562 B.n561 585
R287 B.n559 B.n324 585
R288 B.n324 B.n323 585
R289 B.n553 B.n552 585
R290 B.n551 B.n371 585
R291 B.n550 B.n370 585
R292 B.n555 B.n370 585
R293 B.n549 B.n548 585
R294 B.n547 B.n546 585
R295 B.n545 B.n544 585
R296 B.n543 B.n542 585
R297 B.n541 B.n540 585
R298 B.n539 B.n538 585
R299 B.n537 B.n536 585
R300 B.n535 B.n534 585
R301 B.n533 B.n532 585
R302 B.n531 B.n530 585
R303 B.n529 B.n528 585
R304 B.n527 B.n526 585
R305 B.n525 B.n524 585
R306 B.n523 B.n522 585
R307 B.n521 B.n520 585
R308 B.n519 B.n518 585
R309 B.n517 B.n516 585
R310 B.n515 B.n514 585
R311 B.n513 B.n512 585
R312 B.n511 B.n510 585
R313 B.n509 B.n508 585
R314 B.n507 B.n506 585
R315 B.n505 B.n504 585
R316 B.n503 B.n502 585
R317 B.n501 B.n500 585
R318 B.n499 B.n498 585
R319 B.n497 B.n496 585
R320 B.n495 B.n494 585
R321 B.n493 B.n492 585
R322 B.n491 B.n490 585
R323 B.n489 B.n488 585
R324 B.n487 B.n486 585
R325 B.n485 B.n484 585
R326 B.n483 B.n482 585
R327 B.n481 B.n480 585
R328 B.n479 B.n478 585
R329 B.n477 B.n476 585
R330 B.n475 B.n474 585
R331 B.n473 B.n472 585
R332 B.n471 B.n470 585
R333 B.n469 B.n468 585
R334 B.n467 B.n466 585
R335 B.n465 B.n464 585
R336 B.n463 B.n462 585
R337 B.n461 B.n460 585
R338 B.n459 B.n458 585
R339 B.n457 B.n456 585
R340 B.n454 B.n453 585
R341 B.n452 B.n451 585
R342 B.n450 B.n449 585
R343 B.n448 B.n447 585
R344 B.n446 B.n445 585
R345 B.n444 B.n443 585
R346 B.n442 B.n441 585
R347 B.n440 B.n439 585
R348 B.n438 B.n437 585
R349 B.n436 B.n435 585
R350 B.n434 B.n433 585
R351 B.n432 B.n431 585
R352 B.n430 B.n429 585
R353 B.n428 B.n427 585
R354 B.n426 B.n425 585
R355 B.n424 B.n423 585
R356 B.n422 B.n421 585
R357 B.n420 B.n419 585
R358 B.n418 B.n417 585
R359 B.n416 B.n415 585
R360 B.n414 B.n413 585
R361 B.n412 B.n411 585
R362 B.n410 B.n409 585
R363 B.n408 B.n407 585
R364 B.n406 B.n405 585
R365 B.n404 B.n403 585
R366 B.n402 B.n401 585
R367 B.n400 B.n399 585
R368 B.n398 B.n397 585
R369 B.n396 B.n395 585
R370 B.n394 B.n393 585
R371 B.n392 B.n391 585
R372 B.n390 B.n389 585
R373 B.n388 B.n387 585
R374 B.n386 B.n385 585
R375 B.n384 B.n383 585
R376 B.n382 B.n381 585
R377 B.n380 B.n379 585
R378 B.n378 B.n377 585
R379 B.n326 B.n325 585
R380 B.n558 B.n557 585
R381 B.n322 B.n321 585
R382 B.n323 B.n322 585
R383 B.n564 B.n563 585
R384 B.n563 B.n562 585
R385 B.n565 B.n320 585
R386 B.n320 B.n318 585
R387 B.n567 B.n566 585
R388 B.n568 B.n567 585
R389 B.n314 B.n313 585
R390 B.n319 B.n314 585
R391 B.n576 B.n575 585
R392 B.n575 B.n574 585
R393 B.n577 B.n312 585
R394 B.n312 B.n311 585
R395 B.n579 B.n578 585
R396 B.n580 B.n579 585
R397 B.n306 B.n305 585
R398 B.n307 B.n306 585
R399 B.n589 B.n588 585
R400 B.n588 B.n587 585
R401 B.n590 B.n304 585
R402 B.n586 B.n304 585
R403 B.n592 B.n591 585
R404 B.n593 B.n592 585
R405 B.n299 B.n298 585
R406 B.n300 B.n299 585
R407 B.n601 B.n600 585
R408 B.n600 B.n599 585
R409 B.n602 B.n297 585
R410 B.n297 B.n295 585
R411 B.n604 B.n603 585
R412 B.n605 B.n604 585
R413 B.n291 B.n290 585
R414 B.n296 B.n291 585
R415 B.n613 B.n612 585
R416 B.n612 B.n611 585
R417 B.n614 B.n289 585
R418 B.n289 B.n288 585
R419 B.n616 B.n615 585
R420 B.n617 B.n616 585
R421 B.n283 B.n282 585
R422 B.n284 B.n283 585
R423 B.n626 B.n625 585
R424 B.n625 B.n624 585
R425 B.n627 B.n281 585
R426 B.n281 B.t22 585
R427 B.n629 B.n628 585
R428 B.n630 B.n629 585
R429 B.n2 B.n0 585
R430 B.n4 B.n2 585
R431 B.n3 B.n1 585
R432 B.n717 B.n3 585
R433 B.n715 B.n714 585
R434 B.n716 B.n715 585
R435 B.n713 B.n8 585
R436 B.n8 B.t3 585
R437 B.n712 B.n711 585
R438 B.n711 B.n710 585
R439 B.n10 B.n9 585
R440 B.n709 B.n10 585
R441 B.n707 B.n706 585
R442 B.n708 B.n707 585
R443 B.n705 B.n15 585
R444 B.n15 B.n14 585
R445 B.n704 B.n703 585
R446 B.n703 B.n702 585
R447 B.n17 B.n16 585
R448 B.n701 B.n17 585
R449 B.n699 B.n698 585
R450 B.n700 B.n699 585
R451 B.n697 B.n22 585
R452 B.n22 B.n21 585
R453 B.n696 B.n695 585
R454 B.n695 B.n694 585
R455 B.n24 B.n23 585
R456 B.n693 B.n24 585
R457 B.n691 B.n690 585
R458 B.n692 B.n691 585
R459 B.n689 B.n28 585
R460 B.n31 B.n28 585
R461 B.n688 B.n687 585
R462 B.n687 B.n686 585
R463 B.n30 B.n29 585
R464 B.n685 B.n30 585
R465 B.n683 B.n682 585
R466 B.n684 B.n683 585
R467 B.n681 B.n36 585
R468 B.n36 B.n35 585
R469 B.n680 B.n679 585
R470 B.n679 B.n678 585
R471 B.n38 B.n37 585
R472 B.n677 B.n38 585
R473 B.n675 B.n674 585
R474 B.n676 B.n675 585
R475 B.n673 B.n43 585
R476 B.n43 B.n42 585
R477 B.n672 B.n671 585
R478 B.n671 B.n670 585
R479 B.n45 B.n44 585
R480 B.n669 B.n45 585
R481 B.n720 B.n719 585
R482 B.n719 B.n718 585
R483 B.n553 B.n322 473.281
R484 B.n99 B.n45 473.281
R485 B.n557 B.n324 473.281
R486 B.n667 B.n47 473.281
R487 B.n668 B.n92 256.663
R488 B.n668 B.n91 256.663
R489 B.n668 B.n90 256.663
R490 B.n668 B.n89 256.663
R491 B.n668 B.n88 256.663
R492 B.n668 B.n87 256.663
R493 B.n668 B.n86 256.663
R494 B.n668 B.n85 256.663
R495 B.n668 B.n84 256.663
R496 B.n668 B.n83 256.663
R497 B.n668 B.n82 256.663
R498 B.n668 B.n81 256.663
R499 B.n668 B.n80 256.663
R500 B.n668 B.n79 256.663
R501 B.n668 B.n78 256.663
R502 B.n668 B.n77 256.663
R503 B.n668 B.n76 256.663
R504 B.n668 B.n75 256.663
R505 B.n668 B.n74 256.663
R506 B.n668 B.n73 256.663
R507 B.n668 B.n72 256.663
R508 B.n668 B.n71 256.663
R509 B.n668 B.n70 256.663
R510 B.n668 B.n69 256.663
R511 B.n668 B.n68 256.663
R512 B.n668 B.n67 256.663
R513 B.n668 B.n66 256.663
R514 B.n668 B.n65 256.663
R515 B.n668 B.n64 256.663
R516 B.n668 B.n63 256.663
R517 B.n668 B.n62 256.663
R518 B.n668 B.n61 256.663
R519 B.n668 B.n60 256.663
R520 B.n668 B.n59 256.663
R521 B.n668 B.n58 256.663
R522 B.n668 B.n57 256.663
R523 B.n668 B.n56 256.663
R524 B.n668 B.n55 256.663
R525 B.n668 B.n54 256.663
R526 B.n668 B.n53 256.663
R527 B.n668 B.n52 256.663
R528 B.n668 B.n51 256.663
R529 B.n668 B.n50 256.663
R530 B.n668 B.n49 256.663
R531 B.n668 B.n48 256.663
R532 B.n555 B.n554 256.663
R533 B.n555 B.n327 256.663
R534 B.n555 B.n328 256.663
R535 B.n555 B.n329 256.663
R536 B.n555 B.n330 256.663
R537 B.n555 B.n331 256.663
R538 B.n555 B.n332 256.663
R539 B.n555 B.n333 256.663
R540 B.n555 B.n334 256.663
R541 B.n555 B.n335 256.663
R542 B.n555 B.n336 256.663
R543 B.n555 B.n337 256.663
R544 B.n555 B.n338 256.663
R545 B.n555 B.n339 256.663
R546 B.n555 B.n340 256.663
R547 B.n555 B.n341 256.663
R548 B.n555 B.n342 256.663
R549 B.n555 B.n343 256.663
R550 B.n555 B.n344 256.663
R551 B.n555 B.n345 256.663
R552 B.n555 B.n346 256.663
R553 B.n555 B.n347 256.663
R554 B.n555 B.n348 256.663
R555 B.n555 B.n349 256.663
R556 B.n555 B.n350 256.663
R557 B.n555 B.n351 256.663
R558 B.n555 B.n352 256.663
R559 B.n555 B.n353 256.663
R560 B.n555 B.n354 256.663
R561 B.n555 B.n355 256.663
R562 B.n555 B.n356 256.663
R563 B.n555 B.n357 256.663
R564 B.n555 B.n358 256.663
R565 B.n555 B.n359 256.663
R566 B.n555 B.n360 256.663
R567 B.n555 B.n361 256.663
R568 B.n555 B.n362 256.663
R569 B.n555 B.n363 256.663
R570 B.n555 B.n364 256.663
R571 B.n555 B.n365 256.663
R572 B.n555 B.n366 256.663
R573 B.n555 B.n367 256.663
R574 B.n555 B.n368 256.663
R575 B.n555 B.n369 256.663
R576 B.n556 B.n555 256.663
R577 B.n563 B.n322 163.367
R578 B.n563 B.n320 163.367
R579 B.n567 B.n320 163.367
R580 B.n567 B.n314 163.367
R581 B.n575 B.n314 163.367
R582 B.n575 B.n312 163.367
R583 B.n579 B.n312 163.367
R584 B.n579 B.n306 163.367
R585 B.n588 B.n306 163.367
R586 B.n588 B.n304 163.367
R587 B.n592 B.n304 163.367
R588 B.n592 B.n299 163.367
R589 B.n600 B.n299 163.367
R590 B.n600 B.n297 163.367
R591 B.n604 B.n297 163.367
R592 B.n604 B.n291 163.367
R593 B.n612 B.n291 163.367
R594 B.n612 B.n289 163.367
R595 B.n616 B.n289 163.367
R596 B.n616 B.n283 163.367
R597 B.n625 B.n283 163.367
R598 B.n625 B.n281 163.367
R599 B.n629 B.n281 163.367
R600 B.n629 B.n2 163.367
R601 B.n719 B.n2 163.367
R602 B.n719 B.n3 163.367
R603 B.n715 B.n3 163.367
R604 B.n715 B.n8 163.367
R605 B.n711 B.n8 163.367
R606 B.n711 B.n10 163.367
R607 B.n707 B.n10 163.367
R608 B.n707 B.n15 163.367
R609 B.n703 B.n15 163.367
R610 B.n703 B.n17 163.367
R611 B.n699 B.n17 163.367
R612 B.n699 B.n22 163.367
R613 B.n695 B.n22 163.367
R614 B.n695 B.n24 163.367
R615 B.n691 B.n24 163.367
R616 B.n691 B.n28 163.367
R617 B.n687 B.n28 163.367
R618 B.n687 B.n30 163.367
R619 B.n683 B.n30 163.367
R620 B.n683 B.n36 163.367
R621 B.n679 B.n36 163.367
R622 B.n679 B.n38 163.367
R623 B.n675 B.n38 163.367
R624 B.n675 B.n43 163.367
R625 B.n671 B.n43 163.367
R626 B.n671 B.n45 163.367
R627 B.n371 B.n370 163.367
R628 B.n548 B.n370 163.367
R629 B.n546 B.n545 163.367
R630 B.n542 B.n541 163.367
R631 B.n538 B.n537 163.367
R632 B.n534 B.n533 163.367
R633 B.n530 B.n529 163.367
R634 B.n526 B.n525 163.367
R635 B.n522 B.n521 163.367
R636 B.n518 B.n517 163.367
R637 B.n514 B.n513 163.367
R638 B.n510 B.n509 163.367
R639 B.n506 B.n505 163.367
R640 B.n502 B.n501 163.367
R641 B.n498 B.n497 163.367
R642 B.n494 B.n493 163.367
R643 B.n490 B.n489 163.367
R644 B.n486 B.n485 163.367
R645 B.n482 B.n481 163.367
R646 B.n478 B.n477 163.367
R647 B.n474 B.n473 163.367
R648 B.n470 B.n469 163.367
R649 B.n466 B.n465 163.367
R650 B.n462 B.n461 163.367
R651 B.n458 B.n457 163.367
R652 B.n453 B.n452 163.367
R653 B.n449 B.n448 163.367
R654 B.n445 B.n444 163.367
R655 B.n441 B.n440 163.367
R656 B.n437 B.n436 163.367
R657 B.n433 B.n432 163.367
R658 B.n429 B.n428 163.367
R659 B.n425 B.n424 163.367
R660 B.n421 B.n420 163.367
R661 B.n417 B.n416 163.367
R662 B.n413 B.n412 163.367
R663 B.n409 B.n408 163.367
R664 B.n405 B.n404 163.367
R665 B.n401 B.n400 163.367
R666 B.n397 B.n396 163.367
R667 B.n393 B.n392 163.367
R668 B.n389 B.n388 163.367
R669 B.n385 B.n384 163.367
R670 B.n381 B.n380 163.367
R671 B.n377 B.n326 163.367
R672 B.n561 B.n324 163.367
R673 B.n561 B.n317 163.367
R674 B.n569 B.n317 163.367
R675 B.n569 B.n315 163.367
R676 B.n573 B.n315 163.367
R677 B.n573 B.n310 163.367
R678 B.n581 B.n310 163.367
R679 B.n581 B.n308 163.367
R680 B.n585 B.n308 163.367
R681 B.n585 B.n303 163.367
R682 B.n594 B.n303 163.367
R683 B.n594 B.n301 163.367
R684 B.n598 B.n301 163.367
R685 B.n598 B.n294 163.367
R686 B.n606 B.n294 163.367
R687 B.n606 B.n292 163.367
R688 B.n610 B.n292 163.367
R689 B.n610 B.n287 163.367
R690 B.n618 B.n287 163.367
R691 B.n618 B.n285 163.367
R692 B.n623 B.n285 163.367
R693 B.n623 B.n280 163.367
R694 B.n631 B.n280 163.367
R695 B.n632 B.n631 163.367
R696 B.n632 B.n5 163.367
R697 B.n6 B.n5 163.367
R698 B.n7 B.n6 163.367
R699 B.n637 B.n7 163.367
R700 B.n637 B.n11 163.367
R701 B.n12 B.n11 163.367
R702 B.n13 B.n12 163.367
R703 B.n642 B.n13 163.367
R704 B.n642 B.n18 163.367
R705 B.n19 B.n18 163.367
R706 B.n20 B.n19 163.367
R707 B.n647 B.n20 163.367
R708 B.n647 B.n25 163.367
R709 B.n26 B.n25 163.367
R710 B.n27 B.n26 163.367
R711 B.n652 B.n27 163.367
R712 B.n652 B.n32 163.367
R713 B.n33 B.n32 163.367
R714 B.n34 B.n33 163.367
R715 B.n657 B.n34 163.367
R716 B.n657 B.n39 163.367
R717 B.n40 B.n39 163.367
R718 B.n41 B.n40 163.367
R719 B.n662 B.n41 163.367
R720 B.n662 B.n46 163.367
R721 B.n47 B.n46 163.367
R722 B.n103 B.n102 163.367
R723 B.n107 B.n106 163.367
R724 B.n111 B.n110 163.367
R725 B.n115 B.n114 163.367
R726 B.n119 B.n118 163.367
R727 B.n123 B.n122 163.367
R728 B.n127 B.n126 163.367
R729 B.n131 B.n130 163.367
R730 B.n135 B.n134 163.367
R731 B.n139 B.n138 163.367
R732 B.n143 B.n142 163.367
R733 B.n147 B.n146 163.367
R734 B.n151 B.n150 163.367
R735 B.n155 B.n154 163.367
R736 B.n159 B.n158 163.367
R737 B.n163 B.n162 163.367
R738 B.n167 B.n166 163.367
R739 B.n171 B.n170 163.367
R740 B.n175 B.n174 163.367
R741 B.n179 B.n178 163.367
R742 B.n184 B.n183 163.367
R743 B.n188 B.n187 163.367
R744 B.n192 B.n191 163.367
R745 B.n196 B.n195 163.367
R746 B.n200 B.n199 163.367
R747 B.n204 B.n203 163.367
R748 B.n208 B.n207 163.367
R749 B.n212 B.n211 163.367
R750 B.n216 B.n215 163.367
R751 B.n220 B.n219 163.367
R752 B.n224 B.n223 163.367
R753 B.n228 B.n227 163.367
R754 B.n232 B.n231 163.367
R755 B.n236 B.n235 163.367
R756 B.n240 B.n239 163.367
R757 B.n244 B.n243 163.367
R758 B.n248 B.n247 163.367
R759 B.n252 B.n251 163.367
R760 B.n256 B.n255 163.367
R761 B.n260 B.n259 163.367
R762 B.n264 B.n263 163.367
R763 B.n268 B.n267 163.367
R764 B.n272 B.n271 163.367
R765 B.n276 B.n275 163.367
R766 B.n667 B.n93 163.367
R767 B.n375 B.t13 88.5861
R768 B.n94 B.t19 88.5861
R769 B.n372 B.t10 88.5714
R770 B.n97 B.t16 88.5714
R771 B.n555 B.n323 74.6098
R772 B.n669 B.n668 74.6098
R773 B.n554 B.n553 71.676
R774 B.n548 B.n327 71.676
R775 B.n545 B.n328 71.676
R776 B.n541 B.n329 71.676
R777 B.n537 B.n330 71.676
R778 B.n533 B.n331 71.676
R779 B.n529 B.n332 71.676
R780 B.n525 B.n333 71.676
R781 B.n521 B.n334 71.676
R782 B.n517 B.n335 71.676
R783 B.n513 B.n336 71.676
R784 B.n509 B.n337 71.676
R785 B.n505 B.n338 71.676
R786 B.n501 B.n339 71.676
R787 B.n497 B.n340 71.676
R788 B.n493 B.n341 71.676
R789 B.n489 B.n342 71.676
R790 B.n485 B.n343 71.676
R791 B.n481 B.n344 71.676
R792 B.n477 B.n345 71.676
R793 B.n473 B.n346 71.676
R794 B.n469 B.n347 71.676
R795 B.n465 B.n348 71.676
R796 B.n461 B.n349 71.676
R797 B.n457 B.n350 71.676
R798 B.n452 B.n351 71.676
R799 B.n448 B.n352 71.676
R800 B.n444 B.n353 71.676
R801 B.n440 B.n354 71.676
R802 B.n436 B.n355 71.676
R803 B.n432 B.n356 71.676
R804 B.n428 B.n357 71.676
R805 B.n424 B.n358 71.676
R806 B.n420 B.n359 71.676
R807 B.n416 B.n360 71.676
R808 B.n412 B.n361 71.676
R809 B.n408 B.n362 71.676
R810 B.n404 B.n363 71.676
R811 B.n400 B.n364 71.676
R812 B.n396 B.n365 71.676
R813 B.n392 B.n366 71.676
R814 B.n388 B.n367 71.676
R815 B.n384 B.n368 71.676
R816 B.n380 B.n369 71.676
R817 B.n556 B.n326 71.676
R818 B.n99 B.n48 71.676
R819 B.n103 B.n49 71.676
R820 B.n107 B.n50 71.676
R821 B.n111 B.n51 71.676
R822 B.n115 B.n52 71.676
R823 B.n119 B.n53 71.676
R824 B.n123 B.n54 71.676
R825 B.n127 B.n55 71.676
R826 B.n131 B.n56 71.676
R827 B.n135 B.n57 71.676
R828 B.n139 B.n58 71.676
R829 B.n143 B.n59 71.676
R830 B.n147 B.n60 71.676
R831 B.n151 B.n61 71.676
R832 B.n155 B.n62 71.676
R833 B.n159 B.n63 71.676
R834 B.n163 B.n64 71.676
R835 B.n167 B.n65 71.676
R836 B.n171 B.n66 71.676
R837 B.n175 B.n67 71.676
R838 B.n179 B.n68 71.676
R839 B.n184 B.n69 71.676
R840 B.n188 B.n70 71.676
R841 B.n192 B.n71 71.676
R842 B.n196 B.n72 71.676
R843 B.n200 B.n73 71.676
R844 B.n204 B.n74 71.676
R845 B.n208 B.n75 71.676
R846 B.n212 B.n76 71.676
R847 B.n216 B.n77 71.676
R848 B.n220 B.n78 71.676
R849 B.n224 B.n79 71.676
R850 B.n228 B.n80 71.676
R851 B.n232 B.n81 71.676
R852 B.n236 B.n82 71.676
R853 B.n240 B.n83 71.676
R854 B.n244 B.n84 71.676
R855 B.n248 B.n85 71.676
R856 B.n252 B.n86 71.676
R857 B.n256 B.n87 71.676
R858 B.n260 B.n88 71.676
R859 B.n264 B.n89 71.676
R860 B.n268 B.n90 71.676
R861 B.n272 B.n91 71.676
R862 B.n276 B.n92 71.676
R863 B.n93 B.n92 71.676
R864 B.n275 B.n91 71.676
R865 B.n271 B.n90 71.676
R866 B.n267 B.n89 71.676
R867 B.n263 B.n88 71.676
R868 B.n259 B.n87 71.676
R869 B.n255 B.n86 71.676
R870 B.n251 B.n85 71.676
R871 B.n247 B.n84 71.676
R872 B.n243 B.n83 71.676
R873 B.n239 B.n82 71.676
R874 B.n235 B.n81 71.676
R875 B.n231 B.n80 71.676
R876 B.n227 B.n79 71.676
R877 B.n223 B.n78 71.676
R878 B.n219 B.n77 71.676
R879 B.n215 B.n76 71.676
R880 B.n211 B.n75 71.676
R881 B.n207 B.n74 71.676
R882 B.n203 B.n73 71.676
R883 B.n199 B.n72 71.676
R884 B.n195 B.n71 71.676
R885 B.n191 B.n70 71.676
R886 B.n187 B.n69 71.676
R887 B.n183 B.n68 71.676
R888 B.n178 B.n67 71.676
R889 B.n174 B.n66 71.676
R890 B.n170 B.n65 71.676
R891 B.n166 B.n64 71.676
R892 B.n162 B.n63 71.676
R893 B.n158 B.n62 71.676
R894 B.n154 B.n61 71.676
R895 B.n150 B.n60 71.676
R896 B.n146 B.n59 71.676
R897 B.n142 B.n58 71.676
R898 B.n138 B.n57 71.676
R899 B.n134 B.n56 71.676
R900 B.n130 B.n55 71.676
R901 B.n126 B.n54 71.676
R902 B.n122 B.n53 71.676
R903 B.n118 B.n52 71.676
R904 B.n114 B.n51 71.676
R905 B.n110 B.n50 71.676
R906 B.n106 B.n49 71.676
R907 B.n102 B.n48 71.676
R908 B.n554 B.n371 71.676
R909 B.n546 B.n327 71.676
R910 B.n542 B.n328 71.676
R911 B.n538 B.n329 71.676
R912 B.n534 B.n330 71.676
R913 B.n530 B.n331 71.676
R914 B.n526 B.n332 71.676
R915 B.n522 B.n333 71.676
R916 B.n518 B.n334 71.676
R917 B.n514 B.n335 71.676
R918 B.n510 B.n336 71.676
R919 B.n506 B.n337 71.676
R920 B.n502 B.n338 71.676
R921 B.n498 B.n339 71.676
R922 B.n494 B.n340 71.676
R923 B.n490 B.n341 71.676
R924 B.n486 B.n342 71.676
R925 B.n482 B.n343 71.676
R926 B.n478 B.n344 71.676
R927 B.n474 B.n345 71.676
R928 B.n470 B.n346 71.676
R929 B.n466 B.n347 71.676
R930 B.n462 B.n348 71.676
R931 B.n458 B.n349 71.676
R932 B.n453 B.n350 71.676
R933 B.n449 B.n351 71.676
R934 B.n445 B.n352 71.676
R935 B.n441 B.n353 71.676
R936 B.n437 B.n354 71.676
R937 B.n433 B.n355 71.676
R938 B.n429 B.n356 71.676
R939 B.n425 B.n357 71.676
R940 B.n421 B.n358 71.676
R941 B.n417 B.n359 71.676
R942 B.n413 B.n360 71.676
R943 B.n409 B.n361 71.676
R944 B.n405 B.n362 71.676
R945 B.n401 B.n363 71.676
R946 B.n397 B.n364 71.676
R947 B.n393 B.n365 71.676
R948 B.n389 B.n366 71.676
R949 B.n385 B.n367 71.676
R950 B.n381 B.n368 71.676
R951 B.n377 B.n369 71.676
R952 B.n557 B.n556 71.676
R953 B.n376 B.t12 70.1619
R954 B.n95 B.t20 70.1619
R955 B.n373 B.t9 70.1471
R956 B.n98 B.t17 70.1471
R957 B.n455 B.n376 59.5399
R958 B.n374 B.n373 59.5399
R959 B.n181 B.n98 59.5399
R960 B.n96 B.n95 59.5399
R961 B.n562 B.n323 44.1173
R962 B.n562 B.n318 44.1173
R963 B.n568 B.n318 44.1173
R964 B.n568 B.n319 44.1173
R965 B.n574 B.n311 44.1173
R966 B.n580 B.n311 44.1173
R967 B.n580 B.n307 44.1173
R968 B.n587 B.n307 44.1173
R969 B.n587 B.n586 44.1173
R970 B.n593 B.n300 44.1173
R971 B.n599 B.n300 44.1173
R972 B.n605 B.n295 44.1173
R973 B.n605 B.n296 44.1173
R974 B.n611 B.n288 44.1173
R975 B.n617 B.n288 44.1173
R976 B.n624 B.n284 44.1173
R977 B.n624 B.t22 44.1173
R978 B.n630 B.t22 44.1173
R979 B.n630 B.n4 44.1173
R980 B.n718 B.n4 44.1173
R981 B.n718 B.n717 44.1173
R982 B.n717 B.n716 44.1173
R983 B.n716 B.t3 44.1173
R984 B.n710 B.t3 44.1173
R985 B.n710 B.n709 44.1173
R986 B.n708 B.n14 44.1173
R987 B.n702 B.n14 44.1173
R988 B.n701 B.n700 44.1173
R989 B.n700 B.n21 44.1173
R990 B.n694 B.n693 44.1173
R991 B.n693 B.n692 44.1173
R992 B.n686 B.n31 44.1173
R993 B.n686 B.n685 44.1173
R994 B.n685 B.n684 44.1173
R995 B.n684 B.n35 44.1173
R996 B.n678 B.n35 44.1173
R997 B.n677 B.n676 44.1173
R998 B.n676 B.n42 44.1173
R999 B.n670 B.n42 44.1173
R1000 B.n670 B.n669 44.1173
R1001 B.n319 B.t8 36.332
R1002 B.n586 B.t5 36.332
R1003 B.n31 B.t23 36.332
R1004 B.t15 B.n677 36.332
R1005 B.t6 B.n284 35.0344
R1006 B.n709 B.t21 35.0344
R1007 B.n100 B.n44 30.7517
R1008 B.n666 B.n665 30.7517
R1009 B.n559 B.n558 30.7517
R1010 B.n552 B.n321 30.7517
R1011 B.n599 B.t2 27.2491
R1012 B.n694 B.t4 27.2491
R1013 B.n611 B.t1 25.9515
R1014 B.n702 B.t0 25.9515
R1015 B.n376 B.n375 18.4247
R1016 B.n373 B.n372 18.4247
R1017 B.n98 B.n97 18.4247
R1018 B.n95 B.n94 18.4247
R1019 B.n296 B.t1 18.1662
R1020 B.t0 B.n701 18.1662
R1021 B B.n720 18.0485
R1022 B.t2 B.n295 16.8687
R1023 B.t4 B.n21 16.8687
R1024 B.n101 B.n100 10.6151
R1025 B.n104 B.n101 10.6151
R1026 B.n105 B.n104 10.6151
R1027 B.n108 B.n105 10.6151
R1028 B.n109 B.n108 10.6151
R1029 B.n112 B.n109 10.6151
R1030 B.n113 B.n112 10.6151
R1031 B.n116 B.n113 10.6151
R1032 B.n117 B.n116 10.6151
R1033 B.n120 B.n117 10.6151
R1034 B.n121 B.n120 10.6151
R1035 B.n124 B.n121 10.6151
R1036 B.n125 B.n124 10.6151
R1037 B.n128 B.n125 10.6151
R1038 B.n129 B.n128 10.6151
R1039 B.n132 B.n129 10.6151
R1040 B.n133 B.n132 10.6151
R1041 B.n136 B.n133 10.6151
R1042 B.n137 B.n136 10.6151
R1043 B.n140 B.n137 10.6151
R1044 B.n141 B.n140 10.6151
R1045 B.n144 B.n141 10.6151
R1046 B.n145 B.n144 10.6151
R1047 B.n148 B.n145 10.6151
R1048 B.n149 B.n148 10.6151
R1049 B.n152 B.n149 10.6151
R1050 B.n153 B.n152 10.6151
R1051 B.n156 B.n153 10.6151
R1052 B.n157 B.n156 10.6151
R1053 B.n160 B.n157 10.6151
R1054 B.n161 B.n160 10.6151
R1055 B.n164 B.n161 10.6151
R1056 B.n165 B.n164 10.6151
R1057 B.n168 B.n165 10.6151
R1058 B.n169 B.n168 10.6151
R1059 B.n172 B.n169 10.6151
R1060 B.n173 B.n172 10.6151
R1061 B.n176 B.n173 10.6151
R1062 B.n177 B.n176 10.6151
R1063 B.n180 B.n177 10.6151
R1064 B.n185 B.n182 10.6151
R1065 B.n186 B.n185 10.6151
R1066 B.n189 B.n186 10.6151
R1067 B.n190 B.n189 10.6151
R1068 B.n193 B.n190 10.6151
R1069 B.n194 B.n193 10.6151
R1070 B.n197 B.n194 10.6151
R1071 B.n198 B.n197 10.6151
R1072 B.n202 B.n201 10.6151
R1073 B.n205 B.n202 10.6151
R1074 B.n206 B.n205 10.6151
R1075 B.n209 B.n206 10.6151
R1076 B.n210 B.n209 10.6151
R1077 B.n213 B.n210 10.6151
R1078 B.n214 B.n213 10.6151
R1079 B.n217 B.n214 10.6151
R1080 B.n218 B.n217 10.6151
R1081 B.n221 B.n218 10.6151
R1082 B.n222 B.n221 10.6151
R1083 B.n225 B.n222 10.6151
R1084 B.n226 B.n225 10.6151
R1085 B.n229 B.n226 10.6151
R1086 B.n230 B.n229 10.6151
R1087 B.n233 B.n230 10.6151
R1088 B.n234 B.n233 10.6151
R1089 B.n237 B.n234 10.6151
R1090 B.n238 B.n237 10.6151
R1091 B.n241 B.n238 10.6151
R1092 B.n242 B.n241 10.6151
R1093 B.n245 B.n242 10.6151
R1094 B.n246 B.n245 10.6151
R1095 B.n249 B.n246 10.6151
R1096 B.n250 B.n249 10.6151
R1097 B.n253 B.n250 10.6151
R1098 B.n254 B.n253 10.6151
R1099 B.n257 B.n254 10.6151
R1100 B.n258 B.n257 10.6151
R1101 B.n261 B.n258 10.6151
R1102 B.n262 B.n261 10.6151
R1103 B.n265 B.n262 10.6151
R1104 B.n266 B.n265 10.6151
R1105 B.n269 B.n266 10.6151
R1106 B.n270 B.n269 10.6151
R1107 B.n273 B.n270 10.6151
R1108 B.n274 B.n273 10.6151
R1109 B.n277 B.n274 10.6151
R1110 B.n278 B.n277 10.6151
R1111 B.n666 B.n278 10.6151
R1112 B.n560 B.n559 10.6151
R1113 B.n560 B.n316 10.6151
R1114 B.n570 B.n316 10.6151
R1115 B.n571 B.n570 10.6151
R1116 B.n572 B.n571 10.6151
R1117 B.n572 B.n309 10.6151
R1118 B.n582 B.n309 10.6151
R1119 B.n583 B.n582 10.6151
R1120 B.n584 B.n583 10.6151
R1121 B.n584 B.n302 10.6151
R1122 B.n595 B.n302 10.6151
R1123 B.n596 B.n595 10.6151
R1124 B.n597 B.n596 10.6151
R1125 B.n597 B.n293 10.6151
R1126 B.n607 B.n293 10.6151
R1127 B.n608 B.n607 10.6151
R1128 B.n609 B.n608 10.6151
R1129 B.n609 B.n286 10.6151
R1130 B.n619 B.n286 10.6151
R1131 B.n620 B.n619 10.6151
R1132 B.n622 B.n620 10.6151
R1133 B.n622 B.n621 10.6151
R1134 B.n621 B.n279 10.6151
R1135 B.n633 B.n279 10.6151
R1136 B.n634 B.n633 10.6151
R1137 B.n635 B.n634 10.6151
R1138 B.n636 B.n635 10.6151
R1139 B.n638 B.n636 10.6151
R1140 B.n639 B.n638 10.6151
R1141 B.n640 B.n639 10.6151
R1142 B.n641 B.n640 10.6151
R1143 B.n643 B.n641 10.6151
R1144 B.n644 B.n643 10.6151
R1145 B.n645 B.n644 10.6151
R1146 B.n646 B.n645 10.6151
R1147 B.n648 B.n646 10.6151
R1148 B.n649 B.n648 10.6151
R1149 B.n650 B.n649 10.6151
R1150 B.n651 B.n650 10.6151
R1151 B.n653 B.n651 10.6151
R1152 B.n654 B.n653 10.6151
R1153 B.n655 B.n654 10.6151
R1154 B.n656 B.n655 10.6151
R1155 B.n658 B.n656 10.6151
R1156 B.n659 B.n658 10.6151
R1157 B.n660 B.n659 10.6151
R1158 B.n661 B.n660 10.6151
R1159 B.n663 B.n661 10.6151
R1160 B.n664 B.n663 10.6151
R1161 B.n665 B.n664 10.6151
R1162 B.n552 B.n551 10.6151
R1163 B.n551 B.n550 10.6151
R1164 B.n550 B.n549 10.6151
R1165 B.n549 B.n547 10.6151
R1166 B.n547 B.n544 10.6151
R1167 B.n544 B.n543 10.6151
R1168 B.n543 B.n540 10.6151
R1169 B.n540 B.n539 10.6151
R1170 B.n539 B.n536 10.6151
R1171 B.n536 B.n535 10.6151
R1172 B.n535 B.n532 10.6151
R1173 B.n532 B.n531 10.6151
R1174 B.n531 B.n528 10.6151
R1175 B.n528 B.n527 10.6151
R1176 B.n527 B.n524 10.6151
R1177 B.n524 B.n523 10.6151
R1178 B.n523 B.n520 10.6151
R1179 B.n520 B.n519 10.6151
R1180 B.n519 B.n516 10.6151
R1181 B.n516 B.n515 10.6151
R1182 B.n515 B.n512 10.6151
R1183 B.n512 B.n511 10.6151
R1184 B.n511 B.n508 10.6151
R1185 B.n508 B.n507 10.6151
R1186 B.n507 B.n504 10.6151
R1187 B.n504 B.n503 10.6151
R1188 B.n503 B.n500 10.6151
R1189 B.n500 B.n499 10.6151
R1190 B.n499 B.n496 10.6151
R1191 B.n496 B.n495 10.6151
R1192 B.n495 B.n492 10.6151
R1193 B.n492 B.n491 10.6151
R1194 B.n491 B.n488 10.6151
R1195 B.n488 B.n487 10.6151
R1196 B.n487 B.n484 10.6151
R1197 B.n484 B.n483 10.6151
R1198 B.n483 B.n480 10.6151
R1199 B.n480 B.n479 10.6151
R1200 B.n479 B.n476 10.6151
R1201 B.n476 B.n475 10.6151
R1202 B.n472 B.n471 10.6151
R1203 B.n471 B.n468 10.6151
R1204 B.n468 B.n467 10.6151
R1205 B.n467 B.n464 10.6151
R1206 B.n464 B.n463 10.6151
R1207 B.n463 B.n460 10.6151
R1208 B.n460 B.n459 10.6151
R1209 B.n459 B.n456 10.6151
R1210 B.n454 B.n451 10.6151
R1211 B.n451 B.n450 10.6151
R1212 B.n450 B.n447 10.6151
R1213 B.n447 B.n446 10.6151
R1214 B.n446 B.n443 10.6151
R1215 B.n443 B.n442 10.6151
R1216 B.n442 B.n439 10.6151
R1217 B.n439 B.n438 10.6151
R1218 B.n438 B.n435 10.6151
R1219 B.n435 B.n434 10.6151
R1220 B.n434 B.n431 10.6151
R1221 B.n431 B.n430 10.6151
R1222 B.n430 B.n427 10.6151
R1223 B.n427 B.n426 10.6151
R1224 B.n426 B.n423 10.6151
R1225 B.n423 B.n422 10.6151
R1226 B.n422 B.n419 10.6151
R1227 B.n419 B.n418 10.6151
R1228 B.n418 B.n415 10.6151
R1229 B.n415 B.n414 10.6151
R1230 B.n414 B.n411 10.6151
R1231 B.n411 B.n410 10.6151
R1232 B.n410 B.n407 10.6151
R1233 B.n407 B.n406 10.6151
R1234 B.n406 B.n403 10.6151
R1235 B.n403 B.n402 10.6151
R1236 B.n402 B.n399 10.6151
R1237 B.n399 B.n398 10.6151
R1238 B.n398 B.n395 10.6151
R1239 B.n395 B.n394 10.6151
R1240 B.n394 B.n391 10.6151
R1241 B.n391 B.n390 10.6151
R1242 B.n390 B.n387 10.6151
R1243 B.n387 B.n386 10.6151
R1244 B.n386 B.n383 10.6151
R1245 B.n383 B.n382 10.6151
R1246 B.n382 B.n379 10.6151
R1247 B.n379 B.n378 10.6151
R1248 B.n378 B.n325 10.6151
R1249 B.n558 B.n325 10.6151
R1250 B.n564 B.n321 10.6151
R1251 B.n565 B.n564 10.6151
R1252 B.n566 B.n565 10.6151
R1253 B.n566 B.n313 10.6151
R1254 B.n576 B.n313 10.6151
R1255 B.n577 B.n576 10.6151
R1256 B.n578 B.n577 10.6151
R1257 B.n578 B.n305 10.6151
R1258 B.n589 B.n305 10.6151
R1259 B.n590 B.n589 10.6151
R1260 B.n591 B.n590 10.6151
R1261 B.n591 B.n298 10.6151
R1262 B.n601 B.n298 10.6151
R1263 B.n602 B.n601 10.6151
R1264 B.n603 B.n602 10.6151
R1265 B.n603 B.n290 10.6151
R1266 B.n613 B.n290 10.6151
R1267 B.n614 B.n613 10.6151
R1268 B.n615 B.n614 10.6151
R1269 B.n615 B.n282 10.6151
R1270 B.n626 B.n282 10.6151
R1271 B.n627 B.n626 10.6151
R1272 B.n628 B.n627 10.6151
R1273 B.n628 B.n0 10.6151
R1274 B.n714 B.n1 10.6151
R1275 B.n714 B.n713 10.6151
R1276 B.n713 B.n712 10.6151
R1277 B.n712 B.n9 10.6151
R1278 B.n706 B.n9 10.6151
R1279 B.n706 B.n705 10.6151
R1280 B.n705 B.n704 10.6151
R1281 B.n704 B.n16 10.6151
R1282 B.n698 B.n16 10.6151
R1283 B.n698 B.n697 10.6151
R1284 B.n697 B.n696 10.6151
R1285 B.n696 B.n23 10.6151
R1286 B.n690 B.n23 10.6151
R1287 B.n690 B.n689 10.6151
R1288 B.n689 B.n688 10.6151
R1289 B.n688 B.n29 10.6151
R1290 B.n682 B.n29 10.6151
R1291 B.n682 B.n681 10.6151
R1292 B.n681 B.n680 10.6151
R1293 B.n680 B.n37 10.6151
R1294 B.n674 B.n37 10.6151
R1295 B.n674 B.n673 10.6151
R1296 B.n673 B.n672 10.6151
R1297 B.n672 B.n44 10.6151
R1298 B.n617 B.t6 9.08337
R1299 B.t21 B.n708 9.08337
R1300 B.n574 B.t8 7.78581
R1301 B.n593 B.t5 7.78581
R1302 B.n692 B.t23 7.78581
R1303 B.n678 B.t15 7.78581
R1304 B.n182 B.n181 6.5566
R1305 B.n198 B.n96 6.5566
R1306 B.n472 B.n374 6.5566
R1307 B.n456 B.n455 6.5566
R1308 B.n181 B.n180 4.05904
R1309 B.n201 B.n96 4.05904
R1310 B.n475 B.n374 4.05904
R1311 B.n455 B.n454 4.05904
R1312 B.n720 B.n0 2.81026
R1313 B.n720 B.n1 2.81026
R1314 VP.n4 VP.t3 544.194
R1315 VP.n10 VP.t7 517.374
R1316 VP.n1 VP.t6 517.374
R1317 VP.n14 VP.t5 517.374
R1318 VP.n15 VP.t4 517.374
R1319 VP.n16 VP.t1 517.374
R1320 VP.n8 VP.t9 517.374
R1321 VP.n7 VP.t2 517.374
R1322 VP.n6 VP.t8 517.374
R1323 VP.n5 VP.t0 517.374
R1324 VP.n17 VP.n16 161.3
R1325 VP.n9 VP.n8 161.3
R1326 VP.n11 VP.n10 161.3
R1327 VP.n6 VP.n3 80.6037
R1328 VP.n7 VP.n2 80.6037
R1329 VP.n15 VP.n0 80.6037
R1330 VP.n14 VP.n13 80.6037
R1331 VP.n12 VP.n1 80.6037
R1332 VP.n10 VP.n1 48.2005
R1333 VP.n14 VP.n1 48.2005
R1334 VP.n15 VP.n14 48.2005
R1335 VP.n16 VP.n15 48.2005
R1336 VP.n8 VP.n7 48.2005
R1337 VP.n7 VP.n6 48.2005
R1338 VP.n6 VP.n5 48.2005
R1339 VP.n4 VP.n3 45.2318
R1340 VP.n11 VP.n9 42.1558
R1341 VP.n5 VP.n4 13.3799
R1342 VP.n3 VP.n2 0.380177
R1343 VP.n13 VP.n12 0.380177
R1344 VP.n13 VP.n0 0.380177
R1345 VP.n9 VP.n2 0.285035
R1346 VP.n12 VP.n11 0.285035
R1347 VP.n17 VP.n0 0.285035
R1348 VP VP.n17 0.0516364
R1349 VDD1.n1 VDD1.t6 62.9427
R1350 VDD1.n3 VDD1.t2 62.9425
R1351 VDD1.n5 VDD1.n4 60.9872
R1352 VDD1.n1 VDD1.n0 60.4285
R1353 VDD1.n7 VDD1.n6 60.4283
R1354 VDD1.n3 VDD1.n2 60.4283
R1355 VDD1.n7 VDD1.n5 38.6668
R1356 VDD1.n6 VDD1.t7 1.69571
R1357 VDD1.n6 VDD1.t0 1.69571
R1358 VDD1.n0 VDD1.t9 1.69571
R1359 VDD1.n0 VDD1.t1 1.69571
R1360 VDD1.n4 VDD1.t5 1.69571
R1361 VDD1.n4 VDD1.t8 1.69571
R1362 VDD1.n2 VDD1.t3 1.69571
R1363 VDD1.n2 VDD1.t4 1.69571
R1364 VDD1 VDD1.n7 0.556535
R1365 VDD1 VDD1.n1 0.263431
R1366 VDD1.n5 VDD1.n3 0.149895
C0 VDD2 VDD1 0.923394f
C1 VP VTAIL 5.92042f
C2 VDD1 VTAIL 14.6616f
C3 VP VDD1 6.27791f
C4 VDD2 VN 6.10006f
C5 VN VTAIL 5.9058f
C6 VDD2 VTAIL 14.6951f
C7 VP VN 5.41586f
C8 VN VDD1 0.149293f
C9 VDD2 VP 0.33182f
C10 VDD2 B 4.833187f
C11 VDD1 B 4.747552f
C12 VTAIL B 6.324971f
C13 VN B 9.06921f
C14 VP B 7.085616f
C15 VDD1.t6 B 2.63258f
C16 VDD1.t9 B 0.232042f
C17 VDD1.t1 B 0.232042f
C18 VDD1.n0 B 2.06236f
C19 VDD1.n1 B 0.645778f
C20 VDD1.t2 B 2.63258f
C21 VDD1.t3 B 0.232042f
C22 VDD1.t4 B 0.232042f
C23 VDD1.n2 B 2.06235f
C24 VDD1.n3 B 0.640491f
C25 VDD1.t5 B 0.232042f
C26 VDD1.t8 B 0.232042f
C27 VDD1.n4 B 2.0654f
C28 VDD1.n5 B 1.92915f
C29 VDD1.t7 B 0.232042f
C30 VDD1.t0 B 0.232042f
C31 VDD1.n6 B 2.06235f
C32 VDD1.n7 B 2.34429f
C33 VP.n0 B 0.07525f
C34 VP.t6 B 0.933346f
C35 VP.n1 B 0.386045f
C36 VP.n2 B 0.07525f
C37 VP.t9 B 0.933346f
C38 VP.t2 B 0.933346f
C39 VP.t8 B 0.933346f
C40 VP.n3 B 0.236228f
C41 VP.t0 B 0.933346f
C42 VP.t3 B 0.951874f
C43 VP.n4 B 0.358627f
C44 VP.n5 B 0.386045f
C45 VP.n6 B 0.386045f
C46 VP.n7 B 0.386045f
C47 VP.n8 B 0.375793f
C48 VP.n9 B 1.89139f
C49 VP.t7 B 0.933346f
C50 VP.n10 B 0.375793f
C51 VP.n11 B 1.93003f
C52 VP.n12 B 0.07525f
C53 VP.n13 B 0.090356f
C54 VP.t5 B 0.933346f
C55 VP.n14 B 0.386045f
C56 VP.t4 B 0.933346f
C57 VP.n15 B 0.386045f
C58 VP.t1 B 0.933346f
C59 VP.n16 B 0.375793f
C60 VP.n17 B 0.050118f
C61 VTAIL.t10 B 0.242214f
C62 VTAIL.t9 B 0.242214f
C63 VTAIL.n0 B 2.07129f
C64 VTAIL.n1 B 0.395736f
C65 VTAIL.t19 B 2.639f
C66 VTAIL.n2 B 0.501f
C67 VTAIL.t1 B 0.242214f
C68 VTAIL.t6 B 0.242214f
C69 VTAIL.n3 B 2.07129f
C70 VTAIL.n4 B 0.403025f
C71 VTAIL.t5 B 0.242214f
C72 VTAIL.t2 B 0.242214f
C73 VTAIL.n5 B 2.07129f
C74 VTAIL.n6 B 1.68017f
C75 VTAIL.t14 B 0.242214f
C76 VTAIL.t12 B 0.242214f
C77 VTAIL.n7 B 2.07129f
C78 VTAIL.n8 B 1.68016f
C79 VTAIL.t8 B 0.242214f
C80 VTAIL.t13 B 0.242214f
C81 VTAIL.n9 B 2.07129f
C82 VTAIL.n10 B 0.403018f
C83 VTAIL.t11 B 2.63901f
C84 VTAIL.n11 B 0.500993f
C85 VTAIL.t3 B 0.242214f
C86 VTAIL.t18 B 0.242214f
C87 VTAIL.n12 B 2.07129f
C88 VTAIL.n13 B 0.408121f
C89 VTAIL.t0 B 0.242214f
C90 VTAIL.t4 B 0.242214f
C91 VTAIL.n14 B 2.07129f
C92 VTAIL.n15 B 0.403018f
C93 VTAIL.t17 B 2.639f
C94 VTAIL.n16 B 1.70379f
C95 VTAIL.t15 B 2.639f
C96 VTAIL.n17 B 1.70379f
C97 VTAIL.t7 B 0.242214f
C98 VTAIL.t16 B 0.242214f
C99 VTAIL.n18 B 2.07129f
C100 VTAIL.n19 B 0.346167f
C101 VDD2.t3 B 2.61908f
C102 VDD2.t7 B 0.230852f
C103 VDD2.t2 B 0.230852f
C104 VDD2.n0 B 2.05178f
C105 VDD2.n1 B 0.637209f
C106 VDD2.t9 B 0.230852f
C107 VDD2.t5 B 0.230852f
C108 VDD2.n2 B 2.05481f
C109 VDD2.n3 B 1.84419f
C110 VDD2.t8 B 2.61452f
C111 VDD2.n4 B 2.33702f
C112 VDD2.t1 B 0.230852f
C113 VDD2.t4 B 0.230852f
C114 VDD2.n5 B 2.05179f
C115 VDD2.n6 B 0.295644f
C116 VDD2.t0 B 0.230852f
C117 VDD2.t6 B 0.230852f
C118 VDD2.n7 B 2.05478f
C119 VN.n0 B 0.074127f
C120 VN.t7 B 0.919422f
C121 VN.n1 B 0.380285f
C122 VN.t6 B 0.937673f
C123 VN.n2 B 0.353277f
C124 VN.n3 B 0.232704f
C125 VN.t9 B 0.919422f
C126 VN.n4 B 0.380285f
C127 VN.t0 B 0.919422f
C128 VN.n5 B 0.380285f
C129 VN.t1 B 0.919422f
C130 VN.n6 B 0.370187f
C131 VN.n7 B 0.04937f
C132 VN.n8 B 0.074127f
C133 VN.t3 B 0.919422f
C134 VN.n9 B 0.380285f
C135 VN.t8 B 0.919422f
C136 VN.t5 B 0.937673f
C137 VN.n10 B 0.353277f
C138 VN.n11 B 0.232704f
C139 VN.n12 B 0.380285f
C140 VN.t4 B 0.919422f
C141 VN.n13 B 0.380285f
C142 VN.t2 B 0.919422f
C143 VN.n14 B 0.370187f
C144 VN.n15 B 1.89239f
.ends

