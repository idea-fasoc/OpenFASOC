* File: sky130_osu_sc_12T_hs__addf_1.spice
* Created: Mon Nov 16 20:37:05 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__addf_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__addf_1  GND VDD A B CI CON S CO
*
* CO	CO
* S	S
* CON	CON
* CI	CI
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1013 N_GND_M1013_d N_A_M1013_g N_A_27_115#_M1013_s N_GND_M1013_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75005.3 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_115#_M1001_d N_B_M1001_g N_GND_M1013_d N_GND_M1013_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1003 N_CON_M1003_d N_CI_M1003_g N_A_27_115#_M1001_d N_GND_M1013_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75004.4 A=0.0825 P=1.4 MULT=1
MM1025 A_368_115# N_B_M1025_g N_CON_M1003_d N_GND_M1013_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75004 A=0.0825 P=1.4 MULT=1
MM1027 N_GND_M1027_d N_A_M1027_g A_368_115# N_GND_M1013_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.8
+ SB=75003.6 A=0.0825 P=1.4 MULT=1
MM1022 N_A_526_115#_M1022_d N_A_M1022_g N_GND_M1027_d N_GND_M1013_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.3 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1024 N_GND_M1024_d N_B_M1024_g N_A_526_115#_M1022_d N_GND_M1013_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.7 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1014 N_A_526_115#_M1014_d N_CI_M1014_g N_GND_M1024_d N_GND_M1013_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.1 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1015 N_A_784_115#_M1015_d N_CON_M1015_g N_A_526_115#_M1014_d N_GND_M1013_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75003.6 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1017 A_870_115# N_B_M1017_g N_A_784_115#_M1015_d N_GND_M1013_b NLOWVT L=0.15
+ W=0.55 AD=0.0715 AS=0.077 PD=0.81 PS=0.83 NRD=16.356 NRS=0 M=1 R=3.66667
+ SA=75004 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1008 A_952_115# N_CI_M1008_g A_870_115# N_GND_M1013_b NLOWVT L=0.15 W=0.55
+ AD=0.0715 AS=0.0715 PD=0.81 PS=0.81 NRD=16.356 NRS=16.356 M=1 R=3.66667
+ SA=75004.4 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1004_d N_A_M1004_g A_952_115# N_GND_M1013_b NLOWVT L=0.15 W=0.55
+ AD=0.0935 AS=0.0715 PD=0.89 PS=0.81 NRD=0 NRS=16.356 M=1 R=3.66667 SA=75004.8
+ SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1018 N_S_M1018_d N_A_784_115#_M1018_g N_GND_M1004_d N_GND_M1013_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.0935 PD=1.63 PS=0.89 NRD=0 NRS=13.08 M=1
+ R=3.66667 SA=75005.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1023 N_CO_M1023_d N_CON_M1023_g N_GND_M1023_s N_GND_M1013_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1019 N_A_27_521#_M1019_d N_B_M1019_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1020 N_CON_M1020_d N_CI_M1020_g N_A_27_521#_M1019_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75004.4 A=0.189 P=2.82 MULT=1
MM1012 A_368_521# N_B_M1012_g N_CON_M1020_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004 A=0.189 P=2.82 MULT=1
MM1016 N_VDD_M1016_d N_A_M1016_g A_368_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.8
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1009 N_A_526_521#_M1009_d N_A_M1009_g N_VDD_M1016_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1011 N_VDD_M1011_d N_B_M1011_g N_A_526_521#_M1009_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.7 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1002 N_A_526_521#_M1002_d N_CI_M1002_g N_VDD_M1011_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.1 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 N_A_784_115#_M1005_d N_CON_M1005_g N_A_526_521#_M1002_d N_VDD_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 A_870_521# N_B_M1006_g N_A_784_115#_M1005_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1638 AS=0.1764 PD=1.52 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4
+ SA=75004 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1026 A_952_521# N_CI_M1026_g A_870_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1638 AS=0.1638 PD=1.52 PS=1.52 NRD=11.7215 NRS=11.7215 M=1 R=8.4
+ SA=75004.4 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_VDD_M1021_d N_A_M1021_g A_952_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.2142 AS=0.1638 PD=1.6 PS=1.52 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75004.8
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 N_S_M1007_d N_A_784_115#_M1007_g N_VDD_M1021_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.2142 PD=3.05 PS=1.6 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75005.3 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1010 N_CO_M1010_d N_CON_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref N_GND_M1013_b N_VDD_M1000_b NWDIODE A=14.8732 P=18.56
pX29_noxref noxref_20 A A PROBETYPE=1
pX30_noxref noxref_21 B B PROBETYPE=1
pX31_noxref noxref_22 CI CI PROBETYPE=1
pX32_noxref noxref_23 S S PROBETYPE=1
pX33_noxref noxref_24 CON CON PROBETYPE=1
pX34_noxref noxref_25 CO CO PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__addf_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__addf_l.spice
* Created: Mon Nov 16 20:37:11 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__addf_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__addf_l  GND VDD A B CI CON S CO
*
* CO	CO
* S	S
* CON	CON
* CI	CI
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1012 N_GND_M1012_d N_A_M1012_g N_A_27_115#_M1012_s N_GND_M1012_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75005.3 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_115#_M1001_d N_B_M1001_g N_GND_M1012_d N_GND_M1012_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75004.9 A=0.0825 P=1.4 MULT=1
MM1003 N_CON_M1003_d N_CI_M1003_g N_A_27_115#_M1001_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75004.4 A=0.0825 P=1.4 MULT=1
MM1025 A_368_115# N_B_M1025_g N_CON_M1003_d N_GND_M1012_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75004 A=0.0825 P=1.4 MULT=1
MM1027 N_GND_M1027_d N_A_M1027_g A_368_115# N_GND_M1012_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.8
+ SB=75003.6 A=0.0825 P=1.4 MULT=1
MM1022 N_A_526_115#_M1022_d N_A_M1022_g N_GND_M1027_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.3 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1024 N_GND_M1024_d N_B_M1024_g N_A_526_115#_M1022_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.7 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1013 N_A_526_115#_M1013_d N_CI_M1013_g N_GND_M1024_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.1 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1014 N_A_784_115#_M1014_d N_CON_M1014_g N_A_526_115#_M1013_d N_GND_M1012_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75003.6 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1016 A_870_115# N_B_M1016_g N_A_784_115#_M1014_d N_GND_M1012_b NLOWVT L=0.15
+ W=0.55 AD=0.0715 AS=0.077 PD=0.81 PS=0.83 NRD=16.356 NRS=0 M=1 R=3.66667
+ SA=75004 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1008 A_952_115# N_CI_M1008_g A_870_115# N_GND_M1012_b NLOWVT L=0.15 W=0.55
+ AD=0.0715 AS=0.0715 PD=0.81 PS=0.81 NRD=16.356 NRS=16.356 M=1 R=3.66667
+ SA=75004.4 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1004_d N_A_M1004_g A_952_115# N_GND_M1012_b NLOWVT L=0.15 W=0.55
+ AD=0.0935 AS=0.0715 PD=0.89 PS=0.81 NRD=0 NRS=16.356 M=1 R=3.66667 SA=75004.8
+ SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1017 N_S_M1017_d N_A_784_115#_M1017_g N_GND_M1004_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.0935 PD=1.63 PS=0.89 NRD=0 NRS=13.08 M=1
+ R=3.66667 SA=75005.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1023 N_CO_M1023_d N_CON_M1023_g N_GND_M1023_s N_GND_M1012_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1019 N_A_27_521#_M1019_d N_B_M1019_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.9 A=0.189 P=2.82 MULT=1
MM1020 N_CON_M1020_d N_CI_M1020_g N_A_27_521#_M1019_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75004.4 A=0.189 P=2.82 MULT=1
MM1011 A_368_521# N_B_M1011_g N_CON_M1020_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75004 A=0.189 P=2.82 MULT=1
MM1015 N_VDD_M1015_d N_A_M1015_g A_368_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.8
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1009 N_A_526_521#_M1009_d N_A_M1009_g N_VDD_M1015_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1010 N_VDD_M1010_d N_B_M1010_g N_A_526_521#_M1009_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.7 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1002 N_A_526_521#_M1002_d N_CI_M1002_g N_VDD_M1010_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.1 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1005 N_A_784_115#_M1005_d N_CON_M1005_g N_A_526_521#_M1002_d N_VDD_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 A_870_521# N_B_M1006_g N_A_784_115#_M1005_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1638 AS=0.1764 PD=1.52 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4
+ SA=75004 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1026 A_952_521# N_CI_M1026_g A_870_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1638 AS=0.1638 PD=1.52 PS=1.52 NRD=11.7215 NRS=11.7215 M=1 R=8.4
+ SA=75004.4 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_VDD_M1021_d N_A_M1021_g A_952_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.2142 AS=0.1638 PD=1.6 PS=1.52 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75004.8
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 N_S_M1007_d N_A_784_115#_M1007_g N_VDD_M1021_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.2142 PD=3.05 PS=1.6 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75005.3 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1018 N_CO_M1018_d N_CON_M1018_g N_VDD_M1018_s N_VDD_M1000_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX28_noxref N_GND_M1012_b N_VDD_M1000_b NWDIODE A=14.8732 P=18.56
pX29_noxref noxref_20 A A PROBETYPE=1
pX30_noxref noxref_21 B B PROBETYPE=1
pX31_noxref noxref_22 CI CI PROBETYPE=1
pX32_noxref noxref_23 S S PROBETYPE=1
pX33_noxref noxref_24 CON CON PROBETYPE=1
pX34_noxref noxref_25 CO CO PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__addf_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__addh_1.spice
* Created: Mon Nov 16 20:37:17 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__addh_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__addh_1  GND VDD CON B A S CO
*
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1007 N_GND_M1007_d N_CON_M1007_g N_S_M1007_s N_GND_M1007_b NSHORT L=0.15
+ W=0.55 AD=0.0935 AS=0.14575 PD=0.89 PS=1.63 NRD=13.08 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1008 A_208_115# N_B_M1008_g N_GND_M1007_d N_GND_M1007_b NSHORT L=0.15 W=0.55
+ AD=0.05775 AS=0.0935 PD=0.76 PS=0.89 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.7
+ SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1010 N_A_208_521#_M1010_d N_A_M1010_g A_208_115# N_GND_M1007_b NSHORT L=0.15
+ W=0.55 AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_208_521#_M1002_g N_CO_M1002_s N_GND_M1007_b NSHORT
+ L=0.15 W=0.55 AD=0.0935 AS=0.14575 PD=0.89 PS=1.63 NRD=13.08 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1011 N_CON_M1011_d N_A_208_521#_M1011_g N_GND_M1002_d N_GND_M1007_b NSHORT
+ L=0.15 W=0.55 AD=0.077 AS=0.0935 PD=0.83 PS=0.89 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.7 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1004 N_CON_M1011_d N_B_M1004_g N_CON_M1011_d N_GND_M1007_b NSHORT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1005 N_CON_M1011_d N_A_M1005_g N_CON_M1011_d N_GND_M1007_b NSHORT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_CON_M1000_g N_S_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.2142 AS=0.3339 PD=1.6 PS=3.05 NRD=9.3772 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_208_521#_M1001_d N_B_M1001_g N_VDD_M1000_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.2142 PD=1.54 PS=1.6 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g N_A_208_521#_M1001_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.2142 AS=0.1764 PD=1.6 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1012 N_CO_M1012_d N_A_208_521#_M1012_g N_VDD_M1003_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.2142 PD=3.05 PS=1.6 NRD=0 NRS=9.3772 M=1 R=8.4
+ SA=75001.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1013_d N_A_208_521#_M1013_g N_CON_M1013_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1006 A_668_521# N_B_M1006_g N_VDD_M1013_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_CON_M1009_d N_A_M1009_g A_668_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3528 AS=0.1323 PD=3.08 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref N_GND_M1007_b N_VDD_M1000_b NWDIODE A=8.7138 P=12.58
pX15_noxref noxref_11 S S PROBETYPE=1
pX16_noxref noxref_12 CO CO PROBETYPE=1
pX17_noxref noxref_13 B B PROBETYPE=1
pX18_noxref noxref_14 CON CON PROBETYPE=1
pX19_noxref noxref_15 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__addh_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__addh_l.spice
* Created: Mon Nov 16 20:37:22 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__addh_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__addh_l  GND VDD CON B A S CO
*
* CO	CO
* S	S
* A	A
* B	B
* CON	CON
* VDD	VDD
* GND	GND
MM1007 N_GND_M1007_d N_CON_M1007_g N_S_M1007_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.42 AD=0.0767474 AS=0.1113 PD=0.770722 PS=1.37 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1009 A_208_115# N_B_M1009_g N_GND_M1007_d N_GND_M1007_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.100503 PD=0.76 PS=1.00928 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1010 N_A_208_521#_M1010_d N_A_M1010_g A_208_115# N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.9 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_208_521#_M1002_g N_CO_M1002_s N_GND_M1007_b NLOWVT
+ L=0.15 W=0.42 AD=0.0767474 AS=0.1113 PD=0.770722 PS=1.37 NRD=17.136 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1011 N_CON_M1011_d N_A_208_521#_M1011_g N_GND_M1002_d N_GND_M1007_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.100503 PD=0.83 PS=1.00928 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1004 N_CON_M1011_d N_B_M1004_g N_CON_M1011_d N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1005 N_CON_M1011_d N_A_M1005_g N_CON_M1011_d N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.4 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_VDD_M1003_d N_CON_M1003_g N_S_M1003_s N_VDD_M1003_b PSHORT L=0.15
+ W=0.835 AD=0.158042 AS=0.221275 PD=1.27542 PS=2.2 NRD=14.5386 NRS=0 M=1
+ R=5.56667 SA=75000.2 SB=75001.6 A=0.12525 P=1.97 MULT=1
MM1000 N_A_208_521#_M1000_d N_B_M1000_g N_VDD_M1003_d N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.238483 PD=1.54 PS=1.92458 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_208_521#_M1000_d N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.23814 AS=0.1764 PD=1.92 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.9 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1013 N_CO_M1013_d N_A_208_521#_M1013_g N_VDD_M1001_d N_VDD_M1003_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.15876 PD=2.21 PS=1.28 NRD=0 NRS=14.0658 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_VDD_M1012_d N_A_208_521#_M1012_g N_CON_M1012_s N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1006 A_668_521# N_B_M1006_g N_VDD_M1012_d N_VDD_M1003_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_CON_M1008_d N_A_M1008_g A_668_521# N_VDD_M1003_b PSHORT L=0.15 W=1.26
+ AD=0.3528 AS=0.1323 PD=3.08 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref N_GND_M1007_b N_VDD_M1003_b NWDIODE A=8.7138 P=12.58
pX15_noxref noxref_11 S S PROBETYPE=1
pX16_noxref noxref_12 CO CO PROBETYPE=1
pX17_noxref noxref_13 B B PROBETYPE=1
pX18_noxref noxref_14 CON CON PROBETYPE=1
pX19_noxref noxref_15 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__addh_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_1.spice
* Created: Mon Nov 16 20:37:28 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_1  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.09625 PD=1.63 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B_M1004_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_2.spice
* Created: Mon Nov 16 20:37:34 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_2.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_2  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_Y_M1001_d N_A_27_115#_M1007_g N_GND_M1007_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_B_M1005_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1005_d N_A_27_115#_M1003_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_27_115#_M1006_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=4.8513 P=8.83
pX9_noxref noxref_8 A A PROBETYPE=1
pX10_noxref noxref_9 B B PROBETYPE=1
pX11_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_2.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_4.spice
* Created: Mon Nov 16 20:37:39 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_4.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_4  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_B_M1002_g A_110_115# N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75002 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1001_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1010 N_Y_M1010_d N_A_27_115#_M1010_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1010_d N_A_27_115#_M1011_g N_GND_M1011_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_B_M1007_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1007_d N_A_27_115#_M1003_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_27_115#_M1005_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1005_d N_A_27_115#_M1006_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VDD_M1008_d N_A_27_115#_M1008_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_8 A A PROBETYPE=1
pX14_noxref noxref_9 B B PROBETYPE=1
pX15_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_4.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_6.spice
* Created: Mon Nov 16 20:37:45 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_6.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_6  A B Y GND VDD
*
* Y	Y
* B	B
* A	A
MM1006 A_110_115# N_A_M1006_g N_A_27_115#_M1006_s N_noxref_1_M1006_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1002 N_noxref_1_M1002_d N_B_M1002_g A_110_115# N_noxref_1_M1006_b NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_noxref_1_M1002_d N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1
+ R=3.66667 SA=75001.1 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1001_d N_A_27_115#_M1011_g N_noxref_1_M1011_s N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75001.5 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1012 N_Y_M1012_d N_A_27_115#_M1012_g N_noxref_1_M1011_s N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1013 N_Y_M1012_d N_A_27_115#_M1013_g N_noxref_1_M1013_s N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1014 N_Y_M1014_d N_A_27_115#_M1014_g N_noxref_1_M1013_s N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75002.8 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1015 N_Y_M1014_d N_A_27_115#_M1015_g N_noxref_1_M1015_s N_noxref_1_M1006_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75003.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_noxref_2_M1000_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75003.2 A=0.189 P=2.82 MULT=1
MM1009 N_noxref_2_M1009_d N_B_M1009_g N_A_27_115#_M1000_d N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_noxref_2_M1009_d N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1003_d N_A_27_115#_M1004_g N_noxref_2_M1004_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_noxref_2_M1004_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1005_d N_A_27_115#_M1007_g N_noxref_2_M1007_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1008_d N_A_27_115#_M1008_g N_noxref_2_M1007_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1008_d N_A_27_115#_M1010_g N_noxref_2_M1010_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref N_noxref_1_M1006_b N_noxref_2_M1000_b NWDIODE A=8.4769 P=12.35
pX17_noxref noxref_10 A A PROBETYPE=1
pX18_noxref noxref_11 B B PROBETYPE=1
pX19_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_6.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_8.spice
* Created: Mon Nov 16 20:37:51 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_8  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1008 A_110_115# N_A_M1008_g N_A_27_115#_M1008_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1004_d N_B_M1004_g A_110_115# N_GND_M1008_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75000.5
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_GND_M1004_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.09625 PD=0.83 PS=0.9 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75001.1 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1003_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1012 N_Y_M1012_d N_A_27_115#_M1012_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1015 N_Y_M1012_d N_A_27_115#_M1015_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1016 N_Y_M1016_d N_A_27_115#_M1016_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1017 N_Y_M1016_d N_A_27_115#_M1017_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1018 N_Y_M1018_d N_A_27_115#_M1018_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1019 N_Y_M1018_d N_A_27_115#_M1019_g N_GND_M1019_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_27_115#_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1013_d N_B_M1013_g N_A_27_115#_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_VDD_M1013_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1001_d N_A_27_115#_M1002_g N_VDD_M1002_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1002_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_27_115#_M1006_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_27_115#_M1007_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1007_d N_A_27_115#_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A_27_115#_M1011_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1011_d N_A_27_115#_M1014_g N_VDD_M1014_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref N_GND_M1008_b N_VDD_M1000_b NWDIODE A=10.2897 P=14.11
pX21_noxref noxref_8 A A PROBETYPE=1
pX22_noxref noxref_9 B B PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_8.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__and2_l.spice
* Created: Mon Nov 16 20:37:56 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__and2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__and2_l  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1003 A_110_115# N_A_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1003_b NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1001_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0735 PD=1.37 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_27_115#_M1002_d N_A_M1002_g N_VDD_M1002_s N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_VDD_M1004_d N_B_M1004_g N_A_27_115#_M1002_d N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_27_115#_M1005_g N_VDD_M1004_d N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=3.23635 P=7.21
pX7_noxref noxref_8 A A PROBETYPE=1
pX8_noxref noxref_9 B B PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__and2_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__ant.spice
* Created: Mon Nov 16 20:38:05 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__ant.pex.spice"
.subckt sky130_osu_sc_12T_hs__ant  GND VDD A
*
* A	A
* VDD	VDD
* GND	GND
MM1001 N_A_M1001_s N_A_M1001_g N_A_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.1424 P=6.2
pX3_noxref noxref_4 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__ant.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__aoi21_l.spice
* Created: Mon Nov 16 20:38:11 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__aoi21_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__aoi21_l  GND VDD A0 A1 B0 Y
*
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1002 A_110_114# N_A0_M1002_g N_GND_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_110_114# N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.0997655 AS=0.05775 PD=1.00928 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.5 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1003 N_GND_M1003_d N_B0_M1003_g N_Y_M1001_d N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0761845 PD=1.37 PS=0.770722 NRD=0 NRS=17.136 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VDD_M1000_d N_A0_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_27_521#_M1004_d N_A1_M1004_g N_VDD_M1000_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_B0_M1005_g N_A_27_521#_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=3.9552 P=7.96
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__aoi21_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__aoi22_l.spice
* Created: Mon Nov 16 20:38:16 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__aoi22_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__aoi22_l  GND VDD A0 A1 B0 B1 Y
*
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1004 A_110_115# N_A0_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A1_M1002_g A_110_115# N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.09625 AS=0.05775 PD=0.9 PS=0.76 NRD=7.632 NRS=10.908 M=1 R=3.66667
+ SA=75000.5 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 A_282_115# N_B0_M1001_g N_Y_M1002_d N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.09625 PD=0.76 PS=0.9 NRD=10.908 NRS=7.632 M=1 R=3.66667
+ SA=75001.1 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1007 N_GND_M1007_d N_B1_M1007_g A_282_115# N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.4 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A0_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_A_27_521#_M1005_d N_A1_M1005_g N_VDD_M1000_d N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_B0_M1006_g N_A_27_521#_M1005_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_A_27_521#_M1003_d N_B1_M1003_g N_Y_M1006_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=4.8513 P=8.83
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__aoi22_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_1.spice
* Created: Mon Nov 16 20:38:22 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_1  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=3.0591 P=7.09
pX5_noxref noxref_6 A A PROBETYPE=1
pX6_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_2.spice
* Created: Mon Nov 16 20:38:28 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_2.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_2  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_A_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1001_d N_A_27_115#_M1002_g N_GND_M1002_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_A_27_115#_M1004_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1004_d N_A_27_115#_M1005_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9655 P=7.97
pX7_noxref noxref_6 A A PROBETYPE=1
pX8_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_2.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_4.spice
* Created: Mon Nov 16 20:38:33 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_4.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_4  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A_M1004_g N_A_27_115#_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_GND_M1004_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1001_d N_A_27_115#_M1002_g N_GND_M1002_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1008 N_Y_M1008_d N_A_27_115#_M1008_g N_GND_M1002_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1008_d N_A_27_115#_M1009_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1003_d N_A_27_115#_M1005_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A_27_115#_M1006_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1006_d N_A_27_115#_M1007_g N_VDD_M1007_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=5.7783 P=9.73
pX11_noxref noxref_6 A A PROBETYPE=1
pX12_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_4.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_6.spice
* Created: Mon Nov 16 20:38:39 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_6.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_6  A Y GND VDD
*
* Y	Y
* A	A
MM1005 N_noxref_1_M1005_d N_A_M1005_g N_A_27_115#_M1005_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1001 N_Y_M1001_d N_A_27_115#_M1001_g N_noxref_1_M1005_d N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1001_d N_A_27_115#_M1002_g N_noxref_1_M1002_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75001.1 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1010 N_Y_M1010_d N_A_27_115#_M1010_g N_noxref_1_M1002_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75001.5 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1010_d N_A_27_115#_M1011_g N_noxref_1_M1011_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1012 N_Y_M1012_d N_A_27_115#_M1012_g N_noxref_1_M1011_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1013 N_Y_M1012_d N_A_27_115#_M1013_g N_noxref_1_M1013_s N_noxref_1_M1005_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75002.8 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_noxref_2_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.8 A=0.189 P=2.82 MULT=1
MM1003 N_noxref_2_M1000_d N_A_27_115#_M1003_g N_Y_M1003_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1004 N_noxref_2_M1004_d N_A_27_115#_M1004_g N_Y_M1003_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 N_noxref_2_M1004_d N_A_27_115#_M1006_g N_Y_M1006_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1007 N_noxref_2_M1007_d N_A_27_115#_M1007_g N_Y_M1006_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_noxref_2_M1007_d N_A_27_115#_M1008_g N_Y_M1008_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_noxref_2_M1009_d N_A_27_115#_M1009_g N_Y_M1008_s N_noxref_2_M1000_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref N_noxref_1_M1005_b N_noxref_2_M1000_b NWDIODE A=7.5911 P=11.49
pX15_noxref noxref_8 A A PROBETYPE=1
pX16_noxref noxref_9 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_6.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_8.spice
* Created: Mon Nov 16 20:38:45 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_8  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1007 N_GND_M1007_d N_A_M1007_g N_A_27_115#_M1007_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_27_115#_M1002_g N_GND_M1007_d N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1003 N_Y_M1002_d N_A_27_115#_M1003_g N_GND_M1003_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1008 N_Y_M1008_d N_A_27_115#_M1008_g N_GND_M1003_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1013 N_Y_M1008_d N_A_27_115#_M1013_g N_GND_M1013_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1014 N_Y_M1014_d N_A_27_115#_M1014_g N_GND_M1013_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1015 N_Y_M1014_d N_A_27_115#_M1015_g N_GND_M1015_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1016 N_Y_M1016_d N_A_27_115#_M1016_g N_GND_M1015_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1017 N_Y_M1016_d N_A_27_115#_M1017_g N_GND_M1017_s N_GND_M1007_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.6 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1001 N_VDD_M1000_d N_A_27_115#_M1001_g N_Y_M1001_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_27_115#_M1004_g N_Y_M1001_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1004_d N_A_27_115#_M1005_g N_Y_M1005_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_27_115#_M1006_g N_Y_M1005_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_VDD_M1006_d N_A_27_115#_M1009_g N_Y_M1009_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_VDD_M1010_d N_A_27_115#_M1010_g N_Y_M1009_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_VDD_M1010_d N_A_27_115#_M1011_g N_Y_M1011_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_VDD_M1012_d N_A_27_115#_M1012_g N_Y_M1011_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref N_GND_M1007_b N_VDD_M1000_b NWDIODE A=9.4039 P=13.25
pX19_noxref noxref_6 A A PROBETYPE=1
pX20_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_8.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__buf_l.spice
* Created: Mon Nov 16 20:38:50 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__buf_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__buf_l  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_27_115#_M1000_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VDD_M1001_d N_A_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_27_115#_M1003_g N_VDD_M1001_d N_VDD_M1001_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=2.50965 P=6.35
pX5_noxref noxref_6 A A PROBETYPE=1
pX6_noxref noxref_7 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__buf_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dff_1.spice
* Created: Mon Nov 16 20:38:58 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dff_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dff_1  GND VDD D CK ON Q
*
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1008 N_GND_M1008_d N_A_75_248#_M1008_g N_A_32_115#_M1008_s N_GND_M1008_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1007 A_201_115# N_D_M1007_g N_GND_M1008_d N_GND_M1008_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1025 N_A_75_248#_M1025_d N_A_243_89#_M1025_g A_201_115# N_GND_M1008_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75001 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1020 A_393_115# N_CK_M1020_g N_A_75_248#_M1025_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.6 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1013 N_GND_M1013_d N_A_32_115#_M1013_g A_393_115# N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.9 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1015 A_551_115# N_A_32_115#_M1015_g N_GND_M1013_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1012 N_A_623_115#_M1012_d N_CK_M1012_g A_551_115# N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1005 A_743_115# N_A_243_89#_M1005_g N_A_623_115#_M1012_d N_GND_M1008_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75003.3 SB=75001 A=0.0825 P=1.4 MULT=1
MM1000 N_GND_M1000_d N_A_785_89#_M1000_g A_743_115# N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75003.7 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1001 N_A_243_89#_M1001_d N_CK_M1001_g N_GND_M1000_d N_GND_M1008_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1009 N_A_785_89#_M1009_d N_A_623_115#_M1009_g N_GND_M1009_s N_GND_M1008_b
+ NLOWVT L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1010 N_GND_M1010_d N_A_785_89#_M1010_g N_ON_M1010_s N_GND_M1008_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Q_M1002_d N_ON_M1002_g N_GND_M1010_d N_GND_M1008_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1022 N_VDD_M1022_d N_A_75_248#_M1022_g N_A_32_115#_M1022_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1021 A_201_521# N_D_M1021_g N_VDD_M1022_d N_VDD_M1022_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1014 N_A_75_248#_M1014_d N_CK_M1014_g A_201_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1011 A_393_521# N_A_243_89#_M1011_g N_A_75_248#_M1014_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_32_115#_M1004_g A_393_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 A_551_521# N_A_32_115#_M1006_g N_VDD_M1004_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_623_115#_M1003_d N_A_243_89#_M1003_g A_551_521# N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.7 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1019 A_743_521# N_CK_M1019_g N_A_623_115#_M1003_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75003.3 SB=75001 A=0.189 P=2.82 MULT=1
MM1016 N_VDD_M1016_d N_A_785_89#_M1016_g A_743_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_243_89#_M1017_d N_CK_M1017_g N_VDD_M1016_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1023 N_A_785_89#_M1023_d N_A_623_115#_M1023_g N_VDD_M1023_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_VDD_M1024_d N_A_785_89#_M1024_g N_ON_M1024_s N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_Q_M1018_d N_ON_M1018_g N_VDD_M1024_d N_VDD_M1022_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1008_b N_VDD_M1022_b NWDIODE A=15.0895 P=18.77
pX27_noxref noxref_20 D D PROBETYPE=1
pX28_noxref noxref_21 CK CK PROBETYPE=1
pX29_noxref noxref_22 ON ON PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
c_1319 A_551_521# 0 1.57671e-19 $X=2.755 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dff_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dff_l.spice
* Created: Mon Nov 16 20:39:04 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dff_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dff_l  GND VDD D CK Q
*
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1009 N_GND_M1009_d N_A_75_248#_M1009_g N_A_32_115#_M1009_s N_GND_M1009_b
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1008 A_201_115# N_D_M1008_g N_GND_M1009_d N_GND_M1009_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1025 N_A_75_248#_M1025_d N_A_243_89#_M1025_g A_201_115# N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75001 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1020 A_393_115# N_CK_M1020_g N_A_75_248#_M1025_d N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.6 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1014 N_GND_M1014_d N_A_32_115#_M1014_g A_393_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.9 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1016 A_551_115# N_A_32_115#_M1016_g N_GND_M1014_d N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1013 N_A_623_115#_M1013_d N_CK_M1013_g A_551_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.7 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1005 A_743_115# N_A_243_89#_M1005_g N_A_623_115#_M1013_d N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75003.3 SB=75001 A=0.0825 P=1.4 MULT=1
MM1000 N_GND_M1000_d N_A_785_89#_M1000_g A_743_115# N_GND_M1009_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75003.7 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1001 N_A_243_89#_M1001_d N_CK_M1001_g N_GND_M1000_d N_GND_M1009_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1010 N_A_785_89#_M1010_d N_A_623_115#_M1010_g N_GND_M1010_s N_GND_M1009_b
+ NLOWVT L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1011 N_GND_M1011_d N_A_785_89#_M1011_g N_ON_M1011_s N_GND_M1009_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_Q_M1002_d N_ON_M1002_g N_GND_M1011_d N_GND_M1009_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1022 N_VDD_M1022_d N_A_75_248#_M1022_g N_A_32_115#_M1022_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1021 A_201_521# N_D_M1021_g N_VDD_M1022_d N_VDD_M1022_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1015 N_A_75_248#_M1015_d N_CK_M1015_g A_201_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1012 A_393_521# N_A_243_89#_M1012_g N_A_75_248#_M1015_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_32_115#_M1004_g A_393_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1006 A_551_521# N_A_32_115#_M1006_g N_VDD_M1004_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_623_115#_M1003_d N_A_243_89#_M1003_g A_551_521# N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.7 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1019 A_743_521# N_CK_M1019_g N_A_623_115#_M1003_d N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75003.3 SB=75001 A=0.189 P=2.82 MULT=1
MM1017 N_VDD_M1017_d N_A_785_89#_M1017_g A_743_521# N_VDD_M1022_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_A_243_89#_M1018_d N_CK_M1018_g N_VDD_M1017_d N_VDD_M1022_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75004.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_A_785_89#_M1024_d N_A_623_115#_M1024_g N_VDD_M1024_s N_VDD_M1022_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_A_785_89#_M1007_g N_ON_M1007_s N_VDD_M1022_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1023 N_Q_M1023_d N_ON_M1023_g N_VDD_M1007_d N_VDD_M1022_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX26_noxref N_GND_M1009_b N_VDD_M1022_b NWDIODE A=15.0895 P=18.77
pX27_noxref noxref_20 D D PROBETYPE=1
pX28_noxref noxref_21 CK CK PROBETYPE=1
* pX29_noxref noxref_22 ON ON PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
c_1323 A_551_521# 0 1.57671e-19 $X=2.755 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dff_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffr_1.spice
* Created: Mon Nov 16 20:39:09 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffr_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffr_1  GND VDD RN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* RN	RN
* VDD	VDD
* GND	GND
MM1020 N_A_110_115#_M1020_d N_RN_M1020_g N_GND_M1020_s N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1016 N_A_217_605#_M1016_d N_A_110_115#_M1016_g N_GND_M1016_s N_GND_M1020_b
+ NLOWVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_GND_M1006_d N_A_342_442#_M1006_g N_A_217_605#_M1016_d N_GND_M1020_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_576_115# N_D_M1007_g N_GND_M1007_s N_GND_M1020_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1031 N_A_342_442#_M1031_d N_A_618_89#_M1031_g A_576_115# N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1024 A_768_115# N_CK_M1024_g N_A_342_442#_M1031_d N_GND_M1020_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1028 N_GND_M1028_d N_A_217_605#_M1028_g A_768_115# N_GND_M1020_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1023 A_926_115# N_A_217_605#_M1023_g N_GND_M1028_d N_GND_M1020_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1017 N_A_998_115#_M1017_d N_CK_M1017_g A_926_115# N_GND_M1020_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1018 A_1118_115# N_A_618_89#_M1018_g N_A_998_115#_M1017_d N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1021 N_GND_M1021_d N_A_1160_89#_M1021_g A_1118_115# N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1009 N_A_618_89#_M1009_d N_CK_M1009_g N_GND_M1021_d N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1011 N_A_1160_89#_M1011_d N_A_998_115#_M1011_g N_GND_M1011_s N_GND_M1020_b
+ NLOWVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_GND_M1013_d N_A_110_115#_M1013_g N_A_1160_89#_M1011_d N_GND_M1020_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_GND_M1015_d N_A_1160_89#_M1015_g N_QN_M1015_s N_GND_M1020_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_GND_M1015_d N_GND_M1020_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_A_110_115#_M1003_d N_RN_M1003_g N_VDD_M1003_s N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1012 A_300_605# N_A_110_115#_M1012_g N_A_217_605#_M1012_s N_VDD_M1003_b PSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_VDD_M1001_d N_A_342_442#_M1001_g A_300_605# N_VDD_M1003_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 A_576_521# N_D_M1026_g N_VDD_M1026_s N_VDD_M1003_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1022 N_A_342_442#_M1022_d N_CK_M1022_g A_576_521# N_VDD_M1003_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1014 A_768_521# N_A_618_89#_M1014_g N_A_342_442#_M1022_d N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1019 N_VDD_M1019_d N_A_217_605#_M1019_g A_768_521# N_VDD_M1003_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1010 A_926_521# N_A_217_605#_M1010_g N_VDD_M1019_d N_VDD_M1003_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1002 N_A_998_115#_M1002_d N_A_618_89#_M1002_g A_926_521# N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 A_1118_521# N_CK_M1000_g N_A_998_115#_M1002_d N_VDD_M1003_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_1160_89#_M1005_g A_1118_521# N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_618_89#_M1027_d N_CK_M1027_g N_VDD_M1005_d N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1004 A_1466_605# N_A_998_115#_M1004_g N_A_1160_89#_M1004_s N_VDD_M1003_b
+ PSHORT L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1029 N_VDD_M1029_d N_A_110_115#_M1029_g A_1466_605# N_VDD_M1003_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1030 N_VDD_M1030_d N_A_1160_89#_M1030_g N_QN_M1030_s N_VDD_M1003_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_Q_M1025_d N_QN_M1025_g N_VDD_M1030_d N_VDD_M1003_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref N_GND_M1020_b N_VDD_M1003_b NWDIODE A=19.8481 P=23.39
pX33_noxref noxref_24 RN RN PROBETYPE=1
pX34_noxref noxref_25 D D PROBETYPE=1
pX35_noxref noxref_26 CK CK PROBETYPE=1
pX36_noxref noxref_27 QN QN PROBETYPE=1
pX37_noxref noxref_28 Q Q PROBETYPE=1
c_1783 A_926_521# 0 1.57671e-19 $X=4.63 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffr_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffr_l.spice
* Created: Mon Nov 16 20:39:15 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffr_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffr_l  GND VDD RN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* RN	RN
* VDD	VDD
* GND	GND
MM1022 N_A_110_115#_M1022_d N_RN_M1022_g N_GND_M1022_s N_GND_M1022_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1018 N_A_217_605#_M1018_d N_A_110_115#_M1018_g N_GND_M1018_s N_GND_M1022_b
+ NLOWVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_GND_M1007_d N_A_342_442#_M1007_g N_A_217_605#_M1018_d N_GND_M1022_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_576_115# N_D_M1008_g N_GND_M1008_s N_GND_M1022_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1031 N_A_342_442#_M1031_d N_A_618_89#_M1031_g A_576_115# N_GND_M1022_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1026 A_768_115# N_CK_M1026_g N_A_342_442#_M1031_d N_GND_M1022_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1029 N_GND_M1029_d N_A_217_605#_M1029_g A_768_115# N_GND_M1022_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1025 A_926_115# N_A_217_605#_M1025_g N_GND_M1029_d N_GND_M1022_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1019 N_A_998_115#_M1019_d N_CK_M1019_g A_926_115# N_GND_M1022_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1020 A_1118_115# N_A_618_89#_M1020_g N_A_998_115#_M1019_d N_GND_M1022_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1023 N_GND_M1023_d N_A_1160_89#_M1023_g A_1118_115# N_GND_M1022_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_A_618_89#_M1011_d N_CK_M1011_g N_GND_M1023_d N_GND_M1022_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1013 N_A_1160_89#_M1013_d N_A_998_115#_M1013_g N_GND_M1013_s N_GND_M1022_b
+ NLOWVT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_GND_M1015_d N_A_110_115#_M1015_g N_A_1160_89#_M1013_d N_GND_M1022_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_GND_M1017_d N_A_1160_89#_M1017_g N_QN_M1017_s N_GND_M1022_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_Q_M1009_d N_QN_M1009_g N_GND_M1017_d N_GND_M1022_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_110_115#_M1004_d N_RN_M1004_g N_VDD_M1004_s N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1014 A_300_605# N_A_110_115#_M1014_g N_A_217_605#_M1014_s N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_VDD_M1002_d N_A_342_442#_M1002_g A_300_605# N_VDD_M1004_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1027 A_576_521# N_D_M1027_g N_VDD_M1027_s N_VDD_M1004_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1024 N_A_342_442#_M1024_d N_CK_M1024_g A_576_521# N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1016 A_768_521# N_A_618_89#_M1016_g N_A_342_442#_M1024_d N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1021 N_VDD_M1021_d N_A_217_605#_M1021_g A_768_521# N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1012 A_926_521# N_A_217_605#_M1012_g N_VDD_M1021_d N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_998_115#_M1003_d N_A_618_89#_M1003_g A_926_521# N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 A_1118_521# N_CK_M1000_g N_A_998_115#_M1003_d N_VDD_M1004_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_1160_89#_M1006_g A_1118_521# N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1028 N_A_618_89#_M1028_d N_CK_M1028_g N_VDD_M1006_d N_VDD_M1004_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 A_1466_605# N_A_998_115#_M1005_g N_A_1160_89#_M1005_s N_VDD_M1004_b
+ PSHORT L=0.15 W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_VDD_M1030_d N_A_110_115#_M1030_g A_1466_605# N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VDD_M1010_d N_A_1160_89#_M1010_g N_QN_M1010_s N_VDD_M1004_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_Q_M1001_d N_QN_M1001_g N_VDD_M1010_d N_VDD_M1004_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX32_noxref N_GND_M1022_b N_VDD_M1004_b NWDIODE A=19.8481 P=23.39
pX33_noxref noxref_24 RN RN PROBETYPE=1
pX34_noxref noxref_25 D D PROBETYPE=1
pX35_noxref noxref_26 CK CK PROBETYPE=1
pX36_noxref noxref_27 QN QN PROBETYPE=1
pX37_noxref noxref_28 Q Q PROBETYPE=1
c_1778 A_926_521# 0 1.57671e-19 $X=4.63 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffr_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffs_1.spice
* Created: Mon Nov 16 20:39:21 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffs_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffs_1  GND VDD SN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* VDD	VDD
* GND	GND
MM1015 A_110_115# N_SN_M1015_g N_A_27_115#_M1015_s N_GND_M1015_b NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_GND_M1004_d N_A_152_89#_M1004_g A_110_115# N_GND_M1015_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_386_115# N_D_M1005_g N_GND_M1005_s N_GND_M1015_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1025 N_A_152_89#_M1025_d N_A_428_89#_M1025_g A_386_115# N_GND_M1015_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1019 A_578_115# N_CK_M1019_g N_A_152_89#_M1025_d N_GND_M1015_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1023 N_GND_M1023_d N_A_27_115#_M1023_g A_578_115# N_GND_M1015_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1016 A_736_115# N_A_27_115#_M1016_g N_GND_M1023_d N_GND_M1015_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1013 N_A_808_115#_M1013_d N_CK_M1013_g A_736_115# N_GND_M1015_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1006 A_928_115# N_A_428_89#_M1006_g N_A_808_115#_M1013_d N_GND_M1015_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1009 N_GND_M1009_d N_A_970_89#_M1009_g A_928_115# N_GND_M1015_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_A_428_89#_M1007_d N_CK_M1007_g N_GND_M1009_d N_GND_M1015_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1008 A_1276_115# N_A_808_115#_M1008_g N_A_970_89#_M1008_s N_GND_M1015_b NLOWVT
+ L=0.15 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_GND_M1029_d N_SN_M1029_g A_1276_115# N_GND_M1015_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_GND_M1011_d N_A_970_89#_M1011_g N_QN_M1011_s N_GND_M1015_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1000 N_Q_M1000_d N_QN_M1000_g N_GND_M1011_d N_GND_M1015_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1012 N_A_27_115#_M1012_d N_SN_M1012_g N_VDD_M1012_s N_VDD_M1012_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_VDD_M1027_d N_A_152_89#_M1027_g N_A_27_115#_M1012_d N_VDD_M1012_b
+ PSHORT L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 A_386_521# N_D_M1020_g N_VDD_M1020_s N_VDD_M1012_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1017 N_A_152_89#_M1017_d N_CK_M1017_g A_386_521# N_VDD_M1012_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1010 A_578_521# N_A_428_89#_M1010_g N_A_152_89#_M1017_d N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1014 N_VDD_M1014_d N_A_27_115#_M1014_g A_578_521# N_VDD_M1012_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 A_736_521# N_A_27_115#_M1002_g N_VDD_M1014_d N_VDD_M1012_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1028 N_A_808_115#_M1028_d N_A_428_89#_M1028_g A_736_521# N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1021 A_928_521# N_CK_M1021_g N_A_808_115#_M1028_d N_VDD_M1012_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1024 N_VDD_M1024_d N_A_970_89#_M1024_g A_928_521# N_VDD_M1012_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_428_89#_M1022_d N_CK_M1022_g N_VDD_M1024_d N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_970_89#_M1001_d N_A_808_115#_M1001_g N_VDD_M1001_s N_VDD_M1012_b
+ PSHORT L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_VDD_M1003_d N_SN_M1003_g N_A_970_89#_M1001_d N_VDD_M1012_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_VDD_M1026_d N_A_970_89#_M1026_g N_QN_M1026_s N_VDD_M1012_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_Q_M1018_d N_QN_M1018_g N_VDD_M1026_d N_VDD_M1012_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX30_noxref N_GND_M1015_b N_VDD_M1012_b NWDIODE A=18.0409 P=21.64
pX31_noxref noxref_23 SN SN PROBETYPE=1
pX32_noxref noxref_24 D D PROBETYPE=1
pX33_noxref noxref_25 CK CK PROBETYPE=1
pX34_noxref noxref_26 QN QN PROBETYPE=1
pX35_noxref noxref_27 Q Q PROBETYPE=1
c_1608 A_736_521# 0 1.57671e-19 $X=3.68 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffs_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffs_l.spice
* Created: Mon Nov 16 20:39:27 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffs_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffs_l  GND VDD SN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* VDD	VDD
* GND	GND
MM1016 A_110_115# N_SN_M1016_g N_A_27_115#_M1016_s N_GND_M1016_b NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_GND_M1004_d N_A_152_89#_M1004_g A_110_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_386_115# N_D_M1005_g N_GND_M1005_s N_GND_M1016_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1026 N_A_152_89#_M1026_d N_A_428_89#_M1026_g A_386_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1019 A_578_115# N_CK_M1019_g N_A_152_89#_M1026_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1023 N_GND_M1023_d N_A_27_115#_M1023_g A_578_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1017 A_736_115# N_A_27_115#_M1017_g N_GND_M1023_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1014 N_A_808_115#_M1014_d N_CK_M1014_g A_736_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1007 A_928_115# N_A_428_89#_M1007_g N_A_808_115#_M1014_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1
+ R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1010 N_GND_M1010_d N_A_970_89#_M1010_g A_928_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1008 N_A_428_89#_M1008_d N_CK_M1008_g N_GND_M1010_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1009 A_1276_115# N_A_808_115#_M1009_g N_A_970_89#_M1009_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_GND_M1029_d N_SN_M1029_g A_1276_115# N_GND_M1016_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_GND_M1012_d N_A_970_89#_M1012_g N_QN_M1012_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_Q_M1000_d N_QN_M1000_g N_GND_M1012_d N_GND_M1016_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_27_115#_M1013_d N_SN_M1013_g N_VDD_M1013_s N_VDD_M1013_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_VDD_M1027_d N_A_152_89#_M1027_g N_A_27_115#_M1013_d N_VDD_M1013_b
+ PSHORT L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1020 A_386_521# N_D_M1020_g N_VDD_M1020_s N_VDD_M1013_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1018 N_A_152_89#_M1018_d N_CK_M1018_g A_386_521# N_VDD_M1013_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1011 A_578_521# N_A_428_89#_M1011_g N_A_152_89#_M1018_d N_VDD_M1013_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1015 N_VDD_M1015_d N_A_27_115#_M1015_g A_578_521# N_VDD_M1013_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 A_736_521# N_A_27_115#_M1002_g N_VDD_M1015_d N_VDD_M1013_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1028 N_A_808_115#_M1028_d N_A_428_89#_M1028_g A_736_521# N_VDD_M1013_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1021 A_928_521# N_CK_M1021_g N_A_808_115#_M1028_d N_VDD_M1013_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1025 N_VDD_M1025_d N_A_970_89#_M1025_g A_928_521# N_VDD_M1013_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_428_89#_M1022_d N_CK_M1022_g N_VDD_M1025_d N_VDD_M1013_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_970_89#_M1001_d N_A_808_115#_M1001_g N_VDD_M1001_s N_VDD_M1013_b
+ PSHORT L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_VDD_M1003_d N_SN_M1003_g N_A_970_89#_M1001_d N_VDD_M1013_b PSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VDD_M1006_d N_A_970_89#_M1006_g N_QN_M1006_s N_VDD_M1013_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1024 N_Q_M1024_d N_QN_M1024_g N_VDD_M1006_d N_VDD_M1013_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX30_noxref N_GND_M1016_b N_VDD_M1013_b NWDIODE A=18.0409 P=21.64
pX31_noxref noxref_23 SN SN PROBETYPE=1
pX32_noxref noxref_24 D D PROBETYPE=1
pX33_noxref noxref_25 CK CK PROBETYPE=1
pX34_noxref noxref_26 QN QN PROBETYPE=1
pX35_noxref noxref_27 Q Q PROBETYPE=1
c_1617 A_736_521# 0 1.57671e-19 $X=3.68 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffs_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffsr_1.spice
* Created: Mon Nov 16 20:39:32 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffsr_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffsr_1  GND VDD RN SN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* RN	RN
* VDD	VDD
* GND	GND
MM1016 N_A_110_115#_M1016_d N_RN_M1016_g N_GND_M1016_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1034 N_A_217_521#_M1034_d N_A_110_115#_M1034_g N_GND_M1034_s N_GND_M1016_b
+ NLOWVT L=0.15 W=0.42 AD=0.0767474 AS=0.1113 PD=0.770722 PS=1.37 NRD=17.136
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1015 A_400_115# N_SN_M1015_g N_A_217_521#_M1034_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.100503 PD=0.76 PS=1.00928 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1003 N_GND_M1003_d N_A_432_424#_M1003_g A_400_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.9 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1005 A_662_115# N_D_M1005_g N_GND_M1005_s N_GND_M1016_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1035 N_A_432_424#_M1035_d N_A_704_89#_M1035_g A_662_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1026 A_854_115# N_CK_M1026_g N_A_432_424#_M1035_d N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1020 N_GND_M1020_d N_A_217_521#_M1020_g A_854_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1023 A_1012_115# N_A_217_521#_M1023_g N_GND_M1020_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1021 N_A_1084_115#_M1021_d N_CK_M1021_g A_1012_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1017 A_1204_115# N_A_704_89#_M1017_g N_A_1084_115#_M1021_d N_GND_M1016_b
+ NLOWVT L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54
+ M=1 R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1006 N_GND_M1006_d N_A_1246_89#_M1006_g A_1204_115# N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_A_704_89#_M1011_d N_CK_M1011_g N_GND_M1006_d N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1013 A_1552_115# N_A_1084_115#_M1013_g N_GND_M1013_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1004 N_A_1246_89#_M1004_d N_SN_M1004_g A_1552_115# N_GND_M1016_b NLOWVT L=0.15
+ W=0.55 AD=0.100503 AS=0.05775 PD=1.00928 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1022 N_GND_M1022_d N_A_110_115#_M1022_g N_A_1246_89#_M1004_d N_GND_M1016_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0767474 PD=1.37 PS=0.770722 NRD=0
+ NRS=17.136 M=1 R=2.8 SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_GND_M1007_d N_A_1246_89#_M1007_g N_QN_M1007_s N_GND_M1016_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_GND_M1007_d N_GND_M1016_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1001 N_A_110_115#_M1001_d N_RN_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_300_521#_M1000_d N_A_110_115#_M1000_g N_A_217_521#_M1000_s
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0
+ NRS=0 M=1 R=8.4 SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1024 N_VDD_M1024_d N_SN_M1024_g N_A_300_521#_M1000_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_300_521#_M1027_d N_A_432_424#_M1027_g N_VDD_M1024_d N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1028 A_662_521# N_D_M1028_g N_VDD_M1028_s N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1018 N_A_432_424#_M1018_d N_CK_M1018_g A_662_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1014 A_854_521# N_A_704_89#_M1014_g N_A_432_424#_M1018_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1009 N_VDD_M1009_d N_A_217_521#_M1009_g A_854_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1012 A_1012_521# N_A_217_521#_M1012_g N_VDD_M1009_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1010 N_A_1084_115#_M1010_d N_A_704_89#_M1010_g A_1012_521# N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778
+ NRS=7.8012 M=1 R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 A_1204_521# N_CK_M1002_g N_A_1084_115#_M1010_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1029 N_VDD_M1029_d N_A_1246_89#_M1029_g A_1204_521# N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1031 N_A_704_89#_M1031_d N_CK_M1031_g N_VDD_M1029_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1033 N_VDD_M1033_d N_A_1084_115#_M1033_g N_A_1469_521#_M1033_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_A_1469_521#_M1019_d N_SN_M1019_g N_VDD_M1033_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_A_1246_89#_M1025_d N_A_110_115#_M1025_g N_A_1469_521#_M1019_d
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0
+ NRS=0 M=1 R=8.4 SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1030 N_VDD_M1030_d N_A_1246_89#_M1030_g N_QN_M1030_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_Q_M1032_d N_QN_M1032_g N_VDD_M1030_d N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref N_GND_M1016_b N_VDD_M1001_b NWDIODE A=21.63 P=25.12
pX37_noxref noxref_27 RN RN PROBETYPE=1
pX38_noxref noxref_28 D D PROBETYPE=1
pX39_noxref noxref_29 CK CK PROBETYPE=1
pX40_noxref noxref_30 SN SN PROBETYPE=1
pX41_noxref noxref_31 QN QN PROBETYPE=1
pX42_noxref noxref_32 Q Q PROBETYPE=1
c_2169 A_1012_521# 0 1.57671e-19 $X=5.06 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffsr_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dffsr_l.spice
* Created: Mon Nov 16 20:39:38 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__dffsr_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dffsr_l  GND VDD RN SN D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* SN	SN
* RN	RN
* VDD	VDD
* GND	GND
MM1018 N_A_110_115#_M1018_d N_RN_M1018_g N_GND_M1018_s N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1034 N_A_217_521#_M1034_d N_A_110_115#_M1034_g N_GND_M1034_s N_GND_M1018_b
+ NLOWVT L=0.15 W=0.42 AD=0.0767474 AS=0.1113 PD=0.770722 PS=1.37 NRD=17.136
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1017 A_400_115# N_SN_M1017_g N_A_217_521#_M1034_d N_GND_M1018_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.100503 PD=0.76 PS=1.00928 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1005 N_GND_M1005_d N_A_432_424#_M1005_g A_400_115# N_GND_M1018_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.9 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1007 A_662_115# N_D_M1007_g N_GND_M1007_s N_GND_M1018_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.7 A=0.0825 P=1.4 MULT=1
MM1035 N_A_432_424#_M1035_d N_A_704_89#_M1035_g A_662_115# N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1028 A_854_115# N_CK_M1028_g N_A_432_424#_M1035_d N_GND_M1018_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.1 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1022 N_GND_M1022_d N_A_217_521#_M1022_g A_854_115# N_GND_M1018_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75001.5 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1025 A_1012_115# N_A_217_521#_M1025_g N_GND_M1022_d N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1023 N_A_1084_115#_M1023_d N_CK_M1023_g A_1012_115# N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1
+ R=3.66667 SA=75002.3 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1019 A_1204_115# N_A_704_89#_M1019_g N_A_1084_115#_M1023_d N_GND_M1018_b
+ NLOWVT L=0.15 W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54
+ M=1 R=3.66667 SA=75002.9 SB=75001 A=0.0825 P=1.4 MULT=1
MM1008 N_GND_M1008_d N_A_1246_89#_M1008_g A_1204_115# N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75003.3 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1013 N_A_704_89#_M1013_d N_CK_M1013_g N_GND_M1008_d N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1015 A_1552_115# N_A_1084_115#_M1015_g N_GND_M1015_s N_GND_M1018_b NLOWVT
+ L=0.15 W=0.55 AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1006 N_A_1246_89#_M1006_d N_SN_M1006_g A_1552_115# N_GND_M1018_b NLOWVT L=0.15
+ W=0.55 AD=0.100503 AS=0.05775 PD=1.00928 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.5 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1024 N_GND_M1024_d N_A_110_115#_M1024_g N_A_1246_89#_M1006_d N_GND_M1018_b
+ NLOWVT L=0.15 W=0.42 AD=0.1113 AS=0.0767474 PD=1.37 PS=0.770722 NRD=0
+ NRS=17.136 M=1 R=2.8 SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_GND_M1009_d N_A_1246_89#_M1009_g N_QN_M1009_s N_GND_M1018_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_Q_M1010_d N_QN_M1010_g N_GND_M1009_d N_GND_M1018_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_110_115#_M1001_d N_RN_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_300_521#_M1000_d N_A_110_115#_M1000_g N_A_217_521#_M1000_s
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0
+ NRS=0 M=1 R=8.4 SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1026 N_VDD_M1026_d N_SN_M1026_g N_A_300_521#_M1000_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_A_300_521#_M1029_d N_A_432_424#_M1029_g N_VDD_M1026_d N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1030 A_662_521# N_D_M1030_g N_VDD_M1030_s N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1020 N_A_432_424#_M1020_d N_CK_M1020_g A_662_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1016 A_854_521# N_A_704_89#_M1016_g N_A_432_424#_M1020_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.1 SB=75002.7 A=0.189 P=2.82 MULT=1
MM1011 N_VDD_M1011_d N_A_217_521#_M1011_g A_854_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1014 A_1012_521# N_A_217_521#_M1014_g N_VDD_M1011_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1012 N_A_1084_115#_M1012_d N_A_704_89#_M1012_g A_1012_521# N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778
+ NRS=7.8012 M=1 R=8.4 SA=75002.3 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 A_1204_521# N_CK_M1002_g N_A_1084_115#_M1012_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75002.9 SB=75001 A=0.189 P=2.82 MULT=1
MM1031 N_VDD_M1031_d N_A_1246_89#_M1031_g A_1204_521# N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75003.3 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_A_704_89#_M1032_d N_CK_M1032_g N_VDD_M1031_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1033 N_VDD_M1033_d N_A_1084_115#_M1033_g N_A_1469_521#_M1033_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_A_1469_521#_M1021_d N_SN_M1021_g N_VDD_M1033_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_1246_89#_M1027_d N_A_110_115#_M1027_g N_A_1469_521#_M1021_d
+ N_VDD_M1001_b PSHORT L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0
+ NRS=0 M=1 R=8.4 SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_1246_89#_M1003_g N_QN_M1003_s N_VDD_M1001_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1004 N_Q_M1004_d N_QN_M1004_g N_VDD_M1003_d N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX36_noxref N_GND_M1018_b N_VDD_M1001_b NWDIODE A=21.63 P=25.12
pX37_noxref noxref_27 RN RN PROBETYPE=1
pX38_noxref noxref_28 D D PROBETYPE=1
pX39_noxref noxref_29 CK CK PROBETYPE=1
pX40_noxref noxref_30 SN SN PROBETYPE=1
pX41_noxref noxref_31 QN QN PROBETYPE=1
pX42_noxref noxref_32 Q Q PROBETYPE=1
c_2177 A_1012_521# 0 1.57671e-19 $X=5.06 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dffsr_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dlat_1.spice
* Created: Fri Nov 12 15:10:04 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__dlat_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__dlat_1  GND VDD D CK ON Q
*
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1004 A_115_115# N_D_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1015 N_D_M1015_d N_CK_M1015_g A_115_115# N_GND_M1004_b NLOWVT L=0.15 W=0.52
+ AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1013 A_307_115# N_A_157_349#_M1013_g N_D_M1015_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.1 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_349_89#_M1007_g A_307_115# N_GND_M1004_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.5 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_A_157_349#_M1008_d N_CK_M1008_g N_GND_M1007_d N_GND_M1004_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.9 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_A_349_89#_M1010_d N_D_M1010_g N_GND_M1010_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1011 N_GND_M1011_d N_A_349_89#_M1011_g N_ON_M1011_s N_GND_M1004_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1012 N_Q_M1012_d N_ON_M1012_g N_GND_M1011_d N_GND_M1004_b NLOWVT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1014 A_115_521# N_D_M1014_g N_VDD_M1014_s N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_D_M1009_d N_A_157_349#_M1009_g A_115_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1006 A_307_521# N_CK_M1006_g N_D_M1009_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.1 SB=75001 A=0.189 P=2.82 MULT=1
MM1000 N_VDD_M1000_d N_A_349_89#_M1000_g A_307_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_157_349#_M1001_d N_CK_M1001_g N_VDD_M1000_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_349_89#_M1002_d N_D_M1002_g N_VDD_M1002_s N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_349_89#_M1003_g N_ON_M1003_s N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Q_M1005_d N_ON_M1005_g N_VDD_M1003_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref N_GND_M1004_b N_VDD_M1014_b NWDIODE A=10.5987 P=14.41
pX17_noxref noxref_13 D D PROBETYPE=1
pX18_noxref noxref_14 CK CK PROBETYPE=1
pX19_noxref noxref_15 ON ON PROBETYPE=1
pX20_noxref noxref_16 Q Q PROBETYPE=1
c_836 A_115_521# 0 1.57671e-19 $X=0.575 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dlat_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__dlat_l.spice
* Created: Fri Nov 12 15:10:12 2021
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__dlat_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__dlat_l  GND VDD D CK ON Q
*
* Q	Q
* ON	ON
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1003 A_115_115# N_D_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15 W=0.52
+ AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1015 N_D_M1015_d N_CK_M1015_g A_115_115# N_GND_M1003_b NLOWVT L=0.15 W=0.52
+ AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1013 A_307_115# N_A_157_349#_M1013_g N_D_M1015_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.1 SB=75001 A=0.078 P=1.34 MULT=1
MM1006 N_GND_M1006_d N_A_349_89#_M1006_g A_307_115# N_GND_M1003_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.5 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_A_157_349#_M1008_d N_CK_M1008_g N_GND_M1006_d N_GND_M1003_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.9 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_A_349_89#_M1010_d N_D_M1010_g N_GND_M1010_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.52 AD=0.1378 AS=0.1378 PD=1.57 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1011 N_GND_M1011_d N_A_349_89#_M1011_g N_ON_M1011_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.36 AD=0.0504 AS=0.0954 PD=0.64 PS=1.25 NRD=0 NRS=0 M=1 R=2.4
+ SA=75000.2 SB=75000.6 A=0.054 P=1.02 MULT=1
MM1012 N_Q_M1012_d N_ON_M1012_g N_GND_M1011_d N_GND_M1003_b NLOWVT L=0.15 W=0.36
+ AD=0.0954 AS=0.0504 PD=1.25 PS=0.64 NRD=0 NRS=0 M=1 R=2.4 SA=75000.6
+ SB=75000.2 A=0.054 P=1.02 MULT=1
MM1014 A_115_521# N_D_M1014_g N_VDD_M1014_s N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_D_M1009_d N_A_157_349#_M1009_g A_115_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1004 A_307_521# N_CK_M1004_g N_D_M1009_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.1 SB=75001 A=0.189 P=2.82 MULT=1
MM1000 N_VDD_M1000_d N_A_349_89#_M1000_g A_307_521# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_157_349#_M1001_d N_CK_M1001_g N_VDD_M1000_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_A_349_89#_M1002_d N_D_M1002_g N_VDD_M1002_s N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_349_89#_M1005_g N_ON_M1005_s N_VDD_M1014_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_Q_M1007_d N_ON_M1007_g N_VDD_M1005_d N_VDD_M1014_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX16_noxref N_GND_M1003_b N_VDD_M1014_b NWDIODE A=10.5987 P=14.41
pX17_noxref noxref_13 D D PROBETYPE=1
pX18_noxref noxref_14 CK CK PROBETYPE=1
pX19_noxref noxref_15 ON ON PROBETYPE=1
pX20_noxref noxref_16 Q Q PROBETYPE=1
c_838 A_115_521# 0 1.57671e-19 $X=0.575 $Y=2.605
*
.include "sky130_osu_sc_12T_hs__dlat_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_1.spice
* Created: Mon Nov 16 20:39:56 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_1  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_Y_M1001_d N_A_M1001_g N_GND_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.1424 P=6.2
pX3_noxref noxref_5 A A PROBETYPE=1
pX4_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_2.spice
* Created: Mon Nov 16 20:40:01 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_2.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_2  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=3.0488 P=7.08
pX5_noxref noxref_5 A A PROBETYPE=1
pX6_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_2.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_3.spice
* Created: Mon Nov 16 20:40:07 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_3.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_3  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1003 N_GND_M1002_d N_A_M1003_g N_Y_M1003_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1000_d N_A_M1004_g N_VDD_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VDD_M1004_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=3.9552 P=7.96
pX7_noxref noxref_5 A A PROBETYPE=1
pX8_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_3.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_4.spice
* Created: Mon Nov 16 20:40:13 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_4.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_4  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1002_d N_A_M1004_g N_Y_M1004_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_GND_M1007_d N_A_M1007_g N_Y_M1004_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=4.8616 P=8.84
pX9_noxref noxref_5 A A PROBETYPE=1
pX10_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_4.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_6.spice
* Created: Mon Nov 16 20:40:18 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_6.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_6  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1002_d N_A_M1004_g N_Y_M1004_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1009 N_GND_M1009_d N_A_M1009_g N_Y_M1004_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1010 N_GND_M1009_d N_A_M1010_g N_Y_M1010_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_GND_M1011_d N_A_M1011_g N_Y_M1010_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VDD_M1008_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=6.6744 P=10.6
pX13_noxref noxref_5 A A PROBETYPE=1
pX14_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_6.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_8.spice
* Created: Mon Nov 16 20:40:24 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_8  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1006 N_GND_M1002_d N_A_M1006_g N_Y_M1006_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1011 N_GND_M1011_d N_A_M1011_g N_Y_M1006_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1012 N_GND_M1011_d N_A_M1012_g N_Y_M1012_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1013 N_GND_M1013_d N_A_M1013_g N_Y_M1012_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1014 N_GND_M1013_d N_A_M1014_g N_Y_M1014_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1015 N_GND_M1015_d N_A_M1015_g N_Y_M1014_s N_GND_M1001_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1000_d N_A_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1004_d N_A_M1005_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1007_d N_A_M1008_g N_VDD_M1008_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VDD_M1008_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1009_d N_A_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=8.4769 P=12.35
pX17_noxref noxref_5 A A PROBETYPE=1
pX18_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_8.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_10.spice
* Created: Mon Nov 16 20:39:50 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_10.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_10  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_M1002_g N_Y_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1004 N_GND_M1004_d N_A_M1004_g N_Y_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.6 A=0.0825 P=1.4 MULT=1
MM1008 N_GND_M1004_d N_A_M1008_g N_Y_M1008_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1009 N_GND_M1009_d N_A_M1009_g N_Y_M1008_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1012 N_GND_M1009_d N_A_M1012_g N_Y_M1012_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1015 N_GND_M1015_d N_A_M1015_g N_Y_M1012_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1016 N_GND_M1015_d N_A_M1016_g N_Y_M1016_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1017 N_GND_M1017_d N_A_M1017_g N_Y_M1016_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1018 N_GND_M1017_d N_A_M1018_g N_Y_M1018_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1019 N_GND_M1019_d N_A_M1019_g N_Y_M1018_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75004.1
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VDD_M1001_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VDD_M1001_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1003_d N_A_M1005_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VDD_M1005_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VDD_M1007_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1010_d N_A_M1010_g N_VDD_M1007_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1010_d N_A_M1011_g N_VDD_M1011_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VDD_M1011_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1013_d N_A_M1014_g N_VDD_M1014_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=10.2897 P=14.11
pX21_noxref noxref_5 A A PROBETYPE=1
pX22_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_10.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__inv_l.spice
* Created: Mon Nov 16 20:40:30 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__inv_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__inv_l  GND VDD A Y
*
* Y	Y
* A	A
* VDD	VDD
* GND	GND
MM1001 N_Y_M1001_d N_A_M1001_g N_GND_M1001_s N_GND_M1001_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.132 P=6.18
pX3_noxref noxref_5 A A PROBETYPE=1
pX4_noxref noxref_6 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__inv_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__mux2_1.spice
* Created: Mon Nov 16 20:40:35 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__mux2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__mux2_1  GND VDD S0 A0 Y A1
*
* A1	A1
* Y	Y
* A0	A0
* S0	S0
* VDD	VDD
* GND	GND
MM1004 N_A_110_115#_M1004_d N_S0_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_Y_M1003_d N_A_110_115#_M1003_g N_A0_M1003_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_A1_M1002_d N_S0_M1002_g N_Y_M1003_d N_GND_M1004_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1001 N_A_110_115#_M1001_d N_S0_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_S0_M1000_g N_A0_M1000_s N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_A1_M1005_d N_A_110_115#_M1005_g N_Y_M1000_d N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1001_b NWDIODE A=5.7886 P=9.74
pX7_noxref noxref_8 S0 S0 PROBETYPE=1
pX8_noxref noxref_9 A0 A0 PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
pX10_noxref noxref_11 A1 A1 PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__mux2_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__nand2_1.spice
* Created: Mon Nov 16 20:40:41 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__nand2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__nand2_1  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1002 A_110_115# N_A_M1002_g N_Y_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.14575 PD=0.76 PS=1.63 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_B_M1001_g A_110_115# N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667
+ SA=75000.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_B_M1003_g N_Y_M1000_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=3.0385 P=7.07
pX5_noxref noxref_7 A A PROBETYPE=1
pX6_noxref noxref_8 Y Y PROBETYPE=1
pX7_noxref noxref_9 B B PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__nand2_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__nand2_l.spice
* Created: Mon Nov 16 20:40:47 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__nand2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__nand2_l  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1002 A_110_115# N_A_M1002_g N_Y_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_GND_M1000_d N_B_M1000_g A_110_115# N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g N_VDD_M1001_s N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_VDD_M1003_d N_B_M1003_g N_Y_M1001_d N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=2.49275 P=6.33
pX5_noxref noxref_7 A A PROBETYPE=1
pX6_noxref noxref_8 Y Y PROBETYPE=1
pX7_noxref noxref_9 B B PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__nand2_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__ncgate_1.spice
* Created: Tue Apr 26 09:48:41 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__ncgate_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__ncgate_1  GND Q SE E CK ECK
*
* ECK	ECK
* CK	CK
* E	E
* SE	SE
* Q	VDD
* GND	GND
MM1011 N_A_N233_516#_M1011_d N_SE_M1011_g N_GND_M1011_s N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1021 N_GND_M1021_d N_E_M1021_g N_A_N233_516#_M1011_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_A_86_236#_M1001_g N_A_43_110#_M1001_s N_GND_M1011_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1000 A_212_110# N_A_N233_516#_M1000_g N_GND_M1001_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1023 N_A_86_236#_M1023_d N_CK_M1023_g A_212_110# N_GND_M1011_b NLOWVT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1012 A_404_110# N_A_254_419#_M1012_g N_A_86_236#_M1023_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1
+ R=3.46667 SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1004 N_GND_M1004_d N_A_43_110#_M1004_g A_404_110# N_GND_M1011_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1005 N_A_254_419#_M1005_d N_CK_M1005_g N_GND_M1004_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1018 N_GND_M1018_d N_A_43_110#_M1018_g N_A_687_110#_M1018_s N_GND_M1011_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1007 N_A_856_110#_M1007_d N_A_687_110#_M1007_g N_GND_M1018_d N_GND_M1011_b
+ NLOWVT L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1016 N_A_963_516#_M1016_d N_A_687_110#_M1016_g N_GND_M1016_s N_GND_M1011_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1017 N_GND_M1017_d N_CK_M1017_g N_A_963_516#_M1016_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1010 N_ECK_M1010_d N_A_963_516#_M1010_g N_GND_M1017_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1014 A_N150_516# N_SE_M1014_g N_A_N233_516#_M1014_s N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_Q_M1019_d N_E_M1019_g A_N150_516# N_Q_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_Q_M1003_d N_A_86_236#_M1003_g N_A_43_110#_M1003_s N_Q_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 A_212_516# N_A_N233_516#_M1002_g N_Q_M1003_d N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1025 N_A_86_236#_M1025_d N_A_254_419#_M1025_g A_212_516# N_Q_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1015 A_404_516# N_CK_M1015_g N_A_86_236#_M1025_d N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1006 N_Q_M1006_d N_A_43_110#_M1006_g A_404_516# N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_254_419#_M1008_d N_CK_M1008_g N_Q_M1006_d N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_Q_M1024_d N_A_43_110#_M1024_g N_A_687_110#_M1024_s N_Q_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_A_856_110#_M1009_d N_A_687_110#_M1009_g N_Q_M1024_d N_Q_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1020 A_1046_516# N_A_687_110#_M1020_g N_A_963_516#_M1020_s N_Q_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_Q_M1022_d N_CK_M1022_g A_1046_516# N_Q_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_ECK_M1013_d N_A_963_516#_M1013_g N_Q_M1022_d N_Q_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1011_b N_Q_M1014_b NWDIODE A=16.3094 P=19.99
pX27_noxref noxref_20 N_SE_X27_noxref_CONDUCTOR SE PROBETYPE=1
pX28_noxref noxref_21 N_E_X28_noxref_CONDUCTOR E PROBETYPE=1
pX29_noxref noxref_22 CK CK PROBETYPE=1
pX30_noxref noxref_23 ECK ECK PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__ncgate_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__ncgateCKa_new.spice
* Created: Tue Apr 26 09:48:49 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__ncgateCKa_new.pex.spice"
.subckt sky130_osu_sc_12T_hs__ncgateCKa_new  GND VDD SE E CK Q CKA ECK
*
* ECK	ECK
* CKA	CKA
* Q	Q
* CK	CK
* E	E
* SE	SE
* VDD	VDD
* GND	GND
MM1011 N_A_N233_516#_M1011_d N_SE_M1011_g N_GND_M1011_s N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1021 N_GND_M1021_d N_E_M1021_g N_A_N233_516#_M1011_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 N_GND_M1001_d N_A_86_236#_M1001_g N_A_43_110#_M1001_s N_GND_M1011_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1000 A_212_110# N_A_N233_516#_M1000_g N_GND_M1001_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1023 N_A_86_236#_M1023_d N_CK_M1023_g A_212_110# N_GND_M1011_b NLOWVT L=0.15
+ W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1 R=3.46667
+ SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1012 A_404_110# N_A_254_419#_M1012_g N_A_86_236#_M1023_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1
+ R=3.46667 SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1004 N_GND_M1004_d N_A_43_110#_M1004_g A_404_110# N_GND_M1011_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1005 N_A_254_419#_M1005_d N_CK_M1005_g N_GND_M1004_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1018 N_GND_M1018_d N_A_43_110#_M1018_g N_Q_M1018_s N_GND_M1011_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1007 N_Q_M1007_d N_Q_M1007_g N_GND_M1018_d N_GND_M1011_b NLOWVT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1016 N_A_963_516#_M1016_d N_Q_M1016_g N_GND_M1016_s N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1017 N_GND_M1017_d N_CKA_M1017_g N_A_963_516#_M1016_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.0728 PD=0.8 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1010 N_ECK_M1010_d N_A_963_516#_M1010_g N_GND_M1017_d N_GND_M1011_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1014 A_N150_516# N_SE_M1014_g N_A_N233_516#_M1014_s N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_VDD_M1019_d N_E_M1019_g A_N150_516# N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_86_236#_M1003_g N_A_43_110#_M1003_s N_VDD_M1014_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1002 A_212_516# N_A_N233_516#_M1002_g N_VDD_M1003_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1025 N_A_86_236#_M1025_d N_A_254_419#_M1025_g A_212_516# N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1
+ R=8.4 SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1015 A_404_516# N_CK_M1015_g N_A_86_236#_M1025_d N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_43_110#_M1006_g A_404_516# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_254_419#_M1008_d N_CK_M1008_g N_VDD_M1006_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1024 N_VDD_M1024_d N_A_43_110#_M1024_g N_Q_M1024_s N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_Q_M1009_d N_Q_M1009_g N_VDD_M1024_d N_VDD_M1014_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1020 A_1046_516# N_Q_M1020_g N_A_963_516#_M1020_s N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_VDD_M1022_d N_CKA_M1022_g A_1046_516# N_VDD_M1014_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_ECK_M1013_d N_A_963_516#_M1013_g N_VDD_M1022_d N_VDD_M1014_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1011_b N_VDD_M1014_b NWDIODE A=16.3094 P=19.99
pX27_noxref noxref_20 N_SE_X27_noxref_CONDUCTOR SE PROBETYPE=1
pX28_noxref noxref_21 N_E_X28_noxref_CONDUCTOR E PROBETYPE=1
pX29_noxref noxref_22 CK CK PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
pX31_noxref noxref_24 Q Q PROBETYPE=1
pX32_noxref noxref_25 CKA CKA PROBETYPE=1
pX33_noxref noxref_26 ECK ECK PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__ncgateCKa_new.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__ndlat_1.spice
* Created: Tue Apr 26 09:48:58 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__ndlat_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__ndlat_1  GND VDD D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_161_241#_M1002_g N_A_118_115#_M1002_s N_GND_M1002_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1015 A_287_115# N_D_M1015_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15 W=0.52
+ AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1011 N_A_161_241#_M1011_d N_A_329_89#_M1011_g A_287_115# N_GND_M1002_b NLOWVT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1007 A_479_115# N_CK_M1007_g N_A_161_241#_M1011_d N_GND_M1002_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1009 N_GND_M1009_d N_A_118_115#_M1009_g A_479_115# N_GND_M1002_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1004 N_A_329_89#_M1004_d N_CK_M1004_g N_GND_M1009_d N_GND_M1002_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_GND_M1010_d N_A_118_115#_M1010_g N_QN_M1010_s N_GND_M1002_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1012 N_Q_M1012_d N_QN_M1012_g N_GND_M1010_d N_GND_M1002_b NLOWVT L=0.15 W=0.52
+ AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1013 N_VDD_M1013_d N_A_161_241#_M1013_g N_A_118_115#_M1013_s VDD PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1008 A_287_521# N_D_M1008_g N_VDD_M1013_d VDD PSHORT L=0.15 W=1.26 AD=0.1323
+ AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6 SB=75001.9
+ A=0.189 P=2.82 MULT=1
MM1005 N_A_161_241#_M1005_d N_CK_M1005_g A_287_521# VDD PSHORT L=0.15 W=1.26
+ AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 A_479_521# N_A_329_89#_M1000_g N_A_161_241#_M1005_d VDD PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1001 N_VDD_M1001_d N_A_118_115#_M1001_g A_479_521# VDD PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_329_89#_M1014_d N_CK_M1014_g N_VDD_M1001_d VDD PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_118_115#_M1003_g N_QN_M1003_s VDD PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_Q_M1006_d N_QN_M1006_g N_VDD_M1003_d VDD PSHORT L=0.15 W=1.26 AD=0.3339
+ AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75000.2 A=0.189
+ P=2.82 MULT=1
DX16_noxref N_GND_M1002_b VDD NWDIODE A=9.998 P=13.83
pX17_noxref noxref_14 D D PROBETYPE=1
pX18_noxref noxref_15 CK CK PROBETYPE=1
pX19_noxref noxref_16 QN QN PROBETYPE=1
pX20_noxref noxref_17 Q Q PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__ndlat_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__ndlat_l.spice
* Created: Tue Apr 26 09:49:06 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__ndlat_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__ndlat_l  GND VDD D CK QN Q
*
* Q	Q
* QN	QN
* CK	CK
* D	D
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_A_161_241#_M1002_g N_A_118_115#_M1002_s N_GND_M1002_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1015 A_287_115# N_D_M1015_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15 W=0.52
+ AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001.9 A=0.078 P=1.34 MULT=1
MM1011 N_A_161_241#_M1011_d N_A_329_89#_M1011_g A_287_115# N_GND_M1002_b NLOWVT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1005 A_479_115# N_CK_M1005_g N_A_161_241#_M1011_d N_GND_M1002_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1009 N_GND_M1009_d N_A_118_115#_M1009_g A_479_115# N_GND_M1002_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1003 N_A_329_89#_M1003_d N_CK_M1003_g N_GND_M1009_d N_GND_M1002_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_GND_M1010_d N_A_118_115#_M1010_g N_QN_M1010_s N_GND_M1002_b NLOWVT
+ L=0.15 W=0.37 AD=0.0518 AS=0.09805 PD=0.65 PS=1.27 NRD=0 NRS=0 M=1 R=2.46667
+ SA=75000.2 SB=75000.6 A=0.0555 P=1.04 MULT=1
MM1012 N_Q_M1012_d N_QN_M1012_g N_GND_M1010_d N_GND_M1002_b NLOWVT L=0.15 W=0.37
+ AD=0.09805 AS=0.0518 PD=1.27 PS=0.65 NRD=0 NRS=0 M=1 R=2.46667 SA=75000.6
+ SB=75000.2 A=0.0555 P=1.04 MULT=1
MM1013 N_VDD_M1013_d N_A_161_241#_M1013_g N_A_118_115#_M1013_s VDD PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1007 A_287_521# N_D_M1007_g N_VDD_M1013_d VDD PSHORT L=0.15 W=1.26 AD=0.1323
+ AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6 SB=75001.9
+ A=0.189 P=2.82 MULT=1
MM1004 N_A_161_241#_M1004_d N_CK_M1004_g A_287_521# VDD PSHORT L=0.15 W=1.26
+ AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 A_479_521# N_A_329_89#_M1000_g N_A_161_241#_M1004_d VDD PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1001 N_VDD_M1001_d N_A_118_115#_M1001_g A_479_521# VDD PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_A_329_89#_M1014_d N_CK_M1014_g N_VDD_M1001_d VDD PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_118_115#_M1006_g N_QN_M1006_s VDD PSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_Q_M1008_d N_QN_M1008_g N_VDD_M1006_d VDD PSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75000.2 A=0.126
+ P=1.98 MULT=1
DX16_noxref N_GND_M1002_b VDD NWDIODE A=9.9567 P=13.79
pX17_noxref noxref_14 D D PROBETYPE=1
pX18_noxref noxref_15 CK CK PROBETYPE=1
pX19_noxref noxref_16 QN QN PROBETYPE=1
pX20_noxref noxref_17 Q Q PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__ndlat_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__nor2_1.spice
* Created: Mon Nov 16 20:40:52 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__nor2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__nor2_1  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1002 N_Y_M1002_d N_B_M1002_g N_GND_M1002_s N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1002_d N_GND_M1002_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1003_d N_A_M1003_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX4_noxref N_GND_M1002_b N_VDD_M1000_b NWDIODE A=3.0385 P=7.07
pX5_noxref noxref_7 B B PROBETYPE=1
pX6_noxref noxref_8 Y Y PROBETYPE=1
pX7_noxref noxref_9 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__nor2_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__nor2_l.spice
* Created: Mon Nov 16 20:41:03 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__nor2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__nor2_l  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_Y_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_Y_M1003_d N_GND_M1003_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1002 A_110_605# N_B_M1002_g N_Y_M1002_s N_VDD_M1002_b PSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g A_110_605# N_VDD_M1002_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX4_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=2.49275 P=6.33
pX5_noxref noxref_7 Y Y PROBETYPE=1
pX6_noxref noxref_8 B B PROBETYPE=1
pX7_noxref noxref_9 A A PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__nor2_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__oai21_l.spice
* Created: Mon Nov 16 20:41:09 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__oai21_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__oai21_l  GND VDD A0 A1 B0 Y
*
* Y	Y
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1004 N_GND_M1004_d N_A0_M1004_g N_A_27_114#_M1004_s N_GND_M1004_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_114#_M1001_d N_A1_M1001_g N_GND_M1004_d N_GND_M1004_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_114#_M1001_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_A0_M1000_g N_Y_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A1_M1005_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.23814 AS=0.1323 PD=1.92 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1003_d N_B0_M1003_g N_VDD_M1005_d N_VDD_M1000_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.15876 PD=2.21 PS=1.28 NRD=0 NRS=14.0658 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_9 A0 A0 PROBETYPE=1
pX8_noxref noxref_10 A1 A1 PROBETYPE=1
pX9_noxref noxref_11 B0 B0 PROBETYPE=1
pX10_noxref noxref_12 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__oai21_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__oai22_l.spice
* Created: Mon Nov 16 20:41:14 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__oai22_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__oai22_l  GND VDD A0 A1 B0 B1 Y
*
* Y	Y
* B1	B1
* B0	B0
* A1	A1
* A0	A0
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_A0_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 N_A_27_115#_M1001_d N_A1_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_B0_M1002_g N_A_27_115#_M1001_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_A_27_115#_M1007_d N_B1_M1007_g N_Y_M1002_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_A0_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1006_d N_A1_M1006_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.2205 AS=0.1323 PD=1.61 PS=1.47 NRD=5.4569 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 A_282_521# N_B0_M1005_g N_Y_M1006_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2205 PD=1.47 PS=1.61 NRD=7.8012 NRS=5.4569 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B1_M1004_g A_282_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=4.87485 P=8.85
pX9_noxref noxref_11 A0 A0 PROBETYPE=1
pX10_noxref noxref_12 A1 A1 PROBETYPE=1
pX11_noxref noxref_13 B0 B0 PROBETYPE=1
pX12_noxref noxref_14 Y Y PROBETYPE=1
pX13_noxref noxref_15 B1 B1 PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__oai22_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__or2_1.spice
* Created: Mon Nov 16 20:41:20 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__or2_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_1  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_A_27_521#_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_A_27_521#_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_27_521#_M1002_g N_GND_M1001_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_A_M1004_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_521#_M1005_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9449 P=7.95
pX7_noxref noxref_8 B B PROBETYPE=1
pX8_noxref noxref_9 A A PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__or2_2.spice
* Created: Mon Nov 16 20:41:26 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__or2_2.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_2  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1004 N_A_27_521#_M1004_d N_B_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_A_27_521#_M1004_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_27_521#_M1002_g N_GND_M1001_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_Y_M1002_d N_A_27_521#_M1007_g N_GND_M1007_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75001.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_M1005_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1005_d N_A_27_521#_M1003_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_A_27_521#_M1006_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=4.8513 P=8.83
pX9_noxref noxref_8 B B PROBETYPE=1
pX10_noxref noxref_9 A A PROBETYPE=1
pX11_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_2.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__or2_4.spice
* Created: Mon Nov 16 20:41:32 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__or2_4.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_4  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1004 N_A_27_521#_M1004_d N_B_M1004_g N_GND_M1004_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1001 N_GND_M1001_d N_A_M1001_g N_A_27_521#_M1004_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1002 N_Y_M1002_d N_A_27_521#_M1002_g N_GND_M1001_d N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1002_d N_A_27_521#_M1009_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1010 N_Y_M1010_d N_A_27_521#_M1010_g N_GND_M1009_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1010_d N_A_27_521#_M1011_g N_GND_M1011_s N_GND_M1004_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.3 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.3 A=0.189 P=2.82 MULT=1
MM1007 N_VDD_M1007_d N_A_M1007_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_VDD_M1007_d N_A_27_521#_M1003_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_27_521#_M1005_g N_Y_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1005_d N_A_27_521#_M1006_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_VDD_M1008_d N_A_27_521#_M1008_g N_Y_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1004_b N_VDD_M1000_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_8 B B PROBETYPE=1
pX14_noxref noxref_9 A A PROBETYPE=1
pX15_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_4.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__or2_8.spice
* Created: Mon Nov 16 20:41:37 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__or2_8.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_8  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1008 N_A_27_521#_M1008_d N_B_M1008_g N_GND_M1008_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75004.1 A=0.0825 P=1.4 MULT=1
MM1002 N_GND_M1002_d N_A_M1002_g N_A_27_521#_M1008_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75003.6 A=0.0825 P=1.4 MULT=1
MM1004 N_Y_M1004_d N_A_27_521#_M1004_g N_GND_M1002_d N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.1
+ SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1009 N_Y_M1004_d N_A_27_521#_M1009_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.5
+ SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1012 N_Y_M1012_d N_A_27_521#_M1012_g N_GND_M1009_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75001.9
+ SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1015 N_Y_M1012_d N_A_27_521#_M1015_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.3
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1016 N_Y_M1016_d N_A_27_521#_M1016_g N_GND_M1015_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75002.8
+ SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1017 N_Y_M1016_d N_A_27_521#_M1017_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.2
+ SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1018 N_Y_M1018_d N_A_27_521#_M1018_g N_GND_M1017_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.077 PD=0.83 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667 SA=75003.6
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1019 N_Y_M1018_d N_A_27_521#_M1019_g N_GND_M1019_s N_GND_M1008_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75004.1 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 A_110_521# N_B_M1000_g N_A_27_521#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75004.1 A=0.189 P=2.82 MULT=1
MM1013 N_VDD_M1013_d N_A_M1013_g A_110_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=13.2778 M=1 R=8.4 SA=75000.6
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_27_521#_M1001_g N_VDD_M1013_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1003 N_Y_M1001_d N_A_27_521#_M1003_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_521#_M1005_g N_VDD_M1003_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_27_521#_M1006_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1007_d N_A_27_521#_M1007_g N_VDD_M1006_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1007_d N_A_27_521#_M1010_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_A_27_521#_M1011_g N_VDD_M1010_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1011_d N_A_27_521#_M1014_g N_VDD_M1014_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref N_GND_M1008_b N_VDD_M1000_b NWDIODE A=10.2897 P=14.11
pX21_noxref noxref_8 B B PROBETYPE=1
pX22_noxref noxref_9 A A PROBETYPE=1
pX23_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_8.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__or2_l.spice
* Created: Mon Nov 16 20:41:43 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__or2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__or2_l  GND VDD B A Y
*
* Y	Y
* A	A
* B	B
* VDD	VDD
* GND	GND
MM1003 N_A_27_605#_M1003_d N_B_M1003_g N_GND_M1003_s N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_GND_M1000_d N_A_M1000_g N_A_27_605#_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_27_605#_M1001_g N_GND_M1000_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_110_605# N_B_M1002_g N_A_27_605#_M1002_s N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=19.9167 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_VDD_M1004_d N_A_M1004_g A_110_605# N_VDD_M1002_b PSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=19.9167 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1005_d N_A_27_605#_M1005_g N_VDD_M1004_d N_VDD_M1002_b PSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1002_b NWDIODE A=3.23635 P=7.21
pX7_noxref noxref_8 B B PROBETYPE=1
pX8_noxref noxref_9 A A PROBETYPE=1
pX9_noxref noxref_10 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__or2_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__pcgate_1.spice
* Created: Tue Apr 26 09:50:31 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__pcgate_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__pcgate_1  GND VDD SE E CK Q ECK
*
* ECK	ECK
* Q	Q
* CK	CK
* E	E
* SE	SE
* VDD	VDD
* GND	GND
MM1012 N_A_N233_521#_M1012_d N_SE_M1012_g N_GND_M1012_s N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1019 N_GND_M1019_d N_E_M1019_g N_A_N233_521#_M1012_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1025 N_GND_M1025_d N_A_86_241#_M1025_g N_A_43_115#_M1025_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1023 A_212_115# N_A_N233_521#_M1023_g N_GND_M1025_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1020 N_A_86_241#_M1020_d N_A_254_89#_M1020_g A_212_115# N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1013 A_404_115# N_CK_M1013_g N_A_86_241#_M1020_d N_GND_M1012_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_43_115#_M1007_g A_404_115# N_GND_M1012_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_A_254_89#_M1008_d N_CK_M1008_g N_GND_M1007_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1018 N_GND_M1018_d N_A_43_115#_M1018_g N_A_687_115#_M1018_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1010 N_Q_M1010_d N_A_687_115#_M1010_g N_GND_M1018_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1017 A_1046_115# N_A_687_115#_M1017_g N_A_963_115#_M1017_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1014 N_GND_M1014_d N_CK_M1014_g A_1046_115# N_GND_M1012_b NLOWVT L=0.15 W=0.52
+ AD=0.091 AS=0.0546 PD=0.87 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667 SA=75000.5
+ SB=75000.7 A=0.078 P=1.34 MULT=1
MM1011 N_ECK_M1011_d N_A_963_115#_M1011_g N_GND_M1014_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.091 PD=1.57 PS=0.87 NRD=0 NRS=16.152 M=1
+ R=3.46667 SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 A_N150_521# N_SE_M1001_g N_A_N233_521#_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_E_M1004_g A_N150_521# N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1016 N_VDD_M1016_d N_A_86_241#_M1016_g N_A_43_115#_M1016_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1015 A_212_521# N_A_N233_521#_M1015_g N_VDD_M1016_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_A_86_241#_M1009_d N_CK_M1009_g A_212_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 A_404_521# N_A_254_89#_M1002_g N_A_86_241#_M1009_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1021 N_VDD_M1021_d N_A_43_115#_M1021_g A_404_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_254_89#_M1022_d N_CK_M1022_g N_VDD_M1021_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_43_115#_M1005_g N_A_687_115#_M1005_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_Q_M1024_d N_A_687_115#_M1024_g N_VDD_M1005_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_963_115#_M1003_d N_A_687_115#_M1003_g N_VDD_M1003_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_CK_M1006_g N_A_963_115#_M1003_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_ECK_M1000_d N_A_963_115#_M1000_g N_VDD_M1006_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1012_b N_VDD_M1001_b NWDIODE A=16.3422 P=19.99
pX27_noxref noxref_20 N_SE_X27_noxref_CONDUCTOR SE PROBETYPE=1
pX28_noxref noxref_21 E E PROBETYPE=1
pX29_noxref noxref_22 CK CK PROBETYPE=1
pX30_noxref noxref_23 Q Q PROBETYPE=1
pX31_noxref noxref_24 ECK ECK PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__pcgate_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__pcgateCKa_new.spice
* Created: Tue Apr 26 09:50:40 2022
* Program "Calibre xRC"
* Version "v2021.2_28.15"
*
.include "sky130_osu_sc_12T_hs__pcgateCKa_new.pex.spice"
.subckt sky130_osu_sc_12T_hs__pcgateCKa_new  GND VDD SE E CK CKA Q ECK
*
* ECK	ECK
* Q	Q
* CKA	CKA
* CK	CK
* E	E
* SE	SE
* VDD	VDD
* GND	GND
MM1012 N_A_N233_521#_M1012_d N_SE_M1012_g N_GND_M1012_s N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1019 N_GND_M1019_d N_E_M1019_g N_A_N233_521#_M1012_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1025 N_GND_M1025_d N_A_86_241#_M1025_g N_A_43_115#_M1025_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75002.4 A=0.078 P=1.34 MULT=1
MM1023 A_212_115# N_A_N233_521#_M1023_g N_GND_M1025_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.0546 AS=0.0728 PD=0.73 PS=0.8 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75001.9 A=0.078 P=1.34 MULT=1
MM1020 N_A_86_241#_M1020_d N_A_254_89#_M1020_g A_212_115# N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.117 AS=0.0546 PD=0.97 PS=0.73 NRD=19.608 NRS=11.532 M=1
+ R=3.46667 SA=75001 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1013 A_404_115# N_CK_M1013_g N_A_86_241#_M1020_d N_GND_M1012_b NLOWVT L=0.15
+ W=0.52 AD=0.0546 AS=0.117 PD=0.73 PS=0.97 NRD=11.532 NRS=19.608 M=1 R=3.46667
+ SA=75001.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1007 N_GND_M1007_d N_A_43_115#_M1007_g A_404_115# N_GND_M1012_b NLOWVT L=0.15
+ W=0.52 AD=0.0728 AS=0.0546 PD=0.8 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75001.9 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1008 N_A_254_89#_M1008_d N_CK_M1008_g N_GND_M1007_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75002.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1018 N_GND_M1018_d N_A_43_115#_M1018_g N_A_687_115#_M1018_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0728 AS=0.1378 PD=0.8 PS=1.57 NRD=0 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1010 N_Q_M1010_d N_A_687_115#_M1010_g N_GND_M1018_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.0728 PD=1.57 PS=0.8 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1017 A_1046_115# N_A_687_115#_M1017_g N_A_963_115#_M1017_s N_GND_M1012_b
+ NLOWVT L=0.15 W=0.52 AD=0.0546 AS=0.1378 PD=0.73 PS=1.57 NRD=11.532 NRS=0 M=1
+ R=3.46667 SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1014 N_GND_M1014_d N_CKA_M1014_g A_1046_115# N_GND_M1012_b NLOWVT L=0.15
+ W=0.52 AD=0.091 AS=0.0546 PD=0.87 PS=0.73 NRD=0 NRS=11.532 M=1 R=3.46667
+ SA=75000.5 SB=75000.7 A=0.078 P=1.34 MULT=1
MM1011 N_ECK_M1011_d N_A_963_115#_M1011_g N_GND_M1014_d N_GND_M1012_b NLOWVT
+ L=0.15 W=0.52 AD=0.1378 AS=0.091 PD=1.57 PS=0.87 NRD=0 NRS=16.152 M=1
+ R=3.46667 SA=75001 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1001 A_N150_521# N_SE_M1001_g N_A_N233_521#_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_E_M1004_g A_N150_521# N_VDD_M1001_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1016 N_VDD_M1016_d N_A_86_241#_M1016_g N_A_43_115#_M1016_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1015 A_212_521# N_A_N233_521#_M1015_g N_VDD_M1016_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_A_86_241#_M1009_d N_CK_M1009_g A_212_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 A_404_521# N_A_254_89#_M1002_g N_A_86_241#_M1009_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1
+ R=8.4 SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1021 N_VDD_M1021_d N_A_43_115#_M1021_g A_404_521# N_VDD_M1001_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_254_89#_M1022_d N_CK_M1022_g N_VDD_M1021_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_VDD_M1005_d N_A_43_115#_M1005_g N_A_687_115#_M1005_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1024 N_Q_M1024_d N_A_687_115#_M1024_g N_VDD_M1005_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_A_963_115#_M1003_d N_A_687_115#_M1003_g N_VDD_M1003_s N_VDD_M1001_b
+ PSHORT L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VDD_M1006_d N_CKA_M1006_g N_A_963_115#_M1003_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_ECK_M1000_d N_A_963_115#_M1000_g N_VDD_M1006_d N_VDD_M1001_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref N_GND_M1012_b N_VDD_M1001_b NWDIODE A=16.3422 P=19.99
pX27_noxref noxref_21 N_SE_X27_noxref_CONDUCTOR SE PROBETYPE=1
pX28_noxref noxref_22 E E PROBETYPE=1
pX29_noxref noxref_23 CK CK PROBETYPE=1
pX30_noxref noxref_24 Q Q PROBETYPE=1
pX31_noxref noxref_25 Q Q PROBETYPE=1
pX32_noxref noxref_26 CKA CKA PROBETYPE=1
pX33_noxref noxref_27 ECK ECK PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__pcgateCKa_new.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tbufi_1.spice
* Created: Mon Nov 16 20:41:49 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tbufi_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__tbufi_1  GND VDD OE A Y
*
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_OE_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1001 A_196_115# N_OE_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_196_115# N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_OE_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1004 A_196_521# N_A_27_115#_M1004_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_196_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9552 P=7.96
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tbufi_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tbufi_l.spice
* Created: Mon Nov 16 20:41:55 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tbufi_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__tbufi_l  GND VDD OE A Y
*
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_196_115# N_OE_M1000_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_115# N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VDD_M1001_d N_OE_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1005 A_196_605# N_A_27_115#_M1005_g N_VDD_M1001_d N_VDD_M1001_b PSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_196_605# N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=3.2448 P=7.22
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tbufi_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tiehi.spice
* Created: Mon Nov 16 20:42:00 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tiehi.pex.spice"
.subckt sky130_osu_sc_12T_hs__tiehi  GND VDD Y
*
* Y	Y
* VDD	VDD
* GND	GND
MM1001 N_A_80_89#_M1001_d N_A_80_89#_M1001_g N_GND_M1001_s N_GND_M1001_b NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_Y_M1000_d N_A_80_89#_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.1424 P=6.2
pX3_noxref noxref_5 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tiehi.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tielo.spice
* Created: Mon Nov 16 20:42:06 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tielo.pex.spice"
.subckt sky130_osu_sc_12T_hs__tielo  GND VDD Y
*
* Y	Y
* VDD	VDD
* GND	GND
MM1001 N_Y_M1001_d N_A_80_89#_M1001_g N_GND_M1001_s N_GND_M1001_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.14575 PD=1.63 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_80_89#_M1000_d N_A_80_89#_M1000_g N_VDD_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX2_noxref N_GND_M1001_b N_VDD_M1000_b NWDIODE A=2.1424 P=6.2
pX3_noxref noxref_5 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tielo.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tnbufi_1.spice
* Created: Mon Nov 16 20:42:12 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tnbufi_1.pex.spice"
.subckt sky130_osu_sc_12T_hs__tnbufi_1  GND VDD OE A Y
*
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1003 N_GND_M1003_d N_OE_M1003_g N_A_27_115#_M1003_s N_GND_M1003_b NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1001 A_196_115# N_A_27_115#_M1001_g N_GND_M1003_d N_GND_M1003_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.5 A=0.0825 P=1.4 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g A_196_115# N_GND_M1003_b NLOWVT L=0.15 W=0.55
+ AD=0.14575 AS=0.05775 PD=1.63 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_OE_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001 A=0.189 P=2.82 MULT=1
MM1004 A_196_521# N_OE_M1004_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_196_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX6_noxref N_GND_M1003_b N_VDD_M1000_b NWDIODE A=3.9552 P=7.96
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tnbufi_1.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__tnbufi_l.spice
* Created: Mon Nov 16 20:42:17 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__tnbufi_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__tnbufi_l  GND VDD OE A Y
*
* Y	Y
* A	A
* OE	OE
* VDD	VDD
* GND	GND
MM1002 N_GND_M1002_d N_OE_M1002_g N_A_27_115#_M1002_s N_GND_M1002_b NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_196_115# N_A_27_115#_M1000_g N_GND_M1002_d N_GND_M1002_b NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_196_115# N_GND_M1002_b NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VDD_M1001_d N_OE_M1001_g N_A_27_115#_M1001_s N_VDD_M1001_b PSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001 A=0.126 P=1.98 MULT=1
MM1005 A_196_605# N_OE_M1005_g N_VDD_M1001_d N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1176 PD=1.05 PS=1.12 NRD=11.7215 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g A_196_605# N_VDD_M1001_b PSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6 SA=75001
+ SB=75000.2 A=0.126 P=1.98 MULT=1
DX6_noxref N_GND_M1002_b N_VDD_M1001_b NWDIODE A=3.2448 P=7.22
pX7_noxref noxref_9 OE OE PROBETYPE=1
pX8_noxref noxref_10 A A PROBETYPE=1
pX9_noxref noxref_11 Y Y PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__tnbufi_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__xnor2_l.spice
* Created: Mon Nov 16 20:42:23 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__xnor2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__xnor2_l  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_A_M1006_g N_A_27_115#_M1006_s N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1002 A_196_115# N_A_M1002_g N_GND_M1006_d N_GND_M1006_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667 SA=75000.6
+ SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1011_d N_A_238_89#_M1011_g A_196_115# N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75001 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1008 A_388_115# N_A_27_115#_M1008_g N_Y_M1011_d N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.6 SB=75001 A=0.0825 P=1.4 MULT=1
MM1010 N_GND_M1010_d N_B_M1010_g A_388_115# N_GND_M1006_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_A_238_89#_M1007_d N_B_M1007_g N_GND_M1010_d N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1009 A_196_521# N_A_27_115#_M1009_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_238_89#_M1005_g A_196_521# N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1003 A_388_521# N_A_M1003_g N_Y_M1005_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B_M1004_g A_388_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_238_89#_M1001_d N_B_M1001_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1006_b N_VDD_M1000_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_12 A A PROBETYPE=1
pX14_noxref noxref_13 Y Y PROBETYPE=1
pX15_noxref noxref_14 B B PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__xnor2_l.pxi.spice"
*
.ends
*
*


* File: sky130_osu_sc_12T_hs__xor2_l.spice
* Created: Mon Nov 16 20:42:29 2020
* Program "Calibre xRC"
* Version "v2020.2_35.23"
*
.include "sky130_osu_sc_12T_hs__xor2_l.pex.spice"
.subckt sky130_osu_sc_12T_hs__xor2_l  GND VDD A B Y
*
* Y	Y
* B	B
* A	A
* VDD	VDD
* GND	GND
MM1006 N_GND_M1006_d N_A_M1006_g N_A_27_115#_M1006_s N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.14575 PD=0.83 PS=1.63 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.4 A=0.0825 P=1.4 MULT=1
MM1002 A_196_115# N_A_27_115#_M1002_g N_GND_M1006_d N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.05775 AS=0.077 PD=0.76 PS=0.83 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1011 N_Y_M1011_d N_A_238_89#_M1011_g A_196_115# N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.12375 AS=0.05775 PD=1 PS=0.76 NRD=18.54 NRS=10.908 M=1 R=3.66667
+ SA=75001 SB=75001.6 A=0.0825 P=1.4 MULT=1
MM1008 A_388_115# N_A_M1008_g N_Y_M1011_d N_GND_M1006_b NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.12375 PD=0.76 PS=1 NRD=10.908 NRS=18.54 M=1 R=3.66667
+ SA=75001.6 SB=75001 A=0.0825 P=1.4 MULT=1
MM1010 N_GND_M1010_d N_B_M1010_g A_388_115# N_GND_M1006_b NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.05775 PD=0.83 PS=0.76 NRD=0 NRS=10.908 M=1 R=3.66667 SA=75001.9
+ SB=75000.6 A=0.0825 P=1.4 MULT=1
MM1007 N_A_238_89#_M1007_d N_B_M1007_g N_GND_M1010_d N_GND_M1006_b NLOWVT L=0.15
+ W=0.55 AD=0.14575 AS=0.077 PD=1.63 PS=0.83 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75002.4 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1000 N_VDD_M1000_d N_A_M1000_g N_A_27_115#_M1000_s N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1009 A_196_521# N_A_M1009_g N_VDD_M1000_d N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1323 AS=0.1764 PD=1.47 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_238_89#_M1005_g A_196_521# N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.2835 AS=0.1323 PD=1.71 PS=1.47 NRD=13.2778 NRS=7.8012 M=1 R=8.4
+ SA=75001 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1003 A_388_521# N_A_27_115#_M1003_g N_Y_M1005_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.1323 AS=0.2835 PD=1.47 PS=1.71 NRD=7.8012 NRS=13.2778 M=1 R=8.4
+ SA=75001.6 SB=75001 A=0.189 P=2.82 MULT=1
MM1004 N_VDD_M1004_d N_B_M1004_g A_388_521# N_VDD_M1000_b PSHORT L=0.15 W=1.26
+ AD=0.1764 AS=0.1323 PD=1.54 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1001 N_A_238_89#_M1001_d N_B_M1001_g N_VDD_M1004_d N_VDD_M1000_b PSHORT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref N_GND_M1006_b N_VDD_M1000_b NWDIODE A=6.6641 P=10.59
pX13_noxref noxref_12 A A PROBETYPE=1
pX14_noxref noxref_13 Y Y PROBETYPE=1
pX15_noxref noxref_14 B B PROBETYPE=1
*
.include "sky130_osu_sc_12T_hs__xor2_l.pxi.spice"
*
.ends
*
*


.subckt sky130_osu_sc_12T_hs__fill_1  GND VDD
.ends

.subckt sky130_osu_sc_12T_hs__fill_2  GND VDD
.ends

.subckt sky130_osu_sc_12T_hs__fill_4  GND VDD
.ends

.subckt sky130_osu_sc_12T_hs__fill_8  GND VDD
.ends

.subckt sky130_osu_sc_12T_hs__fill_16  GND VDD
.ends

.subckt sky130_osu_sc_12T_hs__fill_32  GND VDD
.ends
