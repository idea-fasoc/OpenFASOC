* NGSPICE file created from diff_pair_sample_0635.ext - technology: sky130A

.subckt diff_pair_sample_0635 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0.56925 ps=3.78 w=3.45 l=0.78
X1 VDD2.t5 VN.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0.56925 ps=3.78 w=3.45 l=0.78
X2 VDD2.t4 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=1.3455 ps=7.68 w=3.45 l=0.78
X3 VTAIL.t6 VP.t1 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.78
X4 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.78
X5 VDD1.t3 VP.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=1.3455 ps=7.68 w=3.45 l=0.78
X6 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.78
X7 VTAIL.t11 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.78
X8 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0.56925 ps=3.78 w=3.45 l=0.78
X9 VDD2.t2 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=1.3455 ps=7.68 w=3.45 l=0.78
X10 VTAIL.t3 VN.t4 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.78
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.78
X12 VDD1.t1 VP.t4 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=1.3455 ps=7.68 w=3.45 l=0.78
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0 ps=0 w=3.45 l=0.78
X14 VDD1.t0 VP.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=1.3455 pd=7.68 as=0.56925 ps=3.78 w=3.45 l=0.78
X15 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.56925 pd=3.78 as=0.56925 ps=3.78 w=3.45 l=0.78
R0 VP.n3 VP.t0 180.388
R1 VP.n15 VP.n14 161.3
R2 VP.n5 VP.n2 161.3
R3 VP.n7 VP.n6 161.3
R4 VP.n13 VP.n0 161.3
R5 VP.n12 VP.n11 161.3
R6 VP.n10 VP.n1 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n8 VP.t5 157.268
R9 VP.n12 VP.t1 157.268
R10 VP.n14 VP.t2 157.268
R11 VP.n6 VP.t4 157.268
R12 VP.n4 VP.t3 157.268
R13 VP.n3 VP.n2 44.8847
R14 VP.n9 VP.n7 35.1179
R15 VP.n8 VP.n1 32.1338
R16 VP.n14 VP.n13 32.1338
R17 VP.n6 VP.n5 32.1338
R18 VP.n4 VP.n3 18.6308
R19 VP.n12 VP.n1 16.0672
R20 VP.n13 VP.n12 16.0672
R21 VP.n5 VP.n4 16.0672
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VTAIL.n7 VTAIL.t1 63.8391
R29 VTAIL.n11 VTAIL.t5 63.839
R30 VTAIL.n2 VTAIL.t7 63.839
R31 VTAIL.n10 VTAIL.t8 63.839
R32 VTAIL.n9 VTAIL.n8 58.1
R33 VTAIL.n6 VTAIL.n5 58.1
R34 VTAIL.n1 VTAIL.n0 58.0998
R35 VTAIL.n4 VTAIL.n3 58.0998
R36 VTAIL.n6 VTAIL.n4 17.2548
R37 VTAIL.n11 VTAIL.n10 16.2979
R38 VTAIL.n0 VTAIL.t0 5.73963
R39 VTAIL.n0 VTAIL.t3 5.73963
R40 VTAIL.n3 VTAIL.t9 5.73963
R41 VTAIL.n3 VTAIL.t6 5.73963
R42 VTAIL.n8 VTAIL.t10 5.73963
R43 VTAIL.n8 VTAIL.t11 5.73963
R44 VTAIL.n5 VTAIL.t4 5.73963
R45 VTAIL.n5 VTAIL.t2 5.73963
R46 VTAIL.n7 VTAIL.n6 0.957397
R47 VTAIL.n10 VTAIL.n9 0.957397
R48 VTAIL.n4 VTAIL.n2 0.957397
R49 VTAIL.n9 VTAIL.n7 0.948776
R50 VTAIL.n2 VTAIL.n1 0.948776
R51 VTAIL VTAIL.n11 0.659983
R52 VTAIL VTAIL.n1 0.297914
R53 VDD1 VDD1.t5 81.2937
R54 VDD1.n1 VDD1.t0 81.1802
R55 VDD1.n1 VDD1.n0 74.9625
R56 VDD1.n3 VDD1.n2 74.7787
R57 VDD1.n3 VDD1.n1 30.8608
R58 VDD1.n2 VDD1.t2 5.73963
R59 VDD1.n2 VDD1.t1 5.73963
R60 VDD1.n0 VDD1.t4 5.73963
R61 VDD1.n0 VDD1.t3 5.73963
R62 VDD1 VDD1.n3 0.181534
R63 B.n397 B.n396 585
R64 B.n398 B.n397 585
R65 B.n152 B.n63 585
R66 B.n151 B.n150 585
R67 B.n149 B.n148 585
R68 B.n147 B.n146 585
R69 B.n145 B.n144 585
R70 B.n143 B.n142 585
R71 B.n141 B.n140 585
R72 B.n139 B.n138 585
R73 B.n137 B.n136 585
R74 B.n135 B.n134 585
R75 B.n133 B.n132 585
R76 B.n131 B.n130 585
R77 B.n129 B.n128 585
R78 B.n127 B.n126 585
R79 B.n125 B.n124 585
R80 B.n123 B.n122 585
R81 B.n121 B.n120 585
R82 B.n119 B.n118 585
R83 B.n117 B.n116 585
R84 B.n115 B.n114 585
R85 B.n113 B.n112 585
R86 B.n111 B.n110 585
R87 B.n109 B.n108 585
R88 B.n107 B.n106 585
R89 B.n105 B.n104 585
R90 B.n102 B.n101 585
R91 B.n100 B.n99 585
R92 B.n98 B.n97 585
R93 B.n96 B.n95 585
R94 B.n94 B.n93 585
R95 B.n92 B.n91 585
R96 B.n90 B.n89 585
R97 B.n88 B.n87 585
R98 B.n86 B.n85 585
R99 B.n84 B.n83 585
R100 B.n82 B.n81 585
R101 B.n80 B.n79 585
R102 B.n78 B.n77 585
R103 B.n76 B.n75 585
R104 B.n74 B.n73 585
R105 B.n72 B.n71 585
R106 B.n70 B.n69 585
R107 B.n395 B.n41 585
R108 B.n399 B.n41 585
R109 B.n394 B.n40 585
R110 B.n400 B.n40 585
R111 B.n393 B.n392 585
R112 B.n392 B.n36 585
R113 B.n391 B.n35 585
R114 B.n406 B.n35 585
R115 B.n390 B.n34 585
R116 B.n407 B.n34 585
R117 B.n389 B.n33 585
R118 B.n408 B.n33 585
R119 B.n388 B.n387 585
R120 B.n387 B.n29 585
R121 B.n386 B.n28 585
R122 B.n414 B.n28 585
R123 B.n385 B.n27 585
R124 B.n415 B.n27 585
R125 B.n384 B.n26 585
R126 B.n416 B.n26 585
R127 B.n383 B.n382 585
R128 B.n382 B.n22 585
R129 B.n381 B.n21 585
R130 B.n422 B.n21 585
R131 B.n380 B.n20 585
R132 B.n423 B.n20 585
R133 B.n379 B.n19 585
R134 B.n424 B.n19 585
R135 B.n378 B.n377 585
R136 B.n377 B.n18 585
R137 B.n376 B.n14 585
R138 B.n430 B.n14 585
R139 B.n375 B.n13 585
R140 B.n431 B.n13 585
R141 B.n374 B.n12 585
R142 B.n432 B.n12 585
R143 B.n373 B.n372 585
R144 B.n372 B.n8 585
R145 B.n371 B.n7 585
R146 B.n438 B.n7 585
R147 B.n370 B.n6 585
R148 B.n439 B.n6 585
R149 B.n369 B.n5 585
R150 B.n440 B.n5 585
R151 B.n368 B.n367 585
R152 B.n367 B.n4 585
R153 B.n366 B.n153 585
R154 B.n366 B.n365 585
R155 B.n356 B.n154 585
R156 B.n155 B.n154 585
R157 B.n358 B.n357 585
R158 B.n359 B.n358 585
R159 B.n355 B.n160 585
R160 B.n160 B.n159 585
R161 B.n354 B.n353 585
R162 B.n353 B.n352 585
R163 B.n162 B.n161 585
R164 B.n345 B.n162 585
R165 B.n344 B.n343 585
R166 B.n346 B.n344 585
R167 B.n342 B.n167 585
R168 B.n167 B.n166 585
R169 B.n341 B.n340 585
R170 B.n340 B.n339 585
R171 B.n169 B.n168 585
R172 B.n170 B.n169 585
R173 B.n332 B.n331 585
R174 B.n333 B.n332 585
R175 B.n330 B.n175 585
R176 B.n175 B.n174 585
R177 B.n329 B.n328 585
R178 B.n328 B.n327 585
R179 B.n177 B.n176 585
R180 B.n178 B.n177 585
R181 B.n320 B.n319 585
R182 B.n321 B.n320 585
R183 B.n318 B.n182 585
R184 B.n186 B.n182 585
R185 B.n317 B.n316 585
R186 B.n316 B.n315 585
R187 B.n184 B.n183 585
R188 B.n185 B.n184 585
R189 B.n308 B.n307 585
R190 B.n309 B.n308 585
R191 B.n306 B.n191 585
R192 B.n191 B.n190 585
R193 B.n300 B.n299 585
R194 B.n298 B.n214 585
R195 B.n297 B.n213 585
R196 B.n302 B.n213 585
R197 B.n296 B.n295 585
R198 B.n294 B.n293 585
R199 B.n292 B.n291 585
R200 B.n290 B.n289 585
R201 B.n288 B.n287 585
R202 B.n286 B.n285 585
R203 B.n284 B.n283 585
R204 B.n282 B.n281 585
R205 B.n280 B.n279 585
R206 B.n278 B.n277 585
R207 B.n276 B.n275 585
R208 B.n274 B.n273 585
R209 B.n272 B.n271 585
R210 B.n270 B.n269 585
R211 B.n268 B.n267 585
R212 B.n266 B.n265 585
R213 B.n264 B.n263 585
R214 B.n262 B.n261 585
R215 B.n260 B.n259 585
R216 B.n258 B.n257 585
R217 B.n256 B.n255 585
R218 B.n254 B.n253 585
R219 B.n252 B.n251 585
R220 B.n249 B.n248 585
R221 B.n247 B.n246 585
R222 B.n245 B.n244 585
R223 B.n243 B.n242 585
R224 B.n241 B.n240 585
R225 B.n239 B.n238 585
R226 B.n237 B.n236 585
R227 B.n235 B.n234 585
R228 B.n233 B.n232 585
R229 B.n231 B.n230 585
R230 B.n229 B.n228 585
R231 B.n227 B.n226 585
R232 B.n225 B.n224 585
R233 B.n223 B.n222 585
R234 B.n221 B.n220 585
R235 B.n193 B.n192 585
R236 B.n305 B.n304 585
R237 B.n189 B.n188 585
R238 B.n190 B.n189 585
R239 B.n311 B.n310 585
R240 B.n310 B.n309 585
R241 B.n312 B.n187 585
R242 B.n187 B.n185 585
R243 B.n314 B.n313 585
R244 B.n315 B.n314 585
R245 B.n181 B.n180 585
R246 B.n186 B.n181 585
R247 B.n323 B.n322 585
R248 B.n322 B.n321 585
R249 B.n324 B.n179 585
R250 B.n179 B.n178 585
R251 B.n326 B.n325 585
R252 B.n327 B.n326 585
R253 B.n173 B.n172 585
R254 B.n174 B.n173 585
R255 B.n335 B.n334 585
R256 B.n334 B.n333 585
R257 B.n336 B.n171 585
R258 B.n171 B.n170 585
R259 B.n338 B.n337 585
R260 B.n339 B.n338 585
R261 B.n165 B.n164 585
R262 B.n166 B.n165 585
R263 B.n348 B.n347 585
R264 B.n347 B.n346 585
R265 B.n349 B.n163 585
R266 B.n345 B.n163 585
R267 B.n351 B.n350 585
R268 B.n352 B.n351 585
R269 B.n158 B.n157 585
R270 B.n159 B.n158 585
R271 B.n361 B.n360 585
R272 B.n360 B.n359 585
R273 B.n362 B.n156 585
R274 B.n156 B.n155 585
R275 B.n364 B.n363 585
R276 B.n365 B.n364 585
R277 B.n2 B.n0 585
R278 B.n4 B.n2 585
R279 B.n3 B.n1 585
R280 B.n439 B.n3 585
R281 B.n437 B.n436 585
R282 B.n438 B.n437 585
R283 B.n435 B.n9 585
R284 B.n9 B.n8 585
R285 B.n434 B.n433 585
R286 B.n433 B.n432 585
R287 B.n11 B.n10 585
R288 B.n431 B.n11 585
R289 B.n429 B.n428 585
R290 B.n430 B.n429 585
R291 B.n427 B.n15 585
R292 B.n18 B.n15 585
R293 B.n426 B.n425 585
R294 B.n425 B.n424 585
R295 B.n17 B.n16 585
R296 B.n423 B.n17 585
R297 B.n421 B.n420 585
R298 B.n422 B.n421 585
R299 B.n419 B.n23 585
R300 B.n23 B.n22 585
R301 B.n418 B.n417 585
R302 B.n417 B.n416 585
R303 B.n25 B.n24 585
R304 B.n415 B.n25 585
R305 B.n413 B.n412 585
R306 B.n414 B.n413 585
R307 B.n411 B.n30 585
R308 B.n30 B.n29 585
R309 B.n410 B.n409 585
R310 B.n409 B.n408 585
R311 B.n32 B.n31 585
R312 B.n407 B.n32 585
R313 B.n405 B.n404 585
R314 B.n406 B.n405 585
R315 B.n403 B.n37 585
R316 B.n37 B.n36 585
R317 B.n402 B.n401 585
R318 B.n401 B.n400 585
R319 B.n39 B.n38 585
R320 B.n399 B.n39 585
R321 B.n442 B.n441 585
R322 B.n441 B.n440 585
R323 B.n300 B.n189 487.695
R324 B.n69 B.n39 487.695
R325 B.n304 B.n191 487.695
R326 B.n397 B.n41 487.695
R327 B.n218 B.t10 308.678
R328 B.n215 B.t17 308.678
R329 B.n67 B.t14 308.678
R330 B.n64 B.t6 308.678
R331 B.n398 B.n62 256.663
R332 B.n398 B.n61 256.663
R333 B.n398 B.n60 256.663
R334 B.n398 B.n59 256.663
R335 B.n398 B.n58 256.663
R336 B.n398 B.n57 256.663
R337 B.n398 B.n56 256.663
R338 B.n398 B.n55 256.663
R339 B.n398 B.n54 256.663
R340 B.n398 B.n53 256.663
R341 B.n398 B.n52 256.663
R342 B.n398 B.n51 256.663
R343 B.n398 B.n50 256.663
R344 B.n398 B.n49 256.663
R345 B.n398 B.n48 256.663
R346 B.n398 B.n47 256.663
R347 B.n398 B.n46 256.663
R348 B.n398 B.n45 256.663
R349 B.n398 B.n44 256.663
R350 B.n398 B.n43 256.663
R351 B.n398 B.n42 256.663
R352 B.n302 B.n301 256.663
R353 B.n302 B.n194 256.663
R354 B.n302 B.n195 256.663
R355 B.n302 B.n196 256.663
R356 B.n302 B.n197 256.663
R357 B.n302 B.n198 256.663
R358 B.n302 B.n199 256.663
R359 B.n302 B.n200 256.663
R360 B.n302 B.n201 256.663
R361 B.n302 B.n202 256.663
R362 B.n302 B.n203 256.663
R363 B.n302 B.n204 256.663
R364 B.n302 B.n205 256.663
R365 B.n302 B.n206 256.663
R366 B.n302 B.n207 256.663
R367 B.n302 B.n208 256.663
R368 B.n302 B.n209 256.663
R369 B.n302 B.n210 256.663
R370 B.n302 B.n211 256.663
R371 B.n302 B.n212 256.663
R372 B.n303 B.n302 256.663
R373 B.n302 B.n190 170.202
R374 B.n399 B.n398 170.202
R375 B.n310 B.n189 163.367
R376 B.n310 B.n187 163.367
R377 B.n314 B.n187 163.367
R378 B.n314 B.n181 163.367
R379 B.n322 B.n181 163.367
R380 B.n322 B.n179 163.367
R381 B.n326 B.n179 163.367
R382 B.n326 B.n173 163.367
R383 B.n334 B.n173 163.367
R384 B.n334 B.n171 163.367
R385 B.n338 B.n171 163.367
R386 B.n338 B.n165 163.367
R387 B.n347 B.n165 163.367
R388 B.n347 B.n163 163.367
R389 B.n351 B.n163 163.367
R390 B.n351 B.n158 163.367
R391 B.n360 B.n158 163.367
R392 B.n360 B.n156 163.367
R393 B.n364 B.n156 163.367
R394 B.n364 B.n2 163.367
R395 B.n441 B.n2 163.367
R396 B.n441 B.n3 163.367
R397 B.n437 B.n3 163.367
R398 B.n437 B.n9 163.367
R399 B.n433 B.n9 163.367
R400 B.n433 B.n11 163.367
R401 B.n429 B.n11 163.367
R402 B.n429 B.n15 163.367
R403 B.n425 B.n15 163.367
R404 B.n425 B.n17 163.367
R405 B.n421 B.n17 163.367
R406 B.n421 B.n23 163.367
R407 B.n417 B.n23 163.367
R408 B.n417 B.n25 163.367
R409 B.n413 B.n25 163.367
R410 B.n413 B.n30 163.367
R411 B.n409 B.n30 163.367
R412 B.n409 B.n32 163.367
R413 B.n405 B.n32 163.367
R414 B.n405 B.n37 163.367
R415 B.n401 B.n37 163.367
R416 B.n401 B.n39 163.367
R417 B.n214 B.n213 163.367
R418 B.n295 B.n213 163.367
R419 B.n293 B.n292 163.367
R420 B.n289 B.n288 163.367
R421 B.n285 B.n284 163.367
R422 B.n281 B.n280 163.367
R423 B.n277 B.n276 163.367
R424 B.n273 B.n272 163.367
R425 B.n269 B.n268 163.367
R426 B.n265 B.n264 163.367
R427 B.n261 B.n260 163.367
R428 B.n257 B.n256 163.367
R429 B.n253 B.n252 163.367
R430 B.n248 B.n247 163.367
R431 B.n244 B.n243 163.367
R432 B.n240 B.n239 163.367
R433 B.n236 B.n235 163.367
R434 B.n232 B.n231 163.367
R435 B.n228 B.n227 163.367
R436 B.n224 B.n223 163.367
R437 B.n220 B.n193 163.367
R438 B.n308 B.n191 163.367
R439 B.n308 B.n184 163.367
R440 B.n316 B.n184 163.367
R441 B.n316 B.n182 163.367
R442 B.n320 B.n182 163.367
R443 B.n320 B.n177 163.367
R444 B.n328 B.n177 163.367
R445 B.n328 B.n175 163.367
R446 B.n332 B.n175 163.367
R447 B.n332 B.n169 163.367
R448 B.n340 B.n169 163.367
R449 B.n340 B.n167 163.367
R450 B.n344 B.n167 163.367
R451 B.n344 B.n162 163.367
R452 B.n353 B.n162 163.367
R453 B.n353 B.n160 163.367
R454 B.n358 B.n160 163.367
R455 B.n358 B.n154 163.367
R456 B.n366 B.n154 163.367
R457 B.n367 B.n366 163.367
R458 B.n367 B.n5 163.367
R459 B.n6 B.n5 163.367
R460 B.n7 B.n6 163.367
R461 B.n372 B.n7 163.367
R462 B.n372 B.n12 163.367
R463 B.n13 B.n12 163.367
R464 B.n14 B.n13 163.367
R465 B.n377 B.n14 163.367
R466 B.n377 B.n19 163.367
R467 B.n20 B.n19 163.367
R468 B.n21 B.n20 163.367
R469 B.n382 B.n21 163.367
R470 B.n382 B.n26 163.367
R471 B.n27 B.n26 163.367
R472 B.n28 B.n27 163.367
R473 B.n387 B.n28 163.367
R474 B.n387 B.n33 163.367
R475 B.n34 B.n33 163.367
R476 B.n35 B.n34 163.367
R477 B.n392 B.n35 163.367
R478 B.n392 B.n40 163.367
R479 B.n41 B.n40 163.367
R480 B.n73 B.n72 163.367
R481 B.n77 B.n76 163.367
R482 B.n81 B.n80 163.367
R483 B.n85 B.n84 163.367
R484 B.n89 B.n88 163.367
R485 B.n93 B.n92 163.367
R486 B.n97 B.n96 163.367
R487 B.n101 B.n100 163.367
R488 B.n106 B.n105 163.367
R489 B.n110 B.n109 163.367
R490 B.n114 B.n113 163.367
R491 B.n118 B.n117 163.367
R492 B.n122 B.n121 163.367
R493 B.n126 B.n125 163.367
R494 B.n130 B.n129 163.367
R495 B.n134 B.n133 163.367
R496 B.n138 B.n137 163.367
R497 B.n142 B.n141 163.367
R498 B.n146 B.n145 163.367
R499 B.n150 B.n149 163.367
R500 B.n397 B.n63 163.367
R501 B.n218 B.t13 95.1977
R502 B.n64 B.t8 95.1977
R503 B.n215 B.t19 95.1948
R504 B.n67 B.t15 95.1948
R505 B.n309 B.n190 85.7312
R506 B.n309 B.n185 85.7312
R507 B.n315 B.n185 85.7312
R508 B.n315 B.n186 85.7312
R509 B.n321 B.n178 85.7312
R510 B.n327 B.n178 85.7312
R511 B.n327 B.n174 85.7312
R512 B.n333 B.n174 85.7312
R513 B.n333 B.n170 85.7312
R514 B.n339 B.n170 85.7312
R515 B.n346 B.n166 85.7312
R516 B.n346 B.n345 85.7312
R517 B.n352 B.n159 85.7312
R518 B.n359 B.n159 85.7312
R519 B.n365 B.n155 85.7312
R520 B.n365 B.n4 85.7312
R521 B.n440 B.n4 85.7312
R522 B.n440 B.n439 85.7312
R523 B.n439 B.n438 85.7312
R524 B.n438 B.n8 85.7312
R525 B.n432 B.n431 85.7312
R526 B.n431 B.n430 85.7312
R527 B.n424 B.n18 85.7312
R528 B.n424 B.n423 85.7312
R529 B.n422 B.n22 85.7312
R530 B.n416 B.n22 85.7312
R531 B.n416 B.n415 85.7312
R532 B.n415 B.n414 85.7312
R533 B.n414 B.n29 85.7312
R534 B.n408 B.n29 85.7312
R535 B.n407 B.n406 85.7312
R536 B.n406 B.n36 85.7312
R537 B.n400 B.n36 85.7312
R538 B.n400 B.n399 85.7312
R539 B.n219 B.t12 73.6704
R540 B.n65 B.t9 73.6704
R541 B.n216 B.t18 73.6675
R542 B.n68 B.t16 73.6675
R543 B.n301 B.n300 71.676
R544 B.n295 B.n194 71.676
R545 B.n292 B.n195 71.676
R546 B.n288 B.n196 71.676
R547 B.n284 B.n197 71.676
R548 B.n280 B.n198 71.676
R549 B.n276 B.n199 71.676
R550 B.n272 B.n200 71.676
R551 B.n268 B.n201 71.676
R552 B.n264 B.n202 71.676
R553 B.n260 B.n203 71.676
R554 B.n256 B.n204 71.676
R555 B.n252 B.n205 71.676
R556 B.n247 B.n206 71.676
R557 B.n243 B.n207 71.676
R558 B.n239 B.n208 71.676
R559 B.n235 B.n209 71.676
R560 B.n231 B.n210 71.676
R561 B.n227 B.n211 71.676
R562 B.n223 B.n212 71.676
R563 B.n303 B.n193 71.676
R564 B.n69 B.n42 71.676
R565 B.n73 B.n43 71.676
R566 B.n77 B.n44 71.676
R567 B.n81 B.n45 71.676
R568 B.n85 B.n46 71.676
R569 B.n89 B.n47 71.676
R570 B.n93 B.n48 71.676
R571 B.n97 B.n49 71.676
R572 B.n101 B.n50 71.676
R573 B.n106 B.n51 71.676
R574 B.n110 B.n52 71.676
R575 B.n114 B.n53 71.676
R576 B.n118 B.n54 71.676
R577 B.n122 B.n55 71.676
R578 B.n126 B.n56 71.676
R579 B.n130 B.n57 71.676
R580 B.n134 B.n58 71.676
R581 B.n138 B.n59 71.676
R582 B.n142 B.n60 71.676
R583 B.n146 B.n61 71.676
R584 B.n150 B.n62 71.676
R585 B.n63 B.n62 71.676
R586 B.n149 B.n61 71.676
R587 B.n145 B.n60 71.676
R588 B.n141 B.n59 71.676
R589 B.n137 B.n58 71.676
R590 B.n133 B.n57 71.676
R591 B.n129 B.n56 71.676
R592 B.n125 B.n55 71.676
R593 B.n121 B.n54 71.676
R594 B.n117 B.n53 71.676
R595 B.n113 B.n52 71.676
R596 B.n109 B.n51 71.676
R597 B.n105 B.n50 71.676
R598 B.n100 B.n49 71.676
R599 B.n96 B.n48 71.676
R600 B.n92 B.n47 71.676
R601 B.n88 B.n46 71.676
R602 B.n84 B.n45 71.676
R603 B.n80 B.n44 71.676
R604 B.n76 B.n43 71.676
R605 B.n72 B.n42 71.676
R606 B.n301 B.n214 71.676
R607 B.n293 B.n194 71.676
R608 B.n289 B.n195 71.676
R609 B.n285 B.n196 71.676
R610 B.n281 B.n197 71.676
R611 B.n277 B.n198 71.676
R612 B.n273 B.n199 71.676
R613 B.n269 B.n200 71.676
R614 B.n265 B.n201 71.676
R615 B.n261 B.n202 71.676
R616 B.n257 B.n203 71.676
R617 B.n253 B.n204 71.676
R618 B.n248 B.n205 71.676
R619 B.n244 B.n206 71.676
R620 B.n240 B.n207 71.676
R621 B.n236 B.n208 71.676
R622 B.n232 B.n209 71.676
R623 B.n228 B.n210 71.676
R624 B.n224 B.n211 71.676
R625 B.n220 B.n212 71.676
R626 B.n304 B.n303 71.676
R627 B.n186 B.t11 65.5592
R628 B.t4 B.n166 65.5592
R629 B.n359 B.t1 65.5592
R630 B.n432 B.t0 65.5592
R631 B.n423 B.t5 65.5592
R632 B.t7 B.n407 65.5592
R633 B.n250 B.n219 59.5399
R634 B.n217 B.n216 59.5399
R635 B.n103 B.n68 59.5399
R636 B.n66 B.n65 59.5399
R637 B.n345 B.t2 42.8658
R638 B.n352 B.t2 42.8658
R639 B.n430 B.t3 42.8658
R640 B.n18 B.t3 42.8658
R641 B.n70 B.n38 31.6883
R642 B.n396 B.n395 31.6883
R643 B.n306 B.n305 31.6883
R644 B.n299 B.n188 31.6883
R645 B.n219 B.n218 21.5278
R646 B.n216 B.n215 21.5278
R647 B.n68 B.n67 21.5278
R648 B.n65 B.n64 21.5278
R649 B.n321 B.t11 20.1724
R650 B.n339 B.t4 20.1724
R651 B.t1 B.n155 20.1724
R652 B.t0 B.n8 20.1724
R653 B.t5 B.n422 20.1724
R654 B.n408 B.t7 20.1724
R655 B B.n442 18.0485
R656 B.n71 B.n70 10.6151
R657 B.n74 B.n71 10.6151
R658 B.n75 B.n74 10.6151
R659 B.n78 B.n75 10.6151
R660 B.n79 B.n78 10.6151
R661 B.n82 B.n79 10.6151
R662 B.n83 B.n82 10.6151
R663 B.n86 B.n83 10.6151
R664 B.n87 B.n86 10.6151
R665 B.n90 B.n87 10.6151
R666 B.n91 B.n90 10.6151
R667 B.n94 B.n91 10.6151
R668 B.n95 B.n94 10.6151
R669 B.n98 B.n95 10.6151
R670 B.n99 B.n98 10.6151
R671 B.n102 B.n99 10.6151
R672 B.n107 B.n104 10.6151
R673 B.n108 B.n107 10.6151
R674 B.n111 B.n108 10.6151
R675 B.n112 B.n111 10.6151
R676 B.n115 B.n112 10.6151
R677 B.n116 B.n115 10.6151
R678 B.n119 B.n116 10.6151
R679 B.n120 B.n119 10.6151
R680 B.n124 B.n123 10.6151
R681 B.n127 B.n124 10.6151
R682 B.n128 B.n127 10.6151
R683 B.n131 B.n128 10.6151
R684 B.n132 B.n131 10.6151
R685 B.n135 B.n132 10.6151
R686 B.n136 B.n135 10.6151
R687 B.n139 B.n136 10.6151
R688 B.n140 B.n139 10.6151
R689 B.n143 B.n140 10.6151
R690 B.n144 B.n143 10.6151
R691 B.n147 B.n144 10.6151
R692 B.n148 B.n147 10.6151
R693 B.n151 B.n148 10.6151
R694 B.n152 B.n151 10.6151
R695 B.n396 B.n152 10.6151
R696 B.n307 B.n306 10.6151
R697 B.n307 B.n183 10.6151
R698 B.n317 B.n183 10.6151
R699 B.n318 B.n317 10.6151
R700 B.n319 B.n318 10.6151
R701 B.n319 B.n176 10.6151
R702 B.n329 B.n176 10.6151
R703 B.n330 B.n329 10.6151
R704 B.n331 B.n330 10.6151
R705 B.n331 B.n168 10.6151
R706 B.n341 B.n168 10.6151
R707 B.n342 B.n341 10.6151
R708 B.n343 B.n342 10.6151
R709 B.n343 B.n161 10.6151
R710 B.n354 B.n161 10.6151
R711 B.n355 B.n354 10.6151
R712 B.n357 B.n355 10.6151
R713 B.n357 B.n356 10.6151
R714 B.n356 B.n153 10.6151
R715 B.n368 B.n153 10.6151
R716 B.n369 B.n368 10.6151
R717 B.n370 B.n369 10.6151
R718 B.n371 B.n370 10.6151
R719 B.n373 B.n371 10.6151
R720 B.n374 B.n373 10.6151
R721 B.n375 B.n374 10.6151
R722 B.n376 B.n375 10.6151
R723 B.n378 B.n376 10.6151
R724 B.n379 B.n378 10.6151
R725 B.n380 B.n379 10.6151
R726 B.n381 B.n380 10.6151
R727 B.n383 B.n381 10.6151
R728 B.n384 B.n383 10.6151
R729 B.n385 B.n384 10.6151
R730 B.n386 B.n385 10.6151
R731 B.n388 B.n386 10.6151
R732 B.n389 B.n388 10.6151
R733 B.n390 B.n389 10.6151
R734 B.n391 B.n390 10.6151
R735 B.n393 B.n391 10.6151
R736 B.n394 B.n393 10.6151
R737 B.n395 B.n394 10.6151
R738 B.n299 B.n298 10.6151
R739 B.n298 B.n297 10.6151
R740 B.n297 B.n296 10.6151
R741 B.n296 B.n294 10.6151
R742 B.n294 B.n291 10.6151
R743 B.n291 B.n290 10.6151
R744 B.n290 B.n287 10.6151
R745 B.n287 B.n286 10.6151
R746 B.n286 B.n283 10.6151
R747 B.n283 B.n282 10.6151
R748 B.n282 B.n279 10.6151
R749 B.n279 B.n278 10.6151
R750 B.n278 B.n275 10.6151
R751 B.n275 B.n274 10.6151
R752 B.n274 B.n271 10.6151
R753 B.n271 B.n270 10.6151
R754 B.n267 B.n266 10.6151
R755 B.n266 B.n263 10.6151
R756 B.n263 B.n262 10.6151
R757 B.n262 B.n259 10.6151
R758 B.n259 B.n258 10.6151
R759 B.n258 B.n255 10.6151
R760 B.n255 B.n254 10.6151
R761 B.n254 B.n251 10.6151
R762 B.n249 B.n246 10.6151
R763 B.n246 B.n245 10.6151
R764 B.n245 B.n242 10.6151
R765 B.n242 B.n241 10.6151
R766 B.n241 B.n238 10.6151
R767 B.n238 B.n237 10.6151
R768 B.n237 B.n234 10.6151
R769 B.n234 B.n233 10.6151
R770 B.n233 B.n230 10.6151
R771 B.n230 B.n229 10.6151
R772 B.n229 B.n226 10.6151
R773 B.n226 B.n225 10.6151
R774 B.n225 B.n222 10.6151
R775 B.n222 B.n221 10.6151
R776 B.n221 B.n192 10.6151
R777 B.n305 B.n192 10.6151
R778 B.n311 B.n188 10.6151
R779 B.n312 B.n311 10.6151
R780 B.n313 B.n312 10.6151
R781 B.n313 B.n180 10.6151
R782 B.n323 B.n180 10.6151
R783 B.n324 B.n323 10.6151
R784 B.n325 B.n324 10.6151
R785 B.n325 B.n172 10.6151
R786 B.n335 B.n172 10.6151
R787 B.n336 B.n335 10.6151
R788 B.n337 B.n336 10.6151
R789 B.n337 B.n164 10.6151
R790 B.n348 B.n164 10.6151
R791 B.n349 B.n348 10.6151
R792 B.n350 B.n349 10.6151
R793 B.n350 B.n157 10.6151
R794 B.n361 B.n157 10.6151
R795 B.n362 B.n361 10.6151
R796 B.n363 B.n362 10.6151
R797 B.n363 B.n0 10.6151
R798 B.n436 B.n1 10.6151
R799 B.n436 B.n435 10.6151
R800 B.n435 B.n434 10.6151
R801 B.n434 B.n10 10.6151
R802 B.n428 B.n10 10.6151
R803 B.n428 B.n427 10.6151
R804 B.n427 B.n426 10.6151
R805 B.n426 B.n16 10.6151
R806 B.n420 B.n16 10.6151
R807 B.n420 B.n419 10.6151
R808 B.n419 B.n418 10.6151
R809 B.n418 B.n24 10.6151
R810 B.n412 B.n24 10.6151
R811 B.n412 B.n411 10.6151
R812 B.n411 B.n410 10.6151
R813 B.n410 B.n31 10.6151
R814 B.n404 B.n31 10.6151
R815 B.n404 B.n403 10.6151
R816 B.n403 B.n402 10.6151
R817 B.n402 B.n38 10.6151
R818 B.n104 B.n103 6.5566
R819 B.n120 B.n66 6.5566
R820 B.n267 B.n217 6.5566
R821 B.n251 B.n250 6.5566
R822 B.n103 B.n102 4.05904
R823 B.n123 B.n66 4.05904
R824 B.n270 B.n217 4.05904
R825 B.n250 B.n249 4.05904
R826 B.n442 B.n0 2.81026
R827 B.n442 B.n1 2.81026
R828 VN.n1 VN.t2 180.388
R829 VN.n7 VN.t3 180.388
R830 VN.n5 VN.n4 161.3
R831 VN.n11 VN.n10 161.3
R832 VN.n9 VN.n6 161.3
R833 VN.n3 VN.n0 161.3
R834 VN.n2 VN.t4 157.268
R835 VN.n4 VN.t1 157.268
R836 VN.n8 VN.t5 157.268
R837 VN.n10 VN.t0 157.268
R838 VN.n7 VN.n6 44.8847
R839 VN.n1 VN.n0 44.8847
R840 VN VN.n11 35.4986
R841 VN.n4 VN.n3 32.1338
R842 VN.n10 VN.n9 32.1338
R843 VN.n2 VN.n1 18.6308
R844 VN.n8 VN.n7 18.6308
R845 VN.n3 VN.n2 16.0672
R846 VN.n9 VN.n8 16.0672
R847 VN.n11 VN.n6 0.189894
R848 VN.n5 VN.n0 0.189894
R849 VN VN.n5 0.0516364
R850 VDD2.n1 VDD2.t3 81.1802
R851 VDD2.n2 VDD2.t5 80.5179
R852 VDD2.n1 VDD2.n0 74.9625
R853 VDD2 VDD2.n3 74.9597
R854 VDD2.n2 VDD2.n1 29.7993
R855 VDD2.n3 VDD2.t0 5.73963
R856 VDD2.n3 VDD2.t2 5.73963
R857 VDD2.n0 VDD2.t1 5.73963
R858 VDD2.n0 VDD2.t4 5.73963
R859 VDD2 VDD2.n2 0.776362
C0 VTAIL VP 1.70706f
C1 VDD1 VP 1.7112f
C2 VDD1 VTAIL 4.12379f
C3 VP VDD2 0.308101f
C4 VN VP 3.57856f
C5 VTAIL VDD2 4.16326f
C6 VDD1 VDD2 0.736494f
C7 VN VTAIL 1.69282f
C8 VDD1 VN 0.152812f
C9 VN VDD2 1.55791f
C10 VDD2 B 2.907036f
C11 VDD1 B 3.113028f
C12 VTAIL B 3.105857f
C13 VN B 6.167353f
C14 VP B 5.291111f
C15 VDD2.t3 B 0.453523f
C16 VDD2.t1 B 0.046489f
C17 VDD2.t4 B 0.046489f
C18 VDD2.n0 B 0.356672f
C19 VDD2.n1 B 1.06841f
C20 VDD2.t5 B 0.451856f
C21 VDD2.n2 B 1.07588f
C22 VDD2.t0 B 0.046489f
C23 VDD2.t2 B 0.046489f
C24 VDD2.n3 B 0.356659f
C25 VN.n0 B 0.105649f
C26 VN.t2 B 0.211236f
C27 VN.n1 B 0.096746f
C28 VN.t4 B 0.19735f
C29 VN.n2 B 0.109838f
C30 VN.n3 B 0.005592f
C31 VN.t1 B 0.19735f
C32 VN.n4 B 0.107175f
C33 VN.n5 B 0.019099f
C34 VN.n6 B 0.105649f
C35 VN.t3 B 0.211236f
C36 VN.n7 B 0.096746f
C37 VN.t5 B 0.19735f
C38 VN.n8 B 0.109838f
C39 VN.n9 B 0.005592f
C40 VN.t0 B 0.19735f
C41 VN.n10 B 0.107175f
C42 VN.n11 B 0.755505f
C43 VDD1.t5 B 0.43651f
C44 VDD1.t0 B 0.436184f
C45 VDD1.t4 B 0.044711f
C46 VDD1.t3 B 0.044711f
C47 VDD1.n0 B 0.343036f
C48 VDD1.n1 B 1.07652f
C49 VDD1.t2 B 0.044711f
C50 VDD1.t1 B 0.044711f
C51 VDD1.n2 B 0.342561f
C52 VDD1.n3 B 1.03557f
C53 VTAIL.t0 B 0.054314f
C54 VTAIL.t3 B 0.054314f
C55 VTAIL.n0 B 0.373768f
C56 VTAIL.n1 B 0.246616f
C57 VTAIL.t7 B 0.47986f
C58 VTAIL.n2 B 0.330987f
C59 VTAIL.t9 B 0.054314f
C60 VTAIL.t6 B 0.054314f
C61 VTAIL.n3 B 0.373768f
C62 VTAIL.n4 B 0.812471f
C63 VTAIL.t4 B 0.054314f
C64 VTAIL.t2 B 0.054314f
C65 VTAIL.n5 B 0.37377f
C66 VTAIL.n6 B 0.812469f
C67 VTAIL.t1 B 0.479863f
C68 VTAIL.n7 B 0.330984f
C69 VTAIL.t10 B 0.054314f
C70 VTAIL.t11 B 0.054314f
C71 VTAIL.n8 B 0.37377f
C72 VTAIL.n9 B 0.288949f
C73 VTAIL.t8 B 0.47986f
C74 VTAIL.n10 B 0.793081f
C75 VTAIL.t5 B 0.47986f
C76 VTAIL.n11 B 0.773989f
C77 VP.n0 B 0.024884f
C78 VP.n1 B 0.005647f
C79 VP.n2 B 0.106676f
C80 VP.t4 B 0.199268f
C81 VP.t3 B 0.199268f
C82 VP.t0 B 0.213289f
C83 VP.n3 B 0.097686f
C84 VP.n4 B 0.110905f
C85 VP.n5 B 0.005647f
C86 VP.n6 B 0.108216f
C87 VP.n7 B 0.746311f
C88 VP.t5 B 0.199268f
C89 VP.n8 B 0.108216f
C90 VP.n9 B 0.771782f
C91 VP.n10 B 0.024884f
C92 VP.n11 B 0.024884f
C93 VP.t1 B 0.199268f
C94 VP.n12 B 0.108216f
C95 VP.n13 B 0.005647f
C96 VP.t2 B 0.199268f
C97 VP.n14 B 0.108216f
C98 VP.n15 B 0.019284f
.ends

