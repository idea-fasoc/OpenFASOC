* NGSPICE file created from diff_pair_sample_0441.ext - technology: sky130A

.subckt diff_pair_sample_0441 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=4.5591 ps=24.16 w=11.69 l=1.98
X1 VTAIL.t14 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X2 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=0 ps=0 w=11.69 l=1.98
X3 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=1.92885 ps=12.02 w=11.69 l=1.98
X4 VDD2.t6 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X5 VDD1.t5 VP.t2 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X6 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=0 ps=0 w=11.69 l=1.98
X7 VTAIL.t8 VP.t3 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=1.92885 ps=12.02 w=11.69 l=1.98
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=0 ps=0 w=11.69 l=1.98
X9 VDD1.t3 VP.t4 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X10 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=1.92885 ps=12.02 w=11.69 l=1.98
X11 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X12 VDD2.t3 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=4.5591 ps=24.16 w=11.69 l=1.98
X13 VTAIL.t7 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=1.92885 ps=12.02 w=11.69 l=1.98
X14 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=4.5591 ps=24.16 w=11.69 l=1.98
X15 VTAIL.t4 VN.t6 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X16 VDD1.t1 VP.t6 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=4.5591 ps=24.16 w=11.69 l=1.98
X17 VTAIL.t10 VP.t7 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X18 VDD2.t0 VN.t7 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.92885 pd=12.02 as=1.92885 ps=12.02 w=11.69 l=1.98
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.5591 pd=24.16 as=0 ps=0 w=11.69 l=1.98
R0 VP.n12 VP.t5 173.139
R1 VP.n14 VP.n11 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n10 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n9 161.3
R6 VP.n23 VP.n22 161.3
R7 VP.n24 VP.n8 161.3
R8 VP.n26 VP.n25 161.3
R9 VP.n27 VP.n7 161.3
R10 VP.n52 VP.n0 161.3
R11 VP.n51 VP.n50 161.3
R12 VP.n49 VP.n1 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n45 VP.n2 161.3
R15 VP.n44 VP.n43 161.3
R16 VP.n42 VP.n3 161.3
R17 VP.n41 VP.n40 161.3
R18 VP.n39 VP.n4 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n5 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n6 161.3
R23 VP.n31 VP.t3 142.287
R24 VP.n38 VP.t4 142.287
R25 VP.n46 VP.t7 142.287
R26 VP.n53 VP.t0 142.287
R27 VP.n28 VP.t6 142.287
R28 VP.n21 VP.t1 142.287
R29 VP.n13 VP.t2 142.287
R30 VP.n31 VP.n30 88.0021
R31 VP.n54 VP.n53 88.0021
R32 VP.n29 VP.n28 88.0021
R33 VP.n13 VP.n12 62.6111
R34 VP.n33 VP.n5 56.5193
R35 VP.n51 VP.n1 56.5193
R36 VP.n26 VP.n8 56.5193
R37 VP.n30 VP.n29 47.8253
R38 VP.n40 VP.n3 40.4934
R39 VP.n44 VP.n3 40.4934
R40 VP.n19 VP.n10 40.4934
R41 VP.n15 VP.n10 40.4934
R42 VP.n33 VP.n32 24.4675
R43 VP.n37 VP.n5 24.4675
R44 VP.n40 VP.n39 24.4675
R45 VP.n45 VP.n44 24.4675
R46 VP.n47 VP.n1 24.4675
R47 VP.n52 VP.n51 24.4675
R48 VP.n27 VP.n26 24.4675
R49 VP.n20 VP.n19 24.4675
R50 VP.n22 VP.n8 24.4675
R51 VP.n15 VP.n14 24.4675
R52 VP.n32 VP.n31 22.7548
R53 VP.n53 VP.n52 22.7548
R54 VP.n28 VP.n27 22.7548
R55 VP.n38 VP.n37 16.8827
R56 VP.n47 VP.n46 16.8827
R57 VP.n22 VP.n21 16.8827
R58 VP.n12 VP.n11 12.915
R59 VP.n39 VP.n38 7.58527
R60 VP.n46 VP.n45 7.58527
R61 VP.n21 VP.n20 7.58527
R62 VP.n14 VP.n13 7.58527
R63 VP.n29 VP.n7 0.278367
R64 VP.n30 VP.n6 0.278367
R65 VP.n54 VP.n0 0.278367
R66 VP.n16 VP.n11 0.189894
R67 VP.n17 VP.n16 0.189894
R68 VP.n18 VP.n17 0.189894
R69 VP.n18 VP.n9 0.189894
R70 VP.n23 VP.n9 0.189894
R71 VP.n24 VP.n23 0.189894
R72 VP.n25 VP.n24 0.189894
R73 VP.n25 VP.n7 0.189894
R74 VP.n34 VP.n6 0.189894
R75 VP.n35 VP.n34 0.189894
R76 VP.n36 VP.n35 0.189894
R77 VP.n36 VP.n4 0.189894
R78 VP.n41 VP.n4 0.189894
R79 VP.n42 VP.n41 0.189894
R80 VP.n43 VP.n42 0.189894
R81 VP.n43 VP.n2 0.189894
R82 VP.n48 VP.n2 0.189894
R83 VP.n49 VP.n48 0.189894
R84 VP.n50 VP.n49 0.189894
R85 VP.n50 VP.n0 0.189894
R86 VP VP.n54 0.153454
R87 VTAIL.n11 VTAIL.t7 45.6374
R88 VTAIL.n10 VTAIL.t5 45.6374
R89 VTAIL.n7 VTAIL.t1 45.6374
R90 VTAIL.n15 VTAIL.t2 45.6372
R91 VTAIL.n2 VTAIL.t0 45.6372
R92 VTAIL.n3 VTAIL.t12 45.6372
R93 VTAIL.n6 VTAIL.t8 45.6372
R94 VTAIL.n14 VTAIL.t9 45.6372
R95 VTAIL.n13 VTAIL.n12 43.9437
R96 VTAIL.n9 VTAIL.n8 43.9437
R97 VTAIL.n1 VTAIL.n0 43.9434
R98 VTAIL.n5 VTAIL.n4 43.9434
R99 VTAIL.n15 VTAIL.n14 24.4358
R100 VTAIL.n7 VTAIL.n6 24.4358
R101 VTAIL.n9 VTAIL.n7 1.99188
R102 VTAIL.n10 VTAIL.n9 1.99188
R103 VTAIL.n13 VTAIL.n11 1.99188
R104 VTAIL.n14 VTAIL.n13 1.99188
R105 VTAIL.n6 VTAIL.n5 1.99188
R106 VTAIL.n5 VTAIL.n3 1.99188
R107 VTAIL.n2 VTAIL.n1 1.99188
R108 VTAIL VTAIL.n15 1.93369
R109 VTAIL.n0 VTAIL.t15 1.69426
R110 VTAIL.n0 VTAIL.t4 1.69426
R111 VTAIL.n4 VTAIL.t11 1.69426
R112 VTAIL.n4 VTAIL.t10 1.69426
R113 VTAIL.n12 VTAIL.t13 1.69426
R114 VTAIL.n12 VTAIL.t14 1.69426
R115 VTAIL.n8 VTAIL.t3 1.69426
R116 VTAIL.n8 VTAIL.t6 1.69426
R117 VTAIL.n11 VTAIL.n10 0.470328
R118 VTAIL.n3 VTAIL.n2 0.470328
R119 VTAIL VTAIL.n1 0.0586897
R120 VDD1 VDD1.n0 61.6763
R121 VDD1.n3 VDD1.n2 61.5626
R122 VDD1.n3 VDD1.n1 61.5626
R123 VDD1.n5 VDD1.n4 60.6223
R124 VDD1.n5 VDD1.n3 43.3371
R125 VDD1.n4 VDD1.t6 1.69426
R126 VDD1.n4 VDD1.t1 1.69426
R127 VDD1.n0 VDD1.t2 1.69426
R128 VDD1.n0 VDD1.t5 1.69426
R129 VDD1.n2 VDD1.t0 1.69426
R130 VDD1.n2 VDD1.t7 1.69426
R131 VDD1.n1 VDD1.t4 1.69426
R132 VDD1.n1 VDD1.t3 1.69426
R133 VDD1 VDD1.n5 0.938
R134 B.n623 B.n129 585
R135 B.n129 B.n78 585
R136 B.n625 B.n624 585
R137 B.n627 B.n128 585
R138 B.n630 B.n629 585
R139 B.n631 B.n127 585
R140 B.n633 B.n632 585
R141 B.n635 B.n126 585
R142 B.n638 B.n637 585
R143 B.n639 B.n125 585
R144 B.n641 B.n640 585
R145 B.n643 B.n124 585
R146 B.n646 B.n645 585
R147 B.n647 B.n123 585
R148 B.n649 B.n648 585
R149 B.n651 B.n122 585
R150 B.n654 B.n653 585
R151 B.n655 B.n121 585
R152 B.n657 B.n656 585
R153 B.n659 B.n120 585
R154 B.n662 B.n661 585
R155 B.n663 B.n119 585
R156 B.n665 B.n664 585
R157 B.n667 B.n118 585
R158 B.n670 B.n669 585
R159 B.n671 B.n117 585
R160 B.n673 B.n672 585
R161 B.n675 B.n116 585
R162 B.n678 B.n677 585
R163 B.n679 B.n115 585
R164 B.n681 B.n680 585
R165 B.n683 B.n114 585
R166 B.n686 B.n685 585
R167 B.n687 B.n113 585
R168 B.n689 B.n688 585
R169 B.n691 B.n112 585
R170 B.n694 B.n693 585
R171 B.n695 B.n111 585
R172 B.n697 B.n696 585
R173 B.n699 B.n110 585
R174 B.n701 B.n700 585
R175 B.n703 B.n702 585
R176 B.n706 B.n705 585
R177 B.n707 B.n105 585
R178 B.n709 B.n708 585
R179 B.n711 B.n104 585
R180 B.n714 B.n713 585
R181 B.n715 B.n103 585
R182 B.n717 B.n716 585
R183 B.n719 B.n102 585
R184 B.n722 B.n721 585
R185 B.n724 B.n99 585
R186 B.n726 B.n725 585
R187 B.n728 B.n98 585
R188 B.n731 B.n730 585
R189 B.n732 B.n97 585
R190 B.n734 B.n733 585
R191 B.n736 B.n96 585
R192 B.n739 B.n738 585
R193 B.n740 B.n95 585
R194 B.n742 B.n741 585
R195 B.n744 B.n94 585
R196 B.n747 B.n746 585
R197 B.n748 B.n93 585
R198 B.n750 B.n749 585
R199 B.n752 B.n92 585
R200 B.n755 B.n754 585
R201 B.n756 B.n91 585
R202 B.n758 B.n757 585
R203 B.n760 B.n90 585
R204 B.n763 B.n762 585
R205 B.n764 B.n89 585
R206 B.n766 B.n765 585
R207 B.n768 B.n88 585
R208 B.n771 B.n770 585
R209 B.n772 B.n87 585
R210 B.n774 B.n773 585
R211 B.n776 B.n86 585
R212 B.n779 B.n778 585
R213 B.n780 B.n85 585
R214 B.n782 B.n781 585
R215 B.n784 B.n84 585
R216 B.n787 B.n786 585
R217 B.n788 B.n83 585
R218 B.n790 B.n789 585
R219 B.n792 B.n82 585
R220 B.n795 B.n794 585
R221 B.n796 B.n81 585
R222 B.n798 B.n797 585
R223 B.n800 B.n80 585
R224 B.n803 B.n802 585
R225 B.n804 B.n79 585
R226 B.n622 B.n77 585
R227 B.n807 B.n77 585
R228 B.n621 B.n76 585
R229 B.n808 B.n76 585
R230 B.n620 B.n75 585
R231 B.n809 B.n75 585
R232 B.n619 B.n618 585
R233 B.n618 B.n71 585
R234 B.n617 B.n70 585
R235 B.n815 B.n70 585
R236 B.n616 B.n69 585
R237 B.n816 B.n69 585
R238 B.n615 B.n68 585
R239 B.n817 B.n68 585
R240 B.n614 B.n613 585
R241 B.n613 B.n64 585
R242 B.n612 B.n63 585
R243 B.n823 B.n63 585
R244 B.n611 B.n62 585
R245 B.n824 B.n62 585
R246 B.n610 B.n61 585
R247 B.n825 B.n61 585
R248 B.n609 B.n608 585
R249 B.n608 B.n57 585
R250 B.n607 B.n56 585
R251 B.n831 B.n56 585
R252 B.n606 B.n55 585
R253 B.n832 B.n55 585
R254 B.n605 B.n54 585
R255 B.n833 B.n54 585
R256 B.n604 B.n603 585
R257 B.n603 B.n50 585
R258 B.n602 B.n49 585
R259 B.n839 B.n49 585
R260 B.n601 B.n48 585
R261 B.n840 B.n48 585
R262 B.n600 B.n47 585
R263 B.n841 B.n47 585
R264 B.n599 B.n598 585
R265 B.n598 B.n43 585
R266 B.n597 B.n42 585
R267 B.n847 B.n42 585
R268 B.n596 B.n41 585
R269 B.n848 B.n41 585
R270 B.n595 B.n40 585
R271 B.n849 B.n40 585
R272 B.n594 B.n593 585
R273 B.n593 B.n39 585
R274 B.n592 B.n35 585
R275 B.n855 B.n35 585
R276 B.n591 B.n34 585
R277 B.n856 B.n34 585
R278 B.n590 B.n33 585
R279 B.n857 B.n33 585
R280 B.n589 B.n588 585
R281 B.n588 B.n29 585
R282 B.n587 B.n28 585
R283 B.n863 B.n28 585
R284 B.n586 B.n27 585
R285 B.n864 B.n27 585
R286 B.n585 B.n26 585
R287 B.n865 B.n26 585
R288 B.n584 B.n583 585
R289 B.n583 B.n22 585
R290 B.n582 B.n21 585
R291 B.n871 B.n21 585
R292 B.n581 B.n20 585
R293 B.n872 B.n20 585
R294 B.n580 B.n19 585
R295 B.n873 B.n19 585
R296 B.n579 B.n578 585
R297 B.n578 B.n15 585
R298 B.n577 B.n14 585
R299 B.n879 B.n14 585
R300 B.n576 B.n13 585
R301 B.t0 B.n13 585
R302 B.n575 B.n12 585
R303 B.n880 B.n12 585
R304 B.n574 B.n573 585
R305 B.n573 B.n8 585
R306 B.n572 B.n7 585
R307 B.n886 B.n7 585
R308 B.n571 B.n6 585
R309 B.n887 B.n6 585
R310 B.n570 B.n5 585
R311 B.n888 B.n5 585
R312 B.n569 B.n568 585
R313 B.n568 B.n4 585
R314 B.n567 B.n130 585
R315 B.n567 B.n566 585
R316 B.n557 B.n131 585
R317 B.n132 B.n131 585
R318 B.n559 B.n558 585
R319 B.n560 B.n559 585
R320 B.n556 B.n136 585
R321 B.n136 B.t5 585
R322 B.n555 B.n554 585
R323 B.n554 B.n553 585
R324 B.n138 B.n137 585
R325 B.n139 B.n138 585
R326 B.n546 B.n545 585
R327 B.n547 B.n546 585
R328 B.n544 B.n144 585
R329 B.n144 B.n143 585
R330 B.n543 B.n542 585
R331 B.n542 B.n541 585
R332 B.n146 B.n145 585
R333 B.n147 B.n146 585
R334 B.n534 B.n533 585
R335 B.n535 B.n534 585
R336 B.n532 B.n152 585
R337 B.n152 B.n151 585
R338 B.n531 B.n530 585
R339 B.n530 B.n529 585
R340 B.n154 B.n153 585
R341 B.n155 B.n154 585
R342 B.n522 B.n521 585
R343 B.n523 B.n522 585
R344 B.n520 B.n160 585
R345 B.n160 B.n159 585
R346 B.n519 B.n518 585
R347 B.n518 B.n517 585
R348 B.n162 B.n161 585
R349 B.n510 B.n162 585
R350 B.n509 B.n508 585
R351 B.n511 B.n509 585
R352 B.n507 B.n167 585
R353 B.n167 B.n166 585
R354 B.n506 B.n505 585
R355 B.n505 B.n504 585
R356 B.n169 B.n168 585
R357 B.n170 B.n169 585
R358 B.n497 B.n496 585
R359 B.n498 B.n497 585
R360 B.n495 B.n175 585
R361 B.n175 B.n174 585
R362 B.n494 B.n493 585
R363 B.n493 B.n492 585
R364 B.n177 B.n176 585
R365 B.n178 B.n177 585
R366 B.n485 B.n484 585
R367 B.n486 B.n485 585
R368 B.n483 B.n183 585
R369 B.n183 B.n182 585
R370 B.n482 B.n481 585
R371 B.n481 B.n480 585
R372 B.n185 B.n184 585
R373 B.n186 B.n185 585
R374 B.n473 B.n472 585
R375 B.n474 B.n473 585
R376 B.n471 B.n191 585
R377 B.n191 B.n190 585
R378 B.n470 B.n469 585
R379 B.n469 B.n468 585
R380 B.n193 B.n192 585
R381 B.n194 B.n193 585
R382 B.n461 B.n460 585
R383 B.n462 B.n461 585
R384 B.n459 B.n199 585
R385 B.n199 B.n198 585
R386 B.n458 B.n457 585
R387 B.n457 B.n456 585
R388 B.n201 B.n200 585
R389 B.n202 B.n201 585
R390 B.n449 B.n448 585
R391 B.n450 B.n449 585
R392 B.n447 B.n207 585
R393 B.n207 B.n206 585
R394 B.n446 B.n445 585
R395 B.n445 B.n444 585
R396 B.n441 B.n211 585
R397 B.n440 B.n439 585
R398 B.n437 B.n212 585
R399 B.n437 B.n210 585
R400 B.n436 B.n435 585
R401 B.n434 B.n433 585
R402 B.n432 B.n214 585
R403 B.n430 B.n429 585
R404 B.n428 B.n215 585
R405 B.n427 B.n426 585
R406 B.n424 B.n216 585
R407 B.n422 B.n421 585
R408 B.n420 B.n217 585
R409 B.n419 B.n418 585
R410 B.n416 B.n218 585
R411 B.n414 B.n413 585
R412 B.n412 B.n219 585
R413 B.n411 B.n410 585
R414 B.n408 B.n220 585
R415 B.n406 B.n405 585
R416 B.n404 B.n221 585
R417 B.n403 B.n402 585
R418 B.n400 B.n222 585
R419 B.n398 B.n397 585
R420 B.n396 B.n223 585
R421 B.n395 B.n394 585
R422 B.n392 B.n224 585
R423 B.n390 B.n389 585
R424 B.n388 B.n225 585
R425 B.n387 B.n386 585
R426 B.n384 B.n226 585
R427 B.n382 B.n381 585
R428 B.n380 B.n227 585
R429 B.n379 B.n378 585
R430 B.n376 B.n228 585
R431 B.n374 B.n373 585
R432 B.n372 B.n229 585
R433 B.n371 B.n370 585
R434 B.n368 B.n230 585
R435 B.n366 B.n365 585
R436 B.n364 B.n231 585
R437 B.n363 B.n362 585
R438 B.n360 B.n359 585
R439 B.n358 B.n357 585
R440 B.n356 B.n236 585
R441 B.n354 B.n353 585
R442 B.n352 B.n237 585
R443 B.n351 B.n350 585
R444 B.n348 B.n238 585
R445 B.n346 B.n345 585
R446 B.n344 B.n239 585
R447 B.n342 B.n341 585
R448 B.n339 B.n242 585
R449 B.n337 B.n336 585
R450 B.n335 B.n243 585
R451 B.n334 B.n333 585
R452 B.n331 B.n244 585
R453 B.n329 B.n328 585
R454 B.n327 B.n245 585
R455 B.n326 B.n325 585
R456 B.n323 B.n246 585
R457 B.n321 B.n320 585
R458 B.n319 B.n247 585
R459 B.n318 B.n317 585
R460 B.n315 B.n248 585
R461 B.n313 B.n312 585
R462 B.n311 B.n249 585
R463 B.n310 B.n309 585
R464 B.n307 B.n250 585
R465 B.n305 B.n304 585
R466 B.n303 B.n251 585
R467 B.n302 B.n301 585
R468 B.n299 B.n252 585
R469 B.n297 B.n296 585
R470 B.n295 B.n253 585
R471 B.n294 B.n293 585
R472 B.n291 B.n254 585
R473 B.n289 B.n288 585
R474 B.n287 B.n255 585
R475 B.n286 B.n285 585
R476 B.n283 B.n256 585
R477 B.n281 B.n280 585
R478 B.n279 B.n257 585
R479 B.n278 B.n277 585
R480 B.n275 B.n258 585
R481 B.n273 B.n272 585
R482 B.n271 B.n259 585
R483 B.n270 B.n269 585
R484 B.n267 B.n260 585
R485 B.n265 B.n264 585
R486 B.n263 B.n262 585
R487 B.n209 B.n208 585
R488 B.n443 B.n442 585
R489 B.n444 B.n443 585
R490 B.n205 B.n204 585
R491 B.n206 B.n205 585
R492 B.n452 B.n451 585
R493 B.n451 B.n450 585
R494 B.n453 B.n203 585
R495 B.n203 B.n202 585
R496 B.n455 B.n454 585
R497 B.n456 B.n455 585
R498 B.n197 B.n196 585
R499 B.n198 B.n197 585
R500 B.n464 B.n463 585
R501 B.n463 B.n462 585
R502 B.n465 B.n195 585
R503 B.n195 B.n194 585
R504 B.n467 B.n466 585
R505 B.n468 B.n467 585
R506 B.n189 B.n188 585
R507 B.n190 B.n189 585
R508 B.n476 B.n475 585
R509 B.n475 B.n474 585
R510 B.n477 B.n187 585
R511 B.n187 B.n186 585
R512 B.n479 B.n478 585
R513 B.n480 B.n479 585
R514 B.n181 B.n180 585
R515 B.n182 B.n181 585
R516 B.n488 B.n487 585
R517 B.n487 B.n486 585
R518 B.n489 B.n179 585
R519 B.n179 B.n178 585
R520 B.n491 B.n490 585
R521 B.n492 B.n491 585
R522 B.n173 B.n172 585
R523 B.n174 B.n173 585
R524 B.n500 B.n499 585
R525 B.n499 B.n498 585
R526 B.n501 B.n171 585
R527 B.n171 B.n170 585
R528 B.n503 B.n502 585
R529 B.n504 B.n503 585
R530 B.n165 B.n164 585
R531 B.n166 B.n165 585
R532 B.n513 B.n512 585
R533 B.n512 B.n511 585
R534 B.n514 B.n163 585
R535 B.n510 B.n163 585
R536 B.n516 B.n515 585
R537 B.n517 B.n516 585
R538 B.n158 B.n157 585
R539 B.n159 B.n158 585
R540 B.n525 B.n524 585
R541 B.n524 B.n523 585
R542 B.n526 B.n156 585
R543 B.n156 B.n155 585
R544 B.n528 B.n527 585
R545 B.n529 B.n528 585
R546 B.n150 B.n149 585
R547 B.n151 B.n150 585
R548 B.n537 B.n536 585
R549 B.n536 B.n535 585
R550 B.n538 B.n148 585
R551 B.n148 B.n147 585
R552 B.n540 B.n539 585
R553 B.n541 B.n540 585
R554 B.n142 B.n141 585
R555 B.n143 B.n142 585
R556 B.n549 B.n548 585
R557 B.n548 B.n547 585
R558 B.n550 B.n140 585
R559 B.n140 B.n139 585
R560 B.n552 B.n551 585
R561 B.n553 B.n552 585
R562 B.n135 B.n134 585
R563 B.t5 B.n135 585
R564 B.n562 B.n561 585
R565 B.n561 B.n560 585
R566 B.n563 B.n133 585
R567 B.n133 B.n132 585
R568 B.n565 B.n564 585
R569 B.n566 B.n565 585
R570 B.n2 B.n0 585
R571 B.n4 B.n2 585
R572 B.n3 B.n1 585
R573 B.n887 B.n3 585
R574 B.n885 B.n884 585
R575 B.n886 B.n885 585
R576 B.n883 B.n9 585
R577 B.n9 B.n8 585
R578 B.n882 B.n881 585
R579 B.n881 B.n880 585
R580 B.n11 B.n10 585
R581 B.t0 B.n11 585
R582 B.n878 B.n877 585
R583 B.n879 B.n878 585
R584 B.n876 B.n16 585
R585 B.n16 B.n15 585
R586 B.n875 B.n874 585
R587 B.n874 B.n873 585
R588 B.n18 B.n17 585
R589 B.n872 B.n18 585
R590 B.n870 B.n869 585
R591 B.n871 B.n870 585
R592 B.n868 B.n23 585
R593 B.n23 B.n22 585
R594 B.n867 B.n866 585
R595 B.n866 B.n865 585
R596 B.n25 B.n24 585
R597 B.n864 B.n25 585
R598 B.n862 B.n861 585
R599 B.n863 B.n862 585
R600 B.n860 B.n30 585
R601 B.n30 B.n29 585
R602 B.n859 B.n858 585
R603 B.n858 B.n857 585
R604 B.n32 B.n31 585
R605 B.n856 B.n32 585
R606 B.n854 B.n853 585
R607 B.n855 B.n854 585
R608 B.n852 B.n36 585
R609 B.n39 B.n36 585
R610 B.n851 B.n850 585
R611 B.n850 B.n849 585
R612 B.n38 B.n37 585
R613 B.n848 B.n38 585
R614 B.n846 B.n845 585
R615 B.n847 B.n846 585
R616 B.n844 B.n44 585
R617 B.n44 B.n43 585
R618 B.n843 B.n842 585
R619 B.n842 B.n841 585
R620 B.n46 B.n45 585
R621 B.n840 B.n46 585
R622 B.n838 B.n837 585
R623 B.n839 B.n838 585
R624 B.n836 B.n51 585
R625 B.n51 B.n50 585
R626 B.n835 B.n834 585
R627 B.n834 B.n833 585
R628 B.n53 B.n52 585
R629 B.n832 B.n53 585
R630 B.n830 B.n829 585
R631 B.n831 B.n830 585
R632 B.n828 B.n58 585
R633 B.n58 B.n57 585
R634 B.n827 B.n826 585
R635 B.n826 B.n825 585
R636 B.n60 B.n59 585
R637 B.n824 B.n60 585
R638 B.n822 B.n821 585
R639 B.n823 B.n822 585
R640 B.n820 B.n65 585
R641 B.n65 B.n64 585
R642 B.n819 B.n818 585
R643 B.n818 B.n817 585
R644 B.n67 B.n66 585
R645 B.n816 B.n67 585
R646 B.n814 B.n813 585
R647 B.n815 B.n814 585
R648 B.n812 B.n72 585
R649 B.n72 B.n71 585
R650 B.n811 B.n810 585
R651 B.n810 B.n809 585
R652 B.n74 B.n73 585
R653 B.n808 B.n74 585
R654 B.n806 B.n805 585
R655 B.n807 B.n806 585
R656 B.n890 B.n889 585
R657 B.n889 B.n888 585
R658 B.n443 B.n211 511.721
R659 B.n806 B.n79 511.721
R660 B.n445 B.n209 511.721
R661 B.n129 B.n77 511.721
R662 B.n240 B.t8 349.158
R663 B.n232 B.t16 349.158
R664 B.n100 B.t19 349.158
R665 B.n106 B.t12 349.158
R666 B.n626 B.n78 256.663
R667 B.n628 B.n78 256.663
R668 B.n634 B.n78 256.663
R669 B.n636 B.n78 256.663
R670 B.n642 B.n78 256.663
R671 B.n644 B.n78 256.663
R672 B.n650 B.n78 256.663
R673 B.n652 B.n78 256.663
R674 B.n658 B.n78 256.663
R675 B.n660 B.n78 256.663
R676 B.n666 B.n78 256.663
R677 B.n668 B.n78 256.663
R678 B.n674 B.n78 256.663
R679 B.n676 B.n78 256.663
R680 B.n682 B.n78 256.663
R681 B.n684 B.n78 256.663
R682 B.n690 B.n78 256.663
R683 B.n692 B.n78 256.663
R684 B.n698 B.n78 256.663
R685 B.n109 B.n78 256.663
R686 B.n704 B.n78 256.663
R687 B.n710 B.n78 256.663
R688 B.n712 B.n78 256.663
R689 B.n718 B.n78 256.663
R690 B.n720 B.n78 256.663
R691 B.n727 B.n78 256.663
R692 B.n729 B.n78 256.663
R693 B.n735 B.n78 256.663
R694 B.n737 B.n78 256.663
R695 B.n743 B.n78 256.663
R696 B.n745 B.n78 256.663
R697 B.n751 B.n78 256.663
R698 B.n753 B.n78 256.663
R699 B.n759 B.n78 256.663
R700 B.n761 B.n78 256.663
R701 B.n767 B.n78 256.663
R702 B.n769 B.n78 256.663
R703 B.n775 B.n78 256.663
R704 B.n777 B.n78 256.663
R705 B.n783 B.n78 256.663
R706 B.n785 B.n78 256.663
R707 B.n791 B.n78 256.663
R708 B.n793 B.n78 256.663
R709 B.n799 B.n78 256.663
R710 B.n801 B.n78 256.663
R711 B.n438 B.n210 256.663
R712 B.n213 B.n210 256.663
R713 B.n431 B.n210 256.663
R714 B.n425 B.n210 256.663
R715 B.n423 B.n210 256.663
R716 B.n417 B.n210 256.663
R717 B.n415 B.n210 256.663
R718 B.n409 B.n210 256.663
R719 B.n407 B.n210 256.663
R720 B.n401 B.n210 256.663
R721 B.n399 B.n210 256.663
R722 B.n393 B.n210 256.663
R723 B.n391 B.n210 256.663
R724 B.n385 B.n210 256.663
R725 B.n383 B.n210 256.663
R726 B.n377 B.n210 256.663
R727 B.n375 B.n210 256.663
R728 B.n369 B.n210 256.663
R729 B.n367 B.n210 256.663
R730 B.n361 B.n210 256.663
R731 B.n235 B.n210 256.663
R732 B.n355 B.n210 256.663
R733 B.n349 B.n210 256.663
R734 B.n347 B.n210 256.663
R735 B.n340 B.n210 256.663
R736 B.n338 B.n210 256.663
R737 B.n332 B.n210 256.663
R738 B.n330 B.n210 256.663
R739 B.n324 B.n210 256.663
R740 B.n322 B.n210 256.663
R741 B.n316 B.n210 256.663
R742 B.n314 B.n210 256.663
R743 B.n308 B.n210 256.663
R744 B.n306 B.n210 256.663
R745 B.n300 B.n210 256.663
R746 B.n298 B.n210 256.663
R747 B.n292 B.n210 256.663
R748 B.n290 B.n210 256.663
R749 B.n284 B.n210 256.663
R750 B.n282 B.n210 256.663
R751 B.n276 B.n210 256.663
R752 B.n274 B.n210 256.663
R753 B.n268 B.n210 256.663
R754 B.n266 B.n210 256.663
R755 B.n261 B.n210 256.663
R756 B.n443 B.n205 163.367
R757 B.n451 B.n205 163.367
R758 B.n451 B.n203 163.367
R759 B.n455 B.n203 163.367
R760 B.n455 B.n197 163.367
R761 B.n463 B.n197 163.367
R762 B.n463 B.n195 163.367
R763 B.n467 B.n195 163.367
R764 B.n467 B.n189 163.367
R765 B.n475 B.n189 163.367
R766 B.n475 B.n187 163.367
R767 B.n479 B.n187 163.367
R768 B.n479 B.n181 163.367
R769 B.n487 B.n181 163.367
R770 B.n487 B.n179 163.367
R771 B.n491 B.n179 163.367
R772 B.n491 B.n173 163.367
R773 B.n499 B.n173 163.367
R774 B.n499 B.n171 163.367
R775 B.n503 B.n171 163.367
R776 B.n503 B.n165 163.367
R777 B.n512 B.n165 163.367
R778 B.n512 B.n163 163.367
R779 B.n516 B.n163 163.367
R780 B.n516 B.n158 163.367
R781 B.n524 B.n158 163.367
R782 B.n524 B.n156 163.367
R783 B.n528 B.n156 163.367
R784 B.n528 B.n150 163.367
R785 B.n536 B.n150 163.367
R786 B.n536 B.n148 163.367
R787 B.n540 B.n148 163.367
R788 B.n540 B.n142 163.367
R789 B.n548 B.n142 163.367
R790 B.n548 B.n140 163.367
R791 B.n552 B.n140 163.367
R792 B.n552 B.n135 163.367
R793 B.n561 B.n135 163.367
R794 B.n561 B.n133 163.367
R795 B.n565 B.n133 163.367
R796 B.n565 B.n2 163.367
R797 B.n889 B.n2 163.367
R798 B.n889 B.n3 163.367
R799 B.n885 B.n3 163.367
R800 B.n885 B.n9 163.367
R801 B.n881 B.n9 163.367
R802 B.n881 B.n11 163.367
R803 B.n878 B.n11 163.367
R804 B.n878 B.n16 163.367
R805 B.n874 B.n16 163.367
R806 B.n874 B.n18 163.367
R807 B.n870 B.n18 163.367
R808 B.n870 B.n23 163.367
R809 B.n866 B.n23 163.367
R810 B.n866 B.n25 163.367
R811 B.n862 B.n25 163.367
R812 B.n862 B.n30 163.367
R813 B.n858 B.n30 163.367
R814 B.n858 B.n32 163.367
R815 B.n854 B.n32 163.367
R816 B.n854 B.n36 163.367
R817 B.n850 B.n36 163.367
R818 B.n850 B.n38 163.367
R819 B.n846 B.n38 163.367
R820 B.n846 B.n44 163.367
R821 B.n842 B.n44 163.367
R822 B.n842 B.n46 163.367
R823 B.n838 B.n46 163.367
R824 B.n838 B.n51 163.367
R825 B.n834 B.n51 163.367
R826 B.n834 B.n53 163.367
R827 B.n830 B.n53 163.367
R828 B.n830 B.n58 163.367
R829 B.n826 B.n58 163.367
R830 B.n826 B.n60 163.367
R831 B.n822 B.n60 163.367
R832 B.n822 B.n65 163.367
R833 B.n818 B.n65 163.367
R834 B.n818 B.n67 163.367
R835 B.n814 B.n67 163.367
R836 B.n814 B.n72 163.367
R837 B.n810 B.n72 163.367
R838 B.n810 B.n74 163.367
R839 B.n806 B.n74 163.367
R840 B.n439 B.n437 163.367
R841 B.n437 B.n436 163.367
R842 B.n433 B.n432 163.367
R843 B.n430 B.n215 163.367
R844 B.n426 B.n424 163.367
R845 B.n422 B.n217 163.367
R846 B.n418 B.n416 163.367
R847 B.n414 B.n219 163.367
R848 B.n410 B.n408 163.367
R849 B.n406 B.n221 163.367
R850 B.n402 B.n400 163.367
R851 B.n398 B.n223 163.367
R852 B.n394 B.n392 163.367
R853 B.n390 B.n225 163.367
R854 B.n386 B.n384 163.367
R855 B.n382 B.n227 163.367
R856 B.n378 B.n376 163.367
R857 B.n374 B.n229 163.367
R858 B.n370 B.n368 163.367
R859 B.n366 B.n231 163.367
R860 B.n362 B.n360 163.367
R861 B.n357 B.n356 163.367
R862 B.n354 B.n237 163.367
R863 B.n350 B.n348 163.367
R864 B.n346 B.n239 163.367
R865 B.n341 B.n339 163.367
R866 B.n337 B.n243 163.367
R867 B.n333 B.n331 163.367
R868 B.n329 B.n245 163.367
R869 B.n325 B.n323 163.367
R870 B.n321 B.n247 163.367
R871 B.n317 B.n315 163.367
R872 B.n313 B.n249 163.367
R873 B.n309 B.n307 163.367
R874 B.n305 B.n251 163.367
R875 B.n301 B.n299 163.367
R876 B.n297 B.n253 163.367
R877 B.n293 B.n291 163.367
R878 B.n289 B.n255 163.367
R879 B.n285 B.n283 163.367
R880 B.n281 B.n257 163.367
R881 B.n277 B.n275 163.367
R882 B.n273 B.n259 163.367
R883 B.n269 B.n267 163.367
R884 B.n265 B.n262 163.367
R885 B.n445 B.n207 163.367
R886 B.n449 B.n207 163.367
R887 B.n449 B.n201 163.367
R888 B.n457 B.n201 163.367
R889 B.n457 B.n199 163.367
R890 B.n461 B.n199 163.367
R891 B.n461 B.n193 163.367
R892 B.n469 B.n193 163.367
R893 B.n469 B.n191 163.367
R894 B.n473 B.n191 163.367
R895 B.n473 B.n185 163.367
R896 B.n481 B.n185 163.367
R897 B.n481 B.n183 163.367
R898 B.n485 B.n183 163.367
R899 B.n485 B.n177 163.367
R900 B.n493 B.n177 163.367
R901 B.n493 B.n175 163.367
R902 B.n497 B.n175 163.367
R903 B.n497 B.n169 163.367
R904 B.n505 B.n169 163.367
R905 B.n505 B.n167 163.367
R906 B.n509 B.n167 163.367
R907 B.n509 B.n162 163.367
R908 B.n518 B.n162 163.367
R909 B.n518 B.n160 163.367
R910 B.n522 B.n160 163.367
R911 B.n522 B.n154 163.367
R912 B.n530 B.n154 163.367
R913 B.n530 B.n152 163.367
R914 B.n534 B.n152 163.367
R915 B.n534 B.n146 163.367
R916 B.n542 B.n146 163.367
R917 B.n542 B.n144 163.367
R918 B.n546 B.n144 163.367
R919 B.n546 B.n138 163.367
R920 B.n554 B.n138 163.367
R921 B.n554 B.n136 163.367
R922 B.n559 B.n136 163.367
R923 B.n559 B.n131 163.367
R924 B.n567 B.n131 163.367
R925 B.n568 B.n567 163.367
R926 B.n568 B.n5 163.367
R927 B.n6 B.n5 163.367
R928 B.n7 B.n6 163.367
R929 B.n573 B.n7 163.367
R930 B.n573 B.n12 163.367
R931 B.n13 B.n12 163.367
R932 B.n14 B.n13 163.367
R933 B.n578 B.n14 163.367
R934 B.n578 B.n19 163.367
R935 B.n20 B.n19 163.367
R936 B.n21 B.n20 163.367
R937 B.n583 B.n21 163.367
R938 B.n583 B.n26 163.367
R939 B.n27 B.n26 163.367
R940 B.n28 B.n27 163.367
R941 B.n588 B.n28 163.367
R942 B.n588 B.n33 163.367
R943 B.n34 B.n33 163.367
R944 B.n35 B.n34 163.367
R945 B.n593 B.n35 163.367
R946 B.n593 B.n40 163.367
R947 B.n41 B.n40 163.367
R948 B.n42 B.n41 163.367
R949 B.n598 B.n42 163.367
R950 B.n598 B.n47 163.367
R951 B.n48 B.n47 163.367
R952 B.n49 B.n48 163.367
R953 B.n603 B.n49 163.367
R954 B.n603 B.n54 163.367
R955 B.n55 B.n54 163.367
R956 B.n56 B.n55 163.367
R957 B.n608 B.n56 163.367
R958 B.n608 B.n61 163.367
R959 B.n62 B.n61 163.367
R960 B.n63 B.n62 163.367
R961 B.n613 B.n63 163.367
R962 B.n613 B.n68 163.367
R963 B.n69 B.n68 163.367
R964 B.n70 B.n69 163.367
R965 B.n618 B.n70 163.367
R966 B.n618 B.n75 163.367
R967 B.n76 B.n75 163.367
R968 B.n77 B.n76 163.367
R969 B.n802 B.n800 163.367
R970 B.n798 B.n81 163.367
R971 B.n794 B.n792 163.367
R972 B.n790 B.n83 163.367
R973 B.n786 B.n784 163.367
R974 B.n782 B.n85 163.367
R975 B.n778 B.n776 163.367
R976 B.n774 B.n87 163.367
R977 B.n770 B.n768 163.367
R978 B.n766 B.n89 163.367
R979 B.n762 B.n760 163.367
R980 B.n758 B.n91 163.367
R981 B.n754 B.n752 163.367
R982 B.n750 B.n93 163.367
R983 B.n746 B.n744 163.367
R984 B.n742 B.n95 163.367
R985 B.n738 B.n736 163.367
R986 B.n734 B.n97 163.367
R987 B.n730 B.n728 163.367
R988 B.n726 B.n99 163.367
R989 B.n721 B.n719 163.367
R990 B.n717 B.n103 163.367
R991 B.n713 B.n711 163.367
R992 B.n709 B.n105 163.367
R993 B.n705 B.n703 163.367
R994 B.n700 B.n699 163.367
R995 B.n697 B.n111 163.367
R996 B.n693 B.n691 163.367
R997 B.n689 B.n113 163.367
R998 B.n685 B.n683 163.367
R999 B.n681 B.n115 163.367
R1000 B.n677 B.n675 163.367
R1001 B.n673 B.n117 163.367
R1002 B.n669 B.n667 163.367
R1003 B.n665 B.n119 163.367
R1004 B.n661 B.n659 163.367
R1005 B.n657 B.n121 163.367
R1006 B.n653 B.n651 163.367
R1007 B.n649 B.n123 163.367
R1008 B.n645 B.n643 163.367
R1009 B.n641 B.n125 163.367
R1010 B.n637 B.n635 163.367
R1011 B.n633 B.n127 163.367
R1012 B.n629 B.n627 163.367
R1013 B.n625 B.n129 163.367
R1014 B.n240 B.t11 115.154
R1015 B.n106 B.t14 115.154
R1016 B.n232 B.t18 115.139
R1017 B.n100 B.t20 115.139
R1018 B.n444 B.n210 83.6433
R1019 B.n807 B.n78 83.6433
R1020 B.n438 B.n211 71.676
R1021 B.n436 B.n213 71.676
R1022 B.n432 B.n431 71.676
R1023 B.n425 B.n215 71.676
R1024 B.n424 B.n423 71.676
R1025 B.n417 B.n217 71.676
R1026 B.n416 B.n415 71.676
R1027 B.n409 B.n219 71.676
R1028 B.n408 B.n407 71.676
R1029 B.n401 B.n221 71.676
R1030 B.n400 B.n399 71.676
R1031 B.n393 B.n223 71.676
R1032 B.n392 B.n391 71.676
R1033 B.n385 B.n225 71.676
R1034 B.n384 B.n383 71.676
R1035 B.n377 B.n227 71.676
R1036 B.n376 B.n375 71.676
R1037 B.n369 B.n229 71.676
R1038 B.n368 B.n367 71.676
R1039 B.n361 B.n231 71.676
R1040 B.n360 B.n235 71.676
R1041 B.n356 B.n355 71.676
R1042 B.n349 B.n237 71.676
R1043 B.n348 B.n347 71.676
R1044 B.n340 B.n239 71.676
R1045 B.n339 B.n338 71.676
R1046 B.n332 B.n243 71.676
R1047 B.n331 B.n330 71.676
R1048 B.n324 B.n245 71.676
R1049 B.n323 B.n322 71.676
R1050 B.n316 B.n247 71.676
R1051 B.n315 B.n314 71.676
R1052 B.n308 B.n249 71.676
R1053 B.n307 B.n306 71.676
R1054 B.n300 B.n251 71.676
R1055 B.n299 B.n298 71.676
R1056 B.n292 B.n253 71.676
R1057 B.n291 B.n290 71.676
R1058 B.n284 B.n255 71.676
R1059 B.n283 B.n282 71.676
R1060 B.n276 B.n257 71.676
R1061 B.n275 B.n274 71.676
R1062 B.n268 B.n259 71.676
R1063 B.n267 B.n266 71.676
R1064 B.n262 B.n261 71.676
R1065 B.n801 B.n79 71.676
R1066 B.n800 B.n799 71.676
R1067 B.n793 B.n81 71.676
R1068 B.n792 B.n791 71.676
R1069 B.n785 B.n83 71.676
R1070 B.n784 B.n783 71.676
R1071 B.n777 B.n85 71.676
R1072 B.n776 B.n775 71.676
R1073 B.n769 B.n87 71.676
R1074 B.n768 B.n767 71.676
R1075 B.n761 B.n89 71.676
R1076 B.n760 B.n759 71.676
R1077 B.n753 B.n91 71.676
R1078 B.n752 B.n751 71.676
R1079 B.n745 B.n93 71.676
R1080 B.n744 B.n743 71.676
R1081 B.n737 B.n95 71.676
R1082 B.n736 B.n735 71.676
R1083 B.n729 B.n97 71.676
R1084 B.n728 B.n727 71.676
R1085 B.n720 B.n99 71.676
R1086 B.n719 B.n718 71.676
R1087 B.n712 B.n103 71.676
R1088 B.n711 B.n710 71.676
R1089 B.n704 B.n105 71.676
R1090 B.n703 B.n109 71.676
R1091 B.n699 B.n698 71.676
R1092 B.n692 B.n111 71.676
R1093 B.n691 B.n690 71.676
R1094 B.n684 B.n113 71.676
R1095 B.n683 B.n682 71.676
R1096 B.n676 B.n115 71.676
R1097 B.n675 B.n674 71.676
R1098 B.n668 B.n117 71.676
R1099 B.n667 B.n666 71.676
R1100 B.n660 B.n119 71.676
R1101 B.n659 B.n658 71.676
R1102 B.n652 B.n121 71.676
R1103 B.n651 B.n650 71.676
R1104 B.n644 B.n123 71.676
R1105 B.n643 B.n642 71.676
R1106 B.n636 B.n125 71.676
R1107 B.n635 B.n634 71.676
R1108 B.n628 B.n127 71.676
R1109 B.n627 B.n626 71.676
R1110 B.n626 B.n625 71.676
R1111 B.n629 B.n628 71.676
R1112 B.n634 B.n633 71.676
R1113 B.n637 B.n636 71.676
R1114 B.n642 B.n641 71.676
R1115 B.n645 B.n644 71.676
R1116 B.n650 B.n649 71.676
R1117 B.n653 B.n652 71.676
R1118 B.n658 B.n657 71.676
R1119 B.n661 B.n660 71.676
R1120 B.n666 B.n665 71.676
R1121 B.n669 B.n668 71.676
R1122 B.n674 B.n673 71.676
R1123 B.n677 B.n676 71.676
R1124 B.n682 B.n681 71.676
R1125 B.n685 B.n684 71.676
R1126 B.n690 B.n689 71.676
R1127 B.n693 B.n692 71.676
R1128 B.n698 B.n697 71.676
R1129 B.n700 B.n109 71.676
R1130 B.n705 B.n704 71.676
R1131 B.n710 B.n709 71.676
R1132 B.n713 B.n712 71.676
R1133 B.n718 B.n717 71.676
R1134 B.n721 B.n720 71.676
R1135 B.n727 B.n726 71.676
R1136 B.n730 B.n729 71.676
R1137 B.n735 B.n734 71.676
R1138 B.n738 B.n737 71.676
R1139 B.n743 B.n742 71.676
R1140 B.n746 B.n745 71.676
R1141 B.n751 B.n750 71.676
R1142 B.n754 B.n753 71.676
R1143 B.n759 B.n758 71.676
R1144 B.n762 B.n761 71.676
R1145 B.n767 B.n766 71.676
R1146 B.n770 B.n769 71.676
R1147 B.n775 B.n774 71.676
R1148 B.n778 B.n777 71.676
R1149 B.n783 B.n782 71.676
R1150 B.n786 B.n785 71.676
R1151 B.n791 B.n790 71.676
R1152 B.n794 B.n793 71.676
R1153 B.n799 B.n798 71.676
R1154 B.n802 B.n801 71.676
R1155 B.n439 B.n438 71.676
R1156 B.n433 B.n213 71.676
R1157 B.n431 B.n430 71.676
R1158 B.n426 B.n425 71.676
R1159 B.n423 B.n422 71.676
R1160 B.n418 B.n417 71.676
R1161 B.n415 B.n414 71.676
R1162 B.n410 B.n409 71.676
R1163 B.n407 B.n406 71.676
R1164 B.n402 B.n401 71.676
R1165 B.n399 B.n398 71.676
R1166 B.n394 B.n393 71.676
R1167 B.n391 B.n390 71.676
R1168 B.n386 B.n385 71.676
R1169 B.n383 B.n382 71.676
R1170 B.n378 B.n377 71.676
R1171 B.n375 B.n374 71.676
R1172 B.n370 B.n369 71.676
R1173 B.n367 B.n366 71.676
R1174 B.n362 B.n361 71.676
R1175 B.n357 B.n235 71.676
R1176 B.n355 B.n354 71.676
R1177 B.n350 B.n349 71.676
R1178 B.n347 B.n346 71.676
R1179 B.n341 B.n340 71.676
R1180 B.n338 B.n337 71.676
R1181 B.n333 B.n332 71.676
R1182 B.n330 B.n329 71.676
R1183 B.n325 B.n324 71.676
R1184 B.n322 B.n321 71.676
R1185 B.n317 B.n316 71.676
R1186 B.n314 B.n313 71.676
R1187 B.n309 B.n308 71.676
R1188 B.n306 B.n305 71.676
R1189 B.n301 B.n300 71.676
R1190 B.n298 B.n297 71.676
R1191 B.n293 B.n292 71.676
R1192 B.n290 B.n289 71.676
R1193 B.n285 B.n284 71.676
R1194 B.n282 B.n281 71.676
R1195 B.n277 B.n276 71.676
R1196 B.n274 B.n273 71.676
R1197 B.n269 B.n268 71.676
R1198 B.n266 B.n265 71.676
R1199 B.n261 B.n209 71.676
R1200 B.n241 B.t10 70.3544
R1201 B.n107 B.t15 70.3544
R1202 B.n233 B.t17 70.3396
R1203 B.n101 B.t21 70.3396
R1204 B.n343 B.n241 59.5399
R1205 B.n234 B.n233 59.5399
R1206 B.n723 B.n101 59.5399
R1207 B.n108 B.n107 59.5399
R1208 B.n241 B.n240 44.8005
R1209 B.n233 B.n232 44.8005
R1210 B.n101 B.n100 44.8005
R1211 B.n107 B.n106 44.8005
R1212 B.n444 B.n206 44.0913
R1213 B.n450 B.n206 44.0913
R1214 B.n450 B.n202 44.0913
R1215 B.n456 B.n202 44.0913
R1216 B.n456 B.n198 44.0913
R1217 B.n462 B.n198 44.0913
R1218 B.n468 B.n194 44.0913
R1219 B.n468 B.n190 44.0913
R1220 B.n474 B.n190 44.0913
R1221 B.n474 B.n186 44.0913
R1222 B.n480 B.n186 44.0913
R1223 B.n480 B.n182 44.0913
R1224 B.n486 B.n182 44.0913
R1225 B.n486 B.n178 44.0913
R1226 B.n492 B.n178 44.0913
R1227 B.n498 B.n174 44.0913
R1228 B.n498 B.n170 44.0913
R1229 B.n504 B.n170 44.0913
R1230 B.n504 B.n166 44.0913
R1231 B.n511 B.n166 44.0913
R1232 B.n511 B.n510 44.0913
R1233 B.n517 B.n159 44.0913
R1234 B.n523 B.n159 44.0913
R1235 B.n523 B.n155 44.0913
R1236 B.n529 B.n155 44.0913
R1237 B.n529 B.n151 44.0913
R1238 B.n535 B.n151 44.0913
R1239 B.n541 B.n147 44.0913
R1240 B.n541 B.n143 44.0913
R1241 B.n547 B.n143 44.0913
R1242 B.n547 B.n139 44.0913
R1243 B.n553 B.n139 44.0913
R1244 B.n553 B.t5 44.0913
R1245 B.n560 B.t5 44.0913
R1246 B.n560 B.n132 44.0913
R1247 B.n566 B.n132 44.0913
R1248 B.n566 B.n4 44.0913
R1249 B.n888 B.n4 44.0913
R1250 B.n888 B.n887 44.0913
R1251 B.n887 B.n886 44.0913
R1252 B.n886 B.n8 44.0913
R1253 B.n880 B.n8 44.0913
R1254 B.n880 B.t0 44.0913
R1255 B.t0 B.n879 44.0913
R1256 B.n879 B.n15 44.0913
R1257 B.n873 B.n15 44.0913
R1258 B.n873 B.n872 44.0913
R1259 B.n872 B.n871 44.0913
R1260 B.n871 B.n22 44.0913
R1261 B.n865 B.n864 44.0913
R1262 B.n864 B.n863 44.0913
R1263 B.n863 B.n29 44.0913
R1264 B.n857 B.n29 44.0913
R1265 B.n857 B.n856 44.0913
R1266 B.n856 B.n855 44.0913
R1267 B.n849 B.n39 44.0913
R1268 B.n849 B.n848 44.0913
R1269 B.n848 B.n847 44.0913
R1270 B.n847 B.n43 44.0913
R1271 B.n841 B.n43 44.0913
R1272 B.n841 B.n840 44.0913
R1273 B.n839 B.n50 44.0913
R1274 B.n833 B.n50 44.0913
R1275 B.n833 B.n832 44.0913
R1276 B.n832 B.n831 44.0913
R1277 B.n831 B.n57 44.0913
R1278 B.n825 B.n57 44.0913
R1279 B.n825 B.n824 44.0913
R1280 B.n824 B.n823 44.0913
R1281 B.n823 B.n64 44.0913
R1282 B.n817 B.n816 44.0913
R1283 B.n816 B.n815 44.0913
R1284 B.n815 B.n71 44.0913
R1285 B.n809 B.n71 44.0913
R1286 B.n809 B.n808 44.0913
R1287 B.n808 B.n807 44.0913
R1288 B.t6 B.n147 35.0138
R1289 B.t7 B.n22 35.0138
R1290 B.n805 B.n804 33.2493
R1291 B.n623 B.n622 33.2493
R1292 B.n446 B.n208 33.2493
R1293 B.n442 B.n441 33.2493
R1294 B.n462 B.t9 27.233
R1295 B.n492 B.t1 27.233
R1296 B.t2 B.n839 27.233
R1297 B.n817 B.t13 27.233
R1298 B.n517 B.t3 25.9362
R1299 B.n855 B.t4 25.9362
R1300 B.n510 B.t3 18.1555
R1301 B.n39 B.t4 18.1555
R1302 B B.n890 18.0485
R1303 B.t9 B.n194 16.8587
R1304 B.t1 B.n174 16.8587
R1305 B.n840 B.t2 16.8587
R1306 B.t13 B.n64 16.8587
R1307 B.n804 B.n803 10.6151
R1308 B.n803 B.n80 10.6151
R1309 B.n797 B.n80 10.6151
R1310 B.n797 B.n796 10.6151
R1311 B.n796 B.n795 10.6151
R1312 B.n795 B.n82 10.6151
R1313 B.n789 B.n82 10.6151
R1314 B.n789 B.n788 10.6151
R1315 B.n788 B.n787 10.6151
R1316 B.n787 B.n84 10.6151
R1317 B.n781 B.n84 10.6151
R1318 B.n781 B.n780 10.6151
R1319 B.n780 B.n779 10.6151
R1320 B.n779 B.n86 10.6151
R1321 B.n773 B.n86 10.6151
R1322 B.n773 B.n772 10.6151
R1323 B.n772 B.n771 10.6151
R1324 B.n771 B.n88 10.6151
R1325 B.n765 B.n88 10.6151
R1326 B.n765 B.n764 10.6151
R1327 B.n764 B.n763 10.6151
R1328 B.n763 B.n90 10.6151
R1329 B.n757 B.n90 10.6151
R1330 B.n757 B.n756 10.6151
R1331 B.n756 B.n755 10.6151
R1332 B.n755 B.n92 10.6151
R1333 B.n749 B.n92 10.6151
R1334 B.n749 B.n748 10.6151
R1335 B.n748 B.n747 10.6151
R1336 B.n747 B.n94 10.6151
R1337 B.n741 B.n94 10.6151
R1338 B.n741 B.n740 10.6151
R1339 B.n740 B.n739 10.6151
R1340 B.n739 B.n96 10.6151
R1341 B.n733 B.n96 10.6151
R1342 B.n733 B.n732 10.6151
R1343 B.n732 B.n731 10.6151
R1344 B.n731 B.n98 10.6151
R1345 B.n725 B.n98 10.6151
R1346 B.n725 B.n724 10.6151
R1347 B.n722 B.n102 10.6151
R1348 B.n716 B.n102 10.6151
R1349 B.n716 B.n715 10.6151
R1350 B.n715 B.n714 10.6151
R1351 B.n714 B.n104 10.6151
R1352 B.n708 B.n104 10.6151
R1353 B.n708 B.n707 10.6151
R1354 B.n707 B.n706 10.6151
R1355 B.n702 B.n701 10.6151
R1356 B.n701 B.n110 10.6151
R1357 B.n696 B.n110 10.6151
R1358 B.n696 B.n695 10.6151
R1359 B.n695 B.n694 10.6151
R1360 B.n694 B.n112 10.6151
R1361 B.n688 B.n112 10.6151
R1362 B.n688 B.n687 10.6151
R1363 B.n687 B.n686 10.6151
R1364 B.n686 B.n114 10.6151
R1365 B.n680 B.n114 10.6151
R1366 B.n680 B.n679 10.6151
R1367 B.n679 B.n678 10.6151
R1368 B.n678 B.n116 10.6151
R1369 B.n672 B.n116 10.6151
R1370 B.n672 B.n671 10.6151
R1371 B.n671 B.n670 10.6151
R1372 B.n670 B.n118 10.6151
R1373 B.n664 B.n118 10.6151
R1374 B.n664 B.n663 10.6151
R1375 B.n663 B.n662 10.6151
R1376 B.n662 B.n120 10.6151
R1377 B.n656 B.n120 10.6151
R1378 B.n656 B.n655 10.6151
R1379 B.n655 B.n654 10.6151
R1380 B.n654 B.n122 10.6151
R1381 B.n648 B.n122 10.6151
R1382 B.n648 B.n647 10.6151
R1383 B.n647 B.n646 10.6151
R1384 B.n646 B.n124 10.6151
R1385 B.n640 B.n124 10.6151
R1386 B.n640 B.n639 10.6151
R1387 B.n639 B.n638 10.6151
R1388 B.n638 B.n126 10.6151
R1389 B.n632 B.n126 10.6151
R1390 B.n632 B.n631 10.6151
R1391 B.n631 B.n630 10.6151
R1392 B.n630 B.n128 10.6151
R1393 B.n624 B.n128 10.6151
R1394 B.n624 B.n623 10.6151
R1395 B.n447 B.n446 10.6151
R1396 B.n448 B.n447 10.6151
R1397 B.n448 B.n200 10.6151
R1398 B.n458 B.n200 10.6151
R1399 B.n459 B.n458 10.6151
R1400 B.n460 B.n459 10.6151
R1401 B.n460 B.n192 10.6151
R1402 B.n470 B.n192 10.6151
R1403 B.n471 B.n470 10.6151
R1404 B.n472 B.n471 10.6151
R1405 B.n472 B.n184 10.6151
R1406 B.n482 B.n184 10.6151
R1407 B.n483 B.n482 10.6151
R1408 B.n484 B.n483 10.6151
R1409 B.n484 B.n176 10.6151
R1410 B.n494 B.n176 10.6151
R1411 B.n495 B.n494 10.6151
R1412 B.n496 B.n495 10.6151
R1413 B.n496 B.n168 10.6151
R1414 B.n506 B.n168 10.6151
R1415 B.n507 B.n506 10.6151
R1416 B.n508 B.n507 10.6151
R1417 B.n508 B.n161 10.6151
R1418 B.n519 B.n161 10.6151
R1419 B.n520 B.n519 10.6151
R1420 B.n521 B.n520 10.6151
R1421 B.n521 B.n153 10.6151
R1422 B.n531 B.n153 10.6151
R1423 B.n532 B.n531 10.6151
R1424 B.n533 B.n532 10.6151
R1425 B.n533 B.n145 10.6151
R1426 B.n543 B.n145 10.6151
R1427 B.n544 B.n543 10.6151
R1428 B.n545 B.n544 10.6151
R1429 B.n545 B.n137 10.6151
R1430 B.n555 B.n137 10.6151
R1431 B.n556 B.n555 10.6151
R1432 B.n558 B.n556 10.6151
R1433 B.n558 B.n557 10.6151
R1434 B.n557 B.n130 10.6151
R1435 B.n569 B.n130 10.6151
R1436 B.n570 B.n569 10.6151
R1437 B.n571 B.n570 10.6151
R1438 B.n572 B.n571 10.6151
R1439 B.n574 B.n572 10.6151
R1440 B.n575 B.n574 10.6151
R1441 B.n576 B.n575 10.6151
R1442 B.n577 B.n576 10.6151
R1443 B.n579 B.n577 10.6151
R1444 B.n580 B.n579 10.6151
R1445 B.n581 B.n580 10.6151
R1446 B.n582 B.n581 10.6151
R1447 B.n584 B.n582 10.6151
R1448 B.n585 B.n584 10.6151
R1449 B.n586 B.n585 10.6151
R1450 B.n587 B.n586 10.6151
R1451 B.n589 B.n587 10.6151
R1452 B.n590 B.n589 10.6151
R1453 B.n591 B.n590 10.6151
R1454 B.n592 B.n591 10.6151
R1455 B.n594 B.n592 10.6151
R1456 B.n595 B.n594 10.6151
R1457 B.n596 B.n595 10.6151
R1458 B.n597 B.n596 10.6151
R1459 B.n599 B.n597 10.6151
R1460 B.n600 B.n599 10.6151
R1461 B.n601 B.n600 10.6151
R1462 B.n602 B.n601 10.6151
R1463 B.n604 B.n602 10.6151
R1464 B.n605 B.n604 10.6151
R1465 B.n606 B.n605 10.6151
R1466 B.n607 B.n606 10.6151
R1467 B.n609 B.n607 10.6151
R1468 B.n610 B.n609 10.6151
R1469 B.n611 B.n610 10.6151
R1470 B.n612 B.n611 10.6151
R1471 B.n614 B.n612 10.6151
R1472 B.n615 B.n614 10.6151
R1473 B.n616 B.n615 10.6151
R1474 B.n617 B.n616 10.6151
R1475 B.n619 B.n617 10.6151
R1476 B.n620 B.n619 10.6151
R1477 B.n621 B.n620 10.6151
R1478 B.n622 B.n621 10.6151
R1479 B.n441 B.n440 10.6151
R1480 B.n440 B.n212 10.6151
R1481 B.n435 B.n212 10.6151
R1482 B.n435 B.n434 10.6151
R1483 B.n434 B.n214 10.6151
R1484 B.n429 B.n214 10.6151
R1485 B.n429 B.n428 10.6151
R1486 B.n428 B.n427 10.6151
R1487 B.n427 B.n216 10.6151
R1488 B.n421 B.n216 10.6151
R1489 B.n421 B.n420 10.6151
R1490 B.n420 B.n419 10.6151
R1491 B.n419 B.n218 10.6151
R1492 B.n413 B.n218 10.6151
R1493 B.n413 B.n412 10.6151
R1494 B.n412 B.n411 10.6151
R1495 B.n411 B.n220 10.6151
R1496 B.n405 B.n220 10.6151
R1497 B.n405 B.n404 10.6151
R1498 B.n404 B.n403 10.6151
R1499 B.n403 B.n222 10.6151
R1500 B.n397 B.n222 10.6151
R1501 B.n397 B.n396 10.6151
R1502 B.n396 B.n395 10.6151
R1503 B.n395 B.n224 10.6151
R1504 B.n389 B.n224 10.6151
R1505 B.n389 B.n388 10.6151
R1506 B.n388 B.n387 10.6151
R1507 B.n387 B.n226 10.6151
R1508 B.n381 B.n226 10.6151
R1509 B.n381 B.n380 10.6151
R1510 B.n380 B.n379 10.6151
R1511 B.n379 B.n228 10.6151
R1512 B.n373 B.n228 10.6151
R1513 B.n373 B.n372 10.6151
R1514 B.n372 B.n371 10.6151
R1515 B.n371 B.n230 10.6151
R1516 B.n365 B.n230 10.6151
R1517 B.n365 B.n364 10.6151
R1518 B.n364 B.n363 10.6151
R1519 B.n359 B.n358 10.6151
R1520 B.n358 B.n236 10.6151
R1521 B.n353 B.n236 10.6151
R1522 B.n353 B.n352 10.6151
R1523 B.n352 B.n351 10.6151
R1524 B.n351 B.n238 10.6151
R1525 B.n345 B.n238 10.6151
R1526 B.n345 B.n344 10.6151
R1527 B.n342 B.n242 10.6151
R1528 B.n336 B.n242 10.6151
R1529 B.n336 B.n335 10.6151
R1530 B.n335 B.n334 10.6151
R1531 B.n334 B.n244 10.6151
R1532 B.n328 B.n244 10.6151
R1533 B.n328 B.n327 10.6151
R1534 B.n327 B.n326 10.6151
R1535 B.n326 B.n246 10.6151
R1536 B.n320 B.n246 10.6151
R1537 B.n320 B.n319 10.6151
R1538 B.n319 B.n318 10.6151
R1539 B.n318 B.n248 10.6151
R1540 B.n312 B.n248 10.6151
R1541 B.n312 B.n311 10.6151
R1542 B.n311 B.n310 10.6151
R1543 B.n310 B.n250 10.6151
R1544 B.n304 B.n250 10.6151
R1545 B.n304 B.n303 10.6151
R1546 B.n303 B.n302 10.6151
R1547 B.n302 B.n252 10.6151
R1548 B.n296 B.n252 10.6151
R1549 B.n296 B.n295 10.6151
R1550 B.n295 B.n294 10.6151
R1551 B.n294 B.n254 10.6151
R1552 B.n288 B.n254 10.6151
R1553 B.n288 B.n287 10.6151
R1554 B.n287 B.n286 10.6151
R1555 B.n286 B.n256 10.6151
R1556 B.n280 B.n256 10.6151
R1557 B.n280 B.n279 10.6151
R1558 B.n279 B.n278 10.6151
R1559 B.n278 B.n258 10.6151
R1560 B.n272 B.n258 10.6151
R1561 B.n272 B.n271 10.6151
R1562 B.n271 B.n270 10.6151
R1563 B.n270 B.n260 10.6151
R1564 B.n264 B.n260 10.6151
R1565 B.n264 B.n263 10.6151
R1566 B.n263 B.n208 10.6151
R1567 B.n442 B.n204 10.6151
R1568 B.n452 B.n204 10.6151
R1569 B.n453 B.n452 10.6151
R1570 B.n454 B.n453 10.6151
R1571 B.n454 B.n196 10.6151
R1572 B.n464 B.n196 10.6151
R1573 B.n465 B.n464 10.6151
R1574 B.n466 B.n465 10.6151
R1575 B.n466 B.n188 10.6151
R1576 B.n476 B.n188 10.6151
R1577 B.n477 B.n476 10.6151
R1578 B.n478 B.n477 10.6151
R1579 B.n478 B.n180 10.6151
R1580 B.n488 B.n180 10.6151
R1581 B.n489 B.n488 10.6151
R1582 B.n490 B.n489 10.6151
R1583 B.n490 B.n172 10.6151
R1584 B.n500 B.n172 10.6151
R1585 B.n501 B.n500 10.6151
R1586 B.n502 B.n501 10.6151
R1587 B.n502 B.n164 10.6151
R1588 B.n513 B.n164 10.6151
R1589 B.n514 B.n513 10.6151
R1590 B.n515 B.n514 10.6151
R1591 B.n515 B.n157 10.6151
R1592 B.n525 B.n157 10.6151
R1593 B.n526 B.n525 10.6151
R1594 B.n527 B.n526 10.6151
R1595 B.n527 B.n149 10.6151
R1596 B.n537 B.n149 10.6151
R1597 B.n538 B.n537 10.6151
R1598 B.n539 B.n538 10.6151
R1599 B.n539 B.n141 10.6151
R1600 B.n549 B.n141 10.6151
R1601 B.n550 B.n549 10.6151
R1602 B.n551 B.n550 10.6151
R1603 B.n551 B.n134 10.6151
R1604 B.n562 B.n134 10.6151
R1605 B.n563 B.n562 10.6151
R1606 B.n564 B.n563 10.6151
R1607 B.n564 B.n0 10.6151
R1608 B.n884 B.n1 10.6151
R1609 B.n884 B.n883 10.6151
R1610 B.n883 B.n882 10.6151
R1611 B.n882 B.n10 10.6151
R1612 B.n877 B.n10 10.6151
R1613 B.n877 B.n876 10.6151
R1614 B.n876 B.n875 10.6151
R1615 B.n875 B.n17 10.6151
R1616 B.n869 B.n17 10.6151
R1617 B.n869 B.n868 10.6151
R1618 B.n868 B.n867 10.6151
R1619 B.n867 B.n24 10.6151
R1620 B.n861 B.n24 10.6151
R1621 B.n861 B.n860 10.6151
R1622 B.n860 B.n859 10.6151
R1623 B.n859 B.n31 10.6151
R1624 B.n853 B.n31 10.6151
R1625 B.n853 B.n852 10.6151
R1626 B.n852 B.n851 10.6151
R1627 B.n851 B.n37 10.6151
R1628 B.n845 B.n37 10.6151
R1629 B.n845 B.n844 10.6151
R1630 B.n844 B.n843 10.6151
R1631 B.n843 B.n45 10.6151
R1632 B.n837 B.n45 10.6151
R1633 B.n837 B.n836 10.6151
R1634 B.n836 B.n835 10.6151
R1635 B.n835 B.n52 10.6151
R1636 B.n829 B.n52 10.6151
R1637 B.n829 B.n828 10.6151
R1638 B.n828 B.n827 10.6151
R1639 B.n827 B.n59 10.6151
R1640 B.n821 B.n59 10.6151
R1641 B.n821 B.n820 10.6151
R1642 B.n820 B.n819 10.6151
R1643 B.n819 B.n66 10.6151
R1644 B.n813 B.n66 10.6151
R1645 B.n813 B.n812 10.6151
R1646 B.n812 B.n811 10.6151
R1647 B.n811 B.n73 10.6151
R1648 B.n805 B.n73 10.6151
R1649 B.n535 B.t6 9.07801
R1650 B.n865 B.t7 9.07801
R1651 B.n723 B.n722 6.5566
R1652 B.n706 B.n108 6.5566
R1653 B.n359 B.n234 6.5566
R1654 B.n344 B.n343 6.5566
R1655 B.n724 B.n723 4.05904
R1656 B.n702 B.n108 4.05904
R1657 B.n363 B.n234 4.05904
R1658 B.n343 B.n342 4.05904
R1659 B.n890 B.n0 2.81026
R1660 B.n890 B.n1 2.81026
R1661 VN.n5 VN.t2 173.139
R1662 VN.n28 VN.t5 173.139
R1663 VN.n43 VN.n23 161.3
R1664 VN.n42 VN.n41 161.3
R1665 VN.n40 VN.n24 161.3
R1666 VN.n39 VN.n38 161.3
R1667 VN.n36 VN.n25 161.3
R1668 VN.n35 VN.n34 161.3
R1669 VN.n33 VN.n26 161.3
R1670 VN.n32 VN.n31 161.3
R1671 VN.n30 VN.n27 161.3
R1672 VN.n20 VN.n0 161.3
R1673 VN.n19 VN.n18 161.3
R1674 VN.n17 VN.n1 161.3
R1675 VN.n16 VN.n15 161.3
R1676 VN.n13 VN.n2 161.3
R1677 VN.n12 VN.n11 161.3
R1678 VN.n10 VN.n3 161.3
R1679 VN.n9 VN.n8 161.3
R1680 VN.n7 VN.n4 161.3
R1681 VN.n6 VN.t7 142.287
R1682 VN.n14 VN.t6 142.287
R1683 VN.n21 VN.t4 142.287
R1684 VN.n29 VN.t3 142.287
R1685 VN.n37 VN.t1 142.287
R1686 VN.n44 VN.t0 142.287
R1687 VN.n22 VN.n21 88.0021
R1688 VN.n45 VN.n44 88.0021
R1689 VN.n6 VN.n5 62.6111
R1690 VN.n29 VN.n28 62.6111
R1691 VN.n19 VN.n1 56.5193
R1692 VN.n42 VN.n24 56.5193
R1693 VN VN.n45 48.1042
R1694 VN.n8 VN.n3 40.4934
R1695 VN.n12 VN.n3 40.4934
R1696 VN.n31 VN.n26 40.4934
R1697 VN.n35 VN.n26 40.4934
R1698 VN.n8 VN.n7 24.4675
R1699 VN.n13 VN.n12 24.4675
R1700 VN.n15 VN.n1 24.4675
R1701 VN.n20 VN.n19 24.4675
R1702 VN.n31 VN.n30 24.4675
R1703 VN.n38 VN.n24 24.4675
R1704 VN.n36 VN.n35 24.4675
R1705 VN.n43 VN.n42 24.4675
R1706 VN.n21 VN.n20 22.7548
R1707 VN.n44 VN.n43 22.7548
R1708 VN.n15 VN.n14 16.8827
R1709 VN.n38 VN.n37 16.8827
R1710 VN.n28 VN.n27 12.915
R1711 VN.n5 VN.n4 12.915
R1712 VN.n7 VN.n6 7.58527
R1713 VN.n14 VN.n13 7.58527
R1714 VN.n30 VN.n29 7.58527
R1715 VN.n37 VN.n36 7.58527
R1716 VN.n45 VN.n23 0.278367
R1717 VN.n22 VN.n0 0.278367
R1718 VN.n41 VN.n23 0.189894
R1719 VN.n41 VN.n40 0.189894
R1720 VN.n40 VN.n39 0.189894
R1721 VN.n39 VN.n25 0.189894
R1722 VN.n34 VN.n25 0.189894
R1723 VN.n34 VN.n33 0.189894
R1724 VN.n33 VN.n32 0.189894
R1725 VN.n32 VN.n27 0.189894
R1726 VN.n9 VN.n4 0.189894
R1727 VN.n10 VN.n9 0.189894
R1728 VN.n11 VN.n10 0.189894
R1729 VN.n11 VN.n2 0.189894
R1730 VN.n16 VN.n2 0.189894
R1731 VN.n17 VN.n16 0.189894
R1732 VN.n18 VN.n17 0.189894
R1733 VN.n18 VN.n0 0.189894
R1734 VN VN.n22 0.153454
R1735 VDD2.n2 VDD2.n1 61.5626
R1736 VDD2.n2 VDD2.n0 61.5626
R1737 VDD2 VDD2.n5 61.5598
R1738 VDD2.n4 VDD2.n3 60.6225
R1739 VDD2.n4 VDD2.n2 42.7541
R1740 VDD2.n5 VDD2.t4 1.69426
R1741 VDD2.n5 VDD2.t2 1.69426
R1742 VDD2.n3 VDD2.t7 1.69426
R1743 VDD2.n3 VDD2.t6 1.69426
R1744 VDD2.n1 VDD2.t1 1.69426
R1745 VDD2.n1 VDD2.t3 1.69426
R1746 VDD2.n0 VDD2.t5 1.69426
R1747 VDD2.n0 VDD2.t0 1.69426
R1748 VDD2 VDD2.n4 1.05438
C0 VDD2 VDD1 1.45537f
C1 VP VDD2 0.453781f
C2 VP VDD1 8.27846f
C3 VN VTAIL 8.19542f
C4 VTAIL VDD2 8.03961f
C5 VTAIL VDD1 7.98935f
C6 VP VTAIL 8.209531f
C7 VN VDD2 7.97645f
C8 VN VDD1 0.150692f
C9 VP VN 6.84695f
C10 VDD2 B 4.732636f
C11 VDD1 B 5.104959f
C12 VTAIL B 9.855159f
C13 VN B 13.13643f
C14 VP B 11.642154f
C15 VDD2.t5 B 0.226636f
C16 VDD2.t0 B 0.226636f
C17 VDD2.n0 B 2.02146f
C18 VDD2.t1 B 0.226636f
C19 VDD2.t3 B 0.226636f
C20 VDD2.n1 B 2.02146f
C21 VDD2.n2 B 2.84893f
C22 VDD2.t7 B 0.226636f
C23 VDD2.t6 B 0.226636f
C24 VDD2.n3 B 2.01464f
C25 VDD2.n4 B 2.66268f
C26 VDD2.t4 B 0.226636f
C27 VDD2.t2 B 0.226636f
C28 VDD2.n5 B 2.02142f
C29 VN.n0 B 0.034684f
C30 VN.t4 B 1.65782f
C31 VN.n1 B 0.042803f
C32 VN.n2 B 0.026308f
C33 VN.t6 B 1.65782f
C34 VN.n3 B 0.021267f
C35 VN.n4 B 0.196398f
C36 VN.t7 B 1.65782f
C37 VN.t2 B 1.78675f
C38 VN.n5 B 0.6613f
C39 VN.n6 B 0.651313f
C40 VN.n7 B 0.032327f
C41 VN.n8 B 0.052286f
C42 VN.n9 B 0.026308f
C43 VN.n10 B 0.026308f
C44 VN.n11 B 0.026308f
C45 VN.n12 B 0.052286f
C46 VN.n13 B 0.032327f
C47 VN.n14 B 0.593032f
C48 VN.n15 B 0.041526f
C49 VN.n16 B 0.026308f
C50 VN.n17 B 0.026308f
C51 VN.n18 B 0.026308f
C52 VN.n19 B 0.034006f
C53 VN.n20 B 0.047335f
C54 VN.n21 B 0.677678f
C55 VN.n22 B 0.02946f
C56 VN.n23 B 0.034684f
C57 VN.t0 B 1.65782f
C58 VN.n24 B 0.042803f
C59 VN.n25 B 0.026308f
C60 VN.t1 B 1.65782f
C61 VN.n26 B 0.021267f
C62 VN.n27 B 0.196398f
C63 VN.t3 B 1.65782f
C64 VN.t5 B 1.78675f
C65 VN.n28 B 0.6613f
C66 VN.n29 B 0.651313f
C67 VN.n30 B 0.032327f
C68 VN.n31 B 0.052286f
C69 VN.n32 B 0.026308f
C70 VN.n33 B 0.026308f
C71 VN.n34 B 0.026308f
C72 VN.n35 B 0.052286f
C73 VN.n36 B 0.032327f
C74 VN.n37 B 0.593032f
C75 VN.n38 B 0.041526f
C76 VN.n39 B 0.026308f
C77 VN.n40 B 0.026308f
C78 VN.n41 B 0.026308f
C79 VN.n42 B 0.034006f
C80 VN.n43 B 0.047335f
C81 VN.n44 B 0.677678f
C82 VN.n45 B 1.37091f
C83 VDD1.t2 B 0.229585f
C84 VDD1.t5 B 0.229585f
C85 VDD1.n0 B 2.04873f
C86 VDD1.t4 B 0.229585f
C87 VDD1.t3 B 0.229585f
C88 VDD1.n1 B 2.04776f
C89 VDD1.t0 B 0.229585f
C90 VDD1.t7 B 0.229585f
C91 VDD1.n2 B 2.04776f
C92 VDD1.n3 B 2.93814f
C93 VDD1.t6 B 0.229585f
C94 VDD1.t1 B 0.229585f
C95 VDD1.n4 B 2.04085f
C96 VDD1.n5 B 2.72767f
C97 VTAIL.t15 B 0.17997f
C98 VTAIL.t4 B 0.17997f
C99 VTAIL.n0 B 1.53965f
C100 VTAIL.n1 B 0.324548f
C101 VTAIL.t0 B 1.9618f
C102 VTAIL.n2 B 0.419069f
C103 VTAIL.t12 B 1.9618f
C104 VTAIL.n3 B 0.419069f
C105 VTAIL.t11 B 0.17997f
C106 VTAIL.t10 B 0.17997f
C107 VTAIL.n4 B 1.53965f
C108 VTAIL.n5 B 0.445905f
C109 VTAIL.t8 B 1.9618f
C110 VTAIL.n6 B 1.41185f
C111 VTAIL.t1 B 1.9618f
C112 VTAIL.n7 B 1.41184f
C113 VTAIL.t3 B 0.17997f
C114 VTAIL.t6 B 0.17997f
C115 VTAIL.n8 B 1.53965f
C116 VTAIL.n9 B 0.4459f
C117 VTAIL.t5 B 1.9618f
C118 VTAIL.n10 B 0.419063f
C119 VTAIL.t7 B 1.9618f
C120 VTAIL.n11 B 0.419063f
C121 VTAIL.t13 B 0.17997f
C122 VTAIL.t14 B 0.17997f
C123 VTAIL.n12 B 1.53965f
C124 VTAIL.n13 B 0.4459f
C125 VTAIL.t9 B 1.9618f
C126 VTAIL.n14 B 1.41185f
C127 VTAIL.t2 B 1.9618f
C128 VTAIL.n15 B 1.40819f
C129 VP.n0 B 0.035193f
C130 VP.t0 B 1.68215f
C131 VP.n1 B 0.043431f
C132 VP.n2 B 0.026694f
C133 VP.t7 B 1.68215f
C134 VP.n3 B 0.021579f
C135 VP.n4 B 0.026694f
C136 VP.t4 B 1.68215f
C137 VP.n5 B 0.043431f
C138 VP.n6 B 0.035193f
C139 VP.t3 B 1.68215f
C140 VP.n7 B 0.035193f
C141 VP.t6 B 1.68215f
C142 VP.n8 B 0.043431f
C143 VP.n9 B 0.026694f
C144 VP.t1 B 1.68215f
C145 VP.n10 B 0.021579f
C146 VP.n11 B 0.19928f
C147 VP.t2 B 1.68215f
C148 VP.t5 B 1.81297f
C149 VP.n12 B 0.671004f
C150 VP.n13 B 0.660871f
C151 VP.n14 B 0.032801f
C152 VP.n15 B 0.053054f
C153 VP.n16 B 0.026694f
C154 VP.n17 B 0.026694f
C155 VP.n18 B 0.026694f
C156 VP.n19 B 0.053054f
C157 VP.n20 B 0.032801f
C158 VP.n21 B 0.601735f
C159 VP.n22 B 0.042135f
C160 VP.n23 B 0.026694f
C161 VP.n24 B 0.026694f
C162 VP.n25 B 0.026694f
C163 VP.n26 B 0.034505f
C164 VP.n27 B 0.04803f
C165 VP.n28 B 0.687623f
C166 VP.n29 B 1.37658f
C167 VP.n30 B 1.39665f
C168 VP.n31 B 0.687623f
C169 VP.n32 B 0.04803f
C170 VP.n33 B 0.034505f
C171 VP.n34 B 0.026694f
C172 VP.n35 B 0.026694f
C173 VP.n36 B 0.026694f
C174 VP.n37 B 0.042135f
C175 VP.n38 B 0.601735f
C176 VP.n39 B 0.032801f
C177 VP.n40 B 0.053054f
C178 VP.n41 B 0.026694f
C179 VP.n42 B 0.026694f
C180 VP.n43 B 0.026694f
C181 VP.n44 B 0.053054f
C182 VP.n45 B 0.032801f
C183 VP.n46 B 0.601735f
C184 VP.n47 B 0.042135f
C185 VP.n48 B 0.026694f
C186 VP.n49 B 0.026694f
C187 VP.n50 B 0.026694f
C188 VP.n51 B 0.034505f
C189 VP.n52 B 0.04803f
C190 VP.n53 B 0.687623f
C191 VP.n54 B 0.029893f
.ends

