* NGSPICE file created from diff_pair_sample_1072.ext - technology: sky130A

.subckt diff_pair_sample_1072 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=0 ps=0 w=5.45 l=0.88
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=2.1255 ps=11.68 w=5.45 l=0.88
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=2.1255 ps=11.68 w=5.45 l=0.88
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=0 ps=0 w=5.45 l=0.88
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=0 ps=0 w=5.45 l=0.88
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=0 ps=0 w=5.45 l=0.88
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=2.1255 ps=11.68 w=5.45 l=0.88
X7 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1255 pd=11.68 as=2.1255 ps=11.68 w=5.45 l=0.88
R0 B.n400 B.n399 585
R1 B.n166 B.n58 585
R2 B.n165 B.n164 585
R3 B.n163 B.n162 585
R4 B.n161 B.n160 585
R5 B.n159 B.n158 585
R6 B.n157 B.n156 585
R7 B.n155 B.n154 585
R8 B.n153 B.n152 585
R9 B.n151 B.n150 585
R10 B.n149 B.n148 585
R11 B.n147 B.n146 585
R12 B.n145 B.n144 585
R13 B.n143 B.n142 585
R14 B.n141 B.n140 585
R15 B.n139 B.n138 585
R16 B.n137 B.n136 585
R17 B.n135 B.n134 585
R18 B.n133 B.n132 585
R19 B.n131 B.n130 585
R20 B.n129 B.n128 585
R21 B.n127 B.n126 585
R22 B.n125 B.n124 585
R23 B.n123 B.n122 585
R24 B.n121 B.n120 585
R25 B.n119 B.n118 585
R26 B.n117 B.n116 585
R27 B.n115 B.n114 585
R28 B.n113 B.n112 585
R29 B.n111 B.n110 585
R30 B.n109 B.n108 585
R31 B.n107 B.n106 585
R32 B.n105 B.n104 585
R33 B.n103 B.n102 585
R34 B.n101 B.n100 585
R35 B.n99 B.n98 585
R36 B.n97 B.n96 585
R37 B.n95 B.n94 585
R38 B.n93 B.n92 585
R39 B.n91 B.n90 585
R40 B.n89 B.n88 585
R41 B.n87 B.n86 585
R42 B.n85 B.n84 585
R43 B.n83 B.n82 585
R44 B.n81 B.n80 585
R45 B.n79 B.n78 585
R46 B.n77 B.n76 585
R47 B.n75 B.n74 585
R48 B.n73 B.n72 585
R49 B.n71 B.n70 585
R50 B.n69 B.n68 585
R51 B.n67 B.n66 585
R52 B.n32 B.n31 585
R53 B.n405 B.n404 585
R54 B.n398 B.n59 585
R55 B.n59 B.n29 585
R56 B.n397 B.n28 585
R57 B.n409 B.n28 585
R58 B.n396 B.n27 585
R59 B.n410 B.n27 585
R60 B.n395 B.n26 585
R61 B.n411 B.n26 585
R62 B.n394 B.n393 585
R63 B.n393 B.n25 585
R64 B.n392 B.n21 585
R65 B.n417 B.n21 585
R66 B.n391 B.n20 585
R67 B.n418 B.n20 585
R68 B.n390 B.n19 585
R69 B.n419 B.n19 585
R70 B.n389 B.n388 585
R71 B.n388 B.n15 585
R72 B.n387 B.n14 585
R73 B.n425 B.n14 585
R74 B.n386 B.n13 585
R75 B.n426 B.n13 585
R76 B.n385 B.n12 585
R77 B.n427 B.n12 585
R78 B.n384 B.n383 585
R79 B.n383 B.n8 585
R80 B.n382 B.n7 585
R81 B.n433 B.n7 585
R82 B.n381 B.n6 585
R83 B.n434 B.n6 585
R84 B.n380 B.n5 585
R85 B.n435 B.n5 585
R86 B.n379 B.n378 585
R87 B.n378 B.n4 585
R88 B.n377 B.n167 585
R89 B.n377 B.n376 585
R90 B.n367 B.n168 585
R91 B.n169 B.n168 585
R92 B.n369 B.n368 585
R93 B.n370 B.n369 585
R94 B.n366 B.n174 585
R95 B.n174 B.n173 585
R96 B.n365 B.n364 585
R97 B.n364 B.n363 585
R98 B.n176 B.n175 585
R99 B.n177 B.n176 585
R100 B.n356 B.n355 585
R101 B.n357 B.n356 585
R102 B.n354 B.n182 585
R103 B.n182 B.n181 585
R104 B.n353 B.n352 585
R105 B.n352 B.n351 585
R106 B.n184 B.n183 585
R107 B.n344 B.n184 585
R108 B.n343 B.n342 585
R109 B.n345 B.n343 585
R110 B.n341 B.n189 585
R111 B.n189 B.n188 585
R112 B.n340 B.n339 585
R113 B.n339 B.n338 585
R114 B.n191 B.n190 585
R115 B.n192 B.n191 585
R116 B.n334 B.n333 585
R117 B.n195 B.n194 585
R118 B.n330 B.n329 585
R119 B.n331 B.n330 585
R120 B.n328 B.n222 585
R121 B.n327 B.n326 585
R122 B.n325 B.n324 585
R123 B.n323 B.n322 585
R124 B.n321 B.n320 585
R125 B.n319 B.n318 585
R126 B.n317 B.n316 585
R127 B.n315 B.n314 585
R128 B.n313 B.n312 585
R129 B.n311 B.n310 585
R130 B.n309 B.n308 585
R131 B.n307 B.n306 585
R132 B.n305 B.n304 585
R133 B.n303 B.n302 585
R134 B.n301 B.n300 585
R135 B.n299 B.n298 585
R136 B.n297 B.n296 585
R137 B.n295 B.n294 585
R138 B.n293 B.n292 585
R139 B.n290 B.n289 585
R140 B.n288 B.n287 585
R141 B.n286 B.n285 585
R142 B.n284 B.n283 585
R143 B.n282 B.n281 585
R144 B.n280 B.n279 585
R145 B.n278 B.n277 585
R146 B.n276 B.n275 585
R147 B.n274 B.n273 585
R148 B.n272 B.n271 585
R149 B.n269 B.n268 585
R150 B.n267 B.n266 585
R151 B.n265 B.n264 585
R152 B.n263 B.n262 585
R153 B.n261 B.n260 585
R154 B.n259 B.n258 585
R155 B.n257 B.n256 585
R156 B.n255 B.n254 585
R157 B.n253 B.n252 585
R158 B.n251 B.n250 585
R159 B.n249 B.n248 585
R160 B.n247 B.n246 585
R161 B.n245 B.n244 585
R162 B.n243 B.n242 585
R163 B.n241 B.n240 585
R164 B.n239 B.n238 585
R165 B.n237 B.n236 585
R166 B.n235 B.n234 585
R167 B.n233 B.n232 585
R168 B.n231 B.n230 585
R169 B.n229 B.n228 585
R170 B.n227 B.n221 585
R171 B.n331 B.n221 585
R172 B.n335 B.n193 585
R173 B.n193 B.n192 585
R174 B.n337 B.n336 585
R175 B.n338 B.n337 585
R176 B.n187 B.n186 585
R177 B.n188 B.n187 585
R178 B.n347 B.n346 585
R179 B.n346 B.n345 585
R180 B.n348 B.n185 585
R181 B.n344 B.n185 585
R182 B.n350 B.n349 585
R183 B.n351 B.n350 585
R184 B.n180 B.n179 585
R185 B.n181 B.n180 585
R186 B.n359 B.n358 585
R187 B.n358 B.n357 585
R188 B.n360 B.n178 585
R189 B.n178 B.n177 585
R190 B.n362 B.n361 585
R191 B.n363 B.n362 585
R192 B.n172 B.n171 585
R193 B.n173 B.n172 585
R194 B.n372 B.n371 585
R195 B.n371 B.n370 585
R196 B.n373 B.n170 585
R197 B.n170 B.n169 585
R198 B.n375 B.n374 585
R199 B.n376 B.n375 585
R200 B.n2 B.n0 585
R201 B.n4 B.n2 585
R202 B.n3 B.n1 585
R203 B.n434 B.n3 585
R204 B.n432 B.n431 585
R205 B.n433 B.n432 585
R206 B.n430 B.n9 585
R207 B.n9 B.n8 585
R208 B.n429 B.n428 585
R209 B.n428 B.n427 585
R210 B.n11 B.n10 585
R211 B.n426 B.n11 585
R212 B.n424 B.n423 585
R213 B.n425 B.n424 585
R214 B.n422 B.n16 585
R215 B.n16 B.n15 585
R216 B.n421 B.n420 585
R217 B.n420 B.n419 585
R218 B.n18 B.n17 585
R219 B.n418 B.n18 585
R220 B.n416 B.n415 585
R221 B.n417 B.n416 585
R222 B.n414 B.n22 585
R223 B.n25 B.n22 585
R224 B.n413 B.n412 585
R225 B.n412 B.n411 585
R226 B.n24 B.n23 585
R227 B.n410 B.n24 585
R228 B.n408 B.n407 585
R229 B.n409 B.n408 585
R230 B.n406 B.n30 585
R231 B.n30 B.n29 585
R232 B.n437 B.n436 585
R233 B.n436 B.n435 585
R234 B.n333 B.n193 569.379
R235 B.n404 B.n30 569.379
R236 B.n221 B.n191 569.379
R237 B.n400 B.n59 569.379
R238 B.n225 B.t10 351.291
R239 B.n223 B.t2 351.291
R240 B.n63 B.t6 351.291
R241 B.n60 B.t13 351.291
R242 B.n402 B.n401 256.663
R243 B.n402 B.n57 256.663
R244 B.n402 B.n56 256.663
R245 B.n402 B.n55 256.663
R246 B.n402 B.n54 256.663
R247 B.n402 B.n53 256.663
R248 B.n402 B.n52 256.663
R249 B.n402 B.n51 256.663
R250 B.n402 B.n50 256.663
R251 B.n402 B.n49 256.663
R252 B.n402 B.n48 256.663
R253 B.n402 B.n47 256.663
R254 B.n402 B.n46 256.663
R255 B.n402 B.n45 256.663
R256 B.n402 B.n44 256.663
R257 B.n402 B.n43 256.663
R258 B.n402 B.n42 256.663
R259 B.n402 B.n41 256.663
R260 B.n402 B.n40 256.663
R261 B.n402 B.n39 256.663
R262 B.n402 B.n38 256.663
R263 B.n402 B.n37 256.663
R264 B.n402 B.n36 256.663
R265 B.n402 B.n35 256.663
R266 B.n402 B.n34 256.663
R267 B.n402 B.n33 256.663
R268 B.n403 B.n402 256.663
R269 B.n332 B.n331 256.663
R270 B.n331 B.n196 256.663
R271 B.n331 B.n197 256.663
R272 B.n331 B.n198 256.663
R273 B.n331 B.n199 256.663
R274 B.n331 B.n200 256.663
R275 B.n331 B.n201 256.663
R276 B.n331 B.n202 256.663
R277 B.n331 B.n203 256.663
R278 B.n331 B.n204 256.663
R279 B.n331 B.n205 256.663
R280 B.n331 B.n206 256.663
R281 B.n331 B.n207 256.663
R282 B.n331 B.n208 256.663
R283 B.n331 B.n209 256.663
R284 B.n331 B.n210 256.663
R285 B.n331 B.n211 256.663
R286 B.n331 B.n212 256.663
R287 B.n331 B.n213 256.663
R288 B.n331 B.n214 256.663
R289 B.n331 B.n215 256.663
R290 B.n331 B.n216 256.663
R291 B.n331 B.n217 256.663
R292 B.n331 B.n218 256.663
R293 B.n331 B.n219 256.663
R294 B.n331 B.n220 256.663
R295 B.n337 B.n193 163.367
R296 B.n337 B.n187 163.367
R297 B.n346 B.n187 163.367
R298 B.n346 B.n185 163.367
R299 B.n350 B.n185 163.367
R300 B.n350 B.n180 163.367
R301 B.n358 B.n180 163.367
R302 B.n358 B.n178 163.367
R303 B.n362 B.n178 163.367
R304 B.n362 B.n172 163.367
R305 B.n371 B.n172 163.367
R306 B.n371 B.n170 163.367
R307 B.n375 B.n170 163.367
R308 B.n375 B.n2 163.367
R309 B.n436 B.n2 163.367
R310 B.n436 B.n3 163.367
R311 B.n432 B.n3 163.367
R312 B.n432 B.n9 163.367
R313 B.n428 B.n9 163.367
R314 B.n428 B.n11 163.367
R315 B.n424 B.n11 163.367
R316 B.n424 B.n16 163.367
R317 B.n420 B.n16 163.367
R318 B.n420 B.n18 163.367
R319 B.n416 B.n18 163.367
R320 B.n416 B.n22 163.367
R321 B.n412 B.n22 163.367
R322 B.n412 B.n24 163.367
R323 B.n408 B.n24 163.367
R324 B.n408 B.n30 163.367
R325 B.n330 B.n195 163.367
R326 B.n330 B.n222 163.367
R327 B.n326 B.n325 163.367
R328 B.n322 B.n321 163.367
R329 B.n318 B.n317 163.367
R330 B.n314 B.n313 163.367
R331 B.n310 B.n309 163.367
R332 B.n306 B.n305 163.367
R333 B.n302 B.n301 163.367
R334 B.n298 B.n297 163.367
R335 B.n294 B.n293 163.367
R336 B.n289 B.n288 163.367
R337 B.n285 B.n284 163.367
R338 B.n281 B.n280 163.367
R339 B.n277 B.n276 163.367
R340 B.n273 B.n272 163.367
R341 B.n268 B.n267 163.367
R342 B.n264 B.n263 163.367
R343 B.n260 B.n259 163.367
R344 B.n256 B.n255 163.367
R345 B.n252 B.n251 163.367
R346 B.n248 B.n247 163.367
R347 B.n244 B.n243 163.367
R348 B.n240 B.n239 163.367
R349 B.n236 B.n235 163.367
R350 B.n232 B.n231 163.367
R351 B.n228 B.n221 163.367
R352 B.n339 B.n191 163.367
R353 B.n339 B.n189 163.367
R354 B.n343 B.n189 163.367
R355 B.n343 B.n184 163.367
R356 B.n352 B.n184 163.367
R357 B.n352 B.n182 163.367
R358 B.n356 B.n182 163.367
R359 B.n356 B.n176 163.367
R360 B.n364 B.n176 163.367
R361 B.n364 B.n174 163.367
R362 B.n369 B.n174 163.367
R363 B.n369 B.n168 163.367
R364 B.n377 B.n168 163.367
R365 B.n378 B.n377 163.367
R366 B.n378 B.n5 163.367
R367 B.n6 B.n5 163.367
R368 B.n7 B.n6 163.367
R369 B.n383 B.n7 163.367
R370 B.n383 B.n12 163.367
R371 B.n13 B.n12 163.367
R372 B.n14 B.n13 163.367
R373 B.n388 B.n14 163.367
R374 B.n388 B.n19 163.367
R375 B.n20 B.n19 163.367
R376 B.n21 B.n20 163.367
R377 B.n393 B.n21 163.367
R378 B.n393 B.n26 163.367
R379 B.n27 B.n26 163.367
R380 B.n28 B.n27 163.367
R381 B.n59 B.n28 163.367
R382 B.n66 B.n32 163.367
R383 B.n70 B.n69 163.367
R384 B.n74 B.n73 163.367
R385 B.n78 B.n77 163.367
R386 B.n82 B.n81 163.367
R387 B.n86 B.n85 163.367
R388 B.n90 B.n89 163.367
R389 B.n94 B.n93 163.367
R390 B.n98 B.n97 163.367
R391 B.n102 B.n101 163.367
R392 B.n106 B.n105 163.367
R393 B.n110 B.n109 163.367
R394 B.n114 B.n113 163.367
R395 B.n118 B.n117 163.367
R396 B.n122 B.n121 163.367
R397 B.n126 B.n125 163.367
R398 B.n130 B.n129 163.367
R399 B.n134 B.n133 163.367
R400 B.n138 B.n137 163.367
R401 B.n142 B.n141 163.367
R402 B.n146 B.n145 163.367
R403 B.n150 B.n149 163.367
R404 B.n154 B.n153 163.367
R405 B.n158 B.n157 163.367
R406 B.n162 B.n161 163.367
R407 B.n164 B.n58 163.367
R408 B.n331 B.n192 142.299
R409 B.n402 B.n29 142.299
R410 B.n225 B.t12 93.458
R411 B.n60 B.t14 93.458
R412 B.n223 B.t5 93.4522
R413 B.n63 B.t8 93.4522
R414 B.n333 B.n332 71.676
R415 B.n222 B.n196 71.676
R416 B.n325 B.n197 71.676
R417 B.n321 B.n198 71.676
R418 B.n317 B.n199 71.676
R419 B.n313 B.n200 71.676
R420 B.n309 B.n201 71.676
R421 B.n305 B.n202 71.676
R422 B.n301 B.n203 71.676
R423 B.n297 B.n204 71.676
R424 B.n293 B.n205 71.676
R425 B.n288 B.n206 71.676
R426 B.n284 B.n207 71.676
R427 B.n280 B.n208 71.676
R428 B.n276 B.n209 71.676
R429 B.n272 B.n210 71.676
R430 B.n267 B.n211 71.676
R431 B.n263 B.n212 71.676
R432 B.n259 B.n213 71.676
R433 B.n255 B.n214 71.676
R434 B.n251 B.n215 71.676
R435 B.n247 B.n216 71.676
R436 B.n243 B.n217 71.676
R437 B.n239 B.n218 71.676
R438 B.n235 B.n219 71.676
R439 B.n231 B.n220 71.676
R440 B.n404 B.n403 71.676
R441 B.n66 B.n33 71.676
R442 B.n70 B.n34 71.676
R443 B.n74 B.n35 71.676
R444 B.n78 B.n36 71.676
R445 B.n82 B.n37 71.676
R446 B.n86 B.n38 71.676
R447 B.n90 B.n39 71.676
R448 B.n94 B.n40 71.676
R449 B.n98 B.n41 71.676
R450 B.n102 B.n42 71.676
R451 B.n106 B.n43 71.676
R452 B.n110 B.n44 71.676
R453 B.n114 B.n45 71.676
R454 B.n118 B.n46 71.676
R455 B.n122 B.n47 71.676
R456 B.n126 B.n48 71.676
R457 B.n130 B.n49 71.676
R458 B.n134 B.n50 71.676
R459 B.n138 B.n51 71.676
R460 B.n142 B.n52 71.676
R461 B.n146 B.n53 71.676
R462 B.n150 B.n54 71.676
R463 B.n154 B.n55 71.676
R464 B.n158 B.n56 71.676
R465 B.n162 B.n57 71.676
R466 B.n401 B.n58 71.676
R467 B.n401 B.n400 71.676
R468 B.n164 B.n57 71.676
R469 B.n161 B.n56 71.676
R470 B.n157 B.n55 71.676
R471 B.n153 B.n54 71.676
R472 B.n149 B.n53 71.676
R473 B.n145 B.n52 71.676
R474 B.n141 B.n51 71.676
R475 B.n137 B.n50 71.676
R476 B.n133 B.n49 71.676
R477 B.n129 B.n48 71.676
R478 B.n125 B.n47 71.676
R479 B.n121 B.n46 71.676
R480 B.n117 B.n45 71.676
R481 B.n113 B.n44 71.676
R482 B.n109 B.n43 71.676
R483 B.n105 B.n42 71.676
R484 B.n101 B.n41 71.676
R485 B.n97 B.n40 71.676
R486 B.n93 B.n39 71.676
R487 B.n89 B.n38 71.676
R488 B.n85 B.n37 71.676
R489 B.n81 B.n36 71.676
R490 B.n77 B.n35 71.676
R491 B.n73 B.n34 71.676
R492 B.n69 B.n33 71.676
R493 B.n403 B.n32 71.676
R494 B.n332 B.n195 71.676
R495 B.n326 B.n196 71.676
R496 B.n322 B.n197 71.676
R497 B.n318 B.n198 71.676
R498 B.n314 B.n199 71.676
R499 B.n310 B.n200 71.676
R500 B.n306 B.n201 71.676
R501 B.n302 B.n202 71.676
R502 B.n298 B.n203 71.676
R503 B.n294 B.n204 71.676
R504 B.n289 B.n205 71.676
R505 B.n285 B.n206 71.676
R506 B.n281 B.n207 71.676
R507 B.n277 B.n208 71.676
R508 B.n273 B.n209 71.676
R509 B.n268 B.n210 71.676
R510 B.n264 B.n211 71.676
R511 B.n260 B.n212 71.676
R512 B.n256 B.n213 71.676
R513 B.n252 B.n214 71.676
R514 B.n248 B.n215 71.676
R515 B.n244 B.n216 71.676
R516 B.n240 B.n217 71.676
R517 B.n236 B.n218 71.676
R518 B.n232 B.n219 71.676
R519 B.n228 B.n220 71.676
R520 B.n226 B.t11 69.9913
R521 B.n61 B.t15 69.9913
R522 B.n224 B.t4 69.9855
R523 B.n64 B.t9 69.9855
R524 B.n338 B.n192 69.6143
R525 B.n338 B.n188 69.6143
R526 B.n345 B.n188 69.6143
R527 B.n345 B.n344 69.6143
R528 B.n351 B.n181 69.6143
R529 B.n357 B.n181 69.6143
R530 B.n357 B.n177 69.6143
R531 B.n363 B.n177 69.6143
R532 B.n363 B.n173 69.6143
R533 B.n370 B.n173 69.6143
R534 B.n376 B.n169 69.6143
R535 B.n376 B.n4 69.6143
R536 B.n435 B.n4 69.6143
R537 B.n435 B.n434 69.6143
R538 B.n434 B.n433 69.6143
R539 B.n433 B.n8 69.6143
R540 B.n427 B.n426 69.6143
R541 B.n426 B.n425 69.6143
R542 B.n425 B.n15 69.6143
R543 B.n419 B.n15 69.6143
R544 B.n419 B.n418 69.6143
R545 B.n418 B.n417 69.6143
R546 B.n411 B.n25 69.6143
R547 B.n411 B.n410 69.6143
R548 B.n410 B.n409 69.6143
R549 B.n409 B.n29 69.6143
R550 B.n270 B.n226 59.5399
R551 B.n291 B.n224 59.5399
R552 B.n65 B.n64 59.5399
R553 B.n62 B.n61 59.5399
R554 B.n344 B.t3 59.377
R555 B.n25 B.t7 59.377
R556 B.n370 B.t0 42.9972
R557 B.n427 B.t1 42.9972
R558 B.n406 B.n405 36.9956
R559 B.n399 B.n398 36.9956
R560 B.n227 B.n190 36.9956
R561 B.n335 B.n334 36.9956
R562 B.t0 B.n169 26.6175
R563 B.t1 B.n8 26.6175
R564 B.n226 B.n225 23.4672
R565 B.n224 B.n223 23.4672
R566 B.n64 B.n63 23.4672
R567 B.n61 B.n60 23.4672
R568 B B.n437 18.0485
R569 B.n405 B.n31 10.6151
R570 B.n67 B.n31 10.6151
R571 B.n68 B.n67 10.6151
R572 B.n71 B.n68 10.6151
R573 B.n72 B.n71 10.6151
R574 B.n75 B.n72 10.6151
R575 B.n76 B.n75 10.6151
R576 B.n79 B.n76 10.6151
R577 B.n80 B.n79 10.6151
R578 B.n83 B.n80 10.6151
R579 B.n84 B.n83 10.6151
R580 B.n87 B.n84 10.6151
R581 B.n88 B.n87 10.6151
R582 B.n91 B.n88 10.6151
R583 B.n92 B.n91 10.6151
R584 B.n95 B.n92 10.6151
R585 B.n96 B.n95 10.6151
R586 B.n99 B.n96 10.6151
R587 B.n100 B.n99 10.6151
R588 B.n103 B.n100 10.6151
R589 B.n104 B.n103 10.6151
R590 B.n108 B.n107 10.6151
R591 B.n111 B.n108 10.6151
R592 B.n112 B.n111 10.6151
R593 B.n115 B.n112 10.6151
R594 B.n116 B.n115 10.6151
R595 B.n119 B.n116 10.6151
R596 B.n120 B.n119 10.6151
R597 B.n123 B.n120 10.6151
R598 B.n124 B.n123 10.6151
R599 B.n128 B.n127 10.6151
R600 B.n131 B.n128 10.6151
R601 B.n132 B.n131 10.6151
R602 B.n135 B.n132 10.6151
R603 B.n136 B.n135 10.6151
R604 B.n139 B.n136 10.6151
R605 B.n140 B.n139 10.6151
R606 B.n143 B.n140 10.6151
R607 B.n144 B.n143 10.6151
R608 B.n147 B.n144 10.6151
R609 B.n148 B.n147 10.6151
R610 B.n151 B.n148 10.6151
R611 B.n152 B.n151 10.6151
R612 B.n155 B.n152 10.6151
R613 B.n156 B.n155 10.6151
R614 B.n159 B.n156 10.6151
R615 B.n160 B.n159 10.6151
R616 B.n163 B.n160 10.6151
R617 B.n165 B.n163 10.6151
R618 B.n166 B.n165 10.6151
R619 B.n399 B.n166 10.6151
R620 B.n340 B.n190 10.6151
R621 B.n341 B.n340 10.6151
R622 B.n342 B.n341 10.6151
R623 B.n342 B.n183 10.6151
R624 B.n353 B.n183 10.6151
R625 B.n354 B.n353 10.6151
R626 B.n355 B.n354 10.6151
R627 B.n355 B.n175 10.6151
R628 B.n365 B.n175 10.6151
R629 B.n366 B.n365 10.6151
R630 B.n368 B.n366 10.6151
R631 B.n368 B.n367 10.6151
R632 B.n367 B.n167 10.6151
R633 B.n379 B.n167 10.6151
R634 B.n380 B.n379 10.6151
R635 B.n381 B.n380 10.6151
R636 B.n382 B.n381 10.6151
R637 B.n384 B.n382 10.6151
R638 B.n385 B.n384 10.6151
R639 B.n386 B.n385 10.6151
R640 B.n387 B.n386 10.6151
R641 B.n389 B.n387 10.6151
R642 B.n390 B.n389 10.6151
R643 B.n391 B.n390 10.6151
R644 B.n392 B.n391 10.6151
R645 B.n394 B.n392 10.6151
R646 B.n395 B.n394 10.6151
R647 B.n396 B.n395 10.6151
R648 B.n397 B.n396 10.6151
R649 B.n398 B.n397 10.6151
R650 B.n334 B.n194 10.6151
R651 B.n329 B.n194 10.6151
R652 B.n329 B.n328 10.6151
R653 B.n328 B.n327 10.6151
R654 B.n327 B.n324 10.6151
R655 B.n324 B.n323 10.6151
R656 B.n323 B.n320 10.6151
R657 B.n320 B.n319 10.6151
R658 B.n319 B.n316 10.6151
R659 B.n316 B.n315 10.6151
R660 B.n315 B.n312 10.6151
R661 B.n312 B.n311 10.6151
R662 B.n311 B.n308 10.6151
R663 B.n308 B.n307 10.6151
R664 B.n307 B.n304 10.6151
R665 B.n304 B.n303 10.6151
R666 B.n303 B.n300 10.6151
R667 B.n300 B.n299 10.6151
R668 B.n299 B.n296 10.6151
R669 B.n296 B.n295 10.6151
R670 B.n295 B.n292 10.6151
R671 B.n290 B.n287 10.6151
R672 B.n287 B.n286 10.6151
R673 B.n286 B.n283 10.6151
R674 B.n283 B.n282 10.6151
R675 B.n282 B.n279 10.6151
R676 B.n279 B.n278 10.6151
R677 B.n278 B.n275 10.6151
R678 B.n275 B.n274 10.6151
R679 B.n274 B.n271 10.6151
R680 B.n269 B.n266 10.6151
R681 B.n266 B.n265 10.6151
R682 B.n265 B.n262 10.6151
R683 B.n262 B.n261 10.6151
R684 B.n261 B.n258 10.6151
R685 B.n258 B.n257 10.6151
R686 B.n257 B.n254 10.6151
R687 B.n254 B.n253 10.6151
R688 B.n253 B.n250 10.6151
R689 B.n250 B.n249 10.6151
R690 B.n249 B.n246 10.6151
R691 B.n246 B.n245 10.6151
R692 B.n245 B.n242 10.6151
R693 B.n242 B.n241 10.6151
R694 B.n241 B.n238 10.6151
R695 B.n238 B.n237 10.6151
R696 B.n237 B.n234 10.6151
R697 B.n234 B.n233 10.6151
R698 B.n233 B.n230 10.6151
R699 B.n230 B.n229 10.6151
R700 B.n229 B.n227 10.6151
R701 B.n336 B.n335 10.6151
R702 B.n336 B.n186 10.6151
R703 B.n347 B.n186 10.6151
R704 B.n348 B.n347 10.6151
R705 B.n349 B.n348 10.6151
R706 B.n349 B.n179 10.6151
R707 B.n359 B.n179 10.6151
R708 B.n360 B.n359 10.6151
R709 B.n361 B.n360 10.6151
R710 B.n361 B.n171 10.6151
R711 B.n372 B.n171 10.6151
R712 B.n373 B.n372 10.6151
R713 B.n374 B.n373 10.6151
R714 B.n374 B.n0 10.6151
R715 B.n431 B.n1 10.6151
R716 B.n431 B.n430 10.6151
R717 B.n430 B.n429 10.6151
R718 B.n429 B.n10 10.6151
R719 B.n423 B.n10 10.6151
R720 B.n423 B.n422 10.6151
R721 B.n422 B.n421 10.6151
R722 B.n421 B.n17 10.6151
R723 B.n415 B.n17 10.6151
R724 B.n415 B.n414 10.6151
R725 B.n414 B.n413 10.6151
R726 B.n413 B.n23 10.6151
R727 B.n407 B.n23 10.6151
R728 B.n407 B.n406 10.6151
R729 B.n351 B.t3 10.2378
R730 B.n417 B.t7 10.2378
R731 B.n104 B.n65 8.74196
R732 B.n127 B.n62 8.74196
R733 B.n292 B.n291 8.74196
R734 B.n270 B.n269 8.74196
R735 B.n437 B.n0 2.81026
R736 B.n437 B.n1 2.81026
R737 B.n107 B.n65 1.87367
R738 B.n124 B.n62 1.87367
R739 B.n291 B.n290 1.87367
R740 B.n271 B.n270 1.87367
R741 VN VN.t0 390.998
R742 VN VN.t1 355.521
R743 VTAIL.n1 VTAIL.t3 57.218
R744 VTAIL.n2 VTAIL.t1 57.217
R745 VTAIL.n3 VTAIL.t2 57.217
R746 VTAIL.n0 VTAIL.t0 57.217
R747 VTAIL.n1 VTAIL.n0 19.1686
R748 VTAIL.n3 VTAIL.n2 18.1255
R749 VTAIL.n2 VTAIL.n1 0.991879
R750 VTAIL VTAIL.n0 0.789293
R751 VTAIL VTAIL.n3 0.203086
R752 VDD2.n0 VDD2.t0 104.356
R753 VDD2.n0 VDD2.t1 73.8958
R754 VDD2 VDD2.n0 0.319466
R755 VP.n0 VP.t0 390.618
R756 VP.n0 VP.t1 355.469
R757 VP VP.n0 0.0516364
R758 VDD1 VDD1.t0 105.142
R759 VDD1 VDD1.t1 74.2148
C0 VP VDD2 0.265356f
C1 VP VTAIL 0.977688f
C2 VTAIL VDD2 3.20246f
C3 VN VDD1 0.148671f
C4 VP VDD1 1.21781f
C5 VN VP 3.4301f
C6 VDD1 VDD2 0.47819f
C7 VN VDD2 1.10689f
C8 VTAIL VDD1 3.16345f
C9 VN VTAIL 0.963379f
C10 VDD2 B 2.618494f
C11 VDD1 B 4.29981f
C12 VTAIL B 3.839462f
C13 VN B 6.01156f
C14 VP B 3.731956f
C15 VDD1.t1 B 0.697776f
C16 VDD1.t0 B 0.919657f
C17 VP.t0 B 0.661624f
C18 VP.t1 B 0.560652f
C19 VP.n0 B 2.16246f
C20 VDD2.t0 B 0.920684f
C21 VDD2.t1 B 0.70958f
C22 VDD2.n0 B 1.52709f
C23 VTAIL.t0 B 0.75218f
C24 VTAIL.n0 B 0.865906f
C25 VTAIL.t3 B 0.75218f
C26 VTAIL.n1 B 0.877393f
C27 VTAIL.t1 B 0.752177f
C28 VTAIL.n2 B 0.818251f
C29 VTAIL.t2 B 0.75218f
C30 VTAIL.n3 B 0.773522f
C31 VN.t1 B 0.553073f
C32 VN.t0 B 0.655615f
.ends

