* NGSPICE file created from diff_pair_sample_0604.ext - technology: sky130A

.subckt diff_pair_sample_0604 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t16 VN.t0 VDD2.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X1 VDD1.t9 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X2 VTAIL.t15 VN.t1 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X3 VDD1.t8 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=2.98485 ps=18.42 w=18.09 l=2.46
X4 VDD2.t0 VN.t2 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X5 VTAIL.t1 VP.t2 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X6 VDD2.t3 VN.t3 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=2.98485 ps=18.42 w=18.09 l=2.46
X7 VDD2.t2 VN.t4 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X8 VDD1.t6 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=7.0551 ps=36.96 w=18.09 l=2.46
X9 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=0 ps=0 w=18.09 l=2.46
X10 VDD2.t7 VN.t5 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=2.98485 ps=18.42 w=18.09 l=2.46
X11 VTAIL.t10 VN.t6 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X12 VDD1.t5 VP.t4 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X13 VTAIL.t3 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X14 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=0 ps=0 w=18.09 l=2.46
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=0 ps=0 w=18.09 l=2.46
X16 VDD1.t3 VP.t6 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=2.98485 ps=18.42 w=18.09 l=2.46
X17 VDD2.t9 VN.t7 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=7.0551 ps=36.96 w=18.09 l=2.46
X18 VTAIL.t19 VP.t7 VDD1.t2 B.t9 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X19 VDD2.t8 VN.t8 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=7.0551 ps=36.96 w=18.09 l=2.46
X20 VDD1.t1 VP.t8 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=7.0551 ps=36.96 w=18.09 l=2.46
X21 VTAIL.t6 VP.t9 VDD1.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X22 VTAIL.t7 VN.t9 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.98485 pd=18.42 as=2.98485 ps=18.42 w=18.09 l=2.46
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.0551 pd=36.96 as=0 ps=0 w=18.09 l=2.46
R0 VN.n10 VN.t3 208.897
R1 VN.n49 VN.t7 208.897
R2 VN.n19 VN.t2 177.224
R3 VN.n9 VN.t9 177.224
R4 VN.n3 VN.t0 177.224
R5 VN.n37 VN.t8 177.224
R6 VN.n58 VN.t4 177.224
R7 VN.n48 VN.t6 177.224
R8 VN.n42 VN.t1 177.224
R9 VN.n76 VN.t5 177.224
R10 VN.n75 VN.n39 161.3
R11 VN.n74 VN.n73 161.3
R12 VN.n72 VN.n40 161.3
R13 VN.n71 VN.n70 161.3
R14 VN.n69 VN.n41 161.3
R15 VN.n68 VN.n67 161.3
R16 VN.n66 VN.n65 161.3
R17 VN.n64 VN.n43 161.3
R18 VN.n63 VN.n62 161.3
R19 VN.n61 VN.n44 161.3
R20 VN.n60 VN.n59 161.3
R21 VN.n58 VN.n45 161.3
R22 VN.n57 VN.n56 161.3
R23 VN.n55 VN.n46 161.3
R24 VN.n54 VN.n53 161.3
R25 VN.n52 VN.n47 161.3
R26 VN.n51 VN.n50 161.3
R27 VN.n36 VN.n0 161.3
R28 VN.n35 VN.n34 161.3
R29 VN.n33 VN.n1 161.3
R30 VN.n32 VN.n31 161.3
R31 VN.n30 VN.n2 161.3
R32 VN.n29 VN.n28 161.3
R33 VN.n27 VN.n26 161.3
R34 VN.n25 VN.n4 161.3
R35 VN.n24 VN.n23 161.3
R36 VN.n22 VN.n5 161.3
R37 VN.n21 VN.n20 161.3
R38 VN.n19 VN.n6 161.3
R39 VN.n18 VN.n17 161.3
R40 VN.n16 VN.n7 161.3
R41 VN.n15 VN.n14 161.3
R42 VN.n13 VN.n8 161.3
R43 VN.n12 VN.n11 161.3
R44 VN.n38 VN.n37 106.841
R45 VN.n77 VN.n76 106.841
R46 VN.n10 VN.n9 57.8794
R47 VN.n49 VN.n48 57.8794
R48 VN VN.n77 57.1383
R49 VN.n31 VN.n1 56.5193
R50 VN.n70 VN.n40 56.5193
R51 VN.n14 VN.n7 50.6917
R52 VN.n24 VN.n5 50.6917
R53 VN.n53 VN.n46 50.6917
R54 VN.n63 VN.n44 50.6917
R55 VN.n14 VN.n13 30.2951
R56 VN.n25 VN.n24 30.2951
R57 VN.n53 VN.n52 30.2951
R58 VN.n64 VN.n63 30.2951
R59 VN.n13 VN.n12 24.4675
R60 VN.n18 VN.n7 24.4675
R61 VN.n19 VN.n18 24.4675
R62 VN.n20 VN.n19 24.4675
R63 VN.n20 VN.n5 24.4675
R64 VN.n26 VN.n25 24.4675
R65 VN.n30 VN.n29 24.4675
R66 VN.n31 VN.n30 24.4675
R67 VN.n35 VN.n1 24.4675
R68 VN.n36 VN.n35 24.4675
R69 VN.n52 VN.n51 24.4675
R70 VN.n59 VN.n44 24.4675
R71 VN.n59 VN.n58 24.4675
R72 VN.n58 VN.n57 24.4675
R73 VN.n57 VN.n46 24.4675
R74 VN.n70 VN.n69 24.4675
R75 VN.n69 VN.n68 24.4675
R76 VN.n65 VN.n64 24.4675
R77 VN.n75 VN.n74 24.4675
R78 VN.n74 VN.n40 24.4675
R79 VN.n12 VN.n9 14.1914
R80 VN.n26 VN.n3 14.1914
R81 VN.n51 VN.n48 14.1914
R82 VN.n65 VN.n42 14.1914
R83 VN.n29 VN.n3 10.2766
R84 VN.n68 VN.n42 10.2766
R85 VN.n50 VN.n49 7.2327
R86 VN.n11 VN.n10 7.2327
R87 VN.n37 VN.n36 3.91522
R88 VN.n76 VN.n75 3.91522
R89 VN.n77 VN.n39 0.278367
R90 VN.n38 VN.n0 0.278367
R91 VN.n73 VN.n39 0.189894
R92 VN.n73 VN.n72 0.189894
R93 VN.n72 VN.n71 0.189894
R94 VN.n71 VN.n41 0.189894
R95 VN.n67 VN.n41 0.189894
R96 VN.n67 VN.n66 0.189894
R97 VN.n66 VN.n43 0.189894
R98 VN.n62 VN.n43 0.189894
R99 VN.n62 VN.n61 0.189894
R100 VN.n61 VN.n60 0.189894
R101 VN.n60 VN.n45 0.189894
R102 VN.n56 VN.n45 0.189894
R103 VN.n56 VN.n55 0.189894
R104 VN.n55 VN.n54 0.189894
R105 VN.n54 VN.n47 0.189894
R106 VN.n50 VN.n47 0.189894
R107 VN.n11 VN.n8 0.189894
R108 VN.n15 VN.n8 0.189894
R109 VN.n16 VN.n15 0.189894
R110 VN.n17 VN.n16 0.189894
R111 VN.n17 VN.n6 0.189894
R112 VN.n21 VN.n6 0.189894
R113 VN.n22 VN.n21 0.189894
R114 VN.n23 VN.n22 0.189894
R115 VN.n23 VN.n4 0.189894
R116 VN.n27 VN.n4 0.189894
R117 VN.n28 VN.n27 0.189894
R118 VN.n28 VN.n2 0.189894
R119 VN.n32 VN.n2 0.189894
R120 VN.n33 VN.n32 0.189894
R121 VN.n34 VN.n33 0.189894
R122 VN.n34 VN.n0 0.189894
R123 VN VN.n38 0.153454
R124 VDD2.n201 VDD2.n200 289.615
R125 VDD2.n98 VDD2.n97 289.615
R126 VDD2.n200 VDD2.n199 185
R127 VDD2.n105 VDD2.n104 185
R128 VDD2.n194 VDD2.n193 185
R129 VDD2.n192 VDD2.n191 185
R130 VDD2.n109 VDD2.n108 185
R131 VDD2.n186 VDD2.n185 185
R132 VDD2.n184 VDD2.n183 185
R133 VDD2.n113 VDD2.n112 185
R134 VDD2.n178 VDD2.n177 185
R135 VDD2.n176 VDD2.n175 185
R136 VDD2.n117 VDD2.n116 185
R137 VDD2.n170 VDD2.n169 185
R138 VDD2.n168 VDD2.n167 185
R139 VDD2.n121 VDD2.n120 185
R140 VDD2.n162 VDD2.n161 185
R141 VDD2.n160 VDD2.n159 185
R142 VDD2.n158 VDD2.n124 185
R143 VDD2.n128 VDD2.n125 185
R144 VDD2.n153 VDD2.n152 185
R145 VDD2.n151 VDD2.n150 185
R146 VDD2.n130 VDD2.n129 185
R147 VDD2.n145 VDD2.n144 185
R148 VDD2.n143 VDD2.n142 185
R149 VDD2.n134 VDD2.n133 185
R150 VDD2.n137 VDD2.n136 185
R151 VDD2.n33 VDD2.n32 185
R152 VDD2.n30 VDD2.n29 185
R153 VDD2.n39 VDD2.n38 185
R154 VDD2.n41 VDD2.n40 185
R155 VDD2.n26 VDD2.n25 185
R156 VDD2.n47 VDD2.n46 185
R157 VDD2.n50 VDD2.n49 185
R158 VDD2.n48 VDD2.n22 185
R159 VDD2.n55 VDD2.n21 185
R160 VDD2.n57 VDD2.n56 185
R161 VDD2.n59 VDD2.n58 185
R162 VDD2.n18 VDD2.n17 185
R163 VDD2.n65 VDD2.n64 185
R164 VDD2.n67 VDD2.n66 185
R165 VDD2.n14 VDD2.n13 185
R166 VDD2.n73 VDD2.n72 185
R167 VDD2.n75 VDD2.n74 185
R168 VDD2.n10 VDD2.n9 185
R169 VDD2.n81 VDD2.n80 185
R170 VDD2.n83 VDD2.n82 185
R171 VDD2.n6 VDD2.n5 185
R172 VDD2.n89 VDD2.n88 185
R173 VDD2.n91 VDD2.n90 185
R174 VDD2.n2 VDD2.n1 185
R175 VDD2.n97 VDD2.n96 185
R176 VDD2.t7 VDD2.n135 149.524
R177 VDD2.t3 VDD2.n31 149.524
R178 VDD2.n200 VDD2.n104 104.615
R179 VDD2.n193 VDD2.n104 104.615
R180 VDD2.n193 VDD2.n192 104.615
R181 VDD2.n192 VDD2.n108 104.615
R182 VDD2.n185 VDD2.n108 104.615
R183 VDD2.n185 VDD2.n184 104.615
R184 VDD2.n184 VDD2.n112 104.615
R185 VDD2.n177 VDD2.n112 104.615
R186 VDD2.n177 VDD2.n176 104.615
R187 VDD2.n176 VDD2.n116 104.615
R188 VDD2.n169 VDD2.n116 104.615
R189 VDD2.n169 VDD2.n168 104.615
R190 VDD2.n168 VDD2.n120 104.615
R191 VDD2.n161 VDD2.n120 104.615
R192 VDD2.n161 VDD2.n160 104.615
R193 VDD2.n160 VDD2.n124 104.615
R194 VDD2.n128 VDD2.n124 104.615
R195 VDD2.n152 VDD2.n128 104.615
R196 VDD2.n152 VDD2.n151 104.615
R197 VDD2.n151 VDD2.n129 104.615
R198 VDD2.n144 VDD2.n129 104.615
R199 VDD2.n144 VDD2.n143 104.615
R200 VDD2.n143 VDD2.n133 104.615
R201 VDD2.n136 VDD2.n133 104.615
R202 VDD2.n32 VDD2.n29 104.615
R203 VDD2.n39 VDD2.n29 104.615
R204 VDD2.n40 VDD2.n39 104.615
R205 VDD2.n40 VDD2.n25 104.615
R206 VDD2.n47 VDD2.n25 104.615
R207 VDD2.n49 VDD2.n47 104.615
R208 VDD2.n49 VDD2.n48 104.615
R209 VDD2.n48 VDD2.n21 104.615
R210 VDD2.n57 VDD2.n21 104.615
R211 VDD2.n58 VDD2.n57 104.615
R212 VDD2.n58 VDD2.n17 104.615
R213 VDD2.n65 VDD2.n17 104.615
R214 VDD2.n66 VDD2.n65 104.615
R215 VDD2.n66 VDD2.n13 104.615
R216 VDD2.n73 VDD2.n13 104.615
R217 VDD2.n74 VDD2.n73 104.615
R218 VDD2.n74 VDD2.n9 104.615
R219 VDD2.n81 VDD2.n9 104.615
R220 VDD2.n82 VDD2.n81 104.615
R221 VDD2.n82 VDD2.n5 104.615
R222 VDD2.n89 VDD2.n5 104.615
R223 VDD2.n90 VDD2.n89 104.615
R224 VDD2.n90 VDD2.n1 104.615
R225 VDD2.n97 VDD2.n1 104.615
R226 VDD2.n102 VDD2.n101 65.928
R227 VDD2 VDD2.n205 65.9242
R228 VDD2.n204 VDD2.n203 64.1796
R229 VDD2.n100 VDD2.n99 64.1795
R230 VDD2.n100 VDD2.n98 54.1784
R231 VDD2.n136 VDD2.t7 52.3082
R232 VDD2.n32 VDD2.t3 52.3082
R233 VDD2.n202 VDD2.n201 51.7732
R234 VDD2.n202 VDD2.n102 50.7347
R235 VDD2.n159 VDD2.n158 13.1884
R236 VDD2.n56 VDD2.n55 13.1884
R237 VDD2.n162 VDD2.n123 12.8005
R238 VDD2.n157 VDD2.n125 12.8005
R239 VDD2.n54 VDD2.n22 12.8005
R240 VDD2.n59 VDD2.n20 12.8005
R241 VDD2.n199 VDD2.n103 12.0247
R242 VDD2.n163 VDD2.n121 12.0247
R243 VDD2.n154 VDD2.n153 12.0247
R244 VDD2.n51 VDD2.n50 12.0247
R245 VDD2.n60 VDD2.n18 12.0247
R246 VDD2.n96 VDD2.n0 12.0247
R247 VDD2.n198 VDD2.n105 11.249
R248 VDD2.n167 VDD2.n166 11.249
R249 VDD2.n150 VDD2.n127 11.249
R250 VDD2.n46 VDD2.n24 11.249
R251 VDD2.n64 VDD2.n63 11.249
R252 VDD2.n95 VDD2.n2 11.249
R253 VDD2.n195 VDD2.n194 10.4732
R254 VDD2.n170 VDD2.n119 10.4732
R255 VDD2.n149 VDD2.n130 10.4732
R256 VDD2.n45 VDD2.n26 10.4732
R257 VDD2.n67 VDD2.n16 10.4732
R258 VDD2.n92 VDD2.n91 10.4732
R259 VDD2.n137 VDD2.n135 10.2747
R260 VDD2.n33 VDD2.n31 10.2747
R261 VDD2.n191 VDD2.n107 9.69747
R262 VDD2.n171 VDD2.n117 9.69747
R263 VDD2.n146 VDD2.n145 9.69747
R264 VDD2.n42 VDD2.n41 9.69747
R265 VDD2.n68 VDD2.n14 9.69747
R266 VDD2.n88 VDD2.n4 9.69747
R267 VDD2.n197 VDD2.n103 9.45567
R268 VDD2.n94 VDD2.n0 9.45567
R269 VDD2.n139 VDD2.n138 9.3005
R270 VDD2.n141 VDD2.n140 9.3005
R271 VDD2.n132 VDD2.n131 9.3005
R272 VDD2.n147 VDD2.n146 9.3005
R273 VDD2.n149 VDD2.n148 9.3005
R274 VDD2.n127 VDD2.n126 9.3005
R275 VDD2.n155 VDD2.n154 9.3005
R276 VDD2.n157 VDD2.n156 9.3005
R277 VDD2.n111 VDD2.n110 9.3005
R278 VDD2.n188 VDD2.n187 9.3005
R279 VDD2.n190 VDD2.n189 9.3005
R280 VDD2.n107 VDD2.n106 9.3005
R281 VDD2.n196 VDD2.n195 9.3005
R282 VDD2.n198 VDD2.n197 9.3005
R283 VDD2.n182 VDD2.n181 9.3005
R284 VDD2.n180 VDD2.n179 9.3005
R285 VDD2.n115 VDD2.n114 9.3005
R286 VDD2.n174 VDD2.n173 9.3005
R287 VDD2.n172 VDD2.n171 9.3005
R288 VDD2.n119 VDD2.n118 9.3005
R289 VDD2.n166 VDD2.n165 9.3005
R290 VDD2.n164 VDD2.n163 9.3005
R291 VDD2.n123 VDD2.n122 9.3005
R292 VDD2.n79 VDD2.n78 9.3005
R293 VDD2.n8 VDD2.n7 9.3005
R294 VDD2.n85 VDD2.n84 9.3005
R295 VDD2.n87 VDD2.n86 9.3005
R296 VDD2.n4 VDD2.n3 9.3005
R297 VDD2.n93 VDD2.n92 9.3005
R298 VDD2.n95 VDD2.n94 9.3005
R299 VDD2.n12 VDD2.n11 9.3005
R300 VDD2.n71 VDD2.n70 9.3005
R301 VDD2.n69 VDD2.n68 9.3005
R302 VDD2.n16 VDD2.n15 9.3005
R303 VDD2.n63 VDD2.n62 9.3005
R304 VDD2.n61 VDD2.n60 9.3005
R305 VDD2.n20 VDD2.n19 9.3005
R306 VDD2.n35 VDD2.n34 9.3005
R307 VDD2.n37 VDD2.n36 9.3005
R308 VDD2.n28 VDD2.n27 9.3005
R309 VDD2.n43 VDD2.n42 9.3005
R310 VDD2.n45 VDD2.n44 9.3005
R311 VDD2.n24 VDD2.n23 9.3005
R312 VDD2.n52 VDD2.n51 9.3005
R313 VDD2.n54 VDD2.n53 9.3005
R314 VDD2.n77 VDD2.n76 9.3005
R315 VDD2.n190 VDD2.n109 8.92171
R316 VDD2.n175 VDD2.n174 8.92171
R317 VDD2.n142 VDD2.n132 8.92171
R318 VDD2.n38 VDD2.n28 8.92171
R319 VDD2.n72 VDD2.n71 8.92171
R320 VDD2.n87 VDD2.n6 8.92171
R321 VDD2.n187 VDD2.n186 8.14595
R322 VDD2.n178 VDD2.n115 8.14595
R323 VDD2.n141 VDD2.n134 8.14595
R324 VDD2.n37 VDD2.n30 8.14595
R325 VDD2.n75 VDD2.n12 8.14595
R326 VDD2.n84 VDD2.n83 8.14595
R327 VDD2.n183 VDD2.n111 7.3702
R328 VDD2.n179 VDD2.n113 7.3702
R329 VDD2.n138 VDD2.n137 7.3702
R330 VDD2.n34 VDD2.n33 7.3702
R331 VDD2.n76 VDD2.n10 7.3702
R332 VDD2.n80 VDD2.n8 7.3702
R333 VDD2.n183 VDD2.n182 6.59444
R334 VDD2.n182 VDD2.n113 6.59444
R335 VDD2.n79 VDD2.n10 6.59444
R336 VDD2.n80 VDD2.n79 6.59444
R337 VDD2.n186 VDD2.n111 5.81868
R338 VDD2.n179 VDD2.n178 5.81868
R339 VDD2.n138 VDD2.n134 5.81868
R340 VDD2.n34 VDD2.n30 5.81868
R341 VDD2.n76 VDD2.n75 5.81868
R342 VDD2.n83 VDD2.n8 5.81868
R343 VDD2.n187 VDD2.n109 5.04292
R344 VDD2.n175 VDD2.n115 5.04292
R345 VDD2.n142 VDD2.n141 5.04292
R346 VDD2.n38 VDD2.n37 5.04292
R347 VDD2.n72 VDD2.n12 5.04292
R348 VDD2.n84 VDD2.n6 5.04292
R349 VDD2.n191 VDD2.n190 4.26717
R350 VDD2.n174 VDD2.n117 4.26717
R351 VDD2.n145 VDD2.n132 4.26717
R352 VDD2.n41 VDD2.n28 4.26717
R353 VDD2.n71 VDD2.n14 4.26717
R354 VDD2.n88 VDD2.n87 4.26717
R355 VDD2.n194 VDD2.n107 3.49141
R356 VDD2.n171 VDD2.n170 3.49141
R357 VDD2.n146 VDD2.n130 3.49141
R358 VDD2.n42 VDD2.n26 3.49141
R359 VDD2.n68 VDD2.n67 3.49141
R360 VDD2.n91 VDD2.n4 3.49141
R361 VDD2.n139 VDD2.n135 2.84303
R362 VDD2.n35 VDD2.n31 2.84303
R363 VDD2.n195 VDD2.n105 2.71565
R364 VDD2.n167 VDD2.n119 2.71565
R365 VDD2.n150 VDD2.n149 2.71565
R366 VDD2.n46 VDD2.n45 2.71565
R367 VDD2.n64 VDD2.n16 2.71565
R368 VDD2.n92 VDD2.n2 2.71565
R369 VDD2.n204 VDD2.n202 2.40567
R370 VDD2.n199 VDD2.n198 1.93989
R371 VDD2.n166 VDD2.n121 1.93989
R372 VDD2.n153 VDD2.n127 1.93989
R373 VDD2.n50 VDD2.n24 1.93989
R374 VDD2.n63 VDD2.n18 1.93989
R375 VDD2.n96 VDD2.n95 1.93989
R376 VDD2.n201 VDD2.n103 1.16414
R377 VDD2.n163 VDD2.n162 1.16414
R378 VDD2.n154 VDD2.n125 1.16414
R379 VDD2.n51 VDD2.n22 1.16414
R380 VDD2.n60 VDD2.n59 1.16414
R381 VDD2.n98 VDD2.n0 1.16414
R382 VDD2.n205 VDD2.t6 1.09503
R383 VDD2.n205 VDD2.t9 1.09503
R384 VDD2.n203 VDD2.t1 1.09503
R385 VDD2.n203 VDD2.t2 1.09503
R386 VDD2.n101 VDD2.t5 1.09503
R387 VDD2.n101 VDD2.t8 1.09503
R388 VDD2.n99 VDD2.t4 1.09503
R389 VDD2.n99 VDD2.t0 1.09503
R390 VDD2 VDD2.n204 0.659983
R391 VDD2.n102 VDD2.n100 0.546447
R392 VDD2.n159 VDD2.n123 0.388379
R393 VDD2.n158 VDD2.n157 0.388379
R394 VDD2.n55 VDD2.n54 0.388379
R395 VDD2.n56 VDD2.n20 0.388379
R396 VDD2.n197 VDD2.n196 0.155672
R397 VDD2.n196 VDD2.n106 0.155672
R398 VDD2.n189 VDD2.n106 0.155672
R399 VDD2.n189 VDD2.n188 0.155672
R400 VDD2.n188 VDD2.n110 0.155672
R401 VDD2.n181 VDD2.n110 0.155672
R402 VDD2.n181 VDD2.n180 0.155672
R403 VDD2.n180 VDD2.n114 0.155672
R404 VDD2.n173 VDD2.n114 0.155672
R405 VDD2.n173 VDD2.n172 0.155672
R406 VDD2.n172 VDD2.n118 0.155672
R407 VDD2.n165 VDD2.n118 0.155672
R408 VDD2.n165 VDD2.n164 0.155672
R409 VDD2.n164 VDD2.n122 0.155672
R410 VDD2.n156 VDD2.n122 0.155672
R411 VDD2.n156 VDD2.n155 0.155672
R412 VDD2.n155 VDD2.n126 0.155672
R413 VDD2.n148 VDD2.n126 0.155672
R414 VDD2.n148 VDD2.n147 0.155672
R415 VDD2.n147 VDD2.n131 0.155672
R416 VDD2.n140 VDD2.n131 0.155672
R417 VDD2.n140 VDD2.n139 0.155672
R418 VDD2.n36 VDD2.n35 0.155672
R419 VDD2.n36 VDD2.n27 0.155672
R420 VDD2.n43 VDD2.n27 0.155672
R421 VDD2.n44 VDD2.n43 0.155672
R422 VDD2.n44 VDD2.n23 0.155672
R423 VDD2.n52 VDD2.n23 0.155672
R424 VDD2.n53 VDD2.n52 0.155672
R425 VDD2.n53 VDD2.n19 0.155672
R426 VDD2.n61 VDD2.n19 0.155672
R427 VDD2.n62 VDD2.n61 0.155672
R428 VDD2.n62 VDD2.n15 0.155672
R429 VDD2.n69 VDD2.n15 0.155672
R430 VDD2.n70 VDD2.n69 0.155672
R431 VDD2.n70 VDD2.n11 0.155672
R432 VDD2.n77 VDD2.n11 0.155672
R433 VDD2.n78 VDD2.n77 0.155672
R434 VDD2.n78 VDD2.n7 0.155672
R435 VDD2.n85 VDD2.n7 0.155672
R436 VDD2.n86 VDD2.n85 0.155672
R437 VDD2.n86 VDD2.n3 0.155672
R438 VDD2.n93 VDD2.n3 0.155672
R439 VDD2.n94 VDD2.n93 0.155672
R440 VTAIL.n412 VTAIL.n411 289.615
R441 VTAIL.n100 VTAIL.n99 289.615
R442 VTAIL.n312 VTAIL.n311 289.615
R443 VTAIL.n208 VTAIL.n207 289.615
R444 VTAIL.n347 VTAIL.n346 185
R445 VTAIL.n344 VTAIL.n343 185
R446 VTAIL.n353 VTAIL.n352 185
R447 VTAIL.n355 VTAIL.n354 185
R448 VTAIL.n340 VTAIL.n339 185
R449 VTAIL.n361 VTAIL.n360 185
R450 VTAIL.n364 VTAIL.n363 185
R451 VTAIL.n362 VTAIL.n336 185
R452 VTAIL.n369 VTAIL.n335 185
R453 VTAIL.n371 VTAIL.n370 185
R454 VTAIL.n373 VTAIL.n372 185
R455 VTAIL.n332 VTAIL.n331 185
R456 VTAIL.n379 VTAIL.n378 185
R457 VTAIL.n381 VTAIL.n380 185
R458 VTAIL.n328 VTAIL.n327 185
R459 VTAIL.n387 VTAIL.n386 185
R460 VTAIL.n389 VTAIL.n388 185
R461 VTAIL.n324 VTAIL.n323 185
R462 VTAIL.n395 VTAIL.n394 185
R463 VTAIL.n397 VTAIL.n396 185
R464 VTAIL.n320 VTAIL.n319 185
R465 VTAIL.n403 VTAIL.n402 185
R466 VTAIL.n405 VTAIL.n404 185
R467 VTAIL.n316 VTAIL.n315 185
R468 VTAIL.n411 VTAIL.n410 185
R469 VTAIL.n35 VTAIL.n34 185
R470 VTAIL.n32 VTAIL.n31 185
R471 VTAIL.n41 VTAIL.n40 185
R472 VTAIL.n43 VTAIL.n42 185
R473 VTAIL.n28 VTAIL.n27 185
R474 VTAIL.n49 VTAIL.n48 185
R475 VTAIL.n52 VTAIL.n51 185
R476 VTAIL.n50 VTAIL.n24 185
R477 VTAIL.n57 VTAIL.n23 185
R478 VTAIL.n59 VTAIL.n58 185
R479 VTAIL.n61 VTAIL.n60 185
R480 VTAIL.n20 VTAIL.n19 185
R481 VTAIL.n67 VTAIL.n66 185
R482 VTAIL.n69 VTAIL.n68 185
R483 VTAIL.n16 VTAIL.n15 185
R484 VTAIL.n75 VTAIL.n74 185
R485 VTAIL.n77 VTAIL.n76 185
R486 VTAIL.n12 VTAIL.n11 185
R487 VTAIL.n83 VTAIL.n82 185
R488 VTAIL.n85 VTAIL.n84 185
R489 VTAIL.n8 VTAIL.n7 185
R490 VTAIL.n91 VTAIL.n90 185
R491 VTAIL.n93 VTAIL.n92 185
R492 VTAIL.n4 VTAIL.n3 185
R493 VTAIL.n99 VTAIL.n98 185
R494 VTAIL.n311 VTAIL.n310 185
R495 VTAIL.n216 VTAIL.n215 185
R496 VTAIL.n305 VTAIL.n304 185
R497 VTAIL.n303 VTAIL.n302 185
R498 VTAIL.n220 VTAIL.n219 185
R499 VTAIL.n297 VTAIL.n296 185
R500 VTAIL.n295 VTAIL.n294 185
R501 VTAIL.n224 VTAIL.n223 185
R502 VTAIL.n289 VTAIL.n288 185
R503 VTAIL.n287 VTAIL.n286 185
R504 VTAIL.n228 VTAIL.n227 185
R505 VTAIL.n281 VTAIL.n280 185
R506 VTAIL.n279 VTAIL.n278 185
R507 VTAIL.n232 VTAIL.n231 185
R508 VTAIL.n273 VTAIL.n272 185
R509 VTAIL.n271 VTAIL.n270 185
R510 VTAIL.n269 VTAIL.n235 185
R511 VTAIL.n239 VTAIL.n236 185
R512 VTAIL.n264 VTAIL.n263 185
R513 VTAIL.n262 VTAIL.n261 185
R514 VTAIL.n241 VTAIL.n240 185
R515 VTAIL.n256 VTAIL.n255 185
R516 VTAIL.n254 VTAIL.n253 185
R517 VTAIL.n245 VTAIL.n244 185
R518 VTAIL.n248 VTAIL.n247 185
R519 VTAIL.n207 VTAIL.n206 185
R520 VTAIL.n112 VTAIL.n111 185
R521 VTAIL.n201 VTAIL.n200 185
R522 VTAIL.n199 VTAIL.n198 185
R523 VTAIL.n116 VTAIL.n115 185
R524 VTAIL.n193 VTAIL.n192 185
R525 VTAIL.n191 VTAIL.n190 185
R526 VTAIL.n120 VTAIL.n119 185
R527 VTAIL.n185 VTAIL.n184 185
R528 VTAIL.n183 VTAIL.n182 185
R529 VTAIL.n124 VTAIL.n123 185
R530 VTAIL.n177 VTAIL.n176 185
R531 VTAIL.n175 VTAIL.n174 185
R532 VTAIL.n128 VTAIL.n127 185
R533 VTAIL.n169 VTAIL.n168 185
R534 VTAIL.n167 VTAIL.n166 185
R535 VTAIL.n165 VTAIL.n131 185
R536 VTAIL.n135 VTAIL.n132 185
R537 VTAIL.n160 VTAIL.n159 185
R538 VTAIL.n158 VTAIL.n157 185
R539 VTAIL.n137 VTAIL.n136 185
R540 VTAIL.n152 VTAIL.n151 185
R541 VTAIL.n150 VTAIL.n149 185
R542 VTAIL.n141 VTAIL.n140 185
R543 VTAIL.n144 VTAIL.n143 185
R544 VTAIL.t8 VTAIL.n345 149.524
R545 VTAIL.t4 VTAIL.n33 149.524
R546 VTAIL.t2 VTAIL.n246 149.524
R547 VTAIL.t9 VTAIL.n142 149.524
R548 VTAIL.n346 VTAIL.n343 104.615
R549 VTAIL.n353 VTAIL.n343 104.615
R550 VTAIL.n354 VTAIL.n353 104.615
R551 VTAIL.n354 VTAIL.n339 104.615
R552 VTAIL.n361 VTAIL.n339 104.615
R553 VTAIL.n363 VTAIL.n361 104.615
R554 VTAIL.n363 VTAIL.n362 104.615
R555 VTAIL.n362 VTAIL.n335 104.615
R556 VTAIL.n371 VTAIL.n335 104.615
R557 VTAIL.n372 VTAIL.n371 104.615
R558 VTAIL.n372 VTAIL.n331 104.615
R559 VTAIL.n379 VTAIL.n331 104.615
R560 VTAIL.n380 VTAIL.n379 104.615
R561 VTAIL.n380 VTAIL.n327 104.615
R562 VTAIL.n387 VTAIL.n327 104.615
R563 VTAIL.n388 VTAIL.n387 104.615
R564 VTAIL.n388 VTAIL.n323 104.615
R565 VTAIL.n395 VTAIL.n323 104.615
R566 VTAIL.n396 VTAIL.n395 104.615
R567 VTAIL.n396 VTAIL.n319 104.615
R568 VTAIL.n403 VTAIL.n319 104.615
R569 VTAIL.n404 VTAIL.n403 104.615
R570 VTAIL.n404 VTAIL.n315 104.615
R571 VTAIL.n411 VTAIL.n315 104.615
R572 VTAIL.n34 VTAIL.n31 104.615
R573 VTAIL.n41 VTAIL.n31 104.615
R574 VTAIL.n42 VTAIL.n41 104.615
R575 VTAIL.n42 VTAIL.n27 104.615
R576 VTAIL.n49 VTAIL.n27 104.615
R577 VTAIL.n51 VTAIL.n49 104.615
R578 VTAIL.n51 VTAIL.n50 104.615
R579 VTAIL.n50 VTAIL.n23 104.615
R580 VTAIL.n59 VTAIL.n23 104.615
R581 VTAIL.n60 VTAIL.n59 104.615
R582 VTAIL.n60 VTAIL.n19 104.615
R583 VTAIL.n67 VTAIL.n19 104.615
R584 VTAIL.n68 VTAIL.n67 104.615
R585 VTAIL.n68 VTAIL.n15 104.615
R586 VTAIL.n75 VTAIL.n15 104.615
R587 VTAIL.n76 VTAIL.n75 104.615
R588 VTAIL.n76 VTAIL.n11 104.615
R589 VTAIL.n83 VTAIL.n11 104.615
R590 VTAIL.n84 VTAIL.n83 104.615
R591 VTAIL.n84 VTAIL.n7 104.615
R592 VTAIL.n91 VTAIL.n7 104.615
R593 VTAIL.n92 VTAIL.n91 104.615
R594 VTAIL.n92 VTAIL.n3 104.615
R595 VTAIL.n99 VTAIL.n3 104.615
R596 VTAIL.n311 VTAIL.n215 104.615
R597 VTAIL.n304 VTAIL.n215 104.615
R598 VTAIL.n304 VTAIL.n303 104.615
R599 VTAIL.n303 VTAIL.n219 104.615
R600 VTAIL.n296 VTAIL.n219 104.615
R601 VTAIL.n296 VTAIL.n295 104.615
R602 VTAIL.n295 VTAIL.n223 104.615
R603 VTAIL.n288 VTAIL.n223 104.615
R604 VTAIL.n288 VTAIL.n287 104.615
R605 VTAIL.n287 VTAIL.n227 104.615
R606 VTAIL.n280 VTAIL.n227 104.615
R607 VTAIL.n280 VTAIL.n279 104.615
R608 VTAIL.n279 VTAIL.n231 104.615
R609 VTAIL.n272 VTAIL.n231 104.615
R610 VTAIL.n272 VTAIL.n271 104.615
R611 VTAIL.n271 VTAIL.n235 104.615
R612 VTAIL.n239 VTAIL.n235 104.615
R613 VTAIL.n263 VTAIL.n239 104.615
R614 VTAIL.n263 VTAIL.n262 104.615
R615 VTAIL.n262 VTAIL.n240 104.615
R616 VTAIL.n255 VTAIL.n240 104.615
R617 VTAIL.n255 VTAIL.n254 104.615
R618 VTAIL.n254 VTAIL.n244 104.615
R619 VTAIL.n247 VTAIL.n244 104.615
R620 VTAIL.n207 VTAIL.n111 104.615
R621 VTAIL.n200 VTAIL.n111 104.615
R622 VTAIL.n200 VTAIL.n199 104.615
R623 VTAIL.n199 VTAIL.n115 104.615
R624 VTAIL.n192 VTAIL.n115 104.615
R625 VTAIL.n192 VTAIL.n191 104.615
R626 VTAIL.n191 VTAIL.n119 104.615
R627 VTAIL.n184 VTAIL.n119 104.615
R628 VTAIL.n184 VTAIL.n183 104.615
R629 VTAIL.n183 VTAIL.n123 104.615
R630 VTAIL.n176 VTAIL.n123 104.615
R631 VTAIL.n176 VTAIL.n175 104.615
R632 VTAIL.n175 VTAIL.n127 104.615
R633 VTAIL.n168 VTAIL.n127 104.615
R634 VTAIL.n168 VTAIL.n167 104.615
R635 VTAIL.n167 VTAIL.n131 104.615
R636 VTAIL.n135 VTAIL.n131 104.615
R637 VTAIL.n159 VTAIL.n135 104.615
R638 VTAIL.n159 VTAIL.n158 104.615
R639 VTAIL.n158 VTAIL.n136 104.615
R640 VTAIL.n151 VTAIL.n136 104.615
R641 VTAIL.n151 VTAIL.n150 104.615
R642 VTAIL.n150 VTAIL.n140 104.615
R643 VTAIL.n143 VTAIL.n140 104.615
R644 VTAIL.n346 VTAIL.t8 52.3082
R645 VTAIL.n34 VTAIL.t4 52.3082
R646 VTAIL.n247 VTAIL.t2 52.3082
R647 VTAIL.n143 VTAIL.t9 52.3082
R648 VTAIL.n213 VTAIL.n212 47.5008
R649 VTAIL.n211 VTAIL.n210 47.5008
R650 VTAIL.n109 VTAIL.n108 47.5008
R651 VTAIL.n107 VTAIL.n106 47.5008
R652 VTAIL.n415 VTAIL.n414 47.5007
R653 VTAIL.n1 VTAIL.n0 47.5007
R654 VTAIL.n103 VTAIL.n102 47.5007
R655 VTAIL.n105 VTAIL.n104 47.5007
R656 VTAIL.n413 VTAIL.n412 35.0944
R657 VTAIL.n101 VTAIL.n100 35.0944
R658 VTAIL.n313 VTAIL.n312 35.0944
R659 VTAIL.n209 VTAIL.n208 35.0944
R660 VTAIL.n107 VTAIL.n105 32.7721
R661 VTAIL.n413 VTAIL.n313 30.3669
R662 VTAIL.n370 VTAIL.n369 13.1884
R663 VTAIL.n58 VTAIL.n57 13.1884
R664 VTAIL.n270 VTAIL.n269 13.1884
R665 VTAIL.n166 VTAIL.n165 13.1884
R666 VTAIL.n368 VTAIL.n336 12.8005
R667 VTAIL.n373 VTAIL.n334 12.8005
R668 VTAIL.n56 VTAIL.n24 12.8005
R669 VTAIL.n61 VTAIL.n22 12.8005
R670 VTAIL.n273 VTAIL.n234 12.8005
R671 VTAIL.n268 VTAIL.n236 12.8005
R672 VTAIL.n169 VTAIL.n130 12.8005
R673 VTAIL.n164 VTAIL.n132 12.8005
R674 VTAIL.n365 VTAIL.n364 12.0247
R675 VTAIL.n374 VTAIL.n332 12.0247
R676 VTAIL.n410 VTAIL.n314 12.0247
R677 VTAIL.n53 VTAIL.n52 12.0247
R678 VTAIL.n62 VTAIL.n20 12.0247
R679 VTAIL.n98 VTAIL.n2 12.0247
R680 VTAIL.n310 VTAIL.n214 12.0247
R681 VTAIL.n274 VTAIL.n232 12.0247
R682 VTAIL.n265 VTAIL.n264 12.0247
R683 VTAIL.n206 VTAIL.n110 12.0247
R684 VTAIL.n170 VTAIL.n128 12.0247
R685 VTAIL.n161 VTAIL.n160 12.0247
R686 VTAIL.n360 VTAIL.n338 11.249
R687 VTAIL.n378 VTAIL.n377 11.249
R688 VTAIL.n409 VTAIL.n316 11.249
R689 VTAIL.n48 VTAIL.n26 11.249
R690 VTAIL.n66 VTAIL.n65 11.249
R691 VTAIL.n97 VTAIL.n4 11.249
R692 VTAIL.n309 VTAIL.n216 11.249
R693 VTAIL.n278 VTAIL.n277 11.249
R694 VTAIL.n261 VTAIL.n238 11.249
R695 VTAIL.n205 VTAIL.n112 11.249
R696 VTAIL.n174 VTAIL.n173 11.249
R697 VTAIL.n157 VTAIL.n134 11.249
R698 VTAIL.n359 VTAIL.n340 10.4732
R699 VTAIL.n381 VTAIL.n330 10.4732
R700 VTAIL.n406 VTAIL.n405 10.4732
R701 VTAIL.n47 VTAIL.n28 10.4732
R702 VTAIL.n69 VTAIL.n18 10.4732
R703 VTAIL.n94 VTAIL.n93 10.4732
R704 VTAIL.n306 VTAIL.n305 10.4732
R705 VTAIL.n281 VTAIL.n230 10.4732
R706 VTAIL.n260 VTAIL.n241 10.4732
R707 VTAIL.n202 VTAIL.n201 10.4732
R708 VTAIL.n177 VTAIL.n126 10.4732
R709 VTAIL.n156 VTAIL.n137 10.4732
R710 VTAIL.n347 VTAIL.n345 10.2747
R711 VTAIL.n35 VTAIL.n33 10.2747
R712 VTAIL.n248 VTAIL.n246 10.2747
R713 VTAIL.n144 VTAIL.n142 10.2747
R714 VTAIL.n356 VTAIL.n355 9.69747
R715 VTAIL.n382 VTAIL.n328 9.69747
R716 VTAIL.n402 VTAIL.n318 9.69747
R717 VTAIL.n44 VTAIL.n43 9.69747
R718 VTAIL.n70 VTAIL.n16 9.69747
R719 VTAIL.n90 VTAIL.n6 9.69747
R720 VTAIL.n302 VTAIL.n218 9.69747
R721 VTAIL.n282 VTAIL.n228 9.69747
R722 VTAIL.n257 VTAIL.n256 9.69747
R723 VTAIL.n198 VTAIL.n114 9.69747
R724 VTAIL.n178 VTAIL.n124 9.69747
R725 VTAIL.n153 VTAIL.n152 9.69747
R726 VTAIL.n408 VTAIL.n314 9.45567
R727 VTAIL.n96 VTAIL.n2 9.45567
R728 VTAIL.n308 VTAIL.n214 9.45567
R729 VTAIL.n204 VTAIL.n110 9.45567
R730 VTAIL.n393 VTAIL.n392 9.3005
R731 VTAIL.n322 VTAIL.n321 9.3005
R732 VTAIL.n399 VTAIL.n398 9.3005
R733 VTAIL.n401 VTAIL.n400 9.3005
R734 VTAIL.n318 VTAIL.n317 9.3005
R735 VTAIL.n407 VTAIL.n406 9.3005
R736 VTAIL.n409 VTAIL.n408 9.3005
R737 VTAIL.n326 VTAIL.n325 9.3005
R738 VTAIL.n385 VTAIL.n384 9.3005
R739 VTAIL.n383 VTAIL.n382 9.3005
R740 VTAIL.n330 VTAIL.n329 9.3005
R741 VTAIL.n377 VTAIL.n376 9.3005
R742 VTAIL.n375 VTAIL.n374 9.3005
R743 VTAIL.n334 VTAIL.n333 9.3005
R744 VTAIL.n349 VTAIL.n348 9.3005
R745 VTAIL.n351 VTAIL.n350 9.3005
R746 VTAIL.n342 VTAIL.n341 9.3005
R747 VTAIL.n357 VTAIL.n356 9.3005
R748 VTAIL.n359 VTAIL.n358 9.3005
R749 VTAIL.n338 VTAIL.n337 9.3005
R750 VTAIL.n366 VTAIL.n365 9.3005
R751 VTAIL.n368 VTAIL.n367 9.3005
R752 VTAIL.n391 VTAIL.n390 9.3005
R753 VTAIL.n81 VTAIL.n80 9.3005
R754 VTAIL.n10 VTAIL.n9 9.3005
R755 VTAIL.n87 VTAIL.n86 9.3005
R756 VTAIL.n89 VTAIL.n88 9.3005
R757 VTAIL.n6 VTAIL.n5 9.3005
R758 VTAIL.n95 VTAIL.n94 9.3005
R759 VTAIL.n97 VTAIL.n96 9.3005
R760 VTAIL.n14 VTAIL.n13 9.3005
R761 VTAIL.n73 VTAIL.n72 9.3005
R762 VTAIL.n71 VTAIL.n70 9.3005
R763 VTAIL.n18 VTAIL.n17 9.3005
R764 VTAIL.n65 VTAIL.n64 9.3005
R765 VTAIL.n63 VTAIL.n62 9.3005
R766 VTAIL.n22 VTAIL.n21 9.3005
R767 VTAIL.n37 VTAIL.n36 9.3005
R768 VTAIL.n39 VTAIL.n38 9.3005
R769 VTAIL.n30 VTAIL.n29 9.3005
R770 VTAIL.n45 VTAIL.n44 9.3005
R771 VTAIL.n47 VTAIL.n46 9.3005
R772 VTAIL.n26 VTAIL.n25 9.3005
R773 VTAIL.n54 VTAIL.n53 9.3005
R774 VTAIL.n56 VTAIL.n55 9.3005
R775 VTAIL.n79 VTAIL.n78 9.3005
R776 VTAIL.n309 VTAIL.n308 9.3005
R777 VTAIL.n307 VTAIL.n306 9.3005
R778 VTAIL.n218 VTAIL.n217 9.3005
R779 VTAIL.n301 VTAIL.n300 9.3005
R780 VTAIL.n299 VTAIL.n298 9.3005
R781 VTAIL.n222 VTAIL.n221 9.3005
R782 VTAIL.n293 VTAIL.n292 9.3005
R783 VTAIL.n291 VTAIL.n290 9.3005
R784 VTAIL.n226 VTAIL.n225 9.3005
R785 VTAIL.n285 VTAIL.n284 9.3005
R786 VTAIL.n283 VTAIL.n282 9.3005
R787 VTAIL.n230 VTAIL.n229 9.3005
R788 VTAIL.n277 VTAIL.n276 9.3005
R789 VTAIL.n275 VTAIL.n274 9.3005
R790 VTAIL.n234 VTAIL.n233 9.3005
R791 VTAIL.n268 VTAIL.n267 9.3005
R792 VTAIL.n266 VTAIL.n265 9.3005
R793 VTAIL.n238 VTAIL.n237 9.3005
R794 VTAIL.n260 VTAIL.n259 9.3005
R795 VTAIL.n258 VTAIL.n257 9.3005
R796 VTAIL.n243 VTAIL.n242 9.3005
R797 VTAIL.n252 VTAIL.n251 9.3005
R798 VTAIL.n250 VTAIL.n249 9.3005
R799 VTAIL.n146 VTAIL.n145 9.3005
R800 VTAIL.n148 VTAIL.n147 9.3005
R801 VTAIL.n139 VTAIL.n138 9.3005
R802 VTAIL.n154 VTAIL.n153 9.3005
R803 VTAIL.n156 VTAIL.n155 9.3005
R804 VTAIL.n134 VTAIL.n133 9.3005
R805 VTAIL.n162 VTAIL.n161 9.3005
R806 VTAIL.n164 VTAIL.n163 9.3005
R807 VTAIL.n118 VTAIL.n117 9.3005
R808 VTAIL.n195 VTAIL.n194 9.3005
R809 VTAIL.n197 VTAIL.n196 9.3005
R810 VTAIL.n114 VTAIL.n113 9.3005
R811 VTAIL.n203 VTAIL.n202 9.3005
R812 VTAIL.n205 VTAIL.n204 9.3005
R813 VTAIL.n189 VTAIL.n188 9.3005
R814 VTAIL.n187 VTAIL.n186 9.3005
R815 VTAIL.n122 VTAIL.n121 9.3005
R816 VTAIL.n181 VTAIL.n180 9.3005
R817 VTAIL.n179 VTAIL.n178 9.3005
R818 VTAIL.n126 VTAIL.n125 9.3005
R819 VTAIL.n173 VTAIL.n172 9.3005
R820 VTAIL.n171 VTAIL.n170 9.3005
R821 VTAIL.n130 VTAIL.n129 9.3005
R822 VTAIL.n352 VTAIL.n342 8.92171
R823 VTAIL.n386 VTAIL.n385 8.92171
R824 VTAIL.n401 VTAIL.n320 8.92171
R825 VTAIL.n40 VTAIL.n30 8.92171
R826 VTAIL.n74 VTAIL.n73 8.92171
R827 VTAIL.n89 VTAIL.n8 8.92171
R828 VTAIL.n301 VTAIL.n220 8.92171
R829 VTAIL.n286 VTAIL.n285 8.92171
R830 VTAIL.n253 VTAIL.n243 8.92171
R831 VTAIL.n197 VTAIL.n116 8.92171
R832 VTAIL.n182 VTAIL.n181 8.92171
R833 VTAIL.n149 VTAIL.n139 8.92171
R834 VTAIL.n351 VTAIL.n344 8.14595
R835 VTAIL.n389 VTAIL.n326 8.14595
R836 VTAIL.n398 VTAIL.n397 8.14595
R837 VTAIL.n39 VTAIL.n32 8.14595
R838 VTAIL.n77 VTAIL.n14 8.14595
R839 VTAIL.n86 VTAIL.n85 8.14595
R840 VTAIL.n298 VTAIL.n297 8.14595
R841 VTAIL.n289 VTAIL.n226 8.14595
R842 VTAIL.n252 VTAIL.n245 8.14595
R843 VTAIL.n194 VTAIL.n193 8.14595
R844 VTAIL.n185 VTAIL.n122 8.14595
R845 VTAIL.n148 VTAIL.n141 8.14595
R846 VTAIL.n348 VTAIL.n347 7.3702
R847 VTAIL.n390 VTAIL.n324 7.3702
R848 VTAIL.n394 VTAIL.n322 7.3702
R849 VTAIL.n36 VTAIL.n35 7.3702
R850 VTAIL.n78 VTAIL.n12 7.3702
R851 VTAIL.n82 VTAIL.n10 7.3702
R852 VTAIL.n294 VTAIL.n222 7.3702
R853 VTAIL.n290 VTAIL.n224 7.3702
R854 VTAIL.n249 VTAIL.n248 7.3702
R855 VTAIL.n190 VTAIL.n118 7.3702
R856 VTAIL.n186 VTAIL.n120 7.3702
R857 VTAIL.n145 VTAIL.n144 7.3702
R858 VTAIL.n393 VTAIL.n324 6.59444
R859 VTAIL.n394 VTAIL.n393 6.59444
R860 VTAIL.n81 VTAIL.n12 6.59444
R861 VTAIL.n82 VTAIL.n81 6.59444
R862 VTAIL.n294 VTAIL.n293 6.59444
R863 VTAIL.n293 VTAIL.n224 6.59444
R864 VTAIL.n190 VTAIL.n189 6.59444
R865 VTAIL.n189 VTAIL.n120 6.59444
R866 VTAIL.n348 VTAIL.n344 5.81868
R867 VTAIL.n390 VTAIL.n389 5.81868
R868 VTAIL.n397 VTAIL.n322 5.81868
R869 VTAIL.n36 VTAIL.n32 5.81868
R870 VTAIL.n78 VTAIL.n77 5.81868
R871 VTAIL.n85 VTAIL.n10 5.81868
R872 VTAIL.n297 VTAIL.n222 5.81868
R873 VTAIL.n290 VTAIL.n289 5.81868
R874 VTAIL.n249 VTAIL.n245 5.81868
R875 VTAIL.n193 VTAIL.n118 5.81868
R876 VTAIL.n186 VTAIL.n185 5.81868
R877 VTAIL.n145 VTAIL.n141 5.81868
R878 VTAIL.n352 VTAIL.n351 5.04292
R879 VTAIL.n386 VTAIL.n326 5.04292
R880 VTAIL.n398 VTAIL.n320 5.04292
R881 VTAIL.n40 VTAIL.n39 5.04292
R882 VTAIL.n74 VTAIL.n14 5.04292
R883 VTAIL.n86 VTAIL.n8 5.04292
R884 VTAIL.n298 VTAIL.n220 5.04292
R885 VTAIL.n286 VTAIL.n226 5.04292
R886 VTAIL.n253 VTAIL.n252 5.04292
R887 VTAIL.n194 VTAIL.n116 5.04292
R888 VTAIL.n182 VTAIL.n122 5.04292
R889 VTAIL.n149 VTAIL.n148 5.04292
R890 VTAIL.n355 VTAIL.n342 4.26717
R891 VTAIL.n385 VTAIL.n328 4.26717
R892 VTAIL.n402 VTAIL.n401 4.26717
R893 VTAIL.n43 VTAIL.n30 4.26717
R894 VTAIL.n73 VTAIL.n16 4.26717
R895 VTAIL.n90 VTAIL.n89 4.26717
R896 VTAIL.n302 VTAIL.n301 4.26717
R897 VTAIL.n285 VTAIL.n228 4.26717
R898 VTAIL.n256 VTAIL.n243 4.26717
R899 VTAIL.n198 VTAIL.n197 4.26717
R900 VTAIL.n181 VTAIL.n124 4.26717
R901 VTAIL.n152 VTAIL.n139 4.26717
R902 VTAIL.n356 VTAIL.n340 3.49141
R903 VTAIL.n382 VTAIL.n381 3.49141
R904 VTAIL.n405 VTAIL.n318 3.49141
R905 VTAIL.n44 VTAIL.n28 3.49141
R906 VTAIL.n70 VTAIL.n69 3.49141
R907 VTAIL.n93 VTAIL.n6 3.49141
R908 VTAIL.n305 VTAIL.n218 3.49141
R909 VTAIL.n282 VTAIL.n281 3.49141
R910 VTAIL.n257 VTAIL.n241 3.49141
R911 VTAIL.n201 VTAIL.n114 3.49141
R912 VTAIL.n178 VTAIL.n177 3.49141
R913 VTAIL.n153 VTAIL.n137 3.49141
R914 VTAIL.n146 VTAIL.n142 2.84303
R915 VTAIL.n349 VTAIL.n345 2.84303
R916 VTAIL.n37 VTAIL.n33 2.84303
R917 VTAIL.n250 VTAIL.n246 2.84303
R918 VTAIL.n360 VTAIL.n359 2.71565
R919 VTAIL.n378 VTAIL.n330 2.71565
R920 VTAIL.n406 VTAIL.n316 2.71565
R921 VTAIL.n48 VTAIL.n47 2.71565
R922 VTAIL.n66 VTAIL.n18 2.71565
R923 VTAIL.n94 VTAIL.n4 2.71565
R924 VTAIL.n306 VTAIL.n216 2.71565
R925 VTAIL.n278 VTAIL.n230 2.71565
R926 VTAIL.n261 VTAIL.n260 2.71565
R927 VTAIL.n202 VTAIL.n112 2.71565
R928 VTAIL.n174 VTAIL.n126 2.71565
R929 VTAIL.n157 VTAIL.n156 2.71565
R930 VTAIL.n109 VTAIL.n107 2.40567
R931 VTAIL.n209 VTAIL.n109 2.40567
R932 VTAIL.n213 VTAIL.n211 2.40567
R933 VTAIL.n313 VTAIL.n213 2.40567
R934 VTAIL.n105 VTAIL.n103 2.40567
R935 VTAIL.n103 VTAIL.n101 2.40567
R936 VTAIL.n415 VTAIL.n413 2.40567
R937 VTAIL.n364 VTAIL.n338 1.93989
R938 VTAIL.n377 VTAIL.n332 1.93989
R939 VTAIL.n410 VTAIL.n409 1.93989
R940 VTAIL.n52 VTAIL.n26 1.93989
R941 VTAIL.n65 VTAIL.n20 1.93989
R942 VTAIL.n98 VTAIL.n97 1.93989
R943 VTAIL.n310 VTAIL.n309 1.93989
R944 VTAIL.n277 VTAIL.n232 1.93989
R945 VTAIL.n264 VTAIL.n238 1.93989
R946 VTAIL.n206 VTAIL.n205 1.93989
R947 VTAIL.n173 VTAIL.n128 1.93989
R948 VTAIL.n160 VTAIL.n134 1.93989
R949 VTAIL VTAIL.n1 1.86257
R950 VTAIL.n211 VTAIL.n209 1.67291
R951 VTAIL.n101 VTAIL.n1 1.67291
R952 VTAIL.n365 VTAIL.n336 1.16414
R953 VTAIL.n374 VTAIL.n373 1.16414
R954 VTAIL.n412 VTAIL.n314 1.16414
R955 VTAIL.n53 VTAIL.n24 1.16414
R956 VTAIL.n62 VTAIL.n61 1.16414
R957 VTAIL.n100 VTAIL.n2 1.16414
R958 VTAIL.n312 VTAIL.n214 1.16414
R959 VTAIL.n274 VTAIL.n273 1.16414
R960 VTAIL.n265 VTAIL.n236 1.16414
R961 VTAIL.n208 VTAIL.n110 1.16414
R962 VTAIL.n170 VTAIL.n169 1.16414
R963 VTAIL.n161 VTAIL.n132 1.16414
R964 VTAIL.n414 VTAIL.t14 1.09503
R965 VTAIL.n414 VTAIL.t16 1.09503
R966 VTAIL.n0 VTAIL.t13 1.09503
R967 VTAIL.n0 VTAIL.t7 1.09503
R968 VTAIL.n102 VTAIL.t17 1.09503
R969 VTAIL.n102 VTAIL.t6 1.09503
R970 VTAIL.n104 VTAIL.t0 1.09503
R971 VTAIL.n104 VTAIL.t3 1.09503
R972 VTAIL.n212 VTAIL.t5 1.09503
R973 VTAIL.n212 VTAIL.t19 1.09503
R974 VTAIL.n210 VTAIL.t18 1.09503
R975 VTAIL.n210 VTAIL.t1 1.09503
R976 VTAIL.n108 VTAIL.t12 1.09503
R977 VTAIL.n108 VTAIL.t10 1.09503
R978 VTAIL.n106 VTAIL.t11 1.09503
R979 VTAIL.n106 VTAIL.t15 1.09503
R980 VTAIL VTAIL.n415 0.543603
R981 VTAIL.n369 VTAIL.n368 0.388379
R982 VTAIL.n370 VTAIL.n334 0.388379
R983 VTAIL.n57 VTAIL.n56 0.388379
R984 VTAIL.n58 VTAIL.n22 0.388379
R985 VTAIL.n270 VTAIL.n234 0.388379
R986 VTAIL.n269 VTAIL.n268 0.388379
R987 VTAIL.n166 VTAIL.n130 0.388379
R988 VTAIL.n165 VTAIL.n164 0.388379
R989 VTAIL.n350 VTAIL.n349 0.155672
R990 VTAIL.n350 VTAIL.n341 0.155672
R991 VTAIL.n357 VTAIL.n341 0.155672
R992 VTAIL.n358 VTAIL.n357 0.155672
R993 VTAIL.n358 VTAIL.n337 0.155672
R994 VTAIL.n366 VTAIL.n337 0.155672
R995 VTAIL.n367 VTAIL.n366 0.155672
R996 VTAIL.n367 VTAIL.n333 0.155672
R997 VTAIL.n375 VTAIL.n333 0.155672
R998 VTAIL.n376 VTAIL.n375 0.155672
R999 VTAIL.n376 VTAIL.n329 0.155672
R1000 VTAIL.n383 VTAIL.n329 0.155672
R1001 VTAIL.n384 VTAIL.n383 0.155672
R1002 VTAIL.n384 VTAIL.n325 0.155672
R1003 VTAIL.n391 VTAIL.n325 0.155672
R1004 VTAIL.n392 VTAIL.n391 0.155672
R1005 VTAIL.n392 VTAIL.n321 0.155672
R1006 VTAIL.n399 VTAIL.n321 0.155672
R1007 VTAIL.n400 VTAIL.n399 0.155672
R1008 VTAIL.n400 VTAIL.n317 0.155672
R1009 VTAIL.n407 VTAIL.n317 0.155672
R1010 VTAIL.n408 VTAIL.n407 0.155672
R1011 VTAIL.n38 VTAIL.n37 0.155672
R1012 VTAIL.n38 VTAIL.n29 0.155672
R1013 VTAIL.n45 VTAIL.n29 0.155672
R1014 VTAIL.n46 VTAIL.n45 0.155672
R1015 VTAIL.n46 VTAIL.n25 0.155672
R1016 VTAIL.n54 VTAIL.n25 0.155672
R1017 VTAIL.n55 VTAIL.n54 0.155672
R1018 VTAIL.n55 VTAIL.n21 0.155672
R1019 VTAIL.n63 VTAIL.n21 0.155672
R1020 VTAIL.n64 VTAIL.n63 0.155672
R1021 VTAIL.n64 VTAIL.n17 0.155672
R1022 VTAIL.n71 VTAIL.n17 0.155672
R1023 VTAIL.n72 VTAIL.n71 0.155672
R1024 VTAIL.n72 VTAIL.n13 0.155672
R1025 VTAIL.n79 VTAIL.n13 0.155672
R1026 VTAIL.n80 VTAIL.n79 0.155672
R1027 VTAIL.n80 VTAIL.n9 0.155672
R1028 VTAIL.n87 VTAIL.n9 0.155672
R1029 VTAIL.n88 VTAIL.n87 0.155672
R1030 VTAIL.n88 VTAIL.n5 0.155672
R1031 VTAIL.n95 VTAIL.n5 0.155672
R1032 VTAIL.n96 VTAIL.n95 0.155672
R1033 VTAIL.n308 VTAIL.n307 0.155672
R1034 VTAIL.n307 VTAIL.n217 0.155672
R1035 VTAIL.n300 VTAIL.n217 0.155672
R1036 VTAIL.n300 VTAIL.n299 0.155672
R1037 VTAIL.n299 VTAIL.n221 0.155672
R1038 VTAIL.n292 VTAIL.n221 0.155672
R1039 VTAIL.n292 VTAIL.n291 0.155672
R1040 VTAIL.n291 VTAIL.n225 0.155672
R1041 VTAIL.n284 VTAIL.n225 0.155672
R1042 VTAIL.n284 VTAIL.n283 0.155672
R1043 VTAIL.n283 VTAIL.n229 0.155672
R1044 VTAIL.n276 VTAIL.n229 0.155672
R1045 VTAIL.n276 VTAIL.n275 0.155672
R1046 VTAIL.n275 VTAIL.n233 0.155672
R1047 VTAIL.n267 VTAIL.n233 0.155672
R1048 VTAIL.n267 VTAIL.n266 0.155672
R1049 VTAIL.n266 VTAIL.n237 0.155672
R1050 VTAIL.n259 VTAIL.n237 0.155672
R1051 VTAIL.n259 VTAIL.n258 0.155672
R1052 VTAIL.n258 VTAIL.n242 0.155672
R1053 VTAIL.n251 VTAIL.n242 0.155672
R1054 VTAIL.n251 VTAIL.n250 0.155672
R1055 VTAIL.n204 VTAIL.n203 0.155672
R1056 VTAIL.n203 VTAIL.n113 0.155672
R1057 VTAIL.n196 VTAIL.n113 0.155672
R1058 VTAIL.n196 VTAIL.n195 0.155672
R1059 VTAIL.n195 VTAIL.n117 0.155672
R1060 VTAIL.n188 VTAIL.n117 0.155672
R1061 VTAIL.n188 VTAIL.n187 0.155672
R1062 VTAIL.n187 VTAIL.n121 0.155672
R1063 VTAIL.n180 VTAIL.n121 0.155672
R1064 VTAIL.n180 VTAIL.n179 0.155672
R1065 VTAIL.n179 VTAIL.n125 0.155672
R1066 VTAIL.n172 VTAIL.n125 0.155672
R1067 VTAIL.n172 VTAIL.n171 0.155672
R1068 VTAIL.n171 VTAIL.n129 0.155672
R1069 VTAIL.n163 VTAIL.n129 0.155672
R1070 VTAIL.n163 VTAIL.n162 0.155672
R1071 VTAIL.n162 VTAIL.n133 0.155672
R1072 VTAIL.n155 VTAIL.n133 0.155672
R1073 VTAIL.n155 VTAIL.n154 0.155672
R1074 VTAIL.n154 VTAIL.n138 0.155672
R1075 VTAIL.n147 VTAIL.n138 0.155672
R1076 VTAIL.n147 VTAIL.n146 0.155672
R1077 B.n1118 B.n1117 585
R1078 B.n1119 B.n1118 585
R1079 B.n431 B.n170 585
R1080 B.n430 B.n429 585
R1081 B.n428 B.n427 585
R1082 B.n426 B.n425 585
R1083 B.n424 B.n423 585
R1084 B.n422 B.n421 585
R1085 B.n420 B.n419 585
R1086 B.n418 B.n417 585
R1087 B.n416 B.n415 585
R1088 B.n414 B.n413 585
R1089 B.n412 B.n411 585
R1090 B.n410 B.n409 585
R1091 B.n408 B.n407 585
R1092 B.n406 B.n405 585
R1093 B.n404 B.n403 585
R1094 B.n402 B.n401 585
R1095 B.n400 B.n399 585
R1096 B.n398 B.n397 585
R1097 B.n396 B.n395 585
R1098 B.n394 B.n393 585
R1099 B.n392 B.n391 585
R1100 B.n390 B.n389 585
R1101 B.n388 B.n387 585
R1102 B.n386 B.n385 585
R1103 B.n384 B.n383 585
R1104 B.n382 B.n381 585
R1105 B.n380 B.n379 585
R1106 B.n378 B.n377 585
R1107 B.n376 B.n375 585
R1108 B.n374 B.n373 585
R1109 B.n372 B.n371 585
R1110 B.n370 B.n369 585
R1111 B.n368 B.n367 585
R1112 B.n366 B.n365 585
R1113 B.n364 B.n363 585
R1114 B.n362 B.n361 585
R1115 B.n360 B.n359 585
R1116 B.n358 B.n357 585
R1117 B.n356 B.n355 585
R1118 B.n354 B.n353 585
R1119 B.n352 B.n351 585
R1120 B.n350 B.n349 585
R1121 B.n348 B.n347 585
R1122 B.n346 B.n345 585
R1123 B.n344 B.n343 585
R1124 B.n342 B.n341 585
R1125 B.n340 B.n339 585
R1126 B.n338 B.n337 585
R1127 B.n336 B.n335 585
R1128 B.n334 B.n333 585
R1129 B.n332 B.n331 585
R1130 B.n330 B.n329 585
R1131 B.n328 B.n327 585
R1132 B.n326 B.n325 585
R1133 B.n324 B.n323 585
R1134 B.n322 B.n321 585
R1135 B.n320 B.n319 585
R1136 B.n318 B.n317 585
R1137 B.n316 B.n315 585
R1138 B.n313 B.n312 585
R1139 B.n311 B.n310 585
R1140 B.n309 B.n308 585
R1141 B.n307 B.n306 585
R1142 B.n305 B.n304 585
R1143 B.n303 B.n302 585
R1144 B.n301 B.n300 585
R1145 B.n299 B.n298 585
R1146 B.n297 B.n296 585
R1147 B.n295 B.n294 585
R1148 B.n293 B.n292 585
R1149 B.n291 B.n290 585
R1150 B.n289 B.n288 585
R1151 B.n287 B.n286 585
R1152 B.n285 B.n284 585
R1153 B.n283 B.n282 585
R1154 B.n281 B.n280 585
R1155 B.n279 B.n278 585
R1156 B.n277 B.n276 585
R1157 B.n275 B.n274 585
R1158 B.n273 B.n272 585
R1159 B.n271 B.n270 585
R1160 B.n269 B.n268 585
R1161 B.n267 B.n266 585
R1162 B.n265 B.n264 585
R1163 B.n263 B.n262 585
R1164 B.n261 B.n260 585
R1165 B.n259 B.n258 585
R1166 B.n257 B.n256 585
R1167 B.n255 B.n254 585
R1168 B.n253 B.n252 585
R1169 B.n251 B.n250 585
R1170 B.n249 B.n248 585
R1171 B.n247 B.n246 585
R1172 B.n245 B.n244 585
R1173 B.n243 B.n242 585
R1174 B.n241 B.n240 585
R1175 B.n239 B.n238 585
R1176 B.n237 B.n236 585
R1177 B.n235 B.n234 585
R1178 B.n233 B.n232 585
R1179 B.n231 B.n230 585
R1180 B.n229 B.n228 585
R1181 B.n227 B.n226 585
R1182 B.n225 B.n224 585
R1183 B.n223 B.n222 585
R1184 B.n221 B.n220 585
R1185 B.n219 B.n218 585
R1186 B.n217 B.n216 585
R1187 B.n215 B.n214 585
R1188 B.n213 B.n212 585
R1189 B.n211 B.n210 585
R1190 B.n209 B.n208 585
R1191 B.n207 B.n206 585
R1192 B.n205 B.n204 585
R1193 B.n203 B.n202 585
R1194 B.n201 B.n200 585
R1195 B.n199 B.n198 585
R1196 B.n197 B.n196 585
R1197 B.n195 B.n194 585
R1198 B.n193 B.n192 585
R1199 B.n191 B.n190 585
R1200 B.n189 B.n188 585
R1201 B.n187 B.n186 585
R1202 B.n185 B.n184 585
R1203 B.n183 B.n182 585
R1204 B.n181 B.n180 585
R1205 B.n179 B.n178 585
R1206 B.n177 B.n176 585
R1207 B.n1116 B.n105 585
R1208 B.n1120 B.n105 585
R1209 B.n1115 B.n104 585
R1210 B.n1121 B.n104 585
R1211 B.n1114 B.n1113 585
R1212 B.n1113 B.n100 585
R1213 B.n1112 B.n99 585
R1214 B.n1127 B.n99 585
R1215 B.n1111 B.n98 585
R1216 B.n1128 B.n98 585
R1217 B.n1110 B.n97 585
R1218 B.n1129 B.n97 585
R1219 B.n1109 B.n1108 585
R1220 B.n1108 B.n93 585
R1221 B.n1107 B.n92 585
R1222 B.n1135 B.n92 585
R1223 B.n1106 B.n91 585
R1224 B.n1136 B.n91 585
R1225 B.n1105 B.n90 585
R1226 B.n1137 B.n90 585
R1227 B.n1104 B.n1103 585
R1228 B.n1103 B.n86 585
R1229 B.n1102 B.n85 585
R1230 B.n1143 B.n85 585
R1231 B.n1101 B.n84 585
R1232 B.n1144 B.n84 585
R1233 B.n1100 B.n83 585
R1234 B.n1145 B.n83 585
R1235 B.n1099 B.n1098 585
R1236 B.n1098 B.n79 585
R1237 B.n1097 B.n78 585
R1238 B.n1151 B.n78 585
R1239 B.n1096 B.n77 585
R1240 B.n1152 B.n77 585
R1241 B.n1095 B.n76 585
R1242 B.n1153 B.n76 585
R1243 B.n1094 B.n1093 585
R1244 B.n1093 B.n75 585
R1245 B.n1092 B.n71 585
R1246 B.n1159 B.n71 585
R1247 B.n1091 B.n70 585
R1248 B.n1160 B.n70 585
R1249 B.n1090 B.n69 585
R1250 B.n1161 B.n69 585
R1251 B.n1089 B.n1088 585
R1252 B.n1088 B.n65 585
R1253 B.n1087 B.n64 585
R1254 B.n1167 B.n64 585
R1255 B.n1086 B.n63 585
R1256 B.n1168 B.n63 585
R1257 B.n1085 B.n62 585
R1258 B.n1169 B.n62 585
R1259 B.n1084 B.n1083 585
R1260 B.n1083 B.n58 585
R1261 B.n1082 B.n57 585
R1262 B.n1175 B.n57 585
R1263 B.n1081 B.n56 585
R1264 B.n1176 B.n56 585
R1265 B.n1080 B.n55 585
R1266 B.n1177 B.n55 585
R1267 B.n1079 B.n1078 585
R1268 B.n1078 B.n51 585
R1269 B.n1077 B.n50 585
R1270 B.n1183 B.n50 585
R1271 B.n1076 B.n49 585
R1272 B.n1184 B.n49 585
R1273 B.n1075 B.n48 585
R1274 B.n1185 B.n48 585
R1275 B.n1074 B.n1073 585
R1276 B.n1073 B.n44 585
R1277 B.n1072 B.n43 585
R1278 B.n1191 B.n43 585
R1279 B.n1071 B.n42 585
R1280 B.n1192 B.n42 585
R1281 B.n1070 B.n41 585
R1282 B.n1193 B.n41 585
R1283 B.n1069 B.n1068 585
R1284 B.n1068 B.n37 585
R1285 B.n1067 B.n36 585
R1286 B.n1199 B.n36 585
R1287 B.n1066 B.n35 585
R1288 B.n1200 B.n35 585
R1289 B.n1065 B.n34 585
R1290 B.n1201 B.n34 585
R1291 B.n1064 B.n1063 585
R1292 B.n1063 B.n30 585
R1293 B.n1062 B.n29 585
R1294 B.n1207 B.n29 585
R1295 B.n1061 B.n28 585
R1296 B.n1208 B.n28 585
R1297 B.n1060 B.n27 585
R1298 B.n1209 B.n27 585
R1299 B.n1059 B.n1058 585
R1300 B.n1058 B.n23 585
R1301 B.n1057 B.n22 585
R1302 B.n1215 B.n22 585
R1303 B.n1056 B.n21 585
R1304 B.n1216 B.n21 585
R1305 B.n1055 B.n20 585
R1306 B.n1217 B.n20 585
R1307 B.n1054 B.n1053 585
R1308 B.n1053 B.n16 585
R1309 B.n1052 B.n15 585
R1310 B.n1223 B.n15 585
R1311 B.n1051 B.n14 585
R1312 B.n1224 B.n14 585
R1313 B.n1050 B.n13 585
R1314 B.n1225 B.n13 585
R1315 B.n1049 B.n1048 585
R1316 B.n1048 B.n12 585
R1317 B.n1047 B.n1046 585
R1318 B.n1047 B.n8 585
R1319 B.n1045 B.n7 585
R1320 B.n1232 B.n7 585
R1321 B.n1044 B.n6 585
R1322 B.n1233 B.n6 585
R1323 B.n1043 B.n5 585
R1324 B.n1234 B.n5 585
R1325 B.n1042 B.n1041 585
R1326 B.n1041 B.n4 585
R1327 B.n1040 B.n432 585
R1328 B.n1040 B.n1039 585
R1329 B.n1030 B.n433 585
R1330 B.n434 B.n433 585
R1331 B.n1032 B.n1031 585
R1332 B.n1033 B.n1032 585
R1333 B.n1029 B.n439 585
R1334 B.n439 B.n438 585
R1335 B.n1028 B.n1027 585
R1336 B.n1027 B.n1026 585
R1337 B.n441 B.n440 585
R1338 B.n442 B.n441 585
R1339 B.n1019 B.n1018 585
R1340 B.n1020 B.n1019 585
R1341 B.n1017 B.n447 585
R1342 B.n447 B.n446 585
R1343 B.n1016 B.n1015 585
R1344 B.n1015 B.n1014 585
R1345 B.n449 B.n448 585
R1346 B.n450 B.n449 585
R1347 B.n1007 B.n1006 585
R1348 B.n1008 B.n1007 585
R1349 B.n1005 B.n455 585
R1350 B.n455 B.n454 585
R1351 B.n1004 B.n1003 585
R1352 B.n1003 B.n1002 585
R1353 B.n457 B.n456 585
R1354 B.n458 B.n457 585
R1355 B.n995 B.n994 585
R1356 B.n996 B.n995 585
R1357 B.n993 B.n463 585
R1358 B.n463 B.n462 585
R1359 B.n992 B.n991 585
R1360 B.n991 B.n990 585
R1361 B.n465 B.n464 585
R1362 B.n466 B.n465 585
R1363 B.n983 B.n982 585
R1364 B.n984 B.n983 585
R1365 B.n981 B.n471 585
R1366 B.n471 B.n470 585
R1367 B.n980 B.n979 585
R1368 B.n979 B.n978 585
R1369 B.n473 B.n472 585
R1370 B.n474 B.n473 585
R1371 B.n971 B.n970 585
R1372 B.n972 B.n971 585
R1373 B.n969 B.n479 585
R1374 B.n479 B.n478 585
R1375 B.n968 B.n967 585
R1376 B.n967 B.n966 585
R1377 B.n481 B.n480 585
R1378 B.n482 B.n481 585
R1379 B.n959 B.n958 585
R1380 B.n960 B.n959 585
R1381 B.n957 B.n487 585
R1382 B.n487 B.n486 585
R1383 B.n956 B.n955 585
R1384 B.n955 B.n954 585
R1385 B.n489 B.n488 585
R1386 B.n490 B.n489 585
R1387 B.n947 B.n946 585
R1388 B.n948 B.n947 585
R1389 B.n945 B.n495 585
R1390 B.n495 B.n494 585
R1391 B.n944 B.n943 585
R1392 B.n943 B.n942 585
R1393 B.n497 B.n496 585
R1394 B.n498 B.n497 585
R1395 B.n935 B.n934 585
R1396 B.n936 B.n935 585
R1397 B.n933 B.n503 585
R1398 B.n503 B.n502 585
R1399 B.n932 B.n931 585
R1400 B.n931 B.n930 585
R1401 B.n505 B.n504 585
R1402 B.n923 B.n505 585
R1403 B.n922 B.n921 585
R1404 B.n924 B.n922 585
R1405 B.n920 B.n510 585
R1406 B.n510 B.n509 585
R1407 B.n919 B.n918 585
R1408 B.n918 B.n917 585
R1409 B.n512 B.n511 585
R1410 B.n513 B.n512 585
R1411 B.n910 B.n909 585
R1412 B.n911 B.n910 585
R1413 B.n908 B.n518 585
R1414 B.n518 B.n517 585
R1415 B.n907 B.n906 585
R1416 B.n906 B.n905 585
R1417 B.n520 B.n519 585
R1418 B.n521 B.n520 585
R1419 B.n898 B.n897 585
R1420 B.n899 B.n898 585
R1421 B.n896 B.n526 585
R1422 B.n526 B.n525 585
R1423 B.n895 B.n894 585
R1424 B.n894 B.n893 585
R1425 B.n528 B.n527 585
R1426 B.n529 B.n528 585
R1427 B.n886 B.n885 585
R1428 B.n887 B.n886 585
R1429 B.n884 B.n534 585
R1430 B.n534 B.n533 585
R1431 B.n883 B.n882 585
R1432 B.n882 B.n881 585
R1433 B.n536 B.n535 585
R1434 B.n537 B.n536 585
R1435 B.n874 B.n873 585
R1436 B.n875 B.n874 585
R1437 B.n872 B.n542 585
R1438 B.n542 B.n541 585
R1439 B.n866 B.n865 585
R1440 B.n864 B.n608 585
R1441 B.n863 B.n607 585
R1442 B.n868 B.n607 585
R1443 B.n862 B.n861 585
R1444 B.n860 B.n859 585
R1445 B.n858 B.n857 585
R1446 B.n856 B.n855 585
R1447 B.n854 B.n853 585
R1448 B.n852 B.n851 585
R1449 B.n850 B.n849 585
R1450 B.n848 B.n847 585
R1451 B.n846 B.n845 585
R1452 B.n844 B.n843 585
R1453 B.n842 B.n841 585
R1454 B.n840 B.n839 585
R1455 B.n838 B.n837 585
R1456 B.n836 B.n835 585
R1457 B.n834 B.n833 585
R1458 B.n832 B.n831 585
R1459 B.n830 B.n829 585
R1460 B.n828 B.n827 585
R1461 B.n826 B.n825 585
R1462 B.n824 B.n823 585
R1463 B.n822 B.n821 585
R1464 B.n820 B.n819 585
R1465 B.n818 B.n817 585
R1466 B.n816 B.n815 585
R1467 B.n814 B.n813 585
R1468 B.n812 B.n811 585
R1469 B.n810 B.n809 585
R1470 B.n808 B.n807 585
R1471 B.n806 B.n805 585
R1472 B.n804 B.n803 585
R1473 B.n802 B.n801 585
R1474 B.n800 B.n799 585
R1475 B.n798 B.n797 585
R1476 B.n796 B.n795 585
R1477 B.n794 B.n793 585
R1478 B.n792 B.n791 585
R1479 B.n790 B.n789 585
R1480 B.n788 B.n787 585
R1481 B.n786 B.n785 585
R1482 B.n784 B.n783 585
R1483 B.n782 B.n781 585
R1484 B.n780 B.n779 585
R1485 B.n778 B.n777 585
R1486 B.n776 B.n775 585
R1487 B.n774 B.n773 585
R1488 B.n772 B.n771 585
R1489 B.n770 B.n769 585
R1490 B.n768 B.n767 585
R1491 B.n766 B.n765 585
R1492 B.n764 B.n763 585
R1493 B.n762 B.n761 585
R1494 B.n760 B.n759 585
R1495 B.n758 B.n757 585
R1496 B.n756 B.n755 585
R1497 B.n754 B.n753 585
R1498 B.n752 B.n751 585
R1499 B.n750 B.n749 585
R1500 B.n747 B.n746 585
R1501 B.n745 B.n744 585
R1502 B.n743 B.n742 585
R1503 B.n741 B.n740 585
R1504 B.n739 B.n738 585
R1505 B.n737 B.n736 585
R1506 B.n735 B.n734 585
R1507 B.n733 B.n732 585
R1508 B.n731 B.n730 585
R1509 B.n729 B.n728 585
R1510 B.n727 B.n726 585
R1511 B.n725 B.n724 585
R1512 B.n723 B.n722 585
R1513 B.n721 B.n720 585
R1514 B.n719 B.n718 585
R1515 B.n717 B.n716 585
R1516 B.n715 B.n714 585
R1517 B.n713 B.n712 585
R1518 B.n711 B.n710 585
R1519 B.n709 B.n708 585
R1520 B.n707 B.n706 585
R1521 B.n705 B.n704 585
R1522 B.n703 B.n702 585
R1523 B.n701 B.n700 585
R1524 B.n699 B.n698 585
R1525 B.n697 B.n696 585
R1526 B.n695 B.n694 585
R1527 B.n693 B.n692 585
R1528 B.n691 B.n690 585
R1529 B.n689 B.n688 585
R1530 B.n687 B.n686 585
R1531 B.n685 B.n684 585
R1532 B.n683 B.n682 585
R1533 B.n681 B.n680 585
R1534 B.n679 B.n678 585
R1535 B.n677 B.n676 585
R1536 B.n675 B.n674 585
R1537 B.n673 B.n672 585
R1538 B.n671 B.n670 585
R1539 B.n669 B.n668 585
R1540 B.n667 B.n666 585
R1541 B.n665 B.n664 585
R1542 B.n663 B.n662 585
R1543 B.n661 B.n660 585
R1544 B.n659 B.n658 585
R1545 B.n657 B.n656 585
R1546 B.n655 B.n654 585
R1547 B.n653 B.n652 585
R1548 B.n651 B.n650 585
R1549 B.n649 B.n648 585
R1550 B.n647 B.n646 585
R1551 B.n645 B.n644 585
R1552 B.n643 B.n642 585
R1553 B.n641 B.n640 585
R1554 B.n639 B.n638 585
R1555 B.n637 B.n636 585
R1556 B.n635 B.n634 585
R1557 B.n633 B.n632 585
R1558 B.n631 B.n630 585
R1559 B.n629 B.n628 585
R1560 B.n627 B.n626 585
R1561 B.n625 B.n624 585
R1562 B.n623 B.n622 585
R1563 B.n621 B.n620 585
R1564 B.n619 B.n618 585
R1565 B.n617 B.n616 585
R1566 B.n615 B.n614 585
R1567 B.n544 B.n543 585
R1568 B.n871 B.n870 585
R1569 B.n540 B.n539 585
R1570 B.n541 B.n540 585
R1571 B.n877 B.n876 585
R1572 B.n876 B.n875 585
R1573 B.n878 B.n538 585
R1574 B.n538 B.n537 585
R1575 B.n880 B.n879 585
R1576 B.n881 B.n880 585
R1577 B.n532 B.n531 585
R1578 B.n533 B.n532 585
R1579 B.n889 B.n888 585
R1580 B.n888 B.n887 585
R1581 B.n890 B.n530 585
R1582 B.n530 B.n529 585
R1583 B.n892 B.n891 585
R1584 B.n893 B.n892 585
R1585 B.n524 B.n523 585
R1586 B.n525 B.n524 585
R1587 B.n901 B.n900 585
R1588 B.n900 B.n899 585
R1589 B.n902 B.n522 585
R1590 B.n522 B.n521 585
R1591 B.n904 B.n903 585
R1592 B.n905 B.n904 585
R1593 B.n516 B.n515 585
R1594 B.n517 B.n516 585
R1595 B.n913 B.n912 585
R1596 B.n912 B.n911 585
R1597 B.n914 B.n514 585
R1598 B.n514 B.n513 585
R1599 B.n916 B.n915 585
R1600 B.n917 B.n916 585
R1601 B.n508 B.n507 585
R1602 B.n509 B.n508 585
R1603 B.n926 B.n925 585
R1604 B.n925 B.n924 585
R1605 B.n927 B.n506 585
R1606 B.n923 B.n506 585
R1607 B.n929 B.n928 585
R1608 B.n930 B.n929 585
R1609 B.n501 B.n500 585
R1610 B.n502 B.n501 585
R1611 B.n938 B.n937 585
R1612 B.n937 B.n936 585
R1613 B.n939 B.n499 585
R1614 B.n499 B.n498 585
R1615 B.n941 B.n940 585
R1616 B.n942 B.n941 585
R1617 B.n493 B.n492 585
R1618 B.n494 B.n493 585
R1619 B.n950 B.n949 585
R1620 B.n949 B.n948 585
R1621 B.n951 B.n491 585
R1622 B.n491 B.n490 585
R1623 B.n953 B.n952 585
R1624 B.n954 B.n953 585
R1625 B.n485 B.n484 585
R1626 B.n486 B.n485 585
R1627 B.n962 B.n961 585
R1628 B.n961 B.n960 585
R1629 B.n963 B.n483 585
R1630 B.n483 B.n482 585
R1631 B.n965 B.n964 585
R1632 B.n966 B.n965 585
R1633 B.n477 B.n476 585
R1634 B.n478 B.n477 585
R1635 B.n974 B.n973 585
R1636 B.n973 B.n972 585
R1637 B.n975 B.n475 585
R1638 B.n475 B.n474 585
R1639 B.n977 B.n976 585
R1640 B.n978 B.n977 585
R1641 B.n469 B.n468 585
R1642 B.n470 B.n469 585
R1643 B.n986 B.n985 585
R1644 B.n985 B.n984 585
R1645 B.n987 B.n467 585
R1646 B.n467 B.n466 585
R1647 B.n989 B.n988 585
R1648 B.n990 B.n989 585
R1649 B.n461 B.n460 585
R1650 B.n462 B.n461 585
R1651 B.n998 B.n997 585
R1652 B.n997 B.n996 585
R1653 B.n999 B.n459 585
R1654 B.n459 B.n458 585
R1655 B.n1001 B.n1000 585
R1656 B.n1002 B.n1001 585
R1657 B.n453 B.n452 585
R1658 B.n454 B.n453 585
R1659 B.n1010 B.n1009 585
R1660 B.n1009 B.n1008 585
R1661 B.n1011 B.n451 585
R1662 B.n451 B.n450 585
R1663 B.n1013 B.n1012 585
R1664 B.n1014 B.n1013 585
R1665 B.n445 B.n444 585
R1666 B.n446 B.n445 585
R1667 B.n1022 B.n1021 585
R1668 B.n1021 B.n1020 585
R1669 B.n1023 B.n443 585
R1670 B.n443 B.n442 585
R1671 B.n1025 B.n1024 585
R1672 B.n1026 B.n1025 585
R1673 B.n437 B.n436 585
R1674 B.n438 B.n437 585
R1675 B.n1035 B.n1034 585
R1676 B.n1034 B.n1033 585
R1677 B.n1036 B.n435 585
R1678 B.n435 B.n434 585
R1679 B.n1038 B.n1037 585
R1680 B.n1039 B.n1038 585
R1681 B.n3 B.n0 585
R1682 B.n4 B.n3 585
R1683 B.n1231 B.n1 585
R1684 B.n1232 B.n1231 585
R1685 B.n1230 B.n1229 585
R1686 B.n1230 B.n8 585
R1687 B.n1228 B.n9 585
R1688 B.n12 B.n9 585
R1689 B.n1227 B.n1226 585
R1690 B.n1226 B.n1225 585
R1691 B.n11 B.n10 585
R1692 B.n1224 B.n11 585
R1693 B.n1222 B.n1221 585
R1694 B.n1223 B.n1222 585
R1695 B.n1220 B.n17 585
R1696 B.n17 B.n16 585
R1697 B.n1219 B.n1218 585
R1698 B.n1218 B.n1217 585
R1699 B.n19 B.n18 585
R1700 B.n1216 B.n19 585
R1701 B.n1214 B.n1213 585
R1702 B.n1215 B.n1214 585
R1703 B.n1212 B.n24 585
R1704 B.n24 B.n23 585
R1705 B.n1211 B.n1210 585
R1706 B.n1210 B.n1209 585
R1707 B.n26 B.n25 585
R1708 B.n1208 B.n26 585
R1709 B.n1206 B.n1205 585
R1710 B.n1207 B.n1206 585
R1711 B.n1204 B.n31 585
R1712 B.n31 B.n30 585
R1713 B.n1203 B.n1202 585
R1714 B.n1202 B.n1201 585
R1715 B.n33 B.n32 585
R1716 B.n1200 B.n33 585
R1717 B.n1198 B.n1197 585
R1718 B.n1199 B.n1198 585
R1719 B.n1196 B.n38 585
R1720 B.n38 B.n37 585
R1721 B.n1195 B.n1194 585
R1722 B.n1194 B.n1193 585
R1723 B.n40 B.n39 585
R1724 B.n1192 B.n40 585
R1725 B.n1190 B.n1189 585
R1726 B.n1191 B.n1190 585
R1727 B.n1188 B.n45 585
R1728 B.n45 B.n44 585
R1729 B.n1187 B.n1186 585
R1730 B.n1186 B.n1185 585
R1731 B.n47 B.n46 585
R1732 B.n1184 B.n47 585
R1733 B.n1182 B.n1181 585
R1734 B.n1183 B.n1182 585
R1735 B.n1180 B.n52 585
R1736 B.n52 B.n51 585
R1737 B.n1179 B.n1178 585
R1738 B.n1178 B.n1177 585
R1739 B.n54 B.n53 585
R1740 B.n1176 B.n54 585
R1741 B.n1174 B.n1173 585
R1742 B.n1175 B.n1174 585
R1743 B.n1172 B.n59 585
R1744 B.n59 B.n58 585
R1745 B.n1171 B.n1170 585
R1746 B.n1170 B.n1169 585
R1747 B.n61 B.n60 585
R1748 B.n1168 B.n61 585
R1749 B.n1166 B.n1165 585
R1750 B.n1167 B.n1166 585
R1751 B.n1164 B.n66 585
R1752 B.n66 B.n65 585
R1753 B.n1163 B.n1162 585
R1754 B.n1162 B.n1161 585
R1755 B.n68 B.n67 585
R1756 B.n1160 B.n68 585
R1757 B.n1158 B.n1157 585
R1758 B.n1159 B.n1158 585
R1759 B.n1156 B.n72 585
R1760 B.n75 B.n72 585
R1761 B.n1155 B.n1154 585
R1762 B.n1154 B.n1153 585
R1763 B.n74 B.n73 585
R1764 B.n1152 B.n74 585
R1765 B.n1150 B.n1149 585
R1766 B.n1151 B.n1150 585
R1767 B.n1148 B.n80 585
R1768 B.n80 B.n79 585
R1769 B.n1147 B.n1146 585
R1770 B.n1146 B.n1145 585
R1771 B.n82 B.n81 585
R1772 B.n1144 B.n82 585
R1773 B.n1142 B.n1141 585
R1774 B.n1143 B.n1142 585
R1775 B.n1140 B.n87 585
R1776 B.n87 B.n86 585
R1777 B.n1139 B.n1138 585
R1778 B.n1138 B.n1137 585
R1779 B.n89 B.n88 585
R1780 B.n1136 B.n89 585
R1781 B.n1134 B.n1133 585
R1782 B.n1135 B.n1134 585
R1783 B.n1132 B.n94 585
R1784 B.n94 B.n93 585
R1785 B.n1131 B.n1130 585
R1786 B.n1130 B.n1129 585
R1787 B.n96 B.n95 585
R1788 B.n1128 B.n96 585
R1789 B.n1126 B.n1125 585
R1790 B.n1127 B.n1126 585
R1791 B.n1124 B.n101 585
R1792 B.n101 B.n100 585
R1793 B.n1123 B.n1122 585
R1794 B.n1122 B.n1121 585
R1795 B.n103 B.n102 585
R1796 B.n1120 B.n103 585
R1797 B.n1235 B.n1234 585
R1798 B.n1233 B.n2 585
R1799 B.n176 B.n103 444.452
R1800 B.n1118 B.n105 444.452
R1801 B.n870 B.n542 444.452
R1802 B.n866 B.n540 444.452
R1803 B.n173 B.t22 440.947
R1804 B.n171 B.t19 440.947
R1805 B.n611 B.t13 440.947
R1806 B.n609 B.t16 440.947
R1807 B.n172 B.t20 386.839
R1808 B.n612 B.t12 386.839
R1809 B.n174 B.t23 386.837
R1810 B.n610 B.t15 386.837
R1811 B.n173 B.t21 385.048
R1812 B.n171 B.t17 385.048
R1813 B.n611 B.t10 385.048
R1814 B.n609 B.t14 385.048
R1815 B.n1119 B.n169 256.663
R1816 B.n1119 B.n168 256.663
R1817 B.n1119 B.n167 256.663
R1818 B.n1119 B.n166 256.663
R1819 B.n1119 B.n165 256.663
R1820 B.n1119 B.n164 256.663
R1821 B.n1119 B.n163 256.663
R1822 B.n1119 B.n162 256.663
R1823 B.n1119 B.n161 256.663
R1824 B.n1119 B.n160 256.663
R1825 B.n1119 B.n159 256.663
R1826 B.n1119 B.n158 256.663
R1827 B.n1119 B.n157 256.663
R1828 B.n1119 B.n156 256.663
R1829 B.n1119 B.n155 256.663
R1830 B.n1119 B.n154 256.663
R1831 B.n1119 B.n153 256.663
R1832 B.n1119 B.n152 256.663
R1833 B.n1119 B.n151 256.663
R1834 B.n1119 B.n150 256.663
R1835 B.n1119 B.n149 256.663
R1836 B.n1119 B.n148 256.663
R1837 B.n1119 B.n147 256.663
R1838 B.n1119 B.n146 256.663
R1839 B.n1119 B.n145 256.663
R1840 B.n1119 B.n144 256.663
R1841 B.n1119 B.n143 256.663
R1842 B.n1119 B.n142 256.663
R1843 B.n1119 B.n141 256.663
R1844 B.n1119 B.n140 256.663
R1845 B.n1119 B.n139 256.663
R1846 B.n1119 B.n138 256.663
R1847 B.n1119 B.n137 256.663
R1848 B.n1119 B.n136 256.663
R1849 B.n1119 B.n135 256.663
R1850 B.n1119 B.n134 256.663
R1851 B.n1119 B.n133 256.663
R1852 B.n1119 B.n132 256.663
R1853 B.n1119 B.n131 256.663
R1854 B.n1119 B.n130 256.663
R1855 B.n1119 B.n129 256.663
R1856 B.n1119 B.n128 256.663
R1857 B.n1119 B.n127 256.663
R1858 B.n1119 B.n126 256.663
R1859 B.n1119 B.n125 256.663
R1860 B.n1119 B.n124 256.663
R1861 B.n1119 B.n123 256.663
R1862 B.n1119 B.n122 256.663
R1863 B.n1119 B.n121 256.663
R1864 B.n1119 B.n120 256.663
R1865 B.n1119 B.n119 256.663
R1866 B.n1119 B.n118 256.663
R1867 B.n1119 B.n117 256.663
R1868 B.n1119 B.n116 256.663
R1869 B.n1119 B.n115 256.663
R1870 B.n1119 B.n114 256.663
R1871 B.n1119 B.n113 256.663
R1872 B.n1119 B.n112 256.663
R1873 B.n1119 B.n111 256.663
R1874 B.n1119 B.n110 256.663
R1875 B.n1119 B.n109 256.663
R1876 B.n1119 B.n108 256.663
R1877 B.n1119 B.n107 256.663
R1878 B.n1119 B.n106 256.663
R1879 B.n868 B.n867 256.663
R1880 B.n868 B.n545 256.663
R1881 B.n868 B.n546 256.663
R1882 B.n868 B.n547 256.663
R1883 B.n868 B.n548 256.663
R1884 B.n868 B.n549 256.663
R1885 B.n868 B.n550 256.663
R1886 B.n868 B.n551 256.663
R1887 B.n868 B.n552 256.663
R1888 B.n868 B.n553 256.663
R1889 B.n868 B.n554 256.663
R1890 B.n868 B.n555 256.663
R1891 B.n868 B.n556 256.663
R1892 B.n868 B.n557 256.663
R1893 B.n868 B.n558 256.663
R1894 B.n868 B.n559 256.663
R1895 B.n868 B.n560 256.663
R1896 B.n868 B.n561 256.663
R1897 B.n868 B.n562 256.663
R1898 B.n868 B.n563 256.663
R1899 B.n868 B.n564 256.663
R1900 B.n868 B.n565 256.663
R1901 B.n868 B.n566 256.663
R1902 B.n868 B.n567 256.663
R1903 B.n868 B.n568 256.663
R1904 B.n868 B.n569 256.663
R1905 B.n868 B.n570 256.663
R1906 B.n868 B.n571 256.663
R1907 B.n868 B.n572 256.663
R1908 B.n868 B.n573 256.663
R1909 B.n868 B.n574 256.663
R1910 B.n868 B.n575 256.663
R1911 B.n868 B.n576 256.663
R1912 B.n868 B.n577 256.663
R1913 B.n868 B.n578 256.663
R1914 B.n868 B.n579 256.663
R1915 B.n868 B.n580 256.663
R1916 B.n868 B.n581 256.663
R1917 B.n868 B.n582 256.663
R1918 B.n868 B.n583 256.663
R1919 B.n868 B.n584 256.663
R1920 B.n868 B.n585 256.663
R1921 B.n868 B.n586 256.663
R1922 B.n868 B.n587 256.663
R1923 B.n868 B.n588 256.663
R1924 B.n868 B.n589 256.663
R1925 B.n868 B.n590 256.663
R1926 B.n868 B.n591 256.663
R1927 B.n868 B.n592 256.663
R1928 B.n868 B.n593 256.663
R1929 B.n868 B.n594 256.663
R1930 B.n868 B.n595 256.663
R1931 B.n868 B.n596 256.663
R1932 B.n868 B.n597 256.663
R1933 B.n868 B.n598 256.663
R1934 B.n868 B.n599 256.663
R1935 B.n868 B.n600 256.663
R1936 B.n868 B.n601 256.663
R1937 B.n868 B.n602 256.663
R1938 B.n868 B.n603 256.663
R1939 B.n868 B.n604 256.663
R1940 B.n868 B.n605 256.663
R1941 B.n868 B.n606 256.663
R1942 B.n869 B.n868 256.663
R1943 B.n1237 B.n1236 256.663
R1944 B.n180 B.n179 163.367
R1945 B.n184 B.n183 163.367
R1946 B.n188 B.n187 163.367
R1947 B.n192 B.n191 163.367
R1948 B.n196 B.n195 163.367
R1949 B.n200 B.n199 163.367
R1950 B.n204 B.n203 163.367
R1951 B.n208 B.n207 163.367
R1952 B.n212 B.n211 163.367
R1953 B.n216 B.n215 163.367
R1954 B.n220 B.n219 163.367
R1955 B.n224 B.n223 163.367
R1956 B.n228 B.n227 163.367
R1957 B.n232 B.n231 163.367
R1958 B.n236 B.n235 163.367
R1959 B.n240 B.n239 163.367
R1960 B.n244 B.n243 163.367
R1961 B.n248 B.n247 163.367
R1962 B.n252 B.n251 163.367
R1963 B.n256 B.n255 163.367
R1964 B.n260 B.n259 163.367
R1965 B.n264 B.n263 163.367
R1966 B.n268 B.n267 163.367
R1967 B.n272 B.n271 163.367
R1968 B.n276 B.n275 163.367
R1969 B.n280 B.n279 163.367
R1970 B.n284 B.n283 163.367
R1971 B.n288 B.n287 163.367
R1972 B.n292 B.n291 163.367
R1973 B.n296 B.n295 163.367
R1974 B.n300 B.n299 163.367
R1975 B.n304 B.n303 163.367
R1976 B.n308 B.n307 163.367
R1977 B.n312 B.n311 163.367
R1978 B.n317 B.n316 163.367
R1979 B.n321 B.n320 163.367
R1980 B.n325 B.n324 163.367
R1981 B.n329 B.n328 163.367
R1982 B.n333 B.n332 163.367
R1983 B.n337 B.n336 163.367
R1984 B.n341 B.n340 163.367
R1985 B.n345 B.n344 163.367
R1986 B.n349 B.n348 163.367
R1987 B.n353 B.n352 163.367
R1988 B.n357 B.n356 163.367
R1989 B.n361 B.n360 163.367
R1990 B.n365 B.n364 163.367
R1991 B.n369 B.n368 163.367
R1992 B.n373 B.n372 163.367
R1993 B.n377 B.n376 163.367
R1994 B.n381 B.n380 163.367
R1995 B.n385 B.n384 163.367
R1996 B.n389 B.n388 163.367
R1997 B.n393 B.n392 163.367
R1998 B.n397 B.n396 163.367
R1999 B.n401 B.n400 163.367
R2000 B.n405 B.n404 163.367
R2001 B.n409 B.n408 163.367
R2002 B.n413 B.n412 163.367
R2003 B.n417 B.n416 163.367
R2004 B.n421 B.n420 163.367
R2005 B.n425 B.n424 163.367
R2006 B.n429 B.n428 163.367
R2007 B.n1118 B.n170 163.367
R2008 B.n874 B.n542 163.367
R2009 B.n874 B.n536 163.367
R2010 B.n882 B.n536 163.367
R2011 B.n882 B.n534 163.367
R2012 B.n886 B.n534 163.367
R2013 B.n886 B.n528 163.367
R2014 B.n894 B.n528 163.367
R2015 B.n894 B.n526 163.367
R2016 B.n898 B.n526 163.367
R2017 B.n898 B.n520 163.367
R2018 B.n906 B.n520 163.367
R2019 B.n906 B.n518 163.367
R2020 B.n910 B.n518 163.367
R2021 B.n910 B.n512 163.367
R2022 B.n918 B.n512 163.367
R2023 B.n918 B.n510 163.367
R2024 B.n922 B.n510 163.367
R2025 B.n922 B.n505 163.367
R2026 B.n931 B.n505 163.367
R2027 B.n931 B.n503 163.367
R2028 B.n935 B.n503 163.367
R2029 B.n935 B.n497 163.367
R2030 B.n943 B.n497 163.367
R2031 B.n943 B.n495 163.367
R2032 B.n947 B.n495 163.367
R2033 B.n947 B.n489 163.367
R2034 B.n955 B.n489 163.367
R2035 B.n955 B.n487 163.367
R2036 B.n959 B.n487 163.367
R2037 B.n959 B.n481 163.367
R2038 B.n967 B.n481 163.367
R2039 B.n967 B.n479 163.367
R2040 B.n971 B.n479 163.367
R2041 B.n971 B.n473 163.367
R2042 B.n979 B.n473 163.367
R2043 B.n979 B.n471 163.367
R2044 B.n983 B.n471 163.367
R2045 B.n983 B.n465 163.367
R2046 B.n991 B.n465 163.367
R2047 B.n991 B.n463 163.367
R2048 B.n995 B.n463 163.367
R2049 B.n995 B.n457 163.367
R2050 B.n1003 B.n457 163.367
R2051 B.n1003 B.n455 163.367
R2052 B.n1007 B.n455 163.367
R2053 B.n1007 B.n449 163.367
R2054 B.n1015 B.n449 163.367
R2055 B.n1015 B.n447 163.367
R2056 B.n1019 B.n447 163.367
R2057 B.n1019 B.n441 163.367
R2058 B.n1027 B.n441 163.367
R2059 B.n1027 B.n439 163.367
R2060 B.n1032 B.n439 163.367
R2061 B.n1032 B.n433 163.367
R2062 B.n1040 B.n433 163.367
R2063 B.n1041 B.n1040 163.367
R2064 B.n1041 B.n5 163.367
R2065 B.n6 B.n5 163.367
R2066 B.n7 B.n6 163.367
R2067 B.n1047 B.n7 163.367
R2068 B.n1048 B.n1047 163.367
R2069 B.n1048 B.n13 163.367
R2070 B.n14 B.n13 163.367
R2071 B.n15 B.n14 163.367
R2072 B.n1053 B.n15 163.367
R2073 B.n1053 B.n20 163.367
R2074 B.n21 B.n20 163.367
R2075 B.n22 B.n21 163.367
R2076 B.n1058 B.n22 163.367
R2077 B.n1058 B.n27 163.367
R2078 B.n28 B.n27 163.367
R2079 B.n29 B.n28 163.367
R2080 B.n1063 B.n29 163.367
R2081 B.n1063 B.n34 163.367
R2082 B.n35 B.n34 163.367
R2083 B.n36 B.n35 163.367
R2084 B.n1068 B.n36 163.367
R2085 B.n1068 B.n41 163.367
R2086 B.n42 B.n41 163.367
R2087 B.n43 B.n42 163.367
R2088 B.n1073 B.n43 163.367
R2089 B.n1073 B.n48 163.367
R2090 B.n49 B.n48 163.367
R2091 B.n50 B.n49 163.367
R2092 B.n1078 B.n50 163.367
R2093 B.n1078 B.n55 163.367
R2094 B.n56 B.n55 163.367
R2095 B.n57 B.n56 163.367
R2096 B.n1083 B.n57 163.367
R2097 B.n1083 B.n62 163.367
R2098 B.n63 B.n62 163.367
R2099 B.n64 B.n63 163.367
R2100 B.n1088 B.n64 163.367
R2101 B.n1088 B.n69 163.367
R2102 B.n70 B.n69 163.367
R2103 B.n71 B.n70 163.367
R2104 B.n1093 B.n71 163.367
R2105 B.n1093 B.n76 163.367
R2106 B.n77 B.n76 163.367
R2107 B.n78 B.n77 163.367
R2108 B.n1098 B.n78 163.367
R2109 B.n1098 B.n83 163.367
R2110 B.n84 B.n83 163.367
R2111 B.n85 B.n84 163.367
R2112 B.n1103 B.n85 163.367
R2113 B.n1103 B.n90 163.367
R2114 B.n91 B.n90 163.367
R2115 B.n92 B.n91 163.367
R2116 B.n1108 B.n92 163.367
R2117 B.n1108 B.n97 163.367
R2118 B.n98 B.n97 163.367
R2119 B.n99 B.n98 163.367
R2120 B.n1113 B.n99 163.367
R2121 B.n1113 B.n104 163.367
R2122 B.n105 B.n104 163.367
R2123 B.n608 B.n607 163.367
R2124 B.n861 B.n607 163.367
R2125 B.n859 B.n858 163.367
R2126 B.n855 B.n854 163.367
R2127 B.n851 B.n850 163.367
R2128 B.n847 B.n846 163.367
R2129 B.n843 B.n842 163.367
R2130 B.n839 B.n838 163.367
R2131 B.n835 B.n834 163.367
R2132 B.n831 B.n830 163.367
R2133 B.n827 B.n826 163.367
R2134 B.n823 B.n822 163.367
R2135 B.n819 B.n818 163.367
R2136 B.n815 B.n814 163.367
R2137 B.n811 B.n810 163.367
R2138 B.n807 B.n806 163.367
R2139 B.n803 B.n802 163.367
R2140 B.n799 B.n798 163.367
R2141 B.n795 B.n794 163.367
R2142 B.n791 B.n790 163.367
R2143 B.n787 B.n786 163.367
R2144 B.n783 B.n782 163.367
R2145 B.n779 B.n778 163.367
R2146 B.n775 B.n774 163.367
R2147 B.n771 B.n770 163.367
R2148 B.n767 B.n766 163.367
R2149 B.n763 B.n762 163.367
R2150 B.n759 B.n758 163.367
R2151 B.n755 B.n754 163.367
R2152 B.n751 B.n750 163.367
R2153 B.n746 B.n745 163.367
R2154 B.n742 B.n741 163.367
R2155 B.n738 B.n737 163.367
R2156 B.n734 B.n733 163.367
R2157 B.n730 B.n729 163.367
R2158 B.n726 B.n725 163.367
R2159 B.n722 B.n721 163.367
R2160 B.n718 B.n717 163.367
R2161 B.n714 B.n713 163.367
R2162 B.n710 B.n709 163.367
R2163 B.n706 B.n705 163.367
R2164 B.n702 B.n701 163.367
R2165 B.n698 B.n697 163.367
R2166 B.n694 B.n693 163.367
R2167 B.n690 B.n689 163.367
R2168 B.n686 B.n685 163.367
R2169 B.n682 B.n681 163.367
R2170 B.n678 B.n677 163.367
R2171 B.n674 B.n673 163.367
R2172 B.n670 B.n669 163.367
R2173 B.n666 B.n665 163.367
R2174 B.n662 B.n661 163.367
R2175 B.n658 B.n657 163.367
R2176 B.n654 B.n653 163.367
R2177 B.n650 B.n649 163.367
R2178 B.n646 B.n645 163.367
R2179 B.n642 B.n641 163.367
R2180 B.n638 B.n637 163.367
R2181 B.n634 B.n633 163.367
R2182 B.n630 B.n629 163.367
R2183 B.n626 B.n625 163.367
R2184 B.n622 B.n621 163.367
R2185 B.n618 B.n617 163.367
R2186 B.n614 B.n544 163.367
R2187 B.n876 B.n540 163.367
R2188 B.n876 B.n538 163.367
R2189 B.n880 B.n538 163.367
R2190 B.n880 B.n532 163.367
R2191 B.n888 B.n532 163.367
R2192 B.n888 B.n530 163.367
R2193 B.n892 B.n530 163.367
R2194 B.n892 B.n524 163.367
R2195 B.n900 B.n524 163.367
R2196 B.n900 B.n522 163.367
R2197 B.n904 B.n522 163.367
R2198 B.n904 B.n516 163.367
R2199 B.n912 B.n516 163.367
R2200 B.n912 B.n514 163.367
R2201 B.n916 B.n514 163.367
R2202 B.n916 B.n508 163.367
R2203 B.n925 B.n508 163.367
R2204 B.n925 B.n506 163.367
R2205 B.n929 B.n506 163.367
R2206 B.n929 B.n501 163.367
R2207 B.n937 B.n501 163.367
R2208 B.n937 B.n499 163.367
R2209 B.n941 B.n499 163.367
R2210 B.n941 B.n493 163.367
R2211 B.n949 B.n493 163.367
R2212 B.n949 B.n491 163.367
R2213 B.n953 B.n491 163.367
R2214 B.n953 B.n485 163.367
R2215 B.n961 B.n485 163.367
R2216 B.n961 B.n483 163.367
R2217 B.n965 B.n483 163.367
R2218 B.n965 B.n477 163.367
R2219 B.n973 B.n477 163.367
R2220 B.n973 B.n475 163.367
R2221 B.n977 B.n475 163.367
R2222 B.n977 B.n469 163.367
R2223 B.n985 B.n469 163.367
R2224 B.n985 B.n467 163.367
R2225 B.n989 B.n467 163.367
R2226 B.n989 B.n461 163.367
R2227 B.n997 B.n461 163.367
R2228 B.n997 B.n459 163.367
R2229 B.n1001 B.n459 163.367
R2230 B.n1001 B.n453 163.367
R2231 B.n1009 B.n453 163.367
R2232 B.n1009 B.n451 163.367
R2233 B.n1013 B.n451 163.367
R2234 B.n1013 B.n445 163.367
R2235 B.n1021 B.n445 163.367
R2236 B.n1021 B.n443 163.367
R2237 B.n1025 B.n443 163.367
R2238 B.n1025 B.n437 163.367
R2239 B.n1034 B.n437 163.367
R2240 B.n1034 B.n435 163.367
R2241 B.n1038 B.n435 163.367
R2242 B.n1038 B.n3 163.367
R2243 B.n1235 B.n3 163.367
R2244 B.n1231 B.n2 163.367
R2245 B.n1231 B.n1230 163.367
R2246 B.n1230 B.n9 163.367
R2247 B.n1226 B.n9 163.367
R2248 B.n1226 B.n11 163.367
R2249 B.n1222 B.n11 163.367
R2250 B.n1222 B.n17 163.367
R2251 B.n1218 B.n17 163.367
R2252 B.n1218 B.n19 163.367
R2253 B.n1214 B.n19 163.367
R2254 B.n1214 B.n24 163.367
R2255 B.n1210 B.n24 163.367
R2256 B.n1210 B.n26 163.367
R2257 B.n1206 B.n26 163.367
R2258 B.n1206 B.n31 163.367
R2259 B.n1202 B.n31 163.367
R2260 B.n1202 B.n33 163.367
R2261 B.n1198 B.n33 163.367
R2262 B.n1198 B.n38 163.367
R2263 B.n1194 B.n38 163.367
R2264 B.n1194 B.n40 163.367
R2265 B.n1190 B.n40 163.367
R2266 B.n1190 B.n45 163.367
R2267 B.n1186 B.n45 163.367
R2268 B.n1186 B.n47 163.367
R2269 B.n1182 B.n47 163.367
R2270 B.n1182 B.n52 163.367
R2271 B.n1178 B.n52 163.367
R2272 B.n1178 B.n54 163.367
R2273 B.n1174 B.n54 163.367
R2274 B.n1174 B.n59 163.367
R2275 B.n1170 B.n59 163.367
R2276 B.n1170 B.n61 163.367
R2277 B.n1166 B.n61 163.367
R2278 B.n1166 B.n66 163.367
R2279 B.n1162 B.n66 163.367
R2280 B.n1162 B.n68 163.367
R2281 B.n1158 B.n68 163.367
R2282 B.n1158 B.n72 163.367
R2283 B.n1154 B.n72 163.367
R2284 B.n1154 B.n74 163.367
R2285 B.n1150 B.n74 163.367
R2286 B.n1150 B.n80 163.367
R2287 B.n1146 B.n80 163.367
R2288 B.n1146 B.n82 163.367
R2289 B.n1142 B.n82 163.367
R2290 B.n1142 B.n87 163.367
R2291 B.n1138 B.n87 163.367
R2292 B.n1138 B.n89 163.367
R2293 B.n1134 B.n89 163.367
R2294 B.n1134 B.n94 163.367
R2295 B.n1130 B.n94 163.367
R2296 B.n1130 B.n96 163.367
R2297 B.n1126 B.n96 163.367
R2298 B.n1126 B.n101 163.367
R2299 B.n1122 B.n101 163.367
R2300 B.n1122 B.n103 163.367
R2301 B.n176 B.n106 71.676
R2302 B.n180 B.n107 71.676
R2303 B.n184 B.n108 71.676
R2304 B.n188 B.n109 71.676
R2305 B.n192 B.n110 71.676
R2306 B.n196 B.n111 71.676
R2307 B.n200 B.n112 71.676
R2308 B.n204 B.n113 71.676
R2309 B.n208 B.n114 71.676
R2310 B.n212 B.n115 71.676
R2311 B.n216 B.n116 71.676
R2312 B.n220 B.n117 71.676
R2313 B.n224 B.n118 71.676
R2314 B.n228 B.n119 71.676
R2315 B.n232 B.n120 71.676
R2316 B.n236 B.n121 71.676
R2317 B.n240 B.n122 71.676
R2318 B.n244 B.n123 71.676
R2319 B.n248 B.n124 71.676
R2320 B.n252 B.n125 71.676
R2321 B.n256 B.n126 71.676
R2322 B.n260 B.n127 71.676
R2323 B.n264 B.n128 71.676
R2324 B.n268 B.n129 71.676
R2325 B.n272 B.n130 71.676
R2326 B.n276 B.n131 71.676
R2327 B.n280 B.n132 71.676
R2328 B.n284 B.n133 71.676
R2329 B.n288 B.n134 71.676
R2330 B.n292 B.n135 71.676
R2331 B.n296 B.n136 71.676
R2332 B.n300 B.n137 71.676
R2333 B.n304 B.n138 71.676
R2334 B.n308 B.n139 71.676
R2335 B.n312 B.n140 71.676
R2336 B.n317 B.n141 71.676
R2337 B.n321 B.n142 71.676
R2338 B.n325 B.n143 71.676
R2339 B.n329 B.n144 71.676
R2340 B.n333 B.n145 71.676
R2341 B.n337 B.n146 71.676
R2342 B.n341 B.n147 71.676
R2343 B.n345 B.n148 71.676
R2344 B.n349 B.n149 71.676
R2345 B.n353 B.n150 71.676
R2346 B.n357 B.n151 71.676
R2347 B.n361 B.n152 71.676
R2348 B.n365 B.n153 71.676
R2349 B.n369 B.n154 71.676
R2350 B.n373 B.n155 71.676
R2351 B.n377 B.n156 71.676
R2352 B.n381 B.n157 71.676
R2353 B.n385 B.n158 71.676
R2354 B.n389 B.n159 71.676
R2355 B.n393 B.n160 71.676
R2356 B.n397 B.n161 71.676
R2357 B.n401 B.n162 71.676
R2358 B.n405 B.n163 71.676
R2359 B.n409 B.n164 71.676
R2360 B.n413 B.n165 71.676
R2361 B.n417 B.n166 71.676
R2362 B.n421 B.n167 71.676
R2363 B.n425 B.n168 71.676
R2364 B.n429 B.n169 71.676
R2365 B.n170 B.n169 71.676
R2366 B.n428 B.n168 71.676
R2367 B.n424 B.n167 71.676
R2368 B.n420 B.n166 71.676
R2369 B.n416 B.n165 71.676
R2370 B.n412 B.n164 71.676
R2371 B.n408 B.n163 71.676
R2372 B.n404 B.n162 71.676
R2373 B.n400 B.n161 71.676
R2374 B.n396 B.n160 71.676
R2375 B.n392 B.n159 71.676
R2376 B.n388 B.n158 71.676
R2377 B.n384 B.n157 71.676
R2378 B.n380 B.n156 71.676
R2379 B.n376 B.n155 71.676
R2380 B.n372 B.n154 71.676
R2381 B.n368 B.n153 71.676
R2382 B.n364 B.n152 71.676
R2383 B.n360 B.n151 71.676
R2384 B.n356 B.n150 71.676
R2385 B.n352 B.n149 71.676
R2386 B.n348 B.n148 71.676
R2387 B.n344 B.n147 71.676
R2388 B.n340 B.n146 71.676
R2389 B.n336 B.n145 71.676
R2390 B.n332 B.n144 71.676
R2391 B.n328 B.n143 71.676
R2392 B.n324 B.n142 71.676
R2393 B.n320 B.n141 71.676
R2394 B.n316 B.n140 71.676
R2395 B.n311 B.n139 71.676
R2396 B.n307 B.n138 71.676
R2397 B.n303 B.n137 71.676
R2398 B.n299 B.n136 71.676
R2399 B.n295 B.n135 71.676
R2400 B.n291 B.n134 71.676
R2401 B.n287 B.n133 71.676
R2402 B.n283 B.n132 71.676
R2403 B.n279 B.n131 71.676
R2404 B.n275 B.n130 71.676
R2405 B.n271 B.n129 71.676
R2406 B.n267 B.n128 71.676
R2407 B.n263 B.n127 71.676
R2408 B.n259 B.n126 71.676
R2409 B.n255 B.n125 71.676
R2410 B.n251 B.n124 71.676
R2411 B.n247 B.n123 71.676
R2412 B.n243 B.n122 71.676
R2413 B.n239 B.n121 71.676
R2414 B.n235 B.n120 71.676
R2415 B.n231 B.n119 71.676
R2416 B.n227 B.n118 71.676
R2417 B.n223 B.n117 71.676
R2418 B.n219 B.n116 71.676
R2419 B.n215 B.n115 71.676
R2420 B.n211 B.n114 71.676
R2421 B.n207 B.n113 71.676
R2422 B.n203 B.n112 71.676
R2423 B.n199 B.n111 71.676
R2424 B.n195 B.n110 71.676
R2425 B.n191 B.n109 71.676
R2426 B.n187 B.n108 71.676
R2427 B.n183 B.n107 71.676
R2428 B.n179 B.n106 71.676
R2429 B.n867 B.n866 71.676
R2430 B.n861 B.n545 71.676
R2431 B.n858 B.n546 71.676
R2432 B.n854 B.n547 71.676
R2433 B.n850 B.n548 71.676
R2434 B.n846 B.n549 71.676
R2435 B.n842 B.n550 71.676
R2436 B.n838 B.n551 71.676
R2437 B.n834 B.n552 71.676
R2438 B.n830 B.n553 71.676
R2439 B.n826 B.n554 71.676
R2440 B.n822 B.n555 71.676
R2441 B.n818 B.n556 71.676
R2442 B.n814 B.n557 71.676
R2443 B.n810 B.n558 71.676
R2444 B.n806 B.n559 71.676
R2445 B.n802 B.n560 71.676
R2446 B.n798 B.n561 71.676
R2447 B.n794 B.n562 71.676
R2448 B.n790 B.n563 71.676
R2449 B.n786 B.n564 71.676
R2450 B.n782 B.n565 71.676
R2451 B.n778 B.n566 71.676
R2452 B.n774 B.n567 71.676
R2453 B.n770 B.n568 71.676
R2454 B.n766 B.n569 71.676
R2455 B.n762 B.n570 71.676
R2456 B.n758 B.n571 71.676
R2457 B.n754 B.n572 71.676
R2458 B.n750 B.n573 71.676
R2459 B.n745 B.n574 71.676
R2460 B.n741 B.n575 71.676
R2461 B.n737 B.n576 71.676
R2462 B.n733 B.n577 71.676
R2463 B.n729 B.n578 71.676
R2464 B.n725 B.n579 71.676
R2465 B.n721 B.n580 71.676
R2466 B.n717 B.n581 71.676
R2467 B.n713 B.n582 71.676
R2468 B.n709 B.n583 71.676
R2469 B.n705 B.n584 71.676
R2470 B.n701 B.n585 71.676
R2471 B.n697 B.n586 71.676
R2472 B.n693 B.n587 71.676
R2473 B.n689 B.n588 71.676
R2474 B.n685 B.n589 71.676
R2475 B.n681 B.n590 71.676
R2476 B.n677 B.n591 71.676
R2477 B.n673 B.n592 71.676
R2478 B.n669 B.n593 71.676
R2479 B.n665 B.n594 71.676
R2480 B.n661 B.n595 71.676
R2481 B.n657 B.n596 71.676
R2482 B.n653 B.n597 71.676
R2483 B.n649 B.n598 71.676
R2484 B.n645 B.n599 71.676
R2485 B.n641 B.n600 71.676
R2486 B.n637 B.n601 71.676
R2487 B.n633 B.n602 71.676
R2488 B.n629 B.n603 71.676
R2489 B.n625 B.n604 71.676
R2490 B.n621 B.n605 71.676
R2491 B.n617 B.n606 71.676
R2492 B.n869 B.n544 71.676
R2493 B.n867 B.n608 71.676
R2494 B.n859 B.n545 71.676
R2495 B.n855 B.n546 71.676
R2496 B.n851 B.n547 71.676
R2497 B.n847 B.n548 71.676
R2498 B.n843 B.n549 71.676
R2499 B.n839 B.n550 71.676
R2500 B.n835 B.n551 71.676
R2501 B.n831 B.n552 71.676
R2502 B.n827 B.n553 71.676
R2503 B.n823 B.n554 71.676
R2504 B.n819 B.n555 71.676
R2505 B.n815 B.n556 71.676
R2506 B.n811 B.n557 71.676
R2507 B.n807 B.n558 71.676
R2508 B.n803 B.n559 71.676
R2509 B.n799 B.n560 71.676
R2510 B.n795 B.n561 71.676
R2511 B.n791 B.n562 71.676
R2512 B.n787 B.n563 71.676
R2513 B.n783 B.n564 71.676
R2514 B.n779 B.n565 71.676
R2515 B.n775 B.n566 71.676
R2516 B.n771 B.n567 71.676
R2517 B.n767 B.n568 71.676
R2518 B.n763 B.n569 71.676
R2519 B.n759 B.n570 71.676
R2520 B.n755 B.n571 71.676
R2521 B.n751 B.n572 71.676
R2522 B.n746 B.n573 71.676
R2523 B.n742 B.n574 71.676
R2524 B.n738 B.n575 71.676
R2525 B.n734 B.n576 71.676
R2526 B.n730 B.n577 71.676
R2527 B.n726 B.n578 71.676
R2528 B.n722 B.n579 71.676
R2529 B.n718 B.n580 71.676
R2530 B.n714 B.n581 71.676
R2531 B.n710 B.n582 71.676
R2532 B.n706 B.n583 71.676
R2533 B.n702 B.n584 71.676
R2534 B.n698 B.n585 71.676
R2535 B.n694 B.n586 71.676
R2536 B.n690 B.n587 71.676
R2537 B.n686 B.n588 71.676
R2538 B.n682 B.n589 71.676
R2539 B.n678 B.n590 71.676
R2540 B.n674 B.n591 71.676
R2541 B.n670 B.n592 71.676
R2542 B.n666 B.n593 71.676
R2543 B.n662 B.n594 71.676
R2544 B.n658 B.n595 71.676
R2545 B.n654 B.n596 71.676
R2546 B.n650 B.n597 71.676
R2547 B.n646 B.n598 71.676
R2548 B.n642 B.n599 71.676
R2549 B.n638 B.n600 71.676
R2550 B.n634 B.n601 71.676
R2551 B.n630 B.n602 71.676
R2552 B.n626 B.n603 71.676
R2553 B.n622 B.n604 71.676
R2554 B.n618 B.n605 71.676
R2555 B.n614 B.n606 71.676
R2556 B.n870 B.n869 71.676
R2557 B.n1236 B.n1235 71.676
R2558 B.n1236 B.n2 71.676
R2559 B.n175 B.n174 59.5399
R2560 B.n314 B.n172 59.5399
R2561 B.n613 B.n612 59.5399
R2562 B.n748 B.n610 59.5399
R2563 B.n174 B.n173 54.1096
R2564 B.n172 B.n171 54.1096
R2565 B.n612 B.n611 54.1096
R2566 B.n610 B.n609 54.1096
R2567 B.n868 B.n541 53.1997
R2568 B.n1120 B.n1119 53.1997
R2569 B.n875 B.n541 32.0142
R2570 B.n875 B.n537 32.0142
R2571 B.n881 B.n537 32.0142
R2572 B.n881 B.n533 32.0142
R2573 B.n887 B.n533 32.0142
R2574 B.n887 B.n529 32.0142
R2575 B.n893 B.n529 32.0142
R2576 B.n899 B.n525 32.0142
R2577 B.n899 B.n521 32.0142
R2578 B.n905 B.n521 32.0142
R2579 B.n905 B.n517 32.0142
R2580 B.n911 B.n517 32.0142
R2581 B.n911 B.n513 32.0142
R2582 B.n917 B.n513 32.0142
R2583 B.n917 B.n509 32.0142
R2584 B.n924 B.n509 32.0142
R2585 B.n924 B.n923 32.0142
R2586 B.n930 B.n502 32.0142
R2587 B.n936 B.n502 32.0142
R2588 B.n936 B.n498 32.0142
R2589 B.n942 B.n498 32.0142
R2590 B.n942 B.n494 32.0142
R2591 B.n948 B.n494 32.0142
R2592 B.n948 B.n490 32.0142
R2593 B.n954 B.n490 32.0142
R2594 B.n960 B.n486 32.0142
R2595 B.n960 B.n482 32.0142
R2596 B.n966 B.n482 32.0142
R2597 B.n966 B.n478 32.0142
R2598 B.n972 B.n478 32.0142
R2599 B.n972 B.n474 32.0142
R2600 B.n978 B.n474 32.0142
R2601 B.n984 B.n470 32.0142
R2602 B.n984 B.n466 32.0142
R2603 B.n990 B.n466 32.0142
R2604 B.n990 B.n462 32.0142
R2605 B.n996 B.n462 32.0142
R2606 B.n996 B.n458 32.0142
R2607 B.n1002 B.n458 32.0142
R2608 B.n1008 B.n454 32.0142
R2609 B.n1008 B.n450 32.0142
R2610 B.n1014 B.n450 32.0142
R2611 B.n1014 B.n446 32.0142
R2612 B.n1020 B.n446 32.0142
R2613 B.n1020 B.n442 32.0142
R2614 B.n1026 B.n442 32.0142
R2615 B.n1033 B.n438 32.0142
R2616 B.n1033 B.n434 32.0142
R2617 B.n1039 B.n434 32.0142
R2618 B.n1039 B.n4 32.0142
R2619 B.n1234 B.n4 32.0142
R2620 B.n1234 B.n1233 32.0142
R2621 B.n1233 B.n1232 32.0142
R2622 B.n1232 B.n8 32.0142
R2623 B.n12 B.n8 32.0142
R2624 B.n1225 B.n12 32.0142
R2625 B.n1225 B.n1224 32.0142
R2626 B.n1223 B.n16 32.0142
R2627 B.n1217 B.n16 32.0142
R2628 B.n1217 B.n1216 32.0142
R2629 B.n1216 B.n1215 32.0142
R2630 B.n1215 B.n23 32.0142
R2631 B.n1209 B.n23 32.0142
R2632 B.n1209 B.n1208 32.0142
R2633 B.n1207 B.n30 32.0142
R2634 B.n1201 B.n30 32.0142
R2635 B.n1201 B.n1200 32.0142
R2636 B.n1200 B.n1199 32.0142
R2637 B.n1199 B.n37 32.0142
R2638 B.n1193 B.n37 32.0142
R2639 B.n1193 B.n1192 32.0142
R2640 B.n1191 B.n44 32.0142
R2641 B.n1185 B.n44 32.0142
R2642 B.n1185 B.n1184 32.0142
R2643 B.n1184 B.n1183 32.0142
R2644 B.n1183 B.n51 32.0142
R2645 B.n1177 B.n51 32.0142
R2646 B.n1177 B.n1176 32.0142
R2647 B.n1175 B.n58 32.0142
R2648 B.n1169 B.n58 32.0142
R2649 B.n1169 B.n1168 32.0142
R2650 B.n1168 B.n1167 32.0142
R2651 B.n1167 B.n65 32.0142
R2652 B.n1161 B.n65 32.0142
R2653 B.n1161 B.n1160 32.0142
R2654 B.n1160 B.n1159 32.0142
R2655 B.n1153 B.n75 32.0142
R2656 B.n1153 B.n1152 32.0142
R2657 B.n1152 B.n1151 32.0142
R2658 B.n1151 B.n79 32.0142
R2659 B.n1145 B.n79 32.0142
R2660 B.n1145 B.n1144 32.0142
R2661 B.n1144 B.n1143 32.0142
R2662 B.n1143 B.n86 32.0142
R2663 B.n1137 B.n86 32.0142
R2664 B.n1137 B.n1136 32.0142
R2665 B.n1135 B.n93 32.0142
R2666 B.n1129 B.n93 32.0142
R2667 B.n1129 B.n1128 32.0142
R2668 B.n1128 B.n1127 32.0142
R2669 B.n1127 B.n100 32.0142
R2670 B.n1121 B.n100 32.0142
R2671 B.n1121 B.n1120 32.0142
R2672 B.n923 B.t0 31.0726
R2673 B.n75 B.t2 31.0726
R2674 B.n865 B.n539 28.8785
R2675 B.n872 B.n871 28.8785
R2676 B.n1117 B.n1116 28.8785
R2677 B.n177 B.n102 28.8785
R2678 B.t3 B.n486 26.3647
R2679 B.n1176 B.t9 26.3647
R2680 B.n1026 B.t4 25.4231
R2681 B.t8 B.n1223 25.4231
R2682 B.t7 B.n470 19.7737
R2683 B.n1192 B.t5 19.7737
R2684 B.n1002 B.t6 18.8321
R2685 B.t1 B.n1207 18.8321
R2686 B B.n1237 18.0485
R2687 B.n893 B.t11 17.8905
R2688 B.t18 B.n1135 17.8905
R2689 B.t11 B.n525 14.1242
R2690 B.n1136 B.t18 14.1242
R2691 B.t6 B.n454 13.1826
R2692 B.n1208 B.t1 13.1826
R2693 B.n978 B.t7 12.241
R2694 B.t5 B.n1191 12.241
R2695 B.n877 B.n539 10.6151
R2696 B.n878 B.n877 10.6151
R2697 B.n879 B.n878 10.6151
R2698 B.n879 B.n531 10.6151
R2699 B.n889 B.n531 10.6151
R2700 B.n890 B.n889 10.6151
R2701 B.n891 B.n890 10.6151
R2702 B.n891 B.n523 10.6151
R2703 B.n901 B.n523 10.6151
R2704 B.n902 B.n901 10.6151
R2705 B.n903 B.n902 10.6151
R2706 B.n903 B.n515 10.6151
R2707 B.n913 B.n515 10.6151
R2708 B.n914 B.n913 10.6151
R2709 B.n915 B.n914 10.6151
R2710 B.n915 B.n507 10.6151
R2711 B.n926 B.n507 10.6151
R2712 B.n927 B.n926 10.6151
R2713 B.n928 B.n927 10.6151
R2714 B.n928 B.n500 10.6151
R2715 B.n938 B.n500 10.6151
R2716 B.n939 B.n938 10.6151
R2717 B.n940 B.n939 10.6151
R2718 B.n940 B.n492 10.6151
R2719 B.n950 B.n492 10.6151
R2720 B.n951 B.n950 10.6151
R2721 B.n952 B.n951 10.6151
R2722 B.n952 B.n484 10.6151
R2723 B.n962 B.n484 10.6151
R2724 B.n963 B.n962 10.6151
R2725 B.n964 B.n963 10.6151
R2726 B.n964 B.n476 10.6151
R2727 B.n974 B.n476 10.6151
R2728 B.n975 B.n974 10.6151
R2729 B.n976 B.n975 10.6151
R2730 B.n976 B.n468 10.6151
R2731 B.n986 B.n468 10.6151
R2732 B.n987 B.n986 10.6151
R2733 B.n988 B.n987 10.6151
R2734 B.n988 B.n460 10.6151
R2735 B.n998 B.n460 10.6151
R2736 B.n999 B.n998 10.6151
R2737 B.n1000 B.n999 10.6151
R2738 B.n1000 B.n452 10.6151
R2739 B.n1010 B.n452 10.6151
R2740 B.n1011 B.n1010 10.6151
R2741 B.n1012 B.n1011 10.6151
R2742 B.n1012 B.n444 10.6151
R2743 B.n1022 B.n444 10.6151
R2744 B.n1023 B.n1022 10.6151
R2745 B.n1024 B.n1023 10.6151
R2746 B.n1024 B.n436 10.6151
R2747 B.n1035 B.n436 10.6151
R2748 B.n1036 B.n1035 10.6151
R2749 B.n1037 B.n1036 10.6151
R2750 B.n1037 B.n0 10.6151
R2751 B.n865 B.n864 10.6151
R2752 B.n864 B.n863 10.6151
R2753 B.n863 B.n862 10.6151
R2754 B.n862 B.n860 10.6151
R2755 B.n860 B.n857 10.6151
R2756 B.n857 B.n856 10.6151
R2757 B.n856 B.n853 10.6151
R2758 B.n853 B.n852 10.6151
R2759 B.n852 B.n849 10.6151
R2760 B.n849 B.n848 10.6151
R2761 B.n848 B.n845 10.6151
R2762 B.n845 B.n844 10.6151
R2763 B.n844 B.n841 10.6151
R2764 B.n841 B.n840 10.6151
R2765 B.n840 B.n837 10.6151
R2766 B.n837 B.n836 10.6151
R2767 B.n836 B.n833 10.6151
R2768 B.n833 B.n832 10.6151
R2769 B.n832 B.n829 10.6151
R2770 B.n829 B.n828 10.6151
R2771 B.n828 B.n825 10.6151
R2772 B.n825 B.n824 10.6151
R2773 B.n824 B.n821 10.6151
R2774 B.n821 B.n820 10.6151
R2775 B.n820 B.n817 10.6151
R2776 B.n817 B.n816 10.6151
R2777 B.n816 B.n813 10.6151
R2778 B.n813 B.n812 10.6151
R2779 B.n812 B.n809 10.6151
R2780 B.n809 B.n808 10.6151
R2781 B.n808 B.n805 10.6151
R2782 B.n805 B.n804 10.6151
R2783 B.n804 B.n801 10.6151
R2784 B.n801 B.n800 10.6151
R2785 B.n800 B.n797 10.6151
R2786 B.n797 B.n796 10.6151
R2787 B.n796 B.n793 10.6151
R2788 B.n793 B.n792 10.6151
R2789 B.n792 B.n789 10.6151
R2790 B.n789 B.n788 10.6151
R2791 B.n788 B.n785 10.6151
R2792 B.n785 B.n784 10.6151
R2793 B.n784 B.n781 10.6151
R2794 B.n781 B.n780 10.6151
R2795 B.n780 B.n777 10.6151
R2796 B.n777 B.n776 10.6151
R2797 B.n776 B.n773 10.6151
R2798 B.n773 B.n772 10.6151
R2799 B.n772 B.n769 10.6151
R2800 B.n769 B.n768 10.6151
R2801 B.n768 B.n765 10.6151
R2802 B.n765 B.n764 10.6151
R2803 B.n764 B.n761 10.6151
R2804 B.n761 B.n760 10.6151
R2805 B.n760 B.n757 10.6151
R2806 B.n757 B.n756 10.6151
R2807 B.n756 B.n753 10.6151
R2808 B.n753 B.n752 10.6151
R2809 B.n752 B.n749 10.6151
R2810 B.n747 B.n744 10.6151
R2811 B.n744 B.n743 10.6151
R2812 B.n743 B.n740 10.6151
R2813 B.n740 B.n739 10.6151
R2814 B.n739 B.n736 10.6151
R2815 B.n736 B.n735 10.6151
R2816 B.n735 B.n732 10.6151
R2817 B.n732 B.n731 10.6151
R2818 B.n728 B.n727 10.6151
R2819 B.n727 B.n724 10.6151
R2820 B.n724 B.n723 10.6151
R2821 B.n723 B.n720 10.6151
R2822 B.n720 B.n719 10.6151
R2823 B.n719 B.n716 10.6151
R2824 B.n716 B.n715 10.6151
R2825 B.n715 B.n712 10.6151
R2826 B.n712 B.n711 10.6151
R2827 B.n711 B.n708 10.6151
R2828 B.n708 B.n707 10.6151
R2829 B.n707 B.n704 10.6151
R2830 B.n704 B.n703 10.6151
R2831 B.n703 B.n700 10.6151
R2832 B.n700 B.n699 10.6151
R2833 B.n699 B.n696 10.6151
R2834 B.n696 B.n695 10.6151
R2835 B.n695 B.n692 10.6151
R2836 B.n692 B.n691 10.6151
R2837 B.n691 B.n688 10.6151
R2838 B.n688 B.n687 10.6151
R2839 B.n687 B.n684 10.6151
R2840 B.n684 B.n683 10.6151
R2841 B.n683 B.n680 10.6151
R2842 B.n680 B.n679 10.6151
R2843 B.n679 B.n676 10.6151
R2844 B.n676 B.n675 10.6151
R2845 B.n675 B.n672 10.6151
R2846 B.n672 B.n671 10.6151
R2847 B.n671 B.n668 10.6151
R2848 B.n668 B.n667 10.6151
R2849 B.n667 B.n664 10.6151
R2850 B.n664 B.n663 10.6151
R2851 B.n663 B.n660 10.6151
R2852 B.n660 B.n659 10.6151
R2853 B.n659 B.n656 10.6151
R2854 B.n656 B.n655 10.6151
R2855 B.n655 B.n652 10.6151
R2856 B.n652 B.n651 10.6151
R2857 B.n651 B.n648 10.6151
R2858 B.n648 B.n647 10.6151
R2859 B.n647 B.n644 10.6151
R2860 B.n644 B.n643 10.6151
R2861 B.n643 B.n640 10.6151
R2862 B.n640 B.n639 10.6151
R2863 B.n639 B.n636 10.6151
R2864 B.n636 B.n635 10.6151
R2865 B.n635 B.n632 10.6151
R2866 B.n632 B.n631 10.6151
R2867 B.n631 B.n628 10.6151
R2868 B.n628 B.n627 10.6151
R2869 B.n627 B.n624 10.6151
R2870 B.n624 B.n623 10.6151
R2871 B.n623 B.n620 10.6151
R2872 B.n620 B.n619 10.6151
R2873 B.n619 B.n616 10.6151
R2874 B.n616 B.n615 10.6151
R2875 B.n615 B.n543 10.6151
R2876 B.n871 B.n543 10.6151
R2877 B.n873 B.n872 10.6151
R2878 B.n873 B.n535 10.6151
R2879 B.n883 B.n535 10.6151
R2880 B.n884 B.n883 10.6151
R2881 B.n885 B.n884 10.6151
R2882 B.n885 B.n527 10.6151
R2883 B.n895 B.n527 10.6151
R2884 B.n896 B.n895 10.6151
R2885 B.n897 B.n896 10.6151
R2886 B.n897 B.n519 10.6151
R2887 B.n907 B.n519 10.6151
R2888 B.n908 B.n907 10.6151
R2889 B.n909 B.n908 10.6151
R2890 B.n909 B.n511 10.6151
R2891 B.n919 B.n511 10.6151
R2892 B.n920 B.n919 10.6151
R2893 B.n921 B.n920 10.6151
R2894 B.n921 B.n504 10.6151
R2895 B.n932 B.n504 10.6151
R2896 B.n933 B.n932 10.6151
R2897 B.n934 B.n933 10.6151
R2898 B.n934 B.n496 10.6151
R2899 B.n944 B.n496 10.6151
R2900 B.n945 B.n944 10.6151
R2901 B.n946 B.n945 10.6151
R2902 B.n946 B.n488 10.6151
R2903 B.n956 B.n488 10.6151
R2904 B.n957 B.n956 10.6151
R2905 B.n958 B.n957 10.6151
R2906 B.n958 B.n480 10.6151
R2907 B.n968 B.n480 10.6151
R2908 B.n969 B.n968 10.6151
R2909 B.n970 B.n969 10.6151
R2910 B.n970 B.n472 10.6151
R2911 B.n980 B.n472 10.6151
R2912 B.n981 B.n980 10.6151
R2913 B.n982 B.n981 10.6151
R2914 B.n982 B.n464 10.6151
R2915 B.n992 B.n464 10.6151
R2916 B.n993 B.n992 10.6151
R2917 B.n994 B.n993 10.6151
R2918 B.n994 B.n456 10.6151
R2919 B.n1004 B.n456 10.6151
R2920 B.n1005 B.n1004 10.6151
R2921 B.n1006 B.n1005 10.6151
R2922 B.n1006 B.n448 10.6151
R2923 B.n1016 B.n448 10.6151
R2924 B.n1017 B.n1016 10.6151
R2925 B.n1018 B.n1017 10.6151
R2926 B.n1018 B.n440 10.6151
R2927 B.n1028 B.n440 10.6151
R2928 B.n1029 B.n1028 10.6151
R2929 B.n1031 B.n1029 10.6151
R2930 B.n1031 B.n1030 10.6151
R2931 B.n1030 B.n432 10.6151
R2932 B.n1042 B.n432 10.6151
R2933 B.n1043 B.n1042 10.6151
R2934 B.n1044 B.n1043 10.6151
R2935 B.n1045 B.n1044 10.6151
R2936 B.n1046 B.n1045 10.6151
R2937 B.n1049 B.n1046 10.6151
R2938 B.n1050 B.n1049 10.6151
R2939 B.n1051 B.n1050 10.6151
R2940 B.n1052 B.n1051 10.6151
R2941 B.n1054 B.n1052 10.6151
R2942 B.n1055 B.n1054 10.6151
R2943 B.n1056 B.n1055 10.6151
R2944 B.n1057 B.n1056 10.6151
R2945 B.n1059 B.n1057 10.6151
R2946 B.n1060 B.n1059 10.6151
R2947 B.n1061 B.n1060 10.6151
R2948 B.n1062 B.n1061 10.6151
R2949 B.n1064 B.n1062 10.6151
R2950 B.n1065 B.n1064 10.6151
R2951 B.n1066 B.n1065 10.6151
R2952 B.n1067 B.n1066 10.6151
R2953 B.n1069 B.n1067 10.6151
R2954 B.n1070 B.n1069 10.6151
R2955 B.n1071 B.n1070 10.6151
R2956 B.n1072 B.n1071 10.6151
R2957 B.n1074 B.n1072 10.6151
R2958 B.n1075 B.n1074 10.6151
R2959 B.n1076 B.n1075 10.6151
R2960 B.n1077 B.n1076 10.6151
R2961 B.n1079 B.n1077 10.6151
R2962 B.n1080 B.n1079 10.6151
R2963 B.n1081 B.n1080 10.6151
R2964 B.n1082 B.n1081 10.6151
R2965 B.n1084 B.n1082 10.6151
R2966 B.n1085 B.n1084 10.6151
R2967 B.n1086 B.n1085 10.6151
R2968 B.n1087 B.n1086 10.6151
R2969 B.n1089 B.n1087 10.6151
R2970 B.n1090 B.n1089 10.6151
R2971 B.n1091 B.n1090 10.6151
R2972 B.n1092 B.n1091 10.6151
R2973 B.n1094 B.n1092 10.6151
R2974 B.n1095 B.n1094 10.6151
R2975 B.n1096 B.n1095 10.6151
R2976 B.n1097 B.n1096 10.6151
R2977 B.n1099 B.n1097 10.6151
R2978 B.n1100 B.n1099 10.6151
R2979 B.n1101 B.n1100 10.6151
R2980 B.n1102 B.n1101 10.6151
R2981 B.n1104 B.n1102 10.6151
R2982 B.n1105 B.n1104 10.6151
R2983 B.n1106 B.n1105 10.6151
R2984 B.n1107 B.n1106 10.6151
R2985 B.n1109 B.n1107 10.6151
R2986 B.n1110 B.n1109 10.6151
R2987 B.n1111 B.n1110 10.6151
R2988 B.n1112 B.n1111 10.6151
R2989 B.n1114 B.n1112 10.6151
R2990 B.n1115 B.n1114 10.6151
R2991 B.n1116 B.n1115 10.6151
R2992 B.n1229 B.n1 10.6151
R2993 B.n1229 B.n1228 10.6151
R2994 B.n1228 B.n1227 10.6151
R2995 B.n1227 B.n10 10.6151
R2996 B.n1221 B.n10 10.6151
R2997 B.n1221 B.n1220 10.6151
R2998 B.n1220 B.n1219 10.6151
R2999 B.n1219 B.n18 10.6151
R3000 B.n1213 B.n18 10.6151
R3001 B.n1213 B.n1212 10.6151
R3002 B.n1212 B.n1211 10.6151
R3003 B.n1211 B.n25 10.6151
R3004 B.n1205 B.n25 10.6151
R3005 B.n1205 B.n1204 10.6151
R3006 B.n1204 B.n1203 10.6151
R3007 B.n1203 B.n32 10.6151
R3008 B.n1197 B.n32 10.6151
R3009 B.n1197 B.n1196 10.6151
R3010 B.n1196 B.n1195 10.6151
R3011 B.n1195 B.n39 10.6151
R3012 B.n1189 B.n39 10.6151
R3013 B.n1189 B.n1188 10.6151
R3014 B.n1188 B.n1187 10.6151
R3015 B.n1187 B.n46 10.6151
R3016 B.n1181 B.n46 10.6151
R3017 B.n1181 B.n1180 10.6151
R3018 B.n1180 B.n1179 10.6151
R3019 B.n1179 B.n53 10.6151
R3020 B.n1173 B.n53 10.6151
R3021 B.n1173 B.n1172 10.6151
R3022 B.n1172 B.n1171 10.6151
R3023 B.n1171 B.n60 10.6151
R3024 B.n1165 B.n60 10.6151
R3025 B.n1165 B.n1164 10.6151
R3026 B.n1164 B.n1163 10.6151
R3027 B.n1163 B.n67 10.6151
R3028 B.n1157 B.n67 10.6151
R3029 B.n1157 B.n1156 10.6151
R3030 B.n1156 B.n1155 10.6151
R3031 B.n1155 B.n73 10.6151
R3032 B.n1149 B.n73 10.6151
R3033 B.n1149 B.n1148 10.6151
R3034 B.n1148 B.n1147 10.6151
R3035 B.n1147 B.n81 10.6151
R3036 B.n1141 B.n81 10.6151
R3037 B.n1141 B.n1140 10.6151
R3038 B.n1140 B.n1139 10.6151
R3039 B.n1139 B.n88 10.6151
R3040 B.n1133 B.n88 10.6151
R3041 B.n1133 B.n1132 10.6151
R3042 B.n1132 B.n1131 10.6151
R3043 B.n1131 B.n95 10.6151
R3044 B.n1125 B.n95 10.6151
R3045 B.n1125 B.n1124 10.6151
R3046 B.n1124 B.n1123 10.6151
R3047 B.n1123 B.n102 10.6151
R3048 B.n178 B.n177 10.6151
R3049 B.n181 B.n178 10.6151
R3050 B.n182 B.n181 10.6151
R3051 B.n185 B.n182 10.6151
R3052 B.n186 B.n185 10.6151
R3053 B.n189 B.n186 10.6151
R3054 B.n190 B.n189 10.6151
R3055 B.n193 B.n190 10.6151
R3056 B.n194 B.n193 10.6151
R3057 B.n197 B.n194 10.6151
R3058 B.n198 B.n197 10.6151
R3059 B.n201 B.n198 10.6151
R3060 B.n202 B.n201 10.6151
R3061 B.n205 B.n202 10.6151
R3062 B.n206 B.n205 10.6151
R3063 B.n209 B.n206 10.6151
R3064 B.n210 B.n209 10.6151
R3065 B.n213 B.n210 10.6151
R3066 B.n214 B.n213 10.6151
R3067 B.n217 B.n214 10.6151
R3068 B.n218 B.n217 10.6151
R3069 B.n221 B.n218 10.6151
R3070 B.n222 B.n221 10.6151
R3071 B.n225 B.n222 10.6151
R3072 B.n226 B.n225 10.6151
R3073 B.n229 B.n226 10.6151
R3074 B.n230 B.n229 10.6151
R3075 B.n233 B.n230 10.6151
R3076 B.n234 B.n233 10.6151
R3077 B.n237 B.n234 10.6151
R3078 B.n238 B.n237 10.6151
R3079 B.n241 B.n238 10.6151
R3080 B.n242 B.n241 10.6151
R3081 B.n245 B.n242 10.6151
R3082 B.n246 B.n245 10.6151
R3083 B.n249 B.n246 10.6151
R3084 B.n250 B.n249 10.6151
R3085 B.n253 B.n250 10.6151
R3086 B.n254 B.n253 10.6151
R3087 B.n257 B.n254 10.6151
R3088 B.n258 B.n257 10.6151
R3089 B.n261 B.n258 10.6151
R3090 B.n262 B.n261 10.6151
R3091 B.n265 B.n262 10.6151
R3092 B.n266 B.n265 10.6151
R3093 B.n269 B.n266 10.6151
R3094 B.n270 B.n269 10.6151
R3095 B.n273 B.n270 10.6151
R3096 B.n274 B.n273 10.6151
R3097 B.n277 B.n274 10.6151
R3098 B.n278 B.n277 10.6151
R3099 B.n281 B.n278 10.6151
R3100 B.n282 B.n281 10.6151
R3101 B.n285 B.n282 10.6151
R3102 B.n286 B.n285 10.6151
R3103 B.n289 B.n286 10.6151
R3104 B.n290 B.n289 10.6151
R3105 B.n293 B.n290 10.6151
R3106 B.n294 B.n293 10.6151
R3107 B.n298 B.n297 10.6151
R3108 B.n301 B.n298 10.6151
R3109 B.n302 B.n301 10.6151
R3110 B.n305 B.n302 10.6151
R3111 B.n306 B.n305 10.6151
R3112 B.n309 B.n306 10.6151
R3113 B.n310 B.n309 10.6151
R3114 B.n313 B.n310 10.6151
R3115 B.n318 B.n315 10.6151
R3116 B.n319 B.n318 10.6151
R3117 B.n322 B.n319 10.6151
R3118 B.n323 B.n322 10.6151
R3119 B.n326 B.n323 10.6151
R3120 B.n327 B.n326 10.6151
R3121 B.n330 B.n327 10.6151
R3122 B.n331 B.n330 10.6151
R3123 B.n334 B.n331 10.6151
R3124 B.n335 B.n334 10.6151
R3125 B.n338 B.n335 10.6151
R3126 B.n339 B.n338 10.6151
R3127 B.n342 B.n339 10.6151
R3128 B.n343 B.n342 10.6151
R3129 B.n346 B.n343 10.6151
R3130 B.n347 B.n346 10.6151
R3131 B.n350 B.n347 10.6151
R3132 B.n351 B.n350 10.6151
R3133 B.n354 B.n351 10.6151
R3134 B.n355 B.n354 10.6151
R3135 B.n358 B.n355 10.6151
R3136 B.n359 B.n358 10.6151
R3137 B.n362 B.n359 10.6151
R3138 B.n363 B.n362 10.6151
R3139 B.n366 B.n363 10.6151
R3140 B.n367 B.n366 10.6151
R3141 B.n370 B.n367 10.6151
R3142 B.n371 B.n370 10.6151
R3143 B.n374 B.n371 10.6151
R3144 B.n375 B.n374 10.6151
R3145 B.n378 B.n375 10.6151
R3146 B.n379 B.n378 10.6151
R3147 B.n382 B.n379 10.6151
R3148 B.n383 B.n382 10.6151
R3149 B.n386 B.n383 10.6151
R3150 B.n387 B.n386 10.6151
R3151 B.n390 B.n387 10.6151
R3152 B.n391 B.n390 10.6151
R3153 B.n394 B.n391 10.6151
R3154 B.n395 B.n394 10.6151
R3155 B.n398 B.n395 10.6151
R3156 B.n399 B.n398 10.6151
R3157 B.n402 B.n399 10.6151
R3158 B.n403 B.n402 10.6151
R3159 B.n406 B.n403 10.6151
R3160 B.n407 B.n406 10.6151
R3161 B.n410 B.n407 10.6151
R3162 B.n411 B.n410 10.6151
R3163 B.n414 B.n411 10.6151
R3164 B.n415 B.n414 10.6151
R3165 B.n418 B.n415 10.6151
R3166 B.n419 B.n418 10.6151
R3167 B.n422 B.n419 10.6151
R3168 B.n423 B.n422 10.6151
R3169 B.n426 B.n423 10.6151
R3170 B.n427 B.n426 10.6151
R3171 B.n430 B.n427 10.6151
R3172 B.n431 B.n430 10.6151
R3173 B.n1117 B.n431 10.6151
R3174 B.n1237 B.n0 8.11757
R3175 B.n1237 B.n1 8.11757
R3176 B.t4 B.n438 6.59156
R3177 B.n1224 B.t8 6.59156
R3178 B.n748 B.n747 6.5566
R3179 B.n731 B.n613 6.5566
R3180 B.n297 B.n175 6.5566
R3181 B.n314 B.n313 6.5566
R3182 B.n954 B.t3 5.64998
R3183 B.t9 B.n1175 5.64998
R3184 B.n749 B.n748 4.05904
R3185 B.n728 B.n613 4.05904
R3186 B.n294 B.n175 4.05904
R3187 B.n315 B.n314 4.05904
R3188 B.n930 B.t0 0.942079
R3189 B.n1159 B.t2 0.942079
R3190 VP.n23 VP.t6 208.897
R3191 VP.n71 VP.t4 177.224
R3192 VP.n53 VP.t1 177.224
R3193 VP.n9 VP.t5 177.224
R3194 VP.n3 VP.t9 177.224
R3195 VP.n89 VP.t8 177.224
R3196 VP.n32 VP.t0 177.224
R3197 VP.n50 VP.t3 177.224
R3198 VP.n16 VP.t7 177.224
R3199 VP.n22 VP.t2 177.224
R3200 VP.n25 VP.n24 161.3
R3201 VP.n26 VP.n21 161.3
R3202 VP.n28 VP.n27 161.3
R3203 VP.n29 VP.n20 161.3
R3204 VP.n31 VP.n30 161.3
R3205 VP.n32 VP.n19 161.3
R3206 VP.n34 VP.n33 161.3
R3207 VP.n35 VP.n18 161.3
R3208 VP.n37 VP.n36 161.3
R3209 VP.n38 VP.n17 161.3
R3210 VP.n40 VP.n39 161.3
R3211 VP.n42 VP.n41 161.3
R3212 VP.n43 VP.n15 161.3
R3213 VP.n45 VP.n44 161.3
R3214 VP.n46 VP.n14 161.3
R3215 VP.n48 VP.n47 161.3
R3216 VP.n49 VP.n13 161.3
R3217 VP.n88 VP.n0 161.3
R3218 VP.n87 VP.n86 161.3
R3219 VP.n85 VP.n1 161.3
R3220 VP.n84 VP.n83 161.3
R3221 VP.n82 VP.n2 161.3
R3222 VP.n81 VP.n80 161.3
R3223 VP.n79 VP.n78 161.3
R3224 VP.n77 VP.n4 161.3
R3225 VP.n76 VP.n75 161.3
R3226 VP.n74 VP.n5 161.3
R3227 VP.n73 VP.n72 161.3
R3228 VP.n71 VP.n6 161.3
R3229 VP.n70 VP.n69 161.3
R3230 VP.n68 VP.n7 161.3
R3231 VP.n67 VP.n66 161.3
R3232 VP.n65 VP.n8 161.3
R3233 VP.n64 VP.n63 161.3
R3234 VP.n62 VP.n61 161.3
R3235 VP.n60 VP.n10 161.3
R3236 VP.n59 VP.n58 161.3
R3237 VP.n57 VP.n11 161.3
R3238 VP.n56 VP.n55 161.3
R3239 VP.n54 VP.n12 161.3
R3240 VP.n53 VP.n52 106.841
R3241 VP.n90 VP.n89 106.841
R3242 VP.n51 VP.n50 106.841
R3243 VP.n23 VP.n22 57.8794
R3244 VP.n52 VP.n51 56.8594
R3245 VP.n59 VP.n11 56.5193
R3246 VP.n83 VP.n1 56.5193
R3247 VP.n44 VP.n14 56.5193
R3248 VP.n66 VP.n7 50.6917
R3249 VP.n76 VP.n5 50.6917
R3250 VP.n37 VP.n18 50.6917
R3251 VP.n27 VP.n20 50.6917
R3252 VP.n66 VP.n65 30.2951
R3253 VP.n77 VP.n76 30.2951
R3254 VP.n38 VP.n37 30.2951
R3255 VP.n27 VP.n26 30.2951
R3256 VP.n55 VP.n54 24.4675
R3257 VP.n55 VP.n11 24.4675
R3258 VP.n60 VP.n59 24.4675
R3259 VP.n61 VP.n60 24.4675
R3260 VP.n65 VP.n64 24.4675
R3261 VP.n70 VP.n7 24.4675
R3262 VP.n71 VP.n70 24.4675
R3263 VP.n72 VP.n71 24.4675
R3264 VP.n72 VP.n5 24.4675
R3265 VP.n78 VP.n77 24.4675
R3266 VP.n82 VP.n81 24.4675
R3267 VP.n83 VP.n82 24.4675
R3268 VP.n87 VP.n1 24.4675
R3269 VP.n88 VP.n87 24.4675
R3270 VP.n48 VP.n14 24.4675
R3271 VP.n49 VP.n48 24.4675
R3272 VP.n39 VP.n38 24.4675
R3273 VP.n43 VP.n42 24.4675
R3274 VP.n44 VP.n43 24.4675
R3275 VP.n31 VP.n20 24.4675
R3276 VP.n32 VP.n31 24.4675
R3277 VP.n33 VP.n32 24.4675
R3278 VP.n33 VP.n18 24.4675
R3279 VP.n26 VP.n25 24.4675
R3280 VP.n64 VP.n9 14.1914
R3281 VP.n78 VP.n3 14.1914
R3282 VP.n39 VP.n16 14.1914
R3283 VP.n25 VP.n22 14.1914
R3284 VP.n61 VP.n9 10.2766
R3285 VP.n81 VP.n3 10.2766
R3286 VP.n42 VP.n16 10.2766
R3287 VP.n24 VP.n23 7.2327
R3288 VP.n54 VP.n53 3.91522
R3289 VP.n89 VP.n88 3.91522
R3290 VP.n50 VP.n49 3.91522
R3291 VP.n51 VP.n13 0.278367
R3292 VP.n52 VP.n12 0.278367
R3293 VP.n90 VP.n0 0.278367
R3294 VP.n24 VP.n21 0.189894
R3295 VP.n28 VP.n21 0.189894
R3296 VP.n29 VP.n28 0.189894
R3297 VP.n30 VP.n29 0.189894
R3298 VP.n30 VP.n19 0.189894
R3299 VP.n34 VP.n19 0.189894
R3300 VP.n35 VP.n34 0.189894
R3301 VP.n36 VP.n35 0.189894
R3302 VP.n36 VP.n17 0.189894
R3303 VP.n40 VP.n17 0.189894
R3304 VP.n41 VP.n40 0.189894
R3305 VP.n41 VP.n15 0.189894
R3306 VP.n45 VP.n15 0.189894
R3307 VP.n46 VP.n45 0.189894
R3308 VP.n47 VP.n46 0.189894
R3309 VP.n47 VP.n13 0.189894
R3310 VP.n56 VP.n12 0.189894
R3311 VP.n57 VP.n56 0.189894
R3312 VP.n58 VP.n57 0.189894
R3313 VP.n58 VP.n10 0.189894
R3314 VP.n62 VP.n10 0.189894
R3315 VP.n63 VP.n62 0.189894
R3316 VP.n63 VP.n8 0.189894
R3317 VP.n67 VP.n8 0.189894
R3318 VP.n68 VP.n67 0.189894
R3319 VP.n69 VP.n68 0.189894
R3320 VP.n69 VP.n6 0.189894
R3321 VP.n73 VP.n6 0.189894
R3322 VP.n74 VP.n73 0.189894
R3323 VP.n75 VP.n74 0.189894
R3324 VP.n75 VP.n4 0.189894
R3325 VP.n79 VP.n4 0.189894
R3326 VP.n80 VP.n79 0.189894
R3327 VP.n80 VP.n2 0.189894
R3328 VP.n84 VP.n2 0.189894
R3329 VP.n85 VP.n84 0.189894
R3330 VP.n86 VP.n85 0.189894
R3331 VP.n86 VP.n0 0.189894
R3332 VP VP.n90 0.153454
R3333 VDD1.n98 VDD1.n97 289.615
R3334 VDD1.n199 VDD1.n198 289.615
R3335 VDD1.n97 VDD1.n96 185
R3336 VDD1.n2 VDD1.n1 185
R3337 VDD1.n91 VDD1.n90 185
R3338 VDD1.n89 VDD1.n88 185
R3339 VDD1.n6 VDD1.n5 185
R3340 VDD1.n83 VDD1.n82 185
R3341 VDD1.n81 VDD1.n80 185
R3342 VDD1.n10 VDD1.n9 185
R3343 VDD1.n75 VDD1.n74 185
R3344 VDD1.n73 VDD1.n72 185
R3345 VDD1.n14 VDD1.n13 185
R3346 VDD1.n67 VDD1.n66 185
R3347 VDD1.n65 VDD1.n64 185
R3348 VDD1.n18 VDD1.n17 185
R3349 VDD1.n59 VDD1.n58 185
R3350 VDD1.n57 VDD1.n56 185
R3351 VDD1.n55 VDD1.n21 185
R3352 VDD1.n25 VDD1.n22 185
R3353 VDD1.n50 VDD1.n49 185
R3354 VDD1.n48 VDD1.n47 185
R3355 VDD1.n27 VDD1.n26 185
R3356 VDD1.n42 VDD1.n41 185
R3357 VDD1.n40 VDD1.n39 185
R3358 VDD1.n31 VDD1.n30 185
R3359 VDD1.n34 VDD1.n33 185
R3360 VDD1.n134 VDD1.n133 185
R3361 VDD1.n131 VDD1.n130 185
R3362 VDD1.n140 VDD1.n139 185
R3363 VDD1.n142 VDD1.n141 185
R3364 VDD1.n127 VDD1.n126 185
R3365 VDD1.n148 VDD1.n147 185
R3366 VDD1.n151 VDD1.n150 185
R3367 VDD1.n149 VDD1.n123 185
R3368 VDD1.n156 VDD1.n122 185
R3369 VDD1.n158 VDD1.n157 185
R3370 VDD1.n160 VDD1.n159 185
R3371 VDD1.n119 VDD1.n118 185
R3372 VDD1.n166 VDD1.n165 185
R3373 VDD1.n168 VDD1.n167 185
R3374 VDD1.n115 VDD1.n114 185
R3375 VDD1.n174 VDD1.n173 185
R3376 VDD1.n176 VDD1.n175 185
R3377 VDD1.n111 VDD1.n110 185
R3378 VDD1.n182 VDD1.n181 185
R3379 VDD1.n184 VDD1.n183 185
R3380 VDD1.n107 VDD1.n106 185
R3381 VDD1.n190 VDD1.n189 185
R3382 VDD1.n192 VDD1.n191 185
R3383 VDD1.n103 VDD1.n102 185
R3384 VDD1.n198 VDD1.n197 185
R3385 VDD1.t3 VDD1.n32 149.524
R3386 VDD1.t8 VDD1.n132 149.524
R3387 VDD1.n97 VDD1.n1 104.615
R3388 VDD1.n90 VDD1.n1 104.615
R3389 VDD1.n90 VDD1.n89 104.615
R3390 VDD1.n89 VDD1.n5 104.615
R3391 VDD1.n82 VDD1.n5 104.615
R3392 VDD1.n82 VDD1.n81 104.615
R3393 VDD1.n81 VDD1.n9 104.615
R3394 VDD1.n74 VDD1.n9 104.615
R3395 VDD1.n74 VDD1.n73 104.615
R3396 VDD1.n73 VDD1.n13 104.615
R3397 VDD1.n66 VDD1.n13 104.615
R3398 VDD1.n66 VDD1.n65 104.615
R3399 VDD1.n65 VDD1.n17 104.615
R3400 VDD1.n58 VDD1.n17 104.615
R3401 VDD1.n58 VDD1.n57 104.615
R3402 VDD1.n57 VDD1.n21 104.615
R3403 VDD1.n25 VDD1.n21 104.615
R3404 VDD1.n49 VDD1.n25 104.615
R3405 VDD1.n49 VDD1.n48 104.615
R3406 VDD1.n48 VDD1.n26 104.615
R3407 VDD1.n41 VDD1.n26 104.615
R3408 VDD1.n41 VDD1.n40 104.615
R3409 VDD1.n40 VDD1.n30 104.615
R3410 VDD1.n33 VDD1.n30 104.615
R3411 VDD1.n133 VDD1.n130 104.615
R3412 VDD1.n140 VDD1.n130 104.615
R3413 VDD1.n141 VDD1.n140 104.615
R3414 VDD1.n141 VDD1.n126 104.615
R3415 VDD1.n148 VDD1.n126 104.615
R3416 VDD1.n150 VDD1.n148 104.615
R3417 VDD1.n150 VDD1.n149 104.615
R3418 VDD1.n149 VDD1.n122 104.615
R3419 VDD1.n158 VDD1.n122 104.615
R3420 VDD1.n159 VDD1.n158 104.615
R3421 VDD1.n159 VDD1.n118 104.615
R3422 VDD1.n166 VDD1.n118 104.615
R3423 VDD1.n167 VDD1.n166 104.615
R3424 VDD1.n167 VDD1.n114 104.615
R3425 VDD1.n174 VDD1.n114 104.615
R3426 VDD1.n175 VDD1.n174 104.615
R3427 VDD1.n175 VDD1.n110 104.615
R3428 VDD1.n182 VDD1.n110 104.615
R3429 VDD1.n183 VDD1.n182 104.615
R3430 VDD1.n183 VDD1.n106 104.615
R3431 VDD1.n190 VDD1.n106 104.615
R3432 VDD1.n191 VDD1.n190 104.615
R3433 VDD1.n191 VDD1.n102 104.615
R3434 VDD1.n198 VDD1.n102 104.615
R3435 VDD1.n203 VDD1.n202 65.928
R3436 VDD1.n100 VDD1.n99 64.1796
R3437 VDD1.n201 VDD1.n200 64.1795
R3438 VDD1.n205 VDD1.n204 64.1785
R3439 VDD1.n100 VDD1.n98 54.1784
R3440 VDD1.n201 VDD1.n199 54.1784
R3441 VDD1.n205 VDD1.n203 52.5203
R3442 VDD1.n33 VDD1.t3 52.3082
R3443 VDD1.n133 VDD1.t8 52.3082
R3444 VDD1.n56 VDD1.n55 13.1884
R3445 VDD1.n157 VDD1.n156 13.1884
R3446 VDD1.n59 VDD1.n20 12.8005
R3447 VDD1.n54 VDD1.n22 12.8005
R3448 VDD1.n155 VDD1.n123 12.8005
R3449 VDD1.n160 VDD1.n121 12.8005
R3450 VDD1.n96 VDD1.n0 12.0247
R3451 VDD1.n60 VDD1.n18 12.0247
R3452 VDD1.n51 VDD1.n50 12.0247
R3453 VDD1.n152 VDD1.n151 12.0247
R3454 VDD1.n161 VDD1.n119 12.0247
R3455 VDD1.n197 VDD1.n101 12.0247
R3456 VDD1.n95 VDD1.n2 11.249
R3457 VDD1.n64 VDD1.n63 11.249
R3458 VDD1.n47 VDD1.n24 11.249
R3459 VDD1.n147 VDD1.n125 11.249
R3460 VDD1.n165 VDD1.n164 11.249
R3461 VDD1.n196 VDD1.n103 11.249
R3462 VDD1.n92 VDD1.n91 10.4732
R3463 VDD1.n67 VDD1.n16 10.4732
R3464 VDD1.n46 VDD1.n27 10.4732
R3465 VDD1.n146 VDD1.n127 10.4732
R3466 VDD1.n168 VDD1.n117 10.4732
R3467 VDD1.n193 VDD1.n192 10.4732
R3468 VDD1.n34 VDD1.n32 10.2747
R3469 VDD1.n134 VDD1.n132 10.2747
R3470 VDD1.n88 VDD1.n4 9.69747
R3471 VDD1.n68 VDD1.n14 9.69747
R3472 VDD1.n43 VDD1.n42 9.69747
R3473 VDD1.n143 VDD1.n142 9.69747
R3474 VDD1.n169 VDD1.n115 9.69747
R3475 VDD1.n189 VDD1.n105 9.69747
R3476 VDD1.n94 VDD1.n0 9.45567
R3477 VDD1.n195 VDD1.n101 9.45567
R3478 VDD1.n36 VDD1.n35 9.3005
R3479 VDD1.n38 VDD1.n37 9.3005
R3480 VDD1.n29 VDD1.n28 9.3005
R3481 VDD1.n44 VDD1.n43 9.3005
R3482 VDD1.n46 VDD1.n45 9.3005
R3483 VDD1.n24 VDD1.n23 9.3005
R3484 VDD1.n52 VDD1.n51 9.3005
R3485 VDD1.n54 VDD1.n53 9.3005
R3486 VDD1.n8 VDD1.n7 9.3005
R3487 VDD1.n85 VDD1.n84 9.3005
R3488 VDD1.n87 VDD1.n86 9.3005
R3489 VDD1.n4 VDD1.n3 9.3005
R3490 VDD1.n93 VDD1.n92 9.3005
R3491 VDD1.n95 VDD1.n94 9.3005
R3492 VDD1.n79 VDD1.n78 9.3005
R3493 VDD1.n77 VDD1.n76 9.3005
R3494 VDD1.n12 VDD1.n11 9.3005
R3495 VDD1.n71 VDD1.n70 9.3005
R3496 VDD1.n69 VDD1.n68 9.3005
R3497 VDD1.n16 VDD1.n15 9.3005
R3498 VDD1.n63 VDD1.n62 9.3005
R3499 VDD1.n61 VDD1.n60 9.3005
R3500 VDD1.n20 VDD1.n19 9.3005
R3501 VDD1.n180 VDD1.n179 9.3005
R3502 VDD1.n109 VDD1.n108 9.3005
R3503 VDD1.n186 VDD1.n185 9.3005
R3504 VDD1.n188 VDD1.n187 9.3005
R3505 VDD1.n105 VDD1.n104 9.3005
R3506 VDD1.n194 VDD1.n193 9.3005
R3507 VDD1.n196 VDD1.n195 9.3005
R3508 VDD1.n113 VDD1.n112 9.3005
R3509 VDD1.n172 VDD1.n171 9.3005
R3510 VDD1.n170 VDD1.n169 9.3005
R3511 VDD1.n117 VDD1.n116 9.3005
R3512 VDD1.n164 VDD1.n163 9.3005
R3513 VDD1.n162 VDD1.n161 9.3005
R3514 VDD1.n121 VDD1.n120 9.3005
R3515 VDD1.n136 VDD1.n135 9.3005
R3516 VDD1.n138 VDD1.n137 9.3005
R3517 VDD1.n129 VDD1.n128 9.3005
R3518 VDD1.n144 VDD1.n143 9.3005
R3519 VDD1.n146 VDD1.n145 9.3005
R3520 VDD1.n125 VDD1.n124 9.3005
R3521 VDD1.n153 VDD1.n152 9.3005
R3522 VDD1.n155 VDD1.n154 9.3005
R3523 VDD1.n178 VDD1.n177 9.3005
R3524 VDD1.n87 VDD1.n6 8.92171
R3525 VDD1.n72 VDD1.n71 8.92171
R3526 VDD1.n39 VDD1.n29 8.92171
R3527 VDD1.n139 VDD1.n129 8.92171
R3528 VDD1.n173 VDD1.n172 8.92171
R3529 VDD1.n188 VDD1.n107 8.92171
R3530 VDD1.n84 VDD1.n83 8.14595
R3531 VDD1.n75 VDD1.n12 8.14595
R3532 VDD1.n38 VDD1.n31 8.14595
R3533 VDD1.n138 VDD1.n131 8.14595
R3534 VDD1.n176 VDD1.n113 8.14595
R3535 VDD1.n185 VDD1.n184 8.14595
R3536 VDD1.n80 VDD1.n8 7.3702
R3537 VDD1.n76 VDD1.n10 7.3702
R3538 VDD1.n35 VDD1.n34 7.3702
R3539 VDD1.n135 VDD1.n134 7.3702
R3540 VDD1.n177 VDD1.n111 7.3702
R3541 VDD1.n181 VDD1.n109 7.3702
R3542 VDD1.n80 VDD1.n79 6.59444
R3543 VDD1.n79 VDD1.n10 6.59444
R3544 VDD1.n180 VDD1.n111 6.59444
R3545 VDD1.n181 VDD1.n180 6.59444
R3546 VDD1.n83 VDD1.n8 5.81868
R3547 VDD1.n76 VDD1.n75 5.81868
R3548 VDD1.n35 VDD1.n31 5.81868
R3549 VDD1.n135 VDD1.n131 5.81868
R3550 VDD1.n177 VDD1.n176 5.81868
R3551 VDD1.n184 VDD1.n109 5.81868
R3552 VDD1.n84 VDD1.n6 5.04292
R3553 VDD1.n72 VDD1.n12 5.04292
R3554 VDD1.n39 VDD1.n38 5.04292
R3555 VDD1.n139 VDD1.n138 5.04292
R3556 VDD1.n173 VDD1.n113 5.04292
R3557 VDD1.n185 VDD1.n107 5.04292
R3558 VDD1.n88 VDD1.n87 4.26717
R3559 VDD1.n71 VDD1.n14 4.26717
R3560 VDD1.n42 VDD1.n29 4.26717
R3561 VDD1.n142 VDD1.n129 4.26717
R3562 VDD1.n172 VDD1.n115 4.26717
R3563 VDD1.n189 VDD1.n188 4.26717
R3564 VDD1.n91 VDD1.n4 3.49141
R3565 VDD1.n68 VDD1.n67 3.49141
R3566 VDD1.n43 VDD1.n27 3.49141
R3567 VDD1.n143 VDD1.n127 3.49141
R3568 VDD1.n169 VDD1.n168 3.49141
R3569 VDD1.n192 VDD1.n105 3.49141
R3570 VDD1.n36 VDD1.n32 2.84303
R3571 VDD1.n136 VDD1.n132 2.84303
R3572 VDD1.n92 VDD1.n2 2.71565
R3573 VDD1.n64 VDD1.n16 2.71565
R3574 VDD1.n47 VDD1.n46 2.71565
R3575 VDD1.n147 VDD1.n146 2.71565
R3576 VDD1.n165 VDD1.n117 2.71565
R3577 VDD1.n193 VDD1.n103 2.71565
R3578 VDD1.n96 VDD1.n95 1.93989
R3579 VDD1.n63 VDD1.n18 1.93989
R3580 VDD1.n50 VDD1.n24 1.93989
R3581 VDD1.n151 VDD1.n125 1.93989
R3582 VDD1.n164 VDD1.n119 1.93989
R3583 VDD1.n197 VDD1.n196 1.93989
R3584 VDD1 VDD1.n205 1.74619
R3585 VDD1.n98 VDD1.n0 1.16414
R3586 VDD1.n60 VDD1.n59 1.16414
R3587 VDD1.n51 VDD1.n22 1.16414
R3588 VDD1.n152 VDD1.n123 1.16414
R3589 VDD1.n161 VDD1.n160 1.16414
R3590 VDD1.n199 VDD1.n101 1.16414
R3591 VDD1.n204 VDD1.t2 1.09503
R3592 VDD1.n204 VDD1.t6 1.09503
R3593 VDD1.n99 VDD1.t7 1.09503
R3594 VDD1.n99 VDD1.t9 1.09503
R3595 VDD1.n202 VDD1.t0 1.09503
R3596 VDD1.n202 VDD1.t1 1.09503
R3597 VDD1.n200 VDD1.t4 1.09503
R3598 VDD1.n200 VDD1.t5 1.09503
R3599 VDD1 VDD1.n100 0.659983
R3600 VDD1.n203 VDD1.n201 0.546447
R3601 VDD1.n56 VDD1.n20 0.388379
R3602 VDD1.n55 VDD1.n54 0.388379
R3603 VDD1.n156 VDD1.n155 0.388379
R3604 VDD1.n157 VDD1.n121 0.388379
R3605 VDD1.n94 VDD1.n93 0.155672
R3606 VDD1.n93 VDD1.n3 0.155672
R3607 VDD1.n86 VDD1.n3 0.155672
R3608 VDD1.n86 VDD1.n85 0.155672
R3609 VDD1.n85 VDD1.n7 0.155672
R3610 VDD1.n78 VDD1.n7 0.155672
R3611 VDD1.n78 VDD1.n77 0.155672
R3612 VDD1.n77 VDD1.n11 0.155672
R3613 VDD1.n70 VDD1.n11 0.155672
R3614 VDD1.n70 VDD1.n69 0.155672
R3615 VDD1.n69 VDD1.n15 0.155672
R3616 VDD1.n62 VDD1.n15 0.155672
R3617 VDD1.n62 VDD1.n61 0.155672
R3618 VDD1.n61 VDD1.n19 0.155672
R3619 VDD1.n53 VDD1.n19 0.155672
R3620 VDD1.n53 VDD1.n52 0.155672
R3621 VDD1.n52 VDD1.n23 0.155672
R3622 VDD1.n45 VDD1.n23 0.155672
R3623 VDD1.n45 VDD1.n44 0.155672
R3624 VDD1.n44 VDD1.n28 0.155672
R3625 VDD1.n37 VDD1.n28 0.155672
R3626 VDD1.n37 VDD1.n36 0.155672
R3627 VDD1.n137 VDD1.n136 0.155672
R3628 VDD1.n137 VDD1.n128 0.155672
R3629 VDD1.n144 VDD1.n128 0.155672
R3630 VDD1.n145 VDD1.n144 0.155672
R3631 VDD1.n145 VDD1.n124 0.155672
R3632 VDD1.n153 VDD1.n124 0.155672
R3633 VDD1.n154 VDD1.n153 0.155672
R3634 VDD1.n154 VDD1.n120 0.155672
R3635 VDD1.n162 VDD1.n120 0.155672
R3636 VDD1.n163 VDD1.n162 0.155672
R3637 VDD1.n163 VDD1.n116 0.155672
R3638 VDD1.n170 VDD1.n116 0.155672
R3639 VDD1.n171 VDD1.n170 0.155672
R3640 VDD1.n171 VDD1.n112 0.155672
R3641 VDD1.n178 VDD1.n112 0.155672
R3642 VDD1.n179 VDD1.n178 0.155672
R3643 VDD1.n179 VDD1.n108 0.155672
R3644 VDD1.n186 VDD1.n108 0.155672
R3645 VDD1.n187 VDD1.n186 0.155672
R3646 VDD1.n187 VDD1.n104 0.155672
R3647 VDD1.n194 VDD1.n104 0.155672
R3648 VDD1.n195 VDD1.n194 0.155672
C0 VDD2 VP 0.566272f
C1 VTAIL VDD2 13.3084f
C2 VDD2 VN 15.640201f
C3 VDD1 VDD2 2.08434f
C4 VTAIL VP 15.968401f
C5 VP VN 9.32495f
C6 VDD1 VP 16.0484f
C7 VTAIL VN 15.954f
C8 VTAIL VDD1 13.26f
C9 VDD1 VN 0.153082f
C10 VDD2 B 8.114809f
C11 VDD1 B 8.098035f
C12 VTAIL B 10.515832f
C13 VN B 18.002869f
C14 VP B 16.41328f
C15 VDD1.n0 B 0.013337f
C16 VDD1.n1 B 0.030033f
C17 VDD1.n2 B 0.013454f
C18 VDD1.n3 B 0.023646f
C19 VDD1.n4 B 0.012706f
C20 VDD1.n5 B 0.030033f
C21 VDD1.n6 B 0.013454f
C22 VDD1.n7 B 0.023646f
C23 VDD1.n8 B 0.012706f
C24 VDD1.n9 B 0.030033f
C25 VDD1.n10 B 0.013454f
C26 VDD1.n11 B 0.023646f
C27 VDD1.n12 B 0.012706f
C28 VDD1.n13 B 0.030033f
C29 VDD1.n14 B 0.013454f
C30 VDD1.n15 B 0.023646f
C31 VDD1.n16 B 0.012706f
C32 VDD1.n17 B 0.030033f
C33 VDD1.n18 B 0.013454f
C34 VDD1.n19 B 0.023646f
C35 VDD1.n20 B 0.012706f
C36 VDD1.n21 B 0.030033f
C37 VDD1.n22 B 0.013454f
C38 VDD1.n23 B 0.023646f
C39 VDD1.n24 B 0.012706f
C40 VDD1.n25 B 0.030033f
C41 VDD1.n26 B 0.030033f
C42 VDD1.n27 B 0.013454f
C43 VDD1.n28 B 0.023646f
C44 VDD1.n29 B 0.012706f
C45 VDD1.n30 B 0.030033f
C46 VDD1.n31 B 0.013454f
C47 VDD1.n32 B 0.225769f
C48 VDD1.t3 B 0.051499f
C49 VDD1.n33 B 0.022525f
C50 VDD1.n34 B 0.021231f
C51 VDD1.n35 B 0.012706f
C52 VDD1.n36 B 1.8334f
C53 VDD1.n37 B 0.023646f
C54 VDD1.n38 B 0.012706f
C55 VDD1.n39 B 0.013454f
C56 VDD1.n40 B 0.030033f
C57 VDD1.n41 B 0.030033f
C58 VDD1.n42 B 0.013454f
C59 VDD1.n43 B 0.012706f
C60 VDD1.n44 B 0.023646f
C61 VDD1.n45 B 0.023646f
C62 VDD1.n46 B 0.012706f
C63 VDD1.n47 B 0.013454f
C64 VDD1.n48 B 0.030033f
C65 VDD1.n49 B 0.030033f
C66 VDD1.n50 B 0.013454f
C67 VDD1.n51 B 0.012706f
C68 VDD1.n52 B 0.023646f
C69 VDD1.n53 B 0.023646f
C70 VDD1.n54 B 0.012706f
C71 VDD1.n55 B 0.01308f
C72 VDD1.n56 B 0.01308f
C73 VDD1.n57 B 0.030033f
C74 VDD1.n58 B 0.030033f
C75 VDD1.n59 B 0.013454f
C76 VDD1.n60 B 0.012706f
C77 VDD1.n61 B 0.023646f
C78 VDD1.n62 B 0.023646f
C79 VDD1.n63 B 0.012706f
C80 VDD1.n64 B 0.013454f
C81 VDD1.n65 B 0.030033f
C82 VDD1.n66 B 0.030033f
C83 VDD1.n67 B 0.013454f
C84 VDD1.n68 B 0.012706f
C85 VDD1.n69 B 0.023646f
C86 VDD1.n70 B 0.023646f
C87 VDD1.n71 B 0.012706f
C88 VDD1.n72 B 0.013454f
C89 VDD1.n73 B 0.030033f
C90 VDD1.n74 B 0.030033f
C91 VDD1.n75 B 0.013454f
C92 VDD1.n76 B 0.012706f
C93 VDD1.n77 B 0.023646f
C94 VDD1.n78 B 0.023646f
C95 VDD1.n79 B 0.012706f
C96 VDD1.n80 B 0.013454f
C97 VDD1.n81 B 0.030033f
C98 VDD1.n82 B 0.030033f
C99 VDD1.n83 B 0.013454f
C100 VDD1.n84 B 0.012706f
C101 VDD1.n85 B 0.023646f
C102 VDD1.n86 B 0.023646f
C103 VDD1.n87 B 0.012706f
C104 VDD1.n88 B 0.013454f
C105 VDD1.n89 B 0.030033f
C106 VDD1.n90 B 0.030033f
C107 VDD1.n91 B 0.013454f
C108 VDD1.n92 B 0.012706f
C109 VDD1.n93 B 0.023646f
C110 VDD1.n94 B 0.06144f
C111 VDD1.n95 B 0.012706f
C112 VDD1.n96 B 0.013454f
C113 VDD1.n97 B 0.060784f
C114 VDD1.n98 B 0.078204f
C115 VDD1.t7 B 0.338023f
C116 VDD1.t9 B 0.338023f
C117 VDD1.n99 B 3.08961f
C118 VDD1.n100 B 0.641678f
C119 VDD1.n101 B 0.013337f
C120 VDD1.n102 B 0.030033f
C121 VDD1.n103 B 0.013454f
C122 VDD1.n104 B 0.023646f
C123 VDD1.n105 B 0.012706f
C124 VDD1.n106 B 0.030033f
C125 VDD1.n107 B 0.013454f
C126 VDD1.n108 B 0.023646f
C127 VDD1.n109 B 0.012706f
C128 VDD1.n110 B 0.030033f
C129 VDD1.n111 B 0.013454f
C130 VDD1.n112 B 0.023646f
C131 VDD1.n113 B 0.012706f
C132 VDD1.n114 B 0.030033f
C133 VDD1.n115 B 0.013454f
C134 VDD1.n116 B 0.023646f
C135 VDD1.n117 B 0.012706f
C136 VDD1.n118 B 0.030033f
C137 VDD1.n119 B 0.013454f
C138 VDD1.n120 B 0.023646f
C139 VDD1.n121 B 0.012706f
C140 VDD1.n122 B 0.030033f
C141 VDD1.n123 B 0.013454f
C142 VDD1.n124 B 0.023646f
C143 VDD1.n125 B 0.012706f
C144 VDD1.n126 B 0.030033f
C145 VDD1.n127 B 0.013454f
C146 VDD1.n128 B 0.023646f
C147 VDD1.n129 B 0.012706f
C148 VDD1.n130 B 0.030033f
C149 VDD1.n131 B 0.013454f
C150 VDD1.n132 B 0.225769f
C151 VDD1.t8 B 0.051499f
C152 VDD1.n133 B 0.022525f
C153 VDD1.n134 B 0.021231f
C154 VDD1.n135 B 0.012706f
C155 VDD1.n136 B 1.8334f
C156 VDD1.n137 B 0.023646f
C157 VDD1.n138 B 0.012706f
C158 VDD1.n139 B 0.013454f
C159 VDD1.n140 B 0.030033f
C160 VDD1.n141 B 0.030033f
C161 VDD1.n142 B 0.013454f
C162 VDD1.n143 B 0.012706f
C163 VDD1.n144 B 0.023646f
C164 VDD1.n145 B 0.023646f
C165 VDD1.n146 B 0.012706f
C166 VDD1.n147 B 0.013454f
C167 VDD1.n148 B 0.030033f
C168 VDD1.n149 B 0.030033f
C169 VDD1.n150 B 0.030033f
C170 VDD1.n151 B 0.013454f
C171 VDD1.n152 B 0.012706f
C172 VDD1.n153 B 0.023646f
C173 VDD1.n154 B 0.023646f
C174 VDD1.n155 B 0.012706f
C175 VDD1.n156 B 0.01308f
C176 VDD1.n157 B 0.01308f
C177 VDD1.n158 B 0.030033f
C178 VDD1.n159 B 0.030033f
C179 VDD1.n160 B 0.013454f
C180 VDD1.n161 B 0.012706f
C181 VDD1.n162 B 0.023646f
C182 VDD1.n163 B 0.023646f
C183 VDD1.n164 B 0.012706f
C184 VDD1.n165 B 0.013454f
C185 VDD1.n166 B 0.030033f
C186 VDD1.n167 B 0.030033f
C187 VDD1.n168 B 0.013454f
C188 VDD1.n169 B 0.012706f
C189 VDD1.n170 B 0.023646f
C190 VDD1.n171 B 0.023646f
C191 VDD1.n172 B 0.012706f
C192 VDD1.n173 B 0.013454f
C193 VDD1.n174 B 0.030033f
C194 VDD1.n175 B 0.030033f
C195 VDD1.n176 B 0.013454f
C196 VDD1.n177 B 0.012706f
C197 VDD1.n178 B 0.023646f
C198 VDD1.n179 B 0.023646f
C199 VDD1.n180 B 0.012706f
C200 VDD1.n181 B 0.013454f
C201 VDD1.n182 B 0.030033f
C202 VDD1.n183 B 0.030033f
C203 VDD1.n184 B 0.013454f
C204 VDD1.n185 B 0.012706f
C205 VDD1.n186 B 0.023646f
C206 VDD1.n187 B 0.023646f
C207 VDD1.n188 B 0.012706f
C208 VDD1.n189 B 0.013454f
C209 VDD1.n190 B 0.030033f
C210 VDD1.n191 B 0.030033f
C211 VDD1.n192 B 0.013454f
C212 VDD1.n193 B 0.012706f
C213 VDD1.n194 B 0.023646f
C214 VDD1.n195 B 0.06144f
C215 VDD1.n196 B 0.012706f
C216 VDD1.n197 B 0.013454f
C217 VDD1.n198 B 0.060784f
C218 VDD1.n199 B 0.078204f
C219 VDD1.t4 B 0.338023f
C220 VDD1.t5 B 0.338023f
C221 VDD1.n200 B 3.08961f
C222 VDD1.n201 B 0.634037f
C223 VDD1.t0 B 0.338023f
C224 VDD1.t1 B 0.338023f
C225 VDD1.n202 B 3.10322f
C226 VDD1.n203 B 3.15021f
C227 VDD1.t2 B 0.338023f
C228 VDD1.t6 B 0.338023f
C229 VDD1.n204 B 3.08961f
C230 VDD1.n205 B 3.37481f
C231 VP.n0 B 0.028386f
C232 VP.t8 B 2.63568f
C233 VP.n1 B 0.035333f
C234 VP.n2 B 0.021531f
C235 VP.t9 B 2.63568f
C236 VP.n3 B 0.914865f
C237 VP.n4 B 0.021531f
C238 VP.n5 B 0.039308f
C239 VP.n6 B 0.021531f
C240 VP.t4 B 2.63568f
C241 VP.n7 B 0.039308f
C242 VP.n8 B 0.021531f
C243 VP.t5 B 2.63568f
C244 VP.n9 B 0.914865f
C245 VP.n10 B 0.021531f
C246 VP.n11 B 0.035333f
C247 VP.n12 B 0.028386f
C248 VP.t1 B 2.63568f
C249 VP.n13 B 0.028386f
C250 VP.t3 B 2.63568f
C251 VP.n14 B 0.035333f
C252 VP.n15 B 0.021531f
C253 VP.t7 B 2.63568f
C254 VP.n16 B 0.914865f
C255 VP.n17 B 0.021531f
C256 VP.n18 B 0.039308f
C257 VP.n19 B 0.021531f
C258 VP.t0 B 2.63568f
C259 VP.n20 B 0.039308f
C260 VP.n21 B 0.021531f
C261 VP.t2 B 2.63568f
C262 VP.n22 B 0.976507f
C263 VP.t6 B 2.79355f
C264 VP.n23 B 0.963382f
C265 VP.n24 B 0.204421f
C266 VP.n25 B 0.031807f
C267 VP.n26 B 0.043024f
C268 VP.n27 B 0.020662f
C269 VP.n28 B 0.021531f
C270 VP.n29 B 0.021531f
C271 VP.n30 B 0.021531f
C272 VP.n31 B 0.040128f
C273 VP.n32 B 0.935181f
C274 VP.n33 B 0.040128f
C275 VP.n34 B 0.021531f
C276 VP.n35 B 0.021531f
C277 VP.n36 B 0.021531f
C278 VP.n37 B 0.020662f
C279 VP.n38 B 0.043024f
C280 VP.n39 B 0.031807f
C281 VP.n40 B 0.021531f
C282 VP.n41 B 0.021531f
C283 VP.n42 B 0.028637f
C284 VP.n43 B 0.040128f
C285 VP.n44 B 0.027533f
C286 VP.n45 B 0.021531f
C287 VP.n46 B 0.021531f
C288 VP.n47 B 0.021531f
C289 VP.n48 B 0.040128f
C290 VP.n49 B 0.023486f
C291 VP.n50 B 0.976187f
C292 VP.n51 B 1.43993f
C293 VP.n52 B 1.45354f
C294 VP.n53 B 0.976187f
C295 VP.n54 B 0.023486f
C296 VP.n55 B 0.040128f
C297 VP.n56 B 0.021531f
C298 VP.n57 B 0.021531f
C299 VP.n58 B 0.021531f
C300 VP.n59 B 0.027533f
C301 VP.n60 B 0.040128f
C302 VP.n61 B 0.028637f
C303 VP.n62 B 0.021531f
C304 VP.n63 B 0.021531f
C305 VP.n64 B 0.031807f
C306 VP.n65 B 0.043024f
C307 VP.n66 B 0.020662f
C308 VP.n67 B 0.021531f
C309 VP.n68 B 0.021531f
C310 VP.n69 B 0.021531f
C311 VP.n70 B 0.040128f
C312 VP.n71 B 0.935181f
C313 VP.n72 B 0.040128f
C314 VP.n73 B 0.021531f
C315 VP.n74 B 0.021531f
C316 VP.n75 B 0.021531f
C317 VP.n76 B 0.020662f
C318 VP.n77 B 0.043024f
C319 VP.n78 B 0.031807f
C320 VP.n79 B 0.021531f
C321 VP.n80 B 0.021531f
C322 VP.n81 B 0.028637f
C323 VP.n82 B 0.040128f
C324 VP.n83 B 0.027533f
C325 VP.n84 B 0.021531f
C326 VP.n85 B 0.021531f
C327 VP.n86 B 0.021531f
C328 VP.n87 B 0.040128f
C329 VP.n88 B 0.023486f
C330 VP.n89 B 0.976187f
C331 VP.n90 B 0.036836f
C332 VTAIL.t13 B 0.337981f
C333 VTAIL.t7 B 0.337981f
C334 VTAIL.n0 B 3.02519f
C335 VTAIL.n1 B 0.488044f
C336 VTAIL.n2 B 0.013335f
C337 VTAIL.n3 B 0.030029f
C338 VTAIL.n4 B 0.013452f
C339 VTAIL.n5 B 0.023643f
C340 VTAIL.n6 B 0.012705f
C341 VTAIL.n7 B 0.030029f
C342 VTAIL.n8 B 0.013452f
C343 VTAIL.n9 B 0.023643f
C344 VTAIL.n10 B 0.012705f
C345 VTAIL.n11 B 0.030029f
C346 VTAIL.n12 B 0.013452f
C347 VTAIL.n13 B 0.023643f
C348 VTAIL.n14 B 0.012705f
C349 VTAIL.n15 B 0.030029f
C350 VTAIL.n16 B 0.013452f
C351 VTAIL.n17 B 0.023643f
C352 VTAIL.n18 B 0.012705f
C353 VTAIL.n19 B 0.030029f
C354 VTAIL.n20 B 0.013452f
C355 VTAIL.n21 B 0.023643f
C356 VTAIL.n22 B 0.012705f
C357 VTAIL.n23 B 0.030029f
C358 VTAIL.n24 B 0.013452f
C359 VTAIL.n25 B 0.023643f
C360 VTAIL.n26 B 0.012705f
C361 VTAIL.n27 B 0.030029f
C362 VTAIL.n28 B 0.013452f
C363 VTAIL.n29 B 0.023643f
C364 VTAIL.n30 B 0.012705f
C365 VTAIL.n31 B 0.030029f
C366 VTAIL.n32 B 0.013452f
C367 VTAIL.n33 B 0.225741f
C368 VTAIL.t4 B 0.051493f
C369 VTAIL.n34 B 0.022522f
C370 VTAIL.n35 B 0.021228f
C371 VTAIL.n36 B 0.012705f
C372 VTAIL.n37 B 1.83317f
C373 VTAIL.n38 B 0.023643f
C374 VTAIL.n39 B 0.012705f
C375 VTAIL.n40 B 0.013452f
C376 VTAIL.n41 B 0.030029f
C377 VTAIL.n42 B 0.030029f
C378 VTAIL.n43 B 0.013452f
C379 VTAIL.n44 B 0.012705f
C380 VTAIL.n45 B 0.023643f
C381 VTAIL.n46 B 0.023643f
C382 VTAIL.n47 B 0.012705f
C383 VTAIL.n48 B 0.013452f
C384 VTAIL.n49 B 0.030029f
C385 VTAIL.n50 B 0.030029f
C386 VTAIL.n51 B 0.030029f
C387 VTAIL.n52 B 0.013452f
C388 VTAIL.n53 B 0.012705f
C389 VTAIL.n54 B 0.023643f
C390 VTAIL.n55 B 0.023643f
C391 VTAIL.n56 B 0.012705f
C392 VTAIL.n57 B 0.013078f
C393 VTAIL.n58 B 0.013078f
C394 VTAIL.n59 B 0.030029f
C395 VTAIL.n60 B 0.030029f
C396 VTAIL.n61 B 0.013452f
C397 VTAIL.n62 B 0.012705f
C398 VTAIL.n63 B 0.023643f
C399 VTAIL.n64 B 0.023643f
C400 VTAIL.n65 B 0.012705f
C401 VTAIL.n66 B 0.013452f
C402 VTAIL.n67 B 0.030029f
C403 VTAIL.n68 B 0.030029f
C404 VTAIL.n69 B 0.013452f
C405 VTAIL.n70 B 0.012705f
C406 VTAIL.n71 B 0.023643f
C407 VTAIL.n72 B 0.023643f
C408 VTAIL.n73 B 0.012705f
C409 VTAIL.n74 B 0.013452f
C410 VTAIL.n75 B 0.030029f
C411 VTAIL.n76 B 0.030029f
C412 VTAIL.n77 B 0.013452f
C413 VTAIL.n78 B 0.012705f
C414 VTAIL.n79 B 0.023643f
C415 VTAIL.n80 B 0.023643f
C416 VTAIL.n81 B 0.012705f
C417 VTAIL.n82 B 0.013452f
C418 VTAIL.n83 B 0.030029f
C419 VTAIL.n84 B 0.030029f
C420 VTAIL.n85 B 0.013452f
C421 VTAIL.n86 B 0.012705f
C422 VTAIL.n87 B 0.023643f
C423 VTAIL.n88 B 0.023643f
C424 VTAIL.n89 B 0.012705f
C425 VTAIL.n90 B 0.013452f
C426 VTAIL.n91 B 0.030029f
C427 VTAIL.n92 B 0.030029f
C428 VTAIL.n93 B 0.013452f
C429 VTAIL.n94 B 0.012705f
C430 VTAIL.n95 B 0.023643f
C431 VTAIL.n96 B 0.061432f
C432 VTAIL.n97 B 0.012705f
C433 VTAIL.n98 B 0.013452f
C434 VTAIL.n99 B 0.060777f
C435 VTAIL.n100 B 0.051626f
C436 VTAIL.n101 B 0.333574f
C437 VTAIL.t17 B 0.337981f
C438 VTAIL.t6 B 0.337981f
C439 VTAIL.n102 B 3.02519f
C440 VTAIL.n103 B 0.585242f
C441 VTAIL.t0 B 0.337981f
C442 VTAIL.t3 B 0.337981f
C443 VTAIL.n104 B 3.02519f
C444 VTAIL.n105 B 2.27769f
C445 VTAIL.t11 B 0.337981f
C446 VTAIL.t15 B 0.337981f
C447 VTAIL.n106 B 3.0252f
C448 VTAIL.n107 B 2.27768f
C449 VTAIL.t12 B 0.337981f
C450 VTAIL.t10 B 0.337981f
C451 VTAIL.n108 B 3.0252f
C452 VTAIL.n109 B 0.585236f
C453 VTAIL.n110 B 0.013335f
C454 VTAIL.n111 B 0.030029f
C455 VTAIL.n112 B 0.013452f
C456 VTAIL.n113 B 0.023643f
C457 VTAIL.n114 B 0.012705f
C458 VTAIL.n115 B 0.030029f
C459 VTAIL.n116 B 0.013452f
C460 VTAIL.n117 B 0.023643f
C461 VTAIL.n118 B 0.012705f
C462 VTAIL.n119 B 0.030029f
C463 VTAIL.n120 B 0.013452f
C464 VTAIL.n121 B 0.023643f
C465 VTAIL.n122 B 0.012705f
C466 VTAIL.n123 B 0.030029f
C467 VTAIL.n124 B 0.013452f
C468 VTAIL.n125 B 0.023643f
C469 VTAIL.n126 B 0.012705f
C470 VTAIL.n127 B 0.030029f
C471 VTAIL.n128 B 0.013452f
C472 VTAIL.n129 B 0.023643f
C473 VTAIL.n130 B 0.012705f
C474 VTAIL.n131 B 0.030029f
C475 VTAIL.n132 B 0.013452f
C476 VTAIL.n133 B 0.023643f
C477 VTAIL.n134 B 0.012705f
C478 VTAIL.n135 B 0.030029f
C479 VTAIL.n136 B 0.030029f
C480 VTAIL.n137 B 0.013452f
C481 VTAIL.n138 B 0.023643f
C482 VTAIL.n139 B 0.012705f
C483 VTAIL.n140 B 0.030029f
C484 VTAIL.n141 B 0.013452f
C485 VTAIL.n142 B 0.225741f
C486 VTAIL.t9 B 0.051493f
C487 VTAIL.n143 B 0.022522f
C488 VTAIL.n144 B 0.021228f
C489 VTAIL.n145 B 0.012705f
C490 VTAIL.n146 B 1.83317f
C491 VTAIL.n147 B 0.023643f
C492 VTAIL.n148 B 0.012705f
C493 VTAIL.n149 B 0.013452f
C494 VTAIL.n150 B 0.030029f
C495 VTAIL.n151 B 0.030029f
C496 VTAIL.n152 B 0.013452f
C497 VTAIL.n153 B 0.012705f
C498 VTAIL.n154 B 0.023643f
C499 VTAIL.n155 B 0.023643f
C500 VTAIL.n156 B 0.012705f
C501 VTAIL.n157 B 0.013452f
C502 VTAIL.n158 B 0.030029f
C503 VTAIL.n159 B 0.030029f
C504 VTAIL.n160 B 0.013452f
C505 VTAIL.n161 B 0.012705f
C506 VTAIL.n162 B 0.023643f
C507 VTAIL.n163 B 0.023643f
C508 VTAIL.n164 B 0.012705f
C509 VTAIL.n165 B 0.013078f
C510 VTAIL.n166 B 0.013078f
C511 VTAIL.n167 B 0.030029f
C512 VTAIL.n168 B 0.030029f
C513 VTAIL.n169 B 0.013452f
C514 VTAIL.n170 B 0.012705f
C515 VTAIL.n171 B 0.023643f
C516 VTAIL.n172 B 0.023643f
C517 VTAIL.n173 B 0.012705f
C518 VTAIL.n174 B 0.013452f
C519 VTAIL.n175 B 0.030029f
C520 VTAIL.n176 B 0.030029f
C521 VTAIL.n177 B 0.013452f
C522 VTAIL.n178 B 0.012705f
C523 VTAIL.n179 B 0.023643f
C524 VTAIL.n180 B 0.023643f
C525 VTAIL.n181 B 0.012705f
C526 VTAIL.n182 B 0.013452f
C527 VTAIL.n183 B 0.030029f
C528 VTAIL.n184 B 0.030029f
C529 VTAIL.n185 B 0.013452f
C530 VTAIL.n186 B 0.012705f
C531 VTAIL.n187 B 0.023643f
C532 VTAIL.n188 B 0.023643f
C533 VTAIL.n189 B 0.012705f
C534 VTAIL.n190 B 0.013452f
C535 VTAIL.n191 B 0.030029f
C536 VTAIL.n192 B 0.030029f
C537 VTAIL.n193 B 0.013452f
C538 VTAIL.n194 B 0.012705f
C539 VTAIL.n195 B 0.023643f
C540 VTAIL.n196 B 0.023643f
C541 VTAIL.n197 B 0.012705f
C542 VTAIL.n198 B 0.013452f
C543 VTAIL.n199 B 0.030029f
C544 VTAIL.n200 B 0.030029f
C545 VTAIL.n201 B 0.013452f
C546 VTAIL.n202 B 0.012705f
C547 VTAIL.n203 B 0.023643f
C548 VTAIL.n204 B 0.061432f
C549 VTAIL.n205 B 0.012705f
C550 VTAIL.n206 B 0.013452f
C551 VTAIL.n207 B 0.060777f
C552 VTAIL.n208 B 0.051626f
C553 VTAIL.n209 B 0.333574f
C554 VTAIL.t18 B 0.337981f
C555 VTAIL.t1 B 0.337981f
C556 VTAIL.n210 B 3.0252f
C557 VTAIL.n211 B 0.529412f
C558 VTAIL.t5 B 0.337981f
C559 VTAIL.t19 B 0.337981f
C560 VTAIL.n212 B 3.0252f
C561 VTAIL.n213 B 0.585236f
C562 VTAIL.n214 B 0.013335f
C563 VTAIL.n215 B 0.030029f
C564 VTAIL.n216 B 0.013452f
C565 VTAIL.n217 B 0.023643f
C566 VTAIL.n218 B 0.012705f
C567 VTAIL.n219 B 0.030029f
C568 VTAIL.n220 B 0.013452f
C569 VTAIL.n221 B 0.023643f
C570 VTAIL.n222 B 0.012705f
C571 VTAIL.n223 B 0.030029f
C572 VTAIL.n224 B 0.013452f
C573 VTAIL.n225 B 0.023643f
C574 VTAIL.n226 B 0.012705f
C575 VTAIL.n227 B 0.030029f
C576 VTAIL.n228 B 0.013452f
C577 VTAIL.n229 B 0.023643f
C578 VTAIL.n230 B 0.012705f
C579 VTAIL.n231 B 0.030029f
C580 VTAIL.n232 B 0.013452f
C581 VTAIL.n233 B 0.023643f
C582 VTAIL.n234 B 0.012705f
C583 VTAIL.n235 B 0.030029f
C584 VTAIL.n236 B 0.013452f
C585 VTAIL.n237 B 0.023643f
C586 VTAIL.n238 B 0.012705f
C587 VTAIL.n239 B 0.030029f
C588 VTAIL.n240 B 0.030029f
C589 VTAIL.n241 B 0.013452f
C590 VTAIL.n242 B 0.023643f
C591 VTAIL.n243 B 0.012705f
C592 VTAIL.n244 B 0.030029f
C593 VTAIL.n245 B 0.013452f
C594 VTAIL.n246 B 0.225741f
C595 VTAIL.t2 B 0.051493f
C596 VTAIL.n247 B 0.022522f
C597 VTAIL.n248 B 0.021228f
C598 VTAIL.n249 B 0.012705f
C599 VTAIL.n250 B 1.83317f
C600 VTAIL.n251 B 0.023643f
C601 VTAIL.n252 B 0.012705f
C602 VTAIL.n253 B 0.013452f
C603 VTAIL.n254 B 0.030029f
C604 VTAIL.n255 B 0.030029f
C605 VTAIL.n256 B 0.013452f
C606 VTAIL.n257 B 0.012705f
C607 VTAIL.n258 B 0.023643f
C608 VTAIL.n259 B 0.023643f
C609 VTAIL.n260 B 0.012705f
C610 VTAIL.n261 B 0.013452f
C611 VTAIL.n262 B 0.030029f
C612 VTAIL.n263 B 0.030029f
C613 VTAIL.n264 B 0.013452f
C614 VTAIL.n265 B 0.012705f
C615 VTAIL.n266 B 0.023643f
C616 VTAIL.n267 B 0.023643f
C617 VTAIL.n268 B 0.012705f
C618 VTAIL.n269 B 0.013078f
C619 VTAIL.n270 B 0.013078f
C620 VTAIL.n271 B 0.030029f
C621 VTAIL.n272 B 0.030029f
C622 VTAIL.n273 B 0.013452f
C623 VTAIL.n274 B 0.012705f
C624 VTAIL.n275 B 0.023643f
C625 VTAIL.n276 B 0.023643f
C626 VTAIL.n277 B 0.012705f
C627 VTAIL.n278 B 0.013452f
C628 VTAIL.n279 B 0.030029f
C629 VTAIL.n280 B 0.030029f
C630 VTAIL.n281 B 0.013452f
C631 VTAIL.n282 B 0.012705f
C632 VTAIL.n283 B 0.023643f
C633 VTAIL.n284 B 0.023643f
C634 VTAIL.n285 B 0.012705f
C635 VTAIL.n286 B 0.013452f
C636 VTAIL.n287 B 0.030029f
C637 VTAIL.n288 B 0.030029f
C638 VTAIL.n289 B 0.013452f
C639 VTAIL.n290 B 0.012705f
C640 VTAIL.n291 B 0.023643f
C641 VTAIL.n292 B 0.023643f
C642 VTAIL.n293 B 0.012705f
C643 VTAIL.n294 B 0.013452f
C644 VTAIL.n295 B 0.030029f
C645 VTAIL.n296 B 0.030029f
C646 VTAIL.n297 B 0.013452f
C647 VTAIL.n298 B 0.012705f
C648 VTAIL.n299 B 0.023643f
C649 VTAIL.n300 B 0.023643f
C650 VTAIL.n301 B 0.012705f
C651 VTAIL.n302 B 0.013452f
C652 VTAIL.n303 B 0.030029f
C653 VTAIL.n304 B 0.030029f
C654 VTAIL.n305 B 0.013452f
C655 VTAIL.n306 B 0.012705f
C656 VTAIL.n307 B 0.023643f
C657 VTAIL.n308 B 0.061432f
C658 VTAIL.n309 B 0.012705f
C659 VTAIL.n310 B 0.013452f
C660 VTAIL.n311 B 0.060777f
C661 VTAIL.n312 B 0.051626f
C662 VTAIL.n313 B 1.89861f
C663 VTAIL.n314 B 0.013335f
C664 VTAIL.n315 B 0.030029f
C665 VTAIL.n316 B 0.013452f
C666 VTAIL.n317 B 0.023643f
C667 VTAIL.n318 B 0.012705f
C668 VTAIL.n319 B 0.030029f
C669 VTAIL.n320 B 0.013452f
C670 VTAIL.n321 B 0.023643f
C671 VTAIL.n322 B 0.012705f
C672 VTAIL.n323 B 0.030029f
C673 VTAIL.n324 B 0.013452f
C674 VTAIL.n325 B 0.023643f
C675 VTAIL.n326 B 0.012705f
C676 VTAIL.n327 B 0.030029f
C677 VTAIL.n328 B 0.013452f
C678 VTAIL.n329 B 0.023643f
C679 VTAIL.n330 B 0.012705f
C680 VTAIL.n331 B 0.030029f
C681 VTAIL.n332 B 0.013452f
C682 VTAIL.n333 B 0.023643f
C683 VTAIL.n334 B 0.012705f
C684 VTAIL.n335 B 0.030029f
C685 VTAIL.n336 B 0.013452f
C686 VTAIL.n337 B 0.023643f
C687 VTAIL.n338 B 0.012705f
C688 VTAIL.n339 B 0.030029f
C689 VTAIL.n340 B 0.013452f
C690 VTAIL.n341 B 0.023643f
C691 VTAIL.n342 B 0.012705f
C692 VTAIL.n343 B 0.030029f
C693 VTAIL.n344 B 0.013452f
C694 VTAIL.n345 B 0.225741f
C695 VTAIL.t8 B 0.051493f
C696 VTAIL.n346 B 0.022522f
C697 VTAIL.n347 B 0.021228f
C698 VTAIL.n348 B 0.012705f
C699 VTAIL.n349 B 1.83317f
C700 VTAIL.n350 B 0.023643f
C701 VTAIL.n351 B 0.012705f
C702 VTAIL.n352 B 0.013452f
C703 VTAIL.n353 B 0.030029f
C704 VTAIL.n354 B 0.030029f
C705 VTAIL.n355 B 0.013452f
C706 VTAIL.n356 B 0.012705f
C707 VTAIL.n357 B 0.023643f
C708 VTAIL.n358 B 0.023643f
C709 VTAIL.n359 B 0.012705f
C710 VTAIL.n360 B 0.013452f
C711 VTAIL.n361 B 0.030029f
C712 VTAIL.n362 B 0.030029f
C713 VTAIL.n363 B 0.030029f
C714 VTAIL.n364 B 0.013452f
C715 VTAIL.n365 B 0.012705f
C716 VTAIL.n366 B 0.023643f
C717 VTAIL.n367 B 0.023643f
C718 VTAIL.n368 B 0.012705f
C719 VTAIL.n369 B 0.013078f
C720 VTAIL.n370 B 0.013078f
C721 VTAIL.n371 B 0.030029f
C722 VTAIL.n372 B 0.030029f
C723 VTAIL.n373 B 0.013452f
C724 VTAIL.n374 B 0.012705f
C725 VTAIL.n375 B 0.023643f
C726 VTAIL.n376 B 0.023643f
C727 VTAIL.n377 B 0.012705f
C728 VTAIL.n378 B 0.013452f
C729 VTAIL.n379 B 0.030029f
C730 VTAIL.n380 B 0.030029f
C731 VTAIL.n381 B 0.013452f
C732 VTAIL.n382 B 0.012705f
C733 VTAIL.n383 B 0.023643f
C734 VTAIL.n384 B 0.023643f
C735 VTAIL.n385 B 0.012705f
C736 VTAIL.n386 B 0.013452f
C737 VTAIL.n387 B 0.030029f
C738 VTAIL.n388 B 0.030029f
C739 VTAIL.n389 B 0.013452f
C740 VTAIL.n390 B 0.012705f
C741 VTAIL.n391 B 0.023643f
C742 VTAIL.n392 B 0.023643f
C743 VTAIL.n393 B 0.012705f
C744 VTAIL.n394 B 0.013452f
C745 VTAIL.n395 B 0.030029f
C746 VTAIL.n396 B 0.030029f
C747 VTAIL.n397 B 0.013452f
C748 VTAIL.n398 B 0.012705f
C749 VTAIL.n399 B 0.023643f
C750 VTAIL.n400 B 0.023643f
C751 VTAIL.n401 B 0.012705f
C752 VTAIL.n402 B 0.013452f
C753 VTAIL.n403 B 0.030029f
C754 VTAIL.n404 B 0.030029f
C755 VTAIL.n405 B 0.013452f
C756 VTAIL.n406 B 0.012705f
C757 VTAIL.n407 B 0.023643f
C758 VTAIL.n408 B 0.061432f
C759 VTAIL.n409 B 0.012705f
C760 VTAIL.n410 B 0.013452f
C761 VTAIL.n411 B 0.060777f
C762 VTAIL.n412 B 0.051626f
C763 VTAIL.n413 B 1.89861f
C764 VTAIL.t14 B 0.337981f
C765 VTAIL.t16 B 0.337981f
C766 VTAIL.n414 B 3.02519f
C767 VTAIL.n415 B 0.443385f
C768 VDD2.n0 B 0.013204f
C769 VDD2.n1 B 0.029733f
C770 VDD2.n2 B 0.013319f
C771 VDD2.n3 B 0.02341f
C772 VDD2.n4 B 0.012579f
C773 VDD2.n5 B 0.029733f
C774 VDD2.n6 B 0.013319f
C775 VDD2.n7 B 0.02341f
C776 VDD2.n8 B 0.012579f
C777 VDD2.n9 B 0.029733f
C778 VDD2.n10 B 0.013319f
C779 VDD2.n11 B 0.02341f
C780 VDD2.n12 B 0.012579f
C781 VDD2.n13 B 0.029733f
C782 VDD2.n14 B 0.013319f
C783 VDD2.n15 B 0.02341f
C784 VDD2.n16 B 0.012579f
C785 VDD2.n17 B 0.029733f
C786 VDD2.n18 B 0.013319f
C787 VDD2.n19 B 0.02341f
C788 VDD2.n20 B 0.012579f
C789 VDD2.n21 B 0.029733f
C790 VDD2.n22 B 0.013319f
C791 VDD2.n23 B 0.02341f
C792 VDD2.n24 B 0.012579f
C793 VDD2.n25 B 0.029733f
C794 VDD2.n26 B 0.013319f
C795 VDD2.n27 B 0.02341f
C796 VDD2.n28 B 0.012579f
C797 VDD2.n29 B 0.029733f
C798 VDD2.n30 B 0.013319f
C799 VDD2.n31 B 0.223514f
C800 VDD2.t3 B 0.050985f
C801 VDD2.n32 B 0.0223f
C802 VDD2.n33 B 0.021019f
C803 VDD2.n34 B 0.012579f
C804 VDD2.n35 B 1.81509f
C805 VDD2.n36 B 0.02341f
C806 VDD2.n37 B 0.012579f
C807 VDD2.n38 B 0.013319f
C808 VDD2.n39 B 0.029733f
C809 VDD2.n40 B 0.029733f
C810 VDD2.n41 B 0.013319f
C811 VDD2.n42 B 0.012579f
C812 VDD2.n43 B 0.02341f
C813 VDD2.n44 B 0.02341f
C814 VDD2.n45 B 0.012579f
C815 VDD2.n46 B 0.013319f
C816 VDD2.n47 B 0.029733f
C817 VDD2.n48 B 0.029733f
C818 VDD2.n49 B 0.029733f
C819 VDD2.n50 B 0.013319f
C820 VDD2.n51 B 0.012579f
C821 VDD2.n52 B 0.02341f
C822 VDD2.n53 B 0.02341f
C823 VDD2.n54 B 0.012579f
C824 VDD2.n55 B 0.012949f
C825 VDD2.n56 B 0.012949f
C826 VDD2.n57 B 0.029733f
C827 VDD2.n58 B 0.029733f
C828 VDD2.n59 B 0.013319f
C829 VDD2.n60 B 0.012579f
C830 VDD2.n61 B 0.02341f
C831 VDD2.n62 B 0.02341f
C832 VDD2.n63 B 0.012579f
C833 VDD2.n64 B 0.013319f
C834 VDD2.n65 B 0.029733f
C835 VDD2.n66 B 0.029733f
C836 VDD2.n67 B 0.013319f
C837 VDD2.n68 B 0.012579f
C838 VDD2.n69 B 0.02341f
C839 VDD2.n70 B 0.02341f
C840 VDD2.n71 B 0.012579f
C841 VDD2.n72 B 0.013319f
C842 VDD2.n73 B 0.029733f
C843 VDD2.n74 B 0.029733f
C844 VDD2.n75 B 0.013319f
C845 VDD2.n76 B 0.012579f
C846 VDD2.n77 B 0.02341f
C847 VDD2.n78 B 0.02341f
C848 VDD2.n79 B 0.012579f
C849 VDD2.n80 B 0.013319f
C850 VDD2.n81 B 0.029733f
C851 VDD2.n82 B 0.029733f
C852 VDD2.n83 B 0.013319f
C853 VDD2.n84 B 0.012579f
C854 VDD2.n85 B 0.02341f
C855 VDD2.n86 B 0.02341f
C856 VDD2.n87 B 0.012579f
C857 VDD2.n88 B 0.013319f
C858 VDD2.n89 B 0.029733f
C859 VDD2.n90 B 0.029733f
C860 VDD2.n91 B 0.013319f
C861 VDD2.n92 B 0.012579f
C862 VDD2.n93 B 0.02341f
C863 VDD2.n94 B 0.060826f
C864 VDD2.n95 B 0.012579f
C865 VDD2.n96 B 0.013319f
C866 VDD2.n97 B 0.060177f
C867 VDD2.n98 B 0.077423f
C868 VDD2.t4 B 0.334648f
C869 VDD2.t0 B 0.334648f
C870 VDD2.n99 B 3.05876f
C871 VDD2.n100 B 0.627706f
C872 VDD2.t5 B 0.334648f
C873 VDD2.t8 B 0.334648f
C874 VDD2.n101 B 3.07223f
C875 VDD2.n102 B 3.00186f
C876 VDD2.n103 B 0.013204f
C877 VDD2.n104 B 0.029733f
C878 VDD2.n105 B 0.013319f
C879 VDD2.n106 B 0.02341f
C880 VDD2.n107 B 0.012579f
C881 VDD2.n108 B 0.029733f
C882 VDD2.n109 B 0.013319f
C883 VDD2.n110 B 0.02341f
C884 VDD2.n111 B 0.012579f
C885 VDD2.n112 B 0.029733f
C886 VDD2.n113 B 0.013319f
C887 VDD2.n114 B 0.02341f
C888 VDD2.n115 B 0.012579f
C889 VDD2.n116 B 0.029733f
C890 VDD2.n117 B 0.013319f
C891 VDD2.n118 B 0.02341f
C892 VDD2.n119 B 0.012579f
C893 VDD2.n120 B 0.029733f
C894 VDD2.n121 B 0.013319f
C895 VDD2.n122 B 0.02341f
C896 VDD2.n123 B 0.012579f
C897 VDD2.n124 B 0.029733f
C898 VDD2.n125 B 0.013319f
C899 VDD2.n126 B 0.02341f
C900 VDD2.n127 B 0.012579f
C901 VDD2.n128 B 0.029733f
C902 VDD2.n129 B 0.029733f
C903 VDD2.n130 B 0.013319f
C904 VDD2.n131 B 0.02341f
C905 VDD2.n132 B 0.012579f
C906 VDD2.n133 B 0.029733f
C907 VDD2.n134 B 0.013319f
C908 VDD2.n135 B 0.223514f
C909 VDD2.t7 B 0.050985f
C910 VDD2.n136 B 0.0223f
C911 VDD2.n137 B 0.021019f
C912 VDD2.n138 B 0.012579f
C913 VDD2.n139 B 1.81509f
C914 VDD2.n140 B 0.02341f
C915 VDD2.n141 B 0.012579f
C916 VDD2.n142 B 0.013319f
C917 VDD2.n143 B 0.029733f
C918 VDD2.n144 B 0.029733f
C919 VDD2.n145 B 0.013319f
C920 VDD2.n146 B 0.012579f
C921 VDD2.n147 B 0.02341f
C922 VDD2.n148 B 0.02341f
C923 VDD2.n149 B 0.012579f
C924 VDD2.n150 B 0.013319f
C925 VDD2.n151 B 0.029733f
C926 VDD2.n152 B 0.029733f
C927 VDD2.n153 B 0.013319f
C928 VDD2.n154 B 0.012579f
C929 VDD2.n155 B 0.02341f
C930 VDD2.n156 B 0.02341f
C931 VDD2.n157 B 0.012579f
C932 VDD2.n158 B 0.012949f
C933 VDD2.n159 B 0.012949f
C934 VDD2.n160 B 0.029733f
C935 VDD2.n161 B 0.029733f
C936 VDD2.n162 B 0.013319f
C937 VDD2.n163 B 0.012579f
C938 VDD2.n164 B 0.02341f
C939 VDD2.n165 B 0.02341f
C940 VDD2.n166 B 0.012579f
C941 VDD2.n167 B 0.013319f
C942 VDD2.n168 B 0.029733f
C943 VDD2.n169 B 0.029733f
C944 VDD2.n170 B 0.013319f
C945 VDD2.n171 B 0.012579f
C946 VDD2.n172 B 0.02341f
C947 VDD2.n173 B 0.02341f
C948 VDD2.n174 B 0.012579f
C949 VDD2.n175 B 0.013319f
C950 VDD2.n176 B 0.029733f
C951 VDD2.n177 B 0.029733f
C952 VDD2.n178 B 0.013319f
C953 VDD2.n179 B 0.012579f
C954 VDD2.n180 B 0.02341f
C955 VDD2.n181 B 0.02341f
C956 VDD2.n182 B 0.012579f
C957 VDD2.n183 B 0.013319f
C958 VDD2.n184 B 0.029733f
C959 VDD2.n185 B 0.029733f
C960 VDD2.n186 B 0.013319f
C961 VDD2.n187 B 0.012579f
C962 VDD2.n188 B 0.02341f
C963 VDD2.n189 B 0.02341f
C964 VDD2.n190 B 0.012579f
C965 VDD2.n191 B 0.013319f
C966 VDD2.n192 B 0.029733f
C967 VDD2.n193 B 0.029733f
C968 VDD2.n194 B 0.013319f
C969 VDD2.n195 B 0.012579f
C970 VDD2.n196 B 0.02341f
C971 VDD2.n197 B 0.060826f
C972 VDD2.n198 B 0.012579f
C973 VDD2.n199 B 0.013319f
C974 VDD2.n200 B 0.060177f
C975 VDD2.n201 B 0.067246f
C976 VDD2.n202 B 3.09322f
C977 VDD2.t1 B 0.334648f
C978 VDD2.t2 B 0.334648f
C979 VDD2.n203 B 3.05876f
C980 VDD2.n204 B 0.416199f
C981 VDD2.t6 B 0.334648f
C982 VDD2.t9 B 0.334648f
C983 VDD2.n205 B 3.0722f
C984 VN.n0 B 0.02809f
C985 VN.t8 B 2.60824f
C986 VN.n1 B 0.034965f
C987 VN.n2 B 0.021306f
C988 VN.t0 B 2.60824f
C989 VN.n3 B 0.90534f
C990 VN.n4 B 0.021306f
C991 VN.n5 B 0.038898f
C992 VN.n6 B 0.021306f
C993 VN.t2 B 2.60824f
C994 VN.n7 B 0.038898f
C995 VN.n8 B 0.021306f
C996 VN.t9 B 2.60824f
C997 VN.n9 B 0.966341f
C998 VN.t3 B 2.76447f
C999 VN.n10 B 0.953352f
C1000 VN.n11 B 0.202293f
C1001 VN.n12 B 0.031476f
C1002 VN.n13 B 0.042576f
C1003 VN.n14 B 0.020446f
C1004 VN.n15 B 0.021306f
C1005 VN.n16 B 0.021306f
C1006 VN.n17 B 0.021306f
C1007 VN.n18 B 0.03971f
C1008 VN.n19 B 0.925445f
C1009 VN.n20 B 0.03971f
C1010 VN.n21 B 0.021306f
C1011 VN.n22 B 0.021306f
C1012 VN.n23 B 0.021306f
C1013 VN.n24 B 0.020446f
C1014 VN.n25 B 0.042576f
C1015 VN.n26 B 0.031476f
C1016 VN.n27 B 0.021306f
C1017 VN.n28 B 0.021306f
C1018 VN.n29 B 0.028339f
C1019 VN.n30 B 0.03971f
C1020 VN.n31 B 0.027246f
C1021 VN.n32 B 0.021306f
C1022 VN.n33 B 0.021306f
C1023 VN.n34 B 0.021306f
C1024 VN.n35 B 0.03971f
C1025 VN.n36 B 0.023242f
C1026 VN.n37 B 0.966025f
C1027 VN.n38 B 0.036452f
C1028 VN.n39 B 0.02809f
C1029 VN.t5 B 2.60824f
C1030 VN.n40 B 0.034965f
C1031 VN.n41 B 0.021306f
C1032 VN.t1 B 2.60824f
C1033 VN.n42 B 0.90534f
C1034 VN.n43 B 0.021306f
C1035 VN.n44 B 0.038898f
C1036 VN.n45 B 0.021306f
C1037 VN.t4 B 2.60824f
C1038 VN.n46 B 0.038898f
C1039 VN.n47 B 0.021306f
C1040 VN.t6 B 2.60824f
C1041 VN.n48 B 0.966341f
C1042 VN.t7 B 2.76447f
C1043 VN.n49 B 0.953352f
C1044 VN.n50 B 0.202293f
C1045 VN.n51 B 0.031476f
C1046 VN.n52 B 0.042576f
C1047 VN.n53 B 0.020446f
C1048 VN.n54 B 0.021306f
C1049 VN.n55 B 0.021306f
C1050 VN.n56 B 0.021306f
C1051 VN.n57 B 0.03971f
C1052 VN.n58 B 0.925445f
C1053 VN.n59 B 0.03971f
C1054 VN.n60 B 0.021306f
C1055 VN.n61 B 0.021306f
C1056 VN.n62 B 0.021306f
C1057 VN.n63 B 0.020446f
C1058 VN.n64 B 0.042576f
C1059 VN.n65 B 0.031476f
C1060 VN.n66 B 0.021306f
C1061 VN.n67 B 0.021306f
C1062 VN.n68 B 0.028339f
C1063 VN.n69 B 0.03971f
C1064 VN.n70 B 0.027246f
C1065 VN.n71 B 0.021306f
C1066 VN.n72 B 0.021306f
C1067 VN.n73 B 0.021306f
C1068 VN.n74 B 0.03971f
C1069 VN.n75 B 0.023242f
C1070 VN.n76 B 0.966025f
C1071 VN.n77 B 1.43617f
.ends

