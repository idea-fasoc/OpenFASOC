VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_4K
  CLASS BLOCK ;
  FOREIGN DFFRAM_4K ;
  ORIGIN 0.000 0.000 ;
  SIZE 1089.845 BY 1389.360 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.960 1385.360 441.240 1389.360 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.760 1385.360 455.040 1389.360 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.560 1385.360 468.840 1389.360 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.360 1385.360 482.640 1389.360 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.700 1385.360 495.980 1389.360 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.500 1385.360 509.780 1389.360 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.300 1385.360 523.580 1389.360 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.100 1385.360 537.380 1389.360 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.900 1385.360 551.180 1389.360 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.700 1385.360 564.980 1389.360 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.500 1385.360 578.780 1389.360 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.840 1385.360 661.120 1389.360 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.380 1385.360 798.660 1389.360 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.180 1385.360 812.460 1389.360 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.980 1385.360 826.260 1389.360 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.780 1385.360 840.060 1389.360 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.580 1385.360 853.860 1389.360 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.920 1385.360 867.200 1389.360 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.720 1385.360 881.000 1389.360 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.520 1385.360 894.800 1389.360 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.320 1385.360 908.600 1389.360 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.120 1385.360 922.400 1389.360 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.640 1385.360 674.920 1389.360 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.920 1385.360 936.200 1389.360 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.720 1385.360 950.000 1389.360 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.520 1385.360 963.800 1389.360 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.320 1385.360 977.600 1389.360 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.660 1385.360 990.940 1389.360 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.460 1385.360 1004.740 1389.360 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.260 1385.360 1018.540 1389.360 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.060 1385.360 1032.340 1389.360 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.860 1385.360 1046.140 1389.360 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.660 1385.360 1059.940 1389.360 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.440 1385.360 688.720 1389.360 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.460 1385.360 1073.740 1389.360 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.260 1385.360 1087.540 1389.360 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.240 1385.360 702.520 1389.360 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.040 1385.360 716.320 1389.360 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.840 1385.360 730.120 1389.360 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.180 1385.360 743.460 1389.360 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.980 1385.360 757.260 1389.360 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.780 1385.360 771.060 1389.360 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.580 1385.360 784.860 1389.360 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.200 1385.360 1.480 1389.360 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.280 1385.360 138.560 1389.360 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.080 1385.360 152.360 1389.360 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.880 1385.360 166.160 1389.360 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.680 1385.360 179.960 1389.360 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.480 1385.360 193.760 1389.360 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.280 1385.360 207.560 1389.360 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.080 1385.360 221.360 1389.360 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.880 1385.360 235.160 1389.360 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.220 1385.360 248.500 1389.360 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.020 1385.360 262.300 1389.360 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.540 1385.360 14.820 1389.360 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.820 1385.360 276.100 1389.360 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.620 1385.360 289.900 1389.360 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.420 1385.360 303.700 1389.360 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.220 1385.360 317.500 1389.360 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.020 1385.360 331.300 1389.360 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.820 1385.360 345.100 1389.360 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.620 1385.360 358.900 1389.360 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.960 1385.360 372.240 1389.360 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.760 1385.360 386.040 1389.360 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.560 1385.360 399.840 1389.360 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.340 1385.360 28.620 1389.360 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.360 1385.360 413.640 1389.360 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.160 1385.360 427.440 1389.360 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.140 1385.360 42.420 1389.360 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.940 1385.360 56.220 1389.360 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.740 1385.360 70.020 1389.360 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.540 1385.360 83.820 1389.360 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.340 1385.360 97.620 1389.360 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.140 1385.360 111.420 1389.360 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.480 1385.360 124.760 1389.360 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.040 1385.360 647.320 1389.360 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.300 1385.360 592.580 1389.360 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.100 1385.360 606.380 1389.360 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.440 1385.360 619.720 1389.360 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.240 1385.360 633.520 1389.360 ;
    END
  END WE[3]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 937.310 0.000 938.910 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.710 0.000 785.310 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 630.110 0.000 631.710 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 476.510 0.000 478.110 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 322.910 0.000 324.510 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 169.310 0.000 170.910 1376.800 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.710 0.000 17.310 1376.800 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1014.110 0.000 1015.710 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 860.510 0.000 862.110 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 706.910 0.000 708.510 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 553.310 0.000 554.910 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 399.710 0.000 401.310 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.110 0.000 247.710 1376.800 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 92.510 0.000 94.110 1376.800 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 0.190 0.155 1089.785 1376.645 ;
      LAYER met1 ;
        RECT 0.190 0.000 1089.845 1380.260 ;
      LAYER met2 ;
        RECT 1.760 1385.080 14.260 1385.360 ;
        RECT 15.100 1385.080 28.060 1385.360 ;
        RECT 28.900 1385.080 41.860 1385.360 ;
        RECT 42.700 1385.080 55.660 1385.360 ;
        RECT 56.500 1385.080 69.460 1385.360 ;
        RECT 70.300 1385.080 83.260 1385.360 ;
        RECT 84.100 1385.080 97.060 1385.360 ;
        RECT 97.900 1385.080 110.860 1385.360 ;
        RECT 111.700 1385.080 124.200 1385.360 ;
        RECT 125.040 1385.080 138.000 1385.360 ;
        RECT 138.840 1385.080 151.800 1385.360 ;
        RECT 152.640 1385.080 165.600 1385.360 ;
        RECT 166.440 1385.080 179.400 1385.360 ;
        RECT 180.240 1385.080 193.200 1385.360 ;
        RECT 194.040 1385.080 207.000 1385.360 ;
        RECT 207.840 1385.080 220.800 1385.360 ;
        RECT 221.640 1385.080 234.600 1385.360 ;
        RECT 235.440 1385.080 247.940 1385.360 ;
        RECT 248.780 1385.080 261.740 1385.360 ;
        RECT 262.580 1385.080 275.540 1385.360 ;
        RECT 276.380 1385.080 289.340 1385.360 ;
        RECT 290.180 1385.080 303.140 1385.360 ;
        RECT 303.980 1385.080 316.940 1385.360 ;
        RECT 317.780 1385.080 330.740 1385.360 ;
        RECT 331.580 1385.080 344.540 1385.360 ;
        RECT 345.380 1385.080 358.340 1385.360 ;
        RECT 359.180 1385.080 371.680 1385.360 ;
        RECT 372.520 1385.080 385.480 1385.360 ;
        RECT 386.320 1385.080 399.280 1385.360 ;
        RECT 400.120 1385.080 413.080 1385.360 ;
        RECT 413.920 1385.080 426.880 1385.360 ;
        RECT 427.720 1385.080 440.680 1385.360 ;
        RECT 441.520 1385.080 454.480 1385.360 ;
        RECT 455.320 1385.080 468.280 1385.360 ;
        RECT 469.120 1385.080 482.080 1385.360 ;
        RECT 482.920 1385.080 495.420 1385.360 ;
        RECT 496.260 1385.080 509.220 1385.360 ;
        RECT 510.060 1385.080 523.020 1385.360 ;
        RECT 523.860 1385.080 536.820 1385.360 ;
        RECT 537.660 1385.080 550.620 1385.360 ;
        RECT 551.460 1385.080 564.420 1385.360 ;
        RECT 565.260 1385.080 578.220 1385.360 ;
        RECT 579.060 1385.080 592.020 1385.360 ;
        RECT 592.860 1385.080 605.820 1385.360 ;
        RECT 606.660 1385.080 619.160 1385.360 ;
        RECT 620.000 1385.080 632.960 1385.360 ;
        RECT 633.800 1385.080 646.760 1385.360 ;
        RECT 647.600 1385.080 660.560 1385.360 ;
        RECT 661.400 1385.080 674.360 1385.360 ;
        RECT 675.200 1385.080 688.160 1385.360 ;
        RECT 689.000 1385.080 701.960 1385.360 ;
        RECT 702.800 1385.080 715.760 1385.360 ;
        RECT 716.600 1385.080 729.560 1385.360 ;
        RECT 730.400 1385.080 742.900 1385.360 ;
        RECT 743.740 1385.080 756.700 1385.360 ;
        RECT 757.540 1385.080 770.500 1385.360 ;
        RECT 771.340 1385.080 784.300 1385.360 ;
        RECT 785.140 1385.080 798.100 1385.360 ;
        RECT 798.940 1385.080 811.900 1385.360 ;
        RECT 812.740 1385.080 825.700 1385.360 ;
        RECT 826.540 1385.080 839.500 1385.360 ;
        RECT 840.340 1385.080 853.300 1385.360 ;
        RECT 854.140 1385.080 866.640 1385.360 ;
        RECT 867.480 1385.080 880.440 1385.360 ;
        RECT 881.280 1385.080 894.240 1385.360 ;
        RECT 895.080 1385.080 908.040 1385.360 ;
        RECT 908.880 1385.080 921.840 1385.360 ;
        RECT 922.680 1385.080 935.640 1385.360 ;
        RECT 936.480 1385.080 949.440 1385.360 ;
        RECT 950.280 1385.080 963.240 1385.360 ;
        RECT 964.080 1385.080 977.040 1385.360 ;
        RECT 977.880 1385.080 990.380 1385.360 ;
        RECT 991.220 1385.080 1004.180 1385.360 ;
        RECT 1005.020 1385.080 1017.980 1385.360 ;
        RECT 1018.820 1385.080 1031.780 1385.360 ;
        RECT 1032.620 1385.080 1045.580 1385.360 ;
        RECT 1046.420 1385.080 1059.380 1385.360 ;
        RECT 1060.220 1385.080 1073.180 1385.360 ;
        RECT 1074.020 1385.080 1086.980 1385.360 ;
        RECT 1087.820 1385.080 1088.000 1385.360 ;
        RECT 1.210 0.000 1088.000 1385.080 ;
      LAYER met3 ;
        RECT 1.635 0.075 1088.025 1376.725 ;
      LAYER met4 ;
        RECT 11.525 19.455 15.310 1375.025 ;
        RECT 17.710 19.455 92.110 1375.025 ;
        RECT 94.510 19.455 168.910 1375.025 ;
        RECT 171.310 19.455 245.710 1375.025 ;
        RECT 248.110 19.455 322.510 1375.025 ;
        RECT 324.910 19.455 399.310 1375.025 ;
        RECT 401.710 19.455 476.110 1375.025 ;
        RECT 478.510 19.455 552.910 1375.025 ;
        RECT 555.310 19.455 629.710 1375.025 ;
        RECT 632.110 19.455 706.510 1375.025 ;
        RECT 708.910 19.455 783.310 1375.025 ;
        RECT 785.710 19.455 860.110 1375.025 ;
        RECT 862.510 19.455 936.910 1375.025 ;
        RECT 939.310 19.455 1013.710 1375.025 ;
        RECT 1016.110 19.455 1069.855 1375.025 ;
  END
END DFFRAM_4K
END LIBRARY
