* NGSPICE file created from diff_pair_sample_0110.ext - technology: sky130A

.subckt diff_pair_sample_0110 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=3.51
X1 VTAIL.t2 VP.t0 VDD1.t7 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X2 VTAIL.t6 VP.t1 VDD1.t6 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X3 VTAIL.t13 VN.t1 VDD2.t6 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=3.51
X4 VDD2.t5 VN.t2 VTAIL.t10 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X5 B.t11 B.t9 B.t10 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=3.51
X6 VDD2.t4 VN.t3 VTAIL.t11 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X7 B.t8 B.t6 B.t7 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=3.51
X8 B.t5 B.t3 B.t4 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=3.51
X9 VDD2.t3 VN.t4 VTAIL.t8 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=3.51
X10 B.t2 B.t0 B.t1 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=0 ps=0 w=17.64 l=3.51
X11 VDD1.t5 VP.t2 VTAIL.t5 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X12 VTAIL.t15 VN.t5 VDD2.t2 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X13 VDD1.t4 VP.t3 VTAIL.t0 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=3.51
X14 VDD1.t3 VP.t4 VTAIL.t4 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X15 VTAIL.t12 VN.t6 VDD2.t1 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=2.9106 ps=17.97 w=17.64 l=3.51
X16 VTAIL.t9 VN.t7 VDD2.t0 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=3.51
X17 VTAIL.t3 VP.t5 VDD1.t2 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=3.51
X18 VDD1.t1 VP.t6 VTAIL.t7 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=2.9106 pd=17.97 as=6.8796 ps=36.06 w=17.64 l=3.51
X19 VTAIL.t1 VP.t7 VDD1.t0 w_n4810_n4496# sky130_fd_pr__pfet_01v8 ad=6.8796 pd=36.06 as=2.9106 ps=17.97 w=17.64 l=3.51
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n39 161.3
R8 VN.n56 VN.n55 161.3
R9 VN.n54 VN.n40 161.3
R10 VN.n53 VN.n52 161.3
R11 VN.n51 VN.n42 161.3
R12 VN.n50 VN.n49 161.3
R13 VN.n48 VN.n43 161.3
R14 VN.n47 VN.n46 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n4 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n18 VN.n5 161.3
R25 VN.n17 VN.n16 161.3
R26 VN.n15 VN.n6 161.3
R27 VN.n14 VN.n13 161.3
R28 VN.n12 VN.n7 161.3
R29 VN.n11 VN.n10 161.3
R30 VN.n45 VN.t4 154.982
R31 VN.n9 VN.t7 154.982
R32 VN.n8 VN.t2 121.118
R33 VN.n19 VN.t6 121.118
R34 VN.n0 VN.t0 121.118
R35 VN.n44 VN.t5 121.118
R36 VN.n41 VN.t3 121.118
R37 VN.n35 VN.t1 121.118
R38 VN.n34 VN.n0 77.4578
R39 VN.n69 VN.n35 77.4578
R40 VN VN.n69 59.7254
R41 VN.n26 VN.n2 56.0773
R42 VN.n61 VN.n37 56.0773
R43 VN.n45 VN.n44 54.2621
R44 VN.n9 VN.n8 54.2621
R45 VN.n13 VN.n6 40.577
R46 VN.n17 VN.n6 40.577
R47 VN.n49 VN.n42 40.577
R48 VN.n53 VN.n42 40.577
R49 VN.n30 VN.n2 25.0767
R50 VN.n65 VN.n37 25.0767
R51 VN.n12 VN.n11 24.5923
R52 VN.n13 VN.n12 24.5923
R53 VN.n18 VN.n17 24.5923
R54 VN.n20 VN.n18 24.5923
R55 VN.n24 VN.n4 24.5923
R56 VN.n25 VN.n24 24.5923
R57 VN.n26 VN.n25 24.5923
R58 VN.n31 VN.n30 24.5923
R59 VN.n32 VN.n31 24.5923
R60 VN.n49 VN.n48 24.5923
R61 VN.n48 VN.n47 24.5923
R62 VN.n61 VN.n60 24.5923
R63 VN.n60 VN.n59 24.5923
R64 VN.n59 VN.n39 24.5923
R65 VN.n55 VN.n54 24.5923
R66 VN.n54 VN.n53 24.5923
R67 VN.n67 VN.n66 24.5923
R68 VN.n66 VN.n65 24.5923
R69 VN.n11 VN.n8 20.6576
R70 VN.n20 VN.n19 20.6576
R71 VN.n47 VN.n44 20.6576
R72 VN.n55 VN.n41 20.6576
R73 VN.n32 VN.n0 12.7883
R74 VN.n67 VN.n35 12.7883
R75 VN.n19 VN.n4 3.93519
R76 VN.n41 VN.n39 3.93519
R77 VN.n46 VN.n45 3.05448
R78 VN.n10 VN.n9 3.05448
R79 VN.n69 VN.n68 0.354861
R80 VN.n34 VN.n33 0.354861
R81 VN VN.n34 0.267071
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n56 0.189894
R90 VN.n56 VN.n40 0.189894
R91 VN.n52 VN.n40 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n50 0.189894
R94 VN.n50 VN.n43 0.189894
R95 VN.n46 VN.n43 0.189894
R96 VN.n10 VN.n7 0.189894
R97 VN.n14 VN.n7 0.189894
R98 VN.n15 VN.n14 0.189894
R99 VN.n16 VN.n15 0.189894
R100 VN.n16 VN.n5 0.189894
R101 VN.n21 VN.n5 0.189894
R102 VN.n22 VN.n21 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VTAIL.n786 VTAIL.n694 756.745
R111 VTAIL.n94 VTAIL.n2 756.745
R112 VTAIL.n192 VTAIL.n100 756.745
R113 VTAIL.n292 VTAIL.n200 756.745
R114 VTAIL.n688 VTAIL.n596 756.745
R115 VTAIL.n588 VTAIL.n496 756.745
R116 VTAIL.n490 VTAIL.n398 756.745
R117 VTAIL.n390 VTAIL.n298 756.745
R118 VTAIL.n727 VTAIL.n726 585
R119 VTAIL.n729 VTAIL.n728 585
R120 VTAIL.n722 VTAIL.n721 585
R121 VTAIL.n735 VTAIL.n734 585
R122 VTAIL.n737 VTAIL.n736 585
R123 VTAIL.n718 VTAIL.n717 585
R124 VTAIL.n743 VTAIL.n742 585
R125 VTAIL.n745 VTAIL.n744 585
R126 VTAIL.n714 VTAIL.n713 585
R127 VTAIL.n751 VTAIL.n750 585
R128 VTAIL.n753 VTAIL.n752 585
R129 VTAIL.n710 VTAIL.n709 585
R130 VTAIL.n759 VTAIL.n758 585
R131 VTAIL.n761 VTAIL.n760 585
R132 VTAIL.n706 VTAIL.n705 585
R133 VTAIL.n768 VTAIL.n767 585
R134 VTAIL.n769 VTAIL.n704 585
R135 VTAIL.n771 VTAIL.n770 585
R136 VTAIL.n702 VTAIL.n701 585
R137 VTAIL.n777 VTAIL.n776 585
R138 VTAIL.n779 VTAIL.n778 585
R139 VTAIL.n698 VTAIL.n697 585
R140 VTAIL.n785 VTAIL.n784 585
R141 VTAIL.n787 VTAIL.n786 585
R142 VTAIL.n35 VTAIL.n34 585
R143 VTAIL.n37 VTAIL.n36 585
R144 VTAIL.n30 VTAIL.n29 585
R145 VTAIL.n43 VTAIL.n42 585
R146 VTAIL.n45 VTAIL.n44 585
R147 VTAIL.n26 VTAIL.n25 585
R148 VTAIL.n51 VTAIL.n50 585
R149 VTAIL.n53 VTAIL.n52 585
R150 VTAIL.n22 VTAIL.n21 585
R151 VTAIL.n59 VTAIL.n58 585
R152 VTAIL.n61 VTAIL.n60 585
R153 VTAIL.n18 VTAIL.n17 585
R154 VTAIL.n67 VTAIL.n66 585
R155 VTAIL.n69 VTAIL.n68 585
R156 VTAIL.n14 VTAIL.n13 585
R157 VTAIL.n76 VTAIL.n75 585
R158 VTAIL.n77 VTAIL.n12 585
R159 VTAIL.n79 VTAIL.n78 585
R160 VTAIL.n10 VTAIL.n9 585
R161 VTAIL.n85 VTAIL.n84 585
R162 VTAIL.n87 VTAIL.n86 585
R163 VTAIL.n6 VTAIL.n5 585
R164 VTAIL.n93 VTAIL.n92 585
R165 VTAIL.n95 VTAIL.n94 585
R166 VTAIL.n133 VTAIL.n132 585
R167 VTAIL.n135 VTAIL.n134 585
R168 VTAIL.n128 VTAIL.n127 585
R169 VTAIL.n141 VTAIL.n140 585
R170 VTAIL.n143 VTAIL.n142 585
R171 VTAIL.n124 VTAIL.n123 585
R172 VTAIL.n149 VTAIL.n148 585
R173 VTAIL.n151 VTAIL.n150 585
R174 VTAIL.n120 VTAIL.n119 585
R175 VTAIL.n157 VTAIL.n156 585
R176 VTAIL.n159 VTAIL.n158 585
R177 VTAIL.n116 VTAIL.n115 585
R178 VTAIL.n165 VTAIL.n164 585
R179 VTAIL.n167 VTAIL.n166 585
R180 VTAIL.n112 VTAIL.n111 585
R181 VTAIL.n174 VTAIL.n173 585
R182 VTAIL.n175 VTAIL.n110 585
R183 VTAIL.n177 VTAIL.n176 585
R184 VTAIL.n108 VTAIL.n107 585
R185 VTAIL.n183 VTAIL.n182 585
R186 VTAIL.n185 VTAIL.n184 585
R187 VTAIL.n104 VTAIL.n103 585
R188 VTAIL.n191 VTAIL.n190 585
R189 VTAIL.n193 VTAIL.n192 585
R190 VTAIL.n233 VTAIL.n232 585
R191 VTAIL.n235 VTAIL.n234 585
R192 VTAIL.n228 VTAIL.n227 585
R193 VTAIL.n241 VTAIL.n240 585
R194 VTAIL.n243 VTAIL.n242 585
R195 VTAIL.n224 VTAIL.n223 585
R196 VTAIL.n249 VTAIL.n248 585
R197 VTAIL.n251 VTAIL.n250 585
R198 VTAIL.n220 VTAIL.n219 585
R199 VTAIL.n257 VTAIL.n256 585
R200 VTAIL.n259 VTAIL.n258 585
R201 VTAIL.n216 VTAIL.n215 585
R202 VTAIL.n265 VTAIL.n264 585
R203 VTAIL.n267 VTAIL.n266 585
R204 VTAIL.n212 VTAIL.n211 585
R205 VTAIL.n274 VTAIL.n273 585
R206 VTAIL.n275 VTAIL.n210 585
R207 VTAIL.n277 VTAIL.n276 585
R208 VTAIL.n208 VTAIL.n207 585
R209 VTAIL.n283 VTAIL.n282 585
R210 VTAIL.n285 VTAIL.n284 585
R211 VTAIL.n204 VTAIL.n203 585
R212 VTAIL.n291 VTAIL.n290 585
R213 VTAIL.n293 VTAIL.n292 585
R214 VTAIL.n689 VTAIL.n688 585
R215 VTAIL.n687 VTAIL.n686 585
R216 VTAIL.n600 VTAIL.n599 585
R217 VTAIL.n681 VTAIL.n680 585
R218 VTAIL.n679 VTAIL.n678 585
R219 VTAIL.n604 VTAIL.n603 585
R220 VTAIL.n608 VTAIL.n606 585
R221 VTAIL.n673 VTAIL.n672 585
R222 VTAIL.n671 VTAIL.n670 585
R223 VTAIL.n610 VTAIL.n609 585
R224 VTAIL.n665 VTAIL.n664 585
R225 VTAIL.n663 VTAIL.n662 585
R226 VTAIL.n614 VTAIL.n613 585
R227 VTAIL.n657 VTAIL.n656 585
R228 VTAIL.n655 VTAIL.n654 585
R229 VTAIL.n618 VTAIL.n617 585
R230 VTAIL.n649 VTAIL.n648 585
R231 VTAIL.n647 VTAIL.n646 585
R232 VTAIL.n622 VTAIL.n621 585
R233 VTAIL.n641 VTAIL.n640 585
R234 VTAIL.n639 VTAIL.n638 585
R235 VTAIL.n626 VTAIL.n625 585
R236 VTAIL.n633 VTAIL.n632 585
R237 VTAIL.n631 VTAIL.n630 585
R238 VTAIL.n589 VTAIL.n588 585
R239 VTAIL.n587 VTAIL.n586 585
R240 VTAIL.n500 VTAIL.n499 585
R241 VTAIL.n581 VTAIL.n580 585
R242 VTAIL.n579 VTAIL.n578 585
R243 VTAIL.n504 VTAIL.n503 585
R244 VTAIL.n508 VTAIL.n506 585
R245 VTAIL.n573 VTAIL.n572 585
R246 VTAIL.n571 VTAIL.n570 585
R247 VTAIL.n510 VTAIL.n509 585
R248 VTAIL.n565 VTAIL.n564 585
R249 VTAIL.n563 VTAIL.n562 585
R250 VTAIL.n514 VTAIL.n513 585
R251 VTAIL.n557 VTAIL.n556 585
R252 VTAIL.n555 VTAIL.n554 585
R253 VTAIL.n518 VTAIL.n517 585
R254 VTAIL.n549 VTAIL.n548 585
R255 VTAIL.n547 VTAIL.n546 585
R256 VTAIL.n522 VTAIL.n521 585
R257 VTAIL.n541 VTAIL.n540 585
R258 VTAIL.n539 VTAIL.n538 585
R259 VTAIL.n526 VTAIL.n525 585
R260 VTAIL.n533 VTAIL.n532 585
R261 VTAIL.n531 VTAIL.n530 585
R262 VTAIL.n491 VTAIL.n490 585
R263 VTAIL.n489 VTAIL.n488 585
R264 VTAIL.n402 VTAIL.n401 585
R265 VTAIL.n483 VTAIL.n482 585
R266 VTAIL.n481 VTAIL.n480 585
R267 VTAIL.n406 VTAIL.n405 585
R268 VTAIL.n410 VTAIL.n408 585
R269 VTAIL.n475 VTAIL.n474 585
R270 VTAIL.n473 VTAIL.n472 585
R271 VTAIL.n412 VTAIL.n411 585
R272 VTAIL.n467 VTAIL.n466 585
R273 VTAIL.n465 VTAIL.n464 585
R274 VTAIL.n416 VTAIL.n415 585
R275 VTAIL.n459 VTAIL.n458 585
R276 VTAIL.n457 VTAIL.n456 585
R277 VTAIL.n420 VTAIL.n419 585
R278 VTAIL.n451 VTAIL.n450 585
R279 VTAIL.n449 VTAIL.n448 585
R280 VTAIL.n424 VTAIL.n423 585
R281 VTAIL.n443 VTAIL.n442 585
R282 VTAIL.n441 VTAIL.n440 585
R283 VTAIL.n428 VTAIL.n427 585
R284 VTAIL.n435 VTAIL.n434 585
R285 VTAIL.n433 VTAIL.n432 585
R286 VTAIL.n391 VTAIL.n390 585
R287 VTAIL.n389 VTAIL.n388 585
R288 VTAIL.n302 VTAIL.n301 585
R289 VTAIL.n383 VTAIL.n382 585
R290 VTAIL.n381 VTAIL.n380 585
R291 VTAIL.n306 VTAIL.n305 585
R292 VTAIL.n310 VTAIL.n308 585
R293 VTAIL.n375 VTAIL.n374 585
R294 VTAIL.n373 VTAIL.n372 585
R295 VTAIL.n312 VTAIL.n311 585
R296 VTAIL.n367 VTAIL.n366 585
R297 VTAIL.n365 VTAIL.n364 585
R298 VTAIL.n316 VTAIL.n315 585
R299 VTAIL.n359 VTAIL.n358 585
R300 VTAIL.n357 VTAIL.n356 585
R301 VTAIL.n320 VTAIL.n319 585
R302 VTAIL.n351 VTAIL.n350 585
R303 VTAIL.n349 VTAIL.n348 585
R304 VTAIL.n324 VTAIL.n323 585
R305 VTAIL.n343 VTAIL.n342 585
R306 VTAIL.n341 VTAIL.n340 585
R307 VTAIL.n328 VTAIL.n327 585
R308 VTAIL.n335 VTAIL.n334 585
R309 VTAIL.n333 VTAIL.n332 585
R310 VTAIL.n725 VTAIL.t14 327.466
R311 VTAIL.n33 VTAIL.t9 327.466
R312 VTAIL.n131 VTAIL.t0 327.466
R313 VTAIL.n231 VTAIL.t1 327.466
R314 VTAIL.n629 VTAIL.t7 327.466
R315 VTAIL.n529 VTAIL.t3 327.466
R316 VTAIL.n431 VTAIL.t8 327.466
R317 VTAIL.n331 VTAIL.t13 327.466
R318 VTAIL.n728 VTAIL.n727 171.744
R319 VTAIL.n728 VTAIL.n721 171.744
R320 VTAIL.n735 VTAIL.n721 171.744
R321 VTAIL.n736 VTAIL.n735 171.744
R322 VTAIL.n736 VTAIL.n717 171.744
R323 VTAIL.n743 VTAIL.n717 171.744
R324 VTAIL.n744 VTAIL.n743 171.744
R325 VTAIL.n744 VTAIL.n713 171.744
R326 VTAIL.n751 VTAIL.n713 171.744
R327 VTAIL.n752 VTAIL.n751 171.744
R328 VTAIL.n752 VTAIL.n709 171.744
R329 VTAIL.n759 VTAIL.n709 171.744
R330 VTAIL.n760 VTAIL.n759 171.744
R331 VTAIL.n760 VTAIL.n705 171.744
R332 VTAIL.n768 VTAIL.n705 171.744
R333 VTAIL.n769 VTAIL.n768 171.744
R334 VTAIL.n770 VTAIL.n769 171.744
R335 VTAIL.n770 VTAIL.n701 171.744
R336 VTAIL.n777 VTAIL.n701 171.744
R337 VTAIL.n778 VTAIL.n777 171.744
R338 VTAIL.n778 VTAIL.n697 171.744
R339 VTAIL.n785 VTAIL.n697 171.744
R340 VTAIL.n786 VTAIL.n785 171.744
R341 VTAIL.n36 VTAIL.n35 171.744
R342 VTAIL.n36 VTAIL.n29 171.744
R343 VTAIL.n43 VTAIL.n29 171.744
R344 VTAIL.n44 VTAIL.n43 171.744
R345 VTAIL.n44 VTAIL.n25 171.744
R346 VTAIL.n51 VTAIL.n25 171.744
R347 VTAIL.n52 VTAIL.n51 171.744
R348 VTAIL.n52 VTAIL.n21 171.744
R349 VTAIL.n59 VTAIL.n21 171.744
R350 VTAIL.n60 VTAIL.n59 171.744
R351 VTAIL.n60 VTAIL.n17 171.744
R352 VTAIL.n67 VTAIL.n17 171.744
R353 VTAIL.n68 VTAIL.n67 171.744
R354 VTAIL.n68 VTAIL.n13 171.744
R355 VTAIL.n76 VTAIL.n13 171.744
R356 VTAIL.n77 VTAIL.n76 171.744
R357 VTAIL.n78 VTAIL.n77 171.744
R358 VTAIL.n78 VTAIL.n9 171.744
R359 VTAIL.n85 VTAIL.n9 171.744
R360 VTAIL.n86 VTAIL.n85 171.744
R361 VTAIL.n86 VTAIL.n5 171.744
R362 VTAIL.n93 VTAIL.n5 171.744
R363 VTAIL.n94 VTAIL.n93 171.744
R364 VTAIL.n134 VTAIL.n133 171.744
R365 VTAIL.n134 VTAIL.n127 171.744
R366 VTAIL.n141 VTAIL.n127 171.744
R367 VTAIL.n142 VTAIL.n141 171.744
R368 VTAIL.n142 VTAIL.n123 171.744
R369 VTAIL.n149 VTAIL.n123 171.744
R370 VTAIL.n150 VTAIL.n149 171.744
R371 VTAIL.n150 VTAIL.n119 171.744
R372 VTAIL.n157 VTAIL.n119 171.744
R373 VTAIL.n158 VTAIL.n157 171.744
R374 VTAIL.n158 VTAIL.n115 171.744
R375 VTAIL.n165 VTAIL.n115 171.744
R376 VTAIL.n166 VTAIL.n165 171.744
R377 VTAIL.n166 VTAIL.n111 171.744
R378 VTAIL.n174 VTAIL.n111 171.744
R379 VTAIL.n175 VTAIL.n174 171.744
R380 VTAIL.n176 VTAIL.n175 171.744
R381 VTAIL.n176 VTAIL.n107 171.744
R382 VTAIL.n183 VTAIL.n107 171.744
R383 VTAIL.n184 VTAIL.n183 171.744
R384 VTAIL.n184 VTAIL.n103 171.744
R385 VTAIL.n191 VTAIL.n103 171.744
R386 VTAIL.n192 VTAIL.n191 171.744
R387 VTAIL.n234 VTAIL.n233 171.744
R388 VTAIL.n234 VTAIL.n227 171.744
R389 VTAIL.n241 VTAIL.n227 171.744
R390 VTAIL.n242 VTAIL.n241 171.744
R391 VTAIL.n242 VTAIL.n223 171.744
R392 VTAIL.n249 VTAIL.n223 171.744
R393 VTAIL.n250 VTAIL.n249 171.744
R394 VTAIL.n250 VTAIL.n219 171.744
R395 VTAIL.n257 VTAIL.n219 171.744
R396 VTAIL.n258 VTAIL.n257 171.744
R397 VTAIL.n258 VTAIL.n215 171.744
R398 VTAIL.n265 VTAIL.n215 171.744
R399 VTAIL.n266 VTAIL.n265 171.744
R400 VTAIL.n266 VTAIL.n211 171.744
R401 VTAIL.n274 VTAIL.n211 171.744
R402 VTAIL.n275 VTAIL.n274 171.744
R403 VTAIL.n276 VTAIL.n275 171.744
R404 VTAIL.n276 VTAIL.n207 171.744
R405 VTAIL.n283 VTAIL.n207 171.744
R406 VTAIL.n284 VTAIL.n283 171.744
R407 VTAIL.n284 VTAIL.n203 171.744
R408 VTAIL.n291 VTAIL.n203 171.744
R409 VTAIL.n292 VTAIL.n291 171.744
R410 VTAIL.n688 VTAIL.n687 171.744
R411 VTAIL.n687 VTAIL.n599 171.744
R412 VTAIL.n680 VTAIL.n599 171.744
R413 VTAIL.n680 VTAIL.n679 171.744
R414 VTAIL.n679 VTAIL.n603 171.744
R415 VTAIL.n608 VTAIL.n603 171.744
R416 VTAIL.n672 VTAIL.n608 171.744
R417 VTAIL.n672 VTAIL.n671 171.744
R418 VTAIL.n671 VTAIL.n609 171.744
R419 VTAIL.n664 VTAIL.n609 171.744
R420 VTAIL.n664 VTAIL.n663 171.744
R421 VTAIL.n663 VTAIL.n613 171.744
R422 VTAIL.n656 VTAIL.n613 171.744
R423 VTAIL.n656 VTAIL.n655 171.744
R424 VTAIL.n655 VTAIL.n617 171.744
R425 VTAIL.n648 VTAIL.n617 171.744
R426 VTAIL.n648 VTAIL.n647 171.744
R427 VTAIL.n647 VTAIL.n621 171.744
R428 VTAIL.n640 VTAIL.n621 171.744
R429 VTAIL.n640 VTAIL.n639 171.744
R430 VTAIL.n639 VTAIL.n625 171.744
R431 VTAIL.n632 VTAIL.n625 171.744
R432 VTAIL.n632 VTAIL.n631 171.744
R433 VTAIL.n588 VTAIL.n587 171.744
R434 VTAIL.n587 VTAIL.n499 171.744
R435 VTAIL.n580 VTAIL.n499 171.744
R436 VTAIL.n580 VTAIL.n579 171.744
R437 VTAIL.n579 VTAIL.n503 171.744
R438 VTAIL.n508 VTAIL.n503 171.744
R439 VTAIL.n572 VTAIL.n508 171.744
R440 VTAIL.n572 VTAIL.n571 171.744
R441 VTAIL.n571 VTAIL.n509 171.744
R442 VTAIL.n564 VTAIL.n509 171.744
R443 VTAIL.n564 VTAIL.n563 171.744
R444 VTAIL.n563 VTAIL.n513 171.744
R445 VTAIL.n556 VTAIL.n513 171.744
R446 VTAIL.n556 VTAIL.n555 171.744
R447 VTAIL.n555 VTAIL.n517 171.744
R448 VTAIL.n548 VTAIL.n517 171.744
R449 VTAIL.n548 VTAIL.n547 171.744
R450 VTAIL.n547 VTAIL.n521 171.744
R451 VTAIL.n540 VTAIL.n521 171.744
R452 VTAIL.n540 VTAIL.n539 171.744
R453 VTAIL.n539 VTAIL.n525 171.744
R454 VTAIL.n532 VTAIL.n525 171.744
R455 VTAIL.n532 VTAIL.n531 171.744
R456 VTAIL.n490 VTAIL.n489 171.744
R457 VTAIL.n489 VTAIL.n401 171.744
R458 VTAIL.n482 VTAIL.n401 171.744
R459 VTAIL.n482 VTAIL.n481 171.744
R460 VTAIL.n481 VTAIL.n405 171.744
R461 VTAIL.n410 VTAIL.n405 171.744
R462 VTAIL.n474 VTAIL.n410 171.744
R463 VTAIL.n474 VTAIL.n473 171.744
R464 VTAIL.n473 VTAIL.n411 171.744
R465 VTAIL.n466 VTAIL.n411 171.744
R466 VTAIL.n466 VTAIL.n465 171.744
R467 VTAIL.n465 VTAIL.n415 171.744
R468 VTAIL.n458 VTAIL.n415 171.744
R469 VTAIL.n458 VTAIL.n457 171.744
R470 VTAIL.n457 VTAIL.n419 171.744
R471 VTAIL.n450 VTAIL.n419 171.744
R472 VTAIL.n450 VTAIL.n449 171.744
R473 VTAIL.n449 VTAIL.n423 171.744
R474 VTAIL.n442 VTAIL.n423 171.744
R475 VTAIL.n442 VTAIL.n441 171.744
R476 VTAIL.n441 VTAIL.n427 171.744
R477 VTAIL.n434 VTAIL.n427 171.744
R478 VTAIL.n434 VTAIL.n433 171.744
R479 VTAIL.n390 VTAIL.n389 171.744
R480 VTAIL.n389 VTAIL.n301 171.744
R481 VTAIL.n382 VTAIL.n301 171.744
R482 VTAIL.n382 VTAIL.n381 171.744
R483 VTAIL.n381 VTAIL.n305 171.744
R484 VTAIL.n310 VTAIL.n305 171.744
R485 VTAIL.n374 VTAIL.n310 171.744
R486 VTAIL.n374 VTAIL.n373 171.744
R487 VTAIL.n373 VTAIL.n311 171.744
R488 VTAIL.n366 VTAIL.n311 171.744
R489 VTAIL.n366 VTAIL.n365 171.744
R490 VTAIL.n365 VTAIL.n315 171.744
R491 VTAIL.n358 VTAIL.n315 171.744
R492 VTAIL.n358 VTAIL.n357 171.744
R493 VTAIL.n357 VTAIL.n319 171.744
R494 VTAIL.n350 VTAIL.n319 171.744
R495 VTAIL.n350 VTAIL.n349 171.744
R496 VTAIL.n349 VTAIL.n323 171.744
R497 VTAIL.n342 VTAIL.n323 171.744
R498 VTAIL.n342 VTAIL.n341 171.744
R499 VTAIL.n341 VTAIL.n327 171.744
R500 VTAIL.n334 VTAIL.n327 171.744
R501 VTAIL.n334 VTAIL.n333 171.744
R502 VTAIL.n727 VTAIL.t14 85.8723
R503 VTAIL.n35 VTAIL.t9 85.8723
R504 VTAIL.n133 VTAIL.t0 85.8723
R505 VTAIL.n233 VTAIL.t1 85.8723
R506 VTAIL.n631 VTAIL.t7 85.8723
R507 VTAIL.n531 VTAIL.t3 85.8723
R508 VTAIL.n433 VTAIL.t8 85.8723
R509 VTAIL.n333 VTAIL.t13 85.8723
R510 VTAIL.n595 VTAIL.n594 54.6707
R511 VTAIL.n397 VTAIL.n396 54.6707
R512 VTAIL.n1 VTAIL.n0 54.6705
R513 VTAIL.n199 VTAIL.n198 54.6705
R514 VTAIL.n791 VTAIL.n790 34.5126
R515 VTAIL.n99 VTAIL.n98 34.5126
R516 VTAIL.n197 VTAIL.n196 34.5126
R517 VTAIL.n297 VTAIL.n296 34.5126
R518 VTAIL.n693 VTAIL.n692 34.5126
R519 VTAIL.n593 VTAIL.n592 34.5126
R520 VTAIL.n495 VTAIL.n494 34.5126
R521 VTAIL.n395 VTAIL.n394 34.5126
R522 VTAIL.n791 VTAIL.n693 30.8841
R523 VTAIL.n395 VTAIL.n297 30.8841
R524 VTAIL.n726 VTAIL.n725 16.3895
R525 VTAIL.n34 VTAIL.n33 16.3895
R526 VTAIL.n132 VTAIL.n131 16.3895
R527 VTAIL.n232 VTAIL.n231 16.3895
R528 VTAIL.n630 VTAIL.n629 16.3895
R529 VTAIL.n530 VTAIL.n529 16.3895
R530 VTAIL.n432 VTAIL.n431 16.3895
R531 VTAIL.n332 VTAIL.n331 16.3895
R532 VTAIL.n771 VTAIL.n702 13.1884
R533 VTAIL.n79 VTAIL.n10 13.1884
R534 VTAIL.n177 VTAIL.n108 13.1884
R535 VTAIL.n277 VTAIL.n208 13.1884
R536 VTAIL.n606 VTAIL.n604 13.1884
R537 VTAIL.n506 VTAIL.n504 13.1884
R538 VTAIL.n408 VTAIL.n406 13.1884
R539 VTAIL.n308 VTAIL.n306 13.1884
R540 VTAIL.n729 VTAIL.n724 12.8005
R541 VTAIL.n772 VTAIL.n704 12.8005
R542 VTAIL.n776 VTAIL.n775 12.8005
R543 VTAIL.n37 VTAIL.n32 12.8005
R544 VTAIL.n80 VTAIL.n12 12.8005
R545 VTAIL.n84 VTAIL.n83 12.8005
R546 VTAIL.n135 VTAIL.n130 12.8005
R547 VTAIL.n178 VTAIL.n110 12.8005
R548 VTAIL.n182 VTAIL.n181 12.8005
R549 VTAIL.n235 VTAIL.n230 12.8005
R550 VTAIL.n278 VTAIL.n210 12.8005
R551 VTAIL.n282 VTAIL.n281 12.8005
R552 VTAIL.n678 VTAIL.n677 12.8005
R553 VTAIL.n674 VTAIL.n673 12.8005
R554 VTAIL.n633 VTAIL.n628 12.8005
R555 VTAIL.n578 VTAIL.n577 12.8005
R556 VTAIL.n574 VTAIL.n573 12.8005
R557 VTAIL.n533 VTAIL.n528 12.8005
R558 VTAIL.n480 VTAIL.n479 12.8005
R559 VTAIL.n476 VTAIL.n475 12.8005
R560 VTAIL.n435 VTAIL.n430 12.8005
R561 VTAIL.n380 VTAIL.n379 12.8005
R562 VTAIL.n376 VTAIL.n375 12.8005
R563 VTAIL.n335 VTAIL.n330 12.8005
R564 VTAIL.n730 VTAIL.n722 12.0247
R565 VTAIL.n767 VTAIL.n766 12.0247
R566 VTAIL.n779 VTAIL.n700 12.0247
R567 VTAIL.n38 VTAIL.n30 12.0247
R568 VTAIL.n75 VTAIL.n74 12.0247
R569 VTAIL.n87 VTAIL.n8 12.0247
R570 VTAIL.n136 VTAIL.n128 12.0247
R571 VTAIL.n173 VTAIL.n172 12.0247
R572 VTAIL.n185 VTAIL.n106 12.0247
R573 VTAIL.n236 VTAIL.n228 12.0247
R574 VTAIL.n273 VTAIL.n272 12.0247
R575 VTAIL.n285 VTAIL.n206 12.0247
R576 VTAIL.n681 VTAIL.n602 12.0247
R577 VTAIL.n670 VTAIL.n607 12.0247
R578 VTAIL.n634 VTAIL.n626 12.0247
R579 VTAIL.n581 VTAIL.n502 12.0247
R580 VTAIL.n570 VTAIL.n507 12.0247
R581 VTAIL.n534 VTAIL.n526 12.0247
R582 VTAIL.n483 VTAIL.n404 12.0247
R583 VTAIL.n472 VTAIL.n409 12.0247
R584 VTAIL.n436 VTAIL.n428 12.0247
R585 VTAIL.n383 VTAIL.n304 12.0247
R586 VTAIL.n372 VTAIL.n309 12.0247
R587 VTAIL.n336 VTAIL.n328 12.0247
R588 VTAIL.n734 VTAIL.n733 11.249
R589 VTAIL.n765 VTAIL.n706 11.249
R590 VTAIL.n780 VTAIL.n698 11.249
R591 VTAIL.n42 VTAIL.n41 11.249
R592 VTAIL.n73 VTAIL.n14 11.249
R593 VTAIL.n88 VTAIL.n6 11.249
R594 VTAIL.n140 VTAIL.n139 11.249
R595 VTAIL.n171 VTAIL.n112 11.249
R596 VTAIL.n186 VTAIL.n104 11.249
R597 VTAIL.n240 VTAIL.n239 11.249
R598 VTAIL.n271 VTAIL.n212 11.249
R599 VTAIL.n286 VTAIL.n204 11.249
R600 VTAIL.n682 VTAIL.n600 11.249
R601 VTAIL.n669 VTAIL.n610 11.249
R602 VTAIL.n638 VTAIL.n637 11.249
R603 VTAIL.n582 VTAIL.n500 11.249
R604 VTAIL.n569 VTAIL.n510 11.249
R605 VTAIL.n538 VTAIL.n537 11.249
R606 VTAIL.n484 VTAIL.n402 11.249
R607 VTAIL.n471 VTAIL.n412 11.249
R608 VTAIL.n440 VTAIL.n439 11.249
R609 VTAIL.n384 VTAIL.n302 11.249
R610 VTAIL.n371 VTAIL.n312 11.249
R611 VTAIL.n340 VTAIL.n339 11.249
R612 VTAIL.n737 VTAIL.n720 10.4732
R613 VTAIL.n762 VTAIL.n761 10.4732
R614 VTAIL.n784 VTAIL.n783 10.4732
R615 VTAIL.n45 VTAIL.n28 10.4732
R616 VTAIL.n70 VTAIL.n69 10.4732
R617 VTAIL.n92 VTAIL.n91 10.4732
R618 VTAIL.n143 VTAIL.n126 10.4732
R619 VTAIL.n168 VTAIL.n167 10.4732
R620 VTAIL.n190 VTAIL.n189 10.4732
R621 VTAIL.n243 VTAIL.n226 10.4732
R622 VTAIL.n268 VTAIL.n267 10.4732
R623 VTAIL.n290 VTAIL.n289 10.4732
R624 VTAIL.n686 VTAIL.n685 10.4732
R625 VTAIL.n666 VTAIL.n665 10.4732
R626 VTAIL.n641 VTAIL.n624 10.4732
R627 VTAIL.n586 VTAIL.n585 10.4732
R628 VTAIL.n566 VTAIL.n565 10.4732
R629 VTAIL.n541 VTAIL.n524 10.4732
R630 VTAIL.n488 VTAIL.n487 10.4732
R631 VTAIL.n468 VTAIL.n467 10.4732
R632 VTAIL.n443 VTAIL.n426 10.4732
R633 VTAIL.n388 VTAIL.n387 10.4732
R634 VTAIL.n368 VTAIL.n367 10.4732
R635 VTAIL.n343 VTAIL.n326 10.4732
R636 VTAIL.n738 VTAIL.n718 9.69747
R637 VTAIL.n758 VTAIL.n708 9.69747
R638 VTAIL.n787 VTAIL.n696 9.69747
R639 VTAIL.n46 VTAIL.n26 9.69747
R640 VTAIL.n66 VTAIL.n16 9.69747
R641 VTAIL.n95 VTAIL.n4 9.69747
R642 VTAIL.n144 VTAIL.n124 9.69747
R643 VTAIL.n164 VTAIL.n114 9.69747
R644 VTAIL.n193 VTAIL.n102 9.69747
R645 VTAIL.n244 VTAIL.n224 9.69747
R646 VTAIL.n264 VTAIL.n214 9.69747
R647 VTAIL.n293 VTAIL.n202 9.69747
R648 VTAIL.n689 VTAIL.n598 9.69747
R649 VTAIL.n662 VTAIL.n612 9.69747
R650 VTAIL.n642 VTAIL.n622 9.69747
R651 VTAIL.n589 VTAIL.n498 9.69747
R652 VTAIL.n562 VTAIL.n512 9.69747
R653 VTAIL.n542 VTAIL.n522 9.69747
R654 VTAIL.n491 VTAIL.n400 9.69747
R655 VTAIL.n464 VTAIL.n414 9.69747
R656 VTAIL.n444 VTAIL.n424 9.69747
R657 VTAIL.n391 VTAIL.n300 9.69747
R658 VTAIL.n364 VTAIL.n314 9.69747
R659 VTAIL.n344 VTAIL.n324 9.69747
R660 VTAIL.n790 VTAIL.n789 9.45567
R661 VTAIL.n98 VTAIL.n97 9.45567
R662 VTAIL.n196 VTAIL.n195 9.45567
R663 VTAIL.n296 VTAIL.n295 9.45567
R664 VTAIL.n692 VTAIL.n691 9.45567
R665 VTAIL.n592 VTAIL.n591 9.45567
R666 VTAIL.n494 VTAIL.n493 9.45567
R667 VTAIL.n394 VTAIL.n393 9.45567
R668 VTAIL.n789 VTAIL.n788 9.3005
R669 VTAIL.n696 VTAIL.n695 9.3005
R670 VTAIL.n783 VTAIL.n782 9.3005
R671 VTAIL.n781 VTAIL.n780 9.3005
R672 VTAIL.n700 VTAIL.n699 9.3005
R673 VTAIL.n775 VTAIL.n774 9.3005
R674 VTAIL.n747 VTAIL.n746 9.3005
R675 VTAIL.n716 VTAIL.n715 9.3005
R676 VTAIL.n741 VTAIL.n740 9.3005
R677 VTAIL.n739 VTAIL.n738 9.3005
R678 VTAIL.n720 VTAIL.n719 9.3005
R679 VTAIL.n733 VTAIL.n732 9.3005
R680 VTAIL.n731 VTAIL.n730 9.3005
R681 VTAIL.n724 VTAIL.n723 9.3005
R682 VTAIL.n749 VTAIL.n748 9.3005
R683 VTAIL.n712 VTAIL.n711 9.3005
R684 VTAIL.n755 VTAIL.n754 9.3005
R685 VTAIL.n757 VTAIL.n756 9.3005
R686 VTAIL.n708 VTAIL.n707 9.3005
R687 VTAIL.n763 VTAIL.n762 9.3005
R688 VTAIL.n765 VTAIL.n764 9.3005
R689 VTAIL.n766 VTAIL.n703 9.3005
R690 VTAIL.n773 VTAIL.n772 9.3005
R691 VTAIL.n97 VTAIL.n96 9.3005
R692 VTAIL.n4 VTAIL.n3 9.3005
R693 VTAIL.n91 VTAIL.n90 9.3005
R694 VTAIL.n89 VTAIL.n88 9.3005
R695 VTAIL.n8 VTAIL.n7 9.3005
R696 VTAIL.n83 VTAIL.n82 9.3005
R697 VTAIL.n55 VTAIL.n54 9.3005
R698 VTAIL.n24 VTAIL.n23 9.3005
R699 VTAIL.n49 VTAIL.n48 9.3005
R700 VTAIL.n47 VTAIL.n46 9.3005
R701 VTAIL.n28 VTAIL.n27 9.3005
R702 VTAIL.n41 VTAIL.n40 9.3005
R703 VTAIL.n39 VTAIL.n38 9.3005
R704 VTAIL.n32 VTAIL.n31 9.3005
R705 VTAIL.n57 VTAIL.n56 9.3005
R706 VTAIL.n20 VTAIL.n19 9.3005
R707 VTAIL.n63 VTAIL.n62 9.3005
R708 VTAIL.n65 VTAIL.n64 9.3005
R709 VTAIL.n16 VTAIL.n15 9.3005
R710 VTAIL.n71 VTAIL.n70 9.3005
R711 VTAIL.n73 VTAIL.n72 9.3005
R712 VTAIL.n74 VTAIL.n11 9.3005
R713 VTAIL.n81 VTAIL.n80 9.3005
R714 VTAIL.n195 VTAIL.n194 9.3005
R715 VTAIL.n102 VTAIL.n101 9.3005
R716 VTAIL.n189 VTAIL.n188 9.3005
R717 VTAIL.n187 VTAIL.n186 9.3005
R718 VTAIL.n106 VTAIL.n105 9.3005
R719 VTAIL.n181 VTAIL.n180 9.3005
R720 VTAIL.n153 VTAIL.n152 9.3005
R721 VTAIL.n122 VTAIL.n121 9.3005
R722 VTAIL.n147 VTAIL.n146 9.3005
R723 VTAIL.n145 VTAIL.n144 9.3005
R724 VTAIL.n126 VTAIL.n125 9.3005
R725 VTAIL.n139 VTAIL.n138 9.3005
R726 VTAIL.n137 VTAIL.n136 9.3005
R727 VTAIL.n130 VTAIL.n129 9.3005
R728 VTAIL.n155 VTAIL.n154 9.3005
R729 VTAIL.n118 VTAIL.n117 9.3005
R730 VTAIL.n161 VTAIL.n160 9.3005
R731 VTAIL.n163 VTAIL.n162 9.3005
R732 VTAIL.n114 VTAIL.n113 9.3005
R733 VTAIL.n169 VTAIL.n168 9.3005
R734 VTAIL.n171 VTAIL.n170 9.3005
R735 VTAIL.n172 VTAIL.n109 9.3005
R736 VTAIL.n179 VTAIL.n178 9.3005
R737 VTAIL.n295 VTAIL.n294 9.3005
R738 VTAIL.n202 VTAIL.n201 9.3005
R739 VTAIL.n289 VTAIL.n288 9.3005
R740 VTAIL.n287 VTAIL.n286 9.3005
R741 VTAIL.n206 VTAIL.n205 9.3005
R742 VTAIL.n281 VTAIL.n280 9.3005
R743 VTAIL.n253 VTAIL.n252 9.3005
R744 VTAIL.n222 VTAIL.n221 9.3005
R745 VTAIL.n247 VTAIL.n246 9.3005
R746 VTAIL.n245 VTAIL.n244 9.3005
R747 VTAIL.n226 VTAIL.n225 9.3005
R748 VTAIL.n239 VTAIL.n238 9.3005
R749 VTAIL.n237 VTAIL.n236 9.3005
R750 VTAIL.n230 VTAIL.n229 9.3005
R751 VTAIL.n255 VTAIL.n254 9.3005
R752 VTAIL.n218 VTAIL.n217 9.3005
R753 VTAIL.n261 VTAIL.n260 9.3005
R754 VTAIL.n263 VTAIL.n262 9.3005
R755 VTAIL.n214 VTAIL.n213 9.3005
R756 VTAIL.n269 VTAIL.n268 9.3005
R757 VTAIL.n271 VTAIL.n270 9.3005
R758 VTAIL.n272 VTAIL.n209 9.3005
R759 VTAIL.n279 VTAIL.n278 9.3005
R760 VTAIL.n616 VTAIL.n615 9.3005
R761 VTAIL.n659 VTAIL.n658 9.3005
R762 VTAIL.n661 VTAIL.n660 9.3005
R763 VTAIL.n612 VTAIL.n611 9.3005
R764 VTAIL.n667 VTAIL.n666 9.3005
R765 VTAIL.n669 VTAIL.n668 9.3005
R766 VTAIL.n607 VTAIL.n605 9.3005
R767 VTAIL.n675 VTAIL.n674 9.3005
R768 VTAIL.n691 VTAIL.n690 9.3005
R769 VTAIL.n598 VTAIL.n597 9.3005
R770 VTAIL.n685 VTAIL.n684 9.3005
R771 VTAIL.n683 VTAIL.n682 9.3005
R772 VTAIL.n602 VTAIL.n601 9.3005
R773 VTAIL.n677 VTAIL.n676 9.3005
R774 VTAIL.n653 VTAIL.n652 9.3005
R775 VTAIL.n651 VTAIL.n650 9.3005
R776 VTAIL.n620 VTAIL.n619 9.3005
R777 VTAIL.n645 VTAIL.n644 9.3005
R778 VTAIL.n643 VTAIL.n642 9.3005
R779 VTAIL.n624 VTAIL.n623 9.3005
R780 VTAIL.n637 VTAIL.n636 9.3005
R781 VTAIL.n635 VTAIL.n634 9.3005
R782 VTAIL.n628 VTAIL.n627 9.3005
R783 VTAIL.n516 VTAIL.n515 9.3005
R784 VTAIL.n559 VTAIL.n558 9.3005
R785 VTAIL.n561 VTAIL.n560 9.3005
R786 VTAIL.n512 VTAIL.n511 9.3005
R787 VTAIL.n567 VTAIL.n566 9.3005
R788 VTAIL.n569 VTAIL.n568 9.3005
R789 VTAIL.n507 VTAIL.n505 9.3005
R790 VTAIL.n575 VTAIL.n574 9.3005
R791 VTAIL.n591 VTAIL.n590 9.3005
R792 VTAIL.n498 VTAIL.n497 9.3005
R793 VTAIL.n585 VTAIL.n584 9.3005
R794 VTAIL.n583 VTAIL.n582 9.3005
R795 VTAIL.n502 VTAIL.n501 9.3005
R796 VTAIL.n577 VTAIL.n576 9.3005
R797 VTAIL.n553 VTAIL.n552 9.3005
R798 VTAIL.n551 VTAIL.n550 9.3005
R799 VTAIL.n520 VTAIL.n519 9.3005
R800 VTAIL.n545 VTAIL.n544 9.3005
R801 VTAIL.n543 VTAIL.n542 9.3005
R802 VTAIL.n524 VTAIL.n523 9.3005
R803 VTAIL.n537 VTAIL.n536 9.3005
R804 VTAIL.n535 VTAIL.n534 9.3005
R805 VTAIL.n528 VTAIL.n527 9.3005
R806 VTAIL.n418 VTAIL.n417 9.3005
R807 VTAIL.n461 VTAIL.n460 9.3005
R808 VTAIL.n463 VTAIL.n462 9.3005
R809 VTAIL.n414 VTAIL.n413 9.3005
R810 VTAIL.n469 VTAIL.n468 9.3005
R811 VTAIL.n471 VTAIL.n470 9.3005
R812 VTAIL.n409 VTAIL.n407 9.3005
R813 VTAIL.n477 VTAIL.n476 9.3005
R814 VTAIL.n493 VTAIL.n492 9.3005
R815 VTAIL.n400 VTAIL.n399 9.3005
R816 VTAIL.n487 VTAIL.n486 9.3005
R817 VTAIL.n485 VTAIL.n484 9.3005
R818 VTAIL.n404 VTAIL.n403 9.3005
R819 VTAIL.n479 VTAIL.n478 9.3005
R820 VTAIL.n455 VTAIL.n454 9.3005
R821 VTAIL.n453 VTAIL.n452 9.3005
R822 VTAIL.n422 VTAIL.n421 9.3005
R823 VTAIL.n447 VTAIL.n446 9.3005
R824 VTAIL.n445 VTAIL.n444 9.3005
R825 VTAIL.n426 VTAIL.n425 9.3005
R826 VTAIL.n439 VTAIL.n438 9.3005
R827 VTAIL.n437 VTAIL.n436 9.3005
R828 VTAIL.n430 VTAIL.n429 9.3005
R829 VTAIL.n318 VTAIL.n317 9.3005
R830 VTAIL.n361 VTAIL.n360 9.3005
R831 VTAIL.n363 VTAIL.n362 9.3005
R832 VTAIL.n314 VTAIL.n313 9.3005
R833 VTAIL.n369 VTAIL.n368 9.3005
R834 VTAIL.n371 VTAIL.n370 9.3005
R835 VTAIL.n309 VTAIL.n307 9.3005
R836 VTAIL.n377 VTAIL.n376 9.3005
R837 VTAIL.n393 VTAIL.n392 9.3005
R838 VTAIL.n300 VTAIL.n299 9.3005
R839 VTAIL.n387 VTAIL.n386 9.3005
R840 VTAIL.n385 VTAIL.n384 9.3005
R841 VTAIL.n304 VTAIL.n303 9.3005
R842 VTAIL.n379 VTAIL.n378 9.3005
R843 VTAIL.n355 VTAIL.n354 9.3005
R844 VTAIL.n353 VTAIL.n352 9.3005
R845 VTAIL.n322 VTAIL.n321 9.3005
R846 VTAIL.n347 VTAIL.n346 9.3005
R847 VTAIL.n345 VTAIL.n344 9.3005
R848 VTAIL.n326 VTAIL.n325 9.3005
R849 VTAIL.n339 VTAIL.n338 9.3005
R850 VTAIL.n337 VTAIL.n336 9.3005
R851 VTAIL.n330 VTAIL.n329 9.3005
R852 VTAIL.n742 VTAIL.n741 8.92171
R853 VTAIL.n757 VTAIL.n710 8.92171
R854 VTAIL.n788 VTAIL.n694 8.92171
R855 VTAIL.n50 VTAIL.n49 8.92171
R856 VTAIL.n65 VTAIL.n18 8.92171
R857 VTAIL.n96 VTAIL.n2 8.92171
R858 VTAIL.n148 VTAIL.n147 8.92171
R859 VTAIL.n163 VTAIL.n116 8.92171
R860 VTAIL.n194 VTAIL.n100 8.92171
R861 VTAIL.n248 VTAIL.n247 8.92171
R862 VTAIL.n263 VTAIL.n216 8.92171
R863 VTAIL.n294 VTAIL.n200 8.92171
R864 VTAIL.n690 VTAIL.n596 8.92171
R865 VTAIL.n661 VTAIL.n614 8.92171
R866 VTAIL.n646 VTAIL.n645 8.92171
R867 VTAIL.n590 VTAIL.n496 8.92171
R868 VTAIL.n561 VTAIL.n514 8.92171
R869 VTAIL.n546 VTAIL.n545 8.92171
R870 VTAIL.n492 VTAIL.n398 8.92171
R871 VTAIL.n463 VTAIL.n416 8.92171
R872 VTAIL.n448 VTAIL.n447 8.92171
R873 VTAIL.n392 VTAIL.n298 8.92171
R874 VTAIL.n363 VTAIL.n316 8.92171
R875 VTAIL.n348 VTAIL.n347 8.92171
R876 VTAIL.n745 VTAIL.n716 8.14595
R877 VTAIL.n754 VTAIL.n753 8.14595
R878 VTAIL.n53 VTAIL.n24 8.14595
R879 VTAIL.n62 VTAIL.n61 8.14595
R880 VTAIL.n151 VTAIL.n122 8.14595
R881 VTAIL.n160 VTAIL.n159 8.14595
R882 VTAIL.n251 VTAIL.n222 8.14595
R883 VTAIL.n260 VTAIL.n259 8.14595
R884 VTAIL.n658 VTAIL.n657 8.14595
R885 VTAIL.n649 VTAIL.n620 8.14595
R886 VTAIL.n558 VTAIL.n557 8.14595
R887 VTAIL.n549 VTAIL.n520 8.14595
R888 VTAIL.n460 VTAIL.n459 8.14595
R889 VTAIL.n451 VTAIL.n422 8.14595
R890 VTAIL.n360 VTAIL.n359 8.14595
R891 VTAIL.n351 VTAIL.n322 8.14595
R892 VTAIL.n746 VTAIL.n714 7.3702
R893 VTAIL.n750 VTAIL.n712 7.3702
R894 VTAIL.n54 VTAIL.n22 7.3702
R895 VTAIL.n58 VTAIL.n20 7.3702
R896 VTAIL.n152 VTAIL.n120 7.3702
R897 VTAIL.n156 VTAIL.n118 7.3702
R898 VTAIL.n252 VTAIL.n220 7.3702
R899 VTAIL.n256 VTAIL.n218 7.3702
R900 VTAIL.n654 VTAIL.n616 7.3702
R901 VTAIL.n650 VTAIL.n618 7.3702
R902 VTAIL.n554 VTAIL.n516 7.3702
R903 VTAIL.n550 VTAIL.n518 7.3702
R904 VTAIL.n456 VTAIL.n418 7.3702
R905 VTAIL.n452 VTAIL.n420 7.3702
R906 VTAIL.n356 VTAIL.n318 7.3702
R907 VTAIL.n352 VTAIL.n320 7.3702
R908 VTAIL.n749 VTAIL.n714 6.59444
R909 VTAIL.n750 VTAIL.n749 6.59444
R910 VTAIL.n57 VTAIL.n22 6.59444
R911 VTAIL.n58 VTAIL.n57 6.59444
R912 VTAIL.n155 VTAIL.n120 6.59444
R913 VTAIL.n156 VTAIL.n155 6.59444
R914 VTAIL.n255 VTAIL.n220 6.59444
R915 VTAIL.n256 VTAIL.n255 6.59444
R916 VTAIL.n654 VTAIL.n653 6.59444
R917 VTAIL.n653 VTAIL.n618 6.59444
R918 VTAIL.n554 VTAIL.n553 6.59444
R919 VTAIL.n553 VTAIL.n518 6.59444
R920 VTAIL.n456 VTAIL.n455 6.59444
R921 VTAIL.n455 VTAIL.n420 6.59444
R922 VTAIL.n356 VTAIL.n355 6.59444
R923 VTAIL.n355 VTAIL.n320 6.59444
R924 VTAIL.n746 VTAIL.n745 5.81868
R925 VTAIL.n753 VTAIL.n712 5.81868
R926 VTAIL.n54 VTAIL.n53 5.81868
R927 VTAIL.n61 VTAIL.n20 5.81868
R928 VTAIL.n152 VTAIL.n151 5.81868
R929 VTAIL.n159 VTAIL.n118 5.81868
R930 VTAIL.n252 VTAIL.n251 5.81868
R931 VTAIL.n259 VTAIL.n218 5.81868
R932 VTAIL.n657 VTAIL.n616 5.81868
R933 VTAIL.n650 VTAIL.n649 5.81868
R934 VTAIL.n557 VTAIL.n516 5.81868
R935 VTAIL.n550 VTAIL.n549 5.81868
R936 VTAIL.n459 VTAIL.n418 5.81868
R937 VTAIL.n452 VTAIL.n451 5.81868
R938 VTAIL.n359 VTAIL.n318 5.81868
R939 VTAIL.n352 VTAIL.n351 5.81868
R940 VTAIL.n742 VTAIL.n716 5.04292
R941 VTAIL.n754 VTAIL.n710 5.04292
R942 VTAIL.n790 VTAIL.n694 5.04292
R943 VTAIL.n50 VTAIL.n24 5.04292
R944 VTAIL.n62 VTAIL.n18 5.04292
R945 VTAIL.n98 VTAIL.n2 5.04292
R946 VTAIL.n148 VTAIL.n122 5.04292
R947 VTAIL.n160 VTAIL.n116 5.04292
R948 VTAIL.n196 VTAIL.n100 5.04292
R949 VTAIL.n248 VTAIL.n222 5.04292
R950 VTAIL.n260 VTAIL.n216 5.04292
R951 VTAIL.n296 VTAIL.n200 5.04292
R952 VTAIL.n692 VTAIL.n596 5.04292
R953 VTAIL.n658 VTAIL.n614 5.04292
R954 VTAIL.n646 VTAIL.n620 5.04292
R955 VTAIL.n592 VTAIL.n496 5.04292
R956 VTAIL.n558 VTAIL.n514 5.04292
R957 VTAIL.n546 VTAIL.n520 5.04292
R958 VTAIL.n494 VTAIL.n398 5.04292
R959 VTAIL.n460 VTAIL.n416 5.04292
R960 VTAIL.n448 VTAIL.n422 5.04292
R961 VTAIL.n394 VTAIL.n298 5.04292
R962 VTAIL.n360 VTAIL.n316 5.04292
R963 VTAIL.n348 VTAIL.n322 5.04292
R964 VTAIL.n741 VTAIL.n718 4.26717
R965 VTAIL.n758 VTAIL.n757 4.26717
R966 VTAIL.n788 VTAIL.n787 4.26717
R967 VTAIL.n49 VTAIL.n26 4.26717
R968 VTAIL.n66 VTAIL.n65 4.26717
R969 VTAIL.n96 VTAIL.n95 4.26717
R970 VTAIL.n147 VTAIL.n124 4.26717
R971 VTAIL.n164 VTAIL.n163 4.26717
R972 VTAIL.n194 VTAIL.n193 4.26717
R973 VTAIL.n247 VTAIL.n224 4.26717
R974 VTAIL.n264 VTAIL.n263 4.26717
R975 VTAIL.n294 VTAIL.n293 4.26717
R976 VTAIL.n690 VTAIL.n689 4.26717
R977 VTAIL.n662 VTAIL.n661 4.26717
R978 VTAIL.n645 VTAIL.n622 4.26717
R979 VTAIL.n590 VTAIL.n589 4.26717
R980 VTAIL.n562 VTAIL.n561 4.26717
R981 VTAIL.n545 VTAIL.n522 4.26717
R982 VTAIL.n492 VTAIL.n491 4.26717
R983 VTAIL.n464 VTAIL.n463 4.26717
R984 VTAIL.n447 VTAIL.n424 4.26717
R985 VTAIL.n392 VTAIL.n391 4.26717
R986 VTAIL.n364 VTAIL.n363 4.26717
R987 VTAIL.n347 VTAIL.n324 4.26717
R988 VTAIL.n725 VTAIL.n723 3.70982
R989 VTAIL.n33 VTAIL.n31 3.70982
R990 VTAIL.n131 VTAIL.n129 3.70982
R991 VTAIL.n231 VTAIL.n229 3.70982
R992 VTAIL.n629 VTAIL.n627 3.70982
R993 VTAIL.n529 VTAIL.n527 3.70982
R994 VTAIL.n431 VTAIL.n429 3.70982
R995 VTAIL.n331 VTAIL.n329 3.70982
R996 VTAIL.n738 VTAIL.n737 3.49141
R997 VTAIL.n761 VTAIL.n708 3.49141
R998 VTAIL.n784 VTAIL.n696 3.49141
R999 VTAIL.n46 VTAIL.n45 3.49141
R1000 VTAIL.n69 VTAIL.n16 3.49141
R1001 VTAIL.n92 VTAIL.n4 3.49141
R1002 VTAIL.n144 VTAIL.n143 3.49141
R1003 VTAIL.n167 VTAIL.n114 3.49141
R1004 VTAIL.n190 VTAIL.n102 3.49141
R1005 VTAIL.n244 VTAIL.n243 3.49141
R1006 VTAIL.n267 VTAIL.n214 3.49141
R1007 VTAIL.n290 VTAIL.n202 3.49141
R1008 VTAIL.n686 VTAIL.n598 3.49141
R1009 VTAIL.n665 VTAIL.n612 3.49141
R1010 VTAIL.n642 VTAIL.n641 3.49141
R1011 VTAIL.n586 VTAIL.n498 3.49141
R1012 VTAIL.n565 VTAIL.n512 3.49141
R1013 VTAIL.n542 VTAIL.n541 3.49141
R1014 VTAIL.n488 VTAIL.n400 3.49141
R1015 VTAIL.n467 VTAIL.n414 3.49141
R1016 VTAIL.n444 VTAIL.n443 3.49141
R1017 VTAIL.n388 VTAIL.n300 3.49141
R1018 VTAIL.n367 VTAIL.n314 3.49141
R1019 VTAIL.n344 VTAIL.n343 3.49141
R1020 VTAIL.n397 VTAIL.n395 3.31084
R1021 VTAIL.n495 VTAIL.n397 3.31084
R1022 VTAIL.n595 VTAIL.n593 3.31084
R1023 VTAIL.n693 VTAIL.n595 3.31084
R1024 VTAIL.n297 VTAIL.n199 3.31084
R1025 VTAIL.n199 VTAIL.n197 3.31084
R1026 VTAIL.n99 VTAIL.n1 3.31084
R1027 VTAIL VTAIL.n791 3.25266
R1028 VTAIL.n734 VTAIL.n720 2.71565
R1029 VTAIL.n762 VTAIL.n706 2.71565
R1030 VTAIL.n783 VTAIL.n698 2.71565
R1031 VTAIL.n42 VTAIL.n28 2.71565
R1032 VTAIL.n70 VTAIL.n14 2.71565
R1033 VTAIL.n91 VTAIL.n6 2.71565
R1034 VTAIL.n140 VTAIL.n126 2.71565
R1035 VTAIL.n168 VTAIL.n112 2.71565
R1036 VTAIL.n189 VTAIL.n104 2.71565
R1037 VTAIL.n240 VTAIL.n226 2.71565
R1038 VTAIL.n268 VTAIL.n212 2.71565
R1039 VTAIL.n289 VTAIL.n204 2.71565
R1040 VTAIL.n685 VTAIL.n600 2.71565
R1041 VTAIL.n666 VTAIL.n610 2.71565
R1042 VTAIL.n638 VTAIL.n624 2.71565
R1043 VTAIL.n585 VTAIL.n500 2.71565
R1044 VTAIL.n566 VTAIL.n510 2.71565
R1045 VTAIL.n538 VTAIL.n524 2.71565
R1046 VTAIL.n487 VTAIL.n402 2.71565
R1047 VTAIL.n468 VTAIL.n412 2.71565
R1048 VTAIL.n440 VTAIL.n426 2.71565
R1049 VTAIL.n387 VTAIL.n302 2.71565
R1050 VTAIL.n368 VTAIL.n312 2.71565
R1051 VTAIL.n340 VTAIL.n326 2.71565
R1052 VTAIL.n733 VTAIL.n722 1.93989
R1053 VTAIL.n767 VTAIL.n765 1.93989
R1054 VTAIL.n780 VTAIL.n779 1.93989
R1055 VTAIL.n41 VTAIL.n30 1.93989
R1056 VTAIL.n75 VTAIL.n73 1.93989
R1057 VTAIL.n88 VTAIL.n87 1.93989
R1058 VTAIL.n139 VTAIL.n128 1.93989
R1059 VTAIL.n173 VTAIL.n171 1.93989
R1060 VTAIL.n186 VTAIL.n185 1.93989
R1061 VTAIL.n239 VTAIL.n228 1.93989
R1062 VTAIL.n273 VTAIL.n271 1.93989
R1063 VTAIL.n286 VTAIL.n285 1.93989
R1064 VTAIL.n682 VTAIL.n681 1.93989
R1065 VTAIL.n670 VTAIL.n669 1.93989
R1066 VTAIL.n637 VTAIL.n626 1.93989
R1067 VTAIL.n582 VTAIL.n581 1.93989
R1068 VTAIL.n570 VTAIL.n569 1.93989
R1069 VTAIL.n537 VTAIL.n526 1.93989
R1070 VTAIL.n484 VTAIL.n483 1.93989
R1071 VTAIL.n472 VTAIL.n471 1.93989
R1072 VTAIL.n439 VTAIL.n428 1.93989
R1073 VTAIL.n384 VTAIL.n383 1.93989
R1074 VTAIL.n372 VTAIL.n371 1.93989
R1075 VTAIL.n339 VTAIL.n328 1.93989
R1076 VTAIL.n0 VTAIL.t10 1.84319
R1077 VTAIL.n0 VTAIL.t12 1.84319
R1078 VTAIL.n198 VTAIL.t5 1.84319
R1079 VTAIL.n198 VTAIL.t6 1.84319
R1080 VTAIL.n594 VTAIL.t4 1.84319
R1081 VTAIL.n594 VTAIL.t2 1.84319
R1082 VTAIL.n396 VTAIL.t11 1.84319
R1083 VTAIL.n396 VTAIL.t15 1.84319
R1084 VTAIL.n730 VTAIL.n729 1.16414
R1085 VTAIL.n766 VTAIL.n704 1.16414
R1086 VTAIL.n776 VTAIL.n700 1.16414
R1087 VTAIL.n38 VTAIL.n37 1.16414
R1088 VTAIL.n74 VTAIL.n12 1.16414
R1089 VTAIL.n84 VTAIL.n8 1.16414
R1090 VTAIL.n136 VTAIL.n135 1.16414
R1091 VTAIL.n172 VTAIL.n110 1.16414
R1092 VTAIL.n182 VTAIL.n106 1.16414
R1093 VTAIL.n236 VTAIL.n235 1.16414
R1094 VTAIL.n272 VTAIL.n210 1.16414
R1095 VTAIL.n282 VTAIL.n206 1.16414
R1096 VTAIL.n678 VTAIL.n602 1.16414
R1097 VTAIL.n673 VTAIL.n607 1.16414
R1098 VTAIL.n634 VTAIL.n633 1.16414
R1099 VTAIL.n578 VTAIL.n502 1.16414
R1100 VTAIL.n573 VTAIL.n507 1.16414
R1101 VTAIL.n534 VTAIL.n533 1.16414
R1102 VTAIL.n480 VTAIL.n404 1.16414
R1103 VTAIL.n475 VTAIL.n409 1.16414
R1104 VTAIL.n436 VTAIL.n435 1.16414
R1105 VTAIL.n380 VTAIL.n304 1.16414
R1106 VTAIL.n375 VTAIL.n309 1.16414
R1107 VTAIL.n336 VTAIL.n335 1.16414
R1108 VTAIL.n593 VTAIL.n495 0.470328
R1109 VTAIL.n197 VTAIL.n99 0.470328
R1110 VTAIL.n726 VTAIL.n724 0.388379
R1111 VTAIL.n772 VTAIL.n771 0.388379
R1112 VTAIL.n775 VTAIL.n702 0.388379
R1113 VTAIL.n34 VTAIL.n32 0.388379
R1114 VTAIL.n80 VTAIL.n79 0.388379
R1115 VTAIL.n83 VTAIL.n10 0.388379
R1116 VTAIL.n132 VTAIL.n130 0.388379
R1117 VTAIL.n178 VTAIL.n177 0.388379
R1118 VTAIL.n181 VTAIL.n108 0.388379
R1119 VTAIL.n232 VTAIL.n230 0.388379
R1120 VTAIL.n278 VTAIL.n277 0.388379
R1121 VTAIL.n281 VTAIL.n208 0.388379
R1122 VTAIL.n677 VTAIL.n604 0.388379
R1123 VTAIL.n674 VTAIL.n606 0.388379
R1124 VTAIL.n630 VTAIL.n628 0.388379
R1125 VTAIL.n577 VTAIL.n504 0.388379
R1126 VTAIL.n574 VTAIL.n506 0.388379
R1127 VTAIL.n530 VTAIL.n528 0.388379
R1128 VTAIL.n479 VTAIL.n406 0.388379
R1129 VTAIL.n476 VTAIL.n408 0.388379
R1130 VTAIL.n432 VTAIL.n430 0.388379
R1131 VTAIL.n379 VTAIL.n306 0.388379
R1132 VTAIL.n376 VTAIL.n308 0.388379
R1133 VTAIL.n332 VTAIL.n330 0.388379
R1134 VTAIL.n731 VTAIL.n723 0.155672
R1135 VTAIL.n732 VTAIL.n731 0.155672
R1136 VTAIL.n732 VTAIL.n719 0.155672
R1137 VTAIL.n739 VTAIL.n719 0.155672
R1138 VTAIL.n740 VTAIL.n739 0.155672
R1139 VTAIL.n740 VTAIL.n715 0.155672
R1140 VTAIL.n747 VTAIL.n715 0.155672
R1141 VTAIL.n748 VTAIL.n747 0.155672
R1142 VTAIL.n748 VTAIL.n711 0.155672
R1143 VTAIL.n755 VTAIL.n711 0.155672
R1144 VTAIL.n756 VTAIL.n755 0.155672
R1145 VTAIL.n756 VTAIL.n707 0.155672
R1146 VTAIL.n763 VTAIL.n707 0.155672
R1147 VTAIL.n764 VTAIL.n763 0.155672
R1148 VTAIL.n764 VTAIL.n703 0.155672
R1149 VTAIL.n773 VTAIL.n703 0.155672
R1150 VTAIL.n774 VTAIL.n773 0.155672
R1151 VTAIL.n774 VTAIL.n699 0.155672
R1152 VTAIL.n781 VTAIL.n699 0.155672
R1153 VTAIL.n782 VTAIL.n781 0.155672
R1154 VTAIL.n782 VTAIL.n695 0.155672
R1155 VTAIL.n789 VTAIL.n695 0.155672
R1156 VTAIL.n39 VTAIL.n31 0.155672
R1157 VTAIL.n40 VTAIL.n39 0.155672
R1158 VTAIL.n40 VTAIL.n27 0.155672
R1159 VTAIL.n47 VTAIL.n27 0.155672
R1160 VTAIL.n48 VTAIL.n47 0.155672
R1161 VTAIL.n48 VTAIL.n23 0.155672
R1162 VTAIL.n55 VTAIL.n23 0.155672
R1163 VTAIL.n56 VTAIL.n55 0.155672
R1164 VTAIL.n56 VTAIL.n19 0.155672
R1165 VTAIL.n63 VTAIL.n19 0.155672
R1166 VTAIL.n64 VTAIL.n63 0.155672
R1167 VTAIL.n64 VTAIL.n15 0.155672
R1168 VTAIL.n71 VTAIL.n15 0.155672
R1169 VTAIL.n72 VTAIL.n71 0.155672
R1170 VTAIL.n72 VTAIL.n11 0.155672
R1171 VTAIL.n81 VTAIL.n11 0.155672
R1172 VTAIL.n82 VTAIL.n81 0.155672
R1173 VTAIL.n82 VTAIL.n7 0.155672
R1174 VTAIL.n89 VTAIL.n7 0.155672
R1175 VTAIL.n90 VTAIL.n89 0.155672
R1176 VTAIL.n90 VTAIL.n3 0.155672
R1177 VTAIL.n97 VTAIL.n3 0.155672
R1178 VTAIL.n137 VTAIL.n129 0.155672
R1179 VTAIL.n138 VTAIL.n137 0.155672
R1180 VTAIL.n138 VTAIL.n125 0.155672
R1181 VTAIL.n145 VTAIL.n125 0.155672
R1182 VTAIL.n146 VTAIL.n145 0.155672
R1183 VTAIL.n146 VTAIL.n121 0.155672
R1184 VTAIL.n153 VTAIL.n121 0.155672
R1185 VTAIL.n154 VTAIL.n153 0.155672
R1186 VTAIL.n154 VTAIL.n117 0.155672
R1187 VTAIL.n161 VTAIL.n117 0.155672
R1188 VTAIL.n162 VTAIL.n161 0.155672
R1189 VTAIL.n162 VTAIL.n113 0.155672
R1190 VTAIL.n169 VTAIL.n113 0.155672
R1191 VTAIL.n170 VTAIL.n169 0.155672
R1192 VTAIL.n170 VTAIL.n109 0.155672
R1193 VTAIL.n179 VTAIL.n109 0.155672
R1194 VTAIL.n180 VTAIL.n179 0.155672
R1195 VTAIL.n180 VTAIL.n105 0.155672
R1196 VTAIL.n187 VTAIL.n105 0.155672
R1197 VTAIL.n188 VTAIL.n187 0.155672
R1198 VTAIL.n188 VTAIL.n101 0.155672
R1199 VTAIL.n195 VTAIL.n101 0.155672
R1200 VTAIL.n237 VTAIL.n229 0.155672
R1201 VTAIL.n238 VTAIL.n237 0.155672
R1202 VTAIL.n238 VTAIL.n225 0.155672
R1203 VTAIL.n245 VTAIL.n225 0.155672
R1204 VTAIL.n246 VTAIL.n245 0.155672
R1205 VTAIL.n246 VTAIL.n221 0.155672
R1206 VTAIL.n253 VTAIL.n221 0.155672
R1207 VTAIL.n254 VTAIL.n253 0.155672
R1208 VTAIL.n254 VTAIL.n217 0.155672
R1209 VTAIL.n261 VTAIL.n217 0.155672
R1210 VTAIL.n262 VTAIL.n261 0.155672
R1211 VTAIL.n262 VTAIL.n213 0.155672
R1212 VTAIL.n269 VTAIL.n213 0.155672
R1213 VTAIL.n270 VTAIL.n269 0.155672
R1214 VTAIL.n270 VTAIL.n209 0.155672
R1215 VTAIL.n279 VTAIL.n209 0.155672
R1216 VTAIL.n280 VTAIL.n279 0.155672
R1217 VTAIL.n280 VTAIL.n205 0.155672
R1218 VTAIL.n287 VTAIL.n205 0.155672
R1219 VTAIL.n288 VTAIL.n287 0.155672
R1220 VTAIL.n288 VTAIL.n201 0.155672
R1221 VTAIL.n295 VTAIL.n201 0.155672
R1222 VTAIL.n691 VTAIL.n597 0.155672
R1223 VTAIL.n684 VTAIL.n597 0.155672
R1224 VTAIL.n684 VTAIL.n683 0.155672
R1225 VTAIL.n683 VTAIL.n601 0.155672
R1226 VTAIL.n676 VTAIL.n601 0.155672
R1227 VTAIL.n676 VTAIL.n675 0.155672
R1228 VTAIL.n675 VTAIL.n605 0.155672
R1229 VTAIL.n668 VTAIL.n605 0.155672
R1230 VTAIL.n668 VTAIL.n667 0.155672
R1231 VTAIL.n667 VTAIL.n611 0.155672
R1232 VTAIL.n660 VTAIL.n611 0.155672
R1233 VTAIL.n660 VTAIL.n659 0.155672
R1234 VTAIL.n659 VTAIL.n615 0.155672
R1235 VTAIL.n652 VTAIL.n615 0.155672
R1236 VTAIL.n652 VTAIL.n651 0.155672
R1237 VTAIL.n651 VTAIL.n619 0.155672
R1238 VTAIL.n644 VTAIL.n619 0.155672
R1239 VTAIL.n644 VTAIL.n643 0.155672
R1240 VTAIL.n643 VTAIL.n623 0.155672
R1241 VTAIL.n636 VTAIL.n623 0.155672
R1242 VTAIL.n636 VTAIL.n635 0.155672
R1243 VTAIL.n635 VTAIL.n627 0.155672
R1244 VTAIL.n591 VTAIL.n497 0.155672
R1245 VTAIL.n584 VTAIL.n497 0.155672
R1246 VTAIL.n584 VTAIL.n583 0.155672
R1247 VTAIL.n583 VTAIL.n501 0.155672
R1248 VTAIL.n576 VTAIL.n501 0.155672
R1249 VTAIL.n576 VTAIL.n575 0.155672
R1250 VTAIL.n575 VTAIL.n505 0.155672
R1251 VTAIL.n568 VTAIL.n505 0.155672
R1252 VTAIL.n568 VTAIL.n567 0.155672
R1253 VTAIL.n567 VTAIL.n511 0.155672
R1254 VTAIL.n560 VTAIL.n511 0.155672
R1255 VTAIL.n560 VTAIL.n559 0.155672
R1256 VTAIL.n559 VTAIL.n515 0.155672
R1257 VTAIL.n552 VTAIL.n515 0.155672
R1258 VTAIL.n552 VTAIL.n551 0.155672
R1259 VTAIL.n551 VTAIL.n519 0.155672
R1260 VTAIL.n544 VTAIL.n519 0.155672
R1261 VTAIL.n544 VTAIL.n543 0.155672
R1262 VTAIL.n543 VTAIL.n523 0.155672
R1263 VTAIL.n536 VTAIL.n523 0.155672
R1264 VTAIL.n536 VTAIL.n535 0.155672
R1265 VTAIL.n535 VTAIL.n527 0.155672
R1266 VTAIL.n493 VTAIL.n399 0.155672
R1267 VTAIL.n486 VTAIL.n399 0.155672
R1268 VTAIL.n486 VTAIL.n485 0.155672
R1269 VTAIL.n485 VTAIL.n403 0.155672
R1270 VTAIL.n478 VTAIL.n403 0.155672
R1271 VTAIL.n478 VTAIL.n477 0.155672
R1272 VTAIL.n477 VTAIL.n407 0.155672
R1273 VTAIL.n470 VTAIL.n407 0.155672
R1274 VTAIL.n470 VTAIL.n469 0.155672
R1275 VTAIL.n469 VTAIL.n413 0.155672
R1276 VTAIL.n462 VTAIL.n413 0.155672
R1277 VTAIL.n462 VTAIL.n461 0.155672
R1278 VTAIL.n461 VTAIL.n417 0.155672
R1279 VTAIL.n454 VTAIL.n417 0.155672
R1280 VTAIL.n454 VTAIL.n453 0.155672
R1281 VTAIL.n453 VTAIL.n421 0.155672
R1282 VTAIL.n446 VTAIL.n421 0.155672
R1283 VTAIL.n446 VTAIL.n445 0.155672
R1284 VTAIL.n445 VTAIL.n425 0.155672
R1285 VTAIL.n438 VTAIL.n425 0.155672
R1286 VTAIL.n438 VTAIL.n437 0.155672
R1287 VTAIL.n437 VTAIL.n429 0.155672
R1288 VTAIL.n393 VTAIL.n299 0.155672
R1289 VTAIL.n386 VTAIL.n299 0.155672
R1290 VTAIL.n386 VTAIL.n385 0.155672
R1291 VTAIL.n385 VTAIL.n303 0.155672
R1292 VTAIL.n378 VTAIL.n303 0.155672
R1293 VTAIL.n378 VTAIL.n377 0.155672
R1294 VTAIL.n377 VTAIL.n307 0.155672
R1295 VTAIL.n370 VTAIL.n307 0.155672
R1296 VTAIL.n370 VTAIL.n369 0.155672
R1297 VTAIL.n369 VTAIL.n313 0.155672
R1298 VTAIL.n362 VTAIL.n313 0.155672
R1299 VTAIL.n362 VTAIL.n361 0.155672
R1300 VTAIL.n361 VTAIL.n317 0.155672
R1301 VTAIL.n354 VTAIL.n317 0.155672
R1302 VTAIL.n354 VTAIL.n353 0.155672
R1303 VTAIL.n353 VTAIL.n321 0.155672
R1304 VTAIL.n346 VTAIL.n321 0.155672
R1305 VTAIL.n346 VTAIL.n345 0.155672
R1306 VTAIL.n345 VTAIL.n325 0.155672
R1307 VTAIL.n338 VTAIL.n325 0.155672
R1308 VTAIL.n338 VTAIL.n337 0.155672
R1309 VTAIL.n337 VTAIL.n329 0.155672
R1310 VTAIL VTAIL.n1 0.0586897
R1311 VDD2.n2 VDD2.n1 72.9491
R1312 VDD2.n2 VDD2.n0 72.9491
R1313 VDD2 VDD2.n5 72.9463
R1314 VDD2.n4 VDD2.n3 71.3495
R1315 VDD2.n4 VDD2.n2 53.8187
R1316 VDD2.n5 VDD2.t2 1.84319
R1317 VDD2.n5 VDD2.t3 1.84319
R1318 VDD2.n3 VDD2.t6 1.84319
R1319 VDD2.n3 VDD2.t4 1.84319
R1320 VDD2.n1 VDD2.t1 1.84319
R1321 VDD2.n1 VDD2.t7 1.84319
R1322 VDD2.n0 VDD2.t0 1.84319
R1323 VDD2.n0 VDD2.t5 1.84319
R1324 VDD2 VDD2.n4 1.71386
R1325 VP.n24 VP.n23 161.3
R1326 VP.n25 VP.n20 161.3
R1327 VP.n27 VP.n26 161.3
R1328 VP.n28 VP.n19 161.3
R1329 VP.n30 VP.n29 161.3
R1330 VP.n31 VP.n18 161.3
R1331 VP.n34 VP.n33 161.3
R1332 VP.n35 VP.n17 161.3
R1333 VP.n37 VP.n36 161.3
R1334 VP.n38 VP.n16 161.3
R1335 VP.n40 VP.n39 161.3
R1336 VP.n41 VP.n15 161.3
R1337 VP.n43 VP.n42 161.3
R1338 VP.n44 VP.n14 161.3
R1339 VP.n46 VP.n45 161.3
R1340 VP.n85 VP.n84 161.3
R1341 VP.n83 VP.n1 161.3
R1342 VP.n82 VP.n81 161.3
R1343 VP.n80 VP.n2 161.3
R1344 VP.n79 VP.n78 161.3
R1345 VP.n77 VP.n3 161.3
R1346 VP.n76 VP.n75 161.3
R1347 VP.n74 VP.n4 161.3
R1348 VP.n73 VP.n72 161.3
R1349 VP.n70 VP.n5 161.3
R1350 VP.n69 VP.n68 161.3
R1351 VP.n67 VP.n6 161.3
R1352 VP.n66 VP.n65 161.3
R1353 VP.n64 VP.n7 161.3
R1354 VP.n63 VP.n62 161.3
R1355 VP.n61 VP.n60 161.3
R1356 VP.n59 VP.n9 161.3
R1357 VP.n58 VP.n57 161.3
R1358 VP.n56 VP.n10 161.3
R1359 VP.n55 VP.n54 161.3
R1360 VP.n53 VP.n11 161.3
R1361 VP.n52 VP.n51 161.3
R1362 VP.n50 VP.n12 161.3
R1363 VP.n22 VP.t5 154.981
R1364 VP.n48 VP.t7 121.118
R1365 VP.n8 VP.t2 121.118
R1366 VP.n71 VP.t1 121.118
R1367 VP.n0 VP.t3 121.118
R1368 VP.n13 VP.t6 121.118
R1369 VP.n32 VP.t0 121.118
R1370 VP.n21 VP.t4 121.118
R1371 VP.n49 VP.n48 77.4578
R1372 VP.n86 VP.n0 77.4578
R1373 VP.n47 VP.n13 77.4578
R1374 VP.n49 VP.n47 59.5602
R1375 VP.n54 VP.n10 56.0773
R1376 VP.n78 VP.n2 56.0773
R1377 VP.n39 VP.n15 56.0773
R1378 VP.n22 VP.n21 54.2621
R1379 VP.n65 VP.n6 40.577
R1380 VP.n69 VP.n6 40.577
R1381 VP.n30 VP.n19 40.577
R1382 VP.n26 VP.n19 40.577
R1383 VP.n54 VP.n53 25.0767
R1384 VP.n82 VP.n2 25.0767
R1385 VP.n43 VP.n15 25.0767
R1386 VP.n52 VP.n12 24.5923
R1387 VP.n53 VP.n52 24.5923
R1388 VP.n58 VP.n10 24.5923
R1389 VP.n59 VP.n58 24.5923
R1390 VP.n60 VP.n59 24.5923
R1391 VP.n64 VP.n63 24.5923
R1392 VP.n65 VP.n64 24.5923
R1393 VP.n70 VP.n69 24.5923
R1394 VP.n72 VP.n70 24.5923
R1395 VP.n76 VP.n4 24.5923
R1396 VP.n77 VP.n76 24.5923
R1397 VP.n78 VP.n77 24.5923
R1398 VP.n83 VP.n82 24.5923
R1399 VP.n84 VP.n83 24.5923
R1400 VP.n44 VP.n43 24.5923
R1401 VP.n45 VP.n44 24.5923
R1402 VP.n31 VP.n30 24.5923
R1403 VP.n33 VP.n31 24.5923
R1404 VP.n37 VP.n17 24.5923
R1405 VP.n38 VP.n37 24.5923
R1406 VP.n39 VP.n38 24.5923
R1407 VP.n25 VP.n24 24.5923
R1408 VP.n26 VP.n25 24.5923
R1409 VP.n63 VP.n8 20.6576
R1410 VP.n72 VP.n71 20.6576
R1411 VP.n33 VP.n32 20.6576
R1412 VP.n24 VP.n21 20.6576
R1413 VP.n48 VP.n12 12.7883
R1414 VP.n84 VP.n0 12.7883
R1415 VP.n45 VP.n13 12.7883
R1416 VP.n60 VP.n8 3.93519
R1417 VP.n71 VP.n4 3.93519
R1418 VP.n32 VP.n17 3.93519
R1419 VP.n23 VP.n22 3.05446
R1420 VP.n47 VP.n46 0.354861
R1421 VP.n50 VP.n49 0.354861
R1422 VP.n86 VP.n85 0.354861
R1423 VP VP.n86 0.267071
R1424 VP.n23 VP.n20 0.189894
R1425 VP.n27 VP.n20 0.189894
R1426 VP.n28 VP.n27 0.189894
R1427 VP.n29 VP.n28 0.189894
R1428 VP.n29 VP.n18 0.189894
R1429 VP.n34 VP.n18 0.189894
R1430 VP.n35 VP.n34 0.189894
R1431 VP.n36 VP.n35 0.189894
R1432 VP.n36 VP.n16 0.189894
R1433 VP.n40 VP.n16 0.189894
R1434 VP.n41 VP.n40 0.189894
R1435 VP.n42 VP.n41 0.189894
R1436 VP.n42 VP.n14 0.189894
R1437 VP.n46 VP.n14 0.189894
R1438 VP.n51 VP.n50 0.189894
R1439 VP.n51 VP.n11 0.189894
R1440 VP.n55 VP.n11 0.189894
R1441 VP.n56 VP.n55 0.189894
R1442 VP.n57 VP.n56 0.189894
R1443 VP.n57 VP.n9 0.189894
R1444 VP.n61 VP.n9 0.189894
R1445 VP.n62 VP.n61 0.189894
R1446 VP.n62 VP.n7 0.189894
R1447 VP.n66 VP.n7 0.189894
R1448 VP.n67 VP.n66 0.189894
R1449 VP.n68 VP.n67 0.189894
R1450 VP.n68 VP.n5 0.189894
R1451 VP.n73 VP.n5 0.189894
R1452 VP.n74 VP.n73 0.189894
R1453 VP.n75 VP.n74 0.189894
R1454 VP.n75 VP.n3 0.189894
R1455 VP.n79 VP.n3 0.189894
R1456 VP.n80 VP.n79 0.189894
R1457 VP.n81 VP.n80 0.189894
R1458 VP.n81 VP.n1 0.189894
R1459 VP.n85 VP.n1 0.189894
R1460 VDD1 VDD1.n0 73.0629
R1461 VDD1.n3 VDD1.n2 72.9491
R1462 VDD1.n3 VDD1.n1 72.9491
R1463 VDD1.n5 VDD1.n4 71.3493
R1464 VDD1.n5 VDD1.n3 54.4018
R1465 VDD1.n4 VDD1.t7 1.84319
R1466 VDD1.n4 VDD1.t1 1.84319
R1467 VDD1.n0 VDD1.t2 1.84319
R1468 VDD1.n0 VDD1.t3 1.84319
R1469 VDD1.n2 VDD1.t6 1.84319
R1470 VDD1.n2 VDD1.t4 1.84319
R1471 VDD1.n1 VDD1.t0 1.84319
R1472 VDD1.n1 VDD1.t5 1.84319
R1473 VDD1 VDD1.n5 1.59748
R1474 B.n550 B.n549 585
R1475 B.n548 B.n167 585
R1476 B.n547 B.n546 585
R1477 B.n545 B.n168 585
R1478 B.n544 B.n543 585
R1479 B.n542 B.n169 585
R1480 B.n541 B.n540 585
R1481 B.n539 B.n170 585
R1482 B.n538 B.n537 585
R1483 B.n536 B.n171 585
R1484 B.n535 B.n534 585
R1485 B.n533 B.n172 585
R1486 B.n532 B.n531 585
R1487 B.n530 B.n173 585
R1488 B.n529 B.n528 585
R1489 B.n527 B.n174 585
R1490 B.n526 B.n525 585
R1491 B.n524 B.n175 585
R1492 B.n523 B.n522 585
R1493 B.n521 B.n176 585
R1494 B.n520 B.n519 585
R1495 B.n518 B.n177 585
R1496 B.n517 B.n516 585
R1497 B.n515 B.n178 585
R1498 B.n514 B.n513 585
R1499 B.n512 B.n179 585
R1500 B.n511 B.n510 585
R1501 B.n509 B.n180 585
R1502 B.n508 B.n507 585
R1503 B.n506 B.n181 585
R1504 B.n505 B.n504 585
R1505 B.n503 B.n182 585
R1506 B.n502 B.n501 585
R1507 B.n500 B.n183 585
R1508 B.n499 B.n498 585
R1509 B.n497 B.n184 585
R1510 B.n496 B.n495 585
R1511 B.n494 B.n185 585
R1512 B.n493 B.n492 585
R1513 B.n491 B.n186 585
R1514 B.n490 B.n489 585
R1515 B.n488 B.n187 585
R1516 B.n487 B.n486 585
R1517 B.n485 B.n188 585
R1518 B.n484 B.n483 585
R1519 B.n482 B.n189 585
R1520 B.n481 B.n480 585
R1521 B.n479 B.n190 585
R1522 B.n478 B.n477 585
R1523 B.n476 B.n191 585
R1524 B.n475 B.n474 585
R1525 B.n473 B.n192 585
R1526 B.n472 B.n471 585
R1527 B.n470 B.n193 585
R1528 B.n469 B.n468 585
R1529 B.n467 B.n194 585
R1530 B.n466 B.n465 585
R1531 B.n464 B.n195 585
R1532 B.n462 B.n461 585
R1533 B.n460 B.n198 585
R1534 B.n459 B.n458 585
R1535 B.n457 B.n199 585
R1536 B.n456 B.n455 585
R1537 B.n454 B.n200 585
R1538 B.n453 B.n452 585
R1539 B.n451 B.n201 585
R1540 B.n450 B.n449 585
R1541 B.n448 B.n202 585
R1542 B.n447 B.n446 585
R1543 B.n442 B.n203 585
R1544 B.n441 B.n440 585
R1545 B.n439 B.n204 585
R1546 B.n438 B.n437 585
R1547 B.n436 B.n205 585
R1548 B.n435 B.n434 585
R1549 B.n433 B.n206 585
R1550 B.n432 B.n431 585
R1551 B.n430 B.n207 585
R1552 B.n429 B.n428 585
R1553 B.n427 B.n208 585
R1554 B.n426 B.n425 585
R1555 B.n424 B.n209 585
R1556 B.n423 B.n422 585
R1557 B.n421 B.n210 585
R1558 B.n420 B.n419 585
R1559 B.n418 B.n211 585
R1560 B.n417 B.n416 585
R1561 B.n415 B.n212 585
R1562 B.n414 B.n413 585
R1563 B.n412 B.n213 585
R1564 B.n411 B.n410 585
R1565 B.n409 B.n214 585
R1566 B.n408 B.n407 585
R1567 B.n406 B.n215 585
R1568 B.n405 B.n404 585
R1569 B.n403 B.n216 585
R1570 B.n402 B.n401 585
R1571 B.n400 B.n217 585
R1572 B.n399 B.n398 585
R1573 B.n397 B.n218 585
R1574 B.n396 B.n395 585
R1575 B.n394 B.n219 585
R1576 B.n393 B.n392 585
R1577 B.n391 B.n220 585
R1578 B.n390 B.n389 585
R1579 B.n388 B.n221 585
R1580 B.n387 B.n386 585
R1581 B.n385 B.n222 585
R1582 B.n384 B.n383 585
R1583 B.n382 B.n223 585
R1584 B.n381 B.n380 585
R1585 B.n379 B.n224 585
R1586 B.n378 B.n377 585
R1587 B.n376 B.n225 585
R1588 B.n375 B.n374 585
R1589 B.n373 B.n226 585
R1590 B.n372 B.n371 585
R1591 B.n370 B.n227 585
R1592 B.n369 B.n368 585
R1593 B.n367 B.n228 585
R1594 B.n366 B.n365 585
R1595 B.n364 B.n229 585
R1596 B.n363 B.n362 585
R1597 B.n361 B.n230 585
R1598 B.n360 B.n359 585
R1599 B.n358 B.n231 585
R1600 B.n551 B.n166 585
R1601 B.n553 B.n552 585
R1602 B.n554 B.n165 585
R1603 B.n556 B.n555 585
R1604 B.n557 B.n164 585
R1605 B.n559 B.n558 585
R1606 B.n560 B.n163 585
R1607 B.n562 B.n561 585
R1608 B.n563 B.n162 585
R1609 B.n565 B.n564 585
R1610 B.n566 B.n161 585
R1611 B.n568 B.n567 585
R1612 B.n569 B.n160 585
R1613 B.n571 B.n570 585
R1614 B.n572 B.n159 585
R1615 B.n574 B.n573 585
R1616 B.n575 B.n158 585
R1617 B.n577 B.n576 585
R1618 B.n578 B.n157 585
R1619 B.n580 B.n579 585
R1620 B.n581 B.n156 585
R1621 B.n583 B.n582 585
R1622 B.n584 B.n155 585
R1623 B.n586 B.n585 585
R1624 B.n587 B.n154 585
R1625 B.n589 B.n588 585
R1626 B.n590 B.n153 585
R1627 B.n592 B.n591 585
R1628 B.n593 B.n152 585
R1629 B.n595 B.n594 585
R1630 B.n596 B.n151 585
R1631 B.n598 B.n597 585
R1632 B.n599 B.n150 585
R1633 B.n601 B.n600 585
R1634 B.n602 B.n149 585
R1635 B.n604 B.n603 585
R1636 B.n605 B.n148 585
R1637 B.n607 B.n606 585
R1638 B.n608 B.n147 585
R1639 B.n610 B.n609 585
R1640 B.n611 B.n146 585
R1641 B.n613 B.n612 585
R1642 B.n614 B.n145 585
R1643 B.n616 B.n615 585
R1644 B.n617 B.n144 585
R1645 B.n619 B.n618 585
R1646 B.n620 B.n143 585
R1647 B.n622 B.n621 585
R1648 B.n623 B.n142 585
R1649 B.n625 B.n624 585
R1650 B.n626 B.n141 585
R1651 B.n628 B.n627 585
R1652 B.n629 B.n140 585
R1653 B.n631 B.n630 585
R1654 B.n632 B.n139 585
R1655 B.n634 B.n633 585
R1656 B.n635 B.n138 585
R1657 B.n637 B.n636 585
R1658 B.n638 B.n137 585
R1659 B.n640 B.n639 585
R1660 B.n641 B.n136 585
R1661 B.n643 B.n642 585
R1662 B.n644 B.n135 585
R1663 B.n646 B.n645 585
R1664 B.n647 B.n134 585
R1665 B.n649 B.n648 585
R1666 B.n650 B.n133 585
R1667 B.n652 B.n651 585
R1668 B.n653 B.n132 585
R1669 B.n655 B.n654 585
R1670 B.n656 B.n131 585
R1671 B.n658 B.n657 585
R1672 B.n659 B.n130 585
R1673 B.n661 B.n660 585
R1674 B.n662 B.n129 585
R1675 B.n664 B.n663 585
R1676 B.n665 B.n128 585
R1677 B.n667 B.n666 585
R1678 B.n668 B.n127 585
R1679 B.n670 B.n669 585
R1680 B.n671 B.n126 585
R1681 B.n673 B.n672 585
R1682 B.n674 B.n125 585
R1683 B.n676 B.n675 585
R1684 B.n677 B.n124 585
R1685 B.n679 B.n678 585
R1686 B.n680 B.n123 585
R1687 B.n682 B.n681 585
R1688 B.n683 B.n122 585
R1689 B.n685 B.n684 585
R1690 B.n686 B.n121 585
R1691 B.n688 B.n687 585
R1692 B.n689 B.n120 585
R1693 B.n691 B.n690 585
R1694 B.n692 B.n119 585
R1695 B.n694 B.n693 585
R1696 B.n695 B.n118 585
R1697 B.n697 B.n696 585
R1698 B.n698 B.n117 585
R1699 B.n700 B.n699 585
R1700 B.n701 B.n116 585
R1701 B.n703 B.n702 585
R1702 B.n704 B.n115 585
R1703 B.n706 B.n705 585
R1704 B.n707 B.n114 585
R1705 B.n709 B.n708 585
R1706 B.n710 B.n113 585
R1707 B.n712 B.n711 585
R1708 B.n713 B.n112 585
R1709 B.n715 B.n714 585
R1710 B.n716 B.n111 585
R1711 B.n718 B.n717 585
R1712 B.n719 B.n110 585
R1713 B.n721 B.n720 585
R1714 B.n722 B.n109 585
R1715 B.n724 B.n723 585
R1716 B.n725 B.n108 585
R1717 B.n727 B.n726 585
R1718 B.n728 B.n107 585
R1719 B.n730 B.n729 585
R1720 B.n731 B.n106 585
R1721 B.n733 B.n732 585
R1722 B.n734 B.n105 585
R1723 B.n736 B.n735 585
R1724 B.n737 B.n104 585
R1725 B.n739 B.n738 585
R1726 B.n740 B.n103 585
R1727 B.n742 B.n741 585
R1728 B.n743 B.n102 585
R1729 B.n745 B.n744 585
R1730 B.n935 B.n34 585
R1731 B.n934 B.n933 585
R1732 B.n932 B.n35 585
R1733 B.n931 B.n930 585
R1734 B.n929 B.n36 585
R1735 B.n928 B.n927 585
R1736 B.n926 B.n37 585
R1737 B.n925 B.n924 585
R1738 B.n923 B.n38 585
R1739 B.n922 B.n921 585
R1740 B.n920 B.n39 585
R1741 B.n919 B.n918 585
R1742 B.n917 B.n40 585
R1743 B.n916 B.n915 585
R1744 B.n914 B.n41 585
R1745 B.n913 B.n912 585
R1746 B.n911 B.n42 585
R1747 B.n910 B.n909 585
R1748 B.n908 B.n43 585
R1749 B.n907 B.n906 585
R1750 B.n905 B.n44 585
R1751 B.n904 B.n903 585
R1752 B.n902 B.n45 585
R1753 B.n901 B.n900 585
R1754 B.n899 B.n46 585
R1755 B.n898 B.n897 585
R1756 B.n896 B.n47 585
R1757 B.n895 B.n894 585
R1758 B.n893 B.n48 585
R1759 B.n892 B.n891 585
R1760 B.n890 B.n49 585
R1761 B.n889 B.n888 585
R1762 B.n887 B.n50 585
R1763 B.n886 B.n885 585
R1764 B.n884 B.n51 585
R1765 B.n883 B.n882 585
R1766 B.n881 B.n52 585
R1767 B.n880 B.n879 585
R1768 B.n878 B.n53 585
R1769 B.n877 B.n876 585
R1770 B.n875 B.n54 585
R1771 B.n874 B.n873 585
R1772 B.n872 B.n55 585
R1773 B.n871 B.n870 585
R1774 B.n869 B.n56 585
R1775 B.n868 B.n867 585
R1776 B.n866 B.n57 585
R1777 B.n865 B.n864 585
R1778 B.n863 B.n58 585
R1779 B.n862 B.n861 585
R1780 B.n860 B.n59 585
R1781 B.n859 B.n858 585
R1782 B.n857 B.n60 585
R1783 B.n856 B.n855 585
R1784 B.n854 B.n61 585
R1785 B.n853 B.n852 585
R1786 B.n851 B.n62 585
R1787 B.n850 B.n849 585
R1788 B.n847 B.n63 585
R1789 B.n846 B.n845 585
R1790 B.n844 B.n66 585
R1791 B.n843 B.n842 585
R1792 B.n841 B.n67 585
R1793 B.n840 B.n839 585
R1794 B.n838 B.n68 585
R1795 B.n837 B.n836 585
R1796 B.n835 B.n69 585
R1797 B.n834 B.n833 585
R1798 B.n832 B.n831 585
R1799 B.n830 B.n73 585
R1800 B.n829 B.n828 585
R1801 B.n827 B.n74 585
R1802 B.n826 B.n825 585
R1803 B.n824 B.n75 585
R1804 B.n823 B.n822 585
R1805 B.n821 B.n76 585
R1806 B.n820 B.n819 585
R1807 B.n818 B.n77 585
R1808 B.n817 B.n816 585
R1809 B.n815 B.n78 585
R1810 B.n814 B.n813 585
R1811 B.n812 B.n79 585
R1812 B.n811 B.n810 585
R1813 B.n809 B.n80 585
R1814 B.n808 B.n807 585
R1815 B.n806 B.n81 585
R1816 B.n805 B.n804 585
R1817 B.n803 B.n82 585
R1818 B.n802 B.n801 585
R1819 B.n800 B.n83 585
R1820 B.n799 B.n798 585
R1821 B.n797 B.n84 585
R1822 B.n796 B.n795 585
R1823 B.n794 B.n85 585
R1824 B.n793 B.n792 585
R1825 B.n791 B.n86 585
R1826 B.n790 B.n789 585
R1827 B.n788 B.n87 585
R1828 B.n787 B.n786 585
R1829 B.n785 B.n88 585
R1830 B.n784 B.n783 585
R1831 B.n782 B.n89 585
R1832 B.n781 B.n780 585
R1833 B.n779 B.n90 585
R1834 B.n778 B.n777 585
R1835 B.n776 B.n91 585
R1836 B.n775 B.n774 585
R1837 B.n773 B.n92 585
R1838 B.n772 B.n771 585
R1839 B.n770 B.n93 585
R1840 B.n769 B.n768 585
R1841 B.n767 B.n94 585
R1842 B.n766 B.n765 585
R1843 B.n764 B.n95 585
R1844 B.n763 B.n762 585
R1845 B.n761 B.n96 585
R1846 B.n760 B.n759 585
R1847 B.n758 B.n97 585
R1848 B.n757 B.n756 585
R1849 B.n755 B.n98 585
R1850 B.n754 B.n753 585
R1851 B.n752 B.n99 585
R1852 B.n751 B.n750 585
R1853 B.n749 B.n100 585
R1854 B.n748 B.n747 585
R1855 B.n746 B.n101 585
R1856 B.n937 B.n936 585
R1857 B.n938 B.n33 585
R1858 B.n940 B.n939 585
R1859 B.n941 B.n32 585
R1860 B.n943 B.n942 585
R1861 B.n944 B.n31 585
R1862 B.n946 B.n945 585
R1863 B.n947 B.n30 585
R1864 B.n949 B.n948 585
R1865 B.n950 B.n29 585
R1866 B.n952 B.n951 585
R1867 B.n953 B.n28 585
R1868 B.n955 B.n954 585
R1869 B.n956 B.n27 585
R1870 B.n958 B.n957 585
R1871 B.n959 B.n26 585
R1872 B.n961 B.n960 585
R1873 B.n962 B.n25 585
R1874 B.n964 B.n963 585
R1875 B.n965 B.n24 585
R1876 B.n967 B.n966 585
R1877 B.n968 B.n23 585
R1878 B.n970 B.n969 585
R1879 B.n971 B.n22 585
R1880 B.n973 B.n972 585
R1881 B.n974 B.n21 585
R1882 B.n976 B.n975 585
R1883 B.n977 B.n20 585
R1884 B.n979 B.n978 585
R1885 B.n980 B.n19 585
R1886 B.n982 B.n981 585
R1887 B.n983 B.n18 585
R1888 B.n985 B.n984 585
R1889 B.n986 B.n17 585
R1890 B.n988 B.n987 585
R1891 B.n989 B.n16 585
R1892 B.n991 B.n990 585
R1893 B.n992 B.n15 585
R1894 B.n994 B.n993 585
R1895 B.n995 B.n14 585
R1896 B.n997 B.n996 585
R1897 B.n998 B.n13 585
R1898 B.n1000 B.n999 585
R1899 B.n1001 B.n12 585
R1900 B.n1003 B.n1002 585
R1901 B.n1004 B.n11 585
R1902 B.n1006 B.n1005 585
R1903 B.n1007 B.n10 585
R1904 B.n1009 B.n1008 585
R1905 B.n1010 B.n9 585
R1906 B.n1012 B.n1011 585
R1907 B.n1013 B.n8 585
R1908 B.n1015 B.n1014 585
R1909 B.n1016 B.n7 585
R1910 B.n1018 B.n1017 585
R1911 B.n1019 B.n6 585
R1912 B.n1021 B.n1020 585
R1913 B.n1022 B.n5 585
R1914 B.n1024 B.n1023 585
R1915 B.n1025 B.n4 585
R1916 B.n1027 B.n1026 585
R1917 B.n1028 B.n3 585
R1918 B.n1030 B.n1029 585
R1919 B.n1031 B.n0 585
R1920 B.n2 B.n1 585
R1921 B.n264 B.n263 585
R1922 B.n265 B.n262 585
R1923 B.n267 B.n266 585
R1924 B.n268 B.n261 585
R1925 B.n270 B.n269 585
R1926 B.n271 B.n260 585
R1927 B.n273 B.n272 585
R1928 B.n274 B.n259 585
R1929 B.n276 B.n275 585
R1930 B.n277 B.n258 585
R1931 B.n279 B.n278 585
R1932 B.n280 B.n257 585
R1933 B.n282 B.n281 585
R1934 B.n283 B.n256 585
R1935 B.n285 B.n284 585
R1936 B.n286 B.n255 585
R1937 B.n288 B.n287 585
R1938 B.n289 B.n254 585
R1939 B.n291 B.n290 585
R1940 B.n292 B.n253 585
R1941 B.n294 B.n293 585
R1942 B.n295 B.n252 585
R1943 B.n297 B.n296 585
R1944 B.n298 B.n251 585
R1945 B.n300 B.n299 585
R1946 B.n301 B.n250 585
R1947 B.n303 B.n302 585
R1948 B.n304 B.n249 585
R1949 B.n306 B.n305 585
R1950 B.n307 B.n248 585
R1951 B.n309 B.n308 585
R1952 B.n310 B.n247 585
R1953 B.n312 B.n311 585
R1954 B.n313 B.n246 585
R1955 B.n315 B.n314 585
R1956 B.n316 B.n245 585
R1957 B.n318 B.n317 585
R1958 B.n319 B.n244 585
R1959 B.n321 B.n320 585
R1960 B.n322 B.n243 585
R1961 B.n324 B.n323 585
R1962 B.n325 B.n242 585
R1963 B.n327 B.n326 585
R1964 B.n328 B.n241 585
R1965 B.n330 B.n329 585
R1966 B.n331 B.n240 585
R1967 B.n333 B.n332 585
R1968 B.n334 B.n239 585
R1969 B.n336 B.n335 585
R1970 B.n337 B.n238 585
R1971 B.n339 B.n338 585
R1972 B.n340 B.n237 585
R1973 B.n342 B.n341 585
R1974 B.n343 B.n236 585
R1975 B.n345 B.n344 585
R1976 B.n346 B.n235 585
R1977 B.n348 B.n347 585
R1978 B.n349 B.n234 585
R1979 B.n351 B.n350 585
R1980 B.n352 B.n233 585
R1981 B.n354 B.n353 585
R1982 B.n355 B.n232 585
R1983 B.n357 B.n356 585
R1984 B.n196 B.t1 551.865
R1985 B.n70 B.t8 551.865
R1986 B.n443 B.t10 551.865
R1987 B.n64 B.t5 551.865
R1988 B.n356 B.n231 511.721
R1989 B.n551 B.n550 511.721
R1990 B.n744 B.n101 511.721
R1991 B.n936 B.n935 511.721
R1992 B.n197 B.t2 477.392
R1993 B.n71 B.t7 477.392
R1994 B.n444 B.t11 477.392
R1995 B.n65 B.t4 477.392
R1996 B.n443 B.t9 330.221
R1997 B.n196 B.t0 330.221
R1998 B.n70 B.t6 330.221
R1999 B.n64 B.t3 330.221
R2000 B.n1033 B.n1032 256.663
R2001 B.n1032 B.n1031 235.042
R2002 B.n1032 B.n2 235.042
R2003 B.n360 B.n231 163.367
R2004 B.n361 B.n360 163.367
R2005 B.n362 B.n361 163.367
R2006 B.n362 B.n229 163.367
R2007 B.n366 B.n229 163.367
R2008 B.n367 B.n366 163.367
R2009 B.n368 B.n367 163.367
R2010 B.n368 B.n227 163.367
R2011 B.n372 B.n227 163.367
R2012 B.n373 B.n372 163.367
R2013 B.n374 B.n373 163.367
R2014 B.n374 B.n225 163.367
R2015 B.n378 B.n225 163.367
R2016 B.n379 B.n378 163.367
R2017 B.n380 B.n379 163.367
R2018 B.n380 B.n223 163.367
R2019 B.n384 B.n223 163.367
R2020 B.n385 B.n384 163.367
R2021 B.n386 B.n385 163.367
R2022 B.n386 B.n221 163.367
R2023 B.n390 B.n221 163.367
R2024 B.n391 B.n390 163.367
R2025 B.n392 B.n391 163.367
R2026 B.n392 B.n219 163.367
R2027 B.n396 B.n219 163.367
R2028 B.n397 B.n396 163.367
R2029 B.n398 B.n397 163.367
R2030 B.n398 B.n217 163.367
R2031 B.n402 B.n217 163.367
R2032 B.n403 B.n402 163.367
R2033 B.n404 B.n403 163.367
R2034 B.n404 B.n215 163.367
R2035 B.n408 B.n215 163.367
R2036 B.n409 B.n408 163.367
R2037 B.n410 B.n409 163.367
R2038 B.n410 B.n213 163.367
R2039 B.n414 B.n213 163.367
R2040 B.n415 B.n414 163.367
R2041 B.n416 B.n415 163.367
R2042 B.n416 B.n211 163.367
R2043 B.n420 B.n211 163.367
R2044 B.n421 B.n420 163.367
R2045 B.n422 B.n421 163.367
R2046 B.n422 B.n209 163.367
R2047 B.n426 B.n209 163.367
R2048 B.n427 B.n426 163.367
R2049 B.n428 B.n427 163.367
R2050 B.n428 B.n207 163.367
R2051 B.n432 B.n207 163.367
R2052 B.n433 B.n432 163.367
R2053 B.n434 B.n433 163.367
R2054 B.n434 B.n205 163.367
R2055 B.n438 B.n205 163.367
R2056 B.n439 B.n438 163.367
R2057 B.n440 B.n439 163.367
R2058 B.n440 B.n203 163.367
R2059 B.n447 B.n203 163.367
R2060 B.n448 B.n447 163.367
R2061 B.n449 B.n448 163.367
R2062 B.n449 B.n201 163.367
R2063 B.n453 B.n201 163.367
R2064 B.n454 B.n453 163.367
R2065 B.n455 B.n454 163.367
R2066 B.n455 B.n199 163.367
R2067 B.n459 B.n199 163.367
R2068 B.n460 B.n459 163.367
R2069 B.n461 B.n460 163.367
R2070 B.n461 B.n195 163.367
R2071 B.n466 B.n195 163.367
R2072 B.n467 B.n466 163.367
R2073 B.n468 B.n467 163.367
R2074 B.n468 B.n193 163.367
R2075 B.n472 B.n193 163.367
R2076 B.n473 B.n472 163.367
R2077 B.n474 B.n473 163.367
R2078 B.n474 B.n191 163.367
R2079 B.n478 B.n191 163.367
R2080 B.n479 B.n478 163.367
R2081 B.n480 B.n479 163.367
R2082 B.n480 B.n189 163.367
R2083 B.n484 B.n189 163.367
R2084 B.n485 B.n484 163.367
R2085 B.n486 B.n485 163.367
R2086 B.n486 B.n187 163.367
R2087 B.n490 B.n187 163.367
R2088 B.n491 B.n490 163.367
R2089 B.n492 B.n491 163.367
R2090 B.n492 B.n185 163.367
R2091 B.n496 B.n185 163.367
R2092 B.n497 B.n496 163.367
R2093 B.n498 B.n497 163.367
R2094 B.n498 B.n183 163.367
R2095 B.n502 B.n183 163.367
R2096 B.n503 B.n502 163.367
R2097 B.n504 B.n503 163.367
R2098 B.n504 B.n181 163.367
R2099 B.n508 B.n181 163.367
R2100 B.n509 B.n508 163.367
R2101 B.n510 B.n509 163.367
R2102 B.n510 B.n179 163.367
R2103 B.n514 B.n179 163.367
R2104 B.n515 B.n514 163.367
R2105 B.n516 B.n515 163.367
R2106 B.n516 B.n177 163.367
R2107 B.n520 B.n177 163.367
R2108 B.n521 B.n520 163.367
R2109 B.n522 B.n521 163.367
R2110 B.n522 B.n175 163.367
R2111 B.n526 B.n175 163.367
R2112 B.n527 B.n526 163.367
R2113 B.n528 B.n527 163.367
R2114 B.n528 B.n173 163.367
R2115 B.n532 B.n173 163.367
R2116 B.n533 B.n532 163.367
R2117 B.n534 B.n533 163.367
R2118 B.n534 B.n171 163.367
R2119 B.n538 B.n171 163.367
R2120 B.n539 B.n538 163.367
R2121 B.n540 B.n539 163.367
R2122 B.n540 B.n169 163.367
R2123 B.n544 B.n169 163.367
R2124 B.n545 B.n544 163.367
R2125 B.n546 B.n545 163.367
R2126 B.n546 B.n167 163.367
R2127 B.n550 B.n167 163.367
R2128 B.n744 B.n743 163.367
R2129 B.n743 B.n742 163.367
R2130 B.n742 B.n103 163.367
R2131 B.n738 B.n103 163.367
R2132 B.n738 B.n737 163.367
R2133 B.n737 B.n736 163.367
R2134 B.n736 B.n105 163.367
R2135 B.n732 B.n105 163.367
R2136 B.n732 B.n731 163.367
R2137 B.n731 B.n730 163.367
R2138 B.n730 B.n107 163.367
R2139 B.n726 B.n107 163.367
R2140 B.n726 B.n725 163.367
R2141 B.n725 B.n724 163.367
R2142 B.n724 B.n109 163.367
R2143 B.n720 B.n109 163.367
R2144 B.n720 B.n719 163.367
R2145 B.n719 B.n718 163.367
R2146 B.n718 B.n111 163.367
R2147 B.n714 B.n111 163.367
R2148 B.n714 B.n713 163.367
R2149 B.n713 B.n712 163.367
R2150 B.n712 B.n113 163.367
R2151 B.n708 B.n113 163.367
R2152 B.n708 B.n707 163.367
R2153 B.n707 B.n706 163.367
R2154 B.n706 B.n115 163.367
R2155 B.n702 B.n115 163.367
R2156 B.n702 B.n701 163.367
R2157 B.n701 B.n700 163.367
R2158 B.n700 B.n117 163.367
R2159 B.n696 B.n117 163.367
R2160 B.n696 B.n695 163.367
R2161 B.n695 B.n694 163.367
R2162 B.n694 B.n119 163.367
R2163 B.n690 B.n119 163.367
R2164 B.n690 B.n689 163.367
R2165 B.n689 B.n688 163.367
R2166 B.n688 B.n121 163.367
R2167 B.n684 B.n121 163.367
R2168 B.n684 B.n683 163.367
R2169 B.n683 B.n682 163.367
R2170 B.n682 B.n123 163.367
R2171 B.n678 B.n123 163.367
R2172 B.n678 B.n677 163.367
R2173 B.n677 B.n676 163.367
R2174 B.n676 B.n125 163.367
R2175 B.n672 B.n125 163.367
R2176 B.n672 B.n671 163.367
R2177 B.n671 B.n670 163.367
R2178 B.n670 B.n127 163.367
R2179 B.n666 B.n127 163.367
R2180 B.n666 B.n665 163.367
R2181 B.n665 B.n664 163.367
R2182 B.n664 B.n129 163.367
R2183 B.n660 B.n129 163.367
R2184 B.n660 B.n659 163.367
R2185 B.n659 B.n658 163.367
R2186 B.n658 B.n131 163.367
R2187 B.n654 B.n131 163.367
R2188 B.n654 B.n653 163.367
R2189 B.n653 B.n652 163.367
R2190 B.n652 B.n133 163.367
R2191 B.n648 B.n133 163.367
R2192 B.n648 B.n647 163.367
R2193 B.n647 B.n646 163.367
R2194 B.n646 B.n135 163.367
R2195 B.n642 B.n135 163.367
R2196 B.n642 B.n641 163.367
R2197 B.n641 B.n640 163.367
R2198 B.n640 B.n137 163.367
R2199 B.n636 B.n137 163.367
R2200 B.n636 B.n635 163.367
R2201 B.n635 B.n634 163.367
R2202 B.n634 B.n139 163.367
R2203 B.n630 B.n139 163.367
R2204 B.n630 B.n629 163.367
R2205 B.n629 B.n628 163.367
R2206 B.n628 B.n141 163.367
R2207 B.n624 B.n141 163.367
R2208 B.n624 B.n623 163.367
R2209 B.n623 B.n622 163.367
R2210 B.n622 B.n143 163.367
R2211 B.n618 B.n143 163.367
R2212 B.n618 B.n617 163.367
R2213 B.n617 B.n616 163.367
R2214 B.n616 B.n145 163.367
R2215 B.n612 B.n145 163.367
R2216 B.n612 B.n611 163.367
R2217 B.n611 B.n610 163.367
R2218 B.n610 B.n147 163.367
R2219 B.n606 B.n147 163.367
R2220 B.n606 B.n605 163.367
R2221 B.n605 B.n604 163.367
R2222 B.n604 B.n149 163.367
R2223 B.n600 B.n149 163.367
R2224 B.n600 B.n599 163.367
R2225 B.n599 B.n598 163.367
R2226 B.n598 B.n151 163.367
R2227 B.n594 B.n151 163.367
R2228 B.n594 B.n593 163.367
R2229 B.n593 B.n592 163.367
R2230 B.n592 B.n153 163.367
R2231 B.n588 B.n153 163.367
R2232 B.n588 B.n587 163.367
R2233 B.n587 B.n586 163.367
R2234 B.n586 B.n155 163.367
R2235 B.n582 B.n155 163.367
R2236 B.n582 B.n581 163.367
R2237 B.n581 B.n580 163.367
R2238 B.n580 B.n157 163.367
R2239 B.n576 B.n157 163.367
R2240 B.n576 B.n575 163.367
R2241 B.n575 B.n574 163.367
R2242 B.n574 B.n159 163.367
R2243 B.n570 B.n159 163.367
R2244 B.n570 B.n569 163.367
R2245 B.n569 B.n568 163.367
R2246 B.n568 B.n161 163.367
R2247 B.n564 B.n161 163.367
R2248 B.n564 B.n563 163.367
R2249 B.n563 B.n562 163.367
R2250 B.n562 B.n163 163.367
R2251 B.n558 B.n163 163.367
R2252 B.n558 B.n557 163.367
R2253 B.n557 B.n556 163.367
R2254 B.n556 B.n165 163.367
R2255 B.n552 B.n165 163.367
R2256 B.n552 B.n551 163.367
R2257 B.n935 B.n934 163.367
R2258 B.n934 B.n35 163.367
R2259 B.n930 B.n35 163.367
R2260 B.n930 B.n929 163.367
R2261 B.n929 B.n928 163.367
R2262 B.n928 B.n37 163.367
R2263 B.n924 B.n37 163.367
R2264 B.n924 B.n923 163.367
R2265 B.n923 B.n922 163.367
R2266 B.n922 B.n39 163.367
R2267 B.n918 B.n39 163.367
R2268 B.n918 B.n917 163.367
R2269 B.n917 B.n916 163.367
R2270 B.n916 B.n41 163.367
R2271 B.n912 B.n41 163.367
R2272 B.n912 B.n911 163.367
R2273 B.n911 B.n910 163.367
R2274 B.n910 B.n43 163.367
R2275 B.n906 B.n43 163.367
R2276 B.n906 B.n905 163.367
R2277 B.n905 B.n904 163.367
R2278 B.n904 B.n45 163.367
R2279 B.n900 B.n45 163.367
R2280 B.n900 B.n899 163.367
R2281 B.n899 B.n898 163.367
R2282 B.n898 B.n47 163.367
R2283 B.n894 B.n47 163.367
R2284 B.n894 B.n893 163.367
R2285 B.n893 B.n892 163.367
R2286 B.n892 B.n49 163.367
R2287 B.n888 B.n49 163.367
R2288 B.n888 B.n887 163.367
R2289 B.n887 B.n886 163.367
R2290 B.n886 B.n51 163.367
R2291 B.n882 B.n51 163.367
R2292 B.n882 B.n881 163.367
R2293 B.n881 B.n880 163.367
R2294 B.n880 B.n53 163.367
R2295 B.n876 B.n53 163.367
R2296 B.n876 B.n875 163.367
R2297 B.n875 B.n874 163.367
R2298 B.n874 B.n55 163.367
R2299 B.n870 B.n55 163.367
R2300 B.n870 B.n869 163.367
R2301 B.n869 B.n868 163.367
R2302 B.n868 B.n57 163.367
R2303 B.n864 B.n57 163.367
R2304 B.n864 B.n863 163.367
R2305 B.n863 B.n862 163.367
R2306 B.n862 B.n59 163.367
R2307 B.n858 B.n59 163.367
R2308 B.n858 B.n857 163.367
R2309 B.n857 B.n856 163.367
R2310 B.n856 B.n61 163.367
R2311 B.n852 B.n61 163.367
R2312 B.n852 B.n851 163.367
R2313 B.n851 B.n850 163.367
R2314 B.n850 B.n63 163.367
R2315 B.n845 B.n63 163.367
R2316 B.n845 B.n844 163.367
R2317 B.n844 B.n843 163.367
R2318 B.n843 B.n67 163.367
R2319 B.n839 B.n67 163.367
R2320 B.n839 B.n838 163.367
R2321 B.n838 B.n837 163.367
R2322 B.n837 B.n69 163.367
R2323 B.n833 B.n69 163.367
R2324 B.n833 B.n832 163.367
R2325 B.n832 B.n73 163.367
R2326 B.n828 B.n73 163.367
R2327 B.n828 B.n827 163.367
R2328 B.n827 B.n826 163.367
R2329 B.n826 B.n75 163.367
R2330 B.n822 B.n75 163.367
R2331 B.n822 B.n821 163.367
R2332 B.n821 B.n820 163.367
R2333 B.n820 B.n77 163.367
R2334 B.n816 B.n77 163.367
R2335 B.n816 B.n815 163.367
R2336 B.n815 B.n814 163.367
R2337 B.n814 B.n79 163.367
R2338 B.n810 B.n79 163.367
R2339 B.n810 B.n809 163.367
R2340 B.n809 B.n808 163.367
R2341 B.n808 B.n81 163.367
R2342 B.n804 B.n81 163.367
R2343 B.n804 B.n803 163.367
R2344 B.n803 B.n802 163.367
R2345 B.n802 B.n83 163.367
R2346 B.n798 B.n83 163.367
R2347 B.n798 B.n797 163.367
R2348 B.n797 B.n796 163.367
R2349 B.n796 B.n85 163.367
R2350 B.n792 B.n85 163.367
R2351 B.n792 B.n791 163.367
R2352 B.n791 B.n790 163.367
R2353 B.n790 B.n87 163.367
R2354 B.n786 B.n87 163.367
R2355 B.n786 B.n785 163.367
R2356 B.n785 B.n784 163.367
R2357 B.n784 B.n89 163.367
R2358 B.n780 B.n89 163.367
R2359 B.n780 B.n779 163.367
R2360 B.n779 B.n778 163.367
R2361 B.n778 B.n91 163.367
R2362 B.n774 B.n91 163.367
R2363 B.n774 B.n773 163.367
R2364 B.n773 B.n772 163.367
R2365 B.n772 B.n93 163.367
R2366 B.n768 B.n93 163.367
R2367 B.n768 B.n767 163.367
R2368 B.n767 B.n766 163.367
R2369 B.n766 B.n95 163.367
R2370 B.n762 B.n95 163.367
R2371 B.n762 B.n761 163.367
R2372 B.n761 B.n760 163.367
R2373 B.n760 B.n97 163.367
R2374 B.n756 B.n97 163.367
R2375 B.n756 B.n755 163.367
R2376 B.n755 B.n754 163.367
R2377 B.n754 B.n99 163.367
R2378 B.n750 B.n99 163.367
R2379 B.n750 B.n749 163.367
R2380 B.n749 B.n748 163.367
R2381 B.n748 B.n101 163.367
R2382 B.n936 B.n33 163.367
R2383 B.n940 B.n33 163.367
R2384 B.n941 B.n940 163.367
R2385 B.n942 B.n941 163.367
R2386 B.n942 B.n31 163.367
R2387 B.n946 B.n31 163.367
R2388 B.n947 B.n946 163.367
R2389 B.n948 B.n947 163.367
R2390 B.n948 B.n29 163.367
R2391 B.n952 B.n29 163.367
R2392 B.n953 B.n952 163.367
R2393 B.n954 B.n953 163.367
R2394 B.n954 B.n27 163.367
R2395 B.n958 B.n27 163.367
R2396 B.n959 B.n958 163.367
R2397 B.n960 B.n959 163.367
R2398 B.n960 B.n25 163.367
R2399 B.n964 B.n25 163.367
R2400 B.n965 B.n964 163.367
R2401 B.n966 B.n965 163.367
R2402 B.n966 B.n23 163.367
R2403 B.n970 B.n23 163.367
R2404 B.n971 B.n970 163.367
R2405 B.n972 B.n971 163.367
R2406 B.n972 B.n21 163.367
R2407 B.n976 B.n21 163.367
R2408 B.n977 B.n976 163.367
R2409 B.n978 B.n977 163.367
R2410 B.n978 B.n19 163.367
R2411 B.n982 B.n19 163.367
R2412 B.n983 B.n982 163.367
R2413 B.n984 B.n983 163.367
R2414 B.n984 B.n17 163.367
R2415 B.n988 B.n17 163.367
R2416 B.n989 B.n988 163.367
R2417 B.n990 B.n989 163.367
R2418 B.n990 B.n15 163.367
R2419 B.n994 B.n15 163.367
R2420 B.n995 B.n994 163.367
R2421 B.n996 B.n995 163.367
R2422 B.n996 B.n13 163.367
R2423 B.n1000 B.n13 163.367
R2424 B.n1001 B.n1000 163.367
R2425 B.n1002 B.n1001 163.367
R2426 B.n1002 B.n11 163.367
R2427 B.n1006 B.n11 163.367
R2428 B.n1007 B.n1006 163.367
R2429 B.n1008 B.n1007 163.367
R2430 B.n1008 B.n9 163.367
R2431 B.n1012 B.n9 163.367
R2432 B.n1013 B.n1012 163.367
R2433 B.n1014 B.n1013 163.367
R2434 B.n1014 B.n7 163.367
R2435 B.n1018 B.n7 163.367
R2436 B.n1019 B.n1018 163.367
R2437 B.n1020 B.n1019 163.367
R2438 B.n1020 B.n5 163.367
R2439 B.n1024 B.n5 163.367
R2440 B.n1025 B.n1024 163.367
R2441 B.n1026 B.n1025 163.367
R2442 B.n1026 B.n3 163.367
R2443 B.n1030 B.n3 163.367
R2444 B.n1031 B.n1030 163.367
R2445 B.n264 B.n2 163.367
R2446 B.n265 B.n264 163.367
R2447 B.n266 B.n265 163.367
R2448 B.n266 B.n261 163.367
R2449 B.n270 B.n261 163.367
R2450 B.n271 B.n270 163.367
R2451 B.n272 B.n271 163.367
R2452 B.n272 B.n259 163.367
R2453 B.n276 B.n259 163.367
R2454 B.n277 B.n276 163.367
R2455 B.n278 B.n277 163.367
R2456 B.n278 B.n257 163.367
R2457 B.n282 B.n257 163.367
R2458 B.n283 B.n282 163.367
R2459 B.n284 B.n283 163.367
R2460 B.n284 B.n255 163.367
R2461 B.n288 B.n255 163.367
R2462 B.n289 B.n288 163.367
R2463 B.n290 B.n289 163.367
R2464 B.n290 B.n253 163.367
R2465 B.n294 B.n253 163.367
R2466 B.n295 B.n294 163.367
R2467 B.n296 B.n295 163.367
R2468 B.n296 B.n251 163.367
R2469 B.n300 B.n251 163.367
R2470 B.n301 B.n300 163.367
R2471 B.n302 B.n301 163.367
R2472 B.n302 B.n249 163.367
R2473 B.n306 B.n249 163.367
R2474 B.n307 B.n306 163.367
R2475 B.n308 B.n307 163.367
R2476 B.n308 B.n247 163.367
R2477 B.n312 B.n247 163.367
R2478 B.n313 B.n312 163.367
R2479 B.n314 B.n313 163.367
R2480 B.n314 B.n245 163.367
R2481 B.n318 B.n245 163.367
R2482 B.n319 B.n318 163.367
R2483 B.n320 B.n319 163.367
R2484 B.n320 B.n243 163.367
R2485 B.n324 B.n243 163.367
R2486 B.n325 B.n324 163.367
R2487 B.n326 B.n325 163.367
R2488 B.n326 B.n241 163.367
R2489 B.n330 B.n241 163.367
R2490 B.n331 B.n330 163.367
R2491 B.n332 B.n331 163.367
R2492 B.n332 B.n239 163.367
R2493 B.n336 B.n239 163.367
R2494 B.n337 B.n336 163.367
R2495 B.n338 B.n337 163.367
R2496 B.n338 B.n237 163.367
R2497 B.n342 B.n237 163.367
R2498 B.n343 B.n342 163.367
R2499 B.n344 B.n343 163.367
R2500 B.n344 B.n235 163.367
R2501 B.n348 B.n235 163.367
R2502 B.n349 B.n348 163.367
R2503 B.n350 B.n349 163.367
R2504 B.n350 B.n233 163.367
R2505 B.n354 B.n233 163.367
R2506 B.n355 B.n354 163.367
R2507 B.n356 B.n355 163.367
R2508 B.n444 B.n443 74.4732
R2509 B.n197 B.n196 74.4732
R2510 B.n71 B.n70 74.4732
R2511 B.n65 B.n64 74.4732
R2512 B.n445 B.n444 59.5399
R2513 B.n463 B.n197 59.5399
R2514 B.n72 B.n71 59.5399
R2515 B.n848 B.n65 59.5399
R2516 B.n937 B.n34 33.2493
R2517 B.n746 B.n745 33.2493
R2518 B.n549 B.n166 33.2493
R2519 B.n358 B.n357 33.2493
R2520 B B.n1033 18.0485
R2521 B.n938 B.n937 10.6151
R2522 B.n939 B.n938 10.6151
R2523 B.n939 B.n32 10.6151
R2524 B.n943 B.n32 10.6151
R2525 B.n944 B.n943 10.6151
R2526 B.n945 B.n944 10.6151
R2527 B.n945 B.n30 10.6151
R2528 B.n949 B.n30 10.6151
R2529 B.n950 B.n949 10.6151
R2530 B.n951 B.n950 10.6151
R2531 B.n951 B.n28 10.6151
R2532 B.n955 B.n28 10.6151
R2533 B.n956 B.n955 10.6151
R2534 B.n957 B.n956 10.6151
R2535 B.n957 B.n26 10.6151
R2536 B.n961 B.n26 10.6151
R2537 B.n962 B.n961 10.6151
R2538 B.n963 B.n962 10.6151
R2539 B.n963 B.n24 10.6151
R2540 B.n967 B.n24 10.6151
R2541 B.n968 B.n967 10.6151
R2542 B.n969 B.n968 10.6151
R2543 B.n969 B.n22 10.6151
R2544 B.n973 B.n22 10.6151
R2545 B.n974 B.n973 10.6151
R2546 B.n975 B.n974 10.6151
R2547 B.n975 B.n20 10.6151
R2548 B.n979 B.n20 10.6151
R2549 B.n980 B.n979 10.6151
R2550 B.n981 B.n980 10.6151
R2551 B.n981 B.n18 10.6151
R2552 B.n985 B.n18 10.6151
R2553 B.n986 B.n985 10.6151
R2554 B.n987 B.n986 10.6151
R2555 B.n987 B.n16 10.6151
R2556 B.n991 B.n16 10.6151
R2557 B.n992 B.n991 10.6151
R2558 B.n993 B.n992 10.6151
R2559 B.n993 B.n14 10.6151
R2560 B.n997 B.n14 10.6151
R2561 B.n998 B.n997 10.6151
R2562 B.n999 B.n998 10.6151
R2563 B.n999 B.n12 10.6151
R2564 B.n1003 B.n12 10.6151
R2565 B.n1004 B.n1003 10.6151
R2566 B.n1005 B.n1004 10.6151
R2567 B.n1005 B.n10 10.6151
R2568 B.n1009 B.n10 10.6151
R2569 B.n1010 B.n1009 10.6151
R2570 B.n1011 B.n1010 10.6151
R2571 B.n1011 B.n8 10.6151
R2572 B.n1015 B.n8 10.6151
R2573 B.n1016 B.n1015 10.6151
R2574 B.n1017 B.n1016 10.6151
R2575 B.n1017 B.n6 10.6151
R2576 B.n1021 B.n6 10.6151
R2577 B.n1022 B.n1021 10.6151
R2578 B.n1023 B.n1022 10.6151
R2579 B.n1023 B.n4 10.6151
R2580 B.n1027 B.n4 10.6151
R2581 B.n1028 B.n1027 10.6151
R2582 B.n1029 B.n1028 10.6151
R2583 B.n1029 B.n0 10.6151
R2584 B.n933 B.n34 10.6151
R2585 B.n933 B.n932 10.6151
R2586 B.n932 B.n931 10.6151
R2587 B.n931 B.n36 10.6151
R2588 B.n927 B.n36 10.6151
R2589 B.n927 B.n926 10.6151
R2590 B.n926 B.n925 10.6151
R2591 B.n925 B.n38 10.6151
R2592 B.n921 B.n38 10.6151
R2593 B.n921 B.n920 10.6151
R2594 B.n920 B.n919 10.6151
R2595 B.n919 B.n40 10.6151
R2596 B.n915 B.n40 10.6151
R2597 B.n915 B.n914 10.6151
R2598 B.n914 B.n913 10.6151
R2599 B.n913 B.n42 10.6151
R2600 B.n909 B.n42 10.6151
R2601 B.n909 B.n908 10.6151
R2602 B.n908 B.n907 10.6151
R2603 B.n907 B.n44 10.6151
R2604 B.n903 B.n44 10.6151
R2605 B.n903 B.n902 10.6151
R2606 B.n902 B.n901 10.6151
R2607 B.n901 B.n46 10.6151
R2608 B.n897 B.n46 10.6151
R2609 B.n897 B.n896 10.6151
R2610 B.n896 B.n895 10.6151
R2611 B.n895 B.n48 10.6151
R2612 B.n891 B.n48 10.6151
R2613 B.n891 B.n890 10.6151
R2614 B.n890 B.n889 10.6151
R2615 B.n889 B.n50 10.6151
R2616 B.n885 B.n50 10.6151
R2617 B.n885 B.n884 10.6151
R2618 B.n884 B.n883 10.6151
R2619 B.n883 B.n52 10.6151
R2620 B.n879 B.n52 10.6151
R2621 B.n879 B.n878 10.6151
R2622 B.n878 B.n877 10.6151
R2623 B.n877 B.n54 10.6151
R2624 B.n873 B.n54 10.6151
R2625 B.n873 B.n872 10.6151
R2626 B.n872 B.n871 10.6151
R2627 B.n871 B.n56 10.6151
R2628 B.n867 B.n56 10.6151
R2629 B.n867 B.n866 10.6151
R2630 B.n866 B.n865 10.6151
R2631 B.n865 B.n58 10.6151
R2632 B.n861 B.n58 10.6151
R2633 B.n861 B.n860 10.6151
R2634 B.n860 B.n859 10.6151
R2635 B.n859 B.n60 10.6151
R2636 B.n855 B.n60 10.6151
R2637 B.n855 B.n854 10.6151
R2638 B.n854 B.n853 10.6151
R2639 B.n853 B.n62 10.6151
R2640 B.n849 B.n62 10.6151
R2641 B.n847 B.n846 10.6151
R2642 B.n846 B.n66 10.6151
R2643 B.n842 B.n66 10.6151
R2644 B.n842 B.n841 10.6151
R2645 B.n841 B.n840 10.6151
R2646 B.n840 B.n68 10.6151
R2647 B.n836 B.n68 10.6151
R2648 B.n836 B.n835 10.6151
R2649 B.n835 B.n834 10.6151
R2650 B.n831 B.n830 10.6151
R2651 B.n830 B.n829 10.6151
R2652 B.n829 B.n74 10.6151
R2653 B.n825 B.n74 10.6151
R2654 B.n825 B.n824 10.6151
R2655 B.n824 B.n823 10.6151
R2656 B.n823 B.n76 10.6151
R2657 B.n819 B.n76 10.6151
R2658 B.n819 B.n818 10.6151
R2659 B.n818 B.n817 10.6151
R2660 B.n817 B.n78 10.6151
R2661 B.n813 B.n78 10.6151
R2662 B.n813 B.n812 10.6151
R2663 B.n812 B.n811 10.6151
R2664 B.n811 B.n80 10.6151
R2665 B.n807 B.n80 10.6151
R2666 B.n807 B.n806 10.6151
R2667 B.n806 B.n805 10.6151
R2668 B.n805 B.n82 10.6151
R2669 B.n801 B.n82 10.6151
R2670 B.n801 B.n800 10.6151
R2671 B.n800 B.n799 10.6151
R2672 B.n799 B.n84 10.6151
R2673 B.n795 B.n84 10.6151
R2674 B.n795 B.n794 10.6151
R2675 B.n794 B.n793 10.6151
R2676 B.n793 B.n86 10.6151
R2677 B.n789 B.n86 10.6151
R2678 B.n789 B.n788 10.6151
R2679 B.n788 B.n787 10.6151
R2680 B.n787 B.n88 10.6151
R2681 B.n783 B.n88 10.6151
R2682 B.n783 B.n782 10.6151
R2683 B.n782 B.n781 10.6151
R2684 B.n781 B.n90 10.6151
R2685 B.n777 B.n90 10.6151
R2686 B.n777 B.n776 10.6151
R2687 B.n776 B.n775 10.6151
R2688 B.n775 B.n92 10.6151
R2689 B.n771 B.n92 10.6151
R2690 B.n771 B.n770 10.6151
R2691 B.n770 B.n769 10.6151
R2692 B.n769 B.n94 10.6151
R2693 B.n765 B.n94 10.6151
R2694 B.n765 B.n764 10.6151
R2695 B.n764 B.n763 10.6151
R2696 B.n763 B.n96 10.6151
R2697 B.n759 B.n96 10.6151
R2698 B.n759 B.n758 10.6151
R2699 B.n758 B.n757 10.6151
R2700 B.n757 B.n98 10.6151
R2701 B.n753 B.n98 10.6151
R2702 B.n753 B.n752 10.6151
R2703 B.n752 B.n751 10.6151
R2704 B.n751 B.n100 10.6151
R2705 B.n747 B.n100 10.6151
R2706 B.n747 B.n746 10.6151
R2707 B.n745 B.n102 10.6151
R2708 B.n741 B.n102 10.6151
R2709 B.n741 B.n740 10.6151
R2710 B.n740 B.n739 10.6151
R2711 B.n739 B.n104 10.6151
R2712 B.n735 B.n104 10.6151
R2713 B.n735 B.n734 10.6151
R2714 B.n734 B.n733 10.6151
R2715 B.n733 B.n106 10.6151
R2716 B.n729 B.n106 10.6151
R2717 B.n729 B.n728 10.6151
R2718 B.n728 B.n727 10.6151
R2719 B.n727 B.n108 10.6151
R2720 B.n723 B.n108 10.6151
R2721 B.n723 B.n722 10.6151
R2722 B.n722 B.n721 10.6151
R2723 B.n721 B.n110 10.6151
R2724 B.n717 B.n110 10.6151
R2725 B.n717 B.n716 10.6151
R2726 B.n716 B.n715 10.6151
R2727 B.n715 B.n112 10.6151
R2728 B.n711 B.n112 10.6151
R2729 B.n711 B.n710 10.6151
R2730 B.n710 B.n709 10.6151
R2731 B.n709 B.n114 10.6151
R2732 B.n705 B.n114 10.6151
R2733 B.n705 B.n704 10.6151
R2734 B.n704 B.n703 10.6151
R2735 B.n703 B.n116 10.6151
R2736 B.n699 B.n116 10.6151
R2737 B.n699 B.n698 10.6151
R2738 B.n698 B.n697 10.6151
R2739 B.n697 B.n118 10.6151
R2740 B.n693 B.n118 10.6151
R2741 B.n693 B.n692 10.6151
R2742 B.n692 B.n691 10.6151
R2743 B.n691 B.n120 10.6151
R2744 B.n687 B.n120 10.6151
R2745 B.n687 B.n686 10.6151
R2746 B.n686 B.n685 10.6151
R2747 B.n685 B.n122 10.6151
R2748 B.n681 B.n122 10.6151
R2749 B.n681 B.n680 10.6151
R2750 B.n680 B.n679 10.6151
R2751 B.n679 B.n124 10.6151
R2752 B.n675 B.n124 10.6151
R2753 B.n675 B.n674 10.6151
R2754 B.n674 B.n673 10.6151
R2755 B.n673 B.n126 10.6151
R2756 B.n669 B.n126 10.6151
R2757 B.n669 B.n668 10.6151
R2758 B.n668 B.n667 10.6151
R2759 B.n667 B.n128 10.6151
R2760 B.n663 B.n128 10.6151
R2761 B.n663 B.n662 10.6151
R2762 B.n662 B.n661 10.6151
R2763 B.n661 B.n130 10.6151
R2764 B.n657 B.n130 10.6151
R2765 B.n657 B.n656 10.6151
R2766 B.n656 B.n655 10.6151
R2767 B.n655 B.n132 10.6151
R2768 B.n651 B.n132 10.6151
R2769 B.n651 B.n650 10.6151
R2770 B.n650 B.n649 10.6151
R2771 B.n649 B.n134 10.6151
R2772 B.n645 B.n134 10.6151
R2773 B.n645 B.n644 10.6151
R2774 B.n644 B.n643 10.6151
R2775 B.n643 B.n136 10.6151
R2776 B.n639 B.n136 10.6151
R2777 B.n639 B.n638 10.6151
R2778 B.n638 B.n637 10.6151
R2779 B.n637 B.n138 10.6151
R2780 B.n633 B.n138 10.6151
R2781 B.n633 B.n632 10.6151
R2782 B.n632 B.n631 10.6151
R2783 B.n631 B.n140 10.6151
R2784 B.n627 B.n140 10.6151
R2785 B.n627 B.n626 10.6151
R2786 B.n626 B.n625 10.6151
R2787 B.n625 B.n142 10.6151
R2788 B.n621 B.n142 10.6151
R2789 B.n621 B.n620 10.6151
R2790 B.n620 B.n619 10.6151
R2791 B.n619 B.n144 10.6151
R2792 B.n615 B.n144 10.6151
R2793 B.n615 B.n614 10.6151
R2794 B.n614 B.n613 10.6151
R2795 B.n613 B.n146 10.6151
R2796 B.n609 B.n146 10.6151
R2797 B.n609 B.n608 10.6151
R2798 B.n608 B.n607 10.6151
R2799 B.n607 B.n148 10.6151
R2800 B.n603 B.n148 10.6151
R2801 B.n603 B.n602 10.6151
R2802 B.n602 B.n601 10.6151
R2803 B.n601 B.n150 10.6151
R2804 B.n597 B.n150 10.6151
R2805 B.n597 B.n596 10.6151
R2806 B.n596 B.n595 10.6151
R2807 B.n595 B.n152 10.6151
R2808 B.n591 B.n152 10.6151
R2809 B.n591 B.n590 10.6151
R2810 B.n590 B.n589 10.6151
R2811 B.n589 B.n154 10.6151
R2812 B.n585 B.n154 10.6151
R2813 B.n585 B.n584 10.6151
R2814 B.n584 B.n583 10.6151
R2815 B.n583 B.n156 10.6151
R2816 B.n579 B.n156 10.6151
R2817 B.n579 B.n578 10.6151
R2818 B.n578 B.n577 10.6151
R2819 B.n577 B.n158 10.6151
R2820 B.n573 B.n158 10.6151
R2821 B.n573 B.n572 10.6151
R2822 B.n572 B.n571 10.6151
R2823 B.n571 B.n160 10.6151
R2824 B.n567 B.n160 10.6151
R2825 B.n567 B.n566 10.6151
R2826 B.n566 B.n565 10.6151
R2827 B.n565 B.n162 10.6151
R2828 B.n561 B.n162 10.6151
R2829 B.n561 B.n560 10.6151
R2830 B.n560 B.n559 10.6151
R2831 B.n559 B.n164 10.6151
R2832 B.n555 B.n164 10.6151
R2833 B.n555 B.n554 10.6151
R2834 B.n554 B.n553 10.6151
R2835 B.n553 B.n166 10.6151
R2836 B.n263 B.n1 10.6151
R2837 B.n263 B.n262 10.6151
R2838 B.n267 B.n262 10.6151
R2839 B.n268 B.n267 10.6151
R2840 B.n269 B.n268 10.6151
R2841 B.n269 B.n260 10.6151
R2842 B.n273 B.n260 10.6151
R2843 B.n274 B.n273 10.6151
R2844 B.n275 B.n274 10.6151
R2845 B.n275 B.n258 10.6151
R2846 B.n279 B.n258 10.6151
R2847 B.n280 B.n279 10.6151
R2848 B.n281 B.n280 10.6151
R2849 B.n281 B.n256 10.6151
R2850 B.n285 B.n256 10.6151
R2851 B.n286 B.n285 10.6151
R2852 B.n287 B.n286 10.6151
R2853 B.n287 B.n254 10.6151
R2854 B.n291 B.n254 10.6151
R2855 B.n292 B.n291 10.6151
R2856 B.n293 B.n292 10.6151
R2857 B.n293 B.n252 10.6151
R2858 B.n297 B.n252 10.6151
R2859 B.n298 B.n297 10.6151
R2860 B.n299 B.n298 10.6151
R2861 B.n299 B.n250 10.6151
R2862 B.n303 B.n250 10.6151
R2863 B.n304 B.n303 10.6151
R2864 B.n305 B.n304 10.6151
R2865 B.n305 B.n248 10.6151
R2866 B.n309 B.n248 10.6151
R2867 B.n310 B.n309 10.6151
R2868 B.n311 B.n310 10.6151
R2869 B.n311 B.n246 10.6151
R2870 B.n315 B.n246 10.6151
R2871 B.n316 B.n315 10.6151
R2872 B.n317 B.n316 10.6151
R2873 B.n317 B.n244 10.6151
R2874 B.n321 B.n244 10.6151
R2875 B.n322 B.n321 10.6151
R2876 B.n323 B.n322 10.6151
R2877 B.n323 B.n242 10.6151
R2878 B.n327 B.n242 10.6151
R2879 B.n328 B.n327 10.6151
R2880 B.n329 B.n328 10.6151
R2881 B.n329 B.n240 10.6151
R2882 B.n333 B.n240 10.6151
R2883 B.n334 B.n333 10.6151
R2884 B.n335 B.n334 10.6151
R2885 B.n335 B.n238 10.6151
R2886 B.n339 B.n238 10.6151
R2887 B.n340 B.n339 10.6151
R2888 B.n341 B.n340 10.6151
R2889 B.n341 B.n236 10.6151
R2890 B.n345 B.n236 10.6151
R2891 B.n346 B.n345 10.6151
R2892 B.n347 B.n346 10.6151
R2893 B.n347 B.n234 10.6151
R2894 B.n351 B.n234 10.6151
R2895 B.n352 B.n351 10.6151
R2896 B.n353 B.n352 10.6151
R2897 B.n353 B.n232 10.6151
R2898 B.n357 B.n232 10.6151
R2899 B.n359 B.n358 10.6151
R2900 B.n359 B.n230 10.6151
R2901 B.n363 B.n230 10.6151
R2902 B.n364 B.n363 10.6151
R2903 B.n365 B.n364 10.6151
R2904 B.n365 B.n228 10.6151
R2905 B.n369 B.n228 10.6151
R2906 B.n370 B.n369 10.6151
R2907 B.n371 B.n370 10.6151
R2908 B.n371 B.n226 10.6151
R2909 B.n375 B.n226 10.6151
R2910 B.n376 B.n375 10.6151
R2911 B.n377 B.n376 10.6151
R2912 B.n377 B.n224 10.6151
R2913 B.n381 B.n224 10.6151
R2914 B.n382 B.n381 10.6151
R2915 B.n383 B.n382 10.6151
R2916 B.n383 B.n222 10.6151
R2917 B.n387 B.n222 10.6151
R2918 B.n388 B.n387 10.6151
R2919 B.n389 B.n388 10.6151
R2920 B.n389 B.n220 10.6151
R2921 B.n393 B.n220 10.6151
R2922 B.n394 B.n393 10.6151
R2923 B.n395 B.n394 10.6151
R2924 B.n395 B.n218 10.6151
R2925 B.n399 B.n218 10.6151
R2926 B.n400 B.n399 10.6151
R2927 B.n401 B.n400 10.6151
R2928 B.n401 B.n216 10.6151
R2929 B.n405 B.n216 10.6151
R2930 B.n406 B.n405 10.6151
R2931 B.n407 B.n406 10.6151
R2932 B.n407 B.n214 10.6151
R2933 B.n411 B.n214 10.6151
R2934 B.n412 B.n411 10.6151
R2935 B.n413 B.n412 10.6151
R2936 B.n413 B.n212 10.6151
R2937 B.n417 B.n212 10.6151
R2938 B.n418 B.n417 10.6151
R2939 B.n419 B.n418 10.6151
R2940 B.n419 B.n210 10.6151
R2941 B.n423 B.n210 10.6151
R2942 B.n424 B.n423 10.6151
R2943 B.n425 B.n424 10.6151
R2944 B.n425 B.n208 10.6151
R2945 B.n429 B.n208 10.6151
R2946 B.n430 B.n429 10.6151
R2947 B.n431 B.n430 10.6151
R2948 B.n431 B.n206 10.6151
R2949 B.n435 B.n206 10.6151
R2950 B.n436 B.n435 10.6151
R2951 B.n437 B.n436 10.6151
R2952 B.n437 B.n204 10.6151
R2953 B.n441 B.n204 10.6151
R2954 B.n442 B.n441 10.6151
R2955 B.n446 B.n442 10.6151
R2956 B.n450 B.n202 10.6151
R2957 B.n451 B.n450 10.6151
R2958 B.n452 B.n451 10.6151
R2959 B.n452 B.n200 10.6151
R2960 B.n456 B.n200 10.6151
R2961 B.n457 B.n456 10.6151
R2962 B.n458 B.n457 10.6151
R2963 B.n458 B.n198 10.6151
R2964 B.n462 B.n198 10.6151
R2965 B.n465 B.n464 10.6151
R2966 B.n465 B.n194 10.6151
R2967 B.n469 B.n194 10.6151
R2968 B.n470 B.n469 10.6151
R2969 B.n471 B.n470 10.6151
R2970 B.n471 B.n192 10.6151
R2971 B.n475 B.n192 10.6151
R2972 B.n476 B.n475 10.6151
R2973 B.n477 B.n476 10.6151
R2974 B.n477 B.n190 10.6151
R2975 B.n481 B.n190 10.6151
R2976 B.n482 B.n481 10.6151
R2977 B.n483 B.n482 10.6151
R2978 B.n483 B.n188 10.6151
R2979 B.n487 B.n188 10.6151
R2980 B.n488 B.n487 10.6151
R2981 B.n489 B.n488 10.6151
R2982 B.n489 B.n186 10.6151
R2983 B.n493 B.n186 10.6151
R2984 B.n494 B.n493 10.6151
R2985 B.n495 B.n494 10.6151
R2986 B.n495 B.n184 10.6151
R2987 B.n499 B.n184 10.6151
R2988 B.n500 B.n499 10.6151
R2989 B.n501 B.n500 10.6151
R2990 B.n501 B.n182 10.6151
R2991 B.n505 B.n182 10.6151
R2992 B.n506 B.n505 10.6151
R2993 B.n507 B.n506 10.6151
R2994 B.n507 B.n180 10.6151
R2995 B.n511 B.n180 10.6151
R2996 B.n512 B.n511 10.6151
R2997 B.n513 B.n512 10.6151
R2998 B.n513 B.n178 10.6151
R2999 B.n517 B.n178 10.6151
R3000 B.n518 B.n517 10.6151
R3001 B.n519 B.n518 10.6151
R3002 B.n519 B.n176 10.6151
R3003 B.n523 B.n176 10.6151
R3004 B.n524 B.n523 10.6151
R3005 B.n525 B.n524 10.6151
R3006 B.n525 B.n174 10.6151
R3007 B.n529 B.n174 10.6151
R3008 B.n530 B.n529 10.6151
R3009 B.n531 B.n530 10.6151
R3010 B.n531 B.n172 10.6151
R3011 B.n535 B.n172 10.6151
R3012 B.n536 B.n535 10.6151
R3013 B.n537 B.n536 10.6151
R3014 B.n537 B.n170 10.6151
R3015 B.n541 B.n170 10.6151
R3016 B.n542 B.n541 10.6151
R3017 B.n543 B.n542 10.6151
R3018 B.n543 B.n168 10.6151
R3019 B.n547 B.n168 10.6151
R3020 B.n548 B.n547 10.6151
R3021 B.n549 B.n548 10.6151
R3022 B.n849 B.n848 9.36635
R3023 B.n831 B.n72 9.36635
R3024 B.n446 B.n445 9.36635
R3025 B.n464 B.n463 9.36635
R3026 B.n1033 B.n0 8.11757
R3027 B.n1033 B.n1 8.11757
R3028 B.n848 B.n847 1.24928
R3029 B.n834 B.n72 1.24928
R3030 B.n445 B.n202 1.24928
R3031 B.n463 B.n462 1.24928
C0 VN VDD2 13.2316f
C1 VTAIL VDD1 10.0591f
C2 w_n4810_n4496# B 13.0896f
C3 B VP 2.56394f
C4 VTAIL w_n4810_n4496# 5.52169f
C5 B VN 1.50782f
C6 VTAIL VP 13.6899f
C7 VDD1 w_n4810_n4496# 2.40061f
C8 B VDD2 2.20373f
C9 VTAIL VN 13.6758f
C10 VDD1 VP 13.6929f
C11 VDD1 VN 0.153808f
C12 VTAIL VDD2 10.1196f
C13 VDD1 VDD2 2.24969f
C14 w_n4810_n4496# VP 10.7584f
C15 w_n4810_n4496# VN 10.1313f
C16 VTAIL B 7.29754f
C17 VP VN 9.81173f
C18 w_n4810_n4496# VDD2 2.5535f
C19 VDD1 B 2.07907f
C20 VP VDD2 0.616939f
C21 VDD2 VSUBS 2.48053f
C22 VDD1 VSUBS 3.28563f
C23 VTAIL VSUBS 1.741621f
C24 VN VSUBS 8.142449f
C25 VP VSUBS 4.727406f
C26 B VSUBS 6.495272f
C27 w_n4810_n4496# VSUBS 0.264531p
C28 B.n0 VSUBS 0.006666f
C29 B.n1 VSUBS 0.006666f
C30 B.n2 VSUBS 0.009859f
C31 B.n3 VSUBS 0.007555f
C32 B.n4 VSUBS 0.007555f
C33 B.n5 VSUBS 0.007555f
C34 B.n6 VSUBS 0.007555f
C35 B.n7 VSUBS 0.007555f
C36 B.n8 VSUBS 0.007555f
C37 B.n9 VSUBS 0.007555f
C38 B.n10 VSUBS 0.007555f
C39 B.n11 VSUBS 0.007555f
C40 B.n12 VSUBS 0.007555f
C41 B.n13 VSUBS 0.007555f
C42 B.n14 VSUBS 0.007555f
C43 B.n15 VSUBS 0.007555f
C44 B.n16 VSUBS 0.007555f
C45 B.n17 VSUBS 0.007555f
C46 B.n18 VSUBS 0.007555f
C47 B.n19 VSUBS 0.007555f
C48 B.n20 VSUBS 0.007555f
C49 B.n21 VSUBS 0.007555f
C50 B.n22 VSUBS 0.007555f
C51 B.n23 VSUBS 0.007555f
C52 B.n24 VSUBS 0.007555f
C53 B.n25 VSUBS 0.007555f
C54 B.n26 VSUBS 0.007555f
C55 B.n27 VSUBS 0.007555f
C56 B.n28 VSUBS 0.007555f
C57 B.n29 VSUBS 0.007555f
C58 B.n30 VSUBS 0.007555f
C59 B.n31 VSUBS 0.007555f
C60 B.n32 VSUBS 0.007555f
C61 B.n33 VSUBS 0.007555f
C62 B.n34 VSUBS 0.018369f
C63 B.n35 VSUBS 0.007555f
C64 B.n36 VSUBS 0.007555f
C65 B.n37 VSUBS 0.007555f
C66 B.n38 VSUBS 0.007555f
C67 B.n39 VSUBS 0.007555f
C68 B.n40 VSUBS 0.007555f
C69 B.n41 VSUBS 0.007555f
C70 B.n42 VSUBS 0.007555f
C71 B.n43 VSUBS 0.007555f
C72 B.n44 VSUBS 0.007555f
C73 B.n45 VSUBS 0.007555f
C74 B.n46 VSUBS 0.007555f
C75 B.n47 VSUBS 0.007555f
C76 B.n48 VSUBS 0.007555f
C77 B.n49 VSUBS 0.007555f
C78 B.n50 VSUBS 0.007555f
C79 B.n51 VSUBS 0.007555f
C80 B.n52 VSUBS 0.007555f
C81 B.n53 VSUBS 0.007555f
C82 B.n54 VSUBS 0.007555f
C83 B.n55 VSUBS 0.007555f
C84 B.n56 VSUBS 0.007555f
C85 B.n57 VSUBS 0.007555f
C86 B.n58 VSUBS 0.007555f
C87 B.n59 VSUBS 0.007555f
C88 B.n60 VSUBS 0.007555f
C89 B.n61 VSUBS 0.007555f
C90 B.n62 VSUBS 0.007555f
C91 B.n63 VSUBS 0.007555f
C92 B.t4 VSUBS 0.369729f
C93 B.t5 VSUBS 0.416042f
C94 B.t3 VSUBS 3.03262f
C95 B.n64 VSUBS 0.660128f
C96 B.n65 VSUBS 0.353972f
C97 B.n66 VSUBS 0.007555f
C98 B.n67 VSUBS 0.007555f
C99 B.n68 VSUBS 0.007555f
C100 B.n69 VSUBS 0.007555f
C101 B.t7 VSUBS 0.369732f
C102 B.t8 VSUBS 0.416045f
C103 B.t6 VSUBS 3.03262f
C104 B.n70 VSUBS 0.660125f
C105 B.n71 VSUBS 0.353968f
C106 B.n72 VSUBS 0.017504f
C107 B.n73 VSUBS 0.007555f
C108 B.n74 VSUBS 0.007555f
C109 B.n75 VSUBS 0.007555f
C110 B.n76 VSUBS 0.007555f
C111 B.n77 VSUBS 0.007555f
C112 B.n78 VSUBS 0.007555f
C113 B.n79 VSUBS 0.007555f
C114 B.n80 VSUBS 0.007555f
C115 B.n81 VSUBS 0.007555f
C116 B.n82 VSUBS 0.007555f
C117 B.n83 VSUBS 0.007555f
C118 B.n84 VSUBS 0.007555f
C119 B.n85 VSUBS 0.007555f
C120 B.n86 VSUBS 0.007555f
C121 B.n87 VSUBS 0.007555f
C122 B.n88 VSUBS 0.007555f
C123 B.n89 VSUBS 0.007555f
C124 B.n90 VSUBS 0.007555f
C125 B.n91 VSUBS 0.007555f
C126 B.n92 VSUBS 0.007555f
C127 B.n93 VSUBS 0.007555f
C128 B.n94 VSUBS 0.007555f
C129 B.n95 VSUBS 0.007555f
C130 B.n96 VSUBS 0.007555f
C131 B.n97 VSUBS 0.007555f
C132 B.n98 VSUBS 0.007555f
C133 B.n99 VSUBS 0.007555f
C134 B.n100 VSUBS 0.007555f
C135 B.n101 VSUBS 0.018369f
C136 B.n102 VSUBS 0.007555f
C137 B.n103 VSUBS 0.007555f
C138 B.n104 VSUBS 0.007555f
C139 B.n105 VSUBS 0.007555f
C140 B.n106 VSUBS 0.007555f
C141 B.n107 VSUBS 0.007555f
C142 B.n108 VSUBS 0.007555f
C143 B.n109 VSUBS 0.007555f
C144 B.n110 VSUBS 0.007555f
C145 B.n111 VSUBS 0.007555f
C146 B.n112 VSUBS 0.007555f
C147 B.n113 VSUBS 0.007555f
C148 B.n114 VSUBS 0.007555f
C149 B.n115 VSUBS 0.007555f
C150 B.n116 VSUBS 0.007555f
C151 B.n117 VSUBS 0.007555f
C152 B.n118 VSUBS 0.007555f
C153 B.n119 VSUBS 0.007555f
C154 B.n120 VSUBS 0.007555f
C155 B.n121 VSUBS 0.007555f
C156 B.n122 VSUBS 0.007555f
C157 B.n123 VSUBS 0.007555f
C158 B.n124 VSUBS 0.007555f
C159 B.n125 VSUBS 0.007555f
C160 B.n126 VSUBS 0.007555f
C161 B.n127 VSUBS 0.007555f
C162 B.n128 VSUBS 0.007555f
C163 B.n129 VSUBS 0.007555f
C164 B.n130 VSUBS 0.007555f
C165 B.n131 VSUBS 0.007555f
C166 B.n132 VSUBS 0.007555f
C167 B.n133 VSUBS 0.007555f
C168 B.n134 VSUBS 0.007555f
C169 B.n135 VSUBS 0.007555f
C170 B.n136 VSUBS 0.007555f
C171 B.n137 VSUBS 0.007555f
C172 B.n138 VSUBS 0.007555f
C173 B.n139 VSUBS 0.007555f
C174 B.n140 VSUBS 0.007555f
C175 B.n141 VSUBS 0.007555f
C176 B.n142 VSUBS 0.007555f
C177 B.n143 VSUBS 0.007555f
C178 B.n144 VSUBS 0.007555f
C179 B.n145 VSUBS 0.007555f
C180 B.n146 VSUBS 0.007555f
C181 B.n147 VSUBS 0.007555f
C182 B.n148 VSUBS 0.007555f
C183 B.n149 VSUBS 0.007555f
C184 B.n150 VSUBS 0.007555f
C185 B.n151 VSUBS 0.007555f
C186 B.n152 VSUBS 0.007555f
C187 B.n153 VSUBS 0.007555f
C188 B.n154 VSUBS 0.007555f
C189 B.n155 VSUBS 0.007555f
C190 B.n156 VSUBS 0.007555f
C191 B.n157 VSUBS 0.007555f
C192 B.n158 VSUBS 0.007555f
C193 B.n159 VSUBS 0.007555f
C194 B.n160 VSUBS 0.007555f
C195 B.n161 VSUBS 0.007555f
C196 B.n162 VSUBS 0.007555f
C197 B.n163 VSUBS 0.007555f
C198 B.n164 VSUBS 0.007555f
C199 B.n165 VSUBS 0.007555f
C200 B.n166 VSUBS 0.018283f
C201 B.n167 VSUBS 0.007555f
C202 B.n168 VSUBS 0.007555f
C203 B.n169 VSUBS 0.007555f
C204 B.n170 VSUBS 0.007555f
C205 B.n171 VSUBS 0.007555f
C206 B.n172 VSUBS 0.007555f
C207 B.n173 VSUBS 0.007555f
C208 B.n174 VSUBS 0.007555f
C209 B.n175 VSUBS 0.007555f
C210 B.n176 VSUBS 0.007555f
C211 B.n177 VSUBS 0.007555f
C212 B.n178 VSUBS 0.007555f
C213 B.n179 VSUBS 0.007555f
C214 B.n180 VSUBS 0.007555f
C215 B.n181 VSUBS 0.007555f
C216 B.n182 VSUBS 0.007555f
C217 B.n183 VSUBS 0.007555f
C218 B.n184 VSUBS 0.007555f
C219 B.n185 VSUBS 0.007555f
C220 B.n186 VSUBS 0.007555f
C221 B.n187 VSUBS 0.007555f
C222 B.n188 VSUBS 0.007555f
C223 B.n189 VSUBS 0.007555f
C224 B.n190 VSUBS 0.007555f
C225 B.n191 VSUBS 0.007555f
C226 B.n192 VSUBS 0.007555f
C227 B.n193 VSUBS 0.007555f
C228 B.n194 VSUBS 0.007555f
C229 B.n195 VSUBS 0.007555f
C230 B.t2 VSUBS 0.369732f
C231 B.t1 VSUBS 0.416045f
C232 B.t0 VSUBS 3.03262f
C233 B.n196 VSUBS 0.660125f
C234 B.n197 VSUBS 0.353968f
C235 B.n198 VSUBS 0.007555f
C236 B.n199 VSUBS 0.007555f
C237 B.n200 VSUBS 0.007555f
C238 B.n201 VSUBS 0.007555f
C239 B.n202 VSUBS 0.004222f
C240 B.n203 VSUBS 0.007555f
C241 B.n204 VSUBS 0.007555f
C242 B.n205 VSUBS 0.007555f
C243 B.n206 VSUBS 0.007555f
C244 B.n207 VSUBS 0.007555f
C245 B.n208 VSUBS 0.007555f
C246 B.n209 VSUBS 0.007555f
C247 B.n210 VSUBS 0.007555f
C248 B.n211 VSUBS 0.007555f
C249 B.n212 VSUBS 0.007555f
C250 B.n213 VSUBS 0.007555f
C251 B.n214 VSUBS 0.007555f
C252 B.n215 VSUBS 0.007555f
C253 B.n216 VSUBS 0.007555f
C254 B.n217 VSUBS 0.007555f
C255 B.n218 VSUBS 0.007555f
C256 B.n219 VSUBS 0.007555f
C257 B.n220 VSUBS 0.007555f
C258 B.n221 VSUBS 0.007555f
C259 B.n222 VSUBS 0.007555f
C260 B.n223 VSUBS 0.007555f
C261 B.n224 VSUBS 0.007555f
C262 B.n225 VSUBS 0.007555f
C263 B.n226 VSUBS 0.007555f
C264 B.n227 VSUBS 0.007555f
C265 B.n228 VSUBS 0.007555f
C266 B.n229 VSUBS 0.007555f
C267 B.n230 VSUBS 0.007555f
C268 B.n231 VSUBS 0.018369f
C269 B.n232 VSUBS 0.007555f
C270 B.n233 VSUBS 0.007555f
C271 B.n234 VSUBS 0.007555f
C272 B.n235 VSUBS 0.007555f
C273 B.n236 VSUBS 0.007555f
C274 B.n237 VSUBS 0.007555f
C275 B.n238 VSUBS 0.007555f
C276 B.n239 VSUBS 0.007555f
C277 B.n240 VSUBS 0.007555f
C278 B.n241 VSUBS 0.007555f
C279 B.n242 VSUBS 0.007555f
C280 B.n243 VSUBS 0.007555f
C281 B.n244 VSUBS 0.007555f
C282 B.n245 VSUBS 0.007555f
C283 B.n246 VSUBS 0.007555f
C284 B.n247 VSUBS 0.007555f
C285 B.n248 VSUBS 0.007555f
C286 B.n249 VSUBS 0.007555f
C287 B.n250 VSUBS 0.007555f
C288 B.n251 VSUBS 0.007555f
C289 B.n252 VSUBS 0.007555f
C290 B.n253 VSUBS 0.007555f
C291 B.n254 VSUBS 0.007555f
C292 B.n255 VSUBS 0.007555f
C293 B.n256 VSUBS 0.007555f
C294 B.n257 VSUBS 0.007555f
C295 B.n258 VSUBS 0.007555f
C296 B.n259 VSUBS 0.007555f
C297 B.n260 VSUBS 0.007555f
C298 B.n261 VSUBS 0.007555f
C299 B.n262 VSUBS 0.007555f
C300 B.n263 VSUBS 0.007555f
C301 B.n264 VSUBS 0.007555f
C302 B.n265 VSUBS 0.007555f
C303 B.n266 VSUBS 0.007555f
C304 B.n267 VSUBS 0.007555f
C305 B.n268 VSUBS 0.007555f
C306 B.n269 VSUBS 0.007555f
C307 B.n270 VSUBS 0.007555f
C308 B.n271 VSUBS 0.007555f
C309 B.n272 VSUBS 0.007555f
C310 B.n273 VSUBS 0.007555f
C311 B.n274 VSUBS 0.007555f
C312 B.n275 VSUBS 0.007555f
C313 B.n276 VSUBS 0.007555f
C314 B.n277 VSUBS 0.007555f
C315 B.n278 VSUBS 0.007555f
C316 B.n279 VSUBS 0.007555f
C317 B.n280 VSUBS 0.007555f
C318 B.n281 VSUBS 0.007555f
C319 B.n282 VSUBS 0.007555f
C320 B.n283 VSUBS 0.007555f
C321 B.n284 VSUBS 0.007555f
C322 B.n285 VSUBS 0.007555f
C323 B.n286 VSUBS 0.007555f
C324 B.n287 VSUBS 0.007555f
C325 B.n288 VSUBS 0.007555f
C326 B.n289 VSUBS 0.007555f
C327 B.n290 VSUBS 0.007555f
C328 B.n291 VSUBS 0.007555f
C329 B.n292 VSUBS 0.007555f
C330 B.n293 VSUBS 0.007555f
C331 B.n294 VSUBS 0.007555f
C332 B.n295 VSUBS 0.007555f
C333 B.n296 VSUBS 0.007555f
C334 B.n297 VSUBS 0.007555f
C335 B.n298 VSUBS 0.007555f
C336 B.n299 VSUBS 0.007555f
C337 B.n300 VSUBS 0.007555f
C338 B.n301 VSUBS 0.007555f
C339 B.n302 VSUBS 0.007555f
C340 B.n303 VSUBS 0.007555f
C341 B.n304 VSUBS 0.007555f
C342 B.n305 VSUBS 0.007555f
C343 B.n306 VSUBS 0.007555f
C344 B.n307 VSUBS 0.007555f
C345 B.n308 VSUBS 0.007555f
C346 B.n309 VSUBS 0.007555f
C347 B.n310 VSUBS 0.007555f
C348 B.n311 VSUBS 0.007555f
C349 B.n312 VSUBS 0.007555f
C350 B.n313 VSUBS 0.007555f
C351 B.n314 VSUBS 0.007555f
C352 B.n315 VSUBS 0.007555f
C353 B.n316 VSUBS 0.007555f
C354 B.n317 VSUBS 0.007555f
C355 B.n318 VSUBS 0.007555f
C356 B.n319 VSUBS 0.007555f
C357 B.n320 VSUBS 0.007555f
C358 B.n321 VSUBS 0.007555f
C359 B.n322 VSUBS 0.007555f
C360 B.n323 VSUBS 0.007555f
C361 B.n324 VSUBS 0.007555f
C362 B.n325 VSUBS 0.007555f
C363 B.n326 VSUBS 0.007555f
C364 B.n327 VSUBS 0.007555f
C365 B.n328 VSUBS 0.007555f
C366 B.n329 VSUBS 0.007555f
C367 B.n330 VSUBS 0.007555f
C368 B.n331 VSUBS 0.007555f
C369 B.n332 VSUBS 0.007555f
C370 B.n333 VSUBS 0.007555f
C371 B.n334 VSUBS 0.007555f
C372 B.n335 VSUBS 0.007555f
C373 B.n336 VSUBS 0.007555f
C374 B.n337 VSUBS 0.007555f
C375 B.n338 VSUBS 0.007555f
C376 B.n339 VSUBS 0.007555f
C377 B.n340 VSUBS 0.007555f
C378 B.n341 VSUBS 0.007555f
C379 B.n342 VSUBS 0.007555f
C380 B.n343 VSUBS 0.007555f
C381 B.n344 VSUBS 0.007555f
C382 B.n345 VSUBS 0.007555f
C383 B.n346 VSUBS 0.007555f
C384 B.n347 VSUBS 0.007555f
C385 B.n348 VSUBS 0.007555f
C386 B.n349 VSUBS 0.007555f
C387 B.n350 VSUBS 0.007555f
C388 B.n351 VSUBS 0.007555f
C389 B.n352 VSUBS 0.007555f
C390 B.n353 VSUBS 0.007555f
C391 B.n354 VSUBS 0.007555f
C392 B.n355 VSUBS 0.007555f
C393 B.n356 VSUBS 0.017406f
C394 B.n357 VSUBS 0.017406f
C395 B.n358 VSUBS 0.018369f
C396 B.n359 VSUBS 0.007555f
C397 B.n360 VSUBS 0.007555f
C398 B.n361 VSUBS 0.007555f
C399 B.n362 VSUBS 0.007555f
C400 B.n363 VSUBS 0.007555f
C401 B.n364 VSUBS 0.007555f
C402 B.n365 VSUBS 0.007555f
C403 B.n366 VSUBS 0.007555f
C404 B.n367 VSUBS 0.007555f
C405 B.n368 VSUBS 0.007555f
C406 B.n369 VSUBS 0.007555f
C407 B.n370 VSUBS 0.007555f
C408 B.n371 VSUBS 0.007555f
C409 B.n372 VSUBS 0.007555f
C410 B.n373 VSUBS 0.007555f
C411 B.n374 VSUBS 0.007555f
C412 B.n375 VSUBS 0.007555f
C413 B.n376 VSUBS 0.007555f
C414 B.n377 VSUBS 0.007555f
C415 B.n378 VSUBS 0.007555f
C416 B.n379 VSUBS 0.007555f
C417 B.n380 VSUBS 0.007555f
C418 B.n381 VSUBS 0.007555f
C419 B.n382 VSUBS 0.007555f
C420 B.n383 VSUBS 0.007555f
C421 B.n384 VSUBS 0.007555f
C422 B.n385 VSUBS 0.007555f
C423 B.n386 VSUBS 0.007555f
C424 B.n387 VSUBS 0.007555f
C425 B.n388 VSUBS 0.007555f
C426 B.n389 VSUBS 0.007555f
C427 B.n390 VSUBS 0.007555f
C428 B.n391 VSUBS 0.007555f
C429 B.n392 VSUBS 0.007555f
C430 B.n393 VSUBS 0.007555f
C431 B.n394 VSUBS 0.007555f
C432 B.n395 VSUBS 0.007555f
C433 B.n396 VSUBS 0.007555f
C434 B.n397 VSUBS 0.007555f
C435 B.n398 VSUBS 0.007555f
C436 B.n399 VSUBS 0.007555f
C437 B.n400 VSUBS 0.007555f
C438 B.n401 VSUBS 0.007555f
C439 B.n402 VSUBS 0.007555f
C440 B.n403 VSUBS 0.007555f
C441 B.n404 VSUBS 0.007555f
C442 B.n405 VSUBS 0.007555f
C443 B.n406 VSUBS 0.007555f
C444 B.n407 VSUBS 0.007555f
C445 B.n408 VSUBS 0.007555f
C446 B.n409 VSUBS 0.007555f
C447 B.n410 VSUBS 0.007555f
C448 B.n411 VSUBS 0.007555f
C449 B.n412 VSUBS 0.007555f
C450 B.n413 VSUBS 0.007555f
C451 B.n414 VSUBS 0.007555f
C452 B.n415 VSUBS 0.007555f
C453 B.n416 VSUBS 0.007555f
C454 B.n417 VSUBS 0.007555f
C455 B.n418 VSUBS 0.007555f
C456 B.n419 VSUBS 0.007555f
C457 B.n420 VSUBS 0.007555f
C458 B.n421 VSUBS 0.007555f
C459 B.n422 VSUBS 0.007555f
C460 B.n423 VSUBS 0.007555f
C461 B.n424 VSUBS 0.007555f
C462 B.n425 VSUBS 0.007555f
C463 B.n426 VSUBS 0.007555f
C464 B.n427 VSUBS 0.007555f
C465 B.n428 VSUBS 0.007555f
C466 B.n429 VSUBS 0.007555f
C467 B.n430 VSUBS 0.007555f
C468 B.n431 VSUBS 0.007555f
C469 B.n432 VSUBS 0.007555f
C470 B.n433 VSUBS 0.007555f
C471 B.n434 VSUBS 0.007555f
C472 B.n435 VSUBS 0.007555f
C473 B.n436 VSUBS 0.007555f
C474 B.n437 VSUBS 0.007555f
C475 B.n438 VSUBS 0.007555f
C476 B.n439 VSUBS 0.007555f
C477 B.n440 VSUBS 0.007555f
C478 B.n441 VSUBS 0.007555f
C479 B.n442 VSUBS 0.007555f
C480 B.t11 VSUBS 0.369729f
C481 B.t10 VSUBS 0.416042f
C482 B.t9 VSUBS 3.03262f
C483 B.n443 VSUBS 0.660128f
C484 B.n444 VSUBS 0.353972f
C485 B.n445 VSUBS 0.017504f
C486 B.n446 VSUBS 0.007111f
C487 B.n447 VSUBS 0.007555f
C488 B.n448 VSUBS 0.007555f
C489 B.n449 VSUBS 0.007555f
C490 B.n450 VSUBS 0.007555f
C491 B.n451 VSUBS 0.007555f
C492 B.n452 VSUBS 0.007555f
C493 B.n453 VSUBS 0.007555f
C494 B.n454 VSUBS 0.007555f
C495 B.n455 VSUBS 0.007555f
C496 B.n456 VSUBS 0.007555f
C497 B.n457 VSUBS 0.007555f
C498 B.n458 VSUBS 0.007555f
C499 B.n459 VSUBS 0.007555f
C500 B.n460 VSUBS 0.007555f
C501 B.n461 VSUBS 0.007555f
C502 B.n462 VSUBS 0.004222f
C503 B.n463 VSUBS 0.017504f
C504 B.n464 VSUBS 0.007111f
C505 B.n465 VSUBS 0.007555f
C506 B.n466 VSUBS 0.007555f
C507 B.n467 VSUBS 0.007555f
C508 B.n468 VSUBS 0.007555f
C509 B.n469 VSUBS 0.007555f
C510 B.n470 VSUBS 0.007555f
C511 B.n471 VSUBS 0.007555f
C512 B.n472 VSUBS 0.007555f
C513 B.n473 VSUBS 0.007555f
C514 B.n474 VSUBS 0.007555f
C515 B.n475 VSUBS 0.007555f
C516 B.n476 VSUBS 0.007555f
C517 B.n477 VSUBS 0.007555f
C518 B.n478 VSUBS 0.007555f
C519 B.n479 VSUBS 0.007555f
C520 B.n480 VSUBS 0.007555f
C521 B.n481 VSUBS 0.007555f
C522 B.n482 VSUBS 0.007555f
C523 B.n483 VSUBS 0.007555f
C524 B.n484 VSUBS 0.007555f
C525 B.n485 VSUBS 0.007555f
C526 B.n486 VSUBS 0.007555f
C527 B.n487 VSUBS 0.007555f
C528 B.n488 VSUBS 0.007555f
C529 B.n489 VSUBS 0.007555f
C530 B.n490 VSUBS 0.007555f
C531 B.n491 VSUBS 0.007555f
C532 B.n492 VSUBS 0.007555f
C533 B.n493 VSUBS 0.007555f
C534 B.n494 VSUBS 0.007555f
C535 B.n495 VSUBS 0.007555f
C536 B.n496 VSUBS 0.007555f
C537 B.n497 VSUBS 0.007555f
C538 B.n498 VSUBS 0.007555f
C539 B.n499 VSUBS 0.007555f
C540 B.n500 VSUBS 0.007555f
C541 B.n501 VSUBS 0.007555f
C542 B.n502 VSUBS 0.007555f
C543 B.n503 VSUBS 0.007555f
C544 B.n504 VSUBS 0.007555f
C545 B.n505 VSUBS 0.007555f
C546 B.n506 VSUBS 0.007555f
C547 B.n507 VSUBS 0.007555f
C548 B.n508 VSUBS 0.007555f
C549 B.n509 VSUBS 0.007555f
C550 B.n510 VSUBS 0.007555f
C551 B.n511 VSUBS 0.007555f
C552 B.n512 VSUBS 0.007555f
C553 B.n513 VSUBS 0.007555f
C554 B.n514 VSUBS 0.007555f
C555 B.n515 VSUBS 0.007555f
C556 B.n516 VSUBS 0.007555f
C557 B.n517 VSUBS 0.007555f
C558 B.n518 VSUBS 0.007555f
C559 B.n519 VSUBS 0.007555f
C560 B.n520 VSUBS 0.007555f
C561 B.n521 VSUBS 0.007555f
C562 B.n522 VSUBS 0.007555f
C563 B.n523 VSUBS 0.007555f
C564 B.n524 VSUBS 0.007555f
C565 B.n525 VSUBS 0.007555f
C566 B.n526 VSUBS 0.007555f
C567 B.n527 VSUBS 0.007555f
C568 B.n528 VSUBS 0.007555f
C569 B.n529 VSUBS 0.007555f
C570 B.n530 VSUBS 0.007555f
C571 B.n531 VSUBS 0.007555f
C572 B.n532 VSUBS 0.007555f
C573 B.n533 VSUBS 0.007555f
C574 B.n534 VSUBS 0.007555f
C575 B.n535 VSUBS 0.007555f
C576 B.n536 VSUBS 0.007555f
C577 B.n537 VSUBS 0.007555f
C578 B.n538 VSUBS 0.007555f
C579 B.n539 VSUBS 0.007555f
C580 B.n540 VSUBS 0.007555f
C581 B.n541 VSUBS 0.007555f
C582 B.n542 VSUBS 0.007555f
C583 B.n543 VSUBS 0.007555f
C584 B.n544 VSUBS 0.007555f
C585 B.n545 VSUBS 0.007555f
C586 B.n546 VSUBS 0.007555f
C587 B.n547 VSUBS 0.007555f
C588 B.n548 VSUBS 0.007555f
C589 B.n549 VSUBS 0.017492f
C590 B.n550 VSUBS 0.018369f
C591 B.n551 VSUBS 0.017406f
C592 B.n552 VSUBS 0.007555f
C593 B.n553 VSUBS 0.007555f
C594 B.n554 VSUBS 0.007555f
C595 B.n555 VSUBS 0.007555f
C596 B.n556 VSUBS 0.007555f
C597 B.n557 VSUBS 0.007555f
C598 B.n558 VSUBS 0.007555f
C599 B.n559 VSUBS 0.007555f
C600 B.n560 VSUBS 0.007555f
C601 B.n561 VSUBS 0.007555f
C602 B.n562 VSUBS 0.007555f
C603 B.n563 VSUBS 0.007555f
C604 B.n564 VSUBS 0.007555f
C605 B.n565 VSUBS 0.007555f
C606 B.n566 VSUBS 0.007555f
C607 B.n567 VSUBS 0.007555f
C608 B.n568 VSUBS 0.007555f
C609 B.n569 VSUBS 0.007555f
C610 B.n570 VSUBS 0.007555f
C611 B.n571 VSUBS 0.007555f
C612 B.n572 VSUBS 0.007555f
C613 B.n573 VSUBS 0.007555f
C614 B.n574 VSUBS 0.007555f
C615 B.n575 VSUBS 0.007555f
C616 B.n576 VSUBS 0.007555f
C617 B.n577 VSUBS 0.007555f
C618 B.n578 VSUBS 0.007555f
C619 B.n579 VSUBS 0.007555f
C620 B.n580 VSUBS 0.007555f
C621 B.n581 VSUBS 0.007555f
C622 B.n582 VSUBS 0.007555f
C623 B.n583 VSUBS 0.007555f
C624 B.n584 VSUBS 0.007555f
C625 B.n585 VSUBS 0.007555f
C626 B.n586 VSUBS 0.007555f
C627 B.n587 VSUBS 0.007555f
C628 B.n588 VSUBS 0.007555f
C629 B.n589 VSUBS 0.007555f
C630 B.n590 VSUBS 0.007555f
C631 B.n591 VSUBS 0.007555f
C632 B.n592 VSUBS 0.007555f
C633 B.n593 VSUBS 0.007555f
C634 B.n594 VSUBS 0.007555f
C635 B.n595 VSUBS 0.007555f
C636 B.n596 VSUBS 0.007555f
C637 B.n597 VSUBS 0.007555f
C638 B.n598 VSUBS 0.007555f
C639 B.n599 VSUBS 0.007555f
C640 B.n600 VSUBS 0.007555f
C641 B.n601 VSUBS 0.007555f
C642 B.n602 VSUBS 0.007555f
C643 B.n603 VSUBS 0.007555f
C644 B.n604 VSUBS 0.007555f
C645 B.n605 VSUBS 0.007555f
C646 B.n606 VSUBS 0.007555f
C647 B.n607 VSUBS 0.007555f
C648 B.n608 VSUBS 0.007555f
C649 B.n609 VSUBS 0.007555f
C650 B.n610 VSUBS 0.007555f
C651 B.n611 VSUBS 0.007555f
C652 B.n612 VSUBS 0.007555f
C653 B.n613 VSUBS 0.007555f
C654 B.n614 VSUBS 0.007555f
C655 B.n615 VSUBS 0.007555f
C656 B.n616 VSUBS 0.007555f
C657 B.n617 VSUBS 0.007555f
C658 B.n618 VSUBS 0.007555f
C659 B.n619 VSUBS 0.007555f
C660 B.n620 VSUBS 0.007555f
C661 B.n621 VSUBS 0.007555f
C662 B.n622 VSUBS 0.007555f
C663 B.n623 VSUBS 0.007555f
C664 B.n624 VSUBS 0.007555f
C665 B.n625 VSUBS 0.007555f
C666 B.n626 VSUBS 0.007555f
C667 B.n627 VSUBS 0.007555f
C668 B.n628 VSUBS 0.007555f
C669 B.n629 VSUBS 0.007555f
C670 B.n630 VSUBS 0.007555f
C671 B.n631 VSUBS 0.007555f
C672 B.n632 VSUBS 0.007555f
C673 B.n633 VSUBS 0.007555f
C674 B.n634 VSUBS 0.007555f
C675 B.n635 VSUBS 0.007555f
C676 B.n636 VSUBS 0.007555f
C677 B.n637 VSUBS 0.007555f
C678 B.n638 VSUBS 0.007555f
C679 B.n639 VSUBS 0.007555f
C680 B.n640 VSUBS 0.007555f
C681 B.n641 VSUBS 0.007555f
C682 B.n642 VSUBS 0.007555f
C683 B.n643 VSUBS 0.007555f
C684 B.n644 VSUBS 0.007555f
C685 B.n645 VSUBS 0.007555f
C686 B.n646 VSUBS 0.007555f
C687 B.n647 VSUBS 0.007555f
C688 B.n648 VSUBS 0.007555f
C689 B.n649 VSUBS 0.007555f
C690 B.n650 VSUBS 0.007555f
C691 B.n651 VSUBS 0.007555f
C692 B.n652 VSUBS 0.007555f
C693 B.n653 VSUBS 0.007555f
C694 B.n654 VSUBS 0.007555f
C695 B.n655 VSUBS 0.007555f
C696 B.n656 VSUBS 0.007555f
C697 B.n657 VSUBS 0.007555f
C698 B.n658 VSUBS 0.007555f
C699 B.n659 VSUBS 0.007555f
C700 B.n660 VSUBS 0.007555f
C701 B.n661 VSUBS 0.007555f
C702 B.n662 VSUBS 0.007555f
C703 B.n663 VSUBS 0.007555f
C704 B.n664 VSUBS 0.007555f
C705 B.n665 VSUBS 0.007555f
C706 B.n666 VSUBS 0.007555f
C707 B.n667 VSUBS 0.007555f
C708 B.n668 VSUBS 0.007555f
C709 B.n669 VSUBS 0.007555f
C710 B.n670 VSUBS 0.007555f
C711 B.n671 VSUBS 0.007555f
C712 B.n672 VSUBS 0.007555f
C713 B.n673 VSUBS 0.007555f
C714 B.n674 VSUBS 0.007555f
C715 B.n675 VSUBS 0.007555f
C716 B.n676 VSUBS 0.007555f
C717 B.n677 VSUBS 0.007555f
C718 B.n678 VSUBS 0.007555f
C719 B.n679 VSUBS 0.007555f
C720 B.n680 VSUBS 0.007555f
C721 B.n681 VSUBS 0.007555f
C722 B.n682 VSUBS 0.007555f
C723 B.n683 VSUBS 0.007555f
C724 B.n684 VSUBS 0.007555f
C725 B.n685 VSUBS 0.007555f
C726 B.n686 VSUBS 0.007555f
C727 B.n687 VSUBS 0.007555f
C728 B.n688 VSUBS 0.007555f
C729 B.n689 VSUBS 0.007555f
C730 B.n690 VSUBS 0.007555f
C731 B.n691 VSUBS 0.007555f
C732 B.n692 VSUBS 0.007555f
C733 B.n693 VSUBS 0.007555f
C734 B.n694 VSUBS 0.007555f
C735 B.n695 VSUBS 0.007555f
C736 B.n696 VSUBS 0.007555f
C737 B.n697 VSUBS 0.007555f
C738 B.n698 VSUBS 0.007555f
C739 B.n699 VSUBS 0.007555f
C740 B.n700 VSUBS 0.007555f
C741 B.n701 VSUBS 0.007555f
C742 B.n702 VSUBS 0.007555f
C743 B.n703 VSUBS 0.007555f
C744 B.n704 VSUBS 0.007555f
C745 B.n705 VSUBS 0.007555f
C746 B.n706 VSUBS 0.007555f
C747 B.n707 VSUBS 0.007555f
C748 B.n708 VSUBS 0.007555f
C749 B.n709 VSUBS 0.007555f
C750 B.n710 VSUBS 0.007555f
C751 B.n711 VSUBS 0.007555f
C752 B.n712 VSUBS 0.007555f
C753 B.n713 VSUBS 0.007555f
C754 B.n714 VSUBS 0.007555f
C755 B.n715 VSUBS 0.007555f
C756 B.n716 VSUBS 0.007555f
C757 B.n717 VSUBS 0.007555f
C758 B.n718 VSUBS 0.007555f
C759 B.n719 VSUBS 0.007555f
C760 B.n720 VSUBS 0.007555f
C761 B.n721 VSUBS 0.007555f
C762 B.n722 VSUBS 0.007555f
C763 B.n723 VSUBS 0.007555f
C764 B.n724 VSUBS 0.007555f
C765 B.n725 VSUBS 0.007555f
C766 B.n726 VSUBS 0.007555f
C767 B.n727 VSUBS 0.007555f
C768 B.n728 VSUBS 0.007555f
C769 B.n729 VSUBS 0.007555f
C770 B.n730 VSUBS 0.007555f
C771 B.n731 VSUBS 0.007555f
C772 B.n732 VSUBS 0.007555f
C773 B.n733 VSUBS 0.007555f
C774 B.n734 VSUBS 0.007555f
C775 B.n735 VSUBS 0.007555f
C776 B.n736 VSUBS 0.007555f
C777 B.n737 VSUBS 0.007555f
C778 B.n738 VSUBS 0.007555f
C779 B.n739 VSUBS 0.007555f
C780 B.n740 VSUBS 0.007555f
C781 B.n741 VSUBS 0.007555f
C782 B.n742 VSUBS 0.007555f
C783 B.n743 VSUBS 0.007555f
C784 B.n744 VSUBS 0.017406f
C785 B.n745 VSUBS 0.017406f
C786 B.n746 VSUBS 0.018369f
C787 B.n747 VSUBS 0.007555f
C788 B.n748 VSUBS 0.007555f
C789 B.n749 VSUBS 0.007555f
C790 B.n750 VSUBS 0.007555f
C791 B.n751 VSUBS 0.007555f
C792 B.n752 VSUBS 0.007555f
C793 B.n753 VSUBS 0.007555f
C794 B.n754 VSUBS 0.007555f
C795 B.n755 VSUBS 0.007555f
C796 B.n756 VSUBS 0.007555f
C797 B.n757 VSUBS 0.007555f
C798 B.n758 VSUBS 0.007555f
C799 B.n759 VSUBS 0.007555f
C800 B.n760 VSUBS 0.007555f
C801 B.n761 VSUBS 0.007555f
C802 B.n762 VSUBS 0.007555f
C803 B.n763 VSUBS 0.007555f
C804 B.n764 VSUBS 0.007555f
C805 B.n765 VSUBS 0.007555f
C806 B.n766 VSUBS 0.007555f
C807 B.n767 VSUBS 0.007555f
C808 B.n768 VSUBS 0.007555f
C809 B.n769 VSUBS 0.007555f
C810 B.n770 VSUBS 0.007555f
C811 B.n771 VSUBS 0.007555f
C812 B.n772 VSUBS 0.007555f
C813 B.n773 VSUBS 0.007555f
C814 B.n774 VSUBS 0.007555f
C815 B.n775 VSUBS 0.007555f
C816 B.n776 VSUBS 0.007555f
C817 B.n777 VSUBS 0.007555f
C818 B.n778 VSUBS 0.007555f
C819 B.n779 VSUBS 0.007555f
C820 B.n780 VSUBS 0.007555f
C821 B.n781 VSUBS 0.007555f
C822 B.n782 VSUBS 0.007555f
C823 B.n783 VSUBS 0.007555f
C824 B.n784 VSUBS 0.007555f
C825 B.n785 VSUBS 0.007555f
C826 B.n786 VSUBS 0.007555f
C827 B.n787 VSUBS 0.007555f
C828 B.n788 VSUBS 0.007555f
C829 B.n789 VSUBS 0.007555f
C830 B.n790 VSUBS 0.007555f
C831 B.n791 VSUBS 0.007555f
C832 B.n792 VSUBS 0.007555f
C833 B.n793 VSUBS 0.007555f
C834 B.n794 VSUBS 0.007555f
C835 B.n795 VSUBS 0.007555f
C836 B.n796 VSUBS 0.007555f
C837 B.n797 VSUBS 0.007555f
C838 B.n798 VSUBS 0.007555f
C839 B.n799 VSUBS 0.007555f
C840 B.n800 VSUBS 0.007555f
C841 B.n801 VSUBS 0.007555f
C842 B.n802 VSUBS 0.007555f
C843 B.n803 VSUBS 0.007555f
C844 B.n804 VSUBS 0.007555f
C845 B.n805 VSUBS 0.007555f
C846 B.n806 VSUBS 0.007555f
C847 B.n807 VSUBS 0.007555f
C848 B.n808 VSUBS 0.007555f
C849 B.n809 VSUBS 0.007555f
C850 B.n810 VSUBS 0.007555f
C851 B.n811 VSUBS 0.007555f
C852 B.n812 VSUBS 0.007555f
C853 B.n813 VSUBS 0.007555f
C854 B.n814 VSUBS 0.007555f
C855 B.n815 VSUBS 0.007555f
C856 B.n816 VSUBS 0.007555f
C857 B.n817 VSUBS 0.007555f
C858 B.n818 VSUBS 0.007555f
C859 B.n819 VSUBS 0.007555f
C860 B.n820 VSUBS 0.007555f
C861 B.n821 VSUBS 0.007555f
C862 B.n822 VSUBS 0.007555f
C863 B.n823 VSUBS 0.007555f
C864 B.n824 VSUBS 0.007555f
C865 B.n825 VSUBS 0.007555f
C866 B.n826 VSUBS 0.007555f
C867 B.n827 VSUBS 0.007555f
C868 B.n828 VSUBS 0.007555f
C869 B.n829 VSUBS 0.007555f
C870 B.n830 VSUBS 0.007555f
C871 B.n831 VSUBS 0.007111f
C872 B.n832 VSUBS 0.007555f
C873 B.n833 VSUBS 0.007555f
C874 B.n834 VSUBS 0.004222f
C875 B.n835 VSUBS 0.007555f
C876 B.n836 VSUBS 0.007555f
C877 B.n837 VSUBS 0.007555f
C878 B.n838 VSUBS 0.007555f
C879 B.n839 VSUBS 0.007555f
C880 B.n840 VSUBS 0.007555f
C881 B.n841 VSUBS 0.007555f
C882 B.n842 VSUBS 0.007555f
C883 B.n843 VSUBS 0.007555f
C884 B.n844 VSUBS 0.007555f
C885 B.n845 VSUBS 0.007555f
C886 B.n846 VSUBS 0.007555f
C887 B.n847 VSUBS 0.004222f
C888 B.n848 VSUBS 0.017504f
C889 B.n849 VSUBS 0.007111f
C890 B.n850 VSUBS 0.007555f
C891 B.n851 VSUBS 0.007555f
C892 B.n852 VSUBS 0.007555f
C893 B.n853 VSUBS 0.007555f
C894 B.n854 VSUBS 0.007555f
C895 B.n855 VSUBS 0.007555f
C896 B.n856 VSUBS 0.007555f
C897 B.n857 VSUBS 0.007555f
C898 B.n858 VSUBS 0.007555f
C899 B.n859 VSUBS 0.007555f
C900 B.n860 VSUBS 0.007555f
C901 B.n861 VSUBS 0.007555f
C902 B.n862 VSUBS 0.007555f
C903 B.n863 VSUBS 0.007555f
C904 B.n864 VSUBS 0.007555f
C905 B.n865 VSUBS 0.007555f
C906 B.n866 VSUBS 0.007555f
C907 B.n867 VSUBS 0.007555f
C908 B.n868 VSUBS 0.007555f
C909 B.n869 VSUBS 0.007555f
C910 B.n870 VSUBS 0.007555f
C911 B.n871 VSUBS 0.007555f
C912 B.n872 VSUBS 0.007555f
C913 B.n873 VSUBS 0.007555f
C914 B.n874 VSUBS 0.007555f
C915 B.n875 VSUBS 0.007555f
C916 B.n876 VSUBS 0.007555f
C917 B.n877 VSUBS 0.007555f
C918 B.n878 VSUBS 0.007555f
C919 B.n879 VSUBS 0.007555f
C920 B.n880 VSUBS 0.007555f
C921 B.n881 VSUBS 0.007555f
C922 B.n882 VSUBS 0.007555f
C923 B.n883 VSUBS 0.007555f
C924 B.n884 VSUBS 0.007555f
C925 B.n885 VSUBS 0.007555f
C926 B.n886 VSUBS 0.007555f
C927 B.n887 VSUBS 0.007555f
C928 B.n888 VSUBS 0.007555f
C929 B.n889 VSUBS 0.007555f
C930 B.n890 VSUBS 0.007555f
C931 B.n891 VSUBS 0.007555f
C932 B.n892 VSUBS 0.007555f
C933 B.n893 VSUBS 0.007555f
C934 B.n894 VSUBS 0.007555f
C935 B.n895 VSUBS 0.007555f
C936 B.n896 VSUBS 0.007555f
C937 B.n897 VSUBS 0.007555f
C938 B.n898 VSUBS 0.007555f
C939 B.n899 VSUBS 0.007555f
C940 B.n900 VSUBS 0.007555f
C941 B.n901 VSUBS 0.007555f
C942 B.n902 VSUBS 0.007555f
C943 B.n903 VSUBS 0.007555f
C944 B.n904 VSUBS 0.007555f
C945 B.n905 VSUBS 0.007555f
C946 B.n906 VSUBS 0.007555f
C947 B.n907 VSUBS 0.007555f
C948 B.n908 VSUBS 0.007555f
C949 B.n909 VSUBS 0.007555f
C950 B.n910 VSUBS 0.007555f
C951 B.n911 VSUBS 0.007555f
C952 B.n912 VSUBS 0.007555f
C953 B.n913 VSUBS 0.007555f
C954 B.n914 VSUBS 0.007555f
C955 B.n915 VSUBS 0.007555f
C956 B.n916 VSUBS 0.007555f
C957 B.n917 VSUBS 0.007555f
C958 B.n918 VSUBS 0.007555f
C959 B.n919 VSUBS 0.007555f
C960 B.n920 VSUBS 0.007555f
C961 B.n921 VSUBS 0.007555f
C962 B.n922 VSUBS 0.007555f
C963 B.n923 VSUBS 0.007555f
C964 B.n924 VSUBS 0.007555f
C965 B.n925 VSUBS 0.007555f
C966 B.n926 VSUBS 0.007555f
C967 B.n927 VSUBS 0.007555f
C968 B.n928 VSUBS 0.007555f
C969 B.n929 VSUBS 0.007555f
C970 B.n930 VSUBS 0.007555f
C971 B.n931 VSUBS 0.007555f
C972 B.n932 VSUBS 0.007555f
C973 B.n933 VSUBS 0.007555f
C974 B.n934 VSUBS 0.007555f
C975 B.n935 VSUBS 0.018369f
C976 B.n936 VSUBS 0.017406f
C977 B.n937 VSUBS 0.017406f
C978 B.n938 VSUBS 0.007555f
C979 B.n939 VSUBS 0.007555f
C980 B.n940 VSUBS 0.007555f
C981 B.n941 VSUBS 0.007555f
C982 B.n942 VSUBS 0.007555f
C983 B.n943 VSUBS 0.007555f
C984 B.n944 VSUBS 0.007555f
C985 B.n945 VSUBS 0.007555f
C986 B.n946 VSUBS 0.007555f
C987 B.n947 VSUBS 0.007555f
C988 B.n948 VSUBS 0.007555f
C989 B.n949 VSUBS 0.007555f
C990 B.n950 VSUBS 0.007555f
C991 B.n951 VSUBS 0.007555f
C992 B.n952 VSUBS 0.007555f
C993 B.n953 VSUBS 0.007555f
C994 B.n954 VSUBS 0.007555f
C995 B.n955 VSUBS 0.007555f
C996 B.n956 VSUBS 0.007555f
C997 B.n957 VSUBS 0.007555f
C998 B.n958 VSUBS 0.007555f
C999 B.n959 VSUBS 0.007555f
C1000 B.n960 VSUBS 0.007555f
C1001 B.n961 VSUBS 0.007555f
C1002 B.n962 VSUBS 0.007555f
C1003 B.n963 VSUBS 0.007555f
C1004 B.n964 VSUBS 0.007555f
C1005 B.n965 VSUBS 0.007555f
C1006 B.n966 VSUBS 0.007555f
C1007 B.n967 VSUBS 0.007555f
C1008 B.n968 VSUBS 0.007555f
C1009 B.n969 VSUBS 0.007555f
C1010 B.n970 VSUBS 0.007555f
C1011 B.n971 VSUBS 0.007555f
C1012 B.n972 VSUBS 0.007555f
C1013 B.n973 VSUBS 0.007555f
C1014 B.n974 VSUBS 0.007555f
C1015 B.n975 VSUBS 0.007555f
C1016 B.n976 VSUBS 0.007555f
C1017 B.n977 VSUBS 0.007555f
C1018 B.n978 VSUBS 0.007555f
C1019 B.n979 VSUBS 0.007555f
C1020 B.n980 VSUBS 0.007555f
C1021 B.n981 VSUBS 0.007555f
C1022 B.n982 VSUBS 0.007555f
C1023 B.n983 VSUBS 0.007555f
C1024 B.n984 VSUBS 0.007555f
C1025 B.n985 VSUBS 0.007555f
C1026 B.n986 VSUBS 0.007555f
C1027 B.n987 VSUBS 0.007555f
C1028 B.n988 VSUBS 0.007555f
C1029 B.n989 VSUBS 0.007555f
C1030 B.n990 VSUBS 0.007555f
C1031 B.n991 VSUBS 0.007555f
C1032 B.n992 VSUBS 0.007555f
C1033 B.n993 VSUBS 0.007555f
C1034 B.n994 VSUBS 0.007555f
C1035 B.n995 VSUBS 0.007555f
C1036 B.n996 VSUBS 0.007555f
C1037 B.n997 VSUBS 0.007555f
C1038 B.n998 VSUBS 0.007555f
C1039 B.n999 VSUBS 0.007555f
C1040 B.n1000 VSUBS 0.007555f
C1041 B.n1001 VSUBS 0.007555f
C1042 B.n1002 VSUBS 0.007555f
C1043 B.n1003 VSUBS 0.007555f
C1044 B.n1004 VSUBS 0.007555f
C1045 B.n1005 VSUBS 0.007555f
C1046 B.n1006 VSUBS 0.007555f
C1047 B.n1007 VSUBS 0.007555f
C1048 B.n1008 VSUBS 0.007555f
C1049 B.n1009 VSUBS 0.007555f
C1050 B.n1010 VSUBS 0.007555f
C1051 B.n1011 VSUBS 0.007555f
C1052 B.n1012 VSUBS 0.007555f
C1053 B.n1013 VSUBS 0.007555f
C1054 B.n1014 VSUBS 0.007555f
C1055 B.n1015 VSUBS 0.007555f
C1056 B.n1016 VSUBS 0.007555f
C1057 B.n1017 VSUBS 0.007555f
C1058 B.n1018 VSUBS 0.007555f
C1059 B.n1019 VSUBS 0.007555f
C1060 B.n1020 VSUBS 0.007555f
C1061 B.n1021 VSUBS 0.007555f
C1062 B.n1022 VSUBS 0.007555f
C1063 B.n1023 VSUBS 0.007555f
C1064 B.n1024 VSUBS 0.007555f
C1065 B.n1025 VSUBS 0.007555f
C1066 B.n1026 VSUBS 0.007555f
C1067 B.n1027 VSUBS 0.007555f
C1068 B.n1028 VSUBS 0.007555f
C1069 B.n1029 VSUBS 0.007555f
C1070 B.n1030 VSUBS 0.007555f
C1071 B.n1031 VSUBS 0.009859f
C1072 B.n1032 VSUBS 0.010502f
C1073 B.n1033 VSUBS 0.020885f
C1074 VDD1.t2 VSUBS 0.436739f
C1075 VDD1.t3 VSUBS 0.436739f
C1076 VDD1.n0 VSUBS 3.65736f
C1077 VDD1.t0 VSUBS 0.436739f
C1078 VDD1.t5 VSUBS 0.436739f
C1079 VDD1.n1 VSUBS 3.65539f
C1080 VDD1.t6 VSUBS 0.436739f
C1081 VDD1.t4 VSUBS 0.436739f
C1082 VDD1.n2 VSUBS 3.65539f
C1083 VDD1.n3 VSUBS 5.96371f
C1084 VDD1.t7 VSUBS 0.436739f
C1085 VDD1.t1 VSUBS 0.436739f
C1086 VDD1.n4 VSUBS 3.63098f
C1087 VDD1.n5 VSUBS 5.01127f
C1088 VP.t3 VSUBS 4.04973f
C1089 VP.n0 VSUBS 1.49304f
C1090 VP.n1 VSUBS 0.023788f
C1091 VP.n2 VSUBS 0.028303f
C1092 VP.n3 VSUBS 0.023788f
C1093 VP.n4 VSUBS 0.02582f
C1094 VP.n5 VSUBS 0.023788f
C1095 VP.n6 VSUBS 0.019213f
C1096 VP.n7 VSUBS 0.023788f
C1097 VP.t2 VSUBS 4.04973f
C1098 VP.n8 VSUBS 1.39769f
C1099 VP.n9 VSUBS 0.023788f
C1100 VP.n10 VSUBS 0.040445f
C1101 VP.n11 VSUBS 0.023788f
C1102 VP.n12 VSUBS 0.03366f
C1103 VP.t6 VSUBS 4.04973f
C1104 VP.n13 VSUBS 1.49304f
C1105 VP.n14 VSUBS 0.023788f
C1106 VP.n15 VSUBS 0.028303f
C1107 VP.n16 VSUBS 0.023788f
C1108 VP.n17 VSUBS 0.02582f
C1109 VP.n18 VSUBS 0.023788f
C1110 VP.n19 VSUBS 0.019213f
C1111 VP.n20 VSUBS 0.023788f
C1112 VP.t4 VSUBS 4.04973f
C1113 VP.n21 VSUBS 1.48753f
C1114 VP.t5 VSUBS 4.39429f
C1115 VP.n22 VSUBS 1.41301f
C1116 VP.n23 VSUBS 0.292702f
C1117 VP.n24 VSUBS 0.040629f
C1118 VP.n25 VSUBS 0.044113f
C1119 VP.n26 VSUBS 0.04703f
C1120 VP.n27 VSUBS 0.023788f
C1121 VP.n28 VSUBS 0.023788f
C1122 VP.n29 VSUBS 0.023788f
C1123 VP.n30 VSUBS 0.04703f
C1124 VP.n31 VSUBS 0.044113f
C1125 VP.t0 VSUBS 4.04973f
C1126 VP.n32 VSUBS 1.39769f
C1127 VP.n33 VSUBS 0.040629f
C1128 VP.n34 VSUBS 0.023788f
C1129 VP.n35 VSUBS 0.023788f
C1130 VP.n36 VSUBS 0.023788f
C1131 VP.n37 VSUBS 0.044113f
C1132 VP.n38 VSUBS 0.044113f
C1133 VP.n39 VSUBS 0.040445f
C1134 VP.n40 VSUBS 0.023788f
C1135 VP.n41 VSUBS 0.023788f
C1136 VP.n42 VSUBS 0.023788f
C1137 VP.n43 VSUBS 0.044526f
C1138 VP.n44 VSUBS 0.044113f
C1139 VP.n45 VSUBS 0.03366f
C1140 VP.n46 VSUBS 0.038388f
C1141 VP.n47 VSUBS 1.72985f
C1142 VP.t7 VSUBS 4.04973f
C1143 VP.n48 VSUBS 1.49304f
C1144 VP.n49 VSUBS 1.74425f
C1145 VP.n50 VSUBS 0.038388f
C1146 VP.n51 VSUBS 0.023788f
C1147 VP.n52 VSUBS 0.044113f
C1148 VP.n53 VSUBS 0.044526f
C1149 VP.n54 VSUBS 0.028303f
C1150 VP.n55 VSUBS 0.023788f
C1151 VP.n56 VSUBS 0.023788f
C1152 VP.n57 VSUBS 0.023788f
C1153 VP.n58 VSUBS 0.044113f
C1154 VP.n59 VSUBS 0.044113f
C1155 VP.n60 VSUBS 0.02582f
C1156 VP.n61 VSUBS 0.023788f
C1157 VP.n62 VSUBS 0.023788f
C1158 VP.n63 VSUBS 0.040629f
C1159 VP.n64 VSUBS 0.044113f
C1160 VP.n65 VSUBS 0.04703f
C1161 VP.n66 VSUBS 0.023788f
C1162 VP.n67 VSUBS 0.023788f
C1163 VP.n68 VSUBS 0.023788f
C1164 VP.n69 VSUBS 0.04703f
C1165 VP.n70 VSUBS 0.044113f
C1166 VP.t1 VSUBS 4.04973f
C1167 VP.n71 VSUBS 1.39769f
C1168 VP.n72 VSUBS 0.040629f
C1169 VP.n73 VSUBS 0.023788f
C1170 VP.n74 VSUBS 0.023788f
C1171 VP.n75 VSUBS 0.023788f
C1172 VP.n76 VSUBS 0.044113f
C1173 VP.n77 VSUBS 0.044113f
C1174 VP.n78 VSUBS 0.040445f
C1175 VP.n79 VSUBS 0.023788f
C1176 VP.n80 VSUBS 0.023788f
C1177 VP.n81 VSUBS 0.023788f
C1178 VP.n82 VSUBS 0.044526f
C1179 VP.n83 VSUBS 0.044113f
C1180 VP.n84 VSUBS 0.03366f
C1181 VP.n85 VSUBS 0.038388f
C1182 VP.n86 VSUBS 0.061487f
C1183 VDD2.t0 VSUBS 0.435528f
C1184 VDD2.t5 VSUBS 0.435528f
C1185 VDD2.n0 VSUBS 3.64526f
C1186 VDD2.t1 VSUBS 0.435528f
C1187 VDD2.t7 VSUBS 0.435528f
C1188 VDD2.n1 VSUBS 3.64526f
C1189 VDD2.n2 VSUBS 5.88294f
C1190 VDD2.t6 VSUBS 0.435528f
C1191 VDD2.t4 VSUBS 0.435528f
C1192 VDD2.n3 VSUBS 3.62093f
C1193 VDD2.n4 VSUBS 4.9579f
C1194 VDD2.t2 VSUBS 0.435528f
C1195 VDD2.t3 VSUBS 0.435528f
C1196 VDD2.n5 VSUBS 3.6452f
C1197 VTAIL.t10 VSUBS 0.337964f
C1198 VTAIL.t12 VSUBS 0.337964f
C1199 VTAIL.n0 VSUBS 2.66851f
C1200 VTAIL.n1 VSUBS 0.839165f
C1201 VTAIL.n2 VSUBS 0.027361f
C1202 VTAIL.n3 VSUBS 0.024245f
C1203 VTAIL.n4 VSUBS 0.013028f
C1204 VTAIL.n5 VSUBS 0.030794f
C1205 VTAIL.n6 VSUBS 0.013794f
C1206 VTAIL.n7 VSUBS 0.024245f
C1207 VTAIL.n8 VSUBS 0.013028f
C1208 VTAIL.n9 VSUBS 0.030794f
C1209 VTAIL.n10 VSUBS 0.013411f
C1210 VTAIL.n11 VSUBS 0.024245f
C1211 VTAIL.n12 VSUBS 0.013794f
C1212 VTAIL.n13 VSUBS 0.030794f
C1213 VTAIL.n14 VSUBS 0.013794f
C1214 VTAIL.n15 VSUBS 0.024245f
C1215 VTAIL.n16 VSUBS 0.013028f
C1216 VTAIL.n17 VSUBS 0.030794f
C1217 VTAIL.n18 VSUBS 0.013794f
C1218 VTAIL.n19 VSUBS 0.024245f
C1219 VTAIL.n20 VSUBS 0.013028f
C1220 VTAIL.n21 VSUBS 0.030794f
C1221 VTAIL.n22 VSUBS 0.013794f
C1222 VTAIL.n23 VSUBS 0.024245f
C1223 VTAIL.n24 VSUBS 0.013028f
C1224 VTAIL.n25 VSUBS 0.030794f
C1225 VTAIL.n26 VSUBS 0.013794f
C1226 VTAIL.n27 VSUBS 0.024245f
C1227 VTAIL.n28 VSUBS 0.013028f
C1228 VTAIL.n29 VSUBS 0.030794f
C1229 VTAIL.n30 VSUBS 0.013794f
C1230 VTAIL.n31 VSUBS 1.83865f
C1231 VTAIL.n32 VSUBS 0.013028f
C1232 VTAIL.t9 VSUBS 0.066082f
C1233 VTAIL.n33 VSUBS 0.189784f
C1234 VTAIL.n34 VSUBS 0.01959f
C1235 VTAIL.n35 VSUBS 0.023095f
C1236 VTAIL.n36 VSUBS 0.030794f
C1237 VTAIL.n37 VSUBS 0.013794f
C1238 VTAIL.n38 VSUBS 0.013028f
C1239 VTAIL.n39 VSUBS 0.024245f
C1240 VTAIL.n40 VSUBS 0.024245f
C1241 VTAIL.n41 VSUBS 0.013028f
C1242 VTAIL.n42 VSUBS 0.013794f
C1243 VTAIL.n43 VSUBS 0.030794f
C1244 VTAIL.n44 VSUBS 0.030794f
C1245 VTAIL.n45 VSUBS 0.013794f
C1246 VTAIL.n46 VSUBS 0.013028f
C1247 VTAIL.n47 VSUBS 0.024245f
C1248 VTAIL.n48 VSUBS 0.024245f
C1249 VTAIL.n49 VSUBS 0.013028f
C1250 VTAIL.n50 VSUBS 0.013794f
C1251 VTAIL.n51 VSUBS 0.030794f
C1252 VTAIL.n52 VSUBS 0.030794f
C1253 VTAIL.n53 VSUBS 0.013794f
C1254 VTAIL.n54 VSUBS 0.013028f
C1255 VTAIL.n55 VSUBS 0.024245f
C1256 VTAIL.n56 VSUBS 0.024245f
C1257 VTAIL.n57 VSUBS 0.013028f
C1258 VTAIL.n58 VSUBS 0.013794f
C1259 VTAIL.n59 VSUBS 0.030794f
C1260 VTAIL.n60 VSUBS 0.030794f
C1261 VTAIL.n61 VSUBS 0.013794f
C1262 VTAIL.n62 VSUBS 0.013028f
C1263 VTAIL.n63 VSUBS 0.024245f
C1264 VTAIL.n64 VSUBS 0.024245f
C1265 VTAIL.n65 VSUBS 0.013028f
C1266 VTAIL.n66 VSUBS 0.013794f
C1267 VTAIL.n67 VSUBS 0.030794f
C1268 VTAIL.n68 VSUBS 0.030794f
C1269 VTAIL.n69 VSUBS 0.013794f
C1270 VTAIL.n70 VSUBS 0.013028f
C1271 VTAIL.n71 VSUBS 0.024245f
C1272 VTAIL.n72 VSUBS 0.024245f
C1273 VTAIL.n73 VSUBS 0.013028f
C1274 VTAIL.n74 VSUBS 0.013028f
C1275 VTAIL.n75 VSUBS 0.013794f
C1276 VTAIL.n76 VSUBS 0.030794f
C1277 VTAIL.n77 VSUBS 0.030794f
C1278 VTAIL.n78 VSUBS 0.030794f
C1279 VTAIL.n79 VSUBS 0.013411f
C1280 VTAIL.n80 VSUBS 0.013028f
C1281 VTAIL.n81 VSUBS 0.024245f
C1282 VTAIL.n82 VSUBS 0.024245f
C1283 VTAIL.n83 VSUBS 0.013028f
C1284 VTAIL.n84 VSUBS 0.013794f
C1285 VTAIL.n85 VSUBS 0.030794f
C1286 VTAIL.n86 VSUBS 0.030794f
C1287 VTAIL.n87 VSUBS 0.013794f
C1288 VTAIL.n88 VSUBS 0.013028f
C1289 VTAIL.n89 VSUBS 0.024245f
C1290 VTAIL.n90 VSUBS 0.024245f
C1291 VTAIL.n91 VSUBS 0.013028f
C1292 VTAIL.n92 VSUBS 0.013794f
C1293 VTAIL.n93 VSUBS 0.030794f
C1294 VTAIL.n94 VSUBS 0.077003f
C1295 VTAIL.n95 VSUBS 0.013794f
C1296 VTAIL.n96 VSUBS 0.013028f
C1297 VTAIL.n97 VSUBS 0.060015f
C1298 VTAIL.n98 VSUBS 0.038952f
C1299 VTAIL.n99 VSUBS 0.318269f
C1300 VTAIL.n100 VSUBS 0.027361f
C1301 VTAIL.n101 VSUBS 0.024245f
C1302 VTAIL.n102 VSUBS 0.013028f
C1303 VTAIL.n103 VSUBS 0.030794f
C1304 VTAIL.n104 VSUBS 0.013794f
C1305 VTAIL.n105 VSUBS 0.024245f
C1306 VTAIL.n106 VSUBS 0.013028f
C1307 VTAIL.n107 VSUBS 0.030794f
C1308 VTAIL.n108 VSUBS 0.013411f
C1309 VTAIL.n109 VSUBS 0.024245f
C1310 VTAIL.n110 VSUBS 0.013794f
C1311 VTAIL.n111 VSUBS 0.030794f
C1312 VTAIL.n112 VSUBS 0.013794f
C1313 VTAIL.n113 VSUBS 0.024245f
C1314 VTAIL.n114 VSUBS 0.013028f
C1315 VTAIL.n115 VSUBS 0.030794f
C1316 VTAIL.n116 VSUBS 0.013794f
C1317 VTAIL.n117 VSUBS 0.024245f
C1318 VTAIL.n118 VSUBS 0.013028f
C1319 VTAIL.n119 VSUBS 0.030794f
C1320 VTAIL.n120 VSUBS 0.013794f
C1321 VTAIL.n121 VSUBS 0.024245f
C1322 VTAIL.n122 VSUBS 0.013028f
C1323 VTAIL.n123 VSUBS 0.030794f
C1324 VTAIL.n124 VSUBS 0.013794f
C1325 VTAIL.n125 VSUBS 0.024245f
C1326 VTAIL.n126 VSUBS 0.013028f
C1327 VTAIL.n127 VSUBS 0.030794f
C1328 VTAIL.n128 VSUBS 0.013794f
C1329 VTAIL.n129 VSUBS 1.83865f
C1330 VTAIL.n130 VSUBS 0.013028f
C1331 VTAIL.t0 VSUBS 0.066082f
C1332 VTAIL.n131 VSUBS 0.189784f
C1333 VTAIL.n132 VSUBS 0.01959f
C1334 VTAIL.n133 VSUBS 0.023095f
C1335 VTAIL.n134 VSUBS 0.030794f
C1336 VTAIL.n135 VSUBS 0.013794f
C1337 VTAIL.n136 VSUBS 0.013028f
C1338 VTAIL.n137 VSUBS 0.024245f
C1339 VTAIL.n138 VSUBS 0.024245f
C1340 VTAIL.n139 VSUBS 0.013028f
C1341 VTAIL.n140 VSUBS 0.013794f
C1342 VTAIL.n141 VSUBS 0.030794f
C1343 VTAIL.n142 VSUBS 0.030794f
C1344 VTAIL.n143 VSUBS 0.013794f
C1345 VTAIL.n144 VSUBS 0.013028f
C1346 VTAIL.n145 VSUBS 0.024245f
C1347 VTAIL.n146 VSUBS 0.024245f
C1348 VTAIL.n147 VSUBS 0.013028f
C1349 VTAIL.n148 VSUBS 0.013794f
C1350 VTAIL.n149 VSUBS 0.030794f
C1351 VTAIL.n150 VSUBS 0.030794f
C1352 VTAIL.n151 VSUBS 0.013794f
C1353 VTAIL.n152 VSUBS 0.013028f
C1354 VTAIL.n153 VSUBS 0.024245f
C1355 VTAIL.n154 VSUBS 0.024245f
C1356 VTAIL.n155 VSUBS 0.013028f
C1357 VTAIL.n156 VSUBS 0.013794f
C1358 VTAIL.n157 VSUBS 0.030794f
C1359 VTAIL.n158 VSUBS 0.030794f
C1360 VTAIL.n159 VSUBS 0.013794f
C1361 VTAIL.n160 VSUBS 0.013028f
C1362 VTAIL.n161 VSUBS 0.024245f
C1363 VTAIL.n162 VSUBS 0.024245f
C1364 VTAIL.n163 VSUBS 0.013028f
C1365 VTAIL.n164 VSUBS 0.013794f
C1366 VTAIL.n165 VSUBS 0.030794f
C1367 VTAIL.n166 VSUBS 0.030794f
C1368 VTAIL.n167 VSUBS 0.013794f
C1369 VTAIL.n168 VSUBS 0.013028f
C1370 VTAIL.n169 VSUBS 0.024245f
C1371 VTAIL.n170 VSUBS 0.024245f
C1372 VTAIL.n171 VSUBS 0.013028f
C1373 VTAIL.n172 VSUBS 0.013028f
C1374 VTAIL.n173 VSUBS 0.013794f
C1375 VTAIL.n174 VSUBS 0.030794f
C1376 VTAIL.n175 VSUBS 0.030794f
C1377 VTAIL.n176 VSUBS 0.030794f
C1378 VTAIL.n177 VSUBS 0.013411f
C1379 VTAIL.n178 VSUBS 0.013028f
C1380 VTAIL.n179 VSUBS 0.024245f
C1381 VTAIL.n180 VSUBS 0.024245f
C1382 VTAIL.n181 VSUBS 0.013028f
C1383 VTAIL.n182 VSUBS 0.013794f
C1384 VTAIL.n183 VSUBS 0.030794f
C1385 VTAIL.n184 VSUBS 0.030794f
C1386 VTAIL.n185 VSUBS 0.013794f
C1387 VTAIL.n186 VSUBS 0.013028f
C1388 VTAIL.n187 VSUBS 0.024245f
C1389 VTAIL.n188 VSUBS 0.024245f
C1390 VTAIL.n189 VSUBS 0.013028f
C1391 VTAIL.n190 VSUBS 0.013794f
C1392 VTAIL.n191 VSUBS 0.030794f
C1393 VTAIL.n192 VSUBS 0.077003f
C1394 VTAIL.n193 VSUBS 0.013794f
C1395 VTAIL.n194 VSUBS 0.013028f
C1396 VTAIL.n195 VSUBS 0.060015f
C1397 VTAIL.n196 VSUBS 0.038952f
C1398 VTAIL.n197 VSUBS 0.318269f
C1399 VTAIL.t5 VSUBS 0.337964f
C1400 VTAIL.t6 VSUBS 0.337964f
C1401 VTAIL.n198 VSUBS 2.66851f
C1402 VTAIL.n199 VSUBS 1.09323f
C1403 VTAIL.n200 VSUBS 0.027361f
C1404 VTAIL.n201 VSUBS 0.024245f
C1405 VTAIL.n202 VSUBS 0.013028f
C1406 VTAIL.n203 VSUBS 0.030794f
C1407 VTAIL.n204 VSUBS 0.013794f
C1408 VTAIL.n205 VSUBS 0.024245f
C1409 VTAIL.n206 VSUBS 0.013028f
C1410 VTAIL.n207 VSUBS 0.030794f
C1411 VTAIL.n208 VSUBS 0.013411f
C1412 VTAIL.n209 VSUBS 0.024245f
C1413 VTAIL.n210 VSUBS 0.013794f
C1414 VTAIL.n211 VSUBS 0.030794f
C1415 VTAIL.n212 VSUBS 0.013794f
C1416 VTAIL.n213 VSUBS 0.024245f
C1417 VTAIL.n214 VSUBS 0.013028f
C1418 VTAIL.n215 VSUBS 0.030794f
C1419 VTAIL.n216 VSUBS 0.013794f
C1420 VTAIL.n217 VSUBS 0.024245f
C1421 VTAIL.n218 VSUBS 0.013028f
C1422 VTAIL.n219 VSUBS 0.030794f
C1423 VTAIL.n220 VSUBS 0.013794f
C1424 VTAIL.n221 VSUBS 0.024245f
C1425 VTAIL.n222 VSUBS 0.013028f
C1426 VTAIL.n223 VSUBS 0.030794f
C1427 VTAIL.n224 VSUBS 0.013794f
C1428 VTAIL.n225 VSUBS 0.024245f
C1429 VTAIL.n226 VSUBS 0.013028f
C1430 VTAIL.n227 VSUBS 0.030794f
C1431 VTAIL.n228 VSUBS 0.013794f
C1432 VTAIL.n229 VSUBS 1.83865f
C1433 VTAIL.n230 VSUBS 0.013028f
C1434 VTAIL.t1 VSUBS 0.066082f
C1435 VTAIL.n231 VSUBS 0.189784f
C1436 VTAIL.n232 VSUBS 0.01959f
C1437 VTAIL.n233 VSUBS 0.023095f
C1438 VTAIL.n234 VSUBS 0.030794f
C1439 VTAIL.n235 VSUBS 0.013794f
C1440 VTAIL.n236 VSUBS 0.013028f
C1441 VTAIL.n237 VSUBS 0.024245f
C1442 VTAIL.n238 VSUBS 0.024245f
C1443 VTAIL.n239 VSUBS 0.013028f
C1444 VTAIL.n240 VSUBS 0.013794f
C1445 VTAIL.n241 VSUBS 0.030794f
C1446 VTAIL.n242 VSUBS 0.030794f
C1447 VTAIL.n243 VSUBS 0.013794f
C1448 VTAIL.n244 VSUBS 0.013028f
C1449 VTAIL.n245 VSUBS 0.024245f
C1450 VTAIL.n246 VSUBS 0.024245f
C1451 VTAIL.n247 VSUBS 0.013028f
C1452 VTAIL.n248 VSUBS 0.013794f
C1453 VTAIL.n249 VSUBS 0.030794f
C1454 VTAIL.n250 VSUBS 0.030794f
C1455 VTAIL.n251 VSUBS 0.013794f
C1456 VTAIL.n252 VSUBS 0.013028f
C1457 VTAIL.n253 VSUBS 0.024245f
C1458 VTAIL.n254 VSUBS 0.024245f
C1459 VTAIL.n255 VSUBS 0.013028f
C1460 VTAIL.n256 VSUBS 0.013794f
C1461 VTAIL.n257 VSUBS 0.030794f
C1462 VTAIL.n258 VSUBS 0.030794f
C1463 VTAIL.n259 VSUBS 0.013794f
C1464 VTAIL.n260 VSUBS 0.013028f
C1465 VTAIL.n261 VSUBS 0.024245f
C1466 VTAIL.n262 VSUBS 0.024245f
C1467 VTAIL.n263 VSUBS 0.013028f
C1468 VTAIL.n264 VSUBS 0.013794f
C1469 VTAIL.n265 VSUBS 0.030794f
C1470 VTAIL.n266 VSUBS 0.030794f
C1471 VTAIL.n267 VSUBS 0.013794f
C1472 VTAIL.n268 VSUBS 0.013028f
C1473 VTAIL.n269 VSUBS 0.024245f
C1474 VTAIL.n270 VSUBS 0.024245f
C1475 VTAIL.n271 VSUBS 0.013028f
C1476 VTAIL.n272 VSUBS 0.013028f
C1477 VTAIL.n273 VSUBS 0.013794f
C1478 VTAIL.n274 VSUBS 0.030794f
C1479 VTAIL.n275 VSUBS 0.030794f
C1480 VTAIL.n276 VSUBS 0.030794f
C1481 VTAIL.n277 VSUBS 0.013411f
C1482 VTAIL.n278 VSUBS 0.013028f
C1483 VTAIL.n279 VSUBS 0.024245f
C1484 VTAIL.n280 VSUBS 0.024245f
C1485 VTAIL.n281 VSUBS 0.013028f
C1486 VTAIL.n282 VSUBS 0.013794f
C1487 VTAIL.n283 VSUBS 0.030794f
C1488 VTAIL.n284 VSUBS 0.030794f
C1489 VTAIL.n285 VSUBS 0.013794f
C1490 VTAIL.n286 VSUBS 0.013028f
C1491 VTAIL.n287 VSUBS 0.024245f
C1492 VTAIL.n288 VSUBS 0.024245f
C1493 VTAIL.n289 VSUBS 0.013028f
C1494 VTAIL.n290 VSUBS 0.013794f
C1495 VTAIL.n291 VSUBS 0.030794f
C1496 VTAIL.n292 VSUBS 0.077003f
C1497 VTAIL.n293 VSUBS 0.013794f
C1498 VTAIL.n294 VSUBS 0.013028f
C1499 VTAIL.n295 VSUBS 0.060015f
C1500 VTAIL.n296 VSUBS 0.038952f
C1501 VTAIL.n297 VSUBS 2.05751f
C1502 VTAIL.n298 VSUBS 0.027361f
C1503 VTAIL.n299 VSUBS 0.024245f
C1504 VTAIL.n300 VSUBS 0.013028f
C1505 VTAIL.n301 VSUBS 0.030794f
C1506 VTAIL.n302 VSUBS 0.013794f
C1507 VTAIL.n303 VSUBS 0.024245f
C1508 VTAIL.n304 VSUBS 0.013028f
C1509 VTAIL.n305 VSUBS 0.030794f
C1510 VTAIL.n306 VSUBS 0.013411f
C1511 VTAIL.n307 VSUBS 0.024245f
C1512 VTAIL.n308 VSUBS 0.013411f
C1513 VTAIL.n309 VSUBS 0.013028f
C1514 VTAIL.n310 VSUBS 0.030794f
C1515 VTAIL.n311 VSUBS 0.030794f
C1516 VTAIL.n312 VSUBS 0.013794f
C1517 VTAIL.n313 VSUBS 0.024245f
C1518 VTAIL.n314 VSUBS 0.013028f
C1519 VTAIL.n315 VSUBS 0.030794f
C1520 VTAIL.n316 VSUBS 0.013794f
C1521 VTAIL.n317 VSUBS 0.024245f
C1522 VTAIL.n318 VSUBS 0.013028f
C1523 VTAIL.n319 VSUBS 0.030794f
C1524 VTAIL.n320 VSUBS 0.013794f
C1525 VTAIL.n321 VSUBS 0.024245f
C1526 VTAIL.n322 VSUBS 0.013028f
C1527 VTAIL.n323 VSUBS 0.030794f
C1528 VTAIL.n324 VSUBS 0.013794f
C1529 VTAIL.n325 VSUBS 0.024245f
C1530 VTAIL.n326 VSUBS 0.013028f
C1531 VTAIL.n327 VSUBS 0.030794f
C1532 VTAIL.n328 VSUBS 0.013794f
C1533 VTAIL.n329 VSUBS 1.83865f
C1534 VTAIL.n330 VSUBS 0.013028f
C1535 VTAIL.t13 VSUBS 0.066082f
C1536 VTAIL.n331 VSUBS 0.189784f
C1537 VTAIL.n332 VSUBS 0.01959f
C1538 VTAIL.n333 VSUBS 0.023095f
C1539 VTAIL.n334 VSUBS 0.030794f
C1540 VTAIL.n335 VSUBS 0.013794f
C1541 VTAIL.n336 VSUBS 0.013028f
C1542 VTAIL.n337 VSUBS 0.024245f
C1543 VTAIL.n338 VSUBS 0.024245f
C1544 VTAIL.n339 VSUBS 0.013028f
C1545 VTAIL.n340 VSUBS 0.013794f
C1546 VTAIL.n341 VSUBS 0.030794f
C1547 VTAIL.n342 VSUBS 0.030794f
C1548 VTAIL.n343 VSUBS 0.013794f
C1549 VTAIL.n344 VSUBS 0.013028f
C1550 VTAIL.n345 VSUBS 0.024245f
C1551 VTAIL.n346 VSUBS 0.024245f
C1552 VTAIL.n347 VSUBS 0.013028f
C1553 VTAIL.n348 VSUBS 0.013794f
C1554 VTAIL.n349 VSUBS 0.030794f
C1555 VTAIL.n350 VSUBS 0.030794f
C1556 VTAIL.n351 VSUBS 0.013794f
C1557 VTAIL.n352 VSUBS 0.013028f
C1558 VTAIL.n353 VSUBS 0.024245f
C1559 VTAIL.n354 VSUBS 0.024245f
C1560 VTAIL.n355 VSUBS 0.013028f
C1561 VTAIL.n356 VSUBS 0.013794f
C1562 VTAIL.n357 VSUBS 0.030794f
C1563 VTAIL.n358 VSUBS 0.030794f
C1564 VTAIL.n359 VSUBS 0.013794f
C1565 VTAIL.n360 VSUBS 0.013028f
C1566 VTAIL.n361 VSUBS 0.024245f
C1567 VTAIL.n362 VSUBS 0.024245f
C1568 VTAIL.n363 VSUBS 0.013028f
C1569 VTAIL.n364 VSUBS 0.013794f
C1570 VTAIL.n365 VSUBS 0.030794f
C1571 VTAIL.n366 VSUBS 0.030794f
C1572 VTAIL.n367 VSUBS 0.013794f
C1573 VTAIL.n368 VSUBS 0.013028f
C1574 VTAIL.n369 VSUBS 0.024245f
C1575 VTAIL.n370 VSUBS 0.024245f
C1576 VTAIL.n371 VSUBS 0.013028f
C1577 VTAIL.n372 VSUBS 0.013794f
C1578 VTAIL.n373 VSUBS 0.030794f
C1579 VTAIL.n374 VSUBS 0.030794f
C1580 VTAIL.n375 VSUBS 0.013794f
C1581 VTAIL.n376 VSUBS 0.013028f
C1582 VTAIL.n377 VSUBS 0.024245f
C1583 VTAIL.n378 VSUBS 0.024245f
C1584 VTAIL.n379 VSUBS 0.013028f
C1585 VTAIL.n380 VSUBS 0.013794f
C1586 VTAIL.n381 VSUBS 0.030794f
C1587 VTAIL.n382 VSUBS 0.030794f
C1588 VTAIL.n383 VSUBS 0.013794f
C1589 VTAIL.n384 VSUBS 0.013028f
C1590 VTAIL.n385 VSUBS 0.024245f
C1591 VTAIL.n386 VSUBS 0.024245f
C1592 VTAIL.n387 VSUBS 0.013028f
C1593 VTAIL.n388 VSUBS 0.013794f
C1594 VTAIL.n389 VSUBS 0.030794f
C1595 VTAIL.n390 VSUBS 0.077003f
C1596 VTAIL.n391 VSUBS 0.013794f
C1597 VTAIL.n392 VSUBS 0.013028f
C1598 VTAIL.n393 VSUBS 0.060015f
C1599 VTAIL.n394 VSUBS 0.038952f
C1600 VTAIL.n395 VSUBS 2.05751f
C1601 VTAIL.t11 VSUBS 0.337964f
C1602 VTAIL.t15 VSUBS 0.337964f
C1603 VTAIL.n396 VSUBS 2.66852f
C1604 VTAIL.n397 VSUBS 1.09322f
C1605 VTAIL.n398 VSUBS 0.027361f
C1606 VTAIL.n399 VSUBS 0.024245f
C1607 VTAIL.n400 VSUBS 0.013028f
C1608 VTAIL.n401 VSUBS 0.030794f
C1609 VTAIL.n402 VSUBS 0.013794f
C1610 VTAIL.n403 VSUBS 0.024245f
C1611 VTAIL.n404 VSUBS 0.013028f
C1612 VTAIL.n405 VSUBS 0.030794f
C1613 VTAIL.n406 VSUBS 0.013411f
C1614 VTAIL.n407 VSUBS 0.024245f
C1615 VTAIL.n408 VSUBS 0.013411f
C1616 VTAIL.n409 VSUBS 0.013028f
C1617 VTAIL.n410 VSUBS 0.030794f
C1618 VTAIL.n411 VSUBS 0.030794f
C1619 VTAIL.n412 VSUBS 0.013794f
C1620 VTAIL.n413 VSUBS 0.024245f
C1621 VTAIL.n414 VSUBS 0.013028f
C1622 VTAIL.n415 VSUBS 0.030794f
C1623 VTAIL.n416 VSUBS 0.013794f
C1624 VTAIL.n417 VSUBS 0.024245f
C1625 VTAIL.n418 VSUBS 0.013028f
C1626 VTAIL.n419 VSUBS 0.030794f
C1627 VTAIL.n420 VSUBS 0.013794f
C1628 VTAIL.n421 VSUBS 0.024245f
C1629 VTAIL.n422 VSUBS 0.013028f
C1630 VTAIL.n423 VSUBS 0.030794f
C1631 VTAIL.n424 VSUBS 0.013794f
C1632 VTAIL.n425 VSUBS 0.024245f
C1633 VTAIL.n426 VSUBS 0.013028f
C1634 VTAIL.n427 VSUBS 0.030794f
C1635 VTAIL.n428 VSUBS 0.013794f
C1636 VTAIL.n429 VSUBS 1.83865f
C1637 VTAIL.n430 VSUBS 0.013028f
C1638 VTAIL.t8 VSUBS 0.066082f
C1639 VTAIL.n431 VSUBS 0.189784f
C1640 VTAIL.n432 VSUBS 0.01959f
C1641 VTAIL.n433 VSUBS 0.023095f
C1642 VTAIL.n434 VSUBS 0.030794f
C1643 VTAIL.n435 VSUBS 0.013794f
C1644 VTAIL.n436 VSUBS 0.013028f
C1645 VTAIL.n437 VSUBS 0.024245f
C1646 VTAIL.n438 VSUBS 0.024245f
C1647 VTAIL.n439 VSUBS 0.013028f
C1648 VTAIL.n440 VSUBS 0.013794f
C1649 VTAIL.n441 VSUBS 0.030794f
C1650 VTAIL.n442 VSUBS 0.030794f
C1651 VTAIL.n443 VSUBS 0.013794f
C1652 VTAIL.n444 VSUBS 0.013028f
C1653 VTAIL.n445 VSUBS 0.024245f
C1654 VTAIL.n446 VSUBS 0.024245f
C1655 VTAIL.n447 VSUBS 0.013028f
C1656 VTAIL.n448 VSUBS 0.013794f
C1657 VTAIL.n449 VSUBS 0.030794f
C1658 VTAIL.n450 VSUBS 0.030794f
C1659 VTAIL.n451 VSUBS 0.013794f
C1660 VTAIL.n452 VSUBS 0.013028f
C1661 VTAIL.n453 VSUBS 0.024245f
C1662 VTAIL.n454 VSUBS 0.024245f
C1663 VTAIL.n455 VSUBS 0.013028f
C1664 VTAIL.n456 VSUBS 0.013794f
C1665 VTAIL.n457 VSUBS 0.030794f
C1666 VTAIL.n458 VSUBS 0.030794f
C1667 VTAIL.n459 VSUBS 0.013794f
C1668 VTAIL.n460 VSUBS 0.013028f
C1669 VTAIL.n461 VSUBS 0.024245f
C1670 VTAIL.n462 VSUBS 0.024245f
C1671 VTAIL.n463 VSUBS 0.013028f
C1672 VTAIL.n464 VSUBS 0.013794f
C1673 VTAIL.n465 VSUBS 0.030794f
C1674 VTAIL.n466 VSUBS 0.030794f
C1675 VTAIL.n467 VSUBS 0.013794f
C1676 VTAIL.n468 VSUBS 0.013028f
C1677 VTAIL.n469 VSUBS 0.024245f
C1678 VTAIL.n470 VSUBS 0.024245f
C1679 VTAIL.n471 VSUBS 0.013028f
C1680 VTAIL.n472 VSUBS 0.013794f
C1681 VTAIL.n473 VSUBS 0.030794f
C1682 VTAIL.n474 VSUBS 0.030794f
C1683 VTAIL.n475 VSUBS 0.013794f
C1684 VTAIL.n476 VSUBS 0.013028f
C1685 VTAIL.n477 VSUBS 0.024245f
C1686 VTAIL.n478 VSUBS 0.024245f
C1687 VTAIL.n479 VSUBS 0.013028f
C1688 VTAIL.n480 VSUBS 0.013794f
C1689 VTAIL.n481 VSUBS 0.030794f
C1690 VTAIL.n482 VSUBS 0.030794f
C1691 VTAIL.n483 VSUBS 0.013794f
C1692 VTAIL.n484 VSUBS 0.013028f
C1693 VTAIL.n485 VSUBS 0.024245f
C1694 VTAIL.n486 VSUBS 0.024245f
C1695 VTAIL.n487 VSUBS 0.013028f
C1696 VTAIL.n488 VSUBS 0.013794f
C1697 VTAIL.n489 VSUBS 0.030794f
C1698 VTAIL.n490 VSUBS 0.077003f
C1699 VTAIL.n491 VSUBS 0.013794f
C1700 VTAIL.n492 VSUBS 0.013028f
C1701 VTAIL.n493 VSUBS 0.060015f
C1702 VTAIL.n494 VSUBS 0.038952f
C1703 VTAIL.n495 VSUBS 0.318269f
C1704 VTAIL.n496 VSUBS 0.027361f
C1705 VTAIL.n497 VSUBS 0.024245f
C1706 VTAIL.n498 VSUBS 0.013028f
C1707 VTAIL.n499 VSUBS 0.030794f
C1708 VTAIL.n500 VSUBS 0.013794f
C1709 VTAIL.n501 VSUBS 0.024245f
C1710 VTAIL.n502 VSUBS 0.013028f
C1711 VTAIL.n503 VSUBS 0.030794f
C1712 VTAIL.n504 VSUBS 0.013411f
C1713 VTAIL.n505 VSUBS 0.024245f
C1714 VTAIL.n506 VSUBS 0.013411f
C1715 VTAIL.n507 VSUBS 0.013028f
C1716 VTAIL.n508 VSUBS 0.030794f
C1717 VTAIL.n509 VSUBS 0.030794f
C1718 VTAIL.n510 VSUBS 0.013794f
C1719 VTAIL.n511 VSUBS 0.024245f
C1720 VTAIL.n512 VSUBS 0.013028f
C1721 VTAIL.n513 VSUBS 0.030794f
C1722 VTAIL.n514 VSUBS 0.013794f
C1723 VTAIL.n515 VSUBS 0.024245f
C1724 VTAIL.n516 VSUBS 0.013028f
C1725 VTAIL.n517 VSUBS 0.030794f
C1726 VTAIL.n518 VSUBS 0.013794f
C1727 VTAIL.n519 VSUBS 0.024245f
C1728 VTAIL.n520 VSUBS 0.013028f
C1729 VTAIL.n521 VSUBS 0.030794f
C1730 VTAIL.n522 VSUBS 0.013794f
C1731 VTAIL.n523 VSUBS 0.024245f
C1732 VTAIL.n524 VSUBS 0.013028f
C1733 VTAIL.n525 VSUBS 0.030794f
C1734 VTAIL.n526 VSUBS 0.013794f
C1735 VTAIL.n527 VSUBS 1.83865f
C1736 VTAIL.n528 VSUBS 0.013028f
C1737 VTAIL.t3 VSUBS 0.066082f
C1738 VTAIL.n529 VSUBS 0.189784f
C1739 VTAIL.n530 VSUBS 0.01959f
C1740 VTAIL.n531 VSUBS 0.023095f
C1741 VTAIL.n532 VSUBS 0.030794f
C1742 VTAIL.n533 VSUBS 0.013794f
C1743 VTAIL.n534 VSUBS 0.013028f
C1744 VTAIL.n535 VSUBS 0.024245f
C1745 VTAIL.n536 VSUBS 0.024245f
C1746 VTAIL.n537 VSUBS 0.013028f
C1747 VTAIL.n538 VSUBS 0.013794f
C1748 VTAIL.n539 VSUBS 0.030794f
C1749 VTAIL.n540 VSUBS 0.030794f
C1750 VTAIL.n541 VSUBS 0.013794f
C1751 VTAIL.n542 VSUBS 0.013028f
C1752 VTAIL.n543 VSUBS 0.024245f
C1753 VTAIL.n544 VSUBS 0.024245f
C1754 VTAIL.n545 VSUBS 0.013028f
C1755 VTAIL.n546 VSUBS 0.013794f
C1756 VTAIL.n547 VSUBS 0.030794f
C1757 VTAIL.n548 VSUBS 0.030794f
C1758 VTAIL.n549 VSUBS 0.013794f
C1759 VTAIL.n550 VSUBS 0.013028f
C1760 VTAIL.n551 VSUBS 0.024245f
C1761 VTAIL.n552 VSUBS 0.024245f
C1762 VTAIL.n553 VSUBS 0.013028f
C1763 VTAIL.n554 VSUBS 0.013794f
C1764 VTAIL.n555 VSUBS 0.030794f
C1765 VTAIL.n556 VSUBS 0.030794f
C1766 VTAIL.n557 VSUBS 0.013794f
C1767 VTAIL.n558 VSUBS 0.013028f
C1768 VTAIL.n559 VSUBS 0.024245f
C1769 VTAIL.n560 VSUBS 0.024245f
C1770 VTAIL.n561 VSUBS 0.013028f
C1771 VTAIL.n562 VSUBS 0.013794f
C1772 VTAIL.n563 VSUBS 0.030794f
C1773 VTAIL.n564 VSUBS 0.030794f
C1774 VTAIL.n565 VSUBS 0.013794f
C1775 VTAIL.n566 VSUBS 0.013028f
C1776 VTAIL.n567 VSUBS 0.024245f
C1777 VTAIL.n568 VSUBS 0.024245f
C1778 VTAIL.n569 VSUBS 0.013028f
C1779 VTAIL.n570 VSUBS 0.013794f
C1780 VTAIL.n571 VSUBS 0.030794f
C1781 VTAIL.n572 VSUBS 0.030794f
C1782 VTAIL.n573 VSUBS 0.013794f
C1783 VTAIL.n574 VSUBS 0.013028f
C1784 VTAIL.n575 VSUBS 0.024245f
C1785 VTAIL.n576 VSUBS 0.024245f
C1786 VTAIL.n577 VSUBS 0.013028f
C1787 VTAIL.n578 VSUBS 0.013794f
C1788 VTAIL.n579 VSUBS 0.030794f
C1789 VTAIL.n580 VSUBS 0.030794f
C1790 VTAIL.n581 VSUBS 0.013794f
C1791 VTAIL.n582 VSUBS 0.013028f
C1792 VTAIL.n583 VSUBS 0.024245f
C1793 VTAIL.n584 VSUBS 0.024245f
C1794 VTAIL.n585 VSUBS 0.013028f
C1795 VTAIL.n586 VSUBS 0.013794f
C1796 VTAIL.n587 VSUBS 0.030794f
C1797 VTAIL.n588 VSUBS 0.077003f
C1798 VTAIL.n589 VSUBS 0.013794f
C1799 VTAIL.n590 VSUBS 0.013028f
C1800 VTAIL.n591 VSUBS 0.060015f
C1801 VTAIL.n592 VSUBS 0.038952f
C1802 VTAIL.n593 VSUBS 0.318269f
C1803 VTAIL.t4 VSUBS 0.337964f
C1804 VTAIL.t2 VSUBS 0.337964f
C1805 VTAIL.n594 VSUBS 2.66852f
C1806 VTAIL.n595 VSUBS 1.09322f
C1807 VTAIL.n596 VSUBS 0.027361f
C1808 VTAIL.n597 VSUBS 0.024245f
C1809 VTAIL.n598 VSUBS 0.013028f
C1810 VTAIL.n599 VSUBS 0.030794f
C1811 VTAIL.n600 VSUBS 0.013794f
C1812 VTAIL.n601 VSUBS 0.024245f
C1813 VTAIL.n602 VSUBS 0.013028f
C1814 VTAIL.n603 VSUBS 0.030794f
C1815 VTAIL.n604 VSUBS 0.013411f
C1816 VTAIL.n605 VSUBS 0.024245f
C1817 VTAIL.n606 VSUBS 0.013411f
C1818 VTAIL.n607 VSUBS 0.013028f
C1819 VTAIL.n608 VSUBS 0.030794f
C1820 VTAIL.n609 VSUBS 0.030794f
C1821 VTAIL.n610 VSUBS 0.013794f
C1822 VTAIL.n611 VSUBS 0.024245f
C1823 VTAIL.n612 VSUBS 0.013028f
C1824 VTAIL.n613 VSUBS 0.030794f
C1825 VTAIL.n614 VSUBS 0.013794f
C1826 VTAIL.n615 VSUBS 0.024245f
C1827 VTAIL.n616 VSUBS 0.013028f
C1828 VTAIL.n617 VSUBS 0.030794f
C1829 VTAIL.n618 VSUBS 0.013794f
C1830 VTAIL.n619 VSUBS 0.024245f
C1831 VTAIL.n620 VSUBS 0.013028f
C1832 VTAIL.n621 VSUBS 0.030794f
C1833 VTAIL.n622 VSUBS 0.013794f
C1834 VTAIL.n623 VSUBS 0.024245f
C1835 VTAIL.n624 VSUBS 0.013028f
C1836 VTAIL.n625 VSUBS 0.030794f
C1837 VTAIL.n626 VSUBS 0.013794f
C1838 VTAIL.n627 VSUBS 1.83865f
C1839 VTAIL.n628 VSUBS 0.013028f
C1840 VTAIL.t7 VSUBS 0.066082f
C1841 VTAIL.n629 VSUBS 0.189784f
C1842 VTAIL.n630 VSUBS 0.01959f
C1843 VTAIL.n631 VSUBS 0.023095f
C1844 VTAIL.n632 VSUBS 0.030794f
C1845 VTAIL.n633 VSUBS 0.013794f
C1846 VTAIL.n634 VSUBS 0.013028f
C1847 VTAIL.n635 VSUBS 0.024245f
C1848 VTAIL.n636 VSUBS 0.024245f
C1849 VTAIL.n637 VSUBS 0.013028f
C1850 VTAIL.n638 VSUBS 0.013794f
C1851 VTAIL.n639 VSUBS 0.030794f
C1852 VTAIL.n640 VSUBS 0.030794f
C1853 VTAIL.n641 VSUBS 0.013794f
C1854 VTAIL.n642 VSUBS 0.013028f
C1855 VTAIL.n643 VSUBS 0.024245f
C1856 VTAIL.n644 VSUBS 0.024245f
C1857 VTAIL.n645 VSUBS 0.013028f
C1858 VTAIL.n646 VSUBS 0.013794f
C1859 VTAIL.n647 VSUBS 0.030794f
C1860 VTAIL.n648 VSUBS 0.030794f
C1861 VTAIL.n649 VSUBS 0.013794f
C1862 VTAIL.n650 VSUBS 0.013028f
C1863 VTAIL.n651 VSUBS 0.024245f
C1864 VTAIL.n652 VSUBS 0.024245f
C1865 VTAIL.n653 VSUBS 0.013028f
C1866 VTAIL.n654 VSUBS 0.013794f
C1867 VTAIL.n655 VSUBS 0.030794f
C1868 VTAIL.n656 VSUBS 0.030794f
C1869 VTAIL.n657 VSUBS 0.013794f
C1870 VTAIL.n658 VSUBS 0.013028f
C1871 VTAIL.n659 VSUBS 0.024245f
C1872 VTAIL.n660 VSUBS 0.024245f
C1873 VTAIL.n661 VSUBS 0.013028f
C1874 VTAIL.n662 VSUBS 0.013794f
C1875 VTAIL.n663 VSUBS 0.030794f
C1876 VTAIL.n664 VSUBS 0.030794f
C1877 VTAIL.n665 VSUBS 0.013794f
C1878 VTAIL.n666 VSUBS 0.013028f
C1879 VTAIL.n667 VSUBS 0.024245f
C1880 VTAIL.n668 VSUBS 0.024245f
C1881 VTAIL.n669 VSUBS 0.013028f
C1882 VTAIL.n670 VSUBS 0.013794f
C1883 VTAIL.n671 VSUBS 0.030794f
C1884 VTAIL.n672 VSUBS 0.030794f
C1885 VTAIL.n673 VSUBS 0.013794f
C1886 VTAIL.n674 VSUBS 0.013028f
C1887 VTAIL.n675 VSUBS 0.024245f
C1888 VTAIL.n676 VSUBS 0.024245f
C1889 VTAIL.n677 VSUBS 0.013028f
C1890 VTAIL.n678 VSUBS 0.013794f
C1891 VTAIL.n679 VSUBS 0.030794f
C1892 VTAIL.n680 VSUBS 0.030794f
C1893 VTAIL.n681 VSUBS 0.013794f
C1894 VTAIL.n682 VSUBS 0.013028f
C1895 VTAIL.n683 VSUBS 0.024245f
C1896 VTAIL.n684 VSUBS 0.024245f
C1897 VTAIL.n685 VSUBS 0.013028f
C1898 VTAIL.n686 VSUBS 0.013794f
C1899 VTAIL.n687 VSUBS 0.030794f
C1900 VTAIL.n688 VSUBS 0.077003f
C1901 VTAIL.n689 VSUBS 0.013794f
C1902 VTAIL.n690 VSUBS 0.013028f
C1903 VTAIL.n691 VSUBS 0.060015f
C1904 VTAIL.n692 VSUBS 0.038952f
C1905 VTAIL.n693 VSUBS 2.05751f
C1906 VTAIL.n694 VSUBS 0.027361f
C1907 VTAIL.n695 VSUBS 0.024245f
C1908 VTAIL.n696 VSUBS 0.013028f
C1909 VTAIL.n697 VSUBS 0.030794f
C1910 VTAIL.n698 VSUBS 0.013794f
C1911 VTAIL.n699 VSUBS 0.024245f
C1912 VTAIL.n700 VSUBS 0.013028f
C1913 VTAIL.n701 VSUBS 0.030794f
C1914 VTAIL.n702 VSUBS 0.013411f
C1915 VTAIL.n703 VSUBS 0.024245f
C1916 VTAIL.n704 VSUBS 0.013794f
C1917 VTAIL.n705 VSUBS 0.030794f
C1918 VTAIL.n706 VSUBS 0.013794f
C1919 VTAIL.n707 VSUBS 0.024245f
C1920 VTAIL.n708 VSUBS 0.013028f
C1921 VTAIL.n709 VSUBS 0.030794f
C1922 VTAIL.n710 VSUBS 0.013794f
C1923 VTAIL.n711 VSUBS 0.024245f
C1924 VTAIL.n712 VSUBS 0.013028f
C1925 VTAIL.n713 VSUBS 0.030794f
C1926 VTAIL.n714 VSUBS 0.013794f
C1927 VTAIL.n715 VSUBS 0.024245f
C1928 VTAIL.n716 VSUBS 0.013028f
C1929 VTAIL.n717 VSUBS 0.030794f
C1930 VTAIL.n718 VSUBS 0.013794f
C1931 VTAIL.n719 VSUBS 0.024245f
C1932 VTAIL.n720 VSUBS 0.013028f
C1933 VTAIL.n721 VSUBS 0.030794f
C1934 VTAIL.n722 VSUBS 0.013794f
C1935 VTAIL.n723 VSUBS 1.83865f
C1936 VTAIL.n724 VSUBS 0.013028f
C1937 VTAIL.t14 VSUBS 0.066082f
C1938 VTAIL.n725 VSUBS 0.189784f
C1939 VTAIL.n726 VSUBS 0.01959f
C1940 VTAIL.n727 VSUBS 0.023095f
C1941 VTAIL.n728 VSUBS 0.030794f
C1942 VTAIL.n729 VSUBS 0.013794f
C1943 VTAIL.n730 VSUBS 0.013028f
C1944 VTAIL.n731 VSUBS 0.024245f
C1945 VTAIL.n732 VSUBS 0.024245f
C1946 VTAIL.n733 VSUBS 0.013028f
C1947 VTAIL.n734 VSUBS 0.013794f
C1948 VTAIL.n735 VSUBS 0.030794f
C1949 VTAIL.n736 VSUBS 0.030794f
C1950 VTAIL.n737 VSUBS 0.013794f
C1951 VTAIL.n738 VSUBS 0.013028f
C1952 VTAIL.n739 VSUBS 0.024245f
C1953 VTAIL.n740 VSUBS 0.024245f
C1954 VTAIL.n741 VSUBS 0.013028f
C1955 VTAIL.n742 VSUBS 0.013794f
C1956 VTAIL.n743 VSUBS 0.030794f
C1957 VTAIL.n744 VSUBS 0.030794f
C1958 VTAIL.n745 VSUBS 0.013794f
C1959 VTAIL.n746 VSUBS 0.013028f
C1960 VTAIL.n747 VSUBS 0.024245f
C1961 VTAIL.n748 VSUBS 0.024245f
C1962 VTAIL.n749 VSUBS 0.013028f
C1963 VTAIL.n750 VSUBS 0.013794f
C1964 VTAIL.n751 VSUBS 0.030794f
C1965 VTAIL.n752 VSUBS 0.030794f
C1966 VTAIL.n753 VSUBS 0.013794f
C1967 VTAIL.n754 VSUBS 0.013028f
C1968 VTAIL.n755 VSUBS 0.024245f
C1969 VTAIL.n756 VSUBS 0.024245f
C1970 VTAIL.n757 VSUBS 0.013028f
C1971 VTAIL.n758 VSUBS 0.013794f
C1972 VTAIL.n759 VSUBS 0.030794f
C1973 VTAIL.n760 VSUBS 0.030794f
C1974 VTAIL.n761 VSUBS 0.013794f
C1975 VTAIL.n762 VSUBS 0.013028f
C1976 VTAIL.n763 VSUBS 0.024245f
C1977 VTAIL.n764 VSUBS 0.024245f
C1978 VTAIL.n765 VSUBS 0.013028f
C1979 VTAIL.n766 VSUBS 0.013028f
C1980 VTAIL.n767 VSUBS 0.013794f
C1981 VTAIL.n768 VSUBS 0.030794f
C1982 VTAIL.n769 VSUBS 0.030794f
C1983 VTAIL.n770 VSUBS 0.030794f
C1984 VTAIL.n771 VSUBS 0.013411f
C1985 VTAIL.n772 VSUBS 0.013028f
C1986 VTAIL.n773 VSUBS 0.024245f
C1987 VTAIL.n774 VSUBS 0.024245f
C1988 VTAIL.n775 VSUBS 0.013028f
C1989 VTAIL.n776 VSUBS 0.013794f
C1990 VTAIL.n777 VSUBS 0.030794f
C1991 VTAIL.n778 VSUBS 0.030794f
C1992 VTAIL.n779 VSUBS 0.013794f
C1993 VTAIL.n780 VSUBS 0.013028f
C1994 VTAIL.n781 VSUBS 0.024245f
C1995 VTAIL.n782 VSUBS 0.024245f
C1996 VTAIL.n783 VSUBS 0.013028f
C1997 VTAIL.n784 VSUBS 0.013794f
C1998 VTAIL.n785 VSUBS 0.030794f
C1999 VTAIL.n786 VSUBS 0.077003f
C2000 VTAIL.n787 VSUBS 0.013794f
C2001 VTAIL.n788 VSUBS 0.013028f
C2002 VTAIL.n789 VSUBS 0.060015f
C2003 VTAIL.n790 VSUBS 0.038952f
C2004 VTAIL.n791 VSUBS 2.05296f
C2005 VN.t0 VSUBS 3.74313f
C2006 VN.n0 VSUBS 1.38001f
C2007 VN.n1 VSUBS 0.021987f
C2008 VN.n2 VSUBS 0.02616f
C2009 VN.n3 VSUBS 0.021987f
C2010 VN.n4 VSUBS 0.023865f
C2011 VN.n5 VSUBS 0.021987f
C2012 VN.n6 VSUBS 0.017758f
C2013 VN.n7 VSUBS 0.021987f
C2014 VN.t2 VSUBS 3.74313f
C2015 VN.n8 VSUBS 1.37491f
C2016 VN.t7 VSUBS 4.0616f
C2017 VN.n9 VSUBS 1.30603f
C2018 VN.n10 VSUBS 0.270541f
C2019 VN.n11 VSUBS 0.037553f
C2020 VN.n12 VSUBS 0.040774f
C2021 VN.n13 VSUBS 0.04347f
C2022 VN.n14 VSUBS 0.021987f
C2023 VN.n15 VSUBS 0.021987f
C2024 VN.n16 VSUBS 0.021987f
C2025 VN.n17 VSUBS 0.04347f
C2026 VN.n18 VSUBS 0.040774f
C2027 VN.t6 VSUBS 3.74313f
C2028 VN.n19 VSUBS 1.29187f
C2029 VN.n20 VSUBS 0.037553f
C2030 VN.n21 VSUBS 0.021987f
C2031 VN.n22 VSUBS 0.021987f
C2032 VN.n23 VSUBS 0.021987f
C2033 VN.n24 VSUBS 0.040774f
C2034 VN.n25 VSUBS 0.040774f
C2035 VN.n26 VSUBS 0.037383f
C2036 VN.n27 VSUBS 0.021987f
C2037 VN.n28 VSUBS 0.021987f
C2038 VN.n29 VSUBS 0.021987f
C2039 VN.n30 VSUBS 0.041155f
C2040 VN.n31 VSUBS 0.040774f
C2041 VN.n32 VSUBS 0.031112f
C2042 VN.n33 VSUBS 0.035481f
C2043 VN.n34 VSUBS 0.056832f
C2044 VN.t1 VSUBS 3.74313f
C2045 VN.n35 VSUBS 1.38001f
C2046 VN.n36 VSUBS 0.021987f
C2047 VN.n37 VSUBS 0.02616f
C2048 VN.n38 VSUBS 0.021987f
C2049 VN.n39 VSUBS 0.023865f
C2050 VN.n40 VSUBS 0.021987f
C2051 VN.t3 VSUBS 3.74313f
C2052 VN.n41 VSUBS 1.29187f
C2053 VN.n42 VSUBS 0.017758f
C2054 VN.n43 VSUBS 0.021987f
C2055 VN.t5 VSUBS 3.74313f
C2056 VN.n44 VSUBS 1.37491f
C2057 VN.t4 VSUBS 4.0616f
C2058 VN.n45 VSUBS 1.30603f
C2059 VN.n46 VSUBS 0.270541f
C2060 VN.n47 VSUBS 0.037553f
C2061 VN.n48 VSUBS 0.040774f
C2062 VN.n49 VSUBS 0.04347f
C2063 VN.n50 VSUBS 0.021987f
C2064 VN.n51 VSUBS 0.021987f
C2065 VN.n52 VSUBS 0.021987f
C2066 VN.n53 VSUBS 0.04347f
C2067 VN.n54 VSUBS 0.040774f
C2068 VN.n55 VSUBS 0.037553f
C2069 VN.n56 VSUBS 0.021987f
C2070 VN.n57 VSUBS 0.021987f
C2071 VN.n58 VSUBS 0.021987f
C2072 VN.n59 VSUBS 0.040774f
C2073 VN.n60 VSUBS 0.040774f
C2074 VN.n61 VSUBS 0.037383f
C2075 VN.n62 VSUBS 0.021987f
C2076 VN.n63 VSUBS 0.021987f
C2077 VN.n64 VSUBS 0.021987f
C2078 VN.n65 VSUBS 0.041155f
C2079 VN.n66 VSUBS 0.040774f
C2080 VN.n67 VSUBS 0.031112f
C2081 VN.n68 VSUBS 0.035481f
C2082 VN.n69 VSUBS 1.60738f
.ends

