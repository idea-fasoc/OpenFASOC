* NGSPICE file created from diff_pair_sample_0142.ext - technology: sky130A

.subckt diff_pair_sample_0142 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=3.23
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=3.23
X2 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=5.1402 ps=27.14 w=13.18 l=3.23
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=3.23
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=5.1402 ps=27.14 w=13.18 l=3.23
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=5.1402 ps=27.14 w=13.18 l=3.23
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=0 ps=0 w=13.18 l=3.23
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.1402 pd=27.14 as=5.1402 ps=27.14 w=13.18 l=3.23
R0 B.n745 B.n744 585
R1 B.n308 B.n105 585
R2 B.n307 B.n306 585
R3 B.n305 B.n304 585
R4 B.n303 B.n302 585
R5 B.n301 B.n300 585
R6 B.n299 B.n298 585
R7 B.n297 B.n296 585
R8 B.n295 B.n294 585
R9 B.n293 B.n292 585
R10 B.n291 B.n290 585
R11 B.n289 B.n288 585
R12 B.n287 B.n286 585
R13 B.n285 B.n284 585
R14 B.n283 B.n282 585
R15 B.n281 B.n280 585
R16 B.n279 B.n278 585
R17 B.n277 B.n276 585
R18 B.n275 B.n274 585
R19 B.n273 B.n272 585
R20 B.n271 B.n270 585
R21 B.n269 B.n268 585
R22 B.n267 B.n266 585
R23 B.n265 B.n264 585
R24 B.n263 B.n262 585
R25 B.n261 B.n260 585
R26 B.n259 B.n258 585
R27 B.n257 B.n256 585
R28 B.n255 B.n254 585
R29 B.n253 B.n252 585
R30 B.n251 B.n250 585
R31 B.n249 B.n248 585
R32 B.n247 B.n246 585
R33 B.n245 B.n244 585
R34 B.n243 B.n242 585
R35 B.n241 B.n240 585
R36 B.n239 B.n238 585
R37 B.n237 B.n236 585
R38 B.n235 B.n234 585
R39 B.n233 B.n232 585
R40 B.n231 B.n230 585
R41 B.n229 B.n228 585
R42 B.n227 B.n226 585
R43 B.n225 B.n224 585
R44 B.n223 B.n222 585
R45 B.n220 B.n219 585
R46 B.n218 B.n217 585
R47 B.n216 B.n215 585
R48 B.n214 B.n213 585
R49 B.n212 B.n211 585
R50 B.n210 B.n209 585
R51 B.n208 B.n207 585
R52 B.n206 B.n205 585
R53 B.n204 B.n203 585
R54 B.n202 B.n201 585
R55 B.n199 B.n198 585
R56 B.n197 B.n196 585
R57 B.n195 B.n194 585
R58 B.n193 B.n192 585
R59 B.n191 B.n190 585
R60 B.n189 B.n188 585
R61 B.n187 B.n186 585
R62 B.n185 B.n184 585
R63 B.n183 B.n182 585
R64 B.n181 B.n180 585
R65 B.n179 B.n178 585
R66 B.n177 B.n176 585
R67 B.n175 B.n174 585
R68 B.n173 B.n172 585
R69 B.n171 B.n170 585
R70 B.n169 B.n168 585
R71 B.n167 B.n166 585
R72 B.n165 B.n164 585
R73 B.n163 B.n162 585
R74 B.n161 B.n160 585
R75 B.n159 B.n158 585
R76 B.n157 B.n156 585
R77 B.n155 B.n154 585
R78 B.n153 B.n152 585
R79 B.n151 B.n150 585
R80 B.n149 B.n148 585
R81 B.n147 B.n146 585
R82 B.n145 B.n144 585
R83 B.n143 B.n142 585
R84 B.n141 B.n140 585
R85 B.n139 B.n138 585
R86 B.n137 B.n136 585
R87 B.n135 B.n134 585
R88 B.n133 B.n132 585
R89 B.n131 B.n130 585
R90 B.n129 B.n128 585
R91 B.n127 B.n126 585
R92 B.n125 B.n124 585
R93 B.n123 B.n122 585
R94 B.n121 B.n120 585
R95 B.n119 B.n118 585
R96 B.n117 B.n116 585
R97 B.n115 B.n114 585
R98 B.n113 B.n112 585
R99 B.n111 B.n110 585
R100 B.n743 B.n55 585
R101 B.n748 B.n55 585
R102 B.n742 B.n54 585
R103 B.n749 B.n54 585
R104 B.n741 B.n740 585
R105 B.n740 B.n50 585
R106 B.n739 B.n49 585
R107 B.n755 B.n49 585
R108 B.n738 B.n48 585
R109 B.n756 B.n48 585
R110 B.n737 B.n47 585
R111 B.n757 B.n47 585
R112 B.n736 B.n735 585
R113 B.n735 B.n43 585
R114 B.n734 B.n42 585
R115 B.n763 B.n42 585
R116 B.n733 B.n41 585
R117 B.n764 B.n41 585
R118 B.n732 B.n40 585
R119 B.n765 B.n40 585
R120 B.n731 B.n730 585
R121 B.n730 B.n36 585
R122 B.n729 B.n35 585
R123 B.n771 B.n35 585
R124 B.n728 B.n34 585
R125 B.n772 B.n34 585
R126 B.n727 B.n33 585
R127 B.n773 B.n33 585
R128 B.n726 B.n725 585
R129 B.n725 B.n29 585
R130 B.n724 B.n28 585
R131 B.n779 B.n28 585
R132 B.n723 B.n27 585
R133 B.n780 B.n27 585
R134 B.n722 B.n26 585
R135 B.n781 B.n26 585
R136 B.n721 B.n720 585
R137 B.n720 B.n22 585
R138 B.n719 B.n21 585
R139 B.n787 B.n21 585
R140 B.n718 B.n20 585
R141 B.n788 B.n20 585
R142 B.n717 B.n19 585
R143 B.n789 B.n19 585
R144 B.n716 B.n715 585
R145 B.n715 B.n18 585
R146 B.n714 B.n14 585
R147 B.n795 B.n14 585
R148 B.n713 B.n13 585
R149 B.n796 B.n13 585
R150 B.n712 B.n12 585
R151 B.n797 B.n12 585
R152 B.n711 B.n710 585
R153 B.n710 B.n8 585
R154 B.n709 B.n7 585
R155 B.n803 B.n7 585
R156 B.n708 B.n6 585
R157 B.n804 B.n6 585
R158 B.n707 B.n5 585
R159 B.n805 B.n5 585
R160 B.n706 B.n705 585
R161 B.n705 B.n4 585
R162 B.n704 B.n309 585
R163 B.n704 B.n703 585
R164 B.n694 B.n310 585
R165 B.n311 B.n310 585
R166 B.n696 B.n695 585
R167 B.n697 B.n696 585
R168 B.n693 B.n316 585
R169 B.n316 B.n315 585
R170 B.n692 B.n691 585
R171 B.n691 B.n690 585
R172 B.n318 B.n317 585
R173 B.n683 B.n318 585
R174 B.n682 B.n681 585
R175 B.n684 B.n682 585
R176 B.n680 B.n323 585
R177 B.n323 B.n322 585
R178 B.n679 B.n678 585
R179 B.n678 B.n677 585
R180 B.n325 B.n324 585
R181 B.n326 B.n325 585
R182 B.n670 B.n669 585
R183 B.n671 B.n670 585
R184 B.n668 B.n331 585
R185 B.n331 B.n330 585
R186 B.n667 B.n666 585
R187 B.n666 B.n665 585
R188 B.n333 B.n332 585
R189 B.n334 B.n333 585
R190 B.n658 B.n657 585
R191 B.n659 B.n658 585
R192 B.n656 B.n339 585
R193 B.n339 B.n338 585
R194 B.n655 B.n654 585
R195 B.n654 B.n653 585
R196 B.n341 B.n340 585
R197 B.n342 B.n341 585
R198 B.n646 B.n645 585
R199 B.n647 B.n646 585
R200 B.n644 B.n346 585
R201 B.n350 B.n346 585
R202 B.n643 B.n642 585
R203 B.n642 B.n641 585
R204 B.n348 B.n347 585
R205 B.n349 B.n348 585
R206 B.n634 B.n633 585
R207 B.n635 B.n634 585
R208 B.n632 B.n355 585
R209 B.n355 B.n354 585
R210 B.n631 B.n630 585
R211 B.n630 B.n629 585
R212 B.n357 B.n356 585
R213 B.n358 B.n357 585
R214 B.n622 B.n621 585
R215 B.n623 B.n622 585
R216 B.n620 B.n363 585
R217 B.n363 B.n362 585
R218 B.n615 B.n614 585
R219 B.n613 B.n415 585
R220 B.n612 B.n414 585
R221 B.n617 B.n414 585
R222 B.n611 B.n610 585
R223 B.n609 B.n608 585
R224 B.n607 B.n606 585
R225 B.n605 B.n604 585
R226 B.n603 B.n602 585
R227 B.n601 B.n600 585
R228 B.n599 B.n598 585
R229 B.n597 B.n596 585
R230 B.n595 B.n594 585
R231 B.n593 B.n592 585
R232 B.n591 B.n590 585
R233 B.n589 B.n588 585
R234 B.n587 B.n586 585
R235 B.n585 B.n584 585
R236 B.n583 B.n582 585
R237 B.n581 B.n580 585
R238 B.n579 B.n578 585
R239 B.n577 B.n576 585
R240 B.n575 B.n574 585
R241 B.n573 B.n572 585
R242 B.n571 B.n570 585
R243 B.n569 B.n568 585
R244 B.n567 B.n566 585
R245 B.n565 B.n564 585
R246 B.n563 B.n562 585
R247 B.n561 B.n560 585
R248 B.n559 B.n558 585
R249 B.n557 B.n556 585
R250 B.n555 B.n554 585
R251 B.n553 B.n552 585
R252 B.n551 B.n550 585
R253 B.n549 B.n548 585
R254 B.n547 B.n546 585
R255 B.n545 B.n544 585
R256 B.n543 B.n542 585
R257 B.n541 B.n540 585
R258 B.n539 B.n538 585
R259 B.n537 B.n536 585
R260 B.n535 B.n534 585
R261 B.n533 B.n532 585
R262 B.n531 B.n530 585
R263 B.n529 B.n528 585
R264 B.n527 B.n526 585
R265 B.n525 B.n524 585
R266 B.n523 B.n522 585
R267 B.n521 B.n520 585
R268 B.n519 B.n518 585
R269 B.n517 B.n516 585
R270 B.n515 B.n514 585
R271 B.n513 B.n512 585
R272 B.n511 B.n510 585
R273 B.n509 B.n508 585
R274 B.n507 B.n506 585
R275 B.n505 B.n504 585
R276 B.n503 B.n502 585
R277 B.n501 B.n500 585
R278 B.n499 B.n498 585
R279 B.n497 B.n496 585
R280 B.n495 B.n494 585
R281 B.n493 B.n492 585
R282 B.n491 B.n490 585
R283 B.n489 B.n488 585
R284 B.n487 B.n486 585
R285 B.n485 B.n484 585
R286 B.n483 B.n482 585
R287 B.n481 B.n480 585
R288 B.n479 B.n478 585
R289 B.n477 B.n476 585
R290 B.n475 B.n474 585
R291 B.n473 B.n472 585
R292 B.n471 B.n470 585
R293 B.n469 B.n468 585
R294 B.n467 B.n466 585
R295 B.n465 B.n464 585
R296 B.n463 B.n462 585
R297 B.n461 B.n460 585
R298 B.n459 B.n458 585
R299 B.n457 B.n456 585
R300 B.n455 B.n454 585
R301 B.n453 B.n452 585
R302 B.n451 B.n450 585
R303 B.n449 B.n448 585
R304 B.n447 B.n446 585
R305 B.n445 B.n444 585
R306 B.n443 B.n442 585
R307 B.n441 B.n440 585
R308 B.n439 B.n438 585
R309 B.n437 B.n436 585
R310 B.n435 B.n434 585
R311 B.n433 B.n432 585
R312 B.n431 B.n430 585
R313 B.n429 B.n428 585
R314 B.n427 B.n426 585
R315 B.n425 B.n424 585
R316 B.n423 B.n422 585
R317 B.n365 B.n364 585
R318 B.n619 B.n618 585
R319 B.n618 B.n617 585
R320 B.n361 B.n360 585
R321 B.n362 B.n361 585
R322 B.n625 B.n624 585
R323 B.n624 B.n623 585
R324 B.n626 B.n359 585
R325 B.n359 B.n358 585
R326 B.n628 B.n627 585
R327 B.n629 B.n628 585
R328 B.n353 B.n352 585
R329 B.n354 B.n353 585
R330 B.n637 B.n636 585
R331 B.n636 B.n635 585
R332 B.n638 B.n351 585
R333 B.n351 B.n349 585
R334 B.n640 B.n639 585
R335 B.n641 B.n640 585
R336 B.n345 B.n344 585
R337 B.n350 B.n345 585
R338 B.n649 B.n648 585
R339 B.n648 B.n647 585
R340 B.n650 B.n343 585
R341 B.n343 B.n342 585
R342 B.n652 B.n651 585
R343 B.n653 B.n652 585
R344 B.n337 B.n336 585
R345 B.n338 B.n337 585
R346 B.n661 B.n660 585
R347 B.n660 B.n659 585
R348 B.n662 B.n335 585
R349 B.n335 B.n334 585
R350 B.n664 B.n663 585
R351 B.n665 B.n664 585
R352 B.n329 B.n328 585
R353 B.n330 B.n329 585
R354 B.n673 B.n672 585
R355 B.n672 B.n671 585
R356 B.n674 B.n327 585
R357 B.n327 B.n326 585
R358 B.n676 B.n675 585
R359 B.n677 B.n676 585
R360 B.n321 B.n320 585
R361 B.n322 B.n321 585
R362 B.n686 B.n685 585
R363 B.n685 B.n684 585
R364 B.n687 B.n319 585
R365 B.n683 B.n319 585
R366 B.n689 B.n688 585
R367 B.n690 B.n689 585
R368 B.n314 B.n313 585
R369 B.n315 B.n314 585
R370 B.n699 B.n698 585
R371 B.n698 B.n697 585
R372 B.n700 B.n312 585
R373 B.n312 B.n311 585
R374 B.n702 B.n701 585
R375 B.n703 B.n702 585
R376 B.n2 B.n0 585
R377 B.n4 B.n2 585
R378 B.n3 B.n1 585
R379 B.n804 B.n3 585
R380 B.n802 B.n801 585
R381 B.n803 B.n802 585
R382 B.n800 B.n9 585
R383 B.n9 B.n8 585
R384 B.n799 B.n798 585
R385 B.n798 B.n797 585
R386 B.n11 B.n10 585
R387 B.n796 B.n11 585
R388 B.n794 B.n793 585
R389 B.n795 B.n794 585
R390 B.n792 B.n15 585
R391 B.n18 B.n15 585
R392 B.n791 B.n790 585
R393 B.n790 B.n789 585
R394 B.n17 B.n16 585
R395 B.n788 B.n17 585
R396 B.n786 B.n785 585
R397 B.n787 B.n786 585
R398 B.n784 B.n23 585
R399 B.n23 B.n22 585
R400 B.n783 B.n782 585
R401 B.n782 B.n781 585
R402 B.n25 B.n24 585
R403 B.n780 B.n25 585
R404 B.n778 B.n777 585
R405 B.n779 B.n778 585
R406 B.n776 B.n30 585
R407 B.n30 B.n29 585
R408 B.n775 B.n774 585
R409 B.n774 B.n773 585
R410 B.n32 B.n31 585
R411 B.n772 B.n32 585
R412 B.n770 B.n769 585
R413 B.n771 B.n770 585
R414 B.n768 B.n37 585
R415 B.n37 B.n36 585
R416 B.n767 B.n766 585
R417 B.n766 B.n765 585
R418 B.n39 B.n38 585
R419 B.n764 B.n39 585
R420 B.n762 B.n761 585
R421 B.n763 B.n762 585
R422 B.n760 B.n44 585
R423 B.n44 B.n43 585
R424 B.n759 B.n758 585
R425 B.n758 B.n757 585
R426 B.n46 B.n45 585
R427 B.n756 B.n46 585
R428 B.n754 B.n753 585
R429 B.n755 B.n754 585
R430 B.n752 B.n51 585
R431 B.n51 B.n50 585
R432 B.n751 B.n750 585
R433 B.n750 B.n749 585
R434 B.n53 B.n52 585
R435 B.n748 B.n53 585
R436 B.n807 B.n806 585
R437 B.n806 B.n805 585
R438 B.n615 B.n361 487.695
R439 B.n110 B.n53 487.695
R440 B.n618 B.n363 487.695
R441 B.n745 B.n55 487.695
R442 B.n419 B.t2 307.173
R443 B.n416 B.t10 307.173
R444 B.n108 B.t6 307.173
R445 B.n106 B.t13 307.173
R446 B.n747 B.n746 256.663
R447 B.n747 B.n104 256.663
R448 B.n747 B.n103 256.663
R449 B.n747 B.n102 256.663
R450 B.n747 B.n101 256.663
R451 B.n747 B.n100 256.663
R452 B.n747 B.n99 256.663
R453 B.n747 B.n98 256.663
R454 B.n747 B.n97 256.663
R455 B.n747 B.n96 256.663
R456 B.n747 B.n95 256.663
R457 B.n747 B.n94 256.663
R458 B.n747 B.n93 256.663
R459 B.n747 B.n92 256.663
R460 B.n747 B.n91 256.663
R461 B.n747 B.n90 256.663
R462 B.n747 B.n89 256.663
R463 B.n747 B.n88 256.663
R464 B.n747 B.n87 256.663
R465 B.n747 B.n86 256.663
R466 B.n747 B.n85 256.663
R467 B.n747 B.n84 256.663
R468 B.n747 B.n83 256.663
R469 B.n747 B.n82 256.663
R470 B.n747 B.n81 256.663
R471 B.n747 B.n80 256.663
R472 B.n747 B.n79 256.663
R473 B.n747 B.n78 256.663
R474 B.n747 B.n77 256.663
R475 B.n747 B.n76 256.663
R476 B.n747 B.n75 256.663
R477 B.n747 B.n74 256.663
R478 B.n747 B.n73 256.663
R479 B.n747 B.n72 256.663
R480 B.n747 B.n71 256.663
R481 B.n747 B.n70 256.663
R482 B.n747 B.n69 256.663
R483 B.n747 B.n68 256.663
R484 B.n747 B.n67 256.663
R485 B.n747 B.n66 256.663
R486 B.n747 B.n65 256.663
R487 B.n747 B.n64 256.663
R488 B.n747 B.n63 256.663
R489 B.n747 B.n62 256.663
R490 B.n747 B.n61 256.663
R491 B.n747 B.n60 256.663
R492 B.n747 B.n59 256.663
R493 B.n747 B.n58 256.663
R494 B.n747 B.n57 256.663
R495 B.n747 B.n56 256.663
R496 B.n617 B.n616 256.663
R497 B.n617 B.n366 256.663
R498 B.n617 B.n367 256.663
R499 B.n617 B.n368 256.663
R500 B.n617 B.n369 256.663
R501 B.n617 B.n370 256.663
R502 B.n617 B.n371 256.663
R503 B.n617 B.n372 256.663
R504 B.n617 B.n373 256.663
R505 B.n617 B.n374 256.663
R506 B.n617 B.n375 256.663
R507 B.n617 B.n376 256.663
R508 B.n617 B.n377 256.663
R509 B.n617 B.n378 256.663
R510 B.n617 B.n379 256.663
R511 B.n617 B.n380 256.663
R512 B.n617 B.n381 256.663
R513 B.n617 B.n382 256.663
R514 B.n617 B.n383 256.663
R515 B.n617 B.n384 256.663
R516 B.n617 B.n385 256.663
R517 B.n617 B.n386 256.663
R518 B.n617 B.n387 256.663
R519 B.n617 B.n388 256.663
R520 B.n617 B.n389 256.663
R521 B.n617 B.n390 256.663
R522 B.n617 B.n391 256.663
R523 B.n617 B.n392 256.663
R524 B.n617 B.n393 256.663
R525 B.n617 B.n394 256.663
R526 B.n617 B.n395 256.663
R527 B.n617 B.n396 256.663
R528 B.n617 B.n397 256.663
R529 B.n617 B.n398 256.663
R530 B.n617 B.n399 256.663
R531 B.n617 B.n400 256.663
R532 B.n617 B.n401 256.663
R533 B.n617 B.n402 256.663
R534 B.n617 B.n403 256.663
R535 B.n617 B.n404 256.663
R536 B.n617 B.n405 256.663
R537 B.n617 B.n406 256.663
R538 B.n617 B.n407 256.663
R539 B.n617 B.n408 256.663
R540 B.n617 B.n409 256.663
R541 B.n617 B.n410 256.663
R542 B.n617 B.n411 256.663
R543 B.n617 B.n412 256.663
R544 B.n617 B.n413 256.663
R545 B.n624 B.n361 163.367
R546 B.n624 B.n359 163.367
R547 B.n628 B.n359 163.367
R548 B.n628 B.n353 163.367
R549 B.n636 B.n353 163.367
R550 B.n636 B.n351 163.367
R551 B.n640 B.n351 163.367
R552 B.n640 B.n345 163.367
R553 B.n648 B.n345 163.367
R554 B.n648 B.n343 163.367
R555 B.n652 B.n343 163.367
R556 B.n652 B.n337 163.367
R557 B.n660 B.n337 163.367
R558 B.n660 B.n335 163.367
R559 B.n664 B.n335 163.367
R560 B.n664 B.n329 163.367
R561 B.n672 B.n329 163.367
R562 B.n672 B.n327 163.367
R563 B.n676 B.n327 163.367
R564 B.n676 B.n321 163.367
R565 B.n685 B.n321 163.367
R566 B.n685 B.n319 163.367
R567 B.n689 B.n319 163.367
R568 B.n689 B.n314 163.367
R569 B.n698 B.n314 163.367
R570 B.n698 B.n312 163.367
R571 B.n702 B.n312 163.367
R572 B.n702 B.n2 163.367
R573 B.n806 B.n2 163.367
R574 B.n806 B.n3 163.367
R575 B.n802 B.n3 163.367
R576 B.n802 B.n9 163.367
R577 B.n798 B.n9 163.367
R578 B.n798 B.n11 163.367
R579 B.n794 B.n11 163.367
R580 B.n794 B.n15 163.367
R581 B.n790 B.n15 163.367
R582 B.n790 B.n17 163.367
R583 B.n786 B.n17 163.367
R584 B.n786 B.n23 163.367
R585 B.n782 B.n23 163.367
R586 B.n782 B.n25 163.367
R587 B.n778 B.n25 163.367
R588 B.n778 B.n30 163.367
R589 B.n774 B.n30 163.367
R590 B.n774 B.n32 163.367
R591 B.n770 B.n32 163.367
R592 B.n770 B.n37 163.367
R593 B.n766 B.n37 163.367
R594 B.n766 B.n39 163.367
R595 B.n762 B.n39 163.367
R596 B.n762 B.n44 163.367
R597 B.n758 B.n44 163.367
R598 B.n758 B.n46 163.367
R599 B.n754 B.n46 163.367
R600 B.n754 B.n51 163.367
R601 B.n750 B.n51 163.367
R602 B.n750 B.n53 163.367
R603 B.n415 B.n414 163.367
R604 B.n610 B.n414 163.367
R605 B.n608 B.n607 163.367
R606 B.n604 B.n603 163.367
R607 B.n600 B.n599 163.367
R608 B.n596 B.n595 163.367
R609 B.n592 B.n591 163.367
R610 B.n588 B.n587 163.367
R611 B.n584 B.n583 163.367
R612 B.n580 B.n579 163.367
R613 B.n576 B.n575 163.367
R614 B.n572 B.n571 163.367
R615 B.n568 B.n567 163.367
R616 B.n564 B.n563 163.367
R617 B.n560 B.n559 163.367
R618 B.n556 B.n555 163.367
R619 B.n552 B.n551 163.367
R620 B.n548 B.n547 163.367
R621 B.n544 B.n543 163.367
R622 B.n540 B.n539 163.367
R623 B.n536 B.n535 163.367
R624 B.n532 B.n531 163.367
R625 B.n528 B.n527 163.367
R626 B.n524 B.n523 163.367
R627 B.n520 B.n519 163.367
R628 B.n516 B.n515 163.367
R629 B.n512 B.n511 163.367
R630 B.n508 B.n507 163.367
R631 B.n504 B.n503 163.367
R632 B.n500 B.n499 163.367
R633 B.n496 B.n495 163.367
R634 B.n492 B.n491 163.367
R635 B.n488 B.n487 163.367
R636 B.n484 B.n483 163.367
R637 B.n480 B.n479 163.367
R638 B.n476 B.n475 163.367
R639 B.n472 B.n471 163.367
R640 B.n468 B.n467 163.367
R641 B.n464 B.n463 163.367
R642 B.n460 B.n459 163.367
R643 B.n456 B.n455 163.367
R644 B.n452 B.n451 163.367
R645 B.n448 B.n447 163.367
R646 B.n444 B.n443 163.367
R647 B.n440 B.n439 163.367
R648 B.n436 B.n435 163.367
R649 B.n432 B.n431 163.367
R650 B.n428 B.n427 163.367
R651 B.n424 B.n423 163.367
R652 B.n618 B.n365 163.367
R653 B.n622 B.n363 163.367
R654 B.n622 B.n357 163.367
R655 B.n630 B.n357 163.367
R656 B.n630 B.n355 163.367
R657 B.n634 B.n355 163.367
R658 B.n634 B.n348 163.367
R659 B.n642 B.n348 163.367
R660 B.n642 B.n346 163.367
R661 B.n646 B.n346 163.367
R662 B.n646 B.n341 163.367
R663 B.n654 B.n341 163.367
R664 B.n654 B.n339 163.367
R665 B.n658 B.n339 163.367
R666 B.n658 B.n333 163.367
R667 B.n666 B.n333 163.367
R668 B.n666 B.n331 163.367
R669 B.n670 B.n331 163.367
R670 B.n670 B.n325 163.367
R671 B.n678 B.n325 163.367
R672 B.n678 B.n323 163.367
R673 B.n682 B.n323 163.367
R674 B.n682 B.n318 163.367
R675 B.n691 B.n318 163.367
R676 B.n691 B.n316 163.367
R677 B.n696 B.n316 163.367
R678 B.n696 B.n310 163.367
R679 B.n704 B.n310 163.367
R680 B.n705 B.n704 163.367
R681 B.n705 B.n5 163.367
R682 B.n6 B.n5 163.367
R683 B.n7 B.n6 163.367
R684 B.n710 B.n7 163.367
R685 B.n710 B.n12 163.367
R686 B.n13 B.n12 163.367
R687 B.n14 B.n13 163.367
R688 B.n715 B.n14 163.367
R689 B.n715 B.n19 163.367
R690 B.n20 B.n19 163.367
R691 B.n21 B.n20 163.367
R692 B.n720 B.n21 163.367
R693 B.n720 B.n26 163.367
R694 B.n27 B.n26 163.367
R695 B.n28 B.n27 163.367
R696 B.n725 B.n28 163.367
R697 B.n725 B.n33 163.367
R698 B.n34 B.n33 163.367
R699 B.n35 B.n34 163.367
R700 B.n730 B.n35 163.367
R701 B.n730 B.n40 163.367
R702 B.n41 B.n40 163.367
R703 B.n42 B.n41 163.367
R704 B.n735 B.n42 163.367
R705 B.n735 B.n47 163.367
R706 B.n48 B.n47 163.367
R707 B.n49 B.n48 163.367
R708 B.n740 B.n49 163.367
R709 B.n740 B.n54 163.367
R710 B.n55 B.n54 163.367
R711 B.n114 B.n113 163.367
R712 B.n118 B.n117 163.367
R713 B.n122 B.n121 163.367
R714 B.n126 B.n125 163.367
R715 B.n130 B.n129 163.367
R716 B.n134 B.n133 163.367
R717 B.n138 B.n137 163.367
R718 B.n142 B.n141 163.367
R719 B.n146 B.n145 163.367
R720 B.n150 B.n149 163.367
R721 B.n154 B.n153 163.367
R722 B.n158 B.n157 163.367
R723 B.n162 B.n161 163.367
R724 B.n166 B.n165 163.367
R725 B.n170 B.n169 163.367
R726 B.n174 B.n173 163.367
R727 B.n178 B.n177 163.367
R728 B.n182 B.n181 163.367
R729 B.n186 B.n185 163.367
R730 B.n190 B.n189 163.367
R731 B.n194 B.n193 163.367
R732 B.n198 B.n197 163.367
R733 B.n203 B.n202 163.367
R734 B.n207 B.n206 163.367
R735 B.n211 B.n210 163.367
R736 B.n215 B.n214 163.367
R737 B.n219 B.n218 163.367
R738 B.n224 B.n223 163.367
R739 B.n228 B.n227 163.367
R740 B.n232 B.n231 163.367
R741 B.n236 B.n235 163.367
R742 B.n240 B.n239 163.367
R743 B.n244 B.n243 163.367
R744 B.n248 B.n247 163.367
R745 B.n252 B.n251 163.367
R746 B.n256 B.n255 163.367
R747 B.n260 B.n259 163.367
R748 B.n264 B.n263 163.367
R749 B.n268 B.n267 163.367
R750 B.n272 B.n271 163.367
R751 B.n276 B.n275 163.367
R752 B.n280 B.n279 163.367
R753 B.n284 B.n283 163.367
R754 B.n288 B.n287 163.367
R755 B.n292 B.n291 163.367
R756 B.n296 B.n295 163.367
R757 B.n300 B.n299 163.367
R758 B.n304 B.n303 163.367
R759 B.n306 B.n105 163.367
R760 B.n419 B.t5 141.728
R761 B.n106 B.t14 141.728
R762 B.n416 B.t12 141.712
R763 B.n108 B.t8 141.712
R764 B.n617 B.n362 75.6981
R765 B.n748 B.n747 75.6981
R766 B.n420 B.t4 72.6861
R767 B.n107 B.t15 72.6861
R768 B.n417 B.t11 72.6694
R769 B.n109 B.t9 72.6694
R770 B.n616 B.n615 71.676
R771 B.n610 B.n366 71.676
R772 B.n607 B.n367 71.676
R773 B.n603 B.n368 71.676
R774 B.n599 B.n369 71.676
R775 B.n595 B.n370 71.676
R776 B.n591 B.n371 71.676
R777 B.n587 B.n372 71.676
R778 B.n583 B.n373 71.676
R779 B.n579 B.n374 71.676
R780 B.n575 B.n375 71.676
R781 B.n571 B.n376 71.676
R782 B.n567 B.n377 71.676
R783 B.n563 B.n378 71.676
R784 B.n559 B.n379 71.676
R785 B.n555 B.n380 71.676
R786 B.n551 B.n381 71.676
R787 B.n547 B.n382 71.676
R788 B.n543 B.n383 71.676
R789 B.n539 B.n384 71.676
R790 B.n535 B.n385 71.676
R791 B.n531 B.n386 71.676
R792 B.n527 B.n387 71.676
R793 B.n523 B.n388 71.676
R794 B.n519 B.n389 71.676
R795 B.n515 B.n390 71.676
R796 B.n511 B.n391 71.676
R797 B.n507 B.n392 71.676
R798 B.n503 B.n393 71.676
R799 B.n499 B.n394 71.676
R800 B.n495 B.n395 71.676
R801 B.n491 B.n396 71.676
R802 B.n487 B.n397 71.676
R803 B.n483 B.n398 71.676
R804 B.n479 B.n399 71.676
R805 B.n475 B.n400 71.676
R806 B.n471 B.n401 71.676
R807 B.n467 B.n402 71.676
R808 B.n463 B.n403 71.676
R809 B.n459 B.n404 71.676
R810 B.n455 B.n405 71.676
R811 B.n451 B.n406 71.676
R812 B.n447 B.n407 71.676
R813 B.n443 B.n408 71.676
R814 B.n439 B.n409 71.676
R815 B.n435 B.n410 71.676
R816 B.n431 B.n411 71.676
R817 B.n427 B.n412 71.676
R818 B.n423 B.n413 71.676
R819 B.n110 B.n56 71.676
R820 B.n114 B.n57 71.676
R821 B.n118 B.n58 71.676
R822 B.n122 B.n59 71.676
R823 B.n126 B.n60 71.676
R824 B.n130 B.n61 71.676
R825 B.n134 B.n62 71.676
R826 B.n138 B.n63 71.676
R827 B.n142 B.n64 71.676
R828 B.n146 B.n65 71.676
R829 B.n150 B.n66 71.676
R830 B.n154 B.n67 71.676
R831 B.n158 B.n68 71.676
R832 B.n162 B.n69 71.676
R833 B.n166 B.n70 71.676
R834 B.n170 B.n71 71.676
R835 B.n174 B.n72 71.676
R836 B.n178 B.n73 71.676
R837 B.n182 B.n74 71.676
R838 B.n186 B.n75 71.676
R839 B.n190 B.n76 71.676
R840 B.n194 B.n77 71.676
R841 B.n198 B.n78 71.676
R842 B.n203 B.n79 71.676
R843 B.n207 B.n80 71.676
R844 B.n211 B.n81 71.676
R845 B.n215 B.n82 71.676
R846 B.n219 B.n83 71.676
R847 B.n224 B.n84 71.676
R848 B.n228 B.n85 71.676
R849 B.n232 B.n86 71.676
R850 B.n236 B.n87 71.676
R851 B.n240 B.n88 71.676
R852 B.n244 B.n89 71.676
R853 B.n248 B.n90 71.676
R854 B.n252 B.n91 71.676
R855 B.n256 B.n92 71.676
R856 B.n260 B.n93 71.676
R857 B.n264 B.n94 71.676
R858 B.n268 B.n95 71.676
R859 B.n272 B.n96 71.676
R860 B.n276 B.n97 71.676
R861 B.n280 B.n98 71.676
R862 B.n284 B.n99 71.676
R863 B.n288 B.n100 71.676
R864 B.n292 B.n101 71.676
R865 B.n296 B.n102 71.676
R866 B.n300 B.n103 71.676
R867 B.n304 B.n104 71.676
R868 B.n746 B.n105 71.676
R869 B.n746 B.n745 71.676
R870 B.n306 B.n104 71.676
R871 B.n303 B.n103 71.676
R872 B.n299 B.n102 71.676
R873 B.n295 B.n101 71.676
R874 B.n291 B.n100 71.676
R875 B.n287 B.n99 71.676
R876 B.n283 B.n98 71.676
R877 B.n279 B.n97 71.676
R878 B.n275 B.n96 71.676
R879 B.n271 B.n95 71.676
R880 B.n267 B.n94 71.676
R881 B.n263 B.n93 71.676
R882 B.n259 B.n92 71.676
R883 B.n255 B.n91 71.676
R884 B.n251 B.n90 71.676
R885 B.n247 B.n89 71.676
R886 B.n243 B.n88 71.676
R887 B.n239 B.n87 71.676
R888 B.n235 B.n86 71.676
R889 B.n231 B.n85 71.676
R890 B.n227 B.n84 71.676
R891 B.n223 B.n83 71.676
R892 B.n218 B.n82 71.676
R893 B.n214 B.n81 71.676
R894 B.n210 B.n80 71.676
R895 B.n206 B.n79 71.676
R896 B.n202 B.n78 71.676
R897 B.n197 B.n77 71.676
R898 B.n193 B.n76 71.676
R899 B.n189 B.n75 71.676
R900 B.n185 B.n74 71.676
R901 B.n181 B.n73 71.676
R902 B.n177 B.n72 71.676
R903 B.n173 B.n71 71.676
R904 B.n169 B.n70 71.676
R905 B.n165 B.n69 71.676
R906 B.n161 B.n68 71.676
R907 B.n157 B.n67 71.676
R908 B.n153 B.n66 71.676
R909 B.n149 B.n65 71.676
R910 B.n145 B.n64 71.676
R911 B.n141 B.n63 71.676
R912 B.n137 B.n62 71.676
R913 B.n133 B.n61 71.676
R914 B.n129 B.n60 71.676
R915 B.n125 B.n59 71.676
R916 B.n121 B.n58 71.676
R917 B.n117 B.n57 71.676
R918 B.n113 B.n56 71.676
R919 B.n616 B.n415 71.676
R920 B.n608 B.n366 71.676
R921 B.n604 B.n367 71.676
R922 B.n600 B.n368 71.676
R923 B.n596 B.n369 71.676
R924 B.n592 B.n370 71.676
R925 B.n588 B.n371 71.676
R926 B.n584 B.n372 71.676
R927 B.n580 B.n373 71.676
R928 B.n576 B.n374 71.676
R929 B.n572 B.n375 71.676
R930 B.n568 B.n376 71.676
R931 B.n564 B.n377 71.676
R932 B.n560 B.n378 71.676
R933 B.n556 B.n379 71.676
R934 B.n552 B.n380 71.676
R935 B.n548 B.n381 71.676
R936 B.n544 B.n382 71.676
R937 B.n540 B.n383 71.676
R938 B.n536 B.n384 71.676
R939 B.n532 B.n385 71.676
R940 B.n528 B.n386 71.676
R941 B.n524 B.n387 71.676
R942 B.n520 B.n388 71.676
R943 B.n516 B.n389 71.676
R944 B.n512 B.n390 71.676
R945 B.n508 B.n391 71.676
R946 B.n504 B.n392 71.676
R947 B.n500 B.n393 71.676
R948 B.n496 B.n394 71.676
R949 B.n492 B.n395 71.676
R950 B.n488 B.n396 71.676
R951 B.n484 B.n397 71.676
R952 B.n480 B.n398 71.676
R953 B.n476 B.n399 71.676
R954 B.n472 B.n400 71.676
R955 B.n468 B.n401 71.676
R956 B.n464 B.n402 71.676
R957 B.n460 B.n403 71.676
R958 B.n456 B.n404 71.676
R959 B.n452 B.n405 71.676
R960 B.n448 B.n406 71.676
R961 B.n444 B.n407 71.676
R962 B.n440 B.n408 71.676
R963 B.n436 B.n409 71.676
R964 B.n432 B.n410 71.676
R965 B.n428 B.n411 71.676
R966 B.n424 B.n412 71.676
R967 B.n413 B.n365 71.676
R968 B.n420 B.n419 69.0429
R969 B.n417 B.n416 69.0429
R970 B.n109 B.n108 69.0429
R971 B.n107 B.n106 69.0429
R972 B.n421 B.n420 59.5399
R973 B.n418 B.n417 59.5399
R974 B.n200 B.n109 59.5399
R975 B.n221 B.n107 59.5399
R976 B.n623 B.n362 40.5315
R977 B.n623 B.n358 40.5315
R978 B.n629 B.n358 40.5315
R979 B.n629 B.n354 40.5315
R980 B.n635 B.n354 40.5315
R981 B.n635 B.n349 40.5315
R982 B.n641 B.n349 40.5315
R983 B.n641 B.n350 40.5315
R984 B.n647 B.n342 40.5315
R985 B.n653 B.n342 40.5315
R986 B.n653 B.n338 40.5315
R987 B.n659 B.n338 40.5315
R988 B.n659 B.n334 40.5315
R989 B.n665 B.n334 40.5315
R990 B.n665 B.n330 40.5315
R991 B.n671 B.n330 40.5315
R992 B.n671 B.n326 40.5315
R993 B.n677 B.n326 40.5315
R994 B.n677 B.n322 40.5315
R995 B.n684 B.n322 40.5315
R996 B.n684 B.n683 40.5315
R997 B.n690 B.n315 40.5315
R998 B.n697 B.n315 40.5315
R999 B.n697 B.n311 40.5315
R1000 B.n703 B.n311 40.5315
R1001 B.n703 B.n4 40.5315
R1002 B.n805 B.n4 40.5315
R1003 B.n805 B.n804 40.5315
R1004 B.n804 B.n803 40.5315
R1005 B.n803 B.n8 40.5315
R1006 B.n797 B.n8 40.5315
R1007 B.n797 B.n796 40.5315
R1008 B.n796 B.n795 40.5315
R1009 B.n789 B.n18 40.5315
R1010 B.n789 B.n788 40.5315
R1011 B.n788 B.n787 40.5315
R1012 B.n787 B.n22 40.5315
R1013 B.n781 B.n22 40.5315
R1014 B.n781 B.n780 40.5315
R1015 B.n780 B.n779 40.5315
R1016 B.n779 B.n29 40.5315
R1017 B.n773 B.n29 40.5315
R1018 B.n773 B.n772 40.5315
R1019 B.n772 B.n771 40.5315
R1020 B.n771 B.n36 40.5315
R1021 B.n765 B.n36 40.5315
R1022 B.n764 B.n763 40.5315
R1023 B.n763 B.n43 40.5315
R1024 B.n757 B.n43 40.5315
R1025 B.n757 B.n756 40.5315
R1026 B.n756 B.n755 40.5315
R1027 B.n755 B.n50 40.5315
R1028 B.n749 B.n50 40.5315
R1029 B.n749 B.n748 40.5315
R1030 B.n690 B.t0 33.975
R1031 B.n795 B.t1 33.975
R1032 B.n111 B.n52 31.6883
R1033 B.n744 B.n743 31.6883
R1034 B.n620 B.n619 31.6883
R1035 B.n614 B.n360 31.6883
R1036 B.n647 B.t3 20.8621
R1037 B.n765 B.t7 20.8621
R1038 B.n350 B.t3 19.67
R1039 B.t7 B.n764 19.67
R1040 B B.n807 18.0485
R1041 B.n112 B.n111 10.6151
R1042 B.n115 B.n112 10.6151
R1043 B.n116 B.n115 10.6151
R1044 B.n119 B.n116 10.6151
R1045 B.n120 B.n119 10.6151
R1046 B.n123 B.n120 10.6151
R1047 B.n124 B.n123 10.6151
R1048 B.n127 B.n124 10.6151
R1049 B.n128 B.n127 10.6151
R1050 B.n131 B.n128 10.6151
R1051 B.n132 B.n131 10.6151
R1052 B.n135 B.n132 10.6151
R1053 B.n136 B.n135 10.6151
R1054 B.n139 B.n136 10.6151
R1055 B.n140 B.n139 10.6151
R1056 B.n143 B.n140 10.6151
R1057 B.n144 B.n143 10.6151
R1058 B.n147 B.n144 10.6151
R1059 B.n148 B.n147 10.6151
R1060 B.n151 B.n148 10.6151
R1061 B.n152 B.n151 10.6151
R1062 B.n155 B.n152 10.6151
R1063 B.n156 B.n155 10.6151
R1064 B.n159 B.n156 10.6151
R1065 B.n160 B.n159 10.6151
R1066 B.n163 B.n160 10.6151
R1067 B.n164 B.n163 10.6151
R1068 B.n167 B.n164 10.6151
R1069 B.n168 B.n167 10.6151
R1070 B.n171 B.n168 10.6151
R1071 B.n172 B.n171 10.6151
R1072 B.n175 B.n172 10.6151
R1073 B.n176 B.n175 10.6151
R1074 B.n179 B.n176 10.6151
R1075 B.n180 B.n179 10.6151
R1076 B.n183 B.n180 10.6151
R1077 B.n184 B.n183 10.6151
R1078 B.n187 B.n184 10.6151
R1079 B.n188 B.n187 10.6151
R1080 B.n191 B.n188 10.6151
R1081 B.n192 B.n191 10.6151
R1082 B.n195 B.n192 10.6151
R1083 B.n196 B.n195 10.6151
R1084 B.n199 B.n196 10.6151
R1085 B.n204 B.n201 10.6151
R1086 B.n205 B.n204 10.6151
R1087 B.n208 B.n205 10.6151
R1088 B.n209 B.n208 10.6151
R1089 B.n212 B.n209 10.6151
R1090 B.n213 B.n212 10.6151
R1091 B.n216 B.n213 10.6151
R1092 B.n217 B.n216 10.6151
R1093 B.n220 B.n217 10.6151
R1094 B.n225 B.n222 10.6151
R1095 B.n226 B.n225 10.6151
R1096 B.n229 B.n226 10.6151
R1097 B.n230 B.n229 10.6151
R1098 B.n233 B.n230 10.6151
R1099 B.n234 B.n233 10.6151
R1100 B.n237 B.n234 10.6151
R1101 B.n238 B.n237 10.6151
R1102 B.n241 B.n238 10.6151
R1103 B.n242 B.n241 10.6151
R1104 B.n245 B.n242 10.6151
R1105 B.n246 B.n245 10.6151
R1106 B.n249 B.n246 10.6151
R1107 B.n250 B.n249 10.6151
R1108 B.n253 B.n250 10.6151
R1109 B.n254 B.n253 10.6151
R1110 B.n257 B.n254 10.6151
R1111 B.n258 B.n257 10.6151
R1112 B.n261 B.n258 10.6151
R1113 B.n262 B.n261 10.6151
R1114 B.n265 B.n262 10.6151
R1115 B.n266 B.n265 10.6151
R1116 B.n269 B.n266 10.6151
R1117 B.n270 B.n269 10.6151
R1118 B.n273 B.n270 10.6151
R1119 B.n274 B.n273 10.6151
R1120 B.n277 B.n274 10.6151
R1121 B.n278 B.n277 10.6151
R1122 B.n281 B.n278 10.6151
R1123 B.n282 B.n281 10.6151
R1124 B.n285 B.n282 10.6151
R1125 B.n286 B.n285 10.6151
R1126 B.n289 B.n286 10.6151
R1127 B.n290 B.n289 10.6151
R1128 B.n293 B.n290 10.6151
R1129 B.n294 B.n293 10.6151
R1130 B.n297 B.n294 10.6151
R1131 B.n298 B.n297 10.6151
R1132 B.n301 B.n298 10.6151
R1133 B.n302 B.n301 10.6151
R1134 B.n305 B.n302 10.6151
R1135 B.n307 B.n305 10.6151
R1136 B.n308 B.n307 10.6151
R1137 B.n744 B.n308 10.6151
R1138 B.n621 B.n620 10.6151
R1139 B.n621 B.n356 10.6151
R1140 B.n631 B.n356 10.6151
R1141 B.n632 B.n631 10.6151
R1142 B.n633 B.n632 10.6151
R1143 B.n633 B.n347 10.6151
R1144 B.n643 B.n347 10.6151
R1145 B.n644 B.n643 10.6151
R1146 B.n645 B.n644 10.6151
R1147 B.n645 B.n340 10.6151
R1148 B.n655 B.n340 10.6151
R1149 B.n656 B.n655 10.6151
R1150 B.n657 B.n656 10.6151
R1151 B.n657 B.n332 10.6151
R1152 B.n667 B.n332 10.6151
R1153 B.n668 B.n667 10.6151
R1154 B.n669 B.n668 10.6151
R1155 B.n669 B.n324 10.6151
R1156 B.n679 B.n324 10.6151
R1157 B.n680 B.n679 10.6151
R1158 B.n681 B.n680 10.6151
R1159 B.n681 B.n317 10.6151
R1160 B.n692 B.n317 10.6151
R1161 B.n693 B.n692 10.6151
R1162 B.n695 B.n693 10.6151
R1163 B.n695 B.n694 10.6151
R1164 B.n694 B.n309 10.6151
R1165 B.n706 B.n309 10.6151
R1166 B.n707 B.n706 10.6151
R1167 B.n708 B.n707 10.6151
R1168 B.n709 B.n708 10.6151
R1169 B.n711 B.n709 10.6151
R1170 B.n712 B.n711 10.6151
R1171 B.n713 B.n712 10.6151
R1172 B.n714 B.n713 10.6151
R1173 B.n716 B.n714 10.6151
R1174 B.n717 B.n716 10.6151
R1175 B.n718 B.n717 10.6151
R1176 B.n719 B.n718 10.6151
R1177 B.n721 B.n719 10.6151
R1178 B.n722 B.n721 10.6151
R1179 B.n723 B.n722 10.6151
R1180 B.n724 B.n723 10.6151
R1181 B.n726 B.n724 10.6151
R1182 B.n727 B.n726 10.6151
R1183 B.n728 B.n727 10.6151
R1184 B.n729 B.n728 10.6151
R1185 B.n731 B.n729 10.6151
R1186 B.n732 B.n731 10.6151
R1187 B.n733 B.n732 10.6151
R1188 B.n734 B.n733 10.6151
R1189 B.n736 B.n734 10.6151
R1190 B.n737 B.n736 10.6151
R1191 B.n738 B.n737 10.6151
R1192 B.n739 B.n738 10.6151
R1193 B.n741 B.n739 10.6151
R1194 B.n742 B.n741 10.6151
R1195 B.n743 B.n742 10.6151
R1196 B.n614 B.n613 10.6151
R1197 B.n613 B.n612 10.6151
R1198 B.n612 B.n611 10.6151
R1199 B.n611 B.n609 10.6151
R1200 B.n609 B.n606 10.6151
R1201 B.n606 B.n605 10.6151
R1202 B.n605 B.n602 10.6151
R1203 B.n602 B.n601 10.6151
R1204 B.n601 B.n598 10.6151
R1205 B.n598 B.n597 10.6151
R1206 B.n597 B.n594 10.6151
R1207 B.n594 B.n593 10.6151
R1208 B.n593 B.n590 10.6151
R1209 B.n590 B.n589 10.6151
R1210 B.n589 B.n586 10.6151
R1211 B.n586 B.n585 10.6151
R1212 B.n585 B.n582 10.6151
R1213 B.n582 B.n581 10.6151
R1214 B.n581 B.n578 10.6151
R1215 B.n578 B.n577 10.6151
R1216 B.n577 B.n574 10.6151
R1217 B.n574 B.n573 10.6151
R1218 B.n573 B.n570 10.6151
R1219 B.n570 B.n569 10.6151
R1220 B.n569 B.n566 10.6151
R1221 B.n566 B.n565 10.6151
R1222 B.n565 B.n562 10.6151
R1223 B.n562 B.n561 10.6151
R1224 B.n561 B.n558 10.6151
R1225 B.n558 B.n557 10.6151
R1226 B.n557 B.n554 10.6151
R1227 B.n554 B.n553 10.6151
R1228 B.n553 B.n550 10.6151
R1229 B.n550 B.n549 10.6151
R1230 B.n549 B.n546 10.6151
R1231 B.n546 B.n545 10.6151
R1232 B.n545 B.n542 10.6151
R1233 B.n542 B.n541 10.6151
R1234 B.n541 B.n538 10.6151
R1235 B.n538 B.n537 10.6151
R1236 B.n537 B.n534 10.6151
R1237 B.n534 B.n533 10.6151
R1238 B.n533 B.n530 10.6151
R1239 B.n530 B.n529 10.6151
R1240 B.n526 B.n525 10.6151
R1241 B.n525 B.n522 10.6151
R1242 B.n522 B.n521 10.6151
R1243 B.n521 B.n518 10.6151
R1244 B.n518 B.n517 10.6151
R1245 B.n517 B.n514 10.6151
R1246 B.n514 B.n513 10.6151
R1247 B.n513 B.n510 10.6151
R1248 B.n510 B.n509 10.6151
R1249 B.n506 B.n505 10.6151
R1250 B.n505 B.n502 10.6151
R1251 B.n502 B.n501 10.6151
R1252 B.n501 B.n498 10.6151
R1253 B.n498 B.n497 10.6151
R1254 B.n497 B.n494 10.6151
R1255 B.n494 B.n493 10.6151
R1256 B.n493 B.n490 10.6151
R1257 B.n490 B.n489 10.6151
R1258 B.n489 B.n486 10.6151
R1259 B.n486 B.n485 10.6151
R1260 B.n485 B.n482 10.6151
R1261 B.n482 B.n481 10.6151
R1262 B.n481 B.n478 10.6151
R1263 B.n478 B.n477 10.6151
R1264 B.n477 B.n474 10.6151
R1265 B.n474 B.n473 10.6151
R1266 B.n473 B.n470 10.6151
R1267 B.n470 B.n469 10.6151
R1268 B.n469 B.n466 10.6151
R1269 B.n466 B.n465 10.6151
R1270 B.n465 B.n462 10.6151
R1271 B.n462 B.n461 10.6151
R1272 B.n461 B.n458 10.6151
R1273 B.n458 B.n457 10.6151
R1274 B.n457 B.n454 10.6151
R1275 B.n454 B.n453 10.6151
R1276 B.n453 B.n450 10.6151
R1277 B.n450 B.n449 10.6151
R1278 B.n449 B.n446 10.6151
R1279 B.n446 B.n445 10.6151
R1280 B.n445 B.n442 10.6151
R1281 B.n442 B.n441 10.6151
R1282 B.n441 B.n438 10.6151
R1283 B.n438 B.n437 10.6151
R1284 B.n437 B.n434 10.6151
R1285 B.n434 B.n433 10.6151
R1286 B.n433 B.n430 10.6151
R1287 B.n430 B.n429 10.6151
R1288 B.n429 B.n426 10.6151
R1289 B.n426 B.n425 10.6151
R1290 B.n425 B.n422 10.6151
R1291 B.n422 B.n364 10.6151
R1292 B.n619 B.n364 10.6151
R1293 B.n625 B.n360 10.6151
R1294 B.n626 B.n625 10.6151
R1295 B.n627 B.n626 10.6151
R1296 B.n627 B.n352 10.6151
R1297 B.n637 B.n352 10.6151
R1298 B.n638 B.n637 10.6151
R1299 B.n639 B.n638 10.6151
R1300 B.n639 B.n344 10.6151
R1301 B.n649 B.n344 10.6151
R1302 B.n650 B.n649 10.6151
R1303 B.n651 B.n650 10.6151
R1304 B.n651 B.n336 10.6151
R1305 B.n661 B.n336 10.6151
R1306 B.n662 B.n661 10.6151
R1307 B.n663 B.n662 10.6151
R1308 B.n663 B.n328 10.6151
R1309 B.n673 B.n328 10.6151
R1310 B.n674 B.n673 10.6151
R1311 B.n675 B.n674 10.6151
R1312 B.n675 B.n320 10.6151
R1313 B.n686 B.n320 10.6151
R1314 B.n687 B.n686 10.6151
R1315 B.n688 B.n687 10.6151
R1316 B.n688 B.n313 10.6151
R1317 B.n699 B.n313 10.6151
R1318 B.n700 B.n699 10.6151
R1319 B.n701 B.n700 10.6151
R1320 B.n701 B.n0 10.6151
R1321 B.n801 B.n1 10.6151
R1322 B.n801 B.n800 10.6151
R1323 B.n800 B.n799 10.6151
R1324 B.n799 B.n10 10.6151
R1325 B.n793 B.n10 10.6151
R1326 B.n793 B.n792 10.6151
R1327 B.n792 B.n791 10.6151
R1328 B.n791 B.n16 10.6151
R1329 B.n785 B.n16 10.6151
R1330 B.n785 B.n784 10.6151
R1331 B.n784 B.n783 10.6151
R1332 B.n783 B.n24 10.6151
R1333 B.n777 B.n24 10.6151
R1334 B.n777 B.n776 10.6151
R1335 B.n776 B.n775 10.6151
R1336 B.n775 B.n31 10.6151
R1337 B.n769 B.n31 10.6151
R1338 B.n769 B.n768 10.6151
R1339 B.n768 B.n767 10.6151
R1340 B.n767 B.n38 10.6151
R1341 B.n761 B.n38 10.6151
R1342 B.n761 B.n760 10.6151
R1343 B.n760 B.n759 10.6151
R1344 B.n759 B.n45 10.6151
R1345 B.n753 B.n45 10.6151
R1346 B.n753 B.n752 10.6151
R1347 B.n752 B.n751 10.6151
R1348 B.n751 B.n52 10.6151
R1349 B.n200 B.n199 9.36635
R1350 B.n222 B.n221 9.36635
R1351 B.n529 B.n418 9.36635
R1352 B.n506 B.n421 9.36635
R1353 B.n683 B.t0 6.55699
R1354 B.n18 B.t1 6.55699
R1355 B.n807 B.n0 2.81026
R1356 B.n807 B.n1 2.81026
R1357 B.n201 B.n200 1.24928
R1358 B.n221 B.n220 1.24928
R1359 B.n526 B.n418 1.24928
R1360 B.n509 B.n421 1.24928
R1361 VN VN.t1 184.315
R1362 VN VN.t0 137.712
R1363 VTAIL.n1 VTAIL.t2 46.0609
R1364 VTAIL.n3 VTAIL.t1 46.0607
R1365 VTAIL.n0 VTAIL.t0 46.0607
R1366 VTAIL.n2 VTAIL.t3 46.0607
R1367 VTAIL.n1 VTAIL.n0 29.8669
R1368 VTAIL.n3 VTAIL.n2 26.7979
R1369 VTAIL.n2 VTAIL.n1 2.00481
R1370 VTAIL VTAIL.n0 1.29576
R1371 VTAIL VTAIL.n3 0.709552
R1372 VDD2.n0 VDD2.t1 103.898
R1373 VDD2.n0 VDD2.t0 62.7395
R1374 VDD2 VDD2.n0 0.825931
R1375 VP.n0 VP.t1 184.407
R1376 VP.n0 VP.t0 137.186
R1377 VP VP.n0 0.526373
R1378 VDD1 VDD1.t1 105.191
R1379 VDD1 VDD1.t0 63.5649
C0 VDD2 VP 0.359943f
C1 VDD1 VN 0.148745f
C2 VDD2 VN 3.12216f
C3 VDD1 VTAIL 5.4804f
C4 VDD2 VTAIL 5.53559f
C5 VN VP 5.96953f
C6 VDD2 VDD1 0.751439f
C7 VTAIL VP 2.79107f
C8 VTAIL VN 2.77681f
C9 VDD1 VP 3.33093f
C10 VDD2 B 4.860137f
C11 VDD1 B 8.20104f
C12 VTAIL B 8.1496f
C13 VN B 11.63024f
C14 VP B 7.271983f
C15 VDD1.t0 B 2.4351f
C16 VDD1.t1 B 3.09123f
C17 VP.t1 B 4.18209f
C18 VP.t0 B 3.54271f
C19 VP.n0 B 4.28209f
C20 VDD2.t1 B 3.00566f
C21 VDD2.t0 B 2.39665f
C22 VDD2.n0 B 3.04402f
C23 VTAIL.t0 B 2.38614f
C24 VTAIL.n0 B 1.819f
C25 VTAIL.t2 B 2.38614f
C26 VTAIL.n1 B 1.86636f
C27 VTAIL.t3 B 2.38614f
C28 VTAIL.n2 B 1.66136f
C29 VTAIL.t1 B 2.38614f
C30 VTAIL.n3 B 1.57483f
C31 VN.t0 B 3.47733f
C32 VN.t1 B 4.09991f
.ends

