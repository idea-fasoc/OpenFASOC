* NGSPICE file created from diff_pair_sample_1538.ext - technology: sky130A

.subckt diff_pair_sample_1538 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=0 ps=0 w=8.69 l=2.93
X1 VDD1.t5 VP.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=1.43385 ps=9.02 w=8.69 l=2.93
X2 VDD1.t4 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=1.43385 ps=9.02 w=8.69 l=2.93
X3 VDD2.t5 VN.t0 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=1.43385 ps=9.02 w=8.69 l=2.93
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=0 ps=0 w=8.69 l=2.93
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=0 ps=0 w=8.69 l=2.93
X6 VTAIL.t7 VP.t2 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=1.43385 ps=9.02 w=8.69 l=2.93
X7 VTAIL.t8 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=1.43385 ps=9.02 w=8.69 l=2.93
X8 VDD2.t4 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=1.43385 ps=9.02 w=8.69 l=2.93
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=3.3891 ps=18.16 w=8.69 l=2.93
X10 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=3.3891 ps=18.16 w=8.69 l=2.93
X11 VDD1.t1 VP.t4 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=3.3891 ps=18.16 w=8.69 l=2.93
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3891 pd=18.16 as=0 ps=0 w=8.69 l=2.93
X13 VDD1.t0 VP.t5 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=3.3891 ps=18.16 w=8.69 l=2.93
X14 VTAIL.t4 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=1.43385 ps=9.02 w=8.69 l=2.93
X15 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.43385 pd=9.02 as=1.43385 ps=9.02 w=8.69 l=2.93
R0 B.n604 B.n127 585
R1 B.n127 B.n86 585
R2 B.n606 B.n605 585
R3 B.n608 B.n126 585
R4 B.n611 B.n610 585
R5 B.n612 B.n125 585
R6 B.n614 B.n613 585
R7 B.n616 B.n124 585
R8 B.n619 B.n618 585
R9 B.n620 B.n123 585
R10 B.n622 B.n621 585
R11 B.n624 B.n122 585
R12 B.n627 B.n626 585
R13 B.n628 B.n121 585
R14 B.n630 B.n629 585
R15 B.n632 B.n120 585
R16 B.n635 B.n634 585
R17 B.n636 B.n119 585
R18 B.n638 B.n637 585
R19 B.n640 B.n118 585
R20 B.n643 B.n642 585
R21 B.n644 B.n117 585
R22 B.n646 B.n645 585
R23 B.n648 B.n116 585
R24 B.n651 B.n650 585
R25 B.n652 B.n115 585
R26 B.n654 B.n653 585
R27 B.n656 B.n114 585
R28 B.n659 B.n658 585
R29 B.n660 B.n113 585
R30 B.n662 B.n661 585
R31 B.n664 B.n112 585
R32 B.n667 B.n666 585
R33 B.n669 B.n109 585
R34 B.n671 B.n670 585
R35 B.n673 B.n108 585
R36 B.n676 B.n675 585
R37 B.n677 B.n107 585
R38 B.n679 B.n678 585
R39 B.n681 B.n106 585
R40 B.n684 B.n683 585
R41 B.n685 B.n103 585
R42 B.n688 B.n687 585
R43 B.n690 B.n102 585
R44 B.n693 B.n692 585
R45 B.n694 B.n101 585
R46 B.n696 B.n695 585
R47 B.n698 B.n100 585
R48 B.n701 B.n700 585
R49 B.n702 B.n99 585
R50 B.n704 B.n703 585
R51 B.n706 B.n98 585
R52 B.n709 B.n708 585
R53 B.n710 B.n97 585
R54 B.n712 B.n711 585
R55 B.n714 B.n96 585
R56 B.n717 B.n716 585
R57 B.n718 B.n95 585
R58 B.n720 B.n719 585
R59 B.n722 B.n94 585
R60 B.n725 B.n724 585
R61 B.n726 B.n93 585
R62 B.n728 B.n727 585
R63 B.n730 B.n92 585
R64 B.n733 B.n732 585
R65 B.n734 B.n91 585
R66 B.n736 B.n735 585
R67 B.n738 B.n90 585
R68 B.n741 B.n740 585
R69 B.n742 B.n89 585
R70 B.n744 B.n743 585
R71 B.n746 B.n88 585
R72 B.n749 B.n748 585
R73 B.n750 B.n87 585
R74 B.n603 B.n85 585
R75 B.n753 B.n85 585
R76 B.n602 B.n84 585
R77 B.n754 B.n84 585
R78 B.n601 B.n83 585
R79 B.n755 B.n83 585
R80 B.n600 B.n599 585
R81 B.n599 B.n79 585
R82 B.n598 B.n78 585
R83 B.n761 B.n78 585
R84 B.n597 B.n77 585
R85 B.n762 B.n77 585
R86 B.n596 B.n76 585
R87 B.n763 B.n76 585
R88 B.n595 B.n594 585
R89 B.n594 B.n72 585
R90 B.n593 B.n71 585
R91 B.n769 B.n71 585
R92 B.n592 B.n70 585
R93 B.n770 B.n70 585
R94 B.n591 B.n69 585
R95 B.n771 B.n69 585
R96 B.n590 B.n589 585
R97 B.n589 B.n65 585
R98 B.n588 B.n64 585
R99 B.n777 B.n64 585
R100 B.n587 B.n63 585
R101 B.n778 B.n63 585
R102 B.n586 B.n62 585
R103 B.n779 B.n62 585
R104 B.n585 B.n584 585
R105 B.n584 B.n58 585
R106 B.n583 B.n57 585
R107 B.n785 B.n57 585
R108 B.n582 B.n56 585
R109 B.n786 B.n56 585
R110 B.n581 B.n55 585
R111 B.n787 B.n55 585
R112 B.n580 B.n579 585
R113 B.n579 B.n51 585
R114 B.n578 B.n50 585
R115 B.n793 B.n50 585
R116 B.n577 B.n49 585
R117 B.n794 B.n49 585
R118 B.n576 B.n48 585
R119 B.n795 B.n48 585
R120 B.n575 B.n574 585
R121 B.n574 B.n44 585
R122 B.n573 B.n43 585
R123 B.n801 B.n43 585
R124 B.n572 B.n42 585
R125 B.n802 B.n42 585
R126 B.n571 B.n41 585
R127 B.n803 B.n41 585
R128 B.n570 B.n569 585
R129 B.n569 B.n37 585
R130 B.n568 B.n36 585
R131 B.n809 B.n36 585
R132 B.n567 B.n35 585
R133 B.n810 B.n35 585
R134 B.n566 B.n34 585
R135 B.n811 B.n34 585
R136 B.n565 B.n564 585
R137 B.n564 B.n30 585
R138 B.n563 B.n29 585
R139 B.n817 B.n29 585
R140 B.n562 B.n28 585
R141 B.n818 B.n28 585
R142 B.n561 B.n27 585
R143 B.n819 B.n27 585
R144 B.n560 B.n559 585
R145 B.n559 B.n23 585
R146 B.n558 B.n22 585
R147 B.n825 B.n22 585
R148 B.n557 B.n21 585
R149 B.n826 B.n21 585
R150 B.n556 B.n20 585
R151 B.n827 B.n20 585
R152 B.n555 B.n554 585
R153 B.n554 B.n16 585
R154 B.n553 B.n15 585
R155 B.n833 B.n15 585
R156 B.n552 B.n14 585
R157 B.n834 B.n14 585
R158 B.n551 B.n13 585
R159 B.n835 B.n13 585
R160 B.n550 B.n549 585
R161 B.n549 B.n12 585
R162 B.n548 B.n547 585
R163 B.n548 B.n8 585
R164 B.n546 B.n7 585
R165 B.n842 B.n7 585
R166 B.n545 B.n6 585
R167 B.n843 B.n6 585
R168 B.n544 B.n5 585
R169 B.n844 B.n5 585
R170 B.n543 B.n542 585
R171 B.n542 B.n4 585
R172 B.n541 B.n128 585
R173 B.n541 B.n540 585
R174 B.n531 B.n129 585
R175 B.n130 B.n129 585
R176 B.n533 B.n532 585
R177 B.n534 B.n533 585
R178 B.n530 B.n135 585
R179 B.n135 B.n134 585
R180 B.n529 B.n528 585
R181 B.n528 B.n527 585
R182 B.n137 B.n136 585
R183 B.n138 B.n137 585
R184 B.n520 B.n519 585
R185 B.n521 B.n520 585
R186 B.n518 B.n143 585
R187 B.n143 B.n142 585
R188 B.n517 B.n516 585
R189 B.n516 B.n515 585
R190 B.n145 B.n144 585
R191 B.n146 B.n145 585
R192 B.n508 B.n507 585
R193 B.n509 B.n508 585
R194 B.n506 B.n151 585
R195 B.n151 B.n150 585
R196 B.n505 B.n504 585
R197 B.n504 B.n503 585
R198 B.n153 B.n152 585
R199 B.n154 B.n153 585
R200 B.n496 B.n495 585
R201 B.n497 B.n496 585
R202 B.n494 B.n159 585
R203 B.n159 B.n158 585
R204 B.n493 B.n492 585
R205 B.n492 B.n491 585
R206 B.n161 B.n160 585
R207 B.n162 B.n161 585
R208 B.n484 B.n483 585
R209 B.n485 B.n484 585
R210 B.n482 B.n167 585
R211 B.n167 B.n166 585
R212 B.n481 B.n480 585
R213 B.n480 B.n479 585
R214 B.n169 B.n168 585
R215 B.n170 B.n169 585
R216 B.n472 B.n471 585
R217 B.n473 B.n472 585
R218 B.n470 B.n175 585
R219 B.n175 B.n174 585
R220 B.n469 B.n468 585
R221 B.n468 B.n467 585
R222 B.n177 B.n176 585
R223 B.n178 B.n177 585
R224 B.n460 B.n459 585
R225 B.n461 B.n460 585
R226 B.n458 B.n183 585
R227 B.n183 B.n182 585
R228 B.n457 B.n456 585
R229 B.n456 B.n455 585
R230 B.n185 B.n184 585
R231 B.n186 B.n185 585
R232 B.n448 B.n447 585
R233 B.n449 B.n448 585
R234 B.n446 B.n191 585
R235 B.n191 B.n190 585
R236 B.n445 B.n444 585
R237 B.n444 B.n443 585
R238 B.n193 B.n192 585
R239 B.n194 B.n193 585
R240 B.n436 B.n435 585
R241 B.n437 B.n436 585
R242 B.n434 B.n199 585
R243 B.n199 B.n198 585
R244 B.n433 B.n432 585
R245 B.n432 B.n431 585
R246 B.n201 B.n200 585
R247 B.n202 B.n201 585
R248 B.n424 B.n423 585
R249 B.n425 B.n424 585
R250 B.n422 B.n207 585
R251 B.n207 B.n206 585
R252 B.n421 B.n420 585
R253 B.n420 B.n419 585
R254 B.n209 B.n208 585
R255 B.n210 B.n209 585
R256 B.n412 B.n411 585
R257 B.n413 B.n412 585
R258 B.n410 B.n215 585
R259 B.n215 B.n214 585
R260 B.n409 B.n408 585
R261 B.n408 B.n407 585
R262 B.n404 B.n219 585
R263 B.n403 B.n402 585
R264 B.n400 B.n220 585
R265 B.n400 B.n218 585
R266 B.n399 B.n398 585
R267 B.n397 B.n396 585
R268 B.n395 B.n222 585
R269 B.n393 B.n392 585
R270 B.n391 B.n223 585
R271 B.n390 B.n389 585
R272 B.n387 B.n224 585
R273 B.n385 B.n384 585
R274 B.n383 B.n225 585
R275 B.n382 B.n381 585
R276 B.n379 B.n226 585
R277 B.n377 B.n376 585
R278 B.n375 B.n227 585
R279 B.n374 B.n373 585
R280 B.n371 B.n228 585
R281 B.n369 B.n368 585
R282 B.n367 B.n229 585
R283 B.n366 B.n365 585
R284 B.n363 B.n230 585
R285 B.n361 B.n360 585
R286 B.n359 B.n231 585
R287 B.n358 B.n357 585
R288 B.n355 B.n232 585
R289 B.n353 B.n352 585
R290 B.n351 B.n233 585
R291 B.n350 B.n349 585
R292 B.n347 B.n234 585
R293 B.n345 B.n344 585
R294 B.n343 B.n235 585
R295 B.n341 B.n340 585
R296 B.n338 B.n238 585
R297 B.n336 B.n335 585
R298 B.n334 B.n239 585
R299 B.n333 B.n332 585
R300 B.n330 B.n240 585
R301 B.n328 B.n327 585
R302 B.n326 B.n241 585
R303 B.n325 B.n324 585
R304 B.n322 B.n321 585
R305 B.n320 B.n319 585
R306 B.n318 B.n246 585
R307 B.n316 B.n315 585
R308 B.n314 B.n247 585
R309 B.n313 B.n312 585
R310 B.n310 B.n248 585
R311 B.n308 B.n307 585
R312 B.n306 B.n249 585
R313 B.n305 B.n304 585
R314 B.n302 B.n250 585
R315 B.n300 B.n299 585
R316 B.n298 B.n251 585
R317 B.n297 B.n296 585
R318 B.n294 B.n252 585
R319 B.n292 B.n291 585
R320 B.n290 B.n253 585
R321 B.n289 B.n288 585
R322 B.n286 B.n254 585
R323 B.n284 B.n283 585
R324 B.n282 B.n255 585
R325 B.n281 B.n280 585
R326 B.n278 B.n256 585
R327 B.n276 B.n275 585
R328 B.n274 B.n257 585
R329 B.n273 B.n272 585
R330 B.n270 B.n258 585
R331 B.n268 B.n267 585
R332 B.n266 B.n259 585
R333 B.n265 B.n264 585
R334 B.n262 B.n260 585
R335 B.n217 B.n216 585
R336 B.n406 B.n405 585
R337 B.n407 B.n406 585
R338 B.n213 B.n212 585
R339 B.n214 B.n213 585
R340 B.n415 B.n414 585
R341 B.n414 B.n413 585
R342 B.n416 B.n211 585
R343 B.n211 B.n210 585
R344 B.n418 B.n417 585
R345 B.n419 B.n418 585
R346 B.n205 B.n204 585
R347 B.n206 B.n205 585
R348 B.n427 B.n426 585
R349 B.n426 B.n425 585
R350 B.n428 B.n203 585
R351 B.n203 B.n202 585
R352 B.n430 B.n429 585
R353 B.n431 B.n430 585
R354 B.n197 B.n196 585
R355 B.n198 B.n197 585
R356 B.n439 B.n438 585
R357 B.n438 B.n437 585
R358 B.n440 B.n195 585
R359 B.n195 B.n194 585
R360 B.n442 B.n441 585
R361 B.n443 B.n442 585
R362 B.n189 B.n188 585
R363 B.n190 B.n189 585
R364 B.n451 B.n450 585
R365 B.n450 B.n449 585
R366 B.n452 B.n187 585
R367 B.n187 B.n186 585
R368 B.n454 B.n453 585
R369 B.n455 B.n454 585
R370 B.n181 B.n180 585
R371 B.n182 B.n181 585
R372 B.n463 B.n462 585
R373 B.n462 B.n461 585
R374 B.n464 B.n179 585
R375 B.n179 B.n178 585
R376 B.n466 B.n465 585
R377 B.n467 B.n466 585
R378 B.n173 B.n172 585
R379 B.n174 B.n173 585
R380 B.n475 B.n474 585
R381 B.n474 B.n473 585
R382 B.n476 B.n171 585
R383 B.n171 B.n170 585
R384 B.n478 B.n477 585
R385 B.n479 B.n478 585
R386 B.n165 B.n164 585
R387 B.n166 B.n165 585
R388 B.n487 B.n486 585
R389 B.n486 B.n485 585
R390 B.n488 B.n163 585
R391 B.n163 B.n162 585
R392 B.n490 B.n489 585
R393 B.n491 B.n490 585
R394 B.n157 B.n156 585
R395 B.n158 B.n157 585
R396 B.n499 B.n498 585
R397 B.n498 B.n497 585
R398 B.n500 B.n155 585
R399 B.n155 B.n154 585
R400 B.n502 B.n501 585
R401 B.n503 B.n502 585
R402 B.n149 B.n148 585
R403 B.n150 B.n149 585
R404 B.n511 B.n510 585
R405 B.n510 B.n509 585
R406 B.n512 B.n147 585
R407 B.n147 B.n146 585
R408 B.n514 B.n513 585
R409 B.n515 B.n514 585
R410 B.n141 B.n140 585
R411 B.n142 B.n141 585
R412 B.n523 B.n522 585
R413 B.n522 B.n521 585
R414 B.n524 B.n139 585
R415 B.n139 B.n138 585
R416 B.n526 B.n525 585
R417 B.n527 B.n526 585
R418 B.n133 B.n132 585
R419 B.n134 B.n133 585
R420 B.n536 B.n535 585
R421 B.n535 B.n534 585
R422 B.n537 B.n131 585
R423 B.n131 B.n130 585
R424 B.n539 B.n538 585
R425 B.n540 B.n539 585
R426 B.n3 B.n0 585
R427 B.n4 B.n3 585
R428 B.n841 B.n1 585
R429 B.n842 B.n841 585
R430 B.n840 B.n839 585
R431 B.n840 B.n8 585
R432 B.n838 B.n9 585
R433 B.n12 B.n9 585
R434 B.n837 B.n836 585
R435 B.n836 B.n835 585
R436 B.n11 B.n10 585
R437 B.n834 B.n11 585
R438 B.n832 B.n831 585
R439 B.n833 B.n832 585
R440 B.n830 B.n17 585
R441 B.n17 B.n16 585
R442 B.n829 B.n828 585
R443 B.n828 B.n827 585
R444 B.n19 B.n18 585
R445 B.n826 B.n19 585
R446 B.n824 B.n823 585
R447 B.n825 B.n824 585
R448 B.n822 B.n24 585
R449 B.n24 B.n23 585
R450 B.n821 B.n820 585
R451 B.n820 B.n819 585
R452 B.n26 B.n25 585
R453 B.n818 B.n26 585
R454 B.n816 B.n815 585
R455 B.n817 B.n816 585
R456 B.n814 B.n31 585
R457 B.n31 B.n30 585
R458 B.n813 B.n812 585
R459 B.n812 B.n811 585
R460 B.n33 B.n32 585
R461 B.n810 B.n33 585
R462 B.n808 B.n807 585
R463 B.n809 B.n808 585
R464 B.n806 B.n38 585
R465 B.n38 B.n37 585
R466 B.n805 B.n804 585
R467 B.n804 B.n803 585
R468 B.n40 B.n39 585
R469 B.n802 B.n40 585
R470 B.n800 B.n799 585
R471 B.n801 B.n800 585
R472 B.n798 B.n45 585
R473 B.n45 B.n44 585
R474 B.n797 B.n796 585
R475 B.n796 B.n795 585
R476 B.n47 B.n46 585
R477 B.n794 B.n47 585
R478 B.n792 B.n791 585
R479 B.n793 B.n792 585
R480 B.n790 B.n52 585
R481 B.n52 B.n51 585
R482 B.n789 B.n788 585
R483 B.n788 B.n787 585
R484 B.n54 B.n53 585
R485 B.n786 B.n54 585
R486 B.n784 B.n783 585
R487 B.n785 B.n784 585
R488 B.n782 B.n59 585
R489 B.n59 B.n58 585
R490 B.n781 B.n780 585
R491 B.n780 B.n779 585
R492 B.n61 B.n60 585
R493 B.n778 B.n61 585
R494 B.n776 B.n775 585
R495 B.n777 B.n776 585
R496 B.n774 B.n66 585
R497 B.n66 B.n65 585
R498 B.n773 B.n772 585
R499 B.n772 B.n771 585
R500 B.n68 B.n67 585
R501 B.n770 B.n68 585
R502 B.n768 B.n767 585
R503 B.n769 B.n768 585
R504 B.n766 B.n73 585
R505 B.n73 B.n72 585
R506 B.n765 B.n764 585
R507 B.n764 B.n763 585
R508 B.n75 B.n74 585
R509 B.n762 B.n75 585
R510 B.n760 B.n759 585
R511 B.n761 B.n760 585
R512 B.n758 B.n80 585
R513 B.n80 B.n79 585
R514 B.n757 B.n756 585
R515 B.n756 B.n755 585
R516 B.n82 B.n81 585
R517 B.n754 B.n82 585
R518 B.n752 B.n751 585
R519 B.n753 B.n752 585
R520 B.n845 B.n844 585
R521 B.n843 B.n2 585
R522 B.n752 B.n87 521.33
R523 B.n127 B.n85 521.33
R524 B.n408 B.n217 521.33
R525 B.n406 B.n219 521.33
R526 B.n110 B.t11 288.418
R527 B.n242 B.t19 288.418
R528 B.n104 B.t8 288.418
R529 B.n236 B.t16 288.418
R530 B.n104 B.t6 279.974
R531 B.n110 B.t10 279.974
R532 B.n242 B.t17 279.974
R533 B.n236 B.t13 279.974
R534 B.n607 B.n86 256.663
R535 B.n609 B.n86 256.663
R536 B.n615 B.n86 256.663
R537 B.n617 B.n86 256.663
R538 B.n623 B.n86 256.663
R539 B.n625 B.n86 256.663
R540 B.n631 B.n86 256.663
R541 B.n633 B.n86 256.663
R542 B.n639 B.n86 256.663
R543 B.n641 B.n86 256.663
R544 B.n647 B.n86 256.663
R545 B.n649 B.n86 256.663
R546 B.n655 B.n86 256.663
R547 B.n657 B.n86 256.663
R548 B.n663 B.n86 256.663
R549 B.n665 B.n86 256.663
R550 B.n672 B.n86 256.663
R551 B.n674 B.n86 256.663
R552 B.n680 B.n86 256.663
R553 B.n682 B.n86 256.663
R554 B.n689 B.n86 256.663
R555 B.n691 B.n86 256.663
R556 B.n697 B.n86 256.663
R557 B.n699 B.n86 256.663
R558 B.n705 B.n86 256.663
R559 B.n707 B.n86 256.663
R560 B.n713 B.n86 256.663
R561 B.n715 B.n86 256.663
R562 B.n721 B.n86 256.663
R563 B.n723 B.n86 256.663
R564 B.n729 B.n86 256.663
R565 B.n731 B.n86 256.663
R566 B.n737 B.n86 256.663
R567 B.n739 B.n86 256.663
R568 B.n745 B.n86 256.663
R569 B.n747 B.n86 256.663
R570 B.n401 B.n218 256.663
R571 B.n221 B.n218 256.663
R572 B.n394 B.n218 256.663
R573 B.n388 B.n218 256.663
R574 B.n386 B.n218 256.663
R575 B.n380 B.n218 256.663
R576 B.n378 B.n218 256.663
R577 B.n372 B.n218 256.663
R578 B.n370 B.n218 256.663
R579 B.n364 B.n218 256.663
R580 B.n362 B.n218 256.663
R581 B.n356 B.n218 256.663
R582 B.n354 B.n218 256.663
R583 B.n348 B.n218 256.663
R584 B.n346 B.n218 256.663
R585 B.n339 B.n218 256.663
R586 B.n337 B.n218 256.663
R587 B.n331 B.n218 256.663
R588 B.n329 B.n218 256.663
R589 B.n323 B.n218 256.663
R590 B.n245 B.n218 256.663
R591 B.n317 B.n218 256.663
R592 B.n311 B.n218 256.663
R593 B.n309 B.n218 256.663
R594 B.n303 B.n218 256.663
R595 B.n301 B.n218 256.663
R596 B.n295 B.n218 256.663
R597 B.n293 B.n218 256.663
R598 B.n287 B.n218 256.663
R599 B.n285 B.n218 256.663
R600 B.n279 B.n218 256.663
R601 B.n277 B.n218 256.663
R602 B.n271 B.n218 256.663
R603 B.n269 B.n218 256.663
R604 B.n263 B.n218 256.663
R605 B.n261 B.n218 256.663
R606 B.n847 B.n846 256.663
R607 B.n111 B.t12 225.195
R608 B.n243 B.t18 225.195
R609 B.n105 B.t9 225.195
R610 B.n237 B.t15 225.195
R611 B.n748 B.n746 163.367
R612 B.n744 B.n89 163.367
R613 B.n740 B.n738 163.367
R614 B.n736 B.n91 163.367
R615 B.n732 B.n730 163.367
R616 B.n728 B.n93 163.367
R617 B.n724 B.n722 163.367
R618 B.n720 B.n95 163.367
R619 B.n716 B.n714 163.367
R620 B.n712 B.n97 163.367
R621 B.n708 B.n706 163.367
R622 B.n704 B.n99 163.367
R623 B.n700 B.n698 163.367
R624 B.n696 B.n101 163.367
R625 B.n692 B.n690 163.367
R626 B.n688 B.n103 163.367
R627 B.n683 B.n681 163.367
R628 B.n679 B.n107 163.367
R629 B.n675 B.n673 163.367
R630 B.n671 B.n109 163.367
R631 B.n666 B.n664 163.367
R632 B.n662 B.n113 163.367
R633 B.n658 B.n656 163.367
R634 B.n654 B.n115 163.367
R635 B.n650 B.n648 163.367
R636 B.n646 B.n117 163.367
R637 B.n642 B.n640 163.367
R638 B.n638 B.n119 163.367
R639 B.n634 B.n632 163.367
R640 B.n630 B.n121 163.367
R641 B.n626 B.n624 163.367
R642 B.n622 B.n123 163.367
R643 B.n618 B.n616 163.367
R644 B.n614 B.n125 163.367
R645 B.n610 B.n608 163.367
R646 B.n606 B.n127 163.367
R647 B.n408 B.n215 163.367
R648 B.n412 B.n215 163.367
R649 B.n412 B.n209 163.367
R650 B.n420 B.n209 163.367
R651 B.n420 B.n207 163.367
R652 B.n424 B.n207 163.367
R653 B.n424 B.n201 163.367
R654 B.n432 B.n201 163.367
R655 B.n432 B.n199 163.367
R656 B.n436 B.n199 163.367
R657 B.n436 B.n193 163.367
R658 B.n444 B.n193 163.367
R659 B.n444 B.n191 163.367
R660 B.n448 B.n191 163.367
R661 B.n448 B.n185 163.367
R662 B.n456 B.n185 163.367
R663 B.n456 B.n183 163.367
R664 B.n460 B.n183 163.367
R665 B.n460 B.n177 163.367
R666 B.n468 B.n177 163.367
R667 B.n468 B.n175 163.367
R668 B.n472 B.n175 163.367
R669 B.n472 B.n169 163.367
R670 B.n480 B.n169 163.367
R671 B.n480 B.n167 163.367
R672 B.n484 B.n167 163.367
R673 B.n484 B.n161 163.367
R674 B.n492 B.n161 163.367
R675 B.n492 B.n159 163.367
R676 B.n496 B.n159 163.367
R677 B.n496 B.n153 163.367
R678 B.n504 B.n153 163.367
R679 B.n504 B.n151 163.367
R680 B.n508 B.n151 163.367
R681 B.n508 B.n145 163.367
R682 B.n516 B.n145 163.367
R683 B.n516 B.n143 163.367
R684 B.n520 B.n143 163.367
R685 B.n520 B.n137 163.367
R686 B.n528 B.n137 163.367
R687 B.n528 B.n135 163.367
R688 B.n533 B.n135 163.367
R689 B.n533 B.n129 163.367
R690 B.n541 B.n129 163.367
R691 B.n542 B.n541 163.367
R692 B.n542 B.n5 163.367
R693 B.n6 B.n5 163.367
R694 B.n7 B.n6 163.367
R695 B.n548 B.n7 163.367
R696 B.n549 B.n548 163.367
R697 B.n549 B.n13 163.367
R698 B.n14 B.n13 163.367
R699 B.n15 B.n14 163.367
R700 B.n554 B.n15 163.367
R701 B.n554 B.n20 163.367
R702 B.n21 B.n20 163.367
R703 B.n22 B.n21 163.367
R704 B.n559 B.n22 163.367
R705 B.n559 B.n27 163.367
R706 B.n28 B.n27 163.367
R707 B.n29 B.n28 163.367
R708 B.n564 B.n29 163.367
R709 B.n564 B.n34 163.367
R710 B.n35 B.n34 163.367
R711 B.n36 B.n35 163.367
R712 B.n569 B.n36 163.367
R713 B.n569 B.n41 163.367
R714 B.n42 B.n41 163.367
R715 B.n43 B.n42 163.367
R716 B.n574 B.n43 163.367
R717 B.n574 B.n48 163.367
R718 B.n49 B.n48 163.367
R719 B.n50 B.n49 163.367
R720 B.n579 B.n50 163.367
R721 B.n579 B.n55 163.367
R722 B.n56 B.n55 163.367
R723 B.n57 B.n56 163.367
R724 B.n584 B.n57 163.367
R725 B.n584 B.n62 163.367
R726 B.n63 B.n62 163.367
R727 B.n64 B.n63 163.367
R728 B.n589 B.n64 163.367
R729 B.n589 B.n69 163.367
R730 B.n70 B.n69 163.367
R731 B.n71 B.n70 163.367
R732 B.n594 B.n71 163.367
R733 B.n594 B.n76 163.367
R734 B.n77 B.n76 163.367
R735 B.n78 B.n77 163.367
R736 B.n599 B.n78 163.367
R737 B.n599 B.n83 163.367
R738 B.n84 B.n83 163.367
R739 B.n85 B.n84 163.367
R740 B.n402 B.n400 163.367
R741 B.n400 B.n399 163.367
R742 B.n396 B.n395 163.367
R743 B.n393 B.n223 163.367
R744 B.n389 B.n387 163.367
R745 B.n385 B.n225 163.367
R746 B.n381 B.n379 163.367
R747 B.n377 B.n227 163.367
R748 B.n373 B.n371 163.367
R749 B.n369 B.n229 163.367
R750 B.n365 B.n363 163.367
R751 B.n361 B.n231 163.367
R752 B.n357 B.n355 163.367
R753 B.n353 B.n233 163.367
R754 B.n349 B.n347 163.367
R755 B.n345 B.n235 163.367
R756 B.n340 B.n338 163.367
R757 B.n336 B.n239 163.367
R758 B.n332 B.n330 163.367
R759 B.n328 B.n241 163.367
R760 B.n324 B.n322 163.367
R761 B.n319 B.n318 163.367
R762 B.n316 B.n247 163.367
R763 B.n312 B.n310 163.367
R764 B.n308 B.n249 163.367
R765 B.n304 B.n302 163.367
R766 B.n300 B.n251 163.367
R767 B.n296 B.n294 163.367
R768 B.n292 B.n253 163.367
R769 B.n288 B.n286 163.367
R770 B.n284 B.n255 163.367
R771 B.n280 B.n278 163.367
R772 B.n276 B.n257 163.367
R773 B.n272 B.n270 163.367
R774 B.n268 B.n259 163.367
R775 B.n264 B.n262 163.367
R776 B.n406 B.n213 163.367
R777 B.n414 B.n213 163.367
R778 B.n414 B.n211 163.367
R779 B.n418 B.n211 163.367
R780 B.n418 B.n205 163.367
R781 B.n426 B.n205 163.367
R782 B.n426 B.n203 163.367
R783 B.n430 B.n203 163.367
R784 B.n430 B.n197 163.367
R785 B.n438 B.n197 163.367
R786 B.n438 B.n195 163.367
R787 B.n442 B.n195 163.367
R788 B.n442 B.n189 163.367
R789 B.n450 B.n189 163.367
R790 B.n450 B.n187 163.367
R791 B.n454 B.n187 163.367
R792 B.n454 B.n181 163.367
R793 B.n462 B.n181 163.367
R794 B.n462 B.n179 163.367
R795 B.n466 B.n179 163.367
R796 B.n466 B.n173 163.367
R797 B.n474 B.n173 163.367
R798 B.n474 B.n171 163.367
R799 B.n478 B.n171 163.367
R800 B.n478 B.n165 163.367
R801 B.n486 B.n165 163.367
R802 B.n486 B.n163 163.367
R803 B.n490 B.n163 163.367
R804 B.n490 B.n157 163.367
R805 B.n498 B.n157 163.367
R806 B.n498 B.n155 163.367
R807 B.n502 B.n155 163.367
R808 B.n502 B.n149 163.367
R809 B.n510 B.n149 163.367
R810 B.n510 B.n147 163.367
R811 B.n514 B.n147 163.367
R812 B.n514 B.n141 163.367
R813 B.n522 B.n141 163.367
R814 B.n522 B.n139 163.367
R815 B.n526 B.n139 163.367
R816 B.n526 B.n133 163.367
R817 B.n535 B.n133 163.367
R818 B.n535 B.n131 163.367
R819 B.n539 B.n131 163.367
R820 B.n539 B.n3 163.367
R821 B.n845 B.n3 163.367
R822 B.n841 B.n2 163.367
R823 B.n841 B.n840 163.367
R824 B.n840 B.n9 163.367
R825 B.n836 B.n9 163.367
R826 B.n836 B.n11 163.367
R827 B.n832 B.n11 163.367
R828 B.n832 B.n17 163.367
R829 B.n828 B.n17 163.367
R830 B.n828 B.n19 163.367
R831 B.n824 B.n19 163.367
R832 B.n824 B.n24 163.367
R833 B.n820 B.n24 163.367
R834 B.n820 B.n26 163.367
R835 B.n816 B.n26 163.367
R836 B.n816 B.n31 163.367
R837 B.n812 B.n31 163.367
R838 B.n812 B.n33 163.367
R839 B.n808 B.n33 163.367
R840 B.n808 B.n38 163.367
R841 B.n804 B.n38 163.367
R842 B.n804 B.n40 163.367
R843 B.n800 B.n40 163.367
R844 B.n800 B.n45 163.367
R845 B.n796 B.n45 163.367
R846 B.n796 B.n47 163.367
R847 B.n792 B.n47 163.367
R848 B.n792 B.n52 163.367
R849 B.n788 B.n52 163.367
R850 B.n788 B.n54 163.367
R851 B.n784 B.n54 163.367
R852 B.n784 B.n59 163.367
R853 B.n780 B.n59 163.367
R854 B.n780 B.n61 163.367
R855 B.n776 B.n61 163.367
R856 B.n776 B.n66 163.367
R857 B.n772 B.n66 163.367
R858 B.n772 B.n68 163.367
R859 B.n768 B.n68 163.367
R860 B.n768 B.n73 163.367
R861 B.n764 B.n73 163.367
R862 B.n764 B.n75 163.367
R863 B.n760 B.n75 163.367
R864 B.n760 B.n80 163.367
R865 B.n756 B.n80 163.367
R866 B.n756 B.n82 163.367
R867 B.n752 B.n82 163.367
R868 B.n407 B.n218 95.3102
R869 B.n753 B.n86 95.3102
R870 B.n747 B.n87 71.676
R871 B.n746 B.n745 71.676
R872 B.n739 B.n89 71.676
R873 B.n738 B.n737 71.676
R874 B.n731 B.n91 71.676
R875 B.n730 B.n729 71.676
R876 B.n723 B.n93 71.676
R877 B.n722 B.n721 71.676
R878 B.n715 B.n95 71.676
R879 B.n714 B.n713 71.676
R880 B.n707 B.n97 71.676
R881 B.n706 B.n705 71.676
R882 B.n699 B.n99 71.676
R883 B.n698 B.n697 71.676
R884 B.n691 B.n101 71.676
R885 B.n690 B.n689 71.676
R886 B.n682 B.n103 71.676
R887 B.n681 B.n680 71.676
R888 B.n674 B.n107 71.676
R889 B.n673 B.n672 71.676
R890 B.n665 B.n109 71.676
R891 B.n664 B.n663 71.676
R892 B.n657 B.n113 71.676
R893 B.n656 B.n655 71.676
R894 B.n649 B.n115 71.676
R895 B.n648 B.n647 71.676
R896 B.n641 B.n117 71.676
R897 B.n640 B.n639 71.676
R898 B.n633 B.n119 71.676
R899 B.n632 B.n631 71.676
R900 B.n625 B.n121 71.676
R901 B.n624 B.n623 71.676
R902 B.n617 B.n123 71.676
R903 B.n616 B.n615 71.676
R904 B.n609 B.n125 71.676
R905 B.n608 B.n607 71.676
R906 B.n607 B.n606 71.676
R907 B.n610 B.n609 71.676
R908 B.n615 B.n614 71.676
R909 B.n618 B.n617 71.676
R910 B.n623 B.n622 71.676
R911 B.n626 B.n625 71.676
R912 B.n631 B.n630 71.676
R913 B.n634 B.n633 71.676
R914 B.n639 B.n638 71.676
R915 B.n642 B.n641 71.676
R916 B.n647 B.n646 71.676
R917 B.n650 B.n649 71.676
R918 B.n655 B.n654 71.676
R919 B.n658 B.n657 71.676
R920 B.n663 B.n662 71.676
R921 B.n666 B.n665 71.676
R922 B.n672 B.n671 71.676
R923 B.n675 B.n674 71.676
R924 B.n680 B.n679 71.676
R925 B.n683 B.n682 71.676
R926 B.n689 B.n688 71.676
R927 B.n692 B.n691 71.676
R928 B.n697 B.n696 71.676
R929 B.n700 B.n699 71.676
R930 B.n705 B.n704 71.676
R931 B.n708 B.n707 71.676
R932 B.n713 B.n712 71.676
R933 B.n716 B.n715 71.676
R934 B.n721 B.n720 71.676
R935 B.n724 B.n723 71.676
R936 B.n729 B.n728 71.676
R937 B.n732 B.n731 71.676
R938 B.n737 B.n736 71.676
R939 B.n740 B.n739 71.676
R940 B.n745 B.n744 71.676
R941 B.n748 B.n747 71.676
R942 B.n401 B.n219 71.676
R943 B.n399 B.n221 71.676
R944 B.n395 B.n394 71.676
R945 B.n388 B.n223 71.676
R946 B.n387 B.n386 71.676
R947 B.n380 B.n225 71.676
R948 B.n379 B.n378 71.676
R949 B.n372 B.n227 71.676
R950 B.n371 B.n370 71.676
R951 B.n364 B.n229 71.676
R952 B.n363 B.n362 71.676
R953 B.n356 B.n231 71.676
R954 B.n355 B.n354 71.676
R955 B.n348 B.n233 71.676
R956 B.n347 B.n346 71.676
R957 B.n339 B.n235 71.676
R958 B.n338 B.n337 71.676
R959 B.n331 B.n239 71.676
R960 B.n330 B.n329 71.676
R961 B.n323 B.n241 71.676
R962 B.n322 B.n245 71.676
R963 B.n318 B.n317 71.676
R964 B.n311 B.n247 71.676
R965 B.n310 B.n309 71.676
R966 B.n303 B.n249 71.676
R967 B.n302 B.n301 71.676
R968 B.n295 B.n251 71.676
R969 B.n294 B.n293 71.676
R970 B.n287 B.n253 71.676
R971 B.n286 B.n285 71.676
R972 B.n279 B.n255 71.676
R973 B.n278 B.n277 71.676
R974 B.n271 B.n257 71.676
R975 B.n270 B.n269 71.676
R976 B.n263 B.n259 71.676
R977 B.n262 B.n261 71.676
R978 B.n402 B.n401 71.676
R979 B.n396 B.n221 71.676
R980 B.n394 B.n393 71.676
R981 B.n389 B.n388 71.676
R982 B.n386 B.n385 71.676
R983 B.n381 B.n380 71.676
R984 B.n378 B.n377 71.676
R985 B.n373 B.n372 71.676
R986 B.n370 B.n369 71.676
R987 B.n365 B.n364 71.676
R988 B.n362 B.n361 71.676
R989 B.n357 B.n356 71.676
R990 B.n354 B.n353 71.676
R991 B.n349 B.n348 71.676
R992 B.n346 B.n345 71.676
R993 B.n340 B.n339 71.676
R994 B.n337 B.n336 71.676
R995 B.n332 B.n331 71.676
R996 B.n329 B.n328 71.676
R997 B.n324 B.n323 71.676
R998 B.n319 B.n245 71.676
R999 B.n317 B.n316 71.676
R1000 B.n312 B.n311 71.676
R1001 B.n309 B.n308 71.676
R1002 B.n304 B.n303 71.676
R1003 B.n301 B.n300 71.676
R1004 B.n296 B.n295 71.676
R1005 B.n293 B.n292 71.676
R1006 B.n288 B.n287 71.676
R1007 B.n285 B.n284 71.676
R1008 B.n280 B.n279 71.676
R1009 B.n277 B.n276 71.676
R1010 B.n272 B.n271 71.676
R1011 B.n269 B.n268 71.676
R1012 B.n264 B.n263 71.676
R1013 B.n261 B.n217 71.676
R1014 B.n846 B.n845 71.676
R1015 B.n846 B.n2 71.676
R1016 B.n105 B.n104 63.2247
R1017 B.n111 B.n110 63.2247
R1018 B.n243 B.n242 63.2247
R1019 B.n237 B.n236 63.2247
R1020 B.n686 B.n105 59.5399
R1021 B.n668 B.n111 59.5399
R1022 B.n244 B.n243 59.5399
R1023 B.n342 B.n237 59.5399
R1024 B.n407 B.n214 53.563
R1025 B.n413 B.n214 53.563
R1026 B.n413 B.n210 53.563
R1027 B.n419 B.n210 53.563
R1028 B.n419 B.n206 53.563
R1029 B.n425 B.n206 53.563
R1030 B.n425 B.n202 53.563
R1031 B.n431 B.n202 53.563
R1032 B.n437 B.n198 53.563
R1033 B.n437 B.n194 53.563
R1034 B.n443 B.n194 53.563
R1035 B.n443 B.n190 53.563
R1036 B.n449 B.n190 53.563
R1037 B.n449 B.n186 53.563
R1038 B.n455 B.n186 53.563
R1039 B.n455 B.n182 53.563
R1040 B.n461 B.n182 53.563
R1041 B.n461 B.n178 53.563
R1042 B.n467 B.n178 53.563
R1043 B.n473 B.n174 53.563
R1044 B.n473 B.n170 53.563
R1045 B.n479 B.n170 53.563
R1046 B.n479 B.n166 53.563
R1047 B.n485 B.n166 53.563
R1048 B.n485 B.n162 53.563
R1049 B.n491 B.n162 53.563
R1050 B.n491 B.n158 53.563
R1051 B.n497 B.n158 53.563
R1052 B.n503 B.n154 53.563
R1053 B.n503 B.n150 53.563
R1054 B.n509 B.n150 53.563
R1055 B.n509 B.n146 53.563
R1056 B.n515 B.n146 53.563
R1057 B.n515 B.n142 53.563
R1058 B.n521 B.n142 53.563
R1059 B.n521 B.n138 53.563
R1060 B.n527 B.n138 53.563
R1061 B.n534 B.n134 53.563
R1062 B.n534 B.n130 53.563
R1063 B.n540 B.n130 53.563
R1064 B.n540 B.n4 53.563
R1065 B.n844 B.n4 53.563
R1066 B.n844 B.n843 53.563
R1067 B.n843 B.n842 53.563
R1068 B.n842 B.n8 53.563
R1069 B.n12 B.n8 53.563
R1070 B.n835 B.n12 53.563
R1071 B.n835 B.n834 53.563
R1072 B.n833 B.n16 53.563
R1073 B.n827 B.n16 53.563
R1074 B.n827 B.n826 53.563
R1075 B.n826 B.n825 53.563
R1076 B.n825 B.n23 53.563
R1077 B.n819 B.n23 53.563
R1078 B.n819 B.n818 53.563
R1079 B.n818 B.n817 53.563
R1080 B.n817 B.n30 53.563
R1081 B.n811 B.n810 53.563
R1082 B.n810 B.n809 53.563
R1083 B.n809 B.n37 53.563
R1084 B.n803 B.n37 53.563
R1085 B.n803 B.n802 53.563
R1086 B.n802 B.n801 53.563
R1087 B.n801 B.n44 53.563
R1088 B.n795 B.n44 53.563
R1089 B.n795 B.n794 53.563
R1090 B.n793 B.n51 53.563
R1091 B.n787 B.n51 53.563
R1092 B.n787 B.n786 53.563
R1093 B.n786 B.n785 53.563
R1094 B.n785 B.n58 53.563
R1095 B.n779 B.n58 53.563
R1096 B.n779 B.n778 53.563
R1097 B.n778 B.n777 53.563
R1098 B.n777 B.n65 53.563
R1099 B.n771 B.n65 53.563
R1100 B.n771 B.n770 53.563
R1101 B.n769 B.n72 53.563
R1102 B.n763 B.n72 53.563
R1103 B.n763 B.n762 53.563
R1104 B.n762 B.n761 53.563
R1105 B.n761 B.n79 53.563
R1106 B.n755 B.n79 53.563
R1107 B.n755 B.n754 53.563
R1108 B.n754 B.n753 53.563
R1109 B.n467 B.t1 49.6246
R1110 B.t2 B.n793 49.6246
R1111 B.t3 B.n134 48.0492
R1112 B.n834 B.t4 48.0492
R1113 B.t14 B.n198 46.4738
R1114 B.n770 B.t7 46.4738
R1115 B.n405 B.n404 33.8737
R1116 B.n409 B.n216 33.8737
R1117 B.n604 B.n603 33.8737
R1118 B.n751 B.n750 33.8737
R1119 B.n497 B.t5 27.5694
R1120 B.n811 B.t0 27.5694
R1121 B.t5 B.n154 25.9941
R1122 B.t0 B.n30 25.9941
R1123 B B.n847 18.0485
R1124 B.n405 B.n212 10.6151
R1125 B.n415 B.n212 10.6151
R1126 B.n416 B.n415 10.6151
R1127 B.n417 B.n416 10.6151
R1128 B.n417 B.n204 10.6151
R1129 B.n427 B.n204 10.6151
R1130 B.n428 B.n427 10.6151
R1131 B.n429 B.n428 10.6151
R1132 B.n429 B.n196 10.6151
R1133 B.n439 B.n196 10.6151
R1134 B.n440 B.n439 10.6151
R1135 B.n441 B.n440 10.6151
R1136 B.n441 B.n188 10.6151
R1137 B.n451 B.n188 10.6151
R1138 B.n452 B.n451 10.6151
R1139 B.n453 B.n452 10.6151
R1140 B.n453 B.n180 10.6151
R1141 B.n463 B.n180 10.6151
R1142 B.n464 B.n463 10.6151
R1143 B.n465 B.n464 10.6151
R1144 B.n465 B.n172 10.6151
R1145 B.n475 B.n172 10.6151
R1146 B.n476 B.n475 10.6151
R1147 B.n477 B.n476 10.6151
R1148 B.n477 B.n164 10.6151
R1149 B.n487 B.n164 10.6151
R1150 B.n488 B.n487 10.6151
R1151 B.n489 B.n488 10.6151
R1152 B.n489 B.n156 10.6151
R1153 B.n499 B.n156 10.6151
R1154 B.n500 B.n499 10.6151
R1155 B.n501 B.n500 10.6151
R1156 B.n501 B.n148 10.6151
R1157 B.n511 B.n148 10.6151
R1158 B.n512 B.n511 10.6151
R1159 B.n513 B.n512 10.6151
R1160 B.n513 B.n140 10.6151
R1161 B.n523 B.n140 10.6151
R1162 B.n524 B.n523 10.6151
R1163 B.n525 B.n524 10.6151
R1164 B.n525 B.n132 10.6151
R1165 B.n536 B.n132 10.6151
R1166 B.n537 B.n536 10.6151
R1167 B.n538 B.n537 10.6151
R1168 B.n538 B.n0 10.6151
R1169 B.n404 B.n403 10.6151
R1170 B.n403 B.n220 10.6151
R1171 B.n398 B.n220 10.6151
R1172 B.n398 B.n397 10.6151
R1173 B.n397 B.n222 10.6151
R1174 B.n392 B.n222 10.6151
R1175 B.n392 B.n391 10.6151
R1176 B.n391 B.n390 10.6151
R1177 B.n390 B.n224 10.6151
R1178 B.n384 B.n224 10.6151
R1179 B.n384 B.n383 10.6151
R1180 B.n383 B.n382 10.6151
R1181 B.n382 B.n226 10.6151
R1182 B.n376 B.n226 10.6151
R1183 B.n376 B.n375 10.6151
R1184 B.n375 B.n374 10.6151
R1185 B.n374 B.n228 10.6151
R1186 B.n368 B.n228 10.6151
R1187 B.n368 B.n367 10.6151
R1188 B.n367 B.n366 10.6151
R1189 B.n366 B.n230 10.6151
R1190 B.n360 B.n230 10.6151
R1191 B.n360 B.n359 10.6151
R1192 B.n359 B.n358 10.6151
R1193 B.n358 B.n232 10.6151
R1194 B.n352 B.n232 10.6151
R1195 B.n352 B.n351 10.6151
R1196 B.n351 B.n350 10.6151
R1197 B.n350 B.n234 10.6151
R1198 B.n344 B.n234 10.6151
R1199 B.n344 B.n343 10.6151
R1200 B.n341 B.n238 10.6151
R1201 B.n335 B.n238 10.6151
R1202 B.n335 B.n334 10.6151
R1203 B.n334 B.n333 10.6151
R1204 B.n333 B.n240 10.6151
R1205 B.n327 B.n240 10.6151
R1206 B.n327 B.n326 10.6151
R1207 B.n326 B.n325 10.6151
R1208 B.n321 B.n320 10.6151
R1209 B.n320 B.n246 10.6151
R1210 B.n315 B.n246 10.6151
R1211 B.n315 B.n314 10.6151
R1212 B.n314 B.n313 10.6151
R1213 B.n313 B.n248 10.6151
R1214 B.n307 B.n248 10.6151
R1215 B.n307 B.n306 10.6151
R1216 B.n306 B.n305 10.6151
R1217 B.n305 B.n250 10.6151
R1218 B.n299 B.n250 10.6151
R1219 B.n299 B.n298 10.6151
R1220 B.n298 B.n297 10.6151
R1221 B.n297 B.n252 10.6151
R1222 B.n291 B.n252 10.6151
R1223 B.n291 B.n290 10.6151
R1224 B.n290 B.n289 10.6151
R1225 B.n289 B.n254 10.6151
R1226 B.n283 B.n254 10.6151
R1227 B.n283 B.n282 10.6151
R1228 B.n282 B.n281 10.6151
R1229 B.n281 B.n256 10.6151
R1230 B.n275 B.n256 10.6151
R1231 B.n275 B.n274 10.6151
R1232 B.n274 B.n273 10.6151
R1233 B.n273 B.n258 10.6151
R1234 B.n267 B.n258 10.6151
R1235 B.n267 B.n266 10.6151
R1236 B.n266 B.n265 10.6151
R1237 B.n265 B.n260 10.6151
R1238 B.n260 B.n216 10.6151
R1239 B.n410 B.n409 10.6151
R1240 B.n411 B.n410 10.6151
R1241 B.n411 B.n208 10.6151
R1242 B.n421 B.n208 10.6151
R1243 B.n422 B.n421 10.6151
R1244 B.n423 B.n422 10.6151
R1245 B.n423 B.n200 10.6151
R1246 B.n433 B.n200 10.6151
R1247 B.n434 B.n433 10.6151
R1248 B.n435 B.n434 10.6151
R1249 B.n435 B.n192 10.6151
R1250 B.n445 B.n192 10.6151
R1251 B.n446 B.n445 10.6151
R1252 B.n447 B.n446 10.6151
R1253 B.n447 B.n184 10.6151
R1254 B.n457 B.n184 10.6151
R1255 B.n458 B.n457 10.6151
R1256 B.n459 B.n458 10.6151
R1257 B.n459 B.n176 10.6151
R1258 B.n469 B.n176 10.6151
R1259 B.n470 B.n469 10.6151
R1260 B.n471 B.n470 10.6151
R1261 B.n471 B.n168 10.6151
R1262 B.n481 B.n168 10.6151
R1263 B.n482 B.n481 10.6151
R1264 B.n483 B.n482 10.6151
R1265 B.n483 B.n160 10.6151
R1266 B.n493 B.n160 10.6151
R1267 B.n494 B.n493 10.6151
R1268 B.n495 B.n494 10.6151
R1269 B.n495 B.n152 10.6151
R1270 B.n505 B.n152 10.6151
R1271 B.n506 B.n505 10.6151
R1272 B.n507 B.n506 10.6151
R1273 B.n507 B.n144 10.6151
R1274 B.n517 B.n144 10.6151
R1275 B.n518 B.n517 10.6151
R1276 B.n519 B.n518 10.6151
R1277 B.n519 B.n136 10.6151
R1278 B.n529 B.n136 10.6151
R1279 B.n530 B.n529 10.6151
R1280 B.n532 B.n530 10.6151
R1281 B.n532 B.n531 10.6151
R1282 B.n531 B.n128 10.6151
R1283 B.n543 B.n128 10.6151
R1284 B.n544 B.n543 10.6151
R1285 B.n545 B.n544 10.6151
R1286 B.n546 B.n545 10.6151
R1287 B.n547 B.n546 10.6151
R1288 B.n550 B.n547 10.6151
R1289 B.n551 B.n550 10.6151
R1290 B.n552 B.n551 10.6151
R1291 B.n553 B.n552 10.6151
R1292 B.n555 B.n553 10.6151
R1293 B.n556 B.n555 10.6151
R1294 B.n557 B.n556 10.6151
R1295 B.n558 B.n557 10.6151
R1296 B.n560 B.n558 10.6151
R1297 B.n561 B.n560 10.6151
R1298 B.n562 B.n561 10.6151
R1299 B.n563 B.n562 10.6151
R1300 B.n565 B.n563 10.6151
R1301 B.n566 B.n565 10.6151
R1302 B.n567 B.n566 10.6151
R1303 B.n568 B.n567 10.6151
R1304 B.n570 B.n568 10.6151
R1305 B.n571 B.n570 10.6151
R1306 B.n572 B.n571 10.6151
R1307 B.n573 B.n572 10.6151
R1308 B.n575 B.n573 10.6151
R1309 B.n576 B.n575 10.6151
R1310 B.n577 B.n576 10.6151
R1311 B.n578 B.n577 10.6151
R1312 B.n580 B.n578 10.6151
R1313 B.n581 B.n580 10.6151
R1314 B.n582 B.n581 10.6151
R1315 B.n583 B.n582 10.6151
R1316 B.n585 B.n583 10.6151
R1317 B.n586 B.n585 10.6151
R1318 B.n587 B.n586 10.6151
R1319 B.n588 B.n587 10.6151
R1320 B.n590 B.n588 10.6151
R1321 B.n591 B.n590 10.6151
R1322 B.n592 B.n591 10.6151
R1323 B.n593 B.n592 10.6151
R1324 B.n595 B.n593 10.6151
R1325 B.n596 B.n595 10.6151
R1326 B.n597 B.n596 10.6151
R1327 B.n598 B.n597 10.6151
R1328 B.n600 B.n598 10.6151
R1329 B.n601 B.n600 10.6151
R1330 B.n602 B.n601 10.6151
R1331 B.n603 B.n602 10.6151
R1332 B.n839 B.n1 10.6151
R1333 B.n839 B.n838 10.6151
R1334 B.n838 B.n837 10.6151
R1335 B.n837 B.n10 10.6151
R1336 B.n831 B.n10 10.6151
R1337 B.n831 B.n830 10.6151
R1338 B.n830 B.n829 10.6151
R1339 B.n829 B.n18 10.6151
R1340 B.n823 B.n18 10.6151
R1341 B.n823 B.n822 10.6151
R1342 B.n822 B.n821 10.6151
R1343 B.n821 B.n25 10.6151
R1344 B.n815 B.n25 10.6151
R1345 B.n815 B.n814 10.6151
R1346 B.n814 B.n813 10.6151
R1347 B.n813 B.n32 10.6151
R1348 B.n807 B.n32 10.6151
R1349 B.n807 B.n806 10.6151
R1350 B.n806 B.n805 10.6151
R1351 B.n805 B.n39 10.6151
R1352 B.n799 B.n39 10.6151
R1353 B.n799 B.n798 10.6151
R1354 B.n798 B.n797 10.6151
R1355 B.n797 B.n46 10.6151
R1356 B.n791 B.n46 10.6151
R1357 B.n791 B.n790 10.6151
R1358 B.n790 B.n789 10.6151
R1359 B.n789 B.n53 10.6151
R1360 B.n783 B.n53 10.6151
R1361 B.n783 B.n782 10.6151
R1362 B.n782 B.n781 10.6151
R1363 B.n781 B.n60 10.6151
R1364 B.n775 B.n60 10.6151
R1365 B.n775 B.n774 10.6151
R1366 B.n774 B.n773 10.6151
R1367 B.n773 B.n67 10.6151
R1368 B.n767 B.n67 10.6151
R1369 B.n767 B.n766 10.6151
R1370 B.n766 B.n765 10.6151
R1371 B.n765 B.n74 10.6151
R1372 B.n759 B.n74 10.6151
R1373 B.n759 B.n758 10.6151
R1374 B.n758 B.n757 10.6151
R1375 B.n757 B.n81 10.6151
R1376 B.n751 B.n81 10.6151
R1377 B.n750 B.n749 10.6151
R1378 B.n749 B.n88 10.6151
R1379 B.n743 B.n88 10.6151
R1380 B.n743 B.n742 10.6151
R1381 B.n742 B.n741 10.6151
R1382 B.n741 B.n90 10.6151
R1383 B.n735 B.n90 10.6151
R1384 B.n735 B.n734 10.6151
R1385 B.n734 B.n733 10.6151
R1386 B.n733 B.n92 10.6151
R1387 B.n727 B.n92 10.6151
R1388 B.n727 B.n726 10.6151
R1389 B.n726 B.n725 10.6151
R1390 B.n725 B.n94 10.6151
R1391 B.n719 B.n94 10.6151
R1392 B.n719 B.n718 10.6151
R1393 B.n718 B.n717 10.6151
R1394 B.n717 B.n96 10.6151
R1395 B.n711 B.n96 10.6151
R1396 B.n711 B.n710 10.6151
R1397 B.n710 B.n709 10.6151
R1398 B.n709 B.n98 10.6151
R1399 B.n703 B.n98 10.6151
R1400 B.n703 B.n702 10.6151
R1401 B.n702 B.n701 10.6151
R1402 B.n701 B.n100 10.6151
R1403 B.n695 B.n100 10.6151
R1404 B.n695 B.n694 10.6151
R1405 B.n694 B.n693 10.6151
R1406 B.n693 B.n102 10.6151
R1407 B.n687 B.n102 10.6151
R1408 B.n685 B.n684 10.6151
R1409 B.n684 B.n106 10.6151
R1410 B.n678 B.n106 10.6151
R1411 B.n678 B.n677 10.6151
R1412 B.n677 B.n676 10.6151
R1413 B.n676 B.n108 10.6151
R1414 B.n670 B.n108 10.6151
R1415 B.n670 B.n669 10.6151
R1416 B.n667 B.n112 10.6151
R1417 B.n661 B.n112 10.6151
R1418 B.n661 B.n660 10.6151
R1419 B.n660 B.n659 10.6151
R1420 B.n659 B.n114 10.6151
R1421 B.n653 B.n114 10.6151
R1422 B.n653 B.n652 10.6151
R1423 B.n652 B.n651 10.6151
R1424 B.n651 B.n116 10.6151
R1425 B.n645 B.n116 10.6151
R1426 B.n645 B.n644 10.6151
R1427 B.n644 B.n643 10.6151
R1428 B.n643 B.n118 10.6151
R1429 B.n637 B.n118 10.6151
R1430 B.n637 B.n636 10.6151
R1431 B.n636 B.n635 10.6151
R1432 B.n635 B.n120 10.6151
R1433 B.n629 B.n120 10.6151
R1434 B.n629 B.n628 10.6151
R1435 B.n628 B.n627 10.6151
R1436 B.n627 B.n122 10.6151
R1437 B.n621 B.n122 10.6151
R1438 B.n621 B.n620 10.6151
R1439 B.n620 B.n619 10.6151
R1440 B.n619 B.n124 10.6151
R1441 B.n613 B.n124 10.6151
R1442 B.n613 B.n612 10.6151
R1443 B.n612 B.n611 10.6151
R1444 B.n611 B.n126 10.6151
R1445 B.n605 B.n126 10.6151
R1446 B.n605 B.n604 10.6151
R1447 B.n847 B.n0 8.11757
R1448 B.n847 B.n1 8.11757
R1449 B.n431 B.t14 7.08965
R1450 B.t7 B.n769 7.08965
R1451 B.n342 B.n341 6.5566
R1452 B.n325 B.n244 6.5566
R1453 B.n686 B.n685 6.5566
R1454 B.n669 B.n668 6.5566
R1455 B.n527 B.t3 5.51428
R1456 B.t4 B.n833 5.51428
R1457 B.n343 B.n342 4.05904
R1458 B.n321 B.n244 4.05904
R1459 B.n687 B.n686 4.05904
R1460 B.n668 B.n667 4.05904
R1461 B.t1 B.n174 3.93892
R1462 B.n794 B.t2 3.93892
R1463 VP.n14 VP.n11 161.3
R1464 VP.n16 VP.n15 161.3
R1465 VP.n17 VP.n10 161.3
R1466 VP.n19 VP.n18 161.3
R1467 VP.n20 VP.n9 161.3
R1468 VP.n22 VP.n21 161.3
R1469 VP.n23 VP.n8 161.3
R1470 VP.n48 VP.n0 161.3
R1471 VP.n47 VP.n46 161.3
R1472 VP.n45 VP.n1 161.3
R1473 VP.n44 VP.n43 161.3
R1474 VP.n42 VP.n2 161.3
R1475 VP.n41 VP.n40 161.3
R1476 VP.n39 VP.n3 161.3
R1477 VP.n38 VP.n37 161.3
R1478 VP.n35 VP.n4 161.3
R1479 VP.n34 VP.n33 161.3
R1480 VP.n32 VP.n5 161.3
R1481 VP.n31 VP.n30 161.3
R1482 VP.n29 VP.n6 161.3
R1483 VP.n28 VP.n27 161.3
R1484 VP.n26 VP.n7 110.267
R1485 VP.n50 VP.n49 110.267
R1486 VP.n25 VP.n24 110.267
R1487 VP.n13 VP.t0 103.543
R1488 VP.n7 VP.t1 71.478
R1489 VP.n36 VP.t3 71.478
R1490 VP.n49 VP.t5 71.478
R1491 VP.n24 VP.t4 71.478
R1492 VP.n12 VP.t2 71.478
R1493 VP.n13 VP.n12 61.624
R1494 VP.n34 VP.n5 52.1486
R1495 VP.n43 VP.n42 52.1486
R1496 VP.n18 VP.n17 52.1486
R1497 VP.n26 VP.n25 47.4163
R1498 VP.n30 VP.n5 28.8382
R1499 VP.n43 VP.n1 28.8382
R1500 VP.n18 VP.n9 28.8382
R1501 VP.n29 VP.n28 24.4675
R1502 VP.n30 VP.n29 24.4675
R1503 VP.n35 VP.n34 24.4675
R1504 VP.n37 VP.n35 24.4675
R1505 VP.n41 VP.n3 24.4675
R1506 VP.n42 VP.n41 24.4675
R1507 VP.n47 VP.n1 24.4675
R1508 VP.n48 VP.n47 24.4675
R1509 VP.n22 VP.n9 24.4675
R1510 VP.n23 VP.n22 24.4675
R1511 VP.n16 VP.n11 24.4675
R1512 VP.n17 VP.n16 24.4675
R1513 VP.n37 VP.n36 12.234
R1514 VP.n36 VP.n3 12.234
R1515 VP.n12 VP.n11 12.234
R1516 VP.n14 VP.n13 5.19435
R1517 VP.n28 VP.n7 0.48984
R1518 VP.n49 VP.n48 0.48984
R1519 VP.n24 VP.n23 0.48984
R1520 VP.n25 VP.n8 0.278367
R1521 VP.n27 VP.n26 0.278367
R1522 VP.n50 VP.n0 0.278367
R1523 VP.n15 VP.n14 0.189894
R1524 VP.n15 VP.n10 0.189894
R1525 VP.n19 VP.n10 0.189894
R1526 VP.n20 VP.n19 0.189894
R1527 VP.n21 VP.n20 0.189894
R1528 VP.n21 VP.n8 0.189894
R1529 VP.n27 VP.n6 0.189894
R1530 VP.n31 VP.n6 0.189894
R1531 VP.n32 VP.n31 0.189894
R1532 VP.n33 VP.n32 0.189894
R1533 VP.n33 VP.n4 0.189894
R1534 VP.n38 VP.n4 0.189894
R1535 VP.n39 VP.n38 0.189894
R1536 VP.n40 VP.n39 0.189894
R1537 VP.n40 VP.n2 0.189894
R1538 VP.n44 VP.n2 0.189894
R1539 VP.n45 VP.n44 0.189894
R1540 VP.n46 VP.n45 0.189894
R1541 VP.n46 VP.n0 0.189894
R1542 VP VP.n50 0.153454
R1543 VTAIL.n186 VTAIL.n146 289.615
R1544 VTAIL.n42 VTAIL.n2 289.615
R1545 VTAIL.n140 VTAIL.n100 289.615
R1546 VTAIL.n92 VTAIL.n52 289.615
R1547 VTAIL.n161 VTAIL.n160 185
R1548 VTAIL.n158 VTAIL.n157 185
R1549 VTAIL.n167 VTAIL.n166 185
R1550 VTAIL.n169 VTAIL.n168 185
R1551 VTAIL.n154 VTAIL.n153 185
R1552 VTAIL.n175 VTAIL.n174 185
R1553 VTAIL.n178 VTAIL.n177 185
R1554 VTAIL.n176 VTAIL.n150 185
R1555 VTAIL.n183 VTAIL.n149 185
R1556 VTAIL.n185 VTAIL.n184 185
R1557 VTAIL.n187 VTAIL.n186 185
R1558 VTAIL.n17 VTAIL.n16 185
R1559 VTAIL.n14 VTAIL.n13 185
R1560 VTAIL.n23 VTAIL.n22 185
R1561 VTAIL.n25 VTAIL.n24 185
R1562 VTAIL.n10 VTAIL.n9 185
R1563 VTAIL.n31 VTAIL.n30 185
R1564 VTAIL.n34 VTAIL.n33 185
R1565 VTAIL.n32 VTAIL.n6 185
R1566 VTAIL.n39 VTAIL.n5 185
R1567 VTAIL.n41 VTAIL.n40 185
R1568 VTAIL.n43 VTAIL.n42 185
R1569 VTAIL.n141 VTAIL.n140 185
R1570 VTAIL.n139 VTAIL.n138 185
R1571 VTAIL.n137 VTAIL.n103 185
R1572 VTAIL.n107 VTAIL.n104 185
R1573 VTAIL.n132 VTAIL.n131 185
R1574 VTAIL.n130 VTAIL.n129 185
R1575 VTAIL.n109 VTAIL.n108 185
R1576 VTAIL.n124 VTAIL.n123 185
R1577 VTAIL.n122 VTAIL.n121 185
R1578 VTAIL.n113 VTAIL.n112 185
R1579 VTAIL.n116 VTAIL.n115 185
R1580 VTAIL.n93 VTAIL.n92 185
R1581 VTAIL.n91 VTAIL.n90 185
R1582 VTAIL.n89 VTAIL.n55 185
R1583 VTAIL.n59 VTAIL.n56 185
R1584 VTAIL.n84 VTAIL.n83 185
R1585 VTAIL.n82 VTAIL.n81 185
R1586 VTAIL.n61 VTAIL.n60 185
R1587 VTAIL.n76 VTAIL.n75 185
R1588 VTAIL.n74 VTAIL.n73 185
R1589 VTAIL.n65 VTAIL.n64 185
R1590 VTAIL.n68 VTAIL.n67 185
R1591 VTAIL.t1 VTAIL.n159 149.524
R1592 VTAIL.t10 VTAIL.n15 149.524
R1593 VTAIL.t11 VTAIL.n114 149.524
R1594 VTAIL.t3 VTAIL.n66 149.524
R1595 VTAIL.n160 VTAIL.n157 104.615
R1596 VTAIL.n167 VTAIL.n157 104.615
R1597 VTAIL.n168 VTAIL.n167 104.615
R1598 VTAIL.n168 VTAIL.n153 104.615
R1599 VTAIL.n175 VTAIL.n153 104.615
R1600 VTAIL.n177 VTAIL.n175 104.615
R1601 VTAIL.n177 VTAIL.n176 104.615
R1602 VTAIL.n176 VTAIL.n149 104.615
R1603 VTAIL.n185 VTAIL.n149 104.615
R1604 VTAIL.n186 VTAIL.n185 104.615
R1605 VTAIL.n16 VTAIL.n13 104.615
R1606 VTAIL.n23 VTAIL.n13 104.615
R1607 VTAIL.n24 VTAIL.n23 104.615
R1608 VTAIL.n24 VTAIL.n9 104.615
R1609 VTAIL.n31 VTAIL.n9 104.615
R1610 VTAIL.n33 VTAIL.n31 104.615
R1611 VTAIL.n33 VTAIL.n32 104.615
R1612 VTAIL.n32 VTAIL.n5 104.615
R1613 VTAIL.n41 VTAIL.n5 104.615
R1614 VTAIL.n42 VTAIL.n41 104.615
R1615 VTAIL.n140 VTAIL.n139 104.615
R1616 VTAIL.n139 VTAIL.n103 104.615
R1617 VTAIL.n107 VTAIL.n103 104.615
R1618 VTAIL.n131 VTAIL.n107 104.615
R1619 VTAIL.n131 VTAIL.n130 104.615
R1620 VTAIL.n130 VTAIL.n108 104.615
R1621 VTAIL.n123 VTAIL.n108 104.615
R1622 VTAIL.n123 VTAIL.n122 104.615
R1623 VTAIL.n122 VTAIL.n112 104.615
R1624 VTAIL.n115 VTAIL.n112 104.615
R1625 VTAIL.n92 VTAIL.n91 104.615
R1626 VTAIL.n91 VTAIL.n55 104.615
R1627 VTAIL.n59 VTAIL.n55 104.615
R1628 VTAIL.n83 VTAIL.n59 104.615
R1629 VTAIL.n83 VTAIL.n82 104.615
R1630 VTAIL.n82 VTAIL.n60 104.615
R1631 VTAIL.n75 VTAIL.n60 104.615
R1632 VTAIL.n75 VTAIL.n74 104.615
R1633 VTAIL.n74 VTAIL.n64 104.615
R1634 VTAIL.n67 VTAIL.n64 104.615
R1635 VTAIL.n160 VTAIL.t1 52.3082
R1636 VTAIL.n16 VTAIL.t10 52.3082
R1637 VTAIL.n115 VTAIL.t11 52.3082
R1638 VTAIL.n67 VTAIL.t3 52.3082
R1639 VTAIL.n99 VTAIL.n98 50.0594
R1640 VTAIL.n51 VTAIL.n50 50.0594
R1641 VTAIL.n1 VTAIL.n0 50.0592
R1642 VTAIL.n49 VTAIL.n48 50.0592
R1643 VTAIL.n191 VTAIL.n190 35.4823
R1644 VTAIL.n47 VTAIL.n46 35.4823
R1645 VTAIL.n145 VTAIL.n144 35.4823
R1646 VTAIL.n97 VTAIL.n96 35.4823
R1647 VTAIL.n51 VTAIL.n49 25.4789
R1648 VTAIL.n191 VTAIL.n145 22.6686
R1649 VTAIL.n184 VTAIL.n183 13.1884
R1650 VTAIL.n40 VTAIL.n39 13.1884
R1651 VTAIL.n138 VTAIL.n137 13.1884
R1652 VTAIL.n90 VTAIL.n89 13.1884
R1653 VTAIL.n182 VTAIL.n150 12.8005
R1654 VTAIL.n187 VTAIL.n148 12.8005
R1655 VTAIL.n38 VTAIL.n6 12.8005
R1656 VTAIL.n43 VTAIL.n4 12.8005
R1657 VTAIL.n141 VTAIL.n102 12.8005
R1658 VTAIL.n136 VTAIL.n104 12.8005
R1659 VTAIL.n93 VTAIL.n54 12.8005
R1660 VTAIL.n88 VTAIL.n56 12.8005
R1661 VTAIL.n179 VTAIL.n178 12.0247
R1662 VTAIL.n188 VTAIL.n146 12.0247
R1663 VTAIL.n35 VTAIL.n34 12.0247
R1664 VTAIL.n44 VTAIL.n2 12.0247
R1665 VTAIL.n142 VTAIL.n100 12.0247
R1666 VTAIL.n133 VTAIL.n132 12.0247
R1667 VTAIL.n94 VTAIL.n52 12.0247
R1668 VTAIL.n85 VTAIL.n84 12.0247
R1669 VTAIL.n174 VTAIL.n152 11.249
R1670 VTAIL.n30 VTAIL.n8 11.249
R1671 VTAIL.n129 VTAIL.n106 11.249
R1672 VTAIL.n81 VTAIL.n58 11.249
R1673 VTAIL.n173 VTAIL.n154 10.4732
R1674 VTAIL.n29 VTAIL.n10 10.4732
R1675 VTAIL.n128 VTAIL.n109 10.4732
R1676 VTAIL.n80 VTAIL.n61 10.4732
R1677 VTAIL.n161 VTAIL.n159 10.2747
R1678 VTAIL.n17 VTAIL.n15 10.2747
R1679 VTAIL.n116 VTAIL.n114 10.2747
R1680 VTAIL.n68 VTAIL.n66 10.2747
R1681 VTAIL.n170 VTAIL.n169 9.69747
R1682 VTAIL.n26 VTAIL.n25 9.69747
R1683 VTAIL.n125 VTAIL.n124 9.69747
R1684 VTAIL.n77 VTAIL.n76 9.69747
R1685 VTAIL.n190 VTAIL.n189 9.45567
R1686 VTAIL.n46 VTAIL.n45 9.45567
R1687 VTAIL.n144 VTAIL.n143 9.45567
R1688 VTAIL.n96 VTAIL.n95 9.45567
R1689 VTAIL.n189 VTAIL.n188 9.3005
R1690 VTAIL.n148 VTAIL.n147 9.3005
R1691 VTAIL.n163 VTAIL.n162 9.3005
R1692 VTAIL.n165 VTAIL.n164 9.3005
R1693 VTAIL.n156 VTAIL.n155 9.3005
R1694 VTAIL.n171 VTAIL.n170 9.3005
R1695 VTAIL.n173 VTAIL.n172 9.3005
R1696 VTAIL.n152 VTAIL.n151 9.3005
R1697 VTAIL.n180 VTAIL.n179 9.3005
R1698 VTAIL.n182 VTAIL.n181 9.3005
R1699 VTAIL.n45 VTAIL.n44 9.3005
R1700 VTAIL.n4 VTAIL.n3 9.3005
R1701 VTAIL.n19 VTAIL.n18 9.3005
R1702 VTAIL.n21 VTAIL.n20 9.3005
R1703 VTAIL.n12 VTAIL.n11 9.3005
R1704 VTAIL.n27 VTAIL.n26 9.3005
R1705 VTAIL.n29 VTAIL.n28 9.3005
R1706 VTAIL.n8 VTAIL.n7 9.3005
R1707 VTAIL.n36 VTAIL.n35 9.3005
R1708 VTAIL.n38 VTAIL.n37 9.3005
R1709 VTAIL.n118 VTAIL.n117 9.3005
R1710 VTAIL.n120 VTAIL.n119 9.3005
R1711 VTAIL.n111 VTAIL.n110 9.3005
R1712 VTAIL.n126 VTAIL.n125 9.3005
R1713 VTAIL.n128 VTAIL.n127 9.3005
R1714 VTAIL.n106 VTAIL.n105 9.3005
R1715 VTAIL.n134 VTAIL.n133 9.3005
R1716 VTAIL.n136 VTAIL.n135 9.3005
R1717 VTAIL.n143 VTAIL.n142 9.3005
R1718 VTAIL.n102 VTAIL.n101 9.3005
R1719 VTAIL.n70 VTAIL.n69 9.3005
R1720 VTAIL.n72 VTAIL.n71 9.3005
R1721 VTAIL.n63 VTAIL.n62 9.3005
R1722 VTAIL.n78 VTAIL.n77 9.3005
R1723 VTAIL.n80 VTAIL.n79 9.3005
R1724 VTAIL.n58 VTAIL.n57 9.3005
R1725 VTAIL.n86 VTAIL.n85 9.3005
R1726 VTAIL.n88 VTAIL.n87 9.3005
R1727 VTAIL.n95 VTAIL.n94 9.3005
R1728 VTAIL.n54 VTAIL.n53 9.3005
R1729 VTAIL.n166 VTAIL.n156 8.92171
R1730 VTAIL.n22 VTAIL.n12 8.92171
R1731 VTAIL.n121 VTAIL.n111 8.92171
R1732 VTAIL.n73 VTAIL.n63 8.92171
R1733 VTAIL.n165 VTAIL.n158 8.14595
R1734 VTAIL.n21 VTAIL.n14 8.14595
R1735 VTAIL.n120 VTAIL.n113 8.14595
R1736 VTAIL.n72 VTAIL.n65 8.14595
R1737 VTAIL.n162 VTAIL.n161 7.3702
R1738 VTAIL.n18 VTAIL.n17 7.3702
R1739 VTAIL.n117 VTAIL.n116 7.3702
R1740 VTAIL.n69 VTAIL.n68 7.3702
R1741 VTAIL.n162 VTAIL.n158 5.81868
R1742 VTAIL.n18 VTAIL.n14 5.81868
R1743 VTAIL.n117 VTAIL.n113 5.81868
R1744 VTAIL.n69 VTAIL.n65 5.81868
R1745 VTAIL.n166 VTAIL.n165 5.04292
R1746 VTAIL.n22 VTAIL.n21 5.04292
R1747 VTAIL.n121 VTAIL.n120 5.04292
R1748 VTAIL.n73 VTAIL.n72 5.04292
R1749 VTAIL.n169 VTAIL.n156 4.26717
R1750 VTAIL.n25 VTAIL.n12 4.26717
R1751 VTAIL.n124 VTAIL.n111 4.26717
R1752 VTAIL.n76 VTAIL.n63 4.26717
R1753 VTAIL.n170 VTAIL.n154 3.49141
R1754 VTAIL.n26 VTAIL.n10 3.49141
R1755 VTAIL.n125 VTAIL.n109 3.49141
R1756 VTAIL.n77 VTAIL.n61 3.49141
R1757 VTAIL.n163 VTAIL.n159 2.84303
R1758 VTAIL.n19 VTAIL.n15 2.84303
R1759 VTAIL.n118 VTAIL.n114 2.84303
R1760 VTAIL.n70 VTAIL.n66 2.84303
R1761 VTAIL.n97 VTAIL.n51 2.81084
R1762 VTAIL.n145 VTAIL.n99 2.81084
R1763 VTAIL.n49 VTAIL.n47 2.81084
R1764 VTAIL.n174 VTAIL.n173 2.71565
R1765 VTAIL.n30 VTAIL.n29 2.71565
R1766 VTAIL.n129 VTAIL.n128 2.71565
R1767 VTAIL.n81 VTAIL.n80 2.71565
R1768 VTAIL.n0 VTAIL.t5 2.27898
R1769 VTAIL.n0 VTAIL.t0 2.27898
R1770 VTAIL.n48 VTAIL.t6 2.27898
R1771 VTAIL.n48 VTAIL.t8 2.27898
R1772 VTAIL.n98 VTAIL.t9 2.27898
R1773 VTAIL.n98 VTAIL.t7 2.27898
R1774 VTAIL.n50 VTAIL.t2 2.27898
R1775 VTAIL.n50 VTAIL.t4 2.27898
R1776 VTAIL VTAIL.n191 2.05007
R1777 VTAIL.n178 VTAIL.n152 1.93989
R1778 VTAIL.n190 VTAIL.n146 1.93989
R1779 VTAIL.n34 VTAIL.n8 1.93989
R1780 VTAIL.n46 VTAIL.n2 1.93989
R1781 VTAIL.n144 VTAIL.n100 1.93989
R1782 VTAIL.n132 VTAIL.n106 1.93989
R1783 VTAIL.n96 VTAIL.n52 1.93989
R1784 VTAIL.n84 VTAIL.n58 1.93989
R1785 VTAIL.n99 VTAIL.n97 1.8755
R1786 VTAIL.n47 VTAIL.n1 1.8755
R1787 VTAIL.n179 VTAIL.n150 1.16414
R1788 VTAIL.n188 VTAIL.n187 1.16414
R1789 VTAIL.n35 VTAIL.n6 1.16414
R1790 VTAIL.n44 VTAIL.n43 1.16414
R1791 VTAIL.n142 VTAIL.n141 1.16414
R1792 VTAIL.n133 VTAIL.n104 1.16414
R1793 VTAIL.n94 VTAIL.n93 1.16414
R1794 VTAIL.n85 VTAIL.n56 1.16414
R1795 VTAIL VTAIL.n1 0.761276
R1796 VTAIL.n183 VTAIL.n182 0.388379
R1797 VTAIL.n184 VTAIL.n148 0.388379
R1798 VTAIL.n39 VTAIL.n38 0.388379
R1799 VTAIL.n40 VTAIL.n4 0.388379
R1800 VTAIL.n138 VTAIL.n102 0.388379
R1801 VTAIL.n137 VTAIL.n136 0.388379
R1802 VTAIL.n90 VTAIL.n54 0.388379
R1803 VTAIL.n89 VTAIL.n88 0.388379
R1804 VTAIL.n164 VTAIL.n163 0.155672
R1805 VTAIL.n164 VTAIL.n155 0.155672
R1806 VTAIL.n171 VTAIL.n155 0.155672
R1807 VTAIL.n172 VTAIL.n171 0.155672
R1808 VTAIL.n172 VTAIL.n151 0.155672
R1809 VTAIL.n180 VTAIL.n151 0.155672
R1810 VTAIL.n181 VTAIL.n180 0.155672
R1811 VTAIL.n181 VTAIL.n147 0.155672
R1812 VTAIL.n189 VTAIL.n147 0.155672
R1813 VTAIL.n20 VTAIL.n19 0.155672
R1814 VTAIL.n20 VTAIL.n11 0.155672
R1815 VTAIL.n27 VTAIL.n11 0.155672
R1816 VTAIL.n28 VTAIL.n27 0.155672
R1817 VTAIL.n28 VTAIL.n7 0.155672
R1818 VTAIL.n36 VTAIL.n7 0.155672
R1819 VTAIL.n37 VTAIL.n36 0.155672
R1820 VTAIL.n37 VTAIL.n3 0.155672
R1821 VTAIL.n45 VTAIL.n3 0.155672
R1822 VTAIL.n143 VTAIL.n101 0.155672
R1823 VTAIL.n135 VTAIL.n101 0.155672
R1824 VTAIL.n135 VTAIL.n134 0.155672
R1825 VTAIL.n134 VTAIL.n105 0.155672
R1826 VTAIL.n127 VTAIL.n105 0.155672
R1827 VTAIL.n127 VTAIL.n126 0.155672
R1828 VTAIL.n126 VTAIL.n110 0.155672
R1829 VTAIL.n119 VTAIL.n110 0.155672
R1830 VTAIL.n119 VTAIL.n118 0.155672
R1831 VTAIL.n95 VTAIL.n53 0.155672
R1832 VTAIL.n87 VTAIL.n53 0.155672
R1833 VTAIL.n87 VTAIL.n86 0.155672
R1834 VTAIL.n86 VTAIL.n57 0.155672
R1835 VTAIL.n79 VTAIL.n57 0.155672
R1836 VTAIL.n79 VTAIL.n78 0.155672
R1837 VTAIL.n78 VTAIL.n62 0.155672
R1838 VTAIL.n71 VTAIL.n62 0.155672
R1839 VTAIL.n71 VTAIL.n70 0.155672
R1840 VDD1.n40 VDD1.n0 289.615
R1841 VDD1.n85 VDD1.n45 289.615
R1842 VDD1.n41 VDD1.n40 185
R1843 VDD1.n39 VDD1.n38 185
R1844 VDD1.n37 VDD1.n3 185
R1845 VDD1.n7 VDD1.n4 185
R1846 VDD1.n32 VDD1.n31 185
R1847 VDD1.n30 VDD1.n29 185
R1848 VDD1.n9 VDD1.n8 185
R1849 VDD1.n24 VDD1.n23 185
R1850 VDD1.n22 VDD1.n21 185
R1851 VDD1.n13 VDD1.n12 185
R1852 VDD1.n16 VDD1.n15 185
R1853 VDD1.n60 VDD1.n59 185
R1854 VDD1.n57 VDD1.n56 185
R1855 VDD1.n66 VDD1.n65 185
R1856 VDD1.n68 VDD1.n67 185
R1857 VDD1.n53 VDD1.n52 185
R1858 VDD1.n74 VDD1.n73 185
R1859 VDD1.n77 VDD1.n76 185
R1860 VDD1.n75 VDD1.n49 185
R1861 VDD1.n82 VDD1.n48 185
R1862 VDD1.n84 VDD1.n83 185
R1863 VDD1.n86 VDD1.n85 185
R1864 VDD1.t5 VDD1.n14 149.524
R1865 VDD1.t4 VDD1.n58 149.524
R1866 VDD1.n40 VDD1.n39 104.615
R1867 VDD1.n39 VDD1.n3 104.615
R1868 VDD1.n7 VDD1.n3 104.615
R1869 VDD1.n31 VDD1.n7 104.615
R1870 VDD1.n31 VDD1.n30 104.615
R1871 VDD1.n30 VDD1.n8 104.615
R1872 VDD1.n23 VDD1.n8 104.615
R1873 VDD1.n23 VDD1.n22 104.615
R1874 VDD1.n22 VDD1.n12 104.615
R1875 VDD1.n15 VDD1.n12 104.615
R1876 VDD1.n59 VDD1.n56 104.615
R1877 VDD1.n66 VDD1.n56 104.615
R1878 VDD1.n67 VDD1.n66 104.615
R1879 VDD1.n67 VDD1.n52 104.615
R1880 VDD1.n74 VDD1.n52 104.615
R1881 VDD1.n76 VDD1.n74 104.615
R1882 VDD1.n76 VDD1.n75 104.615
R1883 VDD1.n75 VDD1.n48 104.615
R1884 VDD1.n84 VDD1.n48 104.615
R1885 VDD1.n85 VDD1.n84 104.615
R1886 VDD1.n91 VDD1.n90 67.3852
R1887 VDD1.n93 VDD1.n92 66.738
R1888 VDD1 VDD1.n44 54.3271
R1889 VDD1.n91 VDD1.n89 54.2135
R1890 VDD1.n15 VDD1.t5 52.3082
R1891 VDD1.n59 VDD1.t4 52.3082
R1892 VDD1.n93 VDD1.n91 42.3285
R1893 VDD1.n38 VDD1.n37 13.1884
R1894 VDD1.n83 VDD1.n82 13.1884
R1895 VDD1.n41 VDD1.n2 12.8005
R1896 VDD1.n36 VDD1.n4 12.8005
R1897 VDD1.n81 VDD1.n49 12.8005
R1898 VDD1.n86 VDD1.n47 12.8005
R1899 VDD1.n42 VDD1.n0 12.0247
R1900 VDD1.n33 VDD1.n32 12.0247
R1901 VDD1.n78 VDD1.n77 12.0247
R1902 VDD1.n87 VDD1.n45 12.0247
R1903 VDD1.n29 VDD1.n6 11.249
R1904 VDD1.n73 VDD1.n51 11.249
R1905 VDD1.n28 VDD1.n9 10.4732
R1906 VDD1.n72 VDD1.n53 10.4732
R1907 VDD1.n16 VDD1.n14 10.2747
R1908 VDD1.n60 VDD1.n58 10.2747
R1909 VDD1.n25 VDD1.n24 9.69747
R1910 VDD1.n69 VDD1.n68 9.69747
R1911 VDD1.n44 VDD1.n43 9.45567
R1912 VDD1.n89 VDD1.n88 9.45567
R1913 VDD1.n18 VDD1.n17 9.3005
R1914 VDD1.n20 VDD1.n19 9.3005
R1915 VDD1.n11 VDD1.n10 9.3005
R1916 VDD1.n26 VDD1.n25 9.3005
R1917 VDD1.n28 VDD1.n27 9.3005
R1918 VDD1.n6 VDD1.n5 9.3005
R1919 VDD1.n34 VDD1.n33 9.3005
R1920 VDD1.n36 VDD1.n35 9.3005
R1921 VDD1.n43 VDD1.n42 9.3005
R1922 VDD1.n2 VDD1.n1 9.3005
R1923 VDD1.n88 VDD1.n87 9.3005
R1924 VDD1.n47 VDD1.n46 9.3005
R1925 VDD1.n62 VDD1.n61 9.3005
R1926 VDD1.n64 VDD1.n63 9.3005
R1927 VDD1.n55 VDD1.n54 9.3005
R1928 VDD1.n70 VDD1.n69 9.3005
R1929 VDD1.n72 VDD1.n71 9.3005
R1930 VDD1.n51 VDD1.n50 9.3005
R1931 VDD1.n79 VDD1.n78 9.3005
R1932 VDD1.n81 VDD1.n80 9.3005
R1933 VDD1.n21 VDD1.n11 8.92171
R1934 VDD1.n65 VDD1.n55 8.92171
R1935 VDD1.n20 VDD1.n13 8.14595
R1936 VDD1.n64 VDD1.n57 8.14595
R1937 VDD1.n17 VDD1.n16 7.3702
R1938 VDD1.n61 VDD1.n60 7.3702
R1939 VDD1.n17 VDD1.n13 5.81868
R1940 VDD1.n61 VDD1.n57 5.81868
R1941 VDD1.n21 VDD1.n20 5.04292
R1942 VDD1.n65 VDD1.n64 5.04292
R1943 VDD1.n24 VDD1.n11 4.26717
R1944 VDD1.n68 VDD1.n55 4.26717
R1945 VDD1.n25 VDD1.n9 3.49141
R1946 VDD1.n69 VDD1.n53 3.49141
R1947 VDD1.n62 VDD1.n58 2.84303
R1948 VDD1.n18 VDD1.n14 2.84303
R1949 VDD1.n29 VDD1.n28 2.71565
R1950 VDD1.n73 VDD1.n72 2.71565
R1951 VDD1.n92 VDD1.t3 2.27898
R1952 VDD1.n92 VDD1.t1 2.27898
R1953 VDD1.n90 VDD1.t2 2.27898
R1954 VDD1.n90 VDD1.t0 2.27898
R1955 VDD1.n44 VDD1.n0 1.93989
R1956 VDD1.n32 VDD1.n6 1.93989
R1957 VDD1.n77 VDD1.n51 1.93989
R1958 VDD1.n89 VDD1.n45 1.93989
R1959 VDD1.n42 VDD1.n41 1.16414
R1960 VDD1.n33 VDD1.n4 1.16414
R1961 VDD1.n78 VDD1.n49 1.16414
R1962 VDD1.n87 VDD1.n86 1.16414
R1963 VDD1 VDD1.n93 0.644897
R1964 VDD1.n38 VDD1.n2 0.388379
R1965 VDD1.n37 VDD1.n36 0.388379
R1966 VDD1.n82 VDD1.n81 0.388379
R1967 VDD1.n83 VDD1.n47 0.388379
R1968 VDD1.n43 VDD1.n1 0.155672
R1969 VDD1.n35 VDD1.n1 0.155672
R1970 VDD1.n35 VDD1.n34 0.155672
R1971 VDD1.n34 VDD1.n5 0.155672
R1972 VDD1.n27 VDD1.n5 0.155672
R1973 VDD1.n27 VDD1.n26 0.155672
R1974 VDD1.n26 VDD1.n10 0.155672
R1975 VDD1.n19 VDD1.n10 0.155672
R1976 VDD1.n19 VDD1.n18 0.155672
R1977 VDD1.n63 VDD1.n62 0.155672
R1978 VDD1.n63 VDD1.n54 0.155672
R1979 VDD1.n70 VDD1.n54 0.155672
R1980 VDD1.n71 VDD1.n70 0.155672
R1981 VDD1.n71 VDD1.n50 0.155672
R1982 VDD1.n79 VDD1.n50 0.155672
R1983 VDD1.n80 VDD1.n79 0.155672
R1984 VDD1.n80 VDD1.n46 0.155672
R1985 VDD1.n88 VDD1.n46 0.155672
R1986 VN.n33 VN.n18 161.3
R1987 VN.n32 VN.n31 161.3
R1988 VN.n30 VN.n19 161.3
R1989 VN.n29 VN.n28 161.3
R1990 VN.n27 VN.n20 161.3
R1991 VN.n26 VN.n25 161.3
R1992 VN.n24 VN.n21 161.3
R1993 VN.n15 VN.n0 161.3
R1994 VN.n14 VN.n13 161.3
R1995 VN.n12 VN.n1 161.3
R1996 VN.n11 VN.n10 161.3
R1997 VN.n9 VN.n2 161.3
R1998 VN.n8 VN.n7 161.3
R1999 VN.n6 VN.n3 161.3
R2000 VN.n17 VN.n16 110.267
R2001 VN.n35 VN.n34 110.267
R2002 VN.n5 VN.t0 103.543
R2003 VN.n23 VN.t3 103.543
R2004 VN.n4 VN.t5 71.478
R2005 VN.n16 VN.t2 71.478
R2006 VN.n22 VN.t4 71.478
R2007 VN.n34 VN.t1 71.478
R2008 VN.n5 VN.n4 61.624
R2009 VN.n23 VN.n22 61.624
R2010 VN.n10 VN.n9 52.1486
R2011 VN.n28 VN.n27 52.1486
R2012 VN VN.n35 47.6951
R2013 VN.n10 VN.n1 28.8382
R2014 VN.n28 VN.n19 28.8382
R2015 VN.n8 VN.n3 24.4675
R2016 VN.n9 VN.n8 24.4675
R2017 VN.n14 VN.n1 24.4675
R2018 VN.n15 VN.n14 24.4675
R2019 VN.n27 VN.n26 24.4675
R2020 VN.n26 VN.n21 24.4675
R2021 VN.n33 VN.n32 24.4675
R2022 VN.n32 VN.n19 24.4675
R2023 VN.n4 VN.n3 12.234
R2024 VN.n22 VN.n21 12.234
R2025 VN.n24 VN.n23 5.19435
R2026 VN.n6 VN.n5 5.19435
R2027 VN.n16 VN.n15 0.48984
R2028 VN.n34 VN.n33 0.48984
R2029 VN.n35 VN.n18 0.278367
R2030 VN.n17 VN.n0 0.278367
R2031 VN.n31 VN.n18 0.189894
R2032 VN.n31 VN.n30 0.189894
R2033 VN.n30 VN.n29 0.189894
R2034 VN.n29 VN.n20 0.189894
R2035 VN.n25 VN.n20 0.189894
R2036 VN.n25 VN.n24 0.189894
R2037 VN.n7 VN.n6 0.189894
R2038 VN.n7 VN.n2 0.189894
R2039 VN.n11 VN.n2 0.189894
R2040 VN.n12 VN.n11 0.189894
R2041 VN.n13 VN.n12 0.189894
R2042 VN.n13 VN.n0 0.189894
R2043 VN VN.n17 0.153454
R2044 VDD2.n87 VDD2.n47 289.615
R2045 VDD2.n40 VDD2.n0 289.615
R2046 VDD2.n88 VDD2.n87 185
R2047 VDD2.n86 VDD2.n85 185
R2048 VDD2.n84 VDD2.n50 185
R2049 VDD2.n54 VDD2.n51 185
R2050 VDD2.n79 VDD2.n78 185
R2051 VDD2.n77 VDD2.n76 185
R2052 VDD2.n56 VDD2.n55 185
R2053 VDD2.n71 VDD2.n70 185
R2054 VDD2.n69 VDD2.n68 185
R2055 VDD2.n60 VDD2.n59 185
R2056 VDD2.n63 VDD2.n62 185
R2057 VDD2.n15 VDD2.n14 185
R2058 VDD2.n12 VDD2.n11 185
R2059 VDD2.n21 VDD2.n20 185
R2060 VDD2.n23 VDD2.n22 185
R2061 VDD2.n8 VDD2.n7 185
R2062 VDD2.n29 VDD2.n28 185
R2063 VDD2.n32 VDD2.n31 185
R2064 VDD2.n30 VDD2.n4 185
R2065 VDD2.n37 VDD2.n3 185
R2066 VDD2.n39 VDD2.n38 185
R2067 VDD2.n41 VDD2.n40 185
R2068 VDD2.t4 VDD2.n61 149.524
R2069 VDD2.t5 VDD2.n13 149.524
R2070 VDD2.n87 VDD2.n86 104.615
R2071 VDD2.n86 VDD2.n50 104.615
R2072 VDD2.n54 VDD2.n50 104.615
R2073 VDD2.n78 VDD2.n54 104.615
R2074 VDD2.n78 VDD2.n77 104.615
R2075 VDD2.n77 VDD2.n55 104.615
R2076 VDD2.n70 VDD2.n55 104.615
R2077 VDD2.n70 VDD2.n69 104.615
R2078 VDD2.n69 VDD2.n59 104.615
R2079 VDD2.n62 VDD2.n59 104.615
R2080 VDD2.n14 VDD2.n11 104.615
R2081 VDD2.n21 VDD2.n11 104.615
R2082 VDD2.n22 VDD2.n21 104.615
R2083 VDD2.n22 VDD2.n7 104.615
R2084 VDD2.n29 VDD2.n7 104.615
R2085 VDD2.n31 VDD2.n29 104.615
R2086 VDD2.n31 VDD2.n30 104.615
R2087 VDD2.n30 VDD2.n3 104.615
R2088 VDD2.n39 VDD2.n3 104.615
R2089 VDD2.n40 VDD2.n39 104.615
R2090 VDD2.n46 VDD2.n45 67.3852
R2091 VDD2 VDD2.n93 67.3824
R2092 VDD2.n46 VDD2.n44 54.2135
R2093 VDD2.n62 VDD2.t4 52.3082
R2094 VDD2.n14 VDD2.t5 52.3082
R2095 VDD2.n92 VDD2.n91 52.1611
R2096 VDD2.n92 VDD2.n46 40.3403
R2097 VDD2.n85 VDD2.n84 13.1884
R2098 VDD2.n38 VDD2.n37 13.1884
R2099 VDD2.n88 VDD2.n49 12.8005
R2100 VDD2.n83 VDD2.n51 12.8005
R2101 VDD2.n36 VDD2.n4 12.8005
R2102 VDD2.n41 VDD2.n2 12.8005
R2103 VDD2.n89 VDD2.n47 12.0247
R2104 VDD2.n80 VDD2.n79 12.0247
R2105 VDD2.n33 VDD2.n32 12.0247
R2106 VDD2.n42 VDD2.n0 12.0247
R2107 VDD2.n76 VDD2.n53 11.249
R2108 VDD2.n28 VDD2.n6 11.249
R2109 VDD2.n75 VDD2.n56 10.4732
R2110 VDD2.n27 VDD2.n8 10.4732
R2111 VDD2.n63 VDD2.n61 10.2747
R2112 VDD2.n15 VDD2.n13 10.2747
R2113 VDD2.n72 VDD2.n71 9.69747
R2114 VDD2.n24 VDD2.n23 9.69747
R2115 VDD2.n91 VDD2.n90 9.45567
R2116 VDD2.n44 VDD2.n43 9.45567
R2117 VDD2.n65 VDD2.n64 9.3005
R2118 VDD2.n67 VDD2.n66 9.3005
R2119 VDD2.n58 VDD2.n57 9.3005
R2120 VDD2.n73 VDD2.n72 9.3005
R2121 VDD2.n75 VDD2.n74 9.3005
R2122 VDD2.n53 VDD2.n52 9.3005
R2123 VDD2.n81 VDD2.n80 9.3005
R2124 VDD2.n83 VDD2.n82 9.3005
R2125 VDD2.n90 VDD2.n89 9.3005
R2126 VDD2.n49 VDD2.n48 9.3005
R2127 VDD2.n43 VDD2.n42 9.3005
R2128 VDD2.n2 VDD2.n1 9.3005
R2129 VDD2.n17 VDD2.n16 9.3005
R2130 VDD2.n19 VDD2.n18 9.3005
R2131 VDD2.n10 VDD2.n9 9.3005
R2132 VDD2.n25 VDD2.n24 9.3005
R2133 VDD2.n27 VDD2.n26 9.3005
R2134 VDD2.n6 VDD2.n5 9.3005
R2135 VDD2.n34 VDD2.n33 9.3005
R2136 VDD2.n36 VDD2.n35 9.3005
R2137 VDD2.n68 VDD2.n58 8.92171
R2138 VDD2.n20 VDD2.n10 8.92171
R2139 VDD2.n67 VDD2.n60 8.14595
R2140 VDD2.n19 VDD2.n12 8.14595
R2141 VDD2.n64 VDD2.n63 7.3702
R2142 VDD2.n16 VDD2.n15 7.3702
R2143 VDD2.n64 VDD2.n60 5.81868
R2144 VDD2.n16 VDD2.n12 5.81868
R2145 VDD2.n68 VDD2.n67 5.04292
R2146 VDD2.n20 VDD2.n19 5.04292
R2147 VDD2.n71 VDD2.n58 4.26717
R2148 VDD2.n23 VDD2.n10 4.26717
R2149 VDD2.n72 VDD2.n56 3.49141
R2150 VDD2.n24 VDD2.n8 3.49141
R2151 VDD2.n17 VDD2.n13 2.84303
R2152 VDD2.n65 VDD2.n61 2.84303
R2153 VDD2.n76 VDD2.n75 2.71565
R2154 VDD2.n28 VDD2.n27 2.71565
R2155 VDD2.n93 VDD2.t1 2.27898
R2156 VDD2.n93 VDD2.t2 2.27898
R2157 VDD2.n45 VDD2.t0 2.27898
R2158 VDD2.n45 VDD2.t3 2.27898
R2159 VDD2 VDD2.n92 2.16645
R2160 VDD2.n91 VDD2.n47 1.93989
R2161 VDD2.n79 VDD2.n53 1.93989
R2162 VDD2.n32 VDD2.n6 1.93989
R2163 VDD2.n44 VDD2.n0 1.93989
R2164 VDD2.n89 VDD2.n88 1.16414
R2165 VDD2.n80 VDD2.n51 1.16414
R2166 VDD2.n33 VDD2.n4 1.16414
R2167 VDD2.n42 VDD2.n41 1.16414
R2168 VDD2.n85 VDD2.n49 0.388379
R2169 VDD2.n84 VDD2.n83 0.388379
R2170 VDD2.n37 VDD2.n36 0.388379
R2171 VDD2.n38 VDD2.n2 0.388379
R2172 VDD2.n90 VDD2.n48 0.155672
R2173 VDD2.n82 VDD2.n48 0.155672
R2174 VDD2.n82 VDD2.n81 0.155672
R2175 VDD2.n81 VDD2.n52 0.155672
R2176 VDD2.n74 VDD2.n52 0.155672
R2177 VDD2.n74 VDD2.n73 0.155672
R2178 VDD2.n73 VDD2.n57 0.155672
R2179 VDD2.n66 VDD2.n57 0.155672
R2180 VDD2.n66 VDD2.n65 0.155672
R2181 VDD2.n18 VDD2.n17 0.155672
R2182 VDD2.n18 VDD2.n9 0.155672
R2183 VDD2.n25 VDD2.n9 0.155672
R2184 VDD2.n26 VDD2.n25 0.155672
R2185 VDD2.n26 VDD2.n5 0.155672
R2186 VDD2.n34 VDD2.n5 0.155672
R2187 VDD2.n35 VDD2.n34 0.155672
R2188 VDD2.n35 VDD2.n1 0.155672
R2189 VDD2.n43 VDD2.n1 0.155672
C0 VTAIL VDD1 6.65848f
C1 VTAIL VP 5.48574f
C2 VDD2 VTAIL 6.71254f
C3 VP VDD1 5.41377f
C4 VN VTAIL 5.471529f
C5 VDD2 VDD1 1.5353f
C6 VDD2 VP 0.486053f
C7 VN VDD1 0.151188f
C8 VN VP 6.63442f
C9 VDD2 VN 5.0815f
C10 VDD2 B 5.64821f
C11 VDD1 B 5.799511f
C12 VTAIL B 6.706151f
C13 VN B 13.585031f
C14 VP B 12.280816f
C15 VDD2.n0 B 0.029895f
C16 VDD2.n1 B 0.021579f
C17 VDD2.n2 B 0.011596f
C18 VDD2.n3 B 0.027408f
C19 VDD2.n4 B 0.012278f
C20 VDD2.n5 B 0.021579f
C21 VDD2.n6 B 0.011596f
C22 VDD2.n7 B 0.027408f
C23 VDD2.n8 B 0.012278f
C24 VDD2.n9 B 0.021579f
C25 VDD2.n10 B 0.011596f
C26 VDD2.n11 B 0.027408f
C27 VDD2.n12 B 0.012278f
C28 VDD2.n13 B 0.128177f
C29 VDD2.t5 B 0.045914f
C30 VDD2.n14 B 0.020556f
C31 VDD2.n15 B 0.019375f
C32 VDD2.n16 B 0.011596f
C33 VDD2.n17 B 0.770914f
C34 VDD2.n18 B 0.021579f
C35 VDD2.n19 B 0.011596f
C36 VDD2.n20 B 0.012278f
C37 VDD2.n21 B 0.027408f
C38 VDD2.n22 B 0.027408f
C39 VDD2.n23 B 0.012278f
C40 VDD2.n24 B 0.011596f
C41 VDD2.n25 B 0.021579f
C42 VDD2.n26 B 0.021579f
C43 VDD2.n27 B 0.011596f
C44 VDD2.n28 B 0.012278f
C45 VDD2.n29 B 0.027408f
C46 VDD2.n30 B 0.027408f
C47 VDD2.n31 B 0.027408f
C48 VDD2.n32 B 0.012278f
C49 VDD2.n33 B 0.011596f
C50 VDD2.n34 B 0.021579f
C51 VDD2.n35 B 0.021579f
C52 VDD2.n36 B 0.011596f
C53 VDD2.n37 B 0.011937f
C54 VDD2.n38 B 0.011937f
C55 VDD2.n39 B 0.027408f
C56 VDD2.n40 B 0.058562f
C57 VDD2.n41 B 0.012278f
C58 VDD2.n42 B 0.011596f
C59 VDD2.n43 B 0.054891f
C60 VDD2.n44 B 0.054794f
C61 VDD2.t0 B 0.148187f
C62 VDD2.t3 B 0.148187f
C63 VDD2.n45 B 1.29713f
C64 VDD2.n46 B 2.25735f
C65 VDD2.n47 B 0.029895f
C66 VDD2.n48 B 0.021579f
C67 VDD2.n49 B 0.011596f
C68 VDD2.n50 B 0.027408f
C69 VDD2.n51 B 0.012278f
C70 VDD2.n52 B 0.021579f
C71 VDD2.n53 B 0.011596f
C72 VDD2.n54 B 0.027408f
C73 VDD2.n55 B 0.027408f
C74 VDD2.n56 B 0.012278f
C75 VDD2.n57 B 0.021579f
C76 VDD2.n58 B 0.011596f
C77 VDD2.n59 B 0.027408f
C78 VDD2.n60 B 0.012278f
C79 VDD2.n61 B 0.128177f
C80 VDD2.t4 B 0.045914f
C81 VDD2.n62 B 0.020556f
C82 VDD2.n63 B 0.019375f
C83 VDD2.n64 B 0.011596f
C84 VDD2.n65 B 0.770914f
C85 VDD2.n66 B 0.021579f
C86 VDD2.n67 B 0.011596f
C87 VDD2.n68 B 0.012278f
C88 VDD2.n69 B 0.027408f
C89 VDD2.n70 B 0.027408f
C90 VDD2.n71 B 0.012278f
C91 VDD2.n72 B 0.011596f
C92 VDD2.n73 B 0.021579f
C93 VDD2.n74 B 0.021579f
C94 VDD2.n75 B 0.011596f
C95 VDD2.n76 B 0.012278f
C96 VDD2.n77 B 0.027408f
C97 VDD2.n78 B 0.027408f
C98 VDD2.n79 B 0.012278f
C99 VDD2.n80 B 0.011596f
C100 VDD2.n81 B 0.021579f
C101 VDD2.n82 B 0.021579f
C102 VDD2.n83 B 0.011596f
C103 VDD2.n84 B 0.011937f
C104 VDD2.n85 B 0.011937f
C105 VDD2.n86 B 0.027408f
C106 VDD2.n87 B 0.058562f
C107 VDD2.n88 B 0.012278f
C108 VDD2.n89 B 0.011596f
C109 VDD2.n90 B 0.054891f
C110 VDD2.n91 B 0.0477f
C111 VDD2.n92 B 2.06973f
C112 VDD2.t1 B 0.148187f
C113 VDD2.t2 B 0.148187f
C114 VDD2.n93 B 1.2971f
C115 VN.n0 B 0.029919f
C116 VN.t2 B 1.55717f
C117 VN.n1 B 0.044888f
C118 VN.n2 B 0.022693f
C119 VN.n3 B 0.031854f
C120 VN.t0 B 1.77874f
C121 VN.t5 B 1.55717f
C122 VN.n4 B 0.631952f
C123 VN.n5 B 0.609297f
C124 VN.n6 B 0.24148f
C125 VN.n7 B 0.022693f
C126 VN.n8 B 0.042294f
C127 VN.n9 B 0.040741f
C128 VN.n10 B 0.022921f
C129 VN.n11 B 0.022693f
C130 VN.n12 B 0.022693f
C131 VN.n13 B 0.022693f
C132 VN.n14 B 0.042294f
C133 VN.n15 B 0.021831f
C134 VN.n16 B 0.63492f
C135 VN.n17 B 0.044677f
C136 VN.n18 B 0.029919f
C137 VN.t1 B 1.55717f
C138 VN.n19 B 0.044888f
C139 VN.n20 B 0.022693f
C140 VN.n21 B 0.031854f
C141 VN.t3 B 1.77874f
C142 VN.t4 B 1.55717f
C143 VN.n22 B 0.631952f
C144 VN.n23 B 0.609297f
C145 VN.n24 B 0.24148f
C146 VN.n25 B 0.022693f
C147 VN.n26 B 0.042294f
C148 VN.n27 B 0.040741f
C149 VN.n28 B 0.022921f
C150 VN.n29 B 0.022693f
C151 VN.n30 B 0.022693f
C152 VN.n31 B 0.022693f
C153 VN.n32 B 0.042294f
C154 VN.n33 B 0.021831f
C155 VN.n34 B 0.63492f
C156 VN.n35 B 1.1868f
C157 VDD1.n0 B 0.030449f
C158 VDD1.n1 B 0.021979f
C159 VDD1.n2 B 0.011811f
C160 VDD1.n3 B 0.027916f
C161 VDD1.n4 B 0.012506f
C162 VDD1.n5 B 0.021979f
C163 VDD1.n6 B 0.011811f
C164 VDD1.n7 B 0.027916f
C165 VDD1.n8 B 0.027916f
C166 VDD1.n9 B 0.012506f
C167 VDD1.n10 B 0.021979f
C168 VDD1.n11 B 0.011811f
C169 VDD1.n12 B 0.027916f
C170 VDD1.n13 B 0.012506f
C171 VDD1.n14 B 0.130553f
C172 VDD1.t5 B 0.046766f
C173 VDD1.n15 B 0.020937f
C174 VDD1.n16 B 0.019735f
C175 VDD1.n17 B 0.011811f
C176 VDD1.n18 B 0.78521f
C177 VDD1.n19 B 0.021979f
C178 VDD1.n20 B 0.011811f
C179 VDD1.n21 B 0.012506f
C180 VDD1.n22 B 0.027916f
C181 VDD1.n23 B 0.027916f
C182 VDD1.n24 B 0.012506f
C183 VDD1.n25 B 0.011811f
C184 VDD1.n26 B 0.021979f
C185 VDD1.n27 B 0.021979f
C186 VDD1.n28 B 0.011811f
C187 VDD1.n29 B 0.012506f
C188 VDD1.n30 B 0.027916f
C189 VDD1.n31 B 0.027916f
C190 VDD1.n32 B 0.012506f
C191 VDD1.n33 B 0.011811f
C192 VDD1.n34 B 0.021979f
C193 VDD1.n35 B 0.021979f
C194 VDD1.n36 B 0.011811f
C195 VDD1.n37 B 0.012158f
C196 VDD1.n38 B 0.012158f
C197 VDD1.n39 B 0.027916f
C198 VDD1.n40 B 0.059648f
C199 VDD1.n41 B 0.012506f
C200 VDD1.n42 B 0.011811f
C201 VDD1.n43 B 0.055909f
C202 VDD1.n44 B 0.056505f
C203 VDD1.n45 B 0.030449f
C204 VDD1.n46 B 0.021979f
C205 VDD1.n47 B 0.011811f
C206 VDD1.n48 B 0.027916f
C207 VDD1.n49 B 0.012506f
C208 VDD1.n50 B 0.021979f
C209 VDD1.n51 B 0.011811f
C210 VDD1.n52 B 0.027916f
C211 VDD1.n53 B 0.012506f
C212 VDD1.n54 B 0.021979f
C213 VDD1.n55 B 0.011811f
C214 VDD1.n56 B 0.027916f
C215 VDD1.n57 B 0.012506f
C216 VDD1.n58 B 0.130553f
C217 VDD1.t4 B 0.046766f
C218 VDD1.n59 B 0.020937f
C219 VDD1.n60 B 0.019735f
C220 VDD1.n61 B 0.011811f
C221 VDD1.n62 B 0.78521f
C222 VDD1.n63 B 0.021979f
C223 VDD1.n64 B 0.011811f
C224 VDD1.n65 B 0.012506f
C225 VDD1.n66 B 0.027916f
C226 VDD1.n67 B 0.027916f
C227 VDD1.n68 B 0.012506f
C228 VDD1.n69 B 0.011811f
C229 VDD1.n70 B 0.021979f
C230 VDD1.n71 B 0.021979f
C231 VDD1.n72 B 0.011811f
C232 VDD1.n73 B 0.012506f
C233 VDD1.n74 B 0.027916f
C234 VDD1.n75 B 0.027916f
C235 VDD1.n76 B 0.027916f
C236 VDD1.n77 B 0.012506f
C237 VDD1.n78 B 0.011811f
C238 VDD1.n79 B 0.021979f
C239 VDD1.n80 B 0.021979f
C240 VDD1.n81 B 0.011811f
C241 VDD1.n82 B 0.012158f
C242 VDD1.n83 B 0.012158f
C243 VDD1.n84 B 0.027916f
C244 VDD1.n85 B 0.059648f
C245 VDD1.n86 B 0.012506f
C246 VDD1.n87 B 0.011811f
C247 VDD1.n88 B 0.055909f
C248 VDD1.n89 B 0.05581f
C249 VDD1.t2 B 0.150935f
C250 VDD1.t0 B 0.150935f
C251 VDD1.n90 B 1.32118f
C252 VDD1.n91 B 2.4133f
C253 VDD1.t3 B 0.150935f
C254 VDD1.t1 B 0.150935f
C255 VDD1.n92 B 1.31706f
C256 VDD1.n93 B 2.30512f
C257 VTAIL.t5 B 0.173833f
C258 VTAIL.t0 B 0.173833f
C259 VTAIL.n0 B 1.4513f
C260 VTAIL.n1 B 0.447739f
C261 VTAIL.n2 B 0.035068f
C262 VTAIL.n3 B 0.025314f
C263 VTAIL.n4 B 0.013602f
C264 VTAIL.n5 B 0.032152f
C265 VTAIL.n6 B 0.014403f
C266 VTAIL.n7 B 0.025314f
C267 VTAIL.n8 B 0.013602f
C268 VTAIL.n9 B 0.032152f
C269 VTAIL.n10 B 0.014403f
C270 VTAIL.n11 B 0.025314f
C271 VTAIL.n12 B 0.013602f
C272 VTAIL.n13 B 0.032152f
C273 VTAIL.n14 B 0.014403f
C274 VTAIL.n15 B 0.150359f
C275 VTAIL.t10 B 0.05386f
C276 VTAIL.n16 B 0.024114f
C277 VTAIL.n17 B 0.022729f
C278 VTAIL.n18 B 0.013602f
C279 VTAIL.n19 B 0.90433f
C280 VTAIL.n20 B 0.025314f
C281 VTAIL.n21 B 0.013602f
C282 VTAIL.n22 B 0.014403f
C283 VTAIL.n23 B 0.032152f
C284 VTAIL.n24 B 0.032152f
C285 VTAIL.n25 B 0.014403f
C286 VTAIL.n26 B 0.013602f
C287 VTAIL.n27 B 0.025314f
C288 VTAIL.n28 B 0.025314f
C289 VTAIL.n29 B 0.013602f
C290 VTAIL.n30 B 0.014403f
C291 VTAIL.n31 B 0.032152f
C292 VTAIL.n32 B 0.032152f
C293 VTAIL.n33 B 0.032152f
C294 VTAIL.n34 B 0.014403f
C295 VTAIL.n35 B 0.013602f
C296 VTAIL.n36 B 0.025314f
C297 VTAIL.n37 B 0.025314f
C298 VTAIL.n38 B 0.013602f
C299 VTAIL.n39 B 0.014003f
C300 VTAIL.n40 B 0.014003f
C301 VTAIL.n41 B 0.032152f
C302 VTAIL.n42 B 0.068696f
C303 VTAIL.n43 B 0.014403f
C304 VTAIL.n44 B 0.013602f
C305 VTAIL.n45 B 0.064391f
C306 VTAIL.n46 B 0.038518f
C307 VTAIL.n47 B 0.407114f
C308 VTAIL.t6 B 0.173833f
C309 VTAIL.t8 B 0.173833f
C310 VTAIL.n48 B 1.4513f
C311 VTAIL.n49 B 1.87534f
C312 VTAIL.t2 B 0.173833f
C313 VTAIL.t4 B 0.173833f
C314 VTAIL.n50 B 1.45131f
C315 VTAIL.n51 B 1.87534f
C316 VTAIL.n52 B 0.035068f
C317 VTAIL.n53 B 0.025314f
C318 VTAIL.n54 B 0.013602f
C319 VTAIL.n55 B 0.032152f
C320 VTAIL.n56 B 0.014403f
C321 VTAIL.n57 B 0.025314f
C322 VTAIL.n58 B 0.013602f
C323 VTAIL.n59 B 0.032152f
C324 VTAIL.n60 B 0.032152f
C325 VTAIL.n61 B 0.014403f
C326 VTAIL.n62 B 0.025314f
C327 VTAIL.n63 B 0.013602f
C328 VTAIL.n64 B 0.032152f
C329 VTAIL.n65 B 0.014403f
C330 VTAIL.n66 B 0.150359f
C331 VTAIL.t3 B 0.05386f
C332 VTAIL.n67 B 0.024114f
C333 VTAIL.n68 B 0.022729f
C334 VTAIL.n69 B 0.013602f
C335 VTAIL.n70 B 0.90433f
C336 VTAIL.n71 B 0.025314f
C337 VTAIL.n72 B 0.013602f
C338 VTAIL.n73 B 0.014403f
C339 VTAIL.n74 B 0.032152f
C340 VTAIL.n75 B 0.032152f
C341 VTAIL.n76 B 0.014403f
C342 VTAIL.n77 B 0.013602f
C343 VTAIL.n78 B 0.025314f
C344 VTAIL.n79 B 0.025314f
C345 VTAIL.n80 B 0.013602f
C346 VTAIL.n81 B 0.014403f
C347 VTAIL.n82 B 0.032152f
C348 VTAIL.n83 B 0.032152f
C349 VTAIL.n84 B 0.014403f
C350 VTAIL.n85 B 0.013602f
C351 VTAIL.n86 B 0.025314f
C352 VTAIL.n87 B 0.025314f
C353 VTAIL.n88 B 0.013602f
C354 VTAIL.n89 B 0.014003f
C355 VTAIL.n90 B 0.014003f
C356 VTAIL.n91 B 0.032152f
C357 VTAIL.n92 B 0.068696f
C358 VTAIL.n93 B 0.014403f
C359 VTAIL.n94 B 0.013602f
C360 VTAIL.n95 B 0.064391f
C361 VTAIL.n96 B 0.038518f
C362 VTAIL.n97 B 0.407114f
C363 VTAIL.t9 B 0.173833f
C364 VTAIL.t7 B 0.173833f
C365 VTAIL.n98 B 1.45131f
C366 VTAIL.n99 B 0.614907f
C367 VTAIL.n100 B 0.035068f
C368 VTAIL.n101 B 0.025314f
C369 VTAIL.n102 B 0.013602f
C370 VTAIL.n103 B 0.032152f
C371 VTAIL.n104 B 0.014403f
C372 VTAIL.n105 B 0.025314f
C373 VTAIL.n106 B 0.013602f
C374 VTAIL.n107 B 0.032152f
C375 VTAIL.n108 B 0.032152f
C376 VTAIL.n109 B 0.014403f
C377 VTAIL.n110 B 0.025314f
C378 VTAIL.n111 B 0.013602f
C379 VTAIL.n112 B 0.032152f
C380 VTAIL.n113 B 0.014403f
C381 VTAIL.n114 B 0.150359f
C382 VTAIL.t11 B 0.05386f
C383 VTAIL.n115 B 0.024114f
C384 VTAIL.n116 B 0.022729f
C385 VTAIL.n117 B 0.013602f
C386 VTAIL.n118 B 0.90433f
C387 VTAIL.n119 B 0.025314f
C388 VTAIL.n120 B 0.013602f
C389 VTAIL.n121 B 0.014403f
C390 VTAIL.n122 B 0.032152f
C391 VTAIL.n123 B 0.032152f
C392 VTAIL.n124 B 0.014403f
C393 VTAIL.n125 B 0.013602f
C394 VTAIL.n126 B 0.025314f
C395 VTAIL.n127 B 0.025314f
C396 VTAIL.n128 B 0.013602f
C397 VTAIL.n129 B 0.014403f
C398 VTAIL.n130 B 0.032152f
C399 VTAIL.n131 B 0.032152f
C400 VTAIL.n132 B 0.014403f
C401 VTAIL.n133 B 0.013602f
C402 VTAIL.n134 B 0.025314f
C403 VTAIL.n135 B 0.025314f
C404 VTAIL.n136 B 0.013602f
C405 VTAIL.n137 B 0.014003f
C406 VTAIL.n138 B 0.014003f
C407 VTAIL.n139 B 0.032152f
C408 VTAIL.n140 B 0.068696f
C409 VTAIL.n141 B 0.014403f
C410 VTAIL.n142 B 0.013602f
C411 VTAIL.n143 B 0.064391f
C412 VTAIL.n144 B 0.038518f
C413 VTAIL.n145 B 1.43831f
C414 VTAIL.n146 B 0.035068f
C415 VTAIL.n147 B 0.025314f
C416 VTAIL.n148 B 0.013602f
C417 VTAIL.n149 B 0.032152f
C418 VTAIL.n150 B 0.014403f
C419 VTAIL.n151 B 0.025314f
C420 VTAIL.n152 B 0.013602f
C421 VTAIL.n153 B 0.032152f
C422 VTAIL.n154 B 0.014403f
C423 VTAIL.n155 B 0.025314f
C424 VTAIL.n156 B 0.013602f
C425 VTAIL.n157 B 0.032152f
C426 VTAIL.n158 B 0.014403f
C427 VTAIL.n159 B 0.150359f
C428 VTAIL.t1 B 0.05386f
C429 VTAIL.n160 B 0.024114f
C430 VTAIL.n161 B 0.022729f
C431 VTAIL.n162 B 0.013602f
C432 VTAIL.n163 B 0.90433f
C433 VTAIL.n164 B 0.025314f
C434 VTAIL.n165 B 0.013602f
C435 VTAIL.n166 B 0.014403f
C436 VTAIL.n167 B 0.032152f
C437 VTAIL.n168 B 0.032152f
C438 VTAIL.n169 B 0.014403f
C439 VTAIL.n170 B 0.013602f
C440 VTAIL.n171 B 0.025314f
C441 VTAIL.n172 B 0.025314f
C442 VTAIL.n173 B 0.013602f
C443 VTAIL.n174 B 0.014403f
C444 VTAIL.n175 B 0.032152f
C445 VTAIL.n176 B 0.032152f
C446 VTAIL.n177 B 0.032152f
C447 VTAIL.n178 B 0.014403f
C448 VTAIL.n179 B 0.013602f
C449 VTAIL.n180 B 0.025314f
C450 VTAIL.n181 B 0.025314f
C451 VTAIL.n182 B 0.013602f
C452 VTAIL.n183 B 0.014003f
C453 VTAIL.n184 B 0.014003f
C454 VTAIL.n185 B 0.032152f
C455 VTAIL.n186 B 0.068696f
C456 VTAIL.n187 B 0.014403f
C457 VTAIL.n188 B 0.013602f
C458 VTAIL.n189 B 0.064391f
C459 VTAIL.n190 B 0.038518f
C460 VTAIL.n191 B 1.37626f
C461 VP.n0 B 0.030497f
C462 VP.t5 B 1.58728f
C463 VP.n1 B 0.045756f
C464 VP.n2 B 0.023132f
C465 VP.n3 B 0.03247f
C466 VP.n4 B 0.023132f
C467 VP.n5 B 0.023365f
C468 VP.n6 B 0.023132f
C469 VP.t1 B 1.58728f
C470 VP.n7 B 0.647195f
C471 VP.n8 B 0.030497f
C472 VP.t4 B 1.58728f
C473 VP.n9 B 0.045756f
C474 VP.n10 B 0.023132f
C475 VP.n11 B 0.03247f
C476 VP.t0 B 1.81313f
C477 VP.t2 B 1.58728f
C478 VP.n12 B 0.64417f
C479 VP.n13 B 0.621076f
C480 VP.n14 B 0.246148f
C481 VP.n15 B 0.023132f
C482 VP.n16 B 0.043112f
C483 VP.n17 B 0.041528f
C484 VP.n18 B 0.023365f
C485 VP.n19 B 0.023132f
C486 VP.n20 B 0.023132f
C487 VP.n21 B 0.023132f
C488 VP.n22 B 0.043112f
C489 VP.n23 B 0.022253f
C490 VP.n24 B 0.647195f
C491 VP.n25 B 1.19721f
C492 VP.n26 B 1.21475f
C493 VP.n27 B 0.030497f
C494 VP.n28 B 0.022253f
C495 VP.n29 B 0.043112f
C496 VP.n30 B 0.045756f
C497 VP.n31 B 0.023132f
C498 VP.n32 B 0.023132f
C499 VP.n33 B 0.023132f
C500 VP.n34 B 0.041528f
C501 VP.n35 B 0.043112f
C502 VP.t3 B 1.58728f
C503 VP.n36 B 0.571481f
C504 VP.n37 B 0.03247f
C505 VP.n38 B 0.023132f
C506 VP.n39 B 0.023132f
C507 VP.n40 B 0.023132f
C508 VP.n41 B 0.043112f
C509 VP.n42 B 0.041528f
C510 VP.n43 B 0.023365f
C511 VP.n44 B 0.023132f
C512 VP.n45 B 0.023132f
C513 VP.n46 B 0.023132f
C514 VP.n47 B 0.043112f
C515 VP.n48 B 0.022253f
C516 VP.n49 B 0.647195f
C517 VP.n50 B 0.045541f
.ends

