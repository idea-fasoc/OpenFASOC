* NGSPICE file created from diff_pair_sample_0551.ext - technology: sky130A

.subckt diff_pair_sample_0551 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X1 VTAIL.t3 VN.t0 VDD2.t7 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X2 B.t11 B.t9 B.t10 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=0 ps=0 w=15.95 l=1.17
X3 VTAIL.t9 VP.t1 VDD1.t6 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X4 VDD2.t6 VN.t1 VTAIL.t5 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=6.2205 ps=32.68 w=15.95 l=1.17
X5 B.t8 B.t6 B.t7 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=0 ps=0 w=15.95 l=1.17
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X7 B.t5 B.t3 B.t4 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=0 ps=0 w=15.95 l=1.17
X8 VTAIL.t2 VN.t3 VDD2.t4 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X9 B.t2 B.t0 B.t1 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=0 ps=0 w=15.95 l=1.17
X10 VDD1.t5 VP.t2 VTAIL.t11 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=6.2205 ps=32.68 w=15.95 l=1.17
X11 VTAIL.t15 VP.t3 VDD1.t4 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=2.63175 ps=16.28 w=15.95 l=1.17
X12 VDD2.t3 VN.t4 VTAIL.t4 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X13 VTAIL.t10 VP.t4 VDD1.t3 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=2.63175 ps=16.28 w=15.95 l=1.17
X14 VTAIL.t0 VN.t5 VDD2.t2 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=2.63175 ps=16.28 w=15.95 l=1.17
X15 VDD1.t2 VP.t5 VTAIL.t14 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X16 VTAIL.t6 VN.t6 VDD2.t1 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=6.2205 pd=32.68 as=2.63175 ps=16.28 w=15.95 l=1.17
X17 VDD1.t1 VP.t6 VTAIL.t13 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=6.2205 ps=32.68 w=15.95 l=1.17
X18 VTAIL.t12 VP.t7 VDD1.t0 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=2.63175 ps=16.28 w=15.95 l=1.17
X19 VDD2.t0 VN.t7 VTAIL.t7 w_n2470_n4158# sky130_fd_pr__pfet_01v8 ad=2.63175 pd=16.28 as=6.2205 ps=32.68 w=15.95 l=1.17
R0 VP.n10 VP.t4 358.652
R1 VP.n5 VP.t3 328.543
R2 VP.n3 VP.t0 328.543
R3 VP.n32 VP.t1 328.543
R4 VP.n39 VP.t2 328.543
R5 VP.n21 VP.t6 328.543
R6 VP.n14 VP.t7 328.543
R7 VP.n9 VP.t5 328.543
R8 VP.n23 VP.n5 173.534
R9 VP.n40 VP.n39 173.534
R10 VP.n22 VP.n21 173.534
R11 VP.n12 VP.n11 161.3
R12 VP.n13 VP.n8 161.3
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n7 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n20 VP.n6 161.3
R17 VP.n38 VP.n0 161.3
R18 VP.n37 VP.n36 161.3
R19 VP.n35 VP.n1 161.3
R20 VP.n34 VP.n33 161.3
R21 VP.n31 VP.n2 161.3
R22 VP.n30 VP.n29 161.3
R23 VP.n28 VP.n27 161.3
R24 VP.n26 VP.n4 161.3
R25 VP.n25 VP.n24 161.3
R26 VP.n10 VP.n9 51.4127
R27 VP.n23 VP.n22 47.0763
R28 VP.n26 VP.n25 40.4934
R29 VP.n27 VP.n26 40.4934
R30 VP.n31 VP.n30 40.4934
R31 VP.n33 VP.n31 40.4934
R32 VP.n37 VP.n1 40.4934
R33 VP.n38 VP.n37 40.4934
R34 VP.n20 VP.n19 40.4934
R35 VP.n19 VP.n7 40.4934
R36 VP.n15 VP.n13 40.4934
R37 VP.n13 VP.n12 40.4934
R38 VP.n11 VP.n10 27.0291
R39 VP.n25 VP.n5 12.234
R40 VP.n27 VP.n3 12.234
R41 VP.n30 VP.n3 12.234
R42 VP.n33 VP.n32 12.234
R43 VP.n32 VP.n1 12.234
R44 VP.n39 VP.n38 12.234
R45 VP.n21 VP.n20 12.234
R46 VP.n15 VP.n14 12.234
R47 VP.n14 VP.n7 12.234
R48 VP.n12 VP.n9 12.234
R49 VP.n11 VP.n8 0.189894
R50 VP.n16 VP.n8 0.189894
R51 VP.n17 VP.n16 0.189894
R52 VP.n18 VP.n17 0.189894
R53 VP.n18 VP.n6 0.189894
R54 VP.n22 VP.n6 0.189894
R55 VP.n24 VP.n23 0.189894
R56 VP.n24 VP.n4 0.189894
R57 VP.n28 VP.n4 0.189894
R58 VP.n29 VP.n28 0.189894
R59 VP.n29 VP.n2 0.189894
R60 VP.n34 VP.n2 0.189894
R61 VP.n35 VP.n34 0.189894
R62 VP.n36 VP.n35 0.189894
R63 VP.n36 VP.n0 0.189894
R64 VP.n40 VP.n0 0.189894
R65 VP VP.n40 0.0516364
R66 VTAIL.n11 VTAIL.t10 59.8434
R67 VTAIL.n10 VTAIL.t5 59.8434
R68 VTAIL.n7 VTAIL.t6 59.8434
R69 VTAIL.n14 VTAIL.t13 59.8433
R70 VTAIL.n15 VTAIL.t7 59.8433
R71 VTAIL.n2 VTAIL.t0 59.8433
R72 VTAIL.n3 VTAIL.t11 59.8433
R73 VTAIL.n6 VTAIL.t15 59.8433
R74 VTAIL.n13 VTAIL.n12 57.8056
R75 VTAIL.n9 VTAIL.n8 57.8056
R76 VTAIL.n1 VTAIL.n0 57.8053
R77 VTAIL.n5 VTAIL.n4 57.8053
R78 VTAIL.n15 VTAIL.n14 27.41
R79 VTAIL.n7 VTAIL.n6 27.41
R80 VTAIL.n0 VTAIL.t1 2.03843
R81 VTAIL.n0 VTAIL.t3 2.03843
R82 VTAIL.n4 VTAIL.t8 2.03843
R83 VTAIL.n4 VTAIL.t9 2.03843
R84 VTAIL.n12 VTAIL.t14 2.03843
R85 VTAIL.n12 VTAIL.t12 2.03843
R86 VTAIL.n8 VTAIL.t4 2.03843
R87 VTAIL.n8 VTAIL.t2 2.03843
R88 VTAIL.n9 VTAIL.n7 1.2936
R89 VTAIL.n10 VTAIL.n9 1.2936
R90 VTAIL.n13 VTAIL.n11 1.2936
R91 VTAIL.n14 VTAIL.n13 1.2936
R92 VTAIL.n6 VTAIL.n5 1.2936
R93 VTAIL.n5 VTAIL.n3 1.2936
R94 VTAIL.n2 VTAIL.n1 1.2936
R95 VTAIL VTAIL.n15 1.23541
R96 VTAIL.n11 VTAIL.n10 0.470328
R97 VTAIL.n3 VTAIL.n2 0.470328
R98 VTAIL VTAIL.n1 0.0586897
R99 VDD1 VDD1.n0 75.1891
R100 VDD1.n3 VDD1.n2 75.0753
R101 VDD1.n3 VDD1.n1 75.0753
R102 VDD1.n5 VDD1.n4 74.4842
R103 VDD1.n5 VDD1.n3 43.8673
R104 VDD1.n4 VDD1.t0 2.03843
R105 VDD1.n4 VDD1.t1 2.03843
R106 VDD1.n0 VDD1.t3 2.03843
R107 VDD1.n0 VDD1.t2 2.03843
R108 VDD1.n2 VDD1.t6 2.03843
R109 VDD1.n2 VDD1.t5 2.03843
R110 VDD1.n1 VDD1.t4 2.03843
R111 VDD1.n1 VDD1.t7 2.03843
R112 VDD1 VDD1.n5 0.588862
R113 VN.n4 VN.t5 358.652
R114 VN.n22 VN.t1 358.652
R115 VN.n3 VN.t2 328.543
R116 VN.n8 VN.t0 328.543
R117 VN.n15 VN.t7 328.543
R118 VN.n21 VN.t3 328.543
R119 VN.n20 VN.t4 328.543
R120 VN.n32 VN.t6 328.543
R121 VN.n16 VN.n15 173.534
R122 VN.n33 VN.n32 173.534
R123 VN.n31 VN.n17 161.3
R124 VN.n30 VN.n29 161.3
R125 VN.n28 VN.n18 161.3
R126 VN.n27 VN.n26 161.3
R127 VN.n25 VN.n19 161.3
R128 VN.n24 VN.n23 161.3
R129 VN.n14 VN.n0 161.3
R130 VN.n13 VN.n12 161.3
R131 VN.n11 VN.n1 161.3
R132 VN.n10 VN.n9 161.3
R133 VN.n7 VN.n2 161.3
R134 VN.n6 VN.n5 161.3
R135 VN.n4 VN.n3 51.4127
R136 VN.n22 VN.n21 51.4127
R137 VN VN.n33 47.4569
R138 VN.n7 VN.n6 40.4934
R139 VN.n9 VN.n7 40.4934
R140 VN.n13 VN.n1 40.4934
R141 VN.n14 VN.n13 40.4934
R142 VN.n25 VN.n24 40.4934
R143 VN.n26 VN.n25 40.4934
R144 VN.n30 VN.n18 40.4934
R145 VN.n31 VN.n30 40.4934
R146 VN.n23 VN.n22 27.0291
R147 VN.n5 VN.n4 27.0291
R148 VN.n6 VN.n3 12.234
R149 VN.n9 VN.n8 12.234
R150 VN.n8 VN.n1 12.234
R151 VN.n15 VN.n14 12.234
R152 VN.n24 VN.n21 12.234
R153 VN.n20 VN.n18 12.234
R154 VN.n26 VN.n20 12.234
R155 VN.n32 VN.n31 12.234
R156 VN.n33 VN.n17 0.189894
R157 VN.n29 VN.n17 0.189894
R158 VN.n29 VN.n28 0.189894
R159 VN.n28 VN.n27 0.189894
R160 VN.n27 VN.n19 0.189894
R161 VN.n23 VN.n19 0.189894
R162 VN.n5 VN.n2 0.189894
R163 VN.n10 VN.n2 0.189894
R164 VN.n11 VN.n10 0.189894
R165 VN.n12 VN.n11 0.189894
R166 VN.n12 VN.n0 0.189894
R167 VN.n16 VN.n0 0.189894
R168 VN VN.n16 0.0516364
R169 VDD2.n2 VDD2.n1 75.0753
R170 VDD2.n2 VDD2.n0 75.0753
R171 VDD2 VDD2.n5 75.0726
R172 VDD2.n4 VDD2.n3 74.4844
R173 VDD2.n4 VDD2.n2 43.2843
R174 VDD2.n5 VDD2.t4 2.03843
R175 VDD2.n5 VDD2.t6 2.03843
R176 VDD2.n3 VDD2.t1 2.03843
R177 VDD2.n3 VDD2.t3 2.03843
R178 VDD2.n1 VDD2.t7 2.03843
R179 VDD2.n1 VDD2.t0 2.03843
R180 VDD2.n0 VDD2.t2 2.03843
R181 VDD2.n0 VDD2.t5 2.03843
R182 VDD2 VDD2.n4 0.705241
R183 B.n499 B.n498 585
R184 B.n500 B.n79 585
R185 B.n502 B.n501 585
R186 B.n503 B.n78 585
R187 B.n505 B.n504 585
R188 B.n506 B.n77 585
R189 B.n508 B.n507 585
R190 B.n509 B.n76 585
R191 B.n511 B.n510 585
R192 B.n512 B.n75 585
R193 B.n514 B.n513 585
R194 B.n515 B.n74 585
R195 B.n517 B.n516 585
R196 B.n518 B.n73 585
R197 B.n520 B.n519 585
R198 B.n521 B.n72 585
R199 B.n523 B.n522 585
R200 B.n524 B.n71 585
R201 B.n526 B.n525 585
R202 B.n527 B.n70 585
R203 B.n529 B.n528 585
R204 B.n530 B.n69 585
R205 B.n532 B.n531 585
R206 B.n533 B.n68 585
R207 B.n535 B.n534 585
R208 B.n536 B.n67 585
R209 B.n538 B.n537 585
R210 B.n539 B.n66 585
R211 B.n541 B.n540 585
R212 B.n542 B.n65 585
R213 B.n544 B.n543 585
R214 B.n545 B.n64 585
R215 B.n547 B.n546 585
R216 B.n548 B.n63 585
R217 B.n550 B.n549 585
R218 B.n551 B.n62 585
R219 B.n553 B.n552 585
R220 B.n554 B.n61 585
R221 B.n556 B.n555 585
R222 B.n557 B.n60 585
R223 B.n559 B.n558 585
R224 B.n560 B.n59 585
R225 B.n562 B.n561 585
R226 B.n563 B.n58 585
R227 B.n565 B.n564 585
R228 B.n566 B.n57 585
R229 B.n568 B.n567 585
R230 B.n569 B.n56 585
R231 B.n571 B.n570 585
R232 B.n572 B.n55 585
R233 B.n574 B.n573 585
R234 B.n575 B.n51 585
R235 B.n577 B.n576 585
R236 B.n578 B.n50 585
R237 B.n580 B.n579 585
R238 B.n581 B.n49 585
R239 B.n583 B.n582 585
R240 B.n584 B.n48 585
R241 B.n586 B.n585 585
R242 B.n587 B.n47 585
R243 B.n589 B.n588 585
R244 B.n590 B.n46 585
R245 B.n592 B.n591 585
R246 B.n594 B.n43 585
R247 B.n596 B.n595 585
R248 B.n597 B.n42 585
R249 B.n599 B.n598 585
R250 B.n600 B.n41 585
R251 B.n602 B.n601 585
R252 B.n603 B.n40 585
R253 B.n605 B.n604 585
R254 B.n606 B.n39 585
R255 B.n608 B.n607 585
R256 B.n609 B.n38 585
R257 B.n611 B.n610 585
R258 B.n612 B.n37 585
R259 B.n614 B.n613 585
R260 B.n615 B.n36 585
R261 B.n617 B.n616 585
R262 B.n618 B.n35 585
R263 B.n620 B.n619 585
R264 B.n621 B.n34 585
R265 B.n623 B.n622 585
R266 B.n624 B.n33 585
R267 B.n626 B.n625 585
R268 B.n627 B.n32 585
R269 B.n629 B.n628 585
R270 B.n630 B.n31 585
R271 B.n632 B.n631 585
R272 B.n633 B.n30 585
R273 B.n635 B.n634 585
R274 B.n636 B.n29 585
R275 B.n638 B.n637 585
R276 B.n639 B.n28 585
R277 B.n641 B.n640 585
R278 B.n642 B.n27 585
R279 B.n644 B.n643 585
R280 B.n645 B.n26 585
R281 B.n647 B.n646 585
R282 B.n648 B.n25 585
R283 B.n650 B.n649 585
R284 B.n651 B.n24 585
R285 B.n653 B.n652 585
R286 B.n654 B.n23 585
R287 B.n656 B.n655 585
R288 B.n657 B.n22 585
R289 B.n659 B.n658 585
R290 B.n660 B.n21 585
R291 B.n662 B.n661 585
R292 B.n663 B.n20 585
R293 B.n665 B.n664 585
R294 B.n666 B.n19 585
R295 B.n668 B.n667 585
R296 B.n669 B.n18 585
R297 B.n671 B.n670 585
R298 B.n672 B.n17 585
R299 B.n497 B.n80 585
R300 B.n496 B.n495 585
R301 B.n494 B.n81 585
R302 B.n493 B.n492 585
R303 B.n491 B.n82 585
R304 B.n490 B.n489 585
R305 B.n488 B.n83 585
R306 B.n487 B.n486 585
R307 B.n485 B.n84 585
R308 B.n484 B.n483 585
R309 B.n482 B.n85 585
R310 B.n481 B.n480 585
R311 B.n479 B.n86 585
R312 B.n478 B.n477 585
R313 B.n476 B.n87 585
R314 B.n475 B.n474 585
R315 B.n473 B.n88 585
R316 B.n472 B.n471 585
R317 B.n470 B.n89 585
R318 B.n469 B.n468 585
R319 B.n467 B.n90 585
R320 B.n466 B.n465 585
R321 B.n464 B.n91 585
R322 B.n463 B.n462 585
R323 B.n461 B.n92 585
R324 B.n460 B.n459 585
R325 B.n458 B.n93 585
R326 B.n457 B.n456 585
R327 B.n455 B.n94 585
R328 B.n454 B.n453 585
R329 B.n452 B.n95 585
R330 B.n451 B.n450 585
R331 B.n449 B.n96 585
R332 B.n448 B.n447 585
R333 B.n446 B.n97 585
R334 B.n445 B.n444 585
R335 B.n443 B.n98 585
R336 B.n442 B.n441 585
R337 B.n440 B.n99 585
R338 B.n439 B.n438 585
R339 B.n437 B.n100 585
R340 B.n436 B.n435 585
R341 B.n434 B.n101 585
R342 B.n433 B.n432 585
R343 B.n431 B.n102 585
R344 B.n430 B.n429 585
R345 B.n428 B.n103 585
R346 B.n427 B.n426 585
R347 B.n425 B.n104 585
R348 B.n424 B.n423 585
R349 B.n422 B.n105 585
R350 B.n421 B.n420 585
R351 B.n419 B.n106 585
R352 B.n418 B.n417 585
R353 B.n416 B.n107 585
R354 B.n415 B.n414 585
R355 B.n413 B.n108 585
R356 B.n412 B.n411 585
R357 B.n410 B.n109 585
R358 B.n409 B.n408 585
R359 B.n407 B.n110 585
R360 B.n232 B.n231 585
R361 B.n233 B.n172 585
R362 B.n235 B.n234 585
R363 B.n236 B.n171 585
R364 B.n238 B.n237 585
R365 B.n239 B.n170 585
R366 B.n241 B.n240 585
R367 B.n242 B.n169 585
R368 B.n244 B.n243 585
R369 B.n245 B.n168 585
R370 B.n247 B.n246 585
R371 B.n248 B.n167 585
R372 B.n250 B.n249 585
R373 B.n251 B.n166 585
R374 B.n253 B.n252 585
R375 B.n254 B.n165 585
R376 B.n256 B.n255 585
R377 B.n257 B.n164 585
R378 B.n259 B.n258 585
R379 B.n260 B.n163 585
R380 B.n262 B.n261 585
R381 B.n263 B.n162 585
R382 B.n265 B.n264 585
R383 B.n266 B.n161 585
R384 B.n268 B.n267 585
R385 B.n269 B.n160 585
R386 B.n271 B.n270 585
R387 B.n272 B.n159 585
R388 B.n274 B.n273 585
R389 B.n275 B.n158 585
R390 B.n277 B.n276 585
R391 B.n278 B.n157 585
R392 B.n280 B.n279 585
R393 B.n281 B.n156 585
R394 B.n283 B.n282 585
R395 B.n284 B.n155 585
R396 B.n286 B.n285 585
R397 B.n287 B.n154 585
R398 B.n289 B.n288 585
R399 B.n290 B.n153 585
R400 B.n292 B.n291 585
R401 B.n293 B.n152 585
R402 B.n295 B.n294 585
R403 B.n296 B.n151 585
R404 B.n298 B.n297 585
R405 B.n299 B.n150 585
R406 B.n301 B.n300 585
R407 B.n302 B.n149 585
R408 B.n304 B.n303 585
R409 B.n305 B.n148 585
R410 B.n307 B.n306 585
R411 B.n308 B.n147 585
R412 B.n310 B.n309 585
R413 B.n312 B.n144 585
R414 B.n314 B.n313 585
R415 B.n315 B.n143 585
R416 B.n317 B.n316 585
R417 B.n318 B.n142 585
R418 B.n320 B.n319 585
R419 B.n321 B.n141 585
R420 B.n323 B.n322 585
R421 B.n324 B.n140 585
R422 B.n326 B.n325 585
R423 B.n328 B.n327 585
R424 B.n329 B.n136 585
R425 B.n331 B.n330 585
R426 B.n332 B.n135 585
R427 B.n334 B.n333 585
R428 B.n335 B.n134 585
R429 B.n337 B.n336 585
R430 B.n338 B.n133 585
R431 B.n340 B.n339 585
R432 B.n341 B.n132 585
R433 B.n343 B.n342 585
R434 B.n344 B.n131 585
R435 B.n346 B.n345 585
R436 B.n347 B.n130 585
R437 B.n349 B.n348 585
R438 B.n350 B.n129 585
R439 B.n352 B.n351 585
R440 B.n353 B.n128 585
R441 B.n355 B.n354 585
R442 B.n356 B.n127 585
R443 B.n358 B.n357 585
R444 B.n359 B.n126 585
R445 B.n361 B.n360 585
R446 B.n362 B.n125 585
R447 B.n364 B.n363 585
R448 B.n365 B.n124 585
R449 B.n367 B.n366 585
R450 B.n368 B.n123 585
R451 B.n370 B.n369 585
R452 B.n371 B.n122 585
R453 B.n373 B.n372 585
R454 B.n374 B.n121 585
R455 B.n376 B.n375 585
R456 B.n377 B.n120 585
R457 B.n379 B.n378 585
R458 B.n380 B.n119 585
R459 B.n382 B.n381 585
R460 B.n383 B.n118 585
R461 B.n385 B.n384 585
R462 B.n386 B.n117 585
R463 B.n388 B.n387 585
R464 B.n389 B.n116 585
R465 B.n391 B.n390 585
R466 B.n392 B.n115 585
R467 B.n394 B.n393 585
R468 B.n395 B.n114 585
R469 B.n397 B.n396 585
R470 B.n398 B.n113 585
R471 B.n400 B.n399 585
R472 B.n401 B.n112 585
R473 B.n403 B.n402 585
R474 B.n404 B.n111 585
R475 B.n406 B.n405 585
R476 B.n230 B.n173 585
R477 B.n229 B.n228 585
R478 B.n227 B.n174 585
R479 B.n226 B.n225 585
R480 B.n224 B.n175 585
R481 B.n223 B.n222 585
R482 B.n221 B.n176 585
R483 B.n220 B.n219 585
R484 B.n218 B.n177 585
R485 B.n217 B.n216 585
R486 B.n215 B.n178 585
R487 B.n214 B.n213 585
R488 B.n212 B.n179 585
R489 B.n211 B.n210 585
R490 B.n209 B.n180 585
R491 B.n208 B.n207 585
R492 B.n206 B.n181 585
R493 B.n205 B.n204 585
R494 B.n203 B.n182 585
R495 B.n202 B.n201 585
R496 B.n200 B.n183 585
R497 B.n199 B.n198 585
R498 B.n197 B.n184 585
R499 B.n196 B.n195 585
R500 B.n194 B.n185 585
R501 B.n193 B.n192 585
R502 B.n191 B.n186 585
R503 B.n190 B.n189 585
R504 B.n188 B.n187 585
R505 B.n2 B.n0 585
R506 B.n717 B.n1 585
R507 B.n716 B.n715 585
R508 B.n714 B.n3 585
R509 B.n713 B.n712 585
R510 B.n711 B.n4 585
R511 B.n710 B.n709 585
R512 B.n708 B.n5 585
R513 B.n707 B.n706 585
R514 B.n705 B.n6 585
R515 B.n704 B.n703 585
R516 B.n702 B.n7 585
R517 B.n701 B.n700 585
R518 B.n699 B.n8 585
R519 B.n698 B.n697 585
R520 B.n696 B.n9 585
R521 B.n695 B.n694 585
R522 B.n693 B.n10 585
R523 B.n692 B.n691 585
R524 B.n690 B.n11 585
R525 B.n689 B.n688 585
R526 B.n687 B.n12 585
R527 B.n686 B.n685 585
R528 B.n684 B.n13 585
R529 B.n683 B.n682 585
R530 B.n681 B.n14 585
R531 B.n680 B.n679 585
R532 B.n678 B.n15 585
R533 B.n677 B.n676 585
R534 B.n675 B.n16 585
R535 B.n674 B.n673 585
R536 B.n719 B.n718 585
R537 B.n137 B.t9 532.5
R538 B.n145 B.t6 532.5
R539 B.n44 B.t3 532.5
R540 B.n52 B.t0 532.5
R541 B.n231 B.n230 530.939
R542 B.n674 B.n17 530.939
R543 B.n405 B.n110 530.939
R544 B.n499 B.n80 530.939
R545 B.n230 B.n229 163.367
R546 B.n229 B.n174 163.367
R547 B.n225 B.n174 163.367
R548 B.n225 B.n224 163.367
R549 B.n224 B.n223 163.367
R550 B.n223 B.n176 163.367
R551 B.n219 B.n176 163.367
R552 B.n219 B.n218 163.367
R553 B.n218 B.n217 163.367
R554 B.n217 B.n178 163.367
R555 B.n213 B.n178 163.367
R556 B.n213 B.n212 163.367
R557 B.n212 B.n211 163.367
R558 B.n211 B.n180 163.367
R559 B.n207 B.n180 163.367
R560 B.n207 B.n206 163.367
R561 B.n206 B.n205 163.367
R562 B.n205 B.n182 163.367
R563 B.n201 B.n182 163.367
R564 B.n201 B.n200 163.367
R565 B.n200 B.n199 163.367
R566 B.n199 B.n184 163.367
R567 B.n195 B.n184 163.367
R568 B.n195 B.n194 163.367
R569 B.n194 B.n193 163.367
R570 B.n193 B.n186 163.367
R571 B.n189 B.n186 163.367
R572 B.n189 B.n188 163.367
R573 B.n188 B.n2 163.367
R574 B.n718 B.n2 163.367
R575 B.n718 B.n717 163.367
R576 B.n717 B.n716 163.367
R577 B.n716 B.n3 163.367
R578 B.n712 B.n3 163.367
R579 B.n712 B.n711 163.367
R580 B.n711 B.n710 163.367
R581 B.n710 B.n5 163.367
R582 B.n706 B.n5 163.367
R583 B.n706 B.n705 163.367
R584 B.n705 B.n704 163.367
R585 B.n704 B.n7 163.367
R586 B.n700 B.n7 163.367
R587 B.n700 B.n699 163.367
R588 B.n699 B.n698 163.367
R589 B.n698 B.n9 163.367
R590 B.n694 B.n9 163.367
R591 B.n694 B.n693 163.367
R592 B.n693 B.n692 163.367
R593 B.n692 B.n11 163.367
R594 B.n688 B.n11 163.367
R595 B.n688 B.n687 163.367
R596 B.n687 B.n686 163.367
R597 B.n686 B.n13 163.367
R598 B.n682 B.n13 163.367
R599 B.n682 B.n681 163.367
R600 B.n681 B.n680 163.367
R601 B.n680 B.n15 163.367
R602 B.n676 B.n15 163.367
R603 B.n676 B.n675 163.367
R604 B.n675 B.n674 163.367
R605 B.n231 B.n172 163.367
R606 B.n235 B.n172 163.367
R607 B.n236 B.n235 163.367
R608 B.n237 B.n236 163.367
R609 B.n237 B.n170 163.367
R610 B.n241 B.n170 163.367
R611 B.n242 B.n241 163.367
R612 B.n243 B.n242 163.367
R613 B.n243 B.n168 163.367
R614 B.n247 B.n168 163.367
R615 B.n248 B.n247 163.367
R616 B.n249 B.n248 163.367
R617 B.n249 B.n166 163.367
R618 B.n253 B.n166 163.367
R619 B.n254 B.n253 163.367
R620 B.n255 B.n254 163.367
R621 B.n255 B.n164 163.367
R622 B.n259 B.n164 163.367
R623 B.n260 B.n259 163.367
R624 B.n261 B.n260 163.367
R625 B.n261 B.n162 163.367
R626 B.n265 B.n162 163.367
R627 B.n266 B.n265 163.367
R628 B.n267 B.n266 163.367
R629 B.n267 B.n160 163.367
R630 B.n271 B.n160 163.367
R631 B.n272 B.n271 163.367
R632 B.n273 B.n272 163.367
R633 B.n273 B.n158 163.367
R634 B.n277 B.n158 163.367
R635 B.n278 B.n277 163.367
R636 B.n279 B.n278 163.367
R637 B.n279 B.n156 163.367
R638 B.n283 B.n156 163.367
R639 B.n284 B.n283 163.367
R640 B.n285 B.n284 163.367
R641 B.n285 B.n154 163.367
R642 B.n289 B.n154 163.367
R643 B.n290 B.n289 163.367
R644 B.n291 B.n290 163.367
R645 B.n291 B.n152 163.367
R646 B.n295 B.n152 163.367
R647 B.n296 B.n295 163.367
R648 B.n297 B.n296 163.367
R649 B.n297 B.n150 163.367
R650 B.n301 B.n150 163.367
R651 B.n302 B.n301 163.367
R652 B.n303 B.n302 163.367
R653 B.n303 B.n148 163.367
R654 B.n307 B.n148 163.367
R655 B.n308 B.n307 163.367
R656 B.n309 B.n308 163.367
R657 B.n309 B.n144 163.367
R658 B.n314 B.n144 163.367
R659 B.n315 B.n314 163.367
R660 B.n316 B.n315 163.367
R661 B.n316 B.n142 163.367
R662 B.n320 B.n142 163.367
R663 B.n321 B.n320 163.367
R664 B.n322 B.n321 163.367
R665 B.n322 B.n140 163.367
R666 B.n326 B.n140 163.367
R667 B.n327 B.n326 163.367
R668 B.n327 B.n136 163.367
R669 B.n331 B.n136 163.367
R670 B.n332 B.n331 163.367
R671 B.n333 B.n332 163.367
R672 B.n333 B.n134 163.367
R673 B.n337 B.n134 163.367
R674 B.n338 B.n337 163.367
R675 B.n339 B.n338 163.367
R676 B.n339 B.n132 163.367
R677 B.n343 B.n132 163.367
R678 B.n344 B.n343 163.367
R679 B.n345 B.n344 163.367
R680 B.n345 B.n130 163.367
R681 B.n349 B.n130 163.367
R682 B.n350 B.n349 163.367
R683 B.n351 B.n350 163.367
R684 B.n351 B.n128 163.367
R685 B.n355 B.n128 163.367
R686 B.n356 B.n355 163.367
R687 B.n357 B.n356 163.367
R688 B.n357 B.n126 163.367
R689 B.n361 B.n126 163.367
R690 B.n362 B.n361 163.367
R691 B.n363 B.n362 163.367
R692 B.n363 B.n124 163.367
R693 B.n367 B.n124 163.367
R694 B.n368 B.n367 163.367
R695 B.n369 B.n368 163.367
R696 B.n369 B.n122 163.367
R697 B.n373 B.n122 163.367
R698 B.n374 B.n373 163.367
R699 B.n375 B.n374 163.367
R700 B.n375 B.n120 163.367
R701 B.n379 B.n120 163.367
R702 B.n380 B.n379 163.367
R703 B.n381 B.n380 163.367
R704 B.n381 B.n118 163.367
R705 B.n385 B.n118 163.367
R706 B.n386 B.n385 163.367
R707 B.n387 B.n386 163.367
R708 B.n387 B.n116 163.367
R709 B.n391 B.n116 163.367
R710 B.n392 B.n391 163.367
R711 B.n393 B.n392 163.367
R712 B.n393 B.n114 163.367
R713 B.n397 B.n114 163.367
R714 B.n398 B.n397 163.367
R715 B.n399 B.n398 163.367
R716 B.n399 B.n112 163.367
R717 B.n403 B.n112 163.367
R718 B.n404 B.n403 163.367
R719 B.n405 B.n404 163.367
R720 B.n409 B.n110 163.367
R721 B.n410 B.n409 163.367
R722 B.n411 B.n410 163.367
R723 B.n411 B.n108 163.367
R724 B.n415 B.n108 163.367
R725 B.n416 B.n415 163.367
R726 B.n417 B.n416 163.367
R727 B.n417 B.n106 163.367
R728 B.n421 B.n106 163.367
R729 B.n422 B.n421 163.367
R730 B.n423 B.n422 163.367
R731 B.n423 B.n104 163.367
R732 B.n427 B.n104 163.367
R733 B.n428 B.n427 163.367
R734 B.n429 B.n428 163.367
R735 B.n429 B.n102 163.367
R736 B.n433 B.n102 163.367
R737 B.n434 B.n433 163.367
R738 B.n435 B.n434 163.367
R739 B.n435 B.n100 163.367
R740 B.n439 B.n100 163.367
R741 B.n440 B.n439 163.367
R742 B.n441 B.n440 163.367
R743 B.n441 B.n98 163.367
R744 B.n445 B.n98 163.367
R745 B.n446 B.n445 163.367
R746 B.n447 B.n446 163.367
R747 B.n447 B.n96 163.367
R748 B.n451 B.n96 163.367
R749 B.n452 B.n451 163.367
R750 B.n453 B.n452 163.367
R751 B.n453 B.n94 163.367
R752 B.n457 B.n94 163.367
R753 B.n458 B.n457 163.367
R754 B.n459 B.n458 163.367
R755 B.n459 B.n92 163.367
R756 B.n463 B.n92 163.367
R757 B.n464 B.n463 163.367
R758 B.n465 B.n464 163.367
R759 B.n465 B.n90 163.367
R760 B.n469 B.n90 163.367
R761 B.n470 B.n469 163.367
R762 B.n471 B.n470 163.367
R763 B.n471 B.n88 163.367
R764 B.n475 B.n88 163.367
R765 B.n476 B.n475 163.367
R766 B.n477 B.n476 163.367
R767 B.n477 B.n86 163.367
R768 B.n481 B.n86 163.367
R769 B.n482 B.n481 163.367
R770 B.n483 B.n482 163.367
R771 B.n483 B.n84 163.367
R772 B.n487 B.n84 163.367
R773 B.n488 B.n487 163.367
R774 B.n489 B.n488 163.367
R775 B.n489 B.n82 163.367
R776 B.n493 B.n82 163.367
R777 B.n494 B.n493 163.367
R778 B.n495 B.n494 163.367
R779 B.n495 B.n80 163.367
R780 B.n670 B.n17 163.367
R781 B.n670 B.n669 163.367
R782 B.n669 B.n668 163.367
R783 B.n668 B.n19 163.367
R784 B.n664 B.n19 163.367
R785 B.n664 B.n663 163.367
R786 B.n663 B.n662 163.367
R787 B.n662 B.n21 163.367
R788 B.n658 B.n21 163.367
R789 B.n658 B.n657 163.367
R790 B.n657 B.n656 163.367
R791 B.n656 B.n23 163.367
R792 B.n652 B.n23 163.367
R793 B.n652 B.n651 163.367
R794 B.n651 B.n650 163.367
R795 B.n650 B.n25 163.367
R796 B.n646 B.n25 163.367
R797 B.n646 B.n645 163.367
R798 B.n645 B.n644 163.367
R799 B.n644 B.n27 163.367
R800 B.n640 B.n27 163.367
R801 B.n640 B.n639 163.367
R802 B.n639 B.n638 163.367
R803 B.n638 B.n29 163.367
R804 B.n634 B.n29 163.367
R805 B.n634 B.n633 163.367
R806 B.n633 B.n632 163.367
R807 B.n632 B.n31 163.367
R808 B.n628 B.n31 163.367
R809 B.n628 B.n627 163.367
R810 B.n627 B.n626 163.367
R811 B.n626 B.n33 163.367
R812 B.n622 B.n33 163.367
R813 B.n622 B.n621 163.367
R814 B.n621 B.n620 163.367
R815 B.n620 B.n35 163.367
R816 B.n616 B.n35 163.367
R817 B.n616 B.n615 163.367
R818 B.n615 B.n614 163.367
R819 B.n614 B.n37 163.367
R820 B.n610 B.n37 163.367
R821 B.n610 B.n609 163.367
R822 B.n609 B.n608 163.367
R823 B.n608 B.n39 163.367
R824 B.n604 B.n39 163.367
R825 B.n604 B.n603 163.367
R826 B.n603 B.n602 163.367
R827 B.n602 B.n41 163.367
R828 B.n598 B.n41 163.367
R829 B.n598 B.n597 163.367
R830 B.n597 B.n596 163.367
R831 B.n596 B.n43 163.367
R832 B.n591 B.n43 163.367
R833 B.n591 B.n590 163.367
R834 B.n590 B.n589 163.367
R835 B.n589 B.n47 163.367
R836 B.n585 B.n47 163.367
R837 B.n585 B.n584 163.367
R838 B.n584 B.n583 163.367
R839 B.n583 B.n49 163.367
R840 B.n579 B.n49 163.367
R841 B.n579 B.n578 163.367
R842 B.n578 B.n577 163.367
R843 B.n577 B.n51 163.367
R844 B.n573 B.n51 163.367
R845 B.n573 B.n572 163.367
R846 B.n572 B.n571 163.367
R847 B.n571 B.n56 163.367
R848 B.n567 B.n56 163.367
R849 B.n567 B.n566 163.367
R850 B.n566 B.n565 163.367
R851 B.n565 B.n58 163.367
R852 B.n561 B.n58 163.367
R853 B.n561 B.n560 163.367
R854 B.n560 B.n559 163.367
R855 B.n559 B.n60 163.367
R856 B.n555 B.n60 163.367
R857 B.n555 B.n554 163.367
R858 B.n554 B.n553 163.367
R859 B.n553 B.n62 163.367
R860 B.n549 B.n62 163.367
R861 B.n549 B.n548 163.367
R862 B.n548 B.n547 163.367
R863 B.n547 B.n64 163.367
R864 B.n543 B.n64 163.367
R865 B.n543 B.n542 163.367
R866 B.n542 B.n541 163.367
R867 B.n541 B.n66 163.367
R868 B.n537 B.n66 163.367
R869 B.n537 B.n536 163.367
R870 B.n536 B.n535 163.367
R871 B.n535 B.n68 163.367
R872 B.n531 B.n68 163.367
R873 B.n531 B.n530 163.367
R874 B.n530 B.n529 163.367
R875 B.n529 B.n70 163.367
R876 B.n525 B.n70 163.367
R877 B.n525 B.n524 163.367
R878 B.n524 B.n523 163.367
R879 B.n523 B.n72 163.367
R880 B.n519 B.n72 163.367
R881 B.n519 B.n518 163.367
R882 B.n518 B.n517 163.367
R883 B.n517 B.n74 163.367
R884 B.n513 B.n74 163.367
R885 B.n513 B.n512 163.367
R886 B.n512 B.n511 163.367
R887 B.n511 B.n76 163.367
R888 B.n507 B.n76 163.367
R889 B.n507 B.n506 163.367
R890 B.n506 B.n505 163.367
R891 B.n505 B.n78 163.367
R892 B.n501 B.n78 163.367
R893 B.n501 B.n500 163.367
R894 B.n500 B.n499 163.367
R895 B.n137 B.t11 141.536
R896 B.n52 B.t1 141.536
R897 B.n145 B.t8 141.517
R898 B.n44 B.t4 141.517
R899 B.n138 B.t10 112.445
R900 B.n53 B.t2 112.445
R901 B.n146 B.t7 112.425
R902 B.n45 B.t5 112.425
R903 B.n139 B.n138 59.5399
R904 B.n311 B.n146 59.5399
R905 B.n593 B.n45 59.5399
R906 B.n54 B.n53 59.5399
R907 B.n673 B.n672 34.4981
R908 B.n498 B.n497 34.4981
R909 B.n407 B.n406 34.4981
R910 B.n232 B.n173 34.4981
R911 B.n138 B.n137 29.0914
R912 B.n146 B.n145 29.0914
R913 B.n45 B.n44 29.0914
R914 B.n53 B.n52 29.0914
R915 B B.n719 18.0485
R916 B.n672 B.n671 10.6151
R917 B.n671 B.n18 10.6151
R918 B.n667 B.n18 10.6151
R919 B.n667 B.n666 10.6151
R920 B.n666 B.n665 10.6151
R921 B.n665 B.n20 10.6151
R922 B.n661 B.n20 10.6151
R923 B.n661 B.n660 10.6151
R924 B.n660 B.n659 10.6151
R925 B.n659 B.n22 10.6151
R926 B.n655 B.n22 10.6151
R927 B.n655 B.n654 10.6151
R928 B.n654 B.n653 10.6151
R929 B.n653 B.n24 10.6151
R930 B.n649 B.n24 10.6151
R931 B.n649 B.n648 10.6151
R932 B.n648 B.n647 10.6151
R933 B.n647 B.n26 10.6151
R934 B.n643 B.n26 10.6151
R935 B.n643 B.n642 10.6151
R936 B.n642 B.n641 10.6151
R937 B.n641 B.n28 10.6151
R938 B.n637 B.n28 10.6151
R939 B.n637 B.n636 10.6151
R940 B.n636 B.n635 10.6151
R941 B.n635 B.n30 10.6151
R942 B.n631 B.n30 10.6151
R943 B.n631 B.n630 10.6151
R944 B.n630 B.n629 10.6151
R945 B.n629 B.n32 10.6151
R946 B.n625 B.n32 10.6151
R947 B.n625 B.n624 10.6151
R948 B.n624 B.n623 10.6151
R949 B.n623 B.n34 10.6151
R950 B.n619 B.n34 10.6151
R951 B.n619 B.n618 10.6151
R952 B.n618 B.n617 10.6151
R953 B.n617 B.n36 10.6151
R954 B.n613 B.n36 10.6151
R955 B.n613 B.n612 10.6151
R956 B.n612 B.n611 10.6151
R957 B.n611 B.n38 10.6151
R958 B.n607 B.n38 10.6151
R959 B.n607 B.n606 10.6151
R960 B.n606 B.n605 10.6151
R961 B.n605 B.n40 10.6151
R962 B.n601 B.n40 10.6151
R963 B.n601 B.n600 10.6151
R964 B.n600 B.n599 10.6151
R965 B.n599 B.n42 10.6151
R966 B.n595 B.n42 10.6151
R967 B.n595 B.n594 10.6151
R968 B.n592 B.n46 10.6151
R969 B.n588 B.n46 10.6151
R970 B.n588 B.n587 10.6151
R971 B.n587 B.n586 10.6151
R972 B.n586 B.n48 10.6151
R973 B.n582 B.n48 10.6151
R974 B.n582 B.n581 10.6151
R975 B.n581 B.n580 10.6151
R976 B.n580 B.n50 10.6151
R977 B.n576 B.n575 10.6151
R978 B.n575 B.n574 10.6151
R979 B.n574 B.n55 10.6151
R980 B.n570 B.n55 10.6151
R981 B.n570 B.n569 10.6151
R982 B.n569 B.n568 10.6151
R983 B.n568 B.n57 10.6151
R984 B.n564 B.n57 10.6151
R985 B.n564 B.n563 10.6151
R986 B.n563 B.n562 10.6151
R987 B.n562 B.n59 10.6151
R988 B.n558 B.n59 10.6151
R989 B.n558 B.n557 10.6151
R990 B.n557 B.n556 10.6151
R991 B.n556 B.n61 10.6151
R992 B.n552 B.n61 10.6151
R993 B.n552 B.n551 10.6151
R994 B.n551 B.n550 10.6151
R995 B.n550 B.n63 10.6151
R996 B.n546 B.n63 10.6151
R997 B.n546 B.n545 10.6151
R998 B.n545 B.n544 10.6151
R999 B.n544 B.n65 10.6151
R1000 B.n540 B.n65 10.6151
R1001 B.n540 B.n539 10.6151
R1002 B.n539 B.n538 10.6151
R1003 B.n538 B.n67 10.6151
R1004 B.n534 B.n67 10.6151
R1005 B.n534 B.n533 10.6151
R1006 B.n533 B.n532 10.6151
R1007 B.n532 B.n69 10.6151
R1008 B.n528 B.n69 10.6151
R1009 B.n528 B.n527 10.6151
R1010 B.n527 B.n526 10.6151
R1011 B.n526 B.n71 10.6151
R1012 B.n522 B.n71 10.6151
R1013 B.n522 B.n521 10.6151
R1014 B.n521 B.n520 10.6151
R1015 B.n520 B.n73 10.6151
R1016 B.n516 B.n73 10.6151
R1017 B.n516 B.n515 10.6151
R1018 B.n515 B.n514 10.6151
R1019 B.n514 B.n75 10.6151
R1020 B.n510 B.n75 10.6151
R1021 B.n510 B.n509 10.6151
R1022 B.n509 B.n508 10.6151
R1023 B.n508 B.n77 10.6151
R1024 B.n504 B.n77 10.6151
R1025 B.n504 B.n503 10.6151
R1026 B.n503 B.n502 10.6151
R1027 B.n502 B.n79 10.6151
R1028 B.n498 B.n79 10.6151
R1029 B.n408 B.n407 10.6151
R1030 B.n408 B.n109 10.6151
R1031 B.n412 B.n109 10.6151
R1032 B.n413 B.n412 10.6151
R1033 B.n414 B.n413 10.6151
R1034 B.n414 B.n107 10.6151
R1035 B.n418 B.n107 10.6151
R1036 B.n419 B.n418 10.6151
R1037 B.n420 B.n419 10.6151
R1038 B.n420 B.n105 10.6151
R1039 B.n424 B.n105 10.6151
R1040 B.n425 B.n424 10.6151
R1041 B.n426 B.n425 10.6151
R1042 B.n426 B.n103 10.6151
R1043 B.n430 B.n103 10.6151
R1044 B.n431 B.n430 10.6151
R1045 B.n432 B.n431 10.6151
R1046 B.n432 B.n101 10.6151
R1047 B.n436 B.n101 10.6151
R1048 B.n437 B.n436 10.6151
R1049 B.n438 B.n437 10.6151
R1050 B.n438 B.n99 10.6151
R1051 B.n442 B.n99 10.6151
R1052 B.n443 B.n442 10.6151
R1053 B.n444 B.n443 10.6151
R1054 B.n444 B.n97 10.6151
R1055 B.n448 B.n97 10.6151
R1056 B.n449 B.n448 10.6151
R1057 B.n450 B.n449 10.6151
R1058 B.n450 B.n95 10.6151
R1059 B.n454 B.n95 10.6151
R1060 B.n455 B.n454 10.6151
R1061 B.n456 B.n455 10.6151
R1062 B.n456 B.n93 10.6151
R1063 B.n460 B.n93 10.6151
R1064 B.n461 B.n460 10.6151
R1065 B.n462 B.n461 10.6151
R1066 B.n462 B.n91 10.6151
R1067 B.n466 B.n91 10.6151
R1068 B.n467 B.n466 10.6151
R1069 B.n468 B.n467 10.6151
R1070 B.n468 B.n89 10.6151
R1071 B.n472 B.n89 10.6151
R1072 B.n473 B.n472 10.6151
R1073 B.n474 B.n473 10.6151
R1074 B.n474 B.n87 10.6151
R1075 B.n478 B.n87 10.6151
R1076 B.n479 B.n478 10.6151
R1077 B.n480 B.n479 10.6151
R1078 B.n480 B.n85 10.6151
R1079 B.n484 B.n85 10.6151
R1080 B.n485 B.n484 10.6151
R1081 B.n486 B.n485 10.6151
R1082 B.n486 B.n83 10.6151
R1083 B.n490 B.n83 10.6151
R1084 B.n491 B.n490 10.6151
R1085 B.n492 B.n491 10.6151
R1086 B.n492 B.n81 10.6151
R1087 B.n496 B.n81 10.6151
R1088 B.n497 B.n496 10.6151
R1089 B.n233 B.n232 10.6151
R1090 B.n234 B.n233 10.6151
R1091 B.n234 B.n171 10.6151
R1092 B.n238 B.n171 10.6151
R1093 B.n239 B.n238 10.6151
R1094 B.n240 B.n239 10.6151
R1095 B.n240 B.n169 10.6151
R1096 B.n244 B.n169 10.6151
R1097 B.n245 B.n244 10.6151
R1098 B.n246 B.n245 10.6151
R1099 B.n246 B.n167 10.6151
R1100 B.n250 B.n167 10.6151
R1101 B.n251 B.n250 10.6151
R1102 B.n252 B.n251 10.6151
R1103 B.n252 B.n165 10.6151
R1104 B.n256 B.n165 10.6151
R1105 B.n257 B.n256 10.6151
R1106 B.n258 B.n257 10.6151
R1107 B.n258 B.n163 10.6151
R1108 B.n262 B.n163 10.6151
R1109 B.n263 B.n262 10.6151
R1110 B.n264 B.n263 10.6151
R1111 B.n264 B.n161 10.6151
R1112 B.n268 B.n161 10.6151
R1113 B.n269 B.n268 10.6151
R1114 B.n270 B.n269 10.6151
R1115 B.n270 B.n159 10.6151
R1116 B.n274 B.n159 10.6151
R1117 B.n275 B.n274 10.6151
R1118 B.n276 B.n275 10.6151
R1119 B.n276 B.n157 10.6151
R1120 B.n280 B.n157 10.6151
R1121 B.n281 B.n280 10.6151
R1122 B.n282 B.n281 10.6151
R1123 B.n282 B.n155 10.6151
R1124 B.n286 B.n155 10.6151
R1125 B.n287 B.n286 10.6151
R1126 B.n288 B.n287 10.6151
R1127 B.n288 B.n153 10.6151
R1128 B.n292 B.n153 10.6151
R1129 B.n293 B.n292 10.6151
R1130 B.n294 B.n293 10.6151
R1131 B.n294 B.n151 10.6151
R1132 B.n298 B.n151 10.6151
R1133 B.n299 B.n298 10.6151
R1134 B.n300 B.n299 10.6151
R1135 B.n300 B.n149 10.6151
R1136 B.n304 B.n149 10.6151
R1137 B.n305 B.n304 10.6151
R1138 B.n306 B.n305 10.6151
R1139 B.n306 B.n147 10.6151
R1140 B.n310 B.n147 10.6151
R1141 B.n313 B.n312 10.6151
R1142 B.n313 B.n143 10.6151
R1143 B.n317 B.n143 10.6151
R1144 B.n318 B.n317 10.6151
R1145 B.n319 B.n318 10.6151
R1146 B.n319 B.n141 10.6151
R1147 B.n323 B.n141 10.6151
R1148 B.n324 B.n323 10.6151
R1149 B.n325 B.n324 10.6151
R1150 B.n329 B.n328 10.6151
R1151 B.n330 B.n329 10.6151
R1152 B.n330 B.n135 10.6151
R1153 B.n334 B.n135 10.6151
R1154 B.n335 B.n334 10.6151
R1155 B.n336 B.n335 10.6151
R1156 B.n336 B.n133 10.6151
R1157 B.n340 B.n133 10.6151
R1158 B.n341 B.n340 10.6151
R1159 B.n342 B.n341 10.6151
R1160 B.n342 B.n131 10.6151
R1161 B.n346 B.n131 10.6151
R1162 B.n347 B.n346 10.6151
R1163 B.n348 B.n347 10.6151
R1164 B.n348 B.n129 10.6151
R1165 B.n352 B.n129 10.6151
R1166 B.n353 B.n352 10.6151
R1167 B.n354 B.n353 10.6151
R1168 B.n354 B.n127 10.6151
R1169 B.n358 B.n127 10.6151
R1170 B.n359 B.n358 10.6151
R1171 B.n360 B.n359 10.6151
R1172 B.n360 B.n125 10.6151
R1173 B.n364 B.n125 10.6151
R1174 B.n365 B.n364 10.6151
R1175 B.n366 B.n365 10.6151
R1176 B.n366 B.n123 10.6151
R1177 B.n370 B.n123 10.6151
R1178 B.n371 B.n370 10.6151
R1179 B.n372 B.n371 10.6151
R1180 B.n372 B.n121 10.6151
R1181 B.n376 B.n121 10.6151
R1182 B.n377 B.n376 10.6151
R1183 B.n378 B.n377 10.6151
R1184 B.n378 B.n119 10.6151
R1185 B.n382 B.n119 10.6151
R1186 B.n383 B.n382 10.6151
R1187 B.n384 B.n383 10.6151
R1188 B.n384 B.n117 10.6151
R1189 B.n388 B.n117 10.6151
R1190 B.n389 B.n388 10.6151
R1191 B.n390 B.n389 10.6151
R1192 B.n390 B.n115 10.6151
R1193 B.n394 B.n115 10.6151
R1194 B.n395 B.n394 10.6151
R1195 B.n396 B.n395 10.6151
R1196 B.n396 B.n113 10.6151
R1197 B.n400 B.n113 10.6151
R1198 B.n401 B.n400 10.6151
R1199 B.n402 B.n401 10.6151
R1200 B.n402 B.n111 10.6151
R1201 B.n406 B.n111 10.6151
R1202 B.n228 B.n173 10.6151
R1203 B.n228 B.n227 10.6151
R1204 B.n227 B.n226 10.6151
R1205 B.n226 B.n175 10.6151
R1206 B.n222 B.n175 10.6151
R1207 B.n222 B.n221 10.6151
R1208 B.n221 B.n220 10.6151
R1209 B.n220 B.n177 10.6151
R1210 B.n216 B.n177 10.6151
R1211 B.n216 B.n215 10.6151
R1212 B.n215 B.n214 10.6151
R1213 B.n214 B.n179 10.6151
R1214 B.n210 B.n179 10.6151
R1215 B.n210 B.n209 10.6151
R1216 B.n209 B.n208 10.6151
R1217 B.n208 B.n181 10.6151
R1218 B.n204 B.n181 10.6151
R1219 B.n204 B.n203 10.6151
R1220 B.n203 B.n202 10.6151
R1221 B.n202 B.n183 10.6151
R1222 B.n198 B.n183 10.6151
R1223 B.n198 B.n197 10.6151
R1224 B.n197 B.n196 10.6151
R1225 B.n196 B.n185 10.6151
R1226 B.n192 B.n185 10.6151
R1227 B.n192 B.n191 10.6151
R1228 B.n191 B.n190 10.6151
R1229 B.n190 B.n187 10.6151
R1230 B.n187 B.n0 10.6151
R1231 B.n715 B.n1 10.6151
R1232 B.n715 B.n714 10.6151
R1233 B.n714 B.n713 10.6151
R1234 B.n713 B.n4 10.6151
R1235 B.n709 B.n4 10.6151
R1236 B.n709 B.n708 10.6151
R1237 B.n708 B.n707 10.6151
R1238 B.n707 B.n6 10.6151
R1239 B.n703 B.n6 10.6151
R1240 B.n703 B.n702 10.6151
R1241 B.n702 B.n701 10.6151
R1242 B.n701 B.n8 10.6151
R1243 B.n697 B.n8 10.6151
R1244 B.n697 B.n696 10.6151
R1245 B.n696 B.n695 10.6151
R1246 B.n695 B.n10 10.6151
R1247 B.n691 B.n10 10.6151
R1248 B.n691 B.n690 10.6151
R1249 B.n690 B.n689 10.6151
R1250 B.n689 B.n12 10.6151
R1251 B.n685 B.n12 10.6151
R1252 B.n685 B.n684 10.6151
R1253 B.n684 B.n683 10.6151
R1254 B.n683 B.n14 10.6151
R1255 B.n679 B.n14 10.6151
R1256 B.n679 B.n678 10.6151
R1257 B.n678 B.n677 10.6151
R1258 B.n677 B.n16 10.6151
R1259 B.n673 B.n16 10.6151
R1260 B.n594 B.n593 9.36635
R1261 B.n576 B.n54 9.36635
R1262 B.n311 B.n310 9.36635
R1263 B.n328 B.n139 9.36635
R1264 B.n719 B.n0 2.81026
R1265 B.n719 B.n1 2.81026
R1266 B.n593 B.n592 1.24928
R1267 B.n54 B.n50 1.24928
R1268 B.n312 B.n311 1.24928
R1269 B.n325 B.n139 1.24928
C0 VTAIL w_n2470_n4158# 5.09992f
C1 VDD1 VN 0.148599f
C2 VDD2 w_n2470_n4158# 1.62739f
C3 VP B 1.46102f
C4 VTAIL VDD1 11.1998f
C5 VDD2 VDD1 1.05764f
C6 VDD1 w_n2470_n4158# 1.57282f
C7 B VN 0.938182f
C8 VP VN 6.6486f
C9 VTAIL B 5.3332f
C10 VDD2 B 1.3713f
C11 VTAIL VP 8.885321f
C12 B w_n2470_n4158# 9.033821f
C13 VDD2 VP 0.36696f
C14 VP w_n2470_n4158# 5.03448f
C15 VDD1 B 1.32008f
C16 VDD1 VP 9.316441f
C17 VTAIL VN 8.87122f
C18 VDD2 VN 9.09875f
C19 w_n2470_n4158# VN 4.71804f
C20 VTAIL VDD2 11.2447f
C21 VDD2 VSUBS 1.507236f
C22 VDD1 VSUBS 1.898173f
C23 VTAIL VSUBS 1.230684f
C24 VN VSUBS 5.29562f
C25 VP VSUBS 2.25609f
C26 B VSUBS 3.74278f
C27 w_n2470_n4158# VSUBS 0.125822p
C28 B.n0 VSUBS 0.004601f
C29 B.n1 VSUBS 0.004601f
C30 B.n2 VSUBS 0.007276f
C31 B.n3 VSUBS 0.007276f
C32 B.n4 VSUBS 0.007276f
C33 B.n5 VSUBS 0.007276f
C34 B.n6 VSUBS 0.007276f
C35 B.n7 VSUBS 0.007276f
C36 B.n8 VSUBS 0.007276f
C37 B.n9 VSUBS 0.007276f
C38 B.n10 VSUBS 0.007276f
C39 B.n11 VSUBS 0.007276f
C40 B.n12 VSUBS 0.007276f
C41 B.n13 VSUBS 0.007276f
C42 B.n14 VSUBS 0.007276f
C43 B.n15 VSUBS 0.007276f
C44 B.n16 VSUBS 0.007276f
C45 B.n17 VSUBS 0.018142f
C46 B.n18 VSUBS 0.007276f
C47 B.n19 VSUBS 0.007276f
C48 B.n20 VSUBS 0.007276f
C49 B.n21 VSUBS 0.007276f
C50 B.n22 VSUBS 0.007276f
C51 B.n23 VSUBS 0.007276f
C52 B.n24 VSUBS 0.007276f
C53 B.n25 VSUBS 0.007276f
C54 B.n26 VSUBS 0.007276f
C55 B.n27 VSUBS 0.007276f
C56 B.n28 VSUBS 0.007276f
C57 B.n29 VSUBS 0.007276f
C58 B.n30 VSUBS 0.007276f
C59 B.n31 VSUBS 0.007276f
C60 B.n32 VSUBS 0.007276f
C61 B.n33 VSUBS 0.007276f
C62 B.n34 VSUBS 0.007276f
C63 B.n35 VSUBS 0.007276f
C64 B.n36 VSUBS 0.007276f
C65 B.n37 VSUBS 0.007276f
C66 B.n38 VSUBS 0.007276f
C67 B.n39 VSUBS 0.007276f
C68 B.n40 VSUBS 0.007276f
C69 B.n41 VSUBS 0.007276f
C70 B.n42 VSUBS 0.007276f
C71 B.n43 VSUBS 0.007276f
C72 B.t5 VSUBS 0.55472f
C73 B.t4 VSUBS 0.566707f
C74 B.t3 VSUBS 0.815944f
C75 B.n44 VSUBS 0.223051f
C76 B.n45 VSUBS 0.068691f
C77 B.n46 VSUBS 0.007276f
C78 B.n47 VSUBS 0.007276f
C79 B.n48 VSUBS 0.007276f
C80 B.n49 VSUBS 0.007276f
C81 B.n50 VSUBS 0.004066f
C82 B.n51 VSUBS 0.007276f
C83 B.t2 VSUBS 0.554704f
C84 B.t1 VSUBS 0.566693f
C85 B.t0 VSUBS 0.815944f
C86 B.n52 VSUBS 0.223066f
C87 B.n53 VSUBS 0.068707f
C88 B.n54 VSUBS 0.016858f
C89 B.n55 VSUBS 0.007276f
C90 B.n56 VSUBS 0.007276f
C91 B.n57 VSUBS 0.007276f
C92 B.n58 VSUBS 0.007276f
C93 B.n59 VSUBS 0.007276f
C94 B.n60 VSUBS 0.007276f
C95 B.n61 VSUBS 0.007276f
C96 B.n62 VSUBS 0.007276f
C97 B.n63 VSUBS 0.007276f
C98 B.n64 VSUBS 0.007276f
C99 B.n65 VSUBS 0.007276f
C100 B.n66 VSUBS 0.007276f
C101 B.n67 VSUBS 0.007276f
C102 B.n68 VSUBS 0.007276f
C103 B.n69 VSUBS 0.007276f
C104 B.n70 VSUBS 0.007276f
C105 B.n71 VSUBS 0.007276f
C106 B.n72 VSUBS 0.007276f
C107 B.n73 VSUBS 0.007276f
C108 B.n74 VSUBS 0.007276f
C109 B.n75 VSUBS 0.007276f
C110 B.n76 VSUBS 0.007276f
C111 B.n77 VSUBS 0.007276f
C112 B.n78 VSUBS 0.007276f
C113 B.n79 VSUBS 0.007276f
C114 B.n80 VSUBS 0.017169f
C115 B.n81 VSUBS 0.007276f
C116 B.n82 VSUBS 0.007276f
C117 B.n83 VSUBS 0.007276f
C118 B.n84 VSUBS 0.007276f
C119 B.n85 VSUBS 0.007276f
C120 B.n86 VSUBS 0.007276f
C121 B.n87 VSUBS 0.007276f
C122 B.n88 VSUBS 0.007276f
C123 B.n89 VSUBS 0.007276f
C124 B.n90 VSUBS 0.007276f
C125 B.n91 VSUBS 0.007276f
C126 B.n92 VSUBS 0.007276f
C127 B.n93 VSUBS 0.007276f
C128 B.n94 VSUBS 0.007276f
C129 B.n95 VSUBS 0.007276f
C130 B.n96 VSUBS 0.007276f
C131 B.n97 VSUBS 0.007276f
C132 B.n98 VSUBS 0.007276f
C133 B.n99 VSUBS 0.007276f
C134 B.n100 VSUBS 0.007276f
C135 B.n101 VSUBS 0.007276f
C136 B.n102 VSUBS 0.007276f
C137 B.n103 VSUBS 0.007276f
C138 B.n104 VSUBS 0.007276f
C139 B.n105 VSUBS 0.007276f
C140 B.n106 VSUBS 0.007276f
C141 B.n107 VSUBS 0.007276f
C142 B.n108 VSUBS 0.007276f
C143 B.n109 VSUBS 0.007276f
C144 B.n110 VSUBS 0.017169f
C145 B.n111 VSUBS 0.007276f
C146 B.n112 VSUBS 0.007276f
C147 B.n113 VSUBS 0.007276f
C148 B.n114 VSUBS 0.007276f
C149 B.n115 VSUBS 0.007276f
C150 B.n116 VSUBS 0.007276f
C151 B.n117 VSUBS 0.007276f
C152 B.n118 VSUBS 0.007276f
C153 B.n119 VSUBS 0.007276f
C154 B.n120 VSUBS 0.007276f
C155 B.n121 VSUBS 0.007276f
C156 B.n122 VSUBS 0.007276f
C157 B.n123 VSUBS 0.007276f
C158 B.n124 VSUBS 0.007276f
C159 B.n125 VSUBS 0.007276f
C160 B.n126 VSUBS 0.007276f
C161 B.n127 VSUBS 0.007276f
C162 B.n128 VSUBS 0.007276f
C163 B.n129 VSUBS 0.007276f
C164 B.n130 VSUBS 0.007276f
C165 B.n131 VSUBS 0.007276f
C166 B.n132 VSUBS 0.007276f
C167 B.n133 VSUBS 0.007276f
C168 B.n134 VSUBS 0.007276f
C169 B.n135 VSUBS 0.007276f
C170 B.n136 VSUBS 0.007276f
C171 B.t10 VSUBS 0.554704f
C172 B.t11 VSUBS 0.566693f
C173 B.t9 VSUBS 0.815944f
C174 B.n137 VSUBS 0.223066f
C175 B.n138 VSUBS 0.068707f
C176 B.n139 VSUBS 0.016858f
C177 B.n140 VSUBS 0.007276f
C178 B.n141 VSUBS 0.007276f
C179 B.n142 VSUBS 0.007276f
C180 B.n143 VSUBS 0.007276f
C181 B.n144 VSUBS 0.007276f
C182 B.t7 VSUBS 0.55472f
C183 B.t8 VSUBS 0.566707f
C184 B.t6 VSUBS 0.815944f
C185 B.n145 VSUBS 0.223051f
C186 B.n146 VSUBS 0.068691f
C187 B.n147 VSUBS 0.007276f
C188 B.n148 VSUBS 0.007276f
C189 B.n149 VSUBS 0.007276f
C190 B.n150 VSUBS 0.007276f
C191 B.n151 VSUBS 0.007276f
C192 B.n152 VSUBS 0.007276f
C193 B.n153 VSUBS 0.007276f
C194 B.n154 VSUBS 0.007276f
C195 B.n155 VSUBS 0.007276f
C196 B.n156 VSUBS 0.007276f
C197 B.n157 VSUBS 0.007276f
C198 B.n158 VSUBS 0.007276f
C199 B.n159 VSUBS 0.007276f
C200 B.n160 VSUBS 0.007276f
C201 B.n161 VSUBS 0.007276f
C202 B.n162 VSUBS 0.007276f
C203 B.n163 VSUBS 0.007276f
C204 B.n164 VSUBS 0.007276f
C205 B.n165 VSUBS 0.007276f
C206 B.n166 VSUBS 0.007276f
C207 B.n167 VSUBS 0.007276f
C208 B.n168 VSUBS 0.007276f
C209 B.n169 VSUBS 0.007276f
C210 B.n170 VSUBS 0.007276f
C211 B.n171 VSUBS 0.007276f
C212 B.n172 VSUBS 0.007276f
C213 B.n173 VSUBS 0.017169f
C214 B.n174 VSUBS 0.007276f
C215 B.n175 VSUBS 0.007276f
C216 B.n176 VSUBS 0.007276f
C217 B.n177 VSUBS 0.007276f
C218 B.n178 VSUBS 0.007276f
C219 B.n179 VSUBS 0.007276f
C220 B.n180 VSUBS 0.007276f
C221 B.n181 VSUBS 0.007276f
C222 B.n182 VSUBS 0.007276f
C223 B.n183 VSUBS 0.007276f
C224 B.n184 VSUBS 0.007276f
C225 B.n185 VSUBS 0.007276f
C226 B.n186 VSUBS 0.007276f
C227 B.n187 VSUBS 0.007276f
C228 B.n188 VSUBS 0.007276f
C229 B.n189 VSUBS 0.007276f
C230 B.n190 VSUBS 0.007276f
C231 B.n191 VSUBS 0.007276f
C232 B.n192 VSUBS 0.007276f
C233 B.n193 VSUBS 0.007276f
C234 B.n194 VSUBS 0.007276f
C235 B.n195 VSUBS 0.007276f
C236 B.n196 VSUBS 0.007276f
C237 B.n197 VSUBS 0.007276f
C238 B.n198 VSUBS 0.007276f
C239 B.n199 VSUBS 0.007276f
C240 B.n200 VSUBS 0.007276f
C241 B.n201 VSUBS 0.007276f
C242 B.n202 VSUBS 0.007276f
C243 B.n203 VSUBS 0.007276f
C244 B.n204 VSUBS 0.007276f
C245 B.n205 VSUBS 0.007276f
C246 B.n206 VSUBS 0.007276f
C247 B.n207 VSUBS 0.007276f
C248 B.n208 VSUBS 0.007276f
C249 B.n209 VSUBS 0.007276f
C250 B.n210 VSUBS 0.007276f
C251 B.n211 VSUBS 0.007276f
C252 B.n212 VSUBS 0.007276f
C253 B.n213 VSUBS 0.007276f
C254 B.n214 VSUBS 0.007276f
C255 B.n215 VSUBS 0.007276f
C256 B.n216 VSUBS 0.007276f
C257 B.n217 VSUBS 0.007276f
C258 B.n218 VSUBS 0.007276f
C259 B.n219 VSUBS 0.007276f
C260 B.n220 VSUBS 0.007276f
C261 B.n221 VSUBS 0.007276f
C262 B.n222 VSUBS 0.007276f
C263 B.n223 VSUBS 0.007276f
C264 B.n224 VSUBS 0.007276f
C265 B.n225 VSUBS 0.007276f
C266 B.n226 VSUBS 0.007276f
C267 B.n227 VSUBS 0.007276f
C268 B.n228 VSUBS 0.007276f
C269 B.n229 VSUBS 0.007276f
C270 B.n230 VSUBS 0.017169f
C271 B.n231 VSUBS 0.018142f
C272 B.n232 VSUBS 0.018142f
C273 B.n233 VSUBS 0.007276f
C274 B.n234 VSUBS 0.007276f
C275 B.n235 VSUBS 0.007276f
C276 B.n236 VSUBS 0.007276f
C277 B.n237 VSUBS 0.007276f
C278 B.n238 VSUBS 0.007276f
C279 B.n239 VSUBS 0.007276f
C280 B.n240 VSUBS 0.007276f
C281 B.n241 VSUBS 0.007276f
C282 B.n242 VSUBS 0.007276f
C283 B.n243 VSUBS 0.007276f
C284 B.n244 VSUBS 0.007276f
C285 B.n245 VSUBS 0.007276f
C286 B.n246 VSUBS 0.007276f
C287 B.n247 VSUBS 0.007276f
C288 B.n248 VSUBS 0.007276f
C289 B.n249 VSUBS 0.007276f
C290 B.n250 VSUBS 0.007276f
C291 B.n251 VSUBS 0.007276f
C292 B.n252 VSUBS 0.007276f
C293 B.n253 VSUBS 0.007276f
C294 B.n254 VSUBS 0.007276f
C295 B.n255 VSUBS 0.007276f
C296 B.n256 VSUBS 0.007276f
C297 B.n257 VSUBS 0.007276f
C298 B.n258 VSUBS 0.007276f
C299 B.n259 VSUBS 0.007276f
C300 B.n260 VSUBS 0.007276f
C301 B.n261 VSUBS 0.007276f
C302 B.n262 VSUBS 0.007276f
C303 B.n263 VSUBS 0.007276f
C304 B.n264 VSUBS 0.007276f
C305 B.n265 VSUBS 0.007276f
C306 B.n266 VSUBS 0.007276f
C307 B.n267 VSUBS 0.007276f
C308 B.n268 VSUBS 0.007276f
C309 B.n269 VSUBS 0.007276f
C310 B.n270 VSUBS 0.007276f
C311 B.n271 VSUBS 0.007276f
C312 B.n272 VSUBS 0.007276f
C313 B.n273 VSUBS 0.007276f
C314 B.n274 VSUBS 0.007276f
C315 B.n275 VSUBS 0.007276f
C316 B.n276 VSUBS 0.007276f
C317 B.n277 VSUBS 0.007276f
C318 B.n278 VSUBS 0.007276f
C319 B.n279 VSUBS 0.007276f
C320 B.n280 VSUBS 0.007276f
C321 B.n281 VSUBS 0.007276f
C322 B.n282 VSUBS 0.007276f
C323 B.n283 VSUBS 0.007276f
C324 B.n284 VSUBS 0.007276f
C325 B.n285 VSUBS 0.007276f
C326 B.n286 VSUBS 0.007276f
C327 B.n287 VSUBS 0.007276f
C328 B.n288 VSUBS 0.007276f
C329 B.n289 VSUBS 0.007276f
C330 B.n290 VSUBS 0.007276f
C331 B.n291 VSUBS 0.007276f
C332 B.n292 VSUBS 0.007276f
C333 B.n293 VSUBS 0.007276f
C334 B.n294 VSUBS 0.007276f
C335 B.n295 VSUBS 0.007276f
C336 B.n296 VSUBS 0.007276f
C337 B.n297 VSUBS 0.007276f
C338 B.n298 VSUBS 0.007276f
C339 B.n299 VSUBS 0.007276f
C340 B.n300 VSUBS 0.007276f
C341 B.n301 VSUBS 0.007276f
C342 B.n302 VSUBS 0.007276f
C343 B.n303 VSUBS 0.007276f
C344 B.n304 VSUBS 0.007276f
C345 B.n305 VSUBS 0.007276f
C346 B.n306 VSUBS 0.007276f
C347 B.n307 VSUBS 0.007276f
C348 B.n308 VSUBS 0.007276f
C349 B.n309 VSUBS 0.007276f
C350 B.n310 VSUBS 0.006848f
C351 B.n311 VSUBS 0.016858f
C352 B.n312 VSUBS 0.004066f
C353 B.n313 VSUBS 0.007276f
C354 B.n314 VSUBS 0.007276f
C355 B.n315 VSUBS 0.007276f
C356 B.n316 VSUBS 0.007276f
C357 B.n317 VSUBS 0.007276f
C358 B.n318 VSUBS 0.007276f
C359 B.n319 VSUBS 0.007276f
C360 B.n320 VSUBS 0.007276f
C361 B.n321 VSUBS 0.007276f
C362 B.n322 VSUBS 0.007276f
C363 B.n323 VSUBS 0.007276f
C364 B.n324 VSUBS 0.007276f
C365 B.n325 VSUBS 0.004066f
C366 B.n326 VSUBS 0.007276f
C367 B.n327 VSUBS 0.007276f
C368 B.n328 VSUBS 0.006848f
C369 B.n329 VSUBS 0.007276f
C370 B.n330 VSUBS 0.007276f
C371 B.n331 VSUBS 0.007276f
C372 B.n332 VSUBS 0.007276f
C373 B.n333 VSUBS 0.007276f
C374 B.n334 VSUBS 0.007276f
C375 B.n335 VSUBS 0.007276f
C376 B.n336 VSUBS 0.007276f
C377 B.n337 VSUBS 0.007276f
C378 B.n338 VSUBS 0.007276f
C379 B.n339 VSUBS 0.007276f
C380 B.n340 VSUBS 0.007276f
C381 B.n341 VSUBS 0.007276f
C382 B.n342 VSUBS 0.007276f
C383 B.n343 VSUBS 0.007276f
C384 B.n344 VSUBS 0.007276f
C385 B.n345 VSUBS 0.007276f
C386 B.n346 VSUBS 0.007276f
C387 B.n347 VSUBS 0.007276f
C388 B.n348 VSUBS 0.007276f
C389 B.n349 VSUBS 0.007276f
C390 B.n350 VSUBS 0.007276f
C391 B.n351 VSUBS 0.007276f
C392 B.n352 VSUBS 0.007276f
C393 B.n353 VSUBS 0.007276f
C394 B.n354 VSUBS 0.007276f
C395 B.n355 VSUBS 0.007276f
C396 B.n356 VSUBS 0.007276f
C397 B.n357 VSUBS 0.007276f
C398 B.n358 VSUBS 0.007276f
C399 B.n359 VSUBS 0.007276f
C400 B.n360 VSUBS 0.007276f
C401 B.n361 VSUBS 0.007276f
C402 B.n362 VSUBS 0.007276f
C403 B.n363 VSUBS 0.007276f
C404 B.n364 VSUBS 0.007276f
C405 B.n365 VSUBS 0.007276f
C406 B.n366 VSUBS 0.007276f
C407 B.n367 VSUBS 0.007276f
C408 B.n368 VSUBS 0.007276f
C409 B.n369 VSUBS 0.007276f
C410 B.n370 VSUBS 0.007276f
C411 B.n371 VSUBS 0.007276f
C412 B.n372 VSUBS 0.007276f
C413 B.n373 VSUBS 0.007276f
C414 B.n374 VSUBS 0.007276f
C415 B.n375 VSUBS 0.007276f
C416 B.n376 VSUBS 0.007276f
C417 B.n377 VSUBS 0.007276f
C418 B.n378 VSUBS 0.007276f
C419 B.n379 VSUBS 0.007276f
C420 B.n380 VSUBS 0.007276f
C421 B.n381 VSUBS 0.007276f
C422 B.n382 VSUBS 0.007276f
C423 B.n383 VSUBS 0.007276f
C424 B.n384 VSUBS 0.007276f
C425 B.n385 VSUBS 0.007276f
C426 B.n386 VSUBS 0.007276f
C427 B.n387 VSUBS 0.007276f
C428 B.n388 VSUBS 0.007276f
C429 B.n389 VSUBS 0.007276f
C430 B.n390 VSUBS 0.007276f
C431 B.n391 VSUBS 0.007276f
C432 B.n392 VSUBS 0.007276f
C433 B.n393 VSUBS 0.007276f
C434 B.n394 VSUBS 0.007276f
C435 B.n395 VSUBS 0.007276f
C436 B.n396 VSUBS 0.007276f
C437 B.n397 VSUBS 0.007276f
C438 B.n398 VSUBS 0.007276f
C439 B.n399 VSUBS 0.007276f
C440 B.n400 VSUBS 0.007276f
C441 B.n401 VSUBS 0.007276f
C442 B.n402 VSUBS 0.007276f
C443 B.n403 VSUBS 0.007276f
C444 B.n404 VSUBS 0.007276f
C445 B.n405 VSUBS 0.018142f
C446 B.n406 VSUBS 0.018142f
C447 B.n407 VSUBS 0.017169f
C448 B.n408 VSUBS 0.007276f
C449 B.n409 VSUBS 0.007276f
C450 B.n410 VSUBS 0.007276f
C451 B.n411 VSUBS 0.007276f
C452 B.n412 VSUBS 0.007276f
C453 B.n413 VSUBS 0.007276f
C454 B.n414 VSUBS 0.007276f
C455 B.n415 VSUBS 0.007276f
C456 B.n416 VSUBS 0.007276f
C457 B.n417 VSUBS 0.007276f
C458 B.n418 VSUBS 0.007276f
C459 B.n419 VSUBS 0.007276f
C460 B.n420 VSUBS 0.007276f
C461 B.n421 VSUBS 0.007276f
C462 B.n422 VSUBS 0.007276f
C463 B.n423 VSUBS 0.007276f
C464 B.n424 VSUBS 0.007276f
C465 B.n425 VSUBS 0.007276f
C466 B.n426 VSUBS 0.007276f
C467 B.n427 VSUBS 0.007276f
C468 B.n428 VSUBS 0.007276f
C469 B.n429 VSUBS 0.007276f
C470 B.n430 VSUBS 0.007276f
C471 B.n431 VSUBS 0.007276f
C472 B.n432 VSUBS 0.007276f
C473 B.n433 VSUBS 0.007276f
C474 B.n434 VSUBS 0.007276f
C475 B.n435 VSUBS 0.007276f
C476 B.n436 VSUBS 0.007276f
C477 B.n437 VSUBS 0.007276f
C478 B.n438 VSUBS 0.007276f
C479 B.n439 VSUBS 0.007276f
C480 B.n440 VSUBS 0.007276f
C481 B.n441 VSUBS 0.007276f
C482 B.n442 VSUBS 0.007276f
C483 B.n443 VSUBS 0.007276f
C484 B.n444 VSUBS 0.007276f
C485 B.n445 VSUBS 0.007276f
C486 B.n446 VSUBS 0.007276f
C487 B.n447 VSUBS 0.007276f
C488 B.n448 VSUBS 0.007276f
C489 B.n449 VSUBS 0.007276f
C490 B.n450 VSUBS 0.007276f
C491 B.n451 VSUBS 0.007276f
C492 B.n452 VSUBS 0.007276f
C493 B.n453 VSUBS 0.007276f
C494 B.n454 VSUBS 0.007276f
C495 B.n455 VSUBS 0.007276f
C496 B.n456 VSUBS 0.007276f
C497 B.n457 VSUBS 0.007276f
C498 B.n458 VSUBS 0.007276f
C499 B.n459 VSUBS 0.007276f
C500 B.n460 VSUBS 0.007276f
C501 B.n461 VSUBS 0.007276f
C502 B.n462 VSUBS 0.007276f
C503 B.n463 VSUBS 0.007276f
C504 B.n464 VSUBS 0.007276f
C505 B.n465 VSUBS 0.007276f
C506 B.n466 VSUBS 0.007276f
C507 B.n467 VSUBS 0.007276f
C508 B.n468 VSUBS 0.007276f
C509 B.n469 VSUBS 0.007276f
C510 B.n470 VSUBS 0.007276f
C511 B.n471 VSUBS 0.007276f
C512 B.n472 VSUBS 0.007276f
C513 B.n473 VSUBS 0.007276f
C514 B.n474 VSUBS 0.007276f
C515 B.n475 VSUBS 0.007276f
C516 B.n476 VSUBS 0.007276f
C517 B.n477 VSUBS 0.007276f
C518 B.n478 VSUBS 0.007276f
C519 B.n479 VSUBS 0.007276f
C520 B.n480 VSUBS 0.007276f
C521 B.n481 VSUBS 0.007276f
C522 B.n482 VSUBS 0.007276f
C523 B.n483 VSUBS 0.007276f
C524 B.n484 VSUBS 0.007276f
C525 B.n485 VSUBS 0.007276f
C526 B.n486 VSUBS 0.007276f
C527 B.n487 VSUBS 0.007276f
C528 B.n488 VSUBS 0.007276f
C529 B.n489 VSUBS 0.007276f
C530 B.n490 VSUBS 0.007276f
C531 B.n491 VSUBS 0.007276f
C532 B.n492 VSUBS 0.007276f
C533 B.n493 VSUBS 0.007276f
C534 B.n494 VSUBS 0.007276f
C535 B.n495 VSUBS 0.007276f
C536 B.n496 VSUBS 0.007276f
C537 B.n497 VSUBS 0.017983f
C538 B.n498 VSUBS 0.017328f
C539 B.n499 VSUBS 0.018142f
C540 B.n500 VSUBS 0.007276f
C541 B.n501 VSUBS 0.007276f
C542 B.n502 VSUBS 0.007276f
C543 B.n503 VSUBS 0.007276f
C544 B.n504 VSUBS 0.007276f
C545 B.n505 VSUBS 0.007276f
C546 B.n506 VSUBS 0.007276f
C547 B.n507 VSUBS 0.007276f
C548 B.n508 VSUBS 0.007276f
C549 B.n509 VSUBS 0.007276f
C550 B.n510 VSUBS 0.007276f
C551 B.n511 VSUBS 0.007276f
C552 B.n512 VSUBS 0.007276f
C553 B.n513 VSUBS 0.007276f
C554 B.n514 VSUBS 0.007276f
C555 B.n515 VSUBS 0.007276f
C556 B.n516 VSUBS 0.007276f
C557 B.n517 VSUBS 0.007276f
C558 B.n518 VSUBS 0.007276f
C559 B.n519 VSUBS 0.007276f
C560 B.n520 VSUBS 0.007276f
C561 B.n521 VSUBS 0.007276f
C562 B.n522 VSUBS 0.007276f
C563 B.n523 VSUBS 0.007276f
C564 B.n524 VSUBS 0.007276f
C565 B.n525 VSUBS 0.007276f
C566 B.n526 VSUBS 0.007276f
C567 B.n527 VSUBS 0.007276f
C568 B.n528 VSUBS 0.007276f
C569 B.n529 VSUBS 0.007276f
C570 B.n530 VSUBS 0.007276f
C571 B.n531 VSUBS 0.007276f
C572 B.n532 VSUBS 0.007276f
C573 B.n533 VSUBS 0.007276f
C574 B.n534 VSUBS 0.007276f
C575 B.n535 VSUBS 0.007276f
C576 B.n536 VSUBS 0.007276f
C577 B.n537 VSUBS 0.007276f
C578 B.n538 VSUBS 0.007276f
C579 B.n539 VSUBS 0.007276f
C580 B.n540 VSUBS 0.007276f
C581 B.n541 VSUBS 0.007276f
C582 B.n542 VSUBS 0.007276f
C583 B.n543 VSUBS 0.007276f
C584 B.n544 VSUBS 0.007276f
C585 B.n545 VSUBS 0.007276f
C586 B.n546 VSUBS 0.007276f
C587 B.n547 VSUBS 0.007276f
C588 B.n548 VSUBS 0.007276f
C589 B.n549 VSUBS 0.007276f
C590 B.n550 VSUBS 0.007276f
C591 B.n551 VSUBS 0.007276f
C592 B.n552 VSUBS 0.007276f
C593 B.n553 VSUBS 0.007276f
C594 B.n554 VSUBS 0.007276f
C595 B.n555 VSUBS 0.007276f
C596 B.n556 VSUBS 0.007276f
C597 B.n557 VSUBS 0.007276f
C598 B.n558 VSUBS 0.007276f
C599 B.n559 VSUBS 0.007276f
C600 B.n560 VSUBS 0.007276f
C601 B.n561 VSUBS 0.007276f
C602 B.n562 VSUBS 0.007276f
C603 B.n563 VSUBS 0.007276f
C604 B.n564 VSUBS 0.007276f
C605 B.n565 VSUBS 0.007276f
C606 B.n566 VSUBS 0.007276f
C607 B.n567 VSUBS 0.007276f
C608 B.n568 VSUBS 0.007276f
C609 B.n569 VSUBS 0.007276f
C610 B.n570 VSUBS 0.007276f
C611 B.n571 VSUBS 0.007276f
C612 B.n572 VSUBS 0.007276f
C613 B.n573 VSUBS 0.007276f
C614 B.n574 VSUBS 0.007276f
C615 B.n575 VSUBS 0.007276f
C616 B.n576 VSUBS 0.006848f
C617 B.n577 VSUBS 0.007276f
C618 B.n578 VSUBS 0.007276f
C619 B.n579 VSUBS 0.007276f
C620 B.n580 VSUBS 0.007276f
C621 B.n581 VSUBS 0.007276f
C622 B.n582 VSUBS 0.007276f
C623 B.n583 VSUBS 0.007276f
C624 B.n584 VSUBS 0.007276f
C625 B.n585 VSUBS 0.007276f
C626 B.n586 VSUBS 0.007276f
C627 B.n587 VSUBS 0.007276f
C628 B.n588 VSUBS 0.007276f
C629 B.n589 VSUBS 0.007276f
C630 B.n590 VSUBS 0.007276f
C631 B.n591 VSUBS 0.007276f
C632 B.n592 VSUBS 0.004066f
C633 B.n593 VSUBS 0.016858f
C634 B.n594 VSUBS 0.006848f
C635 B.n595 VSUBS 0.007276f
C636 B.n596 VSUBS 0.007276f
C637 B.n597 VSUBS 0.007276f
C638 B.n598 VSUBS 0.007276f
C639 B.n599 VSUBS 0.007276f
C640 B.n600 VSUBS 0.007276f
C641 B.n601 VSUBS 0.007276f
C642 B.n602 VSUBS 0.007276f
C643 B.n603 VSUBS 0.007276f
C644 B.n604 VSUBS 0.007276f
C645 B.n605 VSUBS 0.007276f
C646 B.n606 VSUBS 0.007276f
C647 B.n607 VSUBS 0.007276f
C648 B.n608 VSUBS 0.007276f
C649 B.n609 VSUBS 0.007276f
C650 B.n610 VSUBS 0.007276f
C651 B.n611 VSUBS 0.007276f
C652 B.n612 VSUBS 0.007276f
C653 B.n613 VSUBS 0.007276f
C654 B.n614 VSUBS 0.007276f
C655 B.n615 VSUBS 0.007276f
C656 B.n616 VSUBS 0.007276f
C657 B.n617 VSUBS 0.007276f
C658 B.n618 VSUBS 0.007276f
C659 B.n619 VSUBS 0.007276f
C660 B.n620 VSUBS 0.007276f
C661 B.n621 VSUBS 0.007276f
C662 B.n622 VSUBS 0.007276f
C663 B.n623 VSUBS 0.007276f
C664 B.n624 VSUBS 0.007276f
C665 B.n625 VSUBS 0.007276f
C666 B.n626 VSUBS 0.007276f
C667 B.n627 VSUBS 0.007276f
C668 B.n628 VSUBS 0.007276f
C669 B.n629 VSUBS 0.007276f
C670 B.n630 VSUBS 0.007276f
C671 B.n631 VSUBS 0.007276f
C672 B.n632 VSUBS 0.007276f
C673 B.n633 VSUBS 0.007276f
C674 B.n634 VSUBS 0.007276f
C675 B.n635 VSUBS 0.007276f
C676 B.n636 VSUBS 0.007276f
C677 B.n637 VSUBS 0.007276f
C678 B.n638 VSUBS 0.007276f
C679 B.n639 VSUBS 0.007276f
C680 B.n640 VSUBS 0.007276f
C681 B.n641 VSUBS 0.007276f
C682 B.n642 VSUBS 0.007276f
C683 B.n643 VSUBS 0.007276f
C684 B.n644 VSUBS 0.007276f
C685 B.n645 VSUBS 0.007276f
C686 B.n646 VSUBS 0.007276f
C687 B.n647 VSUBS 0.007276f
C688 B.n648 VSUBS 0.007276f
C689 B.n649 VSUBS 0.007276f
C690 B.n650 VSUBS 0.007276f
C691 B.n651 VSUBS 0.007276f
C692 B.n652 VSUBS 0.007276f
C693 B.n653 VSUBS 0.007276f
C694 B.n654 VSUBS 0.007276f
C695 B.n655 VSUBS 0.007276f
C696 B.n656 VSUBS 0.007276f
C697 B.n657 VSUBS 0.007276f
C698 B.n658 VSUBS 0.007276f
C699 B.n659 VSUBS 0.007276f
C700 B.n660 VSUBS 0.007276f
C701 B.n661 VSUBS 0.007276f
C702 B.n662 VSUBS 0.007276f
C703 B.n663 VSUBS 0.007276f
C704 B.n664 VSUBS 0.007276f
C705 B.n665 VSUBS 0.007276f
C706 B.n666 VSUBS 0.007276f
C707 B.n667 VSUBS 0.007276f
C708 B.n668 VSUBS 0.007276f
C709 B.n669 VSUBS 0.007276f
C710 B.n670 VSUBS 0.007276f
C711 B.n671 VSUBS 0.007276f
C712 B.n672 VSUBS 0.018142f
C713 B.n673 VSUBS 0.017169f
C714 B.n674 VSUBS 0.017169f
C715 B.n675 VSUBS 0.007276f
C716 B.n676 VSUBS 0.007276f
C717 B.n677 VSUBS 0.007276f
C718 B.n678 VSUBS 0.007276f
C719 B.n679 VSUBS 0.007276f
C720 B.n680 VSUBS 0.007276f
C721 B.n681 VSUBS 0.007276f
C722 B.n682 VSUBS 0.007276f
C723 B.n683 VSUBS 0.007276f
C724 B.n684 VSUBS 0.007276f
C725 B.n685 VSUBS 0.007276f
C726 B.n686 VSUBS 0.007276f
C727 B.n687 VSUBS 0.007276f
C728 B.n688 VSUBS 0.007276f
C729 B.n689 VSUBS 0.007276f
C730 B.n690 VSUBS 0.007276f
C731 B.n691 VSUBS 0.007276f
C732 B.n692 VSUBS 0.007276f
C733 B.n693 VSUBS 0.007276f
C734 B.n694 VSUBS 0.007276f
C735 B.n695 VSUBS 0.007276f
C736 B.n696 VSUBS 0.007276f
C737 B.n697 VSUBS 0.007276f
C738 B.n698 VSUBS 0.007276f
C739 B.n699 VSUBS 0.007276f
C740 B.n700 VSUBS 0.007276f
C741 B.n701 VSUBS 0.007276f
C742 B.n702 VSUBS 0.007276f
C743 B.n703 VSUBS 0.007276f
C744 B.n704 VSUBS 0.007276f
C745 B.n705 VSUBS 0.007276f
C746 B.n706 VSUBS 0.007276f
C747 B.n707 VSUBS 0.007276f
C748 B.n708 VSUBS 0.007276f
C749 B.n709 VSUBS 0.007276f
C750 B.n710 VSUBS 0.007276f
C751 B.n711 VSUBS 0.007276f
C752 B.n712 VSUBS 0.007276f
C753 B.n713 VSUBS 0.007276f
C754 B.n714 VSUBS 0.007276f
C755 B.n715 VSUBS 0.007276f
C756 B.n716 VSUBS 0.007276f
C757 B.n717 VSUBS 0.007276f
C758 B.n718 VSUBS 0.007276f
C759 B.n719 VSUBS 0.016476f
C760 VDD2.t2 VSUBS 0.321886f
C761 VDD2.t5 VSUBS 0.321886f
C762 VDD2.n0 VSUBS 2.65591f
C763 VDD2.t7 VSUBS 0.321886f
C764 VDD2.t0 VSUBS 0.321886f
C765 VDD2.n1 VSUBS 2.65591f
C766 VDD2.n2 VSUBS 3.2804f
C767 VDD2.t1 VSUBS 0.321886f
C768 VDD2.t3 VSUBS 0.321886f
C769 VDD2.n3 VSUBS 2.65084f
C770 VDD2.n4 VSUBS 3.08255f
C771 VDD2.t4 VSUBS 0.321886f
C772 VDD2.t6 VSUBS 0.321886f
C773 VDD2.n5 VSUBS 2.65586f
C774 VN.n0 VSUBS 0.041381f
C775 VN.t7 VSUBS 2.11891f
C776 VN.n1 VSUBS 0.063206f
C777 VN.n2 VSUBS 0.041381f
C778 VN.t2 VSUBS 2.11891f
C779 VN.n3 VSUBS 0.819857f
C780 VN.t5 VSUBS 2.19272f
C781 VN.n4 VSUBS 0.853166f
C782 VN.n5 VSUBS 0.214202f
C783 VN.n6 VSUBS 0.063206f
C784 VN.n7 VSUBS 0.033452f
C785 VN.t0 VSUBS 2.11891f
C786 VN.n8 VSUBS 0.759454f
C787 VN.n9 VSUBS 0.063206f
C788 VN.n10 VSUBS 0.041381f
C789 VN.n11 VSUBS 0.041381f
C790 VN.n12 VSUBS 0.041381f
C791 VN.n13 VSUBS 0.033452f
C792 VN.n14 VSUBS 0.063206f
C793 VN.n15 VSUBS 0.825477f
C794 VN.n16 VSUBS 0.037076f
C795 VN.n17 VSUBS 0.041381f
C796 VN.t6 VSUBS 2.11891f
C797 VN.n18 VSUBS 0.063206f
C798 VN.n19 VSUBS 0.041381f
C799 VN.t4 VSUBS 2.11891f
C800 VN.n20 VSUBS 0.759454f
C801 VN.t3 VSUBS 2.11891f
C802 VN.n21 VSUBS 0.819857f
C803 VN.t1 VSUBS 2.19272f
C804 VN.n22 VSUBS 0.853166f
C805 VN.n23 VSUBS 0.214202f
C806 VN.n24 VSUBS 0.063206f
C807 VN.n25 VSUBS 0.033452f
C808 VN.n26 VSUBS 0.063206f
C809 VN.n27 VSUBS 0.041381f
C810 VN.n28 VSUBS 0.041381f
C811 VN.n29 VSUBS 0.041381f
C812 VN.n30 VSUBS 0.033452f
C813 VN.n31 VSUBS 0.063206f
C814 VN.n32 VSUBS 0.825477f
C815 VN.n33 VSUBS 2.08387f
C816 VDD1.t3 VSUBS 0.323554f
C817 VDD1.t2 VSUBS 0.323554f
C818 VDD1.n0 VSUBS 2.67072f
C819 VDD1.t4 VSUBS 0.323554f
C820 VDD1.t7 VSUBS 0.323554f
C821 VDD1.n1 VSUBS 2.66967f
C822 VDD1.t6 VSUBS 0.323554f
C823 VDD1.t5 VSUBS 0.323554f
C824 VDD1.n2 VSUBS 2.66967f
C825 VDD1.n3 VSUBS 3.35159f
C826 VDD1.t0 VSUBS 0.323554f
C827 VDD1.t1 VSUBS 0.323554f
C828 VDD1.n4 VSUBS 2.66457f
C829 VDD1.n5 VSUBS 3.12953f
C830 VTAIL.t1 VSUBS 0.296614f
C831 VTAIL.t3 VSUBS 0.296614f
C832 VTAIL.n0 VSUBS 2.3172f
C833 VTAIL.n1 VSUBS 0.635493f
C834 VTAIL.t0 VSUBS 3.02978f
C835 VTAIL.n2 VSUBS 0.763075f
C836 VTAIL.t11 VSUBS 3.02978f
C837 VTAIL.n3 VSUBS 0.763075f
C838 VTAIL.t8 VSUBS 0.296614f
C839 VTAIL.t9 VSUBS 0.296614f
C840 VTAIL.n4 VSUBS 2.3172f
C841 VTAIL.n5 VSUBS 0.729135f
C842 VTAIL.t15 VSUBS 3.02978f
C843 VTAIL.n6 VSUBS 2.18781f
C844 VTAIL.t6 VSUBS 3.0298f
C845 VTAIL.n7 VSUBS 2.18779f
C846 VTAIL.t4 VSUBS 0.296614f
C847 VTAIL.t2 VSUBS 0.296614f
C848 VTAIL.n8 VSUBS 2.3172f
C849 VTAIL.n9 VSUBS 0.729131f
C850 VTAIL.t5 VSUBS 3.0298f
C851 VTAIL.n10 VSUBS 0.763053f
C852 VTAIL.t10 VSUBS 3.0298f
C853 VTAIL.n11 VSUBS 0.763053f
C854 VTAIL.t14 VSUBS 0.296614f
C855 VTAIL.t12 VSUBS 0.296614f
C856 VTAIL.n12 VSUBS 2.3172f
C857 VTAIL.n13 VSUBS 0.729131f
C858 VTAIL.t13 VSUBS 3.02978f
C859 VTAIL.n14 VSUBS 2.18781f
C860 VTAIL.t7 VSUBS 3.02978f
C861 VTAIL.n15 VSUBS 2.1834f
C862 VP.n0 VSUBS 0.042171f
C863 VP.t2 VSUBS 2.15935f
C864 VP.n1 VSUBS 0.064412f
C865 VP.n2 VSUBS 0.042171f
C866 VP.t0 VSUBS 2.15935f
C867 VP.n3 VSUBS 0.77395f
C868 VP.n4 VSUBS 0.042171f
C869 VP.t3 VSUBS 2.15935f
C870 VP.n5 VSUBS 0.841234f
C871 VP.n6 VSUBS 0.042171f
C872 VP.t6 VSUBS 2.15935f
C873 VP.n7 VSUBS 0.064412f
C874 VP.n8 VSUBS 0.042171f
C875 VP.t5 VSUBS 2.15935f
C876 VP.n9 VSUBS 0.835506f
C877 VP.t4 VSUBS 2.23458f
C878 VP.n10 VSUBS 0.869451f
C879 VP.n11 VSUBS 0.218291f
C880 VP.n12 VSUBS 0.064412f
C881 VP.n13 VSUBS 0.034091f
C882 VP.t7 VSUBS 2.15935f
C883 VP.n14 VSUBS 0.77395f
C884 VP.n15 VSUBS 0.064412f
C885 VP.n16 VSUBS 0.042171f
C886 VP.n17 VSUBS 0.042171f
C887 VP.n18 VSUBS 0.042171f
C888 VP.n19 VSUBS 0.034091f
C889 VP.n20 VSUBS 0.064412f
C890 VP.n21 VSUBS 0.841234f
C891 VP.n22 VSUBS 2.09615f
C892 VP.n23 VSUBS 2.12835f
C893 VP.n24 VSUBS 0.042171f
C894 VP.n25 VSUBS 0.064412f
C895 VP.n26 VSUBS 0.034091f
C896 VP.n27 VSUBS 0.064412f
C897 VP.n28 VSUBS 0.042171f
C898 VP.n29 VSUBS 0.042171f
C899 VP.n30 VSUBS 0.064412f
C900 VP.n31 VSUBS 0.034091f
C901 VP.t1 VSUBS 2.15935f
C902 VP.n32 VSUBS 0.77395f
C903 VP.n33 VSUBS 0.064412f
C904 VP.n34 VSUBS 0.042171f
C905 VP.n35 VSUBS 0.042171f
C906 VP.n36 VSUBS 0.042171f
C907 VP.n37 VSUBS 0.034091f
C908 VP.n38 VSUBS 0.064412f
C909 VP.n39 VSUBS 0.841234f
C910 VP.n40 VSUBS 0.037783f
.ends

