* NGSPICE file created from diff_pair_sample_0683.ext - technology: sky130A

.subckt diff_pair_sample_0683 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0 ps=0 w=0.61 l=0.77
X1 B.t8 B.t6 B.t7 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0 ps=0 w=0.61 l=0.77
X2 VTAIL.t7 VN.t0 VDD2.t0 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0.10065 ps=0.94 w=0.61 l=0.77
X3 VTAIL.t3 VP.t0 VDD1.t3 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0.10065 ps=0.94 w=0.61 l=0.77
X4 VDD2.t2 VN.t1 VTAIL.t6 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.10065 pd=0.94 as=0.2379 ps=2 w=0.61 l=0.77
X5 VTAIL.t2 VP.t1 VDD1.t2 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0.10065 ps=0.94 w=0.61 l=0.77
X6 VDD1.t1 VP.t2 VTAIL.t0 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.10065 pd=0.94 as=0.2379 ps=2 w=0.61 l=0.77
X7 B.t5 B.t3 B.t4 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0 ps=0 w=0.61 l=0.77
X8 VDD2.t3 VN.t2 VTAIL.t5 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.10065 pd=0.94 as=0.2379 ps=2 w=0.61 l=0.77
X9 VDD1.t0 VP.t3 VTAIL.t1 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.10065 pd=0.94 as=0.2379 ps=2 w=0.61 l=0.77
X10 B.t2 B.t0 B.t1 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0 ps=0 w=0.61 l=0.77
X11 VTAIL.t4 VN.t3 VDD2.t1 w_n1630_n1090# sky130_fd_pr__pfet_01v8 ad=0.2379 pd=2 as=0.10065 ps=0.94 w=0.61 l=0.77
R0 B.n52 B.t5 681.149
R1 B.n58 B.t8 681.149
R2 B.n16 B.t10 681.149
R3 B.n22 B.t1 681.149
R4 B.n53 B.t4 659.814
R5 B.n59 B.t7 659.814
R6 B.n17 B.t11 659.814
R7 B.n23 B.t2 659.814
R8 B.n195 B.n28 585
R9 B.n197 B.n196 585
R10 B.n198 B.n27 585
R11 B.n200 B.n199 585
R12 B.n201 B.n26 585
R13 B.n203 B.n202 585
R14 B.n204 B.n25 585
R15 B.n206 B.n205 585
R16 B.n208 B.n207 585
R17 B.n209 B.n21 585
R18 B.n211 B.n210 585
R19 B.n212 B.n20 585
R20 B.n214 B.n213 585
R21 B.n215 B.n19 585
R22 B.n217 B.n216 585
R23 B.n218 B.n18 585
R24 B.n220 B.n219 585
R25 B.n221 B.n15 585
R26 B.n224 B.n223 585
R27 B.n225 B.n14 585
R28 B.n227 B.n226 585
R29 B.n228 B.n13 585
R30 B.n230 B.n229 585
R31 B.n231 B.n12 585
R32 B.n233 B.n232 585
R33 B.n234 B.n11 585
R34 B.n194 B.n193 585
R35 B.n192 B.n29 585
R36 B.n191 B.n190 585
R37 B.n189 B.n30 585
R38 B.n188 B.n187 585
R39 B.n186 B.n31 585
R40 B.n185 B.n184 585
R41 B.n183 B.n32 585
R42 B.n182 B.n181 585
R43 B.n180 B.n33 585
R44 B.n179 B.n178 585
R45 B.n177 B.n34 585
R46 B.n176 B.n175 585
R47 B.n174 B.n35 585
R48 B.n173 B.n172 585
R49 B.n171 B.n36 585
R50 B.n170 B.n169 585
R51 B.n168 B.n37 585
R52 B.n167 B.n166 585
R53 B.n165 B.n38 585
R54 B.n164 B.n163 585
R55 B.n162 B.n39 585
R56 B.n161 B.n160 585
R57 B.n159 B.n40 585
R58 B.n158 B.n157 585
R59 B.n156 B.n41 585
R60 B.n155 B.n154 585
R61 B.n153 B.n42 585
R62 B.n152 B.n151 585
R63 B.n150 B.n43 585
R64 B.n149 B.n148 585
R65 B.n147 B.n44 585
R66 B.n146 B.n145 585
R67 B.n144 B.n45 585
R68 B.n143 B.n142 585
R69 B.n141 B.n46 585
R70 B.n140 B.n139 585
R71 B.n99 B.n64 585
R72 B.n101 B.n100 585
R73 B.n102 B.n63 585
R74 B.n104 B.n103 585
R75 B.n105 B.n62 585
R76 B.n107 B.n106 585
R77 B.n108 B.n61 585
R78 B.n110 B.n109 585
R79 B.n112 B.n111 585
R80 B.n113 B.n57 585
R81 B.n115 B.n114 585
R82 B.n116 B.n56 585
R83 B.n118 B.n117 585
R84 B.n119 B.n55 585
R85 B.n121 B.n120 585
R86 B.n122 B.n54 585
R87 B.n124 B.n123 585
R88 B.n125 B.n51 585
R89 B.n128 B.n127 585
R90 B.n129 B.n50 585
R91 B.n131 B.n130 585
R92 B.n132 B.n49 585
R93 B.n134 B.n133 585
R94 B.n135 B.n48 585
R95 B.n137 B.n136 585
R96 B.n138 B.n47 585
R97 B.n98 B.n97 585
R98 B.n96 B.n65 585
R99 B.n95 B.n94 585
R100 B.n93 B.n66 585
R101 B.n92 B.n91 585
R102 B.n90 B.n67 585
R103 B.n89 B.n88 585
R104 B.n87 B.n68 585
R105 B.n86 B.n85 585
R106 B.n84 B.n69 585
R107 B.n83 B.n82 585
R108 B.n81 B.n70 585
R109 B.n80 B.n79 585
R110 B.n78 B.n71 585
R111 B.n77 B.n76 585
R112 B.n75 B.n72 585
R113 B.n74 B.n73 585
R114 B.n2 B.n0 585
R115 B.n261 B.n1 585
R116 B.n260 B.n259 585
R117 B.n258 B.n3 585
R118 B.n257 B.n256 585
R119 B.n255 B.n4 585
R120 B.n254 B.n253 585
R121 B.n252 B.n5 585
R122 B.n251 B.n250 585
R123 B.n249 B.n6 585
R124 B.n248 B.n247 585
R125 B.n246 B.n7 585
R126 B.n245 B.n244 585
R127 B.n243 B.n8 585
R128 B.n242 B.n241 585
R129 B.n240 B.n9 585
R130 B.n239 B.n238 585
R131 B.n237 B.n10 585
R132 B.n236 B.n235 585
R133 B.n263 B.n262 585
R134 B.n99 B.n98 454.062
R135 B.n236 B.n11 454.062
R136 B.n140 B.n47 454.062
R137 B.n195 B.n194 454.062
R138 B.n52 B.t3 221.274
R139 B.n58 B.t6 221.274
R140 B.n16 B.t9 221.274
R141 B.n22 B.t0 221.274
R142 B.n98 B.n65 163.367
R143 B.n94 B.n65 163.367
R144 B.n94 B.n93 163.367
R145 B.n93 B.n92 163.367
R146 B.n92 B.n67 163.367
R147 B.n88 B.n67 163.367
R148 B.n88 B.n87 163.367
R149 B.n87 B.n86 163.367
R150 B.n86 B.n69 163.367
R151 B.n82 B.n69 163.367
R152 B.n82 B.n81 163.367
R153 B.n81 B.n80 163.367
R154 B.n80 B.n71 163.367
R155 B.n76 B.n71 163.367
R156 B.n76 B.n75 163.367
R157 B.n75 B.n74 163.367
R158 B.n74 B.n2 163.367
R159 B.n262 B.n2 163.367
R160 B.n262 B.n261 163.367
R161 B.n261 B.n260 163.367
R162 B.n260 B.n3 163.367
R163 B.n256 B.n3 163.367
R164 B.n256 B.n255 163.367
R165 B.n255 B.n254 163.367
R166 B.n254 B.n5 163.367
R167 B.n250 B.n5 163.367
R168 B.n250 B.n249 163.367
R169 B.n249 B.n248 163.367
R170 B.n248 B.n7 163.367
R171 B.n244 B.n7 163.367
R172 B.n244 B.n243 163.367
R173 B.n243 B.n242 163.367
R174 B.n242 B.n9 163.367
R175 B.n238 B.n9 163.367
R176 B.n238 B.n237 163.367
R177 B.n237 B.n236 163.367
R178 B.n100 B.n99 163.367
R179 B.n100 B.n63 163.367
R180 B.n104 B.n63 163.367
R181 B.n105 B.n104 163.367
R182 B.n106 B.n105 163.367
R183 B.n106 B.n61 163.367
R184 B.n110 B.n61 163.367
R185 B.n111 B.n110 163.367
R186 B.n111 B.n57 163.367
R187 B.n115 B.n57 163.367
R188 B.n116 B.n115 163.367
R189 B.n117 B.n116 163.367
R190 B.n117 B.n55 163.367
R191 B.n121 B.n55 163.367
R192 B.n122 B.n121 163.367
R193 B.n123 B.n122 163.367
R194 B.n123 B.n51 163.367
R195 B.n128 B.n51 163.367
R196 B.n129 B.n128 163.367
R197 B.n130 B.n129 163.367
R198 B.n130 B.n49 163.367
R199 B.n134 B.n49 163.367
R200 B.n135 B.n134 163.367
R201 B.n136 B.n135 163.367
R202 B.n136 B.n47 163.367
R203 B.n141 B.n140 163.367
R204 B.n142 B.n141 163.367
R205 B.n142 B.n45 163.367
R206 B.n146 B.n45 163.367
R207 B.n147 B.n146 163.367
R208 B.n148 B.n147 163.367
R209 B.n148 B.n43 163.367
R210 B.n152 B.n43 163.367
R211 B.n153 B.n152 163.367
R212 B.n154 B.n153 163.367
R213 B.n154 B.n41 163.367
R214 B.n158 B.n41 163.367
R215 B.n159 B.n158 163.367
R216 B.n160 B.n159 163.367
R217 B.n160 B.n39 163.367
R218 B.n164 B.n39 163.367
R219 B.n165 B.n164 163.367
R220 B.n166 B.n165 163.367
R221 B.n166 B.n37 163.367
R222 B.n170 B.n37 163.367
R223 B.n171 B.n170 163.367
R224 B.n172 B.n171 163.367
R225 B.n172 B.n35 163.367
R226 B.n176 B.n35 163.367
R227 B.n177 B.n176 163.367
R228 B.n178 B.n177 163.367
R229 B.n178 B.n33 163.367
R230 B.n182 B.n33 163.367
R231 B.n183 B.n182 163.367
R232 B.n184 B.n183 163.367
R233 B.n184 B.n31 163.367
R234 B.n188 B.n31 163.367
R235 B.n189 B.n188 163.367
R236 B.n190 B.n189 163.367
R237 B.n190 B.n29 163.367
R238 B.n194 B.n29 163.367
R239 B.n232 B.n11 163.367
R240 B.n232 B.n231 163.367
R241 B.n231 B.n230 163.367
R242 B.n230 B.n13 163.367
R243 B.n226 B.n13 163.367
R244 B.n226 B.n225 163.367
R245 B.n225 B.n224 163.367
R246 B.n224 B.n15 163.367
R247 B.n219 B.n15 163.367
R248 B.n219 B.n218 163.367
R249 B.n218 B.n217 163.367
R250 B.n217 B.n19 163.367
R251 B.n213 B.n19 163.367
R252 B.n213 B.n212 163.367
R253 B.n212 B.n211 163.367
R254 B.n211 B.n21 163.367
R255 B.n207 B.n21 163.367
R256 B.n207 B.n206 163.367
R257 B.n206 B.n25 163.367
R258 B.n202 B.n25 163.367
R259 B.n202 B.n201 163.367
R260 B.n201 B.n200 163.367
R261 B.n200 B.n27 163.367
R262 B.n196 B.n27 163.367
R263 B.n196 B.n195 163.367
R264 B.n126 B.n53 59.5399
R265 B.n60 B.n59 59.5399
R266 B.n222 B.n17 59.5399
R267 B.n24 B.n23 59.5399
R268 B.n235 B.n234 29.5029
R269 B.n139 B.n138 29.5029
R270 B.n97 B.n64 29.5029
R271 B.n193 B.n28 29.5029
R272 B.n53 B.n52 21.3338
R273 B.n59 B.n58 21.3338
R274 B.n17 B.n16 21.3338
R275 B.n23 B.n22 21.3338
R276 B B.n263 18.0485
R277 B.n234 B.n233 10.6151
R278 B.n233 B.n12 10.6151
R279 B.n229 B.n12 10.6151
R280 B.n229 B.n228 10.6151
R281 B.n228 B.n227 10.6151
R282 B.n227 B.n14 10.6151
R283 B.n223 B.n14 10.6151
R284 B.n221 B.n220 10.6151
R285 B.n220 B.n18 10.6151
R286 B.n216 B.n18 10.6151
R287 B.n216 B.n215 10.6151
R288 B.n215 B.n214 10.6151
R289 B.n214 B.n20 10.6151
R290 B.n210 B.n20 10.6151
R291 B.n210 B.n209 10.6151
R292 B.n209 B.n208 10.6151
R293 B.n205 B.n204 10.6151
R294 B.n204 B.n203 10.6151
R295 B.n203 B.n26 10.6151
R296 B.n199 B.n26 10.6151
R297 B.n199 B.n198 10.6151
R298 B.n198 B.n197 10.6151
R299 B.n197 B.n28 10.6151
R300 B.n139 B.n46 10.6151
R301 B.n143 B.n46 10.6151
R302 B.n144 B.n143 10.6151
R303 B.n145 B.n144 10.6151
R304 B.n145 B.n44 10.6151
R305 B.n149 B.n44 10.6151
R306 B.n150 B.n149 10.6151
R307 B.n151 B.n150 10.6151
R308 B.n151 B.n42 10.6151
R309 B.n155 B.n42 10.6151
R310 B.n156 B.n155 10.6151
R311 B.n157 B.n156 10.6151
R312 B.n157 B.n40 10.6151
R313 B.n161 B.n40 10.6151
R314 B.n162 B.n161 10.6151
R315 B.n163 B.n162 10.6151
R316 B.n163 B.n38 10.6151
R317 B.n167 B.n38 10.6151
R318 B.n168 B.n167 10.6151
R319 B.n169 B.n168 10.6151
R320 B.n169 B.n36 10.6151
R321 B.n173 B.n36 10.6151
R322 B.n174 B.n173 10.6151
R323 B.n175 B.n174 10.6151
R324 B.n175 B.n34 10.6151
R325 B.n179 B.n34 10.6151
R326 B.n180 B.n179 10.6151
R327 B.n181 B.n180 10.6151
R328 B.n181 B.n32 10.6151
R329 B.n185 B.n32 10.6151
R330 B.n186 B.n185 10.6151
R331 B.n187 B.n186 10.6151
R332 B.n187 B.n30 10.6151
R333 B.n191 B.n30 10.6151
R334 B.n192 B.n191 10.6151
R335 B.n193 B.n192 10.6151
R336 B.n101 B.n64 10.6151
R337 B.n102 B.n101 10.6151
R338 B.n103 B.n102 10.6151
R339 B.n103 B.n62 10.6151
R340 B.n107 B.n62 10.6151
R341 B.n108 B.n107 10.6151
R342 B.n109 B.n108 10.6151
R343 B.n113 B.n112 10.6151
R344 B.n114 B.n113 10.6151
R345 B.n114 B.n56 10.6151
R346 B.n118 B.n56 10.6151
R347 B.n119 B.n118 10.6151
R348 B.n120 B.n119 10.6151
R349 B.n120 B.n54 10.6151
R350 B.n124 B.n54 10.6151
R351 B.n125 B.n124 10.6151
R352 B.n127 B.n50 10.6151
R353 B.n131 B.n50 10.6151
R354 B.n132 B.n131 10.6151
R355 B.n133 B.n132 10.6151
R356 B.n133 B.n48 10.6151
R357 B.n137 B.n48 10.6151
R358 B.n138 B.n137 10.6151
R359 B.n97 B.n96 10.6151
R360 B.n96 B.n95 10.6151
R361 B.n95 B.n66 10.6151
R362 B.n91 B.n66 10.6151
R363 B.n91 B.n90 10.6151
R364 B.n90 B.n89 10.6151
R365 B.n89 B.n68 10.6151
R366 B.n85 B.n68 10.6151
R367 B.n85 B.n84 10.6151
R368 B.n84 B.n83 10.6151
R369 B.n83 B.n70 10.6151
R370 B.n79 B.n70 10.6151
R371 B.n79 B.n78 10.6151
R372 B.n78 B.n77 10.6151
R373 B.n77 B.n72 10.6151
R374 B.n73 B.n72 10.6151
R375 B.n73 B.n0 10.6151
R376 B.n259 B.n1 10.6151
R377 B.n259 B.n258 10.6151
R378 B.n258 B.n257 10.6151
R379 B.n257 B.n4 10.6151
R380 B.n253 B.n4 10.6151
R381 B.n253 B.n252 10.6151
R382 B.n252 B.n251 10.6151
R383 B.n251 B.n6 10.6151
R384 B.n247 B.n6 10.6151
R385 B.n247 B.n246 10.6151
R386 B.n246 B.n245 10.6151
R387 B.n245 B.n8 10.6151
R388 B.n241 B.n8 10.6151
R389 B.n241 B.n240 10.6151
R390 B.n240 B.n239 10.6151
R391 B.n239 B.n10 10.6151
R392 B.n235 B.n10 10.6151
R393 B.n223 B.n222 9.36635
R394 B.n205 B.n24 9.36635
R395 B.n109 B.n60 9.36635
R396 B.n127 B.n126 9.36635
R397 B.n263 B.n0 2.81026
R398 B.n263 B.n1 2.81026
R399 B.n222 B.n221 1.24928
R400 B.n208 B.n24 1.24928
R401 B.n112 B.n60 1.24928
R402 B.n126 B.n125 1.24928
R403 VN.n0 VN.t3 91.4188
R404 VN.n1 VN.t1 91.4188
R405 VN.n0 VN.t2 91.3692
R406 VN.n1 VN.t0 91.3692
R407 VN VN.n1 77.0882
R408 VN VN.n0 44.7132
R409 VDD2.n2 VDD2.n0 661.144
R410 VDD2.n2 VDD2.n1 634.058
R411 VDD2.n1 VDD2.t0 53.2874
R412 VDD2.n1 VDD2.t2 53.2874
R413 VDD2.n0 VDD2.t1 53.2874
R414 VDD2.n0 VDD2.t3 53.2874
R415 VDD2 VDD2.n2 0.0586897
R416 VTAIL.n7 VTAIL.t5 670.667
R417 VTAIL.n0 VTAIL.t4 670.667
R418 VTAIL.n1 VTAIL.t0 670.667
R419 VTAIL.n2 VTAIL.t3 670.667
R420 VTAIL.n6 VTAIL.t1 670.667
R421 VTAIL.n5 VTAIL.t2 670.667
R422 VTAIL.n4 VTAIL.t6 670.667
R423 VTAIL.n3 VTAIL.t7 670.667
R424 VTAIL.n7 VTAIL.n6 13.841
R425 VTAIL.n3 VTAIL.n2 13.841
R426 VTAIL.n4 VTAIL.n3 0.948776
R427 VTAIL.n6 VTAIL.n5 0.948776
R428 VTAIL.n2 VTAIL.n1 0.948776
R429 VTAIL VTAIL.n0 0.532828
R430 VTAIL.n5 VTAIL.n4 0.470328
R431 VTAIL.n1 VTAIL.n0 0.470328
R432 VTAIL VTAIL.n7 0.416448
R433 VP.n6 VP.n5 161.3
R434 VP.n4 VP.n0 161.3
R435 VP.n3 VP.n2 161.3
R436 VP.n1 VP.t1 91.4188
R437 VP.n1 VP.t3 91.3692
R438 VP.n2 VP.n1 76.7075
R439 VP.n3 VP.t0 70.4226
R440 VP.n5 VP.t2 70.4226
R441 VP.n4 VP.n3 24.1005
R442 VP.n5 VP.n4 24.1005
R443 VP.n2 VP.n0 0.189894
R444 VP.n6 VP.n0 0.189894
R445 VP VP.n6 0.0516364
R446 VDD1 VDD1.n1 661.668
R447 VDD1 VDD1.n0 634.116
R448 VDD1.n0 VDD1.t2 53.2874
R449 VDD1.n0 VDD1.t0 53.2874
R450 VDD1.n1 VDD1.t3 53.2874
R451 VDD1.n1 VDD1.t1 53.2874
C0 w_n1630_n1090# B 3.78443f
C1 VDD1 VN 0.15483f
C2 VTAIL VP 0.722508f
C3 w_n1630_n1090# VN 2.144f
C4 VDD1 VP 0.582603f
C5 w_n1630_n1090# VP 2.33973f
C6 VDD2 B 0.652979f
C7 VDD2 VN 0.452402f
C8 VDD1 VTAIL 1.76201f
C9 w_n1630_n1090# VTAIL 1.13825f
C10 VDD2 VP 0.286656f
C11 VDD1 w_n1630_n1090# 0.760935f
C12 VDD2 VTAIL 1.80395f
C13 VDD1 VDD2 0.582999f
C14 VDD2 w_n1630_n1090# 0.775544f
C15 VN B 0.585049f
C16 B VP 0.91506f
C17 VN VP 2.77266f
C18 VTAIL B 0.679832f
C19 VN VTAIL 0.708401f
C20 VDD1 B 0.630084f
C21 VDD2 VSUBS 0.316139f
C22 VDD1 VSUBS 0.518386f
C23 VTAIL VSUBS 0.194962f
C24 VN VSUBS 4.460701f
C25 VP VSUBS 0.822026f
C26 B VSUBS 1.63402f
C27 w_n1630_n1090# VSUBS 23.0221f
C28 VP.n0 VSUBS 0.070936f
C29 VP.t3 VSUBS 0.163276f
C30 VP.t1 VSUBS 0.163412f
C31 VP.n1 VSUBS 1.06165f
C32 VP.n2 VSUBS 2.97073f
C33 VP.t0 VSUBS 0.12603f
C34 VP.n3 VSUBS 0.157361f
C35 VP.n4 VSUBS 0.016097f
C36 VP.t2 VSUBS 0.12603f
C37 VP.n5 VSUBS 0.157361f
C38 VP.n6 VSUBS 0.054972f
C39 VN.t3 VSUBS 0.153993f
C40 VN.t2 VSUBS 0.153865f
C41 VN.n0 VSUBS 0.242122f
C42 VN.t1 VSUBS 0.153993f
C43 VN.t0 VSUBS 0.153865f
C44 VN.n1 VSUBS 1.0245f
C45 B.n0 VSUBS 0.006947f
C46 B.n1 VSUBS 0.006947f
C47 B.n2 VSUBS 0.010986f
C48 B.n3 VSUBS 0.010986f
C49 B.n4 VSUBS 0.010986f
C50 B.n5 VSUBS 0.010986f
C51 B.n6 VSUBS 0.010986f
C52 B.n7 VSUBS 0.010986f
C53 B.n8 VSUBS 0.010986f
C54 B.n9 VSUBS 0.010986f
C55 B.n10 VSUBS 0.010986f
C56 B.n11 VSUBS 0.02465f
C57 B.n12 VSUBS 0.010986f
C58 B.n13 VSUBS 0.010986f
C59 B.n14 VSUBS 0.010986f
C60 B.n15 VSUBS 0.010986f
C61 B.t11 VSUBS 0.018048f
C62 B.t10 VSUBS 0.019129f
C63 B.t9 VSUBS 0.0405f
C64 B.n16 VSUBS 0.052827f
C65 B.n17 VSUBS 0.050176f
C66 B.n18 VSUBS 0.010986f
C67 B.n19 VSUBS 0.010986f
C68 B.n20 VSUBS 0.010986f
C69 B.n21 VSUBS 0.010986f
C70 B.t2 VSUBS 0.018048f
C71 B.t1 VSUBS 0.019129f
C72 B.t0 VSUBS 0.0405f
C73 B.n22 VSUBS 0.052827f
C74 B.n23 VSUBS 0.050176f
C75 B.n24 VSUBS 0.025452f
C76 B.n25 VSUBS 0.010986f
C77 B.n26 VSUBS 0.010986f
C78 B.n27 VSUBS 0.010986f
C79 B.n28 VSUBS 0.023213f
C80 B.n29 VSUBS 0.010986f
C81 B.n30 VSUBS 0.010986f
C82 B.n31 VSUBS 0.010986f
C83 B.n32 VSUBS 0.010986f
C84 B.n33 VSUBS 0.010986f
C85 B.n34 VSUBS 0.010986f
C86 B.n35 VSUBS 0.010986f
C87 B.n36 VSUBS 0.010986f
C88 B.n37 VSUBS 0.010986f
C89 B.n38 VSUBS 0.010986f
C90 B.n39 VSUBS 0.010986f
C91 B.n40 VSUBS 0.010986f
C92 B.n41 VSUBS 0.010986f
C93 B.n42 VSUBS 0.010986f
C94 B.n43 VSUBS 0.010986f
C95 B.n44 VSUBS 0.010986f
C96 B.n45 VSUBS 0.010986f
C97 B.n46 VSUBS 0.010986f
C98 B.n47 VSUBS 0.02465f
C99 B.n48 VSUBS 0.010986f
C100 B.n49 VSUBS 0.010986f
C101 B.n50 VSUBS 0.010986f
C102 B.n51 VSUBS 0.010986f
C103 B.t4 VSUBS 0.018048f
C104 B.t5 VSUBS 0.019129f
C105 B.t3 VSUBS 0.0405f
C106 B.n52 VSUBS 0.052827f
C107 B.n53 VSUBS 0.050176f
C108 B.n54 VSUBS 0.010986f
C109 B.n55 VSUBS 0.010986f
C110 B.n56 VSUBS 0.010986f
C111 B.n57 VSUBS 0.010986f
C112 B.t7 VSUBS 0.018048f
C113 B.t8 VSUBS 0.019129f
C114 B.t6 VSUBS 0.0405f
C115 B.n58 VSUBS 0.052827f
C116 B.n59 VSUBS 0.050176f
C117 B.n60 VSUBS 0.025452f
C118 B.n61 VSUBS 0.010986f
C119 B.n62 VSUBS 0.010986f
C120 B.n63 VSUBS 0.010986f
C121 B.n64 VSUBS 0.02465f
C122 B.n65 VSUBS 0.010986f
C123 B.n66 VSUBS 0.010986f
C124 B.n67 VSUBS 0.010986f
C125 B.n68 VSUBS 0.010986f
C126 B.n69 VSUBS 0.010986f
C127 B.n70 VSUBS 0.010986f
C128 B.n71 VSUBS 0.010986f
C129 B.n72 VSUBS 0.010986f
C130 B.n73 VSUBS 0.010986f
C131 B.n74 VSUBS 0.010986f
C132 B.n75 VSUBS 0.010986f
C133 B.n76 VSUBS 0.010986f
C134 B.n77 VSUBS 0.010986f
C135 B.n78 VSUBS 0.010986f
C136 B.n79 VSUBS 0.010986f
C137 B.n80 VSUBS 0.010986f
C138 B.n81 VSUBS 0.010986f
C139 B.n82 VSUBS 0.010986f
C140 B.n83 VSUBS 0.010986f
C141 B.n84 VSUBS 0.010986f
C142 B.n85 VSUBS 0.010986f
C143 B.n86 VSUBS 0.010986f
C144 B.n87 VSUBS 0.010986f
C145 B.n88 VSUBS 0.010986f
C146 B.n89 VSUBS 0.010986f
C147 B.n90 VSUBS 0.010986f
C148 B.n91 VSUBS 0.010986f
C149 B.n92 VSUBS 0.010986f
C150 B.n93 VSUBS 0.010986f
C151 B.n94 VSUBS 0.010986f
C152 B.n95 VSUBS 0.010986f
C153 B.n96 VSUBS 0.010986f
C154 B.n97 VSUBS 0.023493f
C155 B.n98 VSUBS 0.023493f
C156 B.n99 VSUBS 0.02465f
C157 B.n100 VSUBS 0.010986f
C158 B.n101 VSUBS 0.010986f
C159 B.n102 VSUBS 0.010986f
C160 B.n103 VSUBS 0.010986f
C161 B.n104 VSUBS 0.010986f
C162 B.n105 VSUBS 0.010986f
C163 B.n106 VSUBS 0.010986f
C164 B.n107 VSUBS 0.010986f
C165 B.n108 VSUBS 0.010986f
C166 B.n109 VSUBS 0.010339f
C167 B.n110 VSUBS 0.010986f
C168 B.n111 VSUBS 0.010986f
C169 B.n112 VSUBS 0.006139f
C170 B.n113 VSUBS 0.010986f
C171 B.n114 VSUBS 0.010986f
C172 B.n115 VSUBS 0.010986f
C173 B.n116 VSUBS 0.010986f
C174 B.n117 VSUBS 0.010986f
C175 B.n118 VSUBS 0.010986f
C176 B.n119 VSUBS 0.010986f
C177 B.n120 VSUBS 0.010986f
C178 B.n121 VSUBS 0.010986f
C179 B.n122 VSUBS 0.010986f
C180 B.n123 VSUBS 0.010986f
C181 B.n124 VSUBS 0.010986f
C182 B.n125 VSUBS 0.006139f
C183 B.n126 VSUBS 0.025452f
C184 B.n127 VSUBS 0.010339f
C185 B.n128 VSUBS 0.010986f
C186 B.n129 VSUBS 0.010986f
C187 B.n130 VSUBS 0.010986f
C188 B.n131 VSUBS 0.010986f
C189 B.n132 VSUBS 0.010986f
C190 B.n133 VSUBS 0.010986f
C191 B.n134 VSUBS 0.010986f
C192 B.n135 VSUBS 0.010986f
C193 B.n136 VSUBS 0.010986f
C194 B.n137 VSUBS 0.010986f
C195 B.n138 VSUBS 0.02465f
C196 B.n139 VSUBS 0.023493f
C197 B.n140 VSUBS 0.023493f
C198 B.n141 VSUBS 0.010986f
C199 B.n142 VSUBS 0.010986f
C200 B.n143 VSUBS 0.010986f
C201 B.n144 VSUBS 0.010986f
C202 B.n145 VSUBS 0.010986f
C203 B.n146 VSUBS 0.010986f
C204 B.n147 VSUBS 0.010986f
C205 B.n148 VSUBS 0.010986f
C206 B.n149 VSUBS 0.010986f
C207 B.n150 VSUBS 0.010986f
C208 B.n151 VSUBS 0.010986f
C209 B.n152 VSUBS 0.010986f
C210 B.n153 VSUBS 0.010986f
C211 B.n154 VSUBS 0.010986f
C212 B.n155 VSUBS 0.010986f
C213 B.n156 VSUBS 0.010986f
C214 B.n157 VSUBS 0.010986f
C215 B.n158 VSUBS 0.010986f
C216 B.n159 VSUBS 0.010986f
C217 B.n160 VSUBS 0.010986f
C218 B.n161 VSUBS 0.010986f
C219 B.n162 VSUBS 0.010986f
C220 B.n163 VSUBS 0.010986f
C221 B.n164 VSUBS 0.010986f
C222 B.n165 VSUBS 0.010986f
C223 B.n166 VSUBS 0.010986f
C224 B.n167 VSUBS 0.010986f
C225 B.n168 VSUBS 0.010986f
C226 B.n169 VSUBS 0.010986f
C227 B.n170 VSUBS 0.010986f
C228 B.n171 VSUBS 0.010986f
C229 B.n172 VSUBS 0.010986f
C230 B.n173 VSUBS 0.010986f
C231 B.n174 VSUBS 0.010986f
C232 B.n175 VSUBS 0.010986f
C233 B.n176 VSUBS 0.010986f
C234 B.n177 VSUBS 0.010986f
C235 B.n178 VSUBS 0.010986f
C236 B.n179 VSUBS 0.010986f
C237 B.n180 VSUBS 0.010986f
C238 B.n181 VSUBS 0.010986f
C239 B.n182 VSUBS 0.010986f
C240 B.n183 VSUBS 0.010986f
C241 B.n184 VSUBS 0.010986f
C242 B.n185 VSUBS 0.010986f
C243 B.n186 VSUBS 0.010986f
C244 B.n187 VSUBS 0.010986f
C245 B.n188 VSUBS 0.010986f
C246 B.n189 VSUBS 0.010986f
C247 B.n190 VSUBS 0.010986f
C248 B.n191 VSUBS 0.010986f
C249 B.n192 VSUBS 0.010986f
C250 B.n193 VSUBS 0.02493f
C251 B.n194 VSUBS 0.023493f
C252 B.n195 VSUBS 0.02465f
C253 B.n196 VSUBS 0.010986f
C254 B.n197 VSUBS 0.010986f
C255 B.n198 VSUBS 0.010986f
C256 B.n199 VSUBS 0.010986f
C257 B.n200 VSUBS 0.010986f
C258 B.n201 VSUBS 0.010986f
C259 B.n202 VSUBS 0.010986f
C260 B.n203 VSUBS 0.010986f
C261 B.n204 VSUBS 0.010986f
C262 B.n205 VSUBS 0.010339f
C263 B.n206 VSUBS 0.010986f
C264 B.n207 VSUBS 0.010986f
C265 B.n208 VSUBS 0.006139f
C266 B.n209 VSUBS 0.010986f
C267 B.n210 VSUBS 0.010986f
C268 B.n211 VSUBS 0.010986f
C269 B.n212 VSUBS 0.010986f
C270 B.n213 VSUBS 0.010986f
C271 B.n214 VSUBS 0.010986f
C272 B.n215 VSUBS 0.010986f
C273 B.n216 VSUBS 0.010986f
C274 B.n217 VSUBS 0.010986f
C275 B.n218 VSUBS 0.010986f
C276 B.n219 VSUBS 0.010986f
C277 B.n220 VSUBS 0.010986f
C278 B.n221 VSUBS 0.006139f
C279 B.n222 VSUBS 0.025452f
C280 B.n223 VSUBS 0.010339f
C281 B.n224 VSUBS 0.010986f
C282 B.n225 VSUBS 0.010986f
C283 B.n226 VSUBS 0.010986f
C284 B.n227 VSUBS 0.010986f
C285 B.n228 VSUBS 0.010986f
C286 B.n229 VSUBS 0.010986f
C287 B.n230 VSUBS 0.010986f
C288 B.n231 VSUBS 0.010986f
C289 B.n232 VSUBS 0.010986f
C290 B.n233 VSUBS 0.010986f
C291 B.n234 VSUBS 0.02465f
C292 B.n235 VSUBS 0.023493f
C293 B.n236 VSUBS 0.023493f
C294 B.n237 VSUBS 0.010986f
C295 B.n238 VSUBS 0.010986f
C296 B.n239 VSUBS 0.010986f
C297 B.n240 VSUBS 0.010986f
C298 B.n241 VSUBS 0.010986f
C299 B.n242 VSUBS 0.010986f
C300 B.n243 VSUBS 0.010986f
C301 B.n244 VSUBS 0.010986f
C302 B.n245 VSUBS 0.010986f
C303 B.n246 VSUBS 0.010986f
C304 B.n247 VSUBS 0.010986f
C305 B.n248 VSUBS 0.010986f
C306 B.n249 VSUBS 0.010986f
C307 B.n250 VSUBS 0.010986f
C308 B.n251 VSUBS 0.010986f
C309 B.n252 VSUBS 0.010986f
C310 B.n253 VSUBS 0.010986f
C311 B.n254 VSUBS 0.010986f
C312 B.n255 VSUBS 0.010986f
C313 B.n256 VSUBS 0.010986f
C314 B.n257 VSUBS 0.010986f
C315 B.n258 VSUBS 0.010986f
C316 B.n259 VSUBS 0.010986f
C317 B.n260 VSUBS 0.010986f
C318 B.n261 VSUBS 0.010986f
C319 B.n262 VSUBS 0.010986f
C320 B.n263 VSUBS 0.024875f
.ends

