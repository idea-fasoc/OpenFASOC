* NGSPICE file created from diff_pair_sample_1705.ext - technology: sky130A

.subckt diff_pair_sample_1705 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.2607 ps=1.91 w=1.58 l=1.92
X1 VDD1.t5 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.6162 ps=3.94 w=1.58 l=1.92
X2 VTAIL.t5 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.2607 ps=1.91 w=1.58 l=1.92
X3 VTAIL.t10 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.2607 ps=1.91 w=1.58 l=1.92
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=1.92
X5 VTAIL.t11 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.2607 ps=1.91 w=1.58 l=1.92
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=1.92
X7 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.2607 ps=1.91 w=1.58 l=1.92
X8 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.2607 ps=1.91 w=1.58 l=1.92
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=1.92
X10 VDD2.t2 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.6162 ps=3.94 w=1.58 l=1.92
X11 VDD2.t1 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.6162 ps=3.94 w=1.58 l=1.92
X12 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2607 pd=1.91 as=0.6162 ps=3.94 w=1.58 l=1.92
X13 VDD2.t0 VN.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.2607 ps=1.91 w=1.58 l=1.92
X14 VDD1.t0 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.2607 ps=1.91 w=1.58 l=1.92
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=1.92
R0 VN.n21 VN.n12 161.3
R1 VN.n20 VN.n19 161.3
R2 VN.n18 VN.n13 161.3
R3 VN.n17 VN.n16 161.3
R4 VN.n9 VN.n0 161.3
R5 VN.n8 VN.n7 161.3
R6 VN.n6 VN.n1 161.3
R7 VN.n5 VN.n4 161.3
R8 VN.n11 VN.n10 86.3164
R9 VN.n23 VN.n22 86.3164
R10 VN.n3 VN.n2 58.0791
R11 VN.n15 VN.n14 58.0791
R12 VN.n8 VN.n1 52.6866
R13 VN.n20 VN.n13 52.6866
R14 VN.n2 VN.t5 51.332
R15 VN.n14 VN.t3 51.332
R16 VN VN.n23 38.4717
R17 VN.n9 VN.n8 28.4674
R18 VN.n21 VN.n20 28.4674
R19 VN.n4 VN.n1 24.5923
R20 VN.n10 VN.n9 24.5923
R21 VN.n16 VN.n13 24.5923
R22 VN.n22 VN.n21 24.5923
R23 VN.n10 VN.t4 19.8328
R24 VN.n3 VN.t2 19.8328
R25 VN.n22 VN.t0 19.8328
R26 VN.n15 VN.t1 19.8328
R27 VN.n17 VN.n14 12.6034
R28 VN.n5 VN.n2 12.6034
R29 VN.n4 VN.n3 12.2964
R30 VN.n16 VN.n15 12.2964
R31 VN.n23 VN.n12 0.278335
R32 VN.n11 VN.n0 0.278335
R33 VN.n19 VN.n12 0.189894
R34 VN.n19 VN.n18 0.189894
R35 VN.n18 VN.n17 0.189894
R36 VN.n6 VN.n5 0.189894
R37 VN.n7 VN.n6 0.189894
R38 VN.n7 VN.n0 0.189894
R39 VN VN.n11 0.153485
R40 VTAIL.n11 VTAIL.t7 110.665
R41 VTAIL.n2 VTAIL.t4 110.665
R42 VTAIL.n10 VTAIL.t1 110.665
R43 VTAIL.n7 VTAIL.t8 110.665
R44 VTAIL.n1 VTAIL.n0 98.1339
R45 VTAIL.n4 VTAIL.n3 98.1339
R46 VTAIL.n9 VTAIL.n8 98.1339
R47 VTAIL.n6 VTAIL.n5 98.1339
R48 VTAIL.n6 VTAIL.n4 17.6083
R49 VTAIL.n11 VTAIL.n10 15.6686
R50 VTAIL.n0 VTAIL.t6 12.5321
R51 VTAIL.n0 VTAIL.t11 12.5321
R52 VTAIL.n3 VTAIL.t3 12.5321
R53 VTAIL.n3 VTAIL.t0 12.5321
R54 VTAIL.n8 VTAIL.t2 12.5321
R55 VTAIL.n8 VTAIL.t5 12.5321
R56 VTAIL.n5 VTAIL.t9 12.5321
R57 VTAIL.n5 VTAIL.t10 12.5321
R58 VTAIL.n7 VTAIL.n6 1.94016
R59 VTAIL.n10 VTAIL.n9 1.94016
R60 VTAIL.n4 VTAIL.n2 1.94016
R61 VTAIL.n9 VTAIL.n7 1.44016
R62 VTAIL.n2 VTAIL.n1 1.44016
R63 VTAIL VTAIL.n11 1.39705
R64 VTAIL VTAIL.n1 0.543603
R65 VDD2.n1 VDD2.t0 128.744
R66 VDD2.n2 VDD2.t5 127.344
R67 VDD2.n1 VDD2.n0 115.243
R68 VDD2 VDD2.n3 115.24
R69 VDD2.n2 VDD2.n1 31.3812
R70 VDD2.n3 VDD2.t4 12.5321
R71 VDD2.n3 VDD2.t2 12.5321
R72 VDD2.n0 VDD2.t3 12.5321
R73 VDD2.n0 VDD2.t1 12.5321
R74 VDD2 VDD2.n2 1.51343
R75 B.n386 B.n385 585
R76 B.n388 B.n86 585
R77 B.n391 B.n390 585
R78 B.n392 B.n85 585
R79 B.n394 B.n393 585
R80 B.n396 B.n84 585
R81 B.n399 B.n398 585
R82 B.n400 B.n83 585
R83 B.n402 B.n401 585
R84 B.n404 B.n82 585
R85 B.n407 B.n406 585
R86 B.n409 B.n79 585
R87 B.n411 B.n410 585
R88 B.n413 B.n78 585
R89 B.n416 B.n415 585
R90 B.n417 B.n77 585
R91 B.n419 B.n418 585
R92 B.n421 B.n76 585
R93 B.n424 B.n423 585
R94 B.n425 B.n72 585
R95 B.n427 B.n426 585
R96 B.n429 B.n71 585
R97 B.n432 B.n431 585
R98 B.n433 B.n70 585
R99 B.n435 B.n434 585
R100 B.n437 B.n69 585
R101 B.n440 B.n439 585
R102 B.n441 B.n68 585
R103 B.n443 B.n442 585
R104 B.n445 B.n67 585
R105 B.n448 B.n447 585
R106 B.n449 B.n66 585
R107 B.n384 B.n64 585
R108 B.n452 B.n64 585
R109 B.n383 B.n63 585
R110 B.n453 B.n63 585
R111 B.n382 B.n62 585
R112 B.n454 B.n62 585
R113 B.n381 B.n380 585
R114 B.n380 B.n58 585
R115 B.n379 B.n57 585
R116 B.n460 B.n57 585
R117 B.n378 B.n56 585
R118 B.n461 B.n56 585
R119 B.n377 B.n55 585
R120 B.n462 B.n55 585
R121 B.n376 B.n375 585
R122 B.n375 B.n51 585
R123 B.n374 B.n50 585
R124 B.n468 B.n50 585
R125 B.n373 B.n49 585
R126 B.n469 B.n49 585
R127 B.n372 B.n48 585
R128 B.n470 B.n48 585
R129 B.n371 B.n370 585
R130 B.n370 B.n44 585
R131 B.n369 B.n43 585
R132 B.n476 B.n43 585
R133 B.n368 B.n42 585
R134 B.n477 B.n42 585
R135 B.n367 B.n41 585
R136 B.n478 B.n41 585
R137 B.n366 B.n365 585
R138 B.n365 B.n37 585
R139 B.n364 B.n36 585
R140 B.n484 B.n36 585
R141 B.n363 B.n35 585
R142 B.n485 B.n35 585
R143 B.n362 B.n34 585
R144 B.n486 B.n34 585
R145 B.n361 B.n360 585
R146 B.n360 B.n30 585
R147 B.n359 B.n29 585
R148 B.n492 B.n29 585
R149 B.n358 B.n28 585
R150 B.n493 B.n28 585
R151 B.n357 B.n27 585
R152 B.n494 B.n27 585
R153 B.n356 B.n355 585
R154 B.n355 B.n23 585
R155 B.n354 B.n22 585
R156 B.n500 B.n22 585
R157 B.n353 B.n21 585
R158 B.n501 B.n21 585
R159 B.n352 B.n20 585
R160 B.n502 B.n20 585
R161 B.n351 B.n350 585
R162 B.n350 B.n16 585
R163 B.n349 B.n15 585
R164 B.n508 B.n15 585
R165 B.n348 B.n14 585
R166 B.n509 B.n14 585
R167 B.n347 B.n13 585
R168 B.n510 B.n13 585
R169 B.n346 B.n345 585
R170 B.n345 B.n12 585
R171 B.n344 B.n343 585
R172 B.n344 B.n8 585
R173 B.n342 B.n7 585
R174 B.n517 B.n7 585
R175 B.n341 B.n6 585
R176 B.n518 B.n6 585
R177 B.n340 B.n5 585
R178 B.n519 B.n5 585
R179 B.n339 B.n338 585
R180 B.n338 B.n4 585
R181 B.n337 B.n87 585
R182 B.n337 B.n336 585
R183 B.n327 B.n88 585
R184 B.n89 B.n88 585
R185 B.n329 B.n328 585
R186 B.n330 B.n329 585
R187 B.n326 B.n93 585
R188 B.n97 B.n93 585
R189 B.n325 B.n324 585
R190 B.n324 B.n323 585
R191 B.n95 B.n94 585
R192 B.n96 B.n95 585
R193 B.n316 B.n315 585
R194 B.n317 B.n316 585
R195 B.n314 B.n102 585
R196 B.n102 B.n101 585
R197 B.n313 B.n312 585
R198 B.n312 B.n311 585
R199 B.n104 B.n103 585
R200 B.n105 B.n104 585
R201 B.n304 B.n303 585
R202 B.n305 B.n304 585
R203 B.n302 B.n110 585
R204 B.n110 B.n109 585
R205 B.n301 B.n300 585
R206 B.n300 B.n299 585
R207 B.n112 B.n111 585
R208 B.n113 B.n112 585
R209 B.n292 B.n291 585
R210 B.n293 B.n292 585
R211 B.n290 B.n118 585
R212 B.n118 B.n117 585
R213 B.n289 B.n288 585
R214 B.n288 B.n287 585
R215 B.n120 B.n119 585
R216 B.n121 B.n120 585
R217 B.n280 B.n279 585
R218 B.n281 B.n280 585
R219 B.n278 B.n126 585
R220 B.n126 B.n125 585
R221 B.n277 B.n276 585
R222 B.n276 B.n275 585
R223 B.n128 B.n127 585
R224 B.n129 B.n128 585
R225 B.n268 B.n267 585
R226 B.n269 B.n268 585
R227 B.n266 B.n134 585
R228 B.n134 B.n133 585
R229 B.n265 B.n264 585
R230 B.n264 B.n263 585
R231 B.n136 B.n135 585
R232 B.n137 B.n136 585
R233 B.n256 B.n255 585
R234 B.n257 B.n256 585
R235 B.n254 B.n142 585
R236 B.n142 B.n141 585
R237 B.n253 B.n252 585
R238 B.n252 B.n251 585
R239 B.n144 B.n143 585
R240 B.n145 B.n144 585
R241 B.n244 B.n243 585
R242 B.n245 B.n244 585
R243 B.n242 B.n150 585
R244 B.n150 B.n149 585
R245 B.n241 B.n240 585
R246 B.n240 B.n239 585
R247 B.n236 B.n154 585
R248 B.n235 B.n234 585
R249 B.n232 B.n155 585
R250 B.n232 B.n153 585
R251 B.n231 B.n230 585
R252 B.n229 B.n228 585
R253 B.n227 B.n157 585
R254 B.n225 B.n224 585
R255 B.n223 B.n158 585
R256 B.n222 B.n221 585
R257 B.n219 B.n159 585
R258 B.n217 B.n216 585
R259 B.n214 B.n160 585
R260 B.n213 B.n212 585
R261 B.n210 B.n163 585
R262 B.n208 B.n207 585
R263 B.n206 B.n164 585
R264 B.n205 B.n204 585
R265 B.n202 B.n165 585
R266 B.n200 B.n199 585
R267 B.n198 B.n166 585
R268 B.n197 B.n196 585
R269 B.n194 B.n193 585
R270 B.n192 B.n191 585
R271 B.n190 B.n171 585
R272 B.n188 B.n187 585
R273 B.n186 B.n172 585
R274 B.n185 B.n184 585
R275 B.n182 B.n173 585
R276 B.n180 B.n179 585
R277 B.n178 B.n174 585
R278 B.n177 B.n176 585
R279 B.n152 B.n151 585
R280 B.n153 B.n152 585
R281 B.n238 B.n237 585
R282 B.n239 B.n238 585
R283 B.n148 B.n147 585
R284 B.n149 B.n148 585
R285 B.n247 B.n246 585
R286 B.n246 B.n245 585
R287 B.n248 B.n146 585
R288 B.n146 B.n145 585
R289 B.n250 B.n249 585
R290 B.n251 B.n250 585
R291 B.n140 B.n139 585
R292 B.n141 B.n140 585
R293 B.n259 B.n258 585
R294 B.n258 B.n257 585
R295 B.n260 B.n138 585
R296 B.n138 B.n137 585
R297 B.n262 B.n261 585
R298 B.n263 B.n262 585
R299 B.n132 B.n131 585
R300 B.n133 B.n132 585
R301 B.n271 B.n270 585
R302 B.n270 B.n269 585
R303 B.n272 B.n130 585
R304 B.n130 B.n129 585
R305 B.n274 B.n273 585
R306 B.n275 B.n274 585
R307 B.n124 B.n123 585
R308 B.n125 B.n124 585
R309 B.n283 B.n282 585
R310 B.n282 B.n281 585
R311 B.n284 B.n122 585
R312 B.n122 B.n121 585
R313 B.n286 B.n285 585
R314 B.n287 B.n286 585
R315 B.n116 B.n115 585
R316 B.n117 B.n116 585
R317 B.n295 B.n294 585
R318 B.n294 B.n293 585
R319 B.n296 B.n114 585
R320 B.n114 B.n113 585
R321 B.n298 B.n297 585
R322 B.n299 B.n298 585
R323 B.n108 B.n107 585
R324 B.n109 B.n108 585
R325 B.n307 B.n306 585
R326 B.n306 B.n305 585
R327 B.n308 B.n106 585
R328 B.n106 B.n105 585
R329 B.n310 B.n309 585
R330 B.n311 B.n310 585
R331 B.n100 B.n99 585
R332 B.n101 B.n100 585
R333 B.n319 B.n318 585
R334 B.n318 B.n317 585
R335 B.n320 B.n98 585
R336 B.n98 B.n96 585
R337 B.n322 B.n321 585
R338 B.n323 B.n322 585
R339 B.n92 B.n91 585
R340 B.n97 B.n92 585
R341 B.n332 B.n331 585
R342 B.n331 B.n330 585
R343 B.n333 B.n90 585
R344 B.n90 B.n89 585
R345 B.n335 B.n334 585
R346 B.n336 B.n335 585
R347 B.n3 B.n0 585
R348 B.n4 B.n3 585
R349 B.n516 B.n1 585
R350 B.n517 B.n516 585
R351 B.n515 B.n514 585
R352 B.n515 B.n8 585
R353 B.n513 B.n9 585
R354 B.n12 B.n9 585
R355 B.n512 B.n511 585
R356 B.n511 B.n510 585
R357 B.n11 B.n10 585
R358 B.n509 B.n11 585
R359 B.n507 B.n506 585
R360 B.n508 B.n507 585
R361 B.n505 B.n17 585
R362 B.n17 B.n16 585
R363 B.n504 B.n503 585
R364 B.n503 B.n502 585
R365 B.n19 B.n18 585
R366 B.n501 B.n19 585
R367 B.n499 B.n498 585
R368 B.n500 B.n499 585
R369 B.n497 B.n24 585
R370 B.n24 B.n23 585
R371 B.n496 B.n495 585
R372 B.n495 B.n494 585
R373 B.n26 B.n25 585
R374 B.n493 B.n26 585
R375 B.n491 B.n490 585
R376 B.n492 B.n491 585
R377 B.n489 B.n31 585
R378 B.n31 B.n30 585
R379 B.n488 B.n487 585
R380 B.n487 B.n486 585
R381 B.n33 B.n32 585
R382 B.n485 B.n33 585
R383 B.n483 B.n482 585
R384 B.n484 B.n483 585
R385 B.n481 B.n38 585
R386 B.n38 B.n37 585
R387 B.n480 B.n479 585
R388 B.n479 B.n478 585
R389 B.n40 B.n39 585
R390 B.n477 B.n40 585
R391 B.n475 B.n474 585
R392 B.n476 B.n475 585
R393 B.n473 B.n45 585
R394 B.n45 B.n44 585
R395 B.n472 B.n471 585
R396 B.n471 B.n470 585
R397 B.n47 B.n46 585
R398 B.n469 B.n47 585
R399 B.n467 B.n466 585
R400 B.n468 B.n467 585
R401 B.n465 B.n52 585
R402 B.n52 B.n51 585
R403 B.n464 B.n463 585
R404 B.n463 B.n462 585
R405 B.n54 B.n53 585
R406 B.n461 B.n54 585
R407 B.n459 B.n458 585
R408 B.n460 B.n459 585
R409 B.n457 B.n59 585
R410 B.n59 B.n58 585
R411 B.n456 B.n455 585
R412 B.n455 B.n454 585
R413 B.n61 B.n60 585
R414 B.n453 B.n61 585
R415 B.n451 B.n450 585
R416 B.n452 B.n451 585
R417 B.n520 B.n519 585
R418 B.n518 B.n2 585
R419 B.n451 B.n66 473.281
R420 B.n386 B.n64 473.281
R421 B.n240 B.n152 473.281
R422 B.n238 B.n154 473.281
R423 B.n387 B.n65 256.663
R424 B.n389 B.n65 256.663
R425 B.n395 B.n65 256.663
R426 B.n397 B.n65 256.663
R427 B.n403 B.n65 256.663
R428 B.n405 B.n65 256.663
R429 B.n412 B.n65 256.663
R430 B.n414 B.n65 256.663
R431 B.n420 B.n65 256.663
R432 B.n422 B.n65 256.663
R433 B.n428 B.n65 256.663
R434 B.n430 B.n65 256.663
R435 B.n436 B.n65 256.663
R436 B.n438 B.n65 256.663
R437 B.n444 B.n65 256.663
R438 B.n446 B.n65 256.663
R439 B.n233 B.n153 256.663
R440 B.n156 B.n153 256.663
R441 B.n226 B.n153 256.663
R442 B.n220 B.n153 256.663
R443 B.n218 B.n153 256.663
R444 B.n211 B.n153 256.663
R445 B.n209 B.n153 256.663
R446 B.n203 B.n153 256.663
R447 B.n201 B.n153 256.663
R448 B.n195 B.n153 256.663
R449 B.n170 B.n153 256.663
R450 B.n189 B.n153 256.663
R451 B.n183 B.n153 256.663
R452 B.n181 B.n153 256.663
R453 B.n175 B.n153 256.663
R454 B.n522 B.n521 256.663
R455 B.n73 B.t10 226.555
R456 B.n80 B.t6 226.555
R457 B.n167 B.t13 226.555
R458 B.n161 B.t17 226.555
R459 B.n239 B.n153 207.002
R460 B.n452 B.n65 207.002
R461 B.n447 B.n445 163.367
R462 B.n443 B.n68 163.367
R463 B.n439 B.n437 163.367
R464 B.n435 B.n70 163.367
R465 B.n431 B.n429 163.367
R466 B.n427 B.n72 163.367
R467 B.n423 B.n421 163.367
R468 B.n419 B.n77 163.367
R469 B.n415 B.n413 163.367
R470 B.n411 B.n79 163.367
R471 B.n406 B.n404 163.367
R472 B.n402 B.n83 163.367
R473 B.n398 B.n396 163.367
R474 B.n394 B.n85 163.367
R475 B.n390 B.n388 163.367
R476 B.n240 B.n150 163.367
R477 B.n244 B.n150 163.367
R478 B.n244 B.n144 163.367
R479 B.n252 B.n144 163.367
R480 B.n252 B.n142 163.367
R481 B.n256 B.n142 163.367
R482 B.n256 B.n136 163.367
R483 B.n264 B.n136 163.367
R484 B.n264 B.n134 163.367
R485 B.n268 B.n134 163.367
R486 B.n268 B.n128 163.367
R487 B.n276 B.n128 163.367
R488 B.n276 B.n126 163.367
R489 B.n280 B.n126 163.367
R490 B.n280 B.n120 163.367
R491 B.n288 B.n120 163.367
R492 B.n288 B.n118 163.367
R493 B.n292 B.n118 163.367
R494 B.n292 B.n112 163.367
R495 B.n300 B.n112 163.367
R496 B.n300 B.n110 163.367
R497 B.n304 B.n110 163.367
R498 B.n304 B.n104 163.367
R499 B.n312 B.n104 163.367
R500 B.n312 B.n102 163.367
R501 B.n316 B.n102 163.367
R502 B.n316 B.n95 163.367
R503 B.n324 B.n95 163.367
R504 B.n324 B.n93 163.367
R505 B.n329 B.n93 163.367
R506 B.n329 B.n88 163.367
R507 B.n337 B.n88 163.367
R508 B.n338 B.n337 163.367
R509 B.n338 B.n5 163.367
R510 B.n6 B.n5 163.367
R511 B.n7 B.n6 163.367
R512 B.n344 B.n7 163.367
R513 B.n345 B.n344 163.367
R514 B.n345 B.n13 163.367
R515 B.n14 B.n13 163.367
R516 B.n15 B.n14 163.367
R517 B.n350 B.n15 163.367
R518 B.n350 B.n20 163.367
R519 B.n21 B.n20 163.367
R520 B.n22 B.n21 163.367
R521 B.n355 B.n22 163.367
R522 B.n355 B.n27 163.367
R523 B.n28 B.n27 163.367
R524 B.n29 B.n28 163.367
R525 B.n360 B.n29 163.367
R526 B.n360 B.n34 163.367
R527 B.n35 B.n34 163.367
R528 B.n36 B.n35 163.367
R529 B.n365 B.n36 163.367
R530 B.n365 B.n41 163.367
R531 B.n42 B.n41 163.367
R532 B.n43 B.n42 163.367
R533 B.n370 B.n43 163.367
R534 B.n370 B.n48 163.367
R535 B.n49 B.n48 163.367
R536 B.n50 B.n49 163.367
R537 B.n375 B.n50 163.367
R538 B.n375 B.n55 163.367
R539 B.n56 B.n55 163.367
R540 B.n57 B.n56 163.367
R541 B.n380 B.n57 163.367
R542 B.n380 B.n62 163.367
R543 B.n63 B.n62 163.367
R544 B.n64 B.n63 163.367
R545 B.n234 B.n232 163.367
R546 B.n232 B.n231 163.367
R547 B.n228 B.n227 163.367
R548 B.n225 B.n158 163.367
R549 B.n221 B.n219 163.367
R550 B.n217 B.n160 163.367
R551 B.n212 B.n210 163.367
R552 B.n208 B.n164 163.367
R553 B.n204 B.n202 163.367
R554 B.n200 B.n166 163.367
R555 B.n196 B.n194 163.367
R556 B.n191 B.n190 163.367
R557 B.n188 B.n172 163.367
R558 B.n184 B.n182 163.367
R559 B.n180 B.n174 163.367
R560 B.n176 B.n152 163.367
R561 B.n238 B.n148 163.367
R562 B.n246 B.n148 163.367
R563 B.n246 B.n146 163.367
R564 B.n250 B.n146 163.367
R565 B.n250 B.n140 163.367
R566 B.n258 B.n140 163.367
R567 B.n258 B.n138 163.367
R568 B.n262 B.n138 163.367
R569 B.n262 B.n132 163.367
R570 B.n270 B.n132 163.367
R571 B.n270 B.n130 163.367
R572 B.n274 B.n130 163.367
R573 B.n274 B.n124 163.367
R574 B.n282 B.n124 163.367
R575 B.n282 B.n122 163.367
R576 B.n286 B.n122 163.367
R577 B.n286 B.n116 163.367
R578 B.n294 B.n116 163.367
R579 B.n294 B.n114 163.367
R580 B.n298 B.n114 163.367
R581 B.n298 B.n108 163.367
R582 B.n306 B.n108 163.367
R583 B.n306 B.n106 163.367
R584 B.n310 B.n106 163.367
R585 B.n310 B.n100 163.367
R586 B.n318 B.n100 163.367
R587 B.n318 B.n98 163.367
R588 B.n322 B.n98 163.367
R589 B.n322 B.n92 163.367
R590 B.n331 B.n92 163.367
R591 B.n331 B.n90 163.367
R592 B.n335 B.n90 163.367
R593 B.n335 B.n3 163.367
R594 B.n520 B.n3 163.367
R595 B.n516 B.n2 163.367
R596 B.n516 B.n515 163.367
R597 B.n515 B.n9 163.367
R598 B.n511 B.n9 163.367
R599 B.n511 B.n11 163.367
R600 B.n507 B.n11 163.367
R601 B.n507 B.n17 163.367
R602 B.n503 B.n17 163.367
R603 B.n503 B.n19 163.367
R604 B.n499 B.n19 163.367
R605 B.n499 B.n24 163.367
R606 B.n495 B.n24 163.367
R607 B.n495 B.n26 163.367
R608 B.n491 B.n26 163.367
R609 B.n491 B.n31 163.367
R610 B.n487 B.n31 163.367
R611 B.n487 B.n33 163.367
R612 B.n483 B.n33 163.367
R613 B.n483 B.n38 163.367
R614 B.n479 B.n38 163.367
R615 B.n479 B.n40 163.367
R616 B.n475 B.n40 163.367
R617 B.n475 B.n45 163.367
R618 B.n471 B.n45 163.367
R619 B.n471 B.n47 163.367
R620 B.n467 B.n47 163.367
R621 B.n467 B.n52 163.367
R622 B.n463 B.n52 163.367
R623 B.n463 B.n54 163.367
R624 B.n459 B.n54 163.367
R625 B.n459 B.n59 163.367
R626 B.n455 B.n59 163.367
R627 B.n455 B.n61 163.367
R628 B.n451 B.n61 163.367
R629 B.n80 B.t8 151.858
R630 B.n167 B.t16 151.858
R631 B.n73 B.t11 151.858
R632 B.n161 B.t19 151.858
R633 B.n239 B.n149 109.118
R634 B.n245 B.n149 109.118
R635 B.n245 B.n145 109.118
R636 B.n251 B.n145 109.118
R637 B.n251 B.n141 109.118
R638 B.n257 B.n141 109.118
R639 B.n263 B.n137 109.118
R640 B.n263 B.n133 109.118
R641 B.n269 B.n133 109.118
R642 B.n269 B.n129 109.118
R643 B.n275 B.n129 109.118
R644 B.n275 B.n125 109.118
R645 B.n281 B.n125 109.118
R646 B.n281 B.n121 109.118
R647 B.n287 B.n121 109.118
R648 B.n293 B.n117 109.118
R649 B.n293 B.n113 109.118
R650 B.n299 B.n113 109.118
R651 B.n299 B.n109 109.118
R652 B.n305 B.n109 109.118
R653 B.n311 B.n105 109.118
R654 B.n311 B.n101 109.118
R655 B.n317 B.n101 109.118
R656 B.n317 B.n96 109.118
R657 B.n323 B.n96 109.118
R658 B.n323 B.n97 109.118
R659 B.n330 B.n89 109.118
R660 B.n336 B.n89 109.118
R661 B.n336 B.n4 109.118
R662 B.n519 B.n4 109.118
R663 B.n519 B.n518 109.118
R664 B.n518 B.n517 109.118
R665 B.n517 B.n8 109.118
R666 B.n12 B.n8 109.118
R667 B.n510 B.n12 109.118
R668 B.n509 B.n508 109.118
R669 B.n508 B.n16 109.118
R670 B.n502 B.n16 109.118
R671 B.n502 B.n501 109.118
R672 B.n501 B.n500 109.118
R673 B.n500 B.n23 109.118
R674 B.n494 B.n493 109.118
R675 B.n493 B.n492 109.118
R676 B.n492 B.n30 109.118
R677 B.n486 B.n30 109.118
R678 B.n486 B.n485 109.118
R679 B.n484 B.n37 109.118
R680 B.n478 B.n37 109.118
R681 B.n478 B.n477 109.118
R682 B.n477 B.n476 109.118
R683 B.n476 B.n44 109.118
R684 B.n470 B.n44 109.118
R685 B.n470 B.n469 109.118
R686 B.n469 B.n468 109.118
R687 B.n468 B.n51 109.118
R688 B.n462 B.n461 109.118
R689 B.n461 B.n460 109.118
R690 B.n460 B.n58 109.118
R691 B.n454 B.n58 109.118
R692 B.n454 B.n453 109.118
R693 B.n453 B.n452 109.118
R694 B.n81 B.t9 108.222
R695 B.n168 B.t15 108.222
R696 B.n74 B.t12 108.222
R697 B.n162 B.t18 108.222
R698 B.n305 B.t0 105.909
R699 B.n494 B.t5 105.909
R700 B.n446 B.n66 71.676
R701 B.n445 B.n444 71.676
R702 B.n438 B.n68 71.676
R703 B.n437 B.n436 71.676
R704 B.n430 B.n70 71.676
R705 B.n429 B.n428 71.676
R706 B.n422 B.n72 71.676
R707 B.n421 B.n420 71.676
R708 B.n414 B.n77 71.676
R709 B.n413 B.n412 71.676
R710 B.n405 B.n79 71.676
R711 B.n404 B.n403 71.676
R712 B.n397 B.n83 71.676
R713 B.n396 B.n395 71.676
R714 B.n389 B.n85 71.676
R715 B.n388 B.n387 71.676
R716 B.n387 B.n386 71.676
R717 B.n390 B.n389 71.676
R718 B.n395 B.n394 71.676
R719 B.n398 B.n397 71.676
R720 B.n403 B.n402 71.676
R721 B.n406 B.n405 71.676
R722 B.n412 B.n411 71.676
R723 B.n415 B.n414 71.676
R724 B.n420 B.n419 71.676
R725 B.n423 B.n422 71.676
R726 B.n428 B.n427 71.676
R727 B.n431 B.n430 71.676
R728 B.n436 B.n435 71.676
R729 B.n439 B.n438 71.676
R730 B.n444 B.n443 71.676
R731 B.n447 B.n446 71.676
R732 B.n233 B.n154 71.676
R733 B.n231 B.n156 71.676
R734 B.n227 B.n226 71.676
R735 B.n220 B.n158 71.676
R736 B.n219 B.n218 71.676
R737 B.n211 B.n160 71.676
R738 B.n210 B.n209 71.676
R739 B.n203 B.n164 71.676
R740 B.n202 B.n201 71.676
R741 B.n195 B.n166 71.676
R742 B.n194 B.n170 71.676
R743 B.n190 B.n189 71.676
R744 B.n183 B.n172 71.676
R745 B.n182 B.n181 71.676
R746 B.n175 B.n174 71.676
R747 B.n234 B.n233 71.676
R748 B.n228 B.n156 71.676
R749 B.n226 B.n225 71.676
R750 B.n221 B.n220 71.676
R751 B.n218 B.n217 71.676
R752 B.n212 B.n211 71.676
R753 B.n209 B.n208 71.676
R754 B.n204 B.n203 71.676
R755 B.n201 B.n200 71.676
R756 B.n196 B.n195 71.676
R757 B.n191 B.n170 71.676
R758 B.n189 B.n188 71.676
R759 B.n184 B.n183 71.676
R760 B.n181 B.n180 71.676
R761 B.n176 B.n175 71.676
R762 B.n521 B.n520 71.676
R763 B.n521 B.n2 71.676
R764 B.t3 B.n117 70.6059
R765 B.n485 B.t1 70.6059
R766 B.n97 B.t4 64.1872
R767 B.t2 B.n509 64.1872
R768 B.n75 B.n74 59.5399
R769 B.n408 B.n81 59.5399
R770 B.n169 B.n168 59.5399
R771 B.n215 B.n162 59.5399
R772 B.n257 B.t14 57.7686
R773 B.n462 B.t7 57.7686
R774 B.t14 B.n137 51.3499
R775 B.t7 B.n51 51.3499
R776 B.n330 B.t4 44.9312
R777 B.n510 B.t2 44.9312
R778 B.n74 B.n73 43.6369
R779 B.n81 B.n80 43.6369
R780 B.n168 B.n167 43.6369
R781 B.n162 B.n161 43.6369
R782 B.n287 B.t3 38.5125
R783 B.t1 B.n484 38.5125
R784 B.n237 B.n236 30.7517
R785 B.n241 B.n151 30.7517
R786 B.n385 B.n384 30.7517
R787 B.n450 B.n449 30.7517
R788 B B.n522 18.0485
R789 B.n237 B.n147 10.6151
R790 B.n247 B.n147 10.6151
R791 B.n248 B.n247 10.6151
R792 B.n249 B.n248 10.6151
R793 B.n249 B.n139 10.6151
R794 B.n259 B.n139 10.6151
R795 B.n260 B.n259 10.6151
R796 B.n261 B.n260 10.6151
R797 B.n261 B.n131 10.6151
R798 B.n271 B.n131 10.6151
R799 B.n272 B.n271 10.6151
R800 B.n273 B.n272 10.6151
R801 B.n273 B.n123 10.6151
R802 B.n283 B.n123 10.6151
R803 B.n284 B.n283 10.6151
R804 B.n285 B.n284 10.6151
R805 B.n285 B.n115 10.6151
R806 B.n295 B.n115 10.6151
R807 B.n296 B.n295 10.6151
R808 B.n297 B.n296 10.6151
R809 B.n297 B.n107 10.6151
R810 B.n307 B.n107 10.6151
R811 B.n308 B.n307 10.6151
R812 B.n309 B.n308 10.6151
R813 B.n309 B.n99 10.6151
R814 B.n319 B.n99 10.6151
R815 B.n320 B.n319 10.6151
R816 B.n321 B.n320 10.6151
R817 B.n321 B.n91 10.6151
R818 B.n332 B.n91 10.6151
R819 B.n333 B.n332 10.6151
R820 B.n334 B.n333 10.6151
R821 B.n334 B.n0 10.6151
R822 B.n236 B.n235 10.6151
R823 B.n235 B.n155 10.6151
R824 B.n230 B.n155 10.6151
R825 B.n230 B.n229 10.6151
R826 B.n229 B.n157 10.6151
R827 B.n224 B.n157 10.6151
R828 B.n224 B.n223 10.6151
R829 B.n223 B.n222 10.6151
R830 B.n222 B.n159 10.6151
R831 B.n216 B.n159 10.6151
R832 B.n214 B.n213 10.6151
R833 B.n213 B.n163 10.6151
R834 B.n207 B.n163 10.6151
R835 B.n207 B.n206 10.6151
R836 B.n206 B.n205 10.6151
R837 B.n205 B.n165 10.6151
R838 B.n199 B.n165 10.6151
R839 B.n199 B.n198 10.6151
R840 B.n198 B.n197 10.6151
R841 B.n193 B.n192 10.6151
R842 B.n192 B.n171 10.6151
R843 B.n187 B.n171 10.6151
R844 B.n187 B.n186 10.6151
R845 B.n186 B.n185 10.6151
R846 B.n185 B.n173 10.6151
R847 B.n179 B.n173 10.6151
R848 B.n179 B.n178 10.6151
R849 B.n178 B.n177 10.6151
R850 B.n177 B.n151 10.6151
R851 B.n242 B.n241 10.6151
R852 B.n243 B.n242 10.6151
R853 B.n243 B.n143 10.6151
R854 B.n253 B.n143 10.6151
R855 B.n254 B.n253 10.6151
R856 B.n255 B.n254 10.6151
R857 B.n255 B.n135 10.6151
R858 B.n265 B.n135 10.6151
R859 B.n266 B.n265 10.6151
R860 B.n267 B.n266 10.6151
R861 B.n267 B.n127 10.6151
R862 B.n277 B.n127 10.6151
R863 B.n278 B.n277 10.6151
R864 B.n279 B.n278 10.6151
R865 B.n279 B.n119 10.6151
R866 B.n289 B.n119 10.6151
R867 B.n290 B.n289 10.6151
R868 B.n291 B.n290 10.6151
R869 B.n291 B.n111 10.6151
R870 B.n301 B.n111 10.6151
R871 B.n302 B.n301 10.6151
R872 B.n303 B.n302 10.6151
R873 B.n303 B.n103 10.6151
R874 B.n313 B.n103 10.6151
R875 B.n314 B.n313 10.6151
R876 B.n315 B.n314 10.6151
R877 B.n315 B.n94 10.6151
R878 B.n325 B.n94 10.6151
R879 B.n326 B.n325 10.6151
R880 B.n328 B.n326 10.6151
R881 B.n328 B.n327 10.6151
R882 B.n327 B.n87 10.6151
R883 B.n339 B.n87 10.6151
R884 B.n340 B.n339 10.6151
R885 B.n341 B.n340 10.6151
R886 B.n342 B.n341 10.6151
R887 B.n343 B.n342 10.6151
R888 B.n346 B.n343 10.6151
R889 B.n347 B.n346 10.6151
R890 B.n348 B.n347 10.6151
R891 B.n349 B.n348 10.6151
R892 B.n351 B.n349 10.6151
R893 B.n352 B.n351 10.6151
R894 B.n353 B.n352 10.6151
R895 B.n354 B.n353 10.6151
R896 B.n356 B.n354 10.6151
R897 B.n357 B.n356 10.6151
R898 B.n358 B.n357 10.6151
R899 B.n359 B.n358 10.6151
R900 B.n361 B.n359 10.6151
R901 B.n362 B.n361 10.6151
R902 B.n363 B.n362 10.6151
R903 B.n364 B.n363 10.6151
R904 B.n366 B.n364 10.6151
R905 B.n367 B.n366 10.6151
R906 B.n368 B.n367 10.6151
R907 B.n369 B.n368 10.6151
R908 B.n371 B.n369 10.6151
R909 B.n372 B.n371 10.6151
R910 B.n373 B.n372 10.6151
R911 B.n374 B.n373 10.6151
R912 B.n376 B.n374 10.6151
R913 B.n377 B.n376 10.6151
R914 B.n378 B.n377 10.6151
R915 B.n379 B.n378 10.6151
R916 B.n381 B.n379 10.6151
R917 B.n382 B.n381 10.6151
R918 B.n383 B.n382 10.6151
R919 B.n384 B.n383 10.6151
R920 B.n514 B.n1 10.6151
R921 B.n514 B.n513 10.6151
R922 B.n513 B.n512 10.6151
R923 B.n512 B.n10 10.6151
R924 B.n506 B.n10 10.6151
R925 B.n506 B.n505 10.6151
R926 B.n505 B.n504 10.6151
R927 B.n504 B.n18 10.6151
R928 B.n498 B.n18 10.6151
R929 B.n498 B.n497 10.6151
R930 B.n497 B.n496 10.6151
R931 B.n496 B.n25 10.6151
R932 B.n490 B.n25 10.6151
R933 B.n490 B.n489 10.6151
R934 B.n489 B.n488 10.6151
R935 B.n488 B.n32 10.6151
R936 B.n482 B.n32 10.6151
R937 B.n482 B.n481 10.6151
R938 B.n481 B.n480 10.6151
R939 B.n480 B.n39 10.6151
R940 B.n474 B.n39 10.6151
R941 B.n474 B.n473 10.6151
R942 B.n473 B.n472 10.6151
R943 B.n472 B.n46 10.6151
R944 B.n466 B.n46 10.6151
R945 B.n466 B.n465 10.6151
R946 B.n465 B.n464 10.6151
R947 B.n464 B.n53 10.6151
R948 B.n458 B.n53 10.6151
R949 B.n458 B.n457 10.6151
R950 B.n457 B.n456 10.6151
R951 B.n456 B.n60 10.6151
R952 B.n450 B.n60 10.6151
R953 B.n449 B.n448 10.6151
R954 B.n448 B.n67 10.6151
R955 B.n442 B.n67 10.6151
R956 B.n442 B.n441 10.6151
R957 B.n441 B.n440 10.6151
R958 B.n440 B.n69 10.6151
R959 B.n434 B.n69 10.6151
R960 B.n434 B.n433 10.6151
R961 B.n433 B.n432 10.6151
R962 B.n432 B.n71 10.6151
R963 B.n426 B.n425 10.6151
R964 B.n425 B.n424 10.6151
R965 B.n424 B.n76 10.6151
R966 B.n418 B.n76 10.6151
R967 B.n418 B.n417 10.6151
R968 B.n417 B.n416 10.6151
R969 B.n416 B.n78 10.6151
R970 B.n410 B.n78 10.6151
R971 B.n410 B.n409 10.6151
R972 B.n407 B.n82 10.6151
R973 B.n401 B.n82 10.6151
R974 B.n401 B.n400 10.6151
R975 B.n400 B.n399 10.6151
R976 B.n399 B.n84 10.6151
R977 B.n393 B.n84 10.6151
R978 B.n393 B.n392 10.6151
R979 B.n392 B.n391 10.6151
R980 B.n391 B.n86 10.6151
R981 B.n385 B.n86 10.6151
R982 B.n216 B.n215 9.36635
R983 B.n193 B.n169 9.36635
R984 B.n75 B.n71 9.36635
R985 B.n408 B.n407 9.36635
R986 B.n522 B.n0 8.11757
R987 B.n522 B.n1 8.11757
R988 B.t0 B.n105 3.20984
R989 B.t5 B.n23 3.20984
R990 B.n215 B.n214 1.24928
R991 B.n197 B.n169 1.24928
R992 B.n426 B.n75 1.24928
R993 B.n409 B.n408 1.24928
R994 VP.n9 VP.n8 161.3
R995 VP.n10 VP.n5 161.3
R996 VP.n12 VP.n11 161.3
R997 VP.n13 VP.n4 161.3
R998 VP.n30 VP.n0 161.3
R999 VP.n29 VP.n28 161.3
R1000 VP.n27 VP.n1 161.3
R1001 VP.n26 VP.n25 161.3
R1002 VP.n23 VP.n2 161.3
R1003 VP.n22 VP.n21 161.3
R1004 VP.n20 VP.n3 161.3
R1005 VP.n19 VP.n18 161.3
R1006 VP.n17 VP.n16 86.3164
R1007 VP.n32 VP.n31 86.3164
R1008 VP.n15 VP.n14 86.3164
R1009 VP.n7 VP.n6 58.0791
R1010 VP.n22 VP.n3 52.6866
R1011 VP.n29 VP.n1 52.6866
R1012 VP.n12 VP.n5 52.6866
R1013 VP.n6 VP.t2 51.332
R1014 VP.n16 VP.n15 38.1928
R1015 VP.n18 VP.n3 28.4674
R1016 VP.n30 VP.n29 28.4674
R1017 VP.n13 VP.n12 28.4674
R1018 VP.n18 VP.n17 24.5923
R1019 VP.n23 VP.n22 24.5923
R1020 VP.n25 VP.n1 24.5923
R1021 VP.n31 VP.n30 24.5923
R1022 VP.n14 VP.n13 24.5923
R1023 VP.n8 VP.n5 24.5923
R1024 VP.n31 VP.t0 19.8328
R1025 VP.n17 VP.t5 19.8328
R1026 VP.n24 VP.t3 19.8328
R1027 VP.n14 VP.t4 19.8328
R1028 VP.n7 VP.t1 19.8328
R1029 VP.n9 VP.n6 12.6034
R1030 VP.n24 VP.n23 12.2964
R1031 VP.n25 VP.n24 12.2964
R1032 VP.n8 VP.n7 12.2964
R1033 VP.n15 VP.n4 0.278335
R1034 VP.n19 VP.n16 0.278335
R1035 VP.n32 VP.n0 0.278335
R1036 VP.n10 VP.n9 0.189894
R1037 VP.n11 VP.n10 0.189894
R1038 VP.n11 VP.n4 0.189894
R1039 VP.n20 VP.n19 0.189894
R1040 VP.n21 VP.n20 0.189894
R1041 VP.n21 VP.n2 0.189894
R1042 VP.n26 VP.n2 0.189894
R1043 VP.n27 VP.n26 0.189894
R1044 VP.n28 VP.n27 0.189894
R1045 VP.n28 VP.n0 0.189894
R1046 VP VP.n32 0.153485
R1047 VDD1 VDD1.t3 128.857
R1048 VDD1.n1 VDD1.t0 128.744
R1049 VDD1.n1 VDD1.n0 115.243
R1050 VDD1.n3 VDD1.n2 114.812
R1051 VDD1.n3 VDD1.n1 32.9341
R1052 VDD1.n2 VDD1.t4 12.5321
R1053 VDD1.n2 VDD1.t1 12.5321
R1054 VDD1.n0 VDD1.t2 12.5321
R1055 VDD1.n0 VDD1.t5 12.5321
R1056 VDD1 VDD1.n3 0.427224
C0 VDD1 VP 1.40266f
C1 VDD2 VP 0.408162f
C2 VN VTAIL 1.81772f
C3 VDD1 VDD2 1.16467f
C4 VP VTAIL 1.83186f
C5 VP VN 4.34002f
C6 VDD1 VTAIL 3.47748f
C7 VDD2 VTAIL 3.52603f
C8 VDD1 VN 0.157162f
C9 VDD2 VN 1.15415f
C10 VDD2 B 3.440033f
C11 VDD1 B 3.69623f
C12 VTAIL B 2.835236f
C13 VN B 9.453265f
C14 VP B 8.520335f
C15 VDD1.t3 B 0.164246f
C16 VDD1.t0 B 0.163986f
C17 VDD1.t2 B 0.020911f
C18 VDD1.t5 B 0.020911f
C19 VDD1.n0 B 0.120883f
C20 VDD1.n1 B 1.34654f
C21 VDD1.t4 B 0.020911f
C22 VDD1.t1 B 0.020911f
C23 VDD1.n2 B 0.119925f
C24 VDD1.n3 B 1.17334f
C25 VP.n0 B 0.029146f
C26 VP.t0 B 0.148302f
C27 VP.n1 B 0.039271f
C28 VP.n2 B 0.022108f
C29 VP.t3 B 0.148302f
C30 VP.n3 B 0.02269f
C31 VP.n4 B 0.029146f
C32 VP.t4 B 0.148302f
C33 VP.n5 B 0.039271f
C34 VP.t2 B 0.265678f
C35 VP.n6 B 0.125913f
C36 VP.t1 B 0.148302f
C37 VP.n7 B 0.134131f
C38 VP.n8 B 0.030878f
C39 VP.n9 B 0.163752f
C40 VP.n10 B 0.022108f
C41 VP.n11 B 0.022108f
C42 VP.n12 B 0.02269f
C43 VP.n13 B 0.043312f
C44 VP.n14 B 0.153975f
C45 VP.n15 B 0.789999f
C46 VP.n16 B 0.810867f
C47 VP.t5 B 0.148302f
C48 VP.n17 B 0.153975f
C49 VP.n18 B 0.043312f
C50 VP.n19 B 0.029146f
C51 VP.n20 B 0.022108f
C52 VP.n21 B 0.022108f
C53 VP.n22 B 0.039271f
C54 VP.n23 B 0.030878f
C55 VP.n24 B 0.082891f
C56 VP.n25 B 0.030878f
C57 VP.n26 B 0.022108f
C58 VP.n27 B 0.022108f
C59 VP.n28 B 0.022108f
C60 VP.n29 B 0.02269f
C61 VP.n30 B 0.043312f
C62 VP.n31 B 0.153975f
C63 VP.n32 B 0.023362f
C64 VDD2.t0 B 0.166936f
C65 VDD2.t3 B 0.021287f
C66 VDD2.t1 B 0.021287f
C67 VDD2.n0 B 0.123058f
C68 VDD2.n1 B 1.30461f
C69 VDD2.t5 B 0.164507f
C70 VDD2.n2 B 1.16637f
C71 VDD2.t4 B 0.021287f
C72 VDD2.t2 B 0.021287f
C73 VDD2.n3 B 0.123048f
C74 VTAIL.t6 B 0.028554f
C75 VTAIL.t11 B 0.028554f
C76 VTAIL.n0 B 0.136264f
C77 VTAIL.n1 B 0.308657f
C78 VTAIL.t4 B 0.193124f
C79 VTAIL.n2 B 0.432586f
C80 VTAIL.t3 B 0.028554f
C81 VTAIL.t0 B 0.028554f
C82 VTAIL.n3 B 0.136264f
C83 VTAIL.n4 B 1.00239f
C84 VTAIL.t9 B 0.028554f
C85 VTAIL.t10 B 0.028554f
C86 VTAIL.n5 B 0.136264f
C87 VTAIL.n6 B 1.00238f
C88 VTAIL.t8 B 0.193124f
C89 VTAIL.n7 B 0.432586f
C90 VTAIL.t2 B 0.028554f
C91 VTAIL.t5 B 0.028554f
C92 VTAIL.n8 B 0.136264f
C93 VTAIL.n9 B 0.41157f
C94 VTAIL.t1 B 0.193124f
C95 VTAIL.n10 B 0.880464f
C96 VTAIL.t7 B 0.193124f
C97 VTAIL.n11 B 0.840442f
C98 VN.n0 B 0.028937f
C99 VN.t4 B 0.147238f
C100 VN.n1 B 0.038989f
C101 VN.t5 B 0.263772f
C102 VN.n2 B 0.12501f
C103 VN.t2 B 0.147238f
C104 VN.n3 B 0.133168f
C105 VN.n4 B 0.030656f
C106 VN.n5 B 0.162577f
C107 VN.n6 B 0.02195f
C108 VN.n7 B 0.02195f
C109 VN.n8 B 0.022527f
C110 VN.n9 B 0.043001f
C111 VN.n10 B 0.15287f
C112 VN.n11 B 0.023194f
C113 VN.n12 B 0.028937f
C114 VN.t0 B 0.147238f
C115 VN.n13 B 0.038989f
C116 VN.t3 B 0.263772f
C117 VN.n14 B 0.12501f
C118 VN.t1 B 0.147238f
C119 VN.n15 B 0.133168f
C120 VN.n16 B 0.030656f
C121 VN.n17 B 0.162577f
C122 VN.n18 B 0.02195f
C123 VN.n19 B 0.02195f
C124 VN.n20 B 0.022527f
C125 VN.n21 B 0.043001f
C126 VN.n22 B 0.15287f
C127 VN.n23 B 0.796704f
.ends

