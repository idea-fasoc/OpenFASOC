* NGSPICE file created from diff_pair_sample_0772.ext - technology: sky130A

.subckt diff_pair_sample_0772 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t5 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X1 VDD2.t0 VN.t1 VTAIL.t17 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X2 VTAIL.t16 VN.t2 VDD2.t1 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X3 VDD1.t9 VP.t0 VTAIL.t0 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=4.3836 ps=23.26 w=11.24 l=1.52
X4 VDD1.t8 VP.t1 VTAIL.t2 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=1.8546 ps=11.57 w=11.24 l=1.52
X5 VTAIL.t7 VP.t2 VDD1.t7 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X6 VDD1.t6 VP.t3 VTAIL.t6 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X7 VDD2.t3 VN.t3 VTAIL.t15 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X8 B.t11 B.t9 B.t10 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=0 ps=0 w=11.24 l=1.52
X9 VTAIL.t14 VN.t4 VDD2.t2 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X10 VTAIL.t8 VP.t4 VDD1.t5 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X11 VDD2.t6 VN.t5 VTAIL.t13 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=4.3836 ps=23.26 w=11.24 l=1.52
X12 VTAIL.t5 VP.t5 VDD1.t4 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X13 VDD2.t9 VN.t6 VTAIL.t12 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=1.8546 ps=11.57 w=11.24 l=1.52
X14 VDD2.t8 VN.t7 VTAIL.t11 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=1.8546 ps=11.57 w=11.24 l=1.52
X15 VTAIL.t19 VP.t6 VDD1.t3 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X16 VDD2.t7 VN.t8 VTAIL.t10 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=4.3836 ps=23.26 w=11.24 l=1.52
X17 VDD1.t2 VP.t7 VTAIL.t1 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=1.8546 ps=11.57 w=11.24 l=1.52
X18 VDD1.t1 VP.t8 VTAIL.t3 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=4.3836 ps=23.26 w=11.24 l=1.52
X19 B.t8 B.t6 B.t7 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=0 ps=0 w=11.24 l=1.52
X20 VDD1.t0 VP.t9 VTAIL.t4 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
X21 B.t5 B.t3 B.t4 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=0 ps=0 w=11.24 l=1.52
X22 B.t2 B.t0 B.t1 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=4.3836 pd=23.26 as=0 ps=0 w=11.24 l=1.52
X23 VTAIL.t9 VN.t9 VDD2.t4 w_n3190_n3216# sky130_fd_pr__pfet_01v8 ad=1.8546 pd=11.57 as=1.8546 ps=11.57 w=11.24 l=1.52
R0 VN.n7 VN.t7 211.75
R1 VN.n34 VN.t5 211.75
R2 VN.n12 VN.t1 178.214
R3 VN.n6 VN.t2 178.214
R4 VN.n18 VN.t4 178.214
R5 VN.n25 VN.t8 178.214
R6 VN.n39 VN.t3 178.214
R7 VN.n33 VN.t0 178.214
R8 VN.n45 VN.t9 178.214
R9 VN.n52 VN.t6 178.214
R10 VN.n26 VN.n25 175.906
R11 VN.n53 VN.n52 175.906
R12 VN.n51 VN.n27 161.3
R13 VN.n50 VN.n49 161.3
R14 VN.n48 VN.n28 161.3
R15 VN.n47 VN.n46 161.3
R16 VN.n44 VN.n29 161.3
R17 VN.n43 VN.n42 161.3
R18 VN.n41 VN.n30 161.3
R19 VN.n40 VN.n39 161.3
R20 VN.n38 VN.n31 161.3
R21 VN.n37 VN.n36 161.3
R22 VN.n35 VN.n32 161.3
R23 VN.n24 VN.n0 161.3
R24 VN.n23 VN.n22 161.3
R25 VN.n21 VN.n1 161.3
R26 VN.n20 VN.n19 161.3
R27 VN.n17 VN.n2 161.3
R28 VN.n16 VN.n15 161.3
R29 VN.n14 VN.n3 161.3
R30 VN.n13 VN.n12 161.3
R31 VN.n11 VN.n4 161.3
R32 VN.n10 VN.n9 161.3
R33 VN.n8 VN.n5 161.3
R34 VN.n23 VN.n1 56.4773
R35 VN.n50 VN.n28 56.4773
R36 VN.n7 VN.n6 49.1005
R37 VN.n34 VN.n33 49.1005
R38 VN.n11 VN.n10 47.7136
R39 VN.n16 VN.n3 47.7136
R40 VN.n38 VN.n37 47.7136
R41 VN.n43 VN.n30 47.7136
R42 VN VN.n53 46.9759
R43 VN.n10 VN.n5 33.1076
R44 VN.n17 VN.n16 33.1076
R45 VN.n37 VN.n32 33.1076
R46 VN.n44 VN.n43 33.1076
R47 VN.n12 VN.n11 24.3439
R48 VN.n12 VN.n3 24.3439
R49 VN.n19 VN.n1 24.3439
R50 VN.n24 VN.n23 24.3439
R51 VN.n39 VN.n30 24.3439
R52 VN.n39 VN.n38 24.3439
R53 VN.n46 VN.n28 24.3439
R54 VN.n51 VN.n50 24.3439
R55 VN.n35 VN.n34 17.831
R56 VN.n8 VN.n7 17.831
R57 VN.n6 VN.n5 17.0409
R58 VN.n18 VN.n17 17.0409
R59 VN.n33 VN.n32 17.0409
R60 VN.n45 VN.n44 17.0409
R61 VN.n25 VN.n24 9.73787
R62 VN.n52 VN.n51 9.73787
R63 VN.n19 VN.n18 7.30353
R64 VN.n46 VN.n45 7.30353
R65 VN.n53 VN.n27 0.189894
R66 VN.n49 VN.n27 0.189894
R67 VN.n49 VN.n48 0.189894
R68 VN.n48 VN.n47 0.189894
R69 VN.n47 VN.n29 0.189894
R70 VN.n42 VN.n29 0.189894
R71 VN.n42 VN.n41 0.189894
R72 VN.n41 VN.n40 0.189894
R73 VN.n40 VN.n31 0.189894
R74 VN.n36 VN.n31 0.189894
R75 VN.n36 VN.n35 0.189894
R76 VN.n9 VN.n8 0.189894
R77 VN.n9 VN.n4 0.189894
R78 VN.n13 VN.n4 0.189894
R79 VN.n14 VN.n13 0.189894
R80 VN.n15 VN.n14 0.189894
R81 VN.n15 VN.n2 0.189894
R82 VN.n20 VN.n2 0.189894
R83 VN.n21 VN.n20 0.189894
R84 VN.n22 VN.n21 0.189894
R85 VN.n22 VN.n0 0.189894
R86 VN.n26 VN.n0 0.189894
R87 VN VN.n26 0.0516364
R88 VDD2.n125 VDD2.n124 756.745
R89 VDD2.n60 VDD2.n59 756.745
R90 VDD2.n124 VDD2.n123 585
R91 VDD2.n67 VDD2.n66 585
R92 VDD2.n118 VDD2.n117 585
R93 VDD2.n116 VDD2.n115 585
R94 VDD2.n71 VDD2.n70 585
R95 VDD2.n110 VDD2.n109 585
R96 VDD2.n108 VDD2.n107 585
R97 VDD2.n75 VDD2.n74 585
R98 VDD2.n102 VDD2.n101 585
R99 VDD2.n100 VDD2.n99 585
R100 VDD2.n79 VDD2.n78 585
R101 VDD2.n94 VDD2.n93 585
R102 VDD2.n92 VDD2.n91 585
R103 VDD2.n83 VDD2.n82 585
R104 VDD2.n86 VDD2.n85 585
R105 VDD2.n21 VDD2.n20 585
R106 VDD2.n18 VDD2.n17 585
R107 VDD2.n27 VDD2.n26 585
R108 VDD2.n29 VDD2.n28 585
R109 VDD2.n14 VDD2.n13 585
R110 VDD2.n35 VDD2.n34 585
R111 VDD2.n37 VDD2.n36 585
R112 VDD2.n10 VDD2.n9 585
R113 VDD2.n43 VDD2.n42 585
R114 VDD2.n45 VDD2.n44 585
R115 VDD2.n6 VDD2.n5 585
R116 VDD2.n51 VDD2.n50 585
R117 VDD2.n53 VDD2.n52 585
R118 VDD2.n2 VDD2.n1 585
R119 VDD2.n59 VDD2.n58 585
R120 VDD2.t9 VDD2.n84 327.466
R121 VDD2.t8 VDD2.n19 327.466
R122 VDD2.n124 VDD2.n66 171.744
R123 VDD2.n117 VDD2.n66 171.744
R124 VDD2.n117 VDD2.n116 171.744
R125 VDD2.n116 VDD2.n70 171.744
R126 VDD2.n109 VDD2.n70 171.744
R127 VDD2.n109 VDD2.n108 171.744
R128 VDD2.n108 VDD2.n74 171.744
R129 VDD2.n101 VDD2.n74 171.744
R130 VDD2.n101 VDD2.n100 171.744
R131 VDD2.n100 VDD2.n78 171.744
R132 VDD2.n93 VDD2.n78 171.744
R133 VDD2.n93 VDD2.n92 171.744
R134 VDD2.n92 VDD2.n82 171.744
R135 VDD2.n85 VDD2.n82 171.744
R136 VDD2.n20 VDD2.n17 171.744
R137 VDD2.n27 VDD2.n17 171.744
R138 VDD2.n28 VDD2.n27 171.744
R139 VDD2.n28 VDD2.n13 171.744
R140 VDD2.n35 VDD2.n13 171.744
R141 VDD2.n36 VDD2.n35 171.744
R142 VDD2.n36 VDD2.n9 171.744
R143 VDD2.n43 VDD2.n9 171.744
R144 VDD2.n44 VDD2.n43 171.744
R145 VDD2.n44 VDD2.n5 171.744
R146 VDD2.n51 VDD2.n5 171.744
R147 VDD2.n52 VDD2.n51 171.744
R148 VDD2.n52 VDD2.n1 171.744
R149 VDD2.n59 VDD2.n1 171.744
R150 VDD2.n85 VDD2.t9 85.8723
R151 VDD2.n20 VDD2.t8 85.8723
R152 VDD2.n64 VDD2.n63 79.3036
R153 VDD2 VDD2.n129 79.2998
R154 VDD2.n128 VDD2.n127 78.163
R155 VDD2.n62 VDD2.n61 78.1628
R156 VDD2.n62 VDD2.n60 52.3984
R157 VDD2.n126 VDD2.n125 50.8035
R158 VDD2.n126 VDD2.n64 40.9804
R159 VDD2.n86 VDD2.n84 16.3895
R160 VDD2.n21 VDD2.n19 16.3895
R161 VDD2.n87 VDD2.n83 12.8005
R162 VDD2.n22 VDD2.n18 12.8005
R163 VDD2.n91 VDD2.n90 12.0247
R164 VDD2.n26 VDD2.n25 12.0247
R165 VDD2.n123 VDD2.n65 11.249
R166 VDD2.n94 VDD2.n81 11.249
R167 VDD2.n29 VDD2.n16 11.249
R168 VDD2.n58 VDD2.n0 11.249
R169 VDD2.n122 VDD2.n67 10.4732
R170 VDD2.n95 VDD2.n79 10.4732
R171 VDD2.n30 VDD2.n14 10.4732
R172 VDD2.n57 VDD2.n2 10.4732
R173 VDD2.n119 VDD2.n118 9.69747
R174 VDD2.n99 VDD2.n98 9.69747
R175 VDD2.n34 VDD2.n33 9.69747
R176 VDD2.n54 VDD2.n53 9.69747
R177 VDD2.n121 VDD2.n65 9.45567
R178 VDD2.n56 VDD2.n0 9.45567
R179 VDD2.n112 VDD2.n111 9.3005
R180 VDD2.n114 VDD2.n113 9.3005
R181 VDD2.n69 VDD2.n68 9.3005
R182 VDD2.n120 VDD2.n119 9.3005
R183 VDD2.n122 VDD2.n121 9.3005
R184 VDD2.n73 VDD2.n72 9.3005
R185 VDD2.n106 VDD2.n105 9.3005
R186 VDD2.n104 VDD2.n103 9.3005
R187 VDD2.n77 VDD2.n76 9.3005
R188 VDD2.n98 VDD2.n97 9.3005
R189 VDD2.n96 VDD2.n95 9.3005
R190 VDD2.n81 VDD2.n80 9.3005
R191 VDD2.n90 VDD2.n89 9.3005
R192 VDD2.n88 VDD2.n87 9.3005
R193 VDD2.n8 VDD2.n7 9.3005
R194 VDD2.n47 VDD2.n46 9.3005
R195 VDD2.n49 VDD2.n48 9.3005
R196 VDD2.n4 VDD2.n3 9.3005
R197 VDD2.n55 VDD2.n54 9.3005
R198 VDD2.n57 VDD2.n56 9.3005
R199 VDD2.n39 VDD2.n38 9.3005
R200 VDD2.n12 VDD2.n11 9.3005
R201 VDD2.n33 VDD2.n32 9.3005
R202 VDD2.n31 VDD2.n30 9.3005
R203 VDD2.n16 VDD2.n15 9.3005
R204 VDD2.n25 VDD2.n24 9.3005
R205 VDD2.n23 VDD2.n22 9.3005
R206 VDD2.n41 VDD2.n40 9.3005
R207 VDD2.n115 VDD2.n69 8.92171
R208 VDD2.n102 VDD2.n77 8.92171
R209 VDD2.n37 VDD2.n12 8.92171
R210 VDD2.n50 VDD2.n4 8.92171
R211 VDD2.n114 VDD2.n71 8.14595
R212 VDD2.n103 VDD2.n75 8.14595
R213 VDD2.n38 VDD2.n10 8.14595
R214 VDD2.n49 VDD2.n6 8.14595
R215 VDD2.n111 VDD2.n110 7.3702
R216 VDD2.n107 VDD2.n106 7.3702
R217 VDD2.n42 VDD2.n41 7.3702
R218 VDD2.n46 VDD2.n45 7.3702
R219 VDD2.n110 VDD2.n73 6.59444
R220 VDD2.n107 VDD2.n73 6.59444
R221 VDD2.n42 VDD2.n8 6.59444
R222 VDD2.n45 VDD2.n8 6.59444
R223 VDD2.n111 VDD2.n71 5.81868
R224 VDD2.n106 VDD2.n75 5.81868
R225 VDD2.n41 VDD2.n10 5.81868
R226 VDD2.n46 VDD2.n6 5.81868
R227 VDD2.n115 VDD2.n114 5.04292
R228 VDD2.n103 VDD2.n102 5.04292
R229 VDD2.n38 VDD2.n37 5.04292
R230 VDD2.n50 VDD2.n49 5.04292
R231 VDD2.n118 VDD2.n69 4.26717
R232 VDD2.n99 VDD2.n77 4.26717
R233 VDD2.n34 VDD2.n12 4.26717
R234 VDD2.n53 VDD2.n4 4.26717
R235 VDD2.n88 VDD2.n84 3.70982
R236 VDD2.n23 VDD2.n19 3.70982
R237 VDD2.n119 VDD2.n67 3.49141
R238 VDD2.n98 VDD2.n79 3.49141
R239 VDD2.n33 VDD2.n14 3.49141
R240 VDD2.n54 VDD2.n2 3.49141
R241 VDD2.n129 VDD2.t5 2.8924
R242 VDD2.n129 VDD2.t6 2.8924
R243 VDD2.n127 VDD2.t4 2.8924
R244 VDD2.n127 VDD2.t3 2.8924
R245 VDD2.n63 VDD2.t2 2.8924
R246 VDD2.n63 VDD2.t7 2.8924
R247 VDD2.n61 VDD2.t1 2.8924
R248 VDD2.n61 VDD2.t0 2.8924
R249 VDD2.n123 VDD2.n122 2.71565
R250 VDD2.n95 VDD2.n94 2.71565
R251 VDD2.n30 VDD2.n29 2.71565
R252 VDD2.n58 VDD2.n57 2.71565
R253 VDD2.n125 VDD2.n65 1.93989
R254 VDD2.n91 VDD2.n81 1.93989
R255 VDD2.n26 VDD2.n16 1.93989
R256 VDD2.n60 VDD2.n0 1.93989
R257 VDD2.n128 VDD2.n126 1.59533
R258 VDD2.n90 VDD2.n83 1.16414
R259 VDD2.n25 VDD2.n18 1.16414
R260 VDD2 VDD2.n128 0.457397
R261 VDD2.n87 VDD2.n86 0.388379
R262 VDD2.n22 VDD2.n21 0.388379
R263 VDD2.n64 VDD2.n62 0.343861
R264 VDD2.n121 VDD2.n120 0.155672
R265 VDD2.n120 VDD2.n68 0.155672
R266 VDD2.n113 VDD2.n68 0.155672
R267 VDD2.n113 VDD2.n112 0.155672
R268 VDD2.n112 VDD2.n72 0.155672
R269 VDD2.n105 VDD2.n72 0.155672
R270 VDD2.n105 VDD2.n104 0.155672
R271 VDD2.n104 VDD2.n76 0.155672
R272 VDD2.n97 VDD2.n76 0.155672
R273 VDD2.n97 VDD2.n96 0.155672
R274 VDD2.n96 VDD2.n80 0.155672
R275 VDD2.n89 VDD2.n80 0.155672
R276 VDD2.n89 VDD2.n88 0.155672
R277 VDD2.n24 VDD2.n23 0.155672
R278 VDD2.n24 VDD2.n15 0.155672
R279 VDD2.n31 VDD2.n15 0.155672
R280 VDD2.n32 VDD2.n31 0.155672
R281 VDD2.n32 VDD2.n11 0.155672
R282 VDD2.n39 VDD2.n11 0.155672
R283 VDD2.n40 VDD2.n39 0.155672
R284 VDD2.n40 VDD2.n7 0.155672
R285 VDD2.n47 VDD2.n7 0.155672
R286 VDD2.n48 VDD2.n47 0.155672
R287 VDD2.n48 VDD2.n3 0.155672
R288 VDD2.n55 VDD2.n3 0.155672
R289 VDD2.n56 VDD2.n55 0.155672
R290 VTAIL.n260 VTAIL.n259 756.745
R291 VTAIL.n62 VTAIL.n61 756.745
R292 VTAIL.n198 VTAIL.n197 756.745
R293 VTAIL.n132 VTAIL.n131 756.745
R294 VTAIL.n221 VTAIL.n220 585
R295 VTAIL.n218 VTAIL.n217 585
R296 VTAIL.n227 VTAIL.n226 585
R297 VTAIL.n229 VTAIL.n228 585
R298 VTAIL.n214 VTAIL.n213 585
R299 VTAIL.n235 VTAIL.n234 585
R300 VTAIL.n237 VTAIL.n236 585
R301 VTAIL.n210 VTAIL.n209 585
R302 VTAIL.n243 VTAIL.n242 585
R303 VTAIL.n245 VTAIL.n244 585
R304 VTAIL.n206 VTAIL.n205 585
R305 VTAIL.n251 VTAIL.n250 585
R306 VTAIL.n253 VTAIL.n252 585
R307 VTAIL.n202 VTAIL.n201 585
R308 VTAIL.n259 VTAIL.n258 585
R309 VTAIL.n23 VTAIL.n22 585
R310 VTAIL.n20 VTAIL.n19 585
R311 VTAIL.n29 VTAIL.n28 585
R312 VTAIL.n31 VTAIL.n30 585
R313 VTAIL.n16 VTAIL.n15 585
R314 VTAIL.n37 VTAIL.n36 585
R315 VTAIL.n39 VTAIL.n38 585
R316 VTAIL.n12 VTAIL.n11 585
R317 VTAIL.n45 VTAIL.n44 585
R318 VTAIL.n47 VTAIL.n46 585
R319 VTAIL.n8 VTAIL.n7 585
R320 VTAIL.n53 VTAIL.n52 585
R321 VTAIL.n55 VTAIL.n54 585
R322 VTAIL.n4 VTAIL.n3 585
R323 VTAIL.n61 VTAIL.n60 585
R324 VTAIL.n197 VTAIL.n196 585
R325 VTAIL.n140 VTAIL.n139 585
R326 VTAIL.n191 VTAIL.n190 585
R327 VTAIL.n189 VTAIL.n188 585
R328 VTAIL.n144 VTAIL.n143 585
R329 VTAIL.n183 VTAIL.n182 585
R330 VTAIL.n181 VTAIL.n180 585
R331 VTAIL.n148 VTAIL.n147 585
R332 VTAIL.n175 VTAIL.n174 585
R333 VTAIL.n173 VTAIL.n172 585
R334 VTAIL.n152 VTAIL.n151 585
R335 VTAIL.n167 VTAIL.n166 585
R336 VTAIL.n165 VTAIL.n164 585
R337 VTAIL.n156 VTAIL.n155 585
R338 VTAIL.n159 VTAIL.n158 585
R339 VTAIL.n131 VTAIL.n130 585
R340 VTAIL.n74 VTAIL.n73 585
R341 VTAIL.n125 VTAIL.n124 585
R342 VTAIL.n123 VTAIL.n122 585
R343 VTAIL.n78 VTAIL.n77 585
R344 VTAIL.n117 VTAIL.n116 585
R345 VTAIL.n115 VTAIL.n114 585
R346 VTAIL.n82 VTAIL.n81 585
R347 VTAIL.n109 VTAIL.n108 585
R348 VTAIL.n107 VTAIL.n106 585
R349 VTAIL.n86 VTAIL.n85 585
R350 VTAIL.n101 VTAIL.n100 585
R351 VTAIL.n99 VTAIL.n98 585
R352 VTAIL.n90 VTAIL.n89 585
R353 VTAIL.n93 VTAIL.n92 585
R354 VTAIL.t10 VTAIL.n219 327.466
R355 VTAIL.t3 VTAIL.n21 327.466
R356 VTAIL.t0 VTAIL.n157 327.466
R357 VTAIL.t13 VTAIL.n91 327.466
R358 VTAIL.n220 VTAIL.n217 171.744
R359 VTAIL.n227 VTAIL.n217 171.744
R360 VTAIL.n228 VTAIL.n227 171.744
R361 VTAIL.n228 VTAIL.n213 171.744
R362 VTAIL.n235 VTAIL.n213 171.744
R363 VTAIL.n236 VTAIL.n235 171.744
R364 VTAIL.n236 VTAIL.n209 171.744
R365 VTAIL.n243 VTAIL.n209 171.744
R366 VTAIL.n244 VTAIL.n243 171.744
R367 VTAIL.n244 VTAIL.n205 171.744
R368 VTAIL.n251 VTAIL.n205 171.744
R369 VTAIL.n252 VTAIL.n251 171.744
R370 VTAIL.n252 VTAIL.n201 171.744
R371 VTAIL.n259 VTAIL.n201 171.744
R372 VTAIL.n22 VTAIL.n19 171.744
R373 VTAIL.n29 VTAIL.n19 171.744
R374 VTAIL.n30 VTAIL.n29 171.744
R375 VTAIL.n30 VTAIL.n15 171.744
R376 VTAIL.n37 VTAIL.n15 171.744
R377 VTAIL.n38 VTAIL.n37 171.744
R378 VTAIL.n38 VTAIL.n11 171.744
R379 VTAIL.n45 VTAIL.n11 171.744
R380 VTAIL.n46 VTAIL.n45 171.744
R381 VTAIL.n46 VTAIL.n7 171.744
R382 VTAIL.n53 VTAIL.n7 171.744
R383 VTAIL.n54 VTAIL.n53 171.744
R384 VTAIL.n54 VTAIL.n3 171.744
R385 VTAIL.n61 VTAIL.n3 171.744
R386 VTAIL.n197 VTAIL.n139 171.744
R387 VTAIL.n190 VTAIL.n139 171.744
R388 VTAIL.n190 VTAIL.n189 171.744
R389 VTAIL.n189 VTAIL.n143 171.744
R390 VTAIL.n182 VTAIL.n143 171.744
R391 VTAIL.n182 VTAIL.n181 171.744
R392 VTAIL.n181 VTAIL.n147 171.744
R393 VTAIL.n174 VTAIL.n147 171.744
R394 VTAIL.n174 VTAIL.n173 171.744
R395 VTAIL.n173 VTAIL.n151 171.744
R396 VTAIL.n166 VTAIL.n151 171.744
R397 VTAIL.n166 VTAIL.n165 171.744
R398 VTAIL.n165 VTAIL.n155 171.744
R399 VTAIL.n158 VTAIL.n155 171.744
R400 VTAIL.n131 VTAIL.n73 171.744
R401 VTAIL.n124 VTAIL.n73 171.744
R402 VTAIL.n124 VTAIL.n123 171.744
R403 VTAIL.n123 VTAIL.n77 171.744
R404 VTAIL.n116 VTAIL.n77 171.744
R405 VTAIL.n116 VTAIL.n115 171.744
R406 VTAIL.n115 VTAIL.n81 171.744
R407 VTAIL.n108 VTAIL.n81 171.744
R408 VTAIL.n108 VTAIL.n107 171.744
R409 VTAIL.n107 VTAIL.n85 171.744
R410 VTAIL.n100 VTAIL.n85 171.744
R411 VTAIL.n100 VTAIL.n99 171.744
R412 VTAIL.n99 VTAIL.n89 171.744
R413 VTAIL.n92 VTAIL.n89 171.744
R414 VTAIL.n220 VTAIL.t10 85.8723
R415 VTAIL.n22 VTAIL.t3 85.8723
R416 VTAIL.n158 VTAIL.t0 85.8723
R417 VTAIL.n92 VTAIL.t13 85.8723
R418 VTAIL.n137 VTAIL.n136 61.4842
R419 VTAIL.n135 VTAIL.n134 61.4842
R420 VTAIL.n71 VTAIL.n70 61.4842
R421 VTAIL.n69 VTAIL.n68 61.4842
R422 VTAIL.n263 VTAIL.n262 61.484
R423 VTAIL.n1 VTAIL.n0 61.484
R424 VTAIL.n65 VTAIL.n64 61.484
R425 VTAIL.n67 VTAIL.n66 61.484
R426 VTAIL.n261 VTAIL.n260 34.1247
R427 VTAIL.n63 VTAIL.n62 34.1247
R428 VTAIL.n199 VTAIL.n198 34.1247
R429 VTAIL.n133 VTAIL.n132 34.1247
R430 VTAIL.n69 VTAIL.n67 25.2462
R431 VTAIL.n261 VTAIL.n199 23.6514
R432 VTAIL.n221 VTAIL.n219 16.3895
R433 VTAIL.n23 VTAIL.n21 16.3895
R434 VTAIL.n159 VTAIL.n157 16.3895
R435 VTAIL.n93 VTAIL.n91 16.3895
R436 VTAIL.n222 VTAIL.n218 12.8005
R437 VTAIL.n24 VTAIL.n20 12.8005
R438 VTAIL.n160 VTAIL.n156 12.8005
R439 VTAIL.n94 VTAIL.n90 12.8005
R440 VTAIL.n226 VTAIL.n225 12.0247
R441 VTAIL.n28 VTAIL.n27 12.0247
R442 VTAIL.n164 VTAIL.n163 12.0247
R443 VTAIL.n98 VTAIL.n97 12.0247
R444 VTAIL.n229 VTAIL.n216 11.249
R445 VTAIL.n258 VTAIL.n200 11.249
R446 VTAIL.n31 VTAIL.n18 11.249
R447 VTAIL.n60 VTAIL.n2 11.249
R448 VTAIL.n196 VTAIL.n138 11.249
R449 VTAIL.n167 VTAIL.n154 11.249
R450 VTAIL.n130 VTAIL.n72 11.249
R451 VTAIL.n101 VTAIL.n88 11.249
R452 VTAIL.n230 VTAIL.n214 10.4732
R453 VTAIL.n257 VTAIL.n202 10.4732
R454 VTAIL.n32 VTAIL.n16 10.4732
R455 VTAIL.n59 VTAIL.n4 10.4732
R456 VTAIL.n195 VTAIL.n140 10.4732
R457 VTAIL.n168 VTAIL.n152 10.4732
R458 VTAIL.n129 VTAIL.n74 10.4732
R459 VTAIL.n102 VTAIL.n86 10.4732
R460 VTAIL.n234 VTAIL.n233 9.69747
R461 VTAIL.n254 VTAIL.n253 9.69747
R462 VTAIL.n36 VTAIL.n35 9.69747
R463 VTAIL.n56 VTAIL.n55 9.69747
R464 VTAIL.n192 VTAIL.n191 9.69747
R465 VTAIL.n172 VTAIL.n171 9.69747
R466 VTAIL.n126 VTAIL.n125 9.69747
R467 VTAIL.n106 VTAIL.n105 9.69747
R468 VTAIL.n256 VTAIL.n200 9.45567
R469 VTAIL.n58 VTAIL.n2 9.45567
R470 VTAIL.n194 VTAIL.n138 9.45567
R471 VTAIL.n128 VTAIL.n72 9.45567
R472 VTAIL.n208 VTAIL.n207 9.3005
R473 VTAIL.n247 VTAIL.n246 9.3005
R474 VTAIL.n249 VTAIL.n248 9.3005
R475 VTAIL.n204 VTAIL.n203 9.3005
R476 VTAIL.n255 VTAIL.n254 9.3005
R477 VTAIL.n257 VTAIL.n256 9.3005
R478 VTAIL.n239 VTAIL.n238 9.3005
R479 VTAIL.n212 VTAIL.n211 9.3005
R480 VTAIL.n233 VTAIL.n232 9.3005
R481 VTAIL.n231 VTAIL.n230 9.3005
R482 VTAIL.n216 VTAIL.n215 9.3005
R483 VTAIL.n225 VTAIL.n224 9.3005
R484 VTAIL.n223 VTAIL.n222 9.3005
R485 VTAIL.n241 VTAIL.n240 9.3005
R486 VTAIL.n10 VTAIL.n9 9.3005
R487 VTAIL.n49 VTAIL.n48 9.3005
R488 VTAIL.n51 VTAIL.n50 9.3005
R489 VTAIL.n6 VTAIL.n5 9.3005
R490 VTAIL.n57 VTAIL.n56 9.3005
R491 VTAIL.n59 VTAIL.n58 9.3005
R492 VTAIL.n41 VTAIL.n40 9.3005
R493 VTAIL.n14 VTAIL.n13 9.3005
R494 VTAIL.n35 VTAIL.n34 9.3005
R495 VTAIL.n33 VTAIL.n32 9.3005
R496 VTAIL.n18 VTAIL.n17 9.3005
R497 VTAIL.n27 VTAIL.n26 9.3005
R498 VTAIL.n25 VTAIL.n24 9.3005
R499 VTAIL.n43 VTAIL.n42 9.3005
R500 VTAIL.n195 VTAIL.n194 9.3005
R501 VTAIL.n193 VTAIL.n192 9.3005
R502 VTAIL.n142 VTAIL.n141 9.3005
R503 VTAIL.n187 VTAIL.n186 9.3005
R504 VTAIL.n185 VTAIL.n184 9.3005
R505 VTAIL.n146 VTAIL.n145 9.3005
R506 VTAIL.n179 VTAIL.n178 9.3005
R507 VTAIL.n177 VTAIL.n176 9.3005
R508 VTAIL.n150 VTAIL.n149 9.3005
R509 VTAIL.n171 VTAIL.n170 9.3005
R510 VTAIL.n169 VTAIL.n168 9.3005
R511 VTAIL.n154 VTAIL.n153 9.3005
R512 VTAIL.n163 VTAIL.n162 9.3005
R513 VTAIL.n161 VTAIL.n160 9.3005
R514 VTAIL.n119 VTAIL.n118 9.3005
R515 VTAIL.n121 VTAIL.n120 9.3005
R516 VTAIL.n76 VTAIL.n75 9.3005
R517 VTAIL.n127 VTAIL.n126 9.3005
R518 VTAIL.n129 VTAIL.n128 9.3005
R519 VTAIL.n80 VTAIL.n79 9.3005
R520 VTAIL.n113 VTAIL.n112 9.3005
R521 VTAIL.n111 VTAIL.n110 9.3005
R522 VTAIL.n84 VTAIL.n83 9.3005
R523 VTAIL.n105 VTAIL.n104 9.3005
R524 VTAIL.n103 VTAIL.n102 9.3005
R525 VTAIL.n88 VTAIL.n87 9.3005
R526 VTAIL.n97 VTAIL.n96 9.3005
R527 VTAIL.n95 VTAIL.n94 9.3005
R528 VTAIL.n237 VTAIL.n212 8.92171
R529 VTAIL.n250 VTAIL.n204 8.92171
R530 VTAIL.n39 VTAIL.n14 8.92171
R531 VTAIL.n52 VTAIL.n6 8.92171
R532 VTAIL.n188 VTAIL.n142 8.92171
R533 VTAIL.n175 VTAIL.n150 8.92171
R534 VTAIL.n122 VTAIL.n76 8.92171
R535 VTAIL.n109 VTAIL.n84 8.92171
R536 VTAIL.n238 VTAIL.n210 8.14595
R537 VTAIL.n249 VTAIL.n206 8.14595
R538 VTAIL.n40 VTAIL.n12 8.14595
R539 VTAIL.n51 VTAIL.n8 8.14595
R540 VTAIL.n187 VTAIL.n144 8.14595
R541 VTAIL.n176 VTAIL.n148 8.14595
R542 VTAIL.n121 VTAIL.n78 8.14595
R543 VTAIL.n110 VTAIL.n82 8.14595
R544 VTAIL.n242 VTAIL.n241 7.3702
R545 VTAIL.n246 VTAIL.n245 7.3702
R546 VTAIL.n44 VTAIL.n43 7.3702
R547 VTAIL.n48 VTAIL.n47 7.3702
R548 VTAIL.n184 VTAIL.n183 7.3702
R549 VTAIL.n180 VTAIL.n179 7.3702
R550 VTAIL.n118 VTAIL.n117 7.3702
R551 VTAIL.n114 VTAIL.n113 7.3702
R552 VTAIL.n242 VTAIL.n208 6.59444
R553 VTAIL.n245 VTAIL.n208 6.59444
R554 VTAIL.n44 VTAIL.n10 6.59444
R555 VTAIL.n47 VTAIL.n10 6.59444
R556 VTAIL.n183 VTAIL.n146 6.59444
R557 VTAIL.n180 VTAIL.n146 6.59444
R558 VTAIL.n117 VTAIL.n80 6.59444
R559 VTAIL.n114 VTAIL.n80 6.59444
R560 VTAIL.n241 VTAIL.n210 5.81868
R561 VTAIL.n246 VTAIL.n206 5.81868
R562 VTAIL.n43 VTAIL.n12 5.81868
R563 VTAIL.n48 VTAIL.n8 5.81868
R564 VTAIL.n184 VTAIL.n144 5.81868
R565 VTAIL.n179 VTAIL.n148 5.81868
R566 VTAIL.n118 VTAIL.n78 5.81868
R567 VTAIL.n113 VTAIL.n82 5.81868
R568 VTAIL.n238 VTAIL.n237 5.04292
R569 VTAIL.n250 VTAIL.n249 5.04292
R570 VTAIL.n40 VTAIL.n39 5.04292
R571 VTAIL.n52 VTAIL.n51 5.04292
R572 VTAIL.n188 VTAIL.n187 5.04292
R573 VTAIL.n176 VTAIL.n175 5.04292
R574 VTAIL.n122 VTAIL.n121 5.04292
R575 VTAIL.n110 VTAIL.n109 5.04292
R576 VTAIL.n234 VTAIL.n212 4.26717
R577 VTAIL.n253 VTAIL.n204 4.26717
R578 VTAIL.n36 VTAIL.n14 4.26717
R579 VTAIL.n55 VTAIL.n6 4.26717
R580 VTAIL.n191 VTAIL.n142 4.26717
R581 VTAIL.n172 VTAIL.n150 4.26717
R582 VTAIL.n125 VTAIL.n76 4.26717
R583 VTAIL.n106 VTAIL.n84 4.26717
R584 VTAIL.n223 VTAIL.n219 3.70982
R585 VTAIL.n25 VTAIL.n21 3.70982
R586 VTAIL.n161 VTAIL.n157 3.70982
R587 VTAIL.n95 VTAIL.n91 3.70982
R588 VTAIL.n233 VTAIL.n214 3.49141
R589 VTAIL.n254 VTAIL.n202 3.49141
R590 VTAIL.n35 VTAIL.n16 3.49141
R591 VTAIL.n56 VTAIL.n4 3.49141
R592 VTAIL.n192 VTAIL.n140 3.49141
R593 VTAIL.n171 VTAIL.n152 3.49141
R594 VTAIL.n126 VTAIL.n74 3.49141
R595 VTAIL.n105 VTAIL.n86 3.49141
R596 VTAIL.n262 VTAIL.t17 2.8924
R597 VTAIL.n262 VTAIL.t14 2.8924
R598 VTAIL.n0 VTAIL.t11 2.8924
R599 VTAIL.n0 VTAIL.t16 2.8924
R600 VTAIL.n64 VTAIL.t6 2.8924
R601 VTAIL.n64 VTAIL.t7 2.8924
R602 VTAIL.n66 VTAIL.t1 2.8924
R603 VTAIL.n66 VTAIL.t8 2.8924
R604 VTAIL.n136 VTAIL.t4 2.8924
R605 VTAIL.n136 VTAIL.t5 2.8924
R606 VTAIL.n134 VTAIL.t2 2.8924
R607 VTAIL.n134 VTAIL.t19 2.8924
R608 VTAIL.n70 VTAIL.t15 2.8924
R609 VTAIL.n70 VTAIL.t18 2.8924
R610 VTAIL.n68 VTAIL.t12 2.8924
R611 VTAIL.n68 VTAIL.t9 2.8924
R612 VTAIL.n230 VTAIL.n229 2.71565
R613 VTAIL.n258 VTAIL.n257 2.71565
R614 VTAIL.n32 VTAIL.n31 2.71565
R615 VTAIL.n60 VTAIL.n59 2.71565
R616 VTAIL.n196 VTAIL.n195 2.71565
R617 VTAIL.n168 VTAIL.n167 2.71565
R618 VTAIL.n130 VTAIL.n129 2.71565
R619 VTAIL.n102 VTAIL.n101 2.71565
R620 VTAIL.n226 VTAIL.n216 1.93989
R621 VTAIL.n260 VTAIL.n200 1.93989
R622 VTAIL.n28 VTAIL.n18 1.93989
R623 VTAIL.n62 VTAIL.n2 1.93989
R624 VTAIL.n198 VTAIL.n138 1.93989
R625 VTAIL.n164 VTAIL.n154 1.93989
R626 VTAIL.n132 VTAIL.n72 1.93989
R627 VTAIL.n98 VTAIL.n88 1.93989
R628 VTAIL.n71 VTAIL.n69 1.59533
R629 VTAIL.n133 VTAIL.n71 1.59533
R630 VTAIL.n137 VTAIL.n135 1.59533
R631 VTAIL.n199 VTAIL.n137 1.59533
R632 VTAIL.n67 VTAIL.n65 1.59533
R633 VTAIL.n65 VTAIL.n63 1.59533
R634 VTAIL.n263 VTAIL.n261 1.59533
R635 VTAIL.n135 VTAIL.n133 1.26774
R636 VTAIL.n63 VTAIL.n1 1.26774
R637 VTAIL VTAIL.n1 1.25481
R638 VTAIL.n225 VTAIL.n218 1.16414
R639 VTAIL.n27 VTAIL.n20 1.16414
R640 VTAIL.n163 VTAIL.n156 1.16414
R641 VTAIL.n97 VTAIL.n90 1.16414
R642 VTAIL.n222 VTAIL.n221 0.388379
R643 VTAIL.n24 VTAIL.n23 0.388379
R644 VTAIL.n160 VTAIL.n159 0.388379
R645 VTAIL.n94 VTAIL.n93 0.388379
R646 VTAIL VTAIL.n263 0.341017
R647 VTAIL.n224 VTAIL.n223 0.155672
R648 VTAIL.n224 VTAIL.n215 0.155672
R649 VTAIL.n231 VTAIL.n215 0.155672
R650 VTAIL.n232 VTAIL.n231 0.155672
R651 VTAIL.n232 VTAIL.n211 0.155672
R652 VTAIL.n239 VTAIL.n211 0.155672
R653 VTAIL.n240 VTAIL.n239 0.155672
R654 VTAIL.n240 VTAIL.n207 0.155672
R655 VTAIL.n247 VTAIL.n207 0.155672
R656 VTAIL.n248 VTAIL.n247 0.155672
R657 VTAIL.n248 VTAIL.n203 0.155672
R658 VTAIL.n255 VTAIL.n203 0.155672
R659 VTAIL.n256 VTAIL.n255 0.155672
R660 VTAIL.n26 VTAIL.n25 0.155672
R661 VTAIL.n26 VTAIL.n17 0.155672
R662 VTAIL.n33 VTAIL.n17 0.155672
R663 VTAIL.n34 VTAIL.n33 0.155672
R664 VTAIL.n34 VTAIL.n13 0.155672
R665 VTAIL.n41 VTAIL.n13 0.155672
R666 VTAIL.n42 VTAIL.n41 0.155672
R667 VTAIL.n42 VTAIL.n9 0.155672
R668 VTAIL.n49 VTAIL.n9 0.155672
R669 VTAIL.n50 VTAIL.n49 0.155672
R670 VTAIL.n50 VTAIL.n5 0.155672
R671 VTAIL.n57 VTAIL.n5 0.155672
R672 VTAIL.n58 VTAIL.n57 0.155672
R673 VTAIL.n194 VTAIL.n193 0.155672
R674 VTAIL.n193 VTAIL.n141 0.155672
R675 VTAIL.n186 VTAIL.n141 0.155672
R676 VTAIL.n186 VTAIL.n185 0.155672
R677 VTAIL.n185 VTAIL.n145 0.155672
R678 VTAIL.n178 VTAIL.n145 0.155672
R679 VTAIL.n178 VTAIL.n177 0.155672
R680 VTAIL.n177 VTAIL.n149 0.155672
R681 VTAIL.n170 VTAIL.n149 0.155672
R682 VTAIL.n170 VTAIL.n169 0.155672
R683 VTAIL.n169 VTAIL.n153 0.155672
R684 VTAIL.n162 VTAIL.n153 0.155672
R685 VTAIL.n162 VTAIL.n161 0.155672
R686 VTAIL.n128 VTAIL.n127 0.155672
R687 VTAIL.n127 VTAIL.n75 0.155672
R688 VTAIL.n120 VTAIL.n75 0.155672
R689 VTAIL.n120 VTAIL.n119 0.155672
R690 VTAIL.n119 VTAIL.n79 0.155672
R691 VTAIL.n112 VTAIL.n79 0.155672
R692 VTAIL.n112 VTAIL.n111 0.155672
R693 VTAIL.n111 VTAIL.n83 0.155672
R694 VTAIL.n104 VTAIL.n83 0.155672
R695 VTAIL.n104 VTAIL.n103 0.155672
R696 VTAIL.n103 VTAIL.n87 0.155672
R697 VTAIL.n96 VTAIL.n87 0.155672
R698 VTAIL.n96 VTAIL.n95 0.155672
R699 VP.n15 VP.t1 211.75
R700 VP.n48 VP.t3 178.214
R701 VP.n35 VP.t7 178.214
R702 VP.n41 VP.t4 178.214
R703 VP.n54 VP.t2 178.214
R704 VP.n61 VP.t8 178.214
R705 VP.n20 VP.t9 178.214
R706 VP.n33 VP.t0 178.214
R707 VP.n26 VP.t5 178.214
R708 VP.n14 VP.t6 178.214
R709 VP.n36 VP.n35 175.906
R710 VP.n62 VP.n61 175.906
R711 VP.n34 VP.n33 175.906
R712 VP.n16 VP.n13 161.3
R713 VP.n18 VP.n17 161.3
R714 VP.n19 VP.n12 161.3
R715 VP.n21 VP.n20 161.3
R716 VP.n22 VP.n11 161.3
R717 VP.n24 VP.n23 161.3
R718 VP.n25 VP.n10 161.3
R719 VP.n28 VP.n27 161.3
R720 VP.n29 VP.n9 161.3
R721 VP.n31 VP.n30 161.3
R722 VP.n32 VP.n8 161.3
R723 VP.n60 VP.n0 161.3
R724 VP.n59 VP.n58 161.3
R725 VP.n57 VP.n1 161.3
R726 VP.n56 VP.n55 161.3
R727 VP.n53 VP.n2 161.3
R728 VP.n52 VP.n51 161.3
R729 VP.n50 VP.n3 161.3
R730 VP.n49 VP.n48 161.3
R731 VP.n47 VP.n4 161.3
R732 VP.n46 VP.n45 161.3
R733 VP.n44 VP.n5 161.3
R734 VP.n43 VP.n42 161.3
R735 VP.n40 VP.n6 161.3
R736 VP.n39 VP.n38 161.3
R737 VP.n37 VP.n7 161.3
R738 VP.n40 VP.n39 56.4773
R739 VP.n59 VP.n1 56.4773
R740 VP.n31 VP.n9 56.4773
R741 VP.n15 VP.n14 49.1005
R742 VP.n47 VP.n46 47.7136
R743 VP.n52 VP.n3 47.7136
R744 VP.n24 VP.n11 47.7136
R745 VP.n19 VP.n18 47.7136
R746 VP.n36 VP.n34 46.5952
R747 VP.n46 VP.n5 33.1076
R748 VP.n53 VP.n52 33.1076
R749 VP.n25 VP.n24 33.1076
R750 VP.n18 VP.n13 33.1076
R751 VP.n39 VP.n7 24.3439
R752 VP.n42 VP.n40 24.3439
R753 VP.n48 VP.n47 24.3439
R754 VP.n48 VP.n3 24.3439
R755 VP.n55 VP.n1 24.3439
R756 VP.n60 VP.n59 24.3439
R757 VP.n32 VP.n31 24.3439
R758 VP.n27 VP.n9 24.3439
R759 VP.n20 VP.n19 24.3439
R760 VP.n20 VP.n11 24.3439
R761 VP.n16 VP.n15 17.8309
R762 VP.n41 VP.n5 17.0409
R763 VP.n54 VP.n53 17.0409
R764 VP.n26 VP.n25 17.0409
R765 VP.n14 VP.n13 17.0409
R766 VP.n35 VP.n7 9.73787
R767 VP.n61 VP.n60 9.73787
R768 VP.n33 VP.n32 9.73787
R769 VP.n42 VP.n41 7.30353
R770 VP.n55 VP.n54 7.30353
R771 VP.n27 VP.n26 7.30353
R772 VP.n17 VP.n16 0.189894
R773 VP.n17 VP.n12 0.189894
R774 VP.n21 VP.n12 0.189894
R775 VP.n22 VP.n21 0.189894
R776 VP.n23 VP.n22 0.189894
R777 VP.n23 VP.n10 0.189894
R778 VP.n28 VP.n10 0.189894
R779 VP.n29 VP.n28 0.189894
R780 VP.n30 VP.n29 0.189894
R781 VP.n30 VP.n8 0.189894
R782 VP.n34 VP.n8 0.189894
R783 VP.n37 VP.n36 0.189894
R784 VP.n38 VP.n37 0.189894
R785 VP.n38 VP.n6 0.189894
R786 VP.n43 VP.n6 0.189894
R787 VP.n44 VP.n43 0.189894
R788 VP.n45 VP.n44 0.189894
R789 VP.n45 VP.n4 0.189894
R790 VP.n49 VP.n4 0.189894
R791 VP.n50 VP.n49 0.189894
R792 VP.n51 VP.n50 0.189894
R793 VP.n51 VP.n2 0.189894
R794 VP.n56 VP.n2 0.189894
R795 VP.n57 VP.n56 0.189894
R796 VP.n58 VP.n57 0.189894
R797 VP.n58 VP.n0 0.189894
R798 VP.n62 VP.n0 0.189894
R799 VP VP.n62 0.0516364
R800 VDD1.n60 VDD1.n59 756.745
R801 VDD1.n123 VDD1.n122 756.745
R802 VDD1.n59 VDD1.n58 585
R803 VDD1.n2 VDD1.n1 585
R804 VDD1.n53 VDD1.n52 585
R805 VDD1.n51 VDD1.n50 585
R806 VDD1.n6 VDD1.n5 585
R807 VDD1.n45 VDD1.n44 585
R808 VDD1.n43 VDD1.n42 585
R809 VDD1.n10 VDD1.n9 585
R810 VDD1.n37 VDD1.n36 585
R811 VDD1.n35 VDD1.n34 585
R812 VDD1.n14 VDD1.n13 585
R813 VDD1.n29 VDD1.n28 585
R814 VDD1.n27 VDD1.n26 585
R815 VDD1.n18 VDD1.n17 585
R816 VDD1.n21 VDD1.n20 585
R817 VDD1.n84 VDD1.n83 585
R818 VDD1.n81 VDD1.n80 585
R819 VDD1.n90 VDD1.n89 585
R820 VDD1.n92 VDD1.n91 585
R821 VDD1.n77 VDD1.n76 585
R822 VDD1.n98 VDD1.n97 585
R823 VDD1.n100 VDD1.n99 585
R824 VDD1.n73 VDD1.n72 585
R825 VDD1.n106 VDD1.n105 585
R826 VDD1.n108 VDD1.n107 585
R827 VDD1.n69 VDD1.n68 585
R828 VDD1.n114 VDD1.n113 585
R829 VDD1.n116 VDD1.n115 585
R830 VDD1.n65 VDD1.n64 585
R831 VDD1.n122 VDD1.n121 585
R832 VDD1.t8 VDD1.n19 327.466
R833 VDD1.t2 VDD1.n82 327.466
R834 VDD1.n59 VDD1.n1 171.744
R835 VDD1.n52 VDD1.n1 171.744
R836 VDD1.n52 VDD1.n51 171.744
R837 VDD1.n51 VDD1.n5 171.744
R838 VDD1.n44 VDD1.n5 171.744
R839 VDD1.n44 VDD1.n43 171.744
R840 VDD1.n43 VDD1.n9 171.744
R841 VDD1.n36 VDD1.n9 171.744
R842 VDD1.n36 VDD1.n35 171.744
R843 VDD1.n35 VDD1.n13 171.744
R844 VDD1.n28 VDD1.n13 171.744
R845 VDD1.n28 VDD1.n27 171.744
R846 VDD1.n27 VDD1.n17 171.744
R847 VDD1.n20 VDD1.n17 171.744
R848 VDD1.n83 VDD1.n80 171.744
R849 VDD1.n90 VDD1.n80 171.744
R850 VDD1.n91 VDD1.n90 171.744
R851 VDD1.n91 VDD1.n76 171.744
R852 VDD1.n98 VDD1.n76 171.744
R853 VDD1.n99 VDD1.n98 171.744
R854 VDD1.n99 VDD1.n72 171.744
R855 VDD1.n106 VDD1.n72 171.744
R856 VDD1.n107 VDD1.n106 171.744
R857 VDD1.n107 VDD1.n68 171.744
R858 VDD1.n114 VDD1.n68 171.744
R859 VDD1.n115 VDD1.n114 171.744
R860 VDD1.n115 VDD1.n64 171.744
R861 VDD1.n122 VDD1.n64 171.744
R862 VDD1.n20 VDD1.t8 85.8723
R863 VDD1.n83 VDD1.t2 85.8723
R864 VDD1.n127 VDD1.n126 79.3036
R865 VDD1.n62 VDD1.n61 78.163
R866 VDD1.n125 VDD1.n124 78.1628
R867 VDD1.n129 VDD1.n128 78.1619
R868 VDD1.n62 VDD1.n60 52.3984
R869 VDD1.n125 VDD1.n123 52.3984
R870 VDD1.n129 VDD1.n127 42.3608
R871 VDD1.n21 VDD1.n19 16.3895
R872 VDD1.n84 VDD1.n82 16.3895
R873 VDD1.n22 VDD1.n18 12.8005
R874 VDD1.n85 VDD1.n81 12.8005
R875 VDD1.n26 VDD1.n25 12.0247
R876 VDD1.n89 VDD1.n88 12.0247
R877 VDD1.n58 VDD1.n0 11.249
R878 VDD1.n29 VDD1.n16 11.249
R879 VDD1.n92 VDD1.n79 11.249
R880 VDD1.n121 VDD1.n63 11.249
R881 VDD1.n57 VDD1.n2 10.4732
R882 VDD1.n30 VDD1.n14 10.4732
R883 VDD1.n93 VDD1.n77 10.4732
R884 VDD1.n120 VDD1.n65 10.4732
R885 VDD1.n54 VDD1.n53 9.69747
R886 VDD1.n34 VDD1.n33 9.69747
R887 VDD1.n97 VDD1.n96 9.69747
R888 VDD1.n117 VDD1.n116 9.69747
R889 VDD1.n56 VDD1.n0 9.45567
R890 VDD1.n119 VDD1.n63 9.45567
R891 VDD1.n47 VDD1.n46 9.3005
R892 VDD1.n49 VDD1.n48 9.3005
R893 VDD1.n4 VDD1.n3 9.3005
R894 VDD1.n55 VDD1.n54 9.3005
R895 VDD1.n57 VDD1.n56 9.3005
R896 VDD1.n8 VDD1.n7 9.3005
R897 VDD1.n41 VDD1.n40 9.3005
R898 VDD1.n39 VDD1.n38 9.3005
R899 VDD1.n12 VDD1.n11 9.3005
R900 VDD1.n33 VDD1.n32 9.3005
R901 VDD1.n31 VDD1.n30 9.3005
R902 VDD1.n16 VDD1.n15 9.3005
R903 VDD1.n25 VDD1.n24 9.3005
R904 VDD1.n23 VDD1.n22 9.3005
R905 VDD1.n71 VDD1.n70 9.3005
R906 VDD1.n110 VDD1.n109 9.3005
R907 VDD1.n112 VDD1.n111 9.3005
R908 VDD1.n67 VDD1.n66 9.3005
R909 VDD1.n118 VDD1.n117 9.3005
R910 VDD1.n120 VDD1.n119 9.3005
R911 VDD1.n102 VDD1.n101 9.3005
R912 VDD1.n75 VDD1.n74 9.3005
R913 VDD1.n96 VDD1.n95 9.3005
R914 VDD1.n94 VDD1.n93 9.3005
R915 VDD1.n79 VDD1.n78 9.3005
R916 VDD1.n88 VDD1.n87 9.3005
R917 VDD1.n86 VDD1.n85 9.3005
R918 VDD1.n104 VDD1.n103 9.3005
R919 VDD1.n50 VDD1.n4 8.92171
R920 VDD1.n37 VDD1.n12 8.92171
R921 VDD1.n100 VDD1.n75 8.92171
R922 VDD1.n113 VDD1.n67 8.92171
R923 VDD1.n49 VDD1.n6 8.14595
R924 VDD1.n38 VDD1.n10 8.14595
R925 VDD1.n101 VDD1.n73 8.14595
R926 VDD1.n112 VDD1.n69 8.14595
R927 VDD1.n46 VDD1.n45 7.3702
R928 VDD1.n42 VDD1.n41 7.3702
R929 VDD1.n105 VDD1.n104 7.3702
R930 VDD1.n109 VDD1.n108 7.3702
R931 VDD1.n45 VDD1.n8 6.59444
R932 VDD1.n42 VDD1.n8 6.59444
R933 VDD1.n105 VDD1.n71 6.59444
R934 VDD1.n108 VDD1.n71 6.59444
R935 VDD1.n46 VDD1.n6 5.81868
R936 VDD1.n41 VDD1.n10 5.81868
R937 VDD1.n104 VDD1.n73 5.81868
R938 VDD1.n109 VDD1.n69 5.81868
R939 VDD1.n50 VDD1.n49 5.04292
R940 VDD1.n38 VDD1.n37 5.04292
R941 VDD1.n101 VDD1.n100 5.04292
R942 VDD1.n113 VDD1.n112 5.04292
R943 VDD1.n53 VDD1.n4 4.26717
R944 VDD1.n34 VDD1.n12 4.26717
R945 VDD1.n97 VDD1.n75 4.26717
R946 VDD1.n116 VDD1.n67 4.26717
R947 VDD1.n23 VDD1.n19 3.70982
R948 VDD1.n86 VDD1.n82 3.70982
R949 VDD1.n54 VDD1.n2 3.49141
R950 VDD1.n33 VDD1.n14 3.49141
R951 VDD1.n96 VDD1.n77 3.49141
R952 VDD1.n117 VDD1.n65 3.49141
R953 VDD1.n128 VDD1.t4 2.8924
R954 VDD1.n128 VDD1.t9 2.8924
R955 VDD1.n61 VDD1.t3 2.8924
R956 VDD1.n61 VDD1.t0 2.8924
R957 VDD1.n126 VDD1.t7 2.8924
R958 VDD1.n126 VDD1.t1 2.8924
R959 VDD1.n124 VDD1.t5 2.8924
R960 VDD1.n124 VDD1.t6 2.8924
R961 VDD1.n58 VDD1.n57 2.71565
R962 VDD1.n30 VDD1.n29 2.71565
R963 VDD1.n93 VDD1.n92 2.71565
R964 VDD1.n121 VDD1.n120 2.71565
R965 VDD1.n60 VDD1.n0 1.93989
R966 VDD1.n26 VDD1.n16 1.93989
R967 VDD1.n89 VDD1.n79 1.93989
R968 VDD1.n123 VDD1.n63 1.93989
R969 VDD1.n25 VDD1.n18 1.16414
R970 VDD1.n88 VDD1.n81 1.16414
R971 VDD1 VDD1.n129 1.13843
R972 VDD1 VDD1.n62 0.457397
R973 VDD1.n22 VDD1.n21 0.388379
R974 VDD1.n85 VDD1.n84 0.388379
R975 VDD1.n127 VDD1.n125 0.343861
R976 VDD1.n56 VDD1.n55 0.155672
R977 VDD1.n55 VDD1.n3 0.155672
R978 VDD1.n48 VDD1.n3 0.155672
R979 VDD1.n48 VDD1.n47 0.155672
R980 VDD1.n47 VDD1.n7 0.155672
R981 VDD1.n40 VDD1.n7 0.155672
R982 VDD1.n40 VDD1.n39 0.155672
R983 VDD1.n39 VDD1.n11 0.155672
R984 VDD1.n32 VDD1.n11 0.155672
R985 VDD1.n32 VDD1.n31 0.155672
R986 VDD1.n31 VDD1.n15 0.155672
R987 VDD1.n24 VDD1.n15 0.155672
R988 VDD1.n24 VDD1.n23 0.155672
R989 VDD1.n87 VDD1.n86 0.155672
R990 VDD1.n87 VDD1.n78 0.155672
R991 VDD1.n94 VDD1.n78 0.155672
R992 VDD1.n95 VDD1.n94 0.155672
R993 VDD1.n95 VDD1.n74 0.155672
R994 VDD1.n102 VDD1.n74 0.155672
R995 VDD1.n103 VDD1.n102 0.155672
R996 VDD1.n103 VDD1.n70 0.155672
R997 VDD1.n110 VDD1.n70 0.155672
R998 VDD1.n111 VDD1.n110 0.155672
R999 VDD1.n111 VDD1.n66 0.155672
R1000 VDD1.n118 VDD1.n66 0.155672
R1001 VDD1.n119 VDD1.n118 0.155672
R1002 B.n371 B.n112 585
R1003 B.n370 B.n369 585
R1004 B.n368 B.n113 585
R1005 B.n367 B.n366 585
R1006 B.n365 B.n114 585
R1007 B.n364 B.n363 585
R1008 B.n362 B.n115 585
R1009 B.n361 B.n360 585
R1010 B.n359 B.n116 585
R1011 B.n358 B.n357 585
R1012 B.n356 B.n117 585
R1013 B.n355 B.n354 585
R1014 B.n353 B.n118 585
R1015 B.n352 B.n351 585
R1016 B.n350 B.n119 585
R1017 B.n349 B.n348 585
R1018 B.n347 B.n120 585
R1019 B.n346 B.n345 585
R1020 B.n344 B.n121 585
R1021 B.n343 B.n342 585
R1022 B.n341 B.n122 585
R1023 B.n340 B.n339 585
R1024 B.n338 B.n123 585
R1025 B.n337 B.n336 585
R1026 B.n335 B.n124 585
R1027 B.n334 B.n333 585
R1028 B.n332 B.n125 585
R1029 B.n331 B.n330 585
R1030 B.n329 B.n126 585
R1031 B.n328 B.n327 585
R1032 B.n326 B.n127 585
R1033 B.n325 B.n324 585
R1034 B.n323 B.n128 585
R1035 B.n322 B.n321 585
R1036 B.n320 B.n129 585
R1037 B.n319 B.n318 585
R1038 B.n317 B.n130 585
R1039 B.n316 B.n315 585
R1040 B.n314 B.n131 585
R1041 B.n313 B.n312 585
R1042 B.n308 B.n132 585
R1043 B.n307 B.n306 585
R1044 B.n305 B.n133 585
R1045 B.n304 B.n303 585
R1046 B.n302 B.n134 585
R1047 B.n301 B.n300 585
R1048 B.n299 B.n135 585
R1049 B.n298 B.n297 585
R1050 B.n296 B.n136 585
R1051 B.n294 B.n293 585
R1052 B.n292 B.n139 585
R1053 B.n291 B.n290 585
R1054 B.n289 B.n140 585
R1055 B.n288 B.n287 585
R1056 B.n286 B.n141 585
R1057 B.n285 B.n284 585
R1058 B.n283 B.n142 585
R1059 B.n282 B.n281 585
R1060 B.n280 B.n143 585
R1061 B.n279 B.n278 585
R1062 B.n277 B.n144 585
R1063 B.n276 B.n275 585
R1064 B.n274 B.n145 585
R1065 B.n273 B.n272 585
R1066 B.n271 B.n146 585
R1067 B.n270 B.n269 585
R1068 B.n268 B.n147 585
R1069 B.n267 B.n266 585
R1070 B.n265 B.n148 585
R1071 B.n264 B.n263 585
R1072 B.n262 B.n149 585
R1073 B.n261 B.n260 585
R1074 B.n259 B.n150 585
R1075 B.n258 B.n257 585
R1076 B.n256 B.n151 585
R1077 B.n255 B.n254 585
R1078 B.n253 B.n152 585
R1079 B.n252 B.n251 585
R1080 B.n250 B.n153 585
R1081 B.n249 B.n248 585
R1082 B.n247 B.n154 585
R1083 B.n246 B.n245 585
R1084 B.n244 B.n155 585
R1085 B.n243 B.n242 585
R1086 B.n241 B.n156 585
R1087 B.n240 B.n239 585
R1088 B.n238 B.n157 585
R1089 B.n237 B.n236 585
R1090 B.n373 B.n372 585
R1091 B.n374 B.n111 585
R1092 B.n376 B.n375 585
R1093 B.n377 B.n110 585
R1094 B.n379 B.n378 585
R1095 B.n380 B.n109 585
R1096 B.n382 B.n381 585
R1097 B.n383 B.n108 585
R1098 B.n385 B.n384 585
R1099 B.n386 B.n107 585
R1100 B.n388 B.n387 585
R1101 B.n389 B.n106 585
R1102 B.n391 B.n390 585
R1103 B.n392 B.n105 585
R1104 B.n394 B.n393 585
R1105 B.n395 B.n104 585
R1106 B.n397 B.n396 585
R1107 B.n398 B.n103 585
R1108 B.n400 B.n399 585
R1109 B.n401 B.n102 585
R1110 B.n403 B.n402 585
R1111 B.n404 B.n101 585
R1112 B.n406 B.n405 585
R1113 B.n407 B.n100 585
R1114 B.n409 B.n408 585
R1115 B.n410 B.n99 585
R1116 B.n412 B.n411 585
R1117 B.n413 B.n98 585
R1118 B.n415 B.n414 585
R1119 B.n416 B.n97 585
R1120 B.n418 B.n417 585
R1121 B.n419 B.n96 585
R1122 B.n421 B.n420 585
R1123 B.n422 B.n95 585
R1124 B.n424 B.n423 585
R1125 B.n425 B.n94 585
R1126 B.n427 B.n426 585
R1127 B.n428 B.n93 585
R1128 B.n430 B.n429 585
R1129 B.n431 B.n92 585
R1130 B.n433 B.n432 585
R1131 B.n434 B.n91 585
R1132 B.n436 B.n435 585
R1133 B.n437 B.n90 585
R1134 B.n439 B.n438 585
R1135 B.n440 B.n89 585
R1136 B.n442 B.n441 585
R1137 B.n443 B.n88 585
R1138 B.n445 B.n444 585
R1139 B.n446 B.n87 585
R1140 B.n448 B.n447 585
R1141 B.n449 B.n86 585
R1142 B.n451 B.n450 585
R1143 B.n452 B.n85 585
R1144 B.n454 B.n453 585
R1145 B.n455 B.n84 585
R1146 B.n457 B.n456 585
R1147 B.n458 B.n83 585
R1148 B.n460 B.n459 585
R1149 B.n461 B.n82 585
R1150 B.n463 B.n462 585
R1151 B.n464 B.n81 585
R1152 B.n466 B.n465 585
R1153 B.n467 B.n80 585
R1154 B.n469 B.n468 585
R1155 B.n470 B.n79 585
R1156 B.n472 B.n471 585
R1157 B.n473 B.n78 585
R1158 B.n475 B.n474 585
R1159 B.n476 B.n77 585
R1160 B.n478 B.n477 585
R1161 B.n479 B.n76 585
R1162 B.n481 B.n480 585
R1163 B.n482 B.n75 585
R1164 B.n484 B.n483 585
R1165 B.n485 B.n74 585
R1166 B.n487 B.n486 585
R1167 B.n488 B.n73 585
R1168 B.n490 B.n489 585
R1169 B.n491 B.n72 585
R1170 B.n493 B.n492 585
R1171 B.n494 B.n71 585
R1172 B.n627 B.n22 585
R1173 B.n626 B.n625 585
R1174 B.n624 B.n23 585
R1175 B.n623 B.n622 585
R1176 B.n621 B.n24 585
R1177 B.n620 B.n619 585
R1178 B.n618 B.n25 585
R1179 B.n617 B.n616 585
R1180 B.n615 B.n26 585
R1181 B.n614 B.n613 585
R1182 B.n612 B.n27 585
R1183 B.n611 B.n610 585
R1184 B.n609 B.n28 585
R1185 B.n608 B.n607 585
R1186 B.n606 B.n29 585
R1187 B.n605 B.n604 585
R1188 B.n603 B.n30 585
R1189 B.n602 B.n601 585
R1190 B.n600 B.n31 585
R1191 B.n599 B.n598 585
R1192 B.n597 B.n32 585
R1193 B.n596 B.n595 585
R1194 B.n594 B.n33 585
R1195 B.n593 B.n592 585
R1196 B.n591 B.n34 585
R1197 B.n590 B.n589 585
R1198 B.n588 B.n35 585
R1199 B.n587 B.n586 585
R1200 B.n585 B.n36 585
R1201 B.n584 B.n583 585
R1202 B.n582 B.n37 585
R1203 B.n581 B.n580 585
R1204 B.n579 B.n38 585
R1205 B.n578 B.n577 585
R1206 B.n576 B.n39 585
R1207 B.n575 B.n574 585
R1208 B.n573 B.n40 585
R1209 B.n572 B.n571 585
R1210 B.n570 B.n41 585
R1211 B.n568 B.n567 585
R1212 B.n566 B.n44 585
R1213 B.n565 B.n564 585
R1214 B.n563 B.n45 585
R1215 B.n562 B.n561 585
R1216 B.n560 B.n46 585
R1217 B.n559 B.n558 585
R1218 B.n557 B.n47 585
R1219 B.n556 B.n555 585
R1220 B.n554 B.n48 585
R1221 B.n553 B.n552 585
R1222 B.n551 B.n49 585
R1223 B.n550 B.n549 585
R1224 B.n548 B.n53 585
R1225 B.n547 B.n546 585
R1226 B.n545 B.n54 585
R1227 B.n544 B.n543 585
R1228 B.n542 B.n55 585
R1229 B.n541 B.n540 585
R1230 B.n539 B.n56 585
R1231 B.n538 B.n537 585
R1232 B.n536 B.n57 585
R1233 B.n535 B.n534 585
R1234 B.n533 B.n58 585
R1235 B.n532 B.n531 585
R1236 B.n530 B.n59 585
R1237 B.n529 B.n528 585
R1238 B.n527 B.n60 585
R1239 B.n526 B.n525 585
R1240 B.n524 B.n61 585
R1241 B.n523 B.n522 585
R1242 B.n521 B.n62 585
R1243 B.n520 B.n519 585
R1244 B.n518 B.n63 585
R1245 B.n517 B.n516 585
R1246 B.n515 B.n64 585
R1247 B.n514 B.n513 585
R1248 B.n512 B.n65 585
R1249 B.n511 B.n510 585
R1250 B.n509 B.n66 585
R1251 B.n508 B.n507 585
R1252 B.n506 B.n67 585
R1253 B.n505 B.n504 585
R1254 B.n503 B.n68 585
R1255 B.n502 B.n501 585
R1256 B.n500 B.n69 585
R1257 B.n499 B.n498 585
R1258 B.n497 B.n70 585
R1259 B.n496 B.n495 585
R1260 B.n629 B.n628 585
R1261 B.n630 B.n21 585
R1262 B.n632 B.n631 585
R1263 B.n633 B.n20 585
R1264 B.n635 B.n634 585
R1265 B.n636 B.n19 585
R1266 B.n638 B.n637 585
R1267 B.n639 B.n18 585
R1268 B.n641 B.n640 585
R1269 B.n642 B.n17 585
R1270 B.n644 B.n643 585
R1271 B.n645 B.n16 585
R1272 B.n647 B.n646 585
R1273 B.n648 B.n15 585
R1274 B.n650 B.n649 585
R1275 B.n651 B.n14 585
R1276 B.n653 B.n652 585
R1277 B.n654 B.n13 585
R1278 B.n656 B.n655 585
R1279 B.n657 B.n12 585
R1280 B.n659 B.n658 585
R1281 B.n660 B.n11 585
R1282 B.n662 B.n661 585
R1283 B.n663 B.n10 585
R1284 B.n665 B.n664 585
R1285 B.n666 B.n9 585
R1286 B.n668 B.n667 585
R1287 B.n669 B.n8 585
R1288 B.n671 B.n670 585
R1289 B.n672 B.n7 585
R1290 B.n674 B.n673 585
R1291 B.n675 B.n6 585
R1292 B.n677 B.n676 585
R1293 B.n678 B.n5 585
R1294 B.n680 B.n679 585
R1295 B.n681 B.n4 585
R1296 B.n683 B.n682 585
R1297 B.n684 B.n3 585
R1298 B.n686 B.n685 585
R1299 B.n687 B.n0 585
R1300 B.n2 B.n1 585
R1301 B.n178 B.n177 585
R1302 B.n180 B.n179 585
R1303 B.n181 B.n176 585
R1304 B.n183 B.n182 585
R1305 B.n184 B.n175 585
R1306 B.n186 B.n185 585
R1307 B.n187 B.n174 585
R1308 B.n189 B.n188 585
R1309 B.n190 B.n173 585
R1310 B.n192 B.n191 585
R1311 B.n193 B.n172 585
R1312 B.n195 B.n194 585
R1313 B.n196 B.n171 585
R1314 B.n198 B.n197 585
R1315 B.n199 B.n170 585
R1316 B.n201 B.n200 585
R1317 B.n202 B.n169 585
R1318 B.n204 B.n203 585
R1319 B.n205 B.n168 585
R1320 B.n207 B.n206 585
R1321 B.n208 B.n167 585
R1322 B.n210 B.n209 585
R1323 B.n211 B.n166 585
R1324 B.n213 B.n212 585
R1325 B.n214 B.n165 585
R1326 B.n216 B.n215 585
R1327 B.n217 B.n164 585
R1328 B.n219 B.n218 585
R1329 B.n220 B.n163 585
R1330 B.n222 B.n221 585
R1331 B.n223 B.n162 585
R1332 B.n225 B.n224 585
R1333 B.n226 B.n161 585
R1334 B.n228 B.n227 585
R1335 B.n229 B.n160 585
R1336 B.n231 B.n230 585
R1337 B.n232 B.n159 585
R1338 B.n234 B.n233 585
R1339 B.n235 B.n158 585
R1340 B.n237 B.n158 569.379
R1341 B.n373 B.n112 569.379
R1342 B.n495 B.n494 569.379
R1343 B.n628 B.n627 569.379
R1344 B.n309 B.t4 397.611
R1345 B.n50 B.t2 397.611
R1346 B.n137 B.t7 397.611
R1347 B.n42 B.t11 397.611
R1348 B.n137 B.t6 383.726
R1349 B.n309 B.t3 383.726
R1350 B.n50 B.t0 383.726
R1351 B.n42 B.t9 383.726
R1352 B.n310 B.t5 361.733
R1353 B.n51 B.t1 361.733
R1354 B.n138 B.t8 361.733
R1355 B.n43 B.t10 361.733
R1356 B.n689 B.n688 256.663
R1357 B.n688 B.n687 235.042
R1358 B.n688 B.n2 235.042
R1359 B.n238 B.n237 163.367
R1360 B.n239 B.n238 163.367
R1361 B.n239 B.n156 163.367
R1362 B.n243 B.n156 163.367
R1363 B.n244 B.n243 163.367
R1364 B.n245 B.n244 163.367
R1365 B.n245 B.n154 163.367
R1366 B.n249 B.n154 163.367
R1367 B.n250 B.n249 163.367
R1368 B.n251 B.n250 163.367
R1369 B.n251 B.n152 163.367
R1370 B.n255 B.n152 163.367
R1371 B.n256 B.n255 163.367
R1372 B.n257 B.n256 163.367
R1373 B.n257 B.n150 163.367
R1374 B.n261 B.n150 163.367
R1375 B.n262 B.n261 163.367
R1376 B.n263 B.n262 163.367
R1377 B.n263 B.n148 163.367
R1378 B.n267 B.n148 163.367
R1379 B.n268 B.n267 163.367
R1380 B.n269 B.n268 163.367
R1381 B.n269 B.n146 163.367
R1382 B.n273 B.n146 163.367
R1383 B.n274 B.n273 163.367
R1384 B.n275 B.n274 163.367
R1385 B.n275 B.n144 163.367
R1386 B.n279 B.n144 163.367
R1387 B.n280 B.n279 163.367
R1388 B.n281 B.n280 163.367
R1389 B.n281 B.n142 163.367
R1390 B.n285 B.n142 163.367
R1391 B.n286 B.n285 163.367
R1392 B.n287 B.n286 163.367
R1393 B.n287 B.n140 163.367
R1394 B.n291 B.n140 163.367
R1395 B.n292 B.n291 163.367
R1396 B.n293 B.n292 163.367
R1397 B.n293 B.n136 163.367
R1398 B.n298 B.n136 163.367
R1399 B.n299 B.n298 163.367
R1400 B.n300 B.n299 163.367
R1401 B.n300 B.n134 163.367
R1402 B.n304 B.n134 163.367
R1403 B.n305 B.n304 163.367
R1404 B.n306 B.n305 163.367
R1405 B.n306 B.n132 163.367
R1406 B.n313 B.n132 163.367
R1407 B.n314 B.n313 163.367
R1408 B.n315 B.n314 163.367
R1409 B.n315 B.n130 163.367
R1410 B.n319 B.n130 163.367
R1411 B.n320 B.n319 163.367
R1412 B.n321 B.n320 163.367
R1413 B.n321 B.n128 163.367
R1414 B.n325 B.n128 163.367
R1415 B.n326 B.n325 163.367
R1416 B.n327 B.n326 163.367
R1417 B.n327 B.n126 163.367
R1418 B.n331 B.n126 163.367
R1419 B.n332 B.n331 163.367
R1420 B.n333 B.n332 163.367
R1421 B.n333 B.n124 163.367
R1422 B.n337 B.n124 163.367
R1423 B.n338 B.n337 163.367
R1424 B.n339 B.n338 163.367
R1425 B.n339 B.n122 163.367
R1426 B.n343 B.n122 163.367
R1427 B.n344 B.n343 163.367
R1428 B.n345 B.n344 163.367
R1429 B.n345 B.n120 163.367
R1430 B.n349 B.n120 163.367
R1431 B.n350 B.n349 163.367
R1432 B.n351 B.n350 163.367
R1433 B.n351 B.n118 163.367
R1434 B.n355 B.n118 163.367
R1435 B.n356 B.n355 163.367
R1436 B.n357 B.n356 163.367
R1437 B.n357 B.n116 163.367
R1438 B.n361 B.n116 163.367
R1439 B.n362 B.n361 163.367
R1440 B.n363 B.n362 163.367
R1441 B.n363 B.n114 163.367
R1442 B.n367 B.n114 163.367
R1443 B.n368 B.n367 163.367
R1444 B.n369 B.n368 163.367
R1445 B.n369 B.n112 163.367
R1446 B.n494 B.n493 163.367
R1447 B.n493 B.n72 163.367
R1448 B.n489 B.n72 163.367
R1449 B.n489 B.n488 163.367
R1450 B.n488 B.n487 163.367
R1451 B.n487 B.n74 163.367
R1452 B.n483 B.n74 163.367
R1453 B.n483 B.n482 163.367
R1454 B.n482 B.n481 163.367
R1455 B.n481 B.n76 163.367
R1456 B.n477 B.n76 163.367
R1457 B.n477 B.n476 163.367
R1458 B.n476 B.n475 163.367
R1459 B.n475 B.n78 163.367
R1460 B.n471 B.n78 163.367
R1461 B.n471 B.n470 163.367
R1462 B.n470 B.n469 163.367
R1463 B.n469 B.n80 163.367
R1464 B.n465 B.n80 163.367
R1465 B.n465 B.n464 163.367
R1466 B.n464 B.n463 163.367
R1467 B.n463 B.n82 163.367
R1468 B.n459 B.n82 163.367
R1469 B.n459 B.n458 163.367
R1470 B.n458 B.n457 163.367
R1471 B.n457 B.n84 163.367
R1472 B.n453 B.n84 163.367
R1473 B.n453 B.n452 163.367
R1474 B.n452 B.n451 163.367
R1475 B.n451 B.n86 163.367
R1476 B.n447 B.n86 163.367
R1477 B.n447 B.n446 163.367
R1478 B.n446 B.n445 163.367
R1479 B.n445 B.n88 163.367
R1480 B.n441 B.n88 163.367
R1481 B.n441 B.n440 163.367
R1482 B.n440 B.n439 163.367
R1483 B.n439 B.n90 163.367
R1484 B.n435 B.n90 163.367
R1485 B.n435 B.n434 163.367
R1486 B.n434 B.n433 163.367
R1487 B.n433 B.n92 163.367
R1488 B.n429 B.n92 163.367
R1489 B.n429 B.n428 163.367
R1490 B.n428 B.n427 163.367
R1491 B.n427 B.n94 163.367
R1492 B.n423 B.n94 163.367
R1493 B.n423 B.n422 163.367
R1494 B.n422 B.n421 163.367
R1495 B.n421 B.n96 163.367
R1496 B.n417 B.n96 163.367
R1497 B.n417 B.n416 163.367
R1498 B.n416 B.n415 163.367
R1499 B.n415 B.n98 163.367
R1500 B.n411 B.n98 163.367
R1501 B.n411 B.n410 163.367
R1502 B.n410 B.n409 163.367
R1503 B.n409 B.n100 163.367
R1504 B.n405 B.n100 163.367
R1505 B.n405 B.n404 163.367
R1506 B.n404 B.n403 163.367
R1507 B.n403 B.n102 163.367
R1508 B.n399 B.n102 163.367
R1509 B.n399 B.n398 163.367
R1510 B.n398 B.n397 163.367
R1511 B.n397 B.n104 163.367
R1512 B.n393 B.n104 163.367
R1513 B.n393 B.n392 163.367
R1514 B.n392 B.n391 163.367
R1515 B.n391 B.n106 163.367
R1516 B.n387 B.n106 163.367
R1517 B.n387 B.n386 163.367
R1518 B.n386 B.n385 163.367
R1519 B.n385 B.n108 163.367
R1520 B.n381 B.n108 163.367
R1521 B.n381 B.n380 163.367
R1522 B.n380 B.n379 163.367
R1523 B.n379 B.n110 163.367
R1524 B.n375 B.n110 163.367
R1525 B.n375 B.n374 163.367
R1526 B.n374 B.n373 163.367
R1527 B.n627 B.n626 163.367
R1528 B.n626 B.n23 163.367
R1529 B.n622 B.n23 163.367
R1530 B.n622 B.n621 163.367
R1531 B.n621 B.n620 163.367
R1532 B.n620 B.n25 163.367
R1533 B.n616 B.n25 163.367
R1534 B.n616 B.n615 163.367
R1535 B.n615 B.n614 163.367
R1536 B.n614 B.n27 163.367
R1537 B.n610 B.n27 163.367
R1538 B.n610 B.n609 163.367
R1539 B.n609 B.n608 163.367
R1540 B.n608 B.n29 163.367
R1541 B.n604 B.n29 163.367
R1542 B.n604 B.n603 163.367
R1543 B.n603 B.n602 163.367
R1544 B.n602 B.n31 163.367
R1545 B.n598 B.n31 163.367
R1546 B.n598 B.n597 163.367
R1547 B.n597 B.n596 163.367
R1548 B.n596 B.n33 163.367
R1549 B.n592 B.n33 163.367
R1550 B.n592 B.n591 163.367
R1551 B.n591 B.n590 163.367
R1552 B.n590 B.n35 163.367
R1553 B.n586 B.n35 163.367
R1554 B.n586 B.n585 163.367
R1555 B.n585 B.n584 163.367
R1556 B.n584 B.n37 163.367
R1557 B.n580 B.n37 163.367
R1558 B.n580 B.n579 163.367
R1559 B.n579 B.n578 163.367
R1560 B.n578 B.n39 163.367
R1561 B.n574 B.n39 163.367
R1562 B.n574 B.n573 163.367
R1563 B.n573 B.n572 163.367
R1564 B.n572 B.n41 163.367
R1565 B.n567 B.n41 163.367
R1566 B.n567 B.n566 163.367
R1567 B.n566 B.n565 163.367
R1568 B.n565 B.n45 163.367
R1569 B.n561 B.n45 163.367
R1570 B.n561 B.n560 163.367
R1571 B.n560 B.n559 163.367
R1572 B.n559 B.n47 163.367
R1573 B.n555 B.n47 163.367
R1574 B.n555 B.n554 163.367
R1575 B.n554 B.n553 163.367
R1576 B.n553 B.n49 163.367
R1577 B.n549 B.n49 163.367
R1578 B.n549 B.n548 163.367
R1579 B.n548 B.n547 163.367
R1580 B.n547 B.n54 163.367
R1581 B.n543 B.n54 163.367
R1582 B.n543 B.n542 163.367
R1583 B.n542 B.n541 163.367
R1584 B.n541 B.n56 163.367
R1585 B.n537 B.n56 163.367
R1586 B.n537 B.n536 163.367
R1587 B.n536 B.n535 163.367
R1588 B.n535 B.n58 163.367
R1589 B.n531 B.n58 163.367
R1590 B.n531 B.n530 163.367
R1591 B.n530 B.n529 163.367
R1592 B.n529 B.n60 163.367
R1593 B.n525 B.n60 163.367
R1594 B.n525 B.n524 163.367
R1595 B.n524 B.n523 163.367
R1596 B.n523 B.n62 163.367
R1597 B.n519 B.n62 163.367
R1598 B.n519 B.n518 163.367
R1599 B.n518 B.n517 163.367
R1600 B.n517 B.n64 163.367
R1601 B.n513 B.n64 163.367
R1602 B.n513 B.n512 163.367
R1603 B.n512 B.n511 163.367
R1604 B.n511 B.n66 163.367
R1605 B.n507 B.n66 163.367
R1606 B.n507 B.n506 163.367
R1607 B.n506 B.n505 163.367
R1608 B.n505 B.n68 163.367
R1609 B.n501 B.n68 163.367
R1610 B.n501 B.n500 163.367
R1611 B.n500 B.n499 163.367
R1612 B.n499 B.n70 163.367
R1613 B.n495 B.n70 163.367
R1614 B.n628 B.n21 163.367
R1615 B.n632 B.n21 163.367
R1616 B.n633 B.n632 163.367
R1617 B.n634 B.n633 163.367
R1618 B.n634 B.n19 163.367
R1619 B.n638 B.n19 163.367
R1620 B.n639 B.n638 163.367
R1621 B.n640 B.n639 163.367
R1622 B.n640 B.n17 163.367
R1623 B.n644 B.n17 163.367
R1624 B.n645 B.n644 163.367
R1625 B.n646 B.n645 163.367
R1626 B.n646 B.n15 163.367
R1627 B.n650 B.n15 163.367
R1628 B.n651 B.n650 163.367
R1629 B.n652 B.n651 163.367
R1630 B.n652 B.n13 163.367
R1631 B.n656 B.n13 163.367
R1632 B.n657 B.n656 163.367
R1633 B.n658 B.n657 163.367
R1634 B.n658 B.n11 163.367
R1635 B.n662 B.n11 163.367
R1636 B.n663 B.n662 163.367
R1637 B.n664 B.n663 163.367
R1638 B.n664 B.n9 163.367
R1639 B.n668 B.n9 163.367
R1640 B.n669 B.n668 163.367
R1641 B.n670 B.n669 163.367
R1642 B.n670 B.n7 163.367
R1643 B.n674 B.n7 163.367
R1644 B.n675 B.n674 163.367
R1645 B.n676 B.n675 163.367
R1646 B.n676 B.n5 163.367
R1647 B.n680 B.n5 163.367
R1648 B.n681 B.n680 163.367
R1649 B.n682 B.n681 163.367
R1650 B.n682 B.n3 163.367
R1651 B.n686 B.n3 163.367
R1652 B.n687 B.n686 163.367
R1653 B.n178 B.n2 163.367
R1654 B.n179 B.n178 163.367
R1655 B.n179 B.n176 163.367
R1656 B.n183 B.n176 163.367
R1657 B.n184 B.n183 163.367
R1658 B.n185 B.n184 163.367
R1659 B.n185 B.n174 163.367
R1660 B.n189 B.n174 163.367
R1661 B.n190 B.n189 163.367
R1662 B.n191 B.n190 163.367
R1663 B.n191 B.n172 163.367
R1664 B.n195 B.n172 163.367
R1665 B.n196 B.n195 163.367
R1666 B.n197 B.n196 163.367
R1667 B.n197 B.n170 163.367
R1668 B.n201 B.n170 163.367
R1669 B.n202 B.n201 163.367
R1670 B.n203 B.n202 163.367
R1671 B.n203 B.n168 163.367
R1672 B.n207 B.n168 163.367
R1673 B.n208 B.n207 163.367
R1674 B.n209 B.n208 163.367
R1675 B.n209 B.n166 163.367
R1676 B.n213 B.n166 163.367
R1677 B.n214 B.n213 163.367
R1678 B.n215 B.n214 163.367
R1679 B.n215 B.n164 163.367
R1680 B.n219 B.n164 163.367
R1681 B.n220 B.n219 163.367
R1682 B.n221 B.n220 163.367
R1683 B.n221 B.n162 163.367
R1684 B.n225 B.n162 163.367
R1685 B.n226 B.n225 163.367
R1686 B.n227 B.n226 163.367
R1687 B.n227 B.n160 163.367
R1688 B.n231 B.n160 163.367
R1689 B.n232 B.n231 163.367
R1690 B.n233 B.n232 163.367
R1691 B.n233 B.n158 163.367
R1692 B.n295 B.n138 59.5399
R1693 B.n311 B.n310 59.5399
R1694 B.n52 B.n51 59.5399
R1695 B.n569 B.n43 59.5399
R1696 B.n629 B.n22 36.9956
R1697 B.n496 B.n71 36.9956
R1698 B.n372 B.n371 36.9956
R1699 B.n236 B.n235 36.9956
R1700 B.n138 B.n137 35.8793
R1701 B.n310 B.n309 35.8793
R1702 B.n51 B.n50 35.8793
R1703 B.n43 B.n42 35.8793
R1704 B B.n689 18.0485
R1705 B.n630 B.n629 10.6151
R1706 B.n631 B.n630 10.6151
R1707 B.n631 B.n20 10.6151
R1708 B.n635 B.n20 10.6151
R1709 B.n636 B.n635 10.6151
R1710 B.n637 B.n636 10.6151
R1711 B.n637 B.n18 10.6151
R1712 B.n641 B.n18 10.6151
R1713 B.n642 B.n641 10.6151
R1714 B.n643 B.n642 10.6151
R1715 B.n643 B.n16 10.6151
R1716 B.n647 B.n16 10.6151
R1717 B.n648 B.n647 10.6151
R1718 B.n649 B.n648 10.6151
R1719 B.n649 B.n14 10.6151
R1720 B.n653 B.n14 10.6151
R1721 B.n654 B.n653 10.6151
R1722 B.n655 B.n654 10.6151
R1723 B.n655 B.n12 10.6151
R1724 B.n659 B.n12 10.6151
R1725 B.n660 B.n659 10.6151
R1726 B.n661 B.n660 10.6151
R1727 B.n661 B.n10 10.6151
R1728 B.n665 B.n10 10.6151
R1729 B.n666 B.n665 10.6151
R1730 B.n667 B.n666 10.6151
R1731 B.n667 B.n8 10.6151
R1732 B.n671 B.n8 10.6151
R1733 B.n672 B.n671 10.6151
R1734 B.n673 B.n672 10.6151
R1735 B.n673 B.n6 10.6151
R1736 B.n677 B.n6 10.6151
R1737 B.n678 B.n677 10.6151
R1738 B.n679 B.n678 10.6151
R1739 B.n679 B.n4 10.6151
R1740 B.n683 B.n4 10.6151
R1741 B.n684 B.n683 10.6151
R1742 B.n685 B.n684 10.6151
R1743 B.n685 B.n0 10.6151
R1744 B.n625 B.n22 10.6151
R1745 B.n625 B.n624 10.6151
R1746 B.n624 B.n623 10.6151
R1747 B.n623 B.n24 10.6151
R1748 B.n619 B.n24 10.6151
R1749 B.n619 B.n618 10.6151
R1750 B.n618 B.n617 10.6151
R1751 B.n617 B.n26 10.6151
R1752 B.n613 B.n26 10.6151
R1753 B.n613 B.n612 10.6151
R1754 B.n612 B.n611 10.6151
R1755 B.n611 B.n28 10.6151
R1756 B.n607 B.n28 10.6151
R1757 B.n607 B.n606 10.6151
R1758 B.n606 B.n605 10.6151
R1759 B.n605 B.n30 10.6151
R1760 B.n601 B.n30 10.6151
R1761 B.n601 B.n600 10.6151
R1762 B.n600 B.n599 10.6151
R1763 B.n599 B.n32 10.6151
R1764 B.n595 B.n32 10.6151
R1765 B.n595 B.n594 10.6151
R1766 B.n594 B.n593 10.6151
R1767 B.n593 B.n34 10.6151
R1768 B.n589 B.n34 10.6151
R1769 B.n589 B.n588 10.6151
R1770 B.n588 B.n587 10.6151
R1771 B.n587 B.n36 10.6151
R1772 B.n583 B.n36 10.6151
R1773 B.n583 B.n582 10.6151
R1774 B.n582 B.n581 10.6151
R1775 B.n581 B.n38 10.6151
R1776 B.n577 B.n38 10.6151
R1777 B.n577 B.n576 10.6151
R1778 B.n576 B.n575 10.6151
R1779 B.n575 B.n40 10.6151
R1780 B.n571 B.n40 10.6151
R1781 B.n571 B.n570 10.6151
R1782 B.n568 B.n44 10.6151
R1783 B.n564 B.n44 10.6151
R1784 B.n564 B.n563 10.6151
R1785 B.n563 B.n562 10.6151
R1786 B.n562 B.n46 10.6151
R1787 B.n558 B.n46 10.6151
R1788 B.n558 B.n557 10.6151
R1789 B.n557 B.n556 10.6151
R1790 B.n556 B.n48 10.6151
R1791 B.n552 B.n551 10.6151
R1792 B.n551 B.n550 10.6151
R1793 B.n550 B.n53 10.6151
R1794 B.n546 B.n53 10.6151
R1795 B.n546 B.n545 10.6151
R1796 B.n545 B.n544 10.6151
R1797 B.n544 B.n55 10.6151
R1798 B.n540 B.n55 10.6151
R1799 B.n540 B.n539 10.6151
R1800 B.n539 B.n538 10.6151
R1801 B.n538 B.n57 10.6151
R1802 B.n534 B.n57 10.6151
R1803 B.n534 B.n533 10.6151
R1804 B.n533 B.n532 10.6151
R1805 B.n532 B.n59 10.6151
R1806 B.n528 B.n59 10.6151
R1807 B.n528 B.n527 10.6151
R1808 B.n527 B.n526 10.6151
R1809 B.n526 B.n61 10.6151
R1810 B.n522 B.n61 10.6151
R1811 B.n522 B.n521 10.6151
R1812 B.n521 B.n520 10.6151
R1813 B.n520 B.n63 10.6151
R1814 B.n516 B.n63 10.6151
R1815 B.n516 B.n515 10.6151
R1816 B.n515 B.n514 10.6151
R1817 B.n514 B.n65 10.6151
R1818 B.n510 B.n65 10.6151
R1819 B.n510 B.n509 10.6151
R1820 B.n509 B.n508 10.6151
R1821 B.n508 B.n67 10.6151
R1822 B.n504 B.n67 10.6151
R1823 B.n504 B.n503 10.6151
R1824 B.n503 B.n502 10.6151
R1825 B.n502 B.n69 10.6151
R1826 B.n498 B.n69 10.6151
R1827 B.n498 B.n497 10.6151
R1828 B.n497 B.n496 10.6151
R1829 B.n492 B.n71 10.6151
R1830 B.n492 B.n491 10.6151
R1831 B.n491 B.n490 10.6151
R1832 B.n490 B.n73 10.6151
R1833 B.n486 B.n73 10.6151
R1834 B.n486 B.n485 10.6151
R1835 B.n485 B.n484 10.6151
R1836 B.n484 B.n75 10.6151
R1837 B.n480 B.n75 10.6151
R1838 B.n480 B.n479 10.6151
R1839 B.n479 B.n478 10.6151
R1840 B.n478 B.n77 10.6151
R1841 B.n474 B.n77 10.6151
R1842 B.n474 B.n473 10.6151
R1843 B.n473 B.n472 10.6151
R1844 B.n472 B.n79 10.6151
R1845 B.n468 B.n79 10.6151
R1846 B.n468 B.n467 10.6151
R1847 B.n467 B.n466 10.6151
R1848 B.n466 B.n81 10.6151
R1849 B.n462 B.n81 10.6151
R1850 B.n462 B.n461 10.6151
R1851 B.n461 B.n460 10.6151
R1852 B.n460 B.n83 10.6151
R1853 B.n456 B.n83 10.6151
R1854 B.n456 B.n455 10.6151
R1855 B.n455 B.n454 10.6151
R1856 B.n454 B.n85 10.6151
R1857 B.n450 B.n85 10.6151
R1858 B.n450 B.n449 10.6151
R1859 B.n449 B.n448 10.6151
R1860 B.n448 B.n87 10.6151
R1861 B.n444 B.n87 10.6151
R1862 B.n444 B.n443 10.6151
R1863 B.n443 B.n442 10.6151
R1864 B.n442 B.n89 10.6151
R1865 B.n438 B.n89 10.6151
R1866 B.n438 B.n437 10.6151
R1867 B.n437 B.n436 10.6151
R1868 B.n436 B.n91 10.6151
R1869 B.n432 B.n91 10.6151
R1870 B.n432 B.n431 10.6151
R1871 B.n431 B.n430 10.6151
R1872 B.n430 B.n93 10.6151
R1873 B.n426 B.n93 10.6151
R1874 B.n426 B.n425 10.6151
R1875 B.n425 B.n424 10.6151
R1876 B.n424 B.n95 10.6151
R1877 B.n420 B.n95 10.6151
R1878 B.n420 B.n419 10.6151
R1879 B.n419 B.n418 10.6151
R1880 B.n418 B.n97 10.6151
R1881 B.n414 B.n97 10.6151
R1882 B.n414 B.n413 10.6151
R1883 B.n413 B.n412 10.6151
R1884 B.n412 B.n99 10.6151
R1885 B.n408 B.n99 10.6151
R1886 B.n408 B.n407 10.6151
R1887 B.n407 B.n406 10.6151
R1888 B.n406 B.n101 10.6151
R1889 B.n402 B.n101 10.6151
R1890 B.n402 B.n401 10.6151
R1891 B.n401 B.n400 10.6151
R1892 B.n400 B.n103 10.6151
R1893 B.n396 B.n103 10.6151
R1894 B.n396 B.n395 10.6151
R1895 B.n395 B.n394 10.6151
R1896 B.n394 B.n105 10.6151
R1897 B.n390 B.n105 10.6151
R1898 B.n390 B.n389 10.6151
R1899 B.n389 B.n388 10.6151
R1900 B.n388 B.n107 10.6151
R1901 B.n384 B.n107 10.6151
R1902 B.n384 B.n383 10.6151
R1903 B.n383 B.n382 10.6151
R1904 B.n382 B.n109 10.6151
R1905 B.n378 B.n109 10.6151
R1906 B.n378 B.n377 10.6151
R1907 B.n377 B.n376 10.6151
R1908 B.n376 B.n111 10.6151
R1909 B.n372 B.n111 10.6151
R1910 B.n177 B.n1 10.6151
R1911 B.n180 B.n177 10.6151
R1912 B.n181 B.n180 10.6151
R1913 B.n182 B.n181 10.6151
R1914 B.n182 B.n175 10.6151
R1915 B.n186 B.n175 10.6151
R1916 B.n187 B.n186 10.6151
R1917 B.n188 B.n187 10.6151
R1918 B.n188 B.n173 10.6151
R1919 B.n192 B.n173 10.6151
R1920 B.n193 B.n192 10.6151
R1921 B.n194 B.n193 10.6151
R1922 B.n194 B.n171 10.6151
R1923 B.n198 B.n171 10.6151
R1924 B.n199 B.n198 10.6151
R1925 B.n200 B.n199 10.6151
R1926 B.n200 B.n169 10.6151
R1927 B.n204 B.n169 10.6151
R1928 B.n205 B.n204 10.6151
R1929 B.n206 B.n205 10.6151
R1930 B.n206 B.n167 10.6151
R1931 B.n210 B.n167 10.6151
R1932 B.n211 B.n210 10.6151
R1933 B.n212 B.n211 10.6151
R1934 B.n212 B.n165 10.6151
R1935 B.n216 B.n165 10.6151
R1936 B.n217 B.n216 10.6151
R1937 B.n218 B.n217 10.6151
R1938 B.n218 B.n163 10.6151
R1939 B.n222 B.n163 10.6151
R1940 B.n223 B.n222 10.6151
R1941 B.n224 B.n223 10.6151
R1942 B.n224 B.n161 10.6151
R1943 B.n228 B.n161 10.6151
R1944 B.n229 B.n228 10.6151
R1945 B.n230 B.n229 10.6151
R1946 B.n230 B.n159 10.6151
R1947 B.n234 B.n159 10.6151
R1948 B.n235 B.n234 10.6151
R1949 B.n236 B.n157 10.6151
R1950 B.n240 B.n157 10.6151
R1951 B.n241 B.n240 10.6151
R1952 B.n242 B.n241 10.6151
R1953 B.n242 B.n155 10.6151
R1954 B.n246 B.n155 10.6151
R1955 B.n247 B.n246 10.6151
R1956 B.n248 B.n247 10.6151
R1957 B.n248 B.n153 10.6151
R1958 B.n252 B.n153 10.6151
R1959 B.n253 B.n252 10.6151
R1960 B.n254 B.n253 10.6151
R1961 B.n254 B.n151 10.6151
R1962 B.n258 B.n151 10.6151
R1963 B.n259 B.n258 10.6151
R1964 B.n260 B.n259 10.6151
R1965 B.n260 B.n149 10.6151
R1966 B.n264 B.n149 10.6151
R1967 B.n265 B.n264 10.6151
R1968 B.n266 B.n265 10.6151
R1969 B.n266 B.n147 10.6151
R1970 B.n270 B.n147 10.6151
R1971 B.n271 B.n270 10.6151
R1972 B.n272 B.n271 10.6151
R1973 B.n272 B.n145 10.6151
R1974 B.n276 B.n145 10.6151
R1975 B.n277 B.n276 10.6151
R1976 B.n278 B.n277 10.6151
R1977 B.n278 B.n143 10.6151
R1978 B.n282 B.n143 10.6151
R1979 B.n283 B.n282 10.6151
R1980 B.n284 B.n283 10.6151
R1981 B.n284 B.n141 10.6151
R1982 B.n288 B.n141 10.6151
R1983 B.n289 B.n288 10.6151
R1984 B.n290 B.n289 10.6151
R1985 B.n290 B.n139 10.6151
R1986 B.n294 B.n139 10.6151
R1987 B.n297 B.n296 10.6151
R1988 B.n297 B.n135 10.6151
R1989 B.n301 B.n135 10.6151
R1990 B.n302 B.n301 10.6151
R1991 B.n303 B.n302 10.6151
R1992 B.n303 B.n133 10.6151
R1993 B.n307 B.n133 10.6151
R1994 B.n308 B.n307 10.6151
R1995 B.n312 B.n308 10.6151
R1996 B.n316 B.n131 10.6151
R1997 B.n317 B.n316 10.6151
R1998 B.n318 B.n317 10.6151
R1999 B.n318 B.n129 10.6151
R2000 B.n322 B.n129 10.6151
R2001 B.n323 B.n322 10.6151
R2002 B.n324 B.n323 10.6151
R2003 B.n324 B.n127 10.6151
R2004 B.n328 B.n127 10.6151
R2005 B.n329 B.n328 10.6151
R2006 B.n330 B.n329 10.6151
R2007 B.n330 B.n125 10.6151
R2008 B.n334 B.n125 10.6151
R2009 B.n335 B.n334 10.6151
R2010 B.n336 B.n335 10.6151
R2011 B.n336 B.n123 10.6151
R2012 B.n340 B.n123 10.6151
R2013 B.n341 B.n340 10.6151
R2014 B.n342 B.n341 10.6151
R2015 B.n342 B.n121 10.6151
R2016 B.n346 B.n121 10.6151
R2017 B.n347 B.n346 10.6151
R2018 B.n348 B.n347 10.6151
R2019 B.n348 B.n119 10.6151
R2020 B.n352 B.n119 10.6151
R2021 B.n353 B.n352 10.6151
R2022 B.n354 B.n353 10.6151
R2023 B.n354 B.n117 10.6151
R2024 B.n358 B.n117 10.6151
R2025 B.n359 B.n358 10.6151
R2026 B.n360 B.n359 10.6151
R2027 B.n360 B.n115 10.6151
R2028 B.n364 B.n115 10.6151
R2029 B.n365 B.n364 10.6151
R2030 B.n366 B.n365 10.6151
R2031 B.n366 B.n113 10.6151
R2032 B.n370 B.n113 10.6151
R2033 B.n371 B.n370 10.6151
R2034 B.n570 B.n569 9.36635
R2035 B.n552 B.n52 9.36635
R2036 B.n295 B.n294 9.36635
R2037 B.n311 B.n131 9.36635
R2038 B.n689 B.n0 8.11757
R2039 B.n689 B.n1 8.11757
R2040 B.n569 B.n568 1.24928
R2041 B.n52 B.n48 1.24928
R2042 B.n296 B.n295 1.24928
R2043 B.n312 B.n311 1.24928
C0 VN VDD2 8.736389f
C1 VN VDD1 0.150532f
C2 VDD2 VDD1 1.4719f
C3 VTAIL VN 8.958269f
C4 VN w_n3190_n3216# 6.48658f
C5 VTAIL VDD2 10.4677f
C6 VN B 0.996745f
C7 VTAIL VDD1 10.4254f
C8 w_n3190_n3216# VDD2 2.40921f
C9 B VDD2 2.06727f
C10 VN VP 6.67006f
C11 w_n3190_n3216# VDD1 2.32174f
C12 B VDD1 1.99141f
C13 VP VDD2 0.445471f
C14 VP VDD1 9.027451f
C15 VTAIL w_n3190_n3216# 2.96921f
C16 VTAIL B 3.07082f
C17 w_n3190_n3216# B 8.51712f
C18 VTAIL VP 8.97267f
C19 w_n3190_n3216# VP 6.89857f
C20 B VP 1.68357f
C21 VDD2 VSUBS 1.708054f
C22 VDD1 VSUBS 1.479807f
C23 VTAIL VSUBS 1.006542f
C24 VN VSUBS 5.93227f
C25 VP VSUBS 2.823187f
C26 B VSUBS 3.961893f
C27 w_n3190_n3216# VSUBS 0.126439p
C28 B.n0 VSUBS 0.0071f
C29 B.n1 VSUBS 0.0071f
C30 B.n2 VSUBS 0.0105f
C31 B.n3 VSUBS 0.008046f
C32 B.n4 VSUBS 0.008046f
C33 B.n5 VSUBS 0.008046f
C34 B.n6 VSUBS 0.008046f
C35 B.n7 VSUBS 0.008046f
C36 B.n8 VSUBS 0.008046f
C37 B.n9 VSUBS 0.008046f
C38 B.n10 VSUBS 0.008046f
C39 B.n11 VSUBS 0.008046f
C40 B.n12 VSUBS 0.008046f
C41 B.n13 VSUBS 0.008046f
C42 B.n14 VSUBS 0.008046f
C43 B.n15 VSUBS 0.008046f
C44 B.n16 VSUBS 0.008046f
C45 B.n17 VSUBS 0.008046f
C46 B.n18 VSUBS 0.008046f
C47 B.n19 VSUBS 0.008046f
C48 B.n20 VSUBS 0.008046f
C49 B.n21 VSUBS 0.008046f
C50 B.n22 VSUBS 0.020931f
C51 B.n23 VSUBS 0.008046f
C52 B.n24 VSUBS 0.008046f
C53 B.n25 VSUBS 0.008046f
C54 B.n26 VSUBS 0.008046f
C55 B.n27 VSUBS 0.008046f
C56 B.n28 VSUBS 0.008046f
C57 B.n29 VSUBS 0.008046f
C58 B.n30 VSUBS 0.008046f
C59 B.n31 VSUBS 0.008046f
C60 B.n32 VSUBS 0.008046f
C61 B.n33 VSUBS 0.008046f
C62 B.n34 VSUBS 0.008046f
C63 B.n35 VSUBS 0.008046f
C64 B.n36 VSUBS 0.008046f
C65 B.n37 VSUBS 0.008046f
C66 B.n38 VSUBS 0.008046f
C67 B.n39 VSUBS 0.008046f
C68 B.n40 VSUBS 0.008046f
C69 B.n41 VSUBS 0.008046f
C70 B.t10 VSUBS 0.223001f
C71 B.t11 VSUBS 0.246538f
C72 B.t9 VSUBS 0.863767f
C73 B.n42 VSUBS 0.383588f
C74 B.n43 VSUBS 0.272313f
C75 B.n44 VSUBS 0.008046f
C76 B.n45 VSUBS 0.008046f
C77 B.n46 VSUBS 0.008046f
C78 B.n47 VSUBS 0.008046f
C79 B.n48 VSUBS 0.004496f
C80 B.n49 VSUBS 0.008046f
C81 B.t1 VSUBS 0.223004f
C82 B.t2 VSUBS 0.246541f
C83 B.t0 VSUBS 0.863767f
C84 B.n50 VSUBS 0.383585f
C85 B.n51 VSUBS 0.27231f
C86 B.n52 VSUBS 0.018642f
C87 B.n53 VSUBS 0.008046f
C88 B.n54 VSUBS 0.008046f
C89 B.n55 VSUBS 0.008046f
C90 B.n56 VSUBS 0.008046f
C91 B.n57 VSUBS 0.008046f
C92 B.n58 VSUBS 0.008046f
C93 B.n59 VSUBS 0.008046f
C94 B.n60 VSUBS 0.008046f
C95 B.n61 VSUBS 0.008046f
C96 B.n62 VSUBS 0.008046f
C97 B.n63 VSUBS 0.008046f
C98 B.n64 VSUBS 0.008046f
C99 B.n65 VSUBS 0.008046f
C100 B.n66 VSUBS 0.008046f
C101 B.n67 VSUBS 0.008046f
C102 B.n68 VSUBS 0.008046f
C103 B.n69 VSUBS 0.008046f
C104 B.n70 VSUBS 0.008046f
C105 B.n71 VSUBS 0.02001f
C106 B.n72 VSUBS 0.008046f
C107 B.n73 VSUBS 0.008046f
C108 B.n74 VSUBS 0.008046f
C109 B.n75 VSUBS 0.008046f
C110 B.n76 VSUBS 0.008046f
C111 B.n77 VSUBS 0.008046f
C112 B.n78 VSUBS 0.008046f
C113 B.n79 VSUBS 0.008046f
C114 B.n80 VSUBS 0.008046f
C115 B.n81 VSUBS 0.008046f
C116 B.n82 VSUBS 0.008046f
C117 B.n83 VSUBS 0.008046f
C118 B.n84 VSUBS 0.008046f
C119 B.n85 VSUBS 0.008046f
C120 B.n86 VSUBS 0.008046f
C121 B.n87 VSUBS 0.008046f
C122 B.n88 VSUBS 0.008046f
C123 B.n89 VSUBS 0.008046f
C124 B.n90 VSUBS 0.008046f
C125 B.n91 VSUBS 0.008046f
C126 B.n92 VSUBS 0.008046f
C127 B.n93 VSUBS 0.008046f
C128 B.n94 VSUBS 0.008046f
C129 B.n95 VSUBS 0.008046f
C130 B.n96 VSUBS 0.008046f
C131 B.n97 VSUBS 0.008046f
C132 B.n98 VSUBS 0.008046f
C133 B.n99 VSUBS 0.008046f
C134 B.n100 VSUBS 0.008046f
C135 B.n101 VSUBS 0.008046f
C136 B.n102 VSUBS 0.008046f
C137 B.n103 VSUBS 0.008046f
C138 B.n104 VSUBS 0.008046f
C139 B.n105 VSUBS 0.008046f
C140 B.n106 VSUBS 0.008046f
C141 B.n107 VSUBS 0.008046f
C142 B.n108 VSUBS 0.008046f
C143 B.n109 VSUBS 0.008046f
C144 B.n110 VSUBS 0.008046f
C145 B.n111 VSUBS 0.008046f
C146 B.n112 VSUBS 0.020931f
C147 B.n113 VSUBS 0.008046f
C148 B.n114 VSUBS 0.008046f
C149 B.n115 VSUBS 0.008046f
C150 B.n116 VSUBS 0.008046f
C151 B.n117 VSUBS 0.008046f
C152 B.n118 VSUBS 0.008046f
C153 B.n119 VSUBS 0.008046f
C154 B.n120 VSUBS 0.008046f
C155 B.n121 VSUBS 0.008046f
C156 B.n122 VSUBS 0.008046f
C157 B.n123 VSUBS 0.008046f
C158 B.n124 VSUBS 0.008046f
C159 B.n125 VSUBS 0.008046f
C160 B.n126 VSUBS 0.008046f
C161 B.n127 VSUBS 0.008046f
C162 B.n128 VSUBS 0.008046f
C163 B.n129 VSUBS 0.008046f
C164 B.n130 VSUBS 0.008046f
C165 B.n131 VSUBS 0.007573f
C166 B.n132 VSUBS 0.008046f
C167 B.n133 VSUBS 0.008046f
C168 B.n134 VSUBS 0.008046f
C169 B.n135 VSUBS 0.008046f
C170 B.n136 VSUBS 0.008046f
C171 B.t8 VSUBS 0.223001f
C172 B.t7 VSUBS 0.246538f
C173 B.t6 VSUBS 0.863767f
C174 B.n137 VSUBS 0.383588f
C175 B.n138 VSUBS 0.272313f
C176 B.n139 VSUBS 0.008046f
C177 B.n140 VSUBS 0.008046f
C178 B.n141 VSUBS 0.008046f
C179 B.n142 VSUBS 0.008046f
C180 B.n143 VSUBS 0.008046f
C181 B.n144 VSUBS 0.008046f
C182 B.n145 VSUBS 0.008046f
C183 B.n146 VSUBS 0.008046f
C184 B.n147 VSUBS 0.008046f
C185 B.n148 VSUBS 0.008046f
C186 B.n149 VSUBS 0.008046f
C187 B.n150 VSUBS 0.008046f
C188 B.n151 VSUBS 0.008046f
C189 B.n152 VSUBS 0.008046f
C190 B.n153 VSUBS 0.008046f
C191 B.n154 VSUBS 0.008046f
C192 B.n155 VSUBS 0.008046f
C193 B.n156 VSUBS 0.008046f
C194 B.n157 VSUBS 0.008046f
C195 B.n158 VSUBS 0.02001f
C196 B.n159 VSUBS 0.008046f
C197 B.n160 VSUBS 0.008046f
C198 B.n161 VSUBS 0.008046f
C199 B.n162 VSUBS 0.008046f
C200 B.n163 VSUBS 0.008046f
C201 B.n164 VSUBS 0.008046f
C202 B.n165 VSUBS 0.008046f
C203 B.n166 VSUBS 0.008046f
C204 B.n167 VSUBS 0.008046f
C205 B.n168 VSUBS 0.008046f
C206 B.n169 VSUBS 0.008046f
C207 B.n170 VSUBS 0.008046f
C208 B.n171 VSUBS 0.008046f
C209 B.n172 VSUBS 0.008046f
C210 B.n173 VSUBS 0.008046f
C211 B.n174 VSUBS 0.008046f
C212 B.n175 VSUBS 0.008046f
C213 B.n176 VSUBS 0.008046f
C214 B.n177 VSUBS 0.008046f
C215 B.n178 VSUBS 0.008046f
C216 B.n179 VSUBS 0.008046f
C217 B.n180 VSUBS 0.008046f
C218 B.n181 VSUBS 0.008046f
C219 B.n182 VSUBS 0.008046f
C220 B.n183 VSUBS 0.008046f
C221 B.n184 VSUBS 0.008046f
C222 B.n185 VSUBS 0.008046f
C223 B.n186 VSUBS 0.008046f
C224 B.n187 VSUBS 0.008046f
C225 B.n188 VSUBS 0.008046f
C226 B.n189 VSUBS 0.008046f
C227 B.n190 VSUBS 0.008046f
C228 B.n191 VSUBS 0.008046f
C229 B.n192 VSUBS 0.008046f
C230 B.n193 VSUBS 0.008046f
C231 B.n194 VSUBS 0.008046f
C232 B.n195 VSUBS 0.008046f
C233 B.n196 VSUBS 0.008046f
C234 B.n197 VSUBS 0.008046f
C235 B.n198 VSUBS 0.008046f
C236 B.n199 VSUBS 0.008046f
C237 B.n200 VSUBS 0.008046f
C238 B.n201 VSUBS 0.008046f
C239 B.n202 VSUBS 0.008046f
C240 B.n203 VSUBS 0.008046f
C241 B.n204 VSUBS 0.008046f
C242 B.n205 VSUBS 0.008046f
C243 B.n206 VSUBS 0.008046f
C244 B.n207 VSUBS 0.008046f
C245 B.n208 VSUBS 0.008046f
C246 B.n209 VSUBS 0.008046f
C247 B.n210 VSUBS 0.008046f
C248 B.n211 VSUBS 0.008046f
C249 B.n212 VSUBS 0.008046f
C250 B.n213 VSUBS 0.008046f
C251 B.n214 VSUBS 0.008046f
C252 B.n215 VSUBS 0.008046f
C253 B.n216 VSUBS 0.008046f
C254 B.n217 VSUBS 0.008046f
C255 B.n218 VSUBS 0.008046f
C256 B.n219 VSUBS 0.008046f
C257 B.n220 VSUBS 0.008046f
C258 B.n221 VSUBS 0.008046f
C259 B.n222 VSUBS 0.008046f
C260 B.n223 VSUBS 0.008046f
C261 B.n224 VSUBS 0.008046f
C262 B.n225 VSUBS 0.008046f
C263 B.n226 VSUBS 0.008046f
C264 B.n227 VSUBS 0.008046f
C265 B.n228 VSUBS 0.008046f
C266 B.n229 VSUBS 0.008046f
C267 B.n230 VSUBS 0.008046f
C268 B.n231 VSUBS 0.008046f
C269 B.n232 VSUBS 0.008046f
C270 B.n233 VSUBS 0.008046f
C271 B.n234 VSUBS 0.008046f
C272 B.n235 VSUBS 0.02001f
C273 B.n236 VSUBS 0.020931f
C274 B.n237 VSUBS 0.020931f
C275 B.n238 VSUBS 0.008046f
C276 B.n239 VSUBS 0.008046f
C277 B.n240 VSUBS 0.008046f
C278 B.n241 VSUBS 0.008046f
C279 B.n242 VSUBS 0.008046f
C280 B.n243 VSUBS 0.008046f
C281 B.n244 VSUBS 0.008046f
C282 B.n245 VSUBS 0.008046f
C283 B.n246 VSUBS 0.008046f
C284 B.n247 VSUBS 0.008046f
C285 B.n248 VSUBS 0.008046f
C286 B.n249 VSUBS 0.008046f
C287 B.n250 VSUBS 0.008046f
C288 B.n251 VSUBS 0.008046f
C289 B.n252 VSUBS 0.008046f
C290 B.n253 VSUBS 0.008046f
C291 B.n254 VSUBS 0.008046f
C292 B.n255 VSUBS 0.008046f
C293 B.n256 VSUBS 0.008046f
C294 B.n257 VSUBS 0.008046f
C295 B.n258 VSUBS 0.008046f
C296 B.n259 VSUBS 0.008046f
C297 B.n260 VSUBS 0.008046f
C298 B.n261 VSUBS 0.008046f
C299 B.n262 VSUBS 0.008046f
C300 B.n263 VSUBS 0.008046f
C301 B.n264 VSUBS 0.008046f
C302 B.n265 VSUBS 0.008046f
C303 B.n266 VSUBS 0.008046f
C304 B.n267 VSUBS 0.008046f
C305 B.n268 VSUBS 0.008046f
C306 B.n269 VSUBS 0.008046f
C307 B.n270 VSUBS 0.008046f
C308 B.n271 VSUBS 0.008046f
C309 B.n272 VSUBS 0.008046f
C310 B.n273 VSUBS 0.008046f
C311 B.n274 VSUBS 0.008046f
C312 B.n275 VSUBS 0.008046f
C313 B.n276 VSUBS 0.008046f
C314 B.n277 VSUBS 0.008046f
C315 B.n278 VSUBS 0.008046f
C316 B.n279 VSUBS 0.008046f
C317 B.n280 VSUBS 0.008046f
C318 B.n281 VSUBS 0.008046f
C319 B.n282 VSUBS 0.008046f
C320 B.n283 VSUBS 0.008046f
C321 B.n284 VSUBS 0.008046f
C322 B.n285 VSUBS 0.008046f
C323 B.n286 VSUBS 0.008046f
C324 B.n287 VSUBS 0.008046f
C325 B.n288 VSUBS 0.008046f
C326 B.n289 VSUBS 0.008046f
C327 B.n290 VSUBS 0.008046f
C328 B.n291 VSUBS 0.008046f
C329 B.n292 VSUBS 0.008046f
C330 B.n293 VSUBS 0.008046f
C331 B.n294 VSUBS 0.007573f
C332 B.n295 VSUBS 0.018642f
C333 B.n296 VSUBS 0.004496f
C334 B.n297 VSUBS 0.008046f
C335 B.n298 VSUBS 0.008046f
C336 B.n299 VSUBS 0.008046f
C337 B.n300 VSUBS 0.008046f
C338 B.n301 VSUBS 0.008046f
C339 B.n302 VSUBS 0.008046f
C340 B.n303 VSUBS 0.008046f
C341 B.n304 VSUBS 0.008046f
C342 B.n305 VSUBS 0.008046f
C343 B.n306 VSUBS 0.008046f
C344 B.n307 VSUBS 0.008046f
C345 B.n308 VSUBS 0.008046f
C346 B.t5 VSUBS 0.223004f
C347 B.t4 VSUBS 0.246541f
C348 B.t3 VSUBS 0.863767f
C349 B.n309 VSUBS 0.383585f
C350 B.n310 VSUBS 0.27231f
C351 B.n311 VSUBS 0.018642f
C352 B.n312 VSUBS 0.004496f
C353 B.n313 VSUBS 0.008046f
C354 B.n314 VSUBS 0.008046f
C355 B.n315 VSUBS 0.008046f
C356 B.n316 VSUBS 0.008046f
C357 B.n317 VSUBS 0.008046f
C358 B.n318 VSUBS 0.008046f
C359 B.n319 VSUBS 0.008046f
C360 B.n320 VSUBS 0.008046f
C361 B.n321 VSUBS 0.008046f
C362 B.n322 VSUBS 0.008046f
C363 B.n323 VSUBS 0.008046f
C364 B.n324 VSUBS 0.008046f
C365 B.n325 VSUBS 0.008046f
C366 B.n326 VSUBS 0.008046f
C367 B.n327 VSUBS 0.008046f
C368 B.n328 VSUBS 0.008046f
C369 B.n329 VSUBS 0.008046f
C370 B.n330 VSUBS 0.008046f
C371 B.n331 VSUBS 0.008046f
C372 B.n332 VSUBS 0.008046f
C373 B.n333 VSUBS 0.008046f
C374 B.n334 VSUBS 0.008046f
C375 B.n335 VSUBS 0.008046f
C376 B.n336 VSUBS 0.008046f
C377 B.n337 VSUBS 0.008046f
C378 B.n338 VSUBS 0.008046f
C379 B.n339 VSUBS 0.008046f
C380 B.n340 VSUBS 0.008046f
C381 B.n341 VSUBS 0.008046f
C382 B.n342 VSUBS 0.008046f
C383 B.n343 VSUBS 0.008046f
C384 B.n344 VSUBS 0.008046f
C385 B.n345 VSUBS 0.008046f
C386 B.n346 VSUBS 0.008046f
C387 B.n347 VSUBS 0.008046f
C388 B.n348 VSUBS 0.008046f
C389 B.n349 VSUBS 0.008046f
C390 B.n350 VSUBS 0.008046f
C391 B.n351 VSUBS 0.008046f
C392 B.n352 VSUBS 0.008046f
C393 B.n353 VSUBS 0.008046f
C394 B.n354 VSUBS 0.008046f
C395 B.n355 VSUBS 0.008046f
C396 B.n356 VSUBS 0.008046f
C397 B.n357 VSUBS 0.008046f
C398 B.n358 VSUBS 0.008046f
C399 B.n359 VSUBS 0.008046f
C400 B.n360 VSUBS 0.008046f
C401 B.n361 VSUBS 0.008046f
C402 B.n362 VSUBS 0.008046f
C403 B.n363 VSUBS 0.008046f
C404 B.n364 VSUBS 0.008046f
C405 B.n365 VSUBS 0.008046f
C406 B.n366 VSUBS 0.008046f
C407 B.n367 VSUBS 0.008046f
C408 B.n368 VSUBS 0.008046f
C409 B.n369 VSUBS 0.008046f
C410 B.n370 VSUBS 0.008046f
C411 B.n371 VSUBS 0.020092f
C412 B.n372 VSUBS 0.020849f
C413 B.n373 VSUBS 0.02001f
C414 B.n374 VSUBS 0.008046f
C415 B.n375 VSUBS 0.008046f
C416 B.n376 VSUBS 0.008046f
C417 B.n377 VSUBS 0.008046f
C418 B.n378 VSUBS 0.008046f
C419 B.n379 VSUBS 0.008046f
C420 B.n380 VSUBS 0.008046f
C421 B.n381 VSUBS 0.008046f
C422 B.n382 VSUBS 0.008046f
C423 B.n383 VSUBS 0.008046f
C424 B.n384 VSUBS 0.008046f
C425 B.n385 VSUBS 0.008046f
C426 B.n386 VSUBS 0.008046f
C427 B.n387 VSUBS 0.008046f
C428 B.n388 VSUBS 0.008046f
C429 B.n389 VSUBS 0.008046f
C430 B.n390 VSUBS 0.008046f
C431 B.n391 VSUBS 0.008046f
C432 B.n392 VSUBS 0.008046f
C433 B.n393 VSUBS 0.008046f
C434 B.n394 VSUBS 0.008046f
C435 B.n395 VSUBS 0.008046f
C436 B.n396 VSUBS 0.008046f
C437 B.n397 VSUBS 0.008046f
C438 B.n398 VSUBS 0.008046f
C439 B.n399 VSUBS 0.008046f
C440 B.n400 VSUBS 0.008046f
C441 B.n401 VSUBS 0.008046f
C442 B.n402 VSUBS 0.008046f
C443 B.n403 VSUBS 0.008046f
C444 B.n404 VSUBS 0.008046f
C445 B.n405 VSUBS 0.008046f
C446 B.n406 VSUBS 0.008046f
C447 B.n407 VSUBS 0.008046f
C448 B.n408 VSUBS 0.008046f
C449 B.n409 VSUBS 0.008046f
C450 B.n410 VSUBS 0.008046f
C451 B.n411 VSUBS 0.008046f
C452 B.n412 VSUBS 0.008046f
C453 B.n413 VSUBS 0.008046f
C454 B.n414 VSUBS 0.008046f
C455 B.n415 VSUBS 0.008046f
C456 B.n416 VSUBS 0.008046f
C457 B.n417 VSUBS 0.008046f
C458 B.n418 VSUBS 0.008046f
C459 B.n419 VSUBS 0.008046f
C460 B.n420 VSUBS 0.008046f
C461 B.n421 VSUBS 0.008046f
C462 B.n422 VSUBS 0.008046f
C463 B.n423 VSUBS 0.008046f
C464 B.n424 VSUBS 0.008046f
C465 B.n425 VSUBS 0.008046f
C466 B.n426 VSUBS 0.008046f
C467 B.n427 VSUBS 0.008046f
C468 B.n428 VSUBS 0.008046f
C469 B.n429 VSUBS 0.008046f
C470 B.n430 VSUBS 0.008046f
C471 B.n431 VSUBS 0.008046f
C472 B.n432 VSUBS 0.008046f
C473 B.n433 VSUBS 0.008046f
C474 B.n434 VSUBS 0.008046f
C475 B.n435 VSUBS 0.008046f
C476 B.n436 VSUBS 0.008046f
C477 B.n437 VSUBS 0.008046f
C478 B.n438 VSUBS 0.008046f
C479 B.n439 VSUBS 0.008046f
C480 B.n440 VSUBS 0.008046f
C481 B.n441 VSUBS 0.008046f
C482 B.n442 VSUBS 0.008046f
C483 B.n443 VSUBS 0.008046f
C484 B.n444 VSUBS 0.008046f
C485 B.n445 VSUBS 0.008046f
C486 B.n446 VSUBS 0.008046f
C487 B.n447 VSUBS 0.008046f
C488 B.n448 VSUBS 0.008046f
C489 B.n449 VSUBS 0.008046f
C490 B.n450 VSUBS 0.008046f
C491 B.n451 VSUBS 0.008046f
C492 B.n452 VSUBS 0.008046f
C493 B.n453 VSUBS 0.008046f
C494 B.n454 VSUBS 0.008046f
C495 B.n455 VSUBS 0.008046f
C496 B.n456 VSUBS 0.008046f
C497 B.n457 VSUBS 0.008046f
C498 B.n458 VSUBS 0.008046f
C499 B.n459 VSUBS 0.008046f
C500 B.n460 VSUBS 0.008046f
C501 B.n461 VSUBS 0.008046f
C502 B.n462 VSUBS 0.008046f
C503 B.n463 VSUBS 0.008046f
C504 B.n464 VSUBS 0.008046f
C505 B.n465 VSUBS 0.008046f
C506 B.n466 VSUBS 0.008046f
C507 B.n467 VSUBS 0.008046f
C508 B.n468 VSUBS 0.008046f
C509 B.n469 VSUBS 0.008046f
C510 B.n470 VSUBS 0.008046f
C511 B.n471 VSUBS 0.008046f
C512 B.n472 VSUBS 0.008046f
C513 B.n473 VSUBS 0.008046f
C514 B.n474 VSUBS 0.008046f
C515 B.n475 VSUBS 0.008046f
C516 B.n476 VSUBS 0.008046f
C517 B.n477 VSUBS 0.008046f
C518 B.n478 VSUBS 0.008046f
C519 B.n479 VSUBS 0.008046f
C520 B.n480 VSUBS 0.008046f
C521 B.n481 VSUBS 0.008046f
C522 B.n482 VSUBS 0.008046f
C523 B.n483 VSUBS 0.008046f
C524 B.n484 VSUBS 0.008046f
C525 B.n485 VSUBS 0.008046f
C526 B.n486 VSUBS 0.008046f
C527 B.n487 VSUBS 0.008046f
C528 B.n488 VSUBS 0.008046f
C529 B.n489 VSUBS 0.008046f
C530 B.n490 VSUBS 0.008046f
C531 B.n491 VSUBS 0.008046f
C532 B.n492 VSUBS 0.008046f
C533 B.n493 VSUBS 0.008046f
C534 B.n494 VSUBS 0.02001f
C535 B.n495 VSUBS 0.020931f
C536 B.n496 VSUBS 0.020931f
C537 B.n497 VSUBS 0.008046f
C538 B.n498 VSUBS 0.008046f
C539 B.n499 VSUBS 0.008046f
C540 B.n500 VSUBS 0.008046f
C541 B.n501 VSUBS 0.008046f
C542 B.n502 VSUBS 0.008046f
C543 B.n503 VSUBS 0.008046f
C544 B.n504 VSUBS 0.008046f
C545 B.n505 VSUBS 0.008046f
C546 B.n506 VSUBS 0.008046f
C547 B.n507 VSUBS 0.008046f
C548 B.n508 VSUBS 0.008046f
C549 B.n509 VSUBS 0.008046f
C550 B.n510 VSUBS 0.008046f
C551 B.n511 VSUBS 0.008046f
C552 B.n512 VSUBS 0.008046f
C553 B.n513 VSUBS 0.008046f
C554 B.n514 VSUBS 0.008046f
C555 B.n515 VSUBS 0.008046f
C556 B.n516 VSUBS 0.008046f
C557 B.n517 VSUBS 0.008046f
C558 B.n518 VSUBS 0.008046f
C559 B.n519 VSUBS 0.008046f
C560 B.n520 VSUBS 0.008046f
C561 B.n521 VSUBS 0.008046f
C562 B.n522 VSUBS 0.008046f
C563 B.n523 VSUBS 0.008046f
C564 B.n524 VSUBS 0.008046f
C565 B.n525 VSUBS 0.008046f
C566 B.n526 VSUBS 0.008046f
C567 B.n527 VSUBS 0.008046f
C568 B.n528 VSUBS 0.008046f
C569 B.n529 VSUBS 0.008046f
C570 B.n530 VSUBS 0.008046f
C571 B.n531 VSUBS 0.008046f
C572 B.n532 VSUBS 0.008046f
C573 B.n533 VSUBS 0.008046f
C574 B.n534 VSUBS 0.008046f
C575 B.n535 VSUBS 0.008046f
C576 B.n536 VSUBS 0.008046f
C577 B.n537 VSUBS 0.008046f
C578 B.n538 VSUBS 0.008046f
C579 B.n539 VSUBS 0.008046f
C580 B.n540 VSUBS 0.008046f
C581 B.n541 VSUBS 0.008046f
C582 B.n542 VSUBS 0.008046f
C583 B.n543 VSUBS 0.008046f
C584 B.n544 VSUBS 0.008046f
C585 B.n545 VSUBS 0.008046f
C586 B.n546 VSUBS 0.008046f
C587 B.n547 VSUBS 0.008046f
C588 B.n548 VSUBS 0.008046f
C589 B.n549 VSUBS 0.008046f
C590 B.n550 VSUBS 0.008046f
C591 B.n551 VSUBS 0.008046f
C592 B.n552 VSUBS 0.007573f
C593 B.n553 VSUBS 0.008046f
C594 B.n554 VSUBS 0.008046f
C595 B.n555 VSUBS 0.008046f
C596 B.n556 VSUBS 0.008046f
C597 B.n557 VSUBS 0.008046f
C598 B.n558 VSUBS 0.008046f
C599 B.n559 VSUBS 0.008046f
C600 B.n560 VSUBS 0.008046f
C601 B.n561 VSUBS 0.008046f
C602 B.n562 VSUBS 0.008046f
C603 B.n563 VSUBS 0.008046f
C604 B.n564 VSUBS 0.008046f
C605 B.n565 VSUBS 0.008046f
C606 B.n566 VSUBS 0.008046f
C607 B.n567 VSUBS 0.008046f
C608 B.n568 VSUBS 0.004496f
C609 B.n569 VSUBS 0.018642f
C610 B.n570 VSUBS 0.007573f
C611 B.n571 VSUBS 0.008046f
C612 B.n572 VSUBS 0.008046f
C613 B.n573 VSUBS 0.008046f
C614 B.n574 VSUBS 0.008046f
C615 B.n575 VSUBS 0.008046f
C616 B.n576 VSUBS 0.008046f
C617 B.n577 VSUBS 0.008046f
C618 B.n578 VSUBS 0.008046f
C619 B.n579 VSUBS 0.008046f
C620 B.n580 VSUBS 0.008046f
C621 B.n581 VSUBS 0.008046f
C622 B.n582 VSUBS 0.008046f
C623 B.n583 VSUBS 0.008046f
C624 B.n584 VSUBS 0.008046f
C625 B.n585 VSUBS 0.008046f
C626 B.n586 VSUBS 0.008046f
C627 B.n587 VSUBS 0.008046f
C628 B.n588 VSUBS 0.008046f
C629 B.n589 VSUBS 0.008046f
C630 B.n590 VSUBS 0.008046f
C631 B.n591 VSUBS 0.008046f
C632 B.n592 VSUBS 0.008046f
C633 B.n593 VSUBS 0.008046f
C634 B.n594 VSUBS 0.008046f
C635 B.n595 VSUBS 0.008046f
C636 B.n596 VSUBS 0.008046f
C637 B.n597 VSUBS 0.008046f
C638 B.n598 VSUBS 0.008046f
C639 B.n599 VSUBS 0.008046f
C640 B.n600 VSUBS 0.008046f
C641 B.n601 VSUBS 0.008046f
C642 B.n602 VSUBS 0.008046f
C643 B.n603 VSUBS 0.008046f
C644 B.n604 VSUBS 0.008046f
C645 B.n605 VSUBS 0.008046f
C646 B.n606 VSUBS 0.008046f
C647 B.n607 VSUBS 0.008046f
C648 B.n608 VSUBS 0.008046f
C649 B.n609 VSUBS 0.008046f
C650 B.n610 VSUBS 0.008046f
C651 B.n611 VSUBS 0.008046f
C652 B.n612 VSUBS 0.008046f
C653 B.n613 VSUBS 0.008046f
C654 B.n614 VSUBS 0.008046f
C655 B.n615 VSUBS 0.008046f
C656 B.n616 VSUBS 0.008046f
C657 B.n617 VSUBS 0.008046f
C658 B.n618 VSUBS 0.008046f
C659 B.n619 VSUBS 0.008046f
C660 B.n620 VSUBS 0.008046f
C661 B.n621 VSUBS 0.008046f
C662 B.n622 VSUBS 0.008046f
C663 B.n623 VSUBS 0.008046f
C664 B.n624 VSUBS 0.008046f
C665 B.n625 VSUBS 0.008046f
C666 B.n626 VSUBS 0.008046f
C667 B.n627 VSUBS 0.020931f
C668 B.n628 VSUBS 0.02001f
C669 B.n629 VSUBS 0.02001f
C670 B.n630 VSUBS 0.008046f
C671 B.n631 VSUBS 0.008046f
C672 B.n632 VSUBS 0.008046f
C673 B.n633 VSUBS 0.008046f
C674 B.n634 VSUBS 0.008046f
C675 B.n635 VSUBS 0.008046f
C676 B.n636 VSUBS 0.008046f
C677 B.n637 VSUBS 0.008046f
C678 B.n638 VSUBS 0.008046f
C679 B.n639 VSUBS 0.008046f
C680 B.n640 VSUBS 0.008046f
C681 B.n641 VSUBS 0.008046f
C682 B.n642 VSUBS 0.008046f
C683 B.n643 VSUBS 0.008046f
C684 B.n644 VSUBS 0.008046f
C685 B.n645 VSUBS 0.008046f
C686 B.n646 VSUBS 0.008046f
C687 B.n647 VSUBS 0.008046f
C688 B.n648 VSUBS 0.008046f
C689 B.n649 VSUBS 0.008046f
C690 B.n650 VSUBS 0.008046f
C691 B.n651 VSUBS 0.008046f
C692 B.n652 VSUBS 0.008046f
C693 B.n653 VSUBS 0.008046f
C694 B.n654 VSUBS 0.008046f
C695 B.n655 VSUBS 0.008046f
C696 B.n656 VSUBS 0.008046f
C697 B.n657 VSUBS 0.008046f
C698 B.n658 VSUBS 0.008046f
C699 B.n659 VSUBS 0.008046f
C700 B.n660 VSUBS 0.008046f
C701 B.n661 VSUBS 0.008046f
C702 B.n662 VSUBS 0.008046f
C703 B.n663 VSUBS 0.008046f
C704 B.n664 VSUBS 0.008046f
C705 B.n665 VSUBS 0.008046f
C706 B.n666 VSUBS 0.008046f
C707 B.n667 VSUBS 0.008046f
C708 B.n668 VSUBS 0.008046f
C709 B.n669 VSUBS 0.008046f
C710 B.n670 VSUBS 0.008046f
C711 B.n671 VSUBS 0.008046f
C712 B.n672 VSUBS 0.008046f
C713 B.n673 VSUBS 0.008046f
C714 B.n674 VSUBS 0.008046f
C715 B.n675 VSUBS 0.008046f
C716 B.n676 VSUBS 0.008046f
C717 B.n677 VSUBS 0.008046f
C718 B.n678 VSUBS 0.008046f
C719 B.n679 VSUBS 0.008046f
C720 B.n680 VSUBS 0.008046f
C721 B.n681 VSUBS 0.008046f
C722 B.n682 VSUBS 0.008046f
C723 B.n683 VSUBS 0.008046f
C724 B.n684 VSUBS 0.008046f
C725 B.n685 VSUBS 0.008046f
C726 B.n686 VSUBS 0.008046f
C727 B.n687 VSUBS 0.0105f
C728 B.n688 VSUBS 0.011185f
C729 B.n689 VSUBS 0.022243f
C730 VDD1.n0 VSUBS 0.014274f
C731 VDD1.n1 VSUBS 0.032157f
C732 VDD1.n2 VSUBS 0.014405f
C733 VDD1.n3 VSUBS 0.025318f
C734 VDD1.n4 VSUBS 0.013605f
C735 VDD1.n5 VSUBS 0.032157f
C736 VDD1.n6 VSUBS 0.014405f
C737 VDD1.n7 VSUBS 0.025318f
C738 VDD1.n8 VSUBS 0.013605f
C739 VDD1.n9 VSUBS 0.032157f
C740 VDD1.n10 VSUBS 0.014405f
C741 VDD1.n11 VSUBS 0.025318f
C742 VDD1.n12 VSUBS 0.013605f
C743 VDD1.n13 VSUBS 0.032157f
C744 VDD1.n14 VSUBS 0.014405f
C745 VDD1.n15 VSUBS 0.025318f
C746 VDD1.n16 VSUBS 0.013605f
C747 VDD1.n17 VSUBS 0.032157f
C748 VDD1.n18 VSUBS 0.014405f
C749 VDD1.n19 VSUBS 0.150399f
C750 VDD1.t8 VSUBS 0.068612f
C751 VDD1.n20 VSUBS 0.024118f
C752 VDD1.n21 VSUBS 0.020457f
C753 VDD1.n22 VSUBS 0.013605f
C754 VDD1.n23 VSUBS 1.18444f
C755 VDD1.n24 VSUBS 0.025318f
C756 VDD1.n25 VSUBS 0.013605f
C757 VDD1.n26 VSUBS 0.014405f
C758 VDD1.n27 VSUBS 0.032157f
C759 VDD1.n28 VSUBS 0.032157f
C760 VDD1.n29 VSUBS 0.014405f
C761 VDD1.n30 VSUBS 0.013605f
C762 VDD1.n31 VSUBS 0.025318f
C763 VDD1.n32 VSUBS 0.025318f
C764 VDD1.n33 VSUBS 0.013605f
C765 VDD1.n34 VSUBS 0.014405f
C766 VDD1.n35 VSUBS 0.032157f
C767 VDD1.n36 VSUBS 0.032157f
C768 VDD1.n37 VSUBS 0.014405f
C769 VDD1.n38 VSUBS 0.013605f
C770 VDD1.n39 VSUBS 0.025318f
C771 VDD1.n40 VSUBS 0.025318f
C772 VDD1.n41 VSUBS 0.013605f
C773 VDD1.n42 VSUBS 0.014405f
C774 VDD1.n43 VSUBS 0.032157f
C775 VDD1.n44 VSUBS 0.032157f
C776 VDD1.n45 VSUBS 0.014405f
C777 VDD1.n46 VSUBS 0.013605f
C778 VDD1.n47 VSUBS 0.025318f
C779 VDD1.n48 VSUBS 0.025318f
C780 VDD1.n49 VSUBS 0.013605f
C781 VDD1.n50 VSUBS 0.014405f
C782 VDD1.n51 VSUBS 0.032157f
C783 VDD1.n52 VSUBS 0.032157f
C784 VDD1.n53 VSUBS 0.014405f
C785 VDD1.n54 VSUBS 0.013605f
C786 VDD1.n55 VSUBS 0.025318f
C787 VDD1.n56 VSUBS 0.065439f
C788 VDD1.n57 VSUBS 0.013605f
C789 VDD1.n58 VSUBS 0.014405f
C790 VDD1.n59 VSUBS 0.070177f
C791 VDD1.n60 VSUBS 0.070565f
C792 VDD1.t3 VSUBS 0.224881f
C793 VDD1.t0 VSUBS 0.224881f
C794 VDD1.n61 VSUBS 1.7581f
C795 VDD1.n62 VSUBS 0.788819f
C796 VDD1.n63 VSUBS 0.014274f
C797 VDD1.n64 VSUBS 0.032157f
C798 VDD1.n65 VSUBS 0.014405f
C799 VDD1.n66 VSUBS 0.025318f
C800 VDD1.n67 VSUBS 0.013605f
C801 VDD1.n68 VSUBS 0.032157f
C802 VDD1.n69 VSUBS 0.014405f
C803 VDD1.n70 VSUBS 0.025318f
C804 VDD1.n71 VSUBS 0.013605f
C805 VDD1.n72 VSUBS 0.032157f
C806 VDD1.n73 VSUBS 0.014405f
C807 VDD1.n74 VSUBS 0.025318f
C808 VDD1.n75 VSUBS 0.013605f
C809 VDD1.n76 VSUBS 0.032157f
C810 VDD1.n77 VSUBS 0.014405f
C811 VDD1.n78 VSUBS 0.025318f
C812 VDD1.n79 VSUBS 0.013605f
C813 VDD1.n80 VSUBS 0.032157f
C814 VDD1.n81 VSUBS 0.014405f
C815 VDD1.n82 VSUBS 0.150399f
C816 VDD1.t2 VSUBS 0.068612f
C817 VDD1.n83 VSUBS 0.024118f
C818 VDD1.n84 VSUBS 0.020457f
C819 VDD1.n85 VSUBS 0.013605f
C820 VDD1.n86 VSUBS 1.18444f
C821 VDD1.n87 VSUBS 0.025318f
C822 VDD1.n88 VSUBS 0.013605f
C823 VDD1.n89 VSUBS 0.014405f
C824 VDD1.n90 VSUBS 0.032157f
C825 VDD1.n91 VSUBS 0.032157f
C826 VDD1.n92 VSUBS 0.014405f
C827 VDD1.n93 VSUBS 0.013605f
C828 VDD1.n94 VSUBS 0.025318f
C829 VDD1.n95 VSUBS 0.025318f
C830 VDD1.n96 VSUBS 0.013605f
C831 VDD1.n97 VSUBS 0.014405f
C832 VDD1.n98 VSUBS 0.032157f
C833 VDD1.n99 VSUBS 0.032157f
C834 VDD1.n100 VSUBS 0.014405f
C835 VDD1.n101 VSUBS 0.013605f
C836 VDD1.n102 VSUBS 0.025318f
C837 VDD1.n103 VSUBS 0.025318f
C838 VDD1.n104 VSUBS 0.013605f
C839 VDD1.n105 VSUBS 0.014405f
C840 VDD1.n106 VSUBS 0.032157f
C841 VDD1.n107 VSUBS 0.032157f
C842 VDD1.n108 VSUBS 0.014405f
C843 VDD1.n109 VSUBS 0.013605f
C844 VDD1.n110 VSUBS 0.025318f
C845 VDD1.n111 VSUBS 0.025318f
C846 VDD1.n112 VSUBS 0.013605f
C847 VDD1.n113 VSUBS 0.014405f
C848 VDD1.n114 VSUBS 0.032157f
C849 VDD1.n115 VSUBS 0.032157f
C850 VDD1.n116 VSUBS 0.014405f
C851 VDD1.n117 VSUBS 0.013605f
C852 VDD1.n118 VSUBS 0.025318f
C853 VDD1.n119 VSUBS 0.065439f
C854 VDD1.n120 VSUBS 0.013605f
C855 VDD1.n121 VSUBS 0.014405f
C856 VDD1.n122 VSUBS 0.070177f
C857 VDD1.n123 VSUBS 0.070565f
C858 VDD1.t5 VSUBS 0.224881f
C859 VDD1.t6 VSUBS 0.224881f
C860 VDD1.n124 VSUBS 1.75809f
C861 VDD1.n125 VSUBS 0.781273f
C862 VDD1.t7 VSUBS 0.224881f
C863 VDD1.t1 VSUBS 0.224881f
C864 VDD1.n126 VSUBS 1.76787f
C865 VDD1.n127 VSUBS 2.65483f
C866 VDD1.t4 VSUBS 0.224881f
C867 VDD1.t9 VSUBS 0.224881f
C868 VDD1.n128 VSUBS 1.75809f
C869 VDD1.n129 VSUBS 2.9388f
C870 VP.n0 VSUBS 0.038756f
C871 VP.t8 VSUBS 1.80058f
C872 VP.n1 VSUBS 0.059542f
C873 VP.n2 VSUBS 0.038756f
C874 VP.t2 VSUBS 1.80058f
C875 VP.n3 VSUBS 0.073295f
C876 VP.n4 VSUBS 0.038756f
C877 VP.t3 VSUBS 1.80058f
C878 VP.n5 VSUBS 0.067912f
C879 VP.n6 VSUBS 0.038756f
C880 VP.n7 VSUBS 0.051088f
C881 VP.n8 VSUBS 0.038756f
C882 VP.t0 VSUBS 1.80058f
C883 VP.n9 VSUBS 0.059542f
C884 VP.n10 VSUBS 0.038756f
C885 VP.t5 VSUBS 1.80058f
C886 VP.n11 VSUBS 0.073295f
C887 VP.n12 VSUBS 0.038756f
C888 VP.t9 VSUBS 1.80058f
C889 VP.n13 VSUBS 0.067912f
C890 VP.t1 VSUBS 1.9284f
C891 VP.t6 VSUBS 1.80058f
C892 VP.n14 VSUBS 0.73463f
C893 VP.n15 VSUBS 0.743747f
C894 VP.n16 VSUBS 0.245724f
C895 VP.n17 VSUBS 0.038756f
C896 VP.n18 VSUBS 0.034278f
C897 VP.n19 VSUBS 0.073295f
C898 VP.n20 VSUBS 0.691129f
C899 VP.n21 VSUBS 0.038756f
C900 VP.n22 VSUBS 0.038756f
C901 VP.n23 VSUBS 0.038756f
C902 VP.n24 VSUBS 0.034278f
C903 VP.n25 VSUBS 0.067912f
C904 VP.n26 VSUBS 0.654378f
C905 VP.n27 VSUBS 0.047504f
C906 VP.n28 VSUBS 0.038756f
C907 VP.n29 VSUBS 0.038756f
C908 VP.n30 VSUBS 0.038756f
C909 VP.n31 VSUBS 0.054104f
C910 VP.n32 VSUBS 0.051088f
C911 VP.n33 VSUBS 0.735404f
C912 VP.n34 VSUBS 1.8986f
C913 VP.t7 VSUBS 1.80058f
C914 VP.n35 VSUBS 0.735404f
C915 VP.n36 VSUBS 1.92842f
C916 VP.n37 VSUBS 0.038756f
C917 VP.n38 VSUBS 0.038756f
C918 VP.n39 VSUBS 0.054104f
C919 VP.n40 VSUBS 0.059542f
C920 VP.t4 VSUBS 1.80058f
C921 VP.n41 VSUBS 0.654378f
C922 VP.n42 VSUBS 0.047504f
C923 VP.n43 VSUBS 0.038756f
C924 VP.n44 VSUBS 0.038756f
C925 VP.n45 VSUBS 0.038756f
C926 VP.n46 VSUBS 0.034278f
C927 VP.n47 VSUBS 0.073295f
C928 VP.n48 VSUBS 0.691129f
C929 VP.n49 VSUBS 0.038756f
C930 VP.n50 VSUBS 0.038756f
C931 VP.n51 VSUBS 0.038756f
C932 VP.n52 VSUBS 0.034278f
C933 VP.n53 VSUBS 0.067912f
C934 VP.n54 VSUBS 0.654378f
C935 VP.n55 VSUBS 0.047504f
C936 VP.n56 VSUBS 0.038756f
C937 VP.n57 VSUBS 0.038756f
C938 VP.n58 VSUBS 0.038756f
C939 VP.n59 VSUBS 0.054104f
C940 VP.n60 VSUBS 0.051088f
C941 VP.n61 VSUBS 0.735404f
C942 VP.n62 VSUBS 0.037371f
C943 VTAIL.t11 VSUBS 0.25361f
C944 VTAIL.t16 VSUBS 0.25361f
C945 VTAIL.n0 VSUBS 1.84769f
C946 VTAIL.n1 VSUBS 0.831285f
C947 VTAIL.n2 VSUBS 0.016098f
C948 VTAIL.n3 VSUBS 0.036265f
C949 VTAIL.n4 VSUBS 0.016246f
C950 VTAIL.n5 VSUBS 0.028553f
C951 VTAIL.n6 VSUBS 0.015343f
C952 VTAIL.n7 VSUBS 0.036265f
C953 VTAIL.n8 VSUBS 0.016246f
C954 VTAIL.n9 VSUBS 0.028553f
C955 VTAIL.n10 VSUBS 0.015343f
C956 VTAIL.n11 VSUBS 0.036265f
C957 VTAIL.n12 VSUBS 0.016246f
C958 VTAIL.n13 VSUBS 0.028553f
C959 VTAIL.n14 VSUBS 0.015343f
C960 VTAIL.n15 VSUBS 0.036265f
C961 VTAIL.n16 VSUBS 0.016246f
C962 VTAIL.n17 VSUBS 0.028553f
C963 VTAIL.n18 VSUBS 0.015343f
C964 VTAIL.n19 VSUBS 0.036265f
C965 VTAIL.n20 VSUBS 0.016246f
C966 VTAIL.n21 VSUBS 0.169613f
C967 VTAIL.t3 VSUBS 0.077377f
C968 VTAIL.n22 VSUBS 0.027199f
C969 VTAIL.n23 VSUBS 0.02307f
C970 VTAIL.n24 VSUBS 0.015343f
C971 VTAIL.n25 VSUBS 1.33576f
C972 VTAIL.n26 VSUBS 0.028553f
C973 VTAIL.n27 VSUBS 0.015343f
C974 VTAIL.n28 VSUBS 0.016246f
C975 VTAIL.n29 VSUBS 0.036265f
C976 VTAIL.n30 VSUBS 0.036265f
C977 VTAIL.n31 VSUBS 0.016246f
C978 VTAIL.n32 VSUBS 0.015343f
C979 VTAIL.n33 VSUBS 0.028553f
C980 VTAIL.n34 VSUBS 0.028553f
C981 VTAIL.n35 VSUBS 0.015343f
C982 VTAIL.n36 VSUBS 0.016246f
C983 VTAIL.n37 VSUBS 0.036265f
C984 VTAIL.n38 VSUBS 0.036265f
C985 VTAIL.n39 VSUBS 0.016246f
C986 VTAIL.n40 VSUBS 0.015343f
C987 VTAIL.n41 VSUBS 0.028553f
C988 VTAIL.n42 VSUBS 0.028553f
C989 VTAIL.n43 VSUBS 0.015343f
C990 VTAIL.n44 VSUBS 0.016246f
C991 VTAIL.n45 VSUBS 0.036265f
C992 VTAIL.n46 VSUBS 0.036265f
C993 VTAIL.n47 VSUBS 0.016246f
C994 VTAIL.n48 VSUBS 0.015343f
C995 VTAIL.n49 VSUBS 0.028553f
C996 VTAIL.n50 VSUBS 0.028553f
C997 VTAIL.n51 VSUBS 0.015343f
C998 VTAIL.n52 VSUBS 0.016246f
C999 VTAIL.n53 VSUBS 0.036265f
C1000 VTAIL.n54 VSUBS 0.036265f
C1001 VTAIL.n55 VSUBS 0.016246f
C1002 VTAIL.n56 VSUBS 0.015343f
C1003 VTAIL.n57 VSUBS 0.028553f
C1004 VTAIL.n58 VSUBS 0.073799f
C1005 VTAIL.n59 VSUBS 0.015343f
C1006 VTAIL.n60 VSUBS 0.016246f
C1007 VTAIL.n61 VSUBS 0.079142f
C1008 VTAIL.n62 VSUBS 0.053687f
C1009 VTAIL.n63 VSUBS 0.28991f
C1010 VTAIL.t6 VSUBS 0.25361f
C1011 VTAIL.t7 VSUBS 0.25361f
C1012 VTAIL.n64 VSUBS 1.84769f
C1013 VTAIL.n65 VSUBS 0.892753f
C1014 VTAIL.t1 VSUBS 0.25361f
C1015 VTAIL.t8 VSUBS 0.25361f
C1016 VTAIL.n66 VSUBS 1.84769f
C1017 VTAIL.n67 VSUBS 2.31882f
C1018 VTAIL.t12 VSUBS 0.25361f
C1019 VTAIL.t9 VSUBS 0.25361f
C1020 VTAIL.n68 VSUBS 1.8477f
C1021 VTAIL.n69 VSUBS 2.31881f
C1022 VTAIL.t15 VSUBS 0.25361f
C1023 VTAIL.t18 VSUBS 0.25361f
C1024 VTAIL.n70 VSUBS 1.8477f
C1025 VTAIL.n71 VSUBS 0.892743f
C1026 VTAIL.n72 VSUBS 0.016098f
C1027 VTAIL.n73 VSUBS 0.036265f
C1028 VTAIL.n74 VSUBS 0.016246f
C1029 VTAIL.n75 VSUBS 0.028553f
C1030 VTAIL.n76 VSUBS 0.015343f
C1031 VTAIL.n77 VSUBS 0.036265f
C1032 VTAIL.n78 VSUBS 0.016246f
C1033 VTAIL.n79 VSUBS 0.028553f
C1034 VTAIL.n80 VSUBS 0.015343f
C1035 VTAIL.n81 VSUBS 0.036265f
C1036 VTAIL.n82 VSUBS 0.016246f
C1037 VTAIL.n83 VSUBS 0.028553f
C1038 VTAIL.n84 VSUBS 0.015343f
C1039 VTAIL.n85 VSUBS 0.036265f
C1040 VTAIL.n86 VSUBS 0.016246f
C1041 VTAIL.n87 VSUBS 0.028553f
C1042 VTAIL.n88 VSUBS 0.015343f
C1043 VTAIL.n89 VSUBS 0.036265f
C1044 VTAIL.n90 VSUBS 0.016246f
C1045 VTAIL.n91 VSUBS 0.169613f
C1046 VTAIL.t13 VSUBS 0.077377f
C1047 VTAIL.n92 VSUBS 0.027199f
C1048 VTAIL.n93 VSUBS 0.02307f
C1049 VTAIL.n94 VSUBS 0.015343f
C1050 VTAIL.n95 VSUBS 1.33576f
C1051 VTAIL.n96 VSUBS 0.028553f
C1052 VTAIL.n97 VSUBS 0.015343f
C1053 VTAIL.n98 VSUBS 0.016246f
C1054 VTAIL.n99 VSUBS 0.036265f
C1055 VTAIL.n100 VSUBS 0.036265f
C1056 VTAIL.n101 VSUBS 0.016246f
C1057 VTAIL.n102 VSUBS 0.015343f
C1058 VTAIL.n103 VSUBS 0.028553f
C1059 VTAIL.n104 VSUBS 0.028553f
C1060 VTAIL.n105 VSUBS 0.015343f
C1061 VTAIL.n106 VSUBS 0.016246f
C1062 VTAIL.n107 VSUBS 0.036265f
C1063 VTAIL.n108 VSUBS 0.036265f
C1064 VTAIL.n109 VSUBS 0.016246f
C1065 VTAIL.n110 VSUBS 0.015343f
C1066 VTAIL.n111 VSUBS 0.028553f
C1067 VTAIL.n112 VSUBS 0.028553f
C1068 VTAIL.n113 VSUBS 0.015343f
C1069 VTAIL.n114 VSUBS 0.016246f
C1070 VTAIL.n115 VSUBS 0.036265f
C1071 VTAIL.n116 VSUBS 0.036265f
C1072 VTAIL.n117 VSUBS 0.016246f
C1073 VTAIL.n118 VSUBS 0.015343f
C1074 VTAIL.n119 VSUBS 0.028553f
C1075 VTAIL.n120 VSUBS 0.028553f
C1076 VTAIL.n121 VSUBS 0.015343f
C1077 VTAIL.n122 VSUBS 0.016246f
C1078 VTAIL.n123 VSUBS 0.036265f
C1079 VTAIL.n124 VSUBS 0.036265f
C1080 VTAIL.n125 VSUBS 0.016246f
C1081 VTAIL.n126 VSUBS 0.015343f
C1082 VTAIL.n127 VSUBS 0.028553f
C1083 VTAIL.n128 VSUBS 0.073799f
C1084 VTAIL.n129 VSUBS 0.015343f
C1085 VTAIL.n130 VSUBS 0.016246f
C1086 VTAIL.n131 VSUBS 0.079142f
C1087 VTAIL.n132 VSUBS 0.053687f
C1088 VTAIL.n133 VSUBS 0.28991f
C1089 VTAIL.t2 VSUBS 0.25361f
C1090 VTAIL.t19 VSUBS 0.25361f
C1091 VTAIL.n134 VSUBS 1.8477f
C1092 VTAIL.n135 VSUBS 0.862604f
C1093 VTAIL.t4 VSUBS 0.25361f
C1094 VTAIL.t5 VSUBS 0.25361f
C1095 VTAIL.n136 VSUBS 1.8477f
C1096 VTAIL.n137 VSUBS 0.892743f
C1097 VTAIL.n138 VSUBS 0.016098f
C1098 VTAIL.n139 VSUBS 0.036265f
C1099 VTAIL.n140 VSUBS 0.016246f
C1100 VTAIL.n141 VSUBS 0.028553f
C1101 VTAIL.n142 VSUBS 0.015343f
C1102 VTAIL.n143 VSUBS 0.036265f
C1103 VTAIL.n144 VSUBS 0.016246f
C1104 VTAIL.n145 VSUBS 0.028553f
C1105 VTAIL.n146 VSUBS 0.015343f
C1106 VTAIL.n147 VSUBS 0.036265f
C1107 VTAIL.n148 VSUBS 0.016246f
C1108 VTAIL.n149 VSUBS 0.028553f
C1109 VTAIL.n150 VSUBS 0.015343f
C1110 VTAIL.n151 VSUBS 0.036265f
C1111 VTAIL.n152 VSUBS 0.016246f
C1112 VTAIL.n153 VSUBS 0.028553f
C1113 VTAIL.n154 VSUBS 0.015343f
C1114 VTAIL.n155 VSUBS 0.036265f
C1115 VTAIL.n156 VSUBS 0.016246f
C1116 VTAIL.n157 VSUBS 0.169613f
C1117 VTAIL.t0 VSUBS 0.077377f
C1118 VTAIL.n158 VSUBS 0.027199f
C1119 VTAIL.n159 VSUBS 0.02307f
C1120 VTAIL.n160 VSUBS 0.015343f
C1121 VTAIL.n161 VSUBS 1.33576f
C1122 VTAIL.n162 VSUBS 0.028553f
C1123 VTAIL.n163 VSUBS 0.015343f
C1124 VTAIL.n164 VSUBS 0.016246f
C1125 VTAIL.n165 VSUBS 0.036265f
C1126 VTAIL.n166 VSUBS 0.036265f
C1127 VTAIL.n167 VSUBS 0.016246f
C1128 VTAIL.n168 VSUBS 0.015343f
C1129 VTAIL.n169 VSUBS 0.028553f
C1130 VTAIL.n170 VSUBS 0.028553f
C1131 VTAIL.n171 VSUBS 0.015343f
C1132 VTAIL.n172 VSUBS 0.016246f
C1133 VTAIL.n173 VSUBS 0.036265f
C1134 VTAIL.n174 VSUBS 0.036265f
C1135 VTAIL.n175 VSUBS 0.016246f
C1136 VTAIL.n176 VSUBS 0.015343f
C1137 VTAIL.n177 VSUBS 0.028553f
C1138 VTAIL.n178 VSUBS 0.028553f
C1139 VTAIL.n179 VSUBS 0.015343f
C1140 VTAIL.n180 VSUBS 0.016246f
C1141 VTAIL.n181 VSUBS 0.036265f
C1142 VTAIL.n182 VSUBS 0.036265f
C1143 VTAIL.n183 VSUBS 0.016246f
C1144 VTAIL.n184 VSUBS 0.015343f
C1145 VTAIL.n185 VSUBS 0.028553f
C1146 VTAIL.n186 VSUBS 0.028553f
C1147 VTAIL.n187 VSUBS 0.015343f
C1148 VTAIL.n188 VSUBS 0.016246f
C1149 VTAIL.n189 VSUBS 0.036265f
C1150 VTAIL.n190 VSUBS 0.036265f
C1151 VTAIL.n191 VSUBS 0.016246f
C1152 VTAIL.n192 VSUBS 0.015343f
C1153 VTAIL.n193 VSUBS 0.028553f
C1154 VTAIL.n194 VSUBS 0.073799f
C1155 VTAIL.n195 VSUBS 0.015343f
C1156 VTAIL.n196 VSUBS 0.016246f
C1157 VTAIL.n197 VSUBS 0.079142f
C1158 VTAIL.n198 VSUBS 0.053687f
C1159 VTAIL.n199 VSUBS 1.59938f
C1160 VTAIL.n200 VSUBS 0.016098f
C1161 VTAIL.n201 VSUBS 0.036265f
C1162 VTAIL.n202 VSUBS 0.016246f
C1163 VTAIL.n203 VSUBS 0.028553f
C1164 VTAIL.n204 VSUBS 0.015343f
C1165 VTAIL.n205 VSUBS 0.036265f
C1166 VTAIL.n206 VSUBS 0.016246f
C1167 VTAIL.n207 VSUBS 0.028553f
C1168 VTAIL.n208 VSUBS 0.015343f
C1169 VTAIL.n209 VSUBS 0.036265f
C1170 VTAIL.n210 VSUBS 0.016246f
C1171 VTAIL.n211 VSUBS 0.028553f
C1172 VTAIL.n212 VSUBS 0.015343f
C1173 VTAIL.n213 VSUBS 0.036265f
C1174 VTAIL.n214 VSUBS 0.016246f
C1175 VTAIL.n215 VSUBS 0.028553f
C1176 VTAIL.n216 VSUBS 0.015343f
C1177 VTAIL.n217 VSUBS 0.036265f
C1178 VTAIL.n218 VSUBS 0.016246f
C1179 VTAIL.n219 VSUBS 0.169613f
C1180 VTAIL.t10 VSUBS 0.077377f
C1181 VTAIL.n220 VSUBS 0.027199f
C1182 VTAIL.n221 VSUBS 0.02307f
C1183 VTAIL.n222 VSUBS 0.015343f
C1184 VTAIL.n223 VSUBS 1.33576f
C1185 VTAIL.n224 VSUBS 0.028553f
C1186 VTAIL.n225 VSUBS 0.015343f
C1187 VTAIL.n226 VSUBS 0.016246f
C1188 VTAIL.n227 VSUBS 0.036265f
C1189 VTAIL.n228 VSUBS 0.036265f
C1190 VTAIL.n229 VSUBS 0.016246f
C1191 VTAIL.n230 VSUBS 0.015343f
C1192 VTAIL.n231 VSUBS 0.028553f
C1193 VTAIL.n232 VSUBS 0.028553f
C1194 VTAIL.n233 VSUBS 0.015343f
C1195 VTAIL.n234 VSUBS 0.016246f
C1196 VTAIL.n235 VSUBS 0.036265f
C1197 VTAIL.n236 VSUBS 0.036265f
C1198 VTAIL.n237 VSUBS 0.016246f
C1199 VTAIL.n238 VSUBS 0.015343f
C1200 VTAIL.n239 VSUBS 0.028553f
C1201 VTAIL.n240 VSUBS 0.028553f
C1202 VTAIL.n241 VSUBS 0.015343f
C1203 VTAIL.n242 VSUBS 0.016246f
C1204 VTAIL.n243 VSUBS 0.036265f
C1205 VTAIL.n244 VSUBS 0.036265f
C1206 VTAIL.n245 VSUBS 0.016246f
C1207 VTAIL.n246 VSUBS 0.015343f
C1208 VTAIL.n247 VSUBS 0.028553f
C1209 VTAIL.n248 VSUBS 0.028553f
C1210 VTAIL.n249 VSUBS 0.015343f
C1211 VTAIL.n250 VSUBS 0.016246f
C1212 VTAIL.n251 VSUBS 0.036265f
C1213 VTAIL.n252 VSUBS 0.036265f
C1214 VTAIL.n253 VSUBS 0.016246f
C1215 VTAIL.n254 VSUBS 0.015343f
C1216 VTAIL.n255 VSUBS 0.028553f
C1217 VTAIL.n256 VSUBS 0.073799f
C1218 VTAIL.n257 VSUBS 0.015343f
C1219 VTAIL.n258 VSUBS 0.016246f
C1220 VTAIL.n259 VSUBS 0.079142f
C1221 VTAIL.n260 VSUBS 0.053687f
C1222 VTAIL.n261 VSUBS 1.59938f
C1223 VTAIL.t17 VSUBS 0.25361f
C1224 VTAIL.t14 VSUBS 0.25361f
C1225 VTAIL.n262 VSUBS 1.84769f
C1226 VTAIL.n263 VSUBS 0.777352f
C1227 VDD2.n0 VSUBS 0.015657f
C1228 VDD2.n1 VSUBS 0.035273f
C1229 VDD2.n2 VSUBS 0.015801f
C1230 VDD2.n3 VSUBS 0.027771f
C1231 VDD2.n4 VSUBS 0.014923f
C1232 VDD2.n5 VSUBS 0.035273f
C1233 VDD2.n6 VSUBS 0.015801f
C1234 VDD2.n7 VSUBS 0.027771f
C1235 VDD2.n8 VSUBS 0.014923f
C1236 VDD2.n9 VSUBS 0.035273f
C1237 VDD2.n10 VSUBS 0.015801f
C1238 VDD2.n11 VSUBS 0.027771f
C1239 VDD2.n12 VSUBS 0.014923f
C1240 VDD2.n13 VSUBS 0.035273f
C1241 VDD2.n14 VSUBS 0.015801f
C1242 VDD2.n15 VSUBS 0.027771f
C1243 VDD2.n16 VSUBS 0.014923f
C1244 VDD2.n17 VSUBS 0.035273f
C1245 VDD2.n18 VSUBS 0.015801f
C1246 VDD2.n19 VSUBS 0.164972f
C1247 VDD2.t8 VSUBS 0.075259f
C1248 VDD2.n20 VSUBS 0.026455f
C1249 VDD2.n21 VSUBS 0.022439f
C1250 VDD2.n22 VSUBS 0.014923f
C1251 VDD2.n23 VSUBS 1.2992f
C1252 VDD2.n24 VSUBS 0.027771f
C1253 VDD2.n25 VSUBS 0.014923f
C1254 VDD2.n26 VSUBS 0.015801f
C1255 VDD2.n27 VSUBS 0.035273f
C1256 VDD2.n28 VSUBS 0.035273f
C1257 VDD2.n29 VSUBS 0.015801f
C1258 VDD2.n30 VSUBS 0.014923f
C1259 VDD2.n31 VSUBS 0.027771f
C1260 VDD2.n32 VSUBS 0.027771f
C1261 VDD2.n33 VSUBS 0.014923f
C1262 VDD2.n34 VSUBS 0.015801f
C1263 VDD2.n35 VSUBS 0.035273f
C1264 VDD2.n36 VSUBS 0.035273f
C1265 VDD2.n37 VSUBS 0.015801f
C1266 VDD2.n38 VSUBS 0.014923f
C1267 VDD2.n39 VSUBS 0.027771f
C1268 VDD2.n40 VSUBS 0.027771f
C1269 VDD2.n41 VSUBS 0.014923f
C1270 VDD2.n42 VSUBS 0.015801f
C1271 VDD2.n43 VSUBS 0.035273f
C1272 VDD2.n44 VSUBS 0.035273f
C1273 VDD2.n45 VSUBS 0.015801f
C1274 VDD2.n46 VSUBS 0.014923f
C1275 VDD2.n47 VSUBS 0.027771f
C1276 VDD2.n48 VSUBS 0.027771f
C1277 VDD2.n49 VSUBS 0.014923f
C1278 VDD2.n50 VSUBS 0.015801f
C1279 VDD2.n51 VSUBS 0.035273f
C1280 VDD2.n52 VSUBS 0.035273f
C1281 VDD2.n53 VSUBS 0.015801f
C1282 VDD2.n54 VSUBS 0.014923f
C1283 VDD2.n55 VSUBS 0.027771f
C1284 VDD2.n56 VSUBS 0.07178f
C1285 VDD2.n57 VSUBS 0.014923f
C1286 VDD2.n58 VSUBS 0.015801f
C1287 VDD2.n59 VSUBS 0.076976f
C1288 VDD2.n60 VSUBS 0.077402f
C1289 VDD2.t1 VSUBS 0.24667f
C1290 VDD2.t0 VSUBS 0.24667f
C1291 VDD2.n61 VSUBS 1.92844f
C1292 VDD2.n62 VSUBS 0.856972f
C1293 VDD2.t2 VSUBS 0.24667f
C1294 VDD2.t7 VSUBS 0.24667f
C1295 VDD2.n63 VSUBS 1.93917f
C1296 VDD2.n64 VSUBS 2.80483f
C1297 VDD2.n65 VSUBS 0.015657f
C1298 VDD2.n66 VSUBS 0.035273f
C1299 VDD2.n67 VSUBS 0.015801f
C1300 VDD2.n68 VSUBS 0.027771f
C1301 VDD2.n69 VSUBS 0.014923f
C1302 VDD2.n70 VSUBS 0.035273f
C1303 VDD2.n71 VSUBS 0.015801f
C1304 VDD2.n72 VSUBS 0.027771f
C1305 VDD2.n73 VSUBS 0.014923f
C1306 VDD2.n74 VSUBS 0.035273f
C1307 VDD2.n75 VSUBS 0.015801f
C1308 VDD2.n76 VSUBS 0.027771f
C1309 VDD2.n77 VSUBS 0.014923f
C1310 VDD2.n78 VSUBS 0.035273f
C1311 VDD2.n79 VSUBS 0.015801f
C1312 VDD2.n80 VSUBS 0.027771f
C1313 VDD2.n81 VSUBS 0.014923f
C1314 VDD2.n82 VSUBS 0.035273f
C1315 VDD2.n83 VSUBS 0.015801f
C1316 VDD2.n84 VSUBS 0.164972f
C1317 VDD2.t9 VSUBS 0.07526f
C1318 VDD2.n85 VSUBS 0.026455f
C1319 VDD2.n86 VSUBS 0.022439f
C1320 VDD2.n87 VSUBS 0.014923f
C1321 VDD2.n88 VSUBS 1.2992f
C1322 VDD2.n89 VSUBS 0.027771f
C1323 VDD2.n90 VSUBS 0.014923f
C1324 VDD2.n91 VSUBS 0.015801f
C1325 VDD2.n92 VSUBS 0.035273f
C1326 VDD2.n93 VSUBS 0.035273f
C1327 VDD2.n94 VSUBS 0.015801f
C1328 VDD2.n95 VSUBS 0.014923f
C1329 VDD2.n96 VSUBS 0.027771f
C1330 VDD2.n97 VSUBS 0.027771f
C1331 VDD2.n98 VSUBS 0.014923f
C1332 VDD2.n99 VSUBS 0.015801f
C1333 VDD2.n100 VSUBS 0.035273f
C1334 VDD2.n101 VSUBS 0.035273f
C1335 VDD2.n102 VSUBS 0.015801f
C1336 VDD2.n103 VSUBS 0.014923f
C1337 VDD2.n104 VSUBS 0.027771f
C1338 VDD2.n105 VSUBS 0.027771f
C1339 VDD2.n106 VSUBS 0.014923f
C1340 VDD2.n107 VSUBS 0.015801f
C1341 VDD2.n108 VSUBS 0.035273f
C1342 VDD2.n109 VSUBS 0.035273f
C1343 VDD2.n110 VSUBS 0.015801f
C1344 VDD2.n111 VSUBS 0.014923f
C1345 VDD2.n112 VSUBS 0.027771f
C1346 VDD2.n113 VSUBS 0.027771f
C1347 VDD2.n114 VSUBS 0.014923f
C1348 VDD2.n115 VSUBS 0.015801f
C1349 VDD2.n116 VSUBS 0.035273f
C1350 VDD2.n117 VSUBS 0.035273f
C1351 VDD2.n118 VSUBS 0.015801f
C1352 VDD2.n119 VSUBS 0.014923f
C1353 VDD2.n120 VSUBS 0.027771f
C1354 VDD2.n121 VSUBS 0.07178f
C1355 VDD2.n122 VSUBS 0.014923f
C1356 VDD2.n123 VSUBS 0.015801f
C1357 VDD2.n124 VSUBS 0.076976f
C1358 VDD2.n125 VSUBS 0.071365f
C1359 VDD2.n126 VSUBS 2.68152f
C1360 VDD2.t4 VSUBS 0.24667f
C1361 VDD2.t3 VSUBS 0.24667f
C1362 VDD2.n127 VSUBS 1.92845f
C1363 VDD2.n128 VSUBS 0.672926f
C1364 VDD2.t5 VSUBS 0.24667f
C1365 VDD2.t6 VSUBS 0.24667f
C1366 VDD2.n129 VSUBS 1.93913f
C1367 VN.n0 VSUBS 0.037832f
C1368 VN.t8 VSUBS 1.75766f
C1369 VN.n1 VSUBS 0.058122f
C1370 VN.n2 VSUBS 0.037832f
C1371 VN.t4 VSUBS 1.75766f
C1372 VN.n3 VSUBS 0.071548f
C1373 VN.n4 VSUBS 0.037832f
C1374 VN.t1 VSUBS 1.75766f
C1375 VN.n5 VSUBS 0.066294f
C1376 VN.t7 VSUBS 1.88244f
C1377 VN.t2 VSUBS 1.75766f
C1378 VN.n6 VSUBS 0.71712f
C1379 VN.n7 VSUBS 0.72602f
C1380 VN.n8 VSUBS 0.239868f
C1381 VN.n9 VSUBS 0.037832f
C1382 VN.n10 VSUBS 0.033461f
C1383 VN.n11 VSUBS 0.071548f
C1384 VN.n12 VSUBS 0.674656f
C1385 VN.n13 VSUBS 0.037832f
C1386 VN.n14 VSUBS 0.037832f
C1387 VN.n15 VSUBS 0.037832f
C1388 VN.n16 VSUBS 0.033461f
C1389 VN.n17 VSUBS 0.066294f
C1390 VN.n18 VSUBS 0.638781f
C1391 VN.n19 VSUBS 0.046371f
C1392 VN.n20 VSUBS 0.037832f
C1393 VN.n21 VSUBS 0.037832f
C1394 VN.n22 VSUBS 0.037832f
C1395 VN.n23 VSUBS 0.052814f
C1396 VN.n24 VSUBS 0.04987f
C1397 VN.n25 VSUBS 0.717876f
C1398 VN.n26 VSUBS 0.03648f
C1399 VN.n27 VSUBS 0.037832f
C1400 VN.t6 VSUBS 1.75766f
C1401 VN.n28 VSUBS 0.058122f
C1402 VN.n29 VSUBS 0.037832f
C1403 VN.t9 VSUBS 1.75766f
C1404 VN.n30 VSUBS 0.071548f
C1405 VN.n31 VSUBS 0.037832f
C1406 VN.t3 VSUBS 1.75766f
C1407 VN.n32 VSUBS 0.066294f
C1408 VN.t5 VSUBS 1.88244f
C1409 VN.t0 VSUBS 1.75766f
C1410 VN.n33 VSUBS 0.71712f
C1411 VN.n34 VSUBS 0.72602f
C1412 VN.n35 VSUBS 0.239868f
C1413 VN.n36 VSUBS 0.037832f
C1414 VN.n37 VSUBS 0.033461f
C1415 VN.n38 VSUBS 0.071548f
C1416 VN.n39 VSUBS 0.674656f
C1417 VN.n40 VSUBS 0.037832f
C1418 VN.n41 VSUBS 0.037832f
C1419 VN.n42 VSUBS 0.037832f
C1420 VN.n43 VSUBS 0.033461f
C1421 VN.n44 VSUBS 0.066294f
C1422 VN.n45 VSUBS 0.638781f
C1423 VN.n46 VSUBS 0.046371f
C1424 VN.n47 VSUBS 0.037832f
C1425 VN.n48 VSUBS 0.037832f
C1426 VN.n49 VSUBS 0.037832f
C1427 VN.n50 VSUBS 0.052814f
C1428 VN.n51 VSUBS 0.04987f
C1429 VN.n52 VSUBS 0.717876f
C1430 VN.n53 VSUBS 1.87804f
.ends

