* NGSPICE file created from diff_pair_sample_1655.ext - technology: sky130A

.subckt diff_pair_sample_1655 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t7 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X1 VDD1.t1 VP.t1 VTAIL.t17 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X2 VTAIL.t1 VN.t0 VDD2.t9 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X3 VTAIL.t5 VN.t1 VDD2.t8 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X4 B.t11 B.t9 B.t10 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=0 ps=0 w=12.58 l=3.04
X5 VDD1.t0 VP.t2 VTAIL.t16 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=4.9062 ps=25.94 w=12.58 l=3.04
X6 VDD1.t6 VP.t3 VTAIL.t15 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X7 VTAIL.t2 VN.t2 VDD2.t7 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X8 VTAIL.t14 VP.t4 VDD1.t5 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X9 B.t8 B.t6 B.t7 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=0 ps=0 w=12.58 l=3.04
X10 B.t5 B.t3 B.t4 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=0 ps=0 w=12.58 l=3.04
X11 VDD2.t6 VN.t3 VTAIL.t7 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=4.9062 ps=25.94 w=12.58 l=3.04
X12 VTAIL.t13 VP.t5 VDD1.t9 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X13 VDD2.t5 VN.t4 VTAIL.t19 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=2.0757 ps=12.91 w=12.58 l=3.04
X14 VDD2.t4 VN.t5 VTAIL.t4 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=2.0757 ps=12.91 w=12.58 l=3.04
X15 VDD1.t8 VP.t6 VTAIL.t12 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=4.9062 ps=25.94 w=12.58 l=3.04
X16 VDD2.t3 VN.t6 VTAIL.t0 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X17 B.t2 B.t0 B.t1 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=0 ps=0 w=12.58 l=3.04
X18 VTAIL.t3 VN.t7 VDD2.t2 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X19 VDD1.t4 VP.t7 VTAIL.t11 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=2.0757 ps=12.91 w=12.58 l=3.04
X20 VDD1.t3 VP.t8 VTAIL.t10 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=4.9062 pd=25.94 as=2.0757 ps=12.91 w=12.58 l=3.04
X21 VTAIL.t9 VP.t9 VDD1.t2 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X22 VDD2.t1 VN.t8 VTAIL.t6 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=2.0757 ps=12.91 w=12.58 l=3.04
X23 VDD2.t0 VN.t9 VTAIL.t8 w_n5014_n3484# sky130_fd_pr__pfet_01v8 ad=2.0757 pd=12.91 as=4.9062 ps=25.94 w=12.58 l=3.04
R0 VP.n27 VP.n24 161.3
R1 VP.n29 VP.n28 161.3
R2 VP.n30 VP.n23 161.3
R3 VP.n32 VP.n31 161.3
R4 VP.n33 VP.n22 161.3
R5 VP.n35 VP.n34 161.3
R6 VP.n36 VP.n21 161.3
R7 VP.n39 VP.n38 161.3
R8 VP.n40 VP.n20 161.3
R9 VP.n42 VP.n41 161.3
R10 VP.n43 VP.n19 161.3
R11 VP.n45 VP.n44 161.3
R12 VP.n46 VP.n18 161.3
R13 VP.n48 VP.n47 161.3
R14 VP.n50 VP.n17 161.3
R15 VP.n52 VP.n51 161.3
R16 VP.n53 VP.n16 161.3
R17 VP.n55 VP.n54 161.3
R18 VP.n56 VP.n15 161.3
R19 VP.n58 VP.n57 161.3
R20 VP.n103 VP.n102 161.3
R21 VP.n101 VP.n1 161.3
R22 VP.n100 VP.n99 161.3
R23 VP.n98 VP.n2 161.3
R24 VP.n97 VP.n96 161.3
R25 VP.n95 VP.n3 161.3
R26 VP.n93 VP.n92 161.3
R27 VP.n91 VP.n4 161.3
R28 VP.n90 VP.n89 161.3
R29 VP.n88 VP.n5 161.3
R30 VP.n87 VP.n86 161.3
R31 VP.n85 VP.n6 161.3
R32 VP.n84 VP.n83 161.3
R33 VP.n81 VP.n7 161.3
R34 VP.n80 VP.n79 161.3
R35 VP.n78 VP.n8 161.3
R36 VP.n77 VP.n76 161.3
R37 VP.n75 VP.n9 161.3
R38 VP.n74 VP.n73 161.3
R39 VP.n72 VP.n10 161.3
R40 VP.n71 VP.n70 161.3
R41 VP.n68 VP.n11 161.3
R42 VP.n67 VP.n66 161.3
R43 VP.n65 VP.n12 161.3
R44 VP.n64 VP.n63 161.3
R45 VP.n62 VP.n13 161.3
R46 VP.n26 VP.t8 131.565
R47 VP.n61 VP.t7 99.7301
R48 VP.n69 VP.t9 99.7301
R49 VP.n82 VP.t3 99.7301
R50 VP.n94 VP.t0 99.7301
R51 VP.n0 VP.t2 99.7301
R52 VP.n14 VP.t6 99.7301
R53 VP.n49 VP.t5 99.7301
R54 VP.n37 VP.t1 99.7301
R55 VP.n25 VP.t4 99.7301
R56 VP.n26 VP.n25 68.2679
R57 VP.n61 VP.n60 66.1456
R58 VP.n104 VP.n0 66.1456
R59 VP.n59 VP.n14 66.1456
R60 VP.n67 VP.n12 56.5617
R61 VP.n100 VP.n2 56.5617
R62 VP.n55 VP.n16 56.5617
R63 VP.n60 VP.n59 56.1397
R64 VP.n76 VP.n8 46.874
R65 VP.n88 VP.n87 46.874
R66 VP.n43 VP.n42 46.874
R67 VP.n31 VP.n22 46.874
R68 VP.n76 VP.n75 34.28
R69 VP.n89 VP.n88 34.28
R70 VP.n44 VP.n43 34.28
R71 VP.n31 VP.n30 34.28
R72 VP.n63 VP.n62 24.5923
R73 VP.n63 VP.n12 24.5923
R74 VP.n68 VP.n67 24.5923
R75 VP.n70 VP.n68 24.5923
R76 VP.n74 VP.n10 24.5923
R77 VP.n75 VP.n74 24.5923
R78 VP.n80 VP.n8 24.5923
R79 VP.n81 VP.n80 24.5923
R80 VP.n83 VP.n6 24.5923
R81 VP.n87 VP.n6 24.5923
R82 VP.n89 VP.n4 24.5923
R83 VP.n93 VP.n4 24.5923
R84 VP.n96 VP.n95 24.5923
R85 VP.n96 VP.n2 24.5923
R86 VP.n101 VP.n100 24.5923
R87 VP.n102 VP.n101 24.5923
R88 VP.n56 VP.n55 24.5923
R89 VP.n57 VP.n56 24.5923
R90 VP.n44 VP.n18 24.5923
R91 VP.n48 VP.n18 24.5923
R92 VP.n51 VP.n50 24.5923
R93 VP.n51 VP.n16 24.5923
R94 VP.n35 VP.n22 24.5923
R95 VP.n36 VP.n35 24.5923
R96 VP.n38 VP.n20 24.5923
R97 VP.n42 VP.n20 24.5923
R98 VP.n29 VP.n24 24.5923
R99 VP.n30 VP.n29 24.5923
R100 VP.n62 VP.n61 24.1005
R101 VP.n102 VP.n0 24.1005
R102 VP.n57 VP.n14 24.1005
R103 VP.n70 VP.n69 18.6903
R104 VP.n95 VP.n94 18.6903
R105 VP.n50 VP.n49 18.6903
R106 VP.n82 VP.n81 12.2964
R107 VP.n83 VP.n82 12.2964
R108 VP.n37 VP.n36 12.2964
R109 VP.n38 VP.n37 12.2964
R110 VP.n69 VP.n10 5.90254
R111 VP.n94 VP.n93 5.90254
R112 VP.n49 VP.n48 5.90254
R113 VP.n25 VP.n24 5.90254
R114 VP.n27 VP.n26 5.25066
R115 VP.n59 VP.n58 0.354861
R116 VP.n60 VP.n13 0.354861
R117 VP.n104 VP.n103 0.354861
R118 VP VP.n104 0.267071
R119 VP.n28 VP.n27 0.189894
R120 VP.n28 VP.n23 0.189894
R121 VP.n32 VP.n23 0.189894
R122 VP.n33 VP.n32 0.189894
R123 VP.n34 VP.n33 0.189894
R124 VP.n34 VP.n21 0.189894
R125 VP.n39 VP.n21 0.189894
R126 VP.n40 VP.n39 0.189894
R127 VP.n41 VP.n40 0.189894
R128 VP.n41 VP.n19 0.189894
R129 VP.n45 VP.n19 0.189894
R130 VP.n46 VP.n45 0.189894
R131 VP.n47 VP.n46 0.189894
R132 VP.n47 VP.n17 0.189894
R133 VP.n52 VP.n17 0.189894
R134 VP.n53 VP.n52 0.189894
R135 VP.n54 VP.n53 0.189894
R136 VP.n54 VP.n15 0.189894
R137 VP.n58 VP.n15 0.189894
R138 VP.n64 VP.n13 0.189894
R139 VP.n65 VP.n64 0.189894
R140 VP.n66 VP.n65 0.189894
R141 VP.n66 VP.n11 0.189894
R142 VP.n71 VP.n11 0.189894
R143 VP.n72 VP.n71 0.189894
R144 VP.n73 VP.n72 0.189894
R145 VP.n73 VP.n9 0.189894
R146 VP.n77 VP.n9 0.189894
R147 VP.n78 VP.n77 0.189894
R148 VP.n79 VP.n78 0.189894
R149 VP.n79 VP.n7 0.189894
R150 VP.n84 VP.n7 0.189894
R151 VP.n85 VP.n84 0.189894
R152 VP.n86 VP.n85 0.189894
R153 VP.n86 VP.n5 0.189894
R154 VP.n90 VP.n5 0.189894
R155 VP.n91 VP.n90 0.189894
R156 VP.n92 VP.n91 0.189894
R157 VP.n92 VP.n3 0.189894
R158 VP.n97 VP.n3 0.189894
R159 VP.n98 VP.n97 0.189894
R160 VP.n99 VP.n98 0.189894
R161 VP.n99 VP.n1 0.189894
R162 VP.n103 VP.n1 0.189894
R163 VDD1.n68 VDD1.n67 756.745
R164 VDD1.n139 VDD1.n138 756.745
R165 VDD1.n67 VDD1.n66 585
R166 VDD1.n2 VDD1.n1 585
R167 VDD1.n61 VDD1.n60 585
R168 VDD1.n59 VDD1.n58 585
R169 VDD1.n6 VDD1.n5 585
R170 VDD1.n53 VDD1.n52 585
R171 VDD1.n51 VDD1.n50 585
R172 VDD1.n10 VDD1.n9 585
R173 VDD1.n45 VDD1.n44 585
R174 VDD1.n43 VDD1.n42 585
R175 VDD1.n14 VDD1.n13 585
R176 VDD1.n37 VDD1.n36 585
R177 VDD1.n35 VDD1.n34 585
R178 VDD1.n18 VDD1.n17 585
R179 VDD1.n29 VDD1.n28 585
R180 VDD1.n27 VDD1.n26 585
R181 VDD1.n22 VDD1.n21 585
R182 VDD1.n93 VDD1.n92 585
R183 VDD1.n98 VDD1.n97 585
R184 VDD1.n100 VDD1.n99 585
R185 VDD1.n89 VDD1.n88 585
R186 VDD1.n106 VDD1.n105 585
R187 VDD1.n108 VDD1.n107 585
R188 VDD1.n85 VDD1.n84 585
R189 VDD1.n114 VDD1.n113 585
R190 VDD1.n116 VDD1.n115 585
R191 VDD1.n81 VDD1.n80 585
R192 VDD1.n122 VDD1.n121 585
R193 VDD1.n124 VDD1.n123 585
R194 VDD1.n77 VDD1.n76 585
R195 VDD1.n130 VDD1.n129 585
R196 VDD1.n132 VDD1.n131 585
R197 VDD1.n73 VDD1.n72 585
R198 VDD1.n138 VDD1.n137 585
R199 VDD1.n23 VDD1.t3 327.466
R200 VDD1.n94 VDD1.t4 327.466
R201 VDD1.n67 VDD1.n1 171.744
R202 VDD1.n60 VDD1.n1 171.744
R203 VDD1.n60 VDD1.n59 171.744
R204 VDD1.n59 VDD1.n5 171.744
R205 VDD1.n52 VDD1.n5 171.744
R206 VDD1.n52 VDD1.n51 171.744
R207 VDD1.n51 VDD1.n9 171.744
R208 VDD1.n44 VDD1.n9 171.744
R209 VDD1.n44 VDD1.n43 171.744
R210 VDD1.n43 VDD1.n13 171.744
R211 VDD1.n36 VDD1.n13 171.744
R212 VDD1.n36 VDD1.n35 171.744
R213 VDD1.n35 VDD1.n17 171.744
R214 VDD1.n28 VDD1.n17 171.744
R215 VDD1.n28 VDD1.n27 171.744
R216 VDD1.n27 VDD1.n21 171.744
R217 VDD1.n98 VDD1.n92 171.744
R218 VDD1.n99 VDD1.n98 171.744
R219 VDD1.n99 VDD1.n88 171.744
R220 VDD1.n106 VDD1.n88 171.744
R221 VDD1.n107 VDD1.n106 171.744
R222 VDD1.n107 VDD1.n84 171.744
R223 VDD1.n114 VDD1.n84 171.744
R224 VDD1.n115 VDD1.n114 171.744
R225 VDD1.n115 VDD1.n80 171.744
R226 VDD1.n122 VDD1.n80 171.744
R227 VDD1.n123 VDD1.n122 171.744
R228 VDD1.n123 VDD1.n76 171.744
R229 VDD1.n130 VDD1.n76 171.744
R230 VDD1.n131 VDD1.n130 171.744
R231 VDD1.n131 VDD1.n72 171.744
R232 VDD1.n138 VDD1.n72 171.744
R233 VDD1.t3 VDD1.n21 85.8723
R234 VDD1.t4 VDD1.n92 85.8723
R235 VDD1.n143 VDD1.n142 76.7177
R236 VDD1.n70 VDD1.n69 74.5952
R237 VDD1.n141 VDD1.n140 74.5942
R238 VDD1.n145 VDD1.n144 74.5941
R239 VDD1.n70 VDD1.n68 53.3208
R240 VDD1.n141 VDD1.n139 53.3208
R241 VDD1.n145 VDD1.n143 50.3953
R242 VDD1.n23 VDD1.n22 16.3895
R243 VDD1.n94 VDD1.n93 16.3895
R244 VDD1.n66 VDD1.n0 12.8005
R245 VDD1.n26 VDD1.n25 12.8005
R246 VDD1.n97 VDD1.n96 12.8005
R247 VDD1.n137 VDD1.n71 12.8005
R248 VDD1.n65 VDD1.n2 12.0247
R249 VDD1.n29 VDD1.n20 12.0247
R250 VDD1.n100 VDD1.n91 12.0247
R251 VDD1.n136 VDD1.n73 12.0247
R252 VDD1.n62 VDD1.n61 11.249
R253 VDD1.n30 VDD1.n18 11.249
R254 VDD1.n101 VDD1.n89 11.249
R255 VDD1.n133 VDD1.n132 11.249
R256 VDD1.n58 VDD1.n4 10.4732
R257 VDD1.n34 VDD1.n33 10.4732
R258 VDD1.n105 VDD1.n104 10.4732
R259 VDD1.n129 VDD1.n75 10.4732
R260 VDD1.n57 VDD1.n6 9.69747
R261 VDD1.n37 VDD1.n16 9.69747
R262 VDD1.n108 VDD1.n87 9.69747
R263 VDD1.n128 VDD1.n77 9.69747
R264 VDD1.n64 VDD1.n0 9.45567
R265 VDD1.n135 VDD1.n71 9.45567
R266 VDD1.n49 VDD1.n48 9.3005
R267 VDD1.n8 VDD1.n7 9.3005
R268 VDD1.n55 VDD1.n54 9.3005
R269 VDD1.n57 VDD1.n56 9.3005
R270 VDD1.n4 VDD1.n3 9.3005
R271 VDD1.n63 VDD1.n62 9.3005
R272 VDD1.n65 VDD1.n64 9.3005
R273 VDD1.n47 VDD1.n46 9.3005
R274 VDD1.n12 VDD1.n11 9.3005
R275 VDD1.n41 VDD1.n40 9.3005
R276 VDD1.n39 VDD1.n38 9.3005
R277 VDD1.n16 VDD1.n15 9.3005
R278 VDD1.n33 VDD1.n32 9.3005
R279 VDD1.n31 VDD1.n30 9.3005
R280 VDD1.n20 VDD1.n19 9.3005
R281 VDD1.n25 VDD1.n24 9.3005
R282 VDD1.n118 VDD1.n117 9.3005
R283 VDD1.n120 VDD1.n119 9.3005
R284 VDD1.n79 VDD1.n78 9.3005
R285 VDD1.n126 VDD1.n125 9.3005
R286 VDD1.n128 VDD1.n127 9.3005
R287 VDD1.n75 VDD1.n74 9.3005
R288 VDD1.n134 VDD1.n133 9.3005
R289 VDD1.n136 VDD1.n135 9.3005
R290 VDD1.n112 VDD1.n111 9.3005
R291 VDD1.n110 VDD1.n109 9.3005
R292 VDD1.n87 VDD1.n86 9.3005
R293 VDD1.n104 VDD1.n103 9.3005
R294 VDD1.n102 VDD1.n101 9.3005
R295 VDD1.n91 VDD1.n90 9.3005
R296 VDD1.n96 VDD1.n95 9.3005
R297 VDD1.n83 VDD1.n82 9.3005
R298 VDD1.n54 VDD1.n53 8.92171
R299 VDD1.n38 VDD1.n14 8.92171
R300 VDD1.n109 VDD1.n85 8.92171
R301 VDD1.n125 VDD1.n124 8.92171
R302 VDD1.n50 VDD1.n8 8.14595
R303 VDD1.n42 VDD1.n41 8.14595
R304 VDD1.n113 VDD1.n112 8.14595
R305 VDD1.n121 VDD1.n79 8.14595
R306 VDD1.n49 VDD1.n10 7.3702
R307 VDD1.n45 VDD1.n12 7.3702
R308 VDD1.n116 VDD1.n83 7.3702
R309 VDD1.n120 VDD1.n81 7.3702
R310 VDD1.n46 VDD1.n10 6.59444
R311 VDD1.n46 VDD1.n45 6.59444
R312 VDD1.n117 VDD1.n116 6.59444
R313 VDD1.n117 VDD1.n81 6.59444
R314 VDD1.n50 VDD1.n49 5.81868
R315 VDD1.n42 VDD1.n12 5.81868
R316 VDD1.n113 VDD1.n83 5.81868
R317 VDD1.n121 VDD1.n120 5.81868
R318 VDD1.n53 VDD1.n8 5.04292
R319 VDD1.n41 VDD1.n14 5.04292
R320 VDD1.n112 VDD1.n85 5.04292
R321 VDD1.n124 VDD1.n79 5.04292
R322 VDD1.n54 VDD1.n6 4.26717
R323 VDD1.n38 VDD1.n37 4.26717
R324 VDD1.n109 VDD1.n108 4.26717
R325 VDD1.n125 VDD1.n77 4.26717
R326 VDD1.n24 VDD1.n23 3.70982
R327 VDD1.n95 VDD1.n94 3.70982
R328 VDD1.n58 VDD1.n57 3.49141
R329 VDD1.n34 VDD1.n16 3.49141
R330 VDD1.n105 VDD1.n87 3.49141
R331 VDD1.n129 VDD1.n128 3.49141
R332 VDD1.n61 VDD1.n4 2.71565
R333 VDD1.n33 VDD1.n18 2.71565
R334 VDD1.n104 VDD1.n89 2.71565
R335 VDD1.n132 VDD1.n75 2.71565
R336 VDD1.n144 VDD1.t9 2.58436
R337 VDD1.n144 VDD1.t8 2.58436
R338 VDD1.n69 VDD1.t5 2.58436
R339 VDD1.n69 VDD1.t1 2.58436
R340 VDD1.n142 VDD1.t7 2.58436
R341 VDD1.n142 VDD1.t0 2.58436
R342 VDD1.n140 VDD1.t2 2.58436
R343 VDD1.n140 VDD1.t6 2.58436
R344 VDD1 VDD1.n145 2.12119
R345 VDD1.n62 VDD1.n2 1.93989
R346 VDD1.n30 VDD1.n29 1.93989
R347 VDD1.n101 VDD1.n100 1.93989
R348 VDD1.n133 VDD1.n73 1.93989
R349 VDD1.n66 VDD1.n65 1.16414
R350 VDD1.n26 VDD1.n20 1.16414
R351 VDD1.n97 VDD1.n91 1.16414
R352 VDD1.n137 VDD1.n136 1.16414
R353 VDD1 VDD1.n70 0.784983
R354 VDD1.n143 VDD1.n141 0.671447
R355 VDD1.n68 VDD1.n0 0.388379
R356 VDD1.n25 VDD1.n22 0.388379
R357 VDD1.n96 VDD1.n93 0.388379
R358 VDD1.n139 VDD1.n71 0.388379
R359 VDD1.n64 VDD1.n63 0.155672
R360 VDD1.n63 VDD1.n3 0.155672
R361 VDD1.n56 VDD1.n3 0.155672
R362 VDD1.n56 VDD1.n55 0.155672
R363 VDD1.n55 VDD1.n7 0.155672
R364 VDD1.n48 VDD1.n7 0.155672
R365 VDD1.n48 VDD1.n47 0.155672
R366 VDD1.n47 VDD1.n11 0.155672
R367 VDD1.n40 VDD1.n11 0.155672
R368 VDD1.n40 VDD1.n39 0.155672
R369 VDD1.n39 VDD1.n15 0.155672
R370 VDD1.n32 VDD1.n15 0.155672
R371 VDD1.n32 VDD1.n31 0.155672
R372 VDD1.n31 VDD1.n19 0.155672
R373 VDD1.n24 VDD1.n19 0.155672
R374 VDD1.n95 VDD1.n90 0.155672
R375 VDD1.n102 VDD1.n90 0.155672
R376 VDD1.n103 VDD1.n102 0.155672
R377 VDD1.n103 VDD1.n86 0.155672
R378 VDD1.n110 VDD1.n86 0.155672
R379 VDD1.n111 VDD1.n110 0.155672
R380 VDD1.n111 VDD1.n82 0.155672
R381 VDD1.n118 VDD1.n82 0.155672
R382 VDD1.n119 VDD1.n118 0.155672
R383 VDD1.n119 VDD1.n78 0.155672
R384 VDD1.n126 VDD1.n78 0.155672
R385 VDD1.n127 VDD1.n126 0.155672
R386 VDD1.n127 VDD1.n74 0.155672
R387 VDD1.n134 VDD1.n74 0.155672
R388 VDD1.n135 VDD1.n134 0.155672
R389 VTAIL.n292 VTAIL.n291 756.745
R390 VTAIL.n70 VTAIL.n69 756.745
R391 VTAIL.n222 VTAIL.n221 756.745
R392 VTAIL.n148 VTAIL.n147 756.745
R393 VTAIL.n246 VTAIL.n245 585
R394 VTAIL.n251 VTAIL.n250 585
R395 VTAIL.n253 VTAIL.n252 585
R396 VTAIL.n242 VTAIL.n241 585
R397 VTAIL.n259 VTAIL.n258 585
R398 VTAIL.n261 VTAIL.n260 585
R399 VTAIL.n238 VTAIL.n237 585
R400 VTAIL.n267 VTAIL.n266 585
R401 VTAIL.n269 VTAIL.n268 585
R402 VTAIL.n234 VTAIL.n233 585
R403 VTAIL.n275 VTAIL.n274 585
R404 VTAIL.n277 VTAIL.n276 585
R405 VTAIL.n230 VTAIL.n229 585
R406 VTAIL.n283 VTAIL.n282 585
R407 VTAIL.n285 VTAIL.n284 585
R408 VTAIL.n226 VTAIL.n225 585
R409 VTAIL.n291 VTAIL.n290 585
R410 VTAIL.n24 VTAIL.n23 585
R411 VTAIL.n29 VTAIL.n28 585
R412 VTAIL.n31 VTAIL.n30 585
R413 VTAIL.n20 VTAIL.n19 585
R414 VTAIL.n37 VTAIL.n36 585
R415 VTAIL.n39 VTAIL.n38 585
R416 VTAIL.n16 VTAIL.n15 585
R417 VTAIL.n45 VTAIL.n44 585
R418 VTAIL.n47 VTAIL.n46 585
R419 VTAIL.n12 VTAIL.n11 585
R420 VTAIL.n53 VTAIL.n52 585
R421 VTAIL.n55 VTAIL.n54 585
R422 VTAIL.n8 VTAIL.n7 585
R423 VTAIL.n61 VTAIL.n60 585
R424 VTAIL.n63 VTAIL.n62 585
R425 VTAIL.n4 VTAIL.n3 585
R426 VTAIL.n69 VTAIL.n68 585
R427 VTAIL.n221 VTAIL.n220 585
R428 VTAIL.n156 VTAIL.n155 585
R429 VTAIL.n215 VTAIL.n214 585
R430 VTAIL.n213 VTAIL.n212 585
R431 VTAIL.n160 VTAIL.n159 585
R432 VTAIL.n207 VTAIL.n206 585
R433 VTAIL.n205 VTAIL.n204 585
R434 VTAIL.n164 VTAIL.n163 585
R435 VTAIL.n199 VTAIL.n198 585
R436 VTAIL.n197 VTAIL.n196 585
R437 VTAIL.n168 VTAIL.n167 585
R438 VTAIL.n191 VTAIL.n190 585
R439 VTAIL.n189 VTAIL.n188 585
R440 VTAIL.n172 VTAIL.n171 585
R441 VTAIL.n183 VTAIL.n182 585
R442 VTAIL.n181 VTAIL.n180 585
R443 VTAIL.n176 VTAIL.n175 585
R444 VTAIL.n147 VTAIL.n146 585
R445 VTAIL.n82 VTAIL.n81 585
R446 VTAIL.n141 VTAIL.n140 585
R447 VTAIL.n139 VTAIL.n138 585
R448 VTAIL.n86 VTAIL.n85 585
R449 VTAIL.n133 VTAIL.n132 585
R450 VTAIL.n131 VTAIL.n130 585
R451 VTAIL.n90 VTAIL.n89 585
R452 VTAIL.n125 VTAIL.n124 585
R453 VTAIL.n123 VTAIL.n122 585
R454 VTAIL.n94 VTAIL.n93 585
R455 VTAIL.n117 VTAIL.n116 585
R456 VTAIL.n115 VTAIL.n114 585
R457 VTAIL.n98 VTAIL.n97 585
R458 VTAIL.n109 VTAIL.n108 585
R459 VTAIL.n107 VTAIL.n106 585
R460 VTAIL.n102 VTAIL.n101 585
R461 VTAIL.n247 VTAIL.t8 327.466
R462 VTAIL.n25 VTAIL.t16 327.466
R463 VTAIL.n177 VTAIL.t12 327.466
R464 VTAIL.n103 VTAIL.t7 327.466
R465 VTAIL.n251 VTAIL.n245 171.744
R466 VTAIL.n252 VTAIL.n251 171.744
R467 VTAIL.n252 VTAIL.n241 171.744
R468 VTAIL.n259 VTAIL.n241 171.744
R469 VTAIL.n260 VTAIL.n259 171.744
R470 VTAIL.n260 VTAIL.n237 171.744
R471 VTAIL.n267 VTAIL.n237 171.744
R472 VTAIL.n268 VTAIL.n267 171.744
R473 VTAIL.n268 VTAIL.n233 171.744
R474 VTAIL.n275 VTAIL.n233 171.744
R475 VTAIL.n276 VTAIL.n275 171.744
R476 VTAIL.n276 VTAIL.n229 171.744
R477 VTAIL.n283 VTAIL.n229 171.744
R478 VTAIL.n284 VTAIL.n283 171.744
R479 VTAIL.n284 VTAIL.n225 171.744
R480 VTAIL.n291 VTAIL.n225 171.744
R481 VTAIL.n29 VTAIL.n23 171.744
R482 VTAIL.n30 VTAIL.n29 171.744
R483 VTAIL.n30 VTAIL.n19 171.744
R484 VTAIL.n37 VTAIL.n19 171.744
R485 VTAIL.n38 VTAIL.n37 171.744
R486 VTAIL.n38 VTAIL.n15 171.744
R487 VTAIL.n45 VTAIL.n15 171.744
R488 VTAIL.n46 VTAIL.n45 171.744
R489 VTAIL.n46 VTAIL.n11 171.744
R490 VTAIL.n53 VTAIL.n11 171.744
R491 VTAIL.n54 VTAIL.n53 171.744
R492 VTAIL.n54 VTAIL.n7 171.744
R493 VTAIL.n61 VTAIL.n7 171.744
R494 VTAIL.n62 VTAIL.n61 171.744
R495 VTAIL.n62 VTAIL.n3 171.744
R496 VTAIL.n69 VTAIL.n3 171.744
R497 VTAIL.n221 VTAIL.n155 171.744
R498 VTAIL.n214 VTAIL.n155 171.744
R499 VTAIL.n214 VTAIL.n213 171.744
R500 VTAIL.n213 VTAIL.n159 171.744
R501 VTAIL.n206 VTAIL.n159 171.744
R502 VTAIL.n206 VTAIL.n205 171.744
R503 VTAIL.n205 VTAIL.n163 171.744
R504 VTAIL.n198 VTAIL.n163 171.744
R505 VTAIL.n198 VTAIL.n197 171.744
R506 VTAIL.n197 VTAIL.n167 171.744
R507 VTAIL.n190 VTAIL.n167 171.744
R508 VTAIL.n190 VTAIL.n189 171.744
R509 VTAIL.n189 VTAIL.n171 171.744
R510 VTAIL.n182 VTAIL.n171 171.744
R511 VTAIL.n182 VTAIL.n181 171.744
R512 VTAIL.n181 VTAIL.n175 171.744
R513 VTAIL.n147 VTAIL.n81 171.744
R514 VTAIL.n140 VTAIL.n81 171.744
R515 VTAIL.n140 VTAIL.n139 171.744
R516 VTAIL.n139 VTAIL.n85 171.744
R517 VTAIL.n132 VTAIL.n85 171.744
R518 VTAIL.n132 VTAIL.n131 171.744
R519 VTAIL.n131 VTAIL.n89 171.744
R520 VTAIL.n124 VTAIL.n89 171.744
R521 VTAIL.n124 VTAIL.n123 171.744
R522 VTAIL.n123 VTAIL.n93 171.744
R523 VTAIL.n116 VTAIL.n93 171.744
R524 VTAIL.n116 VTAIL.n115 171.744
R525 VTAIL.n115 VTAIL.n97 171.744
R526 VTAIL.n108 VTAIL.n97 171.744
R527 VTAIL.n108 VTAIL.n107 171.744
R528 VTAIL.n107 VTAIL.n101 171.744
R529 VTAIL.t8 VTAIL.n245 85.8723
R530 VTAIL.t16 VTAIL.n23 85.8723
R531 VTAIL.t12 VTAIL.n175 85.8723
R532 VTAIL.t7 VTAIL.n101 85.8723
R533 VTAIL.n153 VTAIL.n152 57.9164
R534 VTAIL.n151 VTAIL.n150 57.9164
R535 VTAIL.n79 VTAIL.n78 57.9164
R536 VTAIL.n77 VTAIL.n76 57.9164
R537 VTAIL.n295 VTAIL.n294 57.9154
R538 VTAIL.n1 VTAIL.n0 57.9154
R539 VTAIL.n73 VTAIL.n72 57.9154
R540 VTAIL.n75 VTAIL.n74 57.9154
R541 VTAIL.n293 VTAIL.n292 33.7369
R542 VTAIL.n71 VTAIL.n70 33.7369
R543 VTAIL.n223 VTAIL.n222 33.7369
R544 VTAIL.n149 VTAIL.n148 33.7369
R545 VTAIL.n77 VTAIL.n75 29.0221
R546 VTAIL.n293 VTAIL.n223 26.1169
R547 VTAIL.n247 VTAIL.n246 16.3895
R548 VTAIL.n25 VTAIL.n24 16.3895
R549 VTAIL.n177 VTAIL.n176 16.3895
R550 VTAIL.n103 VTAIL.n102 16.3895
R551 VTAIL.n250 VTAIL.n249 12.8005
R552 VTAIL.n290 VTAIL.n224 12.8005
R553 VTAIL.n28 VTAIL.n27 12.8005
R554 VTAIL.n68 VTAIL.n2 12.8005
R555 VTAIL.n220 VTAIL.n154 12.8005
R556 VTAIL.n180 VTAIL.n179 12.8005
R557 VTAIL.n146 VTAIL.n80 12.8005
R558 VTAIL.n106 VTAIL.n105 12.8005
R559 VTAIL.n253 VTAIL.n244 12.0247
R560 VTAIL.n289 VTAIL.n226 12.0247
R561 VTAIL.n31 VTAIL.n22 12.0247
R562 VTAIL.n67 VTAIL.n4 12.0247
R563 VTAIL.n219 VTAIL.n156 12.0247
R564 VTAIL.n183 VTAIL.n174 12.0247
R565 VTAIL.n145 VTAIL.n82 12.0247
R566 VTAIL.n109 VTAIL.n100 12.0247
R567 VTAIL.n254 VTAIL.n242 11.249
R568 VTAIL.n286 VTAIL.n285 11.249
R569 VTAIL.n32 VTAIL.n20 11.249
R570 VTAIL.n64 VTAIL.n63 11.249
R571 VTAIL.n216 VTAIL.n215 11.249
R572 VTAIL.n184 VTAIL.n172 11.249
R573 VTAIL.n142 VTAIL.n141 11.249
R574 VTAIL.n110 VTAIL.n98 11.249
R575 VTAIL.n258 VTAIL.n257 10.4732
R576 VTAIL.n282 VTAIL.n228 10.4732
R577 VTAIL.n36 VTAIL.n35 10.4732
R578 VTAIL.n60 VTAIL.n6 10.4732
R579 VTAIL.n212 VTAIL.n158 10.4732
R580 VTAIL.n188 VTAIL.n187 10.4732
R581 VTAIL.n138 VTAIL.n84 10.4732
R582 VTAIL.n114 VTAIL.n113 10.4732
R583 VTAIL.n261 VTAIL.n240 9.69747
R584 VTAIL.n281 VTAIL.n230 9.69747
R585 VTAIL.n39 VTAIL.n18 9.69747
R586 VTAIL.n59 VTAIL.n8 9.69747
R587 VTAIL.n211 VTAIL.n160 9.69747
R588 VTAIL.n191 VTAIL.n170 9.69747
R589 VTAIL.n137 VTAIL.n86 9.69747
R590 VTAIL.n117 VTAIL.n96 9.69747
R591 VTAIL.n288 VTAIL.n224 9.45567
R592 VTAIL.n66 VTAIL.n2 9.45567
R593 VTAIL.n218 VTAIL.n154 9.45567
R594 VTAIL.n144 VTAIL.n80 9.45567
R595 VTAIL.n271 VTAIL.n270 9.3005
R596 VTAIL.n273 VTAIL.n272 9.3005
R597 VTAIL.n232 VTAIL.n231 9.3005
R598 VTAIL.n279 VTAIL.n278 9.3005
R599 VTAIL.n281 VTAIL.n280 9.3005
R600 VTAIL.n228 VTAIL.n227 9.3005
R601 VTAIL.n287 VTAIL.n286 9.3005
R602 VTAIL.n289 VTAIL.n288 9.3005
R603 VTAIL.n265 VTAIL.n264 9.3005
R604 VTAIL.n263 VTAIL.n262 9.3005
R605 VTAIL.n240 VTAIL.n239 9.3005
R606 VTAIL.n257 VTAIL.n256 9.3005
R607 VTAIL.n255 VTAIL.n254 9.3005
R608 VTAIL.n244 VTAIL.n243 9.3005
R609 VTAIL.n249 VTAIL.n248 9.3005
R610 VTAIL.n236 VTAIL.n235 9.3005
R611 VTAIL.n49 VTAIL.n48 9.3005
R612 VTAIL.n51 VTAIL.n50 9.3005
R613 VTAIL.n10 VTAIL.n9 9.3005
R614 VTAIL.n57 VTAIL.n56 9.3005
R615 VTAIL.n59 VTAIL.n58 9.3005
R616 VTAIL.n6 VTAIL.n5 9.3005
R617 VTAIL.n65 VTAIL.n64 9.3005
R618 VTAIL.n67 VTAIL.n66 9.3005
R619 VTAIL.n43 VTAIL.n42 9.3005
R620 VTAIL.n41 VTAIL.n40 9.3005
R621 VTAIL.n18 VTAIL.n17 9.3005
R622 VTAIL.n35 VTAIL.n34 9.3005
R623 VTAIL.n33 VTAIL.n32 9.3005
R624 VTAIL.n22 VTAIL.n21 9.3005
R625 VTAIL.n27 VTAIL.n26 9.3005
R626 VTAIL.n14 VTAIL.n13 9.3005
R627 VTAIL.n219 VTAIL.n218 9.3005
R628 VTAIL.n217 VTAIL.n216 9.3005
R629 VTAIL.n158 VTAIL.n157 9.3005
R630 VTAIL.n211 VTAIL.n210 9.3005
R631 VTAIL.n209 VTAIL.n208 9.3005
R632 VTAIL.n162 VTAIL.n161 9.3005
R633 VTAIL.n203 VTAIL.n202 9.3005
R634 VTAIL.n201 VTAIL.n200 9.3005
R635 VTAIL.n166 VTAIL.n165 9.3005
R636 VTAIL.n195 VTAIL.n194 9.3005
R637 VTAIL.n193 VTAIL.n192 9.3005
R638 VTAIL.n170 VTAIL.n169 9.3005
R639 VTAIL.n187 VTAIL.n186 9.3005
R640 VTAIL.n185 VTAIL.n184 9.3005
R641 VTAIL.n174 VTAIL.n173 9.3005
R642 VTAIL.n179 VTAIL.n178 9.3005
R643 VTAIL.n129 VTAIL.n128 9.3005
R644 VTAIL.n88 VTAIL.n87 9.3005
R645 VTAIL.n135 VTAIL.n134 9.3005
R646 VTAIL.n137 VTAIL.n136 9.3005
R647 VTAIL.n84 VTAIL.n83 9.3005
R648 VTAIL.n143 VTAIL.n142 9.3005
R649 VTAIL.n145 VTAIL.n144 9.3005
R650 VTAIL.n127 VTAIL.n126 9.3005
R651 VTAIL.n92 VTAIL.n91 9.3005
R652 VTAIL.n121 VTAIL.n120 9.3005
R653 VTAIL.n119 VTAIL.n118 9.3005
R654 VTAIL.n96 VTAIL.n95 9.3005
R655 VTAIL.n113 VTAIL.n112 9.3005
R656 VTAIL.n111 VTAIL.n110 9.3005
R657 VTAIL.n100 VTAIL.n99 9.3005
R658 VTAIL.n105 VTAIL.n104 9.3005
R659 VTAIL.n262 VTAIL.n238 8.92171
R660 VTAIL.n278 VTAIL.n277 8.92171
R661 VTAIL.n40 VTAIL.n16 8.92171
R662 VTAIL.n56 VTAIL.n55 8.92171
R663 VTAIL.n208 VTAIL.n207 8.92171
R664 VTAIL.n192 VTAIL.n168 8.92171
R665 VTAIL.n134 VTAIL.n133 8.92171
R666 VTAIL.n118 VTAIL.n94 8.92171
R667 VTAIL.n266 VTAIL.n265 8.14595
R668 VTAIL.n274 VTAIL.n232 8.14595
R669 VTAIL.n44 VTAIL.n43 8.14595
R670 VTAIL.n52 VTAIL.n10 8.14595
R671 VTAIL.n204 VTAIL.n162 8.14595
R672 VTAIL.n196 VTAIL.n195 8.14595
R673 VTAIL.n130 VTAIL.n88 8.14595
R674 VTAIL.n122 VTAIL.n121 8.14595
R675 VTAIL.n269 VTAIL.n236 7.3702
R676 VTAIL.n273 VTAIL.n234 7.3702
R677 VTAIL.n47 VTAIL.n14 7.3702
R678 VTAIL.n51 VTAIL.n12 7.3702
R679 VTAIL.n203 VTAIL.n164 7.3702
R680 VTAIL.n199 VTAIL.n166 7.3702
R681 VTAIL.n129 VTAIL.n90 7.3702
R682 VTAIL.n125 VTAIL.n92 7.3702
R683 VTAIL.n270 VTAIL.n269 6.59444
R684 VTAIL.n270 VTAIL.n234 6.59444
R685 VTAIL.n48 VTAIL.n47 6.59444
R686 VTAIL.n48 VTAIL.n12 6.59444
R687 VTAIL.n200 VTAIL.n164 6.59444
R688 VTAIL.n200 VTAIL.n199 6.59444
R689 VTAIL.n126 VTAIL.n90 6.59444
R690 VTAIL.n126 VTAIL.n125 6.59444
R691 VTAIL.n266 VTAIL.n236 5.81868
R692 VTAIL.n274 VTAIL.n273 5.81868
R693 VTAIL.n44 VTAIL.n14 5.81868
R694 VTAIL.n52 VTAIL.n51 5.81868
R695 VTAIL.n204 VTAIL.n203 5.81868
R696 VTAIL.n196 VTAIL.n166 5.81868
R697 VTAIL.n130 VTAIL.n129 5.81868
R698 VTAIL.n122 VTAIL.n92 5.81868
R699 VTAIL.n265 VTAIL.n238 5.04292
R700 VTAIL.n277 VTAIL.n232 5.04292
R701 VTAIL.n43 VTAIL.n16 5.04292
R702 VTAIL.n55 VTAIL.n10 5.04292
R703 VTAIL.n207 VTAIL.n162 5.04292
R704 VTAIL.n195 VTAIL.n168 5.04292
R705 VTAIL.n133 VTAIL.n88 5.04292
R706 VTAIL.n121 VTAIL.n94 5.04292
R707 VTAIL.n262 VTAIL.n261 4.26717
R708 VTAIL.n278 VTAIL.n230 4.26717
R709 VTAIL.n40 VTAIL.n39 4.26717
R710 VTAIL.n56 VTAIL.n8 4.26717
R711 VTAIL.n208 VTAIL.n160 4.26717
R712 VTAIL.n192 VTAIL.n191 4.26717
R713 VTAIL.n134 VTAIL.n86 4.26717
R714 VTAIL.n118 VTAIL.n117 4.26717
R715 VTAIL.n248 VTAIL.n247 3.70982
R716 VTAIL.n26 VTAIL.n25 3.70982
R717 VTAIL.n178 VTAIL.n177 3.70982
R718 VTAIL.n104 VTAIL.n103 3.70982
R719 VTAIL.n258 VTAIL.n240 3.49141
R720 VTAIL.n282 VTAIL.n281 3.49141
R721 VTAIL.n36 VTAIL.n18 3.49141
R722 VTAIL.n60 VTAIL.n59 3.49141
R723 VTAIL.n212 VTAIL.n211 3.49141
R724 VTAIL.n188 VTAIL.n170 3.49141
R725 VTAIL.n138 VTAIL.n137 3.49141
R726 VTAIL.n114 VTAIL.n96 3.49141
R727 VTAIL.n79 VTAIL.n77 2.90567
R728 VTAIL.n149 VTAIL.n79 2.90567
R729 VTAIL.n153 VTAIL.n151 2.90567
R730 VTAIL.n223 VTAIL.n153 2.90567
R731 VTAIL.n75 VTAIL.n73 2.90567
R732 VTAIL.n73 VTAIL.n71 2.90567
R733 VTAIL.n295 VTAIL.n293 2.90567
R734 VTAIL.n257 VTAIL.n242 2.71565
R735 VTAIL.n285 VTAIL.n228 2.71565
R736 VTAIL.n35 VTAIL.n20 2.71565
R737 VTAIL.n63 VTAIL.n6 2.71565
R738 VTAIL.n215 VTAIL.n158 2.71565
R739 VTAIL.n187 VTAIL.n172 2.71565
R740 VTAIL.n141 VTAIL.n84 2.71565
R741 VTAIL.n113 VTAIL.n98 2.71565
R742 VTAIL.n294 VTAIL.t0 2.58436
R743 VTAIL.n294 VTAIL.t2 2.58436
R744 VTAIL.n0 VTAIL.t4 2.58436
R745 VTAIL.n0 VTAIL.t1 2.58436
R746 VTAIL.n72 VTAIL.t15 2.58436
R747 VTAIL.n72 VTAIL.t18 2.58436
R748 VTAIL.n74 VTAIL.t11 2.58436
R749 VTAIL.n74 VTAIL.t9 2.58436
R750 VTAIL.n152 VTAIL.t17 2.58436
R751 VTAIL.n152 VTAIL.t13 2.58436
R752 VTAIL.n150 VTAIL.t10 2.58436
R753 VTAIL.n150 VTAIL.t14 2.58436
R754 VTAIL.n78 VTAIL.t6 2.58436
R755 VTAIL.n78 VTAIL.t3 2.58436
R756 VTAIL.n76 VTAIL.t19 2.58436
R757 VTAIL.n76 VTAIL.t5 2.58436
R758 VTAIL VTAIL.n1 2.23757
R759 VTAIL.n254 VTAIL.n253 1.93989
R760 VTAIL.n286 VTAIL.n226 1.93989
R761 VTAIL.n32 VTAIL.n31 1.93989
R762 VTAIL.n64 VTAIL.n4 1.93989
R763 VTAIL.n216 VTAIL.n156 1.93989
R764 VTAIL.n184 VTAIL.n183 1.93989
R765 VTAIL.n142 VTAIL.n82 1.93989
R766 VTAIL.n110 VTAIL.n109 1.93989
R767 VTAIL.n151 VTAIL.n149 1.92291
R768 VTAIL.n71 VTAIL.n1 1.92291
R769 VTAIL.n250 VTAIL.n244 1.16414
R770 VTAIL.n290 VTAIL.n289 1.16414
R771 VTAIL.n28 VTAIL.n22 1.16414
R772 VTAIL.n68 VTAIL.n67 1.16414
R773 VTAIL.n220 VTAIL.n219 1.16414
R774 VTAIL.n180 VTAIL.n174 1.16414
R775 VTAIL.n146 VTAIL.n145 1.16414
R776 VTAIL.n106 VTAIL.n100 1.16414
R777 VTAIL VTAIL.n295 0.668603
R778 VTAIL.n249 VTAIL.n246 0.388379
R779 VTAIL.n292 VTAIL.n224 0.388379
R780 VTAIL.n27 VTAIL.n24 0.388379
R781 VTAIL.n70 VTAIL.n2 0.388379
R782 VTAIL.n222 VTAIL.n154 0.388379
R783 VTAIL.n179 VTAIL.n176 0.388379
R784 VTAIL.n148 VTAIL.n80 0.388379
R785 VTAIL.n105 VTAIL.n102 0.388379
R786 VTAIL.n248 VTAIL.n243 0.155672
R787 VTAIL.n255 VTAIL.n243 0.155672
R788 VTAIL.n256 VTAIL.n255 0.155672
R789 VTAIL.n256 VTAIL.n239 0.155672
R790 VTAIL.n263 VTAIL.n239 0.155672
R791 VTAIL.n264 VTAIL.n263 0.155672
R792 VTAIL.n264 VTAIL.n235 0.155672
R793 VTAIL.n271 VTAIL.n235 0.155672
R794 VTAIL.n272 VTAIL.n271 0.155672
R795 VTAIL.n272 VTAIL.n231 0.155672
R796 VTAIL.n279 VTAIL.n231 0.155672
R797 VTAIL.n280 VTAIL.n279 0.155672
R798 VTAIL.n280 VTAIL.n227 0.155672
R799 VTAIL.n287 VTAIL.n227 0.155672
R800 VTAIL.n288 VTAIL.n287 0.155672
R801 VTAIL.n26 VTAIL.n21 0.155672
R802 VTAIL.n33 VTAIL.n21 0.155672
R803 VTAIL.n34 VTAIL.n33 0.155672
R804 VTAIL.n34 VTAIL.n17 0.155672
R805 VTAIL.n41 VTAIL.n17 0.155672
R806 VTAIL.n42 VTAIL.n41 0.155672
R807 VTAIL.n42 VTAIL.n13 0.155672
R808 VTAIL.n49 VTAIL.n13 0.155672
R809 VTAIL.n50 VTAIL.n49 0.155672
R810 VTAIL.n50 VTAIL.n9 0.155672
R811 VTAIL.n57 VTAIL.n9 0.155672
R812 VTAIL.n58 VTAIL.n57 0.155672
R813 VTAIL.n58 VTAIL.n5 0.155672
R814 VTAIL.n65 VTAIL.n5 0.155672
R815 VTAIL.n66 VTAIL.n65 0.155672
R816 VTAIL.n218 VTAIL.n217 0.155672
R817 VTAIL.n217 VTAIL.n157 0.155672
R818 VTAIL.n210 VTAIL.n157 0.155672
R819 VTAIL.n210 VTAIL.n209 0.155672
R820 VTAIL.n209 VTAIL.n161 0.155672
R821 VTAIL.n202 VTAIL.n161 0.155672
R822 VTAIL.n202 VTAIL.n201 0.155672
R823 VTAIL.n201 VTAIL.n165 0.155672
R824 VTAIL.n194 VTAIL.n165 0.155672
R825 VTAIL.n194 VTAIL.n193 0.155672
R826 VTAIL.n193 VTAIL.n169 0.155672
R827 VTAIL.n186 VTAIL.n169 0.155672
R828 VTAIL.n186 VTAIL.n185 0.155672
R829 VTAIL.n185 VTAIL.n173 0.155672
R830 VTAIL.n178 VTAIL.n173 0.155672
R831 VTAIL.n144 VTAIL.n143 0.155672
R832 VTAIL.n143 VTAIL.n83 0.155672
R833 VTAIL.n136 VTAIL.n83 0.155672
R834 VTAIL.n136 VTAIL.n135 0.155672
R835 VTAIL.n135 VTAIL.n87 0.155672
R836 VTAIL.n128 VTAIL.n87 0.155672
R837 VTAIL.n128 VTAIL.n127 0.155672
R838 VTAIL.n127 VTAIL.n91 0.155672
R839 VTAIL.n120 VTAIL.n91 0.155672
R840 VTAIL.n120 VTAIL.n119 0.155672
R841 VTAIL.n119 VTAIL.n95 0.155672
R842 VTAIL.n112 VTAIL.n95 0.155672
R843 VTAIL.n112 VTAIL.n111 0.155672
R844 VTAIL.n111 VTAIL.n99 0.155672
R845 VTAIL.n104 VTAIL.n99 0.155672
R846 VN.n90 VN.n89 161.3
R847 VN.n88 VN.n47 161.3
R848 VN.n87 VN.n86 161.3
R849 VN.n85 VN.n48 161.3
R850 VN.n84 VN.n83 161.3
R851 VN.n82 VN.n49 161.3
R852 VN.n80 VN.n79 161.3
R853 VN.n78 VN.n50 161.3
R854 VN.n77 VN.n76 161.3
R855 VN.n75 VN.n51 161.3
R856 VN.n74 VN.n73 161.3
R857 VN.n72 VN.n52 161.3
R858 VN.n71 VN.n70 161.3
R859 VN.n68 VN.n53 161.3
R860 VN.n67 VN.n66 161.3
R861 VN.n65 VN.n54 161.3
R862 VN.n64 VN.n63 161.3
R863 VN.n62 VN.n55 161.3
R864 VN.n61 VN.n60 161.3
R865 VN.n59 VN.n56 161.3
R866 VN.n44 VN.n43 161.3
R867 VN.n42 VN.n1 161.3
R868 VN.n41 VN.n40 161.3
R869 VN.n39 VN.n2 161.3
R870 VN.n38 VN.n37 161.3
R871 VN.n36 VN.n3 161.3
R872 VN.n34 VN.n33 161.3
R873 VN.n32 VN.n4 161.3
R874 VN.n31 VN.n30 161.3
R875 VN.n29 VN.n5 161.3
R876 VN.n28 VN.n27 161.3
R877 VN.n26 VN.n6 161.3
R878 VN.n25 VN.n24 161.3
R879 VN.n22 VN.n7 161.3
R880 VN.n21 VN.n20 161.3
R881 VN.n19 VN.n8 161.3
R882 VN.n18 VN.n17 161.3
R883 VN.n16 VN.n9 161.3
R884 VN.n15 VN.n14 161.3
R885 VN.n13 VN.n10 161.3
R886 VN.n58 VN.t3 131.565
R887 VN.n12 VN.t5 131.565
R888 VN.n11 VN.t0 99.7301
R889 VN.n23 VN.t6 99.7301
R890 VN.n35 VN.t2 99.7301
R891 VN.n0 VN.t9 99.7301
R892 VN.n57 VN.t7 99.7301
R893 VN.n69 VN.t8 99.7301
R894 VN.n81 VN.t1 99.7301
R895 VN.n46 VN.t4 99.7301
R896 VN.n12 VN.n11 68.2679
R897 VN.n58 VN.n57 68.2679
R898 VN.n45 VN.n0 66.1456
R899 VN.n91 VN.n46 66.1456
R900 VN.n41 VN.n2 56.5617
R901 VN.n87 VN.n48 56.5617
R902 VN VN.n91 56.305
R903 VN.n17 VN.n8 46.874
R904 VN.n29 VN.n28 46.874
R905 VN.n63 VN.n54 46.874
R906 VN.n75 VN.n74 46.874
R907 VN.n17 VN.n16 34.28
R908 VN.n30 VN.n29 34.28
R909 VN.n63 VN.n62 34.28
R910 VN.n76 VN.n75 34.28
R911 VN.n15 VN.n10 24.5923
R912 VN.n16 VN.n15 24.5923
R913 VN.n21 VN.n8 24.5923
R914 VN.n22 VN.n21 24.5923
R915 VN.n24 VN.n6 24.5923
R916 VN.n28 VN.n6 24.5923
R917 VN.n30 VN.n4 24.5923
R918 VN.n34 VN.n4 24.5923
R919 VN.n37 VN.n36 24.5923
R920 VN.n37 VN.n2 24.5923
R921 VN.n42 VN.n41 24.5923
R922 VN.n43 VN.n42 24.5923
R923 VN.n62 VN.n61 24.5923
R924 VN.n61 VN.n56 24.5923
R925 VN.n74 VN.n52 24.5923
R926 VN.n70 VN.n52 24.5923
R927 VN.n68 VN.n67 24.5923
R928 VN.n67 VN.n54 24.5923
R929 VN.n83 VN.n48 24.5923
R930 VN.n83 VN.n82 24.5923
R931 VN.n80 VN.n50 24.5923
R932 VN.n76 VN.n50 24.5923
R933 VN.n89 VN.n88 24.5923
R934 VN.n88 VN.n87 24.5923
R935 VN.n43 VN.n0 24.1005
R936 VN.n89 VN.n46 24.1005
R937 VN.n36 VN.n35 18.6903
R938 VN.n82 VN.n81 18.6903
R939 VN.n23 VN.n22 12.2964
R940 VN.n24 VN.n23 12.2964
R941 VN.n70 VN.n69 12.2964
R942 VN.n69 VN.n68 12.2964
R943 VN.n11 VN.n10 5.90254
R944 VN.n35 VN.n34 5.90254
R945 VN.n57 VN.n56 5.90254
R946 VN.n81 VN.n80 5.90254
R947 VN.n13 VN.n12 5.2507
R948 VN.n59 VN.n58 5.2507
R949 VN.n91 VN.n90 0.354861
R950 VN.n45 VN.n44 0.354861
R951 VN VN.n45 0.267071
R952 VN.n90 VN.n47 0.189894
R953 VN.n86 VN.n47 0.189894
R954 VN.n86 VN.n85 0.189894
R955 VN.n85 VN.n84 0.189894
R956 VN.n84 VN.n49 0.189894
R957 VN.n79 VN.n49 0.189894
R958 VN.n79 VN.n78 0.189894
R959 VN.n78 VN.n77 0.189894
R960 VN.n77 VN.n51 0.189894
R961 VN.n73 VN.n51 0.189894
R962 VN.n73 VN.n72 0.189894
R963 VN.n72 VN.n71 0.189894
R964 VN.n71 VN.n53 0.189894
R965 VN.n66 VN.n53 0.189894
R966 VN.n66 VN.n65 0.189894
R967 VN.n65 VN.n64 0.189894
R968 VN.n64 VN.n55 0.189894
R969 VN.n60 VN.n55 0.189894
R970 VN.n60 VN.n59 0.189894
R971 VN.n14 VN.n13 0.189894
R972 VN.n14 VN.n9 0.189894
R973 VN.n18 VN.n9 0.189894
R974 VN.n19 VN.n18 0.189894
R975 VN.n20 VN.n19 0.189894
R976 VN.n20 VN.n7 0.189894
R977 VN.n25 VN.n7 0.189894
R978 VN.n26 VN.n25 0.189894
R979 VN.n27 VN.n26 0.189894
R980 VN.n27 VN.n5 0.189894
R981 VN.n31 VN.n5 0.189894
R982 VN.n32 VN.n31 0.189894
R983 VN.n33 VN.n32 0.189894
R984 VN.n33 VN.n3 0.189894
R985 VN.n38 VN.n3 0.189894
R986 VN.n39 VN.n38 0.189894
R987 VN.n40 VN.n39 0.189894
R988 VN.n40 VN.n1 0.189894
R989 VN.n44 VN.n1 0.189894
R990 VDD2.n141 VDD2.n140 756.745
R991 VDD2.n68 VDD2.n67 756.745
R992 VDD2.n140 VDD2.n139 585
R993 VDD2.n75 VDD2.n74 585
R994 VDD2.n134 VDD2.n133 585
R995 VDD2.n132 VDD2.n131 585
R996 VDD2.n79 VDD2.n78 585
R997 VDD2.n126 VDD2.n125 585
R998 VDD2.n124 VDD2.n123 585
R999 VDD2.n83 VDD2.n82 585
R1000 VDD2.n118 VDD2.n117 585
R1001 VDD2.n116 VDD2.n115 585
R1002 VDD2.n87 VDD2.n86 585
R1003 VDD2.n110 VDD2.n109 585
R1004 VDD2.n108 VDD2.n107 585
R1005 VDD2.n91 VDD2.n90 585
R1006 VDD2.n102 VDD2.n101 585
R1007 VDD2.n100 VDD2.n99 585
R1008 VDD2.n95 VDD2.n94 585
R1009 VDD2.n22 VDD2.n21 585
R1010 VDD2.n27 VDD2.n26 585
R1011 VDD2.n29 VDD2.n28 585
R1012 VDD2.n18 VDD2.n17 585
R1013 VDD2.n35 VDD2.n34 585
R1014 VDD2.n37 VDD2.n36 585
R1015 VDD2.n14 VDD2.n13 585
R1016 VDD2.n43 VDD2.n42 585
R1017 VDD2.n45 VDD2.n44 585
R1018 VDD2.n10 VDD2.n9 585
R1019 VDD2.n51 VDD2.n50 585
R1020 VDD2.n53 VDD2.n52 585
R1021 VDD2.n6 VDD2.n5 585
R1022 VDD2.n59 VDD2.n58 585
R1023 VDD2.n61 VDD2.n60 585
R1024 VDD2.n2 VDD2.n1 585
R1025 VDD2.n67 VDD2.n66 585
R1026 VDD2.n96 VDD2.t5 327.466
R1027 VDD2.n23 VDD2.t4 327.466
R1028 VDD2.n140 VDD2.n74 171.744
R1029 VDD2.n133 VDD2.n74 171.744
R1030 VDD2.n133 VDD2.n132 171.744
R1031 VDD2.n132 VDD2.n78 171.744
R1032 VDD2.n125 VDD2.n78 171.744
R1033 VDD2.n125 VDD2.n124 171.744
R1034 VDD2.n124 VDD2.n82 171.744
R1035 VDD2.n117 VDD2.n82 171.744
R1036 VDD2.n117 VDD2.n116 171.744
R1037 VDD2.n116 VDD2.n86 171.744
R1038 VDD2.n109 VDD2.n86 171.744
R1039 VDD2.n109 VDD2.n108 171.744
R1040 VDD2.n108 VDD2.n90 171.744
R1041 VDD2.n101 VDD2.n90 171.744
R1042 VDD2.n101 VDD2.n100 171.744
R1043 VDD2.n100 VDD2.n94 171.744
R1044 VDD2.n27 VDD2.n21 171.744
R1045 VDD2.n28 VDD2.n27 171.744
R1046 VDD2.n28 VDD2.n17 171.744
R1047 VDD2.n35 VDD2.n17 171.744
R1048 VDD2.n36 VDD2.n35 171.744
R1049 VDD2.n36 VDD2.n13 171.744
R1050 VDD2.n43 VDD2.n13 171.744
R1051 VDD2.n44 VDD2.n43 171.744
R1052 VDD2.n44 VDD2.n9 171.744
R1053 VDD2.n51 VDD2.n9 171.744
R1054 VDD2.n52 VDD2.n51 171.744
R1055 VDD2.n52 VDD2.n5 171.744
R1056 VDD2.n59 VDD2.n5 171.744
R1057 VDD2.n60 VDD2.n59 171.744
R1058 VDD2.n60 VDD2.n1 171.744
R1059 VDD2.n67 VDD2.n1 171.744
R1060 VDD2.t5 VDD2.n94 85.8723
R1061 VDD2.t4 VDD2.n21 85.8723
R1062 VDD2.n72 VDD2.n71 76.7177
R1063 VDD2 VDD2.n145 76.7148
R1064 VDD2.n144 VDD2.n143 74.5952
R1065 VDD2.n70 VDD2.n69 74.5942
R1066 VDD2.n70 VDD2.n68 53.3208
R1067 VDD2.n142 VDD2.n141 50.4157
R1068 VDD2.n142 VDD2.n72 48.3597
R1069 VDD2.n96 VDD2.n95 16.3895
R1070 VDD2.n23 VDD2.n22 16.3895
R1071 VDD2.n139 VDD2.n73 12.8005
R1072 VDD2.n99 VDD2.n98 12.8005
R1073 VDD2.n26 VDD2.n25 12.8005
R1074 VDD2.n66 VDD2.n0 12.8005
R1075 VDD2.n138 VDD2.n75 12.0247
R1076 VDD2.n102 VDD2.n93 12.0247
R1077 VDD2.n29 VDD2.n20 12.0247
R1078 VDD2.n65 VDD2.n2 12.0247
R1079 VDD2.n135 VDD2.n134 11.249
R1080 VDD2.n103 VDD2.n91 11.249
R1081 VDD2.n30 VDD2.n18 11.249
R1082 VDD2.n62 VDD2.n61 11.249
R1083 VDD2.n131 VDD2.n77 10.4732
R1084 VDD2.n107 VDD2.n106 10.4732
R1085 VDD2.n34 VDD2.n33 10.4732
R1086 VDD2.n58 VDD2.n4 10.4732
R1087 VDD2.n130 VDD2.n79 9.69747
R1088 VDD2.n110 VDD2.n89 9.69747
R1089 VDD2.n37 VDD2.n16 9.69747
R1090 VDD2.n57 VDD2.n6 9.69747
R1091 VDD2.n137 VDD2.n73 9.45567
R1092 VDD2.n64 VDD2.n0 9.45567
R1093 VDD2.n122 VDD2.n121 9.3005
R1094 VDD2.n81 VDD2.n80 9.3005
R1095 VDD2.n128 VDD2.n127 9.3005
R1096 VDD2.n130 VDD2.n129 9.3005
R1097 VDD2.n77 VDD2.n76 9.3005
R1098 VDD2.n136 VDD2.n135 9.3005
R1099 VDD2.n138 VDD2.n137 9.3005
R1100 VDD2.n120 VDD2.n119 9.3005
R1101 VDD2.n85 VDD2.n84 9.3005
R1102 VDD2.n114 VDD2.n113 9.3005
R1103 VDD2.n112 VDD2.n111 9.3005
R1104 VDD2.n89 VDD2.n88 9.3005
R1105 VDD2.n106 VDD2.n105 9.3005
R1106 VDD2.n104 VDD2.n103 9.3005
R1107 VDD2.n93 VDD2.n92 9.3005
R1108 VDD2.n98 VDD2.n97 9.3005
R1109 VDD2.n47 VDD2.n46 9.3005
R1110 VDD2.n49 VDD2.n48 9.3005
R1111 VDD2.n8 VDD2.n7 9.3005
R1112 VDD2.n55 VDD2.n54 9.3005
R1113 VDD2.n57 VDD2.n56 9.3005
R1114 VDD2.n4 VDD2.n3 9.3005
R1115 VDD2.n63 VDD2.n62 9.3005
R1116 VDD2.n65 VDD2.n64 9.3005
R1117 VDD2.n41 VDD2.n40 9.3005
R1118 VDD2.n39 VDD2.n38 9.3005
R1119 VDD2.n16 VDD2.n15 9.3005
R1120 VDD2.n33 VDD2.n32 9.3005
R1121 VDD2.n31 VDD2.n30 9.3005
R1122 VDD2.n20 VDD2.n19 9.3005
R1123 VDD2.n25 VDD2.n24 9.3005
R1124 VDD2.n12 VDD2.n11 9.3005
R1125 VDD2.n127 VDD2.n126 8.92171
R1126 VDD2.n111 VDD2.n87 8.92171
R1127 VDD2.n38 VDD2.n14 8.92171
R1128 VDD2.n54 VDD2.n53 8.92171
R1129 VDD2.n123 VDD2.n81 8.14595
R1130 VDD2.n115 VDD2.n114 8.14595
R1131 VDD2.n42 VDD2.n41 8.14595
R1132 VDD2.n50 VDD2.n8 8.14595
R1133 VDD2.n122 VDD2.n83 7.3702
R1134 VDD2.n118 VDD2.n85 7.3702
R1135 VDD2.n45 VDD2.n12 7.3702
R1136 VDD2.n49 VDD2.n10 7.3702
R1137 VDD2.n119 VDD2.n83 6.59444
R1138 VDD2.n119 VDD2.n118 6.59444
R1139 VDD2.n46 VDD2.n45 6.59444
R1140 VDD2.n46 VDD2.n10 6.59444
R1141 VDD2.n123 VDD2.n122 5.81868
R1142 VDD2.n115 VDD2.n85 5.81868
R1143 VDD2.n42 VDD2.n12 5.81868
R1144 VDD2.n50 VDD2.n49 5.81868
R1145 VDD2.n126 VDD2.n81 5.04292
R1146 VDD2.n114 VDD2.n87 5.04292
R1147 VDD2.n41 VDD2.n14 5.04292
R1148 VDD2.n53 VDD2.n8 5.04292
R1149 VDD2.n127 VDD2.n79 4.26717
R1150 VDD2.n111 VDD2.n110 4.26717
R1151 VDD2.n38 VDD2.n37 4.26717
R1152 VDD2.n54 VDD2.n6 4.26717
R1153 VDD2.n97 VDD2.n96 3.70982
R1154 VDD2.n24 VDD2.n23 3.70982
R1155 VDD2.n131 VDD2.n130 3.49141
R1156 VDD2.n107 VDD2.n89 3.49141
R1157 VDD2.n34 VDD2.n16 3.49141
R1158 VDD2.n58 VDD2.n57 3.49141
R1159 VDD2.n144 VDD2.n142 2.90567
R1160 VDD2.n134 VDD2.n77 2.71565
R1161 VDD2.n106 VDD2.n91 2.71565
R1162 VDD2.n33 VDD2.n18 2.71565
R1163 VDD2.n61 VDD2.n4 2.71565
R1164 VDD2.n145 VDD2.t2 2.58436
R1165 VDD2.n145 VDD2.t6 2.58436
R1166 VDD2.n143 VDD2.t8 2.58436
R1167 VDD2.n143 VDD2.t1 2.58436
R1168 VDD2.n71 VDD2.t7 2.58436
R1169 VDD2.n71 VDD2.t0 2.58436
R1170 VDD2.n69 VDD2.t9 2.58436
R1171 VDD2.n69 VDD2.t3 2.58436
R1172 VDD2.n135 VDD2.n75 1.93989
R1173 VDD2.n103 VDD2.n102 1.93989
R1174 VDD2.n30 VDD2.n29 1.93989
R1175 VDD2.n62 VDD2.n2 1.93989
R1176 VDD2.n139 VDD2.n138 1.16414
R1177 VDD2.n99 VDD2.n93 1.16414
R1178 VDD2.n26 VDD2.n20 1.16414
R1179 VDD2.n66 VDD2.n65 1.16414
R1180 VDD2 VDD2.n144 0.784983
R1181 VDD2.n72 VDD2.n70 0.671447
R1182 VDD2.n141 VDD2.n73 0.388379
R1183 VDD2.n98 VDD2.n95 0.388379
R1184 VDD2.n25 VDD2.n22 0.388379
R1185 VDD2.n68 VDD2.n0 0.388379
R1186 VDD2.n137 VDD2.n136 0.155672
R1187 VDD2.n136 VDD2.n76 0.155672
R1188 VDD2.n129 VDD2.n76 0.155672
R1189 VDD2.n129 VDD2.n128 0.155672
R1190 VDD2.n128 VDD2.n80 0.155672
R1191 VDD2.n121 VDD2.n80 0.155672
R1192 VDD2.n121 VDD2.n120 0.155672
R1193 VDD2.n120 VDD2.n84 0.155672
R1194 VDD2.n113 VDD2.n84 0.155672
R1195 VDD2.n113 VDD2.n112 0.155672
R1196 VDD2.n112 VDD2.n88 0.155672
R1197 VDD2.n105 VDD2.n88 0.155672
R1198 VDD2.n105 VDD2.n104 0.155672
R1199 VDD2.n104 VDD2.n92 0.155672
R1200 VDD2.n97 VDD2.n92 0.155672
R1201 VDD2.n24 VDD2.n19 0.155672
R1202 VDD2.n31 VDD2.n19 0.155672
R1203 VDD2.n32 VDD2.n31 0.155672
R1204 VDD2.n32 VDD2.n15 0.155672
R1205 VDD2.n39 VDD2.n15 0.155672
R1206 VDD2.n40 VDD2.n39 0.155672
R1207 VDD2.n40 VDD2.n11 0.155672
R1208 VDD2.n47 VDD2.n11 0.155672
R1209 VDD2.n48 VDD2.n47 0.155672
R1210 VDD2.n48 VDD2.n7 0.155672
R1211 VDD2.n55 VDD2.n7 0.155672
R1212 VDD2.n56 VDD2.n55 0.155672
R1213 VDD2.n56 VDD2.n3 0.155672
R1214 VDD2.n63 VDD2.n3 0.155672
R1215 VDD2.n64 VDD2.n63 0.155672
R1216 B.n485 B.n156 585
R1217 B.n484 B.n483 585
R1218 B.n482 B.n157 585
R1219 B.n481 B.n480 585
R1220 B.n479 B.n158 585
R1221 B.n478 B.n477 585
R1222 B.n476 B.n159 585
R1223 B.n475 B.n474 585
R1224 B.n473 B.n160 585
R1225 B.n472 B.n471 585
R1226 B.n470 B.n161 585
R1227 B.n469 B.n468 585
R1228 B.n467 B.n162 585
R1229 B.n466 B.n465 585
R1230 B.n464 B.n163 585
R1231 B.n463 B.n462 585
R1232 B.n461 B.n164 585
R1233 B.n460 B.n459 585
R1234 B.n458 B.n165 585
R1235 B.n457 B.n456 585
R1236 B.n455 B.n166 585
R1237 B.n454 B.n453 585
R1238 B.n452 B.n167 585
R1239 B.n451 B.n450 585
R1240 B.n449 B.n168 585
R1241 B.n448 B.n447 585
R1242 B.n446 B.n169 585
R1243 B.n445 B.n444 585
R1244 B.n443 B.n170 585
R1245 B.n442 B.n441 585
R1246 B.n440 B.n171 585
R1247 B.n439 B.n438 585
R1248 B.n437 B.n172 585
R1249 B.n436 B.n435 585
R1250 B.n434 B.n173 585
R1251 B.n433 B.n432 585
R1252 B.n431 B.n174 585
R1253 B.n430 B.n429 585
R1254 B.n428 B.n175 585
R1255 B.n427 B.n426 585
R1256 B.n425 B.n176 585
R1257 B.n424 B.n423 585
R1258 B.n422 B.n177 585
R1259 B.n420 B.n419 585
R1260 B.n418 B.n180 585
R1261 B.n417 B.n416 585
R1262 B.n415 B.n181 585
R1263 B.n414 B.n413 585
R1264 B.n412 B.n182 585
R1265 B.n411 B.n410 585
R1266 B.n409 B.n183 585
R1267 B.n408 B.n407 585
R1268 B.n406 B.n184 585
R1269 B.n405 B.n404 585
R1270 B.n400 B.n185 585
R1271 B.n399 B.n398 585
R1272 B.n397 B.n186 585
R1273 B.n396 B.n395 585
R1274 B.n394 B.n187 585
R1275 B.n393 B.n392 585
R1276 B.n391 B.n188 585
R1277 B.n390 B.n389 585
R1278 B.n388 B.n189 585
R1279 B.n387 B.n386 585
R1280 B.n385 B.n190 585
R1281 B.n384 B.n383 585
R1282 B.n382 B.n191 585
R1283 B.n381 B.n380 585
R1284 B.n379 B.n192 585
R1285 B.n378 B.n377 585
R1286 B.n376 B.n193 585
R1287 B.n375 B.n374 585
R1288 B.n373 B.n194 585
R1289 B.n372 B.n371 585
R1290 B.n370 B.n195 585
R1291 B.n369 B.n368 585
R1292 B.n367 B.n196 585
R1293 B.n366 B.n365 585
R1294 B.n364 B.n197 585
R1295 B.n363 B.n362 585
R1296 B.n361 B.n198 585
R1297 B.n360 B.n359 585
R1298 B.n358 B.n199 585
R1299 B.n357 B.n356 585
R1300 B.n355 B.n200 585
R1301 B.n354 B.n353 585
R1302 B.n352 B.n201 585
R1303 B.n351 B.n350 585
R1304 B.n349 B.n202 585
R1305 B.n348 B.n347 585
R1306 B.n346 B.n203 585
R1307 B.n345 B.n344 585
R1308 B.n343 B.n204 585
R1309 B.n342 B.n341 585
R1310 B.n340 B.n205 585
R1311 B.n339 B.n338 585
R1312 B.n487 B.n486 585
R1313 B.n488 B.n155 585
R1314 B.n490 B.n489 585
R1315 B.n491 B.n154 585
R1316 B.n493 B.n492 585
R1317 B.n494 B.n153 585
R1318 B.n496 B.n495 585
R1319 B.n497 B.n152 585
R1320 B.n499 B.n498 585
R1321 B.n500 B.n151 585
R1322 B.n502 B.n501 585
R1323 B.n503 B.n150 585
R1324 B.n505 B.n504 585
R1325 B.n506 B.n149 585
R1326 B.n508 B.n507 585
R1327 B.n509 B.n148 585
R1328 B.n511 B.n510 585
R1329 B.n512 B.n147 585
R1330 B.n514 B.n513 585
R1331 B.n515 B.n146 585
R1332 B.n517 B.n516 585
R1333 B.n518 B.n145 585
R1334 B.n520 B.n519 585
R1335 B.n521 B.n144 585
R1336 B.n523 B.n522 585
R1337 B.n524 B.n143 585
R1338 B.n526 B.n525 585
R1339 B.n527 B.n142 585
R1340 B.n529 B.n528 585
R1341 B.n530 B.n141 585
R1342 B.n532 B.n531 585
R1343 B.n533 B.n140 585
R1344 B.n535 B.n534 585
R1345 B.n536 B.n139 585
R1346 B.n538 B.n537 585
R1347 B.n539 B.n138 585
R1348 B.n541 B.n540 585
R1349 B.n542 B.n137 585
R1350 B.n544 B.n543 585
R1351 B.n545 B.n136 585
R1352 B.n547 B.n546 585
R1353 B.n548 B.n135 585
R1354 B.n550 B.n549 585
R1355 B.n551 B.n134 585
R1356 B.n553 B.n552 585
R1357 B.n554 B.n133 585
R1358 B.n556 B.n555 585
R1359 B.n557 B.n132 585
R1360 B.n559 B.n558 585
R1361 B.n560 B.n131 585
R1362 B.n562 B.n561 585
R1363 B.n563 B.n130 585
R1364 B.n565 B.n564 585
R1365 B.n566 B.n129 585
R1366 B.n568 B.n567 585
R1367 B.n569 B.n128 585
R1368 B.n571 B.n570 585
R1369 B.n572 B.n127 585
R1370 B.n574 B.n573 585
R1371 B.n575 B.n126 585
R1372 B.n577 B.n576 585
R1373 B.n578 B.n125 585
R1374 B.n580 B.n579 585
R1375 B.n581 B.n124 585
R1376 B.n583 B.n582 585
R1377 B.n584 B.n123 585
R1378 B.n586 B.n585 585
R1379 B.n587 B.n122 585
R1380 B.n589 B.n588 585
R1381 B.n590 B.n121 585
R1382 B.n592 B.n591 585
R1383 B.n593 B.n120 585
R1384 B.n595 B.n594 585
R1385 B.n596 B.n119 585
R1386 B.n598 B.n597 585
R1387 B.n599 B.n118 585
R1388 B.n601 B.n600 585
R1389 B.n602 B.n117 585
R1390 B.n604 B.n603 585
R1391 B.n605 B.n116 585
R1392 B.n607 B.n606 585
R1393 B.n608 B.n115 585
R1394 B.n610 B.n609 585
R1395 B.n611 B.n114 585
R1396 B.n613 B.n612 585
R1397 B.n614 B.n113 585
R1398 B.n616 B.n615 585
R1399 B.n617 B.n112 585
R1400 B.n619 B.n618 585
R1401 B.n620 B.n111 585
R1402 B.n622 B.n621 585
R1403 B.n623 B.n110 585
R1404 B.n625 B.n624 585
R1405 B.n626 B.n109 585
R1406 B.n628 B.n627 585
R1407 B.n629 B.n108 585
R1408 B.n631 B.n630 585
R1409 B.n632 B.n107 585
R1410 B.n634 B.n633 585
R1411 B.n635 B.n106 585
R1412 B.n637 B.n636 585
R1413 B.n638 B.n105 585
R1414 B.n640 B.n639 585
R1415 B.n641 B.n104 585
R1416 B.n643 B.n642 585
R1417 B.n644 B.n103 585
R1418 B.n646 B.n645 585
R1419 B.n647 B.n102 585
R1420 B.n649 B.n648 585
R1421 B.n650 B.n101 585
R1422 B.n652 B.n651 585
R1423 B.n653 B.n100 585
R1424 B.n655 B.n654 585
R1425 B.n656 B.n99 585
R1426 B.n658 B.n657 585
R1427 B.n659 B.n98 585
R1428 B.n661 B.n660 585
R1429 B.n662 B.n97 585
R1430 B.n664 B.n663 585
R1431 B.n665 B.n96 585
R1432 B.n667 B.n666 585
R1433 B.n668 B.n95 585
R1434 B.n670 B.n669 585
R1435 B.n671 B.n94 585
R1436 B.n673 B.n672 585
R1437 B.n674 B.n93 585
R1438 B.n676 B.n675 585
R1439 B.n677 B.n92 585
R1440 B.n679 B.n678 585
R1441 B.n680 B.n91 585
R1442 B.n682 B.n681 585
R1443 B.n683 B.n90 585
R1444 B.n685 B.n684 585
R1445 B.n686 B.n89 585
R1446 B.n688 B.n687 585
R1447 B.n689 B.n88 585
R1448 B.n835 B.n834 585
R1449 B.n833 B.n36 585
R1450 B.n832 B.n831 585
R1451 B.n830 B.n37 585
R1452 B.n829 B.n828 585
R1453 B.n827 B.n38 585
R1454 B.n826 B.n825 585
R1455 B.n824 B.n39 585
R1456 B.n823 B.n822 585
R1457 B.n821 B.n40 585
R1458 B.n820 B.n819 585
R1459 B.n818 B.n41 585
R1460 B.n817 B.n816 585
R1461 B.n815 B.n42 585
R1462 B.n814 B.n813 585
R1463 B.n812 B.n43 585
R1464 B.n811 B.n810 585
R1465 B.n809 B.n44 585
R1466 B.n808 B.n807 585
R1467 B.n806 B.n45 585
R1468 B.n805 B.n804 585
R1469 B.n803 B.n46 585
R1470 B.n802 B.n801 585
R1471 B.n800 B.n47 585
R1472 B.n799 B.n798 585
R1473 B.n797 B.n48 585
R1474 B.n796 B.n795 585
R1475 B.n794 B.n49 585
R1476 B.n793 B.n792 585
R1477 B.n791 B.n50 585
R1478 B.n790 B.n789 585
R1479 B.n788 B.n51 585
R1480 B.n787 B.n786 585
R1481 B.n785 B.n52 585
R1482 B.n784 B.n783 585
R1483 B.n782 B.n53 585
R1484 B.n781 B.n780 585
R1485 B.n779 B.n54 585
R1486 B.n778 B.n777 585
R1487 B.n776 B.n55 585
R1488 B.n775 B.n774 585
R1489 B.n773 B.n56 585
R1490 B.n772 B.n771 585
R1491 B.n769 B.n57 585
R1492 B.n768 B.n767 585
R1493 B.n766 B.n60 585
R1494 B.n765 B.n764 585
R1495 B.n763 B.n61 585
R1496 B.n762 B.n761 585
R1497 B.n760 B.n62 585
R1498 B.n759 B.n758 585
R1499 B.n757 B.n63 585
R1500 B.n756 B.n755 585
R1501 B.n754 B.n753 585
R1502 B.n752 B.n67 585
R1503 B.n751 B.n750 585
R1504 B.n749 B.n68 585
R1505 B.n748 B.n747 585
R1506 B.n746 B.n69 585
R1507 B.n745 B.n744 585
R1508 B.n743 B.n70 585
R1509 B.n742 B.n741 585
R1510 B.n740 B.n71 585
R1511 B.n739 B.n738 585
R1512 B.n737 B.n72 585
R1513 B.n736 B.n735 585
R1514 B.n734 B.n73 585
R1515 B.n733 B.n732 585
R1516 B.n731 B.n74 585
R1517 B.n730 B.n729 585
R1518 B.n728 B.n75 585
R1519 B.n727 B.n726 585
R1520 B.n725 B.n76 585
R1521 B.n724 B.n723 585
R1522 B.n722 B.n77 585
R1523 B.n721 B.n720 585
R1524 B.n719 B.n78 585
R1525 B.n718 B.n717 585
R1526 B.n716 B.n79 585
R1527 B.n715 B.n714 585
R1528 B.n713 B.n80 585
R1529 B.n712 B.n711 585
R1530 B.n710 B.n81 585
R1531 B.n709 B.n708 585
R1532 B.n707 B.n82 585
R1533 B.n706 B.n705 585
R1534 B.n704 B.n83 585
R1535 B.n703 B.n702 585
R1536 B.n701 B.n84 585
R1537 B.n700 B.n699 585
R1538 B.n698 B.n85 585
R1539 B.n697 B.n696 585
R1540 B.n695 B.n86 585
R1541 B.n694 B.n693 585
R1542 B.n692 B.n87 585
R1543 B.n691 B.n690 585
R1544 B.n836 B.n35 585
R1545 B.n838 B.n837 585
R1546 B.n839 B.n34 585
R1547 B.n841 B.n840 585
R1548 B.n842 B.n33 585
R1549 B.n844 B.n843 585
R1550 B.n845 B.n32 585
R1551 B.n847 B.n846 585
R1552 B.n848 B.n31 585
R1553 B.n850 B.n849 585
R1554 B.n851 B.n30 585
R1555 B.n853 B.n852 585
R1556 B.n854 B.n29 585
R1557 B.n856 B.n855 585
R1558 B.n857 B.n28 585
R1559 B.n859 B.n858 585
R1560 B.n860 B.n27 585
R1561 B.n862 B.n861 585
R1562 B.n863 B.n26 585
R1563 B.n865 B.n864 585
R1564 B.n866 B.n25 585
R1565 B.n868 B.n867 585
R1566 B.n869 B.n24 585
R1567 B.n871 B.n870 585
R1568 B.n872 B.n23 585
R1569 B.n874 B.n873 585
R1570 B.n875 B.n22 585
R1571 B.n877 B.n876 585
R1572 B.n878 B.n21 585
R1573 B.n880 B.n879 585
R1574 B.n881 B.n20 585
R1575 B.n883 B.n882 585
R1576 B.n884 B.n19 585
R1577 B.n886 B.n885 585
R1578 B.n887 B.n18 585
R1579 B.n889 B.n888 585
R1580 B.n890 B.n17 585
R1581 B.n892 B.n891 585
R1582 B.n893 B.n16 585
R1583 B.n895 B.n894 585
R1584 B.n896 B.n15 585
R1585 B.n898 B.n897 585
R1586 B.n899 B.n14 585
R1587 B.n901 B.n900 585
R1588 B.n902 B.n13 585
R1589 B.n904 B.n903 585
R1590 B.n905 B.n12 585
R1591 B.n907 B.n906 585
R1592 B.n908 B.n11 585
R1593 B.n910 B.n909 585
R1594 B.n911 B.n10 585
R1595 B.n913 B.n912 585
R1596 B.n914 B.n9 585
R1597 B.n916 B.n915 585
R1598 B.n917 B.n8 585
R1599 B.n919 B.n918 585
R1600 B.n920 B.n7 585
R1601 B.n922 B.n921 585
R1602 B.n923 B.n6 585
R1603 B.n925 B.n924 585
R1604 B.n926 B.n5 585
R1605 B.n928 B.n927 585
R1606 B.n929 B.n4 585
R1607 B.n931 B.n930 585
R1608 B.n932 B.n3 585
R1609 B.n934 B.n933 585
R1610 B.n935 B.n0 585
R1611 B.n2 B.n1 585
R1612 B.n240 B.n239 585
R1613 B.n241 B.n238 585
R1614 B.n243 B.n242 585
R1615 B.n244 B.n237 585
R1616 B.n246 B.n245 585
R1617 B.n247 B.n236 585
R1618 B.n249 B.n248 585
R1619 B.n250 B.n235 585
R1620 B.n252 B.n251 585
R1621 B.n253 B.n234 585
R1622 B.n255 B.n254 585
R1623 B.n256 B.n233 585
R1624 B.n258 B.n257 585
R1625 B.n259 B.n232 585
R1626 B.n261 B.n260 585
R1627 B.n262 B.n231 585
R1628 B.n264 B.n263 585
R1629 B.n265 B.n230 585
R1630 B.n267 B.n266 585
R1631 B.n268 B.n229 585
R1632 B.n270 B.n269 585
R1633 B.n271 B.n228 585
R1634 B.n273 B.n272 585
R1635 B.n274 B.n227 585
R1636 B.n276 B.n275 585
R1637 B.n277 B.n226 585
R1638 B.n279 B.n278 585
R1639 B.n280 B.n225 585
R1640 B.n282 B.n281 585
R1641 B.n283 B.n224 585
R1642 B.n285 B.n284 585
R1643 B.n286 B.n223 585
R1644 B.n288 B.n287 585
R1645 B.n289 B.n222 585
R1646 B.n291 B.n290 585
R1647 B.n292 B.n221 585
R1648 B.n294 B.n293 585
R1649 B.n295 B.n220 585
R1650 B.n297 B.n296 585
R1651 B.n298 B.n219 585
R1652 B.n300 B.n299 585
R1653 B.n301 B.n218 585
R1654 B.n303 B.n302 585
R1655 B.n304 B.n217 585
R1656 B.n306 B.n305 585
R1657 B.n307 B.n216 585
R1658 B.n309 B.n308 585
R1659 B.n310 B.n215 585
R1660 B.n312 B.n311 585
R1661 B.n313 B.n214 585
R1662 B.n315 B.n314 585
R1663 B.n316 B.n213 585
R1664 B.n318 B.n317 585
R1665 B.n319 B.n212 585
R1666 B.n321 B.n320 585
R1667 B.n322 B.n211 585
R1668 B.n324 B.n323 585
R1669 B.n325 B.n210 585
R1670 B.n327 B.n326 585
R1671 B.n328 B.n209 585
R1672 B.n330 B.n329 585
R1673 B.n331 B.n208 585
R1674 B.n333 B.n332 585
R1675 B.n334 B.n207 585
R1676 B.n336 B.n335 585
R1677 B.n337 B.n206 585
R1678 B.n338 B.n337 530.939
R1679 B.n486 B.n485 530.939
R1680 B.n690 B.n689 530.939
R1681 B.n834 B.n35 530.939
R1682 B.n178 B.t1 451.195
R1683 B.n64 B.t5 451.195
R1684 B.n401 B.t7 451.195
R1685 B.n58 B.t11 451.195
R1686 B.n179 B.t2 385.837
R1687 B.n65 B.t4 385.837
R1688 B.n402 B.t8 385.837
R1689 B.n59 B.t10 385.837
R1690 B.n401 B.t6 308.356
R1691 B.n178 B.t0 308.356
R1692 B.n64 B.t3 308.356
R1693 B.n58 B.t9 308.356
R1694 B.n937 B.n936 256.663
R1695 B.n936 B.n935 235.042
R1696 B.n936 B.n2 235.042
R1697 B.n338 B.n205 163.367
R1698 B.n342 B.n205 163.367
R1699 B.n343 B.n342 163.367
R1700 B.n344 B.n343 163.367
R1701 B.n344 B.n203 163.367
R1702 B.n348 B.n203 163.367
R1703 B.n349 B.n348 163.367
R1704 B.n350 B.n349 163.367
R1705 B.n350 B.n201 163.367
R1706 B.n354 B.n201 163.367
R1707 B.n355 B.n354 163.367
R1708 B.n356 B.n355 163.367
R1709 B.n356 B.n199 163.367
R1710 B.n360 B.n199 163.367
R1711 B.n361 B.n360 163.367
R1712 B.n362 B.n361 163.367
R1713 B.n362 B.n197 163.367
R1714 B.n366 B.n197 163.367
R1715 B.n367 B.n366 163.367
R1716 B.n368 B.n367 163.367
R1717 B.n368 B.n195 163.367
R1718 B.n372 B.n195 163.367
R1719 B.n373 B.n372 163.367
R1720 B.n374 B.n373 163.367
R1721 B.n374 B.n193 163.367
R1722 B.n378 B.n193 163.367
R1723 B.n379 B.n378 163.367
R1724 B.n380 B.n379 163.367
R1725 B.n380 B.n191 163.367
R1726 B.n384 B.n191 163.367
R1727 B.n385 B.n384 163.367
R1728 B.n386 B.n385 163.367
R1729 B.n386 B.n189 163.367
R1730 B.n390 B.n189 163.367
R1731 B.n391 B.n390 163.367
R1732 B.n392 B.n391 163.367
R1733 B.n392 B.n187 163.367
R1734 B.n396 B.n187 163.367
R1735 B.n397 B.n396 163.367
R1736 B.n398 B.n397 163.367
R1737 B.n398 B.n185 163.367
R1738 B.n405 B.n185 163.367
R1739 B.n406 B.n405 163.367
R1740 B.n407 B.n406 163.367
R1741 B.n407 B.n183 163.367
R1742 B.n411 B.n183 163.367
R1743 B.n412 B.n411 163.367
R1744 B.n413 B.n412 163.367
R1745 B.n413 B.n181 163.367
R1746 B.n417 B.n181 163.367
R1747 B.n418 B.n417 163.367
R1748 B.n419 B.n418 163.367
R1749 B.n419 B.n177 163.367
R1750 B.n424 B.n177 163.367
R1751 B.n425 B.n424 163.367
R1752 B.n426 B.n425 163.367
R1753 B.n426 B.n175 163.367
R1754 B.n430 B.n175 163.367
R1755 B.n431 B.n430 163.367
R1756 B.n432 B.n431 163.367
R1757 B.n432 B.n173 163.367
R1758 B.n436 B.n173 163.367
R1759 B.n437 B.n436 163.367
R1760 B.n438 B.n437 163.367
R1761 B.n438 B.n171 163.367
R1762 B.n442 B.n171 163.367
R1763 B.n443 B.n442 163.367
R1764 B.n444 B.n443 163.367
R1765 B.n444 B.n169 163.367
R1766 B.n448 B.n169 163.367
R1767 B.n449 B.n448 163.367
R1768 B.n450 B.n449 163.367
R1769 B.n450 B.n167 163.367
R1770 B.n454 B.n167 163.367
R1771 B.n455 B.n454 163.367
R1772 B.n456 B.n455 163.367
R1773 B.n456 B.n165 163.367
R1774 B.n460 B.n165 163.367
R1775 B.n461 B.n460 163.367
R1776 B.n462 B.n461 163.367
R1777 B.n462 B.n163 163.367
R1778 B.n466 B.n163 163.367
R1779 B.n467 B.n466 163.367
R1780 B.n468 B.n467 163.367
R1781 B.n468 B.n161 163.367
R1782 B.n472 B.n161 163.367
R1783 B.n473 B.n472 163.367
R1784 B.n474 B.n473 163.367
R1785 B.n474 B.n159 163.367
R1786 B.n478 B.n159 163.367
R1787 B.n479 B.n478 163.367
R1788 B.n480 B.n479 163.367
R1789 B.n480 B.n157 163.367
R1790 B.n484 B.n157 163.367
R1791 B.n485 B.n484 163.367
R1792 B.n689 B.n688 163.367
R1793 B.n688 B.n89 163.367
R1794 B.n684 B.n89 163.367
R1795 B.n684 B.n683 163.367
R1796 B.n683 B.n682 163.367
R1797 B.n682 B.n91 163.367
R1798 B.n678 B.n91 163.367
R1799 B.n678 B.n677 163.367
R1800 B.n677 B.n676 163.367
R1801 B.n676 B.n93 163.367
R1802 B.n672 B.n93 163.367
R1803 B.n672 B.n671 163.367
R1804 B.n671 B.n670 163.367
R1805 B.n670 B.n95 163.367
R1806 B.n666 B.n95 163.367
R1807 B.n666 B.n665 163.367
R1808 B.n665 B.n664 163.367
R1809 B.n664 B.n97 163.367
R1810 B.n660 B.n97 163.367
R1811 B.n660 B.n659 163.367
R1812 B.n659 B.n658 163.367
R1813 B.n658 B.n99 163.367
R1814 B.n654 B.n99 163.367
R1815 B.n654 B.n653 163.367
R1816 B.n653 B.n652 163.367
R1817 B.n652 B.n101 163.367
R1818 B.n648 B.n101 163.367
R1819 B.n648 B.n647 163.367
R1820 B.n647 B.n646 163.367
R1821 B.n646 B.n103 163.367
R1822 B.n642 B.n103 163.367
R1823 B.n642 B.n641 163.367
R1824 B.n641 B.n640 163.367
R1825 B.n640 B.n105 163.367
R1826 B.n636 B.n105 163.367
R1827 B.n636 B.n635 163.367
R1828 B.n635 B.n634 163.367
R1829 B.n634 B.n107 163.367
R1830 B.n630 B.n107 163.367
R1831 B.n630 B.n629 163.367
R1832 B.n629 B.n628 163.367
R1833 B.n628 B.n109 163.367
R1834 B.n624 B.n109 163.367
R1835 B.n624 B.n623 163.367
R1836 B.n623 B.n622 163.367
R1837 B.n622 B.n111 163.367
R1838 B.n618 B.n111 163.367
R1839 B.n618 B.n617 163.367
R1840 B.n617 B.n616 163.367
R1841 B.n616 B.n113 163.367
R1842 B.n612 B.n113 163.367
R1843 B.n612 B.n611 163.367
R1844 B.n611 B.n610 163.367
R1845 B.n610 B.n115 163.367
R1846 B.n606 B.n115 163.367
R1847 B.n606 B.n605 163.367
R1848 B.n605 B.n604 163.367
R1849 B.n604 B.n117 163.367
R1850 B.n600 B.n117 163.367
R1851 B.n600 B.n599 163.367
R1852 B.n599 B.n598 163.367
R1853 B.n598 B.n119 163.367
R1854 B.n594 B.n119 163.367
R1855 B.n594 B.n593 163.367
R1856 B.n593 B.n592 163.367
R1857 B.n592 B.n121 163.367
R1858 B.n588 B.n121 163.367
R1859 B.n588 B.n587 163.367
R1860 B.n587 B.n586 163.367
R1861 B.n586 B.n123 163.367
R1862 B.n582 B.n123 163.367
R1863 B.n582 B.n581 163.367
R1864 B.n581 B.n580 163.367
R1865 B.n580 B.n125 163.367
R1866 B.n576 B.n125 163.367
R1867 B.n576 B.n575 163.367
R1868 B.n575 B.n574 163.367
R1869 B.n574 B.n127 163.367
R1870 B.n570 B.n127 163.367
R1871 B.n570 B.n569 163.367
R1872 B.n569 B.n568 163.367
R1873 B.n568 B.n129 163.367
R1874 B.n564 B.n129 163.367
R1875 B.n564 B.n563 163.367
R1876 B.n563 B.n562 163.367
R1877 B.n562 B.n131 163.367
R1878 B.n558 B.n131 163.367
R1879 B.n558 B.n557 163.367
R1880 B.n557 B.n556 163.367
R1881 B.n556 B.n133 163.367
R1882 B.n552 B.n133 163.367
R1883 B.n552 B.n551 163.367
R1884 B.n551 B.n550 163.367
R1885 B.n550 B.n135 163.367
R1886 B.n546 B.n135 163.367
R1887 B.n546 B.n545 163.367
R1888 B.n545 B.n544 163.367
R1889 B.n544 B.n137 163.367
R1890 B.n540 B.n137 163.367
R1891 B.n540 B.n539 163.367
R1892 B.n539 B.n538 163.367
R1893 B.n538 B.n139 163.367
R1894 B.n534 B.n139 163.367
R1895 B.n534 B.n533 163.367
R1896 B.n533 B.n532 163.367
R1897 B.n532 B.n141 163.367
R1898 B.n528 B.n141 163.367
R1899 B.n528 B.n527 163.367
R1900 B.n527 B.n526 163.367
R1901 B.n526 B.n143 163.367
R1902 B.n522 B.n143 163.367
R1903 B.n522 B.n521 163.367
R1904 B.n521 B.n520 163.367
R1905 B.n520 B.n145 163.367
R1906 B.n516 B.n145 163.367
R1907 B.n516 B.n515 163.367
R1908 B.n515 B.n514 163.367
R1909 B.n514 B.n147 163.367
R1910 B.n510 B.n147 163.367
R1911 B.n510 B.n509 163.367
R1912 B.n509 B.n508 163.367
R1913 B.n508 B.n149 163.367
R1914 B.n504 B.n149 163.367
R1915 B.n504 B.n503 163.367
R1916 B.n503 B.n502 163.367
R1917 B.n502 B.n151 163.367
R1918 B.n498 B.n151 163.367
R1919 B.n498 B.n497 163.367
R1920 B.n497 B.n496 163.367
R1921 B.n496 B.n153 163.367
R1922 B.n492 B.n153 163.367
R1923 B.n492 B.n491 163.367
R1924 B.n491 B.n490 163.367
R1925 B.n490 B.n155 163.367
R1926 B.n486 B.n155 163.367
R1927 B.n834 B.n833 163.367
R1928 B.n833 B.n832 163.367
R1929 B.n832 B.n37 163.367
R1930 B.n828 B.n37 163.367
R1931 B.n828 B.n827 163.367
R1932 B.n827 B.n826 163.367
R1933 B.n826 B.n39 163.367
R1934 B.n822 B.n39 163.367
R1935 B.n822 B.n821 163.367
R1936 B.n821 B.n820 163.367
R1937 B.n820 B.n41 163.367
R1938 B.n816 B.n41 163.367
R1939 B.n816 B.n815 163.367
R1940 B.n815 B.n814 163.367
R1941 B.n814 B.n43 163.367
R1942 B.n810 B.n43 163.367
R1943 B.n810 B.n809 163.367
R1944 B.n809 B.n808 163.367
R1945 B.n808 B.n45 163.367
R1946 B.n804 B.n45 163.367
R1947 B.n804 B.n803 163.367
R1948 B.n803 B.n802 163.367
R1949 B.n802 B.n47 163.367
R1950 B.n798 B.n47 163.367
R1951 B.n798 B.n797 163.367
R1952 B.n797 B.n796 163.367
R1953 B.n796 B.n49 163.367
R1954 B.n792 B.n49 163.367
R1955 B.n792 B.n791 163.367
R1956 B.n791 B.n790 163.367
R1957 B.n790 B.n51 163.367
R1958 B.n786 B.n51 163.367
R1959 B.n786 B.n785 163.367
R1960 B.n785 B.n784 163.367
R1961 B.n784 B.n53 163.367
R1962 B.n780 B.n53 163.367
R1963 B.n780 B.n779 163.367
R1964 B.n779 B.n778 163.367
R1965 B.n778 B.n55 163.367
R1966 B.n774 B.n55 163.367
R1967 B.n774 B.n773 163.367
R1968 B.n773 B.n772 163.367
R1969 B.n772 B.n57 163.367
R1970 B.n767 B.n57 163.367
R1971 B.n767 B.n766 163.367
R1972 B.n766 B.n765 163.367
R1973 B.n765 B.n61 163.367
R1974 B.n761 B.n61 163.367
R1975 B.n761 B.n760 163.367
R1976 B.n760 B.n759 163.367
R1977 B.n759 B.n63 163.367
R1978 B.n755 B.n63 163.367
R1979 B.n755 B.n754 163.367
R1980 B.n754 B.n67 163.367
R1981 B.n750 B.n67 163.367
R1982 B.n750 B.n749 163.367
R1983 B.n749 B.n748 163.367
R1984 B.n748 B.n69 163.367
R1985 B.n744 B.n69 163.367
R1986 B.n744 B.n743 163.367
R1987 B.n743 B.n742 163.367
R1988 B.n742 B.n71 163.367
R1989 B.n738 B.n71 163.367
R1990 B.n738 B.n737 163.367
R1991 B.n737 B.n736 163.367
R1992 B.n736 B.n73 163.367
R1993 B.n732 B.n73 163.367
R1994 B.n732 B.n731 163.367
R1995 B.n731 B.n730 163.367
R1996 B.n730 B.n75 163.367
R1997 B.n726 B.n75 163.367
R1998 B.n726 B.n725 163.367
R1999 B.n725 B.n724 163.367
R2000 B.n724 B.n77 163.367
R2001 B.n720 B.n77 163.367
R2002 B.n720 B.n719 163.367
R2003 B.n719 B.n718 163.367
R2004 B.n718 B.n79 163.367
R2005 B.n714 B.n79 163.367
R2006 B.n714 B.n713 163.367
R2007 B.n713 B.n712 163.367
R2008 B.n712 B.n81 163.367
R2009 B.n708 B.n81 163.367
R2010 B.n708 B.n707 163.367
R2011 B.n707 B.n706 163.367
R2012 B.n706 B.n83 163.367
R2013 B.n702 B.n83 163.367
R2014 B.n702 B.n701 163.367
R2015 B.n701 B.n700 163.367
R2016 B.n700 B.n85 163.367
R2017 B.n696 B.n85 163.367
R2018 B.n696 B.n695 163.367
R2019 B.n695 B.n694 163.367
R2020 B.n694 B.n87 163.367
R2021 B.n690 B.n87 163.367
R2022 B.n838 B.n35 163.367
R2023 B.n839 B.n838 163.367
R2024 B.n840 B.n839 163.367
R2025 B.n840 B.n33 163.367
R2026 B.n844 B.n33 163.367
R2027 B.n845 B.n844 163.367
R2028 B.n846 B.n845 163.367
R2029 B.n846 B.n31 163.367
R2030 B.n850 B.n31 163.367
R2031 B.n851 B.n850 163.367
R2032 B.n852 B.n851 163.367
R2033 B.n852 B.n29 163.367
R2034 B.n856 B.n29 163.367
R2035 B.n857 B.n856 163.367
R2036 B.n858 B.n857 163.367
R2037 B.n858 B.n27 163.367
R2038 B.n862 B.n27 163.367
R2039 B.n863 B.n862 163.367
R2040 B.n864 B.n863 163.367
R2041 B.n864 B.n25 163.367
R2042 B.n868 B.n25 163.367
R2043 B.n869 B.n868 163.367
R2044 B.n870 B.n869 163.367
R2045 B.n870 B.n23 163.367
R2046 B.n874 B.n23 163.367
R2047 B.n875 B.n874 163.367
R2048 B.n876 B.n875 163.367
R2049 B.n876 B.n21 163.367
R2050 B.n880 B.n21 163.367
R2051 B.n881 B.n880 163.367
R2052 B.n882 B.n881 163.367
R2053 B.n882 B.n19 163.367
R2054 B.n886 B.n19 163.367
R2055 B.n887 B.n886 163.367
R2056 B.n888 B.n887 163.367
R2057 B.n888 B.n17 163.367
R2058 B.n892 B.n17 163.367
R2059 B.n893 B.n892 163.367
R2060 B.n894 B.n893 163.367
R2061 B.n894 B.n15 163.367
R2062 B.n898 B.n15 163.367
R2063 B.n899 B.n898 163.367
R2064 B.n900 B.n899 163.367
R2065 B.n900 B.n13 163.367
R2066 B.n904 B.n13 163.367
R2067 B.n905 B.n904 163.367
R2068 B.n906 B.n905 163.367
R2069 B.n906 B.n11 163.367
R2070 B.n910 B.n11 163.367
R2071 B.n911 B.n910 163.367
R2072 B.n912 B.n911 163.367
R2073 B.n912 B.n9 163.367
R2074 B.n916 B.n9 163.367
R2075 B.n917 B.n916 163.367
R2076 B.n918 B.n917 163.367
R2077 B.n918 B.n7 163.367
R2078 B.n922 B.n7 163.367
R2079 B.n923 B.n922 163.367
R2080 B.n924 B.n923 163.367
R2081 B.n924 B.n5 163.367
R2082 B.n928 B.n5 163.367
R2083 B.n929 B.n928 163.367
R2084 B.n930 B.n929 163.367
R2085 B.n930 B.n3 163.367
R2086 B.n934 B.n3 163.367
R2087 B.n935 B.n934 163.367
R2088 B.n240 B.n2 163.367
R2089 B.n241 B.n240 163.367
R2090 B.n242 B.n241 163.367
R2091 B.n242 B.n237 163.367
R2092 B.n246 B.n237 163.367
R2093 B.n247 B.n246 163.367
R2094 B.n248 B.n247 163.367
R2095 B.n248 B.n235 163.367
R2096 B.n252 B.n235 163.367
R2097 B.n253 B.n252 163.367
R2098 B.n254 B.n253 163.367
R2099 B.n254 B.n233 163.367
R2100 B.n258 B.n233 163.367
R2101 B.n259 B.n258 163.367
R2102 B.n260 B.n259 163.367
R2103 B.n260 B.n231 163.367
R2104 B.n264 B.n231 163.367
R2105 B.n265 B.n264 163.367
R2106 B.n266 B.n265 163.367
R2107 B.n266 B.n229 163.367
R2108 B.n270 B.n229 163.367
R2109 B.n271 B.n270 163.367
R2110 B.n272 B.n271 163.367
R2111 B.n272 B.n227 163.367
R2112 B.n276 B.n227 163.367
R2113 B.n277 B.n276 163.367
R2114 B.n278 B.n277 163.367
R2115 B.n278 B.n225 163.367
R2116 B.n282 B.n225 163.367
R2117 B.n283 B.n282 163.367
R2118 B.n284 B.n283 163.367
R2119 B.n284 B.n223 163.367
R2120 B.n288 B.n223 163.367
R2121 B.n289 B.n288 163.367
R2122 B.n290 B.n289 163.367
R2123 B.n290 B.n221 163.367
R2124 B.n294 B.n221 163.367
R2125 B.n295 B.n294 163.367
R2126 B.n296 B.n295 163.367
R2127 B.n296 B.n219 163.367
R2128 B.n300 B.n219 163.367
R2129 B.n301 B.n300 163.367
R2130 B.n302 B.n301 163.367
R2131 B.n302 B.n217 163.367
R2132 B.n306 B.n217 163.367
R2133 B.n307 B.n306 163.367
R2134 B.n308 B.n307 163.367
R2135 B.n308 B.n215 163.367
R2136 B.n312 B.n215 163.367
R2137 B.n313 B.n312 163.367
R2138 B.n314 B.n313 163.367
R2139 B.n314 B.n213 163.367
R2140 B.n318 B.n213 163.367
R2141 B.n319 B.n318 163.367
R2142 B.n320 B.n319 163.367
R2143 B.n320 B.n211 163.367
R2144 B.n324 B.n211 163.367
R2145 B.n325 B.n324 163.367
R2146 B.n326 B.n325 163.367
R2147 B.n326 B.n209 163.367
R2148 B.n330 B.n209 163.367
R2149 B.n331 B.n330 163.367
R2150 B.n332 B.n331 163.367
R2151 B.n332 B.n207 163.367
R2152 B.n336 B.n207 163.367
R2153 B.n337 B.n336 163.367
R2154 B.n402 B.n401 65.3581
R2155 B.n179 B.n178 65.3581
R2156 B.n65 B.n64 65.3581
R2157 B.n59 B.n58 65.3581
R2158 B.n403 B.n402 59.5399
R2159 B.n421 B.n179 59.5399
R2160 B.n66 B.n65 59.5399
R2161 B.n770 B.n59 59.5399
R2162 B.n836 B.n835 34.4981
R2163 B.n691 B.n88 34.4981
R2164 B.n487 B.n156 34.4981
R2165 B.n339 B.n206 34.4981
R2166 B B.n937 18.0485
R2167 B.n837 B.n836 10.6151
R2168 B.n837 B.n34 10.6151
R2169 B.n841 B.n34 10.6151
R2170 B.n842 B.n841 10.6151
R2171 B.n843 B.n842 10.6151
R2172 B.n843 B.n32 10.6151
R2173 B.n847 B.n32 10.6151
R2174 B.n848 B.n847 10.6151
R2175 B.n849 B.n848 10.6151
R2176 B.n849 B.n30 10.6151
R2177 B.n853 B.n30 10.6151
R2178 B.n854 B.n853 10.6151
R2179 B.n855 B.n854 10.6151
R2180 B.n855 B.n28 10.6151
R2181 B.n859 B.n28 10.6151
R2182 B.n860 B.n859 10.6151
R2183 B.n861 B.n860 10.6151
R2184 B.n861 B.n26 10.6151
R2185 B.n865 B.n26 10.6151
R2186 B.n866 B.n865 10.6151
R2187 B.n867 B.n866 10.6151
R2188 B.n867 B.n24 10.6151
R2189 B.n871 B.n24 10.6151
R2190 B.n872 B.n871 10.6151
R2191 B.n873 B.n872 10.6151
R2192 B.n873 B.n22 10.6151
R2193 B.n877 B.n22 10.6151
R2194 B.n878 B.n877 10.6151
R2195 B.n879 B.n878 10.6151
R2196 B.n879 B.n20 10.6151
R2197 B.n883 B.n20 10.6151
R2198 B.n884 B.n883 10.6151
R2199 B.n885 B.n884 10.6151
R2200 B.n885 B.n18 10.6151
R2201 B.n889 B.n18 10.6151
R2202 B.n890 B.n889 10.6151
R2203 B.n891 B.n890 10.6151
R2204 B.n891 B.n16 10.6151
R2205 B.n895 B.n16 10.6151
R2206 B.n896 B.n895 10.6151
R2207 B.n897 B.n896 10.6151
R2208 B.n897 B.n14 10.6151
R2209 B.n901 B.n14 10.6151
R2210 B.n902 B.n901 10.6151
R2211 B.n903 B.n902 10.6151
R2212 B.n903 B.n12 10.6151
R2213 B.n907 B.n12 10.6151
R2214 B.n908 B.n907 10.6151
R2215 B.n909 B.n908 10.6151
R2216 B.n909 B.n10 10.6151
R2217 B.n913 B.n10 10.6151
R2218 B.n914 B.n913 10.6151
R2219 B.n915 B.n914 10.6151
R2220 B.n915 B.n8 10.6151
R2221 B.n919 B.n8 10.6151
R2222 B.n920 B.n919 10.6151
R2223 B.n921 B.n920 10.6151
R2224 B.n921 B.n6 10.6151
R2225 B.n925 B.n6 10.6151
R2226 B.n926 B.n925 10.6151
R2227 B.n927 B.n926 10.6151
R2228 B.n927 B.n4 10.6151
R2229 B.n931 B.n4 10.6151
R2230 B.n932 B.n931 10.6151
R2231 B.n933 B.n932 10.6151
R2232 B.n933 B.n0 10.6151
R2233 B.n835 B.n36 10.6151
R2234 B.n831 B.n36 10.6151
R2235 B.n831 B.n830 10.6151
R2236 B.n830 B.n829 10.6151
R2237 B.n829 B.n38 10.6151
R2238 B.n825 B.n38 10.6151
R2239 B.n825 B.n824 10.6151
R2240 B.n824 B.n823 10.6151
R2241 B.n823 B.n40 10.6151
R2242 B.n819 B.n40 10.6151
R2243 B.n819 B.n818 10.6151
R2244 B.n818 B.n817 10.6151
R2245 B.n817 B.n42 10.6151
R2246 B.n813 B.n42 10.6151
R2247 B.n813 B.n812 10.6151
R2248 B.n812 B.n811 10.6151
R2249 B.n811 B.n44 10.6151
R2250 B.n807 B.n44 10.6151
R2251 B.n807 B.n806 10.6151
R2252 B.n806 B.n805 10.6151
R2253 B.n805 B.n46 10.6151
R2254 B.n801 B.n46 10.6151
R2255 B.n801 B.n800 10.6151
R2256 B.n800 B.n799 10.6151
R2257 B.n799 B.n48 10.6151
R2258 B.n795 B.n48 10.6151
R2259 B.n795 B.n794 10.6151
R2260 B.n794 B.n793 10.6151
R2261 B.n793 B.n50 10.6151
R2262 B.n789 B.n50 10.6151
R2263 B.n789 B.n788 10.6151
R2264 B.n788 B.n787 10.6151
R2265 B.n787 B.n52 10.6151
R2266 B.n783 B.n52 10.6151
R2267 B.n783 B.n782 10.6151
R2268 B.n782 B.n781 10.6151
R2269 B.n781 B.n54 10.6151
R2270 B.n777 B.n54 10.6151
R2271 B.n777 B.n776 10.6151
R2272 B.n776 B.n775 10.6151
R2273 B.n775 B.n56 10.6151
R2274 B.n771 B.n56 10.6151
R2275 B.n769 B.n768 10.6151
R2276 B.n768 B.n60 10.6151
R2277 B.n764 B.n60 10.6151
R2278 B.n764 B.n763 10.6151
R2279 B.n763 B.n762 10.6151
R2280 B.n762 B.n62 10.6151
R2281 B.n758 B.n62 10.6151
R2282 B.n758 B.n757 10.6151
R2283 B.n757 B.n756 10.6151
R2284 B.n753 B.n752 10.6151
R2285 B.n752 B.n751 10.6151
R2286 B.n751 B.n68 10.6151
R2287 B.n747 B.n68 10.6151
R2288 B.n747 B.n746 10.6151
R2289 B.n746 B.n745 10.6151
R2290 B.n745 B.n70 10.6151
R2291 B.n741 B.n70 10.6151
R2292 B.n741 B.n740 10.6151
R2293 B.n740 B.n739 10.6151
R2294 B.n739 B.n72 10.6151
R2295 B.n735 B.n72 10.6151
R2296 B.n735 B.n734 10.6151
R2297 B.n734 B.n733 10.6151
R2298 B.n733 B.n74 10.6151
R2299 B.n729 B.n74 10.6151
R2300 B.n729 B.n728 10.6151
R2301 B.n728 B.n727 10.6151
R2302 B.n727 B.n76 10.6151
R2303 B.n723 B.n76 10.6151
R2304 B.n723 B.n722 10.6151
R2305 B.n722 B.n721 10.6151
R2306 B.n721 B.n78 10.6151
R2307 B.n717 B.n78 10.6151
R2308 B.n717 B.n716 10.6151
R2309 B.n716 B.n715 10.6151
R2310 B.n715 B.n80 10.6151
R2311 B.n711 B.n80 10.6151
R2312 B.n711 B.n710 10.6151
R2313 B.n710 B.n709 10.6151
R2314 B.n709 B.n82 10.6151
R2315 B.n705 B.n82 10.6151
R2316 B.n705 B.n704 10.6151
R2317 B.n704 B.n703 10.6151
R2318 B.n703 B.n84 10.6151
R2319 B.n699 B.n84 10.6151
R2320 B.n699 B.n698 10.6151
R2321 B.n698 B.n697 10.6151
R2322 B.n697 B.n86 10.6151
R2323 B.n693 B.n86 10.6151
R2324 B.n693 B.n692 10.6151
R2325 B.n692 B.n691 10.6151
R2326 B.n687 B.n88 10.6151
R2327 B.n687 B.n686 10.6151
R2328 B.n686 B.n685 10.6151
R2329 B.n685 B.n90 10.6151
R2330 B.n681 B.n90 10.6151
R2331 B.n681 B.n680 10.6151
R2332 B.n680 B.n679 10.6151
R2333 B.n679 B.n92 10.6151
R2334 B.n675 B.n92 10.6151
R2335 B.n675 B.n674 10.6151
R2336 B.n674 B.n673 10.6151
R2337 B.n673 B.n94 10.6151
R2338 B.n669 B.n94 10.6151
R2339 B.n669 B.n668 10.6151
R2340 B.n668 B.n667 10.6151
R2341 B.n667 B.n96 10.6151
R2342 B.n663 B.n96 10.6151
R2343 B.n663 B.n662 10.6151
R2344 B.n662 B.n661 10.6151
R2345 B.n661 B.n98 10.6151
R2346 B.n657 B.n98 10.6151
R2347 B.n657 B.n656 10.6151
R2348 B.n656 B.n655 10.6151
R2349 B.n655 B.n100 10.6151
R2350 B.n651 B.n100 10.6151
R2351 B.n651 B.n650 10.6151
R2352 B.n650 B.n649 10.6151
R2353 B.n649 B.n102 10.6151
R2354 B.n645 B.n102 10.6151
R2355 B.n645 B.n644 10.6151
R2356 B.n644 B.n643 10.6151
R2357 B.n643 B.n104 10.6151
R2358 B.n639 B.n104 10.6151
R2359 B.n639 B.n638 10.6151
R2360 B.n638 B.n637 10.6151
R2361 B.n637 B.n106 10.6151
R2362 B.n633 B.n106 10.6151
R2363 B.n633 B.n632 10.6151
R2364 B.n632 B.n631 10.6151
R2365 B.n631 B.n108 10.6151
R2366 B.n627 B.n108 10.6151
R2367 B.n627 B.n626 10.6151
R2368 B.n626 B.n625 10.6151
R2369 B.n625 B.n110 10.6151
R2370 B.n621 B.n110 10.6151
R2371 B.n621 B.n620 10.6151
R2372 B.n620 B.n619 10.6151
R2373 B.n619 B.n112 10.6151
R2374 B.n615 B.n112 10.6151
R2375 B.n615 B.n614 10.6151
R2376 B.n614 B.n613 10.6151
R2377 B.n613 B.n114 10.6151
R2378 B.n609 B.n114 10.6151
R2379 B.n609 B.n608 10.6151
R2380 B.n608 B.n607 10.6151
R2381 B.n607 B.n116 10.6151
R2382 B.n603 B.n116 10.6151
R2383 B.n603 B.n602 10.6151
R2384 B.n602 B.n601 10.6151
R2385 B.n601 B.n118 10.6151
R2386 B.n597 B.n118 10.6151
R2387 B.n597 B.n596 10.6151
R2388 B.n596 B.n595 10.6151
R2389 B.n595 B.n120 10.6151
R2390 B.n591 B.n120 10.6151
R2391 B.n591 B.n590 10.6151
R2392 B.n590 B.n589 10.6151
R2393 B.n589 B.n122 10.6151
R2394 B.n585 B.n122 10.6151
R2395 B.n585 B.n584 10.6151
R2396 B.n584 B.n583 10.6151
R2397 B.n583 B.n124 10.6151
R2398 B.n579 B.n124 10.6151
R2399 B.n579 B.n578 10.6151
R2400 B.n578 B.n577 10.6151
R2401 B.n577 B.n126 10.6151
R2402 B.n573 B.n126 10.6151
R2403 B.n573 B.n572 10.6151
R2404 B.n572 B.n571 10.6151
R2405 B.n571 B.n128 10.6151
R2406 B.n567 B.n128 10.6151
R2407 B.n567 B.n566 10.6151
R2408 B.n566 B.n565 10.6151
R2409 B.n565 B.n130 10.6151
R2410 B.n561 B.n130 10.6151
R2411 B.n561 B.n560 10.6151
R2412 B.n560 B.n559 10.6151
R2413 B.n559 B.n132 10.6151
R2414 B.n555 B.n132 10.6151
R2415 B.n555 B.n554 10.6151
R2416 B.n554 B.n553 10.6151
R2417 B.n553 B.n134 10.6151
R2418 B.n549 B.n134 10.6151
R2419 B.n549 B.n548 10.6151
R2420 B.n548 B.n547 10.6151
R2421 B.n547 B.n136 10.6151
R2422 B.n543 B.n136 10.6151
R2423 B.n543 B.n542 10.6151
R2424 B.n542 B.n541 10.6151
R2425 B.n541 B.n138 10.6151
R2426 B.n537 B.n138 10.6151
R2427 B.n537 B.n536 10.6151
R2428 B.n536 B.n535 10.6151
R2429 B.n535 B.n140 10.6151
R2430 B.n531 B.n140 10.6151
R2431 B.n531 B.n530 10.6151
R2432 B.n530 B.n529 10.6151
R2433 B.n529 B.n142 10.6151
R2434 B.n525 B.n142 10.6151
R2435 B.n525 B.n524 10.6151
R2436 B.n524 B.n523 10.6151
R2437 B.n523 B.n144 10.6151
R2438 B.n519 B.n144 10.6151
R2439 B.n519 B.n518 10.6151
R2440 B.n518 B.n517 10.6151
R2441 B.n517 B.n146 10.6151
R2442 B.n513 B.n146 10.6151
R2443 B.n513 B.n512 10.6151
R2444 B.n512 B.n511 10.6151
R2445 B.n511 B.n148 10.6151
R2446 B.n507 B.n148 10.6151
R2447 B.n507 B.n506 10.6151
R2448 B.n506 B.n505 10.6151
R2449 B.n505 B.n150 10.6151
R2450 B.n501 B.n150 10.6151
R2451 B.n501 B.n500 10.6151
R2452 B.n500 B.n499 10.6151
R2453 B.n499 B.n152 10.6151
R2454 B.n495 B.n152 10.6151
R2455 B.n495 B.n494 10.6151
R2456 B.n494 B.n493 10.6151
R2457 B.n493 B.n154 10.6151
R2458 B.n489 B.n154 10.6151
R2459 B.n489 B.n488 10.6151
R2460 B.n488 B.n487 10.6151
R2461 B.n239 B.n1 10.6151
R2462 B.n239 B.n238 10.6151
R2463 B.n243 B.n238 10.6151
R2464 B.n244 B.n243 10.6151
R2465 B.n245 B.n244 10.6151
R2466 B.n245 B.n236 10.6151
R2467 B.n249 B.n236 10.6151
R2468 B.n250 B.n249 10.6151
R2469 B.n251 B.n250 10.6151
R2470 B.n251 B.n234 10.6151
R2471 B.n255 B.n234 10.6151
R2472 B.n256 B.n255 10.6151
R2473 B.n257 B.n256 10.6151
R2474 B.n257 B.n232 10.6151
R2475 B.n261 B.n232 10.6151
R2476 B.n262 B.n261 10.6151
R2477 B.n263 B.n262 10.6151
R2478 B.n263 B.n230 10.6151
R2479 B.n267 B.n230 10.6151
R2480 B.n268 B.n267 10.6151
R2481 B.n269 B.n268 10.6151
R2482 B.n269 B.n228 10.6151
R2483 B.n273 B.n228 10.6151
R2484 B.n274 B.n273 10.6151
R2485 B.n275 B.n274 10.6151
R2486 B.n275 B.n226 10.6151
R2487 B.n279 B.n226 10.6151
R2488 B.n280 B.n279 10.6151
R2489 B.n281 B.n280 10.6151
R2490 B.n281 B.n224 10.6151
R2491 B.n285 B.n224 10.6151
R2492 B.n286 B.n285 10.6151
R2493 B.n287 B.n286 10.6151
R2494 B.n287 B.n222 10.6151
R2495 B.n291 B.n222 10.6151
R2496 B.n292 B.n291 10.6151
R2497 B.n293 B.n292 10.6151
R2498 B.n293 B.n220 10.6151
R2499 B.n297 B.n220 10.6151
R2500 B.n298 B.n297 10.6151
R2501 B.n299 B.n298 10.6151
R2502 B.n299 B.n218 10.6151
R2503 B.n303 B.n218 10.6151
R2504 B.n304 B.n303 10.6151
R2505 B.n305 B.n304 10.6151
R2506 B.n305 B.n216 10.6151
R2507 B.n309 B.n216 10.6151
R2508 B.n310 B.n309 10.6151
R2509 B.n311 B.n310 10.6151
R2510 B.n311 B.n214 10.6151
R2511 B.n315 B.n214 10.6151
R2512 B.n316 B.n315 10.6151
R2513 B.n317 B.n316 10.6151
R2514 B.n317 B.n212 10.6151
R2515 B.n321 B.n212 10.6151
R2516 B.n322 B.n321 10.6151
R2517 B.n323 B.n322 10.6151
R2518 B.n323 B.n210 10.6151
R2519 B.n327 B.n210 10.6151
R2520 B.n328 B.n327 10.6151
R2521 B.n329 B.n328 10.6151
R2522 B.n329 B.n208 10.6151
R2523 B.n333 B.n208 10.6151
R2524 B.n334 B.n333 10.6151
R2525 B.n335 B.n334 10.6151
R2526 B.n335 B.n206 10.6151
R2527 B.n340 B.n339 10.6151
R2528 B.n341 B.n340 10.6151
R2529 B.n341 B.n204 10.6151
R2530 B.n345 B.n204 10.6151
R2531 B.n346 B.n345 10.6151
R2532 B.n347 B.n346 10.6151
R2533 B.n347 B.n202 10.6151
R2534 B.n351 B.n202 10.6151
R2535 B.n352 B.n351 10.6151
R2536 B.n353 B.n352 10.6151
R2537 B.n353 B.n200 10.6151
R2538 B.n357 B.n200 10.6151
R2539 B.n358 B.n357 10.6151
R2540 B.n359 B.n358 10.6151
R2541 B.n359 B.n198 10.6151
R2542 B.n363 B.n198 10.6151
R2543 B.n364 B.n363 10.6151
R2544 B.n365 B.n364 10.6151
R2545 B.n365 B.n196 10.6151
R2546 B.n369 B.n196 10.6151
R2547 B.n370 B.n369 10.6151
R2548 B.n371 B.n370 10.6151
R2549 B.n371 B.n194 10.6151
R2550 B.n375 B.n194 10.6151
R2551 B.n376 B.n375 10.6151
R2552 B.n377 B.n376 10.6151
R2553 B.n377 B.n192 10.6151
R2554 B.n381 B.n192 10.6151
R2555 B.n382 B.n381 10.6151
R2556 B.n383 B.n382 10.6151
R2557 B.n383 B.n190 10.6151
R2558 B.n387 B.n190 10.6151
R2559 B.n388 B.n387 10.6151
R2560 B.n389 B.n388 10.6151
R2561 B.n389 B.n188 10.6151
R2562 B.n393 B.n188 10.6151
R2563 B.n394 B.n393 10.6151
R2564 B.n395 B.n394 10.6151
R2565 B.n395 B.n186 10.6151
R2566 B.n399 B.n186 10.6151
R2567 B.n400 B.n399 10.6151
R2568 B.n404 B.n400 10.6151
R2569 B.n408 B.n184 10.6151
R2570 B.n409 B.n408 10.6151
R2571 B.n410 B.n409 10.6151
R2572 B.n410 B.n182 10.6151
R2573 B.n414 B.n182 10.6151
R2574 B.n415 B.n414 10.6151
R2575 B.n416 B.n415 10.6151
R2576 B.n416 B.n180 10.6151
R2577 B.n420 B.n180 10.6151
R2578 B.n423 B.n422 10.6151
R2579 B.n423 B.n176 10.6151
R2580 B.n427 B.n176 10.6151
R2581 B.n428 B.n427 10.6151
R2582 B.n429 B.n428 10.6151
R2583 B.n429 B.n174 10.6151
R2584 B.n433 B.n174 10.6151
R2585 B.n434 B.n433 10.6151
R2586 B.n435 B.n434 10.6151
R2587 B.n435 B.n172 10.6151
R2588 B.n439 B.n172 10.6151
R2589 B.n440 B.n439 10.6151
R2590 B.n441 B.n440 10.6151
R2591 B.n441 B.n170 10.6151
R2592 B.n445 B.n170 10.6151
R2593 B.n446 B.n445 10.6151
R2594 B.n447 B.n446 10.6151
R2595 B.n447 B.n168 10.6151
R2596 B.n451 B.n168 10.6151
R2597 B.n452 B.n451 10.6151
R2598 B.n453 B.n452 10.6151
R2599 B.n453 B.n166 10.6151
R2600 B.n457 B.n166 10.6151
R2601 B.n458 B.n457 10.6151
R2602 B.n459 B.n458 10.6151
R2603 B.n459 B.n164 10.6151
R2604 B.n463 B.n164 10.6151
R2605 B.n464 B.n463 10.6151
R2606 B.n465 B.n464 10.6151
R2607 B.n465 B.n162 10.6151
R2608 B.n469 B.n162 10.6151
R2609 B.n470 B.n469 10.6151
R2610 B.n471 B.n470 10.6151
R2611 B.n471 B.n160 10.6151
R2612 B.n475 B.n160 10.6151
R2613 B.n476 B.n475 10.6151
R2614 B.n477 B.n476 10.6151
R2615 B.n477 B.n158 10.6151
R2616 B.n481 B.n158 10.6151
R2617 B.n482 B.n481 10.6151
R2618 B.n483 B.n482 10.6151
R2619 B.n483 B.n156 10.6151
R2620 B.n771 B.n770 9.36635
R2621 B.n753 B.n66 9.36635
R2622 B.n404 B.n403 9.36635
R2623 B.n422 B.n421 9.36635
R2624 B.n937 B.n0 8.11757
R2625 B.n937 B.n1 8.11757
R2626 B.n770 B.n769 1.24928
R2627 B.n756 B.n66 1.24928
R2628 B.n403 B.n184 1.24928
R2629 B.n421 B.n420 1.24928
C0 VTAIL w_n5014_n3484# 3.35149f
C1 VDD2 B 2.8336f
C2 VDD1 VN 0.15468f
C3 VTAIL VP 12.309f
C4 VDD1 w_n5014_n3484# 2.99569f
C5 B VN 1.4062f
C6 w_n5014_n3484# B 11.4495f
C7 VDD1 VP 11.97f
C8 VTAIL VDD1 10.790599f
C9 VDD2 VN 11.488501f
C10 B VP 2.50862f
C11 VTAIL B 4.0401f
C12 VDD2 w_n5014_n3484# 3.16211f
C13 w_n5014_n3484# VN 10.850599f
C14 VDD2 VP 0.640066f
C15 VDD1 B 2.69855f
C16 VDD2 VTAIL 10.8448f
C17 VP VN 9.145809f
C18 VTAIL VN 12.294701f
C19 w_n5014_n3484# VP 11.5048f
C20 VDD2 VDD1 2.46087f
C21 VDD2 VSUBS 2.33028f
C22 VDD1 VSUBS 2.156237f
C23 VTAIL VSUBS 1.431258f
C24 VN VSUBS 8.439281f
C25 VP VSUBS 4.833511f
C26 B VSUBS 5.961848f
C27 w_n5014_n3484# VSUBS 0.21486p
C28 B.n0 VSUBS 0.007864f
C29 B.n1 VSUBS 0.007864f
C30 B.n2 VSUBS 0.01163f
C31 B.n3 VSUBS 0.008912f
C32 B.n4 VSUBS 0.008912f
C33 B.n5 VSUBS 0.008912f
C34 B.n6 VSUBS 0.008912f
C35 B.n7 VSUBS 0.008912f
C36 B.n8 VSUBS 0.008912f
C37 B.n9 VSUBS 0.008912f
C38 B.n10 VSUBS 0.008912f
C39 B.n11 VSUBS 0.008912f
C40 B.n12 VSUBS 0.008912f
C41 B.n13 VSUBS 0.008912f
C42 B.n14 VSUBS 0.008912f
C43 B.n15 VSUBS 0.008912f
C44 B.n16 VSUBS 0.008912f
C45 B.n17 VSUBS 0.008912f
C46 B.n18 VSUBS 0.008912f
C47 B.n19 VSUBS 0.008912f
C48 B.n20 VSUBS 0.008912f
C49 B.n21 VSUBS 0.008912f
C50 B.n22 VSUBS 0.008912f
C51 B.n23 VSUBS 0.008912f
C52 B.n24 VSUBS 0.008912f
C53 B.n25 VSUBS 0.008912f
C54 B.n26 VSUBS 0.008912f
C55 B.n27 VSUBS 0.008912f
C56 B.n28 VSUBS 0.008912f
C57 B.n29 VSUBS 0.008912f
C58 B.n30 VSUBS 0.008912f
C59 B.n31 VSUBS 0.008912f
C60 B.n32 VSUBS 0.008912f
C61 B.n33 VSUBS 0.008912f
C62 B.n34 VSUBS 0.008912f
C63 B.n35 VSUBS 0.021175f
C64 B.n36 VSUBS 0.008912f
C65 B.n37 VSUBS 0.008912f
C66 B.n38 VSUBS 0.008912f
C67 B.n39 VSUBS 0.008912f
C68 B.n40 VSUBS 0.008912f
C69 B.n41 VSUBS 0.008912f
C70 B.n42 VSUBS 0.008912f
C71 B.n43 VSUBS 0.008912f
C72 B.n44 VSUBS 0.008912f
C73 B.n45 VSUBS 0.008912f
C74 B.n46 VSUBS 0.008912f
C75 B.n47 VSUBS 0.008912f
C76 B.n48 VSUBS 0.008912f
C77 B.n49 VSUBS 0.008912f
C78 B.n50 VSUBS 0.008912f
C79 B.n51 VSUBS 0.008912f
C80 B.n52 VSUBS 0.008912f
C81 B.n53 VSUBS 0.008912f
C82 B.n54 VSUBS 0.008912f
C83 B.n55 VSUBS 0.008912f
C84 B.n56 VSUBS 0.008912f
C85 B.n57 VSUBS 0.008912f
C86 B.t10 VSUBS 0.284852f
C87 B.t11 VSUBS 0.331313f
C88 B.t9 VSUBS 2.23435f
C89 B.n58 VSUBS 0.527392f
C90 B.n59 VSUBS 0.333456f
C91 B.n60 VSUBS 0.008912f
C92 B.n61 VSUBS 0.008912f
C93 B.n62 VSUBS 0.008912f
C94 B.n63 VSUBS 0.008912f
C95 B.t4 VSUBS 0.284856f
C96 B.t5 VSUBS 0.331317f
C97 B.t3 VSUBS 2.23435f
C98 B.n64 VSUBS 0.527388f
C99 B.n65 VSUBS 0.333452f
C100 B.n66 VSUBS 0.020648f
C101 B.n67 VSUBS 0.008912f
C102 B.n68 VSUBS 0.008912f
C103 B.n69 VSUBS 0.008912f
C104 B.n70 VSUBS 0.008912f
C105 B.n71 VSUBS 0.008912f
C106 B.n72 VSUBS 0.008912f
C107 B.n73 VSUBS 0.008912f
C108 B.n74 VSUBS 0.008912f
C109 B.n75 VSUBS 0.008912f
C110 B.n76 VSUBS 0.008912f
C111 B.n77 VSUBS 0.008912f
C112 B.n78 VSUBS 0.008912f
C113 B.n79 VSUBS 0.008912f
C114 B.n80 VSUBS 0.008912f
C115 B.n81 VSUBS 0.008912f
C116 B.n82 VSUBS 0.008912f
C117 B.n83 VSUBS 0.008912f
C118 B.n84 VSUBS 0.008912f
C119 B.n85 VSUBS 0.008912f
C120 B.n86 VSUBS 0.008912f
C121 B.n87 VSUBS 0.008912f
C122 B.n88 VSUBS 0.021175f
C123 B.n89 VSUBS 0.008912f
C124 B.n90 VSUBS 0.008912f
C125 B.n91 VSUBS 0.008912f
C126 B.n92 VSUBS 0.008912f
C127 B.n93 VSUBS 0.008912f
C128 B.n94 VSUBS 0.008912f
C129 B.n95 VSUBS 0.008912f
C130 B.n96 VSUBS 0.008912f
C131 B.n97 VSUBS 0.008912f
C132 B.n98 VSUBS 0.008912f
C133 B.n99 VSUBS 0.008912f
C134 B.n100 VSUBS 0.008912f
C135 B.n101 VSUBS 0.008912f
C136 B.n102 VSUBS 0.008912f
C137 B.n103 VSUBS 0.008912f
C138 B.n104 VSUBS 0.008912f
C139 B.n105 VSUBS 0.008912f
C140 B.n106 VSUBS 0.008912f
C141 B.n107 VSUBS 0.008912f
C142 B.n108 VSUBS 0.008912f
C143 B.n109 VSUBS 0.008912f
C144 B.n110 VSUBS 0.008912f
C145 B.n111 VSUBS 0.008912f
C146 B.n112 VSUBS 0.008912f
C147 B.n113 VSUBS 0.008912f
C148 B.n114 VSUBS 0.008912f
C149 B.n115 VSUBS 0.008912f
C150 B.n116 VSUBS 0.008912f
C151 B.n117 VSUBS 0.008912f
C152 B.n118 VSUBS 0.008912f
C153 B.n119 VSUBS 0.008912f
C154 B.n120 VSUBS 0.008912f
C155 B.n121 VSUBS 0.008912f
C156 B.n122 VSUBS 0.008912f
C157 B.n123 VSUBS 0.008912f
C158 B.n124 VSUBS 0.008912f
C159 B.n125 VSUBS 0.008912f
C160 B.n126 VSUBS 0.008912f
C161 B.n127 VSUBS 0.008912f
C162 B.n128 VSUBS 0.008912f
C163 B.n129 VSUBS 0.008912f
C164 B.n130 VSUBS 0.008912f
C165 B.n131 VSUBS 0.008912f
C166 B.n132 VSUBS 0.008912f
C167 B.n133 VSUBS 0.008912f
C168 B.n134 VSUBS 0.008912f
C169 B.n135 VSUBS 0.008912f
C170 B.n136 VSUBS 0.008912f
C171 B.n137 VSUBS 0.008912f
C172 B.n138 VSUBS 0.008912f
C173 B.n139 VSUBS 0.008912f
C174 B.n140 VSUBS 0.008912f
C175 B.n141 VSUBS 0.008912f
C176 B.n142 VSUBS 0.008912f
C177 B.n143 VSUBS 0.008912f
C178 B.n144 VSUBS 0.008912f
C179 B.n145 VSUBS 0.008912f
C180 B.n146 VSUBS 0.008912f
C181 B.n147 VSUBS 0.008912f
C182 B.n148 VSUBS 0.008912f
C183 B.n149 VSUBS 0.008912f
C184 B.n150 VSUBS 0.008912f
C185 B.n151 VSUBS 0.008912f
C186 B.n152 VSUBS 0.008912f
C187 B.n153 VSUBS 0.008912f
C188 B.n154 VSUBS 0.008912f
C189 B.n155 VSUBS 0.008912f
C190 B.n156 VSUBS 0.021078f
C191 B.n157 VSUBS 0.008912f
C192 B.n158 VSUBS 0.008912f
C193 B.n159 VSUBS 0.008912f
C194 B.n160 VSUBS 0.008912f
C195 B.n161 VSUBS 0.008912f
C196 B.n162 VSUBS 0.008912f
C197 B.n163 VSUBS 0.008912f
C198 B.n164 VSUBS 0.008912f
C199 B.n165 VSUBS 0.008912f
C200 B.n166 VSUBS 0.008912f
C201 B.n167 VSUBS 0.008912f
C202 B.n168 VSUBS 0.008912f
C203 B.n169 VSUBS 0.008912f
C204 B.n170 VSUBS 0.008912f
C205 B.n171 VSUBS 0.008912f
C206 B.n172 VSUBS 0.008912f
C207 B.n173 VSUBS 0.008912f
C208 B.n174 VSUBS 0.008912f
C209 B.n175 VSUBS 0.008912f
C210 B.n176 VSUBS 0.008912f
C211 B.n177 VSUBS 0.008912f
C212 B.t2 VSUBS 0.284856f
C213 B.t1 VSUBS 0.331317f
C214 B.t0 VSUBS 2.23435f
C215 B.n178 VSUBS 0.527388f
C216 B.n179 VSUBS 0.333452f
C217 B.n180 VSUBS 0.008912f
C218 B.n181 VSUBS 0.008912f
C219 B.n182 VSUBS 0.008912f
C220 B.n183 VSUBS 0.008912f
C221 B.n184 VSUBS 0.00498f
C222 B.n185 VSUBS 0.008912f
C223 B.n186 VSUBS 0.008912f
C224 B.n187 VSUBS 0.008912f
C225 B.n188 VSUBS 0.008912f
C226 B.n189 VSUBS 0.008912f
C227 B.n190 VSUBS 0.008912f
C228 B.n191 VSUBS 0.008912f
C229 B.n192 VSUBS 0.008912f
C230 B.n193 VSUBS 0.008912f
C231 B.n194 VSUBS 0.008912f
C232 B.n195 VSUBS 0.008912f
C233 B.n196 VSUBS 0.008912f
C234 B.n197 VSUBS 0.008912f
C235 B.n198 VSUBS 0.008912f
C236 B.n199 VSUBS 0.008912f
C237 B.n200 VSUBS 0.008912f
C238 B.n201 VSUBS 0.008912f
C239 B.n202 VSUBS 0.008912f
C240 B.n203 VSUBS 0.008912f
C241 B.n204 VSUBS 0.008912f
C242 B.n205 VSUBS 0.008912f
C243 B.n206 VSUBS 0.021175f
C244 B.n207 VSUBS 0.008912f
C245 B.n208 VSUBS 0.008912f
C246 B.n209 VSUBS 0.008912f
C247 B.n210 VSUBS 0.008912f
C248 B.n211 VSUBS 0.008912f
C249 B.n212 VSUBS 0.008912f
C250 B.n213 VSUBS 0.008912f
C251 B.n214 VSUBS 0.008912f
C252 B.n215 VSUBS 0.008912f
C253 B.n216 VSUBS 0.008912f
C254 B.n217 VSUBS 0.008912f
C255 B.n218 VSUBS 0.008912f
C256 B.n219 VSUBS 0.008912f
C257 B.n220 VSUBS 0.008912f
C258 B.n221 VSUBS 0.008912f
C259 B.n222 VSUBS 0.008912f
C260 B.n223 VSUBS 0.008912f
C261 B.n224 VSUBS 0.008912f
C262 B.n225 VSUBS 0.008912f
C263 B.n226 VSUBS 0.008912f
C264 B.n227 VSUBS 0.008912f
C265 B.n228 VSUBS 0.008912f
C266 B.n229 VSUBS 0.008912f
C267 B.n230 VSUBS 0.008912f
C268 B.n231 VSUBS 0.008912f
C269 B.n232 VSUBS 0.008912f
C270 B.n233 VSUBS 0.008912f
C271 B.n234 VSUBS 0.008912f
C272 B.n235 VSUBS 0.008912f
C273 B.n236 VSUBS 0.008912f
C274 B.n237 VSUBS 0.008912f
C275 B.n238 VSUBS 0.008912f
C276 B.n239 VSUBS 0.008912f
C277 B.n240 VSUBS 0.008912f
C278 B.n241 VSUBS 0.008912f
C279 B.n242 VSUBS 0.008912f
C280 B.n243 VSUBS 0.008912f
C281 B.n244 VSUBS 0.008912f
C282 B.n245 VSUBS 0.008912f
C283 B.n246 VSUBS 0.008912f
C284 B.n247 VSUBS 0.008912f
C285 B.n248 VSUBS 0.008912f
C286 B.n249 VSUBS 0.008912f
C287 B.n250 VSUBS 0.008912f
C288 B.n251 VSUBS 0.008912f
C289 B.n252 VSUBS 0.008912f
C290 B.n253 VSUBS 0.008912f
C291 B.n254 VSUBS 0.008912f
C292 B.n255 VSUBS 0.008912f
C293 B.n256 VSUBS 0.008912f
C294 B.n257 VSUBS 0.008912f
C295 B.n258 VSUBS 0.008912f
C296 B.n259 VSUBS 0.008912f
C297 B.n260 VSUBS 0.008912f
C298 B.n261 VSUBS 0.008912f
C299 B.n262 VSUBS 0.008912f
C300 B.n263 VSUBS 0.008912f
C301 B.n264 VSUBS 0.008912f
C302 B.n265 VSUBS 0.008912f
C303 B.n266 VSUBS 0.008912f
C304 B.n267 VSUBS 0.008912f
C305 B.n268 VSUBS 0.008912f
C306 B.n269 VSUBS 0.008912f
C307 B.n270 VSUBS 0.008912f
C308 B.n271 VSUBS 0.008912f
C309 B.n272 VSUBS 0.008912f
C310 B.n273 VSUBS 0.008912f
C311 B.n274 VSUBS 0.008912f
C312 B.n275 VSUBS 0.008912f
C313 B.n276 VSUBS 0.008912f
C314 B.n277 VSUBS 0.008912f
C315 B.n278 VSUBS 0.008912f
C316 B.n279 VSUBS 0.008912f
C317 B.n280 VSUBS 0.008912f
C318 B.n281 VSUBS 0.008912f
C319 B.n282 VSUBS 0.008912f
C320 B.n283 VSUBS 0.008912f
C321 B.n284 VSUBS 0.008912f
C322 B.n285 VSUBS 0.008912f
C323 B.n286 VSUBS 0.008912f
C324 B.n287 VSUBS 0.008912f
C325 B.n288 VSUBS 0.008912f
C326 B.n289 VSUBS 0.008912f
C327 B.n290 VSUBS 0.008912f
C328 B.n291 VSUBS 0.008912f
C329 B.n292 VSUBS 0.008912f
C330 B.n293 VSUBS 0.008912f
C331 B.n294 VSUBS 0.008912f
C332 B.n295 VSUBS 0.008912f
C333 B.n296 VSUBS 0.008912f
C334 B.n297 VSUBS 0.008912f
C335 B.n298 VSUBS 0.008912f
C336 B.n299 VSUBS 0.008912f
C337 B.n300 VSUBS 0.008912f
C338 B.n301 VSUBS 0.008912f
C339 B.n302 VSUBS 0.008912f
C340 B.n303 VSUBS 0.008912f
C341 B.n304 VSUBS 0.008912f
C342 B.n305 VSUBS 0.008912f
C343 B.n306 VSUBS 0.008912f
C344 B.n307 VSUBS 0.008912f
C345 B.n308 VSUBS 0.008912f
C346 B.n309 VSUBS 0.008912f
C347 B.n310 VSUBS 0.008912f
C348 B.n311 VSUBS 0.008912f
C349 B.n312 VSUBS 0.008912f
C350 B.n313 VSUBS 0.008912f
C351 B.n314 VSUBS 0.008912f
C352 B.n315 VSUBS 0.008912f
C353 B.n316 VSUBS 0.008912f
C354 B.n317 VSUBS 0.008912f
C355 B.n318 VSUBS 0.008912f
C356 B.n319 VSUBS 0.008912f
C357 B.n320 VSUBS 0.008912f
C358 B.n321 VSUBS 0.008912f
C359 B.n322 VSUBS 0.008912f
C360 B.n323 VSUBS 0.008912f
C361 B.n324 VSUBS 0.008912f
C362 B.n325 VSUBS 0.008912f
C363 B.n326 VSUBS 0.008912f
C364 B.n327 VSUBS 0.008912f
C365 B.n328 VSUBS 0.008912f
C366 B.n329 VSUBS 0.008912f
C367 B.n330 VSUBS 0.008912f
C368 B.n331 VSUBS 0.008912f
C369 B.n332 VSUBS 0.008912f
C370 B.n333 VSUBS 0.008912f
C371 B.n334 VSUBS 0.008912f
C372 B.n335 VSUBS 0.008912f
C373 B.n336 VSUBS 0.008912f
C374 B.n337 VSUBS 0.021175f
C375 B.n338 VSUBS 0.022075f
C376 B.n339 VSUBS 0.022075f
C377 B.n340 VSUBS 0.008912f
C378 B.n341 VSUBS 0.008912f
C379 B.n342 VSUBS 0.008912f
C380 B.n343 VSUBS 0.008912f
C381 B.n344 VSUBS 0.008912f
C382 B.n345 VSUBS 0.008912f
C383 B.n346 VSUBS 0.008912f
C384 B.n347 VSUBS 0.008912f
C385 B.n348 VSUBS 0.008912f
C386 B.n349 VSUBS 0.008912f
C387 B.n350 VSUBS 0.008912f
C388 B.n351 VSUBS 0.008912f
C389 B.n352 VSUBS 0.008912f
C390 B.n353 VSUBS 0.008912f
C391 B.n354 VSUBS 0.008912f
C392 B.n355 VSUBS 0.008912f
C393 B.n356 VSUBS 0.008912f
C394 B.n357 VSUBS 0.008912f
C395 B.n358 VSUBS 0.008912f
C396 B.n359 VSUBS 0.008912f
C397 B.n360 VSUBS 0.008912f
C398 B.n361 VSUBS 0.008912f
C399 B.n362 VSUBS 0.008912f
C400 B.n363 VSUBS 0.008912f
C401 B.n364 VSUBS 0.008912f
C402 B.n365 VSUBS 0.008912f
C403 B.n366 VSUBS 0.008912f
C404 B.n367 VSUBS 0.008912f
C405 B.n368 VSUBS 0.008912f
C406 B.n369 VSUBS 0.008912f
C407 B.n370 VSUBS 0.008912f
C408 B.n371 VSUBS 0.008912f
C409 B.n372 VSUBS 0.008912f
C410 B.n373 VSUBS 0.008912f
C411 B.n374 VSUBS 0.008912f
C412 B.n375 VSUBS 0.008912f
C413 B.n376 VSUBS 0.008912f
C414 B.n377 VSUBS 0.008912f
C415 B.n378 VSUBS 0.008912f
C416 B.n379 VSUBS 0.008912f
C417 B.n380 VSUBS 0.008912f
C418 B.n381 VSUBS 0.008912f
C419 B.n382 VSUBS 0.008912f
C420 B.n383 VSUBS 0.008912f
C421 B.n384 VSUBS 0.008912f
C422 B.n385 VSUBS 0.008912f
C423 B.n386 VSUBS 0.008912f
C424 B.n387 VSUBS 0.008912f
C425 B.n388 VSUBS 0.008912f
C426 B.n389 VSUBS 0.008912f
C427 B.n390 VSUBS 0.008912f
C428 B.n391 VSUBS 0.008912f
C429 B.n392 VSUBS 0.008912f
C430 B.n393 VSUBS 0.008912f
C431 B.n394 VSUBS 0.008912f
C432 B.n395 VSUBS 0.008912f
C433 B.n396 VSUBS 0.008912f
C434 B.n397 VSUBS 0.008912f
C435 B.n398 VSUBS 0.008912f
C436 B.n399 VSUBS 0.008912f
C437 B.n400 VSUBS 0.008912f
C438 B.t8 VSUBS 0.284852f
C439 B.t7 VSUBS 0.331313f
C440 B.t6 VSUBS 2.23435f
C441 B.n401 VSUBS 0.527392f
C442 B.n402 VSUBS 0.333456f
C443 B.n403 VSUBS 0.020648f
C444 B.n404 VSUBS 0.008388f
C445 B.n405 VSUBS 0.008912f
C446 B.n406 VSUBS 0.008912f
C447 B.n407 VSUBS 0.008912f
C448 B.n408 VSUBS 0.008912f
C449 B.n409 VSUBS 0.008912f
C450 B.n410 VSUBS 0.008912f
C451 B.n411 VSUBS 0.008912f
C452 B.n412 VSUBS 0.008912f
C453 B.n413 VSUBS 0.008912f
C454 B.n414 VSUBS 0.008912f
C455 B.n415 VSUBS 0.008912f
C456 B.n416 VSUBS 0.008912f
C457 B.n417 VSUBS 0.008912f
C458 B.n418 VSUBS 0.008912f
C459 B.n419 VSUBS 0.008912f
C460 B.n420 VSUBS 0.00498f
C461 B.n421 VSUBS 0.020648f
C462 B.n422 VSUBS 0.008388f
C463 B.n423 VSUBS 0.008912f
C464 B.n424 VSUBS 0.008912f
C465 B.n425 VSUBS 0.008912f
C466 B.n426 VSUBS 0.008912f
C467 B.n427 VSUBS 0.008912f
C468 B.n428 VSUBS 0.008912f
C469 B.n429 VSUBS 0.008912f
C470 B.n430 VSUBS 0.008912f
C471 B.n431 VSUBS 0.008912f
C472 B.n432 VSUBS 0.008912f
C473 B.n433 VSUBS 0.008912f
C474 B.n434 VSUBS 0.008912f
C475 B.n435 VSUBS 0.008912f
C476 B.n436 VSUBS 0.008912f
C477 B.n437 VSUBS 0.008912f
C478 B.n438 VSUBS 0.008912f
C479 B.n439 VSUBS 0.008912f
C480 B.n440 VSUBS 0.008912f
C481 B.n441 VSUBS 0.008912f
C482 B.n442 VSUBS 0.008912f
C483 B.n443 VSUBS 0.008912f
C484 B.n444 VSUBS 0.008912f
C485 B.n445 VSUBS 0.008912f
C486 B.n446 VSUBS 0.008912f
C487 B.n447 VSUBS 0.008912f
C488 B.n448 VSUBS 0.008912f
C489 B.n449 VSUBS 0.008912f
C490 B.n450 VSUBS 0.008912f
C491 B.n451 VSUBS 0.008912f
C492 B.n452 VSUBS 0.008912f
C493 B.n453 VSUBS 0.008912f
C494 B.n454 VSUBS 0.008912f
C495 B.n455 VSUBS 0.008912f
C496 B.n456 VSUBS 0.008912f
C497 B.n457 VSUBS 0.008912f
C498 B.n458 VSUBS 0.008912f
C499 B.n459 VSUBS 0.008912f
C500 B.n460 VSUBS 0.008912f
C501 B.n461 VSUBS 0.008912f
C502 B.n462 VSUBS 0.008912f
C503 B.n463 VSUBS 0.008912f
C504 B.n464 VSUBS 0.008912f
C505 B.n465 VSUBS 0.008912f
C506 B.n466 VSUBS 0.008912f
C507 B.n467 VSUBS 0.008912f
C508 B.n468 VSUBS 0.008912f
C509 B.n469 VSUBS 0.008912f
C510 B.n470 VSUBS 0.008912f
C511 B.n471 VSUBS 0.008912f
C512 B.n472 VSUBS 0.008912f
C513 B.n473 VSUBS 0.008912f
C514 B.n474 VSUBS 0.008912f
C515 B.n475 VSUBS 0.008912f
C516 B.n476 VSUBS 0.008912f
C517 B.n477 VSUBS 0.008912f
C518 B.n478 VSUBS 0.008912f
C519 B.n479 VSUBS 0.008912f
C520 B.n480 VSUBS 0.008912f
C521 B.n481 VSUBS 0.008912f
C522 B.n482 VSUBS 0.008912f
C523 B.n483 VSUBS 0.008912f
C524 B.n484 VSUBS 0.008912f
C525 B.n485 VSUBS 0.022075f
C526 B.n486 VSUBS 0.021175f
C527 B.n487 VSUBS 0.022172f
C528 B.n488 VSUBS 0.008912f
C529 B.n489 VSUBS 0.008912f
C530 B.n490 VSUBS 0.008912f
C531 B.n491 VSUBS 0.008912f
C532 B.n492 VSUBS 0.008912f
C533 B.n493 VSUBS 0.008912f
C534 B.n494 VSUBS 0.008912f
C535 B.n495 VSUBS 0.008912f
C536 B.n496 VSUBS 0.008912f
C537 B.n497 VSUBS 0.008912f
C538 B.n498 VSUBS 0.008912f
C539 B.n499 VSUBS 0.008912f
C540 B.n500 VSUBS 0.008912f
C541 B.n501 VSUBS 0.008912f
C542 B.n502 VSUBS 0.008912f
C543 B.n503 VSUBS 0.008912f
C544 B.n504 VSUBS 0.008912f
C545 B.n505 VSUBS 0.008912f
C546 B.n506 VSUBS 0.008912f
C547 B.n507 VSUBS 0.008912f
C548 B.n508 VSUBS 0.008912f
C549 B.n509 VSUBS 0.008912f
C550 B.n510 VSUBS 0.008912f
C551 B.n511 VSUBS 0.008912f
C552 B.n512 VSUBS 0.008912f
C553 B.n513 VSUBS 0.008912f
C554 B.n514 VSUBS 0.008912f
C555 B.n515 VSUBS 0.008912f
C556 B.n516 VSUBS 0.008912f
C557 B.n517 VSUBS 0.008912f
C558 B.n518 VSUBS 0.008912f
C559 B.n519 VSUBS 0.008912f
C560 B.n520 VSUBS 0.008912f
C561 B.n521 VSUBS 0.008912f
C562 B.n522 VSUBS 0.008912f
C563 B.n523 VSUBS 0.008912f
C564 B.n524 VSUBS 0.008912f
C565 B.n525 VSUBS 0.008912f
C566 B.n526 VSUBS 0.008912f
C567 B.n527 VSUBS 0.008912f
C568 B.n528 VSUBS 0.008912f
C569 B.n529 VSUBS 0.008912f
C570 B.n530 VSUBS 0.008912f
C571 B.n531 VSUBS 0.008912f
C572 B.n532 VSUBS 0.008912f
C573 B.n533 VSUBS 0.008912f
C574 B.n534 VSUBS 0.008912f
C575 B.n535 VSUBS 0.008912f
C576 B.n536 VSUBS 0.008912f
C577 B.n537 VSUBS 0.008912f
C578 B.n538 VSUBS 0.008912f
C579 B.n539 VSUBS 0.008912f
C580 B.n540 VSUBS 0.008912f
C581 B.n541 VSUBS 0.008912f
C582 B.n542 VSUBS 0.008912f
C583 B.n543 VSUBS 0.008912f
C584 B.n544 VSUBS 0.008912f
C585 B.n545 VSUBS 0.008912f
C586 B.n546 VSUBS 0.008912f
C587 B.n547 VSUBS 0.008912f
C588 B.n548 VSUBS 0.008912f
C589 B.n549 VSUBS 0.008912f
C590 B.n550 VSUBS 0.008912f
C591 B.n551 VSUBS 0.008912f
C592 B.n552 VSUBS 0.008912f
C593 B.n553 VSUBS 0.008912f
C594 B.n554 VSUBS 0.008912f
C595 B.n555 VSUBS 0.008912f
C596 B.n556 VSUBS 0.008912f
C597 B.n557 VSUBS 0.008912f
C598 B.n558 VSUBS 0.008912f
C599 B.n559 VSUBS 0.008912f
C600 B.n560 VSUBS 0.008912f
C601 B.n561 VSUBS 0.008912f
C602 B.n562 VSUBS 0.008912f
C603 B.n563 VSUBS 0.008912f
C604 B.n564 VSUBS 0.008912f
C605 B.n565 VSUBS 0.008912f
C606 B.n566 VSUBS 0.008912f
C607 B.n567 VSUBS 0.008912f
C608 B.n568 VSUBS 0.008912f
C609 B.n569 VSUBS 0.008912f
C610 B.n570 VSUBS 0.008912f
C611 B.n571 VSUBS 0.008912f
C612 B.n572 VSUBS 0.008912f
C613 B.n573 VSUBS 0.008912f
C614 B.n574 VSUBS 0.008912f
C615 B.n575 VSUBS 0.008912f
C616 B.n576 VSUBS 0.008912f
C617 B.n577 VSUBS 0.008912f
C618 B.n578 VSUBS 0.008912f
C619 B.n579 VSUBS 0.008912f
C620 B.n580 VSUBS 0.008912f
C621 B.n581 VSUBS 0.008912f
C622 B.n582 VSUBS 0.008912f
C623 B.n583 VSUBS 0.008912f
C624 B.n584 VSUBS 0.008912f
C625 B.n585 VSUBS 0.008912f
C626 B.n586 VSUBS 0.008912f
C627 B.n587 VSUBS 0.008912f
C628 B.n588 VSUBS 0.008912f
C629 B.n589 VSUBS 0.008912f
C630 B.n590 VSUBS 0.008912f
C631 B.n591 VSUBS 0.008912f
C632 B.n592 VSUBS 0.008912f
C633 B.n593 VSUBS 0.008912f
C634 B.n594 VSUBS 0.008912f
C635 B.n595 VSUBS 0.008912f
C636 B.n596 VSUBS 0.008912f
C637 B.n597 VSUBS 0.008912f
C638 B.n598 VSUBS 0.008912f
C639 B.n599 VSUBS 0.008912f
C640 B.n600 VSUBS 0.008912f
C641 B.n601 VSUBS 0.008912f
C642 B.n602 VSUBS 0.008912f
C643 B.n603 VSUBS 0.008912f
C644 B.n604 VSUBS 0.008912f
C645 B.n605 VSUBS 0.008912f
C646 B.n606 VSUBS 0.008912f
C647 B.n607 VSUBS 0.008912f
C648 B.n608 VSUBS 0.008912f
C649 B.n609 VSUBS 0.008912f
C650 B.n610 VSUBS 0.008912f
C651 B.n611 VSUBS 0.008912f
C652 B.n612 VSUBS 0.008912f
C653 B.n613 VSUBS 0.008912f
C654 B.n614 VSUBS 0.008912f
C655 B.n615 VSUBS 0.008912f
C656 B.n616 VSUBS 0.008912f
C657 B.n617 VSUBS 0.008912f
C658 B.n618 VSUBS 0.008912f
C659 B.n619 VSUBS 0.008912f
C660 B.n620 VSUBS 0.008912f
C661 B.n621 VSUBS 0.008912f
C662 B.n622 VSUBS 0.008912f
C663 B.n623 VSUBS 0.008912f
C664 B.n624 VSUBS 0.008912f
C665 B.n625 VSUBS 0.008912f
C666 B.n626 VSUBS 0.008912f
C667 B.n627 VSUBS 0.008912f
C668 B.n628 VSUBS 0.008912f
C669 B.n629 VSUBS 0.008912f
C670 B.n630 VSUBS 0.008912f
C671 B.n631 VSUBS 0.008912f
C672 B.n632 VSUBS 0.008912f
C673 B.n633 VSUBS 0.008912f
C674 B.n634 VSUBS 0.008912f
C675 B.n635 VSUBS 0.008912f
C676 B.n636 VSUBS 0.008912f
C677 B.n637 VSUBS 0.008912f
C678 B.n638 VSUBS 0.008912f
C679 B.n639 VSUBS 0.008912f
C680 B.n640 VSUBS 0.008912f
C681 B.n641 VSUBS 0.008912f
C682 B.n642 VSUBS 0.008912f
C683 B.n643 VSUBS 0.008912f
C684 B.n644 VSUBS 0.008912f
C685 B.n645 VSUBS 0.008912f
C686 B.n646 VSUBS 0.008912f
C687 B.n647 VSUBS 0.008912f
C688 B.n648 VSUBS 0.008912f
C689 B.n649 VSUBS 0.008912f
C690 B.n650 VSUBS 0.008912f
C691 B.n651 VSUBS 0.008912f
C692 B.n652 VSUBS 0.008912f
C693 B.n653 VSUBS 0.008912f
C694 B.n654 VSUBS 0.008912f
C695 B.n655 VSUBS 0.008912f
C696 B.n656 VSUBS 0.008912f
C697 B.n657 VSUBS 0.008912f
C698 B.n658 VSUBS 0.008912f
C699 B.n659 VSUBS 0.008912f
C700 B.n660 VSUBS 0.008912f
C701 B.n661 VSUBS 0.008912f
C702 B.n662 VSUBS 0.008912f
C703 B.n663 VSUBS 0.008912f
C704 B.n664 VSUBS 0.008912f
C705 B.n665 VSUBS 0.008912f
C706 B.n666 VSUBS 0.008912f
C707 B.n667 VSUBS 0.008912f
C708 B.n668 VSUBS 0.008912f
C709 B.n669 VSUBS 0.008912f
C710 B.n670 VSUBS 0.008912f
C711 B.n671 VSUBS 0.008912f
C712 B.n672 VSUBS 0.008912f
C713 B.n673 VSUBS 0.008912f
C714 B.n674 VSUBS 0.008912f
C715 B.n675 VSUBS 0.008912f
C716 B.n676 VSUBS 0.008912f
C717 B.n677 VSUBS 0.008912f
C718 B.n678 VSUBS 0.008912f
C719 B.n679 VSUBS 0.008912f
C720 B.n680 VSUBS 0.008912f
C721 B.n681 VSUBS 0.008912f
C722 B.n682 VSUBS 0.008912f
C723 B.n683 VSUBS 0.008912f
C724 B.n684 VSUBS 0.008912f
C725 B.n685 VSUBS 0.008912f
C726 B.n686 VSUBS 0.008912f
C727 B.n687 VSUBS 0.008912f
C728 B.n688 VSUBS 0.008912f
C729 B.n689 VSUBS 0.021175f
C730 B.n690 VSUBS 0.022075f
C731 B.n691 VSUBS 0.022075f
C732 B.n692 VSUBS 0.008912f
C733 B.n693 VSUBS 0.008912f
C734 B.n694 VSUBS 0.008912f
C735 B.n695 VSUBS 0.008912f
C736 B.n696 VSUBS 0.008912f
C737 B.n697 VSUBS 0.008912f
C738 B.n698 VSUBS 0.008912f
C739 B.n699 VSUBS 0.008912f
C740 B.n700 VSUBS 0.008912f
C741 B.n701 VSUBS 0.008912f
C742 B.n702 VSUBS 0.008912f
C743 B.n703 VSUBS 0.008912f
C744 B.n704 VSUBS 0.008912f
C745 B.n705 VSUBS 0.008912f
C746 B.n706 VSUBS 0.008912f
C747 B.n707 VSUBS 0.008912f
C748 B.n708 VSUBS 0.008912f
C749 B.n709 VSUBS 0.008912f
C750 B.n710 VSUBS 0.008912f
C751 B.n711 VSUBS 0.008912f
C752 B.n712 VSUBS 0.008912f
C753 B.n713 VSUBS 0.008912f
C754 B.n714 VSUBS 0.008912f
C755 B.n715 VSUBS 0.008912f
C756 B.n716 VSUBS 0.008912f
C757 B.n717 VSUBS 0.008912f
C758 B.n718 VSUBS 0.008912f
C759 B.n719 VSUBS 0.008912f
C760 B.n720 VSUBS 0.008912f
C761 B.n721 VSUBS 0.008912f
C762 B.n722 VSUBS 0.008912f
C763 B.n723 VSUBS 0.008912f
C764 B.n724 VSUBS 0.008912f
C765 B.n725 VSUBS 0.008912f
C766 B.n726 VSUBS 0.008912f
C767 B.n727 VSUBS 0.008912f
C768 B.n728 VSUBS 0.008912f
C769 B.n729 VSUBS 0.008912f
C770 B.n730 VSUBS 0.008912f
C771 B.n731 VSUBS 0.008912f
C772 B.n732 VSUBS 0.008912f
C773 B.n733 VSUBS 0.008912f
C774 B.n734 VSUBS 0.008912f
C775 B.n735 VSUBS 0.008912f
C776 B.n736 VSUBS 0.008912f
C777 B.n737 VSUBS 0.008912f
C778 B.n738 VSUBS 0.008912f
C779 B.n739 VSUBS 0.008912f
C780 B.n740 VSUBS 0.008912f
C781 B.n741 VSUBS 0.008912f
C782 B.n742 VSUBS 0.008912f
C783 B.n743 VSUBS 0.008912f
C784 B.n744 VSUBS 0.008912f
C785 B.n745 VSUBS 0.008912f
C786 B.n746 VSUBS 0.008912f
C787 B.n747 VSUBS 0.008912f
C788 B.n748 VSUBS 0.008912f
C789 B.n749 VSUBS 0.008912f
C790 B.n750 VSUBS 0.008912f
C791 B.n751 VSUBS 0.008912f
C792 B.n752 VSUBS 0.008912f
C793 B.n753 VSUBS 0.008388f
C794 B.n754 VSUBS 0.008912f
C795 B.n755 VSUBS 0.008912f
C796 B.n756 VSUBS 0.00498f
C797 B.n757 VSUBS 0.008912f
C798 B.n758 VSUBS 0.008912f
C799 B.n759 VSUBS 0.008912f
C800 B.n760 VSUBS 0.008912f
C801 B.n761 VSUBS 0.008912f
C802 B.n762 VSUBS 0.008912f
C803 B.n763 VSUBS 0.008912f
C804 B.n764 VSUBS 0.008912f
C805 B.n765 VSUBS 0.008912f
C806 B.n766 VSUBS 0.008912f
C807 B.n767 VSUBS 0.008912f
C808 B.n768 VSUBS 0.008912f
C809 B.n769 VSUBS 0.00498f
C810 B.n770 VSUBS 0.020648f
C811 B.n771 VSUBS 0.008388f
C812 B.n772 VSUBS 0.008912f
C813 B.n773 VSUBS 0.008912f
C814 B.n774 VSUBS 0.008912f
C815 B.n775 VSUBS 0.008912f
C816 B.n776 VSUBS 0.008912f
C817 B.n777 VSUBS 0.008912f
C818 B.n778 VSUBS 0.008912f
C819 B.n779 VSUBS 0.008912f
C820 B.n780 VSUBS 0.008912f
C821 B.n781 VSUBS 0.008912f
C822 B.n782 VSUBS 0.008912f
C823 B.n783 VSUBS 0.008912f
C824 B.n784 VSUBS 0.008912f
C825 B.n785 VSUBS 0.008912f
C826 B.n786 VSUBS 0.008912f
C827 B.n787 VSUBS 0.008912f
C828 B.n788 VSUBS 0.008912f
C829 B.n789 VSUBS 0.008912f
C830 B.n790 VSUBS 0.008912f
C831 B.n791 VSUBS 0.008912f
C832 B.n792 VSUBS 0.008912f
C833 B.n793 VSUBS 0.008912f
C834 B.n794 VSUBS 0.008912f
C835 B.n795 VSUBS 0.008912f
C836 B.n796 VSUBS 0.008912f
C837 B.n797 VSUBS 0.008912f
C838 B.n798 VSUBS 0.008912f
C839 B.n799 VSUBS 0.008912f
C840 B.n800 VSUBS 0.008912f
C841 B.n801 VSUBS 0.008912f
C842 B.n802 VSUBS 0.008912f
C843 B.n803 VSUBS 0.008912f
C844 B.n804 VSUBS 0.008912f
C845 B.n805 VSUBS 0.008912f
C846 B.n806 VSUBS 0.008912f
C847 B.n807 VSUBS 0.008912f
C848 B.n808 VSUBS 0.008912f
C849 B.n809 VSUBS 0.008912f
C850 B.n810 VSUBS 0.008912f
C851 B.n811 VSUBS 0.008912f
C852 B.n812 VSUBS 0.008912f
C853 B.n813 VSUBS 0.008912f
C854 B.n814 VSUBS 0.008912f
C855 B.n815 VSUBS 0.008912f
C856 B.n816 VSUBS 0.008912f
C857 B.n817 VSUBS 0.008912f
C858 B.n818 VSUBS 0.008912f
C859 B.n819 VSUBS 0.008912f
C860 B.n820 VSUBS 0.008912f
C861 B.n821 VSUBS 0.008912f
C862 B.n822 VSUBS 0.008912f
C863 B.n823 VSUBS 0.008912f
C864 B.n824 VSUBS 0.008912f
C865 B.n825 VSUBS 0.008912f
C866 B.n826 VSUBS 0.008912f
C867 B.n827 VSUBS 0.008912f
C868 B.n828 VSUBS 0.008912f
C869 B.n829 VSUBS 0.008912f
C870 B.n830 VSUBS 0.008912f
C871 B.n831 VSUBS 0.008912f
C872 B.n832 VSUBS 0.008912f
C873 B.n833 VSUBS 0.008912f
C874 B.n834 VSUBS 0.022075f
C875 B.n835 VSUBS 0.022075f
C876 B.n836 VSUBS 0.021175f
C877 B.n837 VSUBS 0.008912f
C878 B.n838 VSUBS 0.008912f
C879 B.n839 VSUBS 0.008912f
C880 B.n840 VSUBS 0.008912f
C881 B.n841 VSUBS 0.008912f
C882 B.n842 VSUBS 0.008912f
C883 B.n843 VSUBS 0.008912f
C884 B.n844 VSUBS 0.008912f
C885 B.n845 VSUBS 0.008912f
C886 B.n846 VSUBS 0.008912f
C887 B.n847 VSUBS 0.008912f
C888 B.n848 VSUBS 0.008912f
C889 B.n849 VSUBS 0.008912f
C890 B.n850 VSUBS 0.008912f
C891 B.n851 VSUBS 0.008912f
C892 B.n852 VSUBS 0.008912f
C893 B.n853 VSUBS 0.008912f
C894 B.n854 VSUBS 0.008912f
C895 B.n855 VSUBS 0.008912f
C896 B.n856 VSUBS 0.008912f
C897 B.n857 VSUBS 0.008912f
C898 B.n858 VSUBS 0.008912f
C899 B.n859 VSUBS 0.008912f
C900 B.n860 VSUBS 0.008912f
C901 B.n861 VSUBS 0.008912f
C902 B.n862 VSUBS 0.008912f
C903 B.n863 VSUBS 0.008912f
C904 B.n864 VSUBS 0.008912f
C905 B.n865 VSUBS 0.008912f
C906 B.n866 VSUBS 0.008912f
C907 B.n867 VSUBS 0.008912f
C908 B.n868 VSUBS 0.008912f
C909 B.n869 VSUBS 0.008912f
C910 B.n870 VSUBS 0.008912f
C911 B.n871 VSUBS 0.008912f
C912 B.n872 VSUBS 0.008912f
C913 B.n873 VSUBS 0.008912f
C914 B.n874 VSUBS 0.008912f
C915 B.n875 VSUBS 0.008912f
C916 B.n876 VSUBS 0.008912f
C917 B.n877 VSUBS 0.008912f
C918 B.n878 VSUBS 0.008912f
C919 B.n879 VSUBS 0.008912f
C920 B.n880 VSUBS 0.008912f
C921 B.n881 VSUBS 0.008912f
C922 B.n882 VSUBS 0.008912f
C923 B.n883 VSUBS 0.008912f
C924 B.n884 VSUBS 0.008912f
C925 B.n885 VSUBS 0.008912f
C926 B.n886 VSUBS 0.008912f
C927 B.n887 VSUBS 0.008912f
C928 B.n888 VSUBS 0.008912f
C929 B.n889 VSUBS 0.008912f
C930 B.n890 VSUBS 0.008912f
C931 B.n891 VSUBS 0.008912f
C932 B.n892 VSUBS 0.008912f
C933 B.n893 VSUBS 0.008912f
C934 B.n894 VSUBS 0.008912f
C935 B.n895 VSUBS 0.008912f
C936 B.n896 VSUBS 0.008912f
C937 B.n897 VSUBS 0.008912f
C938 B.n898 VSUBS 0.008912f
C939 B.n899 VSUBS 0.008912f
C940 B.n900 VSUBS 0.008912f
C941 B.n901 VSUBS 0.008912f
C942 B.n902 VSUBS 0.008912f
C943 B.n903 VSUBS 0.008912f
C944 B.n904 VSUBS 0.008912f
C945 B.n905 VSUBS 0.008912f
C946 B.n906 VSUBS 0.008912f
C947 B.n907 VSUBS 0.008912f
C948 B.n908 VSUBS 0.008912f
C949 B.n909 VSUBS 0.008912f
C950 B.n910 VSUBS 0.008912f
C951 B.n911 VSUBS 0.008912f
C952 B.n912 VSUBS 0.008912f
C953 B.n913 VSUBS 0.008912f
C954 B.n914 VSUBS 0.008912f
C955 B.n915 VSUBS 0.008912f
C956 B.n916 VSUBS 0.008912f
C957 B.n917 VSUBS 0.008912f
C958 B.n918 VSUBS 0.008912f
C959 B.n919 VSUBS 0.008912f
C960 B.n920 VSUBS 0.008912f
C961 B.n921 VSUBS 0.008912f
C962 B.n922 VSUBS 0.008912f
C963 B.n923 VSUBS 0.008912f
C964 B.n924 VSUBS 0.008912f
C965 B.n925 VSUBS 0.008912f
C966 B.n926 VSUBS 0.008912f
C967 B.n927 VSUBS 0.008912f
C968 B.n928 VSUBS 0.008912f
C969 B.n929 VSUBS 0.008912f
C970 B.n930 VSUBS 0.008912f
C971 B.n931 VSUBS 0.008912f
C972 B.n932 VSUBS 0.008912f
C973 B.n933 VSUBS 0.008912f
C974 B.n934 VSUBS 0.008912f
C975 B.n935 VSUBS 0.01163f
C976 B.n936 VSUBS 0.012389f
C977 B.n937 VSUBS 0.024636f
C978 VDD2.n0 VSUBS 0.016991f
C979 VDD2.n1 VSUBS 0.038432f
C980 VDD2.n2 VSUBS 0.017216f
C981 VDD2.n3 VSUBS 0.030259f
C982 VDD2.n4 VSUBS 0.01626f
C983 VDD2.n5 VSUBS 0.038432f
C984 VDD2.n6 VSUBS 0.017216f
C985 VDD2.n7 VSUBS 0.030259f
C986 VDD2.n8 VSUBS 0.01626f
C987 VDD2.n9 VSUBS 0.038432f
C988 VDD2.n10 VSUBS 0.017216f
C989 VDD2.n11 VSUBS 0.030259f
C990 VDD2.n12 VSUBS 0.01626f
C991 VDD2.n13 VSUBS 0.038432f
C992 VDD2.n14 VSUBS 0.017216f
C993 VDD2.n15 VSUBS 0.030259f
C994 VDD2.n16 VSUBS 0.01626f
C995 VDD2.n17 VSUBS 0.038432f
C996 VDD2.n18 VSUBS 0.017216f
C997 VDD2.n19 VSUBS 0.030259f
C998 VDD2.n20 VSUBS 0.01626f
C999 VDD2.n21 VSUBS 0.028824f
C1000 VDD2.n22 VSUBS 0.024449f
C1001 VDD2.t4 VSUBS 0.082096f
C1002 VDD2.n23 VSUBS 0.191703f
C1003 VDD2.n24 VSUBS 1.59967f
C1004 VDD2.n25 VSUBS 0.01626f
C1005 VDD2.n26 VSUBS 0.017216f
C1006 VDD2.n27 VSUBS 0.038432f
C1007 VDD2.n28 VSUBS 0.038432f
C1008 VDD2.n29 VSUBS 0.017216f
C1009 VDD2.n30 VSUBS 0.01626f
C1010 VDD2.n31 VSUBS 0.030259f
C1011 VDD2.n32 VSUBS 0.030259f
C1012 VDD2.n33 VSUBS 0.01626f
C1013 VDD2.n34 VSUBS 0.017216f
C1014 VDD2.n35 VSUBS 0.038432f
C1015 VDD2.n36 VSUBS 0.038432f
C1016 VDD2.n37 VSUBS 0.017216f
C1017 VDD2.n38 VSUBS 0.01626f
C1018 VDD2.n39 VSUBS 0.030259f
C1019 VDD2.n40 VSUBS 0.030259f
C1020 VDD2.n41 VSUBS 0.01626f
C1021 VDD2.n42 VSUBS 0.017216f
C1022 VDD2.n43 VSUBS 0.038432f
C1023 VDD2.n44 VSUBS 0.038432f
C1024 VDD2.n45 VSUBS 0.017216f
C1025 VDD2.n46 VSUBS 0.01626f
C1026 VDD2.n47 VSUBS 0.030259f
C1027 VDD2.n48 VSUBS 0.030259f
C1028 VDD2.n49 VSUBS 0.01626f
C1029 VDD2.n50 VSUBS 0.017216f
C1030 VDD2.n51 VSUBS 0.038432f
C1031 VDD2.n52 VSUBS 0.038432f
C1032 VDD2.n53 VSUBS 0.017216f
C1033 VDD2.n54 VSUBS 0.01626f
C1034 VDD2.n55 VSUBS 0.030259f
C1035 VDD2.n56 VSUBS 0.030259f
C1036 VDD2.n57 VSUBS 0.01626f
C1037 VDD2.n58 VSUBS 0.017216f
C1038 VDD2.n59 VSUBS 0.038432f
C1039 VDD2.n60 VSUBS 0.038432f
C1040 VDD2.n61 VSUBS 0.017216f
C1041 VDD2.n62 VSUBS 0.01626f
C1042 VDD2.n63 VSUBS 0.030259f
C1043 VDD2.n64 VSUBS 0.074076f
C1044 VDD2.n65 VSUBS 0.01626f
C1045 VDD2.n66 VSUBS 0.017216f
C1046 VDD2.n67 VSUBS 0.082998f
C1047 VDD2.n68 VSUBS 0.093816f
C1048 VDD2.t9 VSUBS 0.300808f
C1049 VDD2.t3 VSUBS 0.300808f
C1050 VDD2.n69 VSUBS 2.38623f
C1051 VDD2.n70 VSUBS 1.22743f
C1052 VDD2.t7 VSUBS 0.300808f
C1053 VDD2.t0 VSUBS 0.300808f
C1054 VDD2.n71 VSUBS 2.41545f
C1055 VDD2.n72 VSUBS 4.13725f
C1056 VDD2.n73 VSUBS 0.016991f
C1057 VDD2.n74 VSUBS 0.038432f
C1058 VDD2.n75 VSUBS 0.017216f
C1059 VDD2.n76 VSUBS 0.030259f
C1060 VDD2.n77 VSUBS 0.01626f
C1061 VDD2.n78 VSUBS 0.038432f
C1062 VDD2.n79 VSUBS 0.017216f
C1063 VDD2.n80 VSUBS 0.030259f
C1064 VDD2.n81 VSUBS 0.01626f
C1065 VDD2.n82 VSUBS 0.038432f
C1066 VDD2.n83 VSUBS 0.017216f
C1067 VDD2.n84 VSUBS 0.030259f
C1068 VDD2.n85 VSUBS 0.01626f
C1069 VDD2.n86 VSUBS 0.038432f
C1070 VDD2.n87 VSUBS 0.017216f
C1071 VDD2.n88 VSUBS 0.030259f
C1072 VDD2.n89 VSUBS 0.01626f
C1073 VDD2.n90 VSUBS 0.038432f
C1074 VDD2.n91 VSUBS 0.017216f
C1075 VDD2.n92 VSUBS 0.030259f
C1076 VDD2.n93 VSUBS 0.01626f
C1077 VDD2.n94 VSUBS 0.028824f
C1078 VDD2.n95 VSUBS 0.024449f
C1079 VDD2.t5 VSUBS 0.082096f
C1080 VDD2.n96 VSUBS 0.191703f
C1081 VDD2.n97 VSUBS 1.59967f
C1082 VDD2.n98 VSUBS 0.01626f
C1083 VDD2.n99 VSUBS 0.017216f
C1084 VDD2.n100 VSUBS 0.038432f
C1085 VDD2.n101 VSUBS 0.038432f
C1086 VDD2.n102 VSUBS 0.017216f
C1087 VDD2.n103 VSUBS 0.01626f
C1088 VDD2.n104 VSUBS 0.030259f
C1089 VDD2.n105 VSUBS 0.030259f
C1090 VDD2.n106 VSUBS 0.01626f
C1091 VDD2.n107 VSUBS 0.017216f
C1092 VDD2.n108 VSUBS 0.038432f
C1093 VDD2.n109 VSUBS 0.038432f
C1094 VDD2.n110 VSUBS 0.017216f
C1095 VDD2.n111 VSUBS 0.01626f
C1096 VDD2.n112 VSUBS 0.030259f
C1097 VDD2.n113 VSUBS 0.030259f
C1098 VDD2.n114 VSUBS 0.01626f
C1099 VDD2.n115 VSUBS 0.017216f
C1100 VDD2.n116 VSUBS 0.038432f
C1101 VDD2.n117 VSUBS 0.038432f
C1102 VDD2.n118 VSUBS 0.017216f
C1103 VDD2.n119 VSUBS 0.01626f
C1104 VDD2.n120 VSUBS 0.030259f
C1105 VDD2.n121 VSUBS 0.030259f
C1106 VDD2.n122 VSUBS 0.01626f
C1107 VDD2.n123 VSUBS 0.017216f
C1108 VDD2.n124 VSUBS 0.038432f
C1109 VDD2.n125 VSUBS 0.038432f
C1110 VDD2.n126 VSUBS 0.017216f
C1111 VDD2.n127 VSUBS 0.01626f
C1112 VDD2.n128 VSUBS 0.030259f
C1113 VDD2.n129 VSUBS 0.030259f
C1114 VDD2.n130 VSUBS 0.01626f
C1115 VDD2.n131 VSUBS 0.017216f
C1116 VDD2.n132 VSUBS 0.038432f
C1117 VDD2.n133 VSUBS 0.038432f
C1118 VDD2.n134 VSUBS 0.017216f
C1119 VDD2.n135 VSUBS 0.01626f
C1120 VDD2.n136 VSUBS 0.030259f
C1121 VDD2.n137 VSUBS 0.074076f
C1122 VDD2.n138 VSUBS 0.01626f
C1123 VDD2.n139 VSUBS 0.017216f
C1124 VDD2.n140 VSUBS 0.082998f
C1125 VDD2.n141 VSUBS 0.075105f
C1126 VDD2.n142 VSUBS 3.76147f
C1127 VDD2.t8 VSUBS 0.300808f
C1128 VDD2.t1 VSUBS 0.300808f
C1129 VDD2.n143 VSUBS 2.38623f
C1130 VDD2.n144 VSUBS 0.912751f
C1131 VDD2.t2 VSUBS 0.300808f
C1132 VDD2.t6 VSUBS 0.300808f
C1133 VDD2.n145 VSUBS 2.41539f
C1134 VN.t9 VSUBS 2.67438f
C1135 VN.n0 VSUBS 1.04848f
C1136 VN.n1 VSUBS 0.025632f
C1137 VN.n2 VSUBS 0.041161f
C1138 VN.n3 VSUBS 0.025632f
C1139 VN.t2 VSUBS 2.67438f
C1140 VN.n4 VSUBS 0.047533f
C1141 VN.n5 VSUBS 0.025632f
C1142 VN.n6 VSUBS 0.047533f
C1143 VN.n7 VSUBS 0.025632f
C1144 VN.t6 VSUBS 2.67438f
C1145 VN.n8 VSUBS 0.048425f
C1146 VN.n9 VSUBS 0.025632f
C1147 VN.n10 VSUBS 0.029699f
C1148 VN.t0 VSUBS 2.67438f
C1149 VN.n11 VSUBS 1.01513f
C1150 VN.t5 VSUBS 2.94445f
C1151 VN.n12 VSUBS 0.984137f
C1152 VN.n13 VSUBS 0.276148f
C1153 VN.n14 VSUBS 0.025632f
C1154 VN.n15 VSUBS 0.047533f
C1155 VN.n16 VSUBS 0.051512f
C1156 VN.n17 VSUBS 0.022117f
C1157 VN.n18 VSUBS 0.025632f
C1158 VN.n19 VSUBS 0.025632f
C1159 VN.n20 VSUBS 0.025632f
C1160 VN.n21 VSUBS 0.047533f
C1161 VN.n22 VSUBS 0.0358f
C1162 VN.n23 VSUBS 0.93919f
C1163 VN.n24 VSUBS 0.0358f
C1164 VN.n25 VSUBS 0.025632f
C1165 VN.n26 VSUBS 0.025632f
C1166 VN.n27 VSUBS 0.025632f
C1167 VN.n28 VSUBS 0.048425f
C1168 VN.n29 VSUBS 0.022117f
C1169 VN.n30 VSUBS 0.051512f
C1170 VN.n31 VSUBS 0.025632f
C1171 VN.n32 VSUBS 0.025632f
C1172 VN.n33 VSUBS 0.025632f
C1173 VN.n34 VSUBS 0.029699f
C1174 VN.n35 VSUBS 0.93919f
C1175 VN.n36 VSUBS 0.041901f
C1176 VN.n37 VSUBS 0.047533f
C1177 VN.n38 VSUBS 0.025632f
C1178 VN.n39 VSUBS 0.025632f
C1179 VN.n40 VSUBS 0.025632f
C1180 VN.n41 VSUBS 0.03336f
C1181 VN.n42 VSUBS 0.047533f
C1182 VN.n43 VSUBS 0.047064f
C1183 VN.n44 VSUBS 0.041364f
C1184 VN.n45 VSUBS 0.048535f
C1185 VN.t4 VSUBS 2.67438f
C1186 VN.n46 VSUBS 1.04848f
C1187 VN.n47 VSUBS 0.025632f
C1188 VN.n48 VSUBS 0.041161f
C1189 VN.n49 VSUBS 0.025632f
C1190 VN.t1 VSUBS 2.67438f
C1191 VN.n50 VSUBS 0.047533f
C1192 VN.n51 VSUBS 0.025632f
C1193 VN.n52 VSUBS 0.047533f
C1194 VN.n53 VSUBS 0.025632f
C1195 VN.t8 VSUBS 2.67438f
C1196 VN.n54 VSUBS 0.048425f
C1197 VN.n55 VSUBS 0.025632f
C1198 VN.n56 VSUBS 0.029699f
C1199 VN.t3 VSUBS 2.94445f
C1200 VN.t7 VSUBS 2.67438f
C1201 VN.n57 VSUBS 1.01513f
C1202 VN.n58 VSUBS 0.984137f
C1203 VN.n59 VSUBS 0.276148f
C1204 VN.n60 VSUBS 0.025632f
C1205 VN.n61 VSUBS 0.047533f
C1206 VN.n62 VSUBS 0.051512f
C1207 VN.n63 VSUBS 0.022117f
C1208 VN.n64 VSUBS 0.025632f
C1209 VN.n65 VSUBS 0.025632f
C1210 VN.n66 VSUBS 0.025632f
C1211 VN.n67 VSUBS 0.047533f
C1212 VN.n68 VSUBS 0.0358f
C1213 VN.n69 VSUBS 0.93919f
C1214 VN.n70 VSUBS 0.0358f
C1215 VN.n71 VSUBS 0.025632f
C1216 VN.n72 VSUBS 0.025632f
C1217 VN.n73 VSUBS 0.025632f
C1218 VN.n74 VSUBS 0.048425f
C1219 VN.n75 VSUBS 0.022117f
C1220 VN.n76 VSUBS 0.051512f
C1221 VN.n77 VSUBS 0.025632f
C1222 VN.n78 VSUBS 0.025632f
C1223 VN.n79 VSUBS 0.025632f
C1224 VN.n80 VSUBS 0.029699f
C1225 VN.n81 VSUBS 0.93919f
C1226 VN.n82 VSUBS 0.041901f
C1227 VN.n83 VSUBS 0.047533f
C1228 VN.n84 VSUBS 0.025632f
C1229 VN.n85 VSUBS 0.025632f
C1230 VN.n86 VSUBS 0.025632f
C1231 VN.n87 VSUBS 0.03336f
C1232 VN.n88 VSUBS 0.047533f
C1233 VN.n89 VSUBS 0.047064f
C1234 VN.n90 VSUBS 0.041364f
C1235 VN.n91 VSUBS 1.71305f
C1236 VTAIL.t4 VSUBS 0.289328f
C1237 VTAIL.t1 VSUBS 0.289328f
C1238 VTAIL.n0 VSUBS 2.14357f
C1239 VTAIL.n1 VSUBS 1.034f
C1240 VTAIL.n2 VSUBS 0.016343f
C1241 VTAIL.n3 VSUBS 0.036966f
C1242 VTAIL.n4 VSUBS 0.016559f
C1243 VTAIL.n5 VSUBS 0.029104f
C1244 VTAIL.n6 VSUBS 0.015639f
C1245 VTAIL.n7 VSUBS 0.036966f
C1246 VTAIL.n8 VSUBS 0.016559f
C1247 VTAIL.n9 VSUBS 0.029104f
C1248 VTAIL.n10 VSUBS 0.015639f
C1249 VTAIL.n11 VSUBS 0.036966f
C1250 VTAIL.n12 VSUBS 0.016559f
C1251 VTAIL.n13 VSUBS 0.029104f
C1252 VTAIL.n14 VSUBS 0.015639f
C1253 VTAIL.n15 VSUBS 0.036966f
C1254 VTAIL.n16 VSUBS 0.016559f
C1255 VTAIL.n17 VSUBS 0.029104f
C1256 VTAIL.n18 VSUBS 0.015639f
C1257 VTAIL.n19 VSUBS 0.036966f
C1258 VTAIL.n20 VSUBS 0.016559f
C1259 VTAIL.n21 VSUBS 0.029104f
C1260 VTAIL.n22 VSUBS 0.015639f
C1261 VTAIL.n23 VSUBS 0.027724f
C1262 VTAIL.n24 VSUBS 0.023516f
C1263 VTAIL.t16 VSUBS 0.078963f
C1264 VTAIL.n25 VSUBS 0.184387f
C1265 VTAIL.n26 VSUBS 1.53862f
C1266 VTAIL.n27 VSUBS 0.015639f
C1267 VTAIL.n28 VSUBS 0.016559f
C1268 VTAIL.n29 VSUBS 0.036966f
C1269 VTAIL.n30 VSUBS 0.036966f
C1270 VTAIL.n31 VSUBS 0.016559f
C1271 VTAIL.n32 VSUBS 0.015639f
C1272 VTAIL.n33 VSUBS 0.029104f
C1273 VTAIL.n34 VSUBS 0.029104f
C1274 VTAIL.n35 VSUBS 0.015639f
C1275 VTAIL.n36 VSUBS 0.016559f
C1276 VTAIL.n37 VSUBS 0.036966f
C1277 VTAIL.n38 VSUBS 0.036966f
C1278 VTAIL.n39 VSUBS 0.016559f
C1279 VTAIL.n40 VSUBS 0.015639f
C1280 VTAIL.n41 VSUBS 0.029104f
C1281 VTAIL.n42 VSUBS 0.029104f
C1282 VTAIL.n43 VSUBS 0.015639f
C1283 VTAIL.n44 VSUBS 0.016559f
C1284 VTAIL.n45 VSUBS 0.036966f
C1285 VTAIL.n46 VSUBS 0.036966f
C1286 VTAIL.n47 VSUBS 0.016559f
C1287 VTAIL.n48 VSUBS 0.015639f
C1288 VTAIL.n49 VSUBS 0.029104f
C1289 VTAIL.n50 VSUBS 0.029104f
C1290 VTAIL.n51 VSUBS 0.015639f
C1291 VTAIL.n52 VSUBS 0.016559f
C1292 VTAIL.n53 VSUBS 0.036966f
C1293 VTAIL.n54 VSUBS 0.036966f
C1294 VTAIL.n55 VSUBS 0.016559f
C1295 VTAIL.n56 VSUBS 0.015639f
C1296 VTAIL.n57 VSUBS 0.029104f
C1297 VTAIL.n58 VSUBS 0.029104f
C1298 VTAIL.n59 VSUBS 0.015639f
C1299 VTAIL.n60 VSUBS 0.016559f
C1300 VTAIL.n61 VSUBS 0.036966f
C1301 VTAIL.n62 VSUBS 0.036966f
C1302 VTAIL.n63 VSUBS 0.016559f
C1303 VTAIL.n64 VSUBS 0.015639f
C1304 VTAIL.n65 VSUBS 0.029104f
C1305 VTAIL.n66 VSUBS 0.071249f
C1306 VTAIL.n67 VSUBS 0.015639f
C1307 VTAIL.n68 VSUBS 0.016559f
C1308 VTAIL.n69 VSUBS 0.07983f
C1309 VTAIL.n70 VSUBS 0.052167f
C1310 VTAIL.n71 VSUBS 0.479387f
C1311 VTAIL.t15 VSUBS 0.289328f
C1312 VTAIL.t18 VSUBS 0.289328f
C1313 VTAIL.n72 VSUBS 2.14357f
C1314 VTAIL.n73 VSUBS 1.18882f
C1315 VTAIL.t11 VSUBS 0.289328f
C1316 VTAIL.t9 VSUBS 0.289328f
C1317 VTAIL.n74 VSUBS 2.14357f
C1318 VTAIL.n75 VSUBS 2.87365f
C1319 VTAIL.t19 VSUBS 0.289328f
C1320 VTAIL.t5 VSUBS 0.289328f
C1321 VTAIL.n76 VSUBS 2.14357f
C1322 VTAIL.n77 VSUBS 2.87364f
C1323 VTAIL.t6 VSUBS 0.289328f
C1324 VTAIL.t3 VSUBS 0.289328f
C1325 VTAIL.n78 VSUBS 2.14357f
C1326 VTAIL.n79 VSUBS 1.18882f
C1327 VTAIL.n80 VSUBS 0.016343f
C1328 VTAIL.n81 VSUBS 0.036966f
C1329 VTAIL.n82 VSUBS 0.016559f
C1330 VTAIL.n83 VSUBS 0.029104f
C1331 VTAIL.n84 VSUBS 0.015639f
C1332 VTAIL.n85 VSUBS 0.036966f
C1333 VTAIL.n86 VSUBS 0.016559f
C1334 VTAIL.n87 VSUBS 0.029104f
C1335 VTAIL.n88 VSUBS 0.015639f
C1336 VTAIL.n89 VSUBS 0.036966f
C1337 VTAIL.n90 VSUBS 0.016559f
C1338 VTAIL.n91 VSUBS 0.029104f
C1339 VTAIL.n92 VSUBS 0.015639f
C1340 VTAIL.n93 VSUBS 0.036966f
C1341 VTAIL.n94 VSUBS 0.016559f
C1342 VTAIL.n95 VSUBS 0.029104f
C1343 VTAIL.n96 VSUBS 0.015639f
C1344 VTAIL.n97 VSUBS 0.036966f
C1345 VTAIL.n98 VSUBS 0.016559f
C1346 VTAIL.n99 VSUBS 0.029104f
C1347 VTAIL.n100 VSUBS 0.015639f
C1348 VTAIL.n101 VSUBS 0.027724f
C1349 VTAIL.n102 VSUBS 0.023516f
C1350 VTAIL.t7 VSUBS 0.078963f
C1351 VTAIL.n103 VSUBS 0.184387f
C1352 VTAIL.n104 VSUBS 1.53862f
C1353 VTAIL.n105 VSUBS 0.015639f
C1354 VTAIL.n106 VSUBS 0.016559f
C1355 VTAIL.n107 VSUBS 0.036966f
C1356 VTAIL.n108 VSUBS 0.036966f
C1357 VTAIL.n109 VSUBS 0.016559f
C1358 VTAIL.n110 VSUBS 0.015639f
C1359 VTAIL.n111 VSUBS 0.029104f
C1360 VTAIL.n112 VSUBS 0.029104f
C1361 VTAIL.n113 VSUBS 0.015639f
C1362 VTAIL.n114 VSUBS 0.016559f
C1363 VTAIL.n115 VSUBS 0.036966f
C1364 VTAIL.n116 VSUBS 0.036966f
C1365 VTAIL.n117 VSUBS 0.016559f
C1366 VTAIL.n118 VSUBS 0.015639f
C1367 VTAIL.n119 VSUBS 0.029104f
C1368 VTAIL.n120 VSUBS 0.029104f
C1369 VTAIL.n121 VSUBS 0.015639f
C1370 VTAIL.n122 VSUBS 0.016559f
C1371 VTAIL.n123 VSUBS 0.036966f
C1372 VTAIL.n124 VSUBS 0.036966f
C1373 VTAIL.n125 VSUBS 0.016559f
C1374 VTAIL.n126 VSUBS 0.015639f
C1375 VTAIL.n127 VSUBS 0.029104f
C1376 VTAIL.n128 VSUBS 0.029104f
C1377 VTAIL.n129 VSUBS 0.015639f
C1378 VTAIL.n130 VSUBS 0.016559f
C1379 VTAIL.n131 VSUBS 0.036966f
C1380 VTAIL.n132 VSUBS 0.036966f
C1381 VTAIL.n133 VSUBS 0.016559f
C1382 VTAIL.n134 VSUBS 0.015639f
C1383 VTAIL.n135 VSUBS 0.029104f
C1384 VTAIL.n136 VSUBS 0.029104f
C1385 VTAIL.n137 VSUBS 0.015639f
C1386 VTAIL.n138 VSUBS 0.016559f
C1387 VTAIL.n139 VSUBS 0.036966f
C1388 VTAIL.n140 VSUBS 0.036966f
C1389 VTAIL.n141 VSUBS 0.016559f
C1390 VTAIL.n142 VSUBS 0.015639f
C1391 VTAIL.n143 VSUBS 0.029104f
C1392 VTAIL.n144 VSUBS 0.071249f
C1393 VTAIL.n145 VSUBS 0.015639f
C1394 VTAIL.n146 VSUBS 0.016559f
C1395 VTAIL.n147 VSUBS 0.07983f
C1396 VTAIL.n148 VSUBS 0.052167f
C1397 VTAIL.n149 VSUBS 0.479387f
C1398 VTAIL.t10 VSUBS 0.289328f
C1399 VTAIL.t14 VSUBS 0.289328f
C1400 VTAIL.n150 VSUBS 2.14357f
C1401 VTAIL.n151 VSUBS 1.09665f
C1402 VTAIL.t17 VSUBS 0.289328f
C1403 VTAIL.t13 VSUBS 0.289328f
C1404 VTAIL.n152 VSUBS 2.14357f
C1405 VTAIL.n153 VSUBS 1.18882f
C1406 VTAIL.n154 VSUBS 0.016343f
C1407 VTAIL.n155 VSUBS 0.036966f
C1408 VTAIL.n156 VSUBS 0.016559f
C1409 VTAIL.n157 VSUBS 0.029104f
C1410 VTAIL.n158 VSUBS 0.015639f
C1411 VTAIL.n159 VSUBS 0.036966f
C1412 VTAIL.n160 VSUBS 0.016559f
C1413 VTAIL.n161 VSUBS 0.029104f
C1414 VTAIL.n162 VSUBS 0.015639f
C1415 VTAIL.n163 VSUBS 0.036966f
C1416 VTAIL.n164 VSUBS 0.016559f
C1417 VTAIL.n165 VSUBS 0.029104f
C1418 VTAIL.n166 VSUBS 0.015639f
C1419 VTAIL.n167 VSUBS 0.036966f
C1420 VTAIL.n168 VSUBS 0.016559f
C1421 VTAIL.n169 VSUBS 0.029104f
C1422 VTAIL.n170 VSUBS 0.015639f
C1423 VTAIL.n171 VSUBS 0.036966f
C1424 VTAIL.n172 VSUBS 0.016559f
C1425 VTAIL.n173 VSUBS 0.029104f
C1426 VTAIL.n174 VSUBS 0.015639f
C1427 VTAIL.n175 VSUBS 0.027724f
C1428 VTAIL.n176 VSUBS 0.023516f
C1429 VTAIL.t12 VSUBS 0.078963f
C1430 VTAIL.n177 VSUBS 0.184387f
C1431 VTAIL.n178 VSUBS 1.53862f
C1432 VTAIL.n179 VSUBS 0.015639f
C1433 VTAIL.n180 VSUBS 0.016559f
C1434 VTAIL.n181 VSUBS 0.036966f
C1435 VTAIL.n182 VSUBS 0.036966f
C1436 VTAIL.n183 VSUBS 0.016559f
C1437 VTAIL.n184 VSUBS 0.015639f
C1438 VTAIL.n185 VSUBS 0.029104f
C1439 VTAIL.n186 VSUBS 0.029104f
C1440 VTAIL.n187 VSUBS 0.015639f
C1441 VTAIL.n188 VSUBS 0.016559f
C1442 VTAIL.n189 VSUBS 0.036966f
C1443 VTAIL.n190 VSUBS 0.036966f
C1444 VTAIL.n191 VSUBS 0.016559f
C1445 VTAIL.n192 VSUBS 0.015639f
C1446 VTAIL.n193 VSUBS 0.029104f
C1447 VTAIL.n194 VSUBS 0.029104f
C1448 VTAIL.n195 VSUBS 0.015639f
C1449 VTAIL.n196 VSUBS 0.016559f
C1450 VTAIL.n197 VSUBS 0.036966f
C1451 VTAIL.n198 VSUBS 0.036966f
C1452 VTAIL.n199 VSUBS 0.016559f
C1453 VTAIL.n200 VSUBS 0.015639f
C1454 VTAIL.n201 VSUBS 0.029104f
C1455 VTAIL.n202 VSUBS 0.029104f
C1456 VTAIL.n203 VSUBS 0.015639f
C1457 VTAIL.n204 VSUBS 0.016559f
C1458 VTAIL.n205 VSUBS 0.036966f
C1459 VTAIL.n206 VSUBS 0.036966f
C1460 VTAIL.n207 VSUBS 0.016559f
C1461 VTAIL.n208 VSUBS 0.015639f
C1462 VTAIL.n209 VSUBS 0.029104f
C1463 VTAIL.n210 VSUBS 0.029104f
C1464 VTAIL.n211 VSUBS 0.015639f
C1465 VTAIL.n212 VSUBS 0.016559f
C1466 VTAIL.n213 VSUBS 0.036966f
C1467 VTAIL.n214 VSUBS 0.036966f
C1468 VTAIL.n215 VSUBS 0.016559f
C1469 VTAIL.n216 VSUBS 0.015639f
C1470 VTAIL.n217 VSUBS 0.029104f
C1471 VTAIL.n218 VSUBS 0.071249f
C1472 VTAIL.n219 VSUBS 0.015639f
C1473 VTAIL.n220 VSUBS 0.016559f
C1474 VTAIL.n221 VSUBS 0.07983f
C1475 VTAIL.n222 VSUBS 0.052167f
C1476 VTAIL.n223 VSUBS 1.98393f
C1477 VTAIL.n224 VSUBS 0.016343f
C1478 VTAIL.n225 VSUBS 0.036966f
C1479 VTAIL.n226 VSUBS 0.016559f
C1480 VTAIL.n227 VSUBS 0.029104f
C1481 VTAIL.n228 VSUBS 0.015639f
C1482 VTAIL.n229 VSUBS 0.036966f
C1483 VTAIL.n230 VSUBS 0.016559f
C1484 VTAIL.n231 VSUBS 0.029104f
C1485 VTAIL.n232 VSUBS 0.015639f
C1486 VTAIL.n233 VSUBS 0.036966f
C1487 VTAIL.n234 VSUBS 0.016559f
C1488 VTAIL.n235 VSUBS 0.029104f
C1489 VTAIL.n236 VSUBS 0.015639f
C1490 VTAIL.n237 VSUBS 0.036966f
C1491 VTAIL.n238 VSUBS 0.016559f
C1492 VTAIL.n239 VSUBS 0.029104f
C1493 VTAIL.n240 VSUBS 0.015639f
C1494 VTAIL.n241 VSUBS 0.036966f
C1495 VTAIL.n242 VSUBS 0.016559f
C1496 VTAIL.n243 VSUBS 0.029104f
C1497 VTAIL.n244 VSUBS 0.015639f
C1498 VTAIL.n245 VSUBS 0.027724f
C1499 VTAIL.n246 VSUBS 0.023516f
C1500 VTAIL.t8 VSUBS 0.078963f
C1501 VTAIL.n247 VSUBS 0.184387f
C1502 VTAIL.n248 VSUBS 1.53862f
C1503 VTAIL.n249 VSUBS 0.015639f
C1504 VTAIL.n250 VSUBS 0.016559f
C1505 VTAIL.n251 VSUBS 0.036966f
C1506 VTAIL.n252 VSUBS 0.036966f
C1507 VTAIL.n253 VSUBS 0.016559f
C1508 VTAIL.n254 VSUBS 0.015639f
C1509 VTAIL.n255 VSUBS 0.029104f
C1510 VTAIL.n256 VSUBS 0.029104f
C1511 VTAIL.n257 VSUBS 0.015639f
C1512 VTAIL.n258 VSUBS 0.016559f
C1513 VTAIL.n259 VSUBS 0.036966f
C1514 VTAIL.n260 VSUBS 0.036966f
C1515 VTAIL.n261 VSUBS 0.016559f
C1516 VTAIL.n262 VSUBS 0.015639f
C1517 VTAIL.n263 VSUBS 0.029104f
C1518 VTAIL.n264 VSUBS 0.029104f
C1519 VTAIL.n265 VSUBS 0.015639f
C1520 VTAIL.n266 VSUBS 0.016559f
C1521 VTAIL.n267 VSUBS 0.036966f
C1522 VTAIL.n268 VSUBS 0.036966f
C1523 VTAIL.n269 VSUBS 0.016559f
C1524 VTAIL.n270 VSUBS 0.015639f
C1525 VTAIL.n271 VSUBS 0.029104f
C1526 VTAIL.n272 VSUBS 0.029104f
C1527 VTAIL.n273 VSUBS 0.015639f
C1528 VTAIL.n274 VSUBS 0.016559f
C1529 VTAIL.n275 VSUBS 0.036966f
C1530 VTAIL.n276 VSUBS 0.036966f
C1531 VTAIL.n277 VSUBS 0.016559f
C1532 VTAIL.n278 VSUBS 0.015639f
C1533 VTAIL.n279 VSUBS 0.029104f
C1534 VTAIL.n280 VSUBS 0.029104f
C1535 VTAIL.n281 VSUBS 0.015639f
C1536 VTAIL.n282 VSUBS 0.016559f
C1537 VTAIL.n283 VSUBS 0.036966f
C1538 VTAIL.n284 VSUBS 0.036966f
C1539 VTAIL.n285 VSUBS 0.016559f
C1540 VTAIL.n286 VSUBS 0.015639f
C1541 VTAIL.n287 VSUBS 0.029104f
C1542 VTAIL.n288 VSUBS 0.071249f
C1543 VTAIL.n289 VSUBS 0.015639f
C1544 VTAIL.n290 VSUBS 0.016559f
C1545 VTAIL.n291 VSUBS 0.07983f
C1546 VTAIL.n292 VSUBS 0.052167f
C1547 VTAIL.n293 VSUBS 1.98393f
C1548 VTAIL.t0 VSUBS 0.289328f
C1549 VTAIL.t2 VSUBS 0.289328f
C1550 VTAIL.n294 VSUBS 2.14357f
C1551 VTAIL.n295 VSUBS 0.979028f
C1552 VDD1.n0 VSUBS 0.017039f
C1553 VDD1.n1 VSUBS 0.038542f
C1554 VDD1.n2 VSUBS 0.017265f
C1555 VDD1.n3 VSUBS 0.030346f
C1556 VDD1.n4 VSUBS 0.016306f
C1557 VDD1.n5 VSUBS 0.038542f
C1558 VDD1.n6 VSUBS 0.017265f
C1559 VDD1.n7 VSUBS 0.030346f
C1560 VDD1.n8 VSUBS 0.016306f
C1561 VDD1.n9 VSUBS 0.038542f
C1562 VDD1.n10 VSUBS 0.017265f
C1563 VDD1.n11 VSUBS 0.030346f
C1564 VDD1.n12 VSUBS 0.016306f
C1565 VDD1.n13 VSUBS 0.038542f
C1566 VDD1.n14 VSUBS 0.017265f
C1567 VDD1.n15 VSUBS 0.030346f
C1568 VDD1.n16 VSUBS 0.016306f
C1569 VDD1.n17 VSUBS 0.038542f
C1570 VDD1.n18 VSUBS 0.017265f
C1571 VDD1.n19 VSUBS 0.030346f
C1572 VDD1.n20 VSUBS 0.016306f
C1573 VDD1.n21 VSUBS 0.028907f
C1574 VDD1.n22 VSUBS 0.024519f
C1575 VDD1.t3 VSUBS 0.082331f
C1576 VDD1.n23 VSUBS 0.192251f
C1577 VDD1.n24 VSUBS 1.60424f
C1578 VDD1.n25 VSUBS 0.016306f
C1579 VDD1.n26 VSUBS 0.017265f
C1580 VDD1.n27 VSUBS 0.038542f
C1581 VDD1.n28 VSUBS 0.038542f
C1582 VDD1.n29 VSUBS 0.017265f
C1583 VDD1.n30 VSUBS 0.016306f
C1584 VDD1.n31 VSUBS 0.030346f
C1585 VDD1.n32 VSUBS 0.030346f
C1586 VDD1.n33 VSUBS 0.016306f
C1587 VDD1.n34 VSUBS 0.017265f
C1588 VDD1.n35 VSUBS 0.038542f
C1589 VDD1.n36 VSUBS 0.038542f
C1590 VDD1.n37 VSUBS 0.017265f
C1591 VDD1.n38 VSUBS 0.016306f
C1592 VDD1.n39 VSUBS 0.030346f
C1593 VDD1.n40 VSUBS 0.030346f
C1594 VDD1.n41 VSUBS 0.016306f
C1595 VDD1.n42 VSUBS 0.017265f
C1596 VDD1.n43 VSUBS 0.038542f
C1597 VDD1.n44 VSUBS 0.038542f
C1598 VDD1.n45 VSUBS 0.017265f
C1599 VDD1.n46 VSUBS 0.016306f
C1600 VDD1.n47 VSUBS 0.030346f
C1601 VDD1.n48 VSUBS 0.030346f
C1602 VDD1.n49 VSUBS 0.016306f
C1603 VDD1.n50 VSUBS 0.017265f
C1604 VDD1.n51 VSUBS 0.038542f
C1605 VDD1.n52 VSUBS 0.038542f
C1606 VDD1.n53 VSUBS 0.017265f
C1607 VDD1.n54 VSUBS 0.016306f
C1608 VDD1.n55 VSUBS 0.030346f
C1609 VDD1.n56 VSUBS 0.030346f
C1610 VDD1.n57 VSUBS 0.016306f
C1611 VDD1.n58 VSUBS 0.017265f
C1612 VDD1.n59 VSUBS 0.038542f
C1613 VDD1.n60 VSUBS 0.038542f
C1614 VDD1.n61 VSUBS 0.017265f
C1615 VDD1.n62 VSUBS 0.016306f
C1616 VDD1.n63 VSUBS 0.030346f
C1617 VDD1.n64 VSUBS 0.074288f
C1618 VDD1.n65 VSUBS 0.016306f
C1619 VDD1.n66 VSUBS 0.017265f
C1620 VDD1.n67 VSUBS 0.083235f
C1621 VDD1.n68 VSUBS 0.094084f
C1622 VDD1.t5 VSUBS 0.301667f
C1623 VDD1.t1 VSUBS 0.301667f
C1624 VDD1.n69 VSUBS 2.39304f
C1625 VDD1.n70 VSUBS 1.24099f
C1626 VDD1.n71 VSUBS 0.017039f
C1627 VDD1.n72 VSUBS 0.038542f
C1628 VDD1.n73 VSUBS 0.017265f
C1629 VDD1.n74 VSUBS 0.030346f
C1630 VDD1.n75 VSUBS 0.016306f
C1631 VDD1.n76 VSUBS 0.038542f
C1632 VDD1.n77 VSUBS 0.017265f
C1633 VDD1.n78 VSUBS 0.030346f
C1634 VDD1.n79 VSUBS 0.016306f
C1635 VDD1.n80 VSUBS 0.038542f
C1636 VDD1.n81 VSUBS 0.017265f
C1637 VDD1.n82 VSUBS 0.030346f
C1638 VDD1.n83 VSUBS 0.016306f
C1639 VDD1.n84 VSUBS 0.038542f
C1640 VDD1.n85 VSUBS 0.017265f
C1641 VDD1.n86 VSUBS 0.030346f
C1642 VDD1.n87 VSUBS 0.016306f
C1643 VDD1.n88 VSUBS 0.038542f
C1644 VDD1.n89 VSUBS 0.017265f
C1645 VDD1.n90 VSUBS 0.030346f
C1646 VDD1.n91 VSUBS 0.016306f
C1647 VDD1.n92 VSUBS 0.028907f
C1648 VDD1.n93 VSUBS 0.024519f
C1649 VDD1.t4 VSUBS 0.082331f
C1650 VDD1.n94 VSUBS 0.192251f
C1651 VDD1.n95 VSUBS 1.60424f
C1652 VDD1.n96 VSUBS 0.016306f
C1653 VDD1.n97 VSUBS 0.017265f
C1654 VDD1.n98 VSUBS 0.038542f
C1655 VDD1.n99 VSUBS 0.038542f
C1656 VDD1.n100 VSUBS 0.017265f
C1657 VDD1.n101 VSUBS 0.016306f
C1658 VDD1.n102 VSUBS 0.030346f
C1659 VDD1.n103 VSUBS 0.030346f
C1660 VDD1.n104 VSUBS 0.016306f
C1661 VDD1.n105 VSUBS 0.017265f
C1662 VDD1.n106 VSUBS 0.038542f
C1663 VDD1.n107 VSUBS 0.038542f
C1664 VDD1.n108 VSUBS 0.017265f
C1665 VDD1.n109 VSUBS 0.016306f
C1666 VDD1.n110 VSUBS 0.030346f
C1667 VDD1.n111 VSUBS 0.030346f
C1668 VDD1.n112 VSUBS 0.016306f
C1669 VDD1.n113 VSUBS 0.017265f
C1670 VDD1.n114 VSUBS 0.038542f
C1671 VDD1.n115 VSUBS 0.038542f
C1672 VDD1.n116 VSUBS 0.017265f
C1673 VDD1.n117 VSUBS 0.016306f
C1674 VDD1.n118 VSUBS 0.030346f
C1675 VDD1.n119 VSUBS 0.030346f
C1676 VDD1.n120 VSUBS 0.016306f
C1677 VDD1.n121 VSUBS 0.017265f
C1678 VDD1.n122 VSUBS 0.038542f
C1679 VDD1.n123 VSUBS 0.038542f
C1680 VDD1.n124 VSUBS 0.017265f
C1681 VDD1.n125 VSUBS 0.016306f
C1682 VDD1.n126 VSUBS 0.030346f
C1683 VDD1.n127 VSUBS 0.030346f
C1684 VDD1.n128 VSUBS 0.016306f
C1685 VDD1.n129 VSUBS 0.017265f
C1686 VDD1.n130 VSUBS 0.038542f
C1687 VDD1.n131 VSUBS 0.038542f
C1688 VDD1.n132 VSUBS 0.017265f
C1689 VDD1.n133 VSUBS 0.016306f
C1690 VDD1.n134 VSUBS 0.030346f
C1691 VDD1.n135 VSUBS 0.074288f
C1692 VDD1.n136 VSUBS 0.016306f
C1693 VDD1.n137 VSUBS 0.017265f
C1694 VDD1.n138 VSUBS 0.083235f
C1695 VDD1.n139 VSUBS 0.094084f
C1696 VDD1.t2 VSUBS 0.301667f
C1697 VDD1.t6 VSUBS 0.301667f
C1698 VDD1.n140 VSUBS 2.39304f
C1699 VDD1.n141 VSUBS 1.23094f
C1700 VDD1.t7 VSUBS 0.301667f
C1701 VDD1.t0 VSUBS 0.301667f
C1702 VDD1.n142 VSUBS 2.42235f
C1703 VDD1.n143 VSUBS 4.31589f
C1704 VDD1.t9 VSUBS 0.301667f
C1705 VDD1.t8 VSUBS 0.301667f
C1706 VDD1.n144 VSUBS 2.39303f
C1707 VDD1.n145 VSUBS 4.43131f
C1708 VP.t2 VSUBS 2.89657f
C1709 VP.n0 VSUBS 1.13559f
C1710 VP.n1 VSUBS 0.027762f
C1711 VP.n2 VSUBS 0.044581f
C1712 VP.n3 VSUBS 0.027762f
C1713 VP.t0 VSUBS 2.89657f
C1714 VP.n4 VSUBS 0.051482f
C1715 VP.n5 VSUBS 0.027762f
C1716 VP.n6 VSUBS 0.051482f
C1717 VP.n7 VSUBS 0.027762f
C1718 VP.t3 VSUBS 2.89657f
C1719 VP.n8 VSUBS 0.052449f
C1720 VP.n9 VSUBS 0.027762f
C1721 VP.n10 VSUBS 0.032166f
C1722 VP.n11 VSUBS 0.027762f
C1723 VP.n12 VSUBS 0.036132f
C1724 VP.n13 VSUBS 0.0448f
C1725 VP.t7 VSUBS 2.89657f
C1726 VP.t6 VSUBS 2.89657f
C1727 VP.n14 VSUBS 1.13559f
C1728 VP.n15 VSUBS 0.027762f
C1729 VP.n16 VSUBS 0.044581f
C1730 VP.n17 VSUBS 0.027762f
C1731 VP.t5 VSUBS 2.89657f
C1732 VP.n18 VSUBS 0.051482f
C1733 VP.n19 VSUBS 0.027762f
C1734 VP.n20 VSUBS 0.051482f
C1735 VP.n21 VSUBS 0.027762f
C1736 VP.t1 VSUBS 2.89657f
C1737 VP.n22 VSUBS 0.052449f
C1738 VP.n23 VSUBS 0.027762f
C1739 VP.n24 VSUBS 0.032166f
C1740 VP.t8 VSUBS 3.18908f
C1741 VP.t4 VSUBS 2.89657f
C1742 VP.n25 VSUBS 1.09947f
C1743 VP.n26 VSUBS 1.0659f
C1744 VP.n27 VSUBS 0.299092f
C1745 VP.n28 VSUBS 0.027762f
C1746 VP.n29 VSUBS 0.051482f
C1747 VP.n30 VSUBS 0.055792f
C1748 VP.n31 VSUBS 0.023955f
C1749 VP.n32 VSUBS 0.027762f
C1750 VP.n33 VSUBS 0.027762f
C1751 VP.n34 VSUBS 0.027762f
C1752 VP.n35 VSUBS 0.051482f
C1753 VP.n36 VSUBS 0.038775f
C1754 VP.n37 VSUBS 1.01722f
C1755 VP.n38 VSUBS 0.038775f
C1756 VP.n39 VSUBS 0.027762f
C1757 VP.n40 VSUBS 0.027762f
C1758 VP.n41 VSUBS 0.027762f
C1759 VP.n42 VSUBS 0.052449f
C1760 VP.n43 VSUBS 0.023955f
C1761 VP.n44 VSUBS 0.055792f
C1762 VP.n45 VSUBS 0.027762f
C1763 VP.n46 VSUBS 0.027762f
C1764 VP.n47 VSUBS 0.027762f
C1765 VP.n48 VSUBS 0.032166f
C1766 VP.n49 VSUBS 1.01722f
C1767 VP.n50 VSUBS 0.045383f
C1768 VP.n51 VSUBS 0.051482f
C1769 VP.n52 VSUBS 0.027762f
C1770 VP.n53 VSUBS 0.027762f
C1771 VP.n54 VSUBS 0.027762f
C1772 VP.n55 VSUBS 0.036132f
C1773 VP.n56 VSUBS 0.051482f
C1774 VP.n57 VSUBS 0.050974f
C1775 VP.n58 VSUBS 0.0448f
C1776 VP.n59 VSUBS 1.84446f
C1777 VP.n60 VSUBS 1.86228f
C1778 VP.n61 VSUBS 1.13559f
C1779 VP.n62 VSUBS 0.050974f
C1780 VP.n63 VSUBS 0.051482f
C1781 VP.n64 VSUBS 0.027762f
C1782 VP.n65 VSUBS 0.027762f
C1783 VP.n66 VSUBS 0.027762f
C1784 VP.n67 VSUBS 0.044581f
C1785 VP.n68 VSUBS 0.051482f
C1786 VP.t9 VSUBS 2.89657f
C1787 VP.n69 VSUBS 1.01722f
C1788 VP.n70 VSUBS 0.045383f
C1789 VP.n71 VSUBS 0.027762f
C1790 VP.n72 VSUBS 0.027762f
C1791 VP.n73 VSUBS 0.027762f
C1792 VP.n74 VSUBS 0.051482f
C1793 VP.n75 VSUBS 0.055792f
C1794 VP.n76 VSUBS 0.023955f
C1795 VP.n77 VSUBS 0.027762f
C1796 VP.n78 VSUBS 0.027762f
C1797 VP.n79 VSUBS 0.027762f
C1798 VP.n80 VSUBS 0.051482f
C1799 VP.n81 VSUBS 0.038775f
C1800 VP.n82 VSUBS 1.01722f
C1801 VP.n83 VSUBS 0.038775f
C1802 VP.n84 VSUBS 0.027762f
C1803 VP.n85 VSUBS 0.027762f
C1804 VP.n86 VSUBS 0.027762f
C1805 VP.n87 VSUBS 0.052449f
C1806 VP.n88 VSUBS 0.023955f
C1807 VP.n89 VSUBS 0.055792f
C1808 VP.n90 VSUBS 0.027762f
C1809 VP.n91 VSUBS 0.027762f
C1810 VP.n92 VSUBS 0.027762f
C1811 VP.n93 VSUBS 0.032166f
C1812 VP.n94 VSUBS 1.01722f
C1813 VP.n95 VSUBS 0.045383f
C1814 VP.n96 VSUBS 0.051482f
C1815 VP.n97 VSUBS 0.027762f
C1816 VP.n98 VSUBS 0.027762f
C1817 VP.n99 VSUBS 0.027762f
C1818 VP.n100 VSUBS 0.036132f
C1819 VP.n101 VSUBS 0.051482f
C1820 VP.n102 VSUBS 0.050974f
C1821 VP.n103 VSUBS 0.0448f
C1822 VP.n104 VSUBS 0.052568f
.ends

