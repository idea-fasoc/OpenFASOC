* NGSPICE file created from diff_pair_sample_0350.ext - technology: sky130A

.subckt diff_pair_sample_0350 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0 ps=0 w=1.07 l=0.39
X1 B.t8 B.t6 B.t7 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0 ps=0 w=1.07 l=0.39
X2 B.t5 B.t3 B.t4 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0 ps=0 w=1.07 l=0.39
X3 VTAIL.t7 VN.t0 VDD2.t2 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0.17655 ps=1.4 w=1.07 l=0.39
X4 VTAIL.t3 VP.t0 VDD1.t3 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0.17655 ps=1.4 w=1.07 l=0.39
X5 VDD2.t1 VN.t1 VTAIL.t6 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.4173 ps=2.92 w=1.07 l=0.39
X6 B.t2 B.t0 B.t1 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0 ps=0 w=1.07 l=0.39
X7 VTAIL.t5 VN.t2 VDD2.t0 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0.17655 ps=1.4 w=1.07 l=0.39
X8 VTAIL.t1 VP.t1 VDD1.t2 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.4173 pd=2.92 as=0.17655 ps=1.4 w=1.07 l=0.39
X9 VDD1.t1 VP.t2 VTAIL.t2 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.4173 ps=2.92 w=1.07 l=0.39
X10 VDD2.t3 VN.t3 VTAIL.t4 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.4173 ps=2.92 w=1.07 l=0.39
X11 VDD1.t0 VP.t3 VTAIL.t0 w_n1402_n1186# sky130_fd_pr__pfet_01v8 ad=0.17655 pd=1.4 as=0.4173 ps=2.92 w=1.07 l=0.39
R0 B.n132 B.n43 585
R1 B.n131 B.n130 585
R2 B.n129 B.n44 585
R3 B.n128 B.n127 585
R4 B.n126 B.n45 585
R5 B.n125 B.n124 585
R6 B.n123 B.n46 585
R7 B.n122 B.n121 585
R8 B.n120 B.n47 585
R9 B.n119 B.n118 585
R10 B.n117 B.n116 585
R11 B.n115 B.n51 585
R12 B.n114 B.n113 585
R13 B.n112 B.n52 585
R14 B.n111 B.n110 585
R15 B.n109 B.n53 585
R16 B.n108 B.n107 585
R17 B.n106 B.n54 585
R18 B.n105 B.n104 585
R19 B.n102 B.n55 585
R20 B.n101 B.n100 585
R21 B.n99 B.n58 585
R22 B.n98 B.n97 585
R23 B.n96 B.n59 585
R24 B.n95 B.n94 585
R25 B.n93 B.n60 585
R26 B.n92 B.n91 585
R27 B.n90 B.n61 585
R28 B.n89 B.n88 585
R29 B.n134 B.n133 585
R30 B.n135 B.n42 585
R31 B.n137 B.n136 585
R32 B.n138 B.n41 585
R33 B.n140 B.n139 585
R34 B.n141 B.n40 585
R35 B.n143 B.n142 585
R36 B.n144 B.n39 585
R37 B.n146 B.n145 585
R38 B.n147 B.n38 585
R39 B.n149 B.n148 585
R40 B.n150 B.n37 585
R41 B.n152 B.n151 585
R42 B.n153 B.n36 585
R43 B.n155 B.n154 585
R44 B.n156 B.n35 585
R45 B.n158 B.n157 585
R46 B.n159 B.n34 585
R47 B.n161 B.n160 585
R48 B.n162 B.n33 585
R49 B.n164 B.n163 585
R50 B.n165 B.n32 585
R51 B.n167 B.n166 585
R52 B.n168 B.n31 585
R53 B.n170 B.n169 585
R54 B.n171 B.n30 585
R55 B.n173 B.n172 585
R56 B.n174 B.n29 585
R57 B.n176 B.n175 585
R58 B.n177 B.n28 585
R59 B.n222 B.n9 585
R60 B.n221 B.n220 585
R61 B.n219 B.n10 585
R62 B.n218 B.n217 585
R63 B.n216 B.n11 585
R64 B.n215 B.n214 585
R65 B.n213 B.n12 585
R66 B.n212 B.n211 585
R67 B.n210 B.n13 585
R68 B.n209 B.n208 585
R69 B.n207 B.n206 585
R70 B.n205 B.n17 585
R71 B.n204 B.n203 585
R72 B.n202 B.n18 585
R73 B.n201 B.n200 585
R74 B.n199 B.n19 585
R75 B.n198 B.n197 585
R76 B.n196 B.n20 585
R77 B.n195 B.n194 585
R78 B.n192 B.n21 585
R79 B.n191 B.n190 585
R80 B.n189 B.n24 585
R81 B.n188 B.n187 585
R82 B.n186 B.n25 585
R83 B.n185 B.n184 585
R84 B.n183 B.n26 585
R85 B.n182 B.n181 585
R86 B.n180 B.n27 585
R87 B.n179 B.n178 585
R88 B.n224 B.n223 585
R89 B.n225 B.n8 585
R90 B.n227 B.n226 585
R91 B.n228 B.n7 585
R92 B.n230 B.n229 585
R93 B.n231 B.n6 585
R94 B.n233 B.n232 585
R95 B.n234 B.n5 585
R96 B.n236 B.n235 585
R97 B.n237 B.n4 585
R98 B.n239 B.n238 585
R99 B.n240 B.n3 585
R100 B.n242 B.n241 585
R101 B.n243 B.n0 585
R102 B.n2 B.n1 585
R103 B.n69 B.n68 585
R104 B.n71 B.n70 585
R105 B.n72 B.n67 585
R106 B.n74 B.n73 585
R107 B.n75 B.n66 585
R108 B.n77 B.n76 585
R109 B.n78 B.n65 585
R110 B.n80 B.n79 585
R111 B.n81 B.n64 585
R112 B.n83 B.n82 585
R113 B.n84 B.n63 585
R114 B.n86 B.n85 585
R115 B.n87 B.n62 585
R116 B.n88 B.n87 463.671
R117 B.n134 B.n43 463.671
R118 B.n178 B.n177 463.671
R119 B.n224 B.n9 463.671
R120 B.n56 B.t4 376.521
R121 B.n48 B.t7 376.521
R122 B.n22 B.t11 376.521
R123 B.n14 B.t2 376.521
R124 B.n57 B.t5 362.557
R125 B.n49 B.t8 362.557
R126 B.n23 B.t10 362.557
R127 B.n15 B.t1 362.557
R128 B.n56 B.t3 275.928
R129 B.n48 B.t6 275.928
R130 B.n22 B.t9 275.928
R131 B.n14 B.t0 275.928
R132 B.n245 B.n244 256.663
R133 B.n244 B.n243 235.042
R134 B.n244 B.n2 235.042
R135 B.n88 B.n61 163.367
R136 B.n92 B.n61 163.367
R137 B.n93 B.n92 163.367
R138 B.n94 B.n93 163.367
R139 B.n94 B.n59 163.367
R140 B.n98 B.n59 163.367
R141 B.n99 B.n98 163.367
R142 B.n100 B.n99 163.367
R143 B.n100 B.n55 163.367
R144 B.n105 B.n55 163.367
R145 B.n106 B.n105 163.367
R146 B.n107 B.n106 163.367
R147 B.n107 B.n53 163.367
R148 B.n111 B.n53 163.367
R149 B.n112 B.n111 163.367
R150 B.n113 B.n112 163.367
R151 B.n113 B.n51 163.367
R152 B.n117 B.n51 163.367
R153 B.n118 B.n117 163.367
R154 B.n118 B.n47 163.367
R155 B.n122 B.n47 163.367
R156 B.n123 B.n122 163.367
R157 B.n124 B.n123 163.367
R158 B.n124 B.n45 163.367
R159 B.n128 B.n45 163.367
R160 B.n129 B.n128 163.367
R161 B.n130 B.n129 163.367
R162 B.n130 B.n43 163.367
R163 B.n177 B.n176 163.367
R164 B.n176 B.n29 163.367
R165 B.n172 B.n29 163.367
R166 B.n172 B.n171 163.367
R167 B.n171 B.n170 163.367
R168 B.n170 B.n31 163.367
R169 B.n166 B.n31 163.367
R170 B.n166 B.n165 163.367
R171 B.n165 B.n164 163.367
R172 B.n164 B.n33 163.367
R173 B.n160 B.n33 163.367
R174 B.n160 B.n159 163.367
R175 B.n159 B.n158 163.367
R176 B.n158 B.n35 163.367
R177 B.n154 B.n35 163.367
R178 B.n154 B.n153 163.367
R179 B.n153 B.n152 163.367
R180 B.n152 B.n37 163.367
R181 B.n148 B.n37 163.367
R182 B.n148 B.n147 163.367
R183 B.n147 B.n146 163.367
R184 B.n146 B.n39 163.367
R185 B.n142 B.n39 163.367
R186 B.n142 B.n141 163.367
R187 B.n141 B.n140 163.367
R188 B.n140 B.n41 163.367
R189 B.n136 B.n41 163.367
R190 B.n136 B.n135 163.367
R191 B.n135 B.n134 163.367
R192 B.n220 B.n9 163.367
R193 B.n220 B.n219 163.367
R194 B.n219 B.n218 163.367
R195 B.n218 B.n11 163.367
R196 B.n214 B.n11 163.367
R197 B.n214 B.n213 163.367
R198 B.n213 B.n212 163.367
R199 B.n212 B.n13 163.367
R200 B.n208 B.n13 163.367
R201 B.n208 B.n207 163.367
R202 B.n207 B.n17 163.367
R203 B.n203 B.n17 163.367
R204 B.n203 B.n202 163.367
R205 B.n202 B.n201 163.367
R206 B.n201 B.n19 163.367
R207 B.n197 B.n19 163.367
R208 B.n197 B.n196 163.367
R209 B.n196 B.n195 163.367
R210 B.n195 B.n21 163.367
R211 B.n190 B.n21 163.367
R212 B.n190 B.n189 163.367
R213 B.n189 B.n188 163.367
R214 B.n188 B.n25 163.367
R215 B.n184 B.n25 163.367
R216 B.n184 B.n183 163.367
R217 B.n183 B.n182 163.367
R218 B.n182 B.n27 163.367
R219 B.n178 B.n27 163.367
R220 B.n225 B.n224 163.367
R221 B.n226 B.n225 163.367
R222 B.n226 B.n7 163.367
R223 B.n230 B.n7 163.367
R224 B.n231 B.n230 163.367
R225 B.n232 B.n231 163.367
R226 B.n232 B.n5 163.367
R227 B.n236 B.n5 163.367
R228 B.n237 B.n236 163.367
R229 B.n238 B.n237 163.367
R230 B.n238 B.n3 163.367
R231 B.n242 B.n3 163.367
R232 B.n243 B.n242 163.367
R233 B.n69 B.n2 163.367
R234 B.n70 B.n69 163.367
R235 B.n70 B.n67 163.367
R236 B.n74 B.n67 163.367
R237 B.n75 B.n74 163.367
R238 B.n76 B.n75 163.367
R239 B.n76 B.n65 163.367
R240 B.n80 B.n65 163.367
R241 B.n81 B.n80 163.367
R242 B.n82 B.n81 163.367
R243 B.n82 B.n63 163.367
R244 B.n86 B.n63 163.367
R245 B.n87 B.n86 163.367
R246 B.n103 B.n57 59.5399
R247 B.n50 B.n49 59.5399
R248 B.n193 B.n23 59.5399
R249 B.n16 B.n15 59.5399
R250 B.n223 B.n222 30.1273
R251 B.n179 B.n28 30.1273
R252 B.n133 B.n132 30.1273
R253 B.n89 B.n62 30.1273
R254 B B.n245 18.0485
R255 B.n57 B.n56 13.9641
R256 B.n49 B.n48 13.9641
R257 B.n23 B.n22 13.9641
R258 B.n15 B.n14 13.9641
R259 B.n223 B.n8 10.6151
R260 B.n227 B.n8 10.6151
R261 B.n228 B.n227 10.6151
R262 B.n229 B.n228 10.6151
R263 B.n229 B.n6 10.6151
R264 B.n233 B.n6 10.6151
R265 B.n234 B.n233 10.6151
R266 B.n235 B.n234 10.6151
R267 B.n235 B.n4 10.6151
R268 B.n239 B.n4 10.6151
R269 B.n240 B.n239 10.6151
R270 B.n241 B.n240 10.6151
R271 B.n241 B.n0 10.6151
R272 B.n222 B.n221 10.6151
R273 B.n221 B.n10 10.6151
R274 B.n217 B.n10 10.6151
R275 B.n217 B.n216 10.6151
R276 B.n216 B.n215 10.6151
R277 B.n215 B.n12 10.6151
R278 B.n211 B.n12 10.6151
R279 B.n211 B.n210 10.6151
R280 B.n210 B.n209 10.6151
R281 B.n206 B.n205 10.6151
R282 B.n205 B.n204 10.6151
R283 B.n204 B.n18 10.6151
R284 B.n200 B.n18 10.6151
R285 B.n200 B.n199 10.6151
R286 B.n199 B.n198 10.6151
R287 B.n198 B.n20 10.6151
R288 B.n194 B.n20 10.6151
R289 B.n192 B.n191 10.6151
R290 B.n191 B.n24 10.6151
R291 B.n187 B.n24 10.6151
R292 B.n187 B.n186 10.6151
R293 B.n186 B.n185 10.6151
R294 B.n185 B.n26 10.6151
R295 B.n181 B.n26 10.6151
R296 B.n181 B.n180 10.6151
R297 B.n180 B.n179 10.6151
R298 B.n175 B.n28 10.6151
R299 B.n175 B.n174 10.6151
R300 B.n174 B.n173 10.6151
R301 B.n173 B.n30 10.6151
R302 B.n169 B.n30 10.6151
R303 B.n169 B.n168 10.6151
R304 B.n168 B.n167 10.6151
R305 B.n167 B.n32 10.6151
R306 B.n163 B.n32 10.6151
R307 B.n163 B.n162 10.6151
R308 B.n162 B.n161 10.6151
R309 B.n161 B.n34 10.6151
R310 B.n157 B.n34 10.6151
R311 B.n157 B.n156 10.6151
R312 B.n156 B.n155 10.6151
R313 B.n155 B.n36 10.6151
R314 B.n151 B.n36 10.6151
R315 B.n151 B.n150 10.6151
R316 B.n150 B.n149 10.6151
R317 B.n149 B.n38 10.6151
R318 B.n145 B.n38 10.6151
R319 B.n145 B.n144 10.6151
R320 B.n144 B.n143 10.6151
R321 B.n143 B.n40 10.6151
R322 B.n139 B.n40 10.6151
R323 B.n139 B.n138 10.6151
R324 B.n138 B.n137 10.6151
R325 B.n137 B.n42 10.6151
R326 B.n133 B.n42 10.6151
R327 B.n68 B.n1 10.6151
R328 B.n71 B.n68 10.6151
R329 B.n72 B.n71 10.6151
R330 B.n73 B.n72 10.6151
R331 B.n73 B.n66 10.6151
R332 B.n77 B.n66 10.6151
R333 B.n78 B.n77 10.6151
R334 B.n79 B.n78 10.6151
R335 B.n79 B.n64 10.6151
R336 B.n83 B.n64 10.6151
R337 B.n84 B.n83 10.6151
R338 B.n85 B.n84 10.6151
R339 B.n85 B.n62 10.6151
R340 B.n90 B.n89 10.6151
R341 B.n91 B.n90 10.6151
R342 B.n91 B.n60 10.6151
R343 B.n95 B.n60 10.6151
R344 B.n96 B.n95 10.6151
R345 B.n97 B.n96 10.6151
R346 B.n97 B.n58 10.6151
R347 B.n101 B.n58 10.6151
R348 B.n102 B.n101 10.6151
R349 B.n104 B.n54 10.6151
R350 B.n108 B.n54 10.6151
R351 B.n109 B.n108 10.6151
R352 B.n110 B.n109 10.6151
R353 B.n110 B.n52 10.6151
R354 B.n114 B.n52 10.6151
R355 B.n115 B.n114 10.6151
R356 B.n116 B.n115 10.6151
R357 B.n120 B.n119 10.6151
R358 B.n121 B.n120 10.6151
R359 B.n121 B.n46 10.6151
R360 B.n125 B.n46 10.6151
R361 B.n126 B.n125 10.6151
R362 B.n127 B.n126 10.6151
R363 B.n127 B.n44 10.6151
R364 B.n131 B.n44 10.6151
R365 B.n132 B.n131 10.6151
R366 B.n245 B.n0 8.11757
R367 B.n245 B.n1 8.11757
R368 B.n206 B.n16 7.18099
R369 B.n194 B.n193 7.18099
R370 B.n104 B.n103 7.18099
R371 B.n116 B.n50 7.18099
R372 B.n209 B.n16 3.43465
R373 B.n193 B.n192 3.43465
R374 B.n103 B.n102 3.43465
R375 B.n119 B.n50 3.43465
R376 VN VN.n1 193.03
R377 VN.n0 VN.t1 191.565
R378 VN.n0 VN.t2 191.565
R379 VN.n1 VN.t3 191.565
R380 VN.n1 VN.t0 191.565
R381 VN VN.n0 161.351
R382 VDD2.n2 VDD2.n0 372.199
R383 VDD2.n2 VDD2.n1 345.683
R384 VDD2.n1 VDD2.t2 30.379
R385 VDD2.n1 VDD2.t3 30.379
R386 VDD2.n0 VDD2.t0 30.379
R387 VDD2.n0 VDD2.t1 30.379
R388 VDD2 VDD2.n2 0.0586897
R389 VTAIL.n7 VTAIL.t6 371.94
R390 VTAIL.n0 VTAIL.t5 371.94
R391 VTAIL.n1 VTAIL.t2 371.94
R392 VTAIL.n2 VTAIL.t3 371.94
R393 VTAIL.n6 VTAIL.t0 371.94
R394 VTAIL.n5 VTAIL.t1 371.94
R395 VTAIL.n4 VTAIL.t4 371.94
R396 VTAIL.n3 VTAIL.t7 371.94
R397 VTAIL.n7 VTAIL.n6 13.9272
R398 VTAIL.n3 VTAIL.n2 13.9272
R399 VTAIL.n4 VTAIL.n3 0.62119
R400 VTAIL.n6 VTAIL.n5 0.62119
R401 VTAIL.n2 VTAIL.n1 0.62119
R402 VTAIL.n5 VTAIL.n4 0.470328
R403 VTAIL.n1 VTAIL.n0 0.470328
R404 VTAIL VTAIL.n0 0.369034
R405 VTAIL VTAIL.n7 0.252655
R406 VP.n2 VP.n0 192.649
R407 VP.n1 VP.t2 191.565
R408 VP.n1 VP.t0 191.565
R409 VP.n0 VP.t3 191.565
R410 VP.n0 VP.t1 191.565
R411 VP.n2 VP.n1 161.3
R412 VP VP.n2 0.0516364
R413 VDD1 VDD1.n1 372.724
R414 VDD1 VDD1.n0 345.74
R415 VDD1.n0 VDD1.t2 30.379
R416 VDD1.n0 VDD1.t0 30.379
R417 VDD1.n1 VDD1.t3 30.379
R418 VDD1.n1 VDD1.t1 30.379
C0 VN B 0.53203f
C1 VDD1 B 0.574623f
C2 VP VDD2 0.262665f
C3 VTAIL VP 0.575803f
C4 VP w_n1402_n1186# 1.86025f
C5 VTAIL VDD2 1.9908f
C6 VP VN 2.57445f
C7 w_n1402_n1186# VDD2 0.695598f
C8 VP VDD1 0.575954f
C9 VN VDD2 0.469433f
C10 VTAIL w_n1402_n1186# 1.25897f
C11 VDD1 VDD2 0.497989f
C12 VTAIL VN 0.561697f
C13 VN w_n1402_n1186# 1.69309f
C14 VTAIL VDD1 1.95141f
C15 VDD1 w_n1402_n1186# 0.688093f
C16 VP B 0.810355f
C17 VDD1 VN 0.155047f
C18 B VDD2 0.592063f
C19 VTAIL B 0.72997f
C20 B w_n1402_n1186# 3.43851f
C21 VDD2 VSUBS 0.305044f
C22 VDD1 VSUBS 0.470574f
C23 VTAIL VSUBS 0.206943f
C24 VN VSUBS 3.14774f
C25 VP VSUBS 0.655378f
C26 B VSUBS 1.371726f
C27 w_n1402_n1186# VSUBS 21.417f
C28 VP.t1 VSUBS 0.067055f
C29 VP.t3 VSUBS 0.067055f
C30 VP.n0 VSUBS 0.276931f
C31 VP.t0 VSUBS 0.067055f
C32 VP.t2 VSUBS 0.067055f
C33 VP.n1 VSUBS 0.108977f
C34 VP.n2 VSUBS 1.9202f
C35 VN.t2 VSUBS 0.065541f
C36 VN.t1 VSUBS 0.065541f
C37 VN.n0 VSUBS 0.106533f
C38 VN.t0 VSUBS 0.065541f
C39 VN.t3 VSUBS 0.065541f
C40 VN.n1 VSUBS 0.276949f
C41 B.n0 VSUBS 0.008714f
C42 B.n1 VSUBS 0.008714f
C43 B.n2 VSUBS 0.012887f
C44 B.n3 VSUBS 0.009876f
C45 B.n4 VSUBS 0.009876f
C46 B.n5 VSUBS 0.009876f
C47 B.n6 VSUBS 0.009876f
C48 B.n7 VSUBS 0.009876f
C49 B.n8 VSUBS 0.009876f
C50 B.n9 VSUBS 0.022685f
C51 B.n10 VSUBS 0.009876f
C52 B.n11 VSUBS 0.009876f
C53 B.n12 VSUBS 0.009876f
C54 B.n13 VSUBS 0.009876f
C55 B.t1 VSUBS 0.028401f
C56 B.t2 VSUBS 0.029888f
C57 B.t0 VSUBS 0.030168f
C58 B.n14 VSUBS 0.054126f
C59 B.n15 VSUBS 0.054172f
C60 B.n16 VSUBS 0.022881f
C61 B.n17 VSUBS 0.009876f
C62 B.n18 VSUBS 0.009876f
C63 B.n19 VSUBS 0.009876f
C64 B.n20 VSUBS 0.009876f
C65 B.n21 VSUBS 0.009876f
C66 B.t10 VSUBS 0.028401f
C67 B.t11 VSUBS 0.029888f
C68 B.t9 VSUBS 0.030168f
C69 B.n22 VSUBS 0.054126f
C70 B.n23 VSUBS 0.054172f
C71 B.n24 VSUBS 0.009876f
C72 B.n25 VSUBS 0.009876f
C73 B.n26 VSUBS 0.009876f
C74 B.n27 VSUBS 0.009876f
C75 B.n28 VSUBS 0.021174f
C76 B.n29 VSUBS 0.009876f
C77 B.n30 VSUBS 0.009876f
C78 B.n31 VSUBS 0.009876f
C79 B.n32 VSUBS 0.009876f
C80 B.n33 VSUBS 0.009876f
C81 B.n34 VSUBS 0.009876f
C82 B.n35 VSUBS 0.009876f
C83 B.n36 VSUBS 0.009876f
C84 B.n37 VSUBS 0.009876f
C85 B.n38 VSUBS 0.009876f
C86 B.n39 VSUBS 0.009876f
C87 B.n40 VSUBS 0.009876f
C88 B.n41 VSUBS 0.009876f
C89 B.n42 VSUBS 0.009876f
C90 B.n43 VSUBS 0.022685f
C91 B.n44 VSUBS 0.009876f
C92 B.n45 VSUBS 0.009876f
C93 B.n46 VSUBS 0.009876f
C94 B.n47 VSUBS 0.009876f
C95 B.t8 VSUBS 0.028401f
C96 B.t7 VSUBS 0.029888f
C97 B.t6 VSUBS 0.030168f
C98 B.n48 VSUBS 0.054126f
C99 B.n49 VSUBS 0.054172f
C100 B.n50 VSUBS 0.022881f
C101 B.n51 VSUBS 0.009876f
C102 B.n52 VSUBS 0.009876f
C103 B.n53 VSUBS 0.009876f
C104 B.n54 VSUBS 0.009876f
C105 B.n55 VSUBS 0.009876f
C106 B.t5 VSUBS 0.028401f
C107 B.t4 VSUBS 0.029888f
C108 B.t3 VSUBS 0.030168f
C109 B.n56 VSUBS 0.054126f
C110 B.n57 VSUBS 0.054172f
C111 B.n58 VSUBS 0.009876f
C112 B.n59 VSUBS 0.009876f
C113 B.n60 VSUBS 0.009876f
C114 B.n61 VSUBS 0.009876f
C115 B.n62 VSUBS 0.021174f
C116 B.n63 VSUBS 0.009876f
C117 B.n64 VSUBS 0.009876f
C118 B.n65 VSUBS 0.009876f
C119 B.n66 VSUBS 0.009876f
C120 B.n67 VSUBS 0.009876f
C121 B.n68 VSUBS 0.009876f
C122 B.n69 VSUBS 0.009876f
C123 B.n70 VSUBS 0.009876f
C124 B.n71 VSUBS 0.009876f
C125 B.n72 VSUBS 0.009876f
C126 B.n73 VSUBS 0.009876f
C127 B.n74 VSUBS 0.009876f
C128 B.n75 VSUBS 0.009876f
C129 B.n76 VSUBS 0.009876f
C130 B.n77 VSUBS 0.009876f
C131 B.n78 VSUBS 0.009876f
C132 B.n79 VSUBS 0.009876f
C133 B.n80 VSUBS 0.009876f
C134 B.n81 VSUBS 0.009876f
C135 B.n82 VSUBS 0.009876f
C136 B.n83 VSUBS 0.009876f
C137 B.n84 VSUBS 0.009876f
C138 B.n85 VSUBS 0.009876f
C139 B.n86 VSUBS 0.009876f
C140 B.n87 VSUBS 0.021174f
C141 B.n88 VSUBS 0.022685f
C142 B.n89 VSUBS 0.022685f
C143 B.n90 VSUBS 0.009876f
C144 B.n91 VSUBS 0.009876f
C145 B.n92 VSUBS 0.009876f
C146 B.n93 VSUBS 0.009876f
C147 B.n94 VSUBS 0.009876f
C148 B.n95 VSUBS 0.009876f
C149 B.n96 VSUBS 0.009876f
C150 B.n97 VSUBS 0.009876f
C151 B.n98 VSUBS 0.009876f
C152 B.n99 VSUBS 0.009876f
C153 B.n100 VSUBS 0.009876f
C154 B.n101 VSUBS 0.009876f
C155 B.n102 VSUBS 0.006535f
C156 B.n103 VSUBS 0.022881f
C157 B.n104 VSUBS 0.008278f
C158 B.n105 VSUBS 0.009876f
C159 B.n106 VSUBS 0.009876f
C160 B.n107 VSUBS 0.009876f
C161 B.n108 VSUBS 0.009876f
C162 B.n109 VSUBS 0.009876f
C163 B.n110 VSUBS 0.009876f
C164 B.n111 VSUBS 0.009876f
C165 B.n112 VSUBS 0.009876f
C166 B.n113 VSUBS 0.009876f
C167 B.n114 VSUBS 0.009876f
C168 B.n115 VSUBS 0.009876f
C169 B.n116 VSUBS 0.008278f
C170 B.n117 VSUBS 0.009876f
C171 B.n118 VSUBS 0.009876f
C172 B.n119 VSUBS 0.006535f
C173 B.n120 VSUBS 0.009876f
C174 B.n121 VSUBS 0.009876f
C175 B.n122 VSUBS 0.009876f
C176 B.n123 VSUBS 0.009876f
C177 B.n124 VSUBS 0.009876f
C178 B.n125 VSUBS 0.009876f
C179 B.n126 VSUBS 0.009876f
C180 B.n127 VSUBS 0.009876f
C181 B.n128 VSUBS 0.009876f
C182 B.n129 VSUBS 0.009876f
C183 B.n130 VSUBS 0.009876f
C184 B.n131 VSUBS 0.009876f
C185 B.n132 VSUBS 0.021421f
C186 B.n133 VSUBS 0.022439f
C187 B.n134 VSUBS 0.021174f
C188 B.n135 VSUBS 0.009876f
C189 B.n136 VSUBS 0.009876f
C190 B.n137 VSUBS 0.009876f
C191 B.n138 VSUBS 0.009876f
C192 B.n139 VSUBS 0.009876f
C193 B.n140 VSUBS 0.009876f
C194 B.n141 VSUBS 0.009876f
C195 B.n142 VSUBS 0.009876f
C196 B.n143 VSUBS 0.009876f
C197 B.n144 VSUBS 0.009876f
C198 B.n145 VSUBS 0.009876f
C199 B.n146 VSUBS 0.009876f
C200 B.n147 VSUBS 0.009876f
C201 B.n148 VSUBS 0.009876f
C202 B.n149 VSUBS 0.009876f
C203 B.n150 VSUBS 0.009876f
C204 B.n151 VSUBS 0.009876f
C205 B.n152 VSUBS 0.009876f
C206 B.n153 VSUBS 0.009876f
C207 B.n154 VSUBS 0.009876f
C208 B.n155 VSUBS 0.009876f
C209 B.n156 VSUBS 0.009876f
C210 B.n157 VSUBS 0.009876f
C211 B.n158 VSUBS 0.009876f
C212 B.n159 VSUBS 0.009876f
C213 B.n160 VSUBS 0.009876f
C214 B.n161 VSUBS 0.009876f
C215 B.n162 VSUBS 0.009876f
C216 B.n163 VSUBS 0.009876f
C217 B.n164 VSUBS 0.009876f
C218 B.n165 VSUBS 0.009876f
C219 B.n166 VSUBS 0.009876f
C220 B.n167 VSUBS 0.009876f
C221 B.n168 VSUBS 0.009876f
C222 B.n169 VSUBS 0.009876f
C223 B.n170 VSUBS 0.009876f
C224 B.n171 VSUBS 0.009876f
C225 B.n172 VSUBS 0.009876f
C226 B.n173 VSUBS 0.009876f
C227 B.n174 VSUBS 0.009876f
C228 B.n175 VSUBS 0.009876f
C229 B.n176 VSUBS 0.009876f
C230 B.n177 VSUBS 0.021174f
C231 B.n178 VSUBS 0.022685f
C232 B.n179 VSUBS 0.022685f
C233 B.n180 VSUBS 0.009876f
C234 B.n181 VSUBS 0.009876f
C235 B.n182 VSUBS 0.009876f
C236 B.n183 VSUBS 0.009876f
C237 B.n184 VSUBS 0.009876f
C238 B.n185 VSUBS 0.009876f
C239 B.n186 VSUBS 0.009876f
C240 B.n187 VSUBS 0.009876f
C241 B.n188 VSUBS 0.009876f
C242 B.n189 VSUBS 0.009876f
C243 B.n190 VSUBS 0.009876f
C244 B.n191 VSUBS 0.009876f
C245 B.n192 VSUBS 0.006535f
C246 B.n193 VSUBS 0.022881f
C247 B.n194 VSUBS 0.008278f
C248 B.n195 VSUBS 0.009876f
C249 B.n196 VSUBS 0.009876f
C250 B.n197 VSUBS 0.009876f
C251 B.n198 VSUBS 0.009876f
C252 B.n199 VSUBS 0.009876f
C253 B.n200 VSUBS 0.009876f
C254 B.n201 VSUBS 0.009876f
C255 B.n202 VSUBS 0.009876f
C256 B.n203 VSUBS 0.009876f
C257 B.n204 VSUBS 0.009876f
C258 B.n205 VSUBS 0.009876f
C259 B.n206 VSUBS 0.008278f
C260 B.n207 VSUBS 0.009876f
C261 B.n208 VSUBS 0.009876f
C262 B.n209 VSUBS 0.006535f
C263 B.n210 VSUBS 0.009876f
C264 B.n211 VSUBS 0.009876f
C265 B.n212 VSUBS 0.009876f
C266 B.n213 VSUBS 0.009876f
C267 B.n214 VSUBS 0.009876f
C268 B.n215 VSUBS 0.009876f
C269 B.n216 VSUBS 0.009876f
C270 B.n217 VSUBS 0.009876f
C271 B.n218 VSUBS 0.009876f
C272 B.n219 VSUBS 0.009876f
C273 B.n220 VSUBS 0.009876f
C274 B.n221 VSUBS 0.009876f
C275 B.n222 VSUBS 0.022685f
C276 B.n223 VSUBS 0.021174f
C277 B.n224 VSUBS 0.021174f
C278 B.n225 VSUBS 0.009876f
C279 B.n226 VSUBS 0.009876f
C280 B.n227 VSUBS 0.009876f
C281 B.n228 VSUBS 0.009876f
C282 B.n229 VSUBS 0.009876f
C283 B.n230 VSUBS 0.009876f
C284 B.n231 VSUBS 0.009876f
C285 B.n232 VSUBS 0.009876f
C286 B.n233 VSUBS 0.009876f
C287 B.n234 VSUBS 0.009876f
C288 B.n235 VSUBS 0.009876f
C289 B.n236 VSUBS 0.009876f
C290 B.n237 VSUBS 0.009876f
C291 B.n238 VSUBS 0.009876f
C292 B.n239 VSUBS 0.009876f
C293 B.n240 VSUBS 0.009876f
C294 B.n241 VSUBS 0.009876f
C295 B.n242 VSUBS 0.009876f
C296 B.n243 VSUBS 0.012887f
C297 B.n244 VSUBS 0.013728f
C298 B.n245 VSUBS 0.027299f
.ends

