* NGSPICE file created from diff_pair_sample_1029.ext - technology: sky130A

.subckt diff_pair_sample_1029 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=1.63185 ps=10.22 w=9.89 l=1.53
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=1.63185 ps=10.22 w=9.89 l=1.53
X2 VDD2.t4 VN.t1 VTAIL.t11 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=1.63185 ps=10.22 w=9.89 l=1.53
X3 VTAIL.t7 VN.t2 VDD2.t3 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=1.63185 ps=10.22 w=9.89 l=1.53
X4 VTAIL.t2 VP.t1 VDD1.t4 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=1.63185 ps=10.22 w=9.89 l=1.53
X5 VDD2.t2 VN.t3 VTAIL.t6 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=3.8571 ps=20.56 w=9.89 l=1.53
X6 B.t11 B.t9 B.t10 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=0 ps=0 w=9.89 l=1.53
X7 VDD1.t3 VP.t2 VTAIL.t0 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=1.63185 ps=10.22 w=9.89 l=1.53
X8 B.t8 B.t6 B.t7 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=0 ps=0 w=9.89 l=1.53
X9 B.t5 B.t3 B.t4 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=0 ps=0 w=9.89 l=1.53
X10 VTAIL.t3 VP.t3 VDD1.t2 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=1.63185 ps=10.22 w=9.89 l=1.53
X11 B.t2 B.t0 B.t1 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=3.8571 pd=20.56 as=0 ps=0 w=9.89 l=1.53
X12 VTAIL.t9 VN.t4 VDD2.t1 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=1.63185 ps=10.22 w=9.89 l=1.53
X13 VDD1.t1 VP.t4 VTAIL.t4 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=3.8571 ps=20.56 w=9.89 l=1.53
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=3.8571 ps=20.56 w=9.89 l=1.53
X15 VDD2.t0 VN.t5 VTAIL.t10 w_n2458_n2946# sky130_fd_pr__pfet_01v8 ad=1.63185 pd=10.22 as=3.8571 ps=20.56 w=9.89 l=1.53
R0 VN.n2 VN.t1 187.026
R1 VN.n14 VN.t3 187.026
R2 VN.n11 VN.n10 180.385
R3 VN.n23 VN.n22 180.385
R4 VN.n21 VN.n12 161.3
R5 VN.n20 VN.n19 161.3
R6 VN.n18 VN.n13 161.3
R7 VN.n17 VN.n16 161.3
R8 VN.n9 VN.n0 161.3
R9 VN.n8 VN.n7 161.3
R10 VN.n6 VN.n1 161.3
R11 VN.n5 VN.n4 161.3
R12 VN.n3 VN.t4 155.785
R13 VN.n10 VN.t5 155.785
R14 VN.n15 VN.t2 155.785
R15 VN.n22 VN.t0 155.785
R16 VN.n8 VN.n1 56.5193
R17 VN.n20 VN.n13 56.5193
R18 VN.n3 VN.n2 53.6827
R19 VN.n15 VN.n14 53.6827
R20 VN VN.n23 43.1236
R21 VN.n4 VN.n1 24.4675
R22 VN.n9 VN.n8 24.4675
R23 VN.n16 VN.n13 24.4675
R24 VN.n21 VN.n20 24.4675
R25 VN.n17 VN.n14 18.2406
R26 VN.n5 VN.n2 18.2406
R27 VN.n4 VN.n3 12.234
R28 VN.n16 VN.n15 12.234
R29 VN.n10 VN.n9 5.38324
R30 VN.n22 VN.n21 5.38324
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n218 VTAIL.n170 756.745
R41 VTAIL.n50 VTAIL.n2 756.745
R42 VTAIL.n164 VTAIL.n116 756.745
R43 VTAIL.n108 VTAIL.n60 756.745
R44 VTAIL.n186 VTAIL.n185 585
R45 VTAIL.n191 VTAIL.n190 585
R46 VTAIL.n193 VTAIL.n192 585
R47 VTAIL.n182 VTAIL.n181 585
R48 VTAIL.n199 VTAIL.n198 585
R49 VTAIL.n201 VTAIL.n200 585
R50 VTAIL.n178 VTAIL.n177 585
R51 VTAIL.n208 VTAIL.n207 585
R52 VTAIL.n209 VTAIL.n176 585
R53 VTAIL.n211 VTAIL.n210 585
R54 VTAIL.n174 VTAIL.n173 585
R55 VTAIL.n217 VTAIL.n216 585
R56 VTAIL.n219 VTAIL.n218 585
R57 VTAIL.n18 VTAIL.n17 585
R58 VTAIL.n23 VTAIL.n22 585
R59 VTAIL.n25 VTAIL.n24 585
R60 VTAIL.n14 VTAIL.n13 585
R61 VTAIL.n31 VTAIL.n30 585
R62 VTAIL.n33 VTAIL.n32 585
R63 VTAIL.n10 VTAIL.n9 585
R64 VTAIL.n40 VTAIL.n39 585
R65 VTAIL.n41 VTAIL.n8 585
R66 VTAIL.n43 VTAIL.n42 585
R67 VTAIL.n6 VTAIL.n5 585
R68 VTAIL.n49 VTAIL.n48 585
R69 VTAIL.n51 VTAIL.n50 585
R70 VTAIL.n165 VTAIL.n164 585
R71 VTAIL.n163 VTAIL.n162 585
R72 VTAIL.n120 VTAIL.n119 585
R73 VTAIL.n157 VTAIL.n156 585
R74 VTAIL.n155 VTAIL.n122 585
R75 VTAIL.n154 VTAIL.n153 585
R76 VTAIL.n125 VTAIL.n123 585
R77 VTAIL.n148 VTAIL.n147 585
R78 VTAIL.n146 VTAIL.n145 585
R79 VTAIL.n129 VTAIL.n128 585
R80 VTAIL.n140 VTAIL.n139 585
R81 VTAIL.n138 VTAIL.n137 585
R82 VTAIL.n133 VTAIL.n132 585
R83 VTAIL.n109 VTAIL.n108 585
R84 VTAIL.n107 VTAIL.n106 585
R85 VTAIL.n64 VTAIL.n63 585
R86 VTAIL.n101 VTAIL.n100 585
R87 VTAIL.n99 VTAIL.n66 585
R88 VTAIL.n98 VTAIL.n97 585
R89 VTAIL.n69 VTAIL.n67 585
R90 VTAIL.n92 VTAIL.n91 585
R91 VTAIL.n90 VTAIL.n89 585
R92 VTAIL.n73 VTAIL.n72 585
R93 VTAIL.n84 VTAIL.n83 585
R94 VTAIL.n82 VTAIL.n81 585
R95 VTAIL.n77 VTAIL.n76 585
R96 VTAIL.n187 VTAIL.t10 329.038
R97 VTAIL.n19 VTAIL.t4 329.038
R98 VTAIL.n134 VTAIL.t1 329.038
R99 VTAIL.n78 VTAIL.t6 329.038
R100 VTAIL.n191 VTAIL.n185 171.744
R101 VTAIL.n192 VTAIL.n191 171.744
R102 VTAIL.n192 VTAIL.n181 171.744
R103 VTAIL.n199 VTAIL.n181 171.744
R104 VTAIL.n200 VTAIL.n199 171.744
R105 VTAIL.n200 VTAIL.n177 171.744
R106 VTAIL.n208 VTAIL.n177 171.744
R107 VTAIL.n209 VTAIL.n208 171.744
R108 VTAIL.n210 VTAIL.n209 171.744
R109 VTAIL.n210 VTAIL.n173 171.744
R110 VTAIL.n217 VTAIL.n173 171.744
R111 VTAIL.n218 VTAIL.n217 171.744
R112 VTAIL.n23 VTAIL.n17 171.744
R113 VTAIL.n24 VTAIL.n23 171.744
R114 VTAIL.n24 VTAIL.n13 171.744
R115 VTAIL.n31 VTAIL.n13 171.744
R116 VTAIL.n32 VTAIL.n31 171.744
R117 VTAIL.n32 VTAIL.n9 171.744
R118 VTAIL.n40 VTAIL.n9 171.744
R119 VTAIL.n41 VTAIL.n40 171.744
R120 VTAIL.n42 VTAIL.n41 171.744
R121 VTAIL.n42 VTAIL.n5 171.744
R122 VTAIL.n49 VTAIL.n5 171.744
R123 VTAIL.n50 VTAIL.n49 171.744
R124 VTAIL.n164 VTAIL.n163 171.744
R125 VTAIL.n163 VTAIL.n119 171.744
R126 VTAIL.n156 VTAIL.n119 171.744
R127 VTAIL.n156 VTAIL.n155 171.744
R128 VTAIL.n155 VTAIL.n154 171.744
R129 VTAIL.n154 VTAIL.n123 171.744
R130 VTAIL.n147 VTAIL.n123 171.744
R131 VTAIL.n147 VTAIL.n146 171.744
R132 VTAIL.n146 VTAIL.n128 171.744
R133 VTAIL.n139 VTAIL.n128 171.744
R134 VTAIL.n139 VTAIL.n138 171.744
R135 VTAIL.n138 VTAIL.n132 171.744
R136 VTAIL.n108 VTAIL.n107 171.744
R137 VTAIL.n107 VTAIL.n63 171.744
R138 VTAIL.n100 VTAIL.n63 171.744
R139 VTAIL.n100 VTAIL.n99 171.744
R140 VTAIL.n99 VTAIL.n98 171.744
R141 VTAIL.n98 VTAIL.n67 171.744
R142 VTAIL.n91 VTAIL.n67 171.744
R143 VTAIL.n91 VTAIL.n90 171.744
R144 VTAIL.n90 VTAIL.n72 171.744
R145 VTAIL.n83 VTAIL.n72 171.744
R146 VTAIL.n83 VTAIL.n82 171.744
R147 VTAIL.n82 VTAIL.n76 171.744
R148 VTAIL.t10 VTAIL.n185 85.8723
R149 VTAIL.t4 VTAIL.n17 85.8723
R150 VTAIL.t1 VTAIL.n132 85.8723
R151 VTAIL.t6 VTAIL.n76 85.8723
R152 VTAIL.n115 VTAIL.n114 59.0826
R153 VTAIL.n59 VTAIL.n58 59.0826
R154 VTAIL.n1 VTAIL.n0 59.0824
R155 VTAIL.n57 VTAIL.n56 59.0824
R156 VTAIL.n223 VTAIL.n222 30.8278
R157 VTAIL.n55 VTAIL.n54 30.8278
R158 VTAIL.n169 VTAIL.n168 30.8278
R159 VTAIL.n113 VTAIL.n112 30.8278
R160 VTAIL.n59 VTAIL.n57 24.0996
R161 VTAIL.n223 VTAIL.n169 22.4962
R162 VTAIL.n211 VTAIL.n176 13.1884
R163 VTAIL.n43 VTAIL.n8 13.1884
R164 VTAIL.n157 VTAIL.n122 13.1884
R165 VTAIL.n101 VTAIL.n66 13.1884
R166 VTAIL.n207 VTAIL.n206 12.8005
R167 VTAIL.n212 VTAIL.n174 12.8005
R168 VTAIL.n39 VTAIL.n38 12.8005
R169 VTAIL.n44 VTAIL.n6 12.8005
R170 VTAIL.n158 VTAIL.n120 12.8005
R171 VTAIL.n153 VTAIL.n124 12.8005
R172 VTAIL.n102 VTAIL.n64 12.8005
R173 VTAIL.n97 VTAIL.n68 12.8005
R174 VTAIL.n205 VTAIL.n178 12.0247
R175 VTAIL.n216 VTAIL.n215 12.0247
R176 VTAIL.n37 VTAIL.n10 12.0247
R177 VTAIL.n48 VTAIL.n47 12.0247
R178 VTAIL.n162 VTAIL.n161 12.0247
R179 VTAIL.n152 VTAIL.n125 12.0247
R180 VTAIL.n106 VTAIL.n105 12.0247
R181 VTAIL.n96 VTAIL.n69 12.0247
R182 VTAIL.n202 VTAIL.n201 11.249
R183 VTAIL.n219 VTAIL.n172 11.249
R184 VTAIL.n34 VTAIL.n33 11.249
R185 VTAIL.n51 VTAIL.n4 11.249
R186 VTAIL.n165 VTAIL.n118 11.249
R187 VTAIL.n149 VTAIL.n148 11.249
R188 VTAIL.n109 VTAIL.n62 11.249
R189 VTAIL.n93 VTAIL.n92 11.249
R190 VTAIL.n187 VTAIL.n186 10.7239
R191 VTAIL.n19 VTAIL.n18 10.7239
R192 VTAIL.n134 VTAIL.n133 10.7239
R193 VTAIL.n78 VTAIL.n77 10.7239
R194 VTAIL.n198 VTAIL.n180 10.4732
R195 VTAIL.n220 VTAIL.n170 10.4732
R196 VTAIL.n30 VTAIL.n12 10.4732
R197 VTAIL.n52 VTAIL.n2 10.4732
R198 VTAIL.n166 VTAIL.n116 10.4732
R199 VTAIL.n145 VTAIL.n127 10.4732
R200 VTAIL.n110 VTAIL.n60 10.4732
R201 VTAIL.n89 VTAIL.n71 10.4732
R202 VTAIL.n197 VTAIL.n182 9.69747
R203 VTAIL.n29 VTAIL.n14 9.69747
R204 VTAIL.n144 VTAIL.n129 9.69747
R205 VTAIL.n88 VTAIL.n73 9.69747
R206 VTAIL.n222 VTAIL.n221 9.45567
R207 VTAIL.n54 VTAIL.n53 9.45567
R208 VTAIL.n168 VTAIL.n167 9.45567
R209 VTAIL.n112 VTAIL.n111 9.45567
R210 VTAIL.n221 VTAIL.n220 9.3005
R211 VTAIL.n172 VTAIL.n171 9.3005
R212 VTAIL.n215 VTAIL.n214 9.3005
R213 VTAIL.n213 VTAIL.n212 9.3005
R214 VTAIL.n189 VTAIL.n188 9.3005
R215 VTAIL.n184 VTAIL.n183 9.3005
R216 VTAIL.n195 VTAIL.n194 9.3005
R217 VTAIL.n197 VTAIL.n196 9.3005
R218 VTAIL.n180 VTAIL.n179 9.3005
R219 VTAIL.n203 VTAIL.n202 9.3005
R220 VTAIL.n205 VTAIL.n204 9.3005
R221 VTAIL.n206 VTAIL.n175 9.3005
R222 VTAIL.n53 VTAIL.n52 9.3005
R223 VTAIL.n4 VTAIL.n3 9.3005
R224 VTAIL.n47 VTAIL.n46 9.3005
R225 VTAIL.n45 VTAIL.n44 9.3005
R226 VTAIL.n21 VTAIL.n20 9.3005
R227 VTAIL.n16 VTAIL.n15 9.3005
R228 VTAIL.n27 VTAIL.n26 9.3005
R229 VTAIL.n29 VTAIL.n28 9.3005
R230 VTAIL.n12 VTAIL.n11 9.3005
R231 VTAIL.n35 VTAIL.n34 9.3005
R232 VTAIL.n37 VTAIL.n36 9.3005
R233 VTAIL.n38 VTAIL.n7 9.3005
R234 VTAIL.n136 VTAIL.n135 9.3005
R235 VTAIL.n131 VTAIL.n130 9.3005
R236 VTAIL.n142 VTAIL.n141 9.3005
R237 VTAIL.n144 VTAIL.n143 9.3005
R238 VTAIL.n127 VTAIL.n126 9.3005
R239 VTAIL.n150 VTAIL.n149 9.3005
R240 VTAIL.n152 VTAIL.n151 9.3005
R241 VTAIL.n124 VTAIL.n121 9.3005
R242 VTAIL.n167 VTAIL.n166 9.3005
R243 VTAIL.n118 VTAIL.n117 9.3005
R244 VTAIL.n161 VTAIL.n160 9.3005
R245 VTAIL.n159 VTAIL.n158 9.3005
R246 VTAIL.n80 VTAIL.n79 9.3005
R247 VTAIL.n75 VTAIL.n74 9.3005
R248 VTAIL.n86 VTAIL.n85 9.3005
R249 VTAIL.n88 VTAIL.n87 9.3005
R250 VTAIL.n71 VTAIL.n70 9.3005
R251 VTAIL.n94 VTAIL.n93 9.3005
R252 VTAIL.n96 VTAIL.n95 9.3005
R253 VTAIL.n68 VTAIL.n65 9.3005
R254 VTAIL.n111 VTAIL.n110 9.3005
R255 VTAIL.n62 VTAIL.n61 9.3005
R256 VTAIL.n105 VTAIL.n104 9.3005
R257 VTAIL.n103 VTAIL.n102 9.3005
R258 VTAIL.n194 VTAIL.n193 8.92171
R259 VTAIL.n26 VTAIL.n25 8.92171
R260 VTAIL.n141 VTAIL.n140 8.92171
R261 VTAIL.n85 VTAIL.n84 8.92171
R262 VTAIL.n190 VTAIL.n184 8.14595
R263 VTAIL.n22 VTAIL.n16 8.14595
R264 VTAIL.n137 VTAIL.n131 8.14595
R265 VTAIL.n81 VTAIL.n75 8.14595
R266 VTAIL.n189 VTAIL.n186 7.3702
R267 VTAIL.n21 VTAIL.n18 7.3702
R268 VTAIL.n136 VTAIL.n133 7.3702
R269 VTAIL.n80 VTAIL.n77 7.3702
R270 VTAIL.n190 VTAIL.n189 5.81868
R271 VTAIL.n22 VTAIL.n21 5.81868
R272 VTAIL.n137 VTAIL.n136 5.81868
R273 VTAIL.n81 VTAIL.n80 5.81868
R274 VTAIL.n193 VTAIL.n184 5.04292
R275 VTAIL.n25 VTAIL.n16 5.04292
R276 VTAIL.n140 VTAIL.n131 5.04292
R277 VTAIL.n84 VTAIL.n75 5.04292
R278 VTAIL.n194 VTAIL.n182 4.26717
R279 VTAIL.n26 VTAIL.n14 4.26717
R280 VTAIL.n141 VTAIL.n129 4.26717
R281 VTAIL.n85 VTAIL.n73 4.26717
R282 VTAIL.n198 VTAIL.n197 3.49141
R283 VTAIL.n222 VTAIL.n170 3.49141
R284 VTAIL.n30 VTAIL.n29 3.49141
R285 VTAIL.n54 VTAIL.n2 3.49141
R286 VTAIL.n168 VTAIL.n116 3.49141
R287 VTAIL.n145 VTAIL.n144 3.49141
R288 VTAIL.n112 VTAIL.n60 3.49141
R289 VTAIL.n89 VTAIL.n88 3.49141
R290 VTAIL.n0 VTAIL.t11 3.28715
R291 VTAIL.n0 VTAIL.t9 3.28715
R292 VTAIL.n56 VTAIL.t5 3.28715
R293 VTAIL.n56 VTAIL.t3 3.28715
R294 VTAIL.n114 VTAIL.t0 3.28715
R295 VTAIL.n114 VTAIL.t2 3.28715
R296 VTAIL.n58 VTAIL.t8 3.28715
R297 VTAIL.n58 VTAIL.t7 3.28715
R298 VTAIL.n201 VTAIL.n180 2.71565
R299 VTAIL.n220 VTAIL.n219 2.71565
R300 VTAIL.n33 VTAIL.n12 2.71565
R301 VTAIL.n52 VTAIL.n51 2.71565
R302 VTAIL.n166 VTAIL.n165 2.71565
R303 VTAIL.n148 VTAIL.n127 2.71565
R304 VTAIL.n110 VTAIL.n109 2.71565
R305 VTAIL.n92 VTAIL.n71 2.71565
R306 VTAIL.n188 VTAIL.n187 2.41283
R307 VTAIL.n20 VTAIL.n19 2.41283
R308 VTAIL.n135 VTAIL.n134 2.41283
R309 VTAIL.n79 VTAIL.n78 2.41283
R310 VTAIL.n202 VTAIL.n178 1.93989
R311 VTAIL.n216 VTAIL.n172 1.93989
R312 VTAIL.n34 VTAIL.n10 1.93989
R313 VTAIL.n48 VTAIL.n4 1.93989
R314 VTAIL.n162 VTAIL.n118 1.93989
R315 VTAIL.n149 VTAIL.n125 1.93989
R316 VTAIL.n106 VTAIL.n62 1.93989
R317 VTAIL.n93 VTAIL.n69 1.93989
R318 VTAIL.n113 VTAIL.n59 1.60395
R319 VTAIL.n169 VTAIL.n115 1.60395
R320 VTAIL.n57 VTAIL.n55 1.60395
R321 VTAIL.n115 VTAIL.n113 1.27205
R322 VTAIL.n55 VTAIL.n1 1.27205
R323 VTAIL.n207 VTAIL.n205 1.16414
R324 VTAIL.n215 VTAIL.n174 1.16414
R325 VTAIL.n39 VTAIL.n37 1.16414
R326 VTAIL.n47 VTAIL.n6 1.16414
R327 VTAIL.n161 VTAIL.n120 1.16414
R328 VTAIL.n153 VTAIL.n152 1.16414
R329 VTAIL.n105 VTAIL.n64 1.16414
R330 VTAIL.n97 VTAIL.n96 1.16414
R331 VTAIL VTAIL.n223 1.1449
R332 VTAIL VTAIL.n1 0.459552
R333 VTAIL.n206 VTAIL.n176 0.388379
R334 VTAIL.n212 VTAIL.n211 0.388379
R335 VTAIL.n38 VTAIL.n8 0.388379
R336 VTAIL.n44 VTAIL.n43 0.388379
R337 VTAIL.n158 VTAIL.n157 0.388379
R338 VTAIL.n124 VTAIL.n122 0.388379
R339 VTAIL.n102 VTAIL.n101 0.388379
R340 VTAIL.n68 VTAIL.n66 0.388379
R341 VTAIL.n188 VTAIL.n183 0.155672
R342 VTAIL.n195 VTAIL.n183 0.155672
R343 VTAIL.n196 VTAIL.n195 0.155672
R344 VTAIL.n196 VTAIL.n179 0.155672
R345 VTAIL.n203 VTAIL.n179 0.155672
R346 VTAIL.n204 VTAIL.n203 0.155672
R347 VTAIL.n204 VTAIL.n175 0.155672
R348 VTAIL.n213 VTAIL.n175 0.155672
R349 VTAIL.n214 VTAIL.n213 0.155672
R350 VTAIL.n214 VTAIL.n171 0.155672
R351 VTAIL.n221 VTAIL.n171 0.155672
R352 VTAIL.n20 VTAIL.n15 0.155672
R353 VTAIL.n27 VTAIL.n15 0.155672
R354 VTAIL.n28 VTAIL.n27 0.155672
R355 VTAIL.n28 VTAIL.n11 0.155672
R356 VTAIL.n35 VTAIL.n11 0.155672
R357 VTAIL.n36 VTAIL.n35 0.155672
R358 VTAIL.n36 VTAIL.n7 0.155672
R359 VTAIL.n45 VTAIL.n7 0.155672
R360 VTAIL.n46 VTAIL.n45 0.155672
R361 VTAIL.n46 VTAIL.n3 0.155672
R362 VTAIL.n53 VTAIL.n3 0.155672
R363 VTAIL.n167 VTAIL.n117 0.155672
R364 VTAIL.n160 VTAIL.n117 0.155672
R365 VTAIL.n160 VTAIL.n159 0.155672
R366 VTAIL.n159 VTAIL.n121 0.155672
R367 VTAIL.n151 VTAIL.n121 0.155672
R368 VTAIL.n151 VTAIL.n150 0.155672
R369 VTAIL.n150 VTAIL.n126 0.155672
R370 VTAIL.n143 VTAIL.n126 0.155672
R371 VTAIL.n143 VTAIL.n142 0.155672
R372 VTAIL.n142 VTAIL.n130 0.155672
R373 VTAIL.n135 VTAIL.n130 0.155672
R374 VTAIL.n111 VTAIL.n61 0.155672
R375 VTAIL.n104 VTAIL.n61 0.155672
R376 VTAIL.n104 VTAIL.n103 0.155672
R377 VTAIL.n103 VTAIL.n65 0.155672
R378 VTAIL.n95 VTAIL.n65 0.155672
R379 VTAIL.n95 VTAIL.n94 0.155672
R380 VTAIL.n94 VTAIL.n70 0.155672
R381 VTAIL.n87 VTAIL.n70 0.155672
R382 VTAIL.n87 VTAIL.n86 0.155672
R383 VTAIL.n86 VTAIL.n74 0.155672
R384 VTAIL.n79 VTAIL.n74 0.155672
R385 VDD2.n103 VDD2.n55 756.745
R386 VDD2.n48 VDD2.n0 756.745
R387 VDD2.n104 VDD2.n103 585
R388 VDD2.n102 VDD2.n101 585
R389 VDD2.n59 VDD2.n58 585
R390 VDD2.n96 VDD2.n95 585
R391 VDD2.n94 VDD2.n61 585
R392 VDD2.n93 VDD2.n92 585
R393 VDD2.n64 VDD2.n62 585
R394 VDD2.n87 VDD2.n86 585
R395 VDD2.n85 VDD2.n84 585
R396 VDD2.n68 VDD2.n67 585
R397 VDD2.n79 VDD2.n78 585
R398 VDD2.n77 VDD2.n76 585
R399 VDD2.n72 VDD2.n71 585
R400 VDD2.n16 VDD2.n15 585
R401 VDD2.n21 VDD2.n20 585
R402 VDD2.n23 VDD2.n22 585
R403 VDD2.n12 VDD2.n11 585
R404 VDD2.n29 VDD2.n28 585
R405 VDD2.n31 VDD2.n30 585
R406 VDD2.n8 VDD2.n7 585
R407 VDD2.n38 VDD2.n37 585
R408 VDD2.n39 VDD2.n6 585
R409 VDD2.n41 VDD2.n40 585
R410 VDD2.n4 VDD2.n3 585
R411 VDD2.n47 VDD2.n46 585
R412 VDD2.n49 VDD2.n48 585
R413 VDD2.n17 VDD2.t4 329.038
R414 VDD2.n73 VDD2.t5 329.038
R415 VDD2.n103 VDD2.n102 171.744
R416 VDD2.n102 VDD2.n58 171.744
R417 VDD2.n95 VDD2.n58 171.744
R418 VDD2.n95 VDD2.n94 171.744
R419 VDD2.n94 VDD2.n93 171.744
R420 VDD2.n93 VDD2.n62 171.744
R421 VDD2.n86 VDD2.n62 171.744
R422 VDD2.n86 VDD2.n85 171.744
R423 VDD2.n85 VDD2.n67 171.744
R424 VDD2.n78 VDD2.n67 171.744
R425 VDD2.n78 VDD2.n77 171.744
R426 VDD2.n77 VDD2.n71 171.744
R427 VDD2.n21 VDD2.n15 171.744
R428 VDD2.n22 VDD2.n21 171.744
R429 VDD2.n22 VDD2.n11 171.744
R430 VDD2.n29 VDD2.n11 171.744
R431 VDD2.n30 VDD2.n29 171.744
R432 VDD2.n30 VDD2.n7 171.744
R433 VDD2.n38 VDD2.n7 171.744
R434 VDD2.n39 VDD2.n38 171.744
R435 VDD2.n40 VDD2.n39 171.744
R436 VDD2.n40 VDD2.n3 171.744
R437 VDD2.n47 VDD2.n3 171.744
R438 VDD2.n48 VDD2.n47 171.744
R439 VDD2.t5 VDD2.n71 85.8723
R440 VDD2.t4 VDD2.n15 85.8723
R441 VDD2.n54 VDD2.n53 76.1067
R442 VDD2 VDD2.n109 76.1039
R443 VDD2.n54 VDD2.n52 48.6538
R444 VDD2.n108 VDD2.n107 47.5066
R445 VDD2.n108 VDD2.n54 37.4524
R446 VDD2.n96 VDD2.n61 13.1884
R447 VDD2.n41 VDD2.n6 13.1884
R448 VDD2.n97 VDD2.n59 12.8005
R449 VDD2.n92 VDD2.n63 12.8005
R450 VDD2.n37 VDD2.n36 12.8005
R451 VDD2.n42 VDD2.n4 12.8005
R452 VDD2.n101 VDD2.n100 12.0247
R453 VDD2.n91 VDD2.n64 12.0247
R454 VDD2.n35 VDD2.n8 12.0247
R455 VDD2.n46 VDD2.n45 12.0247
R456 VDD2.n104 VDD2.n57 11.249
R457 VDD2.n88 VDD2.n87 11.249
R458 VDD2.n32 VDD2.n31 11.249
R459 VDD2.n49 VDD2.n2 11.249
R460 VDD2.n73 VDD2.n72 10.7239
R461 VDD2.n17 VDD2.n16 10.7239
R462 VDD2.n105 VDD2.n55 10.4732
R463 VDD2.n84 VDD2.n66 10.4732
R464 VDD2.n28 VDD2.n10 10.4732
R465 VDD2.n50 VDD2.n0 10.4732
R466 VDD2.n83 VDD2.n68 9.69747
R467 VDD2.n27 VDD2.n12 9.69747
R468 VDD2.n107 VDD2.n106 9.45567
R469 VDD2.n52 VDD2.n51 9.45567
R470 VDD2.n75 VDD2.n74 9.3005
R471 VDD2.n70 VDD2.n69 9.3005
R472 VDD2.n81 VDD2.n80 9.3005
R473 VDD2.n83 VDD2.n82 9.3005
R474 VDD2.n66 VDD2.n65 9.3005
R475 VDD2.n89 VDD2.n88 9.3005
R476 VDD2.n91 VDD2.n90 9.3005
R477 VDD2.n63 VDD2.n60 9.3005
R478 VDD2.n106 VDD2.n105 9.3005
R479 VDD2.n57 VDD2.n56 9.3005
R480 VDD2.n100 VDD2.n99 9.3005
R481 VDD2.n98 VDD2.n97 9.3005
R482 VDD2.n51 VDD2.n50 9.3005
R483 VDD2.n2 VDD2.n1 9.3005
R484 VDD2.n45 VDD2.n44 9.3005
R485 VDD2.n43 VDD2.n42 9.3005
R486 VDD2.n19 VDD2.n18 9.3005
R487 VDD2.n14 VDD2.n13 9.3005
R488 VDD2.n25 VDD2.n24 9.3005
R489 VDD2.n27 VDD2.n26 9.3005
R490 VDD2.n10 VDD2.n9 9.3005
R491 VDD2.n33 VDD2.n32 9.3005
R492 VDD2.n35 VDD2.n34 9.3005
R493 VDD2.n36 VDD2.n5 9.3005
R494 VDD2.n80 VDD2.n79 8.92171
R495 VDD2.n24 VDD2.n23 8.92171
R496 VDD2.n76 VDD2.n70 8.14595
R497 VDD2.n20 VDD2.n14 8.14595
R498 VDD2.n75 VDD2.n72 7.3702
R499 VDD2.n19 VDD2.n16 7.3702
R500 VDD2.n76 VDD2.n75 5.81868
R501 VDD2.n20 VDD2.n19 5.81868
R502 VDD2.n79 VDD2.n70 5.04292
R503 VDD2.n23 VDD2.n14 5.04292
R504 VDD2.n80 VDD2.n68 4.26717
R505 VDD2.n24 VDD2.n12 4.26717
R506 VDD2.n107 VDD2.n55 3.49141
R507 VDD2.n84 VDD2.n83 3.49141
R508 VDD2.n28 VDD2.n27 3.49141
R509 VDD2.n52 VDD2.n0 3.49141
R510 VDD2.n109 VDD2.t3 3.28715
R511 VDD2.n109 VDD2.t2 3.28715
R512 VDD2.n53 VDD2.t1 3.28715
R513 VDD2.n53 VDD2.t0 3.28715
R514 VDD2.n105 VDD2.n104 2.71565
R515 VDD2.n87 VDD2.n66 2.71565
R516 VDD2.n31 VDD2.n10 2.71565
R517 VDD2.n50 VDD2.n49 2.71565
R518 VDD2.n74 VDD2.n73 2.41283
R519 VDD2.n18 VDD2.n17 2.41283
R520 VDD2.n101 VDD2.n57 1.93989
R521 VDD2.n88 VDD2.n64 1.93989
R522 VDD2.n32 VDD2.n8 1.93989
R523 VDD2.n46 VDD2.n2 1.93989
R524 VDD2 VDD2.n108 1.26128
R525 VDD2.n100 VDD2.n59 1.16414
R526 VDD2.n92 VDD2.n91 1.16414
R527 VDD2.n37 VDD2.n35 1.16414
R528 VDD2.n45 VDD2.n4 1.16414
R529 VDD2.n97 VDD2.n96 0.388379
R530 VDD2.n63 VDD2.n61 0.388379
R531 VDD2.n36 VDD2.n6 0.388379
R532 VDD2.n42 VDD2.n41 0.388379
R533 VDD2.n106 VDD2.n56 0.155672
R534 VDD2.n99 VDD2.n56 0.155672
R535 VDD2.n99 VDD2.n98 0.155672
R536 VDD2.n98 VDD2.n60 0.155672
R537 VDD2.n90 VDD2.n60 0.155672
R538 VDD2.n90 VDD2.n89 0.155672
R539 VDD2.n89 VDD2.n65 0.155672
R540 VDD2.n82 VDD2.n65 0.155672
R541 VDD2.n82 VDD2.n81 0.155672
R542 VDD2.n81 VDD2.n69 0.155672
R543 VDD2.n74 VDD2.n69 0.155672
R544 VDD2.n18 VDD2.n13 0.155672
R545 VDD2.n25 VDD2.n13 0.155672
R546 VDD2.n26 VDD2.n25 0.155672
R547 VDD2.n26 VDD2.n9 0.155672
R548 VDD2.n33 VDD2.n9 0.155672
R549 VDD2.n34 VDD2.n33 0.155672
R550 VDD2.n34 VDD2.n5 0.155672
R551 VDD2.n43 VDD2.n5 0.155672
R552 VDD2.n44 VDD2.n43 0.155672
R553 VDD2.n44 VDD2.n1 0.155672
R554 VDD2.n51 VDD2.n1 0.155672
R555 VP.n6 VP.t2 187.026
R556 VP.n17 VP.n16 180.385
R557 VP.n32 VP.n31 180.385
R558 VP.n15 VP.n14 180.385
R559 VP.n9 VP.n8 161.3
R560 VP.n10 VP.n5 161.3
R561 VP.n12 VP.n11 161.3
R562 VP.n13 VP.n4 161.3
R563 VP.n30 VP.n0 161.3
R564 VP.n29 VP.n28 161.3
R565 VP.n27 VP.n1 161.3
R566 VP.n26 VP.n25 161.3
R567 VP.n23 VP.n2 161.3
R568 VP.n22 VP.n21 161.3
R569 VP.n20 VP.n3 161.3
R570 VP.n19 VP.n18 161.3
R571 VP.n17 VP.t0 155.785
R572 VP.n24 VP.t3 155.785
R573 VP.n31 VP.t4 155.785
R574 VP.n14 VP.t5 155.785
R575 VP.n7 VP.t1 155.785
R576 VP.n29 VP.n1 56.5193
R577 VP.n22 VP.n3 56.5193
R578 VP.n12 VP.n5 56.5193
R579 VP.n7 VP.n6 53.6827
R580 VP.n16 VP.n15 42.7429
R581 VP.n18 VP.n3 24.4675
R582 VP.n23 VP.n22 24.4675
R583 VP.n25 VP.n1 24.4675
R584 VP.n30 VP.n29 24.4675
R585 VP.n13 VP.n12 24.4675
R586 VP.n8 VP.n5 24.4675
R587 VP.n9 VP.n6 18.2406
R588 VP.n24 VP.n23 12.234
R589 VP.n25 VP.n24 12.234
R590 VP.n8 VP.n7 12.234
R591 VP.n18 VP.n17 5.38324
R592 VP.n31 VP.n30 5.38324
R593 VP.n14 VP.n13 5.38324
R594 VP.n10 VP.n9 0.189894
R595 VP.n11 VP.n10 0.189894
R596 VP.n11 VP.n4 0.189894
R597 VP.n15 VP.n4 0.189894
R598 VP.n19 VP.n16 0.189894
R599 VP.n20 VP.n19 0.189894
R600 VP.n21 VP.n20 0.189894
R601 VP.n21 VP.n2 0.189894
R602 VP.n26 VP.n2 0.189894
R603 VP.n27 VP.n26 0.189894
R604 VP.n28 VP.n27 0.189894
R605 VP.n28 VP.n0 0.189894
R606 VP.n32 VP.n0 0.189894
R607 VP VP.n32 0.0516364
R608 VDD1.n48 VDD1.n0 756.745
R609 VDD1.n101 VDD1.n53 756.745
R610 VDD1.n49 VDD1.n48 585
R611 VDD1.n47 VDD1.n46 585
R612 VDD1.n4 VDD1.n3 585
R613 VDD1.n41 VDD1.n40 585
R614 VDD1.n39 VDD1.n6 585
R615 VDD1.n38 VDD1.n37 585
R616 VDD1.n9 VDD1.n7 585
R617 VDD1.n32 VDD1.n31 585
R618 VDD1.n30 VDD1.n29 585
R619 VDD1.n13 VDD1.n12 585
R620 VDD1.n24 VDD1.n23 585
R621 VDD1.n22 VDD1.n21 585
R622 VDD1.n17 VDD1.n16 585
R623 VDD1.n69 VDD1.n68 585
R624 VDD1.n74 VDD1.n73 585
R625 VDD1.n76 VDD1.n75 585
R626 VDD1.n65 VDD1.n64 585
R627 VDD1.n82 VDD1.n81 585
R628 VDD1.n84 VDD1.n83 585
R629 VDD1.n61 VDD1.n60 585
R630 VDD1.n91 VDD1.n90 585
R631 VDD1.n92 VDD1.n59 585
R632 VDD1.n94 VDD1.n93 585
R633 VDD1.n57 VDD1.n56 585
R634 VDD1.n100 VDD1.n99 585
R635 VDD1.n102 VDD1.n101 585
R636 VDD1.n70 VDD1.t5 329.038
R637 VDD1.n18 VDD1.t3 329.038
R638 VDD1.n48 VDD1.n47 171.744
R639 VDD1.n47 VDD1.n3 171.744
R640 VDD1.n40 VDD1.n3 171.744
R641 VDD1.n40 VDD1.n39 171.744
R642 VDD1.n39 VDD1.n38 171.744
R643 VDD1.n38 VDD1.n7 171.744
R644 VDD1.n31 VDD1.n7 171.744
R645 VDD1.n31 VDD1.n30 171.744
R646 VDD1.n30 VDD1.n12 171.744
R647 VDD1.n23 VDD1.n12 171.744
R648 VDD1.n23 VDD1.n22 171.744
R649 VDD1.n22 VDD1.n16 171.744
R650 VDD1.n74 VDD1.n68 171.744
R651 VDD1.n75 VDD1.n74 171.744
R652 VDD1.n75 VDD1.n64 171.744
R653 VDD1.n82 VDD1.n64 171.744
R654 VDD1.n83 VDD1.n82 171.744
R655 VDD1.n83 VDD1.n60 171.744
R656 VDD1.n91 VDD1.n60 171.744
R657 VDD1.n92 VDD1.n91 171.744
R658 VDD1.n93 VDD1.n92 171.744
R659 VDD1.n93 VDD1.n56 171.744
R660 VDD1.n100 VDD1.n56 171.744
R661 VDD1.n101 VDD1.n100 171.744
R662 VDD1.t3 VDD1.n16 85.8723
R663 VDD1.t5 VDD1.n68 85.8723
R664 VDD1.n107 VDD1.n106 76.1067
R665 VDD1.n109 VDD1.n108 75.7612
R666 VDD1 VDD1.n52 48.7673
R667 VDD1.n107 VDD1.n105 48.6538
R668 VDD1.n109 VDD1.n107 38.8371
R669 VDD1.n41 VDD1.n6 13.1884
R670 VDD1.n94 VDD1.n59 13.1884
R671 VDD1.n42 VDD1.n4 12.8005
R672 VDD1.n37 VDD1.n8 12.8005
R673 VDD1.n90 VDD1.n89 12.8005
R674 VDD1.n95 VDD1.n57 12.8005
R675 VDD1.n46 VDD1.n45 12.0247
R676 VDD1.n36 VDD1.n9 12.0247
R677 VDD1.n88 VDD1.n61 12.0247
R678 VDD1.n99 VDD1.n98 12.0247
R679 VDD1.n49 VDD1.n2 11.249
R680 VDD1.n33 VDD1.n32 11.249
R681 VDD1.n85 VDD1.n84 11.249
R682 VDD1.n102 VDD1.n55 11.249
R683 VDD1.n18 VDD1.n17 10.7239
R684 VDD1.n70 VDD1.n69 10.7239
R685 VDD1.n50 VDD1.n0 10.4732
R686 VDD1.n29 VDD1.n11 10.4732
R687 VDD1.n81 VDD1.n63 10.4732
R688 VDD1.n103 VDD1.n53 10.4732
R689 VDD1.n28 VDD1.n13 9.69747
R690 VDD1.n80 VDD1.n65 9.69747
R691 VDD1.n52 VDD1.n51 9.45567
R692 VDD1.n105 VDD1.n104 9.45567
R693 VDD1.n20 VDD1.n19 9.3005
R694 VDD1.n15 VDD1.n14 9.3005
R695 VDD1.n26 VDD1.n25 9.3005
R696 VDD1.n28 VDD1.n27 9.3005
R697 VDD1.n11 VDD1.n10 9.3005
R698 VDD1.n34 VDD1.n33 9.3005
R699 VDD1.n36 VDD1.n35 9.3005
R700 VDD1.n8 VDD1.n5 9.3005
R701 VDD1.n51 VDD1.n50 9.3005
R702 VDD1.n2 VDD1.n1 9.3005
R703 VDD1.n45 VDD1.n44 9.3005
R704 VDD1.n43 VDD1.n42 9.3005
R705 VDD1.n104 VDD1.n103 9.3005
R706 VDD1.n55 VDD1.n54 9.3005
R707 VDD1.n98 VDD1.n97 9.3005
R708 VDD1.n96 VDD1.n95 9.3005
R709 VDD1.n72 VDD1.n71 9.3005
R710 VDD1.n67 VDD1.n66 9.3005
R711 VDD1.n78 VDD1.n77 9.3005
R712 VDD1.n80 VDD1.n79 9.3005
R713 VDD1.n63 VDD1.n62 9.3005
R714 VDD1.n86 VDD1.n85 9.3005
R715 VDD1.n88 VDD1.n87 9.3005
R716 VDD1.n89 VDD1.n58 9.3005
R717 VDD1.n25 VDD1.n24 8.92171
R718 VDD1.n77 VDD1.n76 8.92171
R719 VDD1.n21 VDD1.n15 8.14595
R720 VDD1.n73 VDD1.n67 8.14595
R721 VDD1.n20 VDD1.n17 7.3702
R722 VDD1.n72 VDD1.n69 7.3702
R723 VDD1.n21 VDD1.n20 5.81868
R724 VDD1.n73 VDD1.n72 5.81868
R725 VDD1.n24 VDD1.n15 5.04292
R726 VDD1.n76 VDD1.n67 5.04292
R727 VDD1.n25 VDD1.n13 4.26717
R728 VDD1.n77 VDD1.n65 4.26717
R729 VDD1.n52 VDD1.n0 3.49141
R730 VDD1.n29 VDD1.n28 3.49141
R731 VDD1.n81 VDD1.n80 3.49141
R732 VDD1.n105 VDD1.n53 3.49141
R733 VDD1.n108 VDD1.t4 3.28715
R734 VDD1.n108 VDD1.t0 3.28715
R735 VDD1.n106 VDD1.t2 3.28715
R736 VDD1.n106 VDD1.t1 3.28715
R737 VDD1.n50 VDD1.n49 2.71565
R738 VDD1.n32 VDD1.n11 2.71565
R739 VDD1.n84 VDD1.n63 2.71565
R740 VDD1.n103 VDD1.n102 2.71565
R741 VDD1.n19 VDD1.n18 2.41283
R742 VDD1.n71 VDD1.n70 2.41283
R743 VDD1.n46 VDD1.n2 1.93989
R744 VDD1.n33 VDD1.n9 1.93989
R745 VDD1.n85 VDD1.n61 1.93989
R746 VDD1.n99 VDD1.n55 1.93989
R747 VDD1.n45 VDD1.n4 1.16414
R748 VDD1.n37 VDD1.n36 1.16414
R749 VDD1.n90 VDD1.n88 1.16414
R750 VDD1.n98 VDD1.n57 1.16414
R751 VDD1.n42 VDD1.n41 0.388379
R752 VDD1.n8 VDD1.n6 0.388379
R753 VDD1.n89 VDD1.n59 0.388379
R754 VDD1.n95 VDD1.n94 0.388379
R755 VDD1 VDD1.n109 0.343172
R756 VDD1.n51 VDD1.n1 0.155672
R757 VDD1.n44 VDD1.n1 0.155672
R758 VDD1.n44 VDD1.n43 0.155672
R759 VDD1.n43 VDD1.n5 0.155672
R760 VDD1.n35 VDD1.n5 0.155672
R761 VDD1.n35 VDD1.n34 0.155672
R762 VDD1.n34 VDD1.n10 0.155672
R763 VDD1.n27 VDD1.n10 0.155672
R764 VDD1.n27 VDD1.n26 0.155672
R765 VDD1.n26 VDD1.n14 0.155672
R766 VDD1.n19 VDD1.n14 0.155672
R767 VDD1.n71 VDD1.n66 0.155672
R768 VDD1.n78 VDD1.n66 0.155672
R769 VDD1.n79 VDD1.n78 0.155672
R770 VDD1.n79 VDD1.n62 0.155672
R771 VDD1.n86 VDD1.n62 0.155672
R772 VDD1.n87 VDD1.n86 0.155672
R773 VDD1.n87 VDD1.n58 0.155672
R774 VDD1.n96 VDD1.n58 0.155672
R775 VDD1.n97 VDD1.n96 0.155672
R776 VDD1.n97 VDD1.n54 0.155672
R777 VDD1.n104 VDD1.n54 0.155672
R778 B.n409 B.n408 585
R779 B.n410 B.n61 585
R780 B.n412 B.n411 585
R781 B.n413 B.n60 585
R782 B.n415 B.n414 585
R783 B.n416 B.n59 585
R784 B.n418 B.n417 585
R785 B.n419 B.n58 585
R786 B.n421 B.n420 585
R787 B.n422 B.n57 585
R788 B.n424 B.n423 585
R789 B.n425 B.n56 585
R790 B.n427 B.n426 585
R791 B.n428 B.n55 585
R792 B.n430 B.n429 585
R793 B.n431 B.n54 585
R794 B.n433 B.n432 585
R795 B.n434 B.n53 585
R796 B.n436 B.n435 585
R797 B.n437 B.n52 585
R798 B.n439 B.n438 585
R799 B.n440 B.n51 585
R800 B.n442 B.n441 585
R801 B.n443 B.n50 585
R802 B.n445 B.n444 585
R803 B.n446 B.n49 585
R804 B.n448 B.n447 585
R805 B.n449 B.n48 585
R806 B.n451 B.n450 585
R807 B.n452 B.n47 585
R808 B.n454 B.n453 585
R809 B.n455 B.n46 585
R810 B.n457 B.n456 585
R811 B.n458 B.n45 585
R812 B.n460 B.n459 585
R813 B.n462 B.n42 585
R814 B.n464 B.n463 585
R815 B.n465 B.n41 585
R816 B.n467 B.n466 585
R817 B.n468 B.n40 585
R818 B.n470 B.n469 585
R819 B.n471 B.n39 585
R820 B.n473 B.n472 585
R821 B.n474 B.n35 585
R822 B.n476 B.n475 585
R823 B.n477 B.n34 585
R824 B.n479 B.n478 585
R825 B.n480 B.n33 585
R826 B.n482 B.n481 585
R827 B.n483 B.n32 585
R828 B.n485 B.n484 585
R829 B.n486 B.n31 585
R830 B.n488 B.n487 585
R831 B.n489 B.n30 585
R832 B.n491 B.n490 585
R833 B.n492 B.n29 585
R834 B.n494 B.n493 585
R835 B.n495 B.n28 585
R836 B.n497 B.n496 585
R837 B.n498 B.n27 585
R838 B.n500 B.n499 585
R839 B.n501 B.n26 585
R840 B.n503 B.n502 585
R841 B.n504 B.n25 585
R842 B.n506 B.n505 585
R843 B.n507 B.n24 585
R844 B.n509 B.n508 585
R845 B.n510 B.n23 585
R846 B.n512 B.n511 585
R847 B.n513 B.n22 585
R848 B.n515 B.n514 585
R849 B.n516 B.n21 585
R850 B.n518 B.n517 585
R851 B.n519 B.n20 585
R852 B.n521 B.n520 585
R853 B.n522 B.n19 585
R854 B.n524 B.n523 585
R855 B.n525 B.n18 585
R856 B.n527 B.n526 585
R857 B.n528 B.n17 585
R858 B.n407 B.n62 585
R859 B.n406 B.n405 585
R860 B.n404 B.n63 585
R861 B.n403 B.n402 585
R862 B.n401 B.n64 585
R863 B.n400 B.n399 585
R864 B.n398 B.n65 585
R865 B.n397 B.n396 585
R866 B.n395 B.n66 585
R867 B.n394 B.n393 585
R868 B.n392 B.n67 585
R869 B.n391 B.n390 585
R870 B.n389 B.n68 585
R871 B.n388 B.n387 585
R872 B.n386 B.n69 585
R873 B.n385 B.n384 585
R874 B.n383 B.n70 585
R875 B.n382 B.n381 585
R876 B.n380 B.n71 585
R877 B.n379 B.n378 585
R878 B.n377 B.n72 585
R879 B.n376 B.n375 585
R880 B.n374 B.n73 585
R881 B.n373 B.n372 585
R882 B.n371 B.n74 585
R883 B.n370 B.n369 585
R884 B.n368 B.n75 585
R885 B.n367 B.n366 585
R886 B.n365 B.n76 585
R887 B.n364 B.n363 585
R888 B.n362 B.n77 585
R889 B.n361 B.n360 585
R890 B.n359 B.n78 585
R891 B.n358 B.n357 585
R892 B.n356 B.n79 585
R893 B.n355 B.n354 585
R894 B.n353 B.n80 585
R895 B.n352 B.n351 585
R896 B.n350 B.n81 585
R897 B.n349 B.n348 585
R898 B.n347 B.n82 585
R899 B.n346 B.n345 585
R900 B.n344 B.n83 585
R901 B.n343 B.n342 585
R902 B.n341 B.n84 585
R903 B.n340 B.n339 585
R904 B.n338 B.n85 585
R905 B.n337 B.n336 585
R906 B.n335 B.n86 585
R907 B.n334 B.n333 585
R908 B.n332 B.n87 585
R909 B.n331 B.n330 585
R910 B.n329 B.n88 585
R911 B.n328 B.n327 585
R912 B.n326 B.n89 585
R913 B.n325 B.n324 585
R914 B.n323 B.n90 585
R915 B.n322 B.n321 585
R916 B.n320 B.n91 585
R917 B.n319 B.n318 585
R918 B.n317 B.n92 585
R919 B.n196 B.n195 585
R920 B.n197 B.n136 585
R921 B.n199 B.n198 585
R922 B.n200 B.n135 585
R923 B.n202 B.n201 585
R924 B.n203 B.n134 585
R925 B.n205 B.n204 585
R926 B.n206 B.n133 585
R927 B.n208 B.n207 585
R928 B.n209 B.n132 585
R929 B.n211 B.n210 585
R930 B.n212 B.n131 585
R931 B.n214 B.n213 585
R932 B.n215 B.n130 585
R933 B.n217 B.n216 585
R934 B.n218 B.n129 585
R935 B.n220 B.n219 585
R936 B.n221 B.n128 585
R937 B.n223 B.n222 585
R938 B.n224 B.n127 585
R939 B.n226 B.n225 585
R940 B.n227 B.n126 585
R941 B.n229 B.n228 585
R942 B.n230 B.n125 585
R943 B.n232 B.n231 585
R944 B.n233 B.n124 585
R945 B.n235 B.n234 585
R946 B.n236 B.n123 585
R947 B.n238 B.n237 585
R948 B.n239 B.n122 585
R949 B.n241 B.n240 585
R950 B.n242 B.n121 585
R951 B.n244 B.n243 585
R952 B.n245 B.n120 585
R953 B.n247 B.n246 585
R954 B.n249 B.n248 585
R955 B.n250 B.n116 585
R956 B.n252 B.n251 585
R957 B.n253 B.n115 585
R958 B.n255 B.n254 585
R959 B.n256 B.n114 585
R960 B.n258 B.n257 585
R961 B.n259 B.n113 585
R962 B.n261 B.n260 585
R963 B.n262 B.n110 585
R964 B.n265 B.n264 585
R965 B.n266 B.n109 585
R966 B.n268 B.n267 585
R967 B.n269 B.n108 585
R968 B.n271 B.n270 585
R969 B.n272 B.n107 585
R970 B.n274 B.n273 585
R971 B.n275 B.n106 585
R972 B.n277 B.n276 585
R973 B.n278 B.n105 585
R974 B.n280 B.n279 585
R975 B.n281 B.n104 585
R976 B.n283 B.n282 585
R977 B.n284 B.n103 585
R978 B.n286 B.n285 585
R979 B.n287 B.n102 585
R980 B.n289 B.n288 585
R981 B.n290 B.n101 585
R982 B.n292 B.n291 585
R983 B.n293 B.n100 585
R984 B.n295 B.n294 585
R985 B.n296 B.n99 585
R986 B.n298 B.n297 585
R987 B.n299 B.n98 585
R988 B.n301 B.n300 585
R989 B.n302 B.n97 585
R990 B.n304 B.n303 585
R991 B.n305 B.n96 585
R992 B.n307 B.n306 585
R993 B.n308 B.n95 585
R994 B.n310 B.n309 585
R995 B.n311 B.n94 585
R996 B.n313 B.n312 585
R997 B.n314 B.n93 585
R998 B.n316 B.n315 585
R999 B.n194 B.n137 585
R1000 B.n193 B.n192 585
R1001 B.n191 B.n138 585
R1002 B.n190 B.n189 585
R1003 B.n188 B.n139 585
R1004 B.n187 B.n186 585
R1005 B.n185 B.n140 585
R1006 B.n184 B.n183 585
R1007 B.n182 B.n141 585
R1008 B.n181 B.n180 585
R1009 B.n179 B.n142 585
R1010 B.n178 B.n177 585
R1011 B.n176 B.n143 585
R1012 B.n175 B.n174 585
R1013 B.n173 B.n144 585
R1014 B.n172 B.n171 585
R1015 B.n170 B.n145 585
R1016 B.n169 B.n168 585
R1017 B.n167 B.n146 585
R1018 B.n166 B.n165 585
R1019 B.n164 B.n147 585
R1020 B.n163 B.n162 585
R1021 B.n161 B.n148 585
R1022 B.n160 B.n159 585
R1023 B.n158 B.n149 585
R1024 B.n157 B.n156 585
R1025 B.n155 B.n150 585
R1026 B.n154 B.n153 585
R1027 B.n152 B.n151 585
R1028 B.n2 B.n0 585
R1029 B.n573 B.n1 585
R1030 B.n572 B.n571 585
R1031 B.n570 B.n3 585
R1032 B.n569 B.n568 585
R1033 B.n567 B.n4 585
R1034 B.n566 B.n565 585
R1035 B.n564 B.n5 585
R1036 B.n563 B.n562 585
R1037 B.n561 B.n6 585
R1038 B.n560 B.n559 585
R1039 B.n558 B.n7 585
R1040 B.n557 B.n556 585
R1041 B.n555 B.n8 585
R1042 B.n554 B.n553 585
R1043 B.n552 B.n9 585
R1044 B.n551 B.n550 585
R1045 B.n549 B.n10 585
R1046 B.n548 B.n547 585
R1047 B.n546 B.n11 585
R1048 B.n545 B.n544 585
R1049 B.n543 B.n12 585
R1050 B.n542 B.n541 585
R1051 B.n540 B.n13 585
R1052 B.n539 B.n538 585
R1053 B.n537 B.n14 585
R1054 B.n536 B.n535 585
R1055 B.n534 B.n15 585
R1056 B.n533 B.n532 585
R1057 B.n531 B.n16 585
R1058 B.n530 B.n529 585
R1059 B.n575 B.n574 585
R1060 B.n195 B.n194 530.939
R1061 B.n530 B.n17 530.939
R1062 B.n315 B.n92 530.939
R1063 B.n409 B.n62 530.939
R1064 B.n111 B.t8 373.515
R1065 B.n43 B.t1 373.515
R1066 B.n117 B.t5 373.515
R1067 B.n36 B.t10 373.515
R1068 B.n111 B.t6 361.334
R1069 B.n117 B.t3 361.334
R1070 B.n36 B.t9 361.334
R1071 B.n43 B.t0 361.334
R1072 B.n112 B.t7 337.442
R1073 B.n44 B.t2 337.442
R1074 B.n118 B.t4 337.442
R1075 B.n37 B.t11 337.442
R1076 B.n194 B.n193 163.367
R1077 B.n193 B.n138 163.367
R1078 B.n189 B.n138 163.367
R1079 B.n189 B.n188 163.367
R1080 B.n188 B.n187 163.367
R1081 B.n187 B.n140 163.367
R1082 B.n183 B.n140 163.367
R1083 B.n183 B.n182 163.367
R1084 B.n182 B.n181 163.367
R1085 B.n181 B.n142 163.367
R1086 B.n177 B.n142 163.367
R1087 B.n177 B.n176 163.367
R1088 B.n176 B.n175 163.367
R1089 B.n175 B.n144 163.367
R1090 B.n171 B.n144 163.367
R1091 B.n171 B.n170 163.367
R1092 B.n170 B.n169 163.367
R1093 B.n169 B.n146 163.367
R1094 B.n165 B.n146 163.367
R1095 B.n165 B.n164 163.367
R1096 B.n164 B.n163 163.367
R1097 B.n163 B.n148 163.367
R1098 B.n159 B.n148 163.367
R1099 B.n159 B.n158 163.367
R1100 B.n158 B.n157 163.367
R1101 B.n157 B.n150 163.367
R1102 B.n153 B.n150 163.367
R1103 B.n153 B.n152 163.367
R1104 B.n152 B.n2 163.367
R1105 B.n574 B.n2 163.367
R1106 B.n574 B.n573 163.367
R1107 B.n573 B.n572 163.367
R1108 B.n572 B.n3 163.367
R1109 B.n568 B.n3 163.367
R1110 B.n568 B.n567 163.367
R1111 B.n567 B.n566 163.367
R1112 B.n566 B.n5 163.367
R1113 B.n562 B.n5 163.367
R1114 B.n562 B.n561 163.367
R1115 B.n561 B.n560 163.367
R1116 B.n560 B.n7 163.367
R1117 B.n556 B.n7 163.367
R1118 B.n556 B.n555 163.367
R1119 B.n555 B.n554 163.367
R1120 B.n554 B.n9 163.367
R1121 B.n550 B.n9 163.367
R1122 B.n550 B.n549 163.367
R1123 B.n549 B.n548 163.367
R1124 B.n548 B.n11 163.367
R1125 B.n544 B.n11 163.367
R1126 B.n544 B.n543 163.367
R1127 B.n543 B.n542 163.367
R1128 B.n542 B.n13 163.367
R1129 B.n538 B.n13 163.367
R1130 B.n538 B.n537 163.367
R1131 B.n537 B.n536 163.367
R1132 B.n536 B.n15 163.367
R1133 B.n532 B.n15 163.367
R1134 B.n532 B.n531 163.367
R1135 B.n531 B.n530 163.367
R1136 B.n195 B.n136 163.367
R1137 B.n199 B.n136 163.367
R1138 B.n200 B.n199 163.367
R1139 B.n201 B.n200 163.367
R1140 B.n201 B.n134 163.367
R1141 B.n205 B.n134 163.367
R1142 B.n206 B.n205 163.367
R1143 B.n207 B.n206 163.367
R1144 B.n207 B.n132 163.367
R1145 B.n211 B.n132 163.367
R1146 B.n212 B.n211 163.367
R1147 B.n213 B.n212 163.367
R1148 B.n213 B.n130 163.367
R1149 B.n217 B.n130 163.367
R1150 B.n218 B.n217 163.367
R1151 B.n219 B.n218 163.367
R1152 B.n219 B.n128 163.367
R1153 B.n223 B.n128 163.367
R1154 B.n224 B.n223 163.367
R1155 B.n225 B.n224 163.367
R1156 B.n225 B.n126 163.367
R1157 B.n229 B.n126 163.367
R1158 B.n230 B.n229 163.367
R1159 B.n231 B.n230 163.367
R1160 B.n231 B.n124 163.367
R1161 B.n235 B.n124 163.367
R1162 B.n236 B.n235 163.367
R1163 B.n237 B.n236 163.367
R1164 B.n237 B.n122 163.367
R1165 B.n241 B.n122 163.367
R1166 B.n242 B.n241 163.367
R1167 B.n243 B.n242 163.367
R1168 B.n243 B.n120 163.367
R1169 B.n247 B.n120 163.367
R1170 B.n248 B.n247 163.367
R1171 B.n248 B.n116 163.367
R1172 B.n252 B.n116 163.367
R1173 B.n253 B.n252 163.367
R1174 B.n254 B.n253 163.367
R1175 B.n254 B.n114 163.367
R1176 B.n258 B.n114 163.367
R1177 B.n259 B.n258 163.367
R1178 B.n260 B.n259 163.367
R1179 B.n260 B.n110 163.367
R1180 B.n265 B.n110 163.367
R1181 B.n266 B.n265 163.367
R1182 B.n267 B.n266 163.367
R1183 B.n267 B.n108 163.367
R1184 B.n271 B.n108 163.367
R1185 B.n272 B.n271 163.367
R1186 B.n273 B.n272 163.367
R1187 B.n273 B.n106 163.367
R1188 B.n277 B.n106 163.367
R1189 B.n278 B.n277 163.367
R1190 B.n279 B.n278 163.367
R1191 B.n279 B.n104 163.367
R1192 B.n283 B.n104 163.367
R1193 B.n284 B.n283 163.367
R1194 B.n285 B.n284 163.367
R1195 B.n285 B.n102 163.367
R1196 B.n289 B.n102 163.367
R1197 B.n290 B.n289 163.367
R1198 B.n291 B.n290 163.367
R1199 B.n291 B.n100 163.367
R1200 B.n295 B.n100 163.367
R1201 B.n296 B.n295 163.367
R1202 B.n297 B.n296 163.367
R1203 B.n297 B.n98 163.367
R1204 B.n301 B.n98 163.367
R1205 B.n302 B.n301 163.367
R1206 B.n303 B.n302 163.367
R1207 B.n303 B.n96 163.367
R1208 B.n307 B.n96 163.367
R1209 B.n308 B.n307 163.367
R1210 B.n309 B.n308 163.367
R1211 B.n309 B.n94 163.367
R1212 B.n313 B.n94 163.367
R1213 B.n314 B.n313 163.367
R1214 B.n315 B.n314 163.367
R1215 B.n319 B.n92 163.367
R1216 B.n320 B.n319 163.367
R1217 B.n321 B.n320 163.367
R1218 B.n321 B.n90 163.367
R1219 B.n325 B.n90 163.367
R1220 B.n326 B.n325 163.367
R1221 B.n327 B.n326 163.367
R1222 B.n327 B.n88 163.367
R1223 B.n331 B.n88 163.367
R1224 B.n332 B.n331 163.367
R1225 B.n333 B.n332 163.367
R1226 B.n333 B.n86 163.367
R1227 B.n337 B.n86 163.367
R1228 B.n338 B.n337 163.367
R1229 B.n339 B.n338 163.367
R1230 B.n339 B.n84 163.367
R1231 B.n343 B.n84 163.367
R1232 B.n344 B.n343 163.367
R1233 B.n345 B.n344 163.367
R1234 B.n345 B.n82 163.367
R1235 B.n349 B.n82 163.367
R1236 B.n350 B.n349 163.367
R1237 B.n351 B.n350 163.367
R1238 B.n351 B.n80 163.367
R1239 B.n355 B.n80 163.367
R1240 B.n356 B.n355 163.367
R1241 B.n357 B.n356 163.367
R1242 B.n357 B.n78 163.367
R1243 B.n361 B.n78 163.367
R1244 B.n362 B.n361 163.367
R1245 B.n363 B.n362 163.367
R1246 B.n363 B.n76 163.367
R1247 B.n367 B.n76 163.367
R1248 B.n368 B.n367 163.367
R1249 B.n369 B.n368 163.367
R1250 B.n369 B.n74 163.367
R1251 B.n373 B.n74 163.367
R1252 B.n374 B.n373 163.367
R1253 B.n375 B.n374 163.367
R1254 B.n375 B.n72 163.367
R1255 B.n379 B.n72 163.367
R1256 B.n380 B.n379 163.367
R1257 B.n381 B.n380 163.367
R1258 B.n381 B.n70 163.367
R1259 B.n385 B.n70 163.367
R1260 B.n386 B.n385 163.367
R1261 B.n387 B.n386 163.367
R1262 B.n387 B.n68 163.367
R1263 B.n391 B.n68 163.367
R1264 B.n392 B.n391 163.367
R1265 B.n393 B.n392 163.367
R1266 B.n393 B.n66 163.367
R1267 B.n397 B.n66 163.367
R1268 B.n398 B.n397 163.367
R1269 B.n399 B.n398 163.367
R1270 B.n399 B.n64 163.367
R1271 B.n403 B.n64 163.367
R1272 B.n404 B.n403 163.367
R1273 B.n405 B.n404 163.367
R1274 B.n405 B.n62 163.367
R1275 B.n526 B.n17 163.367
R1276 B.n526 B.n525 163.367
R1277 B.n525 B.n524 163.367
R1278 B.n524 B.n19 163.367
R1279 B.n520 B.n19 163.367
R1280 B.n520 B.n519 163.367
R1281 B.n519 B.n518 163.367
R1282 B.n518 B.n21 163.367
R1283 B.n514 B.n21 163.367
R1284 B.n514 B.n513 163.367
R1285 B.n513 B.n512 163.367
R1286 B.n512 B.n23 163.367
R1287 B.n508 B.n23 163.367
R1288 B.n508 B.n507 163.367
R1289 B.n507 B.n506 163.367
R1290 B.n506 B.n25 163.367
R1291 B.n502 B.n25 163.367
R1292 B.n502 B.n501 163.367
R1293 B.n501 B.n500 163.367
R1294 B.n500 B.n27 163.367
R1295 B.n496 B.n27 163.367
R1296 B.n496 B.n495 163.367
R1297 B.n495 B.n494 163.367
R1298 B.n494 B.n29 163.367
R1299 B.n490 B.n29 163.367
R1300 B.n490 B.n489 163.367
R1301 B.n489 B.n488 163.367
R1302 B.n488 B.n31 163.367
R1303 B.n484 B.n31 163.367
R1304 B.n484 B.n483 163.367
R1305 B.n483 B.n482 163.367
R1306 B.n482 B.n33 163.367
R1307 B.n478 B.n33 163.367
R1308 B.n478 B.n477 163.367
R1309 B.n477 B.n476 163.367
R1310 B.n476 B.n35 163.367
R1311 B.n472 B.n35 163.367
R1312 B.n472 B.n471 163.367
R1313 B.n471 B.n470 163.367
R1314 B.n470 B.n40 163.367
R1315 B.n466 B.n40 163.367
R1316 B.n466 B.n465 163.367
R1317 B.n465 B.n464 163.367
R1318 B.n464 B.n42 163.367
R1319 B.n459 B.n42 163.367
R1320 B.n459 B.n458 163.367
R1321 B.n458 B.n457 163.367
R1322 B.n457 B.n46 163.367
R1323 B.n453 B.n46 163.367
R1324 B.n453 B.n452 163.367
R1325 B.n452 B.n451 163.367
R1326 B.n451 B.n48 163.367
R1327 B.n447 B.n48 163.367
R1328 B.n447 B.n446 163.367
R1329 B.n446 B.n445 163.367
R1330 B.n445 B.n50 163.367
R1331 B.n441 B.n50 163.367
R1332 B.n441 B.n440 163.367
R1333 B.n440 B.n439 163.367
R1334 B.n439 B.n52 163.367
R1335 B.n435 B.n52 163.367
R1336 B.n435 B.n434 163.367
R1337 B.n434 B.n433 163.367
R1338 B.n433 B.n54 163.367
R1339 B.n429 B.n54 163.367
R1340 B.n429 B.n428 163.367
R1341 B.n428 B.n427 163.367
R1342 B.n427 B.n56 163.367
R1343 B.n423 B.n56 163.367
R1344 B.n423 B.n422 163.367
R1345 B.n422 B.n421 163.367
R1346 B.n421 B.n58 163.367
R1347 B.n417 B.n58 163.367
R1348 B.n417 B.n416 163.367
R1349 B.n416 B.n415 163.367
R1350 B.n415 B.n60 163.367
R1351 B.n411 B.n60 163.367
R1352 B.n411 B.n410 163.367
R1353 B.n410 B.n409 163.367
R1354 B.n263 B.n112 59.5399
R1355 B.n119 B.n118 59.5399
R1356 B.n38 B.n37 59.5399
R1357 B.n461 B.n44 59.5399
R1358 B.n112 B.n111 36.0732
R1359 B.n118 B.n117 36.0732
R1360 B.n37 B.n36 36.0732
R1361 B.n44 B.n43 36.0732
R1362 B.n529 B.n528 34.4981
R1363 B.n408 B.n407 34.4981
R1364 B.n317 B.n316 34.4981
R1365 B.n196 B.n137 34.4981
R1366 B B.n575 18.0485
R1367 B.n528 B.n527 10.6151
R1368 B.n527 B.n18 10.6151
R1369 B.n523 B.n18 10.6151
R1370 B.n523 B.n522 10.6151
R1371 B.n522 B.n521 10.6151
R1372 B.n521 B.n20 10.6151
R1373 B.n517 B.n20 10.6151
R1374 B.n517 B.n516 10.6151
R1375 B.n516 B.n515 10.6151
R1376 B.n515 B.n22 10.6151
R1377 B.n511 B.n22 10.6151
R1378 B.n511 B.n510 10.6151
R1379 B.n510 B.n509 10.6151
R1380 B.n509 B.n24 10.6151
R1381 B.n505 B.n24 10.6151
R1382 B.n505 B.n504 10.6151
R1383 B.n504 B.n503 10.6151
R1384 B.n503 B.n26 10.6151
R1385 B.n499 B.n26 10.6151
R1386 B.n499 B.n498 10.6151
R1387 B.n498 B.n497 10.6151
R1388 B.n497 B.n28 10.6151
R1389 B.n493 B.n28 10.6151
R1390 B.n493 B.n492 10.6151
R1391 B.n492 B.n491 10.6151
R1392 B.n491 B.n30 10.6151
R1393 B.n487 B.n30 10.6151
R1394 B.n487 B.n486 10.6151
R1395 B.n486 B.n485 10.6151
R1396 B.n485 B.n32 10.6151
R1397 B.n481 B.n32 10.6151
R1398 B.n481 B.n480 10.6151
R1399 B.n480 B.n479 10.6151
R1400 B.n479 B.n34 10.6151
R1401 B.n475 B.n474 10.6151
R1402 B.n474 B.n473 10.6151
R1403 B.n473 B.n39 10.6151
R1404 B.n469 B.n39 10.6151
R1405 B.n469 B.n468 10.6151
R1406 B.n468 B.n467 10.6151
R1407 B.n467 B.n41 10.6151
R1408 B.n463 B.n41 10.6151
R1409 B.n463 B.n462 10.6151
R1410 B.n460 B.n45 10.6151
R1411 B.n456 B.n45 10.6151
R1412 B.n456 B.n455 10.6151
R1413 B.n455 B.n454 10.6151
R1414 B.n454 B.n47 10.6151
R1415 B.n450 B.n47 10.6151
R1416 B.n450 B.n449 10.6151
R1417 B.n449 B.n448 10.6151
R1418 B.n448 B.n49 10.6151
R1419 B.n444 B.n49 10.6151
R1420 B.n444 B.n443 10.6151
R1421 B.n443 B.n442 10.6151
R1422 B.n442 B.n51 10.6151
R1423 B.n438 B.n51 10.6151
R1424 B.n438 B.n437 10.6151
R1425 B.n437 B.n436 10.6151
R1426 B.n436 B.n53 10.6151
R1427 B.n432 B.n53 10.6151
R1428 B.n432 B.n431 10.6151
R1429 B.n431 B.n430 10.6151
R1430 B.n430 B.n55 10.6151
R1431 B.n426 B.n55 10.6151
R1432 B.n426 B.n425 10.6151
R1433 B.n425 B.n424 10.6151
R1434 B.n424 B.n57 10.6151
R1435 B.n420 B.n57 10.6151
R1436 B.n420 B.n419 10.6151
R1437 B.n419 B.n418 10.6151
R1438 B.n418 B.n59 10.6151
R1439 B.n414 B.n59 10.6151
R1440 B.n414 B.n413 10.6151
R1441 B.n413 B.n412 10.6151
R1442 B.n412 B.n61 10.6151
R1443 B.n408 B.n61 10.6151
R1444 B.n318 B.n317 10.6151
R1445 B.n318 B.n91 10.6151
R1446 B.n322 B.n91 10.6151
R1447 B.n323 B.n322 10.6151
R1448 B.n324 B.n323 10.6151
R1449 B.n324 B.n89 10.6151
R1450 B.n328 B.n89 10.6151
R1451 B.n329 B.n328 10.6151
R1452 B.n330 B.n329 10.6151
R1453 B.n330 B.n87 10.6151
R1454 B.n334 B.n87 10.6151
R1455 B.n335 B.n334 10.6151
R1456 B.n336 B.n335 10.6151
R1457 B.n336 B.n85 10.6151
R1458 B.n340 B.n85 10.6151
R1459 B.n341 B.n340 10.6151
R1460 B.n342 B.n341 10.6151
R1461 B.n342 B.n83 10.6151
R1462 B.n346 B.n83 10.6151
R1463 B.n347 B.n346 10.6151
R1464 B.n348 B.n347 10.6151
R1465 B.n348 B.n81 10.6151
R1466 B.n352 B.n81 10.6151
R1467 B.n353 B.n352 10.6151
R1468 B.n354 B.n353 10.6151
R1469 B.n354 B.n79 10.6151
R1470 B.n358 B.n79 10.6151
R1471 B.n359 B.n358 10.6151
R1472 B.n360 B.n359 10.6151
R1473 B.n360 B.n77 10.6151
R1474 B.n364 B.n77 10.6151
R1475 B.n365 B.n364 10.6151
R1476 B.n366 B.n365 10.6151
R1477 B.n366 B.n75 10.6151
R1478 B.n370 B.n75 10.6151
R1479 B.n371 B.n370 10.6151
R1480 B.n372 B.n371 10.6151
R1481 B.n372 B.n73 10.6151
R1482 B.n376 B.n73 10.6151
R1483 B.n377 B.n376 10.6151
R1484 B.n378 B.n377 10.6151
R1485 B.n378 B.n71 10.6151
R1486 B.n382 B.n71 10.6151
R1487 B.n383 B.n382 10.6151
R1488 B.n384 B.n383 10.6151
R1489 B.n384 B.n69 10.6151
R1490 B.n388 B.n69 10.6151
R1491 B.n389 B.n388 10.6151
R1492 B.n390 B.n389 10.6151
R1493 B.n390 B.n67 10.6151
R1494 B.n394 B.n67 10.6151
R1495 B.n395 B.n394 10.6151
R1496 B.n396 B.n395 10.6151
R1497 B.n396 B.n65 10.6151
R1498 B.n400 B.n65 10.6151
R1499 B.n401 B.n400 10.6151
R1500 B.n402 B.n401 10.6151
R1501 B.n402 B.n63 10.6151
R1502 B.n406 B.n63 10.6151
R1503 B.n407 B.n406 10.6151
R1504 B.n197 B.n196 10.6151
R1505 B.n198 B.n197 10.6151
R1506 B.n198 B.n135 10.6151
R1507 B.n202 B.n135 10.6151
R1508 B.n203 B.n202 10.6151
R1509 B.n204 B.n203 10.6151
R1510 B.n204 B.n133 10.6151
R1511 B.n208 B.n133 10.6151
R1512 B.n209 B.n208 10.6151
R1513 B.n210 B.n209 10.6151
R1514 B.n210 B.n131 10.6151
R1515 B.n214 B.n131 10.6151
R1516 B.n215 B.n214 10.6151
R1517 B.n216 B.n215 10.6151
R1518 B.n216 B.n129 10.6151
R1519 B.n220 B.n129 10.6151
R1520 B.n221 B.n220 10.6151
R1521 B.n222 B.n221 10.6151
R1522 B.n222 B.n127 10.6151
R1523 B.n226 B.n127 10.6151
R1524 B.n227 B.n226 10.6151
R1525 B.n228 B.n227 10.6151
R1526 B.n228 B.n125 10.6151
R1527 B.n232 B.n125 10.6151
R1528 B.n233 B.n232 10.6151
R1529 B.n234 B.n233 10.6151
R1530 B.n234 B.n123 10.6151
R1531 B.n238 B.n123 10.6151
R1532 B.n239 B.n238 10.6151
R1533 B.n240 B.n239 10.6151
R1534 B.n240 B.n121 10.6151
R1535 B.n244 B.n121 10.6151
R1536 B.n245 B.n244 10.6151
R1537 B.n246 B.n245 10.6151
R1538 B.n250 B.n249 10.6151
R1539 B.n251 B.n250 10.6151
R1540 B.n251 B.n115 10.6151
R1541 B.n255 B.n115 10.6151
R1542 B.n256 B.n255 10.6151
R1543 B.n257 B.n256 10.6151
R1544 B.n257 B.n113 10.6151
R1545 B.n261 B.n113 10.6151
R1546 B.n262 B.n261 10.6151
R1547 B.n264 B.n109 10.6151
R1548 B.n268 B.n109 10.6151
R1549 B.n269 B.n268 10.6151
R1550 B.n270 B.n269 10.6151
R1551 B.n270 B.n107 10.6151
R1552 B.n274 B.n107 10.6151
R1553 B.n275 B.n274 10.6151
R1554 B.n276 B.n275 10.6151
R1555 B.n276 B.n105 10.6151
R1556 B.n280 B.n105 10.6151
R1557 B.n281 B.n280 10.6151
R1558 B.n282 B.n281 10.6151
R1559 B.n282 B.n103 10.6151
R1560 B.n286 B.n103 10.6151
R1561 B.n287 B.n286 10.6151
R1562 B.n288 B.n287 10.6151
R1563 B.n288 B.n101 10.6151
R1564 B.n292 B.n101 10.6151
R1565 B.n293 B.n292 10.6151
R1566 B.n294 B.n293 10.6151
R1567 B.n294 B.n99 10.6151
R1568 B.n298 B.n99 10.6151
R1569 B.n299 B.n298 10.6151
R1570 B.n300 B.n299 10.6151
R1571 B.n300 B.n97 10.6151
R1572 B.n304 B.n97 10.6151
R1573 B.n305 B.n304 10.6151
R1574 B.n306 B.n305 10.6151
R1575 B.n306 B.n95 10.6151
R1576 B.n310 B.n95 10.6151
R1577 B.n311 B.n310 10.6151
R1578 B.n312 B.n311 10.6151
R1579 B.n312 B.n93 10.6151
R1580 B.n316 B.n93 10.6151
R1581 B.n192 B.n137 10.6151
R1582 B.n192 B.n191 10.6151
R1583 B.n191 B.n190 10.6151
R1584 B.n190 B.n139 10.6151
R1585 B.n186 B.n139 10.6151
R1586 B.n186 B.n185 10.6151
R1587 B.n185 B.n184 10.6151
R1588 B.n184 B.n141 10.6151
R1589 B.n180 B.n141 10.6151
R1590 B.n180 B.n179 10.6151
R1591 B.n179 B.n178 10.6151
R1592 B.n178 B.n143 10.6151
R1593 B.n174 B.n143 10.6151
R1594 B.n174 B.n173 10.6151
R1595 B.n173 B.n172 10.6151
R1596 B.n172 B.n145 10.6151
R1597 B.n168 B.n145 10.6151
R1598 B.n168 B.n167 10.6151
R1599 B.n167 B.n166 10.6151
R1600 B.n166 B.n147 10.6151
R1601 B.n162 B.n147 10.6151
R1602 B.n162 B.n161 10.6151
R1603 B.n161 B.n160 10.6151
R1604 B.n160 B.n149 10.6151
R1605 B.n156 B.n149 10.6151
R1606 B.n156 B.n155 10.6151
R1607 B.n155 B.n154 10.6151
R1608 B.n154 B.n151 10.6151
R1609 B.n151 B.n0 10.6151
R1610 B.n571 B.n1 10.6151
R1611 B.n571 B.n570 10.6151
R1612 B.n570 B.n569 10.6151
R1613 B.n569 B.n4 10.6151
R1614 B.n565 B.n4 10.6151
R1615 B.n565 B.n564 10.6151
R1616 B.n564 B.n563 10.6151
R1617 B.n563 B.n6 10.6151
R1618 B.n559 B.n6 10.6151
R1619 B.n559 B.n558 10.6151
R1620 B.n558 B.n557 10.6151
R1621 B.n557 B.n8 10.6151
R1622 B.n553 B.n8 10.6151
R1623 B.n553 B.n552 10.6151
R1624 B.n552 B.n551 10.6151
R1625 B.n551 B.n10 10.6151
R1626 B.n547 B.n10 10.6151
R1627 B.n547 B.n546 10.6151
R1628 B.n546 B.n545 10.6151
R1629 B.n545 B.n12 10.6151
R1630 B.n541 B.n12 10.6151
R1631 B.n541 B.n540 10.6151
R1632 B.n540 B.n539 10.6151
R1633 B.n539 B.n14 10.6151
R1634 B.n535 B.n14 10.6151
R1635 B.n535 B.n534 10.6151
R1636 B.n534 B.n533 10.6151
R1637 B.n533 B.n16 10.6151
R1638 B.n529 B.n16 10.6151
R1639 B.n38 B.n34 9.36635
R1640 B.n461 B.n460 9.36635
R1641 B.n246 B.n119 9.36635
R1642 B.n264 B.n263 9.36635
R1643 B.n575 B.n0 2.81026
R1644 B.n575 B.n1 2.81026
R1645 B.n475 B.n38 1.24928
R1646 B.n462 B.n461 1.24928
R1647 B.n249 B.n119 1.24928
R1648 B.n263 B.n262 1.24928
C0 VP B 1.43623f
C1 VDD2 w_n2458_n2946# 1.92938f
C2 VDD2 VTAIL 7.0524f
C3 VN VDD2 4.93359f
C4 VDD2 VDD1 1.01854f
C5 VDD2 B 1.69077f
C6 VDD2 VP 0.367552f
C7 w_n2458_n2946# VTAIL 2.60231f
C8 VN w_n2458_n2946# 4.36179f
C9 VN VTAIL 4.92937f
C10 w_n2458_n2946# VDD1 1.87872f
C11 VDD1 VTAIL 7.0096f
C12 w_n2458_n2946# B 7.60702f
C13 VTAIL B 2.77246f
C14 VN VDD1 0.149343f
C15 VN B 0.916022f
C16 VP w_n2458_n2946# 4.67659f
C17 VP VTAIL 4.94373f
C18 VDD1 B 1.64223f
C19 VN VP 5.49855f
C20 VP VDD1 5.14864f
C21 VDD2 VSUBS 1.359732f
C22 VDD1 VSUBS 1.309498f
C23 VTAIL VSUBS 0.901408f
C24 VN VSUBS 4.772679f
C25 VP VSUBS 2.015573f
C26 B VSUBS 3.400907f
C27 w_n2458_n2946# VSUBS 89.461395f
C28 B.n0 VSUBS 0.004465f
C29 B.n1 VSUBS 0.004465f
C30 B.n2 VSUBS 0.00706f
C31 B.n3 VSUBS 0.00706f
C32 B.n4 VSUBS 0.00706f
C33 B.n5 VSUBS 0.00706f
C34 B.n6 VSUBS 0.00706f
C35 B.n7 VSUBS 0.00706f
C36 B.n8 VSUBS 0.00706f
C37 B.n9 VSUBS 0.00706f
C38 B.n10 VSUBS 0.00706f
C39 B.n11 VSUBS 0.00706f
C40 B.n12 VSUBS 0.00706f
C41 B.n13 VSUBS 0.00706f
C42 B.n14 VSUBS 0.00706f
C43 B.n15 VSUBS 0.00706f
C44 B.n16 VSUBS 0.00706f
C45 B.n17 VSUBS 0.017372f
C46 B.n18 VSUBS 0.00706f
C47 B.n19 VSUBS 0.00706f
C48 B.n20 VSUBS 0.00706f
C49 B.n21 VSUBS 0.00706f
C50 B.n22 VSUBS 0.00706f
C51 B.n23 VSUBS 0.00706f
C52 B.n24 VSUBS 0.00706f
C53 B.n25 VSUBS 0.00706f
C54 B.n26 VSUBS 0.00706f
C55 B.n27 VSUBS 0.00706f
C56 B.n28 VSUBS 0.00706f
C57 B.n29 VSUBS 0.00706f
C58 B.n30 VSUBS 0.00706f
C59 B.n31 VSUBS 0.00706f
C60 B.n32 VSUBS 0.00706f
C61 B.n33 VSUBS 0.00706f
C62 B.n34 VSUBS 0.006645f
C63 B.n35 VSUBS 0.00706f
C64 B.t11 VSUBS 0.166404f
C65 B.t10 VSUBS 0.186584f
C66 B.t9 VSUBS 0.67757f
C67 B.n36 VSUBS 0.298644f
C68 B.n37 VSUBS 0.219024f
C69 B.n38 VSUBS 0.016358f
C70 B.n39 VSUBS 0.00706f
C71 B.n40 VSUBS 0.00706f
C72 B.n41 VSUBS 0.00706f
C73 B.n42 VSUBS 0.00706f
C74 B.t2 VSUBS 0.166407f
C75 B.t1 VSUBS 0.186587f
C76 B.t0 VSUBS 0.67757f
C77 B.n43 VSUBS 0.298642f
C78 B.n44 VSUBS 0.219021f
C79 B.n45 VSUBS 0.00706f
C80 B.n46 VSUBS 0.00706f
C81 B.n47 VSUBS 0.00706f
C82 B.n48 VSUBS 0.00706f
C83 B.n49 VSUBS 0.00706f
C84 B.n50 VSUBS 0.00706f
C85 B.n51 VSUBS 0.00706f
C86 B.n52 VSUBS 0.00706f
C87 B.n53 VSUBS 0.00706f
C88 B.n54 VSUBS 0.00706f
C89 B.n55 VSUBS 0.00706f
C90 B.n56 VSUBS 0.00706f
C91 B.n57 VSUBS 0.00706f
C92 B.n58 VSUBS 0.00706f
C93 B.n59 VSUBS 0.00706f
C94 B.n60 VSUBS 0.00706f
C95 B.n61 VSUBS 0.00706f
C96 B.n62 VSUBS 0.016891f
C97 B.n63 VSUBS 0.00706f
C98 B.n64 VSUBS 0.00706f
C99 B.n65 VSUBS 0.00706f
C100 B.n66 VSUBS 0.00706f
C101 B.n67 VSUBS 0.00706f
C102 B.n68 VSUBS 0.00706f
C103 B.n69 VSUBS 0.00706f
C104 B.n70 VSUBS 0.00706f
C105 B.n71 VSUBS 0.00706f
C106 B.n72 VSUBS 0.00706f
C107 B.n73 VSUBS 0.00706f
C108 B.n74 VSUBS 0.00706f
C109 B.n75 VSUBS 0.00706f
C110 B.n76 VSUBS 0.00706f
C111 B.n77 VSUBS 0.00706f
C112 B.n78 VSUBS 0.00706f
C113 B.n79 VSUBS 0.00706f
C114 B.n80 VSUBS 0.00706f
C115 B.n81 VSUBS 0.00706f
C116 B.n82 VSUBS 0.00706f
C117 B.n83 VSUBS 0.00706f
C118 B.n84 VSUBS 0.00706f
C119 B.n85 VSUBS 0.00706f
C120 B.n86 VSUBS 0.00706f
C121 B.n87 VSUBS 0.00706f
C122 B.n88 VSUBS 0.00706f
C123 B.n89 VSUBS 0.00706f
C124 B.n90 VSUBS 0.00706f
C125 B.n91 VSUBS 0.00706f
C126 B.n92 VSUBS 0.016891f
C127 B.n93 VSUBS 0.00706f
C128 B.n94 VSUBS 0.00706f
C129 B.n95 VSUBS 0.00706f
C130 B.n96 VSUBS 0.00706f
C131 B.n97 VSUBS 0.00706f
C132 B.n98 VSUBS 0.00706f
C133 B.n99 VSUBS 0.00706f
C134 B.n100 VSUBS 0.00706f
C135 B.n101 VSUBS 0.00706f
C136 B.n102 VSUBS 0.00706f
C137 B.n103 VSUBS 0.00706f
C138 B.n104 VSUBS 0.00706f
C139 B.n105 VSUBS 0.00706f
C140 B.n106 VSUBS 0.00706f
C141 B.n107 VSUBS 0.00706f
C142 B.n108 VSUBS 0.00706f
C143 B.n109 VSUBS 0.00706f
C144 B.n110 VSUBS 0.00706f
C145 B.t7 VSUBS 0.166407f
C146 B.t8 VSUBS 0.186587f
C147 B.t6 VSUBS 0.67757f
C148 B.n111 VSUBS 0.298642f
C149 B.n112 VSUBS 0.219021f
C150 B.n113 VSUBS 0.00706f
C151 B.n114 VSUBS 0.00706f
C152 B.n115 VSUBS 0.00706f
C153 B.n116 VSUBS 0.00706f
C154 B.t4 VSUBS 0.166404f
C155 B.t5 VSUBS 0.186584f
C156 B.t3 VSUBS 0.67757f
C157 B.n117 VSUBS 0.298644f
C158 B.n118 VSUBS 0.219024f
C159 B.n119 VSUBS 0.016358f
C160 B.n120 VSUBS 0.00706f
C161 B.n121 VSUBS 0.00706f
C162 B.n122 VSUBS 0.00706f
C163 B.n123 VSUBS 0.00706f
C164 B.n124 VSUBS 0.00706f
C165 B.n125 VSUBS 0.00706f
C166 B.n126 VSUBS 0.00706f
C167 B.n127 VSUBS 0.00706f
C168 B.n128 VSUBS 0.00706f
C169 B.n129 VSUBS 0.00706f
C170 B.n130 VSUBS 0.00706f
C171 B.n131 VSUBS 0.00706f
C172 B.n132 VSUBS 0.00706f
C173 B.n133 VSUBS 0.00706f
C174 B.n134 VSUBS 0.00706f
C175 B.n135 VSUBS 0.00706f
C176 B.n136 VSUBS 0.00706f
C177 B.n137 VSUBS 0.016891f
C178 B.n138 VSUBS 0.00706f
C179 B.n139 VSUBS 0.00706f
C180 B.n140 VSUBS 0.00706f
C181 B.n141 VSUBS 0.00706f
C182 B.n142 VSUBS 0.00706f
C183 B.n143 VSUBS 0.00706f
C184 B.n144 VSUBS 0.00706f
C185 B.n145 VSUBS 0.00706f
C186 B.n146 VSUBS 0.00706f
C187 B.n147 VSUBS 0.00706f
C188 B.n148 VSUBS 0.00706f
C189 B.n149 VSUBS 0.00706f
C190 B.n150 VSUBS 0.00706f
C191 B.n151 VSUBS 0.00706f
C192 B.n152 VSUBS 0.00706f
C193 B.n153 VSUBS 0.00706f
C194 B.n154 VSUBS 0.00706f
C195 B.n155 VSUBS 0.00706f
C196 B.n156 VSUBS 0.00706f
C197 B.n157 VSUBS 0.00706f
C198 B.n158 VSUBS 0.00706f
C199 B.n159 VSUBS 0.00706f
C200 B.n160 VSUBS 0.00706f
C201 B.n161 VSUBS 0.00706f
C202 B.n162 VSUBS 0.00706f
C203 B.n163 VSUBS 0.00706f
C204 B.n164 VSUBS 0.00706f
C205 B.n165 VSUBS 0.00706f
C206 B.n166 VSUBS 0.00706f
C207 B.n167 VSUBS 0.00706f
C208 B.n168 VSUBS 0.00706f
C209 B.n169 VSUBS 0.00706f
C210 B.n170 VSUBS 0.00706f
C211 B.n171 VSUBS 0.00706f
C212 B.n172 VSUBS 0.00706f
C213 B.n173 VSUBS 0.00706f
C214 B.n174 VSUBS 0.00706f
C215 B.n175 VSUBS 0.00706f
C216 B.n176 VSUBS 0.00706f
C217 B.n177 VSUBS 0.00706f
C218 B.n178 VSUBS 0.00706f
C219 B.n179 VSUBS 0.00706f
C220 B.n180 VSUBS 0.00706f
C221 B.n181 VSUBS 0.00706f
C222 B.n182 VSUBS 0.00706f
C223 B.n183 VSUBS 0.00706f
C224 B.n184 VSUBS 0.00706f
C225 B.n185 VSUBS 0.00706f
C226 B.n186 VSUBS 0.00706f
C227 B.n187 VSUBS 0.00706f
C228 B.n188 VSUBS 0.00706f
C229 B.n189 VSUBS 0.00706f
C230 B.n190 VSUBS 0.00706f
C231 B.n191 VSUBS 0.00706f
C232 B.n192 VSUBS 0.00706f
C233 B.n193 VSUBS 0.00706f
C234 B.n194 VSUBS 0.016891f
C235 B.n195 VSUBS 0.017372f
C236 B.n196 VSUBS 0.017372f
C237 B.n197 VSUBS 0.00706f
C238 B.n198 VSUBS 0.00706f
C239 B.n199 VSUBS 0.00706f
C240 B.n200 VSUBS 0.00706f
C241 B.n201 VSUBS 0.00706f
C242 B.n202 VSUBS 0.00706f
C243 B.n203 VSUBS 0.00706f
C244 B.n204 VSUBS 0.00706f
C245 B.n205 VSUBS 0.00706f
C246 B.n206 VSUBS 0.00706f
C247 B.n207 VSUBS 0.00706f
C248 B.n208 VSUBS 0.00706f
C249 B.n209 VSUBS 0.00706f
C250 B.n210 VSUBS 0.00706f
C251 B.n211 VSUBS 0.00706f
C252 B.n212 VSUBS 0.00706f
C253 B.n213 VSUBS 0.00706f
C254 B.n214 VSUBS 0.00706f
C255 B.n215 VSUBS 0.00706f
C256 B.n216 VSUBS 0.00706f
C257 B.n217 VSUBS 0.00706f
C258 B.n218 VSUBS 0.00706f
C259 B.n219 VSUBS 0.00706f
C260 B.n220 VSUBS 0.00706f
C261 B.n221 VSUBS 0.00706f
C262 B.n222 VSUBS 0.00706f
C263 B.n223 VSUBS 0.00706f
C264 B.n224 VSUBS 0.00706f
C265 B.n225 VSUBS 0.00706f
C266 B.n226 VSUBS 0.00706f
C267 B.n227 VSUBS 0.00706f
C268 B.n228 VSUBS 0.00706f
C269 B.n229 VSUBS 0.00706f
C270 B.n230 VSUBS 0.00706f
C271 B.n231 VSUBS 0.00706f
C272 B.n232 VSUBS 0.00706f
C273 B.n233 VSUBS 0.00706f
C274 B.n234 VSUBS 0.00706f
C275 B.n235 VSUBS 0.00706f
C276 B.n236 VSUBS 0.00706f
C277 B.n237 VSUBS 0.00706f
C278 B.n238 VSUBS 0.00706f
C279 B.n239 VSUBS 0.00706f
C280 B.n240 VSUBS 0.00706f
C281 B.n241 VSUBS 0.00706f
C282 B.n242 VSUBS 0.00706f
C283 B.n243 VSUBS 0.00706f
C284 B.n244 VSUBS 0.00706f
C285 B.n245 VSUBS 0.00706f
C286 B.n246 VSUBS 0.006645f
C287 B.n247 VSUBS 0.00706f
C288 B.n248 VSUBS 0.00706f
C289 B.n249 VSUBS 0.003945f
C290 B.n250 VSUBS 0.00706f
C291 B.n251 VSUBS 0.00706f
C292 B.n252 VSUBS 0.00706f
C293 B.n253 VSUBS 0.00706f
C294 B.n254 VSUBS 0.00706f
C295 B.n255 VSUBS 0.00706f
C296 B.n256 VSUBS 0.00706f
C297 B.n257 VSUBS 0.00706f
C298 B.n258 VSUBS 0.00706f
C299 B.n259 VSUBS 0.00706f
C300 B.n260 VSUBS 0.00706f
C301 B.n261 VSUBS 0.00706f
C302 B.n262 VSUBS 0.003945f
C303 B.n263 VSUBS 0.016358f
C304 B.n264 VSUBS 0.006645f
C305 B.n265 VSUBS 0.00706f
C306 B.n266 VSUBS 0.00706f
C307 B.n267 VSUBS 0.00706f
C308 B.n268 VSUBS 0.00706f
C309 B.n269 VSUBS 0.00706f
C310 B.n270 VSUBS 0.00706f
C311 B.n271 VSUBS 0.00706f
C312 B.n272 VSUBS 0.00706f
C313 B.n273 VSUBS 0.00706f
C314 B.n274 VSUBS 0.00706f
C315 B.n275 VSUBS 0.00706f
C316 B.n276 VSUBS 0.00706f
C317 B.n277 VSUBS 0.00706f
C318 B.n278 VSUBS 0.00706f
C319 B.n279 VSUBS 0.00706f
C320 B.n280 VSUBS 0.00706f
C321 B.n281 VSUBS 0.00706f
C322 B.n282 VSUBS 0.00706f
C323 B.n283 VSUBS 0.00706f
C324 B.n284 VSUBS 0.00706f
C325 B.n285 VSUBS 0.00706f
C326 B.n286 VSUBS 0.00706f
C327 B.n287 VSUBS 0.00706f
C328 B.n288 VSUBS 0.00706f
C329 B.n289 VSUBS 0.00706f
C330 B.n290 VSUBS 0.00706f
C331 B.n291 VSUBS 0.00706f
C332 B.n292 VSUBS 0.00706f
C333 B.n293 VSUBS 0.00706f
C334 B.n294 VSUBS 0.00706f
C335 B.n295 VSUBS 0.00706f
C336 B.n296 VSUBS 0.00706f
C337 B.n297 VSUBS 0.00706f
C338 B.n298 VSUBS 0.00706f
C339 B.n299 VSUBS 0.00706f
C340 B.n300 VSUBS 0.00706f
C341 B.n301 VSUBS 0.00706f
C342 B.n302 VSUBS 0.00706f
C343 B.n303 VSUBS 0.00706f
C344 B.n304 VSUBS 0.00706f
C345 B.n305 VSUBS 0.00706f
C346 B.n306 VSUBS 0.00706f
C347 B.n307 VSUBS 0.00706f
C348 B.n308 VSUBS 0.00706f
C349 B.n309 VSUBS 0.00706f
C350 B.n310 VSUBS 0.00706f
C351 B.n311 VSUBS 0.00706f
C352 B.n312 VSUBS 0.00706f
C353 B.n313 VSUBS 0.00706f
C354 B.n314 VSUBS 0.00706f
C355 B.n315 VSUBS 0.017372f
C356 B.n316 VSUBS 0.017372f
C357 B.n317 VSUBS 0.016891f
C358 B.n318 VSUBS 0.00706f
C359 B.n319 VSUBS 0.00706f
C360 B.n320 VSUBS 0.00706f
C361 B.n321 VSUBS 0.00706f
C362 B.n322 VSUBS 0.00706f
C363 B.n323 VSUBS 0.00706f
C364 B.n324 VSUBS 0.00706f
C365 B.n325 VSUBS 0.00706f
C366 B.n326 VSUBS 0.00706f
C367 B.n327 VSUBS 0.00706f
C368 B.n328 VSUBS 0.00706f
C369 B.n329 VSUBS 0.00706f
C370 B.n330 VSUBS 0.00706f
C371 B.n331 VSUBS 0.00706f
C372 B.n332 VSUBS 0.00706f
C373 B.n333 VSUBS 0.00706f
C374 B.n334 VSUBS 0.00706f
C375 B.n335 VSUBS 0.00706f
C376 B.n336 VSUBS 0.00706f
C377 B.n337 VSUBS 0.00706f
C378 B.n338 VSUBS 0.00706f
C379 B.n339 VSUBS 0.00706f
C380 B.n340 VSUBS 0.00706f
C381 B.n341 VSUBS 0.00706f
C382 B.n342 VSUBS 0.00706f
C383 B.n343 VSUBS 0.00706f
C384 B.n344 VSUBS 0.00706f
C385 B.n345 VSUBS 0.00706f
C386 B.n346 VSUBS 0.00706f
C387 B.n347 VSUBS 0.00706f
C388 B.n348 VSUBS 0.00706f
C389 B.n349 VSUBS 0.00706f
C390 B.n350 VSUBS 0.00706f
C391 B.n351 VSUBS 0.00706f
C392 B.n352 VSUBS 0.00706f
C393 B.n353 VSUBS 0.00706f
C394 B.n354 VSUBS 0.00706f
C395 B.n355 VSUBS 0.00706f
C396 B.n356 VSUBS 0.00706f
C397 B.n357 VSUBS 0.00706f
C398 B.n358 VSUBS 0.00706f
C399 B.n359 VSUBS 0.00706f
C400 B.n360 VSUBS 0.00706f
C401 B.n361 VSUBS 0.00706f
C402 B.n362 VSUBS 0.00706f
C403 B.n363 VSUBS 0.00706f
C404 B.n364 VSUBS 0.00706f
C405 B.n365 VSUBS 0.00706f
C406 B.n366 VSUBS 0.00706f
C407 B.n367 VSUBS 0.00706f
C408 B.n368 VSUBS 0.00706f
C409 B.n369 VSUBS 0.00706f
C410 B.n370 VSUBS 0.00706f
C411 B.n371 VSUBS 0.00706f
C412 B.n372 VSUBS 0.00706f
C413 B.n373 VSUBS 0.00706f
C414 B.n374 VSUBS 0.00706f
C415 B.n375 VSUBS 0.00706f
C416 B.n376 VSUBS 0.00706f
C417 B.n377 VSUBS 0.00706f
C418 B.n378 VSUBS 0.00706f
C419 B.n379 VSUBS 0.00706f
C420 B.n380 VSUBS 0.00706f
C421 B.n381 VSUBS 0.00706f
C422 B.n382 VSUBS 0.00706f
C423 B.n383 VSUBS 0.00706f
C424 B.n384 VSUBS 0.00706f
C425 B.n385 VSUBS 0.00706f
C426 B.n386 VSUBS 0.00706f
C427 B.n387 VSUBS 0.00706f
C428 B.n388 VSUBS 0.00706f
C429 B.n389 VSUBS 0.00706f
C430 B.n390 VSUBS 0.00706f
C431 B.n391 VSUBS 0.00706f
C432 B.n392 VSUBS 0.00706f
C433 B.n393 VSUBS 0.00706f
C434 B.n394 VSUBS 0.00706f
C435 B.n395 VSUBS 0.00706f
C436 B.n396 VSUBS 0.00706f
C437 B.n397 VSUBS 0.00706f
C438 B.n398 VSUBS 0.00706f
C439 B.n399 VSUBS 0.00706f
C440 B.n400 VSUBS 0.00706f
C441 B.n401 VSUBS 0.00706f
C442 B.n402 VSUBS 0.00706f
C443 B.n403 VSUBS 0.00706f
C444 B.n404 VSUBS 0.00706f
C445 B.n405 VSUBS 0.00706f
C446 B.n406 VSUBS 0.00706f
C447 B.n407 VSUBS 0.01768f
C448 B.n408 VSUBS 0.016583f
C449 B.n409 VSUBS 0.017372f
C450 B.n410 VSUBS 0.00706f
C451 B.n411 VSUBS 0.00706f
C452 B.n412 VSUBS 0.00706f
C453 B.n413 VSUBS 0.00706f
C454 B.n414 VSUBS 0.00706f
C455 B.n415 VSUBS 0.00706f
C456 B.n416 VSUBS 0.00706f
C457 B.n417 VSUBS 0.00706f
C458 B.n418 VSUBS 0.00706f
C459 B.n419 VSUBS 0.00706f
C460 B.n420 VSUBS 0.00706f
C461 B.n421 VSUBS 0.00706f
C462 B.n422 VSUBS 0.00706f
C463 B.n423 VSUBS 0.00706f
C464 B.n424 VSUBS 0.00706f
C465 B.n425 VSUBS 0.00706f
C466 B.n426 VSUBS 0.00706f
C467 B.n427 VSUBS 0.00706f
C468 B.n428 VSUBS 0.00706f
C469 B.n429 VSUBS 0.00706f
C470 B.n430 VSUBS 0.00706f
C471 B.n431 VSUBS 0.00706f
C472 B.n432 VSUBS 0.00706f
C473 B.n433 VSUBS 0.00706f
C474 B.n434 VSUBS 0.00706f
C475 B.n435 VSUBS 0.00706f
C476 B.n436 VSUBS 0.00706f
C477 B.n437 VSUBS 0.00706f
C478 B.n438 VSUBS 0.00706f
C479 B.n439 VSUBS 0.00706f
C480 B.n440 VSUBS 0.00706f
C481 B.n441 VSUBS 0.00706f
C482 B.n442 VSUBS 0.00706f
C483 B.n443 VSUBS 0.00706f
C484 B.n444 VSUBS 0.00706f
C485 B.n445 VSUBS 0.00706f
C486 B.n446 VSUBS 0.00706f
C487 B.n447 VSUBS 0.00706f
C488 B.n448 VSUBS 0.00706f
C489 B.n449 VSUBS 0.00706f
C490 B.n450 VSUBS 0.00706f
C491 B.n451 VSUBS 0.00706f
C492 B.n452 VSUBS 0.00706f
C493 B.n453 VSUBS 0.00706f
C494 B.n454 VSUBS 0.00706f
C495 B.n455 VSUBS 0.00706f
C496 B.n456 VSUBS 0.00706f
C497 B.n457 VSUBS 0.00706f
C498 B.n458 VSUBS 0.00706f
C499 B.n459 VSUBS 0.00706f
C500 B.n460 VSUBS 0.006645f
C501 B.n461 VSUBS 0.016358f
C502 B.n462 VSUBS 0.003945f
C503 B.n463 VSUBS 0.00706f
C504 B.n464 VSUBS 0.00706f
C505 B.n465 VSUBS 0.00706f
C506 B.n466 VSUBS 0.00706f
C507 B.n467 VSUBS 0.00706f
C508 B.n468 VSUBS 0.00706f
C509 B.n469 VSUBS 0.00706f
C510 B.n470 VSUBS 0.00706f
C511 B.n471 VSUBS 0.00706f
C512 B.n472 VSUBS 0.00706f
C513 B.n473 VSUBS 0.00706f
C514 B.n474 VSUBS 0.00706f
C515 B.n475 VSUBS 0.003945f
C516 B.n476 VSUBS 0.00706f
C517 B.n477 VSUBS 0.00706f
C518 B.n478 VSUBS 0.00706f
C519 B.n479 VSUBS 0.00706f
C520 B.n480 VSUBS 0.00706f
C521 B.n481 VSUBS 0.00706f
C522 B.n482 VSUBS 0.00706f
C523 B.n483 VSUBS 0.00706f
C524 B.n484 VSUBS 0.00706f
C525 B.n485 VSUBS 0.00706f
C526 B.n486 VSUBS 0.00706f
C527 B.n487 VSUBS 0.00706f
C528 B.n488 VSUBS 0.00706f
C529 B.n489 VSUBS 0.00706f
C530 B.n490 VSUBS 0.00706f
C531 B.n491 VSUBS 0.00706f
C532 B.n492 VSUBS 0.00706f
C533 B.n493 VSUBS 0.00706f
C534 B.n494 VSUBS 0.00706f
C535 B.n495 VSUBS 0.00706f
C536 B.n496 VSUBS 0.00706f
C537 B.n497 VSUBS 0.00706f
C538 B.n498 VSUBS 0.00706f
C539 B.n499 VSUBS 0.00706f
C540 B.n500 VSUBS 0.00706f
C541 B.n501 VSUBS 0.00706f
C542 B.n502 VSUBS 0.00706f
C543 B.n503 VSUBS 0.00706f
C544 B.n504 VSUBS 0.00706f
C545 B.n505 VSUBS 0.00706f
C546 B.n506 VSUBS 0.00706f
C547 B.n507 VSUBS 0.00706f
C548 B.n508 VSUBS 0.00706f
C549 B.n509 VSUBS 0.00706f
C550 B.n510 VSUBS 0.00706f
C551 B.n511 VSUBS 0.00706f
C552 B.n512 VSUBS 0.00706f
C553 B.n513 VSUBS 0.00706f
C554 B.n514 VSUBS 0.00706f
C555 B.n515 VSUBS 0.00706f
C556 B.n516 VSUBS 0.00706f
C557 B.n517 VSUBS 0.00706f
C558 B.n518 VSUBS 0.00706f
C559 B.n519 VSUBS 0.00706f
C560 B.n520 VSUBS 0.00706f
C561 B.n521 VSUBS 0.00706f
C562 B.n522 VSUBS 0.00706f
C563 B.n523 VSUBS 0.00706f
C564 B.n524 VSUBS 0.00706f
C565 B.n525 VSUBS 0.00706f
C566 B.n526 VSUBS 0.00706f
C567 B.n527 VSUBS 0.00706f
C568 B.n528 VSUBS 0.017372f
C569 B.n529 VSUBS 0.016891f
C570 B.n530 VSUBS 0.016891f
C571 B.n531 VSUBS 0.00706f
C572 B.n532 VSUBS 0.00706f
C573 B.n533 VSUBS 0.00706f
C574 B.n534 VSUBS 0.00706f
C575 B.n535 VSUBS 0.00706f
C576 B.n536 VSUBS 0.00706f
C577 B.n537 VSUBS 0.00706f
C578 B.n538 VSUBS 0.00706f
C579 B.n539 VSUBS 0.00706f
C580 B.n540 VSUBS 0.00706f
C581 B.n541 VSUBS 0.00706f
C582 B.n542 VSUBS 0.00706f
C583 B.n543 VSUBS 0.00706f
C584 B.n544 VSUBS 0.00706f
C585 B.n545 VSUBS 0.00706f
C586 B.n546 VSUBS 0.00706f
C587 B.n547 VSUBS 0.00706f
C588 B.n548 VSUBS 0.00706f
C589 B.n549 VSUBS 0.00706f
C590 B.n550 VSUBS 0.00706f
C591 B.n551 VSUBS 0.00706f
C592 B.n552 VSUBS 0.00706f
C593 B.n553 VSUBS 0.00706f
C594 B.n554 VSUBS 0.00706f
C595 B.n555 VSUBS 0.00706f
C596 B.n556 VSUBS 0.00706f
C597 B.n557 VSUBS 0.00706f
C598 B.n558 VSUBS 0.00706f
C599 B.n559 VSUBS 0.00706f
C600 B.n560 VSUBS 0.00706f
C601 B.n561 VSUBS 0.00706f
C602 B.n562 VSUBS 0.00706f
C603 B.n563 VSUBS 0.00706f
C604 B.n564 VSUBS 0.00706f
C605 B.n565 VSUBS 0.00706f
C606 B.n566 VSUBS 0.00706f
C607 B.n567 VSUBS 0.00706f
C608 B.n568 VSUBS 0.00706f
C609 B.n569 VSUBS 0.00706f
C610 B.n570 VSUBS 0.00706f
C611 B.n571 VSUBS 0.00706f
C612 B.n572 VSUBS 0.00706f
C613 B.n573 VSUBS 0.00706f
C614 B.n574 VSUBS 0.00706f
C615 B.n575 VSUBS 0.015987f
C616 VDD1.n0 VSUBS 0.022163f
C617 VDD1.n1 VSUBS 0.021856f
C618 VDD1.n2 VSUBS 0.011744f
C619 VDD1.n3 VSUBS 0.027759f
C620 VDD1.n4 VSUBS 0.012435f
C621 VDD1.n5 VSUBS 0.021856f
C622 VDD1.n6 VSUBS 0.01209f
C623 VDD1.n7 VSUBS 0.027759f
C624 VDD1.n8 VSUBS 0.011744f
C625 VDD1.n9 VSUBS 0.012435f
C626 VDD1.n10 VSUBS 0.021856f
C627 VDD1.n11 VSUBS 0.011744f
C628 VDD1.n12 VSUBS 0.027759f
C629 VDD1.n13 VSUBS 0.012435f
C630 VDD1.n14 VSUBS 0.021856f
C631 VDD1.n15 VSUBS 0.011744f
C632 VDD1.n16 VSUBS 0.02082f
C633 VDD1.n17 VSUBS 0.020882f
C634 VDD1.t3 VSUBS 0.059674f
C635 VDD1.n18 VSUBS 0.151285f
C636 VDD1.n19 VSUBS 0.871765f
C637 VDD1.n20 VSUBS 0.011744f
C638 VDD1.n21 VSUBS 0.012435f
C639 VDD1.n22 VSUBS 0.027759f
C640 VDD1.n23 VSUBS 0.027759f
C641 VDD1.n24 VSUBS 0.012435f
C642 VDD1.n25 VSUBS 0.011744f
C643 VDD1.n26 VSUBS 0.021856f
C644 VDD1.n27 VSUBS 0.021856f
C645 VDD1.n28 VSUBS 0.011744f
C646 VDD1.n29 VSUBS 0.012435f
C647 VDD1.n30 VSUBS 0.027759f
C648 VDD1.n31 VSUBS 0.027759f
C649 VDD1.n32 VSUBS 0.012435f
C650 VDD1.n33 VSUBS 0.011744f
C651 VDD1.n34 VSUBS 0.021856f
C652 VDD1.n35 VSUBS 0.021856f
C653 VDD1.n36 VSUBS 0.011744f
C654 VDD1.n37 VSUBS 0.012435f
C655 VDD1.n38 VSUBS 0.027759f
C656 VDD1.n39 VSUBS 0.027759f
C657 VDD1.n40 VSUBS 0.027759f
C658 VDD1.n41 VSUBS 0.01209f
C659 VDD1.n42 VSUBS 0.011744f
C660 VDD1.n43 VSUBS 0.021856f
C661 VDD1.n44 VSUBS 0.021856f
C662 VDD1.n45 VSUBS 0.011744f
C663 VDD1.n46 VSUBS 0.012435f
C664 VDD1.n47 VSUBS 0.027759f
C665 VDD1.n48 VSUBS 0.060895f
C666 VDD1.n49 VSUBS 0.012435f
C667 VDD1.n50 VSUBS 0.011744f
C668 VDD1.n51 VSUBS 0.048429f
C669 VDD1.n52 VSUBS 0.048739f
C670 VDD1.n53 VSUBS 0.022163f
C671 VDD1.n54 VSUBS 0.021856f
C672 VDD1.n55 VSUBS 0.011744f
C673 VDD1.n56 VSUBS 0.027759f
C674 VDD1.n57 VSUBS 0.012435f
C675 VDD1.n58 VSUBS 0.021856f
C676 VDD1.n59 VSUBS 0.01209f
C677 VDD1.n60 VSUBS 0.027759f
C678 VDD1.n61 VSUBS 0.012435f
C679 VDD1.n62 VSUBS 0.021856f
C680 VDD1.n63 VSUBS 0.011744f
C681 VDD1.n64 VSUBS 0.027759f
C682 VDD1.n65 VSUBS 0.012435f
C683 VDD1.n66 VSUBS 0.021856f
C684 VDD1.n67 VSUBS 0.011744f
C685 VDD1.n68 VSUBS 0.02082f
C686 VDD1.n69 VSUBS 0.020882f
C687 VDD1.t5 VSUBS 0.059674f
C688 VDD1.n70 VSUBS 0.151285f
C689 VDD1.n71 VSUBS 0.871765f
C690 VDD1.n72 VSUBS 0.011744f
C691 VDD1.n73 VSUBS 0.012435f
C692 VDD1.n74 VSUBS 0.027759f
C693 VDD1.n75 VSUBS 0.027759f
C694 VDD1.n76 VSUBS 0.012435f
C695 VDD1.n77 VSUBS 0.011744f
C696 VDD1.n78 VSUBS 0.021856f
C697 VDD1.n79 VSUBS 0.021856f
C698 VDD1.n80 VSUBS 0.011744f
C699 VDD1.n81 VSUBS 0.012435f
C700 VDD1.n82 VSUBS 0.027759f
C701 VDD1.n83 VSUBS 0.027759f
C702 VDD1.n84 VSUBS 0.012435f
C703 VDD1.n85 VSUBS 0.011744f
C704 VDD1.n86 VSUBS 0.021856f
C705 VDD1.n87 VSUBS 0.021856f
C706 VDD1.n88 VSUBS 0.011744f
C707 VDD1.n89 VSUBS 0.011744f
C708 VDD1.n90 VSUBS 0.012435f
C709 VDD1.n91 VSUBS 0.027759f
C710 VDD1.n92 VSUBS 0.027759f
C711 VDD1.n93 VSUBS 0.027759f
C712 VDD1.n94 VSUBS 0.01209f
C713 VDD1.n95 VSUBS 0.011744f
C714 VDD1.n96 VSUBS 0.021856f
C715 VDD1.n97 VSUBS 0.021856f
C716 VDD1.n98 VSUBS 0.011744f
C717 VDD1.n99 VSUBS 0.012435f
C718 VDD1.n100 VSUBS 0.027759f
C719 VDD1.n101 VSUBS 0.060895f
C720 VDD1.n102 VSUBS 0.012435f
C721 VDD1.n103 VSUBS 0.011744f
C722 VDD1.n104 VSUBS 0.048429f
C723 VDD1.n105 VSUBS 0.048266f
C724 VDD1.t2 VSUBS 0.170812f
C725 VDD1.t1 VSUBS 0.170812f
C726 VDD1.n106 VSUBS 1.28567f
C727 VDD1.n107 VSUBS 2.12319f
C728 VDD1.t4 VSUBS 0.170812f
C729 VDD1.t0 VSUBS 0.170812f
C730 VDD1.n108 VSUBS 1.28319f
C731 VDD1.n109 VSUBS 2.24988f
C732 VP.n0 VSUBS 0.042915f
C733 VP.t4 VSUBS 1.75854f
C734 VP.n1 VSUBS 0.054278f
C735 VP.n2 VSUBS 0.042915f
C736 VP.t3 VSUBS 1.75854f
C737 VP.n3 VSUBS 0.07102f
C738 VP.n4 VSUBS 0.042915f
C739 VP.t5 VSUBS 1.75854f
C740 VP.n5 VSUBS 0.054278f
C741 VP.t2 VSUBS 1.89439f
C742 VP.n6 VSUBS 0.749972f
C743 VP.t1 VSUBS 1.75854f
C744 VP.n7 VSUBS 0.726988f
C745 VP.n8 VSUBS 0.060239f
C746 VP.n9 VSUBS 0.269285f
C747 VP.n10 VSUBS 0.042915f
C748 VP.n11 VSUBS 0.042915f
C749 VP.n12 VSUBS 0.07102f
C750 VP.n13 VSUBS 0.049183f
C751 VP.n14 VSUBS 0.727522f
C752 VP.n15 VSUBS 1.83326f
C753 VP.n16 VSUBS 1.86935f
C754 VP.t0 VSUBS 1.75854f
C755 VP.n17 VSUBS 0.727522f
C756 VP.n18 VSUBS 0.049183f
C757 VP.n19 VSUBS 0.042915f
C758 VP.n20 VSUBS 0.042915f
C759 VP.n21 VSUBS 0.042915f
C760 VP.n22 VSUBS 0.054278f
C761 VP.n23 VSUBS 0.060239f
C762 VP.n24 VSUBS 0.646113f
C763 VP.n25 VSUBS 0.060239f
C764 VP.n26 VSUBS 0.042915f
C765 VP.n27 VSUBS 0.042915f
C766 VP.n28 VSUBS 0.042915f
C767 VP.n29 VSUBS 0.07102f
C768 VP.n30 VSUBS 0.049183f
C769 VP.n31 VSUBS 0.727522f
C770 VP.n32 VSUBS 0.04289f
C771 VDD2.n0 VSUBS 0.022128f
C772 VDD2.n1 VSUBS 0.021821f
C773 VDD2.n2 VSUBS 0.011726f
C774 VDD2.n3 VSUBS 0.027715f
C775 VDD2.n4 VSUBS 0.012415f
C776 VDD2.n5 VSUBS 0.021821f
C777 VDD2.n6 VSUBS 0.01207f
C778 VDD2.n7 VSUBS 0.027715f
C779 VDD2.n8 VSUBS 0.012415f
C780 VDD2.n9 VSUBS 0.021821f
C781 VDD2.n10 VSUBS 0.011726f
C782 VDD2.n11 VSUBS 0.027715f
C783 VDD2.n12 VSUBS 0.012415f
C784 VDD2.n13 VSUBS 0.021821f
C785 VDD2.n14 VSUBS 0.011726f
C786 VDD2.n15 VSUBS 0.020786f
C787 VDD2.n16 VSUBS 0.020849f
C788 VDD2.t4 VSUBS 0.059578f
C789 VDD2.n17 VSUBS 0.151043f
C790 VDD2.n18 VSUBS 0.870367f
C791 VDD2.n19 VSUBS 0.011726f
C792 VDD2.n20 VSUBS 0.012415f
C793 VDD2.n21 VSUBS 0.027715f
C794 VDD2.n22 VSUBS 0.027715f
C795 VDD2.n23 VSUBS 0.012415f
C796 VDD2.n24 VSUBS 0.011726f
C797 VDD2.n25 VSUBS 0.021821f
C798 VDD2.n26 VSUBS 0.021821f
C799 VDD2.n27 VSUBS 0.011726f
C800 VDD2.n28 VSUBS 0.012415f
C801 VDD2.n29 VSUBS 0.027715f
C802 VDD2.n30 VSUBS 0.027715f
C803 VDD2.n31 VSUBS 0.012415f
C804 VDD2.n32 VSUBS 0.011726f
C805 VDD2.n33 VSUBS 0.021821f
C806 VDD2.n34 VSUBS 0.021821f
C807 VDD2.n35 VSUBS 0.011726f
C808 VDD2.n36 VSUBS 0.011726f
C809 VDD2.n37 VSUBS 0.012415f
C810 VDD2.n38 VSUBS 0.027715f
C811 VDD2.n39 VSUBS 0.027715f
C812 VDD2.n40 VSUBS 0.027715f
C813 VDD2.n41 VSUBS 0.01207f
C814 VDD2.n42 VSUBS 0.011726f
C815 VDD2.n43 VSUBS 0.021821f
C816 VDD2.n44 VSUBS 0.021821f
C817 VDD2.n45 VSUBS 0.011726f
C818 VDD2.n46 VSUBS 0.012415f
C819 VDD2.n47 VSUBS 0.027715f
C820 VDD2.n48 VSUBS 0.060798f
C821 VDD2.n49 VSUBS 0.012415f
C822 VDD2.n50 VSUBS 0.011726f
C823 VDD2.n51 VSUBS 0.048351f
C824 VDD2.n52 VSUBS 0.048189f
C825 VDD2.t1 VSUBS 0.170538f
C826 VDD2.t0 VSUBS 0.170538f
C827 VDD2.n53 VSUBS 1.2836f
C828 VDD2.n54 VSUBS 2.03623f
C829 VDD2.n55 VSUBS 0.022128f
C830 VDD2.n56 VSUBS 0.021821f
C831 VDD2.n57 VSUBS 0.011726f
C832 VDD2.n58 VSUBS 0.027715f
C833 VDD2.n59 VSUBS 0.012415f
C834 VDD2.n60 VSUBS 0.021821f
C835 VDD2.n61 VSUBS 0.01207f
C836 VDD2.n62 VSUBS 0.027715f
C837 VDD2.n63 VSUBS 0.011726f
C838 VDD2.n64 VSUBS 0.012415f
C839 VDD2.n65 VSUBS 0.021821f
C840 VDD2.n66 VSUBS 0.011726f
C841 VDD2.n67 VSUBS 0.027715f
C842 VDD2.n68 VSUBS 0.012415f
C843 VDD2.n69 VSUBS 0.021821f
C844 VDD2.n70 VSUBS 0.011726f
C845 VDD2.n71 VSUBS 0.020786f
C846 VDD2.n72 VSUBS 0.020849f
C847 VDD2.t5 VSUBS 0.059578f
C848 VDD2.n73 VSUBS 0.151043f
C849 VDD2.n74 VSUBS 0.870367f
C850 VDD2.n75 VSUBS 0.011726f
C851 VDD2.n76 VSUBS 0.012415f
C852 VDD2.n77 VSUBS 0.027715f
C853 VDD2.n78 VSUBS 0.027715f
C854 VDD2.n79 VSUBS 0.012415f
C855 VDD2.n80 VSUBS 0.011726f
C856 VDD2.n81 VSUBS 0.021821f
C857 VDD2.n82 VSUBS 0.021821f
C858 VDD2.n83 VSUBS 0.011726f
C859 VDD2.n84 VSUBS 0.012415f
C860 VDD2.n85 VSUBS 0.027715f
C861 VDD2.n86 VSUBS 0.027715f
C862 VDD2.n87 VSUBS 0.012415f
C863 VDD2.n88 VSUBS 0.011726f
C864 VDD2.n89 VSUBS 0.021821f
C865 VDD2.n90 VSUBS 0.021821f
C866 VDD2.n91 VSUBS 0.011726f
C867 VDD2.n92 VSUBS 0.012415f
C868 VDD2.n93 VSUBS 0.027715f
C869 VDD2.n94 VSUBS 0.027715f
C870 VDD2.n95 VSUBS 0.027715f
C871 VDD2.n96 VSUBS 0.01207f
C872 VDD2.n97 VSUBS 0.011726f
C873 VDD2.n98 VSUBS 0.021821f
C874 VDD2.n99 VSUBS 0.021821f
C875 VDD2.n100 VSUBS 0.011726f
C876 VDD2.n101 VSUBS 0.012415f
C877 VDD2.n102 VSUBS 0.027715f
C878 VDD2.n103 VSUBS 0.060798f
C879 VDD2.n104 VSUBS 0.012415f
C880 VDD2.n105 VSUBS 0.011726f
C881 VDD2.n106 VSUBS 0.048351f
C882 VDD2.n107 VSUBS 0.045314f
C883 VDD2.n108 VSUBS 1.83599f
C884 VDD2.t3 VSUBS 0.170538f
C885 VDD2.t2 VSUBS 0.170538f
C886 VDD2.n109 VSUBS 1.28358f
C887 VTAIL.t11 VSUBS 0.227823f
C888 VTAIL.t9 VSUBS 0.227823f
C889 VTAIL.n0 VSUBS 1.56329f
C890 VTAIL.n1 VSUBS 0.801582f
C891 VTAIL.n2 VSUBS 0.029561f
C892 VTAIL.n3 VSUBS 0.029151f
C893 VTAIL.n4 VSUBS 0.015664f
C894 VTAIL.n5 VSUBS 0.037025f
C895 VTAIL.n6 VSUBS 0.016586f
C896 VTAIL.n7 VSUBS 0.029151f
C897 VTAIL.n8 VSUBS 0.016125f
C898 VTAIL.n9 VSUBS 0.037025f
C899 VTAIL.n10 VSUBS 0.016586f
C900 VTAIL.n11 VSUBS 0.029151f
C901 VTAIL.n12 VSUBS 0.015664f
C902 VTAIL.n13 VSUBS 0.037025f
C903 VTAIL.n14 VSUBS 0.016586f
C904 VTAIL.n15 VSUBS 0.029151f
C905 VTAIL.n16 VSUBS 0.015664f
C906 VTAIL.n17 VSUBS 0.027768f
C907 VTAIL.n18 VSUBS 0.027852f
C908 VTAIL.t4 VSUBS 0.07959f
C909 VTAIL.n19 VSUBS 0.201779f
C910 VTAIL.n20 VSUBS 1.16273f
C911 VTAIL.n21 VSUBS 0.015664f
C912 VTAIL.n22 VSUBS 0.016586f
C913 VTAIL.n23 VSUBS 0.037025f
C914 VTAIL.n24 VSUBS 0.037025f
C915 VTAIL.n25 VSUBS 0.016586f
C916 VTAIL.n26 VSUBS 0.015664f
C917 VTAIL.n27 VSUBS 0.029151f
C918 VTAIL.n28 VSUBS 0.029151f
C919 VTAIL.n29 VSUBS 0.015664f
C920 VTAIL.n30 VSUBS 0.016586f
C921 VTAIL.n31 VSUBS 0.037025f
C922 VTAIL.n32 VSUBS 0.037025f
C923 VTAIL.n33 VSUBS 0.016586f
C924 VTAIL.n34 VSUBS 0.015664f
C925 VTAIL.n35 VSUBS 0.029151f
C926 VTAIL.n36 VSUBS 0.029151f
C927 VTAIL.n37 VSUBS 0.015664f
C928 VTAIL.n38 VSUBS 0.015664f
C929 VTAIL.n39 VSUBS 0.016586f
C930 VTAIL.n40 VSUBS 0.037025f
C931 VTAIL.n41 VSUBS 0.037025f
C932 VTAIL.n42 VSUBS 0.037025f
C933 VTAIL.n43 VSUBS 0.016125f
C934 VTAIL.n44 VSUBS 0.015664f
C935 VTAIL.n45 VSUBS 0.029151f
C936 VTAIL.n46 VSUBS 0.029151f
C937 VTAIL.n47 VSUBS 0.015664f
C938 VTAIL.n48 VSUBS 0.016586f
C939 VTAIL.n49 VSUBS 0.037025f
C940 VTAIL.n50 VSUBS 0.08122f
C941 VTAIL.n51 VSUBS 0.016586f
C942 VTAIL.n52 VSUBS 0.015664f
C943 VTAIL.n53 VSUBS 0.064592f
C944 VTAIL.n54 VSUBS 0.040384f
C945 VTAIL.n55 VSUBS 0.293373f
C946 VTAIL.t5 VSUBS 0.227823f
C947 VTAIL.t3 VSUBS 0.227823f
C948 VTAIL.n56 VSUBS 1.56329f
C949 VTAIL.n57 VSUBS 2.28767f
C950 VTAIL.t8 VSUBS 0.227823f
C951 VTAIL.t7 VSUBS 0.227823f
C952 VTAIL.n58 VSUBS 1.5633f
C953 VTAIL.n59 VSUBS 2.28766f
C954 VTAIL.n60 VSUBS 0.029561f
C955 VTAIL.n61 VSUBS 0.029151f
C956 VTAIL.n62 VSUBS 0.015664f
C957 VTAIL.n63 VSUBS 0.037025f
C958 VTAIL.n64 VSUBS 0.016586f
C959 VTAIL.n65 VSUBS 0.029151f
C960 VTAIL.n66 VSUBS 0.016125f
C961 VTAIL.n67 VSUBS 0.037025f
C962 VTAIL.n68 VSUBS 0.015664f
C963 VTAIL.n69 VSUBS 0.016586f
C964 VTAIL.n70 VSUBS 0.029151f
C965 VTAIL.n71 VSUBS 0.015664f
C966 VTAIL.n72 VSUBS 0.037025f
C967 VTAIL.n73 VSUBS 0.016586f
C968 VTAIL.n74 VSUBS 0.029151f
C969 VTAIL.n75 VSUBS 0.015664f
C970 VTAIL.n76 VSUBS 0.027768f
C971 VTAIL.n77 VSUBS 0.027852f
C972 VTAIL.t6 VSUBS 0.07959f
C973 VTAIL.n78 VSUBS 0.201779f
C974 VTAIL.n79 VSUBS 1.16273f
C975 VTAIL.n80 VSUBS 0.015664f
C976 VTAIL.n81 VSUBS 0.016586f
C977 VTAIL.n82 VSUBS 0.037025f
C978 VTAIL.n83 VSUBS 0.037025f
C979 VTAIL.n84 VSUBS 0.016586f
C980 VTAIL.n85 VSUBS 0.015664f
C981 VTAIL.n86 VSUBS 0.029151f
C982 VTAIL.n87 VSUBS 0.029151f
C983 VTAIL.n88 VSUBS 0.015664f
C984 VTAIL.n89 VSUBS 0.016586f
C985 VTAIL.n90 VSUBS 0.037025f
C986 VTAIL.n91 VSUBS 0.037025f
C987 VTAIL.n92 VSUBS 0.016586f
C988 VTAIL.n93 VSUBS 0.015664f
C989 VTAIL.n94 VSUBS 0.029151f
C990 VTAIL.n95 VSUBS 0.029151f
C991 VTAIL.n96 VSUBS 0.015664f
C992 VTAIL.n97 VSUBS 0.016586f
C993 VTAIL.n98 VSUBS 0.037025f
C994 VTAIL.n99 VSUBS 0.037025f
C995 VTAIL.n100 VSUBS 0.037025f
C996 VTAIL.n101 VSUBS 0.016125f
C997 VTAIL.n102 VSUBS 0.015664f
C998 VTAIL.n103 VSUBS 0.029151f
C999 VTAIL.n104 VSUBS 0.029151f
C1000 VTAIL.n105 VSUBS 0.015664f
C1001 VTAIL.n106 VSUBS 0.016586f
C1002 VTAIL.n107 VSUBS 0.037025f
C1003 VTAIL.n108 VSUBS 0.08122f
C1004 VTAIL.n109 VSUBS 0.016586f
C1005 VTAIL.n110 VSUBS 0.015664f
C1006 VTAIL.n111 VSUBS 0.064592f
C1007 VTAIL.n112 VSUBS 0.040384f
C1008 VTAIL.n113 VSUBS 0.293373f
C1009 VTAIL.t0 VSUBS 0.227823f
C1010 VTAIL.t2 VSUBS 0.227823f
C1011 VTAIL.n114 VSUBS 1.5633f
C1012 VTAIL.n115 VSUBS 0.909063f
C1013 VTAIL.n116 VSUBS 0.029561f
C1014 VTAIL.n117 VSUBS 0.029151f
C1015 VTAIL.n118 VSUBS 0.015664f
C1016 VTAIL.n119 VSUBS 0.037025f
C1017 VTAIL.n120 VSUBS 0.016586f
C1018 VTAIL.n121 VSUBS 0.029151f
C1019 VTAIL.n122 VSUBS 0.016125f
C1020 VTAIL.n123 VSUBS 0.037025f
C1021 VTAIL.n124 VSUBS 0.015664f
C1022 VTAIL.n125 VSUBS 0.016586f
C1023 VTAIL.n126 VSUBS 0.029151f
C1024 VTAIL.n127 VSUBS 0.015664f
C1025 VTAIL.n128 VSUBS 0.037025f
C1026 VTAIL.n129 VSUBS 0.016586f
C1027 VTAIL.n130 VSUBS 0.029151f
C1028 VTAIL.n131 VSUBS 0.015664f
C1029 VTAIL.n132 VSUBS 0.027768f
C1030 VTAIL.n133 VSUBS 0.027852f
C1031 VTAIL.t1 VSUBS 0.07959f
C1032 VTAIL.n134 VSUBS 0.201779f
C1033 VTAIL.n135 VSUBS 1.16273f
C1034 VTAIL.n136 VSUBS 0.015664f
C1035 VTAIL.n137 VSUBS 0.016586f
C1036 VTAIL.n138 VSUBS 0.037025f
C1037 VTAIL.n139 VSUBS 0.037025f
C1038 VTAIL.n140 VSUBS 0.016586f
C1039 VTAIL.n141 VSUBS 0.015664f
C1040 VTAIL.n142 VSUBS 0.029151f
C1041 VTAIL.n143 VSUBS 0.029151f
C1042 VTAIL.n144 VSUBS 0.015664f
C1043 VTAIL.n145 VSUBS 0.016586f
C1044 VTAIL.n146 VSUBS 0.037025f
C1045 VTAIL.n147 VSUBS 0.037025f
C1046 VTAIL.n148 VSUBS 0.016586f
C1047 VTAIL.n149 VSUBS 0.015664f
C1048 VTAIL.n150 VSUBS 0.029151f
C1049 VTAIL.n151 VSUBS 0.029151f
C1050 VTAIL.n152 VSUBS 0.015664f
C1051 VTAIL.n153 VSUBS 0.016586f
C1052 VTAIL.n154 VSUBS 0.037025f
C1053 VTAIL.n155 VSUBS 0.037025f
C1054 VTAIL.n156 VSUBS 0.037025f
C1055 VTAIL.n157 VSUBS 0.016125f
C1056 VTAIL.n158 VSUBS 0.015664f
C1057 VTAIL.n159 VSUBS 0.029151f
C1058 VTAIL.n160 VSUBS 0.029151f
C1059 VTAIL.n161 VSUBS 0.015664f
C1060 VTAIL.n162 VSUBS 0.016586f
C1061 VTAIL.n163 VSUBS 0.037025f
C1062 VTAIL.n164 VSUBS 0.08122f
C1063 VTAIL.n165 VSUBS 0.016586f
C1064 VTAIL.n166 VSUBS 0.015664f
C1065 VTAIL.n167 VSUBS 0.064592f
C1066 VTAIL.n168 VSUBS 0.040384f
C1067 VTAIL.n169 VSUBS 1.52135f
C1068 VTAIL.n170 VSUBS 0.029561f
C1069 VTAIL.n171 VSUBS 0.029151f
C1070 VTAIL.n172 VSUBS 0.015664f
C1071 VTAIL.n173 VSUBS 0.037025f
C1072 VTAIL.n174 VSUBS 0.016586f
C1073 VTAIL.n175 VSUBS 0.029151f
C1074 VTAIL.n176 VSUBS 0.016125f
C1075 VTAIL.n177 VSUBS 0.037025f
C1076 VTAIL.n178 VSUBS 0.016586f
C1077 VTAIL.n179 VSUBS 0.029151f
C1078 VTAIL.n180 VSUBS 0.015664f
C1079 VTAIL.n181 VSUBS 0.037025f
C1080 VTAIL.n182 VSUBS 0.016586f
C1081 VTAIL.n183 VSUBS 0.029151f
C1082 VTAIL.n184 VSUBS 0.015664f
C1083 VTAIL.n185 VSUBS 0.027768f
C1084 VTAIL.n186 VSUBS 0.027852f
C1085 VTAIL.t10 VSUBS 0.07959f
C1086 VTAIL.n187 VSUBS 0.201779f
C1087 VTAIL.n188 VSUBS 1.16273f
C1088 VTAIL.n189 VSUBS 0.015664f
C1089 VTAIL.n190 VSUBS 0.016586f
C1090 VTAIL.n191 VSUBS 0.037025f
C1091 VTAIL.n192 VSUBS 0.037025f
C1092 VTAIL.n193 VSUBS 0.016586f
C1093 VTAIL.n194 VSUBS 0.015664f
C1094 VTAIL.n195 VSUBS 0.029151f
C1095 VTAIL.n196 VSUBS 0.029151f
C1096 VTAIL.n197 VSUBS 0.015664f
C1097 VTAIL.n198 VSUBS 0.016586f
C1098 VTAIL.n199 VSUBS 0.037025f
C1099 VTAIL.n200 VSUBS 0.037025f
C1100 VTAIL.n201 VSUBS 0.016586f
C1101 VTAIL.n202 VSUBS 0.015664f
C1102 VTAIL.n203 VSUBS 0.029151f
C1103 VTAIL.n204 VSUBS 0.029151f
C1104 VTAIL.n205 VSUBS 0.015664f
C1105 VTAIL.n206 VSUBS 0.015664f
C1106 VTAIL.n207 VSUBS 0.016586f
C1107 VTAIL.n208 VSUBS 0.037025f
C1108 VTAIL.n209 VSUBS 0.037025f
C1109 VTAIL.n210 VSUBS 0.037025f
C1110 VTAIL.n211 VSUBS 0.016125f
C1111 VTAIL.n212 VSUBS 0.015664f
C1112 VTAIL.n213 VSUBS 0.029151f
C1113 VTAIL.n214 VSUBS 0.029151f
C1114 VTAIL.n215 VSUBS 0.015664f
C1115 VTAIL.n216 VSUBS 0.016586f
C1116 VTAIL.n217 VSUBS 0.037025f
C1117 VTAIL.n218 VSUBS 0.08122f
C1118 VTAIL.n219 VSUBS 0.016586f
C1119 VTAIL.n220 VSUBS 0.015664f
C1120 VTAIL.n221 VSUBS 0.064592f
C1121 VTAIL.n222 VSUBS 0.040384f
C1122 VTAIL.n223 VSUBS 1.47824f
C1123 VN.n0 VSUBS 0.041729f
C1124 VN.t5 VSUBS 1.7099f
C1125 VN.n1 VSUBS 0.052776f
C1126 VN.t1 VSUBS 1.84199f
C1127 VN.n2 VSUBS 0.72923f
C1128 VN.t4 VSUBS 1.7099f
C1129 VN.n3 VSUBS 0.706882f
C1130 VN.n4 VSUBS 0.058573f
C1131 VN.n5 VSUBS 0.261837f
C1132 VN.n6 VSUBS 0.041729f
C1133 VN.n7 VSUBS 0.041729f
C1134 VN.n8 VSUBS 0.069056f
C1135 VN.n9 VSUBS 0.047822f
C1136 VN.n10 VSUBS 0.707401f
C1137 VN.n11 VSUBS 0.041703f
C1138 VN.n12 VSUBS 0.041729f
C1139 VN.t0 VSUBS 1.7099f
C1140 VN.n13 VSUBS 0.052776f
C1141 VN.t3 VSUBS 1.84199f
C1142 VN.n14 VSUBS 0.72923f
C1143 VN.t2 VSUBS 1.7099f
C1144 VN.n15 VSUBS 0.706882f
C1145 VN.n16 VSUBS 0.058573f
C1146 VN.n17 VSUBS 0.261837f
C1147 VN.n18 VSUBS 0.041729f
C1148 VN.n19 VSUBS 0.041729f
C1149 VN.n20 VSUBS 0.069056f
C1150 VN.n21 VSUBS 0.047822f
C1151 VN.n22 VSUBS 0.707401f
C1152 VN.n23 VSUBS 1.80992f
.ends

