* NGSPICE file created from diff_pair_sample_0985.ext - technology: sky130A

.subckt diff_pair_sample_0985 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=0 ps=0 w=16.13 l=3.42
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=0 ps=0 w=16.13 l=3.42
X2 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=6.2907 ps=33.04 w=16.13 l=3.42
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=6.2907 ps=33.04 w=16.13 l=3.42
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=0 ps=0 w=16.13 l=3.42
X5 VDD2.t0 VN.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=6.2907 ps=33.04 w=16.13 l=3.42
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=0 ps=0 w=16.13 l=3.42
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=6.2907 pd=33.04 as=6.2907 ps=33.04 w=16.13 l=3.42
R0 B.n606 B.n605 585
R1 B.n606 B.n57 585
R2 B.n609 B.n608 585
R3 B.n610 B.n120 585
R4 B.n612 B.n611 585
R5 B.n614 B.n119 585
R6 B.n617 B.n616 585
R7 B.n618 B.n118 585
R8 B.n620 B.n619 585
R9 B.n622 B.n117 585
R10 B.n625 B.n624 585
R11 B.n626 B.n116 585
R12 B.n628 B.n627 585
R13 B.n630 B.n115 585
R14 B.n633 B.n632 585
R15 B.n634 B.n114 585
R16 B.n636 B.n635 585
R17 B.n638 B.n113 585
R18 B.n641 B.n640 585
R19 B.n642 B.n112 585
R20 B.n644 B.n643 585
R21 B.n646 B.n111 585
R22 B.n649 B.n648 585
R23 B.n650 B.n110 585
R24 B.n652 B.n651 585
R25 B.n654 B.n109 585
R26 B.n657 B.n656 585
R27 B.n658 B.n108 585
R28 B.n660 B.n659 585
R29 B.n662 B.n107 585
R30 B.n665 B.n664 585
R31 B.n666 B.n106 585
R32 B.n668 B.n667 585
R33 B.n670 B.n105 585
R34 B.n673 B.n672 585
R35 B.n674 B.n104 585
R36 B.n676 B.n675 585
R37 B.n678 B.n103 585
R38 B.n681 B.n680 585
R39 B.n682 B.n102 585
R40 B.n684 B.n683 585
R41 B.n686 B.n101 585
R42 B.n689 B.n688 585
R43 B.n690 B.n100 585
R44 B.n692 B.n691 585
R45 B.n694 B.n99 585
R46 B.n697 B.n696 585
R47 B.n698 B.n98 585
R48 B.n700 B.n699 585
R49 B.n702 B.n97 585
R50 B.n705 B.n704 585
R51 B.n706 B.n96 585
R52 B.n708 B.n707 585
R53 B.n710 B.n95 585
R54 B.n713 B.n712 585
R55 B.n715 B.n92 585
R56 B.n717 B.n716 585
R57 B.n719 B.n91 585
R58 B.n722 B.n721 585
R59 B.n723 B.n90 585
R60 B.n725 B.n724 585
R61 B.n727 B.n89 585
R62 B.n729 B.n728 585
R63 B.n731 B.n730 585
R64 B.n734 B.n733 585
R65 B.n735 B.n84 585
R66 B.n737 B.n736 585
R67 B.n739 B.n83 585
R68 B.n742 B.n741 585
R69 B.n743 B.n82 585
R70 B.n745 B.n744 585
R71 B.n747 B.n81 585
R72 B.n750 B.n749 585
R73 B.n751 B.n80 585
R74 B.n753 B.n752 585
R75 B.n755 B.n79 585
R76 B.n758 B.n757 585
R77 B.n759 B.n78 585
R78 B.n761 B.n760 585
R79 B.n763 B.n77 585
R80 B.n766 B.n765 585
R81 B.n767 B.n76 585
R82 B.n769 B.n768 585
R83 B.n771 B.n75 585
R84 B.n774 B.n773 585
R85 B.n775 B.n74 585
R86 B.n777 B.n776 585
R87 B.n779 B.n73 585
R88 B.n782 B.n781 585
R89 B.n783 B.n72 585
R90 B.n785 B.n784 585
R91 B.n787 B.n71 585
R92 B.n790 B.n789 585
R93 B.n791 B.n70 585
R94 B.n793 B.n792 585
R95 B.n795 B.n69 585
R96 B.n798 B.n797 585
R97 B.n799 B.n68 585
R98 B.n801 B.n800 585
R99 B.n803 B.n67 585
R100 B.n806 B.n805 585
R101 B.n807 B.n66 585
R102 B.n809 B.n808 585
R103 B.n811 B.n65 585
R104 B.n814 B.n813 585
R105 B.n815 B.n64 585
R106 B.n817 B.n816 585
R107 B.n819 B.n63 585
R108 B.n822 B.n821 585
R109 B.n823 B.n62 585
R110 B.n825 B.n824 585
R111 B.n827 B.n61 585
R112 B.n830 B.n829 585
R113 B.n831 B.n60 585
R114 B.n833 B.n832 585
R115 B.n835 B.n59 585
R116 B.n838 B.n837 585
R117 B.n839 B.n58 585
R118 B.n604 B.n56 585
R119 B.n842 B.n56 585
R120 B.n603 B.n55 585
R121 B.n843 B.n55 585
R122 B.n602 B.n54 585
R123 B.n844 B.n54 585
R124 B.n601 B.n600 585
R125 B.n600 B.n50 585
R126 B.n599 B.n49 585
R127 B.n850 B.n49 585
R128 B.n598 B.n48 585
R129 B.n851 B.n48 585
R130 B.n597 B.n47 585
R131 B.n852 B.n47 585
R132 B.n596 B.n595 585
R133 B.n595 B.n43 585
R134 B.n594 B.n42 585
R135 B.n858 B.n42 585
R136 B.n593 B.n41 585
R137 B.n859 B.n41 585
R138 B.n592 B.n40 585
R139 B.n860 B.n40 585
R140 B.n591 B.n590 585
R141 B.n590 B.n36 585
R142 B.n589 B.n35 585
R143 B.n866 B.n35 585
R144 B.n588 B.n34 585
R145 B.n867 B.n34 585
R146 B.n587 B.n33 585
R147 B.n868 B.n33 585
R148 B.n586 B.n585 585
R149 B.n585 B.n29 585
R150 B.n584 B.n28 585
R151 B.n874 B.n28 585
R152 B.n583 B.n27 585
R153 B.n875 B.n27 585
R154 B.n582 B.n26 585
R155 B.n876 B.n26 585
R156 B.n581 B.n580 585
R157 B.n580 B.n22 585
R158 B.n579 B.n21 585
R159 B.n882 B.n21 585
R160 B.n578 B.n20 585
R161 B.n883 B.n20 585
R162 B.n577 B.n19 585
R163 B.n884 B.n19 585
R164 B.n576 B.n575 585
R165 B.n575 B.n15 585
R166 B.n574 B.n14 585
R167 B.n890 B.n14 585
R168 B.n573 B.n13 585
R169 B.n891 B.n13 585
R170 B.n572 B.n12 585
R171 B.n892 B.n12 585
R172 B.n571 B.n570 585
R173 B.n570 B.n8 585
R174 B.n569 B.n7 585
R175 B.n898 B.n7 585
R176 B.n568 B.n6 585
R177 B.n899 B.n6 585
R178 B.n567 B.n5 585
R179 B.n900 B.n5 585
R180 B.n566 B.n565 585
R181 B.n565 B.n4 585
R182 B.n564 B.n121 585
R183 B.n564 B.n563 585
R184 B.n554 B.n122 585
R185 B.n123 B.n122 585
R186 B.n556 B.n555 585
R187 B.n557 B.n556 585
R188 B.n553 B.n128 585
R189 B.n128 B.n127 585
R190 B.n552 B.n551 585
R191 B.n551 B.n550 585
R192 B.n130 B.n129 585
R193 B.n131 B.n130 585
R194 B.n543 B.n542 585
R195 B.n544 B.n543 585
R196 B.n541 B.n136 585
R197 B.n136 B.n135 585
R198 B.n540 B.n539 585
R199 B.n539 B.n538 585
R200 B.n138 B.n137 585
R201 B.n139 B.n138 585
R202 B.n531 B.n530 585
R203 B.n532 B.n531 585
R204 B.n529 B.n144 585
R205 B.n144 B.n143 585
R206 B.n528 B.n527 585
R207 B.n527 B.n526 585
R208 B.n146 B.n145 585
R209 B.n147 B.n146 585
R210 B.n519 B.n518 585
R211 B.n520 B.n519 585
R212 B.n517 B.n152 585
R213 B.n152 B.n151 585
R214 B.n516 B.n515 585
R215 B.n515 B.n514 585
R216 B.n154 B.n153 585
R217 B.n155 B.n154 585
R218 B.n507 B.n506 585
R219 B.n508 B.n507 585
R220 B.n505 B.n160 585
R221 B.n160 B.n159 585
R222 B.n504 B.n503 585
R223 B.n503 B.n502 585
R224 B.n162 B.n161 585
R225 B.n163 B.n162 585
R226 B.n495 B.n494 585
R227 B.n496 B.n495 585
R228 B.n493 B.n168 585
R229 B.n168 B.n167 585
R230 B.n492 B.n491 585
R231 B.n491 B.n490 585
R232 B.n170 B.n169 585
R233 B.n171 B.n170 585
R234 B.n483 B.n482 585
R235 B.n484 B.n483 585
R236 B.n481 B.n176 585
R237 B.n176 B.n175 585
R238 B.n480 B.n479 585
R239 B.n479 B.n478 585
R240 B.n475 B.n180 585
R241 B.n474 B.n473 585
R242 B.n471 B.n181 585
R243 B.n471 B.n179 585
R244 B.n470 B.n469 585
R245 B.n468 B.n467 585
R246 B.n466 B.n183 585
R247 B.n464 B.n463 585
R248 B.n462 B.n184 585
R249 B.n461 B.n460 585
R250 B.n458 B.n185 585
R251 B.n456 B.n455 585
R252 B.n454 B.n186 585
R253 B.n453 B.n452 585
R254 B.n450 B.n187 585
R255 B.n448 B.n447 585
R256 B.n446 B.n188 585
R257 B.n445 B.n444 585
R258 B.n442 B.n189 585
R259 B.n440 B.n439 585
R260 B.n438 B.n190 585
R261 B.n437 B.n436 585
R262 B.n434 B.n191 585
R263 B.n432 B.n431 585
R264 B.n430 B.n192 585
R265 B.n429 B.n428 585
R266 B.n426 B.n193 585
R267 B.n424 B.n423 585
R268 B.n422 B.n194 585
R269 B.n421 B.n420 585
R270 B.n418 B.n195 585
R271 B.n416 B.n415 585
R272 B.n414 B.n196 585
R273 B.n413 B.n412 585
R274 B.n410 B.n197 585
R275 B.n408 B.n407 585
R276 B.n406 B.n198 585
R277 B.n405 B.n404 585
R278 B.n402 B.n199 585
R279 B.n400 B.n399 585
R280 B.n398 B.n200 585
R281 B.n397 B.n396 585
R282 B.n394 B.n201 585
R283 B.n392 B.n391 585
R284 B.n390 B.n202 585
R285 B.n389 B.n388 585
R286 B.n386 B.n203 585
R287 B.n384 B.n383 585
R288 B.n382 B.n204 585
R289 B.n381 B.n380 585
R290 B.n378 B.n205 585
R291 B.n376 B.n375 585
R292 B.n374 B.n206 585
R293 B.n373 B.n372 585
R294 B.n370 B.n207 585
R295 B.n368 B.n367 585
R296 B.n366 B.n208 585
R297 B.n365 B.n364 585
R298 B.n362 B.n212 585
R299 B.n360 B.n359 585
R300 B.n358 B.n213 585
R301 B.n357 B.n356 585
R302 B.n354 B.n214 585
R303 B.n352 B.n351 585
R304 B.n349 B.n215 585
R305 B.n348 B.n347 585
R306 B.n345 B.n218 585
R307 B.n343 B.n342 585
R308 B.n341 B.n219 585
R309 B.n340 B.n339 585
R310 B.n337 B.n220 585
R311 B.n335 B.n334 585
R312 B.n333 B.n221 585
R313 B.n332 B.n331 585
R314 B.n329 B.n222 585
R315 B.n327 B.n326 585
R316 B.n325 B.n223 585
R317 B.n324 B.n323 585
R318 B.n321 B.n224 585
R319 B.n319 B.n318 585
R320 B.n317 B.n225 585
R321 B.n316 B.n315 585
R322 B.n313 B.n226 585
R323 B.n311 B.n310 585
R324 B.n309 B.n227 585
R325 B.n308 B.n307 585
R326 B.n305 B.n228 585
R327 B.n303 B.n302 585
R328 B.n301 B.n229 585
R329 B.n300 B.n299 585
R330 B.n297 B.n230 585
R331 B.n295 B.n294 585
R332 B.n293 B.n231 585
R333 B.n292 B.n291 585
R334 B.n289 B.n232 585
R335 B.n287 B.n286 585
R336 B.n285 B.n233 585
R337 B.n284 B.n283 585
R338 B.n281 B.n234 585
R339 B.n279 B.n278 585
R340 B.n277 B.n235 585
R341 B.n276 B.n275 585
R342 B.n273 B.n236 585
R343 B.n271 B.n270 585
R344 B.n269 B.n237 585
R345 B.n268 B.n267 585
R346 B.n265 B.n238 585
R347 B.n263 B.n262 585
R348 B.n261 B.n239 585
R349 B.n260 B.n259 585
R350 B.n257 B.n240 585
R351 B.n255 B.n254 585
R352 B.n253 B.n241 585
R353 B.n252 B.n251 585
R354 B.n249 B.n242 585
R355 B.n247 B.n246 585
R356 B.n245 B.n244 585
R357 B.n178 B.n177 585
R358 B.n477 B.n476 585
R359 B.n478 B.n477 585
R360 B.n174 B.n173 585
R361 B.n175 B.n174 585
R362 B.n486 B.n485 585
R363 B.n485 B.n484 585
R364 B.n487 B.n172 585
R365 B.n172 B.n171 585
R366 B.n489 B.n488 585
R367 B.n490 B.n489 585
R368 B.n166 B.n165 585
R369 B.n167 B.n166 585
R370 B.n498 B.n497 585
R371 B.n497 B.n496 585
R372 B.n499 B.n164 585
R373 B.n164 B.n163 585
R374 B.n501 B.n500 585
R375 B.n502 B.n501 585
R376 B.n158 B.n157 585
R377 B.n159 B.n158 585
R378 B.n510 B.n509 585
R379 B.n509 B.n508 585
R380 B.n511 B.n156 585
R381 B.n156 B.n155 585
R382 B.n513 B.n512 585
R383 B.n514 B.n513 585
R384 B.n150 B.n149 585
R385 B.n151 B.n150 585
R386 B.n522 B.n521 585
R387 B.n521 B.n520 585
R388 B.n523 B.n148 585
R389 B.n148 B.n147 585
R390 B.n525 B.n524 585
R391 B.n526 B.n525 585
R392 B.n142 B.n141 585
R393 B.n143 B.n142 585
R394 B.n534 B.n533 585
R395 B.n533 B.n532 585
R396 B.n535 B.n140 585
R397 B.n140 B.n139 585
R398 B.n537 B.n536 585
R399 B.n538 B.n537 585
R400 B.n134 B.n133 585
R401 B.n135 B.n134 585
R402 B.n546 B.n545 585
R403 B.n545 B.n544 585
R404 B.n547 B.n132 585
R405 B.n132 B.n131 585
R406 B.n549 B.n548 585
R407 B.n550 B.n549 585
R408 B.n126 B.n125 585
R409 B.n127 B.n126 585
R410 B.n559 B.n558 585
R411 B.n558 B.n557 585
R412 B.n560 B.n124 585
R413 B.n124 B.n123 585
R414 B.n562 B.n561 585
R415 B.n563 B.n562 585
R416 B.n2 B.n0 585
R417 B.n4 B.n2 585
R418 B.n3 B.n1 585
R419 B.n899 B.n3 585
R420 B.n897 B.n896 585
R421 B.n898 B.n897 585
R422 B.n895 B.n9 585
R423 B.n9 B.n8 585
R424 B.n894 B.n893 585
R425 B.n893 B.n892 585
R426 B.n11 B.n10 585
R427 B.n891 B.n11 585
R428 B.n889 B.n888 585
R429 B.n890 B.n889 585
R430 B.n887 B.n16 585
R431 B.n16 B.n15 585
R432 B.n886 B.n885 585
R433 B.n885 B.n884 585
R434 B.n18 B.n17 585
R435 B.n883 B.n18 585
R436 B.n881 B.n880 585
R437 B.n882 B.n881 585
R438 B.n879 B.n23 585
R439 B.n23 B.n22 585
R440 B.n878 B.n877 585
R441 B.n877 B.n876 585
R442 B.n25 B.n24 585
R443 B.n875 B.n25 585
R444 B.n873 B.n872 585
R445 B.n874 B.n873 585
R446 B.n871 B.n30 585
R447 B.n30 B.n29 585
R448 B.n870 B.n869 585
R449 B.n869 B.n868 585
R450 B.n32 B.n31 585
R451 B.n867 B.n32 585
R452 B.n865 B.n864 585
R453 B.n866 B.n865 585
R454 B.n863 B.n37 585
R455 B.n37 B.n36 585
R456 B.n862 B.n861 585
R457 B.n861 B.n860 585
R458 B.n39 B.n38 585
R459 B.n859 B.n39 585
R460 B.n857 B.n856 585
R461 B.n858 B.n857 585
R462 B.n855 B.n44 585
R463 B.n44 B.n43 585
R464 B.n854 B.n853 585
R465 B.n853 B.n852 585
R466 B.n46 B.n45 585
R467 B.n851 B.n46 585
R468 B.n849 B.n848 585
R469 B.n850 B.n849 585
R470 B.n847 B.n51 585
R471 B.n51 B.n50 585
R472 B.n846 B.n845 585
R473 B.n845 B.n844 585
R474 B.n53 B.n52 585
R475 B.n843 B.n53 585
R476 B.n841 B.n840 585
R477 B.n842 B.n841 585
R478 B.n902 B.n901 585
R479 B.n901 B.n900 585
R480 B.n477 B.n180 535.745
R481 B.n841 B.n58 535.745
R482 B.n479 B.n178 535.745
R483 B.n606 B.n56 535.745
R484 B.n216 B.t12 425.979
R485 B.n209 B.t15 425.979
R486 B.n85 B.t7 425.979
R487 B.n93 B.t4 425.979
R488 B.n217 B.t11 353.252
R489 B.n94 B.t5 353.252
R490 B.n210 B.t14 353.252
R491 B.n86 B.t8 353.252
R492 B.n216 B.t9 322.685
R493 B.n209 B.t13 322.685
R494 B.n85 B.t6 322.685
R495 B.n93 B.t2 322.685
R496 B.n607 B.n57 256.663
R497 B.n613 B.n57 256.663
R498 B.n615 B.n57 256.663
R499 B.n621 B.n57 256.663
R500 B.n623 B.n57 256.663
R501 B.n629 B.n57 256.663
R502 B.n631 B.n57 256.663
R503 B.n637 B.n57 256.663
R504 B.n639 B.n57 256.663
R505 B.n645 B.n57 256.663
R506 B.n647 B.n57 256.663
R507 B.n653 B.n57 256.663
R508 B.n655 B.n57 256.663
R509 B.n661 B.n57 256.663
R510 B.n663 B.n57 256.663
R511 B.n669 B.n57 256.663
R512 B.n671 B.n57 256.663
R513 B.n677 B.n57 256.663
R514 B.n679 B.n57 256.663
R515 B.n685 B.n57 256.663
R516 B.n687 B.n57 256.663
R517 B.n693 B.n57 256.663
R518 B.n695 B.n57 256.663
R519 B.n701 B.n57 256.663
R520 B.n703 B.n57 256.663
R521 B.n709 B.n57 256.663
R522 B.n711 B.n57 256.663
R523 B.n718 B.n57 256.663
R524 B.n720 B.n57 256.663
R525 B.n726 B.n57 256.663
R526 B.n88 B.n57 256.663
R527 B.n732 B.n57 256.663
R528 B.n738 B.n57 256.663
R529 B.n740 B.n57 256.663
R530 B.n746 B.n57 256.663
R531 B.n748 B.n57 256.663
R532 B.n754 B.n57 256.663
R533 B.n756 B.n57 256.663
R534 B.n762 B.n57 256.663
R535 B.n764 B.n57 256.663
R536 B.n770 B.n57 256.663
R537 B.n772 B.n57 256.663
R538 B.n778 B.n57 256.663
R539 B.n780 B.n57 256.663
R540 B.n786 B.n57 256.663
R541 B.n788 B.n57 256.663
R542 B.n794 B.n57 256.663
R543 B.n796 B.n57 256.663
R544 B.n802 B.n57 256.663
R545 B.n804 B.n57 256.663
R546 B.n810 B.n57 256.663
R547 B.n812 B.n57 256.663
R548 B.n818 B.n57 256.663
R549 B.n820 B.n57 256.663
R550 B.n826 B.n57 256.663
R551 B.n828 B.n57 256.663
R552 B.n834 B.n57 256.663
R553 B.n836 B.n57 256.663
R554 B.n472 B.n179 256.663
R555 B.n182 B.n179 256.663
R556 B.n465 B.n179 256.663
R557 B.n459 B.n179 256.663
R558 B.n457 B.n179 256.663
R559 B.n451 B.n179 256.663
R560 B.n449 B.n179 256.663
R561 B.n443 B.n179 256.663
R562 B.n441 B.n179 256.663
R563 B.n435 B.n179 256.663
R564 B.n433 B.n179 256.663
R565 B.n427 B.n179 256.663
R566 B.n425 B.n179 256.663
R567 B.n419 B.n179 256.663
R568 B.n417 B.n179 256.663
R569 B.n411 B.n179 256.663
R570 B.n409 B.n179 256.663
R571 B.n403 B.n179 256.663
R572 B.n401 B.n179 256.663
R573 B.n395 B.n179 256.663
R574 B.n393 B.n179 256.663
R575 B.n387 B.n179 256.663
R576 B.n385 B.n179 256.663
R577 B.n379 B.n179 256.663
R578 B.n377 B.n179 256.663
R579 B.n371 B.n179 256.663
R580 B.n369 B.n179 256.663
R581 B.n363 B.n179 256.663
R582 B.n361 B.n179 256.663
R583 B.n355 B.n179 256.663
R584 B.n353 B.n179 256.663
R585 B.n346 B.n179 256.663
R586 B.n344 B.n179 256.663
R587 B.n338 B.n179 256.663
R588 B.n336 B.n179 256.663
R589 B.n330 B.n179 256.663
R590 B.n328 B.n179 256.663
R591 B.n322 B.n179 256.663
R592 B.n320 B.n179 256.663
R593 B.n314 B.n179 256.663
R594 B.n312 B.n179 256.663
R595 B.n306 B.n179 256.663
R596 B.n304 B.n179 256.663
R597 B.n298 B.n179 256.663
R598 B.n296 B.n179 256.663
R599 B.n290 B.n179 256.663
R600 B.n288 B.n179 256.663
R601 B.n282 B.n179 256.663
R602 B.n280 B.n179 256.663
R603 B.n274 B.n179 256.663
R604 B.n272 B.n179 256.663
R605 B.n266 B.n179 256.663
R606 B.n264 B.n179 256.663
R607 B.n258 B.n179 256.663
R608 B.n256 B.n179 256.663
R609 B.n250 B.n179 256.663
R610 B.n248 B.n179 256.663
R611 B.n243 B.n179 256.663
R612 B.n477 B.n174 163.367
R613 B.n485 B.n174 163.367
R614 B.n485 B.n172 163.367
R615 B.n489 B.n172 163.367
R616 B.n489 B.n166 163.367
R617 B.n497 B.n166 163.367
R618 B.n497 B.n164 163.367
R619 B.n501 B.n164 163.367
R620 B.n501 B.n158 163.367
R621 B.n509 B.n158 163.367
R622 B.n509 B.n156 163.367
R623 B.n513 B.n156 163.367
R624 B.n513 B.n150 163.367
R625 B.n521 B.n150 163.367
R626 B.n521 B.n148 163.367
R627 B.n525 B.n148 163.367
R628 B.n525 B.n142 163.367
R629 B.n533 B.n142 163.367
R630 B.n533 B.n140 163.367
R631 B.n537 B.n140 163.367
R632 B.n537 B.n134 163.367
R633 B.n545 B.n134 163.367
R634 B.n545 B.n132 163.367
R635 B.n549 B.n132 163.367
R636 B.n549 B.n126 163.367
R637 B.n558 B.n126 163.367
R638 B.n558 B.n124 163.367
R639 B.n562 B.n124 163.367
R640 B.n562 B.n2 163.367
R641 B.n901 B.n2 163.367
R642 B.n901 B.n3 163.367
R643 B.n897 B.n3 163.367
R644 B.n897 B.n9 163.367
R645 B.n893 B.n9 163.367
R646 B.n893 B.n11 163.367
R647 B.n889 B.n11 163.367
R648 B.n889 B.n16 163.367
R649 B.n885 B.n16 163.367
R650 B.n885 B.n18 163.367
R651 B.n881 B.n18 163.367
R652 B.n881 B.n23 163.367
R653 B.n877 B.n23 163.367
R654 B.n877 B.n25 163.367
R655 B.n873 B.n25 163.367
R656 B.n873 B.n30 163.367
R657 B.n869 B.n30 163.367
R658 B.n869 B.n32 163.367
R659 B.n865 B.n32 163.367
R660 B.n865 B.n37 163.367
R661 B.n861 B.n37 163.367
R662 B.n861 B.n39 163.367
R663 B.n857 B.n39 163.367
R664 B.n857 B.n44 163.367
R665 B.n853 B.n44 163.367
R666 B.n853 B.n46 163.367
R667 B.n849 B.n46 163.367
R668 B.n849 B.n51 163.367
R669 B.n845 B.n51 163.367
R670 B.n845 B.n53 163.367
R671 B.n841 B.n53 163.367
R672 B.n473 B.n471 163.367
R673 B.n471 B.n470 163.367
R674 B.n467 B.n466 163.367
R675 B.n464 B.n184 163.367
R676 B.n460 B.n458 163.367
R677 B.n456 B.n186 163.367
R678 B.n452 B.n450 163.367
R679 B.n448 B.n188 163.367
R680 B.n444 B.n442 163.367
R681 B.n440 B.n190 163.367
R682 B.n436 B.n434 163.367
R683 B.n432 B.n192 163.367
R684 B.n428 B.n426 163.367
R685 B.n424 B.n194 163.367
R686 B.n420 B.n418 163.367
R687 B.n416 B.n196 163.367
R688 B.n412 B.n410 163.367
R689 B.n408 B.n198 163.367
R690 B.n404 B.n402 163.367
R691 B.n400 B.n200 163.367
R692 B.n396 B.n394 163.367
R693 B.n392 B.n202 163.367
R694 B.n388 B.n386 163.367
R695 B.n384 B.n204 163.367
R696 B.n380 B.n378 163.367
R697 B.n376 B.n206 163.367
R698 B.n372 B.n370 163.367
R699 B.n368 B.n208 163.367
R700 B.n364 B.n362 163.367
R701 B.n360 B.n213 163.367
R702 B.n356 B.n354 163.367
R703 B.n352 B.n215 163.367
R704 B.n347 B.n345 163.367
R705 B.n343 B.n219 163.367
R706 B.n339 B.n337 163.367
R707 B.n335 B.n221 163.367
R708 B.n331 B.n329 163.367
R709 B.n327 B.n223 163.367
R710 B.n323 B.n321 163.367
R711 B.n319 B.n225 163.367
R712 B.n315 B.n313 163.367
R713 B.n311 B.n227 163.367
R714 B.n307 B.n305 163.367
R715 B.n303 B.n229 163.367
R716 B.n299 B.n297 163.367
R717 B.n295 B.n231 163.367
R718 B.n291 B.n289 163.367
R719 B.n287 B.n233 163.367
R720 B.n283 B.n281 163.367
R721 B.n279 B.n235 163.367
R722 B.n275 B.n273 163.367
R723 B.n271 B.n237 163.367
R724 B.n267 B.n265 163.367
R725 B.n263 B.n239 163.367
R726 B.n259 B.n257 163.367
R727 B.n255 B.n241 163.367
R728 B.n251 B.n249 163.367
R729 B.n247 B.n244 163.367
R730 B.n479 B.n176 163.367
R731 B.n483 B.n176 163.367
R732 B.n483 B.n170 163.367
R733 B.n491 B.n170 163.367
R734 B.n491 B.n168 163.367
R735 B.n495 B.n168 163.367
R736 B.n495 B.n162 163.367
R737 B.n503 B.n162 163.367
R738 B.n503 B.n160 163.367
R739 B.n507 B.n160 163.367
R740 B.n507 B.n154 163.367
R741 B.n515 B.n154 163.367
R742 B.n515 B.n152 163.367
R743 B.n519 B.n152 163.367
R744 B.n519 B.n146 163.367
R745 B.n527 B.n146 163.367
R746 B.n527 B.n144 163.367
R747 B.n531 B.n144 163.367
R748 B.n531 B.n138 163.367
R749 B.n539 B.n138 163.367
R750 B.n539 B.n136 163.367
R751 B.n543 B.n136 163.367
R752 B.n543 B.n130 163.367
R753 B.n551 B.n130 163.367
R754 B.n551 B.n128 163.367
R755 B.n556 B.n128 163.367
R756 B.n556 B.n122 163.367
R757 B.n564 B.n122 163.367
R758 B.n565 B.n564 163.367
R759 B.n565 B.n5 163.367
R760 B.n6 B.n5 163.367
R761 B.n7 B.n6 163.367
R762 B.n570 B.n7 163.367
R763 B.n570 B.n12 163.367
R764 B.n13 B.n12 163.367
R765 B.n14 B.n13 163.367
R766 B.n575 B.n14 163.367
R767 B.n575 B.n19 163.367
R768 B.n20 B.n19 163.367
R769 B.n21 B.n20 163.367
R770 B.n580 B.n21 163.367
R771 B.n580 B.n26 163.367
R772 B.n27 B.n26 163.367
R773 B.n28 B.n27 163.367
R774 B.n585 B.n28 163.367
R775 B.n585 B.n33 163.367
R776 B.n34 B.n33 163.367
R777 B.n35 B.n34 163.367
R778 B.n590 B.n35 163.367
R779 B.n590 B.n40 163.367
R780 B.n41 B.n40 163.367
R781 B.n42 B.n41 163.367
R782 B.n595 B.n42 163.367
R783 B.n595 B.n47 163.367
R784 B.n48 B.n47 163.367
R785 B.n49 B.n48 163.367
R786 B.n600 B.n49 163.367
R787 B.n600 B.n54 163.367
R788 B.n55 B.n54 163.367
R789 B.n56 B.n55 163.367
R790 B.n837 B.n835 163.367
R791 B.n833 B.n60 163.367
R792 B.n829 B.n827 163.367
R793 B.n825 B.n62 163.367
R794 B.n821 B.n819 163.367
R795 B.n817 B.n64 163.367
R796 B.n813 B.n811 163.367
R797 B.n809 B.n66 163.367
R798 B.n805 B.n803 163.367
R799 B.n801 B.n68 163.367
R800 B.n797 B.n795 163.367
R801 B.n793 B.n70 163.367
R802 B.n789 B.n787 163.367
R803 B.n785 B.n72 163.367
R804 B.n781 B.n779 163.367
R805 B.n777 B.n74 163.367
R806 B.n773 B.n771 163.367
R807 B.n769 B.n76 163.367
R808 B.n765 B.n763 163.367
R809 B.n761 B.n78 163.367
R810 B.n757 B.n755 163.367
R811 B.n753 B.n80 163.367
R812 B.n749 B.n747 163.367
R813 B.n745 B.n82 163.367
R814 B.n741 B.n739 163.367
R815 B.n737 B.n84 163.367
R816 B.n733 B.n731 163.367
R817 B.n728 B.n727 163.367
R818 B.n725 B.n90 163.367
R819 B.n721 B.n719 163.367
R820 B.n717 B.n92 163.367
R821 B.n712 B.n710 163.367
R822 B.n708 B.n96 163.367
R823 B.n704 B.n702 163.367
R824 B.n700 B.n98 163.367
R825 B.n696 B.n694 163.367
R826 B.n692 B.n100 163.367
R827 B.n688 B.n686 163.367
R828 B.n684 B.n102 163.367
R829 B.n680 B.n678 163.367
R830 B.n676 B.n104 163.367
R831 B.n672 B.n670 163.367
R832 B.n668 B.n106 163.367
R833 B.n664 B.n662 163.367
R834 B.n660 B.n108 163.367
R835 B.n656 B.n654 163.367
R836 B.n652 B.n110 163.367
R837 B.n648 B.n646 163.367
R838 B.n644 B.n112 163.367
R839 B.n640 B.n638 163.367
R840 B.n636 B.n114 163.367
R841 B.n632 B.n630 163.367
R842 B.n628 B.n116 163.367
R843 B.n624 B.n622 163.367
R844 B.n620 B.n118 163.367
R845 B.n616 B.n614 163.367
R846 B.n612 B.n120 163.367
R847 B.n608 B.n606 163.367
R848 B.n217 B.n216 72.7278
R849 B.n210 B.n209 72.7278
R850 B.n86 B.n85 72.7278
R851 B.n94 B.n93 72.7278
R852 B.n472 B.n180 71.676
R853 B.n470 B.n182 71.676
R854 B.n466 B.n465 71.676
R855 B.n459 B.n184 71.676
R856 B.n458 B.n457 71.676
R857 B.n451 B.n186 71.676
R858 B.n450 B.n449 71.676
R859 B.n443 B.n188 71.676
R860 B.n442 B.n441 71.676
R861 B.n435 B.n190 71.676
R862 B.n434 B.n433 71.676
R863 B.n427 B.n192 71.676
R864 B.n426 B.n425 71.676
R865 B.n419 B.n194 71.676
R866 B.n418 B.n417 71.676
R867 B.n411 B.n196 71.676
R868 B.n410 B.n409 71.676
R869 B.n403 B.n198 71.676
R870 B.n402 B.n401 71.676
R871 B.n395 B.n200 71.676
R872 B.n394 B.n393 71.676
R873 B.n387 B.n202 71.676
R874 B.n386 B.n385 71.676
R875 B.n379 B.n204 71.676
R876 B.n378 B.n377 71.676
R877 B.n371 B.n206 71.676
R878 B.n370 B.n369 71.676
R879 B.n363 B.n208 71.676
R880 B.n362 B.n361 71.676
R881 B.n355 B.n213 71.676
R882 B.n354 B.n353 71.676
R883 B.n346 B.n215 71.676
R884 B.n345 B.n344 71.676
R885 B.n338 B.n219 71.676
R886 B.n337 B.n336 71.676
R887 B.n330 B.n221 71.676
R888 B.n329 B.n328 71.676
R889 B.n322 B.n223 71.676
R890 B.n321 B.n320 71.676
R891 B.n314 B.n225 71.676
R892 B.n313 B.n312 71.676
R893 B.n306 B.n227 71.676
R894 B.n305 B.n304 71.676
R895 B.n298 B.n229 71.676
R896 B.n297 B.n296 71.676
R897 B.n290 B.n231 71.676
R898 B.n289 B.n288 71.676
R899 B.n282 B.n233 71.676
R900 B.n281 B.n280 71.676
R901 B.n274 B.n235 71.676
R902 B.n273 B.n272 71.676
R903 B.n266 B.n237 71.676
R904 B.n265 B.n264 71.676
R905 B.n258 B.n239 71.676
R906 B.n257 B.n256 71.676
R907 B.n250 B.n241 71.676
R908 B.n249 B.n248 71.676
R909 B.n244 B.n243 71.676
R910 B.n836 B.n58 71.676
R911 B.n835 B.n834 71.676
R912 B.n828 B.n60 71.676
R913 B.n827 B.n826 71.676
R914 B.n820 B.n62 71.676
R915 B.n819 B.n818 71.676
R916 B.n812 B.n64 71.676
R917 B.n811 B.n810 71.676
R918 B.n804 B.n66 71.676
R919 B.n803 B.n802 71.676
R920 B.n796 B.n68 71.676
R921 B.n795 B.n794 71.676
R922 B.n788 B.n70 71.676
R923 B.n787 B.n786 71.676
R924 B.n780 B.n72 71.676
R925 B.n779 B.n778 71.676
R926 B.n772 B.n74 71.676
R927 B.n771 B.n770 71.676
R928 B.n764 B.n76 71.676
R929 B.n763 B.n762 71.676
R930 B.n756 B.n78 71.676
R931 B.n755 B.n754 71.676
R932 B.n748 B.n80 71.676
R933 B.n747 B.n746 71.676
R934 B.n740 B.n82 71.676
R935 B.n739 B.n738 71.676
R936 B.n732 B.n84 71.676
R937 B.n731 B.n88 71.676
R938 B.n727 B.n726 71.676
R939 B.n720 B.n90 71.676
R940 B.n719 B.n718 71.676
R941 B.n711 B.n92 71.676
R942 B.n710 B.n709 71.676
R943 B.n703 B.n96 71.676
R944 B.n702 B.n701 71.676
R945 B.n695 B.n98 71.676
R946 B.n694 B.n693 71.676
R947 B.n687 B.n100 71.676
R948 B.n686 B.n685 71.676
R949 B.n679 B.n102 71.676
R950 B.n678 B.n677 71.676
R951 B.n671 B.n104 71.676
R952 B.n670 B.n669 71.676
R953 B.n663 B.n106 71.676
R954 B.n662 B.n661 71.676
R955 B.n655 B.n108 71.676
R956 B.n654 B.n653 71.676
R957 B.n647 B.n110 71.676
R958 B.n646 B.n645 71.676
R959 B.n639 B.n112 71.676
R960 B.n638 B.n637 71.676
R961 B.n631 B.n114 71.676
R962 B.n630 B.n629 71.676
R963 B.n623 B.n116 71.676
R964 B.n622 B.n621 71.676
R965 B.n615 B.n118 71.676
R966 B.n614 B.n613 71.676
R967 B.n607 B.n120 71.676
R968 B.n608 B.n607 71.676
R969 B.n613 B.n612 71.676
R970 B.n616 B.n615 71.676
R971 B.n621 B.n620 71.676
R972 B.n624 B.n623 71.676
R973 B.n629 B.n628 71.676
R974 B.n632 B.n631 71.676
R975 B.n637 B.n636 71.676
R976 B.n640 B.n639 71.676
R977 B.n645 B.n644 71.676
R978 B.n648 B.n647 71.676
R979 B.n653 B.n652 71.676
R980 B.n656 B.n655 71.676
R981 B.n661 B.n660 71.676
R982 B.n664 B.n663 71.676
R983 B.n669 B.n668 71.676
R984 B.n672 B.n671 71.676
R985 B.n677 B.n676 71.676
R986 B.n680 B.n679 71.676
R987 B.n685 B.n684 71.676
R988 B.n688 B.n687 71.676
R989 B.n693 B.n692 71.676
R990 B.n696 B.n695 71.676
R991 B.n701 B.n700 71.676
R992 B.n704 B.n703 71.676
R993 B.n709 B.n708 71.676
R994 B.n712 B.n711 71.676
R995 B.n718 B.n717 71.676
R996 B.n721 B.n720 71.676
R997 B.n726 B.n725 71.676
R998 B.n728 B.n88 71.676
R999 B.n733 B.n732 71.676
R1000 B.n738 B.n737 71.676
R1001 B.n741 B.n740 71.676
R1002 B.n746 B.n745 71.676
R1003 B.n749 B.n748 71.676
R1004 B.n754 B.n753 71.676
R1005 B.n757 B.n756 71.676
R1006 B.n762 B.n761 71.676
R1007 B.n765 B.n764 71.676
R1008 B.n770 B.n769 71.676
R1009 B.n773 B.n772 71.676
R1010 B.n778 B.n777 71.676
R1011 B.n781 B.n780 71.676
R1012 B.n786 B.n785 71.676
R1013 B.n789 B.n788 71.676
R1014 B.n794 B.n793 71.676
R1015 B.n797 B.n796 71.676
R1016 B.n802 B.n801 71.676
R1017 B.n805 B.n804 71.676
R1018 B.n810 B.n809 71.676
R1019 B.n813 B.n812 71.676
R1020 B.n818 B.n817 71.676
R1021 B.n821 B.n820 71.676
R1022 B.n826 B.n825 71.676
R1023 B.n829 B.n828 71.676
R1024 B.n834 B.n833 71.676
R1025 B.n837 B.n836 71.676
R1026 B.n473 B.n472 71.676
R1027 B.n467 B.n182 71.676
R1028 B.n465 B.n464 71.676
R1029 B.n460 B.n459 71.676
R1030 B.n457 B.n456 71.676
R1031 B.n452 B.n451 71.676
R1032 B.n449 B.n448 71.676
R1033 B.n444 B.n443 71.676
R1034 B.n441 B.n440 71.676
R1035 B.n436 B.n435 71.676
R1036 B.n433 B.n432 71.676
R1037 B.n428 B.n427 71.676
R1038 B.n425 B.n424 71.676
R1039 B.n420 B.n419 71.676
R1040 B.n417 B.n416 71.676
R1041 B.n412 B.n411 71.676
R1042 B.n409 B.n408 71.676
R1043 B.n404 B.n403 71.676
R1044 B.n401 B.n400 71.676
R1045 B.n396 B.n395 71.676
R1046 B.n393 B.n392 71.676
R1047 B.n388 B.n387 71.676
R1048 B.n385 B.n384 71.676
R1049 B.n380 B.n379 71.676
R1050 B.n377 B.n376 71.676
R1051 B.n372 B.n371 71.676
R1052 B.n369 B.n368 71.676
R1053 B.n364 B.n363 71.676
R1054 B.n361 B.n360 71.676
R1055 B.n356 B.n355 71.676
R1056 B.n353 B.n352 71.676
R1057 B.n347 B.n346 71.676
R1058 B.n344 B.n343 71.676
R1059 B.n339 B.n338 71.676
R1060 B.n336 B.n335 71.676
R1061 B.n331 B.n330 71.676
R1062 B.n328 B.n327 71.676
R1063 B.n323 B.n322 71.676
R1064 B.n320 B.n319 71.676
R1065 B.n315 B.n314 71.676
R1066 B.n312 B.n311 71.676
R1067 B.n307 B.n306 71.676
R1068 B.n304 B.n303 71.676
R1069 B.n299 B.n298 71.676
R1070 B.n296 B.n295 71.676
R1071 B.n291 B.n290 71.676
R1072 B.n288 B.n287 71.676
R1073 B.n283 B.n282 71.676
R1074 B.n280 B.n279 71.676
R1075 B.n275 B.n274 71.676
R1076 B.n272 B.n271 71.676
R1077 B.n267 B.n266 71.676
R1078 B.n264 B.n263 71.676
R1079 B.n259 B.n258 71.676
R1080 B.n256 B.n255 71.676
R1081 B.n251 B.n250 71.676
R1082 B.n248 B.n247 71.676
R1083 B.n243 B.n178 71.676
R1084 B.n478 B.n179 69.3768
R1085 B.n842 B.n57 69.3768
R1086 B.n350 B.n217 59.5399
R1087 B.n211 B.n210 59.5399
R1088 B.n87 B.n86 59.5399
R1089 B.n714 B.n94 59.5399
R1090 B.n478 B.n175 34.9456
R1091 B.n484 B.n175 34.9456
R1092 B.n484 B.n171 34.9456
R1093 B.n490 B.n171 34.9456
R1094 B.n490 B.n167 34.9456
R1095 B.n496 B.n167 34.9456
R1096 B.n496 B.n163 34.9456
R1097 B.n502 B.n163 34.9456
R1098 B.n508 B.n159 34.9456
R1099 B.n508 B.n155 34.9456
R1100 B.n514 B.n155 34.9456
R1101 B.n514 B.n151 34.9456
R1102 B.n520 B.n151 34.9456
R1103 B.n520 B.n147 34.9456
R1104 B.n526 B.n147 34.9456
R1105 B.n526 B.n143 34.9456
R1106 B.n532 B.n143 34.9456
R1107 B.n532 B.n139 34.9456
R1108 B.n538 B.n139 34.9456
R1109 B.n538 B.n135 34.9456
R1110 B.n544 B.n135 34.9456
R1111 B.n550 B.n131 34.9456
R1112 B.n550 B.n127 34.9456
R1113 B.n557 B.n127 34.9456
R1114 B.n557 B.n123 34.9456
R1115 B.n563 B.n123 34.9456
R1116 B.n563 B.n4 34.9456
R1117 B.n900 B.n4 34.9456
R1118 B.n900 B.n899 34.9456
R1119 B.n899 B.n898 34.9456
R1120 B.n898 B.n8 34.9456
R1121 B.n892 B.n8 34.9456
R1122 B.n892 B.n891 34.9456
R1123 B.n891 B.n890 34.9456
R1124 B.n890 B.n15 34.9456
R1125 B.n884 B.n883 34.9456
R1126 B.n883 B.n882 34.9456
R1127 B.n882 B.n22 34.9456
R1128 B.n876 B.n22 34.9456
R1129 B.n876 B.n875 34.9456
R1130 B.n875 B.n874 34.9456
R1131 B.n874 B.n29 34.9456
R1132 B.n868 B.n29 34.9456
R1133 B.n868 B.n867 34.9456
R1134 B.n867 B.n866 34.9456
R1135 B.n866 B.n36 34.9456
R1136 B.n860 B.n36 34.9456
R1137 B.n860 B.n859 34.9456
R1138 B.n858 B.n43 34.9456
R1139 B.n852 B.n43 34.9456
R1140 B.n852 B.n851 34.9456
R1141 B.n851 B.n850 34.9456
R1142 B.n850 B.n50 34.9456
R1143 B.n844 B.n50 34.9456
R1144 B.n844 B.n843 34.9456
R1145 B.n843 B.n842 34.9456
R1146 B.n605 B.n604 34.8103
R1147 B.n840 B.n839 34.8103
R1148 B.n480 B.n177 34.8103
R1149 B.n476 B.n475 34.8103
R1150 B.n544 B.t0 30.8344
R1151 B.n884 B.t1 30.8344
R1152 B.n502 B.t10 22.612
R1153 B.t3 B.n858 22.612
R1154 B B.n902 18.0485
R1155 B.t10 B.n159 12.3341
R1156 B.n859 B.t3 12.3341
R1157 B.n839 B.n838 10.6151
R1158 B.n838 B.n59 10.6151
R1159 B.n832 B.n59 10.6151
R1160 B.n832 B.n831 10.6151
R1161 B.n831 B.n830 10.6151
R1162 B.n830 B.n61 10.6151
R1163 B.n824 B.n61 10.6151
R1164 B.n824 B.n823 10.6151
R1165 B.n823 B.n822 10.6151
R1166 B.n822 B.n63 10.6151
R1167 B.n816 B.n63 10.6151
R1168 B.n816 B.n815 10.6151
R1169 B.n815 B.n814 10.6151
R1170 B.n814 B.n65 10.6151
R1171 B.n808 B.n65 10.6151
R1172 B.n808 B.n807 10.6151
R1173 B.n807 B.n806 10.6151
R1174 B.n806 B.n67 10.6151
R1175 B.n800 B.n67 10.6151
R1176 B.n800 B.n799 10.6151
R1177 B.n799 B.n798 10.6151
R1178 B.n798 B.n69 10.6151
R1179 B.n792 B.n69 10.6151
R1180 B.n792 B.n791 10.6151
R1181 B.n791 B.n790 10.6151
R1182 B.n790 B.n71 10.6151
R1183 B.n784 B.n71 10.6151
R1184 B.n784 B.n783 10.6151
R1185 B.n783 B.n782 10.6151
R1186 B.n782 B.n73 10.6151
R1187 B.n776 B.n73 10.6151
R1188 B.n776 B.n775 10.6151
R1189 B.n775 B.n774 10.6151
R1190 B.n774 B.n75 10.6151
R1191 B.n768 B.n75 10.6151
R1192 B.n768 B.n767 10.6151
R1193 B.n767 B.n766 10.6151
R1194 B.n766 B.n77 10.6151
R1195 B.n760 B.n77 10.6151
R1196 B.n760 B.n759 10.6151
R1197 B.n759 B.n758 10.6151
R1198 B.n758 B.n79 10.6151
R1199 B.n752 B.n79 10.6151
R1200 B.n752 B.n751 10.6151
R1201 B.n751 B.n750 10.6151
R1202 B.n750 B.n81 10.6151
R1203 B.n744 B.n81 10.6151
R1204 B.n744 B.n743 10.6151
R1205 B.n743 B.n742 10.6151
R1206 B.n742 B.n83 10.6151
R1207 B.n736 B.n83 10.6151
R1208 B.n736 B.n735 10.6151
R1209 B.n735 B.n734 10.6151
R1210 B.n730 B.n729 10.6151
R1211 B.n729 B.n89 10.6151
R1212 B.n724 B.n89 10.6151
R1213 B.n724 B.n723 10.6151
R1214 B.n723 B.n722 10.6151
R1215 B.n722 B.n91 10.6151
R1216 B.n716 B.n91 10.6151
R1217 B.n716 B.n715 10.6151
R1218 B.n713 B.n95 10.6151
R1219 B.n707 B.n95 10.6151
R1220 B.n707 B.n706 10.6151
R1221 B.n706 B.n705 10.6151
R1222 B.n705 B.n97 10.6151
R1223 B.n699 B.n97 10.6151
R1224 B.n699 B.n698 10.6151
R1225 B.n698 B.n697 10.6151
R1226 B.n697 B.n99 10.6151
R1227 B.n691 B.n99 10.6151
R1228 B.n691 B.n690 10.6151
R1229 B.n690 B.n689 10.6151
R1230 B.n689 B.n101 10.6151
R1231 B.n683 B.n101 10.6151
R1232 B.n683 B.n682 10.6151
R1233 B.n682 B.n681 10.6151
R1234 B.n681 B.n103 10.6151
R1235 B.n675 B.n103 10.6151
R1236 B.n675 B.n674 10.6151
R1237 B.n674 B.n673 10.6151
R1238 B.n673 B.n105 10.6151
R1239 B.n667 B.n105 10.6151
R1240 B.n667 B.n666 10.6151
R1241 B.n666 B.n665 10.6151
R1242 B.n665 B.n107 10.6151
R1243 B.n659 B.n107 10.6151
R1244 B.n659 B.n658 10.6151
R1245 B.n658 B.n657 10.6151
R1246 B.n657 B.n109 10.6151
R1247 B.n651 B.n109 10.6151
R1248 B.n651 B.n650 10.6151
R1249 B.n650 B.n649 10.6151
R1250 B.n649 B.n111 10.6151
R1251 B.n643 B.n111 10.6151
R1252 B.n643 B.n642 10.6151
R1253 B.n642 B.n641 10.6151
R1254 B.n641 B.n113 10.6151
R1255 B.n635 B.n113 10.6151
R1256 B.n635 B.n634 10.6151
R1257 B.n634 B.n633 10.6151
R1258 B.n633 B.n115 10.6151
R1259 B.n627 B.n115 10.6151
R1260 B.n627 B.n626 10.6151
R1261 B.n626 B.n625 10.6151
R1262 B.n625 B.n117 10.6151
R1263 B.n619 B.n117 10.6151
R1264 B.n619 B.n618 10.6151
R1265 B.n618 B.n617 10.6151
R1266 B.n617 B.n119 10.6151
R1267 B.n611 B.n119 10.6151
R1268 B.n611 B.n610 10.6151
R1269 B.n610 B.n609 10.6151
R1270 B.n609 B.n605 10.6151
R1271 B.n481 B.n480 10.6151
R1272 B.n482 B.n481 10.6151
R1273 B.n482 B.n169 10.6151
R1274 B.n492 B.n169 10.6151
R1275 B.n493 B.n492 10.6151
R1276 B.n494 B.n493 10.6151
R1277 B.n494 B.n161 10.6151
R1278 B.n504 B.n161 10.6151
R1279 B.n505 B.n504 10.6151
R1280 B.n506 B.n505 10.6151
R1281 B.n506 B.n153 10.6151
R1282 B.n516 B.n153 10.6151
R1283 B.n517 B.n516 10.6151
R1284 B.n518 B.n517 10.6151
R1285 B.n518 B.n145 10.6151
R1286 B.n528 B.n145 10.6151
R1287 B.n529 B.n528 10.6151
R1288 B.n530 B.n529 10.6151
R1289 B.n530 B.n137 10.6151
R1290 B.n540 B.n137 10.6151
R1291 B.n541 B.n540 10.6151
R1292 B.n542 B.n541 10.6151
R1293 B.n542 B.n129 10.6151
R1294 B.n552 B.n129 10.6151
R1295 B.n553 B.n552 10.6151
R1296 B.n555 B.n553 10.6151
R1297 B.n555 B.n554 10.6151
R1298 B.n554 B.n121 10.6151
R1299 B.n566 B.n121 10.6151
R1300 B.n567 B.n566 10.6151
R1301 B.n568 B.n567 10.6151
R1302 B.n569 B.n568 10.6151
R1303 B.n571 B.n569 10.6151
R1304 B.n572 B.n571 10.6151
R1305 B.n573 B.n572 10.6151
R1306 B.n574 B.n573 10.6151
R1307 B.n576 B.n574 10.6151
R1308 B.n577 B.n576 10.6151
R1309 B.n578 B.n577 10.6151
R1310 B.n579 B.n578 10.6151
R1311 B.n581 B.n579 10.6151
R1312 B.n582 B.n581 10.6151
R1313 B.n583 B.n582 10.6151
R1314 B.n584 B.n583 10.6151
R1315 B.n586 B.n584 10.6151
R1316 B.n587 B.n586 10.6151
R1317 B.n588 B.n587 10.6151
R1318 B.n589 B.n588 10.6151
R1319 B.n591 B.n589 10.6151
R1320 B.n592 B.n591 10.6151
R1321 B.n593 B.n592 10.6151
R1322 B.n594 B.n593 10.6151
R1323 B.n596 B.n594 10.6151
R1324 B.n597 B.n596 10.6151
R1325 B.n598 B.n597 10.6151
R1326 B.n599 B.n598 10.6151
R1327 B.n601 B.n599 10.6151
R1328 B.n602 B.n601 10.6151
R1329 B.n603 B.n602 10.6151
R1330 B.n604 B.n603 10.6151
R1331 B.n475 B.n474 10.6151
R1332 B.n474 B.n181 10.6151
R1333 B.n469 B.n181 10.6151
R1334 B.n469 B.n468 10.6151
R1335 B.n468 B.n183 10.6151
R1336 B.n463 B.n183 10.6151
R1337 B.n463 B.n462 10.6151
R1338 B.n462 B.n461 10.6151
R1339 B.n461 B.n185 10.6151
R1340 B.n455 B.n185 10.6151
R1341 B.n455 B.n454 10.6151
R1342 B.n454 B.n453 10.6151
R1343 B.n453 B.n187 10.6151
R1344 B.n447 B.n187 10.6151
R1345 B.n447 B.n446 10.6151
R1346 B.n446 B.n445 10.6151
R1347 B.n445 B.n189 10.6151
R1348 B.n439 B.n189 10.6151
R1349 B.n439 B.n438 10.6151
R1350 B.n438 B.n437 10.6151
R1351 B.n437 B.n191 10.6151
R1352 B.n431 B.n191 10.6151
R1353 B.n431 B.n430 10.6151
R1354 B.n430 B.n429 10.6151
R1355 B.n429 B.n193 10.6151
R1356 B.n423 B.n193 10.6151
R1357 B.n423 B.n422 10.6151
R1358 B.n422 B.n421 10.6151
R1359 B.n421 B.n195 10.6151
R1360 B.n415 B.n195 10.6151
R1361 B.n415 B.n414 10.6151
R1362 B.n414 B.n413 10.6151
R1363 B.n413 B.n197 10.6151
R1364 B.n407 B.n197 10.6151
R1365 B.n407 B.n406 10.6151
R1366 B.n406 B.n405 10.6151
R1367 B.n405 B.n199 10.6151
R1368 B.n399 B.n199 10.6151
R1369 B.n399 B.n398 10.6151
R1370 B.n398 B.n397 10.6151
R1371 B.n397 B.n201 10.6151
R1372 B.n391 B.n201 10.6151
R1373 B.n391 B.n390 10.6151
R1374 B.n390 B.n389 10.6151
R1375 B.n389 B.n203 10.6151
R1376 B.n383 B.n203 10.6151
R1377 B.n383 B.n382 10.6151
R1378 B.n382 B.n381 10.6151
R1379 B.n381 B.n205 10.6151
R1380 B.n375 B.n205 10.6151
R1381 B.n375 B.n374 10.6151
R1382 B.n374 B.n373 10.6151
R1383 B.n373 B.n207 10.6151
R1384 B.n367 B.n366 10.6151
R1385 B.n366 B.n365 10.6151
R1386 B.n365 B.n212 10.6151
R1387 B.n359 B.n212 10.6151
R1388 B.n359 B.n358 10.6151
R1389 B.n358 B.n357 10.6151
R1390 B.n357 B.n214 10.6151
R1391 B.n351 B.n214 10.6151
R1392 B.n349 B.n348 10.6151
R1393 B.n348 B.n218 10.6151
R1394 B.n342 B.n218 10.6151
R1395 B.n342 B.n341 10.6151
R1396 B.n341 B.n340 10.6151
R1397 B.n340 B.n220 10.6151
R1398 B.n334 B.n220 10.6151
R1399 B.n334 B.n333 10.6151
R1400 B.n333 B.n332 10.6151
R1401 B.n332 B.n222 10.6151
R1402 B.n326 B.n222 10.6151
R1403 B.n326 B.n325 10.6151
R1404 B.n325 B.n324 10.6151
R1405 B.n324 B.n224 10.6151
R1406 B.n318 B.n224 10.6151
R1407 B.n318 B.n317 10.6151
R1408 B.n317 B.n316 10.6151
R1409 B.n316 B.n226 10.6151
R1410 B.n310 B.n226 10.6151
R1411 B.n310 B.n309 10.6151
R1412 B.n309 B.n308 10.6151
R1413 B.n308 B.n228 10.6151
R1414 B.n302 B.n228 10.6151
R1415 B.n302 B.n301 10.6151
R1416 B.n301 B.n300 10.6151
R1417 B.n300 B.n230 10.6151
R1418 B.n294 B.n230 10.6151
R1419 B.n294 B.n293 10.6151
R1420 B.n293 B.n292 10.6151
R1421 B.n292 B.n232 10.6151
R1422 B.n286 B.n232 10.6151
R1423 B.n286 B.n285 10.6151
R1424 B.n285 B.n284 10.6151
R1425 B.n284 B.n234 10.6151
R1426 B.n278 B.n234 10.6151
R1427 B.n278 B.n277 10.6151
R1428 B.n277 B.n276 10.6151
R1429 B.n276 B.n236 10.6151
R1430 B.n270 B.n236 10.6151
R1431 B.n270 B.n269 10.6151
R1432 B.n269 B.n268 10.6151
R1433 B.n268 B.n238 10.6151
R1434 B.n262 B.n238 10.6151
R1435 B.n262 B.n261 10.6151
R1436 B.n261 B.n260 10.6151
R1437 B.n260 B.n240 10.6151
R1438 B.n254 B.n240 10.6151
R1439 B.n254 B.n253 10.6151
R1440 B.n253 B.n252 10.6151
R1441 B.n252 B.n242 10.6151
R1442 B.n246 B.n242 10.6151
R1443 B.n246 B.n245 10.6151
R1444 B.n245 B.n177 10.6151
R1445 B.n476 B.n173 10.6151
R1446 B.n486 B.n173 10.6151
R1447 B.n487 B.n486 10.6151
R1448 B.n488 B.n487 10.6151
R1449 B.n488 B.n165 10.6151
R1450 B.n498 B.n165 10.6151
R1451 B.n499 B.n498 10.6151
R1452 B.n500 B.n499 10.6151
R1453 B.n500 B.n157 10.6151
R1454 B.n510 B.n157 10.6151
R1455 B.n511 B.n510 10.6151
R1456 B.n512 B.n511 10.6151
R1457 B.n512 B.n149 10.6151
R1458 B.n522 B.n149 10.6151
R1459 B.n523 B.n522 10.6151
R1460 B.n524 B.n523 10.6151
R1461 B.n524 B.n141 10.6151
R1462 B.n534 B.n141 10.6151
R1463 B.n535 B.n534 10.6151
R1464 B.n536 B.n535 10.6151
R1465 B.n536 B.n133 10.6151
R1466 B.n546 B.n133 10.6151
R1467 B.n547 B.n546 10.6151
R1468 B.n548 B.n547 10.6151
R1469 B.n548 B.n125 10.6151
R1470 B.n559 B.n125 10.6151
R1471 B.n560 B.n559 10.6151
R1472 B.n561 B.n560 10.6151
R1473 B.n561 B.n0 10.6151
R1474 B.n896 B.n1 10.6151
R1475 B.n896 B.n895 10.6151
R1476 B.n895 B.n894 10.6151
R1477 B.n894 B.n10 10.6151
R1478 B.n888 B.n10 10.6151
R1479 B.n888 B.n887 10.6151
R1480 B.n887 B.n886 10.6151
R1481 B.n886 B.n17 10.6151
R1482 B.n880 B.n17 10.6151
R1483 B.n880 B.n879 10.6151
R1484 B.n879 B.n878 10.6151
R1485 B.n878 B.n24 10.6151
R1486 B.n872 B.n24 10.6151
R1487 B.n872 B.n871 10.6151
R1488 B.n871 B.n870 10.6151
R1489 B.n870 B.n31 10.6151
R1490 B.n864 B.n31 10.6151
R1491 B.n864 B.n863 10.6151
R1492 B.n863 B.n862 10.6151
R1493 B.n862 B.n38 10.6151
R1494 B.n856 B.n38 10.6151
R1495 B.n856 B.n855 10.6151
R1496 B.n855 B.n854 10.6151
R1497 B.n854 B.n45 10.6151
R1498 B.n848 B.n45 10.6151
R1499 B.n848 B.n847 10.6151
R1500 B.n847 B.n846 10.6151
R1501 B.n846 B.n52 10.6151
R1502 B.n840 B.n52 10.6151
R1503 B.n730 B.n87 6.5566
R1504 B.n715 B.n714 6.5566
R1505 B.n367 B.n211 6.5566
R1506 B.n351 B.n350 6.5566
R1507 B.t0 B.n131 4.11169
R1508 B.t1 B.n15 4.11169
R1509 B.n734 B.n87 4.05904
R1510 B.n714 B.n713 4.05904
R1511 B.n211 B.n207 4.05904
R1512 B.n350 B.n349 4.05904
R1513 B.n902 B.n0 2.81026
R1514 B.n902 B.n1 2.81026
R1515 VP.n0 VP.t0 202.412
R1516 VP.n0 VP.t1 152.452
R1517 VP VP.n0 0.52637
R1518 VTAIL.n354 VTAIL.n270 289.615
R1519 VTAIL.n84 VTAIL.n0 289.615
R1520 VTAIL.n264 VTAIL.n180 289.615
R1521 VTAIL.n174 VTAIL.n90 289.615
R1522 VTAIL.n298 VTAIL.n297 185
R1523 VTAIL.n303 VTAIL.n302 185
R1524 VTAIL.n305 VTAIL.n304 185
R1525 VTAIL.n294 VTAIL.n293 185
R1526 VTAIL.n311 VTAIL.n310 185
R1527 VTAIL.n313 VTAIL.n312 185
R1528 VTAIL.n290 VTAIL.n289 185
R1529 VTAIL.n319 VTAIL.n318 185
R1530 VTAIL.n321 VTAIL.n320 185
R1531 VTAIL.n286 VTAIL.n285 185
R1532 VTAIL.n327 VTAIL.n326 185
R1533 VTAIL.n329 VTAIL.n328 185
R1534 VTAIL.n282 VTAIL.n281 185
R1535 VTAIL.n335 VTAIL.n334 185
R1536 VTAIL.n337 VTAIL.n336 185
R1537 VTAIL.n278 VTAIL.n277 185
R1538 VTAIL.n344 VTAIL.n343 185
R1539 VTAIL.n345 VTAIL.n276 185
R1540 VTAIL.n347 VTAIL.n346 185
R1541 VTAIL.n274 VTAIL.n273 185
R1542 VTAIL.n353 VTAIL.n352 185
R1543 VTAIL.n355 VTAIL.n354 185
R1544 VTAIL.n28 VTAIL.n27 185
R1545 VTAIL.n33 VTAIL.n32 185
R1546 VTAIL.n35 VTAIL.n34 185
R1547 VTAIL.n24 VTAIL.n23 185
R1548 VTAIL.n41 VTAIL.n40 185
R1549 VTAIL.n43 VTAIL.n42 185
R1550 VTAIL.n20 VTAIL.n19 185
R1551 VTAIL.n49 VTAIL.n48 185
R1552 VTAIL.n51 VTAIL.n50 185
R1553 VTAIL.n16 VTAIL.n15 185
R1554 VTAIL.n57 VTAIL.n56 185
R1555 VTAIL.n59 VTAIL.n58 185
R1556 VTAIL.n12 VTAIL.n11 185
R1557 VTAIL.n65 VTAIL.n64 185
R1558 VTAIL.n67 VTAIL.n66 185
R1559 VTAIL.n8 VTAIL.n7 185
R1560 VTAIL.n74 VTAIL.n73 185
R1561 VTAIL.n75 VTAIL.n6 185
R1562 VTAIL.n77 VTAIL.n76 185
R1563 VTAIL.n4 VTAIL.n3 185
R1564 VTAIL.n83 VTAIL.n82 185
R1565 VTAIL.n85 VTAIL.n84 185
R1566 VTAIL.n265 VTAIL.n264 185
R1567 VTAIL.n263 VTAIL.n262 185
R1568 VTAIL.n184 VTAIL.n183 185
R1569 VTAIL.n257 VTAIL.n256 185
R1570 VTAIL.n255 VTAIL.n186 185
R1571 VTAIL.n254 VTAIL.n253 185
R1572 VTAIL.n189 VTAIL.n187 185
R1573 VTAIL.n248 VTAIL.n247 185
R1574 VTAIL.n246 VTAIL.n245 185
R1575 VTAIL.n193 VTAIL.n192 185
R1576 VTAIL.n240 VTAIL.n239 185
R1577 VTAIL.n238 VTAIL.n237 185
R1578 VTAIL.n197 VTAIL.n196 185
R1579 VTAIL.n232 VTAIL.n231 185
R1580 VTAIL.n230 VTAIL.n229 185
R1581 VTAIL.n201 VTAIL.n200 185
R1582 VTAIL.n224 VTAIL.n223 185
R1583 VTAIL.n222 VTAIL.n221 185
R1584 VTAIL.n205 VTAIL.n204 185
R1585 VTAIL.n216 VTAIL.n215 185
R1586 VTAIL.n214 VTAIL.n213 185
R1587 VTAIL.n209 VTAIL.n208 185
R1588 VTAIL.n175 VTAIL.n174 185
R1589 VTAIL.n173 VTAIL.n172 185
R1590 VTAIL.n94 VTAIL.n93 185
R1591 VTAIL.n167 VTAIL.n166 185
R1592 VTAIL.n165 VTAIL.n96 185
R1593 VTAIL.n164 VTAIL.n163 185
R1594 VTAIL.n99 VTAIL.n97 185
R1595 VTAIL.n158 VTAIL.n157 185
R1596 VTAIL.n156 VTAIL.n155 185
R1597 VTAIL.n103 VTAIL.n102 185
R1598 VTAIL.n150 VTAIL.n149 185
R1599 VTAIL.n148 VTAIL.n147 185
R1600 VTAIL.n107 VTAIL.n106 185
R1601 VTAIL.n142 VTAIL.n141 185
R1602 VTAIL.n140 VTAIL.n139 185
R1603 VTAIL.n111 VTAIL.n110 185
R1604 VTAIL.n134 VTAIL.n133 185
R1605 VTAIL.n132 VTAIL.n131 185
R1606 VTAIL.n115 VTAIL.n114 185
R1607 VTAIL.n126 VTAIL.n125 185
R1608 VTAIL.n124 VTAIL.n123 185
R1609 VTAIL.n119 VTAIL.n118 185
R1610 VTAIL.n299 VTAIL.t0 147.659
R1611 VTAIL.n29 VTAIL.t3 147.659
R1612 VTAIL.n210 VTAIL.t2 147.659
R1613 VTAIL.n120 VTAIL.t1 147.659
R1614 VTAIL.n303 VTAIL.n297 104.615
R1615 VTAIL.n304 VTAIL.n303 104.615
R1616 VTAIL.n304 VTAIL.n293 104.615
R1617 VTAIL.n311 VTAIL.n293 104.615
R1618 VTAIL.n312 VTAIL.n311 104.615
R1619 VTAIL.n312 VTAIL.n289 104.615
R1620 VTAIL.n319 VTAIL.n289 104.615
R1621 VTAIL.n320 VTAIL.n319 104.615
R1622 VTAIL.n320 VTAIL.n285 104.615
R1623 VTAIL.n327 VTAIL.n285 104.615
R1624 VTAIL.n328 VTAIL.n327 104.615
R1625 VTAIL.n328 VTAIL.n281 104.615
R1626 VTAIL.n335 VTAIL.n281 104.615
R1627 VTAIL.n336 VTAIL.n335 104.615
R1628 VTAIL.n336 VTAIL.n277 104.615
R1629 VTAIL.n344 VTAIL.n277 104.615
R1630 VTAIL.n345 VTAIL.n344 104.615
R1631 VTAIL.n346 VTAIL.n345 104.615
R1632 VTAIL.n346 VTAIL.n273 104.615
R1633 VTAIL.n353 VTAIL.n273 104.615
R1634 VTAIL.n354 VTAIL.n353 104.615
R1635 VTAIL.n33 VTAIL.n27 104.615
R1636 VTAIL.n34 VTAIL.n33 104.615
R1637 VTAIL.n34 VTAIL.n23 104.615
R1638 VTAIL.n41 VTAIL.n23 104.615
R1639 VTAIL.n42 VTAIL.n41 104.615
R1640 VTAIL.n42 VTAIL.n19 104.615
R1641 VTAIL.n49 VTAIL.n19 104.615
R1642 VTAIL.n50 VTAIL.n49 104.615
R1643 VTAIL.n50 VTAIL.n15 104.615
R1644 VTAIL.n57 VTAIL.n15 104.615
R1645 VTAIL.n58 VTAIL.n57 104.615
R1646 VTAIL.n58 VTAIL.n11 104.615
R1647 VTAIL.n65 VTAIL.n11 104.615
R1648 VTAIL.n66 VTAIL.n65 104.615
R1649 VTAIL.n66 VTAIL.n7 104.615
R1650 VTAIL.n74 VTAIL.n7 104.615
R1651 VTAIL.n75 VTAIL.n74 104.615
R1652 VTAIL.n76 VTAIL.n75 104.615
R1653 VTAIL.n76 VTAIL.n3 104.615
R1654 VTAIL.n83 VTAIL.n3 104.615
R1655 VTAIL.n84 VTAIL.n83 104.615
R1656 VTAIL.n264 VTAIL.n263 104.615
R1657 VTAIL.n263 VTAIL.n183 104.615
R1658 VTAIL.n256 VTAIL.n183 104.615
R1659 VTAIL.n256 VTAIL.n255 104.615
R1660 VTAIL.n255 VTAIL.n254 104.615
R1661 VTAIL.n254 VTAIL.n187 104.615
R1662 VTAIL.n247 VTAIL.n187 104.615
R1663 VTAIL.n247 VTAIL.n246 104.615
R1664 VTAIL.n246 VTAIL.n192 104.615
R1665 VTAIL.n239 VTAIL.n192 104.615
R1666 VTAIL.n239 VTAIL.n238 104.615
R1667 VTAIL.n238 VTAIL.n196 104.615
R1668 VTAIL.n231 VTAIL.n196 104.615
R1669 VTAIL.n231 VTAIL.n230 104.615
R1670 VTAIL.n230 VTAIL.n200 104.615
R1671 VTAIL.n223 VTAIL.n200 104.615
R1672 VTAIL.n223 VTAIL.n222 104.615
R1673 VTAIL.n222 VTAIL.n204 104.615
R1674 VTAIL.n215 VTAIL.n204 104.615
R1675 VTAIL.n215 VTAIL.n214 104.615
R1676 VTAIL.n214 VTAIL.n208 104.615
R1677 VTAIL.n174 VTAIL.n173 104.615
R1678 VTAIL.n173 VTAIL.n93 104.615
R1679 VTAIL.n166 VTAIL.n93 104.615
R1680 VTAIL.n166 VTAIL.n165 104.615
R1681 VTAIL.n165 VTAIL.n164 104.615
R1682 VTAIL.n164 VTAIL.n97 104.615
R1683 VTAIL.n157 VTAIL.n97 104.615
R1684 VTAIL.n157 VTAIL.n156 104.615
R1685 VTAIL.n156 VTAIL.n102 104.615
R1686 VTAIL.n149 VTAIL.n102 104.615
R1687 VTAIL.n149 VTAIL.n148 104.615
R1688 VTAIL.n148 VTAIL.n106 104.615
R1689 VTAIL.n141 VTAIL.n106 104.615
R1690 VTAIL.n141 VTAIL.n140 104.615
R1691 VTAIL.n140 VTAIL.n110 104.615
R1692 VTAIL.n133 VTAIL.n110 104.615
R1693 VTAIL.n133 VTAIL.n132 104.615
R1694 VTAIL.n132 VTAIL.n114 104.615
R1695 VTAIL.n125 VTAIL.n114 104.615
R1696 VTAIL.n125 VTAIL.n124 104.615
R1697 VTAIL.n124 VTAIL.n118 104.615
R1698 VTAIL.t0 VTAIL.n297 52.3082
R1699 VTAIL.t3 VTAIL.n27 52.3082
R1700 VTAIL.t2 VTAIL.n208 52.3082
R1701 VTAIL.t1 VTAIL.n118 52.3082
R1702 VTAIL.n359 VTAIL.n358 33.155
R1703 VTAIL.n89 VTAIL.n88 33.155
R1704 VTAIL.n269 VTAIL.n268 33.155
R1705 VTAIL.n179 VTAIL.n178 33.155
R1706 VTAIL.n179 VTAIL.n89 32.7376
R1707 VTAIL.n359 VTAIL.n269 29.5048
R1708 VTAIL.n299 VTAIL.n298 15.6677
R1709 VTAIL.n29 VTAIL.n28 15.6677
R1710 VTAIL.n210 VTAIL.n209 15.6677
R1711 VTAIL.n120 VTAIL.n119 15.6677
R1712 VTAIL.n347 VTAIL.n276 13.1884
R1713 VTAIL.n77 VTAIL.n6 13.1884
R1714 VTAIL.n257 VTAIL.n186 13.1884
R1715 VTAIL.n167 VTAIL.n96 13.1884
R1716 VTAIL.n302 VTAIL.n301 12.8005
R1717 VTAIL.n343 VTAIL.n342 12.8005
R1718 VTAIL.n348 VTAIL.n274 12.8005
R1719 VTAIL.n32 VTAIL.n31 12.8005
R1720 VTAIL.n73 VTAIL.n72 12.8005
R1721 VTAIL.n78 VTAIL.n4 12.8005
R1722 VTAIL.n258 VTAIL.n184 12.8005
R1723 VTAIL.n253 VTAIL.n188 12.8005
R1724 VTAIL.n213 VTAIL.n212 12.8005
R1725 VTAIL.n168 VTAIL.n94 12.8005
R1726 VTAIL.n163 VTAIL.n98 12.8005
R1727 VTAIL.n123 VTAIL.n122 12.8005
R1728 VTAIL.n305 VTAIL.n296 12.0247
R1729 VTAIL.n341 VTAIL.n278 12.0247
R1730 VTAIL.n352 VTAIL.n351 12.0247
R1731 VTAIL.n35 VTAIL.n26 12.0247
R1732 VTAIL.n71 VTAIL.n8 12.0247
R1733 VTAIL.n82 VTAIL.n81 12.0247
R1734 VTAIL.n262 VTAIL.n261 12.0247
R1735 VTAIL.n252 VTAIL.n189 12.0247
R1736 VTAIL.n216 VTAIL.n207 12.0247
R1737 VTAIL.n172 VTAIL.n171 12.0247
R1738 VTAIL.n162 VTAIL.n99 12.0247
R1739 VTAIL.n126 VTAIL.n117 12.0247
R1740 VTAIL.n306 VTAIL.n294 11.249
R1741 VTAIL.n338 VTAIL.n337 11.249
R1742 VTAIL.n355 VTAIL.n272 11.249
R1743 VTAIL.n36 VTAIL.n24 11.249
R1744 VTAIL.n68 VTAIL.n67 11.249
R1745 VTAIL.n85 VTAIL.n2 11.249
R1746 VTAIL.n265 VTAIL.n182 11.249
R1747 VTAIL.n249 VTAIL.n248 11.249
R1748 VTAIL.n217 VTAIL.n205 11.249
R1749 VTAIL.n175 VTAIL.n92 11.249
R1750 VTAIL.n159 VTAIL.n158 11.249
R1751 VTAIL.n127 VTAIL.n115 11.249
R1752 VTAIL.n310 VTAIL.n309 10.4732
R1753 VTAIL.n334 VTAIL.n280 10.4732
R1754 VTAIL.n356 VTAIL.n270 10.4732
R1755 VTAIL.n40 VTAIL.n39 10.4732
R1756 VTAIL.n64 VTAIL.n10 10.4732
R1757 VTAIL.n86 VTAIL.n0 10.4732
R1758 VTAIL.n266 VTAIL.n180 10.4732
R1759 VTAIL.n245 VTAIL.n191 10.4732
R1760 VTAIL.n221 VTAIL.n220 10.4732
R1761 VTAIL.n176 VTAIL.n90 10.4732
R1762 VTAIL.n155 VTAIL.n101 10.4732
R1763 VTAIL.n131 VTAIL.n130 10.4732
R1764 VTAIL.n313 VTAIL.n292 9.69747
R1765 VTAIL.n333 VTAIL.n282 9.69747
R1766 VTAIL.n43 VTAIL.n22 9.69747
R1767 VTAIL.n63 VTAIL.n12 9.69747
R1768 VTAIL.n244 VTAIL.n193 9.69747
R1769 VTAIL.n224 VTAIL.n203 9.69747
R1770 VTAIL.n154 VTAIL.n103 9.69747
R1771 VTAIL.n134 VTAIL.n113 9.69747
R1772 VTAIL.n358 VTAIL.n357 9.45567
R1773 VTAIL.n88 VTAIL.n87 9.45567
R1774 VTAIL.n268 VTAIL.n267 9.45567
R1775 VTAIL.n178 VTAIL.n177 9.45567
R1776 VTAIL.n357 VTAIL.n356 9.3005
R1777 VTAIL.n272 VTAIL.n271 9.3005
R1778 VTAIL.n351 VTAIL.n350 9.3005
R1779 VTAIL.n349 VTAIL.n348 9.3005
R1780 VTAIL.n288 VTAIL.n287 9.3005
R1781 VTAIL.n317 VTAIL.n316 9.3005
R1782 VTAIL.n315 VTAIL.n314 9.3005
R1783 VTAIL.n292 VTAIL.n291 9.3005
R1784 VTAIL.n309 VTAIL.n308 9.3005
R1785 VTAIL.n307 VTAIL.n306 9.3005
R1786 VTAIL.n296 VTAIL.n295 9.3005
R1787 VTAIL.n301 VTAIL.n300 9.3005
R1788 VTAIL.n323 VTAIL.n322 9.3005
R1789 VTAIL.n325 VTAIL.n324 9.3005
R1790 VTAIL.n284 VTAIL.n283 9.3005
R1791 VTAIL.n331 VTAIL.n330 9.3005
R1792 VTAIL.n333 VTAIL.n332 9.3005
R1793 VTAIL.n280 VTAIL.n279 9.3005
R1794 VTAIL.n339 VTAIL.n338 9.3005
R1795 VTAIL.n341 VTAIL.n340 9.3005
R1796 VTAIL.n342 VTAIL.n275 9.3005
R1797 VTAIL.n87 VTAIL.n86 9.3005
R1798 VTAIL.n2 VTAIL.n1 9.3005
R1799 VTAIL.n81 VTAIL.n80 9.3005
R1800 VTAIL.n79 VTAIL.n78 9.3005
R1801 VTAIL.n18 VTAIL.n17 9.3005
R1802 VTAIL.n47 VTAIL.n46 9.3005
R1803 VTAIL.n45 VTAIL.n44 9.3005
R1804 VTAIL.n22 VTAIL.n21 9.3005
R1805 VTAIL.n39 VTAIL.n38 9.3005
R1806 VTAIL.n37 VTAIL.n36 9.3005
R1807 VTAIL.n26 VTAIL.n25 9.3005
R1808 VTAIL.n31 VTAIL.n30 9.3005
R1809 VTAIL.n53 VTAIL.n52 9.3005
R1810 VTAIL.n55 VTAIL.n54 9.3005
R1811 VTAIL.n14 VTAIL.n13 9.3005
R1812 VTAIL.n61 VTAIL.n60 9.3005
R1813 VTAIL.n63 VTAIL.n62 9.3005
R1814 VTAIL.n10 VTAIL.n9 9.3005
R1815 VTAIL.n69 VTAIL.n68 9.3005
R1816 VTAIL.n71 VTAIL.n70 9.3005
R1817 VTAIL.n72 VTAIL.n5 9.3005
R1818 VTAIL.n236 VTAIL.n235 9.3005
R1819 VTAIL.n195 VTAIL.n194 9.3005
R1820 VTAIL.n242 VTAIL.n241 9.3005
R1821 VTAIL.n244 VTAIL.n243 9.3005
R1822 VTAIL.n191 VTAIL.n190 9.3005
R1823 VTAIL.n250 VTAIL.n249 9.3005
R1824 VTAIL.n252 VTAIL.n251 9.3005
R1825 VTAIL.n188 VTAIL.n185 9.3005
R1826 VTAIL.n267 VTAIL.n266 9.3005
R1827 VTAIL.n182 VTAIL.n181 9.3005
R1828 VTAIL.n261 VTAIL.n260 9.3005
R1829 VTAIL.n259 VTAIL.n258 9.3005
R1830 VTAIL.n234 VTAIL.n233 9.3005
R1831 VTAIL.n199 VTAIL.n198 9.3005
R1832 VTAIL.n228 VTAIL.n227 9.3005
R1833 VTAIL.n226 VTAIL.n225 9.3005
R1834 VTAIL.n203 VTAIL.n202 9.3005
R1835 VTAIL.n220 VTAIL.n219 9.3005
R1836 VTAIL.n218 VTAIL.n217 9.3005
R1837 VTAIL.n207 VTAIL.n206 9.3005
R1838 VTAIL.n212 VTAIL.n211 9.3005
R1839 VTAIL.n146 VTAIL.n145 9.3005
R1840 VTAIL.n105 VTAIL.n104 9.3005
R1841 VTAIL.n152 VTAIL.n151 9.3005
R1842 VTAIL.n154 VTAIL.n153 9.3005
R1843 VTAIL.n101 VTAIL.n100 9.3005
R1844 VTAIL.n160 VTAIL.n159 9.3005
R1845 VTAIL.n162 VTAIL.n161 9.3005
R1846 VTAIL.n98 VTAIL.n95 9.3005
R1847 VTAIL.n177 VTAIL.n176 9.3005
R1848 VTAIL.n92 VTAIL.n91 9.3005
R1849 VTAIL.n171 VTAIL.n170 9.3005
R1850 VTAIL.n169 VTAIL.n168 9.3005
R1851 VTAIL.n144 VTAIL.n143 9.3005
R1852 VTAIL.n109 VTAIL.n108 9.3005
R1853 VTAIL.n138 VTAIL.n137 9.3005
R1854 VTAIL.n136 VTAIL.n135 9.3005
R1855 VTAIL.n113 VTAIL.n112 9.3005
R1856 VTAIL.n130 VTAIL.n129 9.3005
R1857 VTAIL.n128 VTAIL.n127 9.3005
R1858 VTAIL.n117 VTAIL.n116 9.3005
R1859 VTAIL.n122 VTAIL.n121 9.3005
R1860 VTAIL.n314 VTAIL.n290 8.92171
R1861 VTAIL.n330 VTAIL.n329 8.92171
R1862 VTAIL.n44 VTAIL.n20 8.92171
R1863 VTAIL.n60 VTAIL.n59 8.92171
R1864 VTAIL.n241 VTAIL.n240 8.92171
R1865 VTAIL.n225 VTAIL.n201 8.92171
R1866 VTAIL.n151 VTAIL.n150 8.92171
R1867 VTAIL.n135 VTAIL.n111 8.92171
R1868 VTAIL.n318 VTAIL.n317 8.14595
R1869 VTAIL.n326 VTAIL.n284 8.14595
R1870 VTAIL.n48 VTAIL.n47 8.14595
R1871 VTAIL.n56 VTAIL.n14 8.14595
R1872 VTAIL.n237 VTAIL.n195 8.14595
R1873 VTAIL.n229 VTAIL.n228 8.14595
R1874 VTAIL.n147 VTAIL.n105 8.14595
R1875 VTAIL.n139 VTAIL.n138 8.14595
R1876 VTAIL.n321 VTAIL.n288 7.3702
R1877 VTAIL.n325 VTAIL.n286 7.3702
R1878 VTAIL.n51 VTAIL.n18 7.3702
R1879 VTAIL.n55 VTAIL.n16 7.3702
R1880 VTAIL.n236 VTAIL.n197 7.3702
R1881 VTAIL.n232 VTAIL.n199 7.3702
R1882 VTAIL.n146 VTAIL.n107 7.3702
R1883 VTAIL.n142 VTAIL.n109 7.3702
R1884 VTAIL.n322 VTAIL.n321 6.59444
R1885 VTAIL.n322 VTAIL.n286 6.59444
R1886 VTAIL.n52 VTAIL.n51 6.59444
R1887 VTAIL.n52 VTAIL.n16 6.59444
R1888 VTAIL.n233 VTAIL.n197 6.59444
R1889 VTAIL.n233 VTAIL.n232 6.59444
R1890 VTAIL.n143 VTAIL.n107 6.59444
R1891 VTAIL.n143 VTAIL.n142 6.59444
R1892 VTAIL.n318 VTAIL.n288 5.81868
R1893 VTAIL.n326 VTAIL.n325 5.81868
R1894 VTAIL.n48 VTAIL.n18 5.81868
R1895 VTAIL.n56 VTAIL.n55 5.81868
R1896 VTAIL.n237 VTAIL.n236 5.81868
R1897 VTAIL.n229 VTAIL.n199 5.81868
R1898 VTAIL.n147 VTAIL.n146 5.81868
R1899 VTAIL.n139 VTAIL.n109 5.81868
R1900 VTAIL.n317 VTAIL.n290 5.04292
R1901 VTAIL.n329 VTAIL.n284 5.04292
R1902 VTAIL.n47 VTAIL.n20 5.04292
R1903 VTAIL.n59 VTAIL.n14 5.04292
R1904 VTAIL.n240 VTAIL.n195 5.04292
R1905 VTAIL.n228 VTAIL.n201 5.04292
R1906 VTAIL.n150 VTAIL.n105 5.04292
R1907 VTAIL.n138 VTAIL.n111 5.04292
R1908 VTAIL.n300 VTAIL.n299 4.38563
R1909 VTAIL.n30 VTAIL.n29 4.38563
R1910 VTAIL.n211 VTAIL.n210 4.38563
R1911 VTAIL.n121 VTAIL.n120 4.38563
R1912 VTAIL.n314 VTAIL.n313 4.26717
R1913 VTAIL.n330 VTAIL.n282 4.26717
R1914 VTAIL.n44 VTAIL.n43 4.26717
R1915 VTAIL.n60 VTAIL.n12 4.26717
R1916 VTAIL.n241 VTAIL.n193 4.26717
R1917 VTAIL.n225 VTAIL.n224 4.26717
R1918 VTAIL.n151 VTAIL.n103 4.26717
R1919 VTAIL.n135 VTAIL.n134 4.26717
R1920 VTAIL.n310 VTAIL.n292 3.49141
R1921 VTAIL.n334 VTAIL.n333 3.49141
R1922 VTAIL.n358 VTAIL.n270 3.49141
R1923 VTAIL.n40 VTAIL.n22 3.49141
R1924 VTAIL.n64 VTAIL.n63 3.49141
R1925 VTAIL.n88 VTAIL.n0 3.49141
R1926 VTAIL.n268 VTAIL.n180 3.49141
R1927 VTAIL.n245 VTAIL.n244 3.49141
R1928 VTAIL.n221 VTAIL.n203 3.49141
R1929 VTAIL.n178 VTAIL.n90 3.49141
R1930 VTAIL.n155 VTAIL.n154 3.49141
R1931 VTAIL.n131 VTAIL.n113 3.49141
R1932 VTAIL.n309 VTAIL.n294 2.71565
R1933 VTAIL.n337 VTAIL.n280 2.71565
R1934 VTAIL.n356 VTAIL.n355 2.71565
R1935 VTAIL.n39 VTAIL.n24 2.71565
R1936 VTAIL.n67 VTAIL.n10 2.71565
R1937 VTAIL.n86 VTAIL.n85 2.71565
R1938 VTAIL.n266 VTAIL.n265 2.71565
R1939 VTAIL.n248 VTAIL.n191 2.71565
R1940 VTAIL.n220 VTAIL.n205 2.71565
R1941 VTAIL.n176 VTAIL.n175 2.71565
R1942 VTAIL.n158 VTAIL.n101 2.71565
R1943 VTAIL.n130 VTAIL.n115 2.71565
R1944 VTAIL.n269 VTAIL.n179 2.08671
R1945 VTAIL.n306 VTAIL.n305 1.93989
R1946 VTAIL.n338 VTAIL.n278 1.93989
R1947 VTAIL.n352 VTAIL.n272 1.93989
R1948 VTAIL.n36 VTAIL.n35 1.93989
R1949 VTAIL.n68 VTAIL.n8 1.93989
R1950 VTAIL.n82 VTAIL.n2 1.93989
R1951 VTAIL.n262 VTAIL.n182 1.93989
R1952 VTAIL.n249 VTAIL.n189 1.93989
R1953 VTAIL.n217 VTAIL.n216 1.93989
R1954 VTAIL.n172 VTAIL.n92 1.93989
R1955 VTAIL.n159 VTAIL.n99 1.93989
R1956 VTAIL.n127 VTAIL.n126 1.93989
R1957 VTAIL VTAIL.n89 1.33671
R1958 VTAIL.n302 VTAIL.n296 1.16414
R1959 VTAIL.n343 VTAIL.n341 1.16414
R1960 VTAIL.n351 VTAIL.n274 1.16414
R1961 VTAIL.n32 VTAIL.n26 1.16414
R1962 VTAIL.n73 VTAIL.n71 1.16414
R1963 VTAIL.n81 VTAIL.n4 1.16414
R1964 VTAIL.n261 VTAIL.n184 1.16414
R1965 VTAIL.n253 VTAIL.n252 1.16414
R1966 VTAIL.n213 VTAIL.n207 1.16414
R1967 VTAIL.n171 VTAIL.n94 1.16414
R1968 VTAIL.n163 VTAIL.n162 1.16414
R1969 VTAIL.n123 VTAIL.n117 1.16414
R1970 VTAIL VTAIL.n359 0.7505
R1971 VTAIL.n301 VTAIL.n298 0.388379
R1972 VTAIL.n342 VTAIL.n276 0.388379
R1973 VTAIL.n348 VTAIL.n347 0.388379
R1974 VTAIL.n31 VTAIL.n28 0.388379
R1975 VTAIL.n72 VTAIL.n6 0.388379
R1976 VTAIL.n78 VTAIL.n77 0.388379
R1977 VTAIL.n258 VTAIL.n257 0.388379
R1978 VTAIL.n188 VTAIL.n186 0.388379
R1979 VTAIL.n212 VTAIL.n209 0.388379
R1980 VTAIL.n168 VTAIL.n167 0.388379
R1981 VTAIL.n98 VTAIL.n96 0.388379
R1982 VTAIL.n122 VTAIL.n119 0.388379
R1983 VTAIL.n300 VTAIL.n295 0.155672
R1984 VTAIL.n307 VTAIL.n295 0.155672
R1985 VTAIL.n308 VTAIL.n307 0.155672
R1986 VTAIL.n308 VTAIL.n291 0.155672
R1987 VTAIL.n315 VTAIL.n291 0.155672
R1988 VTAIL.n316 VTAIL.n315 0.155672
R1989 VTAIL.n316 VTAIL.n287 0.155672
R1990 VTAIL.n323 VTAIL.n287 0.155672
R1991 VTAIL.n324 VTAIL.n323 0.155672
R1992 VTAIL.n324 VTAIL.n283 0.155672
R1993 VTAIL.n331 VTAIL.n283 0.155672
R1994 VTAIL.n332 VTAIL.n331 0.155672
R1995 VTAIL.n332 VTAIL.n279 0.155672
R1996 VTAIL.n339 VTAIL.n279 0.155672
R1997 VTAIL.n340 VTAIL.n339 0.155672
R1998 VTAIL.n340 VTAIL.n275 0.155672
R1999 VTAIL.n349 VTAIL.n275 0.155672
R2000 VTAIL.n350 VTAIL.n349 0.155672
R2001 VTAIL.n350 VTAIL.n271 0.155672
R2002 VTAIL.n357 VTAIL.n271 0.155672
R2003 VTAIL.n30 VTAIL.n25 0.155672
R2004 VTAIL.n37 VTAIL.n25 0.155672
R2005 VTAIL.n38 VTAIL.n37 0.155672
R2006 VTAIL.n38 VTAIL.n21 0.155672
R2007 VTAIL.n45 VTAIL.n21 0.155672
R2008 VTAIL.n46 VTAIL.n45 0.155672
R2009 VTAIL.n46 VTAIL.n17 0.155672
R2010 VTAIL.n53 VTAIL.n17 0.155672
R2011 VTAIL.n54 VTAIL.n53 0.155672
R2012 VTAIL.n54 VTAIL.n13 0.155672
R2013 VTAIL.n61 VTAIL.n13 0.155672
R2014 VTAIL.n62 VTAIL.n61 0.155672
R2015 VTAIL.n62 VTAIL.n9 0.155672
R2016 VTAIL.n69 VTAIL.n9 0.155672
R2017 VTAIL.n70 VTAIL.n69 0.155672
R2018 VTAIL.n70 VTAIL.n5 0.155672
R2019 VTAIL.n79 VTAIL.n5 0.155672
R2020 VTAIL.n80 VTAIL.n79 0.155672
R2021 VTAIL.n80 VTAIL.n1 0.155672
R2022 VTAIL.n87 VTAIL.n1 0.155672
R2023 VTAIL.n267 VTAIL.n181 0.155672
R2024 VTAIL.n260 VTAIL.n181 0.155672
R2025 VTAIL.n260 VTAIL.n259 0.155672
R2026 VTAIL.n259 VTAIL.n185 0.155672
R2027 VTAIL.n251 VTAIL.n185 0.155672
R2028 VTAIL.n251 VTAIL.n250 0.155672
R2029 VTAIL.n250 VTAIL.n190 0.155672
R2030 VTAIL.n243 VTAIL.n190 0.155672
R2031 VTAIL.n243 VTAIL.n242 0.155672
R2032 VTAIL.n242 VTAIL.n194 0.155672
R2033 VTAIL.n235 VTAIL.n194 0.155672
R2034 VTAIL.n235 VTAIL.n234 0.155672
R2035 VTAIL.n234 VTAIL.n198 0.155672
R2036 VTAIL.n227 VTAIL.n198 0.155672
R2037 VTAIL.n227 VTAIL.n226 0.155672
R2038 VTAIL.n226 VTAIL.n202 0.155672
R2039 VTAIL.n219 VTAIL.n202 0.155672
R2040 VTAIL.n219 VTAIL.n218 0.155672
R2041 VTAIL.n218 VTAIL.n206 0.155672
R2042 VTAIL.n211 VTAIL.n206 0.155672
R2043 VTAIL.n177 VTAIL.n91 0.155672
R2044 VTAIL.n170 VTAIL.n91 0.155672
R2045 VTAIL.n170 VTAIL.n169 0.155672
R2046 VTAIL.n169 VTAIL.n95 0.155672
R2047 VTAIL.n161 VTAIL.n95 0.155672
R2048 VTAIL.n161 VTAIL.n160 0.155672
R2049 VTAIL.n160 VTAIL.n100 0.155672
R2050 VTAIL.n153 VTAIL.n100 0.155672
R2051 VTAIL.n153 VTAIL.n152 0.155672
R2052 VTAIL.n152 VTAIL.n104 0.155672
R2053 VTAIL.n145 VTAIL.n104 0.155672
R2054 VTAIL.n145 VTAIL.n144 0.155672
R2055 VTAIL.n144 VTAIL.n108 0.155672
R2056 VTAIL.n137 VTAIL.n108 0.155672
R2057 VTAIL.n137 VTAIL.n136 0.155672
R2058 VTAIL.n136 VTAIL.n112 0.155672
R2059 VTAIL.n129 VTAIL.n112 0.155672
R2060 VTAIL.n129 VTAIL.n128 0.155672
R2061 VTAIL.n128 VTAIL.n116 0.155672
R2062 VTAIL.n121 VTAIL.n116 0.155672
R2063 VDD1.n84 VDD1.n0 289.615
R2064 VDD1.n173 VDD1.n89 289.615
R2065 VDD1.n85 VDD1.n84 185
R2066 VDD1.n83 VDD1.n82 185
R2067 VDD1.n4 VDD1.n3 185
R2068 VDD1.n77 VDD1.n76 185
R2069 VDD1.n75 VDD1.n6 185
R2070 VDD1.n74 VDD1.n73 185
R2071 VDD1.n9 VDD1.n7 185
R2072 VDD1.n68 VDD1.n67 185
R2073 VDD1.n66 VDD1.n65 185
R2074 VDD1.n13 VDD1.n12 185
R2075 VDD1.n60 VDD1.n59 185
R2076 VDD1.n58 VDD1.n57 185
R2077 VDD1.n17 VDD1.n16 185
R2078 VDD1.n52 VDD1.n51 185
R2079 VDD1.n50 VDD1.n49 185
R2080 VDD1.n21 VDD1.n20 185
R2081 VDD1.n44 VDD1.n43 185
R2082 VDD1.n42 VDD1.n41 185
R2083 VDD1.n25 VDD1.n24 185
R2084 VDD1.n36 VDD1.n35 185
R2085 VDD1.n34 VDD1.n33 185
R2086 VDD1.n29 VDD1.n28 185
R2087 VDD1.n117 VDD1.n116 185
R2088 VDD1.n122 VDD1.n121 185
R2089 VDD1.n124 VDD1.n123 185
R2090 VDD1.n113 VDD1.n112 185
R2091 VDD1.n130 VDD1.n129 185
R2092 VDD1.n132 VDD1.n131 185
R2093 VDD1.n109 VDD1.n108 185
R2094 VDD1.n138 VDD1.n137 185
R2095 VDD1.n140 VDD1.n139 185
R2096 VDD1.n105 VDD1.n104 185
R2097 VDD1.n146 VDD1.n145 185
R2098 VDD1.n148 VDD1.n147 185
R2099 VDD1.n101 VDD1.n100 185
R2100 VDD1.n154 VDD1.n153 185
R2101 VDD1.n156 VDD1.n155 185
R2102 VDD1.n97 VDD1.n96 185
R2103 VDD1.n163 VDD1.n162 185
R2104 VDD1.n164 VDD1.n95 185
R2105 VDD1.n166 VDD1.n165 185
R2106 VDD1.n93 VDD1.n92 185
R2107 VDD1.n172 VDD1.n171 185
R2108 VDD1.n174 VDD1.n173 185
R2109 VDD1.n30 VDD1.t1 147.659
R2110 VDD1.n118 VDD1.t0 147.659
R2111 VDD1.n84 VDD1.n83 104.615
R2112 VDD1.n83 VDD1.n3 104.615
R2113 VDD1.n76 VDD1.n3 104.615
R2114 VDD1.n76 VDD1.n75 104.615
R2115 VDD1.n75 VDD1.n74 104.615
R2116 VDD1.n74 VDD1.n7 104.615
R2117 VDD1.n67 VDD1.n7 104.615
R2118 VDD1.n67 VDD1.n66 104.615
R2119 VDD1.n66 VDD1.n12 104.615
R2120 VDD1.n59 VDD1.n12 104.615
R2121 VDD1.n59 VDD1.n58 104.615
R2122 VDD1.n58 VDD1.n16 104.615
R2123 VDD1.n51 VDD1.n16 104.615
R2124 VDD1.n51 VDD1.n50 104.615
R2125 VDD1.n50 VDD1.n20 104.615
R2126 VDD1.n43 VDD1.n20 104.615
R2127 VDD1.n43 VDD1.n42 104.615
R2128 VDD1.n42 VDD1.n24 104.615
R2129 VDD1.n35 VDD1.n24 104.615
R2130 VDD1.n35 VDD1.n34 104.615
R2131 VDD1.n34 VDD1.n28 104.615
R2132 VDD1.n122 VDD1.n116 104.615
R2133 VDD1.n123 VDD1.n122 104.615
R2134 VDD1.n123 VDD1.n112 104.615
R2135 VDD1.n130 VDD1.n112 104.615
R2136 VDD1.n131 VDD1.n130 104.615
R2137 VDD1.n131 VDD1.n108 104.615
R2138 VDD1.n138 VDD1.n108 104.615
R2139 VDD1.n139 VDD1.n138 104.615
R2140 VDD1.n139 VDD1.n104 104.615
R2141 VDD1.n146 VDD1.n104 104.615
R2142 VDD1.n147 VDD1.n146 104.615
R2143 VDD1.n147 VDD1.n100 104.615
R2144 VDD1.n154 VDD1.n100 104.615
R2145 VDD1.n155 VDD1.n154 104.615
R2146 VDD1.n155 VDD1.n96 104.615
R2147 VDD1.n163 VDD1.n96 104.615
R2148 VDD1.n164 VDD1.n163 104.615
R2149 VDD1.n165 VDD1.n164 104.615
R2150 VDD1.n165 VDD1.n92 104.615
R2151 VDD1.n172 VDD1.n92 104.615
R2152 VDD1.n173 VDD1.n172 104.615
R2153 VDD1 VDD1.n177 95.197
R2154 VDD1.t1 VDD1.n28 52.3082
R2155 VDD1.t0 VDD1.n116 52.3082
R2156 VDD1 VDD1.n88 50.7002
R2157 VDD1.n30 VDD1.n29 15.6677
R2158 VDD1.n118 VDD1.n117 15.6677
R2159 VDD1.n77 VDD1.n6 13.1884
R2160 VDD1.n166 VDD1.n95 13.1884
R2161 VDD1.n78 VDD1.n4 12.8005
R2162 VDD1.n73 VDD1.n8 12.8005
R2163 VDD1.n33 VDD1.n32 12.8005
R2164 VDD1.n121 VDD1.n120 12.8005
R2165 VDD1.n162 VDD1.n161 12.8005
R2166 VDD1.n167 VDD1.n93 12.8005
R2167 VDD1.n82 VDD1.n81 12.0247
R2168 VDD1.n72 VDD1.n9 12.0247
R2169 VDD1.n36 VDD1.n27 12.0247
R2170 VDD1.n124 VDD1.n115 12.0247
R2171 VDD1.n160 VDD1.n97 12.0247
R2172 VDD1.n171 VDD1.n170 12.0247
R2173 VDD1.n85 VDD1.n2 11.249
R2174 VDD1.n69 VDD1.n68 11.249
R2175 VDD1.n37 VDD1.n25 11.249
R2176 VDD1.n125 VDD1.n113 11.249
R2177 VDD1.n157 VDD1.n156 11.249
R2178 VDD1.n174 VDD1.n91 11.249
R2179 VDD1.n86 VDD1.n0 10.4732
R2180 VDD1.n65 VDD1.n11 10.4732
R2181 VDD1.n41 VDD1.n40 10.4732
R2182 VDD1.n129 VDD1.n128 10.4732
R2183 VDD1.n153 VDD1.n99 10.4732
R2184 VDD1.n175 VDD1.n89 10.4732
R2185 VDD1.n64 VDD1.n13 9.69747
R2186 VDD1.n44 VDD1.n23 9.69747
R2187 VDD1.n132 VDD1.n111 9.69747
R2188 VDD1.n152 VDD1.n101 9.69747
R2189 VDD1.n88 VDD1.n87 9.45567
R2190 VDD1.n177 VDD1.n176 9.45567
R2191 VDD1.n56 VDD1.n55 9.3005
R2192 VDD1.n15 VDD1.n14 9.3005
R2193 VDD1.n62 VDD1.n61 9.3005
R2194 VDD1.n64 VDD1.n63 9.3005
R2195 VDD1.n11 VDD1.n10 9.3005
R2196 VDD1.n70 VDD1.n69 9.3005
R2197 VDD1.n72 VDD1.n71 9.3005
R2198 VDD1.n8 VDD1.n5 9.3005
R2199 VDD1.n87 VDD1.n86 9.3005
R2200 VDD1.n2 VDD1.n1 9.3005
R2201 VDD1.n81 VDD1.n80 9.3005
R2202 VDD1.n79 VDD1.n78 9.3005
R2203 VDD1.n54 VDD1.n53 9.3005
R2204 VDD1.n19 VDD1.n18 9.3005
R2205 VDD1.n48 VDD1.n47 9.3005
R2206 VDD1.n46 VDD1.n45 9.3005
R2207 VDD1.n23 VDD1.n22 9.3005
R2208 VDD1.n40 VDD1.n39 9.3005
R2209 VDD1.n38 VDD1.n37 9.3005
R2210 VDD1.n27 VDD1.n26 9.3005
R2211 VDD1.n32 VDD1.n31 9.3005
R2212 VDD1.n176 VDD1.n175 9.3005
R2213 VDD1.n91 VDD1.n90 9.3005
R2214 VDD1.n170 VDD1.n169 9.3005
R2215 VDD1.n168 VDD1.n167 9.3005
R2216 VDD1.n107 VDD1.n106 9.3005
R2217 VDD1.n136 VDD1.n135 9.3005
R2218 VDD1.n134 VDD1.n133 9.3005
R2219 VDD1.n111 VDD1.n110 9.3005
R2220 VDD1.n128 VDD1.n127 9.3005
R2221 VDD1.n126 VDD1.n125 9.3005
R2222 VDD1.n115 VDD1.n114 9.3005
R2223 VDD1.n120 VDD1.n119 9.3005
R2224 VDD1.n142 VDD1.n141 9.3005
R2225 VDD1.n144 VDD1.n143 9.3005
R2226 VDD1.n103 VDD1.n102 9.3005
R2227 VDD1.n150 VDD1.n149 9.3005
R2228 VDD1.n152 VDD1.n151 9.3005
R2229 VDD1.n99 VDD1.n98 9.3005
R2230 VDD1.n158 VDD1.n157 9.3005
R2231 VDD1.n160 VDD1.n159 9.3005
R2232 VDD1.n161 VDD1.n94 9.3005
R2233 VDD1.n61 VDD1.n60 8.92171
R2234 VDD1.n45 VDD1.n21 8.92171
R2235 VDD1.n133 VDD1.n109 8.92171
R2236 VDD1.n149 VDD1.n148 8.92171
R2237 VDD1.n57 VDD1.n15 8.14595
R2238 VDD1.n49 VDD1.n48 8.14595
R2239 VDD1.n137 VDD1.n136 8.14595
R2240 VDD1.n145 VDD1.n103 8.14595
R2241 VDD1.n56 VDD1.n17 7.3702
R2242 VDD1.n52 VDD1.n19 7.3702
R2243 VDD1.n140 VDD1.n107 7.3702
R2244 VDD1.n144 VDD1.n105 7.3702
R2245 VDD1.n53 VDD1.n17 6.59444
R2246 VDD1.n53 VDD1.n52 6.59444
R2247 VDD1.n141 VDD1.n140 6.59444
R2248 VDD1.n141 VDD1.n105 6.59444
R2249 VDD1.n57 VDD1.n56 5.81868
R2250 VDD1.n49 VDD1.n19 5.81868
R2251 VDD1.n137 VDD1.n107 5.81868
R2252 VDD1.n145 VDD1.n144 5.81868
R2253 VDD1.n60 VDD1.n15 5.04292
R2254 VDD1.n48 VDD1.n21 5.04292
R2255 VDD1.n136 VDD1.n109 5.04292
R2256 VDD1.n148 VDD1.n103 5.04292
R2257 VDD1.n31 VDD1.n30 4.38563
R2258 VDD1.n119 VDD1.n118 4.38563
R2259 VDD1.n61 VDD1.n13 4.26717
R2260 VDD1.n45 VDD1.n44 4.26717
R2261 VDD1.n133 VDD1.n132 4.26717
R2262 VDD1.n149 VDD1.n101 4.26717
R2263 VDD1.n88 VDD1.n0 3.49141
R2264 VDD1.n65 VDD1.n64 3.49141
R2265 VDD1.n41 VDD1.n23 3.49141
R2266 VDD1.n129 VDD1.n111 3.49141
R2267 VDD1.n153 VDD1.n152 3.49141
R2268 VDD1.n177 VDD1.n89 3.49141
R2269 VDD1.n86 VDD1.n85 2.71565
R2270 VDD1.n68 VDD1.n11 2.71565
R2271 VDD1.n40 VDD1.n25 2.71565
R2272 VDD1.n128 VDD1.n113 2.71565
R2273 VDD1.n156 VDD1.n99 2.71565
R2274 VDD1.n175 VDD1.n174 2.71565
R2275 VDD1.n82 VDD1.n2 1.93989
R2276 VDD1.n69 VDD1.n9 1.93989
R2277 VDD1.n37 VDD1.n36 1.93989
R2278 VDD1.n125 VDD1.n124 1.93989
R2279 VDD1.n157 VDD1.n97 1.93989
R2280 VDD1.n171 VDD1.n91 1.93989
R2281 VDD1.n81 VDD1.n4 1.16414
R2282 VDD1.n73 VDD1.n72 1.16414
R2283 VDD1.n33 VDD1.n27 1.16414
R2284 VDD1.n121 VDD1.n115 1.16414
R2285 VDD1.n162 VDD1.n160 1.16414
R2286 VDD1.n170 VDD1.n93 1.16414
R2287 VDD1.n78 VDD1.n77 0.388379
R2288 VDD1.n8 VDD1.n6 0.388379
R2289 VDD1.n32 VDD1.n29 0.388379
R2290 VDD1.n120 VDD1.n117 0.388379
R2291 VDD1.n161 VDD1.n95 0.388379
R2292 VDD1.n167 VDD1.n166 0.388379
R2293 VDD1.n87 VDD1.n1 0.155672
R2294 VDD1.n80 VDD1.n1 0.155672
R2295 VDD1.n80 VDD1.n79 0.155672
R2296 VDD1.n79 VDD1.n5 0.155672
R2297 VDD1.n71 VDD1.n5 0.155672
R2298 VDD1.n71 VDD1.n70 0.155672
R2299 VDD1.n70 VDD1.n10 0.155672
R2300 VDD1.n63 VDD1.n10 0.155672
R2301 VDD1.n63 VDD1.n62 0.155672
R2302 VDD1.n62 VDD1.n14 0.155672
R2303 VDD1.n55 VDD1.n14 0.155672
R2304 VDD1.n55 VDD1.n54 0.155672
R2305 VDD1.n54 VDD1.n18 0.155672
R2306 VDD1.n47 VDD1.n18 0.155672
R2307 VDD1.n47 VDD1.n46 0.155672
R2308 VDD1.n46 VDD1.n22 0.155672
R2309 VDD1.n39 VDD1.n22 0.155672
R2310 VDD1.n39 VDD1.n38 0.155672
R2311 VDD1.n38 VDD1.n26 0.155672
R2312 VDD1.n31 VDD1.n26 0.155672
R2313 VDD1.n119 VDD1.n114 0.155672
R2314 VDD1.n126 VDD1.n114 0.155672
R2315 VDD1.n127 VDD1.n126 0.155672
R2316 VDD1.n127 VDD1.n110 0.155672
R2317 VDD1.n134 VDD1.n110 0.155672
R2318 VDD1.n135 VDD1.n134 0.155672
R2319 VDD1.n135 VDD1.n106 0.155672
R2320 VDD1.n142 VDD1.n106 0.155672
R2321 VDD1.n143 VDD1.n142 0.155672
R2322 VDD1.n143 VDD1.n102 0.155672
R2323 VDD1.n150 VDD1.n102 0.155672
R2324 VDD1.n151 VDD1.n150 0.155672
R2325 VDD1.n151 VDD1.n98 0.155672
R2326 VDD1.n158 VDD1.n98 0.155672
R2327 VDD1.n159 VDD1.n158 0.155672
R2328 VDD1.n159 VDD1.n94 0.155672
R2329 VDD1.n168 VDD1.n94 0.155672
R2330 VDD1.n169 VDD1.n168 0.155672
R2331 VDD1.n169 VDD1.n90 0.155672
R2332 VDD1.n176 VDD1.n90 0.155672
R2333 VN VN.t0 202.32
R2334 VN VN.t1 152.978
R2335 VDD2.n173 VDD2.n89 289.615
R2336 VDD2.n84 VDD2.n0 289.615
R2337 VDD2.n174 VDD2.n173 185
R2338 VDD2.n172 VDD2.n171 185
R2339 VDD2.n93 VDD2.n92 185
R2340 VDD2.n166 VDD2.n165 185
R2341 VDD2.n164 VDD2.n95 185
R2342 VDD2.n163 VDD2.n162 185
R2343 VDD2.n98 VDD2.n96 185
R2344 VDD2.n157 VDD2.n156 185
R2345 VDD2.n155 VDD2.n154 185
R2346 VDD2.n102 VDD2.n101 185
R2347 VDD2.n149 VDD2.n148 185
R2348 VDD2.n147 VDD2.n146 185
R2349 VDD2.n106 VDD2.n105 185
R2350 VDD2.n141 VDD2.n140 185
R2351 VDD2.n139 VDD2.n138 185
R2352 VDD2.n110 VDD2.n109 185
R2353 VDD2.n133 VDD2.n132 185
R2354 VDD2.n131 VDD2.n130 185
R2355 VDD2.n114 VDD2.n113 185
R2356 VDD2.n125 VDD2.n124 185
R2357 VDD2.n123 VDD2.n122 185
R2358 VDD2.n118 VDD2.n117 185
R2359 VDD2.n28 VDD2.n27 185
R2360 VDD2.n33 VDD2.n32 185
R2361 VDD2.n35 VDD2.n34 185
R2362 VDD2.n24 VDD2.n23 185
R2363 VDD2.n41 VDD2.n40 185
R2364 VDD2.n43 VDD2.n42 185
R2365 VDD2.n20 VDD2.n19 185
R2366 VDD2.n49 VDD2.n48 185
R2367 VDD2.n51 VDD2.n50 185
R2368 VDD2.n16 VDD2.n15 185
R2369 VDD2.n57 VDD2.n56 185
R2370 VDD2.n59 VDD2.n58 185
R2371 VDD2.n12 VDD2.n11 185
R2372 VDD2.n65 VDD2.n64 185
R2373 VDD2.n67 VDD2.n66 185
R2374 VDD2.n8 VDD2.n7 185
R2375 VDD2.n74 VDD2.n73 185
R2376 VDD2.n75 VDD2.n6 185
R2377 VDD2.n77 VDD2.n76 185
R2378 VDD2.n4 VDD2.n3 185
R2379 VDD2.n83 VDD2.n82 185
R2380 VDD2.n85 VDD2.n84 185
R2381 VDD2.n119 VDD2.t1 147.659
R2382 VDD2.n29 VDD2.t0 147.659
R2383 VDD2.n173 VDD2.n172 104.615
R2384 VDD2.n172 VDD2.n92 104.615
R2385 VDD2.n165 VDD2.n92 104.615
R2386 VDD2.n165 VDD2.n164 104.615
R2387 VDD2.n164 VDD2.n163 104.615
R2388 VDD2.n163 VDD2.n96 104.615
R2389 VDD2.n156 VDD2.n96 104.615
R2390 VDD2.n156 VDD2.n155 104.615
R2391 VDD2.n155 VDD2.n101 104.615
R2392 VDD2.n148 VDD2.n101 104.615
R2393 VDD2.n148 VDD2.n147 104.615
R2394 VDD2.n147 VDD2.n105 104.615
R2395 VDD2.n140 VDD2.n105 104.615
R2396 VDD2.n140 VDD2.n139 104.615
R2397 VDD2.n139 VDD2.n109 104.615
R2398 VDD2.n132 VDD2.n109 104.615
R2399 VDD2.n132 VDD2.n131 104.615
R2400 VDD2.n131 VDD2.n113 104.615
R2401 VDD2.n124 VDD2.n113 104.615
R2402 VDD2.n124 VDD2.n123 104.615
R2403 VDD2.n123 VDD2.n117 104.615
R2404 VDD2.n33 VDD2.n27 104.615
R2405 VDD2.n34 VDD2.n33 104.615
R2406 VDD2.n34 VDD2.n23 104.615
R2407 VDD2.n41 VDD2.n23 104.615
R2408 VDD2.n42 VDD2.n41 104.615
R2409 VDD2.n42 VDD2.n19 104.615
R2410 VDD2.n49 VDD2.n19 104.615
R2411 VDD2.n50 VDD2.n49 104.615
R2412 VDD2.n50 VDD2.n15 104.615
R2413 VDD2.n57 VDD2.n15 104.615
R2414 VDD2.n58 VDD2.n57 104.615
R2415 VDD2.n58 VDD2.n11 104.615
R2416 VDD2.n65 VDD2.n11 104.615
R2417 VDD2.n66 VDD2.n65 104.615
R2418 VDD2.n66 VDD2.n7 104.615
R2419 VDD2.n74 VDD2.n7 104.615
R2420 VDD2.n75 VDD2.n74 104.615
R2421 VDD2.n76 VDD2.n75 104.615
R2422 VDD2.n76 VDD2.n3 104.615
R2423 VDD2.n83 VDD2.n3 104.615
R2424 VDD2.n84 VDD2.n83 104.615
R2425 VDD2.n178 VDD2.n88 93.864
R2426 VDD2.t1 VDD2.n117 52.3082
R2427 VDD2.t0 VDD2.n27 52.3082
R2428 VDD2.n178 VDD2.n177 49.8338
R2429 VDD2.n119 VDD2.n118 15.6677
R2430 VDD2.n29 VDD2.n28 15.6677
R2431 VDD2.n166 VDD2.n95 13.1884
R2432 VDD2.n77 VDD2.n6 13.1884
R2433 VDD2.n167 VDD2.n93 12.8005
R2434 VDD2.n162 VDD2.n97 12.8005
R2435 VDD2.n122 VDD2.n121 12.8005
R2436 VDD2.n32 VDD2.n31 12.8005
R2437 VDD2.n73 VDD2.n72 12.8005
R2438 VDD2.n78 VDD2.n4 12.8005
R2439 VDD2.n171 VDD2.n170 12.0247
R2440 VDD2.n161 VDD2.n98 12.0247
R2441 VDD2.n125 VDD2.n116 12.0247
R2442 VDD2.n35 VDD2.n26 12.0247
R2443 VDD2.n71 VDD2.n8 12.0247
R2444 VDD2.n82 VDD2.n81 12.0247
R2445 VDD2.n174 VDD2.n91 11.249
R2446 VDD2.n158 VDD2.n157 11.249
R2447 VDD2.n126 VDD2.n114 11.249
R2448 VDD2.n36 VDD2.n24 11.249
R2449 VDD2.n68 VDD2.n67 11.249
R2450 VDD2.n85 VDD2.n2 11.249
R2451 VDD2.n175 VDD2.n89 10.4732
R2452 VDD2.n154 VDD2.n100 10.4732
R2453 VDD2.n130 VDD2.n129 10.4732
R2454 VDD2.n40 VDD2.n39 10.4732
R2455 VDD2.n64 VDD2.n10 10.4732
R2456 VDD2.n86 VDD2.n0 10.4732
R2457 VDD2.n153 VDD2.n102 9.69747
R2458 VDD2.n133 VDD2.n112 9.69747
R2459 VDD2.n43 VDD2.n22 9.69747
R2460 VDD2.n63 VDD2.n12 9.69747
R2461 VDD2.n177 VDD2.n176 9.45567
R2462 VDD2.n88 VDD2.n87 9.45567
R2463 VDD2.n145 VDD2.n144 9.3005
R2464 VDD2.n104 VDD2.n103 9.3005
R2465 VDD2.n151 VDD2.n150 9.3005
R2466 VDD2.n153 VDD2.n152 9.3005
R2467 VDD2.n100 VDD2.n99 9.3005
R2468 VDD2.n159 VDD2.n158 9.3005
R2469 VDD2.n161 VDD2.n160 9.3005
R2470 VDD2.n97 VDD2.n94 9.3005
R2471 VDD2.n176 VDD2.n175 9.3005
R2472 VDD2.n91 VDD2.n90 9.3005
R2473 VDD2.n170 VDD2.n169 9.3005
R2474 VDD2.n168 VDD2.n167 9.3005
R2475 VDD2.n143 VDD2.n142 9.3005
R2476 VDD2.n108 VDD2.n107 9.3005
R2477 VDD2.n137 VDD2.n136 9.3005
R2478 VDD2.n135 VDD2.n134 9.3005
R2479 VDD2.n112 VDD2.n111 9.3005
R2480 VDD2.n129 VDD2.n128 9.3005
R2481 VDD2.n127 VDD2.n126 9.3005
R2482 VDD2.n116 VDD2.n115 9.3005
R2483 VDD2.n121 VDD2.n120 9.3005
R2484 VDD2.n87 VDD2.n86 9.3005
R2485 VDD2.n2 VDD2.n1 9.3005
R2486 VDD2.n81 VDD2.n80 9.3005
R2487 VDD2.n79 VDD2.n78 9.3005
R2488 VDD2.n18 VDD2.n17 9.3005
R2489 VDD2.n47 VDD2.n46 9.3005
R2490 VDD2.n45 VDD2.n44 9.3005
R2491 VDD2.n22 VDD2.n21 9.3005
R2492 VDD2.n39 VDD2.n38 9.3005
R2493 VDD2.n37 VDD2.n36 9.3005
R2494 VDD2.n26 VDD2.n25 9.3005
R2495 VDD2.n31 VDD2.n30 9.3005
R2496 VDD2.n53 VDD2.n52 9.3005
R2497 VDD2.n55 VDD2.n54 9.3005
R2498 VDD2.n14 VDD2.n13 9.3005
R2499 VDD2.n61 VDD2.n60 9.3005
R2500 VDD2.n63 VDD2.n62 9.3005
R2501 VDD2.n10 VDD2.n9 9.3005
R2502 VDD2.n69 VDD2.n68 9.3005
R2503 VDD2.n71 VDD2.n70 9.3005
R2504 VDD2.n72 VDD2.n5 9.3005
R2505 VDD2.n150 VDD2.n149 8.92171
R2506 VDD2.n134 VDD2.n110 8.92171
R2507 VDD2.n44 VDD2.n20 8.92171
R2508 VDD2.n60 VDD2.n59 8.92171
R2509 VDD2.n146 VDD2.n104 8.14595
R2510 VDD2.n138 VDD2.n137 8.14595
R2511 VDD2.n48 VDD2.n47 8.14595
R2512 VDD2.n56 VDD2.n14 8.14595
R2513 VDD2.n145 VDD2.n106 7.3702
R2514 VDD2.n141 VDD2.n108 7.3702
R2515 VDD2.n51 VDD2.n18 7.3702
R2516 VDD2.n55 VDD2.n16 7.3702
R2517 VDD2.n142 VDD2.n106 6.59444
R2518 VDD2.n142 VDD2.n141 6.59444
R2519 VDD2.n52 VDD2.n51 6.59444
R2520 VDD2.n52 VDD2.n16 6.59444
R2521 VDD2.n146 VDD2.n145 5.81868
R2522 VDD2.n138 VDD2.n108 5.81868
R2523 VDD2.n48 VDD2.n18 5.81868
R2524 VDD2.n56 VDD2.n55 5.81868
R2525 VDD2.n149 VDD2.n104 5.04292
R2526 VDD2.n137 VDD2.n110 5.04292
R2527 VDD2.n47 VDD2.n20 5.04292
R2528 VDD2.n59 VDD2.n14 5.04292
R2529 VDD2.n120 VDD2.n119 4.38563
R2530 VDD2.n30 VDD2.n29 4.38563
R2531 VDD2.n150 VDD2.n102 4.26717
R2532 VDD2.n134 VDD2.n133 4.26717
R2533 VDD2.n44 VDD2.n43 4.26717
R2534 VDD2.n60 VDD2.n12 4.26717
R2535 VDD2.n177 VDD2.n89 3.49141
R2536 VDD2.n154 VDD2.n153 3.49141
R2537 VDD2.n130 VDD2.n112 3.49141
R2538 VDD2.n40 VDD2.n22 3.49141
R2539 VDD2.n64 VDD2.n63 3.49141
R2540 VDD2.n88 VDD2.n0 3.49141
R2541 VDD2.n175 VDD2.n174 2.71565
R2542 VDD2.n157 VDD2.n100 2.71565
R2543 VDD2.n129 VDD2.n114 2.71565
R2544 VDD2.n39 VDD2.n24 2.71565
R2545 VDD2.n67 VDD2.n10 2.71565
R2546 VDD2.n86 VDD2.n85 2.71565
R2547 VDD2.n171 VDD2.n91 1.93989
R2548 VDD2.n158 VDD2.n98 1.93989
R2549 VDD2.n126 VDD2.n125 1.93989
R2550 VDD2.n36 VDD2.n35 1.93989
R2551 VDD2.n68 VDD2.n8 1.93989
R2552 VDD2.n82 VDD2.n2 1.93989
R2553 VDD2.n170 VDD2.n93 1.16414
R2554 VDD2.n162 VDD2.n161 1.16414
R2555 VDD2.n122 VDD2.n116 1.16414
R2556 VDD2.n32 VDD2.n26 1.16414
R2557 VDD2.n73 VDD2.n71 1.16414
R2558 VDD2.n81 VDD2.n4 1.16414
R2559 VDD2 VDD2.n178 0.866879
R2560 VDD2.n167 VDD2.n166 0.388379
R2561 VDD2.n97 VDD2.n95 0.388379
R2562 VDD2.n121 VDD2.n118 0.388379
R2563 VDD2.n31 VDD2.n28 0.388379
R2564 VDD2.n72 VDD2.n6 0.388379
R2565 VDD2.n78 VDD2.n77 0.388379
R2566 VDD2.n176 VDD2.n90 0.155672
R2567 VDD2.n169 VDD2.n90 0.155672
R2568 VDD2.n169 VDD2.n168 0.155672
R2569 VDD2.n168 VDD2.n94 0.155672
R2570 VDD2.n160 VDD2.n94 0.155672
R2571 VDD2.n160 VDD2.n159 0.155672
R2572 VDD2.n159 VDD2.n99 0.155672
R2573 VDD2.n152 VDD2.n99 0.155672
R2574 VDD2.n152 VDD2.n151 0.155672
R2575 VDD2.n151 VDD2.n103 0.155672
R2576 VDD2.n144 VDD2.n103 0.155672
R2577 VDD2.n144 VDD2.n143 0.155672
R2578 VDD2.n143 VDD2.n107 0.155672
R2579 VDD2.n136 VDD2.n107 0.155672
R2580 VDD2.n136 VDD2.n135 0.155672
R2581 VDD2.n135 VDD2.n111 0.155672
R2582 VDD2.n128 VDD2.n111 0.155672
R2583 VDD2.n128 VDD2.n127 0.155672
R2584 VDD2.n127 VDD2.n115 0.155672
R2585 VDD2.n120 VDD2.n115 0.155672
R2586 VDD2.n30 VDD2.n25 0.155672
R2587 VDD2.n37 VDD2.n25 0.155672
R2588 VDD2.n38 VDD2.n37 0.155672
R2589 VDD2.n38 VDD2.n21 0.155672
R2590 VDD2.n45 VDD2.n21 0.155672
R2591 VDD2.n46 VDD2.n45 0.155672
R2592 VDD2.n46 VDD2.n17 0.155672
R2593 VDD2.n53 VDD2.n17 0.155672
R2594 VDD2.n54 VDD2.n53 0.155672
R2595 VDD2.n54 VDD2.n13 0.155672
R2596 VDD2.n61 VDD2.n13 0.155672
R2597 VDD2.n62 VDD2.n61 0.155672
R2598 VDD2.n62 VDD2.n9 0.155672
R2599 VDD2.n69 VDD2.n9 0.155672
R2600 VDD2.n70 VDD2.n69 0.155672
R2601 VDD2.n70 VDD2.n5 0.155672
R2602 VDD2.n79 VDD2.n5 0.155672
R2603 VDD2.n80 VDD2.n79 0.155672
R2604 VDD2.n80 VDD2.n1 0.155672
R2605 VDD2.n87 VDD2.n1 0.155672
C0 VP VN 6.60534f
C1 VP VTAIL 3.33148f
C2 VN VDD1 0.148499f
C3 VTAIL VDD1 6.26553f
C4 VN VDD2 3.7917f
C5 VTAIL VDD2 6.32164f
C6 VP VDD1 4.00822f
C7 VN VTAIL 3.3172f
C8 VP VDD2 0.367781f
C9 VDD1 VDD2 0.775072f
C10 VDD2 B 5.454754f
C11 VDD1 B 8.66895f
C12 VTAIL B 9.449872f
C13 VN B 12.454269f
C14 VP B 7.692243f
C15 VDD2.n0 B 0.027279f
C16 VDD2.n1 B 0.020082f
C17 VDD2.n2 B 0.010791f
C18 VDD2.n3 B 0.025507f
C19 VDD2.n4 B 0.011426f
C20 VDD2.n5 B 0.020082f
C21 VDD2.n6 B 0.011109f
C22 VDD2.n7 B 0.025507f
C23 VDD2.n8 B 0.011426f
C24 VDD2.n9 B 0.020082f
C25 VDD2.n10 B 0.010791f
C26 VDD2.n11 B 0.025507f
C27 VDD2.n12 B 0.011426f
C28 VDD2.n13 B 0.020082f
C29 VDD2.n14 B 0.010791f
C30 VDD2.n15 B 0.025507f
C31 VDD2.n16 B 0.011426f
C32 VDD2.n17 B 0.020082f
C33 VDD2.n18 B 0.010791f
C34 VDD2.n19 B 0.025507f
C35 VDD2.n20 B 0.011426f
C36 VDD2.n21 B 0.020082f
C37 VDD2.n22 B 0.010791f
C38 VDD2.n23 B 0.025507f
C39 VDD2.n24 B 0.011426f
C40 VDD2.n25 B 0.020082f
C41 VDD2.n26 B 0.010791f
C42 VDD2.n27 B 0.01913f
C43 VDD2.n28 B 0.015067f
C44 VDD2.t0 B 0.042135f
C45 VDD2.n29 B 0.136669f
C46 VDD2.n30 B 1.41057f
C47 VDD2.n31 B 0.010791f
C48 VDD2.n32 B 0.011426f
C49 VDD2.n33 B 0.025507f
C50 VDD2.n34 B 0.025507f
C51 VDD2.n35 B 0.011426f
C52 VDD2.n36 B 0.010791f
C53 VDD2.n37 B 0.020082f
C54 VDD2.n38 B 0.020082f
C55 VDD2.n39 B 0.010791f
C56 VDD2.n40 B 0.011426f
C57 VDD2.n41 B 0.025507f
C58 VDD2.n42 B 0.025507f
C59 VDD2.n43 B 0.011426f
C60 VDD2.n44 B 0.010791f
C61 VDD2.n45 B 0.020082f
C62 VDD2.n46 B 0.020082f
C63 VDD2.n47 B 0.010791f
C64 VDD2.n48 B 0.011426f
C65 VDD2.n49 B 0.025507f
C66 VDD2.n50 B 0.025507f
C67 VDD2.n51 B 0.011426f
C68 VDD2.n52 B 0.010791f
C69 VDD2.n53 B 0.020082f
C70 VDD2.n54 B 0.020082f
C71 VDD2.n55 B 0.010791f
C72 VDD2.n56 B 0.011426f
C73 VDD2.n57 B 0.025507f
C74 VDD2.n58 B 0.025507f
C75 VDD2.n59 B 0.011426f
C76 VDD2.n60 B 0.010791f
C77 VDD2.n61 B 0.020082f
C78 VDD2.n62 B 0.020082f
C79 VDD2.n63 B 0.010791f
C80 VDD2.n64 B 0.011426f
C81 VDD2.n65 B 0.025507f
C82 VDD2.n66 B 0.025507f
C83 VDD2.n67 B 0.011426f
C84 VDD2.n68 B 0.010791f
C85 VDD2.n69 B 0.020082f
C86 VDD2.n70 B 0.020082f
C87 VDD2.n71 B 0.010791f
C88 VDD2.n72 B 0.010791f
C89 VDD2.n73 B 0.011426f
C90 VDD2.n74 B 0.025507f
C91 VDD2.n75 B 0.025507f
C92 VDD2.n76 B 0.025507f
C93 VDD2.n77 B 0.011109f
C94 VDD2.n78 B 0.010791f
C95 VDD2.n79 B 0.020082f
C96 VDD2.n80 B 0.020082f
C97 VDD2.n81 B 0.010791f
C98 VDD2.n82 B 0.011426f
C99 VDD2.n83 B 0.025507f
C100 VDD2.n84 B 0.05354f
C101 VDD2.n85 B 0.011426f
C102 VDD2.n86 B 0.010791f
C103 VDD2.n87 B 0.04779f
C104 VDD2.n88 B 0.750603f
C105 VDD2.n89 B 0.027279f
C106 VDD2.n90 B 0.020082f
C107 VDD2.n91 B 0.010791f
C108 VDD2.n92 B 0.025507f
C109 VDD2.n93 B 0.011426f
C110 VDD2.n94 B 0.020082f
C111 VDD2.n95 B 0.011109f
C112 VDD2.n96 B 0.025507f
C113 VDD2.n97 B 0.010791f
C114 VDD2.n98 B 0.011426f
C115 VDD2.n99 B 0.020082f
C116 VDD2.n100 B 0.010791f
C117 VDD2.n101 B 0.025507f
C118 VDD2.n102 B 0.011426f
C119 VDD2.n103 B 0.020082f
C120 VDD2.n104 B 0.010791f
C121 VDD2.n105 B 0.025507f
C122 VDD2.n106 B 0.011426f
C123 VDD2.n107 B 0.020082f
C124 VDD2.n108 B 0.010791f
C125 VDD2.n109 B 0.025507f
C126 VDD2.n110 B 0.011426f
C127 VDD2.n111 B 0.020082f
C128 VDD2.n112 B 0.010791f
C129 VDD2.n113 B 0.025507f
C130 VDD2.n114 B 0.011426f
C131 VDD2.n115 B 0.020082f
C132 VDD2.n116 B 0.010791f
C133 VDD2.n117 B 0.01913f
C134 VDD2.n118 B 0.015067f
C135 VDD2.t1 B 0.042135f
C136 VDD2.n119 B 0.136669f
C137 VDD2.n120 B 1.41057f
C138 VDD2.n121 B 0.010791f
C139 VDD2.n122 B 0.011426f
C140 VDD2.n123 B 0.025507f
C141 VDD2.n124 B 0.025507f
C142 VDD2.n125 B 0.011426f
C143 VDD2.n126 B 0.010791f
C144 VDD2.n127 B 0.020082f
C145 VDD2.n128 B 0.020082f
C146 VDD2.n129 B 0.010791f
C147 VDD2.n130 B 0.011426f
C148 VDD2.n131 B 0.025507f
C149 VDD2.n132 B 0.025507f
C150 VDD2.n133 B 0.011426f
C151 VDD2.n134 B 0.010791f
C152 VDD2.n135 B 0.020082f
C153 VDD2.n136 B 0.020082f
C154 VDD2.n137 B 0.010791f
C155 VDD2.n138 B 0.011426f
C156 VDD2.n139 B 0.025507f
C157 VDD2.n140 B 0.025507f
C158 VDD2.n141 B 0.011426f
C159 VDD2.n142 B 0.010791f
C160 VDD2.n143 B 0.020082f
C161 VDD2.n144 B 0.020082f
C162 VDD2.n145 B 0.010791f
C163 VDD2.n146 B 0.011426f
C164 VDD2.n147 B 0.025507f
C165 VDD2.n148 B 0.025507f
C166 VDD2.n149 B 0.011426f
C167 VDD2.n150 B 0.010791f
C168 VDD2.n151 B 0.020082f
C169 VDD2.n152 B 0.020082f
C170 VDD2.n153 B 0.010791f
C171 VDD2.n154 B 0.011426f
C172 VDD2.n155 B 0.025507f
C173 VDD2.n156 B 0.025507f
C174 VDD2.n157 B 0.011426f
C175 VDD2.n158 B 0.010791f
C176 VDD2.n159 B 0.020082f
C177 VDD2.n160 B 0.020082f
C178 VDD2.n161 B 0.010791f
C179 VDD2.n162 B 0.011426f
C180 VDD2.n163 B 0.025507f
C181 VDD2.n164 B 0.025507f
C182 VDD2.n165 B 0.025507f
C183 VDD2.n166 B 0.011109f
C184 VDD2.n167 B 0.010791f
C185 VDD2.n168 B 0.020082f
C186 VDD2.n169 B 0.020082f
C187 VDD2.n170 B 0.010791f
C188 VDD2.n171 B 0.011426f
C189 VDD2.n172 B 0.025507f
C190 VDD2.n173 B 0.05354f
C191 VDD2.n174 B 0.011426f
C192 VDD2.n175 B 0.010791f
C193 VDD2.n176 B 0.04779f
C194 VDD2.n177 B 0.043682f
C195 VDD2.n178 B 2.92492f
C196 VN.t1 B 4.1616f
C197 VN.t0 B 4.81502f
C198 VDD1.n0 B 0.027616f
C199 VDD1.n1 B 0.02033f
C200 VDD1.n2 B 0.010925f
C201 VDD1.n3 B 0.025822f
C202 VDD1.n4 B 0.011567f
C203 VDD1.n5 B 0.02033f
C204 VDD1.n6 B 0.011246f
C205 VDD1.n7 B 0.025822f
C206 VDD1.n8 B 0.010925f
C207 VDD1.n9 B 0.011567f
C208 VDD1.n10 B 0.02033f
C209 VDD1.n11 B 0.010925f
C210 VDD1.n12 B 0.025822f
C211 VDD1.n13 B 0.011567f
C212 VDD1.n14 B 0.02033f
C213 VDD1.n15 B 0.010925f
C214 VDD1.n16 B 0.025822f
C215 VDD1.n17 B 0.011567f
C216 VDD1.n18 B 0.02033f
C217 VDD1.n19 B 0.010925f
C218 VDD1.n20 B 0.025822f
C219 VDD1.n21 B 0.011567f
C220 VDD1.n22 B 0.02033f
C221 VDD1.n23 B 0.010925f
C222 VDD1.n24 B 0.025822f
C223 VDD1.n25 B 0.011567f
C224 VDD1.n26 B 0.02033f
C225 VDD1.n27 B 0.010925f
C226 VDD1.n28 B 0.019366f
C227 VDD1.n29 B 0.015254f
C228 VDD1.t1 B 0.042656f
C229 VDD1.n30 B 0.138359f
C230 VDD1.n31 B 1.42801f
C231 VDD1.n32 B 0.010925f
C232 VDD1.n33 B 0.011567f
C233 VDD1.n34 B 0.025822f
C234 VDD1.n35 B 0.025822f
C235 VDD1.n36 B 0.011567f
C236 VDD1.n37 B 0.010925f
C237 VDD1.n38 B 0.02033f
C238 VDD1.n39 B 0.02033f
C239 VDD1.n40 B 0.010925f
C240 VDD1.n41 B 0.011567f
C241 VDD1.n42 B 0.025822f
C242 VDD1.n43 B 0.025822f
C243 VDD1.n44 B 0.011567f
C244 VDD1.n45 B 0.010925f
C245 VDD1.n46 B 0.02033f
C246 VDD1.n47 B 0.02033f
C247 VDD1.n48 B 0.010925f
C248 VDD1.n49 B 0.011567f
C249 VDD1.n50 B 0.025822f
C250 VDD1.n51 B 0.025822f
C251 VDD1.n52 B 0.011567f
C252 VDD1.n53 B 0.010925f
C253 VDD1.n54 B 0.02033f
C254 VDD1.n55 B 0.02033f
C255 VDD1.n56 B 0.010925f
C256 VDD1.n57 B 0.011567f
C257 VDD1.n58 B 0.025822f
C258 VDD1.n59 B 0.025822f
C259 VDD1.n60 B 0.011567f
C260 VDD1.n61 B 0.010925f
C261 VDD1.n62 B 0.02033f
C262 VDD1.n63 B 0.02033f
C263 VDD1.n64 B 0.010925f
C264 VDD1.n65 B 0.011567f
C265 VDD1.n66 B 0.025822f
C266 VDD1.n67 B 0.025822f
C267 VDD1.n68 B 0.011567f
C268 VDD1.n69 B 0.010925f
C269 VDD1.n70 B 0.02033f
C270 VDD1.n71 B 0.02033f
C271 VDD1.n72 B 0.010925f
C272 VDD1.n73 B 0.011567f
C273 VDD1.n74 B 0.025822f
C274 VDD1.n75 B 0.025822f
C275 VDD1.n76 B 0.025822f
C276 VDD1.n77 B 0.011246f
C277 VDD1.n78 B 0.010925f
C278 VDD1.n79 B 0.02033f
C279 VDD1.n80 B 0.02033f
C280 VDD1.n81 B 0.010925f
C281 VDD1.n82 B 0.011567f
C282 VDD1.n83 B 0.025822f
C283 VDD1.n84 B 0.054202f
C284 VDD1.n85 B 0.011567f
C285 VDD1.n86 B 0.010925f
C286 VDD1.n87 B 0.048381f
C287 VDD1.n88 B 0.045875f
C288 VDD1.n89 B 0.027616f
C289 VDD1.n90 B 0.02033f
C290 VDD1.n91 B 0.010925f
C291 VDD1.n92 B 0.025822f
C292 VDD1.n93 B 0.011567f
C293 VDD1.n94 B 0.02033f
C294 VDD1.n95 B 0.011246f
C295 VDD1.n96 B 0.025822f
C296 VDD1.n97 B 0.011567f
C297 VDD1.n98 B 0.02033f
C298 VDD1.n99 B 0.010925f
C299 VDD1.n100 B 0.025822f
C300 VDD1.n101 B 0.011567f
C301 VDD1.n102 B 0.02033f
C302 VDD1.n103 B 0.010925f
C303 VDD1.n104 B 0.025822f
C304 VDD1.n105 B 0.011567f
C305 VDD1.n106 B 0.02033f
C306 VDD1.n107 B 0.010925f
C307 VDD1.n108 B 0.025822f
C308 VDD1.n109 B 0.011567f
C309 VDD1.n110 B 0.02033f
C310 VDD1.n111 B 0.010925f
C311 VDD1.n112 B 0.025822f
C312 VDD1.n113 B 0.011567f
C313 VDD1.n114 B 0.02033f
C314 VDD1.n115 B 0.010925f
C315 VDD1.n116 B 0.019366f
C316 VDD1.n117 B 0.015254f
C317 VDD1.t0 B 0.042656f
C318 VDD1.n118 B 0.138359f
C319 VDD1.n119 B 1.42801f
C320 VDD1.n120 B 0.010925f
C321 VDD1.n121 B 0.011567f
C322 VDD1.n122 B 0.025822f
C323 VDD1.n123 B 0.025822f
C324 VDD1.n124 B 0.011567f
C325 VDD1.n125 B 0.010925f
C326 VDD1.n126 B 0.02033f
C327 VDD1.n127 B 0.02033f
C328 VDD1.n128 B 0.010925f
C329 VDD1.n129 B 0.011567f
C330 VDD1.n130 B 0.025822f
C331 VDD1.n131 B 0.025822f
C332 VDD1.n132 B 0.011567f
C333 VDD1.n133 B 0.010925f
C334 VDD1.n134 B 0.02033f
C335 VDD1.n135 B 0.02033f
C336 VDD1.n136 B 0.010925f
C337 VDD1.n137 B 0.011567f
C338 VDD1.n138 B 0.025822f
C339 VDD1.n139 B 0.025822f
C340 VDD1.n140 B 0.011567f
C341 VDD1.n141 B 0.010925f
C342 VDD1.n142 B 0.02033f
C343 VDD1.n143 B 0.02033f
C344 VDD1.n144 B 0.010925f
C345 VDD1.n145 B 0.011567f
C346 VDD1.n146 B 0.025822f
C347 VDD1.n147 B 0.025822f
C348 VDD1.n148 B 0.011567f
C349 VDD1.n149 B 0.010925f
C350 VDD1.n150 B 0.02033f
C351 VDD1.n151 B 0.02033f
C352 VDD1.n152 B 0.010925f
C353 VDD1.n153 B 0.011567f
C354 VDD1.n154 B 0.025822f
C355 VDD1.n155 B 0.025822f
C356 VDD1.n156 B 0.011567f
C357 VDD1.n157 B 0.010925f
C358 VDD1.n158 B 0.02033f
C359 VDD1.n159 B 0.02033f
C360 VDD1.n160 B 0.010925f
C361 VDD1.n161 B 0.010925f
C362 VDD1.n162 B 0.011567f
C363 VDD1.n163 B 0.025822f
C364 VDD1.n164 B 0.025822f
C365 VDD1.n165 B 0.025822f
C366 VDD1.n166 B 0.011246f
C367 VDD1.n167 B 0.010925f
C368 VDD1.n168 B 0.02033f
C369 VDD1.n169 B 0.02033f
C370 VDD1.n170 B 0.010925f
C371 VDD1.n171 B 0.011567f
C372 VDD1.n172 B 0.025822f
C373 VDD1.n173 B 0.054202f
C374 VDD1.n174 B 0.011567f
C375 VDD1.n175 B 0.010925f
C376 VDD1.n176 B 0.048381f
C377 VDD1.n177 B 0.808446f
C378 VTAIL.n0 B 0.027399f
C379 VTAIL.n1 B 0.020171f
C380 VTAIL.n2 B 0.010839f
C381 VTAIL.n3 B 0.025619f
C382 VTAIL.n4 B 0.011476f
C383 VTAIL.n5 B 0.020171f
C384 VTAIL.n6 B 0.011158f
C385 VTAIL.n7 B 0.025619f
C386 VTAIL.n8 B 0.011476f
C387 VTAIL.n9 B 0.020171f
C388 VTAIL.n10 B 0.010839f
C389 VTAIL.n11 B 0.025619f
C390 VTAIL.n12 B 0.011476f
C391 VTAIL.n13 B 0.020171f
C392 VTAIL.n14 B 0.010839f
C393 VTAIL.n15 B 0.025619f
C394 VTAIL.n16 B 0.011476f
C395 VTAIL.n17 B 0.020171f
C396 VTAIL.n18 B 0.010839f
C397 VTAIL.n19 B 0.025619f
C398 VTAIL.n20 B 0.011476f
C399 VTAIL.n21 B 0.020171f
C400 VTAIL.n22 B 0.010839f
C401 VTAIL.n23 B 0.025619f
C402 VTAIL.n24 B 0.011476f
C403 VTAIL.n25 B 0.020171f
C404 VTAIL.n26 B 0.010839f
C405 VTAIL.n27 B 0.019214f
C406 VTAIL.n28 B 0.015134f
C407 VTAIL.t3 B 0.042321f
C408 VTAIL.n29 B 0.137272f
C409 VTAIL.n30 B 1.41679f
C410 VTAIL.n31 B 0.010839f
C411 VTAIL.n32 B 0.011476f
C412 VTAIL.n33 B 0.025619f
C413 VTAIL.n34 B 0.025619f
C414 VTAIL.n35 B 0.011476f
C415 VTAIL.n36 B 0.010839f
C416 VTAIL.n37 B 0.020171f
C417 VTAIL.n38 B 0.020171f
C418 VTAIL.n39 B 0.010839f
C419 VTAIL.n40 B 0.011476f
C420 VTAIL.n41 B 0.025619f
C421 VTAIL.n42 B 0.025619f
C422 VTAIL.n43 B 0.011476f
C423 VTAIL.n44 B 0.010839f
C424 VTAIL.n45 B 0.020171f
C425 VTAIL.n46 B 0.020171f
C426 VTAIL.n47 B 0.010839f
C427 VTAIL.n48 B 0.011476f
C428 VTAIL.n49 B 0.025619f
C429 VTAIL.n50 B 0.025619f
C430 VTAIL.n51 B 0.011476f
C431 VTAIL.n52 B 0.010839f
C432 VTAIL.n53 B 0.020171f
C433 VTAIL.n54 B 0.020171f
C434 VTAIL.n55 B 0.010839f
C435 VTAIL.n56 B 0.011476f
C436 VTAIL.n57 B 0.025619f
C437 VTAIL.n58 B 0.025619f
C438 VTAIL.n59 B 0.011476f
C439 VTAIL.n60 B 0.010839f
C440 VTAIL.n61 B 0.020171f
C441 VTAIL.n62 B 0.020171f
C442 VTAIL.n63 B 0.010839f
C443 VTAIL.n64 B 0.011476f
C444 VTAIL.n65 B 0.025619f
C445 VTAIL.n66 B 0.025619f
C446 VTAIL.n67 B 0.011476f
C447 VTAIL.n68 B 0.010839f
C448 VTAIL.n69 B 0.020171f
C449 VTAIL.n70 B 0.020171f
C450 VTAIL.n71 B 0.010839f
C451 VTAIL.n72 B 0.010839f
C452 VTAIL.n73 B 0.011476f
C453 VTAIL.n74 B 0.025619f
C454 VTAIL.n75 B 0.025619f
C455 VTAIL.n76 B 0.025619f
C456 VTAIL.n77 B 0.011158f
C457 VTAIL.n78 B 0.010839f
C458 VTAIL.n79 B 0.020171f
C459 VTAIL.n80 B 0.020171f
C460 VTAIL.n81 B 0.010839f
C461 VTAIL.n82 B 0.011476f
C462 VTAIL.n83 B 0.025619f
C463 VTAIL.n84 B 0.053776f
C464 VTAIL.n85 B 0.011476f
C465 VTAIL.n86 B 0.010839f
C466 VTAIL.n87 B 0.048001f
C467 VTAIL.n88 B 0.029959f
C468 VTAIL.n89 B 1.70283f
C469 VTAIL.n90 B 0.027399f
C470 VTAIL.n91 B 0.020171f
C471 VTAIL.n92 B 0.010839f
C472 VTAIL.n93 B 0.025619f
C473 VTAIL.n94 B 0.011476f
C474 VTAIL.n95 B 0.020171f
C475 VTAIL.n96 B 0.011158f
C476 VTAIL.n97 B 0.025619f
C477 VTAIL.n98 B 0.010839f
C478 VTAIL.n99 B 0.011476f
C479 VTAIL.n100 B 0.020171f
C480 VTAIL.n101 B 0.010839f
C481 VTAIL.n102 B 0.025619f
C482 VTAIL.n103 B 0.011476f
C483 VTAIL.n104 B 0.020171f
C484 VTAIL.n105 B 0.010839f
C485 VTAIL.n106 B 0.025619f
C486 VTAIL.n107 B 0.011476f
C487 VTAIL.n108 B 0.020171f
C488 VTAIL.n109 B 0.010839f
C489 VTAIL.n110 B 0.025619f
C490 VTAIL.n111 B 0.011476f
C491 VTAIL.n112 B 0.020171f
C492 VTAIL.n113 B 0.010839f
C493 VTAIL.n114 B 0.025619f
C494 VTAIL.n115 B 0.011476f
C495 VTAIL.n116 B 0.020171f
C496 VTAIL.n117 B 0.010839f
C497 VTAIL.n118 B 0.019214f
C498 VTAIL.n119 B 0.015134f
C499 VTAIL.t1 B 0.042321f
C500 VTAIL.n120 B 0.137272f
C501 VTAIL.n121 B 1.41679f
C502 VTAIL.n122 B 0.010839f
C503 VTAIL.n123 B 0.011476f
C504 VTAIL.n124 B 0.025619f
C505 VTAIL.n125 B 0.025619f
C506 VTAIL.n126 B 0.011476f
C507 VTAIL.n127 B 0.010839f
C508 VTAIL.n128 B 0.020171f
C509 VTAIL.n129 B 0.020171f
C510 VTAIL.n130 B 0.010839f
C511 VTAIL.n131 B 0.011476f
C512 VTAIL.n132 B 0.025619f
C513 VTAIL.n133 B 0.025619f
C514 VTAIL.n134 B 0.011476f
C515 VTAIL.n135 B 0.010839f
C516 VTAIL.n136 B 0.020171f
C517 VTAIL.n137 B 0.020171f
C518 VTAIL.n138 B 0.010839f
C519 VTAIL.n139 B 0.011476f
C520 VTAIL.n140 B 0.025619f
C521 VTAIL.n141 B 0.025619f
C522 VTAIL.n142 B 0.011476f
C523 VTAIL.n143 B 0.010839f
C524 VTAIL.n144 B 0.020171f
C525 VTAIL.n145 B 0.020171f
C526 VTAIL.n146 B 0.010839f
C527 VTAIL.n147 B 0.011476f
C528 VTAIL.n148 B 0.025619f
C529 VTAIL.n149 B 0.025619f
C530 VTAIL.n150 B 0.011476f
C531 VTAIL.n151 B 0.010839f
C532 VTAIL.n152 B 0.020171f
C533 VTAIL.n153 B 0.020171f
C534 VTAIL.n154 B 0.010839f
C535 VTAIL.n155 B 0.011476f
C536 VTAIL.n156 B 0.025619f
C537 VTAIL.n157 B 0.025619f
C538 VTAIL.n158 B 0.011476f
C539 VTAIL.n159 B 0.010839f
C540 VTAIL.n160 B 0.020171f
C541 VTAIL.n161 B 0.020171f
C542 VTAIL.n162 B 0.010839f
C543 VTAIL.n163 B 0.011476f
C544 VTAIL.n164 B 0.025619f
C545 VTAIL.n165 B 0.025619f
C546 VTAIL.n166 B 0.025619f
C547 VTAIL.n167 B 0.011158f
C548 VTAIL.n168 B 0.010839f
C549 VTAIL.n169 B 0.020171f
C550 VTAIL.n170 B 0.020171f
C551 VTAIL.n171 B 0.010839f
C552 VTAIL.n172 B 0.011476f
C553 VTAIL.n173 B 0.025619f
C554 VTAIL.n174 B 0.053776f
C555 VTAIL.n175 B 0.011476f
C556 VTAIL.n176 B 0.010839f
C557 VTAIL.n177 B 0.048001f
C558 VTAIL.n178 B 0.029959f
C559 VTAIL.n179 B 1.75158f
C560 VTAIL.n180 B 0.027399f
C561 VTAIL.n181 B 0.020171f
C562 VTAIL.n182 B 0.010839f
C563 VTAIL.n183 B 0.025619f
C564 VTAIL.n184 B 0.011476f
C565 VTAIL.n185 B 0.020171f
C566 VTAIL.n186 B 0.011158f
C567 VTAIL.n187 B 0.025619f
C568 VTAIL.n188 B 0.010839f
C569 VTAIL.n189 B 0.011476f
C570 VTAIL.n190 B 0.020171f
C571 VTAIL.n191 B 0.010839f
C572 VTAIL.n192 B 0.025619f
C573 VTAIL.n193 B 0.011476f
C574 VTAIL.n194 B 0.020171f
C575 VTAIL.n195 B 0.010839f
C576 VTAIL.n196 B 0.025619f
C577 VTAIL.n197 B 0.011476f
C578 VTAIL.n198 B 0.020171f
C579 VTAIL.n199 B 0.010839f
C580 VTAIL.n200 B 0.025619f
C581 VTAIL.n201 B 0.011476f
C582 VTAIL.n202 B 0.020171f
C583 VTAIL.n203 B 0.010839f
C584 VTAIL.n204 B 0.025619f
C585 VTAIL.n205 B 0.011476f
C586 VTAIL.n206 B 0.020171f
C587 VTAIL.n207 B 0.010839f
C588 VTAIL.n208 B 0.019214f
C589 VTAIL.n209 B 0.015134f
C590 VTAIL.t2 B 0.042321f
C591 VTAIL.n210 B 0.137272f
C592 VTAIL.n211 B 1.41679f
C593 VTAIL.n212 B 0.010839f
C594 VTAIL.n213 B 0.011476f
C595 VTAIL.n214 B 0.025619f
C596 VTAIL.n215 B 0.025619f
C597 VTAIL.n216 B 0.011476f
C598 VTAIL.n217 B 0.010839f
C599 VTAIL.n218 B 0.020171f
C600 VTAIL.n219 B 0.020171f
C601 VTAIL.n220 B 0.010839f
C602 VTAIL.n221 B 0.011476f
C603 VTAIL.n222 B 0.025619f
C604 VTAIL.n223 B 0.025619f
C605 VTAIL.n224 B 0.011476f
C606 VTAIL.n225 B 0.010839f
C607 VTAIL.n226 B 0.020171f
C608 VTAIL.n227 B 0.020171f
C609 VTAIL.n228 B 0.010839f
C610 VTAIL.n229 B 0.011476f
C611 VTAIL.n230 B 0.025619f
C612 VTAIL.n231 B 0.025619f
C613 VTAIL.n232 B 0.011476f
C614 VTAIL.n233 B 0.010839f
C615 VTAIL.n234 B 0.020171f
C616 VTAIL.n235 B 0.020171f
C617 VTAIL.n236 B 0.010839f
C618 VTAIL.n237 B 0.011476f
C619 VTAIL.n238 B 0.025619f
C620 VTAIL.n239 B 0.025619f
C621 VTAIL.n240 B 0.011476f
C622 VTAIL.n241 B 0.010839f
C623 VTAIL.n242 B 0.020171f
C624 VTAIL.n243 B 0.020171f
C625 VTAIL.n244 B 0.010839f
C626 VTAIL.n245 B 0.011476f
C627 VTAIL.n246 B 0.025619f
C628 VTAIL.n247 B 0.025619f
C629 VTAIL.n248 B 0.011476f
C630 VTAIL.n249 B 0.010839f
C631 VTAIL.n250 B 0.020171f
C632 VTAIL.n251 B 0.020171f
C633 VTAIL.n252 B 0.010839f
C634 VTAIL.n253 B 0.011476f
C635 VTAIL.n254 B 0.025619f
C636 VTAIL.n255 B 0.025619f
C637 VTAIL.n256 B 0.025619f
C638 VTAIL.n257 B 0.011158f
C639 VTAIL.n258 B 0.010839f
C640 VTAIL.n259 B 0.020171f
C641 VTAIL.n260 B 0.020171f
C642 VTAIL.n261 B 0.010839f
C643 VTAIL.n262 B 0.011476f
C644 VTAIL.n263 B 0.025619f
C645 VTAIL.n264 B 0.053776f
C646 VTAIL.n265 B 0.011476f
C647 VTAIL.n266 B 0.010839f
C648 VTAIL.n267 B 0.048001f
C649 VTAIL.n268 B 0.029959f
C650 VTAIL.n269 B 1.54146f
C651 VTAIL.n270 B 0.027399f
C652 VTAIL.n271 B 0.020171f
C653 VTAIL.n272 B 0.010839f
C654 VTAIL.n273 B 0.025619f
C655 VTAIL.n274 B 0.011476f
C656 VTAIL.n275 B 0.020171f
C657 VTAIL.n276 B 0.011158f
C658 VTAIL.n277 B 0.025619f
C659 VTAIL.n278 B 0.011476f
C660 VTAIL.n279 B 0.020171f
C661 VTAIL.n280 B 0.010839f
C662 VTAIL.n281 B 0.025619f
C663 VTAIL.n282 B 0.011476f
C664 VTAIL.n283 B 0.020171f
C665 VTAIL.n284 B 0.010839f
C666 VTAIL.n285 B 0.025619f
C667 VTAIL.n286 B 0.011476f
C668 VTAIL.n287 B 0.020171f
C669 VTAIL.n288 B 0.010839f
C670 VTAIL.n289 B 0.025619f
C671 VTAIL.n290 B 0.011476f
C672 VTAIL.n291 B 0.020171f
C673 VTAIL.n292 B 0.010839f
C674 VTAIL.n293 B 0.025619f
C675 VTAIL.n294 B 0.011476f
C676 VTAIL.n295 B 0.020171f
C677 VTAIL.n296 B 0.010839f
C678 VTAIL.n297 B 0.019214f
C679 VTAIL.n298 B 0.015134f
C680 VTAIL.t0 B 0.042321f
C681 VTAIL.n299 B 0.137272f
C682 VTAIL.n300 B 1.41679f
C683 VTAIL.n301 B 0.010839f
C684 VTAIL.n302 B 0.011476f
C685 VTAIL.n303 B 0.025619f
C686 VTAIL.n304 B 0.025619f
C687 VTAIL.n305 B 0.011476f
C688 VTAIL.n306 B 0.010839f
C689 VTAIL.n307 B 0.020171f
C690 VTAIL.n308 B 0.020171f
C691 VTAIL.n309 B 0.010839f
C692 VTAIL.n310 B 0.011476f
C693 VTAIL.n311 B 0.025619f
C694 VTAIL.n312 B 0.025619f
C695 VTAIL.n313 B 0.011476f
C696 VTAIL.n314 B 0.010839f
C697 VTAIL.n315 B 0.020171f
C698 VTAIL.n316 B 0.020171f
C699 VTAIL.n317 B 0.010839f
C700 VTAIL.n318 B 0.011476f
C701 VTAIL.n319 B 0.025619f
C702 VTAIL.n320 B 0.025619f
C703 VTAIL.n321 B 0.011476f
C704 VTAIL.n322 B 0.010839f
C705 VTAIL.n323 B 0.020171f
C706 VTAIL.n324 B 0.020171f
C707 VTAIL.n325 B 0.010839f
C708 VTAIL.n326 B 0.011476f
C709 VTAIL.n327 B 0.025619f
C710 VTAIL.n328 B 0.025619f
C711 VTAIL.n329 B 0.011476f
C712 VTAIL.n330 B 0.010839f
C713 VTAIL.n331 B 0.020171f
C714 VTAIL.n332 B 0.020171f
C715 VTAIL.n333 B 0.010839f
C716 VTAIL.n334 B 0.011476f
C717 VTAIL.n335 B 0.025619f
C718 VTAIL.n336 B 0.025619f
C719 VTAIL.n337 B 0.011476f
C720 VTAIL.n338 B 0.010839f
C721 VTAIL.n339 B 0.020171f
C722 VTAIL.n340 B 0.020171f
C723 VTAIL.n341 B 0.010839f
C724 VTAIL.n342 B 0.010839f
C725 VTAIL.n343 B 0.011476f
C726 VTAIL.n344 B 0.025619f
C727 VTAIL.n345 B 0.025619f
C728 VTAIL.n346 B 0.025619f
C729 VTAIL.n347 B 0.011158f
C730 VTAIL.n348 B 0.010839f
C731 VTAIL.n349 B 0.020171f
C732 VTAIL.n350 B 0.020171f
C733 VTAIL.n351 B 0.010839f
C734 VTAIL.n352 B 0.011476f
C735 VTAIL.n353 B 0.025619f
C736 VTAIL.n354 B 0.053776f
C737 VTAIL.n355 B 0.011476f
C738 VTAIL.n356 B 0.010839f
C739 VTAIL.n357 B 0.048001f
C740 VTAIL.n358 B 0.029959f
C741 VTAIL.n359 B 1.45462f
C742 VP.t0 B 4.89811f
C743 VP.t1 B 4.22867f
C744 VP.n0 B 4.68088f
.ends

