* NGSPICE file created from diff_pair_sample_1197.ext - technology: sky130A

.subckt diff_pair_sample_1197 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=4.1652 ps=22.14 w=10.68 l=3.67
X1 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=0 ps=0 w=10.68 l=3.67
X2 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=0 ps=0 w=10.68 l=3.67
X3 VTAIL.t7 VN.t1 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=1.7622 ps=11.01 w=10.68 l=3.67
X4 VTAIL.t0 VP.t0 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=1.7622 ps=11.01 w=10.68 l=3.67
X5 VDD1.t4 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=4.1652 ps=22.14 w=10.68 l=3.67
X6 VDD1.t3 VP.t2 VTAIL.t11 B.t19 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=1.7622 ps=11.01 w=10.68 l=3.67
X7 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=1.7622 ps=11.01 w=10.68 l=3.67
X8 B.t11 B.t9 B.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=0 ps=0 w=10.68 l=3.67
X9 VDD2.t3 VN.t2 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=4.1652 ps=22.14 w=10.68 l=3.67
X10 VDD2.t2 VN.t3 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=1.7622 ps=11.01 w=10.68 l=3.67
X11 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=0 ps=0 w=10.68 l=3.67
X12 VTAIL.t4 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=1.7622 ps=11.01 w=10.68 l=3.67
X13 VDD2.t1 VN.t4 VTAIL.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=4.1652 pd=22.14 as=1.7622 ps=11.01 w=10.68 l=3.67
X14 VTAIL.t6 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=1.7622 ps=11.01 w=10.68 l=3.67
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.7622 pd=11.01 as=4.1652 ps=22.14 w=10.68 l=3.67
R0 VN.n33 VN.n18 161.3
R1 VN.n32 VN.n31 161.3
R2 VN.n30 VN.n19 161.3
R3 VN.n29 VN.n28 161.3
R4 VN.n27 VN.n20 161.3
R5 VN.n26 VN.n25 161.3
R6 VN.n24 VN.n21 161.3
R7 VN.n15 VN.n0 161.3
R8 VN.n14 VN.n13 161.3
R9 VN.n12 VN.n1 161.3
R10 VN.n11 VN.n10 161.3
R11 VN.n9 VN.n2 161.3
R12 VN.n8 VN.n7 161.3
R13 VN.n6 VN.n3 161.3
R14 VN.n5 VN.t3 102.317
R15 VN.n23 VN.t2 102.317
R16 VN.n16 VN.t0 70.1335
R17 VN.n4 VN.t5 70.1335
R18 VN.n34 VN.t4 70.1335
R19 VN.n22 VN.t1 70.1335
R20 VN.n17 VN.n16 57.7881
R21 VN.n35 VN.n34 57.7881
R22 VN VN.n35 52.1407
R23 VN.n5 VN.n4 50.586
R24 VN.n23 VN.n22 50.586
R25 VN.n10 VN.n9 40.577
R26 VN.n10 VN.n1 40.577
R27 VN.n28 VN.n27 40.577
R28 VN.n28 VN.n19 40.577
R29 VN.n4 VN.n3 24.5923
R30 VN.n8 VN.n3 24.5923
R31 VN.n9 VN.n8 24.5923
R32 VN.n14 VN.n1 24.5923
R33 VN.n15 VN.n14 24.5923
R34 VN.n16 VN.n15 24.5923
R35 VN.n27 VN.n26 24.5923
R36 VN.n26 VN.n21 24.5923
R37 VN.n22 VN.n21 24.5923
R38 VN.n34 VN.n33 24.5923
R39 VN.n33 VN.n32 24.5923
R40 VN.n32 VN.n19 24.5923
R41 VN.n24 VN.n23 2.51557
R42 VN.n6 VN.n5 2.51557
R43 VN.n35 VN.n18 0.417304
R44 VN.n17 VN.n0 0.417304
R45 VN VN.n17 0.394524
R46 VN.n31 VN.n18 0.189894
R47 VN.n31 VN.n30 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n20 0.189894
R50 VN.n25 VN.n20 0.189894
R51 VN.n25 VN.n24 0.189894
R52 VN.n7 VN.n6 0.189894
R53 VN.n7 VN.n2 0.189894
R54 VN.n11 VN.n2 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n13 VN.n12 0.189894
R57 VN.n13 VN.n0 0.189894
R58 VTAIL.n234 VTAIL.n182 289.615
R59 VTAIL.n54 VTAIL.n2 289.615
R60 VTAIL.n176 VTAIL.n124 289.615
R61 VTAIL.n116 VTAIL.n64 289.615
R62 VTAIL.n201 VTAIL.n200 185
R63 VTAIL.n198 VTAIL.n197 185
R64 VTAIL.n207 VTAIL.n206 185
R65 VTAIL.n209 VTAIL.n208 185
R66 VTAIL.n194 VTAIL.n193 185
R67 VTAIL.n215 VTAIL.n214 185
R68 VTAIL.n218 VTAIL.n217 185
R69 VTAIL.n216 VTAIL.n190 185
R70 VTAIL.n223 VTAIL.n189 185
R71 VTAIL.n225 VTAIL.n224 185
R72 VTAIL.n227 VTAIL.n226 185
R73 VTAIL.n186 VTAIL.n185 185
R74 VTAIL.n233 VTAIL.n232 185
R75 VTAIL.n235 VTAIL.n234 185
R76 VTAIL.n21 VTAIL.n20 185
R77 VTAIL.n18 VTAIL.n17 185
R78 VTAIL.n27 VTAIL.n26 185
R79 VTAIL.n29 VTAIL.n28 185
R80 VTAIL.n14 VTAIL.n13 185
R81 VTAIL.n35 VTAIL.n34 185
R82 VTAIL.n38 VTAIL.n37 185
R83 VTAIL.n36 VTAIL.n10 185
R84 VTAIL.n43 VTAIL.n9 185
R85 VTAIL.n45 VTAIL.n44 185
R86 VTAIL.n47 VTAIL.n46 185
R87 VTAIL.n6 VTAIL.n5 185
R88 VTAIL.n53 VTAIL.n52 185
R89 VTAIL.n55 VTAIL.n54 185
R90 VTAIL.n177 VTAIL.n176 185
R91 VTAIL.n175 VTAIL.n174 185
R92 VTAIL.n128 VTAIL.n127 185
R93 VTAIL.n169 VTAIL.n168 185
R94 VTAIL.n167 VTAIL.n166 185
R95 VTAIL.n165 VTAIL.n131 185
R96 VTAIL.n135 VTAIL.n132 185
R97 VTAIL.n160 VTAIL.n159 185
R98 VTAIL.n158 VTAIL.n157 185
R99 VTAIL.n137 VTAIL.n136 185
R100 VTAIL.n152 VTAIL.n151 185
R101 VTAIL.n150 VTAIL.n149 185
R102 VTAIL.n141 VTAIL.n140 185
R103 VTAIL.n144 VTAIL.n143 185
R104 VTAIL.n117 VTAIL.n116 185
R105 VTAIL.n115 VTAIL.n114 185
R106 VTAIL.n68 VTAIL.n67 185
R107 VTAIL.n109 VTAIL.n108 185
R108 VTAIL.n107 VTAIL.n106 185
R109 VTAIL.n105 VTAIL.n71 185
R110 VTAIL.n75 VTAIL.n72 185
R111 VTAIL.n100 VTAIL.n99 185
R112 VTAIL.n98 VTAIL.n97 185
R113 VTAIL.n77 VTAIL.n76 185
R114 VTAIL.n92 VTAIL.n91 185
R115 VTAIL.n90 VTAIL.n89 185
R116 VTAIL.n81 VTAIL.n80 185
R117 VTAIL.n84 VTAIL.n83 185
R118 VTAIL.t8 VTAIL.n199 149.524
R119 VTAIL.t1 VTAIL.n19 149.524
R120 VTAIL.t3 VTAIL.n142 149.524
R121 VTAIL.t10 VTAIL.n82 149.524
R122 VTAIL.n200 VTAIL.n197 104.615
R123 VTAIL.n207 VTAIL.n197 104.615
R124 VTAIL.n208 VTAIL.n207 104.615
R125 VTAIL.n208 VTAIL.n193 104.615
R126 VTAIL.n215 VTAIL.n193 104.615
R127 VTAIL.n217 VTAIL.n215 104.615
R128 VTAIL.n217 VTAIL.n216 104.615
R129 VTAIL.n216 VTAIL.n189 104.615
R130 VTAIL.n225 VTAIL.n189 104.615
R131 VTAIL.n226 VTAIL.n225 104.615
R132 VTAIL.n226 VTAIL.n185 104.615
R133 VTAIL.n233 VTAIL.n185 104.615
R134 VTAIL.n234 VTAIL.n233 104.615
R135 VTAIL.n20 VTAIL.n17 104.615
R136 VTAIL.n27 VTAIL.n17 104.615
R137 VTAIL.n28 VTAIL.n27 104.615
R138 VTAIL.n28 VTAIL.n13 104.615
R139 VTAIL.n35 VTAIL.n13 104.615
R140 VTAIL.n37 VTAIL.n35 104.615
R141 VTAIL.n37 VTAIL.n36 104.615
R142 VTAIL.n36 VTAIL.n9 104.615
R143 VTAIL.n45 VTAIL.n9 104.615
R144 VTAIL.n46 VTAIL.n45 104.615
R145 VTAIL.n46 VTAIL.n5 104.615
R146 VTAIL.n53 VTAIL.n5 104.615
R147 VTAIL.n54 VTAIL.n53 104.615
R148 VTAIL.n176 VTAIL.n175 104.615
R149 VTAIL.n175 VTAIL.n127 104.615
R150 VTAIL.n168 VTAIL.n127 104.615
R151 VTAIL.n168 VTAIL.n167 104.615
R152 VTAIL.n167 VTAIL.n131 104.615
R153 VTAIL.n135 VTAIL.n131 104.615
R154 VTAIL.n159 VTAIL.n135 104.615
R155 VTAIL.n159 VTAIL.n158 104.615
R156 VTAIL.n158 VTAIL.n136 104.615
R157 VTAIL.n151 VTAIL.n136 104.615
R158 VTAIL.n151 VTAIL.n150 104.615
R159 VTAIL.n150 VTAIL.n140 104.615
R160 VTAIL.n143 VTAIL.n140 104.615
R161 VTAIL.n116 VTAIL.n115 104.615
R162 VTAIL.n115 VTAIL.n67 104.615
R163 VTAIL.n108 VTAIL.n67 104.615
R164 VTAIL.n108 VTAIL.n107 104.615
R165 VTAIL.n107 VTAIL.n71 104.615
R166 VTAIL.n75 VTAIL.n71 104.615
R167 VTAIL.n99 VTAIL.n75 104.615
R168 VTAIL.n99 VTAIL.n98 104.615
R169 VTAIL.n98 VTAIL.n76 104.615
R170 VTAIL.n91 VTAIL.n76 104.615
R171 VTAIL.n91 VTAIL.n90 104.615
R172 VTAIL.n90 VTAIL.n80 104.615
R173 VTAIL.n83 VTAIL.n80 104.615
R174 VTAIL.n200 VTAIL.t8 52.3082
R175 VTAIL.n20 VTAIL.t1 52.3082
R176 VTAIL.n143 VTAIL.t3 52.3082
R177 VTAIL.n83 VTAIL.t10 52.3082
R178 VTAIL.n123 VTAIL.n122 45.6615
R179 VTAIL.n63 VTAIL.n62 45.6615
R180 VTAIL.n1 VTAIL.n0 45.6613
R181 VTAIL.n61 VTAIL.n60 45.6613
R182 VTAIL.n239 VTAIL.n238 32.1853
R183 VTAIL.n59 VTAIL.n58 32.1853
R184 VTAIL.n181 VTAIL.n180 32.1853
R185 VTAIL.n121 VTAIL.n120 32.1853
R186 VTAIL.n63 VTAIL.n61 28.4703
R187 VTAIL.n239 VTAIL.n181 25.0221
R188 VTAIL.n224 VTAIL.n223 13.1884
R189 VTAIL.n44 VTAIL.n43 13.1884
R190 VTAIL.n166 VTAIL.n165 13.1884
R191 VTAIL.n106 VTAIL.n105 13.1884
R192 VTAIL.n222 VTAIL.n190 12.8005
R193 VTAIL.n227 VTAIL.n188 12.8005
R194 VTAIL.n42 VTAIL.n10 12.8005
R195 VTAIL.n47 VTAIL.n8 12.8005
R196 VTAIL.n169 VTAIL.n130 12.8005
R197 VTAIL.n164 VTAIL.n132 12.8005
R198 VTAIL.n109 VTAIL.n70 12.8005
R199 VTAIL.n104 VTAIL.n72 12.8005
R200 VTAIL.n219 VTAIL.n218 12.0247
R201 VTAIL.n228 VTAIL.n186 12.0247
R202 VTAIL.n39 VTAIL.n38 12.0247
R203 VTAIL.n48 VTAIL.n6 12.0247
R204 VTAIL.n170 VTAIL.n128 12.0247
R205 VTAIL.n161 VTAIL.n160 12.0247
R206 VTAIL.n110 VTAIL.n68 12.0247
R207 VTAIL.n101 VTAIL.n100 12.0247
R208 VTAIL.n214 VTAIL.n192 11.249
R209 VTAIL.n232 VTAIL.n231 11.249
R210 VTAIL.n34 VTAIL.n12 11.249
R211 VTAIL.n52 VTAIL.n51 11.249
R212 VTAIL.n174 VTAIL.n173 11.249
R213 VTAIL.n157 VTAIL.n134 11.249
R214 VTAIL.n114 VTAIL.n113 11.249
R215 VTAIL.n97 VTAIL.n74 11.249
R216 VTAIL.n213 VTAIL.n194 10.4732
R217 VTAIL.n235 VTAIL.n184 10.4732
R218 VTAIL.n33 VTAIL.n14 10.4732
R219 VTAIL.n55 VTAIL.n4 10.4732
R220 VTAIL.n177 VTAIL.n126 10.4732
R221 VTAIL.n156 VTAIL.n137 10.4732
R222 VTAIL.n117 VTAIL.n66 10.4732
R223 VTAIL.n96 VTAIL.n77 10.4732
R224 VTAIL.n201 VTAIL.n199 10.2747
R225 VTAIL.n21 VTAIL.n19 10.2747
R226 VTAIL.n144 VTAIL.n142 10.2747
R227 VTAIL.n84 VTAIL.n82 10.2747
R228 VTAIL.n210 VTAIL.n209 9.69747
R229 VTAIL.n236 VTAIL.n182 9.69747
R230 VTAIL.n30 VTAIL.n29 9.69747
R231 VTAIL.n56 VTAIL.n2 9.69747
R232 VTAIL.n178 VTAIL.n124 9.69747
R233 VTAIL.n153 VTAIL.n152 9.69747
R234 VTAIL.n118 VTAIL.n64 9.69747
R235 VTAIL.n93 VTAIL.n92 9.69747
R236 VTAIL.n238 VTAIL.n237 9.45567
R237 VTAIL.n58 VTAIL.n57 9.45567
R238 VTAIL.n180 VTAIL.n179 9.45567
R239 VTAIL.n120 VTAIL.n119 9.45567
R240 VTAIL.n237 VTAIL.n236 9.3005
R241 VTAIL.n184 VTAIL.n183 9.3005
R242 VTAIL.n231 VTAIL.n230 9.3005
R243 VTAIL.n229 VTAIL.n228 9.3005
R244 VTAIL.n188 VTAIL.n187 9.3005
R245 VTAIL.n203 VTAIL.n202 9.3005
R246 VTAIL.n205 VTAIL.n204 9.3005
R247 VTAIL.n196 VTAIL.n195 9.3005
R248 VTAIL.n211 VTAIL.n210 9.3005
R249 VTAIL.n213 VTAIL.n212 9.3005
R250 VTAIL.n192 VTAIL.n191 9.3005
R251 VTAIL.n220 VTAIL.n219 9.3005
R252 VTAIL.n222 VTAIL.n221 9.3005
R253 VTAIL.n57 VTAIL.n56 9.3005
R254 VTAIL.n4 VTAIL.n3 9.3005
R255 VTAIL.n51 VTAIL.n50 9.3005
R256 VTAIL.n49 VTAIL.n48 9.3005
R257 VTAIL.n8 VTAIL.n7 9.3005
R258 VTAIL.n23 VTAIL.n22 9.3005
R259 VTAIL.n25 VTAIL.n24 9.3005
R260 VTAIL.n16 VTAIL.n15 9.3005
R261 VTAIL.n31 VTAIL.n30 9.3005
R262 VTAIL.n33 VTAIL.n32 9.3005
R263 VTAIL.n12 VTAIL.n11 9.3005
R264 VTAIL.n40 VTAIL.n39 9.3005
R265 VTAIL.n42 VTAIL.n41 9.3005
R266 VTAIL.n146 VTAIL.n145 9.3005
R267 VTAIL.n148 VTAIL.n147 9.3005
R268 VTAIL.n139 VTAIL.n138 9.3005
R269 VTAIL.n154 VTAIL.n153 9.3005
R270 VTAIL.n156 VTAIL.n155 9.3005
R271 VTAIL.n134 VTAIL.n133 9.3005
R272 VTAIL.n162 VTAIL.n161 9.3005
R273 VTAIL.n164 VTAIL.n163 9.3005
R274 VTAIL.n179 VTAIL.n178 9.3005
R275 VTAIL.n126 VTAIL.n125 9.3005
R276 VTAIL.n173 VTAIL.n172 9.3005
R277 VTAIL.n171 VTAIL.n170 9.3005
R278 VTAIL.n130 VTAIL.n129 9.3005
R279 VTAIL.n86 VTAIL.n85 9.3005
R280 VTAIL.n88 VTAIL.n87 9.3005
R281 VTAIL.n79 VTAIL.n78 9.3005
R282 VTAIL.n94 VTAIL.n93 9.3005
R283 VTAIL.n96 VTAIL.n95 9.3005
R284 VTAIL.n74 VTAIL.n73 9.3005
R285 VTAIL.n102 VTAIL.n101 9.3005
R286 VTAIL.n104 VTAIL.n103 9.3005
R287 VTAIL.n119 VTAIL.n118 9.3005
R288 VTAIL.n66 VTAIL.n65 9.3005
R289 VTAIL.n113 VTAIL.n112 9.3005
R290 VTAIL.n111 VTAIL.n110 9.3005
R291 VTAIL.n70 VTAIL.n69 9.3005
R292 VTAIL.n206 VTAIL.n196 8.92171
R293 VTAIL.n26 VTAIL.n16 8.92171
R294 VTAIL.n149 VTAIL.n139 8.92171
R295 VTAIL.n89 VTAIL.n79 8.92171
R296 VTAIL.n205 VTAIL.n198 8.14595
R297 VTAIL.n25 VTAIL.n18 8.14595
R298 VTAIL.n148 VTAIL.n141 8.14595
R299 VTAIL.n88 VTAIL.n81 8.14595
R300 VTAIL.n202 VTAIL.n201 7.3702
R301 VTAIL.n22 VTAIL.n21 7.3702
R302 VTAIL.n145 VTAIL.n144 7.3702
R303 VTAIL.n85 VTAIL.n84 7.3702
R304 VTAIL.n202 VTAIL.n198 5.81868
R305 VTAIL.n22 VTAIL.n18 5.81868
R306 VTAIL.n145 VTAIL.n141 5.81868
R307 VTAIL.n85 VTAIL.n81 5.81868
R308 VTAIL.n206 VTAIL.n205 5.04292
R309 VTAIL.n26 VTAIL.n25 5.04292
R310 VTAIL.n149 VTAIL.n148 5.04292
R311 VTAIL.n89 VTAIL.n88 5.04292
R312 VTAIL.n209 VTAIL.n196 4.26717
R313 VTAIL.n238 VTAIL.n182 4.26717
R314 VTAIL.n29 VTAIL.n16 4.26717
R315 VTAIL.n58 VTAIL.n2 4.26717
R316 VTAIL.n180 VTAIL.n124 4.26717
R317 VTAIL.n152 VTAIL.n139 4.26717
R318 VTAIL.n120 VTAIL.n64 4.26717
R319 VTAIL.n92 VTAIL.n79 4.26717
R320 VTAIL.n210 VTAIL.n194 3.49141
R321 VTAIL.n236 VTAIL.n235 3.49141
R322 VTAIL.n30 VTAIL.n14 3.49141
R323 VTAIL.n56 VTAIL.n55 3.49141
R324 VTAIL.n178 VTAIL.n177 3.49141
R325 VTAIL.n153 VTAIL.n137 3.49141
R326 VTAIL.n118 VTAIL.n117 3.49141
R327 VTAIL.n93 VTAIL.n77 3.49141
R328 VTAIL.n121 VTAIL.n63 3.44878
R329 VTAIL.n181 VTAIL.n123 3.44878
R330 VTAIL.n61 VTAIL.n59 3.44878
R331 VTAIL.n203 VTAIL.n199 2.84303
R332 VTAIL.n23 VTAIL.n19 2.84303
R333 VTAIL.n146 VTAIL.n142 2.84303
R334 VTAIL.n86 VTAIL.n82 2.84303
R335 VTAIL.n214 VTAIL.n213 2.71565
R336 VTAIL.n232 VTAIL.n184 2.71565
R337 VTAIL.n34 VTAIL.n33 2.71565
R338 VTAIL.n52 VTAIL.n4 2.71565
R339 VTAIL.n174 VTAIL.n126 2.71565
R340 VTAIL.n157 VTAIL.n156 2.71565
R341 VTAIL.n114 VTAIL.n66 2.71565
R342 VTAIL.n97 VTAIL.n96 2.71565
R343 VTAIL VTAIL.n239 2.52852
R344 VTAIL.n123 VTAIL.n121 2.19447
R345 VTAIL.n59 VTAIL.n1 2.19447
R346 VTAIL.n218 VTAIL.n192 1.93989
R347 VTAIL.n231 VTAIL.n186 1.93989
R348 VTAIL.n38 VTAIL.n12 1.93989
R349 VTAIL.n51 VTAIL.n6 1.93989
R350 VTAIL.n173 VTAIL.n128 1.93989
R351 VTAIL.n160 VTAIL.n134 1.93989
R352 VTAIL.n113 VTAIL.n68 1.93989
R353 VTAIL.n100 VTAIL.n74 1.93989
R354 VTAIL.n0 VTAIL.t9 1.85443
R355 VTAIL.n0 VTAIL.t6 1.85443
R356 VTAIL.n60 VTAIL.t11 1.85443
R357 VTAIL.n60 VTAIL.t0 1.85443
R358 VTAIL.n122 VTAIL.t2 1.85443
R359 VTAIL.n122 VTAIL.t4 1.85443
R360 VTAIL.n62 VTAIL.t5 1.85443
R361 VTAIL.n62 VTAIL.t7 1.85443
R362 VTAIL.n219 VTAIL.n190 1.16414
R363 VTAIL.n228 VTAIL.n227 1.16414
R364 VTAIL.n39 VTAIL.n10 1.16414
R365 VTAIL.n48 VTAIL.n47 1.16414
R366 VTAIL.n170 VTAIL.n169 1.16414
R367 VTAIL.n161 VTAIL.n132 1.16414
R368 VTAIL.n110 VTAIL.n109 1.16414
R369 VTAIL.n101 VTAIL.n72 1.16414
R370 VTAIL VTAIL.n1 0.920759
R371 VTAIL.n223 VTAIL.n222 0.388379
R372 VTAIL.n224 VTAIL.n188 0.388379
R373 VTAIL.n43 VTAIL.n42 0.388379
R374 VTAIL.n44 VTAIL.n8 0.388379
R375 VTAIL.n166 VTAIL.n130 0.388379
R376 VTAIL.n165 VTAIL.n164 0.388379
R377 VTAIL.n106 VTAIL.n70 0.388379
R378 VTAIL.n105 VTAIL.n104 0.388379
R379 VTAIL.n204 VTAIL.n203 0.155672
R380 VTAIL.n204 VTAIL.n195 0.155672
R381 VTAIL.n211 VTAIL.n195 0.155672
R382 VTAIL.n212 VTAIL.n211 0.155672
R383 VTAIL.n212 VTAIL.n191 0.155672
R384 VTAIL.n220 VTAIL.n191 0.155672
R385 VTAIL.n221 VTAIL.n220 0.155672
R386 VTAIL.n221 VTAIL.n187 0.155672
R387 VTAIL.n229 VTAIL.n187 0.155672
R388 VTAIL.n230 VTAIL.n229 0.155672
R389 VTAIL.n230 VTAIL.n183 0.155672
R390 VTAIL.n237 VTAIL.n183 0.155672
R391 VTAIL.n24 VTAIL.n23 0.155672
R392 VTAIL.n24 VTAIL.n15 0.155672
R393 VTAIL.n31 VTAIL.n15 0.155672
R394 VTAIL.n32 VTAIL.n31 0.155672
R395 VTAIL.n32 VTAIL.n11 0.155672
R396 VTAIL.n40 VTAIL.n11 0.155672
R397 VTAIL.n41 VTAIL.n40 0.155672
R398 VTAIL.n41 VTAIL.n7 0.155672
R399 VTAIL.n49 VTAIL.n7 0.155672
R400 VTAIL.n50 VTAIL.n49 0.155672
R401 VTAIL.n50 VTAIL.n3 0.155672
R402 VTAIL.n57 VTAIL.n3 0.155672
R403 VTAIL.n179 VTAIL.n125 0.155672
R404 VTAIL.n172 VTAIL.n125 0.155672
R405 VTAIL.n172 VTAIL.n171 0.155672
R406 VTAIL.n171 VTAIL.n129 0.155672
R407 VTAIL.n163 VTAIL.n129 0.155672
R408 VTAIL.n163 VTAIL.n162 0.155672
R409 VTAIL.n162 VTAIL.n133 0.155672
R410 VTAIL.n155 VTAIL.n133 0.155672
R411 VTAIL.n155 VTAIL.n154 0.155672
R412 VTAIL.n154 VTAIL.n138 0.155672
R413 VTAIL.n147 VTAIL.n138 0.155672
R414 VTAIL.n147 VTAIL.n146 0.155672
R415 VTAIL.n119 VTAIL.n65 0.155672
R416 VTAIL.n112 VTAIL.n65 0.155672
R417 VTAIL.n112 VTAIL.n111 0.155672
R418 VTAIL.n111 VTAIL.n69 0.155672
R419 VTAIL.n103 VTAIL.n69 0.155672
R420 VTAIL.n103 VTAIL.n102 0.155672
R421 VTAIL.n102 VTAIL.n73 0.155672
R422 VTAIL.n95 VTAIL.n73 0.155672
R423 VTAIL.n95 VTAIL.n94 0.155672
R424 VTAIL.n94 VTAIL.n78 0.155672
R425 VTAIL.n87 VTAIL.n78 0.155672
R426 VTAIL.n87 VTAIL.n86 0.155672
R427 VDD2.n111 VDD2.n59 289.615
R428 VDD2.n52 VDD2.n0 289.615
R429 VDD2.n112 VDD2.n111 185
R430 VDD2.n110 VDD2.n109 185
R431 VDD2.n63 VDD2.n62 185
R432 VDD2.n104 VDD2.n103 185
R433 VDD2.n102 VDD2.n101 185
R434 VDD2.n100 VDD2.n66 185
R435 VDD2.n70 VDD2.n67 185
R436 VDD2.n95 VDD2.n94 185
R437 VDD2.n93 VDD2.n92 185
R438 VDD2.n72 VDD2.n71 185
R439 VDD2.n87 VDD2.n86 185
R440 VDD2.n85 VDD2.n84 185
R441 VDD2.n76 VDD2.n75 185
R442 VDD2.n79 VDD2.n78 185
R443 VDD2.n19 VDD2.n18 185
R444 VDD2.n16 VDD2.n15 185
R445 VDD2.n25 VDD2.n24 185
R446 VDD2.n27 VDD2.n26 185
R447 VDD2.n12 VDD2.n11 185
R448 VDD2.n33 VDD2.n32 185
R449 VDD2.n36 VDD2.n35 185
R450 VDD2.n34 VDD2.n8 185
R451 VDD2.n41 VDD2.n7 185
R452 VDD2.n43 VDD2.n42 185
R453 VDD2.n45 VDD2.n44 185
R454 VDD2.n4 VDD2.n3 185
R455 VDD2.n51 VDD2.n50 185
R456 VDD2.n53 VDD2.n52 185
R457 VDD2.t1 VDD2.n77 149.524
R458 VDD2.t2 VDD2.n17 149.524
R459 VDD2.n111 VDD2.n110 104.615
R460 VDD2.n110 VDD2.n62 104.615
R461 VDD2.n103 VDD2.n62 104.615
R462 VDD2.n103 VDD2.n102 104.615
R463 VDD2.n102 VDD2.n66 104.615
R464 VDD2.n70 VDD2.n66 104.615
R465 VDD2.n94 VDD2.n70 104.615
R466 VDD2.n94 VDD2.n93 104.615
R467 VDD2.n93 VDD2.n71 104.615
R468 VDD2.n86 VDD2.n71 104.615
R469 VDD2.n86 VDD2.n85 104.615
R470 VDD2.n85 VDD2.n75 104.615
R471 VDD2.n78 VDD2.n75 104.615
R472 VDD2.n18 VDD2.n15 104.615
R473 VDD2.n25 VDD2.n15 104.615
R474 VDD2.n26 VDD2.n25 104.615
R475 VDD2.n26 VDD2.n11 104.615
R476 VDD2.n33 VDD2.n11 104.615
R477 VDD2.n35 VDD2.n33 104.615
R478 VDD2.n35 VDD2.n34 104.615
R479 VDD2.n34 VDD2.n7 104.615
R480 VDD2.n43 VDD2.n7 104.615
R481 VDD2.n44 VDD2.n43 104.615
R482 VDD2.n44 VDD2.n3 104.615
R483 VDD2.n51 VDD2.n3 104.615
R484 VDD2.n52 VDD2.n51 104.615
R485 VDD2.n58 VDD2.n57 63.1468
R486 VDD2 VDD2.n117 63.144
R487 VDD2.n78 VDD2.t1 52.3082
R488 VDD2.n18 VDD2.t2 52.3082
R489 VDD2.n58 VDD2.n56 51.395
R490 VDD2.n116 VDD2.n115 48.8641
R491 VDD2.n116 VDD2.n58 44.1291
R492 VDD2.n101 VDD2.n100 13.1884
R493 VDD2.n42 VDD2.n41 13.1884
R494 VDD2.n104 VDD2.n65 12.8005
R495 VDD2.n99 VDD2.n67 12.8005
R496 VDD2.n40 VDD2.n8 12.8005
R497 VDD2.n45 VDD2.n6 12.8005
R498 VDD2.n105 VDD2.n63 12.0247
R499 VDD2.n96 VDD2.n95 12.0247
R500 VDD2.n37 VDD2.n36 12.0247
R501 VDD2.n46 VDD2.n4 12.0247
R502 VDD2.n109 VDD2.n108 11.249
R503 VDD2.n92 VDD2.n69 11.249
R504 VDD2.n32 VDD2.n10 11.249
R505 VDD2.n50 VDD2.n49 11.249
R506 VDD2.n112 VDD2.n61 10.4732
R507 VDD2.n91 VDD2.n72 10.4732
R508 VDD2.n31 VDD2.n12 10.4732
R509 VDD2.n53 VDD2.n2 10.4732
R510 VDD2.n79 VDD2.n77 10.2747
R511 VDD2.n19 VDD2.n17 10.2747
R512 VDD2.n113 VDD2.n59 9.69747
R513 VDD2.n88 VDD2.n87 9.69747
R514 VDD2.n28 VDD2.n27 9.69747
R515 VDD2.n54 VDD2.n0 9.69747
R516 VDD2.n115 VDD2.n114 9.45567
R517 VDD2.n56 VDD2.n55 9.45567
R518 VDD2.n81 VDD2.n80 9.3005
R519 VDD2.n83 VDD2.n82 9.3005
R520 VDD2.n74 VDD2.n73 9.3005
R521 VDD2.n89 VDD2.n88 9.3005
R522 VDD2.n91 VDD2.n90 9.3005
R523 VDD2.n69 VDD2.n68 9.3005
R524 VDD2.n97 VDD2.n96 9.3005
R525 VDD2.n99 VDD2.n98 9.3005
R526 VDD2.n114 VDD2.n113 9.3005
R527 VDD2.n61 VDD2.n60 9.3005
R528 VDD2.n108 VDD2.n107 9.3005
R529 VDD2.n106 VDD2.n105 9.3005
R530 VDD2.n65 VDD2.n64 9.3005
R531 VDD2.n55 VDD2.n54 9.3005
R532 VDD2.n2 VDD2.n1 9.3005
R533 VDD2.n49 VDD2.n48 9.3005
R534 VDD2.n47 VDD2.n46 9.3005
R535 VDD2.n6 VDD2.n5 9.3005
R536 VDD2.n21 VDD2.n20 9.3005
R537 VDD2.n23 VDD2.n22 9.3005
R538 VDD2.n14 VDD2.n13 9.3005
R539 VDD2.n29 VDD2.n28 9.3005
R540 VDD2.n31 VDD2.n30 9.3005
R541 VDD2.n10 VDD2.n9 9.3005
R542 VDD2.n38 VDD2.n37 9.3005
R543 VDD2.n40 VDD2.n39 9.3005
R544 VDD2.n84 VDD2.n74 8.92171
R545 VDD2.n24 VDD2.n14 8.92171
R546 VDD2.n83 VDD2.n76 8.14595
R547 VDD2.n23 VDD2.n16 8.14595
R548 VDD2.n80 VDD2.n79 7.3702
R549 VDD2.n20 VDD2.n19 7.3702
R550 VDD2.n80 VDD2.n76 5.81868
R551 VDD2.n20 VDD2.n16 5.81868
R552 VDD2.n84 VDD2.n83 5.04292
R553 VDD2.n24 VDD2.n23 5.04292
R554 VDD2.n115 VDD2.n59 4.26717
R555 VDD2.n87 VDD2.n74 4.26717
R556 VDD2.n27 VDD2.n14 4.26717
R557 VDD2.n56 VDD2.n0 4.26717
R558 VDD2.n113 VDD2.n112 3.49141
R559 VDD2.n88 VDD2.n72 3.49141
R560 VDD2.n28 VDD2.n12 3.49141
R561 VDD2.n54 VDD2.n53 3.49141
R562 VDD2.n81 VDD2.n77 2.84303
R563 VDD2.n21 VDD2.n17 2.84303
R564 VDD2.n109 VDD2.n61 2.71565
R565 VDD2.n92 VDD2.n91 2.71565
R566 VDD2.n32 VDD2.n31 2.71565
R567 VDD2.n50 VDD2.n2 2.71565
R568 VDD2 VDD2.n116 2.6449
R569 VDD2.n108 VDD2.n63 1.93989
R570 VDD2.n95 VDD2.n69 1.93989
R571 VDD2.n36 VDD2.n10 1.93989
R572 VDD2.n49 VDD2.n4 1.93989
R573 VDD2.n117 VDD2.t4 1.85443
R574 VDD2.n117 VDD2.t3 1.85443
R575 VDD2.n57 VDD2.t0 1.85443
R576 VDD2.n57 VDD2.t5 1.85443
R577 VDD2.n105 VDD2.n104 1.16414
R578 VDD2.n96 VDD2.n67 1.16414
R579 VDD2.n37 VDD2.n8 1.16414
R580 VDD2.n46 VDD2.n45 1.16414
R581 VDD2.n101 VDD2.n65 0.388379
R582 VDD2.n100 VDD2.n99 0.388379
R583 VDD2.n41 VDD2.n40 0.388379
R584 VDD2.n42 VDD2.n6 0.388379
R585 VDD2.n114 VDD2.n60 0.155672
R586 VDD2.n107 VDD2.n60 0.155672
R587 VDD2.n107 VDD2.n106 0.155672
R588 VDD2.n106 VDD2.n64 0.155672
R589 VDD2.n98 VDD2.n64 0.155672
R590 VDD2.n98 VDD2.n97 0.155672
R591 VDD2.n97 VDD2.n68 0.155672
R592 VDD2.n90 VDD2.n68 0.155672
R593 VDD2.n90 VDD2.n89 0.155672
R594 VDD2.n89 VDD2.n73 0.155672
R595 VDD2.n82 VDD2.n73 0.155672
R596 VDD2.n82 VDD2.n81 0.155672
R597 VDD2.n22 VDD2.n21 0.155672
R598 VDD2.n22 VDD2.n13 0.155672
R599 VDD2.n29 VDD2.n13 0.155672
R600 VDD2.n30 VDD2.n29 0.155672
R601 VDD2.n30 VDD2.n9 0.155672
R602 VDD2.n38 VDD2.n9 0.155672
R603 VDD2.n39 VDD2.n38 0.155672
R604 VDD2.n39 VDD2.n5 0.155672
R605 VDD2.n47 VDD2.n5 0.155672
R606 VDD2.n48 VDD2.n47 0.155672
R607 VDD2.n48 VDD2.n1 0.155672
R608 VDD2.n55 VDD2.n1 0.155672
R609 B.n876 B.n875 585
R610 B.n877 B.n876 585
R611 B.n314 B.n144 585
R612 B.n313 B.n312 585
R613 B.n311 B.n310 585
R614 B.n309 B.n308 585
R615 B.n307 B.n306 585
R616 B.n305 B.n304 585
R617 B.n303 B.n302 585
R618 B.n301 B.n300 585
R619 B.n299 B.n298 585
R620 B.n297 B.n296 585
R621 B.n295 B.n294 585
R622 B.n293 B.n292 585
R623 B.n291 B.n290 585
R624 B.n289 B.n288 585
R625 B.n287 B.n286 585
R626 B.n285 B.n284 585
R627 B.n283 B.n282 585
R628 B.n281 B.n280 585
R629 B.n279 B.n278 585
R630 B.n277 B.n276 585
R631 B.n275 B.n274 585
R632 B.n273 B.n272 585
R633 B.n271 B.n270 585
R634 B.n269 B.n268 585
R635 B.n267 B.n266 585
R636 B.n265 B.n264 585
R637 B.n263 B.n262 585
R638 B.n261 B.n260 585
R639 B.n259 B.n258 585
R640 B.n257 B.n256 585
R641 B.n255 B.n254 585
R642 B.n253 B.n252 585
R643 B.n251 B.n250 585
R644 B.n249 B.n248 585
R645 B.n247 B.n246 585
R646 B.n245 B.n244 585
R647 B.n243 B.n242 585
R648 B.n240 B.n239 585
R649 B.n238 B.n237 585
R650 B.n236 B.n235 585
R651 B.n234 B.n233 585
R652 B.n232 B.n231 585
R653 B.n230 B.n229 585
R654 B.n228 B.n227 585
R655 B.n226 B.n225 585
R656 B.n224 B.n223 585
R657 B.n222 B.n221 585
R658 B.n220 B.n219 585
R659 B.n218 B.n217 585
R660 B.n216 B.n215 585
R661 B.n214 B.n213 585
R662 B.n212 B.n211 585
R663 B.n210 B.n209 585
R664 B.n208 B.n207 585
R665 B.n206 B.n205 585
R666 B.n204 B.n203 585
R667 B.n202 B.n201 585
R668 B.n200 B.n199 585
R669 B.n198 B.n197 585
R670 B.n196 B.n195 585
R671 B.n194 B.n193 585
R672 B.n192 B.n191 585
R673 B.n190 B.n189 585
R674 B.n188 B.n187 585
R675 B.n186 B.n185 585
R676 B.n184 B.n183 585
R677 B.n182 B.n181 585
R678 B.n180 B.n179 585
R679 B.n178 B.n177 585
R680 B.n176 B.n175 585
R681 B.n174 B.n173 585
R682 B.n172 B.n171 585
R683 B.n170 B.n169 585
R684 B.n168 B.n167 585
R685 B.n166 B.n165 585
R686 B.n164 B.n163 585
R687 B.n162 B.n161 585
R688 B.n160 B.n159 585
R689 B.n158 B.n157 585
R690 B.n156 B.n155 585
R691 B.n154 B.n153 585
R692 B.n152 B.n151 585
R693 B.n102 B.n101 585
R694 B.n880 B.n879 585
R695 B.n874 B.n145 585
R696 B.n145 B.n99 585
R697 B.n873 B.n98 585
R698 B.n884 B.n98 585
R699 B.n872 B.n97 585
R700 B.n885 B.n97 585
R701 B.n871 B.n96 585
R702 B.n886 B.n96 585
R703 B.n870 B.n869 585
R704 B.n869 B.n92 585
R705 B.n868 B.n91 585
R706 B.n892 B.n91 585
R707 B.n867 B.n90 585
R708 B.n893 B.n90 585
R709 B.n866 B.n89 585
R710 B.n894 B.n89 585
R711 B.n865 B.n864 585
R712 B.n864 B.n85 585
R713 B.n863 B.n84 585
R714 B.n900 B.n84 585
R715 B.n862 B.n83 585
R716 B.n901 B.n83 585
R717 B.n861 B.n82 585
R718 B.n902 B.n82 585
R719 B.n860 B.n859 585
R720 B.n859 B.n78 585
R721 B.n858 B.n77 585
R722 B.n908 B.n77 585
R723 B.n857 B.n76 585
R724 B.n909 B.n76 585
R725 B.n856 B.n75 585
R726 B.n910 B.n75 585
R727 B.n855 B.n854 585
R728 B.n854 B.n71 585
R729 B.n853 B.n70 585
R730 B.n916 B.n70 585
R731 B.n852 B.n69 585
R732 B.n917 B.n69 585
R733 B.n851 B.n68 585
R734 B.n918 B.n68 585
R735 B.n850 B.n849 585
R736 B.n849 B.n64 585
R737 B.n848 B.n63 585
R738 B.n924 B.n63 585
R739 B.n847 B.n62 585
R740 B.n925 B.n62 585
R741 B.n846 B.n61 585
R742 B.n926 B.n61 585
R743 B.n845 B.n844 585
R744 B.n844 B.n57 585
R745 B.n843 B.n56 585
R746 B.n932 B.n56 585
R747 B.n842 B.n55 585
R748 B.n933 B.n55 585
R749 B.n841 B.n54 585
R750 B.n934 B.n54 585
R751 B.n840 B.n839 585
R752 B.n839 B.n50 585
R753 B.n838 B.n49 585
R754 B.n940 B.n49 585
R755 B.n837 B.n48 585
R756 B.n941 B.n48 585
R757 B.n836 B.n47 585
R758 B.n942 B.n47 585
R759 B.n835 B.n834 585
R760 B.n834 B.n43 585
R761 B.n833 B.n42 585
R762 B.n948 B.n42 585
R763 B.n832 B.n41 585
R764 B.n949 B.n41 585
R765 B.n831 B.n40 585
R766 B.n950 B.n40 585
R767 B.n830 B.n829 585
R768 B.n829 B.n36 585
R769 B.n828 B.n35 585
R770 B.n956 B.n35 585
R771 B.n827 B.n34 585
R772 B.n957 B.n34 585
R773 B.n826 B.n33 585
R774 B.n958 B.n33 585
R775 B.n825 B.n824 585
R776 B.n824 B.n29 585
R777 B.n823 B.n28 585
R778 B.n964 B.n28 585
R779 B.n822 B.n27 585
R780 B.n965 B.n27 585
R781 B.n821 B.n26 585
R782 B.n966 B.n26 585
R783 B.n820 B.n819 585
R784 B.n819 B.n22 585
R785 B.n818 B.n21 585
R786 B.n972 B.n21 585
R787 B.n817 B.n20 585
R788 B.n973 B.n20 585
R789 B.n816 B.n19 585
R790 B.n974 B.n19 585
R791 B.n815 B.n814 585
R792 B.n814 B.n15 585
R793 B.n813 B.n14 585
R794 B.n980 B.n14 585
R795 B.n812 B.n13 585
R796 B.n981 B.n13 585
R797 B.n811 B.n12 585
R798 B.n982 B.n12 585
R799 B.n810 B.n809 585
R800 B.n809 B.n8 585
R801 B.n808 B.n7 585
R802 B.n988 B.n7 585
R803 B.n807 B.n6 585
R804 B.n989 B.n6 585
R805 B.n806 B.n5 585
R806 B.n990 B.n5 585
R807 B.n805 B.n804 585
R808 B.n804 B.n4 585
R809 B.n803 B.n315 585
R810 B.n803 B.n802 585
R811 B.n793 B.n316 585
R812 B.n317 B.n316 585
R813 B.n795 B.n794 585
R814 B.n796 B.n795 585
R815 B.n792 B.n322 585
R816 B.n322 B.n321 585
R817 B.n791 B.n790 585
R818 B.n790 B.n789 585
R819 B.n324 B.n323 585
R820 B.n325 B.n324 585
R821 B.n782 B.n781 585
R822 B.n783 B.n782 585
R823 B.n780 B.n330 585
R824 B.n330 B.n329 585
R825 B.n779 B.n778 585
R826 B.n778 B.n777 585
R827 B.n332 B.n331 585
R828 B.n333 B.n332 585
R829 B.n770 B.n769 585
R830 B.n771 B.n770 585
R831 B.n768 B.n338 585
R832 B.n338 B.n337 585
R833 B.n767 B.n766 585
R834 B.n766 B.n765 585
R835 B.n340 B.n339 585
R836 B.n341 B.n340 585
R837 B.n758 B.n757 585
R838 B.n759 B.n758 585
R839 B.n756 B.n346 585
R840 B.n346 B.n345 585
R841 B.n755 B.n754 585
R842 B.n754 B.n753 585
R843 B.n348 B.n347 585
R844 B.n349 B.n348 585
R845 B.n746 B.n745 585
R846 B.n747 B.n746 585
R847 B.n744 B.n354 585
R848 B.n354 B.n353 585
R849 B.n743 B.n742 585
R850 B.n742 B.n741 585
R851 B.n356 B.n355 585
R852 B.n357 B.n356 585
R853 B.n734 B.n733 585
R854 B.n735 B.n734 585
R855 B.n732 B.n362 585
R856 B.n362 B.n361 585
R857 B.n731 B.n730 585
R858 B.n730 B.n729 585
R859 B.n364 B.n363 585
R860 B.n365 B.n364 585
R861 B.n722 B.n721 585
R862 B.n723 B.n722 585
R863 B.n720 B.n370 585
R864 B.n370 B.n369 585
R865 B.n719 B.n718 585
R866 B.n718 B.n717 585
R867 B.n372 B.n371 585
R868 B.n373 B.n372 585
R869 B.n710 B.n709 585
R870 B.n711 B.n710 585
R871 B.n708 B.n378 585
R872 B.n378 B.n377 585
R873 B.n707 B.n706 585
R874 B.n706 B.n705 585
R875 B.n380 B.n379 585
R876 B.n381 B.n380 585
R877 B.n698 B.n697 585
R878 B.n699 B.n698 585
R879 B.n696 B.n386 585
R880 B.n386 B.n385 585
R881 B.n695 B.n694 585
R882 B.n694 B.n693 585
R883 B.n388 B.n387 585
R884 B.n389 B.n388 585
R885 B.n686 B.n685 585
R886 B.n687 B.n686 585
R887 B.n684 B.n394 585
R888 B.n394 B.n393 585
R889 B.n683 B.n682 585
R890 B.n682 B.n681 585
R891 B.n396 B.n395 585
R892 B.n397 B.n396 585
R893 B.n674 B.n673 585
R894 B.n675 B.n674 585
R895 B.n672 B.n402 585
R896 B.n402 B.n401 585
R897 B.n671 B.n670 585
R898 B.n670 B.n669 585
R899 B.n404 B.n403 585
R900 B.n405 B.n404 585
R901 B.n662 B.n661 585
R902 B.n663 B.n662 585
R903 B.n660 B.n410 585
R904 B.n410 B.n409 585
R905 B.n659 B.n658 585
R906 B.n658 B.n657 585
R907 B.n412 B.n411 585
R908 B.n413 B.n412 585
R909 B.n650 B.n649 585
R910 B.n651 B.n650 585
R911 B.n648 B.n418 585
R912 B.n418 B.n417 585
R913 B.n647 B.n646 585
R914 B.n646 B.n645 585
R915 B.n420 B.n419 585
R916 B.n421 B.n420 585
R917 B.n641 B.n640 585
R918 B.n424 B.n423 585
R919 B.n637 B.n636 585
R920 B.n638 B.n637 585
R921 B.n635 B.n466 585
R922 B.n634 B.n633 585
R923 B.n632 B.n631 585
R924 B.n630 B.n629 585
R925 B.n628 B.n627 585
R926 B.n626 B.n625 585
R927 B.n624 B.n623 585
R928 B.n622 B.n621 585
R929 B.n620 B.n619 585
R930 B.n618 B.n617 585
R931 B.n616 B.n615 585
R932 B.n614 B.n613 585
R933 B.n612 B.n611 585
R934 B.n610 B.n609 585
R935 B.n608 B.n607 585
R936 B.n606 B.n605 585
R937 B.n604 B.n603 585
R938 B.n602 B.n601 585
R939 B.n600 B.n599 585
R940 B.n598 B.n597 585
R941 B.n596 B.n595 585
R942 B.n594 B.n593 585
R943 B.n592 B.n591 585
R944 B.n590 B.n589 585
R945 B.n588 B.n587 585
R946 B.n586 B.n585 585
R947 B.n584 B.n583 585
R948 B.n582 B.n581 585
R949 B.n580 B.n579 585
R950 B.n578 B.n577 585
R951 B.n576 B.n575 585
R952 B.n574 B.n573 585
R953 B.n572 B.n571 585
R954 B.n570 B.n569 585
R955 B.n568 B.n567 585
R956 B.n565 B.n564 585
R957 B.n563 B.n562 585
R958 B.n561 B.n560 585
R959 B.n559 B.n558 585
R960 B.n557 B.n556 585
R961 B.n555 B.n554 585
R962 B.n553 B.n552 585
R963 B.n551 B.n550 585
R964 B.n549 B.n548 585
R965 B.n547 B.n546 585
R966 B.n545 B.n544 585
R967 B.n543 B.n542 585
R968 B.n541 B.n540 585
R969 B.n539 B.n538 585
R970 B.n537 B.n536 585
R971 B.n535 B.n534 585
R972 B.n533 B.n532 585
R973 B.n531 B.n530 585
R974 B.n529 B.n528 585
R975 B.n527 B.n526 585
R976 B.n525 B.n524 585
R977 B.n523 B.n522 585
R978 B.n521 B.n520 585
R979 B.n519 B.n518 585
R980 B.n517 B.n516 585
R981 B.n515 B.n514 585
R982 B.n513 B.n512 585
R983 B.n511 B.n510 585
R984 B.n509 B.n508 585
R985 B.n507 B.n506 585
R986 B.n505 B.n504 585
R987 B.n503 B.n502 585
R988 B.n501 B.n500 585
R989 B.n499 B.n498 585
R990 B.n497 B.n496 585
R991 B.n495 B.n494 585
R992 B.n493 B.n492 585
R993 B.n491 B.n490 585
R994 B.n489 B.n488 585
R995 B.n487 B.n486 585
R996 B.n485 B.n484 585
R997 B.n483 B.n482 585
R998 B.n481 B.n480 585
R999 B.n479 B.n478 585
R1000 B.n477 B.n476 585
R1001 B.n475 B.n474 585
R1002 B.n473 B.n472 585
R1003 B.n642 B.n422 585
R1004 B.n422 B.n421 585
R1005 B.n644 B.n643 585
R1006 B.n645 B.n644 585
R1007 B.n416 B.n415 585
R1008 B.n417 B.n416 585
R1009 B.n653 B.n652 585
R1010 B.n652 B.n651 585
R1011 B.n654 B.n414 585
R1012 B.n414 B.n413 585
R1013 B.n656 B.n655 585
R1014 B.n657 B.n656 585
R1015 B.n408 B.n407 585
R1016 B.n409 B.n408 585
R1017 B.n665 B.n664 585
R1018 B.n664 B.n663 585
R1019 B.n666 B.n406 585
R1020 B.n406 B.n405 585
R1021 B.n668 B.n667 585
R1022 B.n669 B.n668 585
R1023 B.n400 B.n399 585
R1024 B.n401 B.n400 585
R1025 B.n677 B.n676 585
R1026 B.n676 B.n675 585
R1027 B.n678 B.n398 585
R1028 B.n398 B.n397 585
R1029 B.n680 B.n679 585
R1030 B.n681 B.n680 585
R1031 B.n392 B.n391 585
R1032 B.n393 B.n392 585
R1033 B.n689 B.n688 585
R1034 B.n688 B.n687 585
R1035 B.n690 B.n390 585
R1036 B.n390 B.n389 585
R1037 B.n692 B.n691 585
R1038 B.n693 B.n692 585
R1039 B.n384 B.n383 585
R1040 B.n385 B.n384 585
R1041 B.n701 B.n700 585
R1042 B.n700 B.n699 585
R1043 B.n702 B.n382 585
R1044 B.n382 B.n381 585
R1045 B.n704 B.n703 585
R1046 B.n705 B.n704 585
R1047 B.n376 B.n375 585
R1048 B.n377 B.n376 585
R1049 B.n713 B.n712 585
R1050 B.n712 B.n711 585
R1051 B.n714 B.n374 585
R1052 B.n374 B.n373 585
R1053 B.n716 B.n715 585
R1054 B.n717 B.n716 585
R1055 B.n368 B.n367 585
R1056 B.n369 B.n368 585
R1057 B.n725 B.n724 585
R1058 B.n724 B.n723 585
R1059 B.n726 B.n366 585
R1060 B.n366 B.n365 585
R1061 B.n728 B.n727 585
R1062 B.n729 B.n728 585
R1063 B.n360 B.n359 585
R1064 B.n361 B.n360 585
R1065 B.n737 B.n736 585
R1066 B.n736 B.n735 585
R1067 B.n738 B.n358 585
R1068 B.n358 B.n357 585
R1069 B.n740 B.n739 585
R1070 B.n741 B.n740 585
R1071 B.n352 B.n351 585
R1072 B.n353 B.n352 585
R1073 B.n749 B.n748 585
R1074 B.n748 B.n747 585
R1075 B.n750 B.n350 585
R1076 B.n350 B.n349 585
R1077 B.n752 B.n751 585
R1078 B.n753 B.n752 585
R1079 B.n344 B.n343 585
R1080 B.n345 B.n344 585
R1081 B.n761 B.n760 585
R1082 B.n760 B.n759 585
R1083 B.n762 B.n342 585
R1084 B.n342 B.n341 585
R1085 B.n764 B.n763 585
R1086 B.n765 B.n764 585
R1087 B.n336 B.n335 585
R1088 B.n337 B.n336 585
R1089 B.n773 B.n772 585
R1090 B.n772 B.n771 585
R1091 B.n774 B.n334 585
R1092 B.n334 B.n333 585
R1093 B.n776 B.n775 585
R1094 B.n777 B.n776 585
R1095 B.n328 B.n327 585
R1096 B.n329 B.n328 585
R1097 B.n785 B.n784 585
R1098 B.n784 B.n783 585
R1099 B.n786 B.n326 585
R1100 B.n326 B.n325 585
R1101 B.n788 B.n787 585
R1102 B.n789 B.n788 585
R1103 B.n320 B.n319 585
R1104 B.n321 B.n320 585
R1105 B.n798 B.n797 585
R1106 B.n797 B.n796 585
R1107 B.n799 B.n318 585
R1108 B.n318 B.n317 585
R1109 B.n801 B.n800 585
R1110 B.n802 B.n801 585
R1111 B.n2 B.n0 585
R1112 B.n4 B.n2 585
R1113 B.n3 B.n1 585
R1114 B.n989 B.n3 585
R1115 B.n987 B.n986 585
R1116 B.n988 B.n987 585
R1117 B.n985 B.n9 585
R1118 B.n9 B.n8 585
R1119 B.n984 B.n983 585
R1120 B.n983 B.n982 585
R1121 B.n11 B.n10 585
R1122 B.n981 B.n11 585
R1123 B.n979 B.n978 585
R1124 B.n980 B.n979 585
R1125 B.n977 B.n16 585
R1126 B.n16 B.n15 585
R1127 B.n976 B.n975 585
R1128 B.n975 B.n974 585
R1129 B.n18 B.n17 585
R1130 B.n973 B.n18 585
R1131 B.n971 B.n970 585
R1132 B.n972 B.n971 585
R1133 B.n969 B.n23 585
R1134 B.n23 B.n22 585
R1135 B.n968 B.n967 585
R1136 B.n967 B.n966 585
R1137 B.n25 B.n24 585
R1138 B.n965 B.n25 585
R1139 B.n963 B.n962 585
R1140 B.n964 B.n963 585
R1141 B.n961 B.n30 585
R1142 B.n30 B.n29 585
R1143 B.n960 B.n959 585
R1144 B.n959 B.n958 585
R1145 B.n32 B.n31 585
R1146 B.n957 B.n32 585
R1147 B.n955 B.n954 585
R1148 B.n956 B.n955 585
R1149 B.n953 B.n37 585
R1150 B.n37 B.n36 585
R1151 B.n952 B.n951 585
R1152 B.n951 B.n950 585
R1153 B.n39 B.n38 585
R1154 B.n949 B.n39 585
R1155 B.n947 B.n946 585
R1156 B.n948 B.n947 585
R1157 B.n945 B.n44 585
R1158 B.n44 B.n43 585
R1159 B.n944 B.n943 585
R1160 B.n943 B.n942 585
R1161 B.n46 B.n45 585
R1162 B.n941 B.n46 585
R1163 B.n939 B.n938 585
R1164 B.n940 B.n939 585
R1165 B.n937 B.n51 585
R1166 B.n51 B.n50 585
R1167 B.n936 B.n935 585
R1168 B.n935 B.n934 585
R1169 B.n53 B.n52 585
R1170 B.n933 B.n53 585
R1171 B.n931 B.n930 585
R1172 B.n932 B.n931 585
R1173 B.n929 B.n58 585
R1174 B.n58 B.n57 585
R1175 B.n928 B.n927 585
R1176 B.n927 B.n926 585
R1177 B.n60 B.n59 585
R1178 B.n925 B.n60 585
R1179 B.n923 B.n922 585
R1180 B.n924 B.n923 585
R1181 B.n921 B.n65 585
R1182 B.n65 B.n64 585
R1183 B.n920 B.n919 585
R1184 B.n919 B.n918 585
R1185 B.n67 B.n66 585
R1186 B.n917 B.n67 585
R1187 B.n915 B.n914 585
R1188 B.n916 B.n915 585
R1189 B.n913 B.n72 585
R1190 B.n72 B.n71 585
R1191 B.n912 B.n911 585
R1192 B.n911 B.n910 585
R1193 B.n74 B.n73 585
R1194 B.n909 B.n74 585
R1195 B.n907 B.n906 585
R1196 B.n908 B.n907 585
R1197 B.n905 B.n79 585
R1198 B.n79 B.n78 585
R1199 B.n904 B.n903 585
R1200 B.n903 B.n902 585
R1201 B.n81 B.n80 585
R1202 B.n901 B.n81 585
R1203 B.n899 B.n898 585
R1204 B.n900 B.n899 585
R1205 B.n897 B.n86 585
R1206 B.n86 B.n85 585
R1207 B.n896 B.n895 585
R1208 B.n895 B.n894 585
R1209 B.n88 B.n87 585
R1210 B.n893 B.n88 585
R1211 B.n891 B.n890 585
R1212 B.n892 B.n891 585
R1213 B.n889 B.n93 585
R1214 B.n93 B.n92 585
R1215 B.n888 B.n887 585
R1216 B.n887 B.n886 585
R1217 B.n95 B.n94 585
R1218 B.n885 B.n95 585
R1219 B.n883 B.n882 585
R1220 B.n884 B.n883 585
R1221 B.n881 B.n100 585
R1222 B.n100 B.n99 585
R1223 B.n992 B.n991 585
R1224 B.n991 B.n990 585
R1225 B.n640 B.n422 530.939
R1226 B.n879 B.n100 530.939
R1227 B.n472 B.n420 530.939
R1228 B.n876 B.n145 530.939
R1229 B.n469 B.t11 336.935
R1230 B.n146 B.t14 336.935
R1231 B.n467 B.t8 336.935
R1232 B.n148 B.t17 336.935
R1233 B.n469 B.t9 279.373
R1234 B.n467 B.t5 279.373
R1235 B.n148 B.t16 279.373
R1236 B.n146 B.t12 279.373
R1237 B.n470 B.t10 259.36
R1238 B.n147 B.t15 259.36
R1239 B.n468 B.t7 259.36
R1240 B.n149 B.t18 259.36
R1241 B.n877 B.n143 256.663
R1242 B.n877 B.n142 256.663
R1243 B.n877 B.n141 256.663
R1244 B.n877 B.n140 256.663
R1245 B.n877 B.n139 256.663
R1246 B.n877 B.n138 256.663
R1247 B.n877 B.n137 256.663
R1248 B.n877 B.n136 256.663
R1249 B.n877 B.n135 256.663
R1250 B.n877 B.n134 256.663
R1251 B.n877 B.n133 256.663
R1252 B.n877 B.n132 256.663
R1253 B.n877 B.n131 256.663
R1254 B.n877 B.n130 256.663
R1255 B.n877 B.n129 256.663
R1256 B.n877 B.n128 256.663
R1257 B.n877 B.n127 256.663
R1258 B.n877 B.n126 256.663
R1259 B.n877 B.n125 256.663
R1260 B.n877 B.n124 256.663
R1261 B.n877 B.n123 256.663
R1262 B.n877 B.n122 256.663
R1263 B.n877 B.n121 256.663
R1264 B.n877 B.n120 256.663
R1265 B.n877 B.n119 256.663
R1266 B.n877 B.n118 256.663
R1267 B.n877 B.n117 256.663
R1268 B.n877 B.n116 256.663
R1269 B.n877 B.n115 256.663
R1270 B.n877 B.n114 256.663
R1271 B.n877 B.n113 256.663
R1272 B.n877 B.n112 256.663
R1273 B.n877 B.n111 256.663
R1274 B.n877 B.n110 256.663
R1275 B.n877 B.n109 256.663
R1276 B.n877 B.n108 256.663
R1277 B.n877 B.n107 256.663
R1278 B.n877 B.n106 256.663
R1279 B.n877 B.n105 256.663
R1280 B.n877 B.n104 256.663
R1281 B.n877 B.n103 256.663
R1282 B.n878 B.n877 256.663
R1283 B.n639 B.n638 256.663
R1284 B.n638 B.n425 256.663
R1285 B.n638 B.n426 256.663
R1286 B.n638 B.n427 256.663
R1287 B.n638 B.n428 256.663
R1288 B.n638 B.n429 256.663
R1289 B.n638 B.n430 256.663
R1290 B.n638 B.n431 256.663
R1291 B.n638 B.n432 256.663
R1292 B.n638 B.n433 256.663
R1293 B.n638 B.n434 256.663
R1294 B.n638 B.n435 256.663
R1295 B.n638 B.n436 256.663
R1296 B.n638 B.n437 256.663
R1297 B.n638 B.n438 256.663
R1298 B.n638 B.n439 256.663
R1299 B.n638 B.n440 256.663
R1300 B.n638 B.n441 256.663
R1301 B.n638 B.n442 256.663
R1302 B.n638 B.n443 256.663
R1303 B.n638 B.n444 256.663
R1304 B.n638 B.n445 256.663
R1305 B.n638 B.n446 256.663
R1306 B.n638 B.n447 256.663
R1307 B.n638 B.n448 256.663
R1308 B.n638 B.n449 256.663
R1309 B.n638 B.n450 256.663
R1310 B.n638 B.n451 256.663
R1311 B.n638 B.n452 256.663
R1312 B.n638 B.n453 256.663
R1313 B.n638 B.n454 256.663
R1314 B.n638 B.n455 256.663
R1315 B.n638 B.n456 256.663
R1316 B.n638 B.n457 256.663
R1317 B.n638 B.n458 256.663
R1318 B.n638 B.n459 256.663
R1319 B.n638 B.n460 256.663
R1320 B.n638 B.n461 256.663
R1321 B.n638 B.n462 256.663
R1322 B.n638 B.n463 256.663
R1323 B.n638 B.n464 256.663
R1324 B.n638 B.n465 256.663
R1325 B.n644 B.n422 163.367
R1326 B.n644 B.n416 163.367
R1327 B.n652 B.n416 163.367
R1328 B.n652 B.n414 163.367
R1329 B.n656 B.n414 163.367
R1330 B.n656 B.n408 163.367
R1331 B.n664 B.n408 163.367
R1332 B.n664 B.n406 163.367
R1333 B.n668 B.n406 163.367
R1334 B.n668 B.n400 163.367
R1335 B.n676 B.n400 163.367
R1336 B.n676 B.n398 163.367
R1337 B.n680 B.n398 163.367
R1338 B.n680 B.n392 163.367
R1339 B.n688 B.n392 163.367
R1340 B.n688 B.n390 163.367
R1341 B.n692 B.n390 163.367
R1342 B.n692 B.n384 163.367
R1343 B.n700 B.n384 163.367
R1344 B.n700 B.n382 163.367
R1345 B.n704 B.n382 163.367
R1346 B.n704 B.n376 163.367
R1347 B.n712 B.n376 163.367
R1348 B.n712 B.n374 163.367
R1349 B.n716 B.n374 163.367
R1350 B.n716 B.n368 163.367
R1351 B.n724 B.n368 163.367
R1352 B.n724 B.n366 163.367
R1353 B.n728 B.n366 163.367
R1354 B.n728 B.n360 163.367
R1355 B.n736 B.n360 163.367
R1356 B.n736 B.n358 163.367
R1357 B.n740 B.n358 163.367
R1358 B.n740 B.n352 163.367
R1359 B.n748 B.n352 163.367
R1360 B.n748 B.n350 163.367
R1361 B.n752 B.n350 163.367
R1362 B.n752 B.n344 163.367
R1363 B.n760 B.n344 163.367
R1364 B.n760 B.n342 163.367
R1365 B.n764 B.n342 163.367
R1366 B.n764 B.n336 163.367
R1367 B.n772 B.n336 163.367
R1368 B.n772 B.n334 163.367
R1369 B.n776 B.n334 163.367
R1370 B.n776 B.n328 163.367
R1371 B.n784 B.n328 163.367
R1372 B.n784 B.n326 163.367
R1373 B.n788 B.n326 163.367
R1374 B.n788 B.n320 163.367
R1375 B.n797 B.n320 163.367
R1376 B.n797 B.n318 163.367
R1377 B.n801 B.n318 163.367
R1378 B.n801 B.n2 163.367
R1379 B.n991 B.n2 163.367
R1380 B.n991 B.n3 163.367
R1381 B.n987 B.n3 163.367
R1382 B.n987 B.n9 163.367
R1383 B.n983 B.n9 163.367
R1384 B.n983 B.n11 163.367
R1385 B.n979 B.n11 163.367
R1386 B.n979 B.n16 163.367
R1387 B.n975 B.n16 163.367
R1388 B.n975 B.n18 163.367
R1389 B.n971 B.n18 163.367
R1390 B.n971 B.n23 163.367
R1391 B.n967 B.n23 163.367
R1392 B.n967 B.n25 163.367
R1393 B.n963 B.n25 163.367
R1394 B.n963 B.n30 163.367
R1395 B.n959 B.n30 163.367
R1396 B.n959 B.n32 163.367
R1397 B.n955 B.n32 163.367
R1398 B.n955 B.n37 163.367
R1399 B.n951 B.n37 163.367
R1400 B.n951 B.n39 163.367
R1401 B.n947 B.n39 163.367
R1402 B.n947 B.n44 163.367
R1403 B.n943 B.n44 163.367
R1404 B.n943 B.n46 163.367
R1405 B.n939 B.n46 163.367
R1406 B.n939 B.n51 163.367
R1407 B.n935 B.n51 163.367
R1408 B.n935 B.n53 163.367
R1409 B.n931 B.n53 163.367
R1410 B.n931 B.n58 163.367
R1411 B.n927 B.n58 163.367
R1412 B.n927 B.n60 163.367
R1413 B.n923 B.n60 163.367
R1414 B.n923 B.n65 163.367
R1415 B.n919 B.n65 163.367
R1416 B.n919 B.n67 163.367
R1417 B.n915 B.n67 163.367
R1418 B.n915 B.n72 163.367
R1419 B.n911 B.n72 163.367
R1420 B.n911 B.n74 163.367
R1421 B.n907 B.n74 163.367
R1422 B.n907 B.n79 163.367
R1423 B.n903 B.n79 163.367
R1424 B.n903 B.n81 163.367
R1425 B.n899 B.n81 163.367
R1426 B.n899 B.n86 163.367
R1427 B.n895 B.n86 163.367
R1428 B.n895 B.n88 163.367
R1429 B.n891 B.n88 163.367
R1430 B.n891 B.n93 163.367
R1431 B.n887 B.n93 163.367
R1432 B.n887 B.n95 163.367
R1433 B.n883 B.n95 163.367
R1434 B.n883 B.n100 163.367
R1435 B.n637 B.n424 163.367
R1436 B.n637 B.n466 163.367
R1437 B.n633 B.n632 163.367
R1438 B.n629 B.n628 163.367
R1439 B.n625 B.n624 163.367
R1440 B.n621 B.n620 163.367
R1441 B.n617 B.n616 163.367
R1442 B.n613 B.n612 163.367
R1443 B.n609 B.n608 163.367
R1444 B.n605 B.n604 163.367
R1445 B.n601 B.n600 163.367
R1446 B.n597 B.n596 163.367
R1447 B.n593 B.n592 163.367
R1448 B.n589 B.n588 163.367
R1449 B.n585 B.n584 163.367
R1450 B.n581 B.n580 163.367
R1451 B.n577 B.n576 163.367
R1452 B.n573 B.n572 163.367
R1453 B.n569 B.n568 163.367
R1454 B.n564 B.n563 163.367
R1455 B.n560 B.n559 163.367
R1456 B.n556 B.n555 163.367
R1457 B.n552 B.n551 163.367
R1458 B.n548 B.n547 163.367
R1459 B.n544 B.n543 163.367
R1460 B.n540 B.n539 163.367
R1461 B.n536 B.n535 163.367
R1462 B.n532 B.n531 163.367
R1463 B.n528 B.n527 163.367
R1464 B.n524 B.n523 163.367
R1465 B.n520 B.n519 163.367
R1466 B.n516 B.n515 163.367
R1467 B.n512 B.n511 163.367
R1468 B.n508 B.n507 163.367
R1469 B.n504 B.n503 163.367
R1470 B.n500 B.n499 163.367
R1471 B.n496 B.n495 163.367
R1472 B.n492 B.n491 163.367
R1473 B.n488 B.n487 163.367
R1474 B.n484 B.n483 163.367
R1475 B.n480 B.n479 163.367
R1476 B.n476 B.n475 163.367
R1477 B.n646 B.n420 163.367
R1478 B.n646 B.n418 163.367
R1479 B.n650 B.n418 163.367
R1480 B.n650 B.n412 163.367
R1481 B.n658 B.n412 163.367
R1482 B.n658 B.n410 163.367
R1483 B.n662 B.n410 163.367
R1484 B.n662 B.n404 163.367
R1485 B.n670 B.n404 163.367
R1486 B.n670 B.n402 163.367
R1487 B.n674 B.n402 163.367
R1488 B.n674 B.n396 163.367
R1489 B.n682 B.n396 163.367
R1490 B.n682 B.n394 163.367
R1491 B.n686 B.n394 163.367
R1492 B.n686 B.n388 163.367
R1493 B.n694 B.n388 163.367
R1494 B.n694 B.n386 163.367
R1495 B.n698 B.n386 163.367
R1496 B.n698 B.n380 163.367
R1497 B.n706 B.n380 163.367
R1498 B.n706 B.n378 163.367
R1499 B.n710 B.n378 163.367
R1500 B.n710 B.n372 163.367
R1501 B.n718 B.n372 163.367
R1502 B.n718 B.n370 163.367
R1503 B.n722 B.n370 163.367
R1504 B.n722 B.n364 163.367
R1505 B.n730 B.n364 163.367
R1506 B.n730 B.n362 163.367
R1507 B.n734 B.n362 163.367
R1508 B.n734 B.n356 163.367
R1509 B.n742 B.n356 163.367
R1510 B.n742 B.n354 163.367
R1511 B.n746 B.n354 163.367
R1512 B.n746 B.n348 163.367
R1513 B.n754 B.n348 163.367
R1514 B.n754 B.n346 163.367
R1515 B.n758 B.n346 163.367
R1516 B.n758 B.n340 163.367
R1517 B.n766 B.n340 163.367
R1518 B.n766 B.n338 163.367
R1519 B.n770 B.n338 163.367
R1520 B.n770 B.n332 163.367
R1521 B.n778 B.n332 163.367
R1522 B.n778 B.n330 163.367
R1523 B.n782 B.n330 163.367
R1524 B.n782 B.n324 163.367
R1525 B.n790 B.n324 163.367
R1526 B.n790 B.n322 163.367
R1527 B.n795 B.n322 163.367
R1528 B.n795 B.n316 163.367
R1529 B.n803 B.n316 163.367
R1530 B.n804 B.n803 163.367
R1531 B.n804 B.n5 163.367
R1532 B.n6 B.n5 163.367
R1533 B.n7 B.n6 163.367
R1534 B.n809 B.n7 163.367
R1535 B.n809 B.n12 163.367
R1536 B.n13 B.n12 163.367
R1537 B.n14 B.n13 163.367
R1538 B.n814 B.n14 163.367
R1539 B.n814 B.n19 163.367
R1540 B.n20 B.n19 163.367
R1541 B.n21 B.n20 163.367
R1542 B.n819 B.n21 163.367
R1543 B.n819 B.n26 163.367
R1544 B.n27 B.n26 163.367
R1545 B.n28 B.n27 163.367
R1546 B.n824 B.n28 163.367
R1547 B.n824 B.n33 163.367
R1548 B.n34 B.n33 163.367
R1549 B.n35 B.n34 163.367
R1550 B.n829 B.n35 163.367
R1551 B.n829 B.n40 163.367
R1552 B.n41 B.n40 163.367
R1553 B.n42 B.n41 163.367
R1554 B.n834 B.n42 163.367
R1555 B.n834 B.n47 163.367
R1556 B.n48 B.n47 163.367
R1557 B.n49 B.n48 163.367
R1558 B.n839 B.n49 163.367
R1559 B.n839 B.n54 163.367
R1560 B.n55 B.n54 163.367
R1561 B.n56 B.n55 163.367
R1562 B.n844 B.n56 163.367
R1563 B.n844 B.n61 163.367
R1564 B.n62 B.n61 163.367
R1565 B.n63 B.n62 163.367
R1566 B.n849 B.n63 163.367
R1567 B.n849 B.n68 163.367
R1568 B.n69 B.n68 163.367
R1569 B.n70 B.n69 163.367
R1570 B.n854 B.n70 163.367
R1571 B.n854 B.n75 163.367
R1572 B.n76 B.n75 163.367
R1573 B.n77 B.n76 163.367
R1574 B.n859 B.n77 163.367
R1575 B.n859 B.n82 163.367
R1576 B.n83 B.n82 163.367
R1577 B.n84 B.n83 163.367
R1578 B.n864 B.n84 163.367
R1579 B.n864 B.n89 163.367
R1580 B.n90 B.n89 163.367
R1581 B.n91 B.n90 163.367
R1582 B.n869 B.n91 163.367
R1583 B.n869 B.n96 163.367
R1584 B.n97 B.n96 163.367
R1585 B.n98 B.n97 163.367
R1586 B.n145 B.n98 163.367
R1587 B.n151 B.n102 163.367
R1588 B.n155 B.n154 163.367
R1589 B.n159 B.n158 163.367
R1590 B.n163 B.n162 163.367
R1591 B.n167 B.n166 163.367
R1592 B.n171 B.n170 163.367
R1593 B.n175 B.n174 163.367
R1594 B.n179 B.n178 163.367
R1595 B.n183 B.n182 163.367
R1596 B.n187 B.n186 163.367
R1597 B.n191 B.n190 163.367
R1598 B.n195 B.n194 163.367
R1599 B.n199 B.n198 163.367
R1600 B.n203 B.n202 163.367
R1601 B.n207 B.n206 163.367
R1602 B.n211 B.n210 163.367
R1603 B.n215 B.n214 163.367
R1604 B.n219 B.n218 163.367
R1605 B.n223 B.n222 163.367
R1606 B.n227 B.n226 163.367
R1607 B.n231 B.n230 163.367
R1608 B.n235 B.n234 163.367
R1609 B.n239 B.n238 163.367
R1610 B.n244 B.n243 163.367
R1611 B.n248 B.n247 163.367
R1612 B.n252 B.n251 163.367
R1613 B.n256 B.n255 163.367
R1614 B.n260 B.n259 163.367
R1615 B.n264 B.n263 163.367
R1616 B.n268 B.n267 163.367
R1617 B.n272 B.n271 163.367
R1618 B.n276 B.n275 163.367
R1619 B.n280 B.n279 163.367
R1620 B.n284 B.n283 163.367
R1621 B.n288 B.n287 163.367
R1622 B.n292 B.n291 163.367
R1623 B.n296 B.n295 163.367
R1624 B.n300 B.n299 163.367
R1625 B.n304 B.n303 163.367
R1626 B.n308 B.n307 163.367
R1627 B.n312 B.n311 163.367
R1628 B.n876 B.n144 163.367
R1629 B.n638 B.n421 93.0748
R1630 B.n877 B.n99 93.0748
R1631 B.n470 B.n469 77.5763
R1632 B.n468 B.n467 77.5763
R1633 B.n149 B.n148 77.5763
R1634 B.n147 B.n146 77.5763
R1635 B.n640 B.n639 71.676
R1636 B.n466 B.n425 71.676
R1637 B.n632 B.n426 71.676
R1638 B.n628 B.n427 71.676
R1639 B.n624 B.n428 71.676
R1640 B.n620 B.n429 71.676
R1641 B.n616 B.n430 71.676
R1642 B.n612 B.n431 71.676
R1643 B.n608 B.n432 71.676
R1644 B.n604 B.n433 71.676
R1645 B.n600 B.n434 71.676
R1646 B.n596 B.n435 71.676
R1647 B.n592 B.n436 71.676
R1648 B.n588 B.n437 71.676
R1649 B.n584 B.n438 71.676
R1650 B.n580 B.n439 71.676
R1651 B.n576 B.n440 71.676
R1652 B.n572 B.n441 71.676
R1653 B.n568 B.n442 71.676
R1654 B.n563 B.n443 71.676
R1655 B.n559 B.n444 71.676
R1656 B.n555 B.n445 71.676
R1657 B.n551 B.n446 71.676
R1658 B.n547 B.n447 71.676
R1659 B.n543 B.n448 71.676
R1660 B.n539 B.n449 71.676
R1661 B.n535 B.n450 71.676
R1662 B.n531 B.n451 71.676
R1663 B.n527 B.n452 71.676
R1664 B.n523 B.n453 71.676
R1665 B.n519 B.n454 71.676
R1666 B.n515 B.n455 71.676
R1667 B.n511 B.n456 71.676
R1668 B.n507 B.n457 71.676
R1669 B.n503 B.n458 71.676
R1670 B.n499 B.n459 71.676
R1671 B.n495 B.n460 71.676
R1672 B.n491 B.n461 71.676
R1673 B.n487 B.n462 71.676
R1674 B.n483 B.n463 71.676
R1675 B.n479 B.n464 71.676
R1676 B.n475 B.n465 71.676
R1677 B.n879 B.n878 71.676
R1678 B.n151 B.n103 71.676
R1679 B.n155 B.n104 71.676
R1680 B.n159 B.n105 71.676
R1681 B.n163 B.n106 71.676
R1682 B.n167 B.n107 71.676
R1683 B.n171 B.n108 71.676
R1684 B.n175 B.n109 71.676
R1685 B.n179 B.n110 71.676
R1686 B.n183 B.n111 71.676
R1687 B.n187 B.n112 71.676
R1688 B.n191 B.n113 71.676
R1689 B.n195 B.n114 71.676
R1690 B.n199 B.n115 71.676
R1691 B.n203 B.n116 71.676
R1692 B.n207 B.n117 71.676
R1693 B.n211 B.n118 71.676
R1694 B.n215 B.n119 71.676
R1695 B.n219 B.n120 71.676
R1696 B.n223 B.n121 71.676
R1697 B.n227 B.n122 71.676
R1698 B.n231 B.n123 71.676
R1699 B.n235 B.n124 71.676
R1700 B.n239 B.n125 71.676
R1701 B.n244 B.n126 71.676
R1702 B.n248 B.n127 71.676
R1703 B.n252 B.n128 71.676
R1704 B.n256 B.n129 71.676
R1705 B.n260 B.n130 71.676
R1706 B.n264 B.n131 71.676
R1707 B.n268 B.n132 71.676
R1708 B.n272 B.n133 71.676
R1709 B.n276 B.n134 71.676
R1710 B.n280 B.n135 71.676
R1711 B.n284 B.n136 71.676
R1712 B.n288 B.n137 71.676
R1713 B.n292 B.n138 71.676
R1714 B.n296 B.n139 71.676
R1715 B.n300 B.n140 71.676
R1716 B.n304 B.n141 71.676
R1717 B.n308 B.n142 71.676
R1718 B.n312 B.n143 71.676
R1719 B.n144 B.n143 71.676
R1720 B.n311 B.n142 71.676
R1721 B.n307 B.n141 71.676
R1722 B.n303 B.n140 71.676
R1723 B.n299 B.n139 71.676
R1724 B.n295 B.n138 71.676
R1725 B.n291 B.n137 71.676
R1726 B.n287 B.n136 71.676
R1727 B.n283 B.n135 71.676
R1728 B.n279 B.n134 71.676
R1729 B.n275 B.n133 71.676
R1730 B.n271 B.n132 71.676
R1731 B.n267 B.n131 71.676
R1732 B.n263 B.n130 71.676
R1733 B.n259 B.n129 71.676
R1734 B.n255 B.n128 71.676
R1735 B.n251 B.n127 71.676
R1736 B.n247 B.n126 71.676
R1737 B.n243 B.n125 71.676
R1738 B.n238 B.n124 71.676
R1739 B.n234 B.n123 71.676
R1740 B.n230 B.n122 71.676
R1741 B.n226 B.n121 71.676
R1742 B.n222 B.n120 71.676
R1743 B.n218 B.n119 71.676
R1744 B.n214 B.n118 71.676
R1745 B.n210 B.n117 71.676
R1746 B.n206 B.n116 71.676
R1747 B.n202 B.n115 71.676
R1748 B.n198 B.n114 71.676
R1749 B.n194 B.n113 71.676
R1750 B.n190 B.n112 71.676
R1751 B.n186 B.n111 71.676
R1752 B.n182 B.n110 71.676
R1753 B.n178 B.n109 71.676
R1754 B.n174 B.n108 71.676
R1755 B.n170 B.n107 71.676
R1756 B.n166 B.n106 71.676
R1757 B.n162 B.n105 71.676
R1758 B.n158 B.n104 71.676
R1759 B.n154 B.n103 71.676
R1760 B.n878 B.n102 71.676
R1761 B.n639 B.n424 71.676
R1762 B.n633 B.n425 71.676
R1763 B.n629 B.n426 71.676
R1764 B.n625 B.n427 71.676
R1765 B.n621 B.n428 71.676
R1766 B.n617 B.n429 71.676
R1767 B.n613 B.n430 71.676
R1768 B.n609 B.n431 71.676
R1769 B.n605 B.n432 71.676
R1770 B.n601 B.n433 71.676
R1771 B.n597 B.n434 71.676
R1772 B.n593 B.n435 71.676
R1773 B.n589 B.n436 71.676
R1774 B.n585 B.n437 71.676
R1775 B.n581 B.n438 71.676
R1776 B.n577 B.n439 71.676
R1777 B.n573 B.n440 71.676
R1778 B.n569 B.n441 71.676
R1779 B.n564 B.n442 71.676
R1780 B.n560 B.n443 71.676
R1781 B.n556 B.n444 71.676
R1782 B.n552 B.n445 71.676
R1783 B.n548 B.n446 71.676
R1784 B.n544 B.n447 71.676
R1785 B.n540 B.n448 71.676
R1786 B.n536 B.n449 71.676
R1787 B.n532 B.n450 71.676
R1788 B.n528 B.n451 71.676
R1789 B.n524 B.n452 71.676
R1790 B.n520 B.n453 71.676
R1791 B.n516 B.n454 71.676
R1792 B.n512 B.n455 71.676
R1793 B.n508 B.n456 71.676
R1794 B.n504 B.n457 71.676
R1795 B.n500 B.n458 71.676
R1796 B.n496 B.n459 71.676
R1797 B.n492 B.n460 71.676
R1798 B.n488 B.n461 71.676
R1799 B.n484 B.n462 71.676
R1800 B.n480 B.n463 71.676
R1801 B.n476 B.n464 71.676
R1802 B.n472 B.n465 71.676
R1803 B.n471 B.n470 59.5399
R1804 B.n566 B.n468 59.5399
R1805 B.n150 B.n149 59.5399
R1806 B.n241 B.n147 59.5399
R1807 B.n645 B.n421 46.8824
R1808 B.n645 B.n417 46.8824
R1809 B.n651 B.n417 46.8824
R1810 B.n651 B.n413 46.8824
R1811 B.n657 B.n413 46.8824
R1812 B.n657 B.n409 46.8824
R1813 B.n663 B.n409 46.8824
R1814 B.n663 B.n405 46.8824
R1815 B.n669 B.n405 46.8824
R1816 B.n675 B.n401 46.8824
R1817 B.n675 B.n397 46.8824
R1818 B.n681 B.n397 46.8824
R1819 B.n681 B.n393 46.8824
R1820 B.n687 B.n393 46.8824
R1821 B.n687 B.n389 46.8824
R1822 B.n693 B.n389 46.8824
R1823 B.n693 B.n385 46.8824
R1824 B.n699 B.n385 46.8824
R1825 B.n699 B.n381 46.8824
R1826 B.n705 B.n381 46.8824
R1827 B.n705 B.n377 46.8824
R1828 B.n711 B.n377 46.8824
R1829 B.n717 B.n373 46.8824
R1830 B.n717 B.n369 46.8824
R1831 B.n723 B.n369 46.8824
R1832 B.n723 B.n365 46.8824
R1833 B.n729 B.n365 46.8824
R1834 B.n729 B.n361 46.8824
R1835 B.n735 B.n361 46.8824
R1836 B.n735 B.n357 46.8824
R1837 B.n741 B.n357 46.8824
R1838 B.n741 B.n353 46.8824
R1839 B.n747 B.n353 46.8824
R1840 B.n753 B.n349 46.8824
R1841 B.n753 B.n345 46.8824
R1842 B.n759 B.n345 46.8824
R1843 B.n759 B.n341 46.8824
R1844 B.n765 B.n341 46.8824
R1845 B.n765 B.n337 46.8824
R1846 B.n771 B.n337 46.8824
R1847 B.n771 B.n333 46.8824
R1848 B.n777 B.n333 46.8824
R1849 B.n777 B.n329 46.8824
R1850 B.n783 B.n329 46.8824
R1851 B.n789 B.n325 46.8824
R1852 B.n789 B.n321 46.8824
R1853 B.n796 B.n321 46.8824
R1854 B.n796 B.n317 46.8824
R1855 B.n802 B.n317 46.8824
R1856 B.n802 B.n4 46.8824
R1857 B.n990 B.n4 46.8824
R1858 B.n990 B.n989 46.8824
R1859 B.n989 B.n988 46.8824
R1860 B.n988 B.n8 46.8824
R1861 B.n982 B.n8 46.8824
R1862 B.n982 B.n981 46.8824
R1863 B.n981 B.n980 46.8824
R1864 B.n980 B.n15 46.8824
R1865 B.n974 B.n973 46.8824
R1866 B.n973 B.n972 46.8824
R1867 B.n972 B.n22 46.8824
R1868 B.n966 B.n22 46.8824
R1869 B.n966 B.n965 46.8824
R1870 B.n965 B.n964 46.8824
R1871 B.n964 B.n29 46.8824
R1872 B.n958 B.n29 46.8824
R1873 B.n958 B.n957 46.8824
R1874 B.n957 B.n956 46.8824
R1875 B.n956 B.n36 46.8824
R1876 B.n950 B.n949 46.8824
R1877 B.n949 B.n948 46.8824
R1878 B.n948 B.n43 46.8824
R1879 B.n942 B.n43 46.8824
R1880 B.n942 B.n941 46.8824
R1881 B.n941 B.n940 46.8824
R1882 B.n940 B.n50 46.8824
R1883 B.n934 B.n50 46.8824
R1884 B.n934 B.n933 46.8824
R1885 B.n933 B.n932 46.8824
R1886 B.n932 B.n57 46.8824
R1887 B.n926 B.n925 46.8824
R1888 B.n925 B.n924 46.8824
R1889 B.n924 B.n64 46.8824
R1890 B.n918 B.n64 46.8824
R1891 B.n918 B.n917 46.8824
R1892 B.n917 B.n916 46.8824
R1893 B.n916 B.n71 46.8824
R1894 B.n910 B.n71 46.8824
R1895 B.n910 B.n909 46.8824
R1896 B.n909 B.n908 46.8824
R1897 B.n908 B.n78 46.8824
R1898 B.n902 B.n78 46.8824
R1899 B.n902 B.n901 46.8824
R1900 B.n900 B.n85 46.8824
R1901 B.n894 B.n85 46.8824
R1902 B.n894 B.n893 46.8824
R1903 B.n893 B.n892 46.8824
R1904 B.n892 B.n92 46.8824
R1905 B.n886 B.n92 46.8824
R1906 B.n886 B.n885 46.8824
R1907 B.n885 B.n884 46.8824
R1908 B.n884 B.n99 46.8824
R1909 B.t6 B.n401 46.1929
R1910 B.n711 B.t19 46.1929
R1911 B.n926 B.t3 46.1929
R1912 B.n901 B.t13 46.1929
R1913 B.n747 B.t0 35.1619
R1914 B.n950 B.t4 35.1619
R1915 B.n881 B.n880 34.4981
R1916 B.n875 B.n874 34.4981
R1917 B.n473 B.n419 34.4981
R1918 B.n642 B.n641 34.4981
R1919 B.n783 B.t1 24.1309
R1920 B.n974 B.t2 24.1309
R1921 B.t1 B.n325 22.752
R1922 B.t2 B.n15 22.752
R1923 B B.n992 18.0485
R1924 B.t0 B.n349 11.721
R1925 B.t4 B.n36 11.721
R1926 B.n880 B.n101 10.6151
R1927 B.n152 B.n101 10.6151
R1928 B.n153 B.n152 10.6151
R1929 B.n156 B.n153 10.6151
R1930 B.n157 B.n156 10.6151
R1931 B.n160 B.n157 10.6151
R1932 B.n161 B.n160 10.6151
R1933 B.n164 B.n161 10.6151
R1934 B.n165 B.n164 10.6151
R1935 B.n168 B.n165 10.6151
R1936 B.n169 B.n168 10.6151
R1937 B.n172 B.n169 10.6151
R1938 B.n173 B.n172 10.6151
R1939 B.n176 B.n173 10.6151
R1940 B.n177 B.n176 10.6151
R1941 B.n180 B.n177 10.6151
R1942 B.n181 B.n180 10.6151
R1943 B.n184 B.n181 10.6151
R1944 B.n185 B.n184 10.6151
R1945 B.n188 B.n185 10.6151
R1946 B.n189 B.n188 10.6151
R1947 B.n192 B.n189 10.6151
R1948 B.n193 B.n192 10.6151
R1949 B.n196 B.n193 10.6151
R1950 B.n197 B.n196 10.6151
R1951 B.n200 B.n197 10.6151
R1952 B.n201 B.n200 10.6151
R1953 B.n204 B.n201 10.6151
R1954 B.n205 B.n204 10.6151
R1955 B.n208 B.n205 10.6151
R1956 B.n209 B.n208 10.6151
R1957 B.n212 B.n209 10.6151
R1958 B.n213 B.n212 10.6151
R1959 B.n216 B.n213 10.6151
R1960 B.n217 B.n216 10.6151
R1961 B.n220 B.n217 10.6151
R1962 B.n221 B.n220 10.6151
R1963 B.n225 B.n224 10.6151
R1964 B.n228 B.n225 10.6151
R1965 B.n229 B.n228 10.6151
R1966 B.n232 B.n229 10.6151
R1967 B.n233 B.n232 10.6151
R1968 B.n236 B.n233 10.6151
R1969 B.n237 B.n236 10.6151
R1970 B.n240 B.n237 10.6151
R1971 B.n245 B.n242 10.6151
R1972 B.n246 B.n245 10.6151
R1973 B.n249 B.n246 10.6151
R1974 B.n250 B.n249 10.6151
R1975 B.n253 B.n250 10.6151
R1976 B.n254 B.n253 10.6151
R1977 B.n257 B.n254 10.6151
R1978 B.n258 B.n257 10.6151
R1979 B.n261 B.n258 10.6151
R1980 B.n262 B.n261 10.6151
R1981 B.n265 B.n262 10.6151
R1982 B.n266 B.n265 10.6151
R1983 B.n269 B.n266 10.6151
R1984 B.n270 B.n269 10.6151
R1985 B.n273 B.n270 10.6151
R1986 B.n274 B.n273 10.6151
R1987 B.n277 B.n274 10.6151
R1988 B.n278 B.n277 10.6151
R1989 B.n281 B.n278 10.6151
R1990 B.n282 B.n281 10.6151
R1991 B.n285 B.n282 10.6151
R1992 B.n286 B.n285 10.6151
R1993 B.n289 B.n286 10.6151
R1994 B.n290 B.n289 10.6151
R1995 B.n293 B.n290 10.6151
R1996 B.n294 B.n293 10.6151
R1997 B.n297 B.n294 10.6151
R1998 B.n298 B.n297 10.6151
R1999 B.n301 B.n298 10.6151
R2000 B.n302 B.n301 10.6151
R2001 B.n305 B.n302 10.6151
R2002 B.n306 B.n305 10.6151
R2003 B.n309 B.n306 10.6151
R2004 B.n310 B.n309 10.6151
R2005 B.n313 B.n310 10.6151
R2006 B.n314 B.n313 10.6151
R2007 B.n875 B.n314 10.6151
R2008 B.n647 B.n419 10.6151
R2009 B.n648 B.n647 10.6151
R2010 B.n649 B.n648 10.6151
R2011 B.n649 B.n411 10.6151
R2012 B.n659 B.n411 10.6151
R2013 B.n660 B.n659 10.6151
R2014 B.n661 B.n660 10.6151
R2015 B.n661 B.n403 10.6151
R2016 B.n671 B.n403 10.6151
R2017 B.n672 B.n671 10.6151
R2018 B.n673 B.n672 10.6151
R2019 B.n673 B.n395 10.6151
R2020 B.n683 B.n395 10.6151
R2021 B.n684 B.n683 10.6151
R2022 B.n685 B.n684 10.6151
R2023 B.n685 B.n387 10.6151
R2024 B.n695 B.n387 10.6151
R2025 B.n696 B.n695 10.6151
R2026 B.n697 B.n696 10.6151
R2027 B.n697 B.n379 10.6151
R2028 B.n707 B.n379 10.6151
R2029 B.n708 B.n707 10.6151
R2030 B.n709 B.n708 10.6151
R2031 B.n709 B.n371 10.6151
R2032 B.n719 B.n371 10.6151
R2033 B.n720 B.n719 10.6151
R2034 B.n721 B.n720 10.6151
R2035 B.n721 B.n363 10.6151
R2036 B.n731 B.n363 10.6151
R2037 B.n732 B.n731 10.6151
R2038 B.n733 B.n732 10.6151
R2039 B.n733 B.n355 10.6151
R2040 B.n743 B.n355 10.6151
R2041 B.n744 B.n743 10.6151
R2042 B.n745 B.n744 10.6151
R2043 B.n745 B.n347 10.6151
R2044 B.n755 B.n347 10.6151
R2045 B.n756 B.n755 10.6151
R2046 B.n757 B.n756 10.6151
R2047 B.n757 B.n339 10.6151
R2048 B.n767 B.n339 10.6151
R2049 B.n768 B.n767 10.6151
R2050 B.n769 B.n768 10.6151
R2051 B.n769 B.n331 10.6151
R2052 B.n779 B.n331 10.6151
R2053 B.n780 B.n779 10.6151
R2054 B.n781 B.n780 10.6151
R2055 B.n781 B.n323 10.6151
R2056 B.n791 B.n323 10.6151
R2057 B.n792 B.n791 10.6151
R2058 B.n794 B.n792 10.6151
R2059 B.n794 B.n793 10.6151
R2060 B.n793 B.n315 10.6151
R2061 B.n805 B.n315 10.6151
R2062 B.n806 B.n805 10.6151
R2063 B.n807 B.n806 10.6151
R2064 B.n808 B.n807 10.6151
R2065 B.n810 B.n808 10.6151
R2066 B.n811 B.n810 10.6151
R2067 B.n812 B.n811 10.6151
R2068 B.n813 B.n812 10.6151
R2069 B.n815 B.n813 10.6151
R2070 B.n816 B.n815 10.6151
R2071 B.n817 B.n816 10.6151
R2072 B.n818 B.n817 10.6151
R2073 B.n820 B.n818 10.6151
R2074 B.n821 B.n820 10.6151
R2075 B.n822 B.n821 10.6151
R2076 B.n823 B.n822 10.6151
R2077 B.n825 B.n823 10.6151
R2078 B.n826 B.n825 10.6151
R2079 B.n827 B.n826 10.6151
R2080 B.n828 B.n827 10.6151
R2081 B.n830 B.n828 10.6151
R2082 B.n831 B.n830 10.6151
R2083 B.n832 B.n831 10.6151
R2084 B.n833 B.n832 10.6151
R2085 B.n835 B.n833 10.6151
R2086 B.n836 B.n835 10.6151
R2087 B.n837 B.n836 10.6151
R2088 B.n838 B.n837 10.6151
R2089 B.n840 B.n838 10.6151
R2090 B.n841 B.n840 10.6151
R2091 B.n842 B.n841 10.6151
R2092 B.n843 B.n842 10.6151
R2093 B.n845 B.n843 10.6151
R2094 B.n846 B.n845 10.6151
R2095 B.n847 B.n846 10.6151
R2096 B.n848 B.n847 10.6151
R2097 B.n850 B.n848 10.6151
R2098 B.n851 B.n850 10.6151
R2099 B.n852 B.n851 10.6151
R2100 B.n853 B.n852 10.6151
R2101 B.n855 B.n853 10.6151
R2102 B.n856 B.n855 10.6151
R2103 B.n857 B.n856 10.6151
R2104 B.n858 B.n857 10.6151
R2105 B.n860 B.n858 10.6151
R2106 B.n861 B.n860 10.6151
R2107 B.n862 B.n861 10.6151
R2108 B.n863 B.n862 10.6151
R2109 B.n865 B.n863 10.6151
R2110 B.n866 B.n865 10.6151
R2111 B.n867 B.n866 10.6151
R2112 B.n868 B.n867 10.6151
R2113 B.n870 B.n868 10.6151
R2114 B.n871 B.n870 10.6151
R2115 B.n872 B.n871 10.6151
R2116 B.n873 B.n872 10.6151
R2117 B.n874 B.n873 10.6151
R2118 B.n641 B.n423 10.6151
R2119 B.n636 B.n423 10.6151
R2120 B.n636 B.n635 10.6151
R2121 B.n635 B.n634 10.6151
R2122 B.n634 B.n631 10.6151
R2123 B.n631 B.n630 10.6151
R2124 B.n630 B.n627 10.6151
R2125 B.n627 B.n626 10.6151
R2126 B.n626 B.n623 10.6151
R2127 B.n623 B.n622 10.6151
R2128 B.n622 B.n619 10.6151
R2129 B.n619 B.n618 10.6151
R2130 B.n618 B.n615 10.6151
R2131 B.n615 B.n614 10.6151
R2132 B.n614 B.n611 10.6151
R2133 B.n611 B.n610 10.6151
R2134 B.n610 B.n607 10.6151
R2135 B.n607 B.n606 10.6151
R2136 B.n606 B.n603 10.6151
R2137 B.n603 B.n602 10.6151
R2138 B.n602 B.n599 10.6151
R2139 B.n599 B.n598 10.6151
R2140 B.n598 B.n595 10.6151
R2141 B.n595 B.n594 10.6151
R2142 B.n594 B.n591 10.6151
R2143 B.n591 B.n590 10.6151
R2144 B.n590 B.n587 10.6151
R2145 B.n587 B.n586 10.6151
R2146 B.n586 B.n583 10.6151
R2147 B.n583 B.n582 10.6151
R2148 B.n582 B.n579 10.6151
R2149 B.n579 B.n578 10.6151
R2150 B.n578 B.n575 10.6151
R2151 B.n575 B.n574 10.6151
R2152 B.n574 B.n571 10.6151
R2153 B.n571 B.n570 10.6151
R2154 B.n570 B.n567 10.6151
R2155 B.n565 B.n562 10.6151
R2156 B.n562 B.n561 10.6151
R2157 B.n561 B.n558 10.6151
R2158 B.n558 B.n557 10.6151
R2159 B.n557 B.n554 10.6151
R2160 B.n554 B.n553 10.6151
R2161 B.n553 B.n550 10.6151
R2162 B.n550 B.n549 10.6151
R2163 B.n546 B.n545 10.6151
R2164 B.n545 B.n542 10.6151
R2165 B.n542 B.n541 10.6151
R2166 B.n541 B.n538 10.6151
R2167 B.n538 B.n537 10.6151
R2168 B.n537 B.n534 10.6151
R2169 B.n534 B.n533 10.6151
R2170 B.n533 B.n530 10.6151
R2171 B.n530 B.n529 10.6151
R2172 B.n529 B.n526 10.6151
R2173 B.n526 B.n525 10.6151
R2174 B.n525 B.n522 10.6151
R2175 B.n522 B.n521 10.6151
R2176 B.n521 B.n518 10.6151
R2177 B.n518 B.n517 10.6151
R2178 B.n517 B.n514 10.6151
R2179 B.n514 B.n513 10.6151
R2180 B.n513 B.n510 10.6151
R2181 B.n510 B.n509 10.6151
R2182 B.n509 B.n506 10.6151
R2183 B.n506 B.n505 10.6151
R2184 B.n505 B.n502 10.6151
R2185 B.n502 B.n501 10.6151
R2186 B.n501 B.n498 10.6151
R2187 B.n498 B.n497 10.6151
R2188 B.n497 B.n494 10.6151
R2189 B.n494 B.n493 10.6151
R2190 B.n493 B.n490 10.6151
R2191 B.n490 B.n489 10.6151
R2192 B.n489 B.n486 10.6151
R2193 B.n486 B.n485 10.6151
R2194 B.n485 B.n482 10.6151
R2195 B.n482 B.n481 10.6151
R2196 B.n481 B.n478 10.6151
R2197 B.n478 B.n477 10.6151
R2198 B.n477 B.n474 10.6151
R2199 B.n474 B.n473 10.6151
R2200 B.n643 B.n642 10.6151
R2201 B.n643 B.n415 10.6151
R2202 B.n653 B.n415 10.6151
R2203 B.n654 B.n653 10.6151
R2204 B.n655 B.n654 10.6151
R2205 B.n655 B.n407 10.6151
R2206 B.n665 B.n407 10.6151
R2207 B.n666 B.n665 10.6151
R2208 B.n667 B.n666 10.6151
R2209 B.n667 B.n399 10.6151
R2210 B.n677 B.n399 10.6151
R2211 B.n678 B.n677 10.6151
R2212 B.n679 B.n678 10.6151
R2213 B.n679 B.n391 10.6151
R2214 B.n689 B.n391 10.6151
R2215 B.n690 B.n689 10.6151
R2216 B.n691 B.n690 10.6151
R2217 B.n691 B.n383 10.6151
R2218 B.n701 B.n383 10.6151
R2219 B.n702 B.n701 10.6151
R2220 B.n703 B.n702 10.6151
R2221 B.n703 B.n375 10.6151
R2222 B.n713 B.n375 10.6151
R2223 B.n714 B.n713 10.6151
R2224 B.n715 B.n714 10.6151
R2225 B.n715 B.n367 10.6151
R2226 B.n725 B.n367 10.6151
R2227 B.n726 B.n725 10.6151
R2228 B.n727 B.n726 10.6151
R2229 B.n727 B.n359 10.6151
R2230 B.n737 B.n359 10.6151
R2231 B.n738 B.n737 10.6151
R2232 B.n739 B.n738 10.6151
R2233 B.n739 B.n351 10.6151
R2234 B.n749 B.n351 10.6151
R2235 B.n750 B.n749 10.6151
R2236 B.n751 B.n750 10.6151
R2237 B.n751 B.n343 10.6151
R2238 B.n761 B.n343 10.6151
R2239 B.n762 B.n761 10.6151
R2240 B.n763 B.n762 10.6151
R2241 B.n763 B.n335 10.6151
R2242 B.n773 B.n335 10.6151
R2243 B.n774 B.n773 10.6151
R2244 B.n775 B.n774 10.6151
R2245 B.n775 B.n327 10.6151
R2246 B.n785 B.n327 10.6151
R2247 B.n786 B.n785 10.6151
R2248 B.n787 B.n786 10.6151
R2249 B.n787 B.n319 10.6151
R2250 B.n798 B.n319 10.6151
R2251 B.n799 B.n798 10.6151
R2252 B.n800 B.n799 10.6151
R2253 B.n800 B.n0 10.6151
R2254 B.n986 B.n1 10.6151
R2255 B.n986 B.n985 10.6151
R2256 B.n985 B.n984 10.6151
R2257 B.n984 B.n10 10.6151
R2258 B.n978 B.n10 10.6151
R2259 B.n978 B.n977 10.6151
R2260 B.n977 B.n976 10.6151
R2261 B.n976 B.n17 10.6151
R2262 B.n970 B.n17 10.6151
R2263 B.n970 B.n969 10.6151
R2264 B.n969 B.n968 10.6151
R2265 B.n968 B.n24 10.6151
R2266 B.n962 B.n24 10.6151
R2267 B.n962 B.n961 10.6151
R2268 B.n961 B.n960 10.6151
R2269 B.n960 B.n31 10.6151
R2270 B.n954 B.n31 10.6151
R2271 B.n954 B.n953 10.6151
R2272 B.n953 B.n952 10.6151
R2273 B.n952 B.n38 10.6151
R2274 B.n946 B.n38 10.6151
R2275 B.n946 B.n945 10.6151
R2276 B.n945 B.n944 10.6151
R2277 B.n944 B.n45 10.6151
R2278 B.n938 B.n45 10.6151
R2279 B.n938 B.n937 10.6151
R2280 B.n937 B.n936 10.6151
R2281 B.n936 B.n52 10.6151
R2282 B.n930 B.n52 10.6151
R2283 B.n930 B.n929 10.6151
R2284 B.n929 B.n928 10.6151
R2285 B.n928 B.n59 10.6151
R2286 B.n922 B.n59 10.6151
R2287 B.n922 B.n921 10.6151
R2288 B.n921 B.n920 10.6151
R2289 B.n920 B.n66 10.6151
R2290 B.n914 B.n66 10.6151
R2291 B.n914 B.n913 10.6151
R2292 B.n913 B.n912 10.6151
R2293 B.n912 B.n73 10.6151
R2294 B.n906 B.n73 10.6151
R2295 B.n906 B.n905 10.6151
R2296 B.n905 B.n904 10.6151
R2297 B.n904 B.n80 10.6151
R2298 B.n898 B.n80 10.6151
R2299 B.n898 B.n897 10.6151
R2300 B.n897 B.n896 10.6151
R2301 B.n896 B.n87 10.6151
R2302 B.n890 B.n87 10.6151
R2303 B.n890 B.n889 10.6151
R2304 B.n889 B.n888 10.6151
R2305 B.n888 B.n94 10.6151
R2306 B.n882 B.n94 10.6151
R2307 B.n882 B.n881 10.6151
R2308 B.n224 B.n150 6.5566
R2309 B.n241 B.n240 6.5566
R2310 B.n566 B.n565 6.5566
R2311 B.n549 B.n471 6.5566
R2312 B.n221 B.n150 4.05904
R2313 B.n242 B.n241 4.05904
R2314 B.n567 B.n566 4.05904
R2315 B.n546 B.n471 4.05904
R2316 B.n992 B.n0 2.81026
R2317 B.n992 B.n1 2.81026
R2318 B.n669 B.t6 0.689939
R2319 B.t19 B.n373 0.689939
R2320 B.t3 B.n57 0.689939
R2321 B.t13 B.n900 0.689939
R2322 VP.n14 VP.n11 161.3
R2323 VP.n16 VP.n15 161.3
R2324 VP.n17 VP.n10 161.3
R2325 VP.n19 VP.n18 161.3
R2326 VP.n20 VP.n9 161.3
R2327 VP.n22 VP.n21 161.3
R2328 VP.n23 VP.n8 161.3
R2329 VP.n49 VP.n0 161.3
R2330 VP.n48 VP.n47 161.3
R2331 VP.n46 VP.n1 161.3
R2332 VP.n45 VP.n44 161.3
R2333 VP.n43 VP.n2 161.3
R2334 VP.n42 VP.n41 161.3
R2335 VP.n40 VP.n3 161.3
R2336 VP.n39 VP.n38 161.3
R2337 VP.n37 VP.n4 161.3
R2338 VP.n36 VP.n35 161.3
R2339 VP.n34 VP.n5 161.3
R2340 VP.n33 VP.n32 161.3
R2341 VP.n31 VP.n6 161.3
R2342 VP.n30 VP.n29 161.3
R2343 VP.n28 VP.n7 161.3
R2344 VP.n13 VP.t3 102.317
R2345 VP.n50 VP.t5 70.1335
R2346 VP.n38 VP.t0 70.1335
R2347 VP.n26 VP.t2 70.1335
R2348 VP.n12 VP.t4 70.1335
R2349 VP.n24 VP.t1 70.1335
R2350 VP.n27 VP.n26 57.7881
R2351 VP.n51 VP.n50 57.7881
R2352 VP.n25 VP.n24 57.7881
R2353 VP.n27 VP.n25 52.1029
R2354 VP.n13 VP.n12 50.586
R2355 VP.n32 VP.n31 40.577
R2356 VP.n32 VP.n5 40.577
R2357 VP.n44 VP.n43 40.577
R2358 VP.n44 VP.n1 40.577
R2359 VP.n18 VP.n9 40.577
R2360 VP.n18 VP.n17 40.577
R2361 VP.n26 VP.n7 24.5923
R2362 VP.n30 VP.n7 24.5923
R2363 VP.n31 VP.n30 24.5923
R2364 VP.n36 VP.n5 24.5923
R2365 VP.n37 VP.n36 24.5923
R2366 VP.n38 VP.n37 24.5923
R2367 VP.n38 VP.n3 24.5923
R2368 VP.n42 VP.n3 24.5923
R2369 VP.n43 VP.n42 24.5923
R2370 VP.n48 VP.n1 24.5923
R2371 VP.n49 VP.n48 24.5923
R2372 VP.n50 VP.n49 24.5923
R2373 VP.n22 VP.n9 24.5923
R2374 VP.n23 VP.n22 24.5923
R2375 VP.n24 VP.n23 24.5923
R2376 VP.n12 VP.n11 24.5923
R2377 VP.n16 VP.n11 24.5923
R2378 VP.n17 VP.n16 24.5923
R2379 VP.n14 VP.n13 2.51554
R2380 VP.n25 VP.n8 0.417304
R2381 VP.n28 VP.n27 0.417304
R2382 VP.n51 VP.n0 0.417304
R2383 VP VP.n51 0.394524
R2384 VP.n15 VP.n14 0.189894
R2385 VP.n15 VP.n10 0.189894
R2386 VP.n19 VP.n10 0.189894
R2387 VP.n20 VP.n19 0.189894
R2388 VP.n21 VP.n20 0.189894
R2389 VP.n21 VP.n8 0.189894
R2390 VP.n29 VP.n28 0.189894
R2391 VP.n29 VP.n6 0.189894
R2392 VP.n33 VP.n6 0.189894
R2393 VP.n34 VP.n33 0.189894
R2394 VP.n35 VP.n34 0.189894
R2395 VP.n35 VP.n4 0.189894
R2396 VP.n39 VP.n4 0.189894
R2397 VP.n40 VP.n39 0.189894
R2398 VP.n41 VP.n40 0.189894
R2399 VP.n41 VP.n2 0.189894
R2400 VP.n45 VP.n2 0.189894
R2401 VP.n46 VP.n45 0.189894
R2402 VP.n47 VP.n46 0.189894
R2403 VP.n47 VP.n0 0.189894
R2404 VDD1.n52 VDD1.n0 289.615
R2405 VDD1.n109 VDD1.n57 289.615
R2406 VDD1.n53 VDD1.n52 185
R2407 VDD1.n51 VDD1.n50 185
R2408 VDD1.n4 VDD1.n3 185
R2409 VDD1.n45 VDD1.n44 185
R2410 VDD1.n43 VDD1.n42 185
R2411 VDD1.n41 VDD1.n7 185
R2412 VDD1.n11 VDD1.n8 185
R2413 VDD1.n36 VDD1.n35 185
R2414 VDD1.n34 VDD1.n33 185
R2415 VDD1.n13 VDD1.n12 185
R2416 VDD1.n28 VDD1.n27 185
R2417 VDD1.n26 VDD1.n25 185
R2418 VDD1.n17 VDD1.n16 185
R2419 VDD1.n20 VDD1.n19 185
R2420 VDD1.n76 VDD1.n75 185
R2421 VDD1.n73 VDD1.n72 185
R2422 VDD1.n82 VDD1.n81 185
R2423 VDD1.n84 VDD1.n83 185
R2424 VDD1.n69 VDD1.n68 185
R2425 VDD1.n90 VDD1.n89 185
R2426 VDD1.n93 VDD1.n92 185
R2427 VDD1.n91 VDD1.n65 185
R2428 VDD1.n98 VDD1.n64 185
R2429 VDD1.n100 VDD1.n99 185
R2430 VDD1.n102 VDD1.n101 185
R2431 VDD1.n61 VDD1.n60 185
R2432 VDD1.n108 VDD1.n107 185
R2433 VDD1.n110 VDD1.n109 185
R2434 VDD1.t2 VDD1.n18 149.524
R2435 VDD1.t3 VDD1.n74 149.524
R2436 VDD1.n52 VDD1.n51 104.615
R2437 VDD1.n51 VDD1.n3 104.615
R2438 VDD1.n44 VDD1.n3 104.615
R2439 VDD1.n44 VDD1.n43 104.615
R2440 VDD1.n43 VDD1.n7 104.615
R2441 VDD1.n11 VDD1.n7 104.615
R2442 VDD1.n35 VDD1.n11 104.615
R2443 VDD1.n35 VDD1.n34 104.615
R2444 VDD1.n34 VDD1.n12 104.615
R2445 VDD1.n27 VDD1.n12 104.615
R2446 VDD1.n27 VDD1.n26 104.615
R2447 VDD1.n26 VDD1.n16 104.615
R2448 VDD1.n19 VDD1.n16 104.615
R2449 VDD1.n75 VDD1.n72 104.615
R2450 VDD1.n82 VDD1.n72 104.615
R2451 VDD1.n83 VDD1.n82 104.615
R2452 VDD1.n83 VDD1.n68 104.615
R2453 VDD1.n90 VDD1.n68 104.615
R2454 VDD1.n92 VDD1.n90 104.615
R2455 VDD1.n92 VDD1.n91 104.615
R2456 VDD1.n91 VDD1.n64 104.615
R2457 VDD1.n100 VDD1.n64 104.615
R2458 VDD1.n101 VDD1.n100 104.615
R2459 VDD1.n101 VDD1.n60 104.615
R2460 VDD1.n108 VDD1.n60 104.615
R2461 VDD1.n109 VDD1.n108 104.615
R2462 VDD1.n115 VDD1.n114 63.1468
R2463 VDD1.n117 VDD1.n116 62.3401
R2464 VDD1.n19 VDD1.t2 52.3082
R2465 VDD1.n75 VDD1.t3 52.3082
R2466 VDD1 VDD1.n56 51.5085
R2467 VDD1.n115 VDD1.n113 51.395
R2468 VDD1.n117 VDD1.n115 46.4362
R2469 VDD1.n42 VDD1.n41 13.1884
R2470 VDD1.n99 VDD1.n98 13.1884
R2471 VDD1.n45 VDD1.n6 12.8005
R2472 VDD1.n40 VDD1.n8 12.8005
R2473 VDD1.n97 VDD1.n65 12.8005
R2474 VDD1.n102 VDD1.n63 12.8005
R2475 VDD1.n46 VDD1.n4 12.0247
R2476 VDD1.n37 VDD1.n36 12.0247
R2477 VDD1.n94 VDD1.n93 12.0247
R2478 VDD1.n103 VDD1.n61 12.0247
R2479 VDD1.n50 VDD1.n49 11.249
R2480 VDD1.n33 VDD1.n10 11.249
R2481 VDD1.n89 VDD1.n67 11.249
R2482 VDD1.n107 VDD1.n106 11.249
R2483 VDD1.n53 VDD1.n2 10.4732
R2484 VDD1.n32 VDD1.n13 10.4732
R2485 VDD1.n88 VDD1.n69 10.4732
R2486 VDD1.n110 VDD1.n59 10.4732
R2487 VDD1.n20 VDD1.n18 10.2747
R2488 VDD1.n76 VDD1.n74 10.2747
R2489 VDD1.n54 VDD1.n0 9.69747
R2490 VDD1.n29 VDD1.n28 9.69747
R2491 VDD1.n85 VDD1.n84 9.69747
R2492 VDD1.n111 VDD1.n57 9.69747
R2493 VDD1.n56 VDD1.n55 9.45567
R2494 VDD1.n113 VDD1.n112 9.45567
R2495 VDD1.n22 VDD1.n21 9.3005
R2496 VDD1.n24 VDD1.n23 9.3005
R2497 VDD1.n15 VDD1.n14 9.3005
R2498 VDD1.n30 VDD1.n29 9.3005
R2499 VDD1.n32 VDD1.n31 9.3005
R2500 VDD1.n10 VDD1.n9 9.3005
R2501 VDD1.n38 VDD1.n37 9.3005
R2502 VDD1.n40 VDD1.n39 9.3005
R2503 VDD1.n55 VDD1.n54 9.3005
R2504 VDD1.n2 VDD1.n1 9.3005
R2505 VDD1.n49 VDD1.n48 9.3005
R2506 VDD1.n47 VDD1.n46 9.3005
R2507 VDD1.n6 VDD1.n5 9.3005
R2508 VDD1.n112 VDD1.n111 9.3005
R2509 VDD1.n59 VDD1.n58 9.3005
R2510 VDD1.n106 VDD1.n105 9.3005
R2511 VDD1.n104 VDD1.n103 9.3005
R2512 VDD1.n63 VDD1.n62 9.3005
R2513 VDD1.n78 VDD1.n77 9.3005
R2514 VDD1.n80 VDD1.n79 9.3005
R2515 VDD1.n71 VDD1.n70 9.3005
R2516 VDD1.n86 VDD1.n85 9.3005
R2517 VDD1.n88 VDD1.n87 9.3005
R2518 VDD1.n67 VDD1.n66 9.3005
R2519 VDD1.n95 VDD1.n94 9.3005
R2520 VDD1.n97 VDD1.n96 9.3005
R2521 VDD1.n25 VDD1.n15 8.92171
R2522 VDD1.n81 VDD1.n71 8.92171
R2523 VDD1.n24 VDD1.n17 8.14595
R2524 VDD1.n80 VDD1.n73 8.14595
R2525 VDD1.n21 VDD1.n20 7.3702
R2526 VDD1.n77 VDD1.n76 7.3702
R2527 VDD1.n21 VDD1.n17 5.81868
R2528 VDD1.n77 VDD1.n73 5.81868
R2529 VDD1.n25 VDD1.n24 5.04292
R2530 VDD1.n81 VDD1.n80 5.04292
R2531 VDD1.n56 VDD1.n0 4.26717
R2532 VDD1.n28 VDD1.n15 4.26717
R2533 VDD1.n84 VDD1.n71 4.26717
R2534 VDD1.n113 VDD1.n57 4.26717
R2535 VDD1.n54 VDD1.n53 3.49141
R2536 VDD1.n29 VDD1.n13 3.49141
R2537 VDD1.n85 VDD1.n69 3.49141
R2538 VDD1.n111 VDD1.n110 3.49141
R2539 VDD1.n22 VDD1.n18 2.84303
R2540 VDD1.n78 VDD1.n74 2.84303
R2541 VDD1.n50 VDD1.n2 2.71565
R2542 VDD1.n33 VDD1.n32 2.71565
R2543 VDD1.n89 VDD1.n88 2.71565
R2544 VDD1.n107 VDD1.n59 2.71565
R2545 VDD1.n49 VDD1.n4 1.93989
R2546 VDD1.n36 VDD1.n10 1.93989
R2547 VDD1.n93 VDD1.n67 1.93989
R2548 VDD1.n106 VDD1.n61 1.93989
R2549 VDD1.n116 VDD1.t1 1.85443
R2550 VDD1.n116 VDD1.t4 1.85443
R2551 VDD1.n114 VDD1.t5 1.85443
R2552 VDD1.n114 VDD1.t0 1.85443
R2553 VDD1.n46 VDD1.n45 1.16414
R2554 VDD1.n37 VDD1.n8 1.16414
R2555 VDD1.n94 VDD1.n65 1.16414
R2556 VDD1.n103 VDD1.n102 1.16414
R2557 VDD1 VDD1.n117 0.804379
R2558 VDD1.n42 VDD1.n6 0.388379
R2559 VDD1.n41 VDD1.n40 0.388379
R2560 VDD1.n98 VDD1.n97 0.388379
R2561 VDD1.n99 VDD1.n63 0.388379
R2562 VDD1.n55 VDD1.n1 0.155672
R2563 VDD1.n48 VDD1.n1 0.155672
R2564 VDD1.n48 VDD1.n47 0.155672
R2565 VDD1.n47 VDD1.n5 0.155672
R2566 VDD1.n39 VDD1.n5 0.155672
R2567 VDD1.n39 VDD1.n38 0.155672
R2568 VDD1.n38 VDD1.n9 0.155672
R2569 VDD1.n31 VDD1.n9 0.155672
R2570 VDD1.n31 VDD1.n30 0.155672
R2571 VDD1.n30 VDD1.n14 0.155672
R2572 VDD1.n23 VDD1.n14 0.155672
R2573 VDD1.n23 VDD1.n22 0.155672
R2574 VDD1.n79 VDD1.n78 0.155672
R2575 VDD1.n79 VDD1.n70 0.155672
R2576 VDD1.n86 VDD1.n70 0.155672
R2577 VDD1.n87 VDD1.n86 0.155672
R2578 VDD1.n87 VDD1.n66 0.155672
R2579 VDD1.n95 VDD1.n66 0.155672
R2580 VDD1.n96 VDD1.n95 0.155672
R2581 VDD1.n96 VDD1.n62 0.155672
R2582 VDD1.n104 VDD1.n62 0.155672
R2583 VDD1.n105 VDD1.n104 0.155672
R2584 VDD1.n105 VDD1.n58 0.155672
R2585 VDD1.n112 VDD1.n58 0.155672
C0 VDD2 VP 0.54891f
C1 VDD2 VTAIL 7.73394f
C2 VDD2 VN 6.37967f
C3 VDD2 VDD1 1.82296f
C4 VP VTAIL 6.87376f
C5 VP VN 7.72088f
C6 VN VTAIL 6.85934f
C7 VP VDD1 6.77357f
C8 VTAIL VDD1 7.67484f
C9 VN VDD1 0.152332f
C10 VDD2 B 6.561971f
C11 VDD1 B 6.744185f
C12 VTAIL B 7.950747f
C13 VN B 15.96767f
C14 VP B 14.688359f
C15 VDD1.n0 B 0.029605f
C16 VDD1.n1 B 0.021904f
C17 VDD1.n2 B 0.01177f
C18 VDD1.n3 B 0.02782f
C19 VDD1.n4 B 0.012462f
C20 VDD1.n5 B 0.021904f
C21 VDD1.n6 B 0.01177f
C22 VDD1.n7 B 0.02782f
C23 VDD1.n8 B 0.012462f
C24 VDD1.n9 B 0.021904f
C25 VDD1.n10 B 0.01177f
C26 VDD1.n11 B 0.02782f
C27 VDD1.n12 B 0.02782f
C28 VDD1.n13 B 0.012462f
C29 VDD1.n14 B 0.021904f
C30 VDD1.n15 B 0.01177f
C31 VDD1.n16 B 0.02782f
C32 VDD1.n17 B 0.012462f
C33 VDD1.n18 B 0.146825f
C34 VDD1.t2 B 0.046832f
C35 VDD1.n19 B 0.020865f
C36 VDD1.n20 B 0.019667f
C37 VDD1.n21 B 0.01177f
C38 VDD1.n22 B 0.976407f
C39 VDD1.n23 B 0.021904f
C40 VDD1.n24 B 0.01177f
C41 VDD1.n25 B 0.012462f
C42 VDD1.n26 B 0.02782f
C43 VDD1.n27 B 0.02782f
C44 VDD1.n28 B 0.012462f
C45 VDD1.n29 B 0.01177f
C46 VDD1.n30 B 0.021904f
C47 VDD1.n31 B 0.021904f
C48 VDD1.n32 B 0.01177f
C49 VDD1.n33 B 0.012462f
C50 VDD1.n34 B 0.02782f
C51 VDD1.n35 B 0.02782f
C52 VDD1.n36 B 0.012462f
C53 VDD1.n37 B 0.01177f
C54 VDD1.n38 B 0.021904f
C55 VDD1.n39 B 0.021904f
C56 VDD1.n40 B 0.01177f
C57 VDD1.n41 B 0.012116f
C58 VDD1.n42 B 0.012116f
C59 VDD1.n43 B 0.02782f
C60 VDD1.n44 B 0.02782f
C61 VDD1.n45 B 0.012462f
C62 VDD1.n46 B 0.01177f
C63 VDD1.n47 B 0.021904f
C64 VDD1.n48 B 0.021904f
C65 VDD1.n49 B 0.01177f
C66 VDD1.n50 B 0.012462f
C67 VDD1.n51 B 0.02782f
C68 VDD1.n52 B 0.058136f
C69 VDD1.n53 B 0.012462f
C70 VDD1.n54 B 0.01177f
C71 VDD1.n55 B 0.05063f
C72 VDD1.n56 B 0.059186f
C73 VDD1.n57 B 0.029605f
C74 VDD1.n58 B 0.021904f
C75 VDD1.n59 B 0.01177f
C76 VDD1.n60 B 0.02782f
C77 VDD1.n61 B 0.012462f
C78 VDD1.n62 B 0.021904f
C79 VDD1.n63 B 0.01177f
C80 VDD1.n64 B 0.02782f
C81 VDD1.n65 B 0.012462f
C82 VDD1.n66 B 0.021904f
C83 VDD1.n67 B 0.01177f
C84 VDD1.n68 B 0.02782f
C85 VDD1.n69 B 0.012462f
C86 VDD1.n70 B 0.021904f
C87 VDD1.n71 B 0.01177f
C88 VDD1.n72 B 0.02782f
C89 VDD1.n73 B 0.012462f
C90 VDD1.n74 B 0.146825f
C91 VDD1.t3 B 0.046832f
C92 VDD1.n75 B 0.020865f
C93 VDD1.n76 B 0.019667f
C94 VDD1.n77 B 0.01177f
C95 VDD1.n78 B 0.976407f
C96 VDD1.n79 B 0.021904f
C97 VDD1.n80 B 0.01177f
C98 VDD1.n81 B 0.012462f
C99 VDD1.n82 B 0.02782f
C100 VDD1.n83 B 0.02782f
C101 VDD1.n84 B 0.012462f
C102 VDD1.n85 B 0.01177f
C103 VDD1.n86 B 0.021904f
C104 VDD1.n87 B 0.021904f
C105 VDD1.n88 B 0.01177f
C106 VDD1.n89 B 0.012462f
C107 VDD1.n90 B 0.02782f
C108 VDD1.n91 B 0.02782f
C109 VDD1.n92 B 0.02782f
C110 VDD1.n93 B 0.012462f
C111 VDD1.n94 B 0.01177f
C112 VDD1.n95 B 0.021904f
C113 VDD1.n96 B 0.021904f
C114 VDD1.n97 B 0.01177f
C115 VDD1.n98 B 0.012116f
C116 VDD1.n99 B 0.012116f
C117 VDD1.n100 B 0.02782f
C118 VDD1.n101 B 0.02782f
C119 VDD1.n102 B 0.012462f
C120 VDD1.n103 B 0.01177f
C121 VDD1.n104 B 0.021904f
C122 VDD1.n105 B 0.021904f
C123 VDD1.n106 B 0.01177f
C124 VDD1.n107 B 0.012462f
C125 VDD1.n108 B 0.02782f
C126 VDD1.n109 B 0.058136f
C127 VDD1.n110 B 0.012462f
C128 VDD1.n111 B 0.01177f
C129 VDD1.n112 B 0.05063f
C130 VDD1.n113 B 0.058321f
C131 VDD1.t5 B 0.184861f
C132 VDD1.t0 B 0.184861f
C133 VDD1.n114 B 1.64127f
C134 VDD1.n115 B 2.81071f
C135 VDD1.t1 B 0.184861f
C136 VDD1.t4 B 0.184861f
C137 VDD1.n116 B 1.63502f
C138 VDD1.n117 B 2.61943f
C139 VP.n0 B 0.03659f
C140 VP.t5 B 2.07065f
C141 VP.n1 B 0.038469f
C142 VP.n2 B 0.019458f
C143 VP.n3 B 0.036083f
C144 VP.n4 B 0.019458f
C145 VP.t0 B 2.07065f
C146 VP.n5 B 0.038469f
C147 VP.n6 B 0.019458f
C148 VP.n7 B 0.036083f
C149 VP.n8 B 0.03659f
C150 VP.t1 B 2.07065f
C151 VP.n9 B 0.038469f
C152 VP.n10 B 0.019458f
C153 VP.n11 B 0.036083f
C154 VP.t3 B 2.3479f
C155 VP.t4 B 2.07065f
C156 VP.n12 B 0.809176f
C157 VP.n13 B 0.769215f
C158 VP.n14 B 0.247713f
C159 VP.n15 B 0.019458f
C160 VP.n16 B 0.036083f
C161 VP.n17 B 0.038469f
C162 VP.n18 B 0.015716f
C163 VP.n19 B 0.019458f
C164 VP.n20 B 0.019458f
C165 VP.n21 B 0.019458f
C166 VP.n22 B 0.036083f
C167 VP.n23 B 0.036083f
C168 VP.n24 B 0.815918f
C169 VP.n25 B 1.19118f
C170 VP.t2 B 2.07065f
C171 VP.n26 B 0.815918f
C172 VP.n27 B 1.20465f
C173 VP.n28 B 0.03659f
C174 VP.n29 B 0.019458f
C175 VP.n30 B 0.036083f
C176 VP.n31 B 0.038469f
C177 VP.n32 B 0.015716f
C178 VP.n33 B 0.019458f
C179 VP.n34 B 0.019458f
C180 VP.n35 B 0.019458f
C181 VP.n36 B 0.036083f
C182 VP.n37 B 0.036083f
C183 VP.n38 B 0.748535f
C184 VP.n39 B 0.019458f
C185 VP.n40 B 0.019458f
C186 VP.n41 B 0.019458f
C187 VP.n42 B 0.036083f
C188 VP.n43 B 0.038469f
C189 VP.n44 B 0.015716f
C190 VP.n45 B 0.019458f
C191 VP.n46 B 0.019458f
C192 VP.n47 B 0.019458f
C193 VP.n48 B 0.036083f
C194 VP.n49 B 0.036083f
C195 VP.n50 B 0.815918f
C196 VP.n51 B 0.054704f
C197 VDD2.n0 B 0.02895f
C198 VDD2.n1 B 0.021419f
C199 VDD2.n2 B 0.01151f
C200 VDD2.n3 B 0.027205f
C201 VDD2.n4 B 0.012187f
C202 VDD2.n5 B 0.021419f
C203 VDD2.n6 B 0.01151f
C204 VDD2.n7 B 0.027205f
C205 VDD2.n8 B 0.012187f
C206 VDD2.n9 B 0.021419f
C207 VDD2.n10 B 0.01151f
C208 VDD2.n11 B 0.027205f
C209 VDD2.n12 B 0.012187f
C210 VDD2.n13 B 0.021419f
C211 VDD2.n14 B 0.01151f
C212 VDD2.n15 B 0.027205f
C213 VDD2.n16 B 0.012187f
C214 VDD2.n17 B 0.143576f
C215 VDD2.t2 B 0.045795f
C216 VDD2.n18 B 0.020404f
C217 VDD2.n19 B 0.019232f
C218 VDD2.n20 B 0.01151f
C219 VDD2.n21 B 0.954799f
C220 VDD2.n22 B 0.021419f
C221 VDD2.n23 B 0.01151f
C222 VDD2.n24 B 0.012187f
C223 VDD2.n25 B 0.027205f
C224 VDD2.n26 B 0.027205f
C225 VDD2.n27 B 0.012187f
C226 VDD2.n28 B 0.01151f
C227 VDD2.n29 B 0.021419f
C228 VDD2.n30 B 0.021419f
C229 VDD2.n31 B 0.01151f
C230 VDD2.n32 B 0.012187f
C231 VDD2.n33 B 0.027205f
C232 VDD2.n34 B 0.027205f
C233 VDD2.n35 B 0.027205f
C234 VDD2.n36 B 0.012187f
C235 VDD2.n37 B 0.01151f
C236 VDD2.n38 B 0.021419f
C237 VDD2.n39 B 0.021419f
C238 VDD2.n40 B 0.01151f
C239 VDD2.n41 B 0.011848f
C240 VDD2.n42 B 0.011848f
C241 VDD2.n43 B 0.027205f
C242 VDD2.n44 B 0.027205f
C243 VDD2.n45 B 0.012187f
C244 VDD2.n46 B 0.01151f
C245 VDD2.n47 B 0.021419f
C246 VDD2.n48 B 0.021419f
C247 VDD2.n49 B 0.01151f
C248 VDD2.n50 B 0.012187f
C249 VDD2.n51 B 0.027205f
C250 VDD2.n52 B 0.056849f
C251 VDD2.n53 B 0.012187f
C252 VDD2.n54 B 0.01151f
C253 VDD2.n55 B 0.049509f
C254 VDD2.n56 B 0.057031f
C255 VDD2.t0 B 0.18077f
C256 VDD2.t5 B 0.18077f
C257 VDD2.n57 B 1.60495f
C258 VDD2.n58 B 2.61882f
C259 VDD2.n59 B 0.02895f
C260 VDD2.n60 B 0.021419f
C261 VDD2.n61 B 0.01151f
C262 VDD2.n62 B 0.027205f
C263 VDD2.n63 B 0.012187f
C264 VDD2.n64 B 0.021419f
C265 VDD2.n65 B 0.01151f
C266 VDD2.n66 B 0.027205f
C267 VDD2.n67 B 0.012187f
C268 VDD2.n68 B 0.021419f
C269 VDD2.n69 B 0.01151f
C270 VDD2.n70 B 0.027205f
C271 VDD2.n71 B 0.027205f
C272 VDD2.n72 B 0.012187f
C273 VDD2.n73 B 0.021419f
C274 VDD2.n74 B 0.01151f
C275 VDD2.n75 B 0.027205f
C276 VDD2.n76 B 0.012187f
C277 VDD2.n77 B 0.143576f
C278 VDD2.t1 B 0.045795f
C279 VDD2.n78 B 0.020404f
C280 VDD2.n79 B 0.019232f
C281 VDD2.n80 B 0.01151f
C282 VDD2.n81 B 0.954799f
C283 VDD2.n82 B 0.021419f
C284 VDD2.n83 B 0.01151f
C285 VDD2.n84 B 0.012187f
C286 VDD2.n85 B 0.027205f
C287 VDD2.n86 B 0.027205f
C288 VDD2.n87 B 0.012187f
C289 VDD2.n88 B 0.01151f
C290 VDD2.n89 B 0.021419f
C291 VDD2.n90 B 0.021419f
C292 VDD2.n91 B 0.01151f
C293 VDD2.n92 B 0.012187f
C294 VDD2.n93 B 0.027205f
C295 VDD2.n94 B 0.027205f
C296 VDD2.n95 B 0.012187f
C297 VDD2.n96 B 0.01151f
C298 VDD2.n97 B 0.021419f
C299 VDD2.n98 B 0.021419f
C300 VDD2.n99 B 0.01151f
C301 VDD2.n100 B 0.011848f
C302 VDD2.n101 B 0.011848f
C303 VDD2.n102 B 0.027205f
C304 VDD2.n103 B 0.027205f
C305 VDD2.n104 B 0.012187f
C306 VDD2.n105 B 0.01151f
C307 VDD2.n106 B 0.021419f
C308 VDD2.n107 B 0.021419f
C309 VDD2.n108 B 0.01151f
C310 VDD2.n109 B 0.012187f
C311 VDD2.n110 B 0.027205f
C312 VDD2.n111 B 0.056849f
C313 VDD2.n112 B 0.012187f
C314 VDD2.n113 B 0.01151f
C315 VDD2.n114 B 0.049509f
C316 VDD2.n115 B 0.046388f
C317 VDD2.n116 B 2.35797f
C318 VDD2.t4 B 0.18077f
C319 VDD2.t3 B 0.18077f
C320 VDD2.n117 B 1.60492f
C321 VTAIL.t9 B 0.21093f
C322 VTAIL.t6 B 0.21093f
C323 VTAIL.n0 B 1.79244f
C324 VTAIL.n1 B 0.495013f
C325 VTAIL.n2 B 0.03378f
C326 VTAIL.n3 B 0.024993f
C327 VTAIL.n4 B 0.01343f
C328 VTAIL.n5 B 0.031744f
C329 VTAIL.n6 B 0.01422f
C330 VTAIL.n7 B 0.024993f
C331 VTAIL.n8 B 0.01343f
C332 VTAIL.n9 B 0.031744f
C333 VTAIL.n10 B 0.01422f
C334 VTAIL.n11 B 0.024993f
C335 VTAIL.n12 B 0.01343f
C336 VTAIL.n13 B 0.031744f
C337 VTAIL.n14 B 0.01422f
C338 VTAIL.n15 B 0.024993f
C339 VTAIL.n16 B 0.01343f
C340 VTAIL.n17 B 0.031744f
C341 VTAIL.n18 B 0.01422f
C342 VTAIL.n19 B 0.16753f
C343 VTAIL.t1 B 0.053436f
C344 VTAIL.n20 B 0.023808f
C345 VTAIL.n21 B 0.02244f
C346 VTAIL.n22 B 0.01343f
C347 VTAIL.n23 B 1.1141f
C348 VTAIL.n24 B 0.024993f
C349 VTAIL.n25 B 0.01343f
C350 VTAIL.n26 B 0.01422f
C351 VTAIL.n27 B 0.031744f
C352 VTAIL.n28 B 0.031744f
C353 VTAIL.n29 B 0.01422f
C354 VTAIL.n30 B 0.01343f
C355 VTAIL.n31 B 0.024993f
C356 VTAIL.n32 B 0.024993f
C357 VTAIL.n33 B 0.01343f
C358 VTAIL.n34 B 0.01422f
C359 VTAIL.n35 B 0.031744f
C360 VTAIL.n36 B 0.031744f
C361 VTAIL.n37 B 0.031744f
C362 VTAIL.n38 B 0.01422f
C363 VTAIL.n39 B 0.01343f
C364 VTAIL.n40 B 0.024993f
C365 VTAIL.n41 B 0.024993f
C366 VTAIL.n42 B 0.01343f
C367 VTAIL.n43 B 0.013825f
C368 VTAIL.n44 B 0.013825f
C369 VTAIL.n45 B 0.031744f
C370 VTAIL.n46 B 0.031744f
C371 VTAIL.n47 B 0.01422f
C372 VTAIL.n48 B 0.01343f
C373 VTAIL.n49 B 0.024993f
C374 VTAIL.n50 B 0.024993f
C375 VTAIL.n51 B 0.01343f
C376 VTAIL.n52 B 0.01422f
C377 VTAIL.n53 B 0.031744f
C378 VTAIL.n54 B 0.066334f
C379 VTAIL.n55 B 0.01422f
C380 VTAIL.n56 B 0.01343f
C381 VTAIL.n57 B 0.057769f
C382 VTAIL.n58 B 0.036871f
C383 VTAIL.n59 B 0.475727f
C384 VTAIL.t11 B 0.21093f
C385 VTAIL.t0 B 0.21093f
C386 VTAIL.n60 B 1.79244f
C387 VTAIL.n61 B 2.15825f
C388 VTAIL.t5 B 0.21093f
C389 VTAIL.t7 B 0.21093f
C390 VTAIL.n62 B 1.79245f
C391 VTAIL.n63 B 2.15824f
C392 VTAIL.n64 B 0.03378f
C393 VTAIL.n65 B 0.024993f
C394 VTAIL.n66 B 0.01343f
C395 VTAIL.n67 B 0.031744f
C396 VTAIL.n68 B 0.01422f
C397 VTAIL.n69 B 0.024993f
C398 VTAIL.n70 B 0.01343f
C399 VTAIL.n71 B 0.031744f
C400 VTAIL.n72 B 0.01422f
C401 VTAIL.n73 B 0.024993f
C402 VTAIL.n74 B 0.01343f
C403 VTAIL.n75 B 0.031744f
C404 VTAIL.n76 B 0.031744f
C405 VTAIL.n77 B 0.01422f
C406 VTAIL.n78 B 0.024993f
C407 VTAIL.n79 B 0.01343f
C408 VTAIL.n80 B 0.031744f
C409 VTAIL.n81 B 0.01422f
C410 VTAIL.n82 B 0.16753f
C411 VTAIL.t10 B 0.053436f
C412 VTAIL.n83 B 0.023808f
C413 VTAIL.n84 B 0.02244f
C414 VTAIL.n85 B 0.01343f
C415 VTAIL.n86 B 1.1141f
C416 VTAIL.n87 B 0.024993f
C417 VTAIL.n88 B 0.01343f
C418 VTAIL.n89 B 0.01422f
C419 VTAIL.n90 B 0.031744f
C420 VTAIL.n91 B 0.031744f
C421 VTAIL.n92 B 0.01422f
C422 VTAIL.n93 B 0.01343f
C423 VTAIL.n94 B 0.024993f
C424 VTAIL.n95 B 0.024993f
C425 VTAIL.n96 B 0.01343f
C426 VTAIL.n97 B 0.01422f
C427 VTAIL.n98 B 0.031744f
C428 VTAIL.n99 B 0.031744f
C429 VTAIL.n100 B 0.01422f
C430 VTAIL.n101 B 0.01343f
C431 VTAIL.n102 B 0.024993f
C432 VTAIL.n103 B 0.024993f
C433 VTAIL.n104 B 0.01343f
C434 VTAIL.n105 B 0.013825f
C435 VTAIL.n106 B 0.013825f
C436 VTAIL.n107 B 0.031744f
C437 VTAIL.n108 B 0.031744f
C438 VTAIL.n109 B 0.01422f
C439 VTAIL.n110 B 0.01343f
C440 VTAIL.n111 B 0.024993f
C441 VTAIL.n112 B 0.024993f
C442 VTAIL.n113 B 0.01343f
C443 VTAIL.n114 B 0.01422f
C444 VTAIL.n115 B 0.031744f
C445 VTAIL.n116 B 0.066334f
C446 VTAIL.n117 B 0.01422f
C447 VTAIL.n118 B 0.01343f
C448 VTAIL.n119 B 0.057769f
C449 VTAIL.n120 B 0.036871f
C450 VTAIL.n121 B 0.475727f
C451 VTAIL.t2 B 0.21093f
C452 VTAIL.t4 B 0.21093f
C453 VTAIL.n122 B 1.79245f
C454 VTAIL.n123 B 0.698589f
C455 VTAIL.n124 B 0.03378f
C456 VTAIL.n125 B 0.024993f
C457 VTAIL.n126 B 0.01343f
C458 VTAIL.n127 B 0.031744f
C459 VTAIL.n128 B 0.01422f
C460 VTAIL.n129 B 0.024993f
C461 VTAIL.n130 B 0.01343f
C462 VTAIL.n131 B 0.031744f
C463 VTAIL.n132 B 0.01422f
C464 VTAIL.n133 B 0.024993f
C465 VTAIL.n134 B 0.01343f
C466 VTAIL.n135 B 0.031744f
C467 VTAIL.n136 B 0.031744f
C468 VTAIL.n137 B 0.01422f
C469 VTAIL.n138 B 0.024993f
C470 VTAIL.n139 B 0.01343f
C471 VTAIL.n140 B 0.031744f
C472 VTAIL.n141 B 0.01422f
C473 VTAIL.n142 B 0.16753f
C474 VTAIL.t3 B 0.053436f
C475 VTAIL.n143 B 0.023808f
C476 VTAIL.n144 B 0.02244f
C477 VTAIL.n145 B 0.01343f
C478 VTAIL.n146 B 1.1141f
C479 VTAIL.n147 B 0.024993f
C480 VTAIL.n148 B 0.01343f
C481 VTAIL.n149 B 0.01422f
C482 VTAIL.n150 B 0.031744f
C483 VTAIL.n151 B 0.031744f
C484 VTAIL.n152 B 0.01422f
C485 VTAIL.n153 B 0.01343f
C486 VTAIL.n154 B 0.024993f
C487 VTAIL.n155 B 0.024993f
C488 VTAIL.n156 B 0.01343f
C489 VTAIL.n157 B 0.01422f
C490 VTAIL.n158 B 0.031744f
C491 VTAIL.n159 B 0.031744f
C492 VTAIL.n160 B 0.01422f
C493 VTAIL.n161 B 0.01343f
C494 VTAIL.n162 B 0.024993f
C495 VTAIL.n163 B 0.024993f
C496 VTAIL.n164 B 0.01343f
C497 VTAIL.n165 B 0.013825f
C498 VTAIL.n166 B 0.013825f
C499 VTAIL.n167 B 0.031744f
C500 VTAIL.n168 B 0.031744f
C501 VTAIL.n169 B 0.01422f
C502 VTAIL.n170 B 0.01343f
C503 VTAIL.n171 B 0.024993f
C504 VTAIL.n172 B 0.024993f
C505 VTAIL.n173 B 0.01343f
C506 VTAIL.n174 B 0.01422f
C507 VTAIL.n175 B 0.031744f
C508 VTAIL.n176 B 0.066334f
C509 VTAIL.n177 B 0.01422f
C510 VTAIL.n178 B 0.01343f
C511 VTAIL.n179 B 0.057769f
C512 VTAIL.n180 B 0.036871f
C513 VTAIL.n181 B 1.65769f
C514 VTAIL.n182 B 0.03378f
C515 VTAIL.n183 B 0.024993f
C516 VTAIL.n184 B 0.01343f
C517 VTAIL.n185 B 0.031744f
C518 VTAIL.n186 B 0.01422f
C519 VTAIL.n187 B 0.024993f
C520 VTAIL.n188 B 0.01343f
C521 VTAIL.n189 B 0.031744f
C522 VTAIL.n190 B 0.01422f
C523 VTAIL.n191 B 0.024993f
C524 VTAIL.n192 B 0.01343f
C525 VTAIL.n193 B 0.031744f
C526 VTAIL.n194 B 0.01422f
C527 VTAIL.n195 B 0.024993f
C528 VTAIL.n196 B 0.01343f
C529 VTAIL.n197 B 0.031744f
C530 VTAIL.n198 B 0.01422f
C531 VTAIL.n199 B 0.16753f
C532 VTAIL.t8 B 0.053436f
C533 VTAIL.n200 B 0.023808f
C534 VTAIL.n201 B 0.02244f
C535 VTAIL.n202 B 0.01343f
C536 VTAIL.n203 B 1.1141f
C537 VTAIL.n204 B 0.024993f
C538 VTAIL.n205 B 0.01343f
C539 VTAIL.n206 B 0.01422f
C540 VTAIL.n207 B 0.031744f
C541 VTAIL.n208 B 0.031744f
C542 VTAIL.n209 B 0.01422f
C543 VTAIL.n210 B 0.01343f
C544 VTAIL.n211 B 0.024993f
C545 VTAIL.n212 B 0.024993f
C546 VTAIL.n213 B 0.01343f
C547 VTAIL.n214 B 0.01422f
C548 VTAIL.n215 B 0.031744f
C549 VTAIL.n216 B 0.031744f
C550 VTAIL.n217 B 0.031744f
C551 VTAIL.n218 B 0.01422f
C552 VTAIL.n219 B 0.01343f
C553 VTAIL.n220 B 0.024993f
C554 VTAIL.n221 B 0.024993f
C555 VTAIL.n222 B 0.01343f
C556 VTAIL.n223 B 0.013825f
C557 VTAIL.n224 B 0.013825f
C558 VTAIL.n225 B 0.031744f
C559 VTAIL.n226 B 0.031744f
C560 VTAIL.n227 B 0.01422f
C561 VTAIL.n228 B 0.01343f
C562 VTAIL.n229 B 0.024993f
C563 VTAIL.n230 B 0.024993f
C564 VTAIL.n231 B 0.01343f
C565 VTAIL.n232 B 0.01422f
C566 VTAIL.n233 B 0.031744f
C567 VTAIL.n234 B 0.066334f
C568 VTAIL.n235 B 0.01422f
C569 VTAIL.n236 B 0.01343f
C570 VTAIL.n237 B 0.057769f
C571 VTAIL.n238 B 0.036871f
C572 VTAIL.n239 B 1.58357f
C573 VN.n0 B 0.03586f
C574 VN.t0 B 2.02935f
C575 VN.n1 B 0.037702f
C576 VN.n2 B 0.01907f
C577 VN.n3 B 0.035363f
C578 VN.t3 B 2.30108f
C579 VN.t5 B 2.02935f
C580 VN.n4 B 0.793037f
C581 VN.n5 B 0.753872f
C582 VN.n6 B 0.242772f
C583 VN.n7 B 0.01907f
C584 VN.n8 B 0.035363f
C585 VN.n9 B 0.037702f
C586 VN.n10 B 0.015402f
C587 VN.n11 B 0.01907f
C588 VN.n12 B 0.01907f
C589 VN.n13 B 0.01907f
C590 VN.n14 B 0.035363f
C591 VN.n15 B 0.035363f
C592 VN.n16 B 0.799645f
C593 VN.n17 B 0.053613f
C594 VN.n18 B 0.03586f
C595 VN.t4 B 2.02935f
C596 VN.n19 B 0.037702f
C597 VN.n20 B 0.01907f
C598 VN.n21 B 0.035363f
C599 VN.t2 B 2.30108f
C600 VN.t1 B 2.02935f
C601 VN.n22 B 0.793037f
C602 VN.n23 B 0.753872f
C603 VN.n24 B 0.242772f
C604 VN.n25 B 0.01907f
C605 VN.n26 B 0.035363f
C606 VN.n27 B 0.037702f
C607 VN.n28 B 0.015402f
C608 VN.n29 B 0.01907f
C609 VN.n30 B 0.01907f
C610 VN.n31 B 0.01907f
C611 VN.n32 B 0.035363f
C612 VN.n33 B 0.035363f
C613 VN.n34 B 0.799645f
C614 VN.n35 B 1.17227f
.ends

