* NGSPICE file created from opamp_sample_0011.ext - technology: sky130A

.subckt opamp_sample_0011 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VOUT.t42 CS_BIAS.t32 GND.t149 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X1 VOUT.t41 CS_BIAS.t33 GND.t148 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X2 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 a_n1431_n2782.t1 GND.t2 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=1.9305 ps=10.68 w=4.95 l=2.4
X3 a_n12440_8296.t10 VN.t2 a_n4178_n267.t3 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X4 VOUT.t40 CS_BIAS.t34 GND.t147 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X5 GND.t146 CS_BIAS.t35 VOUT.t39 GND.t120 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X6 a_n12440_8296.t9 VN.t3 a_n4178_n267.t8 GND.t84 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X7 a_n12440_8296.t8 VN.t4 a_n4178_n267.t10 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=4.7
X8 VOUT.t9 a_n12440_8296.t14 VDD.t104 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=1.3728 ps=7.82 w=3.52 l=4.06
X9 VOUT.t38 CS_BIAS.t36 GND.t144 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X10 CS_BIAS.t19 CS_BIAS.t18 GND.t145 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X11 GND.t81 GND.t78 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.4
X12 GND.t143 CS_BIAS.t37 VOUT.t37 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X13 VN.t1 GND.t75 GND.t77 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X14 VDD.t13 a_n6715_8686.t20 a_n6793_8883.t7 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X15 a_n6793_8883.t13 a_n6715_8686.t14 a_n6715_8686.t15 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X16 GND.t74 GND.t72 GND.t73 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X17 VP.t1 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X18 a_n4178_n267.t2 VP.t2 a_n6715_8686.t2 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=4.7
X19 a_n3792_7061.t14 a_n6715_8686.t21 a_n12440_8296.t12 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X20 VDD.t103 a_n12440_8296.t15 VOUT.t43 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=0.5808 ps=3.85 w=3.52 l=4.06
X21 VDD.t81 VDD.t79 VDD.t80 VDD.t49 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X22 GND.t142 CS_BIAS.t38 VOUT.t36 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X23 VOUT.t2 a_n12440_8296.t16 VDD.t102 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=1.3728 ps=7.82 w=3.52 l=4.06
X24 a_n12440_8296.t13 a_n6715_8686.t22 a_n3792_7061.t13 VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X25 a_n6793_8883.t6 a_n6715_8686.t23 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X26 VDD.t101 a_n12440_8296.t17 VOUT.t0 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=0.5808 ps=3.85 w=3.52 l=4.06
X27 VOUT.t3 a_n12440_8296.t18 VDD.t100 VDD.t90 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0.5808 ps=3.85 w=3.52 l=4.06
X28 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 a_n1431_n2782.t0 GND.t85 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=1.9305 ps=10.68 w=4.95 l=2.4
X29 VDD.t24 a_n6715_8686.t24 a_n3792_7061.t8 VDD.t23 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X30 a_n6793_8883.t12 a_n6715_8686.t10 a_n6715_8686.t11 VDD.t1 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X31 VOUT.t7 a_n12440_8296.t19 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=1.3728 ps=7.82 w=3.52 l=4.06
X32 VDD.t78 VDD.t76 VDD.t77 VDD.t35 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X33 GND.t141 CS_BIAS.t39 VOUT.t35 GND.t90 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X34 a_n3792_7061.t7 a_n6715_8686.t25 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X35 a_6921_8883# a_6921_8883# a_6921_8883# VDD.t109 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=4.1418 ps=22.8 w=5.31 l=3.38
X36 VDD.t75 VDD.t73 VDD.t74 VDD.t67 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X37 VOUT.t8 a_n12440_8296.t20 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=1.3728 ps=7.82 w=3.52 l=4.06
X38 VDD.t95 a_n12440_8296.t21 VOUT.t6 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=0.5808 ps=3.85 w=3.52 l=4.06
X39 GND.t140 CS_BIAS.t40 VOUT.t34 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X40 GND.t68 GND.t66 GND.t67 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X41 VDD.t93 a_n12440_8296.t22 VOUT.t5 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.5808 pd=3.85 as=0.5808 ps=3.85 w=3.52 l=4.06
X42 GND.t139 CS_BIAS.t24 CS_BIAS.t25 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X43 GND.t138 CS_BIAS.t41 VOUT.t33 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X44 VOUT.t1 a_n12440_8296.t23 VDD.t91 VDD.t90 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0.5808 ps=3.85 w=3.52 l=4.06
X45 VDD.t7 a_n6715_8686.t26 a_n3792_7061.t6 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X46 GND.t65 GND.t63 GND.t64 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X47 a_n4178_n267.t0 VP.t3 a_n6715_8686.t0 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=4.7
X48 VDD.t72 VDD.t70 VDD.t71 VDD.t53 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X49 CS_BIAS.t23 CS_BIAS.t22 GND.t137 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X50 VOUT.t32 CS_BIAS.t42 GND.t136 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X51 a_n4178_n267.t1 VP.t4 a_n6715_8686.t1 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X52 GND.t62 GND.t60 GND.t61 GND.t45 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X53 VDD.t69 VDD.t66 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X54 VOUT.t31 CS_BIAS.t43 GND.t133 GND.t105 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X55 GND.t135 CS_BIAS.t20 CS_BIAS.t21 GND.t120 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X56 a_n12440_8296.t11 a_n6715_8686.t27 a_n3792_7061.t12 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X57 VOUT.t30 CS_BIAS.t44 GND.t134 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X58 a_n3792_7061.t5 a_n6715_8686.t28 VDD.t113 VDD.t112 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X59 VDD.t22 a_n6715_8686.t29 a_n6793_8883.t5 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X60 GND.t59 GND.t57 GND.t58 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X61 a_n4178_n267.t11 DIFFPAIR_BIAS.t4 a_n689_n2782.t1 GND.t83 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=1.9305 ps=10.68 w=4.95 l=2.4
X62 VDD.t65 VDD.t63 VDD.t64 VDD.t60 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X63 GND.t132 CS_BIAS.t8 CS_BIAS.t9 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X64 GND.t131 CS_BIAS.t45 VOUT.t29 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X65 a_n6793_8883.t4 a_n6715_8686.t30 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X66 GND.t130 CS_BIAS.t6 CS_BIAS.t7 GND.t90 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X67 GND.t129 CS_BIAS.t46 VOUT.t28 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X68 a_n12440_8296.t7 VN.t5 a_n4178_n267.t5 GND.t82 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=4.7
X69 CS_BIAS.t5 CS_BIAS.t4 GND.t128 GND.t105 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X70 CS_BIAS.t3 CS_BIAS.t2 GND.t127 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X71 a_n4178_n267.t9 VN.t6 a_n12440_8296.t6 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X72 VOUT.t27 CS_BIAS.t47 GND.t126 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X73 GND.t56 GND.t54 GND.t55 GND.t24 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=4.7
X74 a_n12440_8296.t2 a_n6715_8686.t31 a_n3792_7061.t11 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X75 VDD.t62 VDD.t59 VDD.t61 VDD.t60 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X76 GND.t125 CS_BIAS.t0 CS_BIAS.t1 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X77 a_n6715_8686.t9 a_n6715_8686.t8 a_n6793_8883.t11 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X78 GND.t53 GND.t51 GND.t52 GND.t45 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X79 a_n6715_8686.t19 VP.t5 a_n4178_n267.t17 GND.t84 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X80 GND.t50 GND.t48 GND.t49 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=4.7
X81 VOUT.t26 CS_BIAS.t48 GND.t124 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X82 VDD.t86 a_n6715_8686.t32 a_n3792_7061.t4 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X83 GND.t123 CS_BIAS.t49 VOUT.t25 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X84 GND.t47 GND.t44 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X85 GND.t116 CS_BIAS.t50 VOUT.t24 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X86 GND.t43 GND.t41 VP.t0 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X87 GND.t121 CS_BIAS.t51 VOUT.t23 GND.t120 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X88 a_n6793_8883.t10 a_n6715_8686.t4 a_n6715_8686.t5 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X89 GND.t119 CS_BIAS.t16 CS_BIAS.t17 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X90 a_n3792_7061.t3 a_n6715_8686.t33 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X91 VDD.t58 VDD.t56 VDD.t57 VDD.t45 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X92 a_n3792_7061.t2 a_n6715_8686.t34 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X93 CS_BIAS.t15 CS_BIAS.t14 GND.t118 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X94 VOUT.t22 CS_BIAS.t52 GND.t115 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X95 VDD.t83 a_n6715_8686.t35 a_n6793_8883.t3 VDD.t82 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X96 CS_BIAS.t31 CS_BIAS.t30 GND.t114 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X97 GND.t113 CS_BIAS.t28 CS_BIAS.t29 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X98 a_n6715_8686.t7 a_n6715_8686.t6 a_n6793_8883.t9 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X99 a_n6715_8686.t17 VP.t6 a_n4178_n267.t15 GND.t3 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X100 a_n6715_8686.t18 VP.t7 a_n4178_n267.t16 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=4.7
X101 a_n6793_8883.t8 a_n6715_8686.t12 a_n6715_8686.t13 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X102 VDD.t20 a_n6715_8686.t36 a_n3792_7061.t1 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.38
X103 a_n3792_7061.t10 a_n6715_8686.t37 a_n12440_8296.t0 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X104 a_n6793_8883.t2 a_n6715_8686.t38 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X105 GND.t111 CS_BIAS.t53 VOUT.t21 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X106 a_n6793_8883.t1 a_n6715_8686.t39 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X107 VDD.t55 VDD.t52 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X108 a_n4178_n267.t7 VN.t7 a_n12440_8296.t5 GND.t1 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=4.7
X109 VDD.t51 VDD.t48 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X110 a_n4178_n267.t6 VN.t8 a_n12440_8296.t4 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X111 a_n4178_n267.t4 VN.t9 a_n12440_8296.t3 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=4.7
X112 GND.t109 CS_BIAS.t54 VOUT.t20 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X113 GND.t107 CS_BIAS.t26 CS_BIAS.t27 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X114 GND.t40 GND.t37 GND.t39 GND.t38 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=0 ps=0 w=4.95 l=2.4
X115 GND.t36 GND.t33 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X116 VOUT.t19 CS_BIAS.t55 GND.t106 GND.t105 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X117 a_n7753_8883# a_n7753_8883# a_n7753_8883# VDD.t84 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=4.1418 ps=22.8 w=5.31 l=3.38
X118 GND.t32 GND.t30 GND.t31 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X119 CS_BIAS.t11 CS_BIAS.t10 GND.t104 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X120 VOUT.t18 CS_BIAS.t56 GND.t97 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X121 VOUT.t17 CS_BIAS.t57 GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X122 VOUT.t44 a_n3792_7061.t0 sky130_fd_pr__cap_mim_m3_1 l=18.2 w=9.26
X123 VOUT.t16 CS_BIAS.t58 GND.t101 GND.t100 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X124 a_n12440_8296.t1 a_n6715_8686.t40 a_n3792_7061.t9 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.38
X125 GND.t99 CS_BIAS.t59 VOUT.t15 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X126 VDD.t47 VDD.t44 VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X127 GND.t29 GND.t27 GND.t28 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X128 VDD.t43 VDD.t41 VDD.t42 VDD.t31 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X129 VDD.t40 VDD.t38 VDD.t39 VDD.t27 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X130 a_n4178_n267.t12 DIFFPAIR_BIAS.t5 a_n689_n2782.t0 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.9305 pd=10.68 as=1.9305 ps=10.68 w=4.95 l=2.4
X131 a_n6715_8686.t3 VP.t8 a_n4178_n267.t13 GND.t82 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=4.7
X132 a_n4178_n267.t14 VP.t9 a_n6715_8686.t16 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.65175 pd=4.28 as=0.65175 ps=4.28 w=3.95 l=4.7
X133 CS_BIAS.t13 CS_BIAS.t12 GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X134 VOUT.t14 CS_BIAS.t60 GND.t93 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=1.3143 ps=7.52 w=3.37 l=5.45
X135 GND.t26 GND.t23 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=4.7
X136 VDD.t37 VDD.t34 VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.38
X137 VOUT.t4 a_n12440_8296.t24 VDD.t89 VDD.t87 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0.5808 ps=3.85 w=3.52 l=4.06
X138 GND.t22 GND.t19 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X139 GND.t14 GND.t12 VN.t0 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X140 VDD.t33 VDD.t30 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X141 GND.t18 GND.t15 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=4.7
X142 VDD.t29 VDD.t26 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0 ps=0 w=3.52 l=4.06
X143 GND.t11 GND.t8 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0 ps=0 w=3.37 l=5.45
X144 VOUT.t45 a_n3792_7061.t0 sky130_fd_pr__cap_mim_m3_1 l=18.2 w=9.26
X145 VOUT.t10 a_n12440_8296.t25 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=1.3728 pd=7.82 as=0.5808 ps=3.85 w=3.52 l=4.06
X146 GND.t91 CS_BIAS.t61 VOUT.t13 GND.t90 sky130_fd_pr__nfet_01v8 ad=1.3143 pd=7.52 as=0.55605 ps=3.7 w=3.37 l=5.45
X147 GND.t89 CS_BIAS.t62 VOUT.t12 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
X148 VDD.t111 a_n6715_8686.t41 a_n6793_8883.t0 VDD.t110 sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.38
X149 VOUT.t11 CS_BIAS.t63 GND.t87 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.55605 pd=3.7 as=0.55605 ps=3.7 w=3.37 l=5.45
R0 CS_BIAS.n447 CS_BIAS.n446 161.3
R1 CS_BIAS.n445 CS_BIAS.n303 161.3
R2 CS_BIAS.n444 CS_BIAS.n443 161.3
R3 CS_BIAS.n442 CS_BIAS.n304 161.3
R4 CS_BIAS.n441 CS_BIAS.n440 161.3
R5 CS_BIAS.n439 CS_BIAS.n305 161.3
R6 CS_BIAS.n438 CS_BIAS.n437 161.3
R7 CS_BIAS.n436 CS_BIAS.n306 161.3
R8 CS_BIAS.n435 CS_BIAS.n434 161.3
R9 CS_BIAS.n433 CS_BIAS.n307 161.3
R10 CS_BIAS.n432 CS_BIAS.n431 161.3
R11 CS_BIAS.n430 CS_BIAS.n308 161.3
R12 CS_BIAS.n429 CS_BIAS.n428 161.3
R13 CS_BIAS.n427 CS_BIAS.n309 161.3
R14 CS_BIAS.n426 CS_BIAS.n425 161.3
R15 CS_BIAS.n424 CS_BIAS.n311 161.3
R16 CS_BIAS.n423 CS_BIAS.n422 161.3
R17 CS_BIAS.n421 CS_BIAS.n312 161.3
R18 CS_BIAS.n420 CS_BIAS.n419 161.3
R19 CS_BIAS.n418 CS_BIAS.n313 161.3
R20 CS_BIAS.n417 CS_BIAS.n416 161.3
R21 CS_BIAS.n415 CS_BIAS.n314 161.3
R22 CS_BIAS.n414 CS_BIAS.n413 161.3
R23 CS_BIAS.n412 CS_BIAS.n411 161.3
R24 CS_BIAS.n410 CS_BIAS.n316 161.3
R25 CS_BIAS.n409 CS_BIAS.n408 161.3
R26 CS_BIAS.n407 CS_BIAS.n317 161.3
R27 CS_BIAS.n406 CS_BIAS.n405 161.3
R28 CS_BIAS.n404 CS_BIAS.n318 161.3
R29 CS_BIAS.n403 CS_BIAS.n402 161.3
R30 CS_BIAS.n401 CS_BIAS.n319 161.3
R31 CS_BIAS.n400 CS_BIAS.n399 161.3
R32 CS_BIAS.n398 CS_BIAS.n320 161.3
R33 CS_BIAS.n397 CS_BIAS.n396 161.3
R34 CS_BIAS.n395 CS_BIAS.n321 161.3
R35 CS_BIAS.n394 CS_BIAS.n393 161.3
R36 CS_BIAS.n392 CS_BIAS.n322 161.3
R37 CS_BIAS.n391 CS_BIAS.n390 161.3
R38 CS_BIAS.n389 CS_BIAS.n324 161.3
R39 CS_BIAS.n388 CS_BIAS.n387 161.3
R40 CS_BIAS.n386 CS_BIAS.n325 161.3
R41 CS_BIAS.n385 CS_BIAS.n384 161.3
R42 CS_BIAS.n383 CS_BIAS.n326 161.3
R43 CS_BIAS.n382 CS_BIAS.n381 161.3
R44 CS_BIAS.n380 CS_BIAS.n327 161.3
R45 CS_BIAS.n379 CS_BIAS.n378 161.3
R46 CS_BIAS.n377 CS_BIAS.n376 161.3
R47 CS_BIAS.n375 CS_BIAS.n329 161.3
R48 CS_BIAS.n374 CS_BIAS.n373 161.3
R49 CS_BIAS.n372 CS_BIAS.n330 161.3
R50 CS_BIAS.n371 CS_BIAS.n370 161.3
R51 CS_BIAS.n369 CS_BIAS.n331 161.3
R52 CS_BIAS.n368 CS_BIAS.n367 161.3
R53 CS_BIAS.n366 CS_BIAS.n332 161.3
R54 CS_BIAS.n365 CS_BIAS.n364 161.3
R55 CS_BIAS.n363 CS_BIAS.n333 161.3
R56 CS_BIAS.n362 CS_BIAS.n361 161.3
R57 CS_BIAS.n360 CS_BIAS.n334 161.3
R58 CS_BIAS.n359 CS_BIAS.n358 161.3
R59 CS_BIAS.n357 CS_BIAS.n335 161.3
R60 CS_BIAS.n356 CS_BIAS.n355 161.3
R61 CS_BIAS.n354 CS_BIAS.n337 161.3
R62 CS_BIAS.n353 CS_BIAS.n352 161.3
R63 CS_BIAS.n351 CS_BIAS.n338 161.3
R64 CS_BIAS.n350 CS_BIAS.n349 161.3
R65 CS_BIAS.n348 CS_BIAS.n339 161.3
R66 CS_BIAS.n347 CS_BIAS.n346 161.3
R67 CS_BIAS.n345 CS_BIAS.n340 161.3
R68 CS_BIAS.n344 CS_BIAS.n343 161.3
R69 CS_BIAS.n65 CS_BIAS.n64 161.3
R70 CS_BIAS.n66 CS_BIAS.n61 161.3
R71 CS_BIAS.n68 CS_BIAS.n67 161.3
R72 CS_BIAS.n69 CS_BIAS.n60 161.3
R73 CS_BIAS.n71 CS_BIAS.n70 161.3
R74 CS_BIAS.n72 CS_BIAS.n59 161.3
R75 CS_BIAS.n74 CS_BIAS.n73 161.3
R76 CS_BIAS.n75 CS_BIAS.n58 161.3
R77 CS_BIAS.n77 CS_BIAS.n76 161.3
R78 CS_BIAS.n78 CS_BIAS.n56 161.3
R79 CS_BIAS.n80 CS_BIAS.n79 161.3
R80 CS_BIAS.n81 CS_BIAS.n55 161.3
R81 CS_BIAS.n83 CS_BIAS.n82 161.3
R82 CS_BIAS.n84 CS_BIAS.n54 161.3
R83 CS_BIAS.n86 CS_BIAS.n85 161.3
R84 CS_BIAS.n87 CS_BIAS.n53 161.3
R85 CS_BIAS.n89 CS_BIAS.n88 161.3
R86 CS_BIAS.n90 CS_BIAS.n52 161.3
R87 CS_BIAS.n92 CS_BIAS.n91 161.3
R88 CS_BIAS.n93 CS_BIAS.n51 161.3
R89 CS_BIAS.n95 CS_BIAS.n94 161.3
R90 CS_BIAS.n96 CS_BIAS.n50 161.3
R91 CS_BIAS.n98 CS_BIAS.n97 161.3
R92 CS_BIAS.n100 CS_BIAS.n99 161.3
R93 CS_BIAS.n101 CS_BIAS.n48 161.3
R94 CS_BIAS.n103 CS_BIAS.n102 161.3
R95 CS_BIAS.n104 CS_BIAS.n47 161.3
R96 CS_BIAS.n106 CS_BIAS.n105 161.3
R97 CS_BIAS.n107 CS_BIAS.n46 161.3
R98 CS_BIAS.n109 CS_BIAS.n108 161.3
R99 CS_BIAS.n110 CS_BIAS.n45 161.3
R100 CS_BIAS.n112 CS_BIAS.n111 161.3
R101 CS_BIAS.n113 CS_BIAS.n43 161.3
R102 CS_BIAS.n115 CS_BIAS.n114 161.3
R103 CS_BIAS.n116 CS_BIAS.n42 161.3
R104 CS_BIAS.n118 CS_BIAS.n117 161.3
R105 CS_BIAS.n119 CS_BIAS.n41 161.3
R106 CS_BIAS.n121 CS_BIAS.n120 161.3
R107 CS_BIAS.n122 CS_BIAS.n40 161.3
R108 CS_BIAS.n124 CS_BIAS.n123 161.3
R109 CS_BIAS.n125 CS_BIAS.n39 161.3
R110 CS_BIAS.n127 CS_BIAS.n126 161.3
R111 CS_BIAS.n128 CS_BIAS.n38 161.3
R112 CS_BIAS.n130 CS_BIAS.n129 161.3
R113 CS_BIAS.n131 CS_BIAS.n37 161.3
R114 CS_BIAS.n133 CS_BIAS.n132 161.3
R115 CS_BIAS.n135 CS_BIAS.n134 161.3
R116 CS_BIAS.n136 CS_BIAS.n35 161.3
R117 CS_BIAS.n138 CS_BIAS.n137 161.3
R118 CS_BIAS.n139 CS_BIAS.n34 161.3
R119 CS_BIAS.n141 CS_BIAS.n140 161.3
R120 CS_BIAS.n142 CS_BIAS.n33 161.3
R121 CS_BIAS.n144 CS_BIAS.n143 161.3
R122 CS_BIAS.n145 CS_BIAS.n32 161.3
R123 CS_BIAS.n147 CS_BIAS.n146 161.3
R124 CS_BIAS.n148 CS_BIAS.n30 161.3
R125 CS_BIAS.n150 CS_BIAS.n149 161.3
R126 CS_BIAS.n151 CS_BIAS.n29 161.3
R127 CS_BIAS.n153 CS_BIAS.n152 161.3
R128 CS_BIAS.n154 CS_BIAS.n28 161.3
R129 CS_BIAS.n156 CS_BIAS.n155 161.3
R130 CS_BIAS.n157 CS_BIAS.n27 161.3
R131 CS_BIAS.n159 CS_BIAS.n158 161.3
R132 CS_BIAS.n160 CS_BIAS.n26 161.3
R133 CS_BIAS.n162 CS_BIAS.n161 161.3
R134 CS_BIAS.n163 CS_BIAS.n25 161.3
R135 CS_BIAS.n165 CS_BIAS.n164 161.3
R136 CS_BIAS.n166 CS_BIAS.n24 161.3
R137 CS_BIAS.n168 CS_BIAS.n167 161.3
R138 CS_BIAS.n197 CS_BIAS.n196 161.3
R139 CS_BIAS.n198 CS_BIAS.n193 161.3
R140 CS_BIAS.n200 CS_BIAS.n199 161.3
R141 CS_BIAS.n201 CS_BIAS.n192 161.3
R142 CS_BIAS.n203 CS_BIAS.n202 161.3
R143 CS_BIAS.n204 CS_BIAS.n191 161.3
R144 CS_BIAS.n206 CS_BIAS.n205 161.3
R145 CS_BIAS.n207 CS_BIAS.n190 161.3
R146 CS_BIAS.n209 CS_BIAS.n208 161.3
R147 CS_BIAS.n210 CS_BIAS.n188 161.3
R148 CS_BIAS.n212 CS_BIAS.n211 161.3
R149 CS_BIAS.n213 CS_BIAS.n187 161.3
R150 CS_BIAS.n215 CS_BIAS.n214 161.3
R151 CS_BIAS.n216 CS_BIAS.n186 161.3
R152 CS_BIAS.n218 CS_BIAS.n217 161.3
R153 CS_BIAS.n219 CS_BIAS.n185 161.3
R154 CS_BIAS.n221 CS_BIAS.n220 161.3
R155 CS_BIAS.n222 CS_BIAS.n184 161.3
R156 CS_BIAS.n224 CS_BIAS.n223 161.3
R157 CS_BIAS.n225 CS_BIAS.n183 161.3
R158 CS_BIAS.n227 CS_BIAS.n226 161.3
R159 CS_BIAS.n228 CS_BIAS.n182 161.3
R160 CS_BIAS.n230 CS_BIAS.n229 161.3
R161 CS_BIAS.n232 CS_BIAS.n231 161.3
R162 CS_BIAS.n233 CS_BIAS.n180 161.3
R163 CS_BIAS.n235 CS_BIAS.n234 161.3
R164 CS_BIAS.n236 CS_BIAS.n179 161.3
R165 CS_BIAS.n238 CS_BIAS.n237 161.3
R166 CS_BIAS.n239 CS_BIAS.n178 161.3
R167 CS_BIAS.n241 CS_BIAS.n240 161.3
R168 CS_BIAS.n242 CS_BIAS.n22 161.3
R169 CS_BIAS.n244 CS_BIAS.n243 161.3
R170 CS_BIAS.n245 CS_BIAS.n20 161.3
R171 CS_BIAS.n247 CS_BIAS.n246 161.3
R172 CS_BIAS.n248 CS_BIAS.n19 161.3
R173 CS_BIAS.n250 CS_BIAS.n249 161.3
R174 CS_BIAS.n251 CS_BIAS.n18 161.3
R175 CS_BIAS.n253 CS_BIAS.n252 161.3
R176 CS_BIAS.n254 CS_BIAS.n17 161.3
R177 CS_BIAS.n256 CS_BIAS.n255 161.3
R178 CS_BIAS.n257 CS_BIAS.n16 161.3
R179 CS_BIAS.n259 CS_BIAS.n258 161.3
R180 CS_BIAS.n260 CS_BIAS.n15 161.3
R181 CS_BIAS.n262 CS_BIAS.n261 161.3
R182 CS_BIAS.n263 CS_BIAS.n14 161.3
R183 CS_BIAS.n265 CS_BIAS.n264 161.3
R184 CS_BIAS.n267 CS_BIAS.n266 161.3
R185 CS_BIAS.n268 CS_BIAS.n12 161.3
R186 CS_BIAS.n270 CS_BIAS.n269 161.3
R187 CS_BIAS.n271 CS_BIAS.n11 161.3
R188 CS_BIAS.n273 CS_BIAS.n272 161.3
R189 CS_BIAS.n274 CS_BIAS.n10 161.3
R190 CS_BIAS.n276 CS_BIAS.n275 161.3
R191 CS_BIAS.n277 CS_BIAS.n9 161.3
R192 CS_BIAS.n279 CS_BIAS.n278 161.3
R193 CS_BIAS.n280 CS_BIAS.n7 161.3
R194 CS_BIAS.n282 CS_BIAS.n281 161.3
R195 CS_BIAS.n283 CS_BIAS.n6 161.3
R196 CS_BIAS.n285 CS_BIAS.n284 161.3
R197 CS_BIAS.n286 CS_BIAS.n5 161.3
R198 CS_BIAS.n288 CS_BIAS.n287 161.3
R199 CS_BIAS.n289 CS_BIAS.n4 161.3
R200 CS_BIAS.n291 CS_BIAS.n290 161.3
R201 CS_BIAS.n292 CS_BIAS.n3 161.3
R202 CS_BIAS.n294 CS_BIAS.n293 161.3
R203 CS_BIAS.n295 CS_BIAS.n2 161.3
R204 CS_BIAS.n297 CS_BIAS.n296 161.3
R205 CS_BIAS.n298 CS_BIAS.n1 161.3
R206 CS_BIAS.n300 CS_BIAS.n299 161.3
R207 CS_BIAS.n897 CS_BIAS.n896 161.3
R208 CS_BIAS.n895 CS_BIAS.n753 161.3
R209 CS_BIAS.n894 CS_BIAS.n893 161.3
R210 CS_BIAS.n892 CS_BIAS.n754 161.3
R211 CS_BIAS.n891 CS_BIAS.n890 161.3
R212 CS_BIAS.n889 CS_BIAS.n755 161.3
R213 CS_BIAS.n888 CS_BIAS.n887 161.3
R214 CS_BIAS.n886 CS_BIAS.n756 161.3
R215 CS_BIAS.n885 CS_BIAS.n884 161.3
R216 CS_BIAS.n883 CS_BIAS.n757 161.3
R217 CS_BIAS.n882 CS_BIAS.n881 161.3
R218 CS_BIAS.n880 CS_BIAS.n758 161.3
R219 CS_BIAS.n879 CS_BIAS.n878 161.3
R220 CS_BIAS.n876 CS_BIAS.n759 161.3
R221 CS_BIAS.n875 CS_BIAS.n874 161.3
R222 CS_BIAS.n873 CS_BIAS.n760 161.3
R223 CS_BIAS.n872 CS_BIAS.n871 161.3
R224 CS_BIAS.n870 CS_BIAS.n761 161.3
R225 CS_BIAS.n869 CS_BIAS.n868 161.3
R226 CS_BIAS.n867 CS_BIAS.n762 161.3
R227 CS_BIAS.n866 CS_BIAS.n865 161.3
R228 CS_BIAS.n864 CS_BIAS.n763 161.3
R229 CS_BIAS.n863 CS_BIAS.n862 161.3
R230 CS_BIAS.n861 CS_BIAS.n860 161.3
R231 CS_BIAS.n859 CS_BIAS.n765 161.3
R232 CS_BIAS.n858 CS_BIAS.n857 161.3
R233 CS_BIAS.n856 CS_BIAS.n766 161.3
R234 CS_BIAS.n855 CS_BIAS.n854 161.3
R235 CS_BIAS.n853 CS_BIAS.n767 161.3
R236 CS_BIAS.n852 CS_BIAS.n851 161.3
R237 CS_BIAS.n850 CS_BIAS.n768 161.3
R238 CS_BIAS.n849 CS_BIAS.n848 161.3
R239 CS_BIAS.n847 CS_BIAS.n769 161.3
R240 CS_BIAS.n846 CS_BIAS.n845 161.3
R241 CS_BIAS.n844 CS_BIAS.n770 161.3
R242 CS_BIAS.n843 CS_BIAS.n842 161.3
R243 CS_BIAS.n840 CS_BIAS.n771 161.3
R244 CS_BIAS.n839 CS_BIAS.n838 161.3
R245 CS_BIAS.n837 CS_BIAS.n772 161.3
R246 CS_BIAS.n836 CS_BIAS.n835 161.3
R247 CS_BIAS.n834 CS_BIAS.n773 161.3
R248 CS_BIAS.n833 CS_BIAS.n832 161.3
R249 CS_BIAS.n831 CS_BIAS.n774 161.3
R250 CS_BIAS.n830 CS_BIAS.n829 161.3
R251 CS_BIAS.n828 CS_BIAS.n775 161.3
R252 CS_BIAS.n827 CS_BIAS.n826 161.3
R253 CS_BIAS.n825 CS_BIAS.n824 161.3
R254 CS_BIAS.n823 CS_BIAS.n777 161.3
R255 CS_BIAS.n822 CS_BIAS.n821 161.3
R256 CS_BIAS.n820 CS_BIAS.n778 161.3
R257 CS_BIAS.n819 CS_BIAS.n818 161.3
R258 CS_BIAS.n817 CS_BIAS.n779 161.3
R259 CS_BIAS.n816 CS_BIAS.n815 161.3
R260 CS_BIAS.n814 CS_BIAS.n780 161.3
R261 CS_BIAS.n813 CS_BIAS.n812 161.3
R262 CS_BIAS.n811 CS_BIAS.n781 161.3
R263 CS_BIAS.n810 CS_BIAS.n809 161.3
R264 CS_BIAS.n808 CS_BIAS.n782 161.3
R265 CS_BIAS.n807 CS_BIAS.n806 161.3
R266 CS_BIAS.n804 CS_BIAS.n783 161.3
R267 CS_BIAS.n803 CS_BIAS.n802 161.3
R268 CS_BIAS.n801 CS_BIAS.n784 161.3
R269 CS_BIAS.n800 CS_BIAS.n799 161.3
R270 CS_BIAS.n798 CS_BIAS.n785 161.3
R271 CS_BIAS.n797 CS_BIAS.n796 161.3
R272 CS_BIAS.n795 CS_BIAS.n786 161.3
R273 CS_BIAS.n794 CS_BIAS.n793 161.3
R274 CS_BIAS.n792 CS_BIAS.n787 161.3
R275 CS_BIAS.n791 CS_BIAS.n790 161.3
R276 CS_BIAS.n619 CS_BIAS.n618 161.3
R277 CS_BIAS.n617 CS_BIAS.n475 161.3
R278 CS_BIAS.n616 CS_BIAS.n615 161.3
R279 CS_BIAS.n614 CS_BIAS.n476 161.3
R280 CS_BIAS.n613 CS_BIAS.n612 161.3
R281 CS_BIAS.n611 CS_BIAS.n477 161.3
R282 CS_BIAS.n610 CS_BIAS.n609 161.3
R283 CS_BIAS.n608 CS_BIAS.n478 161.3
R284 CS_BIAS.n607 CS_BIAS.n606 161.3
R285 CS_BIAS.n605 CS_BIAS.n479 161.3
R286 CS_BIAS.n604 CS_BIAS.n603 161.3
R287 CS_BIAS.n602 CS_BIAS.n480 161.3
R288 CS_BIAS.n601 CS_BIAS.n600 161.3
R289 CS_BIAS.n598 CS_BIAS.n481 161.3
R290 CS_BIAS.n597 CS_BIAS.n596 161.3
R291 CS_BIAS.n595 CS_BIAS.n482 161.3
R292 CS_BIAS.n594 CS_BIAS.n593 161.3
R293 CS_BIAS.n592 CS_BIAS.n483 161.3
R294 CS_BIAS.n591 CS_BIAS.n590 161.3
R295 CS_BIAS.n589 CS_BIAS.n484 161.3
R296 CS_BIAS.n588 CS_BIAS.n587 161.3
R297 CS_BIAS.n586 CS_BIAS.n485 161.3
R298 CS_BIAS.n585 CS_BIAS.n584 161.3
R299 CS_BIAS.n583 CS_BIAS.n582 161.3
R300 CS_BIAS.n581 CS_BIAS.n487 161.3
R301 CS_BIAS.n580 CS_BIAS.n579 161.3
R302 CS_BIAS.n578 CS_BIAS.n488 161.3
R303 CS_BIAS.n577 CS_BIAS.n576 161.3
R304 CS_BIAS.n575 CS_BIAS.n489 161.3
R305 CS_BIAS.n574 CS_BIAS.n573 161.3
R306 CS_BIAS.n572 CS_BIAS.n490 161.3
R307 CS_BIAS.n571 CS_BIAS.n570 161.3
R308 CS_BIAS.n569 CS_BIAS.n491 161.3
R309 CS_BIAS.n568 CS_BIAS.n567 161.3
R310 CS_BIAS.n566 CS_BIAS.n492 161.3
R311 CS_BIAS.n565 CS_BIAS.n564 161.3
R312 CS_BIAS.n562 CS_BIAS.n493 161.3
R313 CS_BIAS.n561 CS_BIAS.n560 161.3
R314 CS_BIAS.n559 CS_BIAS.n494 161.3
R315 CS_BIAS.n558 CS_BIAS.n557 161.3
R316 CS_BIAS.n556 CS_BIAS.n495 161.3
R317 CS_BIAS.n555 CS_BIAS.n554 161.3
R318 CS_BIAS.n553 CS_BIAS.n496 161.3
R319 CS_BIAS.n552 CS_BIAS.n551 161.3
R320 CS_BIAS.n550 CS_BIAS.n497 161.3
R321 CS_BIAS.n549 CS_BIAS.n548 161.3
R322 CS_BIAS.n547 CS_BIAS.n546 161.3
R323 CS_BIAS.n545 CS_BIAS.n499 161.3
R324 CS_BIAS.n544 CS_BIAS.n543 161.3
R325 CS_BIAS.n542 CS_BIAS.n500 161.3
R326 CS_BIAS.n541 CS_BIAS.n540 161.3
R327 CS_BIAS.n539 CS_BIAS.n501 161.3
R328 CS_BIAS.n538 CS_BIAS.n537 161.3
R329 CS_BIAS.n536 CS_BIAS.n502 161.3
R330 CS_BIAS.n535 CS_BIAS.n534 161.3
R331 CS_BIAS.n533 CS_BIAS.n503 161.3
R332 CS_BIAS.n532 CS_BIAS.n531 161.3
R333 CS_BIAS.n530 CS_BIAS.n504 161.3
R334 CS_BIAS.n529 CS_BIAS.n528 161.3
R335 CS_BIAS.n526 CS_BIAS.n505 161.3
R336 CS_BIAS.n525 CS_BIAS.n524 161.3
R337 CS_BIAS.n523 CS_BIAS.n506 161.3
R338 CS_BIAS.n522 CS_BIAS.n521 161.3
R339 CS_BIAS.n520 CS_BIAS.n507 161.3
R340 CS_BIAS.n519 CS_BIAS.n518 161.3
R341 CS_BIAS.n517 CS_BIAS.n508 161.3
R342 CS_BIAS.n516 CS_BIAS.n515 161.3
R343 CS_BIAS.n514 CS_BIAS.n509 161.3
R344 CS_BIAS.n513 CS_BIAS.n512 161.3
R345 CS_BIAS.n686 CS_BIAS.n685 161.3
R346 CS_BIAS.n684 CS_BIAS.n627 161.3
R347 CS_BIAS.n683 CS_BIAS.n682 161.3
R348 CS_BIAS.n681 CS_BIAS.n628 161.3
R349 CS_BIAS.n680 CS_BIAS.n679 161.3
R350 CS_BIAS.n678 CS_BIAS.n677 161.3
R351 CS_BIAS.n676 CS_BIAS.n630 161.3
R352 CS_BIAS.n675 CS_BIAS.n674 161.3
R353 CS_BIAS.n673 CS_BIAS.n631 161.3
R354 CS_BIAS.n672 CS_BIAS.n671 161.3
R355 CS_BIAS.n670 CS_BIAS.n632 161.3
R356 CS_BIAS.n669 CS_BIAS.n668 161.3
R357 CS_BIAS.n667 CS_BIAS.n633 161.3
R358 CS_BIAS.n666 CS_BIAS.n665 161.3
R359 CS_BIAS.n664 CS_BIAS.n634 161.3
R360 CS_BIAS.n663 CS_BIAS.n662 161.3
R361 CS_BIAS.n661 CS_BIAS.n635 161.3
R362 CS_BIAS.n660 CS_BIAS.n659 161.3
R363 CS_BIAS.n657 CS_BIAS.n636 161.3
R364 CS_BIAS.n656 CS_BIAS.n655 161.3
R365 CS_BIAS.n654 CS_BIAS.n637 161.3
R366 CS_BIAS.n653 CS_BIAS.n652 161.3
R367 CS_BIAS.n651 CS_BIAS.n638 161.3
R368 CS_BIAS.n650 CS_BIAS.n649 161.3
R369 CS_BIAS.n648 CS_BIAS.n639 161.3
R370 CS_BIAS.n647 CS_BIAS.n646 161.3
R371 CS_BIAS.n645 CS_BIAS.n640 161.3
R372 CS_BIAS.n644 CS_BIAS.n643 161.3
R373 CS_BIAS.n687 CS_BIAS.n626 161.3
R374 CS_BIAS.n750 CS_BIAS.n749 161.3
R375 CS_BIAS.n748 CS_BIAS.n451 161.3
R376 CS_BIAS.n747 CS_BIAS.n746 161.3
R377 CS_BIAS.n745 CS_BIAS.n452 161.3
R378 CS_BIAS.n744 CS_BIAS.n743 161.3
R379 CS_BIAS.n742 CS_BIAS.n453 161.3
R380 CS_BIAS.n741 CS_BIAS.n740 161.3
R381 CS_BIAS.n739 CS_BIAS.n454 161.3
R382 CS_BIAS.n738 CS_BIAS.n737 161.3
R383 CS_BIAS.n736 CS_BIAS.n455 161.3
R384 CS_BIAS.n735 CS_BIAS.n734 161.3
R385 CS_BIAS.n733 CS_BIAS.n456 161.3
R386 CS_BIAS.n732 CS_BIAS.n731 161.3
R387 CS_BIAS.n729 CS_BIAS.n457 161.3
R388 CS_BIAS.n728 CS_BIAS.n727 161.3
R389 CS_BIAS.n726 CS_BIAS.n458 161.3
R390 CS_BIAS.n725 CS_BIAS.n724 161.3
R391 CS_BIAS.n723 CS_BIAS.n459 161.3
R392 CS_BIAS.n722 CS_BIAS.n721 161.3
R393 CS_BIAS.n720 CS_BIAS.n460 161.3
R394 CS_BIAS.n719 CS_BIAS.n718 161.3
R395 CS_BIAS.n717 CS_BIAS.n461 161.3
R396 CS_BIAS.n716 CS_BIAS.n715 161.3
R397 CS_BIAS.n714 CS_BIAS.n713 161.3
R398 CS_BIAS.n712 CS_BIAS.n463 161.3
R399 CS_BIAS.n711 CS_BIAS.n710 161.3
R400 CS_BIAS.n709 CS_BIAS.n464 161.3
R401 CS_BIAS.n708 CS_BIAS.n707 161.3
R402 CS_BIAS.n706 CS_BIAS.n465 161.3
R403 CS_BIAS.n705 CS_BIAS.n704 161.3
R404 CS_BIAS.n703 CS_BIAS.n466 161.3
R405 CS_BIAS.n702 CS_BIAS.n701 161.3
R406 CS_BIAS.n700 CS_BIAS.n467 161.3
R407 CS_BIAS.n699 CS_BIAS.n698 161.3
R408 CS_BIAS.n697 CS_BIAS.n468 161.3
R409 CS_BIAS.n696 CS_BIAS.n695 161.3
R410 CS_BIAS.n693 CS_BIAS.n469 161.3
R411 CS_BIAS.n692 CS_BIAS.n691 161.3
R412 CS_BIAS.n690 CS_BIAS.n470 161.3
R413 CS_BIAS.n689 CS_BIAS.n688 161.3
R414 CS_BIAS.n176 CS_BIAS.n174 81.7203
R415 CS_BIAS.n473 CS_BIAS.n471 81.7203
R416 CS_BIAS.n176 CS_BIAS.n175 76.7376
R417 CS_BIAS.n173 CS_BIAS.n172 76.7376
R418 CS_BIAS.n171 CS_BIAS.n170 76.7376
R419 CS_BIAS.n622 CS_BIAS.n621 76.7376
R420 CS_BIAS.n624 CS_BIAS.n623 76.7376
R421 CS_BIAS.n473 CS_BIAS.n472 76.7376
R422 CS_BIAS.n448 CS_BIAS.n302 67.5631
R423 CS_BIAS.n169 CS_BIAS.n23 67.5631
R424 CS_BIAS.n301 CS_BIAS.n0 67.5631
R425 CS_BIAS.n898 CS_BIAS.n752 67.5631
R426 CS_BIAS.n620 CS_BIAS.n474 67.5631
R427 CS_BIAS.n751 CS_BIAS.n450 67.5631
R428 CS_BIAS.n369 CS_BIAS.n368 56.5193
R429 CS_BIAS.n404 CS_BIAS.n403 56.5193
R430 CS_BIAS.n125 CS_BIAS.n124 56.5193
R431 CS_BIAS.n90 CS_BIAS.n89 56.5193
R432 CS_BIAS.n257 CS_BIAS.n256 56.5193
R433 CS_BIAS.n222 CS_BIAS.n221 56.5193
R434 CS_BIAS.n817 CS_BIAS.n816 56.5193
R435 CS_BIAS.n853 CS_BIAS.n852 56.5193
R436 CS_BIAS.n539 CS_BIAS.n538 56.5193
R437 CS_BIAS.n575 CS_BIAS.n574 56.5193
R438 CS_BIAS.n706 CS_BIAS.n705 56.5193
R439 CS_BIAS.n670 CS_BIAS.n669 56.5193
R440 CS_BIAS.n439 CS_BIAS.n438 56.0336
R441 CS_BIAS.n160 CS_BIAS.n159 56.0336
R442 CS_BIAS.n292 CS_BIAS.n291 56.0336
R443 CS_BIAS.n889 CS_BIAS.n888 56.0336
R444 CS_BIAS.n611 CS_BIAS.n610 56.0336
R445 CS_BIAS.n742 CS_BIAS.n741 56.0336
R446 CS_BIAS.n63 CS_BIAS.n62 53.7369
R447 CS_BIAS.n195 CS_BIAS.n194 53.7369
R448 CS_BIAS.n789 CS_BIAS.n788 53.7369
R449 CS_BIAS.n511 CS_BIAS.n510 53.7369
R450 CS_BIAS.n642 CS_BIAS.n641 53.7369
R451 CS_BIAS.n342 CS_BIAS.n341 53.7369
R452 CS_BIAS.n789 CS_BIAS.t39 48.5439
R453 CS_BIAS.n511 CS_BIAS.t6 48.5439
R454 CS_BIAS.n642 CS_BIAS.t61 48.5439
R455 CS_BIAS.n342 CS_BIAS.t47 48.5439
R456 CS_BIAS.n63 CS_BIAS.t12 48.5438
R457 CS_BIAS.n195 CS_BIAS.t52 48.5438
R458 CS_BIAS.n351 CS_BIAS.n350 46.321
R459 CS_BIAS.n422 CS_BIAS.n421 46.321
R460 CS_BIAS.n143 CS_BIAS.n142 46.321
R461 CS_BIAS.n72 CS_BIAS.n71 46.321
R462 CS_BIAS.n275 CS_BIAS.n274 46.321
R463 CS_BIAS.n204 CS_BIAS.n203 46.321
R464 CS_BIAS.n798 CS_BIAS.n797 46.321
R465 CS_BIAS.n871 CS_BIAS.n870 46.321
R466 CS_BIAS.n520 CS_BIAS.n519 46.321
R467 CS_BIAS.n593 CS_BIAS.n592 46.321
R468 CS_BIAS.n724 CS_BIAS.n723 46.321
R469 CS_BIAS.n651 CS_BIAS.n650 46.321
R470 CS_BIAS.n386 CS_BIAS.n385 40.4934
R471 CS_BIAS.n387 CS_BIAS.n386 40.4934
R472 CS_BIAS.n108 CS_BIAS.n107 40.4934
R473 CS_BIAS.n107 CS_BIAS.n106 40.4934
R474 CS_BIAS.n240 CS_BIAS.n239 40.4934
R475 CS_BIAS.n239 CS_BIAS.n238 40.4934
R476 CS_BIAS.n834 CS_BIAS.n833 40.4934
R477 CS_BIAS.n835 CS_BIAS.n834 40.4934
R478 CS_BIAS.n556 CS_BIAS.n555 40.4934
R479 CS_BIAS.n557 CS_BIAS.n556 40.4934
R480 CS_BIAS.n688 CS_BIAS.n687 40.4934
R481 CS_BIAS.n687 CS_BIAS.n686 40.4934
R482 CS_BIAS.n352 CS_BIAS.n351 34.6658
R483 CS_BIAS.n421 CS_BIAS.n420 34.6658
R484 CS_BIAS.n142 CS_BIAS.n141 34.6658
R485 CS_BIAS.n73 CS_BIAS.n72 34.6658
R486 CS_BIAS.n274 CS_BIAS.n273 34.6658
R487 CS_BIAS.n205 CS_BIAS.n204 34.6658
R488 CS_BIAS.n799 CS_BIAS.n798 34.6658
R489 CS_BIAS.n870 CS_BIAS.n869 34.6658
R490 CS_BIAS.n521 CS_BIAS.n520 34.6658
R491 CS_BIAS.n592 CS_BIAS.n591 34.6658
R492 CS_BIAS.n723 CS_BIAS.n722 34.6658
R493 CS_BIAS.n652 CS_BIAS.n651 34.6658
R494 CS_BIAS.n440 CS_BIAS.n439 24.9531
R495 CS_BIAS.n161 CS_BIAS.n160 24.9531
R496 CS_BIAS.n293 CS_BIAS.n292 24.9531
R497 CS_BIAS.n890 CS_BIAS.n889 24.9531
R498 CS_BIAS.n612 CS_BIAS.n611 24.9531
R499 CS_BIAS.n743 CS_BIAS.n742 24.9531
R500 CS_BIAS.n350 CS_BIAS.n339 24.4675
R501 CS_BIAS.n346 CS_BIAS.n339 24.4675
R502 CS_BIAS.n346 CS_BIAS.n345 24.4675
R503 CS_BIAS.n345 CS_BIAS.n344 24.4675
R504 CS_BIAS.n368 CS_BIAS.n332 24.4675
R505 CS_BIAS.n364 CS_BIAS.n332 24.4675
R506 CS_BIAS.n364 CS_BIAS.n363 24.4675
R507 CS_BIAS.n363 CS_BIAS.n362 24.4675
R508 CS_BIAS.n362 CS_BIAS.n334 24.4675
R509 CS_BIAS.n358 CS_BIAS.n357 24.4675
R510 CS_BIAS.n357 CS_BIAS.n356 24.4675
R511 CS_BIAS.n356 CS_BIAS.n337 24.4675
R512 CS_BIAS.n352 CS_BIAS.n337 24.4675
R513 CS_BIAS.n385 CS_BIAS.n326 24.4675
R514 CS_BIAS.n381 CS_BIAS.n326 24.4675
R515 CS_BIAS.n381 CS_BIAS.n380 24.4675
R516 CS_BIAS.n380 CS_BIAS.n379 24.4675
R517 CS_BIAS.n376 CS_BIAS.n375 24.4675
R518 CS_BIAS.n375 CS_BIAS.n374 24.4675
R519 CS_BIAS.n374 CS_BIAS.n330 24.4675
R520 CS_BIAS.n370 CS_BIAS.n330 24.4675
R521 CS_BIAS.n370 CS_BIAS.n369 24.4675
R522 CS_BIAS.n403 CS_BIAS.n319 24.4675
R523 CS_BIAS.n399 CS_BIAS.n319 24.4675
R524 CS_BIAS.n399 CS_BIAS.n398 24.4675
R525 CS_BIAS.n398 CS_BIAS.n397 24.4675
R526 CS_BIAS.n397 CS_BIAS.n321 24.4675
R527 CS_BIAS.n393 CS_BIAS.n392 24.4675
R528 CS_BIAS.n392 CS_BIAS.n391 24.4675
R529 CS_BIAS.n391 CS_BIAS.n324 24.4675
R530 CS_BIAS.n387 CS_BIAS.n324 24.4675
R531 CS_BIAS.n420 CS_BIAS.n313 24.4675
R532 CS_BIAS.n416 CS_BIAS.n313 24.4675
R533 CS_BIAS.n416 CS_BIAS.n415 24.4675
R534 CS_BIAS.n415 CS_BIAS.n414 24.4675
R535 CS_BIAS.n411 CS_BIAS.n410 24.4675
R536 CS_BIAS.n410 CS_BIAS.n409 24.4675
R537 CS_BIAS.n409 CS_BIAS.n317 24.4675
R538 CS_BIAS.n405 CS_BIAS.n317 24.4675
R539 CS_BIAS.n405 CS_BIAS.n404 24.4675
R540 CS_BIAS.n438 CS_BIAS.n306 24.4675
R541 CS_BIAS.n434 CS_BIAS.n306 24.4675
R542 CS_BIAS.n434 CS_BIAS.n433 24.4675
R543 CS_BIAS.n433 CS_BIAS.n432 24.4675
R544 CS_BIAS.n432 CS_BIAS.n308 24.4675
R545 CS_BIAS.n428 CS_BIAS.n427 24.4675
R546 CS_BIAS.n427 CS_BIAS.n426 24.4675
R547 CS_BIAS.n426 CS_BIAS.n311 24.4675
R548 CS_BIAS.n422 CS_BIAS.n311 24.4675
R549 CS_BIAS.n446 CS_BIAS.n445 24.4675
R550 CS_BIAS.n445 CS_BIAS.n444 24.4675
R551 CS_BIAS.n444 CS_BIAS.n304 24.4675
R552 CS_BIAS.n440 CS_BIAS.n304 24.4675
R553 CS_BIAS.n167 CS_BIAS.n166 24.4675
R554 CS_BIAS.n166 CS_BIAS.n165 24.4675
R555 CS_BIAS.n165 CS_BIAS.n25 24.4675
R556 CS_BIAS.n161 CS_BIAS.n25 24.4675
R557 CS_BIAS.n159 CS_BIAS.n27 24.4675
R558 CS_BIAS.n155 CS_BIAS.n27 24.4675
R559 CS_BIAS.n155 CS_BIAS.n154 24.4675
R560 CS_BIAS.n154 CS_BIAS.n153 24.4675
R561 CS_BIAS.n153 CS_BIAS.n29 24.4675
R562 CS_BIAS.n149 CS_BIAS.n148 24.4675
R563 CS_BIAS.n148 CS_BIAS.n147 24.4675
R564 CS_BIAS.n147 CS_BIAS.n32 24.4675
R565 CS_BIAS.n143 CS_BIAS.n32 24.4675
R566 CS_BIAS.n141 CS_BIAS.n34 24.4675
R567 CS_BIAS.n137 CS_BIAS.n34 24.4675
R568 CS_BIAS.n137 CS_BIAS.n136 24.4675
R569 CS_BIAS.n136 CS_BIAS.n135 24.4675
R570 CS_BIAS.n132 CS_BIAS.n131 24.4675
R571 CS_BIAS.n131 CS_BIAS.n130 24.4675
R572 CS_BIAS.n130 CS_BIAS.n38 24.4675
R573 CS_BIAS.n126 CS_BIAS.n38 24.4675
R574 CS_BIAS.n126 CS_BIAS.n125 24.4675
R575 CS_BIAS.n124 CS_BIAS.n40 24.4675
R576 CS_BIAS.n120 CS_BIAS.n40 24.4675
R577 CS_BIAS.n120 CS_BIAS.n119 24.4675
R578 CS_BIAS.n119 CS_BIAS.n118 24.4675
R579 CS_BIAS.n118 CS_BIAS.n42 24.4675
R580 CS_BIAS.n114 CS_BIAS.n113 24.4675
R581 CS_BIAS.n113 CS_BIAS.n112 24.4675
R582 CS_BIAS.n112 CS_BIAS.n45 24.4675
R583 CS_BIAS.n108 CS_BIAS.n45 24.4675
R584 CS_BIAS.n106 CS_BIAS.n47 24.4675
R585 CS_BIAS.n102 CS_BIAS.n47 24.4675
R586 CS_BIAS.n102 CS_BIAS.n101 24.4675
R587 CS_BIAS.n101 CS_BIAS.n100 24.4675
R588 CS_BIAS.n97 CS_BIAS.n96 24.4675
R589 CS_BIAS.n96 CS_BIAS.n95 24.4675
R590 CS_BIAS.n95 CS_BIAS.n51 24.4675
R591 CS_BIAS.n91 CS_BIAS.n51 24.4675
R592 CS_BIAS.n91 CS_BIAS.n90 24.4675
R593 CS_BIAS.n89 CS_BIAS.n53 24.4675
R594 CS_BIAS.n85 CS_BIAS.n53 24.4675
R595 CS_BIAS.n85 CS_BIAS.n84 24.4675
R596 CS_BIAS.n84 CS_BIAS.n83 24.4675
R597 CS_BIAS.n83 CS_BIAS.n55 24.4675
R598 CS_BIAS.n79 CS_BIAS.n78 24.4675
R599 CS_BIAS.n78 CS_BIAS.n77 24.4675
R600 CS_BIAS.n77 CS_BIAS.n58 24.4675
R601 CS_BIAS.n73 CS_BIAS.n58 24.4675
R602 CS_BIAS.n71 CS_BIAS.n60 24.4675
R603 CS_BIAS.n67 CS_BIAS.n60 24.4675
R604 CS_BIAS.n67 CS_BIAS.n66 24.4675
R605 CS_BIAS.n66 CS_BIAS.n65 24.4675
R606 CS_BIAS.n299 CS_BIAS.n298 24.4675
R607 CS_BIAS.n298 CS_BIAS.n297 24.4675
R608 CS_BIAS.n297 CS_BIAS.n2 24.4675
R609 CS_BIAS.n293 CS_BIAS.n2 24.4675
R610 CS_BIAS.n291 CS_BIAS.n4 24.4675
R611 CS_BIAS.n287 CS_BIAS.n4 24.4675
R612 CS_BIAS.n287 CS_BIAS.n286 24.4675
R613 CS_BIAS.n286 CS_BIAS.n285 24.4675
R614 CS_BIAS.n285 CS_BIAS.n6 24.4675
R615 CS_BIAS.n281 CS_BIAS.n280 24.4675
R616 CS_BIAS.n280 CS_BIAS.n279 24.4675
R617 CS_BIAS.n279 CS_BIAS.n9 24.4675
R618 CS_BIAS.n275 CS_BIAS.n9 24.4675
R619 CS_BIAS.n273 CS_BIAS.n11 24.4675
R620 CS_BIAS.n269 CS_BIAS.n11 24.4675
R621 CS_BIAS.n269 CS_BIAS.n268 24.4675
R622 CS_BIAS.n268 CS_BIAS.n267 24.4675
R623 CS_BIAS.n264 CS_BIAS.n263 24.4675
R624 CS_BIAS.n263 CS_BIAS.n262 24.4675
R625 CS_BIAS.n262 CS_BIAS.n15 24.4675
R626 CS_BIAS.n258 CS_BIAS.n15 24.4675
R627 CS_BIAS.n258 CS_BIAS.n257 24.4675
R628 CS_BIAS.n256 CS_BIAS.n17 24.4675
R629 CS_BIAS.n252 CS_BIAS.n17 24.4675
R630 CS_BIAS.n252 CS_BIAS.n251 24.4675
R631 CS_BIAS.n251 CS_BIAS.n250 24.4675
R632 CS_BIAS.n250 CS_BIAS.n19 24.4675
R633 CS_BIAS.n246 CS_BIAS.n245 24.4675
R634 CS_BIAS.n245 CS_BIAS.n244 24.4675
R635 CS_BIAS.n244 CS_BIAS.n22 24.4675
R636 CS_BIAS.n240 CS_BIAS.n22 24.4675
R637 CS_BIAS.n238 CS_BIAS.n179 24.4675
R638 CS_BIAS.n234 CS_BIAS.n179 24.4675
R639 CS_BIAS.n234 CS_BIAS.n233 24.4675
R640 CS_BIAS.n233 CS_BIAS.n232 24.4675
R641 CS_BIAS.n229 CS_BIAS.n228 24.4675
R642 CS_BIAS.n228 CS_BIAS.n227 24.4675
R643 CS_BIAS.n227 CS_BIAS.n183 24.4675
R644 CS_BIAS.n223 CS_BIAS.n183 24.4675
R645 CS_BIAS.n223 CS_BIAS.n222 24.4675
R646 CS_BIAS.n221 CS_BIAS.n185 24.4675
R647 CS_BIAS.n217 CS_BIAS.n185 24.4675
R648 CS_BIAS.n217 CS_BIAS.n216 24.4675
R649 CS_BIAS.n216 CS_BIAS.n215 24.4675
R650 CS_BIAS.n215 CS_BIAS.n187 24.4675
R651 CS_BIAS.n211 CS_BIAS.n210 24.4675
R652 CS_BIAS.n210 CS_BIAS.n209 24.4675
R653 CS_BIAS.n209 CS_BIAS.n190 24.4675
R654 CS_BIAS.n205 CS_BIAS.n190 24.4675
R655 CS_BIAS.n203 CS_BIAS.n192 24.4675
R656 CS_BIAS.n199 CS_BIAS.n192 24.4675
R657 CS_BIAS.n199 CS_BIAS.n198 24.4675
R658 CS_BIAS.n198 CS_BIAS.n197 24.4675
R659 CS_BIAS.n792 CS_BIAS.n791 24.4675
R660 CS_BIAS.n793 CS_BIAS.n792 24.4675
R661 CS_BIAS.n793 CS_BIAS.n786 24.4675
R662 CS_BIAS.n797 CS_BIAS.n786 24.4675
R663 CS_BIAS.n799 CS_BIAS.n784 24.4675
R664 CS_BIAS.n803 CS_BIAS.n784 24.4675
R665 CS_BIAS.n804 CS_BIAS.n803 24.4675
R666 CS_BIAS.n806 CS_BIAS.n804 24.4675
R667 CS_BIAS.n810 CS_BIAS.n782 24.4675
R668 CS_BIAS.n811 CS_BIAS.n810 24.4675
R669 CS_BIAS.n812 CS_BIAS.n811 24.4675
R670 CS_BIAS.n812 CS_BIAS.n780 24.4675
R671 CS_BIAS.n816 CS_BIAS.n780 24.4675
R672 CS_BIAS.n818 CS_BIAS.n817 24.4675
R673 CS_BIAS.n818 CS_BIAS.n778 24.4675
R674 CS_BIAS.n822 CS_BIAS.n778 24.4675
R675 CS_BIAS.n823 CS_BIAS.n822 24.4675
R676 CS_BIAS.n824 CS_BIAS.n823 24.4675
R677 CS_BIAS.n828 CS_BIAS.n827 24.4675
R678 CS_BIAS.n829 CS_BIAS.n828 24.4675
R679 CS_BIAS.n829 CS_BIAS.n774 24.4675
R680 CS_BIAS.n833 CS_BIAS.n774 24.4675
R681 CS_BIAS.n835 CS_BIAS.n772 24.4675
R682 CS_BIAS.n839 CS_BIAS.n772 24.4675
R683 CS_BIAS.n840 CS_BIAS.n839 24.4675
R684 CS_BIAS.n842 CS_BIAS.n840 24.4675
R685 CS_BIAS.n846 CS_BIAS.n770 24.4675
R686 CS_BIAS.n847 CS_BIAS.n846 24.4675
R687 CS_BIAS.n848 CS_BIAS.n847 24.4675
R688 CS_BIAS.n848 CS_BIAS.n768 24.4675
R689 CS_BIAS.n852 CS_BIAS.n768 24.4675
R690 CS_BIAS.n854 CS_BIAS.n853 24.4675
R691 CS_BIAS.n854 CS_BIAS.n766 24.4675
R692 CS_BIAS.n858 CS_BIAS.n766 24.4675
R693 CS_BIAS.n859 CS_BIAS.n858 24.4675
R694 CS_BIAS.n860 CS_BIAS.n859 24.4675
R695 CS_BIAS.n864 CS_BIAS.n863 24.4675
R696 CS_BIAS.n865 CS_BIAS.n864 24.4675
R697 CS_BIAS.n865 CS_BIAS.n762 24.4675
R698 CS_BIAS.n869 CS_BIAS.n762 24.4675
R699 CS_BIAS.n871 CS_BIAS.n760 24.4675
R700 CS_BIAS.n875 CS_BIAS.n760 24.4675
R701 CS_BIAS.n876 CS_BIAS.n875 24.4675
R702 CS_BIAS.n878 CS_BIAS.n876 24.4675
R703 CS_BIAS.n882 CS_BIAS.n758 24.4675
R704 CS_BIAS.n883 CS_BIAS.n882 24.4675
R705 CS_BIAS.n884 CS_BIAS.n883 24.4675
R706 CS_BIAS.n884 CS_BIAS.n756 24.4675
R707 CS_BIAS.n888 CS_BIAS.n756 24.4675
R708 CS_BIAS.n890 CS_BIAS.n754 24.4675
R709 CS_BIAS.n894 CS_BIAS.n754 24.4675
R710 CS_BIAS.n895 CS_BIAS.n894 24.4675
R711 CS_BIAS.n896 CS_BIAS.n895 24.4675
R712 CS_BIAS.n514 CS_BIAS.n513 24.4675
R713 CS_BIAS.n515 CS_BIAS.n514 24.4675
R714 CS_BIAS.n515 CS_BIAS.n508 24.4675
R715 CS_BIAS.n519 CS_BIAS.n508 24.4675
R716 CS_BIAS.n521 CS_BIAS.n506 24.4675
R717 CS_BIAS.n525 CS_BIAS.n506 24.4675
R718 CS_BIAS.n526 CS_BIAS.n525 24.4675
R719 CS_BIAS.n528 CS_BIAS.n526 24.4675
R720 CS_BIAS.n532 CS_BIAS.n504 24.4675
R721 CS_BIAS.n533 CS_BIAS.n532 24.4675
R722 CS_BIAS.n534 CS_BIAS.n533 24.4675
R723 CS_BIAS.n534 CS_BIAS.n502 24.4675
R724 CS_BIAS.n538 CS_BIAS.n502 24.4675
R725 CS_BIAS.n540 CS_BIAS.n539 24.4675
R726 CS_BIAS.n540 CS_BIAS.n500 24.4675
R727 CS_BIAS.n544 CS_BIAS.n500 24.4675
R728 CS_BIAS.n545 CS_BIAS.n544 24.4675
R729 CS_BIAS.n546 CS_BIAS.n545 24.4675
R730 CS_BIAS.n550 CS_BIAS.n549 24.4675
R731 CS_BIAS.n551 CS_BIAS.n550 24.4675
R732 CS_BIAS.n551 CS_BIAS.n496 24.4675
R733 CS_BIAS.n555 CS_BIAS.n496 24.4675
R734 CS_BIAS.n557 CS_BIAS.n494 24.4675
R735 CS_BIAS.n561 CS_BIAS.n494 24.4675
R736 CS_BIAS.n562 CS_BIAS.n561 24.4675
R737 CS_BIAS.n564 CS_BIAS.n562 24.4675
R738 CS_BIAS.n568 CS_BIAS.n492 24.4675
R739 CS_BIAS.n569 CS_BIAS.n568 24.4675
R740 CS_BIAS.n570 CS_BIAS.n569 24.4675
R741 CS_BIAS.n570 CS_BIAS.n490 24.4675
R742 CS_BIAS.n574 CS_BIAS.n490 24.4675
R743 CS_BIAS.n576 CS_BIAS.n575 24.4675
R744 CS_BIAS.n576 CS_BIAS.n488 24.4675
R745 CS_BIAS.n580 CS_BIAS.n488 24.4675
R746 CS_BIAS.n581 CS_BIAS.n580 24.4675
R747 CS_BIAS.n582 CS_BIAS.n581 24.4675
R748 CS_BIAS.n586 CS_BIAS.n585 24.4675
R749 CS_BIAS.n587 CS_BIAS.n586 24.4675
R750 CS_BIAS.n587 CS_BIAS.n484 24.4675
R751 CS_BIAS.n591 CS_BIAS.n484 24.4675
R752 CS_BIAS.n593 CS_BIAS.n482 24.4675
R753 CS_BIAS.n597 CS_BIAS.n482 24.4675
R754 CS_BIAS.n598 CS_BIAS.n597 24.4675
R755 CS_BIAS.n600 CS_BIAS.n598 24.4675
R756 CS_BIAS.n604 CS_BIAS.n480 24.4675
R757 CS_BIAS.n605 CS_BIAS.n604 24.4675
R758 CS_BIAS.n606 CS_BIAS.n605 24.4675
R759 CS_BIAS.n606 CS_BIAS.n478 24.4675
R760 CS_BIAS.n610 CS_BIAS.n478 24.4675
R761 CS_BIAS.n612 CS_BIAS.n476 24.4675
R762 CS_BIAS.n616 CS_BIAS.n476 24.4675
R763 CS_BIAS.n617 CS_BIAS.n616 24.4675
R764 CS_BIAS.n618 CS_BIAS.n617 24.4675
R765 CS_BIAS.n743 CS_BIAS.n452 24.4675
R766 CS_BIAS.n747 CS_BIAS.n452 24.4675
R767 CS_BIAS.n748 CS_BIAS.n747 24.4675
R768 CS_BIAS.n749 CS_BIAS.n748 24.4675
R769 CS_BIAS.n724 CS_BIAS.n458 24.4675
R770 CS_BIAS.n728 CS_BIAS.n458 24.4675
R771 CS_BIAS.n729 CS_BIAS.n728 24.4675
R772 CS_BIAS.n731 CS_BIAS.n729 24.4675
R773 CS_BIAS.n735 CS_BIAS.n456 24.4675
R774 CS_BIAS.n736 CS_BIAS.n735 24.4675
R775 CS_BIAS.n737 CS_BIAS.n736 24.4675
R776 CS_BIAS.n737 CS_BIAS.n454 24.4675
R777 CS_BIAS.n741 CS_BIAS.n454 24.4675
R778 CS_BIAS.n707 CS_BIAS.n706 24.4675
R779 CS_BIAS.n707 CS_BIAS.n464 24.4675
R780 CS_BIAS.n711 CS_BIAS.n464 24.4675
R781 CS_BIAS.n712 CS_BIAS.n711 24.4675
R782 CS_BIAS.n713 CS_BIAS.n712 24.4675
R783 CS_BIAS.n717 CS_BIAS.n716 24.4675
R784 CS_BIAS.n718 CS_BIAS.n717 24.4675
R785 CS_BIAS.n718 CS_BIAS.n460 24.4675
R786 CS_BIAS.n722 CS_BIAS.n460 24.4675
R787 CS_BIAS.n688 CS_BIAS.n470 24.4675
R788 CS_BIAS.n692 CS_BIAS.n470 24.4675
R789 CS_BIAS.n693 CS_BIAS.n692 24.4675
R790 CS_BIAS.n695 CS_BIAS.n693 24.4675
R791 CS_BIAS.n699 CS_BIAS.n468 24.4675
R792 CS_BIAS.n700 CS_BIAS.n699 24.4675
R793 CS_BIAS.n701 CS_BIAS.n700 24.4675
R794 CS_BIAS.n701 CS_BIAS.n466 24.4675
R795 CS_BIAS.n705 CS_BIAS.n466 24.4675
R796 CS_BIAS.n645 CS_BIAS.n644 24.4675
R797 CS_BIAS.n646 CS_BIAS.n645 24.4675
R798 CS_BIAS.n646 CS_BIAS.n639 24.4675
R799 CS_BIAS.n650 CS_BIAS.n639 24.4675
R800 CS_BIAS.n652 CS_BIAS.n637 24.4675
R801 CS_BIAS.n656 CS_BIAS.n637 24.4675
R802 CS_BIAS.n657 CS_BIAS.n656 24.4675
R803 CS_BIAS.n659 CS_BIAS.n657 24.4675
R804 CS_BIAS.n663 CS_BIAS.n635 24.4675
R805 CS_BIAS.n664 CS_BIAS.n663 24.4675
R806 CS_BIAS.n665 CS_BIAS.n664 24.4675
R807 CS_BIAS.n665 CS_BIAS.n633 24.4675
R808 CS_BIAS.n669 CS_BIAS.n633 24.4675
R809 CS_BIAS.n671 CS_BIAS.n670 24.4675
R810 CS_BIAS.n671 CS_BIAS.n631 24.4675
R811 CS_BIAS.n675 CS_BIAS.n631 24.4675
R812 CS_BIAS.n676 CS_BIAS.n675 24.4675
R813 CS_BIAS.n677 CS_BIAS.n676 24.4675
R814 CS_BIAS.n681 CS_BIAS.n680 24.4675
R815 CS_BIAS.n682 CS_BIAS.n681 24.4675
R816 CS_BIAS.n682 CS_BIAS.n627 24.4675
R817 CS_BIAS.n686 CS_BIAS.n627 24.4675
R818 CS_BIAS.n344 CS_BIAS.n341 22.0208
R819 CS_BIAS.n428 CS_BIAS.n310 22.0208
R820 CS_BIAS.n149 CS_BIAS.n31 22.0208
R821 CS_BIAS.n65 CS_BIAS.n62 22.0208
R822 CS_BIAS.n281 CS_BIAS.n8 22.0208
R823 CS_BIAS.n197 CS_BIAS.n194 22.0208
R824 CS_BIAS.n791 CS_BIAS.n788 22.0208
R825 CS_BIAS.n878 CS_BIAS.n877 22.0208
R826 CS_BIAS.n513 CS_BIAS.n510 22.0208
R827 CS_BIAS.n600 CS_BIAS.n599 22.0208
R828 CS_BIAS.n731 CS_BIAS.n730 22.0208
R829 CS_BIAS.n644 CS_BIAS.n641 22.0208
R830 CS_BIAS.n379 CS_BIAS.n328 19.0848
R831 CS_BIAS.n393 CS_BIAS.n323 19.0848
R832 CS_BIAS.n114 CS_BIAS.n44 19.0848
R833 CS_BIAS.n100 CS_BIAS.n49 19.0848
R834 CS_BIAS.n246 CS_BIAS.n21 19.0848
R835 CS_BIAS.n232 CS_BIAS.n181 19.0848
R836 CS_BIAS.n827 CS_BIAS.n776 19.0848
R837 CS_BIAS.n842 CS_BIAS.n841 19.0848
R838 CS_BIAS.n549 CS_BIAS.n498 19.0848
R839 CS_BIAS.n564 CS_BIAS.n563 19.0848
R840 CS_BIAS.n695 CS_BIAS.n694 19.0848
R841 CS_BIAS.n680 CS_BIAS.n629 19.0848
R842 CS_BIAS.n358 CS_BIAS.n336 16.1487
R843 CS_BIAS.n414 CS_BIAS.n315 16.1487
R844 CS_BIAS.n135 CS_BIAS.n36 16.1487
R845 CS_BIAS.n79 CS_BIAS.n57 16.1487
R846 CS_BIAS.n267 CS_BIAS.n13 16.1487
R847 CS_BIAS.n211 CS_BIAS.n189 16.1487
R848 CS_BIAS.n806 CS_BIAS.n805 16.1487
R849 CS_BIAS.n863 CS_BIAS.n764 16.1487
R850 CS_BIAS.n528 CS_BIAS.n527 16.1487
R851 CS_BIAS.n585 CS_BIAS.n486 16.1487
R852 CS_BIAS.n716 CS_BIAS.n462 16.1487
R853 CS_BIAS.n659 CS_BIAS.n658 16.1487
R854 CS_BIAS.n341 CS_BIAS.t40 14.9027
R855 CS_BIAS.n336 CS_BIAS.t57 14.9027
R856 CS_BIAS.n328 CS_BIAS.t49 14.9027
R857 CS_BIAS.n323 CS_BIAS.t33 14.9027
R858 CS_BIAS.n315 CS_BIAS.t59 14.9027
R859 CS_BIAS.n310 CS_BIAS.t44 14.9027
R860 CS_BIAS.n302 CS_BIAS.t35 14.9027
R861 CS_BIAS.n23 CS_BIAS.t20 14.9027
R862 CS_BIAS.n31 CS_BIAS.t14 14.9027
R863 CS_BIAS.n36 CS_BIAS.t16 14.9027
R864 CS_BIAS.n44 CS_BIAS.t2 14.9027
R865 CS_BIAS.n49 CS_BIAS.t8 14.9027
R866 CS_BIAS.n57 CS_BIAS.t22 14.9027
R867 CS_BIAS.n62 CS_BIAS.t24 14.9027
R868 CS_BIAS.n0 CS_BIAS.t51 14.9027
R869 CS_BIAS.n8 CS_BIAS.t48 14.9027
R870 CS_BIAS.n13 CS_BIAS.t38 14.9027
R871 CS_BIAS.n21 CS_BIAS.t58 14.9027
R872 CS_BIAS.n181 CS_BIAS.t46 14.9027
R873 CS_BIAS.n189 CS_BIAS.t34 14.9027
R874 CS_BIAS.n194 CS_BIAS.t54 14.9027
R875 CS_BIAS.n788 CS_BIAS.t55 14.9027
R876 CS_BIAS.n805 CS_BIAS.t41 14.9027
R877 CS_BIAS.n776 CS_BIAS.t63 14.9027
R878 CS_BIAS.n841 CS_BIAS.t50 14.9027
R879 CS_BIAS.n764 CS_BIAS.t42 14.9027
R880 CS_BIAS.n877 CS_BIAS.t37 14.9027
R881 CS_BIAS.n752 CS_BIAS.t60 14.9027
R882 CS_BIAS.n510 CS_BIAS.t4 14.9027
R883 CS_BIAS.n527 CS_BIAS.t0 14.9027
R884 CS_BIAS.n498 CS_BIAS.t30 14.9027
R885 CS_BIAS.n563 CS_BIAS.t28 14.9027
R886 CS_BIAS.n486 CS_BIAS.t10 14.9027
R887 CS_BIAS.n599 CS_BIAS.t26 14.9027
R888 CS_BIAS.n474 CS_BIAS.t18 14.9027
R889 CS_BIAS.n450 CS_BIAS.t36 14.9027
R890 CS_BIAS.n730 CS_BIAS.t62 14.9027
R891 CS_BIAS.n462 CS_BIAS.t56 14.9027
R892 CS_BIAS.n694 CS_BIAS.t45 14.9027
R893 CS_BIAS.n641 CS_BIAS.t43 14.9027
R894 CS_BIAS.n658 CS_BIAS.t53 14.9027
R895 CS_BIAS.n629 CS_BIAS.t32 14.9027
R896 CS_BIAS.n171 CS_BIAS.n169 14.6207
R897 CS_BIAS.n622 CS_BIAS.n620 14.6207
R898 CS_BIAS.n900 CS_BIAS.n449 11.3713
R899 CS_BIAS.n446 CS_BIAS.n302 11.2553
R900 CS_BIAS.n167 CS_BIAS.n23 11.2553
R901 CS_BIAS.n299 CS_BIAS.n0 11.2553
R902 CS_BIAS.n896 CS_BIAS.n752 11.2553
R903 CS_BIAS.n618 CS_BIAS.n474 11.2553
R904 CS_BIAS.n749 CS_BIAS.n450 11.2553
R905 CS_BIAS.n178 CS_BIAS.n177 9.50425
R906 CS_BIAS.n626 CS_BIAS.n625 9.50425
R907 CS_BIAS.n900 CS_BIAS.n899 8.93891
R908 CS_BIAS.n336 CS_BIAS.n334 8.31928
R909 CS_BIAS.n411 CS_BIAS.n315 8.31928
R910 CS_BIAS.n132 CS_BIAS.n36 8.31928
R911 CS_BIAS.n57 CS_BIAS.n55 8.31928
R912 CS_BIAS.n264 CS_BIAS.n13 8.31928
R913 CS_BIAS.n189 CS_BIAS.n187 8.31928
R914 CS_BIAS.n805 CS_BIAS.n782 8.31928
R915 CS_BIAS.n860 CS_BIAS.n764 8.31928
R916 CS_BIAS.n527 CS_BIAS.n504 8.31928
R917 CS_BIAS.n582 CS_BIAS.n486 8.31928
R918 CS_BIAS.n713 CS_BIAS.n462 8.31928
R919 CS_BIAS.n658 CS_BIAS.n635 8.31928
R920 CS_BIAS.n449 CS_BIAS.n301 7.54478
R921 CS_BIAS.n899 CS_BIAS.n751 7.54478
R922 CS_BIAS.n174 CS_BIAS.t25 5.87587
R923 CS_BIAS.n174 CS_BIAS.t13 5.87587
R924 CS_BIAS.n175 CS_BIAS.t9 5.87587
R925 CS_BIAS.n175 CS_BIAS.t23 5.87587
R926 CS_BIAS.n172 CS_BIAS.t17 5.87587
R927 CS_BIAS.n172 CS_BIAS.t3 5.87587
R928 CS_BIAS.n170 CS_BIAS.t21 5.87587
R929 CS_BIAS.n170 CS_BIAS.t15 5.87587
R930 CS_BIAS.n621 CS_BIAS.t27 5.87587
R931 CS_BIAS.n621 CS_BIAS.t19 5.87587
R932 CS_BIAS.n623 CS_BIAS.t29 5.87587
R933 CS_BIAS.n623 CS_BIAS.t11 5.87587
R934 CS_BIAS.n472 CS_BIAS.t1 5.87587
R935 CS_BIAS.n472 CS_BIAS.t31 5.87587
R936 CS_BIAS.n471 CS_BIAS.t7 5.87587
R937 CS_BIAS.n471 CS_BIAS.t5 5.87587
R938 CS_BIAS.n449 CS_BIAS.n448 5.4463
R939 CS_BIAS.n899 CS_BIAS.n898 5.4463
R940 CS_BIAS.n376 CS_BIAS.n328 5.38324
R941 CS_BIAS.n323 CS_BIAS.n321 5.38324
R942 CS_BIAS.n44 CS_BIAS.n42 5.38324
R943 CS_BIAS.n97 CS_BIAS.n49 5.38324
R944 CS_BIAS.n21 CS_BIAS.n19 5.38324
R945 CS_BIAS.n229 CS_BIAS.n181 5.38324
R946 CS_BIAS.n824 CS_BIAS.n776 5.38324
R947 CS_BIAS.n841 CS_BIAS.n770 5.38324
R948 CS_BIAS.n546 CS_BIAS.n498 5.38324
R949 CS_BIAS.n563 CS_BIAS.n492 5.38324
R950 CS_BIAS.n694 CS_BIAS.n468 5.38324
R951 CS_BIAS.n677 CS_BIAS.n629 5.38324
R952 CS_BIAS.n173 CS_BIAS.n171 4.98326
R953 CS_BIAS.n624 CS_BIAS.n622 4.98326
R954 CS_BIAS CS_BIAS.n900 4.69423
R955 CS_BIAS.n177 CS_BIAS.n176 2.46171
R956 CS_BIAS.n177 CS_BIAS.n173 2.46171
R957 CS_BIAS.n625 CS_BIAS.n624 2.46171
R958 CS_BIAS.n625 CS_BIAS.n473 2.46171
R959 CS_BIAS.n310 CS_BIAS.n308 2.4472
R960 CS_BIAS.n31 CS_BIAS.n29 2.4472
R961 CS_BIAS.n8 CS_BIAS.n6 2.4472
R962 CS_BIAS.n877 CS_BIAS.n758 2.4472
R963 CS_BIAS.n599 CS_BIAS.n480 2.4472
R964 CS_BIAS.n730 CS_BIAS.n456 2.4472
R965 CS_BIAS.n343 CS_BIAS.n342 1.07289
R966 CS_BIAS.n790 CS_BIAS.n789 1.07289
R967 CS_BIAS.n512 CS_BIAS.n511 1.07289
R968 CS_BIAS.n643 CS_BIAS.n642 1.07289
R969 CS_BIAS.n64 CS_BIAS.n63 1.07289
R970 CS_BIAS.n196 CS_BIAS.n195 1.07289
R971 CS_BIAS.n448 CS_BIAS.n447 0.466196
R972 CS_BIAS.n169 CS_BIAS.n168 0.466196
R973 CS_BIAS.n301 CS_BIAS.n300 0.466196
R974 CS_BIAS.n898 CS_BIAS.n897 0.466196
R975 CS_BIAS.n620 CS_BIAS.n619 0.466196
R976 CS_BIAS.n751 CS_BIAS.n750 0.466196
R977 CS_BIAS.n447 CS_BIAS.n303 0.189894
R978 CS_BIAS.n443 CS_BIAS.n303 0.189894
R979 CS_BIAS.n443 CS_BIAS.n442 0.189894
R980 CS_BIAS.n442 CS_BIAS.n441 0.189894
R981 CS_BIAS.n441 CS_BIAS.n305 0.189894
R982 CS_BIAS.n437 CS_BIAS.n305 0.189894
R983 CS_BIAS.n437 CS_BIAS.n436 0.189894
R984 CS_BIAS.n436 CS_BIAS.n435 0.189894
R985 CS_BIAS.n435 CS_BIAS.n307 0.189894
R986 CS_BIAS.n431 CS_BIAS.n307 0.189894
R987 CS_BIAS.n431 CS_BIAS.n430 0.189894
R988 CS_BIAS.n430 CS_BIAS.n429 0.189894
R989 CS_BIAS.n429 CS_BIAS.n309 0.189894
R990 CS_BIAS.n425 CS_BIAS.n309 0.189894
R991 CS_BIAS.n425 CS_BIAS.n424 0.189894
R992 CS_BIAS.n424 CS_BIAS.n423 0.189894
R993 CS_BIAS.n423 CS_BIAS.n312 0.189894
R994 CS_BIAS.n419 CS_BIAS.n312 0.189894
R995 CS_BIAS.n419 CS_BIAS.n418 0.189894
R996 CS_BIAS.n418 CS_BIAS.n417 0.189894
R997 CS_BIAS.n417 CS_BIAS.n314 0.189894
R998 CS_BIAS.n413 CS_BIAS.n314 0.189894
R999 CS_BIAS.n413 CS_BIAS.n412 0.189894
R1000 CS_BIAS.n412 CS_BIAS.n316 0.189894
R1001 CS_BIAS.n408 CS_BIAS.n316 0.189894
R1002 CS_BIAS.n408 CS_BIAS.n407 0.189894
R1003 CS_BIAS.n407 CS_BIAS.n406 0.189894
R1004 CS_BIAS.n406 CS_BIAS.n318 0.189894
R1005 CS_BIAS.n402 CS_BIAS.n318 0.189894
R1006 CS_BIAS.n402 CS_BIAS.n401 0.189894
R1007 CS_BIAS.n401 CS_BIAS.n400 0.189894
R1008 CS_BIAS.n400 CS_BIAS.n320 0.189894
R1009 CS_BIAS.n396 CS_BIAS.n320 0.189894
R1010 CS_BIAS.n396 CS_BIAS.n395 0.189894
R1011 CS_BIAS.n395 CS_BIAS.n394 0.189894
R1012 CS_BIAS.n394 CS_BIAS.n322 0.189894
R1013 CS_BIAS.n390 CS_BIAS.n322 0.189894
R1014 CS_BIAS.n390 CS_BIAS.n389 0.189894
R1015 CS_BIAS.n389 CS_BIAS.n388 0.189894
R1016 CS_BIAS.n388 CS_BIAS.n325 0.189894
R1017 CS_BIAS.n384 CS_BIAS.n325 0.189894
R1018 CS_BIAS.n384 CS_BIAS.n383 0.189894
R1019 CS_BIAS.n383 CS_BIAS.n382 0.189894
R1020 CS_BIAS.n382 CS_BIAS.n327 0.189894
R1021 CS_BIAS.n378 CS_BIAS.n327 0.189894
R1022 CS_BIAS.n378 CS_BIAS.n377 0.189894
R1023 CS_BIAS.n377 CS_BIAS.n329 0.189894
R1024 CS_BIAS.n373 CS_BIAS.n329 0.189894
R1025 CS_BIAS.n373 CS_BIAS.n372 0.189894
R1026 CS_BIAS.n372 CS_BIAS.n371 0.189894
R1027 CS_BIAS.n371 CS_BIAS.n331 0.189894
R1028 CS_BIAS.n367 CS_BIAS.n331 0.189894
R1029 CS_BIAS.n367 CS_BIAS.n366 0.189894
R1030 CS_BIAS.n366 CS_BIAS.n365 0.189894
R1031 CS_BIAS.n365 CS_BIAS.n333 0.189894
R1032 CS_BIAS.n361 CS_BIAS.n333 0.189894
R1033 CS_BIAS.n361 CS_BIAS.n360 0.189894
R1034 CS_BIAS.n360 CS_BIAS.n359 0.189894
R1035 CS_BIAS.n359 CS_BIAS.n335 0.189894
R1036 CS_BIAS.n355 CS_BIAS.n335 0.189894
R1037 CS_BIAS.n355 CS_BIAS.n354 0.189894
R1038 CS_BIAS.n354 CS_BIAS.n353 0.189894
R1039 CS_BIAS.n353 CS_BIAS.n338 0.189894
R1040 CS_BIAS.n349 CS_BIAS.n338 0.189894
R1041 CS_BIAS.n349 CS_BIAS.n348 0.189894
R1042 CS_BIAS.n348 CS_BIAS.n347 0.189894
R1043 CS_BIAS.n347 CS_BIAS.n340 0.189894
R1044 CS_BIAS.n343 CS_BIAS.n340 0.189894
R1045 CS_BIAS.n168 CS_BIAS.n24 0.189894
R1046 CS_BIAS.n164 CS_BIAS.n24 0.189894
R1047 CS_BIAS.n164 CS_BIAS.n163 0.189894
R1048 CS_BIAS.n163 CS_BIAS.n162 0.189894
R1049 CS_BIAS.n162 CS_BIAS.n26 0.189894
R1050 CS_BIAS.n158 CS_BIAS.n26 0.189894
R1051 CS_BIAS.n158 CS_BIAS.n157 0.189894
R1052 CS_BIAS.n157 CS_BIAS.n156 0.189894
R1053 CS_BIAS.n156 CS_BIAS.n28 0.189894
R1054 CS_BIAS.n152 CS_BIAS.n28 0.189894
R1055 CS_BIAS.n152 CS_BIAS.n151 0.189894
R1056 CS_BIAS.n151 CS_BIAS.n150 0.189894
R1057 CS_BIAS.n150 CS_BIAS.n30 0.189894
R1058 CS_BIAS.n146 CS_BIAS.n30 0.189894
R1059 CS_BIAS.n146 CS_BIAS.n145 0.189894
R1060 CS_BIAS.n145 CS_BIAS.n144 0.189894
R1061 CS_BIAS.n144 CS_BIAS.n33 0.189894
R1062 CS_BIAS.n140 CS_BIAS.n33 0.189894
R1063 CS_BIAS.n140 CS_BIAS.n139 0.189894
R1064 CS_BIAS.n139 CS_BIAS.n138 0.189894
R1065 CS_BIAS.n138 CS_BIAS.n35 0.189894
R1066 CS_BIAS.n134 CS_BIAS.n35 0.189894
R1067 CS_BIAS.n134 CS_BIAS.n133 0.189894
R1068 CS_BIAS.n133 CS_BIAS.n37 0.189894
R1069 CS_BIAS.n129 CS_BIAS.n37 0.189894
R1070 CS_BIAS.n129 CS_BIAS.n128 0.189894
R1071 CS_BIAS.n128 CS_BIAS.n127 0.189894
R1072 CS_BIAS.n127 CS_BIAS.n39 0.189894
R1073 CS_BIAS.n123 CS_BIAS.n39 0.189894
R1074 CS_BIAS.n123 CS_BIAS.n122 0.189894
R1075 CS_BIAS.n122 CS_BIAS.n121 0.189894
R1076 CS_BIAS.n121 CS_BIAS.n41 0.189894
R1077 CS_BIAS.n117 CS_BIAS.n41 0.189894
R1078 CS_BIAS.n117 CS_BIAS.n116 0.189894
R1079 CS_BIAS.n116 CS_BIAS.n115 0.189894
R1080 CS_BIAS.n115 CS_BIAS.n43 0.189894
R1081 CS_BIAS.n111 CS_BIAS.n43 0.189894
R1082 CS_BIAS.n111 CS_BIAS.n110 0.189894
R1083 CS_BIAS.n110 CS_BIAS.n109 0.189894
R1084 CS_BIAS.n109 CS_BIAS.n46 0.189894
R1085 CS_BIAS.n105 CS_BIAS.n46 0.189894
R1086 CS_BIAS.n105 CS_BIAS.n104 0.189894
R1087 CS_BIAS.n104 CS_BIAS.n103 0.189894
R1088 CS_BIAS.n103 CS_BIAS.n48 0.189894
R1089 CS_BIAS.n99 CS_BIAS.n48 0.189894
R1090 CS_BIAS.n99 CS_BIAS.n98 0.189894
R1091 CS_BIAS.n98 CS_BIAS.n50 0.189894
R1092 CS_BIAS.n94 CS_BIAS.n50 0.189894
R1093 CS_BIAS.n94 CS_BIAS.n93 0.189894
R1094 CS_BIAS.n93 CS_BIAS.n92 0.189894
R1095 CS_BIAS.n92 CS_BIAS.n52 0.189894
R1096 CS_BIAS.n88 CS_BIAS.n52 0.189894
R1097 CS_BIAS.n88 CS_BIAS.n87 0.189894
R1098 CS_BIAS.n87 CS_BIAS.n86 0.189894
R1099 CS_BIAS.n86 CS_BIAS.n54 0.189894
R1100 CS_BIAS.n82 CS_BIAS.n54 0.189894
R1101 CS_BIAS.n82 CS_BIAS.n81 0.189894
R1102 CS_BIAS.n81 CS_BIAS.n80 0.189894
R1103 CS_BIAS.n80 CS_BIAS.n56 0.189894
R1104 CS_BIAS.n76 CS_BIAS.n56 0.189894
R1105 CS_BIAS.n76 CS_BIAS.n75 0.189894
R1106 CS_BIAS.n75 CS_BIAS.n74 0.189894
R1107 CS_BIAS.n74 CS_BIAS.n59 0.189894
R1108 CS_BIAS.n70 CS_BIAS.n59 0.189894
R1109 CS_BIAS.n70 CS_BIAS.n69 0.189894
R1110 CS_BIAS.n69 CS_BIAS.n68 0.189894
R1111 CS_BIAS.n68 CS_BIAS.n61 0.189894
R1112 CS_BIAS.n64 CS_BIAS.n61 0.189894
R1113 CS_BIAS.n237 CS_BIAS.n236 0.189894
R1114 CS_BIAS.n236 CS_BIAS.n235 0.189894
R1115 CS_BIAS.n235 CS_BIAS.n180 0.189894
R1116 CS_BIAS.n231 CS_BIAS.n180 0.189894
R1117 CS_BIAS.n231 CS_BIAS.n230 0.189894
R1118 CS_BIAS.n230 CS_BIAS.n182 0.189894
R1119 CS_BIAS.n226 CS_BIAS.n182 0.189894
R1120 CS_BIAS.n226 CS_BIAS.n225 0.189894
R1121 CS_BIAS.n225 CS_BIAS.n224 0.189894
R1122 CS_BIAS.n224 CS_BIAS.n184 0.189894
R1123 CS_BIAS.n220 CS_BIAS.n184 0.189894
R1124 CS_BIAS.n220 CS_BIAS.n219 0.189894
R1125 CS_BIAS.n219 CS_BIAS.n218 0.189894
R1126 CS_BIAS.n218 CS_BIAS.n186 0.189894
R1127 CS_BIAS.n214 CS_BIAS.n186 0.189894
R1128 CS_BIAS.n214 CS_BIAS.n213 0.189894
R1129 CS_BIAS.n213 CS_BIAS.n212 0.189894
R1130 CS_BIAS.n212 CS_BIAS.n188 0.189894
R1131 CS_BIAS.n208 CS_BIAS.n188 0.189894
R1132 CS_BIAS.n208 CS_BIAS.n207 0.189894
R1133 CS_BIAS.n207 CS_BIAS.n206 0.189894
R1134 CS_BIAS.n206 CS_BIAS.n191 0.189894
R1135 CS_BIAS.n202 CS_BIAS.n191 0.189894
R1136 CS_BIAS.n202 CS_BIAS.n201 0.189894
R1137 CS_BIAS.n201 CS_BIAS.n200 0.189894
R1138 CS_BIAS.n200 CS_BIAS.n193 0.189894
R1139 CS_BIAS.n196 CS_BIAS.n193 0.189894
R1140 CS_BIAS.n300 CS_BIAS.n1 0.189894
R1141 CS_BIAS.n296 CS_BIAS.n1 0.189894
R1142 CS_BIAS.n296 CS_BIAS.n295 0.189894
R1143 CS_BIAS.n295 CS_BIAS.n294 0.189894
R1144 CS_BIAS.n294 CS_BIAS.n3 0.189894
R1145 CS_BIAS.n290 CS_BIAS.n3 0.189894
R1146 CS_BIAS.n290 CS_BIAS.n289 0.189894
R1147 CS_BIAS.n289 CS_BIAS.n288 0.189894
R1148 CS_BIAS.n288 CS_BIAS.n5 0.189894
R1149 CS_BIAS.n284 CS_BIAS.n5 0.189894
R1150 CS_BIAS.n284 CS_BIAS.n283 0.189894
R1151 CS_BIAS.n283 CS_BIAS.n282 0.189894
R1152 CS_BIAS.n282 CS_BIAS.n7 0.189894
R1153 CS_BIAS.n278 CS_BIAS.n7 0.189894
R1154 CS_BIAS.n278 CS_BIAS.n277 0.189894
R1155 CS_BIAS.n277 CS_BIAS.n276 0.189894
R1156 CS_BIAS.n276 CS_BIAS.n10 0.189894
R1157 CS_BIAS.n272 CS_BIAS.n10 0.189894
R1158 CS_BIAS.n272 CS_BIAS.n271 0.189894
R1159 CS_BIAS.n271 CS_BIAS.n270 0.189894
R1160 CS_BIAS.n270 CS_BIAS.n12 0.189894
R1161 CS_BIAS.n266 CS_BIAS.n12 0.189894
R1162 CS_BIAS.n266 CS_BIAS.n265 0.189894
R1163 CS_BIAS.n265 CS_BIAS.n14 0.189894
R1164 CS_BIAS.n261 CS_BIAS.n14 0.189894
R1165 CS_BIAS.n261 CS_BIAS.n260 0.189894
R1166 CS_BIAS.n260 CS_BIAS.n259 0.189894
R1167 CS_BIAS.n259 CS_BIAS.n16 0.189894
R1168 CS_BIAS.n255 CS_BIAS.n16 0.189894
R1169 CS_BIAS.n255 CS_BIAS.n254 0.189894
R1170 CS_BIAS.n254 CS_BIAS.n253 0.189894
R1171 CS_BIAS.n253 CS_BIAS.n18 0.189894
R1172 CS_BIAS.n249 CS_BIAS.n18 0.189894
R1173 CS_BIAS.n249 CS_BIAS.n248 0.189894
R1174 CS_BIAS.n248 CS_BIAS.n247 0.189894
R1175 CS_BIAS.n247 CS_BIAS.n20 0.189894
R1176 CS_BIAS.n243 CS_BIAS.n20 0.189894
R1177 CS_BIAS.n243 CS_BIAS.n242 0.189894
R1178 CS_BIAS.n242 CS_BIAS.n241 0.189894
R1179 CS_BIAS.n790 CS_BIAS.n787 0.189894
R1180 CS_BIAS.n794 CS_BIAS.n787 0.189894
R1181 CS_BIAS.n795 CS_BIAS.n794 0.189894
R1182 CS_BIAS.n796 CS_BIAS.n795 0.189894
R1183 CS_BIAS.n796 CS_BIAS.n785 0.189894
R1184 CS_BIAS.n800 CS_BIAS.n785 0.189894
R1185 CS_BIAS.n801 CS_BIAS.n800 0.189894
R1186 CS_BIAS.n802 CS_BIAS.n801 0.189894
R1187 CS_BIAS.n802 CS_BIAS.n783 0.189894
R1188 CS_BIAS.n807 CS_BIAS.n783 0.189894
R1189 CS_BIAS.n808 CS_BIAS.n807 0.189894
R1190 CS_BIAS.n809 CS_BIAS.n808 0.189894
R1191 CS_BIAS.n809 CS_BIAS.n781 0.189894
R1192 CS_BIAS.n813 CS_BIAS.n781 0.189894
R1193 CS_BIAS.n814 CS_BIAS.n813 0.189894
R1194 CS_BIAS.n815 CS_BIAS.n814 0.189894
R1195 CS_BIAS.n815 CS_BIAS.n779 0.189894
R1196 CS_BIAS.n819 CS_BIAS.n779 0.189894
R1197 CS_BIAS.n820 CS_BIAS.n819 0.189894
R1198 CS_BIAS.n821 CS_BIAS.n820 0.189894
R1199 CS_BIAS.n821 CS_BIAS.n777 0.189894
R1200 CS_BIAS.n825 CS_BIAS.n777 0.189894
R1201 CS_BIAS.n826 CS_BIAS.n825 0.189894
R1202 CS_BIAS.n826 CS_BIAS.n775 0.189894
R1203 CS_BIAS.n830 CS_BIAS.n775 0.189894
R1204 CS_BIAS.n831 CS_BIAS.n830 0.189894
R1205 CS_BIAS.n832 CS_BIAS.n831 0.189894
R1206 CS_BIAS.n832 CS_BIAS.n773 0.189894
R1207 CS_BIAS.n836 CS_BIAS.n773 0.189894
R1208 CS_BIAS.n837 CS_BIAS.n836 0.189894
R1209 CS_BIAS.n838 CS_BIAS.n837 0.189894
R1210 CS_BIAS.n838 CS_BIAS.n771 0.189894
R1211 CS_BIAS.n843 CS_BIAS.n771 0.189894
R1212 CS_BIAS.n844 CS_BIAS.n843 0.189894
R1213 CS_BIAS.n845 CS_BIAS.n844 0.189894
R1214 CS_BIAS.n845 CS_BIAS.n769 0.189894
R1215 CS_BIAS.n849 CS_BIAS.n769 0.189894
R1216 CS_BIAS.n850 CS_BIAS.n849 0.189894
R1217 CS_BIAS.n851 CS_BIAS.n850 0.189894
R1218 CS_BIAS.n851 CS_BIAS.n767 0.189894
R1219 CS_BIAS.n855 CS_BIAS.n767 0.189894
R1220 CS_BIAS.n856 CS_BIAS.n855 0.189894
R1221 CS_BIAS.n857 CS_BIAS.n856 0.189894
R1222 CS_BIAS.n857 CS_BIAS.n765 0.189894
R1223 CS_BIAS.n861 CS_BIAS.n765 0.189894
R1224 CS_BIAS.n862 CS_BIAS.n861 0.189894
R1225 CS_BIAS.n862 CS_BIAS.n763 0.189894
R1226 CS_BIAS.n866 CS_BIAS.n763 0.189894
R1227 CS_BIAS.n867 CS_BIAS.n866 0.189894
R1228 CS_BIAS.n868 CS_BIAS.n867 0.189894
R1229 CS_BIAS.n868 CS_BIAS.n761 0.189894
R1230 CS_BIAS.n872 CS_BIAS.n761 0.189894
R1231 CS_BIAS.n873 CS_BIAS.n872 0.189894
R1232 CS_BIAS.n874 CS_BIAS.n873 0.189894
R1233 CS_BIAS.n874 CS_BIAS.n759 0.189894
R1234 CS_BIAS.n879 CS_BIAS.n759 0.189894
R1235 CS_BIAS.n880 CS_BIAS.n879 0.189894
R1236 CS_BIAS.n881 CS_BIAS.n880 0.189894
R1237 CS_BIAS.n881 CS_BIAS.n757 0.189894
R1238 CS_BIAS.n885 CS_BIAS.n757 0.189894
R1239 CS_BIAS.n886 CS_BIAS.n885 0.189894
R1240 CS_BIAS.n887 CS_BIAS.n886 0.189894
R1241 CS_BIAS.n887 CS_BIAS.n755 0.189894
R1242 CS_BIAS.n891 CS_BIAS.n755 0.189894
R1243 CS_BIAS.n892 CS_BIAS.n891 0.189894
R1244 CS_BIAS.n893 CS_BIAS.n892 0.189894
R1245 CS_BIAS.n893 CS_BIAS.n753 0.189894
R1246 CS_BIAS.n897 CS_BIAS.n753 0.189894
R1247 CS_BIAS.n512 CS_BIAS.n509 0.189894
R1248 CS_BIAS.n516 CS_BIAS.n509 0.189894
R1249 CS_BIAS.n517 CS_BIAS.n516 0.189894
R1250 CS_BIAS.n518 CS_BIAS.n517 0.189894
R1251 CS_BIAS.n518 CS_BIAS.n507 0.189894
R1252 CS_BIAS.n522 CS_BIAS.n507 0.189894
R1253 CS_BIAS.n523 CS_BIAS.n522 0.189894
R1254 CS_BIAS.n524 CS_BIAS.n523 0.189894
R1255 CS_BIAS.n524 CS_BIAS.n505 0.189894
R1256 CS_BIAS.n529 CS_BIAS.n505 0.189894
R1257 CS_BIAS.n530 CS_BIAS.n529 0.189894
R1258 CS_BIAS.n531 CS_BIAS.n530 0.189894
R1259 CS_BIAS.n531 CS_BIAS.n503 0.189894
R1260 CS_BIAS.n535 CS_BIAS.n503 0.189894
R1261 CS_BIAS.n536 CS_BIAS.n535 0.189894
R1262 CS_BIAS.n537 CS_BIAS.n536 0.189894
R1263 CS_BIAS.n537 CS_BIAS.n501 0.189894
R1264 CS_BIAS.n541 CS_BIAS.n501 0.189894
R1265 CS_BIAS.n542 CS_BIAS.n541 0.189894
R1266 CS_BIAS.n543 CS_BIAS.n542 0.189894
R1267 CS_BIAS.n543 CS_BIAS.n499 0.189894
R1268 CS_BIAS.n547 CS_BIAS.n499 0.189894
R1269 CS_BIAS.n548 CS_BIAS.n547 0.189894
R1270 CS_BIAS.n548 CS_BIAS.n497 0.189894
R1271 CS_BIAS.n552 CS_BIAS.n497 0.189894
R1272 CS_BIAS.n553 CS_BIAS.n552 0.189894
R1273 CS_BIAS.n554 CS_BIAS.n553 0.189894
R1274 CS_BIAS.n554 CS_BIAS.n495 0.189894
R1275 CS_BIAS.n558 CS_BIAS.n495 0.189894
R1276 CS_BIAS.n559 CS_BIAS.n558 0.189894
R1277 CS_BIAS.n560 CS_BIAS.n559 0.189894
R1278 CS_BIAS.n560 CS_BIAS.n493 0.189894
R1279 CS_BIAS.n565 CS_BIAS.n493 0.189894
R1280 CS_BIAS.n566 CS_BIAS.n565 0.189894
R1281 CS_BIAS.n567 CS_BIAS.n566 0.189894
R1282 CS_BIAS.n567 CS_BIAS.n491 0.189894
R1283 CS_BIAS.n571 CS_BIAS.n491 0.189894
R1284 CS_BIAS.n572 CS_BIAS.n571 0.189894
R1285 CS_BIAS.n573 CS_BIAS.n572 0.189894
R1286 CS_BIAS.n573 CS_BIAS.n489 0.189894
R1287 CS_BIAS.n577 CS_BIAS.n489 0.189894
R1288 CS_BIAS.n578 CS_BIAS.n577 0.189894
R1289 CS_BIAS.n579 CS_BIAS.n578 0.189894
R1290 CS_BIAS.n579 CS_BIAS.n487 0.189894
R1291 CS_BIAS.n583 CS_BIAS.n487 0.189894
R1292 CS_BIAS.n584 CS_BIAS.n583 0.189894
R1293 CS_BIAS.n584 CS_BIAS.n485 0.189894
R1294 CS_BIAS.n588 CS_BIAS.n485 0.189894
R1295 CS_BIAS.n589 CS_BIAS.n588 0.189894
R1296 CS_BIAS.n590 CS_BIAS.n589 0.189894
R1297 CS_BIAS.n590 CS_BIAS.n483 0.189894
R1298 CS_BIAS.n594 CS_BIAS.n483 0.189894
R1299 CS_BIAS.n595 CS_BIAS.n594 0.189894
R1300 CS_BIAS.n596 CS_BIAS.n595 0.189894
R1301 CS_BIAS.n596 CS_BIAS.n481 0.189894
R1302 CS_BIAS.n601 CS_BIAS.n481 0.189894
R1303 CS_BIAS.n602 CS_BIAS.n601 0.189894
R1304 CS_BIAS.n603 CS_BIAS.n602 0.189894
R1305 CS_BIAS.n603 CS_BIAS.n479 0.189894
R1306 CS_BIAS.n607 CS_BIAS.n479 0.189894
R1307 CS_BIAS.n608 CS_BIAS.n607 0.189894
R1308 CS_BIAS.n609 CS_BIAS.n608 0.189894
R1309 CS_BIAS.n609 CS_BIAS.n477 0.189894
R1310 CS_BIAS.n613 CS_BIAS.n477 0.189894
R1311 CS_BIAS.n614 CS_BIAS.n613 0.189894
R1312 CS_BIAS.n615 CS_BIAS.n614 0.189894
R1313 CS_BIAS.n615 CS_BIAS.n475 0.189894
R1314 CS_BIAS.n619 CS_BIAS.n475 0.189894
R1315 CS_BIAS.n643 CS_BIAS.n640 0.189894
R1316 CS_BIAS.n647 CS_BIAS.n640 0.189894
R1317 CS_BIAS.n648 CS_BIAS.n647 0.189894
R1318 CS_BIAS.n649 CS_BIAS.n648 0.189894
R1319 CS_BIAS.n649 CS_BIAS.n638 0.189894
R1320 CS_BIAS.n653 CS_BIAS.n638 0.189894
R1321 CS_BIAS.n654 CS_BIAS.n653 0.189894
R1322 CS_BIAS.n655 CS_BIAS.n654 0.189894
R1323 CS_BIAS.n655 CS_BIAS.n636 0.189894
R1324 CS_BIAS.n660 CS_BIAS.n636 0.189894
R1325 CS_BIAS.n661 CS_BIAS.n660 0.189894
R1326 CS_BIAS.n662 CS_BIAS.n661 0.189894
R1327 CS_BIAS.n662 CS_BIAS.n634 0.189894
R1328 CS_BIAS.n666 CS_BIAS.n634 0.189894
R1329 CS_BIAS.n667 CS_BIAS.n666 0.189894
R1330 CS_BIAS.n668 CS_BIAS.n667 0.189894
R1331 CS_BIAS.n668 CS_BIAS.n632 0.189894
R1332 CS_BIAS.n672 CS_BIAS.n632 0.189894
R1333 CS_BIAS.n673 CS_BIAS.n672 0.189894
R1334 CS_BIAS.n674 CS_BIAS.n673 0.189894
R1335 CS_BIAS.n674 CS_BIAS.n630 0.189894
R1336 CS_BIAS.n678 CS_BIAS.n630 0.189894
R1337 CS_BIAS.n679 CS_BIAS.n678 0.189894
R1338 CS_BIAS.n679 CS_BIAS.n628 0.189894
R1339 CS_BIAS.n683 CS_BIAS.n628 0.189894
R1340 CS_BIAS.n684 CS_BIAS.n683 0.189894
R1341 CS_BIAS.n685 CS_BIAS.n684 0.189894
R1342 CS_BIAS.n690 CS_BIAS.n689 0.189894
R1343 CS_BIAS.n691 CS_BIAS.n690 0.189894
R1344 CS_BIAS.n691 CS_BIAS.n469 0.189894
R1345 CS_BIAS.n696 CS_BIAS.n469 0.189894
R1346 CS_BIAS.n697 CS_BIAS.n696 0.189894
R1347 CS_BIAS.n698 CS_BIAS.n697 0.189894
R1348 CS_BIAS.n698 CS_BIAS.n467 0.189894
R1349 CS_BIAS.n702 CS_BIAS.n467 0.189894
R1350 CS_BIAS.n703 CS_BIAS.n702 0.189894
R1351 CS_BIAS.n704 CS_BIAS.n703 0.189894
R1352 CS_BIAS.n704 CS_BIAS.n465 0.189894
R1353 CS_BIAS.n708 CS_BIAS.n465 0.189894
R1354 CS_BIAS.n709 CS_BIAS.n708 0.189894
R1355 CS_BIAS.n710 CS_BIAS.n709 0.189894
R1356 CS_BIAS.n710 CS_BIAS.n463 0.189894
R1357 CS_BIAS.n714 CS_BIAS.n463 0.189894
R1358 CS_BIAS.n715 CS_BIAS.n714 0.189894
R1359 CS_BIAS.n715 CS_BIAS.n461 0.189894
R1360 CS_BIAS.n719 CS_BIAS.n461 0.189894
R1361 CS_BIAS.n720 CS_BIAS.n719 0.189894
R1362 CS_BIAS.n721 CS_BIAS.n720 0.189894
R1363 CS_BIAS.n721 CS_BIAS.n459 0.189894
R1364 CS_BIAS.n725 CS_BIAS.n459 0.189894
R1365 CS_BIAS.n726 CS_BIAS.n725 0.189894
R1366 CS_BIAS.n727 CS_BIAS.n726 0.189894
R1367 CS_BIAS.n727 CS_BIAS.n457 0.189894
R1368 CS_BIAS.n732 CS_BIAS.n457 0.189894
R1369 CS_BIAS.n733 CS_BIAS.n732 0.189894
R1370 CS_BIAS.n734 CS_BIAS.n733 0.189894
R1371 CS_BIAS.n734 CS_BIAS.n455 0.189894
R1372 CS_BIAS.n738 CS_BIAS.n455 0.189894
R1373 CS_BIAS.n739 CS_BIAS.n738 0.189894
R1374 CS_BIAS.n740 CS_BIAS.n739 0.189894
R1375 CS_BIAS.n740 CS_BIAS.n453 0.189894
R1376 CS_BIAS.n744 CS_BIAS.n453 0.189894
R1377 CS_BIAS.n745 CS_BIAS.n744 0.189894
R1378 CS_BIAS.n746 CS_BIAS.n745 0.189894
R1379 CS_BIAS.n746 CS_BIAS.n451 0.189894
R1380 CS_BIAS.n750 CS_BIAS.n451 0.189894
R1381 CS_BIAS.n237 CS_BIAS.n178 0.170955
R1382 CS_BIAS.n241 CS_BIAS.n178 0.170955
R1383 CS_BIAS.n685 CS_BIAS.n626 0.170955
R1384 CS_BIAS.n689 CS_BIAS.n626 0.170955
R1385 GND.n5023 GND.n3523 824.038
R1386 GND.n4307 GND.n4078 824.038
R1387 GND.n4191 GND.n295 824.038
R1388 GND.n5033 GND.n2786 824.038
R1389 GND.n7463 GND.n523 766.379
R1390 GND.n7426 GND.n565 766.379
R1391 GND.n6735 GND.n930 766.379
R1392 GND.n6723 GND.n932 766.379
R1393 GND.n5566 GND.n1738 766.379
R1394 GND.n5692 GND.n1736 766.379
R1395 GND.n3186 GND.n3049 766.379
R1396 GND.n3184 GND.n3053 766.379
R1397 GND.n4306 GND.n4305 746.404
R1398 GND.n1340 GND.n1335 739.952
R1399 GND.n6277 GND.n6276 739.952
R1400 GND.n5725 GND.n1684 739.952
R1401 GND.n5820 GND.n1682 739.952
R1402 GND.n7344 GND.n519 713.524
R1403 GND.n7327 GND.n584 713.524
R1404 GND.n950 GND.n934 713.524
R1405 GND.n1345 GND.n933 713.524
R1406 GND.n1776 GND.n1739 713.524
R1407 GND.n1750 GND.n1741 713.524
R1408 GND.n3115 GND.n3051 713.524
R1409 GND.n3135 GND.n3052 713.524
R1410 GND.n1346 GND.n1345 589.749
R1411 GND.n1776 GND.n1726 589.749
R1412 GND.n1370 GND.n950 588.616
R1413 GND.n3482 GND.n2781 585
R1414 GND.n3520 GND.n2781 585
R1415 GND.n2830 GND.n2828 585
R1416 GND.n2828 GND.n2790 585
R1417 GND.n3491 GND.n3490 585
R1418 GND.n3492 GND.n3491 585
R1419 GND.n2829 GND.n2827 585
R1420 GND.n2827 GND.n2824 585
R1421 GND.n2851 GND.n2837 585
R1422 GND.n3477 GND.n2837 585
R1423 GND.n2849 GND.n2847 585
R1424 GND.n2847 GND.n2835 585
R1425 GND.n3468 GND.n3467 585
R1426 GND.n3469 GND.n3468 585
R1427 GND.n2848 GND.n2846 585
R1428 GND.n2846 GND.n2843 585
R1429 GND.n2872 GND.n2858 585
R1430 GND.n3460 GND.n2858 585
R1431 GND.n2870 GND.n2868 585
R1432 GND.n2868 GND.n2856 585
R1433 GND.n3451 GND.n3450 585
R1434 GND.n3452 GND.n3451 585
R1435 GND.n2869 GND.n2867 585
R1436 GND.n2867 GND.n2864 585
R1437 GND.n2893 GND.n2879 585
R1438 GND.n3443 GND.n2879 585
R1439 GND.n2891 GND.n2889 585
R1440 GND.n2889 GND.n2877 585
R1441 GND.n3434 GND.n3433 585
R1442 GND.n3435 GND.n3434 585
R1443 GND.n2890 GND.n2888 585
R1444 GND.n2888 GND.n2885 585
R1445 GND.n2914 GND.n2900 585
R1446 GND.n3426 GND.n2900 585
R1447 GND.n2912 GND.n2910 585
R1448 GND.n2910 GND.n2898 585
R1449 GND.n3417 GND.n3416 585
R1450 GND.n3418 GND.n3417 585
R1451 GND.n2911 GND.n2909 585
R1452 GND.n2909 GND.n2906 585
R1453 GND.n2935 GND.n2921 585
R1454 GND.n3409 GND.n2921 585
R1455 GND.n2933 GND.n2931 585
R1456 GND.n2931 GND.n2919 585
R1457 GND.n3400 GND.n3399 585
R1458 GND.n3401 GND.n3400 585
R1459 GND.n2932 GND.n2930 585
R1460 GND.n2930 GND.n2927 585
R1461 GND.n2956 GND.n2941 585
R1462 GND.n3392 GND.n2941 585
R1463 GND.n2954 GND.n2952 585
R1464 GND.n2952 GND.n2950 585
R1465 GND.n3383 GND.n3382 585
R1466 GND.n3384 GND.n3383 585
R1467 GND.n2953 GND.n2951 585
R1468 GND.n2951 GND.n2947 585
R1469 GND.n2977 GND.n2963 585
R1470 GND.n3375 GND.n2963 585
R1471 GND.n2975 GND.n2973 585
R1472 GND.n2973 GND.n2961 585
R1473 GND.n3366 GND.n3365 585
R1474 GND.n3367 GND.n3366 585
R1475 GND.n2974 GND.n2972 585
R1476 GND.n2972 GND.n2969 585
R1477 GND.n2998 GND.n2984 585
R1478 GND.n3358 GND.n2984 585
R1479 GND.n2996 GND.n2994 585
R1480 GND.n2994 GND.n2982 585
R1481 GND.n3349 GND.n3348 585
R1482 GND.n3350 GND.n3349 585
R1483 GND.n2995 GND.n2993 585
R1484 GND.n2993 GND.n2990 585
R1485 GND.n3018 GND.n3005 585
R1486 GND.n3341 GND.n3005 585
R1487 GND.n3016 GND.n3014 585
R1488 GND.n3014 GND.n3003 585
R1489 GND.n3332 GND.n3331 585
R1490 GND.n3333 GND.n3332 585
R1491 GND.n3015 GND.n3013 585
R1492 GND.n3325 GND.n3013 585
R1493 GND.n3192 GND.n3191 585
R1494 GND.n3191 GND.n3023 585
R1495 GND.n3190 GND.n3032 585
R1496 GND.n3211 GND.n3032 585
R1497 GND.n3045 GND.n3043 585
R1498 GND.n3043 GND.n3030 585
R1499 GND.n3200 GND.n3199 585
R1500 GND.n3201 GND.n3200 585
R1501 GND.n3044 GND.n3042 585
R1502 GND.n3042 GND.n3039 585
R1503 GND.n3089 GND.n3052 585
R1504 GND.n3185 GND.n3052 585
R1505 GND.n3136 GND.n3135 585
R1506 GND.n3133 GND.n3092 585
R1507 GND.n3132 GND.n3131 585
R1508 GND.n3096 GND.n3094 585
R1509 GND.n3127 GND.n3097 585
R1510 GND.n3126 GND.n3099 585
R1511 GND.n3125 GND.n3100 585
R1512 GND.n3104 GND.n3101 585
R1513 GND.n3121 GND.n3105 585
R1514 GND.n3120 GND.n3117 585
R1515 GND.n3115 GND.n3114 585
R1516 GND.n3115 GND.n3050 585
R1517 GND.n3264 GND.n2818 585
R1518 GND.n3520 GND.n2818 585
R1519 GND.n3265 GND.n3253 585
R1520 GND.n3253 GND.n2790 585
R1521 GND.n3251 GND.n2826 585
R1522 GND.n3492 GND.n2826 585
R1523 GND.n3269 GND.n3250 585
R1524 GND.n3250 GND.n2824 585
R1525 GND.n3270 GND.n2836 585
R1526 GND.n3477 GND.n2836 585
R1527 GND.n3271 GND.n3249 585
R1528 GND.n3249 GND.n2835 585
R1529 GND.n3247 GND.n2845 585
R1530 GND.n3469 GND.n2845 585
R1531 GND.n3275 GND.n3246 585
R1532 GND.n3246 GND.n2843 585
R1533 GND.n3276 GND.n2857 585
R1534 GND.n3460 GND.n2857 585
R1535 GND.n3277 GND.n3245 585
R1536 GND.n3245 GND.n2856 585
R1537 GND.n3243 GND.n2866 585
R1538 GND.n3452 GND.n2866 585
R1539 GND.n3281 GND.n3242 585
R1540 GND.n3242 GND.n2864 585
R1541 GND.n3282 GND.n2878 585
R1542 GND.n3443 GND.n2878 585
R1543 GND.n3283 GND.n3241 585
R1544 GND.n3241 GND.n2877 585
R1545 GND.n3239 GND.n2887 585
R1546 GND.n3435 GND.n2887 585
R1547 GND.n3287 GND.n3238 585
R1548 GND.n3238 GND.n2885 585
R1549 GND.n3288 GND.n2899 585
R1550 GND.n3426 GND.n2899 585
R1551 GND.n3289 GND.n3237 585
R1552 GND.n3237 GND.n2898 585
R1553 GND.n3235 GND.n2908 585
R1554 GND.n3418 GND.n2908 585
R1555 GND.n3293 GND.n3234 585
R1556 GND.n3234 GND.n2906 585
R1557 GND.n3294 GND.n2920 585
R1558 GND.n3409 GND.n2920 585
R1559 GND.n3295 GND.n3233 585
R1560 GND.n3233 GND.n2919 585
R1561 GND.n3231 GND.n2929 585
R1562 GND.n3401 GND.n2929 585
R1563 GND.n3299 GND.n3230 585
R1564 GND.n3230 GND.n2927 585
R1565 GND.n3300 GND.n2940 585
R1566 GND.n3392 GND.n2940 585
R1567 GND.n3301 GND.n3229 585
R1568 GND.n3229 GND.n2950 585
R1569 GND.n3227 GND.n2949 585
R1570 GND.n3384 GND.n2949 585
R1571 GND.n3305 GND.n3226 585
R1572 GND.n3226 GND.n2947 585
R1573 GND.n3306 GND.n2962 585
R1574 GND.n3375 GND.n2962 585
R1575 GND.n3307 GND.n3225 585
R1576 GND.n3225 GND.n2961 585
R1577 GND.n3223 GND.n2971 585
R1578 GND.n3367 GND.n2971 585
R1579 GND.n3311 GND.n3222 585
R1580 GND.n3222 GND.n2969 585
R1581 GND.n3312 GND.n2983 585
R1582 GND.n3358 GND.n2983 585
R1583 GND.n3313 GND.n3221 585
R1584 GND.n3221 GND.n2982 585
R1585 GND.n3219 GND.n2992 585
R1586 GND.n3350 GND.n2992 585
R1587 GND.n3317 GND.n3218 585
R1588 GND.n3218 GND.n2990 585
R1589 GND.n3318 GND.n3004 585
R1590 GND.n3341 GND.n3004 585
R1591 GND.n3319 GND.n3217 585
R1592 GND.n3217 GND.n3003 585
R1593 GND.n3026 GND.n3012 585
R1594 GND.n3333 GND.n3012 585
R1595 GND.n3324 GND.n3323 585
R1596 GND.n3325 GND.n3324 585
R1597 GND.n3025 GND.n3024 585
R1598 GND.n3024 GND.n3023 585
R1599 GND.n3213 GND.n3212 585
R1600 GND.n3212 GND.n3211 585
R1601 GND.n3029 GND.n3028 585
R1602 GND.n3030 GND.n3029 585
R1603 GND.n3109 GND.n3041 585
R1604 GND.n3201 GND.n3041 585
R1605 GND.n3110 GND.n3107 585
R1606 GND.n3107 GND.n3039 585
R1607 GND.n3111 GND.n3051 585
R1608 GND.n3185 GND.n3051 585
R1609 GND.n3519 GND.n3518 585
R1610 GND.n3520 GND.n3519 585
R1611 GND.n2820 GND.n2819 585
R1612 GND.n2819 GND.n2790 585
R1613 GND.n3494 GND.n3493 585
R1614 GND.n3493 GND.n3492 585
R1615 GND.n2823 GND.n2822 585
R1616 GND.n2824 GND.n2823 585
R1617 GND.n3476 GND.n3475 585
R1618 GND.n3477 GND.n3476 585
R1619 GND.n2839 GND.n2838 585
R1620 GND.n2838 GND.n2835 585
R1621 GND.n3471 GND.n3470 585
R1622 GND.n3470 GND.n3469 585
R1623 GND.n2842 GND.n2841 585
R1624 GND.n2843 GND.n2842 585
R1625 GND.n3459 GND.n3458 585
R1626 GND.n3460 GND.n3459 585
R1627 GND.n2860 GND.n2859 585
R1628 GND.n2859 GND.n2856 585
R1629 GND.n3454 GND.n3453 585
R1630 GND.n3453 GND.n3452 585
R1631 GND.n2863 GND.n2862 585
R1632 GND.n2864 GND.n2863 585
R1633 GND.n3442 GND.n3441 585
R1634 GND.n3443 GND.n3442 585
R1635 GND.n2881 GND.n2880 585
R1636 GND.n2880 GND.n2877 585
R1637 GND.n3437 GND.n3436 585
R1638 GND.n3436 GND.n3435 585
R1639 GND.n2884 GND.n2883 585
R1640 GND.n2885 GND.n2884 585
R1641 GND.n3425 GND.n3424 585
R1642 GND.n3426 GND.n3425 585
R1643 GND.n2902 GND.n2901 585
R1644 GND.n2901 GND.n2898 585
R1645 GND.n3420 GND.n3419 585
R1646 GND.n3419 GND.n3418 585
R1647 GND.n2905 GND.n2904 585
R1648 GND.n2906 GND.n2905 585
R1649 GND.n3408 GND.n3407 585
R1650 GND.n3409 GND.n3408 585
R1651 GND.n2923 GND.n2922 585
R1652 GND.n2922 GND.n2919 585
R1653 GND.n3403 GND.n3402 585
R1654 GND.n3402 GND.n3401 585
R1655 GND.n2926 GND.n2925 585
R1656 GND.n2927 GND.n2926 585
R1657 GND.n3391 GND.n3390 585
R1658 GND.n3392 GND.n3391 585
R1659 GND.n2943 GND.n2942 585
R1660 GND.n2950 GND.n2942 585
R1661 GND.n3386 GND.n3385 585
R1662 GND.n3385 GND.n3384 585
R1663 GND.n2946 GND.n2945 585
R1664 GND.n2947 GND.n2946 585
R1665 GND.n3374 GND.n3373 585
R1666 GND.n3375 GND.n3374 585
R1667 GND.n2965 GND.n2964 585
R1668 GND.n2964 GND.n2961 585
R1669 GND.n3369 GND.n3368 585
R1670 GND.n3368 GND.n3367 585
R1671 GND.n2968 GND.n2967 585
R1672 GND.n2969 GND.n2968 585
R1673 GND.n3357 GND.n3356 585
R1674 GND.n3358 GND.n3357 585
R1675 GND.n2986 GND.n2985 585
R1676 GND.n2985 GND.n2982 585
R1677 GND.n3352 GND.n3351 585
R1678 GND.n3351 GND.n3350 585
R1679 GND.n2989 GND.n2988 585
R1680 GND.n2990 GND.n2989 585
R1681 GND.n3340 GND.n3339 585
R1682 GND.n3341 GND.n3340 585
R1683 GND.n3007 GND.n3006 585
R1684 GND.n3006 GND.n3003 585
R1685 GND.n3335 GND.n3334 585
R1686 GND.n3334 GND.n3333 585
R1687 GND.n3010 GND.n3009 585
R1688 GND.n3325 GND.n3010 585
R1689 GND.n3208 GND.n3034 585
R1690 GND.n3034 GND.n3023 585
R1691 GND.n3210 GND.n3209 585
R1692 GND.n3211 GND.n3210 585
R1693 GND.n3035 GND.n3033 585
R1694 GND.n3033 GND.n3030 585
R1695 GND.n3203 GND.n3202 585
R1696 GND.n3202 GND.n3201 585
R1697 GND.n3038 GND.n3037 585
R1698 GND.n3039 GND.n3038 585
R1699 GND.n3184 GND.n3183 585
R1700 GND.n3185 GND.n3184 585
R1701 GND.n3180 GND.n3053 585
R1702 GND.n3179 GND.n3178 585
R1703 GND.n3176 GND.n3055 585
R1704 GND.n3176 GND.n3050 585
R1705 GND.n3175 GND.n3174 585
R1706 GND.n3173 GND.n3172 585
R1707 GND.n3171 GND.n3060 585
R1708 GND.n3169 GND.n3168 585
R1709 GND.n3167 GND.n3061 585
R1710 GND.n3166 GND.n3165 585
R1711 GND.n3163 GND.n3068 585
R1712 GND.n3161 GND.n3160 585
R1713 GND.n3159 GND.n3069 585
R1714 GND.n3158 GND.n3157 585
R1715 GND.n3155 GND.n3074 585
R1716 GND.n3153 GND.n3152 585
R1717 GND.n3151 GND.n3075 585
R1718 GND.n3150 GND.n3149 585
R1719 GND.n3147 GND.n3080 585
R1720 GND.n3145 GND.n3144 585
R1721 GND.n3143 GND.n3081 585
R1722 GND.n3088 GND.n3085 585
R1723 GND.n3139 GND.n3049 585
R1724 GND.n3050 GND.n3049 585
R1725 GND.n3486 GND.n2817 585
R1726 GND.n3520 GND.n2817 585
R1727 GND.n3487 GND.n3481 585
R1728 GND.n3481 GND.n2790 585
R1729 GND.n3488 GND.n2825 585
R1730 GND.n3492 GND.n2825 585
R1731 GND.n3480 GND.n3479 585
R1732 GND.n3479 GND.n2824 585
R1733 GND.n3478 GND.n2833 585
R1734 GND.n3478 GND.n3477 585
R1735 GND.n3464 GND.n2834 585
R1736 GND.n2835 GND.n2834 585
R1737 GND.n3465 GND.n2844 585
R1738 GND.n3469 GND.n2844 585
R1739 GND.n3463 GND.n3462 585
R1740 GND.n3462 GND.n2843 585
R1741 GND.n3461 GND.n2854 585
R1742 GND.n3461 GND.n3460 585
R1743 GND.n3447 GND.n2855 585
R1744 GND.n2856 GND.n2855 585
R1745 GND.n3448 GND.n2865 585
R1746 GND.n3452 GND.n2865 585
R1747 GND.n3446 GND.n3445 585
R1748 GND.n3445 GND.n2864 585
R1749 GND.n3444 GND.n2875 585
R1750 GND.n3444 GND.n3443 585
R1751 GND.n3430 GND.n2876 585
R1752 GND.n2877 GND.n2876 585
R1753 GND.n3431 GND.n2886 585
R1754 GND.n3435 GND.n2886 585
R1755 GND.n3429 GND.n3428 585
R1756 GND.n3428 GND.n2885 585
R1757 GND.n3427 GND.n2896 585
R1758 GND.n3427 GND.n3426 585
R1759 GND.n3413 GND.n2897 585
R1760 GND.n2898 GND.n2897 585
R1761 GND.n3414 GND.n2907 585
R1762 GND.n3418 GND.n2907 585
R1763 GND.n3412 GND.n3411 585
R1764 GND.n3411 GND.n2906 585
R1765 GND.n3410 GND.n2917 585
R1766 GND.n3410 GND.n3409 585
R1767 GND.n3396 GND.n2918 585
R1768 GND.n2919 GND.n2918 585
R1769 GND.n3397 GND.n2928 585
R1770 GND.n3401 GND.n2928 585
R1771 GND.n3395 GND.n3394 585
R1772 GND.n3394 GND.n2927 585
R1773 GND.n3393 GND.n2938 585
R1774 GND.n3393 GND.n3392 585
R1775 GND.n3379 GND.n2939 585
R1776 GND.n2950 GND.n2939 585
R1777 GND.n3380 GND.n2948 585
R1778 GND.n3384 GND.n2948 585
R1779 GND.n3378 GND.n3377 585
R1780 GND.n3377 GND.n2947 585
R1781 GND.n3376 GND.n2959 585
R1782 GND.n3376 GND.n3375 585
R1783 GND.n3362 GND.n2960 585
R1784 GND.n2961 GND.n2960 585
R1785 GND.n3363 GND.n2970 585
R1786 GND.n3367 GND.n2970 585
R1787 GND.n3361 GND.n3360 585
R1788 GND.n3360 GND.n2969 585
R1789 GND.n3359 GND.n2980 585
R1790 GND.n3359 GND.n3358 585
R1791 GND.n3345 GND.n2981 585
R1792 GND.n2982 GND.n2981 585
R1793 GND.n3346 GND.n2991 585
R1794 GND.n3350 GND.n2991 585
R1795 GND.n3344 GND.n3343 585
R1796 GND.n3343 GND.n2990 585
R1797 GND.n3342 GND.n3001 585
R1798 GND.n3342 GND.n3341 585
R1799 GND.n3328 GND.n3002 585
R1800 GND.n3003 GND.n3002 585
R1801 GND.n3329 GND.n3011 585
R1802 GND.n3333 GND.n3011 585
R1803 GND.n3327 GND.n3326 585
R1804 GND.n3326 GND.n3325 585
R1805 GND.n3022 GND.n3021 585
R1806 GND.n3023 GND.n3022 585
R1807 GND.n3195 GND.n3031 585
R1808 GND.n3211 GND.n3031 585
R1809 GND.n3196 GND.n3189 585
R1810 GND.n3189 GND.n3030 585
R1811 GND.n3197 GND.n3040 585
R1812 GND.n3201 GND.n3040 585
R1813 GND.n3188 GND.n3187 585
R1814 GND.n3187 GND.n3039 585
R1815 GND.n3186 GND.n3048 585
R1816 GND.n3186 GND.n3185 585
R1817 GND.n5023 GND.n5022 585
R1818 GND.n5021 GND.n3522 585
R1819 GND.n5020 GND.n3521 585
R1820 GND.n5025 GND.n3521 585
R1821 GND.n5019 GND.n5018 585
R1822 GND.n5017 GND.n5016 585
R1823 GND.n5015 GND.n5014 585
R1824 GND.n5013 GND.n5012 585
R1825 GND.n5011 GND.n5010 585
R1826 GND.n5009 GND.n5008 585
R1827 GND.n5007 GND.n5006 585
R1828 GND.n5005 GND.n5004 585
R1829 GND.n5003 GND.n5002 585
R1830 GND.n5001 GND.n5000 585
R1831 GND.n4999 GND.n4998 585
R1832 GND.n4997 GND.n4996 585
R1833 GND.n4995 GND.n4994 585
R1834 GND.n4993 GND.n4992 585
R1835 GND.n4991 GND.n4990 585
R1836 GND.n4989 GND.n4988 585
R1837 GND.n4987 GND.n4986 585
R1838 GND.n4985 GND.n4984 585
R1839 GND.n4983 GND.n4982 585
R1840 GND.n4981 GND.n4980 585
R1841 GND.n4979 GND.n4978 585
R1842 GND.n4977 GND.n4976 585
R1843 GND.n4975 GND.n4974 585
R1844 GND.n4973 GND.n4972 585
R1845 GND.n4971 GND.n4970 585
R1846 GND.n4969 GND.n4968 585
R1847 GND.n4967 GND.n4966 585
R1848 GND.n4965 GND.n4964 585
R1849 GND.n4963 GND.n4962 585
R1850 GND.n4961 GND.n4960 585
R1851 GND.n4959 GND.n4958 585
R1852 GND.n4957 GND.n4956 585
R1853 GND.n4955 GND.n4954 585
R1854 GND.n4953 GND.n4952 585
R1855 GND.n4951 GND.n4950 585
R1856 GND.n4949 GND.n4948 585
R1857 GND.n4947 GND.n4946 585
R1858 GND.n4945 GND.n4944 585
R1859 GND.n4943 GND.n4942 585
R1860 GND.n4941 GND.n4940 585
R1861 GND.n4939 GND.n4938 585
R1862 GND.n4937 GND.n4936 585
R1863 GND.n4935 GND.n4934 585
R1864 GND.n4933 GND.n4932 585
R1865 GND.n4931 GND.n4930 585
R1866 GND.n4929 GND.n4928 585
R1867 GND.n4927 GND.n4926 585
R1868 GND.n4925 GND.n4924 585
R1869 GND.n4923 GND.n4922 585
R1870 GND.n4921 GND.n4920 585
R1871 GND.n4919 GND.n4918 585
R1872 GND.n2789 GND.n2788 585
R1873 GND.n5028 GND.n5027 585
R1874 GND.n5029 GND.n2786 585
R1875 GND.n4861 GND.n3523 585
R1876 GND.n3527 GND.n3523 585
R1877 GND.n4860 GND.n4859 585
R1878 GND.n4859 GND.n4858 585
R1879 GND.n3526 GND.n3525 585
R1880 GND.n4857 GND.n3526 585
R1881 GND.n4855 GND.n4854 585
R1882 GND.n4856 GND.n4855 585
R1883 GND.n4853 GND.n3529 585
R1884 GND.n3529 GND.n3528 585
R1885 GND.n4852 GND.n4851 585
R1886 GND.n4851 GND.n4850 585
R1887 GND.n3535 GND.n3534 585
R1888 GND.n4849 GND.n3535 585
R1889 GND.n4847 GND.n4846 585
R1890 GND.n4848 GND.n4847 585
R1891 GND.n4845 GND.n3537 585
R1892 GND.n3537 GND.n3536 585
R1893 GND.n4844 GND.n4843 585
R1894 GND.n4843 GND.n4842 585
R1895 GND.n3543 GND.n3542 585
R1896 GND.n4841 GND.n3543 585
R1897 GND.n4839 GND.n4838 585
R1898 GND.n4840 GND.n4839 585
R1899 GND.n4837 GND.n3545 585
R1900 GND.n3545 GND.n3544 585
R1901 GND.n4836 GND.n4835 585
R1902 GND.n4835 GND.n4834 585
R1903 GND.n3551 GND.n3550 585
R1904 GND.n4833 GND.n3551 585
R1905 GND.n4831 GND.n4830 585
R1906 GND.n4832 GND.n4831 585
R1907 GND.n4829 GND.n3553 585
R1908 GND.n3553 GND.n3552 585
R1909 GND.n4828 GND.n4827 585
R1910 GND.n4827 GND.n4826 585
R1911 GND.n3559 GND.n3558 585
R1912 GND.n4825 GND.n3559 585
R1913 GND.n4823 GND.n4822 585
R1914 GND.n4824 GND.n4823 585
R1915 GND.n4821 GND.n3561 585
R1916 GND.n3561 GND.n3560 585
R1917 GND.n4820 GND.n4819 585
R1918 GND.n4819 GND.n4818 585
R1919 GND.n3567 GND.n3566 585
R1920 GND.n4817 GND.n3567 585
R1921 GND.n4815 GND.n4814 585
R1922 GND.n4816 GND.n4815 585
R1923 GND.n4813 GND.n3569 585
R1924 GND.n3569 GND.n3568 585
R1925 GND.n4812 GND.n4811 585
R1926 GND.n4811 GND.n4810 585
R1927 GND.n3575 GND.n3574 585
R1928 GND.n4809 GND.n3575 585
R1929 GND.n4807 GND.n4806 585
R1930 GND.n4808 GND.n4807 585
R1931 GND.n4805 GND.n3577 585
R1932 GND.n3577 GND.n3576 585
R1933 GND.n4804 GND.n4803 585
R1934 GND.n4803 GND.n4802 585
R1935 GND.n3583 GND.n3582 585
R1936 GND.n4801 GND.n3583 585
R1937 GND.n4799 GND.n4798 585
R1938 GND.n4800 GND.n4799 585
R1939 GND.n4797 GND.n3585 585
R1940 GND.n3585 GND.n3584 585
R1941 GND.n4796 GND.n4795 585
R1942 GND.n4795 GND.n4794 585
R1943 GND.n3591 GND.n3590 585
R1944 GND.n4793 GND.n3591 585
R1945 GND.n4791 GND.n4790 585
R1946 GND.n4792 GND.n4791 585
R1947 GND.n4789 GND.n3593 585
R1948 GND.n3593 GND.n3592 585
R1949 GND.n4788 GND.n4787 585
R1950 GND.n4787 GND.n4786 585
R1951 GND.n3599 GND.n3598 585
R1952 GND.n4785 GND.n3599 585
R1953 GND.n4783 GND.n4782 585
R1954 GND.n4784 GND.n4783 585
R1955 GND.n4781 GND.n3601 585
R1956 GND.n3601 GND.n3600 585
R1957 GND.n4780 GND.n4779 585
R1958 GND.n4779 GND.n4778 585
R1959 GND.n3607 GND.n3606 585
R1960 GND.n4777 GND.n3607 585
R1961 GND.n4775 GND.n4774 585
R1962 GND.n4776 GND.n4775 585
R1963 GND.n4773 GND.n3609 585
R1964 GND.n3609 GND.n3608 585
R1965 GND.n4772 GND.n4771 585
R1966 GND.n4771 GND.n4770 585
R1967 GND.n3615 GND.n3614 585
R1968 GND.n4769 GND.n3615 585
R1969 GND.n4767 GND.n4766 585
R1970 GND.n4768 GND.n4767 585
R1971 GND.n4765 GND.n3617 585
R1972 GND.n3617 GND.n3616 585
R1973 GND.n4764 GND.n4763 585
R1974 GND.n4763 GND.n4762 585
R1975 GND.n3623 GND.n3622 585
R1976 GND.n4761 GND.n3623 585
R1977 GND.n4759 GND.n4758 585
R1978 GND.n4760 GND.n4759 585
R1979 GND.n4757 GND.n3625 585
R1980 GND.n3625 GND.n3624 585
R1981 GND.n4756 GND.n4755 585
R1982 GND.n4755 GND.n4754 585
R1983 GND.n3631 GND.n3630 585
R1984 GND.n4753 GND.n3631 585
R1985 GND.n4751 GND.n4750 585
R1986 GND.n4752 GND.n4751 585
R1987 GND.n4749 GND.n3633 585
R1988 GND.n3633 GND.n3632 585
R1989 GND.n4748 GND.n4747 585
R1990 GND.n4747 GND.n4746 585
R1991 GND.n3639 GND.n3638 585
R1992 GND.n4745 GND.n3639 585
R1993 GND.n4743 GND.n4742 585
R1994 GND.n4744 GND.n4743 585
R1995 GND.n4741 GND.n3641 585
R1996 GND.n3641 GND.n3640 585
R1997 GND.n4740 GND.n4739 585
R1998 GND.n4739 GND.n4738 585
R1999 GND.n3647 GND.n3646 585
R2000 GND.n4737 GND.n3647 585
R2001 GND.n4735 GND.n4734 585
R2002 GND.n4736 GND.n4735 585
R2003 GND.n4733 GND.n3649 585
R2004 GND.n3649 GND.n3648 585
R2005 GND.n4732 GND.n4731 585
R2006 GND.n4731 GND.n4730 585
R2007 GND.n3655 GND.n3654 585
R2008 GND.n4729 GND.n3655 585
R2009 GND.n4727 GND.n4726 585
R2010 GND.n4728 GND.n4727 585
R2011 GND.n4725 GND.n3657 585
R2012 GND.n3657 GND.n3656 585
R2013 GND.n4724 GND.n4723 585
R2014 GND.n4723 GND.n4722 585
R2015 GND.n3663 GND.n3662 585
R2016 GND.n4721 GND.n3663 585
R2017 GND.n4719 GND.n4718 585
R2018 GND.n4720 GND.n4719 585
R2019 GND.n4717 GND.n3665 585
R2020 GND.n3665 GND.n3664 585
R2021 GND.n4716 GND.n4715 585
R2022 GND.n4715 GND.n4714 585
R2023 GND.n3671 GND.n3670 585
R2024 GND.n4713 GND.n3671 585
R2025 GND.n4711 GND.n4710 585
R2026 GND.n4712 GND.n4711 585
R2027 GND.n4709 GND.n3673 585
R2028 GND.n3673 GND.n3672 585
R2029 GND.n4708 GND.n4707 585
R2030 GND.n4707 GND.n4706 585
R2031 GND.n3679 GND.n3678 585
R2032 GND.n4705 GND.n3679 585
R2033 GND.n4703 GND.n4702 585
R2034 GND.n4704 GND.n4703 585
R2035 GND.n4701 GND.n3681 585
R2036 GND.n3681 GND.n3680 585
R2037 GND.n4700 GND.n4699 585
R2038 GND.n4699 GND.n4698 585
R2039 GND.n3687 GND.n3686 585
R2040 GND.n4697 GND.n3687 585
R2041 GND.n4695 GND.n4694 585
R2042 GND.n4696 GND.n4695 585
R2043 GND.n4693 GND.n3689 585
R2044 GND.n3689 GND.n3688 585
R2045 GND.n4692 GND.n4691 585
R2046 GND.n4691 GND.n4690 585
R2047 GND.n3695 GND.n3694 585
R2048 GND.n4689 GND.n3695 585
R2049 GND.n4687 GND.n4686 585
R2050 GND.n4688 GND.n4687 585
R2051 GND.n4685 GND.n3697 585
R2052 GND.n3697 GND.n3696 585
R2053 GND.n4684 GND.n4683 585
R2054 GND.n4683 GND.n4682 585
R2055 GND.n3703 GND.n3702 585
R2056 GND.n4681 GND.n3703 585
R2057 GND.n4679 GND.n4678 585
R2058 GND.n4680 GND.n4679 585
R2059 GND.n4677 GND.n3705 585
R2060 GND.n3705 GND.n3704 585
R2061 GND.n4676 GND.n4675 585
R2062 GND.n4675 GND.n4674 585
R2063 GND.n3711 GND.n3710 585
R2064 GND.n4673 GND.n3711 585
R2065 GND.n4671 GND.n4670 585
R2066 GND.n4672 GND.n4671 585
R2067 GND.n4669 GND.n3713 585
R2068 GND.n3713 GND.n3712 585
R2069 GND.n4668 GND.n4667 585
R2070 GND.n4667 GND.n4666 585
R2071 GND.n3719 GND.n3718 585
R2072 GND.n4665 GND.n3719 585
R2073 GND.n4663 GND.n4662 585
R2074 GND.n4664 GND.n4663 585
R2075 GND.n4661 GND.n3721 585
R2076 GND.n3721 GND.n3720 585
R2077 GND.n4660 GND.n4659 585
R2078 GND.n4659 GND.n4658 585
R2079 GND.n3727 GND.n3726 585
R2080 GND.n4657 GND.n3727 585
R2081 GND.n4655 GND.n4654 585
R2082 GND.n4656 GND.n4655 585
R2083 GND.n4653 GND.n3729 585
R2084 GND.n3729 GND.n3728 585
R2085 GND.n4652 GND.n4651 585
R2086 GND.n4651 GND.n4650 585
R2087 GND.n3735 GND.n3734 585
R2088 GND.n4649 GND.n3735 585
R2089 GND.n4647 GND.n4646 585
R2090 GND.n4648 GND.n4647 585
R2091 GND.n4645 GND.n3737 585
R2092 GND.n3737 GND.n3736 585
R2093 GND.n4644 GND.n4643 585
R2094 GND.n4643 GND.n4642 585
R2095 GND.n3743 GND.n3742 585
R2096 GND.n4641 GND.n3743 585
R2097 GND.n4639 GND.n4638 585
R2098 GND.n4640 GND.n4639 585
R2099 GND.n4637 GND.n3745 585
R2100 GND.n3745 GND.n3744 585
R2101 GND.n4636 GND.n4635 585
R2102 GND.n4635 GND.n4634 585
R2103 GND.n3751 GND.n3750 585
R2104 GND.n4633 GND.n3751 585
R2105 GND.n4631 GND.n4630 585
R2106 GND.n4632 GND.n4631 585
R2107 GND.n4629 GND.n3753 585
R2108 GND.n3753 GND.n3752 585
R2109 GND.n4628 GND.n4627 585
R2110 GND.n4627 GND.n4626 585
R2111 GND.n3759 GND.n3758 585
R2112 GND.n4625 GND.n3759 585
R2113 GND.n4623 GND.n4622 585
R2114 GND.n4624 GND.n4623 585
R2115 GND.n4621 GND.n3761 585
R2116 GND.n3761 GND.n3760 585
R2117 GND.n4620 GND.n4619 585
R2118 GND.n4619 GND.n4618 585
R2119 GND.n3767 GND.n3766 585
R2120 GND.n4617 GND.n3767 585
R2121 GND.n4615 GND.n4614 585
R2122 GND.n4616 GND.n4615 585
R2123 GND.n4613 GND.n3769 585
R2124 GND.n3769 GND.n3768 585
R2125 GND.n4612 GND.n4611 585
R2126 GND.n4611 GND.n4610 585
R2127 GND.n3775 GND.n3774 585
R2128 GND.n4609 GND.n3775 585
R2129 GND.n4607 GND.n4606 585
R2130 GND.n4608 GND.n4607 585
R2131 GND.n4605 GND.n3777 585
R2132 GND.n3777 GND.n3776 585
R2133 GND.n4604 GND.n4603 585
R2134 GND.n4603 GND.n4602 585
R2135 GND.n3783 GND.n3782 585
R2136 GND.n4601 GND.n3783 585
R2137 GND.n4599 GND.n4598 585
R2138 GND.n4600 GND.n4599 585
R2139 GND.n4597 GND.n3785 585
R2140 GND.n3785 GND.n3784 585
R2141 GND.n4596 GND.n4595 585
R2142 GND.n4595 GND.n4594 585
R2143 GND.n3791 GND.n3790 585
R2144 GND.n4593 GND.n3791 585
R2145 GND.n4591 GND.n4590 585
R2146 GND.n4592 GND.n4591 585
R2147 GND.n4589 GND.n3793 585
R2148 GND.n3793 GND.n3792 585
R2149 GND.n4588 GND.n4587 585
R2150 GND.n4587 GND.n4586 585
R2151 GND.n3799 GND.n3798 585
R2152 GND.n4585 GND.n3799 585
R2153 GND.n4583 GND.n4582 585
R2154 GND.n4584 GND.n4583 585
R2155 GND.n4581 GND.n3801 585
R2156 GND.n3801 GND.n3800 585
R2157 GND.n4580 GND.n4579 585
R2158 GND.n4579 GND.n4578 585
R2159 GND.n3807 GND.n3806 585
R2160 GND.n4577 GND.n3807 585
R2161 GND.n4575 GND.n4574 585
R2162 GND.n4576 GND.n4575 585
R2163 GND.n4573 GND.n3809 585
R2164 GND.n3809 GND.n3808 585
R2165 GND.n4572 GND.n4571 585
R2166 GND.n4571 GND.n4570 585
R2167 GND.n3815 GND.n3814 585
R2168 GND.n4569 GND.n3815 585
R2169 GND.n4567 GND.n4566 585
R2170 GND.n4568 GND.n4567 585
R2171 GND.n4565 GND.n3817 585
R2172 GND.n3817 GND.n3816 585
R2173 GND.n4564 GND.n4563 585
R2174 GND.n4563 GND.n4562 585
R2175 GND.n3823 GND.n3822 585
R2176 GND.n4561 GND.n3823 585
R2177 GND.n4559 GND.n4558 585
R2178 GND.n4560 GND.n4559 585
R2179 GND.n4557 GND.n3825 585
R2180 GND.n3825 GND.n3824 585
R2181 GND.n4556 GND.n4555 585
R2182 GND.n4555 GND.n4554 585
R2183 GND.n3831 GND.n3830 585
R2184 GND.n4553 GND.n3831 585
R2185 GND.n4551 GND.n4550 585
R2186 GND.n4552 GND.n4551 585
R2187 GND.n4549 GND.n3833 585
R2188 GND.n3833 GND.n3832 585
R2189 GND.n4548 GND.n4547 585
R2190 GND.n4547 GND.n4546 585
R2191 GND.n3839 GND.n3838 585
R2192 GND.n4545 GND.n3839 585
R2193 GND.n4543 GND.n4542 585
R2194 GND.n4544 GND.n4543 585
R2195 GND.n4541 GND.n3841 585
R2196 GND.n3841 GND.n3840 585
R2197 GND.n4540 GND.n4539 585
R2198 GND.n4539 GND.n4538 585
R2199 GND.n3847 GND.n3846 585
R2200 GND.n4537 GND.n3847 585
R2201 GND.n4535 GND.n4534 585
R2202 GND.n4536 GND.n4535 585
R2203 GND.n4533 GND.n3849 585
R2204 GND.n3849 GND.n3848 585
R2205 GND.n4532 GND.n4531 585
R2206 GND.n4531 GND.n4530 585
R2207 GND.n3855 GND.n3854 585
R2208 GND.n4529 GND.n3855 585
R2209 GND.n4527 GND.n4526 585
R2210 GND.n4528 GND.n4527 585
R2211 GND.n4525 GND.n3857 585
R2212 GND.n3857 GND.n3856 585
R2213 GND.n4524 GND.n4523 585
R2214 GND.n4523 GND.n4522 585
R2215 GND.n3863 GND.n3862 585
R2216 GND.n4521 GND.n3863 585
R2217 GND.n4519 GND.n4518 585
R2218 GND.n4520 GND.n4519 585
R2219 GND.n4517 GND.n3865 585
R2220 GND.n3865 GND.n3864 585
R2221 GND.n4516 GND.n4515 585
R2222 GND.n4515 GND.n4514 585
R2223 GND.n3871 GND.n3870 585
R2224 GND.n4513 GND.n3871 585
R2225 GND.n4511 GND.n4510 585
R2226 GND.n4512 GND.n4511 585
R2227 GND.n4509 GND.n3873 585
R2228 GND.n3873 GND.n3872 585
R2229 GND.n4508 GND.n4507 585
R2230 GND.n4507 GND.n4506 585
R2231 GND.n3879 GND.n3878 585
R2232 GND.n4505 GND.n3879 585
R2233 GND.n4503 GND.n4502 585
R2234 GND.n4504 GND.n4503 585
R2235 GND.n4501 GND.n3881 585
R2236 GND.n3881 GND.n3880 585
R2237 GND.n4500 GND.n4499 585
R2238 GND.n4499 GND.n4498 585
R2239 GND.n3887 GND.n3886 585
R2240 GND.n4497 GND.n3887 585
R2241 GND.n4495 GND.n4494 585
R2242 GND.n4496 GND.n4495 585
R2243 GND.n4493 GND.n3889 585
R2244 GND.n3889 GND.n3888 585
R2245 GND.n4492 GND.n4491 585
R2246 GND.n4491 GND.n4490 585
R2247 GND.n3895 GND.n3894 585
R2248 GND.n4489 GND.n3895 585
R2249 GND.n4487 GND.n4486 585
R2250 GND.n4488 GND.n4487 585
R2251 GND.n4485 GND.n3897 585
R2252 GND.n3897 GND.n3896 585
R2253 GND.n4484 GND.n4483 585
R2254 GND.n4483 GND.n4482 585
R2255 GND.n3903 GND.n3902 585
R2256 GND.n4481 GND.n3903 585
R2257 GND.n4479 GND.n4478 585
R2258 GND.n4480 GND.n4479 585
R2259 GND.n4477 GND.n3905 585
R2260 GND.n3905 GND.n3904 585
R2261 GND.n4476 GND.n4475 585
R2262 GND.n4475 GND.n4474 585
R2263 GND.n3911 GND.n3910 585
R2264 GND.n4473 GND.n3911 585
R2265 GND.n4471 GND.n4470 585
R2266 GND.n4472 GND.n4471 585
R2267 GND.n4469 GND.n3913 585
R2268 GND.n3913 GND.n3912 585
R2269 GND.n4468 GND.n4467 585
R2270 GND.n4467 GND.n4466 585
R2271 GND.n3919 GND.n3918 585
R2272 GND.n4465 GND.n3919 585
R2273 GND.n4463 GND.n4462 585
R2274 GND.n4464 GND.n4463 585
R2275 GND.n4461 GND.n3921 585
R2276 GND.n3921 GND.n3920 585
R2277 GND.n4460 GND.n4459 585
R2278 GND.n4459 GND.n4458 585
R2279 GND.n3927 GND.n3926 585
R2280 GND.n4457 GND.n3927 585
R2281 GND.n4455 GND.n4454 585
R2282 GND.n4456 GND.n4455 585
R2283 GND.n4453 GND.n3929 585
R2284 GND.n3929 GND.n3928 585
R2285 GND.n4452 GND.n4451 585
R2286 GND.n4451 GND.n4450 585
R2287 GND.n3935 GND.n3934 585
R2288 GND.n4449 GND.n3935 585
R2289 GND.n4447 GND.n4446 585
R2290 GND.n4448 GND.n4447 585
R2291 GND.n4445 GND.n3937 585
R2292 GND.n3937 GND.n3936 585
R2293 GND.n4444 GND.n4443 585
R2294 GND.n4443 GND.n4442 585
R2295 GND.n3943 GND.n3942 585
R2296 GND.n4441 GND.n3943 585
R2297 GND.n4439 GND.n4438 585
R2298 GND.n4440 GND.n4439 585
R2299 GND.n4437 GND.n3945 585
R2300 GND.n3945 GND.n3944 585
R2301 GND.n4436 GND.n4435 585
R2302 GND.n4435 GND.n4434 585
R2303 GND.n3951 GND.n3950 585
R2304 GND.n4433 GND.n3951 585
R2305 GND.n4431 GND.n4430 585
R2306 GND.n4432 GND.n4431 585
R2307 GND.n4429 GND.n3953 585
R2308 GND.n3953 GND.n3952 585
R2309 GND.n4428 GND.n4427 585
R2310 GND.n4427 GND.n4426 585
R2311 GND.n3959 GND.n3958 585
R2312 GND.n4425 GND.n3959 585
R2313 GND.n4423 GND.n4422 585
R2314 GND.n4424 GND.n4423 585
R2315 GND.n4421 GND.n3961 585
R2316 GND.n3961 GND.n3960 585
R2317 GND.n4420 GND.n4419 585
R2318 GND.n4419 GND.n4418 585
R2319 GND.n3967 GND.n3966 585
R2320 GND.n4417 GND.n3967 585
R2321 GND.n4415 GND.n4414 585
R2322 GND.n4416 GND.n4415 585
R2323 GND.n4413 GND.n3969 585
R2324 GND.n3969 GND.n3968 585
R2325 GND.n4412 GND.n4411 585
R2326 GND.n4411 GND.n4410 585
R2327 GND.n3975 GND.n3974 585
R2328 GND.n4409 GND.n3975 585
R2329 GND.n4407 GND.n4406 585
R2330 GND.n4408 GND.n4407 585
R2331 GND.n4405 GND.n3977 585
R2332 GND.n3977 GND.n3976 585
R2333 GND.n4404 GND.n4403 585
R2334 GND.n4403 GND.n4402 585
R2335 GND.n3983 GND.n3982 585
R2336 GND.n4401 GND.n3983 585
R2337 GND.n4399 GND.n4398 585
R2338 GND.n4400 GND.n4399 585
R2339 GND.n4397 GND.n3985 585
R2340 GND.n3985 GND.n3984 585
R2341 GND.n4396 GND.n4395 585
R2342 GND.n4395 GND.n4394 585
R2343 GND.n3991 GND.n3990 585
R2344 GND.n4393 GND.n3991 585
R2345 GND.n4391 GND.n4390 585
R2346 GND.n4392 GND.n4391 585
R2347 GND.n4389 GND.n3993 585
R2348 GND.n3993 GND.n3992 585
R2349 GND.n4388 GND.n4387 585
R2350 GND.n4387 GND.n4386 585
R2351 GND.n3999 GND.n3998 585
R2352 GND.n4385 GND.n3999 585
R2353 GND.n4383 GND.n4382 585
R2354 GND.n4384 GND.n4383 585
R2355 GND.n4381 GND.n4001 585
R2356 GND.n4001 GND.n4000 585
R2357 GND.n4380 GND.n4379 585
R2358 GND.n4379 GND.n4378 585
R2359 GND.n4007 GND.n4006 585
R2360 GND.n4377 GND.n4007 585
R2361 GND.n4375 GND.n4374 585
R2362 GND.n4376 GND.n4375 585
R2363 GND.n4373 GND.n4009 585
R2364 GND.n4009 GND.n4008 585
R2365 GND.n4372 GND.n4371 585
R2366 GND.n4371 GND.n4370 585
R2367 GND.n4015 GND.n4014 585
R2368 GND.n4369 GND.n4015 585
R2369 GND.n4367 GND.n4366 585
R2370 GND.n4368 GND.n4367 585
R2371 GND.n4365 GND.n4017 585
R2372 GND.n4017 GND.n4016 585
R2373 GND.n4364 GND.n4363 585
R2374 GND.n4363 GND.n4362 585
R2375 GND.n4023 GND.n4022 585
R2376 GND.n4361 GND.n4023 585
R2377 GND.n4359 GND.n4358 585
R2378 GND.n4360 GND.n4359 585
R2379 GND.n4357 GND.n4025 585
R2380 GND.n4025 GND.n4024 585
R2381 GND.n4356 GND.n4355 585
R2382 GND.n4355 GND.n4354 585
R2383 GND.n4031 GND.n4030 585
R2384 GND.n4353 GND.n4031 585
R2385 GND.n4351 GND.n4350 585
R2386 GND.n4352 GND.n4351 585
R2387 GND.n4349 GND.n4033 585
R2388 GND.n4033 GND.n4032 585
R2389 GND.n4348 GND.n4347 585
R2390 GND.n4347 GND.n4346 585
R2391 GND.n4039 GND.n4038 585
R2392 GND.n4345 GND.n4039 585
R2393 GND.n4343 GND.n4342 585
R2394 GND.n4344 GND.n4343 585
R2395 GND.n4341 GND.n4041 585
R2396 GND.n4041 GND.n4040 585
R2397 GND.n4340 GND.n4339 585
R2398 GND.n4339 GND.n4338 585
R2399 GND.n4047 GND.n4046 585
R2400 GND.n4337 GND.n4047 585
R2401 GND.n4335 GND.n4334 585
R2402 GND.n4336 GND.n4335 585
R2403 GND.n4333 GND.n4049 585
R2404 GND.n4049 GND.n4048 585
R2405 GND.n4332 GND.n4331 585
R2406 GND.n4331 GND.n4330 585
R2407 GND.n4055 GND.n4054 585
R2408 GND.n4329 GND.n4055 585
R2409 GND.n4327 GND.n4326 585
R2410 GND.n4328 GND.n4327 585
R2411 GND.n4325 GND.n4057 585
R2412 GND.n4057 GND.n4056 585
R2413 GND.n4324 GND.n4323 585
R2414 GND.n4323 GND.n4322 585
R2415 GND.n4063 GND.n4062 585
R2416 GND.n4321 GND.n4063 585
R2417 GND.n4319 GND.n4318 585
R2418 GND.n4320 GND.n4319 585
R2419 GND.n4317 GND.n4065 585
R2420 GND.n4065 GND.n4064 585
R2421 GND.n4316 GND.n4315 585
R2422 GND.n4315 GND.n4314 585
R2423 GND.n4071 GND.n4070 585
R2424 GND.n4313 GND.n4071 585
R2425 GND.n4311 GND.n4310 585
R2426 GND.n4312 GND.n4311 585
R2427 GND.n4309 GND.n4073 585
R2428 GND.n4073 GND.n4072 585
R2429 GND.n4308 GND.n4307 585
R2430 GND.n4307 GND.n4306 585
R2431 GND.n4194 GND.n4193 585
R2432 GND.n4193 GND.n4192 585
R2433 GND.n4195 GND.n4183 585
R2434 GND.n4183 GND.n4182 585
R2435 GND.n4197 GND.n4196 585
R2436 GND.n4198 GND.n4197 585
R2437 GND.n4181 GND.n4180 585
R2438 GND.n4199 GND.n4181 585
R2439 GND.n4202 GND.n4201 585
R2440 GND.n4201 GND.n4200 585
R2441 GND.n4203 GND.n4175 585
R2442 GND.n4175 GND.n4174 585
R2443 GND.n4205 GND.n4204 585
R2444 GND.n4206 GND.n4205 585
R2445 GND.n4173 GND.n4172 585
R2446 GND.n4207 GND.n4173 585
R2447 GND.n4210 GND.n4209 585
R2448 GND.n4209 GND.n4208 585
R2449 GND.n4211 GND.n4167 585
R2450 GND.n4167 GND.n4166 585
R2451 GND.n4213 GND.n4212 585
R2452 GND.n4214 GND.n4213 585
R2453 GND.n4165 GND.n4164 585
R2454 GND.n4215 GND.n4165 585
R2455 GND.n4218 GND.n4217 585
R2456 GND.n4217 GND.n4216 585
R2457 GND.n4219 GND.n4159 585
R2458 GND.n4159 GND.n4158 585
R2459 GND.n4221 GND.n4220 585
R2460 GND.n4222 GND.n4221 585
R2461 GND.n4157 GND.n4156 585
R2462 GND.n4223 GND.n4157 585
R2463 GND.n4226 GND.n4225 585
R2464 GND.n4225 GND.n4224 585
R2465 GND.n4227 GND.n4151 585
R2466 GND.n4151 GND.n4150 585
R2467 GND.n4229 GND.n4228 585
R2468 GND.n4230 GND.n4229 585
R2469 GND.n4149 GND.n4148 585
R2470 GND.n4231 GND.n4149 585
R2471 GND.n4234 GND.n4233 585
R2472 GND.n4233 GND.n4232 585
R2473 GND.n4235 GND.n4143 585
R2474 GND.n4143 GND.n4142 585
R2475 GND.n4237 GND.n4236 585
R2476 GND.n4238 GND.n4237 585
R2477 GND.n4141 GND.n4140 585
R2478 GND.n4239 GND.n4141 585
R2479 GND.n4242 GND.n4241 585
R2480 GND.n4241 GND.n4240 585
R2481 GND.n4243 GND.n4135 585
R2482 GND.n4135 GND.n4134 585
R2483 GND.n4245 GND.n4244 585
R2484 GND.n4246 GND.n4245 585
R2485 GND.n4133 GND.n4132 585
R2486 GND.n4247 GND.n4133 585
R2487 GND.n4250 GND.n4249 585
R2488 GND.n4249 GND.n4248 585
R2489 GND.n4251 GND.n4127 585
R2490 GND.n4127 GND.n4126 585
R2491 GND.n4253 GND.n4252 585
R2492 GND.n4254 GND.n4253 585
R2493 GND.n4125 GND.n4124 585
R2494 GND.n4255 GND.n4125 585
R2495 GND.n4258 GND.n4257 585
R2496 GND.n4257 GND.n4256 585
R2497 GND.n4259 GND.n4119 585
R2498 GND.n4119 GND.n4118 585
R2499 GND.n4261 GND.n4260 585
R2500 GND.n4262 GND.n4261 585
R2501 GND.n4117 GND.n4116 585
R2502 GND.n4263 GND.n4117 585
R2503 GND.n4266 GND.n4265 585
R2504 GND.n4265 GND.n4264 585
R2505 GND.n4267 GND.n4111 585
R2506 GND.n4111 GND.n4110 585
R2507 GND.n4269 GND.n4268 585
R2508 GND.n4270 GND.n4269 585
R2509 GND.n4109 GND.n4108 585
R2510 GND.n4271 GND.n4109 585
R2511 GND.n4274 GND.n4273 585
R2512 GND.n4273 GND.n4272 585
R2513 GND.n4275 GND.n4103 585
R2514 GND.n4103 GND.n4102 585
R2515 GND.n4277 GND.n4276 585
R2516 GND.n4278 GND.n4277 585
R2517 GND.n4101 GND.n4100 585
R2518 GND.n4279 GND.n4101 585
R2519 GND.n4282 GND.n4281 585
R2520 GND.n4281 GND.n4280 585
R2521 GND.n4283 GND.n4095 585
R2522 GND.n4095 GND.n4094 585
R2523 GND.n4285 GND.n4284 585
R2524 GND.n4286 GND.n4285 585
R2525 GND.n4093 GND.n4092 585
R2526 GND.n4287 GND.n4093 585
R2527 GND.n4290 GND.n4289 585
R2528 GND.n4289 GND.n4288 585
R2529 GND.n4291 GND.n4088 585
R2530 GND.n4088 GND.n4087 585
R2531 GND.n4293 GND.n4292 585
R2532 GND.n4294 GND.n4293 585
R2533 GND.n4086 GND.n4085 585
R2534 GND.n4295 GND.n4086 585
R2535 GND.n4298 GND.n4297 585
R2536 GND.n4297 GND.n4296 585
R2537 GND.n4082 GND.n4080 585
R2538 GND.n4080 GND.n4079 585
R2539 GND.n4303 GND.n4302 585
R2540 GND.n4304 GND.n4303 585
R2541 GND.n4081 GND.n4078 585
R2542 GND.n4305 GND.n4078 585
R2543 GND.n1739 GND.n1733 585
R2544 GND.n5691 GND.n1739 585
R2545 GND.n5542 GND.n5541 585
R2546 GND.n5541 GND.n1737 585
R2547 GND.n5543 GND.n2240 585
R2548 GND.n5559 GND.n2240 585
R2549 GND.n5540 GND.n5539 585
R2550 GND.n5539 GND.n2239 585
R2551 GND.n5538 GND.n2250 585
R2552 GND.n5550 GND.n2250 585
R2553 GND.n5537 GND.n5536 585
R2554 GND.n5536 GND.n2248 585
R2555 GND.n5535 GND.n2257 585
R2556 GND.n5535 GND.n5534 585
R2557 GND.n5519 GND.n2258 585
R2558 GND.n2270 GND.n2258 585
R2559 GND.n5518 GND.n2269 585
R2560 GND.n5526 GND.n2269 585
R2561 GND.n5517 GND.n5516 585
R2562 GND.n5516 GND.n2267 585
R2563 GND.n5515 GND.n2277 585
R2564 GND.n5515 GND.n5514 585
R2565 GND.n5499 GND.n2278 585
R2566 GND.n2279 GND.n2278 585
R2567 GND.n5498 GND.n2290 585
R2568 GND.n5506 GND.n2290 585
R2569 GND.n5497 GND.n5496 585
R2570 GND.n5496 GND.n2288 585
R2571 GND.n5495 GND.n2297 585
R2572 GND.n5495 GND.n5494 585
R2573 GND.n5479 GND.n2298 585
R2574 GND.n2299 GND.n2298 585
R2575 GND.n5478 GND.n2310 585
R2576 GND.n5486 GND.n2310 585
R2577 GND.n5477 GND.n5476 585
R2578 GND.n5476 GND.n2308 585
R2579 GND.n5475 GND.n2317 585
R2580 GND.n5475 GND.n5474 585
R2581 GND.n5459 GND.n2318 585
R2582 GND.n2319 GND.n2318 585
R2583 GND.n5458 GND.n2329 585
R2584 GND.n5466 GND.n2329 585
R2585 GND.n5457 GND.n5456 585
R2586 GND.n5456 GND.n5455 585
R2587 GND.n2337 GND.n2336 585
R2588 GND.n2338 GND.n2337 585
R2589 GND.n5376 GND.n2347 585
R2590 GND.n5396 GND.n2347 585
R2591 GND.n5375 GND.n5374 585
R2592 GND.n5374 GND.n2345 585
R2593 GND.n5373 GND.n2357 585
R2594 GND.n5386 GND.n2357 585
R2595 GND.n5372 GND.n5371 585
R2596 GND.n5371 GND.n2355 585
R2597 GND.n5370 GND.n2364 585
R2598 GND.n5370 GND.n5369 585
R2599 GND.n5354 GND.n2365 585
R2600 GND.n2366 GND.n2365 585
R2601 GND.n5353 GND.n2377 585
R2602 GND.n5361 GND.n2377 585
R2603 GND.n5352 GND.n5351 585
R2604 GND.n5351 GND.n2375 585
R2605 GND.n5350 GND.n2384 585
R2606 GND.n5350 GND.n5349 585
R2607 GND.n5334 GND.n2385 585
R2608 GND.n2397 GND.n2385 585
R2609 GND.n5333 GND.n2396 585
R2610 GND.n5341 GND.n2396 585
R2611 GND.n5332 GND.n5331 585
R2612 GND.n5331 GND.n2394 585
R2613 GND.n5330 GND.n2404 585
R2614 GND.n5330 GND.n5329 585
R2615 GND.n5314 GND.n2405 585
R2616 GND.n2406 GND.n2405 585
R2617 GND.n5313 GND.n2417 585
R2618 GND.n5321 GND.n2417 585
R2619 GND.n5312 GND.n5311 585
R2620 GND.n5311 GND.n2415 585
R2621 GND.n5310 GND.n2424 585
R2622 GND.n5310 GND.n5309 585
R2623 GND.n5294 GND.n2425 585
R2624 GND.n2426 GND.n2425 585
R2625 GND.n5293 GND.n2437 585
R2626 GND.n5301 GND.n2437 585
R2627 GND.n5292 GND.n5291 585
R2628 GND.n5291 GND.n2435 585
R2629 GND.n5290 GND.n2444 585
R2630 GND.n5290 GND.n5289 585
R2631 GND.n5274 GND.n2445 585
R2632 GND.n2457 GND.n2445 585
R2633 GND.n5273 GND.n2456 585
R2634 GND.n5281 GND.n2456 585
R2635 GND.n5272 GND.n5271 585
R2636 GND.n5271 GND.n2454 585
R2637 GND.n5270 GND.n2464 585
R2638 GND.n5270 GND.n5269 585
R2639 GND.n5254 GND.n2465 585
R2640 GND.n2466 GND.n2465 585
R2641 GND.n5253 GND.n2477 585
R2642 GND.n5261 GND.n2477 585
R2643 GND.n5252 GND.n5251 585
R2644 GND.n5251 GND.n2475 585
R2645 GND.n5250 GND.n2484 585
R2646 GND.n5250 GND.n5249 585
R2647 GND.n5234 GND.n2485 585
R2648 GND.n2486 GND.n2485 585
R2649 GND.n5233 GND.n2497 585
R2650 GND.n5241 GND.n2497 585
R2651 GND.n5232 GND.n5231 585
R2652 GND.n5231 GND.n2495 585
R2653 GND.n5230 GND.n2504 585
R2654 GND.n5230 GND.n5229 585
R2655 GND.n5185 GND.n2505 585
R2656 GND.n2506 GND.n2505 585
R2657 GND.n5184 GND.n5183 585
R2658 GND.n5183 GND.n5182 585
R2659 GND.n2576 GND.n2575 585
R2660 GND.n2577 GND.n2576 585
R2661 GND.n2720 GND.n2568 585
R2662 GND.n5175 GND.n2720 585
R2663 GND.n2732 GND.n2567 585
R2664 GND.n2732 GND.n2715 585
R2665 GND.n2733 GND.n2566 585
R2666 GND.n5082 GND.n2733 585
R2667 GND.n2748 GND.n2747 585
R2668 GND.n2748 GND.n2727 585
R2669 GND.n2749 GND.n2560 585
R2670 GND.n5075 GND.n2749 585
R2671 GND.n2746 GND.n2559 585
R2672 GND.n2746 GND.n2737 585
R2673 GND.n2745 GND.n2558 585
R2674 GND.n2745 GND.n2530 585
R2675 GND.n2557 GND.n2529 585
R2676 GND.n5220 GND.n2529 585
R2677 GND.n2756 GND.n2552 585
R2678 GND.n2757 GND.n2756 585
R2679 GND.n2755 GND.n2551 585
R2680 GND.n2755 GND.n2543 585
R2681 GND.n2550 GND.n2542 585
R2682 GND.n5210 GND.n2542 585
R2683 GND.n5042 GND.n5041 585
R2684 GND.n5041 GND.n2540 585
R2685 GND.n5043 GND.n2764 585
R2686 GND.n5058 GND.n2764 585
R2687 GND.n5040 GND.n5039 585
R2688 GND.n5039 GND.n2762 585
R2689 GND.n5038 GND.n2773 585
R2690 GND.n5050 GND.n2773 585
R2691 GND.n5037 GND.n5036 585
R2692 GND.n5036 GND.n2771 585
R2693 GND.n5035 GND.n2780 585
R2694 GND.n5035 GND.n5034 585
R2695 GND.n1750 GND.n1730 585
R2696 GND.n1759 GND.n1758 585
R2697 GND.n1761 GND.n1760 585
R2698 GND.n1763 GND.n1762 585
R2699 GND.n1765 GND.n1764 585
R2700 GND.n1767 GND.n1766 585
R2701 GND.n1769 GND.n1768 585
R2702 GND.n1771 GND.n1770 585
R2703 GND.n1773 GND.n1772 585
R2704 GND.n1775 GND.n1774 585
R2705 GND.n1777 GND.n1776 585
R2706 GND.n5422 GND.n1741 585
R2707 GND.n5691 GND.n1741 585
R2708 GND.n5424 GND.n5423 585
R2709 GND.n5423 GND.n1737 585
R2710 GND.n5425 GND.n2241 585
R2711 GND.n5559 GND.n2241 585
R2712 GND.n5427 GND.n5426 585
R2713 GND.n5426 GND.n2239 585
R2714 GND.n5428 GND.n2251 585
R2715 GND.n5550 GND.n2251 585
R2716 GND.n5430 GND.n5429 585
R2717 GND.n5429 GND.n2248 585
R2718 GND.n5431 GND.n2260 585
R2719 GND.n5534 GND.n2260 585
R2720 GND.n5433 GND.n5432 585
R2721 GND.n5432 GND.n2270 585
R2722 GND.n5434 GND.n2271 585
R2723 GND.n5526 GND.n2271 585
R2724 GND.n5436 GND.n5435 585
R2725 GND.n5435 GND.n2267 585
R2726 GND.n5437 GND.n2281 585
R2727 GND.n5514 GND.n2281 585
R2728 GND.n5439 GND.n5438 585
R2729 GND.n5438 GND.n2279 585
R2730 GND.n5440 GND.n2291 585
R2731 GND.n5506 GND.n2291 585
R2732 GND.n5442 GND.n5441 585
R2733 GND.n5441 GND.n2288 585
R2734 GND.n5443 GND.n2301 585
R2735 GND.n5494 GND.n2301 585
R2736 GND.n5445 GND.n5444 585
R2737 GND.n5444 GND.n2299 585
R2738 GND.n5446 GND.n2311 585
R2739 GND.n5486 GND.n2311 585
R2740 GND.n5448 GND.n5447 585
R2741 GND.n5447 GND.n2308 585
R2742 GND.n5449 GND.n2321 585
R2743 GND.n5474 GND.n2321 585
R2744 GND.n5451 GND.n5450 585
R2745 GND.n5450 GND.n2319 585
R2746 GND.n5452 GND.n2330 585
R2747 GND.n5466 GND.n2330 585
R2748 GND.n5454 GND.n5453 585
R2749 GND.n5455 GND.n5454 585
R2750 GND.n2341 GND.n2340 585
R2751 GND.n2340 GND.n2338 585
R2752 GND.n5398 GND.n5397 585
R2753 GND.n5397 GND.n5396 585
R2754 GND.n2344 GND.n2343 585
R2755 GND.n2345 GND.n2344 585
R2756 GND.n5123 GND.n2358 585
R2757 GND.n5386 GND.n2358 585
R2758 GND.n5125 GND.n5124 585
R2759 GND.n5124 GND.n2355 585
R2760 GND.n5126 GND.n2368 585
R2761 GND.n5369 GND.n2368 585
R2762 GND.n5128 GND.n5127 585
R2763 GND.n5127 GND.n2366 585
R2764 GND.n5129 GND.n2378 585
R2765 GND.n5361 GND.n2378 585
R2766 GND.n5131 GND.n5130 585
R2767 GND.n5130 GND.n2375 585
R2768 GND.n5132 GND.n2387 585
R2769 GND.n5349 GND.n2387 585
R2770 GND.n5134 GND.n5133 585
R2771 GND.n5133 GND.n2397 585
R2772 GND.n5135 GND.n2398 585
R2773 GND.n5341 GND.n2398 585
R2774 GND.n5137 GND.n5136 585
R2775 GND.n5136 GND.n2394 585
R2776 GND.n5138 GND.n2408 585
R2777 GND.n5329 GND.n2408 585
R2778 GND.n5140 GND.n5139 585
R2779 GND.n5139 GND.n2406 585
R2780 GND.n5141 GND.n2418 585
R2781 GND.n5321 GND.n2418 585
R2782 GND.n5143 GND.n5142 585
R2783 GND.n5142 GND.n2415 585
R2784 GND.n5144 GND.n2428 585
R2785 GND.n5309 GND.n2428 585
R2786 GND.n5146 GND.n5145 585
R2787 GND.n5145 GND.n2426 585
R2788 GND.n5147 GND.n2438 585
R2789 GND.n5301 GND.n2438 585
R2790 GND.n5149 GND.n5148 585
R2791 GND.n5148 GND.n2435 585
R2792 GND.n5150 GND.n2447 585
R2793 GND.n5289 GND.n2447 585
R2794 GND.n5152 GND.n5151 585
R2795 GND.n5151 GND.n2457 585
R2796 GND.n5153 GND.n2458 585
R2797 GND.n5281 GND.n2458 585
R2798 GND.n5155 GND.n5154 585
R2799 GND.n5154 GND.n2454 585
R2800 GND.n5156 GND.n2468 585
R2801 GND.n5269 GND.n2468 585
R2802 GND.n5158 GND.n5157 585
R2803 GND.n5157 GND.n2466 585
R2804 GND.n5159 GND.n2478 585
R2805 GND.n5261 GND.n2478 585
R2806 GND.n5161 GND.n5160 585
R2807 GND.n5160 GND.n2475 585
R2808 GND.n5162 GND.n2488 585
R2809 GND.n5249 GND.n2488 585
R2810 GND.n5164 GND.n5163 585
R2811 GND.n5163 GND.n2486 585
R2812 GND.n5165 GND.n2498 585
R2813 GND.n5241 GND.n2498 585
R2814 GND.n5167 GND.n5166 585
R2815 GND.n5166 GND.n2495 585
R2816 GND.n5168 GND.n2508 585
R2817 GND.n5229 GND.n2508 585
R2818 GND.n5170 GND.n5169 585
R2819 GND.n5169 GND.n2506 585
R2820 GND.n5171 GND.n2712 585
R2821 GND.n5182 GND.n2712 585
R2822 GND.n5172 GND.n2722 585
R2823 GND.n2722 GND.n2577 585
R2824 GND.n5174 GND.n5173 585
R2825 GND.n5175 GND.n5174 585
R2826 GND.n2723 GND.n2721 585
R2827 GND.n2721 GND.n2715 585
R2828 GND.n5084 GND.n5083 585
R2829 GND.n5083 GND.n5082 585
R2830 GND.n2726 GND.n2725 585
R2831 GND.n2727 GND.n2726 585
R2832 GND.n5074 GND.n5073 585
R2833 GND.n5075 GND.n5074 585
R2834 GND.n2751 GND.n2750 585
R2835 GND.n2750 GND.n2737 585
R2836 GND.n5069 GND.n5068 585
R2837 GND.n5068 GND.n2530 585
R2838 GND.n5067 GND.n2531 585
R2839 GND.n5220 GND.n2531 585
R2840 GND.n5066 GND.n2758 585
R2841 GND.n2758 GND.n2757 585
R2842 GND.n2754 GND.n2753 585
R2843 GND.n2754 GND.n2543 585
R2844 GND.n5062 GND.n2544 585
R2845 GND.n5210 GND.n2544 585
R2846 GND.n5061 GND.n5060 585
R2847 GND.n5060 GND.n2540 585
R2848 GND.n5059 GND.n2760 585
R2849 GND.n5059 GND.n5058 585
R2850 GND.n3258 GND.n2761 585
R2851 GND.n2762 GND.n2761 585
R2852 GND.n3259 GND.n2774 585
R2853 GND.n5050 GND.n2774 585
R2854 GND.n3255 GND.n3254 585
R2855 GND.n3254 GND.n2771 585
R2856 GND.n3263 GND.n2784 585
R2857 GND.n5034 GND.n2784 585
R2858 GND.n519 GND.n518 585
R2859 GND.n522 GND.n519 585
R2860 GND.n7472 GND.n7471 585
R2861 GND.n7471 GND.n7470 585
R2862 GND.n7473 GND.n514 585
R2863 GND.n514 GND.n513 585
R2864 GND.n7475 GND.n7474 585
R2865 GND.n7476 GND.n7475 585
R2866 GND.n499 GND.n498 585
R2867 GND.n503 GND.n499 585
R2868 GND.n7484 GND.n7483 585
R2869 GND.n7483 GND.n7482 585
R2870 GND.n7485 GND.n494 585
R2871 GND.n500 GND.n494 585
R2872 GND.n7487 GND.n7486 585
R2873 GND.n7488 GND.n7487 585
R2874 GND.n481 GND.n480 585
R2875 GND.n484 GND.n481 585
R2876 GND.n7496 GND.n7495 585
R2877 GND.n7495 GND.n7494 585
R2878 GND.n7497 GND.n476 585
R2879 GND.n476 GND.n475 585
R2880 GND.n7499 GND.n7498 585
R2881 GND.n7500 GND.n7499 585
R2882 GND.n462 GND.n461 585
R2883 GND.n465 GND.n462 585
R2884 GND.n7508 GND.n7507 585
R2885 GND.n7507 GND.n7506 585
R2886 GND.n7509 GND.n457 585
R2887 GND.n457 GND.n456 585
R2888 GND.n7511 GND.n7510 585
R2889 GND.n7512 GND.n7511 585
R2890 GND.n442 GND.n441 585
R2891 GND.n445 GND.n442 585
R2892 GND.n7520 GND.n7519 585
R2893 GND.n7519 GND.n7518 585
R2894 GND.n7521 GND.n437 585
R2895 GND.n437 GND.n436 585
R2896 GND.n7523 GND.n7522 585
R2897 GND.n7524 GND.n7523 585
R2898 GND.n423 GND.n422 585
R2899 GND.n433 GND.n423 585
R2900 GND.n7532 GND.n7531 585
R2901 GND.n7531 GND.n7530 585
R2902 GND.n7533 GND.n418 585
R2903 GND.n418 GND.n417 585
R2904 GND.n7535 GND.n7534 585
R2905 GND.n7536 GND.n7535 585
R2906 GND.n404 GND.n403 585
R2907 GND.n407 GND.n404 585
R2908 GND.n7544 GND.n7543 585
R2909 GND.n7543 GND.n7542 585
R2910 GND.n7545 GND.n399 585
R2911 GND.n399 GND.n398 585
R2912 GND.n7547 GND.n7546 585
R2913 GND.n7548 GND.n7547 585
R2914 GND.n385 GND.n384 585
R2915 GND.n388 GND.n385 585
R2916 GND.n7556 GND.n7555 585
R2917 GND.n7555 GND.n7554 585
R2918 GND.n7557 GND.n380 585
R2919 GND.n380 GND.n379 585
R2920 GND.n7559 GND.n7558 585
R2921 GND.n7560 GND.n7559 585
R2922 GND.n366 GND.n365 585
R2923 GND.n369 GND.n366 585
R2924 GND.n7568 GND.n7567 585
R2925 GND.n7567 GND.n7566 585
R2926 GND.n7569 GND.n361 585
R2927 GND.n361 GND.n360 585
R2928 GND.n7571 GND.n7570 585
R2929 GND.n7572 GND.n7571 585
R2930 GND.n347 GND.n346 585
R2931 GND.n350 GND.n347 585
R2932 GND.n7580 GND.n7579 585
R2933 GND.n7579 GND.n7578 585
R2934 GND.n7581 GND.n342 585
R2935 GND.n342 GND.n341 585
R2936 GND.n7583 GND.n7582 585
R2937 GND.n7584 GND.n7583 585
R2938 GND.n328 GND.n327 585
R2939 GND.n331 GND.n328 585
R2940 GND.n7592 GND.n7591 585
R2941 GND.n7591 GND.n7590 585
R2942 GND.n7593 GND.n321 585
R2943 GND.n321 GND.n319 585
R2944 GND.n7595 GND.n7594 585
R2945 GND.n7596 GND.n7595 585
R2946 GND.n322 GND.n320 585
R2947 GND.n7234 GND.n320 585
R2948 GND.n7183 GND.n308 585
R2949 GND.n7602 GND.n308 585
R2950 GND.n7185 GND.n7184 585
R2951 GND.n7184 GND.n298 585
R2952 GND.n7186 GND.n297 585
R2953 GND.n7608 GND.n297 585
R2954 GND.n7188 GND.n7187 585
R2955 GND.n7187 GND.n287 585
R2956 GND.n7189 GND.n286 585
R2957 GND.n7614 GND.n286 585
R2958 GND.n7191 GND.n7190 585
R2959 GND.n7190 GND.n277 585
R2960 GND.n7192 GND.n276 585
R2961 GND.n7620 GND.n276 585
R2962 GND.n7194 GND.n7193 585
R2963 GND.n7193 GND.n267 585
R2964 GND.n7195 GND.n266 585
R2965 GND.n7626 GND.n266 585
R2966 GND.n7197 GND.n7196 585
R2967 GND.n7196 GND.n264 585
R2968 GND.n7198 GND.n254 585
R2969 GND.n7632 GND.n254 585
R2970 GND.n7200 GND.n7199 585
R2971 GND.n7199 GND.n252 585
R2972 GND.n7180 GND.n621 585
R2973 GND.n7208 GND.n621 585
R2974 GND.n7179 GND.n7178 585
R2975 GND.n7178 GND.n619 585
R2976 GND.n7177 GND.n7176 585
R2977 GND.n7177 GND.n236 585
R2978 GND.n625 GND.n235 585
R2979 GND.n7641 GND.n235 585
R2980 GND.n7153 GND.n7152 585
R2981 GND.n7152 GND.n233 585
R2982 GND.n7154 GND.n632 585
R2983 GND.n7168 GND.n632 585
R2984 GND.n7151 GND.n7150 585
R2985 GND.n7150 GND.n630 585
R2986 GND.n7149 GND.n637 585
R2987 GND.n7160 GND.n637 585
R2988 GND.n7148 GND.n7147 585
R2989 GND.n7147 GND.n635 585
R2990 GND.n7146 GND.n642 585
R2991 GND.n7146 GND.n7145 585
R2992 GND.n7087 GND.n644 585
R2993 GND.n7129 GND.n644 585
R2994 GND.n7089 GND.n7088 585
R2995 GND.n7088 GND.n657 585
R2996 GND.n7090 GND.n656 585
R2997 GND.n7135 GND.n656 585
R2998 GND.n7092 GND.n7091 585
R2999 GND.n7091 GND.n654 585
R3000 GND.n7086 GND.n675 585
R3001 GND.n7107 GND.n675 585
R3002 GND.n7085 GND.n7084 585
R3003 GND.n7084 GND.n673 585
R3004 GND.n7083 GND.n684 585
R3005 GND.n7099 GND.n684 585
R3006 GND.n7082 GND.n7081 585
R3007 GND.n7081 GND.n682 585
R3008 GND.n7080 GND.n691 585
R3009 GND.n7080 GND.n7079 585
R3010 GND.n7064 GND.n693 585
R3011 GND.n694 GND.n693 585
R3012 GND.n7063 GND.n704 585
R3013 GND.n7071 GND.n704 585
R3014 GND.n7062 GND.n7061 585
R3015 GND.n7061 GND.n7060 585
R3016 GND.n712 GND.n710 585
R3017 GND.n713 GND.n712 585
R3018 GND.n7018 GND.n722 585
R3019 GND.n7037 GND.n722 585
R3020 GND.n7017 GND.n7016 585
R3021 GND.n7016 GND.n720 585
R3022 GND.n7015 GND.n732 585
R3023 GND.n7027 GND.n732 585
R3024 GND.n7014 GND.n7013 585
R3025 GND.n7013 GND.n730 585
R3026 GND.n7012 GND.n739 585
R3027 GND.n7012 GND.n7011 585
R3028 GND.n6996 GND.n741 585
R3029 GND.n742 GND.n741 585
R3030 GND.n6995 GND.n753 585
R3031 GND.n7003 GND.n753 585
R3032 GND.n6994 GND.n6993 585
R3033 GND.n6993 GND.n751 585
R3034 GND.n6992 GND.n759 585
R3035 GND.n6992 GND.n6991 585
R3036 GND.n6976 GND.n761 585
R3037 GND.n762 GND.n761 585
R3038 GND.n6975 GND.n773 585
R3039 GND.n6983 GND.n773 585
R3040 GND.n6974 GND.n6973 585
R3041 GND.n6973 GND.n771 585
R3042 GND.n6972 GND.n779 585
R3043 GND.n6972 GND.n6971 585
R3044 GND.n6956 GND.n781 585
R3045 GND.n782 GND.n781 585
R3046 GND.n6955 GND.n793 585
R3047 GND.n6963 GND.n793 585
R3048 GND.n6954 GND.n6953 585
R3049 GND.n6953 GND.n791 585
R3050 GND.n6952 GND.n799 585
R3051 GND.n6952 GND.n6951 585
R3052 GND.n6936 GND.n801 585
R3053 GND.n802 GND.n801 585
R3054 GND.n6935 GND.n813 585
R3055 GND.n6943 GND.n813 585
R3056 GND.n6934 GND.n6933 585
R3057 GND.n6933 GND.n811 585
R3058 GND.n6932 GND.n819 585
R3059 GND.n6932 GND.n6931 585
R3060 GND.n6916 GND.n821 585
R3061 GND.n833 GND.n821 585
R3062 GND.n6915 GND.n832 585
R3063 GND.n6923 GND.n832 585
R3064 GND.n6914 GND.n6913 585
R3065 GND.n6913 GND.n830 585
R3066 GND.n6912 GND.n839 585
R3067 GND.n6912 GND.n6911 585
R3068 GND.n6896 GND.n841 585
R3069 GND.n842 GND.n841 585
R3070 GND.n6895 GND.n853 585
R3071 GND.n6903 GND.n853 585
R3072 GND.n6894 GND.n6893 585
R3073 GND.n6893 GND.n851 585
R3074 GND.n6892 GND.n859 585
R3075 GND.n6892 GND.n6891 585
R3076 GND.n6876 GND.n861 585
R3077 GND.n862 GND.n861 585
R3078 GND.n6875 GND.n873 585
R3079 GND.n6883 GND.n873 585
R3080 GND.n6874 GND.n6873 585
R3081 GND.n6873 GND.n871 585
R3082 GND.n6872 GND.n879 585
R3083 GND.n6872 GND.n6871 585
R3084 GND.n6856 GND.n881 585
R3085 GND.n882 GND.n881 585
R3086 GND.n6855 GND.n892 585
R3087 GND.n6863 GND.n892 585
R3088 GND.n6854 GND.n6853 585
R3089 GND.n6853 GND.n6852 585
R3090 GND.n900 GND.n898 585
R3091 GND.n901 GND.n900 585
R3092 GND.n6743 GND.n910 585
R3093 GND.n6762 GND.n910 585
R3094 GND.n6742 GND.n6741 585
R3095 GND.n6741 GND.n908 585
R3096 GND.n6740 GND.n920 585
R3097 GND.n6752 GND.n920 585
R3098 GND.n6739 GND.n928 585
R3099 GND.n928 GND.n918 585
R3100 GND.n933 GND.n927 585
R3101 GND.n6734 GND.n933 585
R3102 GND.n1348 GND.n1347 585
R3103 GND.n1350 GND.n1349 585
R3104 GND.n1353 GND.n1352 585
R3105 GND.n1355 GND.n1354 585
R3106 GND.n1358 GND.n1357 585
R3107 GND.n1360 GND.n1359 585
R3108 GND.n1366 GND.n1365 585
R3109 GND.n1368 GND.n1367 585
R3110 GND.n1369 GND.n1362 585
R3111 GND.n6725 GND.n950 585
R3112 GND.n7327 GND.n7326 585
R3113 GND.n7329 GND.n582 585
R3114 GND.n7331 GND.n7330 585
R3115 GND.n7332 GND.n575 585
R3116 GND.n7334 GND.n7333 585
R3117 GND.n7336 GND.n573 585
R3118 GND.n7338 GND.n7337 585
R3119 GND.n7339 GND.n569 585
R3120 GND.n7341 GND.n7340 585
R3121 GND.n7343 GND.n568 585
R3122 GND.n7345 GND.n7344 585
R3123 GND.n7344 GND.n528 585
R3124 GND.n7323 GND.n584 585
R3125 GND.n584 GND.n522 585
R3126 GND.n7322 GND.n521 585
R3127 GND.n7470 GND.n521 585
R3128 GND.n7321 GND.n7320 585
R3129 GND.n7320 GND.n513 585
R3130 GND.n587 GND.n512 585
R3131 GND.n7476 GND.n512 585
R3132 GND.n7316 GND.n7315 585
R3133 GND.n7315 GND.n503 585
R3134 GND.n7314 GND.n502 585
R3135 GND.n7482 GND.n502 585
R3136 GND.n7313 GND.n7312 585
R3137 GND.n7312 GND.n500 585
R3138 GND.n589 GND.n493 585
R3139 GND.n7488 GND.n493 585
R3140 GND.n7308 GND.n7307 585
R3141 GND.n7307 GND.n484 585
R3142 GND.n7306 GND.n483 585
R3143 GND.n7494 GND.n483 585
R3144 GND.n7305 GND.n7304 585
R3145 GND.n7304 GND.n475 585
R3146 GND.n591 GND.n474 585
R3147 GND.n7500 GND.n474 585
R3148 GND.n7300 GND.n7299 585
R3149 GND.n7299 GND.n465 585
R3150 GND.n7298 GND.n464 585
R3151 GND.n7506 GND.n464 585
R3152 GND.n7297 GND.n7296 585
R3153 GND.n7296 GND.n456 585
R3154 GND.n593 GND.n455 585
R3155 GND.n7512 GND.n455 585
R3156 GND.n7292 GND.n7291 585
R3157 GND.n7291 GND.n445 585
R3158 GND.n7290 GND.n444 585
R3159 GND.n7518 GND.n444 585
R3160 GND.n7289 GND.n7288 585
R3161 GND.n7288 GND.n436 585
R3162 GND.n595 GND.n435 585
R3163 GND.n7524 GND.n435 585
R3164 GND.n7284 GND.n7283 585
R3165 GND.n7283 GND.n433 585
R3166 GND.n7282 GND.n425 585
R3167 GND.n7530 GND.n425 585
R3168 GND.n7281 GND.n7280 585
R3169 GND.n7280 GND.n417 585
R3170 GND.n597 GND.n416 585
R3171 GND.n7536 GND.n416 585
R3172 GND.n7276 GND.n7275 585
R3173 GND.n7275 GND.n407 585
R3174 GND.n7274 GND.n406 585
R3175 GND.n7542 GND.n406 585
R3176 GND.n7273 GND.n7272 585
R3177 GND.n7272 GND.n398 585
R3178 GND.n599 GND.n397 585
R3179 GND.n7548 GND.n397 585
R3180 GND.n7268 GND.n7267 585
R3181 GND.n7267 GND.n388 585
R3182 GND.n7266 GND.n387 585
R3183 GND.n7554 GND.n387 585
R3184 GND.n7265 GND.n7264 585
R3185 GND.n7264 GND.n379 585
R3186 GND.n601 GND.n378 585
R3187 GND.n7560 GND.n378 585
R3188 GND.n7260 GND.n7259 585
R3189 GND.n7259 GND.n369 585
R3190 GND.n7258 GND.n368 585
R3191 GND.n7566 GND.n368 585
R3192 GND.n7257 GND.n7256 585
R3193 GND.n7256 GND.n360 585
R3194 GND.n603 GND.n359 585
R3195 GND.n7572 GND.n359 585
R3196 GND.n7252 GND.n7251 585
R3197 GND.n7251 GND.n350 585
R3198 GND.n7250 GND.n349 585
R3199 GND.n7578 GND.n349 585
R3200 GND.n7249 GND.n7248 585
R3201 GND.n7248 GND.n341 585
R3202 GND.n605 GND.n340 585
R3203 GND.n7584 GND.n340 585
R3204 GND.n7244 GND.n7243 585
R3205 GND.n7243 GND.n331 585
R3206 GND.n7242 GND.n330 585
R3207 GND.n7590 GND.n330 585
R3208 GND.n7241 GND.n7240 585
R3209 GND.n7240 GND.n319 585
R3210 GND.n607 GND.n318 585
R3211 GND.n7596 GND.n318 585
R3212 GND.n7236 GND.n7235 585
R3213 GND.n7235 GND.n7234 585
R3214 GND.n7233 GND.n306 585
R3215 GND.n7602 GND.n306 585
R3216 GND.n7232 GND.n7231 585
R3217 GND.n7231 GND.n298 585
R3218 GND.n609 GND.n299 585
R3219 GND.n7608 GND.n299 585
R3220 GND.n7227 GND.n7226 585
R3221 GND.n7226 GND.n287 585
R3222 GND.n7225 GND.n288 585
R3223 GND.n7614 GND.n288 585
R3224 GND.n7224 GND.n7223 585
R3225 GND.n7223 GND.n277 585
R3226 GND.n611 GND.n278 585
R3227 GND.n7620 GND.n278 585
R3228 GND.n7219 GND.n7218 585
R3229 GND.n7218 GND.n267 585
R3230 GND.n7217 GND.n268 585
R3231 GND.n7626 GND.n268 585
R3232 GND.n7216 GND.n7215 585
R3233 GND.n7215 GND.n264 585
R3234 GND.n613 GND.n255 585
R3235 GND.n7632 GND.n255 585
R3236 GND.n7211 GND.n7210 585
R3237 GND.n7210 GND.n252 585
R3238 GND.n7209 GND.n615 585
R3239 GND.n7209 GND.n7208 585
R3240 GND.n618 GND.n617 585
R3241 GND.n619 GND.n618 585
R3242 GND.n232 GND.n230 585
R3243 GND.n236 GND.n232 585
R3244 GND.n7643 GND.n7642 585
R3245 GND.n7642 GND.n7641 585
R3246 GND.n231 GND.n229 585
R3247 GND.n233 GND.n231 585
R3248 GND.n7120 GND.n633 585
R3249 GND.n7168 GND.n633 585
R3250 GND.n7122 GND.n7121 585
R3251 GND.n7121 GND.n630 585
R3252 GND.n7123 GND.n638 585
R3253 GND.n7160 GND.n638 585
R3254 GND.n7125 GND.n7124 585
R3255 GND.n7124 GND.n635 585
R3256 GND.n7126 GND.n646 585
R3257 GND.n7145 GND.n646 585
R3258 GND.n7128 GND.n7127 585
R3259 GND.n7129 GND.n7128 585
R3260 GND.n669 GND.n668 585
R3261 GND.n668 GND.n657 585
R3262 GND.n7111 GND.n658 585
R3263 GND.n7135 GND.n658 585
R3264 GND.n7110 GND.n7109 585
R3265 GND.n7109 GND.n654 585
R3266 GND.n7108 GND.n671 585
R3267 GND.n7108 GND.n7107 585
R3268 GND.n7050 GND.n672 585
R3269 GND.n673 GND.n672 585
R3270 GND.n7051 GND.n685 585
R3271 GND.n7099 GND.n685 585
R3272 GND.n7053 GND.n7052 585
R3273 GND.n7052 GND.n682 585
R3274 GND.n7054 GND.n696 585
R3275 GND.n7079 GND.n696 585
R3276 GND.n7056 GND.n7055 585
R3277 GND.n7055 GND.n694 585
R3278 GND.n7057 GND.n705 585
R3279 GND.n7071 GND.n705 585
R3280 GND.n7059 GND.n7058 585
R3281 GND.n7060 GND.n7059 585
R3282 GND.n716 GND.n715 585
R3283 GND.n715 GND.n713 585
R3284 GND.n7039 GND.n7038 585
R3285 GND.n7038 GND.n7037 585
R3286 GND.n719 GND.n718 585
R3287 GND.n720 GND.n719 585
R3288 GND.n6801 GND.n733 585
R3289 GND.n7027 GND.n733 585
R3290 GND.n6803 GND.n6802 585
R3291 GND.n6802 GND.n730 585
R3292 GND.n6804 GND.n744 585
R3293 GND.n7011 GND.n744 585
R3294 GND.n6806 GND.n6805 585
R3295 GND.n6805 GND.n742 585
R3296 GND.n6807 GND.n754 585
R3297 GND.n7003 GND.n754 585
R3298 GND.n6809 GND.n6808 585
R3299 GND.n6808 GND.n751 585
R3300 GND.n6810 GND.n764 585
R3301 GND.n6991 GND.n764 585
R3302 GND.n6812 GND.n6811 585
R3303 GND.n6811 GND.n762 585
R3304 GND.n6813 GND.n774 585
R3305 GND.n6983 GND.n774 585
R3306 GND.n6815 GND.n6814 585
R3307 GND.n6814 GND.n771 585
R3308 GND.n6816 GND.n784 585
R3309 GND.n6971 GND.n784 585
R3310 GND.n6818 GND.n6817 585
R3311 GND.n6817 GND.n782 585
R3312 GND.n6819 GND.n794 585
R3313 GND.n6963 GND.n794 585
R3314 GND.n6821 GND.n6820 585
R3315 GND.n6820 GND.n791 585
R3316 GND.n6822 GND.n804 585
R3317 GND.n6951 GND.n804 585
R3318 GND.n6824 GND.n6823 585
R3319 GND.n6823 GND.n802 585
R3320 GND.n6825 GND.n814 585
R3321 GND.n6943 GND.n814 585
R3322 GND.n6827 GND.n6826 585
R3323 GND.n6826 GND.n811 585
R3324 GND.n6828 GND.n823 585
R3325 GND.n6931 GND.n823 585
R3326 GND.n6830 GND.n6829 585
R3327 GND.n6829 GND.n833 585
R3328 GND.n6831 GND.n834 585
R3329 GND.n6923 GND.n834 585
R3330 GND.n6833 GND.n6832 585
R3331 GND.n6832 GND.n830 585
R3332 GND.n6834 GND.n844 585
R3333 GND.n6911 GND.n844 585
R3334 GND.n6836 GND.n6835 585
R3335 GND.n6835 GND.n842 585
R3336 GND.n6837 GND.n854 585
R3337 GND.n6903 GND.n854 585
R3338 GND.n6839 GND.n6838 585
R3339 GND.n6838 GND.n851 585
R3340 GND.n6840 GND.n864 585
R3341 GND.n6891 GND.n864 585
R3342 GND.n6842 GND.n6841 585
R3343 GND.n6841 GND.n862 585
R3344 GND.n6843 GND.n874 585
R3345 GND.n6883 GND.n874 585
R3346 GND.n6845 GND.n6844 585
R3347 GND.n6844 GND.n871 585
R3348 GND.n6846 GND.n884 585
R3349 GND.n6871 GND.n884 585
R3350 GND.n6848 GND.n6847 585
R3351 GND.n6847 GND.n882 585
R3352 GND.n6849 GND.n893 585
R3353 GND.n6863 GND.n893 585
R3354 GND.n6851 GND.n6850 585
R3355 GND.n6852 GND.n6851 585
R3356 GND.n904 GND.n903 585
R3357 GND.n903 GND.n901 585
R3358 GND.n6764 GND.n6763 585
R3359 GND.n6763 GND.n6762 585
R3360 GND.n907 GND.n906 585
R3361 GND.n908 GND.n907 585
R3362 GND.n1374 GND.n921 585
R3363 GND.n6752 GND.n921 585
R3364 GND.n1375 GND.n1372 585
R3365 GND.n1372 GND.n918 585
R3366 GND.n1376 GND.n934 585
R3367 GND.n6734 GND.n934 585
R3368 GND.n5563 GND.n1738 585
R3369 GND.n5691 GND.n1738 585
R3370 GND.n5562 GND.n5561 585
R3371 GND.n5561 GND.n1737 585
R3372 GND.n5560 GND.n2237 585
R3373 GND.n5560 GND.n5559 585
R3374 GND.n2631 GND.n2238 585
R3375 GND.n2239 GND.n2238 585
R3376 GND.n2632 GND.n2249 585
R3377 GND.n5550 GND.n2249 585
R3378 GND.n2634 GND.n2633 585
R3379 GND.n2633 GND.n2248 585
R3380 GND.n2635 GND.n2259 585
R3381 GND.n5534 GND.n2259 585
R3382 GND.n2637 GND.n2636 585
R3383 GND.n2636 GND.n2270 585
R3384 GND.n2638 GND.n2268 585
R3385 GND.n5526 GND.n2268 585
R3386 GND.n2640 GND.n2639 585
R3387 GND.n2639 GND.n2267 585
R3388 GND.n2641 GND.n2280 585
R3389 GND.n5514 GND.n2280 585
R3390 GND.n2643 GND.n2642 585
R3391 GND.n2642 GND.n2279 585
R3392 GND.n2644 GND.n2289 585
R3393 GND.n5506 GND.n2289 585
R3394 GND.n2646 GND.n2645 585
R3395 GND.n2645 GND.n2288 585
R3396 GND.n2647 GND.n2300 585
R3397 GND.n5494 GND.n2300 585
R3398 GND.n2649 GND.n2648 585
R3399 GND.n2648 GND.n2299 585
R3400 GND.n2650 GND.n2309 585
R3401 GND.n5486 GND.n2309 585
R3402 GND.n2652 GND.n2651 585
R3403 GND.n2651 GND.n2308 585
R3404 GND.n2653 GND.n2320 585
R3405 GND.n5474 GND.n2320 585
R3406 GND.n2655 GND.n2654 585
R3407 GND.n2654 GND.n2319 585
R3408 GND.n2656 GND.n2328 585
R3409 GND.n5466 GND.n2328 585
R3410 GND.n2657 GND.n2339 585
R3411 GND.n5455 GND.n2339 585
R3412 GND.n2659 GND.n2658 585
R3413 GND.n2658 GND.n2338 585
R3414 GND.n2660 GND.n2346 585
R3415 GND.n5396 GND.n2346 585
R3416 GND.n2662 GND.n2661 585
R3417 GND.n2661 GND.n2345 585
R3418 GND.n2663 GND.n2356 585
R3419 GND.n5386 GND.n2356 585
R3420 GND.n2665 GND.n2664 585
R3421 GND.n2664 GND.n2355 585
R3422 GND.n2666 GND.n2367 585
R3423 GND.n5369 GND.n2367 585
R3424 GND.n2668 GND.n2667 585
R3425 GND.n2667 GND.n2366 585
R3426 GND.n2669 GND.n2376 585
R3427 GND.n5361 GND.n2376 585
R3428 GND.n2671 GND.n2670 585
R3429 GND.n2670 GND.n2375 585
R3430 GND.n2672 GND.n2386 585
R3431 GND.n5349 GND.n2386 585
R3432 GND.n2674 GND.n2673 585
R3433 GND.n2673 GND.n2397 585
R3434 GND.n2675 GND.n2395 585
R3435 GND.n5341 GND.n2395 585
R3436 GND.n2677 GND.n2676 585
R3437 GND.n2676 GND.n2394 585
R3438 GND.n2678 GND.n2407 585
R3439 GND.n5329 GND.n2407 585
R3440 GND.n2680 GND.n2679 585
R3441 GND.n2679 GND.n2406 585
R3442 GND.n2681 GND.n2416 585
R3443 GND.n5321 GND.n2416 585
R3444 GND.n2683 GND.n2682 585
R3445 GND.n2682 GND.n2415 585
R3446 GND.n2684 GND.n2427 585
R3447 GND.n5309 GND.n2427 585
R3448 GND.n2686 GND.n2685 585
R3449 GND.n2685 GND.n2426 585
R3450 GND.n2687 GND.n2436 585
R3451 GND.n5301 GND.n2436 585
R3452 GND.n2689 GND.n2688 585
R3453 GND.n2688 GND.n2435 585
R3454 GND.n2690 GND.n2446 585
R3455 GND.n5289 GND.n2446 585
R3456 GND.n2692 GND.n2691 585
R3457 GND.n2691 GND.n2457 585
R3458 GND.n2693 GND.n2455 585
R3459 GND.n5281 GND.n2455 585
R3460 GND.n2695 GND.n2694 585
R3461 GND.n2694 GND.n2454 585
R3462 GND.n2696 GND.n2467 585
R3463 GND.n5269 GND.n2467 585
R3464 GND.n2698 GND.n2697 585
R3465 GND.n2697 GND.n2466 585
R3466 GND.n2699 GND.n2476 585
R3467 GND.n5261 GND.n2476 585
R3468 GND.n2701 GND.n2700 585
R3469 GND.n2700 GND.n2475 585
R3470 GND.n2702 GND.n2487 585
R3471 GND.n5249 GND.n2487 585
R3472 GND.n2704 GND.n2703 585
R3473 GND.n2703 GND.n2486 585
R3474 GND.n2705 GND.n2496 585
R3475 GND.n5241 GND.n2496 585
R3476 GND.n2707 GND.n2706 585
R3477 GND.n2706 GND.n2495 585
R3478 GND.n2708 GND.n2507 585
R3479 GND.n5229 GND.n2507 585
R3480 GND.n2710 GND.n2709 585
R3481 GND.n2710 GND.n2506 585
R3482 GND.n2716 GND.n2711 585
R3483 GND.n5182 GND.n2711 585
R3484 GND.n2718 GND.n2717 585
R3485 GND.n2718 GND.n2577 585
R3486 GND.n2728 GND.n2719 585
R3487 GND.n5175 GND.n2719 585
R3488 GND.n2730 GND.n2729 585
R3489 GND.n2730 GND.n2715 585
R3490 GND.n2739 GND.n2731 585
R3491 GND.n5082 GND.n2731 585
R3492 GND.n2741 GND.n2740 585
R3493 GND.n2741 GND.n2727 585
R3494 GND.n2744 GND.n2743 585
R3495 GND.n5075 GND.n2744 585
R3496 GND.n2742 GND.n2738 585
R3497 GND.n2738 GND.n2737 585
R3498 GND.n2528 GND.n2526 585
R3499 GND.n2530 GND.n2528 585
R3500 GND.n5222 GND.n5221 585
R3501 GND.n5221 GND.n5220 585
R3502 GND.n2527 GND.n2525 585
R3503 GND.n2757 GND.n2527 585
R3504 GND.n3507 GND.n3506 585
R3505 GND.n3506 GND.n2543 585
R3506 GND.n3508 GND.n2541 585
R3507 GND.n5210 GND.n2541 585
R3508 GND.n3510 GND.n3509 585
R3509 GND.n3509 GND.n2540 585
R3510 GND.n3511 GND.n2763 585
R3511 GND.n5058 GND.n2763 585
R3512 GND.n3513 GND.n3512 585
R3513 GND.n3512 GND.n2762 585
R3514 GND.n3514 GND.n2772 585
R3515 GND.n5050 GND.n2772 585
R3516 GND.n3516 GND.n3515 585
R3517 GND.n3515 GND.n2771 585
R3518 GND.n3517 GND.n2783 585
R3519 GND.n5034 GND.n2783 585
R3520 GND.n5612 GND.n1736 585
R3521 GND.n5613 GND.n5611 585
R3522 GND.n5609 GND.n5605 585
R3523 GND.n5617 GND.n5604 585
R3524 GND.n5618 GND.n5603 585
R3525 GND.n5619 GND.n5601 585
R3526 GND.n5600 GND.n5597 585
R3527 GND.n5623 GND.n5596 585
R3528 GND.n5624 GND.n5595 585
R3529 GND.n5625 GND.n5593 585
R3530 GND.n5592 GND.n5589 585
R3531 GND.n5629 GND.n5588 585
R3532 GND.n5587 GND.n1777 585
R3533 GND.n5584 GND.n2226 585
R3534 GND.n5583 GND.n5582 585
R3535 GND.n5575 GND.n2231 585
R3536 GND.n5577 GND.n5576 585
R3537 GND.n5573 GND.n2233 585
R3538 GND.n5572 GND.n5571 585
R3539 GND.n5565 GND.n2235 585
R3540 GND.n5567 GND.n5566 585
R3541 GND.n5566 GND.n1777 585
R3542 GND.n5693 GND.n5692 585
R3543 GND.n5692 GND.n5691 585
R3544 GND.n1735 GND.n1734 585
R3545 GND.n1737 GND.n1735 585
R3546 GND.n5544 GND.n2242 585
R3547 GND.n5559 GND.n2242 585
R3548 GND.n2255 GND.n2253 585
R3549 GND.n2253 GND.n2239 585
R3550 GND.n5549 GND.n5548 585
R3551 GND.n5550 GND.n5549 585
R3552 GND.n2254 GND.n2252 585
R3553 GND.n2252 GND.n2248 585
R3554 GND.n5520 GND.n2261 585
R3555 GND.n5534 GND.n2261 585
R3556 GND.n2275 GND.n2273 585
R3557 GND.n2273 GND.n2270 585
R3558 GND.n5525 GND.n5524 585
R3559 GND.n5526 GND.n5525 585
R3560 GND.n2274 GND.n2272 585
R3561 GND.n2272 GND.n2267 585
R3562 GND.n5500 GND.n2282 585
R3563 GND.n5514 GND.n2282 585
R3564 GND.n2295 GND.n2293 585
R3565 GND.n2293 GND.n2279 585
R3566 GND.n5505 GND.n5504 585
R3567 GND.n5506 GND.n5505 585
R3568 GND.n2294 GND.n2292 585
R3569 GND.n2292 GND.n2288 585
R3570 GND.n5480 GND.n2302 585
R3571 GND.n5494 GND.n2302 585
R3572 GND.n2315 GND.n2313 585
R3573 GND.n2313 GND.n2299 585
R3574 GND.n5485 GND.n5484 585
R3575 GND.n5486 GND.n5485 585
R3576 GND.n2314 GND.n2312 585
R3577 GND.n2312 GND.n2308 585
R3578 GND.n5460 GND.n2322 585
R3579 GND.n5474 GND.n2322 585
R3580 GND.n2334 GND.n2332 585
R3581 GND.n2332 GND.n2319 585
R3582 GND.n5465 GND.n5464 585
R3583 GND.n5466 GND.n5465 585
R3584 GND.n2333 GND.n2331 585
R3585 GND.n5455 GND.n2331 585
R3586 GND.n5379 GND.n5378 585
R3587 GND.n5378 GND.n2338 585
R3588 GND.n5380 GND.n2348 585
R3589 GND.n5396 GND.n2348 585
R3590 GND.n2362 GND.n2360 585
R3591 GND.n2360 GND.n2345 585
R3592 GND.n5385 GND.n5384 585
R3593 GND.n5386 GND.n5385 585
R3594 GND.n2361 GND.n2359 585
R3595 GND.n2359 GND.n2355 585
R3596 GND.n5355 GND.n2369 585
R3597 GND.n5369 GND.n2369 585
R3598 GND.n2382 GND.n2380 585
R3599 GND.n2380 GND.n2366 585
R3600 GND.n5360 GND.n5359 585
R3601 GND.n5361 GND.n5360 585
R3602 GND.n2381 GND.n2379 585
R3603 GND.n2379 GND.n2375 585
R3604 GND.n5335 GND.n2388 585
R3605 GND.n5349 GND.n2388 585
R3606 GND.n2402 GND.n2400 585
R3607 GND.n2400 GND.n2397 585
R3608 GND.n5340 GND.n5339 585
R3609 GND.n5341 GND.n5340 585
R3610 GND.n2401 GND.n2399 585
R3611 GND.n2399 GND.n2394 585
R3612 GND.n5315 GND.n2409 585
R3613 GND.n5329 GND.n2409 585
R3614 GND.n2422 GND.n2420 585
R3615 GND.n2420 GND.n2406 585
R3616 GND.n5320 GND.n5319 585
R3617 GND.n5321 GND.n5320 585
R3618 GND.n2421 GND.n2419 585
R3619 GND.n2419 GND.n2415 585
R3620 GND.n5295 GND.n2429 585
R3621 GND.n5309 GND.n2429 585
R3622 GND.n2442 GND.n2440 585
R3623 GND.n2440 GND.n2426 585
R3624 GND.n5300 GND.n5299 585
R3625 GND.n5301 GND.n5300 585
R3626 GND.n2441 GND.n2439 585
R3627 GND.n2439 GND.n2435 585
R3628 GND.n5275 GND.n2448 585
R3629 GND.n5289 GND.n2448 585
R3630 GND.n2462 GND.n2460 585
R3631 GND.n2460 GND.n2457 585
R3632 GND.n5280 GND.n5279 585
R3633 GND.n5281 GND.n5280 585
R3634 GND.n2461 GND.n2459 585
R3635 GND.n2459 GND.n2454 585
R3636 GND.n5255 GND.n2469 585
R3637 GND.n5269 GND.n2469 585
R3638 GND.n2482 GND.n2480 585
R3639 GND.n2480 GND.n2466 585
R3640 GND.n5260 GND.n5259 585
R3641 GND.n5261 GND.n5260 585
R3642 GND.n2481 GND.n2479 585
R3643 GND.n2479 GND.n2475 585
R3644 GND.n5235 GND.n2489 585
R3645 GND.n5249 GND.n2489 585
R3646 GND.n2502 GND.n2500 585
R3647 GND.n2500 GND.n2486 585
R3648 GND.n5240 GND.n5239 585
R3649 GND.n5241 GND.n5240 585
R3650 GND.n2501 GND.n2499 585
R3651 GND.n2499 GND.n2495 585
R3652 GND.n5186 GND.n2509 585
R3653 GND.n5229 GND.n2509 585
R3654 GND.n2574 GND.n2573 585
R3655 GND.n2573 GND.n2506 585
R3656 GND.n5190 GND.n2572 585
R3657 GND.n5182 GND.n2572 585
R3658 GND.n5191 GND.n2571 585
R3659 GND.n2577 GND.n2571 585
R3660 GND.n5192 GND.n2570 585
R3661 GND.n5175 GND.n2570 585
R3662 GND.n2714 GND.n2565 585
R3663 GND.n2715 GND.n2714 585
R3664 GND.n5196 GND.n2564 585
R3665 GND.n5082 GND.n2564 585
R3666 GND.n5197 GND.n2563 585
R3667 GND.n2727 GND.n2563 585
R3668 GND.n5198 GND.n2562 585
R3669 GND.n5075 GND.n2562 585
R3670 GND.n2736 GND.n2556 585
R3671 GND.n2737 GND.n2736 585
R3672 GND.n5202 GND.n2555 585
R3673 GND.n2555 GND.n2530 585
R3674 GND.n5203 GND.n2532 585
R3675 GND.n5220 GND.n2532 585
R3676 GND.n5204 GND.n2554 585
R3677 GND.n2757 GND.n2554 585
R3678 GND.n2548 GND.n2546 585
R3679 GND.n2546 GND.n2543 585
R3680 GND.n5209 GND.n5208 585
R3681 GND.n5210 GND.n5209 585
R3682 GND.n2547 GND.n2545 585
R3683 GND.n2545 GND.n2540 585
R3684 GND.n5044 GND.n2765 585
R3685 GND.n5058 GND.n2765 585
R3686 GND.n2778 GND.n2776 585
R3687 GND.n2776 GND.n2762 585
R3688 GND.n5049 GND.n5048 585
R3689 GND.n5050 GND.n5049 585
R3690 GND.n2777 GND.n2775 585
R3691 GND.n2775 GND.n2771 585
R3692 GND.n3485 GND.n2785 585
R3693 GND.n5034 GND.n2785 585
R3694 GND.n7467 GND.n523 585
R3695 GND.n523 GND.n522 585
R3696 GND.n7469 GND.n7468 585
R3697 GND.n7470 GND.n7469 585
R3698 GND.n510 GND.n509 585
R3699 GND.n513 GND.n510 585
R3700 GND.n7478 GND.n7477 585
R3701 GND.n7477 GND.n7476 585
R3702 GND.n7479 GND.n504 585
R3703 GND.n504 GND.n503 585
R3704 GND.n7481 GND.n7480 585
R3705 GND.n7482 GND.n7481 585
R3706 GND.n491 GND.n490 585
R3707 GND.n500 GND.n491 585
R3708 GND.n7490 GND.n7489 585
R3709 GND.n7489 GND.n7488 585
R3710 GND.n7491 GND.n485 585
R3711 GND.n485 GND.n484 585
R3712 GND.n7493 GND.n7492 585
R3713 GND.n7494 GND.n7493 585
R3714 GND.n472 GND.n471 585
R3715 GND.n475 GND.n472 585
R3716 GND.n7502 GND.n7501 585
R3717 GND.n7501 GND.n7500 585
R3718 GND.n7503 GND.n466 585
R3719 GND.n466 GND.n465 585
R3720 GND.n7505 GND.n7504 585
R3721 GND.n7506 GND.n7505 585
R3722 GND.n452 GND.n451 585
R3723 GND.n456 GND.n452 585
R3724 GND.n7514 GND.n7513 585
R3725 GND.n7513 GND.n7512 585
R3726 GND.n7515 GND.n446 585
R3727 GND.n446 GND.n445 585
R3728 GND.n7517 GND.n7516 585
R3729 GND.n7518 GND.n7517 585
R3730 GND.n432 GND.n431 585
R3731 GND.n436 GND.n432 585
R3732 GND.n7526 GND.n7525 585
R3733 GND.n7525 GND.n7524 585
R3734 GND.n7527 GND.n426 585
R3735 GND.n433 GND.n426 585
R3736 GND.n7529 GND.n7528 585
R3737 GND.n7530 GND.n7529 585
R3738 GND.n414 GND.n413 585
R3739 GND.n417 GND.n414 585
R3740 GND.n7538 GND.n7537 585
R3741 GND.n7537 GND.n7536 585
R3742 GND.n7539 GND.n408 585
R3743 GND.n408 GND.n407 585
R3744 GND.n7541 GND.n7540 585
R3745 GND.n7542 GND.n7541 585
R3746 GND.n395 GND.n394 585
R3747 GND.n398 GND.n395 585
R3748 GND.n7550 GND.n7549 585
R3749 GND.n7549 GND.n7548 585
R3750 GND.n7551 GND.n389 585
R3751 GND.n389 GND.n388 585
R3752 GND.n7553 GND.n7552 585
R3753 GND.n7554 GND.n7553 585
R3754 GND.n376 GND.n375 585
R3755 GND.n379 GND.n376 585
R3756 GND.n7562 GND.n7561 585
R3757 GND.n7561 GND.n7560 585
R3758 GND.n7563 GND.n370 585
R3759 GND.n370 GND.n369 585
R3760 GND.n7565 GND.n7564 585
R3761 GND.n7566 GND.n7565 585
R3762 GND.n357 GND.n356 585
R3763 GND.n360 GND.n357 585
R3764 GND.n7574 GND.n7573 585
R3765 GND.n7573 GND.n7572 585
R3766 GND.n7575 GND.n351 585
R3767 GND.n351 GND.n350 585
R3768 GND.n7577 GND.n7576 585
R3769 GND.n7578 GND.n7577 585
R3770 GND.n338 GND.n337 585
R3771 GND.n341 GND.n338 585
R3772 GND.n7586 GND.n7585 585
R3773 GND.n7585 GND.n7584 585
R3774 GND.n7587 GND.n332 585
R3775 GND.n332 GND.n331 585
R3776 GND.n7589 GND.n7588 585
R3777 GND.n7590 GND.n7589 585
R3778 GND.n316 GND.n315 585
R3779 GND.n319 GND.n316 585
R3780 GND.n7598 GND.n7597 585
R3781 GND.n7597 GND.n7596 585
R3782 GND.n7599 GND.n310 585
R3783 GND.n7234 GND.n310 585
R3784 GND.n7601 GND.n7600 585
R3785 GND.n7602 GND.n7601 585
R3786 GND.n311 GND.n309 585
R3787 GND.n309 GND.n298 585
R3788 GND.n1024 GND.n296 585
R3789 GND.n7608 GND.n296 585
R3790 GND.n1026 GND.n1025 585
R3791 GND.n1025 GND.n287 585
R3792 GND.n1027 GND.n285 585
R3793 GND.n7614 GND.n285 585
R3794 GND.n1029 GND.n1028 585
R3795 GND.n1028 GND.n277 585
R3796 GND.n1030 GND.n275 585
R3797 GND.n7620 GND.n275 585
R3798 GND.n1032 GND.n1031 585
R3799 GND.n1031 GND.n267 585
R3800 GND.n1033 GND.n265 585
R3801 GND.n7626 GND.n265 585
R3802 GND.n1035 GND.n1034 585
R3803 GND.n1034 GND.n264 585
R3804 GND.n1036 GND.n253 585
R3805 GND.n7632 GND.n253 585
R3806 GND.n1038 GND.n1037 585
R3807 GND.n1037 GND.n252 585
R3808 GND.n1039 GND.n620 585
R3809 GND.n7208 GND.n620 585
R3810 GND.n1042 GND.n1041 585
R3811 GND.n1042 GND.n619 585
R3812 GND.n1044 GND.n1043 585
R3813 GND.n1043 GND.n236 585
R3814 GND.n1046 GND.n234 585
R3815 GND.n7641 GND.n234 585
R3816 GND.n1048 GND.n1047 585
R3817 GND.n1047 GND.n233 585
R3818 GND.n1050 GND.n631 585
R3819 GND.n7168 GND.n631 585
R3820 GND.n1052 GND.n1051 585
R3821 GND.n1051 GND.n630 585
R3822 GND.n1053 GND.n636 585
R3823 GND.n7160 GND.n636 585
R3824 GND.n1055 GND.n1013 585
R3825 GND.n1013 GND.n635 585
R3826 GND.n1056 GND.n645 585
R3827 GND.n7145 GND.n645 585
R3828 GND.n1057 GND.n667 585
R3829 GND.n7129 GND.n667 585
R3830 GND.n1059 GND.n1058 585
R3831 GND.n1058 GND.n657 585
R3832 GND.n1060 GND.n655 585
R3833 GND.n7135 GND.n655 585
R3834 GND.n1062 GND.n1061 585
R3835 GND.n1061 GND.n654 585
R3836 GND.n1063 GND.n674 585
R3837 GND.n7107 GND.n674 585
R3838 GND.n1065 GND.n1064 585
R3839 GND.n1064 GND.n673 585
R3840 GND.n1066 GND.n683 585
R3841 GND.n7099 GND.n683 585
R3842 GND.n1068 GND.n1067 585
R3843 GND.n1067 GND.n682 585
R3844 GND.n1069 GND.n695 585
R3845 GND.n7079 GND.n695 585
R3846 GND.n1071 GND.n1070 585
R3847 GND.n1070 GND.n694 585
R3848 GND.n1072 GND.n703 585
R3849 GND.n7071 GND.n703 585
R3850 GND.n1073 GND.n714 585
R3851 GND.n7060 GND.n714 585
R3852 GND.n1075 GND.n1074 585
R3853 GND.n1074 GND.n713 585
R3854 GND.n1076 GND.n721 585
R3855 GND.n7037 GND.n721 585
R3856 GND.n1078 GND.n1077 585
R3857 GND.n1077 GND.n720 585
R3858 GND.n1079 GND.n731 585
R3859 GND.n7027 GND.n731 585
R3860 GND.n1081 GND.n1080 585
R3861 GND.n1080 GND.n730 585
R3862 GND.n1082 GND.n743 585
R3863 GND.n7011 GND.n743 585
R3864 GND.n1084 GND.n1083 585
R3865 GND.n1083 GND.n742 585
R3866 GND.n1085 GND.n752 585
R3867 GND.n7003 GND.n752 585
R3868 GND.n1087 GND.n1086 585
R3869 GND.n1086 GND.n751 585
R3870 GND.n1088 GND.n763 585
R3871 GND.n6991 GND.n763 585
R3872 GND.n1090 GND.n1089 585
R3873 GND.n1089 GND.n762 585
R3874 GND.n1091 GND.n772 585
R3875 GND.n6983 GND.n772 585
R3876 GND.n1093 GND.n1092 585
R3877 GND.n1092 GND.n771 585
R3878 GND.n1094 GND.n783 585
R3879 GND.n6971 GND.n783 585
R3880 GND.n1096 GND.n1095 585
R3881 GND.n1095 GND.n782 585
R3882 GND.n1097 GND.n792 585
R3883 GND.n6963 GND.n792 585
R3884 GND.n1099 GND.n1098 585
R3885 GND.n1098 GND.n791 585
R3886 GND.n1100 GND.n803 585
R3887 GND.n6951 GND.n803 585
R3888 GND.n1102 GND.n1101 585
R3889 GND.n1101 GND.n802 585
R3890 GND.n1103 GND.n812 585
R3891 GND.n6943 GND.n812 585
R3892 GND.n1105 GND.n1104 585
R3893 GND.n1104 GND.n811 585
R3894 GND.n1106 GND.n822 585
R3895 GND.n6931 GND.n822 585
R3896 GND.n1108 GND.n1107 585
R3897 GND.n1107 GND.n833 585
R3898 GND.n1109 GND.n831 585
R3899 GND.n6923 GND.n831 585
R3900 GND.n1111 GND.n1110 585
R3901 GND.n1110 GND.n830 585
R3902 GND.n1112 GND.n843 585
R3903 GND.n6911 GND.n843 585
R3904 GND.n1114 GND.n1113 585
R3905 GND.n1113 GND.n842 585
R3906 GND.n1115 GND.n852 585
R3907 GND.n6903 GND.n852 585
R3908 GND.n1117 GND.n1116 585
R3909 GND.n1116 GND.n851 585
R3910 GND.n1118 GND.n863 585
R3911 GND.n6891 GND.n863 585
R3912 GND.n1120 GND.n1119 585
R3913 GND.n1119 GND.n862 585
R3914 GND.n1121 GND.n872 585
R3915 GND.n6883 GND.n872 585
R3916 GND.n1123 GND.n1122 585
R3917 GND.n1122 GND.n871 585
R3918 GND.n1124 GND.n883 585
R3919 GND.n6871 GND.n883 585
R3920 GND.n1126 GND.n1125 585
R3921 GND.n1125 GND.n882 585
R3922 GND.n1127 GND.n891 585
R3923 GND.n6863 GND.n891 585
R3924 GND.n1128 GND.n902 585
R3925 GND.n6852 GND.n902 585
R3926 GND.n1130 GND.n1129 585
R3927 GND.n1129 GND.n901 585
R3928 GND.n1131 GND.n909 585
R3929 GND.n6762 GND.n909 585
R3930 GND.n1133 GND.n1132 585
R3931 GND.n1132 GND.n908 585
R3932 GND.n1134 GND.n919 585
R3933 GND.n6752 GND.n919 585
R3934 GND.n1136 GND.n1135 585
R3935 GND.n1135 GND.n918 585
R3936 GND.n1137 GND.n932 585
R3937 GND.n6734 GND.n932 585
R3938 GND.n6723 GND.n6722 585
R3939 GND.n6721 GND.n957 585
R3940 GND.n6720 GND.n956 585
R3941 GND.n6725 GND.n956 585
R3942 GND.n6719 GND.n6718 585
R3943 GND.n6717 GND.n6716 585
R3944 GND.n6715 GND.n6714 585
R3945 GND.n6713 GND.n6712 585
R3946 GND.n6711 GND.n6710 585
R3947 GND.n6708 GND.n6707 585
R3948 GND.n6706 GND.n6705 585
R3949 GND.n6704 GND.n6703 585
R3950 GND.n6702 GND.n6701 585
R3951 GND.n6700 GND.n6699 585
R3952 GND.n6698 GND.n6697 585
R3953 GND.n6696 GND.n6695 585
R3954 GND.n6694 GND.n6693 585
R3955 GND.n6692 GND.n6691 585
R3956 GND.n6690 GND.n6689 585
R3957 GND.n6684 GND.n6681 585
R3958 GND.n6685 GND.n930 585
R3959 GND.n6725 GND.n930 585
R3960 GND.n7426 GND.n7425 585
R3961 GND.n7428 GND.n563 585
R3962 GND.n7430 GND.n7429 585
R3963 GND.n7431 GND.n556 585
R3964 GND.n7433 GND.n7432 585
R3965 GND.n7435 GND.n554 585
R3966 GND.n7437 GND.n7436 585
R3967 GND.n7438 GND.n550 585
R3968 GND.n7440 GND.n7439 585
R3969 GND.n7442 GND.n547 585
R3970 GND.n7444 GND.n7443 585
R3971 GND.n548 GND.n541 585
R3972 GND.n7448 GND.n545 585
R3973 GND.n7449 GND.n537 585
R3974 GND.n7451 GND.n7450 585
R3975 GND.n7453 GND.n535 585
R3976 GND.n7455 GND.n7454 585
R3977 GND.n7456 GND.n530 585
R3978 GND.n7458 GND.n7457 585
R3979 GND.n7460 GND.n529 585
R3980 GND.n7461 GND.n527 585
R3981 GND.n7464 GND.n7463 585
R3982 GND.n7421 GND.n565 585
R3983 GND.n565 GND.n522 585
R3984 GND.n7420 GND.n520 585
R3985 GND.n7470 GND.n520 585
R3986 GND.n7419 GND.n7418 585
R3987 GND.n7418 GND.n513 585
R3988 GND.n7417 GND.n511 585
R3989 GND.n7476 GND.n511 585
R3990 GND.n7416 GND.n7415 585
R3991 GND.n7415 GND.n503 585
R3992 GND.n7413 GND.n501 585
R3993 GND.n7482 GND.n501 585
R3994 GND.n7412 GND.n7411 585
R3995 GND.n7411 GND.n500 585
R3996 GND.n7410 GND.n492 585
R3997 GND.n7488 GND.n492 585
R3998 GND.n7409 GND.n7408 585
R3999 GND.n7408 GND.n484 585
R4000 GND.n7406 GND.n482 585
R4001 GND.n7494 GND.n482 585
R4002 GND.n7405 GND.n7404 585
R4003 GND.n7404 GND.n475 585
R4004 GND.n7403 GND.n473 585
R4005 GND.n7500 GND.n473 585
R4006 GND.n7402 GND.n7401 585
R4007 GND.n7401 GND.n465 585
R4008 GND.n7399 GND.n463 585
R4009 GND.n7506 GND.n463 585
R4010 GND.n7398 GND.n7397 585
R4011 GND.n7397 GND.n456 585
R4012 GND.n7396 GND.n454 585
R4013 GND.n7512 GND.n454 585
R4014 GND.n7395 GND.n7394 585
R4015 GND.n7394 GND.n445 585
R4016 GND.n7392 GND.n443 585
R4017 GND.n7518 GND.n443 585
R4018 GND.n7391 GND.n7390 585
R4019 GND.n7390 GND.n436 585
R4020 GND.n7389 GND.n434 585
R4021 GND.n7524 GND.n434 585
R4022 GND.n7388 GND.n7387 585
R4023 GND.n7387 GND.n433 585
R4024 GND.n7385 GND.n424 585
R4025 GND.n7530 GND.n424 585
R4026 GND.n7384 GND.n7383 585
R4027 GND.n7383 GND.n417 585
R4028 GND.n7382 GND.n415 585
R4029 GND.n7536 GND.n415 585
R4030 GND.n7381 GND.n7380 585
R4031 GND.n7380 GND.n407 585
R4032 GND.n7378 GND.n405 585
R4033 GND.n7542 GND.n405 585
R4034 GND.n7377 GND.n7376 585
R4035 GND.n7376 GND.n398 585
R4036 GND.n7375 GND.n396 585
R4037 GND.n7548 GND.n396 585
R4038 GND.n7374 GND.n7373 585
R4039 GND.n7373 GND.n388 585
R4040 GND.n7371 GND.n386 585
R4041 GND.n7554 GND.n386 585
R4042 GND.n7370 GND.n7369 585
R4043 GND.n7369 GND.n379 585
R4044 GND.n7368 GND.n377 585
R4045 GND.n7560 GND.n377 585
R4046 GND.n7367 GND.n7366 585
R4047 GND.n7366 GND.n369 585
R4048 GND.n7364 GND.n367 585
R4049 GND.n7566 GND.n367 585
R4050 GND.n7363 GND.n7362 585
R4051 GND.n7362 GND.n360 585
R4052 GND.n7361 GND.n358 585
R4053 GND.n7572 GND.n358 585
R4054 GND.n7360 GND.n7359 585
R4055 GND.n7359 GND.n350 585
R4056 GND.n7357 GND.n348 585
R4057 GND.n7578 GND.n348 585
R4058 GND.n7356 GND.n7355 585
R4059 GND.n7355 GND.n341 585
R4060 GND.n7354 GND.n339 585
R4061 GND.n7584 GND.n339 585
R4062 GND.n7353 GND.n7352 585
R4063 GND.n7352 GND.n331 585
R4064 GND.n7350 GND.n329 585
R4065 GND.n7590 GND.n329 585
R4066 GND.n7349 GND.n7348 585
R4067 GND.n7348 GND.n319 585
R4068 GND.n7347 GND.n317 585
R4069 GND.n7596 GND.n317 585
R4070 GND.n305 GND.n304 585
R4071 GND.n7234 GND.n305 585
R4072 GND.n7604 GND.n7603 585
R4073 GND.n7603 GND.n7602 585
R4074 GND.n7605 GND.n300 585
R4075 GND.n300 GND.n298 585
R4076 GND.n7607 GND.n7606 585
R4077 GND.n7608 GND.n7607 585
R4078 GND.n284 GND.n283 585
R4079 GND.n287 GND.n284 585
R4080 GND.n7616 GND.n7615 585
R4081 GND.n7615 GND.n7614 585
R4082 GND.n7617 GND.n279 585
R4083 GND.n279 GND.n277 585
R4084 GND.n7619 GND.n7618 585
R4085 GND.n7620 GND.n7619 585
R4086 GND.n263 GND.n262 585
R4087 GND.n267 GND.n263 585
R4088 GND.n7628 GND.n7627 585
R4089 GND.n7627 GND.n7626 585
R4090 GND.n7629 GND.n257 585
R4091 GND.n264 GND.n257 585
R4092 GND.n7631 GND.n7630 585
R4093 GND.n7632 GND.n7631 585
R4094 GND.n258 GND.n256 585
R4095 GND.n256 GND.n252 585
R4096 GND.n7204 GND.n7203 585
R4097 GND.n7208 GND.n7204 585
R4098 GND.n623 GND.n622 585
R4099 GND.n622 GND.n619 585
R4100 GND.n7174 GND.n7173 585
R4101 GND.n7173 GND.n236 585
R4102 GND.n7172 GND.n237 585
R4103 GND.n7641 GND.n237 585
R4104 GND.n7171 GND.n7170 585
R4105 GND.n7170 GND.n233 585
R4106 GND.n7169 GND.n627 585
R4107 GND.n7169 GND.n7168 585
R4108 GND.n7157 GND.n629 585
R4109 GND.n630 GND.n629 585
R4110 GND.n7159 GND.n7158 585
R4111 GND.n7160 GND.n7159 585
R4112 GND.n640 GND.n639 585
R4113 GND.n639 GND.n635 585
R4114 GND.n666 GND.n647 585
R4115 GND.n7145 GND.n647 585
R4116 GND.n7131 GND.n7130 585
R4117 GND.n7130 GND.n7129 585
R4118 GND.n7132 GND.n660 585
R4119 GND.n660 GND.n657 585
R4120 GND.n7134 GND.n7133 585
R4121 GND.n7135 GND.n7134 585
R4122 GND.n661 GND.n659 585
R4123 GND.n659 GND.n654 585
R4124 GND.n7095 GND.n676 585
R4125 GND.n7107 GND.n676 585
R4126 GND.n7096 GND.n687 585
R4127 GND.n687 GND.n673 585
R4128 GND.n7098 GND.n7097 585
R4129 GND.n7099 GND.n7098 585
R4130 GND.n688 GND.n686 585
R4131 GND.n686 GND.n682 585
R4132 GND.n7067 GND.n697 585
R4133 GND.n7079 GND.n697 585
R4134 GND.n7068 GND.n707 585
R4135 GND.n707 GND.n694 585
R4136 GND.n7070 GND.n7069 585
R4137 GND.n7071 GND.n7070 585
R4138 GND.n708 GND.n706 585
R4139 GND.n7060 GND.n706 585
R4140 GND.n7022 GND.n7021 585
R4141 GND.n7021 GND.n713 585
R4142 GND.n7023 GND.n723 585
R4143 GND.n7037 GND.n723 585
R4144 GND.n7024 GND.n735 585
R4145 GND.n735 GND.n720 585
R4146 GND.n7026 GND.n7025 585
R4147 GND.n7027 GND.n7026 585
R4148 GND.n736 GND.n734 585
R4149 GND.n734 GND.n730 585
R4150 GND.n6999 GND.n745 585
R4151 GND.n7011 GND.n745 585
R4152 GND.n7000 GND.n756 585
R4153 GND.n756 GND.n742 585
R4154 GND.n7002 GND.n7001 585
R4155 GND.n7003 GND.n7002 585
R4156 GND.n757 GND.n755 585
R4157 GND.n755 GND.n751 585
R4158 GND.n6979 GND.n765 585
R4159 GND.n6991 GND.n765 585
R4160 GND.n6980 GND.n776 585
R4161 GND.n776 GND.n762 585
R4162 GND.n6982 GND.n6981 585
R4163 GND.n6983 GND.n6982 585
R4164 GND.n777 GND.n775 585
R4165 GND.n775 GND.n771 585
R4166 GND.n6959 GND.n785 585
R4167 GND.n6971 GND.n785 585
R4168 GND.n6960 GND.n796 585
R4169 GND.n796 GND.n782 585
R4170 GND.n6962 GND.n6961 585
R4171 GND.n6963 GND.n6962 585
R4172 GND.n797 GND.n795 585
R4173 GND.n795 GND.n791 585
R4174 GND.n6939 GND.n805 585
R4175 GND.n6951 GND.n805 585
R4176 GND.n6940 GND.n816 585
R4177 GND.n816 GND.n802 585
R4178 GND.n6942 GND.n6941 585
R4179 GND.n6943 GND.n6942 585
R4180 GND.n817 GND.n815 585
R4181 GND.n815 GND.n811 585
R4182 GND.n6919 GND.n824 585
R4183 GND.n6931 GND.n824 585
R4184 GND.n6920 GND.n836 585
R4185 GND.n836 GND.n833 585
R4186 GND.n6922 GND.n6921 585
R4187 GND.n6923 GND.n6922 585
R4188 GND.n837 GND.n835 585
R4189 GND.n835 GND.n830 585
R4190 GND.n6899 GND.n845 585
R4191 GND.n6911 GND.n845 585
R4192 GND.n6900 GND.n856 585
R4193 GND.n856 GND.n842 585
R4194 GND.n6902 GND.n6901 585
R4195 GND.n6903 GND.n6902 585
R4196 GND.n857 GND.n855 585
R4197 GND.n855 GND.n851 585
R4198 GND.n6879 GND.n865 585
R4199 GND.n6891 GND.n865 585
R4200 GND.n6880 GND.n876 585
R4201 GND.n876 GND.n862 585
R4202 GND.n6882 GND.n6881 585
R4203 GND.n6883 GND.n6882 585
R4204 GND.n877 GND.n875 585
R4205 GND.n875 GND.n871 585
R4206 GND.n6859 GND.n885 585
R4207 GND.n6871 GND.n885 585
R4208 GND.n6860 GND.n895 585
R4209 GND.n895 GND.n882 585
R4210 GND.n6862 GND.n6861 585
R4211 GND.n6863 GND.n6862 585
R4212 GND.n896 GND.n894 585
R4213 GND.n6852 GND.n894 585
R4214 GND.n6747 GND.n6746 585
R4215 GND.n6746 GND.n901 585
R4216 GND.n6748 GND.n911 585
R4217 GND.n6762 GND.n911 585
R4218 GND.n6749 GND.n923 585
R4219 GND.n923 GND.n908 585
R4220 GND.n6751 GND.n6750 585
R4221 GND.n6752 GND.n6751 585
R4222 GND.n924 GND.n922 585
R4223 GND.n922 GND.n918 585
R4224 GND.n6736 GND.n6735 585
R4225 GND.n6735 GND.n6734 585
R4226 GND.n6620 GND.n1173 585
R4227 GND.n6576 GND.n1173 585
R4228 GND.n6619 GND.n6618 585
R4229 GND.n6618 GND.n6617 585
R4230 GND.n1181 GND.n1180 585
R4231 GND.n1192 GND.n1181 585
R4232 GND.n6592 GND.n6591 585
R4233 GND.n6593 GND.n6592 585
R4234 GND.n6590 GND.n1193 585
R4235 GND.n1193 GND.n1190 585
R4236 GND.n6589 GND.n6588 585
R4237 GND.n6588 GND.n6587 585
R4238 GND.n1195 GND.n1194 585
R4239 GND.n1196 GND.n1195 585
R4240 GND.n6527 GND.n6526 585
R4241 GND.n6528 GND.n6527 585
R4242 GND.n6525 GND.n1203 585
R4243 GND.n6521 GND.n1203 585
R4244 GND.n6524 GND.n6523 585
R4245 GND.n6523 GND.n6522 585
R4246 GND.n1205 GND.n1204 585
R4247 GND.n1211 GND.n1205 585
R4248 GND.n6514 GND.n6513 585
R4249 GND.n6515 GND.n6514 585
R4250 GND.n6512 GND.n1213 585
R4251 GND.n1213 GND.n1210 585
R4252 GND.n6511 GND.n6510 585
R4253 GND.n6510 GND.n6509 585
R4254 GND.n1215 GND.n1214 585
R4255 GND.n1226 GND.n1215 585
R4256 GND.n6487 GND.n6486 585
R4257 GND.n6488 GND.n6487 585
R4258 GND.n6485 GND.n1227 585
R4259 GND.n1227 GND.n1224 585
R4260 GND.n6484 GND.n6483 585
R4261 GND.n6483 GND.n6482 585
R4262 GND.n1229 GND.n1228 585
R4263 GND.n1230 GND.n1229 585
R4264 GND.n6469 GND.n6468 585
R4265 GND.n6470 GND.n6469 585
R4266 GND.n6467 GND.n1237 585
R4267 GND.n1242 GND.n1237 585
R4268 GND.n6466 GND.n6465 585
R4269 GND.n6465 GND.n6464 585
R4270 GND.n1239 GND.n1238 585
R4271 GND.n1240 GND.n1239 585
R4272 GND.n6448 GND.n6447 585
R4273 GND.n6449 GND.n6448 585
R4274 GND.n6446 GND.n1252 585
R4275 GND.n1252 GND.n1249 585
R4276 GND.n6445 GND.n6444 585
R4277 GND.n6444 GND.n6443 585
R4278 GND.n1254 GND.n1253 585
R4279 GND.n1261 GND.n1254 585
R4280 GND.n6431 GND.n6430 585
R4281 GND.n6432 GND.n6431 585
R4282 GND.n6429 GND.n1263 585
R4283 GND.n1263 GND.n1260 585
R4284 GND.n6428 GND.n6427 585
R4285 GND.n6427 GND.n6426 585
R4286 GND.n1265 GND.n1264 585
R4287 GND.n1276 GND.n1265 585
R4288 GND.n6413 GND.n6412 585
R4289 GND.n6414 GND.n6413 585
R4290 GND.n6411 GND.n1277 585
R4291 GND.n1277 GND.n1274 585
R4292 GND.n6410 GND.n6409 585
R4293 GND.n6409 GND.n6408 585
R4294 GND.n1279 GND.n1278 585
R4295 GND.n1280 GND.n1279 585
R4296 GND.n6395 GND.n6394 585
R4297 GND.n6396 GND.n6395 585
R4298 GND.n6393 GND.n1287 585
R4299 GND.n6389 GND.n1287 585
R4300 GND.n6392 GND.n6391 585
R4301 GND.n6391 GND.n6390 585
R4302 GND.n1289 GND.n1288 585
R4303 GND.n1295 GND.n1289 585
R4304 GND.n6382 GND.n6381 585
R4305 GND.n6383 GND.n6382 585
R4306 GND.n6380 GND.n1297 585
R4307 GND.n1297 GND.n1294 585
R4308 GND.n6379 GND.n6378 585
R4309 GND.n6378 GND.n6377 585
R4310 GND.n1299 GND.n1298 585
R4311 GND.n1309 GND.n1299 585
R4312 GND.n6355 GND.n6354 585
R4313 GND.n6356 GND.n6355 585
R4314 GND.n6353 GND.n1310 585
R4315 GND.n6348 GND.n1310 585
R4316 GND.n6352 GND.n6351 585
R4317 GND.n6351 GND.n6350 585
R4318 GND.n1312 GND.n1311 585
R4319 GND.n6338 GND.n1312 585
R4320 GND.n6336 GND.n6335 585
R4321 GND.n6337 GND.n6336 585
R4322 GND.n6334 GND.n1318 585
R4323 GND.n1323 GND.n1318 585
R4324 GND.n6333 GND.n6332 585
R4325 GND.n6332 GND.n6331 585
R4326 GND.n1320 GND.n1319 585
R4327 GND.n6206 GND.n1320 585
R4328 GND.n6216 GND.n6215 585
R4329 GND.n6215 GND.n1333 585
R4330 GND.n6217 GND.n6214 585
R4331 GND.n6214 GND.n1331 585
R4332 GND.n6219 GND.n6218 585
R4333 GND.n6220 GND.n6219 585
R4334 GND.n1435 GND.n1434 585
R4335 GND.n1435 GND.n1421 585
R4336 GND.n6256 GND.n6255 585
R4337 GND.n6255 GND.n6254 585
R4338 GND.n6257 GND.n1432 585
R4339 GND.n6225 GND.n1432 585
R4340 GND.n6259 GND.n6258 585
R4341 GND.n6260 GND.n6259 585
R4342 GND.n1433 GND.n1431 585
R4343 GND.n6229 GND.n1431 585
R4344 GND.n6242 GND.n6241 585
R4345 GND.n6243 GND.n6242 585
R4346 GND.n6240 GND.n1446 585
R4347 GND.n6235 GND.n1446 585
R4348 GND.n6239 GND.n6238 585
R4349 GND.n6238 GND.n6237 585
R4350 GND.n1448 GND.n1447 585
R4351 GND.n6196 GND.n1448 585
R4352 GND.n6180 GND.n6179 585
R4353 GND.n6179 GND.n6178 585
R4354 GND.n6181 GND.n1462 585
R4355 GND.n6176 GND.n1462 585
R4356 GND.n6183 GND.n6182 585
R4357 GND.n6184 GND.n6183 585
R4358 GND.n1463 GND.n1461 585
R4359 GND.n6170 GND.n1461 585
R4360 GND.n6134 GND.n1490 585
R4361 GND.n6134 GND.n6133 585
R4362 GND.n6136 GND.n6135 585
R4363 GND.n6135 GND.n1477 585
R4364 GND.n6137 GND.n1488 585
R4365 GND.n1488 GND.n1475 585
R4366 GND.n6139 GND.n6138 585
R4367 GND.n6140 GND.n6139 585
R4368 GND.n1489 GND.n1487 585
R4369 GND.n1487 GND.n1483 585
R4370 GND.n6092 GND.n6091 585
R4371 GND.n6091 GND.n1496 585
R4372 GND.n6093 GND.n1507 585
R4373 GND.t1 GND.n1507 585
R4374 GND.n6095 GND.n6094 585
R4375 GND.n6096 GND.n6095 585
R4376 GND.n6090 GND.n1506 585
R4377 GND.n1506 GND.n1502 585
R4378 GND.n6089 GND.n6088 585
R4379 GND.n6088 GND.n6087 585
R4380 GND.n1509 GND.n1508 585
R4381 GND.n6037 GND.n1509 585
R4382 GND.n6074 GND.n6073 585
R4383 GND.n6075 GND.n6074 585
R4384 GND.n6072 GND.n1521 585
R4385 GND.n1521 GND.n1518 585
R4386 GND.n6071 GND.n6070 585
R4387 GND.n6070 GND.n6069 585
R4388 GND.n1523 GND.n1522 585
R4389 GND.n6044 GND.n1523 585
R4390 GND.n6057 GND.n6056 585
R4391 GND.n6058 GND.n6057 585
R4392 GND.n6055 GND.n1538 585
R4393 GND.n6050 GND.n1538 585
R4394 GND.n6054 GND.n6053 585
R4395 GND.n6053 GND.n6052 585
R4396 GND.n1540 GND.n1539 585
R4397 GND.n6015 GND.n1540 585
R4398 GND.n5978 GND.n1569 585
R4399 GND.n5978 GND.n5977 585
R4400 GND.n5979 GND.n1568 585
R4401 GND.n5979 GND.n1555 585
R4402 GND.n5981 GND.n5980 585
R4403 GND.n5980 GND.n1553 585
R4404 GND.n5982 GND.n1566 585
R4405 GND.n1605 GND.n1566 585
R4406 GND.n5984 GND.n5983 585
R4407 GND.n5985 GND.n5984 585
R4408 GND.n1567 GND.n1565 585
R4409 GND.t82 GND.n1565 585
R4410 GND.n5931 GND.n5930 585
R4411 GND.n5931 GND.n1577 585
R4412 GND.n5933 GND.n5932 585
R4413 GND.n5932 GND.n1576 585
R4414 GND.n5934 GND.n1590 585
R4415 GND.n5918 GND.n1590 585
R4416 GND.n5936 GND.n5935 585
R4417 GND.n5937 GND.n5936 585
R4418 GND.n5929 GND.n1589 585
R4419 GND.n5924 GND.n1589 585
R4420 GND.n5928 GND.n5927 585
R4421 GND.n5927 GND.n5926 585
R4422 GND.n1592 GND.n1591 585
R4423 GND.n1621 GND.n1592 585
R4424 GND.n5892 GND.n5891 585
R4425 GND.n5891 GND.n1619 585
R4426 GND.n5893 GND.n1632 585
R4427 GND.n5879 GND.n1632 585
R4428 GND.n5895 GND.n5894 585
R4429 GND.n5896 GND.n5895 585
R4430 GND.n5890 GND.n1631 585
R4431 GND.n5885 GND.n1631 585
R4432 GND.n5889 GND.n5888 585
R4433 GND.n5888 GND.n5887 585
R4434 GND.n1634 GND.n1633 585
R4435 GND.n1649 GND.n1634 585
R4436 GND.n5849 GND.n5848 585
R4437 GND.n5848 GND.n5847 585
R4438 GND.n5850 GND.n1660 585
R4439 GND.n1663 GND.n1660 585
R4440 GND.n5852 GND.n5851 585
R4441 GND.n5853 GND.n5852 585
R4442 GND.n1661 GND.n1659 585
R4443 GND.n5839 GND.n1659 585
R4444 GND.n1692 GND.n1691 585
R4445 GND.n1691 GND.n1668 585
R4446 GND.n5811 GND.n1693 585
R4447 GND.n5811 GND.n5810 585
R4448 GND.n5812 GND.n1690 585
R4449 GND.n5812 GND.n1676 585
R4450 GND.n5814 GND.n5813 585
R4451 GND.n5813 GND.n1675 585
R4452 GND.n5815 GND.n1688 585
R4453 GND.n5781 GND.n1688 585
R4454 GND.n5817 GND.n5816 585
R4455 GND.n5818 GND.n5817 585
R4456 GND.n1689 GND.n1687 585
R4457 GND.n1687 GND.n1683 585
R4458 GND.n5769 GND.n5768 585
R4459 GND.n5770 GND.n5769 585
R4460 GND.n5767 GND.n1707 585
R4461 GND.n5763 GND.n1707 585
R4462 GND.n5766 GND.n5765 585
R4463 GND.n5765 GND.n5764 585
R4464 GND.n1709 GND.n1708 585
R4465 GND.n2076 GND.n1709 585
R4466 GND.n2065 GND.n2064 585
R4467 GND.n2064 GND.n1966 585
R4468 GND.n2067 GND.n2066 585
R4469 GND.n2068 GND.n2067 585
R4470 GND.n1948 GND.n1947 585
R4471 GND.n1951 GND.n1948 585
R4472 GND.n2086 GND.n2085 585
R4473 GND.n2085 GND.n2084 585
R4474 GND.n2087 GND.n1945 585
R4475 GND.n1945 GND.n1943 585
R4476 GND.n2089 GND.n2088 585
R4477 GND.n2090 GND.n2089 585
R4478 GND.n1946 GND.n1944 585
R4479 GND.n1944 GND.n1941 585
R4480 GND.n2052 GND.n2051 585
R4481 GND.n2053 GND.n2052 585
R4482 GND.n1930 GND.n1929 585
R4483 GND.n1933 GND.n1930 585
R4484 GND.n2100 GND.n2099 585
R4485 GND.n2099 GND.n2098 585
R4486 GND.n2101 GND.n1927 585
R4487 GND.n1927 GND.n1925 585
R4488 GND.n2103 GND.n2102 585
R4489 GND.n2104 GND.n2103 585
R4490 GND.n1928 GND.n1926 585
R4491 GND.n1926 GND.n1923 585
R4492 GND.n2039 GND.n2038 585
R4493 GND.n2040 GND.n2039 585
R4494 GND.n1912 GND.n1911 585
R4495 GND.n1915 GND.n1912 585
R4496 GND.n2114 GND.n2113 585
R4497 GND.n2113 GND.n2112 585
R4498 GND.n2115 GND.n1909 585
R4499 GND.n1909 GND.n1907 585
R4500 GND.n2117 GND.n2116 585
R4501 GND.n2118 GND.n2117 585
R4502 GND.n1910 GND.n1908 585
R4503 GND.n1908 GND.n1905 585
R4504 GND.n2026 GND.n2025 585
R4505 GND.n2027 GND.n2026 585
R4506 GND.n1894 GND.n1893 585
R4507 GND.n1897 GND.n1894 585
R4508 GND.n2128 GND.n2127 585
R4509 GND.n2127 GND.n2126 585
R4510 GND.n2129 GND.n1891 585
R4511 GND.n1891 GND.n1889 585
R4512 GND.n2131 GND.n2130 585
R4513 GND.n2132 GND.n2131 585
R4514 GND.n1892 GND.n1890 585
R4515 GND.n1890 GND.n1887 585
R4516 GND.n1875 GND.n1874 585
R4517 GND.n1878 GND.n1875 585
R4518 GND.n2142 GND.n2141 585
R4519 GND.n2141 GND.n2140 585
R4520 GND.n2143 GND.n1872 585
R4521 GND.n1876 GND.n1872 585
R4522 GND.n2145 GND.n2144 585
R4523 GND.n2146 GND.n2145 585
R4524 GND.n1873 GND.n1871 585
R4525 GND.n1871 GND.n1868 585
R4526 GND.n2005 GND.n2004 585
R4527 GND.n2006 GND.n2005 585
R4528 GND.n1856 GND.n1855 585
R4529 GND.n1860 GND.n1856 585
R4530 GND.n2156 GND.n2155 585
R4531 GND.n2155 GND.n2154 585
R4532 GND.n2157 GND.n1853 585
R4533 GND.n1858 GND.n1853 585
R4534 GND.n2159 GND.n2158 585
R4535 GND.n2160 GND.n2159 585
R4536 GND.n1854 GND.n1852 585
R4537 GND.n1852 GND.n1850 585
R4538 GND.n1992 GND.n1991 585
R4539 GND.n1993 GND.n1992 585
R4540 GND.n1839 GND.n1838 585
R4541 GND.n1842 GND.n1839 585
R4542 GND.n2170 GND.n2169 585
R4543 GND.n2169 GND.n2168 585
R4544 GND.n2171 GND.n1836 585
R4545 GND.n1840 GND.n1836 585
R4546 GND.n2173 GND.n2172 585
R4547 GND.n2174 GND.n2173 585
R4548 GND.n1837 GND.n1835 585
R4549 GND.n1835 GND.n1832 585
R4550 GND.n1980 GND.n1979 585
R4551 GND.t13 GND.n1980 585
R4552 GND.n1978 GND.n1976 585
R4553 GND.n1976 GND.n1824 585
R4554 GND.n1977 GND.n1810 585
R4555 GND.n2182 GND.n1810 585
R4556 GND.n5674 GND.n5673 585
R4557 GND.n5672 GND.n1809 585
R4558 GND.n5671 GND.n1808 585
R4559 GND.n5676 GND.n1808 585
R4560 GND.n5670 GND.n5669 585
R4561 GND.n5668 GND.n5667 585
R4562 GND.n5666 GND.n5665 585
R4563 GND.n5664 GND.n5663 585
R4564 GND.n5662 GND.n5661 585
R4565 GND.n5660 GND.n5659 585
R4566 GND.n5658 GND.n5657 585
R4567 GND.n5656 GND.n5655 585
R4568 GND.n5654 GND.n5653 585
R4569 GND.n5652 GND.n5651 585
R4570 GND.n5650 GND.n5649 585
R4571 GND.n5648 GND.n5647 585
R4572 GND.n5646 GND.n5645 585
R4573 GND.n5644 GND.n5643 585
R4574 GND.n5642 GND.n5641 585
R4575 GND.n5639 GND.n5638 585
R4576 GND.n5637 GND.n5636 585
R4577 GND.n5635 GND.n5634 585
R4578 GND.n5633 GND.n5632 585
R4579 GND.n2225 GND.n2224 585
R4580 GND.n2223 GND.n2222 585
R4581 GND.n2221 GND.n2220 585
R4582 GND.n2219 GND.n2218 585
R4583 GND.n2217 GND.n2216 585
R4584 GND.n2215 GND.n2214 585
R4585 GND.n2213 GND.n2212 585
R4586 GND.n2211 GND.n2210 585
R4587 GND.n2209 GND.n2208 585
R4588 GND.n2207 GND.n2206 585
R4589 GND.n2205 GND.n2204 585
R4590 GND.n2203 GND.n2202 585
R4591 GND.n2201 GND.n2200 585
R4592 GND.n2199 GND.n2198 585
R4593 GND.n2197 GND.n2196 585
R4594 GND.n2195 GND.n2194 585
R4595 GND.n2193 GND.n2192 585
R4596 GND.n2191 GND.n2190 585
R4597 GND.n2189 GND.n2188 585
R4598 GND.n2187 GND.n2186 585
R4599 GND.n2185 GND.n2184 585
R4600 GND.n6575 GND.n6574 585
R4601 GND.n6573 GND.n6572 585
R4602 GND.n6571 GND.n6570 585
R4603 GND.n6569 GND.n6568 585
R4604 GND.n6567 GND.n6566 585
R4605 GND.n6565 GND.n6564 585
R4606 GND.n6563 GND.n6562 585
R4607 GND.n6561 GND.n6560 585
R4608 GND.n6559 GND.n6558 585
R4609 GND.n6557 GND.n6556 585
R4610 GND.n6555 GND.n6554 585
R4611 GND.n6553 GND.n6552 585
R4612 GND.n6551 GND.n6550 585
R4613 GND.n6549 GND.n6548 585
R4614 GND.n6547 GND.n6546 585
R4615 GND.n6545 GND.n6544 585
R4616 GND.n6543 GND.n6542 585
R4617 GND.n6541 GND.n6540 585
R4618 GND.n6539 GND.n6538 585
R4619 GND.n6537 GND.n6536 585
R4620 GND.n6535 GND.n1147 585
R4621 GND.n6667 GND.n6666 585
R4622 GND.n1150 GND.n1148 585
R4623 GND.n6625 GND.n6624 585
R4624 GND.n6627 GND.n6626 585
R4625 GND.n6630 GND.n6629 585
R4626 GND.n6632 GND.n6631 585
R4627 GND.n6634 GND.n6633 585
R4628 GND.n6636 GND.n6635 585
R4629 GND.n6638 GND.n6637 585
R4630 GND.n6640 GND.n6639 585
R4631 GND.n6642 GND.n6641 585
R4632 GND.n6644 GND.n6643 585
R4633 GND.n6646 GND.n6645 585
R4634 GND.n6648 GND.n6647 585
R4635 GND.n6650 GND.n6649 585
R4636 GND.n6652 GND.n6651 585
R4637 GND.n6654 GND.n6653 585
R4638 GND.n6656 GND.n6655 585
R4639 GND.n6658 GND.n6657 585
R4640 GND.n6660 GND.n6659 585
R4641 GND.n6661 GND.n1174 585
R4642 GND.n6663 GND.n6662 585
R4643 GND.n6664 GND.n6663 585
R4644 GND.n6578 GND.n6577 585
R4645 GND.n6577 GND.n6576 585
R4646 GND.n6579 GND.n1183 585
R4647 GND.n6617 GND.n1183 585
R4648 GND.n6581 GND.n6580 585
R4649 GND.n6580 GND.n1192 585
R4650 GND.n6582 GND.n1191 585
R4651 GND.n6593 GND.n1191 585
R4652 GND.n6583 GND.n1198 585
R4653 GND.n1198 GND.n1190 585
R4654 GND.n6585 GND.n6584 585
R4655 GND.n6587 GND.n6585 585
R4656 GND.n6531 GND.n1197 585
R4657 GND.n1197 GND.n1196 585
R4658 GND.n6530 GND.n6529 585
R4659 GND.n6529 GND.n6528 585
R4660 GND.n1200 GND.n1199 585
R4661 GND.n6521 GND.n1200 585
R4662 GND.n6520 GND.n6519 585
R4663 GND.n6522 GND.n6520 585
R4664 GND.n6518 GND.n1207 585
R4665 GND.n1211 GND.n1207 585
R4666 GND.n6517 GND.n6516 585
R4667 GND.n6516 GND.n6515 585
R4668 GND.n1209 GND.n1208 585
R4669 GND.n1210 GND.n1209 585
R4670 GND.n6474 GND.n1217 585
R4671 GND.n6509 GND.n1217 585
R4672 GND.n6476 GND.n6475 585
R4673 GND.n6475 GND.n1226 585
R4674 GND.n6477 GND.n1225 585
R4675 GND.n6488 GND.n1225 585
R4676 GND.n6478 GND.n1232 585
R4677 GND.n1232 GND.n1224 585
R4678 GND.n6480 GND.n6479 585
R4679 GND.n6482 GND.n6480 585
R4680 GND.n6473 GND.n1231 585
R4681 GND.n1231 GND.n1230 585
R4682 GND.n6472 GND.n6471 585
R4683 GND.n6471 GND.n6470 585
R4684 GND.n1234 GND.n1233 585
R4685 GND.n1242 GND.n1234 585
R4686 GND.n6436 GND.n1241 585
R4687 GND.n6464 GND.n1241 585
R4688 GND.n6438 GND.n6437 585
R4689 GND.n6437 GND.n1240 585
R4690 GND.n6439 GND.n1250 585
R4691 GND.n6449 GND.n1250 585
R4692 GND.n6440 GND.n1257 585
R4693 GND.n1257 GND.n1249 585
R4694 GND.n6442 GND.n6441 585
R4695 GND.n6443 GND.n6442 585
R4696 GND.n6435 GND.n1256 585
R4697 GND.n1261 GND.n1256 585
R4698 GND.n6434 GND.n6433 585
R4699 GND.n6433 GND.n6432 585
R4700 GND.n1259 GND.n1258 585
R4701 GND.n1260 GND.n1259 585
R4702 GND.n6400 GND.n1267 585
R4703 GND.n6426 GND.n1267 585
R4704 GND.n6402 GND.n6401 585
R4705 GND.n6401 GND.n1276 585
R4706 GND.n6403 GND.n1275 585
R4707 GND.n6414 GND.n1275 585
R4708 GND.n6404 GND.n1282 585
R4709 GND.n1282 GND.n1274 585
R4710 GND.n6406 GND.n6405 585
R4711 GND.n6408 GND.n6406 585
R4712 GND.n6399 GND.n1281 585
R4713 GND.n1281 GND.n1280 585
R4714 GND.n6398 GND.n6397 585
R4715 GND.n6397 GND.n6396 585
R4716 GND.n1284 GND.n1283 585
R4717 GND.n6389 GND.n1284 585
R4718 GND.n6388 GND.n6387 585
R4719 GND.n6390 GND.n6388 585
R4720 GND.n6386 GND.n1291 585
R4721 GND.n1295 GND.n1291 585
R4722 GND.n6385 GND.n6384 585
R4723 GND.n6384 GND.n6383 585
R4724 GND.n1293 GND.n1292 585
R4725 GND.n1294 GND.n1293 585
R4726 GND.n6342 GND.n1301 585
R4727 GND.n6377 GND.n1301 585
R4728 GND.n6344 GND.n6343 585
R4729 GND.n6343 GND.n1309 585
R4730 GND.n6345 GND.n1308 585
R4731 GND.n6356 GND.n1308 585
R4732 GND.n6347 GND.n6346 585
R4733 GND.n6348 GND.n6347 585
R4734 GND.n6341 GND.n1314 585
R4735 GND.n6350 GND.n1314 585
R4736 GND.n6340 GND.n6339 585
R4737 GND.n6339 GND.n6338 585
R4738 GND.n1316 GND.n1315 585
R4739 GND.n6337 GND.n1316 585
R4740 GND.n6203 GND.n6202 585
R4741 GND.n6202 GND.n1323 585
R4742 GND.n6204 GND.n1322 585
R4743 GND.n6331 GND.n1322 585
R4744 GND.n6208 GND.n6207 585
R4745 GND.n6207 GND.n6206 585
R4746 GND.n6209 GND.n6201 585
R4747 GND.n6201 GND.n1333 585
R4748 GND.n6211 GND.n6210 585
R4749 GND.n6211 GND.n1331 585
R4750 GND.n6221 GND.n6200 585
R4751 GND.n6221 GND.n6220 585
R4752 GND.n6223 GND.n6222 585
R4753 GND.n6222 GND.n1421 585
R4754 GND.n6224 GND.n1437 585
R4755 GND.n6254 GND.n1437 585
R4756 GND.n6227 GND.n6226 585
R4757 GND.n6226 GND.n6225 585
R4758 GND.n6228 GND.n1428 585
R4759 GND.n6260 GND.n1428 585
R4760 GND.n6231 GND.n6230 585
R4761 GND.n6230 GND.n6229 585
R4762 GND.n6232 GND.n1444 585
R4763 GND.n6243 GND.n1444 585
R4764 GND.n6234 GND.n6233 585
R4765 GND.n6235 GND.n6234 585
R4766 GND.n6199 GND.n1450 585
R4767 GND.n6237 GND.n1450 585
R4768 GND.n6198 GND.n6197 585
R4769 GND.n6197 GND.n6196 585
R4770 GND.n1452 GND.n1451 585
R4771 GND.n6178 GND.n1452 585
R4772 GND.n6175 GND.n6174 585
R4773 GND.n6176 GND.n6175 585
R4774 GND.n6173 GND.n1459 585
R4775 GND.n6184 GND.n1459 585
R4776 GND.n6172 GND.n6171 585
R4777 GND.n6171 GND.n6170 585
R4778 GND.n1465 GND.n1464 585
R4779 GND.n6133 GND.n1465 585
R4780 GND.n6021 GND.n6020 585
R4781 GND.n6021 GND.n1477 585
R4782 GND.n6023 GND.n6022 585
R4783 GND.n6022 GND.n1475 585
R4784 GND.n6024 GND.n1485 585
R4785 GND.n6140 GND.n1485 585
R4786 GND.n6026 GND.n6025 585
R4787 GND.n6026 GND.n1483 585
R4788 GND.n6027 GND.n6019 585
R4789 GND.n6027 GND.n1496 585
R4790 GND.n6031 GND.n6030 585
R4791 GND.n6030 GND.t1 585
R4792 GND.n6032 GND.n1504 585
R4793 GND.n6096 GND.n1504 585
R4794 GND.n6034 GND.n6033 585
R4795 GND.n6033 GND.n1502 585
R4796 GND.n6035 GND.n1511 585
R4797 GND.n6087 GND.n1511 585
R4798 GND.n6039 GND.n6038 585
R4799 GND.n6038 GND.n6037 585
R4800 GND.n6040 GND.n1519 585
R4801 GND.n6075 GND.n1519 585
R4802 GND.n6042 GND.n6041 585
R4803 GND.n6041 GND.n1518 585
R4804 GND.n6043 GND.n1525 585
R4805 GND.n6069 GND.n1525 585
R4806 GND.n6046 GND.n6045 585
R4807 GND.n6045 GND.n6044 585
R4808 GND.n6047 GND.n1535 585
R4809 GND.n6058 GND.n1535 585
R4810 GND.n6049 GND.n6048 585
R4811 GND.n6050 GND.n6049 585
R4812 GND.n6018 GND.n1542 585
R4813 GND.n6052 GND.n1542 585
R4814 GND.n6017 GND.n6016 585
R4815 GND.n6016 GND.n6015 585
R4816 GND.n1545 GND.n1544 585
R4817 GND.n5977 GND.n1545 585
R4818 GND.n1602 GND.n1601 585
R4819 GND.n1602 GND.n1555 585
R4820 GND.n1603 GND.n1600 585
R4821 GND.n1603 GND.n1553 585
R4822 GND.n1607 GND.n1606 585
R4823 GND.n1606 GND.n1605 585
R4824 GND.n1608 GND.n1563 585
R4825 GND.n5985 GND.n1563 585
R4826 GND.n1609 GND.n1599 585
R4827 GND.n1599 GND.t82 585
R4828 GND.n1611 GND.n1610 585
R4829 GND.n1611 GND.n1577 585
R4830 GND.n1612 GND.n1597 585
R4831 GND.n1612 GND.n1576 585
R4832 GND.n5920 GND.n5919 585
R4833 GND.n5919 GND.n5918 585
R4834 GND.n5921 GND.n1587 585
R4835 GND.n5937 GND.n1587 585
R4836 GND.n5923 GND.n5922 585
R4837 GND.n5924 GND.n5923 585
R4838 GND.n1596 GND.n1594 585
R4839 GND.n5926 GND.n1594 585
R4840 GND.n1641 GND.n1640 585
R4841 GND.n1641 GND.n1621 585
R4842 GND.n1642 GND.n1639 585
R4843 GND.n1642 GND.n1619 585
R4844 GND.n5881 GND.n5880 585
R4845 GND.n5880 GND.n5879 585
R4846 GND.n5882 GND.n1629 585
R4847 GND.n5896 GND.n1629 585
R4848 GND.n5884 GND.n5883 585
R4849 GND.n5885 GND.n5884 585
R4850 GND.n1638 GND.n1636 585
R4851 GND.n5887 GND.n1636 585
R4852 GND.n5844 GND.n1665 585
R4853 GND.n1665 GND.n1649 585
R4854 GND.n5846 GND.n5845 585
R4855 GND.n5847 GND.n5846 585
R4856 GND.n5843 GND.n1664 585
R4857 GND.n1664 GND.n1663 585
R4858 GND.n5842 GND.n1656 585
R4859 GND.n5853 GND.n1656 585
R4860 GND.n5841 GND.n5840 585
R4861 GND.n5840 GND.n5839 585
R4862 GND.n1667 GND.n1666 585
R4863 GND.n1668 GND.n1667 585
R4864 GND.n5775 GND.n1695 585
R4865 GND.n5810 GND.n1695 585
R4866 GND.n5777 GND.n5776 585
R4867 GND.n5776 GND.n1676 585
R4868 GND.n5778 GND.n1702 585
R4869 GND.n1702 GND.n1675 585
R4870 GND.n5780 GND.n5779 585
R4871 GND.n5781 GND.n5780 585
R4872 GND.n5774 GND.n1685 585
R4873 GND.n5818 GND.n1685 585
R4874 GND.n5773 GND.n5772 585
R4875 GND.n5772 GND.n1683 585
R4876 GND.n5771 GND.n1703 585
R4877 GND.n5771 GND.n5770 585
R4878 GND.n2072 GND.n1704 585
R4879 GND.n5763 GND.n1704 585
R4880 GND.n2073 GND.n1711 585
R4881 GND.n5764 GND.n1711 585
R4882 GND.n2075 GND.n2074 585
R4883 GND.n2076 GND.n2075 585
R4884 GND.n2071 GND.n1967 585
R4885 GND.n1967 GND.n1966 585
R4886 GND.n2070 GND.n2069 585
R4887 GND.n2069 GND.n2068 585
R4888 GND.n2062 GND.n2061 585
R4889 GND.n2062 GND.n1951 585
R4890 GND.n2060 GND.n1950 585
R4891 GND.n2084 GND.n1950 585
R4892 GND.n2059 GND.n2058 585
R4893 GND.n2058 GND.n1943 585
R4894 GND.n2057 GND.n1942 585
R4895 GND.n2090 GND.n1942 585
R4896 GND.n2056 GND.n2055 585
R4897 GND.n2055 GND.n1941 585
R4898 GND.n2054 GND.n1968 585
R4899 GND.n2054 GND.n2053 585
R4900 GND.n2049 GND.n2048 585
R4901 GND.n2049 GND.n1933 585
R4902 GND.n2047 GND.n1932 585
R4903 GND.n2098 GND.n1932 585
R4904 GND.n2046 GND.n2045 585
R4905 GND.n2045 GND.n1925 585
R4906 GND.n2044 GND.n1924 585
R4907 GND.n2104 GND.n1924 585
R4908 GND.n2043 GND.n2042 585
R4909 GND.n2042 GND.n1923 585
R4910 GND.n2041 GND.n1969 585
R4911 GND.n2041 GND.n2040 585
R4912 GND.n2036 GND.n2035 585
R4913 GND.n2036 GND.n1915 585
R4914 GND.n2034 GND.n1914 585
R4915 GND.n2112 GND.n1914 585
R4916 GND.n2033 GND.n2032 585
R4917 GND.n2032 GND.n1907 585
R4918 GND.n2031 GND.n1906 585
R4919 GND.n2118 GND.n1906 585
R4920 GND.n2030 GND.n2029 585
R4921 GND.n2029 GND.n1905 585
R4922 GND.n2028 GND.n1970 585
R4923 GND.n2028 GND.n2027 585
R4924 GND.n2023 GND.n2022 585
R4925 GND.n2023 GND.n1897 585
R4926 GND.n2021 GND.n1896 585
R4927 GND.n2126 GND.n1896 585
R4928 GND.n2020 GND.n2019 585
R4929 GND.n2019 GND.n1889 585
R4930 GND.n2018 GND.n1888 585
R4931 GND.n2132 GND.n1888 585
R4932 GND.n2017 GND.n2016 585
R4933 GND.n2016 GND.n1887 585
R4934 GND.n2015 GND.n2014 585
R4935 GND.n2015 GND.n1878 585
R4936 GND.n2013 GND.n1877 585
R4937 GND.n2140 GND.n1877 585
R4938 GND.n2012 GND.n2011 585
R4939 GND.n2011 GND.n1876 585
R4940 GND.n2010 GND.n1869 585
R4941 GND.n2146 GND.n1869 585
R4942 GND.n2009 GND.n2008 585
R4943 GND.n2008 GND.n1868 585
R4944 GND.n2007 GND.n1971 585
R4945 GND.n2007 GND.n2006 585
R4946 GND.n2002 GND.n2001 585
R4947 GND.n2002 GND.n1860 585
R4948 GND.n2000 GND.n1859 585
R4949 GND.n2154 GND.n1859 585
R4950 GND.n1999 GND.n1998 585
R4951 GND.n1998 GND.n1858 585
R4952 GND.n1997 GND.n1851 585
R4953 GND.n2160 GND.n1851 585
R4954 GND.n1996 GND.n1995 585
R4955 GND.n1995 GND.n1850 585
R4956 GND.n1994 GND.n1972 585
R4957 GND.n1994 GND.n1993 585
R4958 GND.n1989 GND.n1988 585
R4959 GND.n1989 GND.n1842 585
R4960 GND.n1987 GND.n1841 585
R4961 GND.n2168 GND.n1841 585
R4962 GND.n1986 GND.n1985 585
R4963 GND.n1985 GND.n1840 585
R4964 GND.n1984 GND.n1833 585
R4965 GND.n2174 GND.n1833 585
R4966 GND.n1983 GND.n1982 585
R4967 GND.n1982 GND.n1832 585
R4968 GND.n1981 GND.n1974 585
R4969 GND.n1981 GND.t13 585
R4970 GND.n1973 GND.n1823 585
R4971 GND.n1824 GND.n1823 585
R4972 GND.n2183 GND.n1822 585
R4973 GND.n2183 GND.n2182 585
R4974 GND.n4191 GND.n4190 585
R4975 GND.n4191 GND.n307 585
R4976 GND.n295 GND.n294 585
R4977 GND.n298 GND.n295 585
R4978 GND.n7610 GND.n7609 585
R4979 GND.n7609 GND.n7608 585
R4980 GND.n7611 GND.n289 585
R4981 GND.n289 GND.n287 585
R4982 GND.n7613 GND.n7612 585
R4983 GND.n7614 GND.n7613 585
R4984 GND.n274 GND.n273 585
R4985 GND.n277 GND.n274 585
R4986 GND.n7622 GND.n7621 585
R4987 GND.n7621 GND.n7620 585
R4988 GND.n7623 GND.n269 585
R4989 GND.n269 GND.n267 585
R4990 GND.n7625 GND.n7624 585
R4991 GND.n7626 GND.n7625 585
R4992 GND.n251 GND.n249 585
R4993 GND.n264 GND.n251 585
R4994 GND.n7634 GND.n7633 585
R4995 GND.n7633 GND.n7632 585
R4996 GND.n250 GND.n248 585
R4997 GND.n252 GND.n250 585
R4998 GND.n7207 GND.n7206 585
R4999 GND.n7208 GND.n7207 585
R5000 GND.n7205 GND.n241 585
R5001 GND.n7205 GND.n619 585
R5002 GND.n7638 GND.n239 585
R5003 GND.n239 GND.n236 585
R5004 GND.n7640 GND.n7639 585
R5005 GND.n7641 GND.n7640 585
R5006 GND.n7165 GND.n238 585
R5007 GND.n238 GND.n233 585
R5008 GND.n7167 GND.n7166 585
R5009 GND.n7168 GND.n7167 585
R5010 GND.n7164 GND.n7163 585
R5011 GND.n7164 GND.n630 585
R5012 GND.n7162 GND.n7161 585
R5013 GND.n7161 GND.n7160 585
R5014 GND.n7142 GND.n634 585
R5015 GND.n635 GND.n634 585
R5016 GND.n7144 GND.n7143 585
R5017 GND.n7145 GND.n7144 585
R5018 GND.n7141 GND.n648 585
R5019 GND.n7129 GND.n648 585
R5020 GND.n653 GND.n649 585
R5021 GND.n657 GND.n653 585
R5022 GND.n7137 GND.n7136 585
R5023 GND.n7136 GND.n7135 585
R5024 GND.n652 GND.n651 585
R5025 GND.n654 GND.n652 585
R5026 GND.n7106 GND.n7105 585
R5027 GND.n7107 GND.n7106 585
R5028 GND.n678 GND.n677 585
R5029 GND.n677 GND.n673 585
R5030 GND.n7101 GND.n7100 585
R5031 GND.n7100 GND.n7099 585
R5032 GND.n681 GND.n680 585
R5033 GND.n682 GND.n681 585
R5034 GND.n7078 GND.n7077 585
R5035 GND.n7079 GND.n7078 585
R5036 GND.n699 GND.n698 585
R5037 GND.n698 GND.n694 585
R5038 GND.n7073 GND.n7072 585
R5039 GND.n7072 GND.n7071 585
R5040 GND.n702 GND.n701 585
R5041 GND.n7060 GND.n702 585
R5042 GND.n7034 GND.n725 585
R5043 GND.n725 GND.n713 585
R5044 GND.n7036 GND.n7035 585
R5045 GND.n7037 GND.n7036 585
R5046 GND.n726 GND.n724 585
R5047 GND.n724 GND.n720 585
R5048 GND.n7029 GND.n7028 585
R5049 GND.n7028 GND.n7027 585
R5050 GND.n729 GND.n728 585
R5051 GND.n730 GND.n729 585
R5052 GND.n7010 GND.n7009 585
R5053 GND.n7011 GND.n7010 585
R5054 GND.n747 GND.n746 585
R5055 GND.n746 GND.n742 585
R5056 GND.n7005 GND.n7004 585
R5057 GND.n7004 GND.n7003 585
R5058 GND.n750 GND.n749 585
R5059 GND.n751 GND.n750 585
R5060 GND.n6990 GND.n6989 585
R5061 GND.n6991 GND.n6990 585
R5062 GND.n767 GND.n766 585
R5063 GND.n766 GND.n762 585
R5064 GND.n6985 GND.n6984 585
R5065 GND.n6984 GND.n6983 585
R5066 GND.n770 GND.n769 585
R5067 GND.n771 GND.n770 585
R5068 GND.n6970 GND.n6969 585
R5069 GND.n6971 GND.n6970 585
R5070 GND.n787 GND.n786 585
R5071 GND.n786 GND.n782 585
R5072 GND.n6965 GND.n6964 585
R5073 GND.n6964 GND.n6963 585
R5074 GND.n790 GND.n789 585
R5075 GND.n791 GND.n790 585
R5076 GND.n6950 GND.n6949 585
R5077 GND.n6951 GND.n6950 585
R5078 GND.n807 GND.n806 585
R5079 GND.n806 GND.n802 585
R5080 GND.n6945 GND.n6944 585
R5081 GND.n6944 GND.n6943 585
R5082 GND.n810 GND.n809 585
R5083 GND.n811 GND.n810 585
R5084 GND.n6930 GND.n6929 585
R5085 GND.n6931 GND.n6930 585
R5086 GND.n826 GND.n825 585
R5087 GND.n833 GND.n825 585
R5088 GND.n6925 GND.n6924 585
R5089 GND.n6924 GND.n6923 585
R5090 GND.n829 GND.n828 585
R5091 GND.n830 GND.n829 585
R5092 GND.n6910 GND.n6909 585
R5093 GND.n6911 GND.n6910 585
R5094 GND.n847 GND.n846 585
R5095 GND.n846 GND.n842 585
R5096 GND.n6905 GND.n6904 585
R5097 GND.n6904 GND.n6903 585
R5098 GND.n850 GND.n849 585
R5099 GND.n851 GND.n850 585
R5100 GND.n6890 GND.n6889 585
R5101 GND.n6891 GND.n6890 585
R5102 GND.n867 GND.n866 585
R5103 GND.n866 GND.n862 585
R5104 GND.n6885 GND.n6884 585
R5105 GND.n6884 GND.n6883 585
R5106 GND.n870 GND.n869 585
R5107 GND.n871 GND.n870 585
R5108 GND.n6870 GND.n6869 585
R5109 GND.n6871 GND.n6870 585
R5110 GND.n887 GND.n886 585
R5111 GND.n886 GND.n882 585
R5112 GND.n6865 GND.n6864 585
R5113 GND.n6864 GND.n6863 585
R5114 GND.n890 GND.n889 585
R5115 GND.n6852 GND.n890 585
R5116 GND.n6759 GND.n913 585
R5117 GND.n913 GND.n901 585
R5118 GND.n6761 GND.n6760 585
R5119 GND.n6762 GND.n6761 585
R5120 GND.n914 GND.n912 585
R5121 GND.n912 GND.n908 585
R5122 GND.n6754 GND.n6753 585
R5123 GND.n6753 GND.n6752 585
R5124 GND.n917 GND.n916 585
R5125 GND.n918 GND.n917 585
R5126 GND.n6733 GND.n6732 585
R5127 GND.n6734 GND.n6733 585
R5128 GND.n936 GND.n935 585
R5129 GND.n935 GND.n931 585
R5130 GND.n6728 GND.n6727 585
R5131 GND.n6727 GND.n6726 585
R5132 GND.n939 GND.n938 585
R5133 GND.n940 GND.n939 585
R5134 GND.n6607 GND.n6606 585
R5135 GND.n6608 GND.n6607 585
R5136 GND.n6603 GND.n6602 585
R5137 GND.n6609 GND.n6603 585
R5138 GND.n6612 GND.n6611 585
R5139 GND.n6611 GND.n6610 585
R5140 GND.n6613 GND.n1185 585
R5141 GND.n1185 GND.n1151 585
R5142 GND.n6615 GND.n6614 585
R5143 GND.n6616 GND.n6615 585
R5144 GND.n1186 GND.n1184 585
R5145 GND.n1184 GND.n1182 585
R5146 GND.n6596 GND.n6595 585
R5147 GND.n6595 GND.n6594 585
R5148 GND.n1189 GND.n1188 585
R5149 GND.n6586 GND.n1189 585
R5150 GND.n6501 GND.n6500 585
R5151 GND.n6501 GND.n1202 585
R5152 GND.n6502 GND.n6497 585
R5153 GND.n6502 GND.n1201 585
R5154 GND.n6504 GND.n6503 585
R5155 GND.n6503 GND.n1206 585
R5156 GND.n6505 GND.n1219 585
R5157 GND.n1219 GND.n1212 585
R5158 GND.n6507 GND.n6506 585
R5159 GND.n6508 GND.n6507 585
R5160 GND.n1220 GND.n1218 585
R5161 GND.n1218 GND.n1216 585
R5162 GND.n6491 GND.n6490 585
R5163 GND.n6490 GND.n6489 585
R5164 GND.n1223 GND.n1222 585
R5165 GND.n6481 GND.n1223 585
R5166 GND.n6459 GND.n6458 585
R5167 GND.n6458 GND.n1236 585
R5168 GND.n6460 GND.n1244 585
R5169 GND.n1244 GND.n1235 585
R5170 GND.n6462 GND.n6461 585
R5171 GND.n6463 GND.n6462 585
R5172 GND.n1245 GND.n1243 585
R5173 GND.n1251 GND.n1243 585
R5174 GND.n6452 GND.n6451 585
R5175 GND.n6451 GND.n6450 585
R5176 GND.n1248 GND.n1247 585
R5177 GND.n1255 GND.n1248 585
R5178 GND.n6422 GND.n1269 585
R5179 GND.n1269 GND.n1262 585
R5180 GND.n6424 GND.n6423 585
R5181 GND.n6425 GND.n6424 585
R5182 GND.n1270 GND.n1268 585
R5183 GND.n1268 GND.n1266 585
R5184 GND.n6417 GND.n6416 585
R5185 GND.n6416 GND.n6415 585
R5186 GND.n1273 GND.n1272 585
R5187 GND.n6407 GND.n1273 585
R5188 GND.n6369 GND.n6368 585
R5189 GND.n6369 GND.n1286 585
R5190 GND.n6370 GND.n6365 585
R5191 GND.n6370 GND.n1285 585
R5192 GND.n6372 GND.n6371 585
R5193 GND.n6371 GND.n1290 585
R5194 GND.n6373 GND.n1303 585
R5195 GND.n1303 GND.n1296 585
R5196 GND.n6375 GND.n6374 585
R5197 GND.n6376 GND.n6375 585
R5198 GND.n1304 GND.n1302 585
R5199 GND.n1302 GND.n1300 585
R5200 GND.n6359 GND.n6358 585
R5201 GND.n6358 GND.n6357 585
R5202 GND.n1307 GND.n1306 585
R5203 GND.n6349 GND.n1307 585
R5204 GND.n6326 GND.n6325 585
R5205 GND.n6325 GND.n1313 585
R5206 GND.n6327 GND.n1326 585
R5207 GND.n1326 GND.n1325 585
R5208 GND.n6329 GND.n6328 585
R5209 GND.n6330 GND.n6329 585
R5210 GND.n1327 GND.n1324 585
R5211 GND.n6205 GND.n1324 585
R5212 GND.n6319 GND.n6318 585
R5213 GND.n6318 GND.n6317 585
R5214 GND.n1330 GND.n1329 585
R5215 GND.n6212 GND.n1330 585
R5216 GND.n6252 GND.n6251 585
R5217 GND.n6253 GND.n6252 585
R5218 GND.n1439 GND.n1438 585
R5219 GND.n1438 GND.n1430 585
R5220 GND.n6247 GND.n6246 585
R5221 GND.n6246 GND.n1427 585
R5222 GND.n6245 GND.n1441 585
R5223 GND.n6245 GND.n6244 585
R5224 GND.n6192 GND.n1442 585
R5225 GND.n6236 GND.n1442 585
R5226 GND.n6194 GND.n6193 585
R5227 GND.n6195 GND.n6194 585
R5228 GND.n1455 GND.n1454 585
R5229 GND.n6177 GND.n1454 585
R5230 GND.n6187 GND.n6186 585
R5231 GND.n6186 GND.n6185 585
R5232 GND.n1458 GND.n1457 585
R5233 GND.n1466 GND.n1458 585
R5234 GND.n6149 GND.n6148 585
R5235 GND.n6150 GND.n6149 585
R5236 GND.n1479 GND.n1478 585
R5237 GND.n1486 GND.n1478 585
R5238 GND.n6144 GND.n6143 585
R5239 GND.n6143 GND.n6142 585
R5240 GND.n1482 GND.n1481 585
R5241 GND.n6029 GND.n1482 585
R5242 GND.n6083 GND.n1513 585
R5243 GND.n1513 GND.n1505 585
R5244 GND.n6085 GND.n6084 585
R5245 GND.n6086 GND.n6085 585
R5246 GND.n1514 GND.n1512 585
R5247 GND.n6036 GND.n1512 585
R5248 GND.n6078 GND.n6077 585
R5249 GND.n6077 GND.n6076 585
R5250 GND.n1517 GND.n1516 585
R5251 GND.n6068 GND.n1517 585
R5252 GND.n5998 GND.n5997 585
R5253 GND.n5998 GND.n1537 585
R5254 GND.n5999 GND.n5994 585
R5255 GND.n5999 GND.n1534 585
R5256 GND.n6001 GND.n6000 585
R5257 GND.n6000 GND.n1541 585
R5258 GND.n6002 GND.n1557 585
R5259 GND.n1557 GND.n1546 585
R5260 GND.n6004 GND.n6003 585
R5261 GND.n6005 GND.n6004 585
R5262 GND.n1558 GND.n1556 585
R5263 GND.n1604 GND.n1556 585
R5264 GND.n5988 GND.n5987 585
R5265 GND.n5987 GND.n5986 585
R5266 GND.n1561 GND.n1560 585
R5267 GND.n1598 GND.n1561 585
R5268 GND.n5915 GND.n5914 585
R5269 GND.n5916 GND.n5915 585
R5270 GND.n1614 GND.n1613 585
R5271 GND.n1613 GND.n1588 585
R5272 GND.n5910 GND.n5909 585
R5273 GND.n5909 GND.n1585 585
R5274 GND.n5908 GND.n1616 585
R5275 GND.n5908 GND.n1593 585
R5276 GND.n5907 GND.n1618 585
R5277 GND.n5907 GND.n5906 585
R5278 GND.n5798 GND.n1617 585
R5279 GND.n1630 GND.n1617 585
R5280 GND.n5799 GND.n5792 585
R5281 GND.n5792 GND.n1627 585
R5282 GND.n5801 GND.n5800 585
R5283 GND.n5801 GND.n1635 585
R5284 GND.n5802 GND.n5791 585
R5285 GND.n5802 GND.n1648 585
R5286 GND.n5804 GND.n5803 585
R5287 GND.n5803 GND.n1658 585
R5288 GND.n5805 GND.n1697 585
R5289 GND.n1697 GND.n1655 585
R5290 GND.n5807 GND.n5806 585
R5291 GND.n5808 GND.n5807 585
R5292 GND.n1698 GND.n1696 585
R5293 GND.n1696 GND.n1694 585
R5294 GND.n5785 GND.n5784 585
R5295 GND.n5784 GND.n5783 585
R5296 GND.n1701 GND.n1700 585
R5297 GND.n1701 GND.n1686 585
R5298 GND.n1962 GND.n1958 585
R5299 GND.n1958 GND.n1706 585
R5300 GND.n1964 GND.n1963 585
R5301 GND.n1964 GND.n1705 585
R5302 GND.n1965 GND.n1957 585
R5303 GND.n1965 GND.n1710 585
R5304 GND.n2079 GND.n2078 585
R5305 GND.n2078 GND.n2077 585
R5306 GND.n2080 GND.n1952 585
R5307 GND.n2063 GND.n1952 585
R5308 GND.n2082 GND.n2081 585
R5309 GND.n2083 GND.n2082 585
R5310 GND.n1940 GND.n1939 585
R5311 GND.n1949 GND.n1940 585
R5312 GND.n2093 GND.n2092 585
R5313 GND.n2092 GND.n2091 585
R5314 GND.n2094 GND.n1934 585
R5315 GND.n2050 GND.n1934 585
R5316 GND.n2096 GND.n2095 585
R5317 GND.n2097 GND.n2096 585
R5318 GND.n1922 GND.n1921 585
R5319 GND.n1931 GND.n1922 585
R5320 GND.n2107 GND.n2106 585
R5321 GND.n2106 GND.n2105 585
R5322 GND.n2108 GND.n1916 585
R5323 GND.n2037 GND.n1916 585
R5324 GND.n2110 GND.n2109 585
R5325 GND.n2111 GND.n2110 585
R5326 GND.n1904 GND.n1903 585
R5327 GND.n1913 GND.n1904 585
R5328 GND.n2121 GND.n2120 585
R5329 GND.n2120 GND.n2119 585
R5330 GND.n2122 GND.n1898 585
R5331 GND.n2024 GND.n1898 585
R5332 GND.n2124 GND.n2123 585
R5333 GND.n2125 GND.n2124 585
R5334 GND.n1885 GND.n1884 585
R5335 GND.n1895 GND.n1885 585
R5336 GND.n2135 GND.n2134 585
R5337 GND.n2134 GND.n2133 585
R5338 GND.n2136 GND.n1879 585
R5339 GND.n1886 GND.n1879 585
R5340 GND.n2138 GND.n2137 585
R5341 GND.n2139 GND.n2138 585
R5342 GND.n1867 GND.n1866 585
R5343 GND.n1870 GND.n1867 585
R5344 GND.n2149 GND.n2148 585
R5345 GND.n2148 GND.n2147 585
R5346 GND.n2150 GND.n1861 585
R5347 GND.n2003 GND.n1861 585
R5348 GND.n2152 GND.n2151 585
R5349 GND.n2153 GND.n2152 585
R5350 GND.n1849 GND.n1848 585
R5351 GND.n1857 GND.n1849 585
R5352 GND.n2163 GND.n2162 585
R5353 GND.n2162 GND.n2161 585
R5354 GND.n2164 GND.n1843 585
R5355 GND.n1990 GND.n1843 585
R5356 GND.n2166 GND.n2165 585
R5357 GND.n2167 GND.n2166 585
R5358 GND.n1831 GND.n1830 585
R5359 GND.n1834 GND.n1831 585
R5360 GND.n2177 GND.n2176 585
R5361 GND.n2176 GND.n2175 585
R5362 GND.n2178 GND.n1825 585
R5363 GND.n1975 GND.n1825 585
R5364 GND.n2180 GND.n2179 585
R5365 GND.n2181 GND.n2180 585
R5366 GND.n1785 GND.n1784 585
R5367 GND.n1807 GND.n1785 585
R5368 GND.n5679 GND.n5678 585
R5369 GND.n5678 GND.n5677 585
R5370 GND.n5680 GND.n1779 585
R5371 GND.n1779 GND.n1778 585
R5372 GND.n5682 GND.n5681 585
R5373 GND.n5683 GND.n5682 585
R5374 GND.n1749 GND.n1748 585
R5375 GND.n5684 GND.n1749 585
R5376 GND.n5687 GND.n5686 585
R5377 GND.n5686 GND.n5685 585
R5378 GND.n5688 GND.n1743 585
R5379 GND.n1743 GND.n1740 585
R5380 GND.n5690 GND.n5689 585
R5381 GND.n5691 GND.n5690 585
R5382 GND.n1744 GND.n1742 585
R5383 GND.n1742 GND.n1737 585
R5384 GND.n5558 GND.n5557 585
R5385 GND.n5559 GND.n5558 585
R5386 GND.n2244 GND.n2243 585
R5387 GND.n2243 GND.n2239 585
R5388 GND.n5552 GND.n5551 585
R5389 GND.n5551 GND.n5550 585
R5390 GND.n2247 GND.n2246 585
R5391 GND.n2248 GND.n2247 585
R5392 GND.n5533 GND.n5532 585
R5393 GND.n5534 GND.n5533 585
R5394 GND.n2263 GND.n2262 585
R5395 GND.n2270 GND.n2262 585
R5396 GND.n5528 GND.n5527 585
R5397 GND.n5527 GND.n5526 585
R5398 GND.n2266 GND.n2265 585
R5399 GND.n2267 GND.n2266 585
R5400 GND.n5513 GND.n5512 585
R5401 GND.n5514 GND.n5513 585
R5402 GND.n2284 GND.n2283 585
R5403 GND.n2283 GND.n2279 585
R5404 GND.n5508 GND.n5507 585
R5405 GND.n5507 GND.n5506 585
R5406 GND.n2287 GND.n2286 585
R5407 GND.n2288 GND.n2287 585
R5408 GND.n5493 GND.n5492 585
R5409 GND.n5494 GND.n5493 585
R5410 GND.n2304 GND.n2303 585
R5411 GND.n2303 GND.n2299 585
R5412 GND.n5488 GND.n5487 585
R5413 GND.n5487 GND.n5486 585
R5414 GND.n2307 GND.n2306 585
R5415 GND.n2308 GND.n2307 585
R5416 GND.n5473 GND.n5472 585
R5417 GND.n5474 GND.n5473 585
R5418 GND.n2324 GND.n2323 585
R5419 GND.n2323 GND.n2319 585
R5420 GND.n5468 GND.n5467 585
R5421 GND.n5467 GND.n5466 585
R5422 GND.n2327 GND.n2326 585
R5423 GND.n5455 GND.n2327 585
R5424 GND.n5393 GND.n2350 585
R5425 GND.n2350 GND.n2338 585
R5426 GND.n5395 GND.n5394 585
R5427 GND.n5396 GND.n5395 585
R5428 GND.n2351 GND.n2349 585
R5429 GND.n2349 GND.n2345 585
R5430 GND.n5388 GND.n5387 585
R5431 GND.n5387 GND.n5386 585
R5432 GND.n2354 GND.n2353 585
R5433 GND.n2355 GND.n2354 585
R5434 GND.n5368 GND.n5367 585
R5435 GND.n5369 GND.n5368 585
R5436 GND.n2371 GND.n2370 585
R5437 GND.n2370 GND.n2366 585
R5438 GND.n5363 GND.n5362 585
R5439 GND.n5362 GND.n5361 585
R5440 GND.n2374 GND.n2373 585
R5441 GND.n2375 GND.n2374 585
R5442 GND.n5348 GND.n5347 585
R5443 GND.n5349 GND.n5348 585
R5444 GND.n2390 GND.n2389 585
R5445 GND.n2397 GND.n2389 585
R5446 GND.n5343 GND.n5342 585
R5447 GND.n5342 GND.n5341 585
R5448 GND.n2393 GND.n2392 585
R5449 GND.n2394 GND.n2393 585
R5450 GND.n5328 GND.n5327 585
R5451 GND.n5329 GND.n5328 585
R5452 GND.n2411 GND.n2410 585
R5453 GND.n2410 GND.n2406 585
R5454 GND.n5323 GND.n5322 585
R5455 GND.n5322 GND.n5321 585
R5456 GND.n2414 GND.n2413 585
R5457 GND.n2415 GND.n2414 585
R5458 GND.n5308 GND.n5307 585
R5459 GND.n5309 GND.n5308 585
R5460 GND.n2431 GND.n2430 585
R5461 GND.n2430 GND.n2426 585
R5462 GND.n5303 GND.n5302 585
R5463 GND.n5302 GND.n5301 585
R5464 GND.n2434 GND.n2433 585
R5465 GND.n2435 GND.n2434 585
R5466 GND.n5288 GND.n5287 585
R5467 GND.n5289 GND.n5288 585
R5468 GND.n2450 GND.n2449 585
R5469 GND.n2457 GND.n2449 585
R5470 GND.n5283 GND.n5282 585
R5471 GND.n5282 GND.n5281 585
R5472 GND.n2453 GND.n2452 585
R5473 GND.n2454 GND.n2453 585
R5474 GND.n5268 GND.n5267 585
R5475 GND.n5269 GND.n5268 585
R5476 GND.n2471 GND.n2470 585
R5477 GND.n2470 GND.n2466 585
R5478 GND.n5263 GND.n5262 585
R5479 GND.n5262 GND.n5261 585
R5480 GND.n2474 GND.n2473 585
R5481 GND.n2475 GND.n2474 585
R5482 GND.n5248 GND.n5247 585
R5483 GND.n5249 GND.n5248 585
R5484 GND.n2491 GND.n2490 585
R5485 GND.n2490 GND.n2486 585
R5486 GND.n5243 GND.n5242 585
R5487 GND.n5242 GND.n5241 585
R5488 GND.n2494 GND.n2493 585
R5489 GND.n2495 GND.n2494 585
R5490 GND.n5228 GND.n5227 585
R5491 GND.n5229 GND.n5228 585
R5492 GND.n2511 GND.n2510 585
R5493 GND.n2510 GND.n2506 585
R5494 GND.n5181 GND.n5180 585
R5495 GND.n5182 GND.n5181 585
R5496 GND.n5179 GND.n5178 585
R5497 GND.n5179 GND.n2577 585
R5498 GND.n5177 GND.n5176 585
R5499 GND.n5176 GND.n5175 585
R5500 GND.n5079 GND.n2713 585
R5501 GND.n2715 GND.n2713 585
R5502 GND.n5081 GND.n5080 585
R5503 GND.n5082 GND.n5081 585
R5504 GND.n5078 GND.n5077 585
R5505 GND.n5078 GND.n2727 585
R5506 GND.n5076 GND.n2516 585
R5507 GND.n5076 GND.n5075 585
R5508 GND.n2735 GND.n2734 585
R5509 GND.n2737 GND.n2735 585
R5510 GND.n5217 GND.n2534 585
R5511 GND.n2534 GND.n2530 585
R5512 GND.n5219 GND.n5218 585
R5513 GND.n5220 GND.n5219 585
R5514 GND.n5216 GND.n2533 585
R5515 GND.n2757 GND.n2533 585
R5516 GND.n2539 GND.n2535 585
R5517 GND.n2543 GND.n2539 585
R5518 GND.n5212 GND.n5211 585
R5519 GND.n5211 GND.n5210 585
R5520 GND.n2538 GND.n2537 585
R5521 GND.n2540 GND.n2538 585
R5522 GND.n5057 GND.n5056 585
R5523 GND.n5058 GND.n5057 585
R5524 GND.n2767 GND.n2766 585
R5525 GND.n2766 GND.n2762 585
R5526 GND.n5052 GND.n5051 585
R5527 GND.n5051 GND.n5050 585
R5528 GND.n2770 GND.n2769 585
R5529 GND.n2771 GND.n2770 585
R5530 GND.n5033 GND.n5032 585
R5531 GND.n5034 GND.n5033 585
R5532 GND.n6278 GND.n6277 585
R5533 GND.n6277 GND.n1317 585
R5534 GND.n1415 GND.n1412 585
R5535 GND.n6282 GND.n1411 585
R5536 GND.n6283 GND.n1410 585
R5537 GND.n6285 GND.n1406 585
R5538 GND.n1405 GND.n1402 585
R5539 GND.n6289 GND.n1401 585
R5540 GND.n6290 GND.n1400 585
R5541 GND.n6291 GND.n1398 585
R5542 GND.n1397 GND.n1394 585
R5543 GND.n6295 GND.n1393 585
R5544 GND.n6296 GND.n1392 585
R5545 GND.n6297 GND.n1390 585
R5546 GND.n1389 GND.n1386 585
R5547 GND.n6301 GND.n1385 585
R5548 GND.n6302 GND.n1384 585
R5549 GND.n6303 GND.n1382 585
R5550 GND.n1381 GND.n1344 585
R5551 GND.n6308 GND.n1343 585
R5552 GND.n6309 GND.n1342 585
R5553 GND.n6310 GND.n1340 585
R5554 GND.n6276 GND.n6275 585
R5555 GND.n6276 GND.n1321 585
R5556 GND.n6274 GND.n1332 585
R5557 GND.n6316 GND.n1332 585
R5558 GND.n1420 GND.n1416 585
R5559 GND.n6213 GND.n1420 585
R5560 GND.n6270 GND.n6269 585
R5561 GND.n6269 GND.n6268 585
R5562 GND.n1419 GND.n1418 585
R5563 GND.n1436 GND.n1419 585
R5564 GND.n6119 GND.n1429 585
R5565 GND.n6260 GND.n1429 585
R5566 GND.n6120 GND.n6118 585
R5567 GND.n6118 GND.n1445 585
R5568 GND.n6117 GND.n6115 585
R5569 GND.n6117 GND.n1443 585
R5570 GND.n6124 GND.n6114 585
R5571 GND.n6114 GND.n1449 585
R5572 GND.n6125 GND.n6113 585
R5573 GND.n6113 GND.n1453 585
R5574 GND.n6126 GND.n6112 585
R5575 GND.n6112 GND.n1460 585
R5576 GND.n1492 GND.n1467 585
R5577 GND.n6169 GND.n1467 585
R5578 GND.n6131 GND.n6130 585
R5579 GND.n6132 GND.n6131 585
R5580 GND.n1491 GND.n1476 585
R5581 GND.n6151 GND.n1476 585
R5582 GND.n6108 GND.n1484 585
R5583 GND.n6141 GND.n1484 585
R5584 GND.n6107 GND.n6106 585
R5585 GND.n6106 GND.n6105 585
R5586 GND.n1495 GND.n1494 585
R5587 GND.n6028 GND.n1495 585
R5588 GND.n5962 GND.n1503 585
R5589 GND.n6097 GND.n1503 585
R5590 GND.n5963 GND.n5959 585
R5591 GND.n5959 GND.n1510 585
R5592 GND.n5964 GND.n5958 585
R5593 GND.n5958 GND.n1520 585
R5594 GND.n5956 GND.n1526 585
R5595 GND.n6067 GND.n1526 585
R5596 GND.n5968 GND.n5955 585
R5597 GND.n5955 GND.n1524 585
R5598 GND.n5969 GND.n1536 585
R5599 GND.n6058 GND.n1536 585
R5600 GND.n5970 GND.n1543 585
R5601 GND.n6051 GND.n1543 585
R5602 GND.n1571 GND.n1547 585
R5603 GND.n6014 GND.n1547 585
R5604 GND.n5975 GND.n5974 585
R5605 GND.n5976 GND.n5975 585
R5606 GND.n1570 GND.n1554 585
R5607 GND.n6006 GND.n1554 585
R5608 GND.n5951 GND.n5950 585
R5609 GND.n5950 GND.n1564 585
R5610 GND.n5949 GND.n1573 585
R5611 GND.n5949 GND.n1562 585
R5612 GND.n5948 GND.n1575 585
R5613 GND.n5948 GND.n5947 585
R5614 GND.n5870 GND.n1574 585
R5615 GND.n5917 GND.n1574 585
R5616 GND.n5871 GND.n1586 585
R5617 GND.n5938 GND.n1586 585
R5618 GND.n5872 GND.n1595 585
R5619 GND.n5925 GND.n1595 585
R5620 GND.n1644 GND.n1620 585
R5621 GND.n5905 GND.n1620 585
R5622 GND.n5877 GND.n5876 585
R5623 GND.n5878 GND.n5877 585
R5624 GND.n1643 GND.n1628 585
R5625 GND.n5897 GND.n1628 585
R5626 GND.n5864 GND.n1637 585
R5627 GND.n5886 GND.n1637 585
R5628 GND.n5863 GND.n5862 585
R5629 GND.n5862 GND.n5861 585
R5630 GND.n1647 GND.n1646 585
R5631 GND.n1662 GND.n1647 585
R5632 GND.n1671 GND.n1657 585
R5633 GND.n5853 GND.n1657 585
R5634 GND.n5837 GND.n5836 585
R5635 GND.n5838 GND.n5837 585
R5636 GND.n1670 GND.n1669 585
R5637 GND.n5809 GND.n1669 585
R5638 GND.n5830 GND.n5829 585
R5639 GND.n5829 GND.n5828 585
R5640 GND.n1674 GND.n1673 585
R5641 GND.n5782 GND.n1674 585
R5642 GND.n5727 GND.n1684 585
R5643 GND.n5819 GND.n1684 585
R5644 GND.n1722 GND.n1682 585
R5645 GND.n5760 GND.n5759 585
R5646 GND.n1723 GND.n1721 585
R5647 GND.n5762 GND.n1721 585
R5648 GND.n5755 GND.n5698 585
R5649 GND.n5754 GND.n5699 585
R5650 GND.n5701 GND.n5700 585
R5651 GND.n5750 GND.n5703 585
R5652 GND.n5749 GND.n5704 585
R5653 GND.n5748 GND.n5705 585
R5654 GND.n5707 GND.n5706 585
R5655 GND.n5744 GND.n5709 585
R5656 GND.n5743 GND.n5710 585
R5657 GND.n5742 GND.n5711 585
R5658 GND.n5713 GND.n5712 585
R5659 GND.n5738 GND.n5715 585
R5660 GND.n5737 GND.n5716 585
R5661 GND.n5736 GND.n5717 585
R5662 GND.n5733 GND.n5722 585
R5663 GND.n5732 GND.n5723 585
R5664 GND.n5731 GND.n5724 585
R5665 GND.n5726 GND.n5725 585
R5666 GND.n1337 GND.n1335 585
R5667 GND.n1335 GND.n1321 585
R5668 GND.n6315 GND.n6314 585
R5669 GND.n6316 GND.n6315 585
R5670 GND.n1336 GND.n1334 585
R5671 GND.n6213 GND.n1334 585
R5672 GND.n6267 GND.n6266 585
R5673 GND.n6268 GND.n6267 585
R5674 GND.n1423 GND.n1422 585
R5675 GND.n1436 GND.n1422 585
R5676 GND.n6262 GND.n6261 585
R5677 GND.n6261 GND.n6260 585
R5678 GND.n1426 GND.n1425 585
R5679 GND.n1445 GND.n1426 585
R5680 GND.n6161 GND.n6159 585
R5681 GND.n6159 GND.n1443 585
R5682 GND.n6162 GND.n6158 585
R5683 GND.n6158 GND.n1449 585
R5684 GND.n6163 GND.n6157 585
R5685 GND.n6157 GND.n1453 585
R5686 GND.n1471 GND.n1469 585
R5687 GND.n1469 GND.n1460 585
R5688 GND.n6168 GND.n6167 585
R5689 GND.n6169 GND.n6168 585
R5690 GND.n1470 GND.n1468 585
R5691 GND.n6132 GND.n1468 585
R5692 GND.n6153 GND.n6152 585
R5693 GND.n6152 GND.n6151 585
R5694 GND.n1474 GND.n1473 585
R5695 GND.n6141 GND.n1474 585
R5696 GND.n6104 GND.n6103 585
R5697 GND.n6105 GND.n6104 585
R5698 GND.n1498 GND.n1497 585
R5699 GND.n6028 GND.n1497 585
R5700 GND.n6099 GND.n6098 585
R5701 GND.n6098 GND.n6097 585
R5702 GND.n1501 GND.n1500 585
R5703 GND.n1510 GND.n1501 585
R5704 GND.n1530 GND.n1528 585
R5705 GND.n1528 GND.n1520 585
R5706 GND.n6066 GND.n6065 585
R5707 GND.n6067 GND.n6066 585
R5708 GND.n1529 GND.n1527 585
R5709 GND.n1527 GND.n1524 585
R5710 GND.n6060 GND.n6059 585
R5711 GND.n6059 GND.n6058 585
R5712 GND.n1533 GND.n1532 585
R5713 GND.n6051 GND.n1533 585
R5714 GND.n6013 GND.n6012 585
R5715 GND.n6014 GND.n6013 585
R5716 GND.n1549 GND.n1548 585
R5717 GND.n5976 GND.n1548 585
R5718 GND.n6008 GND.n6007 585
R5719 GND.n6007 GND.n6006 585
R5720 GND.n1552 GND.n1551 585
R5721 GND.n1564 GND.n1552 585
R5722 GND.n1581 GND.n1579 585
R5723 GND.n1579 GND.n1562 585
R5724 GND.n5946 GND.n5945 585
R5725 GND.n5947 GND.n5946 585
R5726 GND.n1580 GND.n1578 585
R5727 GND.n5917 GND.n1578 585
R5728 GND.n5940 GND.n5939 585
R5729 GND.n5939 GND.n5938 585
R5730 GND.n1584 GND.n1583 585
R5731 GND.n5925 GND.n1584 585
R5732 GND.n5904 GND.n5903 585
R5733 GND.n5905 GND.n5904 585
R5734 GND.n1623 GND.n1622 585
R5735 GND.n5878 GND.n1622 585
R5736 GND.n5899 GND.n5898 585
R5737 GND.n5898 GND.n5897 585
R5738 GND.n1626 GND.n1625 585
R5739 GND.n5886 GND.n1626 585
R5740 GND.n5860 GND.n5859 585
R5741 GND.n5861 GND.n5860 585
R5742 GND.n1651 GND.n1650 585
R5743 GND.n1662 GND.n1650 585
R5744 GND.n5855 GND.n5854 585
R5745 GND.n5854 GND.n5853 585
R5746 GND.n1654 GND.n1653 585
R5747 GND.n5838 GND.n1654 585
R5748 GND.n1680 GND.n1678 585
R5749 GND.n5809 GND.n1678 585
R5750 GND.n5827 GND.n5826 585
R5751 GND.n5828 GND.n5827 585
R5752 GND.n1679 GND.n1677 585
R5753 GND.n5782 GND.n1677 585
R5754 GND.n5821 GND.n5820 585
R5755 GND.n5820 GND.n5819 585
R5756 GND.n6663 GND.n1173 550.159
R5757 GND.n6577 GND.n6575 550.159
R5758 GND.n2184 GND.n2183 550.159
R5759 GND.n5674 GND.n1810 550.159
R5760 GND.n85 GND.n75 289.615
R5761 GND.n106 GND.n96 289.615
R5762 GND.n47 GND.n37 289.615
R5763 GND.n68 GND.n58 289.615
R5764 GND.n10 GND.n0 289.615
R5765 GND.n31 GND.n21 289.615
R5766 GND.n220 GND.n210 289.615
R5767 GND.n199 GND.n189 289.615
R5768 GND.n182 GND.n172 289.615
R5769 GND.n161 GND.n151 289.615
R5770 GND.n145 GND.n135 289.615
R5771 GND.n124 GND.n114 289.615
R5772 GND.n4858 GND.n3527 280.613
R5773 GND.n4858 GND.n4857 280.613
R5774 GND.n4857 GND.n4856 280.613
R5775 GND.n4856 GND.n3528 280.613
R5776 GND.n4850 GND.n3528 280.613
R5777 GND.n4850 GND.n4849 280.613
R5778 GND.n4849 GND.n4848 280.613
R5779 GND.n4848 GND.n3536 280.613
R5780 GND.n4842 GND.n3536 280.613
R5781 GND.n4842 GND.n4841 280.613
R5782 GND.n4841 GND.n4840 280.613
R5783 GND.n4840 GND.n3544 280.613
R5784 GND.n4834 GND.n3544 280.613
R5785 GND.n4834 GND.n4833 280.613
R5786 GND.n4833 GND.n4832 280.613
R5787 GND.n4832 GND.n3552 280.613
R5788 GND.n4826 GND.n3552 280.613
R5789 GND.n4826 GND.n4825 280.613
R5790 GND.n4825 GND.n4824 280.613
R5791 GND.n4824 GND.n3560 280.613
R5792 GND.n4818 GND.n3560 280.613
R5793 GND.n4818 GND.n4817 280.613
R5794 GND.n4817 GND.n4816 280.613
R5795 GND.n4816 GND.n3568 280.613
R5796 GND.n4810 GND.n3568 280.613
R5797 GND.n4810 GND.n4809 280.613
R5798 GND.n4809 GND.n4808 280.613
R5799 GND.n4808 GND.n3576 280.613
R5800 GND.n4802 GND.n3576 280.613
R5801 GND.n4802 GND.n4801 280.613
R5802 GND.n4801 GND.n4800 280.613
R5803 GND.n4800 GND.n3584 280.613
R5804 GND.n4794 GND.n3584 280.613
R5805 GND.n4794 GND.n4793 280.613
R5806 GND.n4793 GND.n4792 280.613
R5807 GND.n4792 GND.n3592 280.613
R5808 GND.n4786 GND.n3592 280.613
R5809 GND.n4786 GND.n4785 280.613
R5810 GND.n4785 GND.n4784 280.613
R5811 GND.n4784 GND.n3600 280.613
R5812 GND.n4778 GND.n3600 280.613
R5813 GND.n4778 GND.n4777 280.613
R5814 GND.n4777 GND.n4776 280.613
R5815 GND.n4776 GND.n3608 280.613
R5816 GND.n4770 GND.n3608 280.613
R5817 GND.n4770 GND.n4769 280.613
R5818 GND.n4769 GND.n4768 280.613
R5819 GND.n4768 GND.n3616 280.613
R5820 GND.n4762 GND.n3616 280.613
R5821 GND.n4762 GND.n4761 280.613
R5822 GND.n4761 GND.n4760 280.613
R5823 GND.n4760 GND.n3624 280.613
R5824 GND.n4754 GND.n3624 280.613
R5825 GND.n4754 GND.n4753 280.613
R5826 GND.n4753 GND.n4752 280.613
R5827 GND.n4752 GND.n3632 280.613
R5828 GND.n4746 GND.n3632 280.613
R5829 GND.n4746 GND.n4745 280.613
R5830 GND.n4745 GND.n4744 280.613
R5831 GND.n4744 GND.n3640 280.613
R5832 GND.n4738 GND.n3640 280.613
R5833 GND.n4738 GND.n4737 280.613
R5834 GND.n4737 GND.n4736 280.613
R5835 GND.n4736 GND.n3648 280.613
R5836 GND.n4730 GND.n3648 280.613
R5837 GND.n4730 GND.n4729 280.613
R5838 GND.n4729 GND.n4728 280.613
R5839 GND.n4728 GND.n3656 280.613
R5840 GND.n4722 GND.n3656 280.613
R5841 GND.n4722 GND.n4721 280.613
R5842 GND.n4721 GND.n4720 280.613
R5843 GND.n4720 GND.n3664 280.613
R5844 GND.n4714 GND.n3664 280.613
R5845 GND.n4714 GND.n4713 280.613
R5846 GND.n4713 GND.n4712 280.613
R5847 GND.n4712 GND.n3672 280.613
R5848 GND.n4706 GND.n3672 280.613
R5849 GND.n4706 GND.n4705 280.613
R5850 GND.n4705 GND.n4704 280.613
R5851 GND.n4704 GND.n3680 280.613
R5852 GND.n4698 GND.n3680 280.613
R5853 GND.n4698 GND.n4697 280.613
R5854 GND.n4697 GND.n4696 280.613
R5855 GND.n4696 GND.n3688 280.613
R5856 GND.n4690 GND.n3688 280.613
R5857 GND.n4690 GND.n4689 280.613
R5858 GND.n4689 GND.n4688 280.613
R5859 GND.n4688 GND.n3696 280.613
R5860 GND.n4682 GND.n3696 280.613
R5861 GND.n4682 GND.n4681 280.613
R5862 GND.n4681 GND.n4680 280.613
R5863 GND.n4680 GND.n3704 280.613
R5864 GND.n4674 GND.n3704 280.613
R5865 GND.n4674 GND.n4673 280.613
R5866 GND.n4673 GND.n4672 280.613
R5867 GND.n4672 GND.n3712 280.613
R5868 GND.n4666 GND.n3712 280.613
R5869 GND.n4666 GND.n4665 280.613
R5870 GND.n4665 GND.n4664 280.613
R5871 GND.n4664 GND.n3720 280.613
R5872 GND.n4658 GND.n3720 280.613
R5873 GND.n4658 GND.n4657 280.613
R5874 GND.n4657 GND.n4656 280.613
R5875 GND.n4656 GND.n3728 280.613
R5876 GND.n4650 GND.n3728 280.613
R5877 GND.n4650 GND.n4649 280.613
R5878 GND.n4649 GND.n4648 280.613
R5879 GND.n4648 GND.n3736 280.613
R5880 GND.n4642 GND.n3736 280.613
R5881 GND.n4642 GND.n4641 280.613
R5882 GND.n4641 GND.n4640 280.613
R5883 GND.n4640 GND.n3744 280.613
R5884 GND.n4634 GND.n3744 280.613
R5885 GND.n4634 GND.n4633 280.613
R5886 GND.n4633 GND.n4632 280.613
R5887 GND.n4632 GND.n3752 280.613
R5888 GND.n4626 GND.n3752 280.613
R5889 GND.n4626 GND.n4625 280.613
R5890 GND.n4625 GND.n4624 280.613
R5891 GND.n4624 GND.n3760 280.613
R5892 GND.n4618 GND.n3760 280.613
R5893 GND.n4618 GND.n4617 280.613
R5894 GND.n4617 GND.n4616 280.613
R5895 GND.n4616 GND.n3768 280.613
R5896 GND.n4610 GND.n3768 280.613
R5897 GND.n4610 GND.n4609 280.613
R5898 GND.n4609 GND.n4608 280.613
R5899 GND.n4608 GND.n3776 280.613
R5900 GND.n4602 GND.n3776 280.613
R5901 GND.n4602 GND.n4601 280.613
R5902 GND.n4601 GND.n4600 280.613
R5903 GND.n4600 GND.n3784 280.613
R5904 GND.n4594 GND.n3784 280.613
R5905 GND.n4594 GND.n4593 280.613
R5906 GND.n4593 GND.n4592 280.613
R5907 GND.n4592 GND.n3792 280.613
R5908 GND.n4586 GND.n3792 280.613
R5909 GND.n4586 GND.n4585 280.613
R5910 GND.n4585 GND.n4584 280.613
R5911 GND.n4584 GND.n3800 280.613
R5912 GND.n4578 GND.n3800 280.613
R5913 GND.n4578 GND.n4577 280.613
R5914 GND.n4577 GND.n4576 280.613
R5915 GND.n4576 GND.n3808 280.613
R5916 GND.n4570 GND.n3808 280.613
R5917 GND.n4570 GND.n4569 280.613
R5918 GND.n4569 GND.n4568 280.613
R5919 GND.n4568 GND.n3816 280.613
R5920 GND.n4562 GND.n3816 280.613
R5921 GND.n4562 GND.n4561 280.613
R5922 GND.n4561 GND.n4560 280.613
R5923 GND.n4560 GND.n3824 280.613
R5924 GND.n4554 GND.n3824 280.613
R5925 GND.n4554 GND.n4553 280.613
R5926 GND.n4553 GND.n4552 280.613
R5927 GND.n4552 GND.n3832 280.613
R5928 GND.n4546 GND.n3832 280.613
R5929 GND.n4546 GND.n4545 280.613
R5930 GND.n4545 GND.n4544 280.613
R5931 GND.n4544 GND.n3840 280.613
R5932 GND.n4538 GND.n3840 280.613
R5933 GND.n4538 GND.n4537 280.613
R5934 GND.n4537 GND.n4536 280.613
R5935 GND.n4536 GND.n3848 280.613
R5936 GND.n4530 GND.n3848 280.613
R5937 GND.n4530 GND.n4529 280.613
R5938 GND.n4529 GND.n4528 280.613
R5939 GND.n4528 GND.n3856 280.613
R5940 GND.n4522 GND.n3856 280.613
R5941 GND.n4522 GND.n4521 280.613
R5942 GND.n4521 GND.n4520 280.613
R5943 GND.n4520 GND.n3864 280.613
R5944 GND.n4514 GND.n3864 280.613
R5945 GND.n4514 GND.n4513 280.613
R5946 GND.n4513 GND.n4512 280.613
R5947 GND.n4512 GND.n3872 280.613
R5948 GND.n4506 GND.n3872 280.613
R5949 GND.n4506 GND.n4505 280.613
R5950 GND.n4505 GND.n4504 280.613
R5951 GND.n4504 GND.n3880 280.613
R5952 GND.n4498 GND.n3880 280.613
R5953 GND.n4498 GND.n4497 280.613
R5954 GND.n4497 GND.n4496 280.613
R5955 GND.n4496 GND.n3888 280.613
R5956 GND.n4490 GND.n3888 280.613
R5957 GND.n4490 GND.n4489 280.613
R5958 GND.n4489 GND.n4488 280.613
R5959 GND.n4488 GND.n3896 280.613
R5960 GND.n4482 GND.n3896 280.613
R5961 GND.n4482 GND.n4481 280.613
R5962 GND.n4481 GND.n4480 280.613
R5963 GND.n4480 GND.n3904 280.613
R5964 GND.n4474 GND.n3904 280.613
R5965 GND.n4474 GND.n4473 280.613
R5966 GND.n4473 GND.n4472 280.613
R5967 GND.n4472 GND.n3912 280.613
R5968 GND.n4466 GND.n3912 280.613
R5969 GND.n4466 GND.n4465 280.613
R5970 GND.n4465 GND.n4464 280.613
R5971 GND.n4464 GND.n3920 280.613
R5972 GND.n4458 GND.n3920 280.613
R5973 GND.n4458 GND.n4457 280.613
R5974 GND.n4457 GND.n4456 280.613
R5975 GND.n4456 GND.n3928 280.613
R5976 GND.n4450 GND.n3928 280.613
R5977 GND.n4450 GND.n4449 280.613
R5978 GND.n4449 GND.n4448 280.613
R5979 GND.n4448 GND.n3936 280.613
R5980 GND.n4442 GND.n3936 280.613
R5981 GND.n4442 GND.n4441 280.613
R5982 GND.n4441 GND.n4440 280.613
R5983 GND.n4440 GND.n3944 280.613
R5984 GND.n4434 GND.n3944 280.613
R5985 GND.n4434 GND.n4433 280.613
R5986 GND.n4433 GND.n4432 280.613
R5987 GND.n4432 GND.n3952 280.613
R5988 GND.n4426 GND.n3952 280.613
R5989 GND.n4426 GND.n4425 280.613
R5990 GND.n4425 GND.n4424 280.613
R5991 GND.n4424 GND.n3960 280.613
R5992 GND.n4418 GND.n3960 280.613
R5993 GND.n4418 GND.n4417 280.613
R5994 GND.n4417 GND.n4416 280.613
R5995 GND.n4416 GND.n3968 280.613
R5996 GND.n4410 GND.n3968 280.613
R5997 GND.n4410 GND.n4409 280.613
R5998 GND.n4409 GND.n4408 280.613
R5999 GND.n4408 GND.n3976 280.613
R6000 GND.n4402 GND.n3976 280.613
R6001 GND.n4402 GND.n4401 280.613
R6002 GND.n4401 GND.n4400 280.613
R6003 GND.n4400 GND.n3984 280.613
R6004 GND.n4394 GND.n3984 280.613
R6005 GND.n4394 GND.n4393 280.613
R6006 GND.n4393 GND.n4392 280.613
R6007 GND.n4392 GND.n3992 280.613
R6008 GND.n4386 GND.n3992 280.613
R6009 GND.n4386 GND.n4385 280.613
R6010 GND.n4385 GND.n4384 280.613
R6011 GND.n4384 GND.n4000 280.613
R6012 GND.n4378 GND.n4000 280.613
R6013 GND.n4378 GND.n4377 280.613
R6014 GND.n4377 GND.n4376 280.613
R6015 GND.n4376 GND.n4008 280.613
R6016 GND.n4370 GND.n4008 280.613
R6017 GND.n4370 GND.n4369 280.613
R6018 GND.n4369 GND.n4368 280.613
R6019 GND.n4368 GND.n4016 280.613
R6020 GND.n4362 GND.n4016 280.613
R6021 GND.n4362 GND.n4361 280.613
R6022 GND.n4361 GND.n4360 280.613
R6023 GND.n4360 GND.n4024 280.613
R6024 GND.n4354 GND.n4024 280.613
R6025 GND.n4354 GND.n4353 280.613
R6026 GND.n4353 GND.n4352 280.613
R6027 GND.n4352 GND.n4032 280.613
R6028 GND.n4346 GND.n4032 280.613
R6029 GND.n4346 GND.n4345 280.613
R6030 GND.n4345 GND.n4344 280.613
R6031 GND.n4344 GND.n4040 280.613
R6032 GND.n4338 GND.n4040 280.613
R6033 GND.n4338 GND.n4337 280.613
R6034 GND.n4337 GND.n4336 280.613
R6035 GND.n4336 GND.n4048 280.613
R6036 GND.n4330 GND.n4048 280.613
R6037 GND.n4330 GND.n4329 280.613
R6038 GND.n4329 GND.n4328 280.613
R6039 GND.n4328 GND.n4056 280.613
R6040 GND.n4322 GND.n4056 280.613
R6041 GND.n4322 GND.n4321 280.613
R6042 GND.n4321 GND.n4320 280.613
R6043 GND.n4320 GND.n4064 280.613
R6044 GND.n4314 GND.n4064 280.613
R6045 GND.n4314 GND.n4313 280.613
R6046 GND.n4313 GND.n4312 280.613
R6047 GND.n4312 GND.n4072 280.613
R6048 GND.n4306 GND.n4072 280.613
R6049 GND.n5718 GND.t37 257.43
R6050 GND.n1407 GND.t78 257.43
R6051 GND.n5676 GND.n5675 256.663
R6052 GND.n5676 GND.n1786 256.663
R6053 GND.n5676 GND.n1787 256.663
R6054 GND.n5676 GND.n1788 256.663
R6055 GND.n5676 GND.n1789 256.663
R6056 GND.n5676 GND.n1790 256.663
R6057 GND.n5676 GND.n1791 256.663
R6058 GND.n5676 GND.n1792 256.663
R6059 GND.n5676 GND.n1793 256.663
R6060 GND.n5676 GND.n1794 256.663
R6061 GND.n5676 GND.n1795 256.663
R6062 GND.n5632 GND.n5631 256.663
R6063 GND.n5676 GND.n1796 256.663
R6064 GND.n5676 GND.n1797 256.663
R6065 GND.n5676 GND.n1798 256.663
R6066 GND.n5676 GND.n1799 256.663
R6067 GND.n5676 GND.n1800 256.663
R6068 GND.n5676 GND.n1801 256.663
R6069 GND.n5676 GND.n1802 256.663
R6070 GND.n5676 GND.n1803 256.663
R6071 GND.n5676 GND.n1804 256.663
R6072 GND.n5676 GND.n1805 256.663
R6073 GND.n5676 GND.n1806 256.663
R6074 GND.n6664 GND.n1152 256.663
R6075 GND.n6664 GND.n1153 256.663
R6076 GND.n6664 GND.n1154 256.663
R6077 GND.n6664 GND.n1155 256.663
R6078 GND.n6664 GND.n1156 256.663
R6079 GND.n6664 GND.n1157 256.663
R6080 GND.n6664 GND.n1158 256.663
R6081 GND.n6664 GND.n1159 256.663
R6082 GND.n6664 GND.n1160 256.663
R6083 GND.n6664 GND.n1161 256.663
R6084 GND.n6664 GND.n1162 256.663
R6085 GND.n6667 GND.n1149 256.663
R6086 GND.n6665 GND.n6664 256.663
R6087 GND.n6664 GND.n1163 256.663
R6088 GND.n6664 GND.n1164 256.663
R6089 GND.n6664 GND.n1165 256.663
R6090 GND.n6664 GND.n1166 256.663
R6091 GND.n6664 GND.n1167 256.663
R6092 GND.n6664 GND.n1168 256.663
R6093 GND.n6664 GND.n1169 256.663
R6094 GND.n6664 GND.n1170 256.663
R6095 GND.n6664 GND.n1171 256.663
R6096 GND.n6664 GND.n1172 256.663
R6097 GND.n2227 GND.t28 247.573
R6098 GND.n5606 GND.t64 247.573
R6099 GND.n1756 GND.t10 247.573
R6100 GND.n6670 GND.t62 247.573
R6101 GND.n6682 GND.t53 247.573
R6102 GND.n561 GND.t31 247.573
R6103 GND.n542 GND.t67 247.573
R6104 GND.n580 GND.t21 247.573
R6105 GND.n1363 GND.t47 247.573
R6106 GND.n3066 GND.t36 247.573
R6107 GND.n3086 GND.t59 247.573
R6108 GND.n3118 GND.t74 247.573
R6109 GND.n3134 GND.n3050 242.672
R6110 GND.n3093 GND.n3050 242.672
R6111 GND.n3098 GND.n3050 242.672
R6112 GND.n3103 GND.n3050 242.672
R6113 GND.n3116 GND.n3050 242.672
R6114 GND.n3177 GND.n3050 242.672
R6115 GND.n3056 GND.n3050 242.672
R6116 GND.n3170 GND.n3050 242.672
R6117 GND.n3164 GND.n3050 242.672
R6118 GND.n3162 GND.n3050 242.672
R6119 GND.n3156 GND.n3050 242.672
R6120 GND.n3154 GND.n3050 242.672
R6121 GND.n3148 GND.n3050 242.672
R6122 GND.n3146 GND.n3050 242.672
R6123 GND.n3084 GND.n3050 242.672
R6124 GND.n5025 GND.n5024 242.672
R6125 GND.n5025 GND.n2791 242.672
R6126 GND.n5025 GND.n2792 242.672
R6127 GND.n5025 GND.n2793 242.672
R6128 GND.n5025 GND.n2794 242.672
R6129 GND.n5025 GND.n2795 242.672
R6130 GND.n5025 GND.n2796 242.672
R6131 GND.n5025 GND.n2797 242.672
R6132 GND.n5025 GND.n2798 242.672
R6133 GND.n5025 GND.n2799 242.672
R6134 GND.n5025 GND.n2800 242.672
R6135 GND.n5025 GND.n2801 242.672
R6136 GND.n5025 GND.n2802 242.672
R6137 GND.n5025 GND.n2803 242.672
R6138 GND.n5025 GND.n2804 242.672
R6139 GND.n5025 GND.n2805 242.672
R6140 GND.n5025 GND.n2806 242.672
R6141 GND.n5025 GND.n2807 242.672
R6142 GND.n5025 GND.n2808 242.672
R6143 GND.n5025 GND.n2809 242.672
R6144 GND.n5025 GND.n2810 242.672
R6145 GND.n5025 GND.n2811 242.672
R6146 GND.n5025 GND.n2812 242.672
R6147 GND.n5025 GND.n2813 242.672
R6148 GND.n5025 GND.n2814 242.672
R6149 GND.n5025 GND.n2815 242.672
R6150 GND.n5025 GND.n2816 242.672
R6151 GND.n5026 GND.n5025 242.672
R6152 GND.n1777 GND.n1751 242.672
R6153 GND.n1777 GND.n1752 242.672
R6154 GND.n1777 GND.n1753 242.672
R6155 GND.n1777 GND.n1754 242.672
R6156 GND.n1777 GND.n1755 242.672
R6157 GND.n6725 GND.n955 242.672
R6158 GND.n6725 GND.n954 242.672
R6159 GND.n6725 GND.n953 242.672
R6160 GND.n6725 GND.n952 242.672
R6161 GND.n6725 GND.n951 242.672
R6162 GND.n7328 GND.n528 242.672
R6163 GND.n583 GND.n528 242.672
R6164 GND.n7335 GND.n528 242.672
R6165 GND.n574 GND.n528 242.672
R6166 GND.n7342 GND.n528 242.672
R6167 GND.n5610 GND.n1777 242.672
R6168 GND.n5608 GND.n1777 242.672
R6169 GND.n5602 GND.n1777 242.672
R6170 GND.n5599 GND.n1777 242.672
R6171 GND.n5594 GND.n1777 242.672
R6172 GND.n5591 GND.n1777 242.672
R6173 GND.n5630 GND.n5586 242.672
R6174 GND.n5585 GND.n1777 242.672
R6175 GND.n2230 GND.n1777 242.672
R6176 GND.n5574 GND.n1777 242.672
R6177 GND.n2234 GND.n1777 242.672
R6178 GND.n6725 GND.n6724 242.672
R6179 GND.n6725 GND.n941 242.672
R6180 GND.n6725 GND.n942 242.672
R6181 GND.n6725 GND.n943 242.672
R6182 GND.n6709 GND.n6668 242.672
R6183 GND.n6725 GND.n944 242.672
R6184 GND.n6725 GND.n945 242.672
R6185 GND.n6725 GND.n946 242.672
R6186 GND.n6725 GND.n947 242.672
R6187 GND.n6725 GND.n948 242.672
R6188 GND.n6725 GND.n949 242.672
R6189 GND.n7427 GND.n528 242.672
R6190 GND.n564 GND.n528 242.672
R6191 GND.n7434 GND.n528 242.672
R6192 GND.n555 GND.n528 242.672
R6193 GND.n7441 GND.n528 242.672
R6194 GND.n549 GND.n528 242.672
R6195 GND.n544 GND.n528 242.672
R6196 GND.n7452 GND.n528 242.672
R6197 GND.n536 GND.n528 242.672
R6198 GND.n7459 GND.n528 242.672
R6199 GND.n7462 GND.n528 242.672
R6200 GND.n1414 GND.n1317 242.672
R6201 GND.n1409 GND.n1317 242.672
R6202 GND.n1404 GND.n1317 242.672
R6203 GND.n1399 GND.n1317 242.672
R6204 GND.n1396 GND.n1317 242.672
R6205 GND.n1391 GND.n1317 242.672
R6206 GND.n1388 GND.n1317 242.672
R6207 GND.n1383 GND.n1317 242.672
R6208 GND.n1380 GND.n1317 242.672
R6209 GND.n1341 GND.n1317 242.672
R6210 GND.n5762 GND.n5761 242.672
R6211 GND.n5762 GND.n1712 242.672
R6212 GND.n5762 GND.n1713 242.672
R6213 GND.n5762 GND.n1714 242.672
R6214 GND.n5762 GND.n1715 242.672
R6215 GND.n5762 GND.n1716 242.672
R6216 GND.n5762 GND.n1717 242.672
R6217 GND.n5762 GND.n1718 242.672
R6218 GND.n5762 GND.n1719 242.672
R6219 GND.n5762 GND.n1720 242.672
R6220 GND.n1819 GND.t50 241.843
R6221 GND.n6532 GND.t55 241.843
R6222 GND.n1817 GND.t18 241.841
R6223 GND.n6622 GND.t25 241.841
R6224 GND.n7461 GND.n7460 240.244
R6225 GND.n7458 GND.n530 240.244
R6226 GND.n7454 GND.n7453 240.244
R6227 GND.n7451 GND.n537 240.244
R6228 GND.n548 GND.n545 240.244
R6229 GND.n7443 GND.n7442 240.244
R6230 GND.n7440 GND.n550 240.244
R6231 GND.n7436 GND.n7435 240.244
R6232 GND.n7433 GND.n556 240.244
R6233 GND.n7429 GND.n7428 240.244
R6234 GND.n6735 GND.n922 240.244
R6235 GND.n6751 GND.n922 240.244
R6236 GND.n6751 GND.n923 240.244
R6237 GND.n923 GND.n911 240.244
R6238 GND.n6746 GND.n911 240.244
R6239 GND.n6746 GND.n894 240.244
R6240 GND.n6862 GND.n894 240.244
R6241 GND.n6862 GND.n895 240.244
R6242 GND.n895 GND.n885 240.244
R6243 GND.n885 GND.n875 240.244
R6244 GND.n6882 GND.n875 240.244
R6245 GND.n6882 GND.n876 240.244
R6246 GND.n876 GND.n865 240.244
R6247 GND.n865 GND.n855 240.244
R6248 GND.n6902 GND.n855 240.244
R6249 GND.n6902 GND.n856 240.244
R6250 GND.n856 GND.n845 240.244
R6251 GND.n845 GND.n835 240.244
R6252 GND.n6922 GND.n835 240.244
R6253 GND.n6922 GND.n836 240.244
R6254 GND.n836 GND.n824 240.244
R6255 GND.n824 GND.n815 240.244
R6256 GND.n6942 GND.n815 240.244
R6257 GND.n6942 GND.n816 240.244
R6258 GND.n816 GND.n805 240.244
R6259 GND.n805 GND.n795 240.244
R6260 GND.n6962 GND.n795 240.244
R6261 GND.n6962 GND.n796 240.244
R6262 GND.n796 GND.n785 240.244
R6263 GND.n785 GND.n775 240.244
R6264 GND.n6982 GND.n775 240.244
R6265 GND.n6982 GND.n776 240.244
R6266 GND.n776 GND.n765 240.244
R6267 GND.n765 GND.n755 240.244
R6268 GND.n7002 GND.n755 240.244
R6269 GND.n7002 GND.n756 240.244
R6270 GND.n756 GND.n745 240.244
R6271 GND.n745 GND.n734 240.244
R6272 GND.n7026 GND.n734 240.244
R6273 GND.n7026 GND.n735 240.244
R6274 GND.n735 GND.n723 240.244
R6275 GND.n7021 GND.n723 240.244
R6276 GND.n7021 GND.n706 240.244
R6277 GND.n7070 GND.n706 240.244
R6278 GND.n7070 GND.n707 240.244
R6279 GND.n707 GND.n697 240.244
R6280 GND.n697 GND.n686 240.244
R6281 GND.n7098 GND.n686 240.244
R6282 GND.n7098 GND.n687 240.244
R6283 GND.n687 GND.n676 240.244
R6284 GND.n676 GND.n659 240.244
R6285 GND.n7134 GND.n659 240.244
R6286 GND.n7134 GND.n660 240.244
R6287 GND.n7130 GND.n660 240.244
R6288 GND.n7130 GND.n647 240.244
R6289 GND.n647 GND.n639 240.244
R6290 GND.n7159 GND.n639 240.244
R6291 GND.n7159 GND.n629 240.244
R6292 GND.n7169 GND.n629 240.244
R6293 GND.n7170 GND.n7169 240.244
R6294 GND.n7170 GND.n237 240.244
R6295 GND.n7173 GND.n237 240.244
R6296 GND.n7173 GND.n622 240.244
R6297 GND.n7204 GND.n622 240.244
R6298 GND.n7204 GND.n256 240.244
R6299 GND.n7631 GND.n256 240.244
R6300 GND.n7631 GND.n257 240.244
R6301 GND.n7627 GND.n257 240.244
R6302 GND.n7627 GND.n263 240.244
R6303 GND.n7619 GND.n263 240.244
R6304 GND.n7619 GND.n279 240.244
R6305 GND.n7615 GND.n279 240.244
R6306 GND.n7615 GND.n284 240.244
R6307 GND.n7607 GND.n284 240.244
R6308 GND.n7607 GND.n300 240.244
R6309 GND.n7603 GND.n300 240.244
R6310 GND.n7603 GND.n305 240.244
R6311 GND.n317 GND.n305 240.244
R6312 GND.n7348 GND.n317 240.244
R6313 GND.n7348 GND.n329 240.244
R6314 GND.n7352 GND.n329 240.244
R6315 GND.n7352 GND.n339 240.244
R6316 GND.n7355 GND.n339 240.244
R6317 GND.n7355 GND.n348 240.244
R6318 GND.n7359 GND.n348 240.244
R6319 GND.n7359 GND.n358 240.244
R6320 GND.n7362 GND.n358 240.244
R6321 GND.n7362 GND.n367 240.244
R6322 GND.n7366 GND.n367 240.244
R6323 GND.n7366 GND.n377 240.244
R6324 GND.n7369 GND.n377 240.244
R6325 GND.n7369 GND.n386 240.244
R6326 GND.n7373 GND.n386 240.244
R6327 GND.n7373 GND.n396 240.244
R6328 GND.n7376 GND.n396 240.244
R6329 GND.n7376 GND.n405 240.244
R6330 GND.n7380 GND.n405 240.244
R6331 GND.n7380 GND.n415 240.244
R6332 GND.n7383 GND.n415 240.244
R6333 GND.n7383 GND.n424 240.244
R6334 GND.n7387 GND.n424 240.244
R6335 GND.n7387 GND.n434 240.244
R6336 GND.n7390 GND.n434 240.244
R6337 GND.n7390 GND.n443 240.244
R6338 GND.n7394 GND.n443 240.244
R6339 GND.n7394 GND.n454 240.244
R6340 GND.n7397 GND.n454 240.244
R6341 GND.n7397 GND.n463 240.244
R6342 GND.n7401 GND.n463 240.244
R6343 GND.n7401 GND.n473 240.244
R6344 GND.n7404 GND.n473 240.244
R6345 GND.n7404 GND.n482 240.244
R6346 GND.n7408 GND.n482 240.244
R6347 GND.n7408 GND.n492 240.244
R6348 GND.n7411 GND.n492 240.244
R6349 GND.n7411 GND.n501 240.244
R6350 GND.n7415 GND.n501 240.244
R6351 GND.n7415 GND.n511 240.244
R6352 GND.n7418 GND.n511 240.244
R6353 GND.n7418 GND.n520 240.244
R6354 GND.n565 GND.n520 240.244
R6355 GND.n957 GND.n956 240.244
R6356 GND.n6718 GND.n956 240.244
R6357 GND.n6716 GND.n6715 240.244
R6358 GND.n6712 GND.n6711 240.244
R6359 GND.n6707 GND.n6706 240.244
R6360 GND.n6703 GND.n6702 240.244
R6361 GND.n6699 GND.n6698 240.244
R6362 GND.n6695 GND.n6694 240.244
R6363 GND.n6691 GND.n6690 240.244
R6364 GND.n6681 GND.n930 240.244
R6365 GND.n1135 GND.n932 240.244
R6366 GND.n1135 GND.n919 240.244
R6367 GND.n1132 GND.n919 240.244
R6368 GND.n1132 GND.n909 240.244
R6369 GND.n1129 GND.n909 240.244
R6370 GND.n1129 GND.n902 240.244
R6371 GND.n902 GND.n891 240.244
R6372 GND.n1125 GND.n891 240.244
R6373 GND.n1125 GND.n883 240.244
R6374 GND.n1122 GND.n883 240.244
R6375 GND.n1122 GND.n872 240.244
R6376 GND.n1119 GND.n872 240.244
R6377 GND.n1119 GND.n863 240.244
R6378 GND.n1116 GND.n863 240.244
R6379 GND.n1116 GND.n852 240.244
R6380 GND.n1113 GND.n852 240.244
R6381 GND.n1113 GND.n843 240.244
R6382 GND.n1110 GND.n843 240.244
R6383 GND.n1110 GND.n831 240.244
R6384 GND.n1107 GND.n831 240.244
R6385 GND.n1107 GND.n822 240.244
R6386 GND.n1104 GND.n822 240.244
R6387 GND.n1104 GND.n812 240.244
R6388 GND.n1101 GND.n812 240.244
R6389 GND.n1101 GND.n803 240.244
R6390 GND.n1098 GND.n803 240.244
R6391 GND.n1098 GND.n792 240.244
R6392 GND.n1095 GND.n792 240.244
R6393 GND.n1095 GND.n783 240.244
R6394 GND.n1092 GND.n783 240.244
R6395 GND.n1092 GND.n772 240.244
R6396 GND.n1089 GND.n772 240.244
R6397 GND.n1089 GND.n763 240.244
R6398 GND.n1086 GND.n763 240.244
R6399 GND.n1086 GND.n752 240.244
R6400 GND.n1083 GND.n752 240.244
R6401 GND.n1083 GND.n743 240.244
R6402 GND.n1080 GND.n743 240.244
R6403 GND.n1080 GND.n731 240.244
R6404 GND.n1077 GND.n731 240.244
R6405 GND.n1077 GND.n721 240.244
R6406 GND.n1074 GND.n721 240.244
R6407 GND.n1074 GND.n714 240.244
R6408 GND.n714 GND.n703 240.244
R6409 GND.n1070 GND.n703 240.244
R6410 GND.n1070 GND.n695 240.244
R6411 GND.n1067 GND.n695 240.244
R6412 GND.n1067 GND.n683 240.244
R6413 GND.n1064 GND.n683 240.244
R6414 GND.n1064 GND.n674 240.244
R6415 GND.n1061 GND.n674 240.244
R6416 GND.n1061 GND.n655 240.244
R6417 GND.n1058 GND.n655 240.244
R6418 GND.n1058 GND.n667 240.244
R6419 GND.n667 GND.n645 240.244
R6420 GND.n1013 GND.n645 240.244
R6421 GND.n1013 GND.n636 240.244
R6422 GND.n1051 GND.n636 240.244
R6423 GND.n1051 GND.n631 240.244
R6424 GND.n1047 GND.n631 240.244
R6425 GND.n1047 GND.n234 240.244
R6426 GND.n1043 GND.n234 240.244
R6427 GND.n1043 GND.n1042 240.244
R6428 GND.n1042 GND.n620 240.244
R6429 GND.n1037 GND.n620 240.244
R6430 GND.n1037 GND.n253 240.244
R6431 GND.n1034 GND.n253 240.244
R6432 GND.n1034 GND.n265 240.244
R6433 GND.n1031 GND.n265 240.244
R6434 GND.n1031 GND.n275 240.244
R6435 GND.n1028 GND.n275 240.244
R6436 GND.n1028 GND.n285 240.244
R6437 GND.n1025 GND.n285 240.244
R6438 GND.n1025 GND.n296 240.244
R6439 GND.n309 GND.n296 240.244
R6440 GND.n7601 GND.n309 240.244
R6441 GND.n7601 GND.n310 240.244
R6442 GND.n7597 GND.n310 240.244
R6443 GND.n7597 GND.n316 240.244
R6444 GND.n7589 GND.n316 240.244
R6445 GND.n7589 GND.n332 240.244
R6446 GND.n7585 GND.n332 240.244
R6447 GND.n7585 GND.n338 240.244
R6448 GND.n7577 GND.n338 240.244
R6449 GND.n7577 GND.n351 240.244
R6450 GND.n7573 GND.n351 240.244
R6451 GND.n7573 GND.n357 240.244
R6452 GND.n7565 GND.n357 240.244
R6453 GND.n7565 GND.n370 240.244
R6454 GND.n7561 GND.n370 240.244
R6455 GND.n7561 GND.n376 240.244
R6456 GND.n7553 GND.n376 240.244
R6457 GND.n7553 GND.n389 240.244
R6458 GND.n7549 GND.n389 240.244
R6459 GND.n7549 GND.n395 240.244
R6460 GND.n7541 GND.n395 240.244
R6461 GND.n7541 GND.n408 240.244
R6462 GND.n7537 GND.n408 240.244
R6463 GND.n7537 GND.n414 240.244
R6464 GND.n7529 GND.n414 240.244
R6465 GND.n7529 GND.n426 240.244
R6466 GND.n7525 GND.n426 240.244
R6467 GND.n7525 GND.n432 240.244
R6468 GND.n7517 GND.n432 240.244
R6469 GND.n7517 GND.n446 240.244
R6470 GND.n7513 GND.n446 240.244
R6471 GND.n7513 GND.n452 240.244
R6472 GND.n7505 GND.n452 240.244
R6473 GND.n7505 GND.n466 240.244
R6474 GND.n7501 GND.n466 240.244
R6475 GND.n7501 GND.n472 240.244
R6476 GND.n7493 GND.n472 240.244
R6477 GND.n7493 GND.n485 240.244
R6478 GND.n7489 GND.n485 240.244
R6479 GND.n7489 GND.n491 240.244
R6480 GND.n7481 GND.n491 240.244
R6481 GND.n7481 GND.n504 240.244
R6482 GND.n7477 GND.n504 240.244
R6483 GND.n7477 GND.n510 240.244
R6484 GND.n7469 GND.n510 240.244
R6485 GND.n7469 GND.n523 240.244
R6486 GND.n7344 GND.n7343 240.244
R6487 GND.n7341 GND.n569 240.244
R6488 GND.n7337 GND.n7336 240.244
R6489 GND.n7334 GND.n575 240.244
R6490 GND.n7330 GND.n7329 240.244
R6491 GND.n1372 GND.n934 240.244
R6492 GND.n1372 GND.n921 240.244
R6493 GND.n921 GND.n907 240.244
R6494 GND.n6763 GND.n907 240.244
R6495 GND.n6763 GND.n903 240.244
R6496 GND.n6851 GND.n903 240.244
R6497 GND.n6851 GND.n893 240.244
R6498 GND.n6847 GND.n893 240.244
R6499 GND.n6847 GND.n884 240.244
R6500 GND.n6844 GND.n884 240.244
R6501 GND.n6844 GND.n874 240.244
R6502 GND.n6841 GND.n874 240.244
R6503 GND.n6841 GND.n864 240.244
R6504 GND.n6838 GND.n864 240.244
R6505 GND.n6838 GND.n854 240.244
R6506 GND.n6835 GND.n854 240.244
R6507 GND.n6835 GND.n844 240.244
R6508 GND.n6832 GND.n844 240.244
R6509 GND.n6832 GND.n834 240.244
R6510 GND.n6829 GND.n834 240.244
R6511 GND.n6829 GND.n823 240.244
R6512 GND.n6826 GND.n823 240.244
R6513 GND.n6826 GND.n814 240.244
R6514 GND.n6823 GND.n814 240.244
R6515 GND.n6823 GND.n804 240.244
R6516 GND.n6820 GND.n804 240.244
R6517 GND.n6820 GND.n794 240.244
R6518 GND.n6817 GND.n794 240.244
R6519 GND.n6817 GND.n784 240.244
R6520 GND.n6814 GND.n784 240.244
R6521 GND.n6814 GND.n774 240.244
R6522 GND.n6811 GND.n774 240.244
R6523 GND.n6811 GND.n764 240.244
R6524 GND.n6808 GND.n764 240.244
R6525 GND.n6808 GND.n754 240.244
R6526 GND.n6805 GND.n754 240.244
R6527 GND.n6805 GND.n744 240.244
R6528 GND.n6802 GND.n744 240.244
R6529 GND.n6802 GND.n733 240.244
R6530 GND.n733 GND.n719 240.244
R6531 GND.n7038 GND.n719 240.244
R6532 GND.n7038 GND.n715 240.244
R6533 GND.n7059 GND.n715 240.244
R6534 GND.n7059 GND.n705 240.244
R6535 GND.n7055 GND.n705 240.244
R6536 GND.n7055 GND.n696 240.244
R6537 GND.n7052 GND.n696 240.244
R6538 GND.n7052 GND.n685 240.244
R6539 GND.n685 GND.n672 240.244
R6540 GND.n7108 GND.n672 240.244
R6541 GND.n7109 GND.n7108 240.244
R6542 GND.n7109 GND.n658 240.244
R6543 GND.n668 GND.n658 240.244
R6544 GND.n7128 GND.n668 240.244
R6545 GND.n7128 GND.n646 240.244
R6546 GND.n7124 GND.n646 240.244
R6547 GND.n7124 GND.n638 240.244
R6548 GND.n7121 GND.n638 240.244
R6549 GND.n7121 GND.n633 240.244
R6550 GND.n633 GND.n231 240.244
R6551 GND.n7642 GND.n231 240.244
R6552 GND.n7642 GND.n232 240.244
R6553 GND.n618 GND.n232 240.244
R6554 GND.n7209 GND.n618 240.244
R6555 GND.n7210 GND.n7209 240.244
R6556 GND.n7210 GND.n255 240.244
R6557 GND.n7215 GND.n255 240.244
R6558 GND.n7215 GND.n268 240.244
R6559 GND.n7218 GND.n268 240.244
R6560 GND.n7218 GND.n278 240.244
R6561 GND.n7223 GND.n278 240.244
R6562 GND.n7223 GND.n288 240.244
R6563 GND.n7226 GND.n288 240.244
R6564 GND.n7226 GND.n299 240.244
R6565 GND.n7231 GND.n299 240.244
R6566 GND.n7231 GND.n306 240.244
R6567 GND.n7235 GND.n306 240.244
R6568 GND.n7235 GND.n318 240.244
R6569 GND.n7240 GND.n318 240.244
R6570 GND.n7240 GND.n330 240.244
R6571 GND.n7243 GND.n330 240.244
R6572 GND.n7243 GND.n340 240.244
R6573 GND.n7248 GND.n340 240.244
R6574 GND.n7248 GND.n349 240.244
R6575 GND.n7251 GND.n349 240.244
R6576 GND.n7251 GND.n359 240.244
R6577 GND.n7256 GND.n359 240.244
R6578 GND.n7256 GND.n368 240.244
R6579 GND.n7259 GND.n368 240.244
R6580 GND.n7259 GND.n378 240.244
R6581 GND.n7264 GND.n378 240.244
R6582 GND.n7264 GND.n387 240.244
R6583 GND.n7267 GND.n387 240.244
R6584 GND.n7267 GND.n397 240.244
R6585 GND.n7272 GND.n397 240.244
R6586 GND.n7272 GND.n406 240.244
R6587 GND.n7275 GND.n406 240.244
R6588 GND.n7275 GND.n416 240.244
R6589 GND.n7280 GND.n416 240.244
R6590 GND.n7280 GND.n425 240.244
R6591 GND.n7283 GND.n425 240.244
R6592 GND.n7283 GND.n435 240.244
R6593 GND.n7288 GND.n435 240.244
R6594 GND.n7288 GND.n444 240.244
R6595 GND.n7291 GND.n444 240.244
R6596 GND.n7291 GND.n455 240.244
R6597 GND.n7296 GND.n455 240.244
R6598 GND.n7296 GND.n464 240.244
R6599 GND.n7299 GND.n464 240.244
R6600 GND.n7299 GND.n474 240.244
R6601 GND.n7304 GND.n474 240.244
R6602 GND.n7304 GND.n483 240.244
R6603 GND.n7307 GND.n483 240.244
R6604 GND.n7307 GND.n493 240.244
R6605 GND.n7312 GND.n493 240.244
R6606 GND.n7312 GND.n502 240.244
R6607 GND.n7315 GND.n502 240.244
R6608 GND.n7315 GND.n512 240.244
R6609 GND.n7320 GND.n512 240.244
R6610 GND.n7320 GND.n521 240.244
R6611 GND.n584 GND.n521 240.244
R6612 GND.n1349 GND.n1348 240.244
R6613 GND.n1354 GND.n1353 240.244
R6614 GND.n1359 GND.n1358 240.244
R6615 GND.n1367 GND.n1366 240.244
R6616 GND.n1362 GND.n950 240.244
R6617 GND.n933 GND.n928 240.244
R6618 GND.n928 GND.n920 240.244
R6619 GND.n6741 GND.n920 240.244
R6620 GND.n6741 GND.n910 240.244
R6621 GND.n910 GND.n900 240.244
R6622 GND.n6853 GND.n900 240.244
R6623 GND.n6853 GND.n892 240.244
R6624 GND.n892 GND.n881 240.244
R6625 GND.n6872 GND.n881 240.244
R6626 GND.n6873 GND.n6872 240.244
R6627 GND.n6873 GND.n873 240.244
R6628 GND.n873 GND.n861 240.244
R6629 GND.n6892 GND.n861 240.244
R6630 GND.n6893 GND.n6892 240.244
R6631 GND.n6893 GND.n853 240.244
R6632 GND.n853 GND.n841 240.244
R6633 GND.n6912 GND.n841 240.244
R6634 GND.n6913 GND.n6912 240.244
R6635 GND.n6913 GND.n832 240.244
R6636 GND.n832 GND.n821 240.244
R6637 GND.n6932 GND.n821 240.244
R6638 GND.n6933 GND.n6932 240.244
R6639 GND.n6933 GND.n813 240.244
R6640 GND.n813 GND.n801 240.244
R6641 GND.n6952 GND.n801 240.244
R6642 GND.n6953 GND.n6952 240.244
R6643 GND.n6953 GND.n793 240.244
R6644 GND.n793 GND.n781 240.244
R6645 GND.n6972 GND.n781 240.244
R6646 GND.n6973 GND.n6972 240.244
R6647 GND.n6973 GND.n773 240.244
R6648 GND.n773 GND.n761 240.244
R6649 GND.n6992 GND.n761 240.244
R6650 GND.n6993 GND.n6992 240.244
R6651 GND.n6993 GND.n753 240.244
R6652 GND.n753 GND.n741 240.244
R6653 GND.n7012 GND.n741 240.244
R6654 GND.n7013 GND.n7012 240.244
R6655 GND.n7013 GND.n732 240.244
R6656 GND.n7016 GND.n732 240.244
R6657 GND.n7016 GND.n722 240.244
R6658 GND.n722 GND.n712 240.244
R6659 GND.n7061 GND.n712 240.244
R6660 GND.n7061 GND.n704 240.244
R6661 GND.n704 GND.n693 240.244
R6662 GND.n7080 GND.n693 240.244
R6663 GND.n7081 GND.n7080 240.244
R6664 GND.n7081 GND.n684 240.244
R6665 GND.n7084 GND.n684 240.244
R6666 GND.n7084 GND.n675 240.244
R6667 GND.n7091 GND.n675 240.244
R6668 GND.n7091 GND.n656 240.244
R6669 GND.n7088 GND.n656 240.244
R6670 GND.n7088 GND.n644 240.244
R6671 GND.n7146 GND.n644 240.244
R6672 GND.n7147 GND.n7146 240.244
R6673 GND.n7147 GND.n637 240.244
R6674 GND.n7150 GND.n637 240.244
R6675 GND.n7150 GND.n632 240.244
R6676 GND.n7152 GND.n632 240.244
R6677 GND.n7152 GND.n235 240.244
R6678 GND.n7177 GND.n235 240.244
R6679 GND.n7178 GND.n7177 240.244
R6680 GND.n7178 GND.n621 240.244
R6681 GND.n7199 GND.n621 240.244
R6682 GND.n7199 GND.n254 240.244
R6683 GND.n7196 GND.n254 240.244
R6684 GND.n7196 GND.n266 240.244
R6685 GND.n7193 GND.n266 240.244
R6686 GND.n7193 GND.n276 240.244
R6687 GND.n7190 GND.n276 240.244
R6688 GND.n7190 GND.n286 240.244
R6689 GND.n7187 GND.n286 240.244
R6690 GND.n7187 GND.n297 240.244
R6691 GND.n7184 GND.n297 240.244
R6692 GND.n7184 GND.n308 240.244
R6693 GND.n320 GND.n308 240.244
R6694 GND.n7595 GND.n320 240.244
R6695 GND.n7595 GND.n321 240.244
R6696 GND.n7591 GND.n321 240.244
R6697 GND.n7591 GND.n328 240.244
R6698 GND.n7583 GND.n328 240.244
R6699 GND.n7583 GND.n342 240.244
R6700 GND.n7579 GND.n342 240.244
R6701 GND.n7579 GND.n347 240.244
R6702 GND.n7571 GND.n347 240.244
R6703 GND.n7571 GND.n361 240.244
R6704 GND.n7567 GND.n361 240.244
R6705 GND.n7567 GND.n366 240.244
R6706 GND.n7559 GND.n366 240.244
R6707 GND.n7559 GND.n380 240.244
R6708 GND.n7555 GND.n380 240.244
R6709 GND.n7555 GND.n385 240.244
R6710 GND.n7547 GND.n385 240.244
R6711 GND.n7547 GND.n399 240.244
R6712 GND.n7543 GND.n399 240.244
R6713 GND.n7543 GND.n404 240.244
R6714 GND.n7535 GND.n404 240.244
R6715 GND.n7535 GND.n418 240.244
R6716 GND.n7531 GND.n418 240.244
R6717 GND.n7531 GND.n423 240.244
R6718 GND.n7523 GND.n423 240.244
R6719 GND.n7523 GND.n437 240.244
R6720 GND.n7519 GND.n437 240.244
R6721 GND.n7519 GND.n442 240.244
R6722 GND.n7511 GND.n442 240.244
R6723 GND.n7511 GND.n457 240.244
R6724 GND.n7507 GND.n457 240.244
R6725 GND.n7507 GND.n462 240.244
R6726 GND.n7499 GND.n462 240.244
R6727 GND.n7499 GND.n476 240.244
R6728 GND.n7495 GND.n476 240.244
R6729 GND.n7495 GND.n481 240.244
R6730 GND.n7487 GND.n481 240.244
R6731 GND.n7487 GND.n494 240.244
R6732 GND.n7483 GND.n494 240.244
R6733 GND.n7483 GND.n499 240.244
R6734 GND.n7475 GND.n499 240.244
R6735 GND.n7475 GND.n514 240.244
R6736 GND.n7471 GND.n514 240.244
R6737 GND.n7471 GND.n519 240.244
R6738 GND.n4859 GND.n3523 240.244
R6739 GND.n4859 GND.n3526 240.244
R6740 GND.n4855 GND.n3526 240.244
R6741 GND.n4855 GND.n3529 240.244
R6742 GND.n4851 GND.n3529 240.244
R6743 GND.n4851 GND.n3535 240.244
R6744 GND.n4847 GND.n3535 240.244
R6745 GND.n4847 GND.n3537 240.244
R6746 GND.n4843 GND.n3537 240.244
R6747 GND.n4843 GND.n3543 240.244
R6748 GND.n4839 GND.n3543 240.244
R6749 GND.n4839 GND.n3545 240.244
R6750 GND.n4835 GND.n3545 240.244
R6751 GND.n4835 GND.n3551 240.244
R6752 GND.n4831 GND.n3551 240.244
R6753 GND.n4831 GND.n3553 240.244
R6754 GND.n4827 GND.n3553 240.244
R6755 GND.n4827 GND.n3559 240.244
R6756 GND.n4823 GND.n3559 240.244
R6757 GND.n4823 GND.n3561 240.244
R6758 GND.n4819 GND.n3561 240.244
R6759 GND.n4819 GND.n3567 240.244
R6760 GND.n4815 GND.n3567 240.244
R6761 GND.n4815 GND.n3569 240.244
R6762 GND.n4811 GND.n3569 240.244
R6763 GND.n4811 GND.n3575 240.244
R6764 GND.n4807 GND.n3575 240.244
R6765 GND.n4807 GND.n3577 240.244
R6766 GND.n4803 GND.n3577 240.244
R6767 GND.n4803 GND.n3583 240.244
R6768 GND.n4799 GND.n3583 240.244
R6769 GND.n4799 GND.n3585 240.244
R6770 GND.n4795 GND.n3585 240.244
R6771 GND.n4795 GND.n3591 240.244
R6772 GND.n4791 GND.n3591 240.244
R6773 GND.n4791 GND.n3593 240.244
R6774 GND.n4787 GND.n3593 240.244
R6775 GND.n4787 GND.n3599 240.244
R6776 GND.n4783 GND.n3599 240.244
R6777 GND.n4783 GND.n3601 240.244
R6778 GND.n4779 GND.n3601 240.244
R6779 GND.n4779 GND.n3607 240.244
R6780 GND.n4775 GND.n3607 240.244
R6781 GND.n4775 GND.n3609 240.244
R6782 GND.n4771 GND.n3609 240.244
R6783 GND.n4771 GND.n3615 240.244
R6784 GND.n4767 GND.n3615 240.244
R6785 GND.n4767 GND.n3617 240.244
R6786 GND.n4763 GND.n3617 240.244
R6787 GND.n4763 GND.n3623 240.244
R6788 GND.n4759 GND.n3623 240.244
R6789 GND.n4759 GND.n3625 240.244
R6790 GND.n4755 GND.n3625 240.244
R6791 GND.n4755 GND.n3631 240.244
R6792 GND.n4751 GND.n3631 240.244
R6793 GND.n4751 GND.n3633 240.244
R6794 GND.n4747 GND.n3633 240.244
R6795 GND.n4747 GND.n3639 240.244
R6796 GND.n4743 GND.n3639 240.244
R6797 GND.n4743 GND.n3641 240.244
R6798 GND.n4739 GND.n3641 240.244
R6799 GND.n4739 GND.n3647 240.244
R6800 GND.n4735 GND.n3647 240.244
R6801 GND.n4735 GND.n3649 240.244
R6802 GND.n4731 GND.n3649 240.244
R6803 GND.n4731 GND.n3655 240.244
R6804 GND.n4727 GND.n3655 240.244
R6805 GND.n4727 GND.n3657 240.244
R6806 GND.n4723 GND.n3657 240.244
R6807 GND.n4723 GND.n3663 240.244
R6808 GND.n4719 GND.n3663 240.244
R6809 GND.n4719 GND.n3665 240.244
R6810 GND.n4715 GND.n3665 240.244
R6811 GND.n4715 GND.n3671 240.244
R6812 GND.n4711 GND.n3671 240.244
R6813 GND.n4711 GND.n3673 240.244
R6814 GND.n4707 GND.n3673 240.244
R6815 GND.n4707 GND.n3679 240.244
R6816 GND.n4703 GND.n3679 240.244
R6817 GND.n4703 GND.n3681 240.244
R6818 GND.n4699 GND.n3681 240.244
R6819 GND.n4699 GND.n3687 240.244
R6820 GND.n4695 GND.n3687 240.244
R6821 GND.n4695 GND.n3689 240.244
R6822 GND.n4691 GND.n3689 240.244
R6823 GND.n4691 GND.n3695 240.244
R6824 GND.n4687 GND.n3695 240.244
R6825 GND.n4687 GND.n3697 240.244
R6826 GND.n4683 GND.n3697 240.244
R6827 GND.n4683 GND.n3703 240.244
R6828 GND.n4679 GND.n3703 240.244
R6829 GND.n4679 GND.n3705 240.244
R6830 GND.n4675 GND.n3705 240.244
R6831 GND.n4675 GND.n3711 240.244
R6832 GND.n4671 GND.n3711 240.244
R6833 GND.n4671 GND.n3713 240.244
R6834 GND.n4667 GND.n3713 240.244
R6835 GND.n4667 GND.n3719 240.244
R6836 GND.n4663 GND.n3719 240.244
R6837 GND.n4663 GND.n3721 240.244
R6838 GND.n4659 GND.n3721 240.244
R6839 GND.n4659 GND.n3727 240.244
R6840 GND.n4655 GND.n3727 240.244
R6841 GND.n4655 GND.n3729 240.244
R6842 GND.n4651 GND.n3729 240.244
R6843 GND.n4651 GND.n3735 240.244
R6844 GND.n4647 GND.n3735 240.244
R6845 GND.n4647 GND.n3737 240.244
R6846 GND.n4643 GND.n3737 240.244
R6847 GND.n4643 GND.n3743 240.244
R6848 GND.n4639 GND.n3743 240.244
R6849 GND.n4639 GND.n3745 240.244
R6850 GND.n4635 GND.n3745 240.244
R6851 GND.n4635 GND.n3751 240.244
R6852 GND.n4631 GND.n3751 240.244
R6853 GND.n4631 GND.n3753 240.244
R6854 GND.n4627 GND.n3753 240.244
R6855 GND.n4627 GND.n3759 240.244
R6856 GND.n4623 GND.n3759 240.244
R6857 GND.n4623 GND.n3761 240.244
R6858 GND.n4619 GND.n3761 240.244
R6859 GND.n4619 GND.n3767 240.244
R6860 GND.n4615 GND.n3767 240.244
R6861 GND.n4615 GND.n3769 240.244
R6862 GND.n4611 GND.n3769 240.244
R6863 GND.n4611 GND.n3775 240.244
R6864 GND.n4607 GND.n3775 240.244
R6865 GND.n4607 GND.n3777 240.244
R6866 GND.n4603 GND.n3777 240.244
R6867 GND.n4603 GND.n3783 240.244
R6868 GND.n4599 GND.n3783 240.244
R6869 GND.n4599 GND.n3785 240.244
R6870 GND.n4595 GND.n3785 240.244
R6871 GND.n4595 GND.n3791 240.244
R6872 GND.n4591 GND.n3791 240.244
R6873 GND.n4591 GND.n3793 240.244
R6874 GND.n4587 GND.n3793 240.244
R6875 GND.n4587 GND.n3799 240.244
R6876 GND.n4583 GND.n3799 240.244
R6877 GND.n4583 GND.n3801 240.244
R6878 GND.n4579 GND.n3801 240.244
R6879 GND.n4579 GND.n3807 240.244
R6880 GND.n4575 GND.n3807 240.244
R6881 GND.n4575 GND.n3809 240.244
R6882 GND.n4571 GND.n3809 240.244
R6883 GND.n4571 GND.n3815 240.244
R6884 GND.n4567 GND.n3815 240.244
R6885 GND.n4567 GND.n3817 240.244
R6886 GND.n4563 GND.n3817 240.244
R6887 GND.n4563 GND.n3823 240.244
R6888 GND.n4559 GND.n3823 240.244
R6889 GND.n4559 GND.n3825 240.244
R6890 GND.n4555 GND.n3825 240.244
R6891 GND.n4555 GND.n3831 240.244
R6892 GND.n4551 GND.n3831 240.244
R6893 GND.n4551 GND.n3833 240.244
R6894 GND.n4547 GND.n3833 240.244
R6895 GND.n4547 GND.n3839 240.244
R6896 GND.n4543 GND.n3839 240.244
R6897 GND.n4543 GND.n3841 240.244
R6898 GND.n4539 GND.n3841 240.244
R6899 GND.n4539 GND.n3847 240.244
R6900 GND.n4535 GND.n3847 240.244
R6901 GND.n4535 GND.n3849 240.244
R6902 GND.n4531 GND.n3849 240.244
R6903 GND.n4531 GND.n3855 240.244
R6904 GND.n4527 GND.n3855 240.244
R6905 GND.n4527 GND.n3857 240.244
R6906 GND.n4523 GND.n3857 240.244
R6907 GND.n4523 GND.n3863 240.244
R6908 GND.n4519 GND.n3863 240.244
R6909 GND.n4519 GND.n3865 240.244
R6910 GND.n4515 GND.n3865 240.244
R6911 GND.n4515 GND.n3871 240.244
R6912 GND.n4511 GND.n3871 240.244
R6913 GND.n4511 GND.n3873 240.244
R6914 GND.n4507 GND.n3873 240.244
R6915 GND.n4507 GND.n3879 240.244
R6916 GND.n4503 GND.n3879 240.244
R6917 GND.n4503 GND.n3881 240.244
R6918 GND.n4499 GND.n3881 240.244
R6919 GND.n4499 GND.n3887 240.244
R6920 GND.n4495 GND.n3887 240.244
R6921 GND.n4495 GND.n3889 240.244
R6922 GND.n4491 GND.n3889 240.244
R6923 GND.n4491 GND.n3895 240.244
R6924 GND.n4487 GND.n3895 240.244
R6925 GND.n4487 GND.n3897 240.244
R6926 GND.n4483 GND.n3897 240.244
R6927 GND.n4483 GND.n3903 240.244
R6928 GND.n4479 GND.n3903 240.244
R6929 GND.n4479 GND.n3905 240.244
R6930 GND.n4475 GND.n3905 240.244
R6931 GND.n4475 GND.n3911 240.244
R6932 GND.n4471 GND.n3911 240.244
R6933 GND.n4471 GND.n3913 240.244
R6934 GND.n4467 GND.n3913 240.244
R6935 GND.n4467 GND.n3919 240.244
R6936 GND.n4463 GND.n3919 240.244
R6937 GND.n4463 GND.n3921 240.244
R6938 GND.n4459 GND.n3921 240.244
R6939 GND.n4459 GND.n3927 240.244
R6940 GND.n4455 GND.n3927 240.244
R6941 GND.n4455 GND.n3929 240.244
R6942 GND.n4451 GND.n3929 240.244
R6943 GND.n4451 GND.n3935 240.244
R6944 GND.n4447 GND.n3935 240.244
R6945 GND.n4447 GND.n3937 240.244
R6946 GND.n4443 GND.n3937 240.244
R6947 GND.n4443 GND.n3943 240.244
R6948 GND.n4439 GND.n3943 240.244
R6949 GND.n4439 GND.n3945 240.244
R6950 GND.n4435 GND.n3945 240.244
R6951 GND.n4435 GND.n3951 240.244
R6952 GND.n4431 GND.n3951 240.244
R6953 GND.n4431 GND.n3953 240.244
R6954 GND.n4427 GND.n3953 240.244
R6955 GND.n4427 GND.n3959 240.244
R6956 GND.n4423 GND.n3959 240.244
R6957 GND.n4423 GND.n3961 240.244
R6958 GND.n4419 GND.n3961 240.244
R6959 GND.n4419 GND.n3967 240.244
R6960 GND.n4415 GND.n3967 240.244
R6961 GND.n4415 GND.n3969 240.244
R6962 GND.n4411 GND.n3969 240.244
R6963 GND.n4411 GND.n3975 240.244
R6964 GND.n4407 GND.n3975 240.244
R6965 GND.n4407 GND.n3977 240.244
R6966 GND.n4403 GND.n3977 240.244
R6967 GND.n4403 GND.n3983 240.244
R6968 GND.n4399 GND.n3983 240.244
R6969 GND.n4399 GND.n3985 240.244
R6970 GND.n4395 GND.n3985 240.244
R6971 GND.n4395 GND.n3991 240.244
R6972 GND.n4391 GND.n3991 240.244
R6973 GND.n4391 GND.n3993 240.244
R6974 GND.n4387 GND.n3993 240.244
R6975 GND.n4387 GND.n3999 240.244
R6976 GND.n4383 GND.n3999 240.244
R6977 GND.n4383 GND.n4001 240.244
R6978 GND.n4379 GND.n4001 240.244
R6979 GND.n4379 GND.n4007 240.244
R6980 GND.n4375 GND.n4007 240.244
R6981 GND.n4375 GND.n4009 240.244
R6982 GND.n4371 GND.n4009 240.244
R6983 GND.n4371 GND.n4015 240.244
R6984 GND.n4367 GND.n4015 240.244
R6985 GND.n4367 GND.n4017 240.244
R6986 GND.n4363 GND.n4017 240.244
R6987 GND.n4363 GND.n4023 240.244
R6988 GND.n4359 GND.n4023 240.244
R6989 GND.n4359 GND.n4025 240.244
R6990 GND.n4355 GND.n4025 240.244
R6991 GND.n4355 GND.n4031 240.244
R6992 GND.n4351 GND.n4031 240.244
R6993 GND.n4351 GND.n4033 240.244
R6994 GND.n4347 GND.n4033 240.244
R6995 GND.n4347 GND.n4039 240.244
R6996 GND.n4343 GND.n4039 240.244
R6997 GND.n4343 GND.n4041 240.244
R6998 GND.n4339 GND.n4041 240.244
R6999 GND.n4339 GND.n4047 240.244
R7000 GND.n4335 GND.n4047 240.244
R7001 GND.n4335 GND.n4049 240.244
R7002 GND.n4331 GND.n4049 240.244
R7003 GND.n4331 GND.n4055 240.244
R7004 GND.n4327 GND.n4055 240.244
R7005 GND.n4327 GND.n4057 240.244
R7006 GND.n4323 GND.n4057 240.244
R7007 GND.n4323 GND.n4063 240.244
R7008 GND.n4319 GND.n4063 240.244
R7009 GND.n4319 GND.n4065 240.244
R7010 GND.n4315 GND.n4065 240.244
R7011 GND.n4315 GND.n4071 240.244
R7012 GND.n4311 GND.n4071 240.244
R7013 GND.n4311 GND.n4073 240.244
R7014 GND.n4307 GND.n4073 240.244
R7015 GND.n4303 GND.n4078 240.244
R7016 GND.n4303 GND.n4080 240.244
R7017 GND.n4297 GND.n4080 240.244
R7018 GND.n4297 GND.n4086 240.244
R7019 GND.n4293 GND.n4086 240.244
R7020 GND.n4293 GND.n4088 240.244
R7021 GND.n4289 GND.n4088 240.244
R7022 GND.n4289 GND.n4093 240.244
R7023 GND.n4285 GND.n4093 240.244
R7024 GND.n4285 GND.n4095 240.244
R7025 GND.n4281 GND.n4095 240.244
R7026 GND.n4281 GND.n4101 240.244
R7027 GND.n4277 GND.n4101 240.244
R7028 GND.n4277 GND.n4103 240.244
R7029 GND.n4273 GND.n4103 240.244
R7030 GND.n4273 GND.n4109 240.244
R7031 GND.n4269 GND.n4109 240.244
R7032 GND.n4269 GND.n4111 240.244
R7033 GND.n4265 GND.n4111 240.244
R7034 GND.n4265 GND.n4117 240.244
R7035 GND.n4261 GND.n4117 240.244
R7036 GND.n4261 GND.n4119 240.244
R7037 GND.n4257 GND.n4119 240.244
R7038 GND.n4257 GND.n4125 240.244
R7039 GND.n4253 GND.n4125 240.244
R7040 GND.n4253 GND.n4127 240.244
R7041 GND.n4249 GND.n4127 240.244
R7042 GND.n4249 GND.n4133 240.244
R7043 GND.n4245 GND.n4133 240.244
R7044 GND.n4245 GND.n4135 240.244
R7045 GND.n4241 GND.n4135 240.244
R7046 GND.n4241 GND.n4141 240.244
R7047 GND.n4237 GND.n4141 240.244
R7048 GND.n4237 GND.n4143 240.244
R7049 GND.n4233 GND.n4143 240.244
R7050 GND.n4233 GND.n4149 240.244
R7051 GND.n4229 GND.n4149 240.244
R7052 GND.n4229 GND.n4151 240.244
R7053 GND.n4225 GND.n4151 240.244
R7054 GND.n4225 GND.n4157 240.244
R7055 GND.n4221 GND.n4157 240.244
R7056 GND.n4221 GND.n4159 240.244
R7057 GND.n4217 GND.n4159 240.244
R7058 GND.n4217 GND.n4165 240.244
R7059 GND.n4213 GND.n4165 240.244
R7060 GND.n4213 GND.n4167 240.244
R7061 GND.n4209 GND.n4167 240.244
R7062 GND.n4209 GND.n4173 240.244
R7063 GND.n4205 GND.n4173 240.244
R7064 GND.n4205 GND.n4175 240.244
R7065 GND.n4201 GND.n4175 240.244
R7066 GND.n4201 GND.n4181 240.244
R7067 GND.n4197 GND.n4181 240.244
R7068 GND.n4197 GND.n4183 240.244
R7069 GND.n4193 GND.n4183 240.244
R7070 GND.n4193 GND.n4191 240.244
R7071 GND.n5033 GND.n2770 240.244
R7072 GND.n5051 GND.n2770 240.244
R7073 GND.n5051 GND.n2766 240.244
R7074 GND.n5057 GND.n2766 240.244
R7075 GND.n5057 GND.n2538 240.244
R7076 GND.n5211 GND.n2538 240.244
R7077 GND.n5211 GND.n2539 240.244
R7078 GND.n2539 GND.n2533 240.244
R7079 GND.n5219 GND.n2533 240.244
R7080 GND.n5219 GND.n2534 240.244
R7081 GND.n2735 GND.n2534 240.244
R7082 GND.n5076 GND.n2735 240.244
R7083 GND.n5078 GND.n5076 240.244
R7084 GND.n5081 GND.n5078 240.244
R7085 GND.n5081 GND.n2713 240.244
R7086 GND.n5176 GND.n2713 240.244
R7087 GND.n5179 GND.n5176 240.244
R7088 GND.n5181 GND.n5179 240.244
R7089 GND.n5181 GND.n2510 240.244
R7090 GND.n5228 GND.n2510 240.244
R7091 GND.n5228 GND.n2494 240.244
R7092 GND.n5242 GND.n2494 240.244
R7093 GND.n5242 GND.n2490 240.244
R7094 GND.n5248 GND.n2490 240.244
R7095 GND.n5248 GND.n2474 240.244
R7096 GND.n5262 GND.n2474 240.244
R7097 GND.n5262 GND.n2470 240.244
R7098 GND.n5268 GND.n2470 240.244
R7099 GND.n5268 GND.n2453 240.244
R7100 GND.n5282 GND.n2453 240.244
R7101 GND.n5282 GND.n2449 240.244
R7102 GND.n5288 GND.n2449 240.244
R7103 GND.n5288 GND.n2434 240.244
R7104 GND.n5302 GND.n2434 240.244
R7105 GND.n5302 GND.n2430 240.244
R7106 GND.n5308 GND.n2430 240.244
R7107 GND.n5308 GND.n2414 240.244
R7108 GND.n5322 GND.n2414 240.244
R7109 GND.n5322 GND.n2410 240.244
R7110 GND.n5328 GND.n2410 240.244
R7111 GND.n5328 GND.n2393 240.244
R7112 GND.n5342 GND.n2393 240.244
R7113 GND.n5342 GND.n2389 240.244
R7114 GND.n5348 GND.n2389 240.244
R7115 GND.n5348 GND.n2374 240.244
R7116 GND.n5362 GND.n2374 240.244
R7117 GND.n5362 GND.n2370 240.244
R7118 GND.n5368 GND.n2370 240.244
R7119 GND.n5368 GND.n2354 240.244
R7120 GND.n5387 GND.n2354 240.244
R7121 GND.n5387 GND.n2349 240.244
R7122 GND.n5395 GND.n2349 240.244
R7123 GND.n5395 GND.n2350 240.244
R7124 GND.n2350 GND.n2327 240.244
R7125 GND.n5467 GND.n2327 240.244
R7126 GND.n5467 GND.n2323 240.244
R7127 GND.n5473 GND.n2323 240.244
R7128 GND.n5473 GND.n2307 240.244
R7129 GND.n5487 GND.n2307 240.244
R7130 GND.n5487 GND.n2303 240.244
R7131 GND.n5493 GND.n2303 240.244
R7132 GND.n5493 GND.n2287 240.244
R7133 GND.n5507 GND.n2287 240.244
R7134 GND.n5507 GND.n2283 240.244
R7135 GND.n5513 GND.n2283 240.244
R7136 GND.n5513 GND.n2266 240.244
R7137 GND.n5527 GND.n2266 240.244
R7138 GND.n5527 GND.n2262 240.244
R7139 GND.n5533 GND.n2262 240.244
R7140 GND.n5533 GND.n2247 240.244
R7141 GND.n5551 GND.n2247 240.244
R7142 GND.n5551 GND.n2243 240.244
R7143 GND.n5558 GND.n2243 240.244
R7144 GND.n5558 GND.n1742 240.244
R7145 GND.n5690 GND.n1742 240.244
R7146 GND.n5690 GND.n1743 240.244
R7147 GND.n5686 GND.n1743 240.244
R7148 GND.n5686 GND.n1749 240.244
R7149 GND.n5682 GND.n1749 240.244
R7150 GND.n5682 GND.n1779 240.244
R7151 GND.n5678 GND.n1779 240.244
R7152 GND.n5678 GND.n1785 240.244
R7153 GND.n2180 GND.n1785 240.244
R7154 GND.n2180 GND.n1825 240.244
R7155 GND.n2176 GND.n1825 240.244
R7156 GND.n2176 GND.n1831 240.244
R7157 GND.n2166 GND.n1831 240.244
R7158 GND.n2166 GND.n1843 240.244
R7159 GND.n2162 GND.n1843 240.244
R7160 GND.n2162 GND.n1849 240.244
R7161 GND.n2152 GND.n1849 240.244
R7162 GND.n2152 GND.n1861 240.244
R7163 GND.n2148 GND.n1861 240.244
R7164 GND.n2148 GND.n1867 240.244
R7165 GND.n2138 GND.n1867 240.244
R7166 GND.n2138 GND.n1879 240.244
R7167 GND.n2134 GND.n1879 240.244
R7168 GND.n2134 GND.n1885 240.244
R7169 GND.n2124 GND.n1885 240.244
R7170 GND.n2124 GND.n1898 240.244
R7171 GND.n2120 GND.n1898 240.244
R7172 GND.n2120 GND.n1904 240.244
R7173 GND.n2110 GND.n1904 240.244
R7174 GND.n2110 GND.n1916 240.244
R7175 GND.n2106 GND.n1916 240.244
R7176 GND.n2106 GND.n1922 240.244
R7177 GND.n2096 GND.n1922 240.244
R7178 GND.n2096 GND.n1934 240.244
R7179 GND.n2092 GND.n1934 240.244
R7180 GND.n2092 GND.n1940 240.244
R7181 GND.n2082 GND.n1940 240.244
R7182 GND.n2082 GND.n1952 240.244
R7183 GND.n2078 GND.n1952 240.244
R7184 GND.n2078 GND.n1965 240.244
R7185 GND.n1965 GND.n1964 240.244
R7186 GND.n1964 GND.n1958 240.244
R7187 GND.n1958 GND.n1701 240.244
R7188 GND.n5784 GND.n1701 240.244
R7189 GND.n5784 GND.n1696 240.244
R7190 GND.n5807 GND.n1696 240.244
R7191 GND.n5807 GND.n1697 240.244
R7192 GND.n5803 GND.n1697 240.244
R7193 GND.n5803 GND.n5802 240.244
R7194 GND.n5802 GND.n5801 240.244
R7195 GND.n5801 GND.n5792 240.244
R7196 GND.n5792 GND.n1617 240.244
R7197 GND.n5907 GND.n1617 240.244
R7198 GND.n5908 GND.n5907 240.244
R7199 GND.n5909 GND.n5908 240.244
R7200 GND.n5909 GND.n1613 240.244
R7201 GND.n5915 GND.n1613 240.244
R7202 GND.n5915 GND.n1561 240.244
R7203 GND.n5987 GND.n1561 240.244
R7204 GND.n5987 GND.n1556 240.244
R7205 GND.n6004 GND.n1556 240.244
R7206 GND.n6004 GND.n1557 240.244
R7207 GND.n6000 GND.n1557 240.244
R7208 GND.n6000 GND.n5999 240.244
R7209 GND.n5999 GND.n5998 240.244
R7210 GND.n5998 GND.n1517 240.244
R7211 GND.n6077 GND.n1517 240.244
R7212 GND.n6077 GND.n1512 240.244
R7213 GND.n6085 GND.n1512 240.244
R7214 GND.n6085 GND.n1513 240.244
R7215 GND.n1513 GND.n1482 240.244
R7216 GND.n6143 GND.n1482 240.244
R7217 GND.n6143 GND.n1478 240.244
R7218 GND.n6149 GND.n1478 240.244
R7219 GND.n6149 GND.n1458 240.244
R7220 GND.n6186 GND.n1458 240.244
R7221 GND.n6186 GND.n1454 240.244
R7222 GND.n6194 GND.n1454 240.244
R7223 GND.n6194 GND.n1442 240.244
R7224 GND.n6245 GND.n1442 240.244
R7225 GND.n6246 GND.n6245 240.244
R7226 GND.n6246 GND.n1438 240.244
R7227 GND.n6252 GND.n1438 240.244
R7228 GND.n6252 GND.n1330 240.244
R7229 GND.n6318 GND.n1330 240.244
R7230 GND.n6318 GND.n1324 240.244
R7231 GND.n6329 GND.n1324 240.244
R7232 GND.n6329 GND.n1326 240.244
R7233 GND.n6325 GND.n1326 240.244
R7234 GND.n6325 GND.n1307 240.244
R7235 GND.n6358 GND.n1307 240.244
R7236 GND.n6358 GND.n1302 240.244
R7237 GND.n6375 GND.n1302 240.244
R7238 GND.n6375 GND.n1303 240.244
R7239 GND.n6371 GND.n1303 240.244
R7240 GND.n6371 GND.n6370 240.244
R7241 GND.n6370 GND.n6369 240.244
R7242 GND.n6369 GND.n1273 240.244
R7243 GND.n6416 GND.n1273 240.244
R7244 GND.n6416 GND.n1268 240.244
R7245 GND.n6424 GND.n1268 240.244
R7246 GND.n6424 GND.n1269 240.244
R7247 GND.n1269 GND.n1248 240.244
R7248 GND.n6451 GND.n1248 240.244
R7249 GND.n6451 GND.n1243 240.244
R7250 GND.n6462 GND.n1243 240.244
R7251 GND.n6462 GND.n1244 240.244
R7252 GND.n6458 GND.n1244 240.244
R7253 GND.n6458 GND.n1223 240.244
R7254 GND.n6490 GND.n1223 240.244
R7255 GND.n6490 GND.n1218 240.244
R7256 GND.n6507 GND.n1218 240.244
R7257 GND.n6507 GND.n1219 240.244
R7258 GND.n6503 GND.n1219 240.244
R7259 GND.n6503 GND.n6502 240.244
R7260 GND.n6502 GND.n6501 240.244
R7261 GND.n6501 GND.n1189 240.244
R7262 GND.n6595 GND.n1189 240.244
R7263 GND.n6595 GND.n1184 240.244
R7264 GND.n6615 GND.n1184 240.244
R7265 GND.n6615 GND.n1185 240.244
R7266 GND.n6611 GND.n1185 240.244
R7267 GND.n6611 GND.n6603 240.244
R7268 GND.n6607 GND.n6603 240.244
R7269 GND.n6607 GND.n939 240.244
R7270 GND.n6727 GND.n939 240.244
R7271 GND.n6727 GND.n935 240.244
R7272 GND.n6733 GND.n935 240.244
R7273 GND.n6733 GND.n917 240.244
R7274 GND.n6753 GND.n917 240.244
R7275 GND.n6753 GND.n912 240.244
R7276 GND.n6761 GND.n912 240.244
R7277 GND.n6761 GND.n913 240.244
R7278 GND.n913 GND.n890 240.244
R7279 GND.n6864 GND.n890 240.244
R7280 GND.n6864 GND.n886 240.244
R7281 GND.n6870 GND.n886 240.244
R7282 GND.n6870 GND.n870 240.244
R7283 GND.n6884 GND.n870 240.244
R7284 GND.n6884 GND.n866 240.244
R7285 GND.n6890 GND.n866 240.244
R7286 GND.n6890 GND.n850 240.244
R7287 GND.n6904 GND.n850 240.244
R7288 GND.n6904 GND.n846 240.244
R7289 GND.n6910 GND.n846 240.244
R7290 GND.n6910 GND.n829 240.244
R7291 GND.n6924 GND.n829 240.244
R7292 GND.n6924 GND.n825 240.244
R7293 GND.n6930 GND.n825 240.244
R7294 GND.n6930 GND.n810 240.244
R7295 GND.n6944 GND.n810 240.244
R7296 GND.n6944 GND.n806 240.244
R7297 GND.n6950 GND.n806 240.244
R7298 GND.n6950 GND.n790 240.244
R7299 GND.n6964 GND.n790 240.244
R7300 GND.n6964 GND.n786 240.244
R7301 GND.n6970 GND.n786 240.244
R7302 GND.n6970 GND.n770 240.244
R7303 GND.n6984 GND.n770 240.244
R7304 GND.n6984 GND.n766 240.244
R7305 GND.n6990 GND.n766 240.244
R7306 GND.n6990 GND.n750 240.244
R7307 GND.n7004 GND.n750 240.244
R7308 GND.n7004 GND.n746 240.244
R7309 GND.n7010 GND.n746 240.244
R7310 GND.n7010 GND.n729 240.244
R7311 GND.n7028 GND.n729 240.244
R7312 GND.n7028 GND.n724 240.244
R7313 GND.n7036 GND.n724 240.244
R7314 GND.n7036 GND.n725 240.244
R7315 GND.n725 GND.n702 240.244
R7316 GND.n7072 GND.n702 240.244
R7317 GND.n7072 GND.n698 240.244
R7318 GND.n7078 GND.n698 240.244
R7319 GND.n7078 GND.n681 240.244
R7320 GND.n7100 GND.n681 240.244
R7321 GND.n7100 GND.n677 240.244
R7322 GND.n7106 GND.n677 240.244
R7323 GND.n7106 GND.n652 240.244
R7324 GND.n7136 GND.n652 240.244
R7325 GND.n7136 GND.n653 240.244
R7326 GND.n653 GND.n648 240.244
R7327 GND.n7144 GND.n648 240.244
R7328 GND.n7144 GND.n634 240.244
R7329 GND.n7161 GND.n634 240.244
R7330 GND.n7164 GND.n7161 240.244
R7331 GND.n7167 GND.n7164 240.244
R7332 GND.n7167 GND.n238 240.244
R7333 GND.n7640 GND.n238 240.244
R7334 GND.n7640 GND.n239 240.244
R7335 GND.n7205 GND.n239 240.244
R7336 GND.n7207 GND.n7205 240.244
R7337 GND.n7207 GND.n250 240.244
R7338 GND.n7633 GND.n250 240.244
R7339 GND.n7633 GND.n251 240.244
R7340 GND.n7625 GND.n251 240.244
R7341 GND.n7625 GND.n269 240.244
R7342 GND.n7621 GND.n269 240.244
R7343 GND.n7621 GND.n274 240.244
R7344 GND.n7613 GND.n274 240.244
R7345 GND.n7613 GND.n289 240.244
R7346 GND.n7609 GND.n289 240.244
R7347 GND.n7609 GND.n295 240.244
R7348 GND.n3522 GND.n3521 240.244
R7349 GND.n5018 GND.n3521 240.244
R7350 GND.n5016 GND.n5015 240.244
R7351 GND.n5012 GND.n5011 240.244
R7352 GND.n5008 GND.n5007 240.244
R7353 GND.n5004 GND.n5003 240.244
R7354 GND.n5000 GND.n4999 240.244
R7355 GND.n4996 GND.n4995 240.244
R7356 GND.n4992 GND.n4991 240.244
R7357 GND.n4988 GND.n4987 240.244
R7358 GND.n4984 GND.n4983 240.244
R7359 GND.n4980 GND.n4979 240.244
R7360 GND.n4976 GND.n4975 240.244
R7361 GND.n4972 GND.n4971 240.244
R7362 GND.n4968 GND.n4967 240.244
R7363 GND.n4964 GND.n4963 240.244
R7364 GND.n4960 GND.n4959 240.244
R7365 GND.n4956 GND.n4955 240.244
R7366 GND.n4952 GND.n4951 240.244
R7367 GND.n4948 GND.n4947 240.244
R7368 GND.n4944 GND.n4943 240.244
R7369 GND.n4940 GND.n4939 240.244
R7370 GND.n4936 GND.n4935 240.244
R7371 GND.n4932 GND.n4931 240.244
R7372 GND.n4928 GND.n4927 240.244
R7373 GND.n4924 GND.n4923 240.244
R7374 GND.n4920 GND.n4919 240.244
R7375 GND.n5027 GND.n2789 240.244
R7376 GND.n5566 GND.n5565 240.244
R7377 GND.n5573 GND.n5572 240.244
R7378 GND.n5576 GND.n5575 240.244
R7379 GND.n5584 GND.n5583 240.244
R7380 GND.n5588 GND.n5587 240.244
R7381 GND.n5593 GND.n5592 240.244
R7382 GND.n5596 GND.n5595 240.244
R7383 GND.n5601 GND.n5600 240.244
R7384 GND.n5604 GND.n5603 240.244
R7385 GND.n5611 GND.n5609 240.244
R7386 GND.n3187 GND.n3186 240.244
R7387 GND.n3187 GND.n3040 240.244
R7388 GND.n3189 GND.n3040 240.244
R7389 GND.n3189 GND.n3031 240.244
R7390 GND.n3031 GND.n3022 240.244
R7391 GND.n3326 GND.n3022 240.244
R7392 GND.n3326 GND.n3011 240.244
R7393 GND.n3011 GND.n3002 240.244
R7394 GND.n3342 GND.n3002 240.244
R7395 GND.n3343 GND.n3342 240.244
R7396 GND.n3343 GND.n2991 240.244
R7397 GND.n2991 GND.n2981 240.244
R7398 GND.n3359 GND.n2981 240.244
R7399 GND.n3360 GND.n3359 240.244
R7400 GND.n3360 GND.n2970 240.244
R7401 GND.n2970 GND.n2960 240.244
R7402 GND.n3376 GND.n2960 240.244
R7403 GND.n3377 GND.n3376 240.244
R7404 GND.n3377 GND.n2948 240.244
R7405 GND.n2948 GND.n2939 240.244
R7406 GND.n3393 GND.n2939 240.244
R7407 GND.n3394 GND.n3393 240.244
R7408 GND.n3394 GND.n2928 240.244
R7409 GND.n2928 GND.n2918 240.244
R7410 GND.n3410 GND.n2918 240.244
R7411 GND.n3411 GND.n3410 240.244
R7412 GND.n3411 GND.n2907 240.244
R7413 GND.n2907 GND.n2897 240.244
R7414 GND.n3427 GND.n2897 240.244
R7415 GND.n3428 GND.n3427 240.244
R7416 GND.n3428 GND.n2886 240.244
R7417 GND.n2886 GND.n2876 240.244
R7418 GND.n3444 GND.n2876 240.244
R7419 GND.n3445 GND.n3444 240.244
R7420 GND.n3445 GND.n2865 240.244
R7421 GND.n2865 GND.n2855 240.244
R7422 GND.n3461 GND.n2855 240.244
R7423 GND.n3462 GND.n3461 240.244
R7424 GND.n3462 GND.n2844 240.244
R7425 GND.n2844 GND.n2834 240.244
R7426 GND.n3478 GND.n2834 240.244
R7427 GND.n3479 GND.n3478 240.244
R7428 GND.n3479 GND.n2825 240.244
R7429 GND.n3481 GND.n2825 240.244
R7430 GND.n3481 GND.n2817 240.244
R7431 GND.n2817 GND.n2785 240.244
R7432 GND.n2785 GND.n2775 240.244
R7433 GND.n5049 GND.n2775 240.244
R7434 GND.n5049 GND.n2776 240.244
R7435 GND.n2776 GND.n2765 240.244
R7436 GND.n2765 GND.n2545 240.244
R7437 GND.n5209 GND.n2545 240.244
R7438 GND.n5209 GND.n2546 240.244
R7439 GND.n2554 GND.n2546 240.244
R7440 GND.n2554 GND.n2532 240.244
R7441 GND.n2555 GND.n2532 240.244
R7442 GND.n2736 GND.n2555 240.244
R7443 GND.n2736 GND.n2562 240.244
R7444 GND.n2563 GND.n2562 240.244
R7445 GND.n2564 GND.n2563 240.244
R7446 GND.n2714 GND.n2564 240.244
R7447 GND.n2714 GND.n2570 240.244
R7448 GND.n2571 GND.n2570 240.244
R7449 GND.n2572 GND.n2571 240.244
R7450 GND.n2573 GND.n2572 240.244
R7451 GND.n2573 GND.n2509 240.244
R7452 GND.n2509 GND.n2499 240.244
R7453 GND.n5240 GND.n2499 240.244
R7454 GND.n5240 GND.n2500 240.244
R7455 GND.n2500 GND.n2489 240.244
R7456 GND.n2489 GND.n2479 240.244
R7457 GND.n5260 GND.n2479 240.244
R7458 GND.n5260 GND.n2480 240.244
R7459 GND.n2480 GND.n2469 240.244
R7460 GND.n2469 GND.n2459 240.244
R7461 GND.n5280 GND.n2459 240.244
R7462 GND.n5280 GND.n2460 240.244
R7463 GND.n2460 GND.n2448 240.244
R7464 GND.n2448 GND.n2439 240.244
R7465 GND.n5300 GND.n2439 240.244
R7466 GND.n5300 GND.n2440 240.244
R7467 GND.n2440 GND.n2429 240.244
R7468 GND.n2429 GND.n2419 240.244
R7469 GND.n5320 GND.n2419 240.244
R7470 GND.n5320 GND.n2420 240.244
R7471 GND.n2420 GND.n2409 240.244
R7472 GND.n2409 GND.n2399 240.244
R7473 GND.n5340 GND.n2399 240.244
R7474 GND.n5340 GND.n2400 240.244
R7475 GND.n2400 GND.n2388 240.244
R7476 GND.n2388 GND.n2379 240.244
R7477 GND.n5360 GND.n2379 240.244
R7478 GND.n5360 GND.n2380 240.244
R7479 GND.n2380 GND.n2369 240.244
R7480 GND.n2369 GND.n2359 240.244
R7481 GND.n5385 GND.n2359 240.244
R7482 GND.n5385 GND.n2360 240.244
R7483 GND.n2360 GND.n2348 240.244
R7484 GND.n5378 GND.n2348 240.244
R7485 GND.n5378 GND.n2331 240.244
R7486 GND.n5465 GND.n2331 240.244
R7487 GND.n5465 GND.n2332 240.244
R7488 GND.n2332 GND.n2322 240.244
R7489 GND.n2322 GND.n2312 240.244
R7490 GND.n5485 GND.n2312 240.244
R7491 GND.n5485 GND.n2313 240.244
R7492 GND.n2313 GND.n2302 240.244
R7493 GND.n2302 GND.n2292 240.244
R7494 GND.n5505 GND.n2292 240.244
R7495 GND.n5505 GND.n2293 240.244
R7496 GND.n2293 GND.n2282 240.244
R7497 GND.n2282 GND.n2272 240.244
R7498 GND.n5525 GND.n2272 240.244
R7499 GND.n5525 GND.n2273 240.244
R7500 GND.n2273 GND.n2261 240.244
R7501 GND.n2261 GND.n2252 240.244
R7502 GND.n5549 GND.n2252 240.244
R7503 GND.n5549 GND.n2253 240.244
R7504 GND.n2253 GND.n2242 240.244
R7505 GND.n2242 GND.n1735 240.244
R7506 GND.n5692 GND.n1735 240.244
R7507 GND.n3178 GND.n3176 240.244
R7508 GND.n3176 GND.n3175 240.244
R7509 GND.n3172 GND.n3171 240.244
R7510 GND.n3169 GND.n3061 240.244
R7511 GND.n3165 GND.n3163 240.244
R7512 GND.n3161 GND.n3069 240.244
R7513 GND.n3157 GND.n3155 240.244
R7514 GND.n3153 GND.n3075 240.244
R7515 GND.n3149 GND.n3147 240.244
R7516 GND.n3145 GND.n3081 240.244
R7517 GND.n3085 GND.n3049 240.244
R7518 GND.n3184 GND.n3038 240.244
R7519 GND.n3202 GND.n3038 240.244
R7520 GND.n3202 GND.n3033 240.244
R7521 GND.n3210 GND.n3033 240.244
R7522 GND.n3210 GND.n3034 240.244
R7523 GND.n3034 GND.n3010 240.244
R7524 GND.n3334 GND.n3010 240.244
R7525 GND.n3334 GND.n3006 240.244
R7526 GND.n3340 GND.n3006 240.244
R7527 GND.n3340 GND.n2989 240.244
R7528 GND.n3351 GND.n2989 240.244
R7529 GND.n3351 GND.n2985 240.244
R7530 GND.n3357 GND.n2985 240.244
R7531 GND.n3357 GND.n2968 240.244
R7532 GND.n3368 GND.n2968 240.244
R7533 GND.n3368 GND.n2964 240.244
R7534 GND.n3374 GND.n2964 240.244
R7535 GND.n3374 GND.n2946 240.244
R7536 GND.n3385 GND.n2946 240.244
R7537 GND.n3385 GND.n2942 240.244
R7538 GND.n3391 GND.n2942 240.244
R7539 GND.n3391 GND.n2926 240.244
R7540 GND.n3402 GND.n2926 240.244
R7541 GND.n3402 GND.n2922 240.244
R7542 GND.n3408 GND.n2922 240.244
R7543 GND.n3408 GND.n2905 240.244
R7544 GND.n3419 GND.n2905 240.244
R7545 GND.n3419 GND.n2901 240.244
R7546 GND.n3425 GND.n2901 240.244
R7547 GND.n3425 GND.n2884 240.244
R7548 GND.n3436 GND.n2884 240.244
R7549 GND.n3436 GND.n2880 240.244
R7550 GND.n3442 GND.n2880 240.244
R7551 GND.n3442 GND.n2863 240.244
R7552 GND.n3453 GND.n2863 240.244
R7553 GND.n3453 GND.n2859 240.244
R7554 GND.n3459 GND.n2859 240.244
R7555 GND.n3459 GND.n2842 240.244
R7556 GND.n3470 GND.n2842 240.244
R7557 GND.n3470 GND.n2838 240.244
R7558 GND.n3476 GND.n2838 240.244
R7559 GND.n3476 GND.n2823 240.244
R7560 GND.n3493 GND.n2823 240.244
R7561 GND.n3493 GND.n2819 240.244
R7562 GND.n3519 GND.n2819 240.244
R7563 GND.n3519 GND.n2783 240.244
R7564 GND.n3515 GND.n2783 240.244
R7565 GND.n3515 GND.n2772 240.244
R7566 GND.n3512 GND.n2772 240.244
R7567 GND.n3512 GND.n2763 240.244
R7568 GND.n3509 GND.n2763 240.244
R7569 GND.n3509 GND.n2541 240.244
R7570 GND.n3506 GND.n2541 240.244
R7571 GND.n3506 GND.n2527 240.244
R7572 GND.n5221 GND.n2527 240.244
R7573 GND.n5221 GND.n2528 240.244
R7574 GND.n2738 GND.n2528 240.244
R7575 GND.n2744 GND.n2738 240.244
R7576 GND.n2744 GND.n2741 240.244
R7577 GND.n2741 GND.n2731 240.244
R7578 GND.n2731 GND.n2730 240.244
R7579 GND.n2730 GND.n2719 240.244
R7580 GND.n2719 GND.n2718 240.244
R7581 GND.n2718 GND.n2711 240.244
R7582 GND.n2711 GND.n2710 240.244
R7583 GND.n2710 GND.n2507 240.244
R7584 GND.n2706 GND.n2507 240.244
R7585 GND.n2706 GND.n2496 240.244
R7586 GND.n2703 GND.n2496 240.244
R7587 GND.n2703 GND.n2487 240.244
R7588 GND.n2700 GND.n2487 240.244
R7589 GND.n2700 GND.n2476 240.244
R7590 GND.n2697 GND.n2476 240.244
R7591 GND.n2697 GND.n2467 240.244
R7592 GND.n2694 GND.n2467 240.244
R7593 GND.n2694 GND.n2455 240.244
R7594 GND.n2691 GND.n2455 240.244
R7595 GND.n2691 GND.n2446 240.244
R7596 GND.n2688 GND.n2446 240.244
R7597 GND.n2688 GND.n2436 240.244
R7598 GND.n2685 GND.n2436 240.244
R7599 GND.n2685 GND.n2427 240.244
R7600 GND.n2682 GND.n2427 240.244
R7601 GND.n2682 GND.n2416 240.244
R7602 GND.n2679 GND.n2416 240.244
R7603 GND.n2679 GND.n2407 240.244
R7604 GND.n2676 GND.n2407 240.244
R7605 GND.n2676 GND.n2395 240.244
R7606 GND.n2673 GND.n2395 240.244
R7607 GND.n2673 GND.n2386 240.244
R7608 GND.n2670 GND.n2386 240.244
R7609 GND.n2670 GND.n2376 240.244
R7610 GND.n2667 GND.n2376 240.244
R7611 GND.n2667 GND.n2367 240.244
R7612 GND.n2664 GND.n2367 240.244
R7613 GND.n2664 GND.n2356 240.244
R7614 GND.n2661 GND.n2356 240.244
R7615 GND.n2661 GND.n2346 240.244
R7616 GND.n2658 GND.n2346 240.244
R7617 GND.n2658 GND.n2339 240.244
R7618 GND.n2339 GND.n2328 240.244
R7619 GND.n2654 GND.n2328 240.244
R7620 GND.n2654 GND.n2320 240.244
R7621 GND.n2651 GND.n2320 240.244
R7622 GND.n2651 GND.n2309 240.244
R7623 GND.n2648 GND.n2309 240.244
R7624 GND.n2648 GND.n2300 240.244
R7625 GND.n2645 GND.n2300 240.244
R7626 GND.n2645 GND.n2289 240.244
R7627 GND.n2642 GND.n2289 240.244
R7628 GND.n2642 GND.n2280 240.244
R7629 GND.n2639 GND.n2280 240.244
R7630 GND.n2639 GND.n2268 240.244
R7631 GND.n2636 GND.n2268 240.244
R7632 GND.n2636 GND.n2259 240.244
R7633 GND.n2633 GND.n2259 240.244
R7634 GND.n2633 GND.n2249 240.244
R7635 GND.n2249 GND.n2238 240.244
R7636 GND.n5560 GND.n2238 240.244
R7637 GND.n5561 GND.n5560 240.244
R7638 GND.n5561 GND.n1738 240.244
R7639 GND.n1776 GND.n1775 240.244
R7640 GND.n1772 GND.n1771 240.244
R7641 GND.n1768 GND.n1767 240.244
R7642 GND.n1764 GND.n1763 240.244
R7643 GND.n1760 GND.n1759 240.244
R7644 GND.n3107 GND.n3051 240.244
R7645 GND.n3107 GND.n3041 240.244
R7646 GND.n3041 GND.n3029 240.244
R7647 GND.n3212 GND.n3029 240.244
R7648 GND.n3212 GND.n3024 240.244
R7649 GND.n3324 GND.n3024 240.244
R7650 GND.n3324 GND.n3012 240.244
R7651 GND.n3217 GND.n3012 240.244
R7652 GND.n3217 GND.n3004 240.244
R7653 GND.n3218 GND.n3004 240.244
R7654 GND.n3218 GND.n2992 240.244
R7655 GND.n3221 GND.n2992 240.244
R7656 GND.n3221 GND.n2983 240.244
R7657 GND.n3222 GND.n2983 240.244
R7658 GND.n3222 GND.n2971 240.244
R7659 GND.n3225 GND.n2971 240.244
R7660 GND.n3225 GND.n2962 240.244
R7661 GND.n3226 GND.n2962 240.244
R7662 GND.n3226 GND.n2949 240.244
R7663 GND.n3229 GND.n2949 240.244
R7664 GND.n3229 GND.n2940 240.244
R7665 GND.n3230 GND.n2940 240.244
R7666 GND.n3230 GND.n2929 240.244
R7667 GND.n3233 GND.n2929 240.244
R7668 GND.n3233 GND.n2920 240.244
R7669 GND.n3234 GND.n2920 240.244
R7670 GND.n3234 GND.n2908 240.244
R7671 GND.n3237 GND.n2908 240.244
R7672 GND.n3237 GND.n2899 240.244
R7673 GND.n3238 GND.n2899 240.244
R7674 GND.n3238 GND.n2887 240.244
R7675 GND.n3241 GND.n2887 240.244
R7676 GND.n3241 GND.n2878 240.244
R7677 GND.n3242 GND.n2878 240.244
R7678 GND.n3242 GND.n2866 240.244
R7679 GND.n3245 GND.n2866 240.244
R7680 GND.n3245 GND.n2857 240.244
R7681 GND.n3246 GND.n2857 240.244
R7682 GND.n3246 GND.n2845 240.244
R7683 GND.n3249 GND.n2845 240.244
R7684 GND.n3249 GND.n2836 240.244
R7685 GND.n3250 GND.n2836 240.244
R7686 GND.n3250 GND.n2826 240.244
R7687 GND.n3253 GND.n2826 240.244
R7688 GND.n3253 GND.n2818 240.244
R7689 GND.n2818 GND.n2784 240.244
R7690 GND.n3254 GND.n2784 240.244
R7691 GND.n3254 GND.n2774 240.244
R7692 GND.n2774 GND.n2761 240.244
R7693 GND.n5059 GND.n2761 240.244
R7694 GND.n5060 GND.n5059 240.244
R7695 GND.n5060 GND.n2544 240.244
R7696 GND.n2754 GND.n2544 240.244
R7697 GND.n2758 GND.n2754 240.244
R7698 GND.n2758 GND.n2531 240.244
R7699 GND.n5068 GND.n2531 240.244
R7700 GND.n5068 GND.n2750 240.244
R7701 GND.n5074 GND.n2750 240.244
R7702 GND.n5074 GND.n2726 240.244
R7703 GND.n5083 GND.n2726 240.244
R7704 GND.n5083 GND.n2721 240.244
R7705 GND.n5174 GND.n2721 240.244
R7706 GND.n5174 GND.n2722 240.244
R7707 GND.n2722 GND.n2712 240.244
R7708 GND.n5169 GND.n2712 240.244
R7709 GND.n5169 GND.n2508 240.244
R7710 GND.n5166 GND.n2508 240.244
R7711 GND.n5166 GND.n2498 240.244
R7712 GND.n5163 GND.n2498 240.244
R7713 GND.n5163 GND.n2488 240.244
R7714 GND.n5160 GND.n2488 240.244
R7715 GND.n5160 GND.n2478 240.244
R7716 GND.n5157 GND.n2478 240.244
R7717 GND.n5157 GND.n2468 240.244
R7718 GND.n5154 GND.n2468 240.244
R7719 GND.n5154 GND.n2458 240.244
R7720 GND.n5151 GND.n2458 240.244
R7721 GND.n5151 GND.n2447 240.244
R7722 GND.n5148 GND.n2447 240.244
R7723 GND.n5148 GND.n2438 240.244
R7724 GND.n5145 GND.n2438 240.244
R7725 GND.n5145 GND.n2428 240.244
R7726 GND.n5142 GND.n2428 240.244
R7727 GND.n5142 GND.n2418 240.244
R7728 GND.n5139 GND.n2418 240.244
R7729 GND.n5139 GND.n2408 240.244
R7730 GND.n5136 GND.n2408 240.244
R7731 GND.n5136 GND.n2398 240.244
R7732 GND.n5133 GND.n2398 240.244
R7733 GND.n5133 GND.n2387 240.244
R7734 GND.n5130 GND.n2387 240.244
R7735 GND.n5130 GND.n2378 240.244
R7736 GND.n5127 GND.n2378 240.244
R7737 GND.n5127 GND.n2368 240.244
R7738 GND.n5124 GND.n2368 240.244
R7739 GND.n5124 GND.n2358 240.244
R7740 GND.n2358 GND.n2344 240.244
R7741 GND.n5397 GND.n2344 240.244
R7742 GND.n5397 GND.n2340 240.244
R7743 GND.n5454 GND.n2340 240.244
R7744 GND.n5454 GND.n2330 240.244
R7745 GND.n5450 GND.n2330 240.244
R7746 GND.n5450 GND.n2321 240.244
R7747 GND.n5447 GND.n2321 240.244
R7748 GND.n5447 GND.n2311 240.244
R7749 GND.n5444 GND.n2311 240.244
R7750 GND.n5444 GND.n2301 240.244
R7751 GND.n5441 GND.n2301 240.244
R7752 GND.n5441 GND.n2291 240.244
R7753 GND.n5438 GND.n2291 240.244
R7754 GND.n5438 GND.n2281 240.244
R7755 GND.n5435 GND.n2281 240.244
R7756 GND.n5435 GND.n2271 240.244
R7757 GND.n5432 GND.n2271 240.244
R7758 GND.n5432 GND.n2260 240.244
R7759 GND.n5429 GND.n2260 240.244
R7760 GND.n5429 GND.n2251 240.244
R7761 GND.n5426 GND.n2251 240.244
R7762 GND.n5426 GND.n2241 240.244
R7763 GND.n5423 GND.n2241 240.244
R7764 GND.n5423 GND.n1741 240.244
R7765 GND.n3133 GND.n3132 240.244
R7766 GND.n3097 GND.n3096 240.244
R7767 GND.n3100 GND.n3099 240.244
R7768 GND.n3105 GND.n3104 240.244
R7769 GND.n3117 GND.n3115 240.244
R7770 GND.n3052 GND.n3042 240.244
R7771 GND.n3200 GND.n3042 240.244
R7772 GND.n3200 GND.n3043 240.244
R7773 GND.n3043 GND.n3032 240.244
R7774 GND.n3191 GND.n3032 240.244
R7775 GND.n3191 GND.n3013 240.244
R7776 GND.n3332 GND.n3013 240.244
R7777 GND.n3332 GND.n3014 240.244
R7778 GND.n3014 GND.n3005 240.244
R7779 GND.n3005 GND.n2993 240.244
R7780 GND.n3349 GND.n2993 240.244
R7781 GND.n3349 GND.n2994 240.244
R7782 GND.n2994 GND.n2984 240.244
R7783 GND.n2984 GND.n2972 240.244
R7784 GND.n3366 GND.n2972 240.244
R7785 GND.n3366 GND.n2973 240.244
R7786 GND.n2973 GND.n2963 240.244
R7787 GND.n2963 GND.n2951 240.244
R7788 GND.n3383 GND.n2951 240.244
R7789 GND.n3383 GND.n2952 240.244
R7790 GND.n2952 GND.n2941 240.244
R7791 GND.n2941 GND.n2930 240.244
R7792 GND.n3400 GND.n2930 240.244
R7793 GND.n3400 GND.n2931 240.244
R7794 GND.n2931 GND.n2921 240.244
R7795 GND.n2921 GND.n2909 240.244
R7796 GND.n3417 GND.n2909 240.244
R7797 GND.n3417 GND.n2910 240.244
R7798 GND.n2910 GND.n2900 240.244
R7799 GND.n2900 GND.n2888 240.244
R7800 GND.n3434 GND.n2888 240.244
R7801 GND.n3434 GND.n2889 240.244
R7802 GND.n2889 GND.n2879 240.244
R7803 GND.n2879 GND.n2867 240.244
R7804 GND.n3451 GND.n2867 240.244
R7805 GND.n3451 GND.n2868 240.244
R7806 GND.n2868 GND.n2858 240.244
R7807 GND.n2858 GND.n2846 240.244
R7808 GND.n3468 GND.n2846 240.244
R7809 GND.n3468 GND.n2847 240.244
R7810 GND.n2847 GND.n2837 240.244
R7811 GND.n2837 GND.n2827 240.244
R7812 GND.n3491 GND.n2827 240.244
R7813 GND.n3491 GND.n2828 240.244
R7814 GND.n2828 GND.n2781 240.244
R7815 GND.n5035 GND.n2781 240.244
R7816 GND.n5036 GND.n5035 240.244
R7817 GND.n5036 GND.n2773 240.244
R7818 GND.n5039 GND.n2773 240.244
R7819 GND.n5039 GND.n2764 240.244
R7820 GND.n5041 GND.n2764 240.244
R7821 GND.n5041 GND.n2542 240.244
R7822 GND.n2755 GND.n2542 240.244
R7823 GND.n2756 GND.n2755 240.244
R7824 GND.n2756 GND.n2529 240.244
R7825 GND.n2745 GND.n2529 240.244
R7826 GND.n2746 GND.n2745 240.244
R7827 GND.n2749 GND.n2746 240.244
R7828 GND.n2749 GND.n2748 240.244
R7829 GND.n2748 GND.n2733 240.244
R7830 GND.n2733 GND.n2732 240.244
R7831 GND.n2732 GND.n2720 240.244
R7832 GND.n2720 GND.n2576 240.244
R7833 GND.n5183 GND.n2576 240.244
R7834 GND.n5183 GND.n2505 240.244
R7835 GND.n5230 GND.n2505 240.244
R7836 GND.n5231 GND.n5230 240.244
R7837 GND.n5231 GND.n2497 240.244
R7838 GND.n2497 GND.n2485 240.244
R7839 GND.n5250 GND.n2485 240.244
R7840 GND.n5251 GND.n5250 240.244
R7841 GND.n5251 GND.n2477 240.244
R7842 GND.n2477 GND.n2465 240.244
R7843 GND.n5270 GND.n2465 240.244
R7844 GND.n5271 GND.n5270 240.244
R7845 GND.n5271 GND.n2456 240.244
R7846 GND.n2456 GND.n2445 240.244
R7847 GND.n5290 GND.n2445 240.244
R7848 GND.n5291 GND.n5290 240.244
R7849 GND.n5291 GND.n2437 240.244
R7850 GND.n2437 GND.n2425 240.244
R7851 GND.n5310 GND.n2425 240.244
R7852 GND.n5311 GND.n5310 240.244
R7853 GND.n5311 GND.n2417 240.244
R7854 GND.n2417 GND.n2405 240.244
R7855 GND.n5330 GND.n2405 240.244
R7856 GND.n5331 GND.n5330 240.244
R7857 GND.n5331 GND.n2396 240.244
R7858 GND.n2396 GND.n2385 240.244
R7859 GND.n5350 GND.n2385 240.244
R7860 GND.n5351 GND.n5350 240.244
R7861 GND.n5351 GND.n2377 240.244
R7862 GND.n2377 GND.n2365 240.244
R7863 GND.n5370 GND.n2365 240.244
R7864 GND.n5371 GND.n5370 240.244
R7865 GND.n5371 GND.n2357 240.244
R7866 GND.n5374 GND.n2357 240.244
R7867 GND.n5374 GND.n2347 240.244
R7868 GND.n2347 GND.n2337 240.244
R7869 GND.n5456 GND.n2337 240.244
R7870 GND.n5456 GND.n2329 240.244
R7871 GND.n2329 GND.n2318 240.244
R7872 GND.n5475 GND.n2318 240.244
R7873 GND.n5476 GND.n5475 240.244
R7874 GND.n5476 GND.n2310 240.244
R7875 GND.n2310 GND.n2298 240.244
R7876 GND.n5495 GND.n2298 240.244
R7877 GND.n5496 GND.n5495 240.244
R7878 GND.n5496 GND.n2290 240.244
R7879 GND.n2290 GND.n2278 240.244
R7880 GND.n5515 GND.n2278 240.244
R7881 GND.n5516 GND.n5515 240.244
R7882 GND.n5516 GND.n2269 240.244
R7883 GND.n2269 GND.n2258 240.244
R7884 GND.n5535 GND.n2258 240.244
R7885 GND.n5536 GND.n5535 240.244
R7886 GND.n5536 GND.n2250 240.244
R7887 GND.n5539 GND.n2250 240.244
R7888 GND.n5539 GND.n2240 240.244
R7889 GND.n5541 GND.n2240 240.244
R7890 GND.n5541 GND.n1739 240.244
R7891 GND.n1343 GND.n1342 240.244
R7892 GND.n1382 GND.n1381 240.244
R7893 GND.n1385 GND.n1384 240.244
R7894 GND.n1390 GND.n1389 240.244
R7895 GND.n1393 GND.n1392 240.244
R7896 GND.n1398 GND.n1397 240.244
R7897 GND.n1401 GND.n1400 240.244
R7898 GND.n1406 GND.n1405 240.244
R7899 GND.n1411 GND.n1410 240.244
R7900 GND.n6277 GND.n1415 240.244
R7901 GND.n1684 GND.n1674 240.244
R7902 GND.n5829 GND.n1674 240.244
R7903 GND.n5829 GND.n1669 240.244
R7904 GND.n5837 GND.n1669 240.244
R7905 GND.n5837 GND.n1657 240.244
R7906 GND.n1657 GND.n1647 240.244
R7907 GND.n5862 GND.n1647 240.244
R7908 GND.n5862 GND.n1637 240.244
R7909 GND.n1637 GND.n1628 240.244
R7910 GND.n5877 GND.n1628 240.244
R7911 GND.n5877 GND.n1620 240.244
R7912 GND.n1620 GND.n1595 240.244
R7913 GND.n1595 GND.n1586 240.244
R7914 GND.n1586 GND.n1574 240.244
R7915 GND.n5948 GND.n1574 240.244
R7916 GND.n5949 GND.n5948 240.244
R7917 GND.n5950 GND.n5949 240.244
R7918 GND.n5950 GND.n1554 240.244
R7919 GND.n5975 GND.n1554 240.244
R7920 GND.n5975 GND.n1547 240.244
R7921 GND.n1547 GND.n1543 240.244
R7922 GND.n1543 GND.n1536 240.244
R7923 GND.n5955 GND.n1536 240.244
R7924 GND.n5955 GND.n1526 240.244
R7925 GND.n5958 GND.n1526 240.244
R7926 GND.n5959 GND.n5958 240.244
R7927 GND.n5959 GND.n1503 240.244
R7928 GND.n1503 GND.n1495 240.244
R7929 GND.n6106 GND.n1495 240.244
R7930 GND.n6106 GND.n1484 240.244
R7931 GND.n1484 GND.n1476 240.244
R7932 GND.n6131 GND.n1476 240.244
R7933 GND.n6131 GND.n1467 240.244
R7934 GND.n6112 GND.n1467 240.244
R7935 GND.n6113 GND.n6112 240.244
R7936 GND.n6114 GND.n6113 240.244
R7937 GND.n6117 GND.n6114 240.244
R7938 GND.n6118 GND.n6117 240.244
R7939 GND.n6118 GND.n1429 240.244
R7940 GND.n1429 GND.n1419 240.244
R7941 GND.n6269 GND.n1419 240.244
R7942 GND.n6269 GND.n1420 240.244
R7943 GND.n1420 GND.n1332 240.244
R7944 GND.n6276 GND.n1332 240.244
R7945 GND.n5760 GND.n1721 240.244
R7946 GND.n5698 GND.n1721 240.244
R7947 GND.n5700 GND.n5699 240.244
R7948 GND.n5704 GND.n5703 240.244
R7949 GND.n5706 GND.n5705 240.244
R7950 GND.n5710 GND.n5709 240.244
R7951 GND.n5712 GND.n5711 240.244
R7952 GND.n5716 GND.n5715 240.244
R7953 GND.n5722 GND.n5717 240.244
R7954 GND.n5724 GND.n5723 240.244
R7955 GND.n5820 GND.n1677 240.244
R7956 GND.n5827 GND.n1677 240.244
R7957 GND.n5827 GND.n1678 240.244
R7958 GND.n1678 GND.n1654 240.244
R7959 GND.n5854 GND.n1654 240.244
R7960 GND.n5854 GND.n1650 240.244
R7961 GND.n5860 GND.n1650 240.244
R7962 GND.n5860 GND.n1626 240.244
R7963 GND.n5898 GND.n1626 240.244
R7964 GND.n5898 GND.n1622 240.244
R7965 GND.n5904 GND.n1622 240.244
R7966 GND.n5904 GND.n1584 240.244
R7967 GND.n5939 GND.n1584 240.244
R7968 GND.n5939 GND.n1578 240.244
R7969 GND.n5946 GND.n1578 240.244
R7970 GND.n5946 GND.n1579 240.244
R7971 GND.n1579 GND.n1552 240.244
R7972 GND.n6007 GND.n1552 240.244
R7973 GND.n6007 GND.n1548 240.244
R7974 GND.n6013 GND.n1548 240.244
R7975 GND.n6013 GND.n1533 240.244
R7976 GND.n6059 GND.n1533 240.244
R7977 GND.n6059 GND.n1527 240.244
R7978 GND.n6066 GND.n1527 240.244
R7979 GND.n6066 GND.n1528 240.244
R7980 GND.n1528 GND.n1501 240.244
R7981 GND.n6098 GND.n1501 240.244
R7982 GND.n6098 GND.n1497 240.244
R7983 GND.n6104 GND.n1497 240.244
R7984 GND.n6104 GND.n1474 240.244
R7985 GND.n6152 GND.n1474 240.244
R7986 GND.n6152 GND.n1468 240.244
R7987 GND.n6168 GND.n1468 240.244
R7988 GND.n6168 GND.n1469 240.244
R7989 GND.n6157 GND.n1469 240.244
R7990 GND.n6158 GND.n6157 240.244
R7991 GND.n6159 GND.n6158 240.244
R7992 GND.n6159 GND.n1426 240.244
R7993 GND.n6261 GND.n1426 240.244
R7994 GND.n6261 GND.n1422 240.244
R7995 GND.n6267 GND.n1422 240.244
R7996 GND.n6267 GND.n1334 240.244
R7997 GND.n6315 GND.n1334 240.244
R7998 GND.n6315 GND.n1335 240.244
R7999 GND.n1819 GND.t48 230.173
R8000 GND.n6532 GND.t54 230.173
R8001 GND.n1817 GND.t15 230.173
R8002 GND.n6622 GND.t23 230.173
R8003 GND.n1812 GND.n1811 228.118
R8004 GND.n1176 GND.n1175 228.118
R8005 GND.n2227 GND.t27 225.165
R8006 GND.n5606 GND.t63 225.165
R8007 GND.n1756 GND.t8 225.165
R8008 GND.n6670 GND.t60 225.165
R8009 GND.n6682 GND.t51 225.165
R8010 GND.n561 GND.t30 225.165
R8011 GND.n542 GND.t66 225.165
R8012 GND.n580 GND.t19 225.165
R8013 GND.n1363 GND.t44 225.165
R8014 GND.n3066 GND.t33 225.165
R8015 GND.n3086 GND.t57 225.165
R8016 GND.n3118 GND.t72 225.165
R8017 GND.n6668 GND.n943 199.319
R8018 GND.n6668 GND.n944 199.319
R8019 GND.n5586 GND.n5585 199.319
R8020 GND.n86 GND.n85 185
R8021 GND.n84 GND.n83 185
R8022 GND.n79 GND.n78 185
R8023 GND.n107 GND.n106 185
R8024 GND.n105 GND.n104 185
R8025 GND.n100 GND.n99 185
R8026 GND.n48 GND.n47 185
R8027 GND.n46 GND.n45 185
R8028 GND.n41 GND.n40 185
R8029 GND.n69 GND.n68 185
R8030 GND.n67 GND.n66 185
R8031 GND.n62 GND.n61 185
R8032 GND.n11 GND.n10 185
R8033 GND.n9 GND.n8 185
R8034 GND.n4 GND.n3 185
R8035 GND.n32 GND.n31 185
R8036 GND.n30 GND.n29 185
R8037 GND.n25 GND.n24 185
R8038 GND.n221 GND.n220 185
R8039 GND.n219 GND.n218 185
R8040 GND.n214 GND.n213 185
R8041 GND.n200 GND.n199 185
R8042 GND.n198 GND.n197 185
R8043 GND.n193 GND.n192 185
R8044 GND.n183 GND.n182 185
R8045 GND.n181 GND.n180 185
R8046 GND.n176 GND.n175 185
R8047 GND.n162 GND.n161 185
R8048 GND.n160 GND.n159 185
R8049 GND.n155 GND.n154 185
R8050 GND.n146 GND.n145 185
R8051 GND.n144 GND.n143 185
R8052 GND.n139 GND.n138 185
R8053 GND.n125 GND.n124 185
R8054 GND.n123 GND.n122 185
R8055 GND.n118 GND.n117 185
R8056 GND.n6663 GND.n1174 163.367
R8057 GND.n6659 GND.n6658 163.367
R8058 GND.n6655 GND.n6654 163.367
R8059 GND.n6651 GND.n6650 163.367
R8060 GND.n6647 GND.n6646 163.367
R8061 GND.n6643 GND.n6642 163.367
R8062 GND.n6639 GND.n6638 163.367
R8063 GND.n6635 GND.n6634 163.367
R8064 GND.n6631 GND.n6630 163.367
R8065 GND.n6626 GND.n6625 163.367
R8066 GND.n6666 GND.n1150 163.367
R8067 GND.n6536 GND.n6535 163.367
R8068 GND.n6540 GND.n6539 163.367
R8069 GND.n6544 GND.n6543 163.367
R8070 GND.n6548 GND.n6547 163.367
R8071 GND.n6552 GND.n6551 163.367
R8072 GND.n6556 GND.n6555 163.367
R8073 GND.n6560 GND.n6559 163.367
R8074 GND.n6564 GND.n6563 163.367
R8075 GND.n6568 GND.n6567 163.367
R8076 GND.n6572 GND.n6571 163.367
R8077 GND.n2183 GND.n1823 163.367
R8078 GND.n1981 GND.n1823 163.367
R8079 GND.n1982 GND.n1981 163.367
R8080 GND.n1982 GND.n1833 163.367
R8081 GND.n1985 GND.n1833 163.367
R8082 GND.n1985 GND.n1841 163.367
R8083 GND.n1989 GND.n1841 163.367
R8084 GND.n1994 GND.n1989 163.367
R8085 GND.n1995 GND.n1994 163.367
R8086 GND.n1995 GND.n1851 163.367
R8087 GND.n1998 GND.n1851 163.367
R8088 GND.n1998 GND.n1859 163.367
R8089 GND.n2002 GND.n1859 163.367
R8090 GND.n2007 GND.n2002 163.367
R8091 GND.n2008 GND.n2007 163.367
R8092 GND.n2008 GND.n1869 163.367
R8093 GND.n2011 GND.n1869 163.367
R8094 GND.n2011 GND.n1877 163.367
R8095 GND.n2015 GND.n1877 163.367
R8096 GND.n2016 GND.n2015 163.367
R8097 GND.n2016 GND.n1888 163.367
R8098 GND.n2019 GND.n1888 163.367
R8099 GND.n2019 GND.n1896 163.367
R8100 GND.n2023 GND.n1896 163.367
R8101 GND.n2028 GND.n2023 163.367
R8102 GND.n2029 GND.n2028 163.367
R8103 GND.n2029 GND.n1906 163.367
R8104 GND.n2032 GND.n1906 163.367
R8105 GND.n2032 GND.n1914 163.367
R8106 GND.n2036 GND.n1914 163.367
R8107 GND.n2041 GND.n2036 163.367
R8108 GND.n2042 GND.n2041 163.367
R8109 GND.n2042 GND.n1924 163.367
R8110 GND.n2045 GND.n1924 163.367
R8111 GND.n2045 GND.n1932 163.367
R8112 GND.n2049 GND.n1932 163.367
R8113 GND.n2054 GND.n2049 163.367
R8114 GND.n2055 GND.n2054 163.367
R8115 GND.n2055 GND.n1942 163.367
R8116 GND.n2058 GND.n1942 163.367
R8117 GND.n2058 GND.n1950 163.367
R8118 GND.n2062 GND.n1950 163.367
R8119 GND.n2069 GND.n2062 163.367
R8120 GND.n2069 GND.n1967 163.367
R8121 GND.n2075 GND.n1967 163.367
R8122 GND.n2075 GND.n1711 163.367
R8123 GND.n1711 GND.n1704 163.367
R8124 GND.n5771 GND.n1704 163.367
R8125 GND.n5772 GND.n5771 163.367
R8126 GND.n5772 GND.n1685 163.367
R8127 GND.n5780 GND.n1685 163.367
R8128 GND.n5780 GND.n1702 163.367
R8129 GND.n5776 GND.n1702 163.367
R8130 GND.n5776 GND.n1695 163.367
R8131 GND.n1695 GND.n1667 163.367
R8132 GND.n5840 GND.n1667 163.367
R8133 GND.n5840 GND.n1656 163.367
R8134 GND.n1664 GND.n1656 163.367
R8135 GND.n5846 GND.n1664 163.367
R8136 GND.n5846 GND.n1665 163.367
R8137 GND.n1665 GND.n1636 163.367
R8138 GND.n5884 GND.n1636 163.367
R8139 GND.n5884 GND.n1629 163.367
R8140 GND.n5880 GND.n1629 163.367
R8141 GND.n5880 GND.n1642 163.367
R8142 GND.n1642 GND.n1641 163.367
R8143 GND.n1641 GND.n1594 163.367
R8144 GND.n5923 GND.n1594 163.367
R8145 GND.n5923 GND.n1587 163.367
R8146 GND.n5919 GND.n1587 163.367
R8147 GND.n5919 GND.n1612 163.367
R8148 GND.n1612 GND.n1611 163.367
R8149 GND.n1611 GND.n1599 163.367
R8150 GND.n1599 GND.n1563 163.367
R8151 GND.n1606 GND.n1563 163.367
R8152 GND.n1606 GND.n1603 163.367
R8153 GND.n1603 GND.n1602 163.367
R8154 GND.n1602 GND.n1545 163.367
R8155 GND.n6016 GND.n1545 163.367
R8156 GND.n6016 GND.n1542 163.367
R8157 GND.n6049 GND.n1542 163.367
R8158 GND.n6049 GND.n1535 163.367
R8159 GND.n6045 GND.n1535 163.367
R8160 GND.n6045 GND.n1525 163.367
R8161 GND.n6041 GND.n1525 163.367
R8162 GND.n6041 GND.n1519 163.367
R8163 GND.n6038 GND.n1519 163.367
R8164 GND.n6038 GND.n1511 163.367
R8165 GND.n6033 GND.n1511 163.367
R8166 GND.n6033 GND.n1504 163.367
R8167 GND.n6030 GND.n1504 163.367
R8168 GND.n6030 GND.n6027 163.367
R8169 GND.n6027 GND.n6026 163.367
R8170 GND.n6026 GND.n1485 163.367
R8171 GND.n6022 GND.n1485 163.367
R8172 GND.n6022 GND.n6021 163.367
R8173 GND.n6021 GND.n1465 163.367
R8174 GND.n6171 GND.n1465 163.367
R8175 GND.n6171 GND.n1459 163.367
R8176 GND.n6175 GND.n1459 163.367
R8177 GND.n6175 GND.n1452 163.367
R8178 GND.n6197 GND.n1452 163.367
R8179 GND.n6197 GND.n1450 163.367
R8180 GND.n6234 GND.n1450 163.367
R8181 GND.n6234 GND.n1444 163.367
R8182 GND.n6230 GND.n1444 163.367
R8183 GND.n6230 GND.n1428 163.367
R8184 GND.n6226 GND.n1428 163.367
R8185 GND.n6226 GND.n1437 163.367
R8186 GND.n6222 GND.n1437 163.367
R8187 GND.n6222 GND.n6221 163.367
R8188 GND.n6221 GND.n6211 163.367
R8189 GND.n6211 GND.n6201 163.367
R8190 GND.n6207 GND.n6201 163.367
R8191 GND.n6207 GND.n1322 163.367
R8192 GND.n6202 GND.n1322 163.367
R8193 GND.n6202 GND.n1316 163.367
R8194 GND.n6339 GND.n1316 163.367
R8195 GND.n6339 GND.n1314 163.367
R8196 GND.n6347 GND.n1314 163.367
R8197 GND.n6347 GND.n1308 163.367
R8198 GND.n6343 GND.n1308 163.367
R8199 GND.n6343 GND.n1301 163.367
R8200 GND.n1301 GND.n1293 163.367
R8201 GND.n6384 GND.n1293 163.367
R8202 GND.n6384 GND.n1291 163.367
R8203 GND.n6388 GND.n1291 163.367
R8204 GND.n6388 GND.n1284 163.367
R8205 GND.n6397 GND.n1284 163.367
R8206 GND.n6397 GND.n1281 163.367
R8207 GND.n6406 GND.n1281 163.367
R8208 GND.n6406 GND.n1282 163.367
R8209 GND.n1282 GND.n1275 163.367
R8210 GND.n6401 GND.n1275 163.367
R8211 GND.n6401 GND.n1267 163.367
R8212 GND.n1267 GND.n1259 163.367
R8213 GND.n6433 GND.n1259 163.367
R8214 GND.n6433 GND.n1256 163.367
R8215 GND.n6442 GND.n1256 163.367
R8216 GND.n6442 GND.n1257 163.367
R8217 GND.n1257 GND.n1250 163.367
R8218 GND.n6437 GND.n1250 163.367
R8219 GND.n6437 GND.n1241 163.367
R8220 GND.n1241 GND.n1234 163.367
R8221 GND.n6471 GND.n1234 163.367
R8222 GND.n6471 GND.n1231 163.367
R8223 GND.n6480 GND.n1231 163.367
R8224 GND.n6480 GND.n1232 163.367
R8225 GND.n1232 GND.n1225 163.367
R8226 GND.n6475 GND.n1225 163.367
R8227 GND.n6475 GND.n1217 163.367
R8228 GND.n1217 GND.n1209 163.367
R8229 GND.n6516 GND.n1209 163.367
R8230 GND.n6516 GND.n1207 163.367
R8231 GND.n6520 GND.n1207 163.367
R8232 GND.n6520 GND.n1200 163.367
R8233 GND.n6529 GND.n1200 163.367
R8234 GND.n6529 GND.n1197 163.367
R8235 GND.n6585 GND.n1197 163.367
R8236 GND.n6585 GND.n1198 163.367
R8237 GND.n1198 GND.n1191 163.367
R8238 GND.n6580 GND.n1191 163.367
R8239 GND.n6580 GND.n1183 163.367
R8240 GND.n6577 GND.n1183 163.367
R8241 GND.n1809 GND.n1808 163.367
R8242 GND.n5669 GND.n1808 163.367
R8243 GND.n5667 GND.n5666 163.367
R8244 GND.n5663 GND.n5662 163.367
R8245 GND.n5659 GND.n5658 163.367
R8246 GND.n5655 GND.n5654 163.367
R8247 GND.n5651 GND.n5650 163.367
R8248 GND.n5647 GND.n5646 163.367
R8249 GND.n5643 GND.n5642 163.367
R8250 GND.n5638 GND.n5637 163.367
R8251 GND.n5634 GND.n5633 163.367
R8252 GND.n2224 GND.n2223 163.367
R8253 GND.n2220 GND.n2219 163.367
R8254 GND.n2216 GND.n2215 163.367
R8255 GND.n2212 GND.n2211 163.367
R8256 GND.n2208 GND.n2207 163.367
R8257 GND.n2204 GND.n2203 163.367
R8258 GND.n2200 GND.n2199 163.367
R8259 GND.n2196 GND.n2195 163.367
R8260 GND.n2192 GND.n2191 163.367
R8261 GND.n2188 GND.n2187 163.367
R8262 GND.n1976 GND.n1810 163.367
R8263 GND.n1980 GND.n1976 163.367
R8264 GND.n1980 GND.n1835 163.367
R8265 GND.n2173 GND.n1835 163.367
R8266 GND.n2173 GND.n1836 163.367
R8267 GND.n2169 GND.n1836 163.367
R8268 GND.n2169 GND.n1839 163.367
R8269 GND.n1992 GND.n1839 163.367
R8270 GND.n1992 GND.n1852 163.367
R8271 GND.n2159 GND.n1852 163.367
R8272 GND.n2159 GND.n1853 163.367
R8273 GND.n2155 GND.n1853 163.367
R8274 GND.n2155 GND.n1856 163.367
R8275 GND.n2005 GND.n1856 163.367
R8276 GND.n2005 GND.n1871 163.367
R8277 GND.n2145 GND.n1871 163.367
R8278 GND.n2145 GND.n1872 163.367
R8279 GND.n2141 GND.n1872 163.367
R8280 GND.n2141 GND.n1875 163.367
R8281 GND.n1890 GND.n1875 163.367
R8282 GND.n2131 GND.n1890 163.367
R8283 GND.n2131 GND.n1891 163.367
R8284 GND.n2127 GND.n1891 163.367
R8285 GND.n2127 GND.n1894 163.367
R8286 GND.n2026 GND.n1894 163.367
R8287 GND.n2026 GND.n1908 163.367
R8288 GND.n2117 GND.n1908 163.367
R8289 GND.n2117 GND.n1909 163.367
R8290 GND.n2113 GND.n1909 163.367
R8291 GND.n2113 GND.n1912 163.367
R8292 GND.n2039 GND.n1912 163.367
R8293 GND.n2039 GND.n1926 163.367
R8294 GND.n2103 GND.n1926 163.367
R8295 GND.n2103 GND.n1927 163.367
R8296 GND.n2099 GND.n1927 163.367
R8297 GND.n2099 GND.n1930 163.367
R8298 GND.n2052 GND.n1930 163.367
R8299 GND.n2052 GND.n1944 163.367
R8300 GND.n2089 GND.n1944 163.367
R8301 GND.n2089 GND.n1945 163.367
R8302 GND.n2085 GND.n1945 163.367
R8303 GND.n2085 GND.n1948 163.367
R8304 GND.n2067 GND.n1948 163.367
R8305 GND.n2067 GND.n2064 163.367
R8306 GND.n2064 GND.n1709 163.367
R8307 GND.n5765 GND.n1709 163.367
R8308 GND.n5765 GND.n1707 163.367
R8309 GND.n5769 GND.n1707 163.367
R8310 GND.n5769 GND.n1687 163.367
R8311 GND.n5817 GND.n1687 163.367
R8312 GND.n5817 GND.n1688 163.367
R8313 GND.n5813 GND.n1688 163.367
R8314 GND.n5813 GND.n5812 163.367
R8315 GND.n5812 GND.n5811 163.367
R8316 GND.n5811 GND.n1691 163.367
R8317 GND.n1691 GND.n1659 163.367
R8318 GND.n5852 GND.n1659 163.367
R8319 GND.n5852 GND.n1660 163.367
R8320 GND.n5848 GND.n1660 163.367
R8321 GND.n5848 GND.n1634 163.367
R8322 GND.n5888 GND.n1634 163.367
R8323 GND.n5888 GND.n1631 163.367
R8324 GND.n5895 GND.n1631 163.367
R8325 GND.n5895 GND.n1632 163.367
R8326 GND.n5891 GND.n1632 163.367
R8327 GND.n5891 GND.n1592 163.367
R8328 GND.n5927 GND.n1592 163.367
R8329 GND.n5927 GND.n1589 163.367
R8330 GND.n5936 GND.n1589 163.367
R8331 GND.n5936 GND.n1590 163.367
R8332 GND.n5932 GND.n1590 163.367
R8333 GND.n5932 GND.n5931 163.367
R8334 GND.n5931 GND.n1565 163.367
R8335 GND.n5984 GND.n1565 163.367
R8336 GND.n5984 GND.n1566 163.367
R8337 GND.n5980 GND.n1566 163.367
R8338 GND.n5980 GND.n5979 163.367
R8339 GND.n5979 GND.n5978 163.367
R8340 GND.n5978 GND.n1540 163.367
R8341 GND.n6053 GND.n1540 163.367
R8342 GND.n6053 GND.n1538 163.367
R8343 GND.n6057 GND.n1538 163.367
R8344 GND.n6057 GND.n1523 163.367
R8345 GND.n6070 GND.n1523 163.367
R8346 GND.n6070 GND.n1521 163.367
R8347 GND.n6074 GND.n1521 163.367
R8348 GND.n6074 GND.n1509 163.367
R8349 GND.n6088 GND.n1509 163.367
R8350 GND.n6088 GND.n1506 163.367
R8351 GND.n6095 GND.n1506 163.367
R8352 GND.n6095 GND.n1507 163.367
R8353 GND.n6091 GND.n1507 163.367
R8354 GND.n6091 GND.n1487 163.367
R8355 GND.n6139 GND.n1487 163.367
R8356 GND.n6139 GND.n1488 163.367
R8357 GND.n6135 GND.n1488 163.367
R8358 GND.n6135 GND.n6134 163.367
R8359 GND.n6134 GND.n1461 163.367
R8360 GND.n6183 GND.n1461 163.367
R8361 GND.n6183 GND.n1462 163.367
R8362 GND.n6179 GND.n1462 163.367
R8363 GND.n6179 GND.n1448 163.367
R8364 GND.n6238 GND.n1448 163.367
R8365 GND.n6238 GND.n1446 163.367
R8366 GND.n6242 GND.n1446 163.367
R8367 GND.n6242 GND.n1431 163.367
R8368 GND.n6259 GND.n1431 163.367
R8369 GND.n6259 GND.n1432 163.367
R8370 GND.n6255 GND.n1432 163.367
R8371 GND.n6255 GND.n1435 163.367
R8372 GND.n6219 GND.n1435 163.367
R8373 GND.n6219 GND.n6214 163.367
R8374 GND.n6215 GND.n6214 163.367
R8375 GND.n6215 GND.n1320 163.367
R8376 GND.n6332 GND.n1320 163.367
R8377 GND.n6332 GND.n1318 163.367
R8378 GND.n6336 GND.n1318 163.367
R8379 GND.n6336 GND.n1312 163.367
R8380 GND.n6351 GND.n1312 163.367
R8381 GND.n6351 GND.n1310 163.367
R8382 GND.n6355 GND.n1310 163.367
R8383 GND.n6355 GND.n1299 163.367
R8384 GND.n6378 GND.n1299 163.367
R8385 GND.n6378 GND.n1297 163.367
R8386 GND.n6382 GND.n1297 163.367
R8387 GND.n6382 GND.n1289 163.367
R8388 GND.n6391 GND.n1289 163.367
R8389 GND.n6391 GND.n1287 163.367
R8390 GND.n6395 GND.n1287 163.367
R8391 GND.n6395 GND.n1279 163.367
R8392 GND.n6409 GND.n1279 163.367
R8393 GND.n6409 GND.n1277 163.367
R8394 GND.n6413 GND.n1277 163.367
R8395 GND.n6413 GND.n1265 163.367
R8396 GND.n6427 GND.n1265 163.367
R8397 GND.n6427 GND.n1263 163.367
R8398 GND.n6431 GND.n1263 163.367
R8399 GND.n6431 GND.n1254 163.367
R8400 GND.n6444 GND.n1254 163.367
R8401 GND.n6444 GND.n1252 163.367
R8402 GND.n6448 GND.n1252 163.367
R8403 GND.n6448 GND.n1239 163.367
R8404 GND.n6465 GND.n1239 163.367
R8405 GND.n6465 GND.n1237 163.367
R8406 GND.n6469 GND.n1237 163.367
R8407 GND.n6469 GND.n1229 163.367
R8408 GND.n6483 GND.n1229 163.367
R8409 GND.n6483 GND.n1227 163.367
R8410 GND.n6487 GND.n1227 163.367
R8411 GND.n6487 GND.n1215 163.367
R8412 GND.n6510 GND.n1215 163.367
R8413 GND.n6510 GND.n1213 163.367
R8414 GND.n6514 GND.n1213 163.367
R8415 GND.n6514 GND.n1205 163.367
R8416 GND.n6523 GND.n1205 163.367
R8417 GND.n6523 GND.n1203 163.367
R8418 GND.n6527 GND.n1203 163.367
R8419 GND.n6527 GND.n1195 163.367
R8420 GND.n6588 GND.n1195 163.367
R8421 GND.n6588 GND.n1193 163.367
R8422 GND.n6592 GND.n1193 163.367
R8423 GND.n6592 GND.n1181 163.367
R8424 GND.n6618 GND.n1181 163.367
R8425 GND.n6618 GND.n1173 163.367
R8426 GND.n1815 GND.n1814 152
R8427 GND.n1179 GND.n1178 152
R8428 GND.n80 GND.t145 150.499
R8429 GND.n101 GND.t130 150.499
R8430 GND.n42 GND.t144 150.499
R8431 GND.n63 GND.t91 150.499
R8432 GND.n5 GND.t93 150.499
R8433 GND.n26 GND.t141 150.499
R8434 GND.n215 GND.t95 150.499
R8435 GND.n194 GND.t135 150.499
R8436 GND.n177 GND.t115 150.499
R8437 GND.n156 GND.t121 150.499
R8438 GND.n140 GND.t126 150.499
R8439 GND.n119 GND.t146 150.499
R8440 GND.n1820 GND.t49 144.291
R8441 GND.n6533 GND.t56 144.291
R8442 GND.n1818 GND.t17 144.291
R8443 GND.n6623 GND.t26 144.291
R8444 GND.n6665 GND.n1149 143.351
R8445 GND.n1162 GND.n1149 143.351
R8446 GND.n5631 GND.n1795 143.351
R8447 GND.n5631 GND.n1796 143.351
R8448 GND.n3527 GND.n2782 140.306
R8449 GND.n1813 GND.t12 138.431
R8450 GND.n1177 GND.t69 138.431
R8451 GND.n2228 GND.t29 135.476
R8452 GND.n5607 GND.t65 135.476
R8453 GND.n1757 GND.t11 135.476
R8454 GND.n6671 GND.t61 135.476
R8455 GND.n6683 GND.t52 135.476
R8456 GND.n562 GND.t32 135.476
R8457 GND.n543 GND.t68 135.476
R8458 GND.n581 GND.t22 135.476
R8459 GND.n1364 GND.t46 135.476
R8460 GND.n3067 GND.t35 135.476
R8461 GND.n3087 GND.t58 135.476
R8462 GND.n3119 GND.t73 135.476
R8463 GND.n5718 GND.t40 126.853
R8464 GND.n1407 GND.t80 126.853
R8465 GND.n1814 GND.t75 126.766
R8466 GND.n1178 GND.t41 126.766
R8467 GND.n2228 GND.n2227 112.097
R8468 GND.n5607 GND.n5606 112.097
R8469 GND.n1757 GND.n1756 112.097
R8470 GND.n6671 GND.n6670 112.097
R8471 GND.n6683 GND.n6682 112.097
R8472 GND.n562 GND.n561 112.097
R8473 GND.n543 GND.n542 112.097
R8474 GND.n581 GND.n580 112.097
R8475 GND.n1364 GND.n1363 112.097
R8476 GND.n3067 GND.n3066 112.097
R8477 GND.n3087 GND.n3086 112.097
R8478 GND.n3119 GND.n3118 112.097
R8479 GND.n85 GND.n84 104.615
R8480 GND.n84 GND.n78 104.615
R8481 GND.n106 GND.n105 104.615
R8482 GND.n105 GND.n99 104.615
R8483 GND.n47 GND.n46 104.615
R8484 GND.n46 GND.n40 104.615
R8485 GND.n68 GND.n67 104.615
R8486 GND.n67 GND.n61 104.615
R8487 GND.n10 GND.n9 104.615
R8488 GND.n9 GND.n3 104.615
R8489 GND.n31 GND.n30 104.615
R8490 GND.n30 GND.n24 104.615
R8491 GND.n220 GND.n219 104.615
R8492 GND.n219 GND.n213 104.615
R8493 GND.n199 GND.n198 104.615
R8494 GND.n198 GND.n192 104.615
R8495 GND.n182 GND.n181 104.615
R8496 GND.n181 GND.n175 104.615
R8497 GND.n161 GND.n160 104.615
R8498 GND.n160 GND.n154 104.615
R8499 GND.n145 GND.n144 104.615
R8500 GND.n144 GND.n138 104.615
R8501 GND.n124 GND.n123 104.615
R8502 GND.n123 GND.n117 104.615
R8503 GND.n7462 GND.n7461 99.6594
R8504 GND.n7459 GND.n7458 99.6594
R8505 GND.n7454 GND.n536 99.6594
R8506 GND.n7452 GND.n7451 99.6594
R8507 GND.n545 GND.n544 99.6594
R8508 GND.n7443 GND.n549 99.6594
R8509 GND.n7441 GND.n7440 99.6594
R8510 GND.n7436 GND.n555 99.6594
R8511 GND.n7434 GND.n7433 99.6594
R8512 GND.n7429 GND.n564 99.6594
R8513 GND.n7427 GND.n7426 99.6594
R8514 GND.n6724 GND.n6723 99.6594
R8515 GND.n6718 GND.n941 99.6594
R8516 GND.n6715 GND.n942 99.6594
R8517 GND.n6711 GND.n943 99.6594
R8518 GND.n6706 GND.n945 99.6594
R8519 GND.n6702 GND.n946 99.6594
R8520 GND.n6698 GND.n947 99.6594
R8521 GND.n6694 GND.n948 99.6594
R8522 GND.n6690 GND.n949 99.6594
R8523 GND.n7342 GND.n7341 99.6594
R8524 GND.n7337 GND.n574 99.6594
R8525 GND.n7335 GND.n7334 99.6594
R8526 GND.n7330 GND.n583 99.6594
R8527 GND.n7328 GND.n7327 99.6594
R8528 GND.n1345 GND.n955 99.6594
R8529 GND.n1349 GND.n954 99.6594
R8530 GND.n1354 GND.n953 99.6594
R8531 GND.n1359 GND.n952 99.6594
R8532 GND.n1367 GND.n951 99.6594
R8533 GND.n5024 GND.n5023 99.6594
R8534 GND.n5018 GND.n2791 99.6594
R8535 GND.n5015 GND.n2792 99.6594
R8536 GND.n5011 GND.n2793 99.6594
R8537 GND.n5007 GND.n2794 99.6594
R8538 GND.n5003 GND.n2795 99.6594
R8539 GND.n4999 GND.n2796 99.6594
R8540 GND.n4995 GND.n2797 99.6594
R8541 GND.n4991 GND.n2798 99.6594
R8542 GND.n4987 GND.n2799 99.6594
R8543 GND.n4983 GND.n2800 99.6594
R8544 GND.n4979 GND.n2801 99.6594
R8545 GND.n4975 GND.n2802 99.6594
R8546 GND.n4971 GND.n2803 99.6594
R8547 GND.n4967 GND.n2804 99.6594
R8548 GND.n4963 GND.n2805 99.6594
R8549 GND.n4959 GND.n2806 99.6594
R8550 GND.n4955 GND.n2807 99.6594
R8551 GND.n4951 GND.n2808 99.6594
R8552 GND.n4947 GND.n2809 99.6594
R8553 GND.n4943 GND.n2810 99.6594
R8554 GND.n4939 GND.n2811 99.6594
R8555 GND.n4935 GND.n2812 99.6594
R8556 GND.n4931 GND.n2813 99.6594
R8557 GND.n4927 GND.n2814 99.6594
R8558 GND.n4923 GND.n2815 99.6594
R8559 GND.n4919 GND.n2816 99.6594
R8560 GND.n5027 GND.n5026 99.6594
R8561 GND.n5572 GND.n2234 99.6594
R8562 GND.n5576 GND.n5574 99.6594
R8563 GND.n5583 GND.n2230 99.6594
R8564 GND.n5592 GND.n5591 99.6594
R8565 GND.n5595 GND.n5594 99.6594
R8566 GND.n5600 GND.n5599 99.6594
R8567 GND.n5603 GND.n5602 99.6594
R8568 GND.n5609 GND.n5608 99.6594
R8569 GND.n5610 GND.n1736 99.6594
R8570 GND.n3177 GND.n3053 99.6594
R8571 GND.n3175 GND.n3056 99.6594
R8572 GND.n3171 GND.n3170 99.6594
R8573 GND.n3164 GND.n3061 99.6594
R8574 GND.n3163 GND.n3162 99.6594
R8575 GND.n3156 GND.n3069 99.6594
R8576 GND.n3155 GND.n3154 99.6594
R8577 GND.n3148 GND.n3075 99.6594
R8578 GND.n3147 GND.n3146 99.6594
R8579 GND.n3084 GND.n3081 99.6594
R8580 GND.n1772 GND.n1755 99.6594
R8581 GND.n1768 GND.n1754 99.6594
R8582 GND.n1764 GND.n1753 99.6594
R8583 GND.n1760 GND.n1752 99.6594
R8584 GND.n1751 GND.n1750 99.6594
R8585 GND.n3135 GND.n3134 99.6594
R8586 GND.n3132 GND.n3093 99.6594
R8587 GND.n3098 GND.n3097 99.6594
R8588 GND.n3103 GND.n3100 99.6594
R8589 GND.n3116 GND.n3105 99.6594
R8590 GND.n3134 GND.n3133 99.6594
R8591 GND.n3096 GND.n3093 99.6594
R8592 GND.n3099 GND.n3098 99.6594
R8593 GND.n3104 GND.n3103 99.6594
R8594 GND.n3117 GND.n3116 99.6594
R8595 GND.n3178 GND.n3177 99.6594
R8596 GND.n3172 GND.n3056 99.6594
R8597 GND.n3170 GND.n3169 99.6594
R8598 GND.n3165 GND.n3164 99.6594
R8599 GND.n3162 GND.n3161 99.6594
R8600 GND.n3157 GND.n3156 99.6594
R8601 GND.n3154 GND.n3153 99.6594
R8602 GND.n3149 GND.n3148 99.6594
R8603 GND.n3146 GND.n3145 99.6594
R8604 GND.n3085 GND.n3084 99.6594
R8605 GND.n5024 GND.n3522 99.6594
R8606 GND.n5016 GND.n2791 99.6594
R8607 GND.n5012 GND.n2792 99.6594
R8608 GND.n5008 GND.n2793 99.6594
R8609 GND.n5004 GND.n2794 99.6594
R8610 GND.n5000 GND.n2795 99.6594
R8611 GND.n4996 GND.n2796 99.6594
R8612 GND.n4992 GND.n2797 99.6594
R8613 GND.n4988 GND.n2798 99.6594
R8614 GND.n4984 GND.n2799 99.6594
R8615 GND.n4980 GND.n2800 99.6594
R8616 GND.n4976 GND.n2801 99.6594
R8617 GND.n4972 GND.n2802 99.6594
R8618 GND.n4968 GND.n2803 99.6594
R8619 GND.n4964 GND.n2804 99.6594
R8620 GND.n4960 GND.n2805 99.6594
R8621 GND.n4956 GND.n2806 99.6594
R8622 GND.n4952 GND.n2807 99.6594
R8623 GND.n4948 GND.n2808 99.6594
R8624 GND.n4944 GND.n2809 99.6594
R8625 GND.n4940 GND.n2810 99.6594
R8626 GND.n4936 GND.n2811 99.6594
R8627 GND.n4932 GND.n2812 99.6594
R8628 GND.n4928 GND.n2813 99.6594
R8629 GND.n4924 GND.n2814 99.6594
R8630 GND.n4920 GND.n2815 99.6594
R8631 GND.n2816 GND.n2789 99.6594
R8632 GND.n5026 GND.n2786 99.6594
R8633 GND.n1759 GND.n1751 99.6594
R8634 GND.n1763 GND.n1752 99.6594
R8635 GND.n1767 GND.n1753 99.6594
R8636 GND.n1771 GND.n1754 99.6594
R8637 GND.n1775 GND.n1755 99.6594
R8638 GND.n1348 GND.n955 99.6594
R8639 GND.n1353 GND.n954 99.6594
R8640 GND.n1358 GND.n953 99.6594
R8641 GND.n1366 GND.n952 99.6594
R8642 GND.n1362 GND.n951 99.6594
R8643 GND.n7329 GND.n7328 99.6594
R8644 GND.n583 GND.n575 99.6594
R8645 GND.n7336 GND.n7335 99.6594
R8646 GND.n574 GND.n569 99.6594
R8647 GND.n7343 GND.n7342 99.6594
R8648 GND.n5611 GND.n5610 99.6594
R8649 GND.n5608 GND.n5604 99.6594
R8650 GND.n5602 GND.n5601 99.6594
R8651 GND.n5599 GND.n5596 99.6594
R8652 GND.n5594 GND.n5593 99.6594
R8653 GND.n5591 GND.n5588 99.6594
R8654 GND.n5587 GND.n5586 99.6594
R8655 GND.n5585 GND.n5584 99.6594
R8656 GND.n5575 GND.n2230 99.6594
R8657 GND.n5574 GND.n5573 99.6594
R8658 GND.n5565 GND.n2234 99.6594
R8659 GND.n6724 GND.n957 99.6594
R8660 GND.n6716 GND.n941 99.6594
R8661 GND.n6712 GND.n942 99.6594
R8662 GND.n6707 GND.n944 99.6594
R8663 GND.n6703 GND.n945 99.6594
R8664 GND.n6699 GND.n946 99.6594
R8665 GND.n6695 GND.n947 99.6594
R8666 GND.n6691 GND.n948 99.6594
R8667 GND.n6681 GND.n949 99.6594
R8668 GND.n7428 GND.n7427 99.6594
R8669 GND.n564 GND.n556 99.6594
R8670 GND.n7435 GND.n7434 99.6594
R8671 GND.n555 GND.n550 99.6594
R8672 GND.n7442 GND.n7441 99.6594
R8673 GND.n549 GND.n548 99.6594
R8674 GND.n544 GND.n537 99.6594
R8675 GND.n7453 GND.n7452 99.6594
R8676 GND.n536 GND.n530 99.6594
R8677 GND.n7460 GND.n7459 99.6594
R8678 GND.n7463 GND.n7462 99.6594
R8679 GND.n1341 GND.n1340 99.6594
R8680 GND.n1380 GND.n1343 99.6594
R8681 GND.n1383 GND.n1382 99.6594
R8682 GND.n1388 GND.n1385 99.6594
R8683 GND.n1391 GND.n1390 99.6594
R8684 GND.n1396 GND.n1393 99.6594
R8685 GND.n1399 GND.n1398 99.6594
R8686 GND.n1404 GND.n1401 99.6594
R8687 GND.n1409 GND.n1406 99.6594
R8688 GND.n1414 GND.n1411 99.6594
R8689 GND.n1415 GND.n1414 99.6594
R8690 GND.n1410 GND.n1409 99.6594
R8691 GND.n1405 GND.n1404 99.6594
R8692 GND.n1400 GND.n1399 99.6594
R8693 GND.n1397 GND.n1396 99.6594
R8694 GND.n1392 GND.n1391 99.6594
R8695 GND.n1389 GND.n1388 99.6594
R8696 GND.n1384 GND.n1383 99.6594
R8697 GND.n1381 GND.n1380 99.6594
R8698 GND.n1342 GND.n1341 99.6594
R8699 GND.n5761 GND.n1682 99.6594
R8700 GND.n5698 GND.n1712 99.6594
R8701 GND.n5700 GND.n1713 99.6594
R8702 GND.n5704 GND.n1714 99.6594
R8703 GND.n5706 GND.n1715 99.6594
R8704 GND.n5710 GND.n1716 99.6594
R8705 GND.n5712 GND.n1717 99.6594
R8706 GND.n5716 GND.n1718 99.6594
R8707 GND.n5722 GND.n1719 99.6594
R8708 GND.n5724 GND.n1720 99.6594
R8709 GND.n5761 GND.n5760 99.6594
R8710 GND.n5699 GND.n1712 99.6594
R8711 GND.n5703 GND.n1713 99.6594
R8712 GND.n5705 GND.n1714 99.6594
R8713 GND.n5709 GND.n1715 99.6594
R8714 GND.n5711 GND.n1716 99.6594
R8715 GND.n5715 GND.n1717 99.6594
R8716 GND.n5717 GND.n1718 99.6594
R8717 GND.n5723 GND.n1719 99.6594
R8718 GND.n5725 GND.n1720 99.6594
R8719 GND.n1820 GND.n1819 97.552
R8720 GND.n6533 GND.n6532 97.552
R8721 GND.n1818 GND.n1817 97.552
R8722 GND.n6623 GND.n6622 97.552
R8723 GND.t110 GND.n2782 89.8748
R8724 GND.n5719 GND.t39 73.9079
R8725 GND.n1408 GND.t81 73.9079
R8726 GND.n1813 GND.n1812 73.571
R8727 GND.n1177 GND.n1176 73.571
R8728 GND.n4305 GND.n4304 72.5001
R8729 GND.n4304 GND.n4079 72.5001
R8730 GND.n4296 GND.n4079 72.5001
R8731 GND.n4296 GND.n4295 72.5001
R8732 GND.n4295 GND.n4294 72.5001
R8733 GND.n4294 GND.n4087 72.5001
R8734 GND.n4288 GND.n4087 72.5001
R8735 GND.n4288 GND.n4287 72.5001
R8736 GND.n4287 GND.n4286 72.5001
R8737 GND.n4286 GND.n4094 72.5001
R8738 GND.n4280 GND.n4094 72.5001
R8739 GND.n4280 GND.n4279 72.5001
R8740 GND.n4279 GND.n4278 72.5001
R8741 GND.n4278 GND.n4102 72.5001
R8742 GND.n4272 GND.n4102 72.5001
R8743 GND.n4272 GND.n4271 72.5001
R8744 GND.n4271 GND.n4270 72.5001
R8745 GND.n4270 GND.n4110 72.5001
R8746 GND.n4264 GND.n4110 72.5001
R8747 GND.n4264 GND.n4263 72.5001
R8748 GND.n4263 GND.n4262 72.5001
R8749 GND.n4262 GND.n4118 72.5001
R8750 GND.n4256 GND.n4118 72.5001
R8751 GND.n4256 GND.n4255 72.5001
R8752 GND.n4255 GND.n4254 72.5001
R8753 GND.n4254 GND.n4126 72.5001
R8754 GND.n4248 GND.n4126 72.5001
R8755 GND.n4248 GND.n4247 72.5001
R8756 GND.n4247 GND.n4246 72.5001
R8757 GND.n4246 GND.n4134 72.5001
R8758 GND.n4240 GND.n4134 72.5001
R8759 GND.n4240 GND.n4239 72.5001
R8760 GND.n4239 GND.n4238 72.5001
R8761 GND.n4238 GND.n4142 72.5001
R8762 GND.n4232 GND.n4142 72.5001
R8763 GND.n4232 GND.n4231 72.5001
R8764 GND.n4231 GND.n4230 72.5001
R8765 GND.n4230 GND.n4150 72.5001
R8766 GND.n4224 GND.n4150 72.5001
R8767 GND.n4224 GND.n4223 72.5001
R8768 GND.n4223 GND.n4222 72.5001
R8769 GND.n4222 GND.n4158 72.5001
R8770 GND.n4216 GND.n4158 72.5001
R8771 GND.n4216 GND.n4215 72.5001
R8772 GND.n4215 GND.n4214 72.5001
R8773 GND.n4214 GND.n4166 72.5001
R8774 GND.n4208 GND.n4166 72.5001
R8775 GND.n4208 GND.n4207 72.5001
R8776 GND.n4207 GND.n4206 72.5001
R8777 GND.n4206 GND.n4174 72.5001
R8778 GND.n4200 GND.n4174 72.5001
R8779 GND.n4200 GND.n4199 72.5001
R8780 GND.n4199 GND.n4198 72.5001
R8781 GND.n4198 GND.n4182 72.5001
R8782 GND.n4192 GND.n4182 72.5001
R8783 GND.n6659 GND.n1172 71.676
R8784 GND.n6655 GND.n1171 71.676
R8785 GND.n6651 GND.n1170 71.676
R8786 GND.n6647 GND.n1169 71.676
R8787 GND.n6643 GND.n1168 71.676
R8788 GND.n6639 GND.n1167 71.676
R8789 GND.n6635 GND.n1166 71.676
R8790 GND.n6631 GND.n1165 71.676
R8791 GND.n6626 GND.n1164 71.676
R8792 GND.n1163 GND.n1150 71.676
R8793 GND.n6535 GND.n1162 71.676
R8794 GND.n6539 GND.n1161 71.676
R8795 GND.n6543 GND.n1160 71.676
R8796 GND.n6547 GND.n1159 71.676
R8797 GND.n6551 GND.n1158 71.676
R8798 GND.n6555 GND.n1157 71.676
R8799 GND.n6559 GND.n1156 71.676
R8800 GND.n6563 GND.n1155 71.676
R8801 GND.n6567 GND.n1154 71.676
R8802 GND.n6571 GND.n1153 71.676
R8803 GND.n6575 GND.n1152 71.676
R8804 GND.n5675 GND.n5674 71.676
R8805 GND.n5669 GND.n1786 71.676
R8806 GND.n5666 GND.n1787 71.676
R8807 GND.n5662 GND.n1788 71.676
R8808 GND.n5658 GND.n1789 71.676
R8809 GND.n5654 GND.n1790 71.676
R8810 GND.n5650 GND.n1791 71.676
R8811 GND.n5646 GND.n1792 71.676
R8812 GND.n5642 GND.n1793 71.676
R8813 GND.n5637 GND.n1794 71.676
R8814 GND.n5633 GND.n1795 71.676
R8815 GND.n2223 GND.n1797 71.676
R8816 GND.n2219 GND.n1798 71.676
R8817 GND.n2215 GND.n1799 71.676
R8818 GND.n2211 GND.n1800 71.676
R8819 GND.n2207 GND.n1801 71.676
R8820 GND.n2203 GND.n1802 71.676
R8821 GND.n2199 GND.n1803 71.676
R8822 GND.n2195 GND.n1804 71.676
R8823 GND.n2191 GND.n1805 71.676
R8824 GND.n2187 GND.n1806 71.676
R8825 GND.n5675 GND.n1809 71.676
R8826 GND.n5667 GND.n1786 71.676
R8827 GND.n5663 GND.n1787 71.676
R8828 GND.n5659 GND.n1788 71.676
R8829 GND.n5655 GND.n1789 71.676
R8830 GND.n5651 GND.n1790 71.676
R8831 GND.n5647 GND.n1791 71.676
R8832 GND.n5643 GND.n1792 71.676
R8833 GND.n5638 GND.n1793 71.676
R8834 GND.n5634 GND.n1794 71.676
R8835 GND.n2224 GND.n1796 71.676
R8836 GND.n2220 GND.n1797 71.676
R8837 GND.n2216 GND.n1798 71.676
R8838 GND.n2212 GND.n1799 71.676
R8839 GND.n2208 GND.n1800 71.676
R8840 GND.n2204 GND.n1801 71.676
R8841 GND.n2200 GND.n1802 71.676
R8842 GND.n2196 GND.n1803 71.676
R8843 GND.n2192 GND.n1804 71.676
R8844 GND.n2188 GND.n1805 71.676
R8845 GND.n2184 GND.n1806 71.676
R8846 GND.n6572 GND.n1152 71.676
R8847 GND.n6568 GND.n1153 71.676
R8848 GND.n6564 GND.n1154 71.676
R8849 GND.n6560 GND.n1155 71.676
R8850 GND.n6556 GND.n1156 71.676
R8851 GND.n6552 GND.n1157 71.676
R8852 GND.n6548 GND.n1158 71.676
R8853 GND.n6544 GND.n1159 71.676
R8854 GND.n6540 GND.n1160 71.676
R8855 GND.n6536 GND.n1161 71.676
R8856 GND.n6666 GND.n6665 71.676
R8857 GND.n6625 GND.n1163 71.676
R8858 GND.n6630 GND.n1164 71.676
R8859 GND.n6634 GND.n1165 71.676
R8860 GND.n6638 GND.n1166 71.676
R8861 GND.n6642 GND.n1167 71.676
R8862 GND.n6646 GND.n1168 71.676
R8863 GND.n6650 GND.n1169 71.676
R8864 GND.n6654 GND.n1170 71.676
R8865 GND.n6658 GND.n1171 71.676
R8866 GND.n1174 GND.n1172 71.676
R8867 GND.n528 GND.n522 63.7575
R8868 GND.n1816 GND.n1815 63.641
R8869 GND.n91 GND.n90 60.0588
R8870 GND.n93 GND.n92 60.0588
R8871 GND.n95 GND.n94 60.0588
R8872 GND.n53 GND.n52 60.0588
R8873 GND.n55 GND.n54 60.0588
R8874 GND.n57 GND.n56 60.0588
R8875 GND.n16 GND.n15 60.0588
R8876 GND.n18 GND.n17 60.0588
R8877 GND.n20 GND.n19 60.0588
R8878 GND.n209 GND.n208 60.0588
R8879 GND.n207 GND.n206 60.0588
R8880 GND.n205 GND.n204 60.0588
R8881 GND.n171 GND.n170 60.0588
R8882 GND.n169 GND.n168 60.0588
R8883 GND.n167 GND.n166 60.0588
R8884 GND.n134 GND.n133 60.0588
R8885 GND.n132 GND.n131 60.0588
R8886 GND.n130 GND.n129 60.0588
R8887 GND.n1821 GND.n1820 59.5399
R8888 GND.n6534 GND.n6533 59.5399
R8889 GND.n5640 GND.n1818 59.5399
R8890 GND.n6628 GND.n6623 59.5399
R8891 GND.n5719 GND.n5718 52.946
R8892 GND.n1408 GND.n1407 52.946
R8893 GND.t145 GND.n78 52.3082
R8894 GND.t130 GND.n99 52.3082
R8895 GND.t144 GND.n40 52.3082
R8896 GND.t91 GND.n61 52.3082
R8897 GND.t93 GND.n3 52.3082
R8898 GND.t141 GND.n24 52.3082
R8899 GND.t95 GND.n213 52.3082
R8900 GND.t135 GND.n192 52.3082
R8901 GND.t115 GND.n175 52.3082
R8902 GND.t121 GND.n154 52.3082
R8903 GND.t126 GND.n138 52.3082
R8904 GND.t146 GND.n117 52.3082
R8905 GND.n6621 GND.n1179 44.3322
R8906 GND.n5720 GND.n5719 42.2793
R8907 GND.n5613 GND.n5607 42.2793
R8908 GND.n1758 GND.n1757 42.2793
R8909 GND.n6684 GND.n6683 42.2793
R8910 GND.n563 GND.n562 42.2793
R8911 GND.n7448 GND.n543 42.2793
R8912 GND.n582 GND.n581 42.2793
R8913 GND.n1369 GND.n1364 42.2793
R8914 GND.n3068 GND.n3067 42.2793
R8915 GND.n3088 GND.n3087 42.2793
R8916 GND.n3120 GND.n3119 42.2793
R8917 GND.n6284 GND.n1408 42.2793
R8918 GND.n3185 GND.n3050 39.2524
R8919 GND.n5034 GND.n2771 38.4083
R8920 GND.n5050 GND.n2771 38.4083
R8921 GND.n5050 GND.n2762 38.4083
R8922 GND.n5058 GND.n2762 38.4083
R8923 GND.n5058 GND.n2540 38.4083
R8924 GND.n5210 GND.n2540 38.4083
R8925 GND.n5210 GND.n2543 38.4083
R8926 GND.n2757 GND.n2543 38.4083
R8927 GND.n5220 GND.n2530 38.4083
R8928 GND.n2737 GND.n2530 38.4083
R8929 GND.n5075 GND.n2737 38.4083
R8930 GND.n5075 GND.n2727 38.4083
R8931 GND.n5082 GND.n2727 38.4083
R8932 GND.n5082 GND.n2715 38.4083
R8933 GND.n5175 GND.n2715 38.4083
R8934 GND.n5175 GND.n2577 38.4083
R8935 GND.n5182 GND.n2577 38.4083
R8936 GND.n5182 GND.n2506 38.4083
R8937 GND.n5229 GND.n2506 38.4083
R8938 GND.n5241 GND.n2495 38.4083
R8939 GND.n5241 GND.n2486 38.4083
R8940 GND.n5249 GND.n2486 38.4083
R8941 GND.n5249 GND.n2475 38.4083
R8942 GND.n5261 GND.n2475 38.4083
R8943 GND.n5261 GND.n2466 38.4083
R8944 GND.n5269 GND.n2466 38.4083
R8945 GND.n5269 GND.n2454 38.4083
R8946 GND.n5281 GND.n2454 38.4083
R8947 GND.n5281 GND.n2457 38.4083
R8948 GND.n5289 GND.n2435 38.4083
R8949 GND.n5301 GND.n2435 38.4083
R8950 GND.n5301 GND.n2426 38.4083
R8951 GND.n5309 GND.n2426 38.4083
R8952 GND.n5309 GND.n2415 38.4083
R8953 GND.n5321 GND.n2415 38.4083
R8954 GND.n5321 GND.n2406 38.4083
R8955 GND.n5329 GND.n2406 38.4083
R8956 GND.n5329 GND.n2394 38.4083
R8957 GND.n5341 GND.n2394 38.4083
R8958 GND.n5341 GND.n2397 38.4083
R8959 GND.n5349 GND.n2375 38.4083
R8960 GND.n5361 GND.n2375 38.4083
R8961 GND.n5361 GND.n2366 38.4083
R8962 GND.n5369 GND.n2366 38.4083
R8963 GND.n5369 GND.n2355 38.4083
R8964 GND.n5386 GND.n2355 38.4083
R8965 GND.n5386 GND.n2345 38.4083
R8966 GND.n5396 GND.n2345 38.4083
R8967 GND.n5396 GND.n2338 38.4083
R8968 GND.n5455 GND.n2338 38.4083
R8969 GND.n5466 GND.n2319 38.4083
R8970 GND.n5474 GND.n2319 38.4083
R8971 GND.n5474 GND.n2308 38.4083
R8972 GND.n5486 GND.n2308 38.4083
R8973 GND.n5486 GND.n2299 38.4083
R8974 GND.n5494 GND.n2299 38.4083
R8975 GND.n5494 GND.n2288 38.4083
R8976 GND.n5506 GND.n2288 38.4083
R8977 GND.n5506 GND.n2279 38.4083
R8978 GND.n5514 GND.n2279 38.4083
R8979 GND.n5514 GND.n2267 38.4083
R8980 GND.n5526 GND.n2267 38.4083
R8981 GND.n5526 GND.n2270 38.4083
R8982 GND.n5534 GND.n2248 38.4083
R8983 GND.n5550 GND.n2248 38.4083
R8984 GND.n5550 GND.n2239 38.4083
R8985 GND.n5559 GND.n2239 38.4083
R8986 GND.n5559 GND.n1737 38.4083
R8987 GND.n5691 GND.n1737 38.4083
R8988 GND.n5691 GND.n1740 38.4083
R8989 GND.n5685 GND.n5684 38.4083
R8990 GND.n5684 GND.n5683 38.4083
R8991 GND.n5683 GND.n1778 38.4083
R8992 GND.n5677 GND.n1778 38.4083
R8993 GND.n6610 GND.n6609 38.4083
R8994 GND.n6609 GND.n6608 38.4083
R8995 GND.n6608 GND.n940 38.4083
R8996 GND.n6726 GND.n940 38.4083
R8997 GND.n6734 GND.n931 38.4083
R8998 GND.n6734 GND.n918 38.4083
R8999 GND.n6752 GND.n918 38.4083
R9000 GND.n6752 GND.n908 38.4083
R9001 GND.n6762 GND.n908 38.4083
R9002 GND.n6762 GND.n901 38.4083
R9003 GND.n6852 GND.n901 38.4083
R9004 GND.n6863 GND.n882 38.4083
R9005 GND.n6871 GND.n882 38.4083
R9006 GND.n6871 GND.n871 38.4083
R9007 GND.n6883 GND.n871 38.4083
R9008 GND.n6883 GND.n862 38.4083
R9009 GND.n6891 GND.n862 38.4083
R9010 GND.n6891 GND.n851 38.4083
R9011 GND.n6903 GND.n851 38.4083
R9012 GND.n6903 GND.n842 38.4083
R9013 GND.n6911 GND.n842 38.4083
R9014 GND.n6911 GND.n830 38.4083
R9015 GND.n6923 GND.n830 38.4083
R9016 GND.n6923 GND.n833 38.4083
R9017 GND.n6931 GND.n811 38.4083
R9018 GND.n6943 GND.n811 38.4083
R9019 GND.n6943 GND.n802 38.4083
R9020 GND.n6951 GND.n802 38.4083
R9021 GND.n6951 GND.n791 38.4083
R9022 GND.n6963 GND.n791 38.4083
R9023 GND.n6963 GND.n782 38.4083
R9024 GND.n6971 GND.n782 38.4083
R9025 GND.n6971 GND.n771 38.4083
R9026 GND.n6983 GND.n771 38.4083
R9027 GND.n6991 GND.n762 38.4083
R9028 GND.n6991 GND.n751 38.4083
R9029 GND.n7003 GND.n751 38.4083
R9030 GND.n7003 GND.n742 38.4083
R9031 GND.n7011 GND.n742 38.4083
R9032 GND.n7011 GND.n730 38.4083
R9033 GND.n7027 GND.n730 38.4083
R9034 GND.n7027 GND.n720 38.4083
R9035 GND.n7037 GND.n720 38.4083
R9036 GND.n7037 GND.n713 38.4083
R9037 GND.n7060 GND.n713 38.4083
R9038 GND.n7071 GND.n694 38.4083
R9039 GND.n7079 GND.n694 38.4083
R9040 GND.n7079 GND.n682 38.4083
R9041 GND.n7099 GND.n682 38.4083
R9042 GND.n7099 GND.n673 38.4083
R9043 GND.n7107 GND.n673 38.4083
R9044 GND.n7107 GND.n654 38.4083
R9045 GND.n7135 GND.n654 38.4083
R9046 GND.n7135 GND.n657 38.4083
R9047 GND.n7129 GND.n657 38.4083
R9048 GND.n7145 GND.n635 38.4083
R9049 GND.n7160 GND.n635 38.4083
R9050 GND.n7160 GND.n630 38.4083
R9051 GND.n7168 GND.n630 38.4083
R9052 GND.n7168 GND.n233 38.4083
R9053 GND.n7641 GND.n233 38.4083
R9054 GND.n7641 GND.n236 38.4083
R9055 GND.n619 GND.n236 38.4083
R9056 GND.n7208 GND.n619 38.4083
R9057 GND.n7208 GND.n252 38.4083
R9058 GND.n7632 GND.n252 38.4083
R9059 GND.n7626 GND.n264 38.4083
R9060 GND.n7626 GND.n267 38.4083
R9061 GND.n7620 GND.n267 38.4083
R9062 GND.n7620 GND.n277 38.4083
R9063 GND.n7614 GND.n277 38.4083
R9064 GND.n7614 GND.n287 38.4083
R9065 GND.n7608 GND.n287 38.4083
R9066 GND.n7608 GND.n298 38.4083
R9067 GND.n7602 GND.n298 38.4083
R9068 GND.n7596 GND.n319 38.4083
R9069 GND.n7590 GND.n319 38.4083
R9070 GND.n7590 GND.n331 38.4083
R9071 GND.n7584 GND.n331 38.4083
R9072 GND.n7584 GND.n341 38.4083
R9073 GND.n7578 GND.n341 38.4083
R9074 GND.n7578 GND.n350 38.4083
R9075 GND.n7572 GND.n350 38.4083
R9076 GND.n7572 GND.n360 38.4083
R9077 GND.n7566 GND.n360 38.4083
R9078 GND.n7566 GND.n369 38.4083
R9079 GND.n7560 GND.n379 38.4083
R9080 GND.n7554 GND.n379 38.4083
R9081 GND.n7554 GND.n388 38.4083
R9082 GND.n7548 GND.n388 38.4083
R9083 GND.n7548 GND.n398 38.4083
R9084 GND.n7542 GND.n398 38.4083
R9085 GND.n7542 GND.n407 38.4083
R9086 GND.n7536 GND.n407 38.4083
R9087 GND.n7536 GND.n417 38.4083
R9088 GND.n7530 GND.n417 38.4083
R9089 GND.n7524 GND.n433 38.4083
R9090 GND.n7524 GND.n436 38.4083
R9091 GND.n7518 GND.n436 38.4083
R9092 GND.n7518 GND.n445 38.4083
R9093 GND.n7512 GND.n456 38.4083
R9094 GND.n7506 GND.n456 38.4083
R9095 GND.n7506 GND.n465 38.4083
R9096 GND.n7500 GND.n465 38.4083
R9097 GND.n7500 GND.n475 38.4083
R9098 GND.n7494 GND.n475 38.4083
R9099 GND.n7494 GND.n484 38.4083
R9100 GND.n7488 GND.n484 38.4083
R9101 GND.n7482 GND.n500 38.4083
R9102 GND.n7482 GND.n503 38.4083
R9103 GND.n7476 GND.n503 38.4083
R9104 GND.n7476 GND.n513 38.4083
R9105 GND.n7470 GND.n513 38.4083
R9106 GND.n7470 GND.n522 38.4083
R9107 GND.n5630 GND.n2228 36.9518
R9108 GND.n6709 GND.n6671 36.9518
R9109 GND.n5455 GND.t92 36.872
R9110 GND.n6931 GND.t120 36.872
R9111 GND.n7530 GND.t94 36.872
R9112 GND.n2185 GND.n1822 35.7468
R9113 GND.n6578 GND.n6574 35.7468
R9114 GND.n91 GND.n89 35.0348
R9115 GND.n53 GND.n51 35.0348
R9116 GND.n16 GND.n14 35.0348
R9117 GND.n205 GND.n203 35.0348
R9118 GND.n167 GND.n165 35.0348
R9119 GND.n130 GND.n128 35.0348
R9120 GND.n7602 GND.n307 34.9516
R9121 GND.n1814 GND.n1813 34.8345
R9122 GND.n1178 GND.n1177 34.8345
R9123 GND.n453 GND.n445 32.6471
R9124 GND.n2457 GND.t96 32.2631
R9125 GND.n7071 GND.t98 32.2631
R9126 GND.n7234 GND.t102 32.2631
R9127 GND.n5632 GND.n5630 30.6565
R9128 GND.n6709 GND.n6667 30.6565
R9129 GND.n111 GND.n110 30.052
R9130 GND.n73 GND.n72 30.052
R9131 GND.n36 GND.n35 30.052
R9132 GND.n225 GND.n224 30.052
R9133 GND.n187 GND.n186 30.052
R9134 GND.n150 GND.n149 30.052
R9135 GND.n6576 GND.n1151 28.4223
R9136 GND.n2757 GND.t86 27.6541
R9137 GND.t112 GND.n2495 27.6541
R9138 GND.n7129 GND.t100 27.6541
R9139 GND.n264 GND.t122 27.6541
R9140 GND.n2270 GND.t9 26.886
R9141 GND.n6863 GND.t45 26.886
R9142 GND.n7488 GND.t20 26.886
R9143 GND.t13 GND.n1832 26.1178
R9144 GND.n2168 GND.n1840 26.1178
R9145 GND.n1993 GND.n1850 26.1178
R9146 GND.n2154 GND.n1858 26.1178
R9147 GND.n2006 GND.n1868 26.1178
R9148 GND.n2140 GND.n1876 26.1178
R9149 GND.n2132 GND.n1889 26.1178
R9150 GND.n2027 GND.n1897 26.1178
R9151 GND.n2118 GND.n1907 26.1178
R9152 GND.n2040 GND.n1915 26.1178
R9153 GND.n2104 GND.n1925 26.1178
R9154 GND.n2053 GND.n1933 26.1178
R9155 GND.n2090 GND.n1943 26.1178
R9156 GND.n2068 GND.n1951 26.1178
R9157 GND.n5764 GND.n5763 26.1178
R9158 GND.n6338 GND.n6337 26.1178
R9159 GND.n6356 GND.n1309 26.1178
R9160 GND.n6383 GND.n1294 26.1178
R9161 GND.n6390 GND.n6389 26.1178
R9162 GND.n6408 GND.n1280 26.1178
R9163 GND.n6414 GND.n1276 26.1178
R9164 GND.n6432 GND.n1260 26.1178
R9165 GND.n6443 GND.n1249 26.1178
R9166 GND.n6464 GND.n1240 26.1178
R9167 GND.n6482 GND.n1230 26.1178
R9168 GND.n6488 GND.n1226 26.1178
R9169 GND.n6515 GND.n1210 26.1178
R9170 GND.n6522 GND.n6521 26.1178
R9171 GND.n6587 GND.n1196 26.1178
R9172 GND.n6593 GND.n1192 26.1178
R9173 GND.n1777 GND.n1740 25.3497
R9174 GND.n2139 GND.n1878 25.3497
R9175 GND.n2133 GND.n1887 25.3497
R9176 GND.n2076 GND.n1710 25.3497
R9177 GND.n6350 GND.n1313 25.3497
R9178 GND.n6463 GND.n1242 25.3497
R9179 GND.n6470 GND.n1236 25.3497
R9180 GND.n6725 GND.n931 25.3497
R9181 GND.n2147 GND.n2146 23.8133
R9182 GND.n2126 GND.n2125 23.8133
R9183 GND.n2084 GND.n1949 23.8133
R9184 GND.n5770 GND.n1706 23.8133
R9185 GND.n6330 GND.n1323 23.8133
R9186 GND.n6377 GND.n6376 23.8133
R9187 GND.n6450 GND.n6449 23.8133
R9188 GND.n6489 GND.n1224 23.8133
R9189 GND.n3185 GND.n3039 23.6462
R9190 GND.n3201 GND.n3039 23.6462
R9191 GND.n3201 GND.n3030 23.6462
R9192 GND.n3211 GND.n3030 23.6462
R9193 GND.n3211 GND.n3023 23.6462
R9194 GND.n3325 GND.n3023 23.6462
R9195 GND.n3333 GND.n3003 23.6462
R9196 GND.n3341 GND.n3003 23.6462
R9197 GND.n3341 GND.n2990 23.6462
R9198 GND.n3350 GND.n2990 23.6462
R9199 GND.n3350 GND.n2982 23.6462
R9200 GND.n3358 GND.n2982 23.6462
R9201 GND.n3358 GND.n2969 23.6462
R9202 GND.n3367 GND.n2969 23.6462
R9203 GND.n3367 GND.n2961 23.6462
R9204 GND.n3375 GND.n2961 23.6462
R9205 GND.n3375 GND.n2947 23.6462
R9206 GND.n3384 GND.n2947 23.6462
R9207 GND.n3384 GND.n2950 23.6462
R9208 GND.n3392 GND.n2927 23.6462
R9209 GND.n3401 GND.n2927 23.6462
R9210 GND.n3401 GND.n2919 23.6462
R9211 GND.n3409 GND.n2919 23.6462
R9212 GND.n3409 GND.n2906 23.6462
R9213 GND.n3418 GND.n2906 23.6462
R9214 GND.n3418 GND.n2898 23.6462
R9215 GND.n3426 GND.n2898 23.6462
R9216 GND.n3426 GND.n2885 23.6462
R9217 GND.n3435 GND.n2885 23.6462
R9218 GND.n3443 GND.n2877 23.6462
R9219 GND.n3443 GND.n2864 23.6462
R9220 GND.n3452 GND.n2864 23.6462
R9221 GND.n3452 GND.n2856 23.6462
R9222 GND.n3460 GND.n2856 23.6462
R9223 GND.n3460 GND.n2843 23.6462
R9224 GND.n3469 GND.n2843 23.6462
R9225 GND.n3469 GND.n2835 23.6462
R9226 GND.n3477 GND.n2835 23.6462
R9227 GND.n3477 GND.n2824 23.6462
R9228 GND.n3492 GND.n2824 23.6462
R9229 GND.n4192 GND.n453 23.2004
R9230 GND.n5349 GND.t88 23.0452
R9231 GND.n6983 GND.t117 23.0452
R9232 GND.n7560 GND.t108 23.0452
R9233 GND.n3392 GND.t90 22.7004
R9234 GND.n1975 GND.n1824 22.277
R9235 GND.n2153 GND.n1860 22.277
R9236 GND.n2119 GND.n1905 22.277
R9237 GND.n2050 GND.n1941 22.277
R9238 GND.n1295 GND.n1290 22.277
R9239 GND.n1262 GND.n1261 22.277
R9240 GND.n6509 GND.n6508 22.277
R9241 GND.n6617 GND.n1182 22.277
R9242 GND.n5025 GND.n3520 21.5181
R9243 GND.n5676 GND.n1807 21.1248
R9244 GND.n6664 GND.n1151 21.1248
R9245 GND.n2174 GND.n1834 20.7407
R9246 GND.n2161 GND.n2160 20.7407
R9247 GND.n2112 GND.n2111 20.7407
R9248 GND.n2098 GND.n1931 20.7407
R9249 GND.n6396 GND.n1286 20.7407
R9250 GND.n6426 GND.n1266 20.7407
R9251 GND.n1211 GND.n1206 20.7407
R9252 GND.n6586 GND.n1190 20.7407
R9253 GND.n1977 GND.n1816 20.1371
R9254 GND.n6621 GND.n6620 20.1371
R9255 GND.t110 GND.n2790 19.8629
R9256 GND.n1811 GND.t77 19.8005
R9257 GND.n1811 GND.t14 19.8005
R9258 GND.n1175 GND.t71 19.8005
R9259 GND.n1175 GND.t43 19.8005
R9260 GND.n5733 GND.n5732 19.3944
R9261 GND.n5732 GND.n5731 19.3944
R9262 GND.n5731 GND.n5726 19.3944
R9263 GND.n5759 GND.n1722 19.3944
R9264 GND.n5759 GND.n1723 19.3944
R9265 GND.n5755 GND.n1723 19.3944
R9266 GND.n5755 GND.n5754 19.3944
R9267 GND.n5754 GND.n5701 19.3944
R9268 GND.n5750 GND.n5701 19.3944
R9269 GND.n5750 GND.n5749 19.3944
R9270 GND.n5749 GND.n5748 19.3944
R9271 GND.n5748 GND.n5707 19.3944
R9272 GND.n5744 GND.n5707 19.3944
R9273 GND.n5744 GND.n5743 19.3944
R9274 GND.n5743 GND.n5742 19.3944
R9275 GND.n5742 GND.n5713 19.3944
R9276 GND.n5738 GND.n5713 19.3944
R9277 GND.n5738 GND.n5737 19.3944
R9278 GND.n5737 GND.n5736 19.3944
R9279 GND.n5727 GND.n1673 19.3944
R9280 GND.n5830 GND.n1673 19.3944
R9281 GND.n5830 GND.n1670 19.3944
R9282 GND.n5836 GND.n1670 19.3944
R9283 GND.n5836 GND.n1671 19.3944
R9284 GND.n1671 GND.n1646 19.3944
R9285 GND.n5863 GND.n1646 19.3944
R9286 GND.n5864 GND.n5863 19.3944
R9287 GND.n5864 GND.n1643 19.3944
R9288 GND.n5876 GND.n1643 19.3944
R9289 GND.n5876 GND.n1644 19.3944
R9290 GND.n5872 GND.n1644 19.3944
R9291 GND.n5872 GND.n5871 19.3944
R9292 GND.n5871 GND.n5870 19.3944
R9293 GND.n5870 GND.n1575 19.3944
R9294 GND.n1575 GND.n1573 19.3944
R9295 GND.n5951 GND.n1573 19.3944
R9296 GND.n5951 GND.n1570 19.3944
R9297 GND.n5974 GND.n1570 19.3944
R9298 GND.n5974 GND.n1571 19.3944
R9299 GND.n5970 GND.n1571 19.3944
R9300 GND.n5970 GND.n5969 19.3944
R9301 GND.n5969 GND.n5968 19.3944
R9302 GND.n5968 GND.n5956 19.3944
R9303 GND.n5964 GND.n5956 19.3944
R9304 GND.n5964 GND.n5963 19.3944
R9305 GND.n5963 GND.n5962 19.3944
R9306 GND.n5962 GND.n1494 19.3944
R9307 GND.n6107 GND.n1494 19.3944
R9308 GND.n6108 GND.n6107 19.3944
R9309 GND.n6108 GND.n1491 19.3944
R9310 GND.n6130 GND.n1491 19.3944
R9311 GND.n6130 GND.n1492 19.3944
R9312 GND.n6126 GND.n1492 19.3944
R9313 GND.n6126 GND.n6125 19.3944
R9314 GND.n6125 GND.n6124 19.3944
R9315 GND.n6124 GND.n6115 19.3944
R9316 GND.n6120 GND.n6115 19.3944
R9317 GND.n6120 GND.n6119 19.3944
R9318 GND.n6119 GND.n1418 19.3944
R9319 GND.n6270 GND.n1418 19.3944
R9320 GND.n6270 GND.n1416 19.3944
R9321 GND.n6274 GND.n1416 19.3944
R9322 GND.n6275 GND.n6274 19.3944
R9323 GND.n5567 GND.n2235 19.3944
R9324 GND.n5571 GND.n2235 19.3944
R9325 GND.n5571 GND.n2233 19.3944
R9326 GND.n5577 GND.n2233 19.3944
R9327 GND.n5577 GND.n2231 19.3944
R9328 GND.n5582 GND.n2231 19.3944
R9329 GND.n5582 GND.n2226 19.3944
R9330 GND.n5629 GND.n5589 19.3944
R9331 GND.n5625 GND.n5589 19.3944
R9332 GND.n5625 GND.n5624 19.3944
R9333 GND.n5624 GND.n5623 19.3944
R9334 GND.n5623 GND.n5597 19.3944
R9335 GND.n5619 GND.n5597 19.3944
R9336 GND.n5619 GND.n5618 19.3944
R9337 GND.n5618 GND.n5617 19.3944
R9338 GND.n5617 GND.n5605 19.3944
R9339 GND.n1774 GND.n1773 19.3944
R9340 GND.n1770 GND.n1769 19.3944
R9341 GND.n1766 GND.n1765 19.3944
R9342 GND.n1762 GND.n1761 19.3944
R9343 GND.n3188 GND.n3048 19.3944
R9344 GND.n3197 GND.n3188 19.3944
R9345 GND.n3197 GND.n3196 19.3944
R9346 GND.n3196 GND.n3195 19.3944
R9347 GND.n3195 GND.n3021 19.3944
R9348 GND.n3327 GND.n3021 19.3944
R9349 GND.n3329 GND.n3327 19.3944
R9350 GND.n3329 GND.n3328 19.3944
R9351 GND.n3328 GND.n3001 19.3944
R9352 GND.n3344 GND.n3001 19.3944
R9353 GND.n3346 GND.n3344 19.3944
R9354 GND.n3346 GND.n3345 19.3944
R9355 GND.n3345 GND.n2980 19.3944
R9356 GND.n3361 GND.n2980 19.3944
R9357 GND.n3363 GND.n3361 19.3944
R9358 GND.n3363 GND.n3362 19.3944
R9359 GND.n3362 GND.n2959 19.3944
R9360 GND.n3378 GND.n2959 19.3944
R9361 GND.n3380 GND.n3378 19.3944
R9362 GND.n3380 GND.n3379 19.3944
R9363 GND.n3379 GND.n2938 19.3944
R9364 GND.n3395 GND.n2938 19.3944
R9365 GND.n3397 GND.n3395 19.3944
R9366 GND.n3397 GND.n3396 19.3944
R9367 GND.n3396 GND.n2917 19.3944
R9368 GND.n3412 GND.n2917 19.3944
R9369 GND.n3414 GND.n3412 19.3944
R9370 GND.n3414 GND.n3413 19.3944
R9371 GND.n3413 GND.n2896 19.3944
R9372 GND.n3429 GND.n2896 19.3944
R9373 GND.n3431 GND.n3429 19.3944
R9374 GND.n3431 GND.n3430 19.3944
R9375 GND.n3430 GND.n2875 19.3944
R9376 GND.n3446 GND.n2875 19.3944
R9377 GND.n3448 GND.n3446 19.3944
R9378 GND.n3448 GND.n3447 19.3944
R9379 GND.n3447 GND.n2854 19.3944
R9380 GND.n3463 GND.n2854 19.3944
R9381 GND.n3465 GND.n3463 19.3944
R9382 GND.n3465 GND.n3464 19.3944
R9383 GND.n3464 GND.n2833 19.3944
R9384 GND.n3480 GND.n2833 19.3944
R9385 GND.n3488 GND.n3480 19.3944
R9386 GND.n3488 GND.n3487 19.3944
R9387 GND.n3487 GND.n3486 19.3944
R9388 GND.n3486 GND.n3485 19.3944
R9389 GND.n3485 GND.n2777 19.3944
R9390 GND.n5048 GND.n2777 19.3944
R9391 GND.n5048 GND.n2778 19.3944
R9392 GND.n5044 GND.n2778 19.3944
R9393 GND.n5044 GND.n2547 19.3944
R9394 GND.n5208 GND.n2547 19.3944
R9395 GND.n5208 GND.n2548 19.3944
R9396 GND.n5204 GND.n2548 19.3944
R9397 GND.n5204 GND.n5203 19.3944
R9398 GND.n5203 GND.n5202 19.3944
R9399 GND.n5202 GND.n2556 19.3944
R9400 GND.n5198 GND.n2556 19.3944
R9401 GND.n5198 GND.n5197 19.3944
R9402 GND.n5197 GND.n5196 19.3944
R9403 GND.n5196 GND.n2565 19.3944
R9404 GND.n5192 GND.n2565 19.3944
R9405 GND.n5192 GND.n5191 19.3944
R9406 GND.n5191 GND.n5190 19.3944
R9407 GND.n5190 GND.n2574 19.3944
R9408 GND.n5186 GND.n2574 19.3944
R9409 GND.n5186 GND.n2501 19.3944
R9410 GND.n5239 GND.n2501 19.3944
R9411 GND.n5239 GND.n2502 19.3944
R9412 GND.n5235 GND.n2502 19.3944
R9413 GND.n5235 GND.n2481 19.3944
R9414 GND.n5259 GND.n2481 19.3944
R9415 GND.n5259 GND.n2482 19.3944
R9416 GND.n5255 GND.n2482 19.3944
R9417 GND.n5255 GND.n2461 19.3944
R9418 GND.n5279 GND.n2461 19.3944
R9419 GND.n5279 GND.n2462 19.3944
R9420 GND.n5275 GND.n2462 19.3944
R9421 GND.n5275 GND.n2441 19.3944
R9422 GND.n5299 GND.n2441 19.3944
R9423 GND.n5299 GND.n2442 19.3944
R9424 GND.n5295 GND.n2442 19.3944
R9425 GND.n5295 GND.n2421 19.3944
R9426 GND.n5319 GND.n2421 19.3944
R9427 GND.n5319 GND.n2422 19.3944
R9428 GND.n5315 GND.n2422 19.3944
R9429 GND.n5315 GND.n2401 19.3944
R9430 GND.n5339 GND.n2401 19.3944
R9431 GND.n5339 GND.n2402 19.3944
R9432 GND.n5335 GND.n2402 19.3944
R9433 GND.n5335 GND.n2381 19.3944
R9434 GND.n5359 GND.n2381 19.3944
R9435 GND.n5359 GND.n2382 19.3944
R9436 GND.n5355 GND.n2382 19.3944
R9437 GND.n5355 GND.n2361 19.3944
R9438 GND.n5384 GND.n2361 19.3944
R9439 GND.n5384 GND.n2362 19.3944
R9440 GND.n5380 GND.n2362 19.3944
R9441 GND.n5380 GND.n5379 19.3944
R9442 GND.n5379 GND.n2333 19.3944
R9443 GND.n5464 GND.n2333 19.3944
R9444 GND.n5464 GND.n2334 19.3944
R9445 GND.n5460 GND.n2334 19.3944
R9446 GND.n5460 GND.n2314 19.3944
R9447 GND.n5484 GND.n2314 19.3944
R9448 GND.n5484 GND.n2315 19.3944
R9449 GND.n5480 GND.n2315 19.3944
R9450 GND.n5480 GND.n2294 19.3944
R9451 GND.n5504 GND.n2294 19.3944
R9452 GND.n5504 GND.n2295 19.3944
R9453 GND.n5500 GND.n2295 19.3944
R9454 GND.n5500 GND.n2274 19.3944
R9455 GND.n5524 GND.n2274 19.3944
R9456 GND.n5524 GND.n2275 19.3944
R9457 GND.n5520 GND.n2275 19.3944
R9458 GND.n5520 GND.n2254 19.3944
R9459 GND.n5548 GND.n2254 19.3944
R9460 GND.n5548 GND.n2255 19.3944
R9461 GND.n5544 GND.n2255 19.3944
R9462 GND.n5544 GND.n1734 19.3944
R9463 GND.n5693 GND.n1734 19.3944
R9464 GND.n5022 GND.n5021 19.3944
R9465 GND.n5021 GND.n5020 19.3944
R9466 GND.n5020 GND.n5019 19.3944
R9467 GND.n5019 GND.n5017 19.3944
R9468 GND.n5017 GND.n5014 19.3944
R9469 GND.n5014 GND.n5013 19.3944
R9470 GND.n5013 GND.n5010 19.3944
R9471 GND.n5010 GND.n5009 19.3944
R9472 GND.n5009 GND.n5006 19.3944
R9473 GND.n5006 GND.n5005 19.3944
R9474 GND.n5005 GND.n5002 19.3944
R9475 GND.n5002 GND.n5001 19.3944
R9476 GND.n5001 GND.n4998 19.3944
R9477 GND.n4998 GND.n4997 19.3944
R9478 GND.n4997 GND.n4994 19.3944
R9479 GND.n4994 GND.n4993 19.3944
R9480 GND.n4993 GND.n4990 19.3944
R9481 GND.n4990 GND.n4989 19.3944
R9482 GND.n4989 GND.n4986 19.3944
R9483 GND.n4986 GND.n4985 19.3944
R9484 GND.n4985 GND.n4982 19.3944
R9485 GND.n4982 GND.n4981 19.3944
R9486 GND.n4981 GND.n4978 19.3944
R9487 GND.n4978 GND.n4977 19.3944
R9488 GND.n4977 GND.n4974 19.3944
R9489 GND.n4974 GND.n4973 19.3944
R9490 GND.n4973 GND.n4970 19.3944
R9491 GND.n4970 GND.n4969 19.3944
R9492 GND.n4969 GND.n4966 19.3944
R9493 GND.n4966 GND.n4965 19.3944
R9494 GND.n4965 GND.n4962 19.3944
R9495 GND.n4962 GND.n4961 19.3944
R9496 GND.n4961 GND.n4958 19.3944
R9497 GND.n4958 GND.n4957 19.3944
R9498 GND.n4957 GND.n4954 19.3944
R9499 GND.n4954 GND.n4953 19.3944
R9500 GND.n4953 GND.n4950 19.3944
R9501 GND.n4950 GND.n4949 19.3944
R9502 GND.n4949 GND.n4946 19.3944
R9503 GND.n4946 GND.n4945 19.3944
R9504 GND.n4945 GND.n4942 19.3944
R9505 GND.n4942 GND.n4941 19.3944
R9506 GND.n4941 GND.n4938 19.3944
R9507 GND.n4938 GND.n4937 19.3944
R9508 GND.n4937 GND.n4934 19.3944
R9509 GND.n4934 GND.n4933 19.3944
R9510 GND.n4933 GND.n4930 19.3944
R9511 GND.n4930 GND.n4929 19.3944
R9512 GND.n4929 GND.n4926 19.3944
R9513 GND.n4926 GND.n4925 19.3944
R9514 GND.n4925 GND.n4922 19.3944
R9515 GND.n4922 GND.n4921 19.3944
R9516 GND.n4921 GND.n4918 19.3944
R9517 GND.n4918 GND.n2788 19.3944
R9518 GND.n5028 GND.n2788 19.3944
R9519 GND.n5029 GND.n5028 19.3944
R9520 GND.n4861 GND.n4860 19.3944
R9521 GND.n4860 GND.n3525 19.3944
R9522 GND.n4854 GND.n3525 19.3944
R9523 GND.n4854 GND.n4853 19.3944
R9524 GND.n4853 GND.n4852 19.3944
R9525 GND.n4852 GND.n3534 19.3944
R9526 GND.n4846 GND.n3534 19.3944
R9527 GND.n4846 GND.n4845 19.3944
R9528 GND.n4845 GND.n4844 19.3944
R9529 GND.n4844 GND.n3542 19.3944
R9530 GND.n4838 GND.n3542 19.3944
R9531 GND.n4838 GND.n4837 19.3944
R9532 GND.n4837 GND.n4836 19.3944
R9533 GND.n4836 GND.n3550 19.3944
R9534 GND.n4830 GND.n3550 19.3944
R9535 GND.n4830 GND.n4829 19.3944
R9536 GND.n4829 GND.n4828 19.3944
R9537 GND.n4828 GND.n3558 19.3944
R9538 GND.n4822 GND.n3558 19.3944
R9539 GND.n4822 GND.n4821 19.3944
R9540 GND.n4821 GND.n4820 19.3944
R9541 GND.n4820 GND.n3566 19.3944
R9542 GND.n4814 GND.n3566 19.3944
R9543 GND.n4814 GND.n4813 19.3944
R9544 GND.n4813 GND.n4812 19.3944
R9545 GND.n4812 GND.n3574 19.3944
R9546 GND.n4806 GND.n3574 19.3944
R9547 GND.n4806 GND.n4805 19.3944
R9548 GND.n4805 GND.n4804 19.3944
R9549 GND.n4804 GND.n3582 19.3944
R9550 GND.n4798 GND.n3582 19.3944
R9551 GND.n4798 GND.n4797 19.3944
R9552 GND.n4797 GND.n4796 19.3944
R9553 GND.n4796 GND.n3590 19.3944
R9554 GND.n4790 GND.n3590 19.3944
R9555 GND.n4790 GND.n4789 19.3944
R9556 GND.n4789 GND.n4788 19.3944
R9557 GND.n4788 GND.n3598 19.3944
R9558 GND.n4782 GND.n3598 19.3944
R9559 GND.n4782 GND.n4781 19.3944
R9560 GND.n4781 GND.n4780 19.3944
R9561 GND.n4780 GND.n3606 19.3944
R9562 GND.n4774 GND.n3606 19.3944
R9563 GND.n4774 GND.n4773 19.3944
R9564 GND.n4773 GND.n4772 19.3944
R9565 GND.n4772 GND.n3614 19.3944
R9566 GND.n4766 GND.n3614 19.3944
R9567 GND.n4766 GND.n4765 19.3944
R9568 GND.n4765 GND.n4764 19.3944
R9569 GND.n4764 GND.n3622 19.3944
R9570 GND.n4758 GND.n3622 19.3944
R9571 GND.n4758 GND.n4757 19.3944
R9572 GND.n4757 GND.n4756 19.3944
R9573 GND.n4756 GND.n3630 19.3944
R9574 GND.n4750 GND.n3630 19.3944
R9575 GND.n4750 GND.n4749 19.3944
R9576 GND.n4749 GND.n4748 19.3944
R9577 GND.n4748 GND.n3638 19.3944
R9578 GND.n4742 GND.n3638 19.3944
R9579 GND.n4742 GND.n4741 19.3944
R9580 GND.n4741 GND.n4740 19.3944
R9581 GND.n4740 GND.n3646 19.3944
R9582 GND.n4734 GND.n3646 19.3944
R9583 GND.n4734 GND.n4733 19.3944
R9584 GND.n4733 GND.n4732 19.3944
R9585 GND.n4732 GND.n3654 19.3944
R9586 GND.n4726 GND.n3654 19.3944
R9587 GND.n4726 GND.n4725 19.3944
R9588 GND.n4725 GND.n4724 19.3944
R9589 GND.n4724 GND.n3662 19.3944
R9590 GND.n4718 GND.n3662 19.3944
R9591 GND.n4718 GND.n4717 19.3944
R9592 GND.n4717 GND.n4716 19.3944
R9593 GND.n4716 GND.n3670 19.3944
R9594 GND.n4710 GND.n3670 19.3944
R9595 GND.n4710 GND.n4709 19.3944
R9596 GND.n4709 GND.n4708 19.3944
R9597 GND.n4708 GND.n3678 19.3944
R9598 GND.n4702 GND.n3678 19.3944
R9599 GND.n4702 GND.n4701 19.3944
R9600 GND.n4701 GND.n4700 19.3944
R9601 GND.n4700 GND.n3686 19.3944
R9602 GND.n4694 GND.n3686 19.3944
R9603 GND.n4694 GND.n4693 19.3944
R9604 GND.n4693 GND.n4692 19.3944
R9605 GND.n4692 GND.n3694 19.3944
R9606 GND.n4686 GND.n3694 19.3944
R9607 GND.n4686 GND.n4685 19.3944
R9608 GND.n4685 GND.n4684 19.3944
R9609 GND.n4684 GND.n3702 19.3944
R9610 GND.n4678 GND.n3702 19.3944
R9611 GND.n4678 GND.n4677 19.3944
R9612 GND.n4677 GND.n4676 19.3944
R9613 GND.n4676 GND.n3710 19.3944
R9614 GND.n4670 GND.n3710 19.3944
R9615 GND.n4670 GND.n4669 19.3944
R9616 GND.n4669 GND.n4668 19.3944
R9617 GND.n4668 GND.n3718 19.3944
R9618 GND.n4662 GND.n3718 19.3944
R9619 GND.n4662 GND.n4661 19.3944
R9620 GND.n4661 GND.n4660 19.3944
R9621 GND.n4660 GND.n3726 19.3944
R9622 GND.n4654 GND.n3726 19.3944
R9623 GND.n4654 GND.n4653 19.3944
R9624 GND.n4653 GND.n4652 19.3944
R9625 GND.n4652 GND.n3734 19.3944
R9626 GND.n4646 GND.n3734 19.3944
R9627 GND.n4646 GND.n4645 19.3944
R9628 GND.n4645 GND.n4644 19.3944
R9629 GND.n4644 GND.n3742 19.3944
R9630 GND.n4638 GND.n3742 19.3944
R9631 GND.n4638 GND.n4637 19.3944
R9632 GND.n4637 GND.n4636 19.3944
R9633 GND.n4636 GND.n3750 19.3944
R9634 GND.n4630 GND.n3750 19.3944
R9635 GND.n4630 GND.n4629 19.3944
R9636 GND.n4629 GND.n4628 19.3944
R9637 GND.n4628 GND.n3758 19.3944
R9638 GND.n4622 GND.n3758 19.3944
R9639 GND.n4622 GND.n4621 19.3944
R9640 GND.n4621 GND.n4620 19.3944
R9641 GND.n4620 GND.n3766 19.3944
R9642 GND.n4614 GND.n3766 19.3944
R9643 GND.n4614 GND.n4613 19.3944
R9644 GND.n4613 GND.n4612 19.3944
R9645 GND.n4612 GND.n3774 19.3944
R9646 GND.n4606 GND.n3774 19.3944
R9647 GND.n4606 GND.n4605 19.3944
R9648 GND.n4605 GND.n4604 19.3944
R9649 GND.n4604 GND.n3782 19.3944
R9650 GND.n4598 GND.n3782 19.3944
R9651 GND.n4598 GND.n4597 19.3944
R9652 GND.n4597 GND.n4596 19.3944
R9653 GND.n4596 GND.n3790 19.3944
R9654 GND.n4590 GND.n3790 19.3944
R9655 GND.n4590 GND.n4589 19.3944
R9656 GND.n4589 GND.n4588 19.3944
R9657 GND.n4588 GND.n3798 19.3944
R9658 GND.n4582 GND.n3798 19.3944
R9659 GND.n4582 GND.n4581 19.3944
R9660 GND.n4581 GND.n4580 19.3944
R9661 GND.n4580 GND.n3806 19.3944
R9662 GND.n4574 GND.n3806 19.3944
R9663 GND.n4574 GND.n4573 19.3944
R9664 GND.n4573 GND.n4572 19.3944
R9665 GND.n4572 GND.n3814 19.3944
R9666 GND.n4566 GND.n3814 19.3944
R9667 GND.n4566 GND.n4565 19.3944
R9668 GND.n4565 GND.n4564 19.3944
R9669 GND.n4564 GND.n3822 19.3944
R9670 GND.n4558 GND.n3822 19.3944
R9671 GND.n4558 GND.n4557 19.3944
R9672 GND.n4557 GND.n4556 19.3944
R9673 GND.n4556 GND.n3830 19.3944
R9674 GND.n4550 GND.n3830 19.3944
R9675 GND.n4550 GND.n4549 19.3944
R9676 GND.n4549 GND.n4548 19.3944
R9677 GND.n4548 GND.n3838 19.3944
R9678 GND.n4542 GND.n3838 19.3944
R9679 GND.n4542 GND.n4541 19.3944
R9680 GND.n4541 GND.n4540 19.3944
R9681 GND.n4540 GND.n3846 19.3944
R9682 GND.n4534 GND.n3846 19.3944
R9683 GND.n4534 GND.n4533 19.3944
R9684 GND.n4533 GND.n4532 19.3944
R9685 GND.n4532 GND.n3854 19.3944
R9686 GND.n4526 GND.n3854 19.3944
R9687 GND.n4526 GND.n4525 19.3944
R9688 GND.n4525 GND.n4524 19.3944
R9689 GND.n4524 GND.n3862 19.3944
R9690 GND.n4518 GND.n3862 19.3944
R9691 GND.n4518 GND.n4517 19.3944
R9692 GND.n4517 GND.n4516 19.3944
R9693 GND.n4516 GND.n3870 19.3944
R9694 GND.n4510 GND.n3870 19.3944
R9695 GND.n4510 GND.n4509 19.3944
R9696 GND.n4509 GND.n4508 19.3944
R9697 GND.n4508 GND.n3878 19.3944
R9698 GND.n4502 GND.n3878 19.3944
R9699 GND.n4502 GND.n4501 19.3944
R9700 GND.n4501 GND.n4500 19.3944
R9701 GND.n4500 GND.n3886 19.3944
R9702 GND.n4494 GND.n3886 19.3944
R9703 GND.n4494 GND.n4493 19.3944
R9704 GND.n4493 GND.n4492 19.3944
R9705 GND.n4492 GND.n3894 19.3944
R9706 GND.n4486 GND.n3894 19.3944
R9707 GND.n4486 GND.n4485 19.3944
R9708 GND.n4485 GND.n4484 19.3944
R9709 GND.n4484 GND.n3902 19.3944
R9710 GND.n4478 GND.n3902 19.3944
R9711 GND.n4478 GND.n4477 19.3944
R9712 GND.n4477 GND.n4476 19.3944
R9713 GND.n4476 GND.n3910 19.3944
R9714 GND.n4470 GND.n3910 19.3944
R9715 GND.n4470 GND.n4469 19.3944
R9716 GND.n4469 GND.n4468 19.3944
R9717 GND.n4468 GND.n3918 19.3944
R9718 GND.n4462 GND.n3918 19.3944
R9719 GND.n4462 GND.n4461 19.3944
R9720 GND.n4461 GND.n4460 19.3944
R9721 GND.n4460 GND.n3926 19.3944
R9722 GND.n4454 GND.n3926 19.3944
R9723 GND.n4454 GND.n4453 19.3944
R9724 GND.n4453 GND.n4452 19.3944
R9725 GND.n4452 GND.n3934 19.3944
R9726 GND.n4446 GND.n3934 19.3944
R9727 GND.n4446 GND.n4445 19.3944
R9728 GND.n4445 GND.n4444 19.3944
R9729 GND.n4444 GND.n3942 19.3944
R9730 GND.n4438 GND.n3942 19.3944
R9731 GND.n4438 GND.n4437 19.3944
R9732 GND.n4437 GND.n4436 19.3944
R9733 GND.n4436 GND.n3950 19.3944
R9734 GND.n4430 GND.n3950 19.3944
R9735 GND.n4430 GND.n4429 19.3944
R9736 GND.n4429 GND.n4428 19.3944
R9737 GND.n4428 GND.n3958 19.3944
R9738 GND.n4422 GND.n3958 19.3944
R9739 GND.n4422 GND.n4421 19.3944
R9740 GND.n4421 GND.n4420 19.3944
R9741 GND.n4420 GND.n3966 19.3944
R9742 GND.n4414 GND.n3966 19.3944
R9743 GND.n4414 GND.n4413 19.3944
R9744 GND.n4413 GND.n4412 19.3944
R9745 GND.n4412 GND.n3974 19.3944
R9746 GND.n4406 GND.n3974 19.3944
R9747 GND.n4406 GND.n4405 19.3944
R9748 GND.n4405 GND.n4404 19.3944
R9749 GND.n4404 GND.n3982 19.3944
R9750 GND.n4398 GND.n3982 19.3944
R9751 GND.n4398 GND.n4397 19.3944
R9752 GND.n4397 GND.n4396 19.3944
R9753 GND.n4396 GND.n3990 19.3944
R9754 GND.n4390 GND.n3990 19.3944
R9755 GND.n4390 GND.n4389 19.3944
R9756 GND.n4389 GND.n4388 19.3944
R9757 GND.n4388 GND.n3998 19.3944
R9758 GND.n4382 GND.n3998 19.3944
R9759 GND.n4382 GND.n4381 19.3944
R9760 GND.n4381 GND.n4380 19.3944
R9761 GND.n4380 GND.n4006 19.3944
R9762 GND.n4374 GND.n4006 19.3944
R9763 GND.n4374 GND.n4373 19.3944
R9764 GND.n4373 GND.n4372 19.3944
R9765 GND.n4372 GND.n4014 19.3944
R9766 GND.n4366 GND.n4014 19.3944
R9767 GND.n4366 GND.n4365 19.3944
R9768 GND.n4365 GND.n4364 19.3944
R9769 GND.n4364 GND.n4022 19.3944
R9770 GND.n4358 GND.n4022 19.3944
R9771 GND.n4358 GND.n4357 19.3944
R9772 GND.n4357 GND.n4356 19.3944
R9773 GND.n4356 GND.n4030 19.3944
R9774 GND.n4350 GND.n4030 19.3944
R9775 GND.n4350 GND.n4349 19.3944
R9776 GND.n4349 GND.n4348 19.3944
R9777 GND.n4348 GND.n4038 19.3944
R9778 GND.n4342 GND.n4038 19.3944
R9779 GND.n4342 GND.n4341 19.3944
R9780 GND.n4341 GND.n4340 19.3944
R9781 GND.n4340 GND.n4046 19.3944
R9782 GND.n4334 GND.n4046 19.3944
R9783 GND.n4334 GND.n4333 19.3944
R9784 GND.n4333 GND.n4332 19.3944
R9785 GND.n4332 GND.n4054 19.3944
R9786 GND.n4326 GND.n4054 19.3944
R9787 GND.n4326 GND.n4325 19.3944
R9788 GND.n4325 GND.n4324 19.3944
R9789 GND.n4324 GND.n4062 19.3944
R9790 GND.n4318 GND.n4062 19.3944
R9791 GND.n4318 GND.n4317 19.3944
R9792 GND.n4317 GND.n4316 19.3944
R9793 GND.n4316 GND.n4070 19.3944
R9794 GND.n4310 GND.n4070 19.3944
R9795 GND.n4310 GND.n4309 19.3944
R9796 GND.n4309 GND.n4308 19.3944
R9797 GND.n4302 GND.n4081 19.3944
R9798 GND.n4302 GND.n4082 19.3944
R9799 GND.n4298 GND.n4082 19.3944
R9800 GND.n4298 GND.n4085 19.3944
R9801 GND.n4292 GND.n4085 19.3944
R9802 GND.n4292 GND.n4291 19.3944
R9803 GND.n4291 GND.n4290 19.3944
R9804 GND.n4290 GND.n4092 19.3944
R9805 GND.n4284 GND.n4092 19.3944
R9806 GND.n4284 GND.n4283 19.3944
R9807 GND.n4283 GND.n4282 19.3944
R9808 GND.n4282 GND.n4100 19.3944
R9809 GND.n4276 GND.n4100 19.3944
R9810 GND.n4276 GND.n4275 19.3944
R9811 GND.n4275 GND.n4274 19.3944
R9812 GND.n4274 GND.n4108 19.3944
R9813 GND.n4268 GND.n4108 19.3944
R9814 GND.n4268 GND.n4267 19.3944
R9815 GND.n4267 GND.n4266 19.3944
R9816 GND.n4266 GND.n4116 19.3944
R9817 GND.n4260 GND.n4116 19.3944
R9818 GND.n4260 GND.n4259 19.3944
R9819 GND.n4259 GND.n4258 19.3944
R9820 GND.n4258 GND.n4124 19.3944
R9821 GND.n4252 GND.n4124 19.3944
R9822 GND.n4252 GND.n4251 19.3944
R9823 GND.n4251 GND.n4250 19.3944
R9824 GND.n4250 GND.n4132 19.3944
R9825 GND.n4244 GND.n4132 19.3944
R9826 GND.n4244 GND.n4243 19.3944
R9827 GND.n4243 GND.n4242 19.3944
R9828 GND.n4242 GND.n4140 19.3944
R9829 GND.n4236 GND.n4140 19.3944
R9830 GND.n4236 GND.n4235 19.3944
R9831 GND.n4235 GND.n4234 19.3944
R9832 GND.n4234 GND.n4148 19.3944
R9833 GND.n4228 GND.n4148 19.3944
R9834 GND.n4228 GND.n4227 19.3944
R9835 GND.n4227 GND.n4226 19.3944
R9836 GND.n4226 GND.n4156 19.3944
R9837 GND.n4220 GND.n4156 19.3944
R9838 GND.n4220 GND.n4219 19.3944
R9839 GND.n4219 GND.n4218 19.3944
R9840 GND.n4218 GND.n4164 19.3944
R9841 GND.n4212 GND.n4164 19.3944
R9842 GND.n4212 GND.n4211 19.3944
R9843 GND.n4211 GND.n4210 19.3944
R9844 GND.n4210 GND.n4172 19.3944
R9845 GND.n4204 GND.n4172 19.3944
R9846 GND.n4204 GND.n4203 19.3944
R9847 GND.n4203 GND.n4202 19.3944
R9848 GND.n4202 GND.n4180 19.3944
R9849 GND.n4196 GND.n4180 19.3944
R9850 GND.n4196 GND.n4195 19.3944
R9851 GND.n4195 GND.n4194 19.3944
R9852 GND.n4194 GND.n4190 19.3944
R9853 GND.n6722 GND.n6721 19.3944
R9854 GND.n6721 GND.n6720 19.3944
R9855 GND.n6720 GND.n6719 19.3944
R9856 GND.n6719 GND.n6717 19.3944
R9857 GND.n6717 GND.n6714 19.3944
R9858 GND.n6714 GND.n6713 19.3944
R9859 GND.n6713 GND.n6710 19.3944
R9860 GND.n6708 GND.n6705 19.3944
R9861 GND.n6705 GND.n6704 19.3944
R9862 GND.n6704 GND.n6701 19.3944
R9863 GND.n6701 GND.n6700 19.3944
R9864 GND.n6700 GND.n6697 19.3944
R9865 GND.n6697 GND.n6696 19.3944
R9866 GND.n6696 GND.n6693 19.3944
R9867 GND.n6693 GND.n6692 19.3944
R9868 GND.n6692 GND.n6689 19.3944
R9869 GND.n6736 GND.n924 19.3944
R9870 GND.n6750 GND.n924 19.3944
R9871 GND.n6750 GND.n6749 19.3944
R9872 GND.n6749 GND.n6748 19.3944
R9873 GND.n6748 GND.n6747 19.3944
R9874 GND.n6747 GND.n896 19.3944
R9875 GND.n6861 GND.n896 19.3944
R9876 GND.n6861 GND.n6860 19.3944
R9877 GND.n6860 GND.n6859 19.3944
R9878 GND.n6859 GND.n877 19.3944
R9879 GND.n6881 GND.n877 19.3944
R9880 GND.n6881 GND.n6880 19.3944
R9881 GND.n6880 GND.n6879 19.3944
R9882 GND.n6879 GND.n857 19.3944
R9883 GND.n6901 GND.n857 19.3944
R9884 GND.n6901 GND.n6900 19.3944
R9885 GND.n6900 GND.n6899 19.3944
R9886 GND.n6899 GND.n837 19.3944
R9887 GND.n6921 GND.n837 19.3944
R9888 GND.n6921 GND.n6920 19.3944
R9889 GND.n6920 GND.n6919 19.3944
R9890 GND.n6919 GND.n817 19.3944
R9891 GND.n6941 GND.n817 19.3944
R9892 GND.n6941 GND.n6940 19.3944
R9893 GND.n6940 GND.n6939 19.3944
R9894 GND.n6939 GND.n797 19.3944
R9895 GND.n6961 GND.n797 19.3944
R9896 GND.n6961 GND.n6960 19.3944
R9897 GND.n6960 GND.n6959 19.3944
R9898 GND.n6959 GND.n777 19.3944
R9899 GND.n6981 GND.n777 19.3944
R9900 GND.n6981 GND.n6980 19.3944
R9901 GND.n6980 GND.n6979 19.3944
R9902 GND.n6979 GND.n757 19.3944
R9903 GND.n7001 GND.n757 19.3944
R9904 GND.n7001 GND.n7000 19.3944
R9905 GND.n7000 GND.n6999 19.3944
R9906 GND.n6999 GND.n736 19.3944
R9907 GND.n7025 GND.n736 19.3944
R9908 GND.n7025 GND.n7024 19.3944
R9909 GND.n7024 GND.n7023 19.3944
R9910 GND.n7023 GND.n7022 19.3944
R9911 GND.n7022 GND.n708 19.3944
R9912 GND.n7069 GND.n708 19.3944
R9913 GND.n7069 GND.n7068 19.3944
R9914 GND.n7068 GND.n7067 19.3944
R9915 GND.n7067 GND.n688 19.3944
R9916 GND.n7097 GND.n688 19.3944
R9917 GND.n7097 GND.n7096 19.3944
R9918 GND.n7096 GND.n7095 19.3944
R9919 GND.n7095 GND.n661 19.3944
R9920 GND.n7133 GND.n661 19.3944
R9921 GND.n7133 GND.n7132 19.3944
R9922 GND.n7132 GND.n7131 19.3944
R9923 GND.n7131 GND.n666 19.3944
R9924 GND.n666 GND.n640 19.3944
R9925 GND.n7158 GND.n640 19.3944
R9926 GND.n7158 GND.n7157 19.3944
R9927 GND.n7157 GND.n627 19.3944
R9928 GND.n7171 GND.n627 19.3944
R9929 GND.n7172 GND.n7171 19.3944
R9930 GND.n7174 GND.n7172 19.3944
R9931 GND.n7174 GND.n623 19.3944
R9932 GND.n7203 GND.n623 19.3944
R9933 GND.n7203 GND.n258 19.3944
R9934 GND.n7630 GND.n258 19.3944
R9935 GND.n7630 GND.n7629 19.3944
R9936 GND.n7629 GND.n7628 19.3944
R9937 GND.n7628 GND.n262 19.3944
R9938 GND.n7618 GND.n262 19.3944
R9939 GND.n7618 GND.n7617 19.3944
R9940 GND.n7617 GND.n7616 19.3944
R9941 GND.n7616 GND.n283 19.3944
R9942 GND.n7606 GND.n283 19.3944
R9943 GND.n7606 GND.n7605 19.3944
R9944 GND.n7605 GND.n7604 19.3944
R9945 GND.n7604 GND.n304 19.3944
R9946 GND.n7347 GND.n304 19.3944
R9947 GND.n7349 GND.n7347 19.3944
R9948 GND.n7350 GND.n7349 19.3944
R9949 GND.n7353 GND.n7350 19.3944
R9950 GND.n7354 GND.n7353 19.3944
R9951 GND.n7356 GND.n7354 19.3944
R9952 GND.n7357 GND.n7356 19.3944
R9953 GND.n7360 GND.n7357 19.3944
R9954 GND.n7361 GND.n7360 19.3944
R9955 GND.n7363 GND.n7361 19.3944
R9956 GND.n7364 GND.n7363 19.3944
R9957 GND.n7367 GND.n7364 19.3944
R9958 GND.n7368 GND.n7367 19.3944
R9959 GND.n7370 GND.n7368 19.3944
R9960 GND.n7371 GND.n7370 19.3944
R9961 GND.n7374 GND.n7371 19.3944
R9962 GND.n7375 GND.n7374 19.3944
R9963 GND.n7377 GND.n7375 19.3944
R9964 GND.n7378 GND.n7377 19.3944
R9965 GND.n7381 GND.n7378 19.3944
R9966 GND.n7382 GND.n7381 19.3944
R9967 GND.n7384 GND.n7382 19.3944
R9968 GND.n7385 GND.n7384 19.3944
R9969 GND.n7388 GND.n7385 19.3944
R9970 GND.n7389 GND.n7388 19.3944
R9971 GND.n7391 GND.n7389 19.3944
R9972 GND.n7392 GND.n7391 19.3944
R9973 GND.n7395 GND.n7392 19.3944
R9974 GND.n7396 GND.n7395 19.3944
R9975 GND.n7398 GND.n7396 19.3944
R9976 GND.n7399 GND.n7398 19.3944
R9977 GND.n7402 GND.n7399 19.3944
R9978 GND.n7403 GND.n7402 19.3944
R9979 GND.n7405 GND.n7403 19.3944
R9980 GND.n7406 GND.n7405 19.3944
R9981 GND.n7409 GND.n7406 19.3944
R9982 GND.n7410 GND.n7409 19.3944
R9983 GND.n7412 GND.n7410 19.3944
R9984 GND.n7413 GND.n7412 19.3944
R9985 GND.n7416 GND.n7413 19.3944
R9986 GND.n7417 GND.n7416 19.3944
R9987 GND.n7419 GND.n7417 19.3944
R9988 GND.n7420 GND.n7419 19.3944
R9989 GND.n7421 GND.n7420 19.3944
R9990 GND.n6739 GND.n927 19.3944
R9991 GND.n6740 GND.n6739 19.3944
R9992 GND.n6742 GND.n6740 19.3944
R9993 GND.n6743 GND.n6742 19.3944
R9994 GND.n6743 GND.n898 19.3944
R9995 GND.n6854 GND.n898 19.3944
R9996 GND.n6855 GND.n6854 19.3944
R9997 GND.n6856 GND.n6855 19.3944
R9998 GND.n6856 GND.n879 19.3944
R9999 GND.n6874 GND.n879 19.3944
R10000 GND.n6875 GND.n6874 19.3944
R10001 GND.n6876 GND.n6875 19.3944
R10002 GND.n6876 GND.n859 19.3944
R10003 GND.n6894 GND.n859 19.3944
R10004 GND.n6895 GND.n6894 19.3944
R10005 GND.n6896 GND.n6895 19.3944
R10006 GND.n6896 GND.n839 19.3944
R10007 GND.n6914 GND.n839 19.3944
R10008 GND.n6915 GND.n6914 19.3944
R10009 GND.n6916 GND.n6915 19.3944
R10010 GND.n6916 GND.n819 19.3944
R10011 GND.n6934 GND.n819 19.3944
R10012 GND.n6935 GND.n6934 19.3944
R10013 GND.n6936 GND.n6935 19.3944
R10014 GND.n6936 GND.n799 19.3944
R10015 GND.n6954 GND.n799 19.3944
R10016 GND.n6955 GND.n6954 19.3944
R10017 GND.n6956 GND.n6955 19.3944
R10018 GND.n6956 GND.n779 19.3944
R10019 GND.n6974 GND.n779 19.3944
R10020 GND.n6975 GND.n6974 19.3944
R10021 GND.n6976 GND.n6975 19.3944
R10022 GND.n6976 GND.n759 19.3944
R10023 GND.n6994 GND.n759 19.3944
R10024 GND.n6995 GND.n6994 19.3944
R10025 GND.n6996 GND.n6995 19.3944
R10026 GND.n6996 GND.n739 19.3944
R10027 GND.n7014 GND.n739 19.3944
R10028 GND.n7015 GND.n7014 19.3944
R10029 GND.n7017 GND.n7015 19.3944
R10030 GND.n7018 GND.n7017 19.3944
R10031 GND.n7018 GND.n710 19.3944
R10032 GND.n7062 GND.n710 19.3944
R10033 GND.n7063 GND.n7062 19.3944
R10034 GND.n7064 GND.n7063 19.3944
R10035 GND.n7064 GND.n691 19.3944
R10036 GND.n7082 GND.n691 19.3944
R10037 GND.n7083 GND.n7082 19.3944
R10038 GND.n7085 GND.n7083 19.3944
R10039 GND.n7086 GND.n7085 19.3944
R10040 GND.n7092 GND.n7086 19.3944
R10041 GND.n7092 GND.n7090 19.3944
R10042 GND.n7090 GND.n7089 19.3944
R10043 GND.n7089 GND.n7087 19.3944
R10044 GND.n7087 GND.n642 19.3944
R10045 GND.n7148 GND.n642 19.3944
R10046 GND.n7149 GND.n7148 19.3944
R10047 GND.n7151 GND.n7149 19.3944
R10048 GND.n7154 GND.n7151 19.3944
R10049 GND.n7154 GND.n7153 19.3944
R10050 GND.n7153 GND.n625 19.3944
R10051 GND.n7176 GND.n625 19.3944
R10052 GND.n7179 GND.n7176 19.3944
R10053 GND.n7180 GND.n7179 19.3944
R10054 GND.n7200 GND.n7180 19.3944
R10055 GND.n7200 GND.n7198 19.3944
R10056 GND.n7198 GND.n7197 19.3944
R10057 GND.n7197 GND.n7195 19.3944
R10058 GND.n7195 GND.n7194 19.3944
R10059 GND.n7194 GND.n7192 19.3944
R10060 GND.n7192 GND.n7191 19.3944
R10061 GND.n7191 GND.n7189 19.3944
R10062 GND.n7189 GND.n7188 19.3944
R10063 GND.n7188 GND.n7186 19.3944
R10064 GND.n7186 GND.n7185 19.3944
R10065 GND.n7185 GND.n7183 19.3944
R10066 GND.n7183 GND.n322 19.3944
R10067 GND.n7594 GND.n322 19.3944
R10068 GND.n7594 GND.n7593 19.3944
R10069 GND.n7593 GND.n7592 19.3944
R10070 GND.n7592 GND.n327 19.3944
R10071 GND.n7582 GND.n327 19.3944
R10072 GND.n7582 GND.n7581 19.3944
R10073 GND.n7581 GND.n7580 19.3944
R10074 GND.n7580 GND.n346 19.3944
R10075 GND.n7570 GND.n346 19.3944
R10076 GND.n7570 GND.n7569 19.3944
R10077 GND.n7569 GND.n7568 19.3944
R10078 GND.n7568 GND.n365 19.3944
R10079 GND.n7558 GND.n365 19.3944
R10080 GND.n7558 GND.n7557 19.3944
R10081 GND.n7557 GND.n7556 19.3944
R10082 GND.n7556 GND.n384 19.3944
R10083 GND.n7546 GND.n384 19.3944
R10084 GND.n7546 GND.n7545 19.3944
R10085 GND.n7545 GND.n7544 19.3944
R10086 GND.n7544 GND.n403 19.3944
R10087 GND.n7534 GND.n403 19.3944
R10088 GND.n7534 GND.n7533 19.3944
R10089 GND.n7533 GND.n7532 19.3944
R10090 GND.n7532 GND.n422 19.3944
R10091 GND.n7522 GND.n422 19.3944
R10092 GND.n7522 GND.n7521 19.3944
R10093 GND.n7521 GND.n7520 19.3944
R10094 GND.n7520 GND.n441 19.3944
R10095 GND.n7510 GND.n441 19.3944
R10096 GND.n7510 GND.n7509 19.3944
R10097 GND.n7509 GND.n7508 19.3944
R10098 GND.n7508 GND.n461 19.3944
R10099 GND.n7498 GND.n461 19.3944
R10100 GND.n7498 GND.n7497 19.3944
R10101 GND.n7497 GND.n7496 19.3944
R10102 GND.n7496 GND.n480 19.3944
R10103 GND.n7486 GND.n480 19.3944
R10104 GND.n7486 GND.n7485 19.3944
R10105 GND.n7485 GND.n7484 19.3944
R10106 GND.n7484 GND.n498 19.3944
R10107 GND.n7474 GND.n498 19.3944
R10108 GND.n7474 GND.n7473 19.3944
R10109 GND.n7473 GND.n7472 19.3944
R10110 GND.n7472 GND.n518 19.3944
R10111 GND.n7444 GND.n541 19.3944
R10112 GND.n7444 GND.n547 19.3944
R10113 GND.n7439 GND.n547 19.3944
R10114 GND.n7439 GND.n7438 19.3944
R10115 GND.n7438 GND.n7437 19.3944
R10116 GND.n7437 GND.n554 19.3944
R10117 GND.n7432 GND.n554 19.3944
R10118 GND.n7432 GND.n7431 19.3944
R10119 GND.n7431 GND.n7430 19.3944
R10120 GND.n7464 GND.n527 19.3944
R10121 GND.n529 GND.n527 19.3944
R10122 GND.n7457 GND.n529 19.3944
R10123 GND.n7457 GND.n7456 19.3944
R10124 GND.n7456 GND.n7455 19.3944
R10125 GND.n7455 GND.n535 19.3944
R10126 GND.n7450 GND.n535 19.3944
R10127 GND.n7450 GND.n7449 19.3944
R10128 GND.n7345 GND.n568 19.3944
R10129 GND.n7340 GND.n568 19.3944
R10130 GND.n7340 GND.n7339 19.3944
R10131 GND.n7339 GND.n7338 19.3944
R10132 GND.n7338 GND.n573 19.3944
R10133 GND.n7333 GND.n573 19.3944
R10134 GND.n7333 GND.n7332 19.3944
R10135 GND.n7332 GND.n7331 19.3944
R10136 GND.n1376 GND.n1375 19.3944
R10137 GND.n1375 GND.n1374 19.3944
R10138 GND.n1374 GND.n906 19.3944
R10139 GND.n6764 GND.n906 19.3944
R10140 GND.n6764 GND.n904 19.3944
R10141 GND.n6850 GND.n904 19.3944
R10142 GND.n6850 GND.n6849 19.3944
R10143 GND.n6849 GND.n6848 19.3944
R10144 GND.n6848 GND.n6846 19.3944
R10145 GND.n6846 GND.n6845 19.3944
R10146 GND.n6845 GND.n6843 19.3944
R10147 GND.n6843 GND.n6842 19.3944
R10148 GND.n6842 GND.n6840 19.3944
R10149 GND.n6840 GND.n6839 19.3944
R10150 GND.n6839 GND.n6837 19.3944
R10151 GND.n6837 GND.n6836 19.3944
R10152 GND.n6836 GND.n6834 19.3944
R10153 GND.n6834 GND.n6833 19.3944
R10154 GND.n6833 GND.n6831 19.3944
R10155 GND.n6831 GND.n6830 19.3944
R10156 GND.n6830 GND.n6828 19.3944
R10157 GND.n6828 GND.n6827 19.3944
R10158 GND.n6827 GND.n6825 19.3944
R10159 GND.n6825 GND.n6824 19.3944
R10160 GND.n6824 GND.n6822 19.3944
R10161 GND.n6822 GND.n6821 19.3944
R10162 GND.n6821 GND.n6819 19.3944
R10163 GND.n6819 GND.n6818 19.3944
R10164 GND.n6818 GND.n6816 19.3944
R10165 GND.n6816 GND.n6815 19.3944
R10166 GND.n6815 GND.n6813 19.3944
R10167 GND.n6813 GND.n6812 19.3944
R10168 GND.n6812 GND.n6810 19.3944
R10169 GND.n6810 GND.n6809 19.3944
R10170 GND.n6809 GND.n6807 19.3944
R10171 GND.n6807 GND.n6806 19.3944
R10172 GND.n6806 GND.n6804 19.3944
R10173 GND.n6804 GND.n6803 19.3944
R10174 GND.n6803 GND.n6801 19.3944
R10175 GND.n6801 GND.n718 19.3944
R10176 GND.n7039 GND.n718 19.3944
R10177 GND.n7039 GND.n716 19.3944
R10178 GND.n7058 GND.n716 19.3944
R10179 GND.n7058 GND.n7057 19.3944
R10180 GND.n7057 GND.n7056 19.3944
R10181 GND.n7056 GND.n7054 19.3944
R10182 GND.n7054 GND.n7053 19.3944
R10183 GND.n7053 GND.n7051 19.3944
R10184 GND.n7051 GND.n7050 19.3944
R10185 GND.n7050 GND.n671 19.3944
R10186 GND.n7110 GND.n671 19.3944
R10187 GND.n7111 GND.n7110 19.3944
R10188 GND.n7111 GND.n669 19.3944
R10189 GND.n7127 GND.n669 19.3944
R10190 GND.n7127 GND.n7126 19.3944
R10191 GND.n7126 GND.n7125 19.3944
R10192 GND.n7125 GND.n7123 19.3944
R10193 GND.n7123 GND.n7122 19.3944
R10194 GND.n7122 GND.n7120 19.3944
R10195 GND.n7120 GND.n229 19.3944
R10196 GND.n7643 GND.n229 19.3944
R10197 GND.n7643 GND.n230 19.3944
R10198 GND.n617 GND.n230 19.3944
R10199 GND.n617 GND.n615 19.3944
R10200 GND.n7211 GND.n615 19.3944
R10201 GND.n7211 GND.n613 19.3944
R10202 GND.n7216 GND.n613 19.3944
R10203 GND.n7217 GND.n7216 19.3944
R10204 GND.n7219 GND.n7217 19.3944
R10205 GND.n7219 GND.n611 19.3944
R10206 GND.n7224 GND.n611 19.3944
R10207 GND.n7225 GND.n7224 19.3944
R10208 GND.n7227 GND.n7225 19.3944
R10209 GND.n7227 GND.n609 19.3944
R10210 GND.n7232 GND.n609 19.3944
R10211 GND.n7233 GND.n7232 19.3944
R10212 GND.n7236 GND.n7233 19.3944
R10213 GND.n7236 GND.n607 19.3944
R10214 GND.n7241 GND.n607 19.3944
R10215 GND.n7242 GND.n7241 19.3944
R10216 GND.n7244 GND.n7242 19.3944
R10217 GND.n7244 GND.n605 19.3944
R10218 GND.n7249 GND.n605 19.3944
R10219 GND.n7250 GND.n7249 19.3944
R10220 GND.n7252 GND.n7250 19.3944
R10221 GND.n7252 GND.n603 19.3944
R10222 GND.n7257 GND.n603 19.3944
R10223 GND.n7258 GND.n7257 19.3944
R10224 GND.n7260 GND.n7258 19.3944
R10225 GND.n7260 GND.n601 19.3944
R10226 GND.n7265 GND.n601 19.3944
R10227 GND.n7266 GND.n7265 19.3944
R10228 GND.n7268 GND.n7266 19.3944
R10229 GND.n7268 GND.n599 19.3944
R10230 GND.n7273 GND.n599 19.3944
R10231 GND.n7274 GND.n7273 19.3944
R10232 GND.n7276 GND.n7274 19.3944
R10233 GND.n7276 GND.n597 19.3944
R10234 GND.n7281 GND.n597 19.3944
R10235 GND.n7282 GND.n7281 19.3944
R10236 GND.n7284 GND.n7282 19.3944
R10237 GND.n7284 GND.n595 19.3944
R10238 GND.n7289 GND.n595 19.3944
R10239 GND.n7290 GND.n7289 19.3944
R10240 GND.n7292 GND.n7290 19.3944
R10241 GND.n7292 GND.n593 19.3944
R10242 GND.n7297 GND.n593 19.3944
R10243 GND.n7298 GND.n7297 19.3944
R10244 GND.n7300 GND.n7298 19.3944
R10245 GND.n7300 GND.n591 19.3944
R10246 GND.n7305 GND.n591 19.3944
R10247 GND.n7306 GND.n7305 19.3944
R10248 GND.n7308 GND.n7306 19.3944
R10249 GND.n7308 GND.n589 19.3944
R10250 GND.n7313 GND.n589 19.3944
R10251 GND.n7314 GND.n7313 19.3944
R10252 GND.n7316 GND.n7314 19.3944
R10253 GND.n7316 GND.n587 19.3944
R10254 GND.n7321 GND.n587 19.3944
R10255 GND.n7322 GND.n7321 19.3944
R10256 GND.n7323 GND.n7322 19.3944
R10257 GND.n1350 GND.n1347 19.3944
R10258 GND.n1355 GND.n1352 19.3944
R10259 GND.n1360 GND.n1357 19.3944
R10260 GND.n1365 GND.n1360 19.3944
R10261 GND.n1137 GND.n1136 19.3944
R10262 GND.n1136 GND.n1134 19.3944
R10263 GND.n1134 GND.n1133 19.3944
R10264 GND.n1133 GND.n1131 19.3944
R10265 GND.n1131 GND.n1130 19.3944
R10266 GND.n1130 GND.n1128 19.3944
R10267 GND.n1128 GND.n1127 19.3944
R10268 GND.n1127 GND.n1126 19.3944
R10269 GND.n1126 GND.n1124 19.3944
R10270 GND.n1124 GND.n1123 19.3944
R10271 GND.n1123 GND.n1121 19.3944
R10272 GND.n1121 GND.n1120 19.3944
R10273 GND.n1120 GND.n1118 19.3944
R10274 GND.n1118 GND.n1117 19.3944
R10275 GND.n1117 GND.n1115 19.3944
R10276 GND.n1115 GND.n1114 19.3944
R10277 GND.n1114 GND.n1112 19.3944
R10278 GND.n1112 GND.n1111 19.3944
R10279 GND.n1111 GND.n1109 19.3944
R10280 GND.n1109 GND.n1108 19.3944
R10281 GND.n1108 GND.n1106 19.3944
R10282 GND.n1106 GND.n1105 19.3944
R10283 GND.n1105 GND.n1103 19.3944
R10284 GND.n1103 GND.n1102 19.3944
R10285 GND.n1102 GND.n1100 19.3944
R10286 GND.n1100 GND.n1099 19.3944
R10287 GND.n1099 GND.n1097 19.3944
R10288 GND.n1097 GND.n1096 19.3944
R10289 GND.n1096 GND.n1094 19.3944
R10290 GND.n1094 GND.n1093 19.3944
R10291 GND.n1093 GND.n1091 19.3944
R10292 GND.n1091 GND.n1090 19.3944
R10293 GND.n1090 GND.n1088 19.3944
R10294 GND.n1088 GND.n1087 19.3944
R10295 GND.n1087 GND.n1085 19.3944
R10296 GND.n1085 GND.n1084 19.3944
R10297 GND.n1084 GND.n1082 19.3944
R10298 GND.n1082 GND.n1081 19.3944
R10299 GND.n1081 GND.n1079 19.3944
R10300 GND.n1079 GND.n1078 19.3944
R10301 GND.n1078 GND.n1076 19.3944
R10302 GND.n1076 GND.n1075 19.3944
R10303 GND.n1075 GND.n1073 19.3944
R10304 GND.n1073 GND.n1072 19.3944
R10305 GND.n1072 GND.n1071 19.3944
R10306 GND.n1071 GND.n1069 19.3944
R10307 GND.n1069 GND.n1068 19.3944
R10308 GND.n1068 GND.n1066 19.3944
R10309 GND.n1066 GND.n1065 19.3944
R10310 GND.n1065 GND.n1063 19.3944
R10311 GND.n1063 GND.n1062 19.3944
R10312 GND.n1062 GND.n1060 19.3944
R10313 GND.n1060 GND.n1059 19.3944
R10314 GND.n1059 GND.n1057 19.3944
R10315 GND.n1057 GND.n1056 19.3944
R10316 GND.n1056 GND.n1055 19.3944
R10317 GND.n1053 GND.n1052 19.3944
R10318 GND.n1052 GND.n1050 19.3944
R10319 GND.n1048 GND.n1046 19.3944
R10320 GND.n1044 GND.n1041 19.3944
R10321 GND.n1039 GND.n1038 19.3944
R10322 GND.n1038 GND.n1036 19.3944
R10323 GND.n1036 GND.n1035 19.3944
R10324 GND.n1035 GND.n1033 19.3944
R10325 GND.n1033 GND.n1032 19.3944
R10326 GND.n1032 GND.n1030 19.3944
R10327 GND.n1030 GND.n1029 19.3944
R10328 GND.n1029 GND.n1027 19.3944
R10329 GND.n1027 GND.n1026 19.3944
R10330 GND.n1026 GND.n1024 19.3944
R10331 GND.n1024 GND.n311 19.3944
R10332 GND.n7600 GND.n311 19.3944
R10333 GND.n7600 GND.n7599 19.3944
R10334 GND.n7599 GND.n7598 19.3944
R10335 GND.n7598 GND.n315 19.3944
R10336 GND.n7588 GND.n315 19.3944
R10337 GND.n7588 GND.n7587 19.3944
R10338 GND.n7587 GND.n7586 19.3944
R10339 GND.n7586 GND.n337 19.3944
R10340 GND.n7576 GND.n337 19.3944
R10341 GND.n7576 GND.n7575 19.3944
R10342 GND.n7575 GND.n7574 19.3944
R10343 GND.n7574 GND.n356 19.3944
R10344 GND.n7564 GND.n356 19.3944
R10345 GND.n7564 GND.n7563 19.3944
R10346 GND.n7563 GND.n7562 19.3944
R10347 GND.n7562 GND.n375 19.3944
R10348 GND.n7552 GND.n375 19.3944
R10349 GND.n7552 GND.n7551 19.3944
R10350 GND.n7551 GND.n7550 19.3944
R10351 GND.n7550 GND.n394 19.3944
R10352 GND.n7540 GND.n394 19.3944
R10353 GND.n7540 GND.n7539 19.3944
R10354 GND.n7539 GND.n7538 19.3944
R10355 GND.n7538 GND.n413 19.3944
R10356 GND.n7528 GND.n413 19.3944
R10357 GND.n7528 GND.n7527 19.3944
R10358 GND.n7527 GND.n7526 19.3944
R10359 GND.n7526 GND.n431 19.3944
R10360 GND.n7516 GND.n431 19.3944
R10361 GND.n7516 GND.n7515 19.3944
R10362 GND.n7515 GND.n7514 19.3944
R10363 GND.n7514 GND.n451 19.3944
R10364 GND.n7504 GND.n451 19.3944
R10365 GND.n7504 GND.n7503 19.3944
R10366 GND.n7503 GND.n7502 19.3944
R10367 GND.n7502 GND.n471 19.3944
R10368 GND.n7492 GND.n471 19.3944
R10369 GND.n7492 GND.n7491 19.3944
R10370 GND.n7491 GND.n7490 19.3944
R10371 GND.n7490 GND.n490 19.3944
R10372 GND.n7480 GND.n490 19.3944
R10373 GND.n7480 GND.n7479 19.3944
R10374 GND.n7479 GND.n7478 19.3944
R10375 GND.n7478 GND.n509 19.3944
R10376 GND.n7468 GND.n509 19.3944
R10377 GND.n7468 GND.n7467 19.3944
R10378 GND.n5032 GND.n2769 19.3944
R10379 GND.n5052 GND.n2769 19.3944
R10380 GND.n5052 GND.n2767 19.3944
R10381 GND.n5056 GND.n2767 19.3944
R10382 GND.n5056 GND.n2537 19.3944
R10383 GND.n5212 GND.n2537 19.3944
R10384 GND.n5212 GND.n2535 19.3944
R10385 GND.n5216 GND.n2535 19.3944
R10386 GND.n5218 GND.n5216 19.3944
R10387 GND.n5218 GND.n5217 19.3944
R10388 GND.n2734 GND.n2516 19.3944
R10389 GND.n5077 GND.n2516 19.3944
R10390 GND.n5080 GND.n5079 19.3944
R10391 GND.n5178 GND.n5177 19.3944
R10392 GND.n5180 GND.n2511 19.3944
R10393 GND.n5227 GND.n2511 19.3944
R10394 GND.n5227 GND.n2493 19.3944
R10395 GND.n5243 GND.n2493 19.3944
R10396 GND.n5243 GND.n2491 19.3944
R10397 GND.n5247 GND.n2491 19.3944
R10398 GND.n5247 GND.n2473 19.3944
R10399 GND.n5263 GND.n2473 19.3944
R10400 GND.n5263 GND.n2471 19.3944
R10401 GND.n5267 GND.n2471 19.3944
R10402 GND.n5267 GND.n2452 19.3944
R10403 GND.n5283 GND.n2452 19.3944
R10404 GND.n5283 GND.n2450 19.3944
R10405 GND.n5287 GND.n2450 19.3944
R10406 GND.n5287 GND.n2433 19.3944
R10407 GND.n5303 GND.n2433 19.3944
R10408 GND.n5303 GND.n2431 19.3944
R10409 GND.n5307 GND.n2431 19.3944
R10410 GND.n5307 GND.n2413 19.3944
R10411 GND.n5323 GND.n2413 19.3944
R10412 GND.n5323 GND.n2411 19.3944
R10413 GND.n5327 GND.n2411 19.3944
R10414 GND.n5327 GND.n2392 19.3944
R10415 GND.n5343 GND.n2392 19.3944
R10416 GND.n5343 GND.n2390 19.3944
R10417 GND.n5347 GND.n2390 19.3944
R10418 GND.n5347 GND.n2373 19.3944
R10419 GND.n5363 GND.n2373 19.3944
R10420 GND.n5363 GND.n2371 19.3944
R10421 GND.n5367 GND.n2371 19.3944
R10422 GND.n5367 GND.n2353 19.3944
R10423 GND.n5388 GND.n2353 19.3944
R10424 GND.n5388 GND.n2351 19.3944
R10425 GND.n5394 GND.n2351 19.3944
R10426 GND.n5394 GND.n5393 19.3944
R10427 GND.n5393 GND.n2326 19.3944
R10428 GND.n5468 GND.n2326 19.3944
R10429 GND.n5468 GND.n2324 19.3944
R10430 GND.n5472 GND.n2324 19.3944
R10431 GND.n5472 GND.n2306 19.3944
R10432 GND.n5488 GND.n2306 19.3944
R10433 GND.n5488 GND.n2304 19.3944
R10434 GND.n5492 GND.n2304 19.3944
R10435 GND.n5492 GND.n2286 19.3944
R10436 GND.n5508 GND.n2286 19.3944
R10437 GND.n5508 GND.n2284 19.3944
R10438 GND.n5512 GND.n2284 19.3944
R10439 GND.n5512 GND.n2265 19.3944
R10440 GND.n5528 GND.n2265 19.3944
R10441 GND.n5528 GND.n2263 19.3944
R10442 GND.n5532 GND.n2263 19.3944
R10443 GND.n5532 GND.n2246 19.3944
R10444 GND.n5552 GND.n2246 19.3944
R10445 GND.n5552 GND.n2244 19.3944
R10446 GND.n5557 GND.n2244 19.3944
R10447 GND.n5557 GND.n1744 19.3944
R10448 GND.n5689 GND.n1744 19.3944
R10449 GND.n5689 GND.n5688 19.3944
R10450 GND.n5688 GND.n5687 19.3944
R10451 GND.n5687 GND.n1748 19.3944
R10452 GND.n5681 GND.n1748 19.3944
R10453 GND.n5681 GND.n5680 19.3944
R10454 GND.n5680 GND.n5679 19.3944
R10455 GND.n5679 GND.n1784 19.3944
R10456 GND.n2179 GND.n1784 19.3944
R10457 GND.n2179 GND.n2178 19.3944
R10458 GND.n2178 GND.n2177 19.3944
R10459 GND.n2177 GND.n1830 19.3944
R10460 GND.n2165 GND.n1830 19.3944
R10461 GND.n2165 GND.n2164 19.3944
R10462 GND.n2164 GND.n2163 19.3944
R10463 GND.n2163 GND.n1848 19.3944
R10464 GND.n2151 GND.n1848 19.3944
R10465 GND.n2151 GND.n2150 19.3944
R10466 GND.n2150 GND.n2149 19.3944
R10467 GND.n2149 GND.n1866 19.3944
R10468 GND.n2137 GND.n1866 19.3944
R10469 GND.n2137 GND.n2136 19.3944
R10470 GND.n2136 GND.n2135 19.3944
R10471 GND.n2135 GND.n1884 19.3944
R10472 GND.n2123 GND.n1884 19.3944
R10473 GND.n2123 GND.n2122 19.3944
R10474 GND.n2122 GND.n2121 19.3944
R10475 GND.n2121 GND.n1903 19.3944
R10476 GND.n2109 GND.n1903 19.3944
R10477 GND.n2109 GND.n2108 19.3944
R10478 GND.n2108 GND.n2107 19.3944
R10479 GND.n2107 GND.n1921 19.3944
R10480 GND.n2095 GND.n1921 19.3944
R10481 GND.n2095 GND.n2094 19.3944
R10482 GND.n2094 GND.n2093 19.3944
R10483 GND.n2093 GND.n1939 19.3944
R10484 GND.n2081 GND.n1939 19.3944
R10485 GND.n2081 GND.n2080 19.3944
R10486 GND.n2080 GND.n2079 19.3944
R10487 GND.n2079 GND.n1957 19.3944
R10488 GND.n1963 GND.n1957 19.3944
R10489 GND.n1963 GND.n1962 19.3944
R10490 GND.n1962 GND.n1700 19.3944
R10491 GND.n5785 GND.n1700 19.3944
R10492 GND.n5785 GND.n1698 19.3944
R10493 GND.n5806 GND.n1698 19.3944
R10494 GND.n5806 GND.n5805 19.3944
R10495 GND.n5805 GND.n5804 19.3944
R10496 GND.n5804 GND.n5791 19.3944
R10497 GND.n5800 GND.n5791 19.3944
R10498 GND.n5800 GND.n5799 19.3944
R10499 GND.n5799 GND.n5798 19.3944
R10500 GND.n5798 GND.n1618 19.3944
R10501 GND.n1618 GND.n1616 19.3944
R10502 GND.n5910 GND.n1616 19.3944
R10503 GND.n5910 GND.n1614 19.3944
R10504 GND.n5914 GND.n1614 19.3944
R10505 GND.n5914 GND.n1560 19.3944
R10506 GND.n5988 GND.n1560 19.3944
R10507 GND.n5988 GND.n1558 19.3944
R10508 GND.n6003 GND.n1558 19.3944
R10509 GND.n6003 GND.n6002 19.3944
R10510 GND.n6002 GND.n6001 19.3944
R10511 GND.n6001 GND.n5994 19.3944
R10512 GND.n5997 GND.n5994 19.3944
R10513 GND.n5997 GND.n1516 19.3944
R10514 GND.n6078 GND.n1516 19.3944
R10515 GND.n6078 GND.n1514 19.3944
R10516 GND.n6084 GND.n1514 19.3944
R10517 GND.n6084 GND.n6083 19.3944
R10518 GND.n6083 GND.n1481 19.3944
R10519 GND.n6144 GND.n1481 19.3944
R10520 GND.n6144 GND.n1479 19.3944
R10521 GND.n6148 GND.n1479 19.3944
R10522 GND.n6148 GND.n1457 19.3944
R10523 GND.n6187 GND.n1457 19.3944
R10524 GND.n6187 GND.n1455 19.3944
R10525 GND.n6193 GND.n1455 19.3944
R10526 GND.n6193 GND.n6192 19.3944
R10527 GND.n6192 GND.n1441 19.3944
R10528 GND.n6247 GND.n1441 19.3944
R10529 GND.n6247 GND.n1439 19.3944
R10530 GND.n6251 GND.n1439 19.3944
R10531 GND.n6251 GND.n1329 19.3944
R10532 GND.n6319 GND.n1329 19.3944
R10533 GND.n6319 GND.n1327 19.3944
R10534 GND.n6328 GND.n1327 19.3944
R10535 GND.n6328 GND.n6327 19.3944
R10536 GND.n6327 GND.n6326 19.3944
R10537 GND.n6326 GND.n1306 19.3944
R10538 GND.n6359 GND.n1306 19.3944
R10539 GND.n6359 GND.n1304 19.3944
R10540 GND.n6374 GND.n1304 19.3944
R10541 GND.n6374 GND.n6373 19.3944
R10542 GND.n6373 GND.n6372 19.3944
R10543 GND.n6372 GND.n6365 19.3944
R10544 GND.n6368 GND.n6365 19.3944
R10545 GND.n6368 GND.n1272 19.3944
R10546 GND.n6417 GND.n1272 19.3944
R10547 GND.n6417 GND.n1270 19.3944
R10548 GND.n6423 GND.n1270 19.3944
R10549 GND.n6423 GND.n6422 19.3944
R10550 GND.n6422 GND.n1247 19.3944
R10551 GND.n6452 GND.n1247 19.3944
R10552 GND.n6452 GND.n1245 19.3944
R10553 GND.n6461 GND.n1245 19.3944
R10554 GND.n6461 GND.n6460 19.3944
R10555 GND.n6460 GND.n6459 19.3944
R10556 GND.n6459 GND.n1222 19.3944
R10557 GND.n6491 GND.n1222 19.3944
R10558 GND.n6491 GND.n1220 19.3944
R10559 GND.n6506 GND.n1220 19.3944
R10560 GND.n6506 GND.n6505 19.3944
R10561 GND.n6505 GND.n6504 19.3944
R10562 GND.n6504 GND.n6497 19.3944
R10563 GND.n6500 GND.n6497 19.3944
R10564 GND.n6500 GND.n1188 19.3944
R10565 GND.n6596 GND.n1188 19.3944
R10566 GND.n6596 GND.n1186 19.3944
R10567 GND.n6614 GND.n1186 19.3944
R10568 GND.n6614 GND.n6613 19.3944
R10569 GND.n6613 GND.n6612 19.3944
R10570 GND.n6612 GND.n6602 19.3944
R10571 GND.n6606 GND.n6602 19.3944
R10572 GND.n6606 GND.n938 19.3944
R10573 GND.n6728 GND.n938 19.3944
R10574 GND.n6728 GND.n936 19.3944
R10575 GND.n6732 GND.n936 19.3944
R10576 GND.n6732 GND.n916 19.3944
R10577 GND.n6754 GND.n916 19.3944
R10578 GND.n6754 GND.n914 19.3944
R10579 GND.n6760 GND.n914 19.3944
R10580 GND.n6760 GND.n6759 19.3944
R10581 GND.n6759 GND.n889 19.3944
R10582 GND.n6865 GND.n889 19.3944
R10583 GND.n6865 GND.n887 19.3944
R10584 GND.n6869 GND.n887 19.3944
R10585 GND.n6869 GND.n869 19.3944
R10586 GND.n6885 GND.n869 19.3944
R10587 GND.n6885 GND.n867 19.3944
R10588 GND.n6889 GND.n867 19.3944
R10589 GND.n6889 GND.n849 19.3944
R10590 GND.n6905 GND.n849 19.3944
R10591 GND.n6905 GND.n847 19.3944
R10592 GND.n6909 GND.n847 19.3944
R10593 GND.n6909 GND.n828 19.3944
R10594 GND.n6925 GND.n828 19.3944
R10595 GND.n6925 GND.n826 19.3944
R10596 GND.n6929 GND.n826 19.3944
R10597 GND.n6929 GND.n809 19.3944
R10598 GND.n6945 GND.n809 19.3944
R10599 GND.n6945 GND.n807 19.3944
R10600 GND.n6949 GND.n807 19.3944
R10601 GND.n6949 GND.n789 19.3944
R10602 GND.n6965 GND.n789 19.3944
R10603 GND.n6965 GND.n787 19.3944
R10604 GND.n6969 GND.n787 19.3944
R10605 GND.n6969 GND.n769 19.3944
R10606 GND.n6985 GND.n769 19.3944
R10607 GND.n6985 GND.n767 19.3944
R10608 GND.n6989 GND.n767 19.3944
R10609 GND.n6989 GND.n749 19.3944
R10610 GND.n7005 GND.n749 19.3944
R10611 GND.n7005 GND.n747 19.3944
R10612 GND.n7009 GND.n747 19.3944
R10613 GND.n7009 GND.n728 19.3944
R10614 GND.n7029 GND.n728 19.3944
R10615 GND.n7029 GND.n726 19.3944
R10616 GND.n7035 GND.n726 19.3944
R10617 GND.n7035 GND.n7034 19.3944
R10618 GND.n7034 GND.n701 19.3944
R10619 GND.n7073 GND.n701 19.3944
R10620 GND.n7073 GND.n699 19.3944
R10621 GND.n7077 GND.n699 19.3944
R10622 GND.n7077 GND.n680 19.3944
R10623 GND.n7101 GND.n680 19.3944
R10624 GND.n7101 GND.n678 19.3944
R10625 GND.n7105 GND.n678 19.3944
R10626 GND.n7105 GND.n651 19.3944
R10627 GND.n7137 GND.n651 19.3944
R10628 GND.n7137 GND.n649 19.3944
R10629 GND.n7141 GND.n649 19.3944
R10630 GND.n7143 GND.n7141 19.3944
R10631 GND.n7143 GND.n7142 19.3944
R10632 GND.n7163 GND.n7162 19.3944
R10633 GND.n7166 GND.n7165 19.3944
R10634 GND.n7639 GND.n7638 19.3944
R10635 GND.n7206 GND.n241 19.3944
R10636 GND.n7634 GND.n248 19.3944
R10637 GND.n7634 GND.n249 19.3944
R10638 GND.n7624 GND.n249 19.3944
R10639 GND.n7624 GND.n7623 19.3944
R10640 GND.n7623 GND.n7622 19.3944
R10641 GND.n7622 GND.n273 19.3944
R10642 GND.n7612 GND.n273 19.3944
R10643 GND.n7612 GND.n7611 19.3944
R10644 GND.n7611 GND.n7610 19.3944
R10645 GND.n7610 GND.n294 19.3944
R10646 GND.n3180 GND.n3179 19.3944
R10647 GND.n3179 GND.n3055 19.3944
R10648 GND.n3174 GND.n3055 19.3944
R10649 GND.n3174 GND.n3173 19.3944
R10650 GND.n3173 GND.n3060 19.3944
R10651 GND.n3168 GND.n3060 19.3944
R10652 GND.n3168 GND.n3167 19.3944
R10653 GND.n3167 GND.n3166 19.3944
R10654 GND.n3160 GND.n3159 19.3944
R10655 GND.n3159 GND.n3158 19.3944
R10656 GND.n3158 GND.n3074 19.3944
R10657 GND.n3152 GND.n3074 19.3944
R10658 GND.n3152 GND.n3151 19.3944
R10659 GND.n3151 GND.n3150 19.3944
R10660 GND.n3150 GND.n3080 19.3944
R10661 GND.n3144 GND.n3080 19.3944
R10662 GND.n3144 GND.n3143 19.3944
R10663 GND.n3183 GND.n3037 19.3944
R10664 GND.n3203 GND.n3037 19.3944
R10665 GND.n3203 GND.n3035 19.3944
R10666 GND.n3209 GND.n3035 19.3944
R10667 GND.n3209 GND.n3208 19.3944
R10668 GND.n3208 GND.n3009 19.3944
R10669 GND.n3335 GND.n3009 19.3944
R10670 GND.n3335 GND.n3007 19.3944
R10671 GND.n3339 GND.n3007 19.3944
R10672 GND.n3339 GND.n2988 19.3944
R10673 GND.n3352 GND.n2988 19.3944
R10674 GND.n3352 GND.n2986 19.3944
R10675 GND.n3356 GND.n2986 19.3944
R10676 GND.n3356 GND.n2967 19.3944
R10677 GND.n3369 GND.n2967 19.3944
R10678 GND.n3369 GND.n2965 19.3944
R10679 GND.n3373 GND.n2965 19.3944
R10680 GND.n3373 GND.n2945 19.3944
R10681 GND.n3386 GND.n2945 19.3944
R10682 GND.n3386 GND.n2943 19.3944
R10683 GND.n3390 GND.n2943 19.3944
R10684 GND.n3390 GND.n2925 19.3944
R10685 GND.n3403 GND.n2925 19.3944
R10686 GND.n3403 GND.n2923 19.3944
R10687 GND.n3407 GND.n2923 19.3944
R10688 GND.n3407 GND.n2904 19.3944
R10689 GND.n3420 GND.n2904 19.3944
R10690 GND.n3420 GND.n2902 19.3944
R10691 GND.n3424 GND.n2902 19.3944
R10692 GND.n3424 GND.n2883 19.3944
R10693 GND.n3437 GND.n2883 19.3944
R10694 GND.n3437 GND.n2881 19.3944
R10695 GND.n3441 GND.n2881 19.3944
R10696 GND.n3441 GND.n2862 19.3944
R10697 GND.n3454 GND.n2862 19.3944
R10698 GND.n3454 GND.n2860 19.3944
R10699 GND.n3458 GND.n2860 19.3944
R10700 GND.n3458 GND.n2841 19.3944
R10701 GND.n3471 GND.n2841 19.3944
R10702 GND.n3471 GND.n2839 19.3944
R10703 GND.n3475 GND.n2839 19.3944
R10704 GND.n3475 GND.n2822 19.3944
R10705 GND.n3494 GND.n2822 19.3944
R10706 GND.n3494 GND.n2820 19.3944
R10707 GND.n3518 GND.n2820 19.3944
R10708 GND.n3518 GND.n3517 19.3944
R10709 GND.n3517 GND.n3516 19.3944
R10710 GND.n3516 GND.n3514 19.3944
R10711 GND.n3514 GND.n3513 19.3944
R10712 GND.n3513 GND.n3511 19.3944
R10713 GND.n3511 GND.n3510 19.3944
R10714 GND.n3510 GND.n3508 19.3944
R10715 GND.n3508 GND.n3507 19.3944
R10716 GND.n3507 GND.n2525 19.3944
R10717 GND.n5222 GND.n2525 19.3944
R10718 GND.n5222 GND.n2526 19.3944
R10719 GND.n2743 GND.n2742 19.3944
R10720 GND.n2740 GND.n2739 19.3944
R10721 GND.n2729 GND.n2728 19.3944
R10722 GND.n2717 GND.n2716 19.3944
R10723 GND.n2709 GND.n2708 19.3944
R10724 GND.n2708 GND.n2707 19.3944
R10725 GND.n2707 GND.n2705 19.3944
R10726 GND.n2705 GND.n2704 19.3944
R10727 GND.n2704 GND.n2702 19.3944
R10728 GND.n2702 GND.n2701 19.3944
R10729 GND.n2701 GND.n2699 19.3944
R10730 GND.n2699 GND.n2698 19.3944
R10731 GND.n2698 GND.n2696 19.3944
R10732 GND.n2696 GND.n2695 19.3944
R10733 GND.n2695 GND.n2693 19.3944
R10734 GND.n2693 GND.n2692 19.3944
R10735 GND.n2692 GND.n2690 19.3944
R10736 GND.n2690 GND.n2689 19.3944
R10737 GND.n2689 GND.n2687 19.3944
R10738 GND.n2687 GND.n2686 19.3944
R10739 GND.n2686 GND.n2684 19.3944
R10740 GND.n2684 GND.n2683 19.3944
R10741 GND.n2683 GND.n2681 19.3944
R10742 GND.n2681 GND.n2680 19.3944
R10743 GND.n2680 GND.n2678 19.3944
R10744 GND.n2678 GND.n2677 19.3944
R10745 GND.n2677 GND.n2675 19.3944
R10746 GND.n2675 GND.n2674 19.3944
R10747 GND.n2674 GND.n2672 19.3944
R10748 GND.n2672 GND.n2671 19.3944
R10749 GND.n2671 GND.n2669 19.3944
R10750 GND.n2669 GND.n2668 19.3944
R10751 GND.n2668 GND.n2666 19.3944
R10752 GND.n2666 GND.n2665 19.3944
R10753 GND.n2665 GND.n2663 19.3944
R10754 GND.n2663 GND.n2662 19.3944
R10755 GND.n2662 GND.n2660 19.3944
R10756 GND.n2660 GND.n2659 19.3944
R10757 GND.n2659 GND.n2657 19.3944
R10758 GND.n2657 GND.n2656 19.3944
R10759 GND.n2656 GND.n2655 19.3944
R10760 GND.n2655 GND.n2653 19.3944
R10761 GND.n2653 GND.n2652 19.3944
R10762 GND.n2652 GND.n2650 19.3944
R10763 GND.n2650 GND.n2649 19.3944
R10764 GND.n2649 GND.n2647 19.3944
R10765 GND.n2647 GND.n2646 19.3944
R10766 GND.n2646 GND.n2644 19.3944
R10767 GND.n2644 GND.n2643 19.3944
R10768 GND.n2643 GND.n2641 19.3944
R10769 GND.n2641 GND.n2640 19.3944
R10770 GND.n2640 GND.n2638 19.3944
R10771 GND.n2638 GND.n2637 19.3944
R10772 GND.n2637 GND.n2635 19.3944
R10773 GND.n2635 GND.n2634 19.3944
R10774 GND.n2634 GND.n2632 19.3944
R10775 GND.n2632 GND.n2631 19.3944
R10776 GND.n2631 GND.n2237 19.3944
R10777 GND.n5562 GND.n2237 19.3944
R10778 GND.n5563 GND.n5562 19.3944
R10779 GND.n3111 GND.n3110 19.3944
R10780 GND.n3110 GND.n3109 19.3944
R10781 GND.n3109 GND.n3028 19.3944
R10782 GND.n3213 GND.n3028 19.3944
R10783 GND.n3213 GND.n3025 19.3944
R10784 GND.n3323 GND.n3025 19.3944
R10785 GND.n3323 GND.n3026 19.3944
R10786 GND.n3319 GND.n3026 19.3944
R10787 GND.n3319 GND.n3318 19.3944
R10788 GND.n3318 GND.n3317 19.3944
R10789 GND.n3317 GND.n3219 19.3944
R10790 GND.n3313 GND.n3219 19.3944
R10791 GND.n3313 GND.n3312 19.3944
R10792 GND.n3312 GND.n3311 19.3944
R10793 GND.n3311 GND.n3223 19.3944
R10794 GND.n3307 GND.n3223 19.3944
R10795 GND.n3307 GND.n3306 19.3944
R10796 GND.n3306 GND.n3305 19.3944
R10797 GND.n3305 GND.n3227 19.3944
R10798 GND.n3301 GND.n3227 19.3944
R10799 GND.n3301 GND.n3300 19.3944
R10800 GND.n3300 GND.n3299 19.3944
R10801 GND.n3299 GND.n3231 19.3944
R10802 GND.n3295 GND.n3231 19.3944
R10803 GND.n3295 GND.n3294 19.3944
R10804 GND.n3294 GND.n3293 19.3944
R10805 GND.n3293 GND.n3235 19.3944
R10806 GND.n3289 GND.n3235 19.3944
R10807 GND.n3289 GND.n3288 19.3944
R10808 GND.n3288 GND.n3287 19.3944
R10809 GND.n3287 GND.n3239 19.3944
R10810 GND.n3283 GND.n3239 19.3944
R10811 GND.n3283 GND.n3282 19.3944
R10812 GND.n3282 GND.n3281 19.3944
R10813 GND.n3281 GND.n3243 19.3944
R10814 GND.n3277 GND.n3243 19.3944
R10815 GND.n3277 GND.n3276 19.3944
R10816 GND.n3276 GND.n3275 19.3944
R10817 GND.n3275 GND.n3247 19.3944
R10818 GND.n3271 GND.n3247 19.3944
R10819 GND.n3271 GND.n3270 19.3944
R10820 GND.n3270 GND.n3269 19.3944
R10821 GND.n3269 GND.n3251 19.3944
R10822 GND.n3265 GND.n3251 19.3944
R10823 GND.n3265 GND.n3264 19.3944
R10824 GND.n3264 GND.n3263 19.3944
R10825 GND.n3263 GND.n3255 19.3944
R10826 GND.n3259 GND.n3255 19.3944
R10827 GND.n3259 GND.n3258 19.3944
R10828 GND.n3258 GND.n2760 19.3944
R10829 GND.n5061 GND.n2760 19.3944
R10830 GND.n5062 GND.n5061 19.3944
R10831 GND.n5062 GND.n2753 19.3944
R10832 GND.n5066 GND.n2753 19.3944
R10833 GND.n5067 GND.n5066 19.3944
R10834 GND.n5069 GND.n5067 19.3944
R10835 GND.n5069 GND.n2751 19.3944
R10836 GND.n5073 GND.n2751 19.3944
R10837 GND.n5073 GND.n2725 19.3944
R10838 GND.n5084 GND.n2725 19.3944
R10839 GND.n5084 GND.n2723 19.3944
R10840 GND.n5173 GND.n2723 19.3944
R10841 GND.n5173 GND.n5172 19.3944
R10842 GND.n5172 GND.n5171 19.3944
R10843 GND.n5171 GND.n5170 19.3944
R10844 GND.n5170 GND.n5168 19.3944
R10845 GND.n5168 GND.n5167 19.3944
R10846 GND.n5167 GND.n5165 19.3944
R10847 GND.n5165 GND.n5164 19.3944
R10848 GND.n5164 GND.n5162 19.3944
R10849 GND.n5162 GND.n5161 19.3944
R10850 GND.n5161 GND.n5159 19.3944
R10851 GND.n5159 GND.n5158 19.3944
R10852 GND.n5158 GND.n5156 19.3944
R10853 GND.n5156 GND.n5155 19.3944
R10854 GND.n5155 GND.n5153 19.3944
R10855 GND.n5153 GND.n5152 19.3944
R10856 GND.n5152 GND.n5150 19.3944
R10857 GND.n5150 GND.n5149 19.3944
R10858 GND.n5149 GND.n5147 19.3944
R10859 GND.n5147 GND.n5146 19.3944
R10860 GND.n5146 GND.n5144 19.3944
R10861 GND.n5144 GND.n5143 19.3944
R10862 GND.n5143 GND.n5141 19.3944
R10863 GND.n5141 GND.n5140 19.3944
R10864 GND.n5140 GND.n5138 19.3944
R10865 GND.n5138 GND.n5137 19.3944
R10866 GND.n5137 GND.n5135 19.3944
R10867 GND.n5135 GND.n5134 19.3944
R10868 GND.n5134 GND.n5132 19.3944
R10869 GND.n5132 GND.n5131 19.3944
R10870 GND.n5131 GND.n5129 19.3944
R10871 GND.n5129 GND.n5128 19.3944
R10872 GND.n5128 GND.n5126 19.3944
R10873 GND.n5126 GND.n5125 19.3944
R10874 GND.n5125 GND.n5123 19.3944
R10875 GND.n5123 GND.n2343 19.3944
R10876 GND.n5398 GND.n2343 19.3944
R10877 GND.n5398 GND.n2341 19.3944
R10878 GND.n5453 GND.n2341 19.3944
R10879 GND.n5453 GND.n5452 19.3944
R10880 GND.n5452 GND.n5451 19.3944
R10881 GND.n5451 GND.n5449 19.3944
R10882 GND.n5449 GND.n5448 19.3944
R10883 GND.n5448 GND.n5446 19.3944
R10884 GND.n5446 GND.n5445 19.3944
R10885 GND.n5445 GND.n5443 19.3944
R10886 GND.n5443 GND.n5442 19.3944
R10887 GND.n5442 GND.n5440 19.3944
R10888 GND.n5440 GND.n5439 19.3944
R10889 GND.n5439 GND.n5437 19.3944
R10890 GND.n5437 GND.n5436 19.3944
R10891 GND.n5436 GND.n5434 19.3944
R10892 GND.n5434 GND.n5433 19.3944
R10893 GND.n5433 GND.n5431 19.3944
R10894 GND.n5431 GND.n5430 19.3944
R10895 GND.n5430 GND.n5428 19.3944
R10896 GND.n5428 GND.n5427 19.3944
R10897 GND.n5427 GND.n5425 19.3944
R10898 GND.n5425 GND.n5424 19.3944
R10899 GND.n5424 GND.n5422 19.3944
R10900 GND.n3136 GND.n3092 19.3944
R10901 GND.n3131 GND.n3092 19.3944
R10902 GND.n3131 GND.n3094 19.3944
R10903 GND.n3127 GND.n3094 19.3944
R10904 GND.n3127 GND.n3126 19.3944
R10905 GND.n3126 GND.n3125 19.3944
R10906 GND.n3125 GND.n3101 19.3944
R10907 GND.n3121 GND.n3101 19.3944
R10908 GND.n3089 GND.n3044 19.3944
R10909 GND.n3199 GND.n3044 19.3944
R10910 GND.n3199 GND.n3045 19.3944
R10911 GND.n3190 GND.n3045 19.3944
R10912 GND.n3192 GND.n3190 19.3944
R10913 GND.n3192 GND.n3015 19.3944
R10914 GND.n3331 GND.n3015 19.3944
R10915 GND.n3331 GND.n3016 19.3944
R10916 GND.n3018 GND.n3016 19.3944
R10917 GND.n3018 GND.n2995 19.3944
R10918 GND.n3348 GND.n2995 19.3944
R10919 GND.n3348 GND.n2996 19.3944
R10920 GND.n2998 GND.n2996 19.3944
R10921 GND.n2998 GND.n2974 19.3944
R10922 GND.n3365 GND.n2974 19.3944
R10923 GND.n3365 GND.n2975 19.3944
R10924 GND.n2977 GND.n2975 19.3944
R10925 GND.n2977 GND.n2953 19.3944
R10926 GND.n3382 GND.n2953 19.3944
R10927 GND.n3382 GND.n2954 19.3944
R10928 GND.n2956 GND.n2954 19.3944
R10929 GND.n2956 GND.n2932 19.3944
R10930 GND.n3399 GND.n2932 19.3944
R10931 GND.n3399 GND.n2933 19.3944
R10932 GND.n2935 GND.n2933 19.3944
R10933 GND.n2935 GND.n2911 19.3944
R10934 GND.n3416 GND.n2911 19.3944
R10935 GND.n3416 GND.n2912 19.3944
R10936 GND.n2914 GND.n2912 19.3944
R10937 GND.n2914 GND.n2890 19.3944
R10938 GND.n3433 GND.n2890 19.3944
R10939 GND.n3433 GND.n2891 19.3944
R10940 GND.n2893 GND.n2891 19.3944
R10941 GND.n2893 GND.n2869 19.3944
R10942 GND.n3450 GND.n2869 19.3944
R10943 GND.n3450 GND.n2870 19.3944
R10944 GND.n2872 GND.n2870 19.3944
R10945 GND.n2872 GND.n2848 19.3944
R10946 GND.n3467 GND.n2848 19.3944
R10947 GND.n3467 GND.n2849 19.3944
R10948 GND.n2851 GND.n2849 19.3944
R10949 GND.n2851 GND.n2829 19.3944
R10950 GND.n3490 GND.n2829 19.3944
R10951 GND.n3490 GND.n2830 19.3944
R10952 GND.n3482 GND.n2830 19.3944
R10953 GND.n3482 GND.n2780 19.3944
R10954 GND.n5037 GND.n2780 19.3944
R10955 GND.n5038 GND.n5037 19.3944
R10956 GND.n5040 GND.n5038 19.3944
R10957 GND.n5043 GND.n5040 19.3944
R10958 GND.n5043 GND.n5042 19.3944
R10959 GND.n5042 GND.n2550 19.3944
R10960 GND.n2551 GND.n2550 19.3944
R10961 GND.n2552 GND.n2551 19.3944
R10962 GND.n2557 GND.n2552 19.3944
R10963 GND.n2558 GND.n2557 19.3944
R10964 GND.n2559 GND.n2558 19.3944
R10965 GND.n2560 GND.n2559 19.3944
R10966 GND.n2747 GND.n2560 19.3944
R10967 GND.n2747 GND.n2566 19.3944
R10968 GND.n2567 GND.n2566 19.3944
R10969 GND.n2568 GND.n2567 19.3944
R10970 GND.n2575 GND.n2568 19.3944
R10971 GND.n5184 GND.n2575 19.3944
R10972 GND.n5185 GND.n5184 19.3944
R10973 GND.n5185 GND.n2504 19.3944
R10974 GND.n5232 GND.n2504 19.3944
R10975 GND.n5233 GND.n5232 19.3944
R10976 GND.n5234 GND.n5233 19.3944
R10977 GND.n5234 GND.n2484 19.3944
R10978 GND.n5252 GND.n2484 19.3944
R10979 GND.n5253 GND.n5252 19.3944
R10980 GND.n5254 GND.n5253 19.3944
R10981 GND.n5254 GND.n2464 19.3944
R10982 GND.n5272 GND.n2464 19.3944
R10983 GND.n5273 GND.n5272 19.3944
R10984 GND.n5274 GND.n5273 19.3944
R10985 GND.n5274 GND.n2444 19.3944
R10986 GND.n5292 GND.n2444 19.3944
R10987 GND.n5293 GND.n5292 19.3944
R10988 GND.n5294 GND.n5293 19.3944
R10989 GND.n5294 GND.n2424 19.3944
R10990 GND.n5312 GND.n2424 19.3944
R10991 GND.n5313 GND.n5312 19.3944
R10992 GND.n5314 GND.n5313 19.3944
R10993 GND.n5314 GND.n2404 19.3944
R10994 GND.n5332 GND.n2404 19.3944
R10995 GND.n5333 GND.n5332 19.3944
R10996 GND.n5334 GND.n5333 19.3944
R10997 GND.n5334 GND.n2384 19.3944
R10998 GND.n5352 GND.n2384 19.3944
R10999 GND.n5353 GND.n5352 19.3944
R11000 GND.n5354 GND.n5353 19.3944
R11001 GND.n5354 GND.n2364 19.3944
R11002 GND.n5372 GND.n2364 19.3944
R11003 GND.n5373 GND.n5372 19.3944
R11004 GND.n5375 GND.n5373 19.3944
R11005 GND.n5376 GND.n5375 19.3944
R11006 GND.n5376 GND.n2336 19.3944
R11007 GND.n5457 GND.n2336 19.3944
R11008 GND.n5458 GND.n5457 19.3944
R11009 GND.n5459 GND.n5458 19.3944
R11010 GND.n5459 GND.n2317 19.3944
R11011 GND.n5477 GND.n2317 19.3944
R11012 GND.n5478 GND.n5477 19.3944
R11013 GND.n5479 GND.n5478 19.3944
R11014 GND.n5479 GND.n2297 19.3944
R11015 GND.n5497 GND.n2297 19.3944
R11016 GND.n5498 GND.n5497 19.3944
R11017 GND.n5499 GND.n5498 19.3944
R11018 GND.n5499 GND.n2277 19.3944
R11019 GND.n5517 GND.n2277 19.3944
R11020 GND.n5518 GND.n5517 19.3944
R11021 GND.n5519 GND.n5518 19.3944
R11022 GND.n5519 GND.n2257 19.3944
R11023 GND.n5537 GND.n2257 19.3944
R11024 GND.n5538 GND.n5537 19.3944
R11025 GND.n5540 GND.n5538 19.3944
R11026 GND.n5543 GND.n5540 19.3944
R11027 GND.n5543 GND.n5542 19.3944
R11028 GND.n5542 GND.n1733 19.3944
R11029 GND.n6310 GND.n6309 19.3944
R11030 GND.n6309 GND.n6308 19.3944
R11031 GND.n6308 GND.n1344 19.3944
R11032 GND.n6303 GND.n1344 19.3944
R11033 GND.n6303 GND.n6302 19.3944
R11034 GND.n6302 GND.n6301 19.3944
R11035 GND.n6301 GND.n1386 19.3944
R11036 GND.n6297 GND.n1386 19.3944
R11037 GND.n6297 GND.n6296 19.3944
R11038 GND.n6296 GND.n6295 19.3944
R11039 GND.n6295 GND.n1394 19.3944
R11040 GND.n6291 GND.n1394 19.3944
R11041 GND.n6291 GND.n6290 19.3944
R11042 GND.n6290 GND.n6289 19.3944
R11043 GND.n6289 GND.n1402 19.3944
R11044 GND.n6285 GND.n1402 19.3944
R11045 GND.n6283 GND.n6282 19.3944
R11046 GND.n6282 GND.n1412 19.3944
R11047 GND.n6278 GND.n1412 19.3944
R11048 GND.n5821 GND.n1679 19.3944
R11049 GND.n5826 GND.n1679 19.3944
R11050 GND.n5826 GND.n1680 19.3944
R11051 GND.n1680 GND.n1653 19.3944
R11052 GND.n5855 GND.n1653 19.3944
R11053 GND.n5855 GND.n1651 19.3944
R11054 GND.n5859 GND.n1651 19.3944
R11055 GND.n5859 GND.n1625 19.3944
R11056 GND.n5899 GND.n1625 19.3944
R11057 GND.n5899 GND.n1623 19.3944
R11058 GND.n5903 GND.n1623 19.3944
R11059 GND.n5903 GND.n1583 19.3944
R11060 GND.n5940 GND.n1583 19.3944
R11061 GND.n5940 GND.n1580 19.3944
R11062 GND.n5945 GND.n1580 19.3944
R11063 GND.n5945 GND.n1581 19.3944
R11064 GND.n1581 GND.n1551 19.3944
R11065 GND.n6008 GND.n1551 19.3944
R11066 GND.n6008 GND.n1549 19.3944
R11067 GND.n6012 GND.n1549 19.3944
R11068 GND.n6012 GND.n1532 19.3944
R11069 GND.n6060 GND.n1532 19.3944
R11070 GND.n6060 GND.n1529 19.3944
R11071 GND.n6065 GND.n1529 19.3944
R11072 GND.n6065 GND.n1530 19.3944
R11073 GND.n1530 GND.n1500 19.3944
R11074 GND.n6099 GND.n1500 19.3944
R11075 GND.n6099 GND.n1498 19.3944
R11076 GND.n6103 GND.n1498 19.3944
R11077 GND.n6103 GND.n1473 19.3944
R11078 GND.n6153 GND.n1473 19.3944
R11079 GND.n6153 GND.n1470 19.3944
R11080 GND.n6167 GND.n1470 19.3944
R11081 GND.n6167 GND.n1471 19.3944
R11082 GND.n6163 GND.n1471 19.3944
R11083 GND.n6163 GND.n6162 19.3944
R11084 GND.n6162 GND.n6161 19.3944
R11085 GND.n6161 GND.n1425 19.3944
R11086 GND.n6262 GND.n1425 19.3944
R11087 GND.n6262 GND.n1423 19.3944
R11088 GND.n6266 GND.n1423 19.3944
R11089 GND.n6266 GND.n1336 19.3944
R11090 GND.n6314 GND.n1336 19.3944
R11091 GND.n6314 GND.n1337 19.3944
R11092 GND.n5034 GND.n2782 19.2044
R11093 GND.n2167 GND.n1842 19.2044
R11094 GND.n1990 GND.n1842 19.2044
R11095 GND.n2037 GND.n1923 19.2044
R11096 GND.n2105 GND.n1923 19.2044
R11097 GND.n5783 GND.n5782 19.2044
R11098 GND.n5853 GND.n1655 19.2044
R11099 GND.n5853 GND.n1658 19.2044
R11100 GND.n5861 GND.n1648 19.2044
R11101 GND.n5897 GND.n1627 19.2044
R11102 GND.n5938 GND.n1585 19.2044
R11103 GND.n5917 GND.n5916 19.2044
R11104 GND.n5986 GND.n1562 19.2044
R11105 GND.n6014 GND.n1541 19.2044
R11106 GND.n6058 GND.n1534 19.2044
R11107 GND.n6058 GND.n1537 19.2044
R11108 GND.n6068 GND.n6067 19.2044
R11109 GND.n6028 GND.n1505 19.2044
R11110 GND.n6142 GND.n6141 19.2044
R11111 GND.n6151 GND.n6150 19.2044
R11112 GND.n6195 GND.n1453 19.2044
R11113 GND.n6244 GND.n1443 19.2044
R11114 GND.n6260 GND.n1427 19.2044
R11115 GND.n6260 GND.n1430 19.2044
R11116 GND.n6317 GND.n6316 19.2044
R11117 GND.n6407 GND.n1274 19.2044
R11118 GND.n6415 GND.n1274 19.2044
R11119 GND.n6528 GND.n1201 19.2044
R11120 GND.n6528 GND.n1202 19.2044
R11121 GND.n5925 GND.n5924 18.4363
R11122 GND.n5947 GND.n1576 18.4363
R11123 GND.n6105 GND.n1483 18.4363
R11124 GND.n6132 GND.n1477 18.4363
R11125 GND.n2175 GND.n2174 17.6681
R11126 GND.n2098 GND.n2097 17.6681
R11127 GND.n5810 GND.n1694 17.6681
R11128 GND.n1649 GND.n1635 17.6681
R11129 GND.n6015 GND.n1546 17.6681
R11130 GND.n6076 GND.n1518 17.6681
R11131 GND.n6236 GND.n6235 17.6681
R11132 GND.n6212 GND.n1421 17.6681
R11133 GND.n6396 GND.n1285 17.6681
R11134 GND.n6594 GND.n1190 17.6681
R11135 GND.n5677 GND.n5676 17.284
R11136 GND.t76 GND.n1807 16.8999
R11137 GND.n5819 GND.n1683 16.8999
R11138 GND.n5878 GND.n1619 16.8999
R11139 GND.n5985 GND.n1564 16.8999
R11140 GND.n6097 GND.n6096 16.8999
R11141 GND.n6184 GND.n1460 16.8999
R11142 GND.n6331 GND.n1321 16.8999
R11143 GND.n3333 GND.t34 16.5525
R11144 GND.n2181 GND.n1824 16.1318
R11145 GND.n2160 GND.t16 16.1318
R11146 GND.n2003 GND.n1860 16.1318
R11147 GND.n2024 GND.n1905 16.1318
R11148 GND.n2091 GND.n1941 16.1318
R11149 GND.n5781 GND.n1686 16.1318
R11150 GND.n5896 GND.n1630 16.1318
R11151 GND.n1604 GND.n1553 16.1318
R11152 GND.n6087 GND.n6086 16.1318
R11153 GND.n6178 GND.n6177 16.1318
R11154 GND.n6205 GND.n1333 16.1318
R11155 GND.n1296 GND.n1295 16.1318
R11156 GND.n1261 GND.n1255 16.1318
R11157 GND.n6509 GND.n1216 16.1318
R11158 GND.t24 GND.n1211 16.1318
R11159 GND.n6617 GND.n6616 16.1318
R11160 GND.n7448 GND.n541 16.0975
R11161 GND.n3160 GND.n3068 16.0975
R11162 GND.n5673 GND.n1816 15.6103
R11163 GND.n6662 GND.n6621 15.6103
R11164 GND.n2397 GND.t88 15.3636
R11165 GND.t84 GND.n1966 15.3636
R11166 GND.n5828 GND.n1675 15.3636
R11167 GND.n5886 GND.n5885 15.3636
R11168 GND.n5976 GND.n1555 15.3636
R11169 GND.n6037 GND.n1520 15.3636
R11170 GND.n6196 GND.n1449 15.3636
R11171 GND.n6213 GND.n1331 15.3636
R11172 GND.n6348 GND.t6 15.3636
R11173 GND.t117 GND.n762 15.3636
R11174 GND.t108 GND.n369 15.3636
R11175 GND.n5613 GND.n5605 15.3217
R11176 GND.n6689 GND.n6684 15.3217
R11177 GND.n7430 GND.n563 15.3217
R11178 GND.n3143 GND.n3088 15.3217
R11179 GND.n2146 GND.n1870 14.5955
R11180 GND.n2126 GND.n1895 14.5955
R11181 GND.n2084 GND.n2083 14.5955
R11182 GND.n5770 GND.n1705 14.5955
R11183 GND.n1621 GND.n1593 14.5955
R11184 GND.t82 GND.n1598 14.5955
R11185 GND.t1 GND.n6029 14.5955
R11186 GND.n6170 GND.n1466 14.5955
R11187 GND.n1325 GND.n1323 14.5955
R11188 GND.n6377 GND.n1300 14.5955
R11189 GND.n6449 GND.n1251 14.5955
R11190 GND.n6481 GND.n1224 14.5955
R11191 GND.n5906 GND.t5 14.2114
R11192 GND.n6185 GND.t85 14.2114
R11193 GND.n3435 GND.t105 14.1879
R11194 GND.n7331 GND.n582 14.1581
R11195 GND.n1369 GND.n1368 14.1581
R11196 GND.n3121 GND.n3120 14.1581
R11197 GND.n5838 GND.n1668 13.8273
R11198 GND.n5847 GND.n1662 13.8273
R11199 GND.n6052 GND.n6051 13.8273
R11200 GND.n6069 GND.n1524 13.8273
R11201 GND.n6243 GND.n1445 13.8273
R11202 GND.n6254 GND.n1436 13.8273
R11203 GND.n1815 GND.n1812 13.1884
R11204 GND.n1179 GND.n1176 13.1884
R11205 GND.n5685 GND.n1777 13.0592
R11206 GND.n1886 GND.n1878 13.0592
R11207 GND.n1887 GND.n1886 13.0592
R11208 GND.n2077 GND.n1966 13.0592
R11209 GND.n2077 GND.n2076 13.0592
R11210 GND.n5937 GND.n1588 13.0592
R11211 GND.n5918 GND.n1588 13.0592
R11212 GND.n6140 GND.n1486 13.0592
R11213 GND.n1486 GND.n1475 13.0592
R11214 GND.n6350 GND.n6349 13.0592
R11215 GND.n6349 GND.n6348 13.0592
R11216 GND.n1242 GND.n1235 13.0592
R11217 GND.n6470 GND.n1235 13.0592
R11218 GND.n6726 GND.n6725 13.0592
R11219 GND.n5839 GND.n5838 12.291
R11220 GND.n6051 GND.n6050 12.291
R11221 GND.n6044 GND.n1524 12.291
R11222 GND.n6225 GND.n1436 12.291
R11223 GND.n1758 GND.n1730 11.8308
R11224 GND.n7326 GND.n582 11.8308
R11225 GND.n3120 GND.n3114 11.8308
R11226 GND.n3520 GND.n2782 11.8234
R11227 GND.n5534 GND.t9 11.5228
R11228 GND.n2182 GND.t76 11.5228
R11229 GND.n1876 GND.n1870 11.5228
R11230 GND.n1895 GND.n1889 11.5228
R11231 GND.n2083 GND.n1951 11.5228
R11232 GND.n5926 GND.n1593 11.5228
R11233 GND.n1598 GND.n1577 11.5228
R11234 GND.n6029 GND.n1496 11.5228
R11235 GND.n6133 GND.n1466 11.5228
R11236 GND.n1309 GND.n1300 11.5228
R11237 GND.n1251 GND.n1240 11.5228
R11238 GND.n6482 GND.n6481 11.5228
R11239 GND.n6610 GND.t42 11.5228
R11240 GND.n6852 GND.t45 11.5228
R11241 GND.n500 GND.t20 11.5228
R11242 GND.n6006 GND.t2 11.1388
R11243 GND.t83 GND.n1510 11.1388
R11244 GND.n5220 GND.t86 10.7547
R11245 GND.n5229 GND.t112 10.7547
R11246 GND.n5828 GND.n1676 10.7547
R11247 GND.n5887 GND.n5886 10.7547
R11248 GND.n5977 GND.n5976 10.7547
R11249 GND.n6075 GND.n1520 10.7547
R11250 GND.n6237 GND.n1449 10.7547
R11251 GND.n6220 GND.n6213 10.7547
R11252 GND.n7145 GND.t100 10.7547
R11253 GND.n7632 GND.t122 10.7547
R11254 GND.n5613 GND.n5612 10.6672
R11255 GND.n6685 GND.n6684 10.6672
R11256 GND.n7425 GND.n563 10.6672
R11257 GND.n3139 GND.n3088 10.6672
R11258 GND.n6537 GND.n1147 10.6151
R11259 GND.n6538 GND.n6537 10.6151
R11260 GND.n6542 GND.n6541 10.6151
R11261 GND.n6545 GND.n6542 10.6151
R11262 GND.n6546 GND.n6545 10.6151
R11263 GND.n6549 GND.n6546 10.6151
R11264 GND.n6550 GND.n6549 10.6151
R11265 GND.n6553 GND.n6550 10.6151
R11266 GND.n6554 GND.n6553 10.6151
R11267 GND.n6557 GND.n6554 10.6151
R11268 GND.n6558 GND.n6557 10.6151
R11269 GND.n6561 GND.n6558 10.6151
R11270 GND.n6562 GND.n6561 10.6151
R11271 GND.n6565 GND.n6562 10.6151
R11272 GND.n6566 GND.n6565 10.6151
R11273 GND.n6569 GND.n6566 10.6151
R11274 GND.n6570 GND.n6569 10.6151
R11275 GND.n6573 GND.n6570 10.6151
R11276 GND.n6574 GND.n6573 10.6151
R11277 GND.n1973 GND.n1822 10.6151
R11278 GND.n1974 GND.n1973 10.6151
R11279 GND.n1983 GND.n1974 10.6151
R11280 GND.n1984 GND.n1983 10.6151
R11281 GND.n1986 GND.n1984 10.6151
R11282 GND.n1987 GND.n1986 10.6151
R11283 GND.n1988 GND.n1987 10.6151
R11284 GND.n1988 GND.n1972 10.6151
R11285 GND.n1996 GND.n1972 10.6151
R11286 GND.n1997 GND.n1996 10.6151
R11287 GND.n1999 GND.n1997 10.6151
R11288 GND.n2000 GND.n1999 10.6151
R11289 GND.n2001 GND.n2000 10.6151
R11290 GND.n2001 GND.n1971 10.6151
R11291 GND.n2009 GND.n1971 10.6151
R11292 GND.n2010 GND.n2009 10.6151
R11293 GND.n2012 GND.n2010 10.6151
R11294 GND.n2013 GND.n2012 10.6151
R11295 GND.n2014 GND.n2013 10.6151
R11296 GND.n2017 GND.n2014 10.6151
R11297 GND.n2018 GND.n2017 10.6151
R11298 GND.n2020 GND.n2018 10.6151
R11299 GND.n2021 GND.n2020 10.6151
R11300 GND.n2022 GND.n2021 10.6151
R11301 GND.n2022 GND.n1970 10.6151
R11302 GND.n2030 GND.n1970 10.6151
R11303 GND.n2031 GND.n2030 10.6151
R11304 GND.n2033 GND.n2031 10.6151
R11305 GND.n2034 GND.n2033 10.6151
R11306 GND.n2035 GND.n2034 10.6151
R11307 GND.n2035 GND.n1969 10.6151
R11308 GND.n2043 GND.n1969 10.6151
R11309 GND.n2044 GND.n2043 10.6151
R11310 GND.n2046 GND.n2044 10.6151
R11311 GND.n2047 GND.n2046 10.6151
R11312 GND.n2048 GND.n2047 10.6151
R11313 GND.n2048 GND.n1968 10.6151
R11314 GND.n2056 GND.n1968 10.6151
R11315 GND.n2057 GND.n2056 10.6151
R11316 GND.n2059 GND.n2057 10.6151
R11317 GND.n2060 GND.n2059 10.6151
R11318 GND.n2061 GND.n2060 10.6151
R11319 GND.n2070 GND.n2061 10.6151
R11320 GND.n2071 GND.n2070 10.6151
R11321 GND.n2074 GND.n2071 10.6151
R11322 GND.n2074 GND.n2073 10.6151
R11323 GND.n2073 GND.n2072 10.6151
R11324 GND.n2072 GND.n1703 10.6151
R11325 GND.n5773 GND.n1703 10.6151
R11326 GND.n5774 GND.n5773 10.6151
R11327 GND.n5779 GND.n5774 10.6151
R11328 GND.n5779 GND.n5778 10.6151
R11329 GND.n5778 GND.n5777 10.6151
R11330 GND.n5777 GND.n5775 10.6151
R11331 GND.n5775 GND.n1666 10.6151
R11332 GND.n5841 GND.n1666 10.6151
R11333 GND.n5842 GND.n5841 10.6151
R11334 GND.n5843 GND.n5842 10.6151
R11335 GND.n5845 GND.n5843 10.6151
R11336 GND.n5845 GND.n5844 10.6151
R11337 GND.n5844 GND.n1638 10.6151
R11338 GND.n5883 GND.n1638 10.6151
R11339 GND.n5883 GND.n5882 10.6151
R11340 GND.n5882 GND.n5881 10.6151
R11341 GND.n5881 GND.n1639 10.6151
R11342 GND.n1640 GND.n1639 10.6151
R11343 GND.n1640 GND.n1596 10.6151
R11344 GND.n5922 GND.n1596 10.6151
R11345 GND.n5922 GND.n5921 10.6151
R11346 GND.n5921 GND.n5920 10.6151
R11347 GND.n5920 GND.n1597 10.6151
R11348 GND.n1610 GND.n1597 10.6151
R11349 GND.n1610 GND.n1609 10.6151
R11350 GND.n1609 GND.n1608 10.6151
R11351 GND.n1608 GND.n1607 10.6151
R11352 GND.n1607 GND.n1600 10.6151
R11353 GND.n1601 GND.n1600 10.6151
R11354 GND.n1601 GND.n1544 10.6151
R11355 GND.n6017 GND.n1544 10.6151
R11356 GND.n6018 GND.n6017 10.6151
R11357 GND.n6048 GND.n6018 10.6151
R11358 GND.n6048 GND.n6047 10.6151
R11359 GND.n6047 GND.n6046 10.6151
R11360 GND.n6046 GND.n6043 10.6151
R11361 GND.n6043 GND.n6042 10.6151
R11362 GND.n6042 GND.n6040 10.6151
R11363 GND.n6040 GND.n6039 10.6151
R11364 GND.n6039 GND.n6035 10.6151
R11365 GND.n6035 GND.n6034 10.6151
R11366 GND.n6034 GND.n6032 10.6151
R11367 GND.n6032 GND.n6031 10.6151
R11368 GND.n6031 GND.n6019 10.6151
R11369 GND.n6025 GND.n6019 10.6151
R11370 GND.n6025 GND.n6024 10.6151
R11371 GND.n6024 GND.n6023 10.6151
R11372 GND.n6023 GND.n6020 10.6151
R11373 GND.n6020 GND.n1464 10.6151
R11374 GND.n6172 GND.n1464 10.6151
R11375 GND.n6173 GND.n6172 10.6151
R11376 GND.n6174 GND.n6173 10.6151
R11377 GND.n6174 GND.n1451 10.6151
R11378 GND.n6198 GND.n1451 10.6151
R11379 GND.n6199 GND.n6198 10.6151
R11380 GND.n6233 GND.n6199 10.6151
R11381 GND.n6233 GND.n6232 10.6151
R11382 GND.n6232 GND.n6231 10.6151
R11383 GND.n6231 GND.n6228 10.6151
R11384 GND.n6228 GND.n6227 10.6151
R11385 GND.n6227 GND.n6224 10.6151
R11386 GND.n6224 GND.n6223 10.6151
R11387 GND.n6223 GND.n6200 10.6151
R11388 GND.n6210 GND.n6200 10.6151
R11389 GND.n6210 GND.n6209 10.6151
R11390 GND.n6209 GND.n6208 10.6151
R11391 GND.n6208 GND.n6204 10.6151
R11392 GND.n6204 GND.n6203 10.6151
R11393 GND.n6203 GND.n1315 10.6151
R11394 GND.n6340 GND.n1315 10.6151
R11395 GND.n6341 GND.n6340 10.6151
R11396 GND.n6346 GND.n6341 10.6151
R11397 GND.n6346 GND.n6345 10.6151
R11398 GND.n6345 GND.n6344 10.6151
R11399 GND.n6344 GND.n6342 10.6151
R11400 GND.n6342 GND.n1292 10.6151
R11401 GND.n6385 GND.n1292 10.6151
R11402 GND.n6386 GND.n6385 10.6151
R11403 GND.n6387 GND.n6386 10.6151
R11404 GND.n6387 GND.n1283 10.6151
R11405 GND.n6398 GND.n1283 10.6151
R11406 GND.n6399 GND.n6398 10.6151
R11407 GND.n6405 GND.n6399 10.6151
R11408 GND.n6405 GND.n6404 10.6151
R11409 GND.n6404 GND.n6403 10.6151
R11410 GND.n6403 GND.n6402 10.6151
R11411 GND.n6402 GND.n6400 10.6151
R11412 GND.n6400 GND.n1258 10.6151
R11413 GND.n6434 GND.n1258 10.6151
R11414 GND.n6435 GND.n6434 10.6151
R11415 GND.n6441 GND.n6435 10.6151
R11416 GND.n6441 GND.n6440 10.6151
R11417 GND.n6440 GND.n6439 10.6151
R11418 GND.n6439 GND.n6438 10.6151
R11419 GND.n6438 GND.n6436 10.6151
R11420 GND.n6436 GND.n1233 10.6151
R11421 GND.n6472 GND.n1233 10.6151
R11422 GND.n6473 GND.n6472 10.6151
R11423 GND.n6479 GND.n6473 10.6151
R11424 GND.n6479 GND.n6478 10.6151
R11425 GND.n6478 GND.n6477 10.6151
R11426 GND.n6477 GND.n6476 10.6151
R11427 GND.n6476 GND.n6474 10.6151
R11428 GND.n6474 GND.n1208 10.6151
R11429 GND.n6517 GND.n1208 10.6151
R11430 GND.n6518 GND.n6517 10.6151
R11431 GND.n6519 GND.n6518 10.6151
R11432 GND.n6519 GND.n1199 10.6151
R11433 GND.n6530 GND.n1199 10.6151
R11434 GND.n6531 GND.n6530 10.6151
R11435 GND.n6584 GND.n6531 10.6151
R11436 GND.n6584 GND.n6583 10.6151
R11437 GND.n6583 GND.n6582 10.6151
R11438 GND.n6582 GND.n6581 10.6151
R11439 GND.n6581 GND.n6579 10.6151
R11440 GND.n6579 GND.n6578 10.6151
R11441 GND.n2225 GND.n2222 10.6151
R11442 GND.n2222 GND.n2221 10.6151
R11443 GND.n2218 GND.n2217 10.6151
R11444 GND.n2217 GND.n2214 10.6151
R11445 GND.n2214 GND.n2213 10.6151
R11446 GND.n2213 GND.n2210 10.6151
R11447 GND.n2210 GND.n2209 10.6151
R11448 GND.n2209 GND.n2206 10.6151
R11449 GND.n2206 GND.n2205 10.6151
R11450 GND.n2205 GND.n2202 10.6151
R11451 GND.n2202 GND.n2201 10.6151
R11452 GND.n2201 GND.n2198 10.6151
R11453 GND.n2198 GND.n2197 10.6151
R11454 GND.n2197 GND.n2194 10.6151
R11455 GND.n2194 GND.n2193 10.6151
R11456 GND.n2193 GND.n2190 10.6151
R11457 GND.n2190 GND.n2189 10.6151
R11458 GND.n2189 GND.n2186 10.6151
R11459 GND.n2186 GND.n2185 10.6151
R11460 GND.n5673 GND.n5672 10.6151
R11461 GND.n5672 GND.n5671 10.6151
R11462 GND.n5671 GND.n5670 10.6151
R11463 GND.n5670 GND.n5668 10.6151
R11464 GND.n5668 GND.n5665 10.6151
R11465 GND.n5665 GND.n5664 10.6151
R11466 GND.n5664 GND.n5661 10.6151
R11467 GND.n5661 GND.n5660 10.6151
R11468 GND.n5660 GND.n5657 10.6151
R11469 GND.n5657 GND.n5656 10.6151
R11470 GND.n5656 GND.n5653 10.6151
R11471 GND.n5653 GND.n5652 10.6151
R11472 GND.n5652 GND.n5649 10.6151
R11473 GND.n5649 GND.n5648 10.6151
R11474 GND.n5648 GND.n5645 10.6151
R11475 GND.n5645 GND.n5644 10.6151
R11476 GND.n5644 GND.n5641 10.6151
R11477 GND.n5639 GND.n5636 10.6151
R11478 GND.n5636 GND.n5635 10.6151
R11479 GND.n6662 GND.n6661 10.6151
R11480 GND.n6661 GND.n6660 10.6151
R11481 GND.n6660 GND.n6657 10.6151
R11482 GND.n6657 GND.n6656 10.6151
R11483 GND.n6656 GND.n6653 10.6151
R11484 GND.n6653 GND.n6652 10.6151
R11485 GND.n6652 GND.n6649 10.6151
R11486 GND.n6649 GND.n6648 10.6151
R11487 GND.n6648 GND.n6645 10.6151
R11488 GND.n6645 GND.n6644 10.6151
R11489 GND.n6644 GND.n6641 10.6151
R11490 GND.n6641 GND.n6640 10.6151
R11491 GND.n6640 GND.n6637 10.6151
R11492 GND.n6637 GND.n6636 10.6151
R11493 GND.n6636 GND.n6633 10.6151
R11494 GND.n6633 GND.n6632 10.6151
R11495 GND.n6632 GND.n6629 10.6151
R11496 GND.n6627 GND.n6624 10.6151
R11497 GND.n6624 GND.n1148 10.6151
R11498 GND.n1978 GND.n1977 10.6151
R11499 GND.n1979 GND.n1978 10.6151
R11500 GND.n1979 GND.n1837 10.6151
R11501 GND.n2172 GND.n1837 10.6151
R11502 GND.n2172 GND.n2171 10.6151
R11503 GND.n2171 GND.n2170 10.6151
R11504 GND.n2170 GND.n1838 10.6151
R11505 GND.n1991 GND.n1838 10.6151
R11506 GND.n1991 GND.n1854 10.6151
R11507 GND.n2158 GND.n1854 10.6151
R11508 GND.n2158 GND.n2157 10.6151
R11509 GND.n2157 GND.n2156 10.6151
R11510 GND.n2156 GND.n1855 10.6151
R11511 GND.n2004 GND.n1855 10.6151
R11512 GND.n2004 GND.n1873 10.6151
R11513 GND.n2144 GND.n1873 10.6151
R11514 GND.n2144 GND.n2143 10.6151
R11515 GND.n2143 GND.n2142 10.6151
R11516 GND.n2142 GND.n1874 10.6151
R11517 GND.n1892 GND.n1874 10.6151
R11518 GND.n2130 GND.n1892 10.6151
R11519 GND.n2130 GND.n2129 10.6151
R11520 GND.n2129 GND.n2128 10.6151
R11521 GND.n2128 GND.n1893 10.6151
R11522 GND.n2025 GND.n1893 10.6151
R11523 GND.n2025 GND.n1910 10.6151
R11524 GND.n2116 GND.n1910 10.6151
R11525 GND.n2116 GND.n2115 10.6151
R11526 GND.n2115 GND.n2114 10.6151
R11527 GND.n2114 GND.n1911 10.6151
R11528 GND.n2038 GND.n1911 10.6151
R11529 GND.n2038 GND.n1928 10.6151
R11530 GND.n2102 GND.n1928 10.6151
R11531 GND.n2102 GND.n2101 10.6151
R11532 GND.n2101 GND.n2100 10.6151
R11533 GND.n2100 GND.n1929 10.6151
R11534 GND.n2051 GND.n1929 10.6151
R11535 GND.n2051 GND.n1946 10.6151
R11536 GND.n2088 GND.n1946 10.6151
R11537 GND.n2088 GND.n2087 10.6151
R11538 GND.n2087 GND.n2086 10.6151
R11539 GND.n2086 GND.n1947 10.6151
R11540 GND.n2066 GND.n1947 10.6151
R11541 GND.n2066 GND.n2065 10.6151
R11542 GND.n2065 GND.n1708 10.6151
R11543 GND.n5766 GND.n1708 10.6151
R11544 GND.n5767 GND.n5766 10.6151
R11545 GND.n5768 GND.n5767 10.6151
R11546 GND.n5768 GND.n1689 10.6151
R11547 GND.n5816 GND.n1689 10.6151
R11548 GND.n5816 GND.n5815 10.6151
R11549 GND.n5815 GND.n5814 10.6151
R11550 GND.n5814 GND.n1690 10.6151
R11551 GND.n1693 GND.n1690 10.6151
R11552 GND.n1693 GND.n1692 10.6151
R11553 GND.n1692 GND.n1661 10.6151
R11554 GND.n5851 GND.n1661 10.6151
R11555 GND.n5851 GND.n5850 10.6151
R11556 GND.n5850 GND.n5849 10.6151
R11557 GND.n5849 GND.n1633 10.6151
R11558 GND.n5889 GND.n1633 10.6151
R11559 GND.n5890 GND.n5889 10.6151
R11560 GND.n5894 GND.n5890 10.6151
R11561 GND.n5894 GND.n5893 10.6151
R11562 GND.n5893 GND.n5892 10.6151
R11563 GND.n5892 GND.n1591 10.6151
R11564 GND.n5928 GND.n1591 10.6151
R11565 GND.n5929 GND.n5928 10.6151
R11566 GND.n5935 GND.n5929 10.6151
R11567 GND.n5935 GND.n5934 10.6151
R11568 GND.n5934 GND.n5933 10.6151
R11569 GND.n5933 GND.n5930 10.6151
R11570 GND.n5930 GND.n1567 10.6151
R11571 GND.n5983 GND.n1567 10.6151
R11572 GND.n5983 GND.n5982 10.6151
R11573 GND.n5982 GND.n5981 10.6151
R11574 GND.n5981 GND.n1568 10.6151
R11575 GND.n1569 GND.n1568 10.6151
R11576 GND.n1569 GND.n1539 10.6151
R11577 GND.n6054 GND.n1539 10.6151
R11578 GND.n6055 GND.n6054 10.6151
R11579 GND.n6056 GND.n6055 10.6151
R11580 GND.n6056 GND.n1522 10.6151
R11581 GND.n6071 GND.n1522 10.6151
R11582 GND.n6072 GND.n6071 10.6151
R11583 GND.n6073 GND.n6072 10.6151
R11584 GND.n6073 GND.n1508 10.6151
R11585 GND.n6089 GND.n1508 10.6151
R11586 GND.n6090 GND.n6089 10.6151
R11587 GND.n6094 GND.n6090 10.6151
R11588 GND.n6094 GND.n6093 10.6151
R11589 GND.n6093 GND.n6092 10.6151
R11590 GND.n6092 GND.n1489 10.6151
R11591 GND.n6138 GND.n1489 10.6151
R11592 GND.n6138 GND.n6137 10.6151
R11593 GND.n6137 GND.n6136 10.6151
R11594 GND.n6136 GND.n1490 10.6151
R11595 GND.n1490 GND.n1463 10.6151
R11596 GND.n6182 GND.n1463 10.6151
R11597 GND.n6182 GND.n6181 10.6151
R11598 GND.n6181 GND.n6180 10.6151
R11599 GND.n6180 GND.n1447 10.6151
R11600 GND.n6239 GND.n1447 10.6151
R11601 GND.n6240 GND.n6239 10.6151
R11602 GND.n6241 GND.n6240 10.6151
R11603 GND.n6241 GND.n1433 10.6151
R11604 GND.n6258 GND.n1433 10.6151
R11605 GND.n6258 GND.n6257 10.6151
R11606 GND.n6257 GND.n6256 10.6151
R11607 GND.n6256 GND.n1434 10.6151
R11608 GND.n6218 GND.n1434 10.6151
R11609 GND.n6218 GND.n6217 10.6151
R11610 GND.n6217 GND.n6216 10.6151
R11611 GND.n6216 GND.n1319 10.6151
R11612 GND.n6333 GND.n1319 10.6151
R11613 GND.n6334 GND.n6333 10.6151
R11614 GND.n6335 GND.n6334 10.6151
R11615 GND.n6335 GND.n1311 10.6151
R11616 GND.n6352 GND.n1311 10.6151
R11617 GND.n6353 GND.n6352 10.6151
R11618 GND.n6354 GND.n6353 10.6151
R11619 GND.n6354 GND.n1298 10.6151
R11620 GND.n6379 GND.n1298 10.6151
R11621 GND.n6380 GND.n6379 10.6151
R11622 GND.n6381 GND.n6380 10.6151
R11623 GND.n6381 GND.n1288 10.6151
R11624 GND.n6392 GND.n1288 10.6151
R11625 GND.n6393 GND.n6392 10.6151
R11626 GND.n6394 GND.n6393 10.6151
R11627 GND.n6394 GND.n1278 10.6151
R11628 GND.n6410 GND.n1278 10.6151
R11629 GND.n6411 GND.n6410 10.6151
R11630 GND.n6412 GND.n6411 10.6151
R11631 GND.n6412 GND.n1264 10.6151
R11632 GND.n6428 GND.n1264 10.6151
R11633 GND.n6429 GND.n6428 10.6151
R11634 GND.n6430 GND.n6429 10.6151
R11635 GND.n6430 GND.n1253 10.6151
R11636 GND.n6445 GND.n1253 10.6151
R11637 GND.n6446 GND.n6445 10.6151
R11638 GND.n6447 GND.n6446 10.6151
R11639 GND.n6447 GND.n1238 10.6151
R11640 GND.n6466 GND.n1238 10.6151
R11641 GND.n6467 GND.n6466 10.6151
R11642 GND.n6468 GND.n6467 10.6151
R11643 GND.n6468 GND.n1228 10.6151
R11644 GND.n6484 GND.n1228 10.6151
R11645 GND.n6485 GND.n6484 10.6151
R11646 GND.n6486 GND.n6485 10.6151
R11647 GND.n6486 GND.n1214 10.6151
R11648 GND.n6511 GND.n1214 10.6151
R11649 GND.n6512 GND.n6511 10.6151
R11650 GND.n6513 GND.n6512 10.6151
R11651 GND.n6513 GND.n1204 10.6151
R11652 GND.n6524 GND.n1204 10.6151
R11653 GND.n6525 GND.n6524 10.6151
R11654 GND.n6526 GND.n6525 10.6151
R11655 GND.n6526 GND.n1194 10.6151
R11656 GND.n6589 GND.n1194 10.6151
R11657 GND.n6590 GND.n6589 10.6151
R11658 GND.n6591 GND.n6590 10.6151
R11659 GND.n6591 GND.n1180 10.6151
R11660 GND.n6619 GND.n1180 10.6151
R11661 GND.n6620 GND.n6619 10.6151
R11662 GND.n5630 GND.n5629 10.4732
R11663 GND.n6709 GND.n6708 10.4732
R11664 GND.t38 GND.n5808 10.3706
R11665 GND.n6253 GND.t79 10.3706
R11666 GND.n80 GND.n79 10.2326
R11667 GND.n101 GND.n100 10.2326
R11668 GND.n42 GND.n41 10.2326
R11669 GND.n63 GND.n62 10.2326
R11670 GND.n5 GND.n4 10.2326
R11671 GND.n26 GND.n25 10.2326
R11672 GND.n215 GND.n214 10.2326
R11673 GND.n194 GND.n193 10.2326
R11674 GND.n177 GND.n176 10.2326
R11675 GND.n156 GND.n155 10.2326
R11676 GND.n140 GND.n139 10.2326
R11677 GND.n119 GND.n118 10.2326
R11678 GND.n2182 GND.n2181 9.98653
R11679 GND.n2006 GND.n2003 9.98653
R11680 GND.n2027 GND.n2024 9.98653
R11681 GND.n2112 GND.t7 9.98653
R11682 GND.n2091 GND.n2090 9.98653
R11683 GND.n2063 GND.t84 9.98653
R11684 GND.n5818 GND.n1686 9.98653
R11685 GND.n5879 GND.n1630 9.98653
R11686 GND.n1605 GND.n1604 9.98653
R11687 GND.n6086 GND.n1502 9.98653
R11688 GND.n6177 GND.n6176 9.98653
R11689 GND.n6206 GND.n6205 9.98653
R11690 GND.n6357 GND.t6 9.98653
R11691 GND.n6383 GND.n1296 9.98653
R11692 GND.n6426 GND.t4 9.98653
R11693 GND.n6443 GND.n1255 9.98653
R11694 GND.n1226 GND.n1216 9.98653
R11695 GND.n7449 GND.n7448 9.89141
R11696 GND.n3166 GND.n3068 9.89141
R11697 GND.n89 GND.n75 9.69747
R11698 GND.n110 GND.n96 9.69747
R11699 GND.n51 GND.n37 9.69747
R11700 GND.n72 GND.n58 9.69747
R11701 GND.n14 GND.n0 9.69747
R11702 GND.n35 GND.n21 9.69747
R11703 GND.n224 GND.n210 9.69747
R11704 GND.n203 GND.n189 9.69747
R11705 GND.n186 GND.n172 9.69747
R11706 GND.n165 GND.n151 9.69747
R11707 GND.n149 GND.n135 9.69747
R11708 GND.n128 GND.n114 9.69747
R11709 GND.n113 GND.n112 9.54346
R11710 GND.n7646 GND.n226 9.54346
R11711 GND.t105 GND.n2877 9.4588
R11712 GND.n89 GND.n88 9.45567
R11713 GND.n110 GND.n109 9.45567
R11714 GND.n51 GND.n50 9.45567
R11715 GND.n72 GND.n71 9.45567
R11716 GND.n14 GND.n13 9.45567
R11717 GND.n35 GND.n34 9.45567
R11718 GND.n224 GND.n223 9.45567
R11719 GND.n203 GND.n202 9.45567
R11720 GND.n186 GND.n185 9.45567
R11721 GND.n165 GND.n164 9.45567
R11722 GND.n149 GND.n148 9.45567
R11723 GND.n128 GND.n127 9.45567
R11724 GND.n77 GND.n76 9.3005
R11725 GND.n88 GND.n87 9.3005
R11726 GND.n82 GND.n81 9.3005
R11727 GND.n98 GND.n97 9.3005
R11728 GND.n109 GND.n108 9.3005
R11729 GND.n103 GND.n102 9.3005
R11730 GND.n39 GND.n38 9.3005
R11731 GND.n50 GND.n49 9.3005
R11732 GND.n44 GND.n43 9.3005
R11733 GND.n60 GND.n59 9.3005
R11734 GND.n71 GND.n70 9.3005
R11735 GND.n65 GND.n64 9.3005
R11736 GND.n2 GND.n1 9.3005
R11737 GND.n13 GND.n12 9.3005
R11738 GND.n7 GND.n6 9.3005
R11739 GND.n23 GND.n22 9.3005
R11740 GND.n34 GND.n33 9.3005
R11741 GND.n28 GND.n27 9.3005
R11742 GND.n212 GND.n211 9.3005
R11743 GND.n223 GND.n222 9.3005
R11744 GND.n217 GND.n216 9.3005
R11745 GND.n191 GND.n190 9.3005
R11746 GND.n202 GND.n201 9.3005
R11747 GND.n196 GND.n195 9.3005
R11748 GND.n174 GND.n173 9.3005
R11749 GND.n185 GND.n184 9.3005
R11750 GND.n179 GND.n178 9.3005
R11751 GND.n153 GND.n152 9.3005
R11752 GND.n164 GND.n163 9.3005
R11753 GND.n158 GND.n157 9.3005
R11754 GND.n137 GND.n136 9.3005
R11755 GND.n148 GND.n147 9.3005
R11756 GND.n142 GND.n141 9.3005
R11757 GND.n116 GND.n115 9.3005
R11758 GND.n127 GND.n126 9.3005
R11759 GND.n121 GND.n120 9.3005
R11760 GND.n1378 GND.n1360 9.3005
R11761 GND.n1375 GND.n1371 9.3005
R11762 GND.n1374 GND.n1373 9.3005
R11763 GND.n906 GND.n905 9.3005
R11764 GND.n6765 GND.n6764 9.3005
R11765 GND.n6766 GND.n904 9.3005
R11766 GND.n6850 GND.n6767 9.3005
R11767 GND.n6849 GND.n6768 9.3005
R11768 GND.n6848 GND.n6769 9.3005
R11769 GND.n6846 GND.n6770 9.3005
R11770 GND.n6845 GND.n6771 9.3005
R11771 GND.n6843 GND.n6772 9.3005
R11772 GND.n6842 GND.n6773 9.3005
R11773 GND.n6840 GND.n6774 9.3005
R11774 GND.n6839 GND.n6775 9.3005
R11775 GND.n6837 GND.n6776 9.3005
R11776 GND.n6836 GND.n6777 9.3005
R11777 GND.n6834 GND.n6778 9.3005
R11778 GND.n6833 GND.n6779 9.3005
R11779 GND.n6831 GND.n6780 9.3005
R11780 GND.n6830 GND.n6781 9.3005
R11781 GND.n6828 GND.n6782 9.3005
R11782 GND.n6827 GND.n6783 9.3005
R11783 GND.n6825 GND.n6784 9.3005
R11784 GND.n6824 GND.n6785 9.3005
R11785 GND.n6822 GND.n6786 9.3005
R11786 GND.n6821 GND.n6787 9.3005
R11787 GND.n6819 GND.n6788 9.3005
R11788 GND.n6818 GND.n6789 9.3005
R11789 GND.n6816 GND.n6790 9.3005
R11790 GND.n6815 GND.n6791 9.3005
R11791 GND.n6813 GND.n6792 9.3005
R11792 GND.n6812 GND.n6793 9.3005
R11793 GND.n6810 GND.n6794 9.3005
R11794 GND.n6809 GND.n6795 9.3005
R11795 GND.n6807 GND.n6796 9.3005
R11796 GND.n6806 GND.n6797 9.3005
R11797 GND.n6804 GND.n6798 9.3005
R11798 GND.n6803 GND.n6799 9.3005
R11799 GND.n6801 GND.n6800 9.3005
R11800 GND.n718 GND.n717 9.3005
R11801 GND.n7040 GND.n7039 9.3005
R11802 GND.n7041 GND.n716 9.3005
R11803 GND.n7058 GND.n7042 9.3005
R11804 GND.n7057 GND.n7043 9.3005
R11805 GND.n7056 GND.n7044 9.3005
R11806 GND.n7054 GND.n7045 9.3005
R11807 GND.n7053 GND.n7046 9.3005
R11808 GND.n7051 GND.n7047 9.3005
R11809 GND.n7050 GND.n7049 9.3005
R11810 GND.n7048 GND.n671 9.3005
R11811 GND.n7110 GND.n670 9.3005
R11812 GND.n7112 GND.n7111 9.3005
R11813 GND.n7113 GND.n669 9.3005
R11814 GND.n7127 GND.n7114 9.3005
R11815 GND.n7126 GND.n7115 9.3005
R11816 GND.n7125 GND.n7116 9.3005
R11817 GND.n7123 GND.n7117 9.3005
R11818 GND.n7122 GND.n7118 9.3005
R11819 GND.n7120 GND.n7119 9.3005
R11820 GND.n229 GND.n227 9.3005
R11821 GND.n1377 GND.n1376 9.3005
R11822 GND.n7644 GND.n7643 9.3005
R11823 GND.n230 GND.n228 9.3005
R11824 GND.n617 GND.n616 9.3005
R11825 GND.n615 GND.n614 9.3005
R11826 GND.n7212 GND.n7211 9.3005
R11827 GND.n7213 GND.n613 9.3005
R11828 GND.n7216 GND.n7214 9.3005
R11829 GND.n7217 GND.n612 9.3005
R11830 GND.n7220 GND.n7219 9.3005
R11831 GND.n7221 GND.n611 9.3005
R11832 GND.n7224 GND.n7222 9.3005
R11833 GND.n7225 GND.n610 9.3005
R11834 GND.n7228 GND.n7227 9.3005
R11835 GND.n7229 GND.n609 9.3005
R11836 GND.n7232 GND.n7230 9.3005
R11837 GND.n7233 GND.n608 9.3005
R11838 GND.n7237 GND.n7236 9.3005
R11839 GND.n7238 GND.n607 9.3005
R11840 GND.n7241 GND.n7239 9.3005
R11841 GND.n7242 GND.n606 9.3005
R11842 GND.n7245 GND.n7244 9.3005
R11843 GND.n7246 GND.n605 9.3005
R11844 GND.n7249 GND.n7247 9.3005
R11845 GND.n7250 GND.n604 9.3005
R11846 GND.n7253 GND.n7252 9.3005
R11847 GND.n7254 GND.n603 9.3005
R11848 GND.n7257 GND.n7255 9.3005
R11849 GND.n7258 GND.n602 9.3005
R11850 GND.n7261 GND.n7260 9.3005
R11851 GND.n7262 GND.n601 9.3005
R11852 GND.n7265 GND.n7263 9.3005
R11853 GND.n7266 GND.n600 9.3005
R11854 GND.n7269 GND.n7268 9.3005
R11855 GND.n7270 GND.n599 9.3005
R11856 GND.n7273 GND.n7271 9.3005
R11857 GND.n7274 GND.n598 9.3005
R11858 GND.n7277 GND.n7276 9.3005
R11859 GND.n7278 GND.n597 9.3005
R11860 GND.n7281 GND.n7279 9.3005
R11861 GND.n7282 GND.n596 9.3005
R11862 GND.n7285 GND.n7284 9.3005
R11863 GND.n7286 GND.n595 9.3005
R11864 GND.n7289 GND.n7287 9.3005
R11865 GND.n7290 GND.n594 9.3005
R11866 GND.n7293 GND.n7292 9.3005
R11867 GND.n7294 GND.n593 9.3005
R11868 GND.n7297 GND.n7295 9.3005
R11869 GND.n7298 GND.n592 9.3005
R11870 GND.n7301 GND.n7300 9.3005
R11871 GND.n7302 GND.n591 9.3005
R11872 GND.n7305 GND.n7303 9.3005
R11873 GND.n7306 GND.n590 9.3005
R11874 GND.n7309 GND.n7308 9.3005
R11875 GND.n7310 GND.n589 9.3005
R11876 GND.n7313 GND.n7311 9.3005
R11877 GND.n7314 GND.n588 9.3005
R11878 GND.n7317 GND.n7316 9.3005
R11879 GND.n7318 GND.n587 9.3005
R11880 GND.n7321 GND.n7319 9.3005
R11881 GND.n7322 GND.n586 9.3005
R11882 GND.n7324 GND.n7323 9.3005
R11883 GND.n568 GND.n567 9.3005
R11884 GND.n7340 GND.n570 9.3005
R11885 GND.n7339 GND.n571 9.3005
R11886 GND.n7338 GND.n572 9.3005
R11887 GND.n576 GND.n573 9.3005
R11888 GND.n7333 GND.n577 9.3005
R11889 GND.n7332 GND.n578 9.3005
R11890 GND.n7331 GND.n579 9.3005
R11891 GND.n585 GND.n582 9.3005
R11892 GND.n7326 GND.n7325 9.3005
R11893 GND.n7346 GND.n7345 9.3005
R11894 GND.n527 GND.n526 9.3005
R11895 GND.n531 GND.n529 9.3005
R11896 GND.n7457 GND.n532 9.3005
R11897 GND.n7456 GND.n533 9.3005
R11898 GND.n7455 GND.n534 9.3005
R11899 GND.n538 GND.n535 9.3005
R11900 GND.n7450 GND.n539 9.3005
R11901 GND.n7449 GND.n540 9.3005
R11902 GND.n7448 GND.n7447 9.3005
R11903 GND.n7446 GND.n541 9.3005
R11904 GND.n7445 GND.n7444 9.3005
R11905 GND.n547 GND.n546 9.3005
R11906 GND.n7439 GND.n551 9.3005
R11907 GND.n7438 GND.n552 9.3005
R11908 GND.n7437 GND.n553 9.3005
R11909 GND.n557 GND.n554 9.3005
R11910 GND.n7432 GND.n558 9.3005
R11911 GND.n7431 GND.n559 9.3005
R11912 GND.n7430 GND.n560 9.3005
R11913 GND.n566 GND.n563 9.3005
R11914 GND.n7425 GND.n7424 9.3005
R11915 GND.n7465 GND.n7464 9.3005
R11916 GND.n6739 GND.n6738 9.3005
R11917 GND.n6740 GND.n925 9.3005
R11918 GND.n6742 GND.n926 9.3005
R11919 GND.n6744 GND.n6743 9.3005
R11920 GND.n6745 GND.n898 9.3005
R11921 GND.n6854 GND.n899 9.3005
R11922 GND.n6855 GND.n897 9.3005
R11923 GND.n6857 GND.n6856 9.3005
R11924 GND.n6858 GND.n879 9.3005
R11925 GND.n6874 GND.n880 9.3005
R11926 GND.n6875 GND.n878 9.3005
R11927 GND.n6877 GND.n6876 9.3005
R11928 GND.n6878 GND.n859 9.3005
R11929 GND.n6894 GND.n860 9.3005
R11930 GND.n6895 GND.n858 9.3005
R11931 GND.n6897 GND.n6896 9.3005
R11932 GND.n6898 GND.n839 9.3005
R11933 GND.n6914 GND.n840 9.3005
R11934 GND.n6915 GND.n838 9.3005
R11935 GND.n6917 GND.n6916 9.3005
R11936 GND.n6918 GND.n819 9.3005
R11937 GND.n6934 GND.n820 9.3005
R11938 GND.n6935 GND.n818 9.3005
R11939 GND.n6937 GND.n6936 9.3005
R11940 GND.n6938 GND.n799 9.3005
R11941 GND.n6954 GND.n800 9.3005
R11942 GND.n6955 GND.n798 9.3005
R11943 GND.n6957 GND.n6956 9.3005
R11944 GND.n6958 GND.n779 9.3005
R11945 GND.n6974 GND.n780 9.3005
R11946 GND.n6975 GND.n778 9.3005
R11947 GND.n6977 GND.n6976 9.3005
R11948 GND.n6978 GND.n759 9.3005
R11949 GND.n6994 GND.n760 9.3005
R11950 GND.n6995 GND.n758 9.3005
R11951 GND.n6997 GND.n6996 9.3005
R11952 GND.n6998 GND.n739 9.3005
R11953 GND.n7014 GND.n740 9.3005
R11954 GND.n7015 GND.n737 9.3005
R11955 GND.n7017 GND.n738 9.3005
R11956 GND.n7019 GND.n7018 9.3005
R11957 GND.n7020 GND.n710 9.3005
R11958 GND.n7062 GND.n711 9.3005
R11959 GND.n7063 GND.n709 9.3005
R11960 GND.n7065 GND.n7064 9.3005
R11961 GND.n7066 GND.n691 9.3005
R11962 GND.n7082 GND.n692 9.3005
R11963 GND.n7083 GND.n689 9.3005
R11964 GND.n7085 GND.n690 9.3005
R11965 GND.n7094 GND.n7086 9.3005
R11966 GND.n7093 GND.n7092 9.3005
R11967 GND.n7090 GND.n662 9.3005
R11968 GND.n7089 GND.n663 9.3005
R11969 GND.n7087 GND.n664 9.3005
R11970 GND.n665 GND.n642 9.3005
R11971 GND.n7148 GND.n643 9.3005
R11972 GND.n7149 GND.n641 9.3005
R11973 GND.n7156 GND.n7151 9.3005
R11974 GND.n7155 GND.n7154 9.3005
R11975 GND.n7153 GND.n628 9.3005
R11976 GND.n626 GND.n625 9.3005
R11977 GND.n7176 GND.n7175 9.3005
R11978 GND.n7179 GND.n624 9.3005
R11979 GND.n7202 GND.n7180 9.3005
R11980 GND.n7201 GND.n7200 9.3005
R11981 GND.n7198 GND.n259 9.3005
R11982 GND.n7197 GND.n260 9.3005
R11983 GND.n7195 GND.n261 9.3005
R11984 GND.n7194 GND.n7181 9.3005
R11985 GND.n7192 GND.n280 9.3005
R11986 GND.n7191 GND.n281 9.3005
R11987 GND.n7189 GND.n282 9.3005
R11988 GND.n7188 GND.n7182 9.3005
R11989 GND.n7186 GND.n301 9.3005
R11990 GND.n7185 GND.n302 9.3005
R11991 GND.n7183 GND.n303 9.3005
R11992 GND.n323 GND.n322 9.3005
R11993 GND.n7594 GND.n324 9.3005
R11994 GND.n7593 GND.n325 9.3005
R11995 GND.n7592 GND.n326 9.3005
R11996 GND.n7351 GND.n327 9.3005
R11997 GND.n7582 GND.n343 9.3005
R11998 GND.n7581 GND.n344 9.3005
R11999 GND.n7580 GND.n345 9.3005
R12000 GND.n7358 GND.n346 9.3005
R12001 GND.n7570 GND.n362 9.3005
R12002 GND.n7569 GND.n363 9.3005
R12003 GND.n7568 GND.n364 9.3005
R12004 GND.n7365 GND.n365 9.3005
R12005 GND.n7558 GND.n381 9.3005
R12006 GND.n7557 GND.n382 9.3005
R12007 GND.n7556 GND.n383 9.3005
R12008 GND.n7372 GND.n384 9.3005
R12009 GND.n7546 GND.n400 9.3005
R12010 GND.n7545 GND.n401 9.3005
R12011 GND.n7544 GND.n402 9.3005
R12012 GND.n7379 GND.n403 9.3005
R12013 GND.n7534 GND.n419 9.3005
R12014 GND.n7533 GND.n420 9.3005
R12015 GND.n7532 GND.n421 9.3005
R12016 GND.n7386 GND.n422 9.3005
R12017 GND.n7522 GND.n438 9.3005
R12018 GND.n7521 GND.n439 9.3005
R12019 GND.n7520 GND.n440 9.3005
R12020 GND.n7393 GND.n441 9.3005
R12021 GND.n7510 GND.n458 9.3005
R12022 GND.n7509 GND.n459 9.3005
R12023 GND.n7508 GND.n460 9.3005
R12024 GND.n7400 GND.n461 9.3005
R12025 GND.n7498 GND.n477 9.3005
R12026 GND.n7497 GND.n478 9.3005
R12027 GND.n7496 GND.n479 9.3005
R12028 GND.n7407 GND.n480 9.3005
R12029 GND.n7486 GND.n495 9.3005
R12030 GND.n7485 GND.n496 9.3005
R12031 GND.n7484 GND.n497 9.3005
R12032 GND.n7414 GND.n498 9.3005
R12033 GND.n7474 GND.n515 9.3005
R12034 GND.n7473 GND.n516 9.3005
R12035 GND.n7472 GND.n517 9.3005
R12036 GND.n7422 GND.n518 9.3005
R12037 GND.n6737 GND.n927 9.3005
R12038 GND.n6738 GND.n924 9.3005
R12039 GND.n6750 GND.n925 9.3005
R12040 GND.n6749 GND.n926 9.3005
R12041 GND.n6748 GND.n6744 9.3005
R12042 GND.n6747 GND.n6745 9.3005
R12043 GND.n899 GND.n896 9.3005
R12044 GND.n6861 GND.n897 9.3005
R12045 GND.n6860 GND.n6857 9.3005
R12046 GND.n6859 GND.n6858 9.3005
R12047 GND.n880 GND.n877 9.3005
R12048 GND.n6881 GND.n878 9.3005
R12049 GND.n6880 GND.n6877 9.3005
R12050 GND.n6879 GND.n6878 9.3005
R12051 GND.n860 GND.n857 9.3005
R12052 GND.n6901 GND.n858 9.3005
R12053 GND.n6900 GND.n6897 9.3005
R12054 GND.n6899 GND.n6898 9.3005
R12055 GND.n840 GND.n837 9.3005
R12056 GND.n6921 GND.n838 9.3005
R12057 GND.n6920 GND.n6917 9.3005
R12058 GND.n6919 GND.n6918 9.3005
R12059 GND.n820 GND.n817 9.3005
R12060 GND.n6941 GND.n818 9.3005
R12061 GND.n6940 GND.n6937 9.3005
R12062 GND.n6939 GND.n6938 9.3005
R12063 GND.n800 GND.n797 9.3005
R12064 GND.n6961 GND.n798 9.3005
R12065 GND.n6960 GND.n6957 9.3005
R12066 GND.n6959 GND.n6958 9.3005
R12067 GND.n780 GND.n777 9.3005
R12068 GND.n6981 GND.n778 9.3005
R12069 GND.n6980 GND.n6977 9.3005
R12070 GND.n6979 GND.n6978 9.3005
R12071 GND.n760 GND.n757 9.3005
R12072 GND.n7001 GND.n758 9.3005
R12073 GND.n7000 GND.n6997 9.3005
R12074 GND.n6999 GND.n6998 9.3005
R12075 GND.n740 GND.n736 9.3005
R12076 GND.n7025 GND.n737 9.3005
R12077 GND.n7024 GND.n738 9.3005
R12078 GND.n7023 GND.n7019 9.3005
R12079 GND.n7022 GND.n7020 9.3005
R12080 GND.n711 GND.n708 9.3005
R12081 GND.n7069 GND.n709 9.3005
R12082 GND.n7068 GND.n7065 9.3005
R12083 GND.n7067 GND.n7066 9.3005
R12084 GND.n692 GND.n688 9.3005
R12085 GND.n7097 GND.n689 9.3005
R12086 GND.n7096 GND.n690 9.3005
R12087 GND.n7095 GND.n7094 9.3005
R12088 GND.n7093 GND.n661 9.3005
R12089 GND.n7133 GND.n662 9.3005
R12090 GND.n7132 GND.n663 9.3005
R12091 GND.n7131 GND.n664 9.3005
R12092 GND.n666 GND.n665 9.3005
R12093 GND.n643 GND.n640 9.3005
R12094 GND.n7158 GND.n641 9.3005
R12095 GND.n7157 GND.n7156 9.3005
R12096 GND.n7155 GND.n627 9.3005
R12097 GND.n7171 GND.n628 9.3005
R12098 GND.n7172 GND.n626 9.3005
R12099 GND.n7175 GND.n7174 9.3005
R12100 GND.n624 GND.n623 9.3005
R12101 GND.n7203 GND.n7202 9.3005
R12102 GND.n7201 GND.n258 9.3005
R12103 GND.n7630 GND.n259 9.3005
R12104 GND.n7629 GND.n260 9.3005
R12105 GND.n7628 GND.n261 9.3005
R12106 GND.n7181 GND.n262 9.3005
R12107 GND.n7618 GND.n280 9.3005
R12108 GND.n7617 GND.n281 9.3005
R12109 GND.n7616 GND.n282 9.3005
R12110 GND.n7182 GND.n283 9.3005
R12111 GND.n7606 GND.n301 9.3005
R12112 GND.n7605 GND.n302 9.3005
R12113 GND.n7604 GND.n303 9.3005
R12114 GND.n323 GND.n304 9.3005
R12115 GND.n7347 GND.n324 9.3005
R12116 GND.n7349 GND.n325 9.3005
R12117 GND.n7350 GND.n326 9.3005
R12118 GND.n7353 GND.n7351 9.3005
R12119 GND.n7354 GND.n343 9.3005
R12120 GND.n7356 GND.n344 9.3005
R12121 GND.n7357 GND.n345 9.3005
R12122 GND.n7360 GND.n7358 9.3005
R12123 GND.n7361 GND.n362 9.3005
R12124 GND.n7363 GND.n363 9.3005
R12125 GND.n7364 GND.n364 9.3005
R12126 GND.n7367 GND.n7365 9.3005
R12127 GND.n7368 GND.n381 9.3005
R12128 GND.n7370 GND.n382 9.3005
R12129 GND.n7371 GND.n383 9.3005
R12130 GND.n7374 GND.n7372 9.3005
R12131 GND.n7375 GND.n400 9.3005
R12132 GND.n7377 GND.n401 9.3005
R12133 GND.n7378 GND.n402 9.3005
R12134 GND.n7381 GND.n7379 9.3005
R12135 GND.n7382 GND.n419 9.3005
R12136 GND.n7384 GND.n420 9.3005
R12137 GND.n7385 GND.n421 9.3005
R12138 GND.n7388 GND.n7386 9.3005
R12139 GND.n7389 GND.n438 9.3005
R12140 GND.n7391 GND.n439 9.3005
R12141 GND.n7392 GND.n440 9.3005
R12142 GND.n7395 GND.n7393 9.3005
R12143 GND.n7396 GND.n458 9.3005
R12144 GND.n7398 GND.n459 9.3005
R12145 GND.n7399 GND.n460 9.3005
R12146 GND.n7402 GND.n7400 9.3005
R12147 GND.n7403 GND.n477 9.3005
R12148 GND.n7405 GND.n478 9.3005
R12149 GND.n7406 GND.n479 9.3005
R12150 GND.n7409 GND.n7407 9.3005
R12151 GND.n7410 GND.n495 9.3005
R12152 GND.n7412 GND.n496 9.3005
R12153 GND.n7413 GND.n497 9.3005
R12154 GND.n7416 GND.n7414 9.3005
R12155 GND.n7417 GND.n515 9.3005
R12156 GND.n7419 GND.n516 9.3005
R12157 GND.n7420 GND.n517 9.3005
R12158 GND.n7422 GND.n7421 9.3005
R12159 GND.n6737 GND.n6736 9.3005
R12160 GND.n6689 GND.n6688 9.3005
R12161 GND.n6692 GND.n6680 9.3005
R12162 GND.n6693 GND.n6679 9.3005
R12163 GND.n6696 GND.n6678 9.3005
R12164 GND.n6697 GND.n6677 9.3005
R12165 GND.n6700 GND.n6676 9.3005
R12166 GND.n6701 GND.n6675 9.3005
R12167 GND.n6704 GND.n6674 9.3005
R12168 GND.n6705 GND.n6673 9.3005
R12169 GND.n6708 GND.n6672 9.3005
R12170 GND.n6710 GND.n1146 9.3005
R12171 GND.n6713 GND.n1145 9.3005
R12172 GND.n6714 GND.n1144 9.3005
R12173 GND.n6717 GND.n1143 9.3005
R12174 GND.n6719 GND.n1142 9.3005
R12175 GND.n6720 GND.n1141 9.3005
R12176 GND.n6721 GND.n1140 9.3005
R12177 GND.n6722 GND.n1139 9.3005
R12178 GND.n6687 GND.n6684 9.3005
R12179 GND.n6686 GND.n6685 9.3005
R12180 GND.n1136 GND.n958 9.3005
R12181 GND.n1134 GND.n959 9.3005
R12182 GND.n1133 GND.n960 9.3005
R12183 GND.n1131 GND.n961 9.3005
R12184 GND.n1130 GND.n962 9.3005
R12185 GND.n1128 GND.n963 9.3005
R12186 GND.n1127 GND.n964 9.3005
R12187 GND.n1126 GND.n965 9.3005
R12188 GND.n1124 GND.n966 9.3005
R12189 GND.n1123 GND.n967 9.3005
R12190 GND.n1121 GND.n968 9.3005
R12191 GND.n1120 GND.n969 9.3005
R12192 GND.n1118 GND.n970 9.3005
R12193 GND.n1117 GND.n971 9.3005
R12194 GND.n1115 GND.n972 9.3005
R12195 GND.n1114 GND.n973 9.3005
R12196 GND.n1112 GND.n974 9.3005
R12197 GND.n1111 GND.n975 9.3005
R12198 GND.n1109 GND.n976 9.3005
R12199 GND.n1108 GND.n977 9.3005
R12200 GND.n1106 GND.n978 9.3005
R12201 GND.n1105 GND.n979 9.3005
R12202 GND.n1103 GND.n980 9.3005
R12203 GND.n1102 GND.n981 9.3005
R12204 GND.n1100 GND.n982 9.3005
R12205 GND.n1099 GND.n983 9.3005
R12206 GND.n1097 GND.n984 9.3005
R12207 GND.n1096 GND.n985 9.3005
R12208 GND.n1094 GND.n986 9.3005
R12209 GND.n1093 GND.n987 9.3005
R12210 GND.n1091 GND.n988 9.3005
R12211 GND.n1090 GND.n989 9.3005
R12212 GND.n1088 GND.n990 9.3005
R12213 GND.n1087 GND.n991 9.3005
R12214 GND.n1085 GND.n992 9.3005
R12215 GND.n1084 GND.n993 9.3005
R12216 GND.n1082 GND.n994 9.3005
R12217 GND.n1081 GND.n995 9.3005
R12218 GND.n1079 GND.n996 9.3005
R12219 GND.n1078 GND.n997 9.3005
R12220 GND.n1076 GND.n998 9.3005
R12221 GND.n1075 GND.n999 9.3005
R12222 GND.n1073 GND.n1000 9.3005
R12223 GND.n1072 GND.n1001 9.3005
R12224 GND.n1071 GND.n1002 9.3005
R12225 GND.n1069 GND.n1003 9.3005
R12226 GND.n1068 GND.n1004 9.3005
R12227 GND.n1066 GND.n1005 9.3005
R12228 GND.n1065 GND.n1006 9.3005
R12229 GND.n1063 GND.n1007 9.3005
R12230 GND.n1062 GND.n1008 9.3005
R12231 GND.n1060 GND.n1009 9.3005
R12232 GND.n1059 GND.n1010 9.3005
R12233 GND.n1057 GND.n1011 9.3005
R12234 GND.n1056 GND.n1012 9.3005
R12235 GND.n1036 GND.n1014 9.3005
R12236 GND.n1035 GND.n1015 9.3005
R12237 GND.n1033 GND.n1016 9.3005
R12238 GND.n1032 GND.n1017 9.3005
R12239 GND.n1030 GND.n1018 9.3005
R12240 GND.n1029 GND.n1019 9.3005
R12241 GND.n1027 GND.n1020 9.3005
R12242 GND.n1026 GND.n1021 9.3005
R12243 GND.n1024 GND.n1023 9.3005
R12244 GND.n1022 GND.n311 9.3005
R12245 GND.n7600 GND.n312 9.3005
R12246 GND.n7599 GND.n313 9.3005
R12247 GND.n7598 GND.n314 9.3005
R12248 GND.n333 GND.n315 9.3005
R12249 GND.n7588 GND.n334 9.3005
R12250 GND.n7587 GND.n335 9.3005
R12251 GND.n7586 GND.n336 9.3005
R12252 GND.n352 GND.n337 9.3005
R12253 GND.n7576 GND.n353 9.3005
R12254 GND.n7575 GND.n354 9.3005
R12255 GND.n7574 GND.n355 9.3005
R12256 GND.n371 GND.n356 9.3005
R12257 GND.n7564 GND.n372 9.3005
R12258 GND.n7563 GND.n373 9.3005
R12259 GND.n7562 GND.n374 9.3005
R12260 GND.n390 GND.n375 9.3005
R12261 GND.n7552 GND.n391 9.3005
R12262 GND.n7551 GND.n392 9.3005
R12263 GND.n7550 GND.n393 9.3005
R12264 GND.n409 GND.n394 9.3005
R12265 GND.n7540 GND.n410 9.3005
R12266 GND.n7539 GND.n411 9.3005
R12267 GND.n7538 GND.n412 9.3005
R12268 GND.n427 GND.n413 9.3005
R12269 GND.n7528 GND.n428 9.3005
R12270 GND.n7527 GND.n429 9.3005
R12271 GND.n7526 GND.n430 9.3005
R12272 GND.n447 GND.n431 9.3005
R12273 GND.n7516 GND.n448 9.3005
R12274 GND.n7515 GND.n449 9.3005
R12275 GND.n7514 GND.n450 9.3005
R12276 GND.n467 GND.n451 9.3005
R12277 GND.n7504 GND.n468 9.3005
R12278 GND.n7503 GND.n469 9.3005
R12279 GND.n7502 GND.n470 9.3005
R12280 GND.n486 GND.n471 9.3005
R12281 GND.n7492 GND.n487 9.3005
R12282 GND.n7491 GND.n488 9.3005
R12283 GND.n7490 GND.n489 9.3005
R12284 GND.n505 GND.n490 9.3005
R12285 GND.n7480 GND.n506 9.3005
R12286 GND.n7479 GND.n507 9.3005
R12287 GND.n7478 GND.n508 9.3005
R12288 GND.n524 GND.n509 9.3005
R12289 GND.n7468 GND.n525 9.3005
R12290 GND.n7467 GND.n7466 9.3005
R12291 GND.n1138 GND.n1137 9.3005
R12292 GND.n1052 GND.n246 9.3005
R12293 GND.n1038 GND.n246 9.3005
R12294 GND.n4302 GND.n4301 9.3005
R12295 GND.n4300 GND.n4082 9.3005
R12296 GND.n4299 GND.n4298 9.3005
R12297 GND.n4085 GND.n4084 9.3005
R12298 GND.n4292 GND.n4089 9.3005
R12299 GND.n4291 GND.n4090 9.3005
R12300 GND.n4290 GND.n4091 9.3005
R12301 GND.n4096 GND.n4092 9.3005
R12302 GND.n4284 GND.n4097 9.3005
R12303 GND.n4283 GND.n4098 9.3005
R12304 GND.n4282 GND.n4099 9.3005
R12305 GND.n4104 GND.n4100 9.3005
R12306 GND.n4276 GND.n4105 9.3005
R12307 GND.n4275 GND.n4106 9.3005
R12308 GND.n4274 GND.n4107 9.3005
R12309 GND.n4112 GND.n4108 9.3005
R12310 GND.n4268 GND.n4113 9.3005
R12311 GND.n4267 GND.n4114 9.3005
R12312 GND.n4266 GND.n4115 9.3005
R12313 GND.n4120 GND.n4116 9.3005
R12314 GND.n4260 GND.n4121 9.3005
R12315 GND.n4259 GND.n4122 9.3005
R12316 GND.n4258 GND.n4123 9.3005
R12317 GND.n4128 GND.n4124 9.3005
R12318 GND.n4252 GND.n4129 9.3005
R12319 GND.n4251 GND.n4130 9.3005
R12320 GND.n4250 GND.n4131 9.3005
R12321 GND.n4136 GND.n4132 9.3005
R12322 GND.n4244 GND.n4137 9.3005
R12323 GND.n4243 GND.n4138 9.3005
R12324 GND.n4242 GND.n4139 9.3005
R12325 GND.n4144 GND.n4140 9.3005
R12326 GND.n4236 GND.n4145 9.3005
R12327 GND.n4235 GND.n4146 9.3005
R12328 GND.n4234 GND.n4147 9.3005
R12329 GND.n4152 GND.n4148 9.3005
R12330 GND.n4228 GND.n4153 9.3005
R12331 GND.n4227 GND.n4154 9.3005
R12332 GND.n4226 GND.n4155 9.3005
R12333 GND.n4160 GND.n4156 9.3005
R12334 GND.n4220 GND.n4161 9.3005
R12335 GND.n4219 GND.n4162 9.3005
R12336 GND.n4218 GND.n4163 9.3005
R12337 GND.n4168 GND.n4164 9.3005
R12338 GND.n4212 GND.n4169 9.3005
R12339 GND.n4211 GND.n4170 9.3005
R12340 GND.n4210 GND.n4171 9.3005
R12341 GND.n4176 GND.n4172 9.3005
R12342 GND.n4204 GND.n4177 9.3005
R12343 GND.n4203 GND.n4178 9.3005
R12344 GND.n4202 GND.n4179 9.3005
R12345 GND.n4184 GND.n4180 9.3005
R12346 GND.n4196 GND.n4185 9.3005
R12347 GND.n4195 GND.n4186 9.3005
R12348 GND.n4194 GND.n4187 9.3005
R12349 GND.n4190 GND.n4189 9.3005
R12350 GND.n4083 GND.n4081 9.3005
R12351 GND.n4862 GND.n4861 9.3005
R12352 GND.n4860 GND.n3524 9.3005
R12353 GND.n3530 GND.n3525 9.3005
R12354 GND.n4854 GND.n3531 9.3005
R12355 GND.n4853 GND.n3532 9.3005
R12356 GND.n4852 GND.n3533 9.3005
R12357 GND.n3538 GND.n3534 9.3005
R12358 GND.n4846 GND.n3539 9.3005
R12359 GND.n4845 GND.n3540 9.3005
R12360 GND.n4844 GND.n3541 9.3005
R12361 GND.n3546 GND.n3542 9.3005
R12362 GND.n4838 GND.n3547 9.3005
R12363 GND.n4837 GND.n3548 9.3005
R12364 GND.n4836 GND.n3549 9.3005
R12365 GND.n3554 GND.n3550 9.3005
R12366 GND.n4830 GND.n3555 9.3005
R12367 GND.n4829 GND.n3556 9.3005
R12368 GND.n4828 GND.n3557 9.3005
R12369 GND.n3562 GND.n3558 9.3005
R12370 GND.n4822 GND.n3563 9.3005
R12371 GND.n4821 GND.n3564 9.3005
R12372 GND.n4820 GND.n3565 9.3005
R12373 GND.n3570 GND.n3566 9.3005
R12374 GND.n4814 GND.n3571 9.3005
R12375 GND.n4813 GND.n3572 9.3005
R12376 GND.n4812 GND.n3573 9.3005
R12377 GND.n3578 GND.n3574 9.3005
R12378 GND.n4806 GND.n3579 9.3005
R12379 GND.n4805 GND.n3580 9.3005
R12380 GND.n4804 GND.n3581 9.3005
R12381 GND.n3586 GND.n3582 9.3005
R12382 GND.n4798 GND.n3587 9.3005
R12383 GND.n4797 GND.n3588 9.3005
R12384 GND.n4796 GND.n3589 9.3005
R12385 GND.n3594 GND.n3590 9.3005
R12386 GND.n4790 GND.n3595 9.3005
R12387 GND.n4789 GND.n3596 9.3005
R12388 GND.n4788 GND.n3597 9.3005
R12389 GND.n3602 GND.n3598 9.3005
R12390 GND.n4782 GND.n3603 9.3005
R12391 GND.n4781 GND.n3604 9.3005
R12392 GND.n4780 GND.n3605 9.3005
R12393 GND.n3610 GND.n3606 9.3005
R12394 GND.n4774 GND.n3611 9.3005
R12395 GND.n4773 GND.n3612 9.3005
R12396 GND.n4772 GND.n3613 9.3005
R12397 GND.n3618 GND.n3614 9.3005
R12398 GND.n4766 GND.n3619 9.3005
R12399 GND.n4765 GND.n3620 9.3005
R12400 GND.n4764 GND.n3621 9.3005
R12401 GND.n3626 GND.n3622 9.3005
R12402 GND.n4758 GND.n3627 9.3005
R12403 GND.n4757 GND.n3628 9.3005
R12404 GND.n4756 GND.n3629 9.3005
R12405 GND.n3634 GND.n3630 9.3005
R12406 GND.n4750 GND.n3635 9.3005
R12407 GND.n4749 GND.n3636 9.3005
R12408 GND.n4748 GND.n3637 9.3005
R12409 GND.n3642 GND.n3638 9.3005
R12410 GND.n4742 GND.n3643 9.3005
R12411 GND.n4741 GND.n3644 9.3005
R12412 GND.n4740 GND.n3645 9.3005
R12413 GND.n3650 GND.n3646 9.3005
R12414 GND.n4734 GND.n3651 9.3005
R12415 GND.n4733 GND.n3652 9.3005
R12416 GND.n4732 GND.n3653 9.3005
R12417 GND.n3658 GND.n3654 9.3005
R12418 GND.n4726 GND.n3659 9.3005
R12419 GND.n4725 GND.n3660 9.3005
R12420 GND.n4724 GND.n3661 9.3005
R12421 GND.n3666 GND.n3662 9.3005
R12422 GND.n4718 GND.n3667 9.3005
R12423 GND.n4717 GND.n3668 9.3005
R12424 GND.n4716 GND.n3669 9.3005
R12425 GND.n3674 GND.n3670 9.3005
R12426 GND.n4710 GND.n3675 9.3005
R12427 GND.n4709 GND.n3676 9.3005
R12428 GND.n4708 GND.n3677 9.3005
R12429 GND.n3682 GND.n3678 9.3005
R12430 GND.n4702 GND.n3683 9.3005
R12431 GND.n4701 GND.n3684 9.3005
R12432 GND.n4700 GND.n3685 9.3005
R12433 GND.n3690 GND.n3686 9.3005
R12434 GND.n4694 GND.n3691 9.3005
R12435 GND.n4693 GND.n3692 9.3005
R12436 GND.n4692 GND.n3693 9.3005
R12437 GND.n3698 GND.n3694 9.3005
R12438 GND.n4686 GND.n3699 9.3005
R12439 GND.n4685 GND.n3700 9.3005
R12440 GND.n4684 GND.n3701 9.3005
R12441 GND.n3706 GND.n3702 9.3005
R12442 GND.n4678 GND.n3707 9.3005
R12443 GND.n4677 GND.n3708 9.3005
R12444 GND.n4676 GND.n3709 9.3005
R12445 GND.n3714 GND.n3710 9.3005
R12446 GND.n4670 GND.n3715 9.3005
R12447 GND.n4669 GND.n3716 9.3005
R12448 GND.n4668 GND.n3717 9.3005
R12449 GND.n3722 GND.n3718 9.3005
R12450 GND.n4662 GND.n3723 9.3005
R12451 GND.n4661 GND.n3724 9.3005
R12452 GND.n4660 GND.n3725 9.3005
R12453 GND.n3730 GND.n3726 9.3005
R12454 GND.n4654 GND.n3731 9.3005
R12455 GND.n4653 GND.n3732 9.3005
R12456 GND.n4652 GND.n3733 9.3005
R12457 GND.n3738 GND.n3734 9.3005
R12458 GND.n4646 GND.n3739 9.3005
R12459 GND.n4645 GND.n3740 9.3005
R12460 GND.n4644 GND.n3741 9.3005
R12461 GND.n3746 GND.n3742 9.3005
R12462 GND.n4638 GND.n3747 9.3005
R12463 GND.n4637 GND.n3748 9.3005
R12464 GND.n4636 GND.n3749 9.3005
R12465 GND.n3754 GND.n3750 9.3005
R12466 GND.n4630 GND.n3755 9.3005
R12467 GND.n4629 GND.n3756 9.3005
R12468 GND.n4628 GND.n3757 9.3005
R12469 GND.n3762 GND.n3758 9.3005
R12470 GND.n4622 GND.n3763 9.3005
R12471 GND.n4621 GND.n3764 9.3005
R12472 GND.n4620 GND.n3765 9.3005
R12473 GND.n3770 GND.n3766 9.3005
R12474 GND.n4614 GND.n3771 9.3005
R12475 GND.n4613 GND.n3772 9.3005
R12476 GND.n4612 GND.n3773 9.3005
R12477 GND.n3778 GND.n3774 9.3005
R12478 GND.n4606 GND.n3779 9.3005
R12479 GND.n4605 GND.n3780 9.3005
R12480 GND.n4604 GND.n3781 9.3005
R12481 GND.n3786 GND.n3782 9.3005
R12482 GND.n4598 GND.n3787 9.3005
R12483 GND.n4597 GND.n3788 9.3005
R12484 GND.n4596 GND.n3789 9.3005
R12485 GND.n3794 GND.n3790 9.3005
R12486 GND.n4590 GND.n3795 9.3005
R12487 GND.n4589 GND.n3796 9.3005
R12488 GND.n4588 GND.n3797 9.3005
R12489 GND.n3802 GND.n3798 9.3005
R12490 GND.n4582 GND.n3803 9.3005
R12491 GND.n4581 GND.n3804 9.3005
R12492 GND.n4580 GND.n3805 9.3005
R12493 GND.n3810 GND.n3806 9.3005
R12494 GND.n4574 GND.n3811 9.3005
R12495 GND.n4573 GND.n3812 9.3005
R12496 GND.n4572 GND.n3813 9.3005
R12497 GND.n3818 GND.n3814 9.3005
R12498 GND.n4566 GND.n3819 9.3005
R12499 GND.n4565 GND.n3820 9.3005
R12500 GND.n4564 GND.n3821 9.3005
R12501 GND.n3826 GND.n3822 9.3005
R12502 GND.n4558 GND.n3827 9.3005
R12503 GND.n4557 GND.n3828 9.3005
R12504 GND.n4556 GND.n3829 9.3005
R12505 GND.n3834 GND.n3830 9.3005
R12506 GND.n4550 GND.n3835 9.3005
R12507 GND.n4549 GND.n3836 9.3005
R12508 GND.n4548 GND.n3837 9.3005
R12509 GND.n3842 GND.n3838 9.3005
R12510 GND.n4542 GND.n3843 9.3005
R12511 GND.n4541 GND.n3844 9.3005
R12512 GND.n4540 GND.n3845 9.3005
R12513 GND.n3850 GND.n3846 9.3005
R12514 GND.n4534 GND.n3851 9.3005
R12515 GND.n4533 GND.n3852 9.3005
R12516 GND.n4532 GND.n3853 9.3005
R12517 GND.n3858 GND.n3854 9.3005
R12518 GND.n4526 GND.n3859 9.3005
R12519 GND.n4525 GND.n3860 9.3005
R12520 GND.n4524 GND.n3861 9.3005
R12521 GND.n3866 GND.n3862 9.3005
R12522 GND.n4518 GND.n3867 9.3005
R12523 GND.n4517 GND.n3868 9.3005
R12524 GND.n4516 GND.n3869 9.3005
R12525 GND.n3874 GND.n3870 9.3005
R12526 GND.n4510 GND.n3875 9.3005
R12527 GND.n4509 GND.n3876 9.3005
R12528 GND.n4508 GND.n3877 9.3005
R12529 GND.n3882 GND.n3878 9.3005
R12530 GND.n4502 GND.n3883 9.3005
R12531 GND.n4501 GND.n3884 9.3005
R12532 GND.n4500 GND.n3885 9.3005
R12533 GND.n3890 GND.n3886 9.3005
R12534 GND.n4494 GND.n3891 9.3005
R12535 GND.n4493 GND.n3892 9.3005
R12536 GND.n4492 GND.n3893 9.3005
R12537 GND.n3898 GND.n3894 9.3005
R12538 GND.n4486 GND.n3899 9.3005
R12539 GND.n4485 GND.n3900 9.3005
R12540 GND.n4484 GND.n3901 9.3005
R12541 GND.n3906 GND.n3902 9.3005
R12542 GND.n4478 GND.n3907 9.3005
R12543 GND.n4477 GND.n3908 9.3005
R12544 GND.n4476 GND.n3909 9.3005
R12545 GND.n3914 GND.n3910 9.3005
R12546 GND.n4470 GND.n3915 9.3005
R12547 GND.n4469 GND.n3916 9.3005
R12548 GND.n4468 GND.n3917 9.3005
R12549 GND.n3922 GND.n3918 9.3005
R12550 GND.n4462 GND.n3923 9.3005
R12551 GND.n4461 GND.n3924 9.3005
R12552 GND.n4460 GND.n3925 9.3005
R12553 GND.n3930 GND.n3926 9.3005
R12554 GND.n4454 GND.n3931 9.3005
R12555 GND.n4453 GND.n3932 9.3005
R12556 GND.n4452 GND.n3933 9.3005
R12557 GND.n3938 GND.n3934 9.3005
R12558 GND.n4446 GND.n3939 9.3005
R12559 GND.n4445 GND.n3940 9.3005
R12560 GND.n4444 GND.n3941 9.3005
R12561 GND.n3946 GND.n3942 9.3005
R12562 GND.n4438 GND.n3947 9.3005
R12563 GND.n4437 GND.n3948 9.3005
R12564 GND.n4436 GND.n3949 9.3005
R12565 GND.n3954 GND.n3950 9.3005
R12566 GND.n4430 GND.n3955 9.3005
R12567 GND.n4429 GND.n3956 9.3005
R12568 GND.n4428 GND.n3957 9.3005
R12569 GND.n3962 GND.n3958 9.3005
R12570 GND.n4422 GND.n3963 9.3005
R12571 GND.n4421 GND.n3964 9.3005
R12572 GND.n4420 GND.n3965 9.3005
R12573 GND.n3970 GND.n3966 9.3005
R12574 GND.n4414 GND.n3971 9.3005
R12575 GND.n4413 GND.n3972 9.3005
R12576 GND.n4412 GND.n3973 9.3005
R12577 GND.n3978 GND.n3974 9.3005
R12578 GND.n4406 GND.n3979 9.3005
R12579 GND.n4405 GND.n3980 9.3005
R12580 GND.n4404 GND.n3981 9.3005
R12581 GND.n3986 GND.n3982 9.3005
R12582 GND.n4398 GND.n3987 9.3005
R12583 GND.n4397 GND.n3988 9.3005
R12584 GND.n4396 GND.n3989 9.3005
R12585 GND.n3994 GND.n3990 9.3005
R12586 GND.n4390 GND.n3995 9.3005
R12587 GND.n4389 GND.n3996 9.3005
R12588 GND.n4388 GND.n3997 9.3005
R12589 GND.n4002 GND.n3998 9.3005
R12590 GND.n4382 GND.n4003 9.3005
R12591 GND.n4381 GND.n4004 9.3005
R12592 GND.n4380 GND.n4005 9.3005
R12593 GND.n4010 GND.n4006 9.3005
R12594 GND.n4374 GND.n4011 9.3005
R12595 GND.n4373 GND.n4012 9.3005
R12596 GND.n4372 GND.n4013 9.3005
R12597 GND.n4018 GND.n4014 9.3005
R12598 GND.n4366 GND.n4019 9.3005
R12599 GND.n4365 GND.n4020 9.3005
R12600 GND.n4364 GND.n4021 9.3005
R12601 GND.n4026 GND.n4022 9.3005
R12602 GND.n4358 GND.n4027 9.3005
R12603 GND.n4357 GND.n4028 9.3005
R12604 GND.n4356 GND.n4029 9.3005
R12605 GND.n4034 GND.n4030 9.3005
R12606 GND.n4350 GND.n4035 9.3005
R12607 GND.n4349 GND.n4036 9.3005
R12608 GND.n4348 GND.n4037 9.3005
R12609 GND.n4042 GND.n4038 9.3005
R12610 GND.n4342 GND.n4043 9.3005
R12611 GND.n4341 GND.n4044 9.3005
R12612 GND.n4340 GND.n4045 9.3005
R12613 GND.n4050 GND.n4046 9.3005
R12614 GND.n4334 GND.n4051 9.3005
R12615 GND.n4333 GND.n4052 9.3005
R12616 GND.n4332 GND.n4053 9.3005
R12617 GND.n4058 GND.n4054 9.3005
R12618 GND.n4326 GND.n4059 9.3005
R12619 GND.n4325 GND.n4060 9.3005
R12620 GND.n4324 GND.n4061 9.3005
R12621 GND.n4066 GND.n4062 9.3005
R12622 GND.n4318 GND.n4067 9.3005
R12623 GND.n4317 GND.n4068 9.3005
R12624 GND.n4316 GND.n4069 9.3005
R12625 GND.n4074 GND.n4070 9.3005
R12626 GND.n4310 GND.n4075 9.3005
R12627 GND.n4309 GND.n4076 9.3005
R12628 GND.n4308 GND.n4077 9.3005
R12629 GND.n5028 GND.n2787 9.3005
R12630 GND.n4916 GND.n2788 9.3005
R12631 GND.n4918 GND.n4917 9.3005
R12632 GND.n4921 GND.n4915 9.3005
R12633 GND.n4922 GND.n4914 9.3005
R12634 GND.n4925 GND.n4913 9.3005
R12635 GND.n4926 GND.n4912 9.3005
R12636 GND.n4929 GND.n4911 9.3005
R12637 GND.n4930 GND.n4910 9.3005
R12638 GND.n4933 GND.n4909 9.3005
R12639 GND.n4934 GND.n4908 9.3005
R12640 GND.n4937 GND.n4907 9.3005
R12641 GND.n4938 GND.n4906 9.3005
R12642 GND.n4941 GND.n4905 9.3005
R12643 GND.n4942 GND.n4904 9.3005
R12644 GND.n4945 GND.n4903 9.3005
R12645 GND.n4946 GND.n4902 9.3005
R12646 GND.n4949 GND.n4901 9.3005
R12647 GND.n4950 GND.n4900 9.3005
R12648 GND.n4953 GND.n4899 9.3005
R12649 GND.n4954 GND.n4898 9.3005
R12650 GND.n4957 GND.n4897 9.3005
R12651 GND.n4958 GND.n4896 9.3005
R12652 GND.n4961 GND.n4895 9.3005
R12653 GND.n4962 GND.n4894 9.3005
R12654 GND.n4965 GND.n4893 9.3005
R12655 GND.n4966 GND.n4892 9.3005
R12656 GND.n4969 GND.n4891 9.3005
R12657 GND.n4970 GND.n4890 9.3005
R12658 GND.n4973 GND.n4889 9.3005
R12659 GND.n4974 GND.n4888 9.3005
R12660 GND.n4977 GND.n4887 9.3005
R12661 GND.n4978 GND.n4886 9.3005
R12662 GND.n4981 GND.n4885 9.3005
R12663 GND.n4982 GND.n4884 9.3005
R12664 GND.n4985 GND.n4883 9.3005
R12665 GND.n4986 GND.n4882 9.3005
R12666 GND.n4989 GND.n4881 9.3005
R12667 GND.n4990 GND.n4880 9.3005
R12668 GND.n4993 GND.n4879 9.3005
R12669 GND.n4994 GND.n4878 9.3005
R12670 GND.n4997 GND.n4877 9.3005
R12671 GND.n4998 GND.n4876 9.3005
R12672 GND.n5001 GND.n4875 9.3005
R12673 GND.n5002 GND.n4874 9.3005
R12674 GND.n5005 GND.n4873 9.3005
R12675 GND.n5006 GND.n4872 9.3005
R12676 GND.n5009 GND.n4871 9.3005
R12677 GND.n5010 GND.n4870 9.3005
R12678 GND.n5013 GND.n4869 9.3005
R12679 GND.n5014 GND.n4868 9.3005
R12680 GND.n5017 GND.n4867 9.3005
R12681 GND.n5019 GND.n4866 9.3005
R12682 GND.n5020 GND.n4865 9.3005
R12683 GND.n5021 GND.n4864 9.3005
R12684 GND.n5022 GND.n4863 9.3005
R12685 GND.n5030 GND.n5029 9.3005
R12686 GND.n2769 GND.n2768 9.3005
R12687 GND.n5053 GND.n5052 9.3005
R12688 GND.n5054 GND.n2767 9.3005
R12689 GND.n5056 GND.n5055 9.3005
R12690 GND.n2537 GND.n2536 9.3005
R12691 GND.n5213 GND.n5212 9.3005
R12692 GND.n5214 GND.n2535 9.3005
R12693 GND.n5216 GND.n5215 9.3005
R12694 GND.n5218 GND.n2512 9.3005
R12695 GND.n5227 GND.n5226 9.3005
R12696 GND.n2493 GND.n2492 9.3005
R12697 GND.n5244 GND.n5243 9.3005
R12698 GND.n5245 GND.n2491 9.3005
R12699 GND.n5247 GND.n5246 9.3005
R12700 GND.n2473 GND.n2472 9.3005
R12701 GND.n5264 GND.n5263 9.3005
R12702 GND.n5265 GND.n2471 9.3005
R12703 GND.n5267 GND.n5266 9.3005
R12704 GND.n2452 GND.n2451 9.3005
R12705 GND.n5284 GND.n5283 9.3005
R12706 GND.n5285 GND.n2450 9.3005
R12707 GND.n5287 GND.n5286 9.3005
R12708 GND.n2433 GND.n2432 9.3005
R12709 GND.n5304 GND.n5303 9.3005
R12710 GND.n5305 GND.n2431 9.3005
R12711 GND.n5307 GND.n5306 9.3005
R12712 GND.n2413 GND.n2412 9.3005
R12713 GND.n5324 GND.n5323 9.3005
R12714 GND.n5325 GND.n2411 9.3005
R12715 GND.n5327 GND.n5326 9.3005
R12716 GND.n2392 GND.n2391 9.3005
R12717 GND.n5344 GND.n5343 9.3005
R12718 GND.n5345 GND.n2390 9.3005
R12719 GND.n5347 GND.n5346 9.3005
R12720 GND.n2373 GND.n2372 9.3005
R12721 GND.n5364 GND.n5363 9.3005
R12722 GND.n5365 GND.n2371 9.3005
R12723 GND.n5367 GND.n5366 9.3005
R12724 GND.n2353 GND.n2352 9.3005
R12725 GND.n5389 GND.n5388 9.3005
R12726 GND.n5390 GND.n2351 9.3005
R12727 GND.n5394 GND.n5391 9.3005
R12728 GND.n5393 GND.n5392 9.3005
R12729 GND.n2326 GND.n2325 9.3005
R12730 GND.n5469 GND.n5468 9.3005
R12731 GND.n5470 GND.n2324 9.3005
R12732 GND.n5472 GND.n5471 9.3005
R12733 GND.n2306 GND.n2305 9.3005
R12734 GND.n5489 GND.n5488 9.3005
R12735 GND.n5490 GND.n2304 9.3005
R12736 GND.n5492 GND.n5491 9.3005
R12737 GND.n2286 GND.n2285 9.3005
R12738 GND.n5509 GND.n5508 9.3005
R12739 GND.n5510 GND.n2284 9.3005
R12740 GND.n5512 GND.n5511 9.3005
R12741 GND.n2265 GND.n2264 9.3005
R12742 GND.n5529 GND.n5528 9.3005
R12743 GND.n5530 GND.n2263 9.3005
R12744 GND.n5532 GND.n5531 9.3005
R12745 GND.n2246 GND.n2245 9.3005
R12746 GND.n5553 GND.n5552 9.3005
R12747 GND.n5554 GND.n2244 9.3005
R12748 GND.n5557 GND.n5556 9.3005
R12749 GND.n5555 GND.n1744 9.3005
R12750 GND.n5689 GND.n1745 9.3005
R12751 GND.n5688 GND.n1746 9.3005
R12752 GND.n5687 GND.n1747 9.3005
R12753 GND.n1780 GND.n1748 9.3005
R12754 GND.n5681 GND.n1781 9.3005
R12755 GND.n5680 GND.n1782 9.3005
R12756 GND.n5679 GND.n1783 9.3005
R12757 GND.n1826 GND.n1784 9.3005
R12758 GND.n2179 GND.n1827 9.3005
R12759 GND.n2178 GND.n1828 9.3005
R12760 GND.n2177 GND.n1829 9.3005
R12761 GND.n1844 GND.n1830 9.3005
R12762 GND.n2165 GND.n1845 9.3005
R12763 GND.n2164 GND.n1846 9.3005
R12764 GND.n2163 GND.n1847 9.3005
R12765 GND.n1862 GND.n1848 9.3005
R12766 GND.n2151 GND.n1863 9.3005
R12767 GND.n2150 GND.n1864 9.3005
R12768 GND.n2149 GND.n1865 9.3005
R12769 GND.n1880 GND.n1866 9.3005
R12770 GND.n2137 GND.n1881 9.3005
R12771 GND.n2136 GND.n1882 9.3005
R12772 GND.n2135 GND.n1883 9.3005
R12773 GND.n1899 GND.n1884 9.3005
R12774 GND.n2123 GND.n1900 9.3005
R12775 GND.n2122 GND.n1901 9.3005
R12776 GND.n2121 GND.n1902 9.3005
R12777 GND.n1917 GND.n1903 9.3005
R12778 GND.n2109 GND.n1918 9.3005
R12779 GND.n2108 GND.n1919 9.3005
R12780 GND.n2107 GND.n1920 9.3005
R12781 GND.n1935 GND.n1921 9.3005
R12782 GND.n2095 GND.n1936 9.3005
R12783 GND.n2094 GND.n1937 9.3005
R12784 GND.n2093 GND.n1938 9.3005
R12785 GND.n1953 GND.n1939 9.3005
R12786 GND.n2081 GND.n1954 9.3005
R12787 GND.n2080 GND.n1955 9.3005
R12788 GND.n2079 GND.n1956 9.3005
R12789 GND.n1959 GND.n1957 9.3005
R12790 GND.n1963 GND.n1960 9.3005
R12791 GND.n1962 GND.n1961 9.3005
R12792 GND.n1700 GND.n1699 9.3005
R12793 GND.n5786 GND.n5785 9.3005
R12794 GND.n5787 GND.n1698 9.3005
R12795 GND.n5806 GND.n5788 9.3005
R12796 GND.n5805 GND.n5789 9.3005
R12797 GND.n5804 GND.n5790 9.3005
R12798 GND.n5793 GND.n5791 9.3005
R12799 GND.n5800 GND.n5794 9.3005
R12800 GND.n5799 GND.n5795 9.3005
R12801 GND.n5798 GND.n5797 9.3005
R12802 GND.n5796 GND.n1618 9.3005
R12803 GND.n1616 GND.n1615 9.3005
R12804 GND.n5911 GND.n5910 9.3005
R12805 GND.n5912 GND.n1614 9.3005
R12806 GND.n5914 GND.n5913 9.3005
R12807 GND.n1560 GND.n1559 9.3005
R12808 GND.n5989 GND.n5988 9.3005
R12809 GND.n5990 GND.n1558 9.3005
R12810 GND.n6003 GND.n5991 9.3005
R12811 GND.n6002 GND.n5992 9.3005
R12812 GND.n6001 GND.n5993 9.3005
R12813 GND.n5995 GND.n5994 9.3005
R12814 GND.n5997 GND.n5996 9.3005
R12815 GND.n1516 GND.n1515 9.3005
R12816 GND.n6079 GND.n6078 9.3005
R12817 GND.n6080 GND.n1514 9.3005
R12818 GND.n6084 GND.n6081 9.3005
R12819 GND.n6083 GND.n6082 9.3005
R12820 GND.n1481 GND.n1480 9.3005
R12821 GND.n6145 GND.n6144 9.3005
R12822 GND.n6146 GND.n1479 9.3005
R12823 GND.n6148 GND.n6147 9.3005
R12824 GND.n1457 GND.n1456 9.3005
R12825 GND.n6188 GND.n6187 9.3005
R12826 GND.n6189 GND.n1455 9.3005
R12827 GND.n6193 GND.n6190 9.3005
R12828 GND.n6192 GND.n6191 9.3005
R12829 GND.n1441 GND.n1440 9.3005
R12830 GND.n6248 GND.n6247 9.3005
R12831 GND.n6249 GND.n1439 9.3005
R12832 GND.n6251 GND.n6250 9.3005
R12833 GND.n1329 GND.n1328 9.3005
R12834 GND.n6320 GND.n6319 9.3005
R12835 GND.n6321 GND.n1327 9.3005
R12836 GND.n6328 GND.n6322 9.3005
R12837 GND.n6327 GND.n6323 9.3005
R12838 GND.n6326 GND.n6324 9.3005
R12839 GND.n1306 GND.n1305 9.3005
R12840 GND.n6360 GND.n6359 9.3005
R12841 GND.n6361 GND.n1304 9.3005
R12842 GND.n6374 GND.n6362 9.3005
R12843 GND.n6373 GND.n6363 9.3005
R12844 GND.n6372 GND.n6364 9.3005
R12845 GND.n6366 GND.n6365 9.3005
R12846 GND.n6368 GND.n6367 9.3005
R12847 GND.n1272 GND.n1271 9.3005
R12848 GND.n6418 GND.n6417 9.3005
R12849 GND.n6419 GND.n1270 9.3005
R12850 GND.n6423 GND.n6420 9.3005
R12851 GND.n6422 GND.n6421 9.3005
R12852 GND.n1247 GND.n1246 9.3005
R12853 GND.n6453 GND.n6452 9.3005
R12854 GND.n6454 GND.n1245 9.3005
R12855 GND.n6461 GND.n6455 9.3005
R12856 GND.n6460 GND.n6456 9.3005
R12857 GND.n6459 GND.n6457 9.3005
R12858 GND.n1222 GND.n1221 9.3005
R12859 GND.n6492 GND.n6491 9.3005
R12860 GND.n6493 GND.n1220 9.3005
R12861 GND.n6506 GND.n6494 9.3005
R12862 GND.n6505 GND.n6495 9.3005
R12863 GND.n6504 GND.n6496 9.3005
R12864 GND.n6498 GND.n6497 9.3005
R12865 GND.n6500 GND.n6499 9.3005
R12866 GND.n1188 GND.n1187 9.3005
R12867 GND.n6597 GND.n6596 9.3005
R12868 GND.n6598 GND.n1186 9.3005
R12869 GND.n6614 GND.n6599 9.3005
R12870 GND.n6613 GND.n6600 9.3005
R12871 GND.n6612 GND.n6601 9.3005
R12872 GND.n6604 GND.n6602 9.3005
R12873 GND.n6606 GND.n6605 9.3005
R12874 GND.n938 GND.n937 9.3005
R12875 GND.n6729 GND.n6728 9.3005
R12876 GND.n6730 GND.n936 9.3005
R12877 GND.n6732 GND.n6731 9.3005
R12878 GND.n916 GND.n915 9.3005
R12879 GND.n6755 GND.n6754 9.3005
R12880 GND.n6756 GND.n914 9.3005
R12881 GND.n6760 GND.n6757 9.3005
R12882 GND.n6759 GND.n6758 9.3005
R12883 GND.n889 GND.n888 9.3005
R12884 GND.n6866 GND.n6865 9.3005
R12885 GND.n6867 GND.n887 9.3005
R12886 GND.n6869 GND.n6868 9.3005
R12887 GND.n869 GND.n868 9.3005
R12888 GND.n6886 GND.n6885 9.3005
R12889 GND.n6887 GND.n867 9.3005
R12890 GND.n6889 GND.n6888 9.3005
R12891 GND.n849 GND.n848 9.3005
R12892 GND.n6906 GND.n6905 9.3005
R12893 GND.n6907 GND.n847 9.3005
R12894 GND.n6909 GND.n6908 9.3005
R12895 GND.n828 GND.n827 9.3005
R12896 GND.n6926 GND.n6925 9.3005
R12897 GND.n6927 GND.n826 9.3005
R12898 GND.n6929 GND.n6928 9.3005
R12899 GND.n809 GND.n808 9.3005
R12900 GND.n6946 GND.n6945 9.3005
R12901 GND.n6947 GND.n807 9.3005
R12902 GND.n6949 GND.n6948 9.3005
R12903 GND.n789 GND.n788 9.3005
R12904 GND.n6966 GND.n6965 9.3005
R12905 GND.n6967 GND.n787 9.3005
R12906 GND.n6969 GND.n6968 9.3005
R12907 GND.n769 GND.n768 9.3005
R12908 GND.n6986 GND.n6985 9.3005
R12909 GND.n6987 GND.n767 9.3005
R12910 GND.n6989 GND.n6988 9.3005
R12911 GND.n749 GND.n748 9.3005
R12912 GND.n7006 GND.n7005 9.3005
R12913 GND.n7007 GND.n747 9.3005
R12914 GND.n7009 GND.n7008 9.3005
R12915 GND.n728 GND.n727 9.3005
R12916 GND.n7030 GND.n7029 9.3005
R12917 GND.n7031 GND.n726 9.3005
R12918 GND.n7035 GND.n7032 9.3005
R12919 GND.n7034 GND.n7033 9.3005
R12920 GND.n701 GND.n700 9.3005
R12921 GND.n7074 GND.n7073 9.3005
R12922 GND.n7075 GND.n699 9.3005
R12923 GND.n7077 GND.n7076 9.3005
R12924 GND.n680 GND.n679 9.3005
R12925 GND.n7102 GND.n7101 9.3005
R12926 GND.n7103 GND.n678 9.3005
R12927 GND.n7105 GND.n7104 9.3005
R12928 GND.n651 GND.n650 9.3005
R12929 GND.n7138 GND.n7137 9.3005
R12930 GND.n7139 GND.n649 9.3005
R12931 GND.n7141 GND.n7140 9.3005
R12932 GND.n7143 GND.n242 9.3005
R12933 GND.n7635 GND.n7634 9.3005
R12934 GND.n249 GND.n247 9.3005
R12935 GND.n7624 GND.n270 9.3005
R12936 GND.n7623 GND.n271 9.3005
R12937 GND.n7622 GND.n272 9.3005
R12938 GND.n290 GND.n273 9.3005
R12939 GND.n7612 GND.n291 9.3005
R12940 GND.n7611 GND.n292 9.3005
R12941 GND.n7610 GND.n293 9.3005
R12942 GND.n4188 GND.n294 9.3005
R12943 GND.n5032 GND.n5031 9.3005
R12944 GND.n5225 GND.n2516 9.3005
R12945 GND.n5225 GND.n2511 9.3005
R12946 GND.n3143 GND.n3142 9.3005
R12947 GND.n3144 GND.n3083 9.3005
R12948 GND.n3082 GND.n3080 9.3005
R12949 GND.n3150 GND.n3079 9.3005
R12950 GND.n3151 GND.n3078 9.3005
R12951 GND.n3152 GND.n3077 9.3005
R12952 GND.n3076 GND.n3074 9.3005
R12953 GND.n3158 GND.n3073 9.3005
R12954 GND.n3159 GND.n3072 9.3005
R12955 GND.n3160 GND.n3071 9.3005
R12956 GND.n3070 GND.n3068 9.3005
R12957 GND.n3166 GND.n3065 9.3005
R12958 GND.n3167 GND.n3064 9.3005
R12959 GND.n3168 GND.n3063 9.3005
R12960 GND.n3062 GND.n3060 9.3005
R12961 GND.n3173 GND.n3059 9.3005
R12962 GND.n3174 GND.n3058 9.3005
R12963 GND.n3057 GND.n3055 9.3005
R12964 GND.n3179 GND.n3054 9.3005
R12965 GND.n3181 GND.n3180 9.3005
R12966 GND.n3141 GND.n3088 9.3005
R12967 GND.n3140 GND.n3139 9.3005
R12968 GND.n3037 GND.n3036 9.3005
R12969 GND.n3204 GND.n3203 9.3005
R12970 GND.n3205 GND.n3035 9.3005
R12971 GND.n3209 GND.n3206 9.3005
R12972 GND.n3208 GND.n3207 9.3005
R12973 GND.n3009 GND.n3008 9.3005
R12974 GND.n3336 GND.n3335 9.3005
R12975 GND.n3337 GND.n3007 9.3005
R12976 GND.n3339 GND.n3338 9.3005
R12977 GND.n2988 GND.n2987 9.3005
R12978 GND.n3353 GND.n3352 9.3005
R12979 GND.n3354 GND.n2986 9.3005
R12980 GND.n3356 GND.n3355 9.3005
R12981 GND.n2967 GND.n2966 9.3005
R12982 GND.n3370 GND.n3369 9.3005
R12983 GND.n3371 GND.n2965 9.3005
R12984 GND.n3373 GND.n3372 9.3005
R12985 GND.n2945 GND.n2944 9.3005
R12986 GND.n3387 GND.n3386 9.3005
R12987 GND.n3388 GND.n2943 9.3005
R12988 GND.n3390 GND.n3389 9.3005
R12989 GND.n2925 GND.n2924 9.3005
R12990 GND.n3404 GND.n3403 9.3005
R12991 GND.n3405 GND.n2923 9.3005
R12992 GND.n3407 GND.n3406 9.3005
R12993 GND.n2904 GND.n2903 9.3005
R12994 GND.n3421 GND.n3420 9.3005
R12995 GND.n3422 GND.n2902 9.3005
R12996 GND.n3424 GND.n3423 9.3005
R12997 GND.n2883 GND.n2882 9.3005
R12998 GND.n3438 GND.n3437 9.3005
R12999 GND.n3439 GND.n2881 9.3005
R13000 GND.n3441 GND.n3440 9.3005
R13001 GND.n2862 GND.n2861 9.3005
R13002 GND.n3455 GND.n3454 9.3005
R13003 GND.n3456 GND.n2860 9.3005
R13004 GND.n3458 GND.n3457 9.3005
R13005 GND.n2841 GND.n2840 9.3005
R13006 GND.n3472 GND.n3471 9.3005
R13007 GND.n3473 GND.n2839 9.3005
R13008 GND.n3475 GND.n3474 9.3005
R13009 GND.n2822 GND.n2821 9.3005
R13010 GND.n3495 GND.n3494 9.3005
R13011 GND.n3496 GND.n2820 9.3005
R13012 GND.n3518 GND.n3497 9.3005
R13013 GND.n3517 GND.n3498 9.3005
R13014 GND.n3516 GND.n3499 9.3005
R13015 GND.n3514 GND.n3500 9.3005
R13016 GND.n3513 GND.n3501 9.3005
R13017 GND.n3511 GND.n3502 9.3005
R13018 GND.n3510 GND.n3503 9.3005
R13019 GND.n3508 GND.n3504 9.3005
R13020 GND.n3507 GND.n3505 9.3005
R13021 GND.n2525 GND.n2524 9.3005
R13022 GND.n5223 GND.n5222 9.3005
R13023 GND.n2708 GND.n2518 9.3005
R13024 GND.n2707 GND.n2578 9.3005
R13025 GND.n2705 GND.n2579 9.3005
R13026 GND.n2704 GND.n2580 9.3005
R13027 GND.n2702 GND.n2581 9.3005
R13028 GND.n2701 GND.n2582 9.3005
R13029 GND.n2699 GND.n2583 9.3005
R13030 GND.n2698 GND.n2584 9.3005
R13031 GND.n2696 GND.n2585 9.3005
R13032 GND.n2695 GND.n2586 9.3005
R13033 GND.n2693 GND.n2587 9.3005
R13034 GND.n2692 GND.n2588 9.3005
R13035 GND.n2690 GND.n2589 9.3005
R13036 GND.n2689 GND.n2590 9.3005
R13037 GND.n2687 GND.n2591 9.3005
R13038 GND.n2686 GND.n2592 9.3005
R13039 GND.n2684 GND.n2593 9.3005
R13040 GND.n2683 GND.n2594 9.3005
R13041 GND.n2681 GND.n2595 9.3005
R13042 GND.n2680 GND.n2596 9.3005
R13043 GND.n2678 GND.n2597 9.3005
R13044 GND.n2677 GND.n2598 9.3005
R13045 GND.n2675 GND.n2599 9.3005
R13046 GND.n2674 GND.n2600 9.3005
R13047 GND.n2672 GND.n2601 9.3005
R13048 GND.n2671 GND.n2602 9.3005
R13049 GND.n2669 GND.n2603 9.3005
R13050 GND.n2668 GND.n2604 9.3005
R13051 GND.n2666 GND.n2605 9.3005
R13052 GND.n2665 GND.n2606 9.3005
R13053 GND.n2663 GND.n2607 9.3005
R13054 GND.n2662 GND.n2608 9.3005
R13055 GND.n2660 GND.n2609 9.3005
R13056 GND.n2659 GND.n2610 9.3005
R13057 GND.n2657 GND.n2611 9.3005
R13058 GND.n2656 GND.n2612 9.3005
R13059 GND.n2655 GND.n2613 9.3005
R13060 GND.n2653 GND.n2614 9.3005
R13061 GND.n2652 GND.n2615 9.3005
R13062 GND.n2650 GND.n2616 9.3005
R13063 GND.n2649 GND.n2617 9.3005
R13064 GND.n2647 GND.n2618 9.3005
R13065 GND.n2646 GND.n2619 9.3005
R13066 GND.n2644 GND.n2620 9.3005
R13067 GND.n2643 GND.n2621 9.3005
R13068 GND.n2641 GND.n2622 9.3005
R13069 GND.n2640 GND.n2623 9.3005
R13070 GND.n2638 GND.n2624 9.3005
R13071 GND.n2637 GND.n2625 9.3005
R13072 GND.n2635 GND.n2626 9.3005
R13073 GND.n2634 GND.n2627 9.3005
R13074 GND.n2632 GND.n2628 9.3005
R13075 GND.n2631 GND.n2630 9.3005
R13076 GND.n2629 GND.n2237 9.3005
R13077 GND.n5562 GND.n2236 9.3005
R13078 GND.n5564 GND.n5563 9.3005
R13079 GND.n3183 GND.n3182 9.3005
R13080 GND.n5087 GND.n2723 9.3005
R13081 GND.n5173 GND.n5088 9.3005
R13082 GND.n5172 GND.n5089 9.3005
R13083 GND.n5171 GND.n5090 9.3005
R13084 GND.n5170 GND.n5091 9.3005
R13085 GND.n5168 GND.n5092 9.3005
R13086 GND.n5167 GND.n5093 9.3005
R13087 GND.n5165 GND.n5094 9.3005
R13088 GND.n5164 GND.n5095 9.3005
R13089 GND.n5162 GND.n5096 9.3005
R13090 GND.n5161 GND.n5097 9.3005
R13091 GND.n5159 GND.n5098 9.3005
R13092 GND.n5158 GND.n5099 9.3005
R13093 GND.n5156 GND.n5100 9.3005
R13094 GND.n5155 GND.n5101 9.3005
R13095 GND.n5153 GND.n5102 9.3005
R13096 GND.n5152 GND.n5103 9.3005
R13097 GND.n5150 GND.n5104 9.3005
R13098 GND.n5149 GND.n5105 9.3005
R13099 GND.n5147 GND.n5106 9.3005
R13100 GND.n5146 GND.n5107 9.3005
R13101 GND.n5144 GND.n5108 9.3005
R13102 GND.n5143 GND.n5109 9.3005
R13103 GND.n5141 GND.n5110 9.3005
R13104 GND.n5140 GND.n5111 9.3005
R13105 GND.n5138 GND.n5112 9.3005
R13106 GND.n5137 GND.n5113 9.3005
R13107 GND.n5135 GND.n5114 9.3005
R13108 GND.n5134 GND.n5115 9.3005
R13109 GND.n5132 GND.n5116 9.3005
R13110 GND.n5131 GND.n5117 9.3005
R13111 GND.n5129 GND.n5118 9.3005
R13112 GND.n5128 GND.n5119 9.3005
R13113 GND.n5126 GND.n5120 9.3005
R13114 GND.n5125 GND.n5121 9.3005
R13115 GND.n5123 GND.n5122 9.3005
R13116 GND.n2343 GND.n2342 9.3005
R13117 GND.n5399 GND.n5398 9.3005
R13118 GND.n5400 GND.n2341 9.3005
R13119 GND.n5453 GND.n5401 9.3005
R13120 GND.n5452 GND.n5402 9.3005
R13121 GND.n5451 GND.n5403 9.3005
R13122 GND.n5449 GND.n5404 9.3005
R13123 GND.n5448 GND.n5405 9.3005
R13124 GND.n5446 GND.n5406 9.3005
R13125 GND.n5445 GND.n5407 9.3005
R13126 GND.n5443 GND.n5408 9.3005
R13127 GND.n5442 GND.n5409 9.3005
R13128 GND.n5440 GND.n5410 9.3005
R13129 GND.n5439 GND.n5411 9.3005
R13130 GND.n5437 GND.n5412 9.3005
R13131 GND.n5436 GND.n5413 9.3005
R13132 GND.n5434 GND.n5414 9.3005
R13133 GND.n5433 GND.n5415 9.3005
R13134 GND.n5431 GND.n5416 9.3005
R13135 GND.n5430 GND.n5417 9.3005
R13136 GND.n5428 GND.n5418 9.3005
R13137 GND.n5427 GND.n5419 9.3005
R13138 GND.n5425 GND.n5420 9.3005
R13139 GND.n5424 GND.n5421 9.3005
R13140 GND.n5422 GND.n1724 9.3005
R13141 GND.n5823 GND.n1679 9.3005
R13142 GND.n5826 GND.n5825 9.3005
R13143 GND.n5824 GND.n1680 9.3005
R13144 GND.n1653 GND.n1652 9.3005
R13145 GND.n5856 GND.n5855 9.3005
R13146 GND.n5857 GND.n1651 9.3005
R13147 GND.n5859 GND.n5858 9.3005
R13148 GND.n1625 GND.n1624 9.3005
R13149 GND.n5900 GND.n5899 9.3005
R13150 GND.n5901 GND.n1623 9.3005
R13151 GND.n5903 GND.n5902 9.3005
R13152 GND.n1583 GND.n1582 9.3005
R13153 GND.n5941 GND.n5940 9.3005
R13154 GND.n5942 GND.n1580 9.3005
R13155 GND.n5945 GND.n5944 9.3005
R13156 GND.n5943 GND.n1581 9.3005
R13157 GND.n1551 GND.n1550 9.3005
R13158 GND.n6009 GND.n6008 9.3005
R13159 GND.n6010 GND.n1549 9.3005
R13160 GND.n6012 GND.n6011 9.3005
R13161 GND.n1532 GND.n1531 9.3005
R13162 GND.n6061 GND.n6060 9.3005
R13163 GND.n6062 GND.n1529 9.3005
R13164 GND.n6065 GND.n6064 9.3005
R13165 GND.n6063 GND.n1530 9.3005
R13166 GND.n1500 GND.n1499 9.3005
R13167 GND.n6100 GND.n6099 9.3005
R13168 GND.n6101 GND.n1498 9.3005
R13169 GND.n6103 GND.n6102 9.3005
R13170 GND.n1473 GND.n1472 9.3005
R13171 GND.n6154 GND.n6153 9.3005
R13172 GND.n6155 GND.n1470 9.3005
R13173 GND.n6167 GND.n6166 9.3005
R13174 GND.n6165 GND.n1471 9.3005
R13175 GND.n6164 GND.n6163 9.3005
R13176 GND.n6162 GND.n6156 9.3005
R13177 GND.n6161 GND.n6160 9.3005
R13178 GND.n1425 GND.n1424 9.3005
R13179 GND.n6263 GND.n6262 9.3005
R13180 GND.n6264 GND.n1423 9.3005
R13181 GND.n6266 GND.n6265 9.3005
R13182 GND.n1338 GND.n1336 9.3005
R13183 GND.n6314 GND.n6313 9.3005
R13184 GND.n6312 GND.n1337 9.3005
R13185 GND.n5822 GND.n5821 9.3005
R13186 GND.n6309 GND.n1339 9.3005
R13187 GND.n6308 GND.n6307 9.3005
R13188 GND.n6306 GND.n1344 9.3005
R13189 GND.n6304 GND.n6303 9.3005
R13190 GND.n6302 GND.n1379 9.3005
R13191 GND.n6301 GND.n6300 9.3005
R13192 GND.n6299 GND.n1386 9.3005
R13193 GND.n6298 GND.n6297 9.3005
R13194 GND.n6296 GND.n1387 9.3005
R13195 GND.n6295 GND.n6294 9.3005
R13196 GND.n6293 GND.n1394 9.3005
R13197 GND.n6292 GND.n6291 9.3005
R13198 GND.n6290 GND.n1395 9.3005
R13199 GND.n6289 GND.n6288 9.3005
R13200 GND.n6287 GND.n1402 9.3005
R13201 GND.n6286 GND.n6285 9.3005
R13202 GND.n6283 GND.n1403 9.3005
R13203 GND.n6282 GND.n6281 9.3005
R13204 GND.n6280 GND.n1412 9.3005
R13205 GND.n6279 GND.n6278 9.3005
R13206 GND.n6311 GND.n6310 9.3005
R13207 GND.n1673 GND.n1672 9.3005
R13208 GND.n5831 GND.n5830 9.3005
R13209 GND.n5832 GND.n1670 9.3005
R13210 GND.n5836 GND.n5835 9.3005
R13211 GND.n5834 GND.n1671 9.3005
R13212 GND.n5833 GND.n1646 9.3005
R13213 GND.n5863 GND.n1645 9.3005
R13214 GND.n5865 GND.n5864 9.3005
R13215 GND.n5866 GND.n1643 9.3005
R13216 GND.n5876 GND.n5875 9.3005
R13217 GND.n5874 GND.n1644 9.3005
R13218 GND.n5873 GND.n5872 9.3005
R13219 GND.n5871 GND.n5867 9.3005
R13220 GND.n5870 GND.n5869 9.3005
R13221 GND.n5868 GND.n1575 9.3005
R13222 GND.n1573 GND.n1572 9.3005
R13223 GND.n5952 GND.n5951 9.3005
R13224 GND.n5953 GND.n1570 9.3005
R13225 GND.n5974 GND.n5973 9.3005
R13226 GND.n5972 GND.n1571 9.3005
R13227 GND.n5971 GND.n5970 9.3005
R13228 GND.n5969 GND.n5954 9.3005
R13229 GND.n5968 GND.n5967 9.3005
R13230 GND.n5966 GND.n5956 9.3005
R13231 GND.n5965 GND.n5964 9.3005
R13232 GND.n5963 GND.n5957 9.3005
R13233 GND.n5962 GND.n5961 9.3005
R13234 GND.n5960 GND.n1494 9.3005
R13235 GND.n6107 GND.n1493 9.3005
R13236 GND.n6109 GND.n6108 9.3005
R13237 GND.n6110 GND.n1491 9.3005
R13238 GND.n6130 GND.n6129 9.3005
R13239 GND.n6128 GND.n1492 9.3005
R13240 GND.n6127 GND.n6126 9.3005
R13241 GND.n6125 GND.n6111 9.3005
R13242 GND.n6124 GND.n6123 9.3005
R13243 GND.n6122 GND.n6115 9.3005
R13244 GND.n6121 GND.n6120 9.3005
R13245 GND.n6119 GND.n6116 9.3005
R13246 GND.n1418 GND.n1417 9.3005
R13247 GND.n6271 GND.n6270 9.3005
R13248 GND.n6272 GND.n1416 9.3005
R13249 GND.n6274 GND.n6273 9.3005
R13250 GND.n6275 GND.n1413 9.3005
R13251 GND.n5728 GND.n5727 9.3005
R13252 GND.n5731 GND.n5730 9.3005
R13253 GND.n5732 GND.n5721 9.3005
R13254 GND.n5734 GND.n5733 9.3005
R13255 GND.n5736 GND.n5735 9.3005
R13256 GND.n5737 GND.n5714 9.3005
R13257 GND.n5739 GND.n5738 9.3005
R13258 GND.n5740 GND.n5713 9.3005
R13259 GND.n5742 GND.n5741 9.3005
R13260 GND.n5743 GND.n5708 9.3005
R13261 GND.n5745 GND.n5744 9.3005
R13262 GND.n5746 GND.n5707 9.3005
R13263 GND.n5748 GND.n5747 9.3005
R13264 GND.n5749 GND.n5702 9.3005
R13265 GND.n5751 GND.n5750 9.3005
R13266 GND.n5752 GND.n5701 9.3005
R13267 GND.n5754 GND.n5753 9.3005
R13268 GND.n5756 GND.n5755 9.3005
R13269 GND.n5757 GND.n1723 9.3005
R13270 GND.n5759 GND.n5758 9.3005
R13271 GND.n1722 GND.n1681 9.3005
R13272 GND.n5729 GND.n5726 9.3005
R13273 GND.n5696 GND.n1730 9.3005
R13274 GND.n5580 GND.n2226 9.3005
R13275 GND.n5582 GND.n5581 9.3005
R13276 GND.n5579 GND.n2231 9.3005
R13277 GND.n5578 GND.n5577 9.3005
R13278 GND.n2233 GND.n2232 9.3005
R13279 GND.n5571 GND.n5570 9.3005
R13280 GND.n5569 GND.n2235 9.3005
R13281 GND.n5568 GND.n5567 9.3005
R13282 GND.n5629 GND.n5628 9.3005
R13283 GND.n5627 GND.n5589 9.3005
R13284 GND.n5626 GND.n5625 9.3005
R13285 GND.n5624 GND.n5590 9.3005
R13286 GND.n5623 GND.n5622 9.3005
R13287 GND.n5621 GND.n5597 9.3005
R13288 GND.n5620 GND.n5619 9.3005
R13289 GND.n5618 GND.n5598 9.3005
R13290 GND.n5617 GND.n5616 9.3005
R13291 GND.n5615 GND.n5605 9.3005
R13292 GND.n5614 GND.n5613 9.3005
R13293 GND.n5612 GND.n1731 9.3005
R13294 GND.n3046 GND.n3044 9.3005
R13295 GND.n3199 GND.n3198 9.3005
R13296 GND.n3047 GND.n3045 9.3005
R13297 GND.n3194 GND.n3190 9.3005
R13298 GND.n3193 GND.n3192 9.3005
R13299 GND.n3017 GND.n3015 9.3005
R13300 GND.n3331 GND.n3330 9.3005
R13301 GND.n3020 GND.n3016 9.3005
R13302 GND.n3019 GND.n3018 9.3005
R13303 GND.n2997 GND.n2995 9.3005
R13304 GND.n3348 GND.n3347 9.3005
R13305 GND.n3000 GND.n2996 9.3005
R13306 GND.n2999 GND.n2998 9.3005
R13307 GND.n2976 GND.n2974 9.3005
R13308 GND.n3365 GND.n3364 9.3005
R13309 GND.n2979 GND.n2975 9.3005
R13310 GND.n2978 GND.n2977 9.3005
R13311 GND.n2955 GND.n2953 9.3005
R13312 GND.n3382 GND.n3381 9.3005
R13313 GND.n2958 GND.n2954 9.3005
R13314 GND.n2957 GND.n2956 9.3005
R13315 GND.n2934 GND.n2932 9.3005
R13316 GND.n3399 GND.n3398 9.3005
R13317 GND.n2937 GND.n2933 9.3005
R13318 GND.n2936 GND.n2935 9.3005
R13319 GND.n2913 GND.n2911 9.3005
R13320 GND.n3416 GND.n3415 9.3005
R13321 GND.n2916 GND.n2912 9.3005
R13322 GND.n2915 GND.n2914 9.3005
R13323 GND.n2892 GND.n2890 9.3005
R13324 GND.n3433 GND.n3432 9.3005
R13325 GND.n2895 GND.n2891 9.3005
R13326 GND.n2894 GND.n2893 9.3005
R13327 GND.n2871 GND.n2869 9.3005
R13328 GND.n3450 GND.n3449 9.3005
R13329 GND.n2874 GND.n2870 9.3005
R13330 GND.n2873 GND.n2872 9.3005
R13331 GND.n2850 GND.n2848 9.3005
R13332 GND.n3467 GND.n3466 9.3005
R13333 GND.n2853 GND.n2849 9.3005
R13334 GND.n2852 GND.n2851 9.3005
R13335 GND.n2831 GND.n2829 9.3005
R13336 GND.n3490 GND.n3489 9.3005
R13337 GND.n2832 GND.n2830 9.3005
R13338 GND.n3483 GND.n3482 9.3005
R13339 GND.n3484 GND.n2780 9.3005
R13340 GND.n5037 GND.n2779 9.3005
R13341 GND.n5047 GND.n5038 9.3005
R13342 GND.n5046 GND.n5040 9.3005
R13343 GND.n5045 GND.n5043 9.3005
R13344 GND.n5042 GND.n2549 9.3005
R13345 GND.n5207 GND.n2550 9.3005
R13346 GND.n5206 GND.n2551 9.3005
R13347 GND.n5205 GND.n2552 9.3005
R13348 GND.n2557 GND.n2553 9.3005
R13349 GND.n5201 GND.n2558 9.3005
R13350 GND.n5200 GND.n2559 9.3005
R13351 GND.n5199 GND.n2560 9.3005
R13352 GND.n2747 GND.n2561 9.3005
R13353 GND.n5195 GND.n2566 9.3005
R13354 GND.n5194 GND.n2567 9.3005
R13355 GND.n5193 GND.n2568 9.3005
R13356 GND.n2575 GND.n2569 9.3005
R13357 GND.n5189 GND.n5184 9.3005
R13358 GND.n5188 GND.n5185 9.3005
R13359 GND.n5187 GND.n2504 9.3005
R13360 GND.n5232 GND.n2503 9.3005
R13361 GND.n5238 GND.n5233 9.3005
R13362 GND.n5237 GND.n5234 9.3005
R13363 GND.n5236 GND.n2484 9.3005
R13364 GND.n5252 GND.n2483 9.3005
R13365 GND.n5258 GND.n5253 9.3005
R13366 GND.n5257 GND.n5254 9.3005
R13367 GND.n5256 GND.n2464 9.3005
R13368 GND.n5272 GND.n2463 9.3005
R13369 GND.n5278 GND.n5273 9.3005
R13370 GND.n5277 GND.n5274 9.3005
R13371 GND.n5276 GND.n2444 9.3005
R13372 GND.n5292 GND.n2443 9.3005
R13373 GND.n5298 GND.n5293 9.3005
R13374 GND.n5297 GND.n5294 9.3005
R13375 GND.n5296 GND.n2424 9.3005
R13376 GND.n5312 GND.n2423 9.3005
R13377 GND.n5318 GND.n5313 9.3005
R13378 GND.n5317 GND.n5314 9.3005
R13379 GND.n5316 GND.n2404 9.3005
R13380 GND.n5332 GND.n2403 9.3005
R13381 GND.n5338 GND.n5333 9.3005
R13382 GND.n5337 GND.n5334 9.3005
R13383 GND.n5336 GND.n2384 9.3005
R13384 GND.n5352 GND.n2383 9.3005
R13385 GND.n5358 GND.n5353 9.3005
R13386 GND.n5357 GND.n5354 9.3005
R13387 GND.n5356 GND.n2364 9.3005
R13388 GND.n5372 GND.n2363 9.3005
R13389 GND.n5383 GND.n5373 9.3005
R13390 GND.n5382 GND.n5375 9.3005
R13391 GND.n5381 GND.n5376 9.3005
R13392 GND.n5377 GND.n2336 9.3005
R13393 GND.n5457 GND.n2335 9.3005
R13394 GND.n5463 GND.n5458 9.3005
R13395 GND.n5462 GND.n5459 9.3005
R13396 GND.n5461 GND.n2317 9.3005
R13397 GND.n5477 GND.n2316 9.3005
R13398 GND.n5483 GND.n5478 9.3005
R13399 GND.n5482 GND.n5479 9.3005
R13400 GND.n5481 GND.n2297 9.3005
R13401 GND.n5497 GND.n2296 9.3005
R13402 GND.n5503 GND.n5498 9.3005
R13403 GND.n5502 GND.n5499 9.3005
R13404 GND.n5501 GND.n2277 9.3005
R13405 GND.n5517 GND.n2276 9.3005
R13406 GND.n5523 GND.n5518 9.3005
R13407 GND.n5522 GND.n5519 9.3005
R13408 GND.n5521 GND.n2257 9.3005
R13409 GND.n5537 GND.n2256 9.3005
R13410 GND.n5547 GND.n5538 9.3005
R13411 GND.n5546 GND.n5540 9.3005
R13412 GND.n5545 GND.n5543 9.3005
R13413 GND.n5542 GND.n1732 9.3005
R13414 GND.n5694 GND.n1733 9.3005
R13415 GND.n3090 GND.n3089 9.3005
R13416 GND.n3188 GND.n3046 9.3005
R13417 GND.n3198 GND.n3197 9.3005
R13418 GND.n3196 GND.n3047 9.3005
R13419 GND.n3195 GND.n3194 9.3005
R13420 GND.n3193 GND.n3021 9.3005
R13421 GND.n3327 GND.n3017 9.3005
R13422 GND.n3330 GND.n3329 9.3005
R13423 GND.n3328 GND.n3020 9.3005
R13424 GND.n3019 GND.n3001 9.3005
R13425 GND.n3344 GND.n2997 9.3005
R13426 GND.n3347 GND.n3346 9.3005
R13427 GND.n3345 GND.n3000 9.3005
R13428 GND.n2999 GND.n2980 9.3005
R13429 GND.n3361 GND.n2976 9.3005
R13430 GND.n3364 GND.n3363 9.3005
R13431 GND.n3362 GND.n2979 9.3005
R13432 GND.n2978 GND.n2959 9.3005
R13433 GND.n3378 GND.n2955 9.3005
R13434 GND.n3381 GND.n3380 9.3005
R13435 GND.n3379 GND.n2958 9.3005
R13436 GND.n2957 GND.n2938 9.3005
R13437 GND.n3395 GND.n2934 9.3005
R13438 GND.n3398 GND.n3397 9.3005
R13439 GND.n3396 GND.n2937 9.3005
R13440 GND.n2936 GND.n2917 9.3005
R13441 GND.n3412 GND.n2913 9.3005
R13442 GND.n3415 GND.n3414 9.3005
R13443 GND.n3413 GND.n2916 9.3005
R13444 GND.n2915 GND.n2896 9.3005
R13445 GND.n3429 GND.n2892 9.3005
R13446 GND.n3432 GND.n3431 9.3005
R13447 GND.n3430 GND.n2895 9.3005
R13448 GND.n2894 GND.n2875 9.3005
R13449 GND.n3446 GND.n2871 9.3005
R13450 GND.n3449 GND.n3448 9.3005
R13451 GND.n3447 GND.n2874 9.3005
R13452 GND.n2873 GND.n2854 9.3005
R13453 GND.n3463 GND.n2850 9.3005
R13454 GND.n3466 GND.n3465 9.3005
R13455 GND.n3464 GND.n2853 9.3005
R13456 GND.n2852 GND.n2833 9.3005
R13457 GND.n3480 GND.n2831 9.3005
R13458 GND.n3489 GND.n3488 9.3005
R13459 GND.n3487 GND.n2832 9.3005
R13460 GND.n3486 GND.n3483 9.3005
R13461 GND.n3485 GND.n3484 9.3005
R13462 GND.n2779 GND.n2777 9.3005
R13463 GND.n5048 GND.n5047 9.3005
R13464 GND.n5046 GND.n2778 9.3005
R13465 GND.n5045 GND.n5044 9.3005
R13466 GND.n2549 GND.n2547 9.3005
R13467 GND.n5208 GND.n5207 9.3005
R13468 GND.n5206 GND.n2548 9.3005
R13469 GND.n5205 GND.n5204 9.3005
R13470 GND.n5203 GND.n2553 9.3005
R13471 GND.n5202 GND.n5201 9.3005
R13472 GND.n5200 GND.n2556 9.3005
R13473 GND.n5199 GND.n5198 9.3005
R13474 GND.n5197 GND.n2561 9.3005
R13475 GND.n5196 GND.n5195 9.3005
R13476 GND.n5194 GND.n2565 9.3005
R13477 GND.n5193 GND.n5192 9.3005
R13478 GND.n5191 GND.n2569 9.3005
R13479 GND.n5190 GND.n5189 9.3005
R13480 GND.n5188 GND.n2574 9.3005
R13481 GND.n5187 GND.n5186 9.3005
R13482 GND.n2503 GND.n2501 9.3005
R13483 GND.n5239 GND.n5238 9.3005
R13484 GND.n5237 GND.n2502 9.3005
R13485 GND.n5236 GND.n5235 9.3005
R13486 GND.n2483 GND.n2481 9.3005
R13487 GND.n5259 GND.n5258 9.3005
R13488 GND.n5257 GND.n2482 9.3005
R13489 GND.n5256 GND.n5255 9.3005
R13490 GND.n2463 GND.n2461 9.3005
R13491 GND.n5279 GND.n5278 9.3005
R13492 GND.n5277 GND.n2462 9.3005
R13493 GND.n5276 GND.n5275 9.3005
R13494 GND.n2443 GND.n2441 9.3005
R13495 GND.n5299 GND.n5298 9.3005
R13496 GND.n5297 GND.n2442 9.3005
R13497 GND.n5296 GND.n5295 9.3005
R13498 GND.n2423 GND.n2421 9.3005
R13499 GND.n5319 GND.n5318 9.3005
R13500 GND.n5317 GND.n2422 9.3005
R13501 GND.n5316 GND.n5315 9.3005
R13502 GND.n2403 GND.n2401 9.3005
R13503 GND.n5339 GND.n5338 9.3005
R13504 GND.n5337 GND.n2402 9.3005
R13505 GND.n5336 GND.n5335 9.3005
R13506 GND.n2383 GND.n2381 9.3005
R13507 GND.n5359 GND.n5358 9.3005
R13508 GND.n5357 GND.n2382 9.3005
R13509 GND.n5356 GND.n5355 9.3005
R13510 GND.n2363 GND.n2361 9.3005
R13511 GND.n5384 GND.n5383 9.3005
R13512 GND.n5382 GND.n2362 9.3005
R13513 GND.n5381 GND.n5380 9.3005
R13514 GND.n5379 GND.n5377 9.3005
R13515 GND.n2335 GND.n2333 9.3005
R13516 GND.n5464 GND.n5463 9.3005
R13517 GND.n5462 GND.n2334 9.3005
R13518 GND.n5461 GND.n5460 9.3005
R13519 GND.n2316 GND.n2314 9.3005
R13520 GND.n5484 GND.n5483 9.3005
R13521 GND.n5482 GND.n2315 9.3005
R13522 GND.n5481 GND.n5480 9.3005
R13523 GND.n2296 GND.n2294 9.3005
R13524 GND.n5504 GND.n5503 9.3005
R13525 GND.n5502 GND.n2295 9.3005
R13526 GND.n5501 GND.n5500 9.3005
R13527 GND.n2276 GND.n2274 9.3005
R13528 GND.n5524 GND.n5523 9.3005
R13529 GND.n5522 GND.n2275 9.3005
R13530 GND.n5521 GND.n5520 9.3005
R13531 GND.n2256 GND.n2254 9.3005
R13532 GND.n5548 GND.n5547 9.3005
R13533 GND.n5546 GND.n2255 9.3005
R13534 GND.n5545 GND.n5544 9.3005
R13535 GND.n1734 GND.n1732 9.3005
R13536 GND.n5694 GND.n5693 9.3005
R13537 GND.n3090 GND.n3048 9.3005
R13538 GND.n3122 GND.n3121 9.3005
R13539 GND.n3123 GND.n3101 9.3005
R13540 GND.n3125 GND.n3124 9.3005
R13541 GND.n3126 GND.n3095 9.3005
R13542 GND.n3128 GND.n3127 9.3005
R13543 GND.n3129 GND.n3094 9.3005
R13544 GND.n3131 GND.n3130 9.3005
R13545 GND.n3092 GND.n3091 9.3005
R13546 GND.n3137 GND.n3136 9.3005
R13547 GND.n3120 GND.n3102 9.3005
R13548 GND.n3114 GND.n3113 9.3005
R13549 GND.n3110 GND.n3106 9.3005
R13550 GND.n3109 GND.n3108 9.3005
R13551 GND.n3028 GND.n3027 9.3005
R13552 GND.n3214 GND.n3213 9.3005
R13553 GND.n3215 GND.n3025 9.3005
R13554 GND.n3323 GND.n3322 9.3005
R13555 GND.n3321 GND.n3026 9.3005
R13556 GND.n3320 GND.n3319 9.3005
R13557 GND.n3318 GND.n3216 9.3005
R13558 GND.n3317 GND.n3316 9.3005
R13559 GND.n3315 GND.n3219 9.3005
R13560 GND.n3314 GND.n3313 9.3005
R13561 GND.n3312 GND.n3220 9.3005
R13562 GND.n3311 GND.n3310 9.3005
R13563 GND.n3309 GND.n3223 9.3005
R13564 GND.n3308 GND.n3307 9.3005
R13565 GND.n3306 GND.n3224 9.3005
R13566 GND.n3305 GND.n3304 9.3005
R13567 GND.n3303 GND.n3227 9.3005
R13568 GND.n3302 GND.n3301 9.3005
R13569 GND.n3300 GND.n3228 9.3005
R13570 GND.n3299 GND.n3298 9.3005
R13571 GND.n3297 GND.n3231 9.3005
R13572 GND.n3296 GND.n3295 9.3005
R13573 GND.n3294 GND.n3232 9.3005
R13574 GND.n3293 GND.n3292 9.3005
R13575 GND.n3291 GND.n3235 9.3005
R13576 GND.n3290 GND.n3289 9.3005
R13577 GND.n3288 GND.n3236 9.3005
R13578 GND.n3287 GND.n3286 9.3005
R13579 GND.n3285 GND.n3239 9.3005
R13580 GND.n3284 GND.n3283 9.3005
R13581 GND.n3282 GND.n3240 9.3005
R13582 GND.n3281 GND.n3280 9.3005
R13583 GND.n3279 GND.n3243 9.3005
R13584 GND.n3278 GND.n3277 9.3005
R13585 GND.n3276 GND.n3244 9.3005
R13586 GND.n3275 GND.n3274 9.3005
R13587 GND.n3273 GND.n3247 9.3005
R13588 GND.n3272 GND.n3271 9.3005
R13589 GND.n3270 GND.n3248 9.3005
R13590 GND.n3269 GND.n3268 9.3005
R13591 GND.n3267 GND.n3251 9.3005
R13592 GND.n3266 GND.n3265 9.3005
R13593 GND.n3264 GND.n3252 9.3005
R13594 GND.n3263 GND.n3262 9.3005
R13595 GND.n3261 GND.n3255 9.3005
R13596 GND.n3260 GND.n3259 9.3005
R13597 GND.n3258 GND.n3257 9.3005
R13598 GND.n3256 GND.n2760 9.3005
R13599 GND.n5061 GND.n2759 9.3005
R13600 GND.n5063 GND.n5062 9.3005
R13601 GND.n5064 GND.n2753 9.3005
R13602 GND.n5066 GND.n5065 9.3005
R13603 GND.n5067 GND.n2752 9.3005
R13604 GND.n5070 GND.n5069 9.3005
R13605 GND.n5071 GND.n2751 9.3005
R13606 GND.n5073 GND.n5072 9.3005
R13607 GND.n2725 GND.n2724 9.3005
R13608 GND.n5085 GND.n5084 9.3005
R13609 GND.n3112 GND.n3111 9.3005
R13610 GND.n5819 GND.n5818 9.21838
R13611 GND.n5879 GND.n5878 9.21838
R13612 GND.n1605 GND.n1564 9.21838
R13613 GND.n6097 GND.n1502 9.21838
R13614 GND.n6176 GND.n1460 9.21838
R13615 GND.n6206 GND.n1321 9.21838
R13616 GND.n87 GND.n86 8.92171
R13617 GND.n108 GND.n107 8.92171
R13618 GND.n49 GND.n48 8.92171
R13619 GND.n70 GND.n69 8.92171
R13620 GND.n12 GND.n11 8.92171
R13621 GND.n33 GND.n32 8.92171
R13622 GND.n5630 GND.n2226 8.92171
R13623 GND.n6710 GND.n6709 8.92171
R13624 GND.n222 GND.n221 8.92171
R13625 GND.n201 GND.n200 8.92171
R13626 GND.n184 GND.n183 8.92171
R13627 GND.n163 GND.n162 8.92171
R13628 GND.n147 GND.n146 8.92171
R13629 GND.n126 GND.n125 8.92171
R13630 GND.n5809 GND.t38 8.8343
R13631 GND.n6268 GND.t79 8.8343
R13632 GND.n2175 GND.n1832 8.45022
R13633 GND.n1858 GND.n1857 8.45022
R13634 GND.n1913 GND.n1907 8.45022
R13635 GND.n2097 GND.n1933 8.45022
R13636 GND.n1694 GND.n1676 8.45022
R13637 GND.n5887 GND.n1635 8.45022
R13638 GND.n5977 GND.n1546 8.45022
R13639 GND.n6076 GND.n6075 8.45022
R13640 GND.n6237 GND.n6236 8.45022
R13641 GND.n6220 GND.n6212 8.45022
R13642 GND.n6389 GND.n1285 8.45022
R13643 GND.n6425 GND.n1260 8.45022
R13644 GND.n6515 GND.n1212 8.45022
R13645 GND.n6594 GND.n6593 8.45022
R13646 GND.n6576 GND.t70 8.45022
R13647 GND.n7646 GND.n7645 8.44769
R13648 GND.n5086 GND.n113 8.44769
R13649 GND.n83 GND.n77 8.14595
R13650 GND.n104 GND.n98 8.14595
R13651 GND.n45 GND.n39 8.14595
R13652 GND.n66 GND.n60 8.14595
R13653 GND.n8 GND.n2 8.14595
R13654 GND.n29 GND.n23 8.14595
R13655 GND.n218 GND.n212 8.14595
R13656 GND.n197 GND.n191 8.14595
R13657 GND.n180 GND.n174 8.14595
R13658 GND.n159 GND.n153 8.14595
R13659 GND.n143 GND.n137 8.14595
R13660 GND.n122 GND.n116 8.14595
R13661 GND.t2 GND.n6005 8.06614
R13662 GND.n6036 GND.t83 8.06614
R13663 GND.t7 GND.n1913 7.68206
R13664 GND.n5926 GND.n5925 7.68206
R13665 GND.n5947 GND.n1577 7.68206
R13666 GND.n6105 GND.n1496 7.68206
R13667 GND.n6133 GND.n6132 7.68206
R13668 GND.t4 GND.n6425 7.68206
R13669 GND.n82 GND.n79 7.3702
R13670 GND.n103 GND.n100 7.3702
R13671 GND.n44 GND.n41 7.3702
R13672 GND.n65 GND.n62 7.3702
R13673 GND.n7 GND.n4 7.3702
R13674 GND.n28 GND.n25 7.3702
R13675 GND.n217 GND.n214 7.3702
R13676 GND.n196 GND.n193 7.3702
R13677 GND.n179 GND.n176 7.3702
R13678 GND.n158 GND.n155 7.3702
R13679 GND.n142 GND.n139 7.3702
R13680 GND.n121 GND.n118 7.3702
R13681 GND.n74 GND.n36 7.25481
R13682 GND.n188 GND.n150 7.25481
R13683 GND.n3325 GND.t34 7.09422
R13684 GND.n2168 GND.n2167 6.91391
R13685 GND.n1993 GND.n1990 6.91391
R13686 GND.n2040 GND.n2037 6.91391
R13687 GND.n2105 GND.n2104 6.91391
R13688 GND.n5762 GND.n1705 6.91391
R13689 GND.n5839 GND.n1655 6.91391
R13690 GND.n1663 GND.n1658 6.91391
R13691 GND.t0 GND.n1662 6.91391
R13692 GND.n6050 GND.n1534 6.91391
R13693 GND.n6044 GND.n1537 6.91391
R13694 GND.t3 GND.n1445 6.91391
R13695 GND.n6229 GND.n1427 6.91391
R13696 GND.n6225 GND.n1430 6.91391
R13697 GND.n1325 GND.n1317 6.91391
R13698 GND.n6408 GND.n6407 6.91391
R13699 GND.n6415 GND.n6414 6.91391
R13700 GND.n6521 GND.n1201 6.91391
R13701 GND.n1202 GND.n1196 6.91391
R13702 GND.n6538 GND.n6534 6.5566
R13703 GND.n2221 GND.n1821 6.5566
R13704 GND.n5640 GND.n5639 6.5566
R13705 GND.n6628 GND.n6627 6.5566
R13706 GND.n5289 GND.t96 6.14575
R13707 GND.n5938 GND.n5937 6.14575
R13708 GND.n5918 GND.n5917 6.14575
R13709 GND.n6141 GND.n6140 6.14575
R13710 GND.n6151 GND.n1475 6.14575
R13711 GND.n7060 GND.t98 6.14575
R13712 GND.n7596 GND.t102 6.14575
R13713 GND.n90 GND.t104 5.87587
R13714 GND.n90 GND.t107 5.87587
R13715 GND.n92 GND.t114 5.87587
R13716 GND.n92 GND.t113 5.87587
R13717 GND.n94 GND.t128 5.87587
R13718 GND.n94 GND.t125 5.87587
R13719 GND.n52 GND.t97 5.87587
R13720 GND.n52 GND.t89 5.87587
R13721 GND.n54 GND.t149 5.87587
R13722 GND.n54 GND.t131 5.87587
R13723 GND.n56 GND.t133 5.87587
R13724 GND.n56 GND.t111 5.87587
R13725 GND.n15 GND.t136 5.87587
R13726 GND.n15 GND.t143 5.87587
R13727 GND.n17 GND.t87 5.87587
R13728 GND.n17 GND.t116 5.87587
R13729 GND.n19 GND.t106 5.87587
R13730 GND.n19 GND.t138 5.87587
R13731 GND.n208 GND.t137 5.87587
R13732 GND.n208 GND.t139 5.87587
R13733 GND.n206 GND.t127 5.87587
R13734 GND.n206 GND.t132 5.87587
R13735 GND.n204 GND.t118 5.87587
R13736 GND.n204 GND.t119 5.87587
R13737 GND.n170 GND.t147 5.87587
R13738 GND.n170 GND.t109 5.87587
R13739 GND.n168 GND.t101 5.87587
R13740 GND.n168 GND.t129 5.87587
R13741 GND.n166 GND.t124 5.87587
R13742 GND.n166 GND.t142 5.87587
R13743 GND.n133 GND.t103 5.87587
R13744 GND.n133 GND.t140 5.87587
R13745 GND.n131 GND.t148 5.87587
R13746 GND.n131 GND.t123 5.87587
R13747 GND.n129 GND.t134 5.87587
R13748 GND.n129 GND.t99 5.87587
R13749 GND.n83 GND.n82 5.81868
R13750 GND.n104 GND.n103 5.81868
R13751 GND.n45 GND.n44 5.81868
R13752 GND.n66 GND.n65 5.81868
R13753 GND.n8 GND.n7 5.81868
R13754 GND.n29 GND.n28 5.81868
R13755 GND.n218 GND.n217 5.81868
R13756 GND.n197 GND.n196 5.81868
R13757 GND.n180 GND.n179 5.81868
R13758 GND.n159 GND.n158 5.81868
R13759 GND.n143 GND.n142 5.81868
R13760 GND.n122 GND.n121 5.81868
R13761 GND.n6664 GND.t42 5.76167
R13762 GND.n7512 GND.n453 5.76167
R13763 GND.n5736 GND.n5720 5.62474
R13764 GND.n6285 GND.n6284 5.62474
R13765 GND.n6667 GND.n1147 5.62001
R13766 GND.n5632 GND.n2225 5.62001
R13767 GND.n5635 GND.n5632 5.62001
R13768 GND.n6667 GND.n1148 5.62001
R13769 GND.n1840 GND.n1834 5.3776
R13770 GND.n2161 GND.n1850 5.3776
R13771 GND.n2111 GND.n1915 5.3776
R13772 GND.n1931 GND.n1925 5.3776
R13773 GND.n5808 GND.n1668 5.3776
R13774 GND.n1663 GND.t0 5.3776
R13775 GND.n5847 GND.n1648 5.3776
R13776 GND.n6052 GND.n1541 5.3776
R13777 GND.n6069 GND.n6068 5.3776
R13778 GND.n6244 GND.n6243 5.3776
R13779 GND.n6229 GND.t3 5.3776
R13780 GND.n6254 GND.n6253 5.3776
R13781 GND.n1286 GND.n1280 5.3776
R13782 GND.n1276 GND.n1266 5.3776
R13783 GND.n6522 GND.n1206 5.3776
R13784 GND.n6587 GND.n6586 5.3776
R13785 GND.n86 GND.n77 5.04292
R13786 GND.n107 GND.n98 5.04292
R13787 GND.n48 GND.n39 5.04292
R13788 GND.n69 GND.n60 5.04292
R13789 GND.n11 GND.n2 5.04292
R13790 GND.n32 GND.n23 5.04292
R13791 GND.n221 GND.n212 5.04292
R13792 GND.n200 GND.n191 5.04292
R13793 GND.n183 GND.n174 5.04292
R13794 GND.n162 GND.n153 5.04292
R13795 GND.n146 GND.n137 5.04292
R13796 GND.n125 GND.n116 5.04292
R13797 GND.t5 GND.n5905 4.99352
R13798 GND.n6169 GND.t85 4.99352
R13799 GND.n111 GND.n95 4.98326
R13800 GND.n95 GND.n93 4.98326
R13801 GND.n93 GND.n91 4.98326
R13802 GND.n73 GND.n57 4.98326
R13803 GND.n57 GND.n55 4.98326
R13804 GND.n55 GND.n53 4.98326
R13805 GND.n36 GND.n20 4.98326
R13806 GND.n20 GND.n18 4.98326
R13807 GND.n18 GND.n16 4.98326
R13808 GND.n207 GND.n205 4.98326
R13809 GND.n209 GND.n207 4.98326
R13810 GND.n225 GND.n209 4.98326
R13811 GND.n169 GND.n167 4.98326
R13812 GND.n171 GND.n169 4.98326
R13813 GND.n187 GND.n171 4.98326
R13814 GND.n132 GND.n130 4.98326
R13815 GND.n134 GND.n132 4.98326
R13816 GND.n150 GND.n134 4.98326
R13817 GND.n112 GND.n111 4.94662
R13818 GND.n226 GND.n225 4.94662
R13819 GND.n74 GND.n73 4.88412
R13820 GND.n188 GND.n187 4.88412
R13821 GND.n1774 GND.n1726 4.74817
R13822 GND.n1773 GND.n1727 4.74817
R13823 GND.n1769 GND.n1728 4.74817
R13824 GND.n1765 GND.n1729 4.74817
R13825 GND.n1351 GND.n1350 4.74817
R13826 GND.n1356 GND.n1355 4.74817
R13827 GND.n1368 GND.n1361 4.74817
R13828 GND.n1365 GND.n1361 4.74817
R13829 GND.n1357 GND.n1356 4.74817
R13830 GND.n1352 GND.n1351 4.74817
R13831 GND.n1347 GND.n1346 4.74817
R13832 GND.n1055 GND.n1054 4.74817
R13833 GND.n1049 GND.n1048 4.74817
R13834 GND.n1045 GND.n1044 4.74817
R13835 GND.n1040 GND.n1039 4.74817
R13836 GND.n1054 GND.n1053 4.74817
R13837 GND.n1050 GND.n1049 4.74817
R13838 GND.n1046 GND.n1045 4.74817
R13839 GND.n1041 GND.n1040 4.74817
R13840 GND.n5217 GND.n2517 4.74817
R13841 GND.n5080 GND.n2515 4.74817
R13842 GND.n5177 GND.n2514 4.74817
R13843 GND.n5180 GND.n2513 4.74817
R13844 GND.n7162 GND.n245 4.74817
R13845 GND.n7166 GND.n244 4.74817
R13846 GND.n7639 GND.n240 4.74817
R13847 GND.n7637 GND.n241 4.74817
R13848 GND.n248 GND.n243 4.74817
R13849 GND.n7142 GND.n245 4.74817
R13850 GND.n7163 GND.n244 4.74817
R13851 GND.n7165 GND.n240 4.74817
R13852 GND.n7638 GND.n7637 4.74817
R13853 GND.n7206 GND.n243 4.74817
R13854 GND.n2734 GND.n2517 4.74817
R13855 GND.n5077 GND.n2515 4.74817
R13856 GND.n5079 GND.n2514 4.74817
R13857 GND.n5178 GND.n2513 4.74817
R13858 GND.n2742 GND.n2523 4.74817
R13859 GND.n2740 GND.n2522 4.74817
R13860 GND.n2729 GND.n2521 4.74817
R13861 GND.n2717 GND.n2520 4.74817
R13862 GND.n2709 GND.n2519 4.74817
R13863 GND.n2526 GND.n2523 4.74817
R13864 GND.n2743 GND.n2522 4.74817
R13865 GND.n2739 GND.n2521 4.74817
R13866 GND.n2728 GND.n2520 4.74817
R13867 GND.n2716 GND.n2519 4.74817
R13868 GND.n1770 GND.n1727 4.74817
R13869 GND.n1766 GND.n1728 4.74817
R13870 GND.n1762 GND.n1729 4.74817
R13871 GND.n6709 GND.n6669 4.6132
R13872 GND.n5630 GND.n2229 4.6132
R13873 GND.n5763 GND.n5762 4.60944
R13874 GND.n5905 GND.n1621 4.60944
R13875 GND.t82 GND.n1562 4.60944
R13876 GND.t1 GND.n6028 4.60944
R13877 GND.n6170 GND.n6169 4.60944
R13878 GND.n6337 GND.n1317 4.60944
R13879 GND.n87 GND.n75 4.26717
R13880 GND.n108 GND.n96 4.26717
R13881 GND.n49 GND.n37 4.26717
R13882 GND.n70 GND.n58 4.26717
R13883 GND.n12 GND.n0 4.26717
R13884 GND.n33 GND.n21 4.26717
R13885 GND.n222 GND.n210 4.26717
R13886 GND.n201 GND.n189 4.26717
R13887 GND.n184 GND.n172 4.26717
R13888 GND.n163 GND.n151 4.26717
R13889 GND.n147 GND.n135 4.26717
R13890 GND.n126 GND.n114 4.26717
R13891 GND.n6541 GND.n6534 4.05904
R13892 GND.n2218 GND.n1821 4.05904
R13893 GND.n5641 GND.n5640 4.05904
R13894 GND.n6629 GND.n6628 4.05904
R13895 GND.n1758 GND.n1725 4.02039
R13896 GND.n1761 GND.n1725 4.02039
R13897 GND.t13 GND.n1975 3.84128
R13898 GND.n2154 GND.n2153 3.84128
R13899 GND.n2119 GND.n2118 3.84128
R13900 GND.n2053 GND.n2050 3.84128
R13901 GND.n5783 GND.n1675 3.84128
R13902 GND.n5885 GND.n1627 3.84128
R13903 GND.n6005 GND.n1555 3.84128
R13904 GND.n6037 GND.n6036 3.84128
R13905 GND.n6196 GND.n6195 3.84128
R13906 GND.n6317 GND.n1331 3.84128
R13907 GND.n6390 GND.n1290 3.84128
R13908 GND.n6432 GND.n1262 3.84128
R13909 GND.n6508 GND.n1210 3.84128
R13910 GND.n1192 GND.n1182 3.84128
R13911 GND.n3492 GND.t110 3.78382
R13912 GND.n1370 GND.n1369 3.61653
R13913 GND.n112 GND.n74 3.46178
R13914 GND.n226 GND.n188 3.46178
R13915 GND.n7234 GND.n307 3.4572
R13916 GND.n5782 GND.n5781 3.07313
R13917 GND.n5897 GND.n5896 3.07313
R13918 GND.n6006 GND.n1553 3.07313
R13919 GND.n6087 GND.n1510 3.07313
R13920 GND.n6178 GND.n1453 3.07313
R13921 GND.n6316 GND.n1333 3.07313
R13922 GND.n81 GND.n80 2.88718
R13923 GND.n102 GND.n101 2.88718
R13924 GND.n43 GND.n42 2.88718
R13925 GND.n64 GND.n63 2.88718
R13926 GND.n6 GND.n5 2.88718
R13927 GND.n27 GND.n26 2.88718
R13928 GND.n216 GND.n215 2.88718
R13929 GND.n195 GND.n194 2.88718
R13930 GND.n178 GND.n177 2.88718
R13931 GND.n157 GND.n156 2.88718
R13932 GND.n141 GND.n140 2.88718
R13933 GND.n120 GND.n119 2.88718
R13934 GND.n1378 GND.n1370 2.84323
R13935 GND.n5696 GND.n1725 2.64131
R13936 GND.n2147 GND.n1868 2.30497
R13937 GND.n2125 GND.n1897 2.30497
R13938 GND.n1949 GND.n1943 2.30497
R13939 GND.n1706 GND.n1683 2.30497
R13940 GND.n5906 GND.n1619 2.30497
R13941 GND.n5986 GND.n5985 2.30497
R13942 GND.n6096 GND.n1505 2.30497
R13943 GND.n6185 GND.n6184 2.30497
R13944 GND.n6331 GND.n6330 2.30497
R13945 GND.n6376 GND.n1294 2.30497
R13946 GND.n6450 GND.n1249 2.30497
R13947 GND.n6489 GND.n6488 2.30497
R13948 GND.n1378 GND.n1361 2.27742
R13949 GND.n1378 GND.n1356 2.27742
R13950 GND.n1378 GND.n1351 2.27742
R13951 GND.n1378 GND.n1346 2.27742
R13952 GND.n1054 GND.n246 2.27742
R13953 GND.n1049 GND.n246 2.27742
R13954 GND.n1045 GND.n246 2.27742
R13955 GND.n1040 GND.n246 2.27742
R13956 GND.n7636 GND.n245 2.27742
R13957 GND.n7636 GND.n244 2.27742
R13958 GND.n7636 GND.n240 2.27742
R13959 GND.n7637 GND.n7636 2.27742
R13960 GND.n7636 GND.n243 2.27742
R13961 GND.n5225 GND.n2517 2.27742
R13962 GND.n5225 GND.n2515 2.27742
R13963 GND.n5225 GND.n2514 2.27742
R13964 GND.n5225 GND.n2513 2.27742
R13965 GND.n5224 GND.n2523 2.27742
R13966 GND.n5224 GND.n2522 2.27742
R13967 GND.n5224 GND.n2521 2.27742
R13968 GND.n5224 GND.n2520 2.27742
R13969 GND.n5224 GND.n2519 2.27742
R13970 GND.n5696 GND.n1726 2.27742
R13971 GND.n5696 GND.n1727 2.27742
R13972 GND.n5696 GND.n1728 2.27742
R13973 GND.n5696 GND.n1729 2.27742
R13974 GND.n5025 GND.n2790 2.12862
R13975 GND GND.n113 1.91967
R13976 GND GND.n7646 1.80224
R13977 GND.n5466 GND.t92 1.53681
R13978 GND.n1857 GND.t16 1.53681
R13979 GND.n5810 GND.n5809 1.53681
R13980 GND.n5861 GND.n1649 1.53681
R13981 GND.n6015 GND.n6014 1.53681
R13982 GND.n6067 GND.n1518 1.53681
R13983 GND.n6235 GND.n1443 1.53681
R13984 GND.n6268 GND.n1421 1.53681
R13985 GND.n1212 GND.t24 1.53681
R13986 GND.n6616 GND.t70 1.53681
R13987 GND.n833 GND.t120 1.53681
R13988 GND.n433 GND.t94 1.53681
R13989 GND.n5733 GND.n5720 0.970197
R13990 GND.n6284 GND.n6283 0.970197
R13991 GND.n2950 GND.t90 0.94633
R13992 GND.n2140 GND.n2139 0.768656
R13993 GND.n2133 GND.n2132 0.768656
R13994 GND.n2068 GND.n2063 0.768656
R13995 GND.n5764 GND.n1710 0.768656
R13996 GND.n5924 GND.n1585 0.768656
R13997 GND.n5916 GND.n1576 0.768656
R13998 GND.n6142 GND.n1483 0.768656
R13999 GND.n6150 GND.n1477 0.768656
R14000 GND.n6338 GND.n1313 0.768656
R14001 GND.n6357 GND.n6356 0.768656
R14002 GND.n6464 GND.n6463 0.768656
R14003 GND.n1236 GND.n1230 0.768656
R14004 GND.n7636 GND.n246 0.548875
R14005 GND.n5225 GND.n5224 0.548875
R14006 GND.n4189 GND.n4188 0.523366
R14007 GND.n4083 GND.n4077 0.523366
R14008 GND.n4863 GND.n4862 0.523366
R14009 GND.n5031 GND.n5030 0.523366
R14010 GND.n5568 GND.n5564 0.486781
R14011 GND.n7466 GND.n7465 0.486781
R14012 GND.n1139 GND.n1138 0.486781
R14013 GND.n3182 GND.n3181 0.486781
R14014 GND.n5822 GND.n1681 0.470012
R14015 GND.n6312 GND.n6311 0.470012
R14016 GND.n6279 GND.n1413 0.470012
R14017 GND.n5729 GND.n5728 0.470012
R14018 GND.n7325 GND.n7324 0.453244
R14019 GND.n3113 GND.n3112 0.453244
R14020 GND.n6305 GND.n1378 0.37441
R14021 GND.n5697 GND.n5696 0.37441
R14022 GND.n7424 GND.n7423 0.296232
R14023 GND.n6686 GND.n929 0.296232
R14024 GND.n3140 GND.n3138 0.296232
R14025 GND.n5695 GND.n1731 0.296232
R14026 GND.n7423 GND.n7346 0.262695
R14027 GND.n3138 GND.n3137 0.262695
R14028 GND.n1378 GND.n1377 0.253549
R14029 GND.n5696 GND.n1724 0.253549
R14030 GND.n6669 GND.n1146 0.229039
R14031 GND.n6672 GND.n6669 0.229039
R14032 GND.n5580 GND.n2229 0.229039
R14033 GND.n5628 GND.n2229 0.229039
R14034 GND.n88 GND.n76 0.155672
R14035 GND.n81 GND.n76 0.155672
R14036 GND.n109 GND.n97 0.155672
R14037 GND.n102 GND.n97 0.155672
R14038 GND.n50 GND.n38 0.155672
R14039 GND.n43 GND.n38 0.155672
R14040 GND.n71 GND.n59 0.155672
R14041 GND.n64 GND.n59 0.155672
R14042 GND.n13 GND.n1 0.155672
R14043 GND.n6 GND.n1 0.155672
R14044 GND.n34 GND.n22 0.155672
R14045 GND.n27 GND.n22 0.155672
R14046 GND.n223 GND.n211 0.155672
R14047 GND.n216 GND.n211 0.155672
R14048 GND.n202 GND.n190 0.155672
R14049 GND.n195 GND.n190 0.155672
R14050 GND.n185 GND.n173 0.155672
R14051 GND.n178 GND.n173 0.155672
R14052 GND.n164 GND.n152 0.155672
R14053 GND.n157 GND.n152 0.155672
R14054 GND.n148 GND.n136 0.155672
R14055 GND.n141 GND.n136 0.155672
R14056 GND.n127 GND.n115 0.155672
R14057 GND.n120 GND.n115 0.155672
R14058 GND.n2578 GND.n2518 0.152939
R14059 GND.n2579 GND.n2578 0.152939
R14060 GND.n2580 GND.n2579 0.152939
R14061 GND.n2581 GND.n2580 0.152939
R14062 GND.n2582 GND.n2581 0.152939
R14063 GND.n2583 GND.n2582 0.152939
R14064 GND.n2584 GND.n2583 0.152939
R14065 GND.n2585 GND.n2584 0.152939
R14066 GND.n2586 GND.n2585 0.152939
R14067 GND.n2587 GND.n2586 0.152939
R14068 GND.n2588 GND.n2587 0.152939
R14069 GND.n2589 GND.n2588 0.152939
R14070 GND.n2590 GND.n2589 0.152939
R14071 GND.n2591 GND.n2590 0.152939
R14072 GND.n2592 GND.n2591 0.152939
R14073 GND.n2593 GND.n2592 0.152939
R14074 GND.n2594 GND.n2593 0.152939
R14075 GND.n2595 GND.n2594 0.152939
R14076 GND.n2596 GND.n2595 0.152939
R14077 GND.n2597 GND.n2596 0.152939
R14078 GND.n2598 GND.n2597 0.152939
R14079 GND.n2599 GND.n2598 0.152939
R14080 GND.n2600 GND.n2599 0.152939
R14081 GND.n2601 GND.n2600 0.152939
R14082 GND.n2602 GND.n2601 0.152939
R14083 GND.n2603 GND.n2602 0.152939
R14084 GND.n2604 GND.n2603 0.152939
R14085 GND.n2605 GND.n2604 0.152939
R14086 GND.n2606 GND.n2605 0.152939
R14087 GND.n2607 GND.n2606 0.152939
R14088 GND.n2608 GND.n2607 0.152939
R14089 GND.n2609 GND.n2608 0.152939
R14090 GND.n2610 GND.n2609 0.152939
R14091 GND.n2611 GND.n2610 0.152939
R14092 GND.n2612 GND.n2611 0.152939
R14093 GND.n2613 GND.n2612 0.152939
R14094 GND.n2614 GND.n2613 0.152939
R14095 GND.n2615 GND.n2614 0.152939
R14096 GND.n2616 GND.n2615 0.152939
R14097 GND.n2617 GND.n2616 0.152939
R14098 GND.n2618 GND.n2617 0.152939
R14099 GND.n2619 GND.n2618 0.152939
R14100 GND.n2620 GND.n2619 0.152939
R14101 GND.n2621 GND.n2620 0.152939
R14102 GND.n2622 GND.n2621 0.152939
R14103 GND.n2623 GND.n2622 0.152939
R14104 GND.n2624 GND.n2623 0.152939
R14105 GND.n2625 GND.n2624 0.152939
R14106 GND.n2626 GND.n2625 0.152939
R14107 GND.n2627 GND.n2626 0.152939
R14108 GND.n2628 GND.n2627 0.152939
R14109 GND.n2630 GND.n2628 0.152939
R14110 GND.n2630 GND.n2629 0.152939
R14111 GND.n2629 GND.n2236 0.152939
R14112 GND.n5564 GND.n2236 0.152939
R14113 GND.n5226 GND.n2492 0.152939
R14114 GND.n5244 GND.n2492 0.152939
R14115 GND.n5245 GND.n5244 0.152939
R14116 GND.n5246 GND.n5245 0.152939
R14117 GND.n5246 GND.n2472 0.152939
R14118 GND.n5264 GND.n2472 0.152939
R14119 GND.n5265 GND.n5264 0.152939
R14120 GND.n5266 GND.n5265 0.152939
R14121 GND.n5266 GND.n2451 0.152939
R14122 GND.n5284 GND.n2451 0.152939
R14123 GND.n5285 GND.n5284 0.152939
R14124 GND.n5286 GND.n5285 0.152939
R14125 GND.n5286 GND.n2432 0.152939
R14126 GND.n5304 GND.n2432 0.152939
R14127 GND.n5305 GND.n5304 0.152939
R14128 GND.n5306 GND.n5305 0.152939
R14129 GND.n5306 GND.n2412 0.152939
R14130 GND.n5324 GND.n2412 0.152939
R14131 GND.n5325 GND.n5324 0.152939
R14132 GND.n5326 GND.n5325 0.152939
R14133 GND.n5326 GND.n2391 0.152939
R14134 GND.n5344 GND.n2391 0.152939
R14135 GND.n5345 GND.n5344 0.152939
R14136 GND.n5346 GND.n5345 0.152939
R14137 GND.n5346 GND.n2372 0.152939
R14138 GND.n5364 GND.n2372 0.152939
R14139 GND.n5365 GND.n5364 0.152939
R14140 GND.n5366 GND.n5365 0.152939
R14141 GND.n5366 GND.n2352 0.152939
R14142 GND.n5389 GND.n2352 0.152939
R14143 GND.n5390 GND.n5389 0.152939
R14144 GND.n5391 GND.n5390 0.152939
R14145 GND.n5392 GND.n5391 0.152939
R14146 GND.n5392 GND.n2325 0.152939
R14147 GND.n5469 GND.n2325 0.152939
R14148 GND.n5470 GND.n5469 0.152939
R14149 GND.n5471 GND.n5470 0.152939
R14150 GND.n5471 GND.n2305 0.152939
R14151 GND.n5489 GND.n2305 0.152939
R14152 GND.n5490 GND.n5489 0.152939
R14153 GND.n5491 GND.n5490 0.152939
R14154 GND.n5491 GND.n2285 0.152939
R14155 GND.n5509 GND.n2285 0.152939
R14156 GND.n5510 GND.n5509 0.152939
R14157 GND.n5511 GND.n5510 0.152939
R14158 GND.n5511 GND.n2264 0.152939
R14159 GND.n5529 GND.n2264 0.152939
R14160 GND.n5530 GND.n5529 0.152939
R14161 GND.n5531 GND.n5530 0.152939
R14162 GND.n5531 GND.n2245 0.152939
R14163 GND.n5553 GND.n2245 0.152939
R14164 GND.n5554 GND.n5553 0.152939
R14165 GND.n5556 GND.n5554 0.152939
R14166 GND.n5556 GND.n5555 0.152939
R14167 GND.n5555 GND.n1745 0.152939
R14168 GND.n1746 GND.n1745 0.152939
R14169 GND.n1747 GND.n1746 0.152939
R14170 GND.n1780 GND.n1747 0.152939
R14171 GND.n1781 GND.n1780 0.152939
R14172 GND.n1782 GND.n1781 0.152939
R14173 GND.n1783 GND.n1782 0.152939
R14174 GND.n1826 GND.n1783 0.152939
R14175 GND.n1827 GND.n1826 0.152939
R14176 GND.n1828 GND.n1827 0.152939
R14177 GND.n1829 GND.n1828 0.152939
R14178 GND.n1844 GND.n1829 0.152939
R14179 GND.n1845 GND.n1844 0.152939
R14180 GND.n1846 GND.n1845 0.152939
R14181 GND.n1847 GND.n1846 0.152939
R14182 GND.n1862 GND.n1847 0.152939
R14183 GND.n1863 GND.n1862 0.152939
R14184 GND.n1864 GND.n1863 0.152939
R14185 GND.n1865 GND.n1864 0.152939
R14186 GND.n1880 GND.n1865 0.152939
R14187 GND.n1881 GND.n1880 0.152939
R14188 GND.n1882 GND.n1881 0.152939
R14189 GND.n1883 GND.n1882 0.152939
R14190 GND.n1899 GND.n1883 0.152939
R14191 GND.n1900 GND.n1899 0.152939
R14192 GND.n1901 GND.n1900 0.152939
R14193 GND.n1902 GND.n1901 0.152939
R14194 GND.n1917 GND.n1902 0.152939
R14195 GND.n1918 GND.n1917 0.152939
R14196 GND.n1919 GND.n1918 0.152939
R14197 GND.n1920 GND.n1919 0.152939
R14198 GND.n1935 GND.n1920 0.152939
R14199 GND.n1936 GND.n1935 0.152939
R14200 GND.n1937 GND.n1936 0.152939
R14201 GND.n1938 GND.n1937 0.152939
R14202 GND.n1953 GND.n1938 0.152939
R14203 GND.n1954 GND.n1953 0.152939
R14204 GND.n1955 GND.n1954 0.152939
R14205 GND.n1956 GND.n1955 0.152939
R14206 GND.n1959 GND.n1956 0.152939
R14207 GND.n1960 GND.n1959 0.152939
R14208 GND.n1961 GND.n1960 0.152939
R14209 GND.n1961 GND.n1699 0.152939
R14210 GND.n5786 GND.n1699 0.152939
R14211 GND.n5787 GND.n5786 0.152939
R14212 GND.n5788 GND.n5787 0.152939
R14213 GND.n5789 GND.n5788 0.152939
R14214 GND.n5790 GND.n5789 0.152939
R14215 GND.n5793 GND.n5790 0.152939
R14216 GND.n5794 GND.n5793 0.152939
R14217 GND.n5795 GND.n5794 0.152939
R14218 GND.n5797 GND.n5795 0.152939
R14219 GND.n5797 GND.n5796 0.152939
R14220 GND.n5796 GND.n1615 0.152939
R14221 GND.n5911 GND.n1615 0.152939
R14222 GND.n5912 GND.n5911 0.152939
R14223 GND.n5913 GND.n5912 0.152939
R14224 GND.n5913 GND.n1559 0.152939
R14225 GND.n5989 GND.n1559 0.152939
R14226 GND.n5990 GND.n5989 0.152939
R14227 GND.n5991 GND.n5990 0.152939
R14228 GND.n5992 GND.n5991 0.152939
R14229 GND.n5993 GND.n5992 0.152939
R14230 GND.n5995 GND.n5993 0.152939
R14231 GND.n5996 GND.n5995 0.152939
R14232 GND.n5996 GND.n1515 0.152939
R14233 GND.n6079 GND.n1515 0.152939
R14234 GND.n6080 GND.n6079 0.152939
R14235 GND.n6081 GND.n6080 0.152939
R14236 GND.n6082 GND.n6081 0.152939
R14237 GND.n6082 GND.n1480 0.152939
R14238 GND.n6145 GND.n1480 0.152939
R14239 GND.n6146 GND.n6145 0.152939
R14240 GND.n6147 GND.n6146 0.152939
R14241 GND.n6147 GND.n1456 0.152939
R14242 GND.n6188 GND.n1456 0.152939
R14243 GND.n6189 GND.n6188 0.152939
R14244 GND.n6190 GND.n6189 0.152939
R14245 GND.n6191 GND.n6190 0.152939
R14246 GND.n6191 GND.n1440 0.152939
R14247 GND.n6248 GND.n1440 0.152939
R14248 GND.n6249 GND.n6248 0.152939
R14249 GND.n6250 GND.n6249 0.152939
R14250 GND.n6250 GND.n1328 0.152939
R14251 GND.n6320 GND.n1328 0.152939
R14252 GND.n6321 GND.n6320 0.152939
R14253 GND.n6322 GND.n6321 0.152939
R14254 GND.n6323 GND.n6322 0.152939
R14255 GND.n6324 GND.n6323 0.152939
R14256 GND.n6324 GND.n1305 0.152939
R14257 GND.n6360 GND.n1305 0.152939
R14258 GND.n6361 GND.n6360 0.152939
R14259 GND.n6362 GND.n6361 0.152939
R14260 GND.n6363 GND.n6362 0.152939
R14261 GND.n6364 GND.n6363 0.152939
R14262 GND.n6366 GND.n6364 0.152939
R14263 GND.n6367 GND.n6366 0.152939
R14264 GND.n6367 GND.n1271 0.152939
R14265 GND.n6418 GND.n1271 0.152939
R14266 GND.n6419 GND.n6418 0.152939
R14267 GND.n6420 GND.n6419 0.152939
R14268 GND.n6421 GND.n6420 0.152939
R14269 GND.n6421 GND.n1246 0.152939
R14270 GND.n6453 GND.n1246 0.152939
R14271 GND.n6454 GND.n6453 0.152939
R14272 GND.n6455 GND.n6454 0.152939
R14273 GND.n6456 GND.n6455 0.152939
R14274 GND.n6457 GND.n6456 0.152939
R14275 GND.n6457 GND.n1221 0.152939
R14276 GND.n6492 GND.n1221 0.152939
R14277 GND.n6493 GND.n6492 0.152939
R14278 GND.n6494 GND.n6493 0.152939
R14279 GND.n6495 GND.n6494 0.152939
R14280 GND.n6496 GND.n6495 0.152939
R14281 GND.n6498 GND.n6496 0.152939
R14282 GND.n6499 GND.n6498 0.152939
R14283 GND.n6499 GND.n1187 0.152939
R14284 GND.n6597 GND.n1187 0.152939
R14285 GND.n6598 GND.n6597 0.152939
R14286 GND.n6599 GND.n6598 0.152939
R14287 GND.n6600 GND.n6599 0.152939
R14288 GND.n6601 GND.n6600 0.152939
R14289 GND.n6604 GND.n6601 0.152939
R14290 GND.n6605 GND.n6604 0.152939
R14291 GND.n6605 GND.n937 0.152939
R14292 GND.n6729 GND.n937 0.152939
R14293 GND.n6730 GND.n6729 0.152939
R14294 GND.n6731 GND.n6730 0.152939
R14295 GND.n6731 GND.n915 0.152939
R14296 GND.n6755 GND.n915 0.152939
R14297 GND.n6756 GND.n6755 0.152939
R14298 GND.n6757 GND.n6756 0.152939
R14299 GND.n6758 GND.n6757 0.152939
R14300 GND.n6758 GND.n888 0.152939
R14301 GND.n6866 GND.n888 0.152939
R14302 GND.n6867 GND.n6866 0.152939
R14303 GND.n6868 GND.n6867 0.152939
R14304 GND.n6868 GND.n868 0.152939
R14305 GND.n6886 GND.n868 0.152939
R14306 GND.n6887 GND.n6886 0.152939
R14307 GND.n6888 GND.n6887 0.152939
R14308 GND.n6888 GND.n848 0.152939
R14309 GND.n6906 GND.n848 0.152939
R14310 GND.n6907 GND.n6906 0.152939
R14311 GND.n6908 GND.n6907 0.152939
R14312 GND.n6908 GND.n827 0.152939
R14313 GND.n6926 GND.n827 0.152939
R14314 GND.n6927 GND.n6926 0.152939
R14315 GND.n6928 GND.n6927 0.152939
R14316 GND.n6928 GND.n808 0.152939
R14317 GND.n6946 GND.n808 0.152939
R14318 GND.n6947 GND.n6946 0.152939
R14319 GND.n6948 GND.n6947 0.152939
R14320 GND.n6948 GND.n788 0.152939
R14321 GND.n6966 GND.n788 0.152939
R14322 GND.n6967 GND.n6966 0.152939
R14323 GND.n6968 GND.n6967 0.152939
R14324 GND.n6968 GND.n768 0.152939
R14325 GND.n6986 GND.n768 0.152939
R14326 GND.n6987 GND.n6986 0.152939
R14327 GND.n6988 GND.n6987 0.152939
R14328 GND.n6988 GND.n748 0.152939
R14329 GND.n7006 GND.n748 0.152939
R14330 GND.n7007 GND.n7006 0.152939
R14331 GND.n7008 GND.n7007 0.152939
R14332 GND.n7008 GND.n727 0.152939
R14333 GND.n7030 GND.n727 0.152939
R14334 GND.n7031 GND.n7030 0.152939
R14335 GND.n7032 GND.n7031 0.152939
R14336 GND.n7033 GND.n7032 0.152939
R14337 GND.n7033 GND.n700 0.152939
R14338 GND.n7074 GND.n700 0.152939
R14339 GND.n7075 GND.n7074 0.152939
R14340 GND.n7076 GND.n7075 0.152939
R14341 GND.n7076 GND.n679 0.152939
R14342 GND.n7102 GND.n679 0.152939
R14343 GND.n7103 GND.n7102 0.152939
R14344 GND.n7104 GND.n7103 0.152939
R14345 GND.n7104 GND.n650 0.152939
R14346 GND.n7138 GND.n650 0.152939
R14347 GND.n7139 GND.n7138 0.152939
R14348 GND.n7140 GND.n7139 0.152939
R14349 GND.n7140 GND.n242 0.152939
R14350 GND.n1015 GND.n1014 0.152939
R14351 GND.n1016 GND.n1015 0.152939
R14352 GND.n1017 GND.n1016 0.152939
R14353 GND.n1018 GND.n1017 0.152939
R14354 GND.n1019 GND.n1018 0.152939
R14355 GND.n1020 GND.n1019 0.152939
R14356 GND.n1021 GND.n1020 0.152939
R14357 GND.n1023 GND.n1021 0.152939
R14358 GND.n1023 GND.n1022 0.152939
R14359 GND.n1022 GND.n312 0.152939
R14360 GND.n313 GND.n312 0.152939
R14361 GND.n314 GND.n313 0.152939
R14362 GND.n333 GND.n314 0.152939
R14363 GND.n334 GND.n333 0.152939
R14364 GND.n335 GND.n334 0.152939
R14365 GND.n336 GND.n335 0.152939
R14366 GND.n352 GND.n336 0.152939
R14367 GND.n353 GND.n352 0.152939
R14368 GND.n354 GND.n353 0.152939
R14369 GND.n355 GND.n354 0.152939
R14370 GND.n371 GND.n355 0.152939
R14371 GND.n372 GND.n371 0.152939
R14372 GND.n373 GND.n372 0.152939
R14373 GND.n374 GND.n373 0.152939
R14374 GND.n390 GND.n374 0.152939
R14375 GND.n391 GND.n390 0.152939
R14376 GND.n392 GND.n391 0.152939
R14377 GND.n393 GND.n392 0.152939
R14378 GND.n409 GND.n393 0.152939
R14379 GND.n410 GND.n409 0.152939
R14380 GND.n411 GND.n410 0.152939
R14381 GND.n412 GND.n411 0.152939
R14382 GND.n427 GND.n412 0.152939
R14383 GND.n428 GND.n427 0.152939
R14384 GND.n429 GND.n428 0.152939
R14385 GND.n430 GND.n429 0.152939
R14386 GND.n447 GND.n430 0.152939
R14387 GND.n448 GND.n447 0.152939
R14388 GND.n449 GND.n448 0.152939
R14389 GND.n450 GND.n449 0.152939
R14390 GND.n467 GND.n450 0.152939
R14391 GND.n468 GND.n467 0.152939
R14392 GND.n469 GND.n468 0.152939
R14393 GND.n470 GND.n469 0.152939
R14394 GND.n486 GND.n470 0.152939
R14395 GND.n487 GND.n486 0.152939
R14396 GND.n488 GND.n487 0.152939
R14397 GND.n489 GND.n488 0.152939
R14398 GND.n505 GND.n489 0.152939
R14399 GND.n506 GND.n505 0.152939
R14400 GND.n507 GND.n506 0.152939
R14401 GND.n508 GND.n507 0.152939
R14402 GND.n524 GND.n508 0.152939
R14403 GND.n525 GND.n524 0.152939
R14404 GND.n7466 GND.n525 0.152939
R14405 GND.n1377 GND.n1371 0.152939
R14406 GND.n1373 GND.n1371 0.152939
R14407 GND.n1373 GND.n905 0.152939
R14408 GND.n6765 GND.n905 0.152939
R14409 GND.n6766 GND.n6765 0.152939
R14410 GND.n6767 GND.n6766 0.152939
R14411 GND.n6768 GND.n6767 0.152939
R14412 GND.n6769 GND.n6768 0.152939
R14413 GND.n6770 GND.n6769 0.152939
R14414 GND.n6771 GND.n6770 0.152939
R14415 GND.n6772 GND.n6771 0.152939
R14416 GND.n6773 GND.n6772 0.152939
R14417 GND.n6774 GND.n6773 0.152939
R14418 GND.n6775 GND.n6774 0.152939
R14419 GND.n6776 GND.n6775 0.152939
R14420 GND.n6777 GND.n6776 0.152939
R14421 GND.n6778 GND.n6777 0.152939
R14422 GND.n6779 GND.n6778 0.152939
R14423 GND.n6780 GND.n6779 0.152939
R14424 GND.n6781 GND.n6780 0.152939
R14425 GND.n6782 GND.n6781 0.152939
R14426 GND.n6783 GND.n6782 0.152939
R14427 GND.n6784 GND.n6783 0.152939
R14428 GND.n6785 GND.n6784 0.152939
R14429 GND.n6786 GND.n6785 0.152939
R14430 GND.n6787 GND.n6786 0.152939
R14431 GND.n6788 GND.n6787 0.152939
R14432 GND.n6789 GND.n6788 0.152939
R14433 GND.n6790 GND.n6789 0.152939
R14434 GND.n6791 GND.n6790 0.152939
R14435 GND.n6792 GND.n6791 0.152939
R14436 GND.n6793 GND.n6792 0.152939
R14437 GND.n6794 GND.n6793 0.152939
R14438 GND.n6795 GND.n6794 0.152939
R14439 GND.n6796 GND.n6795 0.152939
R14440 GND.n6797 GND.n6796 0.152939
R14441 GND.n6798 GND.n6797 0.152939
R14442 GND.n6799 GND.n6798 0.152939
R14443 GND.n6800 GND.n6799 0.152939
R14444 GND.n6800 GND.n717 0.152939
R14445 GND.n7040 GND.n717 0.152939
R14446 GND.n7041 GND.n7040 0.152939
R14447 GND.n7042 GND.n7041 0.152939
R14448 GND.n7043 GND.n7042 0.152939
R14449 GND.n7044 GND.n7043 0.152939
R14450 GND.n7045 GND.n7044 0.152939
R14451 GND.n7046 GND.n7045 0.152939
R14452 GND.n7047 GND.n7046 0.152939
R14453 GND.n7049 GND.n7047 0.152939
R14454 GND.n7049 GND.n7048 0.152939
R14455 GND.n7048 GND.n670 0.152939
R14456 GND.n7112 GND.n670 0.152939
R14457 GND.n7113 GND.n7112 0.152939
R14458 GND.n7114 GND.n7113 0.152939
R14459 GND.n7115 GND.n7114 0.152939
R14460 GND.n7116 GND.n7115 0.152939
R14461 GND.n7117 GND.n7116 0.152939
R14462 GND.n7118 GND.n7117 0.152939
R14463 GND.n7119 GND.n7118 0.152939
R14464 GND.n7119 GND.n227 0.152939
R14465 GND.n7644 GND.n228 0.152939
R14466 GND.n616 GND.n228 0.152939
R14467 GND.n616 GND.n614 0.152939
R14468 GND.n7212 GND.n614 0.152939
R14469 GND.n7213 GND.n7212 0.152939
R14470 GND.n7214 GND.n7213 0.152939
R14471 GND.n7214 GND.n612 0.152939
R14472 GND.n7220 GND.n612 0.152939
R14473 GND.n7221 GND.n7220 0.152939
R14474 GND.n7222 GND.n7221 0.152939
R14475 GND.n7222 GND.n610 0.152939
R14476 GND.n7228 GND.n610 0.152939
R14477 GND.n7229 GND.n7228 0.152939
R14478 GND.n7230 GND.n7229 0.152939
R14479 GND.n7230 GND.n608 0.152939
R14480 GND.n7237 GND.n608 0.152939
R14481 GND.n7238 GND.n7237 0.152939
R14482 GND.n7239 GND.n7238 0.152939
R14483 GND.n7239 GND.n606 0.152939
R14484 GND.n7245 GND.n606 0.152939
R14485 GND.n7246 GND.n7245 0.152939
R14486 GND.n7247 GND.n7246 0.152939
R14487 GND.n7247 GND.n604 0.152939
R14488 GND.n7253 GND.n604 0.152939
R14489 GND.n7254 GND.n7253 0.152939
R14490 GND.n7255 GND.n7254 0.152939
R14491 GND.n7255 GND.n602 0.152939
R14492 GND.n7261 GND.n602 0.152939
R14493 GND.n7262 GND.n7261 0.152939
R14494 GND.n7263 GND.n7262 0.152939
R14495 GND.n7263 GND.n600 0.152939
R14496 GND.n7269 GND.n600 0.152939
R14497 GND.n7270 GND.n7269 0.152939
R14498 GND.n7271 GND.n7270 0.152939
R14499 GND.n7271 GND.n598 0.152939
R14500 GND.n7277 GND.n598 0.152939
R14501 GND.n7278 GND.n7277 0.152939
R14502 GND.n7279 GND.n7278 0.152939
R14503 GND.n7279 GND.n596 0.152939
R14504 GND.n7285 GND.n596 0.152939
R14505 GND.n7286 GND.n7285 0.152939
R14506 GND.n7287 GND.n7286 0.152939
R14507 GND.n7287 GND.n594 0.152939
R14508 GND.n7293 GND.n594 0.152939
R14509 GND.n7294 GND.n7293 0.152939
R14510 GND.n7295 GND.n7294 0.152939
R14511 GND.n7295 GND.n592 0.152939
R14512 GND.n7301 GND.n592 0.152939
R14513 GND.n7302 GND.n7301 0.152939
R14514 GND.n7303 GND.n7302 0.152939
R14515 GND.n7303 GND.n590 0.152939
R14516 GND.n7309 GND.n590 0.152939
R14517 GND.n7310 GND.n7309 0.152939
R14518 GND.n7311 GND.n7310 0.152939
R14519 GND.n7311 GND.n588 0.152939
R14520 GND.n7317 GND.n588 0.152939
R14521 GND.n7318 GND.n7317 0.152939
R14522 GND.n7319 GND.n7318 0.152939
R14523 GND.n7319 GND.n586 0.152939
R14524 GND.n7324 GND.n586 0.152939
R14525 GND.n7346 GND.n567 0.152939
R14526 GND.n570 GND.n567 0.152939
R14527 GND.n571 GND.n570 0.152939
R14528 GND.n572 GND.n571 0.152939
R14529 GND.n576 GND.n572 0.152939
R14530 GND.n577 GND.n576 0.152939
R14531 GND.n578 GND.n577 0.152939
R14532 GND.n579 GND.n578 0.152939
R14533 GND.n585 GND.n579 0.152939
R14534 GND.n7325 GND.n585 0.152939
R14535 GND.n7465 GND.n526 0.152939
R14536 GND.n531 GND.n526 0.152939
R14537 GND.n532 GND.n531 0.152939
R14538 GND.n533 GND.n532 0.152939
R14539 GND.n534 GND.n533 0.152939
R14540 GND.n538 GND.n534 0.152939
R14541 GND.n539 GND.n538 0.152939
R14542 GND.n540 GND.n539 0.152939
R14543 GND.n7447 GND.n540 0.152939
R14544 GND.n7447 GND.n7446 0.152939
R14545 GND.n7446 GND.n7445 0.152939
R14546 GND.n7445 GND.n546 0.152939
R14547 GND.n551 GND.n546 0.152939
R14548 GND.n552 GND.n551 0.152939
R14549 GND.n553 GND.n552 0.152939
R14550 GND.n557 GND.n553 0.152939
R14551 GND.n558 GND.n557 0.152939
R14552 GND.n559 GND.n558 0.152939
R14553 GND.n560 GND.n559 0.152939
R14554 GND.n566 GND.n560 0.152939
R14555 GND.n7424 GND.n566 0.152939
R14556 GND.n1140 GND.n1139 0.152939
R14557 GND.n1141 GND.n1140 0.152939
R14558 GND.n1142 GND.n1141 0.152939
R14559 GND.n1143 GND.n1142 0.152939
R14560 GND.n1144 GND.n1143 0.152939
R14561 GND.n1145 GND.n1144 0.152939
R14562 GND.n1146 GND.n1145 0.152939
R14563 GND.n6673 GND.n6672 0.152939
R14564 GND.n6674 GND.n6673 0.152939
R14565 GND.n6675 GND.n6674 0.152939
R14566 GND.n6676 GND.n6675 0.152939
R14567 GND.n6677 GND.n6676 0.152939
R14568 GND.n6678 GND.n6677 0.152939
R14569 GND.n6679 GND.n6678 0.152939
R14570 GND.n6680 GND.n6679 0.152939
R14571 GND.n6688 GND.n6680 0.152939
R14572 GND.n6688 GND.n6687 0.152939
R14573 GND.n6687 GND.n6686 0.152939
R14574 GND.n1138 GND.n958 0.152939
R14575 GND.n959 GND.n958 0.152939
R14576 GND.n960 GND.n959 0.152939
R14577 GND.n961 GND.n960 0.152939
R14578 GND.n962 GND.n961 0.152939
R14579 GND.n963 GND.n962 0.152939
R14580 GND.n964 GND.n963 0.152939
R14581 GND.n965 GND.n964 0.152939
R14582 GND.n966 GND.n965 0.152939
R14583 GND.n967 GND.n966 0.152939
R14584 GND.n968 GND.n967 0.152939
R14585 GND.n969 GND.n968 0.152939
R14586 GND.n970 GND.n969 0.152939
R14587 GND.n971 GND.n970 0.152939
R14588 GND.n972 GND.n971 0.152939
R14589 GND.n973 GND.n972 0.152939
R14590 GND.n974 GND.n973 0.152939
R14591 GND.n975 GND.n974 0.152939
R14592 GND.n976 GND.n975 0.152939
R14593 GND.n977 GND.n976 0.152939
R14594 GND.n978 GND.n977 0.152939
R14595 GND.n979 GND.n978 0.152939
R14596 GND.n980 GND.n979 0.152939
R14597 GND.n981 GND.n980 0.152939
R14598 GND.n982 GND.n981 0.152939
R14599 GND.n983 GND.n982 0.152939
R14600 GND.n984 GND.n983 0.152939
R14601 GND.n985 GND.n984 0.152939
R14602 GND.n986 GND.n985 0.152939
R14603 GND.n987 GND.n986 0.152939
R14604 GND.n988 GND.n987 0.152939
R14605 GND.n989 GND.n988 0.152939
R14606 GND.n990 GND.n989 0.152939
R14607 GND.n991 GND.n990 0.152939
R14608 GND.n992 GND.n991 0.152939
R14609 GND.n993 GND.n992 0.152939
R14610 GND.n994 GND.n993 0.152939
R14611 GND.n995 GND.n994 0.152939
R14612 GND.n996 GND.n995 0.152939
R14613 GND.n997 GND.n996 0.152939
R14614 GND.n998 GND.n997 0.152939
R14615 GND.n999 GND.n998 0.152939
R14616 GND.n1000 GND.n999 0.152939
R14617 GND.n1001 GND.n1000 0.152939
R14618 GND.n1002 GND.n1001 0.152939
R14619 GND.n1003 GND.n1002 0.152939
R14620 GND.n1004 GND.n1003 0.152939
R14621 GND.n1005 GND.n1004 0.152939
R14622 GND.n1006 GND.n1005 0.152939
R14623 GND.n1007 GND.n1006 0.152939
R14624 GND.n1008 GND.n1007 0.152939
R14625 GND.n1009 GND.n1008 0.152939
R14626 GND.n1010 GND.n1009 0.152939
R14627 GND.n1011 GND.n1010 0.152939
R14628 GND.n1012 GND.n1011 0.152939
R14629 GND.n7635 GND.n247 0.152939
R14630 GND.n270 GND.n247 0.152939
R14631 GND.n271 GND.n270 0.152939
R14632 GND.n272 GND.n271 0.152939
R14633 GND.n290 GND.n272 0.152939
R14634 GND.n291 GND.n290 0.152939
R14635 GND.n292 GND.n291 0.152939
R14636 GND.n293 GND.n292 0.152939
R14637 GND.n4188 GND.n293 0.152939
R14638 GND.n4301 GND.n4083 0.152939
R14639 GND.n4301 GND.n4300 0.152939
R14640 GND.n4300 GND.n4299 0.152939
R14641 GND.n4299 GND.n4084 0.152939
R14642 GND.n4089 GND.n4084 0.152939
R14643 GND.n4090 GND.n4089 0.152939
R14644 GND.n4091 GND.n4090 0.152939
R14645 GND.n4096 GND.n4091 0.152939
R14646 GND.n4097 GND.n4096 0.152939
R14647 GND.n4098 GND.n4097 0.152939
R14648 GND.n4099 GND.n4098 0.152939
R14649 GND.n4104 GND.n4099 0.152939
R14650 GND.n4105 GND.n4104 0.152939
R14651 GND.n4106 GND.n4105 0.152939
R14652 GND.n4107 GND.n4106 0.152939
R14653 GND.n4112 GND.n4107 0.152939
R14654 GND.n4113 GND.n4112 0.152939
R14655 GND.n4114 GND.n4113 0.152939
R14656 GND.n4115 GND.n4114 0.152939
R14657 GND.n4120 GND.n4115 0.152939
R14658 GND.n4121 GND.n4120 0.152939
R14659 GND.n4122 GND.n4121 0.152939
R14660 GND.n4123 GND.n4122 0.152939
R14661 GND.n4128 GND.n4123 0.152939
R14662 GND.n4129 GND.n4128 0.152939
R14663 GND.n4130 GND.n4129 0.152939
R14664 GND.n4131 GND.n4130 0.152939
R14665 GND.n4136 GND.n4131 0.152939
R14666 GND.n4137 GND.n4136 0.152939
R14667 GND.n4138 GND.n4137 0.152939
R14668 GND.n4139 GND.n4138 0.152939
R14669 GND.n4144 GND.n4139 0.152939
R14670 GND.n4145 GND.n4144 0.152939
R14671 GND.n4146 GND.n4145 0.152939
R14672 GND.n4147 GND.n4146 0.152939
R14673 GND.n4152 GND.n4147 0.152939
R14674 GND.n4153 GND.n4152 0.152939
R14675 GND.n4154 GND.n4153 0.152939
R14676 GND.n4155 GND.n4154 0.152939
R14677 GND.n4160 GND.n4155 0.152939
R14678 GND.n4161 GND.n4160 0.152939
R14679 GND.n4162 GND.n4161 0.152939
R14680 GND.n4163 GND.n4162 0.152939
R14681 GND.n4168 GND.n4163 0.152939
R14682 GND.n4169 GND.n4168 0.152939
R14683 GND.n4170 GND.n4169 0.152939
R14684 GND.n4171 GND.n4170 0.152939
R14685 GND.n4176 GND.n4171 0.152939
R14686 GND.n4177 GND.n4176 0.152939
R14687 GND.n4178 GND.n4177 0.152939
R14688 GND.n4179 GND.n4178 0.152939
R14689 GND.n4184 GND.n4179 0.152939
R14690 GND.n4185 GND.n4184 0.152939
R14691 GND.n4186 GND.n4185 0.152939
R14692 GND.n4187 GND.n4186 0.152939
R14693 GND.n4189 GND.n4187 0.152939
R14694 GND.n4862 GND.n3524 0.152939
R14695 GND.n3530 GND.n3524 0.152939
R14696 GND.n3531 GND.n3530 0.152939
R14697 GND.n3532 GND.n3531 0.152939
R14698 GND.n3533 GND.n3532 0.152939
R14699 GND.n3538 GND.n3533 0.152939
R14700 GND.n3539 GND.n3538 0.152939
R14701 GND.n3540 GND.n3539 0.152939
R14702 GND.n3541 GND.n3540 0.152939
R14703 GND.n3546 GND.n3541 0.152939
R14704 GND.n3547 GND.n3546 0.152939
R14705 GND.n3548 GND.n3547 0.152939
R14706 GND.n3549 GND.n3548 0.152939
R14707 GND.n3554 GND.n3549 0.152939
R14708 GND.n3555 GND.n3554 0.152939
R14709 GND.n3556 GND.n3555 0.152939
R14710 GND.n3557 GND.n3556 0.152939
R14711 GND.n3562 GND.n3557 0.152939
R14712 GND.n3563 GND.n3562 0.152939
R14713 GND.n3564 GND.n3563 0.152939
R14714 GND.n3565 GND.n3564 0.152939
R14715 GND.n3570 GND.n3565 0.152939
R14716 GND.n3571 GND.n3570 0.152939
R14717 GND.n3572 GND.n3571 0.152939
R14718 GND.n3573 GND.n3572 0.152939
R14719 GND.n3578 GND.n3573 0.152939
R14720 GND.n3579 GND.n3578 0.152939
R14721 GND.n3580 GND.n3579 0.152939
R14722 GND.n3581 GND.n3580 0.152939
R14723 GND.n3586 GND.n3581 0.152939
R14724 GND.n3587 GND.n3586 0.152939
R14725 GND.n3588 GND.n3587 0.152939
R14726 GND.n3589 GND.n3588 0.152939
R14727 GND.n3594 GND.n3589 0.152939
R14728 GND.n3595 GND.n3594 0.152939
R14729 GND.n3596 GND.n3595 0.152939
R14730 GND.n3597 GND.n3596 0.152939
R14731 GND.n3602 GND.n3597 0.152939
R14732 GND.n3603 GND.n3602 0.152939
R14733 GND.n3604 GND.n3603 0.152939
R14734 GND.n3605 GND.n3604 0.152939
R14735 GND.n3610 GND.n3605 0.152939
R14736 GND.n3611 GND.n3610 0.152939
R14737 GND.n3612 GND.n3611 0.152939
R14738 GND.n3613 GND.n3612 0.152939
R14739 GND.n3618 GND.n3613 0.152939
R14740 GND.n3619 GND.n3618 0.152939
R14741 GND.n3620 GND.n3619 0.152939
R14742 GND.n3621 GND.n3620 0.152939
R14743 GND.n3626 GND.n3621 0.152939
R14744 GND.n3627 GND.n3626 0.152939
R14745 GND.n3628 GND.n3627 0.152939
R14746 GND.n3629 GND.n3628 0.152939
R14747 GND.n3634 GND.n3629 0.152939
R14748 GND.n3635 GND.n3634 0.152939
R14749 GND.n3636 GND.n3635 0.152939
R14750 GND.n3637 GND.n3636 0.152939
R14751 GND.n3642 GND.n3637 0.152939
R14752 GND.n3643 GND.n3642 0.152939
R14753 GND.n3644 GND.n3643 0.152939
R14754 GND.n3645 GND.n3644 0.152939
R14755 GND.n3650 GND.n3645 0.152939
R14756 GND.n3651 GND.n3650 0.152939
R14757 GND.n3652 GND.n3651 0.152939
R14758 GND.n3653 GND.n3652 0.152939
R14759 GND.n3658 GND.n3653 0.152939
R14760 GND.n3659 GND.n3658 0.152939
R14761 GND.n3660 GND.n3659 0.152939
R14762 GND.n3661 GND.n3660 0.152939
R14763 GND.n3666 GND.n3661 0.152939
R14764 GND.n3667 GND.n3666 0.152939
R14765 GND.n3668 GND.n3667 0.152939
R14766 GND.n3669 GND.n3668 0.152939
R14767 GND.n3674 GND.n3669 0.152939
R14768 GND.n3675 GND.n3674 0.152939
R14769 GND.n3676 GND.n3675 0.152939
R14770 GND.n3677 GND.n3676 0.152939
R14771 GND.n3682 GND.n3677 0.152939
R14772 GND.n3683 GND.n3682 0.152939
R14773 GND.n3684 GND.n3683 0.152939
R14774 GND.n3685 GND.n3684 0.152939
R14775 GND.n3690 GND.n3685 0.152939
R14776 GND.n3691 GND.n3690 0.152939
R14777 GND.n3692 GND.n3691 0.152939
R14778 GND.n3693 GND.n3692 0.152939
R14779 GND.n3698 GND.n3693 0.152939
R14780 GND.n3699 GND.n3698 0.152939
R14781 GND.n3700 GND.n3699 0.152939
R14782 GND.n3701 GND.n3700 0.152939
R14783 GND.n3706 GND.n3701 0.152939
R14784 GND.n3707 GND.n3706 0.152939
R14785 GND.n3708 GND.n3707 0.152939
R14786 GND.n3709 GND.n3708 0.152939
R14787 GND.n3714 GND.n3709 0.152939
R14788 GND.n3715 GND.n3714 0.152939
R14789 GND.n3716 GND.n3715 0.152939
R14790 GND.n3717 GND.n3716 0.152939
R14791 GND.n3722 GND.n3717 0.152939
R14792 GND.n3723 GND.n3722 0.152939
R14793 GND.n3724 GND.n3723 0.152939
R14794 GND.n3725 GND.n3724 0.152939
R14795 GND.n3730 GND.n3725 0.152939
R14796 GND.n3731 GND.n3730 0.152939
R14797 GND.n3732 GND.n3731 0.152939
R14798 GND.n3733 GND.n3732 0.152939
R14799 GND.n3738 GND.n3733 0.152939
R14800 GND.n3739 GND.n3738 0.152939
R14801 GND.n3740 GND.n3739 0.152939
R14802 GND.n3741 GND.n3740 0.152939
R14803 GND.n3746 GND.n3741 0.152939
R14804 GND.n3747 GND.n3746 0.152939
R14805 GND.n3748 GND.n3747 0.152939
R14806 GND.n3749 GND.n3748 0.152939
R14807 GND.n3754 GND.n3749 0.152939
R14808 GND.n3755 GND.n3754 0.152939
R14809 GND.n3756 GND.n3755 0.152939
R14810 GND.n3757 GND.n3756 0.152939
R14811 GND.n3762 GND.n3757 0.152939
R14812 GND.n3763 GND.n3762 0.152939
R14813 GND.n3764 GND.n3763 0.152939
R14814 GND.n3765 GND.n3764 0.152939
R14815 GND.n3770 GND.n3765 0.152939
R14816 GND.n3771 GND.n3770 0.152939
R14817 GND.n3772 GND.n3771 0.152939
R14818 GND.n3773 GND.n3772 0.152939
R14819 GND.n3778 GND.n3773 0.152939
R14820 GND.n3779 GND.n3778 0.152939
R14821 GND.n3780 GND.n3779 0.152939
R14822 GND.n3781 GND.n3780 0.152939
R14823 GND.n3786 GND.n3781 0.152939
R14824 GND.n3787 GND.n3786 0.152939
R14825 GND.n3788 GND.n3787 0.152939
R14826 GND.n3789 GND.n3788 0.152939
R14827 GND.n3794 GND.n3789 0.152939
R14828 GND.n3795 GND.n3794 0.152939
R14829 GND.n3796 GND.n3795 0.152939
R14830 GND.n3797 GND.n3796 0.152939
R14831 GND.n3802 GND.n3797 0.152939
R14832 GND.n3803 GND.n3802 0.152939
R14833 GND.n3804 GND.n3803 0.152939
R14834 GND.n3805 GND.n3804 0.152939
R14835 GND.n3810 GND.n3805 0.152939
R14836 GND.n3811 GND.n3810 0.152939
R14837 GND.n3812 GND.n3811 0.152939
R14838 GND.n3813 GND.n3812 0.152939
R14839 GND.n3818 GND.n3813 0.152939
R14840 GND.n3819 GND.n3818 0.152939
R14841 GND.n3820 GND.n3819 0.152939
R14842 GND.n3821 GND.n3820 0.152939
R14843 GND.n3826 GND.n3821 0.152939
R14844 GND.n3827 GND.n3826 0.152939
R14845 GND.n3828 GND.n3827 0.152939
R14846 GND.n3829 GND.n3828 0.152939
R14847 GND.n3834 GND.n3829 0.152939
R14848 GND.n3835 GND.n3834 0.152939
R14849 GND.n3836 GND.n3835 0.152939
R14850 GND.n3837 GND.n3836 0.152939
R14851 GND.n3842 GND.n3837 0.152939
R14852 GND.n3843 GND.n3842 0.152939
R14853 GND.n3844 GND.n3843 0.152939
R14854 GND.n3845 GND.n3844 0.152939
R14855 GND.n3850 GND.n3845 0.152939
R14856 GND.n3851 GND.n3850 0.152939
R14857 GND.n3852 GND.n3851 0.152939
R14858 GND.n3853 GND.n3852 0.152939
R14859 GND.n3858 GND.n3853 0.152939
R14860 GND.n3859 GND.n3858 0.152939
R14861 GND.n3860 GND.n3859 0.152939
R14862 GND.n3861 GND.n3860 0.152939
R14863 GND.n3866 GND.n3861 0.152939
R14864 GND.n3867 GND.n3866 0.152939
R14865 GND.n3868 GND.n3867 0.152939
R14866 GND.n3869 GND.n3868 0.152939
R14867 GND.n3874 GND.n3869 0.152939
R14868 GND.n3875 GND.n3874 0.152939
R14869 GND.n3876 GND.n3875 0.152939
R14870 GND.n3877 GND.n3876 0.152939
R14871 GND.n3882 GND.n3877 0.152939
R14872 GND.n3883 GND.n3882 0.152939
R14873 GND.n3884 GND.n3883 0.152939
R14874 GND.n3885 GND.n3884 0.152939
R14875 GND.n3890 GND.n3885 0.152939
R14876 GND.n3891 GND.n3890 0.152939
R14877 GND.n3892 GND.n3891 0.152939
R14878 GND.n3893 GND.n3892 0.152939
R14879 GND.n3898 GND.n3893 0.152939
R14880 GND.n3899 GND.n3898 0.152939
R14881 GND.n3900 GND.n3899 0.152939
R14882 GND.n3901 GND.n3900 0.152939
R14883 GND.n3906 GND.n3901 0.152939
R14884 GND.n3907 GND.n3906 0.152939
R14885 GND.n3908 GND.n3907 0.152939
R14886 GND.n3909 GND.n3908 0.152939
R14887 GND.n3914 GND.n3909 0.152939
R14888 GND.n3915 GND.n3914 0.152939
R14889 GND.n3916 GND.n3915 0.152939
R14890 GND.n3917 GND.n3916 0.152939
R14891 GND.n3922 GND.n3917 0.152939
R14892 GND.n3923 GND.n3922 0.152939
R14893 GND.n3924 GND.n3923 0.152939
R14894 GND.n3925 GND.n3924 0.152939
R14895 GND.n3930 GND.n3925 0.152939
R14896 GND.n3931 GND.n3930 0.152939
R14897 GND.n3932 GND.n3931 0.152939
R14898 GND.n3933 GND.n3932 0.152939
R14899 GND.n3938 GND.n3933 0.152939
R14900 GND.n3939 GND.n3938 0.152939
R14901 GND.n3940 GND.n3939 0.152939
R14902 GND.n3941 GND.n3940 0.152939
R14903 GND.n3946 GND.n3941 0.152939
R14904 GND.n3947 GND.n3946 0.152939
R14905 GND.n3948 GND.n3947 0.152939
R14906 GND.n3949 GND.n3948 0.152939
R14907 GND.n3954 GND.n3949 0.152939
R14908 GND.n3955 GND.n3954 0.152939
R14909 GND.n3956 GND.n3955 0.152939
R14910 GND.n3957 GND.n3956 0.152939
R14911 GND.n3962 GND.n3957 0.152939
R14912 GND.n3963 GND.n3962 0.152939
R14913 GND.n3964 GND.n3963 0.152939
R14914 GND.n3965 GND.n3964 0.152939
R14915 GND.n3970 GND.n3965 0.152939
R14916 GND.n3971 GND.n3970 0.152939
R14917 GND.n3972 GND.n3971 0.152939
R14918 GND.n3973 GND.n3972 0.152939
R14919 GND.n3978 GND.n3973 0.152939
R14920 GND.n3979 GND.n3978 0.152939
R14921 GND.n3980 GND.n3979 0.152939
R14922 GND.n3981 GND.n3980 0.152939
R14923 GND.n3986 GND.n3981 0.152939
R14924 GND.n3987 GND.n3986 0.152939
R14925 GND.n3988 GND.n3987 0.152939
R14926 GND.n3989 GND.n3988 0.152939
R14927 GND.n3994 GND.n3989 0.152939
R14928 GND.n3995 GND.n3994 0.152939
R14929 GND.n3996 GND.n3995 0.152939
R14930 GND.n3997 GND.n3996 0.152939
R14931 GND.n4002 GND.n3997 0.152939
R14932 GND.n4003 GND.n4002 0.152939
R14933 GND.n4004 GND.n4003 0.152939
R14934 GND.n4005 GND.n4004 0.152939
R14935 GND.n4010 GND.n4005 0.152939
R14936 GND.n4011 GND.n4010 0.152939
R14937 GND.n4012 GND.n4011 0.152939
R14938 GND.n4013 GND.n4012 0.152939
R14939 GND.n4018 GND.n4013 0.152939
R14940 GND.n4019 GND.n4018 0.152939
R14941 GND.n4020 GND.n4019 0.152939
R14942 GND.n4021 GND.n4020 0.152939
R14943 GND.n4026 GND.n4021 0.152939
R14944 GND.n4027 GND.n4026 0.152939
R14945 GND.n4028 GND.n4027 0.152939
R14946 GND.n4029 GND.n4028 0.152939
R14947 GND.n4034 GND.n4029 0.152939
R14948 GND.n4035 GND.n4034 0.152939
R14949 GND.n4036 GND.n4035 0.152939
R14950 GND.n4037 GND.n4036 0.152939
R14951 GND.n4042 GND.n4037 0.152939
R14952 GND.n4043 GND.n4042 0.152939
R14953 GND.n4044 GND.n4043 0.152939
R14954 GND.n4045 GND.n4044 0.152939
R14955 GND.n4050 GND.n4045 0.152939
R14956 GND.n4051 GND.n4050 0.152939
R14957 GND.n4052 GND.n4051 0.152939
R14958 GND.n4053 GND.n4052 0.152939
R14959 GND.n4058 GND.n4053 0.152939
R14960 GND.n4059 GND.n4058 0.152939
R14961 GND.n4060 GND.n4059 0.152939
R14962 GND.n4061 GND.n4060 0.152939
R14963 GND.n4066 GND.n4061 0.152939
R14964 GND.n4067 GND.n4066 0.152939
R14965 GND.n4068 GND.n4067 0.152939
R14966 GND.n4069 GND.n4068 0.152939
R14967 GND.n4074 GND.n4069 0.152939
R14968 GND.n4075 GND.n4074 0.152939
R14969 GND.n4076 GND.n4075 0.152939
R14970 GND.n4077 GND.n4076 0.152939
R14971 GND.n4864 GND.n4863 0.152939
R14972 GND.n4865 GND.n4864 0.152939
R14973 GND.n4866 GND.n4865 0.152939
R14974 GND.n4867 GND.n4866 0.152939
R14975 GND.n4868 GND.n4867 0.152939
R14976 GND.n4869 GND.n4868 0.152939
R14977 GND.n4870 GND.n4869 0.152939
R14978 GND.n4871 GND.n4870 0.152939
R14979 GND.n4872 GND.n4871 0.152939
R14980 GND.n4873 GND.n4872 0.152939
R14981 GND.n4874 GND.n4873 0.152939
R14982 GND.n4875 GND.n4874 0.152939
R14983 GND.n4876 GND.n4875 0.152939
R14984 GND.n4877 GND.n4876 0.152939
R14985 GND.n4878 GND.n4877 0.152939
R14986 GND.n4879 GND.n4878 0.152939
R14987 GND.n4880 GND.n4879 0.152939
R14988 GND.n4881 GND.n4880 0.152939
R14989 GND.n4882 GND.n4881 0.152939
R14990 GND.n4883 GND.n4882 0.152939
R14991 GND.n4884 GND.n4883 0.152939
R14992 GND.n4885 GND.n4884 0.152939
R14993 GND.n4886 GND.n4885 0.152939
R14994 GND.n4887 GND.n4886 0.152939
R14995 GND.n4888 GND.n4887 0.152939
R14996 GND.n4889 GND.n4888 0.152939
R14997 GND.n4890 GND.n4889 0.152939
R14998 GND.n4891 GND.n4890 0.152939
R14999 GND.n4892 GND.n4891 0.152939
R15000 GND.n4893 GND.n4892 0.152939
R15001 GND.n4894 GND.n4893 0.152939
R15002 GND.n4895 GND.n4894 0.152939
R15003 GND.n4896 GND.n4895 0.152939
R15004 GND.n4897 GND.n4896 0.152939
R15005 GND.n4898 GND.n4897 0.152939
R15006 GND.n4899 GND.n4898 0.152939
R15007 GND.n4900 GND.n4899 0.152939
R15008 GND.n4901 GND.n4900 0.152939
R15009 GND.n4902 GND.n4901 0.152939
R15010 GND.n4903 GND.n4902 0.152939
R15011 GND.n4904 GND.n4903 0.152939
R15012 GND.n4905 GND.n4904 0.152939
R15013 GND.n4906 GND.n4905 0.152939
R15014 GND.n4907 GND.n4906 0.152939
R15015 GND.n4908 GND.n4907 0.152939
R15016 GND.n4909 GND.n4908 0.152939
R15017 GND.n4910 GND.n4909 0.152939
R15018 GND.n4911 GND.n4910 0.152939
R15019 GND.n4912 GND.n4911 0.152939
R15020 GND.n4913 GND.n4912 0.152939
R15021 GND.n4914 GND.n4913 0.152939
R15022 GND.n4915 GND.n4914 0.152939
R15023 GND.n4917 GND.n4915 0.152939
R15024 GND.n4917 GND.n4916 0.152939
R15025 GND.n4916 GND.n2787 0.152939
R15026 GND.n5030 GND.n2787 0.152939
R15027 GND.n5031 GND.n2768 0.152939
R15028 GND.n5053 GND.n2768 0.152939
R15029 GND.n5054 GND.n5053 0.152939
R15030 GND.n5055 GND.n5054 0.152939
R15031 GND.n5055 GND.n2536 0.152939
R15032 GND.n5213 GND.n2536 0.152939
R15033 GND.n5214 GND.n5213 0.152939
R15034 GND.n5215 GND.n5214 0.152939
R15035 GND.n5215 GND.n2512 0.152939
R15036 GND.n3181 GND.n3054 0.152939
R15037 GND.n3057 GND.n3054 0.152939
R15038 GND.n3058 GND.n3057 0.152939
R15039 GND.n3059 GND.n3058 0.152939
R15040 GND.n3062 GND.n3059 0.152939
R15041 GND.n3063 GND.n3062 0.152939
R15042 GND.n3064 GND.n3063 0.152939
R15043 GND.n3065 GND.n3064 0.152939
R15044 GND.n3070 GND.n3065 0.152939
R15045 GND.n3071 GND.n3070 0.152939
R15046 GND.n3072 GND.n3071 0.152939
R15047 GND.n3073 GND.n3072 0.152939
R15048 GND.n3076 GND.n3073 0.152939
R15049 GND.n3077 GND.n3076 0.152939
R15050 GND.n3078 GND.n3077 0.152939
R15051 GND.n3079 GND.n3078 0.152939
R15052 GND.n3082 GND.n3079 0.152939
R15053 GND.n3083 GND.n3082 0.152939
R15054 GND.n3142 GND.n3083 0.152939
R15055 GND.n3142 GND.n3141 0.152939
R15056 GND.n3141 GND.n3140 0.152939
R15057 GND.n3182 GND.n3036 0.152939
R15058 GND.n3204 GND.n3036 0.152939
R15059 GND.n3205 GND.n3204 0.152939
R15060 GND.n3206 GND.n3205 0.152939
R15061 GND.n3207 GND.n3206 0.152939
R15062 GND.n3207 GND.n3008 0.152939
R15063 GND.n3336 GND.n3008 0.152939
R15064 GND.n3337 GND.n3336 0.152939
R15065 GND.n3338 GND.n3337 0.152939
R15066 GND.n3338 GND.n2987 0.152939
R15067 GND.n3353 GND.n2987 0.152939
R15068 GND.n3354 GND.n3353 0.152939
R15069 GND.n3355 GND.n3354 0.152939
R15070 GND.n3355 GND.n2966 0.152939
R15071 GND.n3370 GND.n2966 0.152939
R15072 GND.n3371 GND.n3370 0.152939
R15073 GND.n3372 GND.n3371 0.152939
R15074 GND.n3372 GND.n2944 0.152939
R15075 GND.n3387 GND.n2944 0.152939
R15076 GND.n3388 GND.n3387 0.152939
R15077 GND.n3389 GND.n3388 0.152939
R15078 GND.n3389 GND.n2924 0.152939
R15079 GND.n3404 GND.n2924 0.152939
R15080 GND.n3405 GND.n3404 0.152939
R15081 GND.n3406 GND.n3405 0.152939
R15082 GND.n3406 GND.n2903 0.152939
R15083 GND.n3421 GND.n2903 0.152939
R15084 GND.n3422 GND.n3421 0.152939
R15085 GND.n3423 GND.n3422 0.152939
R15086 GND.n3423 GND.n2882 0.152939
R15087 GND.n3438 GND.n2882 0.152939
R15088 GND.n3439 GND.n3438 0.152939
R15089 GND.n3440 GND.n3439 0.152939
R15090 GND.n3440 GND.n2861 0.152939
R15091 GND.n3455 GND.n2861 0.152939
R15092 GND.n3456 GND.n3455 0.152939
R15093 GND.n3457 GND.n3456 0.152939
R15094 GND.n3457 GND.n2840 0.152939
R15095 GND.n3472 GND.n2840 0.152939
R15096 GND.n3473 GND.n3472 0.152939
R15097 GND.n3474 GND.n3473 0.152939
R15098 GND.n3474 GND.n2821 0.152939
R15099 GND.n3495 GND.n2821 0.152939
R15100 GND.n3496 GND.n3495 0.152939
R15101 GND.n3497 GND.n3496 0.152939
R15102 GND.n3498 GND.n3497 0.152939
R15103 GND.n3499 GND.n3498 0.152939
R15104 GND.n3500 GND.n3499 0.152939
R15105 GND.n3501 GND.n3500 0.152939
R15106 GND.n3502 GND.n3501 0.152939
R15107 GND.n3503 GND.n3502 0.152939
R15108 GND.n3504 GND.n3503 0.152939
R15109 GND.n3505 GND.n3504 0.152939
R15110 GND.n3505 GND.n2524 0.152939
R15111 GND.n5223 GND.n2524 0.152939
R15112 GND.n5088 GND.n5087 0.152939
R15113 GND.n5089 GND.n5088 0.152939
R15114 GND.n5090 GND.n5089 0.152939
R15115 GND.n5091 GND.n5090 0.152939
R15116 GND.n5092 GND.n5091 0.152939
R15117 GND.n5093 GND.n5092 0.152939
R15118 GND.n5094 GND.n5093 0.152939
R15119 GND.n5095 GND.n5094 0.152939
R15120 GND.n5096 GND.n5095 0.152939
R15121 GND.n5097 GND.n5096 0.152939
R15122 GND.n5098 GND.n5097 0.152939
R15123 GND.n5099 GND.n5098 0.152939
R15124 GND.n5100 GND.n5099 0.152939
R15125 GND.n5101 GND.n5100 0.152939
R15126 GND.n5102 GND.n5101 0.152939
R15127 GND.n5103 GND.n5102 0.152939
R15128 GND.n5104 GND.n5103 0.152939
R15129 GND.n5105 GND.n5104 0.152939
R15130 GND.n5106 GND.n5105 0.152939
R15131 GND.n5107 GND.n5106 0.152939
R15132 GND.n5108 GND.n5107 0.152939
R15133 GND.n5109 GND.n5108 0.152939
R15134 GND.n5110 GND.n5109 0.152939
R15135 GND.n5111 GND.n5110 0.152939
R15136 GND.n5112 GND.n5111 0.152939
R15137 GND.n5113 GND.n5112 0.152939
R15138 GND.n5114 GND.n5113 0.152939
R15139 GND.n5115 GND.n5114 0.152939
R15140 GND.n5116 GND.n5115 0.152939
R15141 GND.n5117 GND.n5116 0.152939
R15142 GND.n5118 GND.n5117 0.152939
R15143 GND.n5119 GND.n5118 0.152939
R15144 GND.n5120 GND.n5119 0.152939
R15145 GND.n5121 GND.n5120 0.152939
R15146 GND.n5122 GND.n5121 0.152939
R15147 GND.n5122 GND.n2342 0.152939
R15148 GND.n5399 GND.n2342 0.152939
R15149 GND.n5400 GND.n5399 0.152939
R15150 GND.n5401 GND.n5400 0.152939
R15151 GND.n5402 GND.n5401 0.152939
R15152 GND.n5403 GND.n5402 0.152939
R15153 GND.n5404 GND.n5403 0.152939
R15154 GND.n5405 GND.n5404 0.152939
R15155 GND.n5406 GND.n5405 0.152939
R15156 GND.n5407 GND.n5406 0.152939
R15157 GND.n5408 GND.n5407 0.152939
R15158 GND.n5409 GND.n5408 0.152939
R15159 GND.n5410 GND.n5409 0.152939
R15160 GND.n5411 GND.n5410 0.152939
R15161 GND.n5412 GND.n5411 0.152939
R15162 GND.n5413 GND.n5412 0.152939
R15163 GND.n5414 GND.n5413 0.152939
R15164 GND.n5415 GND.n5414 0.152939
R15165 GND.n5416 GND.n5415 0.152939
R15166 GND.n5417 GND.n5416 0.152939
R15167 GND.n5418 GND.n5417 0.152939
R15168 GND.n5419 GND.n5418 0.152939
R15169 GND.n5420 GND.n5419 0.152939
R15170 GND.n5421 GND.n5420 0.152939
R15171 GND.n5421 GND.n1724 0.152939
R15172 GND.n5823 GND.n5822 0.152939
R15173 GND.n5825 GND.n5823 0.152939
R15174 GND.n5825 GND.n5824 0.152939
R15175 GND.n5824 GND.n1652 0.152939
R15176 GND.n5856 GND.n1652 0.152939
R15177 GND.n5857 GND.n5856 0.152939
R15178 GND.n5858 GND.n5857 0.152939
R15179 GND.n5858 GND.n1624 0.152939
R15180 GND.n5900 GND.n1624 0.152939
R15181 GND.n5901 GND.n5900 0.152939
R15182 GND.n5902 GND.n5901 0.152939
R15183 GND.n5902 GND.n1582 0.152939
R15184 GND.n5941 GND.n1582 0.152939
R15185 GND.n5942 GND.n5941 0.152939
R15186 GND.n5944 GND.n5942 0.152939
R15187 GND.n5944 GND.n5943 0.152939
R15188 GND.n5943 GND.n1550 0.152939
R15189 GND.n6009 GND.n1550 0.152939
R15190 GND.n6010 GND.n6009 0.152939
R15191 GND.n6011 GND.n6010 0.152939
R15192 GND.n6011 GND.n1531 0.152939
R15193 GND.n6061 GND.n1531 0.152939
R15194 GND.n6062 GND.n6061 0.152939
R15195 GND.n6064 GND.n6062 0.152939
R15196 GND.n6064 GND.n6063 0.152939
R15197 GND.n6063 GND.n1499 0.152939
R15198 GND.n6100 GND.n1499 0.152939
R15199 GND.n6101 GND.n6100 0.152939
R15200 GND.n6102 GND.n6101 0.152939
R15201 GND.n6102 GND.n1472 0.152939
R15202 GND.n6154 GND.n1472 0.152939
R15203 GND.n6155 GND.n6154 0.152939
R15204 GND.n6166 GND.n6155 0.152939
R15205 GND.n6166 GND.n6165 0.152939
R15206 GND.n6165 GND.n6164 0.152939
R15207 GND.n6164 GND.n6156 0.152939
R15208 GND.n6160 GND.n6156 0.152939
R15209 GND.n6160 GND.n1424 0.152939
R15210 GND.n6263 GND.n1424 0.152939
R15211 GND.n6264 GND.n6263 0.152939
R15212 GND.n6265 GND.n6264 0.152939
R15213 GND.n6265 GND.n1338 0.152939
R15214 GND.n6313 GND.n1338 0.152939
R15215 GND.n6313 GND.n6312 0.152939
R15216 GND.n6311 GND.n1339 0.152939
R15217 GND.n6307 GND.n1339 0.152939
R15218 GND.n6307 GND.n6306 0.152939
R15219 GND.n6304 GND.n1379 0.152939
R15220 GND.n6300 GND.n1379 0.152939
R15221 GND.n6300 GND.n6299 0.152939
R15222 GND.n6299 GND.n6298 0.152939
R15223 GND.n6298 GND.n1387 0.152939
R15224 GND.n6294 GND.n1387 0.152939
R15225 GND.n6294 GND.n6293 0.152939
R15226 GND.n6293 GND.n6292 0.152939
R15227 GND.n6292 GND.n1395 0.152939
R15228 GND.n6288 GND.n1395 0.152939
R15229 GND.n6288 GND.n6287 0.152939
R15230 GND.n6287 GND.n6286 0.152939
R15231 GND.n6286 GND.n1403 0.152939
R15232 GND.n6281 GND.n1403 0.152939
R15233 GND.n6281 GND.n6280 0.152939
R15234 GND.n6280 GND.n6279 0.152939
R15235 GND.n5728 GND.n1672 0.152939
R15236 GND.n5831 GND.n1672 0.152939
R15237 GND.n5832 GND.n5831 0.152939
R15238 GND.n5835 GND.n5832 0.152939
R15239 GND.n5835 GND.n5834 0.152939
R15240 GND.n5834 GND.n5833 0.152939
R15241 GND.n5833 GND.n1645 0.152939
R15242 GND.n5865 GND.n1645 0.152939
R15243 GND.n5866 GND.n5865 0.152939
R15244 GND.n5875 GND.n5866 0.152939
R15245 GND.n5875 GND.n5874 0.152939
R15246 GND.n5874 GND.n5873 0.152939
R15247 GND.n5873 GND.n5867 0.152939
R15248 GND.n5869 GND.n5867 0.152939
R15249 GND.n5869 GND.n5868 0.152939
R15250 GND.n5868 GND.n1572 0.152939
R15251 GND.n5952 GND.n1572 0.152939
R15252 GND.n5953 GND.n5952 0.152939
R15253 GND.n5973 GND.n5953 0.152939
R15254 GND.n5973 GND.n5972 0.152939
R15255 GND.n5972 GND.n5971 0.152939
R15256 GND.n5971 GND.n5954 0.152939
R15257 GND.n5967 GND.n5954 0.152939
R15258 GND.n5967 GND.n5966 0.152939
R15259 GND.n5966 GND.n5965 0.152939
R15260 GND.n5965 GND.n5957 0.152939
R15261 GND.n5961 GND.n5957 0.152939
R15262 GND.n5961 GND.n5960 0.152939
R15263 GND.n5960 GND.n1493 0.152939
R15264 GND.n6109 GND.n1493 0.152939
R15265 GND.n6110 GND.n6109 0.152939
R15266 GND.n6129 GND.n6110 0.152939
R15267 GND.n6129 GND.n6128 0.152939
R15268 GND.n6128 GND.n6127 0.152939
R15269 GND.n6127 GND.n6111 0.152939
R15270 GND.n6123 GND.n6111 0.152939
R15271 GND.n6123 GND.n6122 0.152939
R15272 GND.n6122 GND.n6121 0.152939
R15273 GND.n6121 GND.n6116 0.152939
R15274 GND.n6116 GND.n1417 0.152939
R15275 GND.n6271 GND.n1417 0.152939
R15276 GND.n6272 GND.n6271 0.152939
R15277 GND.n6273 GND.n6272 0.152939
R15278 GND.n6273 GND.n1413 0.152939
R15279 GND.n5758 GND.n1681 0.152939
R15280 GND.n5758 GND.n5757 0.152939
R15281 GND.n5757 GND.n5756 0.152939
R15282 GND.n5753 GND.n5752 0.152939
R15283 GND.n5752 GND.n5751 0.152939
R15284 GND.n5751 GND.n5702 0.152939
R15285 GND.n5747 GND.n5702 0.152939
R15286 GND.n5747 GND.n5746 0.152939
R15287 GND.n5746 GND.n5745 0.152939
R15288 GND.n5745 GND.n5708 0.152939
R15289 GND.n5741 GND.n5708 0.152939
R15290 GND.n5741 GND.n5740 0.152939
R15291 GND.n5740 GND.n5739 0.152939
R15292 GND.n5739 GND.n5714 0.152939
R15293 GND.n5735 GND.n5714 0.152939
R15294 GND.n5735 GND.n5734 0.152939
R15295 GND.n5734 GND.n5721 0.152939
R15296 GND.n5730 GND.n5721 0.152939
R15297 GND.n5730 GND.n5729 0.152939
R15298 GND.n5569 GND.n5568 0.152939
R15299 GND.n5570 GND.n5569 0.152939
R15300 GND.n5570 GND.n2232 0.152939
R15301 GND.n5578 GND.n2232 0.152939
R15302 GND.n5579 GND.n5578 0.152939
R15303 GND.n5581 GND.n5579 0.152939
R15304 GND.n5581 GND.n5580 0.152939
R15305 GND.n5628 GND.n5627 0.152939
R15306 GND.n5627 GND.n5626 0.152939
R15307 GND.n5626 GND.n5590 0.152939
R15308 GND.n5622 GND.n5590 0.152939
R15309 GND.n5622 GND.n5621 0.152939
R15310 GND.n5621 GND.n5620 0.152939
R15311 GND.n5620 GND.n5598 0.152939
R15312 GND.n5616 GND.n5598 0.152939
R15313 GND.n5616 GND.n5615 0.152939
R15314 GND.n5615 GND.n5614 0.152939
R15315 GND.n5614 GND.n1731 0.152939
R15316 GND.n3137 GND.n3091 0.152939
R15317 GND.n3130 GND.n3091 0.152939
R15318 GND.n3130 GND.n3129 0.152939
R15319 GND.n3129 GND.n3128 0.152939
R15320 GND.n3128 GND.n3095 0.152939
R15321 GND.n3124 GND.n3095 0.152939
R15322 GND.n3124 GND.n3123 0.152939
R15323 GND.n3123 GND.n3122 0.152939
R15324 GND.n3122 GND.n3102 0.152939
R15325 GND.n3113 GND.n3102 0.152939
R15326 GND.n3112 GND.n3106 0.152939
R15327 GND.n3108 GND.n3106 0.152939
R15328 GND.n3108 GND.n3027 0.152939
R15329 GND.n3214 GND.n3027 0.152939
R15330 GND.n3215 GND.n3214 0.152939
R15331 GND.n3322 GND.n3215 0.152939
R15332 GND.n3322 GND.n3321 0.152939
R15333 GND.n3321 GND.n3320 0.152939
R15334 GND.n3320 GND.n3216 0.152939
R15335 GND.n3316 GND.n3216 0.152939
R15336 GND.n3316 GND.n3315 0.152939
R15337 GND.n3315 GND.n3314 0.152939
R15338 GND.n3314 GND.n3220 0.152939
R15339 GND.n3310 GND.n3220 0.152939
R15340 GND.n3310 GND.n3309 0.152939
R15341 GND.n3309 GND.n3308 0.152939
R15342 GND.n3308 GND.n3224 0.152939
R15343 GND.n3304 GND.n3224 0.152939
R15344 GND.n3304 GND.n3303 0.152939
R15345 GND.n3303 GND.n3302 0.152939
R15346 GND.n3302 GND.n3228 0.152939
R15347 GND.n3298 GND.n3228 0.152939
R15348 GND.n3298 GND.n3297 0.152939
R15349 GND.n3297 GND.n3296 0.152939
R15350 GND.n3296 GND.n3232 0.152939
R15351 GND.n3292 GND.n3232 0.152939
R15352 GND.n3292 GND.n3291 0.152939
R15353 GND.n3291 GND.n3290 0.152939
R15354 GND.n3290 GND.n3236 0.152939
R15355 GND.n3286 GND.n3236 0.152939
R15356 GND.n3286 GND.n3285 0.152939
R15357 GND.n3285 GND.n3284 0.152939
R15358 GND.n3284 GND.n3240 0.152939
R15359 GND.n3280 GND.n3240 0.152939
R15360 GND.n3280 GND.n3279 0.152939
R15361 GND.n3279 GND.n3278 0.152939
R15362 GND.n3278 GND.n3244 0.152939
R15363 GND.n3274 GND.n3244 0.152939
R15364 GND.n3274 GND.n3273 0.152939
R15365 GND.n3273 GND.n3272 0.152939
R15366 GND.n3272 GND.n3248 0.152939
R15367 GND.n3268 GND.n3248 0.152939
R15368 GND.n3268 GND.n3267 0.152939
R15369 GND.n3267 GND.n3266 0.152939
R15370 GND.n3266 GND.n3252 0.152939
R15371 GND.n3262 GND.n3252 0.152939
R15372 GND.n3262 GND.n3261 0.152939
R15373 GND.n3261 GND.n3260 0.152939
R15374 GND.n3260 GND.n3257 0.152939
R15375 GND.n3257 GND.n3256 0.152939
R15376 GND.n3256 GND.n2759 0.152939
R15377 GND.n5063 GND.n2759 0.152939
R15378 GND.n5064 GND.n5063 0.152939
R15379 GND.n5065 GND.n5064 0.152939
R15380 GND.n5065 GND.n2752 0.152939
R15381 GND.n5070 GND.n2752 0.152939
R15382 GND.n5071 GND.n5070 0.152939
R15383 GND.n5072 GND.n5071 0.152939
R15384 GND.n5072 GND.n2724 0.152939
R15385 GND.n5085 GND.n2724 0.152939
R15386 GND.n6305 GND.n6304 0.0828171
R15387 GND.n5753 GND.n5697 0.0828171
R15388 GND.n5224 GND.n2518 0.0767195
R15389 GND.n5226 GND.n5225 0.0767195
R15390 GND.n7636 GND.n242 0.0767195
R15391 GND.n1014 GND.n246 0.0767195
R15392 GND.n1012 GND.n246 0.0767195
R15393 GND.n7636 GND.n7635 0.0767195
R15394 GND.n5225 GND.n2512 0.0767195
R15395 GND.n5224 GND.n5223 0.0767195
R15396 GND.n6306 GND.n6305 0.070622
R15397 GND.n5756 GND.n5697 0.070622
R15398 GND.n7645 GND.n227 0.0695946
R15399 GND.n7645 GND.n7644 0.0695946
R15400 GND.n5087 GND.n5086 0.0695946
R15401 GND.n5086 GND.n5085 0.0695946
R15402 GND.n1378 GND.n929 0.063
R15403 GND.n5696 GND.n5695 0.063
R15404 GND.n6737 GND.n929 0.0429592
R15405 GND.n7423 GND.n7422 0.0429592
R15406 GND.n3138 GND.n3090 0.0429592
R15407 GND.n5695 GND.n5694 0.0429592
R15408 GND.n6738 GND.n6737 0.0344674
R15409 GND.n6738 GND.n925 0.0344674
R15410 GND.n926 GND.n925 0.0344674
R15411 GND.n6744 GND.n926 0.0344674
R15412 GND.n6745 GND.n6744 0.0344674
R15413 GND.n6745 GND.n899 0.0344674
R15414 GND.n899 GND.n897 0.0344674
R15415 GND.n6857 GND.n897 0.0344674
R15416 GND.n6858 GND.n6857 0.0344674
R15417 GND.n6858 GND.n880 0.0344674
R15418 GND.n880 GND.n878 0.0344674
R15419 GND.n6877 GND.n878 0.0344674
R15420 GND.n6878 GND.n6877 0.0344674
R15421 GND.n6878 GND.n860 0.0344674
R15422 GND.n860 GND.n858 0.0344674
R15423 GND.n6897 GND.n858 0.0344674
R15424 GND.n6898 GND.n6897 0.0344674
R15425 GND.n6898 GND.n840 0.0344674
R15426 GND.n840 GND.n838 0.0344674
R15427 GND.n6917 GND.n838 0.0344674
R15428 GND.n6918 GND.n6917 0.0344674
R15429 GND.n6918 GND.n820 0.0344674
R15430 GND.n820 GND.n818 0.0344674
R15431 GND.n6937 GND.n818 0.0344674
R15432 GND.n6938 GND.n6937 0.0344674
R15433 GND.n6938 GND.n800 0.0344674
R15434 GND.n800 GND.n798 0.0344674
R15435 GND.n6957 GND.n798 0.0344674
R15436 GND.n6958 GND.n6957 0.0344674
R15437 GND.n6958 GND.n780 0.0344674
R15438 GND.n780 GND.n778 0.0344674
R15439 GND.n6977 GND.n778 0.0344674
R15440 GND.n6978 GND.n6977 0.0344674
R15441 GND.n6978 GND.n760 0.0344674
R15442 GND.n760 GND.n758 0.0344674
R15443 GND.n6997 GND.n758 0.0344674
R15444 GND.n6998 GND.n6997 0.0344674
R15445 GND.n6998 GND.n740 0.0344674
R15446 GND.n740 GND.n737 0.0344674
R15447 GND.n738 GND.n737 0.0344674
R15448 GND.n7019 GND.n738 0.0344674
R15449 GND.n7020 GND.n7019 0.0344674
R15450 GND.n7020 GND.n711 0.0344674
R15451 GND.n711 GND.n709 0.0344674
R15452 GND.n7065 GND.n709 0.0344674
R15453 GND.n7066 GND.n7065 0.0344674
R15454 GND.n7066 GND.n692 0.0344674
R15455 GND.n692 GND.n689 0.0344674
R15456 GND.n690 GND.n689 0.0344674
R15457 GND.n7094 GND.n690 0.0344674
R15458 GND.n7094 GND.n7093 0.0344674
R15459 GND.n7093 GND.n662 0.0344674
R15460 GND.n663 GND.n662 0.0344674
R15461 GND.n664 GND.n663 0.0344674
R15462 GND.n665 GND.n664 0.0344674
R15463 GND.n665 GND.n643 0.0344674
R15464 GND.n643 GND.n641 0.0344674
R15465 GND.n7156 GND.n641 0.0344674
R15466 GND.n7156 GND.n7155 0.0344674
R15467 GND.n7155 GND.n628 0.0344674
R15468 GND.n628 GND.n626 0.0344674
R15469 GND.n7175 GND.n626 0.0344674
R15470 GND.n7175 GND.n624 0.0344674
R15471 GND.n7202 GND.n624 0.0344674
R15472 GND.n7202 GND.n7201 0.0344674
R15473 GND.n7201 GND.n259 0.0344674
R15474 GND.n260 GND.n259 0.0344674
R15475 GND.n261 GND.n260 0.0344674
R15476 GND.n7181 GND.n261 0.0344674
R15477 GND.n7181 GND.n280 0.0344674
R15478 GND.n281 GND.n280 0.0344674
R15479 GND.n282 GND.n281 0.0344674
R15480 GND.n7182 GND.n282 0.0344674
R15481 GND.n7182 GND.n301 0.0344674
R15482 GND.n302 GND.n301 0.0344674
R15483 GND.n303 GND.n302 0.0344674
R15484 GND.n323 GND.n303 0.0344674
R15485 GND.n324 GND.n323 0.0344674
R15486 GND.n325 GND.n324 0.0344674
R15487 GND.n326 GND.n325 0.0344674
R15488 GND.n7351 GND.n326 0.0344674
R15489 GND.n7351 GND.n343 0.0344674
R15490 GND.n344 GND.n343 0.0344674
R15491 GND.n345 GND.n344 0.0344674
R15492 GND.n7358 GND.n345 0.0344674
R15493 GND.n7358 GND.n362 0.0344674
R15494 GND.n363 GND.n362 0.0344674
R15495 GND.n364 GND.n363 0.0344674
R15496 GND.n7365 GND.n364 0.0344674
R15497 GND.n7365 GND.n381 0.0344674
R15498 GND.n382 GND.n381 0.0344674
R15499 GND.n383 GND.n382 0.0344674
R15500 GND.n7372 GND.n383 0.0344674
R15501 GND.n7372 GND.n400 0.0344674
R15502 GND.n401 GND.n400 0.0344674
R15503 GND.n402 GND.n401 0.0344674
R15504 GND.n7379 GND.n402 0.0344674
R15505 GND.n7379 GND.n419 0.0344674
R15506 GND.n420 GND.n419 0.0344674
R15507 GND.n421 GND.n420 0.0344674
R15508 GND.n7386 GND.n421 0.0344674
R15509 GND.n7386 GND.n438 0.0344674
R15510 GND.n439 GND.n438 0.0344674
R15511 GND.n440 GND.n439 0.0344674
R15512 GND.n7393 GND.n440 0.0344674
R15513 GND.n7393 GND.n458 0.0344674
R15514 GND.n459 GND.n458 0.0344674
R15515 GND.n460 GND.n459 0.0344674
R15516 GND.n7400 GND.n460 0.0344674
R15517 GND.n7400 GND.n477 0.0344674
R15518 GND.n478 GND.n477 0.0344674
R15519 GND.n479 GND.n478 0.0344674
R15520 GND.n7407 GND.n479 0.0344674
R15521 GND.n7407 GND.n495 0.0344674
R15522 GND.n496 GND.n495 0.0344674
R15523 GND.n497 GND.n496 0.0344674
R15524 GND.n7414 GND.n497 0.0344674
R15525 GND.n7414 GND.n515 0.0344674
R15526 GND.n516 GND.n515 0.0344674
R15527 GND.n517 GND.n516 0.0344674
R15528 GND.n7422 GND.n517 0.0344674
R15529 GND.n3090 GND.n3046 0.0344674
R15530 GND.n3198 GND.n3046 0.0344674
R15531 GND.n3198 GND.n3047 0.0344674
R15532 GND.n3194 GND.n3047 0.0344674
R15533 GND.n3194 GND.n3193 0.0344674
R15534 GND.n3193 GND.n3017 0.0344674
R15535 GND.n3330 GND.n3017 0.0344674
R15536 GND.n3330 GND.n3020 0.0344674
R15537 GND.n3020 GND.n3019 0.0344674
R15538 GND.n3019 GND.n2997 0.0344674
R15539 GND.n3347 GND.n2997 0.0344674
R15540 GND.n3347 GND.n3000 0.0344674
R15541 GND.n3000 GND.n2999 0.0344674
R15542 GND.n2999 GND.n2976 0.0344674
R15543 GND.n3364 GND.n2976 0.0344674
R15544 GND.n3364 GND.n2979 0.0344674
R15545 GND.n2979 GND.n2978 0.0344674
R15546 GND.n2978 GND.n2955 0.0344674
R15547 GND.n3381 GND.n2955 0.0344674
R15548 GND.n3381 GND.n2958 0.0344674
R15549 GND.n2958 GND.n2957 0.0344674
R15550 GND.n2957 GND.n2934 0.0344674
R15551 GND.n3398 GND.n2934 0.0344674
R15552 GND.n3398 GND.n2937 0.0344674
R15553 GND.n2937 GND.n2936 0.0344674
R15554 GND.n2936 GND.n2913 0.0344674
R15555 GND.n3415 GND.n2913 0.0344674
R15556 GND.n3415 GND.n2916 0.0344674
R15557 GND.n2916 GND.n2915 0.0344674
R15558 GND.n2915 GND.n2892 0.0344674
R15559 GND.n3432 GND.n2892 0.0344674
R15560 GND.n3432 GND.n2895 0.0344674
R15561 GND.n2895 GND.n2894 0.0344674
R15562 GND.n2894 GND.n2871 0.0344674
R15563 GND.n3449 GND.n2871 0.0344674
R15564 GND.n3449 GND.n2874 0.0344674
R15565 GND.n2874 GND.n2873 0.0344674
R15566 GND.n2873 GND.n2850 0.0344674
R15567 GND.n3466 GND.n2850 0.0344674
R15568 GND.n3466 GND.n2853 0.0344674
R15569 GND.n2853 GND.n2852 0.0344674
R15570 GND.n2852 GND.n2831 0.0344674
R15571 GND.n3489 GND.n2831 0.0344674
R15572 GND.n3489 GND.n2832 0.0344674
R15573 GND.n3483 GND.n2832 0.0344674
R15574 GND.n3484 GND.n3483 0.0344674
R15575 GND.n3484 GND.n2779 0.0344674
R15576 GND.n5047 GND.n2779 0.0344674
R15577 GND.n5047 GND.n5046 0.0344674
R15578 GND.n5046 GND.n5045 0.0344674
R15579 GND.n5045 GND.n2549 0.0344674
R15580 GND.n5207 GND.n2549 0.0344674
R15581 GND.n5207 GND.n5206 0.0344674
R15582 GND.n5206 GND.n5205 0.0344674
R15583 GND.n5205 GND.n2553 0.0344674
R15584 GND.n5201 GND.n2553 0.0344674
R15585 GND.n5201 GND.n5200 0.0344674
R15586 GND.n5200 GND.n5199 0.0344674
R15587 GND.n5199 GND.n2561 0.0344674
R15588 GND.n5195 GND.n2561 0.0344674
R15589 GND.n5195 GND.n5194 0.0344674
R15590 GND.n5194 GND.n5193 0.0344674
R15591 GND.n5193 GND.n2569 0.0344674
R15592 GND.n5189 GND.n2569 0.0344674
R15593 GND.n5189 GND.n5188 0.0344674
R15594 GND.n5188 GND.n5187 0.0344674
R15595 GND.n5187 GND.n2503 0.0344674
R15596 GND.n5238 GND.n2503 0.0344674
R15597 GND.n5238 GND.n5237 0.0344674
R15598 GND.n5237 GND.n5236 0.0344674
R15599 GND.n5236 GND.n2483 0.0344674
R15600 GND.n5258 GND.n2483 0.0344674
R15601 GND.n5258 GND.n5257 0.0344674
R15602 GND.n5257 GND.n5256 0.0344674
R15603 GND.n5256 GND.n2463 0.0344674
R15604 GND.n5278 GND.n2463 0.0344674
R15605 GND.n5278 GND.n5277 0.0344674
R15606 GND.n5277 GND.n5276 0.0344674
R15607 GND.n5276 GND.n2443 0.0344674
R15608 GND.n5298 GND.n2443 0.0344674
R15609 GND.n5298 GND.n5297 0.0344674
R15610 GND.n5297 GND.n5296 0.0344674
R15611 GND.n5296 GND.n2423 0.0344674
R15612 GND.n5318 GND.n2423 0.0344674
R15613 GND.n5318 GND.n5317 0.0344674
R15614 GND.n5317 GND.n5316 0.0344674
R15615 GND.n5316 GND.n2403 0.0344674
R15616 GND.n5338 GND.n2403 0.0344674
R15617 GND.n5338 GND.n5337 0.0344674
R15618 GND.n5337 GND.n5336 0.0344674
R15619 GND.n5336 GND.n2383 0.0344674
R15620 GND.n5358 GND.n2383 0.0344674
R15621 GND.n5358 GND.n5357 0.0344674
R15622 GND.n5357 GND.n5356 0.0344674
R15623 GND.n5356 GND.n2363 0.0344674
R15624 GND.n5383 GND.n2363 0.0344674
R15625 GND.n5383 GND.n5382 0.0344674
R15626 GND.n5382 GND.n5381 0.0344674
R15627 GND.n5381 GND.n5377 0.0344674
R15628 GND.n5377 GND.n2335 0.0344674
R15629 GND.n5463 GND.n2335 0.0344674
R15630 GND.n5463 GND.n5462 0.0344674
R15631 GND.n5462 GND.n5461 0.0344674
R15632 GND.n5461 GND.n2316 0.0344674
R15633 GND.n5483 GND.n2316 0.0344674
R15634 GND.n5483 GND.n5482 0.0344674
R15635 GND.n5482 GND.n5481 0.0344674
R15636 GND.n5481 GND.n2296 0.0344674
R15637 GND.n5503 GND.n2296 0.0344674
R15638 GND.n5503 GND.n5502 0.0344674
R15639 GND.n5502 GND.n5501 0.0344674
R15640 GND.n5501 GND.n2276 0.0344674
R15641 GND.n5523 GND.n2276 0.0344674
R15642 GND.n5523 GND.n5522 0.0344674
R15643 GND.n5522 GND.n5521 0.0344674
R15644 GND.n5521 GND.n2256 0.0344674
R15645 GND.n5547 GND.n2256 0.0344674
R15646 GND.n5547 GND.n5546 0.0344674
R15647 GND.n5546 GND.n5545 0.0344674
R15648 GND.n5545 GND.n1732 0.0344674
R15649 GND.n5694 GND.n1732 0.0344674
R15650 VOUT.n11 VOUT.t4 133.702
R15651 VOUT.n9 VOUT.t10 133.702
R15652 VOUT.n3 VOUT.t3 129.918
R15653 VOUT.n1 VOUT.t1 129.918
R15654 VOUT.n3 VOUT.n2 124.469
R15655 VOUT.n1 VOUT.n0 124.469
R15656 VOUT.n9 VOUT.n8 120.684
R15657 VOUT.n11 VOUT.n10 120.683
R15658 VOUT.n23 VOUT.n21 81.7203
R15659 VOUT.n16 VOUT.n14 81.7203
R15660 VOUT.n39 VOUT.n37 81.7203
R15661 VOUT.n32 VOUT.n30 81.7203
R15662 VOUT.n27 VOUT.n26 76.7376
R15663 VOUT.n25 VOUT.n24 76.7376
R15664 VOUT.n23 VOUT.n22 76.7376
R15665 VOUT.n20 VOUT.n19 76.7376
R15666 VOUT.n18 VOUT.n17 76.7376
R15667 VOUT.n16 VOUT.n15 76.7376
R15668 VOUT.n39 VOUT.n38 76.7376
R15669 VOUT.n41 VOUT.n40 76.7376
R15670 VOUT.n43 VOUT.n42 76.7376
R15671 VOUT.n32 VOUT.n31 76.7376
R15672 VOUT.n34 VOUT.n33 76.7376
R15673 VOUT.n36 VOUT.n35 76.7376
R15674 VOUT.n28 VOUT.n20 10.2634
R15675 VOUT.n44 VOUT.n36 10.2634
R15676 VOUT.n12 VOUT.n9 9.72464
R15677 VOUT.n10 VOUT.t43 9.23488
R15678 VOUT.n10 VOUT.t2 9.23488
R15679 VOUT.n8 VOUT.t6 9.23488
R15680 VOUT.n8 VOUT.t8 9.23488
R15681 VOUT.n2 VOUT.t0 9.23488
R15682 VOUT.n2 VOUT.t9 9.23488
R15683 VOUT.n0 VOUT.t5 9.23488
R15684 VOUT.n0 VOUT.t7 9.23488
R15685 VOUT.n29 VOUT.n13 9.14649
R15686 VOUT.n13 VOUT.n12 9.04196
R15687 VOUT.n5 VOUT.n4 9.04196
R15688 VOUT.n29 VOUT.n28 8.65403
R15689 VOUT.n45 VOUT.n44 8.65403
R15690 VOUT.n28 VOUT.n27 7.89274
R15691 VOUT.n44 VOUT.n43 7.89274
R15692 VOUT.n4 VOUT.n1 7.8324
R15693 VOUT.n12 VOUT.n11 7.2936
R15694 VOUT.n26 VOUT.t34 5.87587
R15695 VOUT.n26 VOUT.t27 5.87587
R15696 VOUT.n24 VOUT.t25 5.87587
R15697 VOUT.n24 VOUT.t17 5.87587
R15698 VOUT.n22 VOUT.t15 5.87587
R15699 VOUT.n22 VOUT.t41 5.87587
R15700 VOUT.n21 VOUT.t39 5.87587
R15701 VOUT.n21 VOUT.t30 5.87587
R15702 VOUT.n19 VOUT.t20 5.87587
R15703 VOUT.n19 VOUT.t22 5.87587
R15704 VOUT.n17 VOUT.t28 5.87587
R15705 VOUT.n17 VOUT.t40 5.87587
R15706 VOUT.n15 VOUT.t36 5.87587
R15707 VOUT.n15 VOUT.t16 5.87587
R15708 VOUT.n14 VOUT.t23 5.87587
R15709 VOUT.n14 VOUT.t26 5.87587
R15710 VOUT.n37 VOUT.t37 5.87587
R15711 VOUT.n37 VOUT.t14 5.87587
R15712 VOUT.n38 VOUT.t24 5.87587
R15713 VOUT.n38 VOUT.t32 5.87587
R15714 VOUT.n40 VOUT.t33 5.87587
R15715 VOUT.n40 VOUT.t11 5.87587
R15716 VOUT.n42 VOUT.t35 5.87587
R15717 VOUT.n42 VOUT.t19 5.87587
R15718 VOUT.n30 VOUT.t12 5.87587
R15719 VOUT.n30 VOUT.t38 5.87587
R15720 VOUT.n31 VOUT.t29 5.87587
R15721 VOUT.n31 VOUT.t18 5.87587
R15722 VOUT.n33 VOUT.t21 5.87587
R15723 VOUT.n33 VOUT.t42 5.87587
R15724 VOUT.n35 VOUT.t13 5.87587
R15725 VOUT.n35 VOUT.t31 5.87587
R15726 VOUT.n45 VOUT.n29 5.43213
R15727 VOUT.n46 VOUT.n5 5.41399
R15728 VOUT.n4 VOUT.n3 5.40136
R15729 VOUT.n25 VOUT.n23 4.98326
R15730 VOUT.n27 VOUT.n25 4.98326
R15731 VOUT.n18 VOUT.n16 4.98326
R15732 VOUT.n20 VOUT.n18 4.98326
R15733 VOUT.n43 VOUT.n41 4.98326
R15734 VOUT.n41 VOUT.n39 4.98326
R15735 VOUT.n36 VOUT.n34 4.98326
R15736 VOUT.n34 VOUT.n32 4.98326
R15737 VOUT.n13 VOUT.n5 4.08198
R15738 VOUT.n46 VOUT.n45 3.71349
R15739 VOUT.n7 VOUT 3.39155
R15740 VOUT.n7 VOUT.n6 0.362917
R15741 VOUT.n46 VOUT.n7 0.330205
R15742 VOUT.n6 VOUT.t44 0.0919031
R15743 VOUT.n6 VOUT.t45 0.0200581
R15744 VOUT VOUT.n46 0.0099
R15745 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t4 146.666
R15746 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t5 146.27
R15747 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t2 109.995
R15748 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t0 107.835
R15749 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t3 97.0966
R15750 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t1 94.9397
R15751 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 5.38389
R15752 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n0 5.20416
R15753 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 4.34268
R15754 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 1.47354
R15755 DIFFPAIR_BIAS DIFFPAIR_BIAS.n4 0.68425
R15756 a_n1431_n2782.t0 a_n1431_n2782.t1 136.958
R15757 VN.n95 VN.t0 243.97
R15758 VN.n95 VN.t1 243.255
R15759 VN.n91 VN.n47 161.3
R15760 VN.n90 VN.n89 161.3
R15761 VN.n88 VN.n48 161.3
R15762 VN.n87 VN.n86 161.3
R15763 VN.n85 VN.n49 161.3
R15764 VN.n84 VN.n83 161.3
R15765 VN.n82 VN.n50 161.3
R15766 VN.n81 VN.n80 161.3
R15767 VN.n79 VN.n51 161.3
R15768 VN.n78 VN.n77 161.3
R15769 VN.n76 VN.n75 161.3
R15770 VN.n74 VN.n53 161.3
R15771 VN.n73 VN.n72 161.3
R15772 VN.n71 VN.n54 161.3
R15773 VN.n70 VN.n69 161.3
R15774 VN.n68 VN.n55 161.3
R15775 VN.n67 VN.n66 161.3
R15776 VN.n65 VN.n56 161.3
R15777 VN.n64 VN.n63 161.3
R15778 VN.n62 VN.n57 161.3
R15779 VN.n61 VN.n60 161.3
R15780 VN.n14 VN.n13 161.3
R15781 VN.n15 VN.n10 161.3
R15782 VN.n17 VN.n16 161.3
R15783 VN.n18 VN.n9 161.3
R15784 VN.n20 VN.n19 161.3
R15785 VN.n21 VN.n8 161.3
R15786 VN.n23 VN.n22 161.3
R15787 VN.n24 VN.n7 161.3
R15788 VN.n26 VN.n25 161.3
R15789 VN.n27 VN.n6 161.3
R15790 VN.n29 VN.n28 161.3
R15791 VN.n31 VN.n30 161.3
R15792 VN.n32 VN.n4 161.3
R15793 VN.n34 VN.n33 161.3
R15794 VN.n35 VN.n3 161.3
R15795 VN.n37 VN.n36 161.3
R15796 VN.n38 VN.n2 161.3
R15797 VN.n40 VN.n39 161.3
R15798 VN.n41 VN.n1 161.3
R15799 VN.n43 VN.n42 161.3
R15800 VN.n44 VN.n0 161.3
R15801 VN.n93 VN.n92 79.9798
R15802 VN.n46 VN.n45 79.9798
R15803 VN.n12 VN.n11 74.8596
R15804 VN.n59 VN.n58 74.8596
R15805 VN.n59 VN.t7 52.4204
R15806 VN.n12 VN.t5 52.4201
R15807 VN.n85 VN.n84 43.4072
R15808 VN.n38 VN.n37 43.4072
R15809 VN.n94 VN.n93 42.525
R15810 VN.n68 VN.n67 40.4934
R15811 VN.n69 VN.n68 40.4934
R15812 VN.n22 VN.n21 40.4934
R15813 VN.n21 VN.n20 40.4934
R15814 VN.n84 VN.n50 37.5796
R15815 VN.n37 VN.n3 37.5796
R15816 VN.n62 VN.n61 24.4675
R15817 VN.n63 VN.n62 24.4675
R15818 VN.n63 VN.n56 24.4675
R15819 VN.n67 VN.n56 24.4675
R15820 VN.n69 VN.n54 24.4675
R15821 VN.n73 VN.n54 24.4675
R15822 VN.n74 VN.n73 24.4675
R15823 VN.n75 VN.n74 24.4675
R15824 VN.n79 VN.n78 24.4675
R15825 VN.n80 VN.n79 24.4675
R15826 VN.n80 VN.n50 24.4675
R15827 VN.n86 VN.n85 24.4675
R15828 VN.n86 VN.n48 24.4675
R15829 VN.n90 VN.n48 24.4675
R15830 VN.n91 VN.n90 24.4675
R15831 VN.n44 VN.n43 24.4675
R15832 VN.n43 VN.n1 24.4675
R15833 VN.n39 VN.n1 24.4675
R15834 VN.n39 VN.n38 24.4675
R15835 VN.n33 VN.n3 24.4675
R15836 VN.n33 VN.n32 24.4675
R15837 VN.n32 VN.n31 24.4675
R15838 VN.n28 VN.n27 24.4675
R15839 VN.n27 VN.n26 24.4675
R15840 VN.n26 VN.n7 24.4675
R15841 VN.n22 VN.n7 24.4675
R15842 VN.n20 VN.n9 24.4675
R15843 VN.n16 VN.n9 24.4675
R15844 VN.n16 VN.n15 24.4675
R15845 VN.n15 VN.n14 24.4675
R15846 VN.n78 VN.n52 23.7335
R15847 VN.n31 VN.n5 23.7335
R15848 VN.n58 VN.t2 20.2548
R15849 VN.n52 VN.t8 20.2548
R15850 VN.n92 VN.t4 20.2548
R15851 VN.n45 VN.t9 20.2548
R15852 VN.n5 VN.t3 20.2548
R15853 VN.n11 VN.t6 20.2548
R15854 VN VN.n96 17.924
R15855 VN.n94 VN.n46 12.3129
R15856 VN.n96 VN.n95 5.04791
R15857 VN.n92 VN.n91 2.20253
R15858 VN.n45 VN.n44 2.20253
R15859 VN.n60 VN.n59 1.81424
R15860 VN.n13 VN.n12 1.81423
R15861 VN.n96 VN.n94 1.188
R15862 VN.n61 VN.n58 0.73451
R15863 VN.n75 VN.n52 0.73451
R15864 VN.n28 VN.n5 0.73451
R15865 VN.n14 VN.n11 0.73451
R15866 VN.n93 VN.n47 0.417535
R15867 VN.n46 VN.n0 0.417535
R15868 VN.n60 VN.n57 0.189894
R15869 VN.n64 VN.n57 0.189894
R15870 VN.n65 VN.n64 0.189894
R15871 VN.n66 VN.n65 0.189894
R15872 VN.n66 VN.n55 0.189894
R15873 VN.n70 VN.n55 0.189894
R15874 VN.n71 VN.n70 0.189894
R15875 VN.n72 VN.n71 0.189894
R15876 VN.n72 VN.n53 0.189894
R15877 VN.n76 VN.n53 0.189894
R15878 VN.n77 VN.n76 0.189894
R15879 VN.n77 VN.n51 0.189894
R15880 VN.n81 VN.n51 0.189894
R15881 VN.n82 VN.n81 0.189894
R15882 VN.n83 VN.n82 0.189894
R15883 VN.n83 VN.n49 0.189894
R15884 VN.n87 VN.n49 0.189894
R15885 VN.n88 VN.n87 0.189894
R15886 VN.n89 VN.n88 0.189894
R15887 VN.n89 VN.n47 0.189894
R15888 VN.n42 VN.n0 0.189894
R15889 VN.n42 VN.n41 0.189894
R15890 VN.n41 VN.n40 0.189894
R15891 VN.n40 VN.n2 0.189894
R15892 VN.n36 VN.n2 0.189894
R15893 VN.n36 VN.n35 0.189894
R15894 VN.n35 VN.n34 0.189894
R15895 VN.n34 VN.n4 0.189894
R15896 VN.n30 VN.n4 0.189894
R15897 VN.n30 VN.n29 0.189894
R15898 VN.n29 VN.n6 0.189894
R15899 VN.n25 VN.n6 0.189894
R15900 VN.n25 VN.n24 0.189894
R15901 VN.n24 VN.n23 0.189894
R15902 VN.n23 VN.n8 0.189894
R15903 VN.n19 VN.n8 0.189894
R15904 VN.n19 VN.n18 0.189894
R15905 VN.n18 VN.n17 0.189894
R15906 VN.n17 VN.n10 0.189894
R15907 VN.n13 VN.n10 0.189894
R15908 a_n4178_n267.n62 a_n4178_n267.n9 215.069
R15909 a_n4178_n267.n67 a_n4178_n267.n11 215.069
R15910 a_n4178_n267.n70 a_n4178_n267.n13 215.069
R15911 a_n4178_n267.n75 a_n4178_n267.n15 215.069
R15912 a_n4178_n267.n33 a_n4178_n267.n92 187.962
R15913 a_n4178_n267.n42 a_n4178_n267.n41 185
R15914 a_n4178_n267.n93 a_n4178_n267.n18 185
R15915 a_n4178_n267.n0 a_n4178_n267.n1 7.91264
R15916 a_n4178_n267.n34 a_n4178_n267.n87 187.962
R15917 a_n4178_n267.n44 a_n4178_n267.n43 185
R15918 a_n4178_n267.n88 a_n4178_n267.n20 185
R15919 a_n4178_n267.n2 a_n4178_n267.n3 7.91264
R15920 a_n4178_n267.n35 a_n4178_n267.n84 187.962
R15921 a_n4178_n267.n46 a_n4178_n267.n45 185
R15922 a_n4178_n267.n85 a_n4178_n267.n22 185
R15923 a_n4178_n267.n4 a_n4178_n267.n5 7.91264
R15924 a_n4178_n267.n36 a_n4178_n267.n79 187.962
R15925 a_n4178_n267.n48 a_n4178_n267.n47 185
R15926 a_n4178_n267.n80 a_n4178_n267.n24 185
R15927 a_n4178_n267.n6 a_n4178_n267.n7 7.91264
R15928 a_n4178_n267.n8 a_n4178_n267.n9 7.91264
R15929 a_n4178_n267.n62 a_n4178_n267.n26 185
R15930 a_n4178_n267.n50 a_n4178_n267.n49 185
R15931 a_n4178_n267.n37 a_n4178_n267.n61 187.962
R15932 a_n4178_n267.n10 a_n4178_n267.n11 7.91264
R15933 a_n4178_n267.n67 a_n4178_n267.n28 185
R15934 a_n4178_n267.n52 a_n4178_n267.n51 185
R15935 a_n4178_n267.n38 a_n4178_n267.n66 187.962
R15936 a_n4178_n267.n12 a_n4178_n267.n13 7.91264
R15937 a_n4178_n267.n70 a_n4178_n267.n30 185
R15938 a_n4178_n267.n54 a_n4178_n267.n53 185
R15939 a_n4178_n267.n39 a_n4178_n267.n69 187.962
R15940 a_n4178_n267.n14 a_n4178_n267.n15 7.91264
R15941 a_n4178_n267.n75 a_n4178_n267.n32 185
R15942 a_n4178_n267.n56 a_n4178_n267.n55 185
R15943 a_n4178_n267.n40 a_n4178_n267.n74 187.962
R15944 a_n4178_n267.n16 a_n4178_n267.t12 163.207
R15945 a_n4178_n267.t11 a_n4178_n267.n16 163.207
R15946 a_n4178_n267.t16 a_n4178_n267.n17 150.207
R15947 a_n4178_n267.t0 a_n4178_n267.n19 150.207
R15948 a_n4178_n267.t5 a_n4178_n267.n21 150.207
R15949 a_n4178_n267.t4 a_n4178_n267.n23 150.207
R15950 a_n4178_n267.n92 a_n4178_n267.n41 104.615
R15951 a_n4178_n267.n93 a_n4178_n267.n41 104.615
R15952 a_n4178_n267.n1 a_n4178_n267.n93 215.069
R15953 a_n4178_n267.n87 a_n4178_n267.n43 104.615
R15954 a_n4178_n267.n88 a_n4178_n267.n43 104.615
R15955 a_n4178_n267.n3 a_n4178_n267.n88 215.069
R15956 a_n4178_n267.n84 a_n4178_n267.n45 104.615
R15957 a_n4178_n267.n85 a_n4178_n267.n45 104.615
R15958 a_n4178_n267.n5 a_n4178_n267.n85 215.069
R15959 a_n4178_n267.n79 a_n4178_n267.n47 104.615
R15960 a_n4178_n267.n80 a_n4178_n267.n47 104.615
R15961 a_n4178_n267.n7 a_n4178_n267.n80 215.069
R15962 a_n4178_n267.n62 a_n4178_n267.n49 104.615
R15963 a_n4178_n267.n61 a_n4178_n267.n49 104.615
R15964 a_n4178_n267.n67 a_n4178_n267.n51 104.615
R15965 a_n4178_n267.n66 a_n4178_n267.n51 104.615
R15966 a_n4178_n267.n70 a_n4178_n267.n53 104.615
R15967 a_n4178_n267.n69 a_n4178_n267.n53 104.615
R15968 a_n4178_n267.n75 a_n4178_n267.n55 104.615
R15969 a_n4178_n267.n74 a_n4178_n267.n55 104.615
R15970 a_n4178_n267.n57 a_n4178_n267.n65 58.9186
R15971 a_n4178_n267.n73 a_n4178_n267.n72 58.9186
R15972 a_n4178_n267.n91 a_n4178_n267.n90 58.9185
R15973 a_n4178_n267.n59 a_n4178_n267.n83 58.9185
R15974 a_n4178_n267.n92 a_n4178_n267.t16 52.3082
R15975 a_n4178_n267.n87 a_n4178_n267.t0 52.3082
R15976 a_n4178_n267.n84 a_n4178_n267.t5 52.3082
R15977 a_n4178_n267.n79 a_n4178_n267.t4 52.3082
R15978 a_n4178_n267.n61 a_n4178_n267.t10 52.3082
R15979 a_n4178_n267.n66 a_n4178_n267.t7 52.3082
R15980 a_n4178_n267.n69 a_n4178_n267.t13 52.3082
R15981 a_n4178_n267.n74 a_n4178_n267.t2 52.3082
R15982 a_n4178_n267.n95 a_n4178_n267.n94 34.3187
R15983 a_n4178_n267.n60 a_n4178_n267.n89 34.3187
R15984 a_n4178_n267.n60 a_n4178_n267.n86 34.3187
R15985 a_n4178_n267.n82 a_n4178_n267.n81 34.3187
R15986 a_n4178_n267.n64 a_n4178_n267.n63 34.3187
R15987 a_n4178_n267.n58 a_n4178_n267.n68 34.3187
R15988 a_n4178_n267.n58 a_n4178_n267.n71 34.3187
R15989 a_n4178_n267.n77 a_n4178_n267.n76 34.3187
R15990 a_n4178_n267.n33 a_n4178_n267.n42 4.42678
R15991 a_n4178_n267.n34 a_n4178_n267.n44 4.42678
R15992 a_n4178_n267.n35 a_n4178_n267.n46 4.42678
R15993 a_n4178_n267.n36 a_n4178_n267.n48 4.42678
R15994 a_n4178_n267.n37 a_n4178_n267.n50 4.42678
R15995 a_n4178_n267.n38 a_n4178_n267.n52 4.42678
R15996 a_n4178_n267.n39 a_n4178_n267.n54 4.42678
R15997 a_n4178_n267.n40 a_n4178_n267.n56 4.42678
R15998 a_n4178_n267.n96 a_n4178_n267.n64 12.0944
R15999 a_n4178_n267.n78 a_n4178_n267.n77 12.0944
R16000 a_n4178_n267.n18 a_n4178_n267.n42 12.0247
R16001 a_n4178_n267.n20 a_n4178_n267.n44 12.0247
R16002 a_n4178_n267.n22 a_n4178_n267.n46 12.0247
R16003 a_n4178_n267.n24 a_n4178_n267.n48 12.0247
R16004 a_n4178_n267.n26 a_n4178_n267.n50 12.0247
R16005 a_n4178_n267.n28 a_n4178_n267.n52 12.0247
R16006 a_n4178_n267.n30 a_n4178_n267.n54 12.0247
R16007 a_n4178_n267.n32 a_n4178_n267.n56 12.0247
R16008 a_n4178_n267.n1 a_n4178_n267.n94 9.74451
R16009 a_n4178_n267.n3 a_n4178_n267.n89 9.74451
R16010 a_n4178_n267.n5 a_n4178_n267.n86 9.74451
R16011 a_n4178_n267.n7 a_n4178_n267.n81 9.74451
R16012 a_n4178_n267.n16 a_n4178_n267.n96 9.48742
R16013 a_n4178_n267.n94 a_n4178_n267.n17 9.45567
R16014 a_n4178_n267.n89 a_n4178_n267.n19 9.45567
R16015 a_n4178_n267.n86 a_n4178_n267.n21 9.45567
R16016 a_n4178_n267.n81 a_n4178_n267.n23 9.45567
R16017 a_n4178_n267.n63 a_n4178_n267.n25 9.45567
R16018 a_n4178_n267.n68 a_n4178_n267.n27 9.45567
R16019 a_n4178_n267.n71 a_n4178_n267.n29 9.45567
R16020 a_n4178_n267.n76 a_n4178_n267.n31 9.45567
R16021 a_n4178_n267.n82 a_n4178_n267.n78 7.43153
R16022 a_n4178_n267.n96 a_n4178_n267.n95 7.43153
R16023 a_n4178_n267.n90 a_n4178_n267.t15 5.01316
R16024 a_n4178_n267.n90 a_n4178_n267.t1 5.01316
R16025 a_n4178_n267.n83 a_n4178_n267.t8 5.01316
R16026 a_n4178_n267.n83 a_n4178_n267.t9 5.01316
R16027 a_n4178_n267.n65 a_n4178_n267.t3 5.01316
R16028 a_n4178_n267.n65 a_n4178_n267.t6 5.01316
R16029 a_n4178_n267.n72 a_n4178_n267.t17 5.01316
R16030 a_n4178_n267.n72 a_n4178_n267.t14 5.01316
R16031 a_n4178_n267.n25 a_n4178_n267.t10 150.207
R16032 a_n4178_n267.n27 a_n4178_n267.t7 150.207
R16033 a_n4178_n267.n29 a_n4178_n267.t13 150.207
R16034 a_n4178_n267.n31 a_n4178_n267.t2 150.207
R16035 a_n4178_n267.n17 a_n4178_n267.n0 3.91495
R16036 a_n4178_n267.n19 a_n4178_n267.n2 3.91495
R16037 a_n4178_n267.n21 a_n4178_n267.n4 3.91495
R16038 a_n4178_n267.n23 a_n4178_n267.n6 3.91495
R16039 a_n4178_n267.n25 a_n4178_n267.n8 3.91495
R16040 a_n4178_n267.n27 a_n4178_n267.n10 3.91495
R16041 a_n4178_n267.n29 a_n4178_n267.n12 3.91495
R16042 a_n4178_n267.n31 a_n4178_n267.n14 3.91495
R16043 a_n4178_n267.n32 a_n4178_n267.n14 3.6652
R16044 a_n4178_n267.n30 a_n4178_n267.n12 3.6652
R16045 a_n4178_n267.n28 a_n4178_n267.n10 3.6652
R16046 a_n4178_n267.n26 a_n4178_n267.n8 3.6652
R16047 a_n4178_n267.n24 a_n4178_n267.n6 3.6652
R16048 a_n4178_n267.n22 a_n4178_n267.n4 3.6652
R16049 a_n4178_n267.n20 a_n4178_n267.n2 3.6652
R16050 a_n4178_n267.n18 a_n4178_n267.n0 3.6652
R16051 a_n4178_n267.n78 a_n4178_n267.n16 9.7723
R16052 a_n4178_n267.n40 a_n4178_n267.n31 2.42091
R16053 a_n4178_n267.n39 a_n4178_n267.n29 2.42091
R16054 a_n4178_n267.n38 a_n4178_n267.n27 2.42091
R16055 a_n4178_n267.n37 a_n4178_n267.n25 2.42091
R16056 a_n4178_n267.n36 a_n4178_n267.n23 2.42091
R16057 a_n4178_n267.n35 a_n4178_n267.n21 2.42091
R16058 a_n4178_n267.n34 a_n4178_n267.n19 2.42091
R16059 a_n4178_n267.n33 a_n4178_n267.n17 2.42091
R16060 a_n4178_n267.n91 a_n4178_n267.n60 4.80653
R16061 a_n4178_n267.n73 a_n4178_n267.n58 4.80653
R16062 a_n4178_n267.n77 a_n4178_n267.n73 4.33671
R16063 a_n4178_n267.n58 a_n4178_n267.n57 4.33671
R16064 a_n4178_n267.n57 a_n4178_n267.n64 4.33671
R16065 a_n4178_n267.n59 a_n4178_n267.n82 4.33671
R16066 a_n4178_n267.n60 a_n4178_n267.n59 4.33671
R16067 a_n4178_n267.n95 a_n4178_n267.n91 4.33671
R16068 a_n4178_n267.n63 a_n4178_n267.n9 9.74451
R16069 a_n4178_n267.n68 a_n4178_n267.n11 9.74451
R16070 a_n4178_n267.n71 a_n4178_n267.n13 9.74451
R16071 a_n4178_n267.n76 a_n4178_n267.n15 9.74451
R16072 a_n12440_8296.n59 a_n12440_8296.n48 756.745
R16073 a_n12440_8296.n43 a_n12440_8296.n32 756.745
R16074 a_n12440_8296.n60 a_n12440_8296.n59 585
R16075 a_n12440_8296.n58 a_n12440_8296.n57 585
R16076 a_n12440_8296.n51 a_n12440_8296.n50 585
R16077 a_n12440_8296.n54 a_n12440_8296.n53 585
R16078 a_n12440_8296.n52 a_n12440_8296.n1 585
R16079 a_n12440_8296.n21 a_n12440_8296.n20 585
R16080 a_n12440_8296.n44 a_n12440_8296.n43 585
R16081 a_n12440_8296.n42 a_n12440_8296.n41 585
R16082 a_n12440_8296.n35 a_n12440_8296.n34 585
R16083 a_n12440_8296.n38 a_n12440_8296.n37 585
R16084 a_n12440_8296.n36 a_n12440_8296.n3 585
R16085 a_n12440_8296.n24 a_n12440_8296.n23 585
R16086 a_n12440_8296.n59 a_n12440_8296.n58 171.744
R16087 a_n12440_8296.n58 a_n12440_8296.n50 171.744
R16088 a_n12440_8296.n53 a_n12440_8296.n50 171.744
R16089 a_n12440_8296.n53 a_n12440_8296.n52 171.744
R16090 a_n12440_8296.n52 a_n12440_8296.n20 171.744
R16091 a_n12440_8296.n43 a_n12440_8296.n42 171.744
R16092 a_n12440_8296.n42 a_n12440_8296.n34 171.744
R16093 a_n12440_8296.n37 a_n12440_8296.n34 171.744
R16094 a_n12440_8296.n37 a_n12440_8296.n36 171.744
R16095 a_n12440_8296.n36 a_n12440_8296.n23 171.744
R16096 a_n12440_8296.n4 a_n12440_8296.n5 10.6209
R16097 a_n12440_8296.n6 a_n12440_8296.n7 10.6209
R16098 a_n12440_8296.n10 a_n12440_8296.n11 10.6209
R16099 a_n12440_8296.n8 a_n12440_8296.n9 10.6209
R16100 a_n12440_8296.n47 a_n12440_8296.n31 101.111
R16101 a_n12440_8296.n64 a_n12440_8296.n63 97.9127
R16102 a_n12440_8296.t1 a_n12440_8296.n20 85.8723
R16103 a_n12440_8296.t13 a_n12440_8296.n23 85.8723
R16104 a_n12440_8296.n79 a_n12440_8296.n78 77.7261
R16105 a_n12440_8296.n28 a_n12440_8296.n27 77.7101
R16106 a_n12440_8296.n28 a_n12440_8296.n26 77.7101
R16107 a_n12440_8296.n30 a_n12440_8296.n29 75.5974
R16108 a_n12440_8296.n12 a_n12440_8296.n13 28.0669
R16109 a_n12440_8296.n14 a_n12440_8296.n15 28.0669
R16110 a_n12440_8296.n16 a_n12440_8296.n17 28.0669
R16111 a_n12440_8296.n18 a_n12440_8296.n19 28.0669
R16112 a_n12440_8296.n68 a_n12440_8296.t23 54.133
R16113 a_n12440_8296.n66 a_n12440_8296.t18 54.133
R16114 a_n12440_8296.n73 a_n12440_8296.t20 54.1326
R16115 a_n12440_8296.n71 a_n12440_8296.t16 54.1326
R16116 a_n12440_8296.n64 a_n12440_8296.n62 52.6442
R16117 a_n12440_8296.n74 a_n12440_8296.n73 50.7346
R16118 a_n12440_8296.n72 a_n12440_8296.n71 50.7346
R16119 a_n12440_8296.n69 a_n12440_8296.n68 50.7346
R16120 a_n12440_8296.n67 a_n12440_8296.n66 50.7346
R16121 a_n12440_8296.n65 a_n12440_8296.n47 50.4221
R16122 a_n12440_8296.n47 a_n12440_8296.n46 49.446
R16123 a_n12440_8296.n30 a_n12440_8296.n28 46.4774
R16124 a_n12440_8296.n65 a_n12440_8296.n64 36.0305
R16125 a_n12440_8296.n5 a_n12440_8296.n13 97.3931
R16126 a_n12440_8296.n74 a_n12440_8296.n5 67.8434
R16127 a_n12440_8296.n7 a_n12440_8296.n15 97.3931
R16128 a_n12440_8296.n72 a_n12440_8296.n7 67.8434
R16129 a_n12440_8296.n11 a_n12440_8296.n69 67.8434
R16130 a_n12440_8296.n11 a_n12440_8296.n17 97.3931
R16131 a_n12440_8296.n9 a_n12440_8296.n67 67.8434
R16132 a_n12440_8296.n9 a_n12440_8296.n19 97.3931
R16133 a_n12440_8296.n74 a_n12440_8296.t21 20.8951
R16134 a_n12440_8296.n13 a_n12440_8296.t25 32.3586
R16135 a_n12440_8296.n72 a_n12440_8296.t15 20.8951
R16136 a_n12440_8296.n15 a_n12440_8296.t24 32.3586
R16137 a_n12440_8296.n69 a_n12440_8296.t22 20.8951
R16138 a_n12440_8296.n17 a_n12440_8296.t19 32.3586
R16139 a_n12440_8296.n67 a_n12440_8296.t17 20.8951
R16140 a_n12440_8296.n19 a_n12440_8296.t14 32.3586
R16141 a_n12440_8296.n22 a_n12440_8296.n21 5.32867
R16142 a_n12440_8296.n25 a_n12440_8296.n24 5.32867
R16143 a_n12440_8296.n1 a_n12440_8296.n21 12.8005
R16144 a_n12440_8296.n3 a_n12440_8296.n24 12.8005
R16145 a_n12440_8296.n78 a_n12440_8296.n77 12.3049
R16146 a_n12440_8296.n54 a_n12440_8296.n1 12.0247
R16147 a_n12440_8296.n38 a_n12440_8296.n3 12.0247
R16148 a_n12440_8296.n77 a_n12440_8296.n65 11.4887
R16149 a_n12440_8296.n55 a_n12440_8296.n51 11.249
R16150 a_n12440_8296.n39 a_n12440_8296.n35 11.249
R16151 a_n12440_8296.n57 a_n12440_8296.n56 10.4732
R16152 a_n12440_8296.n41 a_n12440_8296.n40 10.4732
R16153 a_n12440_8296.n60 a_n12440_8296.n49 9.69747
R16154 a_n12440_8296.n44 a_n12440_8296.n33 9.69747
R16155 a_n12440_8296.n62 a_n12440_8296.n0 9.45567
R16156 a_n12440_8296.n46 a_n12440_8296.n2 9.45567
R16157 a_n12440_8296.n76 a_n12440_8296.n70 9.30235
R16158 a_n12440_8296.n0 a_n12440_8296.n61 9.3005
R16159 a_n12440_8296.n49 a_n12440_8296.n0 9.3005
R16160 a_n12440_8296.n56 a_n12440_8296.n0 9.3005
R16161 a_n12440_8296.n0 a_n12440_8296.n55 9.3005
R16162 a_n12440_8296.n2 a_n12440_8296.n45 9.3005
R16163 a_n12440_8296.n33 a_n12440_8296.n2 9.3005
R16164 a_n12440_8296.n40 a_n12440_8296.n2 9.3005
R16165 a_n12440_8296.n2 a_n12440_8296.n39 9.3005
R16166 a_n12440_8296.n61 a_n12440_8296.n48 8.92171
R16167 a_n12440_8296.n45 a_n12440_8296.n32 8.92171
R16168 a_n12440_8296.n76 a_n12440_8296.n75 8.63777
R16169 a_n12440_8296.n75 a_n12440_8296.n14 7.44377
R16170 a_n12440_8296.n70 a_n12440_8296.n18 7.44377
R16171 a_n12440_8296.n63 a_n12440_8296.t0 6.12197
R16172 a_n12440_8296.n63 a_n12440_8296.t11 6.12197
R16173 a_n12440_8296.n31 a_n12440_8296.t12 6.12197
R16174 a_n12440_8296.n31 a_n12440_8296.t2 6.12197
R16175 a_n12440_8296.n75 a_n12440_8296.n12 5.29225
R16176 a_n12440_8296.n70 a_n12440_8296.n16 5.29225
R16177 a_n12440_8296.n62 a_n12440_8296.n48 5.04292
R16178 a_n12440_8296.n46 a_n12440_8296.n32 5.04292
R16179 a_n12440_8296.n29 a_n12440_8296.t4 5.01316
R16180 a_n12440_8296.n29 a_n12440_8296.t8 5.01316
R16181 a_n12440_8296.n27 a_n12440_8296.t6 5.01316
R16182 a_n12440_8296.n27 a_n12440_8296.t7 5.01316
R16183 a_n12440_8296.n26 a_n12440_8296.t3 5.01316
R16184 a_n12440_8296.n26 a_n12440_8296.t9 5.01316
R16185 a_n12440_8296.n79 a_n12440_8296.t5 5.01316
R16186 a_n12440_8296.t10 a_n12440_8296.n79 5.01316
R16187 a_n12440_8296.n61 a_n12440_8296.n60 4.26717
R16188 a_n12440_8296.n45 a_n12440_8296.n44 4.26717
R16189 a_n12440_8296.n22 a_n12440_8296.t1 329.901
R16190 a_n12440_8296.n25 a_n12440_8296.t13 329.901
R16191 a_n12440_8296.n3 a_n12440_8296.n2 10.4641
R16192 a_n12440_8296.n1 a_n12440_8296.n0 10.4641
R16193 a_n12440_8296.n57 a_n12440_8296.n49 3.49141
R16194 a_n12440_8296.n41 a_n12440_8296.n33 3.49141
R16195 a_n12440_8296.n77 a_n12440_8296.n76 3.4105
R16196 a_n12440_8296.n56 a_n12440_8296.n51 2.71565
R16197 a_n12440_8296.n40 a_n12440_8296.n35 2.71565
R16198 a_n12440_8296.n78 a_n12440_8296.n30 2.12915
R16199 a_n12440_8296.n10 a_n12440_8296.n68 2.01978
R16200 a_n12440_8296.n8 a_n12440_8296.n66 2.01978
R16201 a_n12440_8296.n4 a_n12440_8296.n73 2.01976
R16202 a_n12440_8296.n6 a_n12440_8296.n71 2.01976
R16203 a_n12440_8296.n25 a_n12440_8296.n2 1.98613
R16204 a_n12440_8296.n22 a_n12440_8296.n0 1.98613
R16205 a_n12440_8296.n55 a_n12440_8296.n54 1.93989
R16206 a_n12440_8296.n39 a_n12440_8296.n38 1.93989
R16207 a_n12440_8296.n16 a_n12440_8296.n10 1.74306
R16208 a_n12440_8296.n18 a_n12440_8296.n8 1.74306
R16209 a_n12440_8296.n14 a_n12440_8296.n6 1.74306
R16210 a_n12440_8296.n12 a_n12440_8296.n4 1.74306
R16211 VDD.n2625 VDD.n90 453.659
R16212 VDD.n2621 VDD.n91 453.659
R16213 VDD.n2473 VDD.n252 453.659
R16214 VDD.n2470 VDD.n250 453.659
R16215 VDD.n1148 VDD.n724 453.659
R16216 VDD.n1221 VDD.n714 453.659
R16217 VDD.n950 VDD.n865 453.659
R16218 VDD.n948 VDD.n867 453.659
R16219 VDD.n1970 VDD.t81 328.182
R16220 VDD.n292 VDD.t71 328.182
R16221 VDD.n1234 VDD.t37 328.182
R16222 VDD.n511 VDD.t57 328.182
R16223 VDD.n1813 VDD.t51 328.182
R16224 VDD.n2279 VDD.t54 328.182
R16225 VDD.n1374 VDD.t78 328.182
R16226 VDD.n1689 VDD.t46 328.182
R16227 VDD.n2106 VDD.n1959 320.488
R16228 VDD.n2386 VDD.n290 320.488
R16229 VDD.n2344 VDD.n2343 320.488
R16230 VDD.n2062 VDD.n1810 320.488
R16231 VDD.n1796 VDD.n509 320.488
R16232 VDD.n1754 VDD.n1753 320.488
R16233 VDD.n1362 VDD.n697 320.488
R16234 VDD.n1516 VDD.n699 320.488
R16235 VDD.n2322 VDD.n2321 320.488
R16236 VDD.n2396 VDD.n281 320.488
R16237 VDD.n1958 VDD.n1811 320.488
R16238 VDD.n2108 VDD.n477 320.488
R16239 VDD.n1732 VDD.n1731 320.488
R16240 VDD.n1806 VDD.n501 320.488
R16241 VDD.n1468 VDD.n698 320.488
R16242 VDD.n1518 VDD.n696 320.488
R16243 VDD.n1971 VDD.t80 256.231
R16244 VDD.n293 VDD.t72 256.231
R16245 VDD.n1235 VDD.t36 256.231
R16246 VDD.n512 VDD.t58 256.231
R16247 VDD.n1814 VDD.t50 256.231
R16248 VDD.n2280 VDD.t55 256.231
R16249 VDD.n1375 VDD.t77 256.231
R16250 VDD.n1690 VDD.t47 256.231
R16251 VDD.n1970 VDD.t79 246.845
R16252 VDD.n292 VDD.t70 246.845
R16253 VDD.n1234 VDD.t34 246.845
R16254 VDD.n511 VDD.t56 246.845
R16255 VDD.n1813 VDD.t48 246.845
R16256 VDD.n2279 VDD.t52 246.845
R16257 VDD.n1374 VDD.t76 246.845
R16258 VDD.n1689 VDD.t44 246.845
R16259 VDD.n906 VDD.t26 230.429
R16260 VDD.n929 VDD.t38 230.429
R16261 VDD.n2420 VDD.t73 230.429
R16262 VDD.n255 VDD.t66 230.429
R16263 VDD.n103 VDD.t30 230.429
R16264 VDD.n111 VDD.t41 230.429
R16265 VDD.n1161 VDD.t63 230.429
R16266 VDD.n715 VDD.t59 230.429
R16267 VDD.n906 VDD.t29 213.767
R16268 VDD.n929 VDD.t40 213.767
R16269 VDD.n2420 VDD.t75 213.767
R16270 VDD.n255 VDD.t69 213.767
R16271 VDD.n103 VDD.t32 213.767
R16272 VDD.n111 VDD.t42 213.767
R16273 VDD.n1161 VDD.t64 213.767
R16274 VDD.n715 VDD.t61 213.767
R16275 VDD.t109 VDD.n1223 206.537
R16276 VDD.n2472 VDD.t84 206.537
R16277 VDD.n1733 VDD.n1732 185
R16278 VDD.n1732 VDD.n478 185
R16279 VDD.n1734 VDD.n507 185
R16280 VDD.n1801 VDD.n507 185
R16281 VDD.n1736 VDD.n1735 185
R16282 VDD.n1735 VDD.n505 185
R16283 VDD.n1737 VDD.n518 185
R16284 VDD.n1747 VDD.n518 185
R16285 VDD.n1738 VDD.n526 185
R16286 VDD.n526 VDD.n516 185
R16287 VDD.n1740 VDD.n1739 185
R16288 VDD.n1741 VDD.n1740 185
R16289 VDD.n1688 VDD.n525 185
R16290 VDD.n525 VDD.n522 185
R16291 VDD.n1687 VDD.n1686 185
R16292 VDD.n1686 VDD.n1685 185
R16293 VDD.n528 VDD.n527 185
R16294 VDD.n529 VDD.n528 185
R16295 VDD.n1678 VDD.n1677 185
R16296 VDD.n1679 VDD.n1678 185
R16297 VDD.n1676 VDD.n538 185
R16298 VDD.n538 VDD.n535 185
R16299 VDD.n1675 VDD.n1674 185
R16300 VDD.n1674 VDD.n1673 185
R16301 VDD.n540 VDD.n539 185
R16302 VDD.n541 VDD.n540 185
R16303 VDD.n1666 VDD.n1665 185
R16304 VDD.n1667 VDD.n1666 185
R16305 VDD.n1664 VDD.n550 185
R16306 VDD.n550 VDD.n547 185
R16307 VDD.n1663 VDD.n1662 185
R16308 VDD.n1662 VDD.n1661 185
R16309 VDD.n552 VDD.n551 185
R16310 VDD.n561 VDD.n552 185
R16311 VDD.n1654 VDD.n1653 185
R16312 VDD.n1655 VDD.n1654 185
R16313 VDD.n1652 VDD.n562 185
R16314 VDD.n562 VDD.n558 185
R16315 VDD.n1651 VDD.n1650 185
R16316 VDD.n1650 VDD.n1649 185
R16317 VDD.n564 VDD.n563 185
R16318 VDD.n565 VDD.n564 185
R16319 VDD.n1642 VDD.n1641 185
R16320 VDD.n1643 VDD.n1642 185
R16321 VDD.n1640 VDD.n574 185
R16322 VDD.n574 VDD.n571 185
R16323 VDD.n1639 VDD.n1638 185
R16324 VDD.n1638 VDD.n1637 185
R16325 VDD.n576 VDD.n575 185
R16326 VDD.n577 VDD.n576 185
R16327 VDD.n1630 VDD.n1629 185
R16328 VDD.n1631 VDD.n1630 185
R16329 VDD.n1628 VDD.n586 185
R16330 VDD.n586 VDD.n583 185
R16331 VDD.n1627 VDD.n1626 185
R16332 VDD.n1626 VDD.n1625 185
R16333 VDD.n588 VDD.n587 185
R16334 VDD.n589 VDD.n588 185
R16335 VDD.n1618 VDD.n1617 185
R16336 VDD.n1619 VDD.n1618 185
R16337 VDD.n1616 VDD.n598 185
R16338 VDD.n598 VDD.n595 185
R16339 VDD.n1615 VDD.n1614 185
R16340 VDD.n1614 VDD.n1613 185
R16341 VDD.n600 VDD.n599 185
R16342 VDD.n609 VDD.n600 185
R16343 VDD.n1606 VDD.n1605 185
R16344 VDD.n1607 VDD.n1606 185
R16345 VDD.n1604 VDD.n610 185
R16346 VDD.n610 VDD.n606 185
R16347 VDD.n1603 VDD.n1602 185
R16348 VDD.n1602 VDD.n1601 185
R16349 VDD.n612 VDD.n611 185
R16350 VDD.n613 VDD.n612 185
R16351 VDD.n1594 VDD.n1593 185
R16352 VDD.n1595 VDD.n1594 185
R16353 VDD.n1592 VDD.n621 185
R16354 VDD.n627 VDD.n621 185
R16355 VDD.n1591 VDD.n1590 185
R16356 VDD.n1590 VDD.n1589 185
R16357 VDD.n623 VDD.n622 185
R16358 VDD.n624 VDD.n623 185
R16359 VDD.n1582 VDD.n1581 185
R16360 VDD.n1583 VDD.n1582 185
R16361 VDD.n1580 VDD.n634 185
R16362 VDD.n634 VDD.n631 185
R16363 VDD.n1579 VDD.n1578 185
R16364 VDD.n1578 VDD.n1577 185
R16365 VDD.n636 VDD.n635 185
R16366 VDD.n637 VDD.n636 185
R16367 VDD.n1570 VDD.n1569 185
R16368 VDD.n1571 VDD.n1570 185
R16369 VDD.n1568 VDD.n646 185
R16370 VDD.n646 VDD.n643 185
R16371 VDD.n1567 VDD.n1566 185
R16372 VDD.n1566 VDD.n1565 185
R16373 VDD.n648 VDD.n647 185
R16374 VDD.n649 VDD.n648 185
R16375 VDD.n1558 VDD.n1557 185
R16376 VDD.n1559 VDD.n1558 185
R16377 VDD.n1556 VDD.n658 185
R16378 VDD.n658 VDD.n655 185
R16379 VDD.n1555 VDD.n1554 185
R16380 VDD.n1554 VDD.n1553 185
R16381 VDD.n660 VDD.n659 185
R16382 VDD.n661 VDD.n660 185
R16383 VDD.n1546 VDD.n1545 185
R16384 VDD.n1547 VDD.n1546 185
R16385 VDD.n1544 VDD.n669 185
R16386 VDD.n675 VDD.n669 185
R16387 VDD.n1543 VDD.n1542 185
R16388 VDD.n1542 VDD.n1541 185
R16389 VDD.n671 VDD.n670 185
R16390 VDD.n672 VDD.n671 185
R16391 VDD.n1534 VDD.n1533 185
R16392 VDD.n1535 VDD.n1534 185
R16393 VDD.n1532 VDD.n682 185
R16394 VDD.n682 VDD.n679 185
R16395 VDD.n1531 VDD.n1530 185
R16396 VDD.n1530 VDD.n1529 185
R16397 VDD.n684 VDD.n683 185
R16398 VDD.n685 VDD.n684 185
R16399 VDD.n1522 VDD.n1521 185
R16400 VDD.n1523 VDD.n1522 185
R16401 VDD.n1520 VDD.n694 185
R16402 VDD.n694 VDD.n691 185
R16403 VDD.n1519 VDD.n1518 185
R16404 VDD.n1518 VDD.n1517 185
R16405 VDD.n696 VDD.n695 185
R16406 VDD.n1508 VDD.n1507 185
R16407 VDD.n1506 VDD.n1373 185
R16408 VDD.n1505 VDD.n1504 185
R16409 VDD.n1503 VDD.n1502 185
R16410 VDD.n1501 VDD.n1500 185
R16411 VDD.n1499 VDD.n1498 185
R16412 VDD.n1497 VDD.n1496 185
R16413 VDD.n1495 VDD.n1494 185
R16414 VDD.n1493 VDD.n1492 185
R16415 VDD.n1491 VDD.n1490 185
R16416 VDD.n1489 VDD.n1488 185
R16417 VDD.n1487 VDD.n1486 185
R16418 VDD.n1485 VDD.n1484 185
R16419 VDD.n1483 VDD.n1482 185
R16420 VDD.n1481 VDD.n1480 185
R16421 VDD.n1479 VDD.n1478 185
R16422 VDD.n1477 VDD.n1476 185
R16423 VDD.n1475 VDD.n1474 185
R16424 VDD.n1473 VDD.n1472 185
R16425 VDD.n1471 VDD.n1470 185
R16426 VDD.n1469 VDD.n1468 185
R16427 VDD.n1806 VDD.n1805 185
R16428 VDD.n502 VDD.n500 185
R16429 VDD.n1693 VDD.n1692 185
R16430 VDD.n1695 VDD.n1694 185
R16431 VDD.n1697 VDD.n1696 185
R16432 VDD.n1699 VDD.n1698 185
R16433 VDD.n1701 VDD.n1700 185
R16434 VDD.n1703 VDD.n1702 185
R16435 VDD.n1705 VDD.n1704 185
R16436 VDD.n1707 VDD.n1706 185
R16437 VDD.n1709 VDD.n1708 185
R16438 VDD.n1711 VDD.n1710 185
R16439 VDD.n1713 VDD.n1712 185
R16440 VDD.n1715 VDD.n1714 185
R16441 VDD.n1717 VDD.n1716 185
R16442 VDD.n1719 VDD.n1718 185
R16443 VDD.n1721 VDD.n1720 185
R16444 VDD.n1723 VDD.n1722 185
R16445 VDD.n1725 VDD.n1724 185
R16446 VDD.n1727 VDD.n1726 185
R16447 VDD.n1729 VDD.n1728 185
R16448 VDD.n1731 VDD.n1730 185
R16449 VDD.n1804 VDD.n501 185
R16450 VDD.n501 VDD.n478 185
R16451 VDD.n1803 VDD.n1802 185
R16452 VDD.n1802 VDD.n1801 185
R16453 VDD.n504 VDD.n503 185
R16454 VDD.n505 VDD.n504 185
R16455 VDD.n1377 VDD.n517 185
R16456 VDD.n1747 VDD.n517 185
R16457 VDD.n1379 VDD.n1378 185
R16458 VDD.n1378 VDD.n516 185
R16459 VDD.n1380 VDD.n524 185
R16460 VDD.n1741 VDD.n524 185
R16461 VDD.n1382 VDD.n1381 185
R16462 VDD.n1381 VDD.n522 185
R16463 VDD.n1383 VDD.n531 185
R16464 VDD.n1685 VDD.n531 185
R16465 VDD.n1385 VDD.n1384 185
R16466 VDD.n1384 VDD.n529 185
R16467 VDD.n1386 VDD.n537 185
R16468 VDD.n1679 VDD.n537 185
R16469 VDD.n1388 VDD.n1387 185
R16470 VDD.n1387 VDD.n535 185
R16471 VDD.n1389 VDD.n543 185
R16472 VDD.n1673 VDD.n543 185
R16473 VDD.n1391 VDD.n1390 185
R16474 VDD.n1390 VDD.n541 185
R16475 VDD.n1392 VDD.n549 185
R16476 VDD.n1667 VDD.n549 185
R16477 VDD.n1394 VDD.n1393 185
R16478 VDD.n1393 VDD.n547 185
R16479 VDD.n1395 VDD.n554 185
R16480 VDD.n1661 VDD.n554 185
R16481 VDD.n1397 VDD.n1396 185
R16482 VDD.n1396 VDD.n561 185
R16483 VDD.n1398 VDD.n560 185
R16484 VDD.n1655 VDD.n560 185
R16485 VDD.n1400 VDD.n1399 185
R16486 VDD.n1399 VDD.n558 185
R16487 VDD.n1401 VDD.n567 185
R16488 VDD.n1649 VDD.n567 185
R16489 VDD.n1403 VDD.n1402 185
R16490 VDD.n1402 VDD.n565 185
R16491 VDD.n1404 VDD.n573 185
R16492 VDD.n1643 VDD.n573 185
R16493 VDD.n1406 VDD.n1405 185
R16494 VDD.n1405 VDD.n571 185
R16495 VDD.n1407 VDD.n579 185
R16496 VDD.n1637 VDD.n579 185
R16497 VDD.n1409 VDD.n1408 185
R16498 VDD.n1408 VDD.n577 185
R16499 VDD.n1410 VDD.n585 185
R16500 VDD.n1631 VDD.n585 185
R16501 VDD.n1412 VDD.n1411 185
R16502 VDD.n1411 VDD.n583 185
R16503 VDD.n1413 VDD.n591 185
R16504 VDD.n1625 VDD.n591 185
R16505 VDD.n1415 VDD.n1414 185
R16506 VDD.n1414 VDD.n589 185
R16507 VDD.n1416 VDD.n597 185
R16508 VDD.n1619 VDD.n597 185
R16509 VDD.n1418 VDD.n1417 185
R16510 VDD.n1417 VDD.n595 185
R16511 VDD.n1419 VDD.n602 185
R16512 VDD.n1613 VDD.n602 185
R16513 VDD.n1421 VDD.n1420 185
R16514 VDD.n1420 VDD.n609 185
R16515 VDD.n1422 VDD.n608 185
R16516 VDD.n1607 VDD.n608 185
R16517 VDD.n1424 VDD.n1423 185
R16518 VDD.n1423 VDD.n606 185
R16519 VDD.n1425 VDD.n615 185
R16520 VDD.n1601 VDD.n615 185
R16521 VDD.n1427 VDD.n1426 185
R16522 VDD.n1426 VDD.n613 185
R16523 VDD.n1428 VDD.n620 185
R16524 VDD.n1595 VDD.n620 185
R16525 VDD.n1430 VDD.n1429 185
R16526 VDD.n1429 VDD.n627 185
R16527 VDD.n1431 VDD.n626 185
R16528 VDD.n1589 VDD.n626 185
R16529 VDD.n1433 VDD.n1432 185
R16530 VDD.n1432 VDD.n624 185
R16531 VDD.n1434 VDD.n633 185
R16532 VDD.n1583 VDD.n633 185
R16533 VDD.n1436 VDD.n1435 185
R16534 VDD.n1435 VDD.n631 185
R16535 VDD.n1437 VDD.n639 185
R16536 VDD.n1577 VDD.n639 185
R16537 VDD.n1439 VDD.n1438 185
R16538 VDD.n1438 VDD.n637 185
R16539 VDD.n1440 VDD.n645 185
R16540 VDD.n1571 VDD.n645 185
R16541 VDD.n1442 VDD.n1441 185
R16542 VDD.n1441 VDD.n643 185
R16543 VDD.n1443 VDD.n651 185
R16544 VDD.n1565 VDD.n651 185
R16545 VDD.n1445 VDD.n1444 185
R16546 VDD.n1444 VDD.n649 185
R16547 VDD.n1446 VDD.n657 185
R16548 VDD.n1559 VDD.n657 185
R16549 VDD.n1448 VDD.n1447 185
R16550 VDD.n1447 VDD.n655 185
R16551 VDD.n1449 VDD.n663 185
R16552 VDD.n1553 VDD.n663 185
R16553 VDD.n1451 VDD.n1450 185
R16554 VDD.n1450 VDD.n661 185
R16555 VDD.n1452 VDD.n668 185
R16556 VDD.n1547 VDD.n668 185
R16557 VDD.n1454 VDD.n1453 185
R16558 VDD.n1453 VDD.n675 185
R16559 VDD.n1455 VDD.n674 185
R16560 VDD.n1541 VDD.n674 185
R16561 VDD.n1457 VDD.n1456 185
R16562 VDD.n1456 VDD.n672 185
R16563 VDD.n1458 VDD.n681 185
R16564 VDD.n1535 VDD.n681 185
R16565 VDD.n1460 VDD.n1459 185
R16566 VDD.n1459 VDD.n679 185
R16567 VDD.n1461 VDD.n687 185
R16568 VDD.n1529 VDD.n687 185
R16569 VDD.n1463 VDD.n1462 185
R16570 VDD.n1462 VDD.n685 185
R16571 VDD.n1464 VDD.n693 185
R16572 VDD.n1523 VDD.n693 185
R16573 VDD.n1466 VDD.n1465 185
R16574 VDD.n1465 VDD.n691 185
R16575 VDD.n1467 VDD.n698 185
R16576 VDD.n1517 VDD.n698 185
R16577 VDD.n2323 VDD.n2322 185
R16578 VDD.n2322 VDD.n287 185
R16579 VDD.n2324 VDD.n288 185
R16580 VDD.n2391 VDD.n288 185
R16581 VDD.n2326 VDD.n2325 185
R16582 VDD.n2325 VDD.n285 185
R16583 VDD.n2327 VDD.n299 185
R16584 VDD.n2337 VDD.n299 185
R16585 VDD.n2328 VDD.n307 185
R16586 VDD.n307 VDD.n297 185
R16587 VDD.n2330 VDD.n2329 185
R16588 VDD.n2331 VDD.n2330 185
R16589 VDD.n2278 VDD.n306 185
R16590 VDD.n306 VDD.n303 185
R16591 VDD.n2277 VDD.n2276 185
R16592 VDD.n2276 VDD.n2275 185
R16593 VDD.n309 VDD.n308 185
R16594 VDD.n310 VDD.n309 185
R16595 VDD.n2268 VDD.n2267 185
R16596 VDD.n2269 VDD.n2268 185
R16597 VDD.n2266 VDD.n318 185
R16598 VDD.n324 VDD.n318 185
R16599 VDD.n2265 VDD.n2264 185
R16600 VDD.n2264 VDD.n2263 185
R16601 VDD.n320 VDD.n319 185
R16602 VDD.n321 VDD.n320 185
R16603 VDD.n2256 VDD.n2255 185
R16604 VDD.n2257 VDD.n2256 185
R16605 VDD.n2254 VDD.n331 185
R16606 VDD.n331 VDD.n328 185
R16607 VDD.n2253 VDD.n2252 185
R16608 VDD.n2252 VDD.n2251 185
R16609 VDD.n333 VDD.n332 185
R16610 VDD.n334 VDD.n333 185
R16611 VDD.n2244 VDD.n2243 185
R16612 VDD.n2245 VDD.n2244 185
R16613 VDD.n2242 VDD.n343 185
R16614 VDD.n343 VDD.n340 185
R16615 VDD.n2241 VDD.n2240 185
R16616 VDD.n2240 VDD.n2239 185
R16617 VDD.n345 VDD.n344 185
R16618 VDD.n346 VDD.n345 185
R16619 VDD.n2232 VDD.n2231 185
R16620 VDD.n2233 VDD.n2232 185
R16621 VDD.n2230 VDD.n355 185
R16622 VDD.n355 VDD.n352 185
R16623 VDD.n2229 VDD.n2228 185
R16624 VDD.n2228 VDD.n2227 185
R16625 VDD.n357 VDD.n356 185
R16626 VDD.n358 VDD.n357 185
R16627 VDD.n2220 VDD.n2219 185
R16628 VDD.n2221 VDD.n2220 185
R16629 VDD.n2218 VDD.n366 185
R16630 VDD.n372 VDD.n366 185
R16631 VDD.n2217 VDD.n2216 185
R16632 VDD.n2216 VDD.n2215 185
R16633 VDD.n368 VDD.n367 185
R16634 VDD.n369 VDD.n368 185
R16635 VDD.n2208 VDD.n2207 185
R16636 VDD.n2209 VDD.n2208 185
R16637 VDD.n2206 VDD.n379 185
R16638 VDD.n379 VDD.n376 185
R16639 VDD.n2205 VDD.n2204 185
R16640 VDD.n2204 VDD.n2203 185
R16641 VDD.n381 VDD.n380 185
R16642 VDD.n390 VDD.n381 185
R16643 VDD.n2196 VDD.n2195 185
R16644 VDD.n2197 VDD.n2196 185
R16645 VDD.n2194 VDD.n391 185
R16646 VDD.n391 VDD.n387 185
R16647 VDD.n2193 VDD.n2192 185
R16648 VDD.n2192 VDD.n2191 185
R16649 VDD.n393 VDD.n392 185
R16650 VDD.n394 VDD.n393 185
R16651 VDD.n2184 VDD.n2183 185
R16652 VDD.n2185 VDD.n2184 185
R16653 VDD.n2182 VDD.n403 185
R16654 VDD.n403 VDD.n400 185
R16655 VDD.n2181 VDD.n2180 185
R16656 VDD.n2180 VDD.n2179 185
R16657 VDD.n405 VDD.n404 185
R16658 VDD.n406 VDD.n405 185
R16659 VDD.n2172 VDD.n2171 185
R16660 VDD.n2173 VDD.n2172 185
R16661 VDD.n2170 VDD.n415 185
R16662 VDD.n415 VDD.n412 185
R16663 VDD.n2169 VDD.n2168 185
R16664 VDD.n2168 VDD.n2167 185
R16665 VDD.n417 VDD.n416 185
R16666 VDD.n418 VDD.n417 185
R16667 VDD.n2160 VDD.n2159 185
R16668 VDD.n2161 VDD.n2160 185
R16669 VDD.n2158 VDD.n427 185
R16670 VDD.n427 VDD.n424 185
R16671 VDD.n2157 VDD.n2156 185
R16672 VDD.n2156 VDD.n2155 185
R16673 VDD.n429 VDD.n428 185
R16674 VDD.n438 VDD.n429 185
R16675 VDD.n2148 VDD.n2147 185
R16676 VDD.n2149 VDD.n2148 185
R16677 VDD.n2146 VDD.n439 185
R16678 VDD.n439 VDD.n435 185
R16679 VDD.n2145 VDD.n2144 185
R16680 VDD.n2144 VDD.n2143 185
R16681 VDD.n441 VDD.n440 185
R16682 VDD.n442 VDD.n441 185
R16683 VDD.n2136 VDD.n2135 185
R16684 VDD.n2137 VDD.n2136 185
R16685 VDD.n2134 VDD.n451 185
R16686 VDD.n451 VDD.n448 185
R16687 VDD.n2133 VDD.n2132 185
R16688 VDD.n2132 VDD.n2131 185
R16689 VDD.n453 VDD.n452 185
R16690 VDD.n454 VDD.n453 185
R16691 VDD.n2124 VDD.n2123 185
R16692 VDD.n2125 VDD.n2124 185
R16693 VDD.n2122 VDD.n463 185
R16694 VDD.n463 VDD.n460 185
R16695 VDD.n2121 VDD.n2120 185
R16696 VDD.n2120 VDD.n2119 185
R16697 VDD.n465 VDD.n464 185
R16698 VDD.n466 VDD.n465 185
R16699 VDD.n2112 VDD.n2111 185
R16700 VDD.n2113 VDD.n2112 185
R16701 VDD.n2110 VDD.n475 185
R16702 VDD.n475 VDD.n472 185
R16703 VDD.n2109 VDD.n2108 185
R16704 VDD.n2108 VDD.n2107 185
R16705 VDD.n477 VDD.n476 185
R16706 VDD.n1827 VDD.n1826 185
R16707 VDD.n1829 VDD.n1828 185
R16708 VDD.n1831 VDD.n1824 185
R16709 VDD.n1834 VDD.n1833 185
R16710 VDD.n1835 VDD.n1823 185
R16711 VDD.n1837 VDD.n1836 185
R16712 VDD.n1839 VDD.n1822 185
R16713 VDD.n1842 VDD.n1841 185
R16714 VDD.n1843 VDD.n1821 185
R16715 VDD.n1845 VDD.n1844 185
R16716 VDD.n1847 VDD.n1820 185
R16717 VDD.n1850 VDD.n1849 185
R16718 VDD.n1851 VDD.n1819 185
R16719 VDD.n1853 VDD.n1852 185
R16720 VDD.n1855 VDD.n1818 185
R16721 VDD.n1858 VDD.n1857 185
R16722 VDD.n1859 VDD.n1817 185
R16723 VDD.n1861 VDD.n1860 185
R16724 VDD.n1863 VDD.n1816 185
R16725 VDD.n1866 VDD.n1865 185
R16726 VDD.n1867 VDD.n1811 185
R16727 VDD.n2396 VDD.n2395 185
R16728 VDD.n282 VDD.n280 185
R16729 VDD.n2283 VDD.n2282 185
R16730 VDD.n2285 VDD.n2284 185
R16731 VDD.n2287 VDD.n2286 185
R16732 VDD.n2289 VDD.n2288 185
R16733 VDD.n2291 VDD.n2290 185
R16734 VDD.n2293 VDD.n2292 185
R16735 VDD.n2295 VDD.n2294 185
R16736 VDD.n2297 VDD.n2296 185
R16737 VDD.n2299 VDD.n2298 185
R16738 VDD.n2301 VDD.n2300 185
R16739 VDD.n2303 VDD.n2302 185
R16740 VDD.n2305 VDD.n2304 185
R16741 VDD.n2307 VDD.n2306 185
R16742 VDD.n2309 VDD.n2308 185
R16743 VDD.n2311 VDD.n2310 185
R16744 VDD.n2313 VDD.n2312 185
R16745 VDD.n2315 VDD.n2314 185
R16746 VDD.n2317 VDD.n2316 185
R16747 VDD.n2319 VDD.n2318 185
R16748 VDD.n2321 VDD.n2320 185
R16749 VDD.n2394 VDD.n281 185
R16750 VDD.n287 VDD.n281 185
R16751 VDD.n2393 VDD.n2392 185
R16752 VDD.n2392 VDD.n2391 185
R16753 VDD.n284 VDD.n283 185
R16754 VDD.n285 VDD.n284 185
R16755 VDD.n1868 VDD.n298 185
R16756 VDD.n2337 VDD.n298 185
R16757 VDD.n1870 VDD.n1869 185
R16758 VDD.n1869 VDD.n297 185
R16759 VDD.n1871 VDD.n305 185
R16760 VDD.n2331 VDD.n305 185
R16761 VDD.n1873 VDD.n1872 185
R16762 VDD.n1872 VDD.n303 185
R16763 VDD.n1874 VDD.n312 185
R16764 VDD.n2275 VDD.n312 185
R16765 VDD.n1876 VDD.n1875 185
R16766 VDD.n1875 VDD.n310 185
R16767 VDD.n1877 VDD.n317 185
R16768 VDD.n2269 VDD.n317 185
R16769 VDD.n1879 VDD.n1878 185
R16770 VDD.n1878 VDD.n324 185
R16771 VDD.n1880 VDD.n323 185
R16772 VDD.n2263 VDD.n323 185
R16773 VDD.n1882 VDD.n1881 185
R16774 VDD.n1881 VDD.n321 185
R16775 VDD.n1883 VDD.n330 185
R16776 VDD.n2257 VDD.n330 185
R16777 VDD.n1885 VDD.n1884 185
R16778 VDD.n1884 VDD.n328 185
R16779 VDD.n1886 VDD.n336 185
R16780 VDD.n2251 VDD.n336 185
R16781 VDD.n1888 VDD.n1887 185
R16782 VDD.n1887 VDD.n334 185
R16783 VDD.n1889 VDD.n342 185
R16784 VDD.n2245 VDD.n342 185
R16785 VDD.n1891 VDD.n1890 185
R16786 VDD.n1890 VDD.n340 185
R16787 VDD.n1892 VDD.n348 185
R16788 VDD.n2239 VDD.n348 185
R16789 VDD.n1894 VDD.n1893 185
R16790 VDD.n1893 VDD.n346 185
R16791 VDD.n1895 VDD.n354 185
R16792 VDD.n2233 VDD.n354 185
R16793 VDD.n1897 VDD.n1896 185
R16794 VDD.n1896 VDD.n352 185
R16795 VDD.n1898 VDD.n360 185
R16796 VDD.n2227 VDD.n360 185
R16797 VDD.n1900 VDD.n1899 185
R16798 VDD.n1899 VDD.n358 185
R16799 VDD.n1901 VDD.n365 185
R16800 VDD.n2221 VDD.n365 185
R16801 VDD.n1903 VDD.n1902 185
R16802 VDD.n1902 VDD.n372 185
R16803 VDD.n1904 VDD.n371 185
R16804 VDD.n2215 VDD.n371 185
R16805 VDD.n1906 VDD.n1905 185
R16806 VDD.n1905 VDD.n369 185
R16807 VDD.n1907 VDD.n378 185
R16808 VDD.n2209 VDD.n378 185
R16809 VDD.n1909 VDD.n1908 185
R16810 VDD.n1908 VDD.n376 185
R16811 VDD.n1910 VDD.n383 185
R16812 VDD.n2203 VDD.n383 185
R16813 VDD.n1912 VDD.n1911 185
R16814 VDD.n1911 VDD.n390 185
R16815 VDD.n1913 VDD.n389 185
R16816 VDD.n2197 VDD.n389 185
R16817 VDD.n1915 VDD.n1914 185
R16818 VDD.n1914 VDD.n387 185
R16819 VDD.n1916 VDD.n396 185
R16820 VDD.n2191 VDD.n396 185
R16821 VDD.n1918 VDD.n1917 185
R16822 VDD.n1917 VDD.n394 185
R16823 VDD.n1919 VDD.n402 185
R16824 VDD.n2185 VDD.n402 185
R16825 VDD.n1921 VDD.n1920 185
R16826 VDD.n1920 VDD.n400 185
R16827 VDD.n1922 VDD.n408 185
R16828 VDD.n2179 VDD.n408 185
R16829 VDD.n1924 VDD.n1923 185
R16830 VDD.n1923 VDD.n406 185
R16831 VDD.n1925 VDD.n414 185
R16832 VDD.n2173 VDD.n414 185
R16833 VDD.n1927 VDD.n1926 185
R16834 VDD.n1926 VDD.n412 185
R16835 VDD.n1928 VDD.n420 185
R16836 VDD.n2167 VDD.n420 185
R16837 VDD.n1930 VDD.n1929 185
R16838 VDD.n1929 VDD.n418 185
R16839 VDD.n1931 VDD.n426 185
R16840 VDD.n2161 VDD.n426 185
R16841 VDD.n1933 VDD.n1932 185
R16842 VDD.n1932 VDD.n424 185
R16843 VDD.n1934 VDD.n431 185
R16844 VDD.n2155 VDD.n431 185
R16845 VDD.n1936 VDD.n1935 185
R16846 VDD.n1935 VDD.n438 185
R16847 VDD.n1937 VDD.n437 185
R16848 VDD.n2149 VDD.n437 185
R16849 VDD.n1939 VDD.n1938 185
R16850 VDD.n1938 VDD.n435 185
R16851 VDD.n1940 VDD.n444 185
R16852 VDD.n2143 VDD.n444 185
R16853 VDD.n1942 VDD.n1941 185
R16854 VDD.n1941 VDD.n442 185
R16855 VDD.n1943 VDD.n450 185
R16856 VDD.n2137 VDD.n450 185
R16857 VDD.n1945 VDD.n1944 185
R16858 VDD.n1944 VDD.n448 185
R16859 VDD.n1946 VDD.n456 185
R16860 VDD.n2131 VDD.n456 185
R16861 VDD.n1948 VDD.n1947 185
R16862 VDD.n1947 VDD.n454 185
R16863 VDD.n1949 VDD.n462 185
R16864 VDD.n2125 VDD.n462 185
R16865 VDD.n1951 VDD.n1950 185
R16866 VDD.n1950 VDD.n460 185
R16867 VDD.n1952 VDD.n468 185
R16868 VDD.n2119 VDD.n468 185
R16869 VDD.n1954 VDD.n1953 185
R16870 VDD.n1953 VDD.n466 185
R16871 VDD.n1955 VDD.n474 185
R16872 VDD.n2113 VDD.n474 185
R16873 VDD.n1956 VDD.n1812 185
R16874 VDD.n1812 VDD.n472 185
R16875 VDD.n1958 VDD.n1957 185
R16876 VDD.n2107 VDD.n1958 185
R16877 VDD.n1798 VDD.n509 185
R16878 VDD.n509 VDD.n478 185
R16879 VDD.n1800 VDD.n1799 185
R16880 VDD.n1801 VDD.n1800 185
R16881 VDD.n510 VDD.n508 185
R16882 VDD.n508 VDD.n505 185
R16883 VDD.n1746 VDD.n1745 185
R16884 VDD.n1747 VDD.n1746 185
R16885 VDD.n1744 VDD.n519 185
R16886 VDD.n519 VDD.n516 185
R16887 VDD.n1743 VDD.n1742 185
R16888 VDD.n1742 VDD.n1741 185
R16889 VDD.n521 VDD.n520 185
R16890 VDD.n522 VDD.n521 185
R16891 VDD.n1684 VDD.n1683 185
R16892 VDD.n1685 VDD.n1684 185
R16893 VDD.n1682 VDD.n532 185
R16894 VDD.n532 VDD.n529 185
R16895 VDD.n1681 VDD.n1680 185
R16896 VDD.n1680 VDD.n1679 185
R16897 VDD.n534 VDD.n533 185
R16898 VDD.n535 VDD.n534 185
R16899 VDD.n1672 VDD.n1671 185
R16900 VDD.n1673 VDD.n1672 185
R16901 VDD.n1670 VDD.n544 185
R16902 VDD.n544 VDD.n541 185
R16903 VDD.n1669 VDD.n1668 185
R16904 VDD.n1668 VDD.n1667 185
R16905 VDD.n546 VDD.n545 185
R16906 VDD.n547 VDD.n546 185
R16907 VDD.n1660 VDD.n1659 185
R16908 VDD.n1661 VDD.n1660 185
R16909 VDD.n1658 VDD.n555 185
R16910 VDD.n561 VDD.n555 185
R16911 VDD.n1657 VDD.n1656 185
R16912 VDD.n1656 VDD.n1655 185
R16913 VDD.n557 VDD.n556 185
R16914 VDD.n558 VDD.n557 185
R16915 VDD.n1648 VDD.n1647 185
R16916 VDD.n1649 VDD.n1648 185
R16917 VDD.n1646 VDD.n568 185
R16918 VDD.n568 VDD.n565 185
R16919 VDD.n1645 VDD.n1644 185
R16920 VDD.n1644 VDD.n1643 185
R16921 VDD.n570 VDD.n569 185
R16922 VDD.n571 VDD.n570 185
R16923 VDD.n1636 VDD.n1635 185
R16924 VDD.n1637 VDD.n1636 185
R16925 VDD.n1634 VDD.n580 185
R16926 VDD.n580 VDD.n577 185
R16927 VDD.n1633 VDD.n1632 185
R16928 VDD.n1632 VDD.n1631 185
R16929 VDD.n582 VDD.n581 185
R16930 VDD.n583 VDD.n582 185
R16931 VDD.n1624 VDD.n1623 185
R16932 VDD.n1625 VDD.n1624 185
R16933 VDD.n1622 VDD.n592 185
R16934 VDD.n592 VDD.n589 185
R16935 VDD.n1621 VDD.n1620 185
R16936 VDD.n1620 VDD.n1619 185
R16937 VDD.n594 VDD.n593 185
R16938 VDD.n595 VDD.n594 185
R16939 VDD.n1612 VDD.n1611 185
R16940 VDD.n1613 VDD.n1612 185
R16941 VDD.n1610 VDD.n603 185
R16942 VDD.n609 VDD.n603 185
R16943 VDD.n1609 VDD.n1608 185
R16944 VDD.n1608 VDD.n1607 185
R16945 VDD.n605 VDD.n604 185
R16946 VDD.n606 VDD.n605 185
R16947 VDD.n1600 VDD.n1599 185
R16948 VDD.n1601 VDD.n1600 185
R16949 VDD.n1598 VDD.n616 185
R16950 VDD.n616 VDD.n613 185
R16951 VDD.n1597 VDD.n1596 185
R16952 VDD.n1596 VDD.n1595 185
R16953 VDD.n618 VDD.n617 185
R16954 VDD.n627 VDD.n618 185
R16955 VDD.n1588 VDD.n1587 185
R16956 VDD.n1589 VDD.n1588 185
R16957 VDD.n1586 VDD.n628 185
R16958 VDD.n628 VDD.n624 185
R16959 VDD.n1585 VDD.n1584 185
R16960 VDD.n1584 VDD.n1583 185
R16961 VDD.n630 VDD.n629 185
R16962 VDD.n631 VDD.n630 185
R16963 VDD.n1576 VDD.n1575 185
R16964 VDD.n1577 VDD.n1576 185
R16965 VDD.n1574 VDD.n640 185
R16966 VDD.n640 VDD.n637 185
R16967 VDD.n1573 VDD.n1572 185
R16968 VDD.n1572 VDD.n1571 185
R16969 VDD.n642 VDD.n641 185
R16970 VDD.n643 VDD.n642 185
R16971 VDD.n1564 VDD.n1563 185
R16972 VDD.n1565 VDD.n1564 185
R16973 VDD.n1562 VDD.n652 185
R16974 VDD.n652 VDD.n649 185
R16975 VDD.n1561 VDD.n1560 185
R16976 VDD.n1560 VDD.n1559 185
R16977 VDD.n654 VDD.n653 185
R16978 VDD.n655 VDD.n654 185
R16979 VDD.n1552 VDD.n1551 185
R16980 VDD.n1553 VDD.n1552 185
R16981 VDD.n1550 VDD.n664 185
R16982 VDD.n664 VDD.n661 185
R16983 VDD.n1549 VDD.n1548 185
R16984 VDD.n1548 VDD.n1547 185
R16985 VDD.n666 VDD.n665 185
R16986 VDD.n675 VDD.n666 185
R16987 VDD.n1540 VDD.n1539 185
R16988 VDD.n1541 VDD.n1540 185
R16989 VDD.n1538 VDD.n676 185
R16990 VDD.n676 VDD.n672 185
R16991 VDD.n1537 VDD.n1536 185
R16992 VDD.n1536 VDD.n1535 185
R16993 VDD.n678 VDD.n677 185
R16994 VDD.n679 VDD.n678 185
R16995 VDD.n1528 VDD.n1527 185
R16996 VDD.n1529 VDD.n1528 185
R16997 VDD.n1526 VDD.n688 185
R16998 VDD.n688 VDD.n685 185
R16999 VDD.n1525 VDD.n1524 185
R17000 VDD.n1524 VDD.n1523 185
R17001 VDD.n690 VDD.n689 185
R17002 VDD.n691 VDD.n690 185
R17003 VDD.n1516 VDD.n1515 185
R17004 VDD.n1517 VDD.n1516 185
R17005 VDD.n1514 VDD.n699 185
R17006 VDD.n1513 VDD.n1512 185
R17007 VDD.n701 VDD.n700 185
R17008 VDD.n1510 VDD.n701 185
R17009 VDD.n1237 VDD.n1236 185
R17010 VDD.n1239 VDD.n1238 185
R17011 VDD.n1241 VDD.n1240 185
R17012 VDD.n1243 VDD.n1242 185
R17013 VDD.n1245 VDD.n1244 185
R17014 VDD.n1247 VDD.n1246 185
R17015 VDD.n1249 VDD.n1248 185
R17016 VDD.n1251 VDD.n1250 185
R17017 VDD.n1253 VDD.n1252 185
R17018 VDD.n1255 VDD.n1254 185
R17019 VDD.n1257 VDD.n1256 185
R17020 VDD.n1259 VDD.n1258 185
R17021 VDD.n1261 VDD.n1260 185
R17022 VDD.n1263 VDD.n1262 185
R17023 VDD.n1265 VDD.n1264 185
R17024 VDD.n1267 VDD.n1266 185
R17025 VDD.n1269 VDD.n1268 185
R17026 VDD.n1271 VDD.n1233 185
R17027 VDD.n1362 VDD.n1361 185
R17028 VDD.n1510 VDD.n1362 185
R17029 VDD.n1755 VDD.n1754 185
R17030 VDD.n1757 VDD.n1756 185
R17031 VDD.n1759 VDD.n1758 185
R17032 VDD.n1761 VDD.n1760 185
R17033 VDD.n1763 VDD.n1762 185
R17034 VDD.n1765 VDD.n1764 185
R17035 VDD.n1767 VDD.n1766 185
R17036 VDD.n1769 VDD.n1768 185
R17037 VDD.n1771 VDD.n1770 185
R17038 VDD.n1773 VDD.n1772 185
R17039 VDD.n1775 VDD.n1774 185
R17040 VDD.n1777 VDD.n1776 185
R17041 VDD.n1779 VDD.n1778 185
R17042 VDD.n1781 VDD.n1780 185
R17043 VDD.n1783 VDD.n1782 185
R17044 VDD.n1785 VDD.n1784 185
R17045 VDD.n1787 VDD.n1786 185
R17046 VDD.n1789 VDD.n1788 185
R17047 VDD.n1791 VDD.n1790 185
R17048 VDD.n1793 VDD.n1792 185
R17049 VDD.n1795 VDD.n1794 185
R17050 VDD.n1797 VDD.n1796 185
R17051 VDD.n1753 VDD.n1752 185
R17052 VDD.n1753 VDD.n478 185
R17053 VDD.n1751 VDD.n506 185
R17054 VDD.n1801 VDD.n506 185
R17055 VDD.n1750 VDD.n1749 185
R17056 VDD.n1749 VDD.n505 185
R17057 VDD.n1748 VDD.n514 185
R17058 VDD.n1748 VDD.n1747 185
R17059 VDD.n1272 VDD.n515 185
R17060 VDD.n516 VDD.n515 185
R17061 VDD.n1273 VDD.n523 185
R17062 VDD.n1741 VDD.n523 185
R17063 VDD.n1275 VDD.n1274 185
R17064 VDD.n1274 VDD.n522 185
R17065 VDD.n1276 VDD.n530 185
R17066 VDD.n1685 VDD.n530 185
R17067 VDD.n1278 VDD.n1277 185
R17068 VDD.n1277 VDD.n529 185
R17069 VDD.n1279 VDD.n536 185
R17070 VDD.n1679 VDD.n536 185
R17071 VDD.n1281 VDD.n1280 185
R17072 VDD.n1280 VDD.n535 185
R17073 VDD.n1282 VDD.n542 185
R17074 VDD.n1673 VDD.n542 185
R17075 VDD.n1284 VDD.n1283 185
R17076 VDD.n1283 VDD.n541 185
R17077 VDD.n1285 VDD.n548 185
R17078 VDD.n1667 VDD.n548 185
R17079 VDD.n1287 VDD.n1286 185
R17080 VDD.n1286 VDD.n547 185
R17081 VDD.n1288 VDD.n553 185
R17082 VDD.n1661 VDD.n553 185
R17083 VDD.n1290 VDD.n1289 185
R17084 VDD.n1289 VDD.n561 185
R17085 VDD.n1291 VDD.n559 185
R17086 VDD.n1655 VDD.n559 185
R17087 VDD.n1293 VDD.n1292 185
R17088 VDD.n1292 VDD.n558 185
R17089 VDD.n1294 VDD.n566 185
R17090 VDD.n1649 VDD.n566 185
R17091 VDD.n1296 VDD.n1295 185
R17092 VDD.n1295 VDD.n565 185
R17093 VDD.n1297 VDD.n572 185
R17094 VDD.n1643 VDD.n572 185
R17095 VDD.n1299 VDD.n1298 185
R17096 VDD.n1298 VDD.n571 185
R17097 VDD.n1300 VDD.n578 185
R17098 VDD.n1637 VDD.n578 185
R17099 VDD.n1302 VDD.n1301 185
R17100 VDD.n1301 VDD.n577 185
R17101 VDD.n1303 VDD.n584 185
R17102 VDD.n1631 VDD.n584 185
R17103 VDD.n1305 VDD.n1304 185
R17104 VDD.n1304 VDD.n583 185
R17105 VDD.n1306 VDD.n590 185
R17106 VDD.n1625 VDD.n590 185
R17107 VDD.n1308 VDD.n1307 185
R17108 VDD.n1307 VDD.n589 185
R17109 VDD.n1309 VDD.n596 185
R17110 VDD.n1619 VDD.n596 185
R17111 VDD.n1311 VDD.n1310 185
R17112 VDD.n1310 VDD.n595 185
R17113 VDD.n1312 VDD.n601 185
R17114 VDD.n1613 VDD.n601 185
R17115 VDD.n1314 VDD.n1313 185
R17116 VDD.n1313 VDD.n609 185
R17117 VDD.n1315 VDD.n607 185
R17118 VDD.n1607 VDD.n607 185
R17119 VDD.n1317 VDD.n1316 185
R17120 VDD.n1316 VDD.n606 185
R17121 VDD.n1318 VDD.n614 185
R17122 VDD.n1601 VDD.n614 185
R17123 VDD.n1320 VDD.n1319 185
R17124 VDD.n1319 VDD.n613 185
R17125 VDD.n1321 VDD.n619 185
R17126 VDD.n1595 VDD.n619 185
R17127 VDD.n1323 VDD.n1322 185
R17128 VDD.n1322 VDD.n627 185
R17129 VDD.n1324 VDD.n625 185
R17130 VDD.n1589 VDD.n625 185
R17131 VDD.n1326 VDD.n1325 185
R17132 VDD.n1325 VDD.n624 185
R17133 VDD.n1327 VDD.n632 185
R17134 VDD.n1583 VDD.n632 185
R17135 VDD.n1329 VDD.n1328 185
R17136 VDD.n1328 VDD.n631 185
R17137 VDD.n1330 VDD.n638 185
R17138 VDD.n1577 VDD.n638 185
R17139 VDD.n1332 VDD.n1331 185
R17140 VDD.n1331 VDD.n637 185
R17141 VDD.n1333 VDD.n644 185
R17142 VDD.n1571 VDD.n644 185
R17143 VDD.n1335 VDD.n1334 185
R17144 VDD.n1334 VDD.n643 185
R17145 VDD.n1336 VDD.n650 185
R17146 VDD.n1565 VDD.n650 185
R17147 VDD.n1338 VDD.n1337 185
R17148 VDD.n1337 VDD.n649 185
R17149 VDD.n1339 VDD.n656 185
R17150 VDD.n1559 VDD.n656 185
R17151 VDD.n1341 VDD.n1340 185
R17152 VDD.n1340 VDD.n655 185
R17153 VDD.n1342 VDD.n662 185
R17154 VDD.n1553 VDD.n662 185
R17155 VDD.n1344 VDD.n1343 185
R17156 VDD.n1343 VDD.n661 185
R17157 VDD.n1345 VDD.n667 185
R17158 VDD.n1547 VDD.n667 185
R17159 VDD.n1347 VDD.n1346 185
R17160 VDD.n1346 VDD.n675 185
R17161 VDD.n1348 VDD.n673 185
R17162 VDD.n1541 VDD.n673 185
R17163 VDD.n1350 VDD.n1349 185
R17164 VDD.n1349 VDD.n672 185
R17165 VDD.n1351 VDD.n680 185
R17166 VDD.n1535 VDD.n680 185
R17167 VDD.n1353 VDD.n1352 185
R17168 VDD.n1352 VDD.n679 185
R17169 VDD.n1354 VDD.n686 185
R17170 VDD.n1529 VDD.n686 185
R17171 VDD.n1356 VDD.n1355 185
R17172 VDD.n1355 VDD.n685 185
R17173 VDD.n1357 VDD.n692 185
R17174 VDD.n1523 VDD.n692 185
R17175 VDD.n1359 VDD.n1358 185
R17176 VDD.n1358 VDD.n691 185
R17177 VDD.n1360 VDD.n697 185
R17178 VDD.n1517 VDD.n697 185
R17179 VDD.n2626 VDD.n2625 185
R17180 VDD.n2625 VDD.n2624 185
R17181 VDD.n2627 VDD.n85 185
R17182 VDD.n85 VDD.n84 185
R17183 VDD.n2629 VDD.n2628 185
R17184 VDD.n2630 VDD.n2629 185
R17185 VDD.n80 VDD.n79 185
R17186 VDD.n2631 VDD.n80 185
R17187 VDD.n2634 VDD.n2633 185
R17188 VDD.n2633 VDD.n2632 185
R17189 VDD.n2635 VDD.n74 185
R17190 VDD.n74 VDD.n73 185
R17191 VDD.n2637 VDD.n2636 185
R17192 VDD.n2638 VDD.n2637 185
R17193 VDD.n69 VDD.n68 185
R17194 VDD.n2639 VDD.n69 185
R17195 VDD.n2642 VDD.n2641 185
R17196 VDD.n2641 VDD.n2640 185
R17197 VDD.n2643 VDD.n63 185
R17198 VDD.n63 VDD.n62 185
R17199 VDD.n2645 VDD.n2644 185
R17200 VDD.n2646 VDD.n2645 185
R17201 VDD.n58 VDD.n57 185
R17202 VDD.n2647 VDD.n58 185
R17203 VDD.n2650 VDD.n2649 185
R17204 VDD.n2649 VDD.n2648 185
R17205 VDD.n2651 VDD.n52 185
R17206 VDD.n52 VDD.n51 185
R17207 VDD.n2653 VDD.n2652 185
R17208 VDD.n2654 VDD.n2653 185
R17209 VDD.n47 VDD.n46 185
R17210 VDD.n2655 VDD.n47 185
R17211 VDD.n2658 VDD.n2657 185
R17212 VDD.n2657 VDD.n2656 185
R17213 VDD.n2659 VDD.n41 185
R17214 VDD.n41 VDD.n40 185
R17215 VDD.n2661 VDD.n2660 185
R17216 VDD.n2662 VDD.n2661 185
R17217 VDD.n36 VDD.n35 185
R17218 VDD.n2663 VDD.n36 185
R17219 VDD.n2666 VDD.n2665 185
R17220 VDD.n2665 VDD.n2664 185
R17221 VDD.n2667 VDD.n31 185
R17222 VDD.n31 VDD.n30 185
R17223 VDD.n2669 VDD.n2668 185
R17224 VDD.n2670 VDD.n2669 185
R17225 VDD.n26 VDD.n24 185
R17226 VDD.n2671 VDD.n26 185
R17227 VDD.n2674 VDD.n2673 185
R17228 VDD.n2673 VDD.n2672 185
R17229 VDD.n25 VDD.n23 185
R17230 VDD.n2572 VDD.n25 185
R17231 VDD.n2570 VDD.n2569 185
R17232 VDD.n2571 VDD.n2570 185
R17233 VDD.n186 VDD.n185 185
R17234 VDD.n185 VDD.n184 185
R17235 VDD.n2565 VDD.n2564 185
R17236 VDD.n2564 VDD.n2563 185
R17237 VDD.n189 VDD.n188 185
R17238 VDD.n190 VDD.n189 185
R17239 VDD.n2551 VDD.n2550 185
R17240 VDD.n2552 VDD.n2551 185
R17241 VDD.n199 VDD.n198 185
R17242 VDD.n198 VDD.n197 185
R17243 VDD.n2546 VDD.n2545 185
R17244 VDD.n2545 VDD.n2544 185
R17245 VDD.n202 VDD.n201 185
R17246 VDD.n203 VDD.n202 185
R17247 VDD.n2535 VDD.n2534 185
R17248 VDD.n2536 VDD.n2535 185
R17249 VDD.n211 VDD.n210 185
R17250 VDD.n210 VDD.n209 185
R17251 VDD.n2530 VDD.n2529 185
R17252 VDD.n2529 VDD.n2528 185
R17253 VDD.n214 VDD.n213 185
R17254 VDD.n215 VDD.n214 185
R17255 VDD.n2519 VDD.n2518 185
R17256 VDD.n2520 VDD.n2519 185
R17257 VDD.n223 VDD.n222 185
R17258 VDD.n222 VDD.n221 185
R17259 VDD.n2514 VDD.n2513 185
R17260 VDD.n2513 VDD.n2512 185
R17261 VDD.n226 VDD.n225 185
R17262 VDD.n227 VDD.n226 185
R17263 VDD.n2503 VDD.n2502 185
R17264 VDD.n2504 VDD.n2503 185
R17265 VDD.n235 VDD.n234 185
R17266 VDD.n234 VDD.n233 185
R17267 VDD.n2498 VDD.n2497 185
R17268 VDD.n2497 VDD.n2496 185
R17269 VDD.n238 VDD.n237 185
R17270 VDD.n245 VDD.n238 185
R17271 VDD.n2487 VDD.n2486 185
R17272 VDD.n2488 VDD.n2487 185
R17273 VDD.n247 VDD.n246 185
R17274 VDD.n246 VDD.n244 185
R17275 VDD.n2482 VDD.n2481 185
R17276 VDD.n2481 VDD.n2480 185
R17277 VDD.n250 VDD.n249 185
R17278 VDD.n251 VDD.n250 185
R17279 VDD.n2470 VDD.n2469 185
R17280 VDD.n2468 VDD.n2409 185
R17281 VDD.n2467 VDD.n2408 185
R17282 VDD.n2472 VDD.n2408 185
R17283 VDD.n2466 VDD.n2465 185
R17284 VDD.n2464 VDD.n2463 185
R17285 VDD.n2462 VDD.n2461 185
R17286 VDD.n2460 VDD.n2459 185
R17287 VDD.n2458 VDD.n2457 185
R17288 VDD.n2456 VDD.n2455 185
R17289 VDD.n2454 VDD.n2453 185
R17290 VDD.n2452 VDD.n2451 185
R17291 VDD.n2450 VDD.n2449 185
R17292 VDD.n2448 VDD.n2447 185
R17293 VDD.n2446 VDD.n2445 185
R17294 VDD.n2444 VDD.n2443 185
R17295 VDD.n2442 VDD.n2441 185
R17296 VDD.n2440 VDD.n2439 185
R17297 VDD.n2438 VDD.n2437 185
R17298 VDD.n2436 VDD.n2435 185
R17299 VDD.n2434 VDD.n2433 185
R17300 VDD.n2432 VDD.n258 185
R17301 VDD.n2474 VDD.n2473 185
R17302 VDD.n2473 VDD.n2472 185
R17303 VDD.n2621 VDD.n2620 185
R17304 VDD.n167 VDD.n102 185
R17305 VDD.n166 VDD.n165 185
R17306 VDD.n164 VDD.n163 185
R17307 VDD.n162 VDD.n107 185
R17308 VDD.n158 VDD.n157 185
R17309 VDD.n156 VDD.n155 185
R17310 VDD.n154 VDD.n153 185
R17311 VDD.n152 VDD.n109 185
R17312 VDD.n148 VDD.n147 185
R17313 VDD.n146 VDD.n145 185
R17314 VDD.n144 VDD.n143 185
R17315 VDD.n142 VDD.n113 185
R17316 VDD.n138 VDD.n137 185
R17317 VDD.n136 VDD.n135 185
R17318 VDD.n134 VDD.n133 185
R17319 VDD.n132 VDD.n115 185
R17320 VDD.n128 VDD.n127 185
R17321 VDD.n126 VDD.n125 185
R17322 VDD.n124 VDD.n123 185
R17323 VDD.n122 VDD.n117 185
R17324 VDD.n118 VDD.n90 185
R17325 VDD.n2617 VDD.n91 185
R17326 VDD.n2624 VDD.n91 185
R17327 VDD.n2616 VDD.n2615 185
R17328 VDD.n2615 VDD.n84 185
R17329 VDD.n2614 VDD.n83 185
R17330 VDD.n2630 VDD.n83 185
R17331 VDD.n170 VDD.n82 185
R17332 VDD.n2631 VDD.n82 185
R17333 VDD.n2610 VDD.n81 185
R17334 VDD.n2632 VDD.n81 185
R17335 VDD.n2609 VDD.n2608 185
R17336 VDD.n2608 VDD.n73 185
R17337 VDD.n2607 VDD.n72 185
R17338 VDD.n2638 VDD.n72 185
R17339 VDD.n172 VDD.n71 185
R17340 VDD.n2639 VDD.n71 185
R17341 VDD.n2603 VDD.n70 185
R17342 VDD.n2640 VDD.n70 185
R17343 VDD.n2602 VDD.n2601 185
R17344 VDD.n2601 VDD.n62 185
R17345 VDD.n2600 VDD.n61 185
R17346 VDD.n2646 VDD.n61 185
R17347 VDD.n174 VDD.n60 185
R17348 VDD.n2647 VDD.n60 185
R17349 VDD.n2596 VDD.n59 185
R17350 VDD.n2648 VDD.n59 185
R17351 VDD.n2595 VDD.n2594 185
R17352 VDD.n2594 VDD.n51 185
R17353 VDD.n2593 VDD.n50 185
R17354 VDD.n2654 VDD.n50 185
R17355 VDD.n176 VDD.n49 185
R17356 VDD.n2655 VDD.n49 185
R17357 VDD.n2589 VDD.n48 185
R17358 VDD.n2656 VDD.n48 185
R17359 VDD.n2588 VDD.n2587 185
R17360 VDD.n2587 VDD.n40 185
R17361 VDD.n2586 VDD.n39 185
R17362 VDD.n2662 VDD.n39 185
R17363 VDD.n178 VDD.n38 185
R17364 VDD.n2663 VDD.n38 185
R17365 VDD.n2582 VDD.n37 185
R17366 VDD.n2664 VDD.n37 185
R17367 VDD.n2581 VDD.n2580 185
R17368 VDD.n2580 VDD.n30 185
R17369 VDD.n2579 VDD.n29 185
R17370 VDD.n2670 VDD.n29 185
R17371 VDD.n180 VDD.n28 185
R17372 VDD.n2671 VDD.n28 185
R17373 VDD.n2575 VDD.n27 185
R17374 VDD.n2672 VDD.n27 185
R17375 VDD.n2574 VDD.n2573 185
R17376 VDD.n2573 VDD.n2572 185
R17377 VDD.n183 VDD.n182 185
R17378 VDD.n2571 VDD.n183 185
R17379 VDD.n2560 VDD.n192 185
R17380 VDD.n192 VDD.n184 185
R17381 VDD.n2562 VDD.n2561 185
R17382 VDD.n2563 VDD.n2562 185
R17383 VDD.n193 VDD.n191 185
R17384 VDD.n191 VDD.n190 185
R17385 VDD.n2554 VDD.n2553 185
R17386 VDD.n2553 VDD.n2552 185
R17387 VDD.n196 VDD.n195 185
R17388 VDD.n197 VDD.n196 185
R17389 VDD.n2543 VDD.n2542 185
R17390 VDD.n2544 VDD.n2543 185
R17391 VDD.n205 VDD.n204 185
R17392 VDD.n204 VDD.n203 185
R17393 VDD.n2538 VDD.n2537 185
R17394 VDD.n2537 VDD.n2536 185
R17395 VDD.n208 VDD.n207 185
R17396 VDD.n209 VDD.n208 185
R17397 VDD.n2527 VDD.n2526 185
R17398 VDD.n2528 VDD.n2527 185
R17399 VDD.n217 VDD.n216 185
R17400 VDD.n216 VDD.n215 185
R17401 VDD.n2522 VDD.n2521 185
R17402 VDD.n2521 VDD.n2520 185
R17403 VDD.n220 VDD.n219 185
R17404 VDD.n221 VDD.n220 185
R17405 VDD.n2511 VDD.n2510 185
R17406 VDD.n2512 VDD.n2511 185
R17407 VDD.n229 VDD.n228 185
R17408 VDD.n228 VDD.n227 185
R17409 VDD.n2506 VDD.n2505 185
R17410 VDD.n2505 VDD.n2504 185
R17411 VDD.n232 VDD.n231 185
R17412 VDD.n233 VDD.n232 185
R17413 VDD.n2495 VDD.n2494 185
R17414 VDD.n2496 VDD.n2495 185
R17415 VDD.n240 VDD.n239 185
R17416 VDD.n245 VDD.n239 185
R17417 VDD.n2490 VDD.n2489 185
R17418 VDD.n2489 VDD.n2488 185
R17419 VDD.n243 VDD.n242 185
R17420 VDD.n244 VDD.n243 185
R17421 VDD.n2479 VDD.n2478 185
R17422 VDD.n2480 VDD.n2479 185
R17423 VDD.n253 VDD.n252 185
R17424 VDD.n252 VDD.n251 185
R17425 VDD.n2104 VDD.n1959 185
R17426 VDD.n2103 VDD.n2102 185
R17427 VDD.n2100 VDD.n1960 185
R17428 VDD.n2100 VDD.n1809 185
R17429 VDD.n2099 VDD.n2098 185
R17430 VDD.n2097 VDD.n2096 185
R17431 VDD.n2095 VDD.n1962 185
R17432 VDD.n2093 VDD.n2092 185
R17433 VDD.n2091 VDD.n1963 185
R17434 VDD.n2090 VDD.n2089 185
R17435 VDD.n2087 VDD.n1964 185
R17436 VDD.n2085 VDD.n2084 185
R17437 VDD.n2083 VDD.n1965 185
R17438 VDD.n2082 VDD.n2081 185
R17439 VDD.n2079 VDD.n1966 185
R17440 VDD.n2077 VDD.n2076 185
R17441 VDD.n2075 VDD.n1967 185
R17442 VDD.n2074 VDD.n2073 185
R17443 VDD.n2071 VDD.n1968 185
R17444 VDD.n2069 VDD.n2068 185
R17445 VDD.n2067 VDD.n1969 185
R17446 VDD.n2065 VDD.n2064 185
R17447 VDD.n2062 VDD.n2061 185
R17448 VDD.n2062 VDD.n1809 185
R17449 VDD.n2345 VDD.n2344 185
R17450 VDD.n2347 VDD.n2346 185
R17451 VDD.n2349 VDD.n2348 185
R17452 VDD.n2351 VDD.n2350 185
R17453 VDD.n2353 VDD.n2352 185
R17454 VDD.n2355 VDD.n2354 185
R17455 VDD.n2357 VDD.n2356 185
R17456 VDD.n2359 VDD.n2358 185
R17457 VDD.n2361 VDD.n2360 185
R17458 VDD.n2363 VDD.n2362 185
R17459 VDD.n2365 VDD.n2364 185
R17460 VDD.n2367 VDD.n2366 185
R17461 VDD.n2369 VDD.n2368 185
R17462 VDD.n2371 VDD.n2370 185
R17463 VDD.n2373 VDD.n2372 185
R17464 VDD.n2375 VDD.n2374 185
R17465 VDD.n2377 VDD.n2376 185
R17466 VDD.n2379 VDD.n2378 185
R17467 VDD.n2381 VDD.n2380 185
R17468 VDD.n2383 VDD.n2382 185
R17469 VDD.n2385 VDD.n2384 185
R17470 VDD.n2387 VDD.n2386 185
R17471 VDD.n2343 VDD.n2342 185
R17472 VDD.n2343 VDD.n287 185
R17473 VDD.n2341 VDD.n286 185
R17474 VDD.n2391 VDD.n286 185
R17475 VDD.n2340 VDD.n2339 185
R17476 VDD.n2339 VDD.n285 185
R17477 VDD.n2338 VDD.n295 185
R17478 VDD.n2338 VDD.n2337 185
R17479 VDD.n1972 VDD.n296 185
R17480 VDD.n297 VDD.n296 185
R17481 VDD.n1973 VDD.n304 185
R17482 VDD.n2331 VDD.n304 185
R17483 VDD.n1975 VDD.n1974 185
R17484 VDD.n1974 VDD.n303 185
R17485 VDD.n1976 VDD.n311 185
R17486 VDD.n2275 VDD.n311 185
R17487 VDD.n1978 VDD.n1977 185
R17488 VDD.n1977 VDD.n310 185
R17489 VDD.n1979 VDD.n316 185
R17490 VDD.n2269 VDD.n316 185
R17491 VDD.n1981 VDD.n1980 185
R17492 VDD.n1980 VDD.n324 185
R17493 VDD.n1982 VDD.n322 185
R17494 VDD.n2263 VDD.n322 185
R17495 VDD.n1984 VDD.n1983 185
R17496 VDD.n1983 VDD.n321 185
R17497 VDD.n1985 VDD.n329 185
R17498 VDD.n2257 VDD.n329 185
R17499 VDD.n1987 VDD.n1986 185
R17500 VDD.n1986 VDD.n328 185
R17501 VDD.n1988 VDD.n335 185
R17502 VDD.n2251 VDD.n335 185
R17503 VDD.n1990 VDD.n1989 185
R17504 VDD.n1989 VDD.n334 185
R17505 VDD.n1991 VDD.n341 185
R17506 VDD.n2245 VDD.n341 185
R17507 VDD.n1993 VDD.n1992 185
R17508 VDD.n1992 VDD.n340 185
R17509 VDD.n1994 VDD.n347 185
R17510 VDD.n2239 VDD.n347 185
R17511 VDD.n1996 VDD.n1995 185
R17512 VDD.n1995 VDD.n346 185
R17513 VDD.n1997 VDD.n353 185
R17514 VDD.n2233 VDD.n353 185
R17515 VDD.n1999 VDD.n1998 185
R17516 VDD.n1998 VDD.n352 185
R17517 VDD.n2000 VDD.n359 185
R17518 VDD.n2227 VDD.n359 185
R17519 VDD.n2002 VDD.n2001 185
R17520 VDD.n2001 VDD.n358 185
R17521 VDD.n2003 VDD.n364 185
R17522 VDD.n2221 VDD.n364 185
R17523 VDD.n2005 VDD.n2004 185
R17524 VDD.n2004 VDD.n372 185
R17525 VDD.n2006 VDD.n370 185
R17526 VDD.n2215 VDD.n370 185
R17527 VDD.n2008 VDD.n2007 185
R17528 VDD.n2007 VDD.n369 185
R17529 VDD.n2009 VDD.n377 185
R17530 VDD.n2209 VDD.n377 185
R17531 VDD.n2011 VDD.n2010 185
R17532 VDD.n2010 VDD.n376 185
R17533 VDD.n2012 VDD.n382 185
R17534 VDD.n2203 VDD.n382 185
R17535 VDD.n2014 VDD.n2013 185
R17536 VDD.n2013 VDD.n390 185
R17537 VDD.n2015 VDD.n388 185
R17538 VDD.n2197 VDD.n388 185
R17539 VDD.n2017 VDD.n2016 185
R17540 VDD.n2016 VDD.n387 185
R17541 VDD.n2018 VDD.n395 185
R17542 VDD.n2191 VDD.n395 185
R17543 VDD.n2020 VDD.n2019 185
R17544 VDD.n2019 VDD.n394 185
R17545 VDD.n2021 VDD.n401 185
R17546 VDD.n2185 VDD.n401 185
R17547 VDD.n2023 VDD.n2022 185
R17548 VDD.n2022 VDD.n400 185
R17549 VDD.n2024 VDD.n407 185
R17550 VDD.n2179 VDD.n407 185
R17551 VDD.n2026 VDD.n2025 185
R17552 VDD.n2025 VDD.n406 185
R17553 VDD.n2027 VDD.n413 185
R17554 VDD.n2173 VDD.n413 185
R17555 VDD.n2029 VDD.n2028 185
R17556 VDD.n2028 VDD.n412 185
R17557 VDD.n2030 VDD.n419 185
R17558 VDD.n2167 VDD.n419 185
R17559 VDD.n2032 VDD.n2031 185
R17560 VDD.n2031 VDD.n418 185
R17561 VDD.n2033 VDD.n425 185
R17562 VDD.n2161 VDD.n425 185
R17563 VDD.n2035 VDD.n2034 185
R17564 VDD.n2034 VDD.n424 185
R17565 VDD.n2036 VDD.n430 185
R17566 VDD.n2155 VDD.n430 185
R17567 VDD.n2038 VDD.n2037 185
R17568 VDD.n2037 VDD.n438 185
R17569 VDD.n2039 VDD.n436 185
R17570 VDD.n2149 VDD.n436 185
R17571 VDD.n2041 VDD.n2040 185
R17572 VDD.n2040 VDD.n435 185
R17573 VDD.n2042 VDD.n443 185
R17574 VDD.n2143 VDD.n443 185
R17575 VDD.n2044 VDD.n2043 185
R17576 VDD.n2043 VDD.n442 185
R17577 VDD.n2045 VDD.n449 185
R17578 VDD.n2137 VDD.n449 185
R17579 VDD.n2047 VDD.n2046 185
R17580 VDD.n2046 VDD.n448 185
R17581 VDD.n2048 VDD.n455 185
R17582 VDD.n2131 VDD.n455 185
R17583 VDD.n2050 VDD.n2049 185
R17584 VDD.n2049 VDD.n454 185
R17585 VDD.n2051 VDD.n461 185
R17586 VDD.n2125 VDD.n461 185
R17587 VDD.n2053 VDD.n2052 185
R17588 VDD.n2052 VDD.n460 185
R17589 VDD.n2054 VDD.n467 185
R17590 VDD.n2119 VDD.n467 185
R17591 VDD.n2056 VDD.n2055 185
R17592 VDD.n2055 VDD.n466 185
R17593 VDD.n2057 VDD.n473 185
R17594 VDD.n2113 VDD.n473 185
R17595 VDD.n2059 VDD.n2058 185
R17596 VDD.n2058 VDD.n472 185
R17597 VDD.n2060 VDD.n1810 185
R17598 VDD.n2107 VDD.n1810 185
R17599 VDD.n2106 VDD.n2105 185
R17600 VDD.n2107 VDD.n2106 185
R17601 VDD.n471 VDD.n470 185
R17602 VDD.n472 VDD.n471 185
R17603 VDD.n2115 VDD.n2114 185
R17604 VDD.n2114 VDD.n2113 185
R17605 VDD.n2116 VDD.n469 185
R17606 VDD.n469 VDD.n466 185
R17607 VDD.n2118 VDD.n2117 185
R17608 VDD.n2119 VDD.n2118 185
R17609 VDD.n459 VDD.n458 185
R17610 VDD.n460 VDD.n459 185
R17611 VDD.n2127 VDD.n2126 185
R17612 VDD.n2126 VDD.n2125 185
R17613 VDD.n2128 VDD.n457 185
R17614 VDD.n457 VDD.n454 185
R17615 VDD.n2130 VDD.n2129 185
R17616 VDD.n2131 VDD.n2130 185
R17617 VDD.n447 VDD.n446 185
R17618 VDD.n448 VDD.n447 185
R17619 VDD.n2139 VDD.n2138 185
R17620 VDD.n2138 VDD.n2137 185
R17621 VDD.n2140 VDD.n445 185
R17622 VDD.n445 VDD.n442 185
R17623 VDD.n2142 VDD.n2141 185
R17624 VDD.n2143 VDD.n2142 185
R17625 VDD.n434 VDD.n433 185
R17626 VDD.n435 VDD.n434 185
R17627 VDD.n2151 VDD.n2150 185
R17628 VDD.n2150 VDD.n2149 185
R17629 VDD.n2152 VDD.n432 185
R17630 VDD.n438 VDD.n432 185
R17631 VDD.n2154 VDD.n2153 185
R17632 VDD.n2155 VDD.n2154 185
R17633 VDD.n423 VDD.n422 185
R17634 VDD.n424 VDD.n423 185
R17635 VDD.n2163 VDD.n2162 185
R17636 VDD.n2162 VDD.n2161 185
R17637 VDD.n2164 VDD.n421 185
R17638 VDD.n421 VDD.n418 185
R17639 VDD.n2166 VDD.n2165 185
R17640 VDD.n2167 VDD.n2166 185
R17641 VDD.n411 VDD.n410 185
R17642 VDD.n412 VDD.n411 185
R17643 VDD.n2175 VDD.n2174 185
R17644 VDD.n2174 VDD.n2173 185
R17645 VDD.n2176 VDD.n409 185
R17646 VDD.n409 VDD.n406 185
R17647 VDD.n2178 VDD.n2177 185
R17648 VDD.n2179 VDD.n2178 185
R17649 VDD.n399 VDD.n398 185
R17650 VDD.n400 VDD.n399 185
R17651 VDD.n2187 VDD.n2186 185
R17652 VDD.n2186 VDD.n2185 185
R17653 VDD.n2188 VDD.n397 185
R17654 VDD.n397 VDD.n394 185
R17655 VDD.n2190 VDD.n2189 185
R17656 VDD.n2191 VDD.n2190 185
R17657 VDD.n386 VDD.n385 185
R17658 VDD.n387 VDD.n386 185
R17659 VDD.n2199 VDD.n2198 185
R17660 VDD.n2198 VDD.n2197 185
R17661 VDD.n2200 VDD.n384 185
R17662 VDD.n390 VDD.n384 185
R17663 VDD.n2202 VDD.n2201 185
R17664 VDD.n2203 VDD.n2202 185
R17665 VDD.n375 VDD.n374 185
R17666 VDD.n376 VDD.n375 185
R17667 VDD.n2211 VDD.n2210 185
R17668 VDD.n2210 VDD.n2209 185
R17669 VDD.n2212 VDD.n373 185
R17670 VDD.n373 VDD.n369 185
R17671 VDD.n2214 VDD.n2213 185
R17672 VDD.n2215 VDD.n2214 185
R17673 VDD.n363 VDD.n362 185
R17674 VDD.n372 VDD.n363 185
R17675 VDD.n2223 VDD.n2222 185
R17676 VDD.n2222 VDD.n2221 185
R17677 VDD.n2224 VDD.n361 185
R17678 VDD.n361 VDD.n358 185
R17679 VDD.n2226 VDD.n2225 185
R17680 VDD.n2227 VDD.n2226 185
R17681 VDD.n351 VDD.n350 185
R17682 VDD.n352 VDD.n351 185
R17683 VDD.n2235 VDD.n2234 185
R17684 VDD.n2234 VDD.n2233 185
R17685 VDD.n2236 VDD.n349 185
R17686 VDD.n349 VDD.n346 185
R17687 VDD.n2238 VDD.n2237 185
R17688 VDD.n2239 VDD.n2238 185
R17689 VDD.n339 VDD.n338 185
R17690 VDD.n340 VDD.n339 185
R17691 VDD.n2247 VDD.n2246 185
R17692 VDD.n2246 VDD.n2245 185
R17693 VDD.n2248 VDD.n337 185
R17694 VDD.n337 VDD.n334 185
R17695 VDD.n2250 VDD.n2249 185
R17696 VDD.n2251 VDD.n2250 185
R17697 VDD.n327 VDD.n326 185
R17698 VDD.n328 VDD.n327 185
R17699 VDD.n2259 VDD.n2258 185
R17700 VDD.n2258 VDD.n2257 185
R17701 VDD.n2260 VDD.n325 185
R17702 VDD.n325 VDD.n321 185
R17703 VDD.n2262 VDD.n2261 185
R17704 VDD.n2263 VDD.n2262 185
R17705 VDD.n315 VDD.n314 185
R17706 VDD.n324 VDD.n315 185
R17707 VDD.n2271 VDD.n2270 185
R17708 VDD.n2270 VDD.n2269 185
R17709 VDD.n2272 VDD.n313 185
R17710 VDD.n313 VDD.n310 185
R17711 VDD.n2274 VDD.n2273 185
R17712 VDD.n2275 VDD.n2274 185
R17713 VDD.n302 VDD.n301 185
R17714 VDD.n303 VDD.n302 185
R17715 VDD.n2333 VDD.n2332 185
R17716 VDD.n2332 VDD.n2331 185
R17717 VDD.n2334 VDD.n300 185
R17718 VDD.n300 VDD.n297 185
R17719 VDD.n2336 VDD.n2335 185
R17720 VDD.n2337 VDD.n2336 185
R17721 VDD.n291 VDD.n289 185
R17722 VDD.n289 VDD.n285 185
R17723 VDD.n2390 VDD.n2389 185
R17724 VDD.n2391 VDD.n2390 185
R17725 VDD.n2388 VDD.n290 185
R17726 VDD.n290 VDD.n287 185
R17727 VDD.n1221 VDD.n1220 185
R17728 VDD.n1178 VDD.n713 185
R17729 VDD.n1179 VDD.n1177 185
R17730 VDD.n1182 VDD.n1176 185
R17731 VDD.n1183 VDD.n1175 185
R17732 VDD.n1184 VDD.n1174 185
R17733 VDD.n1173 VDD.n1171 185
R17734 VDD.n1188 VDD.n1170 185
R17735 VDD.n1189 VDD.n1169 185
R17736 VDD.n1190 VDD.n1168 185
R17737 VDD.n1167 VDD.n1165 185
R17738 VDD.n1194 VDD.n1164 185
R17739 VDD.n1195 VDD.n1163 185
R17740 VDD.n1196 VDD.n1160 185
R17741 VDD.n1159 VDD.n1157 185
R17742 VDD.n1200 VDD.n1156 185
R17743 VDD.n1201 VDD.n1155 185
R17744 VDD.n1202 VDD.n1154 185
R17745 VDD.n1153 VDD.n1151 185
R17746 VDD.n1206 VDD.n1150 185
R17747 VDD.n1207 VDD.n1149 185
R17748 VDD.n1208 VDD.n1148 185
R17749 VDD.n1217 VDD.n714 185
R17750 VDD.n714 VDD.n702 185
R17751 VDD.n1216 VDD.n1215 185
R17752 VDD.n1215 VDD.n1214 185
R17753 VDD.n721 VDD.n720 185
R17754 VDD.n722 VDD.n721 185
R17755 VDD.n1141 VDD.n1140 185
R17756 VDD.n1142 VDD.n1141 185
R17757 VDD.n732 VDD.n731 185
R17758 VDD.n731 VDD.n730 185
R17759 VDD.n1135 VDD.n1134 185
R17760 VDD.n1134 VDD.n1133 185
R17761 VDD.n735 VDD.n734 185
R17762 VDD.n736 VDD.n735 185
R17763 VDD.n1124 VDD.n1123 185
R17764 VDD.n1125 VDD.n1124 185
R17765 VDD.n744 VDD.n743 185
R17766 VDD.n743 VDD.n742 185
R17767 VDD.n1119 VDD.n1118 185
R17768 VDD.n1118 VDD.n1117 185
R17769 VDD.n747 VDD.n746 185
R17770 VDD.n748 VDD.n747 185
R17771 VDD.n1108 VDD.n1107 185
R17772 VDD.n1109 VDD.n1108 185
R17773 VDD.n756 VDD.n755 185
R17774 VDD.n755 VDD.n754 185
R17775 VDD.n1103 VDD.n1102 185
R17776 VDD.n1102 VDD.n1101 185
R17777 VDD.n759 VDD.n758 185
R17778 VDD.n760 VDD.n759 185
R17779 VDD.n1092 VDD.n1091 185
R17780 VDD.n1093 VDD.n1092 185
R17781 VDD.n767 VDD.n766 185
R17782 VDD.n772 VDD.n766 185
R17783 VDD.n1087 VDD.n1086 185
R17784 VDD.n1086 VDD.n1085 185
R17785 VDD.n770 VDD.n769 185
R17786 VDD.n771 VDD.n770 185
R17787 VDD.n1076 VDD.n1075 185
R17788 VDD.n1077 VDD.n1076 185
R17789 VDD.n780 VDD.n779 185
R17790 VDD.n779 VDD.n778 185
R17791 VDD.n1071 VDD.n1070 185
R17792 VDD.n1070 VDD.n1069 185
R17793 VDD.n783 VDD.n782 185
R17794 VDD.n784 VDD.n783 185
R17795 VDD.n1060 VDD.n1059 185
R17796 VDD.n1061 VDD.n1060 185
R17797 VDD.n792 VDD.n791 185
R17798 VDD.n791 VDD.n790 185
R17799 VDD.n1055 VDD.n1054 185
R17800 VDD.n1054 VDD.n1053 185
R17801 VDD.n795 VDD.n794 185
R17802 VDD.n796 VDD.n795 185
R17803 VDD.n1037 VDD.n1036 185
R17804 VDD.n1038 VDD.n1037 185
R17805 VDD.n804 VDD.n803 185
R17806 VDD.n803 VDD.n802 185
R17807 VDD.n1032 VDD.n1031 185
R17808 VDD.n1031 VDD.n1030 185
R17809 VDD.n807 VDD.n806 185
R17810 VDD.n808 VDD.n807 185
R17811 VDD.n1021 VDD.n1020 185
R17812 VDD.n1022 VDD.n1021 185
R17813 VDD.n816 VDD.n815 185
R17814 VDD.n815 VDD.n814 185
R17815 VDD.n1016 VDD.n1015 185
R17816 VDD.n1015 VDD.n1014 185
R17817 VDD.n819 VDD.n818 185
R17818 VDD.n1005 VDD.n819 185
R17819 VDD.n1004 VDD.n1003 185
R17820 VDD.n1006 VDD.n1004 185
R17821 VDD.n827 VDD.n826 185
R17822 VDD.n826 VDD.n825 185
R17823 VDD.n999 VDD.n998 185
R17824 VDD.n998 VDD.n997 185
R17825 VDD.n830 VDD.n829 185
R17826 VDD.n831 VDD.n830 185
R17827 VDD.n988 VDD.n987 185
R17828 VDD.n989 VDD.n988 185
R17829 VDD.n839 VDD.n838 185
R17830 VDD.n838 VDD.n837 185
R17831 VDD.n983 VDD.n982 185
R17832 VDD.n982 VDD.n981 185
R17833 VDD.n842 VDD.n841 185
R17834 VDD.n843 VDD.n842 185
R17835 VDD.n972 VDD.n971 185
R17836 VDD.n973 VDD.n972 185
R17837 VDD.n851 VDD.n850 185
R17838 VDD.n850 VDD.n849 185
R17839 VDD.n967 VDD.n966 185
R17840 VDD.n966 VDD.n965 185
R17841 VDD.n854 VDD.n853 185
R17842 VDD.n855 VDD.n854 185
R17843 VDD.n956 VDD.n955 185
R17844 VDD.n957 VDD.n956 185
R17845 VDD.n863 VDD.n862 185
R17846 VDD.n862 VDD.n861 185
R17847 VDD.n951 VDD.n950 185
R17848 VDD.n950 VDD.n949 185
R17849 VDD.n944 VDD.n867 185
R17850 VDD.n943 VDD.n870 185
R17851 VDD.n942 VDD.n871 185
R17852 VDD.n871 VDD.n866 185
R17853 VDD.n874 VDD.n872 185
R17854 VDD.n938 VDD.n876 185
R17855 VDD.n937 VDD.n877 185
R17856 VDD.n936 VDD.n879 185
R17857 VDD.n882 VDD.n880 185
R17858 VDD.n932 VDD.n884 185
R17859 VDD.n931 VDD.n928 185
R17860 VDD.n926 VDD.n885 185
R17861 VDD.n925 VDD.n924 185
R17862 VDD.n890 VDD.n887 185
R17863 VDD.n920 VDD.n891 185
R17864 VDD.n919 VDD.n893 185
R17865 VDD.n918 VDD.n894 185
R17866 VDD.n898 VDD.n895 185
R17867 VDD.n914 VDD.n899 185
R17868 VDD.n913 VDD.n901 185
R17869 VDD.n912 VDD.n902 185
R17870 VDD.n909 VDD.n904 185
R17871 VDD.n905 VDD.n865 185
R17872 VDD.n866 VDD.n865 185
R17873 VDD.n726 VDD.n724 185
R17874 VDD.n724 VDD.n702 185
R17875 VDD.n1213 VDD.n1212 185
R17876 VDD.n1214 VDD.n1213 185
R17877 VDD.n725 VDD.n723 185
R17878 VDD.n723 VDD.n722 185
R17879 VDD.n1144 VDD.n1143 185
R17880 VDD.n1143 VDD.n1142 185
R17881 VDD.n729 VDD.n728 185
R17882 VDD.n730 VDD.n729 185
R17883 VDD.n1132 VDD.n1131 185
R17884 VDD.n1133 VDD.n1132 185
R17885 VDD.n738 VDD.n737 185
R17886 VDD.n737 VDD.n736 185
R17887 VDD.n1127 VDD.n1126 185
R17888 VDD.n1126 VDD.n1125 185
R17889 VDD.n741 VDD.n740 185
R17890 VDD.n742 VDD.n741 185
R17891 VDD.n1116 VDD.n1115 185
R17892 VDD.n1117 VDD.n1116 185
R17893 VDD.n750 VDD.n749 185
R17894 VDD.n749 VDD.n748 185
R17895 VDD.n1111 VDD.n1110 185
R17896 VDD.n1110 VDD.n1109 185
R17897 VDD.n753 VDD.n752 185
R17898 VDD.n754 VDD.n753 185
R17899 VDD.n1100 VDD.n1099 185
R17900 VDD.n1101 VDD.n1100 185
R17901 VDD.n762 VDD.n761 185
R17902 VDD.n761 VDD.n760 185
R17903 VDD.n1095 VDD.n1094 185
R17904 VDD.n1094 VDD.n1093 185
R17905 VDD.n765 VDD.n764 185
R17906 VDD.n772 VDD.n765 185
R17907 VDD.n1084 VDD.n1083 185
R17908 VDD.n1085 VDD.n1084 185
R17909 VDD.n774 VDD.n773 185
R17910 VDD.n773 VDD.n771 185
R17911 VDD.n1079 VDD.n1078 185
R17912 VDD.n1078 VDD.n1077 185
R17913 VDD.n777 VDD.n776 185
R17914 VDD.n778 VDD.n777 185
R17915 VDD.n1068 VDD.n1067 185
R17916 VDD.n1069 VDD.n1068 185
R17917 VDD.n786 VDD.n785 185
R17918 VDD.n785 VDD.n784 185
R17919 VDD.n1063 VDD.n1062 185
R17920 VDD.n1062 VDD.n1061 185
R17921 VDD.n789 VDD.n788 185
R17922 VDD.n790 VDD.n789 185
R17923 VDD.n1052 VDD.n1051 185
R17924 VDD.n1053 VDD.n1052 185
R17925 VDD.n798 VDD.n797 185
R17926 VDD.n797 VDD.n796 185
R17927 VDD.n1040 VDD.n1039 185
R17928 VDD.n1039 VDD.n1038 185
R17929 VDD.n801 VDD.n800 185
R17930 VDD.n802 VDD.n801 185
R17931 VDD.n1029 VDD.n1028 185
R17932 VDD.n1030 VDD.n1029 185
R17933 VDD.n810 VDD.n809 185
R17934 VDD.n809 VDD.n808 185
R17935 VDD.n1024 VDD.n1023 185
R17936 VDD.n1023 VDD.n1022 185
R17937 VDD.n813 VDD.n812 185
R17938 VDD.n814 VDD.n813 185
R17939 VDD.n1013 VDD.n1012 185
R17940 VDD.n1014 VDD.n1013 185
R17941 VDD.n821 VDD.n820 185
R17942 VDD.n1005 VDD.n820 185
R17943 VDD.n1008 VDD.n1007 185
R17944 VDD.n1007 VDD.n1006 185
R17945 VDD.n824 VDD.n823 185
R17946 VDD.n825 VDD.n824 185
R17947 VDD.n996 VDD.n995 185
R17948 VDD.n997 VDD.n996 185
R17949 VDD.n833 VDD.n832 185
R17950 VDD.n832 VDD.n831 185
R17951 VDD.n991 VDD.n990 185
R17952 VDD.n990 VDD.n989 185
R17953 VDD.n836 VDD.n835 185
R17954 VDD.n837 VDD.n836 185
R17955 VDD.n980 VDD.n979 185
R17956 VDD.n981 VDD.n980 185
R17957 VDD.n845 VDD.n844 185
R17958 VDD.n844 VDD.n843 185
R17959 VDD.n975 VDD.n974 185
R17960 VDD.n974 VDD.n973 185
R17961 VDD.n848 VDD.n847 185
R17962 VDD.n849 VDD.n848 185
R17963 VDD.n964 VDD.n963 185
R17964 VDD.n965 VDD.n964 185
R17965 VDD.n857 VDD.n856 185
R17966 VDD.n856 VDD.n855 185
R17967 VDD.n959 VDD.n958 185
R17968 VDD.n958 VDD.n957 185
R17969 VDD.n860 VDD.n859 185
R17970 VDD.n861 VDD.n860 185
R17971 VDD.n948 VDD.n947 185
R17972 VDD.n949 VDD.n948 185
R17973 VDD.t10 VDD.t109 163.325
R17974 VDD.t84 VDD.t21 163.325
R17975 VDD.n123 VDD.n122 146.341
R17976 VDD.n127 VDD.n126 146.341
R17977 VDD.n133 VDD.n132 146.341
R17978 VDD.n137 VDD.n136 146.341
R17979 VDD.n143 VDD.n142 146.341
R17980 VDD.n147 VDD.n146 146.341
R17981 VDD.n153 VDD.n152 146.341
R17982 VDD.n157 VDD.n156 146.341
R17983 VDD.n163 VDD.n162 146.341
R17984 VDD.n165 VDD.n102 146.341
R17985 VDD.n2479 VDD.n252 146.341
R17986 VDD.n2479 VDD.n243 146.341
R17987 VDD.n2489 VDD.n243 146.341
R17988 VDD.n2489 VDD.n239 146.341
R17989 VDD.n2495 VDD.n239 146.341
R17990 VDD.n2495 VDD.n232 146.341
R17991 VDD.n2505 VDD.n232 146.341
R17992 VDD.n2505 VDD.n228 146.341
R17993 VDD.n2511 VDD.n228 146.341
R17994 VDD.n2511 VDD.n220 146.341
R17995 VDD.n2521 VDD.n220 146.341
R17996 VDD.n2521 VDD.n216 146.341
R17997 VDD.n2527 VDD.n216 146.341
R17998 VDD.n2527 VDD.n208 146.341
R17999 VDD.n2537 VDD.n208 146.341
R18000 VDD.n2537 VDD.n204 146.341
R18001 VDD.n2543 VDD.n204 146.341
R18002 VDD.n2543 VDD.n196 146.341
R18003 VDD.n2553 VDD.n196 146.341
R18004 VDD.n2553 VDD.n191 146.341
R18005 VDD.n2562 VDD.n191 146.341
R18006 VDD.n2562 VDD.n192 146.341
R18007 VDD.n192 VDD.n183 146.341
R18008 VDD.n2573 VDD.n183 146.341
R18009 VDD.n2573 VDD.n27 146.341
R18010 VDD.n28 VDD.n27 146.341
R18011 VDD.n29 VDD.n28 146.341
R18012 VDD.n2580 VDD.n29 146.341
R18013 VDD.n2580 VDD.n37 146.341
R18014 VDD.n38 VDD.n37 146.341
R18015 VDD.n39 VDD.n38 146.341
R18016 VDD.n2587 VDD.n39 146.341
R18017 VDD.n2587 VDD.n48 146.341
R18018 VDD.n49 VDD.n48 146.341
R18019 VDD.n50 VDD.n49 146.341
R18020 VDD.n2594 VDD.n50 146.341
R18021 VDD.n2594 VDD.n59 146.341
R18022 VDD.n60 VDD.n59 146.341
R18023 VDD.n61 VDD.n60 146.341
R18024 VDD.n2601 VDD.n61 146.341
R18025 VDD.n2601 VDD.n70 146.341
R18026 VDD.n71 VDD.n70 146.341
R18027 VDD.n72 VDD.n71 146.341
R18028 VDD.n2608 VDD.n72 146.341
R18029 VDD.n2608 VDD.n81 146.341
R18030 VDD.n82 VDD.n81 146.341
R18031 VDD.n83 VDD.n82 146.341
R18032 VDD.n2615 VDD.n83 146.341
R18033 VDD.n2615 VDD.n91 146.341
R18034 VDD.n2409 VDD.n2408 146.341
R18035 VDD.n2465 VDD.n2408 146.341
R18036 VDD.n2463 VDD.n2462 146.341
R18037 VDD.n2459 VDD.n2458 146.341
R18038 VDD.n2455 VDD.n2454 146.341
R18039 VDD.n2451 VDD.n2450 146.341
R18040 VDD.n2447 VDD.n2446 146.341
R18041 VDD.n2443 VDD.n2442 146.341
R18042 VDD.n2439 VDD.n2438 146.341
R18043 VDD.n2435 VDD.n2434 146.341
R18044 VDD.n2473 VDD.n258 146.341
R18045 VDD.n2481 VDD.n250 146.341
R18046 VDD.n2481 VDD.n246 146.341
R18047 VDD.n2487 VDD.n246 146.341
R18048 VDD.n2487 VDD.n238 146.341
R18049 VDD.n2497 VDD.n238 146.341
R18050 VDD.n2497 VDD.n234 146.341
R18051 VDD.n2503 VDD.n234 146.341
R18052 VDD.n2503 VDD.n226 146.341
R18053 VDD.n2513 VDD.n226 146.341
R18054 VDD.n2513 VDD.n222 146.341
R18055 VDD.n2519 VDD.n222 146.341
R18056 VDD.n2519 VDD.n214 146.341
R18057 VDD.n2529 VDD.n214 146.341
R18058 VDD.n2529 VDD.n210 146.341
R18059 VDD.n2535 VDD.n210 146.341
R18060 VDD.n2535 VDD.n202 146.341
R18061 VDD.n2545 VDD.n202 146.341
R18062 VDD.n2545 VDD.n198 146.341
R18063 VDD.n2551 VDD.n198 146.341
R18064 VDD.n2551 VDD.n189 146.341
R18065 VDD.n2564 VDD.n189 146.341
R18066 VDD.n2564 VDD.n185 146.341
R18067 VDD.n2570 VDD.n185 146.341
R18068 VDD.n2570 VDD.n25 146.341
R18069 VDD.n2673 VDD.n25 146.341
R18070 VDD.n2673 VDD.n26 146.341
R18071 VDD.n2669 VDD.n26 146.341
R18072 VDD.n2669 VDD.n31 146.341
R18073 VDD.n2665 VDD.n31 146.341
R18074 VDD.n2665 VDD.n36 146.341
R18075 VDD.n2661 VDD.n36 146.341
R18076 VDD.n2661 VDD.n41 146.341
R18077 VDD.n2657 VDD.n41 146.341
R18078 VDD.n2657 VDD.n47 146.341
R18079 VDD.n2653 VDD.n47 146.341
R18080 VDD.n2653 VDD.n52 146.341
R18081 VDD.n2649 VDD.n52 146.341
R18082 VDD.n2649 VDD.n58 146.341
R18083 VDD.n2645 VDD.n58 146.341
R18084 VDD.n2645 VDD.n63 146.341
R18085 VDD.n2641 VDD.n63 146.341
R18086 VDD.n2641 VDD.n69 146.341
R18087 VDD.n2637 VDD.n69 146.341
R18088 VDD.n2637 VDD.n74 146.341
R18089 VDD.n2633 VDD.n74 146.341
R18090 VDD.n2633 VDD.n80 146.341
R18091 VDD.n2629 VDD.n80 146.341
R18092 VDD.n2629 VDD.n85 146.341
R18093 VDD.n2625 VDD.n85 146.341
R18094 VDD.n1150 VDD.n1149 146.341
R18095 VDD.n1154 VDD.n1153 146.341
R18096 VDD.n1156 VDD.n1155 146.341
R18097 VDD.n1160 VDD.n1159 146.341
R18098 VDD.n1164 VDD.n1163 146.341
R18099 VDD.n1168 VDD.n1167 146.341
R18100 VDD.n1170 VDD.n1169 146.341
R18101 VDD.n1174 VDD.n1173 146.341
R18102 VDD.n1176 VDD.n1175 146.341
R18103 VDD.n1177 VDD.n713 146.341
R18104 VDD.n950 VDD.n862 146.341
R18105 VDD.n956 VDD.n862 146.341
R18106 VDD.n956 VDD.n854 146.341
R18107 VDD.n966 VDD.n854 146.341
R18108 VDD.n966 VDD.n850 146.341
R18109 VDD.n972 VDD.n850 146.341
R18110 VDD.n972 VDD.n842 146.341
R18111 VDD.n982 VDD.n842 146.341
R18112 VDD.n982 VDD.n838 146.341
R18113 VDD.n988 VDD.n838 146.341
R18114 VDD.n988 VDD.n830 146.341
R18115 VDD.n998 VDD.n830 146.341
R18116 VDD.n998 VDD.n826 146.341
R18117 VDD.n1004 VDD.n826 146.341
R18118 VDD.n1004 VDD.n819 146.341
R18119 VDD.n1015 VDD.n819 146.341
R18120 VDD.n1015 VDD.n815 146.341
R18121 VDD.n1021 VDD.n815 146.341
R18122 VDD.n1021 VDD.n807 146.341
R18123 VDD.n1031 VDD.n807 146.341
R18124 VDD.n1031 VDD.n803 146.341
R18125 VDD.n1037 VDD.n803 146.341
R18126 VDD.n1037 VDD.n795 146.341
R18127 VDD.n1054 VDD.n795 146.341
R18128 VDD.n1054 VDD.n791 146.341
R18129 VDD.n1060 VDD.n791 146.341
R18130 VDD.n1060 VDD.n783 146.341
R18131 VDD.n1070 VDD.n783 146.341
R18132 VDD.n1070 VDD.n779 146.341
R18133 VDD.n1076 VDD.n779 146.341
R18134 VDD.n1076 VDD.n770 146.341
R18135 VDD.n1086 VDD.n770 146.341
R18136 VDD.n1086 VDD.n766 146.341
R18137 VDD.n1092 VDD.n766 146.341
R18138 VDD.n1092 VDD.n759 146.341
R18139 VDD.n1102 VDD.n759 146.341
R18140 VDD.n1102 VDD.n755 146.341
R18141 VDD.n1108 VDD.n755 146.341
R18142 VDD.n1108 VDD.n747 146.341
R18143 VDD.n1118 VDD.n747 146.341
R18144 VDD.n1118 VDD.n743 146.341
R18145 VDD.n1124 VDD.n743 146.341
R18146 VDD.n1124 VDD.n735 146.341
R18147 VDD.n1134 VDD.n735 146.341
R18148 VDD.n1134 VDD.n731 146.341
R18149 VDD.n1141 VDD.n731 146.341
R18150 VDD.n1141 VDD.n721 146.341
R18151 VDD.n1215 VDD.n721 146.341
R18152 VDD.n1215 VDD.n714 146.341
R18153 VDD.n871 VDD.n870 146.341
R18154 VDD.n874 VDD.n871 146.341
R18155 VDD.n877 VDD.n876 146.341
R18156 VDD.n882 VDD.n879 146.341
R18157 VDD.n928 VDD.n884 146.341
R18158 VDD.n926 VDD.n925 146.341
R18159 VDD.n891 VDD.n890 146.341
R18160 VDD.n894 VDD.n893 146.341
R18161 VDD.n899 VDD.n898 146.341
R18162 VDD.n902 VDD.n901 146.341
R18163 VDD.n904 VDD.n865 146.341
R18164 VDD.n948 VDD.n860 146.341
R18165 VDD.n958 VDD.n860 146.341
R18166 VDD.n958 VDD.n856 146.341
R18167 VDD.n964 VDD.n856 146.341
R18168 VDD.n964 VDD.n848 146.341
R18169 VDD.n974 VDD.n848 146.341
R18170 VDD.n974 VDD.n844 146.341
R18171 VDD.n980 VDD.n844 146.341
R18172 VDD.n980 VDD.n836 146.341
R18173 VDD.n990 VDD.n836 146.341
R18174 VDD.n990 VDD.n832 146.341
R18175 VDD.n996 VDD.n832 146.341
R18176 VDD.n996 VDD.n824 146.341
R18177 VDD.n1007 VDD.n824 146.341
R18178 VDD.n1007 VDD.n820 146.341
R18179 VDD.n1013 VDD.n820 146.341
R18180 VDD.n1013 VDD.n813 146.341
R18181 VDD.n1023 VDD.n813 146.341
R18182 VDD.n1023 VDD.n809 146.341
R18183 VDD.n1029 VDD.n809 146.341
R18184 VDD.n1029 VDD.n801 146.341
R18185 VDD.n1039 VDD.n801 146.341
R18186 VDD.n1039 VDD.n797 146.341
R18187 VDD.n1052 VDD.n797 146.341
R18188 VDD.n1052 VDD.n789 146.341
R18189 VDD.n1062 VDD.n789 146.341
R18190 VDD.n1062 VDD.n785 146.341
R18191 VDD.n1068 VDD.n785 146.341
R18192 VDD.n1068 VDD.n777 146.341
R18193 VDD.n1078 VDD.n777 146.341
R18194 VDD.n1078 VDD.n773 146.341
R18195 VDD.n1084 VDD.n773 146.341
R18196 VDD.n1084 VDD.n765 146.341
R18197 VDD.n1094 VDD.n765 146.341
R18198 VDD.n1094 VDD.n761 146.341
R18199 VDD.n1100 VDD.n761 146.341
R18200 VDD.n1100 VDD.n753 146.341
R18201 VDD.n1110 VDD.n753 146.341
R18202 VDD.n1110 VDD.n749 146.341
R18203 VDD.n1116 VDD.n749 146.341
R18204 VDD.n1116 VDD.n741 146.341
R18205 VDD.n1126 VDD.n741 146.341
R18206 VDD.n1126 VDD.n737 146.341
R18207 VDD.n1132 VDD.n737 146.341
R18208 VDD.n1132 VDD.n729 146.341
R18209 VDD.n1143 VDD.n729 146.341
R18210 VDD.n1143 VDD.n723 146.341
R18211 VDD.n1213 VDD.n723 146.341
R18212 VDD.n1213 VDD.n724 146.341
R18213 VDD.n907 VDD.t28 128.627
R18214 VDD.n930 VDD.t39 128.627
R18215 VDD.n2421 VDD.t74 128.627
R18216 VDD.n256 VDD.t68 128.627
R18217 VDD.n104 VDD.t33 128.627
R18218 VDD.n112 VDD.t43 128.627
R18219 VDD.n1162 VDD.t65 128.627
R18220 VDD.n716 VDD.t62 128.627
R18221 VDD.t85 VDD.t10 126.237
R18222 VDD.t21 VDD.t8 126.237
R18223 VDD.n1510 VDD.t85 124.195
R18224 VDD.t8 VDD.n2398 124.195
R18225 VDD.n1809 VDD.n1808 123.514
R18226 VDD.n1046 VDD.t104 117.023
R18227 VDD.n1044 VDD.t99 117.023
R18228 VDD.n19 VDD.t102 113.24
R18229 VDD.n17 VDD.t97 113.24
R18230 VDD.n19 VDD.n18 107.79
R18231 VDD.n17 VDD.n16 107.79
R18232 VDD.n1046 VDD.n1045 104.005
R18233 VDD.n1044 VDD.n1043 104.005
R18234 VDD.n9 VDD.n7 101.112
R18235 VDD.n2 VDD.n0 101.112
R18236 VDD.n2106 VDD.n471 99.5127
R18237 VDD.n2114 VDD.n471 99.5127
R18238 VDD.n2114 VDD.n469 99.5127
R18239 VDD.n2118 VDD.n469 99.5127
R18240 VDD.n2118 VDD.n459 99.5127
R18241 VDD.n2126 VDD.n459 99.5127
R18242 VDD.n2126 VDD.n457 99.5127
R18243 VDD.n2130 VDD.n457 99.5127
R18244 VDD.n2130 VDD.n447 99.5127
R18245 VDD.n2138 VDD.n447 99.5127
R18246 VDD.n2138 VDD.n445 99.5127
R18247 VDD.n2142 VDD.n445 99.5127
R18248 VDD.n2142 VDD.n434 99.5127
R18249 VDD.n2150 VDD.n434 99.5127
R18250 VDD.n2150 VDD.n432 99.5127
R18251 VDD.n2154 VDD.n432 99.5127
R18252 VDD.n2154 VDD.n423 99.5127
R18253 VDD.n2162 VDD.n423 99.5127
R18254 VDD.n2162 VDD.n421 99.5127
R18255 VDD.n2166 VDD.n421 99.5127
R18256 VDD.n2166 VDD.n411 99.5127
R18257 VDD.n2174 VDD.n411 99.5127
R18258 VDD.n2174 VDD.n409 99.5127
R18259 VDD.n2178 VDD.n409 99.5127
R18260 VDD.n2178 VDD.n399 99.5127
R18261 VDD.n2186 VDD.n399 99.5127
R18262 VDD.n2186 VDD.n397 99.5127
R18263 VDD.n2190 VDD.n397 99.5127
R18264 VDD.n2190 VDD.n386 99.5127
R18265 VDD.n2198 VDD.n386 99.5127
R18266 VDD.n2198 VDD.n384 99.5127
R18267 VDD.n2202 VDD.n384 99.5127
R18268 VDD.n2202 VDD.n375 99.5127
R18269 VDD.n2210 VDD.n375 99.5127
R18270 VDD.n2210 VDD.n373 99.5127
R18271 VDD.n2214 VDD.n373 99.5127
R18272 VDD.n2214 VDD.n363 99.5127
R18273 VDD.n2222 VDD.n363 99.5127
R18274 VDD.n2222 VDD.n361 99.5127
R18275 VDD.n2226 VDD.n361 99.5127
R18276 VDD.n2226 VDD.n351 99.5127
R18277 VDD.n2234 VDD.n351 99.5127
R18278 VDD.n2234 VDD.n349 99.5127
R18279 VDD.n2238 VDD.n349 99.5127
R18280 VDD.n2238 VDD.n339 99.5127
R18281 VDD.n2246 VDD.n339 99.5127
R18282 VDD.n2246 VDD.n337 99.5127
R18283 VDD.n2250 VDD.n337 99.5127
R18284 VDD.n2250 VDD.n327 99.5127
R18285 VDD.n2258 VDD.n327 99.5127
R18286 VDD.n2258 VDD.n325 99.5127
R18287 VDD.n2262 VDD.n325 99.5127
R18288 VDD.n2262 VDD.n315 99.5127
R18289 VDD.n2270 VDD.n315 99.5127
R18290 VDD.n2270 VDD.n313 99.5127
R18291 VDD.n2274 VDD.n313 99.5127
R18292 VDD.n2274 VDD.n302 99.5127
R18293 VDD.n2332 VDD.n302 99.5127
R18294 VDD.n2332 VDD.n300 99.5127
R18295 VDD.n2336 VDD.n300 99.5127
R18296 VDD.n2336 VDD.n289 99.5127
R18297 VDD.n2390 VDD.n289 99.5127
R18298 VDD.n2390 VDD.n290 99.5127
R18299 VDD.n2384 VDD.n2383 99.5127
R18300 VDD.n2380 VDD.n2379 99.5127
R18301 VDD.n2376 VDD.n2375 99.5127
R18302 VDD.n2372 VDD.n2371 99.5127
R18303 VDD.n2368 VDD.n2367 99.5127
R18304 VDD.n2364 VDD.n2363 99.5127
R18305 VDD.n2360 VDD.n2359 99.5127
R18306 VDD.n2356 VDD.n2355 99.5127
R18307 VDD.n2352 VDD.n2351 99.5127
R18308 VDD.n2348 VDD.n2347 99.5127
R18309 VDD.n2058 VDD.n1810 99.5127
R18310 VDD.n2058 VDD.n473 99.5127
R18311 VDD.n2055 VDD.n473 99.5127
R18312 VDD.n2055 VDD.n467 99.5127
R18313 VDD.n2052 VDD.n467 99.5127
R18314 VDD.n2052 VDD.n461 99.5127
R18315 VDD.n2049 VDD.n461 99.5127
R18316 VDD.n2049 VDD.n455 99.5127
R18317 VDD.n2046 VDD.n455 99.5127
R18318 VDD.n2046 VDD.n449 99.5127
R18319 VDD.n2043 VDD.n449 99.5127
R18320 VDD.n2043 VDD.n443 99.5127
R18321 VDD.n2040 VDD.n443 99.5127
R18322 VDD.n2040 VDD.n436 99.5127
R18323 VDD.n2037 VDD.n436 99.5127
R18324 VDD.n2037 VDD.n430 99.5127
R18325 VDD.n2034 VDD.n430 99.5127
R18326 VDD.n2034 VDD.n425 99.5127
R18327 VDD.n2031 VDD.n425 99.5127
R18328 VDD.n2031 VDD.n419 99.5127
R18329 VDD.n2028 VDD.n419 99.5127
R18330 VDD.n2028 VDD.n413 99.5127
R18331 VDD.n2025 VDD.n413 99.5127
R18332 VDD.n2025 VDD.n407 99.5127
R18333 VDD.n2022 VDD.n407 99.5127
R18334 VDD.n2022 VDD.n401 99.5127
R18335 VDD.n2019 VDD.n401 99.5127
R18336 VDD.n2019 VDD.n395 99.5127
R18337 VDD.n2016 VDD.n395 99.5127
R18338 VDD.n2016 VDD.n388 99.5127
R18339 VDD.n2013 VDD.n388 99.5127
R18340 VDD.n2013 VDD.n382 99.5127
R18341 VDD.n2010 VDD.n382 99.5127
R18342 VDD.n2010 VDD.n377 99.5127
R18343 VDD.n2007 VDD.n377 99.5127
R18344 VDD.n2007 VDD.n370 99.5127
R18345 VDD.n2004 VDD.n370 99.5127
R18346 VDD.n2004 VDD.n364 99.5127
R18347 VDD.n2001 VDD.n364 99.5127
R18348 VDD.n2001 VDD.n359 99.5127
R18349 VDD.n1998 VDD.n359 99.5127
R18350 VDD.n1998 VDD.n353 99.5127
R18351 VDD.n1995 VDD.n353 99.5127
R18352 VDD.n1995 VDD.n347 99.5127
R18353 VDD.n1992 VDD.n347 99.5127
R18354 VDD.n1992 VDD.n341 99.5127
R18355 VDD.n1989 VDD.n341 99.5127
R18356 VDD.n1989 VDD.n335 99.5127
R18357 VDD.n1986 VDD.n335 99.5127
R18358 VDD.n1986 VDD.n329 99.5127
R18359 VDD.n1983 VDD.n329 99.5127
R18360 VDD.n1983 VDD.n322 99.5127
R18361 VDD.n1980 VDD.n322 99.5127
R18362 VDD.n1980 VDD.n316 99.5127
R18363 VDD.n1977 VDD.n316 99.5127
R18364 VDD.n1977 VDD.n311 99.5127
R18365 VDD.n1974 VDD.n311 99.5127
R18366 VDD.n1974 VDD.n304 99.5127
R18367 VDD.n304 VDD.n296 99.5127
R18368 VDD.n2338 VDD.n296 99.5127
R18369 VDD.n2339 VDD.n2338 99.5127
R18370 VDD.n2339 VDD.n286 99.5127
R18371 VDD.n2343 VDD.n286 99.5127
R18372 VDD.n2102 VDD.n2100 99.5127
R18373 VDD.n2100 VDD.n2099 99.5127
R18374 VDD.n2096 VDD.n2095 99.5127
R18375 VDD.n2093 VDD.n1963 99.5127
R18376 VDD.n2089 VDD.n2087 99.5127
R18377 VDD.n2085 VDD.n1965 99.5127
R18378 VDD.n2081 VDD.n2079 99.5127
R18379 VDD.n2077 VDD.n1967 99.5127
R18380 VDD.n2073 VDD.n2071 99.5127
R18381 VDD.n2069 VDD.n1969 99.5127
R18382 VDD.n2064 VDD.n2062 99.5127
R18383 VDD.n1794 VDD.n1793 99.5127
R18384 VDD.n1790 VDD.n1789 99.5127
R18385 VDD.n1786 VDD.n1785 99.5127
R18386 VDD.n1782 VDD.n1781 99.5127
R18387 VDD.n1778 VDD.n1777 99.5127
R18388 VDD.n1774 VDD.n1773 99.5127
R18389 VDD.n1770 VDD.n1769 99.5127
R18390 VDD.n1766 VDD.n1765 99.5127
R18391 VDD.n1762 VDD.n1761 99.5127
R18392 VDD.n1758 VDD.n1757 99.5127
R18393 VDD.n1358 VDD.n697 99.5127
R18394 VDD.n1358 VDD.n692 99.5127
R18395 VDD.n1355 VDD.n692 99.5127
R18396 VDD.n1355 VDD.n686 99.5127
R18397 VDD.n1352 VDD.n686 99.5127
R18398 VDD.n1352 VDD.n680 99.5127
R18399 VDD.n1349 VDD.n680 99.5127
R18400 VDD.n1349 VDD.n673 99.5127
R18401 VDD.n1346 VDD.n673 99.5127
R18402 VDD.n1346 VDD.n667 99.5127
R18403 VDD.n1343 VDD.n667 99.5127
R18404 VDD.n1343 VDD.n662 99.5127
R18405 VDD.n1340 VDD.n662 99.5127
R18406 VDD.n1340 VDD.n656 99.5127
R18407 VDD.n1337 VDD.n656 99.5127
R18408 VDD.n1337 VDD.n650 99.5127
R18409 VDD.n1334 VDD.n650 99.5127
R18410 VDD.n1334 VDD.n644 99.5127
R18411 VDD.n1331 VDD.n644 99.5127
R18412 VDD.n1331 VDD.n638 99.5127
R18413 VDD.n1328 VDD.n638 99.5127
R18414 VDD.n1328 VDD.n632 99.5127
R18415 VDD.n1325 VDD.n632 99.5127
R18416 VDD.n1325 VDD.n625 99.5127
R18417 VDD.n1322 VDD.n625 99.5127
R18418 VDD.n1322 VDD.n619 99.5127
R18419 VDD.n1319 VDD.n619 99.5127
R18420 VDD.n1319 VDD.n614 99.5127
R18421 VDD.n1316 VDD.n614 99.5127
R18422 VDD.n1316 VDD.n607 99.5127
R18423 VDD.n1313 VDD.n607 99.5127
R18424 VDD.n1313 VDD.n601 99.5127
R18425 VDD.n1310 VDD.n601 99.5127
R18426 VDD.n1310 VDD.n596 99.5127
R18427 VDD.n1307 VDD.n596 99.5127
R18428 VDD.n1307 VDD.n590 99.5127
R18429 VDD.n1304 VDD.n590 99.5127
R18430 VDD.n1304 VDD.n584 99.5127
R18431 VDD.n1301 VDD.n584 99.5127
R18432 VDD.n1301 VDD.n578 99.5127
R18433 VDD.n1298 VDD.n578 99.5127
R18434 VDD.n1298 VDD.n572 99.5127
R18435 VDD.n1295 VDD.n572 99.5127
R18436 VDD.n1295 VDD.n566 99.5127
R18437 VDD.n1292 VDD.n566 99.5127
R18438 VDD.n1292 VDD.n559 99.5127
R18439 VDD.n1289 VDD.n559 99.5127
R18440 VDD.n1289 VDD.n553 99.5127
R18441 VDD.n1286 VDD.n553 99.5127
R18442 VDD.n1286 VDD.n548 99.5127
R18443 VDD.n1283 VDD.n548 99.5127
R18444 VDD.n1283 VDD.n542 99.5127
R18445 VDD.n1280 VDD.n542 99.5127
R18446 VDD.n1280 VDD.n536 99.5127
R18447 VDD.n1277 VDD.n536 99.5127
R18448 VDD.n1277 VDD.n530 99.5127
R18449 VDD.n1274 VDD.n530 99.5127
R18450 VDD.n1274 VDD.n523 99.5127
R18451 VDD.n523 VDD.n515 99.5127
R18452 VDD.n1748 VDD.n515 99.5127
R18453 VDD.n1749 VDD.n1748 99.5127
R18454 VDD.n1749 VDD.n506 99.5127
R18455 VDD.n1753 VDD.n506 99.5127
R18456 VDD.n1512 VDD.n701 99.5127
R18457 VDD.n1236 VDD.n701 99.5127
R18458 VDD.n1240 VDD.n1239 99.5127
R18459 VDD.n1244 VDD.n1243 99.5127
R18460 VDD.n1248 VDD.n1247 99.5127
R18461 VDD.n1252 VDD.n1251 99.5127
R18462 VDD.n1256 VDD.n1255 99.5127
R18463 VDD.n1260 VDD.n1259 99.5127
R18464 VDD.n1264 VDD.n1263 99.5127
R18465 VDD.n1268 VDD.n1267 99.5127
R18466 VDD.n1362 VDD.n1233 99.5127
R18467 VDD.n1516 VDD.n690 99.5127
R18468 VDD.n1524 VDD.n690 99.5127
R18469 VDD.n1524 VDD.n688 99.5127
R18470 VDD.n1528 VDD.n688 99.5127
R18471 VDD.n1528 VDD.n678 99.5127
R18472 VDD.n1536 VDD.n678 99.5127
R18473 VDD.n1536 VDD.n676 99.5127
R18474 VDD.n1540 VDD.n676 99.5127
R18475 VDD.n1540 VDD.n666 99.5127
R18476 VDD.n1548 VDD.n666 99.5127
R18477 VDD.n1548 VDD.n664 99.5127
R18478 VDD.n1552 VDD.n664 99.5127
R18479 VDD.n1552 VDD.n654 99.5127
R18480 VDD.n1560 VDD.n654 99.5127
R18481 VDD.n1560 VDD.n652 99.5127
R18482 VDD.n1564 VDD.n652 99.5127
R18483 VDD.n1564 VDD.n642 99.5127
R18484 VDD.n1572 VDD.n642 99.5127
R18485 VDD.n1572 VDD.n640 99.5127
R18486 VDD.n1576 VDD.n640 99.5127
R18487 VDD.n1576 VDD.n630 99.5127
R18488 VDD.n1584 VDD.n630 99.5127
R18489 VDD.n1584 VDD.n628 99.5127
R18490 VDD.n1588 VDD.n628 99.5127
R18491 VDD.n1588 VDD.n618 99.5127
R18492 VDD.n1596 VDD.n618 99.5127
R18493 VDD.n1596 VDD.n616 99.5127
R18494 VDD.n1600 VDD.n616 99.5127
R18495 VDD.n1600 VDD.n605 99.5127
R18496 VDD.n1608 VDD.n605 99.5127
R18497 VDD.n1608 VDD.n603 99.5127
R18498 VDD.n1612 VDD.n603 99.5127
R18499 VDD.n1612 VDD.n594 99.5127
R18500 VDD.n1620 VDD.n594 99.5127
R18501 VDD.n1620 VDD.n592 99.5127
R18502 VDD.n1624 VDD.n592 99.5127
R18503 VDD.n1624 VDD.n582 99.5127
R18504 VDD.n1632 VDD.n582 99.5127
R18505 VDD.n1632 VDD.n580 99.5127
R18506 VDD.n1636 VDD.n580 99.5127
R18507 VDD.n1636 VDD.n570 99.5127
R18508 VDD.n1644 VDD.n570 99.5127
R18509 VDD.n1644 VDD.n568 99.5127
R18510 VDD.n1648 VDD.n568 99.5127
R18511 VDD.n1648 VDD.n557 99.5127
R18512 VDD.n1656 VDD.n557 99.5127
R18513 VDD.n1656 VDD.n555 99.5127
R18514 VDD.n1660 VDD.n555 99.5127
R18515 VDD.n1660 VDD.n546 99.5127
R18516 VDD.n1668 VDD.n546 99.5127
R18517 VDD.n1668 VDD.n544 99.5127
R18518 VDD.n1672 VDD.n544 99.5127
R18519 VDD.n1672 VDD.n534 99.5127
R18520 VDD.n1680 VDD.n534 99.5127
R18521 VDD.n1680 VDD.n532 99.5127
R18522 VDD.n1684 VDD.n532 99.5127
R18523 VDD.n1684 VDD.n521 99.5127
R18524 VDD.n1742 VDD.n521 99.5127
R18525 VDD.n1742 VDD.n519 99.5127
R18526 VDD.n1746 VDD.n519 99.5127
R18527 VDD.n1746 VDD.n508 99.5127
R18528 VDD.n1800 VDD.n508 99.5127
R18529 VDD.n1800 VDD.n509 99.5127
R18530 VDD.n2318 VDD.n2317 99.5127
R18531 VDD.n2314 VDD.n2313 99.5127
R18532 VDD.n2310 VDD.n2309 99.5127
R18533 VDD.n2306 VDD.n2305 99.5127
R18534 VDD.n2302 VDD.n2301 99.5127
R18535 VDD.n2298 VDD.n2297 99.5127
R18536 VDD.n2294 VDD.n2293 99.5127
R18537 VDD.n2290 VDD.n2289 99.5127
R18538 VDD.n2286 VDD.n2285 99.5127
R18539 VDD.n2282 VDD.n280 99.5127
R18540 VDD.n1958 VDD.n1812 99.5127
R18541 VDD.n1812 VDD.n474 99.5127
R18542 VDD.n1953 VDD.n474 99.5127
R18543 VDD.n1953 VDD.n468 99.5127
R18544 VDD.n1950 VDD.n468 99.5127
R18545 VDD.n1950 VDD.n462 99.5127
R18546 VDD.n1947 VDD.n462 99.5127
R18547 VDD.n1947 VDD.n456 99.5127
R18548 VDD.n1944 VDD.n456 99.5127
R18549 VDD.n1944 VDD.n450 99.5127
R18550 VDD.n1941 VDD.n450 99.5127
R18551 VDD.n1941 VDD.n444 99.5127
R18552 VDD.n1938 VDD.n444 99.5127
R18553 VDD.n1938 VDD.n437 99.5127
R18554 VDD.n1935 VDD.n437 99.5127
R18555 VDD.n1935 VDD.n431 99.5127
R18556 VDD.n1932 VDD.n431 99.5127
R18557 VDD.n1932 VDD.n426 99.5127
R18558 VDD.n1929 VDD.n426 99.5127
R18559 VDD.n1929 VDD.n420 99.5127
R18560 VDD.n1926 VDD.n420 99.5127
R18561 VDD.n1926 VDD.n414 99.5127
R18562 VDD.n1923 VDD.n414 99.5127
R18563 VDD.n1923 VDD.n408 99.5127
R18564 VDD.n1920 VDD.n408 99.5127
R18565 VDD.n1920 VDD.n402 99.5127
R18566 VDD.n1917 VDD.n402 99.5127
R18567 VDD.n1917 VDD.n396 99.5127
R18568 VDD.n1914 VDD.n396 99.5127
R18569 VDD.n1914 VDD.n389 99.5127
R18570 VDD.n1911 VDD.n389 99.5127
R18571 VDD.n1911 VDD.n383 99.5127
R18572 VDD.n1908 VDD.n383 99.5127
R18573 VDD.n1908 VDD.n378 99.5127
R18574 VDD.n1905 VDD.n378 99.5127
R18575 VDD.n1905 VDD.n371 99.5127
R18576 VDD.n1902 VDD.n371 99.5127
R18577 VDD.n1902 VDD.n365 99.5127
R18578 VDD.n1899 VDD.n365 99.5127
R18579 VDD.n1899 VDD.n360 99.5127
R18580 VDD.n1896 VDD.n360 99.5127
R18581 VDD.n1896 VDD.n354 99.5127
R18582 VDD.n1893 VDD.n354 99.5127
R18583 VDD.n1893 VDD.n348 99.5127
R18584 VDD.n1890 VDD.n348 99.5127
R18585 VDD.n1890 VDD.n342 99.5127
R18586 VDD.n1887 VDD.n342 99.5127
R18587 VDD.n1887 VDD.n336 99.5127
R18588 VDD.n1884 VDD.n336 99.5127
R18589 VDD.n1884 VDD.n330 99.5127
R18590 VDD.n1881 VDD.n330 99.5127
R18591 VDD.n1881 VDD.n323 99.5127
R18592 VDD.n1878 VDD.n323 99.5127
R18593 VDD.n1878 VDD.n317 99.5127
R18594 VDD.n1875 VDD.n317 99.5127
R18595 VDD.n1875 VDD.n312 99.5127
R18596 VDD.n1872 VDD.n312 99.5127
R18597 VDD.n1872 VDD.n305 99.5127
R18598 VDD.n1869 VDD.n305 99.5127
R18599 VDD.n1869 VDD.n298 99.5127
R18600 VDD.n298 VDD.n284 99.5127
R18601 VDD.n2392 VDD.n284 99.5127
R18602 VDD.n2392 VDD.n281 99.5127
R18603 VDD.n1829 VDD.n1826 99.5127
R18604 VDD.n1833 VDD.n1831 99.5127
R18605 VDD.n1837 VDD.n1823 99.5127
R18606 VDD.n1841 VDD.n1839 99.5127
R18607 VDD.n1845 VDD.n1821 99.5127
R18608 VDD.n1849 VDD.n1847 99.5127
R18609 VDD.n1853 VDD.n1819 99.5127
R18610 VDD.n1857 VDD.n1855 99.5127
R18611 VDD.n1861 VDD.n1817 99.5127
R18612 VDD.n1865 VDD.n1863 99.5127
R18613 VDD.n2108 VDD.n475 99.5127
R18614 VDD.n2112 VDD.n475 99.5127
R18615 VDD.n2112 VDD.n465 99.5127
R18616 VDD.n2120 VDD.n465 99.5127
R18617 VDD.n2120 VDD.n463 99.5127
R18618 VDD.n2124 VDD.n463 99.5127
R18619 VDD.n2124 VDD.n453 99.5127
R18620 VDD.n2132 VDD.n453 99.5127
R18621 VDD.n2132 VDD.n451 99.5127
R18622 VDD.n2136 VDD.n451 99.5127
R18623 VDD.n2136 VDD.n441 99.5127
R18624 VDD.n2144 VDD.n441 99.5127
R18625 VDD.n2144 VDD.n439 99.5127
R18626 VDD.n2148 VDD.n439 99.5127
R18627 VDD.n2148 VDD.n429 99.5127
R18628 VDD.n2156 VDD.n429 99.5127
R18629 VDD.n2156 VDD.n427 99.5127
R18630 VDD.n2160 VDD.n427 99.5127
R18631 VDD.n2160 VDD.n417 99.5127
R18632 VDD.n2168 VDD.n417 99.5127
R18633 VDD.n2168 VDD.n415 99.5127
R18634 VDD.n2172 VDD.n415 99.5127
R18635 VDD.n2172 VDD.n405 99.5127
R18636 VDD.n2180 VDD.n405 99.5127
R18637 VDD.n2180 VDD.n403 99.5127
R18638 VDD.n2184 VDD.n403 99.5127
R18639 VDD.n2184 VDD.n393 99.5127
R18640 VDD.n2192 VDD.n393 99.5127
R18641 VDD.n2192 VDD.n391 99.5127
R18642 VDD.n2196 VDD.n391 99.5127
R18643 VDD.n2196 VDD.n381 99.5127
R18644 VDD.n2204 VDD.n381 99.5127
R18645 VDD.n2204 VDD.n379 99.5127
R18646 VDD.n2208 VDD.n379 99.5127
R18647 VDD.n2208 VDD.n368 99.5127
R18648 VDD.n2216 VDD.n368 99.5127
R18649 VDD.n2216 VDD.n366 99.5127
R18650 VDD.n2220 VDD.n366 99.5127
R18651 VDD.n2220 VDD.n357 99.5127
R18652 VDD.n2228 VDD.n357 99.5127
R18653 VDD.n2228 VDD.n355 99.5127
R18654 VDD.n2232 VDD.n355 99.5127
R18655 VDD.n2232 VDD.n345 99.5127
R18656 VDD.n2240 VDD.n345 99.5127
R18657 VDD.n2240 VDD.n343 99.5127
R18658 VDD.n2244 VDD.n343 99.5127
R18659 VDD.n2244 VDD.n333 99.5127
R18660 VDD.n2252 VDD.n333 99.5127
R18661 VDD.n2252 VDD.n331 99.5127
R18662 VDD.n2256 VDD.n331 99.5127
R18663 VDD.n2256 VDD.n320 99.5127
R18664 VDD.n2264 VDD.n320 99.5127
R18665 VDD.n2264 VDD.n318 99.5127
R18666 VDD.n2268 VDD.n318 99.5127
R18667 VDD.n2268 VDD.n309 99.5127
R18668 VDD.n2276 VDD.n309 99.5127
R18669 VDD.n2276 VDD.n306 99.5127
R18670 VDD.n2330 VDD.n306 99.5127
R18671 VDD.n2330 VDD.n307 99.5127
R18672 VDD.n307 VDD.n299 99.5127
R18673 VDD.n2325 VDD.n299 99.5127
R18674 VDD.n2325 VDD.n288 99.5127
R18675 VDD.n2322 VDD.n288 99.5127
R18676 VDD.n1728 VDD.n1727 99.5127
R18677 VDD.n1724 VDD.n1723 99.5127
R18678 VDD.n1720 VDD.n1719 99.5127
R18679 VDD.n1716 VDD.n1715 99.5127
R18680 VDD.n1712 VDD.n1711 99.5127
R18681 VDD.n1708 VDD.n1707 99.5127
R18682 VDD.n1704 VDD.n1703 99.5127
R18683 VDD.n1700 VDD.n1699 99.5127
R18684 VDD.n1696 VDD.n1695 99.5127
R18685 VDD.n1692 VDD.n500 99.5127
R18686 VDD.n1465 VDD.n698 99.5127
R18687 VDD.n1465 VDD.n693 99.5127
R18688 VDD.n1462 VDD.n693 99.5127
R18689 VDD.n1462 VDD.n687 99.5127
R18690 VDD.n1459 VDD.n687 99.5127
R18691 VDD.n1459 VDD.n681 99.5127
R18692 VDD.n1456 VDD.n681 99.5127
R18693 VDD.n1456 VDD.n674 99.5127
R18694 VDD.n1453 VDD.n674 99.5127
R18695 VDD.n1453 VDD.n668 99.5127
R18696 VDD.n1450 VDD.n668 99.5127
R18697 VDD.n1450 VDD.n663 99.5127
R18698 VDD.n1447 VDD.n663 99.5127
R18699 VDD.n1447 VDD.n657 99.5127
R18700 VDD.n1444 VDD.n657 99.5127
R18701 VDD.n1444 VDD.n651 99.5127
R18702 VDD.n1441 VDD.n651 99.5127
R18703 VDD.n1441 VDD.n645 99.5127
R18704 VDD.n1438 VDD.n645 99.5127
R18705 VDD.n1438 VDD.n639 99.5127
R18706 VDD.n1435 VDD.n639 99.5127
R18707 VDD.n1435 VDD.n633 99.5127
R18708 VDD.n1432 VDD.n633 99.5127
R18709 VDD.n1432 VDD.n626 99.5127
R18710 VDD.n1429 VDD.n626 99.5127
R18711 VDD.n1429 VDD.n620 99.5127
R18712 VDD.n1426 VDD.n620 99.5127
R18713 VDD.n1426 VDD.n615 99.5127
R18714 VDD.n1423 VDD.n615 99.5127
R18715 VDD.n1423 VDD.n608 99.5127
R18716 VDD.n1420 VDD.n608 99.5127
R18717 VDD.n1420 VDD.n602 99.5127
R18718 VDD.n1417 VDD.n602 99.5127
R18719 VDD.n1417 VDD.n597 99.5127
R18720 VDD.n1414 VDD.n597 99.5127
R18721 VDD.n1414 VDD.n591 99.5127
R18722 VDD.n1411 VDD.n591 99.5127
R18723 VDD.n1411 VDD.n585 99.5127
R18724 VDD.n1408 VDD.n585 99.5127
R18725 VDD.n1408 VDD.n579 99.5127
R18726 VDD.n1405 VDD.n579 99.5127
R18727 VDD.n1405 VDD.n573 99.5127
R18728 VDD.n1402 VDD.n573 99.5127
R18729 VDD.n1402 VDD.n567 99.5127
R18730 VDD.n1399 VDD.n567 99.5127
R18731 VDD.n1399 VDD.n560 99.5127
R18732 VDD.n1396 VDD.n560 99.5127
R18733 VDD.n1396 VDD.n554 99.5127
R18734 VDD.n1393 VDD.n554 99.5127
R18735 VDD.n1393 VDD.n549 99.5127
R18736 VDD.n1390 VDD.n549 99.5127
R18737 VDD.n1390 VDD.n543 99.5127
R18738 VDD.n1387 VDD.n543 99.5127
R18739 VDD.n1387 VDD.n537 99.5127
R18740 VDD.n1384 VDD.n537 99.5127
R18741 VDD.n1384 VDD.n531 99.5127
R18742 VDD.n1381 VDD.n531 99.5127
R18743 VDD.n1381 VDD.n524 99.5127
R18744 VDD.n1378 VDD.n524 99.5127
R18745 VDD.n1378 VDD.n517 99.5127
R18746 VDD.n517 VDD.n504 99.5127
R18747 VDD.n1802 VDD.n504 99.5127
R18748 VDD.n1802 VDD.n501 99.5127
R18749 VDD.n1508 VDD.n1373 99.5127
R18750 VDD.n1504 VDD.n1503 99.5127
R18751 VDD.n1500 VDD.n1499 99.5127
R18752 VDD.n1496 VDD.n1495 99.5127
R18753 VDD.n1492 VDD.n1491 99.5127
R18754 VDD.n1488 VDD.n1487 99.5127
R18755 VDD.n1484 VDD.n1483 99.5127
R18756 VDD.n1480 VDD.n1479 99.5127
R18757 VDD.n1476 VDD.n1475 99.5127
R18758 VDD.n1472 VDD.n1471 99.5127
R18759 VDD.n1518 VDD.n694 99.5127
R18760 VDD.n1522 VDD.n694 99.5127
R18761 VDD.n1522 VDD.n684 99.5127
R18762 VDD.n1530 VDD.n684 99.5127
R18763 VDD.n1530 VDD.n682 99.5127
R18764 VDD.n1534 VDD.n682 99.5127
R18765 VDD.n1534 VDD.n671 99.5127
R18766 VDD.n1542 VDD.n671 99.5127
R18767 VDD.n1542 VDD.n669 99.5127
R18768 VDD.n1546 VDD.n669 99.5127
R18769 VDD.n1546 VDD.n660 99.5127
R18770 VDD.n1554 VDD.n660 99.5127
R18771 VDD.n1554 VDD.n658 99.5127
R18772 VDD.n1558 VDD.n658 99.5127
R18773 VDD.n1558 VDD.n648 99.5127
R18774 VDD.n1566 VDD.n648 99.5127
R18775 VDD.n1566 VDD.n646 99.5127
R18776 VDD.n1570 VDD.n646 99.5127
R18777 VDD.n1570 VDD.n636 99.5127
R18778 VDD.n1578 VDD.n636 99.5127
R18779 VDD.n1578 VDD.n634 99.5127
R18780 VDD.n1582 VDD.n634 99.5127
R18781 VDD.n1582 VDD.n623 99.5127
R18782 VDD.n1590 VDD.n623 99.5127
R18783 VDD.n1590 VDD.n621 99.5127
R18784 VDD.n1594 VDD.n621 99.5127
R18785 VDD.n1594 VDD.n612 99.5127
R18786 VDD.n1602 VDD.n612 99.5127
R18787 VDD.n1602 VDD.n610 99.5127
R18788 VDD.n1606 VDD.n610 99.5127
R18789 VDD.n1606 VDD.n600 99.5127
R18790 VDD.n1614 VDD.n600 99.5127
R18791 VDD.n1614 VDD.n598 99.5127
R18792 VDD.n1618 VDD.n598 99.5127
R18793 VDD.n1618 VDD.n588 99.5127
R18794 VDD.n1626 VDD.n588 99.5127
R18795 VDD.n1626 VDD.n586 99.5127
R18796 VDD.n1630 VDD.n586 99.5127
R18797 VDD.n1630 VDD.n576 99.5127
R18798 VDD.n1638 VDD.n576 99.5127
R18799 VDD.n1638 VDD.n574 99.5127
R18800 VDD.n1642 VDD.n574 99.5127
R18801 VDD.n1642 VDD.n564 99.5127
R18802 VDD.n1650 VDD.n564 99.5127
R18803 VDD.n1650 VDD.n562 99.5127
R18804 VDD.n1654 VDD.n562 99.5127
R18805 VDD.n1654 VDD.n552 99.5127
R18806 VDD.n1662 VDD.n552 99.5127
R18807 VDD.n1662 VDD.n550 99.5127
R18808 VDD.n1666 VDD.n550 99.5127
R18809 VDD.n1666 VDD.n540 99.5127
R18810 VDD.n1674 VDD.n540 99.5127
R18811 VDD.n1674 VDD.n538 99.5127
R18812 VDD.n1678 VDD.n538 99.5127
R18813 VDD.n1678 VDD.n528 99.5127
R18814 VDD.n1686 VDD.n528 99.5127
R18815 VDD.n1686 VDD.n525 99.5127
R18816 VDD.n1740 VDD.n525 99.5127
R18817 VDD.n1740 VDD.n526 99.5127
R18818 VDD.n526 VDD.n518 99.5127
R18819 VDD.n1735 VDD.n518 99.5127
R18820 VDD.n1735 VDD.n507 99.5127
R18821 VDD.n1732 VDD.n507 99.5127
R18822 VDD.n9 VDD.n8 97.9127
R18823 VDD.n11 VDD.n10 97.9127
R18824 VDD.n13 VDD.n12 97.9127
R18825 VDD.n6 VDD.n5 97.9127
R18826 VDD.n4 VDD.n3 97.9127
R18827 VDD.n2 VDD.n1 97.9127
R18828 VDD.n907 VDD.n906 85.1399
R18829 VDD.n930 VDD.n929 85.1399
R18830 VDD.n2421 VDD.n2420 85.1399
R18831 VDD.n256 VDD.n255 85.1399
R18832 VDD.n104 VDD.n103 85.1399
R18833 VDD.n112 VDD.n111 85.1399
R18834 VDD.n1162 VDD.n1161 85.1399
R18835 VDD.n716 VDD.n715 85.1399
R18836 VDD.n1510 VDD.n1509 72.8958
R18837 VDD.n1510 VDD.n1372 72.8958
R18838 VDD.n1510 VDD.n1371 72.8958
R18839 VDD.n1510 VDD.n1370 72.8958
R18840 VDD.n1510 VDD.n1369 72.8958
R18841 VDD.n1510 VDD.n1368 72.8958
R18842 VDD.n1510 VDD.n1367 72.8958
R18843 VDD.n1510 VDD.n1366 72.8958
R18844 VDD.n1510 VDD.n1365 72.8958
R18845 VDD.n1510 VDD.n1364 72.8958
R18846 VDD.n1510 VDD.n1363 72.8958
R18847 VDD.n1808 VDD.n1807 72.8958
R18848 VDD.n1808 VDD.n499 72.8958
R18849 VDD.n1808 VDD.n498 72.8958
R18850 VDD.n1808 VDD.n497 72.8958
R18851 VDD.n1808 VDD.n496 72.8958
R18852 VDD.n1808 VDD.n495 72.8958
R18853 VDD.n1808 VDD.n494 72.8958
R18854 VDD.n1808 VDD.n493 72.8958
R18855 VDD.n1808 VDD.n492 72.8958
R18856 VDD.n1808 VDD.n491 72.8958
R18857 VDD.n1808 VDD.n490 72.8958
R18858 VDD.n1825 VDD.n1809 72.8958
R18859 VDD.n1830 VDD.n1809 72.8958
R18860 VDD.n1832 VDD.n1809 72.8958
R18861 VDD.n1838 VDD.n1809 72.8958
R18862 VDD.n1840 VDD.n1809 72.8958
R18863 VDD.n1846 VDD.n1809 72.8958
R18864 VDD.n1848 VDD.n1809 72.8958
R18865 VDD.n1854 VDD.n1809 72.8958
R18866 VDD.n1856 VDD.n1809 72.8958
R18867 VDD.n1862 VDD.n1809 72.8958
R18868 VDD.n1864 VDD.n1809 72.8958
R18869 VDD.n2398 VDD.n2397 72.8958
R18870 VDD.n2398 VDD.n279 72.8958
R18871 VDD.n2398 VDD.n278 72.8958
R18872 VDD.n2398 VDD.n277 72.8958
R18873 VDD.n2398 VDD.n276 72.8958
R18874 VDD.n2398 VDD.n275 72.8958
R18875 VDD.n2398 VDD.n274 72.8958
R18876 VDD.n2398 VDD.n273 72.8958
R18877 VDD.n2398 VDD.n272 72.8958
R18878 VDD.n2398 VDD.n271 72.8958
R18879 VDD.n2398 VDD.n270 72.8958
R18880 VDD.n1511 VDD.n1510 72.8958
R18881 VDD.n1510 VDD.n1224 72.8958
R18882 VDD.n1510 VDD.n1225 72.8958
R18883 VDD.n1510 VDD.n1226 72.8958
R18884 VDD.n1510 VDD.n1227 72.8958
R18885 VDD.n1510 VDD.n1228 72.8958
R18886 VDD.n1510 VDD.n1229 72.8958
R18887 VDD.n1510 VDD.n1230 72.8958
R18888 VDD.n1510 VDD.n1231 72.8958
R18889 VDD.n1510 VDD.n1232 72.8958
R18890 VDD.n1808 VDD.n489 72.8958
R18891 VDD.n1808 VDD.n488 72.8958
R18892 VDD.n1808 VDD.n487 72.8958
R18893 VDD.n1808 VDD.n486 72.8958
R18894 VDD.n1808 VDD.n485 72.8958
R18895 VDD.n1808 VDD.n484 72.8958
R18896 VDD.n1808 VDD.n483 72.8958
R18897 VDD.n1808 VDD.n482 72.8958
R18898 VDD.n1808 VDD.n481 72.8958
R18899 VDD.n1808 VDD.n480 72.8958
R18900 VDD.n1808 VDD.n479 72.8958
R18901 VDD.n2101 VDD.n1809 72.8958
R18902 VDD.n1961 VDD.n1809 72.8958
R18903 VDD.n2094 VDD.n1809 72.8958
R18904 VDD.n2088 VDD.n1809 72.8958
R18905 VDD.n2086 VDD.n1809 72.8958
R18906 VDD.n2080 VDD.n1809 72.8958
R18907 VDD.n2078 VDD.n1809 72.8958
R18908 VDD.n2072 VDD.n1809 72.8958
R18909 VDD.n2070 VDD.n1809 72.8958
R18910 VDD.n2063 VDD.n1809 72.8958
R18911 VDD.n2398 VDD.n269 72.8958
R18912 VDD.n2398 VDD.n268 72.8958
R18913 VDD.n2398 VDD.n267 72.8958
R18914 VDD.n2398 VDD.n266 72.8958
R18915 VDD.n2398 VDD.n265 72.8958
R18916 VDD.n2398 VDD.n264 72.8958
R18917 VDD.n2398 VDD.n263 72.8958
R18918 VDD.n2398 VDD.n262 72.8958
R18919 VDD.n2398 VDD.n261 72.8958
R18920 VDD.n2398 VDD.n260 72.8958
R18921 VDD.n2398 VDD.n259 72.8958
R18922 VDD.n1971 VDD.n1970 71.952
R18923 VDD.n293 VDD.n292 71.952
R18924 VDD.n1235 VDD.n1234 71.952
R18925 VDD.n512 VDD.n511 71.952
R18926 VDD.n1814 VDD.n1813 71.952
R18927 VDD.n2280 VDD.n2279 71.952
R18928 VDD.n1375 VDD.n1374 71.952
R18929 VDD.n1690 VDD.n1689 71.952
R18930 VDD.n2472 VDD.n2471 66.2847
R18931 VDD.n2472 VDD.n2399 66.2847
R18932 VDD.n2472 VDD.n2400 66.2847
R18933 VDD.n2472 VDD.n2401 66.2847
R18934 VDD.n2472 VDD.n2402 66.2847
R18935 VDD.n2472 VDD.n2403 66.2847
R18936 VDD.n2472 VDD.n2404 66.2847
R18937 VDD.n2472 VDD.n2405 66.2847
R18938 VDD.n2472 VDD.n2406 66.2847
R18939 VDD.n2472 VDD.n2407 66.2847
R18940 VDD.n2623 VDD.n2622 66.2847
R18941 VDD.n2623 VDD.n101 66.2847
R18942 VDD.n2623 VDD.n100 66.2847
R18943 VDD.n2623 VDD.n99 66.2847
R18944 VDD.n2623 VDD.n98 66.2847
R18945 VDD.n2623 VDD.n97 66.2847
R18946 VDD.n2623 VDD.n96 66.2847
R18947 VDD.n2623 VDD.n95 66.2847
R18948 VDD.n2623 VDD.n94 66.2847
R18949 VDD.n2623 VDD.n93 66.2847
R18950 VDD.n2623 VDD.n92 66.2847
R18951 VDD.n1223 VDD.n1222 66.2847
R18952 VDD.n1223 VDD.n712 66.2847
R18953 VDD.n1223 VDD.n711 66.2847
R18954 VDD.n1223 VDD.n710 66.2847
R18955 VDD.n1223 VDD.n709 66.2847
R18956 VDD.n1223 VDD.n708 66.2847
R18957 VDD.n1223 VDD.n707 66.2847
R18958 VDD.n1223 VDD.n706 66.2847
R18959 VDD.n1223 VDD.n705 66.2847
R18960 VDD.n1223 VDD.n704 66.2847
R18961 VDD.n1223 VDD.n703 66.2847
R18962 VDD.n869 VDD.n866 66.2847
R18963 VDD.n875 VDD.n866 66.2847
R18964 VDD.n878 VDD.n866 66.2847
R18965 VDD.n883 VDD.n866 66.2847
R18966 VDD.n927 VDD.n866 66.2847
R18967 VDD.n886 VDD.n866 66.2847
R18968 VDD.n892 VDD.n866 66.2847
R18969 VDD.n897 VDD.n866 66.2847
R18970 VDD.n900 VDD.n866 66.2847
R18971 VDD.n903 VDD.n866 66.2847
R18972 VDD.n122 VDD.n92 52.4337
R18973 VDD.n126 VDD.n93 52.4337
R18974 VDD.n132 VDD.n94 52.4337
R18975 VDD.n136 VDD.n95 52.4337
R18976 VDD.n142 VDD.n96 52.4337
R18977 VDD.n146 VDD.n97 52.4337
R18978 VDD.n152 VDD.n98 52.4337
R18979 VDD.n156 VDD.n99 52.4337
R18980 VDD.n162 VDD.n100 52.4337
R18981 VDD.n165 VDD.n101 52.4337
R18982 VDD.n2622 VDD.n2621 52.4337
R18983 VDD.n2471 VDD.n2470 52.4337
R18984 VDD.n2465 VDD.n2399 52.4337
R18985 VDD.n2462 VDD.n2400 52.4337
R18986 VDD.n2458 VDD.n2401 52.4337
R18987 VDD.n2454 VDD.n2402 52.4337
R18988 VDD.n2450 VDD.n2403 52.4337
R18989 VDD.n2446 VDD.n2404 52.4337
R18990 VDD.n2442 VDD.n2405 52.4337
R18991 VDD.n2438 VDD.n2406 52.4337
R18992 VDD.n2434 VDD.n2407 52.4337
R18993 VDD.n2471 VDD.n2409 52.4337
R18994 VDD.n2463 VDD.n2399 52.4337
R18995 VDD.n2459 VDD.n2400 52.4337
R18996 VDD.n2455 VDD.n2401 52.4337
R18997 VDD.n2451 VDD.n2402 52.4337
R18998 VDD.n2447 VDD.n2403 52.4337
R18999 VDD.n2443 VDD.n2404 52.4337
R19000 VDD.n2439 VDD.n2405 52.4337
R19001 VDD.n2435 VDD.n2406 52.4337
R19002 VDD.n2407 VDD.n258 52.4337
R19003 VDD.n2622 VDD.n102 52.4337
R19004 VDD.n163 VDD.n101 52.4337
R19005 VDD.n157 VDD.n100 52.4337
R19006 VDD.n153 VDD.n99 52.4337
R19007 VDD.n147 VDD.n98 52.4337
R19008 VDD.n143 VDD.n97 52.4337
R19009 VDD.n137 VDD.n96 52.4337
R19010 VDD.n133 VDD.n95 52.4337
R19011 VDD.n127 VDD.n94 52.4337
R19012 VDD.n123 VDD.n93 52.4337
R19013 VDD.n92 VDD.n90 52.4337
R19014 VDD.n1148 VDD.n703 52.4337
R19015 VDD.n1150 VDD.n704 52.4337
R19016 VDD.n1154 VDD.n705 52.4337
R19017 VDD.n1156 VDD.n706 52.4337
R19018 VDD.n1160 VDD.n707 52.4337
R19019 VDD.n1164 VDD.n708 52.4337
R19020 VDD.n1168 VDD.n709 52.4337
R19021 VDD.n1170 VDD.n710 52.4337
R19022 VDD.n1174 VDD.n711 52.4337
R19023 VDD.n1176 VDD.n712 52.4337
R19024 VDD.n1222 VDD.n713 52.4337
R19025 VDD.n1222 VDD.n1221 52.4337
R19026 VDD.n1177 VDD.n712 52.4337
R19027 VDD.n1175 VDD.n711 52.4337
R19028 VDD.n1173 VDD.n710 52.4337
R19029 VDD.n1169 VDD.n709 52.4337
R19030 VDD.n1167 VDD.n708 52.4337
R19031 VDD.n1163 VDD.n707 52.4337
R19032 VDD.n1159 VDD.n706 52.4337
R19033 VDD.n1155 VDD.n705 52.4337
R19034 VDD.n1153 VDD.n704 52.4337
R19035 VDD.n1149 VDD.n703 52.4337
R19036 VDD.n869 VDD.n867 52.4337
R19037 VDD.n875 VDD.n874 52.4337
R19038 VDD.n878 VDD.n877 52.4337
R19039 VDD.n883 VDD.n882 52.4337
R19040 VDD.n928 VDD.n927 52.4337
R19041 VDD.n925 VDD.n886 52.4337
R19042 VDD.n892 VDD.n891 52.4337
R19043 VDD.n897 VDD.n894 52.4337
R19044 VDD.n900 VDD.n899 52.4337
R19045 VDD.n903 VDD.n902 52.4337
R19046 VDD.n870 VDD.n869 52.4337
R19047 VDD.n876 VDD.n875 52.4337
R19048 VDD.n879 VDD.n878 52.4337
R19049 VDD.n884 VDD.n883 52.4337
R19050 VDD.n927 VDD.n926 52.4337
R19051 VDD.n890 VDD.n886 52.4337
R19052 VDD.n893 VDD.n892 52.4337
R19053 VDD.n898 VDD.n897 52.4337
R19054 VDD.n901 VDD.n900 52.4337
R19055 VDD.n904 VDD.n903 52.4337
R19056 VDD.n2384 VDD.n259 39.2114
R19057 VDD.n2380 VDD.n260 39.2114
R19058 VDD.n2376 VDD.n261 39.2114
R19059 VDD.n2372 VDD.n262 39.2114
R19060 VDD.n2368 VDD.n263 39.2114
R19061 VDD.n2364 VDD.n264 39.2114
R19062 VDD.n2360 VDD.n265 39.2114
R19063 VDD.n2356 VDD.n266 39.2114
R19064 VDD.n2352 VDD.n267 39.2114
R19065 VDD.n2348 VDD.n268 39.2114
R19066 VDD.n2344 VDD.n269 39.2114
R19067 VDD.n2101 VDD.n1959 39.2114
R19068 VDD.n2099 VDD.n1961 39.2114
R19069 VDD.n2095 VDD.n2094 39.2114
R19070 VDD.n2088 VDD.n1963 39.2114
R19071 VDD.n2087 VDD.n2086 39.2114
R19072 VDD.n2080 VDD.n1965 39.2114
R19073 VDD.n2079 VDD.n2078 39.2114
R19074 VDD.n2072 VDD.n1967 39.2114
R19075 VDD.n2071 VDD.n2070 39.2114
R19076 VDD.n2063 VDD.n1969 39.2114
R19077 VDD.n1794 VDD.n479 39.2114
R19078 VDD.n1790 VDD.n480 39.2114
R19079 VDD.n1786 VDD.n481 39.2114
R19080 VDD.n1782 VDD.n482 39.2114
R19081 VDD.n1778 VDD.n483 39.2114
R19082 VDD.n1774 VDD.n484 39.2114
R19083 VDD.n1770 VDD.n485 39.2114
R19084 VDD.n1766 VDD.n486 39.2114
R19085 VDD.n1762 VDD.n487 39.2114
R19086 VDD.n1758 VDD.n488 39.2114
R19087 VDD.n1754 VDD.n489 39.2114
R19088 VDD.n1511 VDD.n699 39.2114
R19089 VDD.n1236 VDD.n1224 39.2114
R19090 VDD.n1240 VDD.n1225 39.2114
R19091 VDD.n1244 VDD.n1226 39.2114
R19092 VDD.n1248 VDD.n1227 39.2114
R19093 VDD.n1252 VDD.n1228 39.2114
R19094 VDD.n1256 VDD.n1229 39.2114
R19095 VDD.n1260 VDD.n1230 39.2114
R19096 VDD.n1264 VDD.n1231 39.2114
R19097 VDD.n1268 VDD.n1232 39.2114
R19098 VDD.n2318 VDD.n270 39.2114
R19099 VDD.n2314 VDD.n271 39.2114
R19100 VDD.n2310 VDD.n272 39.2114
R19101 VDD.n2306 VDD.n273 39.2114
R19102 VDD.n2302 VDD.n274 39.2114
R19103 VDD.n2298 VDD.n275 39.2114
R19104 VDD.n2294 VDD.n276 39.2114
R19105 VDD.n2290 VDD.n277 39.2114
R19106 VDD.n2286 VDD.n278 39.2114
R19107 VDD.n2282 VDD.n279 39.2114
R19108 VDD.n2397 VDD.n2396 39.2114
R19109 VDD.n1825 VDD.n477 39.2114
R19110 VDD.n1830 VDD.n1829 39.2114
R19111 VDD.n1833 VDD.n1832 39.2114
R19112 VDD.n1838 VDD.n1837 39.2114
R19113 VDD.n1841 VDD.n1840 39.2114
R19114 VDD.n1846 VDD.n1845 39.2114
R19115 VDD.n1849 VDD.n1848 39.2114
R19116 VDD.n1854 VDD.n1853 39.2114
R19117 VDD.n1857 VDD.n1856 39.2114
R19118 VDD.n1862 VDD.n1861 39.2114
R19119 VDD.n1865 VDD.n1864 39.2114
R19120 VDD.n1728 VDD.n490 39.2114
R19121 VDD.n1724 VDD.n491 39.2114
R19122 VDD.n1720 VDD.n492 39.2114
R19123 VDD.n1716 VDD.n493 39.2114
R19124 VDD.n1712 VDD.n494 39.2114
R19125 VDD.n1708 VDD.n495 39.2114
R19126 VDD.n1704 VDD.n496 39.2114
R19127 VDD.n1700 VDD.n497 39.2114
R19128 VDD.n1696 VDD.n498 39.2114
R19129 VDD.n1692 VDD.n499 39.2114
R19130 VDD.n1807 VDD.n1806 39.2114
R19131 VDD.n1509 VDD.n696 39.2114
R19132 VDD.n1373 VDD.n1372 39.2114
R19133 VDD.n1503 VDD.n1371 39.2114
R19134 VDD.n1499 VDD.n1370 39.2114
R19135 VDD.n1495 VDD.n1369 39.2114
R19136 VDD.n1491 VDD.n1368 39.2114
R19137 VDD.n1487 VDD.n1367 39.2114
R19138 VDD.n1483 VDD.n1366 39.2114
R19139 VDD.n1479 VDD.n1365 39.2114
R19140 VDD.n1475 VDD.n1364 39.2114
R19141 VDD.n1471 VDD.n1363 39.2114
R19142 VDD.n1509 VDD.n1508 39.2114
R19143 VDD.n1504 VDD.n1372 39.2114
R19144 VDD.n1500 VDD.n1371 39.2114
R19145 VDD.n1496 VDD.n1370 39.2114
R19146 VDD.n1492 VDD.n1369 39.2114
R19147 VDD.n1488 VDD.n1368 39.2114
R19148 VDD.n1484 VDD.n1367 39.2114
R19149 VDD.n1480 VDD.n1366 39.2114
R19150 VDD.n1476 VDD.n1365 39.2114
R19151 VDD.n1472 VDD.n1364 39.2114
R19152 VDD.n1468 VDD.n1363 39.2114
R19153 VDD.n1807 VDD.n500 39.2114
R19154 VDD.n1695 VDD.n499 39.2114
R19155 VDD.n1699 VDD.n498 39.2114
R19156 VDD.n1703 VDD.n497 39.2114
R19157 VDD.n1707 VDD.n496 39.2114
R19158 VDD.n1711 VDD.n495 39.2114
R19159 VDD.n1715 VDD.n494 39.2114
R19160 VDD.n1719 VDD.n493 39.2114
R19161 VDD.n1723 VDD.n492 39.2114
R19162 VDD.n1727 VDD.n491 39.2114
R19163 VDD.n1731 VDD.n490 39.2114
R19164 VDD.n1826 VDD.n1825 39.2114
R19165 VDD.n1831 VDD.n1830 39.2114
R19166 VDD.n1832 VDD.n1823 39.2114
R19167 VDD.n1839 VDD.n1838 39.2114
R19168 VDD.n1840 VDD.n1821 39.2114
R19169 VDD.n1847 VDD.n1846 39.2114
R19170 VDD.n1848 VDD.n1819 39.2114
R19171 VDD.n1855 VDD.n1854 39.2114
R19172 VDD.n1856 VDD.n1817 39.2114
R19173 VDD.n1863 VDD.n1862 39.2114
R19174 VDD.n1864 VDD.n1811 39.2114
R19175 VDD.n2397 VDD.n280 39.2114
R19176 VDD.n2285 VDD.n279 39.2114
R19177 VDD.n2289 VDD.n278 39.2114
R19178 VDD.n2293 VDD.n277 39.2114
R19179 VDD.n2297 VDD.n276 39.2114
R19180 VDD.n2301 VDD.n275 39.2114
R19181 VDD.n2305 VDD.n274 39.2114
R19182 VDD.n2309 VDD.n273 39.2114
R19183 VDD.n2313 VDD.n272 39.2114
R19184 VDD.n2317 VDD.n271 39.2114
R19185 VDD.n2321 VDD.n270 39.2114
R19186 VDD.n1512 VDD.n1511 39.2114
R19187 VDD.n1239 VDD.n1224 39.2114
R19188 VDD.n1243 VDD.n1225 39.2114
R19189 VDD.n1247 VDD.n1226 39.2114
R19190 VDD.n1251 VDD.n1227 39.2114
R19191 VDD.n1255 VDD.n1228 39.2114
R19192 VDD.n1259 VDD.n1229 39.2114
R19193 VDD.n1263 VDD.n1230 39.2114
R19194 VDD.n1267 VDD.n1231 39.2114
R19195 VDD.n1233 VDD.n1232 39.2114
R19196 VDD.n1757 VDD.n489 39.2114
R19197 VDD.n1761 VDD.n488 39.2114
R19198 VDD.n1765 VDD.n487 39.2114
R19199 VDD.n1769 VDD.n486 39.2114
R19200 VDD.n1773 VDD.n485 39.2114
R19201 VDD.n1777 VDD.n484 39.2114
R19202 VDD.n1781 VDD.n483 39.2114
R19203 VDD.n1785 VDD.n482 39.2114
R19204 VDD.n1789 VDD.n481 39.2114
R19205 VDD.n1793 VDD.n480 39.2114
R19206 VDD.n1796 VDD.n479 39.2114
R19207 VDD.n2102 VDD.n2101 39.2114
R19208 VDD.n2096 VDD.n1961 39.2114
R19209 VDD.n2094 VDD.n2093 39.2114
R19210 VDD.n2089 VDD.n2088 39.2114
R19211 VDD.n2086 VDD.n2085 39.2114
R19212 VDD.n2081 VDD.n2080 39.2114
R19213 VDD.n2078 VDD.n2077 39.2114
R19214 VDD.n2073 VDD.n2072 39.2114
R19215 VDD.n2070 VDD.n2069 39.2114
R19216 VDD.n2064 VDD.n2063 39.2114
R19217 VDD.n2347 VDD.n269 39.2114
R19218 VDD.n2351 VDD.n268 39.2114
R19219 VDD.n2355 VDD.n267 39.2114
R19220 VDD.n2359 VDD.n266 39.2114
R19221 VDD.n2363 VDD.n265 39.2114
R19222 VDD.n2367 VDD.n264 39.2114
R19223 VDD.n2371 VDD.n263 39.2114
R19224 VDD.n2375 VDD.n262 39.2114
R19225 VDD.n2379 VDD.n261 39.2114
R19226 VDD.n2383 VDD.n260 39.2114
R19227 VDD.n2386 VDD.n259 39.2114
R19228 VDD.n908 VDD.n907 37.2369
R19229 VDD.n931 VDD.n930 37.2369
R19230 VDD.n2453 VDD.n2421 37.2369
R19231 VDD.n257 VDD.n256 37.2369
R19232 VDD.n105 VDD.n104 37.2369
R19233 VDD.n113 VDD.n112 37.2369
R19234 VDD.n1195 VDD.n1162 37.2369
R19235 VDD.n717 VDD.n716 37.2369
R19236 VDD.n2105 VDD.n2104 34.1859
R19237 VDD.n2388 VDD.n2387 34.1859
R19238 VDD.n2345 VDD.n2342 34.1859
R19239 VDD.n2061 VDD.n2060 34.1859
R19240 VDD.n1798 VDD.n1797 34.1859
R19241 VDD.n1755 VDD.n1752 34.1859
R19242 VDD.n1361 VDD.n1360 34.1859
R19243 VDD.n1515 VDD.n1514 34.1859
R19244 VDD.n2323 VDD.n2320 34.1859
R19245 VDD.n2395 VDD.n2394 34.1859
R19246 VDD.n1957 VDD.n1867 34.1859
R19247 VDD.n2109 VDD.n476 34.1859
R19248 VDD.n1733 VDD.n1730 34.1859
R19249 VDD.n1805 VDD.n1804 34.1859
R19250 VDD.n1469 VDD.n1467 34.1859
R19251 VDD.n1519 VDD.n695 34.1859
R19252 VDD.n2066 VDD.n1971 30.449
R19253 VDD.n294 VDD.n293 30.449
R19254 VDD.n1270 VDD.n1235 30.449
R19255 VDD.n513 VDD.n512 30.449
R19256 VDD.n1815 VDD.n1814 30.449
R19257 VDD.n2281 VDD.n2280 30.449
R19258 VDD.n1376 VDD.n1375 30.449
R19259 VDD.n1691 VDD.n1690 30.449
R19260 VDD.n949 VDD.n866 26.3705
R19261 VDD.n1223 VDD.n702 26.3705
R19262 VDD.n2472 VDD.n251 26.3705
R19263 VDD.n2624 VDD.n2623 26.3705
R19264 VDD.n1808 VDD.n478 21.9471
R19265 VDD.n2107 VDD.n1809 21.9471
R19266 VDD.n1517 VDD.t105 19.9056
R19267 VDD.n287 VDD.t12 19.9056
R19268 VDD.n924 VDD.n885 19.3944
R19269 VDD.n924 VDD.n887 19.3944
R19270 VDD.n920 VDD.n887 19.3944
R19271 VDD.n920 VDD.n919 19.3944
R19272 VDD.n919 VDD.n918 19.3944
R19273 VDD.n918 VDD.n895 19.3944
R19274 VDD.n914 VDD.n895 19.3944
R19275 VDD.n914 VDD.n913 19.3944
R19276 VDD.n913 VDD.n912 19.3944
R19277 VDD.n912 VDD.n909 19.3944
R19278 VDD.n944 VDD.n943 19.3944
R19279 VDD.n943 VDD.n942 19.3944
R19280 VDD.n942 VDD.n872 19.3944
R19281 VDD.n938 VDD.n872 19.3944
R19282 VDD.n938 VDD.n937 19.3944
R19283 VDD.n937 VDD.n936 19.3944
R19284 VDD.n936 VDD.n880 19.3944
R19285 VDD.n932 VDD.n880 19.3944
R19286 VDD.n951 VDD.n863 19.3944
R19287 VDD.n955 VDD.n863 19.3944
R19288 VDD.n955 VDD.n853 19.3944
R19289 VDD.n967 VDD.n853 19.3944
R19290 VDD.n967 VDD.n851 19.3944
R19291 VDD.n971 VDD.n851 19.3944
R19292 VDD.n971 VDD.n841 19.3944
R19293 VDD.n983 VDD.n841 19.3944
R19294 VDD.n983 VDD.n839 19.3944
R19295 VDD.n987 VDD.n839 19.3944
R19296 VDD.n987 VDD.n829 19.3944
R19297 VDD.n999 VDD.n829 19.3944
R19298 VDD.n999 VDD.n827 19.3944
R19299 VDD.n1003 VDD.n827 19.3944
R19300 VDD.n1003 VDD.n818 19.3944
R19301 VDD.n1016 VDD.n818 19.3944
R19302 VDD.n1016 VDD.n816 19.3944
R19303 VDD.n1020 VDD.n816 19.3944
R19304 VDD.n1020 VDD.n806 19.3944
R19305 VDD.n1032 VDD.n806 19.3944
R19306 VDD.n1032 VDD.n804 19.3944
R19307 VDD.n1036 VDD.n804 19.3944
R19308 VDD.n1036 VDD.n794 19.3944
R19309 VDD.n1055 VDD.n794 19.3944
R19310 VDD.n1055 VDD.n792 19.3944
R19311 VDD.n1059 VDD.n792 19.3944
R19312 VDD.n1059 VDD.n782 19.3944
R19313 VDD.n1071 VDD.n782 19.3944
R19314 VDD.n1071 VDD.n780 19.3944
R19315 VDD.n1075 VDD.n780 19.3944
R19316 VDD.n1075 VDD.n769 19.3944
R19317 VDD.n1087 VDD.n769 19.3944
R19318 VDD.n1087 VDD.n767 19.3944
R19319 VDD.n1091 VDD.n767 19.3944
R19320 VDD.n1091 VDD.n758 19.3944
R19321 VDD.n1103 VDD.n758 19.3944
R19322 VDD.n1103 VDD.n756 19.3944
R19323 VDD.n1107 VDD.n756 19.3944
R19324 VDD.n1107 VDD.n746 19.3944
R19325 VDD.n1119 VDD.n746 19.3944
R19326 VDD.n1119 VDD.n744 19.3944
R19327 VDD.n1123 VDD.n744 19.3944
R19328 VDD.n1123 VDD.n734 19.3944
R19329 VDD.n1135 VDD.n734 19.3944
R19330 VDD.n1135 VDD.n732 19.3944
R19331 VDD.n1140 VDD.n732 19.3944
R19332 VDD.n1140 VDD.n720 19.3944
R19333 VDD.n1216 VDD.n720 19.3944
R19334 VDD.n1217 VDD.n1216 19.3944
R19335 VDD.n2469 VDD.n2468 19.3944
R19336 VDD.n2468 VDD.n2467 19.3944
R19337 VDD.n2467 VDD.n2466 19.3944
R19338 VDD.n2466 VDD.n2464 19.3944
R19339 VDD.n2464 VDD.n2461 19.3944
R19340 VDD.n2461 VDD.n2460 19.3944
R19341 VDD.n2460 VDD.n2457 19.3944
R19342 VDD.n2457 VDD.n2456 19.3944
R19343 VDD.n2452 VDD.n2449 19.3944
R19344 VDD.n2449 VDD.n2448 19.3944
R19345 VDD.n2448 VDD.n2445 19.3944
R19346 VDD.n2445 VDD.n2444 19.3944
R19347 VDD.n2444 VDD.n2441 19.3944
R19348 VDD.n2441 VDD.n2440 19.3944
R19349 VDD.n2440 VDD.n2437 19.3944
R19350 VDD.n2437 VDD.n2436 19.3944
R19351 VDD.n2436 VDD.n2433 19.3944
R19352 VDD.n2433 VDD.n2432 19.3944
R19353 VDD.n2478 VDD.n253 19.3944
R19354 VDD.n2478 VDD.n242 19.3944
R19355 VDD.n2490 VDD.n242 19.3944
R19356 VDD.n2490 VDD.n240 19.3944
R19357 VDD.n2494 VDD.n240 19.3944
R19358 VDD.n2494 VDD.n231 19.3944
R19359 VDD.n2506 VDD.n231 19.3944
R19360 VDD.n2506 VDD.n229 19.3944
R19361 VDD.n2510 VDD.n229 19.3944
R19362 VDD.n2510 VDD.n219 19.3944
R19363 VDD.n2522 VDD.n219 19.3944
R19364 VDD.n2522 VDD.n217 19.3944
R19365 VDD.n2526 VDD.n217 19.3944
R19366 VDD.n2526 VDD.n207 19.3944
R19367 VDD.n2538 VDD.n207 19.3944
R19368 VDD.n2538 VDD.n205 19.3944
R19369 VDD.n2542 VDD.n205 19.3944
R19370 VDD.n2542 VDD.n195 19.3944
R19371 VDD.n2554 VDD.n195 19.3944
R19372 VDD.n2554 VDD.n193 19.3944
R19373 VDD.n2561 VDD.n193 19.3944
R19374 VDD.n2561 VDD.n2560 19.3944
R19375 VDD.n2560 VDD.n182 19.3944
R19376 VDD.n2574 VDD.n182 19.3944
R19377 VDD.n2575 VDD.n2574 19.3944
R19378 VDD.n2575 VDD.n180 19.3944
R19379 VDD.n2579 VDD.n180 19.3944
R19380 VDD.n2581 VDD.n2579 19.3944
R19381 VDD.n2582 VDD.n2581 19.3944
R19382 VDD.n2582 VDD.n178 19.3944
R19383 VDD.n2586 VDD.n178 19.3944
R19384 VDD.n2588 VDD.n2586 19.3944
R19385 VDD.n2589 VDD.n2588 19.3944
R19386 VDD.n2589 VDD.n176 19.3944
R19387 VDD.n2593 VDD.n176 19.3944
R19388 VDD.n2595 VDD.n2593 19.3944
R19389 VDD.n2596 VDD.n2595 19.3944
R19390 VDD.n2596 VDD.n174 19.3944
R19391 VDD.n2600 VDD.n174 19.3944
R19392 VDD.n2602 VDD.n2600 19.3944
R19393 VDD.n2603 VDD.n2602 19.3944
R19394 VDD.n2603 VDD.n172 19.3944
R19395 VDD.n2607 VDD.n172 19.3944
R19396 VDD.n2609 VDD.n2607 19.3944
R19397 VDD.n2610 VDD.n2609 19.3944
R19398 VDD.n2610 VDD.n170 19.3944
R19399 VDD.n2614 VDD.n170 19.3944
R19400 VDD.n2616 VDD.n2614 19.3944
R19401 VDD.n2617 VDD.n2616 19.3944
R19402 VDD.n145 VDD.n144 19.3944
R19403 VDD.n148 VDD.n145 19.3944
R19404 VDD.n148 VDD.n109 19.3944
R19405 VDD.n154 VDD.n109 19.3944
R19406 VDD.n155 VDD.n154 19.3944
R19407 VDD.n158 VDD.n155 19.3944
R19408 VDD.n158 VDD.n107 19.3944
R19409 VDD.n164 VDD.n107 19.3944
R19410 VDD.n166 VDD.n164 19.3944
R19411 VDD.n167 VDD.n166 19.3944
R19412 VDD.n118 VDD.n117 19.3944
R19413 VDD.n124 VDD.n117 19.3944
R19414 VDD.n125 VDD.n124 19.3944
R19415 VDD.n128 VDD.n125 19.3944
R19416 VDD.n128 VDD.n115 19.3944
R19417 VDD.n134 VDD.n115 19.3944
R19418 VDD.n135 VDD.n134 19.3944
R19419 VDD.n138 VDD.n135 19.3944
R19420 VDD.n2482 VDD.n249 19.3944
R19421 VDD.n2482 VDD.n247 19.3944
R19422 VDD.n2486 VDD.n247 19.3944
R19423 VDD.n2486 VDD.n237 19.3944
R19424 VDD.n2498 VDD.n237 19.3944
R19425 VDD.n2498 VDD.n235 19.3944
R19426 VDD.n2502 VDD.n235 19.3944
R19427 VDD.n2502 VDD.n225 19.3944
R19428 VDD.n2514 VDD.n225 19.3944
R19429 VDD.n2514 VDD.n223 19.3944
R19430 VDD.n2518 VDD.n223 19.3944
R19431 VDD.n2518 VDD.n213 19.3944
R19432 VDD.n2530 VDD.n213 19.3944
R19433 VDD.n2530 VDD.n211 19.3944
R19434 VDD.n2534 VDD.n211 19.3944
R19435 VDD.n2534 VDD.n201 19.3944
R19436 VDD.n2546 VDD.n201 19.3944
R19437 VDD.n2546 VDD.n199 19.3944
R19438 VDD.n2550 VDD.n199 19.3944
R19439 VDD.n2550 VDD.n188 19.3944
R19440 VDD.n2565 VDD.n188 19.3944
R19441 VDD.n2565 VDD.n186 19.3944
R19442 VDD.n2569 VDD.n186 19.3944
R19443 VDD.n2569 VDD.n23 19.3944
R19444 VDD.n2674 VDD.n23 19.3944
R19445 VDD.n2674 VDD.n24 19.3944
R19446 VDD.n2668 VDD.n24 19.3944
R19447 VDD.n2668 VDD.n2667 19.3944
R19448 VDD.n2667 VDD.n2666 19.3944
R19449 VDD.n2666 VDD.n35 19.3944
R19450 VDD.n2660 VDD.n35 19.3944
R19451 VDD.n2660 VDD.n2659 19.3944
R19452 VDD.n2659 VDD.n2658 19.3944
R19453 VDD.n2658 VDD.n46 19.3944
R19454 VDD.n2652 VDD.n46 19.3944
R19455 VDD.n2652 VDD.n2651 19.3944
R19456 VDD.n2651 VDD.n2650 19.3944
R19457 VDD.n2650 VDD.n57 19.3944
R19458 VDD.n2644 VDD.n57 19.3944
R19459 VDD.n2644 VDD.n2643 19.3944
R19460 VDD.n2643 VDD.n2642 19.3944
R19461 VDD.n2642 VDD.n68 19.3944
R19462 VDD.n2636 VDD.n68 19.3944
R19463 VDD.n2636 VDD.n2635 19.3944
R19464 VDD.n2635 VDD.n2634 19.3944
R19465 VDD.n2634 VDD.n79 19.3944
R19466 VDD.n2628 VDD.n79 19.3944
R19467 VDD.n2628 VDD.n2627 19.3944
R19468 VDD.n2627 VDD.n2626 19.3944
R19469 VDD.n1208 VDD.n1207 19.3944
R19470 VDD.n1207 VDD.n1206 19.3944
R19471 VDD.n1206 VDD.n1151 19.3944
R19472 VDD.n1202 VDD.n1151 19.3944
R19473 VDD.n1202 VDD.n1201 19.3944
R19474 VDD.n1201 VDD.n1200 19.3944
R19475 VDD.n1200 VDD.n1157 19.3944
R19476 VDD.n1196 VDD.n1157 19.3944
R19477 VDD.n1194 VDD.n1165 19.3944
R19478 VDD.n1190 VDD.n1165 19.3944
R19479 VDD.n1190 VDD.n1189 19.3944
R19480 VDD.n1189 VDD.n1188 19.3944
R19481 VDD.n1188 VDD.n1171 19.3944
R19482 VDD.n1184 VDD.n1171 19.3944
R19483 VDD.n1184 VDD.n1183 19.3944
R19484 VDD.n1183 VDD.n1182 19.3944
R19485 VDD.n1182 VDD.n1179 19.3944
R19486 VDD.n1179 VDD.n1178 19.3944
R19487 VDD.n947 VDD.n859 19.3944
R19488 VDD.n959 VDD.n859 19.3944
R19489 VDD.n959 VDD.n857 19.3944
R19490 VDD.n963 VDD.n857 19.3944
R19491 VDD.n963 VDD.n847 19.3944
R19492 VDD.n975 VDD.n847 19.3944
R19493 VDD.n975 VDD.n845 19.3944
R19494 VDD.n979 VDD.n845 19.3944
R19495 VDD.n979 VDD.n835 19.3944
R19496 VDD.n991 VDD.n835 19.3944
R19497 VDD.n991 VDD.n833 19.3944
R19498 VDD.n995 VDD.n833 19.3944
R19499 VDD.n995 VDD.n823 19.3944
R19500 VDD.n1008 VDD.n823 19.3944
R19501 VDD.n1008 VDD.n821 19.3944
R19502 VDD.n1012 VDD.n821 19.3944
R19503 VDD.n1012 VDD.n812 19.3944
R19504 VDD.n1024 VDD.n812 19.3944
R19505 VDD.n1024 VDD.n810 19.3944
R19506 VDD.n1028 VDD.n810 19.3944
R19507 VDD.n1028 VDD.n800 19.3944
R19508 VDD.n1040 VDD.n800 19.3944
R19509 VDD.n1040 VDD.n798 19.3944
R19510 VDD.n1051 VDD.n798 19.3944
R19511 VDD.n1051 VDD.n788 19.3944
R19512 VDD.n1063 VDD.n788 19.3944
R19513 VDD.n1063 VDD.n786 19.3944
R19514 VDD.n1067 VDD.n786 19.3944
R19515 VDD.n1067 VDD.n776 19.3944
R19516 VDD.n1079 VDD.n776 19.3944
R19517 VDD.n1079 VDD.n774 19.3944
R19518 VDD.n1083 VDD.n774 19.3944
R19519 VDD.n1083 VDD.n764 19.3944
R19520 VDD.n1095 VDD.n764 19.3944
R19521 VDD.n1095 VDD.n762 19.3944
R19522 VDD.n1099 VDD.n762 19.3944
R19523 VDD.n1099 VDD.n752 19.3944
R19524 VDD.n1111 VDD.n752 19.3944
R19525 VDD.n1111 VDD.n750 19.3944
R19526 VDD.n1115 VDD.n750 19.3944
R19527 VDD.n1115 VDD.n740 19.3944
R19528 VDD.n1127 VDD.n740 19.3944
R19529 VDD.n1127 VDD.n738 19.3944
R19530 VDD.n1131 VDD.n738 19.3944
R19531 VDD.n1131 VDD.n728 19.3944
R19532 VDD.n1144 VDD.n728 19.3944
R19533 VDD.n1144 VDD.n725 19.3944
R19534 VDD.n1212 VDD.n725 19.3944
R19535 VDD.n1212 VDD.n726 19.3944
R19536 VDD.n949 VDD.n861 17.0134
R19537 VDD.n957 VDD.n861 17.0134
R19538 VDD.n957 VDD.n855 17.0134
R19539 VDD.n965 VDD.n855 17.0134
R19540 VDD.n973 VDD.n849 17.0134
R19541 VDD.n973 VDD.n843 17.0134
R19542 VDD.n981 VDD.n843 17.0134
R19543 VDD.n981 VDD.n837 17.0134
R19544 VDD.n989 VDD.n837 17.0134
R19545 VDD.n989 VDD.n831 17.0134
R19546 VDD.n997 VDD.n831 17.0134
R19547 VDD.n997 VDD.n825 17.0134
R19548 VDD.n1006 VDD.n825 17.0134
R19549 VDD.n1006 VDD.n1005 17.0134
R19550 VDD.n1014 VDD.n814 17.0134
R19551 VDD.n1022 VDD.n814 17.0134
R19552 VDD.n1022 VDD.n808 17.0134
R19553 VDD.n1030 VDD.n808 17.0134
R19554 VDD.n1030 VDD.n802 17.0134
R19555 VDD.n1038 VDD.n802 17.0134
R19556 VDD.n1038 VDD.n796 17.0134
R19557 VDD.n1053 VDD.n796 17.0134
R19558 VDD.n1061 VDD.n790 17.0134
R19559 VDD.n1061 VDD.n784 17.0134
R19560 VDD.n1069 VDD.n784 17.0134
R19561 VDD.n1069 VDD.n778 17.0134
R19562 VDD.n1077 VDD.n778 17.0134
R19563 VDD.n1077 VDD.n771 17.0134
R19564 VDD.n1085 VDD.n771 17.0134
R19565 VDD.n1085 VDD.n772 17.0134
R19566 VDD.n1093 VDD.n760 17.0134
R19567 VDD.n1101 VDD.n760 17.0134
R19568 VDD.n1101 VDD.n754 17.0134
R19569 VDD.n1109 VDD.n754 17.0134
R19570 VDD.n1109 VDD.n748 17.0134
R19571 VDD.n1117 VDD.n748 17.0134
R19572 VDD.n1117 VDD.n742 17.0134
R19573 VDD.n1125 VDD.n742 17.0134
R19574 VDD.n1125 VDD.n736 17.0134
R19575 VDD.n1133 VDD.n736 17.0134
R19576 VDD.n1142 VDD.n730 17.0134
R19577 VDD.n1142 VDD.n722 17.0134
R19578 VDD.n1214 VDD.n722 17.0134
R19579 VDD.n1214 VDD.n702 17.0134
R19580 VDD.n2480 VDD.n251 17.0134
R19581 VDD.n2480 VDD.n244 17.0134
R19582 VDD.n2488 VDD.n244 17.0134
R19583 VDD.n2488 VDD.n245 17.0134
R19584 VDD.n2496 VDD.n233 17.0134
R19585 VDD.n2504 VDD.n233 17.0134
R19586 VDD.n2504 VDD.n227 17.0134
R19587 VDD.n2512 VDD.n227 17.0134
R19588 VDD.n2512 VDD.n221 17.0134
R19589 VDD.n2520 VDD.n221 17.0134
R19590 VDD.n2520 VDD.n215 17.0134
R19591 VDD.n2528 VDD.n215 17.0134
R19592 VDD.n2528 VDD.n209 17.0134
R19593 VDD.n2536 VDD.n209 17.0134
R19594 VDD.n2544 VDD.n203 17.0134
R19595 VDD.n2544 VDD.n197 17.0134
R19596 VDD.n2552 VDD.n197 17.0134
R19597 VDD.n2552 VDD.n190 17.0134
R19598 VDD.n2563 VDD.n190 17.0134
R19599 VDD.n2563 VDD.n184 17.0134
R19600 VDD.n2571 VDD.n184 17.0134
R19601 VDD.n2572 VDD.n2571 17.0134
R19602 VDD.n2672 VDD.n2671 17.0134
R19603 VDD.n2671 VDD.n2670 17.0134
R19604 VDD.n2670 VDD.n30 17.0134
R19605 VDD.n2664 VDD.n30 17.0134
R19606 VDD.n2664 VDD.n2663 17.0134
R19607 VDD.n2663 VDD.n2662 17.0134
R19608 VDD.n2662 VDD.n40 17.0134
R19609 VDD.n2656 VDD.n40 17.0134
R19610 VDD.n2655 VDD.n2654 17.0134
R19611 VDD.n2654 VDD.n51 17.0134
R19612 VDD.n2648 VDD.n51 17.0134
R19613 VDD.n2648 VDD.n2647 17.0134
R19614 VDD.n2647 VDD.n2646 17.0134
R19615 VDD.n2646 VDD.n62 17.0134
R19616 VDD.n2640 VDD.n62 17.0134
R19617 VDD.n2640 VDD.n2639 17.0134
R19618 VDD.n2639 VDD.n2638 17.0134
R19619 VDD.n2638 VDD.n73 17.0134
R19620 VDD.n2632 VDD.n2631 17.0134
R19621 VDD.n2631 VDD.n2630 17.0134
R19622 VDD.n2630 VDD.n84 17.0134
R19623 VDD.n2624 VDD.n84 17.0134
R19624 VDD.n931 VDD.n885 15.9035
R19625 VDD.n2453 VDD.n2452 15.9035
R19626 VDD.n144 VDD.n113 15.9035
R19627 VDD.n1195 VDD.n1194 15.9035
R19628 VDD.n965 VDD.t27 12.9303
R19629 VDD.t60 VDD.n730 12.9303
R19630 VDD.n245 VDD.t67 12.9303
R19631 VDD.n2632 VDD.t31 12.9303
R19632 VDD.n1005 VDD.t90 12.2498
R19633 VDD.n1093 VDD.t98 12.2498
R19634 VDD.n2536 VDD.t87 12.2498
R19635 VDD.t96 VDD.n2655 12.2498
R19636 VDD.n1517 VDD.n691 11.5693
R19637 VDD.n1523 VDD.n691 11.5693
R19638 VDD.n1523 VDD.n685 11.5693
R19639 VDD.n1529 VDD.n685 11.5693
R19640 VDD.n1529 VDD.n679 11.5693
R19641 VDD.n1535 VDD.n679 11.5693
R19642 VDD.n1541 VDD.n672 11.5693
R19643 VDD.n1541 VDD.n675 11.5693
R19644 VDD.n1547 VDD.n661 11.5693
R19645 VDD.n1553 VDD.n661 11.5693
R19646 VDD.n1553 VDD.n655 11.5693
R19647 VDD.n1559 VDD.n655 11.5693
R19648 VDD.n1559 VDD.n649 11.5693
R19649 VDD.n1565 VDD.n649 11.5693
R19650 VDD.n1565 VDD.n643 11.5693
R19651 VDD.n1571 VDD.n643 11.5693
R19652 VDD.n1571 VDD.n637 11.5693
R19653 VDD.n1577 VDD.n637 11.5693
R19654 VDD.n1583 VDD.n631 11.5693
R19655 VDD.n1583 VDD.n624 11.5693
R19656 VDD.n1589 VDD.n624 11.5693
R19657 VDD.n1589 VDD.n627 11.5693
R19658 VDD.n1595 VDD.n613 11.5693
R19659 VDD.n1601 VDD.n613 11.5693
R19660 VDD.n1601 VDD.n606 11.5693
R19661 VDD.n1607 VDD.n606 11.5693
R19662 VDD.n1607 VDD.n609 11.5693
R19663 VDD.n1613 VDD.n595 11.5693
R19664 VDD.n1619 VDD.n595 11.5693
R19665 VDD.n1619 VDD.n589 11.5693
R19666 VDD.n1625 VDD.n589 11.5693
R19667 VDD.n1631 VDD.n583 11.5693
R19668 VDD.n1631 VDD.n577 11.5693
R19669 VDD.n1637 VDD.n577 11.5693
R19670 VDD.n1637 VDD.n571 11.5693
R19671 VDD.n1643 VDD.n571 11.5693
R19672 VDD.n1649 VDD.n565 11.5693
R19673 VDD.n1649 VDD.n558 11.5693
R19674 VDD.n1655 VDD.n558 11.5693
R19675 VDD.n1655 VDD.n561 11.5693
R19676 VDD.n1661 VDD.n547 11.5693
R19677 VDD.n1667 VDD.n547 11.5693
R19678 VDD.n1667 VDD.n541 11.5693
R19679 VDD.n1673 VDD.n541 11.5693
R19680 VDD.n1673 VDD.n535 11.5693
R19681 VDD.n1679 VDD.n535 11.5693
R19682 VDD.n1679 VDD.n529 11.5693
R19683 VDD.n1685 VDD.n529 11.5693
R19684 VDD.n1741 VDD.n522 11.5693
R19685 VDD.n1747 VDD.n516 11.5693
R19686 VDD.n1747 VDD.n505 11.5693
R19687 VDD.n1801 VDD.n505 11.5693
R19688 VDD.n1801 VDD.n478 11.5693
R19689 VDD.n2107 VDD.n472 11.5693
R19690 VDD.n2113 VDD.n472 11.5693
R19691 VDD.n2113 VDD.n466 11.5693
R19692 VDD.n2119 VDD.n466 11.5693
R19693 VDD.n2125 VDD.n460 11.5693
R19694 VDD.n2131 VDD.n454 11.5693
R19695 VDD.n2131 VDD.n448 11.5693
R19696 VDD.n2137 VDD.n448 11.5693
R19697 VDD.n2137 VDD.n442 11.5693
R19698 VDD.n2143 VDD.n442 11.5693
R19699 VDD.n2143 VDD.n435 11.5693
R19700 VDD.n2149 VDD.n435 11.5693
R19701 VDD.n2149 VDD.n438 11.5693
R19702 VDD.n2155 VDD.n424 11.5693
R19703 VDD.n2161 VDD.n424 11.5693
R19704 VDD.n2161 VDD.n418 11.5693
R19705 VDD.n2167 VDD.n418 11.5693
R19706 VDD.n2173 VDD.n412 11.5693
R19707 VDD.n2173 VDD.n406 11.5693
R19708 VDD.n2179 VDD.n406 11.5693
R19709 VDD.n2179 VDD.n400 11.5693
R19710 VDD.n2185 VDD.n400 11.5693
R19711 VDD.n2191 VDD.n394 11.5693
R19712 VDD.n2191 VDD.n387 11.5693
R19713 VDD.n2197 VDD.n387 11.5693
R19714 VDD.n2197 VDD.n390 11.5693
R19715 VDD.n2203 VDD.n376 11.5693
R19716 VDD.n2209 VDD.n376 11.5693
R19717 VDD.n2209 VDD.n369 11.5693
R19718 VDD.n2215 VDD.n369 11.5693
R19719 VDD.n2215 VDD.n372 11.5693
R19720 VDD.n2221 VDD.n358 11.5693
R19721 VDD.n2227 VDD.n358 11.5693
R19722 VDD.n2227 VDD.n352 11.5693
R19723 VDD.n2233 VDD.n352 11.5693
R19724 VDD.n2239 VDD.n346 11.5693
R19725 VDD.n2239 VDD.n340 11.5693
R19726 VDD.n2245 VDD.n340 11.5693
R19727 VDD.n2245 VDD.n334 11.5693
R19728 VDD.n2251 VDD.n334 11.5693
R19729 VDD.n2251 VDD.n328 11.5693
R19730 VDD.n2257 VDD.n328 11.5693
R19731 VDD.n2257 VDD.n321 11.5693
R19732 VDD.n2263 VDD.n321 11.5693
R19733 VDD.n2263 VDD.n324 11.5693
R19734 VDD.n2269 VDD.n310 11.5693
R19735 VDD.n2275 VDD.n310 11.5693
R19736 VDD.n2331 VDD.n303 11.5693
R19737 VDD.n2331 VDD.n297 11.5693
R19738 VDD.n2337 VDD.n297 11.5693
R19739 VDD.n2337 VDD.n285 11.5693
R19740 VDD.n2391 VDD.n285 11.5693
R19741 VDD.n2391 VDD.n287 11.5693
R19742 VDD.n2105 VDD.n470 10.6151
R19743 VDD.n2115 VDD.n470 10.6151
R19744 VDD.n2116 VDD.n2115 10.6151
R19745 VDD.n2117 VDD.n2116 10.6151
R19746 VDD.n2117 VDD.n458 10.6151
R19747 VDD.n2127 VDD.n458 10.6151
R19748 VDD.n2128 VDD.n2127 10.6151
R19749 VDD.n2129 VDD.n2128 10.6151
R19750 VDD.n2129 VDD.n446 10.6151
R19751 VDD.n2139 VDD.n446 10.6151
R19752 VDD.n2140 VDD.n2139 10.6151
R19753 VDD.n2141 VDD.n2140 10.6151
R19754 VDD.n2141 VDD.n433 10.6151
R19755 VDD.n2151 VDD.n433 10.6151
R19756 VDD.n2152 VDD.n2151 10.6151
R19757 VDD.n2153 VDD.n2152 10.6151
R19758 VDD.n2153 VDD.n422 10.6151
R19759 VDD.n2163 VDD.n422 10.6151
R19760 VDD.n2164 VDD.n2163 10.6151
R19761 VDD.n2165 VDD.n2164 10.6151
R19762 VDD.n2165 VDD.n410 10.6151
R19763 VDD.n2175 VDD.n410 10.6151
R19764 VDD.n2176 VDD.n2175 10.6151
R19765 VDD.n2177 VDD.n2176 10.6151
R19766 VDD.n2177 VDD.n398 10.6151
R19767 VDD.n2187 VDD.n398 10.6151
R19768 VDD.n2188 VDD.n2187 10.6151
R19769 VDD.n2189 VDD.n2188 10.6151
R19770 VDD.n2189 VDD.n385 10.6151
R19771 VDD.n2199 VDD.n385 10.6151
R19772 VDD.n2200 VDD.n2199 10.6151
R19773 VDD.n2201 VDD.n2200 10.6151
R19774 VDD.n2201 VDD.n374 10.6151
R19775 VDD.n2211 VDD.n374 10.6151
R19776 VDD.n2212 VDD.n2211 10.6151
R19777 VDD.n2213 VDD.n2212 10.6151
R19778 VDD.n2213 VDD.n362 10.6151
R19779 VDD.n2223 VDD.n362 10.6151
R19780 VDD.n2224 VDD.n2223 10.6151
R19781 VDD.n2225 VDD.n2224 10.6151
R19782 VDD.n2225 VDD.n350 10.6151
R19783 VDD.n2235 VDD.n350 10.6151
R19784 VDD.n2236 VDD.n2235 10.6151
R19785 VDD.n2237 VDD.n2236 10.6151
R19786 VDD.n2237 VDD.n338 10.6151
R19787 VDD.n2247 VDD.n338 10.6151
R19788 VDD.n2248 VDD.n2247 10.6151
R19789 VDD.n2249 VDD.n2248 10.6151
R19790 VDD.n2249 VDD.n326 10.6151
R19791 VDD.n2259 VDD.n326 10.6151
R19792 VDD.n2260 VDD.n2259 10.6151
R19793 VDD.n2261 VDD.n2260 10.6151
R19794 VDD.n2261 VDD.n314 10.6151
R19795 VDD.n2271 VDD.n314 10.6151
R19796 VDD.n2272 VDD.n2271 10.6151
R19797 VDD.n2273 VDD.n2272 10.6151
R19798 VDD.n2273 VDD.n301 10.6151
R19799 VDD.n2333 VDD.n301 10.6151
R19800 VDD.n2334 VDD.n2333 10.6151
R19801 VDD.n2335 VDD.n2334 10.6151
R19802 VDD.n2335 VDD.n291 10.6151
R19803 VDD.n2389 VDD.n291 10.6151
R19804 VDD.n2389 VDD.n2388 10.6151
R19805 VDD.n2387 VDD.n2385 10.6151
R19806 VDD.n2385 VDD.n2382 10.6151
R19807 VDD.n2382 VDD.n2381 10.6151
R19808 VDD.n2381 VDD.n2378 10.6151
R19809 VDD.n2378 VDD.n2377 10.6151
R19810 VDD.n2377 VDD.n2374 10.6151
R19811 VDD.n2374 VDD.n2373 10.6151
R19812 VDD.n2373 VDD.n2370 10.6151
R19813 VDD.n2370 VDD.n2369 10.6151
R19814 VDD.n2369 VDD.n2366 10.6151
R19815 VDD.n2366 VDD.n2365 10.6151
R19816 VDD.n2365 VDD.n2362 10.6151
R19817 VDD.n2362 VDD.n2361 10.6151
R19818 VDD.n2361 VDD.n2358 10.6151
R19819 VDD.n2358 VDD.n2357 10.6151
R19820 VDD.n2357 VDD.n2354 10.6151
R19821 VDD.n2354 VDD.n2353 10.6151
R19822 VDD.n2353 VDD.n2350 10.6151
R19823 VDD.n2350 VDD.n2349 10.6151
R19824 VDD.n2346 VDD.n2345 10.6151
R19825 VDD.n2060 VDD.n2059 10.6151
R19826 VDD.n2059 VDD.n2057 10.6151
R19827 VDD.n2057 VDD.n2056 10.6151
R19828 VDD.n2056 VDD.n2054 10.6151
R19829 VDD.n2054 VDD.n2053 10.6151
R19830 VDD.n2053 VDD.n2051 10.6151
R19831 VDD.n2051 VDD.n2050 10.6151
R19832 VDD.n2050 VDD.n2048 10.6151
R19833 VDD.n2048 VDD.n2047 10.6151
R19834 VDD.n2047 VDD.n2045 10.6151
R19835 VDD.n2045 VDD.n2044 10.6151
R19836 VDD.n2044 VDD.n2042 10.6151
R19837 VDD.n2042 VDD.n2041 10.6151
R19838 VDD.n2041 VDD.n2039 10.6151
R19839 VDD.n2039 VDD.n2038 10.6151
R19840 VDD.n2038 VDD.n2036 10.6151
R19841 VDD.n2036 VDD.n2035 10.6151
R19842 VDD.n2035 VDD.n2033 10.6151
R19843 VDD.n2033 VDD.n2032 10.6151
R19844 VDD.n2032 VDD.n2030 10.6151
R19845 VDD.n2030 VDD.n2029 10.6151
R19846 VDD.n2029 VDD.n2027 10.6151
R19847 VDD.n2027 VDD.n2026 10.6151
R19848 VDD.n2026 VDD.n2024 10.6151
R19849 VDD.n2024 VDD.n2023 10.6151
R19850 VDD.n2023 VDD.n2021 10.6151
R19851 VDD.n2021 VDD.n2020 10.6151
R19852 VDD.n2020 VDD.n2018 10.6151
R19853 VDD.n2018 VDD.n2017 10.6151
R19854 VDD.n2017 VDD.n2015 10.6151
R19855 VDD.n2015 VDD.n2014 10.6151
R19856 VDD.n2014 VDD.n2012 10.6151
R19857 VDD.n2012 VDD.n2011 10.6151
R19858 VDD.n2011 VDD.n2009 10.6151
R19859 VDD.n2009 VDD.n2008 10.6151
R19860 VDD.n2008 VDD.n2006 10.6151
R19861 VDD.n2006 VDD.n2005 10.6151
R19862 VDD.n2005 VDD.n2003 10.6151
R19863 VDD.n2003 VDD.n2002 10.6151
R19864 VDD.n2002 VDD.n2000 10.6151
R19865 VDD.n2000 VDD.n1999 10.6151
R19866 VDD.n1999 VDD.n1997 10.6151
R19867 VDD.n1997 VDD.n1996 10.6151
R19868 VDD.n1996 VDD.n1994 10.6151
R19869 VDD.n1994 VDD.n1993 10.6151
R19870 VDD.n1993 VDD.n1991 10.6151
R19871 VDD.n1991 VDD.n1990 10.6151
R19872 VDD.n1990 VDD.n1988 10.6151
R19873 VDD.n1988 VDD.n1987 10.6151
R19874 VDD.n1987 VDD.n1985 10.6151
R19875 VDD.n1985 VDD.n1984 10.6151
R19876 VDD.n1984 VDD.n1982 10.6151
R19877 VDD.n1982 VDD.n1981 10.6151
R19878 VDD.n1981 VDD.n1979 10.6151
R19879 VDD.n1979 VDD.n1978 10.6151
R19880 VDD.n1978 VDD.n1976 10.6151
R19881 VDD.n1976 VDD.n1975 10.6151
R19882 VDD.n1975 VDD.n1973 10.6151
R19883 VDD.n1973 VDD.n1972 10.6151
R19884 VDD.n1972 VDD.n295 10.6151
R19885 VDD.n2340 VDD.n295 10.6151
R19886 VDD.n2341 VDD.n2340 10.6151
R19887 VDD.n2342 VDD.n2341 10.6151
R19888 VDD.n2104 VDD.n2103 10.6151
R19889 VDD.n2103 VDD.n1960 10.6151
R19890 VDD.n2098 VDD.n1960 10.6151
R19891 VDD.n2098 VDD.n2097 10.6151
R19892 VDD.n2097 VDD.n1962 10.6151
R19893 VDD.n2092 VDD.n1962 10.6151
R19894 VDD.n2092 VDD.n2091 10.6151
R19895 VDD.n2091 VDD.n2090 10.6151
R19896 VDD.n2090 VDD.n1964 10.6151
R19897 VDD.n2084 VDD.n1964 10.6151
R19898 VDD.n2084 VDD.n2083 10.6151
R19899 VDD.n2083 VDD.n2082 10.6151
R19900 VDD.n2082 VDD.n1966 10.6151
R19901 VDD.n2076 VDD.n1966 10.6151
R19902 VDD.n2076 VDD.n2075 10.6151
R19903 VDD.n2075 VDD.n2074 10.6151
R19904 VDD.n2074 VDD.n1968 10.6151
R19905 VDD.n2068 VDD.n1968 10.6151
R19906 VDD.n2068 VDD.n2067 10.6151
R19907 VDD.n2065 VDD.n2061 10.6151
R19908 VDD.n1797 VDD.n1795 10.6151
R19909 VDD.n1795 VDD.n1792 10.6151
R19910 VDD.n1792 VDD.n1791 10.6151
R19911 VDD.n1791 VDD.n1788 10.6151
R19912 VDD.n1788 VDD.n1787 10.6151
R19913 VDD.n1787 VDD.n1784 10.6151
R19914 VDD.n1784 VDD.n1783 10.6151
R19915 VDD.n1783 VDD.n1780 10.6151
R19916 VDD.n1780 VDD.n1779 10.6151
R19917 VDD.n1779 VDD.n1776 10.6151
R19918 VDD.n1776 VDD.n1775 10.6151
R19919 VDD.n1775 VDD.n1772 10.6151
R19920 VDD.n1772 VDD.n1771 10.6151
R19921 VDD.n1771 VDD.n1768 10.6151
R19922 VDD.n1768 VDD.n1767 10.6151
R19923 VDD.n1767 VDD.n1764 10.6151
R19924 VDD.n1764 VDD.n1763 10.6151
R19925 VDD.n1763 VDD.n1760 10.6151
R19926 VDD.n1760 VDD.n1759 10.6151
R19927 VDD.n1756 VDD.n1755 10.6151
R19928 VDD.n1360 VDD.n1359 10.6151
R19929 VDD.n1359 VDD.n1357 10.6151
R19930 VDD.n1357 VDD.n1356 10.6151
R19931 VDD.n1356 VDD.n1354 10.6151
R19932 VDD.n1354 VDD.n1353 10.6151
R19933 VDD.n1353 VDD.n1351 10.6151
R19934 VDD.n1351 VDD.n1350 10.6151
R19935 VDD.n1350 VDD.n1348 10.6151
R19936 VDD.n1348 VDD.n1347 10.6151
R19937 VDD.n1347 VDD.n1345 10.6151
R19938 VDD.n1345 VDD.n1344 10.6151
R19939 VDD.n1344 VDD.n1342 10.6151
R19940 VDD.n1342 VDD.n1341 10.6151
R19941 VDD.n1341 VDD.n1339 10.6151
R19942 VDD.n1339 VDD.n1338 10.6151
R19943 VDD.n1338 VDD.n1336 10.6151
R19944 VDD.n1336 VDD.n1335 10.6151
R19945 VDD.n1335 VDD.n1333 10.6151
R19946 VDD.n1333 VDD.n1332 10.6151
R19947 VDD.n1332 VDD.n1330 10.6151
R19948 VDD.n1330 VDD.n1329 10.6151
R19949 VDD.n1329 VDD.n1327 10.6151
R19950 VDD.n1327 VDD.n1326 10.6151
R19951 VDD.n1326 VDD.n1324 10.6151
R19952 VDD.n1324 VDD.n1323 10.6151
R19953 VDD.n1323 VDD.n1321 10.6151
R19954 VDD.n1321 VDD.n1320 10.6151
R19955 VDD.n1320 VDD.n1318 10.6151
R19956 VDD.n1318 VDD.n1317 10.6151
R19957 VDD.n1317 VDD.n1315 10.6151
R19958 VDD.n1315 VDD.n1314 10.6151
R19959 VDD.n1314 VDD.n1312 10.6151
R19960 VDD.n1312 VDD.n1311 10.6151
R19961 VDD.n1311 VDD.n1309 10.6151
R19962 VDD.n1309 VDD.n1308 10.6151
R19963 VDD.n1308 VDD.n1306 10.6151
R19964 VDD.n1306 VDD.n1305 10.6151
R19965 VDD.n1305 VDD.n1303 10.6151
R19966 VDD.n1303 VDD.n1302 10.6151
R19967 VDD.n1302 VDD.n1300 10.6151
R19968 VDD.n1300 VDD.n1299 10.6151
R19969 VDD.n1299 VDD.n1297 10.6151
R19970 VDD.n1297 VDD.n1296 10.6151
R19971 VDD.n1296 VDD.n1294 10.6151
R19972 VDD.n1294 VDD.n1293 10.6151
R19973 VDD.n1293 VDD.n1291 10.6151
R19974 VDD.n1291 VDD.n1290 10.6151
R19975 VDD.n1290 VDD.n1288 10.6151
R19976 VDD.n1288 VDD.n1287 10.6151
R19977 VDD.n1287 VDD.n1285 10.6151
R19978 VDD.n1285 VDD.n1284 10.6151
R19979 VDD.n1284 VDD.n1282 10.6151
R19980 VDD.n1282 VDD.n1281 10.6151
R19981 VDD.n1281 VDD.n1279 10.6151
R19982 VDD.n1279 VDD.n1278 10.6151
R19983 VDD.n1278 VDD.n1276 10.6151
R19984 VDD.n1276 VDD.n1275 10.6151
R19985 VDD.n1275 VDD.n1273 10.6151
R19986 VDD.n1273 VDD.n1272 10.6151
R19987 VDD.n1272 VDD.n514 10.6151
R19988 VDD.n1750 VDD.n514 10.6151
R19989 VDD.n1751 VDD.n1750 10.6151
R19990 VDD.n1752 VDD.n1751 10.6151
R19991 VDD.n1514 VDD.n1513 10.6151
R19992 VDD.n1513 VDD.n700 10.6151
R19993 VDD.n1237 VDD.n700 10.6151
R19994 VDD.n1238 VDD.n1237 10.6151
R19995 VDD.n1241 VDD.n1238 10.6151
R19996 VDD.n1242 VDD.n1241 10.6151
R19997 VDD.n1245 VDD.n1242 10.6151
R19998 VDD.n1246 VDD.n1245 10.6151
R19999 VDD.n1249 VDD.n1246 10.6151
R20000 VDD.n1250 VDD.n1249 10.6151
R20001 VDD.n1253 VDD.n1250 10.6151
R20002 VDD.n1254 VDD.n1253 10.6151
R20003 VDD.n1257 VDD.n1254 10.6151
R20004 VDD.n1258 VDD.n1257 10.6151
R20005 VDD.n1261 VDD.n1258 10.6151
R20006 VDD.n1262 VDD.n1261 10.6151
R20007 VDD.n1265 VDD.n1262 10.6151
R20008 VDD.n1266 VDD.n1265 10.6151
R20009 VDD.n1269 VDD.n1266 10.6151
R20010 VDD.n1361 VDD.n1271 10.6151
R20011 VDD.n1515 VDD.n689 10.6151
R20012 VDD.n1525 VDD.n689 10.6151
R20013 VDD.n1526 VDD.n1525 10.6151
R20014 VDD.n1527 VDD.n1526 10.6151
R20015 VDD.n1527 VDD.n677 10.6151
R20016 VDD.n1537 VDD.n677 10.6151
R20017 VDD.n1538 VDD.n1537 10.6151
R20018 VDD.n1539 VDD.n1538 10.6151
R20019 VDD.n1539 VDD.n665 10.6151
R20020 VDD.n1549 VDD.n665 10.6151
R20021 VDD.n1550 VDD.n1549 10.6151
R20022 VDD.n1551 VDD.n1550 10.6151
R20023 VDD.n1551 VDD.n653 10.6151
R20024 VDD.n1561 VDD.n653 10.6151
R20025 VDD.n1562 VDD.n1561 10.6151
R20026 VDD.n1563 VDD.n1562 10.6151
R20027 VDD.n1563 VDD.n641 10.6151
R20028 VDD.n1573 VDD.n641 10.6151
R20029 VDD.n1574 VDD.n1573 10.6151
R20030 VDD.n1575 VDD.n1574 10.6151
R20031 VDD.n1575 VDD.n629 10.6151
R20032 VDD.n1585 VDD.n629 10.6151
R20033 VDD.n1586 VDD.n1585 10.6151
R20034 VDD.n1587 VDD.n1586 10.6151
R20035 VDD.n1587 VDD.n617 10.6151
R20036 VDD.n1597 VDD.n617 10.6151
R20037 VDD.n1598 VDD.n1597 10.6151
R20038 VDD.n1599 VDD.n1598 10.6151
R20039 VDD.n1599 VDD.n604 10.6151
R20040 VDD.n1609 VDD.n604 10.6151
R20041 VDD.n1610 VDD.n1609 10.6151
R20042 VDD.n1611 VDD.n1610 10.6151
R20043 VDD.n1611 VDD.n593 10.6151
R20044 VDD.n1621 VDD.n593 10.6151
R20045 VDD.n1622 VDD.n1621 10.6151
R20046 VDD.n1623 VDD.n1622 10.6151
R20047 VDD.n1623 VDD.n581 10.6151
R20048 VDD.n1633 VDD.n581 10.6151
R20049 VDD.n1634 VDD.n1633 10.6151
R20050 VDD.n1635 VDD.n1634 10.6151
R20051 VDD.n1635 VDD.n569 10.6151
R20052 VDD.n1645 VDD.n569 10.6151
R20053 VDD.n1646 VDD.n1645 10.6151
R20054 VDD.n1647 VDD.n1646 10.6151
R20055 VDD.n1647 VDD.n556 10.6151
R20056 VDD.n1657 VDD.n556 10.6151
R20057 VDD.n1658 VDD.n1657 10.6151
R20058 VDD.n1659 VDD.n1658 10.6151
R20059 VDD.n1659 VDD.n545 10.6151
R20060 VDD.n1669 VDD.n545 10.6151
R20061 VDD.n1670 VDD.n1669 10.6151
R20062 VDD.n1671 VDD.n1670 10.6151
R20063 VDD.n1671 VDD.n533 10.6151
R20064 VDD.n1681 VDD.n533 10.6151
R20065 VDD.n1682 VDD.n1681 10.6151
R20066 VDD.n1683 VDD.n1682 10.6151
R20067 VDD.n1683 VDD.n520 10.6151
R20068 VDD.n1743 VDD.n520 10.6151
R20069 VDD.n1744 VDD.n1743 10.6151
R20070 VDD.n1745 VDD.n1744 10.6151
R20071 VDD.n1745 VDD.n510 10.6151
R20072 VDD.n1799 VDD.n510 10.6151
R20073 VDD.n1799 VDD.n1798 10.6151
R20074 VDD.n2320 VDD.n2319 10.6151
R20075 VDD.n2319 VDD.n2316 10.6151
R20076 VDD.n2316 VDD.n2315 10.6151
R20077 VDD.n2315 VDD.n2312 10.6151
R20078 VDD.n2312 VDD.n2311 10.6151
R20079 VDD.n2311 VDD.n2308 10.6151
R20080 VDD.n2308 VDD.n2307 10.6151
R20081 VDD.n2307 VDD.n2304 10.6151
R20082 VDD.n2304 VDD.n2303 10.6151
R20083 VDD.n2303 VDD.n2300 10.6151
R20084 VDD.n2300 VDD.n2299 10.6151
R20085 VDD.n2299 VDD.n2296 10.6151
R20086 VDD.n2296 VDD.n2295 10.6151
R20087 VDD.n2295 VDD.n2292 10.6151
R20088 VDD.n2292 VDD.n2291 10.6151
R20089 VDD.n2291 VDD.n2288 10.6151
R20090 VDD.n2288 VDD.n2287 10.6151
R20091 VDD.n2287 VDD.n2284 10.6151
R20092 VDD.n2284 VDD.n2283 10.6151
R20093 VDD.n2395 VDD.n282 10.6151
R20094 VDD.n1957 VDD.n1956 10.6151
R20095 VDD.n1956 VDD.n1955 10.6151
R20096 VDD.n1955 VDD.n1954 10.6151
R20097 VDD.n1954 VDD.n1952 10.6151
R20098 VDD.n1952 VDD.n1951 10.6151
R20099 VDD.n1951 VDD.n1949 10.6151
R20100 VDD.n1949 VDD.n1948 10.6151
R20101 VDD.n1948 VDD.n1946 10.6151
R20102 VDD.n1946 VDD.n1945 10.6151
R20103 VDD.n1945 VDD.n1943 10.6151
R20104 VDD.n1943 VDD.n1942 10.6151
R20105 VDD.n1942 VDD.n1940 10.6151
R20106 VDD.n1940 VDD.n1939 10.6151
R20107 VDD.n1939 VDD.n1937 10.6151
R20108 VDD.n1937 VDD.n1936 10.6151
R20109 VDD.n1936 VDD.n1934 10.6151
R20110 VDD.n1934 VDD.n1933 10.6151
R20111 VDD.n1933 VDD.n1931 10.6151
R20112 VDD.n1931 VDD.n1930 10.6151
R20113 VDD.n1930 VDD.n1928 10.6151
R20114 VDD.n1928 VDD.n1927 10.6151
R20115 VDD.n1927 VDD.n1925 10.6151
R20116 VDD.n1925 VDD.n1924 10.6151
R20117 VDD.n1924 VDD.n1922 10.6151
R20118 VDD.n1922 VDD.n1921 10.6151
R20119 VDD.n1921 VDD.n1919 10.6151
R20120 VDD.n1919 VDD.n1918 10.6151
R20121 VDD.n1918 VDD.n1916 10.6151
R20122 VDD.n1916 VDD.n1915 10.6151
R20123 VDD.n1915 VDD.n1913 10.6151
R20124 VDD.n1913 VDD.n1912 10.6151
R20125 VDD.n1912 VDD.n1910 10.6151
R20126 VDD.n1910 VDD.n1909 10.6151
R20127 VDD.n1909 VDD.n1907 10.6151
R20128 VDD.n1907 VDD.n1906 10.6151
R20129 VDD.n1906 VDD.n1904 10.6151
R20130 VDD.n1904 VDD.n1903 10.6151
R20131 VDD.n1903 VDD.n1901 10.6151
R20132 VDD.n1901 VDD.n1900 10.6151
R20133 VDD.n1900 VDD.n1898 10.6151
R20134 VDD.n1898 VDD.n1897 10.6151
R20135 VDD.n1897 VDD.n1895 10.6151
R20136 VDD.n1895 VDD.n1894 10.6151
R20137 VDD.n1894 VDD.n1892 10.6151
R20138 VDD.n1892 VDD.n1891 10.6151
R20139 VDD.n1891 VDD.n1889 10.6151
R20140 VDD.n1889 VDD.n1888 10.6151
R20141 VDD.n1888 VDD.n1886 10.6151
R20142 VDD.n1886 VDD.n1885 10.6151
R20143 VDD.n1885 VDD.n1883 10.6151
R20144 VDD.n1883 VDD.n1882 10.6151
R20145 VDD.n1882 VDD.n1880 10.6151
R20146 VDD.n1880 VDD.n1879 10.6151
R20147 VDD.n1879 VDD.n1877 10.6151
R20148 VDD.n1877 VDD.n1876 10.6151
R20149 VDD.n1876 VDD.n1874 10.6151
R20150 VDD.n1874 VDD.n1873 10.6151
R20151 VDD.n1873 VDD.n1871 10.6151
R20152 VDD.n1871 VDD.n1870 10.6151
R20153 VDD.n1870 VDD.n1868 10.6151
R20154 VDD.n1868 VDD.n283 10.6151
R20155 VDD.n2393 VDD.n283 10.6151
R20156 VDD.n2394 VDD.n2393 10.6151
R20157 VDD.n1827 VDD.n476 10.6151
R20158 VDD.n1828 VDD.n1827 10.6151
R20159 VDD.n1828 VDD.n1824 10.6151
R20160 VDD.n1834 VDD.n1824 10.6151
R20161 VDD.n1835 VDD.n1834 10.6151
R20162 VDD.n1836 VDD.n1835 10.6151
R20163 VDD.n1836 VDD.n1822 10.6151
R20164 VDD.n1842 VDD.n1822 10.6151
R20165 VDD.n1843 VDD.n1842 10.6151
R20166 VDD.n1844 VDD.n1843 10.6151
R20167 VDD.n1844 VDD.n1820 10.6151
R20168 VDD.n1850 VDD.n1820 10.6151
R20169 VDD.n1851 VDD.n1850 10.6151
R20170 VDD.n1852 VDD.n1851 10.6151
R20171 VDD.n1852 VDD.n1818 10.6151
R20172 VDD.n1858 VDD.n1818 10.6151
R20173 VDD.n1859 VDD.n1858 10.6151
R20174 VDD.n1860 VDD.n1859 10.6151
R20175 VDD.n1860 VDD.n1816 10.6151
R20176 VDD.n1867 VDD.n1866 10.6151
R20177 VDD.n2110 VDD.n2109 10.6151
R20178 VDD.n2111 VDD.n2110 10.6151
R20179 VDD.n2111 VDD.n464 10.6151
R20180 VDD.n2121 VDD.n464 10.6151
R20181 VDD.n2122 VDD.n2121 10.6151
R20182 VDD.n2123 VDD.n2122 10.6151
R20183 VDD.n2123 VDD.n452 10.6151
R20184 VDD.n2133 VDD.n452 10.6151
R20185 VDD.n2134 VDD.n2133 10.6151
R20186 VDD.n2135 VDD.n2134 10.6151
R20187 VDD.n2135 VDD.n440 10.6151
R20188 VDD.n2145 VDD.n440 10.6151
R20189 VDD.n2146 VDD.n2145 10.6151
R20190 VDD.n2147 VDD.n2146 10.6151
R20191 VDD.n2147 VDD.n428 10.6151
R20192 VDD.n2157 VDD.n428 10.6151
R20193 VDD.n2158 VDD.n2157 10.6151
R20194 VDD.n2159 VDD.n2158 10.6151
R20195 VDD.n2159 VDD.n416 10.6151
R20196 VDD.n2169 VDD.n416 10.6151
R20197 VDD.n2170 VDD.n2169 10.6151
R20198 VDD.n2171 VDD.n2170 10.6151
R20199 VDD.n2171 VDD.n404 10.6151
R20200 VDD.n2181 VDD.n404 10.6151
R20201 VDD.n2182 VDD.n2181 10.6151
R20202 VDD.n2183 VDD.n2182 10.6151
R20203 VDD.n2183 VDD.n392 10.6151
R20204 VDD.n2193 VDD.n392 10.6151
R20205 VDD.n2194 VDD.n2193 10.6151
R20206 VDD.n2195 VDD.n2194 10.6151
R20207 VDD.n2195 VDD.n380 10.6151
R20208 VDD.n2205 VDD.n380 10.6151
R20209 VDD.n2206 VDD.n2205 10.6151
R20210 VDD.n2207 VDD.n2206 10.6151
R20211 VDD.n2207 VDD.n367 10.6151
R20212 VDD.n2217 VDD.n367 10.6151
R20213 VDD.n2218 VDD.n2217 10.6151
R20214 VDD.n2219 VDD.n2218 10.6151
R20215 VDD.n2219 VDD.n356 10.6151
R20216 VDD.n2229 VDD.n356 10.6151
R20217 VDD.n2230 VDD.n2229 10.6151
R20218 VDD.n2231 VDD.n2230 10.6151
R20219 VDD.n2231 VDD.n344 10.6151
R20220 VDD.n2241 VDD.n344 10.6151
R20221 VDD.n2242 VDD.n2241 10.6151
R20222 VDD.n2243 VDD.n2242 10.6151
R20223 VDD.n2243 VDD.n332 10.6151
R20224 VDD.n2253 VDD.n332 10.6151
R20225 VDD.n2254 VDD.n2253 10.6151
R20226 VDD.n2255 VDD.n2254 10.6151
R20227 VDD.n2255 VDD.n319 10.6151
R20228 VDD.n2265 VDD.n319 10.6151
R20229 VDD.n2266 VDD.n2265 10.6151
R20230 VDD.n2267 VDD.n2266 10.6151
R20231 VDD.n2267 VDD.n308 10.6151
R20232 VDD.n2277 VDD.n308 10.6151
R20233 VDD.n2278 VDD.n2277 10.6151
R20234 VDD.n2329 VDD.n2278 10.6151
R20235 VDD.n2329 VDD.n2328 10.6151
R20236 VDD.n2328 VDD.n2327 10.6151
R20237 VDD.n2327 VDD.n2326 10.6151
R20238 VDD.n2326 VDD.n2324 10.6151
R20239 VDD.n2324 VDD.n2323 10.6151
R20240 VDD.n1730 VDD.n1729 10.6151
R20241 VDD.n1729 VDD.n1726 10.6151
R20242 VDD.n1726 VDD.n1725 10.6151
R20243 VDD.n1725 VDD.n1722 10.6151
R20244 VDD.n1722 VDD.n1721 10.6151
R20245 VDD.n1721 VDD.n1718 10.6151
R20246 VDD.n1718 VDD.n1717 10.6151
R20247 VDD.n1717 VDD.n1714 10.6151
R20248 VDD.n1714 VDD.n1713 10.6151
R20249 VDD.n1713 VDD.n1710 10.6151
R20250 VDD.n1710 VDD.n1709 10.6151
R20251 VDD.n1709 VDD.n1706 10.6151
R20252 VDD.n1706 VDD.n1705 10.6151
R20253 VDD.n1705 VDD.n1702 10.6151
R20254 VDD.n1702 VDD.n1701 10.6151
R20255 VDD.n1701 VDD.n1698 10.6151
R20256 VDD.n1698 VDD.n1697 10.6151
R20257 VDD.n1697 VDD.n1694 10.6151
R20258 VDD.n1694 VDD.n1693 10.6151
R20259 VDD.n1805 VDD.n502 10.6151
R20260 VDD.n1467 VDD.n1466 10.6151
R20261 VDD.n1466 VDD.n1464 10.6151
R20262 VDD.n1464 VDD.n1463 10.6151
R20263 VDD.n1463 VDD.n1461 10.6151
R20264 VDD.n1461 VDD.n1460 10.6151
R20265 VDD.n1460 VDD.n1458 10.6151
R20266 VDD.n1458 VDD.n1457 10.6151
R20267 VDD.n1457 VDD.n1455 10.6151
R20268 VDD.n1455 VDD.n1454 10.6151
R20269 VDD.n1454 VDD.n1452 10.6151
R20270 VDD.n1452 VDD.n1451 10.6151
R20271 VDD.n1451 VDD.n1449 10.6151
R20272 VDD.n1449 VDD.n1448 10.6151
R20273 VDD.n1448 VDD.n1446 10.6151
R20274 VDD.n1446 VDD.n1445 10.6151
R20275 VDD.n1445 VDD.n1443 10.6151
R20276 VDD.n1443 VDD.n1442 10.6151
R20277 VDD.n1442 VDD.n1440 10.6151
R20278 VDD.n1440 VDD.n1439 10.6151
R20279 VDD.n1439 VDD.n1437 10.6151
R20280 VDD.n1437 VDD.n1436 10.6151
R20281 VDD.n1436 VDD.n1434 10.6151
R20282 VDD.n1434 VDD.n1433 10.6151
R20283 VDD.n1433 VDD.n1431 10.6151
R20284 VDD.n1431 VDD.n1430 10.6151
R20285 VDD.n1430 VDD.n1428 10.6151
R20286 VDD.n1428 VDD.n1427 10.6151
R20287 VDD.n1427 VDD.n1425 10.6151
R20288 VDD.n1425 VDD.n1424 10.6151
R20289 VDD.n1424 VDD.n1422 10.6151
R20290 VDD.n1422 VDD.n1421 10.6151
R20291 VDD.n1421 VDD.n1419 10.6151
R20292 VDD.n1419 VDD.n1418 10.6151
R20293 VDD.n1418 VDD.n1416 10.6151
R20294 VDD.n1416 VDD.n1415 10.6151
R20295 VDD.n1415 VDD.n1413 10.6151
R20296 VDD.n1413 VDD.n1412 10.6151
R20297 VDD.n1412 VDD.n1410 10.6151
R20298 VDD.n1410 VDD.n1409 10.6151
R20299 VDD.n1409 VDD.n1407 10.6151
R20300 VDD.n1407 VDD.n1406 10.6151
R20301 VDD.n1406 VDD.n1404 10.6151
R20302 VDD.n1404 VDD.n1403 10.6151
R20303 VDD.n1403 VDD.n1401 10.6151
R20304 VDD.n1401 VDD.n1400 10.6151
R20305 VDD.n1400 VDD.n1398 10.6151
R20306 VDD.n1398 VDD.n1397 10.6151
R20307 VDD.n1397 VDD.n1395 10.6151
R20308 VDD.n1395 VDD.n1394 10.6151
R20309 VDD.n1394 VDD.n1392 10.6151
R20310 VDD.n1392 VDD.n1391 10.6151
R20311 VDD.n1391 VDD.n1389 10.6151
R20312 VDD.n1389 VDD.n1388 10.6151
R20313 VDD.n1388 VDD.n1386 10.6151
R20314 VDD.n1386 VDD.n1385 10.6151
R20315 VDD.n1385 VDD.n1383 10.6151
R20316 VDD.n1383 VDD.n1382 10.6151
R20317 VDD.n1382 VDD.n1380 10.6151
R20318 VDD.n1380 VDD.n1379 10.6151
R20319 VDD.n1379 VDD.n1377 10.6151
R20320 VDD.n1377 VDD.n503 10.6151
R20321 VDD.n1803 VDD.n503 10.6151
R20322 VDD.n1804 VDD.n1803 10.6151
R20323 VDD.n1507 VDD.n695 10.6151
R20324 VDD.n1507 VDD.n1506 10.6151
R20325 VDD.n1506 VDD.n1505 10.6151
R20326 VDD.n1505 VDD.n1502 10.6151
R20327 VDD.n1502 VDD.n1501 10.6151
R20328 VDD.n1501 VDD.n1498 10.6151
R20329 VDD.n1498 VDD.n1497 10.6151
R20330 VDD.n1497 VDD.n1494 10.6151
R20331 VDD.n1494 VDD.n1493 10.6151
R20332 VDD.n1493 VDD.n1490 10.6151
R20333 VDD.n1490 VDD.n1489 10.6151
R20334 VDD.n1489 VDD.n1486 10.6151
R20335 VDD.n1486 VDD.n1485 10.6151
R20336 VDD.n1485 VDD.n1482 10.6151
R20337 VDD.n1482 VDD.n1481 10.6151
R20338 VDD.n1481 VDD.n1478 10.6151
R20339 VDD.n1478 VDD.n1477 10.6151
R20340 VDD.n1477 VDD.n1474 10.6151
R20341 VDD.n1474 VDD.n1473 10.6151
R20342 VDD.n1470 VDD.n1469 10.6151
R20343 VDD.n1520 VDD.n1519 10.6151
R20344 VDD.n1521 VDD.n1520 10.6151
R20345 VDD.n1521 VDD.n683 10.6151
R20346 VDD.n1531 VDD.n683 10.6151
R20347 VDD.n1532 VDD.n1531 10.6151
R20348 VDD.n1533 VDD.n1532 10.6151
R20349 VDD.n1533 VDD.n670 10.6151
R20350 VDD.n1543 VDD.n670 10.6151
R20351 VDD.n1544 VDD.n1543 10.6151
R20352 VDD.n1545 VDD.n1544 10.6151
R20353 VDD.n1545 VDD.n659 10.6151
R20354 VDD.n1555 VDD.n659 10.6151
R20355 VDD.n1556 VDD.n1555 10.6151
R20356 VDD.n1557 VDD.n1556 10.6151
R20357 VDD.n1557 VDD.n647 10.6151
R20358 VDD.n1567 VDD.n647 10.6151
R20359 VDD.n1568 VDD.n1567 10.6151
R20360 VDD.n1569 VDD.n1568 10.6151
R20361 VDD.n1569 VDD.n635 10.6151
R20362 VDD.n1579 VDD.n635 10.6151
R20363 VDD.n1580 VDD.n1579 10.6151
R20364 VDD.n1581 VDD.n1580 10.6151
R20365 VDD.n1581 VDD.n622 10.6151
R20366 VDD.n1591 VDD.n622 10.6151
R20367 VDD.n1592 VDD.n1591 10.6151
R20368 VDD.n1593 VDD.n1592 10.6151
R20369 VDD.n1593 VDD.n611 10.6151
R20370 VDD.n1603 VDD.n611 10.6151
R20371 VDD.n1604 VDD.n1603 10.6151
R20372 VDD.n1605 VDD.n1604 10.6151
R20373 VDD.n1605 VDD.n599 10.6151
R20374 VDD.n1615 VDD.n599 10.6151
R20375 VDD.n1616 VDD.n1615 10.6151
R20376 VDD.n1617 VDD.n1616 10.6151
R20377 VDD.n1617 VDD.n587 10.6151
R20378 VDD.n1627 VDD.n587 10.6151
R20379 VDD.n1628 VDD.n1627 10.6151
R20380 VDD.n1629 VDD.n1628 10.6151
R20381 VDD.n1629 VDD.n575 10.6151
R20382 VDD.n1639 VDD.n575 10.6151
R20383 VDD.n1640 VDD.n1639 10.6151
R20384 VDD.n1641 VDD.n1640 10.6151
R20385 VDD.n1641 VDD.n563 10.6151
R20386 VDD.n1651 VDD.n563 10.6151
R20387 VDD.n1652 VDD.n1651 10.6151
R20388 VDD.n1653 VDD.n1652 10.6151
R20389 VDD.n1653 VDD.n551 10.6151
R20390 VDD.n1663 VDD.n551 10.6151
R20391 VDD.n1664 VDD.n1663 10.6151
R20392 VDD.n1665 VDD.n1664 10.6151
R20393 VDD.n1665 VDD.n539 10.6151
R20394 VDD.n1675 VDD.n539 10.6151
R20395 VDD.n1676 VDD.n1675 10.6151
R20396 VDD.n1677 VDD.n1676 10.6151
R20397 VDD.n1677 VDD.n527 10.6151
R20398 VDD.n1687 VDD.n527 10.6151
R20399 VDD.n1688 VDD.n1687 10.6151
R20400 VDD.n1739 VDD.n1688 10.6151
R20401 VDD.n1739 VDD.n1738 10.6151
R20402 VDD.n1738 VDD.n1737 10.6151
R20403 VDD.n1737 VDD.n1736 10.6151
R20404 VDD.n1736 VDD.n1734 10.6151
R20405 VDD.n1734 VDD.n1733 10.6151
R20406 VDD.n932 VDD.n931 10.0853
R20407 VDD.n2456 VDD.n2453 10.0853
R20408 VDD.n138 VDD.n113 10.0853
R20409 VDD.n1196 VDD.n1195 10.0853
R20410 VDD.n1547 VDD.t19 9.35759
R20411 VDD.n324 VDD.t17 9.35759
R20412 VDD.n120 VDD.n117 9.3005
R20413 VDD.n124 VDD.n121 9.3005
R20414 VDD.n125 VDD.n116 9.3005
R20415 VDD.n129 VDD.n128 9.3005
R20416 VDD.n130 VDD.n115 9.3005
R20417 VDD.n134 VDD.n131 9.3005
R20418 VDD.n135 VDD.n114 9.3005
R20419 VDD.n139 VDD.n138 9.3005
R20420 VDD.n140 VDD.n113 9.3005
R20421 VDD.n144 VDD.n141 9.3005
R20422 VDD.n145 VDD.n110 9.3005
R20423 VDD.n149 VDD.n148 9.3005
R20424 VDD.n150 VDD.n109 9.3005
R20425 VDD.n154 VDD.n151 9.3005
R20426 VDD.n155 VDD.n108 9.3005
R20427 VDD.n159 VDD.n158 9.3005
R20428 VDD.n160 VDD.n107 9.3005
R20429 VDD.n164 VDD.n161 9.3005
R20430 VDD.n166 VDD.n106 9.3005
R20431 VDD.n168 VDD.n167 9.3005
R20432 VDD.n2620 VDD.n2619 9.3005
R20433 VDD.n119 VDD.n118 9.3005
R20434 VDD.n2478 VDD.n2477 9.3005
R20435 VDD.n242 VDD.n241 9.3005
R20436 VDD.n2491 VDD.n2490 9.3005
R20437 VDD.n2492 VDD.n240 9.3005
R20438 VDD.n2494 VDD.n2493 9.3005
R20439 VDD.n231 VDD.n230 9.3005
R20440 VDD.n2507 VDD.n2506 9.3005
R20441 VDD.n2508 VDD.n229 9.3005
R20442 VDD.n2510 VDD.n2509 9.3005
R20443 VDD.n219 VDD.n218 9.3005
R20444 VDD.n2523 VDD.n2522 9.3005
R20445 VDD.n2524 VDD.n217 9.3005
R20446 VDD.n2526 VDD.n2525 9.3005
R20447 VDD.n207 VDD.n206 9.3005
R20448 VDD.n2539 VDD.n2538 9.3005
R20449 VDD.n2540 VDD.n205 9.3005
R20450 VDD.n2542 VDD.n2541 9.3005
R20451 VDD.n195 VDD.n194 9.3005
R20452 VDD.n2555 VDD.n2554 9.3005
R20453 VDD.n2556 VDD.n193 9.3005
R20454 VDD.n2561 VDD.n2557 9.3005
R20455 VDD.n2560 VDD.n2559 9.3005
R20456 VDD.n2558 VDD.n182 9.3005
R20457 VDD.n2574 VDD.n181 9.3005
R20458 VDD.n2576 VDD.n2575 9.3005
R20459 VDD.n2577 VDD.n180 9.3005
R20460 VDD.n2579 VDD.n2578 9.3005
R20461 VDD.n2581 VDD.n179 9.3005
R20462 VDD.n2583 VDD.n2582 9.3005
R20463 VDD.n2584 VDD.n178 9.3005
R20464 VDD.n2586 VDD.n2585 9.3005
R20465 VDD.n2588 VDD.n177 9.3005
R20466 VDD.n2590 VDD.n2589 9.3005
R20467 VDD.n2591 VDD.n176 9.3005
R20468 VDD.n2593 VDD.n2592 9.3005
R20469 VDD.n2595 VDD.n175 9.3005
R20470 VDD.n2597 VDD.n2596 9.3005
R20471 VDD.n2598 VDD.n174 9.3005
R20472 VDD.n2600 VDD.n2599 9.3005
R20473 VDD.n2602 VDD.n173 9.3005
R20474 VDD.n2604 VDD.n2603 9.3005
R20475 VDD.n2605 VDD.n172 9.3005
R20476 VDD.n2607 VDD.n2606 9.3005
R20477 VDD.n2609 VDD.n171 9.3005
R20478 VDD.n2611 VDD.n2610 9.3005
R20479 VDD.n2612 VDD.n170 9.3005
R20480 VDD.n2614 VDD.n2613 9.3005
R20481 VDD.n2616 VDD.n169 9.3005
R20482 VDD.n2618 VDD.n2617 9.3005
R20483 VDD.n2476 VDD.n253 9.3005
R20484 VDD.n2432 VDD.n254 9.3005
R20485 VDD.n2433 VDD.n2431 9.3005
R20486 VDD.n2436 VDD.n2430 9.3005
R20487 VDD.n2437 VDD.n2429 9.3005
R20488 VDD.n2440 VDD.n2428 9.3005
R20489 VDD.n2441 VDD.n2427 9.3005
R20490 VDD.n2444 VDD.n2426 9.3005
R20491 VDD.n2445 VDD.n2425 9.3005
R20492 VDD.n2448 VDD.n2424 9.3005
R20493 VDD.n2449 VDD.n2423 9.3005
R20494 VDD.n2452 VDD.n2422 9.3005
R20495 VDD.n2453 VDD.n2419 9.3005
R20496 VDD.n2456 VDD.n2418 9.3005
R20497 VDD.n2457 VDD.n2417 9.3005
R20498 VDD.n2460 VDD.n2416 9.3005
R20499 VDD.n2461 VDD.n2415 9.3005
R20500 VDD.n2464 VDD.n2414 9.3005
R20501 VDD.n2466 VDD.n2413 9.3005
R20502 VDD.n2467 VDD.n2412 9.3005
R20503 VDD.n2468 VDD.n2411 9.3005
R20504 VDD.n2469 VDD.n2410 9.3005
R20505 VDD.n2475 VDD.n2474 9.3005
R20506 VDD.n2483 VDD.n2482 9.3005
R20507 VDD.n2484 VDD.n247 9.3005
R20508 VDD.n2486 VDD.n2485 9.3005
R20509 VDD.n237 VDD.n236 9.3005
R20510 VDD.n2499 VDD.n2498 9.3005
R20511 VDD.n2500 VDD.n235 9.3005
R20512 VDD.n2502 VDD.n2501 9.3005
R20513 VDD.n225 VDD.n224 9.3005
R20514 VDD.n2515 VDD.n2514 9.3005
R20515 VDD.n2516 VDD.n223 9.3005
R20516 VDD.n2518 VDD.n2517 9.3005
R20517 VDD.n213 VDD.n212 9.3005
R20518 VDD.n2531 VDD.n2530 9.3005
R20519 VDD.n2532 VDD.n211 9.3005
R20520 VDD.n2534 VDD.n2533 9.3005
R20521 VDD.n201 VDD.n200 9.3005
R20522 VDD.n2547 VDD.n2546 9.3005
R20523 VDD.n2548 VDD.n199 9.3005
R20524 VDD.n2550 VDD.n2549 9.3005
R20525 VDD.n188 VDD.n187 9.3005
R20526 VDD.n2566 VDD.n2565 9.3005
R20527 VDD.n2567 VDD.n186 9.3005
R20528 VDD.n2569 VDD.n2568 9.3005
R20529 VDD.n23 VDD.n21 9.3005
R20530 VDD.n2675 VDD.n2674 9.3005
R20531 VDD.n24 VDD.n22 9.3005
R20532 VDD.n2668 VDD.n32 9.3005
R20533 VDD.n2667 VDD.n33 9.3005
R20534 VDD.n2666 VDD.n34 9.3005
R20535 VDD.n42 VDD.n35 9.3005
R20536 VDD.n2660 VDD.n43 9.3005
R20537 VDD.n2659 VDD.n44 9.3005
R20538 VDD.n2658 VDD.n45 9.3005
R20539 VDD.n53 VDD.n46 9.3005
R20540 VDD.n2652 VDD.n54 9.3005
R20541 VDD.n2651 VDD.n55 9.3005
R20542 VDD.n2650 VDD.n56 9.3005
R20543 VDD.n64 VDD.n57 9.3005
R20544 VDD.n2644 VDD.n65 9.3005
R20545 VDD.n2643 VDD.n66 9.3005
R20546 VDD.n2642 VDD.n67 9.3005
R20547 VDD.n75 VDD.n68 9.3005
R20548 VDD.n2636 VDD.n76 9.3005
R20549 VDD.n2635 VDD.n77 9.3005
R20550 VDD.n2634 VDD.n78 9.3005
R20551 VDD.n86 VDD.n79 9.3005
R20552 VDD.n2628 VDD.n87 9.3005
R20553 VDD.n2627 VDD.n88 9.3005
R20554 VDD.n2626 VDD.n89 9.3005
R20555 VDD.n249 VDD.n248 9.3005
R20556 VDD.n788 VDD.n787 9.3005
R20557 VDD.n1064 VDD.n1063 9.3005
R20558 VDD.n1065 VDD.n786 9.3005
R20559 VDD.n1067 VDD.n1066 9.3005
R20560 VDD.n776 VDD.n775 9.3005
R20561 VDD.n1080 VDD.n1079 9.3005
R20562 VDD.n1081 VDD.n774 9.3005
R20563 VDD.n1083 VDD.n1082 9.3005
R20564 VDD.n764 VDD.n763 9.3005
R20565 VDD.n1096 VDD.n1095 9.3005
R20566 VDD.n1097 VDD.n762 9.3005
R20567 VDD.n1099 VDD.n1098 9.3005
R20568 VDD.n752 VDD.n751 9.3005
R20569 VDD.n1112 VDD.n1111 9.3005
R20570 VDD.n1113 VDD.n750 9.3005
R20571 VDD.n1115 VDD.n1114 9.3005
R20572 VDD.n740 VDD.n739 9.3005
R20573 VDD.n1128 VDD.n1127 9.3005
R20574 VDD.n1129 VDD.n738 9.3005
R20575 VDD.n1131 VDD.n1130 9.3005
R20576 VDD.n728 VDD.n727 9.3005
R20577 VDD.n1145 VDD.n1144 9.3005
R20578 VDD.n1146 VDD.n725 9.3005
R20579 VDD.n1212 VDD.n1211 9.3005
R20580 VDD.n1210 VDD.n726 9.3005
R20581 VDD.n1207 VDD.n1147 9.3005
R20582 VDD.n1206 VDD.n1205 9.3005
R20583 VDD.n1204 VDD.n1151 9.3005
R20584 VDD.n1203 VDD.n1202 9.3005
R20585 VDD.n1201 VDD.n1152 9.3005
R20586 VDD.n1200 VDD.n1199 9.3005
R20587 VDD.n1198 VDD.n1157 9.3005
R20588 VDD.n1197 VDD.n1196 9.3005
R20589 VDD.n1195 VDD.n1158 9.3005
R20590 VDD.n1194 VDD.n1193 9.3005
R20591 VDD.n1192 VDD.n1165 9.3005
R20592 VDD.n1191 VDD.n1190 9.3005
R20593 VDD.n1189 VDD.n1166 9.3005
R20594 VDD.n1188 VDD.n1187 9.3005
R20595 VDD.n1186 VDD.n1171 9.3005
R20596 VDD.n1185 VDD.n1184 9.3005
R20597 VDD.n1183 VDD.n1172 9.3005
R20598 VDD.n1182 VDD.n1181 9.3005
R20599 VDD.n1180 VDD.n1179 9.3005
R20600 VDD.n1178 VDD.n718 9.3005
R20601 VDD.n1220 VDD.n1219 9.3005
R20602 VDD.n1209 VDD.n1208 9.3005
R20603 VDD.n953 VDD.n863 9.3005
R20604 VDD.n955 VDD.n954 9.3005
R20605 VDD.n853 VDD.n852 9.3005
R20606 VDD.n968 VDD.n967 9.3005
R20607 VDD.n969 VDD.n851 9.3005
R20608 VDD.n971 VDD.n970 9.3005
R20609 VDD.n841 VDD.n840 9.3005
R20610 VDD.n984 VDD.n983 9.3005
R20611 VDD.n985 VDD.n839 9.3005
R20612 VDD.n987 VDD.n986 9.3005
R20613 VDD.n829 VDD.n828 9.3005
R20614 VDD.n1000 VDD.n999 9.3005
R20615 VDD.n1001 VDD.n827 9.3005
R20616 VDD.n1003 VDD.n1002 9.3005
R20617 VDD.n818 VDD.n817 9.3005
R20618 VDD.n1017 VDD.n1016 9.3005
R20619 VDD.n1018 VDD.n816 9.3005
R20620 VDD.n1020 VDD.n1019 9.3005
R20621 VDD.n806 VDD.n805 9.3005
R20622 VDD.n1033 VDD.n1032 9.3005
R20623 VDD.n1034 VDD.n804 9.3005
R20624 VDD.n1036 VDD.n1035 9.3005
R20625 VDD.n794 VDD.n793 9.3005
R20626 VDD.n1056 VDD.n1055 9.3005
R20627 VDD.n1057 VDD.n792 9.3005
R20628 VDD.n1059 VDD.n1058 9.3005
R20629 VDD.n782 VDD.n781 9.3005
R20630 VDD.n1072 VDD.n1071 9.3005
R20631 VDD.n1073 VDD.n780 9.3005
R20632 VDD.n1075 VDD.n1074 9.3005
R20633 VDD.n769 VDD.n768 9.3005
R20634 VDD.n1088 VDD.n1087 9.3005
R20635 VDD.n1089 VDD.n767 9.3005
R20636 VDD.n1091 VDD.n1090 9.3005
R20637 VDD.n758 VDD.n757 9.3005
R20638 VDD.n1104 VDD.n1103 9.3005
R20639 VDD.n1105 VDD.n756 9.3005
R20640 VDD.n1107 VDD.n1106 9.3005
R20641 VDD.n746 VDD.n745 9.3005
R20642 VDD.n1120 VDD.n1119 9.3005
R20643 VDD.n1121 VDD.n744 9.3005
R20644 VDD.n1123 VDD.n1122 9.3005
R20645 VDD.n734 VDD.n733 9.3005
R20646 VDD.n1136 VDD.n1135 9.3005
R20647 VDD.n1137 VDD.n732 9.3005
R20648 VDD.n1140 VDD.n1139 9.3005
R20649 VDD.n1138 VDD.n720 9.3005
R20650 VDD.n1216 VDD.n719 9.3005
R20651 VDD.n1218 VDD.n1217 9.3005
R20652 VDD.n952 VDD.n951 9.3005
R20653 VDD.n910 VDD.n909 9.3005
R20654 VDD.n912 VDD.n911 9.3005
R20655 VDD.n913 VDD.n896 9.3005
R20656 VDD.n915 VDD.n914 9.3005
R20657 VDD.n916 VDD.n895 9.3005
R20658 VDD.n918 VDD.n917 9.3005
R20659 VDD.n919 VDD.n889 9.3005
R20660 VDD.n921 VDD.n920 9.3005
R20661 VDD.n922 VDD.n887 9.3005
R20662 VDD.n924 VDD.n923 9.3005
R20663 VDD.n888 VDD.n885 9.3005
R20664 VDD.n931 VDD.n881 9.3005
R20665 VDD.n933 VDD.n932 9.3005
R20666 VDD.n934 VDD.n880 9.3005
R20667 VDD.n936 VDD.n935 9.3005
R20668 VDD.n937 VDD.n873 9.3005
R20669 VDD.n939 VDD.n938 9.3005
R20670 VDD.n940 VDD.n872 9.3005
R20671 VDD.n942 VDD.n941 9.3005
R20672 VDD.n943 VDD.n868 9.3005
R20673 VDD.n945 VDD.n944 9.3005
R20674 VDD.n905 VDD.n864 9.3005
R20675 VDD.n859 VDD.n858 9.3005
R20676 VDD.n960 VDD.n959 9.3005
R20677 VDD.n961 VDD.n857 9.3005
R20678 VDD.n963 VDD.n962 9.3005
R20679 VDD.n847 VDD.n846 9.3005
R20680 VDD.n976 VDD.n975 9.3005
R20681 VDD.n977 VDD.n845 9.3005
R20682 VDD.n979 VDD.n978 9.3005
R20683 VDD.n835 VDD.n834 9.3005
R20684 VDD.n992 VDD.n991 9.3005
R20685 VDD.n993 VDD.n833 9.3005
R20686 VDD.n995 VDD.n994 9.3005
R20687 VDD.n823 VDD.n822 9.3005
R20688 VDD.n1009 VDD.n1008 9.3005
R20689 VDD.n1010 VDD.n821 9.3005
R20690 VDD.n1012 VDD.n1011 9.3005
R20691 VDD.n812 VDD.n811 9.3005
R20692 VDD.n1025 VDD.n1024 9.3005
R20693 VDD.n1026 VDD.n810 9.3005
R20694 VDD.n1028 VDD.n1027 9.3005
R20695 VDD.n800 VDD.n799 9.3005
R20696 VDD.n1041 VDD.n1040 9.3005
R20697 VDD.n1042 VDD.n798 9.3005
R20698 VDD.n1051 VDD.n1050 9.3005
R20699 VDD.n947 VDD.n946 9.3005
R20700 VDD.n18 VDD.t89 9.23488
R20701 VDD.n18 VDD.t103 9.23488
R20702 VDD.n16 VDD.t88 9.23488
R20703 VDD.n16 VDD.t95 9.23488
R20704 VDD.n1045 VDD.t100 9.23488
R20705 VDD.n1045 VDD.t101 9.23488
R20706 VDD.n1043 VDD.t91 9.23488
R20707 VDD.n1043 VDD.t93 9.23488
R20708 VDD.n1047 VDD.n1044 9.2074
R20709 VDD.n1053 VDD.t92 8.50695
R20710 VDD.t92 VDD.n790 8.50695
R20711 VDD.n2572 VDD.t94 8.50695
R20712 VDD.n2672 VDD.t94 8.50695
R20713 VDD.n15 VDD.n14 8.26582
R20714 VDD.n2677 VDD.n2676 8.24962
R20715 VDD.n1049 VDD.n1048 8.24962
R20716 VDD.n627 VDD.t112 7.99656
R20717 VDD.n2221 VDD.t82 7.99656
R20718 VDD.n2677 VDD.n20 7.97925
R20719 VDD.n1048 VDD.n1047 7.97925
R20720 VDD.n20 VDD.n17 7.31515
R20721 VDD.n1625 VDD.t23 6.97579
R20722 VDD.t15 VDD.n394 6.97579
R20723 VDD.n1577 VDD.t1 6.80566
R20724 VDD.t14 VDD.n565 6.80566
R20725 VDD.n2167 VDD.t5 6.80566
R20726 VDD.t0 VDD.n346 6.80566
R20727 VDD.n1047 VDD.n1046 6.77636
R20728 VDD.t6 VDD.n516 6.63553
R20729 VDD.n2119 VDD.t107 6.63553
R20730 VDD.t35 VDD.n672 6.12514
R20731 VDD.n1685 VDD.t45 6.12514
R20732 VDD.t49 VDD.n454 6.12514
R20733 VDD.n2275 VDD.t53 6.12514
R20734 VDD.n7 VDD.t9 6.12197
R20735 VDD.n7 VDD.t22 6.12197
R20736 VDD.n8 VDD.t18 6.12197
R20737 VDD.n8 VDD.t13 6.12197
R20738 VDD.n10 VDD.t16 6.12197
R20739 VDD.n10 VDD.t83 6.12197
R20740 VDD.n12 VDD.t108 6.12197
R20741 VDD.n12 VDD.t111 6.12197
R20742 VDD.n5 VDD.t3 6.12197
R20743 VDD.n5 VDD.t7 6.12197
R20744 VDD.n3 VDD.t113 6.12197
R20745 VDD.n3 VDD.t24 6.12197
R20746 VDD.n1 VDD.t106 6.12197
R20747 VDD.n1 VDD.t20 6.12197
R20748 VDD.n0 VDD.t11 6.12197
R20749 VDD.n0 VDD.t86 6.12197
R20750 VDD.n561 VDD.t2 5.95501
R20751 VDD.n2155 VDD.t110 5.95501
R20752 VDD.n609 VDD.t25 5.78488
R20753 VDD.n1613 VDD.t25 5.78488
R20754 VDD.n390 VDD.t4 5.78488
R20755 VDD.n2203 VDD.t4 5.78488
R20756 VDD.n2349 VDD.n294 5.62001
R20757 VDD.n2067 VDD.n2066 5.62001
R20758 VDD.n1759 VDD.n513 5.62001
R20759 VDD.n1270 VDD.n1269 5.62001
R20760 VDD.n2283 VDD.n2281 5.62001
R20761 VDD.n1816 VDD.n1815 5.62001
R20762 VDD.n1693 VDD.n1691 5.62001
R20763 VDD.n1473 VDD.n1376 5.62001
R20764 VDD.n1661 VDD.t2 5.61475
R20765 VDD.n438 VDD.t110 5.61475
R20766 VDD.n1535 VDD.t35 5.44463
R20767 VDD.t45 VDD.n522 5.44463
R20768 VDD.n2125 VDD.t49 5.44463
R20769 VDD.t53 VDD.n303 5.44463
R20770 VDD.n908 VDD.n905 5.04292
R20771 VDD.n2474 VDD.n257 5.04292
R20772 VDD.n2620 VDD.n105 5.04292
R20773 VDD.n1220 VDD.n717 5.04292
R20774 VDD.n2346 VDD.n294 4.99562
R20775 VDD.n2066 VDD.n2065 4.99562
R20776 VDD.n1756 VDD.n513 4.99562
R20777 VDD.n1271 VDD.n1270 4.99562
R20778 VDD.n2281 VDD.n282 4.99562
R20779 VDD.n1866 VDD.n1815 4.99562
R20780 VDD.n1691 VDD.n502 4.99562
R20781 VDD.n1470 VDD.n1376 4.99562
R20782 VDD.n1741 VDD.t6 4.93424
R20783 VDD.t107 VDD.n460 4.93424
R20784 VDD.n20 VDD.n19 4.88412
R20785 VDD.n1014 VDD.t90 4.76411
R20786 VDD.n772 VDD.t98 4.76411
R20787 VDD.t1 VDD.n631 4.76411
R20788 VDD.n1643 VDD.t14 4.76411
R20789 VDD.t5 VDD.n412 4.76411
R20790 VDD.n2233 VDD.t0 4.76411
R20791 VDD.t87 VDD.n203 4.76411
R20792 VDD.n2656 VDD.t96 4.76411
R20793 VDD.t23 VDD.n583 4.59398
R20794 VDD.n2185 VDD.t15 4.59398
R20795 VDD.t27 VDD.n849 4.08359
R20796 VDD.n1133 VDD.t60 4.08359
R20797 VDD.n2496 VDD.t67 4.08359
R20798 VDD.t31 VDD.n73 4.08359
R20799 VDD.n11 VDD.n9 4.01774
R20800 VDD.n4 VDD.n2 4.01774
R20801 VDD.n1595 VDD.t112 3.57321
R20802 VDD.n372 VDD.t82 3.57321
R20803 VDD.n13 VDD.n11 3.19878
R20804 VDD.n6 VDD.n4 3.19878
R20805 VDD.n14 VDD.n13 2.48474
R20806 VDD.n14 VDD.n6 2.48474
R20807 VDD.n675 VDD.t19 2.21218
R20808 VDD.n2269 VDD.t17 2.21218
R20809 VDD.n1510 VDD.t105 2.04205
R20810 VDD.n2398 VDD.t12 2.04205
R20811 VDD.n1048 VDD.n15 1.70911
R20812 VDD VDD.n2677 1.70127
R20813 VDD.n909 VDD.n908 1.55202
R20814 VDD.n2432 VDD.n257 1.55202
R20815 VDD.n167 VDD.n105 1.55202
R20816 VDD.n1178 VDD.n717 1.55202
R20817 VDD.n119 VDD.n89 0.473061
R20818 VDD.n2619 VDD.n2618 0.473061
R20819 VDD.n2476 VDD.n2475 0.473061
R20820 VDD.n2410 VDD.n248 0.473061
R20821 VDD.n1210 VDD.n1209 0.473061
R20822 VDD.n1219 VDD.n1218 0.473061
R20823 VDD.n952 VDD.n864 0.473061
R20824 VDD.n946 VDD.n945 0.473061
R20825 VDD.n2675 VDD.n22 0.152939
R20826 VDD.n32 VDD.n22 0.152939
R20827 VDD.n33 VDD.n32 0.152939
R20828 VDD.n34 VDD.n33 0.152939
R20829 VDD.n42 VDD.n34 0.152939
R20830 VDD.n43 VDD.n42 0.152939
R20831 VDD.n44 VDD.n43 0.152939
R20832 VDD.n45 VDD.n44 0.152939
R20833 VDD.n53 VDD.n45 0.152939
R20834 VDD.n54 VDD.n53 0.152939
R20835 VDD.n55 VDD.n54 0.152939
R20836 VDD.n56 VDD.n55 0.152939
R20837 VDD.n64 VDD.n56 0.152939
R20838 VDD.n65 VDD.n64 0.152939
R20839 VDD.n66 VDD.n65 0.152939
R20840 VDD.n67 VDD.n66 0.152939
R20841 VDD.n75 VDD.n67 0.152939
R20842 VDD.n76 VDD.n75 0.152939
R20843 VDD.n77 VDD.n76 0.152939
R20844 VDD.n78 VDD.n77 0.152939
R20845 VDD.n86 VDD.n78 0.152939
R20846 VDD.n87 VDD.n86 0.152939
R20847 VDD.n88 VDD.n87 0.152939
R20848 VDD.n89 VDD.n88 0.152939
R20849 VDD.n120 VDD.n119 0.152939
R20850 VDD.n121 VDD.n120 0.152939
R20851 VDD.n121 VDD.n116 0.152939
R20852 VDD.n129 VDD.n116 0.152939
R20853 VDD.n130 VDD.n129 0.152939
R20854 VDD.n131 VDD.n130 0.152939
R20855 VDD.n131 VDD.n114 0.152939
R20856 VDD.n139 VDD.n114 0.152939
R20857 VDD.n140 VDD.n139 0.152939
R20858 VDD.n141 VDD.n140 0.152939
R20859 VDD.n141 VDD.n110 0.152939
R20860 VDD.n149 VDD.n110 0.152939
R20861 VDD.n150 VDD.n149 0.152939
R20862 VDD.n151 VDD.n150 0.152939
R20863 VDD.n151 VDD.n108 0.152939
R20864 VDD.n159 VDD.n108 0.152939
R20865 VDD.n160 VDD.n159 0.152939
R20866 VDD.n161 VDD.n160 0.152939
R20867 VDD.n161 VDD.n106 0.152939
R20868 VDD.n168 VDD.n106 0.152939
R20869 VDD.n2619 VDD.n168 0.152939
R20870 VDD.n2477 VDD.n2476 0.152939
R20871 VDD.n2477 VDD.n241 0.152939
R20872 VDD.n2491 VDD.n241 0.152939
R20873 VDD.n2492 VDD.n2491 0.152939
R20874 VDD.n2493 VDD.n2492 0.152939
R20875 VDD.n2493 VDD.n230 0.152939
R20876 VDD.n2507 VDD.n230 0.152939
R20877 VDD.n2508 VDD.n2507 0.152939
R20878 VDD.n2509 VDD.n2508 0.152939
R20879 VDD.n2509 VDD.n218 0.152939
R20880 VDD.n2523 VDD.n218 0.152939
R20881 VDD.n2524 VDD.n2523 0.152939
R20882 VDD.n2525 VDD.n2524 0.152939
R20883 VDD.n2525 VDD.n206 0.152939
R20884 VDD.n2539 VDD.n206 0.152939
R20885 VDD.n2540 VDD.n2539 0.152939
R20886 VDD.n2541 VDD.n2540 0.152939
R20887 VDD.n2541 VDD.n194 0.152939
R20888 VDD.n2555 VDD.n194 0.152939
R20889 VDD.n2556 VDD.n2555 0.152939
R20890 VDD.n2557 VDD.n2556 0.152939
R20891 VDD.n2559 VDD.n2557 0.152939
R20892 VDD.n2559 VDD.n2558 0.152939
R20893 VDD.n2558 VDD.n181 0.152939
R20894 VDD.n2576 VDD.n181 0.152939
R20895 VDD.n2577 VDD.n2576 0.152939
R20896 VDD.n2578 VDD.n2577 0.152939
R20897 VDD.n2578 VDD.n179 0.152939
R20898 VDD.n2583 VDD.n179 0.152939
R20899 VDD.n2584 VDD.n2583 0.152939
R20900 VDD.n2585 VDD.n2584 0.152939
R20901 VDD.n2585 VDD.n177 0.152939
R20902 VDD.n2590 VDD.n177 0.152939
R20903 VDD.n2591 VDD.n2590 0.152939
R20904 VDD.n2592 VDD.n2591 0.152939
R20905 VDD.n2592 VDD.n175 0.152939
R20906 VDD.n2597 VDD.n175 0.152939
R20907 VDD.n2598 VDD.n2597 0.152939
R20908 VDD.n2599 VDD.n2598 0.152939
R20909 VDD.n2599 VDD.n173 0.152939
R20910 VDD.n2604 VDD.n173 0.152939
R20911 VDD.n2605 VDD.n2604 0.152939
R20912 VDD.n2606 VDD.n2605 0.152939
R20913 VDD.n2606 VDD.n171 0.152939
R20914 VDD.n2611 VDD.n171 0.152939
R20915 VDD.n2612 VDD.n2611 0.152939
R20916 VDD.n2613 VDD.n2612 0.152939
R20917 VDD.n2613 VDD.n169 0.152939
R20918 VDD.n2618 VDD.n169 0.152939
R20919 VDD.n2411 VDD.n2410 0.152939
R20920 VDD.n2412 VDD.n2411 0.152939
R20921 VDD.n2413 VDD.n2412 0.152939
R20922 VDD.n2414 VDD.n2413 0.152939
R20923 VDD.n2415 VDD.n2414 0.152939
R20924 VDD.n2416 VDD.n2415 0.152939
R20925 VDD.n2417 VDD.n2416 0.152939
R20926 VDD.n2418 VDD.n2417 0.152939
R20927 VDD.n2419 VDD.n2418 0.152939
R20928 VDD.n2422 VDD.n2419 0.152939
R20929 VDD.n2423 VDD.n2422 0.152939
R20930 VDD.n2424 VDD.n2423 0.152939
R20931 VDD.n2425 VDD.n2424 0.152939
R20932 VDD.n2426 VDD.n2425 0.152939
R20933 VDD.n2427 VDD.n2426 0.152939
R20934 VDD.n2428 VDD.n2427 0.152939
R20935 VDD.n2429 VDD.n2428 0.152939
R20936 VDD.n2430 VDD.n2429 0.152939
R20937 VDD.n2431 VDD.n2430 0.152939
R20938 VDD.n2431 VDD.n254 0.152939
R20939 VDD.n2475 VDD.n254 0.152939
R20940 VDD.n2483 VDD.n248 0.152939
R20941 VDD.n2484 VDD.n2483 0.152939
R20942 VDD.n2485 VDD.n2484 0.152939
R20943 VDD.n2485 VDD.n236 0.152939
R20944 VDD.n2499 VDD.n236 0.152939
R20945 VDD.n2500 VDD.n2499 0.152939
R20946 VDD.n2501 VDD.n2500 0.152939
R20947 VDD.n2501 VDD.n224 0.152939
R20948 VDD.n2515 VDD.n224 0.152939
R20949 VDD.n2516 VDD.n2515 0.152939
R20950 VDD.n2517 VDD.n2516 0.152939
R20951 VDD.n2517 VDD.n212 0.152939
R20952 VDD.n2531 VDD.n212 0.152939
R20953 VDD.n2532 VDD.n2531 0.152939
R20954 VDD.n2533 VDD.n2532 0.152939
R20955 VDD.n2533 VDD.n200 0.152939
R20956 VDD.n2547 VDD.n200 0.152939
R20957 VDD.n2548 VDD.n2547 0.152939
R20958 VDD.n2549 VDD.n2548 0.152939
R20959 VDD.n2549 VDD.n187 0.152939
R20960 VDD.n2566 VDD.n187 0.152939
R20961 VDD.n2567 VDD.n2566 0.152939
R20962 VDD.n2568 VDD.n2567 0.152939
R20963 VDD.n2568 VDD.n21 0.152939
R20964 VDD.n1064 VDD.n787 0.152939
R20965 VDD.n1065 VDD.n1064 0.152939
R20966 VDD.n1066 VDD.n1065 0.152939
R20967 VDD.n1066 VDD.n775 0.152939
R20968 VDD.n1080 VDD.n775 0.152939
R20969 VDD.n1081 VDD.n1080 0.152939
R20970 VDD.n1082 VDD.n1081 0.152939
R20971 VDD.n1082 VDD.n763 0.152939
R20972 VDD.n1096 VDD.n763 0.152939
R20973 VDD.n1097 VDD.n1096 0.152939
R20974 VDD.n1098 VDD.n1097 0.152939
R20975 VDD.n1098 VDD.n751 0.152939
R20976 VDD.n1112 VDD.n751 0.152939
R20977 VDD.n1113 VDD.n1112 0.152939
R20978 VDD.n1114 VDD.n1113 0.152939
R20979 VDD.n1114 VDD.n739 0.152939
R20980 VDD.n1128 VDD.n739 0.152939
R20981 VDD.n1129 VDD.n1128 0.152939
R20982 VDD.n1130 VDD.n1129 0.152939
R20983 VDD.n1130 VDD.n727 0.152939
R20984 VDD.n1145 VDD.n727 0.152939
R20985 VDD.n1146 VDD.n1145 0.152939
R20986 VDD.n1211 VDD.n1146 0.152939
R20987 VDD.n1211 VDD.n1210 0.152939
R20988 VDD.n1209 VDD.n1147 0.152939
R20989 VDD.n1205 VDD.n1147 0.152939
R20990 VDD.n1205 VDD.n1204 0.152939
R20991 VDD.n1204 VDD.n1203 0.152939
R20992 VDD.n1203 VDD.n1152 0.152939
R20993 VDD.n1199 VDD.n1152 0.152939
R20994 VDD.n1199 VDD.n1198 0.152939
R20995 VDD.n1198 VDD.n1197 0.152939
R20996 VDD.n1197 VDD.n1158 0.152939
R20997 VDD.n1193 VDD.n1158 0.152939
R20998 VDD.n1193 VDD.n1192 0.152939
R20999 VDD.n1192 VDD.n1191 0.152939
R21000 VDD.n1191 VDD.n1166 0.152939
R21001 VDD.n1187 VDD.n1166 0.152939
R21002 VDD.n1187 VDD.n1186 0.152939
R21003 VDD.n1186 VDD.n1185 0.152939
R21004 VDD.n1185 VDD.n1172 0.152939
R21005 VDD.n1181 VDD.n1172 0.152939
R21006 VDD.n1181 VDD.n1180 0.152939
R21007 VDD.n1180 VDD.n718 0.152939
R21008 VDD.n1219 VDD.n718 0.152939
R21009 VDD.n953 VDD.n952 0.152939
R21010 VDD.n954 VDD.n953 0.152939
R21011 VDD.n954 VDD.n852 0.152939
R21012 VDD.n968 VDD.n852 0.152939
R21013 VDD.n969 VDD.n968 0.152939
R21014 VDD.n970 VDD.n969 0.152939
R21015 VDD.n970 VDD.n840 0.152939
R21016 VDD.n984 VDD.n840 0.152939
R21017 VDD.n985 VDD.n984 0.152939
R21018 VDD.n986 VDD.n985 0.152939
R21019 VDD.n986 VDD.n828 0.152939
R21020 VDD.n1000 VDD.n828 0.152939
R21021 VDD.n1001 VDD.n1000 0.152939
R21022 VDD.n1002 VDD.n1001 0.152939
R21023 VDD.n1002 VDD.n817 0.152939
R21024 VDD.n1017 VDD.n817 0.152939
R21025 VDD.n1018 VDD.n1017 0.152939
R21026 VDD.n1019 VDD.n1018 0.152939
R21027 VDD.n1019 VDD.n805 0.152939
R21028 VDD.n1033 VDD.n805 0.152939
R21029 VDD.n1034 VDD.n1033 0.152939
R21030 VDD.n1035 VDD.n1034 0.152939
R21031 VDD.n1035 VDD.n793 0.152939
R21032 VDD.n1056 VDD.n793 0.152939
R21033 VDD.n1057 VDD.n1056 0.152939
R21034 VDD.n1058 VDD.n1057 0.152939
R21035 VDD.n1058 VDD.n781 0.152939
R21036 VDD.n1072 VDD.n781 0.152939
R21037 VDD.n1073 VDD.n1072 0.152939
R21038 VDD.n1074 VDD.n1073 0.152939
R21039 VDD.n1074 VDD.n768 0.152939
R21040 VDD.n1088 VDD.n768 0.152939
R21041 VDD.n1089 VDD.n1088 0.152939
R21042 VDD.n1090 VDD.n1089 0.152939
R21043 VDD.n1090 VDD.n757 0.152939
R21044 VDD.n1104 VDD.n757 0.152939
R21045 VDD.n1105 VDD.n1104 0.152939
R21046 VDD.n1106 VDD.n1105 0.152939
R21047 VDD.n1106 VDD.n745 0.152939
R21048 VDD.n1120 VDD.n745 0.152939
R21049 VDD.n1121 VDD.n1120 0.152939
R21050 VDD.n1122 VDD.n1121 0.152939
R21051 VDD.n1122 VDD.n733 0.152939
R21052 VDD.n1136 VDD.n733 0.152939
R21053 VDD.n1137 VDD.n1136 0.152939
R21054 VDD.n1139 VDD.n1137 0.152939
R21055 VDD.n1139 VDD.n1138 0.152939
R21056 VDD.n1138 VDD.n719 0.152939
R21057 VDD.n1218 VDD.n719 0.152939
R21058 VDD.n945 VDD.n868 0.152939
R21059 VDD.n941 VDD.n868 0.152939
R21060 VDD.n941 VDD.n940 0.152939
R21061 VDD.n940 VDD.n939 0.152939
R21062 VDD.n939 VDD.n873 0.152939
R21063 VDD.n935 VDD.n873 0.152939
R21064 VDD.n935 VDD.n934 0.152939
R21065 VDD.n934 VDD.n933 0.152939
R21066 VDD.n933 VDD.n881 0.152939
R21067 VDD.n888 VDD.n881 0.152939
R21068 VDD.n923 VDD.n888 0.152939
R21069 VDD.n923 VDD.n922 0.152939
R21070 VDD.n922 VDD.n921 0.152939
R21071 VDD.n921 VDD.n889 0.152939
R21072 VDD.n917 VDD.n889 0.152939
R21073 VDD.n917 VDD.n916 0.152939
R21074 VDD.n916 VDD.n915 0.152939
R21075 VDD.n915 VDD.n896 0.152939
R21076 VDD.n911 VDD.n896 0.152939
R21077 VDD.n911 VDD.n910 0.152939
R21078 VDD.n910 VDD.n864 0.152939
R21079 VDD.n946 VDD.n858 0.152939
R21080 VDD.n960 VDD.n858 0.152939
R21081 VDD.n961 VDD.n960 0.152939
R21082 VDD.n962 VDD.n961 0.152939
R21083 VDD.n962 VDD.n846 0.152939
R21084 VDD.n976 VDD.n846 0.152939
R21085 VDD.n977 VDD.n976 0.152939
R21086 VDD.n978 VDD.n977 0.152939
R21087 VDD.n978 VDD.n834 0.152939
R21088 VDD.n992 VDD.n834 0.152939
R21089 VDD.n993 VDD.n992 0.152939
R21090 VDD.n994 VDD.n993 0.152939
R21091 VDD.n994 VDD.n822 0.152939
R21092 VDD.n1009 VDD.n822 0.152939
R21093 VDD.n1010 VDD.n1009 0.152939
R21094 VDD.n1011 VDD.n1010 0.152939
R21095 VDD.n1011 VDD.n811 0.152939
R21096 VDD.n1025 VDD.n811 0.152939
R21097 VDD.n1026 VDD.n1025 0.152939
R21098 VDD.n1027 VDD.n1026 0.152939
R21099 VDD.n1027 VDD.n799 0.152939
R21100 VDD.n1041 VDD.n799 0.152939
R21101 VDD.n1042 VDD.n1041 0.152939
R21102 VDD.n1050 VDD.n1042 0.152939
R21103 VDD.n2676 VDD.n21 0.0695946
R21104 VDD.n2676 VDD.n2675 0.0695946
R21105 VDD.n1049 VDD.n787 0.0695946
R21106 VDD.n1050 VDD.n1049 0.0695946
R21107 VDD VDD.n15 0.00833333
R21108 a_n6715_8686.n44 a_n6715_8686.n41 756.745
R21109 a_n6715_8686.n60 a_n6715_8686.n38 756.745
R21110 a_n6715_8686.n45 a_n6715_8686.n44 585
R21111 a_n6715_8686.n43 a_n6715_8686.n13 585
R21112 a_n6715_8686.n25 a_n6715_8686.n24 585
R21113 a_n6715_8686.n31 a_n6715_8686.n42 585
R21114 a_n6715_8686.n7 a_n6715_8686.n6 113.853
R21115 a_n6715_8686.n60 a_n6715_8686.n59 585
R21116 a_n6715_8686.n15 a_n6715_8686.n61 585
R21117 a_n6715_8686.n27 a_n6715_8686.n26 585
R21118 a_n6715_8686.n62 a_n6715_8686.n32 585
R21119 a_n6715_8686.n8 a_n6715_8686.n9 113.853
R21120 a_n6715_8686.n44 a_n6715_8686.n43 171.744
R21121 a_n6715_8686.n43 a_n6715_8686.n24 171.744
R21122 a_n6715_8686.n42 a_n6715_8686.n24 171.744
R21123 a_n6715_8686.n61 a_n6715_8686.n60 171.744
R21124 a_n6715_8686.n61 a_n6715_8686.n26 171.744
R21125 a_n6715_8686.n62 a_n6715_8686.n26 171.744
R21126 a_n6715_8686.n10 a_n6715_8686.n0 4.72074
R21127 a_n6715_8686.n7 a_n6715_8686.n42 302.252
R21128 a_n6715_8686.n9 a_n6715_8686.n62 302.252
R21129 a_n6715_8686.n48 a_n6715_8686.t15 84.4322
R21130 a_n6715_8686.n56 a_n6715_8686.t11 81.234
R21131 a_n6715_8686.n22 a_n6715_8686.n23 2.62682
R21132 a_n6715_8686.n18 a_n6715_8686.n19 2.62682
R21133 a_n6715_8686.n20 a_n6715_8686.n21 2.62682
R21134 a_n6715_8686.n28 a_n6715_8686.t16 77.7261
R21135 a_n6715_8686.n39 a_n6715_8686.t1 77.7101
R21136 a_n6715_8686.n39 a_n6715_8686.t0 77.7101
R21137 a_n6715_8686.n28 a_n6715_8686.t2 75.5974
R21138 a_n6715_8686.n28 a_n6715_8686.n39 45.9241
R21139 a_n6715_8686.n11 a_n6715_8686.t23 70.1789
R21140 a_n6715_8686.n55 a_n6715_8686.t20 37.8617
R21141 a_n6715_8686.n3 a_n6715_8686.t39 67.0046
R21142 a_n6715_8686.n0 a_n6715_8686.t29 70.1786
R21143 a_n6715_8686.n29 a_n6715_8686.t30 70.1789
R21144 a_n6715_8686.n54 a_n6715_8686.t41 37.8617
R21145 a_n6715_8686.n2 a_n6715_8686.t38 67.0046
R21146 a_n6715_8686.n0 a_n6715_8686.t35 70.1786
R21147 a_n6715_8686.n12 a_n6715_8686.t28 70.1789
R21148 a_n6715_8686.n53 a_n6715_8686.t24 37.8617
R21149 a_n6715_8686.n1 a_n6715_8686.t33 67.0046
R21150 a_n6715_8686.n0 a_n6715_8686.t26 70.1786
R21151 a_n6715_8686.n30 a_n6715_8686.t25 70.1789
R21152 a_n6715_8686.n52 a_n6715_8686.t32 37.8617
R21153 a_n6715_8686.n51 a_n6715_8686.t34 37.8617
R21154 a_n6715_8686.n36 a_n6715_8686.t36 70.1786
R21155 a_n6715_8686.n40 a_n6715_8686.t37 37.8617
R21156 a_n6715_8686.n33 a_n6715_8686.t40 69.3753
R21157 a_n6715_8686.n23 a_n6715_8686.t27 70.5932
R21158 a_n6715_8686.n5 a_n6715_8686.t4 74.8407
R21159 a_n6715_8686.n5 a_n6715_8686.t8 65.7508
R21160 a_n6715_8686.n4 a_n6715_8686.t10 70.5935
R21161 a_n6715_8686.n49 a_n6715_8686.t6 37.8617
R21162 a_n6715_8686.n35 a_n6715_8686.t14 69.3753
R21163 a_n6715_8686.n19 a_n6715_8686.t12 70.5932
R21164 a_n6715_8686.n50 a_n6715_8686.t21 37.8617
R21165 a_n6715_8686.n34 a_n6715_8686.t22 69.3753
R21166 a_n6715_8686.n21 a_n6715_8686.t31 70.5932
R21167 a_n6715_8686.n57 a_n6715_8686.n56 35.9654
R21168 a_n6715_8686.n48 a_n6715_8686.n47 32.7672
R21169 a_n6715_8686.n55 a_n6715_8686.n11 69.6071
R21170 a_n6715_8686.n3 a_n6715_8686.n55 55.5075
R21171 a_n6715_8686.n54 a_n6715_8686.n29 69.6071
R21172 a_n6715_8686.n2 a_n6715_8686.n54 55.5075
R21173 a_n6715_8686.n53 a_n6715_8686.n12 69.6071
R21174 a_n6715_8686.n1 a_n6715_8686.n53 55.5075
R21175 a_n6715_8686.n10 a_n6715_8686.n52 53.5307
R21176 a_n6715_8686.n33 a_n6715_8686.n40 74.8603
R21177 a_n6715_8686.n40 a_n6715_8686.n23 50.3
R21178 a_n6715_8686.n4 a_n6715_8686.n5 3.67326
R21179 a_n6715_8686.n49 a_n6715_8686.n35 74.8603
R21180 a_n6715_8686.n19 a_n6715_8686.n49 50.3
R21181 a_n6715_8686.n50 a_n6715_8686.n34 74.8603
R21182 a_n6715_8686.n21 a_n6715_8686.n50 50.3
R21183 a_n6715_8686.n0 a_n6715_8686.n1 2.57076
R21184 a_n6715_8686.n30 a_n6715_8686.n52 69.6071
R21185 a_n6715_8686.n36 a_n6715_8686.n51 69.6074
R21186 a_n6715_8686.n22 a_n6715_8686.n17 15.9867
R21187 a_n6715_8686.n20 a_n6715_8686.n37 15.9715
R21188 a_n6715_8686.n17 a_n6715_8686.n48 15.5739
R21189 a_n6715_8686.n37 a_n6715_8686.n4 14.9601
R21190 a_n6715_8686.n56 a_n6715_8686.n37 14.7893
R21191 a_n6715_8686.n17 a_n6715_8686.n18 12.5738
R21192 a_n6715_8686.n31 a_n6715_8686.n6 4.008
R21193 a_n6715_8686.n32 a_n6715_8686.n8 4.008
R21194 a_n6715_8686.n31 a_n6715_8686.n25 11.249
R21195 a_n6715_8686.n32 a_n6715_8686.n27 11.249
R21196 a_n6715_8686.n13 a_n6715_8686.n14 3.79806
R21197 a_n6715_8686.n16 a_n6715_8686.n15 3.79806
R21198 a_n6715_8686.n45 a_n6715_8686.n13 9.69747
R21199 a_n6715_8686.n59 a_n6715_8686.n15 9.69747
R21200 a_n6715_8686.n47 a_n6715_8686.n6 9.45567
R21201 a_n6715_8686.n8 a_n6715_8686.n57 9.45567
R21202 a_n6715_8686.n6 a_n6715_8686.n46 9.3005
R21203 a_n6715_8686.n58 a_n6715_8686.n8 9.3005
R21204 a_n6715_8686.n46 a_n6715_8686.n41 8.92171
R21205 a_n6715_8686.n58 a_n6715_8686.n38 8.92171
R21206 a_n6715_8686.n4 a_n6715_8686.n22 6.62054
R21207 a_n6715_8686.n18 a_n6715_8686.n20 6.62054
R21208 a_n6715_8686.t11 a_n6715_8686.t9 6.12197
R21209 a_n6715_8686.t15 a_n6715_8686.t7 6.12197
R21210 a_n6715_8686.n10 a_n6715_8686.n51 53.5304
R21211 a_n6715_8686.n47 a_n6715_8686.n41 5.04292
R21212 a_n6715_8686.n57 a_n6715_8686.n38 5.04292
R21213 a_n6715_8686.t16 a_n6715_8686.t3 5.01316
R21214 a_n6715_8686.t2 a_n6715_8686.t19 5.01316
R21215 a_n6715_8686.t1 a_n6715_8686.t18 5.01316
R21216 a_n6715_8686.t0 a_n6715_8686.t17 5.01316
R21217 a_n6715_8686.n46 a_n6715_8686.n45 4.26717
R21218 a_n6715_8686.n59 a_n6715_8686.n58 4.26717
R21219 a_n6715_8686.n7 a_n6715_8686.t13 70.7672
R21220 a_n6715_8686.t5 a_n6715_8686.n9 70.7672
R21221 a_n6715_8686.n4 a_n6715_8686.n28 25.9906
R21222 a_n6715_8686.n14 a_n6715_8686.n6 4.35729
R21223 a_n6715_8686.n16 a_n6715_8686.n8 4.35729
R21224 a_n6715_8686.n16 a_n6715_8686.n27 3.56777
R21225 a_n6715_8686.n25 a_n6715_8686.n14 3.56777
R21226 a_n6715_8686.n17 a_n6715_8686.n0 10.3276
R21227 a_n6715_8686.n0 a_n6715_8686.n30 9.88709
R21228 a_n6715_8686.n0 a_n6715_8686.n3 8.82765
R21229 a_n6715_8686.n0 a_n6715_8686.n2 8.82765
R21230 a_n6715_8686.n12 a_n6715_8686.n0 8.31641
R21231 a_n6715_8686.n11 a_n6715_8686.n0 8.2638
R21232 a_n6715_8686.n0 a_n6715_8686.n37 7.95635
R21233 a_n6715_8686.n29 a_n6715_8686.n0 7.34713
R21234 a_n6715_8686.n0 a_n6715_8686.n36 7.34713
R21235 a_n6715_8686.n22 a_n6715_8686.n33 7.26955
R21236 a_n6715_8686.n20 a_n6715_8686.n34 7.26955
R21237 a_n6715_8686.n18 a_n6715_8686.n35 7.26955
R21238 a_n6793_8883.n131 a_n6793_8883.n118 756.745
R21239 a_n6793_8883.n74 a_n6793_8883.n61 756.745
R21240 a_n6793_8883.n56 a_n6793_8883.n43 756.745
R21241 a_n6793_8883.n37 a_n6793_8883.n24 756.745
R21242 a_n6793_8883.n92 a_n6793_8883.n79 756.745
R21243 a_n6793_8883.n111 a_n6793_8883.n98 756.745
R21244 a_n6793_8883.n132 a_n6793_8883.n131 585
R21245 a_n6793_8883.n130 a_n6793_8883.n129 585
R21246 a_n6793_8883.n121 a_n6793_8883.n120 585
R21247 a_n6793_8883.n126 a_n6793_8883.n125 585
R21248 a_n6793_8883.n124 a_n6793_8883.n123 585
R21249 a_n6793_8883.n7 a_n6793_8883.n6 585
R21250 a_n6793_8883.n75 a_n6793_8883.n74 585
R21251 a_n6793_8883.n73 a_n6793_8883.n72 585
R21252 a_n6793_8883.n64 a_n6793_8883.n63 585
R21253 a_n6793_8883.n69 a_n6793_8883.n68 585
R21254 a_n6793_8883.n67 a_n6793_8883.n66 585
R21255 a_n6793_8883.n10 a_n6793_8883.n9 585
R21256 a_n6793_8883.n57 a_n6793_8883.n56 585
R21257 a_n6793_8883.n55 a_n6793_8883.n54 585
R21258 a_n6793_8883.n46 a_n6793_8883.n45 585
R21259 a_n6793_8883.n51 a_n6793_8883.n50 585
R21260 a_n6793_8883.n49 a_n6793_8883.n48 585
R21261 a_n6793_8883.n13 a_n6793_8883.n12 585
R21262 a_n6793_8883.n38 a_n6793_8883.n37 585
R21263 a_n6793_8883.n36 a_n6793_8883.n35 585
R21264 a_n6793_8883.n27 a_n6793_8883.n26 585
R21265 a_n6793_8883.n32 a_n6793_8883.n31 585
R21266 a_n6793_8883.n30 a_n6793_8883.n29 585
R21267 a_n6793_8883.n16 a_n6793_8883.n15 585
R21268 a_n6793_8883.n93 a_n6793_8883.n92 585
R21269 a_n6793_8883.n91 a_n6793_8883.n90 585
R21270 a_n6793_8883.n82 a_n6793_8883.n81 585
R21271 a_n6793_8883.n87 a_n6793_8883.n86 585
R21272 a_n6793_8883.n85 a_n6793_8883.n84 585
R21273 a_n6793_8883.n19 a_n6793_8883.n18 585
R21274 a_n6793_8883.n112 a_n6793_8883.n111 585
R21275 a_n6793_8883.n110 a_n6793_8883.n109 585
R21276 a_n6793_8883.n101 a_n6793_8883.n100 585
R21277 a_n6793_8883.n106 a_n6793_8883.n105 585
R21278 a_n6793_8883.n104 a_n6793_8883.n103 585
R21279 a_n6793_8883.n22 a_n6793_8883.n21 585
R21280 a_n6793_8883.n131 a_n6793_8883.n130 171.744
R21281 a_n6793_8883.n130 a_n6793_8883.n120 171.744
R21282 a_n6793_8883.n125 a_n6793_8883.n120 171.744
R21283 a_n6793_8883.n125 a_n6793_8883.n124 171.744
R21284 a_n6793_8883.n124 a_n6793_8883.n6 171.744
R21285 a_n6793_8883.n74 a_n6793_8883.n73 171.744
R21286 a_n6793_8883.n73 a_n6793_8883.n63 171.744
R21287 a_n6793_8883.n68 a_n6793_8883.n63 171.744
R21288 a_n6793_8883.n68 a_n6793_8883.n67 171.744
R21289 a_n6793_8883.n67 a_n6793_8883.n9 171.744
R21290 a_n6793_8883.n56 a_n6793_8883.n55 171.744
R21291 a_n6793_8883.n55 a_n6793_8883.n45 171.744
R21292 a_n6793_8883.n50 a_n6793_8883.n45 171.744
R21293 a_n6793_8883.n50 a_n6793_8883.n49 171.744
R21294 a_n6793_8883.n49 a_n6793_8883.n12 171.744
R21295 a_n6793_8883.n37 a_n6793_8883.n36 171.744
R21296 a_n6793_8883.n36 a_n6793_8883.n26 171.744
R21297 a_n6793_8883.n31 a_n6793_8883.n26 171.744
R21298 a_n6793_8883.n31 a_n6793_8883.n30 171.744
R21299 a_n6793_8883.n30 a_n6793_8883.n15 171.744
R21300 a_n6793_8883.n92 a_n6793_8883.n91 171.744
R21301 a_n6793_8883.n91 a_n6793_8883.n81 171.744
R21302 a_n6793_8883.n86 a_n6793_8883.n81 171.744
R21303 a_n6793_8883.n86 a_n6793_8883.n85 171.744
R21304 a_n6793_8883.n85 a_n6793_8883.n18 171.744
R21305 a_n6793_8883.n111 a_n6793_8883.n110 171.744
R21306 a_n6793_8883.n110 a_n6793_8883.n100 171.744
R21307 a_n6793_8883.n105 a_n6793_8883.n100 171.744
R21308 a_n6793_8883.n105 a_n6793_8883.n104 171.744
R21309 a_n6793_8883.n104 a_n6793_8883.n21 171.744
R21310 a_n6793_8883.n116 a_n6793_8883.n115 97.9127
R21311 a_n6793_8883.n97 a_n6793_8883.n96 97.9126
R21312 a_n6793_8883.t5 a_n6793_8883.n6 85.8723
R21313 a_n6793_8883.t6 a_n6793_8883.n9 85.8723
R21314 a_n6793_8883.t3 a_n6793_8883.n12 85.8723
R21315 a_n6793_8883.t4 a_n6793_8883.n15 85.8723
R21316 a_n6793_8883.t13 a_n6793_8883.n18 85.8723
R21317 a_n6793_8883.t12 a_n6793_8883.n21 85.8723
R21318 a_n6793_8883.n42 a_n6793_8883.n41 81.234
R21319 a_n6793_8883.n137 a_n6793_8883.n136 81.234
R21320 a_n6793_8883.n97 a_n6793_8883.n95 52.6442
R21321 a_n6793_8883.n116 a_n6793_8883.n114 50.5501
R21322 a_n6793_8883.n42 a_n6793_8883.n40 35.9654
R21323 a_n6793_8883.n135 a_n6793_8883.n134 32.7672
R21324 a_n6793_8883.n78 a_n6793_8883.n77 32.7672
R21325 a_n6793_8883.n60 a_n6793_8883.n59 32.7672
R21326 a_n6793_8883.n117 a_n6793_8883.n116 28.4731
R21327 a_n6793_8883.n117 a_n6793_8883.n97 18.6546
R21328 a_n6793_8883.n8 a_n6793_8883.n7 5.32867
R21329 a_n6793_8883.n11 a_n6793_8883.n10 5.32867
R21330 a_n6793_8883.n14 a_n6793_8883.n13 5.32867
R21331 a_n6793_8883.n17 a_n6793_8883.n16 5.32867
R21332 a_n6793_8883.n20 a_n6793_8883.n19 5.32867
R21333 a_n6793_8883.n23 a_n6793_8883.n22 5.32867
R21334 a_n6793_8883.n123 a_n6793_8883.n7 12.8005
R21335 a_n6793_8883.n66 a_n6793_8883.n10 12.8005
R21336 a_n6793_8883.n48 a_n6793_8883.n13 12.8005
R21337 a_n6793_8883.n29 a_n6793_8883.n16 12.8005
R21338 a_n6793_8883.n84 a_n6793_8883.n19 12.8005
R21339 a_n6793_8883.n103 a_n6793_8883.n22 12.8005
R21340 a_n6793_8883.n126 a_n6793_8883.n122 12.0247
R21341 a_n6793_8883.n69 a_n6793_8883.n65 12.0247
R21342 a_n6793_8883.n51 a_n6793_8883.n47 12.0247
R21343 a_n6793_8883.n32 a_n6793_8883.n28 12.0247
R21344 a_n6793_8883.n87 a_n6793_8883.n83 12.0247
R21345 a_n6793_8883.n106 a_n6793_8883.n102 12.0247
R21346 a_n6793_8883.n127 a_n6793_8883.n121 11.249
R21347 a_n6793_8883.n70 a_n6793_8883.n64 11.249
R21348 a_n6793_8883.n52 a_n6793_8883.n46 11.249
R21349 a_n6793_8883.n33 a_n6793_8883.n27 11.249
R21350 a_n6793_8883.n88 a_n6793_8883.n82 11.249
R21351 a_n6793_8883.n107 a_n6793_8883.n101 11.249
R21352 a_n6793_8883.n129 a_n6793_8883.n128 10.4732
R21353 a_n6793_8883.n72 a_n6793_8883.n71 10.4732
R21354 a_n6793_8883.n54 a_n6793_8883.n53 10.4732
R21355 a_n6793_8883.n35 a_n6793_8883.n34 10.4732
R21356 a_n6793_8883.n90 a_n6793_8883.n89 10.4732
R21357 a_n6793_8883.n109 a_n6793_8883.n108 10.4732
R21358 a_n6793_8883.n132 a_n6793_8883.n119 9.69747
R21359 a_n6793_8883.n75 a_n6793_8883.n62 9.69747
R21360 a_n6793_8883.n57 a_n6793_8883.n44 9.69747
R21361 a_n6793_8883.n38 a_n6793_8883.n25 9.69747
R21362 a_n6793_8883.n93 a_n6793_8883.n80 9.69747
R21363 a_n6793_8883.n112 a_n6793_8883.n99 9.69747
R21364 a_n6793_8883.n134 a_n6793_8883.n0 9.45567
R21365 a_n6793_8883.n77 a_n6793_8883.n1 9.45567
R21366 a_n6793_8883.n59 a_n6793_8883.n2 9.45567
R21367 a_n6793_8883.n40 a_n6793_8883.n3 9.45567
R21368 a_n6793_8883.n95 a_n6793_8883.n4 9.45567
R21369 a_n6793_8883.n114 a_n6793_8883.n5 9.45567
R21370 a_n6793_8883.n0 a_n6793_8883.n133 9.3005
R21371 a_n6793_8883.n119 a_n6793_8883.n0 9.3005
R21372 a_n6793_8883.n128 a_n6793_8883.n0 9.3005
R21373 a_n6793_8883.n0 a_n6793_8883.n127 9.3005
R21374 a_n6793_8883.n122 a_n6793_8883.n0 9.3005
R21375 a_n6793_8883.n1 a_n6793_8883.n76 9.3005
R21376 a_n6793_8883.n62 a_n6793_8883.n1 9.3005
R21377 a_n6793_8883.n71 a_n6793_8883.n1 9.3005
R21378 a_n6793_8883.n1 a_n6793_8883.n70 9.3005
R21379 a_n6793_8883.n65 a_n6793_8883.n1 9.3005
R21380 a_n6793_8883.n2 a_n6793_8883.n58 9.3005
R21381 a_n6793_8883.n44 a_n6793_8883.n2 9.3005
R21382 a_n6793_8883.n53 a_n6793_8883.n2 9.3005
R21383 a_n6793_8883.n2 a_n6793_8883.n52 9.3005
R21384 a_n6793_8883.n47 a_n6793_8883.n2 9.3005
R21385 a_n6793_8883.n3 a_n6793_8883.n39 9.3005
R21386 a_n6793_8883.n25 a_n6793_8883.n3 9.3005
R21387 a_n6793_8883.n34 a_n6793_8883.n3 9.3005
R21388 a_n6793_8883.n3 a_n6793_8883.n33 9.3005
R21389 a_n6793_8883.n28 a_n6793_8883.n3 9.3005
R21390 a_n6793_8883.n4 a_n6793_8883.n94 9.3005
R21391 a_n6793_8883.n80 a_n6793_8883.n4 9.3005
R21392 a_n6793_8883.n89 a_n6793_8883.n4 9.3005
R21393 a_n6793_8883.n4 a_n6793_8883.n88 9.3005
R21394 a_n6793_8883.n83 a_n6793_8883.n4 9.3005
R21395 a_n6793_8883.n5 a_n6793_8883.n113 9.3005
R21396 a_n6793_8883.n99 a_n6793_8883.n5 9.3005
R21397 a_n6793_8883.n108 a_n6793_8883.n5 9.3005
R21398 a_n6793_8883.n5 a_n6793_8883.n107 9.3005
R21399 a_n6793_8883.n102 a_n6793_8883.n5 9.3005
R21400 a_n6793_8883.n133 a_n6793_8883.n118 8.92171
R21401 a_n6793_8883.n76 a_n6793_8883.n61 8.92171
R21402 a_n6793_8883.n58 a_n6793_8883.n43 8.92171
R21403 a_n6793_8883.n39 a_n6793_8883.n24 8.92171
R21404 a_n6793_8883.n94 a_n6793_8883.n79 8.92171
R21405 a_n6793_8883.n113 a_n6793_8883.n98 8.92171
R21406 a_n6793_8883.n135 a_n6793_8883.n117 7.08024
R21407 a_n6793_8883.n41 a_n6793_8883.t0 6.12197
R21408 a_n6793_8883.n41 a_n6793_8883.t2 6.12197
R21409 a_n6793_8883.n96 a_n6793_8883.t9 6.12197
R21410 a_n6793_8883.n96 a_n6793_8883.t8 6.12197
R21411 a_n6793_8883.n115 a_n6793_8883.t11 6.12197
R21412 a_n6793_8883.n115 a_n6793_8883.t10 6.12197
R21413 a_n6793_8883.t7 a_n6793_8883.n137 6.12197
R21414 a_n6793_8883.n137 a_n6793_8883.t1 6.12197
R21415 a_n6793_8883.n134 a_n6793_8883.n118 5.04292
R21416 a_n6793_8883.n77 a_n6793_8883.n61 5.04292
R21417 a_n6793_8883.n59 a_n6793_8883.n43 5.04292
R21418 a_n6793_8883.n40 a_n6793_8883.n24 5.04292
R21419 a_n6793_8883.n95 a_n6793_8883.n79 5.04292
R21420 a_n6793_8883.n114 a_n6793_8883.n98 5.04292
R21421 a_n6793_8883.n133 a_n6793_8883.n132 4.26717
R21422 a_n6793_8883.n76 a_n6793_8883.n75 4.26717
R21423 a_n6793_8883.n58 a_n6793_8883.n57 4.26717
R21424 a_n6793_8883.n39 a_n6793_8883.n38 4.26717
R21425 a_n6793_8883.n94 a_n6793_8883.n93 4.26717
R21426 a_n6793_8883.n113 a_n6793_8883.n112 4.26717
R21427 a_n6793_8883.n8 a_n6793_8883.t5 329.901
R21428 a_n6793_8883.n11 a_n6793_8883.t6 329.901
R21429 a_n6793_8883.n14 a_n6793_8883.t3 329.901
R21430 a_n6793_8883.n17 a_n6793_8883.t4 329.901
R21431 a_n6793_8883.n20 a_n6793_8883.t13 329.901
R21432 a_n6793_8883.n23 a_n6793_8883.t12 329.901
R21433 a_n6793_8883.n129 a_n6793_8883.n119 3.49141
R21434 a_n6793_8883.n72 a_n6793_8883.n62 3.49141
R21435 a_n6793_8883.n54 a_n6793_8883.n44 3.49141
R21436 a_n6793_8883.n35 a_n6793_8883.n25 3.49141
R21437 a_n6793_8883.n90 a_n6793_8883.n80 3.49141
R21438 a_n6793_8883.n109 a_n6793_8883.n99 3.49141
R21439 a_n6793_8883.n60 a_n6793_8883.n42 3.19878
R21440 a_n6793_8883.n136 a_n6793_8883.n78 3.19878
R21441 a_n6793_8883.n136 a_n6793_8883.n135 3.19878
R21442 a_n6793_8883.n128 a_n6793_8883.n121 2.71565
R21443 a_n6793_8883.n71 a_n6793_8883.n64 2.71565
R21444 a_n6793_8883.n53 a_n6793_8883.n46 2.71565
R21445 a_n6793_8883.n34 a_n6793_8883.n27 2.71565
R21446 a_n6793_8883.n89 a_n6793_8883.n82 2.71565
R21447 a_n6793_8883.n108 a_n6793_8883.n101 2.71565
R21448 a_n6793_8883.n23 a_n6793_8883.n5 1.98613
R21449 a_n6793_8883.n20 a_n6793_8883.n4 1.98613
R21450 a_n6793_8883.n17 a_n6793_8883.n3 1.98613
R21451 a_n6793_8883.n14 a_n6793_8883.n2 1.98613
R21452 a_n6793_8883.n11 a_n6793_8883.n1 1.98613
R21453 a_n6793_8883.n8 a_n6793_8883.n0 1.98613
R21454 a_n6793_8883.n127 a_n6793_8883.n126 1.93989
R21455 a_n6793_8883.n70 a_n6793_8883.n69 1.93989
R21456 a_n6793_8883.n52 a_n6793_8883.n51 1.93989
R21457 a_n6793_8883.n33 a_n6793_8883.n32 1.93989
R21458 a_n6793_8883.n88 a_n6793_8883.n87 1.93989
R21459 a_n6793_8883.n107 a_n6793_8883.n106 1.93989
R21460 a_n6793_8883.n123 a_n6793_8883.n122 1.16414
R21461 a_n6793_8883.n66 a_n6793_8883.n65 1.16414
R21462 a_n6793_8883.n48 a_n6793_8883.n47 1.16414
R21463 a_n6793_8883.n29 a_n6793_8883.n28 1.16414
R21464 a_n6793_8883.n84 a_n6793_8883.n83 1.16414
R21465 a_n6793_8883.n103 a_n6793_8883.n102 1.16414
R21466 a_n6793_8883.n78 a_n6793_8883.n60 0.819465
R21467 VP.n95 VP.t1 243.97
R21468 VP.n95 VP.t0 243.255
R21469 VP.n61 VP.n60 161.3
R21470 VP.n62 VP.n57 161.3
R21471 VP.n64 VP.n63 161.3
R21472 VP.n65 VP.n56 161.3
R21473 VP.n67 VP.n66 161.3
R21474 VP.n68 VP.n55 161.3
R21475 VP.n70 VP.n69 161.3
R21476 VP.n71 VP.n54 161.3
R21477 VP.n73 VP.n72 161.3
R21478 VP.n74 VP.n53 161.3
R21479 VP.n76 VP.n75 161.3
R21480 VP.n78 VP.n77 161.3
R21481 VP.n79 VP.n51 161.3
R21482 VP.n81 VP.n80 161.3
R21483 VP.n82 VP.n50 161.3
R21484 VP.n84 VP.n83 161.3
R21485 VP.n85 VP.n49 161.3
R21486 VP.n87 VP.n86 161.3
R21487 VP.n88 VP.n48 161.3
R21488 VP.n90 VP.n89 161.3
R21489 VP.n91 VP.n47 161.3
R21490 VP.n44 VP.n0 161.3
R21491 VP.n43 VP.n42 161.3
R21492 VP.n41 VP.n1 161.3
R21493 VP.n40 VP.n39 161.3
R21494 VP.n38 VP.n2 161.3
R21495 VP.n37 VP.n36 161.3
R21496 VP.n35 VP.n3 161.3
R21497 VP.n34 VP.n33 161.3
R21498 VP.n32 VP.n4 161.3
R21499 VP.n31 VP.n30 161.3
R21500 VP.n29 VP.n28 161.3
R21501 VP.n27 VP.n6 161.3
R21502 VP.n26 VP.n25 161.3
R21503 VP.n24 VP.n7 161.3
R21504 VP.n23 VP.n22 161.3
R21505 VP.n21 VP.n8 161.3
R21506 VP.n20 VP.n19 161.3
R21507 VP.n18 VP.n9 161.3
R21508 VP.n17 VP.n16 161.3
R21509 VP.n15 VP.n10 161.3
R21510 VP.n14 VP.n13 161.3
R21511 VP.n93 VP.n92 79.9798
R21512 VP.n46 VP.n45 79.9798
R21513 VP.n59 VP.n58 74.8596
R21514 VP.n12 VP.n11 74.8596
R21515 VP.n12 VP.t3 52.4204
R21516 VP.n59 VP.t8 52.4201
R21517 VP.n85 VP.n84 43.4072
R21518 VP.n38 VP.n37 43.4072
R21519 VP.n94 VP.n93 42.7409
R21520 VP.n69 VP.n68 40.4934
R21521 VP.n68 VP.n67 40.4934
R21522 VP.n21 VP.n20 40.4934
R21523 VP.n22 VP.n21 40.4934
R21524 VP.n84 VP.n50 37.5796
R21525 VP.n37 VP.n3 37.5796
R21526 VP.n91 VP.n90 24.4675
R21527 VP.n90 VP.n48 24.4675
R21528 VP.n86 VP.n48 24.4675
R21529 VP.n86 VP.n85 24.4675
R21530 VP.n80 VP.n50 24.4675
R21531 VP.n80 VP.n79 24.4675
R21532 VP.n79 VP.n78 24.4675
R21533 VP.n75 VP.n74 24.4675
R21534 VP.n74 VP.n73 24.4675
R21535 VP.n73 VP.n54 24.4675
R21536 VP.n69 VP.n54 24.4675
R21537 VP.n67 VP.n56 24.4675
R21538 VP.n63 VP.n56 24.4675
R21539 VP.n63 VP.n62 24.4675
R21540 VP.n62 VP.n61 24.4675
R21541 VP.n15 VP.n14 24.4675
R21542 VP.n16 VP.n15 24.4675
R21543 VP.n16 VP.n9 24.4675
R21544 VP.n20 VP.n9 24.4675
R21545 VP.n22 VP.n7 24.4675
R21546 VP.n26 VP.n7 24.4675
R21547 VP.n27 VP.n26 24.4675
R21548 VP.n28 VP.n27 24.4675
R21549 VP.n32 VP.n31 24.4675
R21550 VP.n33 VP.n32 24.4675
R21551 VP.n33 VP.n3 24.4675
R21552 VP.n39 VP.n38 24.4675
R21553 VP.n39 VP.n1 24.4675
R21554 VP.n43 VP.n1 24.4675
R21555 VP.n44 VP.n43 24.4675
R21556 VP.n78 VP.n52 23.7335
R21557 VP.n31 VP.n5 23.7335
R21558 VP.n92 VP.t2 20.2548
R21559 VP.n52 VP.t5 20.2548
R21560 VP.n58 VP.t9 20.2548
R21561 VP.n11 VP.t6 20.2548
R21562 VP.n5 VP.t4 20.2548
R21563 VP.n45 VP.t7 20.2548
R21564 VP VP.n96 13.2918
R21565 VP.n94 VP.n46 12.5288
R21566 VP.n96 VP.n95 4.80222
R21567 VP.n92 VP.n91 2.20253
R21568 VP.n45 VP.n44 2.20253
R21569 VP.n13 VP.n12 1.81424
R21570 VP.n60 VP.n59 1.81423
R21571 VP.n96 VP.n94 0.972091
R21572 VP.n75 VP.n52 0.73451
R21573 VP.n61 VP.n58 0.73451
R21574 VP.n14 VP.n11 0.73451
R21575 VP.n28 VP.n5 0.73451
R21576 VP.n93 VP.n47 0.417535
R21577 VP.n46 VP.n0 0.417535
R21578 VP.n89 VP.n47 0.189894
R21579 VP.n89 VP.n88 0.189894
R21580 VP.n88 VP.n87 0.189894
R21581 VP.n87 VP.n49 0.189894
R21582 VP.n83 VP.n49 0.189894
R21583 VP.n83 VP.n82 0.189894
R21584 VP.n82 VP.n81 0.189894
R21585 VP.n81 VP.n51 0.189894
R21586 VP.n77 VP.n51 0.189894
R21587 VP.n77 VP.n76 0.189894
R21588 VP.n76 VP.n53 0.189894
R21589 VP.n72 VP.n53 0.189894
R21590 VP.n72 VP.n71 0.189894
R21591 VP.n71 VP.n70 0.189894
R21592 VP.n70 VP.n55 0.189894
R21593 VP.n66 VP.n55 0.189894
R21594 VP.n66 VP.n65 0.189894
R21595 VP.n65 VP.n64 0.189894
R21596 VP.n64 VP.n57 0.189894
R21597 VP.n60 VP.n57 0.189894
R21598 VP.n13 VP.n10 0.189894
R21599 VP.n17 VP.n10 0.189894
R21600 VP.n18 VP.n17 0.189894
R21601 VP.n19 VP.n18 0.189894
R21602 VP.n19 VP.n8 0.189894
R21603 VP.n23 VP.n8 0.189894
R21604 VP.n24 VP.n23 0.189894
R21605 VP.n25 VP.n24 0.189894
R21606 VP.n25 VP.n6 0.189894
R21607 VP.n29 VP.n6 0.189894
R21608 VP.n30 VP.n29 0.189894
R21609 VP.n30 VP.n4 0.189894
R21610 VP.n34 VP.n4 0.189894
R21611 VP.n35 VP.n34 0.189894
R21612 VP.n36 VP.n35 0.189894
R21613 VP.n36 VP.n2 0.189894
R21614 VP.n40 VP.n2 0.189894
R21615 VP.n41 VP.n40 0.189894
R21616 VP.n42 VP.n41 0.189894
R21617 VP.n42 VP.n0 0.189894
R21618 a_n3792_7061.n133 a_n3792_7061.n120 756.745
R21619 a_n3792_7061.n115 a_n3792_7061.n102 756.745
R21620 a_n3792_7061.n97 a_n3792_7061.n84 756.745
R21621 a_n3792_7061.n77 a_n3792_7061.n64 756.745
R21622 a_n3792_7061.n37 a_n3792_7061.n24 756.745
R21623 a_n3792_7061.n57 a_n3792_7061.n44 756.745
R21624 a_n3792_7061.n134 a_n3792_7061.n133 585
R21625 a_n3792_7061.n132 a_n3792_7061.n131 585
R21626 a_n3792_7061.n123 a_n3792_7061.n122 585
R21627 a_n3792_7061.n128 a_n3792_7061.n127 585
R21628 a_n3792_7061.n126 a_n3792_7061.n125 585
R21629 a_n3792_7061.n7 a_n3792_7061.n6 585
R21630 a_n3792_7061.n116 a_n3792_7061.n115 585
R21631 a_n3792_7061.n114 a_n3792_7061.n113 585
R21632 a_n3792_7061.n105 a_n3792_7061.n104 585
R21633 a_n3792_7061.n110 a_n3792_7061.n109 585
R21634 a_n3792_7061.n108 a_n3792_7061.n107 585
R21635 a_n3792_7061.n10 a_n3792_7061.n9 585
R21636 a_n3792_7061.n98 a_n3792_7061.n97 585
R21637 a_n3792_7061.n96 a_n3792_7061.n95 585
R21638 a_n3792_7061.n87 a_n3792_7061.n86 585
R21639 a_n3792_7061.n92 a_n3792_7061.n91 585
R21640 a_n3792_7061.n90 a_n3792_7061.n89 585
R21641 a_n3792_7061.n13 a_n3792_7061.n12 585
R21642 a_n3792_7061.n78 a_n3792_7061.n77 585
R21643 a_n3792_7061.n76 a_n3792_7061.n75 585
R21644 a_n3792_7061.n67 a_n3792_7061.n66 585
R21645 a_n3792_7061.n72 a_n3792_7061.n71 585
R21646 a_n3792_7061.n70 a_n3792_7061.n69 585
R21647 a_n3792_7061.n16 a_n3792_7061.n15 585
R21648 a_n3792_7061.n38 a_n3792_7061.n37 585
R21649 a_n3792_7061.n36 a_n3792_7061.n35 585
R21650 a_n3792_7061.n27 a_n3792_7061.n26 585
R21651 a_n3792_7061.n32 a_n3792_7061.n31 585
R21652 a_n3792_7061.n30 a_n3792_7061.n29 585
R21653 a_n3792_7061.n19 a_n3792_7061.n18 585
R21654 a_n3792_7061.n58 a_n3792_7061.n57 585
R21655 a_n3792_7061.n56 a_n3792_7061.n55 585
R21656 a_n3792_7061.n47 a_n3792_7061.n46 585
R21657 a_n3792_7061.n52 a_n3792_7061.n51 585
R21658 a_n3792_7061.n50 a_n3792_7061.n49 585
R21659 a_n3792_7061.n22 a_n3792_7061.n21 585
R21660 a_n3792_7061.n133 a_n3792_7061.n132 171.744
R21661 a_n3792_7061.n132 a_n3792_7061.n122 171.744
R21662 a_n3792_7061.n127 a_n3792_7061.n122 171.744
R21663 a_n3792_7061.n127 a_n3792_7061.n126 171.744
R21664 a_n3792_7061.n126 a_n3792_7061.n6 171.744
R21665 a_n3792_7061.n115 a_n3792_7061.n114 171.744
R21666 a_n3792_7061.n114 a_n3792_7061.n104 171.744
R21667 a_n3792_7061.n109 a_n3792_7061.n104 171.744
R21668 a_n3792_7061.n109 a_n3792_7061.n108 171.744
R21669 a_n3792_7061.n108 a_n3792_7061.n9 171.744
R21670 a_n3792_7061.n97 a_n3792_7061.n96 171.744
R21671 a_n3792_7061.n96 a_n3792_7061.n86 171.744
R21672 a_n3792_7061.n91 a_n3792_7061.n86 171.744
R21673 a_n3792_7061.n91 a_n3792_7061.n90 171.744
R21674 a_n3792_7061.n90 a_n3792_7061.n12 171.744
R21675 a_n3792_7061.n77 a_n3792_7061.n76 171.744
R21676 a_n3792_7061.n76 a_n3792_7061.n66 171.744
R21677 a_n3792_7061.n71 a_n3792_7061.n66 171.744
R21678 a_n3792_7061.n71 a_n3792_7061.n70 171.744
R21679 a_n3792_7061.n70 a_n3792_7061.n15 171.744
R21680 a_n3792_7061.n37 a_n3792_7061.n36 171.744
R21681 a_n3792_7061.n36 a_n3792_7061.n26 171.744
R21682 a_n3792_7061.n31 a_n3792_7061.n26 171.744
R21683 a_n3792_7061.n31 a_n3792_7061.n30 171.744
R21684 a_n3792_7061.n30 a_n3792_7061.n18 171.744
R21685 a_n3792_7061.n57 a_n3792_7061.n56 171.744
R21686 a_n3792_7061.n56 a_n3792_7061.n46 171.744
R21687 a_n3792_7061.n51 a_n3792_7061.n46 171.744
R21688 a_n3792_7061.n51 a_n3792_7061.n50 171.744
R21689 a_n3792_7061.n50 a_n3792_7061.n21 171.744
R21690 a_n3792_7061.t6 a_n3792_7061.n6 85.8723
R21691 a_n3792_7061.t5 a_n3792_7061.n9 85.8723
R21692 a_n3792_7061.t1 a_n3792_7061.n12 85.8723
R21693 a_n3792_7061.t7 a_n3792_7061.n15 85.8723
R21694 a_n3792_7061.t11 a_n3792_7061.n18 85.8723
R21695 a_n3792_7061.t12 a_n3792_7061.n21 85.8723
R21696 a_n3792_7061.n83 a_n3792_7061.n82 81.234
R21697 a_n3792_7061.n42 a_n3792_7061.n41 81.234
R21698 a_n3792_7061.n62 a_n3792_7061.n61 81.234
R21699 a_n3792_7061.n138 a_n3792_7061.n137 81.234
R21700 a_n3792_7061.n63 a_n3792_7061.n62 38.9042
R21701 a_n3792_7061.n137 a_n3792_7061.n136 35.9654
R21702 a_n3792_7061.n42 a_n3792_7061.n40 35.9654
R21703 a_n3792_7061.n62 a_n3792_7061.n60 35.9654
R21704 a_n3792_7061.n119 a_n3792_7061.n118 32.7672
R21705 a_n3792_7061.n101 a_n3792_7061.n100 32.7672
R21706 a_n3792_7061.n81 a_n3792_7061.n80 32.7672
R21707 a_n3792_7061.n8 a_n3792_7061.n7 5.32867
R21708 a_n3792_7061.n11 a_n3792_7061.n10 5.32867
R21709 a_n3792_7061.n14 a_n3792_7061.n13 5.32867
R21710 a_n3792_7061.n17 a_n3792_7061.n16 5.32867
R21711 a_n3792_7061.n20 a_n3792_7061.n19 5.32867
R21712 a_n3792_7061.n23 a_n3792_7061.n22 5.32867
R21713 a_n3792_7061.n43 a_n3792_7061.n42 15.1471
R21714 a_n3792_7061.n125 a_n3792_7061.n7 12.8005
R21715 a_n3792_7061.n107 a_n3792_7061.n10 12.8005
R21716 a_n3792_7061.n89 a_n3792_7061.n13 12.8005
R21717 a_n3792_7061.n69 a_n3792_7061.n16 12.8005
R21718 a_n3792_7061.n29 a_n3792_7061.n19 12.8005
R21719 a_n3792_7061.n49 a_n3792_7061.n22 12.8005
R21720 a_n3792_7061.n128 a_n3792_7061.n124 12.0247
R21721 a_n3792_7061.n110 a_n3792_7061.n106 12.0247
R21722 a_n3792_7061.n92 a_n3792_7061.n88 12.0247
R21723 a_n3792_7061.n72 a_n3792_7061.n68 12.0247
R21724 a_n3792_7061.n32 a_n3792_7061.n28 12.0247
R21725 a_n3792_7061.n52 a_n3792_7061.n48 12.0247
R21726 a_n3792_7061.n43 a_n3792_7061.t0 11.4334
R21727 a_n3792_7061.n129 a_n3792_7061.n123 11.249
R21728 a_n3792_7061.n111 a_n3792_7061.n105 11.249
R21729 a_n3792_7061.n93 a_n3792_7061.n87 11.249
R21730 a_n3792_7061.n73 a_n3792_7061.n67 11.249
R21731 a_n3792_7061.n33 a_n3792_7061.n27 11.249
R21732 a_n3792_7061.n53 a_n3792_7061.n47 11.249
R21733 a_n3792_7061.n131 a_n3792_7061.n130 10.4732
R21734 a_n3792_7061.n113 a_n3792_7061.n112 10.4732
R21735 a_n3792_7061.n95 a_n3792_7061.n94 10.4732
R21736 a_n3792_7061.n75 a_n3792_7061.n74 10.4732
R21737 a_n3792_7061.n35 a_n3792_7061.n34 10.4732
R21738 a_n3792_7061.n55 a_n3792_7061.n54 10.4732
R21739 a_n3792_7061.n134 a_n3792_7061.n121 9.69747
R21740 a_n3792_7061.n116 a_n3792_7061.n103 9.69747
R21741 a_n3792_7061.n98 a_n3792_7061.n85 9.69747
R21742 a_n3792_7061.n78 a_n3792_7061.n65 9.69747
R21743 a_n3792_7061.n38 a_n3792_7061.n25 9.69747
R21744 a_n3792_7061.n58 a_n3792_7061.n45 9.69747
R21745 a_n3792_7061.n136 a_n3792_7061.n0 9.45567
R21746 a_n3792_7061.n118 a_n3792_7061.n1 9.45567
R21747 a_n3792_7061.n100 a_n3792_7061.n2 9.45567
R21748 a_n3792_7061.n80 a_n3792_7061.n3 9.45567
R21749 a_n3792_7061.n40 a_n3792_7061.n4 9.45567
R21750 a_n3792_7061.n60 a_n3792_7061.n5 9.45567
R21751 a_n3792_7061.n0 a_n3792_7061.n135 9.3005
R21752 a_n3792_7061.n121 a_n3792_7061.n0 9.3005
R21753 a_n3792_7061.n130 a_n3792_7061.n0 9.3005
R21754 a_n3792_7061.n0 a_n3792_7061.n129 9.3005
R21755 a_n3792_7061.n124 a_n3792_7061.n0 9.3005
R21756 a_n3792_7061.n1 a_n3792_7061.n117 9.3005
R21757 a_n3792_7061.n103 a_n3792_7061.n1 9.3005
R21758 a_n3792_7061.n112 a_n3792_7061.n1 9.3005
R21759 a_n3792_7061.n1 a_n3792_7061.n111 9.3005
R21760 a_n3792_7061.n106 a_n3792_7061.n1 9.3005
R21761 a_n3792_7061.n2 a_n3792_7061.n99 9.3005
R21762 a_n3792_7061.n85 a_n3792_7061.n2 9.3005
R21763 a_n3792_7061.n94 a_n3792_7061.n2 9.3005
R21764 a_n3792_7061.n2 a_n3792_7061.n93 9.3005
R21765 a_n3792_7061.n88 a_n3792_7061.n2 9.3005
R21766 a_n3792_7061.n3 a_n3792_7061.n79 9.3005
R21767 a_n3792_7061.n65 a_n3792_7061.n3 9.3005
R21768 a_n3792_7061.n74 a_n3792_7061.n3 9.3005
R21769 a_n3792_7061.n3 a_n3792_7061.n73 9.3005
R21770 a_n3792_7061.n68 a_n3792_7061.n3 9.3005
R21771 a_n3792_7061.n4 a_n3792_7061.n39 9.3005
R21772 a_n3792_7061.n25 a_n3792_7061.n4 9.3005
R21773 a_n3792_7061.n34 a_n3792_7061.n4 9.3005
R21774 a_n3792_7061.n4 a_n3792_7061.n33 9.3005
R21775 a_n3792_7061.n28 a_n3792_7061.n4 9.3005
R21776 a_n3792_7061.n5 a_n3792_7061.n59 9.3005
R21777 a_n3792_7061.n45 a_n3792_7061.n5 9.3005
R21778 a_n3792_7061.n54 a_n3792_7061.n5 9.3005
R21779 a_n3792_7061.n5 a_n3792_7061.n53 9.3005
R21780 a_n3792_7061.n48 a_n3792_7061.n5 9.3005
R21781 a_n3792_7061.n135 a_n3792_7061.n120 8.92171
R21782 a_n3792_7061.n117 a_n3792_7061.n102 8.92171
R21783 a_n3792_7061.n99 a_n3792_7061.n84 8.92171
R21784 a_n3792_7061.n79 a_n3792_7061.n64 8.92171
R21785 a_n3792_7061.n39 a_n3792_7061.n24 8.92171
R21786 a_n3792_7061.n59 a_n3792_7061.n44 8.92171
R21787 a_n3792_7061.n81 a_n3792_7061.n63 7.08024
R21788 a_n3792_7061.n82 a_n3792_7061.t4 6.12197
R21789 a_n3792_7061.n82 a_n3792_7061.t2 6.12197
R21790 a_n3792_7061.n41 a_n3792_7061.t13 6.12197
R21791 a_n3792_7061.n41 a_n3792_7061.t14 6.12197
R21792 a_n3792_7061.n61 a_n3792_7061.t9 6.12197
R21793 a_n3792_7061.n61 a_n3792_7061.t10 6.12197
R21794 a_n3792_7061.t8 a_n3792_7061.n138 6.12197
R21795 a_n3792_7061.n138 a_n3792_7061.t3 6.12197
R21796 a_n3792_7061.n136 a_n3792_7061.n120 5.04292
R21797 a_n3792_7061.n118 a_n3792_7061.n102 5.04292
R21798 a_n3792_7061.n100 a_n3792_7061.n84 5.04292
R21799 a_n3792_7061.n80 a_n3792_7061.n64 5.04292
R21800 a_n3792_7061.n40 a_n3792_7061.n24 5.04292
R21801 a_n3792_7061.n60 a_n3792_7061.n44 5.04292
R21802 a_n3792_7061.n135 a_n3792_7061.n134 4.26717
R21803 a_n3792_7061.n117 a_n3792_7061.n116 4.26717
R21804 a_n3792_7061.n99 a_n3792_7061.n98 4.26717
R21805 a_n3792_7061.n79 a_n3792_7061.n78 4.26717
R21806 a_n3792_7061.n39 a_n3792_7061.n38 4.26717
R21807 a_n3792_7061.n59 a_n3792_7061.n58 4.26717
R21808 a_n3792_7061.n8 a_n3792_7061.t6 329.901
R21809 a_n3792_7061.n11 a_n3792_7061.t5 329.901
R21810 a_n3792_7061.n14 a_n3792_7061.t1 329.901
R21811 a_n3792_7061.n17 a_n3792_7061.t7 329.901
R21812 a_n3792_7061.n20 a_n3792_7061.t11 329.901
R21813 a_n3792_7061.n23 a_n3792_7061.t12 329.901
R21814 a_n3792_7061.n131 a_n3792_7061.n121 3.49141
R21815 a_n3792_7061.n113 a_n3792_7061.n103 3.49141
R21816 a_n3792_7061.n95 a_n3792_7061.n85 3.49141
R21817 a_n3792_7061.n75 a_n3792_7061.n65 3.49141
R21818 a_n3792_7061.n35 a_n3792_7061.n25 3.49141
R21819 a_n3792_7061.n55 a_n3792_7061.n45 3.49141
R21820 a_n3792_7061.n63 a_n3792_7061.n43 3.39823
R21821 a_n3792_7061.n83 a_n3792_7061.n81 3.19878
R21822 a_n3792_7061.n101 a_n3792_7061.n83 3.19878
R21823 a_n3792_7061.n137 a_n3792_7061.n119 3.19878
R21824 a_n3792_7061.n130 a_n3792_7061.n123 2.71565
R21825 a_n3792_7061.n112 a_n3792_7061.n105 2.71565
R21826 a_n3792_7061.n94 a_n3792_7061.n87 2.71565
R21827 a_n3792_7061.n74 a_n3792_7061.n67 2.71565
R21828 a_n3792_7061.n34 a_n3792_7061.n27 2.71565
R21829 a_n3792_7061.n54 a_n3792_7061.n47 2.71565
R21830 a_n3792_7061.n23 a_n3792_7061.n5 1.98613
R21831 a_n3792_7061.n20 a_n3792_7061.n4 1.98613
R21832 a_n3792_7061.n17 a_n3792_7061.n3 1.98613
R21833 a_n3792_7061.n14 a_n3792_7061.n2 1.98613
R21834 a_n3792_7061.n11 a_n3792_7061.n1 1.98613
R21835 a_n3792_7061.n8 a_n3792_7061.n0 1.98613
R21836 a_n3792_7061.n129 a_n3792_7061.n128 1.93989
R21837 a_n3792_7061.n111 a_n3792_7061.n110 1.93989
R21838 a_n3792_7061.n93 a_n3792_7061.n92 1.93989
R21839 a_n3792_7061.n73 a_n3792_7061.n72 1.93989
R21840 a_n3792_7061.n33 a_n3792_7061.n32 1.93989
R21841 a_n3792_7061.n53 a_n3792_7061.n52 1.93989
R21842 a_n3792_7061.n125 a_n3792_7061.n124 1.16414
R21843 a_n3792_7061.n107 a_n3792_7061.n106 1.16414
R21844 a_n3792_7061.n89 a_n3792_7061.n88 1.16414
R21845 a_n3792_7061.n69 a_n3792_7061.n68 1.16414
R21846 a_n3792_7061.n29 a_n3792_7061.n28 1.16414
R21847 a_n3792_7061.n49 a_n3792_7061.n48 1.16414
R21848 a_n3792_7061.n119 a_n3792_7061.n101 0.819465
R21849 a_n689_n2782.t0 a_n689_n2782.t1 273.49
C0 VDD VOUT 20.999699f
C1 a_n7753_8883# VDD 1.34259f
C2 VOUT VP 4.22106f
C3 VDD VN 0.180764f
C4 VOUT VN 1.12158f
C5 VP VN 13.8785f
C6 VOUT CS_BIAS 25.5071f
C7 VP CS_BIAS 0.387033f
C8 VP DIFFPAIR_BIAS 0.010921f
C9 VN CS_BIAS 0.313722f
C10 VN DIFFPAIR_BIAS 0.02354f
C11 a_6921_8883# VDD 1.34208f
C12 DIFFPAIR_BIAS GND 13.506898f
C13 CS_BIAS GND 0.191442p
C14 VN GND 47.124954f
C15 VP GND 38.89248f
C16 VOUT GND 79.60752f
C17 VDD GND 0.478517p
C18 a_6921_8883# GND 0.433531f
C19 a_n7753_8883# GND 0.433531f
C20 a_n689_n2782.t1 GND 1.35069f
C21 a_n689_n2782.t0 GND 1.34931f
C22 a_n3792_7061.n0 GND 0.319828f
C23 a_n3792_7061.n1 GND 0.319828f
C24 a_n3792_7061.n2 GND 0.319828f
C25 a_n3792_7061.n3 GND 0.319828f
C26 a_n3792_7061.n4 GND 0.319828f
C27 a_n3792_7061.n5 GND 0.319828f
C28 a_n3792_7061.n6 GND 0.011661f
C29 a_n3792_7061.n7 GND 0.016454f
C30 a_n3792_7061.n8 GND 0.051497f
C31 a_n3792_7061.n9 GND 0.011661f
C32 a_n3792_7061.n10 GND 0.016454f
C33 a_n3792_7061.n11 GND 0.051497f
C34 a_n3792_7061.n12 GND 0.011661f
C35 a_n3792_7061.n13 GND 0.016454f
C36 a_n3792_7061.n14 GND 0.051497f
C37 a_n3792_7061.n15 GND 0.011661f
C38 a_n3792_7061.n16 GND 0.016454f
C39 a_n3792_7061.n17 GND 0.051497f
C40 a_n3792_7061.n18 GND 0.011661f
C41 a_n3792_7061.n19 GND 0.016454f
C42 a_n3792_7061.n20 GND 0.051497f
C43 a_n3792_7061.n21 GND 0.011661f
C44 a_n3792_7061.n22 GND 0.016454f
C45 a_n3792_7061.n23 GND 0.051497f
C46 a_n3792_7061.t0 GND 51.314396f
C47 a_n3792_7061.n24 GND 0.013348f
C48 a_n3792_7061.n25 GND 0.006578f
C49 a_n3792_7061.n26 GND 0.015548f
C50 a_n3792_7061.n27 GND 0.006965f
C51 a_n3792_7061.n28 GND 0.006578f
C52 a_n3792_7061.t11 GND 0.033882f
C53 a_n3792_7061.n29 GND 0.006965f
C54 a_n3792_7061.n30 GND 0.015548f
C55 a_n3792_7061.n31 GND 0.015548f
C56 a_n3792_7061.n32 GND 0.006965f
C57 a_n3792_7061.n33 GND 0.006578f
C58 a_n3792_7061.n34 GND 0.006578f
C59 a_n3792_7061.n35 GND 0.006965f
C60 a_n3792_7061.n36 GND 0.015548f
C61 a_n3792_7061.n37 GND 0.037289f
C62 a_n3792_7061.n38 GND 0.006965f
C63 a_n3792_7061.n39 GND 0.006578f
C64 a_n3792_7061.n40 GND 0.031364f
C65 a_n3792_7061.t13 GND 0.051366f
C66 a_n3792_7061.t14 GND 0.051366f
C67 a_n3792_7061.n41 GND 0.289994f
C68 a_n3792_7061.n42 GND 1.01833f
C69 a_n3792_7061.n43 GND 5.21359f
C70 a_n3792_7061.n44 GND 0.013348f
C71 a_n3792_7061.n45 GND 0.006578f
C72 a_n3792_7061.n46 GND 0.015548f
C73 a_n3792_7061.n47 GND 0.006965f
C74 a_n3792_7061.n48 GND 0.006578f
C75 a_n3792_7061.t12 GND 0.033882f
C76 a_n3792_7061.n49 GND 0.006965f
C77 a_n3792_7061.n50 GND 0.015548f
C78 a_n3792_7061.n51 GND 0.015548f
C79 a_n3792_7061.n52 GND 0.006965f
C80 a_n3792_7061.n53 GND 0.006578f
C81 a_n3792_7061.n54 GND 0.006578f
C82 a_n3792_7061.n55 GND 0.006965f
C83 a_n3792_7061.n56 GND 0.015548f
C84 a_n3792_7061.n57 GND 0.037289f
C85 a_n3792_7061.n58 GND 0.006965f
C86 a_n3792_7061.n59 GND 0.006578f
C87 a_n3792_7061.n60 GND 0.031364f
C88 a_n3792_7061.t9 GND 0.051366f
C89 a_n3792_7061.t10 GND 0.051366f
C90 a_n3792_7061.n61 GND 0.289994f
C91 a_n3792_7061.n62 GND 1.4351f
C92 a_n3792_7061.n63 GND 1.40144f
C93 a_n3792_7061.n64 GND 0.013348f
C94 a_n3792_7061.n65 GND 0.006578f
C95 a_n3792_7061.n66 GND 0.015548f
C96 a_n3792_7061.n67 GND 0.006965f
C97 a_n3792_7061.n68 GND 0.006578f
C98 a_n3792_7061.t7 GND 0.033882f
C99 a_n3792_7061.n69 GND 0.006965f
C100 a_n3792_7061.n70 GND 0.015548f
C101 a_n3792_7061.n71 GND 0.015548f
C102 a_n3792_7061.n72 GND 0.006965f
C103 a_n3792_7061.n73 GND 0.006578f
C104 a_n3792_7061.n74 GND 0.006578f
C105 a_n3792_7061.n75 GND 0.006965f
C106 a_n3792_7061.n76 GND 0.015548f
C107 a_n3792_7061.n77 GND 0.037289f
C108 a_n3792_7061.n78 GND 0.006965f
C109 a_n3792_7061.n79 GND 0.006578f
C110 a_n3792_7061.n80 GND 0.018752f
C111 a_n3792_7061.n81 GND 0.313997f
C112 a_n3792_7061.t4 GND 0.051366f
C113 a_n3792_7061.t2 GND 0.051366f
C114 a_n3792_7061.n82 GND 0.289994f
C115 a_n3792_7061.n83 GND 0.465576f
C116 a_n3792_7061.n84 GND 0.013348f
C117 a_n3792_7061.n85 GND 0.006578f
C118 a_n3792_7061.n86 GND 0.015548f
C119 a_n3792_7061.n87 GND 0.006965f
C120 a_n3792_7061.n88 GND 0.006578f
C121 a_n3792_7061.t1 GND 0.033882f
C122 a_n3792_7061.n89 GND 0.006965f
C123 a_n3792_7061.n90 GND 0.015548f
C124 a_n3792_7061.n91 GND 0.015548f
C125 a_n3792_7061.n92 GND 0.006965f
C126 a_n3792_7061.n93 GND 0.006578f
C127 a_n3792_7061.n94 GND 0.006578f
C128 a_n3792_7061.n95 GND 0.006965f
C129 a_n3792_7061.n96 GND 0.015548f
C130 a_n3792_7061.n97 GND 0.037289f
C131 a_n3792_7061.n98 GND 0.006965f
C132 a_n3792_7061.n99 GND 0.006578f
C133 a_n3792_7061.n100 GND 0.018752f
C134 a_n3792_7061.n101 GND 0.169195f
C135 a_n3792_7061.n102 GND 0.013348f
C136 a_n3792_7061.n103 GND 0.006578f
C137 a_n3792_7061.n104 GND 0.015548f
C138 a_n3792_7061.n105 GND 0.006965f
C139 a_n3792_7061.n106 GND 0.006578f
C140 a_n3792_7061.t5 GND 0.033882f
C141 a_n3792_7061.n107 GND 0.006965f
C142 a_n3792_7061.n108 GND 0.015548f
C143 a_n3792_7061.n109 GND 0.015548f
C144 a_n3792_7061.n110 GND 0.006965f
C145 a_n3792_7061.n111 GND 0.006578f
C146 a_n3792_7061.n112 GND 0.006578f
C147 a_n3792_7061.n113 GND 0.006965f
C148 a_n3792_7061.n114 GND 0.015548f
C149 a_n3792_7061.n115 GND 0.037289f
C150 a_n3792_7061.n116 GND 0.006965f
C151 a_n3792_7061.n117 GND 0.006578f
C152 a_n3792_7061.n118 GND 0.018752f
C153 a_n3792_7061.n119 GND 0.169195f
C154 a_n3792_7061.n120 GND 0.013348f
C155 a_n3792_7061.n121 GND 0.006578f
C156 a_n3792_7061.n122 GND 0.015548f
C157 a_n3792_7061.n123 GND 0.006965f
C158 a_n3792_7061.n124 GND 0.006578f
C159 a_n3792_7061.t6 GND 0.033882f
C160 a_n3792_7061.n125 GND 0.006965f
C161 a_n3792_7061.n126 GND 0.015548f
C162 a_n3792_7061.n127 GND 0.015548f
C163 a_n3792_7061.n128 GND 0.006965f
C164 a_n3792_7061.n129 GND 0.006578f
C165 a_n3792_7061.n130 GND 0.006578f
C166 a_n3792_7061.n131 GND 0.006965f
C167 a_n3792_7061.n132 GND 0.015548f
C168 a_n3792_7061.n133 GND 0.037289f
C169 a_n3792_7061.n134 GND 0.006965f
C170 a_n3792_7061.n135 GND 0.006578f
C171 a_n3792_7061.n136 GND 0.031364f
C172 a_n3792_7061.n137 GND 0.594786f
C173 a_n3792_7061.t3 GND 0.051366f
C174 a_n3792_7061.n138 GND 0.289994f
C175 a_n3792_7061.t8 GND 0.051366f
C176 VP.n0 GND 0.036172f
C177 VP.t7 GND 0.916063f
C178 VP.n1 GND 0.03584f
C179 VP.n2 GND 0.01923f
C180 VP.n3 GND 0.038678f
C181 VP.n4 GND 0.01923f
C182 VP.t4 GND 0.916063f
C183 VP.n5 GND 0.35119f
C184 VP.n6 GND 0.01923f
C185 VP.n7 GND 0.03584f
C186 VP.n8 GND 0.01923f
C187 VP.n9 GND 0.03584f
C188 VP.n10 GND 0.01923f
C189 VP.t6 GND 0.916063f
C190 VP.n11 GND 0.418472f
C191 VP.t3 GND 1.23294f
C192 VP.n12 GND 0.464278f
C193 VP.n13 GND 0.272901f
C194 VP.n14 GND 0.018675f
C195 VP.n15 GND 0.03584f
C196 VP.n16 GND 0.03584f
C197 VP.n17 GND 0.01923f
C198 VP.n18 GND 0.01923f
C199 VP.n19 GND 0.01923f
C200 VP.n20 GND 0.038219f
C201 VP.n21 GND 0.015546f
C202 VP.n22 GND 0.038219f
C203 VP.n23 GND 0.01923f
C204 VP.n24 GND 0.01923f
C205 VP.n25 GND 0.01923f
C206 VP.n26 GND 0.03584f
C207 VP.n27 GND 0.03584f
C208 VP.n28 GND 0.018675f
C209 VP.n29 GND 0.01923f
C210 VP.n30 GND 0.01923f
C211 VP.n31 GND 0.035308f
C212 VP.n32 GND 0.03584f
C213 VP.n33 GND 0.03584f
C214 VP.n34 GND 0.01923f
C215 VP.n35 GND 0.01923f
C216 VP.n36 GND 0.01923f
C217 VP.n37 GND 0.015769f
C218 VP.n38 GND 0.037537f
C219 VP.n39 GND 0.03584f
C220 VP.n40 GND 0.01923f
C221 VP.n41 GND 0.01923f
C222 VP.n42 GND 0.01923f
C223 VP.n43 GND 0.03584f
C224 VP.n44 GND 0.019737f
C225 VP.n45 GND 0.425807f
C226 VP.n46 GND 0.367208f
C227 VP.n47 GND 0.036172f
C228 VP.t2 GND 0.916063f
C229 VP.n48 GND 0.03584f
C230 VP.n49 GND 0.01923f
C231 VP.n50 GND 0.038678f
C232 VP.n51 GND 0.01923f
C233 VP.t5 GND 0.916063f
C234 VP.n52 GND 0.35119f
C235 VP.n53 GND 0.01923f
C236 VP.n54 GND 0.03584f
C237 VP.n55 GND 0.01923f
C238 VP.n56 GND 0.03584f
C239 VP.n57 GND 0.01923f
C240 VP.t9 GND 0.916063f
C241 VP.n58 GND 0.418472f
C242 VP.t8 GND 1.23294f
C243 VP.n59 GND 0.46428f
C244 VP.n60 GND 0.272902f
C245 VP.n61 GND 0.018675f
C246 VP.n62 GND 0.03584f
C247 VP.n63 GND 0.03584f
C248 VP.n64 GND 0.01923f
C249 VP.n65 GND 0.01923f
C250 VP.n66 GND 0.01923f
C251 VP.n67 GND 0.038219f
C252 VP.n68 GND 0.015546f
C253 VP.n69 GND 0.038219f
C254 VP.n70 GND 0.01923f
C255 VP.n71 GND 0.01923f
C256 VP.n72 GND 0.01923f
C257 VP.n73 GND 0.03584f
C258 VP.n74 GND 0.03584f
C259 VP.n75 GND 0.018675f
C260 VP.n76 GND 0.01923f
C261 VP.n77 GND 0.01923f
C262 VP.n78 GND 0.035308f
C263 VP.n79 GND 0.03584f
C264 VP.n80 GND 0.03584f
C265 VP.n81 GND 0.01923f
C266 VP.n82 GND 0.01923f
C267 VP.n83 GND 0.01923f
C268 VP.n84 GND 0.015769f
C269 VP.n85 GND 0.037537f
C270 VP.n86 GND 0.03584f
C271 VP.n87 GND 0.01923f
C272 VP.n88 GND 0.01923f
C273 VP.n89 GND 0.01923f
C274 VP.n90 GND 0.03584f
C275 VP.n91 GND 0.019737f
C276 VP.n92 GND 0.425807f
C277 VP.n93 GND 1.02051f
C278 VP.n94 GND 1.24497f
C279 VP.t1 GND 0.033196f
C280 VP.t0 GND 0.032995f
C281 VP.n95 GND 0.158124f
C282 VP.n96 GND 2.09918f
C283 a_n6793_8883.n0 GND 0.851849f
C284 a_n6793_8883.n1 GND 0.851849f
C285 a_n6793_8883.n2 GND 0.851849f
C286 a_n6793_8883.n3 GND 0.851849f
C287 a_n6793_8883.n4 GND 0.851849f
C288 a_n6793_8883.n5 GND 0.851849f
C289 a_n6793_8883.n6 GND 0.031058f
C290 a_n6793_8883.n7 GND 0.043824f
C291 a_n6793_8883.n8 GND 0.137161f
C292 a_n6793_8883.n9 GND 0.031058f
C293 a_n6793_8883.n10 GND 0.043824f
C294 a_n6793_8883.n11 GND 0.137161f
C295 a_n6793_8883.n12 GND 0.031058f
C296 a_n6793_8883.n13 GND 0.043824f
C297 a_n6793_8883.n14 GND 0.137161f
C298 a_n6793_8883.n15 GND 0.031058f
C299 a_n6793_8883.n16 GND 0.043824f
C300 a_n6793_8883.n17 GND 0.137161f
C301 a_n6793_8883.n18 GND 0.031058f
C302 a_n6793_8883.n19 GND 0.043824f
C303 a_n6793_8883.n20 GND 0.137161f
C304 a_n6793_8883.n21 GND 0.031058f
C305 a_n6793_8883.n22 GND 0.043824f
C306 a_n6793_8883.n23 GND 0.137161f
C307 a_n6793_8883.n24 GND 0.03555f
C308 a_n6793_8883.n25 GND 0.01752f
C309 a_n6793_8883.n26 GND 0.041411f
C310 a_n6793_8883.n27 GND 0.018551f
C311 a_n6793_8883.n28 GND 0.01752f
C312 a_n6793_8883.t4 GND 0.090242f
C313 a_n6793_8883.n29 GND 0.018551f
C314 a_n6793_8883.n30 GND 0.041411f
C315 a_n6793_8883.n31 GND 0.041411f
C316 a_n6793_8883.n32 GND 0.018551f
C317 a_n6793_8883.n33 GND 0.01752f
C318 a_n6793_8883.n34 GND 0.01752f
C319 a_n6793_8883.n35 GND 0.018551f
C320 a_n6793_8883.n36 GND 0.041411f
C321 a_n6793_8883.n37 GND 0.099316f
C322 a_n6793_8883.n38 GND 0.018551f
C323 a_n6793_8883.n39 GND 0.01752f
C324 a_n6793_8883.n40 GND 0.083536f
C325 a_n6793_8883.t0 GND 0.136811f
C326 a_n6793_8883.t2 GND 0.136811f
C327 a_n6793_8883.n41 GND 0.772387f
C328 a_n6793_8883.n42 GND 1.58419f
C329 a_n6793_8883.n43 GND 0.03555f
C330 a_n6793_8883.n44 GND 0.01752f
C331 a_n6793_8883.n45 GND 0.041411f
C332 a_n6793_8883.n46 GND 0.018551f
C333 a_n6793_8883.n47 GND 0.01752f
C334 a_n6793_8883.t3 GND 0.090242f
C335 a_n6793_8883.n48 GND 0.018551f
C336 a_n6793_8883.n49 GND 0.041411f
C337 a_n6793_8883.n50 GND 0.041411f
C338 a_n6793_8883.n51 GND 0.018551f
C339 a_n6793_8883.n52 GND 0.01752f
C340 a_n6793_8883.n53 GND 0.01752f
C341 a_n6793_8883.n54 GND 0.018551f
C342 a_n6793_8883.n55 GND 0.041411f
C343 a_n6793_8883.n56 GND 0.099316f
C344 a_n6793_8883.n57 GND 0.018551f
C345 a_n6793_8883.n58 GND 0.01752f
C346 a_n6793_8883.n59 GND 0.049945f
C347 a_n6793_8883.n60 GND 0.450643f
C348 a_n6793_8883.n61 GND 0.03555f
C349 a_n6793_8883.n62 GND 0.01752f
C350 a_n6793_8883.n63 GND 0.041411f
C351 a_n6793_8883.n64 GND 0.018551f
C352 a_n6793_8883.n65 GND 0.01752f
C353 a_n6793_8883.t6 GND 0.090242f
C354 a_n6793_8883.n66 GND 0.018551f
C355 a_n6793_8883.n67 GND 0.041411f
C356 a_n6793_8883.n68 GND 0.041411f
C357 a_n6793_8883.n69 GND 0.018551f
C358 a_n6793_8883.n70 GND 0.01752f
C359 a_n6793_8883.n71 GND 0.01752f
C360 a_n6793_8883.n72 GND 0.018551f
C361 a_n6793_8883.n73 GND 0.041411f
C362 a_n6793_8883.n74 GND 0.099316f
C363 a_n6793_8883.n75 GND 0.018551f
C364 a_n6793_8883.n76 GND 0.01752f
C365 a_n6793_8883.n77 GND 0.049945f
C366 a_n6793_8883.n78 GND 0.450643f
C367 a_n6793_8883.n79 GND 0.03555f
C368 a_n6793_8883.n80 GND 0.01752f
C369 a_n6793_8883.n81 GND 0.041411f
C370 a_n6793_8883.n82 GND 0.018551f
C371 a_n6793_8883.n83 GND 0.01752f
C372 a_n6793_8883.t13 GND 0.090242f
C373 a_n6793_8883.n84 GND 0.018551f
C374 a_n6793_8883.n85 GND 0.041411f
C375 a_n6793_8883.n86 GND 0.041411f
C376 a_n6793_8883.n87 GND 0.018551f
C377 a_n6793_8883.n88 GND 0.01752f
C378 a_n6793_8883.n89 GND 0.01752f
C379 a_n6793_8883.n90 GND 0.018551f
C380 a_n6793_8883.n91 GND 0.041411f
C381 a_n6793_8883.n92 GND 0.099316f
C382 a_n6793_8883.n93 GND 0.018551f
C383 a_n6793_8883.n94 GND 0.01752f
C384 a_n6793_8883.n95 GND 0.09672f
C385 a_n6793_8883.t9 GND 0.136811f
C386 a_n6793_8883.t8 GND 0.136811f
C387 a_n6793_8883.n96 GND 0.875636f
C388 a_n6793_8883.n97 GND 2.93112f
C389 a_n6793_8883.n98 GND 0.03555f
C390 a_n6793_8883.n99 GND 0.01752f
C391 a_n6793_8883.n100 GND 0.041411f
C392 a_n6793_8883.n101 GND 0.018551f
C393 a_n6793_8883.n102 GND 0.01752f
C394 a_n6793_8883.t12 GND 0.090242f
C395 a_n6793_8883.n103 GND 0.018551f
C396 a_n6793_8883.n104 GND 0.041411f
C397 a_n6793_8883.n105 GND 0.041411f
C398 a_n6793_8883.n106 GND 0.018551f
C399 a_n6793_8883.n107 GND 0.01752f
C400 a_n6793_8883.n108 GND 0.01752f
C401 a_n6793_8883.n109 GND 0.018551f
C402 a_n6793_8883.n110 GND 0.041411f
C403 a_n6793_8883.n111 GND 0.099316f
C404 a_n6793_8883.n112 GND 0.018551f
C405 a_n6793_8883.n113 GND 0.01752f
C406 a_n6793_8883.n114 GND 0.095638f
C407 a_n6793_8883.t11 GND 0.136811f
C408 a_n6793_8883.t10 GND 0.136811f
C409 a_n6793_8883.n115 GND 0.875641f
C410 a_n6793_8883.n116 GND 6.24398f
C411 a_n6793_8883.n117 GND 4.1368f
C412 a_n6793_8883.n118 GND 0.03555f
C413 a_n6793_8883.n119 GND 0.01752f
C414 a_n6793_8883.n120 GND 0.041411f
C415 a_n6793_8883.n121 GND 0.018551f
C416 a_n6793_8883.n122 GND 0.01752f
C417 a_n6793_8883.t5 GND 0.090242f
C418 a_n6793_8883.n123 GND 0.018551f
C419 a_n6793_8883.n124 GND 0.041411f
C420 a_n6793_8883.n125 GND 0.041411f
C421 a_n6793_8883.n126 GND 0.018551f
C422 a_n6793_8883.n127 GND 0.01752f
C423 a_n6793_8883.n128 GND 0.01752f
C424 a_n6793_8883.n129 GND 0.018551f
C425 a_n6793_8883.n130 GND 0.041411f
C426 a_n6793_8883.n131 GND 0.099316f
C427 a_n6793_8883.n132 GND 0.018551f
C428 a_n6793_8883.n133 GND 0.01752f
C429 a_n6793_8883.n134 GND 0.049945f
C430 a_n6793_8883.n135 GND 0.836318f
C431 a_n6793_8883.n136 GND 1.24004f
C432 a_n6793_8883.t1 GND 0.136811f
C433 a_n6793_8883.n137 GND 0.772387f
C434 a_n6793_8883.t7 GND 0.136811f
C435 a_n6715_8686.n0 GND 7.56642f
C436 a_n6715_8686.n1 GND 0.696739f
C437 a_n6715_8686.n2 GND 0.696739f
C438 a_n6715_8686.n3 GND 0.696739f
C439 a_n6715_8686.n4 GND 4.39005f
C440 a_n6715_8686.n5 GND 1.15377f
C441 a_n6715_8686.n6 GND 0.463734f
C442 a_n6715_8686.n7 GND 0.016399f
C443 a_n6715_8686.n8 GND 0.463734f
C444 a_n6715_8686.n9 GND 0.016399f
C445 a_n6715_8686.n10 GND 0.204955f
C446 a_n6715_8686.n11 GND 0.686626f
C447 a_n6715_8686.n12 GND 0.686626f
C448 a_n6715_8686.n13 GND 0.015664f
C449 a_n6715_8686.n15 GND 0.015664f
C450 a_n6715_8686.n17 GND 1.90276f
C451 a_n6715_8686.n18 GND 1.87855f
C452 a_n6715_8686.n19 GND 0.677343f
C453 a_n6715_8686.n20 GND 1.99058f
C454 a_n6715_8686.n21 GND 0.677343f
C455 a_n6715_8686.n22 GND 1.99116f
C456 a_n6715_8686.n23 GND 0.677343f
C457 a_n6715_8686.n24 GND 0.017983f
C458 a_n6715_8686.n25 GND 0.015664f
C459 a_n6715_8686.n26 GND 0.017983f
C460 a_n6715_8686.n27 GND 0.015664f
C461 a_n6715_8686.n28 GND 4.14952f
C462 a_n6715_8686.n29 GND 0.686626f
C463 a_n6715_8686.n30 GND 0.686626f
C464 a_n6715_8686.t13 GND 0.045505f
C465 a_n6715_8686.n31 GND 0.015664f
C466 a_n6715_8686.n32 GND 0.015664f
C467 a_n6715_8686.n33 GND 0.689236f
C468 a_n6715_8686.n34 GND 0.689236f
C469 a_n6715_8686.n35 GND 0.689236f
C470 a_n6715_8686.n36 GND 0.686627f
C471 a_n6715_8686.n37 GND 1.6682f
C472 a_n6715_8686.n38 GND 0.015438f
C473 a_n6715_8686.t10 GND 2.12744f
C474 a_n6715_8686.t8 GND 2.09016f
C475 a_n6715_8686.t0 GND 0.401772f
C476 a_n6715_8686.t17 GND 0.044194f
C477 a_n6715_8686.t1 GND 0.401772f
C478 a_n6715_8686.t18 GND 0.044194f
C479 a_n6715_8686.n39 GND 2.25462f
C480 a_n6715_8686.t2 GND 0.390622f
C481 a_n6715_8686.t19 GND 0.044194f
C482 a_n6715_8686.t16 GND 0.401874f
C483 a_n6715_8686.t3 GND 0.044194f
C484 a_n6715_8686.t40 GND 2.11555f
C485 a_n6715_8686.t37 GND 1.7109f
C486 a_n6715_8686.n40 GND 0.894132f
C487 a_n6715_8686.t27 GND 2.12744f
C488 a_n6715_8686.t15 GND 0.41543f
C489 a_n6715_8686.t7 GND 0.05941f
C490 a_n6715_8686.n41 GND 0.015438f
C491 a_n6715_8686.n42 GND 0.027171f
C492 a_n6715_8686.n43 GND 0.017983f
C493 a_n6715_8686.n44 GND 0.043128f
C494 a_n6715_8686.n45 GND 0.008056f
C495 a_n6715_8686.n46 GND 0.007608f
C496 a_n6715_8686.n47 GND 0.021688f
C497 a_n6715_8686.n48 GND 1.28596f
C498 a_n6715_8686.t12 GND 2.12744f
C499 a_n6715_8686.t6 GND 1.7109f
C500 a_n6715_8686.n49 GND 0.894132f
C501 a_n6715_8686.t14 GND 2.11555f
C502 a_n6715_8686.t31 GND 2.12744f
C503 a_n6715_8686.t21 GND 1.7109f
C504 a_n6715_8686.n50 GND 0.894132f
C505 a_n6715_8686.t22 GND 2.11555f
C506 a_n6715_8686.t29 GND 2.12438f
C507 a_n6715_8686.t39 GND 2.09506f
C508 a_n6715_8686.t23 GND 2.12438f
C509 a_n6715_8686.t35 GND 2.12438f
C510 a_n6715_8686.t38 GND 2.09506f
C511 a_n6715_8686.t30 GND 2.12438f
C512 a_n6715_8686.t26 GND 2.12438f
C513 a_n6715_8686.t33 GND 2.09506f
C514 a_n6715_8686.t28 GND 2.12438f
C515 a_n6715_8686.t36 GND 2.12438f
C516 a_n6715_8686.t34 GND 1.7109f
C517 a_n6715_8686.n51 GND 0.883241f
C518 a_n6715_8686.t25 GND 2.12438f
C519 a_n6715_8686.t32 GND 1.7109f
C520 a_n6715_8686.n52 GND 0.883241f
C521 a_n6715_8686.t24 GND 1.7109f
C522 a_n6715_8686.n53 GND 0.89054f
C523 a_n6715_8686.t41 GND 1.7109f
C524 a_n6715_8686.n54 GND 0.89054f
C525 a_n6715_8686.t20 GND 1.7109f
C526 a_n6715_8686.n55 GND 0.89054f
C527 a_n6715_8686.t4 GND 2.16588f
C528 a_n6715_8686.t11 GND 0.394816f
C529 a_n6715_8686.t9 GND 0.05941f
C530 a_n6715_8686.n56 GND 1.16014f
C531 a_n6715_8686.n57 GND 0.036275f
C532 a_n6715_8686.n58 GND 0.007608f
C533 a_n6715_8686.n59 GND 0.008056f
C534 a_n6715_8686.n60 GND 0.043128f
C535 a_n6715_8686.n61 GND 0.017983f
C536 a_n6715_8686.n62 GND 0.027171f
C537 a_n6715_8686.t5 GND 0.045505f
C538 VDD.t11 GND 0.01213f
C539 VDD.t86 GND 0.01213f
C540 VDD.n0 GND 0.080985f
C541 VDD.t106 GND 0.01213f
C542 VDD.t20 GND 0.01213f
C543 VDD.n1 GND 0.077636f
C544 VDD.n2 GND 0.214882f
C545 VDD.t113 GND 0.01213f
C546 VDD.t24 GND 0.01213f
C547 VDD.n3 GND 0.077636f
C548 VDD.n4 GND 0.112348f
C549 VDD.t3 GND 0.01213f
C550 VDD.t7 GND 0.01213f
C551 VDD.n5 GND 0.077636f
C552 VDD.n6 GND 0.098092f
C553 VDD.t9 GND 0.01213f
C554 VDD.t22 GND 0.01213f
C555 VDD.n7 GND 0.080985f
C556 VDD.t18 GND 0.01213f
C557 VDD.t13 GND 0.01213f
C558 VDD.n8 GND 0.077636f
C559 VDD.n9 GND 0.214882f
C560 VDD.t16 GND 0.01213f
C561 VDD.t83 GND 0.01213f
C562 VDD.n10 GND 0.077636f
C563 VDD.n11 GND 0.112348f
C564 VDD.t108 GND 0.01213f
C565 VDD.t111 GND 0.01213f
C566 VDD.n12 GND 0.077636f
C567 VDD.n13 GND 0.098092f
C568 VDD.n14 GND 0.067041f
C569 VDD.n15 GND 1.8029f
C570 VDD.t88 GND 0.008041f
C571 VDD.t95 GND 0.008041f
C572 VDD.n16 GND 0.042761f
C573 VDD.t97 GND 0.056434f
C574 VDD.n17 GND 0.20908f
C575 VDD.t89 GND 0.008041f
C576 VDD.t103 GND 0.008041f
C577 VDD.n18 GND 0.042761f
C578 VDD.t102 GND 0.056434f
C579 VDD.n19 GND 0.200046f
C580 VDD.n20 GND 0.135807f
C581 VDD.n21 GND 0.004363f
C582 VDD.n22 GND 0.005676f
C583 VDD.n23 GND 0.004569f
C584 VDD.n24 GND 0.004569f
C585 VDD.n25 GND 0.005676f
C586 VDD.n26 GND 0.005676f
C587 VDD.t94 GND 0.19327f
C588 VDD.n27 GND 0.005676f
C589 VDD.n28 GND 0.005676f
C590 VDD.n29 GND 0.005676f
C591 VDD.n30 GND 0.386541f
C592 VDD.n31 GND 0.005676f
C593 VDD.n32 GND 0.005676f
C594 VDD.n33 GND 0.005676f
C595 VDD.n34 GND 0.005676f
C596 VDD.n35 GND 0.004569f
C597 VDD.n36 GND 0.005676f
C598 VDD.n37 GND 0.005676f
C599 VDD.n38 GND 0.005676f
C600 VDD.n39 GND 0.005676f
C601 VDD.n40 GND 0.386541f
C602 VDD.n41 GND 0.005676f
C603 VDD.n42 GND 0.005676f
C604 VDD.n43 GND 0.005676f
C605 VDD.n44 GND 0.005676f
C606 VDD.n45 GND 0.005676f
C607 VDD.n46 GND 0.004569f
C608 VDD.n47 GND 0.005676f
C609 VDD.n48 GND 0.005676f
C610 VDD.n49 GND 0.005676f
C611 VDD.n50 GND 0.005676f
C612 VDD.n51 GND 0.386541f
C613 VDD.n52 GND 0.005676f
C614 VDD.n53 GND 0.005676f
C615 VDD.n54 GND 0.005676f
C616 VDD.n55 GND 0.005676f
C617 VDD.n56 GND 0.005676f
C618 VDD.n57 GND 0.004569f
C619 VDD.n58 GND 0.005676f
C620 VDD.n59 GND 0.005676f
C621 VDD.n60 GND 0.005676f
C622 VDD.n61 GND 0.005676f
C623 VDD.n62 GND 0.386541f
C624 VDD.n63 GND 0.005676f
C625 VDD.n64 GND 0.005676f
C626 VDD.n65 GND 0.005676f
C627 VDD.n66 GND 0.005676f
C628 VDD.n67 GND 0.005676f
C629 VDD.n68 GND 0.004569f
C630 VDD.n69 GND 0.005676f
C631 VDD.n70 GND 0.005676f
C632 VDD.n71 GND 0.005676f
C633 VDD.n72 GND 0.005676f
C634 VDD.n73 GND 0.239655f
C635 VDD.n74 GND 0.005676f
C636 VDD.n75 GND 0.005676f
C637 VDD.n76 GND 0.005676f
C638 VDD.n77 GND 0.005676f
C639 VDD.n78 GND 0.005676f
C640 VDD.n79 GND 0.004569f
C641 VDD.n80 GND 0.005676f
C642 VDD.t31 GND 0.19327f
C643 VDD.n81 GND 0.005676f
C644 VDD.n82 GND 0.005676f
C645 VDD.n83 GND 0.005676f
C646 VDD.n84 GND 0.386541f
C647 VDD.n85 GND 0.005676f
C648 VDD.n86 GND 0.005676f
C649 VDD.n87 GND 0.005676f
C650 VDD.n88 GND 0.005676f
C651 VDD.n89 GND 0.0128f
C652 VDD.n90 GND 0.0128f
C653 VDD.n91 GND 0.0128f
C654 VDD.n102 GND 0.005676f
C655 VDD.t33 GND 0.049112f
C656 VDD.t32 GND 0.063006f
C657 VDD.t30 GND 0.385677f
C658 VDD.n103 GND 0.054096f
C659 VDD.n104 GND 0.037762f
C660 VDD.n105 GND 0.007036f
C661 VDD.n106 GND 0.005676f
C662 VDD.n107 GND 0.004569f
C663 VDD.n108 GND 0.005676f
C664 VDD.n109 GND 0.004569f
C665 VDD.n110 GND 0.005676f
C666 VDD.t43 GND 0.049112f
C667 VDD.t42 GND 0.063006f
C668 VDD.t41 GND 0.385677f
C669 VDD.n111 GND 0.054096f
C670 VDD.n112 GND 0.037762f
C671 VDD.n113 GND 0.00932f
C672 VDD.n114 GND 0.005676f
C673 VDD.n115 GND 0.004569f
C674 VDD.n116 GND 0.005676f
C675 VDD.n117 GND 0.004569f
C676 VDD.n118 GND 0.003792f
C677 VDD.n119 GND 0.0128f
C678 VDD.n120 GND 0.005676f
C679 VDD.n121 GND 0.005676f
C680 VDD.n122 GND 0.005676f
C681 VDD.n123 GND 0.005676f
C682 VDD.n124 GND 0.004569f
C683 VDD.n125 GND 0.004569f
C684 VDD.n126 GND 0.005676f
C685 VDD.n127 GND 0.005676f
C686 VDD.n128 GND 0.004569f
C687 VDD.n129 GND 0.005676f
C688 VDD.n130 GND 0.005676f
C689 VDD.n131 GND 0.005676f
C690 VDD.n132 GND 0.005676f
C691 VDD.n133 GND 0.005676f
C692 VDD.n134 GND 0.004569f
C693 VDD.n135 GND 0.004569f
C694 VDD.n136 GND 0.005676f
C695 VDD.n137 GND 0.005676f
C696 VDD.n138 GND 0.003472f
C697 VDD.n139 GND 0.005676f
C698 VDD.n140 GND 0.005676f
C699 VDD.n141 GND 0.005676f
C700 VDD.n142 GND 0.005676f
C701 VDD.n143 GND 0.005676f
C702 VDD.n144 GND 0.004158f
C703 VDD.n145 GND 0.004569f
C704 VDD.n146 GND 0.005676f
C705 VDD.n147 GND 0.005676f
C706 VDD.n148 GND 0.004569f
C707 VDD.n149 GND 0.005676f
C708 VDD.n150 GND 0.005676f
C709 VDD.n151 GND 0.005676f
C710 VDD.n152 GND 0.005676f
C711 VDD.n153 GND 0.005676f
C712 VDD.n154 GND 0.004569f
C713 VDD.n155 GND 0.004569f
C714 VDD.n156 GND 0.005676f
C715 VDD.n157 GND 0.005676f
C716 VDD.n158 GND 0.004569f
C717 VDD.n159 GND 0.005676f
C718 VDD.n160 GND 0.005676f
C719 VDD.n161 GND 0.005676f
C720 VDD.n162 GND 0.005676f
C721 VDD.n163 GND 0.005676f
C722 VDD.n164 GND 0.004569f
C723 VDD.n165 GND 0.005676f
C724 VDD.n166 GND 0.004569f
C725 VDD.n167 GND 0.002467f
C726 VDD.n168 GND 0.005676f
C727 VDD.n169 GND 0.005676f
C728 VDD.n170 GND 0.004569f
C729 VDD.n171 GND 0.005676f
C730 VDD.n172 GND 0.004569f
C731 VDD.n173 GND 0.005676f
C732 VDD.n174 GND 0.004569f
C733 VDD.n175 GND 0.005676f
C734 VDD.n176 GND 0.004569f
C735 VDD.n177 GND 0.005676f
C736 VDD.n178 GND 0.004569f
C737 VDD.n179 GND 0.005676f
C738 VDD.n180 GND 0.004569f
C739 VDD.n181 GND 0.005676f
C740 VDD.n182 GND 0.004569f
C741 VDD.n183 GND 0.005676f
C742 VDD.n184 GND 0.386541f
C743 VDD.n185 GND 0.005676f
C744 VDD.n186 GND 0.004569f
C745 VDD.n187 GND 0.005676f
C746 VDD.n188 GND 0.004569f
C747 VDD.n189 GND 0.005676f
C748 VDD.n190 GND 0.386541f
C749 VDD.n191 GND 0.005676f
C750 VDD.n192 GND 0.005676f
C751 VDD.n193 GND 0.004569f
C752 VDD.n194 GND 0.005676f
C753 VDD.n195 GND 0.004569f
C754 VDD.n196 GND 0.005676f
C755 VDD.n197 GND 0.386541f
C756 VDD.n198 GND 0.005676f
C757 VDD.n199 GND 0.004569f
C758 VDD.n200 GND 0.005676f
C759 VDD.n201 GND 0.004569f
C760 VDD.n202 GND 0.005676f
C761 VDD.n203 GND 0.247386f
C762 VDD.n204 GND 0.005676f
C763 VDD.n205 GND 0.004569f
C764 VDD.n206 GND 0.005676f
C765 VDD.n207 GND 0.004569f
C766 VDD.n208 GND 0.005676f
C767 VDD.n209 GND 0.386541f
C768 VDD.t87 GND 0.19327f
C769 VDD.n210 GND 0.005676f
C770 VDD.n211 GND 0.004569f
C771 VDD.n212 GND 0.005676f
C772 VDD.n213 GND 0.004569f
C773 VDD.n214 GND 0.005676f
C774 VDD.n215 GND 0.386541f
C775 VDD.n216 GND 0.005676f
C776 VDD.n217 GND 0.004569f
C777 VDD.n218 GND 0.005676f
C778 VDD.n219 GND 0.004569f
C779 VDD.n220 GND 0.005676f
C780 VDD.n221 GND 0.386541f
C781 VDD.n222 GND 0.005676f
C782 VDD.n223 GND 0.004569f
C783 VDD.n224 GND 0.005676f
C784 VDD.n225 GND 0.004569f
C785 VDD.n226 GND 0.005676f
C786 VDD.n227 GND 0.386541f
C787 VDD.n228 GND 0.005676f
C788 VDD.n229 GND 0.004569f
C789 VDD.n230 GND 0.005676f
C790 VDD.n231 GND 0.004569f
C791 VDD.n232 GND 0.005676f
C792 VDD.n233 GND 0.386541f
C793 VDD.n234 GND 0.005676f
C794 VDD.n235 GND 0.004569f
C795 VDD.n236 GND 0.005676f
C796 VDD.n237 GND 0.004569f
C797 VDD.n238 GND 0.005676f
C798 VDD.t67 GND 0.19327f
C799 VDD.n239 GND 0.005676f
C800 VDD.n240 GND 0.004569f
C801 VDD.n241 GND 0.005676f
C802 VDD.n242 GND 0.004569f
C803 VDD.n243 GND 0.005676f
C804 VDD.n244 GND 0.386541f
C805 VDD.n245 GND 0.340156f
C806 VDD.n246 GND 0.005676f
C807 VDD.n247 GND 0.004569f
C808 VDD.n248 GND 0.0128f
C809 VDD.n249 GND 0.003792f
C810 VDD.n250 GND 0.0128f
C811 VDD.n251 GND 0.49284f
C812 VDD.n252 GND 0.0128f
C813 VDD.n253 GND 0.003792f
C814 VDD.n254 GND 0.005676f
C815 VDD.t68 GND 0.049112f
C816 VDD.t69 GND 0.063006f
C817 VDD.t66 GND 0.385677f
C818 VDD.n255 GND 0.054096f
C819 VDD.n256 GND 0.037762f
C820 VDD.n257 GND 0.007036f
C821 VDD.n258 GND 0.005676f
C822 VDD.t12 GND 0.249319f
C823 VDD.n280 GND 0.00386f
C824 VDD.n281 GND 0.009102f
C825 VDD.n282 GND 0.002838f
C826 VDD.n283 GND 0.00386f
C827 VDD.n284 GND 0.00386f
C828 VDD.n285 GND 0.262848f
C829 VDD.n286 GND 0.00386f
C830 VDD.n287 GND 0.35755f
C831 VDD.n288 GND 0.00386f
C832 VDD.n289 GND 0.00386f
C833 VDD.n290 GND 0.009102f
C834 VDD.n291 GND 0.00386f
C835 VDD.t72 GND 0.042906f
C836 VDD.t71 GND 0.059398f
C837 VDD.t70 GND 0.475789f
C838 VDD.n292 GND 0.099866f
C839 VDD.n293 GND 0.077301f
C840 VDD.n294 GND 0.005516f
C841 VDD.n295 GND 0.00386f
C842 VDD.n296 GND 0.00386f
C843 VDD.n297 GND 0.262848f
C844 VDD.n298 GND 0.00386f
C845 VDD.n299 GND 0.00386f
C846 VDD.n300 GND 0.00386f
C847 VDD.n301 GND 0.00386f
C848 VDD.n302 GND 0.00386f
C849 VDD.n303 GND 0.19327f
C850 VDD.n304 GND 0.00386f
C851 VDD.n305 GND 0.00386f
C852 VDD.n306 GND 0.00386f
C853 VDD.n307 GND 0.00386f
C854 VDD.n308 GND 0.00386f
C855 VDD.n309 GND 0.00386f
C856 VDD.n310 GND 0.262848f
C857 VDD.n311 GND 0.00386f
C858 VDD.n312 GND 0.00386f
C859 VDD.t53 GND 0.131424f
C860 VDD.n313 GND 0.00386f
C861 VDD.n314 GND 0.00386f
C862 VDD.n315 GND 0.00386f
C863 VDD.t17 GND 0.131424f
C864 VDD.n316 GND 0.00386f
C865 VDD.n317 GND 0.00386f
C866 VDD.n318 GND 0.00386f
C867 VDD.n319 GND 0.00386f
C868 VDD.n320 GND 0.00386f
C869 VDD.n321 GND 0.262848f
C870 VDD.n322 GND 0.00386f
C871 VDD.n323 GND 0.00386f
C872 VDD.n324 GND 0.237723f
C873 VDD.n325 GND 0.00386f
C874 VDD.n326 GND 0.00386f
C875 VDD.n327 GND 0.00386f
C876 VDD.n328 GND 0.262848f
C877 VDD.n329 GND 0.00386f
C878 VDD.n330 GND 0.00386f
C879 VDD.n331 GND 0.00386f
C880 VDD.n332 GND 0.00386f
C881 VDD.n333 GND 0.00386f
C882 VDD.n334 GND 0.262848f
C883 VDD.n335 GND 0.00386f
C884 VDD.n336 GND 0.00386f
C885 VDD.n337 GND 0.00386f
C886 VDD.n338 GND 0.00386f
C887 VDD.n339 GND 0.00386f
C888 VDD.n340 GND 0.262848f
C889 VDD.n341 GND 0.00386f
C890 VDD.n342 GND 0.00386f
C891 VDD.n343 GND 0.00386f
C892 VDD.n344 GND 0.00386f
C893 VDD.n345 GND 0.00386f
C894 VDD.n346 GND 0.208732f
C895 VDD.n347 GND 0.00386f
C896 VDD.n348 GND 0.00386f
C897 VDD.n349 GND 0.00386f
C898 VDD.n350 GND 0.00386f
C899 VDD.n351 GND 0.00386f
C900 VDD.n352 GND 0.262848f
C901 VDD.n353 GND 0.00386f
C902 VDD.n354 GND 0.00386f
C903 VDD.t0 GND 0.131424f
C904 VDD.n355 GND 0.00386f
C905 VDD.n356 GND 0.00386f
C906 VDD.n357 GND 0.00386f
C907 VDD.n358 GND 0.262848f
C908 VDD.n359 GND 0.00386f
C909 VDD.n360 GND 0.00386f
C910 VDD.n361 GND 0.00386f
C911 VDD.n362 GND 0.00386f
C912 VDD.n363 GND 0.00386f
C913 VDD.t82 GND 0.131424f
C914 VDD.n364 GND 0.00386f
C915 VDD.n365 GND 0.00386f
C916 VDD.n366 GND 0.00386f
C917 VDD.n367 GND 0.00386f
C918 VDD.n368 GND 0.00386f
C919 VDD.n369 GND 0.262848f
C920 VDD.n370 GND 0.00386f
C921 VDD.n371 GND 0.00386f
C922 VDD.n372 GND 0.172011f
C923 VDD.n373 GND 0.00386f
C924 VDD.n374 GND 0.00386f
C925 VDD.n375 GND 0.00386f
C926 VDD.n376 GND 0.262848f
C927 VDD.n377 GND 0.00386f
C928 VDD.n378 GND 0.00386f
C929 VDD.n379 GND 0.00386f
C930 VDD.n380 GND 0.00386f
C931 VDD.n381 GND 0.00386f
C932 VDD.t4 GND 0.131424f
C933 VDD.n382 GND 0.00386f
C934 VDD.n383 GND 0.00386f
C935 VDD.n384 GND 0.00386f
C936 VDD.n385 GND 0.00386f
C937 VDD.n386 GND 0.00386f
C938 VDD.n387 GND 0.262848f
C939 VDD.n388 GND 0.00386f
C940 VDD.n389 GND 0.00386f
C941 VDD.n390 GND 0.197136f
C942 VDD.n391 GND 0.00386f
C943 VDD.n392 GND 0.00386f
C944 VDD.n393 GND 0.00386f
C945 VDD.n394 GND 0.210665f
C946 VDD.n395 GND 0.00386f
C947 VDD.n396 GND 0.00386f
C948 VDD.n397 GND 0.00386f
C949 VDD.n398 GND 0.00386f
C950 VDD.n399 GND 0.00386f
C951 VDD.n400 GND 0.262848f
C952 VDD.n401 GND 0.00386f
C953 VDD.n402 GND 0.00386f
C954 VDD.t15 GND 0.131424f
C955 VDD.n403 GND 0.00386f
C956 VDD.n404 GND 0.00386f
C957 VDD.n405 GND 0.00386f
C958 VDD.n406 GND 0.262848f
C959 VDD.n407 GND 0.00386f
C960 VDD.n408 GND 0.00386f
C961 VDD.n409 GND 0.00386f
C962 VDD.n410 GND 0.00386f
C963 VDD.n411 GND 0.00386f
C964 VDD.n412 GND 0.18554f
C965 VDD.n413 GND 0.00386f
C966 VDD.n414 GND 0.00386f
C967 VDD.n415 GND 0.00386f
C968 VDD.n416 GND 0.00386f
C969 VDD.n417 GND 0.00386f
C970 VDD.n418 GND 0.262848f
C971 VDD.n419 GND 0.00386f
C972 VDD.n420 GND 0.00386f
C973 VDD.t5 GND 0.131424f
C974 VDD.n421 GND 0.00386f
C975 VDD.n422 GND 0.00386f
C976 VDD.n423 GND 0.00386f
C977 VDD.n424 GND 0.262848f
C978 VDD.n425 GND 0.00386f
C979 VDD.n426 GND 0.00386f
C980 VDD.n427 GND 0.00386f
C981 VDD.n428 GND 0.00386f
C982 VDD.n429 GND 0.00386f
C983 VDD.t110 GND 0.131424f
C984 VDD.n430 GND 0.00386f
C985 VDD.n431 GND 0.00386f
C986 VDD.n432 GND 0.00386f
C987 VDD.n433 GND 0.00386f
C988 VDD.n434 GND 0.00386f
C989 VDD.n435 GND 0.262848f
C990 VDD.n436 GND 0.00386f
C991 VDD.n437 GND 0.00386f
C992 VDD.n438 GND 0.195203f
C993 VDD.n439 GND 0.00386f
C994 VDD.n440 GND 0.00386f
C995 VDD.n441 GND 0.00386f
C996 VDD.n442 GND 0.262848f
C997 VDD.n443 GND 0.00386f
C998 VDD.n444 GND 0.00386f
C999 VDD.n445 GND 0.00386f
C1000 VDD.n446 GND 0.00386f
C1001 VDD.n447 GND 0.00386f
C1002 VDD.n448 GND 0.262848f
C1003 VDD.n449 GND 0.00386f
C1004 VDD.n450 GND 0.00386f
C1005 VDD.n451 GND 0.00386f
C1006 VDD.n452 GND 0.00386f
C1007 VDD.n453 GND 0.00386f
C1008 VDD.n454 GND 0.201001f
C1009 VDD.n455 GND 0.00386f
C1010 VDD.n456 GND 0.00386f
C1011 VDD.n457 GND 0.00386f
C1012 VDD.n458 GND 0.00386f
C1013 VDD.n459 GND 0.00386f
C1014 VDD.n460 GND 0.187472f
C1015 VDD.n461 GND 0.00386f
C1016 VDD.n462 GND 0.00386f
C1017 VDD.t49 GND 0.131424f
C1018 VDD.n463 GND 0.00386f
C1019 VDD.n464 GND 0.00386f
C1020 VDD.n465 GND 0.00386f
C1021 VDD.n466 GND 0.262848f
C1022 VDD.n467 GND 0.00386f
C1023 VDD.n468 GND 0.00386f
C1024 VDD.t107 GND 0.131424f
C1025 VDD.n469 GND 0.00386f
C1026 VDD.n470 GND 0.00386f
C1027 VDD.n471 GND 0.00386f
C1028 VDD.n472 GND 0.262848f
C1029 VDD.n473 GND 0.00386f
C1030 VDD.n474 GND 0.00386f
C1031 VDD.n475 GND 0.00386f
C1032 VDD.n476 GND 0.009516f
C1033 VDD.n477 GND 0.009516f
C1034 VDD.n478 GND 0.380743f
C1035 VDD.n500 GND 0.00386f
C1036 VDD.n501 GND 0.009102f
C1037 VDD.n502 GND 0.002838f
C1038 VDD.n503 GND 0.00386f
C1039 VDD.n504 GND 0.00386f
C1040 VDD.n505 GND 0.262848f
C1041 VDD.n506 GND 0.00386f
C1042 VDD.n507 GND 0.00386f
C1043 VDD.n508 GND 0.00386f
C1044 VDD.n509 GND 0.009102f
C1045 VDD.n510 GND 0.00386f
C1046 VDD.t58 GND 0.042906f
C1047 VDD.t57 GND 0.059398f
C1048 VDD.t56 GND 0.475789f
C1049 VDD.n511 GND 0.099866f
C1050 VDD.n512 GND 0.077301f
C1051 VDD.n513 GND 0.005516f
C1052 VDD.n514 GND 0.00386f
C1053 VDD.n515 GND 0.00386f
C1054 VDD.n516 GND 0.206799f
C1055 VDD.n517 GND 0.00386f
C1056 VDD.n518 GND 0.00386f
C1057 VDD.n519 GND 0.00386f
C1058 VDD.n520 GND 0.00386f
C1059 VDD.n521 GND 0.00386f
C1060 VDD.n522 GND 0.19327f
C1061 VDD.n523 GND 0.00386f
C1062 VDD.n524 GND 0.00386f
C1063 VDD.t6 GND 0.131424f
C1064 VDD.n525 GND 0.00386f
C1065 VDD.n526 GND 0.00386f
C1066 VDD.n527 GND 0.00386f
C1067 VDD.n528 GND 0.00386f
C1068 VDD.n529 GND 0.262848f
C1069 VDD.n530 GND 0.00386f
C1070 VDD.n531 GND 0.00386f
C1071 VDD.t45 GND 0.131424f
C1072 VDD.n532 GND 0.00386f
C1073 VDD.n533 GND 0.00386f
C1074 VDD.n534 GND 0.00386f
C1075 VDD.n535 GND 0.262848f
C1076 VDD.n536 GND 0.00386f
C1077 VDD.n537 GND 0.00386f
C1078 VDD.n538 GND 0.00386f
C1079 VDD.n539 GND 0.00386f
C1080 VDD.n540 GND 0.00386f
C1081 VDD.n541 GND 0.262848f
C1082 VDD.n542 GND 0.00386f
C1083 VDD.n543 GND 0.00386f
C1084 VDD.n544 GND 0.00386f
C1085 VDD.n545 GND 0.00386f
C1086 VDD.n546 GND 0.00386f
C1087 VDD.n547 GND 0.262848f
C1088 VDD.n548 GND 0.00386f
C1089 VDD.n549 GND 0.00386f
C1090 VDD.n550 GND 0.00386f
C1091 VDD.n551 GND 0.00386f
C1092 VDD.n552 GND 0.00386f
C1093 VDD.t2 GND 0.131424f
C1094 VDD.n553 GND 0.00386f
C1095 VDD.n554 GND 0.00386f
C1096 VDD.n555 GND 0.00386f
C1097 VDD.n556 GND 0.00386f
C1098 VDD.n557 GND 0.00386f
C1099 VDD.n558 GND 0.262848f
C1100 VDD.n559 GND 0.00386f
C1101 VDD.n560 GND 0.00386f
C1102 VDD.n561 GND 0.199069f
C1103 VDD.n562 GND 0.00386f
C1104 VDD.n563 GND 0.00386f
C1105 VDD.n564 GND 0.00386f
C1106 VDD.n565 GND 0.208732f
C1107 VDD.n566 GND 0.00386f
C1108 VDD.n567 GND 0.00386f
C1109 VDD.n568 GND 0.00386f
C1110 VDD.n569 GND 0.00386f
C1111 VDD.n570 GND 0.00386f
C1112 VDD.n571 GND 0.262848f
C1113 VDD.n572 GND 0.00386f
C1114 VDD.n573 GND 0.00386f
C1115 VDD.t14 GND 0.131424f
C1116 VDD.n574 GND 0.00386f
C1117 VDD.n575 GND 0.00386f
C1118 VDD.n576 GND 0.00386f
C1119 VDD.n577 GND 0.262848f
C1120 VDD.n578 GND 0.00386f
C1121 VDD.n579 GND 0.00386f
C1122 VDD.n580 GND 0.00386f
C1123 VDD.n581 GND 0.00386f
C1124 VDD.n582 GND 0.00386f
C1125 VDD.n583 GND 0.183607f
C1126 VDD.n584 GND 0.00386f
C1127 VDD.n585 GND 0.00386f
C1128 VDD.n586 GND 0.00386f
C1129 VDD.n587 GND 0.00386f
C1130 VDD.n588 GND 0.00386f
C1131 VDD.n589 GND 0.262848f
C1132 VDD.n590 GND 0.00386f
C1133 VDD.n591 GND 0.00386f
C1134 VDD.t23 GND 0.131424f
C1135 VDD.n592 GND 0.00386f
C1136 VDD.n593 GND 0.00386f
C1137 VDD.n594 GND 0.00386f
C1138 VDD.n595 GND 0.262848f
C1139 VDD.n596 GND 0.00386f
C1140 VDD.n597 GND 0.00386f
C1141 VDD.n598 GND 0.00386f
C1142 VDD.n599 GND 0.00386f
C1143 VDD.n600 GND 0.00386f
C1144 VDD.t25 GND 0.131424f
C1145 VDD.n601 GND 0.00386f
C1146 VDD.n602 GND 0.00386f
C1147 VDD.n603 GND 0.00386f
C1148 VDD.n604 GND 0.00386f
C1149 VDD.n605 GND 0.00386f
C1150 VDD.n606 GND 0.262848f
C1151 VDD.n607 GND 0.00386f
C1152 VDD.n608 GND 0.00386f
C1153 VDD.n609 GND 0.197136f
C1154 VDD.n610 GND 0.00386f
C1155 VDD.n611 GND 0.00386f
C1156 VDD.n612 GND 0.00386f
C1157 VDD.n613 GND 0.262848f
C1158 VDD.n614 GND 0.00386f
C1159 VDD.n615 GND 0.00386f
C1160 VDD.n616 GND 0.00386f
C1161 VDD.n617 GND 0.00386f
C1162 VDD.n618 GND 0.00386f
C1163 VDD.t112 GND 0.131424f
C1164 VDD.n619 GND 0.00386f
C1165 VDD.n620 GND 0.00386f
C1166 VDD.n621 GND 0.00386f
C1167 VDD.n622 GND 0.00386f
C1168 VDD.n623 GND 0.00386f
C1169 VDD.n624 GND 0.262848f
C1170 VDD.n625 GND 0.00386f
C1171 VDD.n626 GND 0.00386f
C1172 VDD.n627 GND 0.222261f
C1173 VDD.n628 GND 0.00386f
C1174 VDD.n629 GND 0.00386f
C1175 VDD.n630 GND 0.00386f
C1176 VDD.n631 GND 0.18554f
C1177 VDD.n632 GND 0.00386f
C1178 VDD.n633 GND 0.00386f
C1179 VDD.n634 GND 0.00386f
C1180 VDD.n635 GND 0.00386f
C1181 VDD.n636 GND 0.00386f
C1182 VDD.n637 GND 0.262848f
C1183 VDD.n638 GND 0.00386f
C1184 VDD.n639 GND 0.00386f
C1185 VDD.t1 GND 0.131424f
C1186 VDD.n640 GND 0.00386f
C1187 VDD.n641 GND 0.00386f
C1188 VDD.n642 GND 0.00386f
C1189 VDD.n643 GND 0.262848f
C1190 VDD.n644 GND 0.00386f
C1191 VDD.n645 GND 0.00386f
C1192 VDD.n646 GND 0.00386f
C1193 VDD.n647 GND 0.00386f
C1194 VDD.n648 GND 0.00386f
C1195 VDD.n649 GND 0.262848f
C1196 VDD.n650 GND 0.00386f
C1197 VDD.n651 GND 0.00386f
C1198 VDD.n652 GND 0.00386f
C1199 VDD.n653 GND 0.00386f
C1200 VDD.n654 GND 0.00386f
C1201 VDD.n655 GND 0.262848f
C1202 VDD.n656 GND 0.00386f
C1203 VDD.n657 GND 0.00386f
C1204 VDD.n658 GND 0.00386f
C1205 VDD.n659 GND 0.00386f
C1206 VDD.n660 GND 0.00386f
C1207 VDD.n661 GND 0.262848f
C1208 VDD.n662 GND 0.00386f
C1209 VDD.n663 GND 0.00386f
C1210 VDD.n664 GND 0.00386f
C1211 VDD.n665 GND 0.00386f
C1212 VDD.n666 GND 0.00386f
C1213 VDD.t19 GND 0.131424f
C1214 VDD.n667 GND 0.00386f
C1215 VDD.n668 GND 0.00386f
C1216 VDD.n669 GND 0.00386f
C1217 VDD.n670 GND 0.00386f
C1218 VDD.n671 GND 0.00386f
C1219 VDD.n672 GND 0.201001f
C1220 VDD.n673 GND 0.00386f
C1221 VDD.n674 GND 0.00386f
C1222 VDD.n675 GND 0.156549f
C1223 VDD.n676 GND 0.00386f
C1224 VDD.n677 GND 0.00386f
C1225 VDD.n678 GND 0.00386f
C1226 VDD.n679 GND 0.262848f
C1227 VDD.n680 GND 0.00386f
C1228 VDD.n681 GND 0.00386f
C1229 VDD.t35 GND 0.131424f
C1230 VDD.n682 GND 0.00386f
C1231 VDD.n683 GND 0.00386f
C1232 VDD.n684 GND 0.00386f
C1233 VDD.n685 GND 0.262848f
C1234 VDD.n686 GND 0.00386f
C1235 VDD.n687 GND 0.00386f
C1236 VDD.n688 GND 0.00386f
C1237 VDD.n689 GND 0.00386f
C1238 VDD.n690 GND 0.00386f
C1239 VDD.n691 GND 0.262848f
C1240 VDD.n692 GND 0.00386f
C1241 VDD.n693 GND 0.00386f
C1242 VDD.n694 GND 0.00386f
C1243 VDD.n695 GND 0.009516f
C1244 VDD.n696 GND 0.009516f
C1245 VDD.t105 GND 0.249319f
C1246 VDD.n697 GND 0.009102f
C1247 VDD.n698 GND 0.009102f
C1248 VDD.n699 GND 0.009516f
C1249 VDD.n700 GND 0.00386f
C1250 VDD.n701 GND 0.00386f
C1251 VDD.n702 GND 0.49284f
C1252 VDD.n713 GND 0.005676f
C1253 VDD.n714 GND 0.0128f
C1254 VDD.t62 GND 0.049112f
C1255 VDD.t61 GND 0.063006f
C1256 VDD.t59 GND 0.385677f
C1257 VDD.n715 GND 0.054096f
C1258 VDD.n716 GND 0.037762f
C1259 VDD.n717 GND 0.007036f
C1260 VDD.n718 GND 0.005676f
C1261 VDD.n719 GND 0.005676f
C1262 VDD.n720 GND 0.004569f
C1263 VDD.n721 GND 0.005676f
C1264 VDD.n722 GND 0.386541f
C1265 VDD.n723 GND 0.005676f
C1266 VDD.n724 GND 0.0128f
C1267 VDD.n725 GND 0.004569f
C1268 VDD.n726 GND 0.003792f
C1269 VDD.n727 GND 0.005676f
C1270 VDD.n728 GND 0.004569f
C1271 VDD.n729 GND 0.005676f
C1272 VDD.n730 GND 0.340156f
C1273 VDD.n731 GND 0.005676f
C1274 VDD.n732 GND 0.004569f
C1275 VDD.n733 GND 0.005676f
C1276 VDD.n734 GND 0.004569f
C1277 VDD.n735 GND 0.005676f
C1278 VDD.n736 GND 0.386541f
C1279 VDD.t60 GND 0.19327f
C1280 VDD.n737 GND 0.005676f
C1281 VDD.n738 GND 0.004569f
C1282 VDD.n739 GND 0.005676f
C1283 VDD.n740 GND 0.004569f
C1284 VDD.n741 GND 0.005676f
C1285 VDD.n742 GND 0.386541f
C1286 VDD.n743 GND 0.005676f
C1287 VDD.n744 GND 0.004569f
C1288 VDD.n745 GND 0.005676f
C1289 VDD.n746 GND 0.004569f
C1290 VDD.n747 GND 0.005676f
C1291 VDD.n748 GND 0.386541f
C1292 VDD.n749 GND 0.005676f
C1293 VDD.n750 GND 0.004569f
C1294 VDD.n751 GND 0.005676f
C1295 VDD.n752 GND 0.004569f
C1296 VDD.n753 GND 0.005676f
C1297 VDD.n754 GND 0.386541f
C1298 VDD.n755 GND 0.005676f
C1299 VDD.n756 GND 0.004569f
C1300 VDD.n757 GND 0.005676f
C1301 VDD.n758 GND 0.004569f
C1302 VDD.n759 GND 0.005676f
C1303 VDD.n760 GND 0.386541f
C1304 VDD.n761 GND 0.005676f
C1305 VDD.n762 GND 0.004569f
C1306 VDD.n763 GND 0.005676f
C1307 VDD.n764 GND 0.004569f
C1308 VDD.n765 GND 0.005676f
C1309 VDD.t98 GND 0.19327f
C1310 VDD.n766 GND 0.005676f
C1311 VDD.n767 GND 0.004569f
C1312 VDD.n768 GND 0.005676f
C1313 VDD.n769 GND 0.004569f
C1314 VDD.n770 GND 0.005676f
C1315 VDD.n771 GND 0.386541f
C1316 VDD.n772 GND 0.247386f
C1317 VDD.n773 GND 0.005676f
C1318 VDD.n774 GND 0.004569f
C1319 VDD.n775 GND 0.005676f
C1320 VDD.n776 GND 0.004569f
C1321 VDD.n777 GND 0.005676f
C1322 VDD.n778 GND 0.386541f
C1323 VDD.n779 GND 0.005676f
C1324 VDD.n780 GND 0.004569f
C1325 VDD.n781 GND 0.005676f
C1326 VDD.n782 GND 0.004569f
C1327 VDD.n783 GND 0.005676f
C1328 VDD.n784 GND 0.386541f
C1329 VDD.n785 GND 0.005676f
C1330 VDD.n786 GND 0.004569f
C1331 VDD.n787 GND 0.004363f
C1332 VDD.n788 GND 0.004569f
C1333 VDD.n789 GND 0.005676f
C1334 VDD.n790 GND 0.289906f
C1335 VDD.n791 GND 0.005676f
C1336 VDD.n792 GND 0.004569f
C1337 VDD.n793 GND 0.005676f
C1338 VDD.n794 GND 0.004569f
C1339 VDD.n795 GND 0.005676f
C1340 VDD.n796 GND 0.386541f
C1341 VDD.t92 GND 0.19327f
C1342 VDD.n797 GND 0.005676f
C1343 VDD.n798 GND 0.004569f
C1344 VDD.n799 GND 0.005676f
C1345 VDD.n800 GND 0.004569f
C1346 VDD.n801 GND 0.005676f
C1347 VDD.n802 GND 0.386541f
C1348 VDD.n803 GND 0.005676f
C1349 VDD.n804 GND 0.004569f
C1350 VDD.n805 GND 0.005676f
C1351 VDD.n806 GND 0.004569f
C1352 VDD.n807 GND 0.005676f
C1353 VDD.n808 GND 0.386541f
C1354 VDD.n809 GND 0.005676f
C1355 VDD.n810 GND 0.004569f
C1356 VDD.n811 GND 0.005676f
C1357 VDD.n812 GND 0.004569f
C1358 VDD.n813 GND 0.005676f
C1359 VDD.n814 GND 0.386541f
C1360 VDD.n815 GND 0.005676f
C1361 VDD.n816 GND 0.004569f
C1362 VDD.n817 GND 0.005676f
C1363 VDD.n818 GND 0.004569f
C1364 VDD.n819 GND 0.005676f
C1365 VDD.t90 GND 0.19327f
C1366 VDD.n820 GND 0.005676f
C1367 VDD.n821 GND 0.004569f
C1368 VDD.n822 GND 0.005676f
C1369 VDD.n823 GND 0.004569f
C1370 VDD.n824 GND 0.005676f
C1371 VDD.n825 GND 0.386541f
C1372 VDD.n826 GND 0.005676f
C1373 VDD.n827 GND 0.004569f
C1374 VDD.n828 GND 0.005676f
C1375 VDD.n829 GND 0.004569f
C1376 VDD.n830 GND 0.005676f
C1377 VDD.n831 GND 0.386541f
C1378 VDD.n832 GND 0.005676f
C1379 VDD.n833 GND 0.004569f
C1380 VDD.n834 GND 0.005676f
C1381 VDD.n835 GND 0.004569f
C1382 VDD.n836 GND 0.005676f
C1383 VDD.n837 GND 0.386541f
C1384 VDD.n838 GND 0.005676f
C1385 VDD.n839 GND 0.004569f
C1386 VDD.n840 GND 0.005676f
C1387 VDD.n841 GND 0.004569f
C1388 VDD.n842 GND 0.005676f
C1389 VDD.n843 GND 0.386541f
C1390 VDD.n844 GND 0.005676f
C1391 VDD.n845 GND 0.004569f
C1392 VDD.n846 GND 0.005676f
C1393 VDD.n847 GND 0.004569f
C1394 VDD.n848 GND 0.005676f
C1395 VDD.n849 GND 0.239655f
C1396 VDD.n850 GND 0.005676f
C1397 VDD.n851 GND 0.004569f
C1398 VDD.n852 GND 0.005676f
C1399 VDD.n853 GND 0.004569f
C1400 VDD.n854 GND 0.005676f
C1401 VDD.n855 GND 0.386541f
C1402 VDD.t27 GND 0.19327f
C1403 VDD.n856 GND 0.005676f
C1404 VDD.n857 GND 0.004569f
C1405 VDD.n858 GND 0.005676f
C1406 VDD.n859 GND 0.004569f
C1407 VDD.n860 GND 0.005676f
C1408 VDD.n861 GND 0.386541f
C1409 VDD.n862 GND 0.005676f
C1410 VDD.n863 GND 0.004569f
C1411 VDD.n864 GND 0.0128f
C1412 VDD.n865 GND 0.0128f
C1413 VDD.n866 GND 0.836861f
C1414 VDD.n867 GND 0.0128f
C1415 VDD.n868 GND 0.005676f
C1416 VDD.n870 GND 0.005676f
C1417 VDD.n871 GND 0.005676f
C1418 VDD.n872 GND 0.004569f
C1419 VDD.n873 GND 0.005676f
C1420 VDD.n874 GND 0.005676f
C1421 VDD.n876 GND 0.005676f
C1422 VDD.n877 GND 0.005676f
C1423 VDD.n879 GND 0.005676f
C1424 VDD.n880 GND 0.004569f
C1425 VDD.n881 GND 0.005676f
C1426 VDD.n882 GND 0.005676f
C1427 VDD.n884 GND 0.005676f
C1428 VDD.n885 GND 0.004158f
C1429 VDD.n887 GND 0.004569f
C1430 VDD.n888 GND 0.005676f
C1431 VDD.n889 GND 0.005676f
C1432 VDD.n890 GND 0.005676f
C1433 VDD.n891 GND 0.005676f
C1434 VDD.n893 GND 0.005676f
C1435 VDD.n894 GND 0.005676f
C1436 VDD.n895 GND 0.004569f
C1437 VDD.n896 GND 0.005676f
C1438 VDD.n898 GND 0.005676f
C1439 VDD.n899 GND 0.005676f
C1440 VDD.n901 GND 0.005676f
C1441 VDD.n902 GND 0.005676f
C1442 VDD.n904 GND 0.005676f
C1443 VDD.n905 GND 0.002102f
C1444 VDD.t28 GND 0.049112f
C1445 VDD.t29 GND 0.063006f
C1446 VDD.t26 GND 0.385677f
C1447 VDD.n906 GND 0.054096f
C1448 VDD.n907 GND 0.037762f
C1449 VDD.n908 GND 0.007036f
C1450 VDD.n909 GND 0.002467f
C1451 VDD.n910 GND 0.005676f
C1452 VDD.n911 GND 0.005676f
C1453 VDD.n912 GND 0.004569f
C1454 VDD.n913 GND 0.004569f
C1455 VDD.n914 GND 0.004569f
C1456 VDD.n915 GND 0.005676f
C1457 VDD.n916 GND 0.005676f
C1458 VDD.n917 GND 0.005676f
C1459 VDD.n918 GND 0.004569f
C1460 VDD.n919 GND 0.004569f
C1461 VDD.n920 GND 0.004569f
C1462 VDD.n921 GND 0.005676f
C1463 VDD.n922 GND 0.005676f
C1464 VDD.n923 GND 0.005676f
C1465 VDD.n924 GND 0.004569f
C1466 VDD.n925 GND 0.005676f
C1467 VDD.n926 GND 0.005676f
C1468 VDD.n928 GND 0.005676f
C1469 VDD.t39 GND 0.049112f
C1470 VDD.t40 GND 0.063006f
C1471 VDD.t38 GND 0.385677f
C1472 VDD.n929 GND 0.054096f
C1473 VDD.n930 GND 0.037762f
C1474 VDD.n931 GND 0.00932f
C1475 VDD.n932 GND 0.003472f
C1476 VDD.n933 GND 0.005676f
C1477 VDD.n934 GND 0.005676f
C1478 VDD.n935 GND 0.005676f
C1479 VDD.n936 GND 0.004569f
C1480 VDD.n937 GND 0.004569f
C1481 VDD.n938 GND 0.004569f
C1482 VDD.n939 GND 0.005676f
C1483 VDD.n940 GND 0.005676f
C1484 VDD.n941 GND 0.005676f
C1485 VDD.n942 GND 0.004569f
C1486 VDD.n943 GND 0.004569f
C1487 VDD.n944 GND 0.003792f
C1488 VDD.n945 GND 0.0128f
C1489 VDD.n946 GND 0.0128f
C1490 VDD.n947 GND 0.003792f
C1491 VDD.n948 GND 0.0128f
C1492 VDD.n949 GND 0.49284f
C1493 VDD.n950 GND 0.0128f
C1494 VDD.n951 GND 0.003792f
C1495 VDD.n952 GND 0.0128f
C1496 VDD.n953 GND 0.005676f
C1497 VDD.n954 GND 0.005676f
C1498 VDD.n955 GND 0.004569f
C1499 VDD.n956 GND 0.005676f
C1500 VDD.n957 GND 0.386541f
C1501 VDD.n958 GND 0.005676f
C1502 VDD.n959 GND 0.004569f
C1503 VDD.n960 GND 0.005676f
C1504 VDD.n961 GND 0.005676f
C1505 VDD.n962 GND 0.005676f
C1506 VDD.n963 GND 0.004569f
C1507 VDD.n964 GND 0.005676f
C1508 VDD.n965 GND 0.340156f
C1509 VDD.n966 GND 0.005676f
C1510 VDD.n967 GND 0.004569f
C1511 VDD.n968 GND 0.005676f
C1512 VDD.n969 GND 0.005676f
C1513 VDD.n970 GND 0.005676f
C1514 VDD.n971 GND 0.004569f
C1515 VDD.n972 GND 0.005676f
C1516 VDD.n973 GND 0.386541f
C1517 VDD.n974 GND 0.005676f
C1518 VDD.n975 GND 0.004569f
C1519 VDD.n976 GND 0.005676f
C1520 VDD.n977 GND 0.005676f
C1521 VDD.n978 GND 0.005676f
C1522 VDD.n979 GND 0.004569f
C1523 VDD.n980 GND 0.005676f
C1524 VDD.n981 GND 0.386541f
C1525 VDD.n982 GND 0.005676f
C1526 VDD.n983 GND 0.004569f
C1527 VDD.n984 GND 0.005676f
C1528 VDD.n985 GND 0.005676f
C1529 VDD.n986 GND 0.005676f
C1530 VDD.n987 GND 0.004569f
C1531 VDD.n988 GND 0.005676f
C1532 VDD.n989 GND 0.386541f
C1533 VDD.n990 GND 0.005676f
C1534 VDD.n991 GND 0.004569f
C1535 VDD.n992 GND 0.005676f
C1536 VDD.n993 GND 0.005676f
C1537 VDD.n994 GND 0.005676f
C1538 VDD.n995 GND 0.004569f
C1539 VDD.n996 GND 0.005676f
C1540 VDD.n997 GND 0.386541f
C1541 VDD.n998 GND 0.005676f
C1542 VDD.n999 GND 0.004569f
C1543 VDD.n1000 GND 0.005676f
C1544 VDD.n1001 GND 0.005676f
C1545 VDD.n1002 GND 0.005676f
C1546 VDD.n1003 GND 0.004569f
C1547 VDD.n1004 GND 0.005676f
C1548 VDD.n1005 GND 0.332425f
C1549 VDD.n1006 GND 0.386541f
C1550 VDD.n1007 GND 0.005676f
C1551 VDD.n1008 GND 0.004569f
C1552 VDD.n1009 GND 0.005676f
C1553 VDD.n1010 GND 0.005676f
C1554 VDD.n1011 GND 0.005676f
C1555 VDD.n1012 GND 0.004569f
C1556 VDD.n1013 GND 0.005676f
C1557 VDD.n1014 GND 0.247386f
C1558 VDD.n1015 GND 0.005676f
C1559 VDD.n1016 GND 0.004569f
C1560 VDD.n1017 GND 0.005676f
C1561 VDD.n1018 GND 0.005676f
C1562 VDD.n1019 GND 0.005676f
C1563 VDD.n1020 GND 0.004569f
C1564 VDD.n1021 GND 0.005676f
C1565 VDD.n1022 GND 0.386541f
C1566 VDD.n1023 GND 0.005676f
C1567 VDD.n1024 GND 0.004569f
C1568 VDD.n1025 GND 0.005676f
C1569 VDD.n1026 GND 0.005676f
C1570 VDD.n1027 GND 0.005676f
C1571 VDD.n1028 GND 0.004569f
C1572 VDD.n1029 GND 0.005676f
C1573 VDD.n1030 GND 0.386541f
C1574 VDD.n1031 GND 0.005676f
C1575 VDD.n1032 GND 0.004569f
C1576 VDD.n1033 GND 0.005676f
C1577 VDD.n1034 GND 0.005676f
C1578 VDD.n1035 GND 0.005676f
C1579 VDD.n1036 GND 0.004569f
C1580 VDD.n1037 GND 0.005676f
C1581 VDD.n1038 GND 0.386541f
C1582 VDD.n1039 GND 0.005676f
C1583 VDD.n1040 GND 0.004569f
C1584 VDD.n1041 GND 0.005676f
C1585 VDD.n1042 GND 0.005676f
C1586 VDD.t99 GND 0.059081f
C1587 VDD.t91 GND 0.008041f
C1588 VDD.t93 GND 0.008041f
C1589 VDD.n1043 GND 0.038801f
C1590 VDD.n1044 GND 0.202753f
C1591 VDD.t104 GND 0.059081f
C1592 VDD.t100 GND 0.008041f
C1593 VDD.t101 GND 0.008041f
C1594 VDD.n1045 GND 0.038801f
C1595 VDD.n1046 GND 0.1935f
C1596 VDD.n1047 GND 0.151308f
C1597 VDD.n1048 GND 2.21347f
C1598 VDD.n1049 GND 0.545011f
C1599 VDD.n1050 GND 0.004363f
C1600 VDD.n1051 GND 0.004569f
C1601 VDD.n1052 GND 0.005676f
C1602 VDD.n1053 GND 0.289906f
C1603 VDD.n1054 GND 0.005676f
C1604 VDD.n1055 GND 0.004569f
C1605 VDD.n1056 GND 0.005676f
C1606 VDD.n1057 GND 0.005676f
C1607 VDD.n1058 GND 0.005676f
C1608 VDD.n1059 GND 0.004569f
C1609 VDD.n1060 GND 0.005676f
C1610 VDD.n1061 GND 0.386541f
C1611 VDD.n1062 GND 0.005676f
C1612 VDD.n1063 GND 0.004569f
C1613 VDD.n1064 GND 0.005676f
C1614 VDD.n1065 GND 0.005676f
C1615 VDD.n1066 GND 0.005676f
C1616 VDD.n1067 GND 0.004569f
C1617 VDD.n1068 GND 0.005676f
C1618 VDD.n1069 GND 0.386541f
C1619 VDD.n1070 GND 0.005676f
C1620 VDD.n1071 GND 0.004569f
C1621 VDD.n1072 GND 0.005676f
C1622 VDD.n1073 GND 0.005676f
C1623 VDD.n1074 GND 0.005676f
C1624 VDD.n1075 GND 0.004569f
C1625 VDD.n1076 GND 0.005676f
C1626 VDD.n1077 GND 0.386541f
C1627 VDD.n1078 GND 0.005676f
C1628 VDD.n1079 GND 0.004569f
C1629 VDD.n1080 GND 0.005676f
C1630 VDD.n1081 GND 0.005676f
C1631 VDD.n1082 GND 0.005676f
C1632 VDD.n1083 GND 0.004569f
C1633 VDD.n1084 GND 0.005676f
C1634 VDD.n1085 GND 0.386541f
C1635 VDD.n1086 GND 0.005676f
C1636 VDD.n1087 GND 0.004569f
C1637 VDD.n1088 GND 0.005676f
C1638 VDD.n1089 GND 0.005676f
C1639 VDD.n1090 GND 0.005676f
C1640 VDD.n1091 GND 0.004569f
C1641 VDD.n1092 GND 0.005676f
C1642 VDD.n1093 GND 0.332425f
C1643 VDD.n1094 GND 0.005676f
C1644 VDD.n1095 GND 0.004569f
C1645 VDD.n1096 GND 0.005676f
C1646 VDD.n1097 GND 0.005676f
C1647 VDD.n1098 GND 0.005676f
C1648 VDD.n1099 GND 0.004569f
C1649 VDD.n1100 GND 0.005676f
C1650 VDD.n1101 GND 0.386541f
C1651 VDD.n1102 GND 0.005676f
C1652 VDD.n1103 GND 0.004569f
C1653 VDD.n1104 GND 0.005676f
C1654 VDD.n1105 GND 0.005676f
C1655 VDD.n1106 GND 0.005676f
C1656 VDD.n1107 GND 0.004569f
C1657 VDD.n1108 GND 0.005676f
C1658 VDD.n1109 GND 0.386541f
C1659 VDD.n1110 GND 0.005676f
C1660 VDD.n1111 GND 0.004569f
C1661 VDD.n1112 GND 0.005676f
C1662 VDD.n1113 GND 0.005676f
C1663 VDD.n1114 GND 0.005676f
C1664 VDD.n1115 GND 0.004569f
C1665 VDD.n1116 GND 0.005676f
C1666 VDD.n1117 GND 0.386541f
C1667 VDD.n1118 GND 0.005676f
C1668 VDD.n1119 GND 0.004569f
C1669 VDD.n1120 GND 0.005676f
C1670 VDD.n1121 GND 0.005676f
C1671 VDD.n1122 GND 0.005676f
C1672 VDD.n1123 GND 0.004569f
C1673 VDD.n1124 GND 0.005676f
C1674 VDD.n1125 GND 0.386541f
C1675 VDD.n1126 GND 0.005676f
C1676 VDD.n1127 GND 0.004569f
C1677 VDD.n1128 GND 0.005676f
C1678 VDD.n1129 GND 0.005676f
C1679 VDD.n1130 GND 0.005676f
C1680 VDD.n1131 GND 0.004569f
C1681 VDD.n1132 GND 0.005676f
C1682 VDD.n1133 GND 0.239655f
C1683 VDD.n1134 GND 0.005676f
C1684 VDD.n1135 GND 0.004569f
C1685 VDD.n1136 GND 0.005676f
C1686 VDD.n1137 GND 0.005676f
C1687 VDD.n1138 GND 0.005676f
C1688 VDD.n1139 GND 0.005676f
C1689 VDD.n1140 GND 0.004569f
C1690 VDD.n1141 GND 0.005676f
C1691 VDD.n1142 GND 0.386541f
C1692 VDD.n1143 GND 0.005676f
C1693 VDD.n1144 GND 0.004569f
C1694 VDD.n1145 GND 0.005676f
C1695 VDD.n1146 GND 0.005676f
C1696 VDD.n1147 GND 0.005676f
C1697 VDD.n1148 GND 0.0128f
C1698 VDD.n1149 GND 0.005676f
C1699 VDD.n1150 GND 0.005676f
C1700 VDD.n1151 GND 0.004569f
C1701 VDD.n1152 GND 0.005676f
C1702 VDD.n1153 GND 0.005676f
C1703 VDD.n1154 GND 0.005676f
C1704 VDD.n1155 GND 0.005676f
C1705 VDD.n1156 GND 0.005676f
C1706 VDD.n1157 GND 0.004569f
C1707 VDD.n1158 GND 0.005676f
C1708 VDD.n1159 GND 0.005676f
C1709 VDD.n1160 GND 0.005676f
C1710 VDD.t65 GND 0.049112f
C1711 VDD.t64 GND 0.063006f
C1712 VDD.t63 GND 0.385677f
C1713 VDD.n1161 GND 0.054096f
C1714 VDD.n1162 GND 0.037762f
C1715 VDD.n1163 GND 0.005676f
C1716 VDD.n1164 GND 0.005676f
C1717 VDD.n1165 GND 0.004569f
C1718 VDD.n1166 GND 0.005676f
C1719 VDD.n1167 GND 0.005676f
C1720 VDD.n1168 GND 0.005676f
C1721 VDD.n1169 GND 0.005676f
C1722 VDD.n1170 GND 0.005676f
C1723 VDD.n1171 GND 0.004569f
C1724 VDD.n1172 GND 0.005676f
C1725 VDD.n1173 GND 0.005676f
C1726 VDD.n1174 GND 0.005676f
C1727 VDD.n1175 GND 0.005676f
C1728 VDD.n1176 GND 0.005676f
C1729 VDD.n1177 GND 0.005676f
C1730 VDD.n1178 GND 0.002467f
C1731 VDD.n1179 GND 0.004569f
C1732 VDD.n1180 GND 0.005676f
C1733 VDD.n1181 GND 0.005676f
C1734 VDD.n1182 GND 0.004569f
C1735 VDD.n1183 GND 0.004569f
C1736 VDD.n1184 GND 0.004569f
C1737 VDD.n1185 GND 0.005676f
C1738 VDD.n1186 GND 0.005676f
C1739 VDD.n1187 GND 0.005676f
C1740 VDD.n1188 GND 0.004569f
C1741 VDD.n1189 GND 0.004569f
C1742 VDD.n1190 GND 0.004569f
C1743 VDD.n1191 GND 0.005676f
C1744 VDD.n1192 GND 0.005676f
C1745 VDD.n1193 GND 0.005676f
C1746 VDD.n1194 GND 0.004158f
C1747 VDD.n1195 GND 0.00932f
C1748 VDD.n1196 GND 0.003472f
C1749 VDD.n1197 GND 0.005676f
C1750 VDD.n1198 GND 0.005676f
C1751 VDD.n1199 GND 0.005676f
C1752 VDD.n1200 GND 0.004569f
C1753 VDD.n1201 GND 0.004569f
C1754 VDD.n1202 GND 0.004569f
C1755 VDD.n1203 GND 0.005676f
C1756 VDD.n1204 GND 0.005676f
C1757 VDD.n1205 GND 0.005676f
C1758 VDD.n1206 GND 0.004569f
C1759 VDD.n1207 GND 0.004569f
C1760 VDD.n1208 GND 0.003792f
C1761 VDD.n1209 GND 0.0128f
C1762 VDD.n1210 GND 0.0128f
C1763 VDD.n1211 GND 0.005676f
C1764 VDD.n1212 GND 0.004569f
C1765 VDD.n1213 GND 0.005676f
C1766 VDD.n1214 GND 0.386541f
C1767 VDD.n1215 GND 0.005676f
C1768 VDD.n1216 GND 0.004569f
C1769 VDD.n1217 GND 0.003792f
C1770 VDD.n1218 GND 0.0128f
C1771 VDD.n1219 GND 0.0128f
C1772 VDD.n1220 GND 0.002102f
C1773 VDD.n1221 GND 0.0128f
C1774 VDD.n1223 GND 2.64587f
C1775 VDD.t109 GND 4.2017f
C1776 VDD.t10 GND 3.28946f
C1777 VDD.t85 GND 2.84494f
C1778 VDD.n1233 GND 0.00386f
C1779 VDD.t36 GND 0.042906f
C1780 VDD.t37 GND 0.059398f
C1781 VDD.t34 GND 0.475789f
C1782 VDD.n1234 GND 0.099866f
C1783 VDD.n1235 GND 0.077301f
C1784 VDD.n1236 GND 0.00386f
C1785 VDD.n1237 GND 0.00386f
C1786 VDD.n1238 GND 0.00386f
C1787 VDD.n1239 GND 0.00386f
C1788 VDD.n1240 GND 0.00386f
C1789 VDD.n1241 GND 0.00386f
C1790 VDD.n1242 GND 0.00386f
C1791 VDD.n1243 GND 0.00386f
C1792 VDD.n1244 GND 0.00386f
C1793 VDD.n1245 GND 0.00386f
C1794 VDD.n1246 GND 0.00386f
C1795 VDD.n1247 GND 0.00386f
C1796 VDD.n1248 GND 0.00386f
C1797 VDD.n1249 GND 0.00386f
C1798 VDD.n1250 GND 0.502957f
C1799 VDD.n1251 GND 0.00386f
C1800 VDD.n1252 GND 0.00386f
C1801 VDD.n1253 GND 0.502957f
C1802 VDD.n1254 GND 0.00386f
C1803 VDD.n1255 GND 0.00386f
C1804 VDD.n1256 GND 0.00386f
C1805 VDD.n1257 GND 0.00386f
C1806 VDD.n1258 GND 0.00386f
C1807 VDD.n1259 GND 0.00386f
C1808 VDD.n1260 GND 0.00386f
C1809 VDD.n1261 GND 0.00386f
C1810 VDD.n1262 GND 0.00386f
C1811 VDD.n1263 GND 0.00386f
C1812 VDD.n1264 GND 0.00386f
C1813 VDD.n1265 GND 0.00386f
C1814 VDD.n1266 GND 0.00386f
C1815 VDD.n1267 GND 0.00386f
C1816 VDD.n1268 GND 0.00386f
C1817 VDD.n1269 GND 0.002952f
C1818 VDD.n1270 GND 0.005516f
C1819 VDD.n1271 GND 0.002838f
C1820 VDD.n1272 GND 0.00386f
C1821 VDD.n1273 GND 0.00386f
C1822 VDD.n1274 GND 0.00386f
C1823 VDD.n1275 GND 0.00386f
C1824 VDD.n1276 GND 0.00386f
C1825 VDD.n1277 GND 0.00386f
C1826 VDD.n1278 GND 0.00386f
C1827 VDD.n1279 GND 0.00386f
C1828 VDD.n1280 GND 0.00386f
C1829 VDD.n1281 GND 0.00386f
C1830 VDD.n1282 GND 0.00386f
C1831 VDD.n1283 GND 0.00386f
C1832 VDD.n1284 GND 0.00386f
C1833 VDD.n1285 GND 0.00386f
C1834 VDD.n1286 GND 0.00386f
C1835 VDD.n1287 GND 0.00386f
C1836 VDD.n1288 GND 0.00386f
C1837 VDD.n1289 GND 0.00386f
C1838 VDD.n1290 GND 0.00386f
C1839 VDD.n1291 GND 0.00386f
C1840 VDD.n1292 GND 0.00386f
C1841 VDD.n1293 GND 0.00386f
C1842 VDD.n1294 GND 0.00386f
C1843 VDD.n1295 GND 0.00386f
C1844 VDD.n1296 GND 0.00386f
C1845 VDD.n1297 GND 0.00386f
C1846 VDD.n1298 GND 0.00386f
C1847 VDD.n1299 GND 0.00386f
C1848 VDD.n1300 GND 0.00386f
C1849 VDD.n1301 GND 0.00386f
C1850 VDD.n1302 GND 0.00386f
C1851 VDD.n1303 GND 0.00386f
C1852 VDD.n1304 GND 0.00386f
C1853 VDD.n1305 GND 0.00386f
C1854 VDD.n1306 GND 0.00386f
C1855 VDD.n1307 GND 0.00386f
C1856 VDD.n1308 GND 0.00386f
C1857 VDD.n1309 GND 0.00386f
C1858 VDD.n1310 GND 0.00386f
C1859 VDD.n1311 GND 0.00386f
C1860 VDD.n1312 GND 0.00386f
C1861 VDD.n1313 GND 0.00386f
C1862 VDD.n1314 GND 0.00386f
C1863 VDD.n1315 GND 0.00386f
C1864 VDD.n1316 GND 0.00386f
C1865 VDD.n1317 GND 0.00386f
C1866 VDD.n1318 GND 0.00386f
C1867 VDD.n1319 GND 0.00386f
C1868 VDD.n1320 GND 0.00386f
C1869 VDD.n1321 GND 0.00386f
C1870 VDD.n1322 GND 0.00386f
C1871 VDD.n1323 GND 0.00386f
C1872 VDD.n1324 GND 0.00386f
C1873 VDD.n1325 GND 0.00386f
C1874 VDD.n1326 GND 0.00386f
C1875 VDD.n1327 GND 0.00386f
C1876 VDD.n1328 GND 0.00386f
C1877 VDD.n1329 GND 0.00386f
C1878 VDD.n1330 GND 0.00386f
C1879 VDD.n1331 GND 0.00386f
C1880 VDD.n1332 GND 0.00386f
C1881 VDD.n1333 GND 0.00386f
C1882 VDD.n1334 GND 0.00386f
C1883 VDD.n1335 GND 0.00386f
C1884 VDD.n1336 GND 0.00386f
C1885 VDD.n1337 GND 0.00386f
C1886 VDD.n1338 GND 0.00386f
C1887 VDD.n1339 GND 0.00386f
C1888 VDD.n1340 GND 0.00386f
C1889 VDD.n1341 GND 0.00386f
C1890 VDD.n1342 GND 0.00386f
C1891 VDD.n1343 GND 0.00386f
C1892 VDD.n1344 GND 0.00386f
C1893 VDD.n1345 GND 0.00386f
C1894 VDD.n1346 GND 0.00386f
C1895 VDD.n1347 GND 0.00386f
C1896 VDD.n1348 GND 0.00386f
C1897 VDD.n1349 GND 0.00386f
C1898 VDD.n1350 GND 0.00386f
C1899 VDD.n1351 GND 0.00386f
C1900 VDD.n1352 GND 0.00386f
C1901 VDD.n1353 GND 0.00386f
C1902 VDD.n1354 GND 0.00386f
C1903 VDD.n1355 GND 0.00386f
C1904 VDD.n1356 GND 0.00386f
C1905 VDD.n1357 GND 0.00386f
C1906 VDD.n1358 GND 0.00386f
C1907 VDD.n1359 GND 0.00386f
C1908 VDD.n1360 GND 0.009102f
C1909 VDD.n1361 GND 0.009516f
C1910 VDD.n1362 GND 0.009516f
C1911 VDD.n1373 GND 0.00386f
C1912 VDD.t77 GND 0.042906f
C1913 VDD.t78 GND 0.059398f
C1914 VDD.t76 GND 0.475789f
C1915 VDD.n1374 GND 0.099866f
C1916 VDD.n1375 GND 0.077301f
C1917 VDD.n1376 GND 0.005516f
C1918 VDD.n1377 GND 0.00386f
C1919 VDD.n1378 GND 0.00386f
C1920 VDD.n1379 GND 0.00386f
C1921 VDD.n1380 GND 0.00386f
C1922 VDD.n1381 GND 0.00386f
C1923 VDD.n1382 GND 0.00386f
C1924 VDD.n1383 GND 0.00386f
C1925 VDD.n1384 GND 0.00386f
C1926 VDD.n1385 GND 0.00386f
C1927 VDD.n1386 GND 0.00386f
C1928 VDD.n1387 GND 0.00386f
C1929 VDD.n1388 GND 0.00386f
C1930 VDD.n1389 GND 0.00386f
C1931 VDD.n1390 GND 0.00386f
C1932 VDD.n1391 GND 0.00386f
C1933 VDD.n1392 GND 0.00386f
C1934 VDD.n1393 GND 0.00386f
C1935 VDD.n1394 GND 0.00386f
C1936 VDD.n1395 GND 0.00386f
C1937 VDD.n1396 GND 0.00386f
C1938 VDD.n1397 GND 0.00386f
C1939 VDD.n1398 GND 0.00386f
C1940 VDD.n1399 GND 0.00386f
C1941 VDD.n1400 GND 0.00386f
C1942 VDD.n1401 GND 0.00386f
C1943 VDD.n1402 GND 0.00386f
C1944 VDD.n1403 GND 0.00386f
C1945 VDD.n1404 GND 0.00386f
C1946 VDD.n1405 GND 0.00386f
C1947 VDD.n1406 GND 0.00386f
C1948 VDD.n1407 GND 0.00386f
C1949 VDD.n1408 GND 0.00386f
C1950 VDD.n1409 GND 0.00386f
C1951 VDD.n1410 GND 0.00386f
C1952 VDD.n1411 GND 0.00386f
C1953 VDD.n1412 GND 0.00386f
C1954 VDD.n1413 GND 0.00386f
C1955 VDD.n1414 GND 0.00386f
C1956 VDD.n1415 GND 0.00386f
C1957 VDD.n1416 GND 0.00386f
C1958 VDD.n1417 GND 0.00386f
C1959 VDD.n1418 GND 0.00386f
C1960 VDD.n1419 GND 0.00386f
C1961 VDD.n1420 GND 0.00386f
C1962 VDD.n1421 GND 0.00386f
C1963 VDD.n1422 GND 0.00386f
C1964 VDD.n1423 GND 0.00386f
C1965 VDD.n1424 GND 0.00386f
C1966 VDD.n1425 GND 0.00386f
C1967 VDD.n1426 GND 0.00386f
C1968 VDD.n1427 GND 0.00386f
C1969 VDD.n1428 GND 0.00386f
C1970 VDD.n1429 GND 0.00386f
C1971 VDD.n1430 GND 0.00386f
C1972 VDD.n1431 GND 0.00386f
C1973 VDD.n1432 GND 0.00386f
C1974 VDD.n1433 GND 0.00386f
C1975 VDD.n1434 GND 0.00386f
C1976 VDD.n1435 GND 0.00386f
C1977 VDD.n1436 GND 0.00386f
C1978 VDD.n1437 GND 0.00386f
C1979 VDD.n1438 GND 0.00386f
C1980 VDD.n1439 GND 0.00386f
C1981 VDD.n1440 GND 0.00386f
C1982 VDD.n1441 GND 0.00386f
C1983 VDD.n1442 GND 0.00386f
C1984 VDD.n1443 GND 0.00386f
C1985 VDD.n1444 GND 0.00386f
C1986 VDD.n1445 GND 0.00386f
C1987 VDD.n1446 GND 0.00386f
C1988 VDD.n1447 GND 0.00386f
C1989 VDD.n1448 GND 0.00386f
C1990 VDD.n1449 GND 0.00386f
C1991 VDD.n1450 GND 0.00386f
C1992 VDD.n1451 GND 0.00386f
C1993 VDD.n1452 GND 0.00386f
C1994 VDD.n1453 GND 0.00386f
C1995 VDD.n1454 GND 0.00386f
C1996 VDD.n1455 GND 0.00386f
C1997 VDD.n1456 GND 0.00386f
C1998 VDD.n1457 GND 0.00386f
C1999 VDD.n1458 GND 0.00386f
C2000 VDD.n1459 GND 0.00386f
C2001 VDD.n1460 GND 0.00386f
C2002 VDD.n1461 GND 0.00386f
C2003 VDD.n1462 GND 0.00386f
C2004 VDD.n1463 GND 0.00386f
C2005 VDD.n1464 GND 0.00386f
C2006 VDD.n1465 GND 0.00386f
C2007 VDD.n1466 GND 0.00386f
C2008 VDD.n1467 GND 0.009102f
C2009 VDD.n1468 GND 0.009516f
C2010 VDD.n1469 GND 0.009516f
C2011 VDD.n1470 GND 0.002838f
C2012 VDD.n1471 GND 0.00386f
C2013 VDD.n1472 GND 0.00386f
C2014 VDD.n1473 GND 0.002952f
C2015 VDD.n1474 GND 0.00386f
C2016 VDD.n1475 GND 0.00386f
C2017 VDD.n1476 GND 0.00386f
C2018 VDD.n1477 GND 0.00386f
C2019 VDD.n1478 GND 0.00386f
C2020 VDD.n1479 GND 0.00386f
C2021 VDD.n1480 GND 0.00386f
C2022 VDD.n1481 GND 0.00386f
C2023 VDD.n1482 GND 0.00386f
C2024 VDD.n1483 GND 0.00386f
C2025 VDD.n1484 GND 0.00386f
C2026 VDD.n1485 GND 0.00386f
C2027 VDD.n1486 GND 0.00386f
C2028 VDD.n1487 GND 0.00386f
C2029 VDD.n1488 GND 0.00386f
C2030 VDD.n1489 GND 0.508633f
C2031 VDD.n1490 GND 0.508633f
C2032 VDD.n1491 GND 0.00386f
C2033 VDD.n1492 GND 0.00386f
C2034 VDD.n1493 GND 0.00386f
C2035 VDD.n1494 GND 0.00386f
C2036 VDD.n1495 GND 0.00386f
C2037 VDD.n1496 GND 0.00386f
C2038 VDD.n1497 GND 0.00386f
C2039 VDD.n1498 GND 0.00386f
C2040 VDD.n1499 GND 0.00386f
C2041 VDD.n1500 GND 0.00386f
C2042 VDD.n1501 GND 0.00386f
C2043 VDD.n1502 GND 0.00386f
C2044 VDD.n1503 GND 0.00386f
C2045 VDD.n1504 GND 0.00386f
C2046 VDD.n1505 GND 0.00386f
C2047 VDD.n1506 GND 0.00386f
C2048 VDD.n1507 GND 0.00386f
C2049 VDD.n1508 GND 0.00386f
C2050 VDD.n1510 GND 1.43407f
C2051 VDD.n1512 GND 0.00386f
C2052 VDD.n1513 GND 0.00386f
C2053 VDD.n1514 GND 0.009516f
C2054 VDD.n1515 GND 0.009102f
C2055 VDD.n1516 GND 0.009102f
C2056 VDD.n1517 GND 0.35755f
C2057 VDD.n1518 GND 0.009102f
C2058 VDD.n1519 GND 0.009102f
C2059 VDD.n1520 GND 0.00386f
C2060 VDD.n1521 GND 0.00386f
C2061 VDD.n1522 GND 0.00386f
C2062 VDD.n1523 GND 0.262848f
C2063 VDD.n1524 GND 0.00386f
C2064 VDD.n1525 GND 0.00386f
C2065 VDD.n1526 GND 0.00386f
C2066 VDD.n1527 GND 0.00386f
C2067 VDD.n1528 GND 0.00386f
C2068 VDD.n1529 GND 0.262848f
C2069 VDD.n1530 GND 0.00386f
C2070 VDD.n1531 GND 0.00386f
C2071 VDD.n1532 GND 0.00386f
C2072 VDD.n1533 GND 0.00386f
C2073 VDD.n1534 GND 0.00386f
C2074 VDD.n1535 GND 0.19327f
C2075 VDD.n1536 GND 0.00386f
C2076 VDD.n1537 GND 0.00386f
C2077 VDD.n1538 GND 0.00386f
C2078 VDD.n1539 GND 0.00386f
C2079 VDD.n1540 GND 0.00386f
C2080 VDD.n1541 GND 0.262848f
C2081 VDD.n1542 GND 0.00386f
C2082 VDD.n1543 GND 0.00386f
C2083 VDD.n1544 GND 0.00386f
C2084 VDD.n1545 GND 0.00386f
C2085 VDD.n1546 GND 0.00386f
C2086 VDD.n1547 GND 0.237723f
C2087 VDD.n1548 GND 0.00386f
C2088 VDD.n1549 GND 0.00386f
C2089 VDD.n1550 GND 0.00386f
C2090 VDD.n1551 GND 0.00386f
C2091 VDD.n1552 GND 0.00386f
C2092 VDD.n1553 GND 0.262848f
C2093 VDD.n1554 GND 0.00386f
C2094 VDD.n1555 GND 0.00386f
C2095 VDD.n1556 GND 0.00386f
C2096 VDD.n1557 GND 0.00386f
C2097 VDD.n1558 GND 0.00386f
C2098 VDD.n1559 GND 0.262848f
C2099 VDD.n1560 GND 0.00386f
C2100 VDD.n1561 GND 0.00386f
C2101 VDD.n1562 GND 0.00386f
C2102 VDD.n1563 GND 0.00386f
C2103 VDD.n1564 GND 0.00386f
C2104 VDD.n1565 GND 0.262848f
C2105 VDD.n1566 GND 0.00386f
C2106 VDD.n1567 GND 0.00386f
C2107 VDD.n1568 GND 0.00386f
C2108 VDD.n1569 GND 0.00386f
C2109 VDD.n1570 GND 0.00386f
C2110 VDD.n1571 GND 0.262848f
C2111 VDD.n1572 GND 0.00386f
C2112 VDD.n1573 GND 0.00386f
C2113 VDD.n1574 GND 0.00386f
C2114 VDD.n1575 GND 0.00386f
C2115 VDD.n1576 GND 0.00386f
C2116 VDD.n1577 GND 0.208732f
C2117 VDD.n1578 GND 0.00386f
C2118 VDD.n1579 GND 0.00386f
C2119 VDD.n1580 GND 0.00386f
C2120 VDD.n1581 GND 0.00386f
C2121 VDD.n1582 GND 0.00386f
C2122 VDD.n1583 GND 0.262848f
C2123 VDD.n1584 GND 0.00386f
C2124 VDD.n1585 GND 0.00386f
C2125 VDD.n1586 GND 0.00386f
C2126 VDD.n1587 GND 0.00386f
C2127 VDD.n1588 GND 0.00386f
C2128 VDD.n1589 GND 0.262848f
C2129 VDD.n1590 GND 0.00386f
C2130 VDD.n1591 GND 0.00386f
C2131 VDD.n1592 GND 0.00386f
C2132 VDD.n1593 GND 0.00386f
C2133 VDD.n1594 GND 0.00386f
C2134 VDD.n1595 GND 0.172011f
C2135 VDD.n1596 GND 0.00386f
C2136 VDD.n1597 GND 0.00386f
C2137 VDD.n1598 GND 0.00386f
C2138 VDD.n1599 GND 0.00386f
C2139 VDD.n1600 GND 0.00386f
C2140 VDD.n1601 GND 0.262848f
C2141 VDD.n1602 GND 0.00386f
C2142 VDD.n1603 GND 0.00386f
C2143 VDD.n1604 GND 0.00386f
C2144 VDD.n1605 GND 0.00386f
C2145 VDD.n1606 GND 0.00386f
C2146 VDD.n1607 GND 0.262848f
C2147 VDD.n1608 GND 0.00386f
C2148 VDD.n1609 GND 0.00386f
C2149 VDD.n1610 GND 0.00386f
C2150 VDD.n1611 GND 0.00386f
C2151 VDD.n1612 GND 0.00386f
C2152 VDD.n1613 GND 0.197136f
C2153 VDD.n1614 GND 0.00386f
C2154 VDD.n1615 GND 0.00386f
C2155 VDD.n1616 GND 0.00386f
C2156 VDD.n1617 GND 0.00386f
C2157 VDD.n1618 GND 0.00386f
C2158 VDD.n1619 GND 0.262848f
C2159 VDD.n1620 GND 0.00386f
C2160 VDD.n1621 GND 0.00386f
C2161 VDD.n1622 GND 0.00386f
C2162 VDD.n1623 GND 0.00386f
C2163 VDD.n1624 GND 0.00386f
C2164 VDD.n1625 GND 0.210665f
C2165 VDD.n1626 GND 0.00386f
C2166 VDD.n1627 GND 0.00386f
C2167 VDD.n1628 GND 0.00386f
C2168 VDD.n1629 GND 0.00386f
C2169 VDD.n1630 GND 0.00386f
C2170 VDD.n1631 GND 0.262848f
C2171 VDD.n1632 GND 0.00386f
C2172 VDD.n1633 GND 0.00386f
C2173 VDD.n1634 GND 0.00386f
C2174 VDD.n1635 GND 0.00386f
C2175 VDD.n1636 GND 0.00386f
C2176 VDD.n1637 GND 0.262848f
C2177 VDD.n1638 GND 0.00386f
C2178 VDD.n1639 GND 0.00386f
C2179 VDD.n1640 GND 0.00386f
C2180 VDD.n1641 GND 0.00386f
C2181 VDD.n1642 GND 0.00386f
C2182 VDD.n1643 GND 0.18554f
C2183 VDD.n1644 GND 0.00386f
C2184 VDD.n1645 GND 0.00386f
C2185 VDD.n1646 GND 0.00386f
C2186 VDD.n1647 GND 0.00386f
C2187 VDD.n1648 GND 0.00386f
C2188 VDD.n1649 GND 0.262848f
C2189 VDD.n1650 GND 0.00386f
C2190 VDD.n1651 GND 0.00386f
C2191 VDD.n1652 GND 0.00386f
C2192 VDD.n1653 GND 0.00386f
C2193 VDD.n1654 GND 0.00386f
C2194 VDD.n1655 GND 0.262848f
C2195 VDD.n1656 GND 0.00386f
C2196 VDD.n1657 GND 0.00386f
C2197 VDD.n1658 GND 0.00386f
C2198 VDD.n1659 GND 0.00386f
C2199 VDD.n1660 GND 0.00386f
C2200 VDD.n1661 GND 0.195203f
C2201 VDD.n1662 GND 0.00386f
C2202 VDD.n1663 GND 0.00386f
C2203 VDD.n1664 GND 0.00386f
C2204 VDD.n1665 GND 0.00386f
C2205 VDD.n1666 GND 0.00386f
C2206 VDD.n1667 GND 0.262848f
C2207 VDD.n1668 GND 0.00386f
C2208 VDD.n1669 GND 0.00386f
C2209 VDD.n1670 GND 0.00386f
C2210 VDD.n1671 GND 0.00386f
C2211 VDD.n1672 GND 0.00386f
C2212 VDD.n1673 GND 0.262848f
C2213 VDD.n1674 GND 0.00386f
C2214 VDD.n1675 GND 0.00386f
C2215 VDD.n1676 GND 0.00386f
C2216 VDD.n1677 GND 0.00386f
C2217 VDD.n1678 GND 0.00386f
C2218 VDD.n1679 GND 0.262848f
C2219 VDD.n1680 GND 0.00386f
C2220 VDD.n1681 GND 0.00386f
C2221 VDD.n1682 GND 0.00386f
C2222 VDD.n1683 GND 0.00386f
C2223 VDD.n1684 GND 0.00386f
C2224 VDD.n1685 GND 0.201001f
C2225 VDD.n1686 GND 0.00386f
C2226 VDD.n1687 GND 0.00386f
C2227 VDD.n1688 GND 0.00386f
C2228 VDD.t47 GND 0.042906f
C2229 VDD.t46 GND 0.059398f
C2230 VDD.t44 GND 0.475789f
C2231 VDD.n1689 GND 0.099866f
C2232 VDD.n1690 GND 0.077301f
C2233 VDD.n1691 GND 0.005516f
C2234 VDD.n1692 GND 0.00386f
C2235 VDD.n1693 GND 0.002952f
C2236 VDD.n1694 GND 0.00386f
C2237 VDD.n1695 GND 0.00386f
C2238 VDD.n1696 GND 0.00386f
C2239 VDD.n1697 GND 0.00386f
C2240 VDD.n1698 GND 0.00386f
C2241 VDD.n1699 GND 0.00386f
C2242 VDD.n1700 GND 0.00386f
C2243 VDD.n1701 GND 0.00386f
C2244 VDD.n1702 GND 0.00386f
C2245 VDD.n1703 GND 0.00386f
C2246 VDD.n1704 GND 0.00386f
C2247 VDD.n1705 GND 0.00386f
C2248 VDD.n1706 GND 0.00386f
C2249 VDD.n1707 GND 0.00386f
C2250 VDD.n1708 GND 0.00386f
C2251 VDD.n1709 GND 0.00386f
C2252 VDD.n1710 GND 0.00386f
C2253 VDD.n1711 GND 0.00386f
C2254 VDD.n1712 GND 0.00386f
C2255 VDD.n1713 GND 0.00386f
C2256 VDD.n1714 GND 0.00386f
C2257 VDD.n1715 GND 0.00386f
C2258 VDD.n1716 GND 0.00386f
C2259 VDD.n1717 GND 0.00386f
C2260 VDD.n1718 GND 0.00386f
C2261 VDD.n1719 GND 0.00386f
C2262 VDD.n1720 GND 0.00386f
C2263 VDD.n1721 GND 0.00386f
C2264 VDD.n1722 GND 0.00386f
C2265 VDD.n1723 GND 0.00386f
C2266 VDD.n1724 GND 0.00386f
C2267 VDD.n1725 GND 0.00386f
C2268 VDD.n1726 GND 0.00386f
C2269 VDD.n1727 GND 0.00386f
C2270 VDD.n1728 GND 0.00386f
C2271 VDD.n1729 GND 0.00386f
C2272 VDD.n1730 GND 0.009516f
C2273 VDD.n1731 GND 0.009516f
C2274 VDD.n1732 GND 0.009102f
C2275 VDD.n1733 GND 0.009102f
C2276 VDD.n1734 GND 0.00386f
C2277 VDD.n1735 GND 0.00386f
C2278 VDD.n1736 GND 0.00386f
C2279 VDD.n1737 GND 0.00386f
C2280 VDD.n1738 GND 0.00386f
C2281 VDD.n1739 GND 0.00386f
C2282 VDD.n1740 GND 0.00386f
C2283 VDD.n1741 GND 0.187472f
C2284 VDD.n1742 GND 0.00386f
C2285 VDD.n1743 GND 0.00386f
C2286 VDD.n1744 GND 0.00386f
C2287 VDD.n1745 GND 0.00386f
C2288 VDD.n1746 GND 0.00386f
C2289 VDD.n1747 GND 0.262848f
C2290 VDD.n1748 GND 0.00386f
C2291 VDD.n1749 GND 0.00386f
C2292 VDD.n1750 GND 0.00386f
C2293 VDD.n1751 GND 0.00386f
C2294 VDD.n1752 GND 0.009538f
C2295 VDD.n1753 GND 0.009102f
C2296 VDD.n1754 GND 0.009516f
C2297 VDD.n1755 GND 0.009081f
C2298 VDD.n1756 GND 0.002838f
C2299 VDD.n1757 GND 0.00386f
C2300 VDD.n1758 GND 0.00386f
C2301 VDD.n1759 GND 0.002952f
C2302 VDD.n1760 GND 0.00386f
C2303 VDD.n1761 GND 0.00386f
C2304 VDD.n1762 GND 0.00386f
C2305 VDD.n1763 GND 0.00386f
C2306 VDD.n1764 GND 0.00386f
C2307 VDD.n1765 GND 0.00386f
C2308 VDD.n1766 GND 0.00386f
C2309 VDD.n1767 GND 0.00386f
C2310 VDD.n1768 GND 0.00386f
C2311 VDD.n1769 GND 0.00386f
C2312 VDD.n1770 GND 0.00386f
C2313 VDD.n1771 GND 0.00386f
C2314 VDD.n1772 GND 0.00386f
C2315 VDD.n1773 GND 0.00386f
C2316 VDD.n1774 GND 0.00386f
C2317 VDD.n1775 GND 0.00386f
C2318 VDD.n1776 GND 0.00386f
C2319 VDD.n1777 GND 0.00386f
C2320 VDD.n1778 GND 0.00386f
C2321 VDD.n1779 GND 0.00386f
C2322 VDD.n1780 GND 0.00386f
C2323 VDD.n1781 GND 0.00386f
C2324 VDD.n1782 GND 0.00386f
C2325 VDD.n1783 GND 0.00386f
C2326 VDD.n1784 GND 0.00386f
C2327 VDD.n1785 GND 0.00386f
C2328 VDD.n1786 GND 0.00386f
C2329 VDD.n1787 GND 0.00386f
C2330 VDD.n1788 GND 0.00386f
C2331 VDD.n1789 GND 0.00386f
C2332 VDD.n1790 GND 0.00386f
C2333 VDD.n1791 GND 0.00386f
C2334 VDD.n1792 GND 0.00386f
C2335 VDD.n1793 GND 0.00386f
C2336 VDD.n1794 GND 0.00386f
C2337 VDD.n1795 GND 0.00386f
C2338 VDD.n1796 GND 0.009516f
C2339 VDD.n1797 GND 0.009516f
C2340 VDD.n1798 GND 0.009102f
C2341 VDD.n1799 GND 0.00386f
C2342 VDD.n1800 GND 0.00386f
C2343 VDD.n1801 GND 0.262848f
C2344 VDD.n1802 GND 0.00386f
C2345 VDD.n1803 GND 0.00386f
C2346 VDD.n1804 GND 0.009538f
C2347 VDD.n1805 GND 0.009081f
C2348 VDD.n1806 GND 0.009516f
C2349 VDD.n1808 GND 1.65246f
C2350 VDD.n1809 GND 1.65246f
C2351 VDD.n1810 GND 0.009102f
C2352 VDD.n1811 GND 0.009516f
C2353 VDD.n1812 GND 0.00386f
C2354 VDD.t50 GND 0.042906f
C2355 VDD.t51 GND 0.059398f
C2356 VDD.t48 GND 0.475789f
C2357 VDD.n1813 GND 0.099866f
C2358 VDD.n1814 GND 0.077301f
C2359 VDD.n1815 GND 0.005516f
C2360 VDD.n1816 GND 0.002952f
C2361 VDD.n1817 GND 0.00386f
C2362 VDD.n1818 GND 0.00386f
C2363 VDD.n1819 GND 0.00386f
C2364 VDD.n1820 GND 0.00386f
C2365 VDD.n1821 GND 0.00386f
C2366 VDD.n1822 GND 0.00386f
C2367 VDD.n1823 GND 0.00386f
C2368 VDD.n1824 GND 0.00386f
C2369 VDD.n1826 GND 0.00386f
C2370 VDD.n1827 GND 0.00386f
C2371 VDD.n1828 GND 0.00386f
C2372 VDD.n1829 GND 0.00386f
C2373 VDD.n1831 GND 0.00386f
C2374 VDD.n1833 GND 0.00386f
C2375 VDD.n1834 GND 0.00386f
C2376 VDD.n1835 GND 0.00386f
C2377 VDD.n1836 GND 0.00386f
C2378 VDD.n1837 GND 0.00386f
C2379 VDD.n1839 GND 0.00386f
C2380 VDD.n1841 GND 0.00386f
C2381 VDD.n1842 GND 0.00386f
C2382 VDD.n1843 GND 0.00386f
C2383 VDD.n1844 GND 0.00386f
C2384 VDD.n1845 GND 0.00386f
C2385 VDD.n1847 GND 0.00386f
C2386 VDD.n1849 GND 0.00386f
C2387 VDD.n1850 GND 0.00386f
C2388 VDD.n1851 GND 0.00386f
C2389 VDD.n1852 GND 0.00386f
C2390 VDD.n1853 GND 0.00386f
C2391 VDD.n1855 GND 0.00386f
C2392 VDD.n1857 GND 0.00386f
C2393 VDD.n1858 GND 0.00386f
C2394 VDD.n1859 GND 0.00386f
C2395 VDD.n1860 GND 0.00386f
C2396 VDD.n1861 GND 0.00386f
C2397 VDD.n1863 GND 0.00386f
C2398 VDD.n1865 GND 0.00386f
C2399 VDD.n1866 GND 0.002838f
C2400 VDD.n1867 GND 0.009516f
C2401 VDD.n1868 GND 0.00386f
C2402 VDD.n1869 GND 0.00386f
C2403 VDD.n1870 GND 0.00386f
C2404 VDD.n1871 GND 0.00386f
C2405 VDD.n1872 GND 0.00386f
C2406 VDD.n1873 GND 0.00386f
C2407 VDD.n1874 GND 0.00386f
C2408 VDD.n1875 GND 0.00386f
C2409 VDD.n1876 GND 0.00386f
C2410 VDD.n1877 GND 0.00386f
C2411 VDD.n1878 GND 0.00386f
C2412 VDD.n1879 GND 0.00386f
C2413 VDD.n1880 GND 0.00386f
C2414 VDD.n1881 GND 0.00386f
C2415 VDD.n1882 GND 0.00386f
C2416 VDD.n1883 GND 0.00386f
C2417 VDD.n1884 GND 0.00386f
C2418 VDD.n1885 GND 0.00386f
C2419 VDD.n1886 GND 0.00386f
C2420 VDD.n1887 GND 0.00386f
C2421 VDD.n1888 GND 0.00386f
C2422 VDD.n1889 GND 0.00386f
C2423 VDD.n1890 GND 0.00386f
C2424 VDD.n1891 GND 0.00386f
C2425 VDD.n1892 GND 0.00386f
C2426 VDD.n1893 GND 0.00386f
C2427 VDD.n1894 GND 0.00386f
C2428 VDD.n1895 GND 0.00386f
C2429 VDD.n1896 GND 0.00386f
C2430 VDD.n1897 GND 0.00386f
C2431 VDD.n1898 GND 0.00386f
C2432 VDD.n1899 GND 0.00386f
C2433 VDD.n1900 GND 0.00386f
C2434 VDD.n1901 GND 0.00386f
C2435 VDD.n1902 GND 0.00386f
C2436 VDD.n1903 GND 0.00386f
C2437 VDD.n1904 GND 0.00386f
C2438 VDD.n1905 GND 0.00386f
C2439 VDD.n1906 GND 0.00386f
C2440 VDD.n1907 GND 0.00386f
C2441 VDD.n1908 GND 0.00386f
C2442 VDD.n1909 GND 0.00386f
C2443 VDD.n1910 GND 0.00386f
C2444 VDD.n1911 GND 0.00386f
C2445 VDD.n1912 GND 0.00386f
C2446 VDD.n1913 GND 0.00386f
C2447 VDD.n1914 GND 0.00386f
C2448 VDD.n1915 GND 0.00386f
C2449 VDD.n1916 GND 0.00386f
C2450 VDD.n1917 GND 0.00386f
C2451 VDD.n1918 GND 0.00386f
C2452 VDD.n1919 GND 0.00386f
C2453 VDD.n1920 GND 0.00386f
C2454 VDD.n1921 GND 0.00386f
C2455 VDD.n1922 GND 0.00386f
C2456 VDD.n1923 GND 0.00386f
C2457 VDD.n1924 GND 0.00386f
C2458 VDD.n1925 GND 0.00386f
C2459 VDD.n1926 GND 0.00386f
C2460 VDD.n1927 GND 0.00386f
C2461 VDD.n1928 GND 0.00386f
C2462 VDD.n1929 GND 0.00386f
C2463 VDD.n1930 GND 0.00386f
C2464 VDD.n1931 GND 0.00386f
C2465 VDD.n1932 GND 0.00386f
C2466 VDD.n1933 GND 0.00386f
C2467 VDD.n1934 GND 0.00386f
C2468 VDD.n1935 GND 0.00386f
C2469 VDD.n1936 GND 0.00386f
C2470 VDD.n1937 GND 0.00386f
C2471 VDD.n1938 GND 0.00386f
C2472 VDD.n1939 GND 0.00386f
C2473 VDD.n1940 GND 0.00386f
C2474 VDD.n1941 GND 0.00386f
C2475 VDD.n1942 GND 0.00386f
C2476 VDD.n1943 GND 0.00386f
C2477 VDD.n1944 GND 0.00386f
C2478 VDD.n1945 GND 0.00386f
C2479 VDD.n1946 GND 0.00386f
C2480 VDD.n1947 GND 0.00386f
C2481 VDD.n1948 GND 0.00386f
C2482 VDD.n1949 GND 0.00386f
C2483 VDD.n1950 GND 0.00386f
C2484 VDD.n1951 GND 0.00386f
C2485 VDD.n1952 GND 0.00386f
C2486 VDD.n1953 GND 0.00386f
C2487 VDD.n1954 GND 0.00386f
C2488 VDD.n1955 GND 0.00386f
C2489 VDD.n1956 GND 0.00386f
C2490 VDD.n1957 GND 0.009102f
C2491 VDD.n1958 GND 0.009102f
C2492 VDD.n1959 GND 0.009516f
C2493 VDD.n1960 GND 0.00386f
C2494 VDD.n1962 GND 0.00386f
C2495 VDD.n1963 GND 0.00386f
C2496 VDD.n1964 GND 0.00386f
C2497 VDD.n1965 GND 0.00386f
C2498 VDD.n1966 GND 0.00386f
C2499 VDD.n1967 GND 0.00386f
C2500 VDD.n1968 GND 0.00386f
C2501 VDD.n1969 GND 0.00386f
C2502 VDD.t80 GND 0.042906f
C2503 VDD.t81 GND 0.059398f
C2504 VDD.t79 GND 0.475789f
C2505 VDD.n1970 GND 0.099866f
C2506 VDD.n1971 GND 0.077301f
C2507 VDD.n1972 GND 0.00386f
C2508 VDD.n1973 GND 0.00386f
C2509 VDD.n1974 GND 0.00386f
C2510 VDD.n1975 GND 0.00386f
C2511 VDD.n1976 GND 0.00386f
C2512 VDD.n1977 GND 0.00386f
C2513 VDD.n1978 GND 0.00386f
C2514 VDD.n1979 GND 0.00386f
C2515 VDD.n1980 GND 0.00386f
C2516 VDD.n1981 GND 0.00386f
C2517 VDD.n1982 GND 0.00386f
C2518 VDD.n1983 GND 0.00386f
C2519 VDD.n1984 GND 0.00386f
C2520 VDD.n1985 GND 0.00386f
C2521 VDD.n1986 GND 0.00386f
C2522 VDD.n1987 GND 0.00386f
C2523 VDD.n1988 GND 0.00386f
C2524 VDD.n1989 GND 0.00386f
C2525 VDD.n1990 GND 0.00386f
C2526 VDD.n1991 GND 0.00386f
C2527 VDD.n1992 GND 0.00386f
C2528 VDD.n1993 GND 0.00386f
C2529 VDD.n1994 GND 0.00386f
C2530 VDD.n1995 GND 0.00386f
C2531 VDD.n1996 GND 0.00386f
C2532 VDD.n1997 GND 0.00386f
C2533 VDD.n1998 GND 0.00386f
C2534 VDD.n1999 GND 0.00386f
C2535 VDD.n2000 GND 0.00386f
C2536 VDD.n2001 GND 0.00386f
C2537 VDD.n2002 GND 0.00386f
C2538 VDD.n2003 GND 0.00386f
C2539 VDD.n2004 GND 0.00386f
C2540 VDD.n2005 GND 0.00386f
C2541 VDD.n2006 GND 0.00386f
C2542 VDD.n2007 GND 0.00386f
C2543 VDD.n2008 GND 0.00386f
C2544 VDD.n2009 GND 0.00386f
C2545 VDD.n2010 GND 0.00386f
C2546 VDD.n2011 GND 0.00386f
C2547 VDD.n2012 GND 0.00386f
C2548 VDD.n2013 GND 0.00386f
C2549 VDD.n2014 GND 0.00386f
C2550 VDD.n2015 GND 0.00386f
C2551 VDD.n2016 GND 0.00386f
C2552 VDD.n2017 GND 0.00386f
C2553 VDD.n2018 GND 0.00386f
C2554 VDD.n2019 GND 0.00386f
C2555 VDD.n2020 GND 0.00386f
C2556 VDD.n2021 GND 0.00386f
C2557 VDD.n2022 GND 0.00386f
C2558 VDD.n2023 GND 0.00386f
C2559 VDD.n2024 GND 0.00386f
C2560 VDD.n2025 GND 0.00386f
C2561 VDD.n2026 GND 0.00386f
C2562 VDD.n2027 GND 0.00386f
C2563 VDD.n2028 GND 0.00386f
C2564 VDD.n2029 GND 0.00386f
C2565 VDD.n2030 GND 0.00386f
C2566 VDD.n2031 GND 0.00386f
C2567 VDD.n2032 GND 0.00386f
C2568 VDD.n2033 GND 0.00386f
C2569 VDD.n2034 GND 0.00386f
C2570 VDD.n2035 GND 0.00386f
C2571 VDD.n2036 GND 0.00386f
C2572 VDD.n2037 GND 0.00386f
C2573 VDD.n2038 GND 0.00386f
C2574 VDD.n2039 GND 0.00386f
C2575 VDD.n2040 GND 0.00386f
C2576 VDD.n2041 GND 0.00386f
C2577 VDD.n2042 GND 0.00386f
C2578 VDD.n2043 GND 0.00386f
C2579 VDD.n2044 GND 0.00386f
C2580 VDD.n2045 GND 0.00386f
C2581 VDD.n2046 GND 0.00386f
C2582 VDD.n2047 GND 0.00386f
C2583 VDD.n2048 GND 0.00386f
C2584 VDD.n2049 GND 0.00386f
C2585 VDD.n2050 GND 0.00386f
C2586 VDD.n2051 GND 0.00386f
C2587 VDD.n2052 GND 0.00386f
C2588 VDD.n2053 GND 0.00386f
C2589 VDD.n2054 GND 0.00386f
C2590 VDD.n2055 GND 0.00386f
C2591 VDD.n2056 GND 0.00386f
C2592 VDD.n2057 GND 0.00386f
C2593 VDD.n2058 GND 0.00386f
C2594 VDD.n2059 GND 0.00386f
C2595 VDD.n2060 GND 0.009102f
C2596 VDD.n2061 GND 0.009516f
C2597 VDD.n2062 GND 0.009516f
C2598 VDD.n2064 GND 0.00386f
C2599 VDD.n2065 GND 0.002838f
C2600 VDD.n2066 GND 0.005516f
C2601 VDD.n2067 GND 0.002952f
C2602 VDD.n2068 GND 0.00386f
C2603 VDD.n2069 GND 0.00386f
C2604 VDD.n2071 GND 0.00386f
C2605 VDD.n2073 GND 0.00386f
C2606 VDD.n2074 GND 0.00386f
C2607 VDD.n2075 GND 0.00386f
C2608 VDD.n2076 GND 0.00386f
C2609 VDD.n2077 GND 0.00386f
C2610 VDD.n2079 GND 0.00386f
C2611 VDD.n2081 GND 0.00386f
C2612 VDD.n2082 GND 0.00386f
C2613 VDD.n2083 GND 0.00386f
C2614 VDD.n2084 GND 0.00386f
C2615 VDD.n2085 GND 0.00386f
C2616 VDD.n2087 GND 0.00386f
C2617 VDD.n2089 GND 0.00386f
C2618 VDD.n2090 GND 0.00386f
C2619 VDD.n2091 GND 0.00386f
C2620 VDD.n2092 GND 0.00386f
C2621 VDD.n2093 GND 0.00386f
C2622 VDD.n2095 GND 0.00386f
C2623 VDD.n2096 GND 0.00386f
C2624 VDD.n2097 GND 0.00386f
C2625 VDD.n2098 GND 0.00386f
C2626 VDD.n2099 GND 0.00386f
C2627 VDD.n2100 GND 0.00386f
C2628 VDD.n2102 GND 0.00386f
C2629 VDD.n2103 GND 0.00386f
C2630 VDD.n2104 GND 0.009516f
C2631 VDD.n2105 GND 0.009102f
C2632 VDD.n2106 GND 0.009102f
C2633 VDD.n2107 GND 0.380743f
C2634 VDD.n2108 GND 0.009102f
C2635 VDD.n2109 GND 0.009102f
C2636 VDD.n2110 GND 0.00386f
C2637 VDD.n2111 GND 0.00386f
C2638 VDD.n2112 GND 0.00386f
C2639 VDD.n2113 GND 0.262848f
C2640 VDD.n2114 GND 0.00386f
C2641 VDD.n2115 GND 0.00386f
C2642 VDD.n2116 GND 0.00386f
C2643 VDD.n2117 GND 0.00386f
C2644 VDD.n2118 GND 0.00386f
C2645 VDD.n2119 GND 0.206799f
C2646 VDD.n2120 GND 0.00386f
C2647 VDD.n2121 GND 0.00386f
C2648 VDD.n2122 GND 0.00386f
C2649 VDD.n2123 GND 0.00386f
C2650 VDD.n2124 GND 0.00386f
C2651 VDD.n2125 GND 0.19327f
C2652 VDD.n2126 GND 0.00386f
C2653 VDD.n2127 GND 0.00386f
C2654 VDD.n2128 GND 0.00386f
C2655 VDD.n2129 GND 0.00386f
C2656 VDD.n2130 GND 0.00386f
C2657 VDD.n2131 GND 0.262848f
C2658 VDD.n2132 GND 0.00386f
C2659 VDD.n2133 GND 0.00386f
C2660 VDD.n2134 GND 0.00386f
C2661 VDD.n2135 GND 0.00386f
C2662 VDD.n2136 GND 0.00386f
C2663 VDD.n2137 GND 0.262848f
C2664 VDD.n2138 GND 0.00386f
C2665 VDD.n2139 GND 0.00386f
C2666 VDD.n2140 GND 0.00386f
C2667 VDD.n2141 GND 0.00386f
C2668 VDD.n2142 GND 0.00386f
C2669 VDD.n2143 GND 0.262848f
C2670 VDD.n2144 GND 0.00386f
C2671 VDD.n2145 GND 0.00386f
C2672 VDD.n2146 GND 0.00386f
C2673 VDD.n2147 GND 0.00386f
C2674 VDD.n2148 GND 0.00386f
C2675 VDD.n2149 GND 0.262848f
C2676 VDD.n2150 GND 0.00386f
C2677 VDD.n2151 GND 0.00386f
C2678 VDD.n2152 GND 0.00386f
C2679 VDD.n2153 GND 0.00386f
C2680 VDD.n2154 GND 0.00386f
C2681 VDD.n2155 GND 0.199069f
C2682 VDD.n2156 GND 0.00386f
C2683 VDD.n2157 GND 0.00386f
C2684 VDD.n2158 GND 0.00386f
C2685 VDD.n2159 GND 0.00386f
C2686 VDD.n2160 GND 0.00386f
C2687 VDD.n2161 GND 0.262848f
C2688 VDD.n2162 GND 0.00386f
C2689 VDD.n2163 GND 0.00386f
C2690 VDD.n2164 GND 0.00386f
C2691 VDD.n2165 GND 0.00386f
C2692 VDD.n2166 GND 0.00386f
C2693 VDD.n2167 GND 0.208732f
C2694 VDD.n2168 GND 0.00386f
C2695 VDD.n2169 GND 0.00386f
C2696 VDD.n2170 GND 0.00386f
C2697 VDD.n2171 GND 0.00386f
C2698 VDD.n2172 GND 0.00386f
C2699 VDD.n2173 GND 0.262848f
C2700 VDD.n2174 GND 0.00386f
C2701 VDD.n2175 GND 0.00386f
C2702 VDD.n2176 GND 0.00386f
C2703 VDD.n2177 GND 0.00386f
C2704 VDD.n2178 GND 0.00386f
C2705 VDD.n2179 GND 0.262848f
C2706 VDD.n2180 GND 0.00386f
C2707 VDD.n2181 GND 0.00386f
C2708 VDD.n2182 GND 0.00386f
C2709 VDD.n2183 GND 0.00386f
C2710 VDD.n2184 GND 0.00386f
C2711 VDD.n2185 GND 0.183607f
C2712 VDD.n2186 GND 0.00386f
C2713 VDD.n2187 GND 0.00386f
C2714 VDD.n2188 GND 0.00386f
C2715 VDD.n2189 GND 0.00386f
C2716 VDD.n2190 GND 0.00386f
C2717 VDD.n2191 GND 0.262848f
C2718 VDD.n2192 GND 0.00386f
C2719 VDD.n2193 GND 0.00386f
C2720 VDD.n2194 GND 0.00386f
C2721 VDD.n2195 GND 0.00386f
C2722 VDD.n2196 GND 0.00386f
C2723 VDD.n2197 GND 0.262848f
C2724 VDD.n2198 GND 0.00386f
C2725 VDD.n2199 GND 0.00386f
C2726 VDD.n2200 GND 0.00386f
C2727 VDD.n2201 GND 0.00386f
C2728 VDD.n2202 GND 0.00386f
C2729 VDD.n2203 GND 0.197136f
C2730 VDD.n2204 GND 0.00386f
C2731 VDD.n2205 GND 0.00386f
C2732 VDD.n2206 GND 0.00386f
C2733 VDD.n2207 GND 0.00386f
C2734 VDD.n2208 GND 0.00386f
C2735 VDD.n2209 GND 0.262848f
C2736 VDD.n2210 GND 0.00386f
C2737 VDD.n2211 GND 0.00386f
C2738 VDD.n2212 GND 0.00386f
C2739 VDD.n2213 GND 0.00386f
C2740 VDD.n2214 GND 0.00386f
C2741 VDD.n2215 GND 0.262848f
C2742 VDD.n2216 GND 0.00386f
C2743 VDD.n2217 GND 0.00386f
C2744 VDD.n2218 GND 0.00386f
C2745 VDD.n2219 GND 0.00386f
C2746 VDD.n2220 GND 0.00386f
C2747 VDD.n2221 GND 0.222261f
C2748 VDD.n2222 GND 0.00386f
C2749 VDD.n2223 GND 0.00386f
C2750 VDD.n2224 GND 0.00386f
C2751 VDD.n2225 GND 0.00386f
C2752 VDD.n2226 GND 0.00386f
C2753 VDD.n2227 GND 0.262848f
C2754 VDD.n2228 GND 0.00386f
C2755 VDD.n2229 GND 0.00386f
C2756 VDD.n2230 GND 0.00386f
C2757 VDD.n2231 GND 0.00386f
C2758 VDD.n2232 GND 0.00386f
C2759 VDD.n2233 GND 0.18554f
C2760 VDD.n2234 GND 0.00386f
C2761 VDD.n2235 GND 0.00386f
C2762 VDD.n2236 GND 0.00386f
C2763 VDD.n2237 GND 0.00386f
C2764 VDD.n2238 GND 0.00386f
C2765 VDD.n2239 GND 0.262848f
C2766 VDD.n2240 GND 0.00386f
C2767 VDD.n2241 GND 0.00386f
C2768 VDD.n2242 GND 0.00386f
C2769 VDD.n2243 GND 0.00386f
C2770 VDD.n2244 GND 0.00386f
C2771 VDD.n2245 GND 0.262848f
C2772 VDD.n2246 GND 0.00386f
C2773 VDD.n2247 GND 0.00386f
C2774 VDD.n2248 GND 0.00386f
C2775 VDD.n2249 GND 0.00386f
C2776 VDD.n2250 GND 0.00386f
C2777 VDD.n2251 GND 0.262848f
C2778 VDD.n2252 GND 0.00386f
C2779 VDD.n2253 GND 0.00386f
C2780 VDD.n2254 GND 0.00386f
C2781 VDD.n2255 GND 0.00386f
C2782 VDD.n2256 GND 0.00386f
C2783 VDD.n2257 GND 0.262848f
C2784 VDD.n2258 GND 0.00386f
C2785 VDD.n2259 GND 0.00386f
C2786 VDD.n2260 GND 0.00386f
C2787 VDD.n2261 GND 0.00386f
C2788 VDD.n2262 GND 0.00386f
C2789 VDD.n2263 GND 0.262848f
C2790 VDD.n2264 GND 0.00386f
C2791 VDD.n2265 GND 0.00386f
C2792 VDD.n2266 GND 0.00386f
C2793 VDD.n2267 GND 0.00386f
C2794 VDD.n2268 GND 0.00386f
C2795 VDD.n2269 GND 0.156549f
C2796 VDD.n2270 GND 0.00386f
C2797 VDD.n2271 GND 0.00386f
C2798 VDD.n2272 GND 0.00386f
C2799 VDD.n2273 GND 0.00386f
C2800 VDD.n2274 GND 0.00386f
C2801 VDD.n2275 GND 0.201001f
C2802 VDD.n2276 GND 0.00386f
C2803 VDD.n2277 GND 0.00386f
C2804 VDD.n2278 GND 0.00386f
C2805 VDD.t55 GND 0.042906f
C2806 VDD.t54 GND 0.059398f
C2807 VDD.t52 GND 0.475789f
C2808 VDD.n2279 GND 0.099866f
C2809 VDD.n2280 GND 0.077301f
C2810 VDD.n2281 GND 0.005516f
C2811 VDD.n2282 GND 0.00386f
C2812 VDD.n2283 GND 0.002952f
C2813 VDD.n2284 GND 0.00386f
C2814 VDD.n2285 GND 0.00386f
C2815 VDD.n2286 GND 0.00386f
C2816 VDD.n2287 GND 0.00386f
C2817 VDD.n2288 GND 0.00386f
C2818 VDD.n2289 GND 0.00386f
C2819 VDD.n2290 GND 0.00386f
C2820 VDD.n2291 GND 0.00386f
C2821 VDD.n2292 GND 0.00386f
C2822 VDD.n2293 GND 0.00386f
C2823 VDD.n2294 GND 0.00386f
C2824 VDD.n2295 GND 0.00386f
C2825 VDD.n2296 GND 0.00386f
C2826 VDD.n2297 GND 0.00386f
C2827 VDD.n2298 GND 0.00386f
C2828 VDD.n2299 GND -0.500914f
C2829 VDD.n2300 GND -0.500914f
C2830 VDD.n2301 GND 0.00386f
C2831 VDD.n2302 GND 0.00386f
C2832 VDD.n2303 GND 0.00386f
C2833 VDD.n2304 GND 0.00386f
C2834 VDD.n2305 GND 0.00386f
C2835 VDD.n2306 GND 0.00386f
C2836 VDD.n2307 GND 0.00386f
C2837 VDD.n2308 GND 0.00386f
C2838 VDD.n2309 GND 0.00386f
C2839 VDD.n2310 GND 0.00386f
C2840 VDD.n2311 GND 0.00386f
C2841 VDD.n2312 GND 0.00386f
C2842 VDD.n2313 GND 0.00386f
C2843 VDD.n2314 GND 0.00386f
C2844 VDD.n2315 GND 0.00386f
C2845 VDD.n2316 GND 0.00386f
C2846 VDD.n2317 GND 0.00386f
C2847 VDD.n2318 GND 0.00386f
C2848 VDD.n2319 GND 0.00386f
C2849 VDD.n2320 GND 0.009516f
C2850 VDD.n2321 GND 0.009516f
C2851 VDD.n2322 GND 0.009102f
C2852 VDD.n2323 GND 0.009102f
C2853 VDD.n2324 GND 0.00386f
C2854 VDD.n2325 GND 0.00386f
C2855 VDD.n2326 GND 0.00386f
C2856 VDD.n2327 GND 0.00386f
C2857 VDD.n2328 GND 0.00386f
C2858 VDD.n2329 GND 0.00386f
C2859 VDD.n2330 GND 0.00386f
C2860 VDD.n2331 GND 0.262848f
C2861 VDD.n2332 GND 0.00386f
C2862 VDD.n2333 GND 0.00386f
C2863 VDD.n2334 GND 0.00386f
C2864 VDD.n2335 GND 0.00386f
C2865 VDD.n2336 GND 0.00386f
C2866 VDD.n2337 GND 0.262848f
C2867 VDD.n2338 GND 0.00386f
C2868 VDD.n2339 GND 0.00386f
C2869 VDD.n2340 GND 0.00386f
C2870 VDD.n2341 GND 0.00386f
C2871 VDD.n2342 GND 0.009538f
C2872 VDD.n2343 GND 0.009102f
C2873 VDD.n2344 GND 0.009516f
C2874 VDD.n2345 GND 0.009081f
C2875 VDD.n2346 GND 0.002838f
C2876 VDD.n2347 GND 0.00386f
C2877 VDD.n2348 GND 0.00386f
C2878 VDD.n2349 GND 0.002952f
C2879 VDD.n2350 GND 0.00386f
C2880 VDD.n2351 GND 0.00386f
C2881 VDD.n2352 GND 0.00386f
C2882 VDD.n2353 GND 0.00386f
C2883 VDD.n2354 GND 0.00386f
C2884 VDD.n2355 GND 0.00386f
C2885 VDD.n2356 GND 0.00386f
C2886 VDD.n2357 GND 0.00386f
C2887 VDD.n2358 GND 0.00386f
C2888 VDD.n2359 GND 0.00386f
C2889 VDD.n2360 GND 0.00386f
C2890 VDD.n2361 GND 0.00386f
C2891 VDD.n2362 GND 0.00386f
C2892 VDD.n2363 GND 0.00386f
C2893 VDD.n2364 GND 0.00386f
C2894 VDD.n2365 GND -0.495237f
C2895 VDD.n2366 GND -0.495237f
C2896 VDD.n2367 GND 0.00386f
C2897 VDD.n2368 GND 0.00386f
C2898 VDD.n2369 GND 0.00386f
C2899 VDD.n2370 GND 0.00386f
C2900 VDD.n2371 GND 0.00386f
C2901 VDD.n2372 GND 0.00386f
C2902 VDD.n2373 GND 0.00386f
C2903 VDD.n2374 GND 0.00386f
C2904 VDD.n2375 GND 0.00386f
C2905 VDD.n2376 GND 0.00386f
C2906 VDD.n2377 GND 0.00386f
C2907 VDD.n2378 GND 0.00386f
C2908 VDD.n2379 GND 0.00386f
C2909 VDD.n2380 GND 0.00386f
C2910 VDD.n2381 GND 0.00386f
C2911 VDD.n2382 GND 0.00386f
C2912 VDD.n2383 GND 0.00386f
C2913 VDD.n2384 GND 0.00386f
C2914 VDD.n2385 GND 0.00386f
C2915 VDD.n2386 GND 0.009516f
C2916 VDD.n2387 GND 0.009516f
C2917 VDD.n2388 GND 0.009102f
C2918 VDD.n2389 GND 0.00386f
C2919 VDD.n2390 GND 0.00386f
C2920 VDD.n2391 GND 0.262848f
C2921 VDD.n2392 GND 0.00386f
C2922 VDD.n2393 GND 0.00386f
C2923 VDD.n2394 GND 0.009538f
C2924 VDD.n2395 GND 0.009081f
C2925 VDD.n2396 GND 0.009516f
C2926 VDD.n2398 GND 1.43407f
C2927 VDD.t8 GND 2.84494f
C2928 VDD.t21 GND 3.28946f
C2929 VDD.t84 GND 4.2017f
C2930 VDD.n2408 GND 0.005676f
C2931 VDD.n2409 GND 0.005676f
C2932 VDD.n2410 GND 0.0128f
C2933 VDD.n2411 GND 0.005676f
C2934 VDD.n2412 GND 0.005676f
C2935 VDD.n2413 GND 0.005676f
C2936 VDD.n2414 GND 0.005676f
C2937 VDD.n2415 GND 0.005676f
C2938 VDD.n2416 GND 0.005676f
C2939 VDD.n2417 GND 0.005676f
C2940 VDD.n2418 GND 0.005676f
C2941 VDD.n2419 GND 0.005676f
C2942 VDD.t74 GND 0.049112f
C2943 VDD.t75 GND 0.063006f
C2944 VDD.t73 GND 0.385677f
C2945 VDD.n2420 GND 0.054096f
C2946 VDD.n2421 GND 0.037762f
C2947 VDD.n2422 GND 0.005676f
C2948 VDD.n2423 GND 0.005676f
C2949 VDD.n2424 GND 0.005676f
C2950 VDD.n2425 GND 0.005676f
C2951 VDD.n2426 GND 0.005676f
C2952 VDD.n2427 GND 0.005676f
C2953 VDD.n2428 GND 0.005676f
C2954 VDD.n2429 GND 0.005676f
C2955 VDD.n2430 GND 0.005676f
C2956 VDD.n2431 GND 0.005676f
C2957 VDD.n2432 GND 0.002467f
C2958 VDD.n2433 GND 0.004569f
C2959 VDD.n2434 GND 0.005676f
C2960 VDD.n2435 GND 0.005676f
C2961 VDD.n2436 GND 0.004569f
C2962 VDD.n2437 GND 0.004569f
C2963 VDD.n2438 GND 0.005676f
C2964 VDD.n2439 GND 0.005676f
C2965 VDD.n2440 GND 0.004569f
C2966 VDD.n2441 GND 0.004569f
C2967 VDD.n2442 GND 0.005676f
C2968 VDD.n2443 GND 0.005676f
C2969 VDD.n2444 GND 0.004569f
C2970 VDD.n2445 GND 0.004569f
C2971 VDD.n2446 GND 0.005676f
C2972 VDD.n2447 GND 0.005676f
C2973 VDD.n2448 GND 0.004569f
C2974 VDD.n2449 GND 0.004569f
C2975 VDD.n2450 GND 0.005676f
C2976 VDD.n2451 GND 0.005676f
C2977 VDD.n2452 GND 0.004158f
C2978 VDD.n2453 GND 0.00932f
C2979 VDD.n2454 GND 0.005676f
C2980 VDD.n2455 GND 0.005676f
C2981 VDD.n2456 GND 0.003472f
C2982 VDD.n2457 GND 0.004569f
C2983 VDD.n2458 GND 0.005676f
C2984 VDD.n2459 GND 0.005676f
C2985 VDD.n2460 GND 0.004569f
C2986 VDD.n2461 GND 0.004569f
C2987 VDD.n2462 GND 0.005676f
C2988 VDD.n2463 GND 0.005676f
C2989 VDD.n2464 GND 0.004569f
C2990 VDD.n2465 GND 0.005676f
C2991 VDD.n2466 GND 0.004569f
C2992 VDD.n2467 GND 0.004569f
C2993 VDD.n2468 GND 0.004569f
C2994 VDD.n2469 GND 0.003792f
C2995 VDD.n2470 GND 0.0128f
C2996 VDD.n2472 GND 2.64587f
C2997 VDD.n2473 GND 0.0128f
C2998 VDD.n2474 GND 0.002102f
C2999 VDD.n2475 GND 0.0128f
C3000 VDD.n2476 GND 0.0128f
C3001 VDD.n2477 GND 0.005676f
C3002 VDD.n2478 GND 0.004569f
C3003 VDD.n2479 GND 0.005676f
C3004 VDD.n2480 GND 0.386541f
C3005 VDD.n2481 GND 0.005676f
C3006 VDD.n2482 GND 0.004569f
C3007 VDD.n2483 GND 0.005676f
C3008 VDD.n2484 GND 0.005676f
C3009 VDD.n2485 GND 0.005676f
C3010 VDD.n2486 GND 0.004569f
C3011 VDD.n2487 GND 0.005676f
C3012 VDD.n2488 GND 0.386541f
C3013 VDD.n2489 GND 0.005676f
C3014 VDD.n2490 GND 0.004569f
C3015 VDD.n2491 GND 0.005676f
C3016 VDD.n2492 GND 0.005676f
C3017 VDD.n2493 GND 0.005676f
C3018 VDD.n2494 GND 0.004569f
C3019 VDD.n2495 GND 0.005676f
C3020 VDD.n2496 GND 0.239655f
C3021 VDD.n2497 GND 0.005676f
C3022 VDD.n2498 GND 0.004569f
C3023 VDD.n2499 GND 0.005676f
C3024 VDD.n2500 GND 0.005676f
C3025 VDD.n2501 GND 0.005676f
C3026 VDD.n2502 GND 0.004569f
C3027 VDD.n2503 GND 0.005676f
C3028 VDD.n2504 GND 0.386541f
C3029 VDD.n2505 GND 0.005676f
C3030 VDD.n2506 GND 0.004569f
C3031 VDD.n2507 GND 0.005676f
C3032 VDD.n2508 GND 0.005676f
C3033 VDD.n2509 GND 0.005676f
C3034 VDD.n2510 GND 0.004569f
C3035 VDD.n2511 GND 0.005676f
C3036 VDD.n2512 GND 0.386541f
C3037 VDD.n2513 GND 0.005676f
C3038 VDD.n2514 GND 0.004569f
C3039 VDD.n2515 GND 0.005676f
C3040 VDD.n2516 GND 0.005676f
C3041 VDD.n2517 GND 0.005676f
C3042 VDD.n2518 GND 0.004569f
C3043 VDD.n2519 GND 0.005676f
C3044 VDD.n2520 GND 0.386541f
C3045 VDD.n2521 GND 0.005676f
C3046 VDD.n2522 GND 0.004569f
C3047 VDD.n2523 GND 0.005676f
C3048 VDD.n2524 GND 0.005676f
C3049 VDD.n2525 GND 0.005676f
C3050 VDD.n2526 GND 0.004569f
C3051 VDD.n2527 GND 0.005676f
C3052 VDD.n2528 GND 0.386541f
C3053 VDD.n2529 GND 0.005676f
C3054 VDD.n2530 GND 0.004569f
C3055 VDD.n2531 GND 0.005676f
C3056 VDD.n2532 GND 0.005676f
C3057 VDD.n2533 GND 0.005676f
C3058 VDD.n2534 GND 0.004569f
C3059 VDD.n2535 GND 0.005676f
C3060 VDD.n2536 GND 0.332425f
C3061 VDD.n2537 GND 0.005676f
C3062 VDD.n2538 GND 0.004569f
C3063 VDD.n2539 GND 0.005676f
C3064 VDD.n2540 GND 0.005676f
C3065 VDD.n2541 GND 0.005676f
C3066 VDD.n2542 GND 0.004569f
C3067 VDD.n2543 GND 0.005676f
C3068 VDD.n2544 GND 0.386541f
C3069 VDD.n2545 GND 0.005676f
C3070 VDD.n2546 GND 0.004569f
C3071 VDD.n2547 GND 0.005676f
C3072 VDD.n2548 GND 0.005676f
C3073 VDD.n2549 GND 0.005676f
C3074 VDD.n2550 GND 0.004569f
C3075 VDD.n2551 GND 0.005676f
C3076 VDD.n2552 GND 0.386541f
C3077 VDD.n2553 GND 0.005676f
C3078 VDD.n2554 GND 0.004569f
C3079 VDD.n2555 GND 0.005676f
C3080 VDD.n2556 GND 0.005676f
C3081 VDD.n2557 GND 0.005676f
C3082 VDD.n2558 GND 0.005676f
C3083 VDD.n2559 GND 0.005676f
C3084 VDD.n2560 GND 0.004569f
C3085 VDD.n2561 GND 0.004569f
C3086 VDD.n2562 GND 0.005676f
C3087 VDD.n2563 GND 0.386541f
C3088 VDD.n2564 GND 0.005676f
C3089 VDD.n2565 GND 0.004569f
C3090 VDD.n2566 GND 0.005676f
C3091 VDD.n2567 GND 0.005676f
C3092 VDD.n2568 GND 0.005676f
C3093 VDD.n2569 GND 0.004569f
C3094 VDD.n2570 GND 0.005676f
C3095 VDD.n2571 GND 0.386541f
C3096 VDD.n2572 GND 0.289906f
C3097 VDD.n2573 GND 0.005676f
C3098 VDD.n2574 GND 0.004569f
C3099 VDD.n2575 GND 0.004569f
C3100 VDD.n2576 GND 0.005676f
C3101 VDD.n2577 GND 0.005676f
C3102 VDD.n2578 GND 0.005676f
C3103 VDD.n2579 GND 0.004569f
C3104 VDD.n2580 GND 0.005676f
C3105 VDD.n2581 GND 0.004569f
C3106 VDD.n2582 GND 0.004569f
C3107 VDD.n2583 GND 0.005676f
C3108 VDD.n2584 GND 0.005676f
C3109 VDD.n2585 GND 0.005676f
C3110 VDD.n2586 GND 0.004569f
C3111 VDD.n2587 GND 0.005676f
C3112 VDD.n2588 GND 0.004569f
C3113 VDD.n2589 GND 0.004569f
C3114 VDD.n2590 GND 0.005676f
C3115 VDD.n2591 GND 0.005676f
C3116 VDD.n2592 GND 0.005676f
C3117 VDD.n2593 GND 0.004569f
C3118 VDD.n2594 GND 0.005676f
C3119 VDD.n2595 GND 0.004569f
C3120 VDD.n2596 GND 0.004569f
C3121 VDD.n2597 GND 0.005676f
C3122 VDD.n2598 GND 0.005676f
C3123 VDD.n2599 GND 0.005676f
C3124 VDD.n2600 GND 0.004569f
C3125 VDD.n2601 GND 0.005676f
C3126 VDD.n2602 GND 0.004569f
C3127 VDD.n2603 GND 0.004569f
C3128 VDD.n2604 GND 0.005676f
C3129 VDD.n2605 GND 0.005676f
C3130 VDD.n2606 GND 0.005676f
C3131 VDD.n2607 GND 0.004569f
C3132 VDD.n2608 GND 0.005676f
C3133 VDD.n2609 GND 0.004569f
C3134 VDD.n2610 GND 0.004569f
C3135 VDD.n2611 GND 0.005676f
C3136 VDD.n2612 GND 0.005676f
C3137 VDD.n2613 GND 0.005676f
C3138 VDD.n2614 GND 0.004569f
C3139 VDD.n2615 GND 0.005676f
C3140 VDD.n2616 GND 0.004569f
C3141 VDD.n2617 GND 0.003792f
C3142 VDD.n2618 GND 0.0128f
C3143 VDD.n2619 GND 0.0128f
C3144 VDD.n2620 GND 0.002102f
C3145 VDD.n2621 GND 0.0128f
C3146 VDD.n2623 GND 0.836861f
C3147 VDD.n2624 GND 0.49284f
C3148 VDD.n2625 GND 0.0128f
C3149 VDD.n2626 GND 0.003792f
C3150 VDD.n2627 GND 0.004569f
C3151 VDD.n2628 GND 0.004569f
C3152 VDD.n2629 GND 0.005676f
C3153 VDD.n2630 GND 0.386541f
C3154 VDD.n2631 GND 0.386541f
C3155 VDD.n2632 GND 0.340156f
C3156 VDD.n2633 GND 0.005676f
C3157 VDD.n2634 GND 0.004569f
C3158 VDD.n2635 GND 0.004569f
C3159 VDD.n2636 GND 0.004569f
C3160 VDD.n2637 GND 0.005676f
C3161 VDD.n2638 GND 0.386541f
C3162 VDD.n2639 GND 0.386541f
C3163 VDD.n2640 GND 0.386541f
C3164 VDD.n2641 GND 0.005676f
C3165 VDD.n2642 GND 0.004569f
C3166 VDD.n2643 GND 0.004569f
C3167 VDD.n2644 GND 0.004569f
C3168 VDD.n2645 GND 0.005676f
C3169 VDD.n2646 GND 0.386541f
C3170 VDD.n2647 GND 0.386541f
C3171 VDD.n2648 GND 0.386541f
C3172 VDD.n2649 GND 0.005676f
C3173 VDD.n2650 GND 0.004569f
C3174 VDD.n2651 GND 0.004569f
C3175 VDD.n2652 GND 0.004569f
C3176 VDD.n2653 GND 0.005676f
C3177 VDD.n2654 GND 0.386541f
C3178 VDD.n2655 GND 0.332425f
C3179 VDD.t96 GND 0.19327f
C3180 VDD.n2656 GND 0.247386f
C3181 VDD.n2657 GND 0.005676f
C3182 VDD.n2658 GND 0.004569f
C3183 VDD.n2659 GND 0.004569f
C3184 VDD.n2660 GND 0.004569f
C3185 VDD.n2661 GND 0.005676f
C3186 VDD.n2662 GND 0.386541f
C3187 VDD.n2663 GND 0.386541f
C3188 VDD.n2664 GND 0.386541f
C3189 VDD.n2665 GND 0.005676f
C3190 VDD.n2666 GND 0.004569f
C3191 VDD.n2667 GND 0.004569f
C3192 VDD.n2668 GND 0.004569f
C3193 VDD.n2669 GND 0.005676f
C3194 VDD.n2670 GND 0.386541f
C3195 VDD.n2671 GND 0.386541f
C3196 VDD.n2672 GND 0.289906f
C3197 VDD.n2673 GND 0.005676f
C3198 VDD.n2674 GND 0.004569f
C3199 VDD.n2675 GND 0.004363f
C3200 VDD.n2676 GND 0.545011f
C3201 VDD.n2677 GND 2.20764f
C3202 a_n12440_8296.n0 GND 0.376134f
C3203 a_n12440_8296.n1 GND 0.015927f
C3204 a_n12440_8296.n2 GND 0.376134f
C3205 a_n12440_8296.n3 GND 0.015927f
C3206 a_n12440_8296.n4 GND 0.672412f
C3207 a_n12440_8296.n5 GND 0.245381f
C3208 a_n12440_8296.n6 GND 0.672412f
C3209 a_n12440_8296.n7 GND 0.245381f
C3210 a_n12440_8296.n8 GND 0.672411f
C3211 a_n12440_8296.n9 GND 0.245381f
C3212 a_n12440_8296.n10 GND 0.672411f
C3213 a_n12440_8296.n11 GND 0.245381f
C3214 a_n12440_8296.n12 GND 0.376476f
C3215 a_n12440_8296.n13 GND 0.60529f
C3216 a_n12440_8296.n14 GND 0.423468f
C3217 a_n12440_8296.n15 GND 0.60529f
C3218 a_n12440_8296.n16 GND 0.376476f
C3219 a_n12440_8296.n17 GND 0.60529f
C3220 a_n12440_8296.n18 GND 0.423468f
C3221 a_n12440_8296.n19 GND 0.60529f
C3222 a_n12440_8296.n20 GND 0.013714f
C3223 a_n12440_8296.n21 GND 0.019351f
C3224 a_n12440_8296.n22 GND 0.060563f
C3225 a_n12440_8296.n23 GND 0.013714f
C3226 a_n12440_8296.n24 GND 0.019351f
C3227 a_n12440_8296.n25 GND 0.060563f
C3228 a_n12440_8296.t5 GND 0.044937f
C3229 a_n12440_8296.t3 GND 0.044937f
C3230 a_n12440_8296.t9 GND 0.044937f
C3231 a_n12440_8296.n26 GND 0.363592f
C3232 a_n12440_8296.t6 GND 0.044937f
C3233 a_n12440_8296.t7 GND 0.044937f
C3234 a_n12440_8296.n27 GND 0.363592f
C3235 a_n12440_8296.n28 GND 2.32233f
C3236 a_n12440_8296.t4 GND 0.044937f
C3237 a_n12440_8296.t8 GND 0.044937f
C3238 a_n12440_8296.n29 GND 0.352255f
C3239 a_n12440_8296.n30 GND 1.83727f
C3240 a_n12440_8296.t12 GND 0.060409f
C3241 a_n12440_8296.t2 GND 0.060409f
C3242 a_n12440_8296.n31 GND 0.403317f
C3243 a_n12440_8296.n32 GND 0.015697f
C3244 a_n12440_8296.n33 GND 0.007736f
C3245 a_n12440_8296.n34 GND 0.018285f
C3246 a_n12440_8296.n35 GND 0.008191f
C3247 a_n12440_8296.t13 GND 0.039847f
C3248 a_n12440_8296.n36 GND 0.018285f
C3249 a_n12440_8296.n37 GND 0.018285f
C3250 a_n12440_8296.n38 GND 0.008191f
C3251 a_n12440_8296.n39 GND 0.007736f
C3252 a_n12440_8296.n40 GND 0.007736f
C3253 a_n12440_8296.n41 GND 0.008191f
C3254 a_n12440_8296.n42 GND 0.018285f
C3255 a_n12440_8296.n43 GND 0.043853f
C3256 a_n12440_8296.n44 GND 0.008191f
C3257 a_n12440_8296.n45 GND 0.007736f
C3258 a_n12440_8296.n46 GND 0.031989f
C3259 a_n12440_8296.n47 GND 2.70253f
C3260 a_n12440_8296.n48 GND 0.015697f
C3261 a_n12440_8296.n49 GND 0.007736f
C3262 a_n12440_8296.n50 GND 0.018285f
C3263 a_n12440_8296.n51 GND 0.008191f
C3264 a_n12440_8296.t1 GND 0.039847f
C3265 a_n12440_8296.n52 GND 0.018285f
C3266 a_n12440_8296.n53 GND 0.018285f
C3267 a_n12440_8296.n54 GND 0.008191f
C3268 a_n12440_8296.n55 GND 0.007736f
C3269 a_n12440_8296.n56 GND 0.007736f
C3270 a_n12440_8296.n57 GND 0.008191f
C3271 a_n12440_8296.n58 GND 0.018285f
C3272 a_n12440_8296.n59 GND 0.043853f
C3273 a_n12440_8296.n60 GND 0.008191f
C3274 a_n12440_8296.n61 GND 0.007736f
C3275 a_n12440_8296.n62 GND 0.042707f
C3276 a_n12440_8296.t0 GND 0.060409f
C3277 a_n12440_8296.t11 GND 0.060409f
C3278 a_n12440_8296.n63 GND 0.386639f
C3279 a_n12440_8296.n64 GND 1.84563f
C3280 a_n12440_8296.n65 GND 3.91069f
C3281 a_n12440_8296.t14 GND 1.5895f
C3282 a_n12440_8296.t18 GND 1.84573f
C3283 a_n12440_8296.n66 GND 0.716388f
C3284 a_n12440_8296.t17 GND 1.33806f
C3285 a_n12440_8296.n67 GND 0.776163f
C3286 a_n12440_8296.t19 GND 1.5895f
C3287 a_n12440_8296.t23 GND 1.84573f
C3288 a_n12440_8296.n68 GND 0.716388f
C3289 a_n12440_8296.t22 GND 1.33806f
C3290 a_n12440_8296.n69 GND 0.776163f
C3291 a_n12440_8296.n70 GND 2.04842f
C3292 a_n12440_8296.t24 GND 1.5895f
C3293 a_n12440_8296.t16 GND 1.84573f
C3294 a_n12440_8296.n71 GND 0.716391f
C3295 a_n12440_8296.t15 GND 1.33806f
C3296 a_n12440_8296.n72 GND 0.776163f
C3297 a_n12440_8296.t25 GND 1.5895f
C3298 a_n12440_8296.t20 GND 1.84573f
C3299 a_n12440_8296.n73 GND 0.716391f
C3300 a_n12440_8296.t21 GND 1.33806f
C3301 a_n12440_8296.n74 GND 0.776163f
C3302 a_n12440_8296.n75 GND 1.34918f
C3303 a_n12440_8296.n76 GND 18.874699f
C3304 a_n12440_8296.n77 GND 3.04405f
C3305 a_n12440_8296.n78 GND 0.856809f
C3306 a_n12440_8296.n79 GND 0.363696f
C3307 a_n12440_8296.t10 GND 0.044937f
C3308 a_n4178_n267.n0 GND 0.011838f
C3309 a_n4178_n267.n1 GND 0.050457f
C3310 a_n4178_n267.n2 GND 0.011838f
C3311 a_n4178_n267.n3 GND 0.050457f
C3312 a_n4178_n267.n4 GND 0.011838f
C3313 a_n4178_n267.n5 GND 0.050457f
C3314 a_n4178_n267.n6 GND 0.011838f
C3315 a_n4178_n267.n7 GND 0.050457f
C3316 a_n4178_n267.n8 GND 0.011838f
C3317 a_n4178_n267.n9 GND 0.050457f
C3318 a_n4178_n267.n10 GND 0.011838f
C3319 a_n4178_n267.n11 GND 0.050457f
C3320 a_n4178_n267.n12 GND 0.011838f
C3321 a_n4178_n267.n13 GND 0.050457f
C3322 a_n4178_n267.n14 GND 0.011838f
C3323 a_n4178_n267.n15 GND 0.050457f
C3324 a_n4178_n267.n16 GND 3.64649f
C3325 a_n4178_n267.n17 GND 0.47738f
C3326 a_n4178_n267.n18 GND 0.023448f
C3327 a_n4178_n267.n19 GND 0.47738f
C3328 a_n4178_n267.n20 GND 0.023448f
C3329 a_n4178_n267.n21 GND 0.47738f
C3330 a_n4178_n267.n22 GND 0.023448f
C3331 a_n4178_n267.n23 GND 0.47738f
C3332 a_n4178_n267.n24 GND 0.023448f
C3333 a_n4178_n267.n25 GND 0.47738f
C3334 a_n4178_n267.n26 GND 0.023448f
C3335 a_n4178_n267.n27 GND 0.47738f
C3336 a_n4178_n267.n28 GND 0.023448f
C3337 a_n4178_n267.n29 GND 0.47738f
C3338 a_n4178_n267.n30 GND 0.023448f
C3339 a_n4178_n267.n31 GND 0.47738f
C3340 a_n4178_n267.n32 GND 0.023448f
C3341 a_n4178_n267.n33 GND 0.026804f
C3342 a_n4178_n267.n34 GND 0.026804f
C3343 a_n4178_n267.n35 GND 0.026804f
C3344 a_n4178_n267.n36 GND 0.026804f
C3345 a_n4178_n267.n37 GND 0.026804f
C3346 a_n4178_n267.n38 GND 0.026804f
C3347 a_n4178_n267.n39 GND 0.026804f
C3348 a_n4178_n267.n40 GND 0.026804f
C3349 a_n4178_n267.n41 GND 0.02692f
C3350 a_n4178_n267.n42 GND 0.023448f
C3351 a_n4178_n267.n43 GND 0.02692f
C3352 a_n4178_n267.n44 GND 0.023448f
C3353 a_n4178_n267.n45 GND 0.02692f
C3354 a_n4178_n267.n46 GND 0.023448f
C3355 a_n4178_n267.n47 GND 0.02692f
C3356 a_n4178_n267.n48 GND 0.023448f
C3357 a_n4178_n267.n49 GND 0.02692f
C3358 a_n4178_n267.n50 GND 0.023448f
C3359 a_n4178_n267.n51 GND 0.02692f
C3360 a_n4178_n267.n52 GND 0.023448f
C3361 a_n4178_n267.n53 GND 0.02692f
C3362 a_n4178_n267.n54 GND 0.023448f
C3363 a_n4178_n267.n55 GND 0.02692f
C3364 a_n4178_n267.n56 GND 0.023448f
C3365 a_n4178_n267.n57 GND 0.773826f
C3366 a_n4178_n267.n58 GND 0.696263f
C3367 a_n4178_n267.n59 GND 0.773829f
C3368 a_n4178_n267.n60 GND 0.696263f
C3369 a_n4178_n267.t12 GND 1.02055f
C3370 a_n4178_n267.t10 GND 0.045961f
C3371 a_n4178_n267.n61 GND 0.020619f
C3372 a_n4178_n267.n62 GND 0.05672f
C3373 a_n4178_n267.n63 GND 0.051563f
C3374 a_n4178_n267.n64 GND 0.85313f
C3375 a_n4178_n267.t3 GND 0.066158f
C3376 a_n4178_n267.t6 GND 0.066158f
C3377 a_n4178_n267.n65 GND 0.473088f
C3378 a_n4178_n267.t7 GND 0.045961f
C3379 a_n4178_n267.n66 GND 0.020619f
C3380 a_n4178_n267.n67 GND 0.05672f
C3381 a_n4178_n267.n68 GND 0.051563f
C3382 a_n4178_n267.t13 GND 0.045961f
C3383 a_n4178_n267.n69 GND 0.020619f
C3384 a_n4178_n267.n70 GND 0.05672f
C3385 a_n4178_n267.n71 GND 0.051563f
C3386 a_n4178_n267.t17 GND 0.066158f
C3387 a_n4178_n267.t14 GND 0.066158f
C3388 a_n4178_n267.n72 GND 0.473088f
C3389 a_n4178_n267.n73 GND 0.773826f
C3390 a_n4178_n267.t2 GND 0.045961f
C3391 a_n4178_n267.n74 GND 0.020619f
C3392 a_n4178_n267.n75 GND 0.05672f
C3393 a_n4178_n267.n76 GND 0.051563f
C3394 a_n4178_n267.n77 GND 0.85313f
C3395 a_n4178_n267.n78 GND 1.79392f
C3396 a_n4178_n267.t4 GND 0.045961f
C3397 a_n4178_n267.n79 GND 0.020619f
C3398 a_n4178_n267.n80 GND 0.05672f
C3399 a_n4178_n267.n81 GND 0.051563f
C3400 a_n4178_n267.n82 GND 0.655045f
C3401 a_n4178_n267.t8 GND 0.066158f
C3402 a_n4178_n267.t9 GND 0.066158f
C3403 a_n4178_n267.n83 GND 0.473085f
C3404 a_n4178_n267.t5 GND 0.045961f
C3405 a_n4178_n267.n84 GND 0.020619f
C3406 a_n4178_n267.n85 GND 0.05672f
C3407 a_n4178_n267.n86 GND 0.051563f
C3408 a_n4178_n267.t0 GND 0.045961f
C3409 a_n4178_n267.n87 GND 0.020619f
C3410 a_n4178_n267.n88 GND 0.05672f
C3411 a_n4178_n267.n89 GND 0.051563f
C3412 a_n4178_n267.t15 GND 0.066158f
C3413 a_n4178_n267.t1 GND 0.066158f
C3414 a_n4178_n267.n90 GND 0.473085f
C3415 a_n4178_n267.n91 GND 0.773829f
C3416 a_n4178_n267.t16 GND 0.045961f
C3417 a_n4178_n267.n92 GND 0.020619f
C3418 a_n4178_n267.n93 GND 0.05672f
C3419 a_n4178_n267.n94 GND 0.051563f
C3420 a_n4178_n267.n95 GND 0.655045f
C3421 a_n4178_n267.n96 GND 2.0714f
C3422 a_n4178_n267.t11 GND 1.02055f
C3423 VN.n0 GND 0.024812f
C3424 VN.t9 GND 0.628387f
C3425 VN.n1 GND 0.024585f
C3426 VN.n2 GND 0.013191f
C3427 VN.n3 GND 0.026532f
C3428 VN.n4 GND 0.013191f
C3429 VN.t3 GND 0.628387f
C3430 VN.n5 GND 0.240904f
C3431 VN.n6 GND 0.013191f
C3432 VN.n7 GND 0.024585f
C3433 VN.n8 GND 0.013191f
C3434 VN.n9 GND 0.024585f
C3435 VN.n10 GND 0.013191f
C3436 VN.t6 GND 0.628387f
C3437 VN.n11 GND 0.287057f
C3438 VN.t5 GND 0.845751f
C3439 VN.n12 GND 0.318479f
C3440 VN.n13 GND 0.187201f
C3441 VN.n14 GND 0.012811f
C3442 VN.n15 GND 0.024585f
C3443 VN.n16 GND 0.024585f
C3444 VN.n17 GND 0.013191f
C3445 VN.n18 GND 0.013191f
C3446 VN.n19 GND 0.013191f
C3447 VN.n20 GND 0.026217f
C3448 VN.n21 GND 0.010664f
C3449 VN.n22 GND 0.026217f
C3450 VN.n23 GND 0.013191f
C3451 VN.n24 GND 0.013191f
C3452 VN.n25 GND 0.013191f
C3453 VN.n26 GND 0.024585f
C3454 VN.n27 GND 0.024585f
C3455 VN.n28 GND 0.012811f
C3456 VN.n29 GND 0.013191f
C3457 VN.n30 GND 0.013191f
C3458 VN.n31 GND 0.02422f
C3459 VN.n32 GND 0.024585f
C3460 VN.n33 GND 0.024585f
C3461 VN.n34 GND 0.013191f
C3462 VN.n35 GND 0.013191f
C3463 VN.n36 GND 0.013191f
C3464 VN.n37 GND 0.010817f
C3465 VN.n38 GND 0.025749f
C3466 VN.n39 GND 0.024585f
C3467 VN.n40 GND 0.013191f
C3468 VN.n41 GND 0.013191f
C3469 VN.n42 GND 0.013191f
C3470 VN.n43 GND 0.024585f
C3471 VN.n44 GND 0.013539f
C3472 VN.n45 GND 0.292089f
C3473 VN.n46 GND 0.248862f
C3474 VN.n47 GND 0.024812f
C3475 VN.t4 GND 0.628387f
C3476 VN.n48 GND 0.024585f
C3477 VN.n49 GND 0.013191f
C3478 VN.n50 GND 0.026532f
C3479 VN.n51 GND 0.013191f
C3480 VN.t8 GND 0.628387f
C3481 VN.n52 GND 0.240904f
C3482 VN.n53 GND 0.013191f
C3483 VN.n54 GND 0.024585f
C3484 VN.n55 GND 0.013191f
C3485 VN.n56 GND 0.024585f
C3486 VN.n57 GND 0.013191f
C3487 VN.t2 GND 0.628387f
C3488 VN.n58 GND 0.287057f
C3489 VN.t7 GND 0.845752f
C3490 VN.n59 GND 0.318479f
C3491 VN.n60 GND 0.187201f
C3492 VN.n61 GND 0.012811f
C3493 VN.n62 GND 0.024585f
C3494 VN.n63 GND 0.024585f
C3495 VN.n64 GND 0.013191f
C3496 VN.n65 GND 0.013191f
C3497 VN.n66 GND 0.013191f
C3498 VN.n67 GND 0.026217f
C3499 VN.n68 GND 0.010664f
C3500 VN.n69 GND 0.026217f
C3501 VN.n70 GND 0.013191f
C3502 VN.n71 GND 0.013191f
C3503 VN.n72 GND 0.013191f
C3504 VN.n73 GND 0.024585f
C3505 VN.n74 GND 0.024585f
C3506 VN.n75 GND 0.012811f
C3507 VN.n76 GND 0.013191f
C3508 VN.n77 GND 0.013191f
C3509 VN.n78 GND 0.02422f
C3510 VN.n79 GND 0.024585f
C3511 VN.n80 GND 0.024585f
C3512 VN.n81 GND 0.013191f
C3513 VN.n82 GND 0.013191f
C3514 VN.n83 GND 0.013191f
C3515 VN.n84 GND 0.010817f
C3516 VN.n85 GND 0.025749f
C3517 VN.n86 GND 0.024585f
C3518 VN.n87 GND 0.013191f
C3519 VN.n88 GND 0.013191f
C3520 VN.n89 GND 0.013191f
C3521 VN.n90 GND 0.024585f
C3522 VN.n91 GND 0.013539f
C3523 VN.n92 GND 0.292089f
C3524 VN.n93 GND 0.694845f
C3525 VN.n94 GND 0.848319f
C3526 VN.t0 GND 0.022772f
C3527 VN.t1 GND 0.022633f
C3528 VN.n95 GND 0.115623f
C3529 VN.n96 GND 3.14509f
C3530 a_n1431_n2782.t1 GND 1.5024f
C3531 a_n1431_n2782.t0 GND 1.4976f
C3532 DIFFPAIR_BIAS.t4 GND 0.545867f
C3533 DIFFPAIR_BIAS.t3 GND 0.194763f
C3534 DIFFPAIR_BIAS.t1 GND 0.190663f
C3535 DIFFPAIR_BIAS.n0 GND 0.408224f
C3536 DIFFPAIR_BIAS.t0 GND 0.519981f
C3537 DIFFPAIR_BIAS.t2 GND 0.525533f
C3538 DIFFPAIR_BIAS.n1 GND 0.638796f
C3539 DIFFPAIR_BIAS.n2 GND 0.638922f
C3540 DIFFPAIR_BIAS.t5 GND 0.545104f
C3541 DIFFPAIR_BIAS.n3 GND 0.285543f
C3542 DIFFPAIR_BIAS.n4 GND 0.477606f
C3543 VOUT.t5 GND 0.016083f
C3544 VOUT.t7 GND 0.016083f
C3545 VOUT.n0 GND 0.096637f
C3546 VOUT.t1 GND 0.12541f
C3547 VOUT.n1 GND 0.42632f
C3548 VOUT.t0 GND 0.016083f
C3549 VOUT.t9 GND 0.016083f
C3550 VOUT.n2 GND 0.096637f
C3551 VOUT.t3 GND 0.12541f
C3552 VOUT.n3 GND 0.408532f
C3553 VOUT.n4 GND 0.285299f
C3554 VOUT.n5 GND 8.423151f
C3555 VOUT.t44 GND 17.0612f
C3556 VOUT.t45 GND 10.529f
C3557 VOUT.n6 GND 11.1799f
C3558 VOUT.n7 GND 1.88444f
C3559 VOUT.t10 GND 0.129911f
C3560 VOUT.t6 GND 0.016083f
C3561 VOUT.t8 GND 0.016083f
C3562 VOUT.n8 GND 0.089912f
C3563 VOUT.n9 GND 0.410949f
C3564 VOUT.t4 GND 0.129911f
C3565 VOUT.t43 GND 0.016083f
C3566 VOUT.t2 GND 0.016083f
C3567 VOUT.n10 GND 0.089912f
C3568 VOUT.n11 GND 0.391912f
C3569 VOUT.n12 GND 0.321738f
C3570 VOUT.n13 GND 10.3756f
C3571 VOUT.t23 GND 0.015398f
C3572 VOUT.t26 GND 0.015398f
C3573 VOUT.n14 GND 0.128572f
C3574 VOUT.t36 GND 0.015398f
C3575 VOUT.t16 GND 0.015398f
C3576 VOUT.n15 GND 0.114245f
C3577 VOUT.n16 GND 0.453287f
C3578 VOUT.t28 GND 0.015398f
C3579 VOUT.t40 GND 0.015398f
C3580 VOUT.n17 GND 0.114245f
C3581 VOUT.n18 GND 0.232642f
C3582 VOUT.t20 GND 0.015398f
C3583 VOUT.t22 GND 0.015398f
C3584 VOUT.n19 GND 0.114245f
C3585 VOUT.n20 GND 0.262655f
C3586 VOUT.t39 GND 0.015398f
C3587 VOUT.t30 GND 0.015398f
C3588 VOUT.n21 GND 0.128572f
C3589 VOUT.t15 GND 0.015398f
C3590 VOUT.t41 GND 0.015398f
C3591 VOUT.n22 GND 0.114245f
C3592 VOUT.n23 GND 0.453287f
C3593 VOUT.t25 GND 0.015398f
C3594 VOUT.t17 GND 0.015398f
C3595 VOUT.n24 GND 0.114245f
C3596 VOUT.n25 GND 0.232642f
C3597 VOUT.t34 GND 0.015398f
C3598 VOUT.t27 GND 0.015398f
C3599 VOUT.n26 GND 0.114245f
C3600 VOUT.n27 GND 0.243567f
C3601 VOUT.n28 GND 0.328428f
C3602 VOUT.n29 GND 10.9936f
C3603 VOUT.t12 GND 0.015398f
C3604 VOUT.t38 GND 0.015398f
C3605 VOUT.n30 GND 0.128572f
C3606 VOUT.t29 GND 0.015398f
C3607 VOUT.t18 GND 0.015398f
C3608 VOUT.n31 GND 0.114245f
C3609 VOUT.n32 GND 0.453287f
C3610 VOUT.t21 GND 0.015398f
C3611 VOUT.t42 GND 0.015398f
C3612 VOUT.n33 GND 0.114245f
C3613 VOUT.n34 GND 0.232642f
C3614 VOUT.t13 GND 0.015398f
C3615 VOUT.t31 GND 0.015398f
C3616 VOUT.n35 GND 0.114245f
C3617 VOUT.n36 GND 0.262655f
C3618 VOUT.t37 GND 0.015398f
C3619 VOUT.t14 GND 0.015398f
C3620 VOUT.n37 GND 0.128572f
C3621 VOUT.t24 GND 0.015398f
C3622 VOUT.t32 GND 0.015398f
C3623 VOUT.n38 GND 0.114245f
C3624 VOUT.n39 GND 0.453287f
C3625 VOUT.t33 GND 0.015398f
C3626 VOUT.t11 GND 0.015398f
C3627 VOUT.n40 GND 0.114245f
C3628 VOUT.n41 GND 0.232642f
C3629 VOUT.t35 GND 0.015398f
C3630 VOUT.t19 GND 0.015398f
C3631 VOUT.n42 GND 0.114245f
C3632 VOUT.n43 GND 0.243567f
C3633 VOUT.n44 GND 0.328428f
C3634 VOUT.n45 GND 8.16125f
C3635 VOUT.n46 GND 4.8739f
C3636 CS_BIAS.t51 GND 0.19437f
C3637 CS_BIAS.n0 GND 0.093799f
C3638 CS_BIAS.n1 GND 0.004191f
C3639 CS_BIAS.n2 GND 0.007811f
C3640 CS_BIAS.n3 GND 0.004191f
C3641 CS_BIAS.n4 GND 0.007811f
C3642 CS_BIAS.n5 GND 0.004191f
C3643 CS_BIAS.n6 GND 0.00434f
C3644 CS_BIAS.n7 GND 0.004191f
C3645 CS_BIAS.t48 GND 0.19437f
C3646 CS_BIAS.n8 GND 0.075758f
C3647 CS_BIAS.n9 GND 0.007811f
C3648 CS_BIAS.n10 GND 0.004191f
C3649 CS_BIAS.n11 GND 0.007811f
C3650 CS_BIAS.n12 GND 0.004191f
C3651 CS_BIAS.t38 GND 0.19437f
C3652 CS_BIAS.n13 GND 0.075758f
C3653 CS_BIAS.n14 GND 0.004191f
C3654 CS_BIAS.n15 GND 0.007811f
C3655 CS_BIAS.n16 GND 0.004191f
C3656 CS_BIAS.n17 GND 0.007811f
C3657 CS_BIAS.n18 GND 0.004191f
C3658 CS_BIAS.n19 GND 0.004803f
C3659 CS_BIAS.n20 GND 0.004191f
C3660 CS_BIAS.t58 GND 0.19437f
C3661 CS_BIAS.n21 GND 0.075758f
C3662 CS_BIAS.n22 GND 0.007811f
C3663 CS_BIAS.t20 GND 0.19437f
C3664 CS_BIAS.n23 GND 0.093799f
C3665 CS_BIAS.n24 GND 0.004191f
C3666 CS_BIAS.n25 GND 0.007811f
C3667 CS_BIAS.n26 GND 0.004191f
C3668 CS_BIAS.n27 GND 0.007811f
C3669 CS_BIAS.n28 GND 0.004191f
C3670 CS_BIAS.n29 GND 0.00434f
C3671 CS_BIAS.n30 GND 0.004191f
C3672 CS_BIAS.t14 GND 0.19437f
C3673 CS_BIAS.n31 GND 0.075758f
C3674 CS_BIAS.n32 GND 0.007811f
C3675 CS_BIAS.n33 GND 0.004191f
C3676 CS_BIAS.n34 GND 0.007811f
C3677 CS_BIAS.n35 GND 0.004191f
C3678 CS_BIAS.t16 GND 0.19437f
C3679 CS_BIAS.n36 GND 0.075758f
C3680 CS_BIAS.n37 GND 0.004191f
C3681 CS_BIAS.n38 GND 0.007811f
C3682 CS_BIAS.n39 GND 0.004191f
C3683 CS_BIAS.n40 GND 0.007811f
C3684 CS_BIAS.n41 GND 0.004191f
C3685 CS_BIAS.n42 GND 0.004803f
C3686 CS_BIAS.n43 GND 0.004191f
C3687 CS_BIAS.t2 GND 0.19437f
C3688 CS_BIAS.n44 GND 0.075758f
C3689 CS_BIAS.n45 GND 0.007811f
C3690 CS_BIAS.n46 GND 0.004191f
C3691 CS_BIAS.n47 GND 0.007811f
C3692 CS_BIAS.n48 GND 0.004191f
C3693 CS_BIAS.t8 GND 0.19437f
C3694 CS_BIAS.n49 GND 0.075758f
C3695 CS_BIAS.n50 GND 0.004191f
C3696 CS_BIAS.n51 GND 0.007811f
C3697 CS_BIAS.n52 GND 0.004191f
C3698 CS_BIAS.n53 GND 0.007811f
C3699 CS_BIAS.n54 GND 0.004191f
C3700 CS_BIAS.n55 GND 0.005266f
C3701 CS_BIAS.n56 GND 0.004191f
C3702 CS_BIAS.t22 GND 0.19437f
C3703 CS_BIAS.n57 GND 0.075758f
C3704 CS_BIAS.n58 GND 0.007811f
C3705 CS_BIAS.n59 GND 0.004191f
C3706 CS_BIAS.n60 GND 0.007811f
C3707 CS_BIAS.n61 GND 0.004191f
C3708 CS_BIAS.t24 GND 0.19437f
C3709 CS_BIAS.n62 GND 0.094402f
C3710 CS_BIAS.t12 GND 0.273902f
C3711 CS_BIAS.n63 GND 0.126453f
C3712 CS_BIAS.n64 GND 0.052852f
C3713 CS_BIAS.n65 GND 0.007425f
C3714 CS_BIAS.n66 GND 0.007811f
C3715 CS_BIAS.n67 GND 0.007811f
C3716 CS_BIAS.n68 GND 0.004191f
C3717 CS_BIAS.n69 GND 0.004191f
C3718 CS_BIAS.n70 GND 0.004191f
C3719 CS_BIAS.n71 GND 0.007992f
C3720 CS_BIAS.n72 GND 0.003586f
C3721 CS_BIAS.n73 GND 0.008468f
C3722 CS_BIAS.n74 GND 0.004191f
C3723 CS_BIAS.n75 GND 0.004191f
C3724 CS_BIAS.n76 GND 0.004191f
C3725 CS_BIAS.n77 GND 0.007811f
C3726 CS_BIAS.n78 GND 0.007811f
C3727 CS_BIAS.n79 GND 0.006499f
C3728 CS_BIAS.n80 GND 0.004191f
C3729 CS_BIAS.n81 GND 0.004191f
C3730 CS_BIAS.n82 GND 0.004191f
C3731 CS_BIAS.n83 GND 0.007811f
C3732 CS_BIAS.n84 GND 0.007811f
C3733 CS_BIAS.n85 GND 0.007811f
C3734 CS_BIAS.n86 GND 0.004191f
C3735 CS_BIAS.n87 GND 0.004191f
C3736 CS_BIAS.n88 GND 0.004191f
C3737 CS_BIAS.n89 GND 0.005767f
C3738 CS_BIAS.n90 GND 0.006468f
C3739 CS_BIAS.n91 GND 0.007811f
C3740 CS_BIAS.n92 GND 0.004191f
C3741 CS_BIAS.n93 GND 0.004191f
C3742 CS_BIAS.n94 GND 0.004191f
C3743 CS_BIAS.n95 GND 0.007811f
C3744 CS_BIAS.n96 GND 0.007811f
C3745 CS_BIAS.n97 GND 0.004803f
C3746 CS_BIAS.n98 GND 0.004191f
C3747 CS_BIAS.n99 GND 0.004191f
C3748 CS_BIAS.n100 GND 0.006962f
C3749 CS_BIAS.n101 GND 0.007811f
C3750 CS_BIAS.n102 GND 0.007811f
C3751 CS_BIAS.n103 GND 0.004191f
C3752 CS_BIAS.n104 GND 0.004191f
C3753 CS_BIAS.n105 GND 0.004191f
C3754 CS_BIAS.n106 GND 0.008329f
C3755 CS_BIAS.n107 GND 0.003388f
C3756 CS_BIAS.n108 GND 0.008329f
C3757 CS_BIAS.n109 GND 0.004191f
C3758 CS_BIAS.n110 GND 0.004191f
C3759 CS_BIAS.n111 GND 0.004191f
C3760 CS_BIAS.n112 GND 0.007811f
C3761 CS_BIAS.n113 GND 0.007811f
C3762 CS_BIAS.n114 GND 0.006962f
C3763 CS_BIAS.n115 GND 0.004191f
C3764 CS_BIAS.n116 GND 0.004191f
C3765 CS_BIAS.n117 GND 0.004191f
C3766 CS_BIAS.n118 GND 0.007811f
C3767 CS_BIAS.n119 GND 0.007811f
C3768 CS_BIAS.n120 GND 0.007811f
C3769 CS_BIAS.n121 GND 0.004191f
C3770 CS_BIAS.n122 GND 0.004191f
C3771 CS_BIAS.n123 GND 0.004191f
C3772 CS_BIAS.n124 GND 0.006468f
C3773 CS_BIAS.n125 GND 0.005767f
C3774 CS_BIAS.n126 GND 0.007811f
C3775 CS_BIAS.n127 GND 0.004191f
C3776 CS_BIAS.n128 GND 0.004191f
C3777 CS_BIAS.n129 GND 0.004191f
C3778 CS_BIAS.n130 GND 0.007811f
C3779 CS_BIAS.n131 GND 0.007811f
C3780 CS_BIAS.n132 GND 0.005266f
C3781 CS_BIAS.n133 GND 0.004191f
C3782 CS_BIAS.n134 GND 0.004191f
C3783 CS_BIAS.n135 GND 0.006499f
C3784 CS_BIAS.n136 GND 0.007811f
C3785 CS_BIAS.n137 GND 0.007811f
C3786 CS_BIAS.n138 GND 0.004191f
C3787 CS_BIAS.n139 GND 0.004191f
C3788 CS_BIAS.n140 GND 0.004191f
C3789 CS_BIAS.n141 GND 0.008468f
C3790 CS_BIAS.n142 GND 0.003586f
C3791 CS_BIAS.n143 GND 0.007992f
C3792 CS_BIAS.n144 GND 0.004191f
C3793 CS_BIAS.n145 GND 0.004191f
C3794 CS_BIAS.n146 GND 0.004191f
C3795 CS_BIAS.n147 GND 0.007811f
C3796 CS_BIAS.n148 GND 0.007811f
C3797 CS_BIAS.n149 GND 0.007425f
C3798 CS_BIAS.n150 GND 0.004191f
C3799 CS_BIAS.n151 GND 0.004191f
C3800 CS_BIAS.n152 GND 0.004191f
C3801 CS_BIAS.n153 GND 0.007811f
C3802 CS_BIAS.n154 GND 0.007811f
C3803 CS_BIAS.n155 GND 0.007811f
C3804 CS_BIAS.n156 GND 0.004191f
C3805 CS_BIAS.n157 GND 0.004191f
C3806 CS_BIAS.n158 GND 0.004191f
C3807 CS_BIAS.n159 GND 0.007159f
C3808 CS_BIAS.n160 GND 0.005004f
C3809 CS_BIAS.n161 GND 0.007884f
C3810 CS_BIAS.n162 GND 0.004191f
C3811 CS_BIAS.n163 GND 0.004191f
C3812 CS_BIAS.n164 GND 0.004191f
C3813 CS_BIAS.n165 GND 0.007811f
C3814 CS_BIAS.n166 GND 0.007811f
C3815 CS_BIAS.n167 GND 0.005728f
C3816 CS_BIAS.n168 GND 0.008868f
C3817 CS_BIAS.n169 GND 0.062806f
C3818 CS_BIAS.t21 GND 0.004354f
C3819 CS_BIAS.t15 GND 0.004354f
C3820 CS_BIAS.n170 GND 0.032303f
C3821 CS_BIAS.n171 GND 0.080555f
C3822 CS_BIAS.t17 GND 0.004354f
C3823 CS_BIAS.t3 GND 0.004354f
C3824 CS_BIAS.n172 GND 0.032303f
C3825 CS_BIAS.n173 GND 0.052507f
C3826 CS_BIAS.t25 GND 0.004354f
C3827 CS_BIAS.t13 GND 0.004354f
C3828 CS_BIAS.n174 GND 0.036354f
C3829 CS_BIAS.t9 GND 0.004354f
C3830 CS_BIAS.t23 GND 0.004354f
C3831 CS_BIAS.n175 GND 0.032303f
C3832 CS_BIAS.n176 GND 0.114894f
C3833 CS_BIAS.n177 GND 0.052918f
C3834 CS_BIAS.n178 GND 0.030334f
C3835 CS_BIAS.n179 GND 0.007811f
C3836 CS_BIAS.n180 GND 0.004191f
C3837 CS_BIAS.t46 GND 0.19437f
C3838 CS_BIAS.n181 GND 0.075758f
C3839 CS_BIAS.n182 GND 0.004191f
C3840 CS_BIAS.n183 GND 0.007811f
C3841 CS_BIAS.n184 GND 0.004191f
C3842 CS_BIAS.n185 GND 0.007811f
C3843 CS_BIAS.n186 GND 0.004191f
C3844 CS_BIAS.n187 GND 0.005266f
C3845 CS_BIAS.n188 GND 0.004191f
C3846 CS_BIAS.t34 GND 0.19437f
C3847 CS_BIAS.n189 GND 0.075758f
C3848 CS_BIAS.n190 GND 0.007811f
C3849 CS_BIAS.n191 GND 0.004191f
C3850 CS_BIAS.n192 GND 0.007811f
C3851 CS_BIAS.n193 GND 0.004191f
C3852 CS_BIAS.t54 GND 0.19437f
C3853 CS_BIAS.n194 GND 0.094402f
C3854 CS_BIAS.t52 GND 0.273902f
C3855 CS_BIAS.n195 GND 0.126453f
C3856 CS_BIAS.n196 GND 0.052852f
C3857 CS_BIAS.n197 GND 0.007425f
C3858 CS_BIAS.n198 GND 0.007811f
C3859 CS_BIAS.n199 GND 0.007811f
C3860 CS_BIAS.n200 GND 0.004191f
C3861 CS_BIAS.n201 GND 0.004191f
C3862 CS_BIAS.n202 GND 0.004191f
C3863 CS_BIAS.n203 GND 0.007992f
C3864 CS_BIAS.n204 GND 0.003586f
C3865 CS_BIAS.n205 GND 0.008468f
C3866 CS_BIAS.n206 GND 0.004191f
C3867 CS_BIAS.n207 GND 0.004191f
C3868 CS_BIAS.n208 GND 0.004191f
C3869 CS_BIAS.n209 GND 0.007811f
C3870 CS_BIAS.n210 GND 0.007811f
C3871 CS_BIAS.n211 GND 0.006499f
C3872 CS_BIAS.n212 GND 0.004191f
C3873 CS_BIAS.n213 GND 0.004191f
C3874 CS_BIAS.n214 GND 0.004191f
C3875 CS_BIAS.n215 GND 0.007811f
C3876 CS_BIAS.n216 GND 0.007811f
C3877 CS_BIAS.n217 GND 0.007811f
C3878 CS_BIAS.n218 GND 0.004191f
C3879 CS_BIAS.n219 GND 0.004191f
C3880 CS_BIAS.n220 GND 0.004191f
C3881 CS_BIAS.n221 GND 0.005767f
C3882 CS_BIAS.n222 GND 0.006468f
C3883 CS_BIAS.n223 GND 0.007811f
C3884 CS_BIAS.n224 GND 0.004191f
C3885 CS_BIAS.n225 GND 0.004191f
C3886 CS_BIAS.n226 GND 0.004191f
C3887 CS_BIAS.n227 GND 0.007811f
C3888 CS_BIAS.n228 GND 0.007811f
C3889 CS_BIAS.n229 GND 0.004803f
C3890 CS_BIAS.n230 GND 0.004191f
C3891 CS_BIAS.n231 GND 0.004191f
C3892 CS_BIAS.n232 GND 0.006962f
C3893 CS_BIAS.n233 GND 0.007811f
C3894 CS_BIAS.n234 GND 0.007811f
C3895 CS_BIAS.n235 GND 0.004191f
C3896 CS_BIAS.n236 GND 0.004191f
C3897 CS_BIAS.n237 GND 0.004171f
C3898 CS_BIAS.n238 GND 0.008329f
C3899 CS_BIAS.n239 GND 0.003388f
C3900 CS_BIAS.n240 GND 0.008329f
C3901 CS_BIAS.n241 GND 0.004171f
C3902 CS_BIAS.n242 GND 0.004191f
C3903 CS_BIAS.n243 GND 0.004191f
C3904 CS_BIAS.n244 GND 0.007811f
C3905 CS_BIAS.n245 GND 0.007811f
C3906 CS_BIAS.n246 GND 0.006962f
C3907 CS_BIAS.n247 GND 0.004191f
C3908 CS_BIAS.n248 GND 0.004191f
C3909 CS_BIAS.n249 GND 0.004191f
C3910 CS_BIAS.n250 GND 0.007811f
C3911 CS_BIAS.n251 GND 0.007811f
C3912 CS_BIAS.n252 GND 0.007811f
C3913 CS_BIAS.n253 GND 0.004191f
C3914 CS_BIAS.n254 GND 0.004191f
C3915 CS_BIAS.n255 GND 0.004191f
C3916 CS_BIAS.n256 GND 0.006468f
C3917 CS_BIAS.n257 GND 0.005767f
C3918 CS_BIAS.n258 GND 0.007811f
C3919 CS_BIAS.n259 GND 0.004191f
C3920 CS_BIAS.n260 GND 0.004191f
C3921 CS_BIAS.n261 GND 0.004191f
C3922 CS_BIAS.n262 GND 0.007811f
C3923 CS_BIAS.n263 GND 0.007811f
C3924 CS_BIAS.n264 GND 0.005266f
C3925 CS_BIAS.n265 GND 0.004191f
C3926 CS_BIAS.n266 GND 0.004191f
C3927 CS_BIAS.n267 GND 0.006499f
C3928 CS_BIAS.n268 GND 0.007811f
C3929 CS_BIAS.n269 GND 0.007811f
C3930 CS_BIAS.n270 GND 0.004191f
C3931 CS_BIAS.n271 GND 0.004191f
C3932 CS_BIAS.n272 GND 0.004191f
C3933 CS_BIAS.n273 GND 0.008468f
C3934 CS_BIAS.n274 GND 0.003586f
C3935 CS_BIAS.n275 GND 0.007992f
C3936 CS_BIAS.n276 GND 0.004191f
C3937 CS_BIAS.n277 GND 0.004191f
C3938 CS_BIAS.n278 GND 0.004191f
C3939 CS_BIAS.n279 GND 0.007811f
C3940 CS_BIAS.n280 GND 0.007811f
C3941 CS_BIAS.n281 GND 0.007425f
C3942 CS_BIAS.n282 GND 0.004191f
C3943 CS_BIAS.n283 GND 0.004191f
C3944 CS_BIAS.n284 GND 0.004191f
C3945 CS_BIAS.n285 GND 0.007811f
C3946 CS_BIAS.n286 GND 0.007811f
C3947 CS_BIAS.n287 GND 0.007811f
C3948 CS_BIAS.n288 GND 0.004191f
C3949 CS_BIAS.n289 GND 0.004191f
C3950 CS_BIAS.n290 GND 0.004191f
C3951 CS_BIAS.n291 GND 0.007159f
C3952 CS_BIAS.n292 GND 0.005004f
C3953 CS_BIAS.n293 GND 0.007884f
C3954 CS_BIAS.n294 GND 0.004191f
C3955 CS_BIAS.n295 GND 0.004191f
C3956 CS_BIAS.n296 GND 0.004191f
C3957 CS_BIAS.n297 GND 0.007811f
C3958 CS_BIAS.n298 GND 0.007811f
C3959 CS_BIAS.n299 GND 0.005728f
C3960 CS_BIAS.n300 GND 0.008868f
C3961 CS_BIAS.n301 GND 0.048316f
C3962 CS_BIAS.t35 GND 0.19437f
C3963 CS_BIAS.n302 GND 0.093799f
C3964 CS_BIAS.n303 GND 0.004191f
C3965 CS_BIAS.n304 GND 0.007811f
C3966 CS_BIAS.n305 GND 0.004191f
C3967 CS_BIAS.n306 GND 0.007811f
C3968 CS_BIAS.n307 GND 0.004191f
C3969 CS_BIAS.n308 GND 0.00434f
C3970 CS_BIAS.n309 GND 0.004191f
C3971 CS_BIAS.t44 GND 0.19437f
C3972 CS_BIAS.n310 GND 0.075758f
C3973 CS_BIAS.n311 GND 0.007811f
C3974 CS_BIAS.n312 GND 0.004191f
C3975 CS_BIAS.n313 GND 0.007811f
C3976 CS_BIAS.n314 GND 0.004191f
C3977 CS_BIAS.t59 GND 0.19437f
C3978 CS_BIAS.n315 GND 0.075758f
C3979 CS_BIAS.n316 GND 0.004191f
C3980 CS_BIAS.n317 GND 0.007811f
C3981 CS_BIAS.n318 GND 0.004191f
C3982 CS_BIAS.n319 GND 0.007811f
C3983 CS_BIAS.n320 GND 0.004191f
C3984 CS_BIAS.n321 GND 0.004803f
C3985 CS_BIAS.n322 GND 0.004191f
C3986 CS_BIAS.t33 GND 0.19437f
C3987 CS_BIAS.n323 GND 0.075758f
C3988 CS_BIAS.n324 GND 0.007811f
C3989 CS_BIAS.n325 GND 0.004191f
C3990 CS_BIAS.n326 GND 0.007811f
C3991 CS_BIAS.n327 GND 0.004191f
C3992 CS_BIAS.t49 GND 0.19437f
C3993 CS_BIAS.n328 GND 0.075758f
C3994 CS_BIAS.n329 GND 0.004191f
C3995 CS_BIAS.n330 GND 0.007811f
C3996 CS_BIAS.n331 GND 0.004191f
C3997 CS_BIAS.n332 GND 0.007811f
C3998 CS_BIAS.n333 GND 0.004191f
C3999 CS_BIAS.n334 GND 0.005266f
C4000 CS_BIAS.n335 GND 0.004191f
C4001 CS_BIAS.t57 GND 0.19437f
C4002 CS_BIAS.n336 GND 0.075758f
C4003 CS_BIAS.n337 GND 0.007811f
C4004 CS_BIAS.n338 GND 0.004191f
C4005 CS_BIAS.n339 GND 0.007811f
C4006 CS_BIAS.n340 GND 0.004191f
C4007 CS_BIAS.t40 GND 0.19437f
C4008 CS_BIAS.n341 GND 0.094402f
C4009 CS_BIAS.t47 GND 0.273902f
C4010 CS_BIAS.n342 GND 0.126453f
C4011 CS_BIAS.n343 GND 0.052852f
C4012 CS_BIAS.n344 GND 0.007425f
C4013 CS_BIAS.n345 GND 0.007811f
C4014 CS_BIAS.n346 GND 0.007811f
C4015 CS_BIAS.n347 GND 0.004191f
C4016 CS_BIAS.n348 GND 0.004191f
C4017 CS_BIAS.n349 GND 0.004191f
C4018 CS_BIAS.n350 GND 0.007992f
C4019 CS_BIAS.n351 GND 0.003586f
C4020 CS_BIAS.n352 GND 0.008468f
C4021 CS_BIAS.n353 GND 0.004191f
C4022 CS_BIAS.n354 GND 0.004191f
C4023 CS_BIAS.n355 GND 0.004191f
C4024 CS_BIAS.n356 GND 0.007811f
C4025 CS_BIAS.n357 GND 0.007811f
C4026 CS_BIAS.n358 GND 0.006499f
C4027 CS_BIAS.n359 GND 0.004191f
C4028 CS_BIAS.n360 GND 0.004191f
C4029 CS_BIAS.n361 GND 0.004191f
C4030 CS_BIAS.n362 GND 0.007811f
C4031 CS_BIAS.n363 GND 0.007811f
C4032 CS_BIAS.n364 GND 0.007811f
C4033 CS_BIAS.n365 GND 0.004191f
C4034 CS_BIAS.n366 GND 0.004191f
C4035 CS_BIAS.n367 GND 0.004191f
C4036 CS_BIAS.n368 GND 0.005767f
C4037 CS_BIAS.n369 GND 0.006468f
C4038 CS_BIAS.n370 GND 0.007811f
C4039 CS_BIAS.n371 GND 0.004191f
C4040 CS_BIAS.n372 GND 0.004191f
C4041 CS_BIAS.n373 GND 0.004191f
C4042 CS_BIAS.n374 GND 0.007811f
C4043 CS_BIAS.n375 GND 0.007811f
C4044 CS_BIAS.n376 GND 0.004803f
C4045 CS_BIAS.n377 GND 0.004191f
C4046 CS_BIAS.n378 GND 0.004191f
C4047 CS_BIAS.n379 GND 0.006962f
C4048 CS_BIAS.n380 GND 0.007811f
C4049 CS_BIAS.n381 GND 0.007811f
C4050 CS_BIAS.n382 GND 0.004191f
C4051 CS_BIAS.n383 GND 0.004191f
C4052 CS_BIAS.n384 GND 0.004191f
C4053 CS_BIAS.n385 GND 0.008329f
C4054 CS_BIAS.n386 GND 0.003388f
C4055 CS_BIAS.n387 GND 0.008329f
C4056 CS_BIAS.n388 GND 0.004191f
C4057 CS_BIAS.n389 GND 0.004191f
C4058 CS_BIAS.n390 GND 0.004191f
C4059 CS_BIAS.n391 GND 0.007811f
C4060 CS_BIAS.n392 GND 0.007811f
C4061 CS_BIAS.n393 GND 0.006962f
C4062 CS_BIAS.n394 GND 0.004191f
C4063 CS_BIAS.n395 GND 0.004191f
C4064 CS_BIAS.n396 GND 0.004191f
C4065 CS_BIAS.n397 GND 0.007811f
C4066 CS_BIAS.n398 GND 0.007811f
C4067 CS_BIAS.n399 GND 0.007811f
C4068 CS_BIAS.n400 GND 0.004191f
C4069 CS_BIAS.n401 GND 0.004191f
C4070 CS_BIAS.n402 GND 0.004191f
C4071 CS_BIAS.n403 GND 0.006468f
C4072 CS_BIAS.n404 GND 0.005767f
C4073 CS_BIAS.n405 GND 0.007811f
C4074 CS_BIAS.n406 GND 0.004191f
C4075 CS_BIAS.n407 GND 0.004191f
C4076 CS_BIAS.n408 GND 0.004191f
C4077 CS_BIAS.n409 GND 0.007811f
C4078 CS_BIAS.n410 GND 0.007811f
C4079 CS_BIAS.n411 GND 0.005266f
C4080 CS_BIAS.n412 GND 0.004191f
C4081 CS_BIAS.n413 GND 0.004191f
C4082 CS_BIAS.n414 GND 0.006499f
C4083 CS_BIAS.n415 GND 0.007811f
C4084 CS_BIAS.n416 GND 0.007811f
C4085 CS_BIAS.n417 GND 0.004191f
C4086 CS_BIAS.n418 GND 0.004191f
C4087 CS_BIAS.n419 GND 0.004191f
C4088 CS_BIAS.n420 GND 0.008468f
C4089 CS_BIAS.n421 GND 0.003586f
C4090 CS_BIAS.n422 GND 0.007992f
C4091 CS_BIAS.n423 GND 0.004191f
C4092 CS_BIAS.n424 GND 0.004191f
C4093 CS_BIAS.n425 GND 0.004191f
C4094 CS_BIAS.n426 GND 0.007811f
C4095 CS_BIAS.n427 GND 0.007811f
C4096 CS_BIAS.n428 GND 0.007425f
C4097 CS_BIAS.n429 GND 0.004191f
C4098 CS_BIAS.n430 GND 0.004191f
C4099 CS_BIAS.n431 GND 0.004191f
C4100 CS_BIAS.n432 GND 0.007811f
C4101 CS_BIAS.n433 GND 0.007811f
C4102 CS_BIAS.n434 GND 0.007811f
C4103 CS_BIAS.n435 GND 0.004191f
C4104 CS_BIAS.n436 GND 0.004191f
C4105 CS_BIAS.n437 GND 0.004191f
C4106 CS_BIAS.n438 GND 0.007159f
C4107 CS_BIAS.n439 GND 0.005004f
C4108 CS_BIAS.n440 GND 0.007884f
C4109 CS_BIAS.n441 GND 0.004191f
C4110 CS_BIAS.n442 GND 0.004191f
C4111 CS_BIAS.n443 GND 0.004191f
C4112 CS_BIAS.n444 GND 0.007811f
C4113 CS_BIAS.n445 GND 0.007811f
C4114 CS_BIAS.n446 GND 0.005728f
C4115 CS_BIAS.n447 GND 0.008868f
C4116 CS_BIAS.n448 GND 0.043009f
C4117 CS_BIAS.n449 GND 0.3056f
C4118 CS_BIAS.t36 GND 0.19437f
C4119 CS_BIAS.n450 GND 0.093799f
C4120 CS_BIAS.n451 GND 0.004191f
C4121 CS_BIAS.n452 GND 0.007811f
C4122 CS_BIAS.n453 GND 0.004191f
C4123 CS_BIAS.n454 GND 0.007811f
C4124 CS_BIAS.n455 GND 0.004191f
C4125 CS_BIAS.n456 GND 0.00434f
C4126 CS_BIAS.n457 GND 0.004191f
C4127 CS_BIAS.n458 GND 0.007811f
C4128 CS_BIAS.n459 GND 0.004191f
C4129 CS_BIAS.n460 GND 0.007811f
C4130 CS_BIAS.n461 GND 0.004191f
C4131 CS_BIAS.t56 GND 0.19437f
C4132 CS_BIAS.n462 GND 0.075758f
C4133 CS_BIAS.n463 GND 0.004191f
C4134 CS_BIAS.n464 GND 0.007811f
C4135 CS_BIAS.n465 GND 0.004191f
C4136 CS_BIAS.n466 GND 0.007811f
C4137 CS_BIAS.n467 GND 0.004191f
C4138 CS_BIAS.n468 GND 0.004803f
C4139 CS_BIAS.n469 GND 0.004191f
C4140 CS_BIAS.n470 GND 0.007811f
C4141 CS_BIAS.t7 GND 0.004354f
C4142 CS_BIAS.t5 GND 0.004354f
C4143 CS_BIAS.n471 GND 0.036354f
C4144 CS_BIAS.t1 GND 0.004354f
C4145 CS_BIAS.t31 GND 0.004354f
C4146 CS_BIAS.n472 GND 0.032303f
C4147 CS_BIAS.n473 GND 0.114894f
C4148 CS_BIAS.t18 GND 0.19437f
C4149 CS_BIAS.n474 GND 0.093799f
C4150 CS_BIAS.n475 GND 0.004191f
C4151 CS_BIAS.n476 GND 0.007811f
C4152 CS_BIAS.n477 GND 0.004191f
C4153 CS_BIAS.n478 GND 0.007811f
C4154 CS_BIAS.n479 GND 0.004191f
C4155 CS_BIAS.n480 GND 0.00434f
C4156 CS_BIAS.n481 GND 0.004191f
C4157 CS_BIAS.n482 GND 0.007811f
C4158 CS_BIAS.n483 GND 0.004191f
C4159 CS_BIAS.n484 GND 0.007811f
C4160 CS_BIAS.n485 GND 0.004191f
C4161 CS_BIAS.t10 GND 0.19437f
C4162 CS_BIAS.n486 GND 0.075758f
C4163 CS_BIAS.n487 GND 0.004191f
C4164 CS_BIAS.n488 GND 0.007811f
C4165 CS_BIAS.n489 GND 0.004191f
C4166 CS_BIAS.n490 GND 0.007811f
C4167 CS_BIAS.n491 GND 0.004191f
C4168 CS_BIAS.n492 GND 0.004803f
C4169 CS_BIAS.n493 GND 0.004191f
C4170 CS_BIAS.n494 GND 0.007811f
C4171 CS_BIAS.n495 GND 0.004191f
C4172 CS_BIAS.n496 GND 0.007811f
C4173 CS_BIAS.n497 GND 0.004191f
C4174 CS_BIAS.t30 GND 0.19437f
C4175 CS_BIAS.n498 GND 0.075758f
C4176 CS_BIAS.n499 GND 0.004191f
C4177 CS_BIAS.n500 GND 0.007811f
C4178 CS_BIAS.n501 GND 0.004191f
C4179 CS_BIAS.n502 GND 0.007811f
C4180 CS_BIAS.n503 GND 0.004191f
C4181 CS_BIAS.n504 GND 0.005266f
C4182 CS_BIAS.n505 GND 0.004191f
C4183 CS_BIAS.n506 GND 0.007811f
C4184 CS_BIAS.n507 GND 0.004191f
C4185 CS_BIAS.n508 GND 0.007811f
C4186 CS_BIAS.n509 GND 0.004191f
C4187 CS_BIAS.t4 GND 0.19437f
C4188 CS_BIAS.n510 GND 0.094402f
C4189 CS_BIAS.t6 GND 0.273902f
C4190 CS_BIAS.n511 GND 0.126453f
C4191 CS_BIAS.n512 GND 0.052852f
C4192 CS_BIAS.n513 GND 0.007425f
C4193 CS_BIAS.n514 GND 0.007811f
C4194 CS_BIAS.n515 GND 0.007811f
C4195 CS_BIAS.n516 GND 0.004191f
C4196 CS_BIAS.n517 GND 0.004191f
C4197 CS_BIAS.n518 GND 0.004191f
C4198 CS_BIAS.n519 GND 0.007992f
C4199 CS_BIAS.n520 GND 0.003586f
C4200 CS_BIAS.n521 GND 0.008468f
C4201 CS_BIAS.n522 GND 0.004191f
C4202 CS_BIAS.n523 GND 0.004191f
C4203 CS_BIAS.n524 GND 0.004191f
C4204 CS_BIAS.n525 GND 0.007811f
C4205 CS_BIAS.n526 GND 0.007811f
C4206 CS_BIAS.t0 GND 0.19437f
C4207 CS_BIAS.n527 GND 0.075758f
C4208 CS_BIAS.n528 GND 0.006499f
C4209 CS_BIAS.n529 GND 0.004191f
C4210 CS_BIAS.n530 GND 0.004191f
C4211 CS_BIAS.n531 GND 0.004191f
C4212 CS_BIAS.n532 GND 0.007811f
C4213 CS_BIAS.n533 GND 0.007811f
C4214 CS_BIAS.n534 GND 0.007811f
C4215 CS_BIAS.n535 GND 0.004191f
C4216 CS_BIAS.n536 GND 0.004191f
C4217 CS_BIAS.n537 GND 0.004191f
C4218 CS_BIAS.n538 GND 0.005767f
C4219 CS_BIAS.n539 GND 0.006468f
C4220 CS_BIAS.n540 GND 0.007811f
C4221 CS_BIAS.n541 GND 0.004191f
C4222 CS_BIAS.n542 GND 0.004191f
C4223 CS_BIAS.n543 GND 0.004191f
C4224 CS_BIAS.n544 GND 0.007811f
C4225 CS_BIAS.n545 GND 0.007811f
C4226 CS_BIAS.n546 GND 0.004803f
C4227 CS_BIAS.n547 GND 0.004191f
C4228 CS_BIAS.n548 GND 0.004191f
C4229 CS_BIAS.n549 GND 0.006962f
C4230 CS_BIAS.n550 GND 0.007811f
C4231 CS_BIAS.n551 GND 0.007811f
C4232 CS_BIAS.n552 GND 0.004191f
C4233 CS_BIAS.n553 GND 0.004191f
C4234 CS_BIAS.n554 GND 0.004191f
C4235 CS_BIAS.n555 GND 0.008329f
C4236 CS_BIAS.n556 GND 0.003388f
C4237 CS_BIAS.n557 GND 0.008329f
C4238 CS_BIAS.n558 GND 0.004191f
C4239 CS_BIAS.n559 GND 0.004191f
C4240 CS_BIAS.n560 GND 0.004191f
C4241 CS_BIAS.n561 GND 0.007811f
C4242 CS_BIAS.n562 GND 0.007811f
C4243 CS_BIAS.t28 GND 0.19437f
C4244 CS_BIAS.n563 GND 0.075758f
C4245 CS_BIAS.n564 GND 0.006962f
C4246 CS_BIAS.n565 GND 0.004191f
C4247 CS_BIAS.n566 GND 0.004191f
C4248 CS_BIAS.n567 GND 0.004191f
C4249 CS_BIAS.n568 GND 0.007811f
C4250 CS_BIAS.n569 GND 0.007811f
C4251 CS_BIAS.n570 GND 0.007811f
C4252 CS_BIAS.n571 GND 0.004191f
C4253 CS_BIAS.n572 GND 0.004191f
C4254 CS_BIAS.n573 GND 0.004191f
C4255 CS_BIAS.n574 GND 0.006468f
C4256 CS_BIAS.n575 GND 0.005767f
C4257 CS_BIAS.n576 GND 0.007811f
C4258 CS_BIAS.n577 GND 0.004191f
C4259 CS_BIAS.n578 GND 0.004191f
C4260 CS_BIAS.n579 GND 0.004191f
C4261 CS_BIAS.n580 GND 0.007811f
C4262 CS_BIAS.n581 GND 0.007811f
C4263 CS_BIAS.n582 GND 0.005266f
C4264 CS_BIAS.n583 GND 0.004191f
C4265 CS_BIAS.n584 GND 0.004191f
C4266 CS_BIAS.n585 GND 0.006499f
C4267 CS_BIAS.n586 GND 0.007811f
C4268 CS_BIAS.n587 GND 0.007811f
C4269 CS_BIAS.n588 GND 0.004191f
C4270 CS_BIAS.n589 GND 0.004191f
C4271 CS_BIAS.n590 GND 0.004191f
C4272 CS_BIAS.n591 GND 0.008468f
C4273 CS_BIAS.n592 GND 0.003586f
C4274 CS_BIAS.n593 GND 0.007992f
C4275 CS_BIAS.n594 GND 0.004191f
C4276 CS_BIAS.n595 GND 0.004191f
C4277 CS_BIAS.n596 GND 0.004191f
C4278 CS_BIAS.n597 GND 0.007811f
C4279 CS_BIAS.n598 GND 0.007811f
C4280 CS_BIAS.t26 GND 0.19437f
C4281 CS_BIAS.n599 GND 0.075758f
C4282 CS_BIAS.n600 GND 0.007425f
C4283 CS_BIAS.n601 GND 0.004191f
C4284 CS_BIAS.n602 GND 0.004191f
C4285 CS_BIAS.n603 GND 0.004191f
C4286 CS_BIAS.n604 GND 0.007811f
C4287 CS_BIAS.n605 GND 0.007811f
C4288 CS_BIAS.n606 GND 0.007811f
C4289 CS_BIAS.n607 GND 0.004191f
C4290 CS_BIAS.n608 GND 0.004191f
C4291 CS_BIAS.n609 GND 0.004191f
C4292 CS_BIAS.n610 GND 0.007159f
C4293 CS_BIAS.n611 GND 0.005004f
C4294 CS_BIAS.n612 GND 0.007884f
C4295 CS_BIAS.n613 GND 0.004191f
C4296 CS_BIAS.n614 GND 0.004191f
C4297 CS_BIAS.n615 GND 0.004191f
C4298 CS_BIAS.n616 GND 0.007811f
C4299 CS_BIAS.n617 GND 0.007811f
C4300 CS_BIAS.n618 GND 0.005728f
C4301 CS_BIAS.n619 GND 0.008868f
C4302 CS_BIAS.n620 GND 0.062806f
C4303 CS_BIAS.t27 GND 0.004354f
C4304 CS_BIAS.t19 GND 0.004354f
C4305 CS_BIAS.n621 GND 0.032303f
C4306 CS_BIAS.n622 GND 0.080555f
C4307 CS_BIAS.t29 GND 0.004354f
C4308 CS_BIAS.t11 GND 0.004354f
C4309 CS_BIAS.n623 GND 0.032303f
C4310 CS_BIAS.n624 GND 0.052507f
C4311 CS_BIAS.n625 GND 0.052918f
C4312 CS_BIAS.n626 GND 0.030334f
C4313 CS_BIAS.n627 GND 0.007811f
C4314 CS_BIAS.n628 GND 0.004191f
C4315 CS_BIAS.t32 GND 0.19437f
C4316 CS_BIAS.n629 GND 0.075758f
C4317 CS_BIAS.n630 GND 0.004191f
C4318 CS_BIAS.n631 GND 0.007811f
C4319 CS_BIAS.n632 GND 0.004191f
C4320 CS_BIAS.n633 GND 0.007811f
C4321 CS_BIAS.n634 GND 0.004191f
C4322 CS_BIAS.n635 GND 0.005266f
C4323 CS_BIAS.n636 GND 0.004191f
C4324 CS_BIAS.n637 GND 0.007811f
C4325 CS_BIAS.n638 GND 0.004191f
C4326 CS_BIAS.n639 GND 0.007811f
C4327 CS_BIAS.n640 GND 0.004191f
C4328 CS_BIAS.t43 GND 0.19437f
C4329 CS_BIAS.n641 GND 0.094402f
C4330 CS_BIAS.t61 GND 0.273902f
C4331 CS_BIAS.n642 GND 0.126453f
C4332 CS_BIAS.n643 GND 0.052852f
C4333 CS_BIAS.n644 GND 0.007425f
C4334 CS_BIAS.n645 GND 0.007811f
C4335 CS_BIAS.n646 GND 0.007811f
C4336 CS_BIAS.n647 GND 0.004191f
C4337 CS_BIAS.n648 GND 0.004191f
C4338 CS_BIAS.n649 GND 0.004191f
C4339 CS_BIAS.n650 GND 0.007992f
C4340 CS_BIAS.n651 GND 0.003586f
C4341 CS_BIAS.n652 GND 0.008468f
C4342 CS_BIAS.n653 GND 0.004191f
C4343 CS_BIAS.n654 GND 0.004191f
C4344 CS_BIAS.n655 GND 0.004191f
C4345 CS_BIAS.n656 GND 0.007811f
C4346 CS_BIAS.n657 GND 0.007811f
C4347 CS_BIAS.t53 GND 0.19437f
C4348 CS_BIAS.n658 GND 0.075758f
C4349 CS_BIAS.n659 GND 0.006499f
C4350 CS_BIAS.n660 GND 0.004191f
C4351 CS_BIAS.n661 GND 0.004191f
C4352 CS_BIAS.n662 GND 0.004191f
C4353 CS_BIAS.n663 GND 0.007811f
C4354 CS_BIAS.n664 GND 0.007811f
C4355 CS_BIAS.n665 GND 0.007811f
C4356 CS_BIAS.n666 GND 0.004191f
C4357 CS_BIAS.n667 GND 0.004191f
C4358 CS_BIAS.n668 GND 0.004191f
C4359 CS_BIAS.n669 GND 0.005767f
C4360 CS_BIAS.n670 GND 0.006468f
C4361 CS_BIAS.n671 GND 0.007811f
C4362 CS_BIAS.n672 GND 0.004191f
C4363 CS_BIAS.n673 GND 0.004191f
C4364 CS_BIAS.n674 GND 0.004191f
C4365 CS_BIAS.n675 GND 0.007811f
C4366 CS_BIAS.n676 GND 0.007811f
C4367 CS_BIAS.n677 GND 0.004803f
C4368 CS_BIAS.n678 GND 0.004191f
C4369 CS_BIAS.n679 GND 0.004191f
C4370 CS_BIAS.n680 GND 0.006962f
C4371 CS_BIAS.n681 GND 0.007811f
C4372 CS_BIAS.n682 GND 0.007811f
C4373 CS_BIAS.n683 GND 0.004191f
C4374 CS_BIAS.n684 GND 0.004191f
C4375 CS_BIAS.n685 GND 0.004171f
C4376 CS_BIAS.n686 GND 0.008329f
C4377 CS_BIAS.n687 GND 0.003388f
C4378 CS_BIAS.n688 GND 0.008329f
C4379 CS_BIAS.n689 GND 0.004171f
C4380 CS_BIAS.n690 GND 0.004191f
C4381 CS_BIAS.n691 GND 0.004191f
C4382 CS_BIAS.n692 GND 0.007811f
C4383 CS_BIAS.n693 GND 0.007811f
C4384 CS_BIAS.t45 GND 0.19437f
C4385 CS_BIAS.n694 GND 0.075758f
C4386 CS_BIAS.n695 GND 0.006962f
C4387 CS_BIAS.n696 GND 0.004191f
C4388 CS_BIAS.n697 GND 0.004191f
C4389 CS_BIAS.n698 GND 0.004191f
C4390 CS_BIAS.n699 GND 0.007811f
C4391 CS_BIAS.n700 GND 0.007811f
C4392 CS_BIAS.n701 GND 0.007811f
C4393 CS_BIAS.n702 GND 0.004191f
C4394 CS_BIAS.n703 GND 0.004191f
C4395 CS_BIAS.n704 GND 0.004191f
C4396 CS_BIAS.n705 GND 0.006468f
C4397 CS_BIAS.n706 GND 0.005767f
C4398 CS_BIAS.n707 GND 0.007811f
C4399 CS_BIAS.n708 GND 0.004191f
C4400 CS_BIAS.n709 GND 0.004191f
C4401 CS_BIAS.n710 GND 0.004191f
C4402 CS_BIAS.n711 GND 0.007811f
C4403 CS_BIAS.n712 GND 0.007811f
C4404 CS_BIAS.n713 GND 0.005266f
C4405 CS_BIAS.n714 GND 0.004191f
C4406 CS_BIAS.n715 GND 0.004191f
C4407 CS_BIAS.n716 GND 0.006499f
C4408 CS_BIAS.n717 GND 0.007811f
C4409 CS_BIAS.n718 GND 0.007811f
C4410 CS_BIAS.n719 GND 0.004191f
C4411 CS_BIAS.n720 GND 0.004191f
C4412 CS_BIAS.n721 GND 0.004191f
C4413 CS_BIAS.n722 GND 0.008468f
C4414 CS_BIAS.n723 GND 0.003586f
C4415 CS_BIAS.n724 GND 0.007992f
C4416 CS_BIAS.n725 GND 0.004191f
C4417 CS_BIAS.n726 GND 0.004191f
C4418 CS_BIAS.n727 GND 0.004191f
C4419 CS_BIAS.n728 GND 0.007811f
C4420 CS_BIAS.n729 GND 0.007811f
C4421 CS_BIAS.t62 GND 0.19437f
C4422 CS_BIAS.n730 GND 0.075758f
C4423 CS_BIAS.n731 GND 0.007425f
C4424 CS_BIAS.n732 GND 0.004191f
C4425 CS_BIAS.n733 GND 0.004191f
C4426 CS_BIAS.n734 GND 0.004191f
C4427 CS_BIAS.n735 GND 0.007811f
C4428 CS_BIAS.n736 GND 0.007811f
C4429 CS_BIAS.n737 GND 0.007811f
C4430 CS_BIAS.n738 GND 0.004191f
C4431 CS_BIAS.n739 GND 0.004191f
C4432 CS_BIAS.n740 GND 0.004191f
C4433 CS_BIAS.n741 GND 0.007159f
C4434 CS_BIAS.n742 GND 0.005004f
C4435 CS_BIAS.n743 GND 0.007884f
C4436 CS_BIAS.n744 GND 0.004191f
C4437 CS_BIAS.n745 GND 0.004191f
C4438 CS_BIAS.n746 GND 0.004191f
C4439 CS_BIAS.n747 GND 0.007811f
C4440 CS_BIAS.n748 GND 0.007811f
C4441 CS_BIAS.n749 GND 0.005728f
C4442 CS_BIAS.n750 GND 0.008868f
C4443 CS_BIAS.n751 GND 0.048316f
C4444 CS_BIAS.t60 GND 0.19437f
C4445 CS_BIAS.n752 GND 0.093799f
C4446 CS_BIAS.n753 GND 0.004191f
C4447 CS_BIAS.n754 GND 0.007811f
C4448 CS_BIAS.n755 GND 0.004191f
C4449 CS_BIAS.n756 GND 0.007811f
C4450 CS_BIAS.n757 GND 0.004191f
C4451 CS_BIAS.n758 GND 0.00434f
C4452 CS_BIAS.n759 GND 0.004191f
C4453 CS_BIAS.n760 GND 0.007811f
C4454 CS_BIAS.n761 GND 0.004191f
C4455 CS_BIAS.n762 GND 0.007811f
C4456 CS_BIAS.n763 GND 0.004191f
C4457 CS_BIAS.t42 GND 0.19437f
C4458 CS_BIAS.n764 GND 0.075758f
C4459 CS_BIAS.n765 GND 0.004191f
C4460 CS_BIAS.n766 GND 0.007811f
C4461 CS_BIAS.n767 GND 0.004191f
C4462 CS_BIAS.n768 GND 0.007811f
C4463 CS_BIAS.n769 GND 0.004191f
C4464 CS_BIAS.n770 GND 0.004803f
C4465 CS_BIAS.n771 GND 0.004191f
C4466 CS_BIAS.n772 GND 0.007811f
C4467 CS_BIAS.n773 GND 0.004191f
C4468 CS_BIAS.n774 GND 0.007811f
C4469 CS_BIAS.n775 GND 0.004191f
C4470 CS_BIAS.t63 GND 0.19437f
C4471 CS_BIAS.n776 GND 0.075758f
C4472 CS_BIAS.n777 GND 0.004191f
C4473 CS_BIAS.n778 GND 0.007811f
C4474 CS_BIAS.n779 GND 0.004191f
C4475 CS_BIAS.n780 GND 0.007811f
C4476 CS_BIAS.n781 GND 0.004191f
C4477 CS_BIAS.n782 GND 0.005266f
C4478 CS_BIAS.n783 GND 0.004191f
C4479 CS_BIAS.n784 GND 0.007811f
C4480 CS_BIAS.n785 GND 0.004191f
C4481 CS_BIAS.n786 GND 0.007811f
C4482 CS_BIAS.n787 GND 0.004191f
C4483 CS_BIAS.t55 GND 0.19437f
C4484 CS_BIAS.n788 GND 0.094402f
C4485 CS_BIAS.t39 GND 0.273902f
C4486 CS_BIAS.n789 GND 0.126453f
C4487 CS_BIAS.n790 GND 0.052852f
C4488 CS_BIAS.n791 GND 0.007425f
C4489 CS_BIAS.n792 GND 0.007811f
C4490 CS_BIAS.n793 GND 0.007811f
C4491 CS_BIAS.n794 GND 0.004191f
C4492 CS_BIAS.n795 GND 0.004191f
C4493 CS_BIAS.n796 GND 0.004191f
C4494 CS_BIAS.n797 GND 0.007992f
C4495 CS_BIAS.n798 GND 0.003586f
C4496 CS_BIAS.n799 GND 0.008468f
C4497 CS_BIAS.n800 GND 0.004191f
C4498 CS_BIAS.n801 GND 0.004191f
C4499 CS_BIAS.n802 GND 0.004191f
C4500 CS_BIAS.n803 GND 0.007811f
C4501 CS_BIAS.n804 GND 0.007811f
C4502 CS_BIAS.t41 GND 0.19437f
C4503 CS_BIAS.n805 GND 0.075758f
C4504 CS_BIAS.n806 GND 0.006499f
C4505 CS_BIAS.n807 GND 0.004191f
C4506 CS_BIAS.n808 GND 0.004191f
C4507 CS_BIAS.n809 GND 0.004191f
C4508 CS_BIAS.n810 GND 0.007811f
C4509 CS_BIAS.n811 GND 0.007811f
C4510 CS_BIAS.n812 GND 0.007811f
C4511 CS_BIAS.n813 GND 0.004191f
C4512 CS_BIAS.n814 GND 0.004191f
C4513 CS_BIAS.n815 GND 0.004191f
C4514 CS_BIAS.n816 GND 0.005767f
C4515 CS_BIAS.n817 GND 0.006468f
C4516 CS_BIAS.n818 GND 0.007811f
C4517 CS_BIAS.n819 GND 0.004191f
C4518 CS_BIAS.n820 GND 0.004191f
C4519 CS_BIAS.n821 GND 0.004191f
C4520 CS_BIAS.n822 GND 0.007811f
C4521 CS_BIAS.n823 GND 0.007811f
C4522 CS_BIAS.n824 GND 0.004803f
C4523 CS_BIAS.n825 GND 0.004191f
C4524 CS_BIAS.n826 GND 0.004191f
C4525 CS_BIAS.n827 GND 0.006962f
C4526 CS_BIAS.n828 GND 0.007811f
C4527 CS_BIAS.n829 GND 0.007811f
C4528 CS_BIAS.n830 GND 0.004191f
C4529 CS_BIAS.n831 GND 0.004191f
C4530 CS_BIAS.n832 GND 0.004191f
C4531 CS_BIAS.n833 GND 0.008329f
C4532 CS_BIAS.n834 GND 0.003388f
C4533 CS_BIAS.n835 GND 0.008329f
C4534 CS_BIAS.n836 GND 0.004191f
C4535 CS_BIAS.n837 GND 0.004191f
C4536 CS_BIAS.n838 GND 0.004191f
C4537 CS_BIAS.n839 GND 0.007811f
C4538 CS_BIAS.n840 GND 0.007811f
C4539 CS_BIAS.t50 GND 0.19437f
C4540 CS_BIAS.n841 GND 0.075758f
C4541 CS_BIAS.n842 GND 0.006962f
C4542 CS_BIAS.n843 GND 0.004191f
C4543 CS_BIAS.n844 GND 0.004191f
C4544 CS_BIAS.n845 GND 0.004191f
C4545 CS_BIAS.n846 GND 0.007811f
C4546 CS_BIAS.n847 GND 0.007811f
C4547 CS_BIAS.n848 GND 0.007811f
C4548 CS_BIAS.n849 GND 0.004191f
C4549 CS_BIAS.n850 GND 0.004191f
C4550 CS_BIAS.n851 GND 0.004191f
C4551 CS_BIAS.n852 GND 0.006468f
C4552 CS_BIAS.n853 GND 0.005767f
C4553 CS_BIAS.n854 GND 0.007811f
C4554 CS_BIAS.n855 GND 0.004191f
C4555 CS_BIAS.n856 GND 0.004191f
C4556 CS_BIAS.n857 GND 0.004191f
C4557 CS_BIAS.n858 GND 0.007811f
C4558 CS_BIAS.n859 GND 0.007811f
C4559 CS_BIAS.n860 GND 0.005266f
C4560 CS_BIAS.n861 GND 0.004191f
C4561 CS_BIAS.n862 GND 0.004191f
C4562 CS_BIAS.n863 GND 0.006499f
C4563 CS_BIAS.n864 GND 0.007811f
C4564 CS_BIAS.n865 GND 0.007811f
C4565 CS_BIAS.n866 GND 0.004191f
C4566 CS_BIAS.n867 GND 0.004191f
C4567 CS_BIAS.n868 GND 0.004191f
C4568 CS_BIAS.n869 GND 0.008468f
C4569 CS_BIAS.n870 GND 0.003586f
C4570 CS_BIAS.n871 GND 0.007992f
C4571 CS_BIAS.n872 GND 0.004191f
C4572 CS_BIAS.n873 GND 0.004191f
C4573 CS_BIAS.n874 GND 0.004191f
C4574 CS_BIAS.n875 GND 0.007811f
C4575 CS_BIAS.n876 GND 0.007811f
C4576 CS_BIAS.t37 GND 0.19437f
C4577 CS_BIAS.n877 GND 0.075758f
C4578 CS_BIAS.n878 GND 0.007425f
C4579 CS_BIAS.n879 GND 0.004191f
C4580 CS_BIAS.n880 GND 0.004191f
C4581 CS_BIAS.n881 GND 0.004191f
C4582 CS_BIAS.n882 GND 0.007811f
C4583 CS_BIAS.n883 GND 0.007811f
C4584 CS_BIAS.n884 GND 0.007811f
C4585 CS_BIAS.n885 GND 0.004191f
C4586 CS_BIAS.n886 GND 0.004191f
C4587 CS_BIAS.n887 GND 0.004191f
C4588 CS_BIAS.n888 GND 0.007159f
C4589 CS_BIAS.n889 GND 0.005004f
C4590 CS_BIAS.n890 GND 0.007884f
C4591 CS_BIAS.n891 GND 0.004191f
C4592 CS_BIAS.n892 GND 0.004191f
C4593 CS_BIAS.n893 GND 0.004191f
C4594 CS_BIAS.n894 GND 0.007811f
C4595 CS_BIAS.n895 GND 0.007811f
C4596 CS_BIAS.n896 GND 0.005728f
C4597 CS_BIAS.n897 GND 0.008868f
C4598 CS_BIAS.n898 GND 0.043009f
C4599 CS_BIAS.n899 GND 0.097271f
C4600 CS_BIAS.n900 GND 3.06527f
.ends

