* NGSPICE file created from diff_pair_sample_1338.ext - technology: sky130A

.subckt diff_pair_sample_1338 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=0 ps=0 w=15.62 l=1.46
X1 VDD2.t1 VN.t0 VTAIL.t2 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=6.0918 ps=32.02 w=15.62 l=1.46
X2 VDD1.t1 VP.t0 VTAIL.t0 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=6.0918 ps=32.02 w=15.62 l=1.46
X3 VDD1.t0 VP.t1 VTAIL.t3 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=6.0918 ps=32.02 w=15.62 l=1.46
X4 B.t8 B.t6 B.t7 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=0 ps=0 w=15.62 l=1.46
X5 VDD2.t0 VN.t1 VTAIL.t1 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=6.0918 ps=32.02 w=15.62 l=1.46
X6 B.t5 B.t3 B.t4 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=0 ps=0 w=15.62 l=1.46
X7 B.t2 B.t0 B.t1 w_n1686_n4092# sky130_fd_pr__pfet_01v8 ad=6.0918 pd=32.02 as=0 ps=0 w=15.62 l=1.46
R0 B.n359 B.n358 585
R1 B.n357 B.n92 585
R2 B.n356 B.n355 585
R3 B.n354 B.n93 585
R4 B.n353 B.n352 585
R5 B.n351 B.n94 585
R6 B.n350 B.n349 585
R7 B.n348 B.n95 585
R8 B.n347 B.n346 585
R9 B.n345 B.n96 585
R10 B.n344 B.n343 585
R11 B.n342 B.n97 585
R12 B.n341 B.n340 585
R13 B.n339 B.n98 585
R14 B.n338 B.n337 585
R15 B.n336 B.n99 585
R16 B.n335 B.n334 585
R17 B.n333 B.n100 585
R18 B.n332 B.n331 585
R19 B.n330 B.n101 585
R20 B.n329 B.n328 585
R21 B.n327 B.n102 585
R22 B.n326 B.n325 585
R23 B.n324 B.n103 585
R24 B.n323 B.n322 585
R25 B.n321 B.n104 585
R26 B.n320 B.n319 585
R27 B.n318 B.n105 585
R28 B.n317 B.n316 585
R29 B.n315 B.n106 585
R30 B.n314 B.n313 585
R31 B.n312 B.n107 585
R32 B.n311 B.n310 585
R33 B.n309 B.n108 585
R34 B.n308 B.n307 585
R35 B.n306 B.n109 585
R36 B.n305 B.n304 585
R37 B.n303 B.n110 585
R38 B.n302 B.n301 585
R39 B.n300 B.n111 585
R40 B.n299 B.n298 585
R41 B.n297 B.n112 585
R42 B.n296 B.n295 585
R43 B.n294 B.n113 585
R44 B.n293 B.n292 585
R45 B.n291 B.n114 585
R46 B.n290 B.n289 585
R47 B.n288 B.n115 585
R48 B.n287 B.n286 585
R49 B.n285 B.n116 585
R50 B.n284 B.n283 585
R51 B.n282 B.n117 585
R52 B.n280 B.n279 585
R53 B.n278 B.n120 585
R54 B.n277 B.n276 585
R55 B.n275 B.n121 585
R56 B.n274 B.n273 585
R57 B.n272 B.n122 585
R58 B.n271 B.n270 585
R59 B.n269 B.n123 585
R60 B.n268 B.n267 585
R61 B.n266 B.n124 585
R62 B.n265 B.n264 585
R63 B.n260 B.n125 585
R64 B.n259 B.n258 585
R65 B.n257 B.n126 585
R66 B.n256 B.n255 585
R67 B.n254 B.n127 585
R68 B.n253 B.n252 585
R69 B.n251 B.n128 585
R70 B.n250 B.n249 585
R71 B.n248 B.n129 585
R72 B.n247 B.n246 585
R73 B.n245 B.n130 585
R74 B.n244 B.n243 585
R75 B.n242 B.n131 585
R76 B.n241 B.n240 585
R77 B.n239 B.n132 585
R78 B.n238 B.n237 585
R79 B.n236 B.n133 585
R80 B.n235 B.n234 585
R81 B.n233 B.n134 585
R82 B.n232 B.n231 585
R83 B.n230 B.n135 585
R84 B.n229 B.n228 585
R85 B.n227 B.n136 585
R86 B.n226 B.n225 585
R87 B.n224 B.n137 585
R88 B.n223 B.n222 585
R89 B.n221 B.n138 585
R90 B.n220 B.n219 585
R91 B.n218 B.n139 585
R92 B.n217 B.n216 585
R93 B.n215 B.n140 585
R94 B.n214 B.n213 585
R95 B.n212 B.n141 585
R96 B.n211 B.n210 585
R97 B.n209 B.n142 585
R98 B.n208 B.n207 585
R99 B.n206 B.n143 585
R100 B.n205 B.n204 585
R101 B.n203 B.n144 585
R102 B.n202 B.n201 585
R103 B.n200 B.n145 585
R104 B.n199 B.n198 585
R105 B.n197 B.n146 585
R106 B.n196 B.n195 585
R107 B.n194 B.n147 585
R108 B.n193 B.n192 585
R109 B.n191 B.n148 585
R110 B.n190 B.n189 585
R111 B.n188 B.n149 585
R112 B.n187 B.n186 585
R113 B.n185 B.n150 585
R114 B.n360 B.n91 585
R115 B.n362 B.n361 585
R116 B.n363 B.n90 585
R117 B.n365 B.n364 585
R118 B.n366 B.n89 585
R119 B.n368 B.n367 585
R120 B.n369 B.n88 585
R121 B.n371 B.n370 585
R122 B.n372 B.n87 585
R123 B.n374 B.n373 585
R124 B.n375 B.n86 585
R125 B.n377 B.n376 585
R126 B.n378 B.n85 585
R127 B.n380 B.n379 585
R128 B.n381 B.n84 585
R129 B.n383 B.n382 585
R130 B.n384 B.n83 585
R131 B.n386 B.n385 585
R132 B.n387 B.n82 585
R133 B.n389 B.n388 585
R134 B.n390 B.n81 585
R135 B.n392 B.n391 585
R136 B.n393 B.n80 585
R137 B.n395 B.n394 585
R138 B.n396 B.n79 585
R139 B.n398 B.n397 585
R140 B.n399 B.n78 585
R141 B.n401 B.n400 585
R142 B.n402 B.n77 585
R143 B.n404 B.n403 585
R144 B.n405 B.n76 585
R145 B.n407 B.n406 585
R146 B.n408 B.n75 585
R147 B.n410 B.n409 585
R148 B.n411 B.n74 585
R149 B.n413 B.n412 585
R150 B.n414 B.n73 585
R151 B.n416 B.n415 585
R152 B.n588 B.n11 585
R153 B.n587 B.n586 585
R154 B.n585 B.n12 585
R155 B.n584 B.n583 585
R156 B.n582 B.n13 585
R157 B.n581 B.n580 585
R158 B.n579 B.n14 585
R159 B.n578 B.n577 585
R160 B.n576 B.n15 585
R161 B.n575 B.n574 585
R162 B.n573 B.n16 585
R163 B.n572 B.n571 585
R164 B.n570 B.n17 585
R165 B.n569 B.n568 585
R166 B.n567 B.n18 585
R167 B.n566 B.n565 585
R168 B.n564 B.n19 585
R169 B.n563 B.n562 585
R170 B.n561 B.n20 585
R171 B.n560 B.n559 585
R172 B.n558 B.n21 585
R173 B.n557 B.n556 585
R174 B.n555 B.n22 585
R175 B.n554 B.n553 585
R176 B.n552 B.n23 585
R177 B.n551 B.n550 585
R178 B.n549 B.n24 585
R179 B.n548 B.n547 585
R180 B.n546 B.n25 585
R181 B.n545 B.n544 585
R182 B.n543 B.n26 585
R183 B.n542 B.n541 585
R184 B.n540 B.n27 585
R185 B.n539 B.n538 585
R186 B.n537 B.n28 585
R187 B.n536 B.n535 585
R188 B.n534 B.n29 585
R189 B.n533 B.n532 585
R190 B.n531 B.n30 585
R191 B.n530 B.n529 585
R192 B.n528 B.n31 585
R193 B.n527 B.n526 585
R194 B.n525 B.n32 585
R195 B.n524 B.n523 585
R196 B.n522 B.n33 585
R197 B.n521 B.n520 585
R198 B.n519 B.n34 585
R199 B.n518 B.n517 585
R200 B.n516 B.n35 585
R201 B.n515 B.n514 585
R202 B.n513 B.n36 585
R203 B.n512 B.n511 585
R204 B.n509 B.n37 585
R205 B.n508 B.n507 585
R206 B.n506 B.n40 585
R207 B.n505 B.n504 585
R208 B.n503 B.n41 585
R209 B.n502 B.n501 585
R210 B.n500 B.n42 585
R211 B.n499 B.n498 585
R212 B.n497 B.n43 585
R213 B.n496 B.n495 585
R214 B.n494 B.n493 585
R215 B.n492 B.n47 585
R216 B.n491 B.n490 585
R217 B.n489 B.n48 585
R218 B.n488 B.n487 585
R219 B.n486 B.n49 585
R220 B.n485 B.n484 585
R221 B.n483 B.n50 585
R222 B.n482 B.n481 585
R223 B.n480 B.n51 585
R224 B.n479 B.n478 585
R225 B.n477 B.n52 585
R226 B.n476 B.n475 585
R227 B.n474 B.n53 585
R228 B.n473 B.n472 585
R229 B.n471 B.n54 585
R230 B.n470 B.n469 585
R231 B.n468 B.n55 585
R232 B.n467 B.n466 585
R233 B.n465 B.n56 585
R234 B.n464 B.n463 585
R235 B.n462 B.n57 585
R236 B.n461 B.n460 585
R237 B.n459 B.n58 585
R238 B.n458 B.n457 585
R239 B.n456 B.n59 585
R240 B.n455 B.n454 585
R241 B.n453 B.n60 585
R242 B.n452 B.n451 585
R243 B.n450 B.n61 585
R244 B.n449 B.n448 585
R245 B.n447 B.n62 585
R246 B.n446 B.n445 585
R247 B.n444 B.n63 585
R248 B.n443 B.n442 585
R249 B.n441 B.n64 585
R250 B.n440 B.n439 585
R251 B.n438 B.n65 585
R252 B.n437 B.n436 585
R253 B.n435 B.n66 585
R254 B.n434 B.n433 585
R255 B.n432 B.n67 585
R256 B.n431 B.n430 585
R257 B.n429 B.n68 585
R258 B.n428 B.n427 585
R259 B.n426 B.n69 585
R260 B.n425 B.n424 585
R261 B.n423 B.n70 585
R262 B.n422 B.n421 585
R263 B.n420 B.n71 585
R264 B.n419 B.n418 585
R265 B.n417 B.n72 585
R266 B.n590 B.n589 585
R267 B.n591 B.n10 585
R268 B.n593 B.n592 585
R269 B.n594 B.n9 585
R270 B.n596 B.n595 585
R271 B.n597 B.n8 585
R272 B.n599 B.n598 585
R273 B.n600 B.n7 585
R274 B.n602 B.n601 585
R275 B.n603 B.n6 585
R276 B.n605 B.n604 585
R277 B.n606 B.n5 585
R278 B.n608 B.n607 585
R279 B.n609 B.n4 585
R280 B.n611 B.n610 585
R281 B.n612 B.n3 585
R282 B.n614 B.n613 585
R283 B.n615 B.n0 585
R284 B.n2 B.n1 585
R285 B.n160 B.n159 585
R286 B.n161 B.n158 585
R287 B.n163 B.n162 585
R288 B.n164 B.n157 585
R289 B.n166 B.n165 585
R290 B.n167 B.n156 585
R291 B.n169 B.n168 585
R292 B.n170 B.n155 585
R293 B.n172 B.n171 585
R294 B.n173 B.n154 585
R295 B.n175 B.n174 585
R296 B.n176 B.n153 585
R297 B.n178 B.n177 585
R298 B.n179 B.n152 585
R299 B.n181 B.n180 585
R300 B.n182 B.n151 585
R301 B.n184 B.n183 585
R302 B.n185 B.n184 530.939
R303 B.n358 B.n91 530.939
R304 B.n417 B.n416 530.939
R305 B.n590 B.n11 530.939
R306 B.n118 B.t7 475.75
R307 B.n44 B.t2 475.75
R308 B.n261 B.t10 475.75
R309 B.n38 B.t5 475.75
R310 B.n261 B.t9 463.125
R311 B.n118 B.t6 463.125
R312 B.n44 B.t0 463.125
R313 B.n38 B.t3 463.125
R314 B.n119 B.t8 441.036
R315 B.n45 B.t1 441.036
R316 B.n262 B.t11 441.034
R317 B.n39 B.t4 441.034
R318 B.n617 B.n616 256.663
R319 B.n616 B.n615 235.042
R320 B.n616 B.n2 235.042
R321 B.n186 B.n185 163.367
R322 B.n186 B.n149 163.367
R323 B.n190 B.n149 163.367
R324 B.n191 B.n190 163.367
R325 B.n192 B.n191 163.367
R326 B.n192 B.n147 163.367
R327 B.n196 B.n147 163.367
R328 B.n197 B.n196 163.367
R329 B.n198 B.n197 163.367
R330 B.n198 B.n145 163.367
R331 B.n202 B.n145 163.367
R332 B.n203 B.n202 163.367
R333 B.n204 B.n203 163.367
R334 B.n204 B.n143 163.367
R335 B.n208 B.n143 163.367
R336 B.n209 B.n208 163.367
R337 B.n210 B.n209 163.367
R338 B.n210 B.n141 163.367
R339 B.n214 B.n141 163.367
R340 B.n215 B.n214 163.367
R341 B.n216 B.n215 163.367
R342 B.n216 B.n139 163.367
R343 B.n220 B.n139 163.367
R344 B.n221 B.n220 163.367
R345 B.n222 B.n221 163.367
R346 B.n222 B.n137 163.367
R347 B.n226 B.n137 163.367
R348 B.n227 B.n226 163.367
R349 B.n228 B.n227 163.367
R350 B.n228 B.n135 163.367
R351 B.n232 B.n135 163.367
R352 B.n233 B.n232 163.367
R353 B.n234 B.n233 163.367
R354 B.n234 B.n133 163.367
R355 B.n238 B.n133 163.367
R356 B.n239 B.n238 163.367
R357 B.n240 B.n239 163.367
R358 B.n240 B.n131 163.367
R359 B.n244 B.n131 163.367
R360 B.n245 B.n244 163.367
R361 B.n246 B.n245 163.367
R362 B.n246 B.n129 163.367
R363 B.n250 B.n129 163.367
R364 B.n251 B.n250 163.367
R365 B.n252 B.n251 163.367
R366 B.n252 B.n127 163.367
R367 B.n256 B.n127 163.367
R368 B.n257 B.n256 163.367
R369 B.n258 B.n257 163.367
R370 B.n258 B.n125 163.367
R371 B.n265 B.n125 163.367
R372 B.n266 B.n265 163.367
R373 B.n267 B.n266 163.367
R374 B.n267 B.n123 163.367
R375 B.n271 B.n123 163.367
R376 B.n272 B.n271 163.367
R377 B.n273 B.n272 163.367
R378 B.n273 B.n121 163.367
R379 B.n277 B.n121 163.367
R380 B.n278 B.n277 163.367
R381 B.n279 B.n278 163.367
R382 B.n279 B.n117 163.367
R383 B.n284 B.n117 163.367
R384 B.n285 B.n284 163.367
R385 B.n286 B.n285 163.367
R386 B.n286 B.n115 163.367
R387 B.n290 B.n115 163.367
R388 B.n291 B.n290 163.367
R389 B.n292 B.n291 163.367
R390 B.n292 B.n113 163.367
R391 B.n296 B.n113 163.367
R392 B.n297 B.n296 163.367
R393 B.n298 B.n297 163.367
R394 B.n298 B.n111 163.367
R395 B.n302 B.n111 163.367
R396 B.n303 B.n302 163.367
R397 B.n304 B.n303 163.367
R398 B.n304 B.n109 163.367
R399 B.n308 B.n109 163.367
R400 B.n309 B.n308 163.367
R401 B.n310 B.n309 163.367
R402 B.n310 B.n107 163.367
R403 B.n314 B.n107 163.367
R404 B.n315 B.n314 163.367
R405 B.n316 B.n315 163.367
R406 B.n316 B.n105 163.367
R407 B.n320 B.n105 163.367
R408 B.n321 B.n320 163.367
R409 B.n322 B.n321 163.367
R410 B.n322 B.n103 163.367
R411 B.n326 B.n103 163.367
R412 B.n327 B.n326 163.367
R413 B.n328 B.n327 163.367
R414 B.n328 B.n101 163.367
R415 B.n332 B.n101 163.367
R416 B.n333 B.n332 163.367
R417 B.n334 B.n333 163.367
R418 B.n334 B.n99 163.367
R419 B.n338 B.n99 163.367
R420 B.n339 B.n338 163.367
R421 B.n340 B.n339 163.367
R422 B.n340 B.n97 163.367
R423 B.n344 B.n97 163.367
R424 B.n345 B.n344 163.367
R425 B.n346 B.n345 163.367
R426 B.n346 B.n95 163.367
R427 B.n350 B.n95 163.367
R428 B.n351 B.n350 163.367
R429 B.n352 B.n351 163.367
R430 B.n352 B.n93 163.367
R431 B.n356 B.n93 163.367
R432 B.n357 B.n356 163.367
R433 B.n358 B.n357 163.367
R434 B.n416 B.n73 163.367
R435 B.n412 B.n73 163.367
R436 B.n412 B.n411 163.367
R437 B.n411 B.n410 163.367
R438 B.n410 B.n75 163.367
R439 B.n406 B.n75 163.367
R440 B.n406 B.n405 163.367
R441 B.n405 B.n404 163.367
R442 B.n404 B.n77 163.367
R443 B.n400 B.n77 163.367
R444 B.n400 B.n399 163.367
R445 B.n399 B.n398 163.367
R446 B.n398 B.n79 163.367
R447 B.n394 B.n79 163.367
R448 B.n394 B.n393 163.367
R449 B.n393 B.n392 163.367
R450 B.n392 B.n81 163.367
R451 B.n388 B.n81 163.367
R452 B.n388 B.n387 163.367
R453 B.n387 B.n386 163.367
R454 B.n386 B.n83 163.367
R455 B.n382 B.n83 163.367
R456 B.n382 B.n381 163.367
R457 B.n381 B.n380 163.367
R458 B.n380 B.n85 163.367
R459 B.n376 B.n85 163.367
R460 B.n376 B.n375 163.367
R461 B.n375 B.n374 163.367
R462 B.n374 B.n87 163.367
R463 B.n370 B.n87 163.367
R464 B.n370 B.n369 163.367
R465 B.n369 B.n368 163.367
R466 B.n368 B.n89 163.367
R467 B.n364 B.n89 163.367
R468 B.n364 B.n363 163.367
R469 B.n363 B.n362 163.367
R470 B.n362 B.n91 163.367
R471 B.n586 B.n11 163.367
R472 B.n586 B.n585 163.367
R473 B.n585 B.n584 163.367
R474 B.n584 B.n13 163.367
R475 B.n580 B.n13 163.367
R476 B.n580 B.n579 163.367
R477 B.n579 B.n578 163.367
R478 B.n578 B.n15 163.367
R479 B.n574 B.n15 163.367
R480 B.n574 B.n573 163.367
R481 B.n573 B.n572 163.367
R482 B.n572 B.n17 163.367
R483 B.n568 B.n17 163.367
R484 B.n568 B.n567 163.367
R485 B.n567 B.n566 163.367
R486 B.n566 B.n19 163.367
R487 B.n562 B.n19 163.367
R488 B.n562 B.n561 163.367
R489 B.n561 B.n560 163.367
R490 B.n560 B.n21 163.367
R491 B.n556 B.n21 163.367
R492 B.n556 B.n555 163.367
R493 B.n555 B.n554 163.367
R494 B.n554 B.n23 163.367
R495 B.n550 B.n23 163.367
R496 B.n550 B.n549 163.367
R497 B.n549 B.n548 163.367
R498 B.n548 B.n25 163.367
R499 B.n544 B.n25 163.367
R500 B.n544 B.n543 163.367
R501 B.n543 B.n542 163.367
R502 B.n542 B.n27 163.367
R503 B.n538 B.n27 163.367
R504 B.n538 B.n537 163.367
R505 B.n537 B.n536 163.367
R506 B.n536 B.n29 163.367
R507 B.n532 B.n29 163.367
R508 B.n532 B.n531 163.367
R509 B.n531 B.n530 163.367
R510 B.n530 B.n31 163.367
R511 B.n526 B.n31 163.367
R512 B.n526 B.n525 163.367
R513 B.n525 B.n524 163.367
R514 B.n524 B.n33 163.367
R515 B.n520 B.n33 163.367
R516 B.n520 B.n519 163.367
R517 B.n519 B.n518 163.367
R518 B.n518 B.n35 163.367
R519 B.n514 B.n35 163.367
R520 B.n514 B.n513 163.367
R521 B.n513 B.n512 163.367
R522 B.n512 B.n37 163.367
R523 B.n507 B.n37 163.367
R524 B.n507 B.n506 163.367
R525 B.n506 B.n505 163.367
R526 B.n505 B.n41 163.367
R527 B.n501 B.n41 163.367
R528 B.n501 B.n500 163.367
R529 B.n500 B.n499 163.367
R530 B.n499 B.n43 163.367
R531 B.n495 B.n43 163.367
R532 B.n495 B.n494 163.367
R533 B.n494 B.n47 163.367
R534 B.n490 B.n47 163.367
R535 B.n490 B.n489 163.367
R536 B.n489 B.n488 163.367
R537 B.n488 B.n49 163.367
R538 B.n484 B.n49 163.367
R539 B.n484 B.n483 163.367
R540 B.n483 B.n482 163.367
R541 B.n482 B.n51 163.367
R542 B.n478 B.n51 163.367
R543 B.n478 B.n477 163.367
R544 B.n477 B.n476 163.367
R545 B.n476 B.n53 163.367
R546 B.n472 B.n53 163.367
R547 B.n472 B.n471 163.367
R548 B.n471 B.n470 163.367
R549 B.n470 B.n55 163.367
R550 B.n466 B.n55 163.367
R551 B.n466 B.n465 163.367
R552 B.n465 B.n464 163.367
R553 B.n464 B.n57 163.367
R554 B.n460 B.n57 163.367
R555 B.n460 B.n459 163.367
R556 B.n459 B.n458 163.367
R557 B.n458 B.n59 163.367
R558 B.n454 B.n59 163.367
R559 B.n454 B.n453 163.367
R560 B.n453 B.n452 163.367
R561 B.n452 B.n61 163.367
R562 B.n448 B.n61 163.367
R563 B.n448 B.n447 163.367
R564 B.n447 B.n446 163.367
R565 B.n446 B.n63 163.367
R566 B.n442 B.n63 163.367
R567 B.n442 B.n441 163.367
R568 B.n441 B.n440 163.367
R569 B.n440 B.n65 163.367
R570 B.n436 B.n65 163.367
R571 B.n436 B.n435 163.367
R572 B.n435 B.n434 163.367
R573 B.n434 B.n67 163.367
R574 B.n430 B.n67 163.367
R575 B.n430 B.n429 163.367
R576 B.n429 B.n428 163.367
R577 B.n428 B.n69 163.367
R578 B.n424 B.n69 163.367
R579 B.n424 B.n423 163.367
R580 B.n423 B.n422 163.367
R581 B.n422 B.n71 163.367
R582 B.n418 B.n71 163.367
R583 B.n418 B.n417 163.367
R584 B.n591 B.n590 163.367
R585 B.n592 B.n591 163.367
R586 B.n592 B.n9 163.367
R587 B.n596 B.n9 163.367
R588 B.n597 B.n596 163.367
R589 B.n598 B.n597 163.367
R590 B.n598 B.n7 163.367
R591 B.n602 B.n7 163.367
R592 B.n603 B.n602 163.367
R593 B.n604 B.n603 163.367
R594 B.n604 B.n5 163.367
R595 B.n608 B.n5 163.367
R596 B.n609 B.n608 163.367
R597 B.n610 B.n609 163.367
R598 B.n610 B.n3 163.367
R599 B.n614 B.n3 163.367
R600 B.n615 B.n614 163.367
R601 B.n160 B.n2 163.367
R602 B.n161 B.n160 163.367
R603 B.n162 B.n161 163.367
R604 B.n162 B.n157 163.367
R605 B.n166 B.n157 163.367
R606 B.n167 B.n166 163.367
R607 B.n168 B.n167 163.367
R608 B.n168 B.n155 163.367
R609 B.n172 B.n155 163.367
R610 B.n173 B.n172 163.367
R611 B.n174 B.n173 163.367
R612 B.n174 B.n153 163.367
R613 B.n178 B.n153 163.367
R614 B.n179 B.n178 163.367
R615 B.n180 B.n179 163.367
R616 B.n180 B.n151 163.367
R617 B.n184 B.n151 163.367
R618 B.n263 B.n262 59.5399
R619 B.n281 B.n119 59.5399
R620 B.n46 B.n45 59.5399
R621 B.n510 B.n39 59.5399
R622 B.n262 B.n261 34.7157
R623 B.n119 B.n118 34.7157
R624 B.n45 B.n44 34.7157
R625 B.n39 B.n38 34.7157
R626 B.n589 B.n588 34.4981
R627 B.n415 B.n72 34.4981
R628 B.n360 B.n359 34.4981
R629 B.n183 B.n150 34.4981
R630 B B.n617 18.0485
R631 B.n589 B.n10 10.6151
R632 B.n593 B.n10 10.6151
R633 B.n594 B.n593 10.6151
R634 B.n595 B.n594 10.6151
R635 B.n595 B.n8 10.6151
R636 B.n599 B.n8 10.6151
R637 B.n600 B.n599 10.6151
R638 B.n601 B.n600 10.6151
R639 B.n601 B.n6 10.6151
R640 B.n605 B.n6 10.6151
R641 B.n606 B.n605 10.6151
R642 B.n607 B.n606 10.6151
R643 B.n607 B.n4 10.6151
R644 B.n611 B.n4 10.6151
R645 B.n612 B.n611 10.6151
R646 B.n613 B.n612 10.6151
R647 B.n613 B.n0 10.6151
R648 B.n588 B.n587 10.6151
R649 B.n587 B.n12 10.6151
R650 B.n583 B.n12 10.6151
R651 B.n583 B.n582 10.6151
R652 B.n582 B.n581 10.6151
R653 B.n581 B.n14 10.6151
R654 B.n577 B.n14 10.6151
R655 B.n577 B.n576 10.6151
R656 B.n576 B.n575 10.6151
R657 B.n575 B.n16 10.6151
R658 B.n571 B.n16 10.6151
R659 B.n571 B.n570 10.6151
R660 B.n570 B.n569 10.6151
R661 B.n569 B.n18 10.6151
R662 B.n565 B.n18 10.6151
R663 B.n565 B.n564 10.6151
R664 B.n564 B.n563 10.6151
R665 B.n563 B.n20 10.6151
R666 B.n559 B.n20 10.6151
R667 B.n559 B.n558 10.6151
R668 B.n558 B.n557 10.6151
R669 B.n557 B.n22 10.6151
R670 B.n553 B.n22 10.6151
R671 B.n553 B.n552 10.6151
R672 B.n552 B.n551 10.6151
R673 B.n551 B.n24 10.6151
R674 B.n547 B.n24 10.6151
R675 B.n547 B.n546 10.6151
R676 B.n546 B.n545 10.6151
R677 B.n545 B.n26 10.6151
R678 B.n541 B.n26 10.6151
R679 B.n541 B.n540 10.6151
R680 B.n540 B.n539 10.6151
R681 B.n539 B.n28 10.6151
R682 B.n535 B.n28 10.6151
R683 B.n535 B.n534 10.6151
R684 B.n534 B.n533 10.6151
R685 B.n533 B.n30 10.6151
R686 B.n529 B.n30 10.6151
R687 B.n529 B.n528 10.6151
R688 B.n528 B.n527 10.6151
R689 B.n527 B.n32 10.6151
R690 B.n523 B.n32 10.6151
R691 B.n523 B.n522 10.6151
R692 B.n522 B.n521 10.6151
R693 B.n521 B.n34 10.6151
R694 B.n517 B.n34 10.6151
R695 B.n517 B.n516 10.6151
R696 B.n516 B.n515 10.6151
R697 B.n515 B.n36 10.6151
R698 B.n511 B.n36 10.6151
R699 B.n509 B.n508 10.6151
R700 B.n508 B.n40 10.6151
R701 B.n504 B.n40 10.6151
R702 B.n504 B.n503 10.6151
R703 B.n503 B.n502 10.6151
R704 B.n502 B.n42 10.6151
R705 B.n498 B.n42 10.6151
R706 B.n498 B.n497 10.6151
R707 B.n497 B.n496 10.6151
R708 B.n493 B.n492 10.6151
R709 B.n492 B.n491 10.6151
R710 B.n491 B.n48 10.6151
R711 B.n487 B.n48 10.6151
R712 B.n487 B.n486 10.6151
R713 B.n486 B.n485 10.6151
R714 B.n485 B.n50 10.6151
R715 B.n481 B.n50 10.6151
R716 B.n481 B.n480 10.6151
R717 B.n480 B.n479 10.6151
R718 B.n479 B.n52 10.6151
R719 B.n475 B.n52 10.6151
R720 B.n475 B.n474 10.6151
R721 B.n474 B.n473 10.6151
R722 B.n473 B.n54 10.6151
R723 B.n469 B.n54 10.6151
R724 B.n469 B.n468 10.6151
R725 B.n468 B.n467 10.6151
R726 B.n467 B.n56 10.6151
R727 B.n463 B.n56 10.6151
R728 B.n463 B.n462 10.6151
R729 B.n462 B.n461 10.6151
R730 B.n461 B.n58 10.6151
R731 B.n457 B.n58 10.6151
R732 B.n457 B.n456 10.6151
R733 B.n456 B.n455 10.6151
R734 B.n455 B.n60 10.6151
R735 B.n451 B.n60 10.6151
R736 B.n451 B.n450 10.6151
R737 B.n450 B.n449 10.6151
R738 B.n449 B.n62 10.6151
R739 B.n445 B.n62 10.6151
R740 B.n445 B.n444 10.6151
R741 B.n444 B.n443 10.6151
R742 B.n443 B.n64 10.6151
R743 B.n439 B.n64 10.6151
R744 B.n439 B.n438 10.6151
R745 B.n438 B.n437 10.6151
R746 B.n437 B.n66 10.6151
R747 B.n433 B.n66 10.6151
R748 B.n433 B.n432 10.6151
R749 B.n432 B.n431 10.6151
R750 B.n431 B.n68 10.6151
R751 B.n427 B.n68 10.6151
R752 B.n427 B.n426 10.6151
R753 B.n426 B.n425 10.6151
R754 B.n425 B.n70 10.6151
R755 B.n421 B.n70 10.6151
R756 B.n421 B.n420 10.6151
R757 B.n420 B.n419 10.6151
R758 B.n419 B.n72 10.6151
R759 B.n415 B.n414 10.6151
R760 B.n414 B.n413 10.6151
R761 B.n413 B.n74 10.6151
R762 B.n409 B.n74 10.6151
R763 B.n409 B.n408 10.6151
R764 B.n408 B.n407 10.6151
R765 B.n407 B.n76 10.6151
R766 B.n403 B.n76 10.6151
R767 B.n403 B.n402 10.6151
R768 B.n402 B.n401 10.6151
R769 B.n401 B.n78 10.6151
R770 B.n397 B.n78 10.6151
R771 B.n397 B.n396 10.6151
R772 B.n396 B.n395 10.6151
R773 B.n395 B.n80 10.6151
R774 B.n391 B.n80 10.6151
R775 B.n391 B.n390 10.6151
R776 B.n390 B.n389 10.6151
R777 B.n389 B.n82 10.6151
R778 B.n385 B.n82 10.6151
R779 B.n385 B.n384 10.6151
R780 B.n384 B.n383 10.6151
R781 B.n383 B.n84 10.6151
R782 B.n379 B.n84 10.6151
R783 B.n379 B.n378 10.6151
R784 B.n378 B.n377 10.6151
R785 B.n377 B.n86 10.6151
R786 B.n373 B.n86 10.6151
R787 B.n373 B.n372 10.6151
R788 B.n372 B.n371 10.6151
R789 B.n371 B.n88 10.6151
R790 B.n367 B.n88 10.6151
R791 B.n367 B.n366 10.6151
R792 B.n366 B.n365 10.6151
R793 B.n365 B.n90 10.6151
R794 B.n361 B.n90 10.6151
R795 B.n361 B.n360 10.6151
R796 B.n159 B.n1 10.6151
R797 B.n159 B.n158 10.6151
R798 B.n163 B.n158 10.6151
R799 B.n164 B.n163 10.6151
R800 B.n165 B.n164 10.6151
R801 B.n165 B.n156 10.6151
R802 B.n169 B.n156 10.6151
R803 B.n170 B.n169 10.6151
R804 B.n171 B.n170 10.6151
R805 B.n171 B.n154 10.6151
R806 B.n175 B.n154 10.6151
R807 B.n176 B.n175 10.6151
R808 B.n177 B.n176 10.6151
R809 B.n177 B.n152 10.6151
R810 B.n181 B.n152 10.6151
R811 B.n182 B.n181 10.6151
R812 B.n183 B.n182 10.6151
R813 B.n187 B.n150 10.6151
R814 B.n188 B.n187 10.6151
R815 B.n189 B.n188 10.6151
R816 B.n189 B.n148 10.6151
R817 B.n193 B.n148 10.6151
R818 B.n194 B.n193 10.6151
R819 B.n195 B.n194 10.6151
R820 B.n195 B.n146 10.6151
R821 B.n199 B.n146 10.6151
R822 B.n200 B.n199 10.6151
R823 B.n201 B.n200 10.6151
R824 B.n201 B.n144 10.6151
R825 B.n205 B.n144 10.6151
R826 B.n206 B.n205 10.6151
R827 B.n207 B.n206 10.6151
R828 B.n207 B.n142 10.6151
R829 B.n211 B.n142 10.6151
R830 B.n212 B.n211 10.6151
R831 B.n213 B.n212 10.6151
R832 B.n213 B.n140 10.6151
R833 B.n217 B.n140 10.6151
R834 B.n218 B.n217 10.6151
R835 B.n219 B.n218 10.6151
R836 B.n219 B.n138 10.6151
R837 B.n223 B.n138 10.6151
R838 B.n224 B.n223 10.6151
R839 B.n225 B.n224 10.6151
R840 B.n225 B.n136 10.6151
R841 B.n229 B.n136 10.6151
R842 B.n230 B.n229 10.6151
R843 B.n231 B.n230 10.6151
R844 B.n231 B.n134 10.6151
R845 B.n235 B.n134 10.6151
R846 B.n236 B.n235 10.6151
R847 B.n237 B.n236 10.6151
R848 B.n237 B.n132 10.6151
R849 B.n241 B.n132 10.6151
R850 B.n242 B.n241 10.6151
R851 B.n243 B.n242 10.6151
R852 B.n243 B.n130 10.6151
R853 B.n247 B.n130 10.6151
R854 B.n248 B.n247 10.6151
R855 B.n249 B.n248 10.6151
R856 B.n249 B.n128 10.6151
R857 B.n253 B.n128 10.6151
R858 B.n254 B.n253 10.6151
R859 B.n255 B.n254 10.6151
R860 B.n255 B.n126 10.6151
R861 B.n259 B.n126 10.6151
R862 B.n260 B.n259 10.6151
R863 B.n264 B.n260 10.6151
R864 B.n268 B.n124 10.6151
R865 B.n269 B.n268 10.6151
R866 B.n270 B.n269 10.6151
R867 B.n270 B.n122 10.6151
R868 B.n274 B.n122 10.6151
R869 B.n275 B.n274 10.6151
R870 B.n276 B.n275 10.6151
R871 B.n276 B.n120 10.6151
R872 B.n280 B.n120 10.6151
R873 B.n283 B.n282 10.6151
R874 B.n283 B.n116 10.6151
R875 B.n287 B.n116 10.6151
R876 B.n288 B.n287 10.6151
R877 B.n289 B.n288 10.6151
R878 B.n289 B.n114 10.6151
R879 B.n293 B.n114 10.6151
R880 B.n294 B.n293 10.6151
R881 B.n295 B.n294 10.6151
R882 B.n295 B.n112 10.6151
R883 B.n299 B.n112 10.6151
R884 B.n300 B.n299 10.6151
R885 B.n301 B.n300 10.6151
R886 B.n301 B.n110 10.6151
R887 B.n305 B.n110 10.6151
R888 B.n306 B.n305 10.6151
R889 B.n307 B.n306 10.6151
R890 B.n307 B.n108 10.6151
R891 B.n311 B.n108 10.6151
R892 B.n312 B.n311 10.6151
R893 B.n313 B.n312 10.6151
R894 B.n313 B.n106 10.6151
R895 B.n317 B.n106 10.6151
R896 B.n318 B.n317 10.6151
R897 B.n319 B.n318 10.6151
R898 B.n319 B.n104 10.6151
R899 B.n323 B.n104 10.6151
R900 B.n324 B.n323 10.6151
R901 B.n325 B.n324 10.6151
R902 B.n325 B.n102 10.6151
R903 B.n329 B.n102 10.6151
R904 B.n330 B.n329 10.6151
R905 B.n331 B.n330 10.6151
R906 B.n331 B.n100 10.6151
R907 B.n335 B.n100 10.6151
R908 B.n336 B.n335 10.6151
R909 B.n337 B.n336 10.6151
R910 B.n337 B.n98 10.6151
R911 B.n341 B.n98 10.6151
R912 B.n342 B.n341 10.6151
R913 B.n343 B.n342 10.6151
R914 B.n343 B.n96 10.6151
R915 B.n347 B.n96 10.6151
R916 B.n348 B.n347 10.6151
R917 B.n349 B.n348 10.6151
R918 B.n349 B.n94 10.6151
R919 B.n353 B.n94 10.6151
R920 B.n354 B.n353 10.6151
R921 B.n355 B.n354 10.6151
R922 B.n355 B.n92 10.6151
R923 B.n359 B.n92 10.6151
R924 B.n511 B.n510 9.36635
R925 B.n493 B.n46 9.36635
R926 B.n264 B.n263 9.36635
R927 B.n282 B.n281 9.36635
R928 B.n617 B.n0 8.11757
R929 B.n617 B.n1 8.11757
R930 B.n510 B.n509 1.24928
R931 B.n496 B.n46 1.24928
R932 B.n263 B.n124 1.24928
R933 B.n281 B.n280 1.24928
R934 VN VN.t1 410.009
R935 VN VN.t0 365.493
R936 VTAIL.n338 VTAIL.n258 756.745
R937 VTAIL.n80 VTAIL.n0 756.745
R938 VTAIL.n252 VTAIL.n172 756.745
R939 VTAIL.n166 VTAIL.n86 756.745
R940 VTAIL.n287 VTAIL.n286 585
R941 VTAIL.n289 VTAIL.n288 585
R942 VTAIL.n282 VTAIL.n281 585
R943 VTAIL.n295 VTAIL.n294 585
R944 VTAIL.n297 VTAIL.n296 585
R945 VTAIL.n278 VTAIL.n277 585
R946 VTAIL.n304 VTAIL.n303 585
R947 VTAIL.n305 VTAIL.n276 585
R948 VTAIL.n307 VTAIL.n306 585
R949 VTAIL.n274 VTAIL.n273 585
R950 VTAIL.n313 VTAIL.n312 585
R951 VTAIL.n315 VTAIL.n314 585
R952 VTAIL.n270 VTAIL.n269 585
R953 VTAIL.n321 VTAIL.n320 585
R954 VTAIL.n323 VTAIL.n322 585
R955 VTAIL.n266 VTAIL.n265 585
R956 VTAIL.n329 VTAIL.n328 585
R957 VTAIL.n331 VTAIL.n330 585
R958 VTAIL.n262 VTAIL.n261 585
R959 VTAIL.n337 VTAIL.n336 585
R960 VTAIL.n339 VTAIL.n338 585
R961 VTAIL.n29 VTAIL.n28 585
R962 VTAIL.n31 VTAIL.n30 585
R963 VTAIL.n24 VTAIL.n23 585
R964 VTAIL.n37 VTAIL.n36 585
R965 VTAIL.n39 VTAIL.n38 585
R966 VTAIL.n20 VTAIL.n19 585
R967 VTAIL.n46 VTAIL.n45 585
R968 VTAIL.n47 VTAIL.n18 585
R969 VTAIL.n49 VTAIL.n48 585
R970 VTAIL.n16 VTAIL.n15 585
R971 VTAIL.n55 VTAIL.n54 585
R972 VTAIL.n57 VTAIL.n56 585
R973 VTAIL.n12 VTAIL.n11 585
R974 VTAIL.n63 VTAIL.n62 585
R975 VTAIL.n65 VTAIL.n64 585
R976 VTAIL.n8 VTAIL.n7 585
R977 VTAIL.n71 VTAIL.n70 585
R978 VTAIL.n73 VTAIL.n72 585
R979 VTAIL.n4 VTAIL.n3 585
R980 VTAIL.n79 VTAIL.n78 585
R981 VTAIL.n81 VTAIL.n80 585
R982 VTAIL.n253 VTAIL.n252 585
R983 VTAIL.n251 VTAIL.n250 585
R984 VTAIL.n176 VTAIL.n175 585
R985 VTAIL.n245 VTAIL.n244 585
R986 VTAIL.n243 VTAIL.n242 585
R987 VTAIL.n180 VTAIL.n179 585
R988 VTAIL.n237 VTAIL.n236 585
R989 VTAIL.n235 VTAIL.n234 585
R990 VTAIL.n184 VTAIL.n183 585
R991 VTAIL.n229 VTAIL.n228 585
R992 VTAIL.n227 VTAIL.n226 585
R993 VTAIL.n188 VTAIL.n187 585
R994 VTAIL.n192 VTAIL.n190 585
R995 VTAIL.n221 VTAIL.n220 585
R996 VTAIL.n219 VTAIL.n218 585
R997 VTAIL.n194 VTAIL.n193 585
R998 VTAIL.n213 VTAIL.n212 585
R999 VTAIL.n211 VTAIL.n210 585
R1000 VTAIL.n198 VTAIL.n197 585
R1001 VTAIL.n205 VTAIL.n204 585
R1002 VTAIL.n203 VTAIL.n202 585
R1003 VTAIL.n167 VTAIL.n166 585
R1004 VTAIL.n165 VTAIL.n164 585
R1005 VTAIL.n90 VTAIL.n89 585
R1006 VTAIL.n159 VTAIL.n158 585
R1007 VTAIL.n157 VTAIL.n156 585
R1008 VTAIL.n94 VTAIL.n93 585
R1009 VTAIL.n151 VTAIL.n150 585
R1010 VTAIL.n149 VTAIL.n148 585
R1011 VTAIL.n98 VTAIL.n97 585
R1012 VTAIL.n143 VTAIL.n142 585
R1013 VTAIL.n141 VTAIL.n140 585
R1014 VTAIL.n102 VTAIL.n101 585
R1015 VTAIL.n106 VTAIL.n104 585
R1016 VTAIL.n135 VTAIL.n134 585
R1017 VTAIL.n133 VTAIL.n132 585
R1018 VTAIL.n108 VTAIL.n107 585
R1019 VTAIL.n127 VTAIL.n126 585
R1020 VTAIL.n125 VTAIL.n124 585
R1021 VTAIL.n112 VTAIL.n111 585
R1022 VTAIL.n119 VTAIL.n118 585
R1023 VTAIL.n117 VTAIL.n116 585
R1024 VTAIL.n285 VTAIL.t2 329.036
R1025 VTAIL.n27 VTAIL.t3 329.036
R1026 VTAIL.n201 VTAIL.t0 329.036
R1027 VTAIL.n115 VTAIL.t1 329.036
R1028 VTAIL.n288 VTAIL.n287 171.744
R1029 VTAIL.n288 VTAIL.n281 171.744
R1030 VTAIL.n295 VTAIL.n281 171.744
R1031 VTAIL.n296 VTAIL.n295 171.744
R1032 VTAIL.n296 VTAIL.n277 171.744
R1033 VTAIL.n304 VTAIL.n277 171.744
R1034 VTAIL.n305 VTAIL.n304 171.744
R1035 VTAIL.n306 VTAIL.n305 171.744
R1036 VTAIL.n306 VTAIL.n273 171.744
R1037 VTAIL.n313 VTAIL.n273 171.744
R1038 VTAIL.n314 VTAIL.n313 171.744
R1039 VTAIL.n314 VTAIL.n269 171.744
R1040 VTAIL.n321 VTAIL.n269 171.744
R1041 VTAIL.n322 VTAIL.n321 171.744
R1042 VTAIL.n322 VTAIL.n265 171.744
R1043 VTAIL.n329 VTAIL.n265 171.744
R1044 VTAIL.n330 VTAIL.n329 171.744
R1045 VTAIL.n330 VTAIL.n261 171.744
R1046 VTAIL.n337 VTAIL.n261 171.744
R1047 VTAIL.n338 VTAIL.n337 171.744
R1048 VTAIL.n30 VTAIL.n29 171.744
R1049 VTAIL.n30 VTAIL.n23 171.744
R1050 VTAIL.n37 VTAIL.n23 171.744
R1051 VTAIL.n38 VTAIL.n37 171.744
R1052 VTAIL.n38 VTAIL.n19 171.744
R1053 VTAIL.n46 VTAIL.n19 171.744
R1054 VTAIL.n47 VTAIL.n46 171.744
R1055 VTAIL.n48 VTAIL.n47 171.744
R1056 VTAIL.n48 VTAIL.n15 171.744
R1057 VTAIL.n55 VTAIL.n15 171.744
R1058 VTAIL.n56 VTAIL.n55 171.744
R1059 VTAIL.n56 VTAIL.n11 171.744
R1060 VTAIL.n63 VTAIL.n11 171.744
R1061 VTAIL.n64 VTAIL.n63 171.744
R1062 VTAIL.n64 VTAIL.n7 171.744
R1063 VTAIL.n71 VTAIL.n7 171.744
R1064 VTAIL.n72 VTAIL.n71 171.744
R1065 VTAIL.n72 VTAIL.n3 171.744
R1066 VTAIL.n79 VTAIL.n3 171.744
R1067 VTAIL.n80 VTAIL.n79 171.744
R1068 VTAIL.n252 VTAIL.n251 171.744
R1069 VTAIL.n251 VTAIL.n175 171.744
R1070 VTAIL.n244 VTAIL.n175 171.744
R1071 VTAIL.n244 VTAIL.n243 171.744
R1072 VTAIL.n243 VTAIL.n179 171.744
R1073 VTAIL.n236 VTAIL.n179 171.744
R1074 VTAIL.n236 VTAIL.n235 171.744
R1075 VTAIL.n235 VTAIL.n183 171.744
R1076 VTAIL.n228 VTAIL.n183 171.744
R1077 VTAIL.n228 VTAIL.n227 171.744
R1078 VTAIL.n227 VTAIL.n187 171.744
R1079 VTAIL.n192 VTAIL.n187 171.744
R1080 VTAIL.n220 VTAIL.n192 171.744
R1081 VTAIL.n220 VTAIL.n219 171.744
R1082 VTAIL.n219 VTAIL.n193 171.744
R1083 VTAIL.n212 VTAIL.n193 171.744
R1084 VTAIL.n212 VTAIL.n211 171.744
R1085 VTAIL.n211 VTAIL.n197 171.744
R1086 VTAIL.n204 VTAIL.n197 171.744
R1087 VTAIL.n204 VTAIL.n203 171.744
R1088 VTAIL.n166 VTAIL.n165 171.744
R1089 VTAIL.n165 VTAIL.n89 171.744
R1090 VTAIL.n158 VTAIL.n89 171.744
R1091 VTAIL.n158 VTAIL.n157 171.744
R1092 VTAIL.n157 VTAIL.n93 171.744
R1093 VTAIL.n150 VTAIL.n93 171.744
R1094 VTAIL.n150 VTAIL.n149 171.744
R1095 VTAIL.n149 VTAIL.n97 171.744
R1096 VTAIL.n142 VTAIL.n97 171.744
R1097 VTAIL.n142 VTAIL.n141 171.744
R1098 VTAIL.n141 VTAIL.n101 171.744
R1099 VTAIL.n106 VTAIL.n101 171.744
R1100 VTAIL.n134 VTAIL.n106 171.744
R1101 VTAIL.n134 VTAIL.n133 171.744
R1102 VTAIL.n133 VTAIL.n107 171.744
R1103 VTAIL.n126 VTAIL.n107 171.744
R1104 VTAIL.n126 VTAIL.n125 171.744
R1105 VTAIL.n125 VTAIL.n111 171.744
R1106 VTAIL.n118 VTAIL.n111 171.744
R1107 VTAIL.n118 VTAIL.n117 171.744
R1108 VTAIL.n287 VTAIL.t2 85.8723
R1109 VTAIL.n29 VTAIL.t3 85.8723
R1110 VTAIL.n203 VTAIL.t0 85.8723
R1111 VTAIL.n117 VTAIL.t1 85.8723
R1112 VTAIL.n343 VTAIL.n342 30.246
R1113 VTAIL.n85 VTAIL.n84 30.246
R1114 VTAIL.n257 VTAIL.n256 30.246
R1115 VTAIL.n171 VTAIL.n170 30.246
R1116 VTAIL.n171 VTAIL.n85 28.9186
R1117 VTAIL.n343 VTAIL.n257 27.3755
R1118 VTAIL.n307 VTAIL.n274 13.1884
R1119 VTAIL.n49 VTAIL.n16 13.1884
R1120 VTAIL.n190 VTAIL.n188 13.1884
R1121 VTAIL.n104 VTAIL.n102 13.1884
R1122 VTAIL.n308 VTAIL.n276 12.8005
R1123 VTAIL.n312 VTAIL.n311 12.8005
R1124 VTAIL.n50 VTAIL.n18 12.8005
R1125 VTAIL.n54 VTAIL.n53 12.8005
R1126 VTAIL.n226 VTAIL.n225 12.8005
R1127 VTAIL.n222 VTAIL.n221 12.8005
R1128 VTAIL.n140 VTAIL.n139 12.8005
R1129 VTAIL.n136 VTAIL.n135 12.8005
R1130 VTAIL.n303 VTAIL.n302 12.0247
R1131 VTAIL.n315 VTAIL.n272 12.0247
R1132 VTAIL.n45 VTAIL.n44 12.0247
R1133 VTAIL.n57 VTAIL.n14 12.0247
R1134 VTAIL.n229 VTAIL.n186 12.0247
R1135 VTAIL.n218 VTAIL.n191 12.0247
R1136 VTAIL.n143 VTAIL.n100 12.0247
R1137 VTAIL.n132 VTAIL.n105 12.0247
R1138 VTAIL.n301 VTAIL.n278 11.249
R1139 VTAIL.n316 VTAIL.n270 11.249
R1140 VTAIL.n43 VTAIL.n20 11.249
R1141 VTAIL.n58 VTAIL.n12 11.249
R1142 VTAIL.n230 VTAIL.n184 11.249
R1143 VTAIL.n217 VTAIL.n194 11.249
R1144 VTAIL.n144 VTAIL.n98 11.249
R1145 VTAIL.n131 VTAIL.n108 11.249
R1146 VTAIL.n286 VTAIL.n285 10.7239
R1147 VTAIL.n28 VTAIL.n27 10.7239
R1148 VTAIL.n202 VTAIL.n201 10.7239
R1149 VTAIL.n116 VTAIL.n115 10.7239
R1150 VTAIL.n298 VTAIL.n297 10.4732
R1151 VTAIL.n320 VTAIL.n319 10.4732
R1152 VTAIL.n40 VTAIL.n39 10.4732
R1153 VTAIL.n62 VTAIL.n61 10.4732
R1154 VTAIL.n234 VTAIL.n233 10.4732
R1155 VTAIL.n214 VTAIL.n213 10.4732
R1156 VTAIL.n148 VTAIL.n147 10.4732
R1157 VTAIL.n128 VTAIL.n127 10.4732
R1158 VTAIL.n294 VTAIL.n280 9.69747
R1159 VTAIL.n323 VTAIL.n268 9.69747
R1160 VTAIL.n342 VTAIL.n258 9.69747
R1161 VTAIL.n36 VTAIL.n22 9.69747
R1162 VTAIL.n65 VTAIL.n10 9.69747
R1163 VTAIL.n84 VTAIL.n0 9.69747
R1164 VTAIL.n256 VTAIL.n172 9.69747
R1165 VTAIL.n237 VTAIL.n182 9.69747
R1166 VTAIL.n210 VTAIL.n196 9.69747
R1167 VTAIL.n170 VTAIL.n86 9.69747
R1168 VTAIL.n151 VTAIL.n96 9.69747
R1169 VTAIL.n124 VTAIL.n110 9.69747
R1170 VTAIL.n342 VTAIL.n341 9.45567
R1171 VTAIL.n84 VTAIL.n83 9.45567
R1172 VTAIL.n256 VTAIL.n255 9.45567
R1173 VTAIL.n170 VTAIL.n169 9.45567
R1174 VTAIL.n333 VTAIL.n332 9.3005
R1175 VTAIL.n335 VTAIL.n334 9.3005
R1176 VTAIL.n260 VTAIL.n259 9.3005
R1177 VTAIL.n341 VTAIL.n340 9.3005
R1178 VTAIL.n327 VTAIL.n326 9.3005
R1179 VTAIL.n325 VTAIL.n324 9.3005
R1180 VTAIL.n268 VTAIL.n267 9.3005
R1181 VTAIL.n319 VTAIL.n318 9.3005
R1182 VTAIL.n317 VTAIL.n316 9.3005
R1183 VTAIL.n272 VTAIL.n271 9.3005
R1184 VTAIL.n311 VTAIL.n310 9.3005
R1185 VTAIL.n284 VTAIL.n283 9.3005
R1186 VTAIL.n291 VTAIL.n290 9.3005
R1187 VTAIL.n293 VTAIL.n292 9.3005
R1188 VTAIL.n280 VTAIL.n279 9.3005
R1189 VTAIL.n299 VTAIL.n298 9.3005
R1190 VTAIL.n301 VTAIL.n300 9.3005
R1191 VTAIL.n302 VTAIL.n275 9.3005
R1192 VTAIL.n309 VTAIL.n308 9.3005
R1193 VTAIL.n264 VTAIL.n263 9.3005
R1194 VTAIL.n75 VTAIL.n74 9.3005
R1195 VTAIL.n77 VTAIL.n76 9.3005
R1196 VTAIL.n2 VTAIL.n1 9.3005
R1197 VTAIL.n83 VTAIL.n82 9.3005
R1198 VTAIL.n69 VTAIL.n68 9.3005
R1199 VTAIL.n67 VTAIL.n66 9.3005
R1200 VTAIL.n10 VTAIL.n9 9.3005
R1201 VTAIL.n61 VTAIL.n60 9.3005
R1202 VTAIL.n59 VTAIL.n58 9.3005
R1203 VTAIL.n14 VTAIL.n13 9.3005
R1204 VTAIL.n53 VTAIL.n52 9.3005
R1205 VTAIL.n26 VTAIL.n25 9.3005
R1206 VTAIL.n33 VTAIL.n32 9.3005
R1207 VTAIL.n35 VTAIL.n34 9.3005
R1208 VTAIL.n22 VTAIL.n21 9.3005
R1209 VTAIL.n41 VTAIL.n40 9.3005
R1210 VTAIL.n43 VTAIL.n42 9.3005
R1211 VTAIL.n44 VTAIL.n17 9.3005
R1212 VTAIL.n51 VTAIL.n50 9.3005
R1213 VTAIL.n6 VTAIL.n5 9.3005
R1214 VTAIL.n174 VTAIL.n173 9.3005
R1215 VTAIL.n249 VTAIL.n248 9.3005
R1216 VTAIL.n247 VTAIL.n246 9.3005
R1217 VTAIL.n178 VTAIL.n177 9.3005
R1218 VTAIL.n241 VTAIL.n240 9.3005
R1219 VTAIL.n239 VTAIL.n238 9.3005
R1220 VTAIL.n182 VTAIL.n181 9.3005
R1221 VTAIL.n233 VTAIL.n232 9.3005
R1222 VTAIL.n231 VTAIL.n230 9.3005
R1223 VTAIL.n186 VTAIL.n185 9.3005
R1224 VTAIL.n225 VTAIL.n224 9.3005
R1225 VTAIL.n223 VTAIL.n222 9.3005
R1226 VTAIL.n191 VTAIL.n189 9.3005
R1227 VTAIL.n217 VTAIL.n216 9.3005
R1228 VTAIL.n215 VTAIL.n214 9.3005
R1229 VTAIL.n196 VTAIL.n195 9.3005
R1230 VTAIL.n209 VTAIL.n208 9.3005
R1231 VTAIL.n207 VTAIL.n206 9.3005
R1232 VTAIL.n200 VTAIL.n199 9.3005
R1233 VTAIL.n255 VTAIL.n254 9.3005
R1234 VTAIL.n114 VTAIL.n113 9.3005
R1235 VTAIL.n121 VTAIL.n120 9.3005
R1236 VTAIL.n123 VTAIL.n122 9.3005
R1237 VTAIL.n110 VTAIL.n109 9.3005
R1238 VTAIL.n129 VTAIL.n128 9.3005
R1239 VTAIL.n131 VTAIL.n130 9.3005
R1240 VTAIL.n105 VTAIL.n103 9.3005
R1241 VTAIL.n137 VTAIL.n136 9.3005
R1242 VTAIL.n163 VTAIL.n162 9.3005
R1243 VTAIL.n88 VTAIL.n87 9.3005
R1244 VTAIL.n169 VTAIL.n168 9.3005
R1245 VTAIL.n161 VTAIL.n160 9.3005
R1246 VTAIL.n92 VTAIL.n91 9.3005
R1247 VTAIL.n155 VTAIL.n154 9.3005
R1248 VTAIL.n153 VTAIL.n152 9.3005
R1249 VTAIL.n96 VTAIL.n95 9.3005
R1250 VTAIL.n147 VTAIL.n146 9.3005
R1251 VTAIL.n145 VTAIL.n144 9.3005
R1252 VTAIL.n100 VTAIL.n99 9.3005
R1253 VTAIL.n139 VTAIL.n138 9.3005
R1254 VTAIL.n293 VTAIL.n282 8.92171
R1255 VTAIL.n324 VTAIL.n266 8.92171
R1256 VTAIL.n340 VTAIL.n339 8.92171
R1257 VTAIL.n35 VTAIL.n24 8.92171
R1258 VTAIL.n66 VTAIL.n8 8.92171
R1259 VTAIL.n82 VTAIL.n81 8.92171
R1260 VTAIL.n254 VTAIL.n253 8.92171
R1261 VTAIL.n238 VTAIL.n180 8.92171
R1262 VTAIL.n209 VTAIL.n198 8.92171
R1263 VTAIL.n168 VTAIL.n167 8.92171
R1264 VTAIL.n152 VTAIL.n94 8.92171
R1265 VTAIL.n123 VTAIL.n112 8.92171
R1266 VTAIL.n290 VTAIL.n289 8.14595
R1267 VTAIL.n328 VTAIL.n327 8.14595
R1268 VTAIL.n336 VTAIL.n260 8.14595
R1269 VTAIL.n32 VTAIL.n31 8.14595
R1270 VTAIL.n70 VTAIL.n69 8.14595
R1271 VTAIL.n78 VTAIL.n2 8.14595
R1272 VTAIL.n250 VTAIL.n174 8.14595
R1273 VTAIL.n242 VTAIL.n241 8.14595
R1274 VTAIL.n206 VTAIL.n205 8.14595
R1275 VTAIL.n164 VTAIL.n88 8.14595
R1276 VTAIL.n156 VTAIL.n155 8.14595
R1277 VTAIL.n120 VTAIL.n119 8.14595
R1278 VTAIL.n286 VTAIL.n284 7.3702
R1279 VTAIL.n331 VTAIL.n264 7.3702
R1280 VTAIL.n335 VTAIL.n262 7.3702
R1281 VTAIL.n28 VTAIL.n26 7.3702
R1282 VTAIL.n73 VTAIL.n6 7.3702
R1283 VTAIL.n77 VTAIL.n4 7.3702
R1284 VTAIL.n249 VTAIL.n176 7.3702
R1285 VTAIL.n245 VTAIL.n178 7.3702
R1286 VTAIL.n202 VTAIL.n200 7.3702
R1287 VTAIL.n163 VTAIL.n90 7.3702
R1288 VTAIL.n159 VTAIL.n92 7.3702
R1289 VTAIL.n116 VTAIL.n114 7.3702
R1290 VTAIL.n332 VTAIL.n331 6.59444
R1291 VTAIL.n332 VTAIL.n262 6.59444
R1292 VTAIL.n74 VTAIL.n73 6.59444
R1293 VTAIL.n74 VTAIL.n4 6.59444
R1294 VTAIL.n246 VTAIL.n176 6.59444
R1295 VTAIL.n246 VTAIL.n245 6.59444
R1296 VTAIL.n160 VTAIL.n90 6.59444
R1297 VTAIL.n160 VTAIL.n159 6.59444
R1298 VTAIL.n289 VTAIL.n284 5.81868
R1299 VTAIL.n328 VTAIL.n264 5.81868
R1300 VTAIL.n336 VTAIL.n335 5.81868
R1301 VTAIL.n31 VTAIL.n26 5.81868
R1302 VTAIL.n70 VTAIL.n6 5.81868
R1303 VTAIL.n78 VTAIL.n77 5.81868
R1304 VTAIL.n250 VTAIL.n249 5.81868
R1305 VTAIL.n242 VTAIL.n178 5.81868
R1306 VTAIL.n205 VTAIL.n200 5.81868
R1307 VTAIL.n164 VTAIL.n163 5.81868
R1308 VTAIL.n156 VTAIL.n92 5.81868
R1309 VTAIL.n119 VTAIL.n114 5.81868
R1310 VTAIL.n290 VTAIL.n282 5.04292
R1311 VTAIL.n327 VTAIL.n266 5.04292
R1312 VTAIL.n339 VTAIL.n260 5.04292
R1313 VTAIL.n32 VTAIL.n24 5.04292
R1314 VTAIL.n69 VTAIL.n8 5.04292
R1315 VTAIL.n81 VTAIL.n2 5.04292
R1316 VTAIL.n253 VTAIL.n174 5.04292
R1317 VTAIL.n241 VTAIL.n180 5.04292
R1318 VTAIL.n206 VTAIL.n198 5.04292
R1319 VTAIL.n167 VTAIL.n88 5.04292
R1320 VTAIL.n155 VTAIL.n94 5.04292
R1321 VTAIL.n120 VTAIL.n112 5.04292
R1322 VTAIL.n294 VTAIL.n293 4.26717
R1323 VTAIL.n324 VTAIL.n323 4.26717
R1324 VTAIL.n340 VTAIL.n258 4.26717
R1325 VTAIL.n36 VTAIL.n35 4.26717
R1326 VTAIL.n66 VTAIL.n65 4.26717
R1327 VTAIL.n82 VTAIL.n0 4.26717
R1328 VTAIL.n254 VTAIL.n172 4.26717
R1329 VTAIL.n238 VTAIL.n237 4.26717
R1330 VTAIL.n210 VTAIL.n209 4.26717
R1331 VTAIL.n168 VTAIL.n86 4.26717
R1332 VTAIL.n152 VTAIL.n151 4.26717
R1333 VTAIL.n124 VTAIL.n123 4.26717
R1334 VTAIL.n297 VTAIL.n280 3.49141
R1335 VTAIL.n320 VTAIL.n268 3.49141
R1336 VTAIL.n39 VTAIL.n22 3.49141
R1337 VTAIL.n62 VTAIL.n10 3.49141
R1338 VTAIL.n234 VTAIL.n182 3.49141
R1339 VTAIL.n213 VTAIL.n196 3.49141
R1340 VTAIL.n148 VTAIL.n96 3.49141
R1341 VTAIL.n127 VTAIL.n110 3.49141
R1342 VTAIL.n298 VTAIL.n278 2.71565
R1343 VTAIL.n319 VTAIL.n270 2.71565
R1344 VTAIL.n40 VTAIL.n20 2.71565
R1345 VTAIL.n61 VTAIL.n12 2.71565
R1346 VTAIL.n233 VTAIL.n184 2.71565
R1347 VTAIL.n214 VTAIL.n194 2.71565
R1348 VTAIL.n147 VTAIL.n98 2.71565
R1349 VTAIL.n128 VTAIL.n108 2.71565
R1350 VTAIL.n285 VTAIL.n283 2.41282
R1351 VTAIL.n27 VTAIL.n25 2.41282
R1352 VTAIL.n201 VTAIL.n199 2.41282
R1353 VTAIL.n115 VTAIL.n113 2.41282
R1354 VTAIL.n303 VTAIL.n301 1.93989
R1355 VTAIL.n316 VTAIL.n315 1.93989
R1356 VTAIL.n45 VTAIL.n43 1.93989
R1357 VTAIL.n58 VTAIL.n57 1.93989
R1358 VTAIL.n230 VTAIL.n229 1.93989
R1359 VTAIL.n218 VTAIL.n217 1.93989
R1360 VTAIL.n144 VTAIL.n143 1.93989
R1361 VTAIL.n132 VTAIL.n131 1.93989
R1362 VTAIL.n257 VTAIL.n171 1.24188
R1363 VTAIL.n302 VTAIL.n276 1.16414
R1364 VTAIL.n312 VTAIL.n272 1.16414
R1365 VTAIL.n44 VTAIL.n18 1.16414
R1366 VTAIL.n54 VTAIL.n14 1.16414
R1367 VTAIL.n226 VTAIL.n186 1.16414
R1368 VTAIL.n221 VTAIL.n191 1.16414
R1369 VTAIL.n140 VTAIL.n100 1.16414
R1370 VTAIL.n135 VTAIL.n105 1.16414
R1371 VTAIL VTAIL.n85 0.914293
R1372 VTAIL.n308 VTAIL.n307 0.388379
R1373 VTAIL.n311 VTAIL.n274 0.388379
R1374 VTAIL.n50 VTAIL.n49 0.388379
R1375 VTAIL.n53 VTAIL.n16 0.388379
R1376 VTAIL.n225 VTAIL.n188 0.388379
R1377 VTAIL.n222 VTAIL.n190 0.388379
R1378 VTAIL.n139 VTAIL.n102 0.388379
R1379 VTAIL.n136 VTAIL.n104 0.388379
R1380 VTAIL VTAIL.n343 0.328086
R1381 VTAIL.n291 VTAIL.n283 0.155672
R1382 VTAIL.n292 VTAIL.n291 0.155672
R1383 VTAIL.n292 VTAIL.n279 0.155672
R1384 VTAIL.n299 VTAIL.n279 0.155672
R1385 VTAIL.n300 VTAIL.n299 0.155672
R1386 VTAIL.n300 VTAIL.n275 0.155672
R1387 VTAIL.n309 VTAIL.n275 0.155672
R1388 VTAIL.n310 VTAIL.n309 0.155672
R1389 VTAIL.n310 VTAIL.n271 0.155672
R1390 VTAIL.n317 VTAIL.n271 0.155672
R1391 VTAIL.n318 VTAIL.n317 0.155672
R1392 VTAIL.n318 VTAIL.n267 0.155672
R1393 VTAIL.n325 VTAIL.n267 0.155672
R1394 VTAIL.n326 VTAIL.n325 0.155672
R1395 VTAIL.n326 VTAIL.n263 0.155672
R1396 VTAIL.n333 VTAIL.n263 0.155672
R1397 VTAIL.n334 VTAIL.n333 0.155672
R1398 VTAIL.n334 VTAIL.n259 0.155672
R1399 VTAIL.n341 VTAIL.n259 0.155672
R1400 VTAIL.n33 VTAIL.n25 0.155672
R1401 VTAIL.n34 VTAIL.n33 0.155672
R1402 VTAIL.n34 VTAIL.n21 0.155672
R1403 VTAIL.n41 VTAIL.n21 0.155672
R1404 VTAIL.n42 VTAIL.n41 0.155672
R1405 VTAIL.n42 VTAIL.n17 0.155672
R1406 VTAIL.n51 VTAIL.n17 0.155672
R1407 VTAIL.n52 VTAIL.n51 0.155672
R1408 VTAIL.n52 VTAIL.n13 0.155672
R1409 VTAIL.n59 VTAIL.n13 0.155672
R1410 VTAIL.n60 VTAIL.n59 0.155672
R1411 VTAIL.n60 VTAIL.n9 0.155672
R1412 VTAIL.n67 VTAIL.n9 0.155672
R1413 VTAIL.n68 VTAIL.n67 0.155672
R1414 VTAIL.n68 VTAIL.n5 0.155672
R1415 VTAIL.n75 VTAIL.n5 0.155672
R1416 VTAIL.n76 VTAIL.n75 0.155672
R1417 VTAIL.n76 VTAIL.n1 0.155672
R1418 VTAIL.n83 VTAIL.n1 0.155672
R1419 VTAIL.n255 VTAIL.n173 0.155672
R1420 VTAIL.n248 VTAIL.n173 0.155672
R1421 VTAIL.n248 VTAIL.n247 0.155672
R1422 VTAIL.n247 VTAIL.n177 0.155672
R1423 VTAIL.n240 VTAIL.n177 0.155672
R1424 VTAIL.n240 VTAIL.n239 0.155672
R1425 VTAIL.n239 VTAIL.n181 0.155672
R1426 VTAIL.n232 VTAIL.n181 0.155672
R1427 VTAIL.n232 VTAIL.n231 0.155672
R1428 VTAIL.n231 VTAIL.n185 0.155672
R1429 VTAIL.n224 VTAIL.n185 0.155672
R1430 VTAIL.n224 VTAIL.n223 0.155672
R1431 VTAIL.n223 VTAIL.n189 0.155672
R1432 VTAIL.n216 VTAIL.n189 0.155672
R1433 VTAIL.n216 VTAIL.n215 0.155672
R1434 VTAIL.n215 VTAIL.n195 0.155672
R1435 VTAIL.n208 VTAIL.n195 0.155672
R1436 VTAIL.n208 VTAIL.n207 0.155672
R1437 VTAIL.n207 VTAIL.n199 0.155672
R1438 VTAIL.n169 VTAIL.n87 0.155672
R1439 VTAIL.n162 VTAIL.n87 0.155672
R1440 VTAIL.n162 VTAIL.n161 0.155672
R1441 VTAIL.n161 VTAIL.n91 0.155672
R1442 VTAIL.n154 VTAIL.n91 0.155672
R1443 VTAIL.n154 VTAIL.n153 0.155672
R1444 VTAIL.n153 VTAIL.n95 0.155672
R1445 VTAIL.n146 VTAIL.n95 0.155672
R1446 VTAIL.n146 VTAIL.n145 0.155672
R1447 VTAIL.n145 VTAIL.n99 0.155672
R1448 VTAIL.n138 VTAIL.n99 0.155672
R1449 VTAIL.n138 VTAIL.n137 0.155672
R1450 VTAIL.n137 VTAIL.n103 0.155672
R1451 VTAIL.n130 VTAIL.n103 0.155672
R1452 VTAIL.n130 VTAIL.n129 0.155672
R1453 VTAIL.n129 VTAIL.n109 0.155672
R1454 VTAIL.n122 VTAIL.n109 0.155672
R1455 VTAIL.n122 VTAIL.n121 0.155672
R1456 VTAIL.n121 VTAIL.n113 0.155672
R1457 VDD2.n165 VDD2.n85 756.745
R1458 VDD2.n80 VDD2.n0 756.745
R1459 VDD2.n166 VDD2.n165 585
R1460 VDD2.n164 VDD2.n163 585
R1461 VDD2.n89 VDD2.n88 585
R1462 VDD2.n158 VDD2.n157 585
R1463 VDD2.n156 VDD2.n155 585
R1464 VDD2.n93 VDD2.n92 585
R1465 VDD2.n150 VDD2.n149 585
R1466 VDD2.n148 VDD2.n147 585
R1467 VDD2.n97 VDD2.n96 585
R1468 VDD2.n142 VDD2.n141 585
R1469 VDD2.n140 VDD2.n139 585
R1470 VDD2.n101 VDD2.n100 585
R1471 VDD2.n105 VDD2.n103 585
R1472 VDD2.n134 VDD2.n133 585
R1473 VDD2.n132 VDD2.n131 585
R1474 VDD2.n107 VDD2.n106 585
R1475 VDD2.n126 VDD2.n125 585
R1476 VDD2.n124 VDD2.n123 585
R1477 VDD2.n111 VDD2.n110 585
R1478 VDD2.n118 VDD2.n117 585
R1479 VDD2.n116 VDD2.n115 585
R1480 VDD2.n29 VDD2.n28 585
R1481 VDD2.n31 VDD2.n30 585
R1482 VDD2.n24 VDD2.n23 585
R1483 VDD2.n37 VDD2.n36 585
R1484 VDD2.n39 VDD2.n38 585
R1485 VDD2.n20 VDD2.n19 585
R1486 VDD2.n46 VDD2.n45 585
R1487 VDD2.n47 VDD2.n18 585
R1488 VDD2.n49 VDD2.n48 585
R1489 VDD2.n16 VDD2.n15 585
R1490 VDD2.n55 VDD2.n54 585
R1491 VDD2.n57 VDD2.n56 585
R1492 VDD2.n12 VDD2.n11 585
R1493 VDD2.n63 VDD2.n62 585
R1494 VDD2.n65 VDD2.n64 585
R1495 VDD2.n8 VDD2.n7 585
R1496 VDD2.n71 VDD2.n70 585
R1497 VDD2.n73 VDD2.n72 585
R1498 VDD2.n4 VDD2.n3 585
R1499 VDD2.n79 VDD2.n78 585
R1500 VDD2.n81 VDD2.n80 585
R1501 VDD2.n114 VDD2.t0 329.036
R1502 VDD2.n27 VDD2.t1 329.036
R1503 VDD2.n165 VDD2.n164 171.744
R1504 VDD2.n164 VDD2.n88 171.744
R1505 VDD2.n157 VDD2.n88 171.744
R1506 VDD2.n157 VDD2.n156 171.744
R1507 VDD2.n156 VDD2.n92 171.744
R1508 VDD2.n149 VDD2.n92 171.744
R1509 VDD2.n149 VDD2.n148 171.744
R1510 VDD2.n148 VDD2.n96 171.744
R1511 VDD2.n141 VDD2.n96 171.744
R1512 VDD2.n141 VDD2.n140 171.744
R1513 VDD2.n140 VDD2.n100 171.744
R1514 VDD2.n105 VDD2.n100 171.744
R1515 VDD2.n133 VDD2.n105 171.744
R1516 VDD2.n133 VDD2.n132 171.744
R1517 VDD2.n132 VDD2.n106 171.744
R1518 VDD2.n125 VDD2.n106 171.744
R1519 VDD2.n125 VDD2.n124 171.744
R1520 VDD2.n124 VDD2.n110 171.744
R1521 VDD2.n117 VDD2.n110 171.744
R1522 VDD2.n117 VDD2.n116 171.744
R1523 VDD2.n30 VDD2.n29 171.744
R1524 VDD2.n30 VDD2.n23 171.744
R1525 VDD2.n37 VDD2.n23 171.744
R1526 VDD2.n38 VDD2.n37 171.744
R1527 VDD2.n38 VDD2.n19 171.744
R1528 VDD2.n46 VDD2.n19 171.744
R1529 VDD2.n47 VDD2.n46 171.744
R1530 VDD2.n48 VDD2.n47 171.744
R1531 VDD2.n48 VDD2.n15 171.744
R1532 VDD2.n55 VDD2.n15 171.744
R1533 VDD2.n56 VDD2.n55 171.744
R1534 VDD2.n56 VDD2.n11 171.744
R1535 VDD2.n63 VDD2.n11 171.744
R1536 VDD2.n64 VDD2.n63 171.744
R1537 VDD2.n64 VDD2.n7 171.744
R1538 VDD2.n71 VDD2.n7 171.744
R1539 VDD2.n72 VDD2.n71 171.744
R1540 VDD2.n72 VDD2.n3 171.744
R1541 VDD2.n79 VDD2.n3 171.744
R1542 VDD2.n80 VDD2.n79 171.744
R1543 VDD2.n170 VDD2.n84 87.1359
R1544 VDD2.n116 VDD2.t0 85.8723
R1545 VDD2.n29 VDD2.t1 85.8723
R1546 VDD2.n170 VDD2.n169 46.9247
R1547 VDD2.n103 VDD2.n101 13.1884
R1548 VDD2.n49 VDD2.n16 13.1884
R1549 VDD2.n139 VDD2.n138 12.8005
R1550 VDD2.n135 VDD2.n134 12.8005
R1551 VDD2.n50 VDD2.n18 12.8005
R1552 VDD2.n54 VDD2.n53 12.8005
R1553 VDD2.n142 VDD2.n99 12.0247
R1554 VDD2.n131 VDD2.n104 12.0247
R1555 VDD2.n45 VDD2.n44 12.0247
R1556 VDD2.n57 VDD2.n14 12.0247
R1557 VDD2.n143 VDD2.n97 11.249
R1558 VDD2.n130 VDD2.n107 11.249
R1559 VDD2.n43 VDD2.n20 11.249
R1560 VDD2.n58 VDD2.n12 11.249
R1561 VDD2.n115 VDD2.n114 10.7239
R1562 VDD2.n28 VDD2.n27 10.7239
R1563 VDD2.n147 VDD2.n146 10.4732
R1564 VDD2.n127 VDD2.n126 10.4732
R1565 VDD2.n40 VDD2.n39 10.4732
R1566 VDD2.n62 VDD2.n61 10.4732
R1567 VDD2.n169 VDD2.n85 9.69747
R1568 VDD2.n150 VDD2.n95 9.69747
R1569 VDD2.n123 VDD2.n109 9.69747
R1570 VDD2.n36 VDD2.n22 9.69747
R1571 VDD2.n65 VDD2.n10 9.69747
R1572 VDD2.n84 VDD2.n0 9.69747
R1573 VDD2.n169 VDD2.n168 9.45567
R1574 VDD2.n84 VDD2.n83 9.45567
R1575 VDD2.n87 VDD2.n86 9.3005
R1576 VDD2.n162 VDD2.n161 9.3005
R1577 VDD2.n160 VDD2.n159 9.3005
R1578 VDD2.n91 VDD2.n90 9.3005
R1579 VDD2.n154 VDD2.n153 9.3005
R1580 VDD2.n152 VDD2.n151 9.3005
R1581 VDD2.n95 VDD2.n94 9.3005
R1582 VDD2.n146 VDD2.n145 9.3005
R1583 VDD2.n144 VDD2.n143 9.3005
R1584 VDD2.n99 VDD2.n98 9.3005
R1585 VDD2.n138 VDD2.n137 9.3005
R1586 VDD2.n136 VDD2.n135 9.3005
R1587 VDD2.n104 VDD2.n102 9.3005
R1588 VDD2.n130 VDD2.n129 9.3005
R1589 VDD2.n128 VDD2.n127 9.3005
R1590 VDD2.n109 VDD2.n108 9.3005
R1591 VDD2.n122 VDD2.n121 9.3005
R1592 VDD2.n120 VDD2.n119 9.3005
R1593 VDD2.n113 VDD2.n112 9.3005
R1594 VDD2.n168 VDD2.n167 9.3005
R1595 VDD2.n75 VDD2.n74 9.3005
R1596 VDD2.n77 VDD2.n76 9.3005
R1597 VDD2.n2 VDD2.n1 9.3005
R1598 VDD2.n83 VDD2.n82 9.3005
R1599 VDD2.n69 VDD2.n68 9.3005
R1600 VDD2.n67 VDD2.n66 9.3005
R1601 VDD2.n10 VDD2.n9 9.3005
R1602 VDD2.n61 VDD2.n60 9.3005
R1603 VDD2.n59 VDD2.n58 9.3005
R1604 VDD2.n14 VDD2.n13 9.3005
R1605 VDD2.n53 VDD2.n52 9.3005
R1606 VDD2.n26 VDD2.n25 9.3005
R1607 VDD2.n33 VDD2.n32 9.3005
R1608 VDD2.n35 VDD2.n34 9.3005
R1609 VDD2.n22 VDD2.n21 9.3005
R1610 VDD2.n41 VDD2.n40 9.3005
R1611 VDD2.n43 VDD2.n42 9.3005
R1612 VDD2.n44 VDD2.n17 9.3005
R1613 VDD2.n51 VDD2.n50 9.3005
R1614 VDD2.n6 VDD2.n5 9.3005
R1615 VDD2.n167 VDD2.n166 8.92171
R1616 VDD2.n151 VDD2.n93 8.92171
R1617 VDD2.n122 VDD2.n111 8.92171
R1618 VDD2.n35 VDD2.n24 8.92171
R1619 VDD2.n66 VDD2.n8 8.92171
R1620 VDD2.n82 VDD2.n81 8.92171
R1621 VDD2.n163 VDD2.n87 8.14595
R1622 VDD2.n155 VDD2.n154 8.14595
R1623 VDD2.n119 VDD2.n118 8.14595
R1624 VDD2.n32 VDD2.n31 8.14595
R1625 VDD2.n70 VDD2.n69 8.14595
R1626 VDD2.n78 VDD2.n2 8.14595
R1627 VDD2.n162 VDD2.n89 7.3702
R1628 VDD2.n158 VDD2.n91 7.3702
R1629 VDD2.n115 VDD2.n113 7.3702
R1630 VDD2.n28 VDD2.n26 7.3702
R1631 VDD2.n73 VDD2.n6 7.3702
R1632 VDD2.n77 VDD2.n4 7.3702
R1633 VDD2.n159 VDD2.n89 6.59444
R1634 VDD2.n159 VDD2.n158 6.59444
R1635 VDD2.n74 VDD2.n73 6.59444
R1636 VDD2.n74 VDD2.n4 6.59444
R1637 VDD2.n163 VDD2.n162 5.81868
R1638 VDD2.n155 VDD2.n91 5.81868
R1639 VDD2.n118 VDD2.n113 5.81868
R1640 VDD2.n31 VDD2.n26 5.81868
R1641 VDD2.n70 VDD2.n6 5.81868
R1642 VDD2.n78 VDD2.n77 5.81868
R1643 VDD2.n166 VDD2.n87 5.04292
R1644 VDD2.n154 VDD2.n93 5.04292
R1645 VDD2.n119 VDD2.n111 5.04292
R1646 VDD2.n32 VDD2.n24 5.04292
R1647 VDD2.n69 VDD2.n8 5.04292
R1648 VDD2.n81 VDD2.n2 5.04292
R1649 VDD2.n167 VDD2.n85 4.26717
R1650 VDD2.n151 VDD2.n150 4.26717
R1651 VDD2.n123 VDD2.n122 4.26717
R1652 VDD2.n36 VDD2.n35 4.26717
R1653 VDD2.n66 VDD2.n65 4.26717
R1654 VDD2.n82 VDD2.n0 4.26717
R1655 VDD2.n147 VDD2.n95 3.49141
R1656 VDD2.n126 VDD2.n109 3.49141
R1657 VDD2.n39 VDD2.n22 3.49141
R1658 VDD2.n62 VDD2.n10 3.49141
R1659 VDD2.n146 VDD2.n97 2.71565
R1660 VDD2.n127 VDD2.n107 2.71565
R1661 VDD2.n40 VDD2.n20 2.71565
R1662 VDD2.n61 VDD2.n12 2.71565
R1663 VDD2.n114 VDD2.n112 2.41282
R1664 VDD2.n27 VDD2.n25 2.41282
R1665 VDD2.n143 VDD2.n142 1.93989
R1666 VDD2.n131 VDD2.n130 1.93989
R1667 VDD2.n45 VDD2.n43 1.93989
R1668 VDD2.n58 VDD2.n57 1.93989
R1669 VDD2.n139 VDD2.n99 1.16414
R1670 VDD2.n134 VDD2.n104 1.16414
R1671 VDD2.n44 VDD2.n18 1.16414
R1672 VDD2.n54 VDD2.n14 1.16414
R1673 VDD2 VDD2.n170 0.444466
R1674 VDD2.n138 VDD2.n101 0.388379
R1675 VDD2.n135 VDD2.n103 0.388379
R1676 VDD2.n50 VDD2.n49 0.388379
R1677 VDD2.n53 VDD2.n16 0.388379
R1678 VDD2.n168 VDD2.n86 0.155672
R1679 VDD2.n161 VDD2.n86 0.155672
R1680 VDD2.n161 VDD2.n160 0.155672
R1681 VDD2.n160 VDD2.n90 0.155672
R1682 VDD2.n153 VDD2.n90 0.155672
R1683 VDD2.n153 VDD2.n152 0.155672
R1684 VDD2.n152 VDD2.n94 0.155672
R1685 VDD2.n145 VDD2.n94 0.155672
R1686 VDD2.n145 VDD2.n144 0.155672
R1687 VDD2.n144 VDD2.n98 0.155672
R1688 VDD2.n137 VDD2.n98 0.155672
R1689 VDD2.n137 VDD2.n136 0.155672
R1690 VDD2.n136 VDD2.n102 0.155672
R1691 VDD2.n129 VDD2.n102 0.155672
R1692 VDD2.n129 VDD2.n128 0.155672
R1693 VDD2.n128 VDD2.n108 0.155672
R1694 VDD2.n121 VDD2.n108 0.155672
R1695 VDD2.n121 VDD2.n120 0.155672
R1696 VDD2.n120 VDD2.n112 0.155672
R1697 VDD2.n33 VDD2.n25 0.155672
R1698 VDD2.n34 VDD2.n33 0.155672
R1699 VDD2.n34 VDD2.n21 0.155672
R1700 VDD2.n41 VDD2.n21 0.155672
R1701 VDD2.n42 VDD2.n41 0.155672
R1702 VDD2.n42 VDD2.n17 0.155672
R1703 VDD2.n51 VDD2.n17 0.155672
R1704 VDD2.n52 VDD2.n51 0.155672
R1705 VDD2.n52 VDD2.n13 0.155672
R1706 VDD2.n59 VDD2.n13 0.155672
R1707 VDD2.n60 VDD2.n59 0.155672
R1708 VDD2.n60 VDD2.n9 0.155672
R1709 VDD2.n67 VDD2.n9 0.155672
R1710 VDD2.n68 VDD2.n67 0.155672
R1711 VDD2.n68 VDD2.n5 0.155672
R1712 VDD2.n75 VDD2.n5 0.155672
R1713 VDD2.n76 VDD2.n75 0.155672
R1714 VDD2.n76 VDD2.n1 0.155672
R1715 VDD2.n83 VDD2.n1 0.155672
R1716 VP.n0 VP.t0 409.723
R1717 VP.n0 VP.t1 365.346
R1718 VP VP.n0 0.146778
R1719 VDD1.n80 VDD1.n0 756.745
R1720 VDD1.n165 VDD1.n85 756.745
R1721 VDD1.n81 VDD1.n80 585
R1722 VDD1.n79 VDD1.n78 585
R1723 VDD1.n4 VDD1.n3 585
R1724 VDD1.n73 VDD1.n72 585
R1725 VDD1.n71 VDD1.n70 585
R1726 VDD1.n8 VDD1.n7 585
R1727 VDD1.n65 VDD1.n64 585
R1728 VDD1.n63 VDD1.n62 585
R1729 VDD1.n12 VDD1.n11 585
R1730 VDD1.n57 VDD1.n56 585
R1731 VDD1.n55 VDD1.n54 585
R1732 VDD1.n16 VDD1.n15 585
R1733 VDD1.n20 VDD1.n18 585
R1734 VDD1.n49 VDD1.n48 585
R1735 VDD1.n47 VDD1.n46 585
R1736 VDD1.n22 VDD1.n21 585
R1737 VDD1.n41 VDD1.n40 585
R1738 VDD1.n39 VDD1.n38 585
R1739 VDD1.n26 VDD1.n25 585
R1740 VDD1.n33 VDD1.n32 585
R1741 VDD1.n31 VDD1.n30 585
R1742 VDD1.n114 VDD1.n113 585
R1743 VDD1.n116 VDD1.n115 585
R1744 VDD1.n109 VDD1.n108 585
R1745 VDD1.n122 VDD1.n121 585
R1746 VDD1.n124 VDD1.n123 585
R1747 VDD1.n105 VDD1.n104 585
R1748 VDD1.n131 VDD1.n130 585
R1749 VDD1.n132 VDD1.n103 585
R1750 VDD1.n134 VDD1.n133 585
R1751 VDD1.n101 VDD1.n100 585
R1752 VDD1.n140 VDD1.n139 585
R1753 VDD1.n142 VDD1.n141 585
R1754 VDD1.n97 VDD1.n96 585
R1755 VDD1.n148 VDD1.n147 585
R1756 VDD1.n150 VDD1.n149 585
R1757 VDD1.n93 VDD1.n92 585
R1758 VDD1.n156 VDD1.n155 585
R1759 VDD1.n158 VDD1.n157 585
R1760 VDD1.n89 VDD1.n88 585
R1761 VDD1.n164 VDD1.n163 585
R1762 VDD1.n166 VDD1.n165 585
R1763 VDD1.n29 VDD1.t1 329.036
R1764 VDD1.n112 VDD1.t0 329.036
R1765 VDD1.n80 VDD1.n79 171.744
R1766 VDD1.n79 VDD1.n3 171.744
R1767 VDD1.n72 VDD1.n3 171.744
R1768 VDD1.n72 VDD1.n71 171.744
R1769 VDD1.n71 VDD1.n7 171.744
R1770 VDD1.n64 VDD1.n7 171.744
R1771 VDD1.n64 VDD1.n63 171.744
R1772 VDD1.n63 VDD1.n11 171.744
R1773 VDD1.n56 VDD1.n11 171.744
R1774 VDD1.n56 VDD1.n55 171.744
R1775 VDD1.n55 VDD1.n15 171.744
R1776 VDD1.n20 VDD1.n15 171.744
R1777 VDD1.n48 VDD1.n20 171.744
R1778 VDD1.n48 VDD1.n47 171.744
R1779 VDD1.n47 VDD1.n21 171.744
R1780 VDD1.n40 VDD1.n21 171.744
R1781 VDD1.n40 VDD1.n39 171.744
R1782 VDD1.n39 VDD1.n25 171.744
R1783 VDD1.n32 VDD1.n25 171.744
R1784 VDD1.n32 VDD1.n31 171.744
R1785 VDD1.n115 VDD1.n114 171.744
R1786 VDD1.n115 VDD1.n108 171.744
R1787 VDD1.n122 VDD1.n108 171.744
R1788 VDD1.n123 VDD1.n122 171.744
R1789 VDD1.n123 VDD1.n104 171.744
R1790 VDD1.n131 VDD1.n104 171.744
R1791 VDD1.n132 VDD1.n131 171.744
R1792 VDD1.n133 VDD1.n132 171.744
R1793 VDD1.n133 VDD1.n100 171.744
R1794 VDD1.n140 VDD1.n100 171.744
R1795 VDD1.n141 VDD1.n140 171.744
R1796 VDD1.n141 VDD1.n96 171.744
R1797 VDD1.n148 VDD1.n96 171.744
R1798 VDD1.n149 VDD1.n148 171.744
R1799 VDD1.n149 VDD1.n92 171.744
R1800 VDD1.n156 VDD1.n92 171.744
R1801 VDD1.n157 VDD1.n156 171.744
R1802 VDD1.n157 VDD1.n88 171.744
R1803 VDD1.n164 VDD1.n88 171.744
R1804 VDD1.n165 VDD1.n164 171.744
R1805 VDD1 VDD1.n169 88.0465
R1806 VDD1.n31 VDD1.t1 85.8723
R1807 VDD1.n114 VDD1.t0 85.8723
R1808 VDD1 VDD1.n84 47.3687
R1809 VDD1.n18 VDD1.n16 13.1884
R1810 VDD1.n134 VDD1.n101 13.1884
R1811 VDD1.n54 VDD1.n53 12.8005
R1812 VDD1.n50 VDD1.n49 12.8005
R1813 VDD1.n135 VDD1.n103 12.8005
R1814 VDD1.n139 VDD1.n138 12.8005
R1815 VDD1.n57 VDD1.n14 12.0247
R1816 VDD1.n46 VDD1.n19 12.0247
R1817 VDD1.n130 VDD1.n129 12.0247
R1818 VDD1.n142 VDD1.n99 12.0247
R1819 VDD1.n58 VDD1.n12 11.249
R1820 VDD1.n45 VDD1.n22 11.249
R1821 VDD1.n128 VDD1.n105 11.249
R1822 VDD1.n143 VDD1.n97 11.249
R1823 VDD1.n30 VDD1.n29 10.7239
R1824 VDD1.n113 VDD1.n112 10.7239
R1825 VDD1.n62 VDD1.n61 10.4732
R1826 VDD1.n42 VDD1.n41 10.4732
R1827 VDD1.n125 VDD1.n124 10.4732
R1828 VDD1.n147 VDD1.n146 10.4732
R1829 VDD1.n84 VDD1.n0 9.69747
R1830 VDD1.n65 VDD1.n10 9.69747
R1831 VDD1.n38 VDD1.n24 9.69747
R1832 VDD1.n121 VDD1.n107 9.69747
R1833 VDD1.n150 VDD1.n95 9.69747
R1834 VDD1.n169 VDD1.n85 9.69747
R1835 VDD1.n84 VDD1.n83 9.45567
R1836 VDD1.n169 VDD1.n168 9.45567
R1837 VDD1.n2 VDD1.n1 9.3005
R1838 VDD1.n77 VDD1.n76 9.3005
R1839 VDD1.n75 VDD1.n74 9.3005
R1840 VDD1.n6 VDD1.n5 9.3005
R1841 VDD1.n69 VDD1.n68 9.3005
R1842 VDD1.n67 VDD1.n66 9.3005
R1843 VDD1.n10 VDD1.n9 9.3005
R1844 VDD1.n61 VDD1.n60 9.3005
R1845 VDD1.n59 VDD1.n58 9.3005
R1846 VDD1.n14 VDD1.n13 9.3005
R1847 VDD1.n53 VDD1.n52 9.3005
R1848 VDD1.n51 VDD1.n50 9.3005
R1849 VDD1.n19 VDD1.n17 9.3005
R1850 VDD1.n45 VDD1.n44 9.3005
R1851 VDD1.n43 VDD1.n42 9.3005
R1852 VDD1.n24 VDD1.n23 9.3005
R1853 VDD1.n37 VDD1.n36 9.3005
R1854 VDD1.n35 VDD1.n34 9.3005
R1855 VDD1.n28 VDD1.n27 9.3005
R1856 VDD1.n83 VDD1.n82 9.3005
R1857 VDD1.n160 VDD1.n159 9.3005
R1858 VDD1.n162 VDD1.n161 9.3005
R1859 VDD1.n87 VDD1.n86 9.3005
R1860 VDD1.n168 VDD1.n167 9.3005
R1861 VDD1.n154 VDD1.n153 9.3005
R1862 VDD1.n152 VDD1.n151 9.3005
R1863 VDD1.n95 VDD1.n94 9.3005
R1864 VDD1.n146 VDD1.n145 9.3005
R1865 VDD1.n144 VDD1.n143 9.3005
R1866 VDD1.n99 VDD1.n98 9.3005
R1867 VDD1.n138 VDD1.n137 9.3005
R1868 VDD1.n111 VDD1.n110 9.3005
R1869 VDD1.n118 VDD1.n117 9.3005
R1870 VDD1.n120 VDD1.n119 9.3005
R1871 VDD1.n107 VDD1.n106 9.3005
R1872 VDD1.n126 VDD1.n125 9.3005
R1873 VDD1.n128 VDD1.n127 9.3005
R1874 VDD1.n129 VDD1.n102 9.3005
R1875 VDD1.n136 VDD1.n135 9.3005
R1876 VDD1.n91 VDD1.n90 9.3005
R1877 VDD1.n82 VDD1.n81 8.92171
R1878 VDD1.n66 VDD1.n8 8.92171
R1879 VDD1.n37 VDD1.n26 8.92171
R1880 VDD1.n120 VDD1.n109 8.92171
R1881 VDD1.n151 VDD1.n93 8.92171
R1882 VDD1.n167 VDD1.n166 8.92171
R1883 VDD1.n78 VDD1.n2 8.14595
R1884 VDD1.n70 VDD1.n69 8.14595
R1885 VDD1.n34 VDD1.n33 8.14595
R1886 VDD1.n117 VDD1.n116 8.14595
R1887 VDD1.n155 VDD1.n154 8.14595
R1888 VDD1.n163 VDD1.n87 8.14595
R1889 VDD1.n77 VDD1.n4 7.3702
R1890 VDD1.n73 VDD1.n6 7.3702
R1891 VDD1.n30 VDD1.n28 7.3702
R1892 VDD1.n113 VDD1.n111 7.3702
R1893 VDD1.n158 VDD1.n91 7.3702
R1894 VDD1.n162 VDD1.n89 7.3702
R1895 VDD1.n74 VDD1.n4 6.59444
R1896 VDD1.n74 VDD1.n73 6.59444
R1897 VDD1.n159 VDD1.n158 6.59444
R1898 VDD1.n159 VDD1.n89 6.59444
R1899 VDD1.n78 VDD1.n77 5.81868
R1900 VDD1.n70 VDD1.n6 5.81868
R1901 VDD1.n33 VDD1.n28 5.81868
R1902 VDD1.n116 VDD1.n111 5.81868
R1903 VDD1.n155 VDD1.n91 5.81868
R1904 VDD1.n163 VDD1.n162 5.81868
R1905 VDD1.n81 VDD1.n2 5.04292
R1906 VDD1.n69 VDD1.n8 5.04292
R1907 VDD1.n34 VDD1.n26 5.04292
R1908 VDD1.n117 VDD1.n109 5.04292
R1909 VDD1.n154 VDD1.n93 5.04292
R1910 VDD1.n166 VDD1.n87 5.04292
R1911 VDD1.n82 VDD1.n0 4.26717
R1912 VDD1.n66 VDD1.n65 4.26717
R1913 VDD1.n38 VDD1.n37 4.26717
R1914 VDD1.n121 VDD1.n120 4.26717
R1915 VDD1.n151 VDD1.n150 4.26717
R1916 VDD1.n167 VDD1.n85 4.26717
R1917 VDD1.n62 VDD1.n10 3.49141
R1918 VDD1.n41 VDD1.n24 3.49141
R1919 VDD1.n124 VDD1.n107 3.49141
R1920 VDD1.n147 VDD1.n95 3.49141
R1921 VDD1.n61 VDD1.n12 2.71565
R1922 VDD1.n42 VDD1.n22 2.71565
R1923 VDD1.n125 VDD1.n105 2.71565
R1924 VDD1.n146 VDD1.n97 2.71565
R1925 VDD1.n29 VDD1.n27 2.41282
R1926 VDD1.n112 VDD1.n110 2.41282
R1927 VDD1.n58 VDD1.n57 1.93989
R1928 VDD1.n46 VDD1.n45 1.93989
R1929 VDD1.n130 VDD1.n128 1.93989
R1930 VDD1.n143 VDD1.n142 1.93989
R1931 VDD1.n54 VDD1.n14 1.16414
R1932 VDD1.n49 VDD1.n19 1.16414
R1933 VDD1.n129 VDD1.n103 1.16414
R1934 VDD1.n139 VDD1.n99 1.16414
R1935 VDD1.n53 VDD1.n16 0.388379
R1936 VDD1.n50 VDD1.n18 0.388379
R1937 VDD1.n135 VDD1.n134 0.388379
R1938 VDD1.n138 VDD1.n101 0.388379
R1939 VDD1.n83 VDD1.n1 0.155672
R1940 VDD1.n76 VDD1.n1 0.155672
R1941 VDD1.n76 VDD1.n75 0.155672
R1942 VDD1.n75 VDD1.n5 0.155672
R1943 VDD1.n68 VDD1.n5 0.155672
R1944 VDD1.n68 VDD1.n67 0.155672
R1945 VDD1.n67 VDD1.n9 0.155672
R1946 VDD1.n60 VDD1.n9 0.155672
R1947 VDD1.n60 VDD1.n59 0.155672
R1948 VDD1.n59 VDD1.n13 0.155672
R1949 VDD1.n52 VDD1.n13 0.155672
R1950 VDD1.n52 VDD1.n51 0.155672
R1951 VDD1.n51 VDD1.n17 0.155672
R1952 VDD1.n44 VDD1.n17 0.155672
R1953 VDD1.n44 VDD1.n43 0.155672
R1954 VDD1.n43 VDD1.n23 0.155672
R1955 VDD1.n36 VDD1.n23 0.155672
R1956 VDD1.n36 VDD1.n35 0.155672
R1957 VDD1.n35 VDD1.n27 0.155672
R1958 VDD1.n118 VDD1.n110 0.155672
R1959 VDD1.n119 VDD1.n118 0.155672
R1960 VDD1.n119 VDD1.n106 0.155672
R1961 VDD1.n126 VDD1.n106 0.155672
R1962 VDD1.n127 VDD1.n126 0.155672
R1963 VDD1.n127 VDD1.n102 0.155672
R1964 VDD1.n136 VDD1.n102 0.155672
R1965 VDD1.n137 VDD1.n136 0.155672
R1966 VDD1.n137 VDD1.n98 0.155672
R1967 VDD1.n144 VDD1.n98 0.155672
R1968 VDD1.n145 VDD1.n144 0.155672
R1969 VDD1.n145 VDD1.n94 0.155672
R1970 VDD1.n152 VDD1.n94 0.155672
R1971 VDD1.n153 VDD1.n152 0.155672
R1972 VDD1.n153 VDD1.n90 0.155672
R1973 VDD1.n160 VDD1.n90 0.155672
R1974 VDD1.n161 VDD1.n160 0.155672
R1975 VDD1.n161 VDD1.n86 0.155672
R1976 VDD1.n168 VDD1.n86 0.155672
C0 VTAIL B 3.86338f
C1 VDD1 VDD2 0.542403f
C2 VDD1 B 1.8177f
C3 w_n1686_n4092# VN 2.2897f
C4 VDD2 B 1.8378f
C5 VP VN 5.5867f
C6 w_n1686_n4092# VP 2.50201f
C7 VTAIL VN 2.59698f
C8 w_n1686_n4092# VTAIL 3.34142f
C9 VTAIL VP 2.6115f
C10 VDD1 VN 0.147933f
C11 VDD2 VN 3.15811f
C12 w_n1686_n4092# VDD1 1.91283f
C13 w_n1686_n4092# VDD2 1.92523f
C14 VDD1 VP 3.29196f
C15 VP VDD2 0.286068f
C16 VN B 0.902473f
C17 VDD1 VTAIL 6.15606f
C18 VTAIL VDD2 6.19591f
C19 w_n1686_n4092# B 8.59134f
C20 VP B 1.24694f
C21 VDD2 VSUBS 0.917945f
C22 VDD1 VSUBS 3.72332f
C23 VTAIL VSUBS 1.014603f
C24 VN VSUBS 8.38399f
C25 VP VSUBS 1.475934f
C26 B VSUBS 3.357009f
C27 w_n1686_n4092# VSUBS 84.5495f
C28 VDD1.n0 VSUBS 0.02301f
C29 VDD1.n1 VSUBS 0.020237f
C30 VDD1.n2 VSUBS 0.010875f
C31 VDD1.n3 VSUBS 0.025704f
C32 VDD1.n4 VSUBS 0.011514f
C33 VDD1.n5 VSUBS 0.020237f
C34 VDD1.n6 VSUBS 0.010875f
C35 VDD1.n7 VSUBS 0.025704f
C36 VDD1.n8 VSUBS 0.011514f
C37 VDD1.n9 VSUBS 0.020237f
C38 VDD1.n10 VSUBS 0.010875f
C39 VDD1.n11 VSUBS 0.025704f
C40 VDD1.n12 VSUBS 0.011514f
C41 VDD1.n13 VSUBS 0.020237f
C42 VDD1.n14 VSUBS 0.010875f
C43 VDD1.n15 VSUBS 0.025704f
C44 VDD1.n16 VSUBS 0.011195f
C45 VDD1.n17 VSUBS 0.020237f
C46 VDD1.n18 VSUBS 0.011195f
C47 VDD1.n19 VSUBS 0.010875f
C48 VDD1.n20 VSUBS 0.025704f
C49 VDD1.n21 VSUBS 0.025704f
C50 VDD1.n22 VSUBS 0.011514f
C51 VDD1.n23 VSUBS 0.020237f
C52 VDD1.n24 VSUBS 0.010875f
C53 VDD1.n25 VSUBS 0.025704f
C54 VDD1.n26 VSUBS 0.011514f
C55 VDD1.n27 VSUBS 1.31532f
C56 VDD1.n28 VSUBS 0.010875f
C57 VDD1.t1 VSUBS 0.055634f
C58 VDD1.n29 VSUBS 0.192504f
C59 VDD1.n30 VSUBS 0.019336f
C60 VDD1.n31 VSUBS 0.019278f
C61 VDD1.n32 VSUBS 0.025704f
C62 VDD1.n33 VSUBS 0.011514f
C63 VDD1.n34 VSUBS 0.010875f
C64 VDD1.n35 VSUBS 0.020237f
C65 VDD1.n36 VSUBS 0.020237f
C66 VDD1.n37 VSUBS 0.010875f
C67 VDD1.n38 VSUBS 0.011514f
C68 VDD1.n39 VSUBS 0.025704f
C69 VDD1.n40 VSUBS 0.025704f
C70 VDD1.n41 VSUBS 0.011514f
C71 VDD1.n42 VSUBS 0.010875f
C72 VDD1.n43 VSUBS 0.020237f
C73 VDD1.n44 VSUBS 0.020237f
C74 VDD1.n45 VSUBS 0.010875f
C75 VDD1.n46 VSUBS 0.011514f
C76 VDD1.n47 VSUBS 0.025704f
C77 VDD1.n48 VSUBS 0.025704f
C78 VDD1.n49 VSUBS 0.011514f
C79 VDD1.n50 VSUBS 0.010875f
C80 VDD1.n51 VSUBS 0.020237f
C81 VDD1.n52 VSUBS 0.020237f
C82 VDD1.n53 VSUBS 0.010875f
C83 VDD1.n54 VSUBS 0.011514f
C84 VDD1.n55 VSUBS 0.025704f
C85 VDD1.n56 VSUBS 0.025704f
C86 VDD1.n57 VSUBS 0.011514f
C87 VDD1.n58 VSUBS 0.010875f
C88 VDD1.n59 VSUBS 0.020237f
C89 VDD1.n60 VSUBS 0.020237f
C90 VDD1.n61 VSUBS 0.010875f
C91 VDD1.n62 VSUBS 0.011514f
C92 VDD1.n63 VSUBS 0.025704f
C93 VDD1.n64 VSUBS 0.025704f
C94 VDD1.n65 VSUBS 0.011514f
C95 VDD1.n66 VSUBS 0.010875f
C96 VDD1.n67 VSUBS 0.020237f
C97 VDD1.n68 VSUBS 0.020237f
C98 VDD1.n69 VSUBS 0.010875f
C99 VDD1.n70 VSUBS 0.011514f
C100 VDD1.n71 VSUBS 0.025704f
C101 VDD1.n72 VSUBS 0.025704f
C102 VDD1.n73 VSUBS 0.011514f
C103 VDD1.n74 VSUBS 0.010875f
C104 VDD1.n75 VSUBS 0.020237f
C105 VDD1.n76 VSUBS 0.020237f
C106 VDD1.n77 VSUBS 0.010875f
C107 VDD1.n78 VSUBS 0.011514f
C108 VDD1.n79 VSUBS 0.025704f
C109 VDD1.n80 VSUBS 0.06486f
C110 VDD1.n81 VSUBS 0.011514f
C111 VDD1.n82 VSUBS 0.010875f
C112 VDD1.n83 VSUBS 0.044013f
C113 VDD1.n84 VSUBS 0.047266f
C114 VDD1.n85 VSUBS 0.02301f
C115 VDD1.n86 VSUBS 0.020237f
C116 VDD1.n87 VSUBS 0.010875f
C117 VDD1.n88 VSUBS 0.025704f
C118 VDD1.n89 VSUBS 0.011514f
C119 VDD1.n90 VSUBS 0.020237f
C120 VDD1.n91 VSUBS 0.010875f
C121 VDD1.n92 VSUBS 0.025704f
C122 VDD1.n93 VSUBS 0.011514f
C123 VDD1.n94 VSUBS 0.020237f
C124 VDD1.n95 VSUBS 0.010875f
C125 VDD1.n96 VSUBS 0.025704f
C126 VDD1.n97 VSUBS 0.011514f
C127 VDD1.n98 VSUBS 0.020237f
C128 VDD1.n99 VSUBS 0.010875f
C129 VDD1.n100 VSUBS 0.025704f
C130 VDD1.n101 VSUBS 0.011195f
C131 VDD1.n102 VSUBS 0.020237f
C132 VDD1.n103 VSUBS 0.011514f
C133 VDD1.n104 VSUBS 0.025704f
C134 VDD1.n105 VSUBS 0.011514f
C135 VDD1.n106 VSUBS 0.020237f
C136 VDD1.n107 VSUBS 0.010875f
C137 VDD1.n108 VSUBS 0.025704f
C138 VDD1.n109 VSUBS 0.011514f
C139 VDD1.n110 VSUBS 1.31532f
C140 VDD1.n111 VSUBS 0.010875f
C141 VDD1.t0 VSUBS 0.055634f
C142 VDD1.n112 VSUBS 0.192504f
C143 VDD1.n113 VSUBS 0.019336f
C144 VDD1.n114 VSUBS 0.019278f
C145 VDD1.n115 VSUBS 0.025704f
C146 VDD1.n116 VSUBS 0.011514f
C147 VDD1.n117 VSUBS 0.010875f
C148 VDD1.n118 VSUBS 0.020237f
C149 VDD1.n119 VSUBS 0.020237f
C150 VDD1.n120 VSUBS 0.010875f
C151 VDD1.n121 VSUBS 0.011514f
C152 VDD1.n122 VSUBS 0.025704f
C153 VDD1.n123 VSUBS 0.025704f
C154 VDD1.n124 VSUBS 0.011514f
C155 VDD1.n125 VSUBS 0.010875f
C156 VDD1.n126 VSUBS 0.020237f
C157 VDD1.n127 VSUBS 0.020237f
C158 VDD1.n128 VSUBS 0.010875f
C159 VDD1.n129 VSUBS 0.010875f
C160 VDD1.n130 VSUBS 0.011514f
C161 VDD1.n131 VSUBS 0.025704f
C162 VDD1.n132 VSUBS 0.025704f
C163 VDD1.n133 VSUBS 0.025704f
C164 VDD1.n134 VSUBS 0.011195f
C165 VDD1.n135 VSUBS 0.010875f
C166 VDD1.n136 VSUBS 0.020237f
C167 VDD1.n137 VSUBS 0.020237f
C168 VDD1.n138 VSUBS 0.010875f
C169 VDD1.n139 VSUBS 0.011514f
C170 VDD1.n140 VSUBS 0.025704f
C171 VDD1.n141 VSUBS 0.025704f
C172 VDD1.n142 VSUBS 0.011514f
C173 VDD1.n143 VSUBS 0.010875f
C174 VDD1.n144 VSUBS 0.020237f
C175 VDD1.n145 VSUBS 0.020237f
C176 VDD1.n146 VSUBS 0.010875f
C177 VDD1.n147 VSUBS 0.011514f
C178 VDD1.n148 VSUBS 0.025704f
C179 VDD1.n149 VSUBS 0.025704f
C180 VDD1.n150 VSUBS 0.011514f
C181 VDD1.n151 VSUBS 0.010875f
C182 VDD1.n152 VSUBS 0.020237f
C183 VDD1.n153 VSUBS 0.020237f
C184 VDD1.n154 VSUBS 0.010875f
C185 VDD1.n155 VSUBS 0.011514f
C186 VDD1.n156 VSUBS 0.025704f
C187 VDD1.n157 VSUBS 0.025704f
C188 VDD1.n158 VSUBS 0.011514f
C189 VDD1.n159 VSUBS 0.010875f
C190 VDD1.n160 VSUBS 0.020237f
C191 VDD1.n161 VSUBS 0.020237f
C192 VDD1.n162 VSUBS 0.010875f
C193 VDD1.n163 VSUBS 0.011514f
C194 VDD1.n164 VSUBS 0.025704f
C195 VDD1.n165 VSUBS 0.06486f
C196 VDD1.n166 VSUBS 0.011514f
C197 VDD1.n167 VSUBS 0.010875f
C198 VDD1.n168 VSUBS 0.044013f
C199 VDD1.n169 VSUBS 0.687749f
C200 VP.t0 VSUBS 3.98135f
C201 VP.t1 VSUBS 3.61724f
C202 VP.n0 VSUBS 6.34921f
C203 VDD2.n0 VSUBS 0.022948f
C204 VDD2.n1 VSUBS 0.020183f
C205 VDD2.n2 VSUBS 0.010846f
C206 VDD2.n3 VSUBS 0.025635f
C207 VDD2.n4 VSUBS 0.011483f
C208 VDD2.n5 VSUBS 0.020183f
C209 VDD2.n6 VSUBS 0.010846f
C210 VDD2.n7 VSUBS 0.025635f
C211 VDD2.n8 VSUBS 0.011483f
C212 VDD2.n9 VSUBS 0.020183f
C213 VDD2.n10 VSUBS 0.010846f
C214 VDD2.n11 VSUBS 0.025635f
C215 VDD2.n12 VSUBS 0.011483f
C216 VDD2.n13 VSUBS 0.020183f
C217 VDD2.n14 VSUBS 0.010846f
C218 VDD2.n15 VSUBS 0.025635f
C219 VDD2.n16 VSUBS 0.011165f
C220 VDD2.n17 VSUBS 0.020183f
C221 VDD2.n18 VSUBS 0.011483f
C222 VDD2.n19 VSUBS 0.025635f
C223 VDD2.n20 VSUBS 0.011483f
C224 VDD2.n21 VSUBS 0.020183f
C225 VDD2.n22 VSUBS 0.010846f
C226 VDD2.n23 VSUBS 0.025635f
C227 VDD2.n24 VSUBS 0.011483f
C228 VDD2.n25 VSUBS 1.3118f
C229 VDD2.n26 VSUBS 0.010846f
C230 VDD2.t1 VSUBS 0.055485f
C231 VDD2.n27 VSUBS 0.191988f
C232 VDD2.n28 VSUBS 0.019284f
C233 VDD2.n29 VSUBS 0.019226f
C234 VDD2.n30 VSUBS 0.025635f
C235 VDD2.n31 VSUBS 0.011483f
C236 VDD2.n32 VSUBS 0.010846f
C237 VDD2.n33 VSUBS 0.020183f
C238 VDD2.n34 VSUBS 0.020183f
C239 VDD2.n35 VSUBS 0.010846f
C240 VDD2.n36 VSUBS 0.011483f
C241 VDD2.n37 VSUBS 0.025635f
C242 VDD2.n38 VSUBS 0.025635f
C243 VDD2.n39 VSUBS 0.011483f
C244 VDD2.n40 VSUBS 0.010846f
C245 VDD2.n41 VSUBS 0.020183f
C246 VDD2.n42 VSUBS 0.020183f
C247 VDD2.n43 VSUBS 0.010846f
C248 VDD2.n44 VSUBS 0.010846f
C249 VDD2.n45 VSUBS 0.011483f
C250 VDD2.n46 VSUBS 0.025635f
C251 VDD2.n47 VSUBS 0.025635f
C252 VDD2.n48 VSUBS 0.025635f
C253 VDD2.n49 VSUBS 0.011165f
C254 VDD2.n50 VSUBS 0.010846f
C255 VDD2.n51 VSUBS 0.020183f
C256 VDD2.n52 VSUBS 0.020183f
C257 VDD2.n53 VSUBS 0.010846f
C258 VDD2.n54 VSUBS 0.011483f
C259 VDD2.n55 VSUBS 0.025635f
C260 VDD2.n56 VSUBS 0.025635f
C261 VDD2.n57 VSUBS 0.011483f
C262 VDD2.n58 VSUBS 0.010846f
C263 VDD2.n59 VSUBS 0.020183f
C264 VDD2.n60 VSUBS 0.020183f
C265 VDD2.n61 VSUBS 0.010846f
C266 VDD2.n62 VSUBS 0.011483f
C267 VDD2.n63 VSUBS 0.025635f
C268 VDD2.n64 VSUBS 0.025635f
C269 VDD2.n65 VSUBS 0.011483f
C270 VDD2.n66 VSUBS 0.010846f
C271 VDD2.n67 VSUBS 0.020183f
C272 VDD2.n68 VSUBS 0.020183f
C273 VDD2.n69 VSUBS 0.010846f
C274 VDD2.n70 VSUBS 0.011483f
C275 VDD2.n71 VSUBS 0.025635f
C276 VDD2.n72 VSUBS 0.025635f
C277 VDD2.n73 VSUBS 0.011483f
C278 VDD2.n74 VSUBS 0.010846f
C279 VDD2.n75 VSUBS 0.020183f
C280 VDD2.n76 VSUBS 0.020183f
C281 VDD2.n77 VSUBS 0.010846f
C282 VDD2.n78 VSUBS 0.011483f
C283 VDD2.n79 VSUBS 0.025635f
C284 VDD2.n80 VSUBS 0.064686f
C285 VDD2.n81 VSUBS 0.011483f
C286 VDD2.n82 VSUBS 0.010846f
C287 VDD2.n83 VSUBS 0.043895f
C288 VDD2.n84 VSUBS 0.651612f
C289 VDD2.n85 VSUBS 0.022948f
C290 VDD2.n86 VSUBS 0.020183f
C291 VDD2.n87 VSUBS 0.010846f
C292 VDD2.n88 VSUBS 0.025635f
C293 VDD2.n89 VSUBS 0.011483f
C294 VDD2.n90 VSUBS 0.020183f
C295 VDD2.n91 VSUBS 0.010846f
C296 VDD2.n92 VSUBS 0.025635f
C297 VDD2.n93 VSUBS 0.011483f
C298 VDD2.n94 VSUBS 0.020183f
C299 VDD2.n95 VSUBS 0.010846f
C300 VDD2.n96 VSUBS 0.025635f
C301 VDD2.n97 VSUBS 0.011483f
C302 VDD2.n98 VSUBS 0.020183f
C303 VDD2.n99 VSUBS 0.010846f
C304 VDD2.n100 VSUBS 0.025635f
C305 VDD2.n101 VSUBS 0.011165f
C306 VDD2.n102 VSUBS 0.020183f
C307 VDD2.n103 VSUBS 0.011165f
C308 VDD2.n104 VSUBS 0.010846f
C309 VDD2.n105 VSUBS 0.025635f
C310 VDD2.n106 VSUBS 0.025635f
C311 VDD2.n107 VSUBS 0.011483f
C312 VDD2.n108 VSUBS 0.020183f
C313 VDD2.n109 VSUBS 0.010846f
C314 VDD2.n110 VSUBS 0.025635f
C315 VDD2.n111 VSUBS 0.011483f
C316 VDD2.n112 VSUBS 1.3118f
C317 VDD2.n113 VSUBS 0.010846f
C318 VDD2.t0 VSUBS 0.055485f
C319 VDD2.n114 VSUBS 0.191988f
C320 VDD2.n115 VSUBS 0.019284f
C321 VDD2.n116 VSUBS 0.019226f
C322 VDD2.n117 VSUBS 0.025635f
C323 VDD2.n118 VSUBS 0.011483f
C324 VDD2.n119 VSUBS 0.010846f
C325 VDD2.n120 VSUBS 0.020183f
C326 VDD2.n121 VSUBS 0.020183f
C327 VDD2.n122 VSUBS 0.010846f
C328 VDD2.n123 VSUBS 0.011483f
C329 VDD2.n124 VSUBS 0.025635f
C330 VDD2.n125 VSUBS 0.025635f
C331 VDD2.n126 VSUBS 0.011483f
C332 VDD2.n127 VSUBS 0.010846f
C333 VDD2.n128 VSUBS 0.020183f
C334 VDD2.n129 VSUBS 0.020183f
C335 VDD2.n130 VSUBS 0.010846f
C336 VDD2.n131 VSUBS 0.011483f
C337 VDD2.n132 VSUBS 0.025635f
C338 VDD2.n133 VSUBS 0.025635f
C339 VDD2.n134 VSUBS 0.011483f
C340 VDD2.n135 VSUBS 0.010846f
C341 VDD2.n136 VSUBS 0.020183f
C342 VDD2.n137 VSUBS 0.020183f
C343 VDD2.n138 VSUBS 0.010846f
C344 VDD2.n139 VSUBS 0.011483f
C345 VDD2.n140 VSUBS 0.025635f
C346 VDD2.n141 VSUBS 0.025635f
C347 VDD2.n142 VSUBS 0.011483f
C348 VDD2.n143 VSUBS 0.010846f
C349 VDD2.n144 VSUBS 0.020183f
C350 VDD2.n145 VSUBS 0.020183f
C351 VDD2.n146 VSUBS 0.010846f
C352 VDD2.n147 VSUBS 0.011483f
C353 VDD2.n148 VSUBS 0.025635f
C354 VDD2.n149 VSUBS 0.025635f
C355 VDD2.n150 VSUBS 0.011483f
C356 VDD2.n151 VSUBS 0.010846f
C357 VDD2.n152 VSUBS 0.020183f
C358 VDD2.n153 VSUBS 0.020183f
C359 VDD2.n154 VSUBS 0.010846f
C360 VDD2.n155 VSUBS 0.011483f
C361 VDD2.n156 VSUBS 0.025635f
C362 VDD2.n157 VSUBS 0.025635f
C363 VDD2.n158 VSUBS 0.011483f
C364 VDD2.n159 VSUBS 0.010846f
C365 VDD2.n160 VSUBS 0.020183f
C366 VDD2.n161 VSUBS 0.020183f
C367 VDD2.n162 VSUBS 0.010846f
C368 VDD2.n163 VSUBS 0.011483f
C369 VDD2.n164 VSUBS 0.025635f
C370 VDD2.n165 VSUBS 0.064686f
C371 VDD2.n166 VSUBS 0.011483f
C372 VDD2.n167 VSUBS 0.010846f
C373 VDD2.n168 VSUBS 0.043895f
C374 VDD2.n169 VSUBS 0.046519f
C375 VDD2.n170 VSUBS 2.57104f
C376 VTAIL.n0 VSUBS 0.031937f
C377 VTAIL.n1 VSUBS 0.028089f
C378 VTAIL.n2 VSUBS 0.015094f
C379 VTAIL.n3 VSUBS 0.035676f
C380 VTAIL.n4 VSUBS 0.015981f
C381 VTAIL.n5 VSUBS 0.028089f
C382 VTAIL.n6 VSUBS 0.015094f
C383 VTAIL.n7 VSUBS 0.035676f
C384 VTAIL.n8 VSUBS 0.015981f
C385 VTAIL.n9 VSUBS 0.028089f
C386 VTAIL.n10 VSUBS 0.015094f
C387 VTAIL.n11 VSUBS 0.035676f
C388 VTAIL.n12 VSUBS 0.015981f
C389 VTAIL.n13 VSUBS 0.028089f
C390 VTAIL.n14 VSUBS 0.015094f
C391 VTAIL.n15 VSUBS 0.035676f
C392 VTAIL.n16 VSUBS 0.015538f
C393 VTAIL.n17 VSUBS 0.028089f
C394 VTAIL.n18 VSUBS 0.015981f
C395 VTAIL.n19 VSUBS 0.035676f
C396 VTAIL.n20 VSUBS 0.015981f
C397 VTAIL.n21 VSUBS 0.028089f
C398 VTAIL.n22 VSUBS 0.015094f
C399 VTAIL.n23 VSUBS 0.035676f
C400 VTAIL.n24 VSUBS 0.015981f
C401 VTAIL.n25 VSUBS 1.82562f
C402 VTAIL.n26 VSUBS 0.015094f
C403 VTAIL.t3 VSUBS 0.077218f
C404 VTAIL.n27 VSUBS 0.267188f
C405 VTAIL.n28 VSUBS 0.026837f
C406 VTAIL.n29 VSUBS 0.026757f
C407 VTAIL.n30 VSUBS 0.035676f
C408 VTAIL.n31 VSUBS 0.015981f
C409 VTAIL.n32 VSUBS 0.015094f
C410 VTAIL.n33 VSUBS 0.028089f
C411 VTAIL.n34 VSUBS 0.028089f
C412 VTAIL.n35 VSUBS 0.015094f
C413 VTAIL.n36 VSUBS 0.015981f
C414 VTAIL.n37 VSUBS 0.035676f
C415 VTAIL.n38 VSUBS 0.035676f
C416 VTAIL.n39 VSUBS 0.015981f
C417 VTAIL.n40 VSUBS 0.015094f
C418 VTAIL.n41 VSUBS 0.028089f
C419 VTAIL.n42 VSUBS 0.028089f
C420 VTAIL.n43 VSUBS 0.015094f
C421 VTAIL.n44 VSUBS 0.015094f
C422 VTAIL.n45 VSUBS 0.015981f
C423 VTAIL.n46 VSUBS 0.035676f
C424 VTAIL.n47 VSUBS 0.035676f
C425 VTAIL.n48 VSUBS 0.035676f
C426 VTAIL.n49 VSUBS 0.015538f
C427 VTAIL.n50 VSUBS 0.015094f
C428 VTAIL.n51 VSUBS 0.028089f
C429 VTAIL.n52 VSUBS 0.028089f
C430 VTAIL.n53 VSUBS 0.015094f
C431 VTAIL.n54 VSUBS 0.015981f
C432 VTAIL.n55 VSUBS 0.035676f
C433 VTAIL.n56 VSUBS 0.035676f
C434 VTAIL.n57 VSUBS 0.015981f
C435 VTAIL.n58 VSUBS 0.015094f
C436 VTAIL.n59 VSUBS 0.028089f
C437 VTAIL.n60 VSUBS 0.028089f
C438 VTAIL.n61 VSUBS 0.015094f
C439 VTAIL.n62 VSUBS 0.015981f
C440 VTAIL.n63 VSUBS 0.035676f
C441 VTAIL.n64 VSUBS 0.035676f
C442 VTAIL.n65 VSUBS 0.015981f
C443 VTAIL.n66 VSUBS 0.015094f
C444 VTAIL.n67 VSUBS 0.028089f
C445 VTAIL.n68 VSUBS 0.028089f
C446 VTAIL.n69 VSUBS 0.015094f
C447 VTAIL.n70 VSUBS 0.015981f
C448 VTAIL.n71 VSUBS 0.035676f
C449 VTAIL.n72 VSUBS 0.035676f
C450 VTAIL.n73 VSUBS 0.015981f
C451 VTAIL.n74 VSUBS 0.015094f
C452 VTAIL.n75 VSUBS 0.028089f
C453 VTAIL.n76 VSUBS 0.028089f
C454 VTAIL.n77 VSUBS 0.015094f
C455 VTAIL.n78 VSUBS 0.015981f
C456 VTAIL.n79 VSUBS 0.035676f
C457 VTAIL.n80 VSUBS 0.090023f
C458 VTAIL.n81 VSUBS 0.015981f
C459 VTAIL.n82 VSUBS 0.015094f
C460 VTAIL.n83 VSUBS 0.061088f
C461 VTAIL.n84 VSUBS 0.045313f
C462 VTAIL.n85 VSUBS 1.98415f
C463 VTAIL.n86 VSUBS 0.031937f
C464 VTAIL.n87 VSUBS 0.028089f
C465 VTAIL.n88 VSUBS 0.015094f
C466 VTAIL.n89 VSUBS 0.035676f
C467 VTAIL.n90 VSUBS 0.015981f
C468 VTAIL.n91 VSUBS 0.028089f
C469 VTAIL.n92 VSUBS 0.015094f
C470 VTAIL.n93 VSUBS 0.035676f
C471 VTAIL.n94 VSUBS 0.015981f
C472 VTAIL.n95 VSUBS 0.028089f
C473 VTAIL.n96 VSUBS 0.015094f
C474 VTAIL.n97 VSUBS 0.035676f
C475 VTAIL.n98 VSUBS 0.015981f
C476 VTAIL.n99 VSUBS 0.028089f
C477 VTAIL.n100 VSUBS 0.015094f
C478 VTAIL.n101 VSUBS 0.035676f
C479 VTAIL.n102 VSUBS 0.015538f
C480 VTAIL.n103 VSUBS 0.028089f
C481 VTAIL.n104 VSUBS 0.015538f
C482 VTAIL.n105 VSUBS 0.015094f
C483 VTAIL.n106 VSUBS 0.035676f
C484 VTAIL.n107 VSUBS 0.035676f
C485 VTAIL.n108 VSUBS 0.015981f
C486 VTAIL.n109 VSUBS 0.028089f
C487 VTAIL.n110 VSUBS 0.015094f
C488 VTAIL.n111 VSUBS 0.035676f
C489 VTAIL.n112 VSUBS 0.015981f
C490 VTAIL.n113 VSUBS 1.82562f
C491 VTAIL.n114 VSUBS 0.015094f
C492 VTAIL.t1 VSUBS 0.077218f
C493 VTAIL.n115 VSUBS 0.267188f
C494 VTAIL.n116 VSUBS 0.026837f
C495 VTAIL.n117 VSUBS 0.026757f
C496 VTAIL.n118 VSUBS 0.035676f
C497 VTAIL.n119 VSUBS 0.015981f
C498 VTAIL.n120 VSUBS 0.015094f
C499 VTAIL.n121 VSUBS 0.028089f
C500 VTAIL.n122 VSUBS 0.028089f
C501 VTAIL.n123 VSUBS 0.015094f
C502 VTAIL.n124 VSUBS 0.015981f
C503 VTAIL.n125 VSUBS 0.035676f
C504 VTAIL.n126 VSUBS 0.035676f
C505 VTAIL.n127 VSUBS 0.015981f
C506 VTAIL.n128 VSUBS 0.015094f
C507 VTAIL.n129 VSUBS 0.028089f
C508 VTAIL.n130 VSUBS 0.028089f
C509 VTAIL.n131 VSUBS 0.015094f
C510 VTAIL.n132 VSUBS 0.015981f
C511 VTAIL.n133 VSUBS 0.035676f
C512 VTAIL.n134 VSUBS 0.035676f
C513 VTAIL.n135 VSUBS 0.015981f
C514 VTAIL.n136 VSUBS 0.015094f
C515 VTAIL.n137 VSUBS 0.028089f
C516 VTAIL.n138 VSUBS 0.028089f
C517 VTAIL.n139 VSUBS 0.015094f
C518 VTAIL.n140 VSUBS 0.015981f
C519 VTAIL.n141 VSUBS 0.035676f
C520 VTAIL.n142 VSUBS 0.035676f
C521 VTAIL.n143 VSUBS 0.015981f
C522 VTAIL.n144 VSUBS 0.015094f
C523 VTAIL.n145 VSUBS 0.028089f
C524 VTAIL.n146 VSUBS 0.028089f
C525 VTAIL.n147 VSUBS 0.015094f
C526 VTAIL.n148 VSUBS 0.015981f
C527 VTAIL.n149 VSUBS 0.035676f
C528 VTAIL.n150 VSUBS 0.035676f
C529 VTAIL.n151 VSUBS 0.015981f
C530 VTAIL.n152 VSUBS 0.015094f
C531 VTAIL.n153 VSUBS 0.028089f
C532 VTAIL.n154 VSUBS 0.028089f
C533 VTAIL.n155 VSUBS 0.015094f
C534 VTAIL.n156 VSUBS 0.015981f
C535 VTAIL.n157 VSUBS 0.035676f
C536 VTAIL.n158 VSUBS 0.035676f
C537 VTAIL.n159 VSUBS 0.015981f
C538 VTAIL.n160 VSUBS 0.015094f
C539 VTAIL.n161 VSUBS 0.028089f
C540 VTAIL.n162 VSUBS 0.028089f
C541 VTAIL.n163 VSUBS 0.015094f
C542 VTAIL.n164 VSUBS 0.015981f
C543 VTAIL.n165 VSUBS 0.035676f
C544 VTAIL.n166 VSUBS 0.090023f
C545 VTAIL.n167 VSUBS 0.015981f
C546 VTAIL.n168 VSUBS 0.015094f
C547 VTAIL.n169 VSUBS 0.061088f
C548 VTAIL.n170 VSUBS 0.045313f
C549 VTAIL.n171 VSUBS 2.0138f
C550 VTAIL.n172 VSUBS 0.031937f
C551 VTAIL.n173 VSUBS 0.028089f
C552 VTAIL.n174 VSUBS 0.015094f
C553 VTAIL.n175 VSUBS 0.035676f
C554 VTAIL.n176 VSUBS 0.015981f
C555 VTAIL.n177 VSUBS 0.028089f
C556 VTAIL.n178 VSUBS 0.015094f
C557 VTAIL.n179 VSUBS 0.035676f
C558 VTAIL.n180 VSUBS 0.015981f
C559 VTAIL.n181 VSUBS 0.028089f
C560 VTAIL.n182 VSUBS 0.015094f
C561 VTAIL.n183 VSUBS 0.035676f
C562 VTAIL.n184 VSUBS 0.015981f
C563 VTAIL.n185 VSUBS 0.028089f
C564 VTAIL.n186 VSUBS 0.015094f
C565 VTAIL.n187 VSUBS 0.035676f
C566 VTAIL.n188 VSUBS 0.015538f
C567 VTAIL.n189 VSUBS 0.028089f
C568 VTAIL.n190 VSUBS 0.015538f
C569 VTAIL.n191 VSUBS 0.015094f
C570 VTAIL.n192 VSUBS 0.035676f
C571 VTAIL.n193 VSUBS 0.035676f
C572 VTAIL.n194 VSUBS 0.015981f
C573 VTAIL.n195 VSUBS 0.028089f
C574 VTAIL.n196 VSUBS 0.015094f
C575 VTAIL.n197 VSUBS 0.035676f
C576 VTAIL.n198 VSUBS 0.015981f
C577 VTAIL.n199 VSUBS 1.82562f
C578 VTAIL.n200 VSUBS 0.015094f
C579 VTAIL.t0 VSUBS 0.077218f
C580 VTAIL.n201 VSUBS 0.267188f
C581 VTAIL.n202 VSUBS 0.026837f
C582 VTAIL.n203 VSUBS 0.026757f
C583 VTAIL.n204 VSUBS 0.035676f
C584 VTAIL.n205 VSUBS 0.015981f
C585 VTAIL.n206 VSUBS 0.015094f
C586 VTAIL.n207 VSUBS 0.028089f
C587 VTAIL.n208 VSUBS 0.028089f
C588 VTAIL.n209 VSUBS 0.015094f
C589 VTAIL.n210 VSUBS 0.015981f
C590 VTAIL.n211 VSUBS 0.035676f
C591 VTAIL.n212 VSUBS 0.035676f
C592 VTAIL.n213 VSUBS 0.015981f
C593 VTAIL.n214 VSUBS 0.015094f
C594 VTAIL.n215 VSUBS 0.028089f
C595 VTAIL.n216 VSUBS 0.028089f
C596 VTAIL.n217 VSUBS 0.015094f
C597 VTAIL.n218 VSUBS 0.015981f
C598 VTAIL.n219 VSUBS 0.035676f
C599 VTAIL.n220 VSUBS 0.035676f
C600 VTAIL.n221 VSUBS 0.015981f
C601 VTAIL.n222 VSUBS 0.015094f
C602 VTAIL.n223 VSUBS 0.028089f
C603 VTAIL.n224 VSUBS 0.028089f
C604 VTAIL.n225 VSUBS 0.015094f
C605 VTAIL.n226 VSUBS 0.015981f
C606 VTAIL.n227 VSUBS 0.035676f
C607 VTAIL.n228 VSUBS 0.035676f
C608 VTAIL.n229 VSUBS 0.015981f
C609 VTAIL.n230 VSUBS 0.015094f
C610 VTAIL.n231 VSUBS 0.028089f
C611 VTAIL.n232 VSUBS 0.028089f
C612 VTAIL.n233 VSUBS 0.015094f
C613 VTAIL.n234 VSUBS 0.015981f
C614 VTAIL.n235 VSUBS 0.035676f
C615 VTAIL.n236 VSUBS 0.035676f
C616 VTAIL.n237 VSUBS 0.015981f
C617 VTAIL.n238 VSUBS 0.015094f
C618 VTAIL.n239 VSUBS 0.028089f
C619 VTAIL.n240 VSUBS 0.028089f
C620 VTAIL.n241 VSUBS 0.015094f
C621 VTAIL.n242 VSUBS 0.015981f
C622 VTAIL.n243 VSUBS 0.035676f
C623 VTAIL.n244 VSUBS 0.035676f
C624 VTAIL.n245 VSUBS 0.015981f
C625 VTAIL.n246 VSUBS 0.015094f
C626 VTAIL.n247 VSUBS 0.028089f
C627 VTAIL.n248 VSUBS 0.028089f
C628 VTAIL.n249 VSUBS 0.015094f
C629 VTAIL.n250 VSUBS 0.015981f
C630 VTAIL.n251 VSUBS 0.035676f
C631 VTAIL.n252 VSUBS 0.090023f
C632 VTAIL.n253 VSUBS 0.015981f
C633 VTAIL.n254 VSUBS 0.015094f
C634 VTAIL.n255 VSUBS 0.061088f
C635 VTAIL.n256 VSUBS 0.045313f
C636 VTAIL.n257 VSUBS 1.87413f
C637 VTAIL.n258 VSUBS 0.031937f
C638 VTAIL.n259 VSUBS 0.028089f
C639 VTAIL.n260 VSUBS 0.015094f
C640 VTAIL.n261 VSUBS 0.035676f
C641 VTAIL.n262 VSUBS 0.015981f
C642 VTAIL.n263 VSUBS 0.028089f
C643 VTAIL.n264 VSUBS 0.015094f
C644 VTAIL.n265 VSUBS 0.035676f
C645 VTAIL.n266 VSUBS 0.015981f
C646 VTAIL.n267 VSUBS 0.028089f
C647 VTAIL.n268 VSUBS 0.015094f
C648 VTAIL.n269 VSUBS 0.035676f
C649 VTAIL.n270 VSUBS 0.015981f
C650 VTAIL.n271 VSUBS 0.028089f
C651 VTAIL.n272 VSUBS 0.015094f
C652 VTAIL.n273 VSUBS 0.035676f
C653 VTAIL.n274 VSUBS 0.015538f
C654 VTAIL.n275 VSUBS 0.028089f
C655 VTAIL.n276 VSUBS 0.015981f
C656 VTAIL.n277 VSUBS 0.035676f
C657 VTAIL.n278 VSUBS 0.015981f
C658 VTAIL.n279 VSUBS 0.028089f
C659 VTAIL.n280 VSUBS 0.015094f
C660 VTAIL.n281 VSUBS 0.035676f
C661 VTAIL.n282 VSUBS 0.015981f
C662 VTAIL.n283 VSUBS 1.82562f
C663 VTAIL.n284 VSUBS 0.015094f
C664 VTAIL.t2 VSUBS 0.077218f
C665 VTAIL.n285 VSUBS 0.267188f
C666 VTAIL.n286 VSUBS 0.026837f
C667 VTAIL.n287 VSUBS 0.026757f
C668 VTAIL.n288 VSUBS 0.035676f
C669 VTAIL.n289 VSUBS 0.015981f
C670 VTAIL.n290 VSUBS 0.015094f
C671 VTAIL.n291 VSUBS 0.028089f
C672 VTAIL.n292 VSUBS 0.028089f
C673 VTAIL.n293 VSUBS 0.015094f
C674 VTAIL.n294 VSUBS 0.015981f
C675 VTAIL.n295 VSUBS 0.035676f
C676 VTAIL.n296 VSUBS 0.035676f
C677 VTAIL.n297 VSUBS 0.015981f
C678 VTAIL.n298 VSUBS 0.015094f
C679 VTAIL.n299 VSUBS 0.028089f
C680 VTAIL.n300 VSUBS 0.028089f
C681 VTAIL.n301 VSUBS 0.015094f
C682 VTAIL.n302 VSUBS 0.015094f
C683 VTAIL.n303 VSUBS 0.015981f
C684 VTAIL.n304 VSUBS 0.035676f
C685 VTAIL.n305 VSUBS 0.035676f
C686 VTAIL.n306 VSUBS 0.035676f
C687 VTAIL.n307 VSUBS 0.015538f
C688 VTAIL.n308 VSUBS 0.015094f
C689 VTAIL.n309 VSUBS 0.028089f
C690 VTAIL.n310 VSUBS 0.028089f
C691 VTAIL.n311 VSUBS 0.015094f
C692 VTAIL.n312 VSUBS 0.015981f
C693 VTAIL.n313 VSUBS 0.035676f
C694 VTAIL.n314 VSUBS 0.035676f
C695 VTAIL.n315 VSUBS 0.015981f
C696 VTAIL.n316 VSUBS 0.015094f
C697 VTAIL.n317 VSUBS 0.028089f
C698 VTAIL.n318 VSUBS 0.028089f
C699 VTAIL.n319 VSUBS 0.015094f
C700 VTAIL.n320 VSUBS 0.015981f
C701 VTAIL.n321 VSUBS 0.035676f
C702 VTAIL.n322 VSUBS 0.035676f
C703 VTAIL.n323 VSUBS 0.015981f
C704 VTAIL.n324 VSUBS 0.015094f
C705 VTAIL.n325 VSUBS 0.028089f
C706 VTAIL.n326 VSUBS 0.028089f
C707 VTAIL.n327 VSUBS 0.015094f
C708 VTAIL.n328 VSUBS 0.015981f
C709 VTAIL.n329 VSUBS 0.035676f
C710 VTAIL.n330 VSUBS 0.035676f
C711 VTAIL.n331 VSUBS 0.015981f
C712 VTAIL.n332 VSUBS 0.015094f
C713 VTAIL.n333 VSUBS 0.028089f
C714 VTAIL.n334 VSUBS 0.028089f
C715 VTAIL.n335 VSUBS 0.015094f
C716 VTAIL.n336 VSUBS 0.015981f
C717 VTAIL.n337 VSUBS 0.035676f
C718 VTAIL.n338 VSUBS 0.090023f
C719 VTAIL.n339 VSUBS 0.015981f
C720 VTAIL.n340 VSUBS 0.015094f
C721 VTAIL.n341 VSUBS 0.061088f
C722 VTAIL.n342 VSUBS 0.045313f
C723 VTAIL.n343 VSUBS 1.79143f
C724 VN.t0 VSUBS 3.52191f
C725 VN.t1 VSUBS 3.88104f
C726 B.n0 VSUBS 0.005589f
C727 B.n1 VSUBS 0.005589f
C728 B.n2 VSUBS 0.008266f
C729 B.n3 VSUBS 0.006334f
C730 B.n4 VSUBS 0.006334f
C731 B.n5 VSUBS 0.006334f
C732 B.n6 VSUBS 0.006334f
C733 B.n7 VSUBS 0.006334f
C734 B.n8 VSUBS 0.006334f
C735 B.n9 VSUBS 0.006334f
C736 B.n10 VSUBS 0.006334f
C737 B.n11 VSUBS 0.015759f
C738 B.n12 VSUBS 0.006334f
C739 B.n13 VSUBS 0.006334f
C740 B.n14 VSUBS 0.006334f
C741 B.n15 VSUBS 0.006334f
C742 B.n16 VSUBS 0.006334f
C743 B.n17 VSUBS 0.006334f
C744 B.n18 VSUBS 0.006334f
C745 B.n19 VSUBS 0.006334f
C746 B.n20 VSUBS 0.006334f
C747 B.n21 VSUBS 0.006334f
C748 B.n22 VSUBS 0.006334f
C749 B.n23 VSUBS 0.006334f
C750 B.n24 VSUBS 0.006334f
C751 B.n25 VSUBS 0.006334f
C752 B.n26 VSUBS 0.006334f
C753 B.n27 VSUBS 0.006334f
C754 B.n28 VSUBS 0.006334f
C755 B.n29 VSUBS 0.006334f
C756 B.n30 VSUBS 0.006334f
C757 B.n31 VSUBS 0.006334f
C758 B.n32 VSUBS 0.006334f
C759 B.n33 VSUBS 0.006334f
C760 B.n34 VSUBS 0.006334f
C761 B.n35 VSUBS 0.006334f
C762 B.n36 VSUBS 0.006334f
C763 B.n37 VSUBS 0.006334f
C764 B.t4 VSUBS 0.266426f
C765 B.t5 VSUBS 0.28522f
C766 B.t3 VSUBS 0.884334f
C767 B.n38 VSUBS 0.409092f
C768 B.n39 VSUBS 0.266592f
C769 B.n40 VSUBS 0.006334f
C770 B.n41 VSUBS 0.006334f
C771 B.n42 VSUBS 0.006334f
C772 B.n43 VSUBS 0.006334f
C773 B.t1 VSUBS 0.266429f
C774 B.t2 VSUBS 0.285222f
C775 B.t0 VSUBS 0.884334f
C776 B.n44 VSUBS 0.40909f
C777 B.n45 VSUBS 0.266589f
C778 B.n46 VSUBS 0.014676f
C779 B.n47 VSUBS 0.006334f
C780 B.n48 VSUBS 0.006334f
C781 B.n49 VSUBS 0.006334f
C782 B.n50 VSUBS 0.006334f
C783 B.n51 VSUBS 0.006334f
C784 B.n52 VSUBS 0.006334f
C785 B.n53 VSUBS 0.006334f
C786 B.n54 VSUBS 0.006334f
C787 B.n55 VSUBS 0.006334f
C788 B.n56 VSUBS 0.006334f
C789 B.n57 VSUBS 0.006334f
C790 B.n58 VSUBS 0.006334f
C791 B.n59 VSUBS 0.006334f
C792 B.n60 VSUBS 0.006334f
C793 B.n61 VSUBS 0.006334f
C794 B.n62 VSUBS 0.006334f
C795 B.n63 VSUBS 0.006334f
C796 B.n64 VSUBS 0.006334f
C797 B.n65 VSUBS 0.006334f
C798 B.n66 VSUBS 0.006334f
C799 B.n67 VSUBS 0.006334f
C800 B.n68 VSUBS 0.006334f
C801 B.n69 VSUBS 0.006334f
C802 B.n70 VSUBS 0.006334f
C803 B.n71 VSUBS 0.006334f
C804 B.n72 VSUBS 0.015759f
C805 B.n73 VSUBS 0.006334f
C806 B.n74 VSUBS 0.006334f
C807 B.n75 VSUBS 0.006334f
C808 B.n76 VSUBS 0.006334f
C809 B.n77 VSUBS 0.006334f
C810 B.n78 VSUBS 0.006334f
C811 B.n79 VSUBS 0.006334f
C812 B.n80 VSUBS 0.006334f
C813 B.n81 VSUBS 0.006334f
C814 B.n82 VSUBS 0.006334f
C815 B.n83 VSUBS 0.006334f
C816 B.n84 VSUBS 0.006334f
C817 B.n85 VSUBS 0.006334f
C818 B.n86 VSUBS 0.006334f
C819 B.n87 VSUBS 0.006334f
C820 B.n88 VSUBS 0.006334f
C821 B.n89 VSUBS 0.006334f
C822 B.n90 VSUBS 0.006334f
C823 B.n91 VSUBS 0.014982f
C824 B.n92 VSUBS 0.006334f
C825 B.n93 VSUBS 0.006334f
C826 B.n94 VSUBS 0.006334f
C827 B.n95 VSUBS 0.006334f
C828 B.n96 VSUBS 0.006334f
C829 B.n97 VSUBS 0.006334f
C830 B.n98 VSUBS 0.006334f
C831 B.n99 VSUBS 0.006334f
C832 B.n100 VSUBS 0.006334f
C833 B.n101 VSUBS 0.006334f
C834 B.n102 VSUBS 0.006334f
C835 B.n103 VSUBS 0.006334f
C836 B.n104 VSUBS 0.006334f
C837 B.n105 VSUBS 0.006334f
C838 B.n106 VSUBS 0.006334f
C839 B.n107 VSUBS 0.006334f
C840 B.n108 VSUBS 0.006334f
C841 B.n109 VSUBS 0.006334f
C842 B.n110 VSUBS 0.006334f
C843 B.n111 VSUBS 0.006334f
C844 B.n112 VSUBS 0.006334f
C845 B.n113 VSUBS 0.006334f
C846 B.n114 VSUBS 0.006334f
C847 B.n115 VSUBS 0.006334f
C848 B.n116 VSUBS 0.006334f
C849 B.n117 VSUBS 0.006334f
C850 B.t8 VSUBS 0.266429f
C851 B.t7 VSUBS 0.285222f
C852 B.t6 VSUBS 0.884334f
C853 B.n118 VSUBS 0.40909f
C854 B.n119 VSUBS 0.266589f
C855 B.n120 VSUBS 0.006334f
C856 B.n121 VSUBS 0.006334f
C857 B.n122 VSUBS 0.006334f
C858 B.n123 VSUBS 0.006334f
C859 B.n124 VSUBS 0.00354f
C860 B.n125 VSUBS 0.006334f
C861 B.n126 VSUBS 0.006334f
C862 B.n127 VSUBS 0.006334f
C863 B.n128 VSUBS 0.006334f
C864 B.n129 VSUBS 0.006334f
C865 B.n130 VSUBS 0.006334f
C866 B.n131 VSUBS 0.006334f
C867 B.n132 VSUBS 0.006334f
C868 B.n133 VSUBS 0.006334f
C869 B.n134 VSUBS 0.006334f
C870 B.n135 VSUBS 0.006334f
C871 B.n136 VSUBS 0.006334f
C872 B.n137 VSUBS 0.006334f
C873 B.n138 VSUBS 0.006334f
C874 B.n139 VSUBS 0.006334f
C875 B.n140 VSUBS 0.006334f
C876 B.n141 VSUBS 0.006334f
C877 B.n142 VSUBS 0.006334f
C878 B.n143 VSUBS 0.006334f
C879 B.n144 VSUBS 0.006334f
C880 B.n145 VSUBS 0.006334f
C881 B.n146 VSUBS 0.006334f
C882 B.n147 VSUBS 0.006334f
C883 B.n148 VSUBS 0.006334f
C884 B.n149 VSUBS 0.006334f
C885 B.n150 VSUBS 0.015759f
C886 B.n151 VSUBS 0.006334f
C887 B.n152 VSUBS 0.006334f
C888 B.n153 VSUBS 0.006334f
C889 B.n154 VSUBS 0.006334f
C890 B.n155 VSUBS 0.006334f
C891 B.n156 VSUBS 0.006334f
C892 B.n157 VSUBS 0.006334f
C893 B.n158 VSUBS 0.006334f
C894 B.n159 VSUBS 0.006334f
C895 B.n160 VSUBS 0.006334f
C896 B.n161 VSUBS 0.006334f
C897 B.n162 VSUBS 0.006334f
C898 B.n163 VSUBS 0.006334f
C899 B.n164 VSUBS 0.006334f
C900 B.n165 VSUBS 0.006334f
C901 B.n166 VSUBS 0.006334f
C902 B.n167 VSUBS 0.006334f
C903 B.n168 VSUBS 0.006334f
C904 B.n169 VSUBS 0.006334f
C905 B.n170 VSUBS 0.006334f
C906 B.n171 VSUBS 0.006334f
C907 B.n172 VSUBS 0.006334f
C908 B.n173 VSUBS 0.006334f
C909 B.n174 VSUBS 0.006334f
C910 B.n175 VSUBS 0.006334f
C911 B.n176 VSUBS 0.006334f
C912 B.n177 VSUBS 0.006334f
C913 B.n178 VSUBS 0.006334f
C914 B.n179 VSUBS 0.006334f
C915 B.n180 VSUBS 0.006334f
C916 B.n181 VSUBS 0.006334f
C917 B.n182 VSUBS 0.006334f
C918 B.n183 VSUBS 0.014982f
C919 B.n184 VSUBS 0.014982f
C920 B.n185 VSUBS 0.015759f
C921 B.n186 VSUBS 0.006334f
C922 B.n187 VSUBS 0.006334f
C923 B.n188 VSUBS 0.006334f
C924 B.n189 VSUBS 0.006334f
C925 B.n190 VSUBS 0.006334f
C926 B.n191 VSUBS 0.006334f
C927 B.n192 VSUBS 0.006334f
C928 B.n193 VSUBS 0.006334f
C929 B.n194 VSUBS 0.006334f
C930 B.n195 VSUBS 0.006334f
C931 B.n196 VSUBS 0.006334f
C932 B.n197 VSUBS 0.006334f
C933 B.n198 VSUBS 0.006334f
C934 B.n199 VSUBS 0.006334f
C935 B.n200 VSUBS 0.006334f
C936 B.n201 VSUBS 0.006334f
C937 B.n202 VSUBS 0.006334f
C938 B.n203 VSUBS 0.006334f
C939 B.n204 VSUBS 0.006334f
C940 B.n205 VSUBS 0.006334f
C941 B.n206 VSUBS 0.006334f
C942 B.n207 VSUBS 0.006334f
C943 B.n208 VSUBS 0.006334f
C944 B.n209 VSUBS 0.006334f
C945 B.n210 VSUBS 0.006334f
C946 B.n211 VSUBS 0.006334f
C947 B.n212 VSUBS 0.006334f
C948 B.n213 VSUBS 0.006334f
C949 B.n214 VSUBS 0.006334f
C950 B.n215 VSUBS 0.006334f
C951 B.n216 VSUBS 0.006334f
C952 B.n217 VSUBS 0.006334f
C953 B.n218 VSUBS 0.006334f
C954 B.n219 VSUBS 0.006334f
C955 B.n220 VSUBS 0.006334f
C956 B.n221 VSUBS 0.006334f
C957 B.n222 VSUBS 0.006334f
C958 B.n223 VSUBS 0.006334f
C959 B.n224 VSUBS 0.006334f
C960 B.n225 VSUBS 0.006334f
C961 B.n226 VSUBS 0.006334f
C962 B.n227 VSUBS 0.006334f
C963 B.n228 VSUBS 0.006334f
C964 B.n229 VSUBS 0.006334f
C965 B.n230 VSUBS 0.006334f
C966 B.n231 VSUBS 0.006334f
C967 B.n232 VSUBS 0.006334f
C968 B.n233 VSUBS 0.006334f
C969 B.n234 VSUBS 0.006334f
C970 B.n235 VSUBS 0.006334f
C971 B.n236 VSUBS 0.006334f
C972 B.n237 VSUBS 0.006334f
C973 B.n238 VSUBS 0.006334f
C974 B.n239 VSUBS 0.006334f
C975 B.n240 VSUBS 0.006334f
C976 B.n241 VSUBS 0.006334f
C977 B.n242 VSUBS 0.006334f
C978 B.n243 VSUBS 0.006334f
C979 B.n244 VSUBS 0.006334f
C980 B.n245 VSUBS 0.006334f
C981 B.n246 VSUBS 0.006334f
C982 B.n247 VSUBS 0.006334f
C983 B.n248 VSUBS 0.006334f
C984 B.n249 VSUBS 0.006334f
C985 B.n250 VSUBS 0.006334f
C986 B.n251 VSUBS 0.006334f
C987 B.n252 VSUBS 0.006334f
C988 B.n253 VSUBS 0.006334f
C989 B.n254 VSUBS 0.006334f
C990 B.n255 VSUBS 0.006334f
C991 B.n256 VSUBS 0.006334f
C992 B.n257 VSUBS 0.006334f
C993 B.n258 VSUBS 0.006334f
C994 B.n259 VSUBS 0.006334f
C995 B.n260 VSUBS 0.006334f
C996 B.t11 VSUBS 0.266426f
C997 B.t10 VSUBS 0.28522f
C998 B.t9 VSUBS 0.884334f
C999 B.n261 VSUBS 0.409092f
C1000 B.n262 VSUBS 0.266592f
C1001 B.n263 VSUBS 0.014676f
C1002 B.n264 VSUBS 0.005962f
C1003 B.n265 VSUBS 0.006334f
C1004 B.n266 VSUBS 0.006334f
C1005 B.n267 VSUBS 0.006334f
C1006 B.n268 VSUBS 0.006334f
C1007 B.n269 VSUBS 0.006334f
C1008 B.n270 VSUBS 0.006334f
C1009 B.n271 VSUBS 0.006334f
C1010 B.n272 VSUBS 0.006334f
C1011 B.n273 VSUBS 0.006334f
C1012 B.n274 VSUBS 0.006334f
C1013 B.n275 VSUBS 0.006334f
C1014 B.n276 VSUBS 0.006334f
C1015 B.n277 VSUBS 0.006334f
C1016 B.n278 VSUBS 0.006334f
C1017 B.n279 VSUBS 0.006334f
C1018 B.n280 VSUBS 0.00354f
C1019 B.n281 VSUBS 0.014676f
C1020 B.n282 VSUBS 0.005962f
C1021 B.n283 VSUBS 0.006334f
C1022 B.n284 VSUBS 0.006334f
C1023 B.n285 VSUBS 0.006334f
C1024 B.n286 VSUBS 0.006334f
C1025 B.n287 VSUBS 0.006334f
C1026 B.n288 VSUBS 0.006334f
C1027 B.n289 VSUBS 0.006334f
C1028 B.n290 VSUBS 0.006334f
C1029 B.n291 VSUBS 0.006334f
C1030 B.n292 VSUBS 0.006334f
C1031 B.n293 VSUBS 0.006334f
C1032 B.n294 VSUBS 0.006334f
C1033 B.n295 VSUBS 0.006334f
C1034 B.n296 VSUBS 0.006334f
C1035 B.n297 VSUBS 0.006334f
C1036 B.n298 VSUBS 0.006334f
C1037 B.n299 VSUBS 0.006334f
C1038 B.n300 VSUBS 0.006334f
C1039 B.n301 VSUBS 0.006334f
C1040 B.n302 VSUBS 0.006334f
C1041 B.n303 VSUBS 0.006334f
C1042 B.n304 VSUBS 0.006334f
C1043 B.n305 VSUBS 0.006334f
C1044 B.n306 VSUBS 0.006334f
C1045 B.n307 VSUBS 0.006334f
C1046 B.n308 VSUBS 0.006334f
C1047 B.n309 VSUBS 0.006334f
C1048 B.n310 VSUBS 0.006334f
C1049 B.n311 VSUBS 0.006334f
C1050 B.n312 VSUBS 0.006334f
C1051 B.n313 VSUBS 0.006334f
C1052 B.n314 VSUBS 0.006334f
C1053 B.n315 VSUBS 0.006334f
C1054 B.n316 VSUBS 0.006334f
C1055 B.n317 VSUBS 0.006334f
C1056 B.n318 VSUBS 0.006334f
C1057 B.n319 VSUBS 0.006334f
C1058 B.n320 VSUBS 0.006334f
C1059 B.n321 VSUBS 0.006334f
C1060 B.n322 VSUBS 0.006334f
C1061 B.n323 VSUBS 0.006334f
C1062 B.n324 VSUBS 0.006334f
C1063 B.n325 VSUBS 0.006334f
C1064 B.n326 VSUBS 0.006334f
C1065 B.n327 VSUBS 0.006334f
C1066 B.n328 VSUBS 0.006334f
C1067 B.n329 VSUBS 0.006334f
C1068 B.n330 VSUBS 0.006334f
C1069 B.n331 VSUBS 0.006334f
C1070 B.n332 VSUBS 0.006334f
C1071 B.n333 VSUBS 0.006334f
C1072 B.n334 VSUBS 0.006334f
C1073 B.n335 VSUBS 0.006334f
C1074 B.n336 VSUBS 0.006334f
C1075 B.n337 VSUBS 0.006334f
C1076 B.n338 VSUBS 0.006334f
C1077 B.n339 VSUBS 0.006334f
C1078 B.n340 VSUBS 0.006334f
C1079 B.n341 VSUBS 0.006334f
C1080 B.n342 VSUBS 0.006334f
C1081 B.n343 VSUBS 0.006334f
C1082 B.n344 VSUBS 0.006334f
C1083 B.n345 VSUBS 0.006334f
C1084 B.n346 VSUBS 0.006334f
C1085 B.n347 VSUBS 0.006334f
C1086 B.n348 VSUBS 0.006334f
C1087 B.n349 VSUBS 0.006334f
C1088 B.n350 VSUBS 0.006334f
C1089 B.n351 VSUBS 0.006334f
C1090 B.n352 VSUBS 0.006334f
C1091 B.n353 VSUBS 0.006334f
C1092 B.n354 VSUBS 0.006334f
C1093 B.n355 VSUBS 0.006334f
C1094 B.n356 VSUBS 0.006334f
C1095 B.n357 VSUBS 0.006334f
C1096 B.n358 VSUBS 0.015759f
C1097 B.n359 VSUBS 0.015051f
C1098 B.n360 VSUBS 0.01569f
C1099 B.n361 VSUBS 0.006334f
C1100 B.n362 VSUBS 0.006334f
C1101 B.n363 VSUBS 0.006334f
C1102 B.n364 VSUBS 0.006334f
C1103 B.n365 VSUBS 0.006334f
C1104 B.n366 VSUBS 0.006334f
C1105 B.n367 VSUBS 0.006334f
C1106 B.n368 VSUBS 0.006334f
C1107 B.n369 VSUBS 0.006334f
C1108 B.n370 VSUBS 0.006334f
C1109 B.n371 VSUBS 0.006334f
C1110 B.n372 VSUBS 0.006334f
C1111 B.n373 VSUBS 0.006334f
C1112 B.n374 VSUBS 0.006334f
C1113 B.n375 VSUBS 0.006334f
C1114 B.n376 VSUBS 0.006334f
C1115 B.n377 VSUBS 0.006334f
C1116 B.n378 VSUBS 0.006334f
C1117 B.n379 VSUBS 0.006334f
C1118 B.n380 VSUBS 0.006334f
C1119 B.n381 VSUBS 0.006334f
C1120 B.n382 VSUBS 0.006334f
C1121 B.n383 VSUBS 0.006334f
C1122 B.n384 VSUBS 0.006334f
C1123 B.n385 VSUBS 0.006334f
C1124 B.n386 VSUBS 0.006334f
C1125 B.n387 VSUBS 0.006334f
C1126 B.n388 VSUBS 0.006334f
C1127 B.n389 VSUBS 0.006334f
C1128 B.n390 VSUBS 0.006334f
C1129 B.n391 VSUBS 0.006334f
C1130 B.n392 VSUBS 0.006334f
C1131 B.n393 VSUBS 0.006334f
C1132 B.n394 VSUBS 0.006334f
C1133 B.n395 VSUBS 0.006334f
C1134 B.n396 VSUBS 0.006334f
C1135 B.n397 VSUBS 0.006334f
C1136 B.n398 VSUBS 0.006334f
C1137 B.n399 VSUBS 0.006334f
C1138 B.n400 VSUBS 0.006334f
C1139 B.n401 VSUBS 0.006334f
C1140 B.n402 VSUBS 0.006334f
C1141 B.n403 VSUBS 0.006334f
C1142 B.n404 VSUBS 0.006334f
C1143 B.n405 VSUBS 0.006334f
C1144 B.n406 VSUBS 0.006334f
C1145 B.n407 VSUBS 0.006334f
C1146 B.n408 VSUBS 0.006334f
C1147 B.n409 VSUBS 0.006334f
C1148 B.n410 VSUBS 0.006334f
C1149 B.n411 VSUBS 0.006334f
C1150 B.n412 VSUBS 0.006334f
C1151 B.n413 VSUBS 0.006334f
C1152 B.n414 VSUBS 0.006334f
C1153 B.n415 VSUBS 0.014982f
C1154 B.n416 VSUBS 0.014982f
C1155 B.n417 VSUBS 0.015759f
C1156 B.n418 VSUBS 0.006334f
C1157 B.n419 VSUBS 0.006334f
C1158 B.n420 VSUBS 0.006334f
C1159 B.n421 VSUBS 0.006334f
C1160 B.n422 VSUBS 0.006334f
C1161 B.n423 VSUBS 0.006334f
C1162 B.n424 VSUBS 0.006334f
C1163 B.n425 VSUBS 0.006334f
C1164 B.n426 VSUBS 0.006334f
C1165 B.n427 VSUBS 0.006334f
C1166 B.n428 VSUBS 0.006334f
C1167 B.n429 VSUBS 0.006334f
C1168 B.n430 VSUBS 0.006334f
C1169 B.n431 VSUBS 0.006334f
C1170 B.n432 VSUBS 0.006334f
C1171 B.n433 VSUBS 0.006334f
C1172 B.n434 VSUBS 0.006334f
C1173 B.n435 VSUBS 0.006334f
C1174 B.n436 VSUBS 0.006334f
C1175 B.n437 VSUBS 0.006334f
C1176 B.n438 VSUBS 0.006334f
C1177 B.n439 VSUBS 0.006334f
C1178 B.n440 VSUBS 0.006334f
C1179 B.n441 VSUBS 0.006334f
C1180 B.n442 VSUBS 0.006334f
C1181 B.n443 VSUBS 0.006334f
C1182 B.n444 VSUBS 0.006334f
C1183 B.n445 VSUBS 0.006334f
C1184 B.n446 VSUBS 0.006334f
C1185 B.n447 VSUBS 0.006334f
C1186 B.n448 VSUBS 0.006334f
C1187 B.n449 VSUBS 0.006334f
C1188 B.n450 VSUBS 0.006334f
C1189 B.n451 VSUBS 0.006334f
C1190 B.n452 VSUBS 0.006334f
C1191 B.n453 VSUBS 0.006334f
C1192 B.n454 VSUBS 0.006334f
C1193 B.n455 VSUBS 0.006334f
C1194 B.n456 VSUBS 0.006334f
C1195 B.n457 VSUBS 0.006334f
C1196 B.n458 VSUBS 0.006334f
C1197 B.n459 VSUBS 0.006334f
C1198 B.n460 VSUBS 0.006334f
C1199 B.n461 VSUBS 0.006334f
C1200 B.n462 VSUBS 0.006334f
C1201 B.n463 VSUBS 0.006334f
C1202 B.n464 VSUBS 0.006334f
C1203 B.n465 VSUBS 0.006334f
C1204 B.n466 VSUBS 0.006334f
C1205 B.n467 VSUBS 0.006334f
C1206 B.n468 VSUBS 0.006334f
C1207 B.n469 VSUBS 0.006334f
C1208 B.n470 VSUBS 0.006334f
C1209 B.n471 VSUBS 0.006334f
C1210 B.n472 VSUBS 0.006334f
C1211 B.n473 VSUBS 0.006334f
C1212 B.n474 VSUBS 0.006334f
C1213 B.n475 VSUBS 0.006334f
C1214 B.n476 VSUBS 0.006334f
C1215 B.n477 VSUBS 0.006334f
C1216 B.n478 VSUBS 0.006334f
C1217 B.n479 VSUBS 0.006334f
C1218 B.n480 VSUBS 0.006334f
C1219 B.n481 VSUBS 0.006334f
C1220 B.n482 VSUBS 0.006334f
C1221 B.n483 VSUBS 0.006334f
C1222 B.n484 VSUBS 0.006334f
C1223 B.n485 VSUBS 0.006334f
C1224 B.n486 VSUBS 0.006334f
C1225 B.n487 VSUBS 0.006334f
C1226 B.n488 VSUBS 0.006334f
C1227 B.n489 VSUBS 0.006334f
C1228 B.n490 VSUBS 0.006334f
C1229 B.n491 VSUBS 0.006334f
C1230 B.n492 VSUBS 0.006334f
C1231 B.n493 VSUBS 0.005962f
C1232 B.n494 VSUBS 0.006334f
C1233 B.n495 VSUBS 0.006334f
C1234 B.n496 VSUBS 0.00354f
C1235 B.n497 VSUBS 0.006334f
C1236 B.n498 VSUBS 0.006334f
C1237 B.n499 VSUBS 0.006334f
C1238 B.n500 VSUBS 0.006334f
C1239 B.n501 VSUBS 0.006334f
C1240 B.n502 VSUBS 0.006334f
C1241 B.n503 VSUBS 0.006334f
C1242 B.n504 VSUBS 0.006334f
C1243 B.n505 VSUBS 0.006334f
C1244 B.n506 VSUBS 0.006334f
C1245 B.n507 VSUBS 0.006334f
C1246 B.n508 VSUBS 0.006334f
C1247 B.n509 VSUBS 0.00354f
C1248 B.n510 VSUBS 0.014676f
C1249 B.n511 VSUBS 0.005962f
C1250 B.n512 VSUBS 0.006334f
C1251 B.n513 VSUBS 0.006334f
C1252 B.n514 VSUBS 0.006334f
C1253 B.n515 VSUBS 0.006334f
C1254 B.n516 VSUBS 0.006334f
C1255 B.n517 VSUBS 0.006334f
C1256 B.n518 VSUBS 0.006334f
C1257 B.n519 VSUBS 0.006334f
C1258 B.n520 VSUBS 0.006334f
C1259 B.n521 VSUBS 0.006334f
C1260 B.n522 VSUBS 0.006334f
C1261 B.n523 VSUBS 0.006334f
C1262 B.n524 VSUBS 0.006334f
C1263 B.n525 VSUBS 0.006334f
C1264 B.n526 VSUBS 0.006334f
C1265 B.n527 VSUBS 0.006334f
C1266 B.n528 VSUBS 0.006334f
C1267 B.n529 VSUBS 0.006334f
C1268 B.n530 VSUBS 0.006334f
C1269 B.n531 VSUBS 0.006334f
C1270 B.n532 VSUBS 0.006334f
C1271 B.n533 VSUBS 0.006334f
C1272 B.n534 VSUBS 0.006334f
C1273 B.n535 VSUBS 0.006334f
C1274 B.n536 VSUBS 0.006334f
C1275 B.n537 VSUBS 0.006334f
C1276 B.n538 VSUBS 0.006334f
C1277 B.n539 VSUBS 0.006334f
C1278 B.n540 VSUBS 0.006334f
C1279 B.n541 VSUBS 0.006334f
C1280 B.n542 VSUBS 0.006334f
C1281 B.n543 VSUBS 0.006334f
C1282 B.n544 VSUBS 0.006334f
C1283 B.n545 VSUBS 0.006334f
C1284 B.n546 VSUBS 0.006334f
C1285 B.n547 VSUBS 0.006334f
C1286 B.n548 VSUBS 0.006334f
C1287 B.n549 VSUBS 0.006334f
C1288 B.n550 VSUBS 0.006334f
C1289 B.n551 VSUBS 0.006334f
C1290 B.n552 VSUBS 0.006334f
C1291 B.n553 VSUBS 0.006334f
C1292 B.n554 VSUBS 0.006334f
C1293 B.n555 VSUBS 0.006334f
C1294 B.n556 VSUBS 0.006334f
C1295 B.n557 VSUBS 0.006334f
C1296 B.n558 VSUBS 0.006334f
C1297 B.n559 VSUBS 0.006334f
C1298 B.n560 VSUBS 0.006334f
C1299 B.n561 VSUBS 0.006334f
C1300 B.n562 VSUBS 0.006334f
C1301 B.n563 VSUBS 0.006334f
C1302 B.n564 VSUBS 0.006334f
C1303 B.n565 VSUBS 0.006334f
C1304 B.n566 VSUBS 0.006334f
C1305 B.n567 VSUBS 0.006334f
C1306 B.n568 VSUBS 0.006334f
C1307 B.n569 VSUBS 0.006334f
C1308 B.n570 VSUBS 0.006334f
C1309 B.n571 VSUBS 0.006334f
C1310 B.n572 VSUBS 0.006334f
C1311 B.n573 VSUBS 0.006334f
C1312 B.n574 VSUBS 0.006334f
C1313 B.n575 VSUBS 0.006334f
C1314 B.n576 VSUBS 0.006334f
C1315 B.n577 VSUBS 0.006334f
C1316 B.n578 VSUBS 0.006334f
C1317 B.n579 VSUBS 0.006334f
C1318 B.n580 VSUBS 0.006334f
C1319 B.n581 VSUBS 0.006334f
C1320 B.n582 VSUBS 0.006334f
C1321 B.n583 VSUBS 0.006334f
C1322 B.n584 VSUBS 0.006334f
C1323 B.n585 VSUBS 0.006334f
C1324 B.n586 VSUBS 0.006334f
C1325 B.n587 VSUBS 0.006334f
C1326 B.n588 VSUBS 0.015759f
C1327 B.n589 VSUBS 0.014982f
C1328 B.n590 VSUBS 0.014982f
C1329 B.n591 VSUBS 0.006334f
C1330 B.n592 VSUBS 0.006334f
C1331 B.n593 VSUBS 0.006334f
C1332 B.n594 VSUBS 0.006334f
C1333 B.n595 VSUBS 0.006334f
C1334 B.n596 VSUBS 0.006334f
C1335 B.n597 VSUBS 0.006334f
C1336 B.n598 VSUBS 0.006334f
C1337 B.n599 VSUBS 0.006334f
C1338 B.n600 VSUBS 0.006334f
C1339 B.n601 VSUBS 0.006334f
C1340 B.n602 VSUBS 0.006334f
C1341 B.n603 VSUBS 0.006334f
C1342 B.n604 VSUBS 0.006334f
C1343 B.n605 VSUBS 0.006334f
C1344 B.n606 VSUBS 0.006334f
C1345 B.n607 VSUBS 0.006334f
C1346 B.n608 VSUBS 0.006334f
C1347 B.n609 VSUBS 0.006334f
C1348 B.n610 VSUBS 0.006334f
C1349 B.n611 VSUBS 0.006334f
C1350 B.n612 VSUBS 0.006334f
C1351 B.n613 VSUBS 0.006334f
C1352 B.n614 VSUBS 0.006334f
C1353 B.n615 VSUBS 0.008266f
C1354 B.n616 VSUBS 0.008806f
C1355 B.n617 VSUBS 0.017511f
.ends

