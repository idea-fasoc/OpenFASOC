* NGSPICE file created from diff_pair_sample_1170.ext - technology: sky130A

.subckt diff_pair_sample_1170 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t6 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0.84315 ps=5.44 w=5.11 l=2.81
X1 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.84315 pd=5.44 as=1.9929 ps=11 w=5.11 l=2.81
X2 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0.84315 ps=5.44 w=5.11 l=2.81
X3 VTAIL.t1 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0.84315 ps=5.44 w=5.11 l=2.81
X4 VDD2.t3 VN.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.84315 pd=5.44 as=1.9929 ps=11 w=5.11 l=2.81
X5 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0 ps=0 w=5.11 l=2.81
X6 VDD2.t0 VN.t2 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.84315 pd=5.44 as=1.9929 ps=11 w=5.11 l=2.81
X7 VTAIL.t3 VN.t3 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0.84315 ps=5.44 w=5.11 l=2.81
X8 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0 ps=0 w=5.11 l=2.81
X9 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0 ps=0 w=5.11 l=2.81
X10 VDD1.t0 VP.t3 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.84315 pd=5.44 as=1.9929 ps=11 w=5.11 l=2.81
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.9929 pd=11 as=0 ps=0 w=5.11 l=2.81
R0 VN.n0 VN.t0 78.8747
R1 VN.n1 VN.t2 78.8747
R2 VN.n0 VN.t1 77.9842
R3 VN.n1 VN.t3 77.9842
R4 VN VN.n1 45.4899
R5 VN VN.n0 3.49365
R6 VDD2.n2 VDD2.n0 107.579
R7 VDD2.n2 VDD2.n1 71.3378
R8 VDD2.n1 VDD2.t1 3.87526
R9 VDD2.n1 VDD2.t0 3.87526
R10 VDD2.n0 VDD2.t2 3.87526
R11 VDD2.n0 VDD2.t3 3.87526
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n206 VTAIL.n205 289.615
R14 VTAIL.n24 VTAIL.n23 289.615
R15 VTAIL.n50 VTAIL.n49 289.615
R16 VTAIL.n76 VTAIL.n75 289.615
R17 VTAIL.n180 VTAIL.n179 289.615
R18 VTAIL.n154 VTAIL.n153 289.615
R19 VTAIL.n128 VTAIL.n127 289.615
R20 VTAIL.n102 VTAIL.n101 289.615
R21 VTAIL.n191 VTAIL.n190 185
R22 VTAIL.n188 VTAIL.n187 185
R23 VTAIL.n197 VTAIL.n196 185
R24 VTAIL.n199 VTAIL.n198 185
R25 VTAIL.n184 VTAIL.n183 185
R26 VTAIL.n205 VTAIL.n204 185
R27 VTAIL.n9 VTAIL.n8 185
R28 VTAIL.n6 VTAIL.n5 185
R29 VTAIL.n15 VTAIL.n14 185
R30 VTAIL.n17 VTAIL.n16 185
R31 VTAIL.n2 VTAIL.n1 185
R32 VTAIL.n23 VTAIL.n22 185
R33 VTAIL.n35 VTAIL.n34 185
R34 VTAIL.n32 VTAIL.n31 185
R35 VTAIL.n41 VTAIL.n40 185
R36 VTAIL.n43 VTAIL.n42 185
R37 VTAIL.n28 VTAIL.n27 185
R38 VTAIL.n49 VTAIL.n48 185
R39 VTAIL.n61 VTAIL.n60 185
R40 VTAIL.n58 VTAIL.n57 185
R41 VTAIL.n67 VTAIL.n66 185
R42 VTAIL.n69 VTAIL.n68 185
R43 VTAIL.n54 VTAIL.n53 185
R44 VTAIL.n75 VTAIL.n74 185
R45 VTAIL.n179 VTAIL.n178 185
R46 VTAIL.n158 VTAIL.n157 185
R47 VTAIL.n173 VTAIL.n172 185
R48 VTAIL.n171 VTAIL.n170 185
R49 VTAIL.n162 VTAIL.n161 185
R50 VTAIL.n165 VTAIL.n164 185
R51 VTAIL.n153 VTAIL.n152 185
R52 VTAIL.n132 VTAIL.n131 185
R53 VTAIL.n147 VTAIL.n146 185
R54 VTAIL.n145 VTAIL.n144 185
R55 VTAIL.n136 VTAIL.n135 185
R56 VTAIL.n139 VTAIL.n138 185
R57 VTAIL.n127 VTAIL.n126 185
R58 VTAIL.n106 VTAIL.n105 185
R59 VTAIL.n121 VTAIL.n120 185
R60 VTAIL.n119 VTAIL.n118 185
R61 VTAIL.n110 VTAIL.n109 185
R62 VTAIL.n113 VTAIL.n112 185
R63 VTAIL.n101 VTAIL.n100 185
R64 VTAIL.n80 VTAIL.n79 185
R65 VTAIL.n95 VTAIL.n94 185
R66 VTAIL.n93 VTAIL.n92 185
R67 VTAIL.n84 VTAIL.n83 185
R68 VTAIL.n87 VTAIL.n86 185
R69 VTAIL.t5 VTAIL.n189 149.54
R70 VTAIL.t6 VTAIL.n7 149.54
R71 VTAIL.t7 VTAIL.n33 149.54
R72 VTAIL.t1 VTAIL.n59 149.54
R73 VTAIL.t0 VTAIL.n137 149.54
R74 VTAIL.t4 VTAIL.n111 149.54
R75 VTAIL.t3 VTAIL.n85 149.54
R76 VTAIL.t2 VTAIL.n163 149.54
R77 VTAIL.n190 VTAIL.n187 104.615
R78 VTAIL.n197 VTAIL.n187 104.615
R79 VTAIL.n198 VTAIL.n197 104.615
R80 VTAIL.n198 VTAIL.n183 104.615
R81 VTAIL.n205 VTAIL.n183 104.615
R82 VTAIL.n8 VTAIL.n5 104.615
R83 VTAIL.n15 VTAIL.n5 104.615
R84 VTAIL.n16 VTAIL.n15 104.615
R85 VTAIL.n16 VTAIL.n1 104.615
R86 VTAIL.n23 VTAIL.n1 104.615
R87 VTAIL.n34 VTAIL.n31 104.615
R88 VTAIL.n41 VTAIL.n31 104.615
R89 VTAIL.n42 VTAIL.n41 104.615
R90 VTAIL.n42 VTAIL.n27 104.615
R91 VTAIL.n49 VTAIL.n27 104.615
R92 VTAIL.n60 VTAIL.n57 104.615
R93 VTAIL.n67 VTAIL.n57 104.615
R94 VTAIL.n68 VTAIL.n67 104.615
R95 VTAIL.n68 VTAIL.n53 104.615
R96 VTAIL.n75 VTAIL.n53 104.615
R97 VTAIL.n179 VTAIL.n157 104.615
R98 VTAIL.n172 VTAIL.n157 104.615
R99 VTAIL.n172 VTAIL.n171 104.615
R100 VTAIL.n171 VTAIL.n161 104.615
R101 VTAIL.n164 VTAIL.n161 104.615
R102 VTAIL.n153 VTAIL.n131 104.615
R103 VTAIL.n146 VTAIL.n131 104.615
R104 VTAIL.n146 VTAIL.n145 104.615
R105 VTAIL.n145 VTAIL.n135 104.615
R106 VTAIL.n138 VTAIL.n135 104.615
R107 VTAIL.n127 VTAIL.n105 104.615
R108 VTAIL.n120 VTAIL.n105 104.615
R109 VTAIL.n120 VTAIL.n119 104.615
R110 VTAIL.n119 VTAIL.n109 104.615
R111 VTAIL.n112 VTAIL.n109 104.615
R112 VTAIL.n101 VTAIL.n79 104.615
R113 VTAIL.n94 VTAIL.n79 104.615
R114 VTAIL.n94 VTAIL.n93 104.615
R115 VTAIL.n93 VTAIL.n83 104.615
R116 VTAIL.n86 VTAIL.n83 104.615
R117 VTAIL.n190 VTAIL.t5 52.3082
R118 VTAIL.n8 VTAIL.t6 52.3082
R119 VTAIL.n34 VTAIL.t7 52.3082
R120 VTAIL.n60 VTAIL.t1 52.3082
R121 VTAIL.n164 VTAIL.t2 52.3082
R122 VTAIL.n138 VTAIL.t0 52.3082
R123 VTAIL.n112 VTAIL.t4 52.3082
R124 VTAIL.n86 VTAIL.t3 52.3082
R125 VTAIL.n207 VTAIL.n206 33.9308
R126 VTAIL.n25 VTAIL.n24 33.9308
R127 VTAIL.n51 VTAIL.n50 33.9308
R128 VTAIL.n77 VTAIL.n76 33.9308
R129 VTAIL.n181 VTAIL.n180 33.9308
R130 VTAIL.n155 VTAIL.n154 33.9308
R131 VTAIL.n129 VTAIL.n128 33.9308
R132 VTAIL.n103 VTAIL.n102 33.9308
R133 VTAIL.n207 VTAIL.n181 19.4789
R134 VTAIL.n103 VTAIL.n77 19.4789
R135 VTAIL.n204 VTAIL.n182 11.249
R136 VTAIL.n22 VTAIL.n0 11.249
R137 VTAIL.n48 VTAIL.n26 11.249
R138 VTAIL.n74 VTAIL.n52 11.249
R139 VTAIL.n178 VTAIL.n156 11.249
R140 VTAIL.n152 VTAIL.n130 11.249
R141 VTAIL.n126 VTAIL.n104 11.249
R142 VTAIL.n100 VTAIL.n78 11.249
R143 VTAIL.n203 VTAIL.n184 10.4732
R144 VTAIL.n21 VTAIL.n2 10.4732
R145 VTAIL.n47 VTAIL.n28 10.4732
R146 VTAIL.n73 VTAIL.n54 10.4732
R147 VTAIL.n177 VTAIL.n158 10.4732
R148 VTAIL.n151 VTAIL.n132 10.4732
R149 VTAIL.n125 VTAIL.n106 10.4732
R150 VTAIL.n99 VTAIL.n80 10.4732
R151 VTAIL.n191 VTAIL.n189 10.2739
R152 VTAIL.n9 VTAIL.n7 10.2739
R153 VTAIL.n35 VTAIL.n33 10.2739
R154 VTAIL.n61 VTAIL.n59 10.2739
R155 VTAIL.n165 VTAIL.n163 10.2739
R156 VTAIL.n139 VTAIL.n137 10.2739
R157 VTAIL.n113 VTAIL.n111 10.2739
R158 VTAIL.n87 VTAIL.n85 10.2739
R159 VTAIL.n200 VTAIL.n199 9.69747
R160 VTAIL.n18 VTAIL.n17 9.69747
R161 VTAIL.n44 VTAIL.n43 9.69747
R162 VTAIL.n70 VTAIL.n69 9.69747
R163 VTAIL.n174 VTAIL.n173 9.69747
R164 VTAIL.n148 VTAIL.n147 9.69747
R165 VTAIL.n122 VTAIL.n121 9.69747
R166 VTAIL.n96 VTAIL.n95 9.69747
R167 VTAIL.n202 VTAIL.n182 9.45567
R168 VTAIL.n20 VTAIL.n0 9.45567
R169 VTAIL.n46 VTAIL.n26 9.45567
R170 VTAIL.n72 VTAIL.n52 9.45567
R171 VTAIL.n176 VTAIL.n156 9.45567
R172 VTAIL.n150 VTAIL.n130 9.45567
R173 VTAIL.n124 VTAIL.n104 9.45567
R174 VTAIL.n98 VTAIL.n78 9.45567
R175 VTAIL.n193 VTAIL.n192 9.3005
R176 VTAIL.n195 VTAIL.n194 9.3005
R177 VTAIL.n186 VTAIL.n185 9.3005
R178 VTAIL.n201 VTAIL.n200 9.3005
R179 VTAIL.n203 VTAIL.n202 9.3005
R180 VTAIL.n11 VTAIL.n10 9.3005
R181 VTAIL.n13 VTAIL.n12 9.3005
R182 VTAIL.n4 VTAIL.n3 9.3005
R183 VTAIL.n19 VTAIL.n18 9.3005
R184 VTAIL.n21 VTAIL.n20 9.3005
R185 VTAIL.n37 VTAIL.n36 9.3005
R186 VTAIL.n39 VTAIL.n38 9.3005
R187 VTAIL.n30 VTAIL.n29 9.3005
R188 VTAIL.n45 VTAIL.n44 9.3005
R189 VTAIL.n47 VTAIL.n46 9.3005
R190 VTAIL.n63 VTAIL.n62 9.3005
R191 VTAIL.n65 VTAIL.n64 9.3005
R192 VTAIL.n56 VTAIL.n55 9.3005
R193 VTAIL.n71 VTAIL.n70 9.3005
R194 VTAIL.n73 VTAIL.n72 9.3005
R195 VTAIL.n177 VTAIL.n176 9.3005
R196 VTAIL.n175 VTAIL.n174 9.3005
R197 VTAIL.n160 VTAIL.n159 9.3005
R198 VTAIL.n169 VTAIL.n168 9.3005
R199 VTAIL.n167 VTAIL.n166 9.3005
R200 VTAIL.n143 VTAIL.n142 9.3005
R201 VTAIL.n134 VTAIL.n133 9.3005
R202 VTAIL.n149 VTAIL.n148 9.3005
R203 VTAIL.n151 VTAIL.n150 9.3005
R204 VTAIL.n141 VTAIL.n140 9.3005
R205 VTAIL.n117 VTAIL.n116 9.3005
R206 VTAIL.n108 VTAIL.n107 9.3005
R207 VTAIL.n123 VTAIL.n122 9.3005
R208 VTAIL.n125 VTAIL.n124 9.3005
R209 VTAIL.n115 VTAIL.n114 9.3005
R210 VTAIL.n91 VTAIL.n90 9.3005
R211 VTAIL.n82 VTAIL.n81 9.3005
R212 VTAIL.n97 VTAIL.n96 9.3005
R213 VTAIL.n99 VTAIL.n98 9.3005
R214 VTAIL.n89 VTAIL.n88 9.3005
R215 VTAIL.n196 VTAIL.n186 8.92171
R216 VTAIL.n14 VTAIL.n4 8.92171
R217 VTAIL.n40 VTAIL.n30 8.92171
R218 VTAIL.n66 VTAIL.n56 8.92171
R219 VTAIL.n170 VTAIL.n160 8.92171
R220 VTAIL.n144 VTAIL.n134 8.92171
R221 VTAIL.n118 VTAIL.n108 8.92171
R222 VTAIL.n92 VTAIL.n82 8.92171
R223 VTAIL.n195 VTAIL.n188 8.14595
R224 VTAIL.n13 VTAIL.n6 8.14595
R225 VTAIL.n39 VTAIL.n32 8.14595
R226 VTAIL.n65 VTAIL.n58 8.14595
R227 VTAIL.n169 VTAIL.n162 8.14595
R228 VTAIL.n143 VTAIL.n136 8.14595
R229 VTAIL.n117 VTAIL.n110 8.14595
R230 VTAIL.n91 VTAIL.n84 8.14595
R231 VTAIL.n192 VTAIL.n191 7.3702
R232 VTAIL.n10 VTAIL.n9 7.3702
R233 VTAIL.n36 VTAIL.n35 7.3702
R234 VTAIL.n62 VTAIL.n61 7.3702
R235 VTAIL.n166 VTAIL.n165 7.3702
R236 VTAIL.n140 VTAIL.n139 7.3702
R237 VTAIL.n114 VTAIL.n113 7.3702
R238 VTAIL.n88 VTAIL.n87 7.3702
R239 VTAIL.n192 VTAIL.n188 5.81868
R240 VTAIL.n10 VTAIL.n6 5.81868
R241 VTAIL.n36 VTAIL.n32 5.81868
R242 VTAIL.n62 VTAIL.n58 5.81868
R243 VTAIL.n166 VTAIL.n162 5.81868
R244 VTAIL.n140 VTAIL.n136 5.81868
R245 VTAIL.n114 VTAIL.n110 5.81868
R246 VTAIL.n88 VTAIL.n84 5.81868
R247 VTAIL.n196 VTAIL.n195 5.04292
R248 VTAIL.n14 VTAIL.n13 5.04292
R249 VTAIL.n40 VTAIL.n39 5.04292
R250 VTAIL.n66 VTAIL.n65 5.04292
R251 VTAIL.n170 VTAIL.n169 5.04292
R252 VTAIL.n144 VTAIL.n143 5.04292
R253 VTAIL.n118 VTAIL.n117 5.04292
R254 VTAIL.n92 VTAIL.n91 5.04292
R255 VTAIL.n199 VTAIL.n186 4.26717
R256 VTAIL.n17 VTAIL.n4 4.26717
R257 VTAIL.n43 VTAIL.n30 4.26717
R258 VTAIL.n69 VTAIL.n56 4.26717
R259 VTAIL.n173 VTAIL.n160 4.26717
R260 VTAIL.n147 VTAIL.n134 4.26717
R261 VTAIL.n121 VTAIL.n108 4.26717
R262 VTAIL.n95 VTAIL.n82 4.26717
R263 VTAIL.n200 VTAIL.n184 3.49141
R264 VTAIL.n18 VTAIL.n2 3.49141
R265 VTAIL.n44 VTAIL.n28 3.49141
R266 VTAIL.n70 VTAIL.n54 3.49141
R267 VTAIL.n174 VTAIL.n158 3.49141
R268 VTAIL.n148 VTAIL.n132 3.49141
R269 VTAIL.n122 VTAIL.n106 3.49141
R270 VTAIL.n96 VTAIL.n80 3.49141
R271 VTAIL.n193 VTAIL.n189 2.84386
R272 VTAIL.n11 VTAIL.n7 2.84386
R273 VTAIL.n37 VTAIL.n33 2.84386
R274 VTAIL.n63 VTAIL.n59 2.84386
R275 VTAIL.n141 VTAIL.n137 2.84386
R276 VTAIL.n115 VTAIL.n111 2.84386
R277 VTAIL.n89 VTAIL.n85 2.84386
R278 VTAIL.n167 VTAIL.n163 2.84386
R279 VTAIL.n204 VTAIL.n203 2.71565
R280 VTAIL.n22 VTAIL.n21 2.71565
R281 VTAIL.n48 VTAIL.n47 2.71565
R282 VTAIL.n74 VTAIL.n73 2.71565
R283 VTAIL.n178 VTAIL.n177 2.71565
R284 VTAIL.n152 VTAIL.n151 2.71565
R285 VTAIL.n126 VTAIL.n125 2.71565
R286 VTAIL.n100 VTAIL.n99 2.71565
R287 VTAIL.n129 VTAIL.n103 2.7074
R288 VTAIL.n181 VTAIL.n155 2.7074
R289 VTAIL.n77 VTAIL.n51 2.7074
R290 VTAIL.n206 VTAIL.n182 1.93989
R291 VTAIL.n24 VTAIL.n0 1.93989
R292 VTAIL.n50 VTAIL.n26 1.93989
R293 VTAIL.n76 VTAIL.n52 1.93989
R294 VTAIL.n180 VTAIL.n156 1.93989
R295 VTAIL.n154 VTAIL.n130 1.93989
R296 VTAIL.n128 VTAIL.n104 1.93989
R297 VTAIL.n102 VTAIL.n78 1.93989
R298 VTAIL VTAIL.n25 1.41214
R299 VTAIL VTAIL.n207 1.29576
R300 VTAIL.n155 VTAIL.n129 0.470328
R301 VTAIL.n51 VTAIL.n25 0.470328
R302 VTAIL.n194 VTAIL.n193 0.155672
R303 VTAIL.n194 VTAIL.n185 0.155672
R304 VTAIL.n201 VTAIL.n185 0.155672
R305 VTAIL.n202 VTAIL.n201 0.155672
R306 VTAIL.n12 VTAIL.n11 0.155672
R307 VTAIL.n12 VTAIL.n3 0.155672
R308 VTAIL.n19 VTAIL.n3 0.155672
R309 VTAIL.n20 VTAIL.n19 0.155672
R310 VTAIL.n38 VTAIL.n37 0.155672
R311 VTAIL.n38 VTAIL.n29 0.155672
R312 VTAIL.n45 VTAIL.n29 0.155672
R313 VTAIL.n46 VTAIL.n45 0.155672
R314 VTAIL.n64 VTAIL.n63 0.155672
R315 VTAIL.n64 VTAIL.n55 0.155672
R316 VTAIL.n71 VTAIL.n55 0.155672
R317 VTAIL.n72 VTAIL.n71 0.155672
R318 VTAIL.n176 VTAIL.n175 0.155672
R319 VTAIL.n175 VTAIL.n159 0.155672
R320 VTAIL.n168 VTAIL.n159 0.155672
R321 VTAIL.n168 VTAIL.n167 0.155672
R322 VTAIL.n150 VTAIL.n149 0.155672
R323 VTAIL.n149 VTAIL.n133 0.155672
R324 VTAIL.n142 VTAIL.n133 0.155672
R325 VTAIL.n142 VTAIL.n141 0.155672
R326 VTAIL.n124 VTAIL.n123 0.155672
R327 VTAIL.n123 VTAIL.n107 0.155672
R328 VTAIL.n116 VTAIL.n107 0.155672
R329 VTAIL.n116 VTAIL.n115 0.155672
R330 VTAIL.n98 VTAIL.n97 0.155672
R331 VTAIL.n97 VTAIL.n81 0.155672
R332 VTAIL.n90 VTAIL.n81 0.155672
R333 VTAIL.n90 VTAIL.n89 0.155672
R334 B.n560 B.n559 585
R335 B.n199 B.n94 585
R336 B.n198 B.n197 585
R337 B.n196 B.n195 585
R338 B.n194 B.n193 585
R339 B.n192 B.n191 585
R340 B.n190 B.n189 585
R341 B.n188 B.n187 585
R342 B.n186 B.n185 585
R343 B.n184 B.n183 585
R344 B.n182 B.n181 585
R345 B.n180 B.n179 585
R346 B.n178 B.n177 585
R347 B.n176 B.n175 585
R348 B.n174 B.n173 585
R349 B.n172 B.n171 585
R350 B.n170 B.n169 585
R351 B.n168 B.n167 585
R352 B.n166 B.n165 585
R353 B.n164 B.n163 585
R354 B.n162 B.n161 585
R355 B.n159 B.n158 585
R356 B.n157 B.n156 585
R357 B.n155 B.n154 585
R358 B.n153 B.n152 585
R359 B.n151 B.n150 585
R360 B.n149 B.n148 585
R361 B.n147 B.n146 585
R362 B.n145 B.n144 585
R363 B.n143 B.n142 585
R364 B.n141 B.n140 585
R365 B.n138 B.n137 585
R366 B.n136 B.n135 585
R367 B.n134 B.n133 585
R368 B.n132 B.n131 585
R369 B.n130 B.n129 585
R370 B.n128 B.n127 585
R371 B.n126 B.n125 585
R372 B.n124 B.n123 585
R373 B.n122 B.n121 585
R374 B.n120 B.n119 585
R375 B.n118 B.n117 585
R376 B.n116 B.n115 585
R377 B.n114 B.n113 585
R378 B.n112 B.n111 585
R379 B.n110 B.n109 585
R380 B.n108 B.n107 585
R381 B.n106 B.n105 585
R382 B.n104 B.n103 585
R383 B.n102 B.n101 585
R384 B.n100 B.n99 585
R385 B.n67 B.n66 585
R386 B.n558 B.n68 585
R387 B.n563 B.n68 585
R388 B.n557 B.n556 585
R389 B.n556 B.n64 585
R390 B.n555 B.n63 585
R391 B.n569 B.n63 585
R392 B.n554 B.n62 585
R393 B.n570 B.n62 585
R394 B.n553 B.n61 585
R395 B.n571 B.n61 585
R396 B.n552 B.n551 585
R397 B.n551 B.n57 585
R398 B.n550 B.n56 585
R399 B.n577 B.n56 585
R400 B.n549 B.n55 585
R401 B.n578 B.n55 585
R402 B.n548 B.n54 585
R403 B.n579 B.n54 585
R404 B.n547 B.n546 585
R405 B.n546 B.n50 585
R406 B.n545 B.n49 585
R407 B.n585 B.n49 585
R408 B.n544 B.n48 585
R409 B.n586 B.n48 585
R410 B.n543 B.n47 585
R411 B.n587 B.n47 585
R412 B.n542 B.n541 585
R413 B.n541 B.n43 585
R414 B.n540 B.n42 585
R415 B.n593 B.n42 585
R416 B.n539 B.n41 585
R417 B.n594 B.n41 585
R418 B.n538 B.n40 585
R419 B.n595 B.n40 585
R420 B.n537 B.n536 585
R421 B.n536 B.n36 585
R422 B.n535 B.n35 585
R423 B.n601 B.n35 585
R424 B.n534 B.n34 585
R425 B.n602 B.n34 585
R426 B.n533 B.n33 585
R427 B.n603 B.n33 585
R428 B.n532 B.n531 585
R429 B.n531 B.n29 585
R430 B.n530 B.n28 585
R431 B.n609 B.n28 585
R432 B.n529 B.n27 585
R433 B.n610 B.n27 585
R434 B.n528 B.n26 585
R435 B.n611 B.n26 585
R436 B.n527 B.n526 585
R437 B.n526 B.n22 585
R438 B.n525 B.n21 585
R439 B.n617 B.n21 585
R440 B.n524 B.n20 585
R441 B.n618 B.n20 585
R442 B.n523 B.n19 585
R443 B.n619 B.n19 585
R444 B.n522 B.n521 585
R445 B.n521 B.n18 585
R446 B.n520 B.n14 585
R447 B.n625 B.n14 585
R448 B.n519 B.n13 585
R449 B.n626 B.n13 585
R450 B.n518 B.n12 585
R451 B.n627 B.n12 585
R452 B.n517 B.n516 585
R453 B.n516 B.n8 585
R454 B.n515 B.n7 585
R455 B.n633 B.n7 585
R456 B.n514 B.n6 585
R457 B.n634 B.n6 585
R458 B.n513 B.n5 585
R459 B.n635 B.n5 585
R460 B.n512 B.n511 585
R461 B.n511 B.n4 585
R462 B.n510 B.n200 585
R463 B.n510 B.n509 585
R464 B.n500 B.n201 585
R465 B.n202 B.n201 585
R466 B.n502 B.n501 585
R467 B.n503 B.n502 585
R468 B.n499 B.n207 585
R469 B.n207 B.n206 585
R470 B.n498 B.n497 585
R471 B.n497 B.n496 585
R472 B.n209 B.n208 585
R473 B.n489 B.n209 585
R474 B.n488 B.n487 585
R475 B.n490 B.n488 585
R476 B.n486 B.n214 585
R477 B.n214 B.n213 585
R478 B.n485 B.n484 585
R479 B.n484 B.n483 585
R480 B.n216 B.n215 585
R481 B.n217 B.n216 585
R482 B.n476 B.n475 585
R483 B.n477 B.n476 585
R484 B.n474 B.n222 585
R485 B.n222 B.n221 585
R486 B.n473 B.n472 585
R487 B.n472 B.n471 585
R488 B.n224 B.n223 585
R489 B.n225 B.n224 585
R490 B.n464 B.n463 585
R491 B.n465 B.n464 585
R492 B.n462 B.n230 585
R493 B.n230 B.n229 585
R494 B.n461 B.n460 585
R495 B.n460 B.n459 585
R496 B.n232 B.n231 585
R497 B.n233 B.n232 585
R498 B.n452 B.n451 585
R499 B.n453 B.n452 585
R500 B.n450 B.n238 585
R501 B.n238 B.n237 585
R502 B.n449 B.n448 585
R503 B.n448 B.n447 585
R504 B.n240 B.n239 585
R505 B.n241 B.n240 585
R506 B.n440 B.n439 585
R507 B.n441 B.n440 585
R508 B.n438 B.n246 585
R509 B.n246 B.n245 585
R510 B.n437 B.n436 585
R511 B.n436 B.n435 585
R512 B.n248 B.n247 585
R513 B.n249 B.n248 585
R514 B.n428 B.n427 585
R515 B.n429 B.n428 585
R516 B.n426 B.n254 585
R517 B.n254 B.n253 585
R518 B.n425 B.n424 585
R519 B.n424 B.n423 585
R520 B.n256 B.n255 585
R521 B.n257 B.n256 585
R522 B.n416 B.n415 585
R523 B.n417 B.n416 585
R524 B.n414 B.n262 585
R525 B.n262 B.n261 585
R526 B.n413 B.n412 585
R527 B.n412 B.n411 585
R528 B.n264 B.n263 585
R529 B.n265 B.n264 585
R530 B.n404 B.n403 585
R531 B.n405 B.n404 585
R532 B.n268 B.n267 585
R533 B.n303 B.n302 585
R534 B.n304 B.n300 585
R535 B.n300 B.n269 585
R536 B.n306 B.n305 585
R537 B.n308 B.n299 585
R538 B.n311 B.n310 585
R539 B.n312 B.n298 585
R540 B.n314 B.n313 585
R541 B.n316 B.n297 585
R542 B.n319 B.n318 585
R543 B.n320 B.n296 585
R544 B.n322 B.n321 585
R545 B.n324 B.n295 585
R546 B.n327 B.n326 585
R547 B.n328 B.n294 585
R548 B.n330 B.n329 585
R549 B.n332 B.n293 585
R550 B.n335 B.n334 585
R551 B.n336 B.n292 585
R552 B.n338 B.n337 585
R553 B.n340 B.n291 585
R554 B.n343 B.n342 585
R555 B.n344 B.n287 585
R556 B.n346 B.n345 585
R557 B.n348 B.n286 585
R558 B.n351 B.n350 585
R559 B.n352 B.n285 585
R560 B.n354 B.n353 585
R561 B.n356 B.n284 585
R562 B.n359 B.n358 585
R563 B.n360 B.n281 585
R564 B.n363 B.n362 585
R565 B.n365 B.n280 585
R566 B.n368 B.n367 585
R567 B.n369 B.n279 585
R568 B.n371 B.n370 585
R569 B.n373 B.n278 585
R570 B.n376 B.n375 585
R571 B.n377 B.n277 585
R572 B.n379 B.n378 585
R573 B.n381 B.n276 585
R574 B.n384 B.n383 585
R575 B.n385 B.n275 585
R576 B.n387 B.n386 585
R577 B.n389 B.n274 585
R578 B.n392 B.n391 585
R579 B.n393 B.n273 585
R580 B.n395 B.n394 585
R581 B.n397 B.n272 585
R582 B.n398 B.n271 585
R583 B.n401 B.n400 585
R584 B.n402 B.n270 585
R585 B.n270 B.n269 585
R586 B.n407 B.n406 585
R587 B.n406 B.n405 585
R588 B.n408 B.n266 585
R589 B.n266 B.n265 585
R590 B.n410 B.n409 585
R591 B.n411 B.n410 585
R592 B.n260 B.n259 585
R593 B.n261 B.n260 585
R594 B.n419 B.n418 585
R595 B.n418 B.n417 585
R596 B.n420 B.n258 585
R597 B.n258 B.n257 585
R598 B.n422 B.n421 585
R599 B.n423 B.n422 585
R600 B.n252 B.n251 585
R601 B.n253 B.n252 585
R602 B.n431 B.n430 585
R603 B.n430 B.n429 585
R604 B.n432 B.n250 585
R605 B.n250 B.n249 585
R606 B.n434 B.n433 585
R607 B.n435 B.n434 585
R608 B.n244 B.n243 585
R609 B.n245 B.n244 585
R610 B.n443 B.n442 585
R611 B.n442 B.n441 585
R612 B.n444 B.n242 585
R613 B.n242 B.n241 585
R614 B.n446 B.n445 585
R615 B.n447 B.n446 585
R616 B.n236 B.n235 585
R617 B.n237 B.n236 585
R618 B.n455 B.n454 585
R619 B.n454 B.n453 585
R620 B.n456 B.n234 585
R621 B.n234 B.n233 585
R622 B.n458 B.n457 585
R623 B.n459 B.n458 585
R624 B.n228 B.n227 585
R625 B.n229 B.n228 585
R626 B.n467 B.n466 585
R627 B.n466 B.n465 585
R628 B.n468 B.n226 585
R629 B.n226 B.n225 585
R630 B.n470 B.n469 585
R631 B.n471 B.n470 585
R632 B.n220 B.n219 585
R633 B.n221 B.n220 585
R634 B.n479 B.n478 585
R635 B.n478 B.n477 585
R636 B.n480 B.n218 585
R637 B.n218 B.n217 585
R638 B.n482 B.n481 585
R639 B.n483 B.n482 585
R640 B.n212 B.n211 585
R641 B.n213 B.n212 585
R642 B.n492 B.n491 585
R643 B.n491 B.n490 585
R644 B.n493 B.n210 585
R645 B.n489 B.n210 585
R646 B.n495 B.n494 585
R647 B.n496 B.n495 585
R648 B.n205 B.n204 585
R649 B.n206 B.n205 585
R650 B.n505 B.n504 585
R651 B.n504 B.n503 585
R652 B.n506 B.n203 585
R653 B.n203 B.n202 585
R654 B.n508 B.n507 585
R655 B.n509 B.n508 585
R656 B.n2 B.n0 585
R657 B.n4 B.n2 585
R658 B.n3 B.n1 585
R659 B.n634 B.n3 585
R660 B.n632 B.n631 585
R661 B.n633 B.n632 585
R662 B.n630 B.n9 585
R663 B.n9 B.n8 585
R664 B.n629 B.n628 585
R665 B.n628 B.n627 585
R666 B.n11 B.n10 585
R667 B.n626 B.n11 585
R668 B.n624 B.n623 585
R669 B.n625 B.n624 585
R670 B.n622 B.n15 585
R671 B.n18 B.n15 585
R672 B.n621 B.n620 585
R673 B.n620 B.n619 585
R674 B.n17 B.n16 585
R675 B.n618 B.n17 585
R676 B.n616 B.n615 585
R677 B.n617 B.n616 585
R678 B.n614 B.n23 585
R679 B.n23 B.n22 585
R680 B.n613 B.n612 585
R681 B.n612 B.n611 585
R682 B.n25 B.n24 585
R683 B.n610 B.n25 585
R684 B.n608 B.n607 585
R685 B.n609 B.n608 585
R686 B.n606 B.n30 585
R687 B.n30 B.n29 585
R688 B.n605 B.n604 585
R689 B.n604 B.n603 585
R690 B.n32 B.n31 585
R691 B.n602 B.n32 585
R692 B.n600 B.n599 585
R693 B.n601 B.n600 585
R694 B.n598 B.n37 585
R695 B.n37 B.n36 585
R696 B.n597 B.n596 585
R697 B.n596 B.n595 585
R698 B.n39 B.n38 585
R699 B.n594 B.n39 585
R700 B.n592 B.n591 585
R701 B.n593 B.n592 585
R702 B.n590 B.n44 585
R703 B.n44 B.n43 585
R704 B.n589 B.n588 585
R705 B.n588 B.n587 585
R706 B.n46 B.n45 585
R707 B.n586 B.n46 585
R708 B.n584 B.n583 585
R709 B.n585 B.n584 585
R710 B.n582 B.n51 585
R711 B.n51 B.n50 585
R712 B.n581 B.n580 585
R713 B.n580 B.n579 585
R714 B.n53 B.n52 585
R715 B.n578 B.n53 585
R716 B.n576 B.n575 585
R717 B.n577 B.n576 585
R718 B.n574 B.n58 585
R719 B.n58 B.n57 585
R720 B.n573 B.n572 585
R721 B.n572 B.n571 585
R722 B.n60 B.n59 585
R723 B.n570 B.n60 585
R724 B.n568 B.n567 585
R725 B.n569 B.n568 585
R726 B.n566 B.n65 585
R727 B.n65 B.n64 585
R728 B.n565 B.n564 585
R729 B.n564 B.n563 585
R730 B.n637 B.n636 585
R731 B.n636 B.n635 585
R732 B.n406 B.n268 492.5
R733 B.n564 B.n67 492.5
R734 B.n404 B.n270 492.5
R735 B.n560 B.n68 492.5
R736 B.n562 B.n561 256.663
R737 B.n562 B.n93 256.663
R738 B.n562 B.n92 256.663
R739 B.n562 B.n91 256.663
R740 B.n562 B.n90 256.663
R741 B.n562 B.n89 256.663
R742 B.n562 B.n88 256.663
R743 B.n562 B.n87 256.663
R744 B.n562 B.n86 256.663
R745 B.n562 B.n85 256.663
R746 B.n562 B.n84 256.663
R747 B.n562 B.n83 256.663
R748 B.n562 B.n82 256.663
R749 B.n562 B.n81 256.663
R750 B.n562 B.n80 256.663
R751 B.n562 B.n79 256.663
R752 B.n562 B.n78 256.663
R753 B.n562 B.n77 256.663
R754 B.n562 B.n76 256.663
R755 B.n562 B.n75 256.663
R756 B.n562 B.n74 256.663
R757 B.n562 B.n73 256.663
R758 B.n562 B.n72 256.663
R759 B.n562 B.n71 256.663
R760 B.n562 B.n70 256.663
R761 B.n562 B.n69 256.663
R762 B.n301 B.n269 256.663
R763 B.n307 B.n269 256.663
R764 B.n309 B.n269 256.663
R765 B.n315 B.n269 256.663
R766 B.n317 B.n269 256.663
R767 B.n323 B.n269 256.663
R768 B.n325 B.n269 256.663
R769 B.n331 B.n269 256.663
R770 B.n333 B.n269 256.663
R771 B.n339 B.n269 256.663
R772 B.n341 B.n269 256.663
R773 B.n347 B.n269 256.663
R774 B.n349 B.n269 256.663
R775 B.n355 B.n269 256.663
R776 B.n357 B.n269 256.663
R777 B.n364 B.n269 256.663
R778 B.n366 B.n269 256.663
R779 B.n372 B.n269 256.663
R780 B.n374 B.n269 256.663
R781 B.n380 B.n269 256.663
R782 B.n382 B.n269 256.663
R783 B.n388 B.n269 256.663
R784 B.n390 B.n269 256.663
R785 B.n396 B.n269 256.663
R786 B.n399 B.n269 256.663
R787 B.n282 B.t4 252.169
R788 B.n288 B.t12 252.169
R789 B.n97 B.t15 252.169
R790 B.n95 B.t8 252.169
R791 B.n282 B.t7 224.173
R792 B.n95 B.t10 224.173
R793 B.n288 B.t14 224.173
R794 B.n97 B.t16 224.173
R795 B.n406 B.n266 163.367
R796 B.n410 B.n266 163.367
R797 B.n410 B.n260 163.367
R798 B.n418 B.n260 163.367
R799 B.n418 B.n258 163.367
R800 B.n422 B.n258 163.367
R801 B.n422 B.n252 163.367
R802 B.n430 B.n252 163.367
R803 B.n430 B.n250 163.367
R804 B.n434 B.n250 163.367
R805 B.n434 B.n244 163.367
R806 B.n442 B.n244 163.367
R807 B.n442 B.n242 163.367
R808 B.n446 B.n242 163.367
R809 B.n446 B.n236 163.367
R810 B.n454 B.n236 163.367
R811 B.n454 B.n234 163.367
R812 B.n458 B.n234 163.367
R813 B.n458 B.n228 163.367
R814 B.n466 B.n228 163.367
R815 B.n466 B.n226 163.367
R816 B.n470 B.n226 163.367
R817 B.n470 B.n220 163.367
R818 B.n478 B.n220 163.367
R819 B.n478 B.n218 163.367
R820 B.n482 B.n218 163.367
R821 B.n482 B.n212 163.367
R822 B.n491 B.n212 163.367
R823 B.n491 B.n210 163.367
R824 B.n495 B.n210 163.367
R825 B.n495 B.n205 163.367
R826 B.n504 B.n205 163.367
R827 B.n504 B.n203 163.367
R828 B.n508 B.n203 163.367
R829 B.n508 B.n2 163.367
R830 B.n636 B.n2 163.367
R831 B.n636 B.n3 163.367
R832 B.n632 B.n3 163.367
R833 B.n632 B.n9 163.367
R834 B.n628 B.n9 163.367
R835 B.n628 B.n11 163.367
R836 B.n624 B.n11 163.367
R837 B.n624 B.n15 163.367
R838 B.n620 B.n15 163.367
R839 B.n620 B.n17 163.367
R840 B.n616 B.n17 163.367
R841 B.n616 B.n23 163.367
R842 B.n612 B.n23 163.367
R843 B.n612 B.n25 163.367
R844 B.n608 B.n25 163.367
R845 B.n608 B.n30 163.367
R846 B.n604 B.n30 163.367
R847 B.n604 B.n32 163.367
R848 B.n600 B.n32 163.367
R849 B.n600 B.n37 163.367
R850 B.n596 B.n37 163.367
R851 B.n596 B.n39 163.367
R852 B.n592 B.n39 163.367
R853 B.n592 B.n44 163.367
R854 B.n588 B.n44 163.367
R855 B.n588 B.n46 163.367
R856 B.n584 B.n46 163.367
R857 B.n584 B.n51 163.367
R858 B.n580 B.n51 163.367
R859 B.n580 B.n53 163.367
R860 B.n576 B.n53 163.367
R861 B.n576 B.n58 163.367
R862 B.n572 B.n58 163.367
R863 B.n572 B.n60 163.367
R864 B.n568 B.n60 163.367
R865 B.n568 B.n65 163.367
R866 B.n564 B.n65 163.367
R867 B.n302 B.n300 163.367
R868 B.n306 B.n300 163.367
R869 B.n310 B.n308 163.367
R870 B.n314 B.n298 163.367
R871 B.n318 B.n316 163.367
R872 B.n322 B.n296 163.367
R873 B.n326 B.n324 163.367
R874 B.n330 B.n294 163.367
R875 B.n334 B.n332 163.367
R876 B.n338 B.n292 163.367
R877 B.n342 B.n340 163.367
R878 B.n346 B.n287 163.367
R879 B.n350 B.n348 163.367
R880 B.n354 B.n285 163.367
R881 B.n358 B.n356 163.367
R882 B.n363 B.n281 163.367
R883 B.n367 B.n365 163.367
R884 B.n371 B.n279 163.367
R885 B.n375 B.n373 163.367
R886 B.n379 B.n277 163.367
R887 B.n383 B.n381 163.367
R888 B.n387 B.n275 163.367
R889 B.n391 B.n389 163.367
R890 B.n395 B.n273 163.367
R891 B.n398 B.n397 163.367
R892 B.n400 B.n270 163.367
R893 B.n404 B.n264 163.367
R894 B.n412 B.n264 163.367
R895 B.n412 B.n262 163.367
R896 B.n416 B.n262 163.367
R897 B.n416 B.n256 163.367
R898 B.n424 B.n256 163.367
R899 B.n424 B.n254 163.367
R900 B.n428 B.n254 163.367
R901 B.n428 B.n248 163.367
R902 B.n436 B.n248 163.367
R903 B.n436 B.n246 163.367
R904 B.n440 B.n246 163.367
R905 B.n440 B.n240 163.367
R906 B.n448 B.n240 163.367
R907 B.n448 B.n238 163.367
R908 B.n452 B.n238 163.367
R909 B.n452 B.n232 163.367
R910 B.n460 B.n232 163.367
R911 B.n460 B.n230 163.367
R912 B.n464 B.n230 163.367
R913 B.n464 B.n224 163.367
R914 B.n472 B.n224 163.367
R915 B.n472 B.n222 163.367
R916 B.n476 B.n222 163.367
R917 B.n476 B.n216 163.367
R918 B.n484 B.n216 163.367
R919 B.n484 B.n214 163.367
R920 B.n488 B.n214 163.367
R921 B.n488 B.n209 163.367
R922 B.n497 B.n209 163.367
R923 B.n497 B.n207 163.367
R924 B.n502 B.n207 163.367
R925 B.n502 B.n201 163.367
R926 B.n510 B.n201 163.367
R927 B.n511 B.n510 163.367
R928 B.n511 B.n5 163.367
R929 B.n6 B.n5 163.367
R930 B.n7 B.n6 163.367
R931 B.n516 B.n7 163.367
R932 B.n516 B.n12 163.367
R933 B.n13 B.n12 163.367
R934 B.n14 B.n13 163.367
R935 B.n521 B.n14 163.367
R936 B.n521 B.n19 163.367
R937 B.n20 B.n19 163.367
R938 B.n21 B.n20 163.367
R939 B.n526 B.n21 163.367
R940 B.n526 B.n26 163.367
R941 B.n27 B.n26 163.367
R942 B.n28 B.n27 163.367
R943 B.n531 B.n28 163.367
R944 B.n531 B.n33 163.367
R945 B.n34 B.n33 163.367
R946 B.n35 B.n34 163.367
R947 B.n536 B.n35 163.367
R948 B.n536 B.n40 163.367
R949 B.n41 B.n40 163.367
R950 B.n42 B.n41 163.367
R951 B.n541 B.n42 163.367
R952 B.n541 B.n47 163.367
R953 B.n48 B.n47 163.367
R954 B.n49 B.n48 163.367
R955 B.n546 B.n49 163.367
R956 B.n546 B.n54 163.367
R957 B.n55 B.n54 163.367
R958 B.n56 B.n55 163.367
R959 B.n551 B.n56 163.367
R960 B.n551 B.n61 163.367
R961 B.n62 B.n61 163.367
R962 B.n63 B.n62 163.367
R963 B.n556 B.n63 163.367
R964 B.n556 B.n68 163.367
R965 B.n101 B.n100 163.367
R966 B.n105 B.n104 163.367
R967 B.n109 B.n108 163.367
R968 B.n113 B.n112 163.367
R969 B.n117 B.n116 163.367
R970 B.n121 B.n120 163.367
R971 B.n125 B.n124 163.367
R972 B.n129 B.n128 163.367
R973 B.n133 B.n132 163.367
R974 B.n137 B.n136 163.367
R975 B.n142 B.n141 163.367
R976 B.n146 B.n145 163.367
R977 B.n150 B.n149 163.367
R978 B.n154 B.n153 163.367
R979 B.n158 B.n157 163.367
R980 B.n163 B.n162 163.367
R981 B.n167 B.n166 163.367
R982 B.n171 B.n170 163.367
R983 B.n175 B.n174 163.367
R984 B.n179 B.n178 163.367
R985 B.n183 B.n182 163.367
R986 B.n187 B.n186 163.367
R987 B.n191 B.n190 163.367
R988 B.n195 B.n194 163.367
R989 B.n197 B.n94 163.367
R990 B.n283 B.t6 163.276
R991 B.n96 B.t11 163.276
R992 B.n289 B.t13 163.276
R993 B.n98 B.t17 163.276
R994 B.n405 B.n269 117.573
R995 B.n563 B.n562 117.573
R996 B.n405 B.n265 72.0275
R997 B.n411 B.n265 72.0275
R998 B.n411 B.n261 72.0275
R999 B.n417 B.n261 72.0275
R1000 B.n417 B.n257 72.0275
R1001 B.n423 B.n257 72.0275
R1002 B.n423 B.n253 72.0275
R1003 B.n429 B.n253 72.0275
R1004 B.n435 B.n249 72.0275
R1005 B.n435 B.n245 72.0275
R1006 B.n441 B.n245 72.0275
R1007 B.n441 B.n241 72.0275
R1008 B.n447 B.n241 72.0275
R1009 B.n447 B.n237 72.0275
R1010 B.n453 B.n237 72.0275
R1011 B.n453 B.n233 72.0275
R1012 B.n459 B.n233 72.0275
R1013 B.n459 B.n229 72.0275
R1014 B.n465 B.n229 72.0275
R1015 B.n471 B.n225 72.0275
R1016 B.n471 B.n221 72.0275
R1017 B.n477 B.n221 72.0275
R1018 B.n477 B.n217 72.0275
R1019 B.n483 B.n217 72.0275
R1020 B.n483 B.n213 72.0275
R1021 B.n490 B.n213 72.0275
R1022 B.n490 B.n489 72.0275
R1023 B.n496 B.n206 72.0275
R1024 B.n503 B.n206 72.0275
R1025 B.n503 B.n202 72.0275
R1026 B.n509 B.n202 72.0275
R1027 B.n509 B.n4 72.0275
R1028 B.n635 B.n4 72.0275
R1029 B.n635 B.n634 72.0275
R1030 B.n634 B.n633 72.0275
R1031 B.n633 B.n8 72.0275
R1032 B.n627 B.n8 72.0275
R1033 B.n627 B.n626 72.0275
R1034 B.n626 B.n625 72.0275
R1035 B.n619 B.n18 72.0275
R1036 B.n619 B.n618 72.0275
R1037 B.n618 B.n617 72.0275
R1038 B.n617 B.n22 72.0275
R1039 B.n611 B.n22 72.0275
R1040 B.n611 B.n610 72.0275
R1041 B.n610 B.n609 72.0275
R1042 B.n609 B.n29 72.0275
R1043 B.n603 B.n602 72.0275
R1044 B.n602 B.n601 72.0275
R1045 B.n601 B.n36 72.0275
R1046 B.n595 B.n36 72.0275
R1047 B.n595 B.n594 72.0275
R1048 B.n594 B.n593 72.0275
R1049 B.n593 B.n43 72.0275
R1050 B.n587 B.n43 72.0275
R1051 B.n587 B.n586 72.0275
R1052 B.n586 B.n585 72.0275
R1053 B.n585 B.n50 72.0275
R1054 B.n579 B.n578 72.0275
R1055 B.n578 B.n577 72.0275
R1056 B.n577 B.n57 72.0275
R1057 B.n571 B.n57 72.0275
R1058 B.n571 B.n570 72.0275
R1059 B.n570 B.n569 72.0275
R1060 B.n569 B.n64 72.0275
R1061 B.n563 B.n64 72.0275
R1062 B.n301 B.n268 71.676
R1063 B.n307 B.n306 71.676
R1064 B.n310 B.n309 71.676
R1065 B.n315 B.n314 71.676
R1066 B.n318 B.n317 71.676
R1067 B.n323 B.n322 71.676
R1068 B.n326 B.n325 71.676
R1069 B.n331 B.n330 71.676
R1070 B.n334 B.n333 71.676
R1071 B.n339 B.n338 71.676
R1072 B.n342 B.n341 71.676
R1073 B.n347 B.n346 71.676
R1074 B.n350 B.n349 71.676
R1075 B.n355 B.n354 71.676
R1076 B.n358 B.n357 71.676
R1077 B.n364 B.n363 71.676
R1078 B.n367 B.n366 71.676
R1079 B.n372 B.n371 71.676
R1080 B.n375 B.n374 71.676
R1081 B.n380 B.n379 71.676
R1082 B.n383 B.n382 71.676
R1083 B.n388 B.n387 71.676
R1084 B.n391 B.n390 71.676
R1085 B.n396 B.n395 71.676
R1086 B.n399 B.n398 71.676
R1087 B.n69 B.n67 71.676
R1088 B.n101 B.n70 71.676
R1089 B.n105 B.n71 71.676
R1090 B.n109 B.n72 71.676
R1091 B.n113 B.n73 71.676
R1092 B.n117 B.n74 71.676
R1093 B.n121 B.n75 71.676
R1094 B.n125 B.n76 71.676
R1095 B.n129 B.n77 71.676
R1096 B.n133 B.n78 71.676
R1097 B.n137 B.n79 71.676
R1098 B.n142 B.n80 71.676
R1099 B.n146 B.n81 71.676
R1100 B.n150 B.n82 71.676
R1101 B.n154 B.n83 71.676
R1102 B.n158 B.n84 71.676
R1103 B.n163 B.n85 71.676
R1104 B.n167 B.n86 71.676
R1105 B.n171 B.n87 71.676
R1106 B.n175 B.n88 71.676
R1107 B.n179 B.n89 71.676
R1108 B.n183 B.n90 71.676
R1109 B.n187 B.n91 71.676
R1110 B.n191 B.n92 71.676
R1111 B.n195 B.n93 71.676
R1112 B.n561 B.n94 71.676
R1113 B.n561 B.n560 71.676
R1114 B.n197 B.n93 71.676
R1115 B.n194 B.n92 71.676
R1116 B.n190 B.n91 71.676
R1117 B.n186 B.n90 71.676
R1118 B.n182 B.n89 71.676
R1119 B.n178 B.n88 71.676
R1120 B.n174 B.n87 71.676
R1121 B.n170 B.n86 71.676
R1122 B.n166 B.n85 71.676
R1123 B.n162 B.n84 71.676
R1124 B.n157 B.n83 71.676
R1125 B.n153 B.n82 71.676
R1126 B.n149 B.n81 71.676
R1127 B.n145 B.n80 71.676
R1128 B.n141 B.n79 71.676
R1129 B.n136 B.n78 71.676
R1130 B.n132 B.n77 71.676
R1131 B.n128 B.n76 71.676
R1132 B.n124 B.n75 71.676
R1133 B.n120 B.n74 71.676
R1134 B.n116 B.n73 71.676
R1135 B.n112 B.n72 71.676
R1136 B.n108 B.n71 71.676
R1137 B.n104 B.n70 71.676
R1138 B.n100 B.n69 71.676
R1139 B.n302 B.n301 71.676
R1140 B.n308 B.n307 71.676
R1141 B.n309 B.n298 71.676
R1142 B.n316 B.n315 71.676
R1143 B.n317 B.n296 71.676
R1144 B.n324 B.n323 71.676
R1145 B.n325 B.n294 71.676
R1146 B.n332 B.n331 71.676
R1147 B.n333 B.n292 71.676
R1148 B.n340 B.n339 71.676
R1149 B.n341 B.n287 71.676
R1150 B.n348 B.n347 71.676
R1151 B.n349 B.n285 71.676
R1152 B.n356 B.n355 71.676
R1153 B.n357 B.n281 71.676
R1154 B.n365 B.n364 71.676
R1155 B.n366 B.n279 71.676
R1156 B.n373 B.n372 71.676
R1157 B.n374 B.n277 71.676
R1158 B.n381 B.n380 71.676
R1159 B.n382 B.n275 71.676
R1160 B.n389 B.n388 71.676
R1161 B.n390 B.n273 71.676
R1162 B.n397 B.n396 71.676
R1163 B.n400 B.n399 71.676
R1164 B.t5 B.n249 64.6129
R1165 B.t9 B.n50 64.6129
R1166 B.n283 B.n282 60.8975
R1167 B.n289 B.n288 60.8975
R1168 B.n98 B.n97 60.8975
R1169 B.n96 B.n95 60.8975
R1170 B.n361 B.n283 59.5399
R1171 B.n290 B.n289 59.5399
R1172 B.n139 B.n98 59.5399
R1173 B.n160 B.n96 59.5399
R1174 B.n489 B.t3 56.1392
R1175 B.n18 B.t0 56.1392
R1176 B.n465 B.t1 39.1916
R1177 B.n603 B.t2 39.1916
R1178 B.t1 B.n225 32.8363
R1179 B.t2 B.n29 32.8363
R1180 B.n565 B.n66 32.0005
R1181 B.n559 B.n558 32.0005
R1182 B.n403 B.n402 32.0005
R1183 B.n407 B.n267 32.0005
R1184 B B.n637 18.0485
R1185 B.n496 B.t3 15.8888
R1186 B.n625 B.t0 15.8888
R1187 B.n99 B.n66 10.6151
R1188 B.n102 B.n99 10.6151
R1189 B.n103 B.n102 10.6151
R1190 B.n106 B.n103 10.6151
R1191 B.n107 B.n106 10.6151
R1192 B.n110 B.n107 10.6151
R1193 B.n111 B.n110 10.6151
R1194 B.n114 B.n111 10.6151
R1195 B.n115 B.n114 10.6151
R1196 B.n118 B.n115 10.6151
R1197 B.n119 B.n118 10.6151
R1198 B.n122 B.n119 10.6151
R1199 B.n123 B.n122 10.6151
R1200 B.n126 B.n123 10.6151
R1201 B.n127 B.n126 10.6151
R1202 B.n130 B.n127 10.6151
R1203 B.n131 B.n130 10.6151
R1204 B.n134 B.n131 10.6151
R1205 B.n135 B.n134 10.6151
R1206 B.n138 B.n135 10.6151
R1207 B.n143 B.n140 10.6151
R1208 B.n144 B.n143 10.6151
R1209 B.n147 B.n144 10.6151
R1210 B.n148 B.n147 10.6151
R1211 B.n151 B.n148 10.6151
R1212 B.n152 B.n151 10.6151
R1213 B.n155 B.n152 10.6151
R1214 B.n156 B.n155 10.6151
R1215 B.n159 B.n156 10.6151
R1216 B.n164 B.n161 10.6151
R1217 B.n165 B.n164 10.6151
R1218 B.n168 B.n165 10.6151
R1219 B.n169 B.n168 10.6151
R1220 B.n172 B.n169 10.6151
R1221 B.n173 B.n172 10.6151
R1222 B.n176 B.n173 10.6151
R1223 B.n177 B.n176 10.6151
R1224 B.n180 B.n177 10.6151
R1225 B.n181 B.n180 10.6151
R1226 B.n184 B.n181 10.6151
R1227 B.n185 B.n184 10.6151
R1228 B.n188 B.n185 10.6151
R1229 B.n189 B.n188 10.6151
R1230 B.n192 B.n189 10.6151
R1231 B.n193 B.n192 10.6151
R1232 B.n196 B.n193 10.6151
R1233 B.n198 B.n196 10.6151
R1234 B.n199 B.n198 10.6151
R1235 B.n559 B.n199 10.6151
R1236 B.n403 B.n263 10.6151
R1237 B.n413 B.n263 10.6151
R1238 B.n414 B.n413 10.6151
R1239 B.n415 B.n414 10.6151
R1240 B.n415 B.n255 10.6151
R1241 B.n425 B.n255 10.6151
R1242 B.n426 B.n425 10.6151
R1243 B.n427 B.n426 10.6151
R1244 B.n427 B.n247 10.6151
R1245 B.n437 B.n247 10.6151
R1246 B.n438 B.n437 10.6151
R1247 B.n439 B.n438 10.6151
R1248 B.n439 B.n239 10.6151
R1249 B.n449 B.n239 10.6151
R1250 B.n450 B.n449 10.6151
R1251 B.n451 B.n450 10.6151
R1252 B.n451 B.n231 10.6151
R1253 B.n461 B.n231 10.6151
R1254 B.n462 B.n461 10.6151
R1255 B.n463 B.n462 10.6151
R1256 B.n463 B.n223 10.6151
R1257 B.n473 B.n223 10.6151
R1258 B.n474 B.n473 10.6151
R1259 B.n475 B.n474 10.6151
R1260 B.n475 B.n215 10.6151
R1261 B.n485 B.n215 10.6151
R1262 B.n486 B.n485 10.6151
R1263 B.n487 B.n486 10.6151
R1264 B.n487 B.n208 10.6151
R1265 B.n498 B.n208 10.6151
R1266 B.n499 B.n498 10.6151
R1267 B.n501 B.n499 10.6151
R1268 B.n501 B.n500 10.6151
R1269 B.n500 B.n200 10.6151
R1270 B.n512 B.n200 10.6151
R1271 B.n513 B.n512 10.6151
R1272 B.n514 B.n513 10.6151
R1273 B.n515 B.n514 10.6151
R1274 B.n517 B.n515 10.6151
R1275 B.n518 B.n517 10.6151
R1276 B.n519 B.n518 10.6151
R1277 B.n520 B.n519 10.6151
R1278 B.n522 B.n520 10.6151
R1279 B.n523 B.n522 10.6151
R1280 B.n524 B.n523 10.6151
R1281 B.n525 B.n524 10.6151
R1282 B.n527 B.n525 10.6151
R1283 B.n528 B.n527 10.6151
R1284 B.n529 B.n528 10.6151
R1285 B.n530 B.n529 10.6151
R1286 B.n532 B.n530 10.6151
R1287 B.n533 B.n532 10.6151
R1288 B.n534 B.n533 10.6151
R1289 B.n535 B.n534 10.6151
R1290 B.n537 B.n535 10.6151
R1291 B.n538 B.n537 10.6151
R1292 B.n539 B.n538 10.6151
R1293 B.n540 B.n539 10.6151
R1294 B.n542 B.n540 10.6151
R1295 B.n543 B.n542 10.6151
R1296 B.n544 B.n543 10.6151
R1297 B.n545 B.n544 10.6151
R1298 B.n547 B.n545 10.6151
R1299 B.n548 B.n547 10.6151
R1300 B.n549 B.n548 10.6151
R1301 B.n550 B.n549 10.6151
R1302 B.n552 B.n550 10.6151
R1303 B.n553 B.n552 10.6151
R1304 B.n554 B.n553 10.6151
R1305 B.n555 B.n554 10.6151
R1306 B.n557 B.n555 10.6151
R1307 B.n558 B.n557 10.6151
R1308 B.n303 B.n267 10.6151
R1309 B.n304 B.n303 10.6151
R1310 B.n305 B.n304 10.6151
R1311 B.n305 B.n299 10.6151
R1312 B.n311 B.n299 10.6151
R1313 B.n312 B.n311 10.6151
R1314 B.n313 B.n312 10.6151
R1315 B.n313 B.n297 10.6151
R1316 B.n319 B.n297 10.6151
R1317 B.n320 B.n319 10.6151
R1318 B.n321 B.n320 10.6151
R1319 B.n321 B.n295 10.6151
R1320 B.n327 B.n295 10.6151
R1321 B.n328 B.n327 10.6151
R1322 B.n329 B.n328 10.6151
R1323 B.n329 B.n293 10.6151
R1324 B.n335 B.n293 10.6151
R1325 B.n336 B.n335 10.6151
R1326 B.n337 B.n336 10.6151
R1327 B.n337 B.n291 10.6151
R1328 B.n344 B.n343 10.6151
R1329 B.n345 B.n344 10.6151
R1330 B.n345 B.n286 10.6151
R1331 B.n351 B.n286 10.6151
R1332 B.n352 B.n351 10.6151
R1333 B.n353 B.n352 10.6151
R1334 B.n353 B.n284 10.6151
R1335 B.n359 B.n284 10.6151
R1336 B.n360 B.n359 10.6151
R1337 B.n362 B.n280 10.6151
R1338 B.n368 B.n280 10.6151
R1339 B.n369 B.n368 10.6151
R1340 B.n370 B.n369 10.6151
R1341 B.n370 B.n278 10.6151
R1342 B.n376 B.n278 10.6151
R1343 B.n377 B.n376 10.6151
R1344 B.n378 B.n377 10.6151
R1345 B.n378 B.n276 10.6151
R1346 B.n384 B.n276 10.6151
R1347 B.n385 B.n384 10.6151
R1348 B.n386 B.n385 10.6151
R1349 B.n386 B.n274 10.6151
R1350 B.n392 B.n274 10.6151
R1351 B.n393 B.n392 10.6151
R1352 B.n394 B.n393 10.6151
R1353 B.n394 B.n272 10.6151
R1354 B.n272 B.n271 10.6151
R1355 B.n401 B.n271 10.6151
R1356 B.n402 B.n401 10.6151
R1357 B.n408 B.n407 10.6151
R1358 B.n409 B.n408 10.6151
R1359 B.n409 B.n259 10.6151
R1360 B.n419 B.n259 10.6151
R1361 B.n420 B.n419 10.6151
R1362 B.n421 B.n420 10.6151
R1363 B.n421 B.n251 10.6151
R1364 B.n431 B.n251 10.6151
R1365 B.n432 B.n431 10.6151
R1366 B.n433 B.n432 10.6151
R1367 B.n433 B.n243 10.6151
R1368 B.n443 B.n243 10.6151
R1369 B.n444 B.n443 10.6151
R1370 B.n445 B.n444 10.6151
R1371 B.n445 B.n235 10.6151
R1372 B.n455 B.n235 10.6151
R1373 B.n456 B.n455 10.6151
R1374 B.n457 B.n456 10.6151
R1375 B.n457 B.n227 10.6151
R1376 B.n467 B.n227 10.6151
R1377 B.n468 B.n467 10.6151
R1378 B.n469 B.n468 10.6151
R1379 B.n469 B.n219 10.6151
R1380 B.n479 B.n219 10.6151
R1381 B.n480 B.n479 10.6151
R1382 B.n481 B.n480 10.6151
R1383 B.n481 B.n211 10.6151
R1384 B.n492 B.n211 10.6151
R1385 B.n493 B.n492 10.6151
R1386 B.n494 B.n493 10.6151
R1387 B.n494 B.n204 10.6151
R1388 B.n505 B.n204 10.6151
R1389 B.n506 B.n505 10.6151
R1390 B.n507 B.n506 10.6151
R1391 B.n507 B.n0 10.6151
R1392 B.n631 B.n1 10.6151
R1393 B.n631 B.n630 10.6151
R1394 B.n630 B.n629 10.6151
R1395 B.n629 B.n10 10.6151
R1396 B.n623 B.n10 10.6151
R1397 B.n623 B.n622 10.6151
R1398 B.n622 B.n621 10.6151
R1399 B.n621 B.n16 10.6151
R1400 B.n615 B.n16 10.6151
R1401 B.n615 B.n614 10.6151
R1402 B.n614 B.n613 10.6151
R1403 B.n613 B.n24 10.6151
R1404 B.n607 B.n24 10.6151
R1405 B.n607 B.n606 10.6151
R1406 B.n606 B.n605 10.6151
R1407 B.n605 B.n31 10.6151
R1408 B.n599 B.n31 10.6151
R1409 B.n599 B.n598 10.6151
R1410 B.n598 B.n597 10.6151
R1411 B.n597 B.n38 10.6151
R1412 B.n591 B.n38 10.6151
R1413 B.n591 B.n590 10.6151
R1414 B.n590 B.n589 10.6151
R1415 B.n589 B.n45 10.6151
R1416 B.n583 B.n45 10.6151
R1417 B.n583 B.n582 10.6151
R1418 B.n582 B.n581 10.6151
R1419 B.n581 B.n52 10.6151
R1420 B.n575 B.n52 10.6151
R1421 B.n575 B.n574 10.6151
R1422 B.n574 B.n573 10.6151
R1423 B.n573 B.n59 10.6151
R1424 B.n567 B.n59 10.6151
R1425 B.n567 B.n566 10.6151
R1426 B.n566 B.n565 10.6151
R1427 B.n139 B.n138 9.36635
R1428 B.n161 B.n160 9.36635
R1429 B.n291 B.n290 9.36635
R1430 B.n362 B.n361 9.36635
R1431 B.n429 B.t5 7.41504
R1432 B.n579 B.t9 7.41504
R1433 B.n637 B.n0 2.81026
R1434 B.n637 B.n1 2.81026
R1435 B.n140 B.n139 1.24928
R1436 B.n160 B.n159 1.24928
R1437 B.n343 B.n290 1.24928
R1438 B.n361 B.n360 1.24928
R1439 VP.n16 VP.n0 161.3
R1440 VP.n15 VP.n14 161.3
R1441 VP.n13 VP.n1 161.3
R1442 VP.n12 VP.n11 161.3
R1443 VP.n10 VP.n2 161.3
R1444 VP.n9 VP.n8 161.3
R1445 VP.n7 VP.n3 161.3
R1446 VP.n6 VP.n5 107.332
R1447 VP.n18 VP.n17 107.332
R1448 VP.n4 VP.t1 78.8747
R1449 VP.n4 VP.t0 77.9842
R1450 VP.n6 VP.n4 45.211
R1451 VP.n5 VP.t2 43.8265
R1452 VP.n17 VP.t3 43.8265
R1453 VP.n11 VP.n10 40.4934
R1454 VP.n11 VP.n1 40.4934
R1455 VP.n9 VP.n3 24.4675
R1456 VP.n10 VP.n9 24.4675
R1457 VP.n15 VP.n1 24.4675
R1458 VP.n16 VP.n15 24.4675
R1459 VP.n5 VP.n3 3.42588
R1460 VP.n17 VP.n16 3.42588
R1461 VP.n7 VP.n6 0.278367
R1462 VP.n18 VP.n0 0.278367
R1463 VP.n8 VP.n7 0.189894
R1464 VP.n8 VP.n2 0.189894
R1465 VP.n12 VP.n2 0.189894
R1466 VP.n13 VP.n12 0.189894
R1467 VP.n14 VP.n13 0.189894
R1468 VP.n14 VP.n0 0.189894
R1469 VP VP.n18 0.153454
R1470 VDD1 VDD1.n1 108.105
R1471 VDD1 VDD1.n0 71.396
R1472 VDD1.n0 VDD1.t2 3.87526
R1473 VDD1.n0 VDD1.t3 3.87526
R1474 VDD1.n1 VDD1.t1 3.87526
R1475 VDD1.n1 VDD1.t0 3.87526
C0 VDD2 VP 0.411581f
C1 VDD2 VTAIL 3.91049f
C2 VDD2 VDD1 1.0723f
C3 VP VN 5.06612f
C4 VN VTAIL 2.62001f
C5 VN VDD1 0.149028f
C6 VP VTAIL 2.63412f
C7 VP VDD1 2.49866f
C8 VDD2 VN 2.24103f
C9 VTAIL VDD1 3.85487f
C10 VDD2 B 3.350941f
C11 VDD1 B 6.95544f
C12 VTAIL B 5.7721f
C13 VN B 10.487041f
C14 VP B 8.760167f
C15 VDD1.t2 B 0.115664f
C16 VDD1.t3 B 0.115664f
C17 VDD1.n0 B 0.957503f
C18 VDD1.t1 B 0.115664f
C19 VDD1.t0 B 0.115664f
C20 VDD1.n1 B 1.41755f
C21 VP.n0 B 0.038455f
C22 VP.t3 B 1.09718f
C23 VP.n1 B 0.057971f
C24 VP.n2 B 0.029168f
C25 VP.n3 B 0.03128f
C26 VP.t0 B 1.3659f
C27 VP.t1 B 1.37268f
C28 VP.n4 B 2.23638f
C29 VP.t2 B 1.09718f
C30 VP.n5 B 0.513581f
C31 VP.n6 B 1.37919f
C32 VP.n7 B 0.038455f
C33 VP.n8 B 0.029168f
C34 VP.n9 B 0.054362f
C35 VP.n10 B 0.057971f
C36 VP.n11 B 0.02358f
C37 VP.n12 B 0.029168f
C38 VP.n13 B 0.029168f
C39 VP.n14 B 0.029168f
C40 VP.n15 B 0.054362f
C41 VP.n16 B 0.03128f
C42 VP.n17 B 0.513581f
C43 VP.n18 B 0.054181f
C44 VTAIL.n0 B 0.011689f
C45 VTAIL.n1 B 0.026342f
C46 VTAIL.n2 B 0.0118f
C47 VTAIL.n3 B 0.02074f
C48 VTAIL.n4 B 0.011145f
C49 VTAIL.n5 B 0.026342f
C50 VTAIL.n6 B 0.0118f
C51 VTAIL.n7 B 0.095049f
C52 VTAIL.t6 B 0.043927f
C53 VTAIL.n8 B 0.019757f
C54 VTAIL.n9 B 0.018618f
C55 VTAIL.n10 B 0.011145f
C56 VTAIL.n11 B 0.410126f
C57 VTAIL.n12 B 0.02074f
C58 VTAIL.n13 B 0.011145f
C59 VTAIL.n14 B 0.0118f
C60 VTAIL.n15 B 0.026342f
C61 VTAIL.n16 B 0.026342f
C62 VTAIL.n17 B 0.0118f
C63 VTAIL.n18 B 0.011145f
C64 VTAIL.n19 B 0.02074f
C65 VTAIL.n20 B 0.053323f
C66 VTAIL.n21 B 0.011145f
C67 VTAIL.n22 B 0.0118f
C68 VTAIL.n23 B 0.05183f
C69 VTAIL.n24 B 0.044099f
C70 VTAIL.n25 B 0.144892f
C71 VTAIL.n26 B 0.011689f
C72 VTAIL.n27 B 0.026342f
C73 VTAIL.n28 B 0.0118f
C74 VTAIL.n29 B 0.02074f
C75 VTAIL.n30 B 0.011145f
C76 VTAIL.n31 B 0.026342f
C77 VTAIL.n32 B 0.0118f
C78 VTAIL.n33 B 0.095049f
C79 VTAIL.t7 B 0.043927f
C80 VTAIL.n34 B 0.019757f
C81 VTAIL.n35 B 0.018618f
C82 VTAIL.n36 B 0.011145f
C83 VTAIL.n37 B 0.410126f
C84 VTAIL.n38 B 0.02074f
C85 VTAIL.n39 B 0.011145f
C86 VTAIL.n40 B 0.0118f
C87 VTAIL.n41 B 0.026342f
C88 VTAIL.n42 B 0.026342f
C89 VTAIL.n43 B 0.0118f
C90 VTAIL.n44 B 0.011145f
C91 VTAIL.n45 B 0.02074f
C92 VTAIL.n46 B 0.053323f
C93 VTAIL.n47 B 0.011145f
C94 VTAIL.n48 B 0.0118f
C95 VTAIL.n49 B 0.05183f
C96 VTAIL.n50 B 0.044099f
C97 VTAIL.n51 B 0.231453f
C98 VTAIL.n52 B 0.011689f
C99 VTAIL.n53 B 0.026342f
C100 VTAIL.n54 B 0.0118f
C101 VTAIL.n55 B 0.02074f
C102 VTAIL.n56 B 0.011145f
C103 VTAIL.n57 B 0.026342f
C104 VTAIL.n58 B 0.0118f
C105 VTAIL.n59 B 0.095049f
C106 VTAIL.t1 B 0.043927f
C107 VTAIL.n60 B 0.019757f
C108 VTAIL.n61 B 0.018618f
C109 VTAIL.n62 B 0.011145f
C110 VTAIL.n63 B 0.410126f
C111 VTAIL.n64 B 0.02074f
C112 VTAIL.n65 B 0.011145f
C113 VTAIL.n66 B 0.0118f
C114 VTAIL.n67 B 0.026342f
C115 VTAIL.n68 B 0.026342f
C116 VTAIL.n69 B 0.0118f
C117 VTAIL.n70 B 0.011145f
C118 VTAIL.n71 B 0.02074f
C119 VTAIL.n72 B 0.053323f
C120 VTAIL.n73 B 0.011145f
C121 VTAIL.n74 B 0.0118f
C122 VTAIL.n75 B 0.05183f
C123 VTAIL.n76 B 0.044099f
C124 VTAIL.n77 B 0.957079f
C125 VTAIL.n78 B 0.011689f
C126 VTAIL.n79 B 0.026342f
C127 VTAIL.n80 B 0.0118f
C128 VTAIL.n81 B 0.02074f
C129 VTAIL.n82 B 0.011145f
C130 VTAIL.n83 B 0.026342f
C131 VTAIL.n84 B 0.0118f
C132 VTAIL.n85 B 0.095049f
C133 VTAIL.t3 B 0.043927f
C134 VTAIL.n86 B 0.019757f
C135 VTAIL.n87 B 0.018618f
C136 VTAIL.n88 B 0.011145f
C137 VTAIL.n89 B 0.410126f
C138 VTAIL.n90 B 0.02074f
C139 VTAIL.n91 B 0.011145f
C140 VTAIL.n92 B 0.0118f
C141 VTAIL.n93 B 0.026342f
C142 VTAIL.n94 B 0.026342f
C143 VTAIL.n95 B 0.0118f
C144 VTAIL.n96 B 0.011145f
C145 VTAIL.n97 B 0.02074f
C146 VTAIL.n98 B 0.053323f
C147 VTAIL.n99 B 0.011145f
C148 VTAIL.n100 B 0.0118f
C149 VTAIL.n101 B 0.05183f
C150 VTAIL.n102 B 0.044099f
C151 VTAIL.n103 B 0.957079f
C152 VTAIL.n104 B 0.011689f
C153 VTAIL.n105 B 0.026342f
C154 VTAIL.n106 B 0.0118f
C155 VTAIL.n107 B 0.02074f
C156 VTAIL.n108 B 0.011145f
C157 VTAIL.n109 B 0.026342f
C158 VTAIL.n110 B 0.0118f
C159 VTAIL.n111 B 0.095049f
C160 VTAIL.t4 B 0.043927f
C161 VTAIL.n112 B 0.019757f
C162 VTAIL.n113 B 0.018618f
C163 VTAIL.n114 B 0.011145f
C164 VTAIL.n115 B 0.410126f
C165 VTAIL.n116 B 0.02074f
C166 VTAIL.n117 B 0.011145f
C167 VTAIL.n118 B 0.0118f
C168 VTAIL.n119 B 0.026342f
C169 VTAIL.n120 B 0.026342f
C170 VTAIL.n121 B 0.0118f
C171 VTAIL.n122 B 0.011145f
C172 VTAIL.n123 B 0.02074f
C173 VTAIL.n124 B 0.053323f
C174 VTAIL.n125 B 0.011145f
C175 VTAIL.n126 B 0.0118f
C176 VTAIL.n127 B 0.05183f
C177 VTAIL.n128 B 0.044099f
C178 VTAIL.n129 B 0.231453f
C179 VTAIL.n130 B 0.011689f
C180 VTAIL.n131 B 0.026342f
C181 VTAIL.n132 B 0.0118f
C182 VTAIL.n133 B 0.02074f
C183 VTAIL.n134 B 0.011145f
C184 VTAIL.n135 B 0.026342f
C185 VTAIL.n136 B 0.0118f
C186 VTAIL.n137 B 0.095049f
C187 VTAIL.t0 B 0.043927f
C188 VTAIL.n138 B 0.019757f
C189 VTAIL.n139 B 0.018618f
C190 VTAIL.n140 B 0.011145f
C191 VTAIL.n141 B 0.410126f
C192 VTAIL.n142 B 0.02074f
C193 VTAIL.n143 B 0.011145f
C194 VTAIL.n144 B 0.0118f
C195 VTAIL.n145 B 0.026342f
C196 VTAIL.n146 B 0.026342f
C197 VTAIL.n147 B 0.0118f
C198 VTAIL.n148 B 0.011145f
C199 VTAIL.n149 B 0.02074f
C200 VTAIL.n150 B 0.053323f
C201 VTAIL.n151 B 0.011145f
C202 VTAIL.n152 B 0.0118f
C203 VTAIL.n153 B 0.05183f
C204 VTAIL.n154 B 0.044099f
C205 VTAIL.n155 B 0.231453f
C206 VTAIL.n156 B 0.011689f
C207 VTAIL.n157 B 0.026342f
C208 VTAIL.n158 B 0.0118f
C209 VTAIL.n159 B 0.02074f
C210 VTAIL.n160 B 0.011145f
C211 VTAIL.n161 B 0.026342f
C212 VTAIL.n162 B 0.0118f
C213 VTAIL.n163 B 0.095049f
C214 VTAIL.t2 B 0.043927f
C215 VTAIL.n164 B 0.019757f
C216 VTAIL.n165 B 0.018618f
C217 VTAIL.n166 B 0.011145f
C218 VTAIL.n167 B 0.410126f
C219 VTAIL.n168 B 0.02074f
C220 VTAIL.n169 B 0.011145f
C221 VTAIL.n170 B 0.0118f
C222 VTAIL.n171 B 0.026342f
C223 VTAIL.n172 B 0.026342f
C224 VTAIL.n173 B 0.0118f
C225 VTAIL.n174 B 0.011145f
C226 VTAIL.n175 B 0.02074f
C227 VTAIL.n176 B 0.053323f
C228 VTAIL.n177 B 0.011145f
C229 VTAIL.n178 B 0.0118f
C230 VTAIL.n179 B 0.05183f
C231 VTAIL.n180 B 0.044099f
C232 VTAIL.n181 B 0.957079f
C233 VTAIL.n182 B 0.011689f
C234 VTAIL.n183 B 0.026342f
C235 VTAIL.n184 B 0.0118f
C236 VTAIL.n185 B 0.02074f
C237 VTAIL.n186 B 0.011145f
C238 VTAIL.n187 B 0.026342f
C239 VTAIL.n188 B 0.0118f
C240 VTAIL.n189 B 0.095049f
C241 VTAIL.t5 B 0.043927f
C242 VTAIL.n190 B 0.019757f
C243 VTAIL.n191 B 0.018618f
C244 VTAIL.n192 B 0.011145f
C245 VTAIL.n193 B 0.410126f
C246 VTAIL.n194 B 0.02074f
C247 VTAIL.n195 B 0.011145f
C248 VTAIL.n196 B 0.0118f
C249 VTAIL.n197 B 0.026342f
C250 VTAIL.n198 B 0.026342f
C251 VTAIL.n199 B 0.0118f
C252 VTAIL.n200 B 0.011145f
C253 VTAIL.n201 B 0.02074f
C254 VTAIL.n202 B 0.053323f
C255 VTAIL.n203 B 0.011145f
C256 VTAIL.n204 B 0.0118f
C257 VTAIL.n205 B 0.05183f
C258 VTAIL.n206 B 0.044099f
C259 VTAIL.n207 B 0.86274f
C260 VDD2.t2 B 0.112095f
C261 VDD2.t3 B 0.112095f
C262 VDD2.n0 B 1.35077f
C263 VDD2.t1 B 0.112095f
C264 VDD2.t0 B 0.112095f
C265 VDD2.n1 B 0.927577f
C266 VDD2.n2 B 3.12517f
C267 VN.t0 B 1.32698f
C268 VN.t1 B 1.32042f
C269 VN.n0 B 0.812597f
C270 VN.t2 B 1.32698f
C271 VN.t3 B 1.32042f
C272 VN.n1 B 2.17705f
.ends

