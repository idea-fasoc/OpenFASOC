* NGSPICE file created from diff_pair_sample_0165.ext - technology: sky130A

.subckt diff_pair_sample_0165 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X1 VTAIL.t4 VP.t0 VDD1.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X2 VDD1.t6 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=4.7034 ps=24.9 w=12.06 l=2.04
X3 VDD2.t7 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X4 VTAIL.t0 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X5 VTAIL.t13 VN.t2 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=1.9899 ps=12.39 w=12.06 l=2.04
X6 VDD1.t4 VP.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X7 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=0 ps=0 w=12.06 l=2.04
X8 VDD2.t4 VN.t3 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X9 VTAIL.t6 VP.t4 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=1.9899 ps=12.39 w=12.06 l=2.04
X10 VTAIL.t11 VN.t4 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=1.9899 ps=12.39 w=12.06 l=2.04
X11 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=0 ps=0 w=12.06 l=2.04
X12 VDD1.t2 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X13 VTAIL.t10 VN.t5 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=1.9899 ps=12.39 w=12.06 l=2.04
X14 VDD2.t0 VN.t6 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=4.7034 ps=24.9 w=12.06 l=2.04
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=0 ps=0 w=12.06 l=2.04
X16 VTAIL.t5 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=1.9899 ps=12.39 w=12.06 l=2.04
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.7034 pd=24.9 as=0 ps=0 w=12.06 l=2.04
X18 VDD2.t1 VN.t7 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=4.7034 ps=24.9 w=12.06 l=2.04
X19 VDD1.t0 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.9899 pd=12.39 as=4.7034 ps=24.9 w=12.06 l=2.04
R0 VN.n5 VN.t4 175.446
R1 VN.n28 VN.t6 175.446
R2 VN.n43 VN.n23 161.3
R3 VN.n42 VN.n41 161.3
R4 VN.n40 VN.n24 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n25 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n33 VN.n26 161.3
R9 VN.n32 VN.n31 161.3
R10 VN.n30 VN.n27 161.3
R11 VN.n20 VN.n0 161.3
R12 VN.n19 VN.n18 161.3
R13 VN.n17 VN.n1 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n14 VN.n2 161.3
R16 VN.n12 VN.n11 161.3
R17 VN.n10 VN.n3 161.3
R18 VN.n9 VN.n8 161.3
R19 VN.n7 VN.n4 161.3
R20 VN.n6 VN.t1 142.475
R21 VN.n13 VN.t0 142.475
R22 VN.n21 VN.t7 142.475
R23 VN.n29 VN.t5 142.475
R24 VN.n36 VN.t3 142.475
R25 VN.n44 VN.t2 142.475
R26 VN.n22 VN.n21 95.7567
R27 VN.n45 VN.n44 95.7567
R28 VN.n8 VN.n3 56.4773
R29 VN.n31 VN.n26 56.4773
R30 VN.n19 VN.n1 52.0954
R31 VN.n42 VN.n24 52.0954
R32 VN.n6 VN.n5 49.1578
R33 VN.n29 VN.n28 49.1578
R34 VN VN.n45 48.5587
R35 VN.n15 VN.n1 28.7258
R36 VN.n38 VN.n24 28.7258
R37 VN.n8 VN.n7 24.3439
R38 VN.n12 VN.n3 24.3439
R39 VN.n15 VN.n14 24.3439
R40 VN.n20 VN.n19 24.3439
R41 VN.n31 VN.n30 24.3439
R42 VN.n38 VN.n37 24.3439
R43 VN.n35 VN.n26 24.3439
R44 VN.n43 VN.n42 24.3439
R45 VN.n7 VN.n6 21.1793
R46 VN.n13 VN.n12 21.1793
R47 VN.n30 VN.n29 21.1793
R48 VN.n36 VN.n35 21.1793
R49 VN.n21 VN.n20 14.85
R50 VN.n44 VN.n43 14.85
R51 VN.n28 VN.n27 9.46412
R52 VN.n5 VN.n4 9.46412
R53 VN.n14 VN.n13 3.16515
R54 VN.n37 VN.n36 3.16515
R55 VN.n45 VN.n23 0.278398
R56 VN.n22 VN.n0 0.278398
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153422
R74 VDD2.n2 VDD2.n1 61.6823
R75 VDD2.n2 VDD2.n0 61.6823
R76 VDD2 VDD2.n5 61.6795
R77 VDD2.n4 VDD2.n3 60.7163
R78 VDD2.n4 VDD2.n2 43.3058
R79 VDD2.n5 VDD2.t3 1.64229
R80 VDD2.n5 VDD2.t0 1.64229
R81 VDD2.n3 VDD2.t6 1.64229
R82 VDD2.n3 VDD2.t4 1.64229
R83 VDD2.n1 VDD2.t5 1.64229
R84 VDD2.n1 VDD2.t1 1.64229
R85 VDD2.n0 VDD2.t2 1.64229
R86 VDD2.n0 VDD2.t7 1.64229
R87 VDD2 VDD2.n4 1.08024
R88 VTAIL.n530 VTAIL.n470 289.615
R89 VTAIL.n62 VTAIL.n2 289.615
R90 VTAIL.n128 VTAIL.n68 289.615
R91 VTAIL.n196 VTAIL.n136 289.615
R92 VTAIL.n464 VTAIL.n404 289.615
R93 VTAIL.n396 VTAIL.n336 289.615
R94 VTAIL.n330 VTAIL.n270 289.615
R95 VTAIL.n262 VTAIL.n202 289.615
R96 VTAIL.n490 VTAIL.n489 185
R97 VTAIL.n495 VTAIL.n494 185
R98 VTAIL.n497 VTAIL.n496 185
R99 VTAIL.n486 VTAIL.n485 185
R100 VTAIL.n503 VTAIL.n502 185
R101 VTAIL.n505 VTAIL.n504 185
R102 VTAIL.n482 VTAIL.n481 185
R103 VTAIL.n512 VTAIL.n511 185
R104 VTAIL.n513 VTAIL.n480 185
R105 VTAIL.n515 VTAIL.n514 185
R106 VTAIL.n478 VTAIL.n477 185
R107 VTAIL.n521 VTAIL.n520 185
R108 VTAIL.n523 VTAIL.n522 185
R109 VTAIL.n474 VTAIL.n473 185
R110 VTAIL.n529 VTAIL.n528 185
R111 VTAIL.n531 VTAIL.n530 185
R112 VTAIL.n22 VTAIL.n21 185
R113 VTAIL.n27 VTAIL.n26 185
R114 VTAIL.n29 VTAIL.n28 185
R115 VTAIL.n18 VTAIL.n17 185
R116 VTAIL.n35 VTAIL.n34 185
R117 VTAIL.n37 VTAIL.n36 185
R118 VTAIL.n14 VTAIL.n13 185
R119 VTAIL.n44 VTAIL.n43 185
R120 VTAIL.n45 VTAIL.n12 185
R121 VTAIL.n47 VTAIL.n46 185
R122 VTAIL.n10 VTAIL.n9 185
R123 VTAIL.n53 VTAIL.n52 185
R124 VTAIL.n55 VTAIL.n54 185
R125 VTAIL.n6 VTAIL.n5 185
R126 VTAIL.n61 VTAIL.n60 185
R127 VTAIL.n63 VTAIL.n62 185
R128 VTAIL.n88 VTAIL.n87 185
R129 VTAIL.n93 VTAIL.n92 185
R130 VTAIL.n95 VTAIL.n94 185
R131 VTAIL.n84 VTAIL.n83 185
R132 VTAIL.n101 VTAIL.n100 185
R133 VTAIL.n103 VTAIL.n102 185
R134 VTAIL.n80 VTAIL.n79 185
R135 VTAIL.n110 VTAIL.n109 185
R136 VTAIL.n111 VTAIL.n78 185
R137 VTAIL.n113 VTAIL.n112 185
R138 VTAIL.n76 VTAIL.n75 185
R139 VTAIL.n119 VTAIL.n118 185
R140 VTAIL.n121 VTAIL.n120 185
R141 VTAIL.n72 VTAIL.n71 185
R142 VTAIL.n127 VTAIL.n126 185
R143 VTAIL.n129 VTAIL.n128 185
R144 VTAIL.n156 VTAIL.n155 185
R145 VTAIL.n161 VTAIL.n160 185
R146 VTAIL.n163 VTAIL.n162 185
R147 VTAIL.n152 VTAIL.n151 185
R148 VTAIL.n169 VTAIL.n168 185
R149 VTAIL.n171 VTAIL.n170 185
R150 VTAIL.n148 VTAIL.n147 185
R151 VTAIL.n178 VTAIL.n177 185
R152 VTAIL.n179 VTAIL.n146 185
R153 VTAIL.n181 VTAIL.n180 185
R154 VTAIL.n144 VTAIL.n143 185
R155 VTAIL.n187 VTAIL.n186 185
R156 VTAIL.n189 VTAIL.n188 185
R157 VTAIL.n140 VTAIL.n139 185
R158 VTAIL.n195 VTAIL.n194 185
R159 VTAIL.n197 VTAIL.n196 185
R160 VTAIL.n465 VTAIL.n464 185
R161 VTAIL.n463 VTAIL.n462 185
R162 VTAIL.n408 VTAIL.n407 185
R163 VTAIL.n457 VTAIL.n456 185
R164 VTAIL.n455 VTAIL.n454 185
R165 VTAIL.n412 VTAIL.n411 185
R166 VTAIL.n449 VTAIL.n448 185
R167 VTAIL.n447 VTAIL.n414 185
R168 VTAIL.n446 VTAIL.n445 185
R169 VTAIL.n417 VTAIL.n415 185
R170 VTAIL.n440 VTAIL.n439 185
R171 VTAIL.n438 VTAIL.n437 185
R172 VTAIL.n421 VTAIL.n420 185
R173 VTAIL.n432 VTAIL.n431 185
R174 VTAIL.n430 VTAIL.n429 185
R175 VTAIL.n425 VTAIL.n424 185
R176 VTAIL.n397 VTAIL.n396 185
R177 VTAIL.n395 VTAIL.n394 185
R178 VTAIL.n340 VTAIL.n339 185
R179 VTAIL.n389 VTAIL.n388 185
R180 VTAIL.n387 VTAIL.n386 185
R181 VTAIL.n344 VTAIL.n343 185
R182 VTAIL.n381 VTAIL.n380 185
R183 VTAIL.n379 VTAIL.n346 185
R184 VTAIL.n378 VTAIL.n377 185
R185 VTAIL.n349 VTAIL.n347 185
R186 VTAIL.n372 VTAIL.n371 185
R187 VTAIL.n370 VTAIL.n369 185
R188 VTAIL.n353 VTAIL.n352 185
R189 VTAIL.n364 VTAIL.n363 185
R190 VTAIL.n362 VTAIL.n361 185
R191 VTAIL.n357 VTAIL.n356 185
R192 VTAIL.n331 VTAIL.n330 185
R193 VTAIL.n329 VTAIL.n328 185
R194 VTAIL.n274 VTAIL.n273 185
R195 VTAIL.n323 VTAIL.n322 185
R196 VTAIL.n321 VTAIL.n320 185
R197 VTAIL.n278 VTAIL.n277 185
R198 VTAIL.n315 VTAIL.n314 185
R199 VTAIL.n313 VTAIL.n280 185
R200 VTAIL.n312 VTAIL.n311 185
R201 VTAIL.n283 VTAIL.n281 185
R202 VTAIL.n306 VTAIL.n305 185
R203 VTAIL.n304 VTAIL.n303 185
R204 VTAIL.n287 VTAIL.n286 185
R205 VTAIL.n298 VTAIL.n297 185
R206 VTAIL.n296 VTAIL.n295 185
R207 VTAIL.n291 VTAIL.n290 185
R208 VTAIL.n263 VTAIL.n262 185
R209 VTAIL.n261 VTAIL.n260 185
R210 VTAIL.n206 VTAIL.n205 185
R211 VTAIL.n255 VTAIL.n254 185
R212 VTAIL.n253 VTAIL.n252 185
R213 VTAIL.n210 VTAIL.n209 185
R214 VTAIL.n247 VTAIL.n246 185
R215 VTAIL.n245 VTAIL.n212 185
R216 VTAIL.n244 VTAIL.n243 185
R217 VTAIL.n215 VTAIL.n213 185
R218 VTAIL.n238 VTAIL.n237 185
R219 VTAIL.n236 VTAIL.n235 185
R220 VTAIL.n219 VTAIL.n218 185
R221 VTAIL.n230 VTAIL.n229 185
R222 VTAIL.n228 VTAIL.n227 185
R223 VTAIL.n223 VTAIL.n222 185
R224 VTAIL.n491 VTAIL.t8 149.524
R225 VTAIL.n23 VTAIL.t11 149.524
R226 VTAIL.n89 VTAIL.t7 149.524
R227 VTAIL.n157 VTAIL.t6 149.524
R228 VTAIL.n426 VTAIL.t2 149.524
R229 VTAIL.n358 VTAIL.t5 149.524
R230 VTAIL.n292 VTAIL.t9 149.524
R231 VTAIL.n224 VTAIL.t13 149.524
R232 VTAIL.n495 VTAIL.n489 104.615
R233 VTAIL.n496 VTAIL.n495 104.615
R234 VTAIL.n496 VTAIL.n485 104.615
R235 VTAIL.n503 VTAIL.n485 104.615
R236 VTAIL.n504 VTAIL.n503 104.615
R237 VTAIL.n504 VTAIL.n481 104.615
R238 VTAIL.n512 VTAIL.n481 104.615
R239 VTAIL.n513 VTAIL.n512 104.615
R240 VTAIL.n514 VTAIL.n513 104.615
R241 VTAIL.n514 VTAIL.n477 104.615
R242 VTAIL.n521 VTAIL.n477 104.615
R243 VTAIL.n522 VTAIL.n521 104.615
R244 VTAIL.n522 VTAIL.n473 104.615
R245 VTAIL.n529 VTAIL.n473 104.615
R246 VTAIL.n530 VTAIL.n529 104.615
R247 VTAIL.n27 VTAIL.n21 104.615
R248 VTAIL.n28 VTAIL.n27 104.615
R249 VTAIL.n28 VTAIL.n17 104.615
R250 VTAIL.n35 VTAIL.n17 104.615
R251 VTAIL.n36 VTAIL.n35 104.615
R252 VTAIL.n36 VTAIL.n13 104.615
R253 VTAIL.n44 VTAIL.n13 104.615
R254 VTAIL.n45 VTAIL.n44 104.615
R255 VTAIL.n46 VTAIL.n45 104.615
R256 VTAIL.n46 VTAIL.n9 104.615
R257 VTAIL.n53 VTAIL.n9 104.615
R258 VTAIL.n54 VTAIL.n53 104.615
R259 VTAIL.n54 VTAIL.n5 104.615
R260 VTAIL.n61 VTAIL.n5 104.615
R261 VTAIL.n62 VTAIL.n61 104.615
R262 VTAIL.n93 VTAIL.n87 104.615
R263 VTAIL.n94 VTAIL.n93 104.615
R264 VTAIL.n94 VTAIL.n83 104.615
R265 VTAIL.n101 VTAIL.n83 104.615
R266 VTAIL.n102 VTAIL.n101 104.615
R267 VTAIL.n102 VTAIL.n79 104.615
R268 VTAIL.n110 VTAIL.n79 104.615
R269 VTAIL.n111 VTAIL.n110 104.615
R270 VTAIL.n112 VTAIL.n111 104.615
R271 VTAIL.n112 VTAIL.n75 104.615
R272 VTAIL.n119 VTAIL.n75 104.615
R273 VTAIL.n120 VTAIL.n119 104.615
R274 VTAIL.n120 VTAIL.n71 104.615
R275 VTAIL.n127 VTAIL.n71 104.615
R276 VTAIL.n128 VTAIL.n127 104.615
R277 VTAIL.n161 VTAIL.n155 104.615
R278 VTAIL.n162 VTAIL.n161 104.615
R279 VTAIL.n162 VTAIL.n151 104.615
R280 VTAIL.n169 VTAIL.n151 104.615
R281 VTAIL.n170 VTAIL.n169 104.615
R282 VTAIL.n170 VTAIL.n147 104.615
R283 VTAIL.n178 VTAIL.n147 104.615
R284 VTAIL.n179 VTAIL.n178 104.615
R285 VTAIL.n180 VTAIL.n179 104.615
R286 VTAIL.n180 VTAIL.n143 104.615
R287 VTAIL.n187 VTAIL.n143 104.615
R288 VTAIL.n188 VTAIL.n187 104.615
R289 VTAIL.n188 VTAIL.n139 104.615
R290 VTAIL.n195 VTAIL.n139 104.615
R291 VTAIL.n196 VTAIL.n195 104.615
R292 VTAIL.n464 VTAIL.n463 104.615
R293 VTAIL.n463 VTAIL.n407 104.615
R294 VTAIL.n456 VTAIL.n407 104.615
R295 VTAIL.n456 VTAIL.n455 104.615
R296 VTAIL.n455 VTAIL.n411 104.615
R297 VTAIL.n448 VTAIL.n411 104.615
R298 VTAIL.n448 VTAIL.n447 104.615
R299 VTAIL.n447 VTAIL.n446 104.615
R300 VTAIL.n446 VTAIL.n415 104.615
R301 VTAIL.n439 VTAIL.n415 104.615
R302 VTAIL.n439 VTAIL.n438 104.615
R303 VTAIL.n438 VTAIL.n420 104.615
R304 VTAIL.n431 VTAIL.n420 104.615
R305 VTAIL.n431 VTAIL.n430 104.615
R306 VTAIL.n430 VTAIL.n424 104.615
R307 VTAIL.n396 VTAIL.n395 104.615
R308 VTAIL.n395 VTAIL.n339 104.615
R309 VTAIL.n388 VTAIL.n339 104.615
R310 VTAIL.n388 VTAIL.n387 104.615
R311 VTAIL.n387 VTAIL.n343 104.615
R312 VTAIL.n380 VTAIL.n343 104.615
R313 VTAIL.n380 VTAIL.n379 104.615
R314 VTAIL.n379 VTAIL.n378 104.615
R315 VTAIL.n378 VTAIL.n347 104.615
R316 VTAIL.n371 VTAIL.n347 104.615
R317 VTAIL.n371 VTAIL.n370 104.615
R318 VTAIL.n370 VTAIL.n352 104.615
R319 VTAIL.n363 VTAIL.n352 104.615
R320 VTAIL.n363 VTAIL.n362 104.615
R321 VTAIL.n362 VTAIL.n356 104.615
R322 VTAIL.n330 VTAIL.n329 104.615
R323 VTAIL.n329 VTAIL.n273 104.615
R324 VTAIL.n322 VTAIL.n273 104.615
R325 VTAIL.n322 VTAIL.n321 104.615
R326 VTAIL.n321 VTAIL.n277 104.615
R327 VTAIL.n314 VTAIL.n277 104.615
R328 VTAIL.n314 VTAIL.n313 104.615
R329 VTAIL.n313 VTAIL.n312 104.615
R330 VTAIL.n312 VTAIL.n281 104.615
R331 VTAIL.n305 VTAIL.n281 104.615
R332 VTAIL.n305 VTAIL.n304 104.615
R333 VTAIL.n304 VTAIL.n286 104.615
R334 VTAIL.n297 VTAIL.n286 104.615
R335 VTAIL.n297 VTAIL.n296 104.615
R336 VTAIL.n296 VTAIL.n290 104.615
R337 VTAIL.n262 VTAIL.n261 104.615
R338 VTAIL.n261 VTAIL.n205 104.615
R339 VTAIL.n254 VTAIL.n205 104.615
R340 VTAIL.n254 VTAIL.n253 104.615
R341 VTAIL.n253 VTAIL.n209 104.615
R342 VTAIL.n246 VTAIL.n209 104.615
R343 VTAIL.n246 VTAIL.n245 104.615
R344 VTAIL.n245 VTAIL.n244 104.615
R345 VTAIL.n244 VTAIL.n213 104.615
R346 VTAIL.n237 VTAIL.n213 104.615
R347 VTAIL.n237 VTAIL.n236 104.615
R348 VTAIL.n236 VTAIL.n218 104.615
R349 VTAIL.n229 VTAIL.n218 104.615
R350 VTAIL.n229 VTAIL.n228 104.615
R351 VTAIL.n228 VTAIL.n222 104.615
R352 VTAIL.t8 VTAIL.n489 52.3082
R353 VTAIL.t11 VTAIL.n21 52.3082
R354 VTAIL.t7 VTAIL.n87 52.3082
R355 VTAIL.t6 VTAIL.n155 52.3082
R356 VTAIL.t2 VTAIL.n424 52.3082
R357 VTAIL.t5 VTAIL.n356 52.3082
R358 VTAIL.t9 VTAIL.n290 52.3082
R359 VTAIL.t13 VTAIL.n222 52.3082
R360 VTAIL.n403 VTAIL.n402 44.0375
R361 VTAIL.n269 VTAIL.n268 44.0375
R362 VTAIL.n1 VTAIL.n0 44.0373
R363 VTAIL.n135 VTAIL.n134 44.0373
R364 VTAIL.n535 VTAIL.n534 31.0217
R365 VTAIL.n67 VTAIL.n66 31.0217
R366 VTAIL.n133 VTAIL.n132 31.0217
R367 VTAIL.n201 VTAIL.n200 31.0217
R368 VTAIL.n469 VTAIL.n468 31.0217
R369 VTAIL.n401 VTAIL.n400 31.0217
R370 VTAIL.n335 VTAIL.n334 31.0217
R371 VTAIL.n267 VTAIL.n266 31.0217
R372 VTAIL.n535 VTAIL.n469 24.8065
R373 VTAIL.n267 VTAIL.n201 24.8065
R374 VTAIL.n515 VTAIL.n480 13.1884
R375 VTAIL.n47 VTAIL.n12 13.1884
R376 VTAIL.n113 VTAIL.n78 13.1884
R377 VTAIL.n181 VTAIL.n146 13.1884
R378 VTAIL.n449 VTAIL.n414 13.1884
R379 VTAIL.n381 VTAIL.n346 13.1884
R380 VTAIL.n315 VTAIL.n280 13.1884
R381 VTAIL.n247 VTAIL.n212 13.1884
R382 VTAIL.n511 VTAIL.n510 12.8005
R383 VTAIL.n516 VTAIL.n478 12.8005
R384 VTAIL.n43 VTAIL.n42 12.8005
R385 VTAIL.n48 VTAIL.n10 12.8005
R386 VTAIL.n109 VTAIL.n108 12.8005
R387 VTAIL.n114 VTAIL.n76 12.8005
R388 VTAIL.n177 VTAIL.n176 12.8005
R389 VTAIL.n182 VTAIL.n144 12.8005
R390 VTAIL.n450 VTAIL.n412 12.8005
R391 VTAIL.n445 VTAIL.n416 12.8005
R392 VTAIL.n382 VTAIL.n344 12.8005
R393 VTAIL.n377 VTAIL.n348 12.8005
R394 VTAIL.n316 VTAIL.n278 12.8005
R395 VTAIL.n311 VTAIL.n282 12.8005
R396 VTAIL.n248 VTAIL.n210 12.8005
R397 VTAIL.n243 VTAIL.n214 12.8005
R398 VTAIL.n509 VTAIL.n482 12.0247
R399 VTAIL.n520 VTAIL.n519 12.0247
R400 VTAIL.n41 VTAIL.n14 12.0247
R401 VTAIL.n52 VTAIL.n51 12.0247
R402 VTAIL.n107 VTAIL.n80 12.0247
R403 VTAIL.n118 VTAIL.n117 12.0247
R404 VTAIL.n175 VTAIL.n148 12.0247
R405 VTAIL.n186 VTAIL.n185 12.0247
R406 VTAIL.n454 VTAIL.n453 12.0247
R407 VTAIL.n444 VTAIL.n417 12.0247
R408 VTAIL.n386 VTAIL.n385 12.0247
R409 VTAIL.n376 VTAIL.n349 12.0247
R410 VTAIL.n320 VTAIL.n319 12.0247
R411 VTAIL.n310 VTAIL.n283 12.0247
R412 VTAIL.n252 VTAIL.n251 12.0247
R413 VTAIL.n242 VTAIL.n215 12.0247
R414 VTAIL.n506 VTAIL.n505 11.249
R415 VTAIL.n523 VTAIL.n476 11.249
R416 VTAIL.n38 VTAIL.n37 11.249
R417 VTAIL.n55 VTAIL.n8 11.249
R418 VTAIL.n104 VTAIL.n103 11.249
R419 VTAIL.n121 VTAIL.n74 11.249
R420 VTAIL.n172 VTAIL.n171 11.249
R421 VTAIL.n189 VTAIL.n142 11.249
R422 VTAIL.n457 VTAIL.n410 11.249
R423 VTAIL.n441 VTAIL.n440 11.249
R424 VTAIL.n389 VTAIL.n342 11.249
R425 VTAIL.n373 VTAIL.n372 11.249
R426 VTAIL.n323 VTAIL.n276 11.249
R427 VTAIL.n307 VTAIL.n306 11.249
R428 VTAIL.n255 VTAIL.n208 11.249
R429 VTAIL.n239 VTAIL.n238 11.249
R430 VTAIL.n502 VTAIL.n484 10.4732
R431 VTAIL.n524 VTAIL.n474 10.4732
R432 VTAIL.n34 VTAIL.n16 10.4732
R433 VTAIL.n56 VTAIL.n6 10.4732
R434 VTAIL.n100 VTAIL.n82 10.4732
R435 VTAIL.n122 VTAIL.n72 10.4732
R436 VTAIL.n168 VTAIL.n150 10.4732
R437 VTAIL.n190 VTAIL.n140 10.4732
R438 VTAIL.n458 VTAIL.n408 10.4732
R439 VTAIL.n437 VTAIL.n419 10.4732
R440 VTAIL.n390 VTAIL.n340 10.4732
R441 VTAIL.n369 VTAIL.n351 10.4732
R442 VTAIL.n324 VTAIL.n274 10.4732
R443 VTAIL.n303 VTAIL.n285 10.4732
R444 VTAIL.n256 VTAIL.n206 10.4732
R445 VTAIL.n235 VTAIL.n217 10.4732
R446 VTAIL.n491 VTAIL.n490 10.2747
R447 VTAIL.n23 VTAIL.n22 10.2747
R448 VTAIL.n89 VTAIL.n88 10.2747
R449 VTAIL.n157 VTAIL.n156 10.2747
R450 VTAIL.n426 VTAIL.n425 10.2747
R451 VTAIL.n358 VTAIL.n357 10.2747
R452 VTAIL.n292 VTAIL.n291 10.2747
R453 VTAIL.n224 VTAIL.n223 10.2747
R454 VTAIL.n501 VTAIL.n486 9.69747
R455 VTAIL.n528 VTAIL.n527 9.69747
R456 VTAIL.n33 VTAIL.n18 9.69747
R457 VTAIL.n60 VTAIL.n59 9.69747
R458 VTAIL.n99 VTAIL.n84 9.69747
R459 VTAIL.n126 VTAIL.n125 9.69747
R460 VTAIL.n167 VTAIL.n152 9.69747
R461 VTAIL.n194 VTAIL.n193 9.69747
R462 VTAIL.n462 VTAIL.n461 9.69747
R463 VTAIL.n436 VTAIL.n421 9.69747
R464 VTAIL.n394 VTAIL.n393 9.69747
R465 VTAIL.n368 VTAIL.n353 9.69747
R466 VTAIL.n328 VTAIL.n327 9.69747
R467 VTAIL.n302 VTAIL.n287 9.69747
R468 VTAIL.n260 VTAIL.n259 9.69747
R469 VTAIL.n234 VTAIL.n219 9.69747
R470 VTAIL.n534 VTAIL.n533 9.45567
R471 VTAIL.n66 VTAIL.n65 9.45567
R472 VTAIL.n132 VTAIL.n131 9.45567
R473 VTAIL.n200 VTAIL.n199 9.45567
R474 VTAIL.n468 VTAIL.n467 9.45567
R475 VTAIL.n400 VTAIL.n399 9.45567
R476 VTAIL.n334 VTAIL.n333 9.45567
R477 VTAIL.n266 VTAIL.n265 9.45567
R478 VTAIL.n533 VTAIL.n532 9.3005
R479 VTAIL.n472 VTAIL.n471 9.3005
R480 VTAIL.n527 VTAIL.n526 9.3005
R481 VTAIL.n525 VTAIL.n524 9.3005
R482 VTAIL.n476 VTAIL.n475 9.3005
R483 VTAIL.n519 VTAIL.n518 9.3005
R484 VTAIL.n517 VTAIL.n516 9.3005
R485 VTAIL.n493 VTAIL.n492 9.3005
R486 VTAIL.n488 VTAIL.n487 9.3005
R487 VTAIL.n499 VTAIL.n498 9.3005
R488 VTAIL.n501 VTAIL.n500 9.3005
R489 VTAIL.n484 VTAIL.n483 9.3005
R490 VTAIL.n507 VTAIL.n506 9.3005
R491 VTAIL.n509 VTAIL.n508 9.3005
R492 VTAIL.n510 VTAIL.n479 9.3005
R493 VTAIL.n65 VTAIL.n64 9.3005
R494 VTAIL.n4 VTAIL.n3 9.3005
R495 VTAIL.n59 VTAIL.n58 9.3005
R496 VTAIL.n57 VTAIL.n56 9.3005
R497 VTAIL.n8 VTAIL.n7 9.3005
R498 VTAIL.n51 VTAIL.n50 9.3005
R499 VTAIL.n49 VTAIL.n48 9.3005
R500 VTAIL.n25 VTAIL.n24 9.3005
R501 VTAIL.n20 VTAIL.n19 9.3005
R502 VTAIL.n31 VTAIL.n30 9.3005
R503 VTAIL.n33 VTAIL.n32 9.3005
R504 VTAIL.n16 VTAIL.n15 9.3005
R505 VTAIL.n39 VTAIL.n38 9.3005
R506 VTAIL.n41 VTAIL.n40 9.3005
R507 VTAIL.n42 VTAIL.n11 9.3005
R508 VTAIL.n131 VTAIL.n130 9.3005
R509 VTAIL.n70 VTAIL.n69 9.3005
R510 VTAIL.n125 VTAIL.n124 9.3005
R511 VTAIL.n123 VTAIL.n122 9.3005
R512 VTAIL.n74 VTAIL.n73 9.3005
R513 VTAIL.n117 VTAIL.n116 9.3005
R514 VTAIL.n115 VTAIL.n114 9.3005
R515 VTAIL.n91 VTAIL.n90 9.3005
R516 VTAIL.n86 VTAIL.n85 9.3005
R517 VTAIL.n97 VTAIL.n96 9.3005
R518 VTAIL.n99 VTAIL.n98 9.3005
R519 VTAIL.n82 VTAIL.n81 9.3005
R520 VTAIL.n105 VTAIL.n104 9.3005
R521 VTAIL.n107 VTAIL.n106 9.3005
R522 VTAIL.n108 VTAIL.n77 9.3005
R523 VTAIL.n199 VTAIL.n198 9.3005
R524 VTAIL.n138 VTAIL.n137 9.3005
R525 VTAIL.n193 VTAIL.n192 9.3005
R526 VTAIL.n191 VTAIL.n190 9.3005
R527 VTAIL.n142 VTAIL.n141 9.3005
R528 VTAIL.n185 VTAIL.n184 9.3005
R529 VTAIL.n183 VTAIL.n182 9.3005
R530 VTAIL.n159 VTAIL.n158 9.3005
R531 VTAIL.n154 VTAIL.n153 9.3005
R532 VTAIL.n165 VTAIL.n164 9.3005
R533 VTAIL.n167 VTAIL.n166 9.3005
R534 VTAIL.n150 VTAIL.n149 9.3005
R535 VTAIL.n173 VTAIL.n172 9.3005
R536 VTAIL.n175 VTAIL.n174 9.3005
R537 VTAIL.n176 VTAIL.n145 9.3005
R538 VTAIL.n428 VTAIL.n427 9.3005
R539 VTAIL.n423 VTAIL.n422 9.3005
R540 VTAIL.n434 VTAIL.n433 9.3005
R541 VTAIL.n436 VTAIL.n435 9.3005
R542 VTAIL.n419 VTAIL.n418 9.3005
R543 VTAIL.n442 VTAIL.n441 9.3005
R544 VTAIL.n444 VTAIL.n443 9.3005
R545 VTAIL.n416 VTAIL.n413 9.3005
R546 VTAIL.n467 VTAIL.n466 9.3005
R547 VTAIL.n406 VTAIL.n405 9.3005
R548 VTAIL.n461 VTAIL.n460 9.3005
R549 VTAIL.n459 VTAIL.n458 9.3005
R550 VTAIL.n410 VTAIL.n409 9.3005
R551 VTAIL.n453 VTAIL.n452 9.3005
R552 VTAIL.n451 VTAIL.n450 9.3005
R553 VTAIL.n360 VTAIL.n359 9.3005
R554 VTAIL.n355 VTAIL.n354 9.3005
R555 VTAIL.n366 VTAIL.n365 9.3005
R556 VTAIL.n368 VTAIL.n367 9.3005
R557 VTAIL.n351 VTAIL.n350 9.3005
R558 VTAIL.n374 VTAIL.n373 9.3005
R559 VTAIL.n376 VTAIL.n375 9.3005
R560 VTAIL.n348 VTAIL.n345 9.3005
R561 VTAIL.n399 VTAIL.n398 9.3005
R562 VTAIL.n338 VTAIL.n337 9.3005
R563 VTAIL.n393 VTAIL.n392 9.3005
R564 VTAIL.n391 VTAIL.n390 9.3005
R565 VTAIL.n342 VTAIL.n341 9.3005
R566 VTAIL.n385 VTAIL.n384 9.3005
R567 VTAIL.n383 VTAIL.n382 9.3005
R568 VTAIL.n294 VTAIL.n293 9.3005
R569 VTAIL.n289 VTAIL.n288 9.3005
R570 VTAIL.n300 VTAIL.n299 9.3005
R571 VTAIL.n302 VTAIL.n301 9.3005
R572 VTAIL.n285 VTAIL.n284 9.3005
R573 VTAIL.n308 VTAIL.n307 9.3005
R574 VTAIL.n310 VTAIL.n309 9.3005
R575 VTAIL.n282 VTAIL.n279 9.3005
R576 VTAIL.n333 VTAIL.n332 9.3005
R577 VTAIL.n272 VTAIL.n271 9.3005
R578 VTAIL.n327 VTAIL.n326 9.3005
R579 VTAIL.n325 VTAIL.n324 9.3005
R580 VTAIL.n276 VTAIL.n275 9.3005
R581 VTAIL.n319 VTAIL.n318 9.3005
R582 VTAIL.n317 VTAIL.n316 9.3005
R583 VTAIL.n226 VTAIL.n225 9.3005
R584 VTAIL.n221 VTAIL.n220 9.3005
R585 VTAIL.n232 VTAIL.n231 9.3005
R586 VTAIL.n234 VTAIL.n233 9.3005
R587 VTAIL.n217 VTAIL.n216 9.3005
R588 VTAIL.n240 VTAIL.n239 9.3005
R589 VTAIL.n242 VTAIL.n241 9.3005
R590 VTAIL.n214 VTAIL.n211 9.3005
R591 VTAIL.n265 VTAIL.n264 9.3005
R592 VTAIL.n204 VTAIL.n203 9.3005
R593 VTAIL.n259 VTAIL.n258 9.3005
R594 VTAIL.n257 VTAIL.n256 9.3005
R595 VTAIL.n208 VTAIL.n207 9.3005
R596 VTAIL.n251 VTAIL.n250 9.3005
R597 VTAIL.n249 VTAIL.n248 9.3005
R598 VTAIL.n498 VTAIL.n497 8.92171
R599 VTAIL.n531 VTAIL.n472 8.92171
R600 VTAIL.n30 VTAIL.n29 8.92171
R601 VTAIL.n63 VTAIL.n4 8.92171
R602 VTAIL.n96 VTAIL.n95 8.92171
R603 VTAIL.n129 VTAIL.n70 8.92171
R604 VTAIL.n164 VTAIL.n163 8.92171
R605 VTAIL.n197 VTAIL.n138 8.92171
R606 VTAIL.n465 VTAIL.n406 8.92171
R607 VTAIL.n433 VTAIL.n432 8.92171
R608 VTAIL.n397 VTAIL.n338 8.92171
R609 VTAIL.n365 VTAIL.n364 8.92171
R610 VTAIL.n331 VTAIL.n272 8.92171
R611 VTAIL.n299 VTAIL.n298 8.92171
R612 VTAIL.n263 VTAIL.n204 8.92171
R613 VTAIL.n231 VTAIL.n230 8.92171
R614 VTAIL.n494 VTAIL.n488 8.14595
R615 VTAIL.n532 VTAIL.n470 8.14595
R616 VTAIL.n26 VTAIL.n20 8.14595
R617 VTAIL.n64 VTAIL.n2 8.14595
R618 VTAIL.n92 VTAIL.n86 8.14595
R619 VTAIL.n130 VTAIL.n68 8.14595
R620 VTAIL.n160 VTAIL.n154 8.14595
R621 VTAIL.n198 VTAIL.n136 8.14595
R622 VTAIL.n466 VTAIL.n404 8.14595
R623 VTAIL.n429 VTAIL.n423 8.14595
R624 VTAIL.n398 VTAIL.n336 8.14595
R625 VTAIL.n361 VTAIL.n355 8.14595
R626 VTAIL.n332 VTAIL.n270 8.14595
R627 VTAIL.n295 VTAIL.n289 8.14595
R628 VTAIL.n264 VTAIL.n202 8.14595
R629 VTAIL.n227 VTAIL.n221 8.14595
R630 VTAIL.n493 VTAIL.n490 7.3702
R631 VTAIL.n25 VTAIL.n22 7.3702
R632 VTAIL.n91 VTAIL.n88 7.3702
R633 VTAIL.n159 VTAIL.n156 7.3702
R634 VTAIL.n428 VTAIL.n425 7.3702
R635 VTAIL.n360 VTAIL.n357 7.3702
R636 VTAIL.n294 VTAIL.n291 7.3702
R637 VTAIL.n226 VTAIL.n223 7.3702
R638 VTAIL.n494 VTAIL.n493 5.81868
R639 VTAIL.n534 VTAIL.n470 5.81868
R640 VTAIL.n26 VTAIL.n25 5.81868
R641 VTAIL.n66 VTAIL.n2 5.81868
R642 VTAIL.n92 VTAIL.n91 5.81868
R643 VTAIL.n132 VTAIL.n68 5.81868
R644 VTAIL.n160 VTAIL.n159 5.81868
R645 VTAIL.n200 VTAIL.n136 5.81868
R646 VTAIL.n468 VTAIL.n404 5.81868
R647 VTAIL.n429 VTAIL.n428 5.81868
R648 VTAIL.n400 VTAIL.n336 5.81868
R649 VTAIL.n361 VTAIL.n360 5.81868
R650 VTAIL.n334 VTAIL.n270 5.81868
R651 VTAIL.n295 VTAIL.n294 5.81868
R652 VTAIL.n266 VTAIL.n202 5.81868
R653 VTAIL.n227 VTAIL.n226 5.81868
R654 VTAIL.n497 VTAIL.n488 5.04292
R655 VTAIL.n532 VTAIL.n531 5.04292
R656 VTAIL.n29 VTAIL.n20 5.04292
R657 VTAIL.n64 VTAIL.n63 5.04292
R658 VTAIL.n95 VTAIL.n86 5.04292
R659 VTAIL.n130 VTAIL.n129 5.04292
R660 VTAIL.n163 VTAIL.n154 5.04292
R661 VTAIL.n198 VTAIL.n197 5.04292
R662 VTAIL.n466 VTAIL.n465 5.04292
R663 VTAIL.n432 VTAIL.n423 5.04292
R664 VTAIL.n398 VTAIL.n397 5.04292
R665 VTAIL.n364 VTAIL.n355 5.04292
R666 VTAIL.n332 VTAIL.n331 5.04292
R667 VTAIL.n298 VTAIL.n289 5.04292
R668 VTAIL.n264 VTAIL.n263 5.04292
R669 VTAIL.n230 VTAIL.n221 5.04292
R670 VTAIL.n498 VTAIL.n486 4.26717
R671 VTAIL.n528 VTAIL.n472 4.26717
R672 VTAIL.n30 VTAIL.n18 4.26717
R673 VTAIL.n60 VTAIL.n4 4.26717
R674 VTAIL.n96 VTAIL.n84 4.26717
R675 VTAIL.n126 VTAIL.n70 4.26717
R676 VTAIL.n164 VTAIL.n152 4.26717
R677 VTAIL.n194 VTAIL.n138 4.26717
R678 VTAIL.n462 VTAIL.n406 4.26717
R679 VTAIL.n433 VTAIL.n421 4.26717
R680 VTAIL.n394 VTAIL.n338 4.26717
R681 VTAIL.n365 VTAIL.n353 4.26717
R682 VTAIL.n328 VTAIL.n272 4.26717
R683 VTAIL.n299 VTAIL.n287 4.26717
R684 VTAIL.n260 VTAIL.n204 4.26717
R685 VTAIL.n231 VTAIL.n219 4.26717
R686 VTAIL.n502 VTAIL.n501 3.49141
R687 VTAIL.n527 VTAIL.n474 3.49141
R688 VTAIL.n34 VTAIL.n33 3.49141
R689 VTAIL.n59 VTAIL.n6 3.49141
R690 VTAIL.n100 VTAIL.n99 3.49141
R691 VTAIL.n125 VTAIL.n72 3.49141
R692 VTAIL.n168 VTAIL.n167 3.49141
R693 VTAIL.n193 VTAIL.n140 3.49141
R694 VTAIL.n461 VTAIL.n408 3.49141
R695 VTAIL.n437 VTAIL.n436 3.49141
R696 VTAIL.n393 VTAIL.n340 3.49141
R697 VTAIL.n369 VTAIL.n368 3.49141
R698 VTAIL.n327 VTAIL.n274 3.49141
R699 VTAIL.n303 VTAIL.n302 3.49141
R700 VTAIL.n259 VTAIL.n206 3.49141
R701 VTAIL.n235 VTAIL.n234 3.49141
R702 VTAIL.n492 VTAIL.n491 2.84303
R703 VTAIL.n24 VTAIL.n23 2.84303
R704 VTAIL.n90 VTAIL.n89 2.84303
R705 VTAIL.n158 VTAIL.n157 2.84303
R706 VTAIL.n427 VTAIL.n426 2.84303
R707 VTAIL.n359 VTAIL.n358 2.84303
R708 VTAIL.n293 VTAIL.n292 2.84303
R709 VTAIL.n225 VTAIL.n224 2.84303
R710 VTAIL.n505 VTAIL.n484 2.71565
R711 VTAIL.n524 VTAIL.n523 2.71565
R712 VTAIL.n37 VTAIL.n16 2.71565
R713 VTAIL.n56 VTAIL.n55 2.71565
R714 VTAIL.n103 VTAIL.n82 2.71565
R715 VTAIL.n122 VTAIL.n121 2.71565
R716 VTAIL.n171 VTAIL.n150 2.71565
R717 VTAIL.n190 VTAIL.n189 2.71565
R718 VTAIL.n458 VTAIL.n457 2.71565
R719 VTAIL.n440 VTAIL.n419 2.71565
R720 VTAIL.n390 VTAIL.n389 2.71565
R721 VTAIL.n372 VTAIL.n351 2.71565
R722 VTAIL.n324 VTAIL.n323 2.71565
R723 VTAIL.n306 VTAIL.n285 2.71565
R724 VTAIL.n256 VTAIL.n255 2.71565
R725 VTAIL.n238 VTAIL.n217 2.71565
R726 VTAIL.n269 VTAIL.n267 2.0436
R727 VTAIL.n335 VTAIL.n269 2.0436
R728 VTAIL.n403 VTAIL.n401 2.0436
R729 VTAIL.n469 VTAIL.n403 2.0436
R730 VTAIL.n201 VTAIL.n135 2.0436
R731 VTAIL.n135 VTAIL.n133 2.0436
R732 VTAIL.n67 VTAIL.n1 2.0436
R733 VTAIL VTAIL.n535 1.98541
R734 VTAIL.n506 VTAIL.n482 1.93989
R735 VTAIL.n520 VTAIL.n476 1.93989
R736 VTAIL.n38 VTAIL.n14 1.93989
R737 VTAIL.n52 VTAIL.n8 1.93989
R738 VTAIL.n104 VTAIL.n80 1.93989
R739 VTAIL.n118 VTAIL.n74 1.93989
R740 VTAIL.n172 VTAIL.n148 1.93989
R741 VTAIL.n186 VTAIL.n142 1.93989
R742 VTAIL.n454 VTAIL.n410 1.93989
R743 VTAIL.n441 VTAIL.n417 1.93989
R744 VTAIL.n386 VTAIL.n342 1.93989
R745 VTAIL.n373 VTAIL.n349 1.93989
R746 VTAIL.n320 VTAIL.n276 1.93989
R747 VTAIL.n307 VTAIL.n283 1.93989
R748 VTAIL.n252 VTAIL.n208 1.93989
R749 VTAIL.n239 VTAIL.n215 1.93989
R750 VTAIL.n0 VTAIL.t14 1.64229
R751 VTAIL.n0 VTAIL.t15 1.64229
R752 VTAIL.n134 VTAIL.t3 1.64229
R753 VTAIL.n134 VTAIL.t4 1.64229
R754 VTAIL.n402 VTAIL.t1 1.64229
R755 VTAIL.n402 VTAIL.t0 1.64229
R756 VTAIL.n268 VTAIL.t12 1.64229
R757 VTAIL.n268 VTAIL.t10 1.64229
R758 VTAIL.n511 VTAIL.n509 1.16414
R759 VTAIL.n519 VTAIL.n478 1.16414
R760 VTAIL.n43 VTAIL.n41 1.16414
R761 VTAIL.n51 VTAIL.n10 1.16414
R762 VTAIL.n109 VTAIL.n107 1.16414
R763 VTAIL.n117 VTAIL.n76 1.16414
R764 VTAIL.n177 VTAIL.n175 1.16414
R765 VTAIL.n185 VTAIL.n144 1.16414
R766 VTAIL.n453 VTAIL.n412 1.16414
R767 VTAIL.n445 VTAIL.n444 1.16414
R768 VTAIL.n385 VTAIL.n344 1.16414
R769 VTAIL.n377 VTAIL.n376 1.16414
R770 VTAIL.n319 VTAIL.n278 1.16414
R771 VTAIL.n311 VTAIL.n310 1.16414
R772 VTAIL.n251 VTAIL.n210 1.16414
R773 VTAIL.n243 VTAIL.n242 1.16414
R774 VTAIL.n401 VTAIL.n335 0.470328
R775 VTAIL.n133 VTAIL.n67 0.470328
R776 VTAIL.n510 VTAIL.n480 0.388379
R777 VTAIL.n516 VTAIL.n515 0.388379
R778 VTAIL.n42 VTAIL.n12 0.388379
R779 VTAIL.n48 VTAIL.n47 0.388379
R780 VTAIL.n108 VTAIL.n78 0.388379
R781 VTAIL.n114 VTAIL.n113 0.388379
R782 VTAIL.n176 VTAIL.n146 0.388379
R783 VTAIL.n182 VTAIL.n181 0.388379
R784 VTAIL.n450 VTAIL.n449 0.388379
R785 VTAIL.n416 VTAIL.n414 0.388379
R786 VTAIL.n382 VTAIL.n381 0.388379
R787 VTAIL.n348 VTAIL.n346 0.388379
R788 VTAIL.n316 VTAIL.n315 0.388379
R789 VTAIL.n282 VTAIL.n280 0.388379
R790 VTAIL.n248 VTAIL.n247 0.388379
R791 VTAIL.n214 VTAIL.n212 0.388379
R792 VTAIL.n492 VTAIL.n487 0.155672
R793 VTAIL.n499 VTAIL.n487 0.155672
R794 VTAIL.n500 VTAIL.n499 0.155672
R795 VTAIL.n500 VTAIL.n483 0.155672
R796 VTAIL.n507 VTAIL.n483 0.155672
R797 VTAIL.n508 VTAIL.n507 0.155672
R798 VTAIL.n508 VTAIL.n479 0.155672
R799 VTAIL.n517 VTAIL.n479 0.155672
R800 VTAIL.n518 VTAIL.n517 0.155672
R801 VTAIL.n518 VTAIL.n475 0.155672
R802 VTAIL.n525 VTAIL.n475 0.155672
R803 VTAIL.n526 VTAIL.n525 0.155672
R804 VTAIL.n526 VTAIL.n471 0.155672
R805 VTAIL.n533 VTAIL.n471 0.155672
R806 VTAIL.n24 VTAIL.n19 0.155672
R807 VTAIL.n31 VTAIL.n19 0.155672
R808 VTAIL.n32 VTAIL.n31 0.155672
R809 VTAIL.n32 VTAIL.n15 0.155672
R810 VTAIL.n39 VTAIL.n15 0.155672
R811 VTAIL.n40 VTAIL.n39 0.155672
R812 VTAIL.n40 VTAIL.n11 0.155672
R813 VTAIL.n49 VTAIL.n11 0.155672
R814 VTAIL.n50 VTAIL.n49 0.155672
R815 VTAIL.n50 VTAIL.n7 0.155672
R816 VTAIL.n57 VTAIL.n7 0.155672
R817 VTAIL.n58 VTAIL.n57 0.155672
R818 VTAIL.n58 VTAIL.n3 0.155672
R819 VTAIL.n65 VTAIL.n3 0.155672
R820 VTAIL.n90 VTAIL.n85 0.155672
R821 VTAIL.n97 VTAIL.n85 0.155672
R822 VTAIL.n98 VTAIL.n97 0.155672
R823 VTAIL.n98 VTAIL.n81 0.155672
R824 VTAIL.n105 VTAIL.n81 0.155672
R825 VTAIL.n106 VTAIL.n105 0.155672
R826 VTAIL.n106 VTAIL.n77 0.155672
R827 VTAIL.n115 VTAIL.n77 0.155672
R828 VTAIL.n116 VTAIL.n115 0.155672
R829 VTAIL.n116 VTAIL.n73 0.155672
R830 VTAIL.n123 VTAIL.n73 0.155672
R831 VTAIL.n124 VTAIL.n123 0.155672
R832 VTAIL.n124 VTAIL.n69 0.155672
R833 VTAIL.n131 VTAIL.n69 0.155672
R834 VTAIL.n158 VTAIL.n153 0.155672
R835 VTAIL.n165 VTAIL.n153 0.155672
R836 VTAIL.n166 VTAIL.n165 0.155672
R837 VTAIL.n166 VTAIL.n149 0.155672
R838 VTAIL.n173 VTAIL.n149 0.155672
R839 VTAIL.n174 VTAIL.n173 0.155672
R840 VTAIL.n174 VTAIL.n145 0.155672
R841 VTAIL.n183 VTAIL.n145 0.155672
R842 VTAIL.n184 VTAIL.n183 0.155672
R843 VTAIL.n184 VTAIL.n141 0.155672
R844 VTAIL.n191 VTAIL.n141 0.155672
R845 VTAIL.n192 VTAIL.n191 0.155672
R846 VTAIL.n192 VTAIL.n137 0.155672
R847 VTAIL.n199 VTAIL.n137 0.155672
R848 VTAIL.n467 VTAIL.n405 0.155672
R849 VTAIL.n460 VTAIL.n405 0.155672
R850 VTAIL.n460 VTAIL.n459 0.155672
R851 VTAIL.n459 VTAIL.n409 0.155672
R852 VTAIL.n452 VTAIL.n409 0.155672
R853 VTAIL.n452 VTAIL.n451 0.155672
R854 VTAIL.n451 VTAIL.n413 0.155672
R855 VTAIL.n443 VTAIL.n413 0.155672
R856 VTAIL.n443 VTAIL.n442 0.155672
R857 VTAIL.n442 VTAIL.n418 0.155672
R858 VTAIL.n435 VTAIL.n418 0.155672
R859 VTAIL.n435 VTAIL.n434 0.155672
R860 VTAIL.n434 VTAIL.n422 0.155672
R861 VTAIL.n427 VTAIL.n422 0.155672
R862 VTAIL.n399 VTAIL.n337 0.155672
R863 VTAIL.n392 VTAIL.n337 0.155672
R864 VTAIL.n392 VTAIL.n391 0.155672
R865 VTAIL.n391 VTAIL.n341 0.155672
R866 VTAIL.n384 VTAIL.n341 0.155672
R867 VTAIL.n384 VTAIL.n383 0.155672
R868 VTAIL.n383 VTAIL.n345 0.155672
R869 VTAIL.n375 VTAIL.n345 0.155672
R870 VTAIL.n375 VTAIL.n374 0.155672
R871 VTAIL.n374 VTAIL.n350 0.155672
R872 VTAIL.n367 VTAIL.n350 0.155672
R873 VTAIL.n367 VTAIL.n366 0.155672
R874 VTAIL.n366 VTAIL.n354 0.155672
R875 VTAIL.n359 VTAIL.n354 0.155672
R876 VTAIL.n333 VTAIL.n271 0.155672
R877 VTAIL.n326 VTAIL.n271 0.155672
R878 VTAIL.n326 VTAIL.n325 0.155672
R879 VTAIL.n325 VTAIL.n275 0.155672
R880 VTAIL.n318 VTAIL.n275 0.155672
R881 VTAIL.n318 VTAIL.n317 0.155672
R882 VTAIL.n317 VTAIL.n279 0.155672
R883 VTAIL.n309 VTAIL.n279 0.155672
R884 VTAIL.n309 VTAIL.n308 0.155672
R885 VTAIL.n308 VTAIL.n284 0.155672
R886 VTAIL.n301 VTAIL.n284 0.155672
R887 VTAIL.n301 VTAIL.n300 0.155672
R888 VTAIL.n300 VTAIL.n288 0.155672
R889 VTAIL.n293 VTAIL.n288 0.155672
R890 VTAIL.n265 VTAIL.n203 0.155672
R891 VTAIL.n258 VTAIL.n203 0.155672
R892 VTAIL.n258 VTAIL.n257 0.155672
R893 VTAIL.n257 VTAIL.n207 0.155672
R894 VTAIL.n250 VTAIL.n207 0.155672
R895 VTAIL.n250 VTAIL.n249 0.155672
R896 VTAIL.n249 VTAIL.n211 0.155672
R897 VTAIL.n241 VTAIL.n211 0.155672
R898 VTAIL.n241 VTAIL.n240 0.155672
R899 VTAIL.n240 VTAIL.n216 0.155672
R900 VTAIL.n233 VTAIL.n216 0.155672
R901 VTAIL.n233 VTAIL.n232 0.155672
R902 VTAIL.n232 VTAIL.n220 0.155672
R903 VTAIL.n225 VTAIL.n220 0.155672
R904 VTAIL VTAIL.n1 0.0586897
R905 B.n819 B.n818 585
R906 B.n820 B.n819 585
R907 B.n313 B.n127 585
R908 B.n312 B.n311 585
R909 B.n310 B.n309 585
R910 B.n308 B.n307 585
R911 B.n306 B.n305 585
R912 B.n304 B.n303 585
R913 B.n302 B.n301 585
R914 B.n300 B.n299 585
R915 B.n298 B.n297 585
R916 B.n296 B.n295 585
R917 B.n294 B.n293 585
R918 B.n292 B.n291 585
R919 B.n290 B.n289 585
R920 B.n288 B.n287 585
R921 B.n286 B.n285 585
R922 B.n284 B.n283 585
R923 B.n282 B.n281 585
R924 B.n280 B.n279 585
R925 B.n278 B.n277 585
R926 B.n276 B.n275 585
R927 B.n274 B.n273 585
R928 B.n272 B.n271 585
R929 B.n270 B.n269 585
R930 B.n268 B.n267 585
R931 B.n266 B.n265 585
R932 B.n264 B.n263 585
R933 B.n262 B.n261 585
R934 B.n260 B.n259 585
R935 B.n258 B.n257 585
R936 B.n256 B.n255 585
R937 B.n254 B.n253 585
R938 B.n252 B.n251 585
R939 B.n250 B.n249 585
R940 B.n248 B.n247 585
R941 B.n246 B.n245 585
R942 B.n244 B.n243 585
R943 B.n242 B.n241 585
R944 B.n240 B.n239 585
R945 B.n238 B.n237 585
R946 B.n236 B.n235 585
R947 B.n234 B.n233 585
R948 B.n231 B.n230 585
R949 B.n229 B.n228 585
R950 B.n227 B.n226 585
R951 B.n225 B.n224 585
R952 B.n223 B.n222 585
R953 B.n221 B.n220 585
R954 B.n219 B.n218 585
R955 B.n217 B.n216 585
R956 B.n215 B.n214 585
R957 B.n213 B.n212 585
R958 B.n211 B.n210 585
R959 B.n209 B.n208 585
R960 B.n207 B.n206 585
R961 B.n205 B.n204 585
R962 B.n203 B.n202 585
R963 B.n201 B.n200 585
R964 B.n199 B.n198 585
R965 B.n197 B.n196 585
R966 B.n195 B.n194 585
R967 B.n193 B.n192 585
R968 B.n191 B.n190 585
R969 B.n189 B.n188 585
R970 B.n187 B.n186 585
R971 B.n185 B.n184 585
R972 B.n183 B.n182 585
R973 B.n181 B.n180 585
R974 B.n179 B.n178 585
R975 B.n177 B.n176 585
R976 B.n175 B.n174 585
R977 B.n173 B.n172 585
R978 B.n171 B.n170 585
R979 B.n169 B.n168 585
R980 B.n167 B.n166 585
R981 B.n165 B.n164 585
R982 B.n163 B.n162 585
R983 B.n161 B.n160 585
R984 B.n159 B.n158 585
R985 B.n157 B.n156 585
R986 B.n155 B.n154 585
R987 B.n153 B.n152 585
R988 B.n151 B.n150 585
R989 B.n149 B.n148 585
R990 B.n147 B.n146 585
R991 B.n145 B.n144 585
R992 B.n143 B.n142 585
R993 B.n141 B.n140 585
R994 B.n139 B.n138 585
R995 B.n137 B.n136 585
R996 B.n135 B.n134 585
R997 B.n81 B.n80 585
R998 B.n823 B.n822 585
R999 B.n817 B.n128 585
R1000 B.n128 B.n78 585
R1001 B.n816 B.n77 585
R1002 B.n827 B.n77 585
R1003 B.n815 B.n76 585
R1004 B.n828 B.n76 585
R1005 B.n814 B.n75 585
R1006 B.n829 B.n75 585
R1007 B.n813 B.n812 585
R1008 B.n812 B.n71 585
R1009 B.n811 B.n70 585
R1010 B.n835 B.n70 585
R1011 B.n810 B.n69 585
R1012 B.n836 B.n69 585
R1013 B.n809 B.n68 585
R1014 B.n837 B.n68 585
R1015 B.n808 B.n807 585
R1016 B.n807 B.n64 585
R1017 B.n806 B.n63 585
R1018 B.n843 B.n63 585
R1019 B.n805 B.n62 585
R1020 B.n844 B.n62 585
R1021 B.n804 B.n61 585
R1022 B.n845 B.n61 585
R1023 B.n803 B.n802 585
R1024 B.n802 B.n57 585
R1025 B.n801 B.n56 585
R1026 B.n851 B.n56 585
R1027 B.n800 B.n55 585
R1028 B.n852 B.n55 585
R1029 B.n799 B.n54 585
R1030 B.n853 B.n54 585
R1031 B.n798 B.n797 585
R1032 B.n797 B.n50 585
R1033 B.n796 B.n49 585
R1034 B.t2 B.n49 585
R1035 B.n795 B.n48 585
R1036 B.n859 B.n48 585
R1037 B.n794 B.n47 585
R1038 B.n860 B.n47 585
R1039 B.n793 B.n792 585
R1040 B.n792 B.n43 585
R1041 B.n791 B.n42 585
R1042 B.n866 B.n42 585
R1043 B.n790 B.n41 585
R1044 B.n867 B.n41 585
R1045 B.n789 B.n40 585
R1046 B.n868 B.n40 585
R1047 B.n788 B.n787 585
R1048 B.n787 B.n36 585
R1049 B.n786 B.n35 585
R1050 B.n874 B.n35 585
R1051 B.n785 B.n34 585
R1052 B.n875 B.n34 585
R1053 B.n784 B.n33 585
R1054 B.n876 B.n33 585
R1055 B.n783 B.n782 585
R1056 B.n782 B.n29 585
R1057 B.n781 B.n28 585
R1058 B.n882 B.n28 585
R1059 B.n780 B.n27 585
R1060 B.n883 B.n27 585
R1061 B.n779 B.n26 585
R1062 B.n884 B.n26 585
R1063 B.n778 B.n777 585
R1064 B.n777 B.n22 585
R1065 B.n776 B.n21 585
R1066 B.n890 B.n21 585
R1067 B.n775 B.n20 585
R1068 B.n891 B.n20 585
R1069 B.n774 B.n19 585
R1070 B.n892 B.n19 585
R1071 B.n773 B.n772 585
R1072 B.n772 B.n15 585
R1073 B.n771 B.n14 585
R1074 B.n898 B.n14 585
R1075 B.n770 B.n13 585
R1076 B.n899 B.n13 585
R1077 B.n769 B.n12 585
R1078 B.n900 B.n12 585
R1079 B.n768 B.n767 585
R1080 B.n767 B.n8 585
R1081 B.n766 B.n7 585
R1082 B.n906 B.n7 585
R1083 B.n765 B.n6 585
R1084 B.n907 B.n6 585
R1085 B.n764 B.n5 585
R1086 B.n908 B.n5 585
R1087 B.n763 B.n762 585
R1088 B.n762 B.n4 585
R1089 B.n761 B.n314 585
R1090 B.n761 B.n760 585
R1091 B.n751 B.n315 585
R1092 B.n316 B.n315 585
R1093 B.n753 B.n752 585
R1094 B.n754 B.n753 585
R1095 B.n750 B.n321 585
R1096 B.n321 B.n320 585
R1097 B.n749 B.n748 585
R1098 B.n748 B.n747 585
R1099 B.n323 B.n322 585
R1100 B.n324 B.n323 585
R1101 B.n740 B.n739 585
R1102 B.n741 B.n740 585
R1103 B.n738 B.n329 585
R1104 B.n329 B.n328 585
R1105 B.n737 B.n736 585
R1106 B.n736 B.n735 585
R1107 B.n331 B.n330 585
R1108 B.n332 B.n331 585
R1109 B.n728 B.n727 585
R1110 B.n729 B.n728 585
R1111 B.n726 B.n336 585
R1112 B.n340 B.n336 585
R1113 B.n725 B.n724 585
R1114 B.n724 B.n723 585
R1115 B.n338 B.n337 585
R1116 B.n339 B.n338 585
R1117 B.n716 B.n715 585
R1118 B.n717 B.n716 585
R1119 B.n714 B.n345 585
R1120 B.n345 B.n344 585
R1121 B.n713 B.n712 585
R1122 B.n712 B.n711 585
R1123 B.n347 B.n346 585
R1124 B.n348 B.n347 585
R1125 B.n704 B.n703 585
R1126 B.n705 B.n704 585
R1127 B.n702 B.n353 585
R1128 B.n353 B.n352 585
R1129 B.n701 B.n700 585
R1130 B.n700 B.n699 585
R1131 B.n355 B.n354 585
R1132 B.n356 B.n355 585
R1133 B.n692 B.n691 585
R1134 B.n693 B.n692 585
R1135 B.n690 B.n361 585
R1136 B.n361 B.n360 585
R1137 B.n689 B.n688 585
R1138 B.n688 B.t6 585
R1139 B.n363 B.n362 585
R1140 B.n364 B.n363 585
R1141 B.n681 B.n680 585
R1142 B.n682 B.n681 585
R1143 B.n679 B.n369 585
R1144 B.n369 B.n368 585
R1145 B.n678 B.n677 585
R1146 B.n677 B.n676 585
R1147 B.n371 B.n370 585
R1148 B.n372 B.n371 585
R1149 B.n669 B.n668 585
R1150 B.n670 B.n669 585
R1151 B.n667 B.n377 585
R1152 B.n377 B.n376 585
R1153 B.n666 B.n665 585
R1154 B.n665 B.n664 585
R1155 B.n379 B.n378 585
R1156 B.n380 B.n379 585
R1157 B.n657 B.n656 585
R1158 B.n658 B.n657 585
R1159 B.n655 B.n384 585
R1160 B.n388 B.n384 585
R1161 B.n654 B.n653 585
R1162 B.n653 B.n652 585
R1163 B.n386 B.n385 585
R1164 B.n387 B.n386 585
R1165 B.n645 B.n644 585
R1166 B.n646 B.n645 585
R1167 B.n643 B.n393 585
R1168 B.n393 B.n392 585
R1169 B.n642 B.n641 585
R1170 B.n641 B.n640 585
R1171 B.n395 B.n394 585
R1172 B.n396 B.n395 585
R1173 B.n636 B.n635 585
R1174 B.n399 B.n398 585
R1175 B.n632 B.n631 585
R1176 B.n633 B.n632 585
R1177 B.n630 B.n445 585
R1178 B.n629 B.n628 585
R1179 B.n627 B.n626 585
R1180 B.n625 B.n624 585
R1181 B.n623 B.n622 585
R1182 B.n621 B.n620 585
R1183 B.n619 B.n618 585
R1184 B.n617 B.n616 585
R1185 B.n615 B.n614 585
R1186 B.n613 B.n612 585
R1187 B.n611 B.n610 585
R1188 B.n609 B.n608 585
R1189 B.n607 B.n606 585
R1190 B.n605 B.n604 585
R1191 B.n603 B.n602 585
R1192 B.n601 B.n600 585
R1193 B.n599 B.n598 585
R1194 B.n597 B.n596 585
R1195 B.n595 B.n594 585
R1196 B.n593 B.n592 585
R1197 B.n591 B.n590 585
R1198 B.n589 B.n588 585
R1199 B.n587 B.n586 585
R1200 B.n585 B.n584 585
R1201 B.n583 B.n582 585
R1202 B.n581 B.n580 585
R1203 B.n579 B.n578 585
R1204 B.n577 B.n576 585
R1205 B.n575 B.n574 585
R1206 B.n573 B.n572 585
R1207 B.n571 B.n570 585
R1208 B.n569 B.n568 585
R1209 B.n567 B.n566 585
R1210 B.n565 B.n564 585
R1211 B.n563 B.n562 585
R1212 B.n561 B.n560 585
R1213 B.n559 B.n558 585
R1214 B.n557 B.n556 585
R1215 B.n555 B.n554 585
R1216 B.n552 B.n551 585
R1217 B.n550 B.n549 585
R1218 B.n548 B.n547 585
R1219 B.n546 B.n545 585
R1220 B.n544 B.n543 585
R1221 B.n542 B.n541 585
R1222 B.n540 B.n539 585
R1223 B.n538 B.n537 585
R1224 B.n536 B.n535 585
R1225 B.n534 B.n533 585
R1226 B.n532 B.n531 585
R1227 B.n530 B.n529 585
R1228 B.n528 B.n527 585
R1229 B.n526 B.n525 585
R1230 B.n524 B.n523 585
R1231 B.n522 B.n521 585
R1232 B.n520 B.n519 585
R1233 B.n518 B.n517 585
R1234 B.n516 B.n515 585
R1235 B.n514 B.n513 585
R1236 B.n512 B.n511 585
R1237 B.n510 B.n509 585
R1238 B.n508 B.n507 585
R1239 B.n506 B.n505 585
R1240 B.n504 B.n503 585
R1241 B.n502 B.n501 585
R1242 B.n500 B.n499 585
R1243 B.n498 B.n497 585
R1244 B.n496 B.n495 585
R1245 B.n494 B.n493 585
R1246 B.n492 B.n491 585
R1247 B.n490 B.n489 585
R1248 B.n488 B.n487 585
R1249 B.n486 B.n485 585
R1250 B.n484 B.n483 585
R1251 B.n482 B.n481 585
R1252 B.n480 B.n479 585
R1253 B.n478 B.n477 585
R1254 B.n476 B.n475 585
R1255 B.n474 B.n473 585
R1256 B.n472 B.n471 585
R1257 B.n470 B.n469 585
R1258 B.n468 B.n467 585
R1259 B.n466 B.n465 585
R1260 B.n464 B.n463 585
R1261 B.n462 B.n461 585
R1262 B.n460 B.n459 585
R1263 B.n458 B.n457 585
R1264 B.n456 B.n455 585
R1265 B.n454 B.n453 585
R1266 B.n452 B.n451 585
R1267 B.n637 B.n397 585
R1268 B.n397 B.n396 585
R1269 B.n639 B.n638 585
R1270 B.n640 B.n639 585
R1271 B.n391 B.n390 585
R1272 B.n392 B.n391 585
R1273 B.n648 B.n647 585
R1274 B.n647 B.n646 585
R1275 B.n649 B.n389 585
R1276 B.n389 B.n387 585
R1277 B.n651 B.n650 585
R1278 B.n652 B.n651 585
R1279 B.n383 B.n382 585
R1280 B.n388 B.n383 585
R1281 B.n660 B.n659 585
R1282 B.n659 B.n658 585
R1283 B.n661 B.n381 585
R1284 B.n381 B.n380 585
R1285 B.n663 B.n662 585
R1286 B.n664 B.n663 585
R1287 B.n375 B.n374 585
R1288 B.n376 B.n375 585
R1289 B.n672 B.n671 585
R1290 B.n671 B.n670 585
R1291 B.n673 B.n373 585
R1292 B.n373 B.n372 585
R1293 B.n675 B.n674 585
R1294 B.n676 B.n675 585
R1295 B.n367 B.n366 585
R1296 B.n368 B.n367 585
R1297 B.n684 B.n683 585
R1298 B.n683 B.n682 585
R1299 B.n685 B.n365 585
R1300 B.n365 B.n364 585
R1301 B.n687 B.n686 585
R1302 B.t6 B.n687 585
R1303 B.n359 B.n358 585
R1304 B.n360 B.n359 585
R1305 B.n695 B.n694 585
R1306 B.n694 B.n693 585
R1307 B.n696 B.n357 585
R1308 B.n357 B.n356 585
R1309 B.n698 B.n697 585
R1310 B.n699 B.n698 585
R1311 B.n351 B.n350 585
R1312 B.n352 B.n351 585
R1313 B.n707 B.n706 585
R1314 B.n706 B.n705 585
R1315 B.n708 B.n349 585
R1316 B.n349 B.n348 585
R1317 B.n710 B.n709 585
R1318 B.n711 B.n710 585
R1319 B.n343 B.n342 585
R1320 B.n344 B.n343 585
R1321 B.n719 B.n718 585
R1322 B.n718 B.n717 585
R1323 B.n720 B.n341 585
R1324 B.n341 B.n339 585
R1325 B.n722 B.n721 585
R1326 B.n723 B.n722 585
R1327 B.n335 B.n334 585
R1328 B.n340 B.n335 585
R1329 B.n731 B.n730 585
R1330 B.n730 B.n729 585
R1331 B.n732 B.n333 585
R1332 B.n333 B.n332 585
R1333 B.n734 B.n733 585
R1334 B.n735 B.n734 585
R1335 B.n327 B.n326 585
R1336 B.n328 B.n327 585
R1337 B.n743 B.n742 585
R1338 B.n742 B.n741 585
R1339 B.n744 B.n325 585
R1340 B.n325 B.n324 585
R1341 B.n746 B.n745 585
R1342 B.n747 B.n746 585
R1343 B.n319 B.n318 585
R1344 B.n320 B.n319 585
R1345 B.n756 B.n755 585
R1346 B.n755 B.n754 585
R1347 B.n757 B.n317 585
R1348 B.n317 B.n316 585
R1349 B.n759 B.n758 585
R1350 B.n760 B.n759 585
R1351 B.n2 B.n0 585
R1352 B.n4 B.n2 585
R1353 B.n3 B.n1 585
R1354 B.n907 B.n3 585
R1355 B.n905 B.n904 585
R1356 B.n906 B.n905 585
R1357 B.n903 B.n9 585
R1358 B.n9 B.n8 585
R1359 B.n902 B.n901 585
R1360 B.n901 B.n900 585
R1361 B.n11 B.n10 585
R1362 B.n899 B.n11 585
R1363 B.n897 B.n896 585
R1364 B.n898 B.n897 585
R1365 B.n895 B.n16 585
R1366 B.n16 B.n15 585
R1367 B.n894 B.n893 585
R1368 B.n893 B.n892 585
R1369 B.n18 B.n17 585
R1370 B.n891 B.n18 585
R1371 B.n889 B.n888 585
R1372 B.n890 B.n889 585
R1373 B.n887 B.n23 585
R1374 B.n23 B.n22 585
R1375 B.n886 B.n885 585
R1376 B.n885 B.n884 585
R1377 B.n25 B.n24 585
R1378 B.n883 B.n25 585
R1379 B.n881 B.n880 585
R1380 B.n882 B.n881 585
R1381 B.n879 B.n30 585
R1382 B.n30 B.n29 585
R1383 B.n878 B.n877 585
R1384 B.n877 B.n876 585
R1385 B.n32 B.n31 585
R1386 B.n875 B.n32 585
R1387 B.n873 B.n872 585
R1388 B.n874 B.n873 585
R1389 B.n871 B.n37 585
R1390 B.n37 B.n36 585
R1391 B.n870 B.n869 585
R1392 B.n869 B.n868 585
R1393 B.n39 B.n38 585
R1394 B.n867 B.n39 585
R1395 B.n865 B.n864 585
R1396 B.n866 B.n865 585
R1397 B.n863 B.n44 585
R1398 B.n44 B.n43 585
R1399 B.n862 B.n861 585
R1400 B.n861 B.n860 585
R1401 B.n46 B.n45 585
R1402 B.n859 B.n46 585
R1403 B.n858 B.n857 585
R1404 B.t2 B.n858 585
R1405 B.n856 B.n51 585
R1406 B.n51 B.n50 585
R1407 B.n855 B.n854 585
R1408 B.n854 B.n853 585
R1409 B.n53 B.n52 585
R1410 B.n852 B.n53 585
R1411 B.n850 B.n849 585
R1412 B.n851 B.n850 585
R1413 B.n848 B.n58 585
R1414 B.n58 B.n57 585
R1415 B.n847 B.n846 585
R1416 B.n846 B.n845 585
R1417 B.n60 B.n59 585
R1418 B.n844 B.n60 585
R1419 B.n842 B.n841 585
R1420 B.n843 B.n842 585
R1421 B.n840 B.n65 585
R1422 B.n65 B.n64 585
R1423 B.n839 B.n838 585
R1424 B.n838 B.n837 585
R1425 B.n67 B.n66 585
R1426 B.n836 B.n67 585
R1427 B.n834 B.n833 585
R1428 B.n835 B.n834 585
R1429 B.n832 B.n72 585
R1430 B.n72 B.n71 585
R1431 B.n831 B.n830 585
R1432 B.n830 B.n829 585
R1433 B.n74 B.n73 585
R1434 B.n828 B.n74 585
R1435 B.n826 B.n825 585
R1436 B.n827 B.n826 585
R1437 B.n824 B.n79 585
R1438 B.n79 B.n78 585
R1439 B.n910 B.n909 585
R1440 B.n909 B.n908 585
R1441 B.n635 B.n397 506.916
R1442 B.n822 B.n79 506.916
R1443 B.n451 B.n395 506.916
R1444 B.n819 B.n128 506.916
R1445 B.n448 B.t19 349.483
R1446 B.n446 B.t12 349.483
R1447 B.n131 B.t16 349.483
R1448 B.n129 B.t8 349.483
R1449 B.n448 B.t21 329.135
R1450 B.n446 B.t15 329.135
R1451 B.n131 B.t17 329.135
R1452 B.n129 B.t10 329.135
R1453 B.n449 B.t20 283.171
R1454 B.n130 B.t11 283.171
R1455 B.n447 B.t14 283.171
R1456 B.n132 B.t18 283.171
R1457 B.n820 B.n126 256.663
R1458 B.n820 B.n125 256.663
R1459 B.n820 B.n124 256.663
R1460 B.n820 B.n123 256.663
R1461 B.n820 B.n122 256.663
R1462 B.n820 B.n121 256.663
R1463 B.n820 B.n120 256.663
R1464 B.n820 B.n119 256.663
R1465 B.n820 B.n118 256.663
R1466 B.n820 B.n117 256.663
R1467 B.n820 B.n116 256.663
R1468 B.n820 B.n115 256.663
R1469 B.n820 B.n114 256.663
R1470 B.n820 B.n113 256.663
R1471 B.n820 B.n112 256.663
R1472 B.n820 B.n111 256.663
R1473 B.n820 B.n110 256.663
R1474 B.n820 B.n109 256.663
R1475 B.n820 B.n108 256.663
R1476 B.n820 B.n107 256.663
R1477 B.n820 B.n106 256.663
R1478 B.n820 B.n105 256.663
R1479 B.n820 B.n104 256.663
R1480 B.n820 B.n103 256.663
R1481 B.n820 B.n102 256.663
R1482 B.n820 B.n101 256.663
R1483 B.n820 B.n100 256.663
R1484 B.n820 B.n99 256.663
R1485 B.n820 B.n98 256.663
R1486 B.n820 B.n97 256.663
R1487 B.n820 B.n96 256.663
R1488 B.n820 B.n95 256.663
R1489 B.n820 B.n94 256.663
R1490 B.n820 B.n93 256.663
R1491 B.n820 B.n92 256.663
R1492 B.n820 B.n91 256.663
R1493 B.n820 B.n90 256.663
R1494 B.n820 B.n89 256.663
R1495 B.n820 B.n88 256.663
R1496 B.n820 B.n87 256.663
R1497 B.n820 B.n86 256.663
R1498 B.n820 B.n85 256.663
R1499 B.n820 B.n84 256.663
R1500 B.n820 B.n83 256.663
R1501 B.n820 B.n82 256.663
R1502 B.n821 B.n820 256.663
R1503 B.n634 B.n633 256.663
R1504 B.n633 B.n400 256.663
R1505 B.n633 B.n401 256.663
R1506 B.n633 B.n402 256.663
R1507 B.n633 B.n403 256.663
R1508 B.n633 B.n404 256.663
R1509 B.n633 B.n405 256.663
R1510 B.n633 B.n406 256.663
R1511 B.n633 B.n407 256.663
R1512 B.n633 B.n408 256.663
R1513 B.n633 B.n409 256.663
R1514 B.n633 B.n410 256.663
R1515 B.n633 B.n411 256.663
R1516 B.n633 B.n412 256.663
R1517 B.n633 B.n413 256.663
R1518 B.n633 B.n414 256.663
R1519 B.n633 B.n415 256.663
R1520 B.n633 B.n416 256.663
R1521 B.n633 B.n417 256.663
R1522 B.n633 B.n418 256.663
R1523 B.n633 B.n419 256.663
R1524 B.n633 B.n420 256.663
R1525 B.n633 B.n421 256.663
R1526 B.n633 B.n422 256.663
R1527 B.n633 B.n423 256.663
R1528 B.n633 B.n424 256.663
R1529 B.n633 B.n425 256.663
R1530 B.n633 B.n426 256.663
R1531 B.n633 B.n427 256.663
R1532 B.n633 B.n428 256.663
R1533 B.n633 B.n429 256.663
R1534 B.n633 B.n430 256.663
R1535 B.n633 B.n431 256.663
R1536 B.n633 B.n432 256.663
R1537 B.n633 B.n433 256.663
R1538 B.n633 B.n434 256.663
R1539 B.n633 B.n435 256.663
R1540 B.n633 B.n436 256.663
R1541 B.n633 B.n437 256.663
R1542 B.n633 B.n438 256.663
R1543 B.n633 B.n439 256.663
R1544 B.n633 B.n440 256.663
R1545 B.n633 B.n441 256.663
R1546 B.n633 B.n442 256.663
R1547 B.n633 B.n443 256.663
R1548 B.n633 B.n444 256.663
R1549 B.n639 B.n397 163.367
R1550 B.n639 B.n391 163.367
R1551 B.n647 B.n391 163.367
R1552 B.n647 B.n389 163.367
R1553 B.n651 B.n389 163.367
R1554 B.n651 B.n383 163.367
R1555 B.n659 B.n383 163.367
R1556 B.n659 B.n381 163.367
R1557 B.n663 B.n381 163.367
R1558 B.n663 B.n375 163.367
R1559 B.n671 B.n375 163.367
R1560 B.n671 B.n373 163.367
R1561 B.n675 B.n373 163.367
R1562 B.n675 B.n367 163.367
R1563 B.n683 B.n367 163.367
R1564 B.n683 B.n365 163.367
R1565 B.n687 B.n365 163.367
R1566 B.n687 B.n359 163.367
R1567 B.n694 B.n359 163.367
R1568 B.n694 B.n357 163.367
R1569 B.n698 B.n357 163.367
R1570 B.n698 B.n351 163.367
R1571 B.n706 B.n351 163.367
R1572 B.n706 B.n349 163.367
R1573 B.n710 B.n349 163.367
R1574 B.n710 B.n343 163.367
R1575 B.n718 B.n343 163.367
R1576 B.n718 B.n341 163.367
R1577 B.n722 B.n341 163.367
R1578 B.n722 B.n335 163.367
R1579 B.n730 B.n335 163.367
R1580 B.n730 B.n333 163.367
R1581 B.n734 B.n333 163.367
R1582 B.n734 B.n327 163.367
R1583 B.n742 B.n327 163.367
R1584 B.n742 B.n325 163.367
R1585 B.n746 B.n325 163.367
R1586 B.n746 B.n319 163.367
R1587 B.n755 B.n319 163.367
R1588 B.n755 B.n317 163.367
R1589 B.n759 B.n317 163.367
R1590 B.n759 B.n2 163.367
R1591 B.n909 B.n2 163.367
R1592 B.n909 B.n3 163.367
R1593 B.n905 B.n3 163.367
R1594 B.n905 B.n9 163.367
R1595 B.n901 B.n9 163.367
R1596 B.n901 B.n11 163.367
R1597 B.n897 B.n11 163.367
R1598 B.n897 B.n16 163.367
R1599 B.n893 B.n16 163.367
R1600 B.n893 B.n18 163.367
R1601 B.n889 B.n18 163.367
R1602 B.n889 B.n23 163.367
R1603 B.n885 B.n23 163.367
R1604 B.n885 B.n25 163.367
R1605 B.n881 B.n25 163.367
R1606 B.n881 B.n30 163.367
R1607 B.n877 B.n30 163.367
R1608 B.n877 B.n32 163.367
R1609 B.n873 B.n32 163.367
R1610 B.n873 B.n37 163.367
R1611 B.n869 B.n37 163.367
R1612 B.n869 B.n39 163.367
R1613 B.n865 B.n39 163.367
R1614 B.n865 B.n44 163.367
R1615 B.n861 B.n44 163.367
R1616 B.n861 B.n46 163.367
R1617 B.n858 B.n46 163.367
R1618 B.n858 B.n51 163.367
R1619 B.n854 B.n51 163.367
R1620 B.n854 B.n53 163.367
R1621 B.n850 B.n53 163.367
R1622 B.n850 B.n58 163.367
R1623 B.n846 B.n58 163.367
R1624 B.n846 B.n60 163.367
R1625 B.n842 B.n60 163.367
R1626 B.n842 B.n65 163.367
R1627 B.n838 B.n65 163.367
R1628 B.n838 B.n67 163.367
R1629 B.n834 B.n67 163.367
R1630 B.n834 B.n72 163.367
R1631 B.n830 B.n72 163.367
R1632 B.n830 B.n74 163.367
R1633 B.n826 B.n74 163.367
R1634 B.n826 B.n79 163.367
R1635 B.n632 B.n399 163.367
R1636 B.n632 B.n445 163.367
R1637 B.n628 B.n627 163.367
R1638 B.n624 B.n623 163.367
R1639 B.n620 B.n619 163.367
R1640 B.n616 B.n615 163.367
R1641 B.n612 B.n611 163.367
R1642 B.n608 B.n607 163.367
R1643 B.n604 B.n603 163.367
R1644 B.n600 B.n599 163.367
R1645 B.n596 B.n595 163.367
R1646 B.n592 B.n591 163.367
R1647 B.n588 B.n587 163.367
R1648 B.n584 B.n583 163.367
R1649 B.n580 B.n579 163.367
R1650 B.n576 B.n575 163.367
R1651 B.n572 B.n571 163.367
R1652 B.n568 B.n567 163.367
R1653 B.n564 B.n563 163.367
R1654 B.n560 B.n559 163.367
R1655 B.n556 B.n555 163.367
R1656 B.n551 B.n550 163.367
R1657 B.n547 B.n546 163.367
R1658 B.n543 B.n542 163.367
R1659 B.n539 B.n538 163.367
R1660 B.n535 B.n534 163.367
R1661 B.n531 B.n530 163.367
R1662 B.n527 B.n526 163.367
R1663 B.n523 B.n522 163.367
R1664 B.n519 B.n518 163.367
R1665 B.n515 B.n514 163.367
R1666 B.n511 B.n510 163.367
R1667 B.n507 B.n506 163.367
R1668 B.n503 B.n502 163.367
R1669 B.n499 B.n498 163.367
R1670 B.n495 B.n494 163.367
R1671 B.n491 B.n490 163.367
R1672 B.n487 B.n486 163.367
R1673 B.n483 B.n482 163.367
R1674 B.n479 B.n478 163.367
R1675 B.n475 B.n474 163.367
R1676 B.n471 B.n470 163.367
R1677 B.n467 B.n466 163.367
R1678 B.n463 B.n462 163.367
R1679 B.n459 B.n458 163.367
R1680 B.n455 B.n454 163.367
R1681 B.n641 B.n395 163.367
R1682 B.n641 B.n393 163.367
R1683 B.n645 B.n393 163.367
R1684 B.n645 B.n386 163.367
R1685 B.n653 B.n386 163.367
R1686 B.n653 B.n384 163.367
R1687 B.n657 B.n384 163.367
R1688 B.n657 B.n379 163.367
R1689 B.n665 B.n379 163.367
R1690 B.n665 B.n377 163.367
R1691 B.n669 B.n377 163.367
R1692 B.n669 B.n371 163.367
R1693 B.n677 B.n371 163.367
R1694 B.n677 B.n369 163.367
R1695 B.n681 B.n369 163.367
R1696 B.n681 B.n363 163.367
R1697 B.n688 B.n363 163.367
R1698 B.n688 B.n361 163.367
R1699 B.n692 B.n361 163.367
R1700 B.n692 B.n355 163.367
R1701 B.n700 B.n355 163.367
R1702 B.n700 B.n353 163.367
R1703 B.n704 B.n353 163.367
R1704 B.n704 B.n347 163.367
R1705 B.n712 B.n347 163.367
R1706 B.n712 B.n345 163.367
R1707 B.n716 B.n345 163.367
R1708 B.n716 B.n338 163.367
R1709 B.n724 B.n338 163.367
R1710 B.n724 B.n336 163.367
R1711 B.n728 B.n336 163.367
R1712 B.n728 B.n331 163.367
R1713 B.n736 B.n331 163.367
R1714 B.n736 B.n329 163.367
R1715 B.n740 B.n329 163.367
R1716 B.n740 B.n323 163.367
R1717 B.n748 B.n323 163.367
R1718 B.n748 B.n321 163.367
R1719 B.n753 B.n321 163.367
R1720 B.n753 B.n315 163.367
R1721 B.n761 B.n315 163.367
R1722 B.n762 B.n761 163.367
R1723 B.n762 B.n5 163.367
R1724 B.n6 B.n5 163.367
R1725 B.n7 B.n6 163.367
R1726 B.n767 B.n7 163.367
R1727 B.n767 B.n12 163.367
R1728 B.n13 B.n12 163.367
R1729 B.n14 B.n13 163.367
R1730 B.n772 B.n14 163.367
R1731 B.n772 B.n19 163.367
R1732 B.n20 B.n19 163.367
R1733 B.n21 B.n20 163.367
R1734 B.n777 B.n21 163.367
R1735 B.n777 B.n26 163.367
R1736 B.n27 B.n26 163.367
R1737 B.n28 B.n27 163.367
R1738 B.n782 B.n28 163.367
R1739 B.n782 B.n33 163.367
R1740 B.n34 B.n33 163.367
R1741 B.n35 B.n34 163.367
R1742 B.n787 B.n35 163.367
R1743 B.n787 B.n40 163.367
R1744 B.n41 B.n40 163.367
R1745 B.n42 B.n41 163.367
R1746 B.n792 B.n42 163.367
R1747 B.n792 B.n47 163.367
R1748 B.n48 B.n47 163.367
R1749 B.n49 B.n48 163.367
R1750 B.n797 B.n49 163.367
R1751 B.n797 B.n54 163.367
R1752 B.n55 B.n54 163.367
R1753 B.n56 B.n55 163.367
R1754 B.n802 B.n56 163.367
R1755 B.n802 B.n61 163.367
R1756 B.n62 B.n61 163.367
R1757 B.n63 B.n62 163.367
R1758 B.n807 B.n63 163.367
R1759 B.n807 B.n68 163.367
R1760 B.n69 B.n68 163.367
R1761 B.n70 B.n69 163.367
R1762 B.n812 B.n70 163.367
R1763 B.n812 B.n75 163.367
R1764 B.n76 B.n75 163.367
R1765 B.n77 B.n76 163.367
R1766 B.n128 B.n77 163.367
R1767 B.n134 B.n81 163.367
R1768 B.n138 B.n137 163.367
R1769 B.n142 B.n141 163.367
R1770 B.n146 B.n145 163.367
R1771 B.n150 B.n149 163.367
R1772 B.n154 B.n153 163.367
R1773 B.n158 B.n157 163.367
R1774 B.n162 B.n161 163.367
R1775 B.n166 B.n165 163.367
R1776 B.n170 B.n169 163.367
R1777 B.n174 B.n173 163.367
R1778 B.n178 B.n177 163.367
R1779 B.n182 B.n181 163.367
R1780 B.n186 B.n185 163.367
R1781 B.n190 B.n189 163.367
R1782 B.n194 B.n193 163.367
R1783 B.n198 B.n197 163.367
R1784 B.n202 B.n201 163.367
R1785 B.n206 B.n205 163.367
R1786 B.n210 B.n209 163.367
R1787 B.n214 B.n213 163.367
R1788 B.n218 B.n217 163.367
R1789 B.n222 B.n221 163.367
R1790 B.n226 B.n225 163.367
R1791 B.n230 B.n229 163.367
R1792 B.n235 B.n234 163.367
R1793 B.n239 B.n238 163.367
R1794 B.n243 B.n242 163.367
R1795 B.n247 B.n246 163.367
R1796 B.n251 B.n250 163.367
R1797 B.n255 B.n254 163.367
R1798 B.n259 B.n258 163.367
R1799 B.n263 B.n262 163.367
R1800 B.n267 B.n266 163.367
R1801 B.n271 B.n270 163.367
R1802 B.n275 B.n274 163.367
R1803 B.n279 B.n278 163.367
R1804 B.n283 B.n282 163.367
R1805 B.n287 B.n286 163.367
R1806 B.n291 B.n290 163.367
R1807 B.n295 B.n294 163.367
R1808 B.n299 B.n298 163.367
R1809 B.n303 B.n302 163.367
R1810 B.n307 B.n306 163.367
R1811 B.n311 B.n310 163.367
R1812 B.n819 B.n127 163.367
R1813 B.n633 B.n396 76.7816
R1814 B.n820 B.n78 76.7816
R1815 B.n635 B.n634 71.676
R1816 B.n445 B.n400 71.676
R1817 B.n627 B.n401 71.676
R1818 B.n623 B.n402 71.676
R1819 B.n619 B.n403 71.676
R1820 B.n615 B.n404 71.676
R1821 B.n611 B.n405 71.676
R1822 B.n607 B.n406 71.676
R1823 B.n603 B.n407 71.676
R1824 B.n599 B.n408 71.676
R1825 B.n595 B.n409 71.676
R1826 B.n591 B.n410 71.676
R1827 B.n587 B.n411 71.676
R1828 B.n583 B.n412 71.676
R1829 B.n579 B.n413 71.676
R1830 B.n575 B.n414 71.676
R1831 B.n571 B.n415 71.676
R1832 B.n567 B.n416 71.676
R1833 B.n563 B.n417 71.676
R1834 B.n559 B.n418 71.676
R1835 B.n555 B.n419 71.676
R1836 B.n550 B.n420 71.676
R1837 B.n546 B.n421 71.676
R1838 B.n542 B.n422 71.676
R1839 B.n538 B.n423 71.676
R1840 B.n534 B.n424 71.676
R1841 B.n530 B.n425 71.676
R1842 B.n526 B.n426 71.676
R1843 B.n522 B.n427 71.676
R1844 B.n518 B.n428 71.676
R1845 B.n514 B.n429 71.676
R1846 B.n510 B.n430 71.676
R1847 B.n506 B.n431 71.676
R1848 B.n502 B.n432 71.676
R1849 B.n498 B.n433 71.676
R1850 B.n494 B.n434 71.676
R1851 B.n490 B.n435 71.676
R1852 B.n486 B.n436 71.676
R1853 B.n482 B.n437 71.676
R1854 B.n478 B.n438 71.676
R1855 B.n474 B.n439 71.676
R1856 B.n470 B.n440 71.676
R1857 B.n466 B.n441 71.676
R1858 B.n462 B.n442 71.676
R1859 B.n458 B.n443 71.676
R1860 B.n454 B.n444 71.676
R1861 B.n822 B.n821 71.676
R1862 B.n134 B.n82 71.676
R1863 B.n138 B.n83 71.676
R1864 B.n142 B.n84 71.676
R1865 B.n146 B.n85 71.676
R1866 B.n150 B.n86 71.676
R1867 B.n154 B.n87 71.676
R1868 B.n158 B.n88 71.676
R1869 B.n162 B.n89 71.676
R1870 B.n166 B.n90 71.676
R1871 B.n170 B.n91 71.676
R1872 B.n174 B.n92 71.676
R1873 B.n178 B.n93 71.676
R1874 B.n182 B.n94 71.676
R1875 B.n186 B.n95 71.676
R1876 B.n190 B.n96 71.676
R1877 B.n194 B.n97 71.676
R1878 B.n198 B.n98 71.676
R1879 B.n202 B.n99 71.676
R1880 B.n206 B.n100 71.676
R1881 B.n210 B.n101 71.676
R1882 B.n214 B.n102 71.676
R1883 B.n218 B.n103 71.676
R1884 B.n222 B.n104 71.676
R1885 B.n226 B.n105 71.676
R1886 B.n230 B.n106 71.676
R1887 B.n235 B.n107 71.676
R1888 B.n239 B.n108 71.676
R1889 B.n243 B.n109 71.676
R1890 B.n247 B.n110 71.676
R1891 B.n251 B.n111 71.676
R1892 B.n255 B.n112 71.676
R1893 B.n259 B.n113 71.676
R1894 B.n263 B.n114 71.676
R1895 B.n267 B.n115 71.676
R1896 B.n271 B.n116 71.676
R1897 B.n275 B.n117 71.676
R1898 B.n279 B.n118 71.676
R1899 B.n283 B.n119 71.676
R1900 B.n287 B.n120 71.676
R1901 B.n291 B.n121 71.676
R1902 B.n295 B.n122 71.676
R1903 B.n299 B.n123 71.676
R1904 B.n303 B.n124 71.676
R1905 B.n307 B.n125 71.676
R1906 B.n311 B.n126 71.676
R1907 B.n127 B.n126 71.676
R1908 B.n310 B.n125 71.676
R1909 B.n306 B.n124 71.676
R1910 B.n302 B.n123 71.676
R1911 B.n298 B.n122 71.676
R1912 B.n294 B.n121 71.676
R1913 B.n290 B.n120 71.676
R1914 B.n286 B.n119 71.676
R1915 B.n282 B.n118 71.676
R1916 B.n278 B.n117 71.676
R1917 B.n274 B.n116 71.676
R1918 B.n270 B.n115 71.676
R1919 B.n266 B.n114 71.676
R1920 B.n262 B.n113 71.676
R1921 B.n258 B.n112 71.676
R1922 B.n254 B.n111 71.676
R1923 B.n250 B.n110 71.676
R1924 B.n246 B.n109 71.676
R1925 B.n242 B.n108 71.676
R1926 B.n238 B.n107 71.676
R1927 B.n234 B.n106 71.676
R1928 B.n229 B.n105 71.676
R1929 B.n225 B.n104 71.676
R1930 B.n221 B.n103 71.676
R1931 B.n217 B.n102 71.676
R1932 B.n213 B.n101 71.676
R1933 B.n209 B.n100 71.676
R1934 B.n205 B.n99 71.676
R1935 B.n201 B.n98 71.676
R1936 B.n197 B.n97 71.676
R1937 B.n193 B.n96 71.676
R1938 B.n189 B.n95 71.676
R1939 B.n185 B.n94 71.676
R1940 B.n181 B.n93 71.676
R1941 B.n177 B.n92 71.676
R1942 B.n173 B.n91 71.676
R1943 B.n169 B.n90 71.676
R1944 B.n165 B.n89 71.676
R1945 B.n161 B.n88 71.676
R1946 B.n157 B.n87 71.676
R1947 B.n153 B.n86 71.676
R1948 B.n149 B.n85 71.676
R1949 B.n145 B.n84 71.676
R1950 B.n141 B.n83 71.676
R1951 B.n137 B.n82 71.676
R1952 B.n821 B.n81 71.676
R1953 B.n634 B.n399 71.676
R1954 B.n628 B.n400 71.676
R1955 B.n624 B.n401 71.676
R1956 B.n620 B.n402 71.676
R1957 B.n616 B.n403 71.676
R1958 B.n612 B.n404 71.676
R1959 B.n608 B.n405 71.676
R1960 B.n604 B.n406 71.676
R1961 B.n600 B.n407 71.676
R1962 B.n596 B.n408 71.676
R1963 B.n592 B.n409 71.676
R1964 B.n588 B.n410 71.676
R1965 B.n584 B.n411 71.676
R1966 B.n580 B.n412 71.676
R1967 B.n576 B.n413 71.676
R1968 B.n572 B.n414 71.676
R1969 B.n568 B.n415 71.676
R1970 B.n564 B.n416 71.676
R1971 B.n560 B.n417 71.676
R1972 B.n556 B.n418 71.676
R1973 B.n551 B.n419 71.676
R1974 B.n547 B.n420 71.676
R1975 B.n543 B.n421 71.676
R1976 B.n539 B.n422 71.676
R1977 B.n535 B.n423 71.676
R1978 B.n531 B.n424 71.676
R1979 B.n527 B.n425 71.676
R1980 B.n523 B.n426 71.676
R1981 B.n519 B.n427 71.676
R1982 B.n515 B.n428 71.676
R1983 B.n511 B.n429 71.676
R1984 B.n507 B.n430 71.676
R1985 B.n503 B.n431 71.676
R1986 B.n499 B.n432 71.676
R1987 B.n495 B.n433 71.676
R1988 B.n491 B.n434 71.676
R1989 B.n487 B.n435 71.676
R1990 B.n483 B.n436 71.676
R1991 B.n479 B.n437 71.676
R1992 B.n475 B.n438 71.676
R1993 B.n471 B.n439 71.676
R1994 B.n467 B.n440 71.676
R1995 B.n463 B.n441 71.676
R1996 B.n459 B.n442 71.676
R1997 B.n455 B.n443 71.676
R1998 B.n451 B.n444 71.676
R1999 B.n450 B.n449 59.5399
R2000 B.n553 B.n447 59.5399
R2001 B.n133 B.n132 59.5399
R2002 B.n232 B.n130 59.5399
R2003 B.n449 B.n448 45.9641
R2004 B.n447 B.n446 45.9641
R2005 B.n132 B.n131 45.9641
R2006 B.n130 B.n129 45.9641
R2007 B.n640 B.n396 43.1502
R2008 B.n640 B.n392 43.1502
R2009 B.n646 B.n392 43.1502
R2010 B.n646 B.n387 43.1502
R2011 B.n652 B.n387 43.1502
R2012 B.n652 B.n388 43.1502
R2013 B.n658 B.n380 43.1502
R2014 B.n664 B.n380 43.1502
R2015 B.n664 B.n376 43.1502
R2016 B.n670 B.n376 43.1502
R2017 B.n670 B.n372 43.1502
R2018 B.n676 B.n372 43.1502
R2019 B.n676 B.n368 43.1502
R2020 B.n682 B.n368 43.1502
R2021 B.n682 B.n364 43.1502
R2022 B.t6 B.n364 43.1502
R2023 B.t6 B.n360 43.1502
R2024 B.n693 B.n360 43.1502
R2025 B.n693 B.n356 43.1502
R2026 B.n699 B.n356 43.1502
R2027 B.n699 B.n352 43.1502
R2028 B.n705 B.n352 43.1502
R2029 B.n711 B.n348 43.1502
R2030 B.n711 B.n344 43.1502
R2031 B.n717 B.n344 43.1502
R2032 B.n717 B.n339 43.1502
R2033 B.n723 B.n339 43.1502
R2034 B.n723 B.n340 43.1502
R2035 B.n729 B.n332 43.1502
R2036 B.n735 B.n332 43.1502
R2037 B.n735 B.n328 43.1502
R2038 B.n741 B.n328 43.1502
R2039 B.n741 B.n324 43.1502
R2040 B.n747 B.n324 43.1502
R2041 B.n754 B.n320 43.1502
R2042 B.n754 B.n316 43.1502
R2043 B.n760 B.n316 43.1502
R2044 B.n760 B.n4 43.1502
R2045 B.n908 B.n4 43.1502
R2046 B.n908 B.n907 43.1502
R2047 B.n907 B.n906 43.1502
R2048 B.n906 B.n8 43.1502
R2049 B.n900 B.n8 43.1502
R2050 B.n900 B.n899 43.1502
R2051 B.n898 B.n15 43.1502
R2052 B.n892 B.n15 43.1502
R2053 B.n892 B.n891 43.1502
R2054 B.n891 B.n890 43.1502
R2055 B.n890 B.n22 43.1502
R2056 B.n884 B.n22 43.1502
R2057 B.n883 B.n882 43.1502
R2058 B.n882 B.n29 43.1502
R2059 B.n876 B.n29 43.1502
R2060 B.n876 B.n875 43.1502
R2061 B.n875 B.n874 43.1502
R2062 B.n874 B.n36 43.1502
R2063 B.n868 B.n867 43.1502
R2064 B.n867 B.n866 43.1502
R2065 B.n866 B.n43 43.1502
R2066 B.n860 B.n43 43.1502
R2067 B.n860 B.n859 43.1502
R2068 B.n859 B.t2 43.1502
R2069 B.t2 B.n50 43.1502
R2070 B.n853 B.n50 43.1502
R2071 B.n853 B.n852 43.1502
R2072 B.n852 B.n851 43.1502
R2073 B.n851 B.n57 43.1502
R2074 B.n845 B.n57 43.1502
R2075 B.n845 B.n844 43.1502
R2076 B.n844 B.n843 43.1502
R2077 B.n843 B.n64 43.1502
R2078 B.n837 B.n64 43.1502
R2079 B.n836 B.n835 43.1502
R2080 B.n835 B.n71 43.1502
R2081 B.n829 B.n71 43.1502
R2082 B.n829 B.n828 43.1502
R2083 B.n828 B.n827 43.1502
R2084 B.n827 B.n78 43.1502
R2085 B.n705 B.t3 41.8811
R2086 B.n868 B.t0 41.8811
R2087 B.n340 B.t4 40.612
R2088 B.t1 B.n883 40.612
R2089 B.n747 B.t7 39.3429
R2090 B.t5 B.n898 39.3429
R2091 B.n388 B.t13 35.5355
R2092 B.t9 B.n836 35.5355
R2093 B.n824 B.n823 32.9371
R2094 B.n818 B.n817 32.9371
R2095 B.n452 B.n394 32.9371
R2096 B.n637 B.n636 32.9371
R2097 B B.n910 18.0485
R2098 B.n823 B.n80 10.6151
R2099 B.n135 B.n80 10.6151
R2100 B.n136 B.n135 10.6151
R2101 B.n139 B.n136 10.6151
R2102 B.n140 B.n139 10.6151
R2103 B.n143 B.n140 10.6151
R2104 B.n144 B.n143 10.6151
R2105 B.n147 B.n144 10.6151
R2106 B.n148 B.n147 10.6151
R2107 B.n151 B.n148 10.6151
R2108 B.n152 B.n151 10.6151
R2109 B.n155 B.n152 10.6151
R2110 B.n156 B.n155 10.6151
R2111 B.n159 B.n156 10.6151
R2112 B.n160 B.n159 10.6151
R2113 B.n163 B.n160 10.6151
R2114 B.n164 B.n163 10.6151
R2115 B.n167 B.n164 10.6151
R2116 B.n168 B.n167 10.6151
R2117 B.n171 B.n168 10.6151
R2118 B.n172 B.n171 10.6151
R2119 B.n175 B.n172 10.6151
R2120 B.n176 B.n175 10.6151
R2121 B.n179 B.n176 10.6151
R2122 B.n180 B.n179 10.6151
R2123 B.n183 B.n180 10.6151
R2124 B.n184 B.n183 10.6151
R2125 B.n187 B.n184 10.6151
R2126 B.n188 B.n187 10.6151
R2127 B.n191 B.n188 10.6151
R2128 B.n192 B.n191 10.6151
R2129 B.n195 B.n192 10.6151
R2130 B.n196 B.n195 10.6151
R2131 B.n199 B.n196 10.6151
R2132 B.n200 B.n199 10.6151
R2133 B.n203 B.n200 10.6151
R2134 B.n204 B.n203 10.6151
R2135 B.n207 B.n204 10.6151
R2136 B.n208 B.n207 10.6151
R2137 B.n211 B.n208 10.6151
R2138 B.n212 B.n211 10.6151
R2139 B.n216 B.n215 10.6151
R2140 B.n219 B.n216 10.6151
R2141 B.n220 B.n219 10.6151
R2142 B.n223 B.n220 10.6151
R2143 B.n224 B.n223 10.6151
R2144 B.n227 B.n224 10.6151
R2145 B.n228 B.n227 10.6151
R2146 B.n231 B.n228 10.6151
R2147 B.n236 B.n233 10.6151
R2148 B.n237 B.n236 10.6151
R2149 B.n240 B.n237 10.6151
R2150 B.n241 B.n240 10.6151
R2151 B.n244 B.n241 10.6151
R2152 B.n245 B.n244 10.6151
R2153 B.n248 B.n245 10.6151
R2154 B.n249 B.n248 10.6151
R2155 B.n252 B.n249 10.6151
R2156 B.n253 B.n252 10.6151
R2157 B.n256 B.n253 10.6151
R2158 B.n257 B.n256 10.6151
R2159 B.n260 B.n257 10.6151
R2160 B.n261 B.n260 10.6151
R2161 B.n264 B.n261 10.6151
R2162 B.n265 B.n264 10.6151
R2163 B.n268 B.n265 10.6151
R2164 B.n269 B.n268 10.6151
R2165 B.n272 B.n269 10.6151
R2166 B.n273 B.n272 10.6151
R2167 B.n276 B.n273 10.6151
R2168 B.n277 B.n276 10.6151
R2169 B.n280 B.n277 10.6151
R2170 B.n281 B.n280 10.6151
R2171 B.n284 B.n281 10.6151
R2172 B.n285 B.n284 10.6151
R2173 B.n288 B.n285 10.6151
R2174 B.n289 B.n288 10.6151
R2175 B.n292 B.n289 10.6151
R2176 B.n293 B.n292 10.6151
R2177 B.n296 B.n293 10.6151
R2178 B.n297 B.n296 10.6151
R2179 B.n300 B.n297 10.6151
R2180 B.n301 B.n300 10.6151
R2181 B.n304 B.n301 10.6151
R2182 B.n305 B.n304 10.6151
R2183 B.n308 B.n305 10.6151
R2184 B.n309 B.n308 10.6151
R2185 B.n312 B.n309 10.6151
R2186 B.n313 B.n312 10.6151
R2187 B.n818 B.n313 10.6151
R2188 B.n642 B.n394 10.6151
R2189 B.n643 B.n642 10.6151
R2190 B.n644 B.n643 10.6151
R2191 B.n644 B.n385 10.6151
R2192 B.n654 B.n385 10.6151
R2193 B.n655 B.n654 10.6151
R2194 B.n656 B.n655 10.6151
R2195 B.n656 B.n378 10.6151
R2196 B.n666 B.n378 10.6151
R2197 B.n667 B.n666 10.6151
R2198 B.n668 B.n667 10.6151
R2199 B.n668 B.n370 10.6151
R2200 B.n678 B.n370 10.6151
R2201 B.n679 B.n678 10.6151
R2202 B.n680 B.n679 10.6151
R2203 B.n680 B.n362 10.6151
R2204 B.n689 B.n362 10.6151
R2205 B.n690 B.n689 10.6151
R2206 B.n691 B.n690 10.6151
R2207 B.n691 B.n354 10.6151
R2208 B.n701 B.n354 10.6151
R2209 B.n702 B.n701 10.6151
R2210 B.n703 B.n702 10.6151
R2211 B.n703 B.n346 10.6151
R2212 B.n713 B.n346 10.6151
R2213 B.n714 B.n713 10.6151
R2214 B.n715 B.n714 10.6151
R2215 B.n715 B.n337 10.6151
R2216 B.n725 B.n337 10.6151
R2217 B.n726 B.n725 10.6151
R2218 B.n727 B.n726 10.6151
R2219 B.n727 B.n330 10.6151
R2220 B.n737 B.n330 10.6151
R2221 B.n738 B.n737 10.6151
R2222 B.n739 B.n738 10.6151
R2223 B.n739 B.n322 10.6151
R2224 B.n749 B.n322 10.6151
R2225 B.n750 B.n749 10.6151
R2226 B.n752 B.n750 10.6151
R2227 B.n752 B.n751 10.6151
R2228 B.n751 B.n314 10.6151
R2229 B.n763 B.n314 10.6151
R2230 B.n764 B.n763 10.6151
R2231 B.n765 B.n764 10.6151
R2232 B.n766 B.n765 10.6151
R2233 B.n768 B.n766 10.6151
R2234 B.n769 B.n768 10.6151
R2235 B.n770 B.n769 10.6151
R2236 B.n771 B.n770 10.6151
R2237 B.n773 B.n771 10.6151
R2238 B.n774 B.n773 10.6151
R2239 B.n775 B.n774 10.6151
R2240 B.n776 B.n775 10.6151
R2241 B.n778 B.n776 10.6151
R2242 B.n779 B.n778 10.6151
R2243 B.n780 B.n779 10.6151
R2244 B.n781 B.n780 10.6151
R2245 B.n783 B.n781 10.6151
R2246 B.n784 B.n783 10.6151
R2247 B.n785 B.n784 10.6151
R2248 B.n786 B.n785 10.6151
R2249 B.n788 B.n786 10.6151
R2250 B.n789 B.n788 10.6151
R2251 B.n790 B.n789 10.6151
R2252 B.n791 B.n790 10.6151
R2253 B.n793 B.n791 10.6151
R2254 B.n794 B.n793 10.6151
R2255 B.n795 B.n794 10.6151
R2256 B.n796 B.n795 10.6151
R2257 B.n798 B.n796 10.6151
R2258 B.n799 B.n798 10.6151
R2259 B.n800 B.n799 10.6151
R2260 B.n801 B.n800 10.6151
R2261 B.n803 B.n801 10.6151
R2262 B.n804 B.n803 10.6151
R2263 B.n805 B.n804 10.6151
R2264 B.n806 B.n805 10.6151
R2265 B.n808 B.n806 10.6151
R2266 B.n809 B.n808 10.6151
R2267 B.n810 B.n809 10.6151
R2268 B.n811 B.n810 10.6151
R2269 B.n813 B.n811 10.6151
R2270 B.n814 B.n813 10.6151
R2271 B.n815 B.n814 10.6151
R2272 B.n816 B.n815 10.6151
R2273 B.n817 B.n816 10.6151
R2274 B.n636 B.n398 10.6151
R2275 B.n631 B.n398 10.6151
R2276 B.n631 B.n630 10.6151
R2277 B.n630 B.n629 10.6151
R2278 B.n629 B.n626 10.6151
R2279 B.n626 B.n625 10.6151
R2280 B.n625 B.n622 10.6151
R2281 B.n622 B.n621 10.6151
R2282 B.n621 B.n618 10.6151
R2283 B.n618 B.n617 10.6151
R2284 B.n617 B.n614 10.6151
R2285 B.n614 B.n613 10.6151
R2286 B.n613 B.n610 10.6151
R2287 B.n610 B.n609 10.6151
R2288 B.n609 B.n606 10.6151
R2289 B.n606 B.n605 10.6151
R2290 B.n605 B.n602 10.6151
R2291 B.n602 B.n601 10.6151
R2292 B.n601 B.n598 10.6151
R2293 B.n598 B.n597 10.6151
R2294 B.n597 B.n594 10.6151
R2295 B.n594 B.n593 10.6151
R2296 B.n593 B.n590 10.6151
R2297 B.n590 B.n589 10.6151
R2298 B.n589 B.n586 10.6151
R2299 B.n586 B.n585 10.6151
R2300 B.n585 B.n582 10.6151
R2301 B.n582 B.n581 10.6151
R2302 B.n581 B.n578 10.6151
R2303 B.n578 B.n577 10.6151
R2304 B.n577 B.n574 10.6151
R2305 B.n574 B.n573 10.6151
R2306 B.n573 B.n570 10.6151
R2307 B.n570 B.n569 10.6151
R2308 B.n569 B.n566 10.6151
R2309 B.n566 B.n565 10.6151
R2310 B.n565 B.n562 10.6151
R2311 B.n562 B.n561 10.6151
R2312 B.n561 B.n558 10.6151
R2313 B.n558 B.n557 10.6151
R2314 B.n557 B.n554 10.6151
R2315 B.n552 B.n549 10.6151
R2316 B.n549 B.n548 10.6151
R2317 B.n548 B.n545 10.6151
R2318 B.n545 B.n544 10.6151
R2319 B.n544 B.n541 10.6151
R2320 B.n541 B.n540 10.6151
R2321 B.n540 B.n537 10.6151
R2322 B.n537 B.n536 10.6151
R2323 B.n533 B.n532 10.6151
R2324 B.n532 B.n529 10.6151
R2325 B.n529 B.n528 10.6151
R2326 B.n528 B.n525 10.6151
R2327 B.n525 B.n524 10.6151
R2328 B.n524 B.n521 10.6151
R2329 B.n521 B.n520 10.6151
R2330 B.n520 B.n517 10.6151
R2331 B.n517 B.n516 10.6151
R2332 B.n516 B.n513 10.6151
R2333 B.n513 B.n512 10.6151
R2334 B.n512 B.n509 10.6151
R2335 B.n509 B.n508 10.6151
R2336 B.n508 B.n505 10.6151
R2337 B.n505 B.n504 10.6151
R2338 B.n504 B.n501 10.6151
R2339 B.n501 B.n500 10.6151
R2340 B.n500 B.n497 10.6151
R2341 B.n497 B.n496 10.6151
R2342 B.n496 B.n493 10.6151
R2343 B.n493 B.n492 10.6151
R2344 B.n492 B.n489 10.6151
R2345 B.n489 B.n488 10.6151
R2346 B.n488 B.n485 10.6151
R2347 B.n485 B.n484 10.6151
R2348 B.n484 B.n481 10.6151
R2349 B.n481 B.n480 10.6151
R2350 B.n480 B.n477 10.6151
R2351 B.n477 B.n476 10.6151
R2352 B.n476 B.n473 10.6151
R2353 B.n473 B.n472 10.6151
R2354 B.n472 B.n469 10.6151
R2355 B.n469 B.n468 10.6151
R2356 B.n468 B.n465 10.6151
R2357 B.n465 B.n464 10.6151
R2358 B.n464 B.n461 10.6151
R2359 B.n461 B.n460 10.6151
R2360 B.n460 B.n457 10.6151
R2361 B.n457 B.n456 10.6151
R2362 B.n456 B.n453 10.6151
R2363 B.n453 B.n452 10.6151
R2364 B.n638 B.n637 10.6151
R2365 B.n638 B.n390 10.6151
R2366 B.n648 B.n390 10.6151
R2367 B.n649 B.n648 10.6151
R2368 B.n650 B.n649 10.6151
R2369 B.n650 B.n382 10.6151
R2370 B.n660 B.n382 10.6151
R2371 B.n661 B.n660 10.6151
R2372 B.n662 B.n661 10.6151
R2373 B.n662 B.n374 10.6151
R2374 B.n672 B.n374 10.6151
R2375 B.n673 B.n672 10.6151
R2376 B.n674 B.n673 10.6151
R2377 B.n674 B.n366 10.6151
R2378 B.n684 B.n366 10.6151
R2379 B.n685 B.n684 10.6151
R2380 B.n686 B.n685 10.6151
R2381 B.n686 B.n358 10.6151
R2382 B.n695 B.n358 10.6151
R2383 B.n696 B.n695 10.6151
R2384 B.n697 B.n696 10.6151
R2385 B.n697 B.n350 10.6151
R2386 B.n707 B.n350 10.6151
R2387 B.n708 B.n707 10.6151
R2388 B.n709 B.n708 10.6151
R2389 B.n709 B.n342 10.6151
R2390 B.n719 B.n342 10.6151
R2391 B.n720 B.n719 10.6151
R2392 B.n721 B.n720 10.6151
R2393 B.n721 B.n334 10.6151
R2394 B.n731 B.n334 10.6151
R2395 B.n732 B.n731 10.6151
R2396 B.n733 B.n732 10.6151
R2397 B.n733 B.n326 10.6151
R2398 B.n743 B.n326 10.6151
R2399 B.n744 B.n743 10.6151
R2400 B.n745 B.n744 10.6151
R2401 B.n745 B.n318 10.6151
R2402 B.n756 B.n318 10.6151
R2403 B.n757 B.n756 10.6151
R2404 B.n758 B.n757 10.6151
R2405 B.n758 B.n0 10.6151
R2406 B.n904 B.n1 10.6151
R2407 B.n904 B.n903 10.6151
R2408 B.n903 B.n902 10.6151
R2409 B.n902 B.n10 10.6151
R2410 B.n896 B.n10 10.6151
R2411 B.n896 B.n895 10.6151
R2412 B.n895 B.n894 10.6151
R2413 B.n894 B.n17 10.6151
R2414 B.n888 B.n17 10.6151
R2415 B.n888 B.n887 10.6151
R2416 B.n887 B.n886 10.6151
R2417 B.n886 B.n24 10.6151
R2418 B.n880 B.n24 10.6151
R2419 B.n880 B.n879 10.6151
R2420 B.n879 B.n878 10.6151
R2421 B.n878 B.n31 10.6151
R2422 B.n872 B.n31 10.6151
R2423 B.n872 B.n871 10.6151
R2424 B.n871 B.n870 10.6151
R2425 B.n870 B.n38 10.6151
R2426 B.n864 B.n38 10.6151
R2427 B.n864 B.n863 10.6151
R2428 B.n863 B.n862 10.6151
R2429 B.n862 B.n45 10.6151
R2430 B.n857 B.n45 10.6151
R2431 B.n857 B.n856 10.6151
R2432 B.n856 B.n855 10.6151
R2433 B.n855 B.n52 10.6151
R2434 B.n849 B.n52 10.6151
R2435 B.n849 B.n848 10.6151
R2436 B.n848 B.n847 10.6151
R2437 B.n847 B.n59 10.6151
R2438 B.n841 B.n59 10.6151
R2439 B.n841 B.n840 10.6151
R2440 B.n840 B.n839 10.6151
R2441 B.n839 B.n66 10.6151
R2442 B.n833 B.n66 10.6151
R2443 B.n833 B.n832 10.6151
R2444 B.n832 B.n831 10.6151
R2445 B.n831 B.n73 10.6151
R2446 B.n825 B.n73 10.6151
R2447 B.n825 B.n824 10.6151
R2448 B.n658 B.t13 7.61515
R2449 B.n837 B.t9 7.61515
R2450 B.n215 B.n133 6.5566
R2451 B.n232 B.n231 6.5566
R2452 B.n553 B.n552 6.5566
R2453 B.n536 B.n450 6.5566
R2454 B.n212 B.n133 4.05904
R2455 B.n233 B.n232 4.05904
R2456 B.n554 B.n553 4.05904
R2457 B.n533 B.n450 4.05904
R2458 B.t7 B.n320 3.80783
R2459 B.n899 B.t5 3.80783
R2460 B.n910 B.n0 2.81026
R2461 B.n910 B.n1 2.81026
R2462 B.n729 B.t4 2.53872
R2463 B.n884 B.t1 2.53872
R2464 B.t3 B.n348 1.26961
R2465 B.t0 B.n36 1.26961
R2466 VP.n13 VP.t6 175.446
R2467 VP.n15 VP.n12 161.3
R2468 VP.n17 VP.n16 161.3
R2469 VP.n18 VP.n11 161.3
R2470 VP.n20 VP.n19 161.3
R2471 VP.n22 VP.n10 161.3
R2472 VP.n24 VP.n23 161.3
R2473 VP.n25 VP.n9 161.3
R2474 VP.n27 VP.n26 161.3
R2475 VP.n28 VP.n8 161.3
R2476 VP.n54 VP.n0 161.3
R2477 VP.n53 VP.n52 161.3
R2478 VP.n51 VP.n1 161.3
R2479 VP.n50 VP.n49 161.3
R2480 VP.n48 VP.n2 161.3
R2481 VP.n46 VP.n45 161.3
R2482 VP.n44 VP.n3 161.3
R2483 VP.n43 VP.n42 161.3
R2484 VP.n41 VP.n4 161.3
R2485 VP.n39 VP.n38 161.3
R2486 VP.n37 VP.n5 161.3
R2487 VP.n36 VP.n35 161.3
R2488 VP.n34 VP.n6 161.3
R2489 VP.n33 VP.n32 161.3
R2490 VP.n7 VP.t4 142.475
R2491 VP.n40 VP.t3 142.475
R2492 VP.n47 VP.t0 142.475
R2493 VP.n55 VP.t7 142.475
R2494 VP.n29 VP.t1 142.475
R2495 VP.n21 VP.t2 142.475
R2496 VP.n14 VP.t5 142.475
R2497 VP.n31 VP.n7 95.7567
R2498 VP.n56 VP.n55 95.7567
R2499 VP.n30 VP.n29 95.7567
R2500 VP.n42 VP.n3 56.4773
R2501 VP.n16 VP.n11 56.4773
R2502 VP.n35 VP.n34 52.0954
R2503 VP.n53 VP.n1 52.0954
R2504 VP.n27 VP.n9 52.0954
R2505 VP.n14 VP.n13 49.1578
R2506 VP.n31 VP.n30 48.2798
R2507 VP.n35 VP.n5 28.7258
R2508 VP.n49 VP.n1 28.7258
R2509 VP.n23 VP.n9 28.7258
R2510 VP.n34 VP.n33 24.3439
R2511 VP.n39 VP.n5 24.3439
R2512 VP.n42 VP.n41 24.3439
R2513 VP.n46 VP.n3 24.3439
R2514 VP.n49 VP.n48 24.3439
R2515 VP.n54 VP.n53 24.3439
R2516 VP.n28 VP.n27 24.3439
R2517 VP.n20 VP.n11 24.3439
R2518 VP.n23 VP.n22 24.3439
R2519 VP.n16 VP.n15 24.3439
R2520 VP.n41 VP.n40 21.1793
R2521 VP.n47 VP.n46 21.1793
R2522 VP.n21 VP.n20 21.1793
R2523 VP.n15 VP.n14 21.1793
R2524 VP.n33 VP.n7 14.85
R2525 VP.n55 VP.n54 14.85
R2526 VP.n29 VP.n28 14.85
R2527 VP.n13 VP.n12 9.46412
R2528 VP.n40 VP.n39 3.16515
R2529 VP.n48 VP.n47 3.16515
R2530 VP.n22 VP.n21 3.16515
R2531 VP.n30 VP.n8 0.278398
R2532 VP.n32 VP.n31 0.278398
R2533 VP.n56 VP.n0 0.278398
R2534 VP.n17 VP.n12 0.189894
R2535 VP.n18 VP.n17 0.189894
R2536 VP.n19 VP.n18 0.189894
R2537 VP.n19 VP.n10 0.189894
R2538 VP.n24 VP.n10 0.189894
R2539 VP.n25 VP.n24 0.189894
R2540 VP.n26 VP.n25 0.189894
R2541 VP.n26 VP.n8 0.189894
R2542 VP.n32 VP.n6 0.189894
R2543 VP.n36 VP.n6 0.189894
R2544 VP.n37 VP.n36 0.189894
R2545 VP.n38 VP.n37 0.189894
R2546 VP.n38 VP.n4 0.189894
R2547 VP.n43 VP.n4 0.189894
R2548 VP.n44 VP.n43 0.189894
R2549 VP.n45 VP.n44 0.189894
R2550 VP.n45 VP.n2 0.189894
R2551 VP.n50 VP.n2 0.189894
R2552 VP.n51 VP.n50 0.189894
R2553 VP.n52 VP.n51 0.189894
R2554 VP.n52 VP.n0 0.189894
R2555 VP VP.n56 0.153422
R2556 VDD1 VDD1.n0 61.7961
R2557 VDD1.n3 VDD1.n2 61.6823
R2558 VDD1.n3 VDD1.n1 61.6823
R2559 VDD1.n5 VDD1.n4 60.7161
R2560 VDD1.n5 VDD1.n3 43.8888
R2561 VDD1.n4 VDD1.t5 1.64229
R2562 VDD1.n4 VDD1.t6 1.64229
R2563 VDD1.n0 VDD1.t1 1.64229
R2564 VDD1.n0 VDD1.t2 1.64229
R2565 VDD1.n2 VDD1.t7 1.64229
R2566 VDD1.n2 VDD1.t0 1.64229
R2567 VDD1.n1 VDD1.t3 1.64229
R2568 VDD1.n1 VDD1.t4 1.64229
R2569 VDD1 VDD1.n5 0.963862
C0 VP VDD2 0.459658f
C1 VDD1 VDD2 1.48535f
C2 VTAIL VP 8.505179f
C3 VTAIL VDD1 8.11463f
C4 VTAIL VDD2 8.1653f
C5 VN VP 6.99829f
C6 VN VDD1 0.150292f
C7 VN VDD2 8.280519f
C8 VN VTAIL 8.49108f
C9 VP VDD1 8.58878f
C10 VDD2 B 4.818894f
C11 VDD1 B 5.193599f
C12 VTAIL B 10.128505f
C13 VN B 13.40628f
C14 VP B 11.912911f
C15 VDD1.t1 B 0.236116f
C16 VDD1.t2 B 0.236116f
C17 VDD1.n0 B 2.11124f
C18 VDD1.t3 B 0.236116f
C19 VDD1.t4 B 0.236116f
C20 VDD1.n1 B 2.11026f
C21 VDD1.t7 B 0.236116f
C22 VDD1.t0 B 0.236116f
C23 VDD1.n2 B 2.11026f
C24 VDD1.n3 B 2.98697f
C25 VDD1.t5 B 0.236116f
C26 VDD1.t6 B 0.236116f
C27 VDD1.n4 B 2.10309f
C28 VDD1.n5 B 2.76839f
C29 VP.n0 B 0.034492f
C30 VP.t7 B 1.75386f
C31 VP.n1 B 0.026489f
C32 VP.n2 B 0.026161f
C33 VP.t0 B 1.75386f
C34 VP.n3 B 0.038356f
C35 VP.n4 B 0.026161f
C36 VP.t3 B 1.75386f
C37 VP.n5 B 0.052028f
C38 VP.n6 B 0.026161f
C39 VP.t4 B 1.75386f
C40 VP.n7 B 0.700317f
C41 VP.n8 B 0.034492f
C42 VP.t1 B 1.75386f
C43 VP.n9 B 0.026489f
C44 VP.n10 B 0.026161f
C45 VP.t2 B 1.75386f
C46 VP.n11 B 0.038356f
C47 VP.n12 B 0.21868f
C48 VP.t5 B 1.75386f
C49 VP.t6 B 1.8967f
C50 VP.n13 B 0.685573f
C51 VP.n14 B 0.699216f
C52 VP.n15 B 0.045856f
C53 VP.n16 B 0.038356f
C54 VP.n17 B 0.026161f
C55 VP.n18 B 0.026161f
C56 VP.n19 B 0.026161f
C57 VP.n20 B 0.045856f
C58 VP.n21 B 0.625433f
C59 VP.n22 B 0.027953f
C60 VP.n23 B 0.052028f
C61 VP.n24 B 0.026161f
C62 VP.n25 B 0.026161f
C63 VP.n26 B 0.026161f
C64 VP.n27 B 0.047197f
C65 VP.n28 B 0.039566f
C66 VP.n29 B 0.700317f
C67 VP.n30 B 1.3735f
C68 VP.n31 B 1.39292f
C69 VP.n32 B 0.034492f
C70 VP.n33 B 0.039566f
C71 VP.n34 B 0.047197f
C72 VP.n35 B 0.026489f
C73 VP.n36 B 0.026161f
C74 VP.n37 B 0.026161f
C75 VP.n38 B 0.026161f
C76 VP.n39 B 0.027953f
C77 VP.n40 B 0.625433f
C78 VP.n41 B 0.045856f
C79 VP.n42 B 0.038356f
C80 VP.n43 B 0.026161f
C81 VP.n44 B 0.026161f
C82 VP.n45 B 0.026161f
C83 VP.n46 B 0.045856f
C84 VP.n47 B 0.625433f
C85 VP.n48 B 0.027953f
C86 VP.n49 B 0.052028f
C87 VP.n50 B 0.026161f
C88 VP.n51 B 0.026161f
C89 VP.n52 B 0.026161f
C90 VP.n53 B 0.047197f
C91 VP.n54 B 0.039566f
C92 VP.n55 B 0.700317f
C93 VP.n56 B 0.035317f
C94 VTAIL.t14 B 0.185303f
C95 VTAIL.t15 B 0.185303f
C96 VTAIL.n0 B 1.59048f
C97 VTAIL.n1 B 0.3274f
C98 VTAIL.n2 B 0.026543f
C99 VTAIL.n3 B 0.019444f
C100 VTAIL.n4 B 0.010448f
C101 VTAIL.n5 B 0.024696f
C102 VTAIL.n6 B 0.011063f
C103 VTAIL.n7 B 0.019444f
C104 VTAIL.n8 B 0.010448f
C105 VTAIL.n9 B 0.024696f
C106 VTAIL.n10 B 0.011063f
C107 VTAIL.n11 B 0.019444f
C108 VTAIL.n12 B 0.010756f
C109 VTAIL.n13 B 0.024696f
C110 VTAIL.n14 B 0.011063f
C111 VTAIL.n15 B 0.019444f
C112 VTAIL.n16 B 0.010448f
C113 VTAIL.n17 B 0.024696f
C114 VTAIL.n18 B 0.011063f
C115 VTAIL.n19 B 0.019444f
C116 VTAIL.n20 B 0.010448f
C117 VTAIL.n21 B 0.018522f
C118 VTAIL.n22 B 0.017458f
C119 VTAIL.t11 B 0.041716f
C120 VTAIL.n23 B 0.140636f
C121 VTAIL.n24 B 0.986096f
C122 VTAIL.n25 B 0.010448f
C123 VTAIL.n26 B 0.011063f
C124 VTAIL.n27 B 0.024696f
C125 VTAIL.n28 B 0.024696f
C126 VTAIL.n29 B 0.011063f
C127 VTAIL.n30 B 0.010448f
C128 VTAIL.n31 B 0.019444f
C129 VTAIL.n32 B 0.019444f
C130 VTAIL.n33 B 0.010448f
C131 VTAIL.n34 B 0.011063f
C132 VTAIL.n35 B 0.024696f
C133 VTAIL.n36 B 0.024696f
C134 VTAIL.n37 B 0.011063f
C135 VTAIL.n38 B 0.010448f
C136 VTAIL.n39 B 0.019444f
C137 VTAIL.n40 B 0.019444f
C138 VTAIL.n41 B 0.010448f
C139 VTAIL.n42 B 0.010448f
C140 VTAIL.n43 B 0.011063f
C141 VTAIL.n44 B 0.024696f
C142 VTAIL.n45 B 0.024696f
C143 VTAIL.n46 B 0.024696f
C144 VTAIL.n47 B 0.010756f
C145 VTAIL.n48 B 0.010448f
C146 VTAIL.n49 B 0.019444f
C147 VTAIL.n50 B 0.019444f
C148 VTAIL.n51 B 0.010448f
C149 VTAIL.n52 B 0.011063f
C150 VTAIL.n53 B 0.024696f
C151 VTAIL.n54 B 0.024696f
C152 VTAIL.n55 B 0.011063f
C153 VTAIL.n56 B 0.010448f
C154 VTAIL.n57 B 0.019444f
C155 VTAIL.n58 B 0.019444f
C156 VTAIL.n59 B 0.010448f
C157 VTAIL.n60 B 0.011063f
C158 VTAIL.n61 B 0.024696f
C159 VTAIL.n62 B 0.05207f
C160 VTAIL.n63 B 0.011063f
C161 VTAIL.n64 B 0.010448f
C162 VTAIL.n65 B 0.04335f
C163 VTAIL.n66 B 0.028943f
C164 VTAIL.n67 B 0.173149f
C165 VTAIL.n68 B 0.026543f
C166 VTAIL.n69 B 0.019444f
C167 VTAIL.n70 B 0.010448f
C168 VTAIL.n71 B 0.024696f
C169 VTAIL.n72 B 0.011063f
C170 VTAIL.n73 B 0.019444f
C171 VTAIL.n74 B 0.010448f
C172 VTAIL.n75 B 0.024696f
C173 VTAIL.n76 B 0.011063f
C174 VTAIL.n77 B 0.019444f
C175 VTAIL.n78 B 0.010756f
C176 VTAIL.n79 B 0.024696f
C177 VTAIL.n80 B 0.011063f
C178 VTAIL.n81 B 0.019444f
C179 VTAIL.n82 B 0.010448f
C180 VTAIL.n83 B 0.024696f
C181 VTAIL.n84 B 0.011063f
C182 VTAIL.n85 B 0.019444f
C183 VTAIL.n86 B 0.010448f
C184 VTAIL.n87 B 0.018522f
C185 VTAIL.n88 B 0.017458f
C186 VTAIL.t7 B 0.041716f
C187 VTAIL.n89 B 0.140636f
C188 VTAIL.n90 B 0.986096f
C189 VTAIL.n91 B 0.010448f
C190 VTAIL.n92 B 0.011063f
C191 VTAIL.n93 B 0.024696f
C192 VTAIL.n94 B 0.024696f
C193 VTAIL.n95 B 0.011063f
C194 VTAIL.n96 B 0.010448f
C195 VTAIL.n97 B 0.019444f
C196 VTAIL.n98 B 0.019444f
C197 VTAIL.n99 B 0.010448f
C198 VTAIL.n100 B 0.011063f
C199 VTAIL.n101 B 0.024696f
C200 VTAIL.n102 B 0.024696f
C201 VTAIL.n103 B 0.011063f
C202 VTAIL.n104 B 0.010448f
C203 VTAIL.n105 B 0.019444f
C204 VTAIL.n106 B 0.019444f
C205 VTAIL.n107 B 0.010448f
C206 VTAIL.n108 B 0.010448f
C207 VTAIL.n109 B 0.011063f
C208 VTAIL.n110 B 0.024696f
C209 VTAIL.n111 B 0.024696f
C210 VTAIL.n112 B 0.024696f
C211 VTAIL.n113 B 0.010756f
C212 VTAIL.n114 B 0.010448f
C213 VTAIL.n115 B 0.019444f
C214 VTAIL.n116 B 0.019444f
C215 VTAIL.n117 B 0.010448f
C216 VTAIL.n118 B 0.011063f
C217 VTAIL.n119 B 0.024696f
C218 VTAIL.n120 B 0.024696f
C219 VTAIL.n121 B 0.011063f
C220 VTAIL.n122 B 0.010448f
C221 VTAIL.n123 B 0.019444f
C222 VTAIL.n124 B 0.019444f
C223 VTAIL.n125 B 0.010448f
C224 VTAIL.n126 B 0.011063f
C225 VTAIL.n127 B 0.024696f
C226 VTAIL.n128 B 0.05207f
C227 VTAIL.n129 B 0.011063f
C228 VTAIL.n130 B 0.010448f
C229 VTAIL.n131 B 0.04335f
C230 VTAIL.n132 B 0.028943f
C231 VTAIL.n133 B 0.173149f
C232 VTAIL.t3 B 0.185303f
C233 VTAIL.t4 B 0.185303f
C234 VTAIL.n134 B 1.59048f
C235 VTAIL.n135 B 0.451759f
C236 VTAIL.n136 B 0.026543f
C237 VTAIL.n137 B 0.019444f
C238 VTAIL.n138 B 0.010448f
C239 VTAIL.n139 B 0.024696f
C240 VTAIL.n140 B 0.011063f
C241 VTAIL.n141 B 0.019444f
C242 VTAIL.n142 B 0.010448f
C243 VTAIL.n143 B 0.024696f
C244 VTAIL.n144 B 0.011063f
C245 VTAIL.n145 B 0.019444f
C246 VTAIL.n146 B 0.010756f
C247 VTAIL.n147 B 0.024696f
C248 VTAIL.n148 B 0.011063f
C249 VTAIL.n149 B 0.019444f
C250 VTAIL.n150 B 0.010448f
C251 VTAIL.n151 B 0.024696f
C252 VTAIL.n152 B 0.011063f
C253 VTAIL.n153 B 0.019444f
C254 VTAIL.n154 B 0.010448f
C255 VTAIL.n155 B 0.018522f
C256 VTAIL.n156 B 0.017458f
C257 VTAIL.t6 B 0.041716f
C258 VTAIL.n157 B 0.140636f
C259 VTAIL.n158 B 0.986096f
C260 VTAIL.n159 B 0.010448f
C261 VTAIL.n160 B 0.011063f
C262 VTAIL.n161 B 0.024696f
C263 VTAIL.n162 B 0.024696f
C264 VTAIL.n163 B 0.011063f
C265 VTAIL.n164 B 0.010448f
C266 VTAIL.n165 B 0.019444f
C267 VTAIL.n166 B 0.019444f
C268 VTAIL.n167 B 0.010448f
C269 VTAIL.n168 B 0.011063f
C270 VTAIL.n169 B 0.024696f
C271 VTAIL.n170 B 0.024696f
C272 VTAIL.n171 B 0.011063f
C273 VTAIL.n172 B 0.010448f
C274 VTAIL.n173 B 0.019444f
C275 VTAIL.n174 B 0.019444f
C276 VTAIL.n175 B 0.010448f
C277 VTAIL.n176 B 0.010448f
C278 VTAIL.n177 B 0.011063f
C279 VTAIL.n178 B 0.024696f
C280 VTAIL.n179 B 0.024696f
C281 VTAIL.n180 B 0.024696f
C282 VTAIL.n181 B 0.010756f
C283 VTAIL.n182 B 0.010448f
C284 VTAIL.n183 B 0.019444f
C285 VTAIL.n184 B 0.019444f
C286 VTAIL.n185 B 0.010448f
C287 VTAIL.n186 B 0.011063f
C288 VTAIL.n187 B 0.024696f
C289 VTAIL.n188 B 0.024696f
C290 VTAIL.n189 B 0.011063f
C291 VTAIL.n190 B 0.010448f
C292 VTAIL.n191 B 0.019444f
C293 VTAIL.n192 B 0.019444f
C294 VTAIL.n193 B 0.010448f
C295 VTAIL.n194 B 0.011063f
C296 VTAIL.n195 B 0.024696f
C297 VTAIL.n196 B 0.05207f
C298 VTAIL.n197 B 0.011063f
C299 VTAIL.n198 B 0.010448f
C300 VTAIL.n199 B 0.04335f
C301 VTAIL.n200 B 0.028943f
C302 VTAIL.n201 B 1.18721f
C303 VTAIL.n202 B 0.026543f
C304 VTAIL.n203 B 0.019444f
C305 VTAIL.n204 B 0.010448f
C306 VTAIL.n205 B 0.024696f
C307 VTAIL.n206 B 0.011063f
C308 VTAIL.n207 B 0.019444f
C309 VTAIL.n208 B 0.010448f
C310 VTAIL.n209 B 0.024696f
C311 VTAIL.n210 B 0.011063f
C312 VTAIL.n211 B 0.019444f
C313 VTAIL.n212 B 0.010756f
C314 VTAIL.n213 B 0.024696f
C315 VTAIL.n214 B 0.010448f
C316 VTAIL.n215 B 0.011063f
C317 VTAIL.n216 B 0.019444f
C318 VTAIL.n217 B 0.010448f
C319 VTAIL.n218 B 0.024696f
C320 VTAIL.n219 B 0.011063f
C321 VTAIL.n220 B 0.019444f
C322 VTAIL.n221 B 0.010448f
C323 VTAIL.n222 B 0.018522f
C324 VTAIL.n223 B 0.017458f
C325 VTAIL.t13 B 0.041716f
C326 VTAIL.n224 B 0.140636f
C327 VTAIL.n225 B 0.986096f
C328 VTAIL.n226 B 0.010448f
C329 VTAIL.n227 B 0.011063f
C330 VTAIL.n228 B 0.024696f
C331 VTAIL.n229 B 0.024696f
C332 VTAIL.n230 B 0.011063f
C333 VTAIL.n231 B 0.010448f
C334 VTAIL.n232 B 0.019444f
C335 VTAIL.n233 B 0.019444f
C336 VTAIL.n234 B 0.010448f
C337 VTAIL.n235 B 0.011063f
C338 VTAIL.n236 B 0.024696f
C339 VTAIL.n237 B 0.024696f
C340 VTAIL.n238 B 0.011063f
C341 VTAIL.n239 B 0.010448f
C342 VTAIL.n240 B 0.019444f
C343 VTAIL.n241 B 0.019444f
C344 VTAIL.n242 B 0.010448f
C345 VTAIL.n243 B 0.011063f
C346 VTAIL.n244 B 0.024696f
C347 VTAIL.n245 B 0.024696f
C348 VTAIL.n246 B 0.024696f
C349 VTAIL.n247 B 0.010756f
C350 VTAIL.n248 B 0.010448f
C351 VTAIL.n249 B 0.019444f
C352 VTAIL.n250 B 0.019444f
C353 VTAIL.n251 B 0.010448f
C354 VTAIL.n252 B 0.011063f
C355 VTAIL.n253 B 0.024696f
C356 VTAIL.n254 B 0.024696f
C357 VTAIL.n255 B 0.011063f
C358 VTAIL.n256 B 0.010448f
C359 VTAIL.n257 B 0.019444f
C360 VTAIL.n258 B 0.019444f
C361 VTAIL.n259 B 0.010448f
C362 VTAIL.n260 B 0.011063f
C363 VTAIL.n261 B 0.024696f
C364 VTAIL.n262 B 0.05207f
C365 VTAIL.n263 B 0.011063f
C366 VTAIL.n264 B 0.010448f
C367 VTAIL.n265 B 0.04335f
C368 VTAIL.n266 B 0.028943f
C369 VTAIL.n267 B 1.18721f
C370 VTAIL.t12 B 0.185303f
C371 VTAIL.t10 B 0.185303f
C372 VTAIL.n268 B 1.59049f
C373 VTAIL.n269 B 0.45175f
C374 VTAIL.n270 B 0.026543f
C375 VTAIL.n271 B 0.019444f
C376 VTAIL.n272 B 0.010448f
C377 VTAIL.n273 B 0.024696f
C378 VTAIL.n274 B 0.011063f
C379 VTAIL.n275 B 0.019444f
C380 VTAIL.n276 B 0.010448f
C381 VTAIL.n277 B 0.024696f
C382 VTAIL.n278 B 0.011063f
C383 VTAIL.n279 B 0.019444f
C384 VTAIL.n280 B 0.010756f
C385 VTAIL.n281 B 0.024696f
C386 VTAIL.n282 B 0.010448f
C387 VTAIL.n283 B 0.011063f
C388 VTAIL.n284 B 0.019444f
C389 VTAIL.n285 B 0.010448f
C390 VTAIL.n286 B 0.024696f
C391 VTAIL.n287 B 0.011063f
C392 VTAIL.n288 B 0.019444f
C393 VTAIL.n289 B 0.010448f
C394 VTAIL.n290 B 0.018522f
C395 VTAIL.n291 B 0.017458f
C396 VTAIL.t9 B 0.041716f
C397 VTAIL.n292 B 0.140636f
C398 VTAIL.n293 B 0.986096f
C399 VTAIL.n294 B 0.010448f
C400 VTAIL.n295 B 0.011063f
C401 VTAIL.n296 B 0.024696f
C402 VTAIL.n297 B 0.024696f
C403 VTAIL.n298 B 0.011063f
C404 VTAIL.n299 B 0.010448f
C405 VTAIL.n300 B 0.019444f
C406 VTAIL.n301 B 0.019444f
C407 VTAIL.n302 B 0.010448f
C408 VTAIL.n303 B 0.011063f
C409 VTAIL.n304 B 0.024696f
C410 VTAIL.n305 B 0.024696f
C411 VTAIL.n306 B 0.011063f
C412 VTAIL.n307 B 0.010448f
C413 VTAIL.n308 B 0.019444f
C414 VTAIL.n309 B 0.019444f
C415 VTAIL.n310 B 0.010448f
C416 VTAIL.n311 B 0.011063f
C417 VTAIL.n312 B 0.024696f
C418 VTAIL.n313 B 0.024696f
C419 VTAIL.n314 B 0.024696f
C420 VTAIL.n315 B 0.010756f
C421 VTAIL.n316 B 0.010448f
C422 VTAIL.n317 B 0.019444f
C423 VTAIL.n318 B 0.019444f
C424 VTAIL.n319 B 0.010448f
C425 VTAIL.n320 B 0.011063f
C426 VTAIL.n321 B 0.024696f
C427 VTAIL.n322 B 0.024696f
C428 VTAIL.n323 B 0.011063f
C429 VTAIL.n324 B 0.010448f
C430 VTAIL.n325 B 0.019444f
C431 VTAIL.n326 B 0.019444f
C432 VTAIL.n327 B 0.010448f
C433 VTAIL.n328 B 0.011063f
C434 VTAIL.n329 B 0.024696f
C435 VTAIL.n330 B 0.05207f
C436 VTAIL.n331 B 0.011063f
C437 VTAIL.n332 B 0.010448f
C438 VTAIL.n333 B 0.04335f
C439 VTAIL.n334 B 0.028943f
C440 VTAIL.n335 B 0.173149f
C441 VTAIL.n336 B 0.026543f
C442 VTAIL.n337 B 0.019444f
C443 VTAIL.n338 B 0.010448f
C444 VTAIL.n339 B 0.024696f
C445 VTAIL.n340 B 0.011063f
C446 VTAIL.n341 B 0.019444f
C447 VTAIL.n342 B 0.010448f
C448 VTAIL.n343 B 0.024696f
C449 VTAIL.n344 B 0.011063f
C450 VTAIL.n345 B 0.019444f
C451 VTAIL.n346 B 0.010756f
C452 VTAIL.n347 B 0.024696f
C453 VTAIL.n348 B 0.010448f
C454 VTAIL.n349 B 0.011063f
C455 VTAIL.n350 B 0.019444f
C456 VTAIL.n351 B 0.010448f
C457 VTAIL.n352 B 0.024696f
C458 VTAIL.n353 B 0.011063f
C459 VTAIL.n354 B 0.019444f
C460 VTAIL.n355 B 0.010448f
C461 VTAIL.n356 B 0.018522f
C462 VTAIL.n357 B 0.017458f
C463 VTAIL.t5 B 0.041716f
C464 VTAIL.n358 B 0.140636f
C465 VTAIL.n359 B 0.986096f
C466 VTAIL.n360 B 0.010448f
C467 VTAIL.n361 B 0.011063f
C468 VTAIL.n362 B 0.024696f
C469 VTAIL.n363 B 0.024696f
C470 VTAIL.n364 B 0.011063f
C471 VTAIL.n365 B 0.010448f
C472 VTAIL.n366 B 0.019444f
C473 VTAIL.n367 B 0.019444f
C474 VTAIL.n368 B 0.010448f
C475 VTAIL.n369 B 0.011063f
C476 VTAIL.n370 B 0.024696f
C477 VTAIL.n371 B 0.024696f
C478 VTAIL.n372 B 0.011063f
C479 VTAIL.n373 B 0.010448f
C480 VTAIL.n374 B 0.019444f
C481 VTAIL.n375 B 0.019444f
C482 VTAIL.n376 B 0.010448f
C483 VTAIL.n377 B 0.011063f
C484 VTAIL.n378 B 0.024696f
C485 VTAIL.n379 B 0.024696f
C486 VTAIL.n380 B 0.024696f
C487 VTAIL.n381 B 0.010756f
C488 VTAIL.n382 B 0.010448f
C489 VTAIL.n383 B 0.019444f
C490 VTAIL.n384 B 0.019444f
C491 VTAIL.n385 B 0.010448f
C492 VTAIL.n386 B 0.011063f
C493 VTAIL.n387 B 0.024696f
C494 VTAIL.n388 B 0.024696f
C495 VTAIL.n389 B 0.011063f
C496 VTAIL.n390 B 0.010448f
C497 VTAIL.n391 B 0.019444f
C498 VTAIL.n392 B 0.019444f
C499 VTAIL.n393 B 0.010448f
C500 VTAIL.n394 B 0.011063f
C501 VTAIL.n395 B 0.024696f
C502 VTAIL.n396 B 0.05207f
C503 VTAIL.n397 B 0.011063f
C504 VTAIL.n398 B 0.010448f
C505 VTAIL.n399 B 0.04335f
C506 VTAIL.n400 B 0.028943f
C507 VTAIL.n401 B 0.173149f
C508 VTAIL.t1 B 0.185303f
C509 VTAIL.t0 B 0.185303f
C510 VTAIL.n402 B 1.59049f
C511 VTAIL.n403 B 0.45175f
C512 VTAIL.n404 B 0.026543f
C513 VTAIL.n405 B 0.019444f
C514 VTAIL.n406 B 0.010448f
C515 VTAIL.n407 B 0.024696f
C516 VTAIL.n408 B 0.011063f
C517 VTAIL.n409 B 0.019444f
C518 VTAIL.n410 B 0.010448f
C519 VTAIL.n411 B 0.024696f
C520 VTAIL.n412 B 0.011063f
C521 VTAIL.n413 B 0.019444f
C522 VTAIL.n414 B 0.010756f
C523 VTAIL.n415 B 0.024696f
C524 VTAIL.n416 B 0.010448f
C525 VTAIL.n417 B 0.011063f
C526 VTAIL.n418 B 0.019444f
C527 VTAIL.n419 B 0.010448f
C528 VTAIL.n420 B 0.024696f
C529 VTAIL.n421 B 0.011063f
C530 VTAIL.n422 B 0.019444f
C531 VTAIL.n423 B 0.010448f
C532 VTAIL.n424 B 0.018522f
C533 VTAIL.n425 B 0.017458f
C534 VTAIL.t2 B 0.041716f
C535 VTAIL.n426 B 0.140636f
C536 VTAIL.n427 B 0.986096f
C537 VTAIL.n428 B 0.010448f
C538 VTAIL.n429 B 0.011063f
C539 VTAIL.n430 B 0.024696f
C540 VTAIL.n431 B 0.024696f
C541 VTAIL.n432 B 0.011063f
C542 VTAIL.n433 B 0.010448f
C543 VTAIL.n434 B 0.019444f
C544 VTAIL.n435 B 0.019444f
C545 VTAIL.n436 B 0.010448f
C546 VTAIL.n437 B 0.011063f
C547 VTAIL.n438 B 0.024696f
C548 VTAIL.n439 B 0.024696f
C549 VTAIL.n440 B 0.011063f
C550 VTAIL.n441 B 0.010448f
C551 VTAIL.n442 B 0.019444f
C552 VTAIL.n443 B 0.019444f
C553 VTAIL.n444 B 0.010448f
C554 VTAIL.n445 B 0.011063f
C555 VTAIL.n446 B 0.024696f
C556 VTAIL.n447 B 0.024696f
C557 VTAIL.n448 B 0.024696f
C558 VTAIL.n449 B 0.010756f
C559 VTAIL.n450 B 0.010448f
C560 VTAIL.n451 B 0.019444f
C561 VTAIL.n452 B 0.019444f
C562 VTAIL.n453 B 0.010448f
C563 VTAIL.n454 B 0.011063f
C564 VTAIL.n455 B 0.024696f
C565 VTAIL.n456 B 0.024696f
C566 VTAIL.n457 B 0.011063f
C567 VTAIL.n458 B 0.010448f
C568 VTAIL.n459 B 0.019444f
C569 VTAIL.n460 B 0.019444f
C570 VTAIL.n461 B 0.010448f
C571 VTAIL.n462 B 0.011063f
C572 VTAIL.n463 B 0.024696f
C573 VTAIL.n464 B 0.05207f
C574 VTAIL.n465 B 0.011063f
C575 VTAIL.n466 B 0.010448f
C576 VTAIL.n467 B 0.04335f
C577 VTAIL.n468 B 0.028943f
C578 VTAIL.n469 B 1.18721f
C579 VTAIL.n470 B 0.026543f
C580 VTAIL.n471 B 0.019444f
C581 VTAIL.n472 B 0.010448f
C582 VTAIL.n473 B 0.024696f
C583 VTAIL.n474 B 0.011063f
C584 VTAIL.n475 B 0.019444f
C585 VTAIL.n476 B 0.010448f
C586 VTAIL.n477 B 0.024696f
C587 VTAIL.n478 B 0.011063f
C588 VTAIL.n479 B 0.019444f
C589 VTAIL.n480 B 0.010756f
C590 VTAIL.n481 B 0.024696f
C591 VTAIL.n482 B 0.011063f
C592 VTAIL.n483 B 0.019444f
C593 VTAIL.n484 B 0.010448f
C594 VTAIL.n485 B 0.024696f
C595 VTAIL.n486 B 0.011063f
C596 VTAIL.n487 B 0.019444f
C597 VTAIL.n488 B 0.010448f
C598 VTAIL.n489 B 0.018522f
C599 VTAIL.n490 B 0.017458f
C600 VTAIL.t8 B 0.041716f
C601 VTAIL.n491 B 0.140636f
C602 VTAIL.n492 B 0.986096f
C603 VTAIL.n493 B 0.010448f
C604 VTAIL.n494 B 0.011063f
C605 VTAIL.n495 B 0.024696f
C606 VTAIL.n496 B 0.024696f
C607 VTAIL.n497 B 0.011063f
C608 VTAIL.n498 B 0.010448f
C609 VTAIL.n499 B 0.019444f
C610 VTAIL.n500 B 0.019444f
C611 VTAIL.n501 B 0.010448f
C612 VTAIL.n502 B 0.011063f
C613 VTAIL.n503 B 0.024696f
C614 VTAIL.n504 B 0.024696f
C615 VTAIL.n505 B 0.011063f
C616 VTAIL.n506 B 0.010448f
C617 VTAIL.n507 B 0.019444f
C618 VTAIL.n508 B 0.019444f
C619 VTAIL.n509 B 0.010448f
C620 VTAIL.n510 B 0.010448f
C621 VTAIL.n511 B 0.011063f
C622 VTAIL.n512 B 0.024696f
C623 VTAIL.n513 B 0.024696f
C624 VTAIL.n514 B 0.024696f
C625 VTAIL.n515 B 0.010756f
C626 VTAIL.n516 B 0.010448f
C627 VTAIL.n517 B 0.019444f
C628 VTAIL.n518 B 0.019444f
C629 VTAIL.n519 B 0.010448f
C630 VTAIL.n520 B 0.011063f
C631 VTAIL.n521 B 0.024696f
C632 VTAIL.n522 B 0.024696f
C633 VTAIL.n523 B 0.011063f
C634 VTAIL.n524 B 0.010448f
C635 VTAIL.n525 B 0.019444f
C636 VTAIL.n526 B 0.019444f
C637 VTAIL.n527 B 0.010448f
C638 VTAIL.n528 B 0.011063f
C639 VTAIL.n529 B 0.024696f
C640 VTAIL.n530 B 0.05207f
C641 VTAIL.n531 B 0.011063f
C642 VTAIL.n532 B 0.010448f
C643 VTAIL.n533 B 0.04335f
C644 VTAIL.n534 B 0.028943f
C645 VTAIL.n535 B 1.18356f
C646 VDD2.t2 B 0.234574f
C647 VDD2.t7 B 0.234574f
C648 VDD2.n0 B 2.09647f
C649 VDD2.t5 B 0.234574f
C650 VDD2.t1 B 0.234574f
C651 VDD2.n1 B 2.09647f
C652 VDD2.n2 B 2.91586f
C653 VDD2.t6 B 0.234574f
C654 VDD2.t4 B 0.234574f
C655 VDD2.n3 B 2.08936f
C656 VDD2.n4 B 2.7202f
C657 VDD2.t3 B 0.234574f
C658 VDD2.t0 B 0.234574f
C659 VDD2.n5 B 2.09644f
C660 VN.n0 B 0.034011f
C661 VN.t7 B 1.72939f
C662 VN.n1 B 0.026119f
C663 VN.n2 B 0.025796f
C664 VN.t0 B 1.72939f
C665 VN.n3 B 0.037821f
C666 VN.n4 B 0.215628f
C667 VN.t1 B 1.72939f
C668 VN.t4 B 1.87024f
C669 VN.n5 B 0.676007f
C670 VN.n6 B 0.68946f
C671 VN.n7 B 0.045216f
C672 VN.n8 B 0.037821f
C673 VN.n9 B 0.025796f
C674 VN.n10 B 0.025796f
C675 VN.n11 B 0.025796f
C676 VN.n12 B 0.045216f
C677 VN.n13 B 0.616707f
C678 VN.n14 B 0.027563f
C679 VN.n15 B 0.051302f
C680 VN.n16 B 0.025796f
C681 VN.n17 B 0.025796f
C682 VN.n18 B 0.025796f
C683 VN.n19 B 0.046539f
C684 VN.n20 B 0.039014f
C685 VN.n21 B 0.690546f
C686 VN.n22 B 0.034824f
C687 VN.n23 B 0.034011f
C688 VN.t2 B 1.72939f
C689 VN.n24 B 0.026119f
C690 VN.n25 B 0.025796f
C691 VN.t3 B 1.72939f
C692 VN.n26 B 0.037821f
C693 VN.n27 B 0.215628f
C694 VN.t5 B 1.72939f
C695 VN.t6 B 1.87024f
C696 VN.n28 B 0.676007f
C697 VN.n29 B 0.68946f
C698 VN.n30 B 0.045216f
C699 VN.n31 B 0.037821f
C700 VN.n32 B 0.025796f
C701 VN.n33 B 0.025796f
C702 VN.n34 B 0.025796f
C703 VN.n35 B 0.045216f
C704 VN.n36 B 0.616707f
C705 VN.n37 B 0.027563f
C706 VN.n38 B 0.051302f
C707 VN.n39 B 0.025796f
C708 VN.n40 B 0.025796f
C709 VN.n41 B 0.025796f
C710 VN.n42 B 0.046539f
C711 VN.n43 B 0.039014f
C712 VN.n44 B 0.690546f
C713 VN.n45 B 1.36828f
.ends

