* NGSPICE file created from diff_pair_sample_0147.ext - technology: sky130A

.subckt diff_pair_sample_0147 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=4.0443 ps=21.52 w=10.37 l=3.84
X1 B.t11 B.t9 B.t10 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=0 ps=0 w=10.37 l=3.84
X2 B.t8 B.t6 B.t7 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=0 ps=0 w=10.37 l=3.84
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=4.0443 ps=21.52 w=10.37 l=3.84
X4 B.t5 B.t3 B.t4 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=0 ps=0 w=10.37 l=3.84
X5 VDD1.t0 VP.t1 VTAIL.t3 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=4.0443 ps=21.52 w=10.37 l=3.84
X6 VDD2.t0 VN.t1 VTAIL.t1 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=4.0443 ps=21.52 w=10.37 l=3.84
X7 B.t2 B.t0 B.t1 w_n2638_n3042# sky130_fd_pr__pfet_01v8 ad=4.0443 pd=21.52 as=0 ps=0 w=10.37 l=3.84
R0 VP.n0 VP.t1 146.831
R1 VP.n0 VP.t0 100.121
R2 VP VP.n0 0.621237
R3 VTAIL.n1 VTAIL.t1 63.8941
R4 VTAIL.n2 VTAIL.t3 63.8939
R5 VTAIL.n3 VTAIL.t0 63.8939
R6 VTAIL.n0 VTAIL.t2 63.8939
R7 VTAIL.n1 VTAIL.n0 28.4962
R8 VTAIL.n3 VTAIL.n2 24.9014
R9 VTAIL.n2 VTAIL.n1 2.26774
R10 VTAIL VTAIL.n0 1.42722
R11 VTAIL VTAIL.n3 0.841017
R12 VDD1 VDD1.t1 121.784
R13 VDD1 VDD1.t0 81.5296
R14 B.n331 B.n330 585
R15 B.n329 B.n98 585
R16 B.n328 B.n327 585
R17 B.n326 B.n99 585
R18 B.n325 B.n324 585
R19 B.n323 B.n100 585
R20 B.n322 B.n321 585
R21 B.n320 B.n101 585
R22 B.n319 B.n318 585
R23 B.n317 B.n102 585
R24 B.n316 B.n315 585
R25 B.n314 B.n103 585
R26 B.n313 B.n312 585
R27 B.n311 B.n104 585
R28 B.n310 B.n309 585
R29 B.n308 B.n105 585
R30 B.n307 B.n306 585
R31 B.n305 B.n106 585
R32 B.n304 B.n303 585
R33 B.n302 B.n107 585
R34 B.n301 B.n300 585
R35 B.n299 B.n108 585
R36 B.n298 B.n297 585
R37 B.n296 B.n109 585
R38 B.n295 B.n294 585
R39 B.n293 B.n110 585
R40 B.n292 B.n291 585
R41 B.n290 B.n111 585
R42 B.n289 B.n288 585
R43 B.n287 B.n112 585
R44 B.n286 B.n285 585
R45 B.n284 B.n113 585
R46 B.n283 B.n282 585
R47 B.n281 B.n114 585
R48 B.n280 B.n279 585
R49 B.n278 B.n115 585
R50 B.n277 B.n276 585
R51 B.n274 B.n116 585
R52 B.n273 B.n272 585
R53 B.n271 B.n119 585
R54 B.n270 B.n269 585
R55 B.n268 B.n120 585
R56 B.n267 B.n266 585
R57 B.n265 B.n121 585
R58 B.n264 B.n263 585
R59 B.n262 B.n122 585
R60 B.n260 B.n259 585
R61 B.n258 B.n125 585
R62 B.n257 B.n256 585
R63 B.n255 B.n126 585
R64 B.n254 B.n253 585
R65 B.n252 B.n127 585
R66 B.n251 B.n250 585
R67 B.n249 B.n128 585
R68 B.n248 B.n247 585
R69 B.n246 B.n129 585
R70 B.n245 B.n244 585
R71 B.n243 B.n130 585
R72 B.n242 B.n241 585
R73 B.n240 B.n131 585
R74 B.n239 B.n238 585
R75 B.n237 B.n132 585
R76 B.n236 B.n235 585
R77 B.n234 B.n133 585
R78 B.n233 B.n232 585
R79 B.n231 B.n134 585
R80 B.n230 B.n229 585
R81 B.n228 B.n135 585
R82 B.n227 B.n226 585
R83 B.n225 B.n136 585
R84 B.n224 B.n223 585
R85 B.n222 B.n137 585
R86 B.n221 B.n220 585
R87 B.n219 B.n138 585
R88 B.n218 B.n217 585
R89 B.n216 B.n139 585
R90 B.n215 B.n214 585
R91 B.n213 B.n140 585
R92 B.n212 B.n211 585
R93 B.n210 B.n141 585
R94 B.n209 B.n208 585
R95 B.n207 B.n142 585
R96 B.n206 B.n205 585
R97 B.n332 B.n97 585
R98 B.n334 B.n333 585
R99 B.n335 B.n96 585
R100 B.n337 B.n336 585
R101 B.n338 B.n95 585
R102 B.n340 B.n339 585
R103 B.n341 B.n94 585
R104 B.n343 B.n342 585
R105 B.n344 B.n93 585
R106 B.n346 B.n345 585
R107 B.n347 B.n92 585
R108 B.n349 B.n348 585
R109 B.n350 B.n91 585
R110 B.n352 B.n351 585
R111 B.n353 B.n90 585
R112 B.n355 B.n354 585
R113 B.n356 B.n89 585
R114 B.n358 B.n357 585
R115 B.n359 B.n88 585
R116 B.n361 B.n360 585
R117 B.n362 B.n87 585
R118 B.n364 B.n363 585
R119 B.n365 B.n86 585
R120 B.n367 B.n366 585
R121 B.n368 B.n85 585
R122 B.n370 B.n369 585
R123 B.n371 B.n84 585
R124 B.n373 B.n372 585
R125 B.n374 B.n83 585
R126 B.n376 B.n375 585
R127 B.n377 B.n82 585
R128 B.n379 B.n378 585
R129 B.n380 B.n81 585
R130 B.n382 B.n381 585
R131 B.n383 B.n80 585
R132 B.n385 B.n384 585
R133 B.n386 B.n79 585
R134 B.n388 B.n387 585
R135 B.n389 B.n78 585
R136 B.n391 B.n390 585
R137 B.n392 B.n77 585
R138 B.n394 B.n393 585
R139 B.n395 B.n76 585
R140 B.n397 B.n396 585
R141 B.n398 B.n75 585
R142 B.n400 B.n399 585
R143 B.n401 B.n74 585
R144 B.n403 B.n402 585
R145 B.n404 B.n73 585
R146 B.n406 B.n405 585
R147 B.n407 B.n72 585
R148 B.n409 B.n408 585
R149 B.n410 B.n71 585
R150 B.n412 B.n411 585
R151 B.n413 B.n70 585
R152 B.n415 B.n414 585
R153 B.n416 B.n69 585
R154 B.n418 B.n417 585
R155 B.n419 B.n68 585
R156 B.n421 B.n420 585
R157 B.n422 B.n67 585
R158 B.n424 B.n423 585
R159 B.n425 B.n66 585
R160 B.n427 B.n426 585
R161 B.n428 B.n65 585
R162 B.n430 B.n429 585
R163 B.n555 B.n18 585
R164 B.n554 B.n553 585
R165 B.n552 B.n19 585
R166 B.n551 B.n550 585
R167 B.n549 B.n20 585
R168 B.n548 B.n547 585
R169 B.n546 B.n21 585
R170 B.n545 B.n544 585
R171 B.n543 B.n22 585
R172 B.n542 B.n541 585
R173 B.n540 B.n23 585
R174 B.n539 B.n538 585
R175 B.n537 B.n24 585
R176 B.n536 B.n535 585
R177 B.n534 B.n25 585
R178 B.n533 B.n532 585
R179 B.n531 B.n26 585
R180 B.n530 B.n529 585
R181 B.n528 B.n27 585
R182 B.n527 B.n526 585
R183 B.n525 B.n28 585
R184 B.n524 B.n523 585
R185 B.n522 B.n29 585
R186 B.n521 B.n520 585
R187 B.n519 B.n30 585
R188 B.n518 B.n517 585
R189 B.n516 B.n31 585
R190 B.n515 B.n514 585
R191 B.n513 B.n32 585
R192 B.n512 B.n511 585
R193 B.n510 B.n33 585
R194 B.n509 B.n508 585
R195 B.n507 B.n34 585
R196 B.n506 B.n505 585
R197 B.n504 B.n35 585
R198 B.n503 B.n502 585
R199 B.n501 B.n36 585
R200 B.n500 B.n499 585
R201 B.n498 B.n37 585
R202 B.n497 B.n496 585
R203 B.n495 B.n41 585
R204 B.n494 B.n493 585
R205 B.n492 B.n42 585
R206 B.n491 B.n490 585
R207 B.n489 B.n43 585
R208 B.n488 B.n487 585
R209 B.n485 B.n44 585
R210 B.n484 B.n483 585
R211 B.n482 B.n47 585
R212 B.n481 B.n480 585
R213 B.n479 B.n48 585
R214 B.n478 B.n477 585
R215 B.n476 B.n49 585
R216 B.n475 B.n474 585
R217 B.n473 B.n50 585
R218 B.n472 B.n471 585
R219 B.n470 B.n51 585
R220 B.n469 B.n468 585
R221 B.n467 B.n52 585
R222 B.n466 B.n465 585
R223 B.n464 B.n53 585
R224 B.n463 B.n462 585
R225 B.n461 B.n54 585
R226 B.n460 B.n459 585
R227 B.n458 B.n55 585
R228 B.n457 B.n456 585
R229 B.n455 B.n56 585
R230 B.n454 B.n453 585
R231 B.n452 B.n57 585
R232 B.n451 B.n450 585
R233 B.n449 B.n58 585
R234 B.n448 B.n447 585
R235 B.n446 B.n59 585
R236 B.n445 B.n444 585
R237 B.n443 B.n60 585
R238 B.n442 B.n441 585
R239 B.n440 B.n61 585
R240 B.n439 B.n438 585
R241 B.n437 B.n62 585
R242 B.n436 B.n435 585
R243 B.n434 B.n63 585
R244 B.n433 B.n432 585
R245 B.n431 B.n64 585
R246 B.n557 B.n556 585
R247 B.n558 B.n17 585
R248 B.n560 B.n559 585
R249 B.n561 B.n16 585
R250 B.n563 B.n562 585
R251 B.n564 B.n15 585
R252 B.n566 B.n565 585
R253 B.n567 B.n14 585
R254 B.n569 B.n568 585
R255 B.n570 B.n13 585
R256 B.n572 B.n571 585
R257 B.n573 B.n12 585
R258 B.n575 B.n574 585
R259 B.n576 B.n11 585
R260 B.n578 B.n577 585
R261 B.n579 B.n10 585
R262 B.n581 B.n580 585
R263 B.n582 B.n9 585
R264 B.n584 B.n583 585
R265 B.n585 B.n8 585
R266 B.n587 B.n586 585
R267 B.n588 B.n7 585
R268 B.n590 B.n589 585
R269 B.n591 B.n6 585
R270 B.n593 B.n592 585
R271 B.n594 B.n5 585
R272 B.n596 B.n595 585
R273 B.n597 B.n4 585
R274 B.n599 B.n598 585
R275 B.n600 B.n3 585
R276 B.n602 B.n601 585
R277 B.n603 B.n0 585
R278 B.n2 B.n1 585
R279 B.n159 B.n158 585
R280 B.n161 B.n160 585
R281 B.n162 B.n157 585
R282 B.n164 B.n163 585
R283 B.n165 B.n156 585
R284 B.n167 B.n166 585
R285 B.n168 B.n155 585
R286 B.n170 B.n169 585
R287 B.n171 B.n154 585
R288 B.n173 B.n172 585
R289 B.n174 B.n153 585
R290 B.n176 B.n175 585
R291 B.n177 B.n152 585
R292 B.n179 B.n178 585
R293 B.n180 B.n151 585
R294 B.n182 B.n181 585
R295 B.n183 B.n150 585
R296 B.n185 B.n184 585
R297 B.n186 B.n149 585
R298 B.n188 B.n187 585
R299 B.n189 B.n148 585
R300 B.n191 B.n190 585
R301 B.n192 B.n147 585
R302 B.n194 B.n193 585
R303 B.n195 B.n146 585
R304 B.n197 B.n196 585
R305 B.n198 B.n145 585
R306 B.n200 B.n199 585
R307 B.n201 B.n144 585
R308 B.n203 B.n202 585
R309 B.n204 B.n143 585
R310 B.n205 B.n204 540.549
R311 B.n332 B.n331 540.549
R312 B.n429 B.n64 540.549
R313 B.n556 B.n555 540.549
R314 B.n123 B.t3 274.457
R315 B.n117 B.t6 274.457
R316 B.n45 B.t9 274.457
R317 B.n38 B.t0 274.457
R318 B.n605 B.n604 256.663
R319 B.n604 B.n603 235.042
R320 B.n604 B.n2 235.042
R321 B.n117 B.t7 191.72
R322 B.n45 B.t11 191.72
R323 B.n123 B.t4 191.708
R324 B.n38 B.t2 191.708
R325 B.n205 B.n142 163.367
R326 B.n209 B.n142 163.367
R327 B.n210 B.n209 163.367
R328 B.n211 B.n210 163.367
R329 B.n211 B.n140 163.367
R330 B.n215 B.n140 163.367
R331 B.n216 B.n215 163.367
R332 B.n217 B.n216 163.367
R333 B.n217 B.n138 163.367
R334 B.n221 B.n138 163.367
R335 B.n222 B.n221 163.367
R336 B.n223 B.n222 163.367
R337 B.n223 B.n136 163.367
R338 B.n227 B.n136 163.367
R339 B.n228 B.n227 163.367
R340 B.n229 B.n228 163.367
R341 B.n229 B.n134 163.367
R342 B.n233 B.n134 163.367
R343 B.n234 B.n233 163.367
R344 B.n235 B.n234 163.367
R345 B.n235 B.n132 163.367
R346 B.n239 B.n132 163.367
R347 B.n240 B.n239 163.367
R348 B.n241 B.n240 163.367
R349 B.n241 B.n130 163.367
R350 B.n245 B.n130 163.367
R351 B.n246 B.n245 163.367
R352 B.n247 B.n246 163.367
R353 B.n247 B.n128 163.367
R354 B.n251 B.n128 163.367
R355 B.n252 B.n251 163.367
R356 B.n253 B.n252 163.367
R357 B.n253 B.n126 163.367
R358 B.n257 B.n126 163.367
R359 B.n258 B.n257 163.367
R360 B.n259 B.n258 163.367
R361 B.n259 B.n122 163.367
R362 B.n264 B.n122 163.367
R363 B.n265 B.n264 163.367
R364 B.n266 B.n265 163.367
R365 B.n266 B.n120 163.367
R366 B.n270 B.n120 163.367
R367 B.n271 B.n270 163.367
R368 B.n272 B.n271 163.367
R369 B.n272 B.n116 163.367
R370 B.n277 B.n116 163.367
R371 B.n278 B.n277 163.367
R372 B.n279 B.n278 163.367
R373 B.n279 B.n114 163.367
R374 B.n283 B.n114 163.367
R375 B.n284 B.n283 163.367
R376 B.n285 B.n284 163.367
R377 B.n285 B.n112 163.367
R378 B.n289 B.n112 163.367
R379 B.n290 B.n289 163.367
R380 B.n291 B.n290 163.367
R381 B.n291 B.n110 163.367
R382 B.n295 B.n110 163.367
R383 B.n296 B.n295 163.367
R384 B.n297 B.n296 163.367
R385 B.n297 B.n108 163.367
R386 B.n301 B.n108 163.367
R387 B.n302 B.n301 163.367
R388 B.n303 B.n302 163.367
R389 B.n303 B.n106 163.367
R390 B.n307 B.n106 163.367
R391 B.n308 B.n307 163.367
R392 B.n309 B.n308 163.367
R393 B.n309 B.n104 163.367
R394 B.n313 B.n104 163.367
R395 B.n314 B.n313 163.367
R396 B.n315 B.n314 163.367
R397 B.n315 B.n102 163.367
R398 B.n319 B.n102 163.367
R399 B.n320 B.n319 163.367
R400 B.n321 B.n320 163.367
R401 B.n321 B.n100 163.367
R402 B.n325 B.n100 163.367
R403 B.n326 B.n325 163.367
R404 B.n327 B.n326 163.367
R405 B.n327 B.n98 163.367
R406 B.n331 B.n98 163.367
R407 B.n429 B.n428 163.367
R408 B.n428 B.n427 163.367
R409 B.n427 B.n66 163.367
R410 B.n423 B.n66 163.367
R411 B.n423 B.n422 163.367
R412 B.n422 B.n421 163.367
R413 B.n421 B.n68 163.367
R414 B.n417 B.n68 163.367
R415 B.n417 B.n416 163.367
R416 B.n416 B.n415 163.367
R417 B.n415 B.n70 163.367
R418 B.n411 B.n70 163.367
R419 B.n411 B.n410 163.367
R420 B.n410 B.n409 163.367
R421 B.n409 B.n72 163.367
R422 B.n405 B.n72 163.367
R423 B.n405 B.n404 163.367
R424 B.n404 B.n403 163.367
R425 B.n403 B.n74 163.367
R426 B.n399 B.n74 163.367
R427 B.n399 B.n398 163.367
R428 B.n398 B.n397 163.367
R429 B.n397 B.n76 163.367
R430 B.n393 B.n76 163.367
R431 B.n393 B.n392 163.367
R432 B.n392 B.n391 163.367
R433 B.n391 B.n78 163.367
R434 B.n387 B.n78 163.367
R435 B.n387 B.n386 163.367
R436 B.n386 B.n385 163.367
R437 B.n385 B.n80 163.367
R438 B.n381 B.n80 163.367
R439 B.n381 B.n380 163.367
R440 B.n380 B.n379 163.367
R441 B.n379 B.n82 163.367
R442 B.n375 B.n82 163.367
R443 B.n375 B.n374 163.367
R444 B.n374 B.n373 163.367
R445 B.n373 B.n84 163.367
R446 B.n369 B.n84 163.367
R447 B.n369 B.n368 163.367
R448 B.n368 B.n367 163.367
R449 B.n367 B.n86 163.367
R450 B.n363 B.n86 163.367
R451 B.n363 B.n362 163.367
R452 B.n362 B.n361 163.367
R453 B.n361 B.n88 163.367
R454 B.n357 B.n88 163.367
R455 B.n357 B.n356 163.367
R456 B.n356 B.n355 163.367
R457 B.n355 B.n90 163.367
R458 B.n351 B.n90 163.367
R459 B.n351 B.n350 163.367
R460 B.n350 B.n349 163.367
R461 B.n349 B.n92 163.367
R462 B.n345 B.n92 163.367
R463 B.n345 B.n344 163.367
R464 B.n344 B.n343 163.367
R465 B.n343 B.n94 163.367
R466 B.n339 B.n94 163.367
R467 B.n339 B.n338 163.367
R468 B.n338 B.n337 163.367
R469 B.n337 B.n96 163.367
R470 B.n333 B.n96 163.367
R471 B.n333 B.n332 163.367
R472 B.n555 B.n554 163.367
R473 B.n554 B.n19 163.367
R474 B.n550 B.n19 163.367
R475 B.n550 B.n549 163.367
R476 B.n549 B.n548 163.367
R477 B.n548 B.n21 163.367
R478 B.n544 B.n21 163.367
R479 B.n544 B.n543 163.367
R480 B.n543 B.n542 163.367
R481 B.n542 B.n23 163.367
R482 B.n538 B.n23 163.367
R483 B.n538 B.n537 163.367
R484 B.n537 B.n536 163.367
R485 B.n536 B.n25 163.367
R486 B.n532 B.n25 163.367
R487 B.n532 B.n531 163.367
R488 B.n531 B.n530 163.367
R489 B.n530 B.n27 163.367
R490 B.n526 B.n27 163.367
R491 B.n526 B.n525 163.367
R492 B.n525 B.n524 163.367
R493 B.n524 B.n29 163.367
R494 B.n520 B.n29 163.367
R495 B.n520 B.n519 163.367
R496 B.n519 B.n518 163.367
R497 B.n518 B.n31 163.367
R498 B.n514 B.n31 163.367
R499 B.n514 B.n513 163.367
R500 B.n513 B.n512 163.367
R501 B.n512 B.n33 163.367
R502 B.n508 B.n33 163.367
R503 B.n508 B.n507 163.367
R504 B.n507 B.n506 163.367
R505 B.n506 B.n35 163.367
R506 B.n502 B.n35 163.367
R507 B.n502 B.n501 163.367
R508 B.n501 B.n500 163.367
R509 B.n500 B.n37 163.367
R510 B.n496 B.n37 163.367
R511 B.n496 B.n495 163.367
R512 B.n495 B.n494 163.367
R513 B.n494 B.n42 163.367
R514 B.n490 B.n42 163.367
R515 B.n490 B.n489 163.367
R516 B.n489 B.n488 163.367
R517 B.n488 B.n44 163.367
R518 B.n483 B.n44 163.367
R519 B.n483 B.n482 163.367
R520 B.n482 B.n481 163.367
R521 B.n481 B.n48 163.367
R522 B.n477 B.n48 163.367
R523 B.n477 B.n476 163.367
R524 B.n476 B.n475 163.367
R525 B.n475 B.n50 163.367
R526 B.n471 B.n50 163.367
R527 B.n471 B.n470 163.367
R528 B.n470 B.n469 163.367
R529 B.n469 B.n52 163.367
R530 B.n465 B.n52 163.367
R531 B.n465 B.n464 163.367
R532 B.n464 B.n463 163.367
R533 B.n463 B.n54 163.367
R534 B.n459 B.n54 163.367
R535 B.n459 B.n458 163.367
R536 B.n458 B.n457 163.367
R537 B.n457 B.n56 163.367
R538 B.n453 B.n56 163.367
R539 B.n453 B.n452 163.367
R540 B.n452 B.n451 163.367
R541 B.n451 B.n58 163.367
R542 B.n447 B.n58 163.367
R543 B.n447 B.n446 163.367
R544 B.n446 B.n445 163.367
R545 B.n445 B.n60 163.367
R546 B.n441 B.n60 163.367
R547 B.n441 B.n440 163.367
R548 B.n440 B.n439 163.367
R549 B.n439 B.n62 163.367
R550 B.n435 B.n62 163.367
R551 B.n435 B.n434 163.367
R552 B.n434 B.n433 163.367
R553 B.n433 B.n64 163.367
R554 B.n556 B.n17 163.367
R555 B.n560 B.n17 163.367
R556 B.n561 B.n560 163.367
R557 B.n562 B.n561 163.367
R558 B.n562 B.n15 163.367
R559 B.n566 B.n15 163.367
R560 B.n567 B.n566 163.367
R561 B.n568 B.n567 163.367
R562 B.n568 B.n13 163.367
R563 B.n572 B.n13 163.367
R564 B.n573 B.n572 163.367
R565 B.n574 B.n573 163.367
R566 B.n574 B.n11 163.367
R567 B.n578 B.n11 163.367
R568 B.n579 B.n578 163.367
R569 B.n580 B.n579 163.367
R570 B.n580 B.n9 163.367
R571 B.n584 B.n9 163.367
R572 B.n585 B.n584 163.367
R573 B.n586 B.n585 163.367
R574 B.n586 B.n7 163.367
R575 B.n590 B.n7 163.367
R576 B.n591 B.n590 163.367
R577 B.n592 B.n591 163.367
R578 B.n592 B.n5 163.367
R579 B.n596 B.n5 163.367
R580 B.n597 B.n596 163.367
R581 B.n598 B.n597 163.367
R582 B.n598 B.n3 163.367
R583 B.n602 B.n3 163.367
R584 B.n603 B.n602 163.367
R585 B.n158 B.n2 163.367
R586 B.n161 B.n158 163.367
R587 B.n162 B.n161 163.367
R588 B.n163 B.n162 163.367
R589 B.n163 B.n156 163.367
R590 B.n167 B.n156 163.367
R591 B.n168 B.n167 163.367
R592 B.n169 B.n168 163.367
R593 B.n169 B.n154 163.367
R594 B.n173 B.n154 163.367
R595 B.n174 B.n173 163.367
R596 B.n175 B.n174 163.367
R597 B.n175 B.n152 163.367
R598 B.n179 B.n152 163.367
R599 B.n180 B.n179 163.367
R600 B.n181 B.n180 163.367
R601 B.n181 B.n150 163.367
R602 B.n185 B.n150 163.367
R603 B.n186 B.n185 163.367
R604 B.n187 B.n186 163.367
R605 B.n187 B.n148 163.367
R606 B.n191 B.n148 163.367
R607 B.n192 B.n191 163.367
R608 B.n193 B.n192 163.367
R609 B.n193 B.n146 163.367
R610 B.n197 B.n146 163.367
R611 B.n198 B.n197 163.367
R612 B.n199 B.n198 163.367
R613 B.n199 B.n144 163.367
R614 B.n203 B.n144 163.367
R615 B.n204 B.n203 163.367
R616 B.n118 B.t8 110.847
R617 B.n46 B.t10 110.847
R618 B.n124 B.t5 110.835
R619 B.n39 B.t1 110.835
R620 B.n124 B.n123 80.8732
R621 B.n118 B.n117 80.8732
R622 B.n46 B.n45 80.8732
R623 B.n39 B.n38 80.8732
R624 B.n261 B.n124 59.5399
R625 B.n275 B.n118 59.5399
R626 B.n486 B.n46 59.5399
R627 B.n40 B.n39 59.5399
R628 B.n557 B.n18 35.1225
R629 B.n431 B.n430 35.1225
R630 B.n330 B.n97 35.1225
R631 B.n206 B.n143 35.1225
R632 B B.n605 18.0485
R633 B.n558 B.n557 10.6151
R634 B.n559 B.n558 10.6151
R635 B.n559 B.n16 10.6151
R636 B.n563 B.n16 10.6151
R637 B.n564 B.n563 10.6151
R638 B.n565 B.n564 10.6151
R639 B.n565 B.n14 10.6151
R640 B.n569 B.n14 10.6151
R641 B.n570 B.n569 10.6151
R642 B.n571 B.n570 10.6151
R643 B.n571 B.n12 10.6151
R644 B.n575 B.n12 10.6151
R645 B.n576 B.n575 10.6151
R646 B.n577 B.n576 10.6151
R647 B.n577 B.n10 10.6151
R648 B.n581 B.n10 10.6151
R649 B.n582 B.n581 10.6151
R650 B.n583 B.n582 10.6151
R651 B.n583 B.n8 10.6151
R652 B.n587 B.n8 10.6151
R653 B.n588 B.n587 10.6151
R654 B.n589 B.n588 10.6151
R655 B.n589 B.n6 10.6151
R656 B.n593 B.n6 10.6151
R657 B.n594 B.n593 10.6151
R658 B.n595 B.n594 10.6151
R659 B.n595 B.n4 10.6151
R660 B.n599 B.n4 10.6151
R661 B.n600 B.n599 10.6151
R662 B.n601 B.n600 10.6151
R663 B.n601 B.n0 10.6151
R664 B.n553 B.n18 10.6151
R665 B.n553 B.n552 10.6151
R666 B.n552 B.n551 10.6151
R667 B.n551 B.n20 10.6151
R668 B.n547 B.n20 10.6151
R669 B.n547 B.n546 10.6151
R670 B.n546 B.n545 10.6151
R671 B.n545 B.n22 10.6151
R672 B.n541 B.n22 10.6151
R673 B.n541 B.n540 10.6151
R674 B.n540 B.n539 10.6151
R675 B.n539 B.n24 10.6151
R676 B.n535 B.n24 10.6151
R677 B.n535 B.n534 10.6151
R678 B.n534 B.n533 10.6151
R679 B.n533 B.n26 10.6151
R680 B.n529 B.n26 10.6151
R681 B.n529 B.n528 10.6151
R682 B.n528 B.n527 10.6151
R683 B.n527 B.n28 10.6151
R684 B.n523 B.n28 10.6151
R685 B.n523 B.n522 10.6151
R686 B.n522 B.n521 10.6151
R687 B.n521 B.n30 10.6151
R688 B.n517 B.n30 10.6151
R689 B.n517 B.n516 10.6151
R690 B.n516 B.n515 10.6151
R691 B.n515 B.n32 10.6151
R692 B.n511 B.n32 10.6151
R693 B.n511 B.n510 10.6151
R694 B.n510 B.n509 10.6151
R695 B.n509 B.n34 10.6151
R696 B.n505 B.n34 10.6151
R697 B.n505 B.n504 10.6151
R698 B.n504 B.n503 10.6151
R699 B.n503 B.n36 10.6151
R700 B.n499 B.n498 10.6151
R701 B.n498 B.n497 10.6151
R702 B.n497 B.n41 10.6151
R703 B.n493 B.n41 10.6151
R704 B.n493 B.n492 10.6151
R705 B.n492 B.n491 10.6151
R706 B.n491 B.n43 10.6151
R707 B.n487 B.n43 10.6151
R708 B.n485 B.n484 10.6151
R709 B.n484 B.n47 10.6151
R710 B.n480 B.n47 10.6151
R711 B.n480 B.n479 10.6151
R712 B.n479 B.n478 10.6151
R713 B.n478 B.n49 10.6151
R714 B.n474 B.n49 10.6151
R715 B.n474 B.n473 10.6151
R716 B.n473 B.n472 10.6151
R717 B.n472 B.n51 10.6151
R718 B.n468 B.n51 10.6151
R719 B.n468 B.n467 10.6151
R720 B.n467 B.n466 10.6151
R721 B.n466 B.n53 10.6151
R722 B.n462 B.n53 10.6151
R723 B.n462 B.n461 10.6151
R724 B.n461 B.n460 10.6151
R725 B.n460 B.n55 10.6151
R726 B.n456 B.n55 10.6151
R727 B.n456 B.n455 10.6151
R728 B.n455 B.n454 10.6151
R729 B.n454 B.n57 10.6151
R730 B.n450 B.n57 10.6151
R731 B.n450 B.n449 10.6151
R732 B.n449 B.n448 10.6151
R733 B.n448 B.n59 10.6151
R734 B.n444 B.n59 10.6151
R735 B.n444 B.n443 10.6151
R736 B.n443 B.n442 10.6151
R737 B.n442 B.n61 10.6151
R738 B.n438 B.n61 10.6151
R739 B.n438 B.n437 10.6151
R740 B.n437 B.n436 10.6151
R741 B.n436 B.n63 10.6151
R742 B.n432 B.n63 10.6151
R743 B.n432 B.n431 10.6151
R744 B.n430 B.n65 10.6151
R745 B.n426 B.n65 10.6151
R746 B.n426 B.n425 10.6151
R747 B.n425 B.n424 10.6151
R748 B.n424 B.n67 10.6151
R749 B.n420 B.n67 10.6151
R750 B.n420 B.n419 10.6151
R751 B.n419 B.n418 10.6151
R752 B.n418 B.n69 10.6151
R753 B.n414 B.n69 10.6151
R754 B.n414 B.n413 10.6151
R755 B.n413 B.n412 10.6151
R756 B.n412 B.n71 10.6151
R757 B.n408 B.n71 10.6151
R758 B.n408 B.n407 10.6151
R759 B.n407 B.n406 10.6151
R760 B.n406 B.n73 10.6151
R761 B.n402 B.n73 10.6151
R762 B.n402 B.n401 10.6151
R763 B.n401 B.n400 10.6151
R764 B.n400 B.n75 10.6151
R765 B.n396 B.n75 10.6151
R766 B.n396 B.n395 10.6151
R767 B.n395 B.n394 10.6151
R768 B.n394 B.n77 10.6151
R769 B.n390 B.n77 10.6151
R770 B.n390 B.n389 10.6151
R771 B.n389 B.n388 10.6151
R772 B.n388 B.n79 10.6151
R773 B.n384 B.n79 10.6151
R774 B.n384 B.n383 10.6151
R775 B.n383 B.n382 10.6151
R776 B.n382 B.n81 10.6151
R777 B.n378 B.n81 10.6151
R778 B.n378 B.n377 10.6151
R779 B.n377 B.n376 10.6151
R780 B.n376 B.n83 10.6151
R781 B.n372 B.n83 10.6151
R782 B.n372 B.n371 10.6151
R783 B.n371 B.n370 10.6151
R784 B.n370 B.n85 10.6151
R785 B.n366 B.n85 10.6151
R786 B.n366 B.n365 10.6151
R787 B.n365 B.n364 10.6151
R788 B.n364 B.n87 10.6151
R789 B.n360 B.n87 10.6151
R790 B.n360 B.n359 10.6151
R791 B.n359 B.n358 10.6151
R792 B.n358 B.n89 10.6151
R793 B.n354 B.n89 10.6151
R794 B.n354 B.n353 10.6151
R795 B.n353 B.n352 10.6151
R796 B.n352 B.n91 10.6151
R797 B.n348 B.n91 10.6151
R798 B.n348 B.n347 10.6151
R799 B.n347 B.n346 10.6151
R800 B.n346 B.n93 10.6151
R801 B.n342 B.n93 10.6151
R802 B.n342 B.n341 10.6151
R803 B.n341 B.n340 10.6151
R804 B.n340 B.n95 10.6151
R805 B.n336 B.n95 10.6151
R806 B.n336 B.n335 10.6151
R807 B.n335 B.n334 10.6151
R808 B.n334 B.n97 10.6151
R809 B.n159 B.n1 10.6151
R810 B.n160 B.n159 10.6151
R811 B.n160 B.n157 10.6151
R812 B.n164 B.n157 10.6151
R813 B.n165 B.n164 10.6151
R814 B.n166 B.n165 10.6151
R815 B.n166 B.n155 10.6151
R816 B.n170 B.n155 10.6151
R817 B.n171 B.n170 10.6151
R818 B.n172 B.n171 10.6151
R819 B.n172 B.n153 10.6151
R820 B.n176 B.n153 10.6151
R821 B.n177 B.n176 10.6151
R822 B.n178 B.n177 10.6151
R823 B.n178 B.n151 10.6151
R824 B.n182 B.n151 10.6151
R825 B.n183 B.n182 10.6151
R826 B.n184 B.n183 10.6151
R827 B.n184 B.n149 10.6151
R828 B.n188 B.n149 10.6151
R829 B.n189 B.n188 10.6151
R830 B.n190 B.n189 10.6151
R831 B.n190 B.n147 10.6151
R832 B.n194 B.n147 10.6151
R833 B.n195 B.n194 10.6151
R834 B.n196 B.n195 10.6151
R835 B.n196 B.n145 10.6151
R836 B.n200 B.n145 10.6151
R837 B.n201 B.n200 10.6151
R838 B.n202 B.n201 10.6151
R839 B.n202 B.n143 10.6151
R840 B.n207 B.n206 10.6151
R841 B.n208 B.n207 10.6151
R842 B.n208 B.n141 10.6151
R843 B.n212 B.n141 10.6151
R844 B.n213 B.n212 10.6151
R845 B.n214 B.n213 10.6151
R846 B.n214 B.n139 10.6151
R847 B.n218 B.n139 10.6151
R848 B.n219 B.n218 10.6151
R849 B.n220 B.n219 10.6151
R850 B.n220 B.n137 10.6151
R851 B.n224 B.n137 10.6151
R852 B.n225 B.n224 10.6151
R853 B.n226 B.n225 10.6151
R854 B.n226 B.n135 10.6151
R855 B.n230 B.n135 10.6151
R856 B.n231 B.n230 10.6151
R857 B.n232 B.n231 10.6151
R858 B.n232 B.n133 10.6151
R859 B.n236 B.n133 10.6151
R860 B.n237 B.n236 10.6151
R861 B.n238 B.n237 10.6151
R862 B.n238 B.n131 10.6151
R863 B.n242 B.n131 10.6151
R864 B.n243 B.n242 10.6151
R865 B.n244 B.n243 10.6151
R866 B.n244 B.n129 10.6151
R867 B.n248 B.n129 10.6151
R868 B.n249 B.n248 10.6151
R869 B.n250 B.n249 10.6151
R870 B.n250 B.n127 10.6151
R871 B.n254 B.n127 10.6151
R872 B.n255 B.n254 10.6151
R873 B.n256 B.n255 10.6151
R874 B.n256 B.n125 10.6151
R875 B.n260 B.n125 10.6151
R876 B.n263 B.n262 10.6151
R877 B.n263 B.n121 10.6151
R878 B.n267 B.n121 10.6151
R879 B.n268 B.n267 10.6151
R880 B.n269 B.n268 10.6151
R881 B.n269 B.n119 10.6151
R882 B.n273 B.n119 10.6151
R883 B.n274 B.n273 10.6151
R884 B.n276 B.n115 10.6151
R885 B.n280 B.n115 10.6151
R886 B.n281 B.n280 10.6151
R887 B.n282 B.n281 10.6151
R888 B.n282 B.n113 10.6151
R889 B.n286 B.n113 10.6151
R890 B.n287 B.n286 10.6151
R891 B.n288 B.n287 10.6151
R892 B.n288 B.n111 10.6151
R893 B.n292 B.n111 10.6151
R894 B.n293 B.n292 10.6151
R895 B.n294 B.n293 10.6151
R896 B.n294 B.n109 10.6151
R897 B.n298 B.n109 10.6151
R898 B.n299 B.n298 10.6151
R899 B.n300 B.n299 10.6151
R900 B.n300 B.n107 10.6151
R901 B.n304 B.n107 10.6151
R902 B.n305 B.n304 10.6151
R903 B.n306 B.n305 10.6151
R904 B.n306 B.n105 10.6151
R905 B.n310 B.n105 10.6151
R906 B.n311 B.n310 10.6151
R907 B.n312 B.n311 10.6151
R908 B.n312 B.n103 10.6151
R909 B.n316 B.n103 10.6151
R910 B.n317 B.n316 10.6151
R911 B.n318 B.n317 10.6151
R912 B.n318 B.n101 10.6151
R913 B.n322 B.n101 10.6151
R914 B.n323 B.n322 10.6151
R915 B.n324 B.n323 10.6151
R916 B.n324 B.n99 10.6151
R917 B.n328 B.n99 10.6151
R918 B.n329 B.n328 10.6151
R919 B.n330 B.n329 10.6151
R920 B.n605 B.n0 8.11757
R921 B.n605 B.n1 8.11757
R922 B.n499 B.n40 6.5566
R923 B.n487 B.n486 6.5566
R924 B.n262 B.n261 6.5566
R925 B.n275 B.n274 6.5566
R926 B.n40 B.n36 4.05904
R927 B.n486 B.n485 4.05904
R928 B.n261 B.n260 4.05904
R929 B.n276 B.n275 4.05904
R930 VN VN.t1 146.643
R931 VN VN.t0 100.74
R932 VDD2.n0 VDD2.t1 120.362
R933 VDD2.n0 VDD2.t0 80.5727
R934 VDD2 VDD2.n0 0.957397
C0 VDD2 B 1.77776f
C1 VN VTAIL 2.3824f
C2 VDD1 VP 2.79604f
C3 VN w_n2638_n3042# 3.73345f
C4 B VP 1.80094f
C5 VTAIL w_n2638_n3042# 2.55884f
C6 VDD2 VP 0.384592f
C7 VDD1 VN 0.148692f
C8 VDD1 VTAIL 4.91811f
C9 B VN 1.23912f
C10 VDD1 w_n2638_n3042# 1.80739f
C11 B VTAIL 3.71465f
C12 VDD2 VN 2.56151f
C13 B w_n2638_n3042# 9.691549f
C14 VDD2 VTAIL 4.97827f
C15 VDD2 w_n2638_n3042# 1.84854f
C16 VN VP 5.73735f
C17 VDD1 B 1.73654f
C18 VTAIL VP 2.3971f
C19 VDD2 VDD1 0.812915f
C20 VP w_n2638_n3042# 4.07215f
C21 VDD2 VSUBS 0.965426f
C22 VDD1 VSUBS 4.76674f
C23 VTAIL VSUBS 1.068127f
C24 VN VSUBS 7.97304f
C25 VP VSUBS 2.0037f
C26 B VSUBS 4.680101f
C27 w_n2638_n3042# VSUBS 99.0516f
C28 VDD2.t1 VSUBS 2.27031f
C29 VDD2.t0 VSUBS 1.70406f
C30 VDD2.n0 VSUBS 3.44012f
C31 VN.t0 VSUBS 4.18881f
C32 VN.t1 VSUBS 5.12724f
C33 B.n0 VSUBS 0.005242f
C34 B.n1 VSUBS 0.005242f
C35 B.n2 VSUBS 0.007752f
C36 B.n3 VSUBS 0.005941f
C37 B.n4 VSUBS 0.005941f
C38 B.n5 VSUBS 0.005941f
C39 B.n6 VSUBS 0.005941f
C40 B.n7 VSUBS 0.005941f
C41 B.n8 VSUBS 0.005941f
C42 B.n9 VSUBS 0.005941f
C43 B.n10 VSUBS 0.005941f
C44 B.n11 VSUBS 0.005941f
C45 B.n12 VSUBS 0.005941f
C46 B.n13 VSUBS 0.005941f
C47 B.n14 VSUBS 0.005941f
C48 B.n15 VSUBS 0.005941f
C49 B.n16 VSUBS 0.005941f
C50 B.n17 VSUBS 0.005941f
C51 B.n18 VSUBS 0.014916f
C52 B.n19 VSUBS 0.005941f
C53 B.n20 VSUBS 0.005941f
C54 B.n21 VSUBS 0.005941f
C55 B.n22 VSUBS 0.005941f
C56 B.n23 VSUBS 0.005941f
C57 B.n24 VSUBS 0.005941f
C58 B.n25 VSUBS 0.005941f
C59 B.n26 VSUBS 0.005941f
C60 B.n27 VSUBS 0.005941f
C61 B.n28 VSUBS 0.005941f
C62 B.n29 VSUBS 0.005941f
C63 B.n30 VSUBS 0.005941f
C64 B.n31 VSUBS 0.005941f
C65 B.n32 VSUBS 0.005941f
C66 B.n33 VSUBS 0.005941f
C67 B.n34 VSUBS 0.005941f
C68 B.n35 VSUBS 0.005941f
C69 B.n36 VSUBS 0.004106f
C70 B.n37 VSUBS 0.005941f
C71 B.t1 VSUBS 0.281979f
C72 B.t2 VSUBS 0.3059f
C73 B.t0 VSUBS 1.58865f
C74 B.n38 VSUBS 0.175092f
C75 B.n39 VSUBS 0.065177f
C76 B.n40 VSUBS 0.013764f
C77 B.n41 VSUBS 0.005941f
C78 B.n42 VSUBS 0.005941f
C79 B.n43 VSUBS 0.005941f
C80 B.n44 VSUBS 0.005941f
C81 B.t10 VSUBS 0.281975f
C82 B.t11 VSUBS 0.305896f
C83 B.t9 VSUBS 1.58865f
C84 B.n45 VSUBS 0.175096f
C85 B.n46 VSUBS 0.065181f
C86 B.n47 VSUBS 0.005941f
C87 B.n48 VSUBS 0.005941f
C88 B.n49 VSUBS 0.005941f
C89 B.n50 VSUBS 0.005941f
C90 B.n51 VSUBS 0.005941f
C91 B.n52 VSUBS 0.005941f
C92 B.n53 VSUBS 0.005941f
C93 B.n54 VSUBS 0.005941f
C94 B.n55 VSUBS 0.005941f
C95 B.n56 VSUBS 0.005941f
C96 B.n57 VSUBS 0.005941f
C97 B.n58 VSUBS 0.005941f
C98 B.n59 VSUBS 0.005941f
C99 B.n60 VSUBS 0.005941f
C100 B.n61 VSUBS 0.005941f
C101 B.n62 VSUBS 0.005941f
C102 B.n63 VSUBS 0.005941f
C103 B.n64 VSUBS 0.014916f
C104 B.n65 VSUBS 0.005941f
C105 B.n66 VSUBS 0.005941f
C106 B.n67 VSUBS 0.005941f
C107 B.n68 VSUBS 0.005941f
C108 B.n69 VSUBS 0.005941f
C109 B.n70 VSUBS 0.005941f
C110 B.n71 VSUBS 0.005941f
C111 B.n72 VSUBS 0.005941f
C112 B.n73 VSUBS 0.005941f
C113 B.n74 VSUBS 0.005941f
C114 B.n75 VSUBS 0.005941f
C115 B.n76 VSUBS 0.005941f
C116 B.n77 VSUBS 0.005941f
C117 B.n78 VSUBS 0.005941f
C118 B.n79 VSUBS 0.005941f
C119 B.n80 VSUBS 0.005941f
C120 B.n81 VSUBS 0.005941f
C121 B.n82 VSUBS 0.005941f
C122 B.n83 VSUBS 0.005941f
C123 B.n84 VSUBS 0.005941f
C124 B.n85 VSUBS 0.005941f
C125 B.n86 VSUBS 0.005941f
C126 B.n87 VSUBS 0.005941f
C127 B.n88 VSUBS 0.005941f
C128 B.n89 VSUBS 0.005941f
C129 B.n90 VSUBS 0.005941f
C130 B.n91 VSUBS 0.005941f
C131 B.n92 VSUBS 0.005941f
C132 B.n93 VSUBS 0.005941f
C133 B.n94 VSUBS 0.005941f
C134 B.n95 VSUBS 0.005941f
C135 B.n96 VSUBS 0.005941f
C136 B.n97 VSUBS 0.014916f
C137 B.n98 VSUBS 0.005941f
C138 B.n99 VSUBS 0.005941f
C139 B.n100 VSUBS 0.005941f
C140 B.n101 VSUBS 0.005941f
C141 B.n102 VSUBS 0.005941f
C142 B.n103 VSUBS 0.005941f
C143 B.n104 VSUBS 0.005941f
C144 B.n105 VSUBS 0.005941f
C145 B.n106 VSUBS 0.005941f
C146 B.n107 VSUBS 0.005941f
C147 B.n108 VSUBS 0.005941f
C148 B.n109 VSUBS 0.005941f
C149 B.n110 VSUBS 0.005941f
C150 B.n111 VSUBS 0.005941f
C151 B.n112 VSUBS 0.005941f
C152 B.n113 VSUBS 0.005941f
C153 B.n114 VSUBS 0.005941f
C154 B.n115 VSUBS 0.005941f
C155 B.n116 VSUBS 0.005941f
C156 B.t8 VSUBS 0.281975f
C157 B.t7 VSUBS 0.305896f
C158 B.t6 VSUBS 1.58865f
C159 B.n117 VSUBS 0.175096f
C160 B.n118 VSUBS 0.065181f
C161 B.n119 VSUBS 0.005941f
C162 B.n120 VSUBS 0.005941f
C163 B.n121 VSUBS 0.005941f
C164 B.n122 VSUBS 0.005941f
C165 B.t5 VSUBS 0.281979f
C166 B.t4 VSUBS 0.3059f
C167 B.t3 VSUBS 1.58865f
C168 B.n123 VSUBS 0.175092f
C169 B.n124 VSUBS 0.065177f
C170 B.n125 VSUBS 0.005941f
C171 B.n126 VSUBS 0.005941f
C172 B.n127 VSUBS 0.005941f
C173 B.n128 VSUBS 0.005941f
C174 B.n129 VSUBS 0.005941f
C175 B.n130 VSUBS 0.005941f
C176 B.n131 VSUBS 0.005941f
C177 B.n132 VSUBS 0.005941f
C178 B.n133 VSUBS 0.005941f
C179 B.n134 VSUBS 0.005941f
C180 B.n135 VSUBS 0.005941f
C181 B.n136 VSUBS 0.005941f
C182 B.n137 VSUBS 0.005941f
C183 B.n138 VSUBS 0.005941f
C184 B.n139 VSUBS 0.005941f
C185 B.n140 VSUBS 0.005941f
C186 B.n141 VSUBS 0.005941f
C187 B.n142 VSUBS 0.005941f
C188 B.n143 VSUBS 0.014263f
C189 B.n144 VSUBS 0.005941f
C190 B.n145 VSUBS 0.005941f
C191 B.n146 VSUBS 0.005941f
C192 B.n147 VSUBS 0.005941f
C193 B.n148 VSUBS 0.005941f
C194 B.n149 VSUBS 0.005941f
C195 B.n150 VSUBS 0.005941f
C196 B.n151 VSUBS 0.005941f
C197 B.n152 VSUBS 0.005941f
C198 B.n153 VSUBS 0.005941f
C199 B.n154 VSUBS 0.005941f
C200 B.n155 VSUBS 0.005941f
C201 B.n156 VSUBS 0.005941f
C202 B.n157 VSUBS 0.005941f
C203 B.n158 VSUBS 0.005941f
C204 B.n159 VSUBS 0.005941f
C205 B.n160 VSUBS 0.005941f
C206 B.n161 VSUBS 0.005941f
C207 B.n162 VSUBS 0.005941f
C208 B.n163 VSUBS 0.005941f
C209 B.n164 VSUBS 0.005941f
C210 B.n165 VSUBS 0.005941f
C211 B.n166 VSUBS 0.005941f
C212 B.n167 VSUBS 0.005941f
C213 B.n168 VSUBS 0.005941f
C214 B.n169 VSUBS 0.005941f
C215 B.n170 VSUBS 0.005941f
C216 B.n171 VSUBS 0.005941f
C217 B.n172 VSUBS 0.005941f
C218 B.n173 VSUBS 0.005941f
C219 B.n174 VSUBS 0.005941f
C220 B.n175 VSUBS 0.005941f
C221 B.n176 VSUBS 0.005941f
C222 B.n177 VSUBS 0.005941f
C223 B.n178 VSUBS 0.005941f
C224 B.n179 VSUBS 0.005941f
C225 B.n180 VSUBS 0.005941f
C226 B.n181 VSUBS 0.005941f
C227 B.n182 VSUBS 0.005941f
C228 B.n183 VSUBS 0.005941f
C229 B.n184 VSUBS 0.005941f
C230 B.n185 VSUBS 0.005941f
C231 B.n186 VSUBS 0.005941f
C232 B.n187 VSUBS 0.005941f
C233 B.n188 VSUBS 0.005941f
C234 B.n189 VSUBS 0.005941f
C235 B.n190 VSUBS 0.005941f
C236 B.n191 VSUBS 0.005941f
C237 B.n192 VSUBS 0.005941f
C238 B.n193 VSUBS 0.005941f
C239 B.n194 VSUBS 0.005941f
C240 B.n195 VSUBS 0.005941f
C241 B.n196 VSUBS 0.005941f
C242 B.n197 VSUBS 0.005941f
C243 B.n198 VSUBS 0.005941f
C244 B.n199 VSUBS 0.005941f
C245 B.n200 VSUBS 0.005941f
C246 B.n201 VSUBS 0.005941f
C247 B.n202 VSUBS 0.005941f
C248 B.n203 VSUBS 0.005941f
C249 B.n204 VSUBS 0.014263f
C250 B.n205 VSUBS 0.014916f
C251 B.n206 VSUBS 0.014916f
C252 B.n207 VSUBS 0.005941f
C253 B.n208 VSUBS 0.005941f
C254 B.n209 VSUBS 0.005941f
C255 B.n210 VSUBS 0.005941f
C256 B.n211 VSUBS 0.005941f
C257 B.n212 VSUBS 0.005941f
C258 B.n213 VSUBS 0.005941f
C259 B.n214 VSUBS 0.005941f
C260 B.n215 VSUBS 0.005941f
C261 B.n216 VSUBS 0.005941f
C262 B.n217 VSUBS 0.005941f
C263 B.n218 VSUBS 0.005941f
C264 B.n219 VSUBS 0.005941f
C265 B.n220 VSUBS 0.005941f
C266 B.n221 VSUBS 0.005941f
C267 B.n222 VSUBS 0.005941f
C268 B.n223 VSUBS 0.005941f
C269 B.n224 VSUBS 0.005941f
C270 B.n225 VSUBS 0.005941f
C271 B.n226 VSUBS 0.005941f
C272 B.n227 VSUBS 0.005941f
C273 B.n228 VSUBS 0.005941f
C274 B.n229 VSUBS 0.005941f
C275 B.n230 VSUBS 0.005941f
C276 B.n231 VSUBS 0.005941f
C277 B.n232 VSUBS 0.005941f
C278 B.n233 VSUBS 0.005941f
C279 B.n234 VSUBS 0.005941f
C280 B.n235 VSUBS 0.005941f
C281 B.n236 VSUBS 0.005941f
C282 B.n237 VSUBS 0.005941f
C283 B.n238 VSUBS 0.005941f
C284 B.n239 VSUBS 0.005941f
C285 B.n240 VSUBS 0.005941f
C286 B.n241 VSUBS 0.005941f
C287 B.n242 VSUBS 0.005941f
C288 B.n243 VSUBS 0.005941f
C289 B.n244 VSUBS 0.005941f
C290 B.n245 VSUBS 0.005941f
C291 B.n246 VSUBS 0.005941f
C292 B.n247 VSUBS 0.005941f
C293 B.n248 VSUBS 0.005941f
C294 B.n249 VSUBS 0.005941f
C295 B.n250 VSUBS 0.005941f
C296 B.n251 VSUBS 0.005941f
C297 B.n252 VSUBS 0.005941f
C298 B.n253 VSUBS 0.005941f
C299 B.n254 VSUBS 0.005941f
C300 B.n255 VSUBS 0.005941f
C301 B.n256 VSUBS 0.005941f
C302 B.n257 VSUBS 0.005941f
C303 B.n258 VSUBS 0.005941f
C304 B.n259 VSUBS 0.005941f
C305 B.n260 VSUBS 0.004106f
C306 B.n261 VSUBS 0.013764f
C307 B.n262 VSUBS 0.004805f
C308 B.n263 VSUBS 0.005941f
C309 B.n264 VSUBS 0.005941f
C310 B.n265 VSUBS 0.005941f
C311 B.n266 VSUBS 0.005941f
C312 B.n267 VSUBS 0.005941f
C313 B.n268 VSUBS 0.005941f
C314 B.n269 VSUBS 0.005941f
C315 B.n270 VSUBS 0.005941f
C316 B.n271 VSUBS 0.005941f
C317 B.n272 VSUBS 0.005941f
C318 B.n273 VSUBS 0.005941f
C319 B.n274 VSUBS 0.004805f
C320 B.n275 VSUBS 0.013764f
C321 B.n276 VSUBS 0.004106f
C322 B.n277 VSUBS 0.005941f
C323 B.n278 VSUBS 0.005941f
C324 B.n279 VSUBS 0.005941f
C325 B.n280 VSUBS 0.005941f
C326 B.n281 VSUBS 0.005941f
C327 B.n282 VSUBS 0.005941f
C328 B.n283 VSUBS 0.005941f
C329 B.n284 VSUBS 0.005941f
C330 B.n285 VSUBS 0.005941f
C331 B.n286 VSUBS 0.005941f
C332 B.n287 VSUBS 0.005941f
C333 B.n288 VSUBS 0.005941f
C334 B.n289 VSUBS 0.005941f
C335 B.n290 VSUBS 0.005941f
C336 B.n291 VSUBS 0.005941f
C337 B.n292 VSUBS 0.005941f
C338 B.n293 VSUBS 0.005941f
C339 B.n294 VSUBS 0.005941f
C340 B.n295 VSUBS 0.005941f
C341 B.n296 VSUBS 0.005941f
C342 B.n297 VSUBS 0.005941f
C343 B.n298 VSUBS 0.005941f
C344 B.n299 VSUBS 0.005941f
C345 B.n300 VSUBS 0.005941f
C346 B.n301 VSUBS 0.005941f
C347 B.n302 VSUBS 0.005941f
C348 B.n303 VSUBS 0.005941f
C349 B.n304 VSUBS 0.005941f
C350 B.n305 VSUBS 0.005941f
C351 B.n306 VSUBS 0.005941f
C352 B.n307 VSUBS 0.005941f
C353 B.n308 VSUBS 0.005941f
C354 B.n309 VSUBS 0.005941f
C355 B.n310 VSUBS 0.005941f
C356 B.n311 VSUBS 0.005941f
C357 B.n312 VSUBS 0.005941f
C358 B.n313 VSUBS 0.005941f
C359 B.n314 VSUBS 0.005941f
C360 B.n315 VSUBS 0.005941f
C361 B.n316 VSUBS 0.005941f
C362 B.n317 VSUBS 0.005941f
C363 B.n318 VSUBS 0.005941f
C364 B.n319 VSUBS 0.005941f
C365 B.n320 VSUBS 0.005941f
C366 B.n321 VSUBS 0.005941f
C367 B.n322 VSUBS 0.005941f
C368 B.n323 VSUBS 0.005941f
C369 B.n324 VSUBS 0.005941f
C370 B.n325 VSUBS 0.005941f
C371 B.n326 VSUBS 0.005941f
C372 B.n327 VSUBS 0.005941f
C373 B.n328 VSUBS 0.005941f
C374 B.n329 VSUBS 0.005941f
C375 B.n330 VSUBS 0.014263f
C376 B.n331 VSUBS 0.014916f
C377 B.n332 VSUBS 0.014263f
C378 B.n333 VSUBS 0.005941f
C379 B.n334 VSUBS 0.005941f
C380 B.n335 VSUBS 0.005941f
C381 B.n336 VSUBS 0.005941f
C382 B.n337 VSUBS 0.005941f
C383 B.n338 VSUBS 0.005941f
C384 B.n339 VSUBS 0.005941f
C385 B.n340 VSUBS 0.005941f
C386 B.n341 VSUBS 0.005941f
C387 B.n342 VSUBS 0.005941f
C388 B.n343 VSUBS 0.005941f
C389 B.n344 VSUBS 0.005941f
C390 B.n345 VSUBS 0.005941f
C391 B.n346 VSUBS 0.005941f
C392 B.n347 VSUBS 0.005941f
C393 B.n348 VSUBS 0.005941f
C394 B.n349 VSUBS 0.005941f
C395 B.n350 VSUBS 0.005941f
C396 B.n351 VSUBS 0.005941f
C397 B.n352 VSUBS 0.005941f
C398 B.n353 VSUBS 0.005941f
C399 B.n354 VSUBS 0.005941f
C400 B.n355 VSUBS 0.005941f
C401 B.n356 VSUBS 0.005941f
C402 B.n357 VSUBS 0.005941f
C403 B.n358 VSUBS 0.005941f
C404 B.n359 VSUBS 0.005941f
C405 B.n360 VSUBS 0.005941f
C406 B.n361 VSUBS 0.005941f
C407 B.n362 VSUBS 0.005941f
C408 B.n363 VSUBS 0.005941f
C409 B.n364 VSUBS 0.005941f
C410 B.n365 VSUBS 0.005941f
C411 B.n366 VSUBS 0.005941f
C412 B.n367 VSUBS 0.005941f
C413 B.n368 VSUBS 0.005941f
C414 B.n369 VSUBS 0.005941f
C415 B.n370 VSUBS 0.005941f
C416 B.n371 VSUBS 0.005941f
C417 B.n372 VSUBS 0.005941f
C418 B.n373 VSUBS 0.005941f
C419 B.n374 VSUBS 0.005941f
C420 B.n375 VSUBS 0.005941f
C421 B.n376 VSUBS 0.005941f
C422 B.n377 VSUBS 0.005941f
C423 B.n378 VSUBS 0.005941f
C424 B.n379 VSUBS 0.005941f
C425 B.n380 VSUBS 0.005941f
C426 B.n381 VSUBS 0.005941f
C427 B.n382 VSUBS 0.005941f
C428 B.n383 VSUBS 0.005941f
C429 B.n384 VSUBS 0.005941f
C430 B.n385 VSUBS 0.005941f
C431 B.n386 VSUBS 0.005941f
C432 B.n387 VSUBS 0.005941f
C433 B.n388 VSUBS 0.005941f
C434 B.n389 VSUBS 0.005941f
C435 B.n390 VSUBS 0.005941f
C436 B.n391 VSUBS 0.005941f
C437 B.n392 VSUBS 0.005941f
C438 B.n393 VSUBS 0.005941f
C439 B.n394 VSUBS 0.005941f
C440 B.n395 VSUBS 0.005941f
C441 B.n396 VSUBS 0.005941f
C442 B.n397 VSUBS 0.005941f
C443 B.n398 VSUBS 0.005941f
C444 B.n399 VSUBS 0.005941f
C445 B.n400 VSUBS 0.005941f
C446 B.n401 VSUBS 0.005941f
C447 B.n402 VSUBS 0.005941f
C448 B.n403 VSUBS 0.005941f
C449 B.n404 VSUBS 0.005941f
C450 B.n405 VSUBS 0.005941f
C451 B.n406 VSUBS 0.005941f
C452 B.n407 VSUBS 0.005941f
C453 B.n408 VSUBS 0.005941f
C454 B.n409 VSUBS 0.005941f
C455 B.n410 VSUBS 0.005941f
C456 B.n411 VSUBS 0.005941f
C457 B.n412 VSUBS 0.005941f
C458 B.n413 VSUBS 0.005941f
C459 B.n414 VSUBS 0.005941f
C460 B.n415 VSUBS 0.005941f
C461 B.n416 VSUBS 0.005941f
C462 B.n417 VSUBS 0.005941f
C463 B.n418 VSUBS 0.005941f
C464 B.n419 VSUBS 0.005941f
C465 B.n420 VSUBS 0.005941f
C466 B.n421 VSUBS 0.005941f
C467 B.n422 VSUBS 0.005941f
C468 B.n423 VSUBS 0.005941f
C469 B.n424 VSUBS 0.005941f
C470 B.n425 VSUBS 0.005941f
C471 B.n426 VSUBS 0.005941f
C472 B.n427 VSUBS 0.005941f
C473 B.n428 VSUBS 0.005941f
C474 B.n429 VSUBS 0.014263f
C475 B.n430 VSUBS 0.014263f
C476 B.n431 VSUBS 0.014916f
C477 B.n432 VSUBS 0.005941f
C478 B.n433 VSUBS 0.005941f
C479 B.n434 VSUBS 0.005941f
C480 B.n435 VSUBS 0.005941f
C481 B.n436 VSUBS 0.005941f
C482 B.n437 VSUBS 0.005941f
C483 B.n438 VSUBS 0.005941f
C484 B.n439 VSUBS 0.005941f
C485 B.n440 VSUBS 0.005941f
C486 B.n441 VSUBS 0.005941f
C487 B.n442 VSUBS 0.005941f
C488 B.n443 VSUBS 0.005941f
C489 B.n444 VSUBS 0.005941f
C490 B.n445 VSUBS 0.005941f
C491 B.n446 VSUBS 0.005941f
C492 B.n447 VSUBS 0.005941f
C493 B.n448 VSUBS 0.005941f
C494 B.n449 VSUBS 0.005941f
C495 B.n450 VSUBS 0.005941f
C496 B.n451 VSUBS 0.005941f
C497 B.n452 VSUBS 0.005941f
C498 B.n453 VSUBS 0.005941f
C499 B.n454 VSUBS 0.005941f
C500 B.n455 VSUBS 0.005941f
C501 B.n456 VSUBS 0.005941f
C502 B.n457 VSUBS 0.005941f
C503 B.n458 VSUBS 0.005941f
C504 B.n459 VSUBS 0.005941f
C505 B.n460 VSUBS 0.005941f
C506 B.n461 VSUBS 0.005941f
C507 B.n462 VSUBS 0.005941f
C508 B.n463 VSUBS 0.005941f
C509 B.n464 VSUBS 0.005941f
C510 B.n465 VSUBS 0.005941f
C511 B.n466 VSUBS 0.005941f
C512 B.n467 VSUBS 0.005941f
C513 B.n468 VSUBS 0.005941f
C514 B.n469 VSUBS 0.005941f
C515 B.n470 VSUBS 0.005941f
C516 B.n471 VSUBS 0.005941f
C517 B.n472 VSUBS 0.005941f
C518 B.n473 VSUBS 0.005941f
C519 B.n474 VSUBS 0.005941f
C520 B.n475 VSUBS 0.005941f
C521 B.n476 VSUBS 0.005941f
C522 B.n477 VSUBS 0.005941f
C523 B.n478 VSUBS 0.005941f
C524 B.n479 VSUBS 0.005941f
C525 B.n480 VSUBS 0.005941f
C526 B.n481 VSUBS 0.005941f
C527 B.n482 VSUBS 0.005941f
C528 B.n483 VSUBS 0.005941f
C529 B.n484 VSUBS 0.005941f
C530 B.n485 VSUBS 0.004106f
C531 B.n486 VSUBS 0.013764f
C532 B.n487 VSUBS 0.004805f
C533 B.n488 VSUBS 0.005941f
C534 B.n489 VSUBS 0.005941f
C535 B.n490 VSUBS 0.005941f
C536 B.n491 VSUBS 0.005941f
C537 B.n492 VSUBS 0.005941f
C538 B.n493 VSUBS 0.005941f
C539 B.n494 VSUBS 0.005941f
C540 B.n495 VSUBS 0.005941f
C541 B.n496 VSUBS 0.005941f
C542 B.n497 VSUBS 0.005941f
C543 B.n498 VSUBS 0.005941f
C544 B.n499 VSUBS 0.004805f
C545 B.n500 VSUBS 0.005941f
C546 B.n501 VSUBS 0.005941f
C547 B.n502 VSUBS 0.005941f
C548 B.n503 VSUBS 0.005941f
C549 B.n504 VSUBS 0.005941f
C550 B.n505 VSUBS 0.005941f
C551 B.n506 VSUBS 0.005941f
C552 B.n507 VSUBS 0.005941f
C553 B.n508 VSUBS 0.005941f
C554 B.n509 VSUBS 0.005941f
C555 B.n510 VSUBS 0.005941f
C556 B.n511 VSUBS 0.005941f
C557 B.n512 VSUBS 0.005941f
C558 B.n513 VSUBS 0.005941f
C559 B.n514 VSUBS 0.005941f
C560 B.n515 VSUBS 0.005941f
C561 B.n516 VSUBS 0.005941f
C562 B.n517 VSUBS 0.005941f
C563 B.n518 VSUBS 0.005941f
C564 B.n519 VSUBS 0.005941f
C565 B.n520 VSUBS 0.005941f
C566 B.n521 VSUBS 0.005941f
C567 B.n522 VSUBS 0.005941f
C568 B.n523 VSUBS 0.005941f
C569 B.n524 VSUBS 0.005941f
C570 B.n525 VSUBS 0.005941f
C571 B.n526 VSUBS 0.005941f
C572 B.n527 VSUBS 0.005941f
C573 B.n528 VSUBS 0.005941f
C574 B.n529 VSUBS 0.005941f
C575 B.n530 VSUBS 0.005941f
C576 B.n531 VSUBS 0.005941f
C577 B.n532 VSUBS 0.005941f
C578 B.n533 VSUBS 0.005941f
C579 B.n534 VSUBS 0.005941f
C580 B.n535 VSUBS 0.005941f
C581 B.n536 VSUBS 0.005941f
C582 B.n537 VSUBS 0.005941f
C583 B.n538 VSUBS 0.005941f
C584 B.n539 VSUBS 0.005941f
C585 B.n540 VSUBS 0.005941f
C586 B.n541 VSUBS 0.005941f
C587 B.n542 VSUBS 0.005941f
C588 B.n543 VSUBS 0.005941f
C589 B.n544 VSUBS 0.005941f
C590 B.n545 VSUBS 0.005941f
C591 B.n546 VSUBS 0.005941f
C592 B.n547 VSUBS 0.005941f
C593 B.n548 VSUBS 0.005941f
C594 B.n549 VSUBS 0.005941f
C595 B.n550 VSUBS 0.005941f
C596 B.n551 VSUBS 0.005941f
C597 B.n552 VSUBS 0.005941f
C598 B.n553 VSUBS 0.005941f
C599 B.n554 VSUBS 0.005941f
C600 B.n555 VSUBS 0.014916f
C601 B.n556 VSUBS 0.014263f
C602 B.n557 VSUBS 0.014263f
C603 B.n558 VSUBS 0.005941f
C604 B.n559 VSUBS 0.005941f
C605 B.n560 VSUBS 0.005941f
C606 B.n561 VSUBS 0.005941f
C607 B.n562 VSUBS 0.005941f
C608 B.n563 VSUBS 0.005941f
C609 B.n564 VSUBS 0.005941f
C610 B.n565 VSUBS 0.005941f
C611 B.n566 VSUBS 0.005941f
C612 B.n567 VSUBS 0.005941f
C613 B.n568 VSUBS 0.005941f
C614 B.n569 VSUBS 0.005941f
C615 B.n570 VSUBS 0.005941f
C616 B.n571 VSUBS 0.005941f
C617 B.n572 VSUBS 0.005941f
C618 B.n573 VSUBS 0.005941f
C619 B.n574 VSUBS 0.005941f
C620 B.n575 VSUBS 0.005941f
C621 B.n576 VSUBS 0.005941f
C622 B.n577 VSUBS 0.005941f
C623 B.n578 VSUBS 0.005941f
C624 B.n579 VSUBS 0.005941f
C625 B.n580 VSUBS 0.005941f
C626 B.n581 VSUBS 0.005941f
C627 B.n582 VSUBS 0.005941f
C628 B.n583 VSUBS 0.005941f
C629 B.n584 VSUBS 0.005941f
C630 B.n585 VSUBS 0.005941f
C631 B.n586 VSUBS 0.005941f
C632 B.n587 VSUBS 0.005941f
C633 B.n588 VSUBS 0.005941f
C634 B.n589 VSUBS 0.005941f
C635 B.n590 VSUBS 0.005941f
C636 B.n591 VSUBS 0.005941f
C637 B.n592 VSUBS 0.005941f
C638 B.n593 VSUBS 0.005941f
C639 B.n594 VSUBS 0.005941f
C640 B.n595 VSUBS 0.005941f
C641 B.n596 VSUBS 0.005941f
C642 B.n597 VSUBS 0.005941f
C643 B.n598 VSUBS 0.005941f
C644 B.n599 VSUBS 0.005941f
C645 B.n600 VSUBS 0.005941f
C646 B.n601 VSUBS 0.005941f
C647 B.n602 VSUBS 0.005941f
C648 B.n603 VSUBS 0.007752f
C649 B.n604 VSUBS 0.008258f
C650 B.n605 VSUBS 0.016422f
C651 VDD1.t0 VSUBS 1.7152f
C652 VDD1.t1 VSUBS 2.31844f
C653 VTAIL.t2 VSUBS 2.37702f
C654 VTAIL.n0 VSUBS 2.969f
C655 VTAIL.t1 VSUBS 2.37703f
C656 VTAIL.n1 VSUBS 3.05334f
C657 VTAIL.t3 VSUBS 2.37702f
C658 VTAIL.n2 VSUBS 2.69261f
C659 VTAIL.t0 VSUBS 2.37702f
C660 VTAIL.n3 VSUBS 2.54944f
C661 VP.t1 VSUBS 5.36102f
C662 VP.t0 VSUBS 4.36941f
C663 VP.n0 VSUBS 5.1182f
.ends

