* NGSPICE file created from diff_pair_sample_1435.ext - technology: sky130A

.subckt diff_pair_sample_1435 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=3.7635 ps=20.08 w=9.65 l=0.69
X1 VDD1.t8 VP.t1 VTAIL.t11 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X2 VDD2.t9 VN.t0 VTAIL.t6 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=3.7635 ps=20.08 w=9.65 l=0.69
X3 VDD2.t8 VN.t1 VTAIL.t2 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X4 VDD2.t7 VN.t2 VTAIL.t4 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=1.59225 ps=9.98 w=9.65 l=0.69
X5 VDD1.t7 VP.t2 VTAIL.t18 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=1.59225 ps=9.98 w=9.65 l=0.69
X6 B.t11 B.t9 B.t10 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=0 ps=0 w=9.65 l=0.69
X7 VDD2.t6 VN.t3 VTAIL.t7 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=3.7635 ps=20.08 w=9.65 l=0.69
X8 VTAIL.t0 VN.t4 VDD2.t5 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X9 VTAIL.t8 VN.t5 VDD2.t4 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X10 VTAIL.t9 VN.t6 VDD2.t3 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X11 B.t8 B.t6 B.t7 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=0 ps=0 w=9.65 l=0.69
X12 VDD2.t2 VN.t7 VTAIL.t1 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X13 VDD1.t6 VP.t3 VTAIL.t17 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=1.59225 ps=9.98 w=9.65 l=0.69
X14 VTAIL.t16 VP.t4 VDD1.t5 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X15 VTAIL.t13 VP.t5 VDD1.t4 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X16 VTAIL.t5 VN.t8 VDD2.t1 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X17 VTAIL.t19 VP.t6 VDD1.t3 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X18 VDD1.t2 VP.t7 VTAIL.t14 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X19 VDD2.t0 VN.t9 VTAIL.t3 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=1.59225 ps=9.98 w=9.65 l=0.69
X20 B.t5 B.t3 B.t4 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=0 ps=0 w=9.65 l=0.69
X21 VTAIL.t15 VP.t8 VDD1.t1 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=1.59225 ps=9.98 w=9.65 l=0.69
X22 VDD1.t0 VP.t9 VTAIL.t10 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=1.59225 pd=9.98 as=3.7635 ps=20.08 w=9.65 l=0.69
X23 B.t2 B.t0 B.t1 w_n2194_n2898# sky130_fd_pr__pfet_01v8 ad=3.7635 pd=20.08 as=0 ps=0 w=9.65 l=0.69
R0 VP.n7 VP.t3 416.51
R1 VP.n18 VP.t2 394.332
R2 VP.n22 VP.t5 394.332
R3 VP.n24 VP.t1 394.332
R4 VP.n28 VP.t4 394.332
R5 VP.n30 VP.t0 394.332
R6 VP.n16 VP.t9 394.332
R7 VP.n14 VP.t8 394.332
R8 VP.n6 VP.t7 394.332
R9 VP.n8 VP.t6 394.332
R10 VP.n31 VP.n30 161.3
R11 VP.n10 VP.n9 161.3
R12 VP.n11 VP.n6 161.3
R13 VP.n13 VP.n12 161.3
R14 VP.n14 VP.n5 161.3
R15 VP.n15 VP.n4 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n29 VP.n0 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.n1 161.3
R20 VP.n25 VP.n24 161.3
R21 VP.n23 VP.n2 161.3
R22 VP.n22 VP.n21 161.3
R23 VP.n20 VP.n3 161.3
R24 VP.n19 VP.n18 161.3
R25 VP.n10 VP.n7 44.862
R26 VP.n19 VP.n17 40.9323
R27 VP.n18 VP.n3 28.4823
R28 VP.n30 VP.n29 28.4823
R29 VP.n16 VP.n15 28.4823
R30 VP.n23 VP.n22 25.5611
R31 VP.n28 VP.n1 25.5611
R32 VP.n14 VP.n13 25.5611
R33 VP.n9 VP.n8 25.5611
R34 VP.n24 VP.n23 22.6399
R35 VP.n24 VP.n1 22.6399
R36 VP.n13 VP.n6 22.6399
R37 VP.n9 VP.n6 22.6399
R38 VP.n22 VP.n3 19.7187
R39 VP.n29 VP.n28 19.7187
R40 VP.n15 VP.n14 19.7187
R41 VP.n8 VP.n7 19.7081
R42 VP.n11 VP.n10 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n5 0.189894
R45 VP.n5 VP.n4 0.189894
R46 VP.n17 VP.n4 0.189894
R47 VP.n20 VP.n19 0.189894
R48 VP.n21 VP.n20 0.189894
R49 VP.n21 VP.n2 0.189894
R50 VP.n25 VP.n2 0.189894
R51 VP.n26 VP.n25 0.189894
R52 VP.n27 VP.n26 0.189894
R53 VP.n27 VP.n0 0.189894
R54 VP.n31 VP.n0 0.189894
R55 VP VP.n31 0.0516364
R56 VTAIL.n11 VTAIL.t7 65.4796
R57 VTAIL.n17 VTAIL.t6 65.4795
R58 VTAIL.n2 VTAIL.t12 65.4795
R59 VTAIL.n16 VTAIL.t10 65.4795
R60 VTAIL.n15 VTAIL.n14 62.1113
R61 VTAIL.n13 VTAIL.n12 62.1113
R62 VTAIL.n10 VTAIL.n9 62.1113
R63 VTAIL.n8 VTAIL.n7 62.1113
R64 VTAIL.n19 VTAIL.n18 62.111
R65 VTAIL.n1 VTAIL.n0 62.111
R66 VTAIL.n4 VTAIL.n3 62.111
R67 VTAIL.n6 VTAIL.n5 62.111
R68 VTAIL.n8 VTAIL.n6 22.4445
R69 VTAIL.n17 VTAIL.n16 21.5652
R70 VTAIL.n18 VTAIL.t2 3.36889
R71 VTAIL.n18 VTAIL.t0 3.36889
R72 VTAIL.n0 VTAIL.t4 3.36889
R73 VTAIL.n0 VTAIL.t8 3.36889
R74 VTAIL.n3 VTAIL.t11 3.36889
R75 VTAIL.n3 VTAIL.t16 3.36889
R76 VTAIL.n5 VTAIL.t18 3.36889
R77 VTAIL.n5 VTAIL.t13 3.36889
R78 VTAIL.n14 VTAIL.t14 3.36889
R79 VTAIL.n14 VTAIL.t15 3.36889
R80 VTAIL.n12 VTAIL.t17 3.36889
R81 VTAIL.n12 VTAIL.t19 3.36889
R82 VTAIL.n9 VTAIL.t1 3.36889
R83 VTAIL.n9 VTAIL.t9 3.36889
R84 VTAIL.n7 VTAIL.t3 3.36889
R85 VTAIL.n7 VTAIL.t5 3.36889
R86 VTAIL.n13 VTAIL.n11 0.909983
R87 VTAIL.n2 VTAIL.n1 0.909983
R88 VTAIL.n10 VTAIL.n8 0.87981
R89 VTAIL.n11 VTAIL.n10 0.87981
R90 VTAIL.n15 VTAIL.n13 0.87981
R91 VTAIL.n16 VTAIL.n15 0.87981
R92 VTAIL.n6 VTAIL.n4 0.87981
R93 VTAIL.n4 VTAIL.n2 0.87981
R94 VTAIL.n19 VTAIL.n17 0.87981
R95 VTAIL VTAIL.n1 0.718172
R96 VTAIL VTAIL.n19 0.162138
R97 VDD1.n1 VDD1.t6 83.0377
R98 VDD1.n3 VDD1.t7 83.0376
R99 VDD1.n5 VDD1.n4 79.394
R100 VDD1.n1 VDD1.n0 78.7901
R101 VDD1.n7 VDD1.n6 78.7899
R102 VDD1.n3 VDD1.n2 78.7898
R103 VDD1.n7 VDD1.n5 37.2337
R104 VDD1.n6 VDD1.t1 3.36889
R105 VDD1.n6 VDD1.t0 3.36889
R106 VDD1.n0 VDD1.t3 3.36889
R107 VDD1.n0 VDD1.t2 3.36889
R108 VDD1.n4 VDD1.t5 3.36889
R109 VDD1.n4 VDD1.t9 3.36889
R110 VDD1.n2 VDD1.t4 3.36889
R111 VDD1.n2 VDD1.t8 3.36889
R112 VDD1 VDD1.n7 0.601793
R113 VDD1 VDD1.n1 0.278517
R114 VDD1.n5 VDD1.n3 0.164982
R115 VN.n3 VN.t2 416.51
R116 VN.n17 VN.t3 416.51
R117 VN.n4 VN.t5 394.332
R118 VN.n6 VN.t1 394.332
R119 VN.n10 VN.t4 394.332
R120 VN.n12 VN.t0 394.332
R121 VN.n18 VN.t6 394.332
R122 VN.n20 VN.t7 394.332
R123 VN.n24 VN.t8 394.332
R124 VN.n26 VN.t9 394.332
R125 VN.n13 VN.n12 161.3
R126 VN.n27 VN.n26 161.3
R127 VN.n25 VN.n14 161.3
R128 VN.n24 VN.n23 161.3
R129 VN.n22 VN.n15 161.3
R130 VN.n21 VN.n20 161.3
R131 VN.n19 VN.n16 161.3
R132 VN.n11 VN.n0 161.3
R133 VN.n10 VN.n9 161.3
R134 VN.n8 VN.n1 161.3
R135 VN.n7 VN.n6 161.3
R136 VN.n5 VN.n2 161.3
R137 VN.n17 VN.n16 44.862
R138 VN.n3 VN.n2 44.862
R139 VN VN.n27 41.313
R140 VN.n12 VN.n11 28.4823
R141 VN.n26 VN.n25 28.4823
R142 VN.n5 VN.n4 25.5611
R143 VN.n10 VN.n1 25.5611
R144 VN.n19 VN.n18 25.5611
R145 VN.n24 VN.n15 25.5611
R146 VN.n6 VN.n5 22.6399
R147 VN.n6 VN.n1 22.6399
R148 VN.n20 VN.n19 22.6399
R149 VN.n20 VN.n15 22.6399
R150 VN.n11 VN.n10 19.7187
R151 VN.n25 VN.n24 19.7187
R152 VN.n4 VN.n3 19.7081
R153 VN.n18 VN.n17 19.7081
R154 VN.n27 VN.n14 0.189894
R155 VN.n23 VN.n14 0.189894
R156 VN.n23 VN.n22 0.189894
R157 VN.n22 VN.n21 0.189894
R158 VN.n21 VN.n16 0.189894
R159 VN.n7 VN.n2 0.189894
R160 VN.n8 VN.n7 0.189894
R161 VN.n9 VN.n8 0.189894
R162 VN.n9 VN.n0 0.189894
R163 VN.n13 VN.n0 0.189894
R164 VN VN.n13 0.0516364
R165 VDD2.n1 VDD2.t7 83.0376
R166 VDD2.n4 VDD2.t0 82.1584
R167 VDD2.n3 VDD2.n2 79.394
R168 VDD2 VDD2.n7 79.3912
R169 VDD2.n6 VDD2.n5 78.7901
R170 VDD2.n1 VDD2.n0 78.7898
R171 VDD2.n4 VDD2.n3 36.211
R172 VDD2.n7 VDD2.t3 3.36889
R173 VDD2.n7 VDD2.t6 3.36889
R174 VDD2.n5 VDD2.t1 3.36889
R175 VDD2.n5 VDD2.t2 3.36889
R176 VDD2.n2 VDD2.t5 3.36889
R177 VDD2.n2 VDD2.t9 3.36889
R178 VDD2.n0 VDD2.t4 3.36889
R179 VDD2.n0 VDD2.t8 3.36889
R180 VDD2.n6 VDD2.n4 0.87981
R181 VDD2 VDD2.n6 0.278517
R182 VDD2.n3 VDD2.n1 0.164982
R183 B.n380 B.n59 585
R184 B.n382 B.n381 585
R185 B.n383 B.n58 585
R186 B.n385 B.n384 585
R187 B.n386 B.n57 585
R188 B.n388 B.n387 585
R189 B.n389 B.n56 585
R190 B.n391 B.n390 585
R191 B.n392 B.n55 585
R192 B.n394 B.n393 585
R193 B.n395 B.n54 585
R194 B.n397 B.n396 585
R195 B.n398 B.n53 585
R196 B.n400 B.n399 585
R197 B.n401 B.n52 585
R198 B.n403 B.n402 585
R199 B.n404 B.n51 585
R200 B.n406 B.n405 585
R201 B.n407 B.n50 585
R202 B.n409 B.n408 585
R203 B.n410 B.n49 585
R204 B.n412 B.n411 585
R205 B.n413 B.n48 585
R206 B.n415 B.n414 585
R207 B.n416 B.n47 585
R208 B.n418 B.n417 585
R209 B.n419 B.n46 585
R210 B.n421 B.n420 585
R211 B.n422 B.n45 585
R212 B.n424 B.n423 585
R213 B.n425 B.n44 585
R214 B.n427 B.n426 585
R215 B.n428 B.n43 585
R216 B.n430 B.n429 585
R217 B.n431 B.n40 585
R218 B.n434 B.n433 585
R219 B.n435 B.n39 585
R220 B.n437 B.n436 585
R221 B.n438 B.n38 585
R222 B.n440 B.n439 585
R223 B.n441 B.n37 585
R224 B.n443 B.n442 585
R225 B.n444 B.n33 585
R226 B.n446 B.n445 585
R227 B.n447 B.n32 585
R228 B.n449 B.n448 585
R229 B.n450 B.n31 585
R230 B.n452 B.n451 585
R231 B.n453 B.n30 585
R232 B.n455 B.n454 585
R233 B.n456 B.n29 585
R234 B.n458 B.n457 585
R235 B.n459 B.n28 585
R236 B.n461 B.n460 585
R237 B.n462 B.n27 585
R238 B.n464 B.n463 585
R239 B.n465 B.n26 585
R240 B.n467 B.n466 585
R241 B.n468 B.n25 585
R242 B.n470 B.n469 585
R243 B.n471 B.n24 585
R244 B.n473 B.n472 585
R245 B.n474 B.n23 585
R246 B.n476 B.n475 585
R247 B.n477 B.n22 585
R248 B.n479 B.n478 585
R249 B.n480 B.n21 585
R250 B.n482 B.n481 585
R251 B.n483 B.n20 585
R252 B.n485 B.n484 585
R253 B.n486 B.n19 585
R254 B.n488 B.n487 585
R255 B.n489 B.n18 585
R256 B.n491 B.n490 585
R257 B.n492 B.n17 585
R258 B.n494 B.n493 585
R259 B.n495 B.n16 585
R260 B.n497 B.n496 585
R261 B.n498 B.n15 585
R262 B.n379 B.n378 585
R263 B.n377 B.n60 585
R264 B.n376 B.n375 585
R265 B.n374 B.n61 585
R266 B.n373 B.n372 585
R267 B.n371 B.n62 585
R268 B.n370 B.n369 585
R269 B.n368 B.n63 585
R270 B.n367 B.n366 585
R271 B.n365 B.n64 585
R272 B.n364 B.n363 585
R273 B.n362 B.n65 585
R274 B.n361 B.n360 585
R275 B.n359 B.n66 585
R276 B.n358 B.n357 585
R277 B.n356 B.n67 585
R278 B.n355 B.n354 585
R279 B.n353 B.n68 585
R280 B.n352 B.n351 585
R281 B.n350 B.n69 585
R282 B.n349 B.n348 585
R283 B.n347 B.n70 585
R284 B.n346 B.n345 585
R285 B.n344 B.n71 585
R286 B.n343 B.n342 585
R287 B.n341 B.n72 585
R288 B.n340 B.n339 585
R289 B.n338 B.n73 585
R290 B.n337 B.n336 585
R291 B.n335 B.n74 585
R292 B.n334 B.n333 585
R293 B.n332 B.n75 585
R294 B.n331 B.n330 585
R295 B.n329 B.n76 585
R296 B.n328 B.n327 585
R297 B.n326 B.n77 585
R298 B.n325 B.n324 585
R299 B.n323 B.n78 585
R300 B.n322 B.n321 585
R301 B.n320 B.n79 585
R302 B.n319 B.n318 585
R303 B.n317 B.n80 585
R304 B.n316 B.n315 585
R305 B.n314 B.n81 585
R306 B.n313 B.n312 585
R307 B.n311 B.n82 585
R308 B.n310 B.n309 585
R309 B.n308 B.n83 585
R310 B.n307 B.n306 585
R311 B.n305 B.n84 585
R312 B.n304 B.n303 585
R313 B.n302 B.n85 585
R314 B.n301 B.n300 585
R315 B.n178 B.n127 585
R316 B.n180 B.n179 585
R317 B.n181 B.n126 585
R318 B.n183 B.n182 585
R319 B.n184 B.n125 585
R320 B.n186 B.n185 585
R321 B.n187 B.n124 585
R322 B.n189 B.n188 585
R323 B.n190 B.n123 585
R324 B.n192 B.n191 585
R325 B.n193 B.n122 585
R326 B.n195 B.n194 585
R327 B.n196 B.n121 585
R328 B.n198 B.n197 585
R329 B.n199 B.n120 585
R330 B.n201 B.n200 585
R331 B.n202 B.n119 585
R332 B.n204 B.n203 585
R333 B.n205 B.n118 585
R334 B.n207 B.n206 585
R335 B.n208 B.n117 585
R336 B.n210 B.n209 585
R337 B.n211 B.n116 585
R338 B.n213 B.n212 585
R339 B.n214 B.n115 585
R340 B.n216 B.n215 585
R341 B.n217 B.n114 585
R342 B.n219 B.n218 585
R343 B.n220 B.n113 585
R344 B.n222 B.n221 585
R345 B.n223 B.n112 585
R346 B.n225 B.n224 585
R347 B.n226 B.n111 585
R348 B.n228 B.n227 585
R349 B.n229 B.n108 585
R350 B.n232 B.n231 585
R351 B.n233 B.n107 585
R352 B.n235 B.n234 585
R353 B.n236 B.n106 585
R354 B.n238 B.n237 585
R355 B.n239 B.n105 585
R356 B.n241 B.n240 585
R357 B.n242 B.n104 585
R358 B.n247 B.n246 585
R359 B.n248 B.n103 585
R360 B.n250 B.n249 585
R361 B.n251 B.n102 585
R362 B.n253 B.n252 585
R363 B.n254 B.n101 585
R364 B.n256 B.n255 585
R365 B.n257 B.n100 585
R366 B.n259 B.n258 585
R367 B.n260 B.n99 585
R368 B.n262 B.n261 585
R369 B.n263 B.n98 585
R370 B.n265 B.n264 585
R371 B.n266 B.n97 585
R372 B.n268 B.n267 585
R373 B.n269 B.n96 585
R374 B.n271 B.n270 585
R375 B.n272 B.n95 585
R376 B.n274 B.n273 585
R377 B.n275 B.n94 585
R378 B.n277 B.n276 585
R379 B.n278 B.n93 585
R380 B.n280 B.n279 585
R381 B.n281 B.n92 585
R382 B.n283 B.n282 585
R383 B.n284 B.n91 585
R384 B.n286 B.n285 585
R385 B.n287 B.n90 585
R386 B.n289 B.n288 585
R387 B.n290 B.n89 585
R388 B.n292 B.n291 585
R389 B.n293 B.n88 585
R390 B.n295 B.n294 585
R391 B.n296 B.n87 585
R392 B.n298 B.n297 585
R393 B.n299 B.n86 585
R394 B.n177 B.n176 585
R395 B.n175 B.n128 585
R396 B.n174 B.n173 585
R397 B.n172 B.n129 585
R398 B.n171 B.n170 585
R399 B.n169 B.n130 585
R400 B.n168 B.n167 585
R401 B.n166 B.n131 585
R402 B.n165 B.n164 585
R403 B.n163 B.n132 585
R404 B.n162 B.n161 585
R405 B.n160 B.n133 585
R406 B.n159 B.n158 585
R407 B.n157 B.n134 585
R408 B.n156 B.n155 585
R409 B.n154 B.n135 585
R410 B.n153 B.n152 585
R411 B.n151 B.n136 585
R412 B.n150 B.n149 585
R413 B.n148 B.n137 585
R414 B.n147 B.n146 585
R415 B.n145 B.n138 585
R416 B.n144 B.n143 585
R417 B.n142 B.n139 585
R418 B.n141 B.n140 585
R419 B.n2 B.n0 585
R420 B.n537 B.n1 585
R421 B.n536 B.n535 585
R422 B.n534 B.n3 585
R423 B.n533 B.n532 585
R424 B.n531 B.n4 585
R425 B.n530 B.n529 585
R426 B.n528 B.n5 585
R427 B.n527 B.n526 585
R428 B.n525 B.n6 585
R429 B.n524 B.n523 585
R430 B.n522 B.n7 585
R431 B.n521 B.n520 585
R432 B.n519 B.n8 585
R433 B.n518 B.n517 585
R434 B.n516 B.n9 585
R435 B.n515 B.n514 585
R436 B.n513 B.n10 585
R437 B.n512 B.n511 585
R438 B.n510 B.n11 585
R439 B.n509 B.n508 585
R440 B.n507 B.n12 585
R441 B.n506 B.n505 585
R442 B.n504 B.n13 585
R443 B.n503 B.n502 585
R444 B.n501 B.n14 585
R445 B.n500 B.n499 585
R446 B.n539 B.n538 585
R447 B.n243 B.t9 540.14
R448 B.n109 B.t6 540.14
R449 B.n34 B.t3 540.14
R450 B.n41 B.t0 540.14
R451 B.n178 B.n177 516.524
R452 B.n500 B.n15 516.524
R453 B.n301 B.n86 516.524
R454 B.n380 B.n379 516.524
R455 B.n177 B.n128 163.367
R456 B.n173 B.n128 163.367
R457 B.n173 B.n172 163.367
R458 B.n172 B.n171 163.367
R459 B.n171 B.n130 163.367
R460 B.n167 B.n130 163.367
R461 B.n167 B.n166 163.367
R462 B.n166 B.n165 163.367
R463 B.n165 B.n132 163.367
R464 B.n161 B.n132 163.367
R465 B.n161 B.n160 163.367
R466 B.n160 B.n159 163.367
R467 B.n159 B.n134 163.367
R468 B.n155 B.n134 163.367
R469 B.n155 B.n154 163.367
R470 B.n154 B.n153 163.367
R471 B.n153 B.n136 163.367
R472 B.n149 B.n136 163.367
R473 B.n149 B.n148 163.367
R474 B.n148 B.n147 163.367
R475 B.n147 B.n138 163.367
R476 B.n143 B.n138 163.367
R477 B.n143 B.n142 163.367
R478 B.n142 B.n141 163.367
R479 B.n141 B.n2 163.367
R480 B.n538 B.n2 163.367
R481 B.n538 B.n537 163.367
R482 B.n537 B.n536 163.367
R483 B.n536 B.n3 163.367
R484 B.n532 B.n3 163.367
R485 B.n532 B.n531 163.367
R486 B.n531 B.n530 163.367
R487 B.n530 B.n5 163.367
R488 B.n526 B.n5 163.367
R489 B.n526 B.n525 163.367
R490 B.n525 B.n524 163.367
R491 B.n524 B.n7 163.367
R492 B.n520 B.n7 163.367
R493 B.n520 B.n519 163.367
R494 B.n519 B.n518 163.367
R495 B.n518 B.n9 163.367
R496 B.n514 B.n9 163.367
R497 B.n514 B.n513 163.367
R498 B.n513 B.n512 163.367
R499 B.n512 B.n11 163.367
R500 B.n508 B.n11 163.367
R501 B.n508 B.n507 163.367
R502 B.n507 B.n506 163.367
R503 B.n506 B.n13 163.367
R504 B.n502 B.n13 163.367
R505 B.n502 B.n501 163.367
R506 B.n501 B.n500 163.367
R507 B.n179 B.n178 163.367
R508 B.n179 B.n126 163.367
R509 B.n183 B.n126 163.367
R510 B.n184 B.n183 163.367
R511 B.n185 B.n184 163.367
R512 B.n185 B.n124 163.367
R513 B.n189 B.n124 163.367
R514 B.n190 B.n189 163.367
R515 B.n191 B.n190 163.367
R516 B.n191 B.n122 163.367
R517 B.n195 B.n122 163.367
R518 B.n196 B.n195 163.367
R519 B.n197 B.n196 163.367
R520 B.n197 B.n120 163.367
R521 B.n201 B.n120 163.367
R522 B.n202 B.n201 163.367
R523 B.n203 B.n202 163.367
R524 B.n203 B.n118 163.367
R525 B.n207 B.n118 163.367
R526 B.n208 B.n207 163.367
R527 B.n209 B.n208 163.367
R528 B.n209 B.n116 163.367
R529 B.n213 B.n116 163.367
R530 B.n214 B.n213 163.367
R531 B.n215 B.n214 163.367
R532 B.n215 B.n114 163.367
R533 B.n219 B.n114 163.367
R534 B.n220 B.n219 163.367
R535 B.n221 B.n220 163.367
R536 B.n221 B.n112 163.367
R537 B.n225 B.n112 163.367
R538 B.n226 B.n225 163.367
R539 B.n227 B.n226 163.367
R540 B.n227 B.n108 163.367
R541 B.n232 B.n108 163.367
R542 B.n233 B.n232 163.367
R543 B.n234 B.n233 163.367
R544 B.n234 B.n106 163.367
R545 B.n238 B.n106 163.367
R546 B.n239 B.n238 163.367
R547 B.n240 B.n239 163.367
R548 B.n240 B.n104 163.367
R549 B.n247 B.n104 163.367
R550 B.n248 B.n247 163.367
R551 B.n249 B.n248 163.367
R552 B.n249 B.n102 163.367
R553 B.n253 B.n102 163.367
R554 B.n254 B.n253 163.367
R555 B.n255 B.n254 163.367
R556 B.n255 B.n100 163.367
R557 B.n259 B.n100 163.367
R558 B.n260 B.n259 163.367
R559 B.n261 B.n260 163.367
R560 B.n261 B.n98 163.367
R561 B.n265 B.n98 163.367
R562 B.n266 B.n265 163.367
R563 B.n267 B.n266 163.367
R564 B.n267 B.n96 163.367
R565 B.n271 B.n96 163.367
R566 B.n272 B.n271 163.367
R567 B.n273 B.n272 163.367
R568 B.n273 B.n94 163.367
R569 B.n277 B.n94 163.367
R570 B.n278 B.n277 163.367
R571 B.n279 B.n278 163.367
R572 B.n279 B.n92 163.367
R573 B.n283 B.n92 163.367
R574 B.n284 B.n283 163.367
R575 B.n285 B.n284 163.367
R576 B.n285 B.n90 163.367
R577 B.n289 B.n90 163.367
R578 B.n290 B.n289 163.367
R579 B.n291 B.n290 163.367
R580 B.n291 B.n88 163.367
R581 B.n295 B.n88 163.367
R582 B.n296 B.n295 163.367
R583 B.n297 B.n296 163.367
R584 B.n297 B.n86 163.367
R585 B.n302 B.n301 163.367
R586 B.n303 B.n302 163.367
R587 B.n303 B.n84 163.367
R588 B.n307 B.n84 163.367
R589 B.n308 B.n307 163.367
R590 B.n309 B.n308 163.367
R591 B.n309 B.n82 163.367
R592 B.n313 B.n82 163.367
R593 B.n314 B.n313 163.367
R594 B.n315 B.n314 163.367
R595 B.n315 B.n80 163.367
R596 B.n319 B.n80 163.367
R597 B.n320 B.n319 163.367
R598 B.n321 B.n320 163.367
R599 B.n321 B.n78 163.367
R600 B.n325 B.n78 163.367
R601 B.n326 B.n325 163.367
R602 B.n327 B.n326 163.367
R603 B.n327 B.n76 163.367
R604 B.n331 B.n76 163.367
R605 B.n332 B.n331 163.367
R606 B.n333 B.n332 163.367
R607 B.n333 B.n74 163.367
R608 B.n337 B.n74 163.367
R609 B.n338 B.n337 163.367
R610 B.n339 B.n338 163.367
R611 B.n339 B.n72 163.367
R612 B.n343 B.n72 163.367
R613 B.n344 B.n343 163.367
R614 B.n345 B.n344 163.367
R615 B.n345 B.n70 163.367
R616 B.n349 B.n70 163.367
R617 B.n350 B.n349 163.367
R618 B.n351 B.n350 163.367
R619 B.n351 B.n68 163.367
R620 B.n355 B.n68 163.367
R621 B.n356 B.n355 163.367
R622 B.n357 B.n356 163.367
R623 B.n357 B.n66 163.367
R624 B.n361 B.n66 163.367
R625 B.n362 B.n361 163.367
R626 B.n363 B.n362 163.367
R627 B.n363 B.n64 163.367
R628 B.n367 B.n64 163.367
R629 B.n368 B.n367 163.367
R630 B.n369 B.n368 163.367
R631 B.n369 B.n62 163.367
R632 B.n373 B.n62 163.367
R633 B.n374 B.n373 163.367
R634 B.n375 B.n374 163.367
R635 B.n375 B.n60 163.367
R636 B.n379 B.n60 163.367
R637 B.n496 B.n15 163.367
R638 B.n496 B.n495 163.367
R639 B.n495 B.n494 163.367
R640 B.n494 B.n17 163.367
R641 B.n490 B.n17 163.367
R642 B.n490 B.n489 163.367
R643 B.n489 B.n488 163.367
R644 B.n488 B.n19 163.367
R645 B.n484 B.n19 163.367
R646 B.n484 B.n483 163.367
R647 B.n483 B.n482 163.367
R648 B.n482 B.n21 163.367
R649 B.n478 B.n21 163.367
R650 B.n478 B.n477 163.367
R651 B.n477 B.n476 163.367
R652 B.n476 B.n23 163.367
R653 B.n472 B.n23 163.367
R654 B.n472 B.n471 163.367
R655 B.n471 B.n470 163.367
R656 B.n470 B.n25 163.367
R657 B.n466 B.n25 163.367
R658 B.n466 B.n465 163.367
R659 B.n465 B.n464 163.367
R660 B.n464 B.n27 163.367
R661 B.n460 B.n27 163.367
R662 B.n460 B.n459 163.367
R663 B.n459 B.n458 163.367
R664 B.n458 B.n29 163.367
R665 B.n454 B.n29 163.367
R666 B.n454 B.n453 163.367
R667 B.n453 B.n452 163.367
R668 B.n452 B.n31 163.367
R669 B.n448 B.n31 163.367
R670 B.n448 B.n447 163.367
R671 B.n447 B.n446 163.367
R672 B.n446 B.n33 163.367
R673 B.n442 B.n33 163.367
R674 B.n442 B.n441 163.367
R675 B.n441 B.n440 163.367
R676 B.n440 B.n38 163.367
R677 B.n436 B.n38 163.367
R678 B.n436 B.n435 163.367
R679 B.n435 B.n434 163.367
R680 B.n434 B.n40 163.367
R681 B.n429 B.n40 163.367
R682 B.n429 B.n428 163.367
R683 B.n428 B.n427 163.367
R684 B.n427 B.n44 163.367
R685 B.n423 B.n44 163.367
R686 B.n423 B.n422 163.367
R687 B.n422 B.n421 163.367
R688 B.n421 B.n46 163.367
R689 B.n417 B.n46 163.367
R690 B.n417 B.n416 163.367
R691 B.n416 B.n415 163.367
R692 B.n415 B.n48 163.367
R693 B.n411 B.n48 163.367
R694 B.n411 B.n410 163.367
R695 B.n410 B.n409 163.367
R696 B.n409 B.n50 163.367
R697 B.n405 B.n50 163.367
R698 B.n405 B.n404 163.367
R699 B.n404 B.n403 163.367
R700 B.n403 B.n52 163.367
R701 B.n399 B.n52 163.367
R702 B.n399 B.n398 163.367
R703 B.n398 B.n397 163.367
R704 B.n397 B.n54 163.367
R705 B.n393 B.n54 163.367
R706 B.n393 B.n392 163.367
R707 B.n392 B.n391 163.367
R708 B.n391 B.n56 163.367
R709 B.n387 B.n56 163.367
R710 B.n387 B.n386 163.367
R711 B.n386 B.n385 163.367
R712 B.n385 B.n58 163.367
R713 B.n381 B.n58 163.367
R714 B.n381 B.n380 163.367
R715 B.n243 B.t11 130.111
R716 B.n41 B.t1 130.111
R717 B.n109 B.t8 130.1
R718 B.n34 B.t4 130.1
R719 B.n244 B.t10 110.329
R720 B.n42 B.t2 110.329
R721 B.n110 B.t7 110.319
R722 B.n35 B.t5 110.319
R723 B.n245 B.n244 59.5399
R724 B.n230 B.n110 59.5399
R725 B.n36 B.n35 59.5399
R726 B.n432 B.n42 59.5399
R727 B.n499 B.n498 33.5615
R728 B.n378 B.n59 33.5615
R729 B.n300 B.n299 33.5615
R730 B.n176 B.n127 33.5615
R731 B.n244 B.n243 19.7823
R732 B.n110 B.n109 19.7823
R733 B.n35 B.n34 19.7823
R734 B.n42 B.n41 19.7823
R735 B B.n539 18.0485
R736 B.n498 B.n497 10.6151
R737 B.n497 B.n16 10.6151
R738 B.n493 B.n16 10.6151
R739 B.n493 B.n492 10.6151
R740 B.n492 B.n491 10.6151
R741 B.n491 B.n18 10.6151
R742 B.n487 B.n18 10.6151
R743 B.n487 B.n486 10.6151
R744 B.n486 B.n485 10.6151
R745 B.n485 B.n20 10.6151
R746 B.n481 B.n20 10.6151
R747 B.n481 B.n480 10.6151
R748 B.n480 B.n479 10.6151
R749 B.n479 B.n22 10.6151
R750 B.n475 B.n22 10.6151
R751 B.n475 B.n474 10.6151
R752 B.n474 B.n473 10.6151
R753 B.n473 B.n24 10.6151
R754 B.n469 B.n24 10.6151
R755 B.n469 B.n468 10.6151
R756 B.n468 B.n467 10.6151
R757 B.n467 B.n26 10.6151
R758 B.n463 B.n26 10.6151
R759 B.n463 B.n462 10.6151
R760 B.n462 B.n461 10.6151
R761 B.n461 B.n28 10.6151
R762 B.n457 B.n28 10.6151
R763 B.n457 B.n456 10.6151
R764 B.n456 B.n455 10.6151
R765 B.n455 B.n30 10.6151
R766 B.n451 B.n30 10.6151
R767 B.n451 B.n450 10.6151
R768 B.n450 B.n449 10.6151
R769 B.n449 B.n32 10.6151
R770 B.n445 B.n444 10.6151
R771 B.n444 B.n443 10.6151
R772 B.n443 B.n37 10.6151
R773 B.n439 B.n37 10.6151
R774 B.n439 B.n438 10.6151
R775 B.n438 B.n437 10.6151
R776 B.n437 B.n39 10.6151
R777 B.n433 B.n39 10.6151
R778 B.n431 B.n430 10.6151
R779 B.n430 B.n43 10.6151
R780 B.n426 B.n43 10.6151
R781 B.n426 B.n425 10.6151
R782 B.n425 B.n424 10.6151
R783 B.n424 B.n45 10.6151
R784 B.n420 B.n45 10.6151
R785 B.n420 B.n419 10.6151
R786 B.n419 B.n418 10.6151
R787 B.n418 B.n47 10.6151
R788 B.n414 B.n47 10.6151
R789 B.n414 B.n413 10.6151
R790 B.n413 B.n412 10.6151
R791 B.n412 B.n49 10.6151
R792 B.n408 B.n49 10.6151
R793 B.n408 B.n407 10.6151
R794 B.n407 B.n406 10.6151
R795 B.n406 B.n51 10.6151
R796 B.n402 B.n51 10.6151
R797 B.n402 B.n401 10.6151
R798 B.n401 B.n400 10.6151
R799 B.n400 B.n53 10.6151
R800 B.n396 B.n53 10.6151
R801 B.n396 B.n395 10.6151
R802 B.n395 B.n394 10.6151
R803 B.n394 B.n55 10.6151
R804 B.n390 B.n55 10.6151
R805 B.n390 B.n389 10.6151
R806 B.n389 B.n388 10.6151
R807 B.n388 B.n57 10.6151
R808 B.n384 B.n57 10.6151
R809 B.n384 B.n383 10.6151
R810 B.n383 B.n382 10.6151
R811 B.n382 B.n59 10.6151
R812 B.n300 B.n85 10.6151
R813 B.n304 B.n85 10.6151
R814 B.n305 B.n304 10.6151
R815 B.n306 B.n305 10.6151
R816 B.n306 B.n83 10.6151
R817 B.n310 B.n83 10.6151
R818 B.n311 B.n310 10.6151
R819 B.n312 B.n311 10.6151
R820 B.n312 B.n81 10.6151
R821 B.n316 B.n81 10.6151
R822 B.n317 B.n316 10.6151
R823 B.n318 B.n317 10.6151
R824 B.n318 B.n79 10.6151
R825 B.n322 B.n79 10.6151
R826 B.n323 B.n322 10.6151
R827 B.n324 B.n323 10.6151
R828 B.n324 B.n77 10.6151
R829 B.n328 B.n77 10.6151
R830 B.n329 B.n328 10.6151
R831 B.n330 B.n329 10.6151
R832 B.n330 B.n75 10.6151
R833 B.n334 B.n75 10.6151
R834 B.n335 B.n334 10.6151
R835 B.n336 B.n335 10.6151
R836 B.n336 B.n73 10.6151
R837 B.n340 B.n73 10.6151
R838 B.n341 B.n340 10.6151
R839 B.n342 B.n341 10.6151
R840 B.n342 B.n71 10.6151
R841 B.n346 B.n71 10.6151
R842 B.n347 B.n346 10.6151
R843 B.n348 B.n347 10.6151
R844 B.n348 B.n69 10.6151
R845 B.n352 B.n69 10.6151
R846 B.n353 B.n352 10.6151
R847 B.n354 B.n353 10.6151
R848 B.n354 B.n67 10.6151
R849 B.n358 B.n67 10.6151
R850 B.n359 B.n358 10.6151
R851 B.n360 B.n359 10.6151
R852 B.n360 B.n65 10.6151
R853 B.n364 B.n65 10.6151
R854 B.n365 B.n364 10.6151
R855 B.n366 B.n365 10.6151
R856 B.n366 B.n63 10.6151
R857 B.n370 B.n63 10.6151
R858 B.n371 B.n370 10.6151
R859 B.n372 B.n371 10.6151
R860 B.n372 B.n61 10.6151
R861 B.n376 B.n61 10.6151
R862 B.n377 B.n376 10.6151
R863 B.n378 B.n377 10.6151
R864 B.n180 B.n127 10.6151
R865 B.n181 B.n180 10.6151
R866 B.n182 B.n181 10.6151
R867 B.n182 B.n125 10.6151
R868 B.n186 B.n125 10.6151
R869 B.n187 B.n186 10.6151
R870 B.n188 B.n187 10.6151
R871 B.n188 B.n123 10.6151
R872 B.n192 B.n123 10.6151
R873 B.n193 B.n192 10.6151
R874 B.n194 B.n193 10.6151
R875 B.n194 B.n121 10.6151
R876 B.n198 B.n121 10.6151
R877 B.n199 B.n198 10.6151
R878 B.n200 B.n199 10.6151
R879 B.n200 B.n119 10.6151
R880 B.n204 B.n119 10.6151
R881 B.n205 B.n204 10.6151
R882 B.n206 B.n205 10.6151
R883 B.n206 B.n117 10.6151
R884 B.n210 B.n117 10.6151
R885 B.n211 B.n210 10.6151
R886 B.n212 B.n211 10.6151
R887 B.n212 B.n115 10.6151
R888 B.n216 B.n115 10.6151
R889 B.n217 B.n216 10.6151
R890 B.n218 B.n217 10.6151
R891 B.n218 B.n113 10.6151
R892 B.n222 B.n113 10.6151
R893 B.n223 B.n222 10.6151
R894 B.n224 B.n223 10.6151
R895 B.n224 B.n111 10.6151
R896 B.n228 B.n111 10.6151
R897 B.n229 B.n228 10.6151
R898 B.n231 B.n107 10.6151
R899 B.n235 B.n107 10.6151
R900 B.n236 B.n235 10.6151
R901 B.n237 B.n236 10.6151
R902 B.n237 B.n105 10.6151
R903 B.n241 B.n105 10.6151
R904 B.n242 B.n241 10.6151
R905 B.n246 B.n242 10.6151
R906 B.n250 B.n103 10.6151
R907 B.n251 B.n250 10.6151
R908 B.n252 B.n251 10.6151
R909 B.n252 B.n101 10.6151
R910 B.n256 B.n101 10.6151
R911 B.n257 B.n256 10.6151
R912 B.n258 B.n257 10.6151
R913 B.n258 B.n99 10.6151
R914 B.n262 B.n99 10.6151
R915 B.n263 B.n262 10.6151
R916 B.n264 B.n263 10.6151
R917 B.n264 B.n97 10.6151
R918 B.n268 B.n97 10.6151
R919 B.n269 B.n268 10.6151
R920 B.n270 B.n269 10.6151
R921 B.n270 B.n95 10.6151
R922 B.n274 B.n95 10.6151
R923 B.n275 B.n274 10.6151
R924 B.n276 B.n275 10.6151
R925 B.n276 B.n93 10.6151
R926 B.n280 B.n93 10.6151
R927 B.n281 B.n280 10.6151
R928 B.n282 B.n281 10.6151
R929 B.n282 B.n91 10.6151
R930 B.n286 B.n91 10.6151
R931 B.n287 B.n286 10.6151
R932 B.n288 B.n287 10.6151
R933 B.n288 B.n89 10.6151
R934 B.n292 B.n89 10.6151
R935 B.n293 B.n292 10.6151
R936 B.n294 B.n293 10.6151
R937 B.n294 B.n87 10.6151
R938 B.n298 B.n87 10.6151
R939 B.n299 B.n298 10.6151
R940 B.n176 B.n175 10.6151
R941 B.n175 B.n174 10.6151
R942 B.n174 B.n129 10.6151
R943 B.n170 B.n129 10.6151
R944 B.n170 B.n169 10.6151
R945 B.n169 B.n168 10.6151
R946 B.n168 B.n131 10.6151
R947 B.n164 B.n131 10.6151
R948 B.n164 B.n163 10.6151
R949 B.n163 B.n162 10.6151
R950 B.n162 B.n133 10.6151
R951 B.n158 B.n133 10.6151
R952 B.n158 B.n157 10.6151
R953 B.n157 B.n156 10.6151
R954 B.n156 B.n135 10.6151
R955 B.n152 B.n135 10.6151
R956 B.n152 B.n151 10.6151
R957 B.n151 B.n150 10.6151
R958 B.n150 B.n137 10.6151
R959 B.n146 B.n137 10.6151
R960 B.n146 B.n145 10.6151
R961 B.n145 B.n144 10.6151
R962 B.n144 B.n139 10.6151
R963 B.n140 B.n139 10.6151
R964 B.n140 B.n0 10.6151
R965 B.n535 B.n1 10.6151
R966 B.n535 B.n534 10.6151
R967 B.n534 B.n533 10.6151
R968 B.n533 B.n4 10.6151
R969 B.n529 B.n4 10.6151
R970 B.n529 B.n528 10.6151
R971 B.n528 B.n527 10.6151
R972 B.n527 B.n6 10.6151
R973 B.n523 B.n6 10.6151
R974 B.n523 B.n522 10.6151
R975 B.n522 B.n521 10.6151
R976 B.n521 B.n8 10.6151
R977 B.n517 B.n8 10.6151
R978 B.n517 B.n516 10.6151
R979 B.n516 B.n515 10.6151
R980 B.n515 B.n10 10.6151
R981 B.n511 B.n10 10.6151
R982 B.n511 B.n510 10.6151
R983 B.n510 B.n509 10.6151
R984 B.n509 B.n12 10.6151
R985 B.n505 B.n12 10.6151
R986 B.n505 B.n504 10.6151
R987 B.n504 B.n503 10.6151
R988 B.n503 B.n14 10.6151
R989 B.n499 B.n14 10.6151
R990 B.n445 B.n36 6.5566
R991 B.n433 B.n432 6.5566
R992 B.n231 B.n230 6.5566
R993 B.n246 B.n245 6.5566
R994 B.n36 B.n32 4.05904
R995 B.n432 B.n431 4.05904
R996 B.n230 B.n229 4.05904
R997 B.n245 B.n103 4.05904
R998 B.n539 B.n0 2.81026
R999 B.n539 B.n1 2.81026
C0 VTAIL VP 5.36637f
C1 B VN 0.768279f
C2 VDD2 B 1.57211f
C3 B w_n2194_n2898# 6.67855f
C4 B VDD1 1.52822f
C5 VN VP 5.14895f
C6 VDD2 VP 0.339545f
C7 w_n2194_n2898# VP 4.35988f
C8 VP VDD1 5.61672f
C9 VTAIL VN 5.35185f
C10 VDD2 VTAIL 12.028701f
C11 VTAIL w_n2194_n2898# 2.63439f
C12 VTAIL VDD1 11.993299f
C13 B VP 1.22817f
C14 VDD2 VN 5.42967f
C15 w_n2194_n2898# VN 4.08013f
C16 VN VDD1 0.148591f
C17 VTAIL B 2.30719f
C18 VDD2 w_n2194_n2898# 1.90099f
C19 VDD2 VDD1 0.962755f
C20 w_n2194_n2898# VDD1 1.8569f
C21 VDD2 VSUBS 1.299713f
C22 VDD1 VSUBS 1.079027f
C23 VTAIL VSUBS 0.700217f
C24 VN VSUBS 4.7451f
C25 VP VSUBS 1.716407f
C26 B VSUBS 2.799472f
C27 w_n2194_n2898# VSUBS 78.589096f
C28 B.n0 VSUBS 0.004842f
C29 B.n1 VSUBS 0.004842f
C30 B.n2 VSUBS 0.007657f
C31 B.n3 VSUBS 0.007657f
C32 B.n4 VSUBS 0.007657f
C33 B.n5 VSUBS 0.007657f
C34 B.n6 VSUBS 0.007657f
C35 B.n7 VSUBS 0.007657f
C36 B.n8 VSUBS 0.007657f
C37 B.n9 VSUBS 0.007657f
C38 B.n10 VSUBS 0.007657f
C39 B.n11 VSUBS 0.007657f
C40 B.n12 VSUBS 0.007657f
C41 B.n13 VSUBS 0.007657f
C42 B.n14 VSUBS 0.007657f
C43 B.n15 VSUBS 0.018747f
C44 B.n16 VSUBS 0.007657f
C45 B.n17 VSUBS 0.007657f
C46 B.n18 VSUBS 0.007657f
C47 B.n19 VSUBS 0.007657f
C48 B.n20 VSUBS 0.007657f
C49 B.n21 VSUBS 0.007657f
C50 B.n22 VSUBS 0.007657f
C51 B.n23 VSUBS 0.007657f
C52 B.n24 VSUBS 0.007657f
C53 B.n25 VSUBS 0.007657f
C54 B.n26 VSUBS 0.007657f
C55 B.n27 VSUBS 0.007657f
C56 B.n28 VSUBS 0.007657f
C57 B.n29 VSUBS 0.007657f
C58 B.n30 VSUBS 0.007657f
C59 B.n31 VSUBS 0.007657f
C60 B.n32 VSUBS 0.005293f
C61 B.n33 VSUBS 0.007657f
C62 B.t5 VSUBS 0.335072f
C63 B.t4 VSUBS 0.344003f
C64 B.t3 VSUBS 0.304386f
C65 B.n34 VSUBS 0.126409f
C66 B.n35 VSUBS 0.06966f
C67 B.n36 VSUBS 0.017742f
C68 B.n37 VSUBS 0.007657f
C69 B.n38 VSUBS 0.007657f
C70 B.n39 VSUBS 0.007657f
C71 B.n40 VSUBS 0.007657f
C72 B.t2 VSUBS 0.335067f
C73 B.t1 VSUBS 0.343998f
C74 B.t0 VSUBS 0.304386f
C75 B.n41 VSUBS 0.126413f
C76 B.n42 VSUBS 0.069664f
C77 B.n43 VSUBS 0.007657f
C78 B.n44 VSUBS 0.007657f
C79 B.n45 VSUBS 0.007657f
C80 B.n46 VSUBS 0.007657f
C81 B.n47 VSUBS 0.007657f
C82 B.n48 VSUBS 0.007657f
C83 B.n49 VSUBS 0.007657f
C84 B.n50 VSUBS 0.007657f
C85 B.n51 VSUBS 0.007657f
C86 B.n52 VSUBS 0.007657f
C87 B.n53 VSUBS 0.007657f
C88 B.n54 VSUBS 0.007657f
C89 B.n55 VSUBS 0.007657f
C90 B.n56 VSUBS 0.007657f
C91 B.n57 VSUBS 0.007657f
C92 B.n58 VSUBS 0.007657f
C93 B.n59 VSUBS 0.017867f
C94 B.n60 VSUBS 0.007657f
C95 B.n61 VSUBS 0.007657f
C96 B.n62 VSUBS 0.007657f
C97 B.n63 VSUBS 0.007657f
C98 B.n64 VSUBS 0.007657f
C99 B.n65 VSUBS 0.007657f
C100 B.n66 VSUBS 0.007657f
C101 B.n67 VSUBS 0.007657f
C102 B.n68 VSUBS 0.007657f
C103 B.n69 VSUBS 0.007657f
C104 B.n70 VSUBS 0.007657f
C105 B.n71 VSUBS 0.007657f
C106 B.n72 VSUBS 0.007657f
C107 B.n73 VSUBS 0.007657f
C108 B.n74 VSUBS 0.007657f
C109 B.n75 VSUBS 0.007657f
C110 B.n76 VSUBS 0.007657f
C111 B.n77 VSUBS 0.007657f
C112 B.n78 VSUBS 0.007657f
C113 B.n79 VSUBS 0.007657f
C114 B.n80 VSUBS 0.007657f
C115 B.n81 VSUBS 0.007657f
C116 B.n82 VSUBS 0.007657f
C117 B.n83 VSUBS 0.007657f
C118 B.n84 VSUBS 0.007657f
C119 B.n85 VSUBS 0.007657f
C120 B.n86 VSUBS 0.018747f
C121 B.n87 VSUBS 0.007657f
C122 B.n88 VSUBS 0.007657f
C123 B.n89 VSUBS 0.007657f
C124 B.n90 VSUBS 0.007657f
C125 B.n91 VSUBS 0.007657f
C126 B.n92 VSUBS 0.007657f
C127 B.n93 VSUBS 0.007657f
C128 B.n94 VSUBS 0.007657f
C129 B.n95 VSUBS 0.007657f
C130 B.n96 VSUBS 0.007657f
C131 B.n97 VSUBS 0.007657f
C132 B.n98 VSUBS 0.007657f
C133 B.n99 VSUBS 0.007657f
C134 B.n100 VSUBS 0.007657f
C135 B.n101 VSUBS 0.007657f
C136 B.n102 VSUBS 0.007657f
C137 B.n103 VSUBS 0.005293f
C138 B.n104 VSUBS 0.007657f
C139 B.n105 VSUBS 0.007657f
C140 B.n106 VSUBS 0.007657f
C141 B.n107 VSUBS 0.007657f
C142 B.n108 VSUBS 0.007657f
C143 B.t7 VSUBS 0.335072f
C144 B.t8 VSUBS 0.344003f
C145 B.t6 VSUBS 0.304386f
C146 B.n109 VSUBS 0.126409f
C147 B.n110 VSUBS 0.06966f
C148 B.n111 VSUBS 0.007657f
C149 B.n112 VSUBS 0.007657f
C150 B.n113 VSUBS 0.007657f
C151 B.n114 VSUBS 0.007657f
C152 B.n115 VSUBS 0.007657f
C153 B.n116 VSUBS 0.007657f
C154 B.n117 VSUBS 0.007657f
C155 B.n118 VSUBS 0.007657f
C156 B.n119 VSUBS 0.007657f
C157 B.n120 VSUBS 0.007657f
C158 B.n121 VSUBS 0.007657f
C159 B.n122 VSUBS 0.007657f
C160 B.n123 VSUBS 0.007657f
C161 B.n124 VSUBS 0.007657f
C162 B.n125 VSUBS 0.007657f
C163 B.n126 VSUBS 0.007657f
C164 B.n127 VSUBS 0.018747f
C165 B.n128 VSUBS 0.007657f
C166 B.n129 VSUBS 0.007657f
C167 B.n130 VSUBS 0.007657f
C168 B.n131 VSUBS 0.007657f
C169 B.n132 VSUBS 0.007657f
C170 B.n133 VSUBS 0.007657f
C171 B.n134 VSUBS 0.007657f
C172 B.n135 VSUBS 0.007657f
C173 B.n136 VSUBS 0.007657f
C174 B.n137 VSUBS 0.007657f
C175 B.n138 VSUBS 0.007657f
C176 B.n139 VSUBS 0.007657f
C177 B.n140 VSUBS 0.007657f
C178 B.n141 VSUBS 0.007657f
C179 B.n142 VSUBS 0.007657f
C180 B.n143 VSUBS 0.007657f
C181 B.n144 VSUBS 0.007657f
C182 B.n145 VSUBS 0.007657f
C183 B.n146 VSUBS 0.007657f
C184 B.n147 VSUBS 0.007657f
C185 B.n148 VSUBS 0.007657f
C186 B.n149 VSUBS 0.007657f
C187 B.n150 VSUBS 0.007657f
C188 B.n151 VSUBS 0.007657f
C189 B.n152 VSUBS 0.007657f
C190 B.n153 VSUBS 0.007657f
C191 B.n154 VSUBS 0.007657f
C192 B.n155 VSUBS 0.007657f
C193 B.n156 VSUBS 0.007657f
C194 B.n157 VSUBS 0.007657f
C195 B.n158 VSUBS 0.007657f
C196 B.n159 VSUBS 0.007657f
C197 B.n160 VSUBS 0.007657f
C198 B.n161 VSUBS 0.007657f
C199 B.n162 VSUBS 0.007657f
C200 B.n163 VSUBS 0.007657f
C201 B.n164 VSUBS 0.007657f
C202 B.n165 VSUBS 0.007657f
C203 B.n166 VSUBS 0.007657f
C204 B.n167 VSUBS 0.007657f
C205 B.n168 VSUBS 0.007657f
C206 B.n169 VSUBS 0.007657f
C207 B.n170 VSUBS 0.007657f
C208 B.n171 VSUBS 0.007657f
C209 B.n172 VSUBS 0.007657f
C210 B.n173 VSUBS 0.007657f
C211 B.n174 VSUBS 0.007657f
C212 B.n175 VSUBS 0.007657f
C213 B.n176 VSUBS 0.017738f
C214 B.n177 VSUBS 0.017738f
C215 B.n178 VSUBS 0.018747f
C216 B.n179 VSUBS 0.007657f
C217 B.n180 VSUBS 0.007657f
C218 B.n181 VSUBS 0.007657f
C219 B.n182 VSUBS 0.007657f
C220 B.n183 VSUBS 0.007657f
C221 B.n184 VSUBS 0.007657f
C222 B.n185 VSUBS 0.007657f
C223 B.n186 VSUBS 0.007657f
C224 B.n187 VSUBS 0.007657f
C225 B.n188 VSUBS 0.007657f
C226 B.n189 VSUBS 0.007657f
C227 B.n190 VSUBS 0.007657f
C228 B.n191 VSUBS 0.007657f
C229 B.n192 VSUBS 0.007657f
C230 B.n193 VSUBS 0.007657f
C231 B.n194 VSUBS 0.007657f
C232 B.n195 VSUBS 0.007657f
C233 B.n196 VSUBS 0.007657f
C234 B.n197 VSUBS 0.007657f
C235 B.n198 VSUBS 0.007657f
C236 B.n199 VSUBS 0.007657f
C237 B.n200 VSUBS 0.007657f
C238 B.n201 VSUBS 0.007657f
C239 B.n202 VSUBS 0.007657f
C240 B.n203 VSUBS 0.007657f
C241 B.n204 VSUBS 0.007657f
C242 B.n205 VSUBS 0.007657f
C243 B.n206 VSUBS 0.007657f
C244 B.n207 VSUBS 0.007657f
C245 B.n208 VSUBS 0.007657f
C246 B.n209 VSUBS 0.007657f
C247 B.n210 VSUBS 0.007657f
C248 B.n211 VSUBS 0.007657f
C249 B.n212 VSUBS 0.007657f
C250 B.n213 VSUBS 0.007657f
C251 B.n214 VSUBS 0.007657f
C252 B.n215 VSUBS 0.007657f
C253 B.n216 VSUBS 0.007657f
C254 B.n217 VSUBS 0.007657f
C255 B.n218 VSUBS 0.007657f
C256 B.n219 VSUBS 0.007657f
C257 B.n220 VSUBS 0.007657f
C258 B.n221 VSUBS 0.007657f
C259 B.n222 VSUBS 0.007657f
C260 B.n223 VSUBS 0.007657f
C261 B.n224 VSUBS 0.007657f
C262 B.n225 VSUBS 0.007657f
C263 B.n226 VSUBS 0.007657f
C264 B.n227 VSUBS 0.007657f
C265 B.n228 VSUBS 0.007657f
C266 B.n229 VSUBS 0.005293f
C267 B.n230 VSUBS 0.017742f
C268 B.n231 VSUBS 0.006194f
C269 B.n232 VSUBS 0.007657f
C270 B.n233 VSUBS 0.007657f
C271 B.n234 VSUBS 0.007657f
C272 B.n235 VSUBS 0.007657f
C273 B.n236 VSUBS 0.007657f
C274 B.n237 VSUBS 0.007657f
C275 B.n238 VSUBS 0.007657f
C276 B.n239 VSUBS 0.007657f
C277 B.n240 VSUBS 0.007657f
C278 B.n241 VSUBS 0.007657f
C279 B.n242 VSUBS 0.007657f
C280 B.t10 VSUBS 0.335067f
C281 B.t11 VSUBS 0.343998f
C282 B.t9 VSUBS 0.304386f
C283 B.n243 VSUBS 0.126413f
C284 B.n244 VSUBS 0.069664f
C285 B.n245 VSUBS 0.017742f
C286 B.n246 VSUBS 0.006194f
C287 B.n247 VSUBS 0.007657f
C288 B.n248 VSUBS 0.007657f
C289 B.n249 VSUBS 0.007657f
C290 B.n250 VSUBS 0.007657f
C291 B.n251 VSUBS 0.007657f
C292 B.n252 VSUBS 0.007657f
C293 B.n253 VSUBS 0.007657f
C294 B.n254 VSUBS 0.007657f
C295 B.n255 VSUBS 0.007657f
C296 B.n256 VSUBS 0.007657f
C297 B.n257 VSUBS 0.007657f
C298 B.n258 VSUBS 0.007657f
C299 B.n259 VSUBS 0.007657f
C300 B.n260 VSUBS 0.007657f
C301 B.n261 VSUBS 0.007657f
C302 B.n262 VSUBS 0.007657f
C303 B.n263 VSUBS 0.007657f
C304 B.n264 VSUBS 0.007657f
C305 B.n265 VSUBS 0.007657f
C306 B.n266 VSUBS 0.007657f
C307 B.n267 VSUBS 0.007657f
C308 B.n268 VSUBS 0.007657f
C309 B.n269 VSUBS 0.007657f
C310 B.n270 VSUBS 0.007657f
C311 B.n271 VSUBS 0.007657f
C312 B.n272 VSUBS 0.007657f
C313 B.n273 VSUBS 0.007657f
C314 B.n274 VSUBS 0.007657f
C315 B.n275 VSUBS 0.007657f
C316 B.n276 VSUBS 0.007657f
C317 B.n277 VSUBS 0.007657f
C318 B.n278 VSUBS 0.007657f
C319 B.n279 VSUBS 0.007657f
C320 B.n280 VSUBS 0.007657f
C321 B.n281 VSUBS 0.007657f
C322 B.n282 VSUBS 0.007657f
C323 B.n283 VSUBS 0.007657f
C324 B.n284 VSUBS 0.007657f
C325 B.n285 VSUBS 0.007657f
C326 B.n286 VSUBS 0.007657f
C327 B.n287 VSUBS 0.007657f
C328 B.n288 VSUBS 0.007657f
C329 B.n289 VSUBS 0.007657f
C330 B.n290 VSUBS 0.007657f
C331 B.n291 VSUBS 0.007657f
C332 B.n292 VSUBS 0.007657f
C333 B.n293 VSUBS 0.007657f
C334 B.n294 VSUBS 0.007657f
C335 B.n295 VSUBS 0.007657f
C336 B.n296 VSUBS 0.007657f
C337 B.n297 VSUBS 0.007657f
C338 B.n298 VSUBS 0.007657f
C339 B.n299 VSUBS 0.018747f
C340 B.n300 VSUBS 0.017738f
C341 B.n301 VSUBS 0.017738f
C342 B.n302 VSUBS 0.007657f
C343 B.n303 VSUBS 0.007657f
C344 B.n304 VSUBS 0.007657f
C345 B.n305 VSUBS 0.007657f
C346 B.n306 VSUBS 0.007657f
C347 B.n307 VSUBS 0.007657f
C348 B.n308 VSUBS 0.007657f
C349 B.n309 VSUBS 0.007657f
C350 B.n310 VSUBS 0.007657f
C351 B.n311 VSUBS 0.007657f
C352 B.n312 VSUBS 0.007657f
C353 B.n313 VSUBS 0.007657f
C354 B.n314 VSUBS 0.007657f
C355 B.n315 VSUBS 0.007657f
C356 B.n316 VSUBS 0.007657f
C357 B.n317 VSUBS 0.007657f
C358 B.n318 VSUBS 0.007657f
C359 B.n319 VSUBS 0.007657f
C360 B.n320 VSUBS 0.007657f
C361 B.n321 VSUBS 0.007657f
C362 B.n322 VSUBS 0.007657f
C363 B.n323 VSUBS 0.007657f
C364 B.n324 VSUBS 0.007657f
C365 B.n325 VSUBS 0.007657f
C366 B.n326 VSUBS 0.007657f
C367 B.n327 VSUBS 0.007657f
C368 B.n328 VSUBS 0.007657f
C369 B.n329 VSUBS 0.007657f
C370 B.n330 VSUBS 0.007657f
C371 B.n331 VSUBS 0.007657f
C372 B.n332 VSUBS 0.007657f
C373 B.n333 VSUBS 0.007657f
C374 B.n334 VSUBS 0.007657f
C375 B.n335 VSUBS 0.007657f
C376 B.n336 VSUBS 0.007657f
C377 B.n337 VSUBS 0.007657f
C378 B.n338 VSUBS 0.007657f
C379 B.n339 VSUBS 0.007657f
C380 B.n340 VSUBS 0.007657f
C381 B.n341 VSUBS 0.007657f
C382 B.n342 VSUBS 0.007657f
C383 B.n343 VSUBS 0.007657f
C384 B.n344 VSUBS 0.007657f
C385 B.n345 VSUBS 0.007657f
C386 B.n346 VSUBS 0.007657f
C387 B.n347 VSUBS 0.007657f
C388 B.n348 VSUBS 0.007657f
C389 B.n349 VSUBS 0.007657f
C390 B.n350 VSUBS 0.007657f
C391 B.n351 VSUBS 0.007657f
C392 B.n352 VSUBS 0.007657f
C393 B.n353 VSUBS 0.007657f
C394 B.n354 VSUBS 0.007657f
C395 B.n355 VSUBS 0.007657f
C396 B.n356 VSUBS 0.007657f
C397 B.n357 VSUBS 0.007657f
C398 B.n358 VSUBS 0.007657f
C399 B.n359 VSUBS 0.007657f
C400 B.n360 VSUBS 0.007657f
C401 B.n361 VSUBS 0.007657f
C402 B.n362 VSUBS 0.007657f
C403 B.n363 VSUBS 0.007657f
C404 B.n364 VSUBS 0.007657f
C405 B.n365 VSUBS 0.007657f
C406 B.n366 VSUBS 0.007657f
C407 B.n367 VSUBS 0.007657f
C408 B.n368 VSUBS 0.007657f
C409 B.n369 VSUBS 0.007657f
C410 B.n370 VSUBS 0.007657f
C411 B.n371 VSUBS 0.007657f
C412 B.n372 VSUBS 0.007657f
C413 B.n373 VSUBS 0.007657f
C414 B.n374 VSUBS 0.007657f
C415 B.n375 VSUBS 0.007657f
C416 B.n376 VSUBS 0.007657f
C417 B.n377 VSUBS 0.007657f
C418 B.n378 VSUBS 0.018619f
C419 B.n379 VSUBS 0.017738f
C420 B.n380 VSUBS 0.018747f
C421 B.n381 VSUBS 0.007657f
C422 B.n382 VSUBS 0.007657f
C423 B.n383 VSUBS 0.007657f
C424 B.n384 VSUBS 0.007657f
C425 B.n385 VSUBS 0.007657f
C426 B.n386 VSUBS 0.007657f
C427 B.n387 VSUBS 0.007657f
C428 B.n388 VSUBS 0.007657f
C429 B.n389 VSUBS 0.007657f
C430 B.n390 VSUBS 0.007657f
C431 B.n391 VSUBS 0.007657f
C432 B.n392 VSUBS 0.007657f
C433 B.n393 VSUBS 0.007657f
C434 B.n394 VSUBS 0.007657f
C435 B.n395 VSUBS 0.007657f
C436 B.n396 VSUBS 0.007657f
C437 B.n397 VSUBS 0.007657f
C438 B.n398 VSUBS 0.007657f
C439 B.n399 VSUBS 0.007657f
C440 B.n400 VSUBS 0.007657f
C441 B.n401 VSUBS 0.007657f
C442 B.n402 VSUBS 0.007657f
C443 B.n403 VSUBS 0.007657f
C444 B.n404 VSUBS 0.007657f
C445 B.n405 VSUBS 0.007657f
C446 B.n406 VSUBS 0.007657f
C447 B.n407 VSUBS 0.007657f
C448 B.n408 VSUBS 0.007657f
C449 B.n409 VSUBS 0.007657f
C450 B.n410 VSUBS 0.007657f
C451 B.n411 VSUBS 0.007657f
C452 B.n412 VSUBS 0.007657f
C453 B.n413 VSUBS 0.007657f
C454 B.n414 VSUBS 0.007657f
C455 B.n415 VSUBS 0.007657f
C456 B.n416 VSUBS 0.007657f
C457 B.n417 VSUBS 0.007657f
C458 B.n418 VSUBS 0.007657f
C459 B.n419 VSUBS 0.007657f
C460 B.n420 VSUBS 0.007657f
C461 B.n421 VSUBS 0.007657f
C462 B.n422 VSUBS 0.007657f
C463 B.n423 VSUBS 0.007657f
C464 B.n424 VSUBS 0.007657f
C465 B.n425 VSUBS 0.007657f
C466 B.n426 VSUBS 0.007657f
C467 B.n427 VSUBS 0.007657f
C468 B.n428 VSUBS 0.007657f
C469 B.n429 VSUBS 0.007657f
C470 B.n430 VSUBS 0.007657f
C471 B.n431 VSUBS 0.005293f
C472 B.n432 VSUBS 0.017742f
C473 B.n433 VSUBS 0.006194f
C474 B.n434 VSUBS 0.007657f
C475 B.n435 VSUBS 0.007657f
C476 B.n436 VSUBS 0.007657f
C477 B.n437 VSUBS 0.007657f
C478 B.n438 VSUBS 0.007657f
C479 B.n439 VSUBS 0.007657f
C480 B.n440 VSUBS 0.007657f
C481 B.n441 VSUBS 0.007657f
C482 B.n442 VSUBS 0.007657f
C483 B.n443 VSUBS 0.007657f
C484 B.n444 VSUBS 0.007657f
C485 B.n445 VSUBS 0.006194f
C486 B.n446 VSUBS 0.007657f
C487 B.n447 VSUBS 0.007657f
C488 B.n448 VSUBS 0.007657f
C489 B.n449 VSUBS 0.007657f
C490 B.n450 VSUBS 0.007657f
C491 B.n451 VSUBS 0.007657f
C492 B.n452 VSUBS 0.007657f
C493 B.n453 VSUBS 0.007657f
C494 B.n454 VSUBS 0.007657f
C495 B.n455 VSUBS 0.007657f
C496 B.n456 VSUBS 0.007657f
C497 B.n457 VSUBS 0.007657f
C498 B.n458 VSUBS 0.007657f
C499 B.n459 VSUBS 0.007657f
C500 B.n460 VSUBS 0.007657f
C501 B.n461 VSUBS 0.007657f
C502 B.n462 VSUBS 0.007657f
C503 B.n463 VSUBS 0.007657f
C504 B.n464 VSUBS 0.007657f
C505 B.n465 VSUBS 0.007657f
C506 B.n466 VSUBS 0.007657f
C507 B.n467 VSUBS 0.007657f
C508 B.n468 VSUBS 0.007657f
C509 B.n469 VSUBS 0.007657f
C510 B.n470 VSUBS 0.007657f
C511 B.n471 VSUBS 0.007657f
C512 B.n472 VSUBS 0.007657f
C513 B.n473 VSUBS 0.007657f
C514 B.n474 VSUBS 0.007657f
C515 B.n475 VSUBS 0.007657f
C516 B.n476 VSUBS 0.007657f
C517 B.n477 VSUBS 0.007657f
C518 B.n478 VSUBS 0.007657f
C519 B.n479 VSUBS 0.007657f
C520 B.n480 VSUBS 0.007657f
C521 B.n481 VSUBS 0.007657f
C522 B.n482 VSUBS 0.007657f
C523 B.n483 VSUBS 0.007657f
C524 B.n484 VSUBS 0.007657f
C525 B.n485 VSUBS 0.007657f
C526 B.n486 VSUBS 0.007657f
C527 B.n487 VSUBS 0.007657f
C528 B.n488 VSUBS 0.007657f
C529 B.n489 VSUBS 0.007657f
C530 B.n490 VSUBS 0.007657f
C531 B.n491 VSUBS 0.007657f
C532 B.n492 VSUBS 0.007657f
C533 B.n493 VSUBS 0.007657f
C534 B.n494 VSUBS 0.007657f
C535 B.n495 VSUBS 0.007657f
C536 B.n496 VSUBS 0.007657f
C537 B.n497 VSUBS 0.007657f
C538 B.n498 VSUBS 0.018747f
C539 B.n499 VSUBS 0.017738f
C540 B.n500 VSUBS 0.017738f
C541 B.n501 VSUBS 0.007657f
C542 B.n502 VSUBS 0.007657f
C543 B.n503 VSUBS 0.007657f
C544 B.n504 VSUBS 0.007657f
C545 B.n505 VSUBS 0.007657f
C546 B.n506 VSUBS 0.007657f
C547 B.n507 VSUBS 0.007657f
C548 B.n508 VSUBS 0.007657f
C549 B.n509 VSUBS 0.007657f
C550 B.n510 VSUBS 0.007657f
C551 B.n511 VSUBS 0.007657f
C552 B.n512 VSUBS 0.007657f
C553 B.n513 VSUBS 0.007657f
C554 B.n514 VSUBS 0.007657f
C555 B.n515 VSUBS 0.007657f
C556 B.n516 VSUBS 0.007657f
C557 B.n517 VSUBS 0.007657f
C558 B.n518 VSUBS 0.007657f
C559 B.n519 VSUBS 0.007657f
C560 B.n520 VSUBS 0.007657f
C561 B.n521 VSUBS 0.007657f
C562 B.n522 VSUBS 0.007657f
C563 B.n523 VSUBS 0.007657f
C564 B.n524 VSUBS 0.007657f
C565 B.n525 VSUBS 0.007657f
C566 B.n526 VSUBS 0.007657f
C567 B.n527 VSUBS 0.007657f
C568 B.n528 VSUBS 0.007657f
C569 B.n529 VSUBS 0.007657f
C570 B.n530 VSUBS 0.007657f
C571 B.n531 VSUBS 0.007657f
C572 B.n532 VSUBS 0.007657f
C573 B.n533 VSUBS 0.007657f
C574 B.n534 VSUBS 0.007657f
C575 B.n535 VSUBS 0.007657f
C576 B.n536 VSUBS 0.007657f
C577 B.n537 VSUBS 0.007657f
C578 B.n538 VSUBS 0.007657f
C579 B.n539 VSUBS 0.017339f
C580 VDD2.t7 VSUBS 1.84649f
C581 VDD2.t4 VSUBS 0.186629f
C582 VDD2.t8 VSUBS 0.186629f
C583 VDD2.n0 VSUBS 1.402f
C584 VDD2.n1 VSUBS 1.10163f
C585 VDD2.t5 VSUBS 0.186629f
C586 VDD2.t9 VSUBS 0.186629f
C587 VDD2.n2 VSUBS 1.40629f
C588 VDD2.n3 VSUBS 1.95255f
C589 VDD2.t0 VSUBS 1.8403f
C590 VDD2.n4 VSUBS 2.39432f
C591 VDD2.t1 VSUBS 0.186629f
C592 VDD2.t2 VSUBS 0.186629f
C593 VDD2.n5 VSUBS 1.402f
C594 VDD2.n6 VSUBS 0.527347f
C595 VDD2.t3 VSUBS 0.186629f
C596 VDD2.t6 VSUBS 0.186629f
C597 VDD2.n7 VSUBS 1.40626f
C598 VN.n0 VSUBS 0.054185f
C599 VN.n1 VSUBS 0.012296f
C600 VN.n2 VSUBS 0.224665f
C601 VN.t2 VSUBS 1.05627f
C602 VN.n3 VSUBS 0.410831f
C603 VN.t5 VSUBS 1.03346f
C604 VN.n4 VSUBS 0.433898f
C605 VN.n5 VSUBS 0.012296f
C606 VN.t1 VSUBS 1.03346f
C607 VN.n6 VSUBS 0.428994f
C608 VN.n7 VSUBS 0.054185f
C609 VN.n8 VSUBS 0.054185f
C610 VN.n9 VSUBS 0.054185f
C611 VN.t4 VSUBS 1.03346f
C612 VN.n10 VSUBS 0.428994f
C613 VN.n11 VSUBS 0.012296f
C614 VN.t0 VSUBS 1.03346f
C615 VN.n12 VSUBS 0.425153f
C616 VN.n13 VSUBS 0.041991f
C617 VN.n14 VSUBS 0.054185f
C618 VN.n15 VSUBS 0.012296f
C619 VN.t8 VSUBS 1.03346f
C620 VN.n16 VSUBS 0.224665f
C621 VN.t3 VSUBS 1.05627f
C622 VN.n17 VSUBS 0.410831f
C623 VN.t6 VSUBS 1.03346f
C624 VN.n18 VSUBS 0.433898f
C625 VN.n19 VSUBS 0.012296f
C626 VN.t7 VSUBS 1.03346f
C627 VN.n20 VSUBS 0.428994f
C628 VN.n21 VSUBS 0.054185f
C629 VN.n22 VSUBS 0.054185f
C630 VN.n23 VSUBS 0.054185f
C631 VN.n24 VSUBS 0.428994f
C632 VN.n25 VSUBS 0.012296f
C633 VN.t9 VSUBS 1.03346f
C634 VN.n26 VSUBS 0.425153f
C635 VN.n27 VSUBS 2.17746f
C636 VDD1.t6 VSUBS 1.85807f
C637 VDD1.t3 VSUBS 0.187799f
C638 VDD1.t2 VSUBS 0.187799f
C639 VDD1.n0 VSUBS 1.41079f
C640 VDD1.n1 VSUBS 1.11406f
C641 VDD1.t7 VSUBS 1.85806f
C642 VDD1.t4 VSUBS 0.187799f
C643 VDD1.t8 VSUBS 0.187799f
C644 VDD1.n2 VSUBS 1.41078f
C645 VDD1.n3 VSUBS 1.10853f
C646 VDD1.t5 VSUBS 0.187799f
C647 VDD1.t9 VSUBS 0.187799f
C648 VDD1.n4 VSUBS 1.4151f
C649 VDD1.n5 VSUBS 2.03961f
C650 VDD1.t1 VSUBS 0.187799f
C651 VDD1.t0 VSUBS 0.187799f
C652 VDD1.n6 VSUBS 1.41078f
C653 VDD1.n7 VSUBS 2.40204f
C654 VTAIL.t4 VSUBS 0.228353f
C655 VTAIL.t8 VSUBS 0.228353f
C656 VTAIL.n0 VSUBS 1.57368f
C657 VTAIL.n1 VSUBS 0.791634f
C658 VTAIL.t12 VSUBS 2.09522f
C659 VTAIL.n2 VSUBS 0.908479f
C660 VTAIL.t11 VSUBS 0.228353f
C661 VTAIL.t16 VSUBS 0.228353f
C662 VTAIL.n3 VSUBS 1.57368f
C663 VTAIL.n4 VSUBS 0.804319f
C664 VTAIL.t18 VSUBS 0.228353f
C665 VTAIL.t13 VSUBS 0.228353f
C666 VTAIL.n5 VSUBS 1.57368f
C667 VTAIL.n6 VSUBS 2.09863f
C668 VTAIL.t3 VSUBS 0.228353f
C669 VTAIL.t5 VSUBS 0.228353f
C670 VTAIL.n7 VSUBS 1.57369f
C671 VTAIL.n8 VSUBS 2.09862f
C672 VTAIL.t1 VSUBS 0.228353f
C673 VTAIL.t9 VSUBS 0.228353f
C674 VTAIL.n9 VSUBS 1.57369f
C675 VTAIL.n10 VSUBS 0.804312f
C676 VTAIL.t7 VSUBS 2.09523f
C677 VTAIL.n11 VSUBS 0.908464f
C678 VTAIL.t17 VSUBS 0.228353f
C679 VTAIL.t19 VSUBS 0.228353f
C680 VTAIL.n12 VSUBS 1.57369f
C681 VTAIL.n13 VSUBS 0.807224f
C682 VTAIL.t14 VSUBS 0.228353f
C683 VTAIL.t15 VSUBS 0.228353f
C684 VTAIL.n14 VSUBS 1.57369f
C685 VTAIL.n15 VSUBS 0.804312f
C686 VTAIL.t10 VSUBS 2.09522f
C687 VTAIL.n16 VSUBS 2.11503f
C688 VTAIL.t6 VSUBS 2.09522f
C689 VTAIL.n17 VSUBS 2.11503f
C690 VTAIL.t2 VSUBS 0.228353f
C691 VTAIL.t0 VSUBS 0.228353f
C692 VTAIL.n18 VSUBS 1.57368f
C693 VTAIL.n19 VSUBS 0.73507f
C694 VP.n0 VSUBS 0.055752f
C695 VP.n1 VSUBS 0.012651f
C696 VP.n2 VSUBS 0.055752f
C697 VP.n3 VSUBS 0.012651f
C698 VP.n4 VSUBS 0.055752f
C699 VP.t9 VSUBS 1.06335f
C700 VP.t8 VSUBS 1.06335f
C701 VP.n5 VSUBS 0.055752f
C702 VP.t7 VSUBS 1.06335f
C703 VP.n6 VSUBS 0.4414f
C704 VP.t3 VSUBS 1.08682f
C705 VP.n7 VSUBS 0.422712f
C706 VP.t6 VSUBS 1.06335f
C707 VP.n8 VSUBS 0.446446f
C708 VP.n9 VSUBS 0.012651f
C709 VP.n10 VSUBS 0.231163f
C710 VP.n11 VSUBS 0.055752f
C711 VP.n12 VSUBS 0.055752f
C712 VP.n13 VSUBS 0.012651f
C713 VP.n14 VSUBS 0.4414f
C714 VP.n15 VSUBS 0.012651f
C715 VP.n16 VSUBS 0.437447f
C716 VP.n17 VSUBS 2.20377f
C717 VP.t2 VSUBS 1.06335f
C718 VP.n18 VSUBS 0.437447f
C719 VP.n19 VSUBS 2.25273f
C720 VP.n20 VSUBS 0.055752f
C721 VP.n21 VSUBS 0.055752f
C722 VP.t5 VSUBS 1.06335f
C723 VP.n22 VSUBS 0.4414f
C724 VP.n23 VSUBS 0.012651f
C725 VP.t1 VSUBS 1.06335f
C726 VP.n24 VSUBS 0.4414f
C727 VP.n25 VSUBS 0.055752f
C728 VP.n26 VSUBS 0.055752f
C729 VP.n27 VSUBS 0.055752f
C730 VP.t4 VSUBS 1.06335f
C731 VP.n28 VSUBS 0.4414f
C732 VP.n29 VSUBS 0.012651f
C733 VP.t0 VSUBS 1.06335f
C734 VP.n30 VSUBS 0.437447f
C735 VP.n31 VSUBS 0.043206f
.ends

