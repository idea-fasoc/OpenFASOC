* NGSPICE file created from diff_pair_sample_0818.ext - technology: sky130A

.subckt diff_pair_sample_0818 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=3.0987 ps=19.11 w=18.78 l=0.68
X1 VDD1.t3 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0987 pd=19.11 as=7.3242 ps=38.34 w=18.78 l=0.68
X2 VTAIL.t6 VN.t1 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=3.0987 ps=19.11 w=18.78 l=0.68
X3 VDD2.t2 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.0987 pd=19.11 as=7.3242 ps=38.34 w=18.78 l=0.68
X4 VTAIL.t1 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=3.0987 ps=19.11 w=18.78 l=0.68
X5 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0987 pd=19.11 as=7.3242 ps=38.34 w=18.78 l=0.68
X6 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=0.68
X7 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=0.68
X8 VDD2.t3 VN.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.0987 pd=19.11 as=7.3242 ps=38.34 w=18.78 l=0.68
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=0.68
X10 VTAIL.t2 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=3.0987 ps=19.11 w=18.78 l=0.68
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.3242 pd=38.34 as=0 ps=0 w=18.78 l=0.68
R0 VN.n0 VN.t0 745.061
R1 VN.n1 VN.t3 745.061
R2 VN.n0 VN.t2 745.01
R3 VN.n1 VN.t1 745.01
R4 VN VN.n1 90.5125
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 106.175
R7 VDD2.n2 VDD2.n1 63.6588
R8 VDD2.n1 VDD2.t1 1.05481
R9 VDD2.n1 VDD2.t3 1.05481
R10 VDD2.n0 VDD2.t0 1.05481
R11 VDD2.n0 VDD2.t2 1.05481
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n830 VTAIL.n829 289.615
R14 VTAIL.n102 VTAIL.n101 289.615
R15 VTAIL.n206 VTAIL.n205 289.615
R16 VTAIL.n310 VTAIL.n309 289.615
R17 VTAIL.n726 VTAIL.n725 289.615
R18 VTAIL.n622 VTAIL.n621 289.615
R19 VTAIL.n518 VTAIL.n517 289.615
R20 VTAIL.n414 VTAIL.n413 289.615
R21 VTAIL.n763 VTAIL.n762 185
R22 VTAIL.n765 VTAIL.n764 185
R23 VTAIL.n758 VTAIL.n757 185
R24 VTAIL.n771 VTAIL.n770 185
R25 VTAIL.n773 VTAIL.n772 185
R26 VTAIL.n754 VTAIL.n753 185
R27 VTAIL.n780 VTAIL.n779 185
R28 VTAIL.n781 VTAIL.n752 185
R29 VTAIL.n783 VTAIL.n782 185
R30 VTAIL.n750 VTAIL.n749 185
R31 VTAIL.n789 VTAIL.n788 185
R32 VTAIL.n791 VTAIL.n790 185
R33 VTAIL.n746 VTAIL.n745 185
R34 VTAIL.n797 VTAIL.n796 185
R35 VTAIL.n799 VTAIL.n798 185
R36 VTAIL.n742 VTAIL.n741 185
R37 VTAIL.n805 VTAIL.n804 185
R38 VTAIL.n807 VTAIL.n806 185
R39 VTAIL.n738 VTAIL.n737 185
R40 VTAIL.n813 VTAIL.n812 185
R41 VTAIL.n815 VTAIL.n814 185
R42 VTAIL.n734 VTAIL.n733 185
R43 VTAIL.n821 VTAIL.n820 185
R44 VTAIL.n823 VTAIL.n822 185
R45 VTAIL.n730 VTAIL.n729 185
R46 VTAIL.n829 VTAIL.n828 185
R47 VTAIL.n35 VTAIL.n34 185
R48 VTAIL.n37 VTAIL.n36 185
R49 VTAIL.n30 VTAIL.n29 185
R50 VTAIL.n43 VTAIL.n42 185
R51 VTAIL.n45 VTAIL.n44 185
R52 VTAIL.n26 VTAIL.n25 185
R53 VTAIL.n52 VTAIL.n51 185
R54 VTAIL.n53 VTAIL.n24 185
R55 VTAIL.n55 VTAIL.n54 185
R56 VTAIL.n22 VTAIL.n21 185
R57 VTAIL.n61 VTAIL.n60 185
R58 VTAIL.n63 VTAIL.n62 185
R59 VTAIL.n18 VTAIL.n17 185
R60 VTAIL.n69 VTAIL.n68 185
R61 VTAIL.n71 VTAIL.n70 185
R62 VTAIL.n14 VTAIL.n13 185
R63 VTAIL.n77 VTAIL.n76 185
R64 VTAIL.n79 VTAIL.n78 185
R65 VTAIL.n10 VTAIL.n9 185
R66 VTAIL.n85 VTAIL.n84 185
R67 VTAIL.n87 VTAIL.n86 185
R68 VTAIL.n6 VTAIL.n5 185
R69 VTAIL.n93 VTAIL.n92 185
R70 VTAIL.n95 VTAIL.n94 185
R71 VTAIL.n2 VTAIL.n1 185
R72 VTAIL.n101 VTAIL.n100 185
R73 VTAIL.n139 VTAIL.n138 185
R74 VTAIL.n141 VTAIL.n140 185
R75 VTAIL.n134 VTAIL.n133 185
R76 VTAIL.n147 VTAIL.n146 185
R77 VTAIL.n149 VTAIL.n148 185
R78 VTAIL.n130 VTAIL.n129 185
R79 VTAIL.n156 VTAIL.n155 185
R80 VTAIL.n157 VTAIL.n128 185
R81 VTAIL.n159 VTAIL.n158 185
R82 VTAIL.n126 VTAIL.n125 185
R83 VTAIL.n165 VTAIL.n164 185
R84 VTAIL.n167 VTAIL.n166 185
R85 VTAIL.n122 VTAIL.n121 185
R86 VTAIL.n173 VTAIL.n172 185
R87 VTAIL.n175 VTAIL.n174 185
R88 VTAIL.n118 VTAIL.n117 185
R89 VTAIL.n181 VTAIL.n180 185
R90 VTAIL.n183 VTAIL.n182 185
R91 VTAIL.n114 VTAIL.n113 185
R92 VTAIL.n189 VTAIL.n188 185
R93 VTAIL.n191 VTAIL.n190 185
R94 VTAIL.n110 VTAIL.n109 185
R95 VTAIL.n197 VTAIL.n196 185
R96 VTAIL.n199 VTAIL.n198 185
R97 VTAIL.n106 VTAIL.n105 185
R98 VTAIL.n205 VTAIL.n204 185
R99 VTAIL.n243 VTAIL.n242 185
R100 VTAIL.n245 VTAIL.n244 185
R101 VTAIL.n238 VTAIL.n237 185
R102 VTAIL.n251 VTAIL.n250 185
R103 VTAIL.n253 VTAIL.n252 185
R104 VTAIL.n234 VTAIL.n233 185
R105 VTAIL.n260 VTAIL.n259 185
R106 VTAIL.n261 VTAIL.n232 185
R107 VTAIL.n263 VTAIL.n262 185
R108 VTAIL.n230 VTAIL.n229 185
R109 VTAIL.n269 VTAIL.n268 185
R110 VTAIL.n271 VTAIL.n270 185
R111 VTAIL.n226 VTAIL.n225 185
R112 VTAIL.n277 VTAIL.n276 185
R113 VTAIL.n279 VTAIL.n278 185
R114 VTAIL.n222 VTAIL.n221 185
R115 VTAIL.n285 VTAIL.n284 185
R116 VTAIL.n287 VTAIL.n286 185
R117 VTAIL.n218 VTAIL.n217 185
R118 VTAIL.n293 VTAIL.n292 185
R119 VTAIL.n295 VTAIL.n294 185
R120 VTAIL.n214 VTAIL.n213 185
R121 VTAIL.n301 VTAIL.n300 185
R122 VTAIL.n303 VTAIL.n302 185
R123 VTAIL.n210 VTAIL.n209 185
R124 VTAIL.n309 VTAIL.n308 185
R125 VTAIL.n725 VTAIL.n724 185
R126 VTAIL.n626 VTAIL.n625 185
R127 VTAIL.n719 VTAIL.n718 185
R128 VTAIL.n717 VTAIL.n716 185
R129 VTAIL.n630 VTAIL.n629 185
R130 VTAIL.n711 VTAIL.n710 185
R131 VTAIL.n709 VTAIL.n708 185
R132 VTAIL.n634 VTAIL.n633 185
R133 VTAIL.n703 VTAIL.n702 185
R134 VTAIL.n701 VTAIL.n700 185
R135 VTAIL.n638 VTAIL.n637 185
R136 VTAIL.n695 VTAIL.n694 185
R137 VTAIL.n693 VTAIL.n692 185
R138 VTAIL.n642 VTAIL.n641 185
R139 VTAIL.n687 VTAIL.n686 185
R140 VTAIL.n685 VTAIL.n684 185
R141 VTAIL.n646 VTAIL.n645 185
R142 VTAIL.n650 VTAIL.n648 185
R143 VTAIL.n679 VTAIL.n678 185
R144 VTAIL.n677 VTAIL.n676 185
R145 VTAIL.n652 VTAIL.n651 185
R146 VTAIL.n671 VTAIL.n670 185
R147 VTAIL.n669 VTAIL.n668 185
R148 VTAIL.n656 VTAIL.n655 185
R149 VTAIL.n663 VTAIL.n662 185
R150 VTAIL.n661 VTAIL.n660 185
R151 VTAIL.n621 VTAIL.n620 185
R152 VTAIL.n522 VTAIL.n521 185
R153 VTAIL.n615 VTAIL.n614 185
R154 VTAIL.n613 VTAIL.n612 185
R155 VTAIL.n526 VTAIL.n525 185
R156 VTAIL.n607 VTAIL.n606 185
R157 VTAIL.n605 VTAIL.n604 185
R158 VTAIL.n530 VTAIL.n529 185
R159 VTAIL.n599 VTAIL.n598 185
R160 VTAIL.n597 VTAIL.n596 185
R161 VTAIL.n534 VTAIL.n533 185
R162 VTAIL.n591 VTAIL.n590 185
R163 VTAIL.n589 VTAIL.n588 185
R164 VTAIL.n538 VTAIL.n537 185
R165 VTAIL.n583 VTAIL.n582 185
R166 VTAIL.n581 VTAIL.n580 185
R167 VTAIL.n542 VTAIL.n541 185
R168 VTAIL.n546 VTAIL.n544 185
R169 VTAIL.n575 VTAIL.n574 185
R170 VTAIL.n573 VTAIL.n572 185
R171 VTAIL.n548 VTAIL.n547 185
R172 VTAIL.n567 VTAIL.n566 185
R173 VTAIL.n565 VTAIL.n564 185
R174 VTAIL.n552 VTAIL.n551 185
R175 VTAIL.n559 VTAIL.n558 185
R176 VTAIL.n557 VTAIL.n556 185
R177 VTAIL.n517 VTAIL.n516 185
R178 VTAIL.n418 VTAIL.n417 185
R179 VTAIL.n511 VTAIL.n510 185
R180 VTAIL.n509 VTAIL.n508 185
R181 VTAIL.n422 VTAIL.n421 185
R182 VTAIL.n503 VTAIL.n502 185
R183 VTAIL.n501 VTAIL.n500 185
R184 VTAIL.n426 VTAIL.n425 185
R185 VTAIL.n495 VTAIL.n494 185
R186 VTAIL.n493 VTAIL.n492 185
R187 VTAIL.n430 VTAIL.n429 185
R188 VTAIL.n487 VTAIL.n486 185
R189 VTAIL.n485 VTAIL.n484 185
R190 VTAIL.n434 VTAIL.n433 185
R191 VTAIL.n479 VTAIL.n478 185
R192 VTAIL.n477 VTAIL.n476 185
R193 VTAIL.n438 VTAIL.n437 185
R194 VTAIL.n442 VTAIL.n440 185
R195 VTAIL.n471 VTAIL.n470 185
R196 VTAIL.n469 VTAIL.n468 185
R197 VTAIL.n444 VTAIL.n443 185
R198 VTAIL.n463 VTAIL.n462 185
R199 VTAIL.n461 VTAIL.n460 185
R200 VTAIL.n448 VTAIL.n447 185
R201 VTAIL.n455 VTAIL.n454 185
R202 VTAIL.n453 VTAIL.n452 185
R203 VTAIL.n413 VTAIL.n412 185
R204 VTAIL.n314 VTAIL.n313 185
R205 VTAIL.n407 VTAIL.n406 185
R206 VTAIL.n405 VTAIL.n404 185
R207 VTAIL.n318 VTAIL.n317 185
R208 VTAIL.n399 VTAIL.n398 185
R209 VTAIL.n397 VTAIL.n396 185
R210 VTAIL.n322 VTAIL.n321 185
R211 VTAIL.n391 VTAIL.n390 185
R212 VTAIL.n389 VTAIL.n388 185
R213 VTAIL.n326 VTAIL.n325 185
R214 VTAIL.n383 VTAIL.n382 185
R215 VTAIL.n381 VTAIL.n380 185
R216 VTAIL.n330 VTAIL.n329 185
R217 VTAIL.n375 VTAIL.n374 185
R218 VTAIL.n373 VTAIL.n372 185
R219 VTAIL.n334 VTAIL.n333 185
R220 VTAIL.n338 VTAIL.n336 185
R221 VTAIL.n367 VTAIL.n366 185
R222 VTAIL.n365 VTAIL.n364 185
R223 VTAIL.n340 VTAIL.n339 185
R224 VTAIL.n359 VTAIL.n358 185
R225 VTAIL.n357 VTAIL.n356 185
R226 VTAIL.n344 VTAIL.n343 185
R227 VTAIL.n351 VTAIL.n350 185
R228 VTAIL.n349 VTAIL.n348 185
R229 VTAIL.n761 VTAIL.t5 149.524
R230 VTAIL.n33 VTAIL.t7 149.524
R231 VTAIL.n137 VTAIL.t3 149.524
R232 VTAIL.n241 VTAIL.t2 149.524
R233 VTAIL.n659 VTAIL.t0 149.524
R234 VTAIL.n555 VTAIL.t1 149.524
R235 VTAIL.n451 VTAIL.t4 149.524
R236 VTAIL.n347 VTAIL.t6 149.524
R237 VTAIL.n764 VTAIL.n763 104.615
R238 VTAIL.n764 VTAIL.n757 104.615
R239 VTAIL.n771 VTAIL.n757 104.615
R240 VTAIL.n772 VTAIL.n771 104.615
R241 VTAIL.n772 VTAIL.n753 104.615
R242 VTAIL.n780 VTAIL.n753 104.615
R243 VTAIL.n781 VTAIL.n780 104.615
R244 VTAIL.n782 VTAIL.n781 104.615
R245 VTAIL.n782 VTAIL.n749 104.615
R246 VTAIL.n789 VTAIL.n749 104.615
R247 VTAIL.n790 VTAIL.n789 104.615
R248 VTAIL.n790 VTAIL.n745 104.615
R249 VTAIL.n797 VTAIL.n745 104.615
R250 VTAIL.n798 VTAIL.n797 104.615
R251 VTAIL.n798 VTAIL.n741 104.615
R252 VTAIL.n805 VTAIL.n741 104.615
R253 VTAIL.n806 VTAIL.n805 104.615
R254 VTAIL.n806 VTAIL.n737 104.615
R255 VTAIL.n813 VTAIL.n737 104.615
R256 VTAIL.n814 VTAIL.n813 104.615
R257 VTAIL.n814 VTAIL.n733 104.615
R258 VTAIL.n821 VTAIL.n733 104.615
R259 VTAIL.n822 VTAIL.n821 104.615
R260 VTAIL.n822 VTAIL.n729 104.615
R261 VTAIL.n829 VTAIL.n729 104.615
R262 VTAIL.n36 VTAIL.n35 104.615
R263 VTAIL.n36 VTAIL.n29 104.615
R264 VTAIL.n43 VTAIL.n29 104.615
R265 VTAIL.n44 VTAIL.n43 104.615
R266 VTAIL.n44 VTAIL.n25 104.615
R267 VTAIL.n52 VTAIL.n25 104.615
R268 VTAIL.n53 VTAIL.n52 104.615
R269 VTAIL.n54 VTAIL.n53 104.615
R270 VTAIL.n54 VTAIL.n21 104.615
R271 VTAIL.n61 VTAIL.n21 104.615
R272 VTAIL.n62 VTAIL.n61 104.615
R273 VTAIL.n62 VTAIL.n17 104.615
R274 VTAIL.n69 VTAIL.n17 104.615
R275 VTAIL.n70 VTAIL.n69 104.615
R276 VTAIL.n70 VTAIL.n13 104.615
R277 VTAIL.n77 VTAIL.n13 104.615
R278 VTAIL.n78 VTAIL.n77 104.615
R279 VTAIL.n78 VTAIL.n9 104.615
R280 VTAIL.n85 VTAIL.n9 104.615
R281 VTAIL.n86 VTAIL.n85 104.615
R282 VTAIL.n86 VTAIL.n5 104.615
R283 VTAIL.n93 VTAIL.n5 104.615
R284 VTAIL.n94 VTAIL.n93 104.615
R285 VTAIL.n94 VTAIL.n1 104.615
R286 VTAIL.n101 VTAIL.n1 104.615
R287 VTAIL.n140 VTAIL.n139 104.615
R288 VTAIL.n140 VTAIL.n133 104.615
R289 VTAIL.n147 VTAIL.n133 104.615
R290 VTAIL.n148 VTAIL.n147 104.615
R291 VTAIL.n148 VTAIL.n129 104.615
R292 VTAIL.n156 VTAIL.n129 104.615
R293 VTAIL.n157 VTAIL.n156 104.615
R294 VTAIL.n158 VTAIL.n157 104.615
R295 VTAIL.n158 VTAIL.n125 104.615
R296 VTAIL.n165 VTAIL.n125 104.615
R297 VTAIL.n166 VTAIL.n165 104.615
R298 VTAIL.n166 VTAIL.n121 104.615
R299 VTAIL.n173 VTAIL.n121 104.615
R300 VTAIL.n174 VTAIL.n173 104.615
R301 VTAIL.n174 VTAIL.n117 104.615
R302 VTAIL.n181 VTAIL.n117 104.615
R303 VTAIL.n182 VTAIL.n181 104.615
R304 VTAIL.n182 VTAIL.n113 104.615
R305 VTAIL.n189 VTAIL.n113 104.615
R306 VTAIL.n190 VTAIL.n189 104.615
R307 VTAIL.n190 VTAIL.n109 104.615
R308 VTAIL.n197 VTAIL.n109 104.615
R309 VTAIL.n198 VTAIL.n197 104.615
R310 VTAIL.n198 VTAIL.n105 104.615
R311 VTAIL.n205 VTAIL.n105 104.615
R312 VTAIL.n244 VTAIL.n243 104.615
R313 VTAIL.n244 VTAIL.n237 104.615
R314 VTAIL.n251 VTAIL.n237 104.615
R315 VTAIL.n252 VTAIL.n251 104.615
R316 VTAIL.n252 VTAIL.n233 104.615
R317 VTAIL.n260 VTAIL.n233 104.615
R318 VTAIL.n261 VTAIL.n260 104.615
R319 VTAIL.n262 VTAIL.n261 104.615
R320 VTAIL.n262 VTAIL.n229 104.615
R321 VTAIL.n269 VTAIL.n229 104.615
R322 VTAIL.n270 VTAIL.n269 104.615
R323 VTAIL.n270 VTAIL.n225 104.615
R324 VTAIL.n277 VTAIL.n225 104.615
R325 VTAIL.n278 VTAIL.n277 104.615
R326 VTAIL.n278 VTAIL.n221 104.615
R327 VTAIL.n285 VTAIL.n221 104.615
R328 VTAIL.n286 VTAIL.n285 104.615
R329 VTAIL.n286 VTAIL.n217 104.615
R330 VTAIL.n293 VTAIL.n217 104.615
R331 VTAIL.n294 VTAIL.n293 104.615
R332 VTAIL.n294 VTAIL.n213 104.615
R333 VTAIL.n301 VTAIL.n213 104.615
R334 VTAIL.n302 VTAIL.n301 104.615
R335 VTAIL.n302 VTAIL.n209 104.615
R336 VTAIL.n309 VTAIL.n209 104.615
R337 VTAIL.n725 VTAIL.n625 104.615
R338 VTAIL.n718 VTAIL.n625 104.615
R339 VTAIL.n718 VTAIL.n717 104.615
R340 VTAIL.n717 VTAIL.n629 104.615
R341 VTAIL.n710 VTAIL.n629 104.615
R342 VTAIL.n710 VTAIL.n709 104.615
R343 VTAIL.n709 VTAIL.n633 104.615
R344 VTAIL.n702 VTAIL.n633 104.615
R345 VTAIL.n702 VTAIL.n701 104.615
R346 VTAIL.n701 VTAIL.n637 104.615
R347 VTAIL.n694 VTAIL.n637 104.615
R348 VTAIL.n694 VTAIL.n693 104.615
R349 VTAIL.n693 VTAIL.n641 104.615
R350 VTAIL.n686 VTAIL.n641 104.615
R351 VTAIL.n686 VTAIL.n685 104.615
R352 VTAIL.n685 VTAIL.n645 104.615
R353 VTAIL.n650 VTAIL.n645 104.615
R354 VTAIL.n678 VTAIL.n650 104.615
R355 VTAIL.n678 VTAIL.n677 104.615
R356 VTAIL.n677 VTAIL.n651 104.615
R357 VTAIL.n670 VTAIL.n651 104.615
R358 VTAIL.n670 VTAIL.n669 104.615
R359 VTAIL.n669 VTAIL.n655 104.615
R360 VTAIL.n662 VTAIL.n655 104.615
R361 VTAIL.n662 VTAIL.n661 104.615
R362 VTAIL.n621 VTAIL.n521 104.615
R363 VTAIL.n614 VTAIL.n521 104.615
R364 VTAIL.n614 VTAIL.n613 104.615
R365 VTAIL.n613 VTAIL.n525 104.615
R366 VTAIL.n606 VTAIL.n525 104.615
R367 VTAIL.n606 VTAIL.n605 104.615
R368 VTAIL.n605 VTAIL.n529 104.615
R369 VTAIL.n598 VTAIL.n529 104.615
R370 VTAIL.n598 VTAIL.n597 104.615
R371 VTAIL.n597 VTAIL.n533 104.615
R372 VTAIL.n590 VTAIL.n533 104.615
R373 VTAIL.n590 VTAIL.n589 104.615
R374 VTAIL.n589 VTAIL.n537 104.615
R375 VTAIL.n582 VTAIL.n537 104.615
R376 VTAIL.n582 VTAIL.n581 104.615
R377 VTAIL.n581 VTAIL.n541 104.615
R378 VTAIL.n546 VTAIL.n541 104.615
R379 VTAIL.n574 VTAIL.n546 104.615
R380 VTAIL.n574 VTAIL.n573 104.615
R381 VTAIL.n573 VTAIL.n547 104.615
R382 VTAIL.n566 VTAIL.n547 104.615
R383 VTAIL.n566 VTAIL.n565 104.615
R384 VTAIL.n565 VTAIL.n551 104.615
R385 VTAIL.n558 VTAIL.n551 104.615
R386 VTAIL.n558 VTAIL.n557 104.615
R387 VTAIL.n517 VTAIL.n417 104.615
R388 VTAIL.n510 VTAIL.n417 104.615
R389 VTAIL.n510 VTAIL.n509 104.615
R390 VTAIL.n509 VTAIL.n421 104.615
R391 VTAIL.n502 VTAIL.n421 104.615
R392 VTAIL.n502 VTAIL.n501 104.615
R393 VTAIL.n501 VTAIL.n425 104.615
R394 VTAIL.n494 VTAIL.n425 104.615
R395 VTAIL.n494 VTAIL.n493 104.615
R396 VTAIL.n493 VTAIL.n429 104.615
R397 VTAIL.n486 VTAIL.n429 104.615
R398 VTAIL.n486 VTAIL.n485 104.615
R399 VTAIL.n485 VTAIL.n433 104.615
R400 VTAIL.n478 VTAIL.n433 104.615
R401 VTAIL.n478 VTAIL.n477 104.615
R402 VTAIL.n477 VTAIL.n437 104.615
R403 VTAIL.n442 VTAIL.n437 104.615
R404 VTAIL.n470 VTAIL.n442 104.615
R405 VTAIL.n470 VTAIL.n469 104.615
R406 VTAIL.n469 VTAIL.n443 104.615
R407 VTAIL.n462 VTAIL.n443 104.615
R408 VTAIL.n462 VTAIL.n461 104.615
R409 VTAIL.n461 VTAIL.n447 104.615
R410 VTAIL.n454 VTAIL.n447 104.615
R411 VTAIL.n454 VTAIL.n453 104.615
R412 VTAIL.n413 VTAIL.n313 104.615
R413 VTAIL.n406 VTAIL.n313 104.615
R414 VTAIL.n406 VTAIL.n405 104.615
R415 VTAIL.n405 VTAIL.n317 104.615
R416 VTAIL.n398 VTAIL.n317 104.615
R417 VTAIL.n398 VTAIL.n397 104.615
R418 VTAIL.n397 VTAIL.n321 104.615
R419 VTAIL.n390 VTAIL.n321 104.615
R420 VTAIL.n390 VTAIL.n389 104.615
R421 VTAIL.n389 VTAIL.n325 104.615
R422 VTAIL.n382 VTAIL.n325 104.615
R423 VTAIL.n382 VTAIL.n381 104.615
R424 VTAIL.n381 VTAIL.n329 104.615
R425 VTAIL.n374 VTAIL.n329 104.615
R426 VTAIL.n374 VTAIL.n373 104.615
R427 VTAIL.n373 VTAIL.n333 104.615
R428 VTAIL.n338 VTAIL.n333 104.615
R429 VTAIL.n366 VTAIL.n338 104.615
R430 VTAIL.n366 VTAIL.n365 104.615
R431 VTAIL.n365 VTAIL.n339 104.615
R432 VTAIL.n358 VTAIL.n339 104.615
R433 VTAIL.n358 VTAIL.n357 104.615
R434 VTAIL.n357 VTAIL.n343 104.615
R435 VTAIL.n350 VTAIL.n343 104.615
R436 VTAIL.n350 VTAIL.n349 104.615
R437 VTAIL.n763 VTAIL.t5 52.3082
R438 VTAIL.n35 VTAIL.t7 52.3082
R439 VTAIL.n139 VTAIL.t3 52.3082
R440 VTAIL.n243 VTAIL.t2 52.3082
R441 VTAIL.n661 VTAIL.t0 52.3082
R442 VTAIL.n557 VTAIL.t1 52.3082
R443 VTAIL.n453 VTAIL.t4 52.3082
R444 VTAIL.n349 VTAIL.t6 52.3082
R445 VTAIL.n831 VTAIL.n830 35.2884
R446 VTAIL.n103 VTAIL.n102 35.2884
R447 VTAIL.n207 VTAIL.n206 35.2884
R448 VTAIL.n311 VTAIL.n310 35.2884
R449 VTAIL.n727 VTAIL.n726 35.2884
R450 VTAIL.n623 VTAIL.n622 35.2884
R451 VTAIL.n519 VTAIL.n518 35.2884
R452 VTAIL.n415 VTAIL.n414 35.2884
R453 VTAIL.n831 VTAIL.n727 29.4272
R454 VTAIL.n415 VTAIL.n311 29.4272
R455 VTAIL.n783 VTAIL.n750 13.1884
R456 VTAIL.n55 VTAIL.n22 13.1884
R457 VTAIL.n159 VTAIL.n126 13.1884
R458 VTAIL.n263 VTAIL.n230 13.1884
R459 VTAIL.n648 VTAIL.n646 13.1884
R460 VTAIL.n544 VTAIL.n542 13.1884
R461 VTAIL.n440 VTAIL.n438 13.1884
R462 VTAIL.n336 VTAIL.n334 13.1884
R463 VTAIL.n784 VTAIL.n752 12.8005
R464 VTAIL.n788 VTAIL.n787 12.8005
R465 VTAIL.n828 VTAIL.n728 12.8005
R466 VTAIL.n56 VTAIL.n24 12.8005
R467 VTAIL.n60 VTAIL.n59 12.8005
R468 VTAIL.n100 VTAIL.n0 12.8005
R469 VTAIL.n160 VTAIL.n128 12.8005
R470 VTAIL.n164 VTAIL.n163 12.8005
R471 VTAIL.n204 VTAIL.n104 12.8005
R472 VTAIL.n264 VTAIL.n232 12.8005
R473 VTAIL.n268 VTAIL.n267 12.8005
R474 VTAIL.n308 VTAIL.n208 12.8005
R475 VTAIL.n724 VTAIL.n624 12.8005
R476 VTAIL.n684 VTAIL.n683 12.8005
R477 VTAIL.n680 VTAIL.n679 12.8005
R478 VTAIL.n620 VTAIL.n520 12.8005
R479 VTAIL.n580 VTAIL.n579 12.8005
R480 VTAIL.n576 VTAIL.n575 12.8005
R481 VTAIL.n516 VTAIL.n416 12.8005
R482 VTAIL.n476 VTAIL.n475 12.8005
R483 VTAIL.n472 VTAIL.n471 12.8005
R484 VTAIL.n412 VTAIL.n312 12.8005
R485 VTAIL.n372 VTAIL.n371 12.8005
R486 VTAIL.n368 VTAIL.n367 12.8005
R487 VTAIL.n779 VTAIL.n778 12.0247
R488 VTAIL.n791 VTAIL.n748 12.0247
R489 VTAIL.n827 VTAIL.n730 12.0247
R490 VTAIL.n51 VTAIL.n50 12.0247
R491 VTAIL.n63 VTAIL.n20 12.0247
R492 VTAIL.n99 VTAIL.n2 12.0247
R493 VTAIL.n155 VTAIL.n154 12.0247
R494 VTAIL.n167 VTAIL.n124 12.0247
R495 VTAIL.n203 VTAIL.n106 12.0247
R496 VTAIL.n259 VTAIL.n258 12.0247
R497 VTAIL.n271 VTAIL.n228 12.0247
R498 VTAIL.n307 VTAIL.n210 12.0247
R499 VTAIL.n723 VTAIL.n626 12.0247
R500 VTAIL.n687 VTAIL.n644 12.0247
R501 VTAIL.n676 VTAIL.n649 12.0247
R502 VTAIL.n619 VTAIL.n522 12.0247
R503 VTAIL.n583 VTAIL.n540 12.0247
R504 VTAIL.n572 VTAIL.n545 12.0247
R505 VTAIL.n515 VTAIL.n418 12.0247
R506 VTAIL.n479 VTAIL.n436 12.0247
R507 VTAIL.n468 VTAIL.n441 12.0247
R508 VTAIL.n411 VTAIL.n314 12.0247
R509 VTAIL.n375 VTAIL.n332 12.0247
R510 VTAIL.n364 VTAIL.n337 12.0247
R511 VTAIL.n777 VTAIL.n754 11.249
R512 VTAIL.n792 VTAIL.n746 11.249
R513 VTAIL.n824 VTAIL.n823 11.249
R514 VTAIL.n49 VTAIL.n26 11.249
R515 VTAIL.n64 VTAIL.n18 11.249
R516 VTAIL.n96 VTAIL.n95 11.249
R517 VTAIL.n153 VTAIL.n130 11.249
R518 VTAIL.n168 VTAIL.n122 11.249
R519 VTAIL.n200 VTAIL.n199 11.249
R520 VTAIL.n257 VTAIL.n234 11.249
R521 VTAIL.n272 VTAIL.n226 11.249
R522 VTAIL.n304 VTAIL.n303 11.249
R523 VTAIL.n720 VTAIL.n719 11.249
R524 VTAIL.n688 VTAIL.n642 11.249
R525 VTAIL.n675 VTAIL.n652 11.249
R526 VTAIL.n616 VTAIL.n615 11.249
R527 VTAIL.n584 VTAIL.n538 11.249
R528 VTAIL.n571 VTAIL.n548 11.249
R529 VTAIL.n512 VTAIL.n511 11.249
R530 VTAIL.n480 VTAIL.n434 11.249
R531 VTAIL.n467 VTAIL.n444 11.249
R532 VTAIL.n408 VTAIL.n407 11.249
R533 VTAIL.n376 VTAIL.n330 11.249
R534 VTAIL.n363 VTAIL.n340 11.249
R535 VTAIL.n774 VTAIL.n773 10.4732
R536 VTAIL.n796 VTAIL.n795 10.4732
R537 VTAIL.n820 VTAIL.n732 10.4732
R538 VTAIL.n46 VTAIL.n45 10.4732
R539 VTAIL.n68 VTAIL.n67 10.4732
R540 VTAIL.n92 VTAIL.n4 10.4732
R541 VTAIL.n150 VTAIL.n149 10.4732
R542 VTAIL.n172 VTAIL.n171 10.4732
R543 VTAIL.n196 VTAIL.n108 10.4732
R544 VTAIL.n254 VTAIL.n253 10.4732
R545 VTAIL.n276 VTAIL.n275 10.4732
R546 VTAIL.n300 VTAIL.n212 10.4732
R547 VTAIL.n716 VTAIL.n628 10.4732
R548 VTAIL.n692 VTAIL.n691 10.4732
R549 VTAIL.n672 VTAIL.n671 10.4732
R550 VTAIL.n612 VTAIL.n524 10.4732
R551 VTAIL.n588 VTAIL.n587 10.4732
R552 VTAIL.n568 VTAIL.n567 10.4732
R553 VTAIL.n508 VTAIL.n420 10.4732
R554 VTAIL.n484 VTAIL.n483 10.4732
R555 VTAIL.n464 VTAIL.n463 10.4732
R556 VTAIL.n404 VTAIL.n316 10.4732
R557 VTAIL.n380 VTAIL.n379 10.4732
R558 VTAIL.n360 VTAIL.n359 10.4732
R559 VTAIL.n762 VTAIL.n761 10.2747
R560 VTAIL.n34 VTAIL.n33 10.2747
R561 VTAIL.n138 VTAIL.n137 10.2747
R562 VTAIL.n242 VTAIL.n241 10.2747
R563 VTAIL.n660 VTAIL.n659 10.2747
R564 VTAIL.n556 VTAIL.n555 10.2747
R565 VTAIL.n452 VTAIL.n451 10.2747
R566 VTAIL.n348 VTAIL.n347 10.2747
R567 VTAIL.n770 VTAIL.n756 9.69747
R568 VTAIL.n799 VTAIL.n744 9.69747
R569 VTAIL.n819 VTAIL.n734 9.69747
R570 VTAIL.n42 VTAIL.n28 9.69747
R571 VTAIL.n71 VTAIL.n16 9.69747
R572 VTAIL.n91 VTAIL.n6 9.69747
R573 VTAIL.n146 VTAIL.n132 9.69747
R574 VTAIL.n175 VTAIL.n120 9.69747
R575 VTAIL.n195 VTAIL.n110 9.69747
R576 VTAIL.n250 VTAIL.n236 9.69747
R577 VTAIL.n279 VTAIL.n224 9.69747
R578 VTAIL.n299 VTAIL.n214 9.69747
R579 VTAIL.n715 VTAIL.n630 9.69747
R580 VTAIL.n695 VTAIL.n640 9.69747
R581 VTAIL.n668 VTAIL.n654 9.69747
R582 VTAIL.n611 VTAIL.n526 9.69747
R583 VTAIL.n591 VTAIL.n536 9.69747
R584 VTAIL.n564 VTAIL.n550 9.69747
R585 VTAIL.n507 VTAIL.n422 9.69747
R586 VTAIL.n487 VTAIL.n432 9.69747
R587 VTAIL.n460 VTAIL.n446 9.69747
R588 VTAIL.n403 VTAIL.n318 9.69747
R589 VTAIL.n383 VTAIL.n328 9.69747
R590 VTAIL.n356 VTAIL.n342 9.69747
R591 VTAIL.n826 VTAIL.n728 9.45567
R592 VTAIL.n98 VTAIL.n0 9.45567
R593 VTAIL.n202 VTAIL.n104 9.45567
R594 VTAIL.n306 VTAIL.n208 9.45567
R595 VTAIL.n722 VTAIL.n624 9.45567
R596 VTAIL.n618 VTAIL.n520 9.45567
R597 VTAIL.n514 VTAIL.n416 9.45567
R598 VTAIL.n410 VTAIL.n312 9.45567
R599 VTAIL.n809 VTAIL.n808 9.3005
R600 VTAIL.n811 VTAIL.n810 9.3005
R601 VTAIL.n736 VTAIL.n735 9.3005
R602 VTAIL.n817 VTAIL.n816 9.3005
R603 VTAIL.n819 VTAIL.n818 9.3005
R604 VTAIL.n732 VTAIL.n731 9.3005
R605 VTAIL.n825 VTAIL.n824 9.3005
R606 VTAIL.n827 VTAIL.n826 9.3005
R607 VTAIL.n803 VTAIL.n802 9.3005
R608 VTAIL.n801 VTAIL.n800 9.3005
R609 VTAIL.n744 VTAIL.n743 9.3005
R610 VTAIL.n795 VTAIL.n794 9.3005
R611 VTAIL.n793 VTAIL.n792 9.3005
R612 VTAIL.n748 VTAIL.n747 9.3005
R613 VTAIL.n787 VTAIL.n786 9.3005
R614 VTAIL.n760 VTAIL.n759 9.3005
R615 VTAIL.n767 VTAIL.n766 9.3005
R616 VTAIL.n769 VTAIL.n768 9.3005
R617 VTAIL.n756 VTAIL.n755 9.3005
R618 VTAIL.n775 VTAIL.n774 9.3005
R619 VTAIL.n777 VTAIL.n776 9.3005
R620 VTAIL.n778 VTAIL.n751 9.3005
R621 VTAIL.n785 VTAIL.n784 9.3005
R622 VTAIL.n740 VTAIL.n739 9.3005
R623 VTAIL.n81 VTAIL.n80 9.3005
R624 VTAIL.n83 VTAIL.n82 9.3005
R625 VTAIL.n8 VTAIL.n7 9.3005
R626 VTAIL.n89 VTAIL.n88 9.3005
R627 VTAIL.n91 VTAIL.n90 9.3005
R628 VTAIL.n4 VTAIL.n3 9.3005
R629 VTAIL.n97 VTAIL.n96 9.3005
R630 VTAIL.n99 VTAIL.n98 9.3005
R631 VTAIL.n75 VTAIL.n74 9.3005
R632 VTAIL.n73 VTAIL.n72 9.3005
R633 VTAIL.n16 VTAIL.n15 9.3005
R634 VTAIL.n67 VTAIL.n66 9.3005
R635 VTAIL.n65 VTAIL.n64 9.3005
R636 VTAIL.n20 VTAIL.n19 9.3005
R637 VTAIL.n59 VTAIL.n58 9.3005
R638 VTAIL.n32 VTAIL.n31 9.3005
R639 VTAIL.n39 VTAIL.n38 9.3005
R640 VTAIL.n41 VTAIL.n40 9.3005
R641 VTAIL.n28 VTAIL.n27 9.3005
R642 VTAIL.n47 VTAIL.n46 9.3005
R643 VTAIL.n49 VTAIL.n48 9.3005
R644 VTAIL.n50 VTAIL.n23 9.3005
R645 VTAIL.n57 VTAIL.n56 9.3005
R646 VTAIL.n12 VTAIL.n11 9.3005
R647 VTAIL.n185 VTAIL.n184 9.3005
R648 VTAIL.n187 VTAIL.n186 9.3005
R649 VTAIL.n112 VTAIL.n111 9.3005
R650 VTAIL.n193 VTAIL.n192 9.3005
R651 VTAIL.n195 VTAIL.n194 9.3005
R652 VTAIL.n108 VTAIL.n107 9.3005
R653 VTAIL.n201 VTAIL.n200 9.3005
R654 VTAIL.n203 VTAIL.n202 9.3005
R655 VTAIL.n179 VTAIL.n178 9.3005
R656 VTAIL.n177 VTAIL.n176 9.3005
R657 VTAIL.n120 VTAIL.n119 9.3005
R658 VTAIL.n171 VTAIL.n170 9.3005
R659 VTAIL.n169 VTAIL.n168 9.3005
R660 VTAIL.n124 VTAIL.n123 9.3005
R661 VTAIL.n163 VTAIL.n162 9.3005
R662 VTAIL.n136 VTAIL.n135 9.3005
R663 VTAIL.n143 VTAIL.n142 9.3005
R664 VTAIL.n145 VTAIL.n144 9.3005
R665 VTAIL.n132 VTAIL.n131 9.3005
R666 VTAIL.n151 VTAIL.n150 9.3005
R667 VTAIL.n153 VTAIL.n152 9.3005
R668 VTAIL.n154 VTAIL.n127 9.3005
R669 VTAIL.n161 VTAIL.n160 9.3005
R670 VTAIL.n116 VTAIL.n115 9.3005
R671 VTAIL.n289 VTAIL.n288 9.3005
R672 VTAIL.n291 VTAIL.n290 9.3005
R673 VTAIL.n216 VTAIL.n215 9.3005
R674 VTAIL.n297 VTAIL.n296 9.3005
R675 VTAIL.n299 VTAIL.n298 9.3005
R676 VTAIL.n212 VTAIL.n211 9.3005
R677 VTAIL.n305 VTAIL.n304 9.3005
R678 VTAIL.n307 VTAIL.n306 9.3005
R679 VTAIL.n283 VTAIL.n282 9.3005
R680 VTAIL.n281 VTAIL.n280 9.3005
R681 VTAIL.n224 VTAIL.n223 9.3005
R682 VTAIL.n275 VTAIL.n274 9.3005
R683 VTAIL.n273 VTAIL.n272 9.3005
R684 VTAIL.n228 VTAIL.n227 9.3005
R685 VTAIL.n267 VTAIL.n266 9.3005
R686 VTAIL.n240 VTAIL.n239 9.3005
R687 VTAIL.n247 VTAIL.n246 9.3005
R688 VTAIL.n249 VTAIL.n248 9.3005
R689 VTAIL.n236 VTAIL.n235 9.3005
R690 VTAIL.n255 VTAIL.n254 9.3005
R691 VTAIL.n257 VTAIL.n256 9.3005
R692 VTAIL.n258 VTAIL.n231 9.3005
R693 VTAIL.n265 VTAIL.n264 9.3005
R694 VTAIL.n220 VTAIL.n219 9.3005
R695 VTAIL.n723 VTAIL.n722 9.3005
R696 VTAIL.n721 VTAIL.n720 9.3005
R697 VTAIL.n628 VTAIL.n627 9.3005
R698 VTAIL.n715 VTAIL.n714 9.3005
R699 VTAIL.n713 VTAIL.n712 9.3005
R700 VTAIL.n632 VTAIL.n631 9.3005
R701 VTAIL.n707 VTAIL.n706 9.3005
R702 VTAIL.n705 VTAIL.n704 9.3005
R703 VTAIL.n636 VTAIL.n635 9.3005
R704 VTAIL.n699 VTAIL.n698 9.3005
R705 VTAIL.n697 VTAIL.n696 9.3005
R706 VTAIL.n640 VTAIL.n639 9.3005
R707 VTAIL.n691 VTAIL.n690 9.3005
R708 VTAIL.n689 VTAIL.n688 9.3005
R709 VTAIL.n644 VTAIL.n643 9.3005
R710 VTAIL.n683 VTAIL.n682 9.3005
R711 VTAIL.n681 VTAIL.n680 9.3005
R712 VTAIL.n649 VTAIL.n647 9.3005
R713 VTAIL.n675 VTAIL.n674 9.3005
R714 VTAIL.n673 VTAIL.n672 9.3005
R715 VTAIL.n654 VTAIL.n653 9.3005
R716 VTAIL.n667 VTAIL.n666 9.3005
R717 VTAIL.n665 VTAIL.n664 9.3005
R718 VTAIL.n658 VTAIL.n657 9.3005
R719 VTAIL.n554 VTAIL.n553 9.3005
R720 VTAIL.n561 VTAIL.n560 9.3005
R721 VTAIL.n563 VTAIL.n562 9.3005
R722 VTAIL.n550 VTAIL.n549 9.3005
R723 VTAIL.n569 VTAIL.n568 9.3005
R724 VTAIL.n571 VTAIL.n570 9.3005
R725 VTAIL.n545 VTAIL.n543 9.3005
R726 VTAIL.n577 VTAIL.n576 9.3005
R727 VTAIL.n603 VTAIL.n602 9.3005
R728 VTAIL.n528 VTAIL.n527 9.3005
R729 VTAIL.n609 VTAIL.n608 9.3005
R730 VTAIL.n611 VTAIL.n610 9.3005
R731 VTAIL.n524 VTAIL.n523 9.3005
R732 VTAIL.n617 VTAIL.n616 9.3005
R733 VTAIL.n619 VTAIL.n618 9.3005
R734 VTAIL.n601 VTAIL.n600 9.3005
R735 VTAIL.n532 VTAIL.n531 9.3005
R736 VTAIL.n595 VTAIL.n594 9.3005
R737 VTAIL.n593 VTAIL.n592 9.3005
R738 VTAIL.n536 VTAIL.n535 9.3005
R739 VTAIL.n587 VTAIL.n586 9.3005
R740 VTAIL.n585 VTAIL.n584 9.3005
R741 VTAIL.n540 VTAIL.n539 9.3005
R742 VTAIL.n579 VTAIL.n578 9.3005
R743 VTAIL.n450 VTAIL.n449 9.3005
R744 VTAIL.n457 VTAIL.n456 9.3005
R745 VTAIL.n459 VTAIL.n458 9.3005
R746 VTAIL.n446 VTAIL.n445 9.3005
R747 VTAIL.n465 VTAIL.n464 9.3005
R748 VTAIL.n467 VTAIL.n466 9.3005
R749 VTAIL.n441 VTAIL.n439 9.3005
R750 VTAIL.n473 VTAIL.n472 9.3005
R751 VTAIL.n499 VTAIL.n498 9.3005
R752 VTAIL.n424 VTAIL.n423 9.3005
R753 VTAIL.n505 VTAIL.n504 9.3005
R754 VTAIL.n507 VTAIL.n506 9.3005
R755 VTAIL.n420 VTAIL.n419 9.3005
R756 VTAIL.n513 VTAIL.n512 9.3005
R757 VTAIL.n515 VTAIL.n514 9.3005
R758 VTAIL.n497 VTAIL.n496 9.3005
R759 VTAIL.n428 VTAIL.n427 9.3005
R760 VTAIL.n491 VTAIL.n490 9.3005
R761 VTAIL.n489 VTAIL.n488 9.3005
R762 VTAIL.n432 VTAIL.n431 9.3005
R763 VTAIL.n483 VTAIL.n482 9.3005
R764 VTAIL.n481 VTAIL.n480 9.3005
R765 VTAIL.n436 VTAIL.n435 9.3005
R766 VTAIL.n475 VTAIL.n474 9.3005
R767 VTAIL.n346 VTAIL.n345 9.3005
R768 VTAIL.n353 VTAIL.n352 9.3005
R769 VTAIL.n355 VTAIL.n354 9.3005
R770 VTAIL.n342 VTAIL.n341 9.3005
R771 VTAIL.n361 VTAIL.n360 9.3005
R772 VTAIL.n363 VTAIL.n362 9.3005
R773 VTAIL.n337 VTAIL.n335 9.3005
R774 VTAIL.n369 VTAIL.n368 9.3005
R775 VTAIL.n395 VTAIL.n394 9.3005
R776 VTAIL.n320 VTAIL.n319 9.3005
R777 VTAIL.n401 VTAIL.n400 9.3005
R778 VTAIL.n403 VTAIL.n402 9.3005
R779 VTAIL.n316 VTAIL.n315 9.3005
R780 VTAIL.n409 VTAIL.n408 9.3005
R781 VTAIL.n411 VTAIL.n410 9.3005
R782 VTAIL.n393 VTAIL.n392 9.3005
R783 VTAIL.n324 VTAIL.n323 9.3005
R784 VTAIL.n387 VTAIL.n386 9.3005
R785 VTAIL.n385 VTAIL.n384 9.3005
R786 VTAIL.n328 VTAIL.n327 9.3005
R787 VTAIL.n379 VTAIL.n378 9.3005
R788 VTAIL.n377 VTAIL.n376 9.3005
R789 VTAIL.n332 VTAIL.n331 9.3005
R790 VTAIL.n371 VTAIL.n370 9.3005
R791 VTAIL.n769 VTAIL.n758 8.92171
R792 VTAIL.n800 VTAIL.n742 8.92171
R793 VTAIL.n816 VTAIL.n815 8.92171
R794 VTAIL.n41 VTAIL.n30 8.92171
R795 VTAIL.n72 VTAIL.n14 8.92171
R796 VTAIL.n88 VTAIL.n87 8.92171
R797 VTAIL.n145 VTAIL.n134 8.92171
R798 VTAIL.n176 VTAIL.n118 8.92171
R799 VTAIL.n192 VTAIL.n191 8.92171
R800 VTAIL.n249 VTAIL.n238 8.92171
R801 VTAIL.n280 VTAIL.n222 8.92171
R802 VTAIL.n296 VTAIL.n295 8.92171
R803 VTAIL.n712 VTAIL.n711 8.92171
R804 VTAIL.n696 VTAIL.n638 8.92171
R805 VTAIL.n667 VTAIL.n656 8.92171
R806 VTAIL.n608 VTAIL.n607 8.92171
R807 VTAIL.n592 VTAIL.n534 8.92171
R808 VTAIL.n563 VTAIL.n552 8.92171
R809 VTAIL.n504 VTAIL.n503 8.92171
R810 VTAIL.n488 VTAIL.n430 8.92171
R811 VTAIL.n459 VTAIL.n448 8.92171
R812 VTAIL.n400 VTAIL.n399 8.92171
R813 VTAIL.n384 VTAIL.n326 8.92171
R814 VTAIL.n355 VTAIL.n344 8.92171
R815 VTAIL.n766 VTAIL.n765 8.14595
R816 VTAIL.n804 VTAIL.n803 8.14595
R817 VTAIL.n812 VTAIL.n736 8.14595
R818 VTAIL.n38 VTAIL.n37 8.14595
R819 VTAIL.n76 VTAIL.n75 8.14595
R820 VTAIL.n84 VTAIL.n8 8.14595
R821 VTAIL.n142 VTAIL.n141 8.14595
R822 VTAIL.n180 VTAIL.n179 8.14595
R823 VTAIL.n188 VTAIL.n112 8.14595
R824 VTAIL.n246 VTAIL.n245 8.14595
R825 VTAIL.n284 VTAIL.n283 8.14595
R826 VTAIL.n292 VTAIL.n216 8.14595
R827 VTAIL.n708 VTAIL.n632 8.14595
R828 VTAIL.n700 VTAIL.n699 8.14595
R829 VTAIL.n664 VTAIL.n663 8.14595
R830 VTAIL.n604 VTAIL.n528 8.14595
R831 VTAIL.n596 VTAIL.n595 8.14595
R832 VTAIL.n560 VTAIL.n559 8.14595
R833 VTAIL.n500 VTAIL.n424 8.14595
R834 VTAIL.n492 VTAIL.n491 8.14595
R835 VTAIL.n456 VTAIL.n455 8.14595
R836 VTAIL.n396 VTAIL.n320 8.14595
R837 VTAIL.n388 VTAIL.n387 8.14595
R838 VTAIL.n352 VTAIL.n351 8.14595
R839 VTAIL.n762 VTAIL.n760 7.3702
R840 VTAIL.n807 VTAIL.n740 7.3702
R841 VTAIL.n811 VTAIL.n738 7.3702
R842 VTAIL.n34 VTAIL.n32 7.3702
R843 VTAIL.n79 VTAIL.n12 7.3702
R844 VTAIL.n83 VTAIL.n10 7.3702
R845 VTAIL.n138 VTAIL.n136 7.3702
R846 VTAIL.n183 VTAIL.n116 7.3702
R847 VTAIL.n187 VTAIL.n114 7.3702
R848 VTAIL.n242 VTAIL.n240 7.3702
R849 VTAIL.n287 VTAIL.n220 7.3702
R850 VTAIL.n291 VTAIL.n218 7.3702
R851 VTAIL.n707 VTAIL.n634 7.3702
R852 VTAIL.n703 VTAIL.n636 7.3702
R853 VTAIL.n660 VTAIL.n658 7.3702
R854 VTAIL.n603 VTAIL.n530 7.3702
R855 VTAIL.n599 VTAIL.n532 7.3702
R856 VTAIL.n556 VTAIL.n554 7.3702
R857 VTAIL.n499 VTAIL.n426 7.3702
R858 VTAIL.n495 VTAIL.n428 7.3702
R859 VTAIL.n452 VTAIL.n450 7.3702
R860 VTAIL.n395 VTAIL.n322 7.3702
R861 VTAIL.n391 VTAIL.n324 7.3702
R862 VTAIL.n348 VTAIL.n346 7.3702
R863 VTAIL.n808 VTAIL.n807 6.59444
R864 VTAIL.n808 VTAIL.n738 6.59444
R865 VTAIL.n80 VTAIL.n79 6.59444
R866 VTAIL.n80 VTAIL.n10 6.59444
R867 VTAIL.n184 VTAIL.n183 6.59444
R868 VTAIL.n184 VTAIL.n114 6.59444
R869 VTAIL.n288 VTAIL.n287 6.59444
R870 VTAIL.n288 VTAIL.n218 6.59444
R871 VTAIL.n704 VTAIL.n634 6.59444
R872 VTAIL.n704 VTAIL.n703 6.59444
R873 VTAIL.n600 VTAIL.n530 6.59444
R874 VTAIL.n600 VTAIL.n599 6.59444
R875 VTAIL.n496 VTAIL.n426 6.59444
R876 VTAIL.n496 VTAIL.n495 6.59444
R877 VTAIL.n392 VTAIL.n322 6.59444
R878 VTAIL.n392 VTAIL.n391 6.59444
R879 VTAIL.n765 VTAIL.n760 5.81868
R880 VTAIL.n804 VTAIL.n740 5.81868
R881 VTAIL.n812 VTAIL.n811 5.81868
R882 VTAIL.n37 VTAIL.n32 5.81868
R883 VTAIL.n76 VTAIL.n12 5.81868
R884 VTAIL.n84 VTAIL.n83 5.81868
R885 VTAIL.n141 VTAIL.n136 5.81868
R886 VTAIL.n180 VTAIL.n116 5.81868
R887 VTAIL.n188 VTAIL.n187 5.81868
R888 VTAIL.n245 VTAIL.n240 5.81868
R889 VTAIL.n284 VTAIL.n220 5.81868
R890 VTAIL.n292 VTAIL.n291 5.81868
R891 VTAIL.n708 VTAIL.n707 5.81868
R892 VTAIL.n700 VTAIL.n636 5.81868
R893 VTAIL.n663 VTAIL.n658 5.81868
R894 VTAIL.n604 VTAIL.n603 5.81868
R895 VTAIL.n596 VTAIL.n532 5.81868
R896 VTAIL.n559 VTAIL.n554 5.81868
R897 VTAIL.n500 VTAIL.n499 5.81868
R898 VTAIL.n492 VTAIL.n428 5.81868
R899 VTAIL.n455 VTAIL.n450 5.81868
R900 VTAIL.n396 VTAIL.n395 5.81868
R901 VTAIL.n388 VTAIL.n324 5.81868
R902 VTAIL.n351 VTAIL.n346 5.81868
R903 VTAIL.n766 VTAIL.n758 5.04292
R904 VTAIL.n803 VTAIL.n742 5.04292
R905 VTAIL.n815 VTAIL.n736 5.04292
R906 VTAIL.n38 VTAIL.n30 5.04292
R907 VTAIL.n75 VTAIL.n14 5.04292
R908 VTAIL.n87 VTAIL.n8 5.04292
R909 VTAIL.n142 VTAIL.n134 5.04292
R910 VTAIL.n179 VTAIL.n118 5.04292
R911 VTAIL.n191 VTAIL.n112 5.04292
R912 VTAIL.n246 VTAIL.n238 5.04292
R913 VTAIL.n283 VTAIL.n222 5.04292
R914 VTAIL.n295 VTAIL.n216 5.04292
R915 VTAIL.n711 VTAIL.n632 5.04292
R916 VTAIL.n699 VTAIL.n638 5.04292
R917 VTAIL.n664 VTAIL.n656 5.04292
R918 VTAIL.n607 VTAIL.n528 5.04292
R919 VTAIL.n595 VTAIL.n534 5.04292
R920 VTAIL.n560 VTAIL.n552 5.04292
R921 VTAIL.n503 VTAIL.n424 5.04292
R922 VTAIL.n491 VTAIL.n430 5.04292
R923 VTAIL.n456 VTAIL.n448 5.04292
R924 VTAIL.n399 VTAIL.n320 5.04292
R925 VTAIL.n387 VTAIL.n326 5.04292
R926 VTAIL.n352 VTAIL.n344 5.04292
R927 VTAIL.n770 VTAIL.n769 4.26717
R928 VTAIL.n800 VTAIL.n799 4.26717
R929 VTAIL.n816 VTAIL.n734 4.26717
R930 VTAIL.n42 VTAIL.n41 4.26717
R931 VTAIL.n72 VTAIL.n71 4.26717
R932 VTAIL.n88 VTAIL.n6 4.26717
R933 VTAIL.n146 VTAIL.n145 4.26717
R934 VTAIL.n176 VTAIL.n175 4.26717
R935 VTAIL.n192 VTAIL.n110 4.26717
R936 VTAIL.n250 VTAIL.n249 4.26717
R937 VTAIL.n280 VTAIL.n279 4.26717
R938 VTAIL.n296 VTAIL.n214 4.26717
R939 VTAIL.n712 VTAIL.n630 4.26717
R940 VTAIL.n696 VTAIL.n695 4.26717
R941 VTAIL.n668 VTAIL.n667 4.26717
R942 VTAIL.n608 VTAIL.n526 4.26717
R943 VTAIL.n592 VTAIL.n591 4.26717
R944 VTAIL.n564 VTAIL.n563 4.26717
R945 VTAIL.n504 VTAIL.n422 4.26717
R946 VTAIL.n488 VTAIL.n487 4.26717
R947 VTAIL.n460 VTAIL.n459 4.26717
R948 VTAIL.n400 VTAIL.n318 4.26717
R949 VTAIL.n384 VTAIL.n383 4.26717
R950 VTAIL.n356 VTAIL.n355 4.26717
R951 VTAIL.n773 VTAIL.n756 3.49141
R952 VTAIL.n796 VTAIL.n744 3.49141
R953 VTAIL.n820 VTAIL.n819 3.49141
R954 VTAIL.n45 VTAIL.n28 3.49141
R955 VTAIL.n68 VTAIL.n16 3.49141
R956 VTAIL.n92 VTAIL.n91 3.49141
R957 VTAIL.n149 VTAIL.n132 3.49141
R958 VTAIL.n172 VTAIL.n120 3.49141
R959 VTAIL.n196 VTAIL.n195 3.49141
R960 VTAIL.n253 VTAIL.n236 3.49141
R961 VTAIL.n276 VTAIL.n224 3.49141
R962 VTAIL.n300 VTAIL.n299 3.49141
R963 VTAIL.n716 VTAIL.n715 3.49141
R964 VTAIL.n692 VTAIL.n640 3.49141
R965 VTAIL.n671 VTAIL.n654 3.49141
R966 VTAIL.n612 VTAIL.n611 3.49141
R967 VTAIL.n588 VTAIL.n536 3.49141
R968 VTAIL.n567 VTAIL.n550 3.49141
R969 VTAIL.n508 VTAIL.n507 3.49141
R970 VTAIL.n484 VTAIL.n432 3.49141
R971 VTAIL.n463 VTAIL.n446 3.49141
R972 VTAIL.n404 VTAIL.n403 3.49141
R973 VTAIL.n380 VTAIL.n328 3.49141
R974 VTAIL.n359 VTAIL.n342 3.49141
R975 VTAIL.n761 VTAIL.n759 2.84303
R976 VTAIL.n33 VTAIL.n31 2.84303
R977 VTAIL.n137 VTAIL.n135 2.84303
R978 VTAIL.n241 VTAIL.n239 2.84303
R979 VTAIL.n659 VTAIL.n657 2.84303
R980 VTAIL.n555 VTAIL.n553 2.84303
R981 VTAIL.n451 VTAIL.n449 2.84303
R982 VTAIL.n347 VTAIL.n345 2.84303
R983 VTAIL.n774 VTAIL.n754 2.71565
R984 VTAIL.n795 VTAIL.n746 2.71565
R985 VTAIL.n823 VTAIL.n732 2.71565
R986 VTAIL.n46 VTAIL.n26 2.71565
R987 VTAIL.n67 VTAIL.n18 2.71565
R988 VTAIL.n95 VTAIL.n4 2.71565
R989 VTAIL.n150 VTAIL.n130 2.71565
R990 VTAIL.n171 VTAIL.n122 2.71565
R991 VTAIL.n199 VTAIL.n108 2.71565
R992 VTAIL.n254 VTAIL.n234 2.71565
R993 VTAIL.n275 VTAIL.n226 2.71565
R994 VTAIL.n303 VTAIL.n212 2.71565
R995 VTAIL.n719 VTAIL.n628 2.71565
R996 VTAIL.n691 VTAIL.n642 2.71565
R997 VTAIL.n672 VTAIL.n652 2.71565
R998 VTAIL.n615 VTAIL.n524 2.71565
R999 VTAIL.n587 VTAIL.n538 2.71565
R1000 VTAIL.n568 VTAIL.n548 2.71565
R1001 VTAIL.n511 VTAIL.n420 2.71565
R1002 VTAIL.n483 VTAIL.n434 2.71565
R1003 VTAIL.n464 VTAIL.n444 2.71565
R1004 VTAIL.n407 VTAIL.n316 2.71565
R1005 VTAIL.n379 VTAIL.n330 2.71565
R1006 VTAIL.n360 VTAIL.n340 2.71565
R1007 VTAIL.n779 VTAIL.n777 1.93989
R1008 VTAIL.n792 VTAIL.n791 1.93989
R1009 VTAIL.n824 VTAIL.n730 1.93989
R1010 VTAIL.n51 VTAIL.n49 1.93989
R1011 VTAIL.n64 VTAIL.n63 1.93989
R1012 VTAIL.n96 VTAIL.n2 1.93989
R1013 VTAIL.n155 VTAIL.n153 1.93989
R1014 VTAIL.n168 VTAIL.n167 1.93989
R1015 VTAIL.n200 VTAIL.n106 1.93989
R1016 VTAIL.n259 VTAIL.n257 1.93989
R1017 VTAIL.n272 VTAIL.n271 1.93989
R1018 VTAIL.n304 VTAIL.n210 1.93989
R1019 VTAIL.n720 VTAIL.n626 1.93989
R1020 VTAIL.n688 VTAIL.n687 1.93989
R1021 VTAIL.n676 VTAIL.n675 1.93989
R1022 VTAIL.n616 VTAIL.n522 1.93989
R1023 VTAIL.n584 VTAIL.n583 1.93989
R1024 VTAIL.n572 VTAIL.n571 1.93989
R1025 VTAIL.n512 VTAIL.n418 1.93989
R1026 VTAIL.n480 VTAIL.n479 1.93989
R1027 VTAIL.n468 VTAIL.n467 1.93989
R1028 VTAIL.n408 VTAIL.n314 1.93989
R1029 VTAIL.n376 VTAIL.n375 1.93989
R1030 VTAIL.n364 VTAIL.n363 1.93989
R1031 VTAIL.n778 VTAIL.n752 1.16414
R1032 VTAIL.n788 VTAIL.n748 1.16414
R1033 VTAIL.n828 VTAIL.n827 1.16414
R1034 VTAIL.n50 VTAIL.n24 1.16414
R1035 VTAIL.n60 VTAIL.n20 1.16414
R1036 VTAIL.n100 VTAIL.n99 1.16414
R1037 VTAIL.n154 VTAIL.n128 1.16414
R1038 VTAIL.n164 VTAIL.n124 1.16414
R1039 VTAIL.n204 VTAIL.n203 1.16414
R1040 VTAIL.n258 VTAIL.n232 1.16414
R1041 VTAIL.n268 VTAIL.n228 1.16414
R1042 VTAIL.n308 VTAIL.n307 1.16414
R1043 VTAIL.n724 VTAIL.n723 1.16414
R1044 VTAIL.n684 VTAIL.n644 1.16414
R1045 VTAIL.n679 VTAIL.n649 1.16414
R1046 VTAIL.n620 VTAIL.n619 1.16414
R1047 VTAIL.n580 VTAIL.n540 1.16414
R1048 VTAIL.n575 VTAIL.n545 1.16414
R1049 VTAIL.n516 VTAIL.n515 1.16414
R1050 VTAIL.n476 VTAIL.n436 1.16414
R1051 VTAIL.n471 VTAIL.n441 1.16414
R1052 VTAIL.n412 VTAIL.n411 1.16414
R1053 VTAIL.n372 VTAIL.n332 1.16414
R1054 VTAIL.n367 VTAIL.n337 1.16414
R1055 VTAIL.n519 VTAIL.n415 0.87119
R1056 VTAIL.n727 VTAIL.n623 0.87119
R1057 VTAIL.n311 VTAIL.n207 0.87119
R1058 VTAIL VTAIL.n103 0.494034
R1059 VTAIL.n623 VTAIL.n519 0.470328
R1060 VTAIL.n207 VTAIL.n103 0.470328
R1061 VTAIL.n784 VTAIL.n783 0.388379
R1062 VTAIL.n787 VTAIL.n750 0.388379
R1063 VTAIL.n830 VTAIL.n728 0.388379
R1064 VTAIL.n56 VTAIL.n55 0.388379
R1065 VTAIL.n59 VTAIL.n22 0.388379
R1066 VTAIL.n102 VTAIL.n0 0.388379
R1067 VTAIL.n160 VTAIL.n159 0.388379
R1068 VTAIL.n163 VTAIL.n126 0.388379
R1069 VTAIL.n206 VTAIL.n104 0.388379
R1070 VTAIL.n264 VTAIL.n263 0.388379
R1071 VTAIL.n267 VTAIL.n230 0.388379
R1072 VTAIL.n310 VTAIL.n208 0.388379
R1073 VTAIL.n726 VTAIL.n624 0.388379
R1074 VTAIL.n683 VTAIL.n646 0.388379
R1075 VTAIL.n680 VTAIL.n648 0.388379
R1076 VTAIL.n622 VTAIL.n520 0.388379
R1077 VTAIL.n579 VTAIL.n542 0.388379
R1078 VTAIL.n576 VTAIL.n544 0.388379
R1079 VTAIL.n518 VTAIL.n416 0.388379
R1080 VTAIL.n475 VTAIL.n438 0.388379
R1081 VTAIL.n472 VTAIL.n440 0.388379
R1082 VTAIL.n414 VTAIL.n312 0.388379
R1083 VTAIL.n371 VTAIL.n334 0.388379
R1084 VTAIL.n368 VTAIL.n336 0.388379
R1085 VTAIL VTAIL.n831 0.377655
R1086 VTAIL.n767 VTAIL.n759 0.155672
R1087 VTAIL.n768 VTAIL.n767 0.155672
R1088 VTAIL.n768 VTAIL.n755 0.155672
R1089 VTAIL.n775 VTAIL.n755 0.155672
R1090 VTAIL.n776 VTAIL.n775 0.155672
R1091 VTAIL.n776 VTAIL.n751 0.155672
R1092 VTAIL.n785 VTAIL.n751 0.155672
R1093 VTAIL.n786 VTAIL.n785 0.155672
R1094 VTAIL.n786 VTAIL.n747 0.155672
R1095 VTAIL.n793 VTAIL.n747 0.155672
R1096 VTAIL.n794 VTAIL.n793 0.155672
R1097 VTAIL.n794 VTAIL.n743 0.155672
R1098 VTAIL.n801 VTAIL.n743 0.155672
R1099 VTAIL.n802 VTAIL.n801 0.155672
R1100 VTAIL.n802 VTAIL.n739 0.155672
R1101 VTAIL.n809 VTAIL.n739 0.155672
R1102 VTAIL.n810 VTAIL.n809 0.155672
R1103 VTAIL.n810 VTAIL.n735 0.155672
R1104 VTAIL.n817 VTAIL.n735 0.155672
R1105 VTAIL.n818 VTAIL.n817 0.155672
R1106 VTAIL.n818 VTAIL.n731 0.155672
R1107 VTAIL.n825 VTAIL.n731 0.155672
R1108 VTAIL.n826 VTAIL.n825 0.155672
R1109 VTAIL.n39 VTAIL.n31 0.155672
R1110 VTAIL.n40 VTAIL.n39 0.155672
R1111 VTAIL.n40 VTAIL.n27 0.155672
R1112 VTAIL.n47 VTAIL.n27 0.155672
R1113 VTAIL.n48 VTAIL.n47 0.155672
R1114 VTAIL.n48 VTAIL.n23 0.155672
R1115 VTAIL.n57 VTAIL.n23 0.155672
R1116 VTAIL.n58 VTAIL.n57 0.155672
R1117 VTAIL.n58 VTAIL.n19 0.155672
R1118 VTAIL.n65 VTAIL.n19 0.155672
R1119 VTAIL.n66 VTAIL.n65 0.155672
R1120 VTAIL.n66 VTAIL.n15 0.155672
R1121 VTAIL.n73 VTAIL.n15 0.155672
R1122 VTAIL.n74 VTAIL.n73 0.155672
R1123 VTAIL.n74 VTAIL.n11 0.155672
R1124 VTAIL.n81 VTAIL.n11 0.155672
R1125 VTAIL.n82 VTAIL.n81 0.155672
R1126 VTAIL.n82 VTAIL.n7 0.155672
R1127 VTAIL.n89 VTAIL.n7 0.155672
R1128 VTAIL.n90 VTAIL.n89 0.155672
R1129 VTAIL.n90 VTAIL.n3 0.155672
R1130 VTAIL.n97 VTAIL.n3 0.155672
R1131 VTAIL.n98 VTAIL.n97 0.155672
R1132 VTAIL.n143 VTAIL.n135 0.155672
R1133 VTAIL.n144 VTAIL.n143 0.155672
R1134 VTAIL.n144 VTAIL.n131 0.155672
R1135 VTAIL.n151 VTAIL.n131 0.155672
R1136 VTAIL.n152 VTAIL.n151 0.155672
R1137 VTAIL.n152 VTAIL.n127 0.155672
R1138 VTAIL.n161 VTAIL.n127 0.155672
R1139 VTAIL.n162 VTAIL.n161 0.155672
R1140 VTAIL.n162 VTAIL.n123 0.155672
R1141 VTAIL.n169 VTAIL.n123 0.155672
R1142 VTAIL.n170 VTAIL.n169 0.155672
R1143 VTAIL.n170 VTAIL.n119 0.155672
R1144 VTAIL.n177 VTAIL.n119 0.155672
R1145 VTAIL.n178 VTAIL.n177 0.155672
R1146 VTAIL.n178 VTAIL.n115 0.155672
R1147 VTAIL.n185 VTAIL.n115 0.155672
R1148 VTAIL.n186 VTAIL.n185 0.155672
R1149 VTAIL.n186 VTAIL.n111 0.155672
R1150 VTAIL.n193 VTAIL.n111 0.155672
R1151 VTAIL.n194 VTAIL.n193 0.155672
R1152 VTAIL.n194 VTAIL.n107 0.155672
R1153 VTAIL.n201 VTAIL.n107 0.155672
R1154 VTAIL.n202 VTAIL.n201 0.155672
R1155 VTAIL.n247 VTAIL.n239 0.155672
R1156 VTAIL.n248 VTAIL.n247 0.155672
R1157 VTAIL.n248 VTAIL.n235 0.155672
R1158 VTAIL.n255 VTAIL.n235 0.155672
R1159 VTAIL.n256 VTAIL.n255 0.155672
R1160 VTAIL.n256 VTAIL.n231 0.155672
R1161 VTAIL.n265 VTAIL.n231 0.155672
R1162 VTAIL.n266 VTAIL.n265 0.155672
R1163 VTAIL.n266 VTAIL.n227 0.155672
R1164 VTAIL.n273 VTAIL.n227 0.155672
R1165 VTAIL.n274 VTAIL.n273 0.155672
R1166 VTAIL.n274 VTAIL.n223 0.155672
R1167 VTAIL.n281 VTAIL.n223 0.155672
R1168 VTAIL.n282 VTAIL.n281 0.155672
R1169 VTAIL.n282 VTAIL.n219 0.155672
R1170 VTAIL.n289 VTAIL.n219 0.155672
R1171 VTAIL.n290 VTAIL.n289 0.155672
R1172 VTAIL.n290 VTAIL.n215 0.155672
R1173 VTAIL.n297 VTAIL.n215 0.155672
R1174 VTAIL.n298 VTAIL.n297 0.155672
R1175 VTAIL.n298 VTAIL.n211 0.155672
R1176 VTAIL.n305 VTAIL.n211 0.155672
R1177 VTAIL.n306 VTAIL.n305 0.155672
R1178 VTAIL.n722 VTAIL.n721 0.155672
R1179 VTAIL.n721 VTAIL.n627 0.155672
R1180 VTAIL.n714 VTAIL.n627 0.155672
R1181 VTAIL.n714 VTAIL.n713 0.155672
R1182 VTAIL.n713 VTAIL.n631 0.155672
R1183 VTAIL.n706 VTAIL.n631 0.155672
R1184 VTAIL.n706 VTAIL.n705 0.155672
R1185 VTAIL.n705 VTAIL.n635 0.155672
R1186 VTAIL.n698 VTAIL.n635 0.155672
R1187 VTAIL.n698 VTAIL.n697 0.155672
R1188 VTAIL.n697 VTAIL.n639 0.155672
R1189 VTAIL.n690 VTAIL.n639 0.155672
R1190 VTAIL.n690 VTAIL.n689 0.155672
R1191 VTAIL.n689 VTAIL.n643 0.155672
R1192 VTAIL.n682 VTAIL.n643 0.155672
R1193 VTAIL.n682 VTAIL.n681 0.155672
R1194 VTAIL.n681 VTAIL.n647 0.155672
R1195 VTAIL.n674 VTAIL.n647 0.155672
R1196 VTAIL.n674 VTAIL.n673 0.155672
R1197 VTAIL.n673 VTAIL.n653 0.155672
R1198 VTAIL.n666 VTAIL.n653 0.155672
R1199 VTAIL.n666 VTAIL.n665 0.155672
R1200 VTAIL.n665 VTAIL.n657 0.155672
R1201 VTAIL.n618 VTAIL.n617 0.155672
R1202 VTAIL.n617 VTAIL.n523 0.155672
R1203 VTAIL.n610 VTAIL.n523 0.155672
R1204 VTAIL.n610 VTAIL.n609 0.155672
R1205 VTAIL.n609 VTAIL.n527 0.155672
R1206 VTAIL.n602 VTAIL.n527 0.155672
R1207 VTAIL.n602 VTAIL.n601 0.155672
R1208 VTAIL.n601 VTAIL.n531 0.155672
R1209 VTAIL.n594 VTAIL.n531 0.155672
R1210 VTAIL.n594 VTAIL.n593 0.155672
R1211 VTAIL.n593 VTAIL.n535 0.155672
R1212 VTAIL.n586 VTAIL.n535 0.155672
R1213 VTAIL.n586 VTAIL.n585 0.155672
R1214 VTAIL.n585 VTAIL.n539 0.155672
R1215 VTAIL.n578 VTAIL.n539 0.155672
R1216 VTAIL.n578 VTAIL.n577 0.155672
R1217 VTAIL.n577 VTAIL.n543 0.155672
R1218 VTAIL.n570 VTAIL.n543 0.155672
R1219 VTAIL.n570 VTAIL.n569 0.155672
R1220 VTAIL.n569 VTAIL.n549 0.155672
R1221 VTAIL.n562 VTAIL.n549 0.155672
R1222 VTAIL.n562 VTAIL.n561 0.155672
R1223 VTAIL.n561 VTAIL.n553 0.155672
R1224 VTAIL.n514 VTAIL.n513 0.155672
R1225 VTAIL.n513 VTAIL.n419 0.155672
R1226 VTAIL.n506 VTAIL.n419 0.155672
R1227 VTAIL.n506 VTAIL.n505 0.155672
R1228 VTAIL.n505 VTAIL.n423 0.155672
R1229 VTAIL.n498 VTAIL.n423 0.155672
R1230 VTAIL.n498 VTAIL.n497 0.155672
R1231 VTAIL.n497 VTAIL.n427 0.155672
R1232 VTAIL.n490 VTAIL.n427 0.155672
R1233 VTAIL.n490 VTAIL.n489 0.155672
R1234 VTAIL.n489 VTAIL.n431 0.155672
R1235 VTAIL.n482 VTAIL.n431 0.155672
R1236 VTAIL.n482 VTAIL.n481 0.155672
R1237 VTAIL.n481 VTAIL.n435 0.155672
R1238 VTAIL.n474 VTAIL.n435 0.155672
R1239 VTAIL.n474 VTAIL.n473 0.155672
R1240 VTAIL.n473 VTAIL.n439 0.155672
R1241 VTAIL.n466 VTAIL.n439 0.155672
R1242 VTAIL.n466 VTAIL.n465 0.155672
R1243 VTAIL.n465 VTAIL.n445 0.155672
R1244 VTAIL.n458 VTAIL.n445 0.155672
R1245 VTAIL.n458 VTAIL.n457 0.155672
R1246 VTAIL.n457 VTAIL.n449 0.155672
R1247 VTAIL.n410 VTAIL.n409 0.155672
R1248 VTAIL.n409 VTAIL.n315 0.155672
R1249 VTAIL.n402 VTAIL.n315 0.155672
R1250 VTAIL.n402 VTAIL.n401 0.155672
R1251 VTAIL.n401 VTAIL.n319 0.155672
R1252 VTAIL.n394 VTAIL.n319 0.155672
R1253 VTAIL.n394 VTAIL.n393 0.155672
R1254 VTAIL.n393 VTAIL.n323 0.155672
R1255 VTAIL.n386 VTAIL.n323 0.155672
R1256 VTAIL.n386 VTAIL.n385 0.155672
R1257 VTAIL.n385 VTAIL.n327 0.155672
R1258 VTAIL.n378 VTAIL.n327 0.155672
R1259 VTAIL.n378 VTAIL.n377 0.155672
R1260 VTAIL.n377 VTAIL.n331 0.155672
R1261 VTAIL.n370 VTAIL.n331 0.155672
R1262 VTAIL.n370 VTAIL.n369 0.155672
R1263 VTAIL.n369 VTAIL.n335 0.155672
R1264 VTAIL.n362 VTAIL.n335 0.155672
R1265 VTAIL.n362 VTAIL.n361 0.155672
R1266 VTAIL.n361 VTAIL.n341 0.155672
R1267 VTAIL.n354 VTAIL.n341 0.155672
R1268 VTAIL.n354 VTAIL.n353 0.155672
R1269 VTAIL.n353 VTAIL.n345 0.155672
R1270 B.n472 B.t4 868.803
R1271 B.n470 B.t8 868.803
R1272 B.n104 B.t11 868.803
R1273 B.n102 B.t15 868.803
R1274 B.n815 B.n814 585
R1275 B.n816 B.n815 585
R1276 B.n370 B.n101 585
R1277 B.n369 B.n368 585
R1278 B.n367 B.n366 585
R1279 B.n365 B.n364 585
R1280 B.n363 B.n362 585
R1281 B.n361 B.n360 585
R1282 B.n359 B.n358 585
R1283 B.n357 B.n356 585
R1284 B.n355 B.n354 585
R1285 B.n353 B.n352 585
R1286 B.n351 B.n350 585
R1287 B.n349 B.n348 585
R1288 B.n347 B.n346 585
R1289 B.n345 B.n344 585
R1290 B.n343 B.n342 585
R1291 B.n341 B.n340 585
R1292 B.n339 B.n338 585
R1293 B.n337 B.n336 585
R1294 B.n335 B.n334 585
R1295 B.n333 B.n332 585
R1296 B.n331 B.n330 585
R1297 B.n329 B.n328 585
R1298 B.n327 B.n326 585
R1299 B.n325 B.n324 585
R1300 B.n323 B.n322 585
R1301 B.n321 B.n320 585
R1302 B.n319 B.n318 585
R1303 B.n317 B.n316 585
R1304 B.n315 B.n314 585
R1305 B.n313 B.n312 585
R1306 B.n311 B.n310 585
R1307 B.n309 B.n308 585
R1308 B.n307 B.n306 585
R1309 B.n305 B.n304 585
R1310 B.n303 B.n302 585
R1311 B.n301 B.n300 585
R1312 B.n299 B.n298 585
R1313 B.n297 B.n296 585
R1314 B.n295 B.n294 585
R1315 B.n293 B.n292 585
R1316 B.n291 B.n290 585
R1317 B.n289 B.n288 585
R1318 B.n287 B.n286 585
R1319 B.n285 B.n284 585
R1320 B.n283 B.n282 585
R1321 B.n281 B.n280 585
R1322 B.n279 B.n278 585
R1323 B.n277 B.n276 585
R1324 B.n275 B.n274 585
R1325 B.n273 B.n272 585
R1326 B.n271 B.n270 585
R1327 B.n269 B.n268 585
R1328 B.n267 B.n266 585
R1329 B.n265 B.n264 585
R1330 B.n263 B.n262 585
R1331 B.n261 B.n260 585
R1332 B.n259 B.n258 585
R1333 B.n257 B.n256 585
R1334 B.n255 B.n254 585
R1335 B.n253 B.n252 585
R1336 B.n251 B.n250 585
R1337 B.n248 B.n247 585
R1338 B.n246 B.n245 585
R1339 B.n244 B.n243 585
R1340 B.n242 B.n241 585
R1341 B.n240 B.n239 585
R1342 B.n238 B.n237 585
R1343 B.n236 B.n235 585
R1344 B.n234 B.n233 585
R1345 B.n232 B.n231 585
R1346 B.n230 B.n229 585
R1347 B.n228 B.n227 585
R1348 B.n226 B.n225 585
R1349 B.n224 B.n223 585
R1350 B.n222 B.n221 585
R1351 B.n220 B.n219 585
R1352 B.n218 B.n217 585
R1353 B.n216 B.n215 585
R1354 B.n214 B.n213 585
R1355 B.n212 B.n211 585
R1356 B.n210 B.n209 585
R1357 B.n208 B.n207 585
R1358 B.n206 B.n205 585
R1359 B.n204 B.n203 585
R1360 B.n202 B.n201 585
R1361 B.n200 B.n199 585
R1362 B.n198 B.n197 585
R1363 B.n196 B.n195 585
R1364 B.n194 B.n193 585
R1365 B.n192 B.n191 585
R1366 B.n190 B.n189 585
R1367 B.n188 B.n187 585
R1368 B.n186 B.n185 585
R1369 B.n184 B.n183 585
R1370 B.n182 B.n181 585
R1371 B.n180 B.n179 585
R1372 B.n178 B.n177 585
R1373 B.n176 B.n175 585
R1374 B.n174 B.n173 585
R1375 B.n172 B.n171 585
R1376 B.n170 B.n169 585
R1377 B.n168 B.n167 585
R1378 B.n166 B.n165 585
R1379 B.n164 B.n163 585
R1380 B.n162 B.n161 585
R1381 B.n160 B.n159 585
R1382 B.n158 B.n157 585
R1383 B.n156 B.n155 585
R1384 B.n154 B.n153 585
R1385 B.n152 B.n151 585
R1386 B.n150 B.n149 585
R1387 B.n148 B.n147 585
R1388 B.n146 B.n145 585
R1389 B.n144 B.n143 585
R1390 B.n142 B.n141 585
R1391 B.n140 B.n139 585
R1392 B.n138 B.n137 585
R1393 B.n136 B.n135 585
R1394 B.n134 B.n133 585
R1395 B.n132 B.n131 585
R1396 B.n130 B.n129 585
R1397 B.n128 B.n127 585
R1398 B.n126 B.n125 585
R1399 B.n124 B.n123 585
R1400 B.n122 B.n121 585
R1401 B.n120 B.n119 585
R1402 B.n118 B.n117 585
R1403 B.n116 B.n115 585
R1404 B.n114 B.n113 585
R1405 B.n112 B.n111 585
R1406 B.n110 B.n109 585
R1407 B.n108 B.n107 585
R1408 B.n813 B.n34 585
R1409 B.n817 B.n34 585
R1410 B.n812 B.n33 585
R1411 B.n818 B.n33 585
R1412 B.n811 B.n810 585
R1413 B.n810 B.n29 585
R1414 B.n809 B.n28 585
R1415 B.n824 B.n28 585
R1416 B.n808 B.n27 585
R1417 B.n825 B.n27 585
R1418 B.n807 B.n26 585
R1419 B.n826 B.n26 585
R1420 B.n806 B.n805 585
R1421 B.n805 B.n22 585
R1422 B.n804 B.n21 585
R1423 B.n832 B.n21 585
R1424 B.n803 B.n20 585
R1425 B.n833 B.n20 585
R1426 B.n802 B.n19 585
R1427 B.n834 B.n19 585
R1428 B.n801 B.n800 585
R1429 B.n800 B.n18 585
R1430 B.n799 B.n14 585
R1431 B.n840 B.n14 585
R1432 B.n798 B.n13 585
R1433 B.n841 B.n13 585
R1434 B.n797 B.n12 585
R1435 B.n842 B.n12 585
R1436 B.n796 B.n795 585
R1437 B.n795 B.n8 585
R1438 B.n794 B.n7 585
R1439 B.n848 B.n7 585
R1440 B.n793 B.n6 585
R1441 B.n849 B.n6 585
R1442 B.n792 B.n5 585
R1443 B.n850 B.n5 585
R1444 B.n791 B.n790 585
R1445 B.n790 B.n4 585
R1446 B.n789 B.n371 585
R1447 B.n789 B.n788 585
R1448 B.n779 B.n372 585
R1449 B.n373 B.n372 585
R1450 B.n781 B.n780 585
R1451 B.n782 B.n781 585
R1452 B.n778 B.n378 585
R1453 B.n378 B.n377 585
R1454 B.n777 B.n776 585
R1455 B.n776 B.n775 585
R1456 B.n380 B.n379 585
R1457 B.n768 B.n380 585
R1458 B.n767 B.n766 585
R1459 B.n769 B.n767 585
R1460 B.n765 B.n385 585
R1461 B.n385 B.n384 585
R1462 B.n764 B.n763 585
R1463 B.n763 B.n762 585
R1464 B.n387 B.n386 585
R1465 B.n388 B.n387 585
R1466 B.n755 B.n754 585
R1467 B.n756 B.n755 585
R1468 B.n753 B.n392 585
R1469 B.n396 B.n392 585
R1470 B.n752 B.n751 585
R1471 B.n751 B.n750 585
R1472 B.n394 B.n393 585
R1473 B.n395 B.n394 585
R1474 B.n743 B.n742 585
R1475 B.n744 B.n743 585
R1476 B.n741 B.n401 585
R1477 B.n401 B.n400 585
R1478 B.n735 B.n734 585
R1479 B.n733 B.n469 585
R1480 B.n732 B.n468 585
R1481 B.n737 B.n468 585
R1482 B.n731 B.n730 585
R1483 B.n729 B.n728 585
R1484 B.n727 B.n726 585
R1485 B.n725 B.n724 585
R1486 B.n723 B.n722 585
R1487 B.n721 B.n720 585
R1488 B.n719 B.n718 585
R1489 B.n717 B.n716 585
R1490 B.n715 B.n714 585
R1491 B.n713 B.n712 585
R1492 B.n711 B.n710 585
R1493 B.n709 B.n708 585
R1494 B.n707 B.n706 585
R1495 B.n705 B.n704 585
R1496 B.n703 B.n702 585
R1497 B.n701 B.n700 585
R1498 B.n699 B.n698 585
R1499 B.n697 B.n696 585
R1500 B.n695 B.n694 585
R1501 B.n693 B.n692 585
R1502 B.n691 B.n690 585
R1503 B.n689 B.n688 585
R1504 B.n687 B.n686 585
R1505 B.n685 B.n684 585
R1506 B.n683 B.n682 585
R1507 B.n681 B.n680 585
R1508 B.n679 B.n678 585
R1509 B.n677 B.n676 585
R1510 B.n675 B.n674 585
R1511 B.n673 B.n672 585
R1512 B.n671 B.n670 585
R1513 B.n669 B.n668 585
R1514 B.n667 B.n666 585
R1515 B.n665 B.n664 585
R1516 B.n663 B.n662 585
R1517 B.n661 B.n660 585
R1518 B.n659 B.n658 585
R1519 B.n657 B.n656 585
R1520 B.n655 B.n654 585
R1521 B.n653 B.n652 585
R1522 B.n651 B.n650 585
R1523 B.n649 B.n648 585
R1524 B.n647 B.n646 585
R1525 B.n645 B.n644 585
R1526 B.n643 B.n642 585
R1527 B.n641 B.n640 585
R1528 B.n639 B.n638 585
R1529 B.n637 B.n636 585
R1530 B.n635 B.n634 585
R1531 B.n633 B.n632 585
R1532 B.n631 B.n630 585
R1533 B.n629 B.n628 585
R1534 B.n627 B.n626 585
R1535 B.n625 B.n624 585
R1536 B.n623 B.n622 585
R1537 B.n621 B.n620 585
R1538 B.n619 B.n618 585
R1539 B.n617 B.n616 585
R1540 B.n615 B.n614 585
R1541 B.n612 B.n611 585
R1542 B.n610 B.n609 585
R1543 B.n608 B.n607 585
R1544 B.n606 B.n605 585
R1545 B.n604 B.n603 585
R1546 B.n602 B.n601 585
R1547 B.n600 B.n599 585
R1548 B.n598 B.n597 585
R1549 B.n596 B.n595 585
R1550 B.n594 B.n593 585
R1551 B.n592 B.n591 585
R1552 B.n590 B.n589 585
R1553 B.n588 B.n587 585
R1554 B.n586 B.n585 585
R1555 B.n584 B.n583 585
R1556 B.n582 B.n581 585
R1557 B.n580 B.n579 585
R1558 B.n578 B.n577 585
R1559 B.n576 B.n575 585
R1560 B.n574 B.n573 585
R1561 B.n572 B.n571 585
R1562 B.n570 B.n569 585
R1563 B.n568 B.n567 585
R1564 B.n566 B.n565 585
R1565 B.n564 B.n563 585
R1566 B.n562 B.n561 585
R1567 B.n560 B.n559 585
R1568 B.n558 B.n557 585
R1569 B.n556 B.n555 585
R1570 B.n554 B.n553 585
R1571 B.n552 B.n551 585
R1572 B.n550 B.n549 585
R1573 B.n548 B.n547 585
R1574 B.n546 B.n545 585
R1575 B.n544 B.n543 585
R1576 B.n542 B.n541 585
R1577 B.n540 B.n539 585
R1578 B.n538 B.n537 585
R1579 B.n536 B.n535 585
R1580 B.n534 B.n533 585
R1581 B.n532 B.n531 585
R1582 B.n530 B.n529 585
R1583 B.n528 B.n527 585
R1584 B.n526 B.n525 585
R1585 B.n524 B.n523 585
R1586 B.n522 B.n521 585
R1587 B.n520 B.n519 585
R1588 B.n518 B.n517 585
R1589 B.n516 B.n515 585
R1590 B.n514 B.n513 585
R1591 B.n512 B.n511 585
R1592 B.n510 B.n509 585
R1593 B.n508 B.n507 585
R1594 B.n506 B.n505 585
R1595 B.n504 B.n503 585
R1596 B.n502 B.n501 585
R1597 B.n500 B.n499 585
R1598 B.n498 B.n497 585
R1599 B.n496 B.n495 585
R1600 B.n494 B.n493 585
R1601 B.n492 B.n491 585
R1602 B.n490 B.n489 585
R1603 B.n488 B.n487 585
R1604 B.n486 B.n485 585
R1605 B.n484 B.n483 585
R1606 B.n482 B.n481 585
R1607 B.n480 B.n479 585
R1608 B.n478 B.n477 585
R1609 B.n476 B.n475 585
R1610 B.n403 B.n402 585
R1611 B.n740 B.n739 585
R1612 B.n399 B.n398 585
R1613 B.n400 B.n399 585
R1614 B.n746 B.n745 585
R1615 B.n745 B.n744 585
R1616 B.n747 B.n397 585
R1617 B.n397 B.n395 585
R1618 B.n749 B.n748 585
R1619 B.n750 B.n749 585
R1620 B.n391 B.n390 585
R1621 B.n396 B.n391 585
R1622 B.n758 B.n757 585
R1623 B.n757 B.n756 585
R1624 B.n759 B.n389 585
R1625 B.n389 B.n388 585
R1626 B.n761 B.n760 585
R1627 B.n762 B.n761 585
R1628 B.n383 B.n382 585
R1629 B.n384 B.n383 585
R1630 B.n771 B.n770 585
R1631 B.n770 B.n769 585
R1632 B.n772 B.n381 585
R1633 B.n768 B.n381 585
R1634 B.n774 B.n773 585
R1635 B.n775 B.n774 585
R1636 B.n376 B.n375 585
R1637 B.n377 B.n376 585
R1638 B.n784 B.n783 585
R1639 B.n783 B.n782 585
R1640 B.n785 B.n374 585
R1641 B.n374 B.n373 585
R1642 B.n787 B.n786 585
R1643 B.n788 B.n787 585
R1644 B.n2 B.n0 585
R1645 B.n4 B.n2 585
R1646 B.n3 B.n1 585
R1647 B.n849 B.n3 585
R1648 B.n847 B.n846 585
R1649 B.n848 B.n847 585
R1650 B.n845 B.n9 585
R1651 B.n9 B.n8 585
R1652 B.n844 B.n843 585
R1653 B.n843 B.n842 585
R1654 B.n11 B.n10 585
R1655 B.n841 B.n11 585
R1656 B.n839 B.n838 585
R1657 B.n840 B.n839 585
R1658 B.n837 B.n15 585
R1659 B.n18 B.n15 585
R1660 B.n836 B.n835 585
R1661 B.n835 B.n834 585
R1662 B.n17 B.n16 585
R1663 B.n833 B.n17 585
R1664 B.n831 B.n830 585
R1665 B.n832 B.n831 585
R1666 B.n829 B.n23 585
R1667 B.n23 B.n22 585
R1668 B.n828 B.n827 585
R1669 B.n827 B.n826 585
R1670 B.n25 B.n24 585
R1671 B.n825 B.n25 585
R1672 B.n823 B.n822 585
R1673 B.n824 B.n823 585
R1674 B.n821 B.n30 585
R1675 B.n30 B.n29 585
R1676 B.n820 B.n819 585
R1677 B.n819 B.n818 585
R1678 B.n32 B.n31 585
R1679 B.n817 B.n32 585
R1680 B.n852 B.n851 585
R1681 B.n851 B.n850 585
R1682 B.n735 B.n399 478.086
R1683 B.n107 B.n32 478.086
R1684 B.n739 B.n401 478.086
R1685 B.n815 B.n34 478.086
R1686 B.n472 B.t7 418.332
R1687 B.n102 B.t16 418.332
R1688 B.n470 B.t10 418.332
R1689 B.n104 B.t13 418.332
R1690 B.n473 B.t6 398.745
R1691 B.n103 B.t17 398.745
R1692 B.n471 B.t9 398.745
R1693 B.n105 B.t14 398.745
R1694 B.n816 B.n100 256.663
R1695 B.n816 B.n99 256.663
R1696 B.n816 B.n98 256.663
R1697 B.n816 B.n97 256.663
R1698 B.n816 B.n96 256.663
R1699 B.n816 B.n95 256.663
R1700 B.n816 B.n94 256.663
R1701 B.n816 B.n93 256.663
R1702 B.n816 B.n92 256.663
R1703 B.n816 B.n91 256.663
R1704 B.n816 B.n90 256.663
R1705 B.n816 B.n89 256.663
R1706 B.n816 B.n88 256.663
R1707 B.n816 B.n87 256.663
R1708 B.n816 B.n86 256.663
R1709 B.n816 B.n85 256.663
R1710 B.n816 B.n84 256.663
R1711 B.n816 B.n83 256.663
R1712 B.n816 B.n82 256.663
R1713 B.n816 B.n81 256.663
R1714 B.n816 B.n80 256.663
R1715 B.n816 B.n79 256.663
R1716 B.n816 B.n78 256.663
R1717 B.n816 B.n77 256.663
R1718 B.n816 B.n76 256.663
R1719 B.n816 B.n75 256.663
R1720 B.n816 B.n74 256.663
R1721 B.n816 B.n73 256.663
R1722 B.n816 B.n72 256.663
R1723 B.n816 B.n71 256.663
R1724 B.n816 B.n70 256.663
R1725 B.n816 B.n69 256.663
R1726 B.n816 B.n68 256.663
R1727 B.n816 B.n67 256.663
R1728 B.n816 B.n66 256.663
R1729 B.n816 B.n65 256.663
R1730 B.n816 B.n64 256.663
R1731 B.n816 B.n63 256.663
R1732 B.n816 B.n62 256.663
R1733 B.n816 B.n61 256.663
R1734 B.n816 B.n60 256.663
R1735 B.n816 B.n59 256.663
R1736 B.n816 B.n58 256.663
R1737 B.n816 B.n57 256.663
R1738 B.n816 B.n56 256.663
R1739 B.n816 B.n55 256.663
R1740 B.n816 B.n54 256.663
R1741 B.n816 B.n53 256.663
R1742 B.n816 B.n52 256.663
R1743 B.n816 B.n51 256.663
R1744 B.n816 B.n50 256.663
R1745 B.n816 B.n49 256.663
R1746 B.n816 B.n48 256.663
R1747 B.n816 B.n47 256.663
R1748 B.n816 B.n46 256.663
R1749 B.n816 B.n45 256.663
R1750 B.n816 B.n44 256.663
R1751 B.n816 B.n43 256.663
R1752 B.n816 B.n42 256.663
R1753 B.n816 B.n41 256.663
R1754 B.n816 B.n40 256.663
R1755 B.n816 B.n39 256.663
R1756 B.n816 B.n38 256.663
R1757 B.n816 B.n37 256.663
R1758 B.n816 B.n36 256.663
R1759 B.n816 B.n35 256.663
R1760 B.n737 B.n736 256.663
R1761 B.n737 B.n404 256.663
R1762 B.n737 B.n405 256.663
R1763 B.n737 B.n406 256.663
R1764 B.n737 B.n407 256.663
R1765 B.n737 B.n408 256.663
R1766 B.n737 B.n409 256.663
R1767 B.n737 B.n410 256.663
R1768 B.n737 B.n411 256.663
R1769 B.n737 B.n412 256.663
R1770 B.n737 B.n413 256.663
R1771 B.n737 B.n414 256.663
R1772 B.n737 B.n415 256.663
R1773 B.n737 B.n416 256.663
R1774 B.n737 B.n417 256.663
R1775 B.n737 B.n418 256.663
R1776 B.n737 B.n419 256.663
R1777 B.n737 B.n420 256.663
R1778 B.n737 B.n421 256.663
R1779 B.n737 B.n422 256.663
R1780 B.n737 B.n423 256.663
R1781 B.n737 B.n424 256.663
R1782 B.n737 B.n425 256.663
R1783 B.n737 B.n426 256.663
R1784 B.n737 B.n427 256.663
R1785 B.n737 B.n428 256.663
R1786 B.n737 B.n429 256.663
R1787 B.n737 B.n430 256.663
R1788 B.n737 B.n431 256.663
R1789 B.n737 B.n432 256.663
R1790 B.n737 B.n433 256.663
R1791 B.n737 B.n434 256.663
R1792 B.n737 B.n435 256.663
R1793 B.n737 B.n436 256.663
R1794 B.n737 B.n437 256.663
R1795 B.n737 B.n438 256.663
R1796 B.n737 B.n439 256.663
R1797 B.n737 B.n440 256.663
R1798 B.n737 B.n441 256.663
R1799 B.n737 B.n442 256.663
R1800 B.n737 B.n443 256.663
R1801 B.n737 B.n444 256.663
R1802 B.n737 B.n445 256.663
R1803 B.n737 B.n446 256.663
R1804 B.n737 B.n447 256.663
R1805 B.n737 B.n448 256.663
R1806 B.n737 B.n449 256.663
R1807 B.n737 B.n450 256.663
R1808 B.n737 B.n451 256.663
R1809 B.n737 B.n452 256.663
R1810 B.n737 B.n453 256.663
R1811 B.n737 B.n454 256.663
R1812 B.n737 B.n455 256.663
R1813 B.n737 B.n456 256.663
R1814 B.n737 B.n457 256.663
R1815 B.n737 B.n458 256.663
R1816 B.n737 B.n459 256.663
R1817 B.n737 B.n460 256.663
R1818 B.n737 B.n461 256.663
R1819 B.n737 B.n462 256.663
R1820 B.n737 B.n463 256.663
R1821 B.n737 B.n464 256.663
R1822 B.n737 B.n465 256.663
R1823 B.n737 B.n466 256.663
R1824 B.n737 B.n467 256.663
R1825 B.n738 B.n737 256.663
R1826 B.n745 B.n399 163.367
R1827 B.n745 B.n397 163.367
R1828 B.n749 B.n397 163.367
R1829 B.n749 B.n391 163.367
R1830 B.n757 B.n391 163.367
R1831 B.n757 B.n389 163.367
R1832 B.n761 B.n389 163.367
R1833 B.n761 B.n383 163.367
R1834 B.n770 B.n383 163.367
R1835 B.n770 B.n381 163.367
R1836 B.n774 B.n381 163.367
R1837 B.n774 B.n376 163.367
R1838 B.n783 B.n376 163.367
R1839 B.n783 B.n374 163.367
R1840 B.n787 B.n374 163.367
R1841 B.n787 B.n2 163.367
R1842 B.n851 B.n2 163.367
R1843 B.n851 B.n3 163.367
R1844 B.n847 B.n3 163.367
R1845 B.n847 B.n9 163.367
R1846 B.n843 B.n9 163.367
R1847 B.n843 B.n11 163.367
R1848 B.n839 B.n11 163.367
R1849 B.n839 B.n15 163.367
R1850 B.n835 B.n15 163.367
R1851 B.n835 B.n17 163.367
R1852 B.n831 B.n17 163.367
R1853 B.n831 B.n23 163.367
R1854 B.n827 B.n23 163.367
R1855 B.n827 B.n25 163.367
R1856 B.n823 B.n25 163.367
R1857 B.n823 B.n30 163.367
R1858 B.n819 B.n30 163.367
R1859 B.n819 B.n32 163.367
R1860 B.n469 B.n468 163.367
R1861 B.n730 B.n468 163.367
R1862 B.n728 B.n727 163.367
R1863 B.n724 B.n723 163.367
R1864 B.n720 B.n719 163.367
R1865 B.n716 B.n715 163.367
R1866 B.n712 B.n711 163.367
R1867 B.n708 B.n707 163.367
R1868 B.n704 B.n703 163.367
R1869 B.n700 B.n699 163.367
R1870 B.n696 B.n695 163.367
R1871 B.n692 B.n691 163.367
R1872 B.n688 B.n687 163.367
R1873 B.n684 B.n683 163.367
R1874 B.n680 B.n679 163.367
R1875 B.n676 B.n675 163.367
R1876 B.n672 B.n671 163.367
R1877 B.n668 B.n667 163.367
R1878 B.n664 B.n663 163.367
R1879 B.n660 B.n659 163.367
R1880 B.n656 B.n655 163.367
R1881 B.n652 B.n651 163.367
R1882 B.n648 B.n647 163.367
R1883 B.n644 B.n643 163.367
R1884 B.n640 B.n639 163.367
R1885 B.n636 B.n635 163.367
R1886 B.n632 B.n631 163.367
R1887 B.n628 B.n627 163.367
R1888 B.n624 B.n623 163.367
R1889 B.n620 B.n619 163.367
R1890 B.n616 B.n615 163.367
R1891 B.n611 B.n610 163.367
R1892 B.n607 B.n606 163.367
R1893 B.n603 B.n602 163.367
R1894 B.n599 B.n598 163.367
R1895 B.n595 B.n594 163.367
R1896 B.n591 B.n590 163.367
R1897 B.n587 B.n586 163.367
R1898 B.n583 B.n582 163.367
R1899 B.n579 B.n578 163.367
R1900 B.n575 B.n574 163.367
R1901 B.n571 B.n570 163.367
R1902 B.n567 B.n566 163.367
R1903 B.n563 B.n562 163.367
R1904 B.n559 B.n558 163.367
R1905 B.n555 B.n554 163.367
R1906 B.n551 B.n550 163.367
R1907 B.n547 B.n546 163.367
R1908 B.n543 B.n542 163.367
R1909 B.n539 B.n538 163.367
R1910 B.n535 B.n534 163.367
R1911 B.n531 B.n530 163.367
R1912 B.n527 B.n526 163.367
R1913 B.n523 B.n522 163.367
R1914 B.n519 B.n518 163.367
R1915 B.n515 B.n514 163.367
R1916 B.n511 B.n510 163.367
R1917 B.n507 B.n506 163.367
R1918 B.n503 B.n502 163.367
R1919 B.n499 B.n498 163.367
R1920 B.n495 B.n494 163.367
R1921 B.n491 B.n490 163.367
R1922 B.n487 B.n486 163.367
R1923 B.n483 B.n482 163.367
R1924 B.n479 B.n478 163.367
R1925 B.n475 B.n403 163.367
R1926 B.n743 B.n401 163.367
R1927 B.n743 B.n394 163.367
R1928 B.n751 B.n394 163.367
R1929 B.n751 B.n392 163.367
R1930 B.n755 B.n392 163.367
R1931 B.n755 B.n387 163.367
R1932 B.n763 B.n387 163.367
R1933 B.n763 B.n385 163.367
R1934 B.n767 B.n385 163.367
R1935 B.n767 B.n380 163.367
R1936 B.n776 B.n380 163.367
R1937 B.n776 B.n378 163.367
R1938 B.n781 B.n378 163.367
R1939 B.n781 B.n372 163.367
R1940 B.n789 B.n372 163.367
R1941 B.n790 B.n789 163.367
R1942 B.n790 B.n5 163.367
R1943 B.n6 B.n5 163.367
R1944 B.n7 B.n6 163.367
R1945 B.n795 B.n7 163.367
R1946 B.n795 B.n12 163.367
R1947 B.n13 B.n12 163.367
R1948 B.n14 B.n13 163.367
R1949 B.n800 B.n14 163.367
R1950 B.n800 B.n19 163.367
R1951 B.n20 B.n19 163.367
R1952 B.n21 B.n20 163.367
R1953 B.n805 B.n21 163.367
R1954 B.n805 B.n26 163.367
R1955 B.n27 B.n26 163.367
R1956 B.n28 B.n27 163.367
R1957 B.n810 B.n28 163.367
R1958 B.n810 B.n33 163.367
R1959 B.n34 B.n33 163.367
R1960 B.n111 B.n110 163.367
R1961 B.n115 B.n114 163.367
R1962 B.n119 B.n118 163.367
R1963 B.n123 B.n122 163.367
R1964 B.n127 B.n126 163.367
R1965 B.n131 B.n130 163.367
R1966 B.n135 B.n134 163.367
R1967 B.n139 B.n138 163.367
R1968 B.n143 B.n142 163.367
R1969 B.n147 B.n146 163.367
R1970 B.n151 B.n150 163.367
R1971 B.n155 B.n154 163.367
R1972 B.n159 B.n158 163.367
R1973 B.n163 B.n162 163.367
R1974 B.n167 B.n166 163.367
R1975 B.n171 B.n170 163.367
R1976 B.n175 B.n174 163.367
R1977 B.n179 B.n178 163.367
R1978 B.n183 B.n182 163.367
R1979 B.n187 B.n186 163.367
R1980 B.n191 B.n190 163.367
R1981 B.n195 B.n194 163.367
R1982 B.n199 B.n198 163.367
R1983 B.n203 B.n202 163.367
R1984 B.n207 B.n206 163.367
R1985 B.n211 B.n210 163.367
R1986 B.n215 B.n214 163.367
R1987 B.n219 B.n218 163.367
R1988 B.n223 B.n222 163.367
R1989 B.n227 B.n226 163.367
R1990 B.n231 B.n230 163.367
R1991 B.n235 B.n234 163.367
R1992 B.n239 B.n238 163.367
R1993 B.n243 B.n242 163.367
R1994 B.n247 B.n246 163.367
R1995 B.n252 B.n251 163.367
R1996 B.n256 B.n255 163.367
R1997 B.n260 B.n259 163.367
R1998 B.n264 B.n263 163.367
R1999 B.n268 B.n267 163.367
R2000 B.n272 B.n271 163.367
R2001 B.n276 B.n275 163.367
R2002 B.n280 B.n279 163.367
R2003 B.n284 B.n283 163.367
R2004 B.n288 B.n287 163.367
R2005 B.n292 B.n291 163.367
R2006 B.n296 B.n295 163.367
R2007 B.n300 B.n299 163.367
R2008 B.n304 B.n303 163.367
R2009 B.n308 B.n307 163.367
R2010 B.n312 B.n311 163.367
R2011 B.n316 B.n315 163.367
R2012 B.n320 B.n319 163.367
R2013 B.n324 B.n323 163.367
R2014 B.n328 B.n327 163.367
R2015 B.n332 B.n331 163.367
R2016 B.n336 B.n335 163.367
R2017 B.n340 B.n339 163.367
R2018 B.n344 B.n343 163.367
R2019 B.n348 B.n347 163.367
R2020 B.n352 B.n351 163.367
R2021 B.n356 B.n355 163.367
R2022 B.n360 B.n359 163.367
R2023 B.n364 B.n363 163.367
R2024 B.n368 B.n367 163.367
R2025 B.n815 B.n101 163.367
R2026 B.n736 B.n735 71.676
R2027 B.n730 B.n404 71.676
R2028 B.n727 B.n405 71.676
R2029 B.n723 B.n406 71.676
R2030 B.n719 B.n407 71.676
R2031 B.n715 B.n408 71.676
R2032 B.n711 B.n409 71.676
R2033 B.n707 B.n410 71.676
R2034 B.n703 B.n411 71.676
R2035 B.n699 B.n412 71.676
R2036 B.n695 B.n413 71.676
R2037 B.n691 B.n414 71.676
R2038 B.n687 B.n415 71.676
R2039 B.n683 B.n416 71.676
R2040 B.n679 B.n417 71.676
R2041 B.n675 B.n418 71.676
R2042 B.n671 B.n419 71.676
R2043 B.n667 B.n420 71.676
R2044 B.n663 B.n421 71.676
R2045 B.n659 B.n422 71.676
R2046 B.n655 B.n423 71.676
R2047 B.n651 B.n424 71.676
R2048 B.n647 B.n425 71.676
R2049 B.n643 B.n426 71.676
R2050 B.n639 B.n427 71.676
R2051 B.n635 B.n428 71.676
R2052 B.n631 B.n429 71.676
R2053 B.n627 B.n430 71.676
R2054 B.n623 B.n431 71.676
R2055 B.n619 B.n432 71.676
R2056 B.n615 B.n433 71.676
R2057 B.n610 B.n434 71.676
R2058 B.n606 B.n435 71.676
R2059 B.n602 B.n436 71.676
R2060 B.n598 B.n437 71.676
R2061 B.n594 B.n438 71.676
R2062 B.n590 B.n439 71.676
R2063 B.n586 B.n440 71.676
R2064 B.n582 B.n441 71.676
R2065 B.n578 B.n442 71.676
R2066 B.n574 B.n443 71.676
R2067 B.n570 B.n444 71.676
R2068 B.n566 B.n445 71.676
R2069 B.n562 B.n446 71.676
R2070 B.n558 B.n447 71.676
R2071 B.n554 B.n448 71.676
R2072 B.n550 B.n449 71.676
R2073 B.n546 B.n450 71.676
R2074 B.n542 B.n451 71.676
R2075 B.n538 B.n452 71.676
R2076 B.n534 B.n453 71.676
R2077 B.n530 B.n454 71.676
R2078 B.n526 B.n455 71.676
R2079 B.n522 B.n456 71.676
R2080 B.n518 B.n457 71.676
R2081 B.n514 B.n458 71.676
R2082 B.n510 B.n459 71.676
R2083 B.n506 B.n460 71.676
R2084 B.n502 B.n461 71.676
R2085 B.n498 B.n462 71.676
R2086 B.n494 B.n463 71.676
R2087 B.n490 B.n464 71.676
R2088 B.n486 B.n465 71.676
R2089 B.n482 B.n466 71.676
R2090 B.n478 B.n467 71.676
R2091 B.n738 B.n403 71.676
R2092 B.n107 B.n35 71.676
R2093 B.n111 B.n36 71.676
R2094 B.n115 B.n37 71.676
R2095 B.n119 B.n38 71.676
R2096 B.n123 B.n39 71.676
R2097 B.n127 B.n40 71.676
R2098 B.n131 B.n41 71.676
R2099 B.n135 B.n42 71.676
R2100 B.n139 B.n43 71.676
R2101 B.n143 B.n44 71.676
R2102 B.n147 B.n45 71.676
R2103 B.n151 B.n46 71.676
R2104 B.n155 B.n47 71.676
R2105 B.n159 B.n48 71.676
R2106 B.n163 B.n49 71.676
R2107 B.n167 B.n50 71.676
R2108 B.n171 B.n51 71.676
R2109 B.n175 B.n52 71.676
R2110 B.n179 B.n53 71.676
R2111 B.n183 B.n54 71.676
R2112 B.n187 B.n55 71.676
R2113 B.n191 B.n56 71.676
R2114 B.n195 B.n57 71.676
R2115 B.n199 B.n58 71.676
R2116 B.n203 B.n59 71.676
R2117 B.n207 B.n60 71.676
R2118 B.n211 B.n61 71.676
R2119 B.n215 B.n62 71.676
R2120 B.n219 B.n63 71.676
R2121 B.n223 B.n64 71.676
R2122 B.n227 B.n65 71.676
R2123 B.n231 B.n66 71.676
R2124 B.n235 B.n67 71.676
R2125 B.n239 B.n68 71.676
R2126 B.n243 B.n69 71.676
R2127 B.n247 B.n70 71.676
R2128 B.n252 B.n71 71.676
R2129 B.n256 B.n72 71.676
R2130 B.n260 B.n73 71.676
R2131 B.n264 B.n74 71.676
R2132 B.n268 B.n75 71.676
R2133 B.n272 B.n76 71.676
R2134 B.n276 B.n77 71.676
R2135 B.n280 B.n78 71.676
R2136 B.n284 B.n79 71.676
R2137 B.n288 B.n80 71.676
R2138 B.n292 B.n81 71.676
R2139 B.n296 B.n82 71.676
R2140 B.n300 B.n83 71.676
R2141 B.n304 B.n84 71.676
R2142 B.n308 B.n85 71.676
R2143 B.n312 B.n86 71.676
R2144 B.n316 B.n87 71.676
R2145 B.n320 B.n88 71.676
R2146 B.n324 B.n89 71.676
R2147 B.n328 B.n90 71.676
R2148 B.n332 B.n91 71.676
R2149 B.n336 B.n92 71.676
R2150 B.n340 B.n93 71.676
R2151 B.n344 B.n94 71.676
R2152 B.n348 B.n95 71.676
R2153 B.n352 B.n96 71.676
R2154 B.n356 B.n97 71.676
R2155 B.n360 B.n98 71.676
R2156 B.n364 B.n99 71.676
R2157 B.n368 B.n100 71.676
R2158 B.n101 B.n100 71.676
R2159 B.n367 B.n99 71.676
R2160 B.n363 B.n98 71.676
R2161 B.n359 B.n97 71.676
R2162 B.n355 B.n96 71.676
R2163 B.n351 B.n95 71.676
R2164 B.n347 B.n94 71.676
R2165 B.n343 B.n93 71.676
R2166 B.n339 B.n92 71.676
R2167 B.n335 B.n91 71.676
R2168 B.n331 B.n90 71.676
R2169 B.n327 B.n89 71.676
R2170 B.n323 B.n88 71.676
R2171 B.n319 B.n87 71.676
R2172 B.n315 B.n86 71.676
R2173 B.n311 B.n85 71.676
R2174 B.n307 B.n84 71.676
R2175 B.n303 B.n83 71.676
R2176 B.n299 B.n82 71.676
R2177 B.n295 B.n81 71.676
R2178 B.n291 B.n80 71.676
R2179 B.n287 B.n79 71.676
R2180 B.n283 B.n78 71.676
R2181 B.n279 B.n77 71.676
R2182 B.n275 B.n76 71.676
R2183 B.n271 B.n75 71.676
R2184 B.n267 B.n74 71.676
R2185 B.n263 B.n73 71.676
R2186 B.n259 B.n72 71.676
R2187 B.n255 B.n71 71.676
R2188 B.n251 B.n70 71.676
R2189 B.n246 B.n69 71.676
R2190 B.n242 B.n68 71.676
R2191 B.n238 B.n67 71.676
R2192 B.n234 B.n66 71.676
R2193 B.n230 B.n65 71.676
R2194 B.n226 B.n64 71.676
R2195 B.n222 B.n63 71.676
R2196 B.n218 B.n62 71.676
R2197 B.n214 B.n61 71.676
R2198 B.n210 B.n60 71.676
R2199 B.n206 B.n59 71.676
R2200 B.n202 B.n58 71.676
R2201 B.n198 B.n57 71.676
R2202 B.n194 B.n56 71.676
R2203 B.n190 B.n55 71.676
R2204 B.n186 B.n54 71.676
R2205 B.n182 B.n53 71.676
R2206 B.n178 B.n52 71.676
R2207 B.n174 B.n51 71.676
R2208 B.n170 B.n50 71.676
R2209 B.n166 B.n49 71.676
R2210 B.n162 B.n48 71.676
R2211 B.n158 B.n47 71.676
R2212 B.n154 B.n46 71.676
R2213 B.n150 B.n45 71.676
R2214 B.n146 B.n44 71.676
R2215 B.n142 B.n43 71.676
R2216 B.n138 B.n42 71.676
R2217 B.n134 B.n41 71.676
R2218 B.n130 B.n40 71.676
R2219 B.n126 B.n39 71.676
R2220 B.n122 B.n38 71.676
R2221 B.n118 B.n37 71.676
R2222 B.n114 B.n36 71.676
R2223 B.n110 B.n35 71.676
R2224 B.n736 B.n469 71.676
R2225 B.n728 B.n404 71.676
R2226 B.n724 B.n405 71.676
R2227 B.n720 B.n406 71.676
R2228 B.n716 B.n407 71.676
R2229 B.n712 B.n408 71.676
R2230 B.n708 B.n409 71.676
R2231 B.n704 B.n410 71.676
R2232 B.n700 B.n411 71.676
R2233 B.n696 B.n412 71.676
R2234 B.n692 B.n413 71.676
R2235 B.n688 B.n414 71.676
R2236 B.n684 B.n415 71.676
R2237 B.n680 B.n416 71.676
R2238 B.n676 B.n417 71.676
R2239 B.n672 B.n418 71.676
R2240 B.n668 B.n419 71.676
R2241 B.n664 B.n420 71.676
R2242 B.n660 B.n421 71.676
R2243 B.n656 B.n422 71.676
R2244 B.n652 B.n423 71.676
R2245 B.n648 B.n424 71.676
R2246 B.n644 B.n425 71.676
R2247 B.n640 B.n426 71.676
R2248 B.n636 B.n427 71.676
R2249 B.n632 B.n428 71.676
R2250 B.n628 B.n429 71.676
R2251 B.n624 B.n430 71.676
R2252 B.n620 B.n431 71.676
R2253 B.n616 B.n432 71.676
R2254 B.n611 B.n433 71.676
R2255 B.n607 B.n434 71.676
R2256 B.n603 B.n435 71.676
R2257 B.n599 B.n436 71.676
R2258 B.n595 B.n437 71.676
R2259 B.n591 B.n438 71.676
R2260 B.n587 B.n439 71.676
R2261 B.n583 B.n440 71.676
R2262 B.n579 B.n441 71.676
R2263 B.n575 B.n442 71.676
R2264 B.n571 B.n443 71.676
R2265 B.n567 B.n444 71.676
R2266 B.n563 B.n445 71.676
R2267 B.n559 B.n446 71.676
R2268 B.n555 B.n447 71.676
R2269 B.n551 B.n448 71.676
R2270 B.n547 B.n449 71.676
R2271 B.n543 B.n450 71.676
R2272 B.n539 B.n451 71.676
R2273 B.n535 B.n452 71.676
R2274 B.n531 B.n453 71.676
R2275 B.n527 B.n454 71.676
R2276 B.n523 B.n455 71.676
R2277 B.n519 B.n456 71.676
R2278 B.n515 B.n457 71.676
R2279 B.n511 B.n458 71.676
R2280 B.n507 B.n459 71.676
R2281 B.n503 B.n460 71.676
R2282 B.n499 B.n461 71.676
R2283 B.n495 B.n462 71.676
R2284 B.n491 B.n463 71.676
R2285 B.n487 B.n464 71.676
R2286 B.n483 B.n465 71.676
R2287 B.n479 B.n466 71.676
R2288 B.n475 B.n467 71.676
R2289 B.n739 B.n738 71.676
R2290 B.n474 B.n473 59.5399
R2291 B.n613 B.n471 59.5399
R2292 B.n106 B.n105 59.5399
R2293 B.n249 B.n103 59.5399
R2294 B.n737 B.n400 57.1612
R2295 B.n817 B.n816 57.1612
R2296 B.n744 B.n400 31.0959
R2297 B.n744 B.n395 31.0959
R2298 B.n750 B.n395 31.0959
R2299 B.n750 B.n396 31.0959
R2300 B.n756 B.n388 31.0959
R2301 B.n762 B.n388 31.0959
R2302 B.n762 B.n384 31.0959
R2303 B.n769 B.n384 31.0959
R2304 B.n769 B.n768 31.0959
R2305 B.n775 B.n377 31.0959
R2306 B.n782 B.n377 31.0959
R2307 B.n788 B.n373 31.0959
R2308 B.n788 B.n4 31.0959
R2309 B.n850 B.n4 31.0959
R2310 B.n850 B.n849 31.0959
R2311 B.n849 B.n848 31.0959
R2312 B.n848 B.n8 31.0959
R2313 B.n842 B.n841 31.0959
R2314 B.n841 B.n840 31.0959
R2315 B.n834 B.n18 31.0959
R2316 B.n834 B.n833 31.0959
R2317 B.n833 B.n832 31.0959
R2318 B.n832 B.n22 31.0959
R2319 B.n826 B.n22 31.0959
R2320 B.n825 B.n824 31.0959
R2321 B.n824 B.n29 31.0959
R2322 B.n818 B.n29 31.0959
R2323 B.n818 B.n817 31.0959
R2324 B.n108 B.n31 31.0639
R2325 B.n814 B.n813 31.0639
R2326 B.n741 B.n740 31.0639
R2327 B.n734 B.n398 31.0639
R2328 B.n768 B.t2 29.2668
R2329 B.n18 B.t0 29.2668
R2330 B.n782 B.t3 28.3522
R2331 B.n842 B.t1 28.3522
R2332 B.n396 B.t5 23.7793
R2333 B.t12 B.n825 23.7793
R2334 B.n473 B.n472 19.5884
R2335 B.n471 B.n470 19.5884
R2336 B.n105 B.n104 19.5884
R2337 B.n103 B.n102 19.5884
R2338 B B.n852 18.0485
R2339 B.n109 B.n108 10.6151
R2340 B.n112 B.n109 10.6151
R2341 B.n113 B.n112 10.6151
R2342 B.n116 B.n113 10.6151
R2343 B.n117 B.n116 10.6151
R2344 B.n120 B.n117 10.6151
R2345 B.n121 B.n120 10.6151
R2346 B.n124 B.n121 10.6151
R2347 B.n125 B.n124 10.6151
R2348 B.n128 B.n125 10.6151
R2349 B.n129 B.n128 10.6151
R2350 B.n132 B.n129 10.6151
R2351 B.n133 B.n132 10.6151
R2352 B.n136 B.n133 10.6151
R2353 B.n137 B.n136 10.6151
R2354 B.n140 B.n137 10.6151
R2355 B.n141 B.n140 10.6151
R2356 B.n144 B.n141 10.6151
R2357 B.n145 B.n144 10.6151
R2358 B.n148 B.n145 10.6151
R2359 B.n149 B.n148 10.6151
R2360 B.n152 B.n149 10.6151
R2361 B.n153 B.n152 10.6151
R2362 B.n156 B.n153 10.6151
R2363 B.n157 B.n156 10.6151
R2364 B.n160 B.n157 10.6151
R2365 B.n161 B.n160 10.6151
R2366 B.n164 B.n161 10.6151
R2367 B.n165 B.n164 10.6151
R2368 B.n168 B.n165 10.6151
R2369 B.n169 B.n168 10.6151
R2370 B.n172 B.n169 10.6151
R2371 B.n173 B.n172 10.6151
R2372 B.n176 B.n173 10.6151
R2373 B.n177 B.n176 10.6151
R2374 B.n180 B.n177 10.6151
R2375 B.n181 B.n180 10.6151
R2376 B.n184 B.n181 10.6151
R2377 B.n185 B.n184 10.6151
R2378 B.n188 B.n185 10.6151
R2379 B.n189 B.n188 10.6151
R2380 B.n192 B.n189 10.6151
R2381 B.n193 B.n192 10.6151
R2382 B.n196 B.n193 10.6151
R2383 B.n197 B.n196 10.6151
R2384 B.n200 B.n197 10.6151
R2385 B.n201 B.n200 10.6151
R2386 B.n204 B.n201 10.6151
R2387 B.n205 B.n204 10.6151
R2388 B.n208 B.n205 10.6151
R2389 B.n209 B.n208 10.6151
R2390 B.n212 B.n209 10.6151
R2391 B.n213 B.n212 10.6151
R2392 B.n216 B.n213 10.6151
R2393 B.n217 B.n216 10.6151
R2394 B.n220 B.n217 10.6151
R2395 B.n221 B.n220 10.6151
R2396 B.n224 B.n221 10.6151
R2397 B.n225 B.n224 10.6151
R2398 B.n228 B.n225 10.6151
R2399 B.n229 B.n228 10.6151
R2400 B.n233 B.n232 10.6151
R2401 B.n236 B.n233 10.6151
R2402 B.n237 B.n236 10.6151
R2403 B.n240 B.n237 10.6151
R2404 B.n241 B.n240 10.6151
R2405 B.n244 B.n241 10.6151
R2406 B.n245 B.n244 10.6151
R2407 B.n248 B.n245 10.6151
R2408 B.n253 B.n250 10.6151
R2409 B.n254 B.n253 10.6151
R2410 B.n257 B.n254 10.6151
R2411 B.n258 B.n257 10.6151
R2412 B.n261 B.n258 10.6151
R2413 B.n262 B.n261 10.6151
R2414 B.n265 B.n262 10.6151
R2415 B.n266 B.n265 10.6151
R2416 B.n269 B.n266 10.6151
R2417 B.n270 B.n269 10.6151
R2418 B.n273 B.n270 10.6151
R2419 B.n274 B.n273 10.6151
R2420 B.n277 B.n274 10.6151
R2421 B.n278 B.n277 10.6151
R2422 B.n281 B.n278 10.6151
R2423 B.n282 B.n281 10.6151
R2424 B.n285 B.n282 10.6151
R2425 B.n286 B.n285 10.6151
R2426 B.n289 B.n286 10.6151
R2427 B.n290 B.n289 10.6151
R2428 B.n293 B.n290 10.6151
R2429 B.n294 B.n293 10.6151
R2430 B.n297 B.n294 10.6151
R2431 B.n298 B.n297 10.6151
R2432 B.n301 B.n298 10.6151
R2433 B.n302 B.n301 10.6151
R2434 B.n305 B.n302 10.6151
R2435 B.n306 B.n305 10.6151
R2436 B.n309 B.n306 10.6151
R2437 B.n310 B.n309 10.6151
R2438 B.n313 B.n310 10.6151
R2439 B.n314 B.n313 10.6151
R2440 B.n317 B.n314 10.6151
R2441 B.n318 B.n317 10.6151
R2442 B.n321 B.n318 10.6151
R2443 B.n322 B.n321 10.6151
R2444 B.n325 B.n322 10.6151
R2445 B.n326 B.n325 10.6151
R2446 B.n329 B.n326 10.6151
R2447 B.n330 B.n329 10.6151
R2448 B.n333 B.n330 10.6151
R2449 B.n334 B.n333 10.6151
R2450 B.n337 B.n334 10.6151
R2451 B.n338 B.n337 10.6151
R2452 B.n341 B.n338 10.6151
R2453 B.n342 B.n341 10.6151
R2454 B.n345 B.n342 10.6151
R2455 B.n346 B.n345 10.6151
R2456 B.n349 B.n346 10.6151
R2457 B.n350 B.n349 10.6151
R2458 B.n353 B.n350 10.6151
R2459 B.n354 B.n353 10.6151
R2460 B.n357 B.n354 10.6151
R2461 B.n358 B.n357 10.6151
R2462 B.n361 B.n358 10.6151
R2463 B.n362 B.n361 10.6151
R2464 B.n365 B.n362 10.6151
R2465 B.n366 B.n365 10.6151
R2466 B.n369 B.n366 10.6151
R2467 B.n370 B.n369 10.6151
R2468 B.n814 B.n370 10.6151
R2469 B.n742 B.n741 10.6151
R2470 B.n742 B.n393 10.6151
R2471 B.n752 B.n393 10.6151
R2472 B.n753 B.n752 10.6151
R2473 B.n754 B.n753 10.6151
R2474 B.n754 B.n386 10.6151
R2475 B.n764 B.n386 10.6151
R2476 B.n765 B.n764 10.6151
R2477 B.n766 B.n765 10.6151
R2478 B.n766 B.n379 10.6151
R2479 B.n777 B.n379 10.6151
R2480 B.n778 B.n777 10.6151
R2481 B.n780 B.n778 10.6151
R2482 B.n780 B.n779 10.6151
R2483 B.n779 B.n371 10.6151
R2484 B.n791 B.n371 10.6151
R2485 B.n792 B.n791 10.6151
R2486 B.n793 B.n792 10.6151
R2487 B.n794 B.n793 10.6151
R2488 B.n796 B.n794 10.6151
R2489 B.n797 B.n796 10.6151
R2490 B.n798 B.n797 10.6151
R2491 B.n799 B.n798 10.6151
R2492 B.n801 B.n799 10.6151
R2493 B.n802 B.n801 10.6151
R2494 B.n803 B.n802 10.6151
R2495 B.n804 B.n803 10.6151
R2496 B.n806 B.n804 10.6151
R2497 B.n807 B.n806 10.6151
R2498 B.n808 B.n807 10.6151
R2499 B.n809 B.n808 10.6151
R2500 B.n811 B.n809 10.6151
R2501 B.n812 B.n811 10.6151
R2502 B.n813 B.n812 10.6151
R2503 B.n734 B.n733 10.6151
R2504 B.n733 B.n732 10.6151
R2505 B.n732 B.n731 10.6151
R2506 B.n731 B.n729 10.6151
R2507 B.n729 B.n726 10.6151
R2508 B.n726 B.n725 10.6151
R2509 B.n725 B.n722 10.6151
R2510 B.n722 B.n721 10.6151
R2511 B.n721 B.n718 10.6151
R2512 B.n718 B.n717 10.6151
R2513 B.n717 B.n714 10.6151
R2514 B.n714 B.n713 10.6151
R2515 B.n713 B.n710 10.6151
R2516 B.n710 B.n709 10.6151
R2517 B.n709 B.n706 10.6151
R2518 B.n706 B.n705 10.6151
R2519 B.n705 B.n702 10.6151
R2520 B.n702 B.n701 10.6151
R2521 B.n701 B.n698 10.6151
R2522 B.n698 B.n697 10.6151
R2523 B.n697 B.n694 10.6151
R2524 B.n694 B.n693 10.6151
R2525 B.n693 B.n690 10.6151
R2526 B.n690 B.n689 10.6151
R2527 B.n689 B.n686 10.6151
R2528 B.n686 B.n685 10.6151
R2529 B.n685 B.n682 10.6151
R2530 B.n682 B.n681 10.6151
R2531 B.n681 B.n678 10.6151
R2532 B.n678 B.n677 10.6151
R2533 B.n677 B.n674 10.6151
R2534 B.n674 B.n673 10.6151
R2535 B.n673 B.n670 10.6151
R2536 B.n670 B.n669 10.6151
R2537 B.n669 B.n666 10.6151
R2538 B.n666 B.n665 10.6151
R2539 B.n665 B.n662 10.6151
R2540 B.n662 B.n661 10.6151
R2541 B.n661 B.n658 10.6151
R2542 B.n658 B.n657 10.6151
R2543 B.n657 B.n654 10.6151
R2544 B.n654 B.n653 10.6151
R2545 B.n653 B.n650 10.6151
R2546 B.n650 B.n649 10.6151
R2547 B.n649 B.n646 10.6151
R2548 B.n646 B.n645 10.6151
R2549 B.n645 B.n642 10.6151
R2550 B.n642 B.n641 10.6151
R2551 B.n641 B.n638 10.6151
R2552 B.n638 B.n637 10.6151
R2553 B.n637 B.n634 10.6151
R2554 B.n634 B.n633 10.6151
R2555 B.n633 B.n630 10.6151
R2556 B.n630 B.n629 10.6151
R2557 B.n629 B.n626 10.6151
R2558 B.n626 B.n625 10.6151
R2559 B.n625 B.n622 10.6151
R2560 B.n622 B.n621 10.6151
R2561 B.n621 B.n618 10.6151
R2562 B.n618 B.n617 10.6151
R2563 B.n617 B.n614 10.6151
R2564 B.n612 B.n609 10.6151
R2565 B.n609 B.n608 10.6151
R2566 B.n608 B.n605 10.6151
R2567 B.n605 B.n604 10.6151
R2568 B.n604 B.n601 10.6151
R2569 B.n601 B.n600 10.6151
R2570 B.n600 B.n597 10.6151
R2571 B.n597 B.n596 10.6151
R2572 B.n593 B.n592 10.6151
R2573 B.n592 B.n589 10.6151
R2574 B.n589 B.n588 10.6151
R2575 B.n588 B.n585 10.6151
R2576 B.n585 B.n584 10.6151
R2577 B.n584 B.n581 10.6151
R2578 B.n581 B.n580 10.6151
R2579 B.n580 B.n577 10.6151
R2580 B.n577 B.n576 10.6151
R2581 B.n576 B.n573 10.6151
R2582 B.n573 B.n572 10.6151
R2583 B.n572 B.n569 10.6151
R2584 B.n569 B.n568 10.6151
R2585 B.n568 B.n565 10.6151
R2586 B.n565 B.n564 10.6151
R2587 B.n564 B.n561 10.6151
R2588 B.n561 B.n560 10.6151
R2589 B.n560 B.n557 10.6151
R2590 B.n557 B.n556 10.6151
R2591 B.n556 B.n553 10.6151
R2592 B.n553 B.n552 10.6151
R2593 B.n552 B.n549 10.6151
R2594 B.n549 B.n548 10.6151
R2595 B.n548 B.n545 10.6151
R2596 B.n545 B.n544 10.6151
R2597 B.n544 B.n541 10.6151
R2598 B.n541 B.n540 10.6151
R2599 B.n540 B.n537 10.6151
R2600 B.n537 B.n536 10.6151
R2601 B.n536 B.n533 10.6151
R2602 B.n533 B.n532 10.6151
R2603 B.n532 B.n529 10.6151
R2604 B.n529 B.n528 10.6151
R2605 B.n528 B.n525 10.6151
R2606 B.n525 B.n524 10.6151
R2607 B.n524 B.n521 10.6151
R2608 B.n521 B.n520 10.6151
R2609 B.n520 B.n517 10.6151
R2610 B.n517 B.n516 10.6151
R2611 B.n516 B.n513 10.6151
R2612 B.n513 B.n512 10.6151
R2613 B.n512 B.n509 10.6151
R2614 B.n509 B.n508 10.6151
R2615 B.n508 B.n505 10.6151
R2616 B.n505 B.n504 10.6151
R2617 B.n504 B.n501 10.6151
R2618 B.n501 B.n500 10.6151
R2619 B.n500 B.n497 10.6151
R2620 B.n497 B.n496 10.6151
R2621 B.n496 B.n493 10.6151
R2622 B.n493 B.n492 10.6151
R2623 B.n492 B.n489 10.6151
R2624 B.n489 B.n488 10.6151
R2625 B.n488 B.n485 10.6151
R2626 B.n485 B.n484 10.6151
R2627 B.n484 B.n481 10.6151
R2628 B.n481 B.n480 10.6151
R2629 B.n480 B.n477 10.6151
R2630 B.n477 B.n476 10.6151
R2631 B.n476 B.n402 10.6151
R2632 B.n740 B.n402 10.6151
R2633 B.n746 B.n398 10.6151
R2634 B.n747 B.n746 10.6151
R2635 B.n748 B.n747 10.6151
R2636 B.n748 B.n390 10.6151
R2637 B.n758 B.n390 10.6151
R2638 B.n759 B.n758 10.6151
R2639 B.n760 B.n759 10.6151
R2640 B.n760 B.n382 10.6151
R2641 B.n771 B.n382 10.6151
R2642 B.n772 B.n771 10.6151
R2643 B.n773 B.n772 10.6151
R2644 B.n773 B.n375 10.6151
R2645 B.n784 B.n375 10.6151
R2646 B.n785 B.n784 10.6151
R2647 B.n786 B.n785 10.6151
R2648 B.n786 B.n0 10.6151
R2649 B.n846 B.n1 10.6151
R2650 B.n846 B.n845 10.6151
R2651 B.n845 B.n844 10.6151
R2652 B.n844 B.n10 10.6151
R2653 B.n838 B.n10 10.6151
R2654 B.n838 B.n837 10.6151
R2655 B.n837 B.n836 10.6151
R2656 B.n836 B.n16 10.6151
R2657 B.n830 B.n16 10.6151
R2658 B.n830 B.n829 10.6151
R2659 B.n829 B.n828 10.6151
R2660 B.n828 B.n24 10.6151
R2661 B.n822 B.n24 10.6151
R2662 B.n822 B.n821 10.6151
R2663 B.n821 B.n820 10.6151
R2664 B.n820 B.n31 10.6151
R2665 B.n756 B.t5 7.31707
R2666 B.n826 B.t12 7.31707
R2667 B.n232 B.n106 6.5566
R2668 B.n249 B.n248 6.5566
R2669 B.n613 B.n612 6.5566
R2670 B.n596 B.n474 6.5566
R2671 B.n229 B.n106 4.05904
R2672 B.n250 B.n249 4.05904
R2673 B.n614 B.n613 4.05904
R2674 B.n593 B.n474 4.05904
R2675 B.n852 B.n0 2.81026
R2676 B.n852 B.n1 2.81026
R2677 B.t3 B.n373 2.74421
R2678 B.t1 B.n8 2.74421
R2679 B.n775 B.t2 1.82964
R2680 B.n840 B.t0 1.82964
R2681 VP.n1 VP.t1 745.061
R2682 VP.n1 VP.t0 745.01
R2683 VP.n3 VP.t3 724.063
R2684 VP.n5 VP.t2 724.063
R2685 VP.n6 VP.n5 161.3
R2686 VP.n4 VP.n0 161.3
R2687 VP.n3 VP.n2 161.3
R2688 VP.n2 VP.n1 90.1318
R2689 VP.n4 VP.n3 24.1005
R2690 VP.n5 VP.n4 24.1005
R2691 VP.n2 VP.n0 0.189894
R2692 VP.n6 VP.n0 0.189894
R2693 VP VP.n6 0.0516364
R2694 VDD1 VDD1.n1 106.701
R2695 VDD1 VDD1.n0 63.717
R2696 VDD1.n0 VDD1.t2 1.05481
R2697 VDD1.n0 VDD1.t3 1.05481
R2698 VDD1.n1 VDD1.t0 1.05481
R2699 VDD1.n1 VDD1.t1 1.05481
C0 VP VTAIL 4.06237f
C1 VDD1 VDD2 0.561847f
C2 VN VTAIL 4.04826f
C3 VP VDD1 4.84887f
C4 VP VDD2 0.271604f
C5 VN VDD1 0.146737f
C6 VTAIL VDD1 9.91241f
C7 VN VDD2 4.72426f
C8 VTAIL VDD2 9.95375f
C9 VP VN 6.06823f
C10 VDD2 B 3.218584f
C11 VDD1 B 7.73539f
C12 VTAIL B 12.57909f
C13 VN B 9.11267f
C14 VP B 5.316017f
C15 VDD1.t2 B 0.420677f
C16 VDD1.t3 B 0.420677f
C17 VDD1.n0 B 3.84939f
C18 VDD1.t0 B 0.420677f
C19 VDD1.t1 B 0.420677f
C20 VDD1.n1 B 4.72126f
C21 VP.n0 B 0.050287f
C22 VP.t0 B 1.83968f
C23 VP.t1 B 1.83973f
C24 VP.n1 B 2.57806f
C25 VP.n2 B 3.62377f
C26 VP.t3 B 1.82046f
C27 VP.n3 B 0.679983f
C28 VP.n4 B 0.011411f
C29 VP.t2 B 1.82046f
C30 VP.n5 B 0.679983f
C31 VP.n6 B 0.03897f
C32 VTAIL.n0 B 0.008933f
C33 VTAIL.n1 B 0.020141f
C34 VTAIL.n2 B 0.009023f
C35 VTAIL.n3 B 0.015858f
C36 VTAIL.n4 B 0.008521f
C37 VTAIL.n5 B 0.020141f
C38 VTAIL.n6 B 0.009023f
C39 VTAIL.n7 B 0.015858f
C40 VTAIL.n8 B 0.008521f
C41 VTAIL.n9 B 0.020141f
C42 VTAIL.n10 B 0.009023f
C43 VTAIL.n11 B 0.015858f
C44 VTAIL.n12 B 0.008521f
C45 VTAIL.n13 B 0.020141f
C46 VTAIL.n14 B 0.009023f
C47 VTAIL.n15 B 0.015858f
C48 VTAIL.n16 B 0.008521f
C49 VTAIL.n17 B 0.020141f
C50 VTAIL.n18 B 0.009023f
C51 VTAIL.n19 B 0.015858f
C52 VTAIL.n20 B 0.008521f
C53 VTAIL.n21 B 0.020141f
C54 VTAIL.n22 B 0.008772f
C55 VTAIL.n23 B 0.015858f
C56 VTAIL.n24 B 0.009023f
C57 VTAIL.n25 B 0.020141f
C58 VTAIL.n26 B 0.009023f
C59 VTAIL.n27 B 0.015858f
C60 VTAIL.n28 B 0.008521f
C61 VTAIL.n29 B 0.020141f
C62 VTAIL.n30 B 0.009023f
C63 VTAIL.n31 B 1.27822f
C64 VTAIL.n32 B 0.008521f
C65 VTAIL.t7 B 0.034597f
C66 VTAIL.n33 B 0.155611f
C67 VTAIL.n34 B 0.014238f
C68 VTAIL.n35 B 0.015106f
C69 VTAIL.n36 B 0.020141f
C70 VTAIL.n37 B 0.009023f
C71 VTAIL.n38 B 0.008521f
C72 VTAIL.n39 B 0.015858f
C73 VTAIL.n40 B 0.015858f
C74 VTAIL.n41 B 0.008521f
C75 VTAIL.n42 B 0.009023f
C76 VTAIL.n43 B 0.020141f
C77 VTAIL.n44 B 0.020141f
C78 VTAIL.n45 B 0.009023f
C79 VTAIL.n46 B 0.008521f
C80 VTAIL.n47 B 0.015858f
C81 VTAIL.n48 B 0.015858f
C82 VTAIL.n49 B 0.008521f
C83 VTAIL.n50 B 0.008521f
C84 VTAIL.n51 B 0.009023f
C85 VTAIL.n52 B 0.020141f
C86 VTAIL.n53 B 0.020141f
C87 VTAIL.n54 B 0.020141f
C88 VTAIL.n55 B 0.008772f
C89 VTAIL.n56 B 0.008521f
C90 VTAIL.n57 B 0.015858f
C91 VTAIL.n58 B 0.015858f
C92 VTAIL.n59 B 0.008521f
C93 VTAIL.n60 B 0.009023f
C94 VTAIL.n61 B 0.020141f
C95 VTAIL.n62 B 0.020141f
C96 VTAIL.n63 B 0.009023f
C97 VTAIL.n64 B 0.008521f
C98 VTAIL.n65 B 0.015858f
C99 VTAIL.n66 B 0.015858f
C100 VTAIL.n67 B 0.008521f
C101 VTAIL.n68 B 0.009023f
C102 VTAIL.n69 B 0.020141f
C103 VTAIL.n70 B 0.020141f
C104 VTAIL.n71 B 0.009023f
C105 VTAIL.n72 B 0.008521f
C106 VTAIL.n73 B 0.015858f
C107 VTAIL.n74 B 0.015858f
C108 VTAIL.n75 B 0.008521f
C109 VTAIL.n76 B 0.009023f
C110 VTAIL.n77 B 0.020141f
C111 VTAIL.n78 B 0.020141f
C112 VTAIL.n79 B 0.009023f
C113 VTAIL.n80 B 0.008521f
C114 VTAIL.n81 B 0.015858f
C115 VTAIL.n82 B 0.015858f
C116 VTAIL.n83 B 0.008521f
C117 VTAIL.n84 B 0.009023f
C118 VTAIL.n85 B 0.020141f
C119 VTAIL.n86 B 0.020141f
C120 VTAIL.n87 B 0.009023f
C121 VTAIL.n88 B 0.008521f
C122 VTAIL.n89 B 0.015858f
C123 VTAIL.n90 B 0.015858f
C124 VTAIL.n91 B 0.008521f
C125 VTAIL.n92 B 0.009023f
C126 VTAIL.n93 B 0.020141f
C127 VTAIL.n94 B 0.020141f
C128 VTAIL.n95 B 0.009023f
C129 VTAIL.n96 B 0.008521f
C130 VTAIL.n97 B 0.015858f
C131 VTAIL.n98 B 0.040554f
C132 VTAIL.n99 B 0.008521f
C133 VTAIL.n100 B 0.009023f
C134 VTAIL.n101 B 0.040954f
C135 VTAIL.n102 B 0.03436f
C136 VTAIL.n103 B 0.06473f
C137 VTAIL.n104 B 0.008933f
C138 VTAIL.n105 B 0.020141f
C139 VTAIL.n106 B 0.009023f
C140 VTAIL.n107 B 0.015858f
C141 VTAIL.n108 B 0.008521f
C142 VTAIL.n109 B 0.020141f
C143 VTAIL.n110 B 0.009023f
C144 VTAIL.n111 B 0.015858f
C145 VTAIL.n112 B 0.008521f
C146 VTAIL.n113 B 0.020141f
C147 VTAIL.n114 B 0.009023f
C148 VTAIL.n115 B 0.015858f
C149 VTAIL.n116 B 0.008521f
C150 VTAIL.n117 B 0.020141f
C151 VTAIL.n118 B 0.009023f
C152 VTAIL.n119 B 0.015858f
C153 VTAIL.n120 B 0.008521f
C154 VTAIL.n121 B 0.020141f
C155 VTAIL.n122 B 0.009023f
C156 VTAIL.n123 B 0.015858f
C157 VTAIL.n124 B 0.008521f
C158 VTAIL.n125 B 0.020141f
C159 VTAIL.n126 B 0.008772f
C160 VTAIL.n127 B 0.015858f
C161 VTAIL.n128 B 0.009023f
C162 VTAIL.n129 B 0.020141f
C163 VTAIL.n130 B 0.009023f
C164 VTAIL.n131 B 0.015858f
C165 VTAIL.n132 B 0.008521f
C166 VTAIL.n133 B 0.020141f
C167 VTAIL.n134 B 0.009023f
C168 VTAIL.n135 B 1.27822f
C169 VTAIL.n136 B 0.008521f
C170 VTAIL.t3 B 0.034597f
C171 VTAIL.n137 B 0.155611f
C172 VTAIL.n138 B 0.014238f
C173 VTAIL.n139 B 0.015106f
C174 VTAIL.n140 B 0.020141f
C175 VTAIL.n141 B 0.009023f
C176 VTAIL.n142 B 0.008521f
C177 VTAIL.n143 B 0.015858f
C178 VTAIL.n144 B 0.015858f
C179 VTAIL.n145 B 0.008521f
C180 VTAIL.n146 B 0.009023f
C181 VTAIL.n147 B 0.020141f
C182 VTAIL.n148 B 0.020141f
C183 VTAIL.n149 B 0.009023f
C184 VTAIL.n150 B 0.008521f
C185 VTAIL.n151 B 0.015858f
C186 VTAIL.n152 B 0.015858f
C187 VTAIL.n153 B 0.008521f
C188 VTAIL.n154 B 0.008521f
C189 VTAIL.n155 B 0.009023f
C190 VTAIL.n156 B 0.020141f
C191 VTAIL.n157 B 0.020141f
C192 VTAIL.n158 B 0.020141f
C193 VTAIL.n159 B 0.008772f
C194 VTAIL.n160 B 0.008521f
C195 VTAIL.n161 B 0.015858f
C196 VTAIL.n162 B 0.015858f
C197 VTAIL.n163 B 0.008521f
C198 VTAIL.n164 B 0.009023f
C199 VTAIL.n165 B 0.020141f
C200 VTAIL.n166 B 0.020141f
C201 VTAIL.n167 B 0.009023f
C202 VTAIL.n168 B 0.008521f
C203 VTAIL.n169 B 0.015858f
C204 VTAIL.n170 B 0.015858f
C205 VTAIL.n171 B 0.008521f
C206 VTAIL.n172 B 0.009023f
C207 VTAIL.n173 B 0.020141f
C208 VTAIL.n174 B 0.020141f
C209 VTAIL.n175 B 0.009023f
C210 VTAIL.n176 B 0.008521f
C211 VTAIL.n177 B 0.015858f
C212 VTAIL.n178 B 0.015858f
C213 VTAIL.n179 B 0.008521f
C214 VTAIL.n180 B 0.009023f
C215 VTAIL.n181 B 0.020141f
C216 VTAIL.n182 B 0.020141f
C217 VTAIL.n183 B 0.009023f
C218 VTAIL.n184 B 0.008521f
C219 VTAIL.n185 B 0.015858f
C220 VTAIL.n186 B 0.015858f
C221 VTAIL.n187 B 0.008521f
C222 VTAIL.n188 B 0.009023f
C223 VTAIL.n189 B 0.020141f
C224 VTAIL.n190 B 0.020141f
C225 VTAIL.n191 B 0.009023f
C226 VTAIL.n192 B 0.008521f
C227 VTAIL.n193 B 0.015858f
C228 VTAIL.n194 B 0.015858f
C229 VTAIL.n195 B 0.008521f
C230 VTAIL.n196 B 0.009023f
C231 VTAIL.n197 B 0.020141f
C232 VTAIL.n198 B 0.020141f
C233 VTAIL.n199 B 0.009023f
C234 VTAIL.n200 B 0.008521f
C235 VTAIL.n201 B 0.015858f
C236 VTAIL.n202 B 0.040554f
C237 VTAIL.n203 B 0.008521f
C238 VTAIL.n204 B 0.009023f
C239 VTAIL.n205 B 0.040954f
C240 VTAIL.n206 B 0.03436f
C241 VTAIL.n207 B 0.084002f
C242 VTAIL.n208 B 0.008933f
C243 VTAIL.n209 B 0.020141f
C244 VTAIL.n210 B 0.009023f
C245 VTAIL.n211 B 0.015858f
C246 VTAIL.n212 B 0.008521f
C247 VTAIL.n213 B 0.020141f
C248 VTAIL.n214 B 0.009023f
C249 VTAIL.n215 B 0.015858f
C250 VTAIL.n216 B 0.008521f
C251 VTAIL.n217 B 0.020141f
C252 VTAIL.n218 B 0.009023f
C253 VTAIL.n219 B 0.015858f
C254 VTAIL.n220 B 0.008521f
C255 VTAIL.n221 B 0.020141f
C256 VTAIL.n222 B 0.009023f
C257 VTAIL.n223 B 0.015858f
C258 VTAIL.n224 B 0.008521f
C259 VTAIL.n225 B 0.020141f
C260 VTAIL.n226 B 0.009023f
C261 VTAIL.n227 B 0.015858f
C262 VTAIL.n228 B 0.008521f
C263 VTAIL.n229 B 0.020141f
C264 VTAIL.n230 B 0.008772f
C265 VTAIL.n231 B 0.015858f
C266 VTAIL.n232 B 0.009023f
C267 VTAIL.n233 B 0.020141f
C268 VTAIL.n234 B 0.009023f
C269 VTAIL.n235 B 0.015858f
C270 VTAIL.n236 B 0.008521f
C271 VTAIL.n237 B 0.020141f
C272 VTAIL.n238 B 0.009023f
C273 VTAIL.n239 B 1.27822f
C274 VTAIL.n240 B 0.008521f
C275 VTAIL.t2 B 0.034597f
C276 VTAIL.n241 B 0.155611f
C277 VTAIL.n242 B 0.014238f
C278 VTAIL.n243 B 0.015106f
C279 VTAIL.n244 B 0.020141f
C280 VTAIL.n245 B 0.009023f
C281 VTAIL.n246 B 0.008521f
C282 VTAIL.n247 B 0.015858f
C283 VTAIL.n248 B 0.015858f
C284 VTAIL.n249 B 0.008521f
C285 VTAIL.n250 B 0.009023f
C286 VTAIL.n251 B 0.020141f
C287 VTAIL.n252 B 0.020141f
C288 VTAIL.n253 B 0.009023f
C289 VTAIL.n254 B 0.008521f
C290 VTAIL.n255 B 0.015858f
C291 VTAIL.n256 B 0.015858f
C292 VTAIL.n257 B 0.008521f
C293 VTAIL.n258 B 0.008521f
C294 VTAIL.n259 B 0.009023f
C295 VTAIL.n260 B 0.020141f
C296 VTAIL.n261 B 0.020141f
C297 VTAIL.n262 B 0.020141f
C298 VTAIL.n263 B 0.008772f
C299 VTAIL.n264 B 0.008521f
C300 VTAIL.n265 B 0.015858f
C301 VTAIL.n266 B 0.015858f
C302 VTAIL.n267 B 0.008521f
C303 VTAIL.n268 B 0.009023f
C304 VTAIL.n269 B 0.020141f
C305 VTAIL.n270 B 0.020141f
C306 VTAIL.n271 B 0.009023f
C307 VTAIL.n272 B 0.008521f
C308 VTAIL.n273 B 0.015858f
C309 VTAIL.n274 B 0.015858f
C310 VTAIL.n275 B 0.008521f
C311 VTAIL.n276 B 0.009023f
C312 VTAIL.n277 B 0.020141f
C313 VTAIL.n278 B 0.020141f
C314 VTAIL.n279 B 0.009023f
C315 VTAIL.n280 B 0.008521f
C316 VTAIL.n281 B 0.015858f
C317 VTAIL.n282 B 0.015858f
C318 VTAIL.n283 B 0.008521f
C319 VTAIL.n284 B 0.009023f
C320 VTAIL.n285 B 0.020141f
C321 VTAIL.n286 B 0.020141f
C322 VTAIL.n287 B 0.009023f
C323 VTAIL.n288 B 0.008521f
C324 VTAIL.n289 B 0.015858f
C325 VTAIL.n290 B 0.015858f
C326 VTAIL.n291 B 0.008521f
C327 VTAIL.n292 B 0.009023f
C328 VTAIL.n293 B 0.020141f
C329 VTAIL.n294 B 0.020141f
C330 VTAIL.n295 B 0.009023f
C331 VTAIL.n296 B 0.008521f
C332 VTAIL.n297 B 0.015858f
C333 VTAIL.n298 B 0.015858f
C334 VTAIL.n299 B 0.008521f
C335 VTAIL.n300 B 0.009023f
C336 VTAIL.n301 B 0.020141f
C337 VTAIL.n302 B 0.020141f
C338 VTAIL.n303 B 0.009023f
C339 VTAIL.n304 B 0.008521f
C340 VTAIL.n305 B 0.015858f
C341 VTAIL.n306 B 0.040554f
C342 VTAIL.n307 B 0.008521f
C343 VTAIL.n308 B 0.009023f
C344 VTAIL.n309 B 0.040954f
C345 VTAIL.n310 B 0.03436f
C346 VTAIL.n311 B 1.14715f
C347 VTAIL.n312 B 0.008933f
C348 VTAIL.n313 B 0.020141f
C349 VTAIL.n314 B 0.009023f
C350 VTAIL.n315 B 0.015858f
C351 VTAIL.n316 B 0.008521f
C352 VTAIL.n317 B 0.020141f
C353 VTAIL.n318 B 0.009023f
C354 VTAIL.n319 B 0.015858f
C355 VTAIL.n320 B 0.008521f
C356 VTAIL.n321 B 0.020141f
C357 VTAIL.n322 B 0.009023f
C358 VTAIL.n323 B 0.015858f
C359 VTAIL.n324 B 0.008521f
C360 VTAIL.n325 B 0.020141f
C361 VTAIL.n326 B 0.009023f
C362 VTAIL.n327 B 0.015858f
C363 VTAIL.n328 B 0.008521f
C364 VTAIL.n329 B 0.020141f
C365 VTAIL.n330 B 0.009023f
C366 VTAIL.n331 B 0.015858f
C367 VTAIL.n332 B 0.008521f
C368 VTAIL.n333 B 0.020141f
C369 VTAIL.n334 B 0.008772f
C370 VTAIL.n335 B 0.015858f
C371 VTAIL.n336 B 0.008772f
C372 VTAIL.n337 B 0.008521f
C373 VTAIL.n338 B 0.020141f
C374 VTAIL.n339 B 0.020141f
C375 VTAIL.n340 B 0.009023f
C376 VTAIL.n341 B 0.015858f
C377 VTAIL.n342 B 0.008521f
C378 VTAIL.n343 B 0.020141f
C379 VTAIL.n344 B 0.009023f
C380 VTAIL.n345 B 1.27822f
C381 VTAIL.n346 B 0.008521f
C382 VTAIL.t6 B 0.034597f
C383 VTAIL.n347 B 0.155611f
C384 VTAIL.n348 B 0.014238f
C385 VTAIL.n349 B 0.015106f
C386 VTAIL.n350 B 0.020141f
C387 VTAIL.n351 B 0.009023f
C388 VTAIL.n352 B 0.008521f
C389 VTAIL.n353 B 0.015858f
C390 VTAIL.n354 B 0.015858f
C391 VTAIL.n355 B 0.008521f
C392 VTAIL.n356 B 0.009023f
C393 VTAIL.n357 B 0.020141f
C394 VTAIL.n358 B 0.020141f
C395 VTAIL.n359 B 0.009023f
C396 VTAIL.n360 B 0.008521f
C397 VTAIL.n361 B 0.015858f
C398 VTAIL.n362 B 0.015858f
C399 VTAIL.n363 B 0.008521f
C400 VTAIL.n364 B 0.009023f
C401 VTAIL.n365 B 0.020141f
C402 VTAIL.n366 B 0.020141f
C403 VTAIL.n367 B 0.009023f
C404 VTAIL.n368 B 0.008521f
C405 VTAIL.n369 B 0.015858f
C406 VTAIL.n370 B 0.015858f
C407 VTAIL.n371 B 0.008521f
C408 VTAIL.n372 B 0.009023f
C409 VTAIL.n373 B 0.020141f
C410 VTAIL.n374 B 0.020141f
C411 VTAIL.n375 B 0.009023f
C412 VTAIL.n376 B 0.008521f
C413 VTAIL.n377 B 0.015858f
C414 VTAIL.n378 B 0.015858f
C415 VTAIL.n379 B 0.008521f
C416 VTAIL.n380 B 0.009023f
C417 VTAIL.n381 B 0.020141f
C418 VTAIL.n382 B 0.020141f
C419 VTAIL.n383 B 0.009023f
C420 VTAIL.n384 B 0.008521f
C421 VTAIL.n385 B 0.015858f
C422 VTAIL.n386 B 0.015858f
C423 VTAIL.n387 B 0.008521f
C424 VTAIL.n388 B 0.009023f
C425 VTAIL.n389 B 0.020141f
C426 VTAIL.n390 B 0.020141f
C427 VTAIL.n391 B 0.009023f
C428 VTAIL.n392 B 0.008521f
C429 VTAIL.n393 B 0.015858f
C430 VTAIL.n394 B 0.015858f
C431 VTAIL.n395 B 0.008521f
C432 VTAIL.n396 B 0.009023f
C433 VTAIL.n397 B 0.020141f
C434 VTAIL.n398 B 0.020141f
C435 VTAIL.n399 B 0.009023f
C436 VTAIL.n400 B 0.008521f
C437 VTAIL.n401 B 0.015858f
C438 VTAIL.n402 B 0.015858f
C439 VTAIL.n403 B 0.008521f
C440 VTAIL.n404 B 0.009023f
C441 VTAIL.n405 B 0.020141f
C442 VTAIL.n406 B 0.020141f
C443 VTAIL.n407 B 0.009023f
C444 VTAIL.n408 B 0.008521f
C445 VTAIL.n409 B 0.015858f
C446 VTAIL.n410 B 0.040554f
C447 VTAIL.n411 B 0.008521f
C448 VTAIL.n412 B 0.009023f
C449 VTAIL.n413 B 0.040954f
C450 VTAIL.n414 B 0.03436f
C451 VTAIL.n415 B 1.14715f
C452 VTAIL.n416 B 0.008933f
C453 VTAIL.n417 B 0.020141f
C454 VTAIL.n418 B 0.009023f
C455 VTAIL.n419 B 0.015858f
C456 VTAIL.n420 B 0.008521f
C457 VTAIL.n421 B 0.020141f
C458 VTAIL.n422 B 0.009023f
C459 VTAIL.n423 B 0.015858f
C460 VTAIL.n424 B 0.008521f
C461 VTAIL.n425 B 0.020141f
C462 VTAIL.n426 B 0.009023f
C463 VTAIL.n427 B 0.015858f
C464 VTAIL.n428 B 0.008521f
C465 VTAIL.n429 B 0.020141f
C466 VTAIL.n430 B 0.009023f
C467 VTAIL.n431 B 0.015858f
C468 VTAIL.n432 B 0.008521f
C469 VTAIL.n433 B 0.020141f
C470 VTAIL.n434 B 0.009023f
C471 VTAIL.n435 B 0.015858f
C472 VTAIL.n436 B 0.008521f
C473 VTAIL.n437 B 0.020141f
C474 VTAIL.n438 B 0.008772f
C475 VTAIL.n439 B 0.015858f
C476 VTAIL.n440 B 0.008772f
C477 VTAIL.n441 B 0.008521f
C478 VTAIL.n442 B 0.020141f
C479 VTAIL.n443 B 0.020141f
C480 VTAIL.n444 B 0.009023f
C481 VTAIL.n445 B 0.015858f
C482 VTAIL.n446 B 0.008521f
C483 VTAIL.n447 B 0.020141f
C484 VTAIL.n448 B 0.009023f
C485 VTAIL.n449 B 1.27822f
C486 VTAIL.n450 B 0.008521f
C487 VTAIL.t4 B 0.034597f
C488 VTAIL.n451 B 0.155611f
C489 VTAIL.n452 B 0.014238f
C490 VTAIL.n453 B 0.015106f
C491 VTAIL.n454 B 0.020141f
C492 VTAIL.n455 B 0.009023f
C493 VTAIL.n456 B 0.008521f
C494 VTAIL.n457 B 0.015858f
C495 VTAIL.n458 B 0.015858f
C496 VTAIL.n459 B 0.008521f
C497 VTAIL.n460 B 0.009023f
C498 VTAIL.n461 B 0.020141f
C499 VTAIL.n462 B 0.020141f
C500 VTAIL.n463 B 0.009023f
C501 VTAIL.n464 B 0.008521f
C502 VTAIL.n465 B 0.015858f
C503 VTAIL.n466 B 0.015858f
C504 VTAIL.n467 B 0.008521f
C505 VTAIL.n468 B 0.009023f
C506 VTAIL.n469 B 0.020141f
C507 VTAIL.n470 B 0.020141f
C508 VTAIL.n471 B 0.009023f
C509 VTAIL.n472 B 0.008521f
C510 VTAIL.n473 B 0.015858f
C511 VTAIL.n474 B 0.015858f
C512 VTAIL.n475 B 0.008521f
C513 VTAIL.n476 B 0.009023f
C514 VTAIL.n477 B 0.020141f
C515 VTAIL.n478 B 0.020141f
C516 VTAIL.n479 B 0.009023f
C517 VTAIL.n480 B 0.008521f
C518 VTAIL.n481 B 0.015858f
C519 VTAIL.n482 B 0.015858f
C520 VTAIL.n483 B 0.008521f
C521 VTAIL.n484 B 0.009023f
C522 VTAIL.n485 B 0.020141f
C523 VTAIL.n486 B 0.020141f
C524 VTAIL.n487 B 0.009023f
C525 VTAIL.n488 B 0.008521f
C526 VTAIL.n489 B 0.015858f
C527 VTAIL.n490 B 0.015858f
C528 VTAIL.n491 B 0.008521f
C529 VTAIL.n492 B 0.009023f
C530 VTAIL.n493 B 0.020141f
C531 VTAIL.n494 B 0.020141f
C532 VTAIL.n495 B 0.009023f
C533 VTAIL.n496 B 0.008521f
C534 VTAIL.n497 B 0.015858f
C535 VTAIL.n498 B 0.015858f
C536 VTAIL.n499 B 0.008521f
C537 VTAIL.n500 B 0.009023f
C538 VTAIL.n501 B 0.020141f
C539 VTAIL.n502 B 0.020141f
C540 VTAIL.n503 B 0.009023f
C541 VTAIL.n504 B 0.008521f
C542 VTAIL.n505 B 0.015858f
C543 VTAIL.n506 B 0.015858f
C544 VTAIL.n507 B 0.008521f
C545 VTAIL.n508 B 0.009023f
C546 VTAIL.n509 B 0.020141f
C547 VTAIL.n510 B 0.020141f
C548 VTAIL.n511 B 0.009023f
C549 VTAIL.n512 B 0.008521f
C550 VTAIL.n513 B 0.015858f
C551 VTAIL.n514 B 0.040554f
C552 VTAIL.n515 B 0.008521f
C553 VTAIL.n516 B 0.009023f
C554 VTAIL.n517 B 0.040954f
C555 VTAIL.n518 B 0.03436f
C556 VTAIL.n519 B 0.084002f
C557 VTAIL.n520 B 0.008933f
C558 VTAIL.n521 B 0.020141f
C559 VTAIL.n522 B 0.009023f
C560 VTAIL.n523 B 0.015858f
C561 VTAIL.n524 B 0.008521f
C562 VTAIL.n525 B 0.020141f
C563 VTAIL.n526 B 0.009023f
C564 VTAIL.n527 B 0.015858f
C565 VTAIL.n528 B 0.008521f
C566 VTAIL.n529 B 0.020141f
C567 VTAIL.n530 B 0.009023f
C568 VTAIL.n531 B 0.015858f
C569 VTAIL.n532 B 0.008521f
C570 VTAIL.n533 B 0.020141f
C571 VTAIL.n534 B 0.009023f
C572 VTAIL.n535 B 0.015858f
C573 VTAIL.n536 B 0.008521f
C574 VTAIL.n537 B 0.020141f
C575 VTAIL.n538 B 0.009023f
C576 VTAIL.n539 B 0.015858f
C577 VTAIL.n540 B 0.008521f
C578 VTAIL.n541 B 0.020141f
C579 VTAIL.n542 B 0.008772f
C580 VTAIL.n543 B 0.015858f
C581 VTAIL.n544 B 0.008772f
C582 VTAIL.n545 B 0.008521f
C583 VTAIL.n546 B 0.020141f
C584 VTAIL.n547 B 0.020141f
C585 VTAIL.n548 B 0.009023f
C586 VTAIL.n549 B 0.015858f
C587 VTAIL.n550 B 0.008521f
C588 VTAIL.n551 B 0.020141f
C589 VTAIL.n552 B 0.009023f
C590 VTAIL.n553 B 1.27822f
C591 VTAIL.n554 B 0.008521f
C592 VTAIL.t1 B 0.034597f
C593 VTAIL.n555 B 0.155611f
C594 VTAIL.n556 B 0.014238f
C595 VTAIL.n557 B 0.015106f
C596 VTAIL.n558 B 0.020141f
C597 VTAIL.n559 B 0.009023f
C598 VTAIL.n560 B 0.008521f
C599 VTAIL.n561 B 0.015858f
C600 VTAIL.n562 B 0.015858f
C601 VTAIL.n563 B 0.008521f
C602 VTAIL.n564 B 0.009023f
C603 VTAIL.n565 B 0.020141f
C604 VTAIL.n566 B 0.020141f
C605 VTAIL.n567 B 0.009023f
C606 VTAIL.n568 B 0.008521f
C607 VTAIL.n569 B 0.015858f
C608 VTAIL.n570 B 0.015858f
C609 VTAIL.n571 B 0.008521f
C610 VTAIL.n572 B 0.009023f
C611 VTAIL.n573 B 0.020141f
C612 VTAIL.n574 B 0.020141f
C613 VTAIL.n575 B 0.009023f
C614 VTAIL.n576 B 0.008521f
C615 VTAIL.n577 B 0.015858f
C616 VTAIL.n578 B 0.015858f
C617 VTAIL.n579 B 0.008521f
C618 VTAIL.n580 B 0.009023f
C619 VTAIL.n581 B 0.020141f
C620 VTAIL.n582 B 0.020141f
C621 VTAIL.n583 B 0.009023f
C622 VTAIL.n584 B 0.008521f
C623 VTAIL.n585 B 0.015858f
C624 VTAIL.n586 B 0.015858f
C625 VTAIL.n587 B 0.008521f
C626 VTAIL.n588 B 0.009023f
C627 VTAIL.n589 B 0.020141f
C628 VTAIL.n590 B 0.020141f
C629 VTAIL.n591 B 0.009023f
C630 VTAIL.n592 B 0.008521f
C631 VTAIL.n593 B 0.015858f
C632 VTAIL.n594 B 0.015858f
C633 VTAIL.n595 B 0.008521f
C634 VTAIL.n596 B 0.009023f
C635 VTAIL.n597 B 0.020141f
C636 VTAIL.n598 B 0.020141f
C637 VTAIL.n599 B 0.009023f
C638 VTAIL.n600 B 0.008521f
C639 VTAIL.n601 B 0.015858f
C640 VTAIL.n602 B 0.015858f
C641 VTAIL.n603 B 0.008521f
C642 VTAIL.n604 B 0.009023f
C643 VTAIL.n605 B 0.020141f
C644 VTAIL.n606 B 0.020141f
C645 VTAIL.n607 B 0.009023f
C646 VTAIL.n608 B 0.008521f
C647 VTAIL.n609 B 0.015858f
C648 VTAIL.n610 B 0.015858f
C649 VTAIL.n611 B 0.008521f
C650 VTAIL.n612 B 0.009023f
C651 VTAIL.n613 B 0.020141f
C652 VTAIL.n614 B 0.020141f
C653 VTAIL.n615 B 0.009023f
C654 VTAIL.n616 B 0.008521f
C655 VTAIL.n617 B 0.015858f
C656 VTAIL.n618 B 0.040554f
C657 VTAIL.n619 B 0.008521f
C658 VTAIL.n620 B 0.009023f
C659 VTAIL.n621 B 0.040954f
C660 VTAIL.n622 B 0.03436f
C661 VTAIL.n623 B 0.084002f
C662 VTAIL.n624 B 0.008933f
C663 VTAIL.n625 B 0.020141f
C664 VTAIL.n626 B 0.009023f
C665 VTAIL.n627 B 0.015858f
C666 VTAIL.n628 B 0.008521f
C667 VTAIL.n629 B 0.020141f
C668 VTAIL.n630 B 0.009023f
C669 VTAIL.n631 B 0.015858f
C670 VTAIL.n632 B 0.008521f
C671 VTAIL.n633 B 0.020141f
C672 VTAIL.n634 B 0.009023f
C673 VTAIL.n635 B 0.015858f
C674 VTAIL.n636 B 0.008521f
C675 VTAIL.n637 B 0.020141f
C676 VTAIL.n638 B 0.009023f
C677 VTAIL.n639 B 0.015858f
C678 VTAIL.n640 B 0.008521f
C679 VTAIL.n641 B 0.020141f
C680 VTAIL.n642 B 0.009023f
C681 VTAIL.n643 B 0.015858f
C682 VTAIL.n644 B 0.008521f
C683 VTAIL.n645 B 0.020141f
C684 VTAIL.n646 B 0.008772f
C685 VTAIL.n647 B 0.015858f
C686 VTAIL.n648 B 0.008772f
C687 VTAIL.n649 B 0.008521f
C688 VTAIL.n650 B 0.020141f
C689 VTAIL.n651 B 0.020141f
C690 VTAIL.n652 B 0.009023f
C691 VTAIL.n653 B 0.015858f
C692 VTAIL.n654 B 0.008521f
C693 VTAIL.n655 B 0.020141f
C694 VTAIL.n656 B 0.009023f
C695 VTAIL.n657 B 1.27822f
C696 VTAIL.n658 B 0.008521f
C697 VTAIL.t0 B 0.034597f
C698 VTAIL.n659 B 0.155611f
C699 VTAIL.n660 B 0.014238f
C700 VTAIL.n661 B 0.015106f
C701 VTAIL.n662 B 0.020141f
C702 VTAIL.n663 B 0.009023f
C703 VTAIL.n664 B 0.008521f
C704 VTAIL.n665 B 0.015858f
C705 VTAIL.n666 B 0.015858f
C706 VTAIL.n667 B 0.008521f
C707 VTAIL.n668 B 0.009023f
C708 VTAIL.n669 B 0.020141f
C709 VTAIL.n670 B 0.020141f
C710 VTAIL.n671 B 0.009023f
C711 VTAIL.n672 B 0.008521f
C712 VTAIL.n673 B 0.015858f
C713 VTAIL.n674 B 0.015858f
C714 VTAIL.n675 B 0.008521f
C715 VTAIL.n676 B 0.009023f
C716 VTAIL.n677 B 0.020141f
C717 VTAIL.n678 B 0.020141f
C718 VTAIL.n679 B 0.009023f
C719 VTAIL.n680 B 0.008521f
C720 VTAIL.n681 B 0.015858f
C721 VTAIL.n682 B 0.015858f
C722 VTAIL.n683 B 0.008521f
C723 VTAIL.n684 B 0.009023f
C724 VTAIL.n685 B 0.020141f
C725 VTAIL.n686 B 0.020141f
C726 VTAIL.n687 B 0.009023f
C727 VTAIL.n688 B 0.008521f
C728 VTAIL.n689 B 0.015858f
C729 VTAIL.n690 B 0.015858f
C730 VTAIL.n691 B 0.008521f
C731 VTAIL.n692 B 0.009023f
C732 VTAIL.n693 B 0.020141f
C733 VTAIL.n694 B 0.020141f
C734 VTAIL.n695 B 0.009023f
C735 VTAIL.n696 B 0.008521f
C736 VTAIL.n697 B 0.015858f
C737 VTAIL.n698 B 0.015858f
C738 VTAIL.n699 B 0.008521f
C739 VTAIL.n700 B 0.009023f
C740 VTAIL.n701 B 0.020141f
C741 VTAIL.n702 B 0.020141f
C742 VTAIL.n703 B 0.009023f
C743 VTAIL.n704 B 0.008521f
C744 VTAIL.n705 B 0.015858f
C745 VTAIL.n706 B 0.015858f
C746 VTAIL.n707 B 0.008521f
C747 VTAIL.n708 B 0.009023f
C748 VTAIL.n709 B 0.020141f
C749 VTAIL.n710 B 0.020141f
C750 VTAIL.n711 B 0.009023f
C751 VTAIL.n712 B 0.008521f
C752 VTAIL.n713 B 0.015858f
C753 VTAIL.n714 B 0.015858f
C754 VTAIL.n715 B 0.008521f
C755 VTAIL.n716 B 0.009023f
C756 VTAIL.n717 B 0.020141f
C757 VTAIL.n718 B 0.020141f
C758 VTAIL.n719 B 0.009023f
C759 VTAIL.n720 B 0.008521f
C760 VTAIL.n721 B 0.015858f
C761 VTAIL.n722 B 0.040554f
C762 VTAIL.n723 B 0.008521f
C763 VTAIL.n724 B 0.009023f
C764 VTAIL.n725 B 0.040954f
C765 VTAIL.n726 B 0.03436f
C766 VTAIL.n727 B 1.14715f
C767 VTAIL.n728 B 0.008933f
C768 VTAIL.n729 B 0.020141f
C769 VTAIL.n730 B 0.009023f
C770 VTAIL.n731 B 0.015858f
C771 VTAIL.n732 B 0.008521f
C772 VTAIL.n733 B 0.020141f
C773 VTAIL.n734 B 0.009023f
C774 VTAIL.n735 B 0.015858f
C775 VTAIL.n736 B 0.008521f
C776 VTAIL.n737 B 0.020141f
C777 VTAIL.n738 B 0.009023f
C778 VTAIL.n739 B 0.015858f
C779 VTAIL.n740 B 0.008521f
C780 VTAIL.n741 B 0.020141f
C781 VTAIL.n742 B 0.009023f
C782 VTAIL.n743 B 0.015858f
C783 VTAIL.n744 B 0.008521f
C784 VTAIL.n745 B 0.020141f
C785 VTAIL.n746 B 0.009023f
C786 VTAIL.n747 B 0.015858f
C787 VTAIL.n748 B 0.008521f
C788 VTAIL.n749 B 0.020141f
C789 VTAIL.n750 B 0.008772f
C790 VTAIL.n751 B 0.015858f
C791 VTAIL.n752 B 0.009023f
C792 VTAIL.n753 B 0.020141f
C793 VTAIL.n754 B 0.009023f
C794 VTAIL.n755 B 0.015858f
C795 VTAIL.n756 B 0.008521f
C796 VTAIL.n757 B 0.020141f
C797 VTAIL.n758 B 0.009023f
C798 VTAIL.n759 B 1.27822f
C799 VTAIL.n760 B 0.008521f
C800 VTAIL.t5 B 0.034597f
C801 VTAIL.n761 B 0.155611f
C802 VTAIL.n762 B 0.014238f
C803 VTAIL.n763 B 0.015106f
C804 VTAIL.n764 B 0.020141f
C805 VTAIL.n765 B 0.009023f
C806 VTAIL.n766 B 0.008521f
C807 VTAIL.n767 B 0.015858f
C808 VTAIL.n768 B 0.015858f
C809 VTAIL.n769 B 0.008521f
C810 VTAIL.n770 B 0.009023f
C811 VTAIL.n771 B 0.020141f
C812 VTAIL.n772 B 0.020141f
C813 VTAIL.n773 B 0.009023f
C814 VTAIL.n774 B 0.008521f
C815 VTAIL.n775 B 0.015858f
C816 VTAIL.n776 B 0.015858f
C817 VTAIL.n777 B 0.008521f
C818 VTAIL.n778 B 0.008521f
C819 VTAIL.n779 B 0.009023f
C820 VTAIL.n780 B 0.020141f
C821 VTAIL.n781 B 0.020141f
C822 VTAIL.n782 B 0.020141f
C823 VTAIL.n783 B 0.008772f
C824 VTAIL.n784 B 0.008521f
C825 VTAIL.n785 B 0.015858f
C826 VTAIL.n786 B 0.015858f
C827 VTAIL.n787 B 0.008521f
C828 VTAIL.n788 B 0.009023f
C829 VTAIL.n789 B 0.020141f
C830 VTAIL.n790 B 0.020141f
C831 VTAIL.n791 B 0.009023f
C832 VTAIL.n792 B 0.008521f
C833 VTAIL.n793 B 0.015858f
C834 VTAIL.n794 B 0.015858f
C835 VTAIL.n795 B 0.008521f
C836 VTAIL.n796 B 0.009023f
C837 VTAIL.n797 B 0.020141f
C838 VTAIL.n798 B 0.020141f
C839 VTAIL.n799 B 0.009023f
C840 VTAIL.n800 B 0.008521f
C841 VTAIL.n801 B 0.015858f
C842 VTAIL.n802 B 0.015858f
C843 VTAIL.n803 B 0.008521f
C844 VTAIL.n804 B 0.009023f
C845 VTAIL.n805 B 0.020141f
C846 VTAIL.n806 B 0.020141f
C847 VTAIL.n807 B 0.009023f
C848 VTAIL.n808 B 0.008521f
C849 VTAIL.n809 B 0.015858f
C850 VTAIL.n810 B 0.015858f
C851 VTAIL.n811 B 0.008521f
C852 VTAIL.n812 B 0.009023f
C853 VTAIL.n813 B 0.020141f
C854 VTAIL.n814 B 0.020141f
C855 VTAIL.n815 B 0.009023f
C856 VTAIL.n816 B 0.008521f
C857 VTAIL.n817 B 0.015858f
C858 VTAIL.n818 B 0.015858f
C859 VTAIL.n819 B 0.008521f
C860 VTAIL.n820 B 0.009023f
C861 VTAIL.n821 B 0.020141f
C862 VTAIL.n822 B 0.020141f
C863 VTAIL.n823 B 0.009023f
C864 VTAIL.n824 B 0.008521f
C865 VTAIL.n825 B 0.015858f
C866 VTAIL.n826 B 0.040554f
C867 VTAIL.n827 B 0.008521f
C868 VTAIL.n828 B 0.009023f
C869 VTAIL.n829 B 0.040954f
C870 VTAIL.n830 B 0.03436f
C871 VTAIL.n831 B 1.12193f
C872 VDD2.t0 B 0.423695f
C873 VDD2.t2 B 0.423695f
C874 VDD2.n0 B 4.72586f
C875 VDD2.t1 B 0.423695f
C876 VDD2.t3 B 0.423695f
C877 VDD2.n1 B 3.87671f
C878 VDD2.n2 B 4.31641f
C879 VN.t0 B 1.80668f
C880 VN.t2 B 1.80664f
C881 VN.n0 B 1.30944f
C882 VN.t3 B 1.80668f
C883 VN.t1 B 1.80664f
C884 VN.n1 B 2.55315f
.ends

