* NGSPICE file created from diff_pair_sample_0835.ext - technology: sky130A

.subckt diff_pair_sample_0835 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=3.88
X1 VTAIL.t7 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=3.88
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=3.88
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=3.88
X4 VTAIL.t6 VN.t1 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=3.88
X5 VDD2.t2 VN.t2 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=3.88
X6 VDD1.t3 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=3.88
X7 VDD2.t1 VN.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=3.88
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0 ps=0 w=2.01 l=3.88
X9 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.33165 pd=2.34 as=0.7839 ps=4.8 w=2.01 l=3.88
X10 VTAIL.t3 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=3.88
X11 VTAIL.t0 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7839 pd=4.8 as=0.33165 ps=2.34 w=2.01 l=3.88
R0 B.n543 B.n542 585
R1 B.n171 B.n100 585
R2 B.n170 B.n169 585
R3 B.n168 B.n167 585
R4 B.n166 B.n165 585
R5 B.n164 B.n163 585
R6 B.n162 B.n161 585
R7 B.n160 B.n159 585
R8 B.n158 B.n157 585
R9 B.n156 B.n155 585
R10 B.n154 B.n153 585
R11 B.n152 B.n151 585
R12 B.n150 B.n149 585
R13 B.n148 B.n147 585
R14 B.n146 B.n145 585
R15 B.n144 B.n143 585
R16 B.n142 B.n141 585
R17 B.n140 B.n139 585
R18 B.n138 B.n137 585
R19 B.n136 B.n135 585
R20 B.n134 B.n133 585
R21 B.n132 B.n131 585
R22 B.n130 B.n129 585
R23 B.n128 B.n127 585
R24 B.n126 B.n125 585
R25 B.n124 B.n123 585
R26 B.n122 B.n121 585
R27 B.n120 B.n119 585
R28 B.n118 B.n117 585
R29 B.n116 B.n115 585
R30 B.n114 B.n113 585
R31 B.n112 B.n111 585
R32 B.n110 B.n109 585
R33 B.n108 B.n107 585
R34 B.n541 B.n83 585
R35 B.n546 B.n83 585
R36 B.n540 B.n82 585
R37 B.n547 B.n82 585
R38 B.n539 B.n538 585
R39 B.n538 B.n78 585
R40 B.n537 B.n77 585
R41 B.n553 B.n77 585
R42 B.n536 B.n76 585
R43 B.n554 B.n76 585
R44 B.n535 B.n75 585
R45 B.n555 B.n75 585
R46 B.n534 B.n533 585
R47 B.n533 B.n71 585
R48 B.n532 B.n70 585
R49 B.n561 B.n70 585
R50 B.n531 B.n69 585
R51 B.n562 B.n69 585
R52 B.n530 B.n68 585
R53 B.n563 B.n68 585
R54 B.n529 B.n528 585
R55 B.n528 B.n64 585
R56 B.n527 B.n63 585
R57 B.n569 B.n63 585
R58 B.n526 B.n62 585
R59 B.n570 B.n62 585
R60 B.n525 B.n61 585
R61 B.n571 B.n61 585
R62 B.n524 B.n523 585
R63 B.n523 B.n57 585
R64 B.n522 B.n56 585
R65 B.n577 B.n56 585
R66 B.n521 B.n55 585
R67 B.n578 B.n55 585
R68 B.n520 B.n54 585
R69 B.n579 B.n54 585
R70 B.n519 B.n518 585
R71 B.n518 B.n50 585
R72 B.n517 B.n49 585
R73 B.n585 B.n49 585
R74 B.n516 B.n48 585
R75 B.n586 B.n48 585
R76 B.n515 B.n47 585
R77 B.n587 B.n47 585
R78 B.n514 B.n513 585
R79 B.n513 B.n43 585
R80 B.n512 B.n42 585
R81 B.n593 B.n42 585
R82 B.n511 B.n41 585
R83 B.n594 B.n41 585
R84 B.n510 B.n40 585
R85 B.n595 B.n40 585
R86 B.n509 B.n508 585
R87 B.n508 B.n36 585
R88 B.n507 B.n35 585
R89 B.n601 B.n35 585
R90 B.n506 B.n34 585
R91 B.n602 B.n34 585
R92 B.n505 B.n33 585
R93 B.n603 B.n33 585
R94 B.n504 B.n503 585
R95 B.n503 B.n29 585
R96 B.n502 B.n28 585
R97 B.n609 B.n28 585
R98 B.n501 B.n27 585
R99 B.n610 B.n27 585
R100 B.n500 B.n26 585
R101 B.n611 B.n26 585
R102 B.n499 B.n498 585
R103 B.n498 B.n22 585
R104 B.n497 B.n21 585
R105 B.n617 B.n21 585
R106 B.n496 B.n20 585
R107 B.n618 B.n20 585
R108 B.n495 B.n19 585
R109 B.n619 B.n19 585
R110 B.n494 B.n493 585
R111 B.n493 B.n15 585
R112 B.n492 B.n14 585
R113 B.n625 B.n14 585
R114 B.n491 B.n13 585
R115 B.n626 B.n13 585
R116 B.n490 B.n12 585
R117 B.n627 B.n12 585
R118 B.n489 B.n488 585
R119 B.n488 B.n8 585
R120 B.n487 B.n7 585
R121 B.n633 B.n7 585
R122 B.n486 B.n6 585
R123 B.n634 B.n6 585
R124 B.n485 B.n5 585
R125 B.n635 B.n5 585
R126 B.n484 B.n483 585
R127 B.n483 B.n4 585
R128 B.n482 B.n172 585
R129 B.n482 B.n481 585
R130 B.n472 B.n173 585
R131 B.n174 B.n173 585
R132 B.n474 B.n473 585
R133 B.n475 B.n474 585
R134 B.n471 B.n179 585
R135 B.n179 B.n178 585
R136 B.n470 B.n469 585
R137 B.n469 B.n468 585
R138 B.n181 B.n180 585
R139 B.n182 B.n181 585
R140 B.n461 B.n460 585
R141 B.n462 B.n461 585
R142 B.n459 B.n187 585
R143 B.n187 B.n186 585
R144 B.n458 B.n457 585
R145 B.n457 B.n456 585
R146 B.n189 B.n188 585
R147 B.n190 B.n189 585
R148 B.n449 B.n448 585
R149 B.n450 B.n449 585
R150 B.n447 B.n195 585
R151 B.n195 B.n194 585
R152 B.n446 B.n445 585
R153 B.n445 B.n444 585
R154 B.n197 B.n196 585
R155 B.n198 B.n197 585
R156 B.n437 B.n436 585
R157 B.n438 B.n437 585
R158 B.n435 B.n203 585
R159 B.n203 B.n202 585
R160 B.n434 B.n433 585
R161 B.n433 B.n432 585
R162 B.n205 B.n204 585
R163 B.n206 B.n205 585
R164 B.n425 B.n424 585
R165 B.n426 B.n425 585
R166 B.n423 B.n210 585
R167 B.n214 B.n210 585
R168 B.n422 B.n421 585
R169 B.n421 B.n420 585
R170 B.n212 B.n211 585
R171 B.n213 B.n212 585
R172 B.n413 B.n412 585
R173 B.n414 B.n413 585
R174 B.n411 B.n219 585
R175 B.n219 B.n218 585
R176 B.n410 B.n409 585
R177 B.n409 B.n408 585
R178 B.n221 B.n220 585
R179 B.n222 B.n221 585
R180 B.n401 B.n400 585
R181 B.n402 B.n401 585
R182 B.n399 B.n227 585
R183 B.n227 B.n226 585
R184 B.n398 B.n397 585
R185 B.n397 B.n396 585
R186 B.n229 B.n228 585
R187 B.n230 B.n229 585
R188 B.n389 B.n388 585
R189 B.n390 B.n389 585
R190 B.n387 B.n235 585
R191 B.n235 B.n234 585
R192 B.n386 B.n385 585
R193 B.n385 B.n384 585
R194 B.n237 B.n236 585
R195 B.n238 B.n237 585
R196 B.n377 B.n376 585
R197 B.n378 B.n377 585
R198 B.n375 B.n243 585
R199 B.n243 B.n242 585
R200 B.n374 B.n373 585
R201 B.n373 B.n372 585
R202 B.n245 B.n244 585
R203 B.n246 B.n245 585
R204 B.n365 B.n364 585
R205 B.n366 B.n365 585
R206 B.n363 B.n251 585
R207 B.n251 B.n250 585
R208 B.n362 B.n361 585
R209 B.n361 B.n360 585
R210 B.n253 B.n252 585
R211 B.n254 B.n253 585
R212 B.n353 B.n352 585
R213 B.n354 B.n353 585
R214 B.n351 B.n259 585
R215 B.n259 B.n258 585
R216 B.n346 B.n345 585
R217 B.n344 B.n278 585
R218 B.n343 B.n277 585
R219 B.n348 B.n277 585
R220 B.n342 B.n341 585
R221 B.n340 B.n339 585
R222 B.n338 B.n337 585
R223 B.n336 B.n335 585
R224 B.n334 B.n333 585
R225 B.n332 B.n331 585
R226 B.n330 B.n329 585
R227 B.n328 B.n327 585
R228 B.n326 B.n325 585
R229 B.n323 B.n322 585
R230 B.n321 B.n320 585
R231 B.n319 B.n318 585
R232 B.n317 B.n316 585
R233 B.n315 B.n314 585
R234 B.n313 B.n312 585
R235 B.n311 B.n310 585
R236 B.n309 B.n308 585
R237 B.n307 B.n306 585
R238 B.n305 B.n304 585
R239 B.n302 B.n301 585
R240 B.n300 B.n299 585
R241 B.n298 B.n297 585
R242 B.n296 B.n295 585
R243 B.n294 B.n293 585
R244 B.n292 B.n291 585
R245 B.n290 B.n289 585
R246 B.n288 B.n287 585
R247 B.n286 B.n285 585
R248 B.n284 B.n283 585
R249 B.n261 B.n260 585
R250 B.n350 B.n349 585
R251 B.n349 B.n348 585
R252 B.n257 B.n256 585
R253 B.n258 B.n257 585
R254 B.n356 B.n355 585
R255 B.n355 B.n354 585
R256 B.n357 B.n255 585
R257 B.n255 B.n254 585
R258 B.n359 B.n358 585
R259 B.n360 B.n359 585
R260 B.n249 B.n248 585
R261 B.n250 B.n249 585
R262 B.n368 B.n367 585
R263 B.n367 B.n366 585
R264 B.n369 B.n247 585
R265 B.n247 B.n246 585
R266 B.n371 B.n370 585
R267 B.n372 B.n371 585
R268 B.n241 B.n240 585
R269 B.n242 B.n241 585
R270 B.n380 B.n379 585
R271 B.n379 B.n378 585
R272 B.n381 B.n239 585
R273 B.n239 B.n238 585
R274 B.n383 B.n382 585
R275 B.n384 B.n383 585
R276 B.n233 B.n232 585
R277 B.n234 B.n233 585
R278 B.n392 B.n391 585
R279 B.n391 B.n390 585
R280 B.n393 B.n231 585
R281 B.n231 B.n230 585
R282 B.n395 B.n394 585
R283 B.n396 B.n395 585
R284 B.n225 B.n224 585
R285 B.n226 B.n225 585
R286 B.n404 B.n403 585
R287 B.n403 B.n402 585
R288 B.n405 B.n223 585
R289 B.n223 B.n222 585
R290 B.n407 B.n406 585
R291 B.n408 B.n407 585
R292 B.n217 B.n216 585
R293 B.n218 B.n217 585
R294 B.n416 B.n415 585
R295 B.n415 B.n414 585
R296 B.n417 B.n215 585
R297 B.n215 B.n213 585
R298 B.n419 B.n418 585
R299 B.n420 B.n419 585
R300 B.n209 B.n208 585
R301 B.n214 B.n209 585
R302 B.n428 B.n427 585
R303 B.n427 B.n426 585
R304 B.n429 B.n207 585
R305 B.n207 B.n206 585
R306 B.n431 B.n430 585
R307 B.n432 B.n431 585
R308 B.n201 B.n200 585
R309 B.n202 B.n201 585
R310 B.n440 B.n439 585
R311 B.n439 B.n438 585
R312 B.n441 B.n199 585
R313 B.n199 B.n198 585
R314 B.n443 B.n442 585
R315 B.n444 B.n443 585
R316 B.n193 B.n192 585
R317 B.n194 B.n193 585
R318 B.n452 B.n451 585
R319 B.n451 B.n450 585
R320 B.n453 B.n191 585
R321 B.n191 B.n190 585
R322 B.n455 B.n454 585
R323 B.n456 B.n455 585
R324 B.n185 B.n184 585
R325 B.n186 B.n185 585
R326 B.n464 B.n463 585
R327 B.n463 B.n462 585
R328 B.n465 B.n183 585
R329 B.n183 B.n182 585
R330 B.n467 B.n466 585
R331 B.n468 B.n467 585
R332 B.n177 B.n176 585
R333 B.n178 B.n177 585
R334 B.n477 B.n476 585
R335 B.n476 B.n475 585
R336 B.n478 B.n175 585
R337 B.n175 B.n174 585
R338 B.n480 B.n479 585
R339 B.n481 B.n480 585
R340 B.n2 B.n0 585
R341 B.n4 B.n2 585
R342 B.n3 B.n1 585
R343 B.n634 B.n3 585
R344 B.n632 B.n631 585
R345 B.n633 B.n632 585
R346 B.n630 B.n9 585
R347 B.n9 B.n8 585
R348 B.n629 B.n628 585
R349 B.n628 B.n627 585
R350 B.n11 B.n10 585
R351 B.n626 B.n11 585
R352 B.n624 B.n623 585
R353 B.n625 B.n624 585
R354 B.n622 B.n16 585
R355 B.n16 B.n15 585
R356 B.n621 B.n620 585
R357 B.n620 B.n619 585
R358 B.n18 B.n17 585
R359 B.n618 B.n18 585
R360 B.n616 B.n615 585
R361 B.n617 B.n616 585
R362 B.n614 B.n23 585
R363 B.n23 B.n22 585
R364 B.n613 B.n612 585
R365 B.n612 B.n611 585
R366 B.n25 B.n24 585
R367 B.n610 B.n25 585
R368 B.n608 B.n607 585
R369 B.n609 B.n608 585
R370 B.n606 B.n30 585
R371 B.n30 B.n29 585
R372 B.n605 B.n604 585
R373 B.n604 B.n603 585
R374 B.n32 B.n31 585
R375 B.n602 B.n32 585
R376 B.n600 B.n599 585
R377 B.n601 B.n600 585
R378 B.n598 B.n37 585
R379 B.n37 B.n36 585
R380 B.n597 B.n596 585
R381 B.n596 B.n595 585
R382 B.n39 B.n38 585
R383 B.n594 B.n39 585
R384 B.n592 B.n591 585
R385 B.n593 B.n592 585
R386 B.n590 B.n44 585
R387 B.n44 B.n43 585
R388 B.n589 B.n588 585
R389 B.n588 B.n587 585
R390 B.n46 B.n45 585
R391 B.n586 B.n46 585
R392 B.n584 B.n583 585
R393 B.n585 B.n584 585
R394 B.n582 B.n51 585
R395 B.n51 B.n50 585
R396 B.n581 B.n580 585
R397 B.n580 B.n579 585
R398 B.n53 B.n52 585
R399 B.n578 B.n53 585
R400 B.n576 B.n575 585
R401 B.n577 B.n576 585
R402 B.n574 B.n58 585
R403 B.n58 B.n57 585
R404 B.n573 B.n572 585
R405 B.n572 B.n571 585
R406 B.n60 B.n59 585
R407 B.n570 B.n60 585
R408 B.n568 B.n567 585
R409 B.n569 B.n568 585
R410 B.n566 B.n65 585
R411 B.n65 B.n64 585
R412 B.n565 B.n564 585
R413 B.n564 B.n563 585
R414 B.n67 B.n66 585
R415 B.n562 B.n67 585
R416 B.n560 B.n559 585
R417 B.n561 B.n560 585
R418 B.n558 B.n72 585
R419 B.n72 B.n71 585
R420 B.n557 B.n556 585
R421 B.n556 B.n555 585
R422 B.n74 B.n73 585
R423 B.n554 B.n74 585
R424 B.n552 B.n551 585
R425 B.n553 B.n552 585
R426 B.n550 B.n79 585
R427 B.n79 B.n78 585
R428 B.n549 B.n548 585
R429 B.n548 B.n547 585
R430 B.n81 B.n80 585
R431 B.n546 B.n81 585
R432 B.n637 B.n636 585
R433 B.n636 B.n635 585
R434 B.n346 B.n257 545.355
R435 B.n107 B.n81 545.355
R436 B.n349 B.n259 545.355
R437 B.n543 B.n83 545.355
R438 B.n545 B.n544 256.663
R439 B.n545 B.n99 256.663
R440 B.n545 B.n98 256.663
R441 B.n545 B.n97 256.663
R442 B.n545 B.n96 256.663
R443 B.n545 B.n95 256.663
R444 B.n545 B.n94 256.663
R445 B.n545 B.n93 256.663
R446 B.n545 B.n92 256.663
R447 B.n545 B.n91 256.663
R448 B.n545 B.n90 256.663
R449 B.n545 B.n89 256.663
R450 B.n545 B.n88 256.663
R451 B.n545 B.n87 256.663
R452 B.n545 B.n86 256.663
R453 B.n545 B.n85 256.663
R454 B.n545 B.n84 256.663
R455 B.n348 B.n347 256.663
R456 B.n348 B.n262 256.663
R457 B.n348 B.n263 256.663
R458 B.n348 B.n264 256.663
R459 B.n348 B.n265 256.663
R460 B.n348 B.n266 256.663
R461 B.n348 B.n267 256.663
R462 B.n348 B.n268 256.663
R463 B.n348 B.n269 256.663
R464 B.n348 B.n270 256.663
R465 B.n348 B.n271 256.663
R466 B.n348 B.n272 256.663
R467 B.n348 B.n273 256.663
R468 B.n348 B.n274 256.663
R469 B.n348 B.n275 256.663
R470 B.n348 B.n276 256.663
R471 B.n348 B.n258 212.904
R472 B.n546 B.n545 212.904
R473 B.n281 B.t4 209.752
R474 B.n279 B.t15 209.752
R475 B.n104 B.t12 209.752
R476 B.n101 B.t8 209.752
R477 B.n281 B.t7 204.861
R478 B.n101 B.t10 204.861
R479 B.n279 B.t17 204.861
R480 B.n104 B.t13 204.861
R481 B.n355 B.n257 163.367
R482 B.n355 B.n255 163.367
R483 B.n359 B.n255 163.367
R484 B.n359 B.n249 163.367
R485 B.n367 B.n249 163.367
R486 B.n367 B.n247 163.367
R487 B.n371 B.n247 163.367
R488 B.n371 B.n241 163.367
R489 B.n379 B.n241 163.367
R490 B.n379 B.n239 163.367
R491 B.n383 B.n239 163.367
R492 B.n383 B.n233 163.367
R493 B.n391 B.n233 163.367
R494 B.n391 B.n231 163.367
R495 B.n395 B.n231 163.367
R496 B.n395 B.n225 163.367
R497 B.n403 B.n225 163.367
R498 B.n403 B.n223 163.367
R499 B.n407 B.n223 163.367
R500 B.n407 B.n217 163.367
R501 B.n415 B.n217 163.367
R502 B.n415 B.n215 163.367
R503 B.n419 B.n215 163.367
R504 B.n419 B.n209 163.367
R505 B.n427 B.n209 163.367
R506 B.n427 B.n207 163.367
R507 B.n431 B.n207 163.367
R508 B.n431 B.n201 163.367
R509 B.n439 B.n201 163.367
R510 B.n439 B.n199 163.367
R511 B.n443 B.n199 163.367
R512 B.n443 B.n193 163.367
R513 B.n451 B.n193 163.367
R514 B.n451 B.n191 163.367
R515 B.n455 B.n191 163.367
R516 B.n455 B.n185 163.367
R517 B.n463 B.n185 163.367
R518 B.n463 B.n183 163.367
R519 B.n467 B.n183 163.367
R520 B.n467 B.n177 163.367
R521 B.n476 B.n177 163.367
R522 B.n476 B.n175 163.367
R523 B.n480 B.n175 163.367
R524 B.n480 B.n2 163.367
R525 B.n636 B.n2 163.367
R526 B.n636 B.n3 163.367
R527 B.n632 B.n3 163.367
R528 B.n632 B.n9 163.367
R529 B.n628 B.n9 163.367
R530 B.n628 B.n11 163.367
R531 B.n624 B.n11 163.367
R532 B.n624 B.n16 163.367
R533 B.n620 B.n16 163.367
R534 B.n620 B.n18 163.367
R535 B.n616 B.n18 163.367
R536 B.n616 B.n23 163.367
R537 B.n612 B.n23 163.367
R538 B.n612 B.n25 163.367
R539 B.n608 B.n25 163.367
R540 B.n608 B.n30 163.367
R541 B.n604 B.n30 163.367
R542 B.n604 B.n32 163.367
R543 B.n600 B.n32 163.367
R544 B.n600 B.n37 163.367
R545 B.n596 B.n37 163.367
R546 B.n596 B.n39 163.367
R547 B.n592 B.n39 163.367
R548 B.n592 B.n44 163.367
R549 B.n588 B.n44 163.367
R550 B.n588 B.n46 163.367
R551 B.n584 B.n46 163.367
R552 B.n584 B.n51 163.367
R553 B.n580 B.n51 163.367
R554 B.n580 B.n53 163.367
R555 B.n576 B.n53 163.367
R556 B.n576 B.n58 163.367
R557 B.n572 B.n58 163.367
R558 B.n572 B.n60 163.367
R559 B.n568 B.n60 163.367
R560 B.n568 B.n65 163.367
R561 B.n564 B.n65 163.367
R562 B.n564 B.n67 163.367
R563 B.n560 B.n67 163.367
R564 B.n560 B.n72 163.367
R565 B.n556 B.n72 163.367
R566 B.n556 B.n74 163.367
R567 B.n552 B.n74 163.367
R568 B.n552 B.n79 163.367
R569 B.n548 B.n79 163.367
R570 B.n548 B.n81 163.367
R571 B.n278 B.n277 163.367
R572 B.n341 B.n277 163.367
R573 B.n339 B.n338 163.367
R574 B.n335 B.n334 163.367
R575 B.n331 B.n330 163.367
R576 B.n327 B.n326 163.367
R577 B.n322 B.n321 163.367
R578 B.n318 B.n317 163.367
R579 B.n314 B.n313 163.367
R580 B.n310 B.n309 163.367
R581 B.n306 B.n305 163.367
R582 B.n301 B.n300 163.367
R583 B.n297 B.n296 163.367
R584 B.n293 B.n292 163.367
R585 B.n289 B.n288 163.367
R586 B.n285 B.n284 163.367
R587 B.n349 B.n261 163.367
R588 B.n353 B.n259 163.367
R589 B.n353 B.n253 163.367
R590 B.n361 B.n253 163.367
R591 B.n361 B.n251 163.367
R592 B.n365 B.n251 163.367
R593 B.n365 B.n245 163.367
R594 B.n373 B.n245 163.367
R595 B.n373 B.n243 163.367
R596 B.n377 B.n243 163.367
R597 B.n377 B.n237 163.367
R598 B.n385 B.n237 163.367
R599 B.n385 B.n235 163.367
R600 B.n389 B.n235 163.367
R601 B.n389 B.n229 163.367
R602 B.n397 B.n229 163.367
R603 B.n397 B.n227 163.367
R604 B.n401 B.n227 163.367
R605 B.n401 B.n221 163.367
R606 B.n409 B.n221 163.367
R607 B.n409 B.n219 163.367
R608 B.n413 B.n219 163.367
R609 B.n413 B.n212 163.367
R610 B.n421 B.n212 163.367
R611 B.n421 B.n210 163.367
R612 B.n425 B.n210 163.367
R613 B.n425 B.n205 163.367
R614 B.n433 B.n205 163.367
R615 B.n433 B.n203 163.367
R616 B.n437 B.n203 163.367
R617 B.n437 B.n197 163.367
R618 B.n445 B.n197 163.367
R619 B.n445 B.n195 163.367
R620 B.n449 B.n195 163.367
R621 B.n449 B.n189 163.367
R622 B.n457 B.n189 163.367
R623 B.n457 B.n187 163.367
R624 B.n461 B.n187 163.367
R625 B.n461 B.n181 163.367
R626 B.n469 B.n181 163.367
R627 B.n469 B.n179 163.367
R628 B.n474 B.n179 163.367
R629 B.n474 B.n173 163.367
R630 B.n482 B.n173 163.367
R631 B.n483 B.n482 163.367
R632 B.n483 B.n5 163.367
R633 B.n6 B.n5 163.367
R634 B.n7 B.n6 163.367
R635 B.n488 B.n7 163.367
R636 B.n488 B.n12 163.367
R637 B.n13 B.n12 163.367
R638 B.n14 B.n13 163.367
R639 B.n493 B.n14 163.367
R640 B.n493 B.n19 163.367
R641 B.n20 B.n19 163.367
R642 B.n21 B.n20 163.367
R643 B.n498 B.n21 163.367
R644 B.n498 B.n26 163.367
R645 B.n27 B.n26 163.367
R646 B.n28 B.n27 163.367
R647 B.n503 B.n28 163.367
R648 B.n503 B.n33 163.367
R649 B.n34 B.n33 163.367
R650 B.n35 B.n34 163.367
R651 B.n508 B.n35 163.367
R652 B.n508 B.n40 163.367
R653 B.n41 B.n40 163.367
R654 B.n42 B.n41 163.367
R655 B.n513 B.n42 163.367
R656 B.n513 B.n47 163.367
R657 B.n48 B.n47 163.367
R658 B.n49 B.n48 163.367
R659 B.n518 B.n49 163.367
R660 B.n518 B.n54 163.367
R661 B.n55 B.n54 163.367
R662 B.n56 B.n55 163.367
R663 B.n523 B.n56 163.367
R664 B.n523 B.n61 163.367
R665 B.n62 B.n61 163.367
R666 B.n63 B.n62 163.367
R667 B.n528 B.n63 163.367
R668 B.n528 B.n68 163.367
R669 B.n69 B.n68 163.367
R670 B.n70 B.n69 163.367
R671 B.n533 B.n70 163.367
R672 B.n533 B.n75 163.367
R673 B.n76 B.n75 163.367
R674 B.n77 B.n76 163.367
R675 B.n538 B.n77 163.367
R676 B.n538 B.n82 163.367
R677 B.n83 B.n82 163.367
R678 B.n111 B.n110 163.367
R679 B.n115 B.n114 163.367
R680 B.n119 B.n118 163.367
R681 B.n123 B.n122 163.367
R682 B.n127 B.n126 163.367
R683 B.n131 B.n130 163.367
R684 B.n135 B.n134 163.367
R685 B.n139 B.n138 163.367
R686 B.n143 B.n142 163.367
R687 B.n147 B.n146 163.367
R688 B.n151 B.n150 163.367
R689 B.n155 B.n154 163.367
R690 B.n159 B.n158 163.367
R691 B.n163 B.n162 163.367
R692 B.n167 B.n166 163.367
R693 B.n169 B.n100 163.367
R694 B.n282 B.t6 123.213
R695 B.n102 B.t11 123.213
R696 B.n280 B.t16 123.213
R697 B.n105 B.t14 123.213
R698 B.n354 B.n258 102.677
R699 B.n354 B.n254 102.677
R700 B.n360 B.n254 102.677
R701 B.n360 B.n250 102.677
R702 B.n366 B.n250 102.677
R703 B.n366 B.n246 102.677
R704 B.n372 B.n246 102.677
R705 B.n372 B.n242 102.677
R706 B.n378 B.n242 102.677
R707 B.n384 B.n238 102.677
R708 B.n384 B.n234 102.677
R709 B.n390 B.n234 102.677
R710 B.n390 B.n230 102.677
R711 B.n396 B.n230 102.677
R712 B.n396 B.n226 102.677
R713 B.n402 B.n226 102.677
R714 B.n402 B.n222 102.677
R715 B.n408 B.n222 102.677
R716 B.n408 B.n218 102.677
R717 B.n414 B.n218 102.677
R718 B.n414 B.n213 102.677
R719 B.n420 B.n213 102.677
R720 B.n420 B.n214 102.677
R721 B.n426 B.n206 102.677
R722 B.n432 B.n206 102.677
R723 B.n432 B.n202 102.677
R724 B.n438 B.n202 102.677
R725 B.n438 B.n198 102.677
R726 B.n444 B.n198 102.677
R727 B.n444 B.n194 102.677
R728 B.n450 B.n194 102.677
R729 B.n450 B.n190 102.677
R730 B.n456 B.n190 102.677
R731 B.n456 B.n186 102.677
R732 B.n462 B.n186 102.677
R733 B.n468 B.n182 102.677
R734 B.n468 B.n178 102.677
R735 B.n475 B.n178 102.677
R736 B.n475 B.n174 102.677
R737 B.n481 B.n174 102.677
R738 B.n481 B.n4 102.677
R739 B.n635 B.n4 102.677
R740 B.n635 B.n634 102.677
R741 B.n634 B.n633 102.677
R742 B.n633 B.n8 102.677
R743 B.n627 B.n8 102.677
R744 B.n627 B.n626 102.677
R745 B.n626 B.n625 102.677
R746 B.n625 B.n15 102.677
R747 B.n619 B.n618 102.677
R748 B.n618 B.n617 102.677
R749 B.n617 B.n22 102.677
R750 B.n611 B.n22 102.677
R751 B.n611 B.n610 102.677
R752 B.n610 B.n609 102.677
R753 B.n609 B.n29 102.677
R754 B.n603 B.n29 102.677
R755 B.n603 B.n602 102.677
R756 B.n602 B.n601 102.677
R757 B.n601 B.n36 102.677
R758 B.n595 B.n36 102.677
R759 B.n594 B.n593 102.677
R760 B.n593 B.n43 102.677
R761 B.n587 B.n43 102.677
R762 B.n587 B.n586 102.677
R763 B.n586 B.n585 102.677
R764 B.n585 B.n50 102.677
R765 B.n579 B.n50 102.677
R766 B.n579 B.n578 102.677
R767 B.n578 B.n577 102.677
R768 B.n577 B.n57 102.677
R769 B.n571 B.n57 102.677
R770 B.n571 B.n570 102.677
R771 B.n570 B.n569 102.677
R772 B.n569 B.n64 102.677
R773 B.n563 B.n562 102.677
R774 B.n562 B.n561 102.677
R775 B.n561 B.n71 102.677
R776 B.n555 B.n71 102.677
R777 B.n555 B.n554 102.677
R778 B.n554 B.n553 102.677
R779 B.n553 B.n78 102.677
R780 B.n547 B.n78 102.677
R781 B.n547 B.n546 102.677
R782 B.n214 B.t1 84.5578
R783 B.t2 B.n594 84.5578
R784 B.n282 B.n281 81.649
R785 B.n280 B.n279 81.649
R786 B.n105 B.n104 81.649
R787 B.n102 B.n101 81.649
R788 B.t0 B.n182 81.5379
R789 B.t3 B.n15 81.5379
R790 B.t5 B.n238 78.518
R791 B.t9 B.n64 78.518
R792 B.n347 B.n346 71.676
R793 B.n341 B.n262 71.676
R794 B.n338 B.n263 71.676
R795 B.n334 B.n264 71.676
R796 B.n330 B.n265 71.676
R797 B.n326 B.n266 71.676
R798 B.n321 B.n267 71.676
R799 B.n317 B.n268 71.676
R800 B.n313 B.n269 71.676
R801 B.n309 B.n270 71.676
R802 B.n305 B.n271 71.676
R803 B.n300 B.n272 71.676
R804 B.n296 B.n273 71.676
R805 B.n292 B.n274 71.676
R806 B.n288 B.n275 71.676
R807 B.n284 B.n276 71.676
R808 B.n107 B.n84 71.676
R809 B.n111 B.n85 71.676
R810 B.n115 B.n86 71.676
R811 B.n119 B.n87 71.676
R812 B.n123 B.n88 71.676
R813 B.n127 B.n89 71.676
R814 B.n131 B.n90 71.676
R815 B.n135 B.n91 71.676
R816 B.n139 B.n92 71.676
R817 B.n143 B.n93 71.676
R818 B.n147 B.n94 71.676
R819 B.n151 B.n95 71.676
R820 B.n155 B.n96 71.676
R821 B.n159 B.n97 71.676
R822 B.n163 B.n98 71.676
R823 B.n167 B.n99 71.676
R824 B.n544 B.n100 71.676
R825 B.n544 B.n543 71.676
R826 B.n169 B.n99 71.676
R827 B.n166 B.n98 71.676
R828 B.n162 B.n97 71.676
R829 B.n158 B.n96 71.676
R830 B.n154 B.n95 71.676
R831 B.n150 B.n94 71.676
R832 B.n146 B.n93 71.676
R833 B.n142 B.n92 71.676
R834 B.n138 B.n91 71.676
R835 B.n134 B.n90 71.676
R836 B.n130 B.n89 71.676
R837 B.n126 B.n88 71.676
R838 B.n122 B.n87 71.676
R839 B.n118 B.n86 71.676
R840 B.n114 B.n85 71.676
R841 B.n110 B.n84 71.676
R842 B.n347 B.n278 71.676
R843 B.n339 B.n262 71.676
R844 B.n335 B.n263 71.676
R845 B.n331 B.n264 71.676
R846 B.n327 B.n265 71.676
R847 B.n322 B.n266 71.676
R848 B.n318 B.n267 71.676
R849 B.n314 B.n268 71.676
R850 B.n310 B.n269 71.676
R851 B.n306 B.n270 71.676
R852 B.n301 B.n271 71.676
R853 B.n297 B.n272 71.676
R854 B.n293 B.n273 71.676
R855 B.n289 B.n274 71.676
R856 B.n285 B.n275 71.676
R857 B.n276 B.n261 71.676
R858 B.n303 B.n282 59.5399
R859 B.n324 B.n280 59.5399
R860 B.n106 B.n105 59.5399
R861 B.n103 B.n102 59.5399
R862 B.n108 B.n80 35.4346
R863 B.n542 B.n541 35.4346
R864 B.n351 B.n350 35.4346
R865 B.n345 B.n256 35.4346
R866 B.n378 B.t5 24.1597
R867 B.n563 B.t9 24.1597
R868 B.n462 B.t0 21.1398
R869 B.n619 B.t3 21.1398
R870 B.n426 B.t1 18.1199
R871 B.n595 B.t2 18.1199
R872 B B.n637 18.0485
R873 B.n109 B.n108 10.6151
R874 B.n112 B.n109 10.6151
R875 B.n113 B.n112 10.6151
R876 B.n116 B.n113 10.6151
R877 B.n117 B.n116 10.6151
R878 B.n120 B.n117 10.6151
R879 B.n121 B.n120 10.6151
R880 B.n124 B.n121 10.6151
R881 B.n125 B.n124 10.6151
R882 B.n128 B.n125 10.6151
R883 B.n129 B.n128 10.6151
R884 B.n133 B.n132 10.6151
R885 B.n136 B.n133 10.6151
R886 B.n137 B.n136 10.6151
R887 B.n140 B.n137 10.6151
R888 B.n141 B.n140 10.6151
R889 B.n144 B.n141 10.6151
R890 B.n145 B.n144 10.6151
R891 B.n148 B.n145 10.6151
R892 B.n149 B.n148 10.6151
R893 B.n153 B.n152 10.6151
R894 B.n156 B.n153 10.6151
R895 B.n157 B.n156 10.6151
R896 B.n160 B.n157 10.6151
R897 B.n161 B.n160 10.6151
R898 B.n164 B.n161 10.6151
R899 B.n165 B.n164 10.6151
R900 B.n168 B.n165 10.6151
R901 B.n170 B.n168 10.6151
R902 B.n171 B.n170 10.6151
R903 B.n542 B.n171 10.6151
R904 B.n352 B.n351 10.6151
R905 B.n352 B.n252 10.6151
R906 B.n362 B.n252 10.6151
R907 B.n363 B.n362 10.6151
R908 B.n364 B.n363 10.6151
R909 B.n364 B.n244 10.6151
R910 B.n374 B.n244 10.6151
R911 B.n375 B.n374 10.6151
R912 B.n376 B.n375 10.6151
R913 B.n376 B.n236 10.6151
R914 B.n386 B.n236 10.6151
R915 B.n387 B.n386 10.6151
R916 B.n388 B.n387 10.6151
R917 B.n388 B.n228 10.6151
R918 B.n398 B.n228 10.6151
R919 B.n399 B.n398 10.6151
R920 B.n400 B.n399 10.6151
R921 B.n400 B.n220 10.6151
R922 B.n410 B.n220 10.6151
R923 B.n411 B.n410 10.6151
R924 B.n412 B.n411 10.6151
R925 B.n412 B.n211 10.6151
R926 B.n422 B.n211 10.6151
R927 B.n423 B.n422 10.6151
R928 B.n424 B.n423 10.6151
R929 B.n424 B.n204 10.6151
R930 B.n434 B.n204 10.6151
R931 B.n435 B.n434 10.6151
R932 B.n436 B.n435 10.6151
R933 B.n436 B.n196 10.6151
R934 B.n446 B.n196 10.6151
R935 B.n447 B.n446 10.6151
R936 B.n448 B.n447 10.6151
R937 B.n448 B.n188 10.6151
R938 B.n458 B.n188 10.6151
R939 B.n459 B.n458 10.6151
R940 B.n460 B.n459 10.6151
R941 B.n460 B.n180 10.6151
R942 B.n470 B.n180 10.6151
R943 B.n471 B.n470 10.6151
R944 B.n473 B.n471 10.6151
R945 B.n473 B.n472 10.6151
R946 B.n472 B.n172 10.6151
R947 B.n484 B.n172 10.6151
R948 B.n485 B.n484 10.6151
R949 B.n486 B.n485 10.6151
R950 B.n487 B.n486 10.6151
R951 B.n489 B.n487 10.6151
R952 B.n490 B.n489 10.6151
R953 B.n491 B.n490 10.6151
R954 B.n492 B.n491 10.6151
R955 B.n494 B.n492 10.6151
R956 B.n495 B.n494 10.6151
R957 B.n496 B.n495 10.6151
R958 B.n497 B.n496 10.6151
R959 B.n499 B.n497 10.6151
R960 B.n500 B.n499 10.6151
R961 B.n501 B.n500 10.6151
R962 B.n502 B.n501 10.6151
R963 B.n504 B.n502 10.6151
R964 B.n505 B.n504 10.6151
R965 B.n506 B.n505 10.6151
R966 B.n507 B.n506 10.6151
R967 B.n509 B.n507 10.6151
R968 B.n510 B.n509 10.6151
R969 B.n511 B.n510 10.6151
R970 B.n512 B.n511 10.6151
R971 B.n514 B.n512 10.6151
R972 B.n515 B.n514 10.6151
R973 B.n516 B.n515 10.6151
R974 B.n517 B.n516 10.6151
R975 B.n519 B.n517 10.6151
R976 B.n520 B.n519 10.6151
R977 B.n521 B.n520 10.6151
R978 B.n522 B.n521 10.6151
R979 B.n524 B.n522 10.6151
R980 B.n525 B.n524 10.6151
R981 B.n526 B.n525 10.6151
R982 B.n527 B.n526 10.6151
R983 B.n529 B.n527 10.6151
R984 B.n530 B.n529 10.6151
R985 B.n531 B.n530 10.6151
R986 B.n532 B.n531 10.6151
R987 B.n534 B.n532 10.6151
R988 B.n535 B.n534 10.6151
R989 B.n536 B.n535 10.6151
R990 B.n537 B.n536 10.6151
R991 B.n539 B.n537 10.6151
R992 B.n540 B.n539 10.6151
R993 B.n541 B.n540 10.6151
R994 B.n345 B.n344 10.6151
R995 B.n344 B.n343 10.6151
R996 B.n343 B.n342 10.6151
R997 B.n342 B.n340 10.6151
R998 B.n340 B.n337 10.6151
R999 B.n337 B.n336 10.6151
R1000 B.n336 B.n333 10.6151
R1001 B.n333 B.n332 10.6151
R1002 B.n332 B.n329 10.6151
R1003 B.n329 B.n328 10.6151
R1004 B.n328 B.n325 10.6151
R1005 B.n323 B.n320 10.6151
R1006 B.n320 B.n319 10.6151
R1007 B.n319 B.n316 10.6151
R1008 B.n316 B.n315 10.6151
R1009 B.n315 B.n312 10.6151
R1010 B.n312 B.n311 10.6151
R1011 B.n311 B.n308 10.6151
R1012 B.n308 B.n307 10.6151
R1013 B.n307 B.n304 10.6151
R1014 B.n302 B.n299 10.6151
R1015 B.n299 B.n298 10.6151
R1016 B.n298 B.n295 10.6151
R1017 B.n295 B.n294 10.6151
R1018 B.n294 B.n291 10.6151
R1019 B.n291 B.n290 10.6151
R1020 B.n290 B.n287 10.6151
R1021 B.n287 B.n286 10.6151
R1022 B.n286 B.n283 10.6151
R1023 B.n283 B.n260 10.6151
R1024 B.n350 B.n260 10.6151
R1025 B.n356 B.n256 10.6151
R1026 B.n357 B.n356 10.6151
R1027 B.n358 B.n357 10.6151
R1028 B.n358 B.n248 10.6151
R1029 B.n368 B.n248 10.6151
R1030 B.n369 B.n368 10.6151
R1031 B.n370 B.n369 10.6151
R1032 B.n370 B.n240 10.6151
R1033 B.n380 B.n240 10.6151
R1034 B.n381 B.n380 10.6151
R1035 B.n382 B.n381 10.6151
R1036 B.n382 B.n232 10.6151
R1037 B.n392 B.n232 10.6151
R1038 B.n393 B.n392 10.6151
R1039 B.n394 B.n393 10.6151
R1040 B.n394 B.n224 10.6151
R1041 B.n404 B.n224 10.6151
R1042 B.n405 B.n404 10.6151
R1043 B.n406 B.n405 10.6151
R1044 B.n406 B.n216 10.6151
R1045 B.n416 B.n216 10.6151
R1046 B.n417 B.n416 10.6151
R1047 B.n418 B.n417 10.6151
R1048 B.n418 B.n208 10.6151
R1049 B.n428 B.n208 10.6151
R1050 B.n429 B.n428 10.6151
R1051 B.n430 B.n429 10.6151
R1052 B.n430 B.n200 10.6151
R1053 B.n440 B.n200 10.6151
R1054 B.n441 B.n440 10.6151
R1055 B.n442 B.n441 10.6151
R1056 B.n442 B.n192 10.6151
R1057 B.n452 B.n192 10.6151
R1058 B.n453 B.n452 10.6151
R1059 B.n454 B.n453 10.6151
R1060 B.n454 B.n184 10.6151
R1061 B.n464 B.n184 10.6151
R1062 B.n465 B.n464 10.6151
R1063 B.n466 B.n465 10.6151
R1064 B.n466 B.n176 10.6151
R1065 B.n477 B.n176 10.6151
R1066 B.n478 B.n477 10.6151
R1067 B.n479 B.n478 10.6151
R1068 B.n479 B.n0 10.6151
R1069 B.n631 B.n1 10.6151
R1070 B.n631 B.n630 10.6151
R1071 B.n630 B.n629 10.6151
R1072 B.n629 B.n10 10.6151
R1073 B.n623 B.n10 10.6151
R1074 B.n623 B.n622 10.6151
R1075 B.n622 B.n621 10.6151
R1076 B.n621 B.n17 10.6151
R1077 B.n615 B.n17 10.6151
R1078 B.n615 B.n614 10.6151
R1079 B.n614 B.n613 10.6151
R1080 B.n613 B.n24 10.6151
R1081 B.n607 B.n24 10.6151
R1082 B.n607 B.n606 10.6151
R1083 B.n606 B.n605 10.6151
R1084 B.n605 B.n31 10.6151
R1085 B.n599 B.n31 10.6151
R1086 B.n599 B.n598 10.6151
R1087 B.n598 B.n597 10.6151
R1088 B.n597 B.n38 10.6151
R1089 B.n591 B.n38 10.6151
R1090 B.n591 B.n590 10.6151
R1091 B.n590 B.n589 10.6151
R1092 B.n589 B.n45 10.6151
R1093 B.n583 B.n45 10.6151
R1094 B.n583 B.n582 10.6151
R1095 B.n582 B.n581 10.6151
R1096 B.n581 B.n52 10.6151
R1097 B.n575 B.n52 10.6151
R1098 B.n575 B.n574 10.6151
R1099 B.n574 B.n573 10.6151
R1100 B.n573 B.n59 10.6151
R1101 B.n567 B.n59 10.6151
R1102 B.n567 B.n566 10.6151
R1103 B.n566 B.n565 10.6151
R1104 B.n565 B.n66 10.6151
R1105 B.n559 B.n66 10.6151
R1106 B.n559 B.n558 10.6151
R1107 B.n558 B.n557 10.6151
R1108 B.n557 B.n73 10.6151
R1109 B.n551 B.n73 10.6151
R1110 B.n551 B.n550 10.6151
R1111 B.n550 B.n549 10.6151
R1112 B.n549 B.n80 10.6151
R1113 B.n129 B.n106 9.36635
R1114 B.n152 B.n103 9.36635
R1115 B.n325 B.n324 9.36635
R1116 B.n303 B.n302 9.36635
R1117 B.n637 B.n0 2.81026
R1118 B.n637 B.n1 2.81026
R1119 B.n132 B.n106 1.24928
R1120 B.n149 B.n103 1.24928
R1121 B.n324 B.n323 1.24928
R1122 B.n304 B.n303 1.24928
R1123 VN.n0 VN.t0 46.8985
R1124 VN.n1 VN.t3 46.8985
R1125 VN.n0 VN.t2 45.5287
R1126 VN.n1 VN.t1 45.5287
R1127 VN VN.n1 44.7395
R1128 VN VN.n0 1.79633
R1129 VDD2.n2 VDD2.n0 137.326
R1130 VDD2.n2 VDD2.n1 100.99
R1131 VDD2.n1 VDD2.t3 9.85125
R1132 VDD2.n1 VDD2.t1 9.85125
R1133 VDD2.n0 VDD2.t0 9.85125
R1134 VDD2.n0 VDD2.t2 9.85125
R1135 VDD2 VDD2.n2 0.0586897
R1136 VTAIL.n58 VTAIL.n56 289.615
R1137 VTAIL.n2 VTAIL.n0 289.615
R1138 VTAIL.n10 VTAIL.n8 289.615
R1139 VTAIL.n18 VTAIL.n16 289.615
R1140 VTAIL.n50 VTAIL.n48 289.615
R1141 VTAIL.n42 VTAIL.n40 289.615
R1142 VTAIL.n34 VTAIL.n32 289.615
R1143 VTAIL.n26 VTAIL.n24 289.615
R1144 VTAIL.n59 VTAIL.n58 185
R1145 VTAIL.n3 VTAIL.n2 185
R1146 VTAIL.n11 VTAIL.n10 185
R1147 VTAIL.n19 VTAIL.n18 185
R1148 VTAIL.n51 VTAIL.n50 185
R1149 VTAIL.n43 VTAIL.n42 185
R1150 VTAIL.n35 VTAIL.n34 185
R1151 VTAIL.n27 VTAIL.n26 185
R1152 VTAIL.t5 VTAIL.n57 167.117
R1153 VTAIL.t7 VTAIL.n1 167.117
R1154 VTAIL.t1 VTAIL.n9 167.117
R1155 VTAIL.t0 VTAIL.n17 167.117
R1156 VTAIL.t2 VTAIL.n49 167.117
R1157 VTAIL.t3 VTAIL.n41 167.117
R1158 VTAIL.t4 VTAIL.n33 167.117
R1159 VTAIL.t6 VTAIL.n25 167.117
R1160 VTAIL.n58 VTAIL.t5 52.3082
R1161 VTAIL.n2 VTAIL.t7 52.3082
R1162 VTAIL.n10 VTAIL.t1 52.3082
R1163 VTAIL.n18 VTAIL.t0 52.3082
R1164 VTAIL.n50 VTAIL.t2 52.3082
R1165 VTAIL.n42 VTAIL.t3 52.3082
R1166 VTAIL.n34 VTAIL.t4 52.3082
R1167 VTAIL.n26 VTAIL.t6 52.3082
R1168 VTAIL.n63 VTAIL.n62 31.6035
R1169 VTAIL.n7 VTAIL.n6 31.6035
R1170 VTAIL.n15 VTAIL.n14 31.6035
R1171 VTAIL.n23 VTAIL.n22 31.6035
R1172 VTAIL.n55 VTAIL.n54 31.6035
R1173 VTAIL.n47 VTAIL.n46 31.6035
R1174 VTAIL.n39 VTAIL.n38 31.6035
R1175 VTAIL.n31 VTAIL.n30 31.6035
R1176 VTAIL.n63 VTAIL.n55 17.7289
R1177 VTAIL.n31 VTAIL.n23 17.7289
R1178 VTAIL.n59 VTAIL.n57 9.71174
R1179 VTAIL.n3 VTAIL.n1 9.71174
R1180 VTAIL.n11 VTAIL.n9 9.71174
R1181 VTAIL.n19 VTAIL.n17 9.71174
R1182 VTAIL.n51 VTAIL.n49 9.71174
R1183 VTAIL.n43 VTAIL.n41 9.71174
R1184 VTAIL.n35 VTAIL.n33 9.71174
R1185 VTAIL.n27 VTAIL.n25 9.71174
R1186 VTAIL.n62 VTAIL.n61 9.45567
R1187 VTAIL.n6 VTAIL.n5 9.45567
R1188 VTAIL.n14 VTAIL.n13 9.45567
R1189 VTAIL.n22 VTAIL.n21 9.45567
R1190 VTAIL.n54 VTAIL.n53 9.45567
R1191 VTAIL.n46 VTAIL.n45 9.45567
R1192 VTAIL.n38 VTAIL.n37 9.45567
R1193 VTAIL.n30 VTAIL.n29 9.45567
R1194 VTAIL.n61 VTAIL.n60 9.3005
R1195 VTAIL.n5 VTAIL.n4 9.3005
R1196 VTAIL.n13 VTAIL.n12 9.3005
R1197 VTAIL.n21 VTAIL.n20 9.3005
R1198 VTAIL.n53 VTAIL.n52 9.3005
R1199 VTAIL.n45 VTAIL.n44 9.3005
R1200 VTAIL.n37 VTAIL.n36 9.3005
R1201 VTAIL.n29 VTAIL.n28 9.3005
R1202 VTAIL.n62 VTAIL.n56 8.14595
R1203 VTAIL.n6 VTAIL.n0 8.14595
R1204 VTAIL.n14 VTAIL.n8 8.14595
R1205 VTAIL.n22 VTAIL.n16 8.14595
R1206 VTAIL.n54 VTAIL.n48 8.14595
R1207 VTAIL.n46 VTAIL.n40 8.14595
R1208 VTAIL.n38 VTAIL.n32 8.14595
R1209 VTAIL.n30 VTAIL.n24 8.14595
R1210 VTAIL.n60 VTAIL.n59 7.3702
R1211 VTAIL.n4 VTAIL.n3 7.3702
R1212 VTAIL.n12 VTAIL.n11 7.3702
R1213 VTAIL.n20 VTAIL.n19 7.3702
R1214 VTAIL.n52 VTAIL.n51 7.3702
R1215 VTAIL.n44 VTAIL.n43 7.3702
R1216 VTAIL.n36 VTAIL.n35 7.3702
R1217 VTAIL.n28 VTAIL.n27 7.3702
R1218 VTAIL.n60 VTAIL.n56 5.81868
R1219 VTAIL.n4 VTAIL.n0 5.81868
R1220 VTAIL.n12 VTAIL.n8 5.81868
R1221 VTAIL.n20 VTAIL.n16 5.81868
R1222 VTAIL.n52 VTAIL.n48 5.81868
R1223 VTAIL.n44 VTAIL.n40 5.81868
R1224 VTAIL.n36 VTAIL.n32 5.81868
R1225 VTAIL.n28 VTAIL.n24 5.81868
R1226 VTAIL.n39 VTAIL.n31 3.62981
R1227 VTAIL.n55 VTAIL.n47 3.62981
R1228 VTAIL.n23 VTAIL.n15 3.62981
R1229 VTAIL.n61 VTAIL.n57 3.44771
R1230 VTAIL.n5 VTAIL.n1 3.44771
R1231 VTAIL.n13 VTAIL.n9 3.44771
R1232 VTAIL.n21 VTAIL.n17 3.44771
R1233 VTAIL.n53 VTAIL.n49 3.44771
R1234 VTAIL.n45 VTAIL.n41 3.44771
R1235 VTAIL.n37 VTAIL.n33 3.44771
R1236 VTAIL.n29 VTAIL.n25 3.44771
R1237 VTAIL VTAIL.n7 1.87334
R1238 VTAIL VTAIL.n63 1.75697
R1239 VTAIL.n47 VTAIL.n39 0.470328
R1240 VTAIL.n15 VTAIL.n7 0.470328
R1241 VP.n21 VP.n20 161.3
R1242 VP.n19 VP.n1 161.3
R1243 VP.n18 VP.n17 161.3
R1244 VP.n16 VP.n2 161.3
R1245 VP.n15 VP.n14 161.3
R1246 VP.n13 VP.n3 161.3
R1247 VP.n12 VP.n11 161.3
R1248 VP.n10 VP.n4 161.3
R1249 VP.n9 VP.n8 161.3
R1250 VP.n7 VP.n6 84.9293
R1251 VP.n22 VP.n0 84.9293
R1252 VP.n5 VP.t2 46.8983
R1253 VP.n5 VP.t1 45.5287
R1254 VP.n6 VP.n5 44.5742
R1255 VP.n14 VP.n13 40.4934
R1256 VP.n14 VP.n2 40.4934
R1257 VP.n8 VP.n4 24.4675
R1258 VP.n12 VP.n4 24.4675
R1259 VP.n13 VP.n12 24.4675
R1260 VP.n18 VP.n2 24.4675
R1261 VP.n19 VP.n18 24.4675
R1262 VP.n20 VP.n19 24.4675
R1263 VP.n7 VP.t3 12.4853
R1264 VP.n0 VP.t0 12.4853
R1265 VP.n8 VP.n7 5.13857
R1266 VP.n20 VP.n0 5.13857
R1267 VP.n9 VP.n6 0.354971
R1268 VP.n22 VP.n21 0.354971
R1269 VP VP.n22 0.26696
R1270 VP.n10 VP.n9 0.189894
R1271 VP.n11 VP.n10 0.189894
R1272 VP.n11 VP.n3 0.189894
R1273 VP.n15 VP.n3 0.189894
R1274 VP.n16 VP.n15 0.189894
R1275 VP.n17 VP.n16 0.189894
R1276 VP.n17 VP.n1 0.189894
R1277 VP.n21 VP.n1 0.189894
R1278 VDD1 VDD1.n1 137.85
R1279 VDD1 VDD1.n0 101.047
R1280 VDD1.n0 VDD1.t1 9.85125
R1281 VDD1.n0 VDD1.t2 9.85125
R1282 VDD1.n1 VDD1.t0 9.85125
R1283 VDD1.n1 VDD1.t3 9.85125
C0 VTAIL VDD1 3.71228f
C1 VN VP 5.26875f
C2 VTAIL VP 2.00457f
C3 VN VTAIL 1.99046f
C4 VDD2 VDD1 1.33877f
C5 VDD2 VP 0.482372f
C6 VN VDD2 1.13282f
C7 VDD2 VTAIL 3.77506f
C8 VDD1 VP 1.45718f
C9 VN VDD1 0.155758f
C10 VDD2 B 3.653999f
C11 VDD1 B 6.56964f
C12 VTAIL B 4.218097f
C13 VN B 11.977301f
C14 VP B 10.705782f
C15 VDD1.t1 B 0.035692f
C16 VDD1.t2 B 0.035692f
C17 VDD1.n0 B 0.224598f
C18 VDD1.t0 B 0.035692f
C19 VDD1.t3 B 0.035692f
C20 VDD1.n1 B 0.47889f
C21 VP.t0 B 0.484238f
C22 VP.n0 B 0.322935f
C23 VP.n1 B 0.026561f
C24 VP.n2 B 0.052789f
C25 VP.n3 B 0.026561f
C26 VP.n4 B 0.049502f
C27 VP.t2 B 0.807858f
C28 VP.t1 B 0.793823f
C29 VP.n5 B 1.98449f
C30 VP.n6 B 1.30212f
C31 VP.t3 B 0.484238f
C32 VP.n7 B 0.322935f
C33 VP.n8 B 0.030194f
C34 VP.n9 B 0.042868f
C35 VP.n10 B 0.026561f
C36 VP.n11 B 0.026561f
C37 VP.n12 B 0.049502f
C38 VP.n13 B 0.052789f
C39 VP.n14 B 0.021472f
C40 VP.n15 B 0.026561f
C41 VP.n16 B 0.026561f
C42 VP.n17 B 0.026561f
C43 VP.n18 B 0.049502f
C44 VP.n19 B 0.049502f
C45 VP.n20 B 0.030194f
C46 VP.n21 B 0.042868f
C47 VP.n22 B 0.080872f
C48 VTAIL.n0 B 0.035892f
C49 VTAIL.n1 B 0.07936f
C50 VTAIL.t7 B 0.059531f
C51 VTAIL.n2 B 0.06216f
C52 VTAIL.n3 B 0.019944f
C53 VTAIL.n4 B 0.013153f
C54 VTAIL.n5 B 0.175249f
C55 VTAIL.n6 B 0.039369f
C56 VTAIL.n7 B 0.205115f
C57 VTAIL.n8 B 0.035892f
C58 VTAIL.n9 B 0.07936f
C59 VTAIL.t1 B 0.059531f
C60 VTAIL.n10 B 0.06216f
C61 VTAIL.n11 B 0.019944f
C62 VTAIL.n12 B 0.013153f
C63 VTAIL.n13 B 0.175249f
C64 VTAIL.n14 B 0.039369f
C65 VTAIL.n15 B 0.343654f
C66 VTAIL.n16 B 0.035892f
C67 VTAIL.n17 B 0.07936f
C68 VTAIL.t0 B 0.059531f
C69 VTAIL.n18 B 0.06216f
C70 VTAIL.n19 B 0.019944f
C71 VTAIL.n20 B 0.013153f
C72 VTAIL.n21 B 0.175249f
C73 VTAIL.n22 B 0.039369f
C74 VTAIL.n23 B 1.06203f
C75 VTAIL.n24 B 0.035892f
C76 VTAIL.n25 B 0.07936f
C77 VTAIL.t6 B 0.059531f
C78 VTAIL.n26 B 0.06216f
C79 VTAIL.n27 B 0.019944f
C80 VTAIL.n28 B 0.013153f
C81 VTAIL.n29 B 0.175249f
C82 VTAIL.n30 B 0.039369f
C83 VTAIL.n31 B 1.06203f
C84 VTAIL.n32 B 0.035892f
C85 VTAIL.n33 B 0.07936f
C86 VTAIL.t4 B 0.059531f
C87 VTAIL.n34 B 0.06216f
C88 VTAIL.n35 B 0.019944f
C89 VTAIL.n36 B 0.013153f
C90 VTAIL.n37 B 0.175249f
C91 VTAIL.n38 B 0.039369f
C92 VTAIL.n39 B 0.343654f
C93 VTAIL.n40 B 0.035892f
C94 VTAIL.n41 B 0.07936f
C95 VTAIL.t3 B 0.059531f
C96 VTAIL.n42 B 0.06216f
C97 VTAIL.n43 B 0.019944f
C98 VTAIL.n44 B 0.013153f
C99 VTAIL.n45 B 0.175249f
C100 VTAIL.n46 B 0.039369f
C101 VTAIL.n47 B 0.343654f
C102 VTAIL.n48 B 0.035892f
C103 VTAIL.n49 B 0.07936f
C104 VTAIL.t2 B 0.059531f
C105 VTAIL.n50 B 0.06216f
C106 VTAIL.n51 B 0.019944f
C107 VTAIL.n52 B 0.013153f
C108 VTAIL.n53 B 0.175249f
C109 VTAIL.n54 B 0.039369f
C110 VTAIL.n55 B 1.06203f
C111 VTAIL.n56 B 0.035892f
C112 VTAIL.n57 B 0.07936f
C113 VTAIL.t5 B 0.059531f
C114 VTAIL.n58 B 0.06216f
C115 VTAIL.n59 B 0.019944f
C116 VTAIL.n60 B 0.013153f
C117 VTAIL.n61 B 0.175249f
C118 VTAIL.n62 B 0.039369f
C119 VTAIL.n63 B 0.914309f
C120 VDD2.t0 B 0.037497f
C121 VDD2.t2 B 0.037497f
C122 VDD2.n0 B 0.487812f
C123 VDD2.t3 B 0.037497f
C124 VDD2.t1 B 0.037497f
C125 VDD2.n1 B 0.23569f
C126 VDD2.n2 B 2.64535f
C127 VN.t2 B 0.573404f
C128 VN.t0 B 0.583543f
C129 VN.n0 B 0.403114f
C130 VN.t1 B 0.573404f
C131 VN.t3 B 0.583543f
C132 VN.n1 B 1.44159f
.ends

