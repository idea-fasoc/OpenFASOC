* NGSPICE file created from diff_pair_sample_0029.ext - technology: sky130A

.subckt diff_pair_sample_0029 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=0 ps=0 w=6.37 l=3.02
X2 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X3 VDD2.t6 VN.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=2.4843 ps=13.52 w=6.37 l=3.02
X4 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=0 ps=0 w=6.37 l=3.02
X5 VTAIL.t14 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X6 VTAIL.t4 VN.t2 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=1.05105 ps=6.7 w=6.37 l=3.02
X7 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X8 VTAIL.t3 VN.t4 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=1.05105 ps=6.7 w=6.37 l=3.02
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=0 ps=0 w=6.37 l=3.02
X10 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X11 VTAIL.t11 VP.t2 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=1.05105 ps=6.7 w=6.37 l=3.02
X12 VTAIL.t15 VP.t3 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=1.05105 ps=6.7 w=6.37 l=3.02
X13 VDD1.t3 VP.t4 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X14 VDD2.t1 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=2.4843 ps=13.52 w=6.37 l=3.02
X15 VDD2.t0 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
X16 VDD1.t2 VP.t5 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=2.4843 ps=13.52 w=6.37 l=3.02
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4843 pd=13.52 as=0 ps=0 w=6.37 l=3.02
X18 VDD1.t1 VP.t6 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=2.4843 ps=13.52 w=6.37 l=3.02
X19 VTAIL.t13 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.05105 pd=6.7 as=1.05105 ps=6.7 w=6.37 l=3.02
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n29 VP.n16 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n15 161.3
R8 VP.n35 VP.n34 161.3
R9 VP.n36 VP.n14 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n39 VP.n13 161.3
R12 VP.n41 VP.n40 161.3
R13 VP.n42 VP.n12 161.3
R14 VP.n78 VP.n0 161.3
R15 VP.n77 VP.n76 161.3
R16 VP.n75 VP.n1 161.3
R17 VP.n74 VP.n73 161.3
R18 VP.n72 VP.n2 161.3
R19 VP.n71 VP.n70 161.3
R20 VP.n69 VP.n3 161.3
R21 VP.n68 VP.n67 161.3
R22 VP.n65 VP.n4 161.3
R23 VP.n64 VP.n63 161.3
R24 VP.n62 VP.n5 161.3
R25 VP.n61 VP.n60 161.3
R26 VP.n59 VP.n6 161.3
R27 VP.n58 VP.n57 161.3
R28 VP.n56 VP.n55 161.3
R29 VP.n54 VP.n8 161.3
R30 VP.n53 VP.n52 161.3
R31 VP.n51 VP.n9 161.3
R32 VP.n50 VP.n49 161.3
R33 VP.n48 VP.n10 161.3
R34 VP.n47 VP.n46 161.3
R35 VP.n45 VP.n11 109.534
R36 VP.n80 VP.n79 109.534
R37 VP.n44 VP.n43 109.534
R38 VP.n20 VP.t2 83.102
R39 VP.n20 VP.n19 65.4202
R40 VP.n53 VP.n9 55.0624
R41 VP.n73 VP.n72 55.0624
R42 VP.n37 VP.n36 55.0624
R43 VP.n11 VP.t3 50.8339
R44 VP.n7 VP.t4 50.8339
R45 VP.n66 VP.t7 50.8339
R46 VP.n79 VP.t5 50.8339
R47 VP.n43 VP.t6 50.8339
R48 VP.n30 VP.t1 50.8339
R49 VP.n19 VP.t0 50.8339
R50 VP.n45 VP.n44 48.5829
R51 VP.n60 VP.n5 40.4934
R52 VP.n64 VP.n5 40.4934
R53 VP.n28 VP.n17 40.4934
R54 VP.n24 VP.n17 40.4934
R55 VP.n49 VP.n9 25.9244
R56 VP.n73 VP.n1 25.9244
R57 VP.n37 VP.n13 25.9244
R58 VP.n48 VP.n47 24.4675
R59 VP.n49 VP.n48 24.4675
R60 VP.n54 VP.n53 24.4675
R61 VP.n55 VP.n54 24.4675
R62 VP.n59 VP.n58 24.4675
R63 VP.n60 VP.n59 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n67 VP.n65 24.4675
R66 VP.n71 VP.n3 24.4675
R67 VP.n72 VP.n71 24.4675
R68 VP.n77 VP.n1 24.4675
R69 VP.n78 VP.n77 24.4675
R70 VP.n41 VP.n13 24.4675
R71 VP.n42 VP.n41 24.4675
R72 VP.n29 VP.n28 24.4675
R73 VP.n31 VP.n29 24.4675
R74 VP.n35 VP.n15 24.4675
R75 VP.n36 VP.n35 24.4675
R76 VP.n23 VP.n22 24.4675
R77 VP.n24 VP.n23 24.4675
R78 VP.n55 VP.n7 15.9041
R79 VP.n66 VP.n3 15.9041
R80 VP.n30 VP.n15 15.9041
R81 VP.n58 VP.n7 8.56395
R82 VP.n67 VP.n66 8.56395
R83 VP.n31 VP.n30 8.56395
R84 VP.n22 VP.n19 8.56395
R85 VP.n21 VP.n20 5.17456
R86 VP.n47 VP.n11 1.22385
R87 VP.n79 VP.n78 1.22385
R88 VP.n43 VP.n42 1.22385
R89 VP.n44 VP.n12 0.278367
R90 VP.n46 VP.n45 0.278367
R91 VP.n80 VP.n0 0.278367
R92 VP.n21 VP.n18 0.189894
R93 VP.n25 VP.n18 0.189894
R94 VP.n26 VP.n25 0.189894
R95 VP.n27 VP.n26 0.189894
R96 VP.n27 VP.n16 0.189894
R97 VP.n32 VP.n16 0.189894
R98 VP.n33 VP.n32 0.189894
R99 VP.n34 VP.n33 0.189894
R100 VP.n34 VP.n14 0.189894
R101 VP.n38 VP.n14 0.189894
R102 VP.n39 VP.n38 0.189894
R103 VP.n40 VP.n39 0.189894
R104 VP.n40 VP.n12 0.189894
R105 VP.n46 VP.n10 0.189894
R106 VP.n50 VP.n10 0.189894
R107 VP.n51 VP.n50 0.189894
R108 VP.n52 VP.n51 0.189894
R109 VP.n52 VP.n8 0.189894
R110 VP.n56 VP.n8 0.189894
R111 VP.n57 VP.n56 0.189894
R112 VP.n57 VP.n6 0.189894
R113 VP.n61 VP.n6 0.189894
R114 VP.n62 VP.n61 0.189894
R115 VP.n63 VP.n62 0.189894
R116 VP.n63 VP.n4 0.189894
R117 VP.n68 VP.n4 0.189894
R118 VP.n69 VP.n68 0.189894
R119 VP.n70 VP.n69 0.189894
R120 VP.n70 VP.n2 0.189894
R121 VP.n74 VP.n2 0.189894
R122 VP.n75 VP.n74 0.189894
R123 VP.n76 VP.n75 0.189894
R124 VP.n76 VP.n0 0.189894
R125 VP VP.n80 0.153454
R126 VTAIL.n11 VTAIL.t11 53.2195
R127 VTAIL.n10 VTAIL.t0 53.2195
R128 VTAIL.n7 VTAIL.t4 53.2195
R129 VTAIL.n15 VTAIL.t7 53.2194
R130 VTAIL.n2 VTAIL.t3 53.2194
R131 VTAIL.n3 VTAIL.t9 53.2194
R132 VTAIL.n6 VTAIL.t15 53.2194
R133 VTAIL.n14 VTAIL.t10 53.2194
R134 VTAIL.n13 VTAIL.n12 50.1112
R135 VTAIL.n9 VTAIL.n8 50.1112
R136 VTAIL.n1 VTAIL.n0 50.111
R137 VTAIL.n5 VTAIL.n4 50.111
R138 VTAIL.n15 VTAIL.n14 20.7462
R139 VTAIL.n7 VTAIL.n6 20.7462
R140 VTAIL.n0 VTAIL.t6 3.10882
R141 VTAIL.n0 VTAIL.t2 3.10882
R142 VTAIL.n4 VTAIL.t8 3.10882
R143 VTAIL.n4 VTAIL.t13 3.10882
R144 VTAIL.n12 VTAIL.t12 3.10882
R145 VTAIL.n12 VTAIL.t14 3.10882
R146 VTAIL.n8 VTAIL.t5 3.10882
R147 VTAIL.n8 VTAIL.t1 3.10882
R148 VTAIL.n9 VTAIL.n7 2.88843
R149 VTAIL.n10 VTAIL.n9 2.88843
R150 VTAIL.n13 VTAIL.n11 2.88843
R151 VTAIL.n14 VTAIL.n13 2.88843
R152 VTAIL.n6 VTAIL.n5 2.88843
R153 VTAIL.n5 VTAIL.n3 2.88843
R154 VTAIL.n2 VTAIL.n1 2.88843
R155 VTAIL VTAIL.n15 2.83024
R156 VTAIL.n11 VTAIL.n10 0.470328
R157 VTAIL.n3 VTAIL.n2 0.470328
R158 VTAIL VTAIL.n1 0.0586897
R159 VDD1 VDD1.n0 68.2921
R160 VDD1.n3 VDD1.n2 68.1784
R161 VDD1.n3 VDD1.n1 68.1784
R162 VDD1.n5 VDD1.n4 66.7898
R163 VDD1.n5 VDD1.n3 42.7854
R164 VDD1.n4 VDD1.t6 3.10882
R165 VDD1.n4 VDD1.t1 3.10882
R166 VDD1.n0 VDD1.t5 3.10882
R167 VDD1.n0 VDD1.t7 3.10882
R168 VDD1.n2 VDD1.t0 3.10882
R169 VDD1.n2 VDD1.t2 3.10882
R170 VDD1.n1 VDD1.t4 3.10882
R171 VDD1.n1 VDD1.t3 3.10882
R172 VDD1 VDD1.n5 1.38628
R173 B.n772 B.n771 585
R174 B.n258 B.n135 585
R175 B.n257 B.n256 585
R176 B.n255 B.n254 585
R177 B.n253 B.n252 585
R178 B.n251 B.n250 585
R179 B.n249 B.n248 585
R180 B.n247 B.n246 585
R181 B.n245 B.n244 585
R182 B.n243 B.n242 585
R183 B.n241 B.n240 585
R184 B.n239 B.n238 585
R185 B.n237 B.n236 585
R186 B.n235 B.n234 585
R187 B.n233 B.n232 585
R188 B.n231 B.n230 585
R189 B.n229 B.n228 585
R190 B.n227 B.n226 585
R191 B.n225 B.n224 585
R192 B.n223 B.n222 585
R193 B.n221 B.n220 585
R194 B.n219 B.n218 585
R195 B.n217 B.n216 585
R196 B.n215 B.n214 585
R197 B.n213 B.n212 585
R198 B.n210 B.n209 585
R199 B.n208 B.n207 585
R200 B.n206 B.n205 585
R201 B.n204 B.n203 585
R202 B.n202 B.n201 585
R203 B.n200 B.n199 585
R204 B.n198 B.n197 585
R205 B.n196 B.n195 585
R206 B.n194 B.n193 585
R207 B.n192 B.n191 585
R208 B.n189 B.n188 585
R209 B.n187 B.n186 585
R210 B.n185 B.n184 585
R211 B.n183 B.n182 585
R212 B.n181 B.n180 585
R213 B.n179 B.n178 585
R214 B.n177 B.n176 585
R215 B.n175 B.n174 585
R216 B.n173 B.n172 585
R217 B.n171 B.n170 585
R218 B.n169 B.n168 585
R219 B.n167 B.n166 585
R220 B.n165 B.n164 585
R221 B.n163 B.n162 585
R222 B.n161 B.n160 585
R223 B.n159 B.n158 585
R224 B.n157 B.n156 585
R225 B.n155 B.n154 585
R226 B.n153 B.n152 585
R227 B.n151 B.n150 585
R228 B.n149 B.n148 585
R229 B.n147 B.n146 585
R230 B.n145 B.n144 585
R231 B.n143 B.n142 585
R232 B.n141 B.n140 585
R233 B.n770 B.n105 585
R234 B.n775 B.n105 585
R235 B.n769 B.n104 585
R236 B.n776 B.n104 585
R237 B.n768 B.n767 585
R238 B.n767 B.n100 585
R239 B.n766 B.n99 585
R240 B.n782 B.n99 585
R241 B.n765 B.n98 585
R242 B.n783 B.n98 585
R243 B.n764 B.n97 585
R244 B.n784 B.n97 585
R245 B.n763 B.n762 585
R246 B.n762 B.n93 585
R247 B.n761 B.n92 585
R248 B.n790 B.n92 585
R249 B.n760 B.n91 585
R250 B.n791 B.n91 585
R251 B.n759 B.n90 585
R252 B.n792 B.n90 585
R253 B.n758 B.n757 585
R254 B.n757 B.n86 585
R255 B.n756 B.n85 585
R256 B.n798 B.n85 585
R257 B.n755 B.n84 585
R258 B.n799 B.n84 585
R259 B.n754 B.n83 585
R260 B.n800 B.n83 585
R261 B.n753 B.n752 585
R262 B.n752 B.n79 585
R263 B.n751 B.n78 585
R264 B.n806 B.n78 585
R265 B.n750 B.n77 585
R266 B.n807 B.n77 585
R267 B.n749 B.n76 585
R268 B.n808 B.n76 585
R269 B.n748 B.n747 585
R270 B.n747 B.n72 585
R271 B.n746 B.n71 585
R272 B.n814 B.n71 585
R273 B.n745 B.n70 585
R274 B.n815 B.n70 585
R275 B.n744 B.n69 585
R276 B.n816 B.n69 585
R277 B.n743 B.n742 585
R278 B.n742 B.n65 585
R279 B.n741 B.n64 585
R280 B.n822 B.n64 585
R281 B.n740 B.n63 585
R282 B.n823 B.n63 585
R283 B.n739 B.n62 585
R284 B.n824 B.n62 585
R285 B.n738 B.n737 585
R286 B.n737 B.n58 585
R287 B.n736 B.n57 585
R288 B.n830 B.n57 585
R289 B.n735 B.n56 585
R290 B.n831 B.n56 585
R291 B.n734 B.n55 585
R292 B.n832 B.n55 585
R293 B.n733 B.n732 585
R294 B.n732 B.n51 585
R295 B.n731 B.n50 585
R296 B.n838 B.n50 585
R297 B.n730 B.n49 585
R298 B.n839 B.n49 585
R299 B.n729 B.n48 585
R300 B.n840 B.n48 585
R301 B.n728 B.n727 585
R302 B.n727 B.n44 585
R303 B.n726 B.n43 585
R304 B.n846 B.n43 585
R305 B.n725 B.n42 585
R306 B.n847 B.n42 585
R307 B.n724 B.n41 585
R308 B.n848 B.n41 585
R309 B.n723 B.n722 585
R310 B.n722 B.n37 585
R311 B.n721 B.n36 585
R312 B.n854 B.n36 585
R313 B.n720 B.n35 585
R314 B.n855 B.n35 585
R315 B.n719 B.n34 585
R316 B.n856 B.n34 585
R317 B.n718 B.n717 585
R318 B.n717 B.n30 585
R319 B.n716 B.n29 585
R320 B.n862 B.n29 585
R321 B.n715 B.n28 585
R322 B.n863 B.n28 585
R323 B.n714 B.n27 585
R324 B.n864 B.n27 585
R325 B.n713 B.n712 585
R326 B.n712 B.n23 585
R327 B.n711 B.n22 585
R328 B.n870 B.n22 585
R329 B.n710 B.n21 585
R330 B.n871 B.n21 585
R331 B.n709 B.n20 585
R332 B.n872 B.n20 585
R333 B.n708 B.n707 585
R334 B.n707 B.n19 585
R335 B.n706 B.n15 585
R336 B.n878 B.n15 585
R337 B.n705 B.n14 585
R338 B.n879 B.n14 585
R339 B.n704 B.n13 585
R340 B.n880 B.n13 585
R341 B.n703 B.n702 585
R342 B.n702 B.n12 585
R343 B.n701 B.n700 585
R344 B.n701 B.n8 585
R345 B.n699 B.n7 585
R346 B.n887 B.n7 585
R347 B.n698 B.n6 585
R348 B.n888 B.n6 585
R349 B.n697 B.n5 585
R350 B.n889 B.n5 585
R351 B.n696 B.n695 585
R352 B.n695 B.n4 585
R353 B.n694 B.n259 585
R354 B.n694 B.n693 585
R355 B.n684 B.n260 585
R356 B.n261 B.n260 585
R357 B.n686 B.n685 585
R358 B.n687 B.n686 585
R359 B.n683 B.n266 585
R360 B.n266 B.n265 585
R361 B.n682 B.n681 585
R362 B.n681 B.n680 585
R363 B.n268 B.n267 585
R364 B.n673 B.n268 585
R365 B.n672 B.n671 585
R366 B.n674 B.n672 585
R367 B.n670 B.n273 585
R368 B.n273 B.n272 585
R369 B.n669 B.n668 585
R370 B.n668 B.n667 585
R371 B.n275 B.n274 585
R372 B.n276 B.n275 585
R373 B.n660 B.n659 585
R374 B.n661 B.n660 585
R375 B.n658 B.n281 585
R376 B.n281 B.n280 585
R377 B.n657 B.n656 585
R378 B.n656 B.n655 585
R379 B.n283 B.n282 585
R380 B.n284 B.n283 585
R381 B.n648 B.n647 585
R382 B.n649 B.n648 585
R383 B.n646 B.n289 585
R384 B.n289 B.n288 585
R385 B.n645 B.n644 585
R386 B.n644 B.n643 585
R387 B.n291 B.n290 585
R388 B.n292 B.n291 585
R389 B.n636 B.n635 585
R390 B.n637 B.n636 585
R391 B.n634 B.n297 585
R392 B.n297 B.n296 585
R393 B.n633 B.n632 585
R394 B.n632 B.n631 585
R395 B.n299 B.n298 585
R396 B.n300 B.n299 585
R397 B.n624 B.n623 585
R398 B.n625 B.n624 585
R399 B.n622 B.n305 585
R400 B.n305 B.n304 585
R401 B.n621 B.n620 585
R402 B.n620 B.n619 585
R403 B.n307 B.n306 585
R404 B.n308 B.n307 585
R405 B.n612 B.n611 585
R406 B.n613 B.n612 585
R407 B.n610 B.n313 585
R408 B.n313 B.n312 585
R409 B.n609 B.n608 585
R410 B.n608 B.n607 585
R411 B.n315 B.n314 585
R412 B.n316 B.n315 585
R413 B.n600 B.n599 585
R414 B.n601 B.n600 585
R415 B.n598 B.n321 585
R416 B.n321 B.n320 585
R417 B.n597 B.n596 585
R418 B.n596 B.n595 585
R419 B.n323 B.n322 585
R420 B.n324 B.n323 585
R421 B.n588 B.n587 585
R422 B.n589 B.n588 585
R423 B.n586 B.n329 585
R424 B.n329 B.n328 585
R425 B.n585 B.n584 585
R426 B.n584 B.n583 585
R427 B.n331 B.n330 585
R428 B.n332 B.n331 585
R429 B.n576 B.n575 585
R430 B.n577 B.n576 585
R431 B.n574 B.n337 585
R432 B.n337 B.n336 585
R433 B.n573 B.n572 585
R434 B.n572 B.n571 585
R435 B.n339 B.n338 585
R436 B.n340 B.n339 585
R437 B.n564 B.n563 585
R438 B.n565 B.n564 585
R439 B.n562 B.n345 585
R440 B.n345 B.n344 585
R441 B.n561 B.n560 585
R442 B.n560 B.n559 585
R443 B.n347 B.n346 585
R444 B.n348 B.n347 585
R445 B.n552 B.n551 585
R446 B.n553 B.n552 585
R447 B.n550 B.n352 585
R448 B.n356 B.n352 585
R449 B.n549 B.n548 585
R450 B.n548 B.n547 585
R451 B.n354 B.n353 585
R452 B.n355 B.n354 585
R453 B.n540 B.n539 585
R454 B.n541 B.n540 585
R455 B.n538 B.n361 585
R456 B.n361 B.n360 585
R457 B.n537 B.n536 585
R458 B.n536 B.n535 585
R459 B.n363 B.n362 585
R460 B.n364 B.n363 585
R461 B.n528 B.n527 585
R462 B.n529 B.n528 585
R463 B.n526 B.n369 585
R464 B.n369 B.n368 585
R465 B.n521 B.n520 585
R466 B.n519 B.n401 585
R467 B.n518 B.n400 585
R468 B.n523 B.n400 585
R469 B.n517 B.n516 585
R470 B.n515 B.n514 585
R471 B.n513 B.n512 585
R472 B.n511 B.n510 585
R473 B.n509 B.n508 585
R474 B.n507 B.n506 585
R475 B.n505 B.n504 585
R476 B.n503 B.n502 585
R477 B.n501 B.n500 585
R478 B.n499 B.n498 585
R479 B.n497 B.n496 585
R480 B.n495 B.n494 585
R481 B.n493 B.n492 585
R482 B.n491 B.n490 585
R483 B.n489 B.n488 585
R484 B.n487 B.n486 585
R485 B.n485 B.n484 585
R486 B.n483 B.n482 585
R487 B.n481 B.n480 585
R488 B.n479 B.n478 585
R489 B.n477 B.n476 585
R490 B.n475 B.n474 585
R491 B.n473 B.n472 585
R492 B.n471 B.n470 585
R493 B.n469 B.n468 585
R494 B.n467 B.n466 585
R495 B.n465 B.n464 585
R496 B.n463 B.n462 585
R497 B.n461 B.n460 585
R498 B.n459 B.n458 585
R499 B.n457 B.n456 585
R500 B.n455 B.n454 585
R501 B.n453 B.n452 585
R502 B.n451 B.n450 585
R503 B.n449 B.n448 585
R504 B.n447 B.n446 585
R505 B.n445 B.n444 585
R506 B.n443 B.n442 585
R507 B.n441 B.n440 585
R508 B.n439 B.n438 585
R509 B.n437 B.n436 585
R510 B.n435 B.n434 585
R511 B.n433 B.n432 585
R512 B.n431 B.n430 585
R513 B.n429 B.n428 585
R514 B.n427 B.n426 585
R515 B.n425 B.n424 585
R516 B.n423 B.n422 585
R517 B.n421 B.n420 585
R518 B.n419 B.n418 585
R519 B.n417 B.n416 585
R520 B.n415 B.n414 585
R521 B.n413 B.n412 585
R522 B.n411 B.n410 585
R523 B.n409 B.n408 585
R524 B.n371 B.n370 585
R525 B.n525 B.n524 585
R526 B.n524 B.n523 585
R527 B.n367 B.n366 585
R528 B.n368 B.n367 585
R529 B.n531 B.n530 585
R530 B.n530 B.n529 585
R531 B.n532 B.n365 585
R532 B.n365 B.n364 585
R533 B.n534 B.n533 585
R534 B.n535 B.n534 585
R535 B.n359 B.n358 585
R536 B.n360 B.n359 585
R537 B.n543 B.n542 585
R538 B.n542 B.n541 585
R539 B.n544 B.n357 585
R540 B.n357 B.n355 585
R541 B.n546 B.n545 585
R542 B.n547 B.n546 585
R543 B.n351 B.n350 585
R544 B.n356 B.n351 585
R545 B.n555 B.n554 585
R546 B.n554 B.n553 585
R547 B.n556 B.n349 585
R548 B.n349 B.n348 585
R549 B.n558 B.n557 585
R550 B.n559 B.n558 585
R551 B.n343 B.n342 585
R552 B.n344 B.n343 585
R553 B.n567 B.n566 585
R554 B.n566 B.n565 585
R555 B.n568 B.n341 585
R556 B.n341 B.n340 585
R557 B.n570 B.n569 585
R558 B.n571 B.n570 585
R559 B.n335 B.n334 585
R560 B.n336 B.n335 585
R561 B.n579 B.n578 585
R562 B.n578 B.n577 585
R563 B.n580 B.n333 585
R564 B.n333 B.n332 585
R565 B.n582 B.n581 585
R566 B.n583 B.n582 585
R567 B.n327 B.n326 585
R568 B.n328 B.n327 585
R569 B.n591 B.n590 585
R570 B.n590 B.n589 585
R571 B.n592 B.n325 585
R572 B.n325 B.n324 585
R573 B.n594 B.n593 585
R574 B.n595 B.n594 585
R575 B.n319 B.n318 585
R576 B.n320 B.n319 585
R577 B.n603 B.n602 585
R578 B.n602 B.n601 585
R579 B.n604 B.n317 585
R580 B.n317 B.n316 585
R581 B.n606 B.n605 585
R582 B.n607 B.n606 585
R583 B.n311 B.n310 585
R584 B.n312 B.n311 585
R585 B.n615 B.n614 585
R586 B.n614 B.n613 585
R587 B.n616 B.n309 585
R588 B.n309 B.n308 585
R589 B.n618 B.n617 585
R590 B.n619 B.n618 585
R591 B.n303 B.n302 585
R592 B.n304 B.n303 585
R593 B.n627 B.n626 585
R594 B.n626 B.n625 585
R595 B.n628 B.n301 585
R596 B.n301 B.n300 585
R597 B.n630 B.n629 585
R598 B.n631 B.n630 585
R599 B.n295 B.n294 585
R600 B.n296 B.n295 585
R601 B.n639 B.n638 585
R602 B.n638 B.n637 585
R603 B.n640 B.n293 585
R604 B.n293 B.n292 585
R605 B.n642 B.n641 585
R606 B.n643 B.n642 585
R607 B.n287 B.n286 585
R608 B.n288 B.n287 585
R609 B.n651 B.n650 585
R610 B.n650 B.n649 585
R611 B.n652 B.n285 585
R612 B.n285 B.n284 585
R613 B.n654 B.n653 585
R614 B.n655 B.n654 585
R615 B.n279 B.n278 585
R616 B.n280 B.n279 585
R617 B.n663 B.n662 585
R618 B.n662 B.n661 585
R619 B.n664 B.n277 585
R620 B.n277 B.n276 585
R621 B.n666 B.n665 585
R622 B.n667 B.n666 585
R623 B.n271 B.n270 585
R624 B.n272 B.n271 585
R625 B.n676 B.n675 585
R626 B.n675 B.n674 585
R627 B.n677 B.n269 585
R628 B.n673 B.n269 585
R629 B.n679 B.n678 585
R630 B.n680 B.n679 585
R631 B.n264 B.n263 585
R632 B.n265 B.n264 585
R633 B.n689 B.n688 585
R634 B.n688 B.n687 585
R635 B.n690 B.n262 585
R636 B.n262 B.n261 585
R637 B.n692 B.n691 585
R638 B.n693 B.n692 585
R639 B.n3 B.n0 585
R640 B.n4 B.n3 585
R641 B.n886 B.n1 585
R642 B.n887 B.n886 585
R643 B.n885 B.n884 585
R644 B.n885 B.n8 585
R645 B.n883 B.n9 585
R646 B.n12 B.n9 585
R647 B.n882 B.n881 585
R648 B.n881 B.n880 585
R649 B.n11 B.n10 585
R650 B.n879 B.n11 585
R651 B.n877 B.n876 585
R652 B.n878 B.n877 585
R653 B.n875 B.n16 585
R654 B.n19 B.n16 585
R655 B.n874 B.n873 585
R656 B.n873 B.n872 585
R657 B.n18 B.n17 585
R658 B.n871 B.n18 585
R659 B.n869 B.n868 585
R660 B.n870 B.n869 585
R661 B.n867 B.n24 585
R662 B.n24 B.n23 585
R663 B.n866 B.n865 585
R664 B.n865 B.n864 585
R665 B.n26 B.n25 585
R666 B.n863 B.n26 585
R667 B.n861 B.n860 585
R668 B.n862 B.n861 585
R669 B.n859 B.n31 585
R670 B.n31 B.n30 585
R671 B.n858 B.n857 585
R672 B.n857 B.n856 585
R673 B.n33 B.n32 585
R674 B.n855 B.n33 585
R675 B.n853 B.n852 585
R676 B.n854 B.n853 585
R677 B.n851 B.n38 585
R678 B.n38 B.n37 585
R679 B.n850 B.n849 585
R680 B.n849 B.n848 585
R681 B.n40 B.n39 585
R682 B.n847 B.n40 585
R683 B.n845 B.n844 585
R684 B.n846 B.n845 585
R685 B.n843 B.n45 585
R686 B.n45 B.n44 585
R687 B.n842 B.n841 585
R688 B.n841 B.n840 585
R689 B.n47 B.n46 585
R690 B.n839 B.n47 585
R691 B.n837 B.n836 585
R692 B.n838 B.n837 585
R693 B.n835 B.n52 585
R694 B.n52 B.n51 585
R695 B.n834 B.n833 585
R696 B.n833 B.n832 585
R697 B.n54 B.n53 585
R698 B.n831 B.n54 585
R699 B.n829 B.n828 585
R700 B.n830 B.n829 585
R701 B.n827 B.n59 585
R702 B.n59 B.n58 585
R703 B.n826 B.n825 585
R704 B.n825 B.n824 585
R705 B.n61 B.n60 585
R706 B.n823 B.n61 585
R707 B.n821 B.n820 585
R708 B.n822 B.n821 585
R709 B.n819 B.n66 585
R710 B.n66 B.n65 585
R711 B.n818 B.n817 585
R712 B.n817 B.n816 585
R713 B.n68 B.n67 585
R714 B.n815 B.n68 585
R715 B.n813 B.n812 585
R716 B.n814 B.n813 585
R717 B.n811 B.n73 585
R718 B.n73 B.n72 585
R719 B.n810 B.n809 585
R720 B.n809 B.n808 585
R721 B.n75 B.n74 585
R722 B.n807 B.n75 585
R723 B.n805 B.n804 585
R724 B.n806 B.n805 585
R725 B.n803 B.n80 585
R726 B.n80 B.n79 585
R727 B.n802 B.n801 585
R728 B.n801 B.n800 585
R729 B.n82 B.n81 585
R730 B.n799 B.n82 585
R731 B.n797 B.n796 585
R732 B.n798 B.n797 585
R733 B.n795 B.n87 585
R734 B.n87 B.n86 585
R735 B.n794 B.n793 585
R736 B.n793 B.n792 585
R737 B.n89 B.n88 585
R738 B.n791 B.n89 585
R739 B.n789 B.n788 585
R740 B.n790 B.n789 585
R741 B.n787 B.n94 585
R742 B.n94 B.n93 585
R743 B.n786 B.n785 585
R744 B.n785 B.n784 585
R745 B.n96 B.n95 585
R746 B.n783 B.n96 585
R747 B.n781 B.n780 585
R748 B.n782 B.n781 585
R749 B.n779 B.n101 585
R750 B.n101 B.n100 585
R751 B.n778 B.n777 585
R752 B.n777 B.n776 585
R753 B.n103 B.n102 585
R754 B.n775 B.n103 585
R755 B.n890 B.n889 585
R756 B.n888 B.n2 585
R757 B.n140 B.n103 454.062
R758 B.n772 B.n105 454.062
R759 B.n524 B.n369 454.062
R760 B.n521 B.n367 454.062
R761 B.n138 B.t8 259.438
R762 B.n136 B.t19 259.438
R763 B.n405 B.t12 259.438
R764 B.n402 B.t16 259.438
R765 B.n774 B.n773 256.663
R766 B.n774 B.n134 256.663
R767 B.n774 B.n133 256.663
R768 B.n774 B.n132 256.663
R769 B.n774 B.n131 256.663
R770 B.n774 B.n130 256.663
R771 B.n774 B.n129 256.663
R772 B.n774 B.n128 256.663
R773 B.n774 B.n127 256.663
R774 B.n774 B.n126 256.663
R775 B.n774 B.n125 256.663
R776 B.n774 B.n124 256.663
R777 B.n774 B.n123 256.663
R778 B.n774 B.n122 256.663
R779 B.n774 B.n121 256.663
R780 B.n774 B.n120 256.663
R781 B.n774 B.n119 256.663
R782 B.n774 B.n118 256.663
R783 B.n774 B.n117 256.663
R784 B.n774 B.n116 256.663
R785 B.n774 B.n115 256.663
R786 B.n774 B.n114 256.663
R787 B.n774 B.n113 256.663
R788 B.n774 B.n112 256.663
R789 B.n774 B.n111 256.663
R790 B.n774 B.n110 256.663
R791 B.n774 B.n109 256.663
R792 B.n774 B.n108 256.663
R793 B.n774 B.n107 256.663
R794 B.n774 B.n106 256.663
R795 B.n523 B.n522 256.663
R796 B.n523 B.n372 256.663
R797 B.n523 B.n373 256.663
R798 B.n523 B.n374 256.663
R799 B.n523 B.n375 256.663
R800 B.n523 B.n376 256.663
R801 B.n523 B.n377 256.663
R802 B.n523 B.n378 256.663
R803 B.n523 B.n379 256.663
R804 B.n523 B.n380 256.663
R805 B.n523 B.n381 256.663
R806 B.n523 B.n382 256.663
R807 B.n523 B.n383 256.663
R808 B.n523 B.n384 256.663
R809 B.n523 B.n385 256.663
R810 B.n523 B.n386 256.663
R811 B.n523 B.n387 256.663
R812 B.n523 B.n388 256.663
R813 B.n523 B.n389 256.663
R814 B.n523 B.n390 256.663
R815 B.n523 B.n391 256.663
R816 B.n523 B.n392 256.663
R817 B.n523 B.n393 256.663
R818 B.n523 B.n394 256.663
R819 B.n523 B.n395 256.663
R820 B.n523 B.n396 256.663
R821 B.n523 B.n397 256.663
R822 B.n523 B.n398 256.663
R823 B.n523 B.n399 256.663
R824 B.n892 B.n891 256.663
R825 B.n144 B.n143 163.367
R826 B.n148 B.n147 163.367
R827 B.n152 B.n151 163.367
R828 B.n156 B.n155 163.367
R829 B.n160 B.n159 163.367
R830 B.n164 B.n163 163.367
R831 B.n168 B.n167 163.367
R832 B.n172 B.n171 163.367
R833 B.n176 B.n175 163.367
R834 B.n180 B.n179 163.367
R835 B.n184 B.n183 163.367
R836 B.n188 B.n187 163.367
R837 B.n193 B.n192 163.367
R838 B.n197 B.n196 163.367
R839 B.n201 B.n200 163.367
R840 B.n205 B.n204 163.367
R841 B.n209 B.n208 163.367
R842 B.n214 B.n213 163.367
R843 B.n218 B.n217 163.367
R844 B.n222 B.n221 163.367
R845 B.n226 B.n225 163.367
R846 B.n230 B.n229 163.367
R847 B.n234 B.n233 163.367
R848 B.n238 B.n237 163.367
R849 B.n242 B.n241 163.367
R850 B.n246 B.n245 163.367
R851 B.n250 B.n249 163.367
R852 B.n254 B.n253 163.367
R853 B.n256 B.n135 163.367
R854 B.n528 B.n369 163.367
R855 B.n528 B.n363 163.367
R856 B.n536 B.n363 163.367
R857 B.n536 B.n361 163.367
R858 B.n540 B.n361 163.367
R859 B.n540 B.n354 163.367
R860 B.n548 B.n354 163.367
R861 B.n548 B.n352 163.367
R862 B.n552 B.n352 163.367
R863 B.n552 B.n347 163.367
R864 B.n560 B.n347 163.367
R865 B.n560 B.n345 163.367
R866 B.n564 B.n345 163.367
R867 B.n564 B.n339 163.367
R868 B.n572 B.n339 163.367
R869 B.n572 B.n337 163.367
R870 B.n576 B.n337 163.367
R871 B.n576 B.n331 163.367
R872 B.n584 B.n331 163.367
R873 B.n584 B.n329 163.367
R874 B.n588 B.n329 163.367
R875 B.n588 B.n323 163.367
R876 B.n596 B.n323 163.367
R877 B.n596 B.n321 163.367
R878 B.n600 B.n321 163.367
R879 B.n600 B.n315 163.367
R880 B.n608 B.n315 163.367
R881 B.n608 B.n313 163.367
R882 B.n612 B.n313 163.367
R883 B.n612 B.n307 163.367
R884 B.n620 B.n307 163.367
R885 B.n620 B.n305 163.367
R886 B.n624 B.n305 163.367
R887 B.n624 B.n299 163.367
R888 B.n632 B.n299 163.367
R889 B.n632 B.n297 163.367
R890 B.n636 B.n297 163.367
R891 B.n636 B.n291 163.367
R892 B.n644 B.n291 163.367
R893 B.n644 B.n289 163.367
R894 B.n648 B.n289 163.367
R895 B.n648 B.n283 163.367
R896 B.n656 B.n283 163.367
R897 B.n656 B.n281 163.367
R898 B.n660 B.n281 163.367
R899 B.n660 B.n275 163.367
R900 B.n668 B.n275 163.367
R901 B.n668 B.n273 163.367
R902 B.n672 B.n273 163.367
R903 B.n672 B.n268 163.367
R904 B.n681 B.n268 163.367
R905 B.n681 B.n266 163.367
R906 B.n686 B.n266 163.367
R907 B.n686 B.n260 163.367
R908 B.n694 B.n260 163.367
R909 B.n695 B.n694 163.367
R910 B.n695 B.n5 163.367
R911 B.n6 B.n5 163.367
R912 B.n7 B.n6 163.367
R913 B.n701 B.n7 163.367
R914 B.n702 B.n701 163.367
R915 B.n702 B.n13 163.367
R916 B.n14 B.n13 163.367
R917 B.n15 B.n14 163.367
R918 B.n707 B.n15 163.367
R919 B.n707 B.n20 163.367
R920 B.n21 B.n20 163.367
R921 B.n22 B.n21 163.367
R922 B.n712 B.n22 163.367
R923 B.n712 B.n27 163.367
R924 B.n28 B.n27 163.367
R925 B.n29 B.n28 163.367
R926 B.n717 B.n29 163.367
R927 B.n717 B.n34 163.367
R928 B.n35 B.n34 163.367
R929 B.n36 B.n35 163.367
R930 B.n722 B.n36 163.367
R931 B.n722 B.n41 163.367
R932 B.n42 B.n41 163.367
R933 B.n43 B.n42 163.367
R934 B.n727 B.n43 163.367
R935 B.n727 B.n48 163.367
R936 B.n49 B.n48 163.367
R937 B.n50 B.n49 163.367
R938 B.n732 B.n50 163.367
R939 B.n732 B.n55 163.367
R940 B.n56 B.n55 163.367
R941 B.n57 B.n56 163.367
R942 B.n737 B.n57 163.367
R943 B.n737 B.n62 163.367
R944 B.n63 B.n62 163.367
R945 B.n64 B.n63 163.367
R946 B.n742 B.n64 163.367
R947 B.n742 B.n69 163.367
R948 B.n70 B.n69 163.367
R949 B.n71 B.n70 163.367
R950 B.n747 B.n71 163.367
R951 B.n747 B.n76 163.367
R952 B.n77 B.n76 163.367
R953 B.n78 B.n77 163.367
R954 B.n752 B.n78 163.367
R955 B.n752 B.n83 163.367
R956 B.n84 B.n83 163.367
R957 B.n85 B.n84 163.367
R958 B.n757 B.n85 163.367
R959 B.n757 B.n90 163.367
R960 B.n91 B.n90 163.367
R961 B.n92 B.n91 163.367
R962 B.n762 B.n92 163.367
R963 B.n762 B.n97 163.367
R964 B.n98 B.n97 163.367
R965 B.n99 B.n98 163.367
R966 B.n767 B.n99 163.367
R967 B.n767 B.n104 163.367
R968 B.n105 B.n104 163.367
R969 B.n401 B.n400 163.367
R970 B.n516 B.n400 163.367
R971 B.n514 B.n513 163.367
R972 B.n510 B.n509 163.367
R973 B.n506 B.n505 163.367
R974 B.n502 B.n501 163.367
R975 B.n498 B.n497 163.367
R976 B.n494 B.n493 163.367
R977 B.n490 B.n489 163.367
R978 B.n486 B.n485 163.367
R979 B.n482 B.n481 163.367
R980 B.n478 B.n477 163.367
R981 B.n474 B.n473 163.367
R982 B.n470 B.n469 163.367
R983 B.n466 B.n465 163.367
R984 B.n462 B.n461 163.367
R985 B.n458 B.n457 163.367
R986 B.n454 B.n453 163.367
R987 B.n450 B.n449 163.367
R988 B.n446 B.n445 163.367
R989 B.n442 B.n441 163.367
R990 B.n438 B.n437 163.367
R991 B.n434 B.n433 163.367
R992 B.n430 B.n429 163.367
R993 B.n426 B.n425 163.367
R994 B.n422 B.n421 163.367
R995 B.n418 B.n417 163.367
R996 B.n414 B.n413 163.367
R997 B.n410 B.n409 163.367
R998 B.n524 B.n371 163.367
R999 B.n530 B.n367 163.367
R1000 B.n530 B.n365 163.367
R1001 B.n534 B.n365 163.367
R1002 B.n534 B.n359 163.367
R1003 B.n542 B.n359 163.367
R1004 B.n542 B.n357 163.367
R1005 B.n546 B.n357 163.367
R1006 B.n546 B.n351 163.367
R1007 B.n554 B.n351 163.367
R1008 B.n554 B.n349 163.367
R1009 B.n558 B.n349 163.367
R1010 B.n558 B.n343 163.367
R1011 B.n566 B.n343 163.367
R1012 B.n566 B.n341 163.367
R1013 B.n570 B.n341 163.367
R1014 B.n570 B.n335 163.367
R1015 B.n578 B.n335 163.367
R1016 B.n578 B.n333 163.367
R1017 B.n582 B.n333 163.367
R1018 B.n582 B.n327 163.367
R1019 B.n590 B.n327 163.367
R1020 B.n590 B.n325 163.367
R1021 B.n594 B.n325 163.367
R1022 B.n594 B.n319 163.367
R1023 B.n602 B.n319 163.367
R1024 B.n602 B.n317 163.367
R1025 B.n606 B.n317 163.367
R1026 B.n606 B.n311 163.367
R1027 B.n614 B.n311 163.367
R1028 B.n614 B.n309 163.367
R1029 B.n618 B.n309 163.367
R1030 B.n618 B.n303 163.367
R1031 B.n626 B.n303 163.367
R1032 B.n626 B.n301 163.367
R1033 B.n630 B.n301 163.367
R1034 B.n630 B.n295 163.367
R1035 B.n638 B.n295 163.367
R1036 B.n638 B.n293 163.367
R1037 B.n642 B.n293 163.367
R1038 B.n642 B.n287 163.367
R1039 B.n650 B.n287 163.367
R1040 B.n650 B.n285 163.367
R1041 B.n654 B.n285 163.367
R1042 B.n654 B.n279 163.367
R1043 B.n662 B.n279 163.367
R1044 B.n662 B.n277 163.367
R1045 B.n666 B.n277 163.367
R1046 B.n666 B.n271 163.367
R1047 B.n675 B.n271 163.367
R1048 B.n675 B.n269 163.367
R1049 B.n679 B.n269 163.367
R1050 B.n679 B.n264 163.367
R1051 B.n688 B.n264 163.367
R1052 B.n688 B.n262 163.367
R1053 B.n692 B.n262 163.367
R1054 B.n692 B.n3 163.367
R1055 B.n890 B.n3 163.367
R1056 B.n886 B.n2 163.367
R1057 B.n886 B.n885 163.367
R1058 B.n885 B.n9 163.367
R1059 B.n881 B.n9 163.367
R1060 B.n881 B.n11 163.367
R1061 B.n877 B.n11 163.367
R1062 B.n877 B.n16 163.367
R1063 B.n873 B.n16 163.367
R1064 B.n873 B.n18 163.367
R1065 B.n869 B.n18 163.367
R1066 B.n869 B.n24 163.367
R1067 B.n865 B.n24 163.367
R1068 B.n865 B.n26 163.367
R1069 B.n861 B.n26 163.367
R1070 B.n861 B.n31 163.367
R1071 B.n857 B.n31 163.367
R1072 B.n857 B.n33 163.367
R1073 B.n853 B.n33 163.367
R1074 B.n853 B.n38 163.367
R1075 B.n849 B.n38 163.367
R1076 B.n849 B.n40 163.367
R1077 B.n845 B.n40 163.367
R1078 B.n845 B.n45 163.367
R1079 B.n841 B.n45 163.367
R1080 B.n841 B.n47 163.367
R1081 B.n837 B.n47 163.367
R1082 B.n837 B.n52 163.367
R1083 B.n833 B.n52 163.367
R1084 B.n833 B.n54 163.367
R1085 B.n829 B.n54 163.367
R1086 B.n829 B.n59 163.367
R1087 B.n825 B.n59 163.367
R1088 B.n825 B.n61 163.367
R1089 B.n821 B.n61 163.367
R1090 B.n821 B.n66 163.367
R1091 B.n817 B.n66 163.367
R1092 B.n817 B.n68 163.367
R1093 B.n813 B.n68 163.367
R1094 B.n813 B.n73 163.367
R1095 B.n809 B.n73 163.367
R1096 B.n809 B.n75 163.367
R1097 B.n805 B.n75 163.367
R1098 B.n805 B.n80 163.367
R1099 B.n801 B.n80 163.367
R1100 B.n801 B.n82 163.367
R1101 B.n797 B.n82 163.367
R1102 B.n797 B.n87 163.367
R1103 B.n793 B.n87 163.367
R1104 B.n793 B.n89 163.367
R1105 B.n789 B.n89 163.367
R1106 B.n789 B.n94 163.367
R1107 B.n785 B.n94 163.367
R1108 B.n785 B.n96 163.367
R1109 B.n781 B.n96 163.367
R1110 B.n781 B.n101 163.367
R1111 B.n777 B.n101 163.367
R1112 B.n777 B.n103 163.367
R1113 B.n136 B.t20 139.07
R1114 B.n405 B.t15 139.07
R1115 B.n138 B.t10 139.062
R1116 B.n402 B.t18 139.062
R1117 B.n523 B.n368 108.63
R1118 B.n775 B.n774 108.63
R1119 B.n137 B.t21 74.0999
R1120 B.n406 B.t14 74.0999
R1121 B.n139 B.t11 74.0932
R1122 B.n403 B.t17 74.0932
R1123 B.n140 B.n106 71.676
R1124 B.n144 B.n107 71.676
R1125 B.n148 B.n108 71.676
R1126 B.n152 B.n109 71.676
R1127 B.n156 B.n110 71.676
R1128 B.n160 B.n111 71.676
R1129 B.n164 B.n112 71.676
R1130 B.n168 B.n113 71.676
R1131 B.n172 B.n114 71.676
R1132 B.n176 B.n115 71.676
R1133 B.n180 B.n116 71.676
R1134 B.n184 B.n117 71.676
R1135 B.n188 B.n118 71.676
R1136 B.n193 B.n119 71.676
R1137 B.n197 B.n120 71.676
R1138 B.n201 B.n121 71.676
R1139 B.n205 B.n122 71.676
R1140 B.n209 B.n123 71.676
R1141 B.n214 B.n124 71.676
R1142 B.n218 B.n125 71.676
R1143 B.n222 B.n126 71.676
R1144 B.n226 B.n127 71.676
R1145 B.n230 B.n128 71.676
R1146 B.n234 B.n129 71.676
R1147 B.n238 B.n130 71.676
R1148 B.n242 B.n131 71.676
R1149 B.n246 B.n132 71.676
R1150 B.n250 B.n133 71.676
R1151 B.n254 B.n134 71.676
R1152 B.n773 B.n135 71.676
R1153 B.n773 B.n772 71.676
R1154 B.n256 B.n134 71.676
R1155 B.n253 B.n133 71.676
R1156 B.n249 B.n132 71.676
R1157 B.n245 B.n131 71.676
R1158 B.n241 B.n130 71.676
R1159 B.n237 B.n129 71.676
R1160 B.n233 B.n128 71.676
R1161 B.n229 B.n127 71.676
R1162 B.n225 B.n126 71.676
R1163 B.n221 B.n125 71.676
R1164 B.n217 B.n124 71.676
R1165 B.n213 B.n123 71.676
R1166 B.n208 B.n122 71.676
R1167 B.n204 B.n121 71.676
R1168 B.n200 B.n120 71.676
R1169 B.n196 B.n119 71.676
R1170 B.n192 B.n118 71.676
R1171 B.n187 B.n117 71.676
R1172 B.n183 B.n116 71.676
R1173 B.n179 B.n115 71.676
R1174 B.n175 B.n114 71.676
R1175 B.n171 B.n113 71.676
R1176 B.n167 B.n112 71.676
R1177 B.n163 B.n111 71.676
R1178 B.n159 B.n110 71.676
R1179 B.n155 B.n109 71.676
R1180 B.n151 B.n108 71.676
R1181 B.n147 B.n107 71.676
R1182 B.n143 B.n106 71.676
R1183 B.n522 B.n521 71.676
R1184 B.n516 B.n372 71.676
R1185 B.n513 B.n373 71.676
R1186 B.n509 B.n374 71.676
R1187 B.n505 B.n375 71.676
R1188 B.n501 B.n376 71.676
R1189 B.n497 B.n377 71.676
R1190 B.n493 B.n378 71.676
R1191 B.n489 B.n379 71.676
R1192 B.n485 B.n380 71.676
R1193 B.n481 B.n381 71.676
R1194 B.n477 B.n382 71.676
R1195 B.n473 B.n383 71.676
R1196 B.n469 B.n384 71.676
R1197 B.n465 B.n385 71.676
R1198 B.n461 B.n386 71.676
R1199 B.n457 B.n387 71.676
R1200 B.n453 B.n388 71.676
R1201 B.n449 B.n389 71.676
R1202 B.n445 B.n390 71.676
R1203 B.n441 B.n391 71.676
R1204 B.n437 B.n392 71.676
R1205 B.n433 B.n393 71.676
R1206 B.n429 B.n394 71.676
R1207 B.n425 B.n395 71.676
R1208 B.n421 B.n396 71.676
R1209 B.n417 B.n397 71.676
R1210 B.n413 B.n398 71.676
R1211 B.n409 B.n399 71.676
R1212 B.n522 B.n401 71.676
R1213 B.n514 B.n372 71.676
R1214 B.n510 B.n373 71.676
R1215 B.n506 B.n374 71.676
R1216 B.n502 B.n375 71.676
R1217 B.n498 B.n376 71.676
R1218 B.n494 B.n377 71.676
R1219 B.n490 B.n378 71.676
R1220 B.n486 B.n379 71.676
R1221 B.n482 B.n380 71.676
R1222 B.n478 B.n381 71.676
R1223 B.n474 B.n382 71.676
R1224 B.n470 B.n383 71.676
R1225 B.n466 B.n384 71.676
R1226 B.n462 B.n385 71.676
R1227 B.n458 B.n386 71.676
R1228 B.n454 B.n387 71.676
R1229 B.n450 B.n388 71.676
R1230 B.n446 B.n389 71.676
R1231 B.n442 B.n390 71.676
R1232 B.n438 B.n391 71.676
R1233 B.n434 B.n392 71.676
R1234 B.n430 B.n393 71.676
R1235 B.n426 B.n394 71.676
R1236 B.n422 B.n395 71.676
R1237 B.n418 B.n396 71.676
R1238 B.n414 B.n397 71.676
R1239 B.n410 B.n398 71.676
R1240 B.n399 B.n371 71.676
R1241 B.n891 B.n890 71.676
R1242 B.n891 B.n2 71.676
R1243 B.n139 B.n138 64.9702
R1244 B.n137 B.n136 64.9702
R1245 B.n406 B.n405 64.9702
R1246 B.n403 B.n402 64.9702
R1247 B.n529 B.n368 64.2341
R1248 B.n529 B.n364 64.2341
R1249 B.n535 B.n364 64.2341
R1250 B.n535 B.n360 64.2341
R1251 B.n541 B.n360 64.2341
R1252 B.n541 B.n355 64.2341
R1253 B.n547 B.n355 64.2341
R1254 B.n547 B.n356 64.2341
R1255 B.n553 B.n348 64.2341
R1256 B.n559 B.n348 64.2341
R1257 B.n559 B.n344 64.2341
R1258 B.n565 B.n344 64.2341
R1259 B.n565 B.n340 64.2341
R1260 B.n571 B.n340 64.2341
R1261 B.n571 B.n336 64.2341
R1262 B.n577 B.n336 64.2341
R1263 B.n577 B.n332 64.2341
R1264 B.n583 B.n332 64.2341
R1265 B.n583 B.n328 64.2341
R1266 B.n589 B.n328 64.2341
R1267 B.n595 B.n324 64.2341
R1268 B.n595 B.n320 64.2341
R1269 B.n601 B.n320 64.2341
R1270 B.n601 B.n316 64.2341
R1271 B.n607 B.n316 64.2341
R1272 B.n607 B.n312 64.2341
R1273 B.n613 B.n312 64.2341
R1274 B.n613 B.n308 64.2341
R1275 B.n619 B.n308 64.2341
R1276 B.n625 B.n304 64.2341
R1277 B.n625 B.n300 64.2341
R1278 B.n631 B.n300 64.2341
R1279 B.n631 B.n296 64.2341
R1280 B.n637 B.n296 64.2341
R1281 B.n637 B.n292 64.2341
R1282 B.n643 B.n292 64.2341
R1283 B.n643 B.n288 64.2341
R1284 B.n649 B.n288 64.2341
R1285 B.n655 B.n284 64.2341
R1286 B.n655 B.n280 64.2341
R1287 B.n661 B.n280 64.2341
R1288 B.n661 B.n276 64.2341
R1289 B.n667 B.n276 64.2341
R1290 B.n667 B.n272 64.2341
R1291 B.n674 B.n272 64.2341
R1292 B.n674 B.n673 64.2341
R1293 B.n680 B.n265 64.2341
R1294 B.n687 B.n265 64.2341
R1295 B.n687 B.n261 64.2341
R1296 B.n693 B.n261 64.2341
R1297 B.n693 B.n4 64.2341
R1298 B.n889 B.n4 64.2341
R1299 B.n889 B.n888 64.2341
R1300 B.n888 B.n887 64.2341
R1301 B.n887 B.n8 64.2341
R1302 B.n12 B.n8 64.2341
R1303 B.n880 B.n12 64.2341
R1304 B.n880 B.n879 64.2341
R1305 B.n879 B.n878 64.2341
R1306 B.n872 B.n19 64.2341
R1307 B.n872 B.n871 64.2341
R1308 B.n871 B.n870 64.2341
R1309 B.n870 B.n23 64.2341
R1310 B.n864 B.n23 64.2341
R1311 B.n864 B.n863 64.2341
R1312 B.n863 B.n862 64.2341
R1313 B.n862 B.n30 64.2341
R1314 B.n856 B.n855 64.2341
R1315 B.n855 B.n854 64.2341
R1316 B.n854 B.n37 64.2341
R1317 B.n848 B.n37 64.2341
R1318 B.n848 B.n847 64.2341
R1319 B.n847 B.n846 64.2341
R1320 B.n846 B.n44 64.2341
R1321 B.n840 B.n44 64.2341
R1322 B.n840 B.n839 64.2341
R1323 B.n838 B.n51 64.2341
R1324 B.n832 B.n51 64.2341
R1325 B.n832 B.n831 64.2341
R1326 B.n831 B.n830 64.2341
R1327 B.n830 B.n58 64.2341
R1328 B.n824 B.n58 64.2341
R1329 B.n824 B.n823 64.2341
R1330 B.n823 B.n822 64.2341
R1331 B.n822 B.n65 64.2341
R1332 B.n816 B.n815 64.2341
R1333 B.n815 B.n814 64.2341
R1334 B.n814 B.n72 64.2341
R1335 B.n808 B.n72 64.2341
R1336 B.n808 B.n807 64.2341
R1337 B.n807 B.n806 64.2341
R1338 B.n806 B.n79 64.2341
R1339 B.n800 B.n79 64.2341
R1340 B.n800 B.n799 64.2341
R1341 B.n799 B.n798 64.2341
R1342 B.n798 B.n86 64.2341
R1343 B.n792 B.n86 64.2341
R1344 B.n791 B.n790 64.2341
R1345 B.n790 B.n93 64.2341
R1346 B.n784 B.n93 64.2341
R1347 B.n784 B.n783 64.2341
R1348 B.n783 B.n782 64.2341
R1349 B.n782 B.n100 64.2341
R1350 B.n776 B.n100 64.2341
R1351 B.n776 B.n775 64.2341
R1352 B.n673 B.t0 62.3449
R1353 B.n19 B.t3 62.3449
R1354 B.n190 B.n139 59.5399
R1355 B.n211 B.n137 59.5399
R1356 B.n407 B.n406 59.5399
R1357 B.n404 B.n403 59.5399
R1358 B.t1 B.n284 56.6772
R1359 B.t6 B.n30 56.6772
R1360 B.t5 B.n304 47.2311
R1361 B.n839 B.t2 47.2311
R1362 B.n553 B.t13 41.5634
R1363 B.n792 B.t9 41.5634
R1364 B.t4 B.n324 37.785
R1365 B.t7 B.n65 37.785
R1366 B.n520 B.n366 29.5029
R1367 B.n526 B.n525 29.5029
R1368 B.n771 B.n770 29.5029
R1369 B.n141 B.n102 29.5029
R1370 B.n589 B.t4 26.4496
R1371 B.n816 B.t7 26.4496
R1372 B.n356 B.t13 22.6712
R1373 B.t9 B.n791 22.6712
R1374 B B.n892 18.0485
R1375 B.n619 B.t5 17.0035
R1376 B.t2 B.n838 17.0035
R1377 B.n531 B.n366 10.6151
R1378 B.n532 B.n531 10.6151
R1379 B.n533 B.n532 10.6151
R1380 B.n533 B.n358 10.6151
R1381 B.n543 B.n358 10.6151
R1382 B.n544 B.n543 10.6151
R1383 B.n545 B.n544 10.6151
R1384 B.n545 B.n350 10.6151
R1385 B.n555 B.n350 10.6151
R1386 B.n556 B.n555 10.6151
R1387 B.n557 B.n556 10.6151
R1388 B.n557 B.n342 10.6151
R1389 B.n567 B.n342 10.6151
R1390 B.n568 B.n567 10.6151
R1391 B.n569 B.n568 10.6151
R1392 B.n569 B.n334 10.6151
R1393 B.n579 B.n334 10.6151
R1394 B.n580 B.n579 10.6151
R1395 B.n581 B.n580 10.6151
R1396 B.n581 B.n326 10.6151
R1397 B.n591 B.n326 10.6151
R1398 B.n592 B.n591 10.6151
R1399 B.n593 B.n592 10.6151
R1400 B.n593 B.n318 10.6151
R1401 B.n603 B.n318 10.6151
R1402 B.n604 B.n603 10.6151
R1403 B.n605 B.n604 10.6151
R1404 B.n605 B.n310 10.6151
R1405 B.n615 B.n310 10.6151
R1406 B.n616 B.n615 10.6151
R1407 B.n617 B.n616 10.6151
R1408 B.n617 B.n302 10.6151
R1409 B.n627 B.n302 10.6151
R1410 B.n628 B.n627 10.6151
R1411 B.n629 B.n628 10.6151
R1412 B.n629 B.n294 10.6151
R1413 B.n639 B.n294 10.6151
R1414 B.n640 B.n639 10.6151
R1415 B.n641 B.n640 10.6151
R1416 B.n641 B.n286 10.6151
R1417 B.n651 B.n286 10.6151
R1418 B.n652 B.n651 10.6151
R1419 B.n653 B.n652 10.6151
R1420 B.n653 B.n278 10.6151
R1421 B.n663 B.n278 10.6151
R1422 B.n664 B.n663 10.6151
R1423 B.n665 B.n664 10.6151
R1424 B.n665 B.n270 10.6151
R1425 B.n676 B.n270 10.6151
R1426 B.n677 B.n676 10.6151
R1427 B.n678 B.n677 10.6151
R1428 B.n678 B.n263 10.6151
R1429 B.n689 B.n263 10.6151
R1430 B.n690 B.n689 10.6151
R1431 B.n691 B.n690 10.6151
R1432 B.n691 B.n0 10.6151
R1433 B.n520 B.n519 10.6151
R1434 B.n519 B.n518 10.6151
R1435 B.n518 B.n517 10.6151
R1436 B.n517 B.n515 10.6151
R1437 B.n515 B.n512 10.6151
R1438 B.n512 B.n511 10.6151
R1439 B.n511 B.n508 10.6151
R1440 B.n508 B.n507 10.6151
R1441 B.n507 B.n504 10.6151
R1442 B.n504 B.n503 10.6151
R1443 B.n503 B.n500 10.6151
R1444 B.n500 B.n499 10.6151
R1445 B.n499 B.n496 10.6151
R1446 B.n496 B.n495 10.6151
R1447 B.n495 B.n492 10.6151
R1448 B.n492 B.n491 10.6151
R1449 B.n491 B.n488 10.6151
R1450 B.n488 B.n487 10.6151
R1451 B.n487 B.n484 10.6151
R1452 B.n484 B.n483 10.6151
R1453 B.n483 B.n480 10.6151
R1454 B.n480 B.n479 10.6151
R1455 B.n479 B.n476 10.6151
R1456 B.n476 B.n475 10.6151
R1457 B.n472 B.n471 10.6151
R1458 B.n471 B.n468 10.6151
R1459 B.n468 B.n467 10.6151
R1460 B.n467 B.n464 10.6151
R1461 B.n464 B.n463 10.6151
R1462 B.n463 B.n460 10.6151
R1463 B.n460 B.n459 10.6151
R1464 B.n459 B.n456 10.6151
R1465 B.n456 B.n455 10.6151
R1466 B.n452 B.n451 10.6151
R1467 B.n451 B.n448 10.6151
R1468 B.n448 B.n447 10.6151
R1469 B.n447 B.n444 10.6151
R1470 B.n444 B.n443 10.6151
R1471 B.n443 B.n440 10.6151
R1472 B.n440 B.n439 10.6151
R1473 B.n439 B.n436 10.6151
R1474 B.n436 B.n435 10.6151
R1475 B.n435 B.n432 10.6151
R1476 B.n432 B.n431 10.6151
R1477 B.n431 B.n428 10.6151
R1478 B.n428 B.n427 10.6151
R1479 B.n427 B.n424 10.6151
R1480 B.n424 B.n423 10.6151
R1481 B.n423 B.n420 10.6151
R1482 B.n420 B.n419 10.6151
R1483 B.n419 B.n416 10.6151
R1484 B.n416 B.n415 10.6151
R1485 B.n415 B.n412 10.6151
R1486 B.n412 B.n411 10.6151
R1487 B.n411 B.n408 10.6151
R1488 B.n408 B.n370 10.6151
R1489 B.n525 B.n370 10.6151
R1490 B.n527 B.n526 10.6151
R1491 B.n527 B.n362 10.6151
R1492 B.n537 B.n362 10.6151
R1493 B.n538 B.n537 10.6151
R1494 B.n539 B.n538 10.6151
R1495 B.n539 B.n353 10.6151
R1496 B.n549 B.n353 10.6151
R1497 B.n550 B.n549 10.6151
R1498 B.n551 B.n550 10.6151
R1499 B.n551 B.n346 10.6151
R1500 B.n561 B.n346 10.6151
R1501 B.n562 B.n561 10.6151
R1502 B.n563 B.n562 10.6151
R1503 B.n563 B.n338 10.6151
R1504 B.n573 B.n338 10.6151
R1505 B.n574 B.n573 10.6151
R1506 B.n575 B.n574 10.6151
R1507 B.n575 B.n330 10.6151
R1508 B.n585 B.n330 10.6151
R1509 B.n586 B.n585 10.6151
R1510 B.n587 B.n586 10.6151
R1511 B.n587 B.n322 10.6151
R1512 B.n597 B.n322 10.6151
R1513 B.n598 B.n597 10.6151
R1514 B.n599 B.n598 10.6151
R1515 B.n599 B.n314 10.6151
R1516 B.n609 B.n314 10.6151
R1517 B.n610 B.n609 10.6151
R1518 B.n611 B.n610 10.6151
R1519 B.n611 B.n306 10.6151
R1520 B.n621 B.n306 10.6151
R1521 B.n622 B.n621 10.6151
R1522 B.n623 B.n622 10.6151
R1523 B.n623 B.n298 10.6151
R1524 B.n633 B.n298 10.6151
R1525 B.n634 B.n633 10.6151
R1526 B.n635 B.n634 10.6151
R1527 B.n635 B.n290 10.6151
R1528 B.n645 B.n290 10.6151
R1529 B.n646 B.n645 10.6151
R1530 B.n647 B.n646 10.6151
R1531 B.n647 B.n282 10.6151
R1532 B.n657 B.n282 10.6151
R1533 B.n658 B.n657 10.6151
R1534 B.n659 B.n658 10.6151
R1535 B.n659 B.n274 10.6151
R1536 B.n669 B.n274 10.6151
R1537 B.n670 B.n669 10.6151
R1538 B.n671 B.n670 10.6151
R1539 B.n671 B.n267 10.6151
R1540 B.n682 B.n267 10.6151
R1541 B.n683 B.n682 10.6151
R1542 B.n685 B.n683 10.6151
R1543 B.n685 B.n684 10.6151
R1544 B.n684 B.n259 10.6151
R1545 B.n696 B.n259 10.6151
R1546 B.n697 B.n696 10.6151
R1547 B.n698 B.n697 10.6151
R1548 B.n699 B.n698 10.6151
R1549 B.n700 B.n699 10.6151
R1550 B.n703 B.n700 10.6151
R1551 B.n704 B.n703 10.6151
R1552 B.n705 B.n704 10.6151
R1553 B.n706 B.n705 10.6151
R1554 B.n708 B.n706 10.6151
R1555 B.n709 B.n708 10.6151
R1556 B.n710 B.n709 10.6151
R1557 B.n711 B.n710 10.6151
R1558 B.n713 B.n711 10.6151
R1559 B.n714 B.n713 10.6151
R1560 B.n715 B.n714 10.6151
R1561 B.n716 B.n715 10.6151
R1562 B.n718 B.n716 10.6151
R1563 B.n719 B.n718 10.6151
R1564 B.n720 B.n719 10.6151
R1565 B.n721 B.n720 10.6151
R1566 B.n723 B.n721 10.6151
R1567 B.n724 B.n723 10.6151
R1568 B.n725 B.n724 10.6151
R1569 B.n726 B.n725 10.6151
R1570 B.n728 B.n726 10.6151
R1571 B.n729 B.n728 10.6151
R1572 B.n730 B.n729 10.6151
R1573 B.n731 B.n730 10.6151
R1574 B.n733 B.n731 10.6151
R1575 B.n734 B.n733 10.6151
R1576 B.n735 B.n734 10.6151
R1577 B.n736 B.n735 10.6151
R1578 B.n738 B.n736 10.6151
R1579 B.n739 B.n738 10.6151
R1580 B.n740 B.n739 10.6151
R1581 B.n741 B.n740 10.6151
R1582 B.n743 B.n741 10.6151
R1583 B.n744 B.n743 10.6151
R1584 B.n745 B.n744 10.6151
R1585 B.n746 B.n745 10.6151
R1586 B.n748 B.n746 10.6151
R1587 B.n749 B.n748 10.6151
R1588 B.n750 B.n749 10.6151
R1589 B.n751 B.n750 10.6151
R1590 B.n753 B.n751 10.6151
R1591 B.n754 B.n753 10.6151
R1592 B.n755 B.n754 10.6151
R1593 B.n756 B.n755 10.6151
R1594 B.n758 B.n756 10.6151
R1595 B.n759 B.n758 10.6151
R1596 B.n760 B.n759 10.6151
R1597 B.n761 B.n760 10.6151
R1598 B.n763 B.n761 10.6151
R1599 B.n764 B.n763 10.6151
R1600 B.n765 B.n764 10.6151
R1601 B.n766 B.n765 10.6151
R1602 B.n768 B.n766 10.6151
R1603 B.n769 B.n768 10.6151
R1604 B.n770 B.n769 10.6151
R1605 B.n884 B.n1 10.6151
R1606 B.n884 B.n883 10.6151
R1607 B.n883 B.n882 10.6151
R1608 B.n882 B.n10 10.6151
R1609 B.n876 B.n10 10.6151
R1610 B.n876 B.n875 10.6151
R1611 B.n875 B.n874 10.6151
R1612 B.n874 B.n17 10.6151
R1613 B.n868 B.n17 10.6151
R1614 B.n868 B.n867 10.6151
R1615 B.n867 B.n866 10.6151
R1616 B.n866 B.n25 10.6151
R1617 B.n860 B.n25 10.6151
R1618 B.n860 B.n859 10.6151
R1619 B.n859 B.n858 10.6151
R1620 B.n858 B.n32 10.6151
R1621 B.n852 B.n32 10.6151
R1622 B.n852 B.n851 10.6151
R1623 B.n851 B.n850 10.6151
R1624 B.n850 B.n39 10.6151
R1625 B.n844 B.n39 10.6151
R1626 B.n844 B.n843 10.6151
R1627 B.n843 B.n842 10.6151
R1628 B.n842 B.n46 10.6151
R1629 B.n836 B.n46 10.6151
R1630 B.n836 B.n835 10.6151
R1631 B.n835 B.n834 10.6151
R1632 B.n834 B.n53 10.6151
R1633 B.n828 B.n53 10.6151
R1634 B.n828 B.n827 10.6151
R1635 B.n827 B.n826 10.6151
R1636 B.n826 B.n60 10.6151
R1637 B.n820 B.n60 10.6151
R1638 B.n820 B.n819 10.6151
R1639 B.n819 B.n818 10.6151
R1640 B.n818 B.n67 10.6151
R1641 B.n812 B.n67 10.6151
R1642 B.n812 B.n811 10.6151
R1643 B.n811 B.n810 10.6151
R1644 B.n810 B.n74 10.6151
R1645 B.n804 B.n74 10.6151
R1646 B.n804 B.n803 10.6151
R1647 B.n803 B.n802 10.6151
R1648 B.n802 B.n81 10.6151
R1649 B.n796 B.n81 10.6151
R1650 B.n796 B.n795 10.6151
R1651 B.n795 B.n794 10.6151
R1652 B.n794 B.n88 10.6151
R1653 B.n788 B.n88 10.6151
R1654 B.n788 B.n787 10.6151
R1655 B.n787 B.n786 10.6151
R1656 B.n786 B.n95 10.6151
R1657 B.n780 B.n95 10.6151
R1658 B.n780 B.n779 10.6151
R1659 B.n779 B.n778 10.6151
R1660 B.n778 B.n102 10.6151
R1661 B.n142 B.n141 10.6151
R1662 B.n145 B.n142 10.6151
R1663 B.n146 B.n145 10.6151
R1664 B.n149 B.n146 10.6151
R1665 B.n150 B.n149 10.6151
R1666 B.n153 B.n150 10.6151
R1667 B.n154 B.n153 10.6151
R1668 B.n157 B.n154 10.6151
R1669 B.n158 B.n157 10.6151
R1670 B.n161 B.n158 10.6151
R1671 B.n162 B.n161 10.6151
R1672 B.n165 B.n162 10.6151
R1673 B.n166 B.n165 10.6151
R1674 B.n169 B.n166 10.6151
R1675 B.n170 B.n169 10.6151
R1676 B.n173 B.n170 10.6151
R1677 B.n174 B.n173 10.6151
R1678 B.n177 B.n174 10.6151
R1679 B.n178 B.n177 10.6151
R1680 B.n181 B.n178 10.6151
R1681 B.n182 B.n181 10.6151
R1682 B.n185 B.n182 10.6151
R1683 B.n186 B.n185 10.6151
R1684 B.n189 B.n186 10.6151
R1685 B.n194 B.n191 10.6151
R1686 B.n195 B.n194 10.6151
R1687 B.n198 B.n195 10.6151
R1688 B.n199 B.n198 10.6151
R1689 B.n202 B.n199 10.6151
R1690 B.n203 B.n202 10.6151
R1691 B.n206 B.n203 10.6151
R1692 B.n207 B.n206 10.6151
R1693 B.n210 B.n207 10.6151
R1694 B.n215 B.n212 10.6151
R1695 B.n216 B.n215 10.6151
R1696 B.n219 B.n216 10.6151
R1697 B.n220 B.n219 10.6151
R1698 B.n223 B.n220 10.6151
R1699 B.n224 B.n223 10.6151
R1700 B.n227 B.n224 10.6151
R1701 B.n228 B.n227 10.6151
R1702 B.n231 B.n228 10.6151
R1703 B.n232 B.n231 10.6151
R1704 B.n235 B.n232 10.6151
R1705 B.n236 B.n235 10.6151
R1706 B.n239 B.n236 10.6151
R1707 B.n240 B.n239 10.6151
R1708 B.n243 B.n240 10.6151
R1709 B.n244 B.n243 10.6151
R1710 B.n247 B.n244 10.6151
R1711 B.n248 B.n247 10.6151
R1712 B.n251 B.n248 10.6151
R1713 B.n252 B.n251 10.6151
R1714 B.n255 B.n252 10.6151
R1715 B.n257 B.n255 10.6151
R1716 B.n258 B.n257 10.6151
R1717 B.n771 B.n258 10.6151
R1718 B.n475 B.n404 9.36635
R1719 B.n452 B.n407 9.36635
R1720 B.n190 B.n189 9.36635
R1721 B.n212 B.n211 9.36635
R1722 B.n892 B.n0 8.11757
R1723 B.n892 B.n1 8.11757
R1724 B.n649 B.t1 7.55739
R1725 B.n856 B.t6 7.55739
R1726 B.n680 B.t0 1.88972
R1727 B.n878 B.t3 1.88972
R1728 B.n472 B.n404 1.24928
R1729 B.n455 B.n407 1.24928
R1730 B.n191 B.n190 1.24928
R1731 B.n211 B.n210 1.24928
R1732 VN.n63 VN.n33 161.3
R1733 VN.n62 VN.n61 161.3
R1734 VN.n60 VN.n34 161.3
R1735 VN.n59 VN.n58 161.3
R1736 VN.n57 VN.n35 161.3
R1737 VN.n56 VN.n55 161.3
R1738 VN.n54 VN.n36 161.3
R1739 VN.n53 VN.n52 161.3
R1740 VN.n51 VN.n37 161.3
R1741 VN.n50 VN.n49 161.3
R1742 VN.n48 VN.n39 161.3
R1743 VN.n47 VN.n46 161.3
R1744 VN.n45 VN.n40 161.3
R1745 VN.n44 VN.n43 161.3
R1746 VN.n30 VN.n0 161.3
R1747 VN.n29 VN.n28 161.3
R1748 VN.n27 VN.n1 161.3
R1749 VN.n26 VN.n25 161.3
R1750 VN.n24 VN.n2 161.3
R1751 VN.n23 VN.n22 161.3
R1752 VN.n21 VN.n3 161.3
R1753 VN.n20 VN.n19 161.3
R1754 VN.n17 VN.n4 161.3
R1755 VN.n16 VN.n15 161.3
R1756 VN.n14 VN.n5 161.3
R1757 VN.n13 VN.n12 161.3
R1758 VN.n11 VN.n6 161.3
R1759 VN.n10 VN.n9 161.3
R1760 VN.n32 VN.n31 109.534
R1761 VN.n65 VN.n64 109.534
R1762 VN.n8 VN.t4 83.102
R1763 VN.n42 VN.t6 83.102
R1764 VN.n8 VN.n7 65.4202
R1765 VN.n42 VN.n41 65.4202
R1766 VN.n25 VN.n24 55.0624
R1767 VN.n58 VN.n57 55.0624
R1768 VN.n7 VN.t5 50.8339
R1769 VN.n18 VN.t0 50.8339
R1770 VN.n31 VN.t1 50.8339
R1771 VN.n41 VN.t3 50.8339
R1772 VN.n38 VN.t7 50.8339
R1773 VN.n64 VN.t2 50.8339
R1774 VN VN.n65 48.8618
R1775 VN.n12 VN.n5 40.4934
R1776 VN.n16 VN.n5 40.4934
R1777 VN.n46 VN.n39 40.4934
R1778 VN.n50 VN.n39 40.4934
R1779 VN.n25 VN.n1 25.9244
R1780 VN.n58 VN.n34 25.9244
R1781 VN.n11 VN.n10 24.4675
R1782 VN.n12 VN.n11 24.4675
R1783 VN.n17 VN.n16 24.4675
R1784 VN.n19 VN.n17 24.4675
R1785 VN.n23 VN.n3 24.4675
R1786 VN.n24 VN.n23 24.4675
R1787 VN.n29 VN.n1 24.4675
R1788 VN.n30 VN.n29 24.4675
R1789 VN.n46 VN.n45 24.4675
R1790 VN.n45 VN.n44 24.4675
R1791 VN.n57 VN.n56 24.4675
R1792 VN.n56 VN.n36 24.4675
R1793 VN.n52 VN.n51 24.4675
R1794 VN.n51 VN.n50 24.4675
R1795 VN.n63 VN.n62 24.4675
R1796 VN.n62 VN.n34 24.4675
R1797 VN.n18 VN.n3 15.9041
R1798 VN.n38 VN.n36 15.9041
R1799 VN.n10 VN.n7 8.56395
R1800 VN.n19 VN.n18 8.56395
R1801 VN.n44 VN.n41 8.56395
R1802 VN.n52 VN.n38 8.56395
R1803 VN.n43 VN.n42 5.17456
R1804 VN.n9 VN.n8 5.17456
R1805 VN.n31 VN.n30 1.22385
R1806 VN.n64 VN.n63 1.22385
R1807 VN.n65 VN.n33 0.278367
R1808 VN.n32 VN.n0 0.278367
R1809 VN.n61 VN.n33 0.189894
R1810 VN.n61 VN.n60 0.189894
R1811 VN.n60 VN.n59 0.189894
R1812 VN.n59 VN.n35 0.189894
R1813 VN.n55 VN.n35 0.189894
R1814 VN.n55 VN.n54 0.189894
R1815 VN.n54 VN.n53 0.189894
R1816 VN.n53 VN.n37 0.189894
R1817 VN.n49 VN.n37 0.189894
R1818 VN.n49 VN.n48 0.189894
R1819 VN.n48 VN.n47 0.189894
R1820 VN.n47 VN.n40 0.189894
R1821 VN.n43 VN.n40 0.189894
R1822 VN.n9 VN.n6 0.189894
R1823 VN.n13 VN.n6 0.189894
R1824 VN.n14 VN.n13 0.189894
R1825 VN.n15 VN.n14 0.189894
R1826 VN.n15 VN.n4 0.189894
R1827 VN.n20 VN.n4 0.189894
R1828 VN.n21 VN.n20 0.189894
R1829 VN.n22 VN.n21 0.189894
R1830 VN.n22 VN.n2 0.189894
R1831 VN.n26 VN.n2 0.189894
R1832 VN.n27 VN.n26 0.189894
R1833 VN.n28 VN.n27 0.189894
R1834 VN.n28 VN.n0 0.189894
R1835 VN VN.n32 0.153454
R1836 VDD2.n2 VDD2.n1 68.1784
R1837 VDD2.n2 VDD2.n0 68.1784
R1838 VDD2 VDD2.n5 68.1756
R1839 VDD2.n4 VDD2.n3 66.79
R1840 VDD2.n4 VDD2.n2 42.2024
R1841 VDD2.n5 VDD2.t4 3.10882
R1842 VDD2.n5 VDD2.t1 3.10882
R1843 VDD2.n3 VDD2.t5 3.10882
R1844 VDD2.n3 VDD2.t0 3.10882
R1845 VDD2.n1 VDD2.t7 3.10882
R1846 VDD2.n1 VDD2.t6 3.10882
R1847 VDD2.n0 VDD2.t3 3.10882
R1848 VDD2.n0 VDD2.t2 3.10882
R1849 VDD2 VDD2.n4 1.50266
C0 VN VDD1 0.152537f
C1 VTAIL VP 5.96607f
C2 VDD2 VP 0.564413f
C3 VN VP 7.13172f
C4 VDD1 VP 5.36853f
C5 VDD2 VTAIL 6.50933f
C6 VTAIL VN 5.95197f
C7 VDD2 VN 4.95827f
C8 VTAIL VDD1 6.4521f
C9 VDD2 VDD1 1.99652f
C10 VDD2 B 5.307961f
C11 VDD1 B 5.79977f
C12 VTAIL B 6.959456f
C13 VN B 16.499208f
C14 VP B 15.132747f
C15 VDD2.t3 B 0.12182f
C16 VDD2.t2 B 0.12182f
C17 VDD2.n0 B 1.0343f
C18 VDD2.t7 B 0.12182f
C19 VDD2.t6 B 0.12182f
C20 VDD2.n1 B 1.0343f
C21 VDD2.n2 B 3.06861f
C22 VDD2.t5 B 0.12182f
C23 VDD2.t0 B 0.12182f
C24 VDD2.n3 B 1.02328f
C25 VDD2.n4 B 2.57602f
C26 VDD2.t4 B 0.12182f
C27 VDD2.t1 B 0.12182f
C28 VDD2.n5 B 1.03426f
C29 VN.n0 B 0.029854f
C30 VN.t1 B 1.15693f
C31 VN.n1 B 0.043303f
C32 VN.n2 B 0.022644f
C33 VN.n3 B 0.03491f
C34 VN.n4 B 0.022644f
C35 VN.n5 B 0.018306f
C36 VN.n6 B 0.022644f
C37 VN.t5 B 1.15693f
C38 VN.n7 B 0.497124f
C39 VN.t4 B 1.38419f
C40 VN.n8 B 0.479446f
C41 VN.n9 B 0.243269f
C42 VN.n10 B 0.028659f
C43 VN.n11 B 0.042204f
C44 VN.n12 B 0.045006f
C45 VN.n13 B 0.022644f
C46 VN.n14 B 0.022644f
C47 VN.n15 B 0.022644f
C48 VN.n16 B 0.045006f
C49 VN.n17 B 0.042204f
C50 VN.t0 B 1.15693f
C51 VN.n18 B 0.427771f
C52 VN.n19 B 0.028659f
C53 VN.n20 B 0.022644f
C54 VN.n21 B 0.022644f
C55 VN.n22 B 0.022644f
C56 VN.n23 B 0.042204f
C57 VN.n24 B 0.039191f
C58 VN.n25 B 0.025823f
C59 VN.n26 B 0.022644f
C60 VN.n27 B 0.022644f
C61 VN.n28 B 0.022644f
C62 VN.n29 B 0.042204f
C63 VN.n30 B 0.022408f
C64 VN.n31 B 0.505313f
C65 VN.n32 B 0.045093f
C66 VN.n33 B 0.029854f
C67 VN.t2 B 1.15693f
C68 VN.n34 B 0.043303f
C69 VN.n35 B 0.022644f
C70 VN.n36 B 0.03491f
C71 VN.n37 B 0.022644f
C72 VN.t7 B 1.15693f
C73 VN.n38 B 0.427771f
C74 VN.n39 B 0.018306f
C75 VN.n40 B 0.022644f
C76 VN.t3 B 1.15693f
C77 VN.n41 B 0.497124f
C78 VN.t6 B 1.38419f
C79 VN.n42 B 0.479446f
C80 VN.n43 B 0.243269f
C81 VN.n44 B 0.028659f
C82 VN.n45 B 0.042204f
C83 VN.n46 B 0.045006f
C84 VN.n47 B 0.022644f
C85 VN.n48 B 0.022644f
C86 VN.n49 B 0.022644f
C87 VN.n50 B 0.045006f
C88 VN.n51 B 0.042204f
C89 VN.n52 B 0.028659f
C90 VN.n53 B 0.022644f
C91 VN.n54 B 0.022644f
C92 VN.n55 B 0.022644f
C93 VN.n56 B 0.042204f
C94 VN.n57 B 0.039191f
C95 VN.n58 B 0.025823f
C96 VN.n59 B 0.022644f
C97 VN.n60 B 0.022644f
C98 VN.n61 B 0.022644f
C99 VN.n62 B 0.042204f
C100 VN.n63 B 0.022408f
C101 VN.n64 B 0.505313f
C102 VN.n65 B 1.22836f
C103 VDD1.t5 B 0.125085f
C104 VDD1.t7 B 0.125085f
C105 VDD1.n0 B 1.06312f
C106 VDD1.t4 B 0.125085f
C107 VDD1.t3 B 0.125085f
C108 VDD1.n1 B 1.06202f
C109 VDD1.t0 B 0.125085f
C110 VDD1.t2 B 0.125085f
C111 VDD1.n2 B 1.06202f
C112 VDD1.n3 B 3.20254f
C113 VDD1.t6 B 0.125085f
C114 VDD1.t1 B 0.125085f
C115 VDD1.n4 B 1.0507f
C116 VDD1.n5 B 2.67584f
C117 VTAIL.t6 B 0.119129f
C118 VTAIL.t2 B 0.119129f
C119 VTAIL.n0 B 0.937904f
C120 VTAIL.n1 B 0.448345f
C121 VTAIL.t3 B 1.196f
C122 VTAIL.n2 B 0.546534f
C123 VTAIL.t9 B 1.196f
C124 VTAIL.n3 B 0.546534f
C125 VTAIL.t8 B 0.119129f
C126 VTAIL.t13 B 0.119129f
C127 VTAIL.n4 B 0.937904f
C128 VTAIL.n5 B 0.664133f
C129 VTAIL.t15 B 1.196f
C130 VTAIL.n6 B 1.47116f
C131 VTAIL.t4 B 1.19601f
C132 VTAIL.n7 B 1.47116f
C133 VTAIL.t5 B 0.119129f
C134 VTAIL.t1 B 0.119129f
C135 VTAIL.n8 B 0.937909f
C136 VTAIL.n9 B 0.664128f
C137 VTAIL.t0 B 1.19601f
C138 VTAIL.n10 B 0.546527f
C139 VTAIL.t11 B 1.19601f
C140 VTAIL.n11 B 0.546527f
C141 VTAIL.t12 B 0.119129f
C142 VTAIL.t14 B 0.119129f
C143 VTAIL.n12 B 0.937909f
C144 VTAIL.n13 B 0.664128f
C145 VTAIL.t10 B 1.196f
C146 VTAIL.n14 B 1.47116f
C147 VTAIL.t7 B 1.196f
C148 VTAIL.n15 B 1.46673f
C149 VP.n0 B 0.030568f
C150 VP.t5 B 1.18458f
C151 VP.n1 B 0.044338f
C152 VP.n2 B 0.023186f
C153 VP.n3 B 0.035744f
C154 VP.n4 B 0.023186f
C155 VP.n5 B 0.018743f
C156 VP.n6 B 0.023186f
C157 VP.t4 B 1.18458f
C158 VP.n7 B 0.437994f
C159 VP.n8 B 0.023186f
C160 VP.n9 B 0.02644f
C161 VP.n10 B 0.023186f
C162 VP.t3 B 1.18458f
C163 VP.n11 B 0.51739f
C164 VP.n12 B 0.030568f
C165 VP.t6 B 1.18458f
C166 VP.n13 B 0.044338f
C167 VP.n14 B 0.023186f
C168 VP.n15 B 0.035744f
C169 VP.n16 B 0.023186f
C170 VP.n17 B 0.018743f
C171 VP.n18 B 0.023186f
C172 VP.t0 B 1.18458f
C173 VP.n19 B 0.509005f
C174 VP.t2 B 1.41727f
C175 VP.n20 B 0.490904f
C176 VP.n21 B 0.249083f
C177 VP.n22 B 0.029344f
C178 VP.n23 B 0.043212f
C179 VP.n24 B 0.046081f
C180 VP.n25 B 0.023186f
C181 VP.n26 B 0.023186f
C182 VP.n27 B 0.023186f
C183 VP.n28 B 0.046081f
C184 VP.n29 B 0.043212f
C185 VP.t1 B 1.18458f
C186 VP.n30 B 0.437994f
C187 VP.n31 B 0.029344f
C188 VP.n32 B 0.023186f
C189 VP.n33 B 0.023186f
C190 VP.n34 B 0.023186f
C191 VP.n35 B 0.043212f
C192 VP.n36 B 0.040128f
C193 VP.n37 B 0.02644f
C194 VP.n38 B 0.023186f
C195 VP.n39 B 0.023186f
C196 VP.n40 B 0.023186f
C197 VP.n41 B 0.043212f
C198 VP.n42 B 0.022944f
C199 VP.n43 B 0.51739f
C200 VP.n44 B 1.24521f
C201 VP.n45 B 1.26236f
C202 VP.n46 B 0.030568f
C203 VP.n47 B 0.022944f
C204 VP.n48 B 0.043212f
C205 VP.n49 B 0.044338f
C206 VP.n50 B 0.023186f
C207 VP.n51 B 0.023186f
C208 VP.n52 B 0.023186f
C209 VP.n53 B 0.040128f
C210 VP.n54 B 0.043212f
C211 VP.n55 B 0.035744f
C212 VP.n56 B 0.023186f
C213 VP.n57 B 0.023186f
C214 VP.n58 B 0.029344f
C215 VP.n59 B 0.043212f
C216 VP.n60 B 0.046081f
C217 VP.n61 B 0.023186f
C218 VP.n62 B 0.023186f
C219 VP.n63 B 0.023186f
C220 VP.n64 B 0.046081f
C221 VP.n65 B 0.043212f
C222 VP.t7 B 1.18458f
C223 VP.n66 B 0.437994f
C224 VP.n67 B 0.029344f
C225 VP.n68 B 0.023186f
C226 VP.n69 B 0.023186f
C227 VP.n70 B 0.023186f
C228 VP.n71 B 0.043212f
C229 VP.n72 B 0.040128f
C230 VP.n73 B 0.02644f
C231 VP.n74 B 0.023186f
C232 VP.n75 B 0.023186f
C233 VP.n76 B 0.023186f
C234 VP.n77 B 0.043212f
C235 VP.n78 B 0.022944f
C236 VP.n79 B 0.51739f
C237 VP.n80 B 0.046171f
.ends

