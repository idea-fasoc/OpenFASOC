* NGSPICE file created from opamp_sample_0005.ext - technology: sky130A

.subckt opamp_sample_0005 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VOUT.t84 a_n7097_7899.t16 VDD.t187 VDD.t154 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X1 VDD.t186 a_n7097_7899.t17 VOUT.t83 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 VOUT.t14 CS_BIAS.t32 GND.t179 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X3 VDD.t96 VDD.t94 VDD.t95 VDD.t71 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X4 VOUT.t82 a_n7097_7899.t18 VDD.t185 VDD.t150 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 VOUT.t85 CS_BIAS.t33 GND.t178 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X6 VDD.t93 VDD.t91 VDD.t92 VDD.t64 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X7 VDD.t90 VDD.t88 VDD.t89 VDD.t51 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 a_n7097_7899.t10 VN.t5 a_n1455_n3628.t19 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X9 VOUT.t81 a_n7097_7899.t19 VDD.t184 VDD.t150 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 VDD.t87 VDD.t85 VDD.t86 VDD.t78 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X11 VDD.t84 VDD.t81 VDD.t83 VDD.t82 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X12 VDD.t183 a_n7097_7899.t20 VOUT.t80 VDD.t147 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 GND.t177 CS_BIAS.t0 CS_BIAS.t1 GND.t145 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X14 VDD.t191 a_n2433_10060.t24 a_n2511_10256.t7 VDD.t190 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X15 VDD.t182 a_n7097_7899.t21 VOUT.t79 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 VOUT.t1 CS_BIAS.t34 GND.t176 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X17 a_n2433_10060.t3 VP.t5 a_n1455_n3628.t4 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X18 a_n2511_10256.t15 a_n2433_10060.t9 a_n2433_10060.t10 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 a_n1455_n3628.t5 DIFFPAIR_BIAS.t8 GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X20 a_n1455_n3628.t3 VP.t6 a_n2433_10060.t2 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X21 VOUT.t2 CS_BIAS.t35 GND.t175 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X22 VOUT.t19 CS_BIAS.t36 GND.t174 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X23 VDD.t181 a_n7097_7899.t22 VOUT.t78 VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 VOUT.t77 a_n7097_7899.t23 VDD.t180 VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 GND.t173 CS_BIAS.t37 VOUT.t0 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X26 VOUT.t76 a_n7097_7899.t24 VDD.t179 VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X28 VN.t4 GND.t113 GND.t115 GND.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 GND.t112 GND.t109 GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X30 VDD.t2 a_n2433_10060.t25 a_n2511_10256.t6 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X31 VDD.t13 a_n2433_10060.t26 a_n2154_8322.t7 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X32 GND.t155 CS_BIAS.t38 VOUT.t17 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X33 VOUT.t75 a_n7097_7899.t25 VDD.t178 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 GND.t108 GND.t106 VP.t4 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X35 GND.t105 GND.t102 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X36 GND.t172 CS_BIAS.t6 CS_BIAS.t7 GND.t140 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X37 GND.t171 CS_BIAS.t39 VOUT.t11 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X38 VOUT.t8 CS_BIAS.t40 GND.t170 GND.t158 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X39 VDD.t80 VDD.t77 VDD.t79 VDD.t78 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X40 VOUT.t74 a_n7097_7899.t26 VDD.t177 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 VDD.t176 a_n7097_7899.t27 VOUT.t73 VDD.t128 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X42 CS_BIAS.t29 CS_BIAS.t28 GND.t169 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X43 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X44 CS_BIAS.t27 CS_BIAS.t26 GND.t168 GND.t158 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X45 a_n1455_n3628.t9 VP.t7 a_n2433_10060.t5 GND.t19 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X46 GND.t101 GND.t99 GND.t100 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X47 GND.t98 GND.t96 VP.t3 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X48 GND.t167 CS_BIAS.t24 CS_BIAS.t25 GND.t136 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X49 VDD.t76 VDD.t74 VDD.t75 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X50 VDD.t8 a_n2433_10060.t27 a_n2154_8322.t6 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X51 VOUT.t72 a_n7097_7899.t28 VDD.t175 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n1455_n3628.t8 DIFFPAIR_BIAS.t9 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X53 VDD.t159 a_n7097_7899.t29 VOUT.t71 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X54 GND.t166 CS_BIAS.t22 CS_BIAS.t23 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X55 a_n7097_7899.t3 VN.t6 a_n1455_n3628.t18 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X56 VOUT.t92 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X57 VDD.t106 a_n2433_10060.t28 a_n2511_10256.t5 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X58 a_n2511_10256.t4 a_n2433_10060.t29 VDD.t193 VDD.t192 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X59 VOUT.t93 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X60 VDD.t73 VDD.t70 VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X61 CS_BIAS.t11 CS_BIAS.t10 GND.t165 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X62 VOUT.t70 a_n7097_7899.t30 VDD.t174 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 VDD.t173 a_n7097_7899.t31 VOUT.t69 VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 VN.t3 GND.t93 GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X65 GND.t164 CS_BIAS.t8 CS_BIAS.t9 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X66 VDD.t172 a_n7097_7899.t32 VOUT.t68 VDD.t133 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 VOUT.t21 CS_BIAS.t41 GND.t163 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X68 GND.t92 GND.t90 GND.t91 GND.t59 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X69 VDD.t69 VDD.t67 VDD.t68 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X70 VDD.t171 a_n7097_7899.t33 VOUT.t67 VDD.t128 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X71 a_n2433_10060.t8 a_n2433_10060.t7 a_n2511_10256.t14 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X72 a_n1455_n3628.t17 VN.t7 a_n7097_7899.t9 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X73 GND.t162 CS_BIAS.t42 VOUT.t20 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X74 VDD.t170 a_n7097_7899.t34 VOUT.t66 VDD.t126 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X75 VDD.t169 a_n7097_7899.t35 VOUT.t65 VDD.t133 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 GND.t161 CS_BIAS.t43 VOUT.t91 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X77 VOUT.t64 a_n7097_7899.t36 VDD.t168 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 GND.t160 CS_BIAS.t20 CS_BIAS.t21 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X79 VOUT.t5 CS_BIAS.t44 GND.t159 GND.t158 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X80 a_n2154_8322.t15 a_n2433_10060.t30 a_n7097_7899.t4 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X81 VOUT.t63 a_n7097_7899.t37 VDD.t165 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 VOUT.t18 CS_BIAS.t45 GND.t153 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X83 VOUT.t62 a_n7097_7899.t38 VDD.t167 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 VDD.t100 a_n2433_10060.t31 a_n2154_8322.t5 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X85 VDD.t166 a_n7097_7899.t39 VOUT.t61 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 CS_BIAS.t19 CS_BIAS.t18 GND.t157 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X87 VOUT.t60 a_n7097_7899.t40 VDD.t164 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 GND.t156 CS_BIAS.t46 VOUT.t90 GND.t145 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X89 GND.t89 GND.t87 GND.t88 GND.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X90 VDD.t163 a_n7097_7899.t41 VOUT.t59 VDD.t116 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n7097_7899.t11 a_n2433_10060.t32 a_n2154_8322.t14 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X92 VDD.t66 VDD.t63 VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X93 GND.t86 GND.t84 GND.t85 GND.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X94 VOUT.t58 a_n7097_7899.t42 VDD.t162 VDD.t154 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 VDD.t161 a_n7097_7899.t43 VOUT.t57 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 VOUT.t9 CS_BIAS.t47 GND.t152 GND.t143 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X97 VDD.t11 a_n2433_10060.t33 a_n2154_8322.t4 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X98 VDD.t62 VDD.t60 VDD.t61 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X99 GND.t83 GND.t81 VN.t2 GND.t82 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X100 a_n7097_7899.t1 VN.t8 a_n1455_n3628.t16 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X101 VOUT.t56 a_n7097_7899.t44 VDD.t160 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 VP.t2 GND.t78 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X103 CS_BIAS.t17 CS_BIAS.t16 GND.t151 GND.t143 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X104 a_n2154_8322.t3 a_n2433_10060.t34 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X105 a_n2511_10256.t3 a_n2433_10060.t35 VDD.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X106 VOUT.t94 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X107 VOUT.t55 a_n7097_7899.t45 VDD.t158 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X108 GND.t150 CS_BIAS.t48 VOUT.t3 GND.t140 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X109 a_n2511_10256.t2 a_n2433_10060.t36 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X110 a_n2154_8322.t13 a_n2433_10060.t37 a_n7097_7899.t2 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X111 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X112 VDD.t157 a_n7097_7899.t46 VOUT.t54 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 VDD.t59 VDD.t57 VDD.t58 VDD.t51 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X114 VOUT.t53 a_n7097_7899.t47 VDD.t156 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 VOUT.t52 a_n7097_7899.t48 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X116 GND.t77 GND.t75 GND.t76 GND.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X117 VDD.t153 a_n7097_7899.t49 VOUT.t51 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 a_n2433_10060.t18 a_n2433_10060.t17 a_n2511_10256.t13 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X119 VOUT.t89 CS_BIAS.t49 GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X120 VDD.t56 VDD.t54 VDD.t55 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X121 GND.t147 CS_BIAS.t50 VOUT.t10 GND.t136 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X122 VOUT.t50 a_n7097_7899.t50 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 a_n1455_n3628.t2 VP.t8 a_n2433_10060.t1 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X124 GND.t146 CS_BIAS.t51 VOUT.t12 GND.t145 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X125 GND.t74 GND.t72 GND.t73 GND.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X126 VDD.t4 a_n2433_10060.t38 a_n2511_10256.t1 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 VDD.t53 VDD.t50 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X128 VDD.t49 VDD.t47 VDD.t48 VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X129 a_n2154_8322.t12 a_n2433_10060.t39 a_n7097_7899.t14 VDD.t102 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X130 GND.t71 GND.t69 VN.t1 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X131 VOUT.t95 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X132 VDD.t149 a_n7097_7899.t51 VOUT.t49 VDD.t147 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 a_n1455_n3628.t7 DIFFPAIR_BIAS.t10 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X134 GND.t68 GND.t66 GND.t67 GND.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X135 a_n2511_10256.t0 a_n2433_10060.t40 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X136 VDD.t148 a_n7097_7899.t52 VOUT.t48 VDD.t147 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 VOUT.t47 a_n7097_7899.t53 VDD.t144 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 VDD.t146 a_n7097_7899.t54 VOUT.t46 VDD.t145 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 VOUT.t87 CS_BIAS.t52 GND.t144 GND.t143 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X140 VDD.t143 a_n7097_7899.t55 VOUT.t45 VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 a_n2154_8322.t11 a_n2433_10060.t41 a_n7097_7899.t5 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X142 a_n2433_10060.t4 VP.t9 a_n1455_n3628.t6 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X143 VOUT.t44 a_n7097_7899.t56 VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 a_n1455_n3628.t15 VN.t9 a_n7097_7899.t15 GND.t19 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X145 a_n2511_10256.t12 a_n2433_10060.t15 a_n2433_10060.t16 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X146 GND.t139 CS_BIAS.t53 VOUT.t88 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X147 GND.t142 CS_BIAS.t54 VOUT.t6 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X148 VOUT.t43 a_n7097_7899.t57 VDD.t139 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n2433_10060.t23 VP.t10 a_n1455_n3628.t11 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X150 a_n7097_7899.t6 VN.t10 a_n1455_n3628.t14 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X151 GND.t141 CS_BIAS.t55 VOUT.t7 GND.t140 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X152 a_n1455_n3628.t13 VN.t11 a_n7097_7899.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X153 a_n7097_7899.t12 a_n2433_10060.t42 a_n2154_8322.t10 VDD.t101 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X154 VDD.t138 a_n7097_7899.t58 VOUT.t42 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 a_n7097_7899.t13 a_n2433_10060.t43 a_n2154_8322.t9 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X156 VDD.t46 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 VDD.t137 a_n7097_7899.t59 VOUT.t41 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 GND.t65 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X159 GND.t61 GND.t58 GND.t60 GND.t59 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X160 a_n2511_10256.t11 a_n2433_10060.t13 a_n2433_10060.t14 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X161 a_n2511_10256.t10 a_n2433_10060.t11 a_n2433_10060.t12 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X162 VDD.t42 VDD.t40 VDD.t41 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X163 CS_BIAS.t15 CS_BIAS.t14 GND.t138 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X164 GND.t137 CS_BIAS.t56 VOUT.t23 GND.t136 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X165 a_n1455_n3628.t1 VP.t11 a_n2433_10060.t0 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X166 GND.t57 GND.t55 GND.t56 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X167 VOUT.t40 a_n7097_7899.t60 VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 VDD.t39 VDD.t36 VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X169 a_n1455_n3628.t0 DIFFPAIR_BIAS.t11 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X170 VOUT.t96 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X171 GND.t54 GND.t52 GND.t53 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X172 VDD.t134 a_n7097_7899.t61 VOUT.t39 VDD.t133 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 GND.t135 CS_BIAS.t4 CS_BIAS.t5 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X174 VDD.t35 VDD.t32 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X175 VDD.t130 a_n7097_7899.t62 VOUT.t38 VDD.t126 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X176 VOUT.t37 a_n7097_7899.t63 VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 VDD.t31 VDD.t29 VDD.t30 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X178 VOUT.t97 a_n2154_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X179 VDD.t129 a_n7097_7899.t64 VOUT.t36 VDD.t128 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X180 VDD.t28 VDD.t25 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X181 VDD.t127 a_n7097_7899.t65 VOUT.t35 VDD.t126 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X182 a_n2154_8322.t2 a_n2433_10060.t44 VDD.t195 VDD.t194 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X183 GND.t134 CS_BIAS.t2 CS_BIAS.t3 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X184 VP.t1 GND.t49 GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X185 GND.t132 CS_BIAS.t57 VOUT.t22 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X186 GND.t130 CS_BIAS.t58 VOUT.t4 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X187 VOUT.t13 CS_BIAS.t59 GND.t128 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X188 VOUT.t34 a_n7097_7899.t66 VDD.t125 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X190 VOUT.t33 a_n7097_7899.t67 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 GND.t48 GND.t46 GND.t47 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X192 VOUT.t15 CS_BIAS.t60 GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X193 a_n2154_8322.t1 a_n2433_10060.t45 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X194 CS_BIAS.t31 CS_BIAS.t30 GND.t124 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X195 VOUT.t32 a_n7097_7899.t68 VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 VOUT.t31 a_n7097_7899.t69 VDD.t121 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 VDD.t118 a_n7097_7899.t70 VOUT.t30 VDD.t116 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 GND.t45 GND.t42 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X199 VDD.t117 a_n7097_7899.t71 VOUT.t29 VDD.t116 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 a_n2433_10060.t22 a_n2433_10060.t21 a_n2511_10256.t9 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X201 VOUT.t86 CS_BIAS.t61 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X202 VOUT.t16 CS_BIAS.t62 GND.t121 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X203 VDD.t24 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 GND.t41 GND.t38 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X205 VOUT.t28 a_n7097_7899.t72 VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 GND.t37 GND.t34 GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X207 GND.t30 GND.t28 VN.t0 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X208 a_n2154_8322.t0 a_n2433_10060.t46 VDD.t189 VDD.t188 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X209 VDD.t113 a_n7097_7899.t73 VOUT.t27 VDD.t112 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 GND.t119 CS_BIAS.t63 VOUT.t24 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X211 a_n2433_10060.t20 a_n2433_10060.t19 a_n2511_10256.t8 VDD.t9 sky130_fd_pr__pfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X212 VOUT.t26 a_n7097_7899.t74 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X213 a_n1455_n3628.t12 VN.t12 a_n7097_7899.t8 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X214 VDD.t109 a_n7097_7899.t75 VOUT.t25 VDD.t108 sky130_fd_pr__pfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 CS_BIAS.t13 CS_BIAS.t12 GND.t117 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X216 a_n2433_10060.t6 VP.t12 a_n1455_n3628.t10 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X217 a_n7097_7899.t0 a_n2433_10060.t47 a_n2154_8322.t8 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X218 GND.t33 GND.t31 VP.t0 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X219 GND.t27 GND.t24 GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
R0 a_n7097_7899.n168 a_n7097_7899.t69 223.136
R1 a_n7097_7899.n156 a_n7097_7899.t45 223.136
R2 a_n7097_7899.n145 a_n7097_7899.t74 223.136
R3 a_n7097_7899.n129 a_n7097_7899.t62 223.136
R4 a_n7097_7899.n114 a_n7097_7899.t34 223.136
R5 a_n7097_7899.n100 a_n7097_7899.t65 223.136
R6 a_n7097_7899.n11 a_n7097_7899.t27 223.097
R7 a_n7097_7899.n10 a_n7097_7899.t33 223.097
R8 a_n7097_7899.n9 a_n7097_7899.t64 223.097
R9 a_n7097_7899.n138 a_n7097_7899.t42 207.983
R10 a_n7097_7899.n123 a_n7097_7899.t16 207.983
R11 a_n7097_7899.n109 a_n7097_7899.t48 207.983
R12 a_n7097_7899.n174 a_n7097_7899.t37 168.701
R13 a_n7097_7899.n173 a_n7097_7899.t70 168.701
R14 a_n7097_7899.n164 a_n7097_7899.t19 168.701
R15 a_n7097_7899.n170 a_n7097_7899.t31 168.701
R16 a_n7097_7899.n169 a_n7097_7899.t63 168.701
R17 a_n7097_7899.n165 a_n7097_7899.t73 168.701
R18 a_n7097_7899.n166 a_n7097_7899.t26 168.701
R19 a_n7097_7899.n167 a_n7097_7899.t39 168.701
R20 a_n7097_7899.n162 a_n7097_7899.t67 168.701
R21 a_n7097_7899.n161 a_n7097_7899.t41 168.701
R22 a_n7097_7899.n152 a_n7097_7899.t18 168.701
R23 a_n7097_7899.n158 a_n7097_7899.t55 168.701
R24 a_n7097_7899.n157 a_n7097_7899.t25 168.701
R25 a_n7097_7899.n153 a_n7097_7899.t59 168.701
R26 a_n7097_7899.n154 a_n7097_7899.t40 168.701
R27 a_n7097_7899.n155 a_n7097_7899.t17 168.701
R28 a_n7097_7899.n151 a_n7097_7899.t38 168.701
R29 a_n7097_7899.n150 a_n7097_7899.t71 168.701
R30 a_n7097_7899.n141 a_n7097_7899.t50 168.701
R31 a_n7097_7899.n149 a_n7097_7899.t22 168.701
R32 a_n7097_7899.n148 a_n7097_7899.t57 168.701
R33 a_n7097_7899.n142 a_n7097_7899.t29 168.701
R34 a_n7097_7899.n143 a_n7097_7899.t68 168.701
R35 a_n7097_7899.n144 a_n7097_7899.t49 168.701
R36 a_n7097_7899.n128 a_n7097_7899.t53 168.701
R37 a_n7097_7899.n127 a_n7097_7899.t43 168.701
R38 a_n7097_7899.n126 a_n7097_7899.t28 168.701
R39 a_n7097_7899.n132 a_n7097_7899.t58 168.701
R40 a_n7097_7899.n133 a_n7097_7899.t47 168.701
R41 a_n7097_7899.n23 a_n7097_7899.t35 168.701
R42 a_n7097_7899.n135 a_n7097_7899.t24 168.701
R43 a_n7097_7899.n136 a_n7097_7899.t52 168.701
R44 a_n7097_7899.n113 a_n7097_7899.t60 168.701
R45 a_n7097_7899.n112 a_n7097_7899.t21 168.701
R46 a_n7097_7899.n111 a_n7097_7899.t44 168.701
R47 a_n7097_7899.n117 a_n7097_7899.t75 168.701
R48 a_n7097_7899.n118 a_n7097_7899.t36 168.701
R49 a_n7097_7899.n25 a_n7097_7899.t61 168.701
R50 a_n7097_7899.n120 a_n7097_7899.t23 168.701
R51 a_n7097_7899.n121 a_n7097_7899.t51 168.701
R52 a_n7097_7899.n99 a_n7097_7899.t30 168.701
R53 a_n7097_7899.n98 a_n7097_7899.t54 168.701
R54 a_n7097_7899.n97 a_n7097_7899.t72 168.701
R55 a_n7097_7899.n103 a_n7097_7899.t46 168.701
R56 a_n7097_7899.n104 a_n7097_7899.t66 168.701
R57 a_n7097_7899.n27 a_n7097_7899.t32 168.701
R58 a_n7097_7899.n106 a_n7097_7899.t56 168.701
R59 a_n7097_7899.n107 a_n7097_7899.t20 168.701
R60 a_n7097_7899.n19 a_n7097_7899.n0 39.6376
R61 a_n7097_7899.n5 a_n7097_7899.n0 39.7274
R62 a_n7097_7899.n29 a_n7097_7899.n0 68.6201
R63 a_n7097_7899.n20 a_n7097_7899.n0 39.6373
R64 a_n7097_7899.n171 a_n7097_7899.n0 161.3
R65 a_n7097_7899.n1 a_n7097_7899.n172 161.3
R66 a_n7097_7899.n21 a_n7097_7899.n1 39.7274
R67 a_n7097_7899.n22 a_n7097_7899.n1 39.6376
R68 a_n7097_7899.n15 a_n7097_7899.n2 39.6376
R69 a_n7097_7899.n6 a_n7097_7899.n2 39.7274
R70 a_n7097_7899.n30 a_n7097_7899.n2 68.6201
R71 a_n7097_7899.n16 a_n7097_7899.n2 39.6373
R72 a_n7097_7899.n159 a_n7097_7899.n2 161.3
R73 a_n7097_7899.n3 a_n7097_7899.n160 161.3
R74 a_n7097_7899.n17 a_n7097_7899.n3 39.7274
R75 a_n7097_7899.n18 a_n7097_7899.n3 39.6376
R76 a_n7097_7899.n35 a_n7097_7899.n33 71.8318
R77 a_n7097_7899.n34 a_n7097_7899.n146 161.3
R78 a_n7097_7899.n147 a_n7097_7899.n34 161.3
R79 a_n7097_7899.n32 a_n7097_7899.n7 74.8341
R80 a_n7097_7899.n31 a_n7097_7899.n4 68.6201
R81 a_n7097_7899.n12 a_n7097_7899.n4 39.6373
R82 a_n7097_7899.n4 a_n7097_7899.n8 68.6201
R83 a_n7097_7899.n13 a_n7097_7899.n4 39.7274
R84 a_n7097_7899.n14 a_n7097_7899.n4 39.6376
R85 a_n7097_7899.n137 a_n7097_7899.n53 161.3
R86 a_n7097_7899.n50 a_n7097_7899.n53 161.3
R87 a_n7097_7899.n52 a_n7097_7899.n51 71.4497
R88 a_n7097_7899.n49 a_n7097_7899.n48 68.7078
R89 a_n7097_7899.n24 a_n7097_7899.n23 11.426
R90 a_n7097_7899.n47 a_n7097_7899.n24 74.9385
R91 a_n7097_7899.n134 a_n7097_7899.n46 161.3
R92 a_n7097_7899.n43 a_n7097_7899.n46 161.3
R93 a_n7097_7899.n45 a_n7097_7899.n44 71.6402
R94 a_n7097_7899.n42 a_n7097_7899.n41 68.6201
R95 a_n7097_7899.n38 a_n7097_7899.n40 74.8341
R96 a_n7097_7899.n131 a_n7097_7899.n39 161.3
R97 a_n7097_7899.n39 a_n7097_7899.n130 161.3
R98 a_n7097_7899.n37 a_n7097_7899.n36 71.8318
R99 a_n7097_7899.n122 a_n7097_7899.n71 161.3
R100 a_n7097_7899.n68 a_n7097_7899.n71 161.3
R101 a_n7097_7899.n70 a_n7097_7899.n69 71.4497
R102 a_n7097_7899.n67 a_n7097_7899.n66 68.7078
R103 a_n7097_7899.n26 a_n7097_7899.n25 11.426
R104 a_n7097_7899.n65 a_n7097_7899.n26 74.9385
R105 a_n7097_7899.n119 a_n7097_7899.n64 161.3
R106 a_n7097_7899.n61 a_n7097_7899.n64 161.3
R107 a_n7097_7899.n63 a_n7097_7899.n62 71.6402
R108 a_n7097_7899.n60 a_n7097_7899.n59 68.6201
R109 a_n7097_7899.n56 a_n7097_7899.n58 74.8341
R110 a_n7097_7899.n116 a_n7097_7899.n57 161.3
R111 a_n7097_7899.n57 a_n7097_7899.n115 161.3
R112 a_n7097_7899.n55 a_n7097_7899.n54 71.8318
R113 a_n7097_7899.n108 a_n7097_7899.n89 161.3
R114 a_n7097_7899.n86 a_n7097_7899.n89 161.3
R115 a_n7097_7899.n88 a_n7097_7899.n87 71.4497
R116 a_n7097_7899.n85 a_n7097_7899.n84 68.7078
R117 a_n7097_7899.n28 a_n7097_7899.n27 11.426
R118 a_n7097_7899.n83 a_n7097_7899.n28 74.9385
R119 a_n7097_7899.n105 a_n7097_7899.n82 161.3
R120 a_n7097_7899.n79 a_n7097_7899.n82 161.3
R121 a_n7097_7899.n81 a_n7097_7899.n80 71.6402
R122 a_n7097_7899.n78 a_n7097_7899.n77 68.6201
R123 a_n7097_7899.n74 a_n7097_7899.n76 74.8341
R124 a_n7097_7899.n102 a_n7097_7899.n75 161.3
R125 a_n7097_7899.n75 a_n7097_7899.n101 161.3
R126 a_n7097_7899.n73 a_n7097_7899.n72 71.8318
R127 a_n7097_7899.n95 a_n7097_7899.n93 119.439
R128 a_n7097_7899.n92 a_n7097_7899.n90 119.439
R129 a_n7097_7899.n95 a_n7097_7899.n94 118.865
R130 a_n7097_7899.n92 a_n7097_7899.n91 118.865
R131 a_n7097_7899.n184 a_n7097_7899.n183 84.3504
R132 a_n7097_7899.n179 a_n7097_7899.n178 84.3502
R133 a_n7097_7899.n183 a_n7097_7899.n182 84.35
R134 a_n7097_7899.n181 a_n7097_7899.n180 84.0635
R135 a_n7097_7899.n1 a_n7097_7899.n11 43.6696
R136 a_n7097_7899.n3 a_n7097_7899.n10 43.6696
R137 a_n7097_7899.n4 a_n7097_7899.n9 43.6696
R138 a_n7097_7899.n139 a_n7097_7899.n138 80.6037
R139 a_n7097_7899.n124 a_n7097_7899.n123 80.6037
R140 a_n7097_7899.n110 a_n7097_7899.n109 80.6037
R141 a_n7097_7899.n172 a_n7097_7899.n171 56.5617
R142 a_n7097_7899.n29 a_n7097_7899.n165 48.4088
R143 a_n7097_7899.n160 a_n7097_7899.n159 56.5617
R144 a_n7097_7899.n30 a_n7097_7899.n153 48.4088
R145 a_n7097_7899.n31 a_n7097_7899.n142 48.4088
R146 a_n7097_7899.n132 a_n7097_7899.n42 40.5394
R147 a_n7097_7899.n24 a_n7097_7899.n134 67.9872
R148 a_n7097_7899.n117 a_n7097_7899.n60 40.5394
R149 a_n7097_7899.n26 a_n7097_7899.n119 67.9872
R150 a_n7097_7899.n103 a_n7097_7899.n78 40.5394
R151 a_n7097_7899.n28 a_n7097_7899.n105 67.9872
R152 a_n7097_7899.n173 a_n7097_7899.n21 51.9316
R153 a_n7097_7899.n161 a_n7097_7899.n17 51.9316
R154 a_n7097_7899.n150 a_n7097_7899.n13 51.9316
R155 a_n7097_7899.n40 a_n7097_7899.n131 67.7116
R156 a_n7097_7899.n135 a_n7097_7899.n49 39.872
R157 a_n7097_7899.n58 a_n7097_7899.n116 67.7116
R158 a_n7097_7899.n120 a_n7097_7899.n67 39.872
R159 a_n7097_7899.n76 a_n7097_7899.n102 67.7116
R160 a_n7097_7899.n106 a_n7097_7899.n85 39.872
R161 a_n7097_7899.n138 a_n7097_7899.n137 55.824
R162 a_n7097_7899.n123 a_n7097_7899.n122 55.824
R163 a_n7097_7899.n109 a_n7097_7899.n108 55.824
R164 a_n7097_7899.n168 a_n7097_7899.n167 47.1841
R165 a_n7097_7899.n156 a_n7097_7899.n155 47.1841
R166 a_n7097_7899.n145 a_n7097_7899.n144 47.1841
R167 a_n7097_7899.n129 a_n7097_7899.n128 47.1841
R168 a_n7097_7899.n114 a_n7097_7899.n113 47.1841
R169 a_n7097_7899.n100 a_n7097_7899.n99 47.1841
R170 a_n7097_7899.n36 a_n7097_7899.n129 43.9713
R171 a_n7097_7899.n54 a_n7097_7899.n114 43.9713
R172 a_n7097_7899.n72 a_n7097_7899.n100 43.9713
R173 a_n7097_7899.n0 a_n7097_7899.n168 43.9713
R174 a_n7097_7899.n2 a_n7097_7899.n156 43.9713
R175 a_n7097_7899.n33 a_n7097_7899.n145 43.9713
R176 a_n7097_7899.n173 a_n7097_7899.n22 41.2665
R177 a_n7097_7899.n161 a_n7097_7899.n18 41.2665
R178 a_n7097_7899.n150 a_n7097_7899.n14 41.2665
R179 a_n7097_7899.n146 a_n7097_7899.n35 59.1846
R180 a_n7097_7899.n130 a_n7097_7899.n37 59.1846
R181 a_n7097_7899.n51 a_n7097_7899.n50 58.0115
R182 a_n7097_7899.n115 a_n7097_7899.n55 59.1846
R183 a_n7097_7899.n69 a_n7097_7899.n68 58.0115
R184 a_n7097_7899.n101 a_n7097_7899.n73 59.1846
R185 a_n7097_7899.n87 a_n7097_7899.n86 58.0115
R186 a_n7097_7899.n169 a_n7097_7899.n20 40.5378
R187 a_n7097_7899.n157 a_n7097_7899.n16 40.5378
R188 a_n7097_7899.n148 a_n7097_7899.n12 40.5378
R189 a_n7097_7899.n44 a_n7097_7899.n43 58.5991
R190 a_n7097_7899.n62 a_n7097_7899.n61 58.5991
R191 a_n7097_7899.n80 a_n7097_7899.n79 58.5991
R192 a_n7097_7899.n19 a_n7097_7899.n167 39.8067
R193 a_n7097_7899.n15 a_n7097_7899.n155 39.8067
R194 a_n7097_7899.n35 a_n7097_7899.n144 25.2628
R195 a_n7097_7899.n183 a_n7097_7899.n181 30.5791
R196 a_n7097_7899.n96 a_n7097_7899.n92 25.6013
R197 a_n7097_7899.n5 a_n7097_7899.n166 51.931
R198 a_n7097_7899.n6 a_n7097_7899.n154 51.931
R199 a_n7097_7899.n32 a_n7097_7899.n147 67.7116
R200 a_n7097_7899.n126 a_n7097_7899.n40 11.8807
R201 a_n7097_7899.n49 a_n7097_7899.n23 48.9635
R202 a_n7097_7899.n111 a_n7097_7899.n58 11.8807
R203 a_n7097_7899.n67 a_n7097_7899.n25 48.9635
R204 a_n7097_7899.n97 a_n7097_7899.n76 11.8807
R205 a_n7097_7899.n85 a_n7097_7899.n27 48.9635
R206 a_n7097_7899.n172 a_n7097_7899.n164 24.3464
R207 a_n7097_7899.n160 a_n7097_7899.n152 24.3464
R208 a_n7097_7899.n8 a_n7097_7899.n141 48.4088
R209 a_n7097_7899.n42 a_n7097_7899.n126 48.4088
R210 a_n7097_7899.n60 a_n7097_7899.n111 48.4088
R211 a_n7097_7899.n78 a_n7097_7899.n97 48.4088
R212 a_n7097_7899.n11 a_n7097_7899.n174 47.213
R213 a_n7097_7899.n10 a_n7097_7899.n162 47.213
R214 a_n7097_7899.n9 a_n7097_7899.n151 47.213
R215 a_n7097_7899.n137 a_n7097_7899.n136 16.9689
R216 a_n7097_7899.n122 a_n7097_7899.n121 16.9689
R217 a_n7097_7899.n108 a_n7097_7899.n107 16.9689
R218 a_n7097_7899.n96 a_n7097_7899.n95 16.7274
R219 a_n7097_7899.n171 a_n7097_7899.n170 16.477
R220 a_n7097_7899.n169 a_n7097_7899.n29 40.5394
R221 a_n7097_7899.n159 a_n7097_7899.n158 16.477
R222 a_n7097_7899.n157 a_n7097_7899.n30 40.5394
R223 a_n7097_7899.n8 a_n7097_7899.n149 40.5394
R224 a_n7097_7899.n148 a_n7097_7899.n31 40.5394
R225 a_n7097_7899.n134 a_n7097_7899.n133 16.477
R226 a_n7097_7899.n119 a_n7097_7899.n118 16.477
R227 a_n7097_7899.n105 a_n7097_7899.n104 16.477
R228 a_n7097_7899.n147 a_n7097_7899.n143 15.9852
R229 a_n7097_7899.n131 a_n7097_7899.n127 15.9852
R230 a_n7097_7899.n116 a_n7097_7899.n112 15.9852
R231 a_n7097_7899.n102 a_n7097_7899.n98 15.9852
R232 a_n7097_7899.n179 a_n7097_7899.n177 12.3788
R233 a_n7097_7899.n177 a_n7097_7899.n96 11.5231
R234 a_n7097_7899.n163 a_n7097_7899.n4 8.76042
R235 a_n7097_7899.n125 a_n7097_7899.n110 8.76042
R236 a_n7097_7899.n19 a_n7097_7899.n166 41.266
R237 a_n7097_7899.n15 a_n7097_7899.n154 41.266
R238 a_n7097_7899.n146 a_n7097_7899.n143 8.60764
R239 a_n7097_7899.n130 a_n7097_7899.n127 8.60764
R240 a_n7097_7899.n51 a_n7097_7899.n135 27.0108
R241 a_n7097_7899.n115 a_n7097_7899.n112 8.60764
R242 a_n7097_7899.n69 a_n7097_7899.n120 27.0108
R243 a_n7097_7899.n101 a_n7097_7899.n98 8.60764
R244 a_n7097_7899.n87 a_n7097_7899.n106 27.0108
R245 a_n7097_7899.n170 a_n7097_7899.n20 40.5373
R246 a_n7097_7899.n158 a_n7097_7899.n16 40.5373
R247 a_n7097_7899.n149 a_n7097_7899.n12 40.5373
R248 a_n7097_7899.n44 a_n7097_7899.n132 26.1378
R249 a_n7097_7899.n133 a_n7097_7899.n43 8.11581
R250 a_n7097_7899.n62 a_n7097_7899.n117 26.1378
R251 a_n7097_7899.n118 a_n7097_7899.n61 8.11581
R252 a_n7097_7899.n80 a_n7097_7899.n103 26.1378
R253 a_n7097_7899.n104 a_n7097_7899.n79 8.11581
R254 a_n7097_7899.n174 a_n7097_7899.n22 39.8062
R255 a_n7097_7899.n162 a_n7097_7899.n18 39.8062
R256 a_n7097_7899.n151 a_n7097_7899.n14 39.8062
R257 a_n7097_7899.n37 a_n7097_7899.n128 25.2628
R258 a_n7097_7899.n136 a_n7097_7899.n50 7.62397
R259 a_n7097_7899.n55 a_n7097_7899.n113 25.2628
R260 a_n7097_7899.n121 a_n7097_7899.n68 7.62397
R261 a_n7097_7899.n73 a_n7097_7899.n99 25.2628
R262 a_n7097_7899.n107 a_n7097_7899.n86 7.62397
R263 a_n7097_7899.n94 a_n7097_7899.t5 6.5015
R264 a_n7097_7899.n94 a_n7097_7899.t11 6.5015
R265 a_n7097_7899.n93 a_n7097_7899.t2 6.5015
R266 a_n7097_7899.n93 a_n7097_7899.t12 6.5015
R267 a_n7097_7899.n90 a_n7097_7899.t4 6.5015
R268 a_n7097_7899.n90 a_n7097_7899.t13 6.5015
R269 a_n7097_7899.n91 a_n7097_7899.t14 6.5015
R270 a_n7097_7899.n91 a_n7097_7899.t0 6.5015
R271 a_n7097_7899.n176 a_n7097_7899.n140 5.3373
R272 a_n7097_7899.n176 a_n7097_7899.n175 5.13645
R273 a_n7097_7899.n175 a_n7097_7899.n1 5.06913
R274 a_n7097_7899.n163 a_n7097_7899.n3 5.06913
R275 a_n7097_7899.n140 a_n7097_7899.n139 5.06913
R276 a_n7097_7899.n125 a_n7097_7899.n124 5.06913
R277 a_n7097_7899.n175 a_n7097_7899.n163 3.69179
R278 a_n7097_7899.n140 a_n7097_7899.n125 3.69179
R279 a_n7097_7899.n177 a_n7097_7899.n176 3.4105
R280 a_n7097_7899.n182 a_n7097_7899.t8 3.3005
R281 a_n7097_7899.n182 a_n7097_7899.t10 3.3005
R282 a_n7097_7899.n180 a_n7097_7899.t7 3.3005
R283 a_n7097_7899.n180 a_n7097_7899.t6 3.3005
R284 a_n7097_7899.n178 a_n7097_7899.t9 3.3005
R285 a_n7097_7899.n178 a_n7097_7899.t3 3.3005
R286 a_n7097_7899.n184 a_n7097_7899.t15 3.3005
R287 a_n7097_7899.t1 a_n7097_7899.n184 3.3005
R288 a_n7097_7899.n75 a_n7097_7899.n72 0.568682
R289 a_n7097_7899.n57 a_n7097_7899.n54 0.568682
R290 a_n7097_7899.n39 a_n7097_7899.n36 0.568682
R291 a_n7097_7899.n89 a_n7097_7899.n88 0.379288
R292 a_n7097_7899.n88 a_n7097_7899.n84 0.379288
R293 a_n7097_7899.n84 a_n7097_7899.n83 0.379288
R294 a_n7097_7899.n83 a_n7097_7899.n82 0.379288
R295 a_n7097_7899.n82 a_n7097_7899.n81 0.379288
R296 a_n7097_7899.n81 a_n7097_7899.n77 0.379288
R297 a_n7097_7899.n77 a_n7097_7899.n74 0.379288
R298 a_n7097_7899.n75 a_n7097_7899.n74 0.379288
R299 a_n7097_7899.n71 a_n7097_7899.n70 0.379288
R300 a_n7097_7899.n70 a_n7097_7899.n66 0.379288
R301 a_n7097_7899.n66 a_n7097_7899.n65 0.379288
R302 a_n7097_7899.n65 a_n7097_7899.n64 0.379288
R303 a_n7097_7899.n64 a_n7097_7899.n63 0.379288
R304 a_n7097_7899.n63 a_n7097_7899.n59 0.379288
R305 a_n7097_7899.n59 a_n7097_7899.n56 0.379288
R306 a_n7097_7899.n57 a_n7097_7899.n56 0.379288
R307 a_n7097_7899.n53 a_n7097_7899.n52 0.379288
R308 a_n7097_7899.n52 a_n7097_7899.n48 0.379288
R309 a_n7097_7899.n48 a_n7097_7899.n47 0.379288
R310 a_n7097_7899.n47 a_n7097_7899.n46 0.379288
R311 a_n7097_7899.n46 a_n7097_7899.n45 0.379288
R312 a_n7097_7899.n45 a_n7097_7899.n41 0.379288
R313 a_n7097_7899.n41 a_n7097_7899.n38 0.379288
R314 a_n7097_7899.n39 a_n7097_7899.n38 0.379288
R315 a_n7097_7899.n34 a_n7097_7899.n33 0.379288
R316 a_n7097_7899.n34 a_n7097_7899.n7 0.379288
R317 a_n7097_7899.n181 a_n7097_7899.n179 0.287138
R318 a_n7097_7899.n139 a_n7097_7899.n53 0.285035
R319 a_n7097_7899.n124 a_n7097_7899.n71 0.285035
R320 a_n7097_7899.n110 a_n7097_7899.n89 0.285035
R321 a_n7097_7899.n164 a_n7097_7899.n21 28.5572
R322 a_n7097_7899.n5 a_n7097_7899.n165 28.5577
R323 a_n7097_7899.n152 a_n7097_7899.n17 28.5572
R324 a_n7097_7899.n6 a_n7097_7899.n153 28.5577
R325 a_n7097_7899.n141 a_n7097_7899.n13 28.5572
R326 a_n7097_7899.n32 a_n7097_7899.n142 11.8807
R327 a_n7097_7899.n3 a_n7097_7899.n2 3.88352
R328 a_n7097_7899.n1 a_n7097_7899.n0 3.88352
R329 a_n7097_7899.n4 a_n7097_7899.n7 3.12594
R330 VDD.n2275 VDD.n270 452.195
R331 VDD.n2489 VDD.n99 452.195
R332 VDD.n2382 VDD.n97 452.195
R333 VDD.n302 VDD.n268 452.195
R334 VDD.n1485 VDD.n648 452.195
R335 VDD.n1487 VDD.n637 452.195
R336 VDD.n818 VDD.n784 452.195
R337 VDD.n995 VDD.n786 452.195
R338 VDD.n900 VDD.t40 371.625
R339 VDD.n933 VDD.t32 371.625
R340 VDD.n966 VDD.t67 371.625
R341 VDD.n1492 VDD.t29 371.625
R342 VDD.n1207 VDD.t60 371.625
R343 VDD.n1172 VDD.t21 371.625
R344 VDD.n199 VDD.t57 371.625
R345 VDD.n166 VDD.t88 371.625
R346 VDD.n131 VDD.t50 371.625
R347 VDD.n340 VDD.t43 371.625
R348 VDD.n2242 VDD.t74 371.625
R349 VDD.n2159 VDD.t54 371.625
R350 VDD.n1348 VDD.t70 323.425
R351 VDD.n525 VDD.t63 323.425
R352 VDD.n1333 VDD.t94 323.425
R353 VDD.n509 VDD.t91 323.425
R354 VDD.n2027 VDD.t81 323.425
R355 VDD.n1790 VDD.t85 323.425
R356 VDD.n388 VDD.t47 323.425
R357 VDD.n1762 VDD.t77 323.425
R358 VDD.n360 VDD.t36 323.425
R359 VDD.n617 VDD.t25 323.425
R360 VDD.n2116 VDD.n372 305.854
R361 VDD.n2077 VDD.n2076 305.854
R362 VDD.n1902 VDD.n1901 305.854
R363 VDD.n1946 VDD.n479 305.854
R364 VDD.n1737 VDD.n506 305.854
R365 VDD.n1692 VDD.n1691 305.854
R366 VDD.n1443 VDD.n614 305.854
R367 VDD.n1533 VDD.n612 305.854
R368 VDD.n2054 VDD.n2053 305.854
R369 VDD.n2126 VDD.n364 305.854
R370 VDD.n1838 VDD.n1760 305.854
R371 VDD.n1793 VDD.n475 305.854
R372 VDD.n1677 VDD.n1676 305.854
R373 VDD.n1630 VDD.n494 305.854
R374 VDD.n1372 VDD.n615 305.854
R375 VDD.n1531 VDD.n616 305.854
R376 VDD.n2055 VDD.n2054 185
R377 VDD.n2054 VDD.n369 185
R378 VDD.n2056 VDD.n370 185
R379 VDD.n2121 VDD.n370 185
R380 VDD.n2058 VDD.n2057 185
R381 VDD.n2057 VDD.n367 185
R382 VDD.n2059 VDD.n394 185
R383 VDD.n2069 VDD.n394 185
R384 VDD.n2060 VDD.n402 185
R385 VDD.n1854 VDD.n402 185
R386 VDD.n2062 VDD.n2061 185
R387 VDD.n2063 VDD.n2062 185
R388 VDD.n2026 VDD.n401 185
R389 VDD.n401 VDD.n398 185
R390 VDD.n2025 VDD.n2024 185
R391 VDD.n2024 VDD.n2023 185
R392 VDD.n404 VDD.n403 185
R393 VDD.n405 VDD.n404 185
R394 VDD.n2016 VDD.n2015 185
R395 VDD.n2017 VDD.n2016 185
R396 VDD.n2014 VDD.n414 185
R397 VDD.n414 VDD.n411 185
R398 VDD.n2013 VDD.n2012 185
R399 VDD.n2012 VDD.n2011 185
R400 VDD.n416 VDD.n415 185
R401 VDD.n417 VDD.n416 185
R402 VDD.n2004 VDD.n2003 185
R403 VDD.n2005 VDD.n2004 185
R404 VDD.n2002 VDD.n426 185
R405 VDD.n426 VDD.n423 185
R406 VDD.n2001 VDD.n2000 185
R407 VDD.n2000 VDD.n1999 185
R408 VDD.n428 VDD.n427 185
R409 VDD.n429 VDD.n428 185
R410 VDD.n1992 VDD.n1991 185
R411 VDD.n1993 VDD.n1992 185
R412 VDD.n1990 VDD.n437 185
R413 VDD.n443 VDD.n437 185
R414 VDD.n1989 VDD.n1988 185
R415 VDD.n1988 VDD.n1987 185
R416 VDD.n439 VDD.n438 185
R417 VDD.n440 VDD.n439 185
R418 VDD.n1980 VDD.n1979 185
R419 VDD.n1981 VDD.n1980 185
R420 VDD.n1978 VDD.n449 185
R421 VDD.n1884 VDD.n449 185
R422 VDD.n1977 VDD.n1976 185
R423 VDD.n1976 VDD.n1975 185
R424 VDD.n451 VDD.n450 185
R425 VDD.n452 VDD.n451 185
R426 VDD.n1968 VDD.n1967 185
R427 VDD.n1969 VDD.n1968 185
R428 VDD.n1966 VDD.n461 185
R429 VDD.n461 VDD.n458 185
R430 VDD.n1965 VDD.n1964 185
R431 VDD.n1964 VDD.n1963 185
R432 VDD.n463 VDD.n462 185
R433 VDD.n464 VDD.n463 185
R434 VDD.n1956 VDD.n1955 185
R435 VDD.n1957 VDD.n1956 185
R436 VDD.n1954 VDD.n473 185
R437 VDD.n473 VDD.n470 185
R438 VDD.n1953 VDD.n1952 185
R439 VDD.n1952 VDD.n1951 185
R440 VDD.n475 VDD.n474 185
R441 VDD.n476 VDD.n475 185
R442 VDD.n1794 VDD.n1793 185
R443 VDD.n1796 VDD.n1795 185
R444 VDD.n1798 VDD.n1797 185
R445 VDD.n1800 VDD.n1799 185
R446 VDD.n1802 VDD.n1801 185
R447 VDD.n1804 VDD.n1803 185
R448 VDD.n1806 VDD.n1805 185
R449 VDD.n1808 VDD.n1807 185
R450 VDD.n1810 VDD.n1809 185
R451 VDD.n1812 VDD.n1811 185
R452 VDD.n1814 VDD.n1813 185
R453 VDD.n1816 VDD.n1815 185
R454 VDD.n1818 VDD.n1817 185
R455 VDD.n1820 VDD.n1819 185
R456 VDD.n1822 VDD.n1821 185
R457 VDD.n1824 VDD.n1823 185
R458 VDD.n1826 VDD.n1825 185
R459 VDD.n1828 VDD.n1827 185
R460 VDD.n1830 VDD.n1829 185
R461 VDD.n1832 VDD.n1831 185
R462 VDD.n1834 VDD.n1833 185
R463 VDD.n1836 VDD.n1835 185
R464 VDD.n1837 VDD.n1760 185
R465 VDD.n1944 VDD.n1760 185
R466 VDD.n2126 VDD.n2125 185
R467 VDD.n2128 VDD.n362 185
R468 VDD.n2130 VDD.n2129 185
R469 VDD.n2132 VDD.n359 185
R470 VDD.n2134 VDD.n2133 185
R471 VDD.n2136 VDD.n357 185
R472 VDD.n2138 VDD.n2137 185
R473 VDD.n2139 VDD.n356 185
R474 VDD.n2141 VDD.n2140 185
R475 VDD.n2143 VDD.n355 185
R476 VDD.n2144 VDD.n352 185
R477 VDD.n2147 VDD.n2146 185
R478 VDD.n353 VDD.n351 185
R479 VDD.n2037 VDD.n2036 185
R480 VDD.n2039 VDD.n2038 185
R481 VDD.n2041 VDD.n2033 185
R482 VDD.n2043 VDD.n2042 185
R483 VDD.n2044 VDD.n2032 185
R484 VDD.n2046 VDD.n2045 185
R485 VDD.n2048 VDD.n2030 185
R486 VDD.n2050 VDD.n2049 185
R487 VDD.n2051 VDD.n2029 185
R488 VDD.n2053 VDD.n2052 185
R489 VDD.n2053 VDD.n354 185
R490 VDD.n2124 VDD.n364 185
R491 VDD.n369 VDD.n364 185
R492 VDD.n2123 VDD.n2122 185
R493 VDD.n2122 VDD.n2121 185
R494 VDD.n366 VDD.n365 185
R495 VDD.n367 VDD.n366 185
R496 VDD.n1853 VDD.n393 185
R497 VDD.n2069 VDD.n393 185
R498 VDD.n1856 VDD.n1855 185
R499 VDD.n1855 VDD.n1854 185
R500 VDD.n1857 VDD.n400 185
R501 VDD.n2063 VDD.n400 185
R502 VDD.n1859 VDD.n1858 185
R503 VDD.n1858 VDD.n398 185
R504 VDD.n1860 VDD.n407 185
R505 VDD.n2023 VDD.n407 185
R506 VDD.n1862 VDD.n1861 185
R507 VDD.n1861 VDD.n405 185
R508 VDD.n1863 VDD.n413 185
R509 VDD.n2017 VDD.n413 185
R510 VDD.n1865 VDD.n1864 185
R511 VDD.n1864 VDD.n411 185
R512 VDD.n1866 VDD.n419 185
R513 VDD.n2011 VDD.n419 185
R514 VDD.n1868 VDD.n1867 185
R515 VDD.n1867 VDD.n417 185
R516 VDD.n1869 VDD.n425 185
R517 VDD.n2005 VDD.n425 185
R518 VDD.n1871 VDD.n1870 185
R519 VDD.n1870 VDD.n423 185
R520 VDD.n1872 VDD.n431 185
R521 VDD.n1999 VDD.n431 185
R522 VDD.n1874 VDD.n1873 185
R523 VDD.n1873 VDD.n429 185
R524 VDD.n1875 VDD.n436 185
R525 VDD.n1993 VDD.n436 185
R526 VDD.n1877 VDD.n1876 185
R527 VDD.n1876 VDD.n443 185
R528 VDD.n1878 VDD.n442 185
R529 VDD.n1987 VDD.n442 185
R530 VDD.n1880 VDD.n1879 185
R531 VDD.n1879 VDD.n440 185
R532 VDD.n1881 VDD.n448 185
R533 VDD.n1981 VDD.n448 185
R534 VDD.n1883 VDD.n1882 185
R535 VDD.n1884 VDD.n1883 185
R536 VDD.n1852 VDD.n454 185
R537 VDD.n1975 VDD.n454 185
R538 VDD.n1851 VDD.n1850 185
R539 VDD.n1850 VDD.n452 185
R540 VDD.n1849 VDD.n460 185
R541 VDD.n1969 VDD.n460 185
R542 VDD.n1848 VDD.n1847 185
R543 VDD.n1847 VDD.n458 185
R544 VDD.n1846 VDD.n466 185
R545 VDD.n1963 VDD.n466 185
R546 VDD.n1845 VDD.n1844 185
R547 VDD.n1844 VDD.n464 185
R548 VDD.n1843 VDD.n472 185
R549 VDD.n1957 VDD.n472 185
R550 VDD.n1842 VDD.n1841 185
R551 VDD.n1841 VDD.n470 185
R552 VDD.n1840 VDD.n478 185
R553 VDD.n1951 VDD.n478 185
R554 VDD.n1839 VDD.n1838 185
R555 VDD.n1838 VDD.n476 185
R556 VDD.n508 VDD.n506 185
R557 VDD.n506 VDD.n482 185
R558 VDD.n1688 VDD.n1687 185
R559 VDD.n1689 VDD.n1688 185
R560 VDD.n1686 VDD.n516 185
R561 VDD.n521 VDD.n516 185
R562 VDD.n1685 VDD.n1684 185
R563 VDD.n1684 VDD.n1683 185
R564 VDD.n518 VDD.n517 185
R565 VDD.n1623 VDD.n518 185
R566 VDD.n1612 VDD.n538 185
R567 VDD.n538 VDD.n530 185
R568 VDD.n1614 VDD.n1613 185
R569 VDD.n1615 VDD.n1614 185
R570 VDD.n1611 VDD.n537 185
R571 VDD.n537 VDD.n534 185
R572 VDD.n1610 VDD.n1609 185
R573 VDD.n1609 VDD.n1608 185
R574 VDD.n540 VDD.n539 185
R575 VDD.n541 VDD.n540 185
R576 VDD.n1597 VDD.n1596 185
R577 VDD.n1598 VDD.n1597 185
R578 VDD.n1595 VDD.n550 185
R579 VDD.n556 VDD.n550 185
R580 VDD.n1594 VDD.n1593 185
R581 VDD.n1593 VDD.n1592 185
R582 VDD.n552 VDD.n551 185
R583 VDD.n553 VDD.n552 185
R584 VDD.n1585 VDD.n1584 185
R585 VDD.n1586 VDD.n1585 185
R586 VDD.n1583 VDD.n562 185
R587 VDD.n1414 VDD.n562 185
R588 VDD.n1582 VDD.n1581 185
R589 VDD.n1581 VDD.n1580 185
R590 VDD.n564 VDD.n563 185
R591 VDD.n565 VDD.n564 185
R592 VDD.n1573 VDD.n1572 185
R593 VDD.n1574 VDD.n1573 185
R594 VDD.n1571 VDD.n574 185
R595 VDD.n574 VDD.n571 185
R596 VDD.n1570 VDD.n1569 185
R597 VDD.n1569 VDD.n1568 185
R598 VDD.n576 VDD.n575 185
R599 VDD.n577 VDD.n576 185
R600 VDD.n1561 VDD.n1560 185
R601 VDD.n1562 VDD.n1561 185
R602 VDD.n1559 VDD.n586 185
R603 VDD.n586 VDD.n583 185
R604 VDD.n1558 VDD.n1557 185
R605 VDD.n1557 VDD.n1556 185
R606 VDD.n588 VDD.n587 185
R607 VDD.n589 VDD.n588 185
R608 VDD.n1549 VDD.n1548 185
R609 VDD.n1550 VDD.n1549 185
R610 VDD.n1547 VDD.n598 185
R611 VDD.n598 VDD.n595 185
R612 VDD.n1546 VDD.n1545 185
R613 VDD.n1545 VDD.n1544 185
R614 VDD.n600 VDD.n599 185
R615 VDD.n609 VDD.n600 185
R616 VDD.n1537 VDD.n1536 185
R617 VDD.n1538 VDD.n1537 185
R618 VDD.n1535 VDD.n610 185
R619 VDD.n610 VDD.n606 185
R620 VDD.n1534 VDD.n1533 185
R621 VDD.n1533 VDD.n1532 185
R622 VDD.n612 VDD.n611 185
R623 VDD.n1310 VDD.n1308 185
R624 VDD.n1311 VDD.n1307 185
R625 VDD.n1311 VDD.n613 185
R626 VDD.n1314 VDD.n1313 185
R627 VDD.n1315 VDD.n1306 185
R628 VDD.n1317 VDD.n1316 185
R629 VDD.n1319 VDD.n1305 185
R630 VDD.n1322 VDD.n1321 185
R631 VDD.n1323 VDD.n1304 185
R632 VDD.n1325 VDD.n1324 185
R633 VDD.n1327 VDD.n1302 185
R634 VDD.n1465 VDD.n1464 185
R635 VDD.n1462 VDD.n1303 185
R636 VDD.n1461 VDD.n1460 185
R637 VDD.n1459 VDD.n1458 185
R638 VDD.n1457 VDD.n1329 185
R639 VDD.n1455 VDD.n1454 185
R640 VDD.n1453 VDD.n1330 185
R641 VDD.n1452 VDD.n1451 185
R642 VDD.n1449 VDD.n1331 185
R643 VDD.n1447 VDD.n1446 185
R644 VDD.n1445 VDD.n1332 185
R645 VDD.n1444 VDD.n1443 185
R646 VDD.n1693 VDD.n1692 185
R647 VDD.n1695 VDD.n1694 185
R648 VDD.n1697 VDD.n1696 185
R649 VDD.n1700 VDD.n1699 185
R650 VDD.n1702 VDD.n1701 185
R651 VDD.n1704 VDD.n1703 185
R652 VDD.n1706 VDD.n1705 185
R653 VDD.n1708 VDD.n1707 185
R654 VDD.n1710 VDD.n1709 185
R655 VDD.n1712 VDD.n1711 185
R656 VDD.n1714 VDD.n1713 185
R657 VDD.n1716 VDD.n1715 185
R658 VDD.n1718 VDD.n1717 185
R659 VDD.n1720 VDD.n1719 185
R660 VDD.n1722 VDD.n1721 185
R661 VDD.n1724 VDD.n1723 185
R662 VDD.n1726 VDD.n1725 185
R663 VDD.n1728 VDD.n1727 185
R664 VDD.n1730 VDD.n1729 185
R665 VDD.n1732 VDD.n1731 185
R666 VDD.n1734 VDD.n1733 185
R667 VDD.n1735 VDD.n507 185
R668 VDD.n1737 VDD.n1736 185
R669 VDD.n1738 VDD.n1737 185
R670 VDD.n1691 VDD.n511 185
R671 VDD.n1691 VDD.n482 185
R672 VDD.n1690 VDD.n513 185
R673 VDD.n1690 VDD.n1689 185
R674 VDD.n1619 VDD.n512 185
R675 VDD.n521 VDD.n512 185
R676 VDD.n1620 VDD.n519 185
R677 VDD.n1683 VDD.n519 185
R678 VDD.n1622 VDD.n1621 185
R679 VDD.n1623 VDD.n1622 185
R680 VDD.n1618 VDD.n531 185
R681 VDD.n531 VDD.n530 185
R682 VDD.n1617 VDD.n1616 185
R683 VDD.n1616 VDD.n1615 185
R684 VDD.n533 VDD.n532 185
R685 VDD.n534 VDD.n533 185
R686 VDD.n1336 VDD.n542 185
R687 VDD.n1608 VDD.n542 185
R688 VDD.n1338 VDD.n1337 185
R689 VDD.n1337 VDD.n541 185
R690 VDD.n1339 VDD.n548 185
R691 VDD.n1598 VDD.n548 185
R692 VDD.n1341 VDD.n1340 185
R693 VDD.n1340 VDD.n556 185
R694 VDD.n1342 VDD.n554 185
R695 VDD.n1592 VDD.n554 185
R696 VDD.n1344 VDD.n1343 185
R697 VDD.n1343 VDD.n553 185
R698 VDD.n1345 VDD.n560 185
R699 VDD.n1586 VDD.n560 185
R700 VDD.n1416 VDD.n1415 185
R701 VDD.n1415 VDD.n1414 185
R702 VDD.n1417 VDD.n566 185
R703 VDD.n1580 VDD.n566 185
R704 VDD.n1419 VDD.n1418 185
R705 VDD.n1418 VDD.n565 185
R706 VDD.n1420 VDD.n572 185
R707 VDD.n1574 VDD.n572 185
R708 VDD.n1422 VDD.n1421 185
R709 VDD.n1421 VDD.n571 185
R710 VDD.n1423 VDD.n578 185
R711 VDD.n1568 VDD.n578 185
R712 VDD.n1425 VDD.n1424 185
R713 VDD.n1424 VDD.n577 185
R714 VDD.n1426 VDD.n584 185
R715 VDD.n1562 VDD.n584 185
R716 VDD.n1428 VDD.n1427 185
R717 VDD.n1427 VDD.n583 185
R718 VDD.n1429 VDD.n590 185
R719 VDD.n1556 VDD.n590 185
R720 VDD.n1431 VDD.n1430 185
R721 VDD.n1430 VDD.n589 185
R722 VDD.n1432 VDD.n596 185
R723 VDD.n1550 VDD.n596 185
R724 VDD.n1434 VDD.n1433 185
R725 VDD.n1433 VDD.n595 185
R726 VDD.n1435 VDD.n601 185
R727 VDD.n1544 VDD.n601 185
R728 VDD.n1437 VDD.n1436 185
R729 VDD.n1436 VDD.n609 185
R730 VDD.n1438 VDD.n607 185
R731 VDD.n1538 VDD.n607 185
R732 VDD.n1440 VDD.n1439 185
R733 VDD.n1439 VDD.n606 185
R734 VDD.n1441 VDD.n614 185
R735 VDD.n1532 VDD.n614 185
R736 VDD.n2118 VDD.n372 185
R737 VDD.n372 VDD.n369 185
R738 VDD.n2120 VDD.n2119 185
R739 VDD.n2121 VDD.n2120 185
R740 VDD.n373 VDD.n371 185
R741 VDD.n371 VDD.n367 185
R742 VDD.n2068 VDD.n2067 185
R743 VDD.n2069 VDD.n2068 185
R744 VDD.n2066 VDD.n395 185
R745 VDD.n1854 VDD.n395 185
R746 VDD.n2065 VDD.n2064 185
R747 VDD.n2064 VDD.n2063 185
R748 VDD.n397 VDD.n396 185
R749 VDD.n398 VDD.n397 185
R750 VDD.n2022 VDD.n2021 185
R751 VDD.n2023 VDD.n2022 185
R752 VDD.n2020 VDD.n408 185
R753 VDD.n408 VDD.n405 185
R754 VDD.n2019 VDD.n2018 185
R755 VDD.n2018 VDD.n2017 185
R756 VDD.n410 VDD.n409 185
R757 VDD.n411 VDD.n410 185
R758 VDD.n2010 VDD.n2009 185
R759 VDD.n2011 VDD.n2010 185
R760 VDD.n2008 VDD.n420 185
R761 VDD.n420 VDD.n417 185
R762 VDD.n2007 VDD.n2006 185
R763 VDD.n2006 VDD.n2005 185
R764 VDD.n422 VDD.n421 185
R765 VDD.n423 VDD.n422 185
R766 VDD.n1998 VDD.n1997 185
R767 VDD.n1999 VDD.n1998 185
R768 VDD.n1996 VDD.n432 185
R769 VDD.n432 VDD.n429 185
R770 VDD.n1995 VDD.n1994 185
R771 VDD.n1994 VDD.n1993 185
R772 VDD.n434 VDD.n433 185
R773 VDD.n443 VDD.n434 185
R774 VDD.n1986 VDD.n1985 185
R775 VDD.n1987 VDD.n1986 185
R776 VDD.n1984 VDD.n444 185
R777 VDD.n444 VDD.n440 185
R778 VDD.n1983 VDD.n1982 185
R779 VDD.n1982 VDD.n1981 185
R780 VDD.n446 VDD.n445 185
R781 VDD.n1884 VDD.n446 185
R782 VDD.n1974 VDD.n1973 185
R783 VDD.n1975 VDD.n1974 185
R784 VDD.n1972 VDD.n455 185
R785 VDD.n455 VDD.n452 185
R786 VDD.n1971 VDD.n1970 185
R787 VDD.n1970 VDD.n1969 185
R788 VDD.n457 VDD.n456 185
R789 VDD.n458 VDD.n457 185
R790 VDD.n1962 VDD.n1961 185
R791 VDD.n1963 VDD.n1962 185
R792 VDD.n1960 VDD.n467 185
R793 VDD.n467 VDD.n464 185
R794 VDD.n1959 VDD.n1958 185
R795 VDD.n1958 VDD.n1957 185
R796 VDD.n469 VDD.n468 185
R797 VDD.n470 VDD.n469 185
R798 VDD.n1950 VDD.n1949 185
R799 VDD.n1951 VDD.n1950 185
R800 VDD.n1948 VDD.n479 185
R801 VDD.n479 VDD.n476 185
R802 VDD.n1947 VDD.n1946 185
R803 VDD.n481 VDD.n480 185
R804 VDD.n1943 VDD.n1942 185
R805 VDD.n1944 VDD.n1943 185
R806 VDD.n1941 VDD.n1761 185
R807 VDD.n1940 VDD.n1939 185
R808 VDD.n1938 VDD.n1937 185
R809 VDD.n1936 VDD.n1935 185
R810 VDD.n1934 VDD.n1933 185
R811 VDD.n1932 VDD.n1931 185
R812 VDD.n1930 VDD.n1929 185
R813 VDD.n1928 VDD.n1927 185
R814 VDD.n1926 VDD.n1925 185
R815 VDD.n1924 VDD.n1923 185
R816 VDD.n1922 VDD.n1921 185
R817 VDD.n1920 VDD.n1919 185
R818 VDD.n1918 VDD.n1917 185
R819 VDD.n1916 VDD.n1915 185
R820 VDD.n1914 VDD.n1913 185
R821 VDD.n1912 VDD.n1911 185
R822 VDD.n1910 VDD.n1909 185
R823 VDD.n1907 VDD.n1906 185
R824 VDD.n1905 VDD.n1904 185
R825 VDD.n1903 VDD.n1902 185
R826 VDD.n2078 VDD.n2077 185
R827 VDD.n2079 VDD.n387 185
R828 VDD.n2081 VDD.n2080 185
R829 VDD.n2083 VDD.n385 185
R830 VDD.n2085 VDD.n2084 185
R831 VDD.n2086 VDD.n384 185
R832 VDD.n2088 VDD.n2087 185
R833 VDD.n2090 VDD.n382 185
R834 VDD.n2092 VDD.n2091 185
R835 VDD.n2093 VDD.n381 185
R836 VDD.n2095 VDD.n2094 185
R837 VDD.n2097 VDD.n311 185
R838 VDD.n2099 VDD.n2098 185
R839 VDD.n2101 VDD.n379 185
R840 VDD.n2103 VDD.n2102 185
R841 VDD.n2104 VDD.n378 185
R842 VDD.n2106 VDD.n2105 185
R843 VDD.n2108 VDD.n376 185
R844 VDD.n2110 VDD.n2109 185
R845 VDD.n2111 VDD.n375 185
R846 VDD.n2113 VDD.n2112 185
R847 VDD.n2115 VDD.n374 185
R848 VDD.n2117 VDD.n2116 185
R849 VDD.n2116 VDD.n354 185
R850 VDD.n2076 VDD.n2074 185
R851 VDD.n2076 VDD.n369 185
R852 VDD.n2073 VDD.n368 185
R853 VDD.n2121 VDD.n368 185
R854 VDD.n2072 VDD.n2071 185
R855 VDD.n2071 VDD.n367 185
R856 VDD.n2070 VDD.n391 185
R857 VDD.n2070 VDD.n2069 185
R858 VDD.n1764 VDD.n392 185
R859 VDD.n1854 VDD.n392 185
R860 VDD.n1765 VDD.n399 185
R861 VDD.n2063 VDD.n399 185
R862 VDD.n1767 VDD.n1766 185
R863 VDD.n1766 VDD.n398 185
R864 VDD.n1768 VDD.n406 185
R865 VDD.n2023 VDD.n406 185
R866 VDD.n1770 VDD.n1769 185
R867 VDD.n1769 VDD.n405 185
R868 VDD.n1771 VDD.n412 185
R869 VDD.n2017 VDD.n412 185
R870 VDD.n1773 VDD.n1772 185
R871 VDD.n1772 VDD.n411 185
R872 VDD.n1774 VDD.n418 185
R873 VDD.n2011 VDD.n418 185
R874 VDD.n1776 VDD.n1775 185
R875 VDD.n1775 VDD.n417 185
R876 VDD.n1777 VDD.n424 185
R877 VDD.n2005 VDD.n424 185
R878 VDD.n1779 VDD.n1778 185
R879 VDD.n1778 VDD.n423 185
R880 VDD.n1780 VDD.n430 185
R881 VDD.n1999 VDD.n430 185
R882 VDD.n1782 VDD.n1781 185
R883 VDD.n1781 VDD.n429 185
R884 VDD.n1783 VDD.n435 185
R885 VDD.n1993 VDD.n435 185
R886 VDD.n1785 VDD.n1784 185
R887 VDD.n1784 VDD.n443 185
R888 VDD.n1786 VDD.n441 185
R889 VDD.n1987 VDD.n441 185
R890 VDD.n1788 VDD.n1787 185
R891 VDD.n1787 VDD.n440 185
R892 VDD.n1789 VDD.n447 185
R893 VDD.n1981 VDD.n447 185
R894 VDD.n1886 VDD.n1885 185
R895 VDD.n1885 VDD.n1884 185
R896 VDD.n1887 VDD.n453 185
R897 VDD.n1975 VDD.n453 185
R898 VDD.n1889 VDD.n1888 185
R899 VDD.n1888 VDD.n452 185
R900 VDD.n1890 VDD.n459 185
R901 VDD.n1969 VDD.n459 185
R902 VDD.n1892 VDD.n1891 185
R903 VDD.n1891 VDD.n458 185
R904 VDD.n1893 VDD.n465 185
R905 VDD.n1963 VDD.n465 185
R906 VDD.n1895 VDD.n1894 185
R907 VDD.n1894 VDD.n464 185
R908 VDD.n1896 VDD.n471 185
R909 VDD.n1957 VDD.n471 185
R910 VDD.n1898 VDD.n1897 185
R911 VDD.n1897 VDD.n470 185
R912 VDD.n1899 VDD.n477 185
R913 VDD.n1951 VDD.n477 185
R914 VDD.n1901 VDD.n1900 185
R915 VDD.n1901 VDD.n476 185
R916 VDD.n1485 VDD.n1484 185
R917 VDD.n1486 VDD.n1485 185
R918 VDD.n649 VDD.n647 185
R919 VDD.n647 VDD.n641 185
R920 VDD.n1141 VDD.n1140 185
R921 VDD.n1140 VDD.n1139 185
R922 VDD.n652 VDD.n651 185
R923 VDD.n653 VDD.n652 185
R924 VDD.n1130 VDD.n1129 185
R925 VDD.n1131 VDD.n1130 185
R926 VDD.n661 VDD.n660 185
R927 VDD.n660 VDD.n659 185
R928 VDD.n1125 VDD.n1124 185
R929 VDD.n1124 VDD.n1123 185
R930 VDD.n664 VDD.n663 185
R931 VDD.n671 VDD.n664 185
R932 VDD.n1114 VDD.n1113 185
R933 VDD.n1115 VDD.n1114 185
R934 VDD.n673 VDD.n672 185
R935 VDD.n672 VDD.n670 185
R936 VDD.n1109 VDD.n1108 185
R937 VDD.n1108 VDD.n1107 185
R938 VDD.n676 VDD.n675 185
R939 VDD.n677 VDD.n676 185
R940 VDD.n1098 VDD.n1097 185
R941 VDD.n1099 VDD.n1098 185
R942 VDD.n685 VDD.n684 185
R943 VDD.n684 VDD.n683 185
R944 VDD.n1093 VDD.n1092 185
R945 VDD.n1092 VDD.n1091 185
R946 VDD.n688 VDD.n687 185
R947 VDD.n695 VDD.n688 185
R948 VDD.n1082 VDD.n1081 185
R949 VDD.n1083 VDD.n1082 185
R950 VDD.n697 VDD.n696 185
R951 VDD.n696 VDD.n694 185
R952 VDD.n1077 VDD.n1076 185
R953 VDD.n1076 VDD.n1075 185
R954 VDD.n730 VDD.n729 185
R955 VDD.n731 VDD.n730 185
R956 VDD.n1066 VDD.n1065 185
R957 VDD.n1067 VDD.n1066 185
R958 VDD.n739 VDD.n738 185
R959 VDD.n738 VDD.n737 185
R960 VDD.n1060 VDD.n1059 185
R961 VDD.n1059 VDD.n1058 185
R962 VDD.n742 VDD.n741 185
R963 VDD.n749 VDD.n742 185
R964 VDD.n1049 VDD.n1048 185
R965 VDD.n1050 VDD.n1049 185
R966 VDD.n751 VDD.n750 185
R967 VDD.n750 VDD.n748 185
R968 VDD.n1044 VDD.n1043 185
R969 VDD.n1043 VDD.n1042 185
R970 VDD.n754 VDD.n753 185
R971 VDD.n755 VDD.n754 185
R972 VDD.n1033 VDD.n1032 185
R973 VDD.n1034 VDD.n1033 185
R974 VDD.n763 VDD.n762 185
R975 VDD.n762 VDD.n761 185
R976 VDD.n1028 VDD.n1027 185
R977 VDD.n1027 VDD.n1026 185
R978 VDD.n766 VDD.n765 185
R979 VDD.n773 VDD.n766 185
R980 VDD.n1017 VDD.n1016 185
R981 VDD.n1018 VDD.n1017 185
R982 VDD.n775 VDD.n774 185
R983 VDD.n774 VDD.n772 185
R984 VDD.n1012 VDD.n1011 185
R985 VDD.n1011 VDD.n1010 185
R986 VDD.n778 VDD.n777 185
R987 VDD.n779 VDD.n778 185
R988 VDD.n1001 VDD.n1000 185
R989 VDD.n1002 VDD.n1001 185
R990 VDD.n787 VDD.n786 185
R991 VDD.n786 VDD.n785 185
R992 VDD.n996 VDD.n995 185
R993 VDD.n790 VDD.n789 185
R994 VDD.n992 VDD.n991 185
R995 VDD.n993 VDD.n992 185
R996 VDD.n820 VDD.n819 185
R997 VDD.n987 VDD.n822 185
R998 VDD.n986 VDD.n823 185
R999 VDD.n985 VDD.n824 185
R1000 VDD.n826 VDD.n825 185
R1001 VDD.n981 VDD.n828 185
R1002 VDD.n980 VDD.n829 185
R1003 VDD.n979 VDD.n830 185
R1004 VDD.n832 VDD.n831 185
R1005 VDD.n975 VDD.n834 185
R1006 VDD.n974 VDD.n835 185
R1007 VDD.n973 VDD.n836 185
R1008 VDD.n838 VDD.n837 185
R1009 VDD.n969 VDD.n840 185
R1010 VDD.n968 VDD.n965 185
R1011 VDD.n964 VDD.n841 185
R1012 VDD.n843 VDD.n842 185
R1013 VDD.n960 VDD.n845 185
R1014 VDD.n959 VDD.n846 185
R1015 VDD.n958 VDD.n847 185
R1016 VDD.n849 VDD.n848 185
R1017 VDD.n954 VDD.n851 185
R1018 VDD.n953 VDD.n852 185
R1019 VDD.n952 VDD.n853 185
R1020 VDD.n855 VDD.n854 185
R1021 VDD.n948 VDD.n857 185
R1022 VDD.n947 VDD.n858 185
R1023 VDD.n946 VDD.n859 185
R1024 VDD.n861 VDD.n860 185
R1025 VDD.n942 VDD.n863 185
R1026 VDD.n941 VDD.n864 185
R1027 VDD.n940 VDD.n865 185
R1028 VDD.n867 VDD.n866 185
R1029 VDD.n936 VDD.n869 185
R1030 VDD.n935 VDD.n932 185
R1031 VDD.n931 VDD.n870 185
R1032 VDD.n872 VDD.n871 185
R1033 VDD.n927 VDD.n874 185
R1034 VDD.n926 VDD.n875 185
R1035 VDD.n925 VDD.n876 185
R1036 VDD.n878 VDD.n877 185
R1037 VDD.n921 VDD.n880 185
R1038 VDD.n920 VDD.n881 185
R1039 VDD.n919 VDD.n882 185
R1040 VDD.n884 VDD.n883 185
R1041 VDD.n915 VDD.n886 185
R1042 VDD.n914 VDD.n887 185
R1043 VDD.n913 VDD.n888 185
R1044 VDD.n890 VDD.n889 185
R1045 VDD.n909 VDD.n892 185
R1046 VDD.n908 VDD.n893 185
R1047 VDD.n907 VDD.n894 185
R1048 VDD.n896 VDD.n895 185
R1049 VDD.n903 VDD.n898 185
R1050 VDD.n899 VDD.n818 185
R1051 VDD.n993 VDD.n818 185
R1052 VDD.n1491 VDD.n637 185
R1053 VDD.n1495 VDD.n636 185
R1054 VDD.n1496 VDD.n635 185
R1055 VDD.n643 VDD.n633 185
R1056 VDD.n1500 VDD.n632 185
R1057 VDD.n1501 VDD.n631 185
R1058 VDD.n1502 VDD.n630 185
R1059 VDD.n1225 VDD.n629 185
R1060 VDD.n1227 VDD.n1226 185
R1061 VDD.n1229 VDD.n1223 185
R1062 VDD.n1231 VDD.n1230 185
R1063 VDD.n1232 VDD.n1219 185
R1064 VDD.n1234 VDD.n1233 185
R1065 VDD.n1236 VDD.n1217 185
R1066 VDD.n1238 VDD.n1237 185
R1067 VDD.n1239 VDD.n1213 185
R1068 VDD.n1241 VDD.n1240 185
R1069 VDD.n1243 VDD.n1211 185
R1070 VDD.n1245 VDD.n1244 185
R1071 VDD.n1206 VDD.n1205 185
R1072 VDD.n1250 VDD.n1249 185
R1073 VDD.n1252 VDD.n1203 185
R1074 VDD.n1254 VDD.n1253 185
R1075 VDD.n1255 VDD.n1198 185
R1076 VDD.n1257 VDD.n1256 185
R1077 VDD.n1259 VDD.n1196 185
R1078 VDD.n1261 VDD.n1260 185
R1079 VDD.n1262 VDD.n1191 185
R1080 VDD.n1264 VDD.n1263 185
R1081 VDD.n1266 VDD.n1189 185
R1082 VDD.n1268 VDD.n1267 185
R1083 VDD.n1269 VDD.n1184 185
R1084 VDD.n1271 VDD.n1270 185
R1085 VDD.n1273 VDD.n1182 185
R1086 VDD.n1275 VDD.n1274 185
R1087 VDD.n1276 VDD.n1178 185
R1088 VDD.n1278 VDD.n1277 185
R1089 VDD.n1280 VDD.n1176 185
R1090 VDD.n1282 VDD.n1281 185
R1091 VDD.n1171 VDD.n1170 185
R1092 VDD.n1287 VDD.n1286 185
R1093 VDD.n1289 VDD.n1168 185
R1094 VDD.n1291 VDD.n1290 185
R1095 VDD.n1292 VDD.n1163 185
R1096 VDD.n1294 VDD.n1293 185
R1097 VDD.n1296 VDD.n1162 185
R1098 VDD.n1297 VDD.n1159 185
R1099 VDD.n1300 VDD.n1299 185
R1100 VDD.n1161 VDD.n1158 185
R1101 VDD.n1155 VDD.n1154 185
R1102 VDD.n1469 VDD.n1468 185
R1103 VDD.n1471 VDD.n1152 185
R1104 VDD.n1473 VDD.n1472 185
R1105 VDD.n1474 VDD.n1147 185
R1106 VDD.n1476 VDD.n1475 185
R1107 VDD.n1478 VDD.n1145 185
R1108 VDD.n1480 VDD.n1479 185
R1109 VDD.n1481 VDD.n648 185
R1110 VDD.n1488 VDD.n1487 185
R1111 VDD.n1487 VDD.n1486 185
R1112 VDD.n640 VDD.n639 185
R1113 VDD.n641 VDD.n640 185
R1114 VDD.n1138 VDD.n1137 185
R1115 VDD.n1139 VDD.n1138 185
R1116 VDD.n655 VDD.n654 185
R1117 VDD.n654 VDD.n653 185
R1118 VDD.n1133 VDD.n1132 185
R1119 VDD.n1132 VDD.n1131 185
R1120 VDD.n658 VDD.n657 185
R1121 VDD.n659 VDD.n658 185
R1122 VDD.n1122 VDD.n1121 185
R1123 VDD.n1123 VDD.n1122 185
R1124 VDD.n666 VDD.n665 185
R1125 VDD.n671 VDD.n665 185
R1126 VDD.n1117 VDD.n1116 185
R1127 VDD.n1116 VDD.n1115 185
R1128 VDD.n669 VDD.n668 185
R1129 VDD.n670 VDD.n669 185
R1130 VDD.n1106 VDD.n1105 185
R1131 VDD.n1107 VDD.n1106 185
R1132 VDD.n679 VDD.n678 185
R1133 VDD.n678 VDD.n677 185
R1134 VDD.n1101 VDD.n1100 185
R1135 VDD.n1100 VDD.n1099 185
R1136 VDD.n682 VDD.n681 185
R1137 VDD.n683 VDD.n682 185
R1138 VDD.n1090 VDD.n1089 185
R1139 VDD.n1091 VDD.n1090 185
R1140 VDD.n690 VDD.n689 185
R1141 VDD.n695 VDD.n689 185
R1142 VDD.n1085 VDD.n1084 185
R1143 VDD.n1084 VDD.n1083 185
R1144 VDD.n693 VDD.n692 185
R1145 VDD.n694 VDD.n693 185
R1146 VDD.n1074 VDD.n1073 185
R1147 VDD.n1075 VDD.n1074 185
R1148 VDD.n733 VDD.n732 185
R1149 VDD.n732 VDD.n731 185
R1150 VDD.n1069 VDD.n1068 185
R1151 VDD.n1068 VDD.n1067 185
R1152 VDD.n736 VDD.n735 185
R1153 VDD.n737 VDD.n736 185
R1154 VDD.n1057 VDD.n1056 185
R1155 VDD.n1058 VDD.n1057 185
R1156 VDD.n744 VDD.n743 185
R1157 VDD.n749 VDD.n743 185
R1158 VDD.n1052 VDD.n1051 185
R1159 VDD.n1051 VDD.n1050 185
R1160 VDD.n747 VDD.n746 185
R1161 VDD.n748 VDD.n747 185
R1162 VDD.n1041 VDD.n1040 185
R1163 VDD.n1042 VDD.n1041 185
R1164 VDD.n757 VDD.n756 185
R1165 VDD.n756 VDD.n755 185
R1166 VDD.n1036 VDD.n1035 185
R1167 VDD.n1035 VDD.n1034 185
R1168 VDD.n760 VDD.n759 185
R1169 VDD.n761 VDD.n760 185
R1170 VDD.n1025 VDD.n1024 185
R1171 VDD.n1026 VDD.n1025 185
R1172 VDD.n768 VDD.n767 185
R1173 VDD.n773 VDD.n767 185
R1174 VDD.n1020 VDD.n1019 185
R1175 VDD.n1019 VDD.n1018 185
R1176 VDD.n771 VDD.n770 185
R1177 VDD.n772 VDD.n771 185
R1178 VDD.n1009 VDD.n1008 185
R1179 VDD.n1010 VDD.n1009 185
R1180 VDD.n781 VDD.n780 185
R1181 VDD.n780 VDD.n779 185
R1182 VDD.n1004 VDD.n1003 185
R1183 VDD.n1003 VDD.n1002 185
R1184 VDD.n784 VDD.n783 185
R1185 VDD.n785 VDD.n784 185
R1186 VDD.n2276 VDD.n2275 185
R1187 VDD.n274 VDD.n273 185
R1188 VDD.n2272 VDD.n2271 185
R1189 VDD.n2273 VDD.n2272 185
R1190 VDD.n2270 VDD.n303 185
R1191 VDD.n2269 VDD.n2268 185
R1192 VDD.n2267 VDD.n2266 185
R1193 VDD.n2265 VDD.n2264 185
R1194 VDD.n2263 VDD.n2262 185
R1195 VDD.n312 VDD.n309 185
R1196 VDD.n314 VDD.n313 185
R1197 VDD.n2258 VDD.n315 185
R1198 VDD.n2257 VDD.n2256 185
R1199 VDD.n2255 VDD.n2254 185
R1200 VDD.n2253 VDD.n2252 185
R1201 VDD.n2251 VDD.n2250 185
R1202 VDD.n2249 VDD.n2248 185
R1203 VDD.n2247 VDD.n2246 185
R1204 VDD.n2245 VDD.n2244 185
R1205 VDD.n2236 VDD.n321 185
R1206 VDD.n2238 VDD.n2237 185
R1207 VDD.n2235 VDD.n2234 185
R1208 VDD.n2233 VDD.n2232 185
R1209 VDD.n2231 VDD.n2230 185
R1210 VDD.n2229 VDD.n2228 185
R1211 VDD.n2227 VDD.n2226 185
R1212 VDD.n2225 VDD.n2224 185
R1213 VDD.n2223 VDD.n2222 185
R1214 VDD.n2221 VDD.n2220 185
R1215 VDD.n2219 VDD.n2218 185
R1216 VDD.n2217 VDD.n2216 185
R1217 VDD.n2215 VDD.n2214 185
R1218 VDD.n2213 VDD.n2212 185
R1219 VDD.n2211 VDD.n2210 185
R1220 VDD.n2209 VDD.n2208 185
R1221 VDD.n2207 VDD.n2206 185
R1222 VDD.n2205 VDD.n2204 185
R1223 VDD.n2203 VDD.n2202 185
R1224 VDD.n2201 VDD.n2200 185
R1225 VDD.n2194 VDD.n339 185
R1226 VDD.n2196 VDD.n2195 185
R1227 VDD.n2193 VDD.n2192 185
R1228 VDD.n2191 VDD.n2190 185
R1229 VDD.n2189 VDD.n2188 185
R1230 VDD.n2187 VDD.n2186 185
R1231 VDD.n2185 VDD.n2184 185
R1232 VDD.n2183 VDD.n2182 185
R1233 VDD.n2181 VDD.n2180 185
R1234 VDD.n2179 VDD.n2178 185
R1235 VDD.n2148 VDD.n349 185
R1236 VDD.n2150 VDD.n2149 185
R1237 VDD.n2174 VDD.n2151 185
R1238 VDD.n2173 VDD.n2172 185
R1239 VDD.n2171 VDD.n2170 185
R1240 VDD.n2169 VDD.n2168 185
R1241 VDD.n2167 VDD.n2166 185
R1242 VDD.n2165 VDD.n2164 185
R1243 VDD.n2163 VDD.n2162 185
R1244 VDD.n2158 VDD.n302 185
R1245 VDD.n2273 VDD.n302 185
R1246 VDD.n2382 VDD.n2381 185
R1247 VDD.n2384 VDD.n197 185
R1248 VDD.n2386 VDD.n2385 185
R1249 VDD.n2387 VDD.n192 185
R1250 VDD.n2389 VDD.n2388 185
R1251 VDD.n2391 VDD.n190 185
R1252 VDD.n2393 VDD.n2392 185
R1253 VDD.n2394 VDD.n185 185
R1254 VDD.n2396 VDD.n2395 185
R1255 VDD.n2398 VDD.n183 185
R1256 VDD.n2400 VDD.n2399 185
R1257 VDD.n2401 VDD.n178 185
R1258 VDD.n2403 VDD.n2402 185
R1259 VDD.n2405 VDD.n176 185
R1260 VDD.n2407 VDD.n2406 185
R1261 VDD.n2408 VDD.n172 185
R1262 VDD.n2410 VDD.n2409 185
R1263 VDD.n2412 VDD.n170 185
R1264 VDD.n2414 VDD.n2413 185
R1265 VDD.n165 VDD.n164 185
R1266 VDD.n2419 VDD.n2418 185
R1267 VDD.n2421 VDD.n162 185
R1268 VDD.n2423 VDD.n2422 185
R1269 VDD.n2424 VDD.n157 185
R1270 VDD.n2426 VDD.n2425 185
R1271 VDD.n2428 VDD.n155 185
R1272 VDD.n2430 VDD.n2429 185
R1273 VDD.n2431 VDD.n150 185
R1274 VDD.n2433 VDD.n2432 185
R1275 VDD.n2435 VDD.n148 185
R1276 VDD.n2437 VDD.n2436 185
R1277 VDD.n2438 VDD.n143 185
R1278 VDD.n2440 VDD.n2439 185
R1279 VDD.n2442 VDD.n141 185
R1280 VDD.n2444 VDD.n2443 185
R1281 VDD.n2445 VDD.n137 185
R1282 VDD.n2447 VDD.n2446 185
R1283 VDD.n2449 VDD.n135 185
R1284 VDD.n2451 VDD.n2450 185
R1285 VDD.n130 VDD.n129 185
R1286 VDD.n2456 VDD.n2455 185
R1287 VDD.n2458 VDD.n127 185
R1288 VDD.n2460 VDD.n2459 185
R1289 VDD.n2461 VDD.n122 185
R1290 VDD.n2463 VDD.n2462 185
R1291 VDD.n2465 VDD.n120 185
R1292 VDD.n2467 VDD.n2466 185
R1293 VDD.n2468 VDD.n115 185
R1294 VDD.n2470 VDD.n2469 185
R1295 VDD.n2472 VDD.n113 185
R1296 VDD.n2474 VDD.n2473 185
R1297 VDD.n2475 VDD.n107 185
R1298 VDD.n2477 VDD.n2476 185
R1299 VDD.n2479 VDD.n106 185
R1300 VDD.n2480 VDD.n105 185
R1301 VDD.n2483 VDD.n2482 185
R1302 VDD.n2484 VDD.n103 185
R1303 VDD.n2485 VDD.n99 185
R1304 VDD.n2378 VDD.n97 185
R1305 VDD.n2490 VDD.n97 185
R1306 VDD.n2377 VDD.n96 185
R1307 VDD.n2491 VDD.n96 185
R1308 VDD.n2376 VDD.n95 185
R1309 VDD.n2492 VDD.n95 185
R1310 VDD.n205 VDD.n204 185
R1311 VDD.n204 VDD.n87 185
R1312 VDD.n2372 VDD.n86 185
R1313 VDD.n2498 VDD.n86 185
R1314 VDD.n2371 VDD.n85 185
R1315 VDD.n2499 VDD.n85 185
R1316 VDD.n2370 VDD.n84 185
R1317 VDD.n2500 VDD.n84 185
R1318 VDD.n208 VDD.n207 185
R1319 VDD.n207 VDD.n76 185
R1320 VDD.n2366 VDD.n75 185
R1321 VDD.n2506 VDD.n75 185
R1322 VDD.n2365 VDD.n74 185
R1323 VDD.n2507 VDD.n74 185
R1324 VDD.n2364 VDD.n73 185
R1325 VDD.n2508 VDD.n73 185
R1326 VDD.n211 VDD.n210 185
R1327 VDD.n210 VDD.n72 185
R1328 VDD.n2360 VDD.n64 185
R1329 VDD.n2514 VDD.n64 185
R1330 VDD.n2359 VDD.n63 185
R1331 VDD.n2515 VDD.n63 185
R1332 VDD.n2358 VDD.n62 185
R1333 VDD.n2516 VDD.n62 185
R1334 VDD.n214 VDD.n213 185
R1335 VDD.n213 VDD.n55 185
R1336 VDD.n2354 VDD.n54 185
R1337 VDD.n2522 VDD.n54 185
R1338 VDD.n2353 VDD.n53 185
R1339 VDD.n2523 VDD.n53 185
R1340 VDD.n2352 VDD.n52 185
R1341 VDD.n2524 VDD.n52 185
R1342 VDD.n220 VDD.n216 185
R1343 VDD.n220 VDD.n51 185
R1344 VDD.n2348 VDD.n2347 185
R1345 VDD.n2347 VDD.n2346 185
R1346 VDD.n219 VDD.n218 185
R1347 VDD.n221 VDD.n219 185
R1348 VDD.n2337 VDD.n2336 185
R1349 VDD.n2338 VDD.n2337 185
R1350 VDD.n228 VDD.n227 185
R1351 VDD.n233 VDD.n227 185
R1352 VDD.n2332 VDD.n2331 185
R1353 VDD.n2331 VDD.n2330 185
R1354 VDD.n231 VDD.n230 185
R1355 VDD.n232 VDD.n231 185
R1356 VDD.n2321 VDD.n2320 185
R1357 VDD.n2322 VDD.n2321 185
R1358 VDD.n241 VDD.n240 185
R1359 VDD.n240 VDD.n239 185
R1360 VDD.n2316 VDD.n2315 185
R1361 VDD.n2315 VDD.n2314 185
R1362 VDD.n244 VDD.n243 185
R1363 VDD.n245 VDD.n244 185
R1364 VDD.n2305 VDD.n2304 185
R1365 VDD.n2306 VDD.n2305 185
R1366 VDD.n252 VDD.n251 185
R1367 VDD.n257 VDD.n251 185
R1368 VDD.n2300 VDD.n2299 185
R1369 VDD.n2299 VDD.n2298 185
R1370 VDD.n255 VDD.n254 185
R1371 VDD.n256 VDD.n255 185
R1372 VDD.n2289 VDD.n2288 185
R1373 VDD.n2290 VDD.n2289 185
R1374 VDD.n265 VDD.n264 185
R1375 VDD.n264 VDD.n263 185
R1376 VDD.n2284 VDD.n2283 185
R1377 VDD.n2283 VDD.n2282 185
R1378 VDD.n268 VDD.n267 185
R1379 VDD.n269 VDD.n268 185
R1380 VDD.n271 VDD.n270 185
R1381 VDD.n270 VDD.n269 185
R1382 VDD.n2281 VDD.n2280 185
R1383 VDD.n2282 VDD.n2281 185
R1384 VDD.n262 VDD.n261 185
R1385 VDD.n263 VDD.n262 185
R1386 VDD.n2292 VDD.n2291 185
R1387 VDD.n2291 VDD.n2290 185
R1388 VDD.n259 VDD.n258 185
R1389 VDD.n258 VDD.n256 185
R1390 VDD.n2297 VDD.n2296 185
R1391 VDD.n2298 VDD.n2297 185
R1392 VDD.n250 VDD.n249 185
R1393 VDD.n257 VDD.n250 185
R1394 VDD.n2308 VDD.n2307 185
R1395 VDD.n2307 VDD.n2306 185
R1396 VDD.n247 VDD.n246 185
R1397 VDD.n246 VDD.n245 185
R1398 VDD.n2313 VDD.n2312 185
R1399 VDD.n2314 VDD.n2313 185
R1400 VDD.n238 VDD.n237 185
R1401 VDD.n239 VDD.n238 185
R1402 VDD.n2324 VDD.n2323 185
R1403 VDD.n2323 VDD.n2322 185
R1404 VDD.n235 VDD.n234 185
R1405 VDD.n234 VDD.n232 185
R1406 VDD.n2329 VDD.n2328 185
R1407 VDD.n2330 VDD.n2329 185
R1408 VDD.n226 VDD.n225 185
R1409 VDD.n233 VDD.n226 185
R1410 VDD.n2340 VDD.n2339 185
R1411 VDD.n2339 VDD.n2338 185
R1412 VDD.n223 VDD.n222 185
R1413 VDD.n222 VDD.n221 185
R1414 VDD.n2345 VDD.n2344 185
R1415 VDD.n2346 VDD.n2345 185
R1416 VDD.n49 VDD.n47 185
R1417 VDD.n51 VDD.n49 185
R1418 VDD.n2526 VDD.n2525 185
R1419 VDD.n2525 VDD.n2524 185
R1420 VDD.n50 VDD.n48 185
R1421 VDD.n2523 VDD.n50 185
R1422 VDD.n2521 VDD.n2520 185
R1423 VDD.n2522 VDD.n2521 185
R1424 VDD.n2519 VDD.n56 185
R1425 VDD.n56 VDD.n55 185
R1426 VDD.n2518 VDD.n2517 185
R1427 VDD.n2517 VDD.n2516 185
R1428 VDD.n61 VDD.n60 185
R1429 VDD.n2515 VDD.n61 185
R1430 VDD.n2513 VDD.n2512 185
R1431 VDD.n2514 VDD.n2513 185
R1432 VDD.n2511 VDD.n65 185
R1433 VDD.n72 VDD.n65 185
R1434 VDD.n2510 VDD.n2509 185
R1435 VDD.n2509 VDD.n2508 185
R1436 VDD.n71 VDD.n70 185
R1437 VDD.n2507 VDD.n71 185
R1438 VDD.n2505 VDD.n2504 185
R1439 VDD.n2506 VDD.n2505 185
R1440 VDD.n2503 VDD.n77 185
R1441 VDD.n77 VDD.n76 185
R1442 VDD.n2502 VDD.n2501 185
R1443 VDD.n2501 VDD.n2500 185
R1444 VDD.n83 VDD.n82 185
R1445 VDD.n2499 VDD.n83 185
R1446 VDD.n2497 VDD.n2496 185
R1447 VDD.n2498 VDD.n2497 185
R1448 VDD.n2495 VDD.n88 185
R1449 VDD.n88 VDD.n87 185
R1450 VDD.n2494 VDD.n2493 185
R1451 VDD.n2493 VDD.n2492 185
R1452 VDD.n94 VDD.n93 185
R1453 VDD.n2491 VDD.n94 185
R1454 VDD.n2489 VDD.n2488 185
R1455 VDD.n2490 VDD.n2489 185
R1456 VDD.n1678 VDD.n1677 185
R1457 VDD.n1677 VDD.n482 185
R1458 VDD.n1679 VDD.n515 185
R1459 VDD.n1689 VDD.n515 185
R1460 VDD.n1680 VDD.n523 185
R1461 VDD.n523 VDD.n521 185
R1462 VDD.n1682 VDD.n1681 185
R1463 VDD.n1683 VDD.n1682 185
R1464 VDD.n524 VDD.n522 185
R1465 VDD.n1623 VDD.n522 185
R1466 VDD.n1603 VDD.n1602 185
R1467 VDD.n1602 VDD.n530 185
R1468 VDD.n1604 VDD.n536 185
R1469 VDD.n1615 VDD.n536 185
R1470 VDD.n1605 VDD.n545 185
R1471 VDD.n545 VDD.n534 185
R1472 VDD.n1607 VDD.n1606 185
R1473 VDD.n1608 VDD.n1607 185
R1474 VDD.n1601 VDD.n544 185
R1475 VDD.n544 VDD.n541 185
R1476 VDD.n1600 VDD.n1599 185
R1477 VDD.n1599 VDD.n1598 185
R1478 VDD.n547 VDD.n546 185
R1479 VDD.n556 VDD.n547 185
R1480 VDD.n1591 VDD.n1590 185
R1481 VDD.n1592 VDD.n1591 185
R1482 VDD.n1589 VDD.n557 185
R1483 VDD.n557 VDD.n553 185
R1484 VDD.n1588 VDD.n1587 185
R1485 VDD.n1587 VDD.n1586 185
R1486 VDD.n559 VDD.n558 185
R1487 VDD.n1414 VDD.n559 185
R1488 VDD.n1579 VDD.n1578 185
R1489 VDD.n1580 VDD.n1579 185
R1490 VDD.n1577 VDD.n568 185
R1491 VDD.n568 VDD.n565 185
R1492 VDD.n1576 VDD.n1575 185
R1493 VDD.n1575 VDD.n1574 185
R1494 VDD.n570 VDD.n569 185
R1495 VDD.n571 VDD.n570 185
R1496 VDD.n1567 VDD.n1566 185
R1497 VDD.n1568 VDD.n1567 185
R1498 VDD.n1565 VDD.n580 185
R1499 VDD.n580 VDD.n577 185
R1500 VDD.n1564 VDD.n1563 185
R1501 VDD.n1563 VDD.n1562 185
R1502 VDD.n582 VDD.n581 185
R1503 VDD.n583 VDD.n582 185
R1504 VDD.n1555 VDD.n1554 185
R1505 VDD.n1556 VDD.n1555 185
R1506 VDD.n1553 VDD.n592 185
R1507 VDD.n592 VDD.n589 185
R1508 VDD.n1552 VDD.n1551 185
R1509 VDD.n1551 VDD.n1550 185
R1510 VDD.n594 VDD.n593 185
R1511 VDD.n595 VDD.n594 185
R1512 VDD.n1543 VDD.n1542 185
R1513 VDD.n1544 VDD.n1543 185
R1514 VDD.n1541 VDD.n603 185
R1515 VDD.n609 VDD.n603 185
R1516 VDD.n1540 VDD.n1539 185
R1517 VDD.n1539 VDD.n1538 185
R1518 VDD.n605 VDD.n604 185
R1519 VDD.n606 VDD.n605 185
R1520 VDD.n1531 VDD.n1530 185
R1521 VDD.n1532 VDD.n1531 185
R1522 VDD.n1632 VDD.n494 185
R1523 VDD.n1738 VDD.n494 185
R1524 VDD.n1634 VDD.n1633 185
R1525 VDD.n1636 VDD.n1635 185
R1526 VDD.n1638 VDD.n1637 185
R1527 VDD.n1640 VDD.n1639 185
R1528 VDD.n1642 VDD.n1641 185
R1529 VDD.n1644 VDD.n1643 185
R1530 VDD.n1646 VDD.n1645 185
R1531 VDD.n1648 VDD.n1647 185
R1532 VDD.n1650 VDD.n1649 185
R1533 VDD.n1652 VDD.n1651 185
R1534 VDD.n1654 VDD.n1653 185
R1535 VDD.n1656 VDD.n1655 185
R1536 VDD.n1658 VDD.n1657 185
R1537 VDD.n1660 VDD.n1659 185
R1538 VDD.n1662 VDD.n1661 185
R1539 VDD.n1664 VDD.n1663 185
R1540 VDD.n1666 VDD.n1665 185
R1541 VDD.n1668 VDD.n1667 185
R1542 VDD.n1670 VDD.n1669 185
R1543 VDD.n1672 VDD.n1671 185
R1544 VDD.n1674 VDD.n1673 185
R1545 VDD.n1676 VDD.n1675 185
R1546 VDD.n1631 VDD.n1630 185
R1547 VDD.n1630 VDD.n482 185
R1548 VDD.n1629 VDD.n514 185
R1549 VDD.n1689 VDD.n514 185
R1550 VDD.n1628 VDD.n1627 185
R1551 VDD.n1627 VDD.n521 185
R1552 VDD.n1626 VDD.n520 185
R1553 VDD.n1683 VDD.n520 185
R1554 VDD.n1625 VDD.n1624 185
R1555 VDD.n1624 VDD.n1623 185
R1556 VDD.n529 VDD.n528 185
R1557 VDD.n530 VDD.n529 185
R1558 VDD.n1399 VDD.n535 185
R1559 VDD.n1615 VDD.n535 185
R1560 VDD.n1401 VDD.n1400 185
R1561 VDD.n1400 VDD.n534 185
R1562 VDD.n1402 VDD.n543 185
R1563 VDD.n1608 VDD.n543 185
R1564 VDD.n1404 VDD.n1403 185
R1565 VDD.n1403 VDD.n541 185
R1566 VDD.n1405 VDD.n549 185
R1567 VDD.n1598 VDD.n549 185
R1568 VDD.n1407 VDD.n1406 185
R1569 VDD.n1406 VDD.n556 185
R1570 VDD.n1408 VDD.n555 185
R1571 VDD.n1592 VDD.n555 185
R1572 VDD.n1410 VDD.n1409 185
R1573 VDD.n1409 VDD.n553 185
R1574 VDD.n1411 VDD.n561 185
R1575 VDD.n1586 VDD.n561 185
R1576 VDD.n1413 VDD.n1412 185
R1577 VDD.n1414 VDD.n1413 185
R1578 VDD.n1398 VDD.n567 185
R1579 VDD.n1580 VDD.n567 185
R1580 VDD.n1397 VDD.n1396 185
R1581 VDD.n1396 VDD.n565 185
R1582 VDD.n1395 VDD.n573 185
R1583 VDD.n1574 VDD.n573 185
R1584 VDD.n1394 VDD.n1393 185
R1585 VDD.n1393 VDD.n571 185
R1586 VDD.n1392 VDD.n579 185
R1587 VDD.n1568 VDD.n579 185
R1588 VDD.n1391 VDD.n1390 185
R1589 VDD.n1390 VDD.n577 185
R1590 VDD.n1389 VDD.n585 185
R1591 VDD.n1562 VDD.n585 185
R1592 VDD.n1388 VDD.n1387 185
R1593 VDD.n1387 VDD.n583 185
R1594 VDD.n1386 VDD.n591 185
R1595 VDD.n1556 VDD.n591 185
R1596 VDD.n1385 VDD.n1384 185
R1597 VDD.n1384 VDD.n589 185
R1598 VDD.n1383 VDD.n597 185
R1599 VDD.n1550 VDD.n597 185
R1600 VDD.n1382 VDD.n1381 185
R1601 VDD.n1381 VDD.n595 185
R1602 VDD.n1380 VDD.n602 185
R1603 VDD.n1544 VDD.n602 185
R1604 VDD.n1379 VDD.n1378 185
R1605 VDD.n1378 VDD.n609 185
R1606 VDD.n1377 VDD.n608 185
R1607 VDD.n1538 VDD.n608 185
R1608 VDD.n1376 VDD.n1375 185
R1609 VDD.n1375 VDD.n606 185
R1610 VDD.n1374 VDD.n615 185
R1611 VDD.n1532 VDD.n615 185
R1612 VDD.n1528 VDD.n616 185
R1613 VDD.n1527 VDD.n1526 185
R1614 VDD.n1524 VDD.n618 185
R1615 VDD.n1522 VDD.n1521 185
R1616 VDD.n1520 VDD.n619 185
R1617 VDD.n1519 VDD.n1518 185
R1618 VDD.n1516 VDD.n620 185
R1619 VDD.n1514 VDD.n1513 185
R1620 VDD.n1512 VDD.n621 185
R1621 VDD.n1511 VDD.n1510 185
R1622 VDD.n1508 VDD.n622 185
R1623 VDD.n1506 VDD.n1505 185
R1624 VDD.n624 VDD.n623 185
R1625 VDD.n1354 VDD.n1352 185
R1626 VDD.n1357 VDD.n1356 185
R1627 VDD.n1358 VDD.n1351 185
R1628 VDD.n1360 VDD.n1359 185
R1629 VDD.n1362 VDD.n1350 185
R1630 VDD.n1365 VDD.n1364 185
R1631 VDD.n1366 VDD.n1347 185
R1632 VDD.n1369 VDD.n1368 185
R1633 VDD.n1371 VDD.n1346 185
R1634 VDD.n1373 VDD.n1372 185
R1635 VDD.n1372 VDD.n613 185
R1636 VDD.n2281 VDD.n270 146.341
R1637 VDD.n2281 VDD.n262 146.341
R1638 VDD.n2291 VDD.n262 146.341
R1639 VDD.n2291 VDD.n258 146.341
R1640 VDD.n2297 VDD.n258 146.341
R1641 VDD.n2297 VDD.n250 146.341
R1642 VDD.n2307 VDD.n250 146.341
R1643 VDD.n2307 VDD.n246 146.341
R1644 VDD.n2313 VDD.n246 146.341
R1645 VDD.n2313 VDD.n238 146.341
R1646 VDD.n2323 VDD.n238 146.341
R1647 VDD.n2323 VDD.n234 146.341
R1648 VDD.n2329 VDD.n234 146.341
R1649 VDD.n2329 VDD.n226 146.341
R1650 VDD.n2339 VDD.n226 146.341
R1651 VDD.n2339 VDD.n222 146.341
R1652 VDD.n2345 VDD.n222 146.341
R1653 VDD.n2345 VDD.n49 146.341
R1654 VDD.n2525 VDD.n49 146.341
R1655 VDD.n2525 VDD.n50 146.341
R1656 VDD.n2521 VDD.n50 146.341
R1657 VDD.n2521 VDD.n56 146.341
R1658 VDD.n2517 VDD.n56 146.341
R1659 VDD.n2517 VDD.n61 146.341
R1660 VDD.n2513 VDD.n61 146.341
R1661 VDD.n2513 VDD.n65 146.341
R1662 VDD.n2509 VDD.n65 146.341
R1663 VDD.n2509 VDD.n71 146.341
R1664 VDD.n2505 VDD.n71 146.341
R1665 VDD.n2505 VDD.n77 146.341
R1666 VDD.n2501 VDD.n77 146.341
R1667 VDD.n2501 VDD.n83 146.341
R1668 VDD.n2497 VDD.n83 146.341
R1669 VDD.n2497 VDD.n88 146.341
R1670 VDD.n2493 VDD.n88 146.341
R1671 VDD.n2493 VDD.n94 146.341
R1672 VDD.n2489 VDD.n94 146.341
R1673 VDD.n2482 VDD.n103 146.341
R1674 VDD.n2480 VDD.n2479 146.341
R1675 VDD.n2477 VDD.n107 146.341
R1676 VDD.n2473 VDD.n2472 146.341
R1677 VDD.n2470 VDD.n115 146.341
R1678 VDD.n2466 VDD.n2465 146.341
R1679 VDD.n2463 VDD.n122 146.341
R1680 VDD.n2459 VDD.n2458 146.341
R1681 VDD.n2456 VDD.n129 146.341
R1682 VDD.n2450 VDD.n2449 146.341
R1683 VDD.n2447 VDD.n137 146.341
R1684 VDD.n2443 VDD.n2442 146.341
R1685 VDD.n2440 VDD.n143 146.341
R1686 VDD.n2436 VDD.n2435 146.341
R1687 VDD.n2433 VDD.n150 146.341
R1688 VDD.n2429 VDD.n2428 146.341
R1689 VDD.n2426 VDD.n157 146.341
R1690 VDD.n2422 VDD.n2421 146.341
R1691 VDD.n2419 VDD.n164 146.341
R1692 VDD.n2413 VDD.n2412 146.341
R1693 VDD.n2410 VDD.n172 146.341
R1694 VDD.n2406 VDD.n2405 146.341
R1695 VDD.n2403 VDD.n178 146.341
R1696 VDD.n2399 VDD.n2398 146.341
R1697 VDD.n2396 VDD.n185 146.341
R1698 VDD.n2392 VDD.n2391 146.341
R1699 VDD.n2389 VDD.n192 146.341
R1700 VDD.n2385 VDD.n2384 146.341
R1701 VDD.n2283 VDD.n268 146.341
R1702 VDD.n2283 VDD.n264 146.341
R1703 VDD.n2289 VDD.n264 146.341
R1704 VDD.n2289 VDD.n255 146.341
R1705 VDD.n2299 VDD.n255 146.341
R1706 VDD.n2299 VDD.n251 146.341
R1707 VDD.n2305 VDD.n251 146.341
R1708 VDD.n2305 VDD.n244 146.341
R1709 VDD.n2315 VDD.n244 146.341
R1710 VDD.n2315 VDD.n240 146.341
R1711 VDD.n2321 VDD.n240 146.341
R1712 VDD.n2321 VDD.n231 146.341
R1713 VDD.n2331 VDD.n231 146.341
R1714 VDD.n2331 VDD.n227 146.341
R1715 VDD.n2337 VDD.n227 146.341
R1716 VDD.n2337 VDD.n219 146.341
R1717 VDD.n2347 VDD.n219 146.341
R1718 VDD.n2347 VDD.n220 146.341
R1719 VDD.n220 VDD.n52 146.341
R1720 VDD.n53 VDD.n52 146.341
R1721 VDD.n54 VDD.n53 146.341
R1722 VDD.n213 VDD.n54 146.341
R1723 VDD.n213 VDD.n62 146.341
R1724 VDD.n63 VDD.n62 146.341
R1725 VDD.n64 VDD.n63 146.341
R1726 VDD.n210 VDD.n64 146.341
R1727 VDD.n210 VDD.n73 146.341
R1728 VDD.n74 VDD.n73 146.341
R1729 VDD.n75 VDD.n74 146.341
R1730 VDD.n207 VDD.n75 146.341
R1731 VDD.n207 VDD.n84 146.341
R1732 VDD.n85 VDD.n84 146.341
R1733 VDD.n86 VDD.n85 146.341
R1734 VDD.n204 VDD.n86 146.341
R1735 VDD.n204 VDD.n95 146.341
R1736 VDD.n96 VDD.n95 146.341
R1737 VDD.n97 VDD.n96 146.341
R1738 VDD.n2272 VDD.n274 146.341
R1739 VDD.n2272 VDD.n303 146.341
R1740 VDD.n2268 VDD.n2267 146.341
R1741 VDD.n2264 VDD.n2263 146.341
R1742 VDD.n313 VDD.n312 146.341
R1743 VDD.n2256 VDD.n315 146.341
R1744 VDD.n2254 VDD.n2253 146.341
R1745 VDD.n2250 VDD.n2249 146.341
R1746 VDD.n2246 VDD.n2245 146.341
R1747 VDD.n2237 VDD.n2236 146.341
R1748 VDD.n2234 VDD.n2233 146.341
R1749 VDD.n2230 VDD.n2229 146.341
R1750 VDD.n2226 VDD.n2225 146.341
R1751 VDD.n2222 VDD.n2221 146.341
R1752 VDD.n2218 VDD.n2217 146.341
R1753 VDD.n2214 VDD.n2213 146.341
R1754 VDD.n2210 VDD.n2209 146.341
R1755 VDD.n2206 VDD.n2205 146.341
R1756 VDD.n2202 VDD.n2201 146.341
R1757 VDD.n2195 VDD.n2194 146.341
R1758 VDD.n2192 VDD.n2191 146.341
R1759 VDD.n2188 VDD.n2187 146.341
R1760 VDD.n2184 VDD.n2183 146.341
R1761 VDD.n2180 VDD.n2179 146.341
R1762 VDD.n2149 VDD.n2148 146.341
R1763 VDD.n2172 VDD.n2151 146.341
R1764 VDD.n2170 VDD.n2169 146.341
R1765 VDD.n2166 VDD.n2165 146.341
R1766 VDD.n2162 VDD.n302 146.341
R1767 VDD.n1479 VDD.n1478 146.341
R1768 VDD.n1476 VDD.n1147 146.341
R1769 VDD.n1472 VDD.n1471 146.341
R1770 VDD.n1469 VDD.n1154 146.341
R1771 VDD.n1299 VDD.n1161 146.341
R1772 VDD.n1297 VDD.n1296 146.341
R1773 VDD.n1294 VDD.n1163 146.341
R1774 VDD.n1290 VDD.n1289 146.341
R1775 VDD.n1287 VDD.n1170 146.341
R1776 VDD.n1281 VDD.n1280 146.341
R1777 VDD.n1278 VDD.n1178 146.341
R1778 VDD.n1274 VDD.n1273 146.341
R1779 VDD.n1271 VDD.n1184 146.341
R1780 VDD.n1267 VDD.n1266 146.341
R1781 VDD.n1264 VDD.n1191 146.341
R1782 VDD.n1260 VDD.n1259 146.341
R1783 VDD.n1257 VDD.n1198 146.341
R1784 VDD.n1253 VDD.n1252 146.341
R1785 VDD.n1250 VDD.n1205 146.341
R1786 VDD.n1244 VDD.n1243 146.341
R1787 VDD.n1241 VDD.n1213 146.341
R1788 VDD.n1237 VDD.n1236 146.341
R1789 VDD.n1234 VDD.n1219 146.341
R1790 VDD.n1230 VDD.n1229 146.341
R1791 VDD.n1227 VDD.n1225 146.341
R1792 VDD.n631 VDD.n630 146.341
R1793 VDD.n643 VDD.n632 146.341
R1794 VDD.n636 VDD.n635 146.341
R1795 VDD.n1003 VDD.n784 146.341
R1796 VDD.n1003 VDD.n780 146.341
R1797 VDD.n1009 VDD.n780 146.341
R1798 VDD.n1009 VDD.n771 146.341
R1799 VDD.n1019 VDD.n771 146.341
R1800 VDD.n1019 VDD.n767 146.341
R1801 VDD.n1025 VDD.n767 146.341
R1802 VDD.n1025 VDD.n760 146.341
R1803 VDD.n1035 VDD.n760 146.341
R1804 VDD.n1035 VDD.n756 146.341
R1805 VDD.n1041 VDD.n756 146.341
R1806 VDD.n1041 VDD.n747 146.341
R1807 VDD.n1051 VDD.n747 146.341
R1808 VDD.n1051 VDD.n743 146.341
R1809 VDD.n1057 VDD.n743 146.341
R1810 VDD.n1057 VDD.n736 146.341
R1811 VDD.n1068 VDD.n736 146.341
R1812 VDD.n1068 VDD.n732 146.341
R1813 VDD.n1074 VDD.n732 146.341
R1814 VDD.n1074 VDD.n693 146.341
R1815 VDD.n1084 VDD.n693 146.341
R1816 VDD.n1084 VDD.n689 146.341
R1817 VDD.n1090 VDD.n689 146.341
R1818 VDD.n1090 VDD.n682 146.341
R1819 VDD.n1100 VDD.n682 146.341
R1820 VDD.n1100 VDD.n678 146.341
R1821 VDD.n1106 VDD.n678 146.341
R1822 VDD.n1106 VDD.n669 146.341
R1823 VDD.n1116 VDD.n669 146.341
R1824 VDD.n1116 VDD.n665 146.341
R1825 VDD.n1122 VDD.n665 146.341
R1826 VDD.n1122 VDD.n658 146.341
R1827 VDD.n1132 VDD.n658 146.341
R1828 VDD.n1132 VDD.n654 146.341
R1829 VDD.n1138 VDD.n654 146.341
R1830 VDD.n1138 VDD.n640 146.341
R1831 VDD.n1487 VDD.n640 146.341
R1832 VDD.n992 VDD.n790 146.341
R1833 VDD.n992 VDD.n819 146.341
R1834 VDD.n823 VDD.n822 146.341
R1835 VDD.n825 VDD.n824 146.341
R1836 VDD.n829 VDD.n828 146.341
R1837 VDD.n831 VDD.n830 146.341
R1838 VDD.n835 VDD.n834 146.341
R1839 VDD.n837 VDD.n836 146.341
R1840 VDD.n965 VDD.n840 146.341
R1841 VDD.n842 VDD.n841 146.341
R1842 VDD.n846 VDD.n845 146.341
R1843 VDD.n848 VDD.n847 146.341
R1844 VDD.n852 VDD.n851 146.341
R1845 VDD.n854 VDD.n853 146.341
R1846 VDD.n858 VDD.n857 146.341
R1847 VDD.n860 VDD.n859 146.341
R1848 VDD.n864 VDD.n863 146.341
R1849 VDD.n866 VDD.n865 146.341
R1850 VDD.n932 VDD.n869 146.341
R1851 VDD.n871 VDD.n870 146.341
R1852 VDD.n875 VDD.n874 146.341
R1853 VDD.n877 VDD.n876 146.341
R1854 VDD.n881 VDD.n880 146.341
R1855 VDD.n883 VDD.n882 146.341
R1856 VDD.n887 VDD.n886 146.341
R1857 VDD.n889 VDD.n888 146.341
R1858 VDD.n893 VDD.n892 146.341
R1859 VDD.n895 VDD.n894 146.341
R1860 VDD.n898 VDD.n818 146.341
R1861 VDD.n1001 VDD.n786 146.341
R1862 VDD.n1001 VDD.n778 146.341
R1863 VDD.n1011 VDD.n778 146.341
R1864 VDD.n1011 VDD.n774 146.341
R1865 VDD.n1017 VDD.n774 146.341
R1866 VDD.n1017 VDD.n766 146.341
R1867 VDD.n1027 VDD.n766 146.341
R1868 VDD.n1027 VDD.n762 146.341
R1869 VDD.n1033 VDD.n762 146.341
R1870 VDD.n1033 VDD.n754 146.341
R1871 VDD.n1043 VDD.n754 146.341
R1872 VDD.n1043 VDD.n750 146.341
R1873 VDD.n1049 VDD.n750 146.341
R1874 VDD.n1049 VDD.n742 146.341
R1875 VDD.n1059 VDD.n742 146.341
R1876 VDD.n1059 VDD.n738 146.341
R1877 VDD.n1066 VDD.n738 146.341
R1878 VDD.n1066 VDD.n730 146.341
R1879 VDD.n1076 VDD.n730 146.341
R1880 VDD.n1076 VDD.n696 146.341
R1881 VDD.n1082 VDD.n696 146.341
R1882 VDD.n1082 VDD.n688 146.341
R1883 VDD.n1092 VDD.n688 146.341
R1884 VDD.n1092 VDD.n684 146.341
R1885 VDD.n1098 VDD.n684 146.341
R1886 VDD.n1098 VDD.n676 146.341
R1887 VDD.n1108 VDD.n676 146.341
R1888 VDD.n1108 VDD.n672 146.341
R1889 VDD.n1114 VDD.n672 146.341
R1890 VDD.n1114 VDD.n664 146.341
R1891 VDD.n1124 VDD.n664 146.341
R1892 VDD.n1124 VDD.n660 146.341
R1893 VDD.n1130 VDD.n660 146.341
R1894 VDD.n1130 VDD.n652 146.341
R1895 VDD.n1140 VDD.n652 146.341
R1896 VDD.n1140 VDD.n647 146.341
R1897 VDD.n1485 VDD.n647 146.341
R1898 VDD.n646 VDD.t26 145.696
R1899 VDD.n2273 VDD.t82 145.696
R1900 VDD.n1348 VDD.t73 144.964
R1901 VDD.n525 VDD.t65 144.964
R1902 VDD.n1333 VDD.t96 144.964
R1903 VDD.n509 VDD.t92 144.964
R1904 VDD.n2027 VDD.t83 144.964
R1905 VDD.n2027 VDD.t84 144.964
R1906 VDD.n1790 VDD.t87 144.964
R1907 VDD.n388 VDD.t48 144.964
R1908 VDD.n1762 VDD.t80 144.964
R1909 VDD.n360 VDD.t38 144.964
R1910 VDD.n617 VDD.t27 144.964
R1911 VDD.n617 VDD.t28 144.964
R1912 VDD.n900 VDD.t42 139.282
R1913 VDD.n933 VDD.t35 139.282
R1914 VDD.n966 VDD.t69 139.282
R1915 VDD.n1492 VDD.t30 139.282
R1916 VDD.n1207 VDD.t61 139.282
R1917 VDD.n1172 VDD.t23 139.282
R1918 VDD.n199 VDD.t58 139.282
R1919 VDD.n166 VDD.t89 139.282
R1920 VDD.n131 VDD.t52 139.282
R1921 VDD.n340 VDD.t46 139.282
R1922 VDD.n2242 VDD.t76 139.282
R1923 VDD.n2159 VDD.t56 139.282
R1924 VDD.n9 VDD.n7 119.439
R1925 VDD.n2 VDD.n0 119.439
R1926 VDD.n1349 VDD.t72 119.169
R1927 VDD.n526 VDD.t66 119.169
R1928 VDD.n1334 VDD.t95 119.169
R1929 VDD.n510 VDD.t93 119.169
R1930 VDD.n1791 VDD.t86 119.169
R1931 VDD.n389 VDD.t49 119.169
R1932 VDD.n1763 VDD.t79 119.169
R1933 VDD.n361 VDD.t39 119.169
R1934 VDD.n9 VDD.n8 118.865
R1935 VDD.n11 VDD.n10 118.865
R1936 VDD.n13 VDD.n12 118.865
R1937 VDD.n6 VDD.n5 118.865
R1938 VDD.n4 VDD.n3 118.865
R1939 VDD.n2 VDD.n1 118.865
R1940 VDD.n901 VDD.t41 113.489
R1941 VDD.n934 VDD.t34 113.489
R1942 VDD.n967 VDD.t68 113.489
R1943 VDD.n1493 VDD.t31 113.489
R1944 VDD.n1208 VDD.t62 113.489
R1945 VDD.n1173 VDD.t24 113.489
R1946 VDD.n200 VDD.t59 113.489
R1947 VDD.n167 VDD.t90 113.489
R1948 VDD.n132 VDD.t53 113.489
R1949 VDD.n341 VDD.t45 113.489
R1950 VDD.n2243 VDD.t75 113.489
R1951 VDD.n2160 VDD.t55 113.489
R1952 VDD.n2116 VDD.n2115 99.5127
R1953 VDD.n2113 VDD.n375 99.5127
R1954 VDD.n2109 VDD.n2108 99.5127
R1955 VDD.n2106 VDD.n378 99.5127
R1956 VDD.n2102 VDD.n2101 99.5127
R1957 VDD.n2099 VDD.n2097 99.5127
R1958 VDD.n2095 VDD.n381 99.5127
R1959 VDD.n2091 VDD.n2090 99.5127
R1960 VDD.n2088 VDD.n384 99.5127
R1961 VDD.n2084 VDD.n2083 99.5127
R1962 VDD.n2081 VDD.n387 99.5127
R1963 VDD.n1901 VDD.n477 99.5127
R1964 VDD.n1897 VDD.n477 99.5127
R1965 VDD.n1897 VDD.n471 99.5127
R1966 VDD.n1894 VDD.n471 99.5127
R1967 VDD.n1894 VDD.n465 99.5127
R1968 VDD.n1891 VDD.n465 99.5127
R1969 VDD.n1891 VDD.n459 99.5127
R1970 VDD.n1888 VDD.n459 99.5127
R1971 VDD.n1888 VDD.n453 99.5127
R1972 VDD.n1885 VDD.n453 99.5127
R1973 VDD.n1885 VDD.n447 99.5127
R1974 VDD.n1787 VDD.n447 99.5127
R1975 VDD.n1787 VDD.n441 99.5127
R1976 VDD.n1784 VDD.n441 99.5127
R1977 VDD.n1784 VDD.n435 99.5127
R1978 VDD.n1781 VDD.n435 99.5127
R1979 VDD.n1781 VDD.n430 99.5127
R1980 VDD.n1778 VDD.n430 99.5127
R1981 VDD.n1778 VDD.n424 99.5127
R1982 VDD.n1775 VDD.n424 99.5127
R1983 VDD.n1775 VDD.n418 99.5127
R1984 VDD.n1772 VDD.n418 99.5127
R1985 VDD.n1772 VDD.n412 99.5127
R1986 VDD.n1769 VDD.n412 99.5127
R1987 VDD.n1769 VDD.n406 99.5127
R1988 VDD.n1766 VDD.n406 99.5127
R1989 VDD.n1766 VDD.n399 99.5127
R1990 VDD.n399 VDD.n392 99.5127
R1991 VDD.n2070 VDD.n392 99.5127
R1992 VDD.n2071 VDD.n2070 99.5127
R1993 VDD.n2071 VDD.n368 99.5127
R1994 VDD.n2076 VDD.n368 99.5127
R1995 VDD.n1943 VDD.n481 99.5127
R1996 VDD.n1943 VDD.n1761 99.5127
R1997 VDD.n1939 VDD.n1938 99.5127
R1998 VDD.n1935 VDD.n1934 99.5127
R1999 VDD.n1931 VDD.n1930 99.5127
R2000 VDD.n1927 VDD.n1926 99.5127
R2001 VDD.n1923 VDD.n1922 99.5127
R2002 VDD.n1919 VDD.n1918 99.5127
R2003 VDD.n1915 VDD.n1914 99.5127
R2004 VDD.n1911 VDD.n1910 99.5127
R2005 VDD.n1906 VDD.n1905 99.5127
R2006 VDD.n1950 VDD.n479 99.5127
R2007 VDD.n1950 VDD.n469 99.5127
R2008 VDD.n1958 VDD.n469 99.5127
R2009 VDD.n1958 VDD.n467 99.5127
R2010 VDD.n1962 VDD.n467 99.5127
R2011 VDD.n1962 VDD.n457 99.5127
R2012 VDD.n1970 VDD.n457 99.5127
R2013 VDD.n1970 VDD.n455 99.5127
R2014 VDD.n1974 VDD.n455 99.5127
R2015 VDD.n1974 VDD.n446 99.5127
R2016 VDD.n1982 VDD.n446 99.5127
R2017 VDD.n1982 VDD.n444 99.5127
R2018 VDD.n1986 VDD.n444 99.5127
R2019 VDD.n1986 VDD.n434 99.5127
R2020 VDD.n1994 VDD.n434 99.5127
R2021 VDD.n1994 VDD.n432 99.5127
R2022 VDD.n1998 VDD.n432 99.5127
R2023 VDD.n1998 VDD.n422 99.5127
R2024 VDD.n2006 VDD.n422 99.5127
R2025 VDD.n2006 VDD.n420 99.5127
R2026 VDD.n2010 VDD.n420 99.5127
R2027 VDD.n2010 VDD.n410 99.5127
R2028 VDD.n2018 VDD.n410 99.5127
R2029 VDD.n2018 VDD.n408 99.5127
R2030 VDD.n2022 VDD.n408 99.5127
R2031 VDD.n2022 VDD.n397 99.5127
R2032 VDD.n2064 VDD.n397 99.5127
R2033 VDD.n2064 VDD.n395 99.5127
R2034 VDD.n2068 VDD.n395 99.5127
R2035 VDD.n2068 VDD.n371 99.5127
R2036 VDD.n2120 VDD.n371 99.5127
R2037 VDD.n2120 VDD.n372 99.5127
R2038 VDD.n1737 VDD.n507 99.5127
R2039 VDD.n1733 VDD.n1732 99.5127
R2040 VDD.n1729 VDD.n1728 99.5127
R2041 VDD.n1725 VDD.n1724 99.5127
R2042 VDD.n1721 VDD.n1720 99.5127
R2043 VDD.n1717 VDD.n1716 99.5127
R2044 VDD.n1713 VDD.n1712 99.5127
R2045 VDD.n1709 VDD.n1708 99.5127
R2046 VDD.n1705 VDD.n1704 99.5127
R2047 VDD.n1701 VDD.n1700 99.5127
R2048 VDD.n1696 VDD.n1695 99.5127
R2049 VDD.n1439 VDD.n614 99.5127
R2050 VDD.n1439 VDD.n607 99.5127
R2051 VDD.n1436 VDD.n607 99.5127
R2052 VDD.n1436 VDD.n601 99.5127
R2053 VDD.n1433 VDD.n601 99.5127
R2054 VDD.n1433 VDD.n596 99.5127
R2055 VDD.n1430 VDD.n596 99.5127
R2056 VDD.n1430 VDD.n590 99.5127
R2057 VDD.n1427 VDD.n590 99.5127
R2058 VDD.n1427 VDD.n584 99.5127
R2059 VDD.n1424 VDD.n584 99.5127
R2060 VDD.n1424 VDD.n578 99.5127
R2061 VDD.n1421 VDD.n578 99.5127
R2062 VDD.n1421 VDD.n572 99.5127
R2063 VDD.n1418 VDD.n572 99.5127
R2064 VDD.n1418 VDD.n566 99.5127
R2065 VDD.n1415 VDD.n566 99.5127
R2066 VDD.n1415 VDD.n560 99.5127
R2067 VDD.n1343 VDD.n560 99.5127
R2068 VDD.n1343 VDD.n554 99.5127
R2069 VDD.n1340 VDD.n554 99.5127
R2070 VDD.n1340 VDD.n548 99.5127
R2071 VDD.n1337 VDD.n548 99.5127
R2072 VDD.n1337 VDD.n542 99.5127
R2073 VDD.n542 VDD.n533 99.5127
R2074 VDD.n1616 VDD.n533 99.5127
R2075 VDD.n1616 VDD.n531 99.5127
R2076 VDD.n1622 VDD.n531 99.5127
R2077 VDD.n1622 VDD.n519 99.5127
R2078 VDD.n519 VDD.n512 99.5127
R2079 VDD.n1690 VDD.n512 99.5127
R2080 VDD.n1691 VDD.n1690 99.5127
R2081 VDD.n1311 VDD.n1310 99.5127
R2082 VDD.n1313 VDD.n1311 99.5127
R2083 VDD.n1317 VDD.n1306 99.5127
R2084 VDD.n1321 VDD.n1319 99.5127
R2085 VDD.n1325 VDD.n1304 99.5127
R2086 VDD.n1464 VDD.n1327 99.5127
R2087 VDD.n1462 VDD.n1461 99.5127
R2088 VDD.n1458 VDD.n1457 99.5127
R2089 VDD.n1455 VDD.n1330 99.5127
R2090 VDD.n1451 VDD.n1449 99.5127
R2091 VDD.n1447 VDD.n1332 99.5127
R2092 VDD.n1533 VDD.n610 99.5127
R2093 VDD.n1537 VDD.n610 99.5127
R2094 VDD.n1537 VDD.n600 99.5127
R2095 VDD.n1545 VDD.n600 99.5127
R2096 VDD.n1545 VDD.n598 99.5127
R2097 VDD.n1549 VDD.n598 99.5127
R2098 VDD.n1549 VDD.n588 99.5127
R2099 VDD.n1557 VDD.n588 99.5127
R2100 VDD.n1557 VDD.n586 99.5127
R2101 VDD.n1561 VDD.n586 99.5127
R2102 VDD.n1561 VDD.n576 99.5127
R2103 VDD.n1569 VDD.n576 99.5127
R2104 VDD.n1569 VDD.n574 99.5127
R2105 VDD.n1573 VDD.n574 99.5127
R2106 VDD.n1573 VDD.n564 99.5127
R2107 VDD.n1581 VDD.n564 99.5127
R2108 VDD.n1581 VDD.n562 99.5127
R2109 VDD.n1585 VDD.n562 99.5127
R2110 VDD.n1585 VDD.n552 99.5127
R2111 VDD.n1593 VDD.n552 99.5127
R2112 VDD.n1593 VDD.n550 99.5127
R2113 VDD.n1597 VDD.n550 99.5127
R2114 VDD.n1597 VDD.n540 99.5127
R2115 VDD.n1609 VDD.n540 99.5127
R2116 VDD.n1609 VDD.n537 99.5127
R2117 VDD.n1614 VDD.n537 99.5127
R2118 VDD.n1614 VDD.n538 99.5127
R2119 VDD.n538 VDD.n518 99.5127
R2120 VDD.n1684 VDD.n518 99.5127
R2121 VDD.n1684 VDD.n516 99.5127
R2122 VDD.n1688 VDD.n516 99.5127
R2123 VDD.n1688 VDD.n506 99.5127
R2124 VDD.n2053 VDD.n2029 99.5127
R2125 VDD.n2049 VDD.n2048 99.5127
R2126 VDD.n2046 VDD.n2032 99.5127
R2127 VDD.n2042 VDD.n2041 99.5127
R2128 VDD.n2039 VDD.n2036 99.5127
R2129 VDD.n2146 VDD.n353 99.5127
R2130 VDD.n2144 VDD.n2143 99.5127
R2131 VDD.n2141 VDD.n356 99.5127
R2132 VDD.n2137 VDD.n2136 99.5127
R2133 VDD.n2134 VDD.n359 99.5127
R2134 VDD.n2129 VDD.n2128 99.5127
R2135 VDD.n1838 VDD.n478 99.5127
R2136 VDD.n1841 VDD.n478 99.5127
R2137 VDD.n1841 VDD.n472 99.5127
R2138 VDD.n1844 VDD.n472 99.5127
R2139 VDD.n1844 VDD.n466 99.5127
R2140 VDD.n1847 VDD.n466 99.5127
R2141 VDD.n1847 VDD.n460 99.5127
R2142 VDD.n1850 VDD.n460 99.5127
R2143 VDD.n1850 VDD.n454 99.5127
R2144 VDD.n1883 VDD.n454 99.5127
R2145 VDD.n1883 VDD.n448 99.5127
R2146 VDD.n1879 VDD.n448 99.5127
R2147 VDD.n1879 VDD.n442 99.5127
R2148 VDD.n1876 VDD.n442 99.5127
R2149 VDD.n1876 VDD.n436 99.5127
R2150 VDD.n1873 VDD.n436 99.5127
R2151 VDD.n1873 VDD.n431 99.5127
R2152 VDD.n1870 VDD.n431 99.5127
R2153 VDD.n1870 VDD.n425 99.5127
R2154 VDD.n1867 VDD.n425 99.5127
R2155 VDD.n1867 VDD.n419 99.5127
R2156 VDD.n1864 VDD.n419 99.5127
R2157 VDD.n1864 VDD.n413 99.5127
R2158 VDD.n1861 VDD.n413 99.5127
R2159 VDD.n1861 VDD.n407 99.5127
R2160 VDD.n1858 VDD.n407 99.5127
R2161 VDD.n1858 VDD.n400 99.5127
R2162 VDD.n1855 VDD.n400 99.5127
R2163 VDD.n1855 VDD.n393 99.5127
R2164 VDD.n393 VDD.n366 99.5127
R2165 VDD.n2122 VDD.n366 99.5127
R2166 VDD.n2122 VDD.n364 99.5127
R2167 VDD.n1797 VDD.n1796 99.5127
R2168 VDD.n1801 VDD.n1800 99.5127
R2169 VDD.n1805 VDD.n1804 99.5127
R2170 VDD.n1809 VDD.n1808 99.5127
R2171 VDD.n1813 VDD.n1812 99.5127
R2172 VDD.n1817 VDD.n1816 99.5127
R2173 VDD.n1821 VDD.n1820 99.5127
R2174 VDD.n1825 VDD.n1824 99.5127
R2175 VDD.n1829 VDD.n1828 99.5127
R2176 VDD.n1833 VDD.n1832 99.5127
R2177 VDD.n1835 VDD.n1760 99.5127
R2178 VDD.n1952 VDD.n475 99.5127
R2179 VDD.n1952 VDD.n473 99.5127
R2180 VDD.n1956 VDD.n473 99.5127
R2181 VDD.n1956 VDD.n463 99.5127
R2182 VDD.n1964 VDD.n463 99.5127
R2183 VDD.n1964 VDD.n461 99.5127
R2184 VDD.n1968 VDD.n461 99.5127
R2185 VDD.n1968 VDD.n451 99.5127
R2186 VDD.n1976 VDD.n451 99.5127
R2187 VDD.n1976 VDD.n449 99.5127
R2188 VDD.n1980 VDD.n449 99.5127
R2189 VDD.n1980 VDD.n439 99.5127
R2190 VDD.n1988 VDD.n439 99.5127
R2191 VDD.n1988 VDD.n437 99.5127
R2192 VDD.n1992 VDD.n437 99.5127
R2193 VDD.n1992 VDD.n428 99.5127
R2194 VDD.n2000 VDD.n428 99.5127
R2195 VDD.n2000 VDD.n426 99.5127
R2196 VDD.n2004 VDD.n426 99.5127
R2197 VDD.n2004 VDD.n416 99.5127
R2198 VDD.n2012 VDD.n416 99.5127
R2199 VDD.n2012 VDD.n414 99.5127
R2200 VDD.n2016 VDD.n414 99.5127
R2201 VDD.n2016 VDD.n404 99.5127
R2202 VDD.n2024 VDD.n404 99.5127
R2203 VDD.n2024 VDD.n401 99.5127
R2204 VDD.n2062 VDD.n401 99.5127
R2205 VDD.n2062 VDD.n402 99.5127
R2206 VDD.n402 VDD.n394 99.5127
R2207 VDD.n2057 VDD.n394 99.5127
R2208 VDD.n2057 VDD.n370 99.5127
R2209 VDD.n2054 VDD.n370 99.5127
R2210 VDD.n1673 VDD.n1672 99.5127
R2211 VDD.n1669 VDD.n1668 99.5127
R2212 VDD.n1665 VDD.n1664 99.5127
R2213 VDD.n1661 VDD.n1660 99.5127
R2214 VDD.n1657 VDD.n1656 99.5127
R2215 VDD.n1653 VDD.n1652 99.5127
R2216 VDD.n1649 VDD.n1648 99.5127
R2217 VDD.n1645 VDD.n1644 99.5127
R2218 VDD.n1641 VDD.n1640 99.5127
R2219 VDD.n1637 VDD.n1636 99.5127
R2220 VDD.n1633 VDD.n494 99.5127
R2221 VDD.n1375 VDD.n615 99.5127
R2222 VDD.n1375 VDD.n608 99.5127
R2223 VDD.n1378 VDD.n608 99.5127
R2224 VDD.n1378 VDD.n602 99.5127
R2225 VDD.n1381 VDD.n602 99.5127
R2226 VDD.n1381 VDD.n597 99.5127
R2227 VDD.n1384 VDD.n597 99.5127
R2228 VDD.n1384 VDD.n591 99.5127
R2229 VDD.n1387 VDD.n591 99.5127
R2230 VDD.n1387 VDD.n585 99.5127
R2231 VDD.n1390 VDD.n585 99.5127
R2232 VDD.n1390 VDD.n579 99.5127
R2233 VDD.n1393 VDD.n579 99.5127
R2234 VDD.n1393 VDD.n573 99.5127
R2235 VDD.n1396 VDD.n573 99.5127
R2236 VDD.n1396 VDD.n567 99.5127
R2237 VDD.n1413 VDD.n567 99.5127
R2238 VDD.n1413 VDD.n561 99.5127
R2239 VDD.n1409 VDD.n561 99.5127
R2240 VDD.n1409 VDD.n555 99.5127
R2241 VDD.n1406 VDD.n555 99.5127
R2242 VDD.n1406 VDD.n549 99.5127
R2243 VDD.n1403 VDD.n549 99.5127
R2244 VDD.n1403 VDD.n543 99.5127
R2245 VDD.n1400 VDD.n543 99.5127
R2246 VDD.n1400 VDD.n535 99.5127
R2247 VDD.n535 VDD.n529 99.5127
R2248 VDD.n1624 VDD.n529 99.5127
R2249 VDD.n1624 VDD.n520 99.5127
R2250 VDD.n1627 VDD.n520 99.5127
R2251 VDD.n1627 VDD.n514 99.5127
R2252 VDD.n1630 VDD.n514 99.5127
R2253 VDD.n1526 VDD.n1524 99.5127
R2254 VDD.n1522 VDD.n619 99.5127
R2255 VDD.n1518 VDD.n1516 99.5127
R2256 VDD.n1514 VDD.n621 99.5127
R2257 VDD.n1510 VDD.n1508 99.5127
R2258 VDD.n1506 VDD.n623 99.5127
R2259 VDD.n1356 VDD.n1354 99.5127
R2260 VDD.n1360 VDD.n1351 99.5127
R2261 VDD.n1364 VDD.n1362 99.5127
R2262 VDD.n1369 VDD.n1347 99.5127
R2263 VDD.n1372 VDD.n1371 99.5127
R2264 VDD.n1531 VDD.n605 99.5127
R2265 VDD.n1539 VDD.n605 99.5127
R2266 VDD.n1539 VDD.n603 99.5127
R2267 VDD.n1543 VDD.n603 99.5127
R2268 VDD.n1543 VDD.n594 99.5127
R2269 VDD.n1551 VDD.n594 99.5127
R2270 VDD.n1551 VDD.n592 99.5127
R2271 VDD.n1555 VDD.n592 99.5127
R2272 VDD.n1555 VDD.n582 99.5127
R2273 VDD.n1563 VDD.n582 99.5127
R2274 VDD.n1563 VDD.n580 99.5127
R2275 VDD.n1567 VDD.n580 99.5127
R2276 VDD.n1567 VDD.n570 99.5127
R2277 VDD.n1575 VDD.n570 99.5127
R2278 VDD.n1575 VDD.n568 99.5127
R2279 VDD.n1579 VDD.n568 99.5127
R2280 VDD.n1579 VDD.n559 99.5127
R2281 VDD.n1587 VDD.n559 99.5127
R2282 VDD.n1587 VDD.n557 99.5127
R2283 VDD.n1591 VDD.n557 99.5127
R2284 VDD.n1591 VDD.n547 99.5127
R2285 VDD.n1599 VDD.n547 99.5127
R2286 VDD.n1599 VDD.n544 99.5127
R2287 VDD.n1607 VDD.n544 99.5127
R2288 VDD.n1607 VDD.n545 99.5127
R2289 VDD.n545 VDD.n536 99.5127
R2290 VDD.n1602 VDD.n536 99.5127
R2291 VDD.n1602 VDD.n522 99.5127
R2292 VDD.n1682 VDD.n522 99.5127
R2293 VDD.n1682 VDD.n523 99.5127
R2294 VDD.n523 VDD.n515 99.5127
R2295 VDD.n1677 VDD.n515 99.5127
R2296 VDD.t192 VDD.t12 97.6278
R2297 VDD.n2028 VDD.n2027 82.6045
R2298 VDD.n1529 VDD.n617 82.6045
R2299 VDD.n36 VDD.t129 79.3769
R2300 VDD.n26 VDD.t171 79.3769
R2301 VDD.n17 VDD.t176 79.3769
R2302 VDD.n718 VDD.t155 79.3769
R2303 VDD.n708 VDD.t187 79.3769
R2304 VDD.n699 VDD.t162 79.3769
R2305 VDD.n43 VDD.t111 78.8036
R2306 VDD.n33 VDD.t158 78.8036
R2307 VDD.n24 VDD.t121 78.8036
R2308 VDD.n725 VDD.t127 78.8036
R2309 VDD.n715 VDD.t170 78.8036
R2310 VDD.n706 VDD.t130 78.8036
R2311 VDD.n42 VDD.n41 74.1601
R2312 VDD.n40 VDD.n39 74.1601
R2313 VDD.n38 VDD.n37 74.1601
R2314 VDD.n36 VDD.n35 74.1601
R2315 VDD.n32 VDD.n31 74.1601
R2316 VDD.n30 VDD.n29 74.1601
R2317 VDD.n28 VDD.n27 74.1601
R2318 VDD.n26 VDD.n25 74.1601
R2319 VDD.n23 VDD.n22 74.1601
R2320 VDD.n21 VDD.n20 74.1601
R2321 VDD.n19 VDD.n18 74.1601
R2322 VDD.n17 VDD.n16 74.1601
R2323 VDD.n718 VDD.n717 74.1601
R2324 VDD.n720 VDD.n719 74.1601
R2325 VDD.n722 VDD.n721 74.1601
R2326 VDD.n724 VDD.n723 74.1601
R2327 VDD.n708 VDD.n707 74.1601
R2328 VDD.n710 VDD.n709 74.1601
R2329 VDD.n712 VDD.n711 74.1601
R2330 VDD.n714 VDD.n713 74.1601
R2331 VDD.n699 VDD.n698 74.1601
R2332 VDD.n701 VDD.n700 74.1601
R2333 VDD.n703 VDD.n702 74.1601
R2334 VDD.n705 VDD.n704 74.1601
R2335 VDD.n1944 VDD.n1749 72.8958
R2336 VDD.n1944 VDD.n1750 72.8958
R2337 VDD.n1944 VDD.n1751 72.8958
R2338 VDD.n1944 VDD.n1752 72.8958
R2339 VDD.n1944 VDD.n1753 72.8958
R2340 VDD.n1944 VDD.n1754 72.8958
R2341 VDD.n1944 VDD.n1755 72.8958
R2342 VDD.n1944 VDD.n1756 72.8958
R2343 VDD.n1944 VDD.n1757 72.8958
R2344 VDD.n1944 VDD.n1758 72.8958
R2345 VDD.n1944 VDD.n1759 72.8958
R2346 VDD.n2127 VDD.n354 72.8958
R2347 VDD.n363 VDD.n354 72.8958
R2348 VDD.n2135 VDD.n354 72.8958
R2349 VDD.n358 VDD.n354 72.8958
R2350 VDD.n2142 VDD.n354 72.8958
R2351 VDD.n2145 VDD.n354 72.8958
R2352 VDD.n2035 VDD.n354 72.8958
R2353 VDD.n2040 VDD.n354 72.8958
R2354 VDD.n2034 VDD.n354 72.8958
R2355 VDD.n2047 VDD.n354 72.8958
R2356 VDD.n2031 VDD.n354 72.8958
R2357 VDD.n1309 VDD.n613 72.8958
R2358 VDD.n1312 VDD.n613 72.8958
R2359 VDD.n1318 VDD.n613 72.8958
R2360 VDD.n1320 VDD.n613 72.8958
R2361 VDD.n1326 VDD.n613 72.8958
R2362 VDD.n1463 VDD.n613 72.8958
R2363 VDD.n1328 VDD.n613 72.8958
R2364 VDD.n1456 VDD.n613 72.8958
R2365 VDD.n1450 VDD.n613 72.8958
R2366 VDD.n1448 VDD.n613 72.8958
R2367 VDD.n1442 VDD.n613 72.8958
R2368 VDD.n1738 VDD.n495 72.8958
R2369 VDD.n1738 VDD.n496 72.8958
R2370 VDD.n1738 VDD.n497 72.8958
R2371 VDD.n1738 VDD.n498 72.8958
R2372 VDD.n1738 VDD.n499 72.8958
R2373 VDD.n1738 VDD.n500 72.8958
R2374 VDD.n1738 VDD.n501 72.8958
R2375 VDD.n1738 VDD.n502 72.8958
R2376 VDD.n1738 VDD.n503 72.8958
R2377 VDD.n1738 VDD.n504 72.8958
R2378 VDD.n1738 VDD.n505 72.8958
R2379 VDD.n1945 VDD.n1944 72.8958
R2380 VDD.n1944 VDD.n1739 72.8958
R2381 VDD.n1944 VDD.n1740 72.8958
R2382 VDD.n1944 VDD.n1741 72.8958
R2383 VDD.n1944 VDD.n1742 72.8958
R2384 VDD.n1944 VDD.n1743 72.8958
R2385 VDD.n1944 VDD.n1744 72.8958
R2386 VDD.n1944 VDD.n1745 72.8958
R2387 VDD.n1944 VDD.n1746 72.8958
R2388 VDD.n1944 VDD.n1747 72.8958
R2389 VDD.n1944 VDD.n1748 72.8958
R2390 VDD.n2075 VDD.n354 72.8958
R2391 VDD.n2082 VDD.n354 72.8958
R2392 VDD.n386 VDD.n354 72.8958
R2393 VDD.n2089 VDD.n354 72.8958
R2394 VDD.n383 VDD.n354 72.8958
R2395 VDD.n2096 VDD.n354 72.8958
R2396 VDD.n2100 VDD.n354 72.8958
R2397 VDD.n380 VDD.n354 72.8958
R2398 VDD.n2107 VDD.n354 72.8958
R2399 VDD.n377 VDD.n354 72.8958
R2400 VDD.n2114 VDD.n354 72.8958
R2401 VDD.n1738 VDD.n493 72.8958
R2402 VDD.n1738 VDD.n492 72.8958
R2403 VDD.n1738 VDD.n491 72.8958
R2404 VDD.n1738 VDD.n490 72.8958
R2405 VDD.n1738 VDD.n489 72.8958
R2406 VDD.n1738 VDD.n488 72.8958
R2407 VDD.n1738 VDD.n487 72.8958
R2408 VDD.n1738 VDD.n486 72.8958
R2409 VDD.n1738 VDD.n485 72.8958
R2410 VDD.n1738 VDD.n484 72.8958
R2411 VDD.n1738 VDD.n483 72.8958
R2412 VDD.n1525 VDD.n613 72.8958
R2413 VDD.n1523 VDD.n613 72.8958
R2414 VDD.n1517 VDD.n613 72.8958
R2415 VDD.n1515 VDD.n613 72.8958
R2416 VDD.n1509 VDD.n613 72.8958
R2417 VDD.n1507 VDD.n613 72.8958
R2418 VDD.n1353 VDD.n613 72.8958
R2419 VDD.n1355 VDD.n613 72.8958
R2420 VDD.n1361 VDD.n613 72.8958
R2421 VDD.n1363 VDD.n613 72.8958
R2422 VDD.n1370 VDD.n613 72.8958
R2423 VDD.n994 VDD.n993 66.2847
R2424 VDD.n993 VDD.n791 66.2847
R2425 VDD.n993 VDD.n792 66.2847
R2426 VDD.n993 VDD.n793 66.2847
R2427 VDD.n993 VDD.n794 66.2847
R2428 VDD.n993 VDD.n795 66.2847
R2429 VDD.n993 VDD.n796 66.2847
R2430 VDD.n993 VDD.n797 66.2847
R2431 VDD.n993 VDD.n798 66.2847
R2432 VDD.n993 VDD.n799 66.2847
R2433 VDD.n993 VDD.n800 66.2847
R2434 VDD.n993 VDD.n801 66.2847
R2435 VDD.n993 VDD.n802 66.2847
R2436 VDD.n993 VDD.n803 66.2847
R2437 VDD.n993 VDD.n804 66.2847
R2438 VDD.n993 VDD.n805 66.2847
R2439 VDD.n993 VDD.n806 66.2847
R2440 VDD.n993 VDD.n807 66.2847
R2441 VDD.n993 VDD.n808 66.2847
R2442 VDD.n993 VDD.n809 66.2847
R2443 VDD.n993 VDD.n810 66.2847
R2444 VDD.n993 VDD.n811 66.2847
R2445 VDD.n993 VDD.n812 66.2847
R2446 VDD.n993 VDD.n813 66.2847
R2447 VDD.n993 VDD.n814 66.2847
R2448 VDD.n993 VDD.n815 66.2847
R2449 VDD.n993 VDD.n816 66.2847
R2450 VDD.n993 VDD.n817 66.2847
R2451 VDD.n646 VDD.n645 66.2847
R2452 VDD.n646 VDD.n644 66.2847
R2453 VDD.n646 VDD.n642 66.2847
R2454 VDD.n1224 VDD.n646 66.2847
R2455 VDD.n1228 VDD.n646 66.2847
R2456 VDD.n1222 VDD.n646 66.2847
R2457 VDD.n1235 VDD.n646 66.2847
R2458 VDD.n1218 VDD.n646 66.2847
R2459 VDD.n1242 VDD.n646 66.2847
R2460 VDD.n1212 VDD.n646 66.2847
R2461 VDD.n1251 VDD.n646 66.2847
R2462 VDD.n1204 VDD.n646 66.2847
R2463 VDD.n1258 VDD.n646 66.2847
R2464 VDD.n1197 VDD.n646 66.2847
R2465 VDD.n1265 VDD.n646 66.2847
R2466 VDD.n1190 VDD.n646 66.2847
R2467 VDD.n1272 VDD.n646 66.2847
R2468 VDD.n1183 VDD.n646 66.2847
R2469 VDD.n1279 VDD.n646 66.2847
R2470 VDD.n1177 VDD.n646 66.2847
R2471 VDD.n1288 VDD.n646 66.2847
R2472 VDD.n1169 VDD.n646 66.2847
R2473 VDD.n1295 VDD.n646 66.2847
R2474 VDD.n1298 VDD.n646 66.2847
R2475 VDD.n1160 VDD.n646 66.2847
R2476 VDD.n1470 VDD.n646 66.2847
R2477 VDD.n1153 VDD.n646 66.2847
R2478 VDD.n1477 VDD.n646 66.2847
R2479 VDD.n1146 VDD.n646 66.2847
R2480 VDD.n2274 VDD.n2273 66.2847
R2481 VDD.n2273 VDD.n275 66.2847
R2482 VDD.n2273 VDD.n276 66.2847
R2483 VDD.n2273 VDD.n277 66.2847
R2484 VDD.n2273 VDD.n278 66.2847
R2485 VDD.n2273 VDD.n279 66.2847
R2486 VDD.n2273 VDD.n280 66.2847
R2487 VDD.n2273 VDD.n281 66.2847
R2488 VDD.n2273 VDD.n282 66.2847
R2489 VDD.n2273 VDD.n283 66.2847
R2490 VDD.n2273 VDD.n284 66.2847
R2491 VDD.n2273 VDD.n285 66.2847
R2492 VDD.n2273 VDD.n286 66.2847
R2493 VDD.n2273 VDD.n287 66.2847
R2494 VDD.n2273 VDD.n288 66.2847
R2495 VDD.n2273 VDD.n289 66.2847
R2496 VDD.n2273 VDD.n290 66.2847
R2497 VDD.n2273 VDD.n291 66.2847
R2498 VDD.n2273 VDD.n292 66.2847
R2499 VDD.n2273 VDD.n293 66.2847
R2500 VDD.n2273 VDD.n294 66.2847
R2501 VDD.n2273 VDD.n295 66.2847
R2502 VDD.n2273 VDD.n296 66.2847
R2503 VDD.n2273 VDD.n297 66.2847
R2504 VDD.n2273 VDD.n298 66.2847
R2505 VDD.n2273 VDD.n299 66.2847
R2506 VDD.n2273 VDD.n300 66.2847
R2507 VDD.n2273 VDD.n301 66.2847
R2508 VDD.n2383 VDD.n98 66.2847
R2509 VDD.n198 VDD.n98 66.2847
R2510 VDD.n2390 VDD.n98 66.2847
R2511 VDD.n191 VDD.n98 66.2847
R2512 VDD.n2397 VDD.n98 66.2847
R2513 VDD.n184 VDD.n98 66.2847
R2514 VDD.n2404 VDD.n98 66.2847
R2515 VDD.n177 VDD.n98 66.2847
R2516 VDD.n2411 VDD.n98 66.2847
R2517 VDD.n171 VDD.n98 66.2847
R2518 VDD.n2420 VDD.n98 66.2847
R2519 VDD.n163 VDD.n98 66.2847
R2520 VDD.n2427 VDD.n98 66.2847
R2521 VDD.n156 VDD.n98 66.2847
R2522 VDD.n2434 VDD.n98 66.2847
R2523 VDD.n149 VDD.n98 66.2847
R2524 VDD.n2441 VDD.n98 66.2847
R2525 VDD.n142 VDD.n98 66.2847
R2526 VDD.n2448 VDD.n98 66.2847
R2527 VDD.n136 VDD.n98 66.2847
R2528 VDD.n2457 VDD.n98 66.2847
R2529 VDD.n128 VDD.n98 66.2847
R2530 VDD.n2464 VDD.n98 66.2847
R2531 VDD.n121 VDD.n98 66.2847
R2532 VDD.n2471 VDD.n98 66.2847
R2533 VDD.n114 VDD.n98 66.2847
R2534 VDD.n2478 VDD.n98 66.2847
R2535 VDD.n2481 VDD.n98 66.2847
R2536 VDD.n102 VDD.n98 66.2847
R2537 VDD.n103 VDD.n102 52.4337
R2538 VDD.n2481 VDD.n2480 52.4337
R2539 VDD.n2478 VDD.n2477 52.4337
R2540 VDD.n2473 VDD.n114 52.4337
R2541 VDD.n2471 VDD.n2470 52.4337
R2542 VDD.n2466 VDD.n121 52.4337
R2543 VDD.n2464 VDD.n2463 52.4337
R2544 VDD.n2459 VDD.n128 52.4337
R2545 VDD.n2457 VDD.n2456 52.4337
R2546 VDD.n2450 VDD.n136 52.4337
R2547 VDD.n2448 VDD.n2447 52.4337
R2548 VDD.n2443 VDD.n142 52.4337
R2549 VDD.n2441 VDD.n2440 52.4337
R2550 VDD.n2436 VDD.n149 52.4337
R2551 VDD.n2434 VDD.n2433 52.4337
R2552 VDD.n2429 VDD.n156 52.4337
R2553 VDD.n2427 VDD.n2426 52.4337
R2554 VDD.n2422 VDD.n163 52.4337
R2555 VDD.n2420 VDD.n2419 52.4337
R2556 VDD.n2413 VDD.n171 52.4337
R2557 VDD.n2411 VDD.n2410 52.4337
R2558 VDD.n2406 VDD.n177 52.4337
R2559 VDD.n2404 VDD.n2403 52.4337
R2560 VDD.n2399 VDD.n184 52.4337
R2561 VDD.n2397 VDD.n2396 52.4337
R2562 VDD.n2392 VDD.n191 52.4337
R2563 VDD.n2390 VDD.n2389 52.4337
R2564 VDD.n2385 VDD.n198 52.4337
R2565 VDD.n2383 VDD.n2382 52.4337
R2566 VDD.n2275 VDD.n2274 52.4337
R2567 VDD.n303 VDD.n275 52.4337
R2568 VDD.n2267 VDD.n276 52.4337
R2569 VDD.n2263 VDD.n277 52.4337
R2570 VDD.n313 VDD.n278 52.4337
R2571 VDD.n2256 VDD.n279 52.4337
R2572 VDD.n2253 VDD.n280 52.4337
R2573 VDD.n2249 VDD.n281 52.4337
R2574 VDD.n2245 VDD.n282 52.4337
R2575 VDD.n2237 VDD.n283 52.4337
R2576 VDD.n2233 VDD.n284 52.4337
R2577 VDD.n2229 VDD.n285 52.4337
R2578 VDD.n2225 VDD.n286 52.4337
R2579 VDD.n2221 VDD.n287 52.4337
R2580 VDD.n2217 VDD.n288 52.4337
R2581 VDD.n2213 VDD.n289 52.4337
R2582 VDD.n2209 VDD.n290 52.4337
R2583 VDD.n2205 VDD.n291 52.4337
R2584 VDD.n2201 VDD.n292 52.4337
R2585 VDD.n2195 VDD.n293 52.4337
R2586 VDD.n2191 VDD.n294 52.4337
R2587 VDD.n2187 VDD.n295 52.4337
R2588 VDD.n2183 VDD.n296 52.4337
R2589 VDD.n2179 VDD.n297 52.4337
R2590 VDD.n2149 VDD.n298 52.4337
R2591 VDD.n2172 VDD.n299 52.4337
R2592 VDD.n2169 VDD.n300 52.4337
R2593 VDD.n2165 VDD.n301 52.4337
R2594 VDD.n1479 VDD.n1146 52.4337
R2595 VDD.n1477 VDD.n1476 52.4337
R2596 VDD.n1472 VDD.n1153 52.4337
R2597 VDD.n1470 VDD.n1469 52.4337
R2598 VDD.n1161 VDD.n1160 52.4337
R2599 VDD.n1298 VDD.n1297 52.4337
R2600 VDD.n1295 VDD.n1294 52.4337
R2601 VDD.n1290 VDD.n1169 52.4337
R2602 VDD.n1288 VDD.n1287 52.4337
R2603 VDD.n1281 VDD.n1177 52.4337
R2604 VDD.n1279 VDD.n1278 52.4337
R2605 VDD.n1274 VDD.n1183 52.4337
R2606 VDD.n1272 VDD.n1271 52.4337
R2607 VDD.n1267 VDD.n1190 52.4337
R2608 VDD.n1265 VDD.n1264 52.4337
R2609 VDD.n1260 VDD.n1197 52.4337
R2610 VDD.n1258 VDD.n1257 52.4337
R2611 VDD.n1253 VDD.n1204 52.4337
R2612 VDD.n1251 VDD.n1250 52.4337
R2613 VDD.n1244 VDD.n1212 52.4337
R2614 VDD.n1242 VDD.n1241 52.4337
R2615 VDD.n1237 VDD.n1218 52.4337
R2616 VDD.n1235 VDD.n1234 52.4337
R2617 VDD.n1230 VDD.n1222 52.4337
R2618 VDD.n1228 VDD.n1227 52.4337
R2619 VDD.n1224 VDD.n630 52.4337
R2620 VDD.n642 VDD.n632 52.4337
R2621 VDD.n644 VDD.n635 52.4337
R2622 VDD.n645 VDD.n637 52.4337
R2623 VDD.n995 VDD.n994 52.4337
R2624 VDD.n819 VDD.n791 52.4337
R2625 VDD.n823 VDD.n792 52.4337
R2626 VDD.n825 VDD.n793 52.4337
R2627 VDD.n829 VDD.n794 52.4337
R2628 VDD.n831 VDD.n795 52.4337
R2629 VDD.n835 VDD.n796 52.4337
R2630 VDD.n837 VDD.n797 52.4337
R2631 VDD.n965 VDD.n798 52.4337
R2632 VDD.n842 VDD.n799 52.4337
R2633 VDD.n846 VDD.n800 52.4337
R2634 VDD.n848 VDD.n801 52.4337
R2635 VDD.n852 VDD.n802 52.4337
R2636 VDD.n854 VDD.n803 52.4337
R2637 VDD.n858 VDD.n804 52.4337
R2638 VDD.n860 VDD.n805 52.4337
R2639 VDD.n864 VDD.n806 52.4337
R2640 VDD.n866 VDD.n807 52.4337
R2641 VDD.n932 VDD.n808 52.4337
R2642 VDD.n871 VDD.n809 52.4337
R2643 VDD.n875 VDD.n810 52.4337
R2644 VDD.n877 VDD.n811 52.4337
R2645 VDD.n881 VDD.n812 52.4337
R2646 VDD.n883 VDD.n813 52.4337
R2647 VDD.n887 VDD.n814 52.4337
R2648 VDD.n889 VDD.n815 52.4337
R2649 VDD.n893 VDD.n816 52.4337
R2650 VDD.n895 VDD.n817 52.4337
R2651 VDD.n994 VDD.n790 52.4337
R2652 VDD.n822 VDD.n791 52.4337
R2653 VDD.n824 VDD.n792 52.4337
R2654 VDD.n828 VDD.n793 52.4337
R2655 VDD.n830 VDD.n794 52.4337
R2656 VDD.n834 VDD.n795 52.4337
R2657 VDD.n836 VDD.n796 52.4337
R2658 VDD.n840 VDD.n797 52.4337
R2659 VDD.n841 VDD.n798 52.4337
R2660 VDD.n845 VDD.n799 52.4337
R2661 VDD.n847 VDD.n800 52.4337
R2662 VDD.n851 VDD.n801 52.4337
R2663 VDD.n853 VDD.n802 52.4337
R2664 VDD.n857 VDD.n803 52.4337
R2665 VDD.n859 VDD.n804 52.4337
R2666 VDD.n863 VDD.n805 52.4337
R2667 VDD.n865 VDD.n806 52.4337
R2668 VDD.n869 VDD.n807 52.4337
R2669 VDD.n870 VDD.n808 52.4337
R2670 VDD.n874 VDD.n809 52.4337
R2671 VDD.n876 VDD.n810 52.4337
R2672 VDD.n880 VDD.n811 52.4337
R2673 VDD.n882 VDD.n812 52.4337
R2674 VDD.n886 VDD.n813 52.4337
R2675 VDD.n888 VDD.n814 52.4337
R2676 VDD.n892 VDD.n815 52.4337
R2677 VDD.n894 VDD.n816 52.4337
R2678 VDD.n898 VDD.n817 52.4337
R2679 VDD.n645 VDD.n636 52.4337
R2680 VDD.n644 VDD.n643 52.4337
R2681 VDD.n642 VDD.n631 52.4337
R2682 VDD.n1225 VDD.n1224 52.4337
R2683 VDD.n1229 VDD.n1228 52.4337
R2684 VDD.n1222 VDD.n1219 52.4337
R2685 VDD.n1236 VDD.n1235 52.4337
R2686 VDD.n1218 VDD.n1213 52.4337
R2687 VDD.n1243 VDD.n1242 52.4337
R2688 VDD.n1212 VDD.n1205 52.4337
R2689 VDD.n1252 VDD.n1251 52.4337
R2690 VDD.n1204 VDD.n1198 52.4337
R2691 VDD.n1259 VDD.n1258 52.4337
R2692 VDD.n1197 VDD.n1191 52.4337
R2693 VDD.n1266 VDD.n1265 52.4337
R2694 VDD.n1190 VDD.n1184 52.4337
R2695 VDD.n1273 VDD.n1272 52.4337
R2696 VDD.n1183 VDD.n1178 52.4337
R2697 VDD.n1280 VDD.n1279 52.4337
R2698 VDD.n1177 VDD.n1170 52.4337
R2699 VDD.n1289 VDD.n1288 52.4337
R2700 VDD.n1169 VDD.n1163 52.4337
R2701 VDD.n1296 VDD.n1295 52.4337
R2702 VDD.n1299 VDD.n1298 52.4337
R2703 VDD.n1160 VDD.n1154 52.4337
R2704 VDD.n1471 VDD.n1470 52.4337
R2705 VDD.n1153 VDD.n1147 52.4337
R2706 VDD.n1478 VDD.n1477 52.4337
R2707 VDD.n1146 VDD.n648 52.4337
R2708 VDD.n2274 VDD.n274 52.4337
R2709 VDD.n2268 VDD.n275 52.4337
R2710 VDD.n2264 VDD.n276 52.4337
R2711 VDD.n312 VDD.n277 52.4337
R2712 VDD.n315 VDD.n278 52.4337
R2713 VDD.n2254 VDD.n279 52.4337
R2714 VDD.n2250 VDD.n280 52.4337
R2715 VDD.n2246 VDD.n281 52.4337
R2716 VDD.n2236 VDD.n282 52.4337
R2717 VDD.n2234 VDD.n283 52.4337
R2718 VDD.n2230 VDD.n284 52.4337
R2719 VDD.n2226 VDD.n285 52.4337
R2720 VDD.n2222 VDD.n286 52.4337
R2721 VDD.n2218 VDD.n287 52.4337
R2722 VDD.n2214 VDD.n288 52.4337
R2723 VDD.n2210 VDD.n289 52.4337
R2724 VDD.n2206 VDD.n290 52.4337
R2725 VDD.n2202 VDD.n291 52.4337
R2726 VDD.n2194 VDD.n292 52.4337
R2727 VDD.n2192 VDD.n293 52.4337
R2728 VDD.n2188 VDD.n294 52.4337
R2729 VDD.n2184 VDD.n295 52.4337
R2730 VDD.n2180 VDD.n296 52.4337
R2731 VDD.n2148 VDD.n297 52.4337
R2732 VDD.n2151 VDD.n298 52.4337
R2733 VDD.n2170 VDD.n299 52.4337
R2734 VDD.n2166 VDD.n300 52.4337
R2735 VDD.n2162 VDD.n301 52.4337
R2736 VDD.n2384 VDD.n2383 52.4337
R2737 VDD.n198 VDD.n192 52.4337
R2738 VDD.n2391 VDD.n2390 52.4337
R2739 VDD.n191 VDD.n185 52.4337
R2740 VDD.n2398 VDD.n2397 52.4337
R2741 VDD.n184 VDD.n178 52.4337
R2742 VDD.n2405 VDD.n2404 52.4337
R2743 VDD.n177 VDD.n172 52.4337
R2744 VDD.n2412 VDD.n2411 52.4337
R2745 VDD.n171 VDD.n164 52.4337
R2746 VDD.n2421 VDD.n2420 52.4337
R2747 VDD.n163 VDD.n157 52.4337
R2748 VDD.n2428 VDD.n2427 52.4337
R2749 VDD.n156 VDD.n150 52.4337
R2750 VDD.n2435 VDD.n2434 52.4337
R2751 VDD.n149 VDD.n143 52.4337
R2752 VDD.n2442 VDD.n2441 52.4337
R2753 VDD.n142 VDD.n137 52.4337
R2754 VDD.n2449 VDD.n2448 52.4337
R2755 VDD.n136 VDD.n129 52.4337
R2756 VDD.n2458 VDD.n2457 52.4337
R2757 VDD.n128 VDD.n122 52.4337
R2758 VDD.n2465 VDD.n2464 52.4337
R2759 VDD.n121 VDD.n115 52.4337
R2760 VDD.n2472 VDD.n2471 52.4337
R2761 VDD.n114 VDD.n107 52.4337
R2762 VDD.n2479 VDD.n2478 52.4337
R2763 VDD.n2482 VDD.n2481 52.4337
R2764 VDD.n102 VDD.n99 52.4337
R2765 VDD.n2114 VDD.n2113 39.2114
R2766 VDD.n2109 VDD.n377 39.2114
R2767 VDD.n2107 VDD.n2106 39.2114
R2768 VDD.n2102 VDD.n380 39.2114
R2769 VDD.n2100 VDD.n2099 39.2114
R2770 VDD.n2096 VDD.n2095 39.2114
R2771 VDD.n2091 VDD.n383 39.2114
R2772 VDD.n2089 VDD.n2088 39.2114
R2773 VDD.n2084 VDD.n386 39.2114
R2774 VDD.n2082 VDD.n2081 39.2114
R2775 VDD.n2077 VDD.n2075 39.2114
R2776 VDD.n1946 VDD.n1945 39.2114
R2777 VDD.n1761 VDD.n1739 39.2114
R2778 VDD.n1938 VDD.n1740 39.2114
R2779 VDD.n1934 VDD.n1741 39.2114
R2780 VDD.n1930 VDD.n1742 39.2114
R2781 VDD.n1926 VDD.n1743 39.2114
R2782 VDD.n1922 VDD.n1744 39.2114
R2783 VDD.n1918 VDD.n1745 39.2114
R2784 VDD.n1914 VDD.n1746 39.2114
R2785 VDD.n1910 VDD.n1747 39.2114
R2786 VDD.n1905 VDD.n1748 39.2114
R2787 VDD.n1733 VDD.n505 39.2114
R2788 VDD.n1729 VDD.n504 39.2114
R2789 VDD.n1725 VDD.n503 39.2114
R2790 VDD.n1721 VDD.n502 39.2114
R2791 VDD.n1717 VDD.n501 39.2114
R2792 VDD.n1713 VDD.n500 39.2114
R2793 VDD.n1709 VDD.n499 39.2114
R2794 VDD.n1705 VDD.n498 39.2114
R2795 VDD.n1701 VDD.n497 39.2114
R2796 VDD.n1696 VDD.n496 39.2114
R2797 VDD.n1692 VDD.n495 39.2114
R2798 VDD.n1309 VDD.n612 39.2114
R2799 VDD.n1313 VDD.n1312 39.2114
R2800 VDD.n1318 VDD.n1317 39.2114
R2801 VDD.n1321 VDD.n1320 39.2114
R2802 VDD.n1326 VDD.n1325 39.2114
R2803 VDD.n1464 VDD.n1463 39.2114
R2804 VDD.n1461 VDD.n1328 39.2114
R2805 VDD.n1457 VDD.n1456 39.2114
R2806 VDD.n1450 VDD.n1330 39.2114
R2807 VDD.n1449 VDD.n1448 39.2114
R2808 VDD.n1442 VDD.n1332 39.2114
R2809 VDD.n2049 VDD.n2031 39.2114
R2810 VDD.n2047 VDD.n2046 39.2114
R2811 VDD.n2042 VDD.n2034 39.2114
R2812 VDD.n2040 VDD.n2039 39.2114
R2813 VDD.n2035 VDD.n353 39.2114
R2814 VDD.n2145 VDD.n2144 39.2114
R2815 VDD.n2142 VDD.n2141 39.2114
R2816 VDD.n2137 VDD.n358 39.2114
R2817 VDD.n2135 VDD.n2134 39.2114
R2818 VDD.n2129 VDD.n363 39.2114
R2819 VDD.n2127 VDD.n2126 39.2114
R2820 VDD.n1793 VDD.n1749 39.2114
R2821 VDD.n1797 VDD.n1750 39.2114
R2822 VDD.n1801 VDD.n1751 39.2114
R2823 VDD.n1805 VDD.n1752 39.2114
R2824 VDD.n1809 VDD.n1753 39.2114
R2825 VDD.n1813 VDD.n1754 39.2114
R2826 VDD.n1817 VDD.n1755 39.2114
R2827 VDD.n1821 VDD.n1756 39.2114
R2828 VDD.n1825 VDD.n1757 39.2114
R2829 VDD.n1829 VDD.n1758 39.2114
R2830 VDD.n1833 VDD.n1759 39.2114
R2831 VDD.n1796 VDD.n1749 39.2114
R2832 VDD.n1800 VDD.n1750 39.2114
R2833 VDD.n1804 VDD.n1751 39.2114
R2834 VDD.n1808 VDD.n1752 39.2114
R2835 VDD.n1812 VDD.n1753 39.2114
R2836 VDD.n1816 VDD.n1754 39.2114
R2837 VDD.n1820 VDD.n1755 39.2114
R2838 VDD.n1824 VDD.n1756 39.2114
R2839 VDD.n1828 VDD.n1757 39.2114
R2840 VDD.n1832 VDD.n1758 39.2114
R2841 VDD.n1835 VDD.n1759 39.2114
R2842 VDD.n2128 VDD.n2127 39.2114
R2843 VDD.n363 VDD.n359 39.2114
R2844 VDD.n2136 VDD.n2135 39.2114
R2845 VDD.n358 VDD.n356 39.2114
R2846 VDD.n2143 VDD.n2142 39.2114
R2847 VDD.n2146 VDD.n2145 39.2114
R2848 VDD.n2036 VDD.n2035 39.2114
R2849 VDD.n2041 VDD.n2040 39.2114
R2850 VDD.n2034 VDD.n2032 39.2114
R2851 VDD.n2048 VDD.n2047 39.2114
R2852 VDD.n2031 VDD.n2029 39.2114
R2853 VDD.n1310 VDD.n1309 39.2114
R2854 VDD.n1312 VDD.n1306 39.2114
R2855 VDD.n1319 VDD.n1318 39.2114
R2856 VDD.n1320 VDD.n1304 39.2114
R2857 VDD.n1327 VDD.n1326 39.2114
R2858 VDD.n1463 VDD.n1462 39.2114
R2859 VDD.n1458 VDD.n1328 39.2114
R2860 VDD.n1456 VDD.n1455 39.2114
R2861 VDD.n1451 VDD.n1450 39.2114
R2862 VDD.n1448 VDD.n1447 39.2114
R2863 VDD.n1443 VDD.n1442 39.2114
R2864 VDD.n1695 VDD.n495 39.2114
R2865 VDD.n1700 VDD.n496 39.2114
R2866 VDD.n1704 VDD.n497 39.2114
R2867 VDD.n1708 VDD.n498 39.2114
R2868 VDD.n1712 VDD.n499 39.2114
R2869 VDD.n1716 VDD.n500 39.2114
R2870 VDD.n1720 VDD.n501 39.2114
R2871 VDD.n1724 VDD.n502 39.2114
R2872 VDD.n1728 VDD.n503 39.2114
R2873 VDD.n1732 VDD.n504 39.2114
R2874 VDD.n507 VDD.n505 39.2114
R2875 VDD.n1945 VDD.n481 39.2114
R2876 VDD.n1939 VDD.n1739 39.2114
R2877 VDD.n1935 VDD.n1740 39.2114
R2878 VDD.n1931 VDD.n1741 39.2114
R2879 VDD.n1927 VDD.n1742 39.2114
R2880 VDD.n1923 VDD.n1743 39.2114
R2881 VDD.n1919 VDD.n1744 39.2114
R2882 VDD.n1915 VDD.n1745 39.2114
R2883 VDD.n1911 VDD.n1746 39.2114
R2884 VDD.n1906 VDD.n1747 39.2114
R2885 VDD.n1902 VDD.n1748 39.2114
R2886 VDD.n2075 VDD.n387 39.2114
R2887 VDD.n2083 VDD.n2082 39.2114
R2888 VDD.n386 VDD.n384 39.2114
R2889 VDD.n2090 VDD.n2089 39.2114
R2890 VDD.n383 VDD.n381 39.2114
R2891 VDD.n2097 VDD.n2096 39.2114
R2892 VDD.n2101 VDD.n2100 39.2114
R2893 VDD.n380 VDD.n378 39.2114
R2894 VDD.n2108 VDD.n2107 39.2114
R2895 VDD.n377 VDD.n375 39.2114
R2896 VDD.n2115 VDD.n2114 39.2114
R2897 VDD.n1676 VDD.n483 39.2114
R2898 VDD.n1672 VDD.n484 39.2114
R2899 VDD.n1668 VDD.n485 39.2114
R2900 VDD.n1664 VDD.n486 39.2114
R2901 VDD.n1660 VDD.n487 39.2114
R2902 VDD.n1656 VDD.n488 39.2114
R2903 VDD.n1652 VDD.n489 39.2114
R2904 VDD.n1648 VDD.n490 39.2114
R2905 VDD.n1644 VDD.n491 39.2114
R2906 VDD.n1640 VDD.n492 39.2114
R2907 VDD.n1636 VDD.n493 39.2114
R2908 VDD.n1525 VDD.n616 39.2114
R2909 VDD.n1524 VDD.n1523 39.2114
R2910 VDD.n1517 VDD.n619 39.2114
R2911 VDD.n1516 VDD.n1515 39.2114
R2912 VDD.n1509 VDD.n621 39.2114
R2913 VDD.n1508 VDD.n1507 39.2114
R2914 VDD.n1353 VDD.n623 39.2114
R2915 VDD.n1356 VDD.n1355 39.2114
R2916 VDD.n1361 VDD.n1360 39.2114
R2917 VDD.n1364 VDD.n1363 39.2114
R2918 VDD.n1370 VDD.n1369 39.2114
R2919 VDD.n1633 VDD.n493 39.2114
R2920 VDD.n1637 VDD.n492 39.2114
R2921 VDD.n1641 VDD.n491 39.2114
R2922 VDD.n1645 VDD.n490 39.2114
R2923 VDD.n1649 VDD.n489 39.2114
R2924 VDD.n1653 VDD.n488 39.2114
R2925 VDD.n1657 VDD.n487 39.2114
R2926 VDD.n1661 VDD.n486 39.2114
R2927 VDD.n1665 VDD.n485 39.2114
R2928 VDD.n1669 VDD.n484 39.2114
R2929 VDD.n1673 VDD.n483 39.2114
R2930 VDD.n1526 VDD.n1525 39.2114
R2931 VDD.n1523 VDD.n1522 39.2114
R2932 VDD.n1518 VDD.n1517 39.2114
R2933 VDD.n1515 VDD.n1514 39.2114
R2934 VDD.n1510 VDD.n1509 39.2114
R2935 VDD.n1507 VDD.n1506 39.2114
R2936 VDD.n1354 VDD.n1353 39.2114
R2937 VDD.n1355 VDD.n1351 39.2114
R2938 VDD.n1362 VDD.n1361 39.2114
R2939 VDD.n1363 VDD.n1347 39.2114
R2940 VDD.n1371 VDD.n1370 39.2114
R2941 VDD.n902 VDD.n901 37.4308
R2942 VDD.n935 VDD.n934 37.4308
R2943 VDD.n968 VDD.n967 37.4308
R2944 VDD.n1494 VDD.n1493 37.4308
R2945 VDD.n1249 VDD.n1208 37.4308
R2946 VDD.n1286 VDD.n1173 37.4308
R2947 VDD.n201 VDD.n200 37.4308
R2948 VDD.n2418 VDD.n167 37.4308
R2949 VDD.n2455 VDD.n132 37.4308
R2950 VDD.n2200 VDD.n341 37.4308
R2951 VDD.n2244 VDD.n2243 37.4308
R2952 VDD.n2161 VDD.n2160 37.4308
R2953 VDD.n1736 VDD.n508 32.6249
R2954 VDD.n1693 VDD.n511 32.6249
R2955 VDD.n1444 VDD.n1441 32.6249
R2956 VDD.n1534 VDD.n611 32.6249
R2957 VDD.n1903 VDD.n1900 32.6249
R2958 VDD.n2078 VDD.n2074 32.6249
R2959 VDD.n1948 VDD.n1947 32.6249
R2960 VDD.n2118 VDD.n2117 32.6249
R2961 VDD.n2125 VDD.n2124 32.6249
R2962 VDD.n1839 VDD.n1837 32.6249
R2963 VDD.n1794 VDD.n474 32.6249
R2964 VDD.n1678 VDD.n1675 32.6249
R2965 VDD.n1632 VDD.n1631 32.6249
R2966 VDD.n1374 VDD.n1373 32.6249
R2967 VDD.n1367 VDD.n1349 30.449
R2968 VDD.n527 VDD.n526 30.449
R2969 VDD.n1335 VDD.n1334 30.449
R2970 VDD.n1698 VDD.n510 30.449
R2971 VDD.n1792 VDD.n1791 30.449
R2972 VDD.n390 VDD.n389 30.449
R2973 VDD.n1908 VDD.n1763 30.449
R2974 VDD.n2131 VDD.n361 30.449
R2975 VDD.n1349 VDD.n1348 25.7944
R2976 VDD.n526 VDD.n525 25.7944
R2977 VDD.n901 VDD.n900 25.7944
R2978 VDD.n934 VDD.n933 25.7944
R2979 VDD.n967 VDD.n966 25.7944
R2980 VDD.n1493 VDD.n1492 25.7944
R2981 VDD.n1208 VDD.n1207 25.7944
R2982 VDD.n1173 VDD.n1172 25.7944
R2983 VDD.n1334 VDD.n1333 25.7944
R2984 VDD.n510 VDD.n509 25.7944
R2985 VDD.n1791 VDD.n1790 25.7944
R2986 VDD.n200 VDD.n199 25.7944
R2987 VDD.n167 VDD.n166 25.7944
R2988 VDD.n132 VDD.n131 25.7944
R2989 VDD.n341 VDD.n340 25.7944
R2990 VDD.n2243 VDD.n2242 25.7944
R2991 VDD.n389 VDD.n388 25.7944
R2992 VDD.n1763 VDD.n1762 25.7944
R2993 VDD.n2160 VDD.n2159 25.7944
R2994 VDD.n361 VDD.n360 25.7944
R2995 VDD.n993 VDD.n785 23.437
R2996 VDD.n1486 VDD.n646 23.437
R2997 VDD.n2273 VDD.n269 23.437
R2998 VDD.n2490 VDD.n98 23.437
R2999 VDD.n2055 VDD.n2028 19.6688
R3000 VDD.n1530 VDD.n1529 19.6688
R3001 VDD.n1004 VDD.n783 19.3944
R3002 VDD.n1004 VDD.n781 19.3944
R3003 VDD.n1008 VDD.n781 19.3944
R3004 VDD.n1008 VDD.n770 19.3944
R3005 VDD.n1020 VDD.n770 19.3944
R3006 VDD.n1020 VDD.n768 19.3944
R3007 VDD.n1024 VDD.n768 19.3944
R3008 VDD.n1024 VDD.n759 19.3944
R3009 VDD.n1036 VDD.n759 19.3944
R3010 VDD.n1036 VDD.n757 19.3944
R3011 VDD.n1040 VDD.n757 19.3944
R3012 VDD.n1040 VDD.n746 19.3944
R3013 VDD.n1052 VDD.n746 19.3944
R3014 VDD.n1052 VDD.n744 19.3944
R3015 VDD.n1056 VDD.n744 19.3944
R3016 VDD.n1056 VDD.n735 19.3944
R3017 VDD.n1069 VDD.n735 19.3944
R3018 VDD.n1069 VDD.n733 19.3944
R3019 VDD.n1073 VDD.n733 19.3944
R3020 VDD.n1073 VDD.n692 19.3944
R3021 VDD.n1085 VDD.n692 19.3944
R3022 VDD.n1085 VDD.n690 19.3944
R3023 VDD.n1089 VDD.n690 19.3944
R3024 VDD.n1089 VDD.n681 19.3944
R3025 VDD.n1101 VDD.n681 19.3944
R3026 VDD.n1101 VDD.n679 19.3944
R3027 VDD.n1105 VDD.n679 19.3944
R3028 VDD.n1105 VDD.n668 19.3944
R3029 VDD.n1117 VDD.n668 19.3944
R3030 VDD.n1117 VDD.n666 19.3944
R3031 VDD.n1121 VDD.n666 19.3944
R3032 VDD.n1121 VDD.n657 19.3944
R3033 VDD.n1133 VDD.n657 19.3944
R3034 VDD.n1133 VDD.n655 19.3944
R3035 VDD.n1137 VDD.n655 19.3944
R3036 VDD.n1137 VDD.n639 19.3944
R3037 VDD.n1488 VDD.n639 19.3944
R3038 VDD.n931 VDD.n872 19.3944
R3039 VDD.n927 VDD.n872 19.3944
R3040 VDD.n927 VDD.n926 19.3944
R3041 VDD.n926 VDD.n925 19.3944
R3042 VDD.n925 VDD.n878 19.3944
R3043 VDD.n921 VDD.n878 19.3944
R3044 VDD.n921 VDD.n920 19.3944
R3045 VDD.n920 VDD.n919 19.3944
R3046 VDD.n919 VDD.n884 19.3944
R3047 VDD.n915 VDD.n884 19.3944
R3048 VDD.n915 VDD.n914 19.3944
R3049 VDD.n914 VDD.n913 19.3944
R3050 VDD.n913 VDD.n890 19.3944
R3051 VDD.n909 VDD.n890 19.3944
R3052 VDD.n909 VDD.n908 19.3944
R3053 VDD.n908 VDD.n907 19.3944
R3054 VDD.n907 VDD.n896 19.3944
R3055 VDD.n903 VDD.n896 19.3944
R3056 VDD.n964 VDD.n843 19.3944
R3057 VDD.n960 VDD.n843 19.3944
R3058 VDD.n960 VDD.n959 19.3944
R3059 VDD.n959 VDD.n958 19.3944
R3060 VDD.n958 VDD.n849 19.3944
R3061 VDD.n954 VDD.n849 19.3944
R3062 VDD.n954 VDD.n953 19.3944
R3063 VDD.n953 VDD.n952 19.3944
R3064 VDD.n952 VDD.n855 19.3944
R3065 VDD.n948 VDD.n855 19.3944
R3066 VDD.n948 VDD.n947 19.3944
R3067 VDD.n947 VDD.n946 19.3944
R3068 VDD.n946 VDD.n861 19.3944
R3069 VDD.n942 VDD.n861 19.3944
R3070 VDD.n942 VDD.n941 19.3944
R3071 VDD.n941 VDD.n940 19.3944
R3072 VDD.n940 VDD.n867 19.3944
R3073 VDD.n936 VDD.n867 19.3944
R3074 VDD.n996 VDD.n789 19.3944
R3075 VDD.n991 VDD.n789 19.3944
R3076 VDD.n991 VDD.n820 19.3944
R3077 VDD.n987 VDD.n820 19.3944
R3078 VDD.n987 VDD.n986 19.3944
R3079 VDD.n986 VDD.n985 19.3944
R3080 VDD.n985 VDD.n826 19.3944
R3081 VDD.n981 VDD.n826 19.3944
R3082 VDD.n981 VDD.n980 19.3944
R3083 VDD.n980 VDD.n979 19.3944
R3084 VDD.n979 VDD.n832 19.3944
R3085 VDD.n975 VDD.n832 19.3944
R3086 VDD.n975 VDD.n974 19.3944
R3087 VDD.n974 VDD.n973 19.3944
R3088 VDD.n973 VDD.n838 19.3944
R3089 VDD.n969 VDD.n838 19.3944
R3090 VDD.n1000 VDD.n787 19.3944
R3091 VDD.n1000 VDD.n777 19.3944
R3092 VDD.n1012 VDD.n777 19.3944
R3093 VDD.n1012 VDD.n775 19.3944
R3094 VDD.n1016 VDD.n775 19.3944
R3095 VDD.n1016 VDD.n765 19.3944
R3096 VDD.n1028 VDD.n765 19.3944
R3097 VDD.n1028 VDD.n763 19.3944
R3098 VDD.n1032 VDD.n763 19.3944
R3099 VDD.n1032 VDD.n753 19.3944
R3100 VDD.n1044 VDD.n753 19.3944
R3101 VDD.n1044 VDD.n751 19.3944
R3102 VDD.n1048 VDD.n751 19.3944
R3103 VDD.n1048 VDD.n741 19.3944
R3104 VDD.n1060 VDD.n741 19.3944
R3105 VDD.n1060 VDD.n739 19.3944
R3106 VDD.n1065 VDD.n739 19.3944
R3107 VDD.n1065 VDD.n729 19.3944
R3108 VDD.n1077 VDD.n729 19.3944
R3109 VDD.n1077 VDD.n697 19.3944
R3110 VDD.n1081 VDD.n697 19.3944
R3111 VDD.n1081 VDD.n687 19.3944
R3112 VDD.n1093 VDD.n687 19.3944
R3113 VDD.n1093 VDD.n685 19.3944
R3114 VDD.n1097 VDD.n685 19.3944
R3115 VDD.n1097 VDD.n675 19.3944
R3116 VDD.n1109 VDD.n675 19.3944
R3117 VDD.n1109 VDD.n673 19.3944
R3118 VDD.n1113 VDD.n673 19.3944
R3119 VDD.n1113 VDD.n663 19.3944
R3120 VDD.n1125 VDD.n663 19.3944
R3121 VDD.n1125 VDD.n661 19.3944
R3122 VDD.n1129 VDD.n661 19.3944
R3123 VDD.n1129 VDD.n651 19.3944
R3124 VDD.n1141 VDD.n651 19.3944
R3125 VDD.n1141 VDD.n649 19.3944
R3126 VDD.n1484 VDD.n649 19.3944
R3127 VDD.n1245 VDD.n1206 19.3944
R3128 VDD.n1245 VDD.n1211 19.3944
R3129 VDD.n1240 VDD.n1211 19.3944
R3130 VDD.n1240 VDD.n1239 19.3944
R3131 VDD.n1239 VDD.n1238 19.3944
R3132 VDD.n1238 VDD.n1217 19.3944
R3133 VDD.n1233 VDD.n1217 19.3944
R3134 VDD.n1233 VDD.n1232 19.3944
R3135 VDD.n1232 VDD.n1231 19.3944
R3136 VDD.n1226 VDD.n1223 19.3944
R3137 VDD.n1502 VDD.n629 19.3944
R3138 VDD.n1502 VDD.n1501 19.3944
R3139 VDD.n1501 VDD.n1500 19.3944
R3140 VDD.n1500 VDD.n633 19.3944
R3141 VDD.n1496 VDD.n633 19.3944
R3142 VDD.n1496 VDD.n1495 19.3944
R3143 VDD.n1282 VDD.n1171 19.3944
R3144 VDD.n1282 VDD.n1176 19.3944
R3145 VDD.n1277 VDD.n1176 19.3944
R3146 VDD.n1277 VDD.n1276 19.3944
R3147 VDD.n1276 VDD.n1275 19.3944
R3148 VDD.n1275 VDD.n1182 19.3944
R3149 VDD.n1270 VDD.n1182 19.3944
R3150 VDD.n1270 VDD.n1269 19.3944
R3151 VDD.n1269 VDD.n1268 19.3944
R3152 VDD.n1268 VDD.n1189 19.3944
R3153 VDD.n1263 VDD.n1189 19.3944
R3154 VDD.n1263 VDD.n1262 19.3944
R3155 VDD.n1262 VDD.n1261 19.3944
R3156 VDD.n1261 VDD.n1196 19.3944
R3157 VDD.n1256 VDD.n1196 19.3944
R3158 VDD.n1256 VDD.n1255 19.3944
R3159 VDD.n1255 VDD.n1254 19.3944
R3160 VDD.n1254 VDD.n1203 19.3944
R3161 VDD.n1481 VDD.n1480 19.3944
R3162 VDD.n1480 VDD.n1145 19.3944
R3163 VDD.n1475 VDD.n1145 19.3944
R3164 VDD.n1475 VDD.n1474 19.3944
R3165 VDD.n1474 VDD.n1473 19.3944
R3166 VDD.n1473 VDD.n1152 19.3944
R3167 VDD.n1468 VDD.n1152 19.3944
R3168 VDD.n1158 VDD.n1155 19.3944
R3169 VDD.n1300 VDD.n1159 19.3944
R3170 VDD.n1162 VDD.n1159 19.3944
R3171 VDD.n1293 VDD.n1162 19.3944
R3172 VDD.n1293 VDD.n1292 19.3944
R3173 VDD.n1292 VDD.n1291 19.3944
R3174 VDD.n1291 VDD.n1168 19.3944
R3175 VDD.n2284 VDD.n267 19.3944
R3176 VDD.n2284 VDD.n265 19.3944
R3177 VDD.n2288 VDD.n265 19.3944
R3178 VDD.n2288 VDD.n254 19.3944
R3179 VDD.n2300 VDD.n254 19.3944
R3180 VDD.n2300 VDD.n252 19.3944
R3181 VDD.n2304 VDD.n252 19.3944
R3182 VDD.n2304 VDD.n243 19.3944
R3183 VDD.n2316 VDD.n243 19.3944
R3184 VDD.n2316 VDD.n241 19.3944
R3185 VDD.n2320 VDD.n241 19.3944
R3186 VDD.n2320 VDD.n230 19.3944
R3187 VDD.n2332 VDD.n230 19.3944
R3188 VDD.n2332 VDD.n228 19.3944
R3189 VDD.n2336 VDD.n228 19.3944
R3190 VDD.n2336 VDD.n218 19.3944
R3191 VDD.n2348 VDD.n218 19.3944
R3192 VDD.n2348 VDD.n216 19.3944
R3193 VDD.n2352 VDD.n216 19.3944
R3194 VDD.n2353 VDD.n2352 19.3944
R3195 VDD.n2354 VDD.n2353 19.3944
R3196 VDD.n2354 VDD.n214 19.3944
R3197 VDD.n2358 VDD.n214 19.3944
R3198 VDD.n2359 VDD.n2358 19.3944
R3199 VDD.n2360 VDD.n2359 19.3944
R3200 VDD.n2360 VDD.n211 19.3944
R3201 VDD.n2364 VDD.n211 19.3944
R3202 VDD.n2365 VDD.n2364 19.3944
R3203 VDD.n2366 VDD.n2365 19.3944
R3204 VDD.n2366 VDD.n208 19.3944
R3205 VDD.n2370 VDD.n208 19.3944
R3206 VDD.n2371 VDD.n2370 19.3944
R3207 VDD.n2372 VDD.n2371 19.3944
R3208 VDD.n2372 VDD.n205 19.3944
R3209 VDD.n2376 VDD.n205 19.3944
R3210 VDD.n2377 VDD.n2376 19.3944
R3211 VDD.n2378 VDD.n2377 19.3944
R3212 VDD.n2414 VDD.n165 19.3944
R3213 VDD.n2414 VDD.n170 19.3944
R3214 VDD.n2409 VDD.n170 19.3944
R3215 VDD.n2409 VDD.n2408 19.3944
R3216 VDD.n2408 VDD.n2407 19.3944
R3217 VDD.n2407 VDD.n176 19.3944
R3218 VDD.n2402 VDD.n176 19.3944
R3219 VDD.n2402 VDD.n2401 19.3944
R3220 VDD.n2401 VDD.n2400 19.3944
R3221 VDD.n2400 VDD.n183 19.3944
R3222 VDD.n2395 VDD.n183 19.3944
R3223 VDD.n2395 VDD.n2394 19.3944
R3224 VDD.n2394 VDD.n2393 19.3944
R3225 VDD.n2393 VDD.n190 19.3944
R3226 VDD.n2388 VDD.n190 19.3944
R3227 VDD.n2388 VDD.n2387 19.3944
R3228 VDD.n2387 VDD.n2386 19.3944
R3229 VDD.n2386 VDD.n197 19.3944
R3230 VDD.n2451 VDD.n130 19.3944
R3231 VDD.n2451 VDD.n135 19.3944
R3232 VDD.n2446 VDD.n135 19.3944
R3233 VDD.n2446 VDD.n2445 19.3944
R3234 VDD.n2445 VDD.n2444 19.3944
R3235 VDD.n2444 VDD.n141 19.3944
R3236 VDD.n2439 VDD.n141 19.3944
R3237 VDD.n2439 VDD.n2438 19.3944
R3238 VDD.n2438 VDD.n2437 19.3944
R3239 VDD.n2437 VDD.n148 19.3944
R3240 VDD.n2432 VDD.n148 19.3944
R3241 VDD.n2432 VDD.n2431 19.3944
R3242 VDD.n2431 VDD.n2430 19.3944
R3243 VDD.n2430 VDD.n155 19.3944
R3244 VDD.n2425 VDD.n155 19.3944
R3245 VDD.n2425 VDD.n2424 19.3944
R3246 VDD.n2424 VDD.n2423 19.3944
R3247 VDD.n2423 VDD.n162 19.3944
R3248 VDD.n2485 VDD.n2484 19.3944
R3249 VDD.n2484 VDD.n2483 19.3944
R3250 VDD.n2483 VDD.n105 19.3944
R3251 VDD.n106 VDD.n105 19.3944
R3252 VDD.n2476 VDD.n106 19.3944
R3253 VDD.n2476 VDD.n2475 19.3944
R3254 VDD.n2475 VDD.n2474 19.3944
R3255 VDD.n2474 VDD.n113 19.3944
R3256 VDD.n2469 VDD.n113 19.3944
R3257 VDD.n2469 VDD.n2468 19.3944
R3258 VDD.n2468 VDD.n2467 19.3944
R3259 VDD.n2467 VDD.n120 19.3944
R3260 VDD.n2462 VDD.n120 19.3944
R3261 VDD.n2462 VDD.n2461 19.3944
R3262 VDD.n2461 VDD.n2460 19.3944
R3263 VDD.n2460 VDD.n127 19.3944
R3264 VDD.n2280 VDD.n271 19.3944
R3265 VDD.n2280 VDD.n261 19.3944
R3266 VDD.n2292 VDD.n261 19.3944
R3267 VDD.n2292 VDD.n259 19.3944
R3268 VDD.n2296 VDD.n259 19.3944
R3269 VDD.n2296 VDD.n249 19.3944
R3270 VDD.n2308 VDD.n249 19.3944
R3271 VDD.n2308 VDD.n247 19.3944
R3272 VDD.n2312 VDD.n247 19.3944
R3273 VDD.n2312 VDD.n237 19.3944
R3274 VDD.n2324 VDD.n237 19.3944
R3275 VDD.n2324 VDD.n235 19.3944
R3276 VDD.n2328 VDD.n235 19.3944
R3277 VDD.n2328 VDD.n225 19.3944
R3278 VDD.n2340 VDD.n225 19.3944
R3279 VDD.n2340 VDD.n223 19.3944
R3280 VDD.n2344 VDD.n223 19.3944
R3281 VDD.n2344 VDD.n47 19.3944
R3282 VDD.n2526 VDD.n47 19.3944
R3283 VDD.n2526 VDD.n48 19.3944
R3284 VDD.n2520 VDD.n48 19.3944
R3285 VDD.n2520 VDD.n2519 19.3944
R3286 VDD.n2519 VDD.n2518 19.3944
R3287 VDD.n2518 VDD.n60 19.3944
R3288 VDD.n2512 VDD.n60 19.3944
R3289 VDD.n2512 VDD.n2511 19.3944
R3290 VDD.n2511 VDD.n2510 19.3944
R3291 VDD.n2510 VDD.n70 19.3944
R3292 VDD.n2504 VDD.n70 19.3944
R3293 VDD.n2504 VDD.n2503 19.3944
R3294 VDD.n2503 VDD.n2502 19.3944
R3295 VDD.n2502 VDD.n82 19.3944
R3296 VDD.n2496 VDD.n82 19.3944
R3297 VDD.n2496 VDD.n2495 19.3944
R3298 VDD.n2495 VDD.n2494 19.3944
R3299 VDD.n2494 VDD.n93 19.3944
R3300 VDD.n2488 VDD.n93 19.3944
R3301 VDD.n2238 VDD.n321 19.3944
R3302 VDD.n2238 VDD.n2235 19.3944
R3303 VDD.n2235 VDD.n2232 19.3944
R3304 VDD.n2232 VDD.n2231 19.3944
R3305 VDD.n2231 VDD.n2228 19.3944
R3306 VDD.n2228 VDD.n2227 19.3944
R3307 VDD.n2227 VDD.n2224 19.3944
R3308 VDD.n2224 VDD.n2223 19.3944
R3309 VDD.n2223 VDD.n2220 19.3944
R3310 VDD.n2220 VDD.n2219 19.3944
R3311 VDD.n2219 VDD.n2216 19.3944
R3312 VDD.n2216 VDD.n2215 19.3944
R3313 VDD.n2215 VDD.n2212 19.3944
R3314 VDD.n2212 VDD.n2211 19.3944
R3315 VDD.n2211 VDD.n2208 19.3944
R3316 VDD.n2208 VDD.n2207 19.3944
R3317 VDD.n2207 VDD.n2204 19.3944
R3318 VDD.n2204 VDD.n2203 19.3944
R3319 VDD.n2276 VDD.n273 19.3944
R3320 VDD.n2271 VDD.n273 19.3944
R3321 VDD.n2271 VDD.n2270 19.3944
R3322 VDD.n2270 VDD.n2269 19.3944
R3323 VDD.n2269 VDD.n2266 19.3944
R3324 VDD.n2266 VDD.n2265 19.3944
R3325 VDD.n2265 VDD.n2262 19.3944
R3326 VDD.n314 VDD.n309 19.3944
R3327 VDD.n2258 VDD.n2257 19.3944
R3328 VDD.n2257 VDD.n2255 19.3944
R3329 VDD.n2255 VDD.n2252 19.3944
R3330 VDD.n2252 VDD.n2251 19.3944
R3331 VDD.n2251 VDD.n2248 19.3944
R3332 VDD.n2248 VDD.n2247 19.3944
R3333 VDD.n2196 VDD.n339 19.3944
R3334 VDD.n2196 VDD.n2193 19.3944
R3335 VDD.n2193 VDD.n2190 19.3944
R3336 VDD.n2190 VDD.n2189 19.3944
R3337 VDD.n2189 VDD.n2186 19.3944
R3338 VDD.n2186 VDD.n2185 19.3944
R3339 VDD.n2185 VDD.n2182 19.3944
R3340 VDD.n2182 VDD.n2181 19.3944
R3341 VDD.n2181 VDD.n2178 19.3944
R3342 VDD.n2150 VDD.n349 19.3944
R3343 VDD.n2174 VDD.n2173 19.3944
R3344 VDD.n2173 VDD.n2171 19.3944
R3345 VDD.n2171 VDD.n2168 19.3944
R3346 VDD.n2168 VDD.n2167 19.3944
R3347 VDD.n2167 VDD.n2164 19.3944
R3348 VDD.n2164 VDD.n2163 19.3944
R3349 VDD.n935 VDD.n931 19.0066
R3350 VDD.n1249 VDD.n1206 19.0066
R3351 VDD.n2418 VDD.n165 19.0066
R3352 VDD.n2200 VDD.n339 19.0066
R3353 VDD.n1532 VDD.n613 18.8094
R3354 VDD.n1738 VDD.n482 18.8094
R3355 VDD.n1944 VDD.n476 18.8094
R3356 VDD.n369 VDD.n354 18.8094
R3357 VDD.n1002 VDD.n785 14.9282
R3358 VDD.n1010 VDD.n779 14.9282
R3359 VDD.n1010 VDD.n772 14.9282
R3360 VDD.n1018 VDD.n772 14.9282
R3361 VDD.n1018 VDD.n773 14.9282
R3362 VDD.n1026 VDD.n761 14.9282
R3363 VDD.n1034 VDD.n761 14.9282
R3364 VDD.n1042 VDD.n755 14.9282
R3365 VDD.n1050 VDD.n748 14.9282
R3366 VDD.n1050 VDD.n749 14.9282
R3367 VDD.n1058 VDD.n737 14.9282
R3368 VDD.n1067 VDD.n737 14.9282
R3369 VDD.n1075 VDD.n731 14.9282
R3370 VDD.n1083 VDD.n694 14.9282
R3371 VDD.n1083 VDD.n695 14.9282
R3372 VDD.n1091 VDD.n683 14.9282
R3373 VDD.n1099 VDD.n683 14.9282
R3374 VDD.n1107 VDD.n677 14.9282
R3375 VDD.n1115 VDD.n670 14.9282
R3376 VDD.n1115 VDD.n671 14.9282
R3377 VDD.n1123 VDD.n659 14.9282
R3378 VDD.n1131 VDD.n659 14.9282
R3379 VDD.n1131 VDD.n653 14.9282
R3380 VDD.n1139 VDD.n653 14.9282
R3381 VDD.n1486 VDD.n641 14.9282
R3382 VDD.n2282 VDD.n269 14.9282
R3383 VDD.n2290 VDD.n263 14.9282
R3384 VDD.n2290 VDD.n256 14.9282
R3385 VDD.n2298 VDD.n256 14.9282
R3386 VDD.n2298 VDD.n257 14.9282
R3387 VDD.n2306 VDD.n245 14.9282
R3388 VDD.n2314 VDD.n245 14.9282
R3389 VDD.n2322 VDD.n239 14.9282
R3390 VDD.n2330 VDD.n232 14.9282
R3391 VDD.n2330 VDD.n233 14.9282
R3392 VDD.n2338 VDD.n221 14.9282
R3393 VDD.n2346 VDD.n221 14.9282
R3394 VDD.n2524 VDD.n51 14.9282
R3395 VDD.n2523 VDD.n2522 14.9282
R3396 VDD.n2522 VDD.n55 14.9282
R3397 VDD.n2516 VDD.n2515 14.9282
R3398 VDD.n2515 VDD.n2514 14.9282
R3399 VDD.n2508 VDD.n72 14.9282
R3400 VDD.n2507 VDD.n2506 14.9282
R3401 VDD.n2506 VDD.n76 14.9282
R3402 VDD.n2500 VDD.n2499 14.9282
R3403 VDD.n2499 VDD.n2498 14.9282
R3404 VDD.n2498 VDD.n87 14.9282
R3405 VDD.n2492 VDD.n87 14.9282
R3406 VDD.n2491 VDD.n2490 14.9282
R3407 VDD.n968 VDD.n964 12.9944
R3408 VDD.n969 VDD.n968 12.9944
R3409 VDD.n1286 VDD.n1171 12.9944
R3410 VDD.n1286 VDD.n1168 12.9944
R3411 VDD.n2455 VDD.n130 12.9944
R3412 VDD.n2455 VDD.n127 12.9944
R3413 VDD.n2244 VDD.n321 12.9944
R3414 VDD.n2247 VDD.n2244 12.9944
R3415 VDD.n2052 VDD.n2028 12.9566
R3416 VDD.n1529 VDD.n1528 12.9566
R3417 VDD.n1042 VDD.t145 12.6891
R3418 VDD.t140 VDD.n677 12.6891
R3419 VDD.n2322 VDD.t116 12.6891
R3420 VDD.n72 VDD.t119 12.6891
R3421 VDD.t108 VDD.n731 12.3905
R3422 VDD.n1075 VDD.t124 12.3905
R3423 VDD.t142 VDD.n51 12.3905
R3424 VDD.n2524 VDD.t131 12.3905
R3425 VDD.t135 VDD.n755 12.092
R3426 VDD.n1107 VDD.t147 12.092
R3427 VDD.t122 VDD.n239 12.092
R3428 VDD.n2508 VDD.t152 12.092
R3429 VDD.n1736 VDD.n1735 10.6151
R3430 VDD.n1735 VDD.n1734 10.6151
R3431 VDD.n1734 VDD.n1731 10.6151
R3432 VDD.n1731 VDD.n1730 10.6151
R3433 VDD.n1730 VDD.n1727 10.6151
R3434 VDD.n1727 VDD.n1726 10.6151
R3435 VDD.n1726 VDD.n1723 10.6151
R3436 VDD.n1723 VDD.n1722 10.6151
R3437 VDD.n1722 VDD.n1719 10.6151
R3438 VDD.n1719 VDD.n1718 10.6151
R3439 VDD.n1718 VDD.n1715 10.6151
R3440 VDD.n1715 VDD.n1714 10.6151
R3441 VDD.n1714 VDD.n1711 10.6151
R3442 VDD.n1711 VDD.n1710 10.6151
R3443 VDD.n1710 VDD.n1707 10.6151
R3444 VDD.n1707 VDD.n1706 10.6151
R3445 VDD.n1706 VDD.n1703 10.6151
R3446 VDD.n1703 VDD.n1702 10.6151
R3447 VDD.n1702 VDD.n1699 10.6151
R3448 VDD.n1697 VDD.n1694 10.6151
R3449 VDD.n1694 VDD.n1693 10.6151
R3450 VDD.n1441 VDD.n1440 10.6151
R3451 VDD.n1440 VDD.n1438 10.6151
R3452 VDD.n1438 VDD.n1437 10.6151
R3453 VDD.n1437 VDD.n1435 10.6151
R3454 VDD.n1435 VDD.n1434 10.6151
R3455 VDD.n1434 VDD.n1432 10.6151
R3456 VDD.n1432 VDD.n1431 10.6151
R3457 VDD.n1431 VDD.n1429 10.6151
R3458 VDD.n1429 VDD.n1428 10.6151
R3459 VDD.n1428 VDD.n1426 10.6151
R3460 VDD.n1426 VDD.n1425 10.6151
R3461 VDD.n1425 VDD.n1423 10.6151
R3462 VDD.n1423 VDD.n1422 10.6151
R3463 VDD.n1422 VDD.n1420 10.6151
R3464 VDD.n1420 VDD.n1419 10.6151
R3465 VDD.n1419 VDD.n1417 10.6151
R3466 VDD.n1417 VDD.n1416 10.6151
R3467 VDD.n1416 VDD.n1345 10.6151
R3468 VDD.n1345 VDD.n1344 10.6151
R3469 VDD.n1344 VDD.n1342 10.6151
R3470 VDD.n1342 VDD.n1341 10.6151
R3471 VDD.n1341 VDD.n1339 10.6151
R3472 VDD.n1339 VDD.n1338 10.6151
R3473 VDD.n1338 VDD.n1336 10.6151
R3474 VDD.n1336 VDD.n532 10.6151
R3475 VDD.n1617 VDD.n532 10.6151
R3476 VDD.n1618 VDD.n1617 10.6151
R3477 VDD.n1621 VDD.n1618 10.6151
R3478 VDD.n1621 VDD.n1620 10.6151
R3479 VDD.n1620 VDD.n1619 10.6151
R3480 VDD.n1619 VDD.n513 10.6151
R3481 VDD.n513 VDD.n511 10.6151
R3482 VDD.n1308 VDD.n611 10.6151
R3483 VDD.n1308 VDD.n1307 10.6151
R3484 VDD.n1314 VDD.n1307 10.6151
R3485 VDD.n1315 VDD.n1314 10.6151
R3486 VDD.n1316 VDD.n1315 10.6151
R3487 VDD.n1316 VDD.n1305 10.6151
R3488 VDD.n1322 VDD.n1305 10.6151
R3489 VDD.n1323 VDD.n1322 10.6151
R3490 VDD.n1324 VDD.n1323 10.6151
R3491 VDD.n1324 VDD.n1302 10.6151
R3492 VDD.n1465 VDD.n1302 10.6151
R3493 VDD.n1465 VDD.n1303 10.6151
R3494 VDD.n1460 VDD.n1303 10.6151
R3495 VDD.n1460 VDD.n1459 10.6151
R3496 VDD.n1459 VDD.n1329 10.6151
R3497 VDD.n1454 VDD.n1329 10.6151
R3498 VDD.n1454 VDD.n1453 10.6151
R3499 VDD.n1453 VDD.n1452 10.6151
R3500 VDD.n1452 VDD.n1331 10.6151
R3501 VDD.n1446 VDD.n1445 10.6151
R3502 VDD.n1445 VDD.n1444 10.6151
R3503 VDD.n1535 VDD.n1534 10.6151
R3504 VDD.n1536 VDD.n1535 10.6151
R3505 VDD.n1536 VDD.n599 10.6151
R3506 VDD.n1546 VDD.n599 10.6151
R3507 VDD.n1547 VDD.n1546 10.6151
R3508 VDD.n1548 VDD.n1547 10.6151
R3509 VDD.n1548 VDD.n587 10.6151
R3510 VDD.n1558 VDD.n587 10.6151
R3511 VDD.n1559 VDD.n1558 10.6151
R3512 VDD.n1560 VDD.n1559 10.6151
R3513 VDD.n1560 VDD.n575 10.6151
R3514 VDD.n1570 VDD.n575 10.6151
R3515 VDD.n1571 VDD.n1570 10.6151
R3516 VDD.n1572 VDD.n1571 10.6151
R3517 VDD.n1572 VDD.n563 10.6151
R3518 VDD.n1582 VDD.n563 10.6151
R3519 VDD.n1583 VDD.n1582 10.6151
R3520 VDD.n1584 VDD.n1583 10.6151
R3521 VDD.n1584 VDD.n551 10.6151
R3522 VDD.n1594 VDD.n551 10.6151
R3523 VDD.n1595 VDD.n1594 10.6151
R3524 VDD.n1596 VDD.n1595 10.6151
R3525 VDD.n1596 VDD.n539 10.6151
R3526 VDD.n1610 VDD.n539 10.6151
R3527 VDD.n1611 VDD.n1610 10.6151
R3528 VDD.n1613 VDD.n1611 10.6151
R3529 VDD.n1613 VDD.n1612 10.6151
R3530 VDD.n1612 VDD.n517 10.6151
R3531 VDD.n1685 VDD.n517 10.6151
R3532 VDD.n1686 VDD.n1685 10.6151
R3533 VDD.n1687 VDD.n1686 10.6151
R3534 VDD.n1687 VDD.n508 10.6151
R3535 VDD.n1900 VDD.n1899 10.6151
R3536 VDD.n1899 VDD.n1898 10.6151
R3537 VDD.n1898 VDD.n1896 10.6151
R3538 VDD.n1896 VDD.n1895 10.6151
R3539 VDD.n1895 VDD.n1893 10.6151
R3540 VDD.n1893 VDD.n1892 10.6151
R3541 VDD.n1892 VDD.n1890 10.6151
R3542 VDD.n1890 VDD.n1889 10.6151
R3543 VDD.n1889 VDD.n1887 10.6151
R3544 VDD.n1887 VDD.n1886 10.6151
R3545 VDD.n1886 VDD.n1789 10.6151
R3546 VDD.n1789 VDD.n1788 10.6151
R3547 VDD.n1788 VDD.n1786 10.6151
R3548 VDD.n1786 VDD.n1785 10.6151
R3549 VDD.n1785 VDD.n1783 10.6151
R3550 VDD.n1783 VDD.n1782 10.6151
R3551 VDD.n1782 VDD.n1780 10.6151
R3552 VDD.n1780 VDD.n1779 10.6151
R3553 VDD.n1779 VDD.n1777 10.6151
R3554 VDD.n1777 VDD.n1776 10.6151
R3555 VDD.n1776 VDD.n1774 10.6151
R3556 VDD.n1774 VDD.n1773 10.6151
R3557 VDD.n1773 VDD.n1771 10.6151
R3558 VDD.n1771 VDD.n1770 10.6151
R3559 VDD.n1770 VDD.n1768 10.6151
R3560 VDD.n1768 VDD.n1767 10.6151
R3561 VDD.n1767 VDD.n1765 10.6151
R3562 VDD.n1765 VDD.n1764 10.6151
R3563 VDD.n1764 VDD.n391 10.6151
R3564 VDD.n2072 VDD.n391 10.6151
R3565 VDD.n2073 VDD.n2072 10.6151
R3566 VDD.n2074 VDD.n2073 10.6151
R3567 VDD.n1947 VDD.n480 10.6151
R3568 VDD.n1942 VDD.n480 10.6151
R3569 VDD.n1942 VDD.n1941 10.6151
R3570 VDD.n1941 VDD.n1940 10.6151
R3571 VDD.n1940 VDD.n1937 10.6151
R3572 VDD.n1937 VDD.n1936 10.6151
R3573 VDD.n1936 VDD.n1933 10.6151
R3574 VDD.n1933 VDD.n1932 10.6151
R3575 VDD.n1932 VDD.n1929 10.6151
R3576 VDD.n1929 VDD.n1928 10.6151
R3577 VDD.n1928 VDD.n1925 10.6151
R3578 VDD.n1925 VDD.n1924 10.6151
R3579 VDD.n1924 VDD.n1921 10.6151
R3580 VDD.n1921 VDD.n1920 10.6151
R3581 VDD.n1920 VDD.n1917 10.6151
R3582 VDD.n1917 VDD.n1916 10.6151
R3583 VDD.n1916 VDD.n1913 10.6151
R3584 VDD.n1913 VDD.n1912 10.6151
R3585 VDD.n1912 VDD.n1909 10.6151
R3586 VDD.n1907 VDD.n1904 10.6151
R3587 VDD.n1904 VDD.n1903 10.6151
R3588 VDD.n1949 VDD.n1948 10.6151
R3589 VDD.n1949 VDD.n468 10.6151
R3590 VDD.n1959 VDD.n468 10.6151
R3591 VDD.n1960 VDD.n1959 10.6151
R3592 VDD.n1961 VDD.n1960 10.6151
R3593 VDD.n1961 VDD.n456 10.6151
R3594 VDD.n1971 VDD.n456 10.6151
R3595 VDD.n1972 VDD.n1971 10.6151
R3596 VDD.n1973 VDD.n1972 10.6151
R3597 VDD.n1973 VDD.n445 10.6151
R3598 VDD.n1983 VDD.n445 10.6151
R3599 VDD.n1984 VDD.n1983 10.6151
R3600 VDD.n1985 VDD.n1984 10.6151
R3601 VDD.n1985 VDD.n433 10.6151
R3602 VDD.n1995 VDD.n433 10.6151
R3603 VDD.n1996 VDD.n1995 10.6151
R3604 VDD.n1997 VDD.n1996 10.6151
R3605 VDD.n1997 VDD.n421 10.6151
R3606 VDD.n2007 VDD.n421 10.6151
R3607 VDD.n2008 VDD.n2007 10.6151
R3608 VDD.n2009 VDD.n2008 10.6151
R3609 VDD.n2009 VDD.n409 10.6151
R3610 VDD.n2019 VDD.n409 10.6151
R3611 VDD.n2020 VDD.n2019 10.6151
R3612 VDD.n2021 VDD.n2020 10.6151
R3613 VDD.n2021 VDD.n396 10.6151
R3614 VDD.n2065 VDD.n396 10.6151
R3615 VDD.n2066 VDD.n2065 10.6151
R3616 VDD.n2067 VDD.n2066 10.6151
R3617 VDD.n2067 VDD.n373 10.6151
R3618 VDD.n2119 VDD.n373 10.6151
R3619 VDD.n2119 VDD.n2118 10.6151
R3620 VDD.n2117 VDD.n374 10.6151
R3621 VDD.n2112 VDD.n374 10.6151
R3622 VDD.n2112 VDD.n2111 10.6151
R3623 VDD.n2111 VDD.n2110 10.6151
R3624 VDD.n2110 VDD.n376 10.6151
R3625 VDD.n2105 VDD.n376 10.6151
R3626 VDD.n2105 VDD.n2104 10.6151
R3627 VDD.n2104 VDD.n2103 10.6151
R3628 VDD.n2103 VDD.n379 10.6151
R3629 VDD.n2098 VDD.n379 10.6151
R3630 VDD.n2098 VDD.n311 10.6151
R3631 VDD.n2094 VDD.n311 10.6151
R3632 VDD.n2094 VDD.n2093 10.6151
R3633 VDD.n2093 VDD.n2092 10.6151
R3634 VDD.n2092 VDD.n382 10.6151
R3635 VDD.n2087 VDD.n382 10.6151
R3636 VDD.n2087 VDD.n2086 10.6151
R3637 VDD.n2086 VDD.n2085 10.6151
R3638 VDD.n2085 VDD.n385 10.6151
R3639 VDD.n2080 VDD.n2079 10.6151
R3640 VDD.n2079 VDD.n2078 10.6151
R3641 VDD.n2052 VDD.n2051 10.6151
R3642 VDD.n2051 VDD.n2050 10.6151
R3643 VDD.n2050 VDD.n2030 10.6151
R3644 VDD.n2045 VDD.n2030 10.6151
R3645 VDD.n2045 VDD.n2044 10.6151
R3646 VDD.n2044 VDD.n2043 10.6151
R3647 VDD.n2043 VDD.n2033 10.6151
R3648 VDD.n2038 VDD.n2033 10.6151
R3649 VDD.n2038 VDD.n2037 10.6151
R3650 VDD.n2037 VDD.n351 10.6151
R3651 VDD.n2147 VDD.n351 10.6151
R3652 VDD.n2147 VDD.n352 10.6151
R3653 VDD.n355 VDD.n352 10.6151
R3654 VDD.n2140 VDD.n355 10.6151
R3655 VDD.n2140 VDD.n2139 10.6151
R3656 VDD.n2139 VDD.n2138 10.6151
R3657 VDD.n2138 VDD.n357 10.6151
R3658 VDD.n2133 VDD.n357 10.6151
R3659 VDD.n2133 VDD.n2132 10.6151
R3660 VDD.n2130 VDD.n362 10.6151
R3661 VDD.n2125 VDD.n362 10.6151
R3662 VDD.n1840 VDD.n1839 10.6151
R3663 VDD.n1842 VDD.n1840 10.6151
R3664 VDD.n1843 VDD.n1842 10.6151
R3665 VDD.n1845 VDD.n1843 10.6151
R3666 VDD.n1846 VDD.n1845 10.6151
R3667 VDD.n1848 VDD.n1846 10.6151
R3668 VDD.n1849 VDD.n1848 10.6151
R3669 VDD.n1851 VDD.n1849 10.6151
R3670 VDD.n1852 VDD.n1851 10.6151
R3671 VDD.n1882 VDD.n1852 10.6151
R3672 VDD.n1882 VDD.n1881 10.6151
R3673 VDD.n1881 VDD.n1880 10.6151
R3674 VDD.n1880 VDD.n1878 10.6151
R3675 VDD.n1878 VDD.n1877 10.6151
R3676 VDD.n1877 VDD.n1875 10.6151
R3677 VDD.n1875 VDD.n1874 10.6151
R3678 VDD.n1874 VDD.n1872 10.6151
R3679 VDD.n1872 VDD.n1871 10.6151
R3680 VDD.n1871 VDD.n1869 10.6151
R3681 VDD.n1869 VDD.n1868 10.6151
R3682 VDD.n1868 VDD.n1866 10.6151
R3683 VDD.n1866 VDD.n1865 10.6151
R3684 VDD.n1865 VDD.n1863 10.6151
R3685 VDD.n1863 VDD.n1862 10.6151
R3686 VDD.n1862 VDD.n1860 10.6151
R3687 VDD.n1860 VDD.n1859 10.6151
R3688 VDD.n1859 VDD.n1857 10.6151
R3689 VDD.n1857 VDD.n1856 10.6151
R3690 VDD.n1856 VDD.n1853 10.6151
R3691 VDD.n1853 VDD.n365 10.6151
R3692 VDD.n2123 VDD.n365 10.6151
R3693 VDD.n2124 VDD.n2123 10.6151
R3694 VDD.n1795 VDD.n1794 10.6151
R3695 VDD.n1798 VDD.n1795 10.6151
R3696 VDD.n1799 VDD.n1798 10.6151
R3697 VDD.n1802 VDD.n1799 10.6151
R3698 VDD.n1803 VDD.n1802 10.6151
R3699 VDD.n1806 VDD.n1803 10.6151
R3700 VDD.n1807 VDD.n1806 10.6151
R3701 VDD.n1810 VDD.n1807 10.6151
R3702 VDD.n1811 VDD.n1810 10.6151
R3703 VDD.n1814 VDD.n1811 10.6151
R3704 VDD.n1815 VDD.n1814 10.6151
R3705 VDD.n1818 VDD.n1815 10.6151
R3706 VDD.n1819 VDD.n1818 10.6151
R3707 VDD.n1822 VDD.n1819 10.6151
R3708 VDD.n1823 VDD.n1822 10.6151
R3709 VDD.n1826 VDD.n1823 10.6151
R3710 VDD.n1827 VDD.n1826 10.6151
R3711 VDD.n1830 VDD.n1827 10.6151
R3712 VDD.n1831 VDD.n1830 10.6151
R3713 VDD.n1836 VDD.n1834 10.6151
R3714 VDD.n1837 VDD.n1836 10.6151
R3715 VDD.n1953 VDD.n474 10.6151
R3716 VDD.n1954 VDD.n1953 10.6151
R3717 VDD.n1955 VDD.n1954 10.6151
R3718 VDD.n1955 VDD.n462 10.6151
R3719 VDD.n1965 VDD.n462 10.6151
R3720 VDD.n1966 VDD.n1965 10.6151
R3721 VDD.n1967 VDD.n1966 10.6151
R3722 VDD.n1967 VDD.n450 10.6151
R3723 VDD.n1977 VDD.n450 10.6151
R3724 VDD.n1978 VDD.n1977 10.6151
R3725 VDD.n1979 VDD.n1978 10.6151
R3726 VDD.n1979 VDD.n438 10.6151
R3727 VDD.n1989 VDD.n438 10.6151
R3728 VDD.n1990 VDD.n1989 10.6151
R3729 VDD.n1991 VDD.n1990 10.6151
R3730 VDD.n1991 VDD.n427 10.6151
R3731 VDD.n2001 VDD.n427 10.6151
R3732 VDD.n2002 VDD.n2001 10.6151
R3733 VDD.n2003 VDD.n2002 10.6151
R3734 VDD.n2003 VDD.n415 10.6151
R3735 VDD.n2013 VDD.n415 10.6151
R3736 VDD.n2014 VDD.n2013 10.6151
R3737 VDD.n2015 VDD.n2014 10.6151
R3738 VDD.n2015 VDD.n403 10.6151
R3739 VDD.n2025 VDD.n403 10.6151
R3740 VDD.n2026 VDD.n2025 10.6151
R3741 VDD.n2061 VDD.n2026 10.6151
R3742 VDD.n2061 VDD.n2060 10.6151
R3743 VDD.n2060 VDD.n2059 10.6151
R3744 VDD.n2059 VDD.n2058 10.6151
R3745 VDD.n2058 VDD.n2056 10.6151
R3746 VDD.n2056 VDD.n2055 10.6151
R3747 VDD.n1530 VDD.n604 10.6151
R3748 VDD.n1540 VDD.n604 10.6151
R3749 VDD.n1541 VDD.n1540 10.6151
R3750 VDD.n1542 VDD.n1541 10.6151
R3751 VDD.n1542 VDD.n593 10.6151
R3752 VDD.n1552 VDD.n593 10.6151
R3753 VDD.n1553 VDD.n1552 10.6151
R3754 VDD.n1554 VDD.n1553 10.6151
R3755 VDD.n1554 VDD.n581 10.6151
R3756 VDD.n1564 VDD.n581 10.6151
R3757 VDD.n1565 VDD.n1564 10.6151
R3758 VDD.n1566 VDD.n1565 10.6151
R3759 VDD.n1566 VDD.n569 10.6151
R3760 VDD.n1576 VDD.n569 10.6151
R3761 VDD.n1577 VDD.n1576 10.6151
R3762 VDD.n1578 VDD.n1577 10.6151
R3763 VDD.n1578 VDD.n558 10.6151
R3764 VDD.n1588 VDD.n558 10.6151
R3765 VDD.n1589 VDD.n1588 10.6151
R3766 VDD.n1590 VDD.n1589 10.6151
R3767 VDD.n1590 VDD.n546 10.6151
R3768 VDD.n1600 VDD.n546 10.6151
R3769 VDD.n1601 VDD.n1600 10.6151
R3770 VDD.n1606 VDD.n1601 10.6151
R3771 VDD.n1606 VDD.n1605 10.6151
R3772 VDD.n1605 VDD.n1604 10.6151
R3773 VDD.n1604 VDD.n1603 10.6151
R3774 VDD.n1603 VDD.n524 10.6151
R3775 VDD.n1681 VDD.n524 10.6151
R3776 VDD.n1681 VDD.n1680 10.6151
R3777 VDD.n1680 VDD.n1679 10.6151
R3778 VDD.n1679 VDD.n1678 10.6151
R3779 VDD.n1675 VDD.n1674 10.6151
R3780 VDD.n1674 VDD.n1671 10.6151
R3781 VDD.n1671 VDD.n1670 10.6151
R3782 VDD.n1670 VDD.n1667 10.6151
R3783 VDD.n1667 VDD.n1666 10.6151
R3784 VDD.n1666 VDD.n1663 10.6151
R3785 VDD.n1663 VDD.n1662 10.6151
R3786 VDD.n1662 VDD.n1659 10.6151
R3787 VDD.n1659 VDD.n1658 10.6151
R3788 VDD.n1658 VDD.n1655 10.6151
R3789 VDD.n1655 VDD.n1654 10.6151
R3790 VDD.n1654 VDD.n1651 10.6151
R3791 VDD.n1651 VDD.n1650 10.6151
R3792 VDD.n1650 VDD.n1647 10.6151
R3793 VDD.n1647 VDD.n1646 10.6151
R3794 VDD.n1646 VDD.n1643 10.6151
R3795 VDD.n1643 VDD.n1642 10.6151
R3796 VDD.n1642 VDD.n1639 10.6151
R3797 VDD.n1639 VDD.n1638 10.6151
R3798 VDD.n1635 VDD.n1634 10.6151
R3799 VDD.n1634 VDD.n1632 10.6151
R3800 VDD.n1376 VDD.n1374 10.6151
R3801 VDD.n1377 VDD.n1376 10.6151
R3802 VDD.n1379 VDD.n1377 10.6151
R3803 VDD.n1380 VDD.n1379 10.6151
R3804 VDD.n1382 VDD.n1380 10.6151
R3805 VDD.n1383 VDD.n1382 10.6151
R3806 VDD.n1385 VDD.n1383 10.6151
R3807 VDD.n1386 VDD.n1385 10.6151
R3808 VDD.n1388 VDD.n1386 10.6151
R3809 VDD.n1389 VDD.n1388 10.6151
R3810 VDD.n1391 VDD.n1389 10.6151
R3811 VDD.n1392 VDD.n1391 10.6151
R3812 VDD.n1394 VDD.n1392 10.6151
R3813 VDD.n1395 VDD.n1394 10.6151
R3814 VDD.n1397 VDD.n1395 10.6151
R3815 VDD.n1398 VDD.n1397 10.6151
R3816 VDD.n1412 VDD.n1398 10.6151
R3817 VDD.n1412 VDD.n1411 10.6151
R3818 VDD.n1411 VDD.n1410 10.6151
R3819 VDD.n1410 VDD.n1408 10.6151
R3820 VDD.n1408 VDD.n1407 10.6151
R3821 VDD.n1407 VDD.n1405 10.6151
R3822 VDD.n1405 VDD.n1404 10.6151
R3823 VDD.n1404 VDD.n1402 10.6151
R3824 VDD.n1402 VDD.n1401 10.6151
R3825 VDD.n1401 VDD.n1399 10.6151
R3826 VDD.n1399 VDD.n528 10.6151
R3827 VDD.n1625 VDD.n528 10.6151
R3828 VDD.n1626 VDD.n1625 10.6151
R3829 VDD.n1628 VDD.n1626 10.6151
R3830 VDD.n1629 VDD.n1628 10.6151
R3831 VDD.n1631 VDD.n1629 10.6151
R3832 VDD.n1528 VDD.n1527 10.6151
R3833 VDD.n1527 VDD.n618 10.6151
R3834 VDD.n1521 VDD.n618 10.6151
R3835 VDD.n1521 VDD.n1520 10.6151
R3836 VDD.n1520 VDD.n1519 10.6151
R3837 VDD.n1519 VDD.n620 10.6151
R3838 VDD.n1513 VDD.n620 10.6151
R3839 VDD.n1513 VDD.n1512 10.6151
R3840 VDD.n1512 VDD.n1511 10.6151
R3841 VDD.n1511 VDD.n622 10.6151
R3842 VDD.n1505 VDD.n622 10.6151
R3843 VDD.n1505 VDD.n624 10.6151
R3844 VDD.n1352 VDD.n624 10.6151
R3845 VDD.n1357 VDD.n1352 10.6151
R3846 VDD.n1358 VDD.n1357 10.6151
R3847 VDD.n1359 VDD.n1358 10.6151
R3848 VDD.n1359 VDD.n1350 10.6151
R3849 VDD.n1365 VDD.n1350 10.6151
R3850 VDD.n1366 VDD.n1365 10.6151
R3851 VDD.n1368 VDD.n1346 10.6151
R3852 VDD.n1373 VDD.n1346 10.6151
R3853 VDD.n1002 VDD.t33 10.3006
R3854 VDD.t22 VDD.n641 10.3006
R3855 VDD.n2282 VDD.t44 10.3006
R3856 VDD.t51 VDD.n2491 10.3006
R3857 VDD.n1532 VDD.n606 10.1513
R3858 VDD.n1538 VDD.n606 10.1513
R3859 VDD.n1538 VDD.n609 10.1513
R3860 VDD.n1550 VDD.n595 10.1513
R3861 VDD.n1550 VDD.n589 10.1513
R3862 VDD.n1556 VDD.n589 10.1513
R3863 VDD.n1562 VDD.n583 10.1513
R3864 VDD.n1568 VDD.n577 10.1513
R3865 VDD.n1574 VDD.n571 10.1513
R3866 VDD.n1580 VDD.n565 10.1513
R3867 VDD.n1586 VDD.n553 10.1513
R3868 VDD.n1592 VDD.n553 10.1513
R3869 VDD.n1592 VDD.n556 10.1513
R3870 VDD.n1608 VDD.n541 10.1513
R3871 VDD.n1608 VDD.n534 10.1513
R3872 VDD.n1615 VDD.n534 10.1513
R3873 VDD.n1623 VDD.n530 10.1513
R3874 VDD.n1683 VDD.n521 10.1513
R3875 VDD.n1689 VDD.n482 10.1513
R3876 VDD.n1951 VDD.n476 10.1513
R3877 VDD.n1957 VDD.n470 10.1513
R3878 VDD.n1963 VDD.n464 10.1513
R3879 VDD.n1969 VDD.n458 10.1513
R3880 VDD.n1969 VDD.n452 10.1513
R3881 VDD.n1975 VDD.n452 10.1513
R3882 VDD.n1981 VDD.n440 10.1513
R3883 VDD.n1987 VDD.n440 10.1513
R3884 VDD.n1987 VDD.n443 10.1513
R3885 VDD.n1999 VDD.n429 10.1513
R3886 VDD.n2005 VDD.n423 10.1513
R3887 VDD.n2011 VDD.n417 10.1513
R3888 VDD.n2017 VDD.n411 10.1513
R3889 VDD.n2023 VDD.n405 10.1513
R3890 VDD.n2023 VDD.n398 10.1513
R3891 VDD.n2063 VDD.n398 10.1513
R3892 VDD.n2069 VDD.n367 10.1513
R3893 VDD.n2121 VDD.n367 10.1513
R3894 VDD.n2121 VDD.n369 10.1513
R3895 VDD.n1544 VDD.t71 10.0021
R3896 VDD.n1623 VDD.t64 10.0021
R3897 VDD.t78 VDD.n464 10.0021
R3898 VDD.n1854 VDD.t37 10.0021
R3899 VDD.t0 VDD.n565 9.70352
R3900 VDD.n1414 VDD.t17 9.70352
R3901 VDD.n1993 VDD.t101 9.70352
R3902 VDD.n1999 VDD.t18 9.70352
R3903 VDD.n1466 VDD.n1465 9.60081
R3904 VDD.n2260 VDD.n311 9.60081
R3905 VDD.n2176 VDD.n2147 9.60081
R3906 VDD.n1505 VDD.n1504 9.60081
R3907 VDD.n1078 VDD.n1077 9.3005
R3908 VDD.n1079 VDD.n697 9.3005
R3909 VDD.n1081 VDD.n1080 9.3005
R3910 VDD.n687 VDD.n686 9.3005
R3911 VDD.n1094 VDD.n1093 9.3005
R3912 VDD.n1095 VDD.n685 9.3005
R3913 VDD.n1097 VDD.n1096 9.3005
R3914 VDD.n675 VDD.n674 9.3005
R3915 VDD.n1110 VDD.n1109 9.3005
R3916 VDD.n1111 VDD.n673 9.3005
R3917 VDD.n1113 VDD.n1112 9.3005
R3918 VDD.n663 VDD.n662 9.3005
R3919 VDD.n1126 VDD.n1125 9.3005
R3920 VDD.n1127 VDD.n661 9.3005
R3921 VDD.n1129 VDD.n1128 9.3005
R3922 VDD.n651 VDD.n650 9.3005
R3923 VDD.n1142 VDD.n1141 9.3005
R3924 VDD.n1143 VDD.n649 9.3005
R3925 VDD.n1484 VDD.n1483 9.3005
R3926 VDD.n1284 VDD.n1171 9.3005
R3927 VDD.n1283 VDD.n1282 9.3005
R3928 VDD.n1176 VDD.n1175 9.3005
R3929 VDD.n1277 VDD.n1179 9.3005
R3930 VDD.n1276 VDD.n1180 9.3005
R3931 VDD.n1275 VDD.n1181 9.3005
R3932 VDD.n1185 VDD.n1182 9.3005
R3933 VDD.n1270 VDD.n1186 9.3005
R3934 VDD.n1269 VDD.n1187 9.3005
R3935 VDD.n1268 VDD.n1188 9.3005
R3936 VDD.n1192 VDD.n1189 9.3005
R3937 VDD.n1263 VDD.n1193 9.3005
R3938 VDD.n1262 VDD.n1194 9.3005
R3939 VDD.n1261 VDD.n1195 9.3005
R3940 VDD.n1199 VDD.n1196 9.3005
R3941 VDD.n1256 VDD.n1200 9.3005
R3942 VDD.n1255 VDD.n1201 9.3005
R3943 VDD.n1254 VDD.n1202 9.3005
R3944 VDD.n1209 VDD.n1203 9.3005
R3945 VDD.n1249 VDD.n1248 9.3005
R3946 VDD.n1247 VDD.n1206 9.3005
R3947 VDD.n1246 VDD.n1245 9.3005
R3948 VDD.n1211 VDD.n1210 9.3005
R3949 VDD.n1240 VDD.n1214 9.3005
R3950 VDD.n1239 VDD.n1215 9.3005
R3951 VDD.n1238 VDD.n1216 9.3005
R3952 VDD.n1220 VDD.n1217 9.3005
R3953 VDD.n1233 VDD.n1221 9.3005
R3954 VDD.n1232 VDD.n625 9.3005
R3955 VDD.n1286 VDD.n1285 9.3005
R3956 VDD.n1480 VDD.n1144 9.3005
R3957 VDD.n1148 VDD.n1145 9.3005
R3958 VDD.n1475 VDD.n1149 9.3005
R3959 VDD.n1474 VDD.n1150 9.3005
R3960 VDD.n1473 VDD.n1151 9.3005
R3961 VDD.n1156 VDD.n1152 9.3005
R3962 VDD.n1159 VDD.n1157 9.3005
R3963 VDD.n1164 VDD.n1162 9.3005
R3964 VDD.n1293 VDD.n1165 9.3005
R3965 VDD.n1292 VDD.n1166 9.3005
R3966 VDD.n1291 VDD.n1167 9.3005
R3967 VDD.n1174 VDD.n1168 9.3005
R3968 VDD.n1482 VDD.n1481 9.3005
R3969 VDD.n2200 VDD.n2199 9.3005
R3970 VDD.n2203 VDD.n338 9.3005
R3971 VDD.n2204 VDD.n337 9.3005
R3972 VDD.n2207 VDD.n336 9.3005
R3973 VDD.n2208 VDD.n335 9.3005
R3974 VDD.n2211 VDD.n334 9.3005
R3975 VDD.n2212 VDD.n333 9.3005
R3976 VDD.n2215 VDD.n332 9.3005
R3977 VDD.n2216 VDD.n331 9.3005
R3978 VDD.n2219 VDD.n330 9.3005
R3979 VDD.n2220 VDD.n329 9.3005
R3980 VDD.n2223 VDD.n328 9.3005
R3981 VDD.n2224 VDD.n327 9.3005
R3982 VDD.n2227 VDD.n326 9.3005
R3983 VDD.n2228 VDD.n325 9.3005
R3984 VDD.n2231 VDD.n324 9.3005
R3985 VDD.n2232 VDD.n323 9.3005
R3986 VDD.n2235 VDD.n322 9.3005
R3987 VDD.n2239 VDD.n2238 9.3005
R3988 VDD.n2240 VDD.n321 9.3005
R3989 VDD.n2244 VDD.n2241 9.3005
R3990 VDD.n2247 VDD.n320 9.3005
R3991 VDD.n2248 VDD.n319 9.3005
R3992 VDD.n2251 VDD.n318 9.3005
R3993 VDD.n2252 VDD.n317 9.3005
R3994 VDD.n2255 VDD.n316 9.3005
R3995 VDD.n2257 VDD.n310 9.3005
R3996 VDD.n2265 VDD.n308 9.3005
R3997 VDD.n2266 VDD.n307 9.3005
R3998 VDD.n2269 VDD.n306 9.3005
R3999 VDD.n2270 VDD.n305 9.3005
R4000 VDD.n2271 VDD.n304 9.3005
R4001 VDD.n273 VDD.n272 9.3005
R4002 VDD.n2277 VDD.n2276 9.3005
R4003 VDD.n2278 VDD.n271 9.3005
R4004 VDD.n2280 VDD.n2279 9.3005
R4005 VDD.n261 VDD.n260 9.3005
R4006 VDD.n2293 VDD.n2292 9.3005
R4007 VDD.n2294 VDD.n259 9.3005
R4008 VDD.n2296 VDD.n2295 9.3005
R4009 VDD.n249 VDD.n248 9.3005
R4010 VDD.n2309 VDD.n2308 9.3005
R4011 VDD.n2310 VDD.n247 9.3005
R4012 VDD.n2312 VDD.n2311 9.3005
R4013 VDD.n237 VDD.n236 9.3005
R4014 VDD.n2325 VDD.n2324 9.3005
R4015 VDD.n2326 VDD.n235 9.3005
R4016 VDD.n2328 VDD.n2327 9.3005
R4017 VDD.n225 VDD.n224 9.3005
R4018 VDD.n2341 VDD.n2340 9.3005
R4019 VDD.n2342 VDD.n223 9.3005
R4020 VDD.n2344 VDD.n2343 9.3005
R4021 VDD.n47 VDD.n45 9.3005
R4022 VDD.n2527 VDD.n2526 9.3005
R4023 VDD.n48 VDD.n46 9.3005
R4024 VDD.n2520 VDD.n57 9.3005
R4025 VDD.n2519 VDD.n58 9.3005
R4026 VDD.n2518 VDD.n59 9.3005
R4027 VDD.n66 VDD.n60 9.3005
R4028 VDD.n2512 VDD.n67 9.3005
R4029 VDD.n2511 VDD.n68 9.3005
R4030 VDD.n2510 VDD.n69 9.3005
R4031 VDD.n78 VDD.n70 9.3005
R4032 VDD.n2504 VDD.n79 9.3005
R4033 VDD.n2503 VDD.n80 9.3005
R4034 VDD.n2502 VDD.n81 9.3005
R4035 VDD.n89 VDD.n82 9.3005
R4036 VDD.n2496 VDD.n90 9.3005
R4037 VDD.n2495 VDD.n91 9.3005
R4038 VDD.n2494 VDD.n92 9.3005
R4039 VDD.n100 VDD.n93 9.3005
R4040 VDD.n2488 VDD.n2487 9.3005
R4041 VDD.n2484 VDD.n101 9.3005
R4042 VDD.n2483 VDD.n104 9.3005
R4043 VDD.n108 VDD.n105 9.3005
R4044 VDD.n109 VDD.n106 9.3005
R4045 VDD.n2476 VDD.n110 9.3005
R4046 VDD.n2475 VDD.n111 9.3005
R4047 VDD.n2474 VDD.n112 9.3005
R4048 VDD.n116 VDD.n113 9.3005
R4049 VDD.n2469 VDD.n117 9.3005
R4050 VDD.n2468 VDD.n118 9.3005
R4051 VDD.n2467 VDD.n119 9.3005
R4052 VDD.n123 VDD.n120 9.3005
R4053 VDD.n2462 VDD.n124 9.3005
R4054 VDD.n2461 VDD.n125 9.3005
R4055 VDD.n2460 VDD.n126 9.3005
R4056 VDD.n133 VDD.n127 9.3005
R4057 VDD.n2455 VDD.n2454 9.3005
R4058 VDD.n2453 VDD.n130 9.3005
R4059 VDD.n2452 VDD.n2451 9.3005
R4060 VDD.n135 VDD.n134 9.3005
R4061 VDD.n2446 VDD.n138 9.3005
R4062 VDD.n2445 VDD.n139 9.3005
R4063 VDD.n2444 VDD.n140 9.3005
R4064 VDD.n144 VDD.n141 9.3005
R4065 VDD.n2439 VDD.n145 9.3005
R4066 VDD.n2438 VDD.n146 9.3005
R4067 VDD.n2437 VDD.n147 9.3005
R4068 VDD.n151 VDD.n148 9.3005
R4069 VDD.n2432 VDD.n152 9.3005
R4070 VDD.n2431 VDD.n153 9.3005
R4071 VDD.n2430 VDD.n154 9.3005
R4072 VDD.n158 VDD.n155 9.3005
R4073 VDD.n2425 VDD.n159 9.3005
R4074 VDD.n2424 VDD.n160 9.3005
R4075 VDD.n2423 VDD.n161 9.3005
R4076 VDD.n168 VDD.n162 9.3005
R4077 VDD.n2418 VDD.n2417 9.3005
R4078 VDD.n2416 VDD.n165 9.3005
R4079 VDD.n2415 VDD.n2414 9.3005
R4080 VDD.n170 VDD.n169 9.3005
R4081 VDD.n2409 VDD.n173 9.3005
R4082 VDD.n2408 VDD.n174 9.3005
R4083 VDD.n2407 VDD.n175 9.3005
R4084 VDD.n179 VDD.n176 9.3005
R4085 VDD.n2402 VDD.n180 9.3005
R4086 VDD.n2401 VDD.n181 9.3005
R4087 VDD.n2400 VDD.n182 9.3005
R4088 VDD.n186 VDD.n183 9.3005
R4089 VDD.n2395 VDD.n187 9.3005
R4090 VDD.n2394 VDD.n188 9.3005
R4091 VDD.n2393 VDD.n189 9.3005
R4092 VDD.n193 VDD.n190 9.3005
R4093 VDD.n2388 VDD.n194 9.3005
R4094 VDD.n2387 VDD.n195 9.3005
R4095 VDD.n2386 VDD.n196 9.3005
R4096 VDD.n202 VDD.n197 9.3005
R4097 VDD.n2381 VDD.n2380 9.3005
R4098 VDD.n2486 VDD.n2485 9.3005
R4099 VDD.n2285 VDD.n2284 9.3005
R4100 VDD.n2286 VDD.n265 9.3005
R4101 VDD.n2288 VDD.n2287 9.3005
R4102 VDD.n254 VDD.n253 9.3005
R4103 VDD.n2301 VDD.n2300 9.3005
R4104 VDD.n2302 VDD.n252 9.3005
R4105 VDD.n2304 VDD.n2303 9.3005
R4106 VDD.n243 VDD.n242 9.3005
R4107 VDD.n2317 VDD.n2316 9.3005
R4108 VDD.n2318 VDD.n241 9.3005
R4109 VDD.n2320 VDD.n2319 9.3005
R4110 VDD.n230 VDD.n229 9.3005
R4111 VDD.n2333 VDD.n2332 9.3005
R4112 VDD.n2334 VDD.n228 9.3005
R4113 VDD.n2336 VDD.n2335 9.3005
R4114 VDD.n218 VDD.n217 9.3005
R4115 VDD.n2349 VDD.n2348 9.3005
R4116 VDD.n2350 VDD.n216 9.3005
R4117 VDD.n2352 VDD.n2351 9.3005
R4118 VDD.n2353 VDD.n215 9.3005
R4119 VDD.n2355 VDD.n2354 9.3005
R4120 VDD.n2356 VDD.n214 9.3005
R4121 VDD.n2358 VDD.n2357 9.3005
R4122 VDD.n2359 VDD.n212 9.3005
R4123 VDD.n2361 VDD.n2360 9.3005
R4124 VDD.n2362 VDD.n211 9.3005
R4125 VDD.n2364 VDD.n2363 9.3005
R4126 VDD.n2365 VDD.n209 9.3005
R4127 VDD.n2367 VDD.n2366 9.3005
R4128 VDD.n2368 VDD.n208 9.3005
R4129 VDD.n2370 VDD.n2369 9.3005
R4130 VDD.n2371 VDD.n206 9.3005
R4131 VDD.n2373 VDD.n2372 9.3005
R4132 VDD.n2374 VDD.n205 9.3005
R4133 VDD.n2376 VDD.n2375 9.3005
R4134 VDD.n2377 VDD.n203 9.3005
R4135 VDD.n2379 VDD.n2378 9.3005
R4136 VDD.n267 VDD.n266 9.3005
R4137 VDD.n2158 VDD.n2157 9.3005
R4138 VDD.n2163 VDD.n2156 9.3005
R4139 VDD.n2164 VDD.n2155 9.3005
R4140 VDD.n2167 VDD.n2154 9.3005
R4141 VDD.n2168 VDD.n2153 9.3005
R4142 VDD.n2171 VDD.n2152 9.3005
R4143 VDD.n2173 VDD.n350 9.3005
R4144 VDD.n2181 VDD.n348 9.3005
R4145 VDD.n2182 VDD.n347 9.3005
R4146 VDD.n2185 VDD.n346 9.3005
R4147 VDD.n2186 VDD.n345 9.3005
R4148 VDD.n2189 VDD.n344 9.3005
R4149 VDD.n2190 VDD.n343 9.3005
R4150 VDD.n2193 VDD.n342 9.3005
R4151 VDD.n2197 VDD.n2196 9.3005
R4152 VDD.n2198 VDD.n339 9.3005
R4153 VDD.n1503 VDD.n1502 9.3005
R4154 VDD.n1501 VDD.n628 9.3005
R4155 VDD.n1500 VDD.n1499 9.3005
R4156 VDD.n1498 VDD.n633 9.3005
R4157 VDD.n1497 VDD.n1496 9.3005
R4158 VDD.n1495 VDD.n634 9.3005
R4159 VDD.n1491 VDD.n1490 9.3005
R4160 VDD.n1005 VDD.n1004 9.3005
R4161 VDD.n1006 VDD.n781 9.3005
R4162 VDD.n1008 VDD.n1007 9.3005
R4163 VDD.n770 VDD.n769 9.3005
R4164 VDD.n1021 VDD.n1020 9.3005
R4165 VDD.n1022 VDD.n768 9.3005
R4166 VDD.n1024 VDD.n1023 9.3005
R4167 VDD.n759 VDD.n758 9.3005
R4168 VDD.n1037 VDD.n1036 9.3005
R4169 VDD.n1038 VDD.n757 9.3005
R4170 VDD.n1040 VDD.n1039 9.3005
R4171 VDD.n746 VDD.n745 9.3005
R4172 VDD.n1053 VDD.n1052 9.3005
R4173 VDD.n1054 VDD.n744 9.3005
R4174 VDD.n1056 VDD.n1055 9.3005
R4175 VDD.n735 VDD.n734 9.3005
R4176 VDD.n1070 VDD.n1069 9.3005
R4177 VDD.n1071 VDD.n733 9.3005
R4178 VDD.n1073 VDD.n1072 9.3005
R4179 VDD.n692 VDD.n691 9.3005
R4180 VDD.n1086 VDD.n1085 9.3005
R4181 VDD.n1087 VDD.n690 9.3005
R4182 VDD.n1089 VDD.n1088 9.3005
R4183 VDD.n681 VDD.n680 9.3005
R4184 VDD.n1102 VDD.n1101 9.3005
R4185 VDD.n1103 VDD.n679 9.3005
R4186 VDD.n1105 VDD.n1104 9.3005
R4187 VDD.n668 VDD.n667 9.3005
R4188 VDD.n1118 VDD.n1117 9.3005
R4189 VDD.n1119 VDD.n666 9.3005
R4190 VDD.n1121 VDD.n1120 9.3005
R4191 VDD.n657 VDD.n656 9.3005
R4192 VDD.n1134 VDD.n1133 9.3005
R4193 VDD.n1135 VDD.n655 9.3005
R4194 VDD.n1137 VDD.n1136 9.3005
R4195 VDD.n639 VDD.n638 9.3005
R4196 VDD.n1489 VDD.n1488 9.3005
R4197 VDD.n783 VDD.n782 9.3005
R4198 VDD.n904 VDD.n903 9.3005
R4199 VDD.n905 VDD.n896 9.3005
R4200 VDD.n907 VDD.n906 9.3005
R4201 VDD.n908 VDD.n891 9.3005
R4202 VDD.n910 VDD.n909 9.3005
R4203 VDD.n911 VDD.n890 9.3005
R4204 VDD.n913 VDD.n912 9.3005
R4205 VDD.n914 VDD.n885 9.3005
R4206 VDD.n916 VDD.n915 9.3005
R4207 VDD.n917 VDD.n884 9.3005
R4208 VDD.n919 VDD.n918 9.3005
R4209 VDD.n920 VDD.n879 9.3005
R4210 VDD.n922 VDD.n921 9.3005
R4211 VDD.n923 VDD.n878 9.3005
R4212 VDD.n925 VDD.n924 9.3005
R4213 VDD.n926 VDD.n873 9.3005
R4214 VDD.n928 VDD.n927 9.3005
R4215 VDD.n929 VDD.n872 9.3005
R4216 VDD.n931 VDD.n930 9.3005
R4217 VDD.n935 VDD.n868 9.3005
R4218 VDD.n937 VDD.n936 9.3005
R4219 VDD.n938 VDD.n867 9.3005
R4220 VDD.n940 VDD.n939 9.3005
R4221 VDD.n941 VDD.n862 9.3005
R4222 VDD.n943 VDD.n942 9.3005
R4223 VDD.n944 VDD.n861 9.3005
R4224 VDD.n946 VDD.n945 9.3005
R4225 VDD.n947 VDD.n856 9.3005
R4226 VDD.n949 VDD.n948 9.3005
R4227 VDD.n950 VDD.n855 9.3005
R4228 VDD.n952 VDD.n951 9.3005
R4229 VDD.n953 VDD.n850 9.3005
R4230 VDD.n955 VDD.n954 9.3005
R4231 VDD.n956 VDD.n849 9.3005
R4232 VDD.n958 VDD.n957 9.3005
R4233 VDD.n959 VDD.n844 9.3005
R4234 VDD.n961 VDD.n960 9.3005
R4235 VDD.n962 VDD.n843 9.3005
R4236 VDD.n964 VDD.n963 9.3005
R4237 VDD.n968 VDD.n839 9.3005
R4238 VDD.n970 VDD.n969 9.3005
R4239 VDD.n971 VDD.n838 9.3005
R4240 VDD.n973 VDD.n972 9.3005
R4241 VDD.n974 VDD.n833 9.3005
R4242 VDD.n976 VDD.n975 9.3005
R4243 VDD.n977 VDD.n832 9.3005
R4244 VDD.n979 VDD.n978 9.3005
R4245 VDD.n980 VDD.n827 9.3005
R4246 VDD.n982 VDD.n981 9.3005
R4247 VDD.n983 VDD.n826 9.3005
R4248 VDD.n985 VDD.n984 9.3005
R4249 VDD.n986 VDD.n821 9.3005
R4250 VDD.n988 VDD.n987 9.3005
R4251 VDD.n989 VDD.n820 9.3005
R4252 VDD.n991 VDD.n990 9.3005
R4253 VDD.n789 VDD.n788 9.3005
R4254 VDD.n997 VDD.n996 9.3005
R4255 VDD.n899 VDD.n897 9.3005
R4256 VDD.n1000 VDD.n999 9.3005
R4257 VDD.n777 VDD.n776 9.3005
R4258 VDD.n1013 VDD.n1012 9.3005
R4259 VDD.n1014 VDD.n775 9.3005
R4260 VDD.n1016 VDD.n1015 9.3005
R4261 VDD.n765 VDD.n764 9.3005
R4262 VDD.n1029 VDD.n1028 9.3005
R4263 VDD.n1030 VDD.n763 9.3005
R4264 VDD.n1032 VDD.n1031 9.3005
R4265 VDD.n753 VDD.n752 9.3005
R4266 VDD.n1045 VDD.n1044 9.3005
R4267 VDD.n1046 VDD.n751 9.3005
R4268 VDD.n1048 VDD.n1047 9.3005
R4269 VDD.n741 VDD.n740 9.3005
R4270 VDD.n1061 VDD.n1060 9.3005
R4271 VDD.n1062 VDD.n739 9.3005
R4272 VDD.n1065 VDD.n1064 9.3005
R4273 VDD.n1063 VDD.n729 9.3005
R4274 VDD.n998 VDD.n787 9.3005
R4275 VDD.n1544 VDD.t188 8.95713
R4276 VDD.n1854 VDD.t105 8.95713
R4277 VDD.t102 VDD.n577 8.80785
R4278 VDD.n556 VDD.t14 8.80785
R4279 VDD.n1981 VDD.t9 8.80785
R4280 VDD.n2011 VDD.t107 8.80785
R4281 VDD.n15 VDD.n14 8.32723
R4282 VDD.n2529 VDD.n2528 8.07375
R4283 VDD.n728 VDD.n727 8.07375
R4284 VDD.n1556 VDD.t10 8.06147
R4285 VDD.t19 VDD.n405 8.06147
R4286 VDD.n773 VDD.t126 7.91219
R4287 VDD.n1123 VDD.t154 7.91219
R4288 VDD.n257 VDD.t128 7.91219
R4289 VDD.n2500 VDD.t110 7.91219
R4290 VDD.n749 VDD.t114 7.61364
R4291 VDD.n1091 VDD.t133 7.61364
R4292 VDD.n233 VDD.t150 7.61364
R4293 VDD.n2516 VDD.t112 7.61364
R4294 VDD.n1058 VDD.t114 7.31508
R4295 VDD.n695 VDD.t133 7.31508
R4296 VDD.n2338 VDD.t150 7.31508
R4297 VDD.t112 VDD.n55 7.31508
R4298 VDD.n1568 VDD.t97 7.1658
R4299 VDD.t1 VDD.n417 7.1658
R4300 VDD.n1026 VDD.t126 7.01653
R4301 VDD.n671 VDD.t154 7.01653
R4302 VDD.n2306 VDD.t128 7.01653
R4303 VDD.t110 VDD.n76 7.01653
R4304 VDD.n936 VDD.n935 6.98232
R4305 VDD.n1249 VDD.n1203 6.98232
R4306 VDD.n2418 VDD.n162 6.98232
R4307 VDD.n2203 VDD.n2200 6.98232
R4308 VDD.n34 VDD.n24 6.82916
R4309 VDD.n716 VDD.n706 6.82916
R4310 VDD.n1598 VDD.t194 6.5687
R4311 VDD.n1884 VDD.t190 6.5687
R4312 VDD.n7 VDD.t20 6.5015
R4313 VDD.n7 VDD.t106 6.5015
R4314 VDD.n8 VDD.t16 6.5015
R4315 VDD.n8 VDD.t2 6.5015
R4316 VDD.n10 VDD.t104 6.5015
R4317 VDD.n10 VDD.t191 6.5015
R4318 VDD.n12 VDD.t193 6.5015
R4319 VDD.n12 VDD.t4 6.5015
R4320 VDD.n5 VDD.t6 6.5015
R4321 VDD.n5 VDD.t13 6.5015
R4322 VDD.n3 VDD.t195 6.5015
R4323 VDD.n3 VDD.t100 6.5015
R4324 VDD.n1 VDD.t98 6.5015
R4325 VDD.n1 VDD.t8 6.5015
R4326 VDD.n0 VDD.t189 6.5015
R4327 VDD.n0 VDD.t11 6.5015
R4328 VDD.n1580 VDD.t7 6.27014
R4329 VDD.t15 VDD.n429 6.27014
R4330 VDD.n1699 VDD.n1698 6.0883
R4331 VDD.n1335 VDD.n1331 6.0883
R4332 VDD.n1909 VDD.n1908 6.0883
R4333 VDD.n390 VDD.n385 6.0883
R4334 VDD.n2132 VDD.n2131 6.0883
R4335 VDD.n1831 VDD.n1792 6.0883
R4336 VDD.n1638 VDD.n527 6.0883
R4337 VDD.n1367 VDD.n1366 6.0883
R4338 VDD.n1615 VDD.t99 5.67303
R4339 VDD.t103 VDD.n458 5.67303
R4340 VDD.n902 VDD.n899 5.62474
R4341 VDD.n1494 VDD.n1491 5.62474
R4342 VDD.n2381 VDD.n201 5.62474
R4343 VDD.n2161 VDD.n2158 5.62474
R4344 VDD.n1689 VDD.t5 5.37448
R4345 VDD.t12 VDD.n1738 5.37448
R4346 VDD.n1944 VDD.t192 5.37448
R4347 VDD.n1951 VDD.t3 5.37448
R4348 VDD.n521 VDD.t5 4.77737
R4349 VDD.t3 VDD.n470 4.77737
R4350 VDD.n1231 VDD.n626 4.74817
R4351 VDD.n1226 VDD.n627 4.74817
R4352 VDD.n1468 VDD.n1467 4.74817
R4353 VDD.n1301 VDD.n1158 4.74817
R4354 VDD.n1467 VDD.n1155 4.74817
R4355 VDD.n1301 VDD.n1300 4.74817
R4356 VDD.n2262 VDD.n2261 4.74817
R4357 VDD.n2259 VDD.n2258 4.74817
R4358 VDD.n2259 VDD.n314 4.74817
R4359 VDD.n2261 VDD.n309 4.74817
R4360 VDD.n2177 VDD.n349 4.74817
R4361 VDD.n2175 VDD.n2174 4.74817
R4362 VDD.n2175 VDD.n2150 4.74817
R4363 VDD.n2178 VDD.n2177 4.74817
R4364 VDD.n1223 VDD.n626 4.74817
R4365 VDD.n629 VDD.n627 4.74817
R4366 VDD.n44 VDD.n43 4.7074
R4367 VDD.n34 VDD.n33 4.7074
R4368 VDD.n726 VDD.n725 4.7074
R4369 VDD.n716 VDD.n715 4.7074
R4370 VDD.n41 VDD.t120 4.64407
R4371 VDD.n41 VDD.t153 4.64407
R4372 VDD.n39 VDD.t139 4.64407
R4373 VDD.n39 VDD.t159 4.64407
R4374 VDD.n37 VDD.t151 4.64407
R4375 VDD.n37 VDD.t181 4.64407
R4376 VDD.n35 VDD.t167 4.64407
R4377 VDD.n35 VDD.t117 4.64407
R4378 VDD.n31 VDD.t164 4.64407
R4379 VDD.n31 VDD.t186 4.64407
R4380 VDD.n29 VDD.t178 4.64407
R4381 VDD.n29 VDD.t137 4.64407
R4382 VDD.n27 VDD.t185 4.64407
R4383 VDD.n27 VDD.t143 4.64407
R4384 VDD.n25 VDD.t123 4.64407
R4385 VDD.n25 VDD.t163 4.64407
R4386 VDD.n22 VDD.t177 4.64407
R4387 VDD.n22 VDD.t166 4.64407
R4388 VDD.n20 VDD.t132 4.64407
R4389 VDD.n20 VDD.t113 4.64407
R4390 VDD.n18 VDD.t184 4.64407
R4391 VDD.n18 VDD.t173 4.64407
R4392 VDD.n16 VDD.t165 4.64407
R4393 VDD.n16 VDD.t118 4.64407
R4394 VDD.n717 VDD.t141 4.64407
R4395 VDD.n717 VDD.t183 4.64407
R4396 VDD.n719 VDD.t125 4.64407
R4397 VDD.n719 VDD.t172 4.64407
R4398 VDD.n721 VDD.t115 4.64407
R4399 VDD.n721 VDD.t157 4.64407
R4400 VDD.n723 VDD.t174 4.64407
R4401 VDD.n723 VDD.t146 4.64407
R4402 VDD.n707 VDD.t180 4.64407
R4403 VDD.n707 VDD.t149 4.64407
R4404 VDD.n709 VDD.t168 4.64407
R4405 VDD.n709 VDD.t134 4.64407
R4406 VDD.n711 VDD.t160 4.64407
R4407 VDD.n711 VDD.t109 4.64407
R4408 VDD.n713 VDD.t136 4.64407
R4409 VDD.n713 VDD.t182 4.64407
R4410 VDD.n698 VDD.t179 4.64407
R4411 VDD.n698 VDD.t148 4.64407
R4412 VDD.n700 VDD.t156 4.64407
R4413 VDD.n700 VDD.t169 4.64407
R4414 VDD.n702 VDD.t175 4.64407
R4415 VDD.n702 VDD.t138 4.64407
R4416 VDD.n704 VDD.t144 4.64407
R4417 VDD.n704 VDD.t161 4.64407
R4418 VDD.t33 VDD.n779 4.62809
R4419 VDD.n1139 VDD.t22 4.62809
R4420 VDD.t44 VDD.n263 4.62809
R4421 VDD.n2492 VDD.t51 4.62809
R4422 VDD.n1698 VDD.n1697 4.52733
R4423 VDD.n1446 VDD.n1335 4.52733
R4424 VDD.n1908 VDD.n1907 4.52733
R4425 VDD.n2080 VDD.n390 4.52733
R4426 VDD.n2131 VDD.n2130 4.52733
R4427 VDD.n1834 VDD.n1792 4.52733
R4428 VDD.n1635 VDD.n527 4.52733
R4429 VDD.n1368 VDD.n1367 4.52733
R4430 VDD.t99 VDD.n530 4.47882
R4431 VDD.n1963 VDD.t103 4.47882
R4432 VDD.n2529 VDD.n44 4.43518
R4433 VDD.n727 VDD.n726 4.43518
R4434 VDD.t26 VDD.n613 3.88171
R4435 VDD.n1414 VDD.t7 3.88171
R4436 VDD.n1993 VDD.t15 3.88171
R4437 VDD.n354 VDD.t82 3.88171
R4438 VDD.t194 VDD.n541 3.58315
R4439 VDD.n1975 VDD.t190 3.58315
R4440 VDD.t97 VDD.n571 2.98604
R4441 VDD.n2005 VDD.t1 2.98604
R4442 VDD.n1034 VDD.t135 2.83677
R4443 VDD.t147 VDD.n670 2.83677
R4444 VDD.n2314 VDD.t122 2.83677
R4445 VDD.t152 VDD.n2507 2.83677
R4446 VDD.n1067 VDD.t108 2.53821
R4447 VDD.t124 VDD.n694 2.53821
R4448 VDD.n2346 VDD.t142 2.53821
R4449 VDD.t131 VDD.n2523 2.53821
R4450 VDD.n1467 VDD.n1466 2.27742
R4451 VDD.n1466 VDD.n1301 2.27742
R4452 VDD.n2260 VDD.n2259 2.27742
R4453 VDD.n2261 VDD.n2260 2.27742
R4454 VDD.n2176 VDD.n2175 2.27742
R4455 VDD.n2177 VDD.n2176 2.27742
R4456 VDD.n1504 VDD.n626 2.27742
R4457 VDD.n1504 VDD.n627 2.27742
R4458 VDD.t145 VDD.n748 2.23966
R4459 VDD.n1099 VDD.t140 2.23966
R4460 VDD.t116 VDD.n232 2.23966
R4461 VDD.n2514 VDD.t119 2.23966
R4462 VDD.n44 VDD.n34 2.12227
R4463 VDD.n726 VDD.n716 2.12227
R4464 VDD.t10 VDD.n583 2.09038
R4465 VDD.n2017 VDD.t19 2.09038
R4466 VDD.n1562 VDD.t102 1.34399
R4467 VDD.n1598 VDD.t14 1.34399
R4468 VDD.n1884 VDD.t9 1.34399
R4469 VDD.t107 VDD.n411 1.34399
R4470 VDD.t188 VDD.n595 1.19472
R4471 VDD.n2063 VDD.t105 1.19472
R4472 VDD.n903 VDD.n902 0.970197
R4473 VDD.n1495 VDD.n1494 0.970197
R4474 VDD.n201 VDD.n197 0.970197
R4475 VDD.n2163 VDD.n2161 0.970197
R4476 VDD.n727 VDD.n15 0.87
R4477 VDD VDD.n2529 0.862167
R4478 VDD.n4 VDD.n2 0.728948
R4479 VDD.n11 VDD.n9 0.728948
R4480 VDD.n38 VDD.n36 0.573776
R4481 VDD.n40 VDD.n38 0.573776
R4482 VDD.n42 VDD.n40 0.573776
R4483 VDD.n43 VDD.n42 0.573776
R4484 VDD.n28 VDD.n26 0.573776
R4485 VDD.n30 VDD.n28 0.573776
R4486 VDD.n32 VDD.n30 0.573776
R4487 VDD.n33 VDD.n32 0.573776
R4488 VDD.n19 VDD.n17 0.573776
R4489 VDD.n21 VDD.n19 0.573776
R4490 VDD.n23 VDD.n21 0.573776
R4491 VDD.n24 VDD.n23 0.573776
R4492 VDD.n725 VDD.n724 0.573776
R4493 VDD.n724 VDD.n722 0.573776
R4494 VDD.n722 VDD.n720 0.573776
R4495 VDD.n720 VDD.n718 0.573776
R4496 VDD.n715 VDD.n714 0.573776
R4497 VDD.n714 VDD.n712 0.573776
R4498 VDD.n712 VDD.n710 0.573776
R4499 VDD.n710 VDD.n708 0.573776
R4500 VDD.n706 VDD.n705 0.573776
R4501 VDD.n705 VDD.n703 0.573776
R4502 VDD.n703 VDD.n701 0.573776
R4503 VDD.n701 VDD.n699 0.573776
R4504 VDD.n6 VDD.n4 0.573776
R4505 VDD.n13 VDD.n11 0.573776
R4506 VDD.n14 VDD.n6 0.49619
R4507 VDD.n14 VDD.n13 0.49619
R4508 VDD.n1483 VDD.n1482 0.471537
R4509 VDD.n2278 VDD.n2277 0.471537
R4510 VDD.n2487 VDD.n2486 0.471537
R4511 VDD.n2380 VDD.n2379 0.471537
R4512 VDD.n2157 VDD.n266 0.471537
R4513 VDD.n1490 VDD.n1489 0.471537
R4514 VDD.n897 VDD.n782 0.471537
R4515 VDD.n998 VDD.n997 0.471537
R4516 VDD.n1574 VDD.t0 0.448332
R4517 VDD.n1586 VDD.t17 0.448332
R4518 VDD.n443 VDD.t101 0.448332
R4519 VDD.t18 VDD.n423 0.448332
R4520 VDD.n1079 VDD.n1078 0.152939
R4521 VDD.n1080 VDD.n1079 0.152939
R4522 VDD.n1080 VDD.n686 0.152939
R4523 VDD.n1094 VDD.n686 0.152939
R4524 VDD.n1095 VDD.n1094 0.152939
R4525 VDD.n1096 VDD.n1095 0.152939
R4526 VDD.n1096 VDD.n674 0.152939
R4527 VDD.n1110 VDD.n674 0.152939
R4528 VDD.n1111 VDD.n1110 0.152939
R4529 VDD.n1112 VDD.n1111 0.152939
R4530 VDD.n1112 VDD.n662 0.152939
R4531 VDD.n1126 VDD.n662 0.152939
R4532 VDD.n1127 VDD.n1126 0.152939
R4533 VDD.n1128 VDD.n1127 0.152939
R4534 VDD.n1128 VDD.n650 0.152939
R4535 VDD.n1142 VDD.n650 0.152939
R4536 VDD.n1143 VDD.n1142 0.152939
R4537 VDD.n1483 VDD.n1143 0.152939
R4538 VDD.n1482 VDD.n1144 0.152939
R4539 VDD.n1148 VDD.n1144 0.152939
R4540 VDD.n1149 VDD.n1148 0.152939
R4541 VDD.n1150 VDD.n1149 0.152939
R4542 VDD.n1151 VDD.n1150 0.152939
R4543 VDD.n1156 VDD.n1151 0.152939
R4544 VDD.n1164 VDD.n1157 0.152939
R4545 VDD.n1165 VDD.n1164 0.152939
R4546 VDD.n1166 VDD.n1165 0.152939
R4547 VDD.n1167 VDD.n1166 0.152939
R4548 VDD.n1174 VDD.n1167 0.152939
R4549 VDD.n1285 VDD.n1174 0.152939
R4550 VDD.n1285 VDD.n1284 0.152939
R4551 VDD.n1284 VDD.n1283 0.152939
R4552 VDD.n1283 VDD.n1175 0.152939
R4553 VDD.n1179 VDD.n1175 0.152939
R4554 VDD.n1180 VDD.n1179 0.152939
R4555 VDD.n1181 VDD.n1180 0.152939
R4556 VDD.n1185 VDD.n1181 0.152939
R4557 VDD.n1186 VDD.n1185 0.152939
R4558 VDD.n1187 VDD.n1186 0.152939
R4559 VDD.n1188 VDD.n1187 0.152939
R4560 VDD.n1192 VDD.n1188 0.152939
R4561 VDD.n1193 VDD.n1192 0.152939
R4562 VDD.n1194 VDD.n1193 0.152939
R4563 VDD.n1195 VDD.n1194 0.152939
R4564 VDD.n1199 VDD.n1195 0.152939
R4565 VDD.n1200 VDD.n1199 0.152939
R4566 VDD.n1201 VDD.n1200 0.152939
R4567 VDD.n1202 VDD.n1201 0.152939
R4568 VDD.n1209 VDD.n1202 0.152939
R4569 VDD.n1248 VDD.n1209 0.152939
R4570 VDD.n1248 VDD.n1247 0.152939
R4571 VDD.n1247 VDD.n1246 0.152939
R4572 VDD.n1246 VDD.n1210 0.152939
R4573 VDD.n1214 VDD.n1210 0.152939
R4574 VDD.n1215 VDD.n1214 0.152939
R4575 VDD.n1216 VDD.n1215 0.152939
R4576 VDD.n1220 VDD.n1216 0.152939
R4577 VDD.n1221 VDD.n1220 0.152939
R4578 VDD.n1221 VDD.n625 0.152939
R4579 VDD.n316 VDD.n310 0.152939
R4580 VDD.n317 VDD.n316 0.152939
R4581 VDD.n318 VDD.n317 0.152939
R4582 VDD.n319 VDD.n318 0.152939
R4583 VDD.n320 VDD.n319 0.152939
R4584 VDD.n2241 VDD.n320 0.152939
R4585 VDD.n2241 VDD.n2240 0.152939
R4586 VDD.n2240 VDD.n2239 0.152939
R4587 VDD.n2239 VDD.n322 0.152939
R4588 VDD.n323 VDD.n322 0.152939
R4589 VDD.n324 VDD.n323 0.152939
R4590 VDD.n325 VDD.n324 0.152939
R4591 VDD.n326 VDD.n325 0.152939
R4592 VDD.n327 VDD.n326 0.152939
R4593 VDD.n328 VDD.n327 0.152939
R4594 VDD.n329 VDD.n328 0.152939
R4595 VDD.n330 VDD.n329 0.152939
R4596 VDD.n331 VDD.n330 0.152939
R4597 VDD.n332 VDD.n331 0.152939
R4598 VDD.n333 VDD.n332 0.152939
R4599 VDD.n334 VDD.n333 0.152939
R4600 VDD.n335 VDD.n334 0.152939
R4601 VDD.n336 VDD.n335 0.152939
R4602 VDD.n337 VDD.n336 0.152939
R4603 VDD.n338 VDD.n337 0.152939
R4604 VDD.n2199 VDD.n338 0.152939
R4605 VDD.n2199 VDD.n2198 0.152939
R4606 VDD.n2198 VDD.n2197 0.152939
R4607 VDD.n2197 VDD.n342 0.152939
R4608 VDD.n343 VDD.n342 0.152939
R4609 VDD.n344 VDD.n343 0.152939
R4610 VDD.n345 VDD.n344 0.152939
R4611 VDD.n346 VDD.n345 0.152939
R4612 VDD.n347 VDD.n346 0.152939
R4613 VDD.n348 VDD.n347 0.152939
R4614 VDD.n2277 VDD.n272 0.152939
R4615 VDD.n304 VDD.n272 0.152939
R4616 VDD.n305 VDD.n304 0.152939
R4617 VDD.n306 VDD.n305 0.152939
R4618 VDD.n307 VDD.n306 0.152939
R4619 VDD.n308 VDD.n307 0.152939
R4620 VDD.n2279 VDD.n2278 0.152939
R4621 VDD.n2279 VDD.n260 0.152939
R4622 VDD.n2293 VDD.n260 0.152939
R4623 VDD.n2294 VDD.n2293 0.152939
R4624 VDD.n2295 VDD.n2294 0.152939
R4625 VDD.n2295 VDD.n248 0.152939
R4626 VDD.n2309 VDD.n248 0.152939
R4627 VDD.n2310 VDD.n2309 0.152939
R4628 VDD.n2311 VDD.n2310 0.152939
R4629 VDD.n2311 VDD.n236 0.152939
R4630 VDD.n2325 VDD.n236 0.152939
R4631 VDD.n2326 VDD.n2325 0.152939
R4632 VDD.n2327 VDD.n2326 0.152939
R4633 VDD.n2327 VDD.n224 0.152939
R4634 VDD.n2341 VDD.n224 0.152939
R4635 VDD.n2342 VDD.n2341 0.152939
R4636 VDD.n2343 VDD.n2342 0.152939
R4637 VDD.n2343 VDD.n45 0.152939
R4638 VDD.n2527 VDD.n46 0.152939
R4639 VDD.n57 VDD.n46 0.152939
R4640 VDD.n58 VDD.n57 0.152939
R4641 VDD.n59 VDD.n58 0.152939
R4642 VDD.n66 VDD.n59 0.152939
R4643 VDD.n67 VDD.n66 0.152939
R4644 VDD.n68 VDD.n67 0.152939
R4645 VDD.n69 VDD.n68 0.152939
R4646 VDD.n78 VDD.n69 0.152939
R4647 VDD.n79 VDD.n78 0.152939
R4648 VDD.n80 VDD.n79 0.152939
R4649 VDD.n81 VDD.n80 0.152939
R4650 VDD.n89 VDD.n81 0.152939
R4651 VDD.n90 VDD.n89 0.152939
R4652 VDD.n91 VDD.n90 0.152939
R4653 VDD.n92 VDD.n91 0.152939
R4654 VDD.n100 VDD.n92 0.152939
R4655 VDD.n2487 VDD.n100 0.152939
R4656 VDD.n2486 VDD.n101 0.152939
R4657 VDD.n104 VDD.n101 0.152939
R4658 VDD.n108 VDD.n104 0.152939
R4659 VDD.n109 VDD.n108 0.152939
R4660 VDD.n110 VDD.n109 0.152939
R4661 VDD.n111 VDD.n110 0.152939
R4662 VDD.n112 VDD.n111 0.152939
R4663 VDD.n116 VDD.n112 0.152939
R4664 VDD.n117 VDD.n116 0.152939
R4665 VDD.n118 VDD.n117 0.152939
R4666 VDD.n119 VDD.n118 0.152939
R4667 VDD.n123 VDD.n119 0.152939
R4668 VDD.n124 VDD.n123 0.152939
R4669 VDD.n125 VDD.n124 0.152939
R4670 VDD.n126 VDD.n125 0.152939
R4671 VDD.n133 VDD.n126 0.152939
R4672 VDD.n2454 VDD.n133 0.152939
R4673 VDD.n2454 VDD.n2453 0.152939
R4674 VDD.n2453 VDD.n2452 0.152939
R4675 VDD.n2452 VDD.n134 0.152939
R4676 VDD.n138 VDD.n134 0.152939
R4677 VDD.n139 VDD.n138 0.152939
R4678 VDD.n140 VDD.n139 0.152939
R4679 VDD.n144 VDD.n140 0.152939
R4680 VDD.n145 VDD.n144 0.152939
R4681 VDD.n146 VDD.n145 0.152939
R4682 VDD.n147 VDD.n146 0.152939
R4683 VDD.n151 VDD.n147 0.152939
R4684 VDD.n152 VDD.n151 0.152939
R4685 VDD.n153 VDD.n152 0.152939
R4686 VDD.n154 VDD.n153 0.152939
R4687 VDD.n158 VDD.n154 0.152939
R4688 VDD.n159 VDD.n158 0.152939
R4689 VDD.n160 VDD.n159 0.152939
R4690 VDD.n161 VDD.n160 0.152939
R4691 VDD.n168 VDD.n161 0.152939
R4692 VDD.n2417 VDD.n168 0.152939
R4693 VDD.n2417 VDD.n2416 0.152939
R4694 VDD.n2416 VDD.n2415 0.152939
R4695 VDD.n2415 VDD.n169 0.152939
R4696 VDD.n173 VDD.n169 0.152939
R4697 VDD.n174 VDD.n173 0.152939
R4698 VDD.n175 VDD.n174 0.152939
R4699 VDD.n179 VDD.n175 0.152939
R4700 VDD.n180 VDD.n179 0.152939
R4701 VDD.n181 VDD.n180 0.152939
R4702 VDD.n182 VDD.n181 0.152939
R4703 VDD.n186 VDD.n182 0.152939
R4704 VDD.n187 VDD.n186 0.152939
R4705 VDD.n188 VDD.n187 0.152939
R4706 VDD.n189 VDD.n188 0.152939
R4707 VDD.n193 VDD.n189 0.152939
R4708 VDD.n194 VDD.n193 0.152939
R4709 VDD.n195 VDD.n194 0.152939
R4710 VDD.n196 VDD.n195 0.152939
R4711 VDD.n202 VDD.n196 0.152939
R4712 VDD.n2380 VDD.n202 0.152939
R4713 VDD.n2285 VDD.n266 0.152939
R4714 VDD.n2286 VDD.n2285 0.152939
R4715 VDD.n2287 VDD.n2286 0.152939
R4716 VDD.n2287 VDD.n253 0.152939
R4717 VDD.n2301 VDD.n253 0.152939
R4718 VDD.n2302 VDD.n2301 0.152939
R4719 VDD.n2303 VDD.n2302 0.152939
R4720 VDD.n2303 VDD.n242 0.152939
R4721 VDD.n2317 VDD.n242 0.152939
R4722 VDD.n2318 VDD.n2317 0.152939
R4723 VDD.n2319 VDD.n2318 0.152939
R4724 VDD.n2319 VDD.n229 0.152939
R4725 VDD.n2333 VDD.n229 0.152939
R4726 VDD.n2334 VDD.n2333 0.152939
R4727 VDD.n2335 VDD.n2334 0.152939
R4728 VDD.n2335 VDD.n217 0.152939
R4729 VDD.n2349 VDD.n217 0.152939
R4730 VDD.n2350 VDD.n2349 0.152939
R4731 VDD.n2351 VDD.n2350 0.152939
R4732 VDD.n2351 VDD.n215 0.152939
R4733 VDD.n2355 VDD.n215 0.152939
R4734 VDD.n2356 VDD.n2355 0.152939
R4735 VDD.n2357 VDD.n2356 0.152939
R4736 VDD.n2357 VDD.n212 0.152939
R4737 VDD.n2361 VDD.n212 0.152939
R4738 VDD.n2362 VDD.n2361 0.152939
R4739 VDD.n2363 VDD.n2362 0.152939
R4740 VDD.n2363 VDD.n209 0.152939
R4741 VDD.n2367 VDD.n209 0.152939
R4742 VDD.n2368 VDD.n2367 0.152939
R4743 VDD.n2369 VDD.n2368 0.152939
R4744 VDD.n2369 VDD.n206 0.152939
R4745 VDD.n2373 VDD.n206 0.152939
R4746 VDD.n2374 VDD.n2373 0.152939
R4747 VDD.n2375 VDD.n2374 0.152939
R4748 VDD.n2375 VDD.n203 0.152939
R4749 VDD.n2379 VDD.n203 0.152939
R4750 VDD.n2152 VDD.n350 0.152939
R4751 VDD.n2153 VDD.n2152 0.152939
R4752 VDD.n2154 VDD.n2153 0.152939
R4753 VDD.n2155 VDD.n2154 0.152939
R4754 VDD.n2156 VDD.n2155 0.152939
R4755 VDD.n2157 VDD.n2156 0.152939
R4756 VDD.n1503 VDD.n628 0.152939
R4757 VDD.n1499 VDD.n628 0.152939
R4758 VDD.n1499 VDD.n1498 0.152939
R4759 VDD.n1498 VDD.n1497 0.152939
R4760 VDD.n1497 VDD.n634 0.152939
R4761 VDD.n1490 VDD.n634 0.152939
R4762 VDD.n1005 VDD.n782 0.152939
R4763 VDD.n1006 VDD.n1005 0.152939
R4764 VDD.n1007 VDD.n1006 0.152939
R4765 VDD.n1007 VDD.n769 0.152939
R4766 VDD.n1021 VDD.n769 0.152939
R4767 VDD.n1022 VDD.n1021 0.152939
R4768 VDD.n1023 VDD.n1022 0.152939
R4769 VDD.n1023 VDD.n758 0.152939
R4770 VDD.n1037 VDD.n758 0.152939
R4771 VDD.n1038 VDD.n1037 0.152939
R4772 VDD.n1039 VDD.n1038 0.152939
R4773 VDD.n1039 VDD.n745 0.152939
R4774 VDD.n1053 VDD.n745 0.152939
R4775 VDD.n1054 VDD.n1053 0.152939
R4776 VDD.n1055 VDD.n1054 0.152939
R4777 VDD.n1055 VDD.n734 0.152939
R4778 VDD.n1070 VDD.n734 0.152939
R4779 VDD.n1071 VDD.n1070 0.152939
R4780 VDD.n1072 VDD.n1071 0.152939
R4781 VDD.n1072 VDD.n691 0.152939
R4782 VDD.n1086 VDD.n691 0.152939
R4783 VDD.n1087 VDD.n1086 0.152939
R4784 VDD.n1088 VDD.n1087 0.152939
R4785 VDD.n1088 VDD.n680 0.152939
R4786 VDD.n1102 VDD.n680 0.152939
R4787 VDD.n1103 VDD.n1102 0.152939
R4788 VDD.n1104 VDD.n1103 0.152939
R4789 VDD.n1104 VDD.n667 0.152939
R4790 VDD.n1118 VDD.n667 0.152939
R4791 VDD.n1119 VDD.n1118 0.152939
R4792 VDD.n1120 VDD.n1119 0.152939
R4793 VDD.n1120 VDD.n656 0.152939
R4794 VDD.n1134 VDD.n656 0.152939
R4795 VDD.n1135 VDD.n1134 0.152939
R4796 VDD.n1136 VDD.n1135 0.152939
R4797 VDD.n1136 VDD.n638 0.152939
R4798 VDD.n1489 VDD.n638 0.152939
R4799 VDD.n997 VDD.n788 0.152939
R4800 VDD.n990 VDD.n788 0.152939
R4801 VDD.n990 VDD.n989 0.152939
R4802 VDD.n989 VDD.n988 0.152939
R4803 VDD.n988 VDD.n821 0.152939
R4804 VDD.n984 VDD.n821 0.152939
R4805 VDD.n984 VDD.n983 0.152939
R4806 VDD.n983 VDD.n982 0.152939
R4807 VDD.n982 VDD.n827 0.152939
R4808 VDD.n978 VDD.n827 0.152939
R4809 VDD.n978 VDD.n977 0.152939
R4810 VDD.n977 VDD.n976 0.152939
R4811 VDD.n976 VDD.n833 0.152939
R4812 VDD.n972 VDD.n833 0.152939
R4813 VDD.n972 VDD.n971 0.152939
R4814 VDD.n971 VDD.n970 0.152939
R4815 VDD.n970 VDD.n839 0.152939
R4816 VDD.n963 VDD.n839 0.152939
R4817 VDD.n963 VDD.n962 0.152939
R4818 VDD.n962 VDD.n961 0.152939
R4819 VDD.n961 VDD.n844 0.152939
R4820 VDD.n957 VDD.n844 0.152939
R4821 VDD.n957 VDD.n956 0.152939
R4822 VDD.n956 VDD.n955 0.152939
R4823 VDD.n955 VDD.n850 0.152939
R4824 VDD.n951 VDD.n850 0.152939
R4825 VDD.n951 VDD.n950 0.152939
R4826 VDD.n950 VDD.n949 0.152939
R4827 VDD.n949 VDD.n856 0.152939
R4828 VDD.n945 VDD.n856 0.152939
R4829 VDD.n945 VDD.n944 0.152939
R4830 VDD.n944 VDD.n943 0.152939
R4831 VDD.n943 VDD.n862 0.152939
R4832 VDD.n939 VDD.n862 0.152939
R4833 VDD.n939 VDD.n938 0.152939
R4834 VDD.n938 VDD.n937 0.152939
R4835 VDD.n937 VDD.n868 0.152939
R4836 VDD.n930 VDD.n868 0.152939
R4837 VDD.n930 VDD.n929 0.152939
R4838 VDD.n929 VDD.n928 0.152939
R4839 VDD.n928 VDD.n873 0.152939
R4840 VDD.n924 VDD.n873 0.152939
R4841 VDD.n924 VDD.n923 0.152939
R4842 VDD.n923 VDD.n922 0.152939
R4843 VDD.n922 VDD.n879 0.152939
R4844 VDD.n918 VDD.n879 0.152939
R4845 VDD.n918 VDD.n917 0.152939
R4846 VDD.n917 VDD.n916 0.152939
R4847 VDD.n916 VDD.n885 0.152939
R4848 VDD.n912 VDD.n885 0.152939
R4849 VDD.n912 VDD.n911 0.152939
R4850 VDD.n911 VDD.n910 0.152939
R4851 VDD.n910 VDD.n891 0.152939
R4852 VDD.n906 VDD.n891 0.152939
R4853 VDD.n906 VDD.n905 0.152939
R4854 VDD.n905 VDD.n904 0.152939
R4855 VDD.n904 VDD.n897 0.152939
R4856 VDD.n999 VDD.n998 0.152939
R4857 VDD.n999 VDD.n776 0.152939
R4858 VDD.n1013 VDD.n776 0.152939
R4859 VDD.n1014 VDD.n1013 0.152939
R4860 VDD.n1015 VDD.n1014 0.152939
R4861 VDD.n1015 VDD.n764 0.152939
R4862 VDD.n1029 VDD.n764 0.152939
R4863 VDD.n1030 VDD.n1029 0.152939
R4864 VDD.n1031 VDD.n1030 0.152939
R4865 VDD.n1031 VDD.n752 0.152939
R4866 VDD.n1045 VDD.n752 0.152939
R4867 VDD.n1046 VDD.n1045 0.152939
R4868 VDD.n1047 VDD.n1046 0.152939
R4869 VDD.n1047 VDD.n740 0.152939
R4870 VDD.n1061 VDD.n740 0.152939
R4871 VDD.n1062 VDD.n1061 0.152939
R4872 VDD.n1064 VDD.n1062 0.152939
R4873 VDD.n1064 VDD.n1063 0.152939
R4874 VDD.n609 VDD.t71 0.149777
R4875 VDD.n1683 VDD.t64 0.149777
R4876 VDD.n1957 VDD.t78 0.149777
R4877 VDD.n2069 VDD.t37 0.149777
R4878 VDD.n1466 VDD.n1156 0.110256
R4879 VDD.n2260 VDD.n308 0.110256
R4880 VDD.n2176 VDD.n350 0.110256
R4881 VDD.n1504 VDD.n1503 0.110256
R4882 VDD.n1078 VDD.n728 0.0695946
R4883 VDD.n2528 VDD.n45 0.0695946
R4884 VDD.n2528 VDD.n2527 0.0695946
R4885 VDD.n1063 VDD.n728 0.0695946
R4886 VDD.n1466 VDD.n1157 0.0431829
R4887 VDD.n1504 VDD.n625 0.0431829
R4888 VDD.n2260 VDD.n310 0.0431829
R4889 VDD.n2176 VDD.n348 0.0431829
R4890 VDD VDD.n15 0.00833333
R4891 VOUT.n202 VOUT.n200 102.66
R4892 VOUT.n192 VOUT.n190 102.66
R4893 VOUT.n183 VOUT.n181 102.66
R4894 VOUT.n21 VOUT.n19 102.66
R4895 VOUT.n11 VOUT.n9 102.66
R4896 VOUT.n2 VOUT.n0 102.66
R4897 VOUT.n206 VOUT.n205 102.088
R4898 VOUT.n204 VOUT.n203 102.088
R4899 VOUT.n202 VOUT.n201 102.088
R4900 VOUT.n198 VOUT.n197 102.088
R4901 VOUT.n196 VOUT.n195 102.088
R4902 VOUT.n194 VOUT.n193 102.088
R4903 VOUT.n192 VOUT.n191 102.088
R4904 VOUT.n189 VOUT.n188 102.088
R4905 VOUT.n187 VOUT.n186 102.088
R4906 VOUT.n185 VOUT.n184 102.088
R4907 VOUT.n183 VOUT.n182 102.088
R4908 VOUT.n21 VOUT.n20 102.088
R4909 VOUT.n23 VOUT.n22 102.088
R4910 VOUT.n25 VOUT.n24 102.088
R4911 VOUT.n27 VOUT.n26 102.088
R4912 VOUT.n11 VOUT.n10 102.088
R4913 VOUT.n13 VOUT.n12 102.088
R4914 VOUT.n15 VOUT.n14 102.088
R4915 VOUT.n17 VOUT.n16 102.088
R4916 VOUT.n2 VOUT.n1 102.088
R4917 VOUT.n4 VOUT.n3 102.088
R4918 VOUT.n6 VOUT.n5 102.088
R4919 VOUT.n8 VOUT.n7 102.088
R4920 VOUT.n208 VOUT.n207 102.088
R4921 VOUT.n220 VOUT.n218 85.0679
R4922 VOUT.n213 VOUT.n211 85.0679
R4923 VOUT.n236 VOUT.n234 85.0679
R4924 VOUT.n229 VOUT.n227 85.0679
R4925 VOUT.n224 VOUT.n223 84.0635
R4926 VOUT.n222 VOUT.n221 84.0635
R4927 VOUT.n220 VOUT.n219 84.0635
R4928 VOUT.n217 VOUT.n216 84.0635
R4929 VOUT.n215 VOUT.n214 84.0635
R4930 VOUT.n213 VOUT.n212 84.0635
R4931 VOUT.n236 VOUT.n235 84.0635
R4932 VOUT.n238 VOUT.n237 84.0635
R4933 VOUT.n240 VOUT.n239 84.0635
R4934 VOUT.n229 VOUT.n228 84.0635
R4935 VOUT.n231 VOUT.n230 84.0635
R4936 VOUT.n233 VOUT.n232 84.0635
R4937 VOUT.n226 VOUT.n210 8.52206
R4938 VOUT.n199 VOUT.n189 7.37442
R4939 VOUT.n18 VOUT.n8 7.37442
R4940 VOUT.n225 VOUT.n217 7.37334
R4941 VOUT.n241 VOUT.n233 7.37334
R4942 VOUT.n226 VOUT.n225 5.98809
R4943 VOUT.n242 VOUT.n241 5.98809
R4944 VOUT.n225 VOUT.n224 5.46817
R4945 VOUT.n241 VOUT.n240 5.46817
R4946 VOUT.n209 VOUT.n208 5.25266
R4947 VOUT.n199 VOUT.n198 5.25266
R4948 VOUT.n28 VOUT.n27 5.25266
R4949 VOUT.n18 VOUT.n17 5.25266
R4950 VOUT.n243 VOUT.n29 4.9022
R4951 VOUT.n210 VOUT.n209 4.78873
R4952 VOUT.n29 VOUT.n28 4.78873
R4953 VOUT.n207 VOUT.t51 4.64407
R4954 VOUT.n207 VOUT.t26 4.64407
R4955 VOUT.n205 VOUT.t71 4.64407
R4956 VOUT.n205 VOUT.t32 4.64407
R4957 VOUT.n203 VOUT.t78 4.64407
R4958 VOUT.n203 VOUT.t43 4.64407
R4959 VOUT.n201 VOUT.t29 4.64407
R4960 VOUT.n201 VOUT.t50 4.64407
R4961 VOUT.n200 VOUT.t36 4.64407
R4962 VOUT.n200 VOUT.t62 4.64407
R4963 VOUT.n197 VOUT.t83 4.64407
R4964 VOUT.n197 VOUT.t55 4.64407
R4965 VOUT.n195 VOUT.t41 4.64407
R4966 VOUT.n195 VOUT.t60 4.64407
R4967 VOUT.n193 VOUT.t45 4.64407
R4968 VOUT.n193 VOUT.t75 4.64407
R4969 VOUT.n191 VOUT.t59 4.64407
R4970 VOUT.n191 VOUT.t82 4.64407
R4971 VOUT.n190 VOUT.t67 4.64407
R4972 VOUT.n190 VOUT.t33 4.64407
R4973 VOUT.n188 VOUT.t61 4.64407
R4974 VOUT.n188 VOUT.t31 4.64407
R4975 VOUT.n186 VOUT.t27 4.64407
R4976 VOUT.n186 VOUT.t74 4.64407
R4977 VOUT.n184 VOUT.t69 4.64407
R4978 VOUT.n184 VOUT.t37 4.64407
R4979 VOUT.n182 VOUT.t30 4.64407
R4980 VOUT.n182 VOUT.t81 4.64407
R4981 VOUT.n181 VOUT.t73 4.64407
R4982 VOUT.n181 VOUT.t63 4.64407
R4983 VOUT.n19 VOUT.t80 4.64407
R4984 VOUT.n19 VOUT.t52 4.64407
R4985 VOUT.n20 VOUT.t68 4.64407
R4986 VOUT.n20 VOUT.t44 4.64407
R4987 VOUT.n22 VOUT.t54 4.64407
R4988 VOUT.n22 VOUT.t34 4.64407
R4989 VOUT.n24 VOUT.t46 4.64407
R4990 VOUT.n24 VOUT.t28 4.64407
R4991 VOUT.n26 VOUT.t35 4.64407
R4992 VOUT.n26 VOUT.t70 4.64407
R4993 VOUT.n9 VOUT.t49 4.64407
R4994 VOUT.n9 VOUT.t84 4.64407
R4995 VOUT.n10 VOUT.t39 4.64407
R4996 VOUT.n10 VOUT.t77 4.64407
R4997 VOUT.n12 VOUT.t25 4.64407
R4998 VOUT.n12 VOUT.t64 4.64407
R4999 VOUT.n14 VOUT.t79 4.64407
R5000 VOUT.n14 VOUT.t56 4.64407
R5001 VOUT.n16 VOUT.t66 4.64407
R5002 VOUT.n16 VOUT.t40 4.64407
R5003 VOUT.n0 VOUT.t48 4.64407
R5004 VOUT.n0 VOUT.t58 4.64407
R5005 VOUT.n1 VOUT.t65 4.64407
R5006 VOUT.n1 VOUT.t76 4.64407
R5007 VOUT.n3 VOUT.t42 4.64407
R5008 VOUT.n3 VOUT.t53 4.64407
R5009 VOUT.n5 VOUT.t57 4.64407
R5010 VOUT.n5 VOUT.t72 4.64407
R5011 VOUT.n7 VOUT.t38 4.64407
R5012 VOUT.n7 VOUT.t47 4.64407
R5013 VOUT.n120 VOUT.n73 4.5005
R5014 VOUT.n89 VOUT.n73 4.5005
R5015 VOUT.n84 VOUT.n68 4.5005
R5016 VOUT.n84 VOUT.n70 4.5005
R5017 VOUT.n84 VOUT.n67 4.5005
R5018 VOUT.n84 VOUT.n71 4.5005
R5019 VOUT.n84 VOUT.n66 4.5005
R5020 VOUT.n84 VOUT.t94 4.5005
R5021 VOUT.n84 VOUT.n65 4.5005
R5022 VOUT.n84 VOUT.n72 4.5005
R5023 VOUT.n84 VOUT.n73 4.5005
R5024 VOUT.n82 VOUT.n68 4.5005
R5025 VOUT.n82 VOUT.n70 4.5005
R5026 VOUT.n82 VOUT.n67 4.5005
R5027 VOUT.n82 VOUT.n71 4.5005
R5028 VOUT.n82 VOUT.n66 4.5005
R5029 VOUT.n82 VOUT.t94 4.5005
R5030 VOUT.n82 VOUT.n65 4.5005
R5031 VOUT.n82 VOUT.n72 4.5005
R5032 VOUT.n82 VOUT.n73 4.5005
R5033 VOUT.n81 VOUT.n68 4.5005
R5034 VOUT.n81 VOUT.n70 4.5005
R5035 VOUT.n81 VOUT.n67 4.5005
R5036 VOUT.n81 VOUT.n71 4.5005
R5037 VOUT.n81 VOUT.n66 4.5005
R5038 VOUT.n81 VOUT.t94 4.5005
R5039 VOUT.n81 VOUT.n65 4.5005
R5040 VOUT.n81 VOUT.n72 4.5005
R5041 VOUT.n81 VOUT.n73 4.5005
R5042 VOUT.n166 VOUT.n68 4.5005
R5043 VOUT.n166 VOUT.n70 4.5005
R5044 VOUT.n166 VOUT.n67 4.5005
R5045 VOUT.n166 VOUT.n71 4.5005
R5046 VOUT.n166 VOUT.n66 4.5005
R5047 VOUT.n166 VOUT.t94 4.5005
R5048 VOUT.n166 VOUT.n65 4.5005
R5049 VOUT.n166 VOUT.n72 4.5005
R5050 VOUT.n166 VOUT.n73 4.5005
R5051 VOUT.n164 VOUT.n68 4.5005
R5052 VOUT.n164 VOUT.n70 4.5005
R5053 VOUT.n164 VOUT.n67 4.5005
R5054 VOUT.n164 VOUT.n71 4.5005
R5055 VOUT.n164 VOUT.n66 4.5005
R5056 VOUT.n164 VOUT.t94 4.5005
R5057 VOUT.n164 VOUT.n65 4.5005
R5058 VOUT.n164 VOUT.n72 4.5005
R5059 VOUT.n162 VOUT.n68 4.5005
R5060 VOUT.n162 VOUT.n70 4.5005
R5061 VOUT.n162 VOUT.n67 4.5005
R5062 VOUT.n162 VOUT.n71 4.5005
R5063 VOUT.n162 VOUT.n66 4.5005
R5064 VOUT.n162 VOUT.t94 4.5005
R5065 VOUT.n162 VOUT.n65 4.5005
R5066 VOUT.n162 VOUT.n72 4.5005
R5067 VOUT.n92 VOUT.n68 4.5005
R5068 VOUT.n92 VOUT.n70 4.5005
R5069 VOUT.n92 VOUT.n67 4.5005
R5070 VOUT.n92 VOUT.n71 4.5005
R5071 VOUT.n92 VOUT.n66 4.5005
R5072 VOUT.n92 VOUT.t94 4.5005
R5073 VOUT.n92 VOUT.n65 4.5005
R5074 VOUT.n92 VOUT.n72 4.5005
R5075 VOUT.n92 VOUT.n73 4.5005
R5076 VOUT.n91 VOUT.n68 4.5005
R5077 VOUT.n91 VOUT.n70 4.5005
R5078 VOUT.n91 VOUT.n67 4.5005
R5079 VOUT.n91 VOUT.n71 4.5005
R5080 VOUT.n91 VOUT.n66 4.5005
R5081 VOUT.n91 VOUT.t94 4.5005
R5082 VOUT.n91 VOUT.n65 4.5005
R5083 VOUT.n91 VOUT.n72 4.5005
R5084 VOUT.n91 VOUT.n73 4.5005
R5085 VOUT.n95 VOUT.n68 4.5005
R5086 VOUT.n95 VOUT.n70 4.5005
R5087 VOUT.n95 VOUT.n67 4.5005
R5088 VOUT.n95 VOUT.n71 4.5005
R5089 VOUT.n95 VOUT.n66 4.5005
R5090 VOUT.n95 VOUT.t94 4.5005
R5091 VOUT.n95 VOUT.n65 4.5005
R5092 VOUT.n95 VOUT.n72 4.5005
R5093 VOUT.n95 VOUT.n73 4.5005
R5094 VOUT.n94 VOUT.n68 4.5005
R5095 VOUT.n94 VOUT.n70 4.5005
R5096 VOUT.n94 VOUT.n67 4.5005
R5097 VOUT.n94 VOUT.n71 4.5005
R5098 VOUT.n94 VOUT.n66 4.5005
R5099 VOUT.n94 VOUT.t94 4.5005
R5100 VOUT.n94 VOUT.n65 4.5005
R5101 VOUT.n94 VOUT.n72 4.5005
R5102 VOUT.n94 VOUT.n73 4.5005
R5103 VOUT.n77 VOUT.n68 4.5005
R5104 VOUT.n77 VOUT.n70 4.5005
R5105 VOUT.n77 VOUT.n67 4.5005
R5106 VOUT.n77 VOUT.n71 4.5005
R5107 VOUT.n77 VOUT.n66 4.5005
R5108 VOUT.n77 VOUT.t94 4.5005
R5109 VOUT.n77 VOUT.n65 4.5005
R5110 VOUT.n77 VOUT.n72 4.5005
R5111 VOUT.n77 VOUT.n73 4.5005
R5112 VOUT.n169 VOUT.n68 4.5005
R5113 VOUT.n169 VOUT.n70 4.5005
R5114 VOUT.n169 VOUT.n67 4.5005
R5115 VOUT.n169 VOUT.n71 4.5005
R5116 VOUT.n169 VOUT.n66 4.5005
R5117 VOUT.n169 VOUT.t94 4.5005
R5118 VOUT.n169 VOUT.n65 4.5005
R5119 VOUT.n169 VOUT.n72 4.5005
R5120 VOUT.n169 VOUT.n73 4.5005
R5121 VOUT.n156 VOUT.n127 4.5005
R5122 VOUT.n156 VOUT.n133 4.5005
R5123 VOUT.n114 VOUT.n103 4.5005
R5124 VOUT.n114 VOUT.n105 4.5005
R5125 VOUT.n114 VOUT.n102 4.5005
R5126 VOUT.n114 VOUT.n106 4.5005
R5127 VOUT.n114 VOUT.n101 4.5005
R5128 VOUT.n114 VOUT.t92 4.5005
R5129 VOUT.n114 VOUT.n100 4.5005
R5130 VOUT.n114 VOUT.n107 4.5005
R5131 VOUT.n156 VOUT.n114 4.5005
R5132 VOUT.n135 VOUT.n103 4.5005
R5133 VOUT.n135 VOUT.n105 4.5005
R5134 VOUT.n135 VOUT.n102 4.5005
R5135 VOUT.n135 VOUT.n106 4.5005
R5136 VOUT.n135 VOUT.n101 4.5005
R5137 VOUT.n135 VOUT.t92 4.5005
R5138 VOUT.n135 VOUT.n100 4.5005
R5139 VOUT.n135 VOUT.n107 4.5005
R5140 VOUT.n156 VOUT.n135 4.5005
R5141 VOUT.n113 VOUT.n103 4.5005
R5142 VOUT.n113 VOUT.n105 4.5005
R5143 VOUT.n113 VOUT.n102 4.5005
R5144 VOUT.n113 VOUT.n106 4.5005
R5145 VOUT.n113 VOUT.n101 4.5005
R5146 VOUT.n113 VOUT.t92 4.5005
R5147 VOUT.n113 VOUT.n100 4.5005
R5148 VOUT.n113 VOUT.n107 4.5005
R5149 VOUT.n156 VOUT.n113 4.5005
R5150 VOUT.n137 VOUT.n103 4.5005
R5151 VOUT.n137 VOUT.n105 4.5005
R5152 VOUT.n137 VOUT.n102 4.5005
R5153 VOUT.n137 VOUT.n106 4.5005
R5154 VOUT.n137 VOUT.n101 4.5005
R5155 VOUT.n137 VOUT.t92 4.5005
R5156 VOUT.n137 VOUT.n100 4.5005
R5157 VOUT.n137 VOUT.n107 4.5005
R5158 VOUT.n156 VOUT.n137 4.5005
R5159 VOUT.n103 VOUT.n98 4.5005
R5160 VOUT.n105 VOUT.n98 4.5005
R5161 VOUT.n102 VOUT.n98 4.5005
R5162 VOUT.n106 VOUT.n98 4.5005
R5163 VOUT.n101 VOUT.n98 4.5005
R5164 VOUT.t92 VOUT.n98 4.5005
R5165 VOUT.n100 VOUT.n98 4.5005
R5166 VOUT.n107 VOUT.n98 4.5005
R5167 VOUT.n159 VOUT.n103 4.5005
R5168 VOUT.n159 VOUT.n105 4.5005
R5169 VOUT.n159 VOUT.n102 4.5005
R5170 VOUT.n159 VOUT.n106 4.5005
R5171 VOUT.n159 VOUT.n101 4.5005
R5172 VOUT.n159 VOUT.t92 4.5005
R5173 VOUT.n159 VOUT.n100 4.5005
R5174 VOUT.n159 VOUT.n107 4.5005
R5175 VOUT.n157 VOUT.n103 4.5005
R5176 VOUT.n157 VOUT.n105 4.5005
R5177 VOUT.n157 VOUT.n102 4.5005
R5178 VOUT.n157 VOUT.n106 4.5005
R5179 VOUT.n157 VOUT.n101 4.5005
R5180 VOUT.n157 VOUT.t92 4.5005
R5181 VOUT.n157 VOUT.n100 4.5005
R5182 VOUT.n157 VOUT.n107 4.5005
R5183 VOUT.n157 VOUT.n156 4.5005
R5184 VOUT.n139 VOUT.n103 4.5005
R5185 VOUT.n139 VOUT.n105 4.5005
R5186 VOUT.n139 VOUT.n102 4.5005
R5187 VOUT.n139 VOUT.n106 4.5005
R5188 VOUT.n139 VOUT.n101 4.5005
R5189 VOUT.n139 VOUT.t92 4.5005
R5190 VOUT.n139 VOUT.n100 4.5005
R5191 VOUT.n139 VOUT.n107 4.5005
R5192 VOUT.n156 VOUT.n139 4.5005
R5193 VOUT.n111 VOUT.n103 4.5005
R5194 VOUT.n111 VOUT.n105 4.5005
R5195 VOUT.n111 VOUT.n102 4.5005
R5196 VOUT.n111 VOUT.n106 4.5005
R5197 VOUT.n111 VOUT.n101 4.5005
R5198 VOUT.n111 VOUT.t92 4.5005
R5199 VOUT.n111 VOUT.n100 4.5005
R5200 VOUT.n111 VOUT.n107 4.5005
R5201 VOUT.n156 VOUT.n111 4.5005
R5202 VOUT.n141 VOUT.n103 4.5005
R5203 VOUT.n141 VOUT.n105 4.5005
R5204 VOUT.n141 VOUT.n102 4.5005
R5205 VOUT.n141 VOUT.n106 4.5005
R5206 VOUT.n141 VOUT.n101 4.5005
R5207 VOUT.n141 VOUT.t92 4.5005
R5208 VOUT.n141 VOUT.n100 4.5005
R5209 VOUT.n141 VOUT.n107 4.5005
R5210 VOUT.n156 VOUT.n141 4.5005
R5211 VOUT.n110 VOUT.n103 4.5005
R5212 VOUT.n110 VOUT.n105 4.5005
R5213 VOUT.n110 VOUT.n102 4.5005
R5214 VOUT.n110 VOUT.n106 4.5005
R5215 VOUT.n110 VOUT.n101 4.5005
R5216 VOUT.n110 VOUT.t92 4.5005
R5217 VOUT.n110 VOUT.n100 4.5005
R5218 VOUT.n110 VOUT.n107 4.5005
R5219 VOUT.n156 VOUT.n110 4.5005
R5220 VOUT.n155 VOUT.n103 4.5005
R5221 VOUT.n155 VOUT.n105 4.5005
R5222 VOUT.n155 VOUT.n102 4.5005
R5223 VOUT.n155 VOUT.n106 4.5005
R5224 VOUT.n155 VOUT.n101 4.5005
R5225 VOUT.n155 VOUT.t92 4.5005
R5226 VOUT.n155 VOUT.n100 4.5005
R5227 VOUT.n155 VOUT.n107 4.5005
R5228 VOUT.n156 VOUT.n155 4.5005
R5229 VOUT.n154 VOUT.n39 4.5005
R5230 VOUT.n55 VOUT.n39 4.5005
R5231 VOUT.n50 VOUT.n34 4.5005
R5232 VOUT.n50 VOUT.n36 4.5005
R5233 VOUT.n50 VOUT.n33 4.5005
R5234 VOUT.n50 VOUT.n37 4.5005
R5235 VOUT.n50 VOUT.n32 4.5005
R5236 VOUT.n50 VOUT.t93 4.5005
R5237 VOUT.n50 VOUT.n31 4.5005
R5238 VOUT.n50 VOUT.n38 4.5005
R5239 VOUT.n50 VOUT.n39 4.5005
R5240 VOUT.n48 VOUT.n34 4.5005
R5241 VOUT.n48 VOUT.n36 4.5005
R5242 VOUT.n48 VOUT.n33 4.5005
R5243 VOUT.n48 VOUT.n37 4.5005
R5244 VOUT.n48 VOUT.n32 4.5005
R5245 VOUT.n48 VOUT.t93 4.5005
R5246 VOUT.n48 VOUT.n31 4.5005
R5247 VOUT.n48 VOUT.n38 4.5005
R5248 VOUT.n48 VOUT.n39 4.5005
R5249 VOUT.n47 VOUT.n34 4.5005
R5250 VOUT.n47 VOUT.n36 4.5005
R5251 VOUT.n47 VOUT.n33 4.5005
R5252 VOUT.n47 VOUT.n37 4.5005
R5253 VOUT.n47 VOUT.n32 4.5005
R5254 VOUT.n47 VOUT.t93 4.5005
R5255 VOUT.n47 VOUT.n31 4.5005
R5256 VOUT.n47 VOUT.n38 4.5005
R5257 VOUT.n47 VOUT.n39 4.5005
R5258 VOUT.n176 VOUT.n34 4.5005
R5259 VOUT.n176 VOUT.n36 4.5005
R5260 VOUT.n176 VOUT.n33 4.5005
R5261 VOUT.n176 VOUT.n37 4.5005
R5262 VOUT.n176 VOUT.n32 4.5005
R5263 VOUT.n176 VOUT.t93 4.5005
R5264 VOUT.n176 VOUT.n31 4.5005
R5265 VOUT.n176 VOUT.n38 4.5005
R5266 VOUT.n176 VOUT.n39 4.5005
R5267 VOUT.n174 VOUT.n34 4.5005
R5268 VOUT.n174 VOUT.n36 4.5005
R5269 VOUT.n174 VOUT.n33 4.5005
R5270 VOUT.n174 VOUT.n37 4.5005
R5271 VOUT.n174 VOUT.n32 4.5005
R5272 VOUT.n174 VOUT.t93 4.5005
R5273 VOUT.n174 VOUT.n31 4.5005
R5274 VOUT.n174 VOUT.n38 4.5005
R5275 VOUT.n172 VOUT.n34 4.5005
R5276 VOUT.n172 VOUT.n36 4.5005
R5277 VOUT.n172 VOUT.n33 4.5005
R5278 VOUT.n172 VOUT.n37 4.5005
R5279 VOUT.n172 VOUT.n32 4.5005
R5280 VOUT.n172 VOUT.t93 4.5005
R5281 VOUT.n172 VOUT.n31 4.5005
R5282 VOUT.n172 VOUT.n38 4.5005
R5283 VOUT.n58 VOUT.n34 4.5005
R5284 VOUT.n58 VOUT.n36 4.5005
R5285 VOUT.n58 VOUT.n33 4.5005
R5286 VOUT.n58 VOUT.n37 4.5005
R5287 VOUT.n58 VOUT.n32 4.5005
R5288 VOUT.n58 VOUT.t93 4.5005
R5289 VOUT.n58 VOUT.n31 4.5005
R5290 VOUT.n58 VOUT.n38 4.5005
R5291 VOUT.n58 VOUT.n39 4.5005
R5292 VOUT.n57 VOUT.n34 4.5005
R5293 VOUT.n57 VOUT.n36 4.5005
R5294 VOUT.n57 VOUT.n33 4.5005
R5295 VOUT.n57 VOUT.n37 4.5005
R5296 VOUT.n57 VOUT.n32 4.5005
R5297 VOUT.n57 VOUT.t93 4.5005
R5298 VOUT.n57 VOUT.n31 4.5005
R5299 VOUT.n57 VOUT.n38 4.5005
R5300 VOUT.n57 VOUT.n39 4.5005
R5301 VOUT.n61 VOUT.n34 4.5005
R5302 VOUT.n61 VOUT.n36 4.5005
R5303 VOUT.n61 VOUT.n33 4.5005
R5304 VOUT.n61 VOUT.n37 4.5005
R5305 VOUT.n61 VOUT.n32 4.5005
R5306 VOUT.n61 VOUT.t93 4.5005
R5307 VOUT.n61 VOUT.n31 4.5005
R5308 VOUT.n61 VOUT.n38 4.5005
R5309 VOUT.n61 VOUT.n39 4.5005
R5310 VOUT.n60 VOUT.n34 4.5005
R5311 VOUT.n60 VOUT.n36 4.5005
R5312 VOUT.n60 VOUT.n33 4.5005
R5313 VOUT.n60 VOUT.n37 4.5005
R5314 VOUT.n60 VOUT.n32 4.5005
R5315 VOUT.n60 VOUT.t93 4.5005
R5316 VOUT.n60 VOUT.n31 4.5005
R5317 VOUT.n60 VOUT.n38 4.5005
R5318 VOUT.n60 VOUT.n39 4.5005
R5319 VOUT.n43 VOUT.n34 4.5005
R5320 VOUT.n43 VOUT.n36 4.5005
R5321 VOUT.n43 VOUT.n33 4.5005
R5322 VOUT.n43 VOUT.n37 4.5005
R5323 VOUT.n43 VOUT.n32 4.5005
R5324 VOUT.n43 VOUT.t93 4.5005
R5325 VOUT.n43 VOUT.n31 4.5005
R5326 VOUT.n43 VOUT.n38 4.5005
R5327 VOUT.n43 VOUT.n39 4.5005
R5328 VOUT.n179 VOUT.n34 4.5005
R5329 VOUT.n179 VOUT.n36 4.5005
R5330 VOUT.n179 VOUT.n33 4.5005
R5331 VOUT.n179 VOUT.n37 4.5005
R5332 VOUT.n179 VOUT.n32 4.5005
R5333 VOUT.n179 VOUT.t93 4.5005
R5334 VOUT.n179 VOUT.n31 4.5005
R5335 VOUT.n179 VOUT.n38 4.5005
R5336 VOUT.n179 VOUT.n39 4.5005
R5337 VOUT.n180 VOUT 3.7135
R5338 VOUT.n243 VOUT.n242 3.60085
R5339 VOUT.n223 VOUT.t0 3.3005
R5340 VOUT.n223 VOUT.t8 3.3005
R5341 VOUT.n221 VOUT.t90 3.3005
R5342 VOUT.n221 VOUT.t9 3.3005
R5343 VOUT.n219 VOUT.t24 3.3005
R5344 VOUT.n219 VOUT.t16 3.3005
R5345 VOUT.n218 VOUT.t3 3.3005
R5346 VOUT.n218 VOUT.t86 3.3005
R5347 VOUT.n216 VOUT.t20 3.3005
R5348 VOUT.n216 VOUT.t5 3.3005
R5349 VOUT.n214 VOUT.t12 3.3005
R5350 VOUT.n214 VOUT.t87 3.3005
R5351 VOUT.n212 VOUT.t11 3.3005
R5352 VOUT.n212 VOUT.t19 3.3005
R5353 VOUT.n211 VOUT.t7 3.3005
R5354 VOUT.n211 VOUT.t2 3.3005
R5355 VOUT.n234 VOUT.t6 3.3005
R5356 VOUT.n234 VOUT.t15 3.3005
R5357 VOUT.n235 VOUT.t88 3.3005
R5358 VOUT.n235 VOUT.t18 3.3005
R5359 VOUT.n237 VOUT.t17 3.3005
R5360 VOUT.n237 VOUT.t1 3.3005
R5361 VOUT.n239 VOUT.t10 3.3005
R5362 VOUT.n239 VOUT.t13 3.3005
R5363 VOUT.n227 VOUT.t4 3.3005
R5364 VOUT.n227 VOUT.t85 3.3005
R5365 VOUT.n228 VOUT.t22 3.3005
R5366 VOUT.n228 VOUT.t89 3.3005
R5367 VOUT.n230 VOUT.t91 3.3005
R5368 VOUT.n230 VOUT.t21 3.3005
R5369 VOUT.n232 VOUT.t23 3.3005
R5370 VOUT.n232 VOUT.t14 3.3005
R5371 VOUT.n242 VOUT.n226 2.72901
R5372 VOUT.n210 VOUT.n29 2.39875
R5373 VOUT.n120 VOUT.n118 2.251
R5374 VOUT.n120 VOUT.n117 2.251
R5375 VOUT.n120 VOUT.n116 2.251
R5376 VOUT.n120 VOUT.n115 2.251
R5377 VOUT.n89 VOUT.n88 2.251
R5378 VOUT.n89 VOUT.n87 2.251
R5379 VOUT.n89 VOUT.n86 2.251
R5380 VOUT.n89 VOUT.n85 2.251
R5381 VOUT.n162 VOUT.n161 2.251
R5382 VOUT.n127 VOUT.n125 2.251
R5383 VOUT.n127 VOUT.n124 2.251
R5384 VOUT.n127 VOUT.n123 2.251
R5385 VOUT.n145 VOUT.n127 2.251
R5386 VOUT.n133 VOUT.n132 2.251
R5387 VOUT.n133 VOUT.n131 2.251
R5388 VOUT.n133 VOUT.n130 2.251
R5389 VOUT.n133 VOUT.n129 2.251
R5390 VOUT.n159 VOUT.n99 2.251
R5391 VOUT.n154 VOUT.n152 2.251
R5392 VOUT.n154 VOUT.n151 2.251
R5393 VOUT.n154 VOUT.n150 2.251
R5394 VOUT.n154 VOUT.n149 2.251
R5395 VOUT.n55 VOUT.n54 2.251
R5396 VOUT.n55 VOUT.n53 2.251
R5397 VOUT.n55 VOUT.n52 2.251
R5398 VOUT.n55 VOUT.n51 2.251
R5399 VOUT.n172 VOUT.n171 2.251
R5400 VOUT.n89 VOUT.n69 2.2505
R5401 VOUT.n84 VOUT.n69 2.2505
R5402 VOUT.n82 VOUT.n69 2.2505
R5403 VOUT.n81 VOUT.n69 2.2505
R5404 VOUT.n166 VOUT.n69 2.2505
R5405 VOUT.n164 VOUT.n69 2.2505
R5406 VOUT.n162 VOUT.n69 2.2505
R5407 VOUT.n92 VOUT.n69 2.2505
R5408 VOUT.n91 VOUT.n69 2.2505
R5409 VOUT.n95 VOUT.n69 2.2505
R5410 VOUT.n94 VOUT.n69 2.2505
R5411 VOUT.n77 VOUT.n69 2.2505
R5412 VOUT.n169 VOUT.n69 2.2505
R5413 VOUT.n169 VOUT.n168 2.2505
R5414 VOUT.n133 VOUT.n104 2.2505
R5415 VOUT.n114 VOUT.n104 2.2505
R5416 VOUT.n135 VOUT.n104 2.2505
R5417 VOUT.n113 VOUT.n104 2.2505
R5418 VOUT.n137 VOUT.n104 2.2505
R5419 VOUT.n104 VOUT.n98 2.2505
R5420 VOUT.n159 VOUT.n104 2.2505
R5421 VOUT.n157 VOUT.n104 2.2505
R5422 VOUT.n139 VOUT.n104 2.2505
R5423 VOUT.n111 VOUT.n104 2.2505
R5424 VOUT.n141 VOUT.n104 2.2505
R5425 VOUT.n110 VOUT.n104 2.2505
R5426 VOUT.n155 VOUT.n104 2.2505
R5427 VOUT.n155 VOUT.n108 2.2505
R5428 VOUT.n55 VOUT.n35 2.2505
R5429 VOUT.n50 VOUT.n35 2.2505
R5430 VOUT.n48 VOUT.n35 2.2505
R5431 VOUT.n47 VOUT.n35 2.2505
R5432 VOUT.n176 VOUT.n35 2.2505
R5433 VOUT.n174 VOUT.n35 2.2505
R5434 VOUT.n172 VOUT.n35 2.2505
R5435 VOUT.n58 VOUT.n35 2.2505
R5436 VOUT.n57 VOUT.n35 2.2505
R5437 VOUT.n61 VOUT.n35 2.2505
R5438 VOUT.n60 VOUT.n35 2.2505
R5439 VOUT.n43 VOUT.n35 2.2505
R5440 VOUT.n179 VOUT.n35 2.2505
R5441 VOUT.n179 VOUT.n178 2.2505
R5442 VOUT.n97 VOUT.n90 2.25024
R5443 VOUT.n97 VOUT.n83 2.25024
R5444 VOUT.n165 VOUT.n97 2.25024
R5445 VOUT.n97 VOUT.n93 2.25024
R5446 VOUT.n97 VOUT.n96 2.25024
R5447 VOUT.n97 VOUT.n64 2.25024
R5448 VOUT.n147 VOUT.n144 2.25024
R5449 VOUT.n147 VOUT.n143 2.25024
R5450 VOUT.n147 VOUT.n142 2.25024
R5451 VOUT.n147 VOUT.n109 2.25024
R5452 VOUT.n147 VOUT.n146 2.25024
R5453 VOUT.n148 VOUT.n147 2.25024
R5454 VOUT.n63 VOUT.n56 2.25024
R5455 VOUT.n63 VOUT.n49 2.25024
R5456 VOUT.n175 VOUT.n63 2.25024
R5457 VOUT.n63 VOUT.n59 2.25024
R5458 VOUT.n63 VOUT.n62 2.25024
R5459 VOUT.n63 VOUT.n30 2.25024
R5460 VOUT.n209 VOUT.n199 2.12227
R5461 VOUT.n28 VOUT.n18 2.12227
R5462 VOUT.n164 VOUT.n74 1.50111
R5463 VOUT.n112 VOUT.n98 1.50111
R5464 VOUT.n174 VOUT.n40 1.50111
R5465 VOUT.n120 VOUT.n119 1.501
R5466 VOUT.n127 VOUT.n126 1.501
R5467 VOUT.n154 VOUT.n153 1.501
R5468 VOUT.n168 VOUT.n79 1.12536
R5469 VOUT.n168 VOUT.n80 1.12536
R5470 VOUT.n168 VOUT.n167 1.12536
R5471 VOUT.n128 VOUT.n108 1.12536
R5472 VOUT.n134 VOUT.n108 1.12536
R5473 VOUT.n136 VOUT.n108 1.12536
R5474 VOUT.n178 VOUT.n45 1.12536
R5475 VOUT.n178 VOUT.n46 1.12536
R5476 VOUT.n178 VOUT.n177 1.12536
R5477 VOUT.n168 VOUT.n75 1.12536
R5478 VOUT.n168 VOUT.n76 1.12536
R5479 VOUT.n168 VOUT.n78 1.12536
R5480 VOUT.n158 VOUT.n108 1.12536
R5481 VOUT.n138 VOUT.n108 1.12536
R5482 VOUT.n140 VOUT.n108 1.12536
R5483 VOUT.n178 VOUT.n41 1.12536
R5484 VOUT.n178 VOUT.n42 1.12536
R5485 VOUT.n178 VOUT.n44 1.12536
R5486 VOUT.n222 VOUT.n220 1.00481
R5487 VOUT.n224 VOUT.n222 1.00481
R5488 VOUT.n215 VOUT.n213 1.00481
R5489 VOUT.n217 VOUT.n215 1.00481
R5490 VOUT.n240 VOUT.n238 1.00481
R5491 VOUT.n238 VOUT.n236 1.00481
R5492 VOUT.n233 VOUT.n231 1.00481
R5493 VOUT.n231 VOUT.n229 1.00481
R5494 VOUT.n204 VOUT.n202 0.573776
R5495 VOUT.n206 VOUT.n204 0.573776
R5496 VOUT.n208 VOUT.n206 0.573776
R5497 VOUT.n194 VOUT.n192 0.573776
R5498 VOUT.n196 VOUT.n194 0.573776
R5499 VOUT.n198 VOUT.n196 0.573776
R5500 VOUT.n185 VOUT.n183 0.573776
R5501 VOUT.n187 VOUT.n185 0.573776
R5502 VOUT.n189 VOUT.n187 0.573776
R5503 VOUT.n27 VOUT.n25 0.573776
R5504 VOUT.n25 VOUT.n23 0.573776
R5505 VOUT.n23 VOUT.n21 0.573776
R5506 VOUT.n17 VOUT.n15 0.573776
R5507 VOUT.n15 VOUT.n13 0.573776
R5508 VOUT.n13 VOUT.n11 0.573776
R5509 VOUT.n8 VOUT.n6 0.573776
R5510 VOUT.n6 VOUT.n4 0.573776
R5511 VOUT.n4 VOUT.n2 0.573776
R5512 VOUT.n180 VOUT.n179 0.373399
R5513 VOUT.n243 VOUT.n180 0.3624
R5514 VOUT.n122 VOUT.n121 0.0910737
R5515 VOUT.n173 VOUT.n170 0.0723685
R5516 VOUT.n127 VOUT.n122 0.0522944
R5517 VOUT.n170 VOUT.n169 0.0499135
R5518 VOUT.n121 VOUT.n120 0.0499135
R5519 VOUT.n155 VOUT.n154 0.0464294
R5520 VOUT.n163 VOUT.n160 0.0391444
R5521 VOUT.n122 VOUT.t95 0.023435
R5522 VOUT.n170 VOUT.t96 0.02262
R5523 VOUT.n121 VOUT.t97 0.02262
R5524 VOUT VOUT.n243 0.0099
R5525 VOUT.n92 VOUT.n75 0.00365111
R5526 VOUT.n95 VOUT.n76 0.00365111
R5527 VOUT.n78 VOUT.n77 0.00365111
R5528 VOUT.n120 VOUT.n79 0.00365111
R5529 VOUT.n84 VOUT.n80 0.00365111
R5530 VOUT.n167 VOUT.n81 0.00365111
R5531 VOUT.n158 VOUT.n157 0.00365111
R5532 VOUT.n138 VOUT.n111 0.00365111
R5533 VOUT.n140 VOUT.n110 0.00365111
R5534 VOUT.n128 VOUT.n127 0.00365111
R5535 VOUT.n134 VOUT.n114 0.00365111
R5536 VOUT.n136 VOUT.n113 0.00365111
R5537 VOUT.n58 VOUT.n41 0.00365111
R5538 VOUT.n61 VOUT.n42 0.00365111
R5539 VOUT.n44 VOUT.n43 0.00365111
R5540 VOUT.n154 VOUT.n45 0.00365111
R5541 VOUT.n50 VOUT.n46 0.00365111
R5542 VOUT.n177 VOUT.n47 0.00365111
R5543 VOUT.n89 VOUT.n79 0.00340054
R5544 VOUT.n82 VOUT.n80 0.00340054
R5545 VOUT.n167 VOUT.n166 0.00340054
R5546 VOUT.n162 VOUT.n75 0.00340054
R5547 VOUT.n91 VOUT.n76 0.00340054
R5548 VOUT.n94 VOUT.n78 0.00340054
R5549 VOUT.n133 VOUT.n128 0.00340054
R5550 VOUT.n135 VOUT.n134 0.00340054
R5551 VOUT.n137 VOUT.n136 0.00340054
R5552 VOUT.n159 VOUT.n158 0.00340054
R5553 VOUT.n139 VOUT.n138 0.00340054
R5554 VOUT.n141 VOUT.n140 0.00340054
R5555 VOUT.n55 VOUT.n45 0.00340054
R5556 VOUT.n48 VOUT.n46 0.00340054
R5557 VOUT.n177 VOUT.n176 0.00340054
R5558 VOUT.n172 VOUT.n41 0.00340054
R5559 VOUT.n57 VOUT.n42 0.00340054
R5560 VOUT.n60 VOUT.n44 0.00340054
R5561 VOUT.n90 VOUT.n84 0.00252698
R5562 VOUT.n83 VOUT.n81 0.00252698
R5563 VOUT.n165 VOUT.n164 0.00252698
R5564 VOUT.n93 VOUT.n91 0.00252698
R5565 VOUT.n96 VOUT.n94 0.00252698
R5566 VOUT.n169 VOUT.n64 0.00252698
R5567 VOUT.n90 VOUT.n89 0.00252698
R5568 VOUT.n83 VOUT.n82 0.00252698
R5569 VOUT.n166 VOUT.n165 0.00252698
R5570 VOUT.n93 VOUT.n92 0.00252698
R5571 VOUT.n96 VOUT.n95 0.00252698
R5572 VOUT.n77 VOUT.n64 0.00252698
R5573 VOUT.n144 VOUT.n114 0.00252698
R5574 VOUT.n143 VOUT.n113 0.00252698
R5575 VOUT.n142 VOUT.n98 0.00252698
R5576 VOUT.n139 VOUT.n109 0.00252698
R5577 VOUT.n146 VOUT.n141 0.00252698
R5578 VOUT.n155 VOUT.n148 0.00252698
R5579 VOUT.n144 VOUT.n133 0.00252698
R5580 VOUT.n143 VOUT.n135 0.00252698
R5581 VOUT.n142 VOUT.n137 0.00252698
R5582 VOUT.n157 VOUT.n109 0.00252698
R5583 VOUT.n146 VOUT.n111 0.00252698
R5584 VOUT.n148 VOUT.n110 0.00252698
R5585 VOUT.n56 VOUT.n50 0.00252698
R5586 VOUT.n49 VOUT.n47 0.00252698
R5587 VOUT.n175 VOUT.n174 0.00252698
R5588 VOUT.n59 VOUT.n57 0.00252698
R5589 VOUT.n62 VOUT.n60 0.00252698
R5590 VOUT.n179 VOUT.n30 0.00252698
R5591 VOUT.n56 VOUT.n55 0.00252698
R5592 VOUT.n49 VOUT.n48 0.00252698
R5593 VOUT.n176 VOUT.n175 0.00252698
R5594 VOUT.n59 VOUT.n58 0.00252698
R5595 VOUT.n62 VOUT.n61 0.00252698
R5596 VOUT.n43 VOUT.n30 0.00252698
R5597 VOUT.n164 VOUT.n163 0.0020275
R5598 VOUT.n163 VOUT.n162 0.0020275
R5599 VOUT.n160 VOUT.n98 0.0020275
R5600 VOUT.n160 VOUT.n159 0.0020275
R5601 VOUT.n174 VOUT.n173 0.0020275
R5602 VOUT.n173 VOUT.n172 0.0020275
R5603 VOUT.n74 VOUT.n73 0.00166668
R5604 VOUT.n156 VOUT.n112 0.00166668
R5605 VOUT.n40 VOUT.n39 0.00166668
R5606 VOUT.n178 VOUT.n40 0.00133328
R5607 VOUT.n112 VOUT.n108 0.00133328
R5608 VOUT.n168 VOUT.n74 0.00133328
R5609 VOUT.n171 VOUT.n63 0.001
R5610 VOUT.n149 VOUT.n63 0.001
R5611 VOUT.n51 VOUT.n31 0.001
R5612 VOUT.n150 VOUT.n31 0.001
R5613 VOUT.n52 VOUT.n32 0.001
R5614 VOUT.n151 VOUT.n32 0.001
R5615 VOUT.n53 VOUT.n33 0.001
R5616 VOUT.n152 VOUT.n33 0.001
R5617 VOUT.n54 VOUT.n34 0.001
R5618 VOUT.n153 VOUT.n34 0.001
R5619 VOUT.n147 VOUT.n99 0.001
R5620 VOUT.n147 VOUT.n145 0.001
R5621 VOUT.n129 VOUT.n100 0.001
R5622 VOUT.n123 VOUT.n100 0.001
R5623 VOUT.n130 VOUT.n101 0.001
R5624 VOUT.n124 VOUT.n101 0.001
R5625 VOUT.n131 VOUT.n102 0.001
R5626 VOUT.n125 VOUT.n102 0.001
R5627 VOUT.n132 VOUT.n103 0.001
R5628 VOUT.n126 VOUT.n103 0.001
R5629 VOUT.n161 VOUT.n97 0.001
R5630 VOUT.n115 VOUT.n97 0.001
R5631 VOUT.n85 VOUT.n65 0.001
R5632 VOUT.n116 VOUT.n65 0.001
R5633 VOUT.n86 VOUT.n66 0.001
R5634 VOUT.n117 VOUT.n66 0.001
R5635 VOUT.n87 VOUT.n67 0.001
R5636 VOUT.n118 VOUT.n67 0.001
R5637 VOUT.n88 VOUT.n68 0.001
R5638 VOUT.n119 VOUT.n68 0.001
R5639 VOUT.n119 VOUT.n69 0.001
R5640 VOUT.n118 VOUT.n70 0.001
R5641 VOUT.n117 VOUT.n71 0.001
R5642 VOUT.n116 VOUT.t94 0.001
R5643 VOUT.n115 VOUT.n72 0.001
R5644 VOUT.n88 VOUT.n70 0.001
R5645 VOUT.n87 VOUT.n71 0.001
R5646 VOUT.n86 VOUT.t94 0.001
R5647 VOUT.n85 VOUT.n72 0.001
R5648 VOUT.n161 VOUT.n73 0.001
R5649 VOUT.n126 VOUT.n104 0.001
R5650 VOUT.n125 VOUT.n105 0.001
R5651 VOUT.n124 VOUT.n106 0.001
R5652 VOUT.n123 VOUT.t92 0.001
R5653 VOUT.n145 VOUT.n107 0.001
R5654 VOUT.n132 VOUT.n105 0.001
R5655 VOUT.n131 VOUT.n106 0.001
R5656 VOUT.n130 VOUT.t92 0.001
R5657 VOUT.n129 VOUT.n107 0.001
R5658 VOUT.n156 VOUT.n99 0.001
R5659 VOUT.n153 VOUT.n35 0.001
R5660 VOUT.n152 VOUT.n36 0.001
R5661 VOUT.n151 VOUT.n37 0.001
R5662 VOUT.n150 VOUT.t93 0.001
R5663 VOUT.n149 VOUT.n38 0.001
R5664 VOUT.n54 VOUT.n36 0.001
R5665 VOUT.n53 VOUT.n37 0.001
R5666 VOUT.n52 VOUT.t93 0.001
R5667 VOUT.n51 VOUT.n38 0.001
R5668 VOUT.n171 VOUT.n39 0.001
R5669 CS_BIAS.n201 CS_BIAS.n139 161.3
R5670 CS_BIAS.n200 CS_BIAS.n199 161.3
R5671 CS_BIAS.n198 CS_BIAS.n140 161.3
R5672 CS_BIAS.n197 CS_BIAS.n196 161.3
R5673 CS_BIAS.n194 CS_BIAS.n141 161.3
R5674 CS_BIAS.n193 CS_BIAS.n192 161.3
R5675 CS_BIAS.n191 CS_BIAS.n142 161.3
R5676 CS_BIAS.n190 CS_BIAS.n189 161.3
R5677 CS_BIAS.n188 CS_BIAS.n143 161.3
R5678 CS_BIAS.n186 CS_BIAS.n185 161.3
R5679 CS_BIAS.n184 CS_BIAS.n144 161.3
R5680 CS_BIAS.n183 CS_BIAS.n182 161.3
R5681 CS_BIAS.n181 CS_BIAS.n145 161.3
R5682 CS_BIAS.n180 CS_BIAS.n179 161.3
R5683 CS_BIAS.n178 CS_BIAS.n177 161.3
R5684 CS_BIAS.n176 CS_BIAS.n147 161.3
R5685 CS_BIAS.n175 CS_BIAS.n174 161.3
R5686 CS_BIAS.n173 CS_BIAS.n148 161.3
R5687 CS_BIAS.n172 CS_BIAS.n171 161.3
R5688 CS_BIAS.n170 CS_BIAS.n149 161.3
R5689 CS_BIAS.n169 CS_BIAS.n168 161.3
R5690 CS_BIAS.n167 CS_BIAS.n151 161.3
R5691 CS_BIAS.n166 CS_BIAS.n165 161.3
R5692 CS_BIAS.n163 CS_BIAS.n152 161.3
R5693 CS_BIAS.n162 CS_BIAS.n161 161.3
R5694 CS_BIAS.n160 CS_BIAS.n153 161.3
R5695 CS_BIAS.n159 CS_BIAS.n158 161.3
R5696 CS_BIAS.n157 CS_BIAS.n154 161.3
R5697 CS_BIAS.n28 CS_BIAS.n25 161.3
R5698 CS_BIAS.n30 CS_BIAS.n29 161.3
R5699 CS_BIAS.n31 CS_BIAS.n24 161.3
R5700 CS_BIAS.n33 CS_BIAS.n32 161.3
R5701 CS_BIAS.n34 CS_BIAS.n23 161.3
R5702 CS_BIAS.n37 CS_BIAS.n36 161.3
R5703 CS_BIAS.n38 CS_BIAS.n22 161.3
R5704 CS_BIAS.n40 CS_BIAS.n39 161.3
R5705 CS_BIAS.n41 CS_BIAS.n20 161.3
R5706 CS_BIAS.n43 CS_BIAS.n42 161.3
R5707 CS_BIAS.n44 CS_BIAS.n19 161.3
R5708 CS_BIAS.n46 CS_BIAS.n45 161.3
R5709 CS_BIAS.n47 CS_BIAS.n18 161.3
R5710 CS_BIAS.n49 CS_BIAS.n48 161.3
R5711 CS_BIAS.n51 CS_BIAS.n50 161.3
R5712 CS_BIAS.n52 CS_BIAS.n16 161.3
R5713 CS_BIAS.n54 CS_BIAS.n53 161.3
R5714 CS_BIAS.n55 CS_BIAS.n15 161.3
R5715 CS_BIAS.n57 CS_BIAS.n56 161.3
R5716 CS_BIAS.n59 CS_BIAS.n14 161.3
R5717 CS_BIAS.n61 CS_BIAS.n60 161.3
R5718 CS_BIAS.n62 CS_BIAS.n13 161.3
R5719 CS_BIAS.n64 CS_BIAS.n63 161.3
R5720 CS_BIAS.n65 CS_BIAS.n12 161.3
R5721 CS_BIAS.n68 CS_BIAS.n67 161.3
R5722 CS_BIAS.n69 CS_BIAS.n11 161.3
R5723 CS_BIAS.n71 CS_BIAS.n70 161.3
R5724 CS_BIAS.n72 CS_BIAS.n10 161.3
R5725 CS_BIAS.n92 CS_BIAS.n89 161.3
R5726 CS_BIAS.n94 CS_BIAS.n93 161.3
R5727 CS_BIAS.n95 CS_BIAS.n88 161.3
R5728 CS_BIAS.n97 CS_BIAS.n96 161.3
R5729 CS_BIAS.n98 CS_BIAS.n87 161.3
R5730 CS_BIAS.n101 CS_BIAS.n100 161.3
R5731 CS_BIAS.n102 CS_BIAS.n86 161.3
R5732 CS_BIAS.n104 CS_BIAS.n103 161.3
R5733 CS_BIAS.n105 CS_BIAS.n84 161.3
R5734 CS_BIAS.n107 CS_BIAS.n106 161.3
R5735 CS_BIAS.n108 CS_BIAS.n9 161.3
R5736 CS_BIAS.n110 CS_BIAS.n109 161.3
R5737 CS_BIAS.n111 CS_BIAS.n8 161.3
R5738 CS_BIAS.n113 CS_BIAS.n112 161.3
R5739 CS_BIAS.n115 CS_BIAS.n114 161.3
R5740 CS_BIAS.n116 CS_BIAS.n6 161.3
R5741 CS_BIAS.n118 CS_BIAS.n117 161.3
R5742 CS_BIAS.n119 CS_BIAS.n5 161.3
R5743 CS_BIAS.n121 CS_BIAS.n120 161.3
R5744 CS_BIAS.n123 CS_BIAS.n4 161.3
R5745 CS_BIAS.n125 CS_BIAS.n124 161.3
R5746 CS_BIAS.n126 CS_BIAS.n3 161.3
R5747 CS_BIAS.n128 CS_BIAS.n127 161.3
R5748 CS_BIAS.n129 CS_BIAS.n2 161.3
R5749 CS_BIAS.n132 CS_BIAS.n131 161.3
R5750 CS_BIAS.n133 CS_BIAS.n1 161.3
R5751 CS_BIAS.n135 CS_BIAS.n134 161.3
R5752 CS_BIAS.n136 CS_BIAS.n0 161.3
R5753 CS_BIAS.n406 CS_BIAS.n344 161.3
R5754 CS_BIAS.n405 CS_BIAS.n404 161.3
R5755 CS_BIAS.n403 CS_BIAS.n345 161.3
R5756 CS_BIAS.n402 CS_BIAS.n401 161.3
R5757 CS_BIAS.n399 CS_BIAS.n346 161.3
R5758 CS_BIAS.n398 CS_BIAS.n397 161.3
R5759 CS_BIAS.n396 CS_BIAS.n347 161.3
R5760 CS_BIAS.n395 CS_BIAS.n394 161.3
R5761 CS_BIAS.n393 CS_BIAS.n348 161.3
R5762 CS_BIAS.n391 CS_BIAS.n390 161.3
R5763 CS_BIAS.n389 CS_BIAS.n349 161.3
R5764 CS_BIAS.n388 CS_BIAS.n387 161.3
R5765 CS_BIAS.n386 CS_BIAS.n350 161.3
R5766 CS_BIAS.n385 CS_BIAS.n384 161.3
R5767 CS_BIAS.n383 CS_BIAS.n382 161.3
R5768 CS_BIAS.n381 CS_BIAS.n352 161.3
R5769 CS_BIAS.n380 CS_BIAS.n379 161.3
R5770 CS_BIAS.n378 CS_BIAS.n353 161.3
R5771 CS_BIAS.n377 CS_BIAS.n376 161.3
R5772 CS_BIAS.n374 CS_BIAS.n354 161.3
R5773 CS_BIAS.n373 CS_BIAS.n372 161.3
R5774 CS_BIAS.n371 CS_BIAS.n355 161.3
R5775 CS_BIAS.n370 CS_BIAS.n369 161.3
R5776 CS_BIAS.n367 CS_BIAS.n356 161.3
R5777 CS_BIAS.n366 CS_BIAS.n365 161.3
R5778 CS_BIAS.n364 CS_BIAS.n357 161.3
R5779 CS_BIAS.n363 CS_BIAS.n362 161.3
R5780 CS_BIAS.n361 CS_BIAS.n358 161.3
R5781 CS_BIAS.n305 CS_BIAS.n243 161.3
R5782 CS_BIAS.n304 CS_BIAS.n303 161.3
R5783 CS_BIAS.n302 CS_BIAS.n244 161.3
R5784 CS_BIAS.n301 CS_BIAS.n300 161.3
R5785 CS_BIAS.n298 CS_BIAS.n245 161.3
R5786 CS_BIAS.n297 CS_BIAS.n296 161.3
R5787 CS_BIAS.n295 CS_BIAS.n246 161.3
R5788 CS_BIAS.n294 CS_BIAS.n293 161.3
R5789 CS_BIAS.n292 CS_BIAS.n247 161.3
R5790 CS_BIAS.n290 CS_BIAS.n289 161.3
R5791 CS_BIAS.n288 CS_BIAS.n248 161.3
R5792 CS_BIAS.n287 CS_BIAS.n286 161.3
R5793 CS_BIAS.n285 CS_BIAS.n249 161.3
R5794 CS_BIAS.n284 CS_BIAS.n283 161.3
R5795 CS_BIAS.n282 CS_BIAS.n281 161.3
R5796 CS_BIAS.n280 CS_BIAS.n251 161.3
R5797 CS_BIAS.n279 CS_BIAS.n278 161.3
R5798 CS_BIAS.n277 CS_BIAS.n252 161.3
R5799 CS_BIAS.n276 CS_BIAS.n275 161.3
R5800 CS_BIAS.n273 CS_BIAS.n253 161.3
R5801 CS_BIAS.n272 CS_BIAS.n271 161.3
R5802 CS_BIAS.n270 CS_BIAS.n254 161.3
R5803 CS_BIAS.n269 CS_BIAS.n268 161.3
R5804 CS_BIAS.n266 CS_BIAS.n255 161.3
R5805 CS_BIAS.n265 CS_BIAS.n264 161.3
R5806 CS_BIAS.n263 CS_BIAS.n256 161.3
R5807 CS_BIAS.n262 CS_BIAS.n261 161.3
R5808 CS_BIAS.n260 CS_BIAS.n257 161.3
R5809 CS_BIAS.n315 CS_BIAS.n314 161.3
R5810 CS_BIAS.n239 CS_BIAS.n214 161.3
R5811 CS_BIAS.n238 CS_BIAS.n237 161.3
R5812 CS_BIAS.n235 CS_BIAS.n215 161.3
R5813 CS_BIAS.n234 CS_BIAS.n233 161.3
R5814 CS_BIAS.n232 CS_BIAS.n216 161.3
R5815 CS_BIAS.n231 CS_BIAS.n230 161.3
R5816 CS_BIAS.n228 CS_BIAS.n217 161.3
R5817 CS_BIAS.n227 CS_BIAS.n226 161.3
R5818 CS_BIAS.n225 CS_BIAS.n218 161.3
R5819 CS_BIAS.n224 CS_BIAS.n223 161.3
R5820 CS_BIAS.n222 CS_BIAS.n219 161.3
R5821 CS_BIAS.n341 CS_BIAS.n205 161.3
R5822 CS_BIAS.n340 CS_BIAS.n339 161.3
R5823 CS_BIAS.n338 CS_BIAS.n206 161.3
R5824 CS_BIAS.n337 CS_BIAS.n336 161.3
R5825 CS_BIAS.n334 CS_BIAS.n207 161.3
R5826 CS_BIAS.n333 CS_BIAS.n332 161.3
R5827 CS_BIAS.n331 CS_BIAS.n208 161.3
R5828 CS_BIAS.n330 CS_BIAS.n329 161.3
R5829 CS_BIAS.n328 CS_BIAS.n209 161.3
R5830 CS_BIAS.n326 CS_BIAS.n325 161.3
R5831 CS_BIAS.n324 CS_BIAS.n210 161.3
R5832 CS_BIAS.n323 CS_BIAS.n322 161.3
R5833 CS_BIAS.n321 CS_BIAS.n211 161.3
R5834 CS_BIAS.n320 CS_BIAS.n319 161.3
R5835 CS_BIAS.n318 CS_BIAS.n317 161.3
R5836 CS_BIAS.n316 CS_BIAS.n213 161.3
R5837 CS_BIAS.n155 CS_BIAS.t40 102.697
R5838 CS_BIAS.n359 CS_BIAS.t50 102.697
R5839 CS_BIAS.n258 CS_BIAS.t24 102.697
R5840 CS_BIAS.n220 CS_BIAS.t56 102.697
R5841 CS_BIAS.n26 CS_BIAS.t26 102.697
R5842 CS_BIAS.n90 CS_BIAS.t44 102.697
R5843 CS_BIAS.n203 CS_BIAS.n202 90.9889
R5844 CS_BIAS.n74 CS_BIAS.n73 90.9889
R5845 CS_BIAS.n138 CS_BIAS.n137 90.9889
R5846 CS_BIAS.n408 CS_BIAS.n407 90.9889
R5847 CS_BIAS.n307 CS_BIAS.n306 90.9889
R5848 CS_BIAS.n343 CS_BIAS.n342 90.9889
R5849 CS_BIAS.n81 CS_BIAS.n79 85.0679
R5850 CS_BIAS.n242 CS_BIAS.n240 85.0679
R5851 CS_BIAS.n81 CS_BIAS.n80 84.0635
R5852 CS_BIAS.n78 CS_BIAS.n77 84.0635
R5853 CS_BIAS.n76 CS_BIAS.n75 84.0635
R5854 CS_BIAS.n309 CS_BIAS.n308 84.0635
R5855 CS_BIAS.n311 CS_BIAS.n310 84.0635
R5856 CS_BIAS.n242 CS_BIAS.n241 84.0635
R5857 CS_BIAS.n156 CS_BIAS.t37 72.3005
R5858 CS_BIAS.n164 CS_BIAS.t47 72.3005
R5859 CS_BIAS.n150 CS_BIAS.t46 72.3005
R5860 CS_BIAS.n146 CS_BIAS.t62 72.3005
R5861 CS_BIAS.n187 CS_BIAS.t63 72.3005
R5862 CS_BIAS.n195 CS_BIAS.t61 72.3005
R5863 CS_BIAS.n202 CS_BIAS.t48 72.3005
R5864 CS_BIAS.n73 CS_BIAS.t6 72.3005
R5865 CS_BIAS.n66 CS_BIAS.t30 72.3005
R5866 CS_BIAS.n58 CS_BIAS.t22 72.3005
R5867 CS_BIAS.n17 CS_BIAS.t18 72.3005
R5868 CS_BIAS.n21 CS_BIAS.t0 72.3005
R5869 CS_BIAS.n35 CS_BIAS.t16 72.3005
R5870 CS_BIAS.n27 CS_BIAS.t2 72.3005
R5871 CS_BIAS.n137 CS_BIAS.t55 72.3005
R5872 CS_BIAS.n130 CS_BIAS.t35 72.3005
R5873 CS_BIAS.n122 CS_BIAS.t39 72.3005
R5874 CS_BIAS.n7 CS_BIAS.t36 72.3005
R5875 CS_BIAS.n85 CS_BIAS.t51 72.3005
R5876 CS_BIAS.n99 CS_BIAS.t52 72.3005
R5877 CS_BIAS.n91 CS_BIAS.t42 72.3005
R5878 CS_BIAS.n360 CS_BIAS.t59 72.3005
R5879 CS_BIAS.n368 CS_BIAS.t38 72.3005
R5880 CS_BIAS.n375 CS_BIAS.t34 72.3005
R5881 CS_BIAS.n351 CS_BIAS.t53 72.3005
R5882 CS_BIAS.n392 CS_BIAS.t45 72.3005
R5883 CS_BIAS.n400 CS_BIAS.t54 72.3005
R5884 CS_BIAS.n407 CS_BIAS.t60 72.3005
R5885 CS_BIAS.n259 CS_BIAS.t14 72.3005
R5886 CS_BIAS.n267 CS_BIAS.t20 72.3005
R5887 CS_BIAS.n274 CS_BIAS.t12 72.3005
R5888 CS_BIAS.n250 CS_BIAS.t8 72.3005
R5889 CS_BIAS.n291 CS_BIAS.t10 72.3005
R5890 CS_BIAS.n299 CS_BIAS.t4 72.3005
R5891 CS_BIAS.n306 CS_BIAS.t28 72.3005
R5892 CS_BIAS.n342 CS_BIAS.t33 72.3005
R5893 CS_BIAS.n335 CS_BIAS.t58 72.3005
R5894 CS_BIAS.n327 CS_BIAS.t49 72.3005
R5895 CS_BIAS.n212 CS_BIAS.t57 72.3005
R5896 CS_BIAS.n221 CS_BIAS.t32 72.3005
R5897 CS_BIAS.n229 CS_BIAS.t43 72.3005
R5898 CS_BIAS.n236 CS_BIAS.t41 72.3005
R5899 CS_BIAS.n27 CS_BIAS.n26 66.3065
R5900 CS_BIAS.n91 CS_BIAS.n90 66.3065
R5901 CS_BIAS.n156 CS_BIAS.n155 66.3065
R5902 CS_BIAS.n360 CS_BIAS.n359 66.3065
R5903 CS_BIAS.n259 CS_BIAS.n258 66.3065
R5904 CS_BIAS.n221 CS_BIAS.n220 66.3065
R5905 CS_BIAS.n176 CS_BIAS.n175 56.5617
R5906 CS_BIAS.n200 CS_BIAS.n140 56.5617
R5907 CS_BIAS.n47 CS_BIAS.n46 56.5617
R5908 CS_BIAS.n111 CS_BIAS.n110 56.5617
R5909 CS_BIAS.n381 CS_BIAS.n380 56.5617
R5910 CS_BIAS.n405 CS_BIAS.n345 56.5617
R5911 CS_BIAS.n280 CS_BIAS.n279 56.5617
R5912 CS_BIAS.n304 CS_BIAS.n244 56.5617
R5913 CS_BIAS.n316 CS_BIAS.n315 56.5617
R5914 CS_BIAS.n71 CS_BIAS.n11 56.5617
R5915 CS_BIAS.n135 CS_BIAS.n1 56.5617
R5916 CS_BIAS.n340 CS_BIAS.n206 56.5617
R5917 CS_BIAS.n162 CS_BIAS.n153 49.296
R5918 CS_BIAS.n189 CS_BIAS.n142 49.296
R5919 CS_BIAS.n60 CS_BIAS.n13 49.296
R5920 CS_BIAS.n33 CS_BIAS.n24 49.296
R5921 CS_BIAS.n124 CS_BIAS.n3 49.296
R5922 CS_BIAS.n97 CS_BIAS.n88 49.296
R5923 CS_BIAS.n366 CS_BIAS.n357 49.296
R5924 CS_BIAS.n394 CS_BIAS.n347 49.296
R5925 CS_BIAS.n265 CS_BIAS.n256 49.296
R5926 CS_BIAS.n293 CS_BIAS.n246 49.296
R5927 CS_BIAS.n329 CS_BIAS.n208 49.296
R5928 CS_BIAS.n227 CS_BIAS.n218 49.296
R5929 CS_BIAS.n169 CS_BIAS.n151 48.3272
R5930 CS_BIAS.n182 CS_BIAS.n144 48.3272
R5931 CS_BIAS.n53 CS_BIAS.n15 48.3272
R5932 CS_BIAS.n40 CS_BIAS.n22 48.3272
R5933 CS_BIAS.n117 CS_BIAS.n5 48.3272
R5934 CS_BIAS.n104 CS_BIAS.n86 48.3272
R5935 CS_BIAS.n373 CS_BIAS.n355 48.3272
R5936 CS_BIAS.n387 CS_BIAS.n349 48.3272
R5937 CS_BIAS.n272 CS_BIAS.n254 48.3272
R5938 CS_BIAS.n286 CS_BIAS.n248 48.3272
R5939 CS_BIAS.n322 CS_BIAS.n210 48.3272
R5940 CS_BIAS.n234 CS_BIAS.n216 48.3272
R5941 CS_BIAS.n170 CS_BIAS.n169 32.8269
R5942 CS_BIAS.n182 CS_BIAS.n181 32.8269
R5943 CS_BIAS.n53 CS_BIAS.n52 32.8269
R5944 CS_BIAS.n41 CS_BIAS.n40 32.8269
R5945 CS_BIAS.n117 CS_BIAS.n116 32.8269
R5946 CS_BIAS.n105 CS_BIAS.n104 32.8269
R5947 CS_BIAS.n374 CS_BIAS.n373 32.8269
R5948 CS_BIAS.n387 CS_BIAS.n386 32.8269
R5949 CS_BIAS.n273 CS_BIAS.n272 32.8269
R5950 CS_BIAS.n286 CS_BIAS.n285 32.8269
R5951 CS_BIAS.n322 CS_BIAS.n321 32.8269
R5952 CS_BIAS.n235 CS_BIAS.n234 32.8269
R5953 CS_BIAS.n158 CS_BIAS.n153 31.8581
R5954 CS_BIAS.n193 CS_BIAS.n142 31.8581
R5955 CS_BIAS.n64 CS_BIAS.n13 31.8581
R5956 CS_BIAS.n29 CS_BIAS.n24 31.8581
R5957 CS_BIAS.n128 CS_BIAS.n3 31.8581
R5958 CS_BIAS.n93 CS_BIAS.n88 31.8581
R5959 CS_BIAS.n362 CS_BIAS.n357 31.8581
R5960 CS_BIAS.n398 CS_BIAS.n347 31.8581
R5961 CS_BIAS.n261 CS_BIAS.n256 31.8581
R5962 CS_BIAS.n297 CS_BIAS.n246 31.8581
R5963 CS_BIAS.n333 CS_BIAS.n208 31.8581
R5964 CS_BIAS.n223 CS_BIAS.n218 31.8581
R5965 CS_BIAS.n158 CS_BIAS.n157 24.5923
R5966 CS_BIAS.n165 CS_BIAS.n151 24.5923
R5967 CS_BIAS.n163 CS_BIAS.n162 24.5923
R5968 CS_BIAS.n175 CS_BIAS.n148 24.5923
R5969 CS_BIAS.n171 CS_BIAS.n170 24.5923
R5970 CS_BIAS.n181 CS_BIAS.n180 24.5923
R5971 CS_BIAS.n177 CS_BIAS.n176 24.5923
R5972 CS_BIAS.n189 CS_BIAS.n188 24.5923
R5973 CS_BIAS.n186 CS_BIAS.n144 24.5923
R5974 CS_BIAS.n196 CS_BIAS.n140 24.5923
R5975 CS_BIAS.n194 CS_BIAS.n193 24.5923
R5976 CS_BIAS.n201 CS_BIAS.n200 24.5923
R5977 CS_BIAS.n72 CS_BIAS.n71 24.5923
R5978 CS_BIAS.n67 CS_BIAS.n11 24.5923
R5979 CS_BIAS.n65 CS_BIAS.n64 24.5923
R5980 CS_BIAS.n60 CS_BIAS.n59 24.5923
R5981 CS_BIAS.n57 CS_BIAS.n15 24.5923
R5982 CS_BIAS.n52 CS_BIAS.n51 24.5923
R5983 CS_BIAS.n48 CS_BIAS.n47 24.5923
R5984 CS_BIAS.n46 CS_BIAS.n19 24.5923
R5985 CS_BIAS.n42 CS_BIAS.n41 24.5923
R5986 CS_BIAS.n36 CS_BIAS.n22 24.5923
R5987 CS_BIAS.n34 CS_BIAS.n33 24.5923
R5988 CS_BIAS.n29 CS_BIAS.n28 24.5923
R5989 CS_BIAS.n136 CS_BIAS.n135 24.5923
R5990 CS_BIAS.n131 CS_BIAS.n1 24.5923
R5991 CS_BIAS.n129 CS_BIAS.n128 24.5923
R5992 CS_BIAS.n124 CS_BIAS.n123 24.5923
R5993 CS_BIAS.n121 CS_BIAS.n5 24.5923
R5994 CS_BIAS.n116 CS_BIAS.n115 24.5923
R5995 CS_BIAS.n112 CS_BIAS.n111 24.5923
R5996 CS_BIAS.n110 CS_BIAS.n9 24.5923
R5997 CS_BIAS.n106 CS_BIAS.n105 24.5923
R5998 CS_BIAS.n100 CS_BIAS.n86 24.5923
R5999 CS_BIAS.n98 CS_BIAS.n97 24.5923
R6000 CS_BIAS.n93 CS_BIAS.n92 24.5923
R6001 CS_BIAS.n362 CS_BIAS.n361 24.5923
R6002 CS_BIAS.n367 CS_BIAS.n366 24.5923
R6003 CS_BIAS.n369 CS_BIAS.n355 24.5923
R6004 CS_BIAS.n376 CS_BIAS.n374 24.5923
R6005 CS_BIAS.n380 CS_BIAS.n353 24.5923
R6006 CS_BIAS.n382 CS_BIAS.n381 24.5923
R6007 CS_BIAS.n386 CS_BIAS.n385 24.5923
R6008 CS_BIAS.n391 CS_BIAS.n349 24.5923
R6009 CS_BIAS.n394 CS_BIAS.n393 24.5923
R6010 CS_BIAS.n399 CS_BIAS.n398 24.5923
R6011 CS_BIAS.n401 CS_BIAS.n345 24.5923
R6012 CS_BIAS.n406 CS_BIAS.n405 24.5923
R6013 CS_BIAS.n261 CS_BIAS.n260 24.5923
R6014 CS_BIAS.n266 CS_BIAS.n265 24.5923
R6015 CS_BIAS.n268 CS_BIAS.n254 24.5923
R6016 CS_BIAS.n275 CS_BIAS.n273 24.5923
R6017 CS_BIAS.n279 CS_BIAS.n252 24.5923
R6018 CS_BIAS.n281 CS_BIAS.n280 24.5923
R6019 CS_BIAS.n285 CS_BIAS.n284 24.5923
R6020 CS_BIAS.n290 CS_BIAS.n248 24.5923
R6021 CS_BIAS.n293 CS_BIAS.n292 24.5923
R6022 CS_BIAS.n298 CS_BIAS.n297 24.5923
R6023 CS_BIAS.n300 CS_BIAS.n244 24.5923
R6024 CS_BIAS.n305 CS_BIAS.n304 24.5923
R6025 CS_BIAS.n341 CS_BIAS.n340 24.5923
R6026 CS_BIAS.n334 CS_BIAS.n333 24.5923
R6027 CS_BIAS.n336 CS_BIAS.n206 24.5923
R6028 CS_BIAS.n326 CS_BIAS.n210 24.5923
R6029 CS_BIAS.n329 CS_BIAS.n328 24.5923
R6030 CS_BIAS.n317 CS_BIAS.n316 24.5923
R6031 CS_BIAS.n321 CS_BIAS.n320 24.5923
R6032 CS_BIAS.n223 CS_BIAS.n222 24.5923
R6033 CS_BIAS.n228 CS_BIAS.n227 24.5923
R6034 CS_BIAS.n230 CS_BIAS.n216 24.5923
R6035 CS_BIAS.n237 CS_BIAS.n235 24.5923
R6036 CS_BIAS.n315 CS_BIAS.n214 24.5923
R6037 CS_BIAS.n196 CS_BIAS.n195 20.9036
R6038 CS_BIAS.n67 CS_BIAS.n66 20.9036
R6039 CS_BIAS.n131 CS_BIAS.n130 20.9036
R6040 CS_BIAS.n401 CS_BIAS.n400 20.9036
R6041 CS_BIAS.n300 CS_BIAS.n299 20.9036
R6042 CS_BIAS.n336 CS_BIAS.n335 20.9036
R6043 CS_BIAS.n150 CS_BIAS.n148 20.4117
R6044 CS_BIAS.n177 CS_BIAS.n146 20.4117
R6045 CS_BIAS.n48 CS_BIAS.n17 20.4117
R6046 CS_BIAS.n21 CS_BIAS.n19 20.4117
R6047 CS_BIAS.n112 CS_BIAS.n7 20.4117
R6048 CS_BIAS.n85 CS_BIAS.n9 20.4117
R6049 CS_BIAS.n375 CS_BIAS.n353 20.4117
R6050 CS_BIAS.n382 CS_BIAS.n351 20.4117
R6051 CS_BIAS.n274 CS_BIAS.n252 20.4117
R6052 CS_BIAS.n281 CS_BIAS.n250 20.4117
R6053 CS_BIAS.n317 CS_BIAS.n212 20.4117
R6054 CS_BIAS.n236 CS_BIAS.n214 20.4117
R6055 CS_BIAS.n202 CS_BIAS.n201 19.9199
R6056 CS_BIAS.n73 CS_BIAS.n72 19.9199
R6057 CS_BIAS.n137 CS_BIAS.n136 19.9199
R6058 CS_BIAS.n407 CS_BIAS.n406 19.9199
R6059 CS_BIAS.n306 CS_BIAS.n305 19.9199
R6060 CS_BIAS.n342 CS_BIAS.n341 19.9199
R6061 CS_BIAS.n155 CS_BIAS.n154 13.3071
R6062 CS_BIAS.n359 CS_BIAS.n358 13.3071
R6063 CS_BIAS.n258 CS_BIAS.n257 13.3071
R6064 CS_BIAS.n220 CS_BIAS.n219 13.3071
R6065 CS_BIAS.n26 CS_BIAS.n25 13.3071
R6066 CS_BIAS.n90 CS_BIAS.n89 13.3071
R6067 CS_BIAS.n76 CS_BIAS.n74 13.0832
R6068 CS_BIAS.n309 CS_BIAS.n307 13.0832
R6069 CS_BIAS.n164 CS_BIAS.n163 12.5423
R6070 CS_BIAS.n188 CS_BIAS.n187 12.5423
R6071 CS_BIAS.n59 CS_BIAS.n58 12.5423
R6072 CS_BIAS.n35 CS_BIAS.n34 12.5423
R6073 CS_BIAS.n123 CS_BIAS.n122 12.5423
R6074 CS_BIAS.n99 CS_BIAS.n98 12.5423
R6075 CS_BIAS.n368 CS_BIAS.n367 12.5423
R6076 CS_BIAS.n393 CS_BIAS.n392 12.5423
R6077 CS_BIAS.n267 CS_BIAS.n266 12.5423
R6078 CS_BIAS.n292 CS_BIAS.n291 12.5423
R6079 CS_BIAS.n328 CS_BIAS.n327 12.5423
R6080 CS_BIAS.n229 CS_BIAS.n228 12.5423
R6081 CS_BIAS.n165 CS_BIAS.n164 12.0505
R6082 CS_BIAS.n187 CS_BIAS.n186 12.0505
R6083 CS_BIAS.n58 CS_BIAS.n57 12.0505
R6084 CS_BIAS.n36 CS_BIAS.n35 12.0505
R6085 CS_BIAS.n122 CS_BIAS.n121 12.0505
R6086 CS_BIAS.n100 CS_BIAS.n99 12.0505
R6087 CS_BIAS.n369 CS_BIAS.n368 12.0505
R6088 CS_BIAS.n392 CS_BIAS.n391 12.0505
R6089 CS_BIAS.n268 CS_BIAS.n267 12.0505
R6090 CS_BIAS.n291 CS_BIAS.n290 12.0505
R6091 CS_BIAS.n327 CS_BIAS.n326 12.0505
R6092 CS_BIAS.n230 CS_BIAS.n229 12.0505
R6093 CS_BIAS.n410 CS_BIAS.n204 11.3868
R6094 CS_BIAS.n410 CS_BIAS.n409 9.93702
R6095 CS_BIAS.n83 CS_BIAS.n82 9.50363
R6096 CS_BIAS.n313 CS_BIAS.n312 9.50363
R6097 CS_BIAS.n204 CS_BIAS.n138 8.35614
R6098 CS_BIAS.n409 CS_BIAS.n343 8.35614
R6099 CS_BIAS.n204 CS_BIAS.n203 5.04553
R6100 CS_BIAS.n409 CS_BIAS.n408 5.04553
R6101 CS_BIAS.n171 CS_BIAS.n150 4.18111
R6102 CS_BIAS.n180 CS_BIAS.n146 4.18111
R6103 CS_BIAS.n51 CS_BIAS.n17 4.18111
R6104 CS_BIAS.n42 CS_BIAS.n21 4.18111
R6105 CS_BIAS.n115 CS_BIAS.n7 4.18111
R6106 CS_BIAS.n106 CS_BIAS.n85 4.18111
R6107 CS_BIAS.n376 CS_BIAS.n375 4.18111
R6108 CS_BIAS.n385 CS_BIAS.n351 4.18111
R6109 CS_BIAS.n275 CS_BIAS.n274 4.18111
R6110 CS_BIAS.n284 CS_BIAS.n250 4.18111
R6111 CS_BIAS.n320 CS_BIAS.n212 4.18111
R6112 CS_BIAS.n237 CS_BIAS.n236 4.18111
R6113 CS_BIAS CS_BIAS.n410 3.92026
R6114 CS_BIAS.n157 CS_BIAS.n156 3.68928
R6115 CS_BIAS.n195 CS_BIAS.n194 3.68928
R6116 CS_BIAS.n66 CS_BIAS.n65 3.68928
R6117 CS_BIAS.n28 CS_BIAS.n27 3.68928
R6118 CS_BIAS.n130 CS_BIAS.n129 3.68928
R6119 CS_BIAS.n92 CS_BIAS.n91 3.68928
R6120 CS_BIAS.n361 CS_BIAS.n360 3.68928
R6121 CS_BIAS.n400 CS_BIAS.n399 3.68928
R6122 CS_BIAS.n260 CS_BIAS.n259 3.68928
R6123 CS_BIAS.n299 CS_BIAS.n298 3.68928
R6124 CS_BIAS.n335 CS_BIAS.n334 3.68928
R6125 CS_BIAS.n222 CS_BIAS.n221 3.68928
R6126 CS_BIAS.n79 CS_BIAS.t3 3.3005
R6127 CS_BIAS.n79 CS_BIAS.t27 3.3005
R6128 CS_BIAS.n80 CS_BIAS.t1 3.3005
R6129 CS_BIAS.n80 CS_BIAS.t17 3.3005
R6130 CS_BIAS.n77 CS_BIAS.t23 3.3005
R6131 CS_BIAS.n77 CS_BIAS.t19 3.3005
R6132 CS_BIAS.n75 CS_BIAS.t7 3.3005
R6133 CS_BIAS.n75 CS_BIAS.t31 3.3005
R6134 CS_BIAS.n308 CS_BIAS.t5 3.3005
R6135 CS_BIAS.n308 CS_BIAS.t29 3.3005
R6136 CS_BIAS.n310 CS_BIAS.t9 3.3005
R6137 CS_BIAS.n310 CS_BIAS.t11 3.3005
R6138 CS_BIAS.n241 CS_BIAS.t21 3.3005
R6139 CS_BIAS.n241 CS_BIAS.t13 3.3005
R6140 CS_BIAS.n240 CS_BIAS.t25 3.3005
R6141 CS_BIAS.n240 CS_BIAS.t15 3.3005
R6142 CS_BIAS.n78 CS_BIAS.n76 1.00481
R6143 CS_BIAS.n311 CS_BIAS.n309 1.00481
R6144 CS_BIAS.n82 CS_BIAS.n78 0.502655
R6145 CS_BIAS.n82 CS_BIAS.n81 0.502655
R6146 CS_BIAS.n312 CS_BIAS.n242 0.502655
R6147 CS_BIAS.n312 CS_BIAS.n311 0.502655
R6148 CS_BIAS.n203 CS_BIAS.n139 0.278335
R6149 CS_BIAS.n74 CS_BIAS.n10 0.278335
R6150 CS_BIAS.n138 CS_BIAS.n0 0.278335
R6151 CS_BIAS.n408 CS_BIAS.n344 0.278335
R6152 CS_BIAS.n307 CS_BIAS.n243 0.278335
R6153 CS_BIAS.n343 CS_BIAS.n205 0.278335
R6154 CS_BIAS.n199 CS_BIAS.n139 0.189894
R6155 CS_BIAS.n199 CS_BIAS.n198 0.189894
R6156 CS_BIAS.n198 CS_BIAS.n197 0.189894
R6157 CS_BIAS.n197 CS_BIAS.n141 0.189894
R6158 CS_BIAS.n192 CS_BIAS.n141 0.189894
R6159 CS_BIAS.n192 CS_BIAS.n191 0.189894
R6160 CS_BIAS.n191 CS_BIAS.n190 0.189894
R6161 CS_BIAS.n190 CS_BIAS.n143 0.189894
R6162 CS_BIAS.n185 CS_BIAS.n143 0.189894
R6163 CS_BIAS.n185 CS_BIAS.n184 0.189894
R6164 CS_BIAS.n184 CS_BIAS.n183 0.189894
R6165 CS_BIAS.n183 CS_BIAS.n145 0.189894
R6166 CS_BIAS.n179 CS_BIAS.n145 0.189894
R6167 CS_BIAS.n179 CS_BIAS.n178 0.189894
R6168 CS_BIAS.n178 CS_BIAS.n147 0.189894
R6169 CS_BIAS.n174 CS_BIAS.n147 0.189894
R6170 CS_BIAS.n174 CS_BIAS.n173 0.189894
R6171 CS_BIAS.n173 CS_BIAS.n172 0.189894
R6172 CS_BIAS.n172 CS_BIAS.n149 0.189894
R6173 CS_BIAS.n168 CS_BIAS.n149 0.189894
R6174 CS_BIAS.n168 CS_BIAS.n167 0.189894
R6175 CS_BIAS.n167 CS_BIAS.n166 0.189894
R6176 CS_BIAS.n166 CS_BIAS.n152 0.189894
R6177 CS_BIAS.n161 CS_BIAS.n152 0.189894
R6178 CS_BIAS.n161 CS_BIAS.n160 0.189894
R6179 CS_BIAS.n160 CS_BIAS.n159 0.189894
R6180 CS_BIAS.n159 CS_BIAS.n154 0.189894
R6181 CS_BIAS.n70 CS_BIAS.n10 0.189894
R6182 CS_BIAS.n70 CS_BIAS.n69 0.189894
R6183 CS_BIAS.n69 CS_BIAS.n68 0.189894
R6184 CS_BIAS.n68 CS_BIAS.n12 0.189894
R6185 CS_BIAS.n63 CS_BIAS.n12 0.189894
R6186 CS_BIAS.n63 CS_BIAS.n62 0.189894
R6187 CS_BIAS.n62 CS_BIAS.n61 0.189894
R6188 CS_BIAS.n61 CS_BIAS.n14 0.189894
R6189 CS_BIAS.n56 CS_BIAS.n14 0.189894
R6190 CS_BIAS.n56 CS_BIAS.n55 0.189894
R6191 CS_BIAS.n55 CS_BIAS.n54 0.189894
R6192 CS_BIAS.n54 CS_BIAS.n16 0.189894
R6193 CS_BIAS.n50 CS_BIAS.n16 0.189894
R6194 CS_BIAS.n50 CS_BIAS.n49 0.189894
R6195 CS_BIAS.n49 CS_BIAS.n18 0.189894
R6196 CS_BIAS.n45 CS_BIAS.n18 0.189894
R6197 CS_BIAS.n45 CS_BIAS.n44 0.189894
R6198 CS_BIAS.n44 CS_BIAS.n43 0.189894
R6199 CS_BIAS.n43 CS_BIAS.n20 0.189894
R6200 CS_BIAS.n39 CS_BIAS.n20 0.189894
R6201 CS_BIAS.n39 CS_BIAS.n38 0.189894
R6202 CS_BIAS.n38 CS_BIAS.n37 0.189894
R6203 CS_BIAS.n37 CS_BIAS.n23 0.189894
R6204 CS_BIAS.n32 CS_BIAS.n23 0.189894
R6205 CS_BIAS.n32 CS_BIAS.n31 0.189894
R6206 CS_BIAS.n31 CS_BIAS.n30 0.189894
R6207 CS_BIAS.n30 CS_BIAS.n25 0.189894
R6208 CS_BIAS.n109 CS_BIAS.n108 0.189894
R6209 CS_BIAS.n108 CS_BIAS.n107 0.189894
R6210 CS_BIAS.n107 CS_BIAS.n84 0.189894
R6211 CS_BIAS.n103 CS_BIAS.n84 0.189894
R6212 CS_BIAS.n103 CS_BIAS.n102 0.189894
R6213 CS_BIAS.n102 CS_BIAS.n101 0.189894
R6214 CS_BIAS.n101 CS_BIAS.n87 0.189894
R6215 CS_BIAS.n96 CS_BIAS.n87 0.189894
R6216 CS_BIAS.n96 CS_BIAS.n95 0.189894
R6217 CS_BIAS.n95 CS_BIAS.n94 0.189894
R6218 CS_BIAS.n94 CS_BIAS.n89 0.189894
R6219 CS_BIAS.n134 CS_BIAS.n0 0.189894
R6220 CS_BIAS.n134 CS_BIAS.n133 0.189894
R6221 CS_BIAS.n133 CS_BIAS.n132 0.189894
R6222 CS_BIAS.n132 CS_BIAS.n2 0.189894
R6223 CS_BIAS.n127 CS_BIAS.n2 0.189894
R6224 CS_BIAS.n127 CS_BIAS.n126 0.189894
R6225 CS_BIAS.n126 CS_BIAS.n125 0.189894
R6226 CS_BIAS.n125 CS_BIAS.n4 0.189894
R6227 CS_BIAS.n120 CS_BIAS.n4 0.189894
R6228 CS_BIAS.n120 CS_BIAS.n119 0.189894
R6229 CS_BIAS.n119 CS_BIAS.n118 0.189894
R6230 CS_BIAS.n118 CS_BIAS.n6 0.189894
R6231 CS_BIAS.n114 CS_BIAS.n6 0.189894
R6232 CS_BIAS.n114 CS_BIAS.n113 0.189894
R6233 CS_BIAS.n113 CS_BIAS.n8 0.189894
R6234 CS_BIAS.n363 CS_BIAS.n358 0.189894
R6235 CS_BIAS.n364 CS_BIAS.n363 0.189894
R6236 CS_BIAS.n365 CS_BIAS.n364 0.189894
R6237 CS_BIAS.n365 CS_BIAS.n356 0.189894
R6238 CS_BIAS.n370 CS_BIAS.n356 0.189894
R6239 CS_BIAS.n371 CS_BIAS.n370 0.189894
R6240 CS_BIAS.n372 CS_BIAS.n371 0.189894
R6241 CS_BIAS.n372 CS_BIAS.n354 0.189894
R6242 CS_BIAS.n377 CS_BIAS.n354 0.189894
R6243 CS_BIAS.n378 CS_BIAS.n377 0.189894
R6244 CS_BIAS.n379 CS_BIAS.n378 0.189894
R6245 CS_BIAS.n379 CS_BIAS.n352 0.189894
R6246 CS_BIAS.n383 CS_BIAS.n352 0.189894
R6247 CS_BIAS.n384 CS_BIAS.n383 0.189894
R6248 CS_BIAS.n384 CS_BIAS.n350 0.189894
R6249 CS_BIAS.n388 CS_BIAS.n350 0.189894
R6250 CS_BIAS.n389 CS_BIAS.n388 0.189894
R6251 CS_BIAS.n390 CS_BIAS.n389 0.189894
R6252 CS_BIAS.n390 CS_BIAS.n348 0.189894
R6253 CS_BIAS.n395 CS_BIAS.n348 0.189894
R6254 CS_BIAS.n396 CS_BIAS.n395 0.189894
R6255 CS_BIAS.n397 CS_BIAS.n396 0.189894
R6256 CS_BIAS.n397 CS_BIAS.n346 0.189894
R6257 CS_BIAS.n402 CS_BIAS.n346 0.189894
R6258 CS_BIAS.n403 CS_BIAS.n402 0.189894
R6259 CS_BIAS.n404 CS_BIAS.n403 0.189894
R6260 CS_BIAS.n404 CS_BIAS.n344 0.189894
R6261 CS_BIAS.n262 CS_BIAS.n257 0.189894
R6262 CS_BIAS.n263 CS_BIAS.n262 0.189894
R6263 CS_BIAS.n264 CS_BIAS.n263 0.189894
R6264 CS_BIAS.n264 CS_BIAS.n255 0.189894
R6265 CS_BIAS.n269 CS_BIAS.n255 0.189894
R6266 CS_BIAS.n270 CS_BIAS.n269 0.189894
R6267 CS_BIAS.n271 CS_BIAS.n270 0.189894
R6268 CS_BIAS.n271 CS_BIAS.n253 0.189894
R6269 CS_BIAS.n276 CS_BIAS.n253 0.189894
R6270 CS_BIAS.n277 CS_BIAS.n276 0.189894
R6271 CS_BIAS.n278 CS_BIAS.n277 0.189894
R6272 CS_BIAS.n278 CS_BIAS.n251 0.189894
R6273 CS_BIAS.n282 CS_BIAS.n251 0.189894
R6274 CS_BIAS.n283 CS_BIAS.n282 0.189894
R6275 CS_BIAS.n283 CS_BIAS.n249 0.189894
R6276 CS_BIAS.n287 CS_BIAS.n249 0.189894
R6277 CS_BIAS.n288 CS_BIAS.n287 0.189894
R6278 CS_BIAS.n289 CS_BIAS.n288 0.189894
R6279 CS_BIAS.n289 CS_BIAS.n247 0.189894
R6280 CS_BIAS.n294 CS_BIAS.n247 0.189894
R6281 CS_BIAS.n295 CS_BIAS.n294 0.189894
R6282 CS_BIAS.n296 CS_BIAS.n295 0.189894
R6283 CS_BIAS.n296 CS_BIAS.n245 0.189894
R6284 CS_BIAS.n301 CS_BIAS.n245 0.189894
R6285 CS_BIAS.n302 CS_BIAS.n301 0.189894
R6286 CS_BIAS.n303 CS_BIAS.n302 0.189894
R6287 CS_BIAS.n303 CS_BIAS.n243 0.189894
R6288 CS_BIAS.n224 CS_BIAS.n219 0.189894
R6289 CS_BIAS.n225 CS_BIAS.n224 0.189894
R6290 CS_BIAS.n226 CS_BIAS.n225 0.189894
R6291 CS_BIAS.n226 CS_BIAS.n217 0.189894
R6292 CS_BIAS.n231 CS_BIAS.n217 0.189894
R6293 CS_BIAS.n232 CS_BIAS.n231 0.189894
R6294 CS_BIAS.n233 CS_BIAS.n232 0.189894
R6295 CS_BIAS.n233 CS_BIAS.n215 0.189894
R6296 CS_BIAS.n238 CS_BIAS.n215 0.189894
R6297 CS_BIAS.n239 CS_BIAS.n238 0.189894
R6298 CS_BIAS.n314 CS_BIAS.n239 0.189894
R6299 CS_BIAS.n318 CS_BIAS.n213 0.189894
R6300 CS_BIAS.n319 CS_BIAS.n318 0.189894
R6301 CS_BIAS.n319 CS_BIAS.n211 0.189894
R6302 CS_BIAS.n323 CS_BIAS.n211 0.189894
R6303 CS_BIAS.n324 CS_BIAS.n323 0.189894
R6304 CS_BIAS.n325 CS_BIAS.n324 0.189894
R6305 CS_BIAS.n325 CS_BIAS.n209 0.189894
R6306 CS_BIAS.n330 CS_BIAS.n209 0.189894
R6307 CS_BIAS.n331 CS_BIAS.n330 0.189894
R6308 CS_BIAS.n332 CS_BIAS.n331 0.189894
R6309 CS_BIAS.n332 CS_BIAS.n207 0.189894
R6310 CS_BIAS.n337 CS_BIAS.n207 0.189894
R6311 CS_BIAS.n338 CS_BIAS.n337 0.189894
R6312 CS_BIAS.n339 CS_BIAS.n338 0.189894
R6313 CS_BIAS.n339 CS_BIAS.n205 0.189894
R6314 CS_BIAS.n109 CS_BIAS.n83 0.0762576
R6315 CS_BIAS.n83 CS_BIAS.n8 0.0762576
R6316 CS_BIAS.n314 CS_BIAS.n313 0.0762576
R6317 CS_BIAS.n313 CS_BIAS.n213 0.0762576
R6318 GND.n5366 GND.n984 1514.84
R6319 GND.n4838 GND.n4837 1118.08
R6320 GND.n4237 GND.n2044 766.379
R6321 GND.n4239 GND.n2107 766.379
R6322 GND.n3264 GND.n1669 766.379
R6323 GND.n4548 GND.n4547 766.379
R6324 GND.n4964 GND.n1222 766.379
R6325 GND.n5365 GND.n985 766.379
R6326 GND.n5526 GND.n889 766.379
R6327 GND.n2789 GND.n1349 766.379
R6328 GND.n1581 GND.n1528 761.573
R6329 GND.n4585 GND.n1526 761.573
R6330 GND.n2872 GND.n1374 761.573
R6331 GND.n2839 GND.n2838 761.573
R6332 GND.n4307 GND.n2039 761.573
R6333 GND.n3917 GND.n2084 761.573
R6334 GND.n5652 GND.n5651 761.573
R6335 GND.n5714 GND.n709 761.573
R6336 GND.n5712 GND.n742 742.355
R6337 GND.n5657 GND.n5656 742.355
R6338 GND.n2169 GND.n2168 742.355
R6339 GND.n2412 GND.n2411 742.355
R6340 GND.n4684 GND.n1530 742.355
R6341 GND.n4686 GND.n1524 742.355
R6342 GND.n4767 GND.n4766 742.355
R6343 GND.n4835 GND.n1378 742.355
R6344 GND.n4964 GND.n4963 585
R6345 GND.n4965 GND.n4964 585
R6346 GND.n4962 GND.n1224 585
R6347 GND.n1224 GND.n1223 585
R6348 GND.n4961 GND.n4960 585
R6349 GND.n4960 GND.n4959 585
R6350 GND.n1229 GND.n1228 585
R6351 GND.n4958 GND.n1229 585
R6352 GND.n4956 GND.n4955 585
R6353 GND.n4957 GND.n4956 585
R6354 GND.n4954 GND.n1231 585
R6355 GND.n1231 GND.n1230 585
R6356 GND.n4953 GND.n4952 585
R6357 GND.n4952 GND.n4951 585
R6358 GND.n1237 GND.n1236 585
R6359 GND.n4950 GND.n1237 585
R6360 GND.n4948 GND.n4947 585
R6361 GND.n4949 GND.n4948 585
R6362 GND.n4946 GND.n1239 585
R6363 GND.n1239 GND.n1238 585
R6364 GND.n4945 GND.n4944 585
R6365 GND.n4944 GND.n4943 585
R6366 GND.n1245 GND.n1244 585
R6367 GND.n4942 GND.n1245 585
R6368 GND.n4940 GND.n4939 585
R6369 GND.n4941 GND.n4940 585
R6370 GND.n4938 GND.n1247 585
R6371 GND.n1247 GND.n1246 585
R6372 GND.n4937 GND.n4936 585
R6373 GND.n4936 GND.n4935 585
R6374 GND.n1253 GND.n1252 585
R6375 GND.n4934 GND.n1253 585
R6376 GND.n4932 GND.n4931 585
R6377 GND.n4933 GND.n4932 585
R6378 GND.n4930 GND.n1255 585
R6379 GND.n1255 GND.n1254 585
R6380 GND.n4929 GND.n4928 585
R6381 GND.n4928 GND.n4927 585
R6382 GND.n1261 GND.n1260 585
R6383 GND.n4926 GND.n1261 585
R6384 GND.n4924 GND.n4923 585
R6385 GND.n4925 GND.n4924 585
R6386 GND.n4922 GND.n1263 585
R6387 GND.n1263 GND.n1262 585
R6388 GND.n4921 GND.n4920 585
R6389 GND.n4920 GND.n4919 585
R6390 GND.n1269 GND.n1268 585
R6391 GND.n4918 GND.n1269 585
R6392 GND.n4916 GND.n4915 585
R6393 GND.n4917 GND.n4916 585
R6394 GND.n4914 GND.n1271 585
R6395 GND.n1271 GND.n1270 585
R6396 GND.n4913 GND.n4912 585
R6397 GND.n4912 GND.n4911 585
R6398 GND.n1277 GND.n1276 585
R6399 GND.n4910 GND.n1277 585
R6400 GND.n4908 GND.n4907 585
R6401 GND.n4909 GND.n4908 585
R6402 GND.n4906 GND.n1279 585
R6403 GND.n1279 GND.n1278 585
R6404 GND.n4905 GND.n4904 585
R6405 GND.n4904 GND.n4903 585
R6406 GND.n1285 GND.n1284 585
R6407 GND.n4902 GND.n1285 585
R6408 GND.n4900 GND.n4899 585
R6409 GND.n4901 GND.n4900 585
R6410 GND.n4898 GND.n1287 585
R6411 GND.n1287 GND.n1286 585
R6412 GND.n4897 GND.n4896 585
R6413 GND.n4896 GND.n4895 585
R6414 GND.n1293 GND.n1292 585
R6415 GND.n4894 GND.n1293 585
R6416 GND.n4892 GND.n4891 585
R6417 GND.n4893 GND.n4892 585
R6418 GND.n4890 GND.n1295 585
R6419 GND.n1295 GND.n1294 585
R6420 GND.n4889 GND.n4888 585
R6421 GND.n4888 GND.n4887 585
R6422 GND.n1301 GND.n1300 585
R6423 GND.n4886 GND.n1301 585
R6424 GND.n4884 GND.n4883 585
R6425 GND.n4885 GND.n4884 585
R6426 GND.n4882 GND.n1303 585
R6427 GND.n1303 GND.n1302 585
R6428 GND.n4881 GND.n4880 585
R6429 GND.n4880 GND.n4879 585
R6430 GND.n1309 GND.n1308 585
R6431 GND.n4878 GND.n1309 585
R6432 GND.n4876 GND.n4875 585
R6433 GND.n4877 GND.n4876 585
R6434 GND.n4874 GND.n1311 585
R6435 GND.n1311 GND.n1310 585
R6436 GND.n4873 GND.n4872 585
R6437 GND.n4872 GND.n4871 585
R6438 GND.n1317 GND.n1316 585
R6439 GND.n4870 GND.n1317 585
R6440 GND.n4868 GND.n4867 585
R6441 GND.n4869 GND.n4868 585
R6442 GND.n4866 GND.n1319 585
R6443 GND.n1319 GND.n1318 585
R6444 GND.n4865 GND.n4864 585
R6445 GND.n4864 GND.n4863 585
R6446 GND.n1325 GND.n1324 585
R6447 GND.n4862 GND.n1325 585
R6448 GND.n4860 GND.n4859 585
R6449 GND.n4861 GND.n4860 585
R6450 GND.n4858 GND.n1327 585
R6451 GND.n1327 GND.n1326 585
R6452 GND.n4857 GND.n4856 585
R6453 GND.n4856 GND.n4855 585
R6454 GND.n1333 GND.n1332 585
R6455 GND.n4854 GND.n1333 585
R6456 GND.n4852 GND.n4851 585
R6457 GND.n4853 GND.n4852 585
R6458 GND.n4850 GND.n1335 585
R6459 GND.n1335 GND.n1334 585
R6460 GND.n4849 GND.n4848 585
R6461 GND.n4848 GND.n4847 585
R6462 GND.n1341 GND.n1340 585
R6463 GND.n4846 GND.n1341 585
R6464 GND.n4844 GND.n4843 585
R6465 GND.n4845 GND.n4844 585
R6466 GND.n4842 GND.n1343 585
R6467 GND.n1343 GND.n1342 585
R6468 GND.n4841 GND.n4840 585
R6469 GND.n4840 GND.n4839 585
R6470 GND.n1349 GND.n1348 585
R6471 GND.n4838 GND.n1349 585
R6472 GND.n1222 GND.n1221 585
R6473 GND.n4966 GND.n1222 585
R6474 GND.n4969 GND.n4968 585
R6475 GND.n4968 GND.n4967 585
R6476 GND.n1219 GND.n1218 585
R6477 GND.n1218 GND.n1217 585
R6478 GND.n4974 GND.n4973 585
R6479 GND.n4975 GND.n4974 585
R6480 GND.n1216 GND.n1215 585
R6481 GND.n4976 GND.n1216 585
R6482 GND.n4979 GND.n4978 585
R6483 GND.n4978 GND.n4977 585
R6484 GND.n1213 GND.n1212 585
R6485 GND.n1212 GND.n1211 585
R6486 GND.n4984 GND.n4983 585
R6487 GND.n4985 GND.n4984 585
R6488 GND.n1210 GND.n1209 585
R6489 GND.n4986 GND.n1210 585
R6490 GND.n4989 GND.n4988 585
R6491 GND.n4988 GND.n4987 585
R6492 GND.n1207 GND.n1206 585
R6493 GND.n1206 GND.n1205 585
R6494 GND.n4994 GND.n4993 585
R6495 GND.n4995 GND.n4994 585
R6496 GND.n1204 GND.n1203 585
R6497 GND.n4996 GND.n1204 585
R6498 GND.n4999 GND.n4998 585
R6499 GND.n4998 GND.n4997 585
R6500 GND.n1201 GND.n1200 585
R6501 GND.n1200 GND.n1199 585
R6502 GND.n5004 GND.n5003 585
R6503 GND.n5005 GND.n5004 585
R6504 GND.n1198 GND.n1197 585
R6505 GND.n5006 GND.n1198 585
R6506 GND.n5009 GND.n5008 585
R6507 GND.n5008 GND.n5007 585
R6508 GND.n1195 GND.n1194 585
R6509 GND.n1194 GND.n1193 585
R6510 GND.n5014 GND.n5013 585
R6511 GND.n5015 GND.n5014 585
R6512 GND.n1192 GND.n1191 585
R6513 GND.n5016 GND.n1192 585
R6514 GND.n5019 GND.n5018 585
R6515 GND.n5018 GND.n5017 585
R6516 GND.n1189 GND.n1188 585
R6517 GND.n1188 GND.n1187 585
R6518 GND.n5024 GND.n5023 585
R6519 GND.n5025 GND.n5024 585
R6520 GND.n1186 GND.n1185 585
R6521 GND.n5026 GND.n1186 585
R6522 GND.n5029 GND.n5028 585
R6523 GND.n5028 GND.n5027 585
R6524 GND.n1183 GND.n1182 585
R6525 GND.n1182 GND.n1181 585
R6526 GND.n5034 GND.n5033 585
R6527 GND.n5035 GND.n5034 585
R6528 GND.n1180 GND.n1179 585
R6529 GND.n5036 GND.n1180 585
R6530 GND.n5039 GND.n5038 585
R6531 GND.n5038 GND.n5037 585
R6532 GND.n1177 GND.n1176 585
R6533 GND.n1176 GND.n1175 585
R6534 GND.n5044 GND.n5043 585
R6535 GND.n5045 GND.n5044 585
R6536 GND.n1174 GND.n1173 585
R6537 GND.n5046 GND.n1174 585
R6538 GND.n5049 GND.n5048 585
R6539 GND.n5048 GND.n5047 585
R6540 GND.n1171 GND.n1170 585
R6541 GND.n1170 GND.n1169 585
R6542 GND.n5054 GND.n5053 585
R6543 GND.n5055 GND.n5054 585
R6544 GND.n1168 GND.n1167 585
R6545 GND.n5056 GND.n1168 585
R6546 GND.n5059 GND.n5058 585
R6547 GND.n5058 GND.n5057 585
R6548 GND.n1165 GND.n1164 585
R6549 GND.n1164 GND.n1163 585
R6550 GND.n5064 GND.n5063 585
R6551 GND.n5065 GND.n5064 585
R6552 GND.n1162 GND.n1161 585
R6553 GND.n5066 GND.n1162 585
R6554 GND.n5069 GND.n5068 585
R6555 GND.n5068 GND.n5067 585
R6556 GND.n1159 GND.n1158 585
R6557 GND.n1158 GND.n1157 585
R6558 GND.n5074 GND.n5073 585
R6559 GND.n5075 GND.n5074 585
R6560 GND.n1156 GND.n1155 585
R6561 GND.n5076 GND.n1156 585
R6562 GND.n5079 GND.n5078 585
R6563 GND.n5078 GND.n5077 585
R6564 GND.n1153 GND.n1152 585
R6565 GND.n1152 GND.n1151 585
R6566 GND.n5084 GND.n5083 585
R6567 GND.n5085 GND.n5084 585
R6568 GND.n1150 GND.n1149 585
R6569 GND.n5086 GND.n1150 585
R6570 GND.n5089 GND.n5088 585
R6571 GND.n5088 GND.n5087 585
R6572 GND.n1147 GND.n1146 585
R6573 GND.n1146 GND.n1145 585
R6574 GND.n5094 GND.n5093 585
R6575 GND.n5095 GND.n5094 585
R6576 GND.n1144 GND.n1143 585
R6577 GND.n5096 GND.n1144 585
R6578 GND.n5099 GND.n5098 585
R6579 GND.n5098 GND.n5097 585
R6580 GND.n1141 GND.n1140 585
R6581 GND.n1140 GND.n1139 585
R6582 GND.n5104 GND.n5103 585
R6583 GND.n5105 GND.n5104 585
R6584 GND.n1138 GND.n1137 585
R6585 GND.n5106 GND.n1138 585
R6586 GND.n5109 GND.n5108 585
R6587 GND.n5108 GND.n5107 585
R6588 GND.n1135 GND.n1134 585
R6589 GND.n1134 GND.n1133 585
R6590 GND.n5114 GND.n5113 585
R6591 GND.n5115 GND.n5114 585
R6592 GND.n1132 GND.n1131 585
R6593 GND.n5116 GND.n1132 585
R6594 GND.n5119 GND.n5118 585
R6595 GND.n5118 GND.n5117 585
R6596 GND.n1129 GND.n1128 585
R6597 GND.n1128 GND.n1127 585
R6598 GND.n5124 GND.n5123 585
R6599 GND.n5125 GND.n5124 585
R6600 GND.n1126 GND.n1125 585
R6601 GND.n5126 GND.n1126 585
R6602 GND.n5129 GND.n5128 585
R6603 GND.n5128 GND.n5127 585
R6604 GND.n1123 GND.n1122 585
R6605 GND.n1122 GND.n1121 585
R6606 GND.n5134 GND.n5133 585
R6607 GND.n5135 GND.n5134 585
R6608 GND.n1120 GND.n1119 585
R6609 GND.n5136 GND.n1120 585
R6610 GND.n5139 GND.n5138 585
R6611 GND.n5138 GND.n5137 585
R6612 GND.n1117 GND.n1116 585
R6613 GND.n1116 GND.n1115 585
R6614 GND.n5144 GND.n5143 585
R6615 GND.n5145 GND.n5144 585
R6616 GND.n1114 GND.n1113 585
R6617 GND.n5146 GND.n1114 585
R6618 GND.n5149 GND.n5148 585
R6619 GND.n5148 GND.n5147 585
R6620 GND.n1111 GND.n1110 585
R6621 GND.n1110 GND.n1109 585
R6622 GND.n5154 GND.n5153 585
R6623 GND.n5155 GND.n5154 585
R6624 GND.n1108 GND.n1107 585
R6625 GND.n5156 GND.n1108 585
R6626 GND.n5159 GND.n5158 585
R6627 GND.n5158 GND.n5157 585
R6628 GND.n1105 GND.n1104 585
R6629 GND.n1104 GND.n1103 585
R6630 GND.n5164 GND.n5163 585
R6631 GND.n5165 GND.n5164 585
R6632 GND.n1102 GND.n1101 585
R6633 GND.n5166 GND.n1102 585
R6634 GND.n5169 GND.n5168 585
R6635 GND.n5168 GND.n5167 585
R6636 GND.n1099 GND.n1098 585
R6637 GND.n1098 GND.n1097 585
R6638 GND.n5174 GND.n5173 585
R6639 GND.n5175 GND.n5174 585
R6640 GND.n1096 GND.n1095 585
R6641 GND.n5176 GND.n1096 585
R6642 GND.n5179 GND.n5178 585
R6643 GND.n5178 GND.n5177 585
R6644 GND.n1093 GND.n1092 585
R6645 GND.n1092 GND.n1091 585
R6646 GND.n5184 GND.n5183 585
R6647 GND.n5185 GND.n5184 585
R6648 GND.n1090 GND.n1089 585
R6649 GND.n5186 GND.n1090 585
R6650 GND.n5189 GND.n5188 585
R6651 GND.n5188 GND.n5187 585
R6652 GND.n1087 GND.n1086 585
R6653 GND.n1086 GND.n1085 585
R6654 GND.n5194 GND.n5193 585
R6655 GND.n5195 GND.n5194 585
R6656 GND.n1084 GND.n1083 585
R6657 GND.n5196 GND.n1084 585
R6658 GND.n5199 GND.n5198 585
R6659 GND.n5198 GND.n5197 585
R6660 GND.n1081 GND.n1080 585
R6661 GND.n1080 GND.n1079 585
R6662 GND.n5204 GND.n5203 585
R6663 GND.n5205 GND.n5204 585
R6664 GND.n1078 GND.n1077 585
R6665 GND.n5206 GND.n1078 585
R6666 GND.n5209 GND.n5208 585
R6667 GND.n5208 GND.n5207 585
R6668 GND.n1075 GND.n1074 585
R6669 GND.n1074 GND.n1073 585
R6670 GND.n5214 GND.n5213 585
R6671 GND.n5215 GND.n5214 585
R6672 GND.n1072 GND.n1071 585
R6673 GND.n5216 GND.n1072 585
R6674 GND.n5219 GND.n5218 585
R6675 GND.n5218 GND.n5217 585
R6676 GND.n1069 GND.n1068 585
R6677 GND.n1068 GND.n1067 585
R6678 GND.n5224 GND.n5223 585
R6679 GND.n5225 GND.n5224 585
R6680 GND.n1066 GND.n1065 585
R6681 GND.n5226 GND.n1066 585
R6682 GND.n5229 GND.n5228 585
R6683 GND.n5228 GND.n5227 585
R6684 GND.n1063 GND.n1062 585
R6685 GND.n1062 GND.n1061 585
R6686 GND.n5234 GND.n5233 585
R6687 GND.n5235 GND.n5234 585
R6688 GND.n1060 GND.n1059 585
R6689 GND.n5236 GND.n1060 585
R6690 GND.n5239 GND.n5238 585
R6691 GND.n5238 GND.n5237 585
R6692 GND.n1057 GND.n1056 585
R6693 GND.n1056 GND.n1055 585
R6694 GND.n5244 GND.n5243 585
R6695 GND.n5245 GND.n5244 585
R6696 GND.n1054 GND.n1053 585
R6697 GND.n5246 GND.n1054 585
R6698 GND.n5249 GND.n5248 585
R6699 GND.n5248 GND.n5247 585
R6700 GND.n1051 GND.n1050 585
R6701 GND.n1050 GND.n1049 585
R6702 GND.n5254 GND.n5253 585
R6703 GND.n5255 GND.n5254 585
R6704 GND.n1048 GND.n1047 585
R6705 GND.n5256 GND.n1048 585
R6706 GND.n5259 GND.n5258 585
R6707 GND.n5258 GND.n5257 585
R6708 GND.n1045 GND.n1044 585
R6709 GND.n1044 GND.n1043 585
R6710 GND.n5264 GND.n5263 585
R6711 GND.n5265 GND.n5264 585
R6712 GND.n1042 GND.n1041 585
R6713 GND.n5266 GND.n1042 585
R6714 GND.n5269 GND.n5268 585
R6715 GND.n5268 GND.n5267 585
R6716 GND.n1039 GND.n1038 585
R6717 GND.n1038 GND.n1037 585
R6718 GND.n5274 GND.n5273 585
R6719 GND.n5275 GND.n5274 585
R6720 GND.n1036 GND.n1035 585
R6721 GND.n5276 GND.n1036 585
R6722 GND.n5279 GND.n5278 585
R6723 GND.n5278 GND.n5277 585
R6724 GND.n1033 GND.n1032 585
R6725 GND.n1032 GND.n1031 585
R6726 GND.n5284 GND.n5283 585
R6727 GND.n5285 GND.n5284 585
R6728 GND.n1030 GND.n1029 585
R6729 GND.n5286 GND.n1030 585
R6730 GND.n5289 GND.n5288 585
R6731 GND.n5288 GND.n5287 585
R6732 GND.n1027 GND.n1026 585
R6733 GND.n1026 GND.n1025 585
R6734 GND.n5294 GND.n5293 585
R6735 GND.n5295 GND.n5294 585
R6736 GND.n1024 GND.n1023 585
R6737 GND.n5296 GND.n1024 585
R6738 GND.n5299 GND.n5298 585
R6739 GND.n5298 GND.n5297 585
R6740 GND.n1021 GND.n1020 585
R6741 GND.n1020 GND.n1019 585
R6742 GND.n5304 GND.n5303 585
R6743 GND.n5305 GND.n5304 585
R6744 GND.n1018 GND.n1017 585
R6745 GND.n5306 GND.n1018 585
R6746 GND.n5309 GND.n5308 585
R6747 GND.n5308 GND.n5307 585
R6748 GND.n1015 GND.n1014 585
R6749 GND.n1014 GND.n1013 585
R6750 GND.n5314 GND.n5313 585
R6751 GND.n5315 GND.n5314 585
R6752 GND.n1012 GND.n1011 585
R6753 GND.n5316 GND.n1012 585
R6754 GND.n5319 GND.n5318 585
R6755 GND.n5318 GND.n5317 585
R6756 GND.n1009 GND.n1008 585
R6757 GND.n1008 GND.n1007 585
R6758 GND.n5324 GND.n5323 585
R6759 GND.n5325 GND.n5324 585
R6760 GND.n1006 GND.n1005 585
R6761 GND.n5326 GND.n1006 585
R6762 GND.n5329 GND.n5328 585
R6763 GND.n5328 GND.n5327 585
R6764 GND.n1003 GND.n1002 585
R6765 GND.n1002 GND.n1001 585
R6766 GND.n5334 GND.n5333 585
R6767 GND.n5335 GND.n5334 585
R6768 GND.n1000 GND.n999 585
R6769 GND.n5336 GND.n1000 585
R6770 GND.n5339 GND.n5338 585
R6771 GND.n5338 GND.n5337 585
R6772 GND.n997 GND.n996 585
R6773 GND.n996 GND.n995 585
R6774 GND.n5344 GND.n5343 585
R6775 GND.n5345 GND.n5344 585
R6776 GND.n994 GND.n993 585
R6777 GND.n5346 GND.n994 585
R6778 GND.n5349 GND.n5348 585
R6779 GND.n5348 GND.n5347 585
R6780 GND.n991 GND.n990 585
R6781 GND.n990 GND.n989 585
R6782 GND.n5355 GND.n5354 585
R6783 GND.n5356 GND.n5355 585
R6784 GND.n988 GND.n987 585
R6785 GND.n5357 GND.n988 585
R6786 GND.n5360 GND.n5359 585
R6787 GND.n5359 GND.n5358 585
R6788 GND.n5361 GND.n985 585
R6789 GND.n985 GND.n984 585
R6790 GND.n5522 GND.n889 585
R6791 GND.n889 GND.n724 585
R6792 GND.n5521 GND.n5520 585
R6793 GND.n5520 GND.n5519 585
R6794 GND.n893 GND.n892 585
R6795 GND.n5518 GND.n893 585
R6796 GND.n5516 GND.n5515 585
R6797 GND.n5517 GND.n5516 585
R6798 GND.n896 GND.n895 585
R6799 GND.n895 GND.n894 585
R6800 GND.n5510 GND.n5509 585
R6801 GND.n5509 GND.n5508 585
R6802 GND.n899 GND.n898 585
R6803 GND.n5507 GND.n899 585
R6804 GND.n5505 GND.n5504 585
R6805 GND.n5506 GND.n5505 585
R6806 GND.n902 GND.n901 585
R6807 GND.n901 GND.n900 585
R6808 GND.n5500 GND.n5499 585
R6809 GND.n5499 GND.n5498 585
R6810 GND.n905 GND.n904 585
R6811 GND.n5497 GND.n905 585
R6812 GND.n5495 GND.n5494 585
R6813 GND.n5496 GND.n5495 585
R6814 GND.n908 GND.n907 585
R6815 GND.n907 GND.n906 585
R6816 GND.n5490 GND.n5489 585
R6817 GND.n5489 GND.n5488 585
R6818 GND.n911 GND.n910 585
R6819 GND.n5487 GND.n911 585
R6820 GND.n5485 GND.n5484 585
R6821 GND.n5486 GND.n5485 585
R6822 GND.n914 GND.n913 585
R6823 GND.n913 GND.n912 585
R6824 GND.n5480 GND.n5479 585
R6825 GND.n5479 GND.n5478 585
R6826 GND.n917 GND.n916 585
R6827 GND.n5477 GND.n917 585
R6828 GND.n5475 GND.n5474 585
R6829 GND.n5476 GND.n5475 585
R6830 GND.n920 GND.n919 585
R6831 GND.n919 GND.n918 585
R6832 GND.n5470 GND.n5469 585
R6833 GND.n5469 GND.n5468 585
R6834 GND.n923 GND.n922 585
R6835 GND.n5467 GND.n923 585
R6836 GND.n5465 GND.n5464 585
R6837 GND.n5466 GND.n5465 585
R6838 GND.n926 GND.n925 585
R6839 GND.n925 GND.n924 585
R6840 GND.n5460 GND.n5459 585
R6841 GND.n5459 GND.n5458 585
R6842 GND.n929 GND.n928 585
R6843 GND.n5457 GND.n929 585
R6844 GND.n5455 GND.n5454 585
R6845 GND.n5456 GND.n5455 585
R6846 GND.n932 GND.n931 585
R6847 GND.n931 GND.n930 585
R6848 GND.n5450 GND.n5449 585
R6849 GND.n5449 GND.n5448 585
R6850 GND.n935 GND.n934 585
R6851 GND.n5447 GND.n935 585
R6852 GND.n5445 GND.n5444 585
R6853 GND.n5446 GND.n5445 585
R6854 GND.n938 GND.n937 585
R6855 GND.n937 GND.n936 585
R6856 GND.n5440 GND.n5439 585
R6857 GND.n5439 GND.n5438 585
R6858 GND.n941 GND.n940 585
R6859 GND.n5437 GND.n941 585
R6860 GND.n5435 GND.n5434 585
R6861 GND.n5436 GND.n5435 585
R6862 GND.n944 GND.n943 585
R6863 GND.n943 GND.n942 585
R6864 GND.n5430 GND.n5429 585
R6865 GND.n5429 GND.n5428 585
R6866 GND.n947 GND.n946 585
R6867 GND.n5427 GND.n947 585
R6868 GND.n5425 GND.n5424 585
R6869 GND.n5426 GND.n5425 585
R6870 GND.n950 GND.n949 585
R6871 GND.n949 GND.n948 585
R6872 GND.n5420 GND.n5419 585
R6873 GND.n5419 GND.n5418 585
R6874 GND.n953 GND.n952 585
R6875 GND.n5417 GND.n953 585
R6876 GND.n5415 GND.n5414 585
R6877 GND.n5416 GND.n5415 585
R6878 GND.n956 GND.n955 585
R6879 GND.n955 GND.n954 585
R6880 GND.n5410 GND.n5409 585
R6881 GND.n5409 GND.n5408 585
R6882 GND.n959 GND.n958 585
R6883 GND.n5407 GND.n959 585
R6884 GND.n5405 GND.n5404 585
R6885 GND.n5406 GND.n5405 585
R6886 GND.n962 GND.n961 585
R6887 GND.n961 GND.n960 585
R6888 GND.n5400 GND.n5399 585
R6889 GND.n5399 GND.n5398 585
R6890 GND.n965 GND.n964 585
R6891 GND.n5397 GND.n965 585
R6892 GND.n5395 GND.n5394 585
R6893 GND.n5396 GND.n5395 585
R6894 GND.n968 GND.n967 585
R6895 GND.n967 GND.n966 585
R6896 GND.n5390 GND.n5389 585
R6897 GND.n5389 GND.n5388 585
R6898 GND.n971 GND.n970 585
R6899 GND.n5387 GND.n971 585
R6900 GND.n5385 GND.n5384 585
R6901 GND.n5386 GND.n5385 585
R6902 GND.n974 GND.n973 585
R6903 GND.n973 GND.n972 585
R6904 GND.n5380 GND.n5379 585
R6905 GND.n5379 GND.n5378 585
R6906 GND.n977 GND.n976 585
R6907 GND.n5377 GND.n977 585
R6908 GND.n5375 GND.n5374 585
R6909 GND.n5376 GND.n5375 585
R6910 GND.n980 GND.n979 585
R6911 GND.n979 GND.n978 585
R6912 GND.n5370 GND.n5369 585
R6913 GND.n5369 GND.n5368 585
R6914 GND.n983 GND.n982 585
R6915 GND.n5367 GND.n983 585
R6916 GND.n5365 GND.n5364 585
R6917 GND.n5366 GND.n5365 585
R6918 GND.n4237 GND.n4236 585
R6919 GND.n4238 GND.n4237 585
R6920 GND.n2111 GND.n2110 585
R6921 GND.n3871 GND.n2110 585
R6922 GND.n3869 GND.n3868 585
R6923 GND.n3870 GND.n3869 585
R6924 GND.n2431 GND.n2430 585
R6925 GND.n2438 GND.n2430 585
R6926 GND.n3864 GND.n3863 585
R6927 GND.n3863 GND.n3862 585
R6928 GND.n2434 GND.n2433 585
R6929 GND.n3852 GND.n2434 585
R6930 GND.n3835 GND.n2454 585
R6931 GND.n2454 GND.n2444 585
R6932 GND.n3837 GND.n3836 585
R6933 GND.n3838 GND.n3837 585
R6934 GND.n2455 GND.n2453 585
R6935 GND.n2460 GND.n2453 585
R6936 GND.n3830 GND.n3829 585
R6937 GND.n3829 GND.n3828 585
R6938 GND.n2458 GND.n2457 585
R6939 GND.n3816 GND.n2458 585
R6940 GND.n3803 GND.n3788 585
R6941 GND.n3788 GND.n2471 585
R6942 GND.n3805 GND.n3804 585
R6943 GND.n3806 GND.n3805 585
R6944 GND.n3789 GND.n3787 585
R6945 GND.n3787 GND.n3786 585
R6946 GND.n3798 GND.n3797 585
R6947 GND.n3797 GND.n1944 585
R6948 GND.n3796 GND.n3791 585
R6949 GND.n3796 GND.n1942 585
R6950 GND.n3795 GND.n3794 585
R6951 GND.n3795 GND.n1928 585
R6952 GND.n1916 GND.n1915 585
R6953 GND.n1926 GND.n1916 585
R6954 GND.n4395 GND.n4394 585
R6955 GND.n4394 GND.n4393 585
R6956 GND.n4396 GND.n1910 585
R6957 GND.n3706 GND.n1910 585
R6958 GND.n4398 GND.n4397 585
R6959 GND.n4399 GND.n4398 585
R6960 GND.n1911 GND.n1909 585
R6961 GND.n3685 GND.n1909 585
R6962 GND.n2494 GND.n2493 585
R6963 GND.n2495 GND.n2494 585
R6964 GND.n1878 GND.n1877 585
R6965 GND.n1888 GND.n1878 585
R6966 GND.n4415 GND.n4414 585
R6967 GND.n4414 GND.n4413 585
R6968 GND.n4416 GND.n1867 585
R6969 GND.n3661 GND.n1867 585
R6970 GND.n4418 GND.n4417 585
R6971 GND.n4419 GND.n4418 585
R6972 GND.n1868 GND.n1866 585
R6973 GND.n1866 GND.n1856 585
R6974 GND.n1871 GND.n1870 585
R6975 GND.n1870 GND.n1854 585
R6976 GND.n1843 GND.n1842 585
R6977 GND.n3647 GND.n1843 585
R6978 GND.n4436 GND.n4435 585
R6979 GND.n4435 GND.n4434 585
R6980 GND.n4437 GND.n1837 585
R6981 GND.n3623 GND.n1837 585
R6982 GND.n4439 GND.n4438 585
R6983 GND.n4440 GND.n4439 585
R6984 GND.n1823 GND.n1822 585
R6985 GND.n3612 GND.n1823 585
R6986 GND.n4450 GND.n4449 585
R6987 GND.n4449 GND.n4448 585
R6988 GND.n4451 GND.n1817 585
R6989 GND.n3557 GND.n1817 585
R6990 GND.n4453 GND.n4452 585
R6991 GND.n4454 GND.n4453 585
R6992 GND.n1805 GND.n1804 585
R6993 GND.n3582 GND.n1805 585
R6994 GND.n4464 GND.n4463 585
R6995 GND.n4463 GND.n4462 585
R6996 GND.n4465 GND.n1799 585
R6997 GND.n3568 GND.n1799 585
R6998 GND.n4467 GND.n4466 585
R6999 GND.n4468 GND.n4467 585
R7000 GND.n1785 GND.n1784 585
R7001 GND.n3549 GND.n1785 585
R7002 GND.n4478 GND.n4477 585
R7003 GND.n4477 GND.n4476 585
R7004 GND.n4479 GND.n1779 585
R7005 GND.n3537 GND.n1779 585
R7006 GND.n4481 GND.n4480 585
R7007 GND.n4482 GND.n4481 585
R7008 GND.n1765 GND.n1764 585
R7009 GND.n3504 GND.n1765 585
R7010 GND.n4492 GND.n4491 585
R7011 GND.n4491 GND.n4490 585
R7012 GND.n4493 GND.n1759 585
R7013 GND.n3515 GND.n1759 585
R7014 GND.n4495 GND.n4494 585
R7015 GND.n4496 GND.n4495 585
R7016 GND.n1745 GND.n1744 585
R7017 GND.n3488 GND.n1745 585
R7018 GND.n4506 GND.n4505 585
R7019 GND.n4505 GND.n4504 585
R7020 GND.n4507 GND.n1737 585
R7021 GND.n3480 GND.n1737 585
R7022 GND.n4509 GND.n4508 585
R7023 GND.n4510 GND.n4509 585
R7024 GND.n1738 GND.n1736 585
R7025 GND.n2575 GND.n1736 585
R7026 GND.n1720 GND.n1719 585
R7027 GND.n1723 GND.n1720 585
R7028 GND.n4520 GND.n4519 585
R7029 GND.n4519 GND.n4518 585
R7030 GND.n4521 GND.n1712 585
R7031 GND.n3287 GND.n1712 585
R7032 GND.n4523 GND.n4522 585
R7033 GND.n4524 GND.n4523 585
R7034 GND.n1713 GND.n1711 585
R7035 GND.n1711 GND.n1708 585
R7036 GND.n1693 GND.n1692 585
R7037 GND.n1696 GND.n1693 585
R7038 GND.n4534 GND.n4533 585
R7039 GND.n4533 GND.n4532 585
R7040 GND.n4535 GND.n1684 585
R7041 GND.n2581 GND.n1684 585
R7042 GND.n4537 GND.n4536 585
R7043 GND.n4538 GND.n4537 585
R7044 GND.n1685 GND.n1683 585
R7045 GND.n3272 GND.n1683 585
R7046 GND.n1686 GND.n1666 585
R7047 GND.n1670 GND.n1666 585
R7048 GND.n4547 GND.n1667 585
R7049 GND.n4547 GND.n4546 585
R7050 GND.n4548 GND.n1587 585
R7051 GND.n4622 GND.n1588 585
R7052 GND.n4621 GND.n1589 585
R7053 GND.n4550 GND.n1589 585
R7054 GND.n1648 GND.n1590 585
R7055 GND.n4614 GND.n1596 585
R7056 GND.n4613 GND.n1597 585
R7057 GND.n1650 GND.n1598 585
R7058 GND.n4606 GND.n1604 585
R7059 GND.n4605 GND.n1605 585
R7060 GND.n1653 GND.n1606 585
R7061 GND.n4598 GND.n1612 585
R7062 GND.n4597 GND.n1613 585
R7063 GND.n1655 GND.n1614 585
R7064 GND.n4590 GND.n1622 585
R7065 GND.n4589 GND.n1623 585
R7066 GND.n1658 GND.n1624 585
R7067 GND.n3238 GND.n3237 585
R7068 GND.n3240 GND.n3239 585
R7069 GND.n3243 GND.n3242 585
R7070 GND.n3241 GND.n2587 585
R7071 GND.n3248 GND.n3247 585
R7072 GND.n3250 GND.n3249 585
R7073 GND.n3256 GND.n3252 585
R7074 GND.n3251 GND.n2585 585
R7075 GND.n3261 GND.n3260 585
R7076 GND.n3263 GND.n3262 585
R7077 GND.n3265 GND.n3264 585
R7078 GND.n2107 GND.n2103 585
R7079 GND.n4244 GND.n2102 585
R7080 GND.n4245 GND.n2101 585
R7081 GND.n4246 GND.n2100 585
R7082 GND.n3884 GND.n2095 585
R7083 GND.n4250 GND.n2094 585
R7084 GND.n4251 GND.n2093 585
R7085 GND.n4252 GND.n2092 585
R7086 GND.n3887 GND.n2089 585
R7087 GND.n4256 GND.n2088 585
R7088 GND.n4257 GND.n2087 585
R7089 GND.n4258 GND.n2086 585
R7090 GND.n3890 GND.n2082 585
R7091 GND.n4269 GND.n2081 585
R7092 GND.n4270 GND.n2080 585
R7093 GND.n3892 GND.n2074 585
R7094 GND.n4277 GND.n2073 585
R7095 GND.n4278 GND.n2072 585
R7096 GND.n3895 GND.n2064 585
R7097 GND.n4285 GND.n2063 585
R7098 GND.n4286 GND.n2062 585
R7099 GND.n3897 GND.n2056 585
R7100 GND.n4293 GND.n2055 585
R7101 GND.n4294 GND.n2054 585
R7102 GND.n3900 GND.n2046 585
R7103 GND.n4301 GND.n2045 585
R7104 GND.n4302 GND.n2044 585
R7105 GND.n3902 GND.n2044 585
R7106 GND.n4240 GND.n4239 585
R7107 GND.n4239 GND.n4238 585
R7108 GND.n2106 GND.n2105 585
R7109 GND.n3871 GND.n2106 585
R7110 GND.n3845 GND.n2429 585
R7111 GND.n3870 GND.n2429 585
R7112 GND.n3846 GND.n3844 585
R7113 GND.n3844 GND.n2438 585
R7114 GND.n2447 GND.n2436 585
R7115 GND.n3862 GND.n2436 585
R7116 GND.n3851 GND.n3850 585
R7117 GND.n3852 GND.n3851 585
R7118 GND.n2446 GND.n2445 585
R7119 GND.n2445 GND.n2444 585
R7120 GND.n3840 GND.n3839 585
R7121 GND.n3839 GND.n3838 585
R7122 GND.n2450 GND.n2449 585
R7123 GND.n2460 GND.n2450 585
R7124 GND.n2474 GND.n2459 585
R7125 GND.n3828 GND.n2459 585
R7126 GND.n3814 GND.n3813 585
R7127 GND.n3816 GND.n3814 585
R7128 GND.n2473 GND.n2472 585
R7129 GND.n2472 GND.n2471 585
R7130 GND.n3808 GND.n3807 585
R7131 GND.n3807 GND.n3806 585
R7132 GND.n2477 GND.n2476 585
R7133 GND.n3786 GND.n2477 585
R7134 GND.n3695 GND.n3694 585
R7135 GND.n3694 GND.n1944 585
R7136 GND.n3698 GND.n3693 585
R7137 GND.n3693 GND.n1942 585
R7138 GND.n3699 GND.n3692 585
R7139 GND.n3692 GND.n1928 585
R7140 GND.n3700 GND.n3691 585
R7141 GND.n3691 GND.n1926 585
R7142 GND.n2485 GND.n1918 585
R7143 GND.n4393 GND.n1918 585
R7144 GND.n3705 GND.n3704 585
R7145 GND.n3706 GND.n3705 585
R7146 GND.n2484 GND.n1907 585
R7147 GND.n4399 GND.n1907 585
R7148 GND.n3687 GND.n3686 585
R7149 GND.n3686 GND.n3685 585
R7150 GND.n2488 GND.n2487 585
R7151 GND.n2495 GND.n2488 585
R7152 GND.n3655 GND.n3654 585
R7153 GND.n3654 GND.n1888 585
R7154 GND.n2503 GND.n1881 585
R7155 GND.n4413 GND.n1881 585
R7156 GND.n3660 GND.n3659 585
R7157 GND.n3661 GND.n3660 585
R7158 GND.n2502 GND.n1864 585
R7159 GND.n4419 GND.n1864 585
R7160 GND.n3651 GND.n3650 585
R7161 GND.n3650 GND.n1856 585
R7162 GND.n3649 GND.n2505 585
R7163 GND.n3649 GND.n1854 585
R7164 GND.n3648 GND.n2506 585
R7165 GND.n3648 GND.n3647 585
R7166 GND.n2517 GND.n1844 585
R7167 GND.n4434 GND.n1844 585
R7168 GND.n3621 GND.n3620 585
R7169 GND.n3623 GND.n3621 585
R7170 GND.n2516 GND.n1835 585
R7171 GND.n4440 GND.n1835 585
R7172 GND.n3614 GND.n3613 585
R7173 GND.n3613 GND.n3612 585
R7174 GND.n2519 GND.n1825 585
R7175 GND.n4448 GND.n1825 585
R7176 GND.n3560 GND.n3558 585
R7177 GND.n3558 GND.n3557 585
R7178 GND.n3561 GND.n1816 585
R7179 GND.n4454 GND.n1816 585
R7180 GND.n3562 GND.n2528 585
R7181 GND.n3582 GND.n2528 585
R7182 GND.n2533 GND.n1807 585
R7183 GND.n4462 GND.n1807 585
R7184 GND.n3567 GND.n3566 585
R7185 GND.n3568 GND.n3567 585
R7186 GND.n2532 GND.n1797 585
R7187 GND.n4468 GND.n1797 585
R7188 GND.n3551 GND.n3550 585
R7189 GND.n3550 GND.n3549 585
R7190 GND.n2535 GND.n1787 585
R7191 GND.n4476 GND.n1787 585
R7192 GND.n3507 GND.n2539 585
R7193 GND.n3537 GND.n2539 585
R7194 GND.n3508 GND.n1777 585
R7195 GND.n4482 GND.n1777 585
R7196 GND.n3509 GND.n3505 585
R7197 GND.n3505 GND.n3504 585
R7198 GND.n2565 GND.n1767 585
R7199 GND.n4490 GND.n1767 585
R7200 GND.n3514 GND.n3513 585
R7201 GND.n3515 GND.n3514 585
R7202 GND.n2564 GND.n1757 585
R7203 GND.n4496 GND.n1757 585
R7204 GND.n3487 GND.n3486 585
R7205 GND.n3488 GND.n3487 585
R7206 GND.n2570 GND.n1747 585
R7207 GND.n4504 GND.n1747 585
R7208 GND.n3482 GND.n3481 585
R7209 GND.n3481 GND.n3480 585
R7210 GND.n3295 GND.n1735 585
R7211 GND.n4510 GND.n1735 585
R7212 GND.n3294 GND.n2576 585
R7213 GND.n2576 GND.n2575 585
R7214 GND.n2573 GND.n2572 585
R7215 GND.n2573 GND.n1723 585
R7216 GND.n3290 GND.n1722 585
R7217 GND.n4518 GND.n1722 585
R7218 GND.n3289 GND.n3288 585
R7219 GND.n3288 GND.n3287 585
R7220 GND.n3286 GND.n1709 585
R7221 GND.n4524 GND.n1709 585
R7222 GND.n3280 GND.n2578 585
R7223 GND.n3280 GND.n1708 585
R7224 GND.n3282 GND.n3281 585
R7225 GND.n3281 GND.n1696 585
R7226 GND.n3279 GND.n1695 585
R7227 GND.n4532 GND.n1695 585
R7228 GND.n3278 GND.n2582 585
R7229 GND.n2582 GND.n2581 585
R7230 GND.n2580 GND.n1681 585
R7231 GND.n4538 GND.n1681 585
R7232 GND.n3274 GND.n3273 585
R7233 GND.n3273 GND.n3272 585
R7234 GND.n3270 GND.n3269 585
R7235 GND.n3270 GND.n1670 585
R7236 GND.n3268 GND.n1669 585
R7237 GND.n4546 GND.n1669 585
R7238 GND.n3227 GND.n1528 585
R7239 GND.n4685 GND.n1528 585
R7240 GND.n3229 GND.n3228 585
R7241 GND.n3230 GND.n3229 585
R7242 GND.n3226 GND.n1519 585
R7243 GND.n3226 GND.n3225 585
R7244 GND.n2593 GND.n1518 585
R7245 GND.n3206 GND.n2593 585
R7246 GND.n3216 GND.n1517 585
R7247 GND.n3217 GND.n3216 585
R7248 GND.n3215 GND.n2603 585
R7249 GND.n3215 GND.n3214 585
R7250 GND.n2602 GND.n1511 585
R7251 GND.n3185 GND.n2602 585
R7252 GND.n3175 GND.n1510 585
R7253 GND.n3175 GND.n2619 585
R7254 GND.n3176 GND.n1509 585
R7255 GND.n3177 GND.n3176 585
R7256 GND.n3174 GND.n2629 585
R7257 GND.n3174 GND.n3173 585
R7258 GND.n2628 GND.n1503 585
R7259 GND.n3040 GND.n2628 585
R7260 GND.n2639 GND.n1502 585
R7261 GND.n3161 GND.n2639 585
R7262 GND.n3148 GND.n1501 585
R7263 GND.n3148 GND.n3147 585
R7264 GND.n3150 GND.n3149 585
R7265 GND.n3151 GND.n3150 585
R7266 GND.n3146 GND.n1495 585
R7267 GND.n3146 GND.n3145 585
R7268 GND.n2649 GND.n1494 585
R7269 GND.n3061 GND.n2649 585
R7270 GND.n2658 GND.n1493 585
R7271 GND.n3136 GND.n2658 585
R7272 GND.n3124 GND.n3122 585
R7273 GND.n3124 GND.n3123 585
R7274 GND.n3125 GND.n1487 585
R7275 GND.n3126 GND.n3125 585
R7276 GND.n3121 GND.n1486 585
R7277 GND.n3121 GND.n3120 585
R7278 GND.n2668 GND.n1485 585
R7279 GND.n3070 GND.n2668 585
R7280 GND.n2679 GND.n2678 585
R7281 GND.n3111 GND.n2679 585
R7282 GND.n2721 GND.n1479 585
R7283 GND.n3021 GND.n2721 585
R7284 GND.n3081 GND.n1478 585
R7285 GND.n3081 GND.n3080 585
R7286 GND.n3082 GND.n1477 585
R7287 GND.n3083 GND.n3082 585
R7288 GND.n2711 GND.n2710 585
R7289 GND.n3088 GND.n2711 585
R7290 GND.n2709 GND.n1471 585
R7291 GND.n2709 GND.n2706 585
R7292 GND.n2696 GND.n1470 585
R7293 GND.n2699 GND.n2696 585
R7294 GND.n3098 GND.n1469 585
R7295 GND.n3098 GND.n3097 585
R7296 GND.n3100 GND.n3099 585
R7297 GND.n3101 GND.n3100 585
R7298 GND.n2695 GND.n1463 585
R7299 GND.n3004 GND.n2695 585
R7300 GND.n2963 GND.n1462 585
R7301 GND.n2963 GND.n2730 585
R7302 GND.n2964 GND.n1461 585
R7303 GND.n2965 GND.n2964 585
R7304 GND.n2741 GND.n2740 585
R7305 GND.n2990 GND.n2741 585
R7306 GND.n2979 GND.n1455 585
R7307 GND.n2979 GND.n2738 585
R7308 GND.n2980 GND.n1454 585
R7309 GND.n2981 GND.n2980 585
R7310 GND.n2978 GND.n1453 585
R7311 GND.n2978 GND.n2977 585
R7312 GND.n2754 GND.n2753 585
R7313 GND.n2766 GND.n2754 585
R7314 GND.n2764 GND.n1447 585
R7315 GND.n2954 GND.n2764 585
R7316 GND.n2942 GND.n1446 585
R7317 GND.n2942 GND.n2941 585
R7318 GND.n2943 GND.n1445 585
R7319 GND.n2944 GND.n2943 585
R7320 GND.n2939 GND.n2938 585
R7321 GND.n2939 GND.n2772 585
R7322 GND.n2937 GND.n1439 585
R7323 GND.n2937 GND.n2936 585
R7324 GND.n2791 GND.n1438 585
R7325 GND.n2801 GND.n2791 585
R7326 GND.n2927 GND.n1437 585
R7327 GND.n2928 GND.n2927 585
R7328 GND.n2926 GND.n2925 585
R7329 GND.n2926 GND.n2798 585
R7330 GND.n2924 GND.n1431 585
R7331 GND.n2924 GND.n2923 585
R7332 GND.n2802 GND.n1430 585
R7333 GND.n2804 GND.n2802 585
R7334 GND.n2914 GND.n1429 585
R7335 GND.n2915 GND.n2914 585
R7336 GND.n2913 GND.n2912 585
R7337 GND.n2913 GND.n2811 585
R7338 GND.n2911 GND.n1423 585
R7339 GND.n2911 GND.n2910 585
R7340 GND.n2813 GND.n1422 585
R7341 GND.n2814 GND.n2813 585
R7342 GND.n2838 GND.n1421 585
R7343 GND.n2838 GND.n1375 585
R7344 GND.n2840 GND.n2839 585
R7345 GND.n2836 GND.n2835 585
R7346 GND.n2844 GND.n2837 585
R7347 GND.n2846 GND.n2845 585
R7348 GND.n2848 GND.n2847 585
R7349 GND.n2832 GND.n2831 585
R7350 GND.n2852 GND.n2833 585
R7351 GND.n2854 GND.n2853 585
R7352 GND.n2856 GND.n2855 585
R7353 GND.n2828 GND.n2827 585
R7354 GND.n2860 GND.n2829 585
R7355 GND.n2862 GND.n2861 585
R7356 GND.n2864 GND.n2863 585
R7357 GND.n2824 GND.n2823 585
R7358 GND.n2868 GND.n2825 585
R7359 GND.n2869 GND.n2820 585
R7360 GND.n2870 GND.n1374 585
R7361 GND.n4837 GND.n1374 585
R7362 GND.n4586 GND.n4585 585
R7363 GND.n1626 GND.n1620 585
R7364 GND.n4593 GND.n1617 585
R7365 GND.n4594 GND.n1616 585
R7366 GND.n1636 GND.n1610 585
R7367 GND.n4601 GND.n1609 585
R7368 GND.n4602 GND.n1608 585
R7369 GND.n1634 GND.n1602 585
R7370 GND.n4609 GND.n1601 585
R7371 GND.n4610 GND.n1600 585
R7372 GND.n1631 GND.n1594 585
R7373 GND.n4617 GND.n1593 585
R7374 GND.n4618 GND.n1592 585
R7375 GND.n1629 GND.n1584 585
R7376 GND.n4625 GND.n1583 585
R7377 GND.n4626 GND.n1582 585
R7378 GND.n4627 GND.n1581 585
R7379 GND.n4583 GND.n1581 585
R7380 GND.n3233 GND.n1526 585
R7381 GND.n4685 GND.n1526 585
R7382 GND.n3232 GND.n3231 585
R7383 GND.n3231 GND.n3230 585
R7384 GND.n2591 GND.n2590 585
R7385 GND.n3225 GND.n2591 585
R7386 GND.n3208 GND.n3207 585
R7387 GND.n3207 GND.n3206 585
R7388 GND.n2607 GND.n2600 585
R7389 GND.n3217 GND.n2600 585
R7390 GND.n3213 GND.n3212 585
R7391 GND.n3214 GND.n3213 585
R7392 GND.n2606 GND.n2605 585
R7393 GND.n3185 GND.n2605 585
R7394 GND.n3167 GND.n3166 585
R7395 GND.n3166 GND.n2619 585
R7396 GND.n2632 GND.n2626 585
R7397 GND.n3177 GND.n2626 585
R7398 GND.n3172 GND.n3171 585
R7399 GND.n3173 GND.n3172 585
R7400 GND.n2631 GND.n2630 585
R7401 GND.n3040 GND.n2630 585
R7402 GND.n3163 GND.n3162 585
R7403 GND.n3162 GND.n3161 585
R7404 GND.n2635 GND.n2634 585
R7405 GND.n3147 GND.n2635 585
R7406 GND.n2652 GND.n2647 585
R7407 GND.n3151 GND.n2647 585
R7408 GND.n3144 GND.n3143 585
R7409 GND.n3145 GND.n3144 585
R7410 GND.n2651 GND.n2650 585
R7411 GND.n3061 GND.n2650 585
R7412 GND.n3138 GND.n3137 585
R7413 GND.n3137 GND.n3136 585
R7414 GND.n2655 GND.n2654 585
R7415 GND.n3123 GND.n2655 585
R7416 GND.n2672 GND.n2666 585
R7417 GND.n3126 GND.n2666 585
R7418 GND.n3119 GND.n3118 585
R7419 GND.n3120 GND.n3119 585
R7420 GND.n2671 GND.n2670 585
R7421 GND.n3070 GND.n2670 585
R7422 GND.n3113 GND.n3112 585
R7423 GND.n3112 GND.n3111 585
R7424 GND.n2675 GND.n2674 585
R7425 GND.n3021 GND.n2675 585
R7426 GND.n3020 GND.n3019 585
R7427 GND.n3080 GND.n3020 585
R7428 GND.n2723 GND.n2719 585
R7429 GND.n3083 GND.n2719 585
R7430 GND.n3015 GND.n2707 585
R7431 GND.n3088 GND.n2707 585
R7432 GND.n3014 GND.n3013 585
R7433 GND.n3013 GND.n2706 585
R7434 GND.n3012 GND.n3011 585
R7435 GND.n3012 GND.n2699 585
R7436 GND.n2725 GND.n2697 585
R7437 GND.n3097 GND.n2697 585
R7438 GND.n3007 GND.n2693 585
R7439 GND.n3101 GND.n2693 585
R7440 GND.n3006 GND.n3005 585
R7441 GND.n3005 GND.n3004 585
R7442 GND.n2728 GND.n2727 585
R7443 GND.n2730 GND.n2728 585
R7444 GND.n2969 GND.n2966 585
R7445 GND.n2966 GND.n2965 585
R7446 GND.n2970 GND.n2739 585
R7447 GND.n2990 GND.n2739 585
R7448 GND.n2971 GND.n2960 585
R7449 GND.n2960 GND.n2738 585
R7450 GND.n2758 GND.n2751 585
R7451 GND.n2981 GND.n2751 585
R7452 GND.n2976 GND.n2975 585
R7453 GND.n2977 GND.n2976 585
R7454 GND.n2757 GND.n2756 585
R7455 GND.n2766 GND.n2756 585
R7456 GND.n2956 GND.n2955 585
R7457 GND.n2955 GND.n2954 585
R7458 GND.n2761 GND.n2760 585
R7459 GND.n2941 GND.n2761 585
R7460 GND.n2884 GND.n2773 585
R7461 GND.n2944 GND.n2773 585
R7462 GND.n2883 GND.n2882 585
R7463 GND.n2882 GND.n2772 585
R7464 GND.n2888 GND.n2792 585
R7465 GND.n2936 GND.n2792 585
R7466 GND.n2889 GND.n2881 585
R7467 GND.n2881 GND.n2801 585
R7468 GND.n2890 GND.n2799 585
R7469 GND.n2928 GND.n2799 585
R7470 GND.n2879 GND.n2878 585
R7471 GND.n2878 GND.n2798 585
R7472 GND.n2894 GND.n2805 585
R7473 GND.n2923 GND.n2805 585
R7474 GND.n2895 GND.n2877 585
R7475 GND.n2877 GND.n2804 585
R7476 GND.n2896 GND.n2812 585
R7477 GND.n2915 GND.n2812 585
R7478 GND.n2818 GND.n2816 585
R7479 GND.n2816 GND.n2811 585
R7480 GND.n2901 GND.n2900 585
R7481 GND.n2910 GND.n2901 585
R7482 GND.n2817 GND.n2815 585
R7483 GND.n2815 GND.n2814 585
R7484 GND.n2873 GND.n2872 585
R7485 GND.n2872 GND.n1375 585
R7486 GND.n4684 GND.n4683 585
R7487 GND.n4685 GND.n4684 585
R7488 GND.n1531 GND.n1529 585
R7489 GND.n3230 GND.n1529 585
R7490 GND.n3224 GND.n3223 585
R7491 GND.n3225 GND.n3224 585
R7492 GND.n2595 GND.n2594 585
R7493 GND.n3206 GND.n2594 585
R7494 GND.n3219 GND.n3218 585
R7495 GND.n3218 GND.n3217 585
R7496 GND.n2598 GND.n2597 585
R7497 GND.n3214 GND.n2598 585
R7498 GND.n3184 GND.n3183 585
R7499 GND.n3185 GND.n3184 585
R7500 GND.n2621 GND.n2620 585
R7501 GND.n2620 GND.n2619 585
R7502 GND.n3179 GND.n3178 585
R7503 GND.n3178 GND.n3177 585
R7504 GND.n2624 GND.n2623 585
R7505 GND.n3173 GND.n2624 585
R7506 GND.n3158 GND.n2641 585
R7507 GND.n3040 GND.n2641 585
R7508 GND.n3160 GND.n3159 585
R7509 GND.n3161 GND.n3160 585
R7510 GND.n2642 GND.n2640 585
R7511 GND.n3147 GND.n2640 585
R7512 GND.n3153 GND.n3152 585
R7513 GND.n3152 GND.n3151 585
R7514 GND.n2645 GND.n2644 585
R7515 GND.n3145 GND.n2645 585
R7516 GND.n3133 GND.n2660 585
R7517 GND.n3061 GND.n2660 585
R7518 GND.n3135 GND.n3134 585
R7519 GND.n3136 GND.n3135 585
R7520 GND.n2661 GND.n2659 585
R7521 GND.n3123 GND.n2659 585
R7522 GND.n3128 GND.n3127 585
R7523 GND.n3127 GND.n3126 585
R7524 GND.n2664 GND.n2663 585
R7525 GND.n3120 GND.n2664 585
R7526 GND.n3108 GND.n2681 585
R7527 GND.n3070 GND.n2681 585
R7528 GND.n3110 GND.n3109 585
R7529 GND.n3111 GND.n3110 585
R7530 GND.n2682 GND.n2680 585
R7531 GND.n3021 GND.n2680 585
R7532 GND.n2717 GND.n2716 585
R7533 GND.n3080 GND.n2716 585
R7534 GND.n3084 GND.n2718 585
R7535 GND.n3084 GND.n3083 585
R7536 GND.n3087 GND.n3086 585
R7537 GND.n3088 GND.n3087 585
R7538 GND.n3085 GND.n2715 585
R7539 GND.n2715 GND.n2706 585
R7540 GND.n2714 GND.n2713 585
R7541 GND.n2714 GND.n2699 585
R7542 GND.n2712 GND.n2691 585
R7543 GND.n3097 GND.n2691 585
R7544 GND.n3103 GND.n3102 585
R7545 GND.n3102 GND.n3101 585
R7546 GND.n3104 GND.n2690 585
R7547 GND.n3004 GND.n2690 585
R7548 GND.n2743 GND.n2689 585
R7549 GND.n2743 GND.n2730 585
R7550 GND.n2987 GND.n2744 585
R7551 GND.n2965 GND.n2744 585
R7552 GND.n2989 GND.n2988 585
R7553 GND.n2990 GND.n2989 585
R7554 GND.n2745 GND.n2742 585
R7555 GND.n2742 GND.n2738 585
R7556 GND.n2983 GND.n2982 585
R7557 GND.n2982 GND.n2981 585
R7558 GND.n2748 GND.n2747 585
R7559 GND.n2977 GND.n2748 585
R7560 GND.n2951 GND.n2767 585
R7561 GND.n2767 GND.n2766 585
R7562 GND.n2953 GND.n2952 585
R7563 GND.n2954 GND.n2953 585
R7564 GND.n2768 GND.n2765 585
R7565 GND.n2941 GND.n2765 585
R7566 GND.n2946 GND.n2945 585
R7567 GND.n2945 GND.n2944 585
R7568 GND.n2771 GND.n2770 585
R7569 GND.n2772 GND.n2771 585
R7570 GND.n2935 GND.n2934 585
R7571 GND.n2936 GND.n2935 585
R7572 GND.n2794 GND.n2793 585
R7573 GND.n2801 GND.n2793 585
R7574 GND.n2930 GND.n2929 585
R7575 GND.n2929 GND.n2928 585
R7576 GND.n2797 GND.n2796 585
R7577 GND.n2798 GND.n2797 585
R7578 GND.n2922 GND.n2921 585
R7579 GND.n2923 GND.n2922 585
R7580 GND.n2807 GND.n2806 585
R7581 GND.n2806 GND.n2804 585
R7582 GND.n2917 GND.n2916 585
R7583 GND.n2916 GND.n2915 585
R7584 GND.n2810 GND.n2809 585
R7585 GND.n2811 GND.n2810 585
R7586 GND.n2909 GND.n2908 585
R7587 GND.n2910 GND.n2909 585
R7588 GND.n2903 GND.n2902 585
R7589 GND.n2902 GND.n2814 585
R7590 GND.n2904 GND.n1378 585
R7591 GND.n1378 GND.n1375 585
R7592 GND.n4835 GND.n4834 585
R7593 GND.n4833 GND.n1377 585
R7594 GND.n4832 GND.n1376 585
R7595 GND.n4837 GND.n1376 585
R7596 GND.n4831 GND.n4830 585
R7597 GND.n4829 GND.n4828 585
R7598 GND.n4827 GND.n4826 585
R7599 GND.n4825 GND.n4824 585
R7600 GND.n4823 GND.n4822 585
R7601 GND.n4821 GND.n4820 585
R7602 GND.n4819 GND.n4818 585
R7603 GND.n4817 GND.n4816 585
R7604 GND.n4815 GND.n4814 585
R7605 GND.n4813 GND.n4812 585
R7606 GND.n4811 GND.n4810 585
R7607 GND.n4809 GND.n4808 585
R7608 GND.n4807 GND.n4806 585
R7609 GND.n4804 GND.n4803 585
R7610 GND.n4802 GND.n4801 585
R7611 GND.n4800 GND.n4799 585
R7612 GND.n4798 GND.n4797 585
R7613 GND.n4796 GND.n4795 585
R7614 GND.n4794 GND.n4793 585
R7615 GND.n4792 GND.n4791 585
R7616 GND.n4790 GND.n4789 585
R7617 GND.n4788 GND.n4787 585
R7618 GND.n4786 GND.n4785 585
R7619 GND.n4784 GND.n4783 585
R7620 GND.n4782 GND.n4781 585
R7621 GND.n4780 GND.n4779 585
R7622 GND.n4778 GND.n4777 585
R7623 GND.n4776 GND.n4775 585
R7624 GND.n4774 GND.n4773 585
R7625 GND.n4772 GND.n1413 585
R7626 GND.n1417 GND.n1414 585
R7627 GND.n4768 GND.n4767 585
R7628 GND.n4631 GND.n1524 585
R7629 GND.n4558 GND.n1578 585
R7630 GND.n4635 GND.n1575 585
R7631 GND.n4636 GND.n1574 585
R7632 GND.n4637 GND.n1573 585
R7633 GND.n4561 GND.n1571 585
R7634 GND.n4641 GND.n1570 585
R7635 GND.n4642 GND.n1569 585
R7636 GND.n4643 GND.n1568 585
R7637 GND.n4564 GND.n1566 585
R7638 GND.n4647 GND.n1565 585
R7639 GND.n4648 GND.n1564 585
R7640 GND.n4649 GND.n1563 585
R7641 GND.n4567 GND.n1561 585
R7642 GND.n4653 GND.n1560 585
R7643 GND.n4654 GND.n1559 585
R7644 GND.n4655 GND.n1558 585
R7645 GND.n4570 GND.n1556 585
R7646 GND.n4659 GND.n1555 585
R7647 GND.n4661 GND.n1549 585
R7648 GND.n4662 GND.n1548 585
R7649 GND.n4574 GND.n1546 585
R7650 GND.n4666 GND.n1545 585
R7651 GND.n4667 GND.n1544 585
R7652 GND.n4668 GND.n1543 585
R7653 GND.n4577 GND.n1541 585
R7654 GND.n4672 GND.n1540 585
R7655 GND.n4673 GND.n1539 585
R7656 GND.n4674 GND.n1538 585
R7657 GND.n4580 GND.n1536 585
R7658 GND.n4678 GND.n1535 585
R7659 GND.n4679 GND.n1534 585
R7660 GND.n4680 GND.n1530 585
R7661 GND.n4583 GND.n1530 585
R7662 GND.n4687 GND.n4686 585
R7663 GND.n4686 GND.n4685 585
R7664 GND.n4688 GND.n1522 585
R7665 GND.n3230 GND.n1522 585
R7666 GND.n4689 GND.n1521 585
R7667 GND.n3225 GND.n1521 585
R7668 GND.n2610 GND.n1516 585
R7669 GND.n3206 GND.n2610 585
R7670 GND.n4693 GND.n1515 585
R7671 GND.n3217 GND.n1515 585
R7672 GND.n4694 GND.n1514 585
R7673 GND.n3214 GND.n1514 585
R7674 GND.n4695 GND.n1513 585
R7675 GND.n3185 GND.n1513 585
R7676 GND.n2618 GND.n1508 585
R7677 GND.n2619 GND.n2618 585
R7678 GND.n4699 GND.n1507 585
R7679 GND.n3177 GND.n1507 585
R7680 GND.n4700 GND.n1506 585
R7681 GND.n3173 GND.n1506 585
R7682 GND.n4701 GND.n1505 585
R7683 GND.n3040 GND.n1505 585
R7684 GND.n2637 GND.n1500 585
R7685 GND.n3161 GND.n2637 585
R7686 GND.n4705 GND.n1499 585
R7687 GND.n3147 GND.n1499 585
R7688 GND.n4706 GND.n1498 585
R7689 GND.n3151 GND.n1498 585
R7690 GND.n4707 GND.n1497 585
R7691 GND.n3145 GND.n1497 585
R7692 GND.n3060 GND.n1492 585
R7693 GND.n3061 GND.n3060 585
R7694 GND.n4711 GND.n1491 585
R7695 GND.n3136 GND.n1491 585
R7696 GND.n4712 GND.n1490 585
R7697 GND.n3123 GND.n1490 585
R7698 GND.n4713 GND.n1489 585
R7699 GND.n3126 GND.n1489 585
R7700 GND.n2669 GND.n1484 585
R7701 GND.n3120 GND.n2669 585
R7702 GND.n4717 GND.n1483 585
R7703 GND.n3070 GND.n1483 585
R7704 GND.n4718 GND.n1482 585
R7705 GND.n3111 GND.n1482 585
R7706 GND.n4719 GND.n1481 585
R7707 GND.n3021 GND.n1481 585
R7708 GND.n2722 GND.n1476 585
R7709 GND.n3080 GND.n2722 585
R7710 GND.n4723 GND.n1475 585
R7711 GND.n3083 GND.n1475 585
R7712 GND.n4724 GND.n1474 585
R7713 GND.n3088 GND.n1474 585
R7714 GND.n4725 GND.n1473 585
R7715 GND.n2706 GND.n1473 585
R7716 GND.n2698 GND.n1468 585
R7717 GND.n2699 GND.n2698 585
R7718 GND.n4729 GND.n1467 585
R7719 GND.n3097 GND.n1467 585
R7720 GND.n4730 GND.n1466 585
R7721 GND.n3101 GND.n1466 585
R7722 GND.n4731 GND.n1465 585
R7723 GND.n3004 GND.n1465 585
R7724 GND.n2729 GND.n1460 585
R7725 GND.n2730 GND.n2729 585
R7726 GND.n4735 GND.n1459 585
R7727 GND.n2965 GND.n1459 585
R7728 GND.n4736 GND.n1458 585
R7729 GND.n2990 GND.n1458 585
R7730 GND.n4737 GND.n1457 585
R7731 GND.n2738 GND.n1457 585
R7732 GND.n2750 GND.n1452 585
R7733 GND.n2981 GND.n2750 585
R7734 GND.n4741 GND.n1451 585
R7735 GND.n2977 GND.n1451 585
R7736 GND.n4742 GND.n1450 585
R7737 GND.n2766 GND.n1450 585
R7738 GND.n4743 GND.n1449 585
R7739 GND.n2954 GND.n1449 585
R7740 GND.n2940 GND.n1444 585
R7741 GND.n2941 GND.n2940 585
R7742 GND.n4747 GND.n1443 585
R7743 GND.n2944 GND.n1443 585
R7744 GND.n4748 GND.n1442 585
R7745 GND.n2772 GND.n1442 585
R7746 GND.n4749 GND.n1441 585
R7747 GND.n2936 GND.n1441 585
R7748 GND.n2800 GND.n1436 585
R7749 GND.n2801 GND.n2800 585
R7750 GND.n4753 GND.n1435 585
R7751 GND.n2928 GND.n1435 585
R7752 GND.n4754 GND.n1434 585
R7753 GND.n2798 GND.n1434 585
R7754 GND.n4755 GND.n1433 585
R7755 GND.n2923 GND.n1433 585
R7756 GND.n2803 GND.n1428 585
R7757 GND.n2804 GND.n2803 585
R7758 GND.n4759 GND.n1427 585
R7759 GND.n2915 GND.n1427 585
R7760 GND.n4760 GND.n1426 585
R7761 GND.n2811 GND.n1426 585
R7762 GND.n4761 GND.n1425 585
R7763 GND.n2910 GND.n1425 585
R7764 GND.n1420 GND.n1419 585
R7765 GND.n2814 GND.n1419 585
R7766 GND.n4766 GND.n4765 585
R7767 GND.n4766 GND.n1375 585
R7768 GND.n5602 GND.n742 585
R7769 GND.n742 GND.n715 585
R7770 GND.n5604 GND.n5603 585
R7771 GND.n5605 GND.n5604 585
R7772 GND.n806 GND.n805 585
R7773 GND.n805 GND.n804 585
R7774 GND.n5598 GND.n5597 585
R7775 GND.n5597 GND.n5596 585
R7776 GND.n809 GND.n808 585
R7777 GND.n810 GND.n809 585
R7778 GND.n5585 GND.n5584 585
R7779 GND.n5586 GND.n5585 585
R7780 GND.n823 GND.n822 585
R7781 GND.n822 GND.n820 585
R7782 GND.n5580 GND.n5579 585
R7783 GND.n5579 GND.n5578 585
R7784 GND.n826 GND.n825 585
R7785 GND.n827 GND.n826 585
R7786 GND.n5568 GND.n5567 585
R7787 GND.n5569 GND.n5568 585
R7788 GND.n842 GND.n841 585
R7789 GND.n849 GND.n841 585
R7790 GND.n5563 GND.n5562 585
R7791 GND.n5562 GND.n5561 585
R7792 GND.n845 GND.n844 585
R7793 GND.n846 GND.n845 585
R7794 GND.n5551 GND.n5550 585
R7795 GND.n5552 GND.n5551 585
R7796 GND.n864 GND.n863 585
R7797 GND.n5528 GND.n863 585
R7798 GND.n5546 GND.n5545 585
R7799 GND.n5545 GND.n5544 585
R7800 GND.n867 GND.n866 585
R7801 GND.n5536 GND.n867 585
R7802 GND.n4172 GND.n2242 585
R7803 GND.n2242 GND.n881 585
R7804 GND.n4174 GND.n4173 585
R7805 GND.n4175 GND.n4174 585
R7806 GND.n2243 GND.n2241 585
R7807 GND.n2249 GND.n2241 585
R7808 GND.n4167 GND.n4166 585
R7809 GND.n4166 GND.n4165 585
R7810 GND.n2246 GND.n2245 585
R7811 GND.n4162 GND.n2246 585
R7812 GND.n4100 GND.n4099 585
R7813 GND.n4100 GND.n2252 585
R7814 GND.n4101 GND.n4097 585
R7815 GND.n4116 GND.n4101 585
R7816 GND.n4121 GND.n4120 585
R7817 GND.n4120 GND.n4119 585
R7818 GND.n4123 GND.n4093 585
R7819 GND.n4104 GND.n4093 585
R7820 GND.n4125 GND.n4124 585
R7821 GND.n4126 GND.n4125 585
R7822 GND.n4095 GND.n4092 585
R7823 GND.n4092 GND.n4084 585
R7824 GND.n4094 GND.n2274 585
R7825 GND.n4133 GND.n2274 585
R7826 GND.n4138 GND.n4137 585
R7827 GND.n4137 GND.n4136 585
R7828 GND.n4139 GND.n2271 585
R7829 GND.n4075 GND.n2271 585
R7830 GND.n4142 GND.n4141 585
R7831 GND.n4143 GND.n4142 585
R7832 GND.n2272 GND.n2270 585
R7833 GND.n2270 GND.n2265 585
R7834 GND.n4064 GND.n2299 585
R7835 GND.n2299 GND.n2298 585
R7836 GND.n4066 GND.n4065 585
R7837 GND.n4067 GND.n4066 585
R7838 GND.n2300 GND.n2293 585
R7839 GND.n4053 GND.n2293 585
R7840 GND.n4058 GND.n4057 585
R7841 GND.n4057 GND.n4056 585
R7842 GND.n2303 GND.n2302 585
R7843 GND.n4050 GND.n2303 585
R7844 GND.n4038 GND.n2322 585
R7845 GND.n2322 GND.n2321 585
R7846 GND.n4040 GND.n4039 585
R7847 GND.n4041 GND.n4040 585
R7848 GND.n2323 GND.n2320 585
R7849 GND.n4028 GND.n2320 585
R7850 GND.n4033 GND.n4032 585
R7851 GND.n4032 GND.n4031 585
R7852 GND.n2326 GND.n2325 585
R7853 GND.n4026 GND.n2326 585
R7854 GND.n4014 GND.n2345 585
R7855 GND.n2345 GND.n2344 585
R7856 GND.n4016 GND.n4015 585
R7857 GND.n4017 GND.n4016 585
R7858 GND.n2346 GND.n2343 585
R7859 GND.n4004 GND.n2343 585
R7860 GND.n4009 GND.n4008 585
R7861 GND.n4008 GND.n4007 585
R7862 GND.n2349 GND.n2348 585
R7863 GND.n4001 GND.n2349 585
R7864 GND.n3989 GND.n2368 585
R7865 GND.n2368 GND.n2367 585
R7866 GND.n3991 GND.n3990 585
R7867 GND.n3992 GND.n3991 585
R7868 GND.n2369 GND.n2366 585
R7869 GND.n3978 GND.n2366 585
R7870 GND.n3984 GND.n3983 585
R7871 GND.n3983 GND.n3982 585
R7872 GND.n2412 GND.n2371 585
R7873 GND.n3918 GND.n2412 585
R7874 GND.n2411 GND.n2410 585
R7875 GND.n2409 GND.n2408 585
R7876 GND.n2407 GND.n2406 585
R7877 GND.n2405 GND.n2404 585
R7878 GND.n2403 GND.n2402 585
R7879 GND.n2401 GND.n2400 585
R7880 GND.n2399 GND.n2398 585
R7881 GND.n2397 GND.n2396 585
R7882 GND.n2395 GND.n2394 585
R7883 GND.n2393 GND.n2392 585
R7884 GND.n2391 GND.n2390 585
R7885 GND.n2389 GND.n2388 585
R7886 GND.n2387 GND.n2386 585
R7887 GND.n2019 GND.n2003 585
R7888 GND.n4308 GND.n2020 585
R7889 GND.n4311 GND.n4310 585
R7890 GND.n2010 GND.n2009 585
R7891 GND.n2131 GND.n2130 585
R7892 GND.n2129 GND.n2127 585
R7893 GND.n2136 GND.n2135 585
R7894 GND.n2138 GND.n2137 585
R7895 GND.n2141 GND.n2140 585
R7896 GND.n2139 GND.n2125 585
R7897 GND.n2146 GND.n2145 585
R7898 GND.n2148 GND.n2147 585
R7899 GND.n2151 GND.n2150 585
R7900 GND.n2149 GND.n2123 585
R7901 GND.n2156 GND.n2155 585
R7902 GND.n2158 GND.n2157 585
R7903 GND.n2161 GND.n2160 585
R7904 GND.n2159 GND.n2120 585
R7905 GND.n2165 GND.n2121 585
R7906 GND.n2166 GND.n2116 585
R7907 GND.n2168 GND.n2167 585
R7908 GND.n5658 GND.n5657 585
R7909 GND.n797 GND.n796 585
R7910 GND.n5662 GND.n793 585
R7911 GND.n5663 GND.n792 585
R7912 GND.n5664 GND.n791 585
R7913 GND.n789 GND.n788 585
R7914 GND.n5668 GND.n787 585
R7915 GND.n5669 GND.n786 585
R7916 GND.n5670 GND.n785 585
R7917 GND.n783 GND.n782 585
R7918 GND.n5674 GND.n781 585
R7919 GND.n5675 GND.n780 585
R7920 GND.n5676 GND.n779 585
R7921 GND.n777 GND.n776 585
R7922 GND.n5680 GND.n775 585
R7923 GND.n5681 GND.n774 585
R7924 GND.n5682 GND.n773 585
R7925 GND.n771 GND.n770 585
R7926 GND.n5686 GND.n769 585
R7927 GND.n5688 GND.n766 585
R7928 GND.n5689 GND.n765 585
R7929 GND.n763 GND.n762 585
R7930 GND.n5693 GND.n761 585
R7931 GND.n5694 GND.n760 585
R7932 GND.n5695 GND.n759 585
R7933 GND.n757 GND.n756 585
R7934 GND.n5699 GND.n755 585
R7935 GND.n5700 GND.n754 585
R7936 GND.n5701 GND.n753 585
R7937 GND.n751 GND.n750 585
R7938 GND.n5705 GND.n749 585
R7939 GND.n5706 GND.n748 585
R7940 GND.n5707 GND.n747 585
R7941 GND.n744 GND.n743 585
R7942 GND.n5712 GND.n5711 585
R7943 GND.n5713 GND.n5712 585
R7944 GND.n5656 GND.n5655 585
R7945 GND.n5656 GND.n715 585
R7946 GND.n800 GND.n799 585
R7947 GND.n5605 GND.n799 585
R7948 GND.n5591 GND.n5590 585
R7949 GND.n5590 GND.n804 585
R7950 GND.n5592 GND.n811 585
R7951 GND.n5596 GND.n811 585
R7952 GND.n5589 GND.n5588 585
R7953 GND.n5588 GND.n810 585
R7954 GND.n5587 GND.n818 585
R7955 GND.n5587 GND.n5586 585
R7956 GND.n5573 GND.n819 585
R7957 GND.n820 GND.n819 585
R7958 GND.n5574 GND.n828 585
R7959 GND.n5578 GND.n828 585
R7960 GND.n5572 GND.n5571 585
R7961 GND.n5571 GND.n827 585
R7962 GND.n5570 GND.n838 585
R7963 GND.n5570 GND.n5569 585
R7964 GND.n5556 GND.n839 585
R7965 GND.n849 GND.n839 585
R7966 GND.n5557 GND.n847 585
R7967 GND.n5561 GND.n847 585
R7968 GND.n5555 GND.n5554 585
R7969 GND.n5554 GND.n846 585
R7970 GND.n5553 GND.n858 585
R7971 GND.n5553 GND.n5552 585
R7972 GND.n5539 GND.n859 585
R7973 GND.n5528 GND.n859 585
R7974 GND.n5540 GND.n869 585
R7975 GND.n5544 GND.n869 585
R7976 GND.n5538 GND.n5537 585
R7977 GND.n5537 GND.n5536 585
R7978 GND.n880 GND.n879 585
R7979 GND.n881 GND.n880 585
R7980 GND.n4181 GND.n2235 585
R7981 GND.n4175 GND.n2235 585
R7982 GND.n4182 GND.n2234 585
R7983 GND.n2249 GND.n2234 585
R7984 GND.n4183 GND.n2233 585
R7985 GND.n4165 GND.n2233 585
R7986 GND.n4161 GND.n2228 585
R7987 GND.n4162 GND.n4161 585
R7988 GND.n4187 GND.n2227 585
R7989 GND.n2252 GND.n2227 585
R7990 GND.n4188 GND.n2226 585
R7991 GND.n4116 GND.n2226 585
R7992 GND.n4189 GND.n2225 585
R7993 GND.n4119 GND.n2225 585
R7994 GND.n4103 GND.n2220 585
R7995 GND.n4104 GND.n4103 585
R7996 GND.n4193 GND.n2219 585
R7997 GND.n4126 GND.n2219 585
R7998 GND.n4194 GND.n2218 585
R7999 GND.n4084 GND.n2218 585
R8000 GND.n4195 GND.n2217 585
R8001 GND.n4133 GND.n2217 585
R8002 GND.n2276 GND.n2212 585
R8003 GND.n4136 GND.n2276 585
R8004 GND.n4199 GND.n2211 585
R8005 GND.n4075 GND.n2211 585
R8006 GND.n4200 GND.n2210 585
R8007 GND.n4143 GND.n2210 585
R8008 GND.n4201 GND.n2209 585
R8009 GND.n2265 GND.n2209 585
R8010 GND.n2294 GND.n2204 585
R8011 GND.n2298 GND.n2294 585
R8012 GND.n4205 GND.n2203 585
R8013 GND.n4067 GND.n2203 585
R8014 GND.n4206 GND.n2202 585
R8015 GND.n4053 GND.n2202 585
R8016 GND.n4207 GND.n2201 585
R8017 GND.n4056 GND.n2201 585
R8018 GND.n2309 GND.n2196 585
R8019 GND.n4050 GND.n2309 585
R8020 GND.n4211 GND.n2195 585
R8021 GND.n2321 GND.n2195 585
R8022 GND.n4212 GND.n2194 585
R8023 GND.n4041 GND.n2194 585
R8024 GND.n4213 GND.n2193 585
R8025 GND.n4028 GND.n2193 585
R8026 GND.n2328 GND.n2188 585
R8027 GND.n4031 GND.n2328 585
R8028 GND.n4217 GND.n2187 585
R8029 GND.n4026 GND.n2187 585
R8030 GND.n4218 GND.n2186 585
R8031 GND.n2344 GND.n2186 585
R8032 GND.n4219 GND.n2185 585
R8033 GND.n4017 GND.n2185 585
R8034 GND.n4003 GND.n2180 585
R8035 GND.n4004 GND.n4003 585
R8036 GND.n4223 GND.n2179 585
R8037 GND.n4007 GND.n2179 585
R8038 GND.n4224 GND.n2178 585
R8039 GND.n4001 GND.n2178 585
R8040 GND.n4225 GND.n2177 585
R8041 GND.n2367 GND.n2177 585
R8042 GND.n2363 GND.n2172 585
R8043 GND.n3992 GND.n2363 585
R8044 GND.n4229 GND.n2171 585
R8045 GND.n3978 GND.n2171 585
R8046 GND.n4230 GND.n2170 585
R8047 GND.n3982 GND.n2170 585
R8048 GND.n4231 GND.n2169 585
R8049 GND.n3918 GND.n2169 585
R8050 GND.n4375 GND.n1946 585
R8051 GND.n3784 GND.n1946 585
R8052 GND.n4377 GND.n4376 585
R8053 GND.n4378 GND.n4377 585
R8054 GND.n1947 GND.n1945 585
R8055 GND.n3719 GND.n1945 585
R8056 GND.n1925 GND.n1924 585
R8057 GND.n3717 GND.n1925 585
R8058 GND.n4388 GND.n4387 585
R8059 GND.n4387 GND.n4386 585
R8060 GND.n4389 GND.n1922 585
R8061 GND.n3711 GND.n1922 585
R8062 GND.n4391 GND.n4390 585
R8063 GND.n4392 GND.n4391 585
R8064 GND.n1923 GND.n1921 585
R8065 GND.n3707 GND.n1921 585
R8066 GND.n3678 GND.n3677 585
R8067 GND.n3678 GND.n2483 585
R8068 GND.n3680 GND.n3679 585
R8069 GND.n3679 GND.n1908 585
R8070 GND.n3681 GND.n3676 585
R8071 GND.n3676 GND.n1906 585
R8072 GND.n3683 GND.n3682 585
R8073 GND.n3684 GND.n3683 585
R8074 GND.n1887 GND.n1886 585
R8075 GND.n2496 GND.n1887 585
R8076 GND.n4409 GND.n4408 585
R8077 GND.n4408 GND.n4407 585
R8078 GND.n4410 GND.n1884 585
R8079 GND.n3666 GND.n1884 585
R8080 GND.n4412 GND.n4411 585
R8081 GND.n4413 GND.n4412 585
R8082 GND.n1885 GND.n1883 585
R8083 GND.n3662 GND.n1883 585
R8084 GND.n1861 GND.n1860 585
R8085 GND.n2501 GND.n1861 585
R8086 GND.n4422 GND.n4421 585
R8087 GND.n4421 GND.n4420 585
R8088 GND.n4423 GND.n1858 585
R8089 GND.n3629 GND.n1858 585
R8090 GND.n4425 GND.n4424 585
R8091 GND.n4426 GND.n4425 585
R8092 GND.n1859 GND.n1857 585
R8093 GND.n3633 GND.n1857 585
R8094 GND.n3645 GND.n3644 585
R8095 GND.n3646 GND.n3645 585
R8096 GND.n3643 GND.n2509 585
R8097 GND.n2509 GND.n1845 585
R8098 GND.n3642 GND.n3641 585
R8099 GND.n3641 GND.n3640 585
R8100 GND.n2511 GND.n2510 585
R8101 GND.n3622 GND.n2511 585
R8102 GND.n1832 GND.n1831 585
R8103 GND.n3624 GND.n1832 585
R8104 GND.n4443 GND.n4442 585
R8105 GND.n4442 GND.n4441 585
R8106 GND.n4444 GND.n1829 585
R8107 GND.n3611 GND.n1829 585
R8108 GND.n4446 GND.n4445 585
R8109 GND.n4447 GND.n4446 585
R8110 GND.n1830 GND.n1828 585
R8111 GND.n1828 GND.n1824 585
R8112 GND.n3603 GND.n3602 585
R8113 GND.n3604 GND.n3603 585
R8114 GND.n1813 GND.n1812 585
R8115 GND.n3555 GND.n1813 585
R8116 GND.n4457 GND.n4456 585
R8117 GND.n4456 GND.n4455 585
R8118 GND.n4458 GND.n1810 585
R8119 GND.n3581 GND.n1810 585
R8120 GND.n4460 GND.n4459 585
R8121 GND.n4461 GND.n4460 585
R8122 GND.n1811 GND.n1809 585
R8123 GND.n1809 GND.n1806 585
R8124 GND.n3571 GND.n3570 585
R8125 GND.n3572 GND.n3571 585
R8126 GND.n1794 GND.n1793 585
R8127 GND.n1798 GND.n1794 585
R8128 GND.n4471 GND.n4470 585
R8129 GND.n4470 GND.n4469 585
R8130 GND.n4472 GND.n1791 585
R8131 GND.n3549 GND.n1791 585
R8132 GND.n4474 GND.n4473 585
R8133 GND.n4475 GND.n4474 585
R8134 GND.n1792 GND.n1790 585
R8135 GND.n1790 GND.n1786 585
R8136 GND.n3539 GND.n3538 585
R8137 GND.n3540 GND.n3539 585
R8138 GND.n1774 GND.n1773 585
R8139 GND.n1778 GND.n1774 585
R8140 GND.n4485 GND.n4484 585
R8141 GND.n4484 GND.n4483 585
R8142 GND.n4486 GND.n1771 585
R8143 GND.n3503 GND.n1771 585
R8144 GND.n4488 GND.n4487 585
R8145 GND.n4489 GND.n4488 585
R8146 GND.n1772 GND.n1770 585
R8147 GND.n1770 GND.n1766 585
R8148 GND.n2562 GND.n2561 585
R8149 GND.n2563 GND.n2562 585
R8150 GND.n1754 GND.n1753 585
R8151 GND.n1758 GND.n1754 585
R8152 GND.n4499 GND.n4498 585
R8153 GND.n4498 GND.n4497 585
R8154 GND.n4500 GND.n1751 585
R8155 GND.n3489 GND.n1751 585
R8156 GND.n4502 GND.n4501 585
R8157 GND.n4503 GND.n4502 585
R8158 GND.n1752 GND.n1750 585
R8159 GND.n3479 GND.n1750 585
R8160 GND.n3355 GND.n3354 585
R8161 GND.n3355 GND.n3297 585
R8162 GND.n3356 GND.n3332 585
R8163 GND.n3359 GND.n3358 585
R8164 GND.n3360 GND.n3331 585
R8165 GND.n3331 GND.n1734 585
R8166 GND.n3362 GND.n3361 585
R8167 GND.n3364 GND.n3330 585
R8168 GND.n3367 GND.n3366 585
R8169 GND.n3368 GND.n3329 585
R8170 GND.n3370 GND.n3369 585
R8171 GND.n3372 GND.n3328 585
R8172 GND.n3375 GND.n3374 585
R8173 GND.n3376 GND.n3327 585
R8174 GND.n3378 GND.n3377 585
R8175 GND.n3380 GND.n3326 585
R8176 GND.n3383 GND.n3382 585
R8177 GND.n3384 GND.n3325 585
R8178 GND.n3386 GND.n3385 585
R8179 GND.n3388 GND.n3324 585
R8180 GND.n3391 GND.n3390 585
R8181 GND.n3392 GND.n3323 585
R8182 GND.n3394 GND.n3393 585
R8183 GND.n3396 GND.n3322 585
R8184 GND.n3399 GND.n3398 585
R8185 GND.n3400 GND.n3321 585
R8186 GND.n3402 GND.n3401 585
R8187 GND.n3404 GND.n3320 585
R8188 GND.n3407 GND.n3406 585
R8189 GND.n3409 GND.n3317 585
R8190 GND.n3411 GND.n3410 585
R8191 GND.n3413 GND.n3316 585
R8192 GND.n3414 GND.n1554 585
R8193 GND.n3419 GND.n3418 585
R8194 GND.n3421 GND.n3420 585
R8195 GND.n3423 GND.n3315 585
R8196 GND.n3426 GND.n3425 585
R8197 GND.n3427 GND.n3311 585
R8198 GND.n3429 GND.n3428 585
R8199 GND.n3431 GND.n3310 585
R8200 GND.n3434 GND.n3433 585
R8201 GND.n3435 GND.n3309 585
R8202 GND.n3437 GND.n3436 585
R8203 GND.n3439 GND.n3308 585
R8204 GND.n3442 GND.n3441 585
R8205 GND.n3443 GND.n3307 585
R8206 GND.n3445 GND.n3444 585
R8207 GND.n3447 GND.n3306 585
R8208 GND.n3450 GND.n3449 585
R8209 GND.n3451 GND.n3305 585
R8210 GND.n3453 GND.n3452 585
R8211 GND.n3455 GND.n3304 585
R8212 GND.n3458 GND.n3457 585
R8213 GND.n3459 GND.n3303 585
R8214 GND.n3461 GND.n3460 585
R8215 GND.n3463 GND.n3302 585
R8216 GND.n3466 GND.n3465 585
R8217 GND.n3467 GND.n3301 585
R8218 GND.n3469 GND.n3468 585
R8219 GND.n3471 GND.n3300 585
R8220 GND.n3472 GND.n3299 585
R8221 GND.n3475 GND.n3474 585
R8222 GND.n3781 GND.n2479 585
R8223 GND.n3780 GND.n3779 585
R8224 GND.n3778 GND.n3777 585
R8225 GND.n3776 GND.n3775 585
R8226 GND.n3774 GND.n3773 585
R8227 GND.n3772 GND.n3771 585
R8228 GND.n3770 GND.n3769 585
R8229 GND.n3768 GND.n3767 585
R8230 GND.n3766 GND.n3765 585
R8231 GND.n3764 GND.n3763 585
R8232 GND.n3762 GND.n3761 585
R8233 GND.n3760 GND.n3759 585
R8234 GND.n3758 GND.n3757 585
R8235 GND.n3756 GND.n3755 585
R8236 GND.n3754 GND.n3753 585
R8237 GND.n3752 GND.n3751 585
R8238 GND.n3750 GND.n3749 585
R8239 GND.n3748 GND.n3747 585
R8240 GND.n3746 GND.n3745 585
R8241 GND.n3744 GND.n3743 585
R8242 GND.n3742 GND.n3741 585
R8243 GND.n3740 GND.n3739 585
R8244 GND.n3738 GND.n3737 585
R8245 GND.n3736 GND.n3735 585
R8246 GND.n3734 GND.n3733 585
R8247 GND.n3732 GND.n3731 585
R8248 GND.n3730 GND.n3729 585
R8249 GND.n3728 GND.n3727 585
R8250 GND.n3726 GND.n2002 585
R8251 GND.n4315 GND.n4314 585
R8252 GND.n4317 GND.n4316 585
R8253 GND.n4319 GND.n4318 585
R8254 GND.n4321 GND.n4320 585
R8255 GND.n4324 GND.n4323 585
R8256 GND.n4326 GND.n4325 585
R8257 GND.n4328 GND.n4327 585
R8258 GND.n4330 GND.n4329 585
R8259 GND.n4332 GND.n4331 585
R8260 GND.n4334 GND.n4333 585
R8261 GND.n4336 GND.n4335 585
R8262 GND.n4338 GND.n4337 585
R8263 GND.n4340 GND.n4339 585
R8264 GND.n4342 GND.n4341 585
R8265 GND.n4344 GND.n4343 585
R8266 GND.n4346 GND.n4345 585
R8267 GND.n4348 GND.n4347 585
R8268 GND.n4350 GND.n4349 585
R8269 GND.n4352 GND.n4351 585
R8270 GND.n4354 GND.n4353 585
R8271 GND.n4356 GND.n4355 585
R8272 GND.n4358 GND.n4357 585
R8273 GND.n4360 GND.n4359 585
R8274 GND.n4362 GND.n4361 585
R8275 GND.n4364 GND.n4363 585
R8276 GND.n4366 GND.n4365 585
R8277 GND.n4367 GND.n1999 585
R8278 GND.n4369 GND.n4368 585
R8279 GND.n1968 GND.n1967 585
R8280 GND.n4373 GND.n4372 585
R8281 GND.n4372 GND.n4371 585
R8282 GND.n3783 GND.n3782 585
R8283 GND.n3784 GND.n3783 585
R8284 GND.n3722 GND.n1943 585
R8285 GND.n4378 GND.n1943 585
R8286 GND.n3721 GND.n3720 585
R8287 GND.n3720 GND.n3719 585
R8288 GND.n3716 GND.n3715 585
R8289 GND.n3717 GND.n3716 585
R8290 GND.n3714 GND.n1927 585
R8291 GND.n4386 GND.n1927 585
R8292 GND.n3713 GND.n3712 585
R8293 GND.n3712 GND.n3711 585
R8294 GND.n3710 GND.n1919 585
R8295 GND.n4392 GND.n1919 585
R8296 GND.n3709 GND.n3708 585
R8297 GND.n3708 GND.n3707 585
R8298 GND.n2481 GND.n2480 585
R8299 GND.n2483 GND.n2481 585
R8300 GND.n3672 GND.n3671 585
R8301 GND.n3671 GND.n1908 585
R8302 GND.n3673 GND.n2498 585
R8303 GND.n2498 GND.n1906 585
R8304 GND.n3675 GND.n3674 585
R8305 GND.n3684 GND.n3675 585
R8306 GND.n3670 GND.n2497 585
R8307 GND.n2497 GND.n2496 585
R8308 GND.n3669 GND.n1889 585
R8309 GND.n4407 GND.n1889 585
R8310 GND.n3668 GND.n3667 585
R8311 GND.n3667 GND.n3666 585
R8312 GND.n3665 GND.n1880 585
R8313 GND.n4413 GND.n1880 585
R8314 GND.n3664 GND.n3663 585
R8315 GND.n3663 GND.n3662 585
R8316 GND.n2500 GND.n2499 585
R8317 GND.n2501 GND.n2500 585
R8318 GND.n3628 GND.n1863 585
R8319 GND.n4420 GND.n1863 585
R8320 GND.n3631 GND.n3630 585
R8321 GND.n3630 GND.n3629 585
R8322 GND.n3632 GND.n1855 585
R8323 GND.n4426 GND.n1855 585
R8324 GND.n3635 GND.n3634 585
R8325 GND.n3634 GND.n3633 585
R8326 GND.n3636 GND.n2507 585
R8327 GND.n3646 GND.n2507 585
R8328 GND.n3637 GND.n2514 585
R8329 GND.n2514 GND.n1845 585
R8330 GND.n3639 GND.n3638 585
R8331 GND.n3640 GND.n3639 585
R8332 GND.n3627 GND.n2513 585
R8333 GND.n3622 GND.n2513 585
R8334 GND.n3626 GND.n3625 585
R8335 GND.n3625 GND.n3624 585
R8336 GND.n2515 GND.n1834 585
R8337 GND.n4441 GND.n1834 585
R8338 GND.n3610 GND.n3609 585
R8339 GND.n3611 GND.n3610 585
R8340 GND.n3608 GND.n1826 585
R8341 GND.n4447 GND.n1826 585
R8342 GND.n3607 GND.n3606 585
R8343 GND.n3606 GND.n1824 585
R8344 GND.n3605 GND.n2520 585
R8345 GND.n3605 GND.n3604 585
R8346 GND.n3577 GND.n2521 585
R8347 GND.n3555 GND.n2521 585
R8348 GND.n3578 GND.n1815 585
R8349 GND.n4455 GND.n1815 585
R8350 GND.n3580 GND.n3579 585
R8351 GND.n3581 GND.n3580 585
R8352 GND.n3576 GND.n1808 585
R8353 GND.n4461 GND.n1808 585
R8354 GND.n3575 GND.n3574 585
R8355 GND.n3574 GND.n1806 585
R8356 GND.n3573 GND.n2529 585
R8357 GND.n3573 GND.n3572 585
R8358 GND.n3545 GND.n2530 585
R8359 GND.n2530 GND.n1798 585
R8360 GND.n3546 GND.n1796 585
R8361 GND.n4469 GND.n1796 585
R8362 GND.n3548 GND.n3547 585
R8363 GND.n3549 GND.n3548 585
R8364 GND.n3544 GND.n1788 585
R8365 GND.n4475 GND.n1788 585
R8366 GND.n3543 GND.n3542 585
R8367 GND.n3542 GND.n1786 585
R8368 GND.n3541 GND.n2536 585
R8369 GND.n3541 GND.n3540 585
R8370 GND.n3499 GND.n2537 585
R8371 GND.n2537 GND.n1778 585
R8372 GND.n3500 GND.n1776 585
R8373 GND.n4483 GND.n1776 585
R8374 GND.n3502 GND.n3501 585
R8375 GND.n3503 GND.n3502 585
R8376 GND.n3498 GND.n1768 585
R8377 GND.n4489 GND.n1768 585
R8378 GND.n3497 GND.n3496 585
R8379 GND.n3496 GND.n1766 585
R8380 GND.n3495 GND.n2568 585
R8381 GND.n3495 GND.n2563 585
R8382 GND.n3494 GND.n3493 585
R8383 GND.n3494 GND.n1758 585
R8384 GND.n3492 GND.n1756 585
R8385 GND.n4497 GND.n1756 585
R8386 GND.n3491 GND.n3490 585
R8387 GND.n3490 GND.n3489 585
R8388 GND.n2569 GND.n1748 585
R8389 GND.n4503 GND.n1748 585
R8390 GND.n3478 GND.n3477 585
R8391 GND.n3479 GND.n3478 585
R8392 GND.n3476 GND.n3298 585
R8393 GND.n3298 GND.n3297 585
R8394 GND.n5526 GND.n5525 585
R8395 GND.n5526 GND.n861 585
R8396 GND.n5527 GND.n888 585
R8397 GND.n5527 GND.n860 585
R8398 GND.n5531 GND.n5530 585
R8399 GND.n5530 GND.n5529 585
R8400 GND.n5532 GND.n883 585
R8401 GND.n883 GND.n868 585
R8402 GND.n5534 GND.n5533 585
R8403 GND.n5535 GND.n5534 585
R8404 GND.n884 GND.n882 585
R8405 GND.n2240 GND.n882 585
R8406 GND.n4154 GND.n4153 585
R8407 GND.n4154 GND.n2239 585
R8408 GND.n4156 GND.n4155 585
R8409 GND.n4155 GND.n2250 585
R8410 GND.n4157 GND.n2254 585
R8411 GND.n2254 GND.n2247 585
R8412 GND.n4159 GND.n4158 585
R8413 GND.n4160 GND.n4159 585
R8414 GND.n4110 GND.n2253 585
R8415 GND.n4115 GND.n2253 585
R8416 GND.n4112 GND.n4111 585
R8417 GND.n4113 GND.n4112 585
R8418 GND.n4109 GND.n4108 585
R8419 GND.n4109 GND.n4102 585
R8420 GND.n4107 GND.n4089 585
R8421 GND.n4090 GND.n4089 585
R8422 GND.n4129 GND.n4128 585
R8423 GND.n4128 GND.n4127 585
R8424 GND.n4131 GND.n4130 585
R8425 GND.n4132 GND.n4131 585
R8426 GND.n4088 GND.n4087 585
R8427 GND.n4088 GND.n2281 585
R8428 GND.n4086 GND.n4085 585
R8429 GND.n4085 GND.n2275 585
R8430 GND.n2264 GND.n2262 585
R8431 GND.n2267 GND.n2264 585
R8432 GND.n4146 GND.n4145 585
R8433 GND.n4145 GND.n4144 585
R8434 GND.n2263 GND.n2261 585
R8435 GND.n2295 GND.n2263 585
R8436 GND.n3950 GND.n3946 585
R8437 GND.n3946 GND.n2291 585
R8438 GND.n3952 GND.n3951 585
R8439 GND.n3952 GND.n2290 585
R8440 GND.n3953 GND.n3945 585
R8441 GND.n3953 GND.n2306 585
R8442 GND.n3955 GND.n3954 585
R8443 GND.n3954 GND.n2304 585
R8444 GND.n3956 GND.n3940 585
R8445 GND.n3940 GND.n2308 585
R8446 GND.n3958 GND.n3957 585
R8447 GND.n3958 GND.n2317 585
R8448 GND.n3959 GND.n3939 585
R8449 GND.n3959 GND.n2316 585
R8450 GND.n3961 GND.n3960 585
R8451 GND.n3960 GND.n2330 585
R8452 GND.n3962 GND.n3934 585
R8453 GND.n3934 GND.n2327 585
R8454 GND.n3964 GND.n3963 585
R8455 GND.n3964 GND.n2333 585
R8456 GND.n3965 GND.n3933 585
R8457 GND.n3965 GND.n2341 585
R8458 GND.n3967 GND.n3966 585
R8459 GND.n3966 GND.n2340 585
R8460 GND.n3968 GND.n3928 585
R8461 GND.n3928 GND.n2352 585
R8462 GND.n3970 GND.n3969 585
R8463 GND.n3970 GND.n2350 585
R8464 GND.n3971 GND.n3927 585
R8465 GND.n3971 GND.n2355 585
R8466 GND.n3973 GND.n3972 585
R8467 GND.n3972 GND.n2364 585
R8468 GND.n3974 GND.n2416 585
R8469 GND.n2416 GND.n2362 585
R8470 GND.n3976 GND.n3975 585
R8471 GND.n3977 GND.n3976 585
R8472 GND.n2417 GND.n2415 585
R8473 GND.n2415 GND.n2413 585
R8474 GND.n3921 GND.n3920 585
R8475 GND.n3920 GND.n3919 585
R8476 GND.n3912 GND.n2419 585
R8477 GND.n3912 GND.n2038 585
R8478 GND.n3911 GND.n3910 585
R8479 GND.n3911 GND.n2011 585
R8480 GND.n2421 GND.n2420 585
R8481 GND.n3903 GND.n2420 585
R8482 GND.n3906 GND.n3905 585
R8483 GND.n3905 GND.n3904 585
R8484 GND.n3880 GND.n2423 585
R8485 GND.n3881 GND.n3880 585
R8486 GND.n3879 GND.n3878 585
R8487 GND.n3879 GND.n2109 585
R8488 GND.n2425 GND.n2424 585
R8489 GND.n2424 GND.n2108 585
R8490 GND.n3874 GND.n3873 585
R8491 GND.n3873 GND.n3872 585
R8492 GND.n2428 GND.n2427 585
R8493 GND.n2437 GND.n2428 585
R8494 GND.n3860 GND.n3859 585
R8495 GND.n3861 GND.n3860 585
R8496 GND.n2440 GND.n2439 585
R8497 GND.n2439 GND.n2435 585
R8498 GND.n3855 GND.n3854 585
R8499 GND.n3854 GND.n3853 585
R8500 GND.n2443 GND.n2442 585
R8501 GND.n2452 GND.n2443 585
R8502 GND.n3824 GND.n2462 585
R8503 GND.n2462 GND.n2451 585
R8504 GND.n3826 GND.n3825 585
R8505 GND.n3827 GND.n3826 585
R8506 GND.n2463 GND.n2461 585
R8507 GND.n3815 GND.n2461 585
R8508 GND.n3819 GND.n3818 585
R8509 GND.n3818 GND.n3817 585
R8510 GND.n2470 GND.n2465 585
R8511 GND.n2478 GND.n2470 585
R8512 GND.n2469 GND.n2468 585
R8513 GND.n2469 GND.n1969 585
R8514 GND.n1941 GND.n1940 585
R8515 GND.n3785 GND.n1941 585
R8516 GND.n4381 GND.n4380 585
R8517 GND.n4380 GND.n4379 585
R8518 GND.n4382 GND.n1930 585
R8519 GND.n3718 GND.n1930 585
R8520 GND.n4384 GND.n4383 585
R8521 GND.n4385 GND.n4384 585
R8522 GND.n1931 GND.n1929 585
R8523 GND.n1929 GND.n1920 585
R8524 GND.n1934 GND.n1933 585
R8525 GND.n1933 GND.n1917 585
R8526 GND.n1905 GND.n1904 585
R8527 GND.n2482 GND.n1905 585
R8528 GND.n4402 GND.n4401 585
R8529 GND.n4401 GND.n4400 585
R8530 GND.n4403 GND.n1891 585
R8531 GND.n2489 GND.n1891 585
R8532 GND.n4405 GND.n4404 585
R8533 GND.n4406 GND.n4405 585
R8534 GND.n1892 GND.n1890 585
R8535 GND.n1890 GND.n1882 585
R8536 GND.n1898 GND.n1897 585
R8537 GND.n1897 GND.n1879 585
R8538 GND.n1896 GND.n1895 585
R8539 GND.n1896 GND.n1865 585
R8540 GND.n1853 GND.n1852 585
R8541 GND.n1862 GND.n1853 585
R8542 GND.n4429 GND.n4428 585
R8543 GND.n4428 GND.n4427 585
R8544 GND.n4430 GND.n1847 585
R8545 GND.n2508 GND.n1847 585
R8546 GND.n4432 GND.n4431 585
R8547 GND.n4433 GND.n4432 585
R8548 GND.n1848 GND.n1846 585
R8549 GND.n2512 GND.n1846 585
R8550 GND.n3595 GND.n3594 585
R8551 GND.n3595 GND.n1836 585
R8552 GND.n3597 GND.n3596 585
R8553 GND.n3596 GND.n1833 585
R8554 GND.n3598 GND.n2523 585
R8555 GND.n2523 GND.n1827 585
R8556 GND.n3600 GND.n3599 585
R8557 GND.n3601 GND.n3600 585
R8558 GND.n2524 GND.n2522 585
R8559 GND.n3556 GND.n2522 585
R8560 GND.n3586 GND.n3585 585
R8561 GND.n3585 GND.n1814 585
R8562 GND.n3584 GND.n2526 585
R8563 GND.n3584 GND.n3583 585
R8564 GND.n3528 GND.n2527 585
R8565 GND.n3569 GND.n2527 585
R8566 GND.n3530 GND.n3529 585
R8567 GND.n3530 GND.n2531 585
R8568 GND.n3532 GND.n3531 585
R8569 GND.n3531 GND.n1795 585
R8570 GND.n3533 GND.n2541 585
R8571 GND.n2541 GND.n1789 585
R8572 GND.n3535 GND.n3534 585
R8573 GND.n3536 GND.n3535 585
R8574 GND.n2542 GND.n2540 585
R8575 GND.n2540 GND.n2538 585
R8576 GND.n3520 GND.n3519 585
R8577 GND.n3519 GND.n1775 585
R8578 GND.n3518 GND.n2544 585
R8579 GND.n3518 GND.n1769 585
R8580 GND.n3517 GND.n2559 585
R8581 GND.n3517 GND.n3516 585
R8582 GND.n2546 GND.n2545 585
R8583 GND.n2560 GND.n2545 585
R8584 GND.n2555 GND.n2554 585
R8585 GND.n2554 GND.n1755 585
R8586 GND.n2553 GND.n2548 585
R8587 GND.n2553 GND.n1749 585
R8588 GND.n2552 GND.n2551 585
R8589 GND.n2552 GND.n1746 585
R8590 GND.n1733 GND.n1732 585
R8591 GND.n3296 GND.n1733 585
R8592 GND.n4513 GND.n4512 585
R8593 GND.n4512 GND.n4511 585
R8594 GND.n4514 GND.n1725 585
R8595 GND.n2574 GND.n1725 585
R8596 GND.n4516 GND.n4515 585
R8597 GND.n4517 GND.n4516 585
R8598 GND.n1726 GND.n1724 585
R8599 GND.n1724 GND.n1721 585
R8600 GND.n1706 GND.n1705 585
R8601 GND.n1710 GND.n1706 585
R8602 GND.n4527 GND.n4526 585
R8603 GND.n4526 GND.n4525 585
R8604 GND.n4528 GND.n1698 585
R8605 GND.n1707 GND.n1698 585
R8606 GND.n4530 GND.n4529 585
R8607 GND.n4531 GND.n4530 585
R8608 GND.n1699 GND.n1697 585
R8609 GND.n1697 GND.n1694 585
R8610 GND.n1680 GND.n1679 585
R8611 GND.n1682 GND.n1680 585
R8612 GND.n4541 GND.n4540 585
R8613 GND.n4540 GND.n4539 585
R8614 GND.n4542 GND.n1672 585
R8615 GND.n3271 GND.n1672 585
R8616 GND.n4544 GND.n4543 585
R8617 GND.n4545 GND.n4544 585
R8618 GND.n1673 GND.n1671 585
R8619 GND.n1671 GND.n1668 585
R8620 GND.n1647 GND.n1646 585
R8621 GND.n1665 GND.n1647 585
R8622 GND.n4553 GND.n4552 585
R8623 GND.n4552 GND.n4551 585
R8624 GND.n4554 GND.n1641 585
R8625 GND.n1641 GND.n1639 585
R8626 GND.n4556 GND.n4555 585
R8627 GND.n4557 GND.n4556 585
R8628 GND.n1642 GND.n1640 585
R8629 GND.n1640 GND.n1627 585
R8630 GND.n3199 GND.n3198 585
R8631 GND.n3199 GND.n1527 585
R8632 GND.n3201 GND.n3200 585
R8633 GND.n3200 GND.n1525 585
R8634 GND.n3202 GND.n2612 585
R8635 GND.n2612 GND.n2592 585
R8636 GND.n3204 GND.n3203 585
R8637 GND.n3205 GND.n3204 585
R8638 GND.n2613 GND.n2611 585
R8639 GND.n2611 GND.n2601 585
R8640 GND.n3190 GND.n3189 585
R8641 GND.n3189 GND.n2599 585
R8642 GND.n3188 GND.n2615 585
R8643 GND.n3188 GND.n2604 585
R8644 GND.n3187 GND.n2617 585
R8645 GND.n3187 GND.n3186 585
R8646 GND.n3049 GND.n2616 585
R8647 GND.n2627 GND.n2616 585
R8648 GND.n3051 GND.n3050 585
R8649 GND.n3050 GND.n2625 585
R8650 GND.n3052 GND.n3042 585
R8651 GND.n3042 GND.n3041 585
R8652 GND.n3054 GND.n3053 585
R8653 GND.n3054 GND.n2638 585
R8654 GND.n3055 GND.n3039 585
R8655 GND.n3055 GND.n2636 585
R8656 GND.n3057 GND.n3056 585
R8657 GND.n3056 GND.n2648 585
R8658 GND.n3058 GND.n3034 585
R8659 GND.n3034 GND.n2646 585
R8660 GND.n3063 GND.n3059 585
R8661 GND.n3063 GND.n3062 585
R8662 GND.n3064 GND.n3033 585
R8663 GND.n3064 GND.n2657 585
R8664 GND.n3066 GND.n3065 585
R8665 GND.n3065 GND.n2656 585
R8666 GND.n3067 GND.n3028 585
R8667 GND.n3028 GND.n2667 585
R8668 GND.n3069 GND.n3068 585
R8669 GND.n3069 GND.n2665 585
R8670 GND.n3072 GND.n3027 585
R8671 GND.n3072 GND.n3071 585
R8672 GND.n3074 GND.n3073 585
R8673 GND.n3073 GND.n2677 585
R8674 GND.n3075 GND.n3023 585
R8675 GND.n3023 GND.n2676 585
R8676 GND.n3078 GND.n3077 585
R8677 GND.n3079 GND.n3078 585
R8678 GND.n3025 GND.n3022 585
R8679 GND.n3022 GND.n2720 585
R8680 GND.n2704 GND.n2703 585
R8681 GND.n2708 GND.n2704 585
R8682 GND.n3091 GND.n3090 585
R8683 GND.n3090 GND.n3089 585
R8684 GND.n3093 GND.n2701 585
R8685 GND.n2705 GND.n2701 585
R8686 GND.n3095 GND.n3094 585
R8687 GND.n3096 GND.n3095 585
R8688 GND.n2998 GND.n2700 585
R8689 GND.n2700 GND.n2694 585
R8690 GND.n2999 GND.n2732 585
R8691 GND.n2732 GND.n2692 585
R8692 GND.n3002 GND.n3001 585
R8693 GND.n3003 GND.n3002 585
R8694 GND.n2997 GND.n2731 585
R8695 GND.n2962 GND.n2731 585
R8696 GND.n2737 GND.n2733 585
R8697 GND.n2961 GND.n2737 585
R8698 GND.n2993 GND.n2992 585
R8699 GND.n2992 GND.n2991 585
R8700 GND.n2736 GND.n2735 585
R8701 GND.n2752 GND.n2736 585
R8702 GND.n2783 GND.n2782 585
R8703 GND.n2783 GND.n2749 585
R8704 GND.n2784 GND.n2779 585
R8705 GND.n2784 GND.n2755 585
R8706 GND.n2786 GND.n2785 585
R8707 GND.n2785 GND.n2763 585
R8708 GND.n2787 GND.n2774 585
R8709 GND.n2774 GND.n2762 585
R8710 GND.n2789 GND.n2788 585
R8711 GND.n2790 GND.n2789 585
R8712 GND.n4307 GND.n4306 585
R8713 GND.n4308 GND.n4307 585
R8714 GND.n4305 GND.n2040 585
R8715 GND.n2048 GND.n2042 585
R8716 GND.n4298 GND.n2049 585
R8717 GND.n4297 GND.n2050 585
R8718 GND.n2052 GND.n2051 585
R8719 GND.n4290 GND.n2058 585
R8720 GND.n4289 GND.n2059 585
R8721 GND.n2066 GND.n2060 585
R8722 GND.n4282 GND.n2067 585
R8723 GND.n4281 GND.n2068 585
R8724 GND.n2070 GND.n2069 585
R8725 GND.n4274 GND.n2076 585
R8726 GND.n4273 GND.n2077 585
R8727 GND.n4262 GND.n2078 585
R8728 GND.n4266 GND.n4263 585
R8729 GND.n4261 GND.n2084 585
R8730 GND.n5653 GND.n5652 585
R8731 GND.n5652 GND.n715 585
R8732 GND.n5606 GND.n802 585
R8733 GND.n5606 GND.n5605 585
R8734 GND.n815 GND.n803 585
R8735 GND.n804 GND.n803 585
R8736 GND.n5595 GND.n5594 585
R8737 GND.n5596 GND.n5595 585
R8738 GND.n814 GND.n813 585
R8739 GND.n813 GND.n810 585
R8740 GND.n835 GND.n821 585
R8741 GND.n5586 GND.n821 585
R8742 GND.n833 GND.n831 585
R8743 GND.n831 GND.n820 585
R8744 GND.n5577 GND.n5576 585
R8745 GND.n5578 GND.n5577 585
R8746 GND.n832 GND.n830 585
R8747 GND.n830 GND.n827 585
R8748 GND.n855 GND.n840 585
R8749 GND.n5569 GND.n840 585
R8750 GND.n853 GND.n851 585
R8751 GND.n851 GND.n849 585
R8752 GND.n5560 GND.n5559 585
R8753 GND.n5561 GND.n5560 585
R8754 GND.n852 GND.n850 585
R8755 GND.n850 GND.n846 585
R8756 GND.n876 GND.n862 585
R8757 GND.n5552 GND.n862 585
R8758 GND.n874 GND.n872 585
R8759 GND.n5528 GND.n872 585
R8760 GND.n5543 GND.n5542 585
R8761 GND.n5544 GND.n5543 585
R8762 GND.n873 GND.n871 585
R8763 GND.n5536 GND.n871 585
R8764 GND.n4178 GND.n4177 585
R8765 GND.n4177 GND.n881 585
R8766 GND.n4176 GND.n2236 585
R8767 GND.n4176 GND.n4175 585
R8768 GND.n2238 GND.n2237 585
R8769 GND.n2249 GND.n2238 585
R8770 GND.n4164 GND.n2231 585
R8771 GND.n4165 GND.n4164 585
R8772 GND.n4163 GND.n2230 585
R8773 GND.n4163 GND.n4162 585
R8774 GND.n2251 GND.n2229 585
R8775 GND.n2252 GND.n2251 585
R8776 GND.n4117 GND.n4106 585
R8777 GND.n4117 GND.n4116 585
R8778 GND.n4118 GND.n2223 585
R8779 GND.n4119 GND.n4118 585
R8780 GND.n4105 GND.n2222 585
R8781 GND.n4105 GND.n4104 585
R8782 GND.n4091 GND.n2221 585
R8783 GND.n4126 GND.n4091 585
R8784 GND.n2280 GND.n2279 585
R8785 GND.n4084 GND.n2280 585
R8786 GND.n4134 GND.n2215 585
R8787 GND.n4134 GND.n4133 585
R8788 GND.n4135 GND.n2214 585
R8789 GND.n4136 GND.n4135 585
R8790 GND.n2278 GND.n2213 585
R8791 GND.n4075 GND.n2278 585
R8792 GND.n2269 GND.n2268 585
R8793 GND.n4143 GND.n2269 585
R8794 GND.n2296 GND.n2207 585
R8795 GND.n2296 GND.n2265 585
R8796 GND.n2297 GND.n2206 585
R8797 GND.n2298 GND.n2297 585
R8798 GND.n2292 GND.n2205 585
R8799 GND.n4067 GND.n2292 585
R8800 GND.n4054 GND.n4052 585
R8801 GND.n4054 GND.n4053 585
R8802 GND.n4055 GND.n2199 585
R8803 GND.n4056 GND.n4055 585
R8804 GND.n4051 GND.n2198 585
R8805 GND.n4051 GND.n4050 585
R8806 GND.n2307 GND.n2197 585
R8807 GND.n2321 GND.n2307 585
R8808 GND.n2319 GND.n2318 585
R8809 GND.n4041 GND.n2319 585
R8810 GND.n4029 GND.n2191 585
R8811 GND.n4029 GND.n4028 585
R8812 GND.n4030 GND.n2190 585
R8813 GND.n4031 GND.n4030 585
R8814 GND.n4027 GND.n2189 585
R8815 GND.n4027 GND.n4026 585
R8816 GND.n2332 GND.n2331 585
R8817 GND.n2344 GND.n2332 585
R8818 GND.n2342 GND.n2183 585
R8819 GND.n4017 GND.n2342 585
R8820 GND.n4005 GND.n2182 585
R8821 GND.n4005 GND.n4004 585
R8822 GND.n4006 GND.n2181 585
R8823 GND.n4007 GND.n4006 585
R8824 GND.n4002 GND.n2354 585
R8825 GND.n4002 GND.n4001 585
R8826 GND.n2353 GND.n2175 585
R8827 GND.n2367 GND.n2353 585
R8828 GND.n2365 GND.n2174 585
R8829 GND.n3992 GND.n2365 585
R8830 GND.n3979 GND.n2173 585
R8831 GND.n3979 GND.n3978 585
R8832 GND.n3981 GND.n3980 585
R8833 GND.n3982 GND.n3981 585
R8834 GND.n2114 GND.n2039 585
R8835 GND.n3918 GND.n2039 585
R8836 GND.n5715 GND.n5714 585
R8837 GND.n5714 GND.n5713 585
R8838 GND.n714 GND.n713 585
R8839 GND.n5628 GND.n5627 585
R8840 GND.n5626 GND.n5625 585
R8841 GND.n5632 GND.n5624 585
R8842 GND.n5633 GND.n5623 585
R8843 GND.n5634 GND.n5622 585
R8844 GND.n5621 GND.n5619 585
R8845 GND.n5638 GND.n5618 585
R8846 GND.n5639 GND.n5617 585
R8847 GND.n5640 GND.n5616 585
R8848 GND.n5615 GND.n5613 585
R8849 GND.n5644 GND.n5612 585
R8850 GND.n5645 GND.n5611 585
R8851 GND.n5646 GND.n5610 585
R8852 GND.n5609 GND.n5607 585
R8853 GND.n5651 GND.n5650 585
R8854 GND.n5718 GND.n709 585
R8855 GND.n715 GND.n709 585
R8856 GND.n5719 GND.n708 585
R8857 GND.n5605 GND.n708 585
R8858 GND.n5720 GND.n707 585
R8859 GND.n804 GND.n707 585
R8860 GND.n812 GND.n705 585
R8861 GND.n5596 GND.n812 585
R8862 GND.n5724 GND.n704 585
R8863 GND.n810 GND.n704 585
R8864 GND.n5725 GND.n703 585
R8865 GND.n5586 GND.n703 585
R8866 GND.n5726 GND.n702 585
R8867 GND.n820 GND.n702 585
R8868 GND.n829 GND.n700 585
R8869 GND.n5578 GND.n829 585
R8870 GND.n5730 GND.n699 585
R8871 GND.n827 GND.n699 585
R8872 GND.n5731 GND.n698 585
R8873 GND.n5569 GND.n698 585
R8874 GND.n5732 GND.n697 585
R8875 GND.n849 GND.n697 585
R8876 GND.n848 GND.n695 585
R8877 GND.n5561 GND.n848 585
R8878 GND.n5736 GND.n694 585
R8879 GND.n846 GND.n694 585
R8880 GND.n5737 GND.n693 585
R8881 GND.n5552 GND.n693 585
R8882 GND.n5738 GND.n692 585
R8883 GND.n5528 GND.n692 585
R8884 GND.n870 GND.n690 585
R8885 GND.n5544 GND.n870 585
R8886 GND.n5742 GND.n689 585
R8887 GND.n5536 GND.n689 585
R8888 GND.n5743 GND.n688 585
R8889 GND.n881 GND.n688 585
R8890 GND.n5744 GND.n687 585
R8891 GND.n4175 GND.n687 585
R8892 GND.n2248 GND.n685 585
R8893 GND.n2249 GND.n2248 585
R8894 GND.n5748 GND.n684 585
R8895 GND.n4165 GND.n684 585
R8896 GND.n5749 GND.n683 585
R8897 GND.n4162 GND.n683 585
R8898 GND.n5750 GND.n682 585
R8899 GND.n2252 GND.n682 585
R8900 GND.n4114 GND.n680 585
R8901 GND.n4116 GND.n4114 585
R8902 GND.n5754 GND.n679 585
R8903 GND.n4119 GND.n679 585
R8904 GND.n5755 GND.n678 585
R8905 GND.n4104 GND.n678 585
R8906 GND.n5756 GND.n677 585
R8907 GND.n4126 GND.n677 585
R8908 GND.n4083 GND.n676 585
R8909 GND.n4084 GND.n4083 585
R8910 GND.n4082 GND.n4081 585
R8911 GND.n4133 GND.n4082 585
R8912 GND.n2282 GND.n2277 585
R8913 GND.n4136 GND.n2277 585
R8914 GND.n4077 GND.n4076 585
R8915 GND.n4076 GND.n4075 585
R8916 GND.n4074 GND.n2266 585
R8917 GND.n4143 GND.n2266 585
R8918 GND.n4073 GND.n2285 585
R8919 GND.n2285 GND.n2265 585
R8920 GND.n2289 GND.n2284 585
R8921 GND.n2298 GND.n2289 585
R8922 GND.n4069 GND.n4068 585
R8923 GND.n4068 GND.n4067 585
R8924 GND.n2288 GND.n2287 585
R8925 GND.n4053 GND.n2288 585
R8926 GND.n2312 GND.n2305 585
R8927 GND.n4056 GND.n2305 585
R8928 GND.n4049 GND.n4048 585
R8929 GND.n4050 GND.n4049 585
R8930 GND.n2311 GND.n2310 585
R8931 GND.n2321 GND.n2310 585
R8932 GND.n4043 GND.n4042 585
R8933 GND.n4042 GND.n4041 585
R8934 GND.n2315 GND.n2314 585
R8935 GND.n4028 GND.n2315 585
R8936 GND.n2336 GND.n2329 585
R8937 GND.n4031 GND.n2329 585
R8938 GND.n4025 GND.n4024 585
R8939 GND.n4026 GND.n4025 585
R8940 GND.n2335 GND.n2334 585
R8941 GND.n2344 GND.n2334 585
R8942 GND.n4019 GND.n4018 585
R8943 GND.n4018 GND.n4017 585
R8944 GND.n2339 GND.n2338 585
R8945 GND.n4004 GND.n2339 585
R8946 GND.n2358 GND.n2351 585
R8947 GND.n4007 GND.n2351 585
R8948 GND.n4000 GND.n3999 585
R8949 GND.n4001 GND.n4000 585
R8950 GND.n2357 GND.n2356 585
R8951 GND.n2367 GND.n2356 585
R8952 GND.n3994 GND.n3993 585
R8953 GND.n3993 GND.n3992 585
R8954 GND.n2361 GND.n2360 585
R8955 GND.n3978 GND.n2361 585
R8956 GND.n3913 GND.n2414 585
R8957 GND.n3982 GND.n2414 585
R8958 GND.n3917 GND.n3916 585
R8959 GND.n3918 GND.n3917 585
R8960 GND.n4966 GND.n4965 523.639
R8961 GND.n4372 GND.n1946 521.33
R8962 GND.n3783 GND.n2479 521.33
R8963 GND.n3474 GND.n3298 521.33
R8964 GND.n3356 GND.n3355 521.33
R8965 GND.n3312 GND.t34 347.526
R8966 GND.n3723 GND.t58 347.526
R8967 GND.n3318 GND.t75 347.526
R8968 GND.n2000 GND.t90 347.526
R8969 GND.n95 GND.n69 289.615
R8970 GND.n132 GND.n106 289.615
R8971 GND.n164 GND.n138 289.615
R8972 GND.n201 GND.n175 289.615
R8973 GND.n26 GND.n0 289.615
R8974 GND.n63 GND.n37 289.615
R8975 GND.n528 GND.n502 289.615
R8976 GND.n491 GND.n465 289.615
R8977 GND.n597 GND.n571 289.615
R8978 GND.n560 GND.n534 289.615
R8979 GND.n667 GND.n641 289.615
R8980 GND.n630 GND.n604 289.615
R8981 GND.n331 GND.n305 289.615
R8982 GND.n299 GND.n273 289.615
R8983 GND.n267 GND.n241 289.615
R8984 GND.n236 GND.n210 289.615
R8985 GND.n458 GND.n432 289.615
R8986 GND.n426 GND.n400 289.615
R8987 GND.n394 GND.n368 289.615
R8988 GND.n363 GND.n337 289.615
R8989 GND.n711 GND.t62 279.217
R8990 GND.n767 GND.t87 279.217
R8991 GND.n794 GND.t72 279.217
R8992 GND.n1550 GND.t84 279.217
R8993 GND.n1576 GND.t66 279.217
R8994 GND.n1618 GND.t42 279.217
R8995 GND.n2821 GND.t55 279.217
R8996 GND.n2097 GND.t109 279.217
R8997 GND.n3253 GND.t102 279.217
R8998 GND.n2006 GND.t24 279.217
R8999 GND.n2118 GND.t99 279.217
R9000 GND.n1395 GND.t52 279.217
R9001 GND.n1415 GND.t38 279.217
R9002 GND.n4264 GND.t46 279.217
R9003 GND.n4967 GND.n4966 270.271
R9004 GND.n4967 GND.n1217 270.271
R9005 GND.n4975 GND.n1217 270.271
R9006 GND.n4976 GND.n4975 270.271
R9007 GND.n4977 GND.n4976 270.271
R9008 GND.n4977 GND.n1211 270.271
R9009 GND.n4985 GND.n1211 270.271
R9010 GND.n4986 GND.n4985 270.271
R9011 GND.n4987 GND.n4986 270.271
R9012 GND.n4987 GND.n1205 270.271
R9013 GND.n4995 GND.n1205 270.271
R9014 GND.n4996 GND.n4995 270.271
R9015 GND.n4997 GND.n4996 270.271
R9016 GND.n4997 GND.n1199 270.271
R9017 GND.n5005 GND.n1199 270.271
R9018 GND.n5006 GND.n5005 270.271
R9019 GND.n5007 GND.n5006 270.271
R9020 GND.n5007 GND.n1193 270.271
R9021 GND.n5015 GND.n1193 270.271
R9022 GND.n5016 GND.n5015 270.271
R9023 GND.n5017 GND.n5016 270.271
R9024 GND.n5017 GND.n1187 270.271
R9025 GND.n5025 GND.n1187 270.271
R9026 GND.n5026 GND.n5025 270.271
R9027 GND.n5027 GND.n5026 270.271
R9028 GND.n5027 GND.n1181 270.271
R9029 GND.n5035 GND.n1181 270.271
R9030 GND.n5036 GND.n5035 270.271
R9031 GND.n5037 GND.n5036 270.271
R9032 GND.n5037 GND.n1175 270.271
R9033 GND.n5045 GND.n1175 270.271
R9034 GND.n5046 GND.n5045 270.271
R9035 GND.n5047 GND.n5046 270.271
R9036 GND.n5047 GND.n1169 270.271
R9037 GND.n5055 GND.n1169 270.271
R9038 GND.n5056 GND.n5055 270.271
R9039 GND.n5057 GND.n5056 270.271
R9040 GND.n5057 GND.n1163 270.271
R9041 GND.n5065 GND.n1163 270.271
R9042 GND.n5066 GND.n5065 270.271
R9043 GND.n5067 GND.n5066 270.271
R9044 GND.n5067 GND.n1157 270.271
R9045 GND.n5075 GND.n1157 270.271
R9046 GND.n5076 GND.n5075 270.271
R9047 GND.n5077 GND.n5076 270.271
R9048 GND.n5077 GND.n1151 270.271
R9049 GND.n5085 GND.n1151 270.271
R9050 GND.n5086 GND.n5085 270.271
R9051 GND.n5087 GND.n5086 270.271
R9052 GND.n5087 GND.n1145 270.271
R9053 GND.n5095 GND.n1145 270.271
R9054 GND.n5096 GND.n5095 270.271
R9055 GND.n5097 GND.n5096 270.271
R9056 GND.n5097 GND.n1139 270.271
R9057 GND.n5105 GND.n1139 270.271
R9058 GND.n5106 GND.n5105 270.271
R9059 GND.n5107 GND.n5106 270.271
R9060 GND.n5107 GND.n1133 270.271
R9061 GND.n5115 GND.n1133 270.271
R9062 GND.n5116 GND.n5115 270.271
R9063 GND.n5117 GND.n5116 270.271
R9064 GND.n5117 GND.n1127 270.271
R9065 GND.n5125 GND.n1127 270.271
R9066 GND.n5126 GND.n5125 270.271
R9067 GND.n5127 GND.n5126 270.271
R9068 GND.n5127 GND.n1121 270.271
R9069 GND.n5135 GND.n1121 270.271
R9070 GND.n5136 GND.n5135 270.271
R9071 GND.n5137 GND.n5136 270.271
R9072 GND.n5137 GND.n1115 270.271
R9073 GND.n5145 GND.n1115 270.271
R9074 GND.n5146 GND.n5145 270.271
R9075 GND.n5147 GND.n5146 270.271
R9076 GND.n5147 GND.n1109 270.271
R9077 GND.n5155 GND.n1109 270.271
R9078 GND.n5156 GND.n5155 270.271
R9079 GND.n5157 GND.n5156 270.271
R9080 GND.n5157 GND.n1103 270.271
R9081 GND.n5165 GND.n1103 270.271
R9082 GND.n5166 GND.n5165 270.271
R9083 GND.n5167 GND.n5166 270.271
R9084 GND.n5167 GND.n1097 270.271
R9085 GND.n5175 GND.n1097 270.271
R9086 GND.n5176 GND.n5175 270.271
R9087 GND.n5177 GND.n5176 270.271
R9088 GND.n5177 GND.n1091 270.271
R9089 GND.n5185 GND.n1091 270.271
R9090 GND.n5186 GND.n5185 270.271
R9091 GND.n5187 GND.n5186 270.271
R9092 GND.n5187 GND.n1085 270.271
R9093 GND.n5195 GND.n1085 270.271
R9094 GND.n5196 GND.n5195 270.271
R9095 GND.n5197 GND.n5196 270.271
R9096 GND.n5197 GND.n1079 270.271
R9097 GND.n5205 GND.n1079 270.271
R9098 GND.n5206 GND.n5205 270.271
R9099 GND.n5207 GND.n5206 270.271
R9100 GND.n5207 GND.n1073 270.271
R9101 GND.n5215 GND.n1073 270.271
R9102 GND.n5216 GND.n5215 270.271
R9103 GND.n5217 GND.n5216 270.271
R9104 GND.n5217 GND.n1067 270.271
R9105 GND.n5225 GND.n1067 270.271
R9106 GND.n5226 GND.n5225 270.271
R9107 GND.n5227 GND.n5226 270.271
R9108 GND.n5227 GND.n1061 270.271
R9109 GND.n5235 GND.n1061 270.271
R9110 GND.n5236 GND.n5235 270.271
R9111 GND.n5237 GND.n5236 270.271
R9112 GND.n5237 GND.n1055 270.271
R9113 GND.n5245 GND.n1055 270.271
R9114 GND.n5246 GND.n5245 270.271
R9115 GND.n5247 GND.n5246 270.271
R9116 GND.n5247 GND.n1049 270.271
R9117 GND.n5255 GND.n1049 270.271
R9118 GND.n5256 GND.n5255 270.271
R9119 GND.n5257 GND.n5256 270.271
R9120 GND.n5257 GND.n1043 270.271
R9121 GND.n5265 GND.n1043 270.271
R9122 GND.n5266 GND.n5265 270.271
R9123 GND.n5267 GND.n5266 270.271
R9124 GND.n5267 GND.n1037 270.271
R9125 GND.n5275 GND.n1037 270.271
R9126 GND.n5276 GND.n5275 270.271
R9127 GND.n5277 GND.n5276 270.271
R9128 GND.n5277 GND.n1031 270.271
R9129 GND.n5285 GND.n1031 270.271
R9130 GND.n5286 GND.n5285 270.271
R9131 GND.n5287 GND.n5286 270.271
R9132 GND.n5287 GND.n1025 270.271
R9133 GND.n5295 GND.n1025 270.271
R9134 GND.n5296 GND.n5295 270.271
R9135 GND.n5297 GND.n5296 270.271
R9136 GND.n5297 GND.n1019 270.271
R9137 GND.n5305 GND.n1019 270.271
R9138 GND.n5306 GND.n5305 270.271
R9139 GND.n5307 GND.n5306 270.271
R9140 GND.n5307 GND.n1013 270.271
R9141 GND.n5315 GND.n1013 270.271
R9142 GND.n5316 GND.n5315 270.271
R9143 GND.n5317 GND.n5316 270.271
R9144 GND.n5317 GND.n1007 270.271
R9145 GND.n5325 GND.n1007 270.271
R9146 GND.n5326 GND.n5325 270.271
R9147 GND.n5327 GND.n5326 270.271
R9148 GND.n5327 GND.n1001 270.271
R9149 GND.n5335 GND.n1001 270.271
R9150 GND.n5336 GND.n5335 270.271
R9151 GND.n5337 GND.n5336 270.271
R9152 GND.n5337 GND.n995 270.271
R9153 GND.n5345 GND.n995 270.271
R9154 GND.n5346 GND.n5345 270.271
R9155 GND.n5347 GND.n5346 270.271
R9156 GND.n5347 GND.n989 270.271
R9157 GND.n5356 GND.n989 270.271
R9158 GND.n5357 GND.n5356 270.271
R9159 GND.n5358 GND.n5357 270.271
R9160 GND.n5358 GND.n984 270.271
R9161 GND.n3339 GND.t83 260.649
R9162 GND.n1959 GND.t108 260.649
R9163 GND.n3357 GND.n1734 256.663
R9164 GND.n3363 GND.n1734 256.663
R9165 GND.n3365 GND.n1734 256.663
R9166 GND.n3371 GND.n1734 256.663
R9167 GND.n3373 GND.n1734 256.663
R9168 GND.n3379 GND.n1734 256.663
R9169 GND.n3381 GND.n1734 256.663
R9170 GND.n3387 GND.n1734 256.663
R9171 GND.n3389 GND.n1734 256.663
R9172 GND.n3395 GND.n1734 256.663
R9173 GND.n3397 GND.n1734 256.663
R9174 GND.n3403 GND.n1734 256.663
R9175 GND.n3405 GND.n1734 256.663
R9176 GND.n3412 GND.n1734 256.663
R9177 GND.n3415 GND.n1734 256.663
R9178 GND.n3416 GND.n1554 256.663
R9179 GND.n3417 GND.n1734 256.663
R9180 GND.n3422 GND.n1734 256.663
R9181 GND.n3424 GND.n1734 256.663
R9182 GND.n3430 GND.n1734 256.663
R9183 GND.n3432 GND.n1734 256.663
R9184 GND.n3438 GND.n1734 256.663
R9185 GND.n3440 GND.n1734 256.663
R9186 GND.n3446 GND.n1734 256.663
R9187 GND.n3448 GND.n1734 256.663
R9188 GND.n3454 GND.n1734 256.663
R9189 GND.n3456 GND.n1734 256.663
R9190 GND.n3462 GND.n1734 256.663
R9191 GND.n3464 GND.n1734 256.663
R9192 GND.n3470 GND.n1734 256.663
R9193 GND.n3473 GND.n1734 256.663
R9194 GND.n4371 GND.n1970 256.663
R9195 GND.n4371 GND.n1971 256.663
R9196 GND.n4371 GND.n1972 256.663
R9197 GND.n4371 GND.n1973 256.663
R9198 GND.n4371 GND.n1974 256.663
R9199 GND.n4371 GND.n1975 256.663
R9200 GND.n4371 GND.n1976 256.663
R9201 GND.n4371 GND.n1977 256.663
R9202 GND.n4371 GND.n1978 256.663
R9203 GND.n4371 GND.n1979 256.663
R9204 GND.n4371 GND.n1980 256.663
R9205 GND.n4371 GND.n1981 256.663
R9206 GND.n4371 GND.n1982 256.663
R9207 GND.n4371 GND.n1983 256.663
R9208 GND.n4371 GND.n1984 256.663
R9209 GND.n4314 GND.n4313 256.663
R9210 GND.n4371 GND.n1985 256.663
R9211 GND.n4371 GND.n1986 256.663
R9212 GND.n4371 GND.n1987 256.663
R9213 GND.n4371 GND.n1988 256.663
R9214 GND.n4371 GND.n1989 256.663
R9215 GND.n4371 GND.n1990 256.663
R9216 GND.n4371 GND.n1991 256.663
R9217 GND.n4371 GND.n1992 256.663
R9218 GND.n4371 GND.n1993 256.663
R9219 GND.n4371 GND.n1994 256.663
R9220 GND.n4371 GND.n1995 256.663
R9221 GND.n4371 GND.n1996 256.663
R9222 GND.n4371 GND.n1997 256.663
R9223 GND.n4371 GND.n1998 256.663
R9224 GND.n4371 GND.n4370 256.663
R9225 GND.n4550 GND.n4549 242.672
R9226 GND.n4550 GND.n1649 242.672
R9227 GND.n4550 GND.n1651 242.672
R9228 GND.n4550 GND.n1652 242.672
R9229 GND.n4550 GND.n1654 242.672
R9230 GND.n4550 GND.n1656 242.672
R9231 GND.n4550 GND.n1657 242.672
R9232 GND.n4550 GND.n1659 242.672
R9233 GND.n4550 GND.n1660 242.672
R9234 GND.n4550 GND.n1661 242.672
R9235 GND.n4550 GND.n1662 242.672
R9236 GND.n4550 GND.n1663 242.672
R9237 GND.n4550 GND.n1664 242.672
R9238 GND.n3902 GND.n3882 242.672
R9239 GND.n3902 GND.n3883 242.672
R9240 GND.n3902 GND.n3885 242.672
R9241 GND.n3902 GND.n3886 242.672
R9242 GND.n3902 GND.n3888 242.672
R9243 GND.n3902 GND.n3889 242.672
R9244 GND.n3902 GND.n3891 242.672
R9245 GND.n3902 GND.n3893 242.672
R9246 GND.n3902 GND.n3894 242.672
R9247 GND.n3902 GND.n3896 242.672
R9248 GND.n3902 GND.n3898 242.672
R9249 GND.n3902 GND.n3899 242.672
R9250 GND.n3902 GND.n3901 242.672
R9251 GND.n4837 GND.n1366 242.672
R9252 GND.n4837 GND.n1367 242.672
R9253 GND.n4837 GND.n1368 242.672
R9254 GND.n4837 GND.n1369 242.672
R9255 GND.n4837 GND.n1370 242.672
R9256 GND.n4837 GND.n1371 242.672
R9257 GND.n4837 GND.n1372 242.672
R9258 GND.n4837 GND.n1373 242.672
R9259 GND.n4584 GND.n4583 242.672
R9260 GND.n4583 GND.n1638 242.672
R9261 GND.n4583 GND.n1637 242.672
R9262 GND.n4583 GND.n1635 242.672
R9263 GND.n4583 GND.n1633 242.672
R9264 GND.n4583 GND.n1632 242.672
R9265 GND.n4583 GND.n1630 242.672
R9266 GND.n4583 GND.n1628 242.672
R9267 GND.n4837 GND.n4836 242.672
R9268 GND.n4837 GND.n1350 242.672
R9269 GND.n4837 GND.n1351 242.672
R9270 GND.n4837 GND.n1352 242.672
R9271 GND.n4837 GND.n1353 242.672
R9272 GND.n4837 GND.n1354 242.672
R9273 GND.n4837 GND.n1355 242.672
R9274 GND.n4837 GND.n1356 242.672
R9275 GND.n4837 GND.n1357 242.672
R9276 GND.n4837 GND.n1358 242.672
R9277 GND.n4837 GND.n1359 242.672
R9278 GND.n4837 GND.n1360 242.672
R9279 GND.n4837 GND.n1361 242.672
R9280 GND.n4837 GND.n1362 242.672
R9281 GND.n4837 GND.n1363 242.672
R9282 GND.n4837 GND.n1364 242.672
R9283 GND.n4837 GND.n1365 242.672
R9284 GND.n4583 GND.n4559 242.672
R9285 GND.n4583 GND.n4560 242.672
R9286 GND.n4583 GND.n4562 242.672
R9287 GND.n4583 GND.n4563 242.672
R9288 GND.n4583 GND.n4565 242.672
R9289 GND.n4583 GND.n4566 242.672
R9290 GND.n4583 GND.n4568 242.672
R9291 GND.n4583 GND.n4569 242.672
R9292 GND.n4583 GND.n4571 242.672
R9293 GND.n4583 GND.n4572 242.672
R9294 GND.n4660 GND.n1553 242.672
R9295 GND.n4583 GND.n4573 242.672
R9296 GND.n4583 GND.n4575 242.672
R9297 GND.n4583 GND.n4576 242.672
R9298 GND.n4583 GND.n4578 242.672
R9299 GND.n4583 GND.n4579 242.672
R9300 GND.n4583 GND.n4581 242.672
R9301 GND.n4583 GND.n4582 242.672
R9302 GND.n4308 GND.n2012 242.672
R9303 GND.n4308 GND.n2013 242.672
R9304 GND.n4308 GND.n2014 242.672
R9305 GND.n4308 GND.n2015 242.672
R9306 GND.n4308 GND.n2016 242.672
R9307 GND.n4308 GND.n2017 242.672
R9308 GND.n4308 GND.n2018 242.672
R9309 GND.n4312 GND.n2004 242.672
R9310 GND.n4309 GND.n4308 242.672
R9311 GND.n4308 GND.n2021 242.672
R9312 GND.n4308 GND.n2022 242.672
R9313 GND.n4308 GND.n2023 242.672
R9314 GND.n4308 GND.n2024 242.672
R9315 GND.n4308 GND.n2025 242.672
R9316 GND.n4308 GND.n2026 242.672
R9317 GND.n4308 GND.n2027 242.672
R9318 GND.n4308 GND.n2028 242.672
R9319 GND.n4308 GND.n2029 242.672
R9320 GND.n5713 GND.n725 242.672
R9321 GND.n5713 GND.n726 242.672
R9322 GND.n5713 GND.n727 242.672
R9323 GND.n5713 GND.n728 242.672
R9324 GND.n5713 GND.n729 242.672
R9325 GND.n5713 GND.n730 242.672
R9326 GND.n5713 GND.n731 242.672
R9327 GND.n5713 GND.n732 242.672
R9328 GND.n5713 GND.n733 242.672
R9329 GND.n5713 GND.n734 242.672
R9330 GND.n5713 GND.n735 242.672
R9331 GND.n5713 GND.n736 242.672
R9332 GND.n5713 GND.n737 242.672
R9333 GND.n5713 GND.n738 242.672
R9334 GND.n5713 GND.n739 242.672
R9335 GND.n5713 GND.n740 242.672
R9336 GND.n5713 GND.n741 242.672
R9337 GND.n4308 GND.n2030 242.672
R9338 GND.n4308 GND.n2031 242.672
R9339 GND.n4308 GND.n2032 242.672
R9340 GND.n4308 GND.n2033 242.672
R9341 GND.n4308 GND.n2034 242.672
R9342 GND.n4308 GND.n2035 242.672
R9343 GND.n4308 GND.n2036 242.672
R9344 GND.n4308 GND.n2037 242.672
R9345 GND.n5713 GND.n723 242.672
R9346 GND.n5713 GND.n722 242.672
R9347 GND.n5713 GND.n721 242.672
R9348 GND.n5713 GND.n720 242.672
R9349 GND.n5713 GND.n719 242.672
R9350 GND.n5713 GND.n718 242.672
R9351 GND.n5713 GND.n717 242.672
R9352 GND.n5713 GND.n716 242.672
R9353 GND.n5712 GND.n743 240.244
R9354 GND.n748 GND.n747 240.244
R9355 GND.n750 GND.n749 240.244
R9356 GND.n754 GND.n753 240.244
R9357 GND.n756 GND.n755 240.244
R9358 GND.n760 GND.n759 240.244
R9359 GND.n762 GND.n761 240.244
R9360 GND.n766 GND.n765 240.244
R9361 GND.n770 GND.n769 240.244
R9362 GND.n774 GND.n773 240.244
R9363 GND.n776 GND.n775 240.244
R9364 GND.n780 GND.n779 240.244
R9365 GND.n782 GND.n781 240.244
R9366 GND.n786 GND.n785 240.244
R9367 GND.n788 GND.n787 240.244
R9368 GND.n792 GND.n791 240.244
R9369 GND.n796 GND.n793 240.244
R9370 GND.n2170 GND.n2169 240.244
R9371 GND.n2171 GND.n2170 240.244
R9372 GND.n2363 GND.n2171 240.244
R9373 GND.n2363 GND.n2177 240.244
R9374 GND.n2178 GND.n2177 240.244
R9375 GND.n2179 GND.n2178 240.244
R9376 GND.n4003 GND.n2179 240.244
R9377 GND.n4003 GND.n2185 240.244
R9378 GND.n2186 GND.n2185 240.244
R9379 GND.n2187 GND.n2186 240.244
R9380 GND.n2328 GND.n2187 240.244
R9381 GND.n2328 GND.n2193 240.244
R9382 GND.n2194 GND.n2193 240.244
R9383 GND.n2195 GND.n2194 240.244
R9384 GND.n2309 GND.n2195 240.244
R9385 GND.n2309 GND.n2201 240.244
R9386 GND.n2202 GND.n2201 240.244
R9387 GND.n2203 GND.n2202 240.244
R9388 GND.n2294 GND.n2203 240.244
R9389 GND.n2294 GND.n2209 240.244
R9390 GND.n2210 GND.n2209 240.244
R9391 GND.n2211 GND.n2210 240.244
R9392 GND.n2276 GND.n2211 240.244
R9393 GND.n2276 GND.n2217 240.244
R9394 GND.n2218 GND.n2217 240.244
R9395 GND.n2219 GND.n2218 240.244
R9396 GND.n4103 GND.n2219 240.244
R9397 GND.n4103 GND.n2225 240.244
R9398 GND.n2226 GND.n2225 240.244
R9399 GND.n2227 GND.n2226 240.244
R9400 GND.n4161 GND.n2227 240.244
R9401 GND.n4161 GND.n2233 240.244
R9402 GND.n2234 GND.n2233 240.244
R9403 GND.n2235 GND.n2234 240.244
R9404 GND.n2235 GND.n880 240.244
R9405 GND.n5537 GND.n880 240.244
R9406 GND.n5537 GND.n869 240.244
R9407 GND.n869 GND.n859 240.244
R9408 GND.n5553 GND.n859 240.244
R9409 GND.n5554 GND.n5553 240.244
R9410 GND.n5554 GND.n847 240.244
R9411 GND.n847 GND.n839 240.244
R9412 GND.n5570 GND.n839 240.244
R9413 GND.n5571 GND.n5570 240.244
R9414 GND.n5571 GND.n828 240.244
R9415 GND.n828 GND.n819 240.244
R9416 GND.n5587 GND.n819 240.244
R9417 GND.n5588 GND.n5587 240.244
R9418 GND.n5588 GND.n811 240.244
R9419 GND.n5590 GND.n811 240.244
R9420 GND.n5590 GND.n799 240.244
R9421 GND.n5656 GND.n799 240.244
R9422 GND.n2408 GND.n2407 240.244
R9423 GND.n2404 GND.n2403 240.244
R9424 GND.n2400 GND.n2399 240.244
R9425 GND.n2396 GND.n2395 240.244
R9426 GND.n2392 GND.n2391 240.244
R9427 GND.n2388 GND.n2387 240.244
R9428 GND.n2020 GND.n2019 240.244
R9429 GND.n4310 GND.n2010 240.244
R9430 GND.n2130 GND.n2129 240.244
R9431 GND.n2137 GND.n2136 240.244
R9432 GND.n2140 GND.n2139 240.244
R9433 GND.n2147 GND.n2146 240.244
R9434 GND.n2150 GND.n2149 240.244
R9435 GND.n2157 GND.n2156 240.244
R9436 GND.n2160 GND.n2159 240.244
R9437 GND.n2121 GND.n2116 240.244
R9438 GND.n3983 GND.n2412 240.244
R9439 GND.n3983 GND.n2366 240.244
R9440 GND.n3991 GND.n2366 240.244
R9441 GND.n3991 GND.n2368 240.244
R9442 GND.n2368 GND.n2349 240.244
R9443 GND.n4008 GND.n2349 240.244
R9444 GND.n4008 GND.n2343 240.244
R9445 GND.n4016 GND.n2343 240.244
R9446 GND.n4016 GND.n2345 240.244
R9447 GND.n2345 GND.n2326 240.244
R9448 GND.n4032 GND.n2326 240.244
R9449 GND.n4032 GND.n2320 240.244
R9450 GND.n4040 GND.n2320 240.244
R9451 GND.n4040 GND.n2322 240.244
R9452 GND.n2322 GND.n2303 240.244
R9453 GND.n4057 GND.n2303 240.244
R9454 GND.n4057 GND.n2293 240.244
R9455 GND.n4066 GND.n2293 240.244
R9456 GND.n4066 GND.n2299 240.244
R9457 GND.n2299 GND.n2270 240.244
R9458 GND.n4142 GND.n2270 240.244
R9459 GND.n4142 GND.n2271 240.244
R9460 GND.n4137 GND.n2271 240.244
R9461 GND.n4137 GND.n2274 240.244
R9462 GND.n4092 GND.n2274 240.244
R9463 GND.n4125 GND.n4092 240.244
R9464 GND.n4125 GND.n4093 240.244
R9465 GND.n4120 GND.n4093 240.244
R9466 GND.n4120 GND.n4101 240.244
R9467 GND.n4101 GND.n4100 240.244
R9468 GND.n4100 GND.n2246 240.244
R9469 GND.n4166 GND.n2246 240.244
R9470 GND.n4166 GND.n2241 240.244
R9471 GND.n4174 GND.n2241 240.244
R9472 GND.n4174 GND.n2242 240.244
R9473 GND.n2242 GND.n867 240.244
R9474 GND.n5545 GND.n867 240.244
R9475 GND.n5545 GND.n863 240.244
R9476 GND.n5551 GND.n863 240.244
R9477 GND.n5551 GND.n845 240.244
R9478 GND.n5562 GND.n845 240.244
R9479 GND.n5562 GND.n841 240.244
R9480 GND.n5568 GND.n841 240.244
R9481 GND.n5568 GND.n826 240.244
R9482 GND.n5579 GND.n826 240.244
R9483 GND.n5579 GND.n822 240.244
R9484 GND.n5585 GND.n822 240.244
R9485 GND.n5585 GND.n809 240.244
R9486 GND.n5597 GND.n809 240.244
R9487 GND.n5597 GND.n805 240.244
R9488 GND.n5604 GND.n805 240.244
R9489 GND.n5604 GND.n742 240.244
R9490 GND.n1534 GND.n1530 240.244
R9491 GND.n4580 GND.n1535 240.244
R9492 GND.n1539 GND.n1538 240.244
R9493 GND.n4577 GND.n1540 240.244
R9494 GND.n1544 GND.n1543 240.244
R9495 GND.n4574 GND.n1545 240.244
R9496 GND.n1549 GND.n1548 240.244
R9497 GND.n4570 GND.n1555 240.244
R9498 GND.n1559 GND.n1558 240.244
R9499 GND.n4567 GND.n1560 240.244
R9500 GND.n1564 GND.n1563 240.244
R9501 GND.n4564 GND.n1565 240.244
R9502 GND.n1569 GND.n1568 240.244
R9503 GND.n4561 GND.n1570 240.244
R9504 GND.n1574 GND.n1573 240.244
R9505 GND.n4558 GND.n1575 240.244
R9506 GND.n4766 GND.n1419 240.244
R9507 GND.n1425 GND.n1419 240.244
R9508 GND.n1426 GND.n1425 240.244
R9509 GND.n1427 GND.n1426 240.244
R9510 GND.n2803 GND.n1427 240.244
R9511 GND.n2803 GND.n1433 240.244
R9512 GND.n1434 GND.n1433 240.244
R9513 GND.n1435 GND.n1434 240.244
R9514 GND.n2800 GND.n1435 240.244
R9515 GND.n2800 GND.n1441 240.244
R9516 GND.n1442 GND.n1441 240.244
R9517 GND.n1443 GND.n1442 240.244
R9518 GND.n2940 GND.n1443 240.244
R9519 GND.n2940 GND.n1449 240.244
R9520 GND.n1450 GND.n1449 240.244
R9521 GND.n1451 GND.n1450 240.244
R9522 GND.n2750 GND.n1451 240.244
R9523 GND.n2750 GND.n1457 240.244
R9524 GND.n1458 GND.n1457 240.244
R9525 GND.n1459 GND.n1458 240.244
R9526 GND.n2729 GND.n1459 240.244
R9527 GND.n2729 GND.n1465 240.244
R9528 GND.n1466 GND.n1465 240.244
R9529 GND.n1467 GND.n1466 240.244
R9530 GND.n2698 GND.n1467 240.244
R9531 GND.n2698 GND.n1473 240.244
R9532 GND.n1474 GND.n1473 240.244
R9533 GND.n1475 GND.n1474 240.244
R9534 GND.n2722 GND.n1475 240.244
R9535 GND.n2722 GND.n1481 240.244
R9536 GND.n1482 GND.n1481 240.244
R9537 GND.n1483 GND.n1482 240.244
R9538 GND.n2669 GND.n1483 240.244
R9539 GND.n2669 GND.n1489 240.244
R9540 GND.n1490 GND.n1489 240.244
R9541 GND.n1491 GND.n1490 240.244
R9542 GND.n3060 GND.n1491 240.244
R9543 GND.n3060 GND.n1497 240.244
R9544 GND.n1498 GND.n1497 240.244
R9545 GND.n1499 GND.n1498 240.244
R9546 GND.n2637 GND.n1499 240.244
R9547 GND.n2637 GND.n1505 240.244
R9548 GND.n1506 GND.n1505 240.244
R9549 GND.n1507 GND.n1506 240.244
R9550 GND.n2618 GND.n1507 240.244
R9551 GND.n2618 GND.n1513 240.244
R9552 GND.n1514 GND.n1513 240.244
R9553 GND.n1515 GND.n1514 240.244
R9554 GND.n2610 GND.n1515 240.244
R9555 GND.n2610 GND.n1521 240.244
R9556 GND.n1522 GND.n1521 240.244
R9557 GND.n4686 GND.n1522 240.244
R9558 GND.n1377 GND.n1376 240.244
R9559 GND.n4830 GND.n1376 240.244
R9560 GND.n4828 GND.n4827 240.244
R9561 GND.n4824 GND.n4823 240.244
R9562 GND.n4820 GND.n4819 240.244
R9563 GND.n4816 GND.n4815 240.244
R9564 GND.n4812 GND.n4811 240.244
R9565 GND.n4808 GND.n4807 240.244
R9566 GND.n4803 GND.n4802 240.244
R9567 GND.n4799 GND.n4798 240.244
R9568 GND.n4795 GND.n4794 240.244
R9569 GND.n4791 GND.n4790 240.244
R9570 GND.n4787 GND.n4786 240.244
R9571 GND.n4783 GND.n4782 240.244
R9572 GND.n4779 GND.n4778 240.244
R9573 GND.n4775 GND.n4774 240.244
R9574 GND.n1414 GND.n1413 240.244
R9575 GND.n2902 GND.n1378 240.244
R9576 GND.n2909 GND.n2902 240.244
R9577 GND.n2909 GND.n2810 240.244
R9578 GND.n2916 GND.n2810 240.244
R9579 GND.n2916 GND.n2806 240.244
R9580 GND.n2922 GND.n2806 240.244
R9581 GND.n2922 GND.n2797 240.244
R9582 GND.n2929 GND.n2797 240.244
R9583 GND.n2929 GND.n2793 240.244
R9584 GND.n2935 GND.n2793 240.244
R9585 GND.n2935 GND.n2771 240.244
R9586 GND.n2945 GND.n2771 240.244
R9587 GND.n2945 GND.n2765 240.244
R9588 GND.n2953 GND.n2765 240.244
R9589 GND.n2953 GND.n2767 240.244
R9590 GND.n2767 GND.n2748 240.244
R9591 GND.n2982 GND.n2748 240.244
R9592 GND.n2982 GND.n2742 240.244
R9593 GND.n2989 GND.n2742 240.244
R9594 GND.n2989 GND.n2744 240.244
R9595 GND.n2744 GND.n2743 240.244
R9596 GND.n2743 GND.n2690 240.244
R9597 GND.n3102 GND.n2690 240.244
R9598 GND.n3102 GND.n2691 240.244
R9599 GND.n2714 GND.n2691 240.244
R9600 GND.n2715 GND.n2714 240.244
R9601 GND.n3087 GND.n2715 240.244
R9602 GND.n3087 GND.n3084 240.244
R9603 GND.n3084 GND.n2716 240.244
R9604 GND.n2716 GND.n2680 240.244
R9605 GND.n3110 GND.n2680 240.244
R9606 GND.n3110 GND.n2681 240.244
R9607 GND.n2681 GND.n2664 240.244
R9608 GND.n3127 GND.n2664 240.244
R9609 GND.n3127 GND.n2659 240.244
R9610 GND.n3135 GND.n2659 240.244
R9611 GND.n3135 GND.n2660 240.244
R9612 GND.n2660 GND.n2645 240.244
R9613 GND.n3152 GND.n2645 240.244
R9614 GND.n3152 GND.n2640 240.244
R9615 GND.n3160 GND.n2640 240.244
R9616 GND.n3160 GND.n2641 240.244
R9617 GND.n2641 GND.n2624 240.244
R9618 GND.n3178 GND.n2624 240.244
R9619 GND.n3178 GND.n2620 240.244
R9620 GND.n3184 GND.n2620 240.244
R9621 GND.n3184 GND.n2598 240.244
R9622 GND.n3218 GND.n2598 240.244
R9623 GND.n3218 GND.n2594 240.244
R9624 GND.n3224 GND.n2594 240.244
R9625 GND.n3224 GND.n1529 240.244
R9626 GND.n4684 GND.n1529 240.244
R9627 GND.n1582 GND.n1581 240.244
R9628 GND.n1629 GND.n1583 240.244
R9629 GND.n1593 GND.n1592 240.244
R9630 GND.n1631 GND.n1600 240.244
R9631 GND.n1634 GND.n1601 240.244
R9632 GND.n1609 GND.n1608 240.244
R9633 GND.n1636 GND.n1616 240.244
R9634 GND.n1626 GND.n1617 240.244
R9635 GND.n2872 GND.n2815 240.244
R9636 GND.n2901 GND.n2815 240.244
R9637 GND.n2901 GND.n2816 240.244
R9638 GND.n2816 GND.n2812 240.244
R9639 GND.n2877 GND.n2812 240.244
R9640 GND.n2877 GND.n2805 240.244
R9641 GND.n2878 GND.n2805 240.244
R9642 GND.n2878 GND.n2799 240.244
R9643 GND.n2881 GND.n2799 240.244
R9644 GND.n2881 GND.n2792 240.244
R9645 GND.n2882 GND.n2792 240.244
R9646 GND.n2882 GND.n2773 240.244
R9647 GND.n2773 GND.n2761 240.244
R9648 GND.n2955 GND.n2761 240.244
R9649 GND.n2955 GND.n2756 240.244
R9650 GND.n2976 GND.n2756 240.244
R9651 GND.n2976 GND.n2751 240.244
R9652 GND.n2960 GND.n2751 240.244
R9653 GND.n2960 GND.n2739 240.244
R9654 GND.n2966 GND.n2739 240.244
R9655 GND.n2966 GND.n2728 240.244
R9656 GND.n3005 GND.n2728 240.244
R9657 GND.n3005 GND.n2693 240.244
R9658 GND.n2697 GND.n2693 240.244
R9659 GND.n3012 GND.n2697 240.244
R9660 GND.n3013 GND.n3012 240.244
R9661 GND.n3013 GND.n2707 240.244
R9662 GND.n2719 GND.n2707 240.244
R9663 GND.n3020 GND.n2719 240.244
R9664 GND.n3020 GND.n2675 240.244
R9665 GND.n3112 GND.n2675 240.244
R9666 GND.n3112 GND.n2670 240.244
R9667 GND.n3119 GND.n2670 240.244
R9668 GND.n3119 GND.n2666 240.244
R9669 GND.n2666 GND.n2655 240.244
R9670 GND.n3137 GND.n2655 240.244
R9671 GND.n3137 GND.n2650 240.244
R9672 GND.n3144 GND.n2650 240.244
R9673 GND.n3144 GND.n2647 240.244
R9674 GND.n2647 GND.n2635 240.244
R9675 GND.n3162 GND.n2635 240.244
R9676 GND.n3162 GND.n2630 240.244
R9677 GND.n3172 GND.n2630 240.244
R9678 GND.n3172 GND.n2626 240.244
R9679 GND.n3166 GND.n2626 240.244
R9680 GND.n3166 GND.n2605 240.244
R9681 GND.n3213 GND.n2605 240.244
R9682 GND.n3213 GND.n2600 240.244
R9683 GND.n3207 GND.n2600 240.244
R9684 GND.n3207 GND.n2591 240.244
R9685 GND.n3231 GND.n2591 240.244
R9686 GND.n3231 GND.n1526 240.244
R9687 GND.n2837 GND.n2836 240.244
R9688 GND.n2847 GND.n2846 240.244
R9689 GND.n2833 GND.n2832 240.244
R9690 GND.n2855 GND.n2854 240.244
R9691 GND.n2829 GND.n2828 240.244
R9692 GND.n2863 GND.n2862 240.244
R9693 GND.n2825 GND.n2824 240.244
R9694 GND.n2820 GND.n1374 240.244
R9695 GND.n2838 GND.n2813 240.244
R9696 GND.n2911 GND.n2813 240.244
R9697 GND.n2913 GND.n2911 240.244
R9698 GND.n2914 GND.n2913 240.244
R9699 GND.n2914 GND.n2802 240.244
R9700 GND.n2924 GND.n2802 240.244
R9701 GND.n2926 GND.n2924 240.244
R9702 GND.n2927 GND.n2926 240.244
R9703 GND.n2927 GND.n2791 240.244
R9704 GND.n2937 GND.n2791 240.244
R9705 GND.n2939 GND.n2937 240.244
R9706 GND.n2943 GND.n2939 240.244
R9707 GND.n2943 GND.n2942 240.244
R9708 GND.n2942 GND.n2764 240.244
R9709 GND.n2764 GND.n2754 240.244
R9710 GND.n2978 GND.n2754 240.244
R9711 GND.n2980 GND.n2978 240.244
R9712 GND.n2980 GND.n2979 240.244
R9713 GND.n2979 GND.n2741 240.244
R9714 GND.n2964 GND.n2741 240.244
R9715 GND.n2964 GND.n2963 240.244
R9716 GND.n2963 GND.n2695 240.244
R9717 GND.n3100 GND.n2695 240.244
R9718 GND.n3100 GND.n3098 240.244
R9719 GND.n3098 GND.n2696 240.244
R9720 GND.n2709 GND.n2696 240.244
R9721 GND.n2711 GND.n2709 240.244
R9722 GND.n3082 GND.n2711 240.244
R9723 GND.n3082 GND.n3081 240.244
R9724 GND.n3081 GND.n2721 240.244
R9725 GND.n2721 GND.n2679 240.244
R9726 GND.n2679 GND.n2668 240.244
R9727 GND.n3121 GND.n2668 240.244
R9728 GND.n3125 GND.n3121 240.244
R9729 GND.n3125 GND.n3124 240.244
R9730 GND.n3124 GND.n2658 240.244
R9731 GND.n2658 GND.n2649 240.244
R9732 GND.n3146 GND.n2649 240.244
R9733 GND.n3150 GND.n3146 240.244
R9734 GND.n3150 GND.n3148 240.244
R9735 GND.n3148 GND.n2639 240.244
R9736 GND.n2639 GND.n2628 240.244
R9737 GND.n3174 GND.n2628 240.244
R9738 GND.n3176 GND.n3174 240.244
R9739 GND.n3176 GND.n3175 240.244
R9740 GND.n3175 GND.n2602 240.244
R9741 GND.n3215 GND.n2602 240.244
R9742 GND.n3216 GND.n3215 240.244
R9743 GND.n3216 GND.n2593 240.244
R9744 GND.n3226 GND.n2593 240.244
R9745 GND.n3229 GND.n3226 240.244
R9746 GND.n3229 GND.n1528 240.244
R9747 GND.n2045 GND.n2044 240.244
R9748 GND.n3900 GND.n2054 240.244
R9749 GND.n3897 GND.n2055 240.244
R9750 GND.n2063 GND.n2062 240.244
R9751 GND.n3895 GND.n2072 240.244
R9752 GND.n3892 GND.n2073 240.244
R9753 GND.n2081 GND.n2080 240.244
R9754 GND.n3890 GND.n2086 240.244
R9755 GND.n2088 GND.n2087 240.244
R9756 GND.n3887 GND.n2092 240.244
R9757 GND.n2094 GND.n2093 240.244
R9758 GND.n3884 GND.n2100 240.244
R9759 GND.n2102 GND.n2101 240.244
R9760 GND.n3270 GND.n1669 240.244
R9761 GND.n3273 GND.n3270 240.244
R9762 GND.n3273 GND.n1681 240.244
R9763 GND.n2582 GND.n1681 240.244
R9764 GND.n2582 GND.n1695 240.244
R9765 GND.n3281 GND.n1695 240.244
R9766 GND.n3281 GND.n3280 240.244
R9767 GND.n3280 GND.n1709 240.244
R9768 GND.n3288 GND.n1709 240.244
R9769 GND.n3288 GND.n1722 240.244
R9770 GND.n2573 GND.n1722 240.244
R9771 GND.n2576 GND.n2573 240.244
R9772 GND.n2576 GND.n1735 240.244
R9773 GND.n3481 GND.n1735 240.244
R9774 GND.n3481 GND.n1747 240.244
R9775 GND.n3487 GND.n1747 240.244
R9776 GND.n3487 GND.n1757 240.244
R9777 GND.n3514 GND.n1757 240.244
R9778 GND.n3514 GND.n1767 240.244
R9779 GND.n3505 GND.n1767 240.244
R9780 GND.n3505 GND.n1777 240.244
R9781 GND.n2539 GND.n1777 240.244
R9782 GND.n2539 GND.n1787 240.244
R9783 GND.n3550 GND.n1787 240.244
R9784 GND.n3550 GND.n1797 240.244
R9785 GND.n3567 GND.n1797 240.244
R9786 GND.n3567 GND.n1807 240.244
R9787 GND.n2528 GND.n1807 240.244
R9788 GND.n2528 GND.n1816 240.244
R9789 GND.n3558 GND.n1816 240.244
R9790 GND.n3558 GND.n1825 240.244
R9791 GND.n3613 GND.n1825 240.244
R9792 GND.n3613 GND.n1835 240.244
R9793 GND.n3621 GND.n1835 240.244
R9794 GND.n3621 GND.n1844 240.244
R9795 GND.n3648 GND.n1844 240.244
R9796 GND.n3649 GND.n3648 240.244
R9797 GND.n3650 GND.n3649 240.244
R9798 GND.n3650 GND.n1864 240.244
R9799 GND.n3660 GND.n1864 240.244
R9800 GND.n3660 GND.n1881 240.244
R9801 GND.n3654 GND.n1881 240.244
R9802 GND.n3654 GND.n2488 240.244
R9803 GND.n3686 GND.n2488 240.244
R9804 GND.n3686 GND.n1907 240.244
R9805 GND.n3705 GND.n1907 240.244
R9806 GND.n3705 GND.n1918 240.244
R9807 GND.n3691 GND.n1918 240.244
R9808 GND.n3692 GND.n3691 240.244
R9809 GND.n3693 GND.n3692 240.244
R9810 GND.n3694 GND.n3693 240.244
R9811 GND.n3694 GND.n2477 240.244
R9812 GND.n3807 GND.n2477 240.244
R9813 GND.n3807 GND.n2472 240.244
R9814 GND.n3814 GND.n2472 240.244
R9815 GND.n3814 GND.n2459 240.244
R9816 GND.n2459 GND.n2450 240.244
R9817 GND.n3839 GND.n2450 240.244
R9818 GND.n3839 GND.n2445 240.244
R9819 GND.n3851 GND.n2445 240.244
R9820 GND.n3851 GND.n2436 240.244
R9821 GND.n3844 GND.n2436 240.244
R9822 GND.n3844 GND.n2429 240.244
R9823 GND.n2429 GND.n2106 240.244
R9824 GND.n4239 GND.n2106 240.244
R9825 GND.n1589 GND.n1588 240.244
R9826 GND.n1648 GND.n1589 240.244
R9827 GND.n1597 GND.n1596 240.244
R9828 GND.n1650 GND.n1604 240.244
R9829 GND.n1653 GND.n1605 240.244
R9830 GND.n1613 GND.n1612 240.244
R9831 GND.n1655 GND.n1622 240.244
R9832 GND.n1658 GND.n1623 240.244
R9833 GND.n3239 GND.n3238 240.244
R9834 GND.n3242 GND.n3241 240.244
R9835 GND.n3249 GND.n3248 240.244
R9836 GND.n3252 GND.n3251 240.244
R9837 GND.n3262 GND.n3261 240.244
R9838 GND.n4547 GND.n1666 240.244
R9839 GND.n1683 GND.n1666 240.244
R9840 GND.n4537 GND.n1683 240.244
R9841 GND.n4537 GND.n1684 240.244
R9842 GND.n4533 GND.n1684 240.244
R9843 GND.n4533 GND.n1693 240.244
R9844 GND.n1711 GND.n1693 240.244
R9845 GND.n4523 GND.n1711 240.244
R9846 GND.n4523 GND.n1712 240.244
R9847 GND.n4519 GND.n1712 240.244
R9848 GND.n4519 GND.n1720 240.244
R9849 GND.n1736 GND.n1720 240.244
R9850 GND.n4509 GND.n1736 240.244
R9851 GND.n4509 GND.n1737 240.244
R9852 GND.n4505 GND.n1737 240.244
R9853 GND.n4505 GND.n1745 240.244
R9854 GND.n4495 GND.n1745 240.244
R9855 GND.n4495 GND.n1759 240.244
R9856 GND.n4491 GND.n1759 240.244
R9857 GND.n4491 GND.n1765 240.244
R9858 GND.n4481 GND.n1765 240.244
R9859 GND.n4481 GND.n1779 240.244
R9860 GND.n4477 GND.n1779 240.244
R9861 GND.n4477 GND.n1785 240.244
R9862 GND.n4467 GND.n1785 240.244
R9863 GND.n4467 GND.n1799 240.244
R9864 GND.n4463 GND.n1799 240.244
R9865 GND.n4463 GND.n1805 240.244
R9866 GND.n4453 GND.n1805 240.244
R9867 GND.n4453 GND.n1817 240.244
R9868 GND.n4449 GND.n1817 240.244
R9869 GND.n4449 GND.n1823 240.244
R9870 GND.n4439 GND.n1823 240.244
R9871 GND.n4439 GND.n1837 240.244
R9872 GND.n4435 GND.n1837 240.244
R9873 GND.n4435 GND.n1843 240.244
R9874 GND.n1870 GND.n1843 240.244
R9875 GND.n1870 GND.n1866 240.244
R9876 GND.n4418 GND.n1866 240.244
R9877 GND.n4418 GND.n1867 240.244
R9878 GND.n4414 GND.n1867 240.244
R9879 GND.n4414 GND.n1878 240.244
R9880 GND.n2494 GND.n1878 240.244
R9881 GND.n2494 GND.n1909 240.244
R9882 GND.n4398 GND.n1909 240.244
R9883 GND.n4398 GND.n1910 240.244
R9884 GND.n4394 GND.n1910 240.244
R9885 GND.n4394 GND.n1916 240.244
R9886 GND.n3795 GND.n1916 240.244
R9887 GND.n3796 GND.n3795 240.244
R9888 GND.n3797 GND.n3796 240.244
R9889 GND.n3797 GND.n3787 240.244
R9890 GND.n3805 GND.n3787 240.244
R9891 GND.n3805 GND.n3788 240.244
R9892 GND.n3788 GND.n2458 240.244
R9893 GND.n3829 GND.n2458 240.244
R9894 GND.n3829 GND.n2453 240.244
R9895 GND.n3837 GND.n2453 240.244
R9896 GND.n3837 GND.n2454 240.244
R9897 GND.n2454 GND.n2434 240.244
R9898 GND.n3863 GND.n2434 240.244
R9899 GND.n3863 GND.n2430 240.244
R9900 GND.n3869 GND.n2430 240.244
R9901 GND.n3869 GND.n2110 240.244
R9902 GND.n4237 GND.n2110 240.244
R9903 GND.n4968 GND.n1222 240.244
R9904 GND.n4968 GND.n1218 240.244
R9905 GND.n4974 GND.n1218 240.244
R9906 GND.n4974 GND.n1216 240.244
R9907 GND.n4978 GND.n1216 240.244
R9908 GND.n4978 GND.n1212 240.244
R9909 GND.n4984 GND.n1212 240.244
R9910 GND.n4984 GND.n1210 240.244
R9911 GND.n4988 GND.n1210 240.244
R9912 GND.n4988 GND.n1206 240.244
R9913 GND.n4994 GND.n1206 240.244
R9914 GND.n4994 GND.n1204 240.244
R9915 GND.n4998 GND.n1204 240.244
R9916 GND.n4998 GND.n1200 240.244
R9917 GND.n5004 GND.n1200 240.244
R9918 GND.n5004 GND.n1198 240.244
R9919 GND.n5008 GND.n1198 240.244
R9920 GND.n5008 GND.n1194 240.244
R9921 GND.n5014 GND.n1194 240.244
R9922 GND.n5014 GND.n1192 240.244
R9923 GND.n5018 GND.n1192 240.244
R9924 GND.n5018 GND.n1188 240.244
R9925 GND.n5024 GND.n1188 240.244
R9926 GND.n5024 GND.n1186 240.244
R9927 GND.n5028 GND.n1186 240.244
R9928 GND.n5028 GND.n1182 240.244
R9929 GND.n5034 GND.n1182 240.244
R9930 GND.n5034 GND.n1180 240.244
R9931 GND.n5038 GND.n1180 240.244
R9932 GND.n5038 GND.n1176 240.244
R9933 GND.n5044 GND.n1176 240.244
R9934 GND.n5044 GND.n1174 240.244
R9935 GND.n5048 GND.n1174 240.244
R9936 GND.n5048 GND.n1170 240.244
R9937 GND.n5054 GND.n1170 240.244
R9938 GND.n5054 GND.n1168 240.244
R9939 GND.n5058 GND.n1168 240.244
R9940 GND.n5058 GND.n1164 240.244
R9941 GND.n5064 GND.n1164 240.244
R9942 GND.n5064 GND.n1162 240.244
R9943 GND.n5068 GND.n1162 240.244
R9944 GND.n5068 GND.n1158 240.244
R9945 GND.n5074 GND.n1158 240.244
R9946 GND.n5074 GND.n1156 240.244
R9947 GND.n5078 GND.n1156 240.244
R9948 GND.n5078 GND.n1152 240.244
R9949 GND.n5084 GND.n1152 240.244
R9950 GND.n5084 GND.n1150 240.244
R9951 GND.n5088 GND.n1150 240.244
R9952 GND.n5088 GND.n1146 240.244
R9953 GND.n5094 GND.n1146 240.244
R9954 GND.n5094 GND.n1144 240.244
R9955 GND.n5098 GND.n1144 240.244
R9956 GND.n5098 GND.n1140 240.244
R9957 GND.n5104 GND.n1140 240.244
R9958 GND.n5104 GND.n1138 240.244
R9959 GND.n5108 GND.n1138 240.244
R9960 GND.n5108 GND.n1134 240.244
R9961 GND.n5114 GND.n1134 240.244
R9962 GND.n5114 GND.n1132 240.244
R9963 GND.n5118 GND.n1132 240.244
R9964 GND.n5118 GND.n1128 240.244
R9965 GND.n5124 GND.n1128 240.244
R9966 GND.n5124 GND.n1126 240.244
R9967 GND.n5128 GND.n1126 240.244
R9968 GND.n5128 GND.n1122 240.244
R9969 GND.n5134 GND.n1122 240.244
R9970 GND.n5134 GND.n1120 240.244
R9971 GND.n5138 GND.n1120 240.244
R9972 GND.n5138 GND.n1116 240.244
R9973 GND.n5144 GND.n1116 240.244
R9974 GND.n5144 GND.n1114 240.244
R9975 GND.n5148 GND.n1114 240.244
R9976 GND.n5148 GND.n1110 240.244
R9977 GND.n5154 GND.n1110 240.244
R9978 GND.n5154 GND.n1108 240.244
R9979 GND.n5158 GND.n1108 240.244
R9980 GND.n5158 GND.n1104 240.244
R9981 GND.n5164 GND.n1104 240.244
R9982 GND.n5164 GND.n1102 240.244
R9983 GND.n5168 GND.n1102 240.244
R9984 GND.n5168 GND.n1098 240.244
R9985 GND.n5174 GND.n1098 240.244
R9986 GND.n5174 GND.n1096 240.244
R9987 GND.n5178 GND.n1096 240.244
R9988 GND.n5178 GND.n1092 240.244
R9989 GND.n5184 GND.n1092 240.244
R9990 GND.n5184 GND.n1090 240.244
R9991 GND.n5188 GND.n1090 240.244
R9992 GND.n5188 GND.n1086 240.244
R9993 GND.n5194 GND.n1086 240.244
R9994 GND.n5194 GND.n1084 240.244
R9995 GND.n5198 GND.n1084 240.244
R9996 GND.n5198 GND.n1080 240.244
R9997 GND.n5204 GND.n1080 240.244
R9998 GND.n5204 GND.n1078 240.244
R9999 GND.n5208 GND.n1078 240.244
R10000 GND.n5208 GND.n1074 240.244
R10001 GND.n5214 GND.n1074 240.244
R10002 GND.n5214 GND.n1072 240.244
R10003 GND.n5218 GND.n1072 240.244
R10004 GND.n5218 GND.n1068 240.244
R10005 GND.n5224 GND.n1068 240.244
R10006 GND.n5224 GND.n1066 240.244
R10007 GND.n5228 GND.n1066 240.244
R10008 GND.n5228 GND.n1062 240.244
R10009 GND.n5234 GND.n1062 240.244
R10010 GND.n5234 GND.n1060 240.244
R10011 GND.n5238 GND.n1060 240.244
R10012 GND.n5238 GND.n1056 240.244
R10013 GND.n5244 GND.n1056 240.244
R10014 GND.n5244 GND.n1054 240.244
R10015 GND.n5248 GND.n1054 240.244
R10016 GND.n5248 GND.n1050 240.244
R10017 GND.n5254 GND.n1050 240.244
R10018 GND.n5254 GND.n1048 240.244
R10019 GND.n5258 GND.n1048 240.244
R10020 GND.n5258 GND.n1044 240.244
R10021 GND.n5264 GND.n1044 240.244
R10022 GND.n5264 GND.n1042 240.244
R10023 GND.n5268 GND.n1042 240.244
R10024 GND.n5268 GND.n1038 240.244
R10025 GND.n5274 GND.n1038 240.244
R10026 GND.n5274 GND.n1036 240.244
R10027 GND.n5278 GND.n1036 240.244
R10028 GND.n5278 GND.n1032 240.244
R10029 GND.n5284 GND.n1032 240.244
R10030 GND.n5284 GND.n1030 240.244
R10031 GND.n5288 GND.n1030 240.244
R10032 GND.n5288 GND.n1026 240.244
R10033 GND.n5294 GND.n1026 240.244
R10034 GND.n5294 GND.n1024 240.244
R10035 GND.n5298 GND.n1024 240.244
R10036 GND.n5298 GND.n1020 240.244
R10037 GND.n5304 GND.n1020 240.244
R10038 GND.n5304 GND.n1018 240.244
R10039 GND.n5308 GND.n1018 240.244
R10040 GND.n5308 GND.n1014 240.244
R10041 GND.n5314 GND.n1014 240.244
R10042 GND.n5314 GND.n1012 240.244
R10043 GND.n5318 GND.n1012 240.244
R10044 GND.n5318 GND.n1008 240.244
R10045 GND.n5324 GND.n1008 240.244
R10046 GND.n5324 GND.n1006 240.244
R10047 GND.n5328 GND.n1006 240.244
R10048 GND.n5328 GND.n1002 240.244
R10049 GND.n5334 GND.n1002 240.244
R10050 GND.n5334 GND.n1000 240.244
R10051 GND.n5338 GND.n1000 240.244
R10052 GND.n5338 GND.n996 240.244
R10053 GND.n5344 GND.n996 240.244
R10054 GND.n5344 GND.n994 240.244
R10055 GND.n5348 GND.n994 240.244
R10056 GND.n5348 GND.n990 240.244
R10057 GND.n5355 GND.n990 240.244
R10058 GND.n5355 GND.n988 240.244
R10059 GND.n5359 GND.n988 240.244
R10060 GND.n5359 GND.n985 240.244
R10061 GND.n5365 GND.n983 240.244
R10062 GND.n5369 GND.n983 240.244
R10063 GND.n5369 GND.n979 240.244
R10064 GND.n5375 GND.n979 240.244
R10065 GND.n5375 GND.n977 240.244
R10066 GND.n5379 GND.n977 240.244
R10067 GND.n5379 GND.n973 240.244
R10068 GND.n5385 GND.n973 240.244
R10069 GND.n5385 GND.n971 240.244
R10070 GND.n5389 GND.n971 240.244
R10071 GND.n5389 GND.n967 240.244
R10072 GND.n5395 GND.n967 240.244
R10073 GND.n5395 GND.n965 240.244
R10074 GND.n5399 GND.n965 240.244
R10075 GND.n5399 GND.n961 240.244
R10076 GND.n5405 GND.n961 240.244
R10077 GND.n5405 GND.n959 240.244
R10078 GND.n5409 GND.n959 240.244
R10079 GND.n5409 GND.n955 240.244
R10080 GND.n5415 GND.n955 240.244
R10081 GND.n5415 GND.n953 240.244
R10082 GND.n5419 GND.n953 240.244
R10083 GND.n5419 GND.n949 240.244
R10084 GND.n5425 GND.n949 240.244
R10085 GND.n5425 GND.n947 240.244
R10086 GND.n5429 GND.n947 240.244
R10087 GND.n5429 GND.n943 240.244
R10088 GND.n5435 GND.n943 240.244
R10089 GND.n5435 GND.n941 240.244
R10090 GND.n5439 GND.n941 240.244
R10091 GND.n5439 GND.n937 240.244
R10092 GND.n5445 GND.n937 240.244
R10093 GND.n5445 GND.n935 240.244
R10094 GND.n5449 GND.n935 240.244
R10095 GND.n5449 GND.n931 240.244
R10096 GND.n5455 GND.n931 240.244
R10097 GND.n5455 GND.n929 240.244
R10098 GND.n5459 GND.n929 240.244
R10099 GND.n5459 GND.n925 240.244
R10100 GND.n5465 GND.n925 240.244
R10101 GND.n5465 GND.n923 240.244
R10102 GND.n5469 GND.n923 240.244
R10103 GND.n5469 GND.n919 240.244
R10104 GND.n5475 GND.n919 240.244
R10105 GND.n5475 GND.n917 240.244
R10106 GND.n5479 GND.n917 240.244
R10107 GND.n5479 GND.n913 240.244
R10108 GND.n5485 GND.n913 240.244
R10109 GND.n5485 GND.n911 240.244
R10110 GND.n5489 GND.n911 240.244
R10111 GND.n5489 GND.n907 240.244
R10112 GND.n5495 GND.n907 240.244
R10113 GND.n5495 GND.n905 240.244
R10114 GND.n5499 GND.n905 240.244
R10115 GND.n5499 GND.n901 240.244
R10116 GND.n5505 GND.n901 240.244
R10117 GND.n5505 GND.n899 240.244
R10118 GND.n5509 GND.n899 240.244
R10119 GND.n5509 GND.n895 240.244
R10120 GND.n5516 GND.n895 240.244
R10121 GND.n5516 GND.n893 240.244
R10122 GND.n5520 GND.n893 240.244
R10123 GND.n5520 GND.n889 240.244
R10124 GND.n2789 GND.n2774 240.244
R10125 GND.n2785 GND.n2774 240.244
R10126 GND.n2785 GND.n2784 240.244
R10127 GND.n2784 GND.n2783 240.244
R10128 GND.n2783 GND.n2736 240.244
R10129 GND.n2992 GND.n2736 240.244
R10130 GND.n2992 GND.n2737 240.244
R10131 GND.n2737 GND.n2731 240.244
R10132 GND.n3002 GND.n2731 240.244
R10133 GND.n3002 GND.n2732 240.244
R10134 GND.n2732 GND.n2700 240.244
R10135 GND.n3095 GND.n2700 240.244
R10136 GND.n3095 GND.n2701 240.244
R10137 GND.n3090 GND.n2701 240.244
R10138 GND.n3090 GND.n2704 240.244
R10139 GND.n3022 GND.n2704 240.244
R10140 GND.n3078 GND.n3022 240.244
R10141 GND.n3078 GND.n3023 240.244
R10142 GND.n3073 GND.n3023 240.244
R10143 GND.n3073 GND.n3072 240.244
R10144 GND.n3072 GND.n3069 240.244
R10145 GND.n3069 GND.n3028 240.244
R10146 GND.n3065 GND.n3028 240.244
R10147 GND.n3065 GND.n3064 240.244
R10148 GND.n3064 GND.n3063 240.244
R10149 GND.n3063 GND.n3034 240.244
R10150 GND.n3056 GND.n3034 240.244
R10151 GND.n3056 GND.n3055 240.244
R10152 GND.n3055 GND.n3054 240.244
R10153 GND.n3054 GND.n3042 240.244
R10154 GND.n3050 GND.n3042 240.244
R10155 GND.n3050 GND.n2616 240.244
R10156 GND.n3187 GND.n2616 240.244
R10157 GND.n3188 GND.n3187 240.244
R10158 GND.n3189 GND.n3188 240.244
R10159 GND.n3189 GND.n2611 240.244
R10160 GND.n3204 GND.n2611 240.244
R10161 GND.n3204 GND.n2612 240.244
R10162 GND.n3200 GND.n2612 240.244
R10163 GND.n3200 GND.n3199 240.244
R10164 GND.n3199 GND.n1640 240.244
R10165 GND.n4556 GND.n1640 240.244
R10166 GND.n4556 GND.n1641 240.244
R10167 GND.n4552 GND.n1641 240.244
R10168 GND.n4552 GND.n1647 240.244
R10169 GND.n1671 GND.n1647 240.244
R10170 GND.n4544 GND.n1671 240.244
R10171 GND.n4544 GND.n1672 240.244
R10172 GND.n4540 GND.n1672 240.244
R10173 GND.n4540 GND.n1680 240.244
R10174 GND.n1697 GND.n1680 240.244
R10175 GND.n4530 GND.n1697 240.244
R10176 GND.n4530 GND.n1698 240.244
R10177 GND.n4526 GND.n1698 240.244
R10178 GND.n4526 GND.n1706 240.244
R10179 GND.n1724 GND.n1706 240.244
R10180 GND.n4516 GND.n1724 240.244
R10181 GND.n4516 GND.n1725 240.244
R10182 GND.n4512 GND.n1725 240.244
R10183 GND.n4512 GND.n1733 240.244
R10184 GND.n2552 GND.n1733 240.244
R10185 GND.n2553 GND.n2552 240.244
R10186 GND.n2554 GND.n2553 240.244
R10187 GND.n2554 GND.n2545 240.244
R10188 GND.n3517 GND.n2545 240.244
R10189 GND.n3518 GND.n3517 240.244
R10190 GND.n3519 GND.n3518 240.244
R10191 GND.n3519 GND.n2540 240.244
R10192 GND.n3535 GND.n2540 240.244
R10193 GND.n3535 GND.n2541 240.244
R10194 GND.n3531 GND.n2541 240.244
R10195 GND.n3531 GND.n3530 240.244
R10196 GND.n3530 GND.n2527 240.244
R10197 GND.n3584 GND.n2527 240.244
R10198 GND.n3585 GND.n3584 240.244
R10199 GND.n3585 GND.n2522 240.244
R10200 GND.n3600 GND.n2522 240.244
R10201 GND.n3600 GND.n2523 240.244
R10202 GND.n3596 GND.n2523 240.244
R10203 GND.n3596 GND.n3595 240.244
R10204 GND.n3595 GND.n1846 240.244
R10205 GND.n4432 GND.n1846 240.244
R10206 GND.n4432 GND.n1847 240.244
R10207 GND.n4428 GND.n1847 240.244
R10208 GND.n4428 GND.n1853 240.244
R10209 GND.n1896 GND.n1853 240.244
R10210 GND.n1897 GND.n1896 240.244
R10211 GND.n1897 GND.n1890 240.244
R10212 GND.n4405 GND.n1890 240.244
R10213 GND.n4405 GND.n1891 240.244
R10214 GND.n4401 GND.n1891 240.244
R10215 GND.n4401 GND.n1905 240.244
R10216 GND.n1933 GND.n1905 240.244
R10217 GND.n1933 GND.n1929 240.244
R10218 GND.n4384 GND.n1929 240.244
R10219 GND.n4384 GND.n1930 240.244
R10220 GND.n4380 GND.n1930 240.244
R10221 GND.n4380 GND.n1941 240.244
R10222 GND.n2469 GND.n1941 240.244
R10223 GND.n2470 GND.n2469 240.244
R10224 GND.n3818 GND.n2470 240.244
R10225 GND.n3818 GND.n2461 240.244
R10226 GND.n3826 GND.n2461 240.244
R10227 GND.n3826 GND.n2462 240.244
R10228 GND.n2462 GND.n2443 240.244
R10229 GND.n3854 GND.n2443 240.244
R10230 GND.n3854 GND.n2439 240.244
R10231 GND.n3860 GND.n2439 240.244
R10232 GND.n3860 GND.n2428 240.244
R10233 GND.n3873 GND.n2428 240.244
R10234 GND.n3873 GND.n2424 240.244
R10235 GND.n3879 GND.n2424 240.244
R10236 GND.n3880 GND.n3879 240.244
R10237 GND.n3905 GND.n3880 240.244
R10238 GND.n3905 GND.n2420 240.244
R10239 GND.n3911 GND.n2420 240.244
R10240 GND.n3912 GND.n3911 240.244
R10241 GND.n3920 GND.n3912 240.244
R10242 GND.n3920 GND.n2415 240.244
R10243 GND.n3976 GND.n2415 240.244
R10244 GND.n3976 GND.n2416 240.244
R10245 GND.n3972 GND.n2416 240.244
R10246 GND.n3972 GND.n3971 240.244
R10247 GND.n3971 GND.n3970 240.244
R10248 GND.n3970 GND.n3928 240.244
R10249 GND.n3966 GND.n3928 240.244
R10250 GND.n3966 GND.n3965 240.244
R10251 GND.n3965 GND.n3964 240.244
R10252 GND.n3964 GND.n3934 240.244
R10253 GND.n3960 GND.n3934 240.244
R10254 GND.n3960 GND.n3959 240.244
R10255 GND.n3959 GND.n3958 240.244
R10256 GND.n3958 GND.n3940 240.244
R10257 GND.n3954 GND.n3940 240.244
R10258 GND.n3954 GND.n3953 240.244
R10259 GND.n3953 GND.n3952 240.244
R10260 GND.n3952 GND.n3946 240.244
R10261 GND.n3946 GND.n2263 240.244
R10262 GND.n4145 GND.n2263 240.244
R10263 GND.n4145 GND.n2264 240.244
R10264 GND.n4085 GND.n2264 240.244
R10265 GND.n4088 GND.n4085 240.244
R10266 GND.n4131 GND.n4088 240.244
R10267 GND.n4131 GND.n4128 240.244
R10268 GND.n4128 GND.n4089 240.244
R10269 GND.n4109 GND.n4089 240.244
R10270 GND.n4112 GND.n4109 240.244
R10271 GND.n4112 GND.n2253 240.244
R10272 GND.n4159 GND.n2253 240.244
R10273 GND.n4159 GND.n2254 240.244
R10274 GND.n4155 GND.n2254 240.244
R10275 GND.n4155 GND.n4154 240.244
R10276 GND.n4154 GND.n882 240.244
R10277 GND.n5534 GND.n882 240.244
R10278 GND.n5534 GND.n883 240.244
R10279 GND.n5530 GND.n883 240.244
R10280 GND.n5530 GND.n5527 240.244
R10281 GND.n5527 GND.n5526 240.244
R10282 GND.n4964 GND.n1224 240.244
R10283 GND.n4960 GND.n1224 240.244
R10284 GND.n4960 GND.n1229 240.244
R10285 GND.n4956 GND.n1229 240.244
R10286 GND.n4956 GND.n1231 240.244
R10287 GND.n4952 GND.n1231 240.244
R10288 GND.n4952 GND.n1237 240.244
R10289 GND.n4948 GND.n1237 240.244
R10290 GND.n4948 GND.n1239 240.244
R10291 GND.n4944 GND.n1239 240.244
R10292 GND.n4944 GND.n1245 240.244
R10293 GND.n4940 GND.n1245 240.244
R10294 GND.n4940 GND.n1247 240.244
R10295 GND.n4936 GND.n1247 240.244
R10296 GND.n4936 GND.n1253 240.244
R10297 GND.n4932 GND.n1253 240.244
R10298 GND.n4932 GND.n1255 240.244
R10299 GND.n4928 GND.n1255 240.244
R10300 GND.n4928 GND.n1261 240.244
R10301 GND.n4924 GND.n1261 240.244
R10302 GND.n4924 GND.n1263 240.244
R10303 GND.n4920 GND.n1263 240.244
R10304 GND.n4920 GND.n1269 240.244
R10305 GND.n4916 GND.n1269 240.244
R10306 GND.n4916 GND.n1271 240.244
R10307 GND.n4912 GND.n1271 240.244
R10308 GND.n4912 GND.n1277 240.244
R10309 GND.n4908 GND.n1277 240.244
R10310 GND.n4908 GND.n1279 240.244
R10311 GND.n4904 GND.n1279 240.244
R10312 GND.n4904 GND.n1285 240.244
R10313 GND.n4900 GND.n1285 240.244
R10314 GND.n4900 GND.n1287 240.244
R10315 GND.n4896 GND.n1287 240.244
R10316 GND.n4896 GND.n1293 240.244
R10317 GND.n4892 GND.n1293 240.244
R10318 GND.n4892 GND.n1295 240.244
R10319 GND.n4888 GND.n1295 240.244
R10320 GND.n4888 GND.n1301 240.244
R10321 GND.n4884 GND.n1301 240.244
R10322 GND.n4884 GND.n1303 240.244
R10323 GND.n4880 GND.n1303 240.244
R10324 GND.n4880 GND.n1309 240.244
R10325 GND.n4876 GND.n1309 240.244
R10326 GND.n4876 GND.n1311 240.244
R10327 GND.n4872 GND.n1311 240.244
R10328 GND.n4872 GND.n1317 240.244
R10329 GND.n4868 GND.n1317 240.244
R10330 GND.n4868 GND.n1319 240.244
R10331 GND.n4864 GND.n1319 240.244
R10332 GND.n4864 GND.n1325 240.244
R10333 GND.n4860 GND.n1325 240.244
R10334 GND.n4860 GND.n1327 240.244
R10335 GND.n4856 GND.n1327 240.244
R10336 GND.n4856 GND.n1333 240.244
R10337 GND.n4852 GND.n1333 240.244
R10338 GND.n4852 GND.n1335 240.244
R10339 GND.n4848 GND.n1335 240.244
R10340 GND.n4848 GND.n1341 240.244
R10341 GND.n4844 GND.n1341 240.244
R10342 GND.n4844 GND.n1343 240.244
R10343 GND.n4840 GND.n1343 240.244
R10344 GND.n4840 GND.n1349 240.244
R10345 GND.n4307 GND.n2040 240.244
R10346 GND.n2049 GND.n2048 240.244
R10347 GND.n2051 GND.n2050 240.244
R10348 GND.n2059 GND.n2058 240.244
R10349 GND.n2067 GND.n2066 240.244
R10350 GND.n2069 GND.n2068 240.244
R10351 GND.n2077 GND.n2076 240.244
R10352 GND.n4263 GND.n4262 240.244
R10353 GND.n3981 GND.n2039 240.244
R10354 GND.n3981 GND.n3979 240.244
R10355 GND.n3979 GND.n2365 240.244
R10356 GND.n2365 GND.n2353 240.244
R10357 GND.n4002 GND.n2353 240.244
R10358 GND.n4006 GND.n4002 240.244
R10359 GND.n4006 GND.n4005 240.244
R10360 GND.n4005 GND.n2342 240.244
R10361 GND.n2342 GND.n2332 240.244
R10362 GND.n4027 GND.n2332 240.244
R10363 GND.n4030 GND.n4027 240.244
R10364 GND.n4030 GND.n4029 240.244
R10365 GND.n4029 GND.n2319 240.244
R10366 GND.n2319 GND.n2307 240.244
R10367 GND.n4051 GND.n2307 240.244
R10368 GND.n4055 GND.n4051 240.244
R10369 GND.n4055 GND.n4054 240.244
R10370 GND.n4054 GND.n2292 240.244
R10371 GND.n2297 GND.n2292 240.244
R10372 GND.n2297 GND.n2296 240.244
R10373 GND.n2296 GND.n2269 240.244
R10374 GND.n2278 GND.n2269 240.244
R10375 GND.n4135 GND.n2278 240.244
R10376 GND.n4135 GND.n4134 240.244
R10377 GND.n4134 GND.n2280 240.244
R10378 GND.n4091 GND.n2280 240.244
R10379 GND.n4105 GND.n4091 240.244
R10380 GND.n4118 GND.n4105 240.244
R10381 GND.n4118 GND.n4117 240.244
R10382 GND.n4117 GND.n2251 240.244
R10383 GND.n4163 GND.n2251 240.244
R10384 GND.n4164 GND.n4163 240.244
R10385 GND.n4164 GND.n2238 240.244
R10386 GND.n4176 GND.n2238 240.244
R10387 GND.n4177 GND.n4176 240.244
R10388 GND.n4177 GND.n871 240.244
R10389 GND.n5543 GND.n871 240.244
R10390 GND.n5543 GND.n872 240.244
R10391 GND.n872 GND.n862 240.244
R10392 GND.n862 GND.n850 240.244
R10393 GND.n5560 GND.n850 240.244
R10394 GND.n5560 GND.n851 240.244
R10395 GND.n851 GND.n840 240.244
R10396 GND.n840 GND.n830 240.244
R10397 GND.n5577 GND.n830 240.244
R10398 GND.n5577 GND.n831 240.244
R10399 GND.n831 GND.n821 240.244
R10400 GND.n821 GND.n813 240.244
R10401 GND.n5595 GND.n813 240.244
R10402 GND.n5595 GND.n803 240.244
R10403 GND.n5606 GND.n803 240.244
R10404 GND.n5652 GND.n5606 240.244
R10405 GND.n5610 GND.n5609 240.244
R10406 GND.n5612 GND.n5611 240.244
R10407 GND.n5616 GND.n5615 240.244
R10408 GND.n5618 GND.n5617 240.244
R10409 GND.n5622 GND.n5621 240.244
R10410 GND.n5624 GND.n5623 240.244
R10411 GND.n5627 GND.n5626 240.244
R10412 GND.n5714 GND.n714 240.244
R10413 GND.n3917 GND.n2414 240.244
R10414 GND.n2414 GND.n2361 240.244
R10415 GND.n3993 GND.n2361 240.244
R10416 GND.n3993 GND.n2356 240.244
R10417 GND.n4000 GND.n2356 240.244
R10418 GND.n4000 GND.n2351 240.244
R10419 GND.n2351 GND.n2339 240.244
R10420 GND.n4018 GND.n2339 240.244
R10421 GND.n4018 GND.n2334 240.244
R10422 GND.n4025 GND.n2334 240.244
R10423 GND.n4025 GND.n2329 240.244
R10424 GND.n2329 GND.n2315 240.244
R10425 GND.n4042 GND.n2315 240.244
R10426 GND.n4042 GND.n2310 240.244
R10427 GND.n4049 GND.n2310 240.244
R10428 GND.n4049 GND.n2305 240.244
R10429 GND.n2305 GND.n2288 240.244
R10430 GND.n4068 GND.n2288 240.244
R10431 GND.n4068 GND.n2289 240.244
R10432 GND.n2289 GND.n2285 240.244
R10433 GND.n2285 GND.n2266 240.244
R10434 GND.n4076 GND.n2266 240.244
R10435 GND.n4076 GND.n2277 240.244
R10436 GND.n4082 GND.n2277 240.244
R10437 GND.n4083 GND.n4082 240.244
R10438 GND.n4083 GND.n677 240.244
R10439 GND.n678 GND.n677 240.244
R10440 GND.n679 GND.n678 240.244
R10441 GND.n4114 GND.n679 240.244
R10442 GND.n4114 GND.n682 240.244
R10443 GND.n683 GND.n682 240.244
R10444 GND.n684 GND.n683 240.244
R10445 GND.n2248 GND.n684 240.244
R10446 GND.n2248 GND.n687 240.244
R10447 GND.n688 GND.n687 240.244
R10448 GND.n689 GND.n688 240.244
R10449 GND.n870 GND.n689 240.244
R10450 GND.n870 GND.n692 240.244
R10451 GND.n693 GND.n692 240.244
R10452 GND.n694 GND.n693 240.244
R10453 GND.n848 GND.n694 240.244
R10454 GND.n848 GND.n697 240.244
R10455 GND.n698 GND.n697 240.244
R10456 GND.n699 GND.n698 240.244
R10457 GND.n829 GND.n699 240.244
R10458 GND.n829 GND.n702 240.244
R10459 GND.n703 GND.n702 240.244
R10460 GND.n704 GND.n703 240.244
R10461 GND.n812 GND.n704 240.244
R10462 GND.n812 GND.n707 240.244
R10463 GND.n708 GND.n707 240.244
R10464 GND.n709 GND.n708 240.244
R10465 GND.n3339 GND.n3338 240.132
R10466 GND.n1959 GND.n1958 240.132
R10467 GND.n711 GND.t64 224.174
R10468 GND.n767 GND.t88 224.174
R10469 GND.n794 GND.t73 224.174
R10470 GND.n1550 GND.t85 224.174
R10471 GND.n1576 GND.t67 224.174
R10472 GND.n1618 GND.t44 224.174
R10473 GND.n2821 GND.t57 224.174
R10474 GND.n2097 GND.t111 224.174
R10475 GND.n3253 GND.t105 224.174
R10476 GND.n2006 GND.t27 224.174
R10477 GND.n2118 GND.t101 224.174
R10478 GND.n1395 GND.t54 224.174
R10479 GND.n1415 GND.t41 224.174
R10480 GND.n4264 GND.t48 224.174
R10481 GND.n3312 GND.t37 204.78
R10482 GND.n3723 GND.t60 204.78
R10483 GND.n3318 GND.t77 204.78
R10484 GND.n2000 GND.t91 204.78
R10485 GND.n4309 GND.n2004 199.319
R10486 GND.n4573 GND.n1553 199.319
R10487 GND.n4572 GND.n1553 199.319
R10488 GND.n3340 GND.n3337 186.49
R10489 GND.n1960 GND.n1957 186.49
R10490 GND.n96 GND.n95 185
R10491 GND.n94 GND.n93 185
R10492 GND.n73 GND.n72 185
R10493 GND.n88 GND.n87 185
R10494 GND.n86 GND.n85 185
R10495 GND.n77 GND.n76 185
R10496 GND.n80 GND.n79 185
R10497 GND.n133 GND.n132 185
R10498 GND.n131 GND.n130 185
R10499 GND.n110 GND.n109 185
R10500 GND.n125 GND.n124 185
R10501 GND.n123 GND.n122 185
R10502 GND.n114 GND.n113 185
R10503 GND.n117 GND.n116 185
R10504 GND.n165 GND.n164 185
R10505 GND.n163 GND.n162 185
R10506 GND.n142 GND.n141 185
R10507 GND.n157 GND.n156 185
R10508 GND.n155 GND.n154 185
R10509 GND.n146 GND.n145 185
R10510 GND.n149 GND.n148 185
R10511 GND.n202 GND.n201 185
R10512 GND.n200 GND.n199 185
R10513 GND.n179 GND.n178 185
R10514 GND.n194 GND.n193 185
R10515 GND.n192 GND.n191 185
R10516 GND.n183 GND.n182 185
R10517 GND.n186 GND.n185 185
R10518 GND.n27 GND.n26 185
R10519 GND.n25 GND.n24 185
R10520 GND.n4 GND.n3 185
R10521 GND.n19 GND.n18 185
R10522 GND.n17 GND.n16 185
R10523 GND.n8 GND.n7 185
R10524 GND.n11 GND.n10 185
R10525 GND.n64 GND.n63 185
R10526 GND.n62 GND.n61 185
R10527 GND.n41 GND.n40 185
R10528 GND.n56 GND.n55 185
R10529 GND.n54 GND.n53 185
R10530 GND.n45 GND.n44 185
R10531 GND.n48 GND.n47 185
R10532 GND.n529 GND.n528 185
R10533 GND.n527 GND.n526 185
R10534 GND.n506 GND.n505 185
R10535 GND.n521 GND.n520 185
R10536 GND.n519 GND.n518 185
R10537 GND.n510 GND.n509 185
R10538 GND.n513 GND.n512 185
R10539 GND.n492 GND.n491 185
R10540 GND.n490 GND.n489 185
R10541 GND.n469 GND.n468 185
R10542 GND.n484 GND.n483 185
R10543 GND.n482 GND.n481 185
R10544 GND.n473 GND.n472 185
R10545 GND.n476 GND.n475 185
R10546 GND.n598 GND.n597 185
R10547 GND.n596 GND.n595 185
R10548 GND.n575 GND.n574 185
R10549 GND.n590 GND.n589 185
R10550 GND.n588 GND.n587 185
R10551 GND.n579 GND.n578 185
R10552 GND.n582 GND.n581 185
R10553 GND.n561 GND.n560 185
R10554 GND.n559 GND.n558 185
R10555 GND.n538 GND.n537 185
R10556 GND.n553 GND.n552 185
R10557 GND.n551 GND.n550 185
R10558 GND.n542 GND.n541 185
R10559 GND.n545 GND.n544 185
R10560 GND.n668 GND.n667 185
R10561 GND.n666 GND.n665 185
R10562 GND.n645 GND.n644 185
R10563 GND.n660 GND.n659 185
R10564 GND.n658 GND.n657 185
R10565 GND.n649 GND.n648 185
R10566 GND.n652 GND.n651 185
R10567 GND.n631 GND.n630 185
R10568 GND.n629 GND.n628 185
R10569 GND.n608 GND.n607 185
R10570 GND.n623 GND.n622 185
R10571 GND.n621 GND.n620 185
R10572 GND.n612 GND.n611 185
R10573 GND.n615 GND.n614 185
R10574 GND.n332 GND.n331 185
R10575 GND.n330 GND.n329 185
R10576 GND.n309 GND.n308 185
R10577 GND.n324 GND.n323 185
R10578 GND.n322 GND.n321 185
R10579 GND.n313 GND.n312 185
R10580 GND.n316 GND.n315 185
R10581 GND.n300 GND.n299 185
R10582 GND.n298 GND.n297 185
R10583 GND.n277 GND.n276 185
R10584 GND.n292 GND.n291 185
R10585 GND.n290 GND.n289 185
R10586 GND.n281 GND.n280 185
R10587 GND.n284 GND.n283 185
R10588 GND.n268 GND.n267 185
R10589 GND.n266 GND.n265 185
R10590 GND.n245 GND.n244 185
R10591 GND.n260 GND.n259 185
R10592 GND.n258 GND.n257 185
R10593 GND.n249 GND.n248 185
R10594 GND.n252 GND.n251 185
R10595 GND.n237 GND.n236 185
R10596 GND.n235 GND.n234 185
R10597 GND.n214 GND.n213 185
R10598 GND.n229 GND.n228 185
R10599 GND.n227 GND.n226 185
R10600 GND.n218 GND.n217 185
R10601 GND.n221 GND.n220 185
R10602 GND.n459 GND.n458 185
R10603 GND.n457 GND.n456 185
R10604 GND.n436 GND.n435 185
R10605 GND.n451 GND.n450 185
R10606 GND.n449 GND.n448 185
R10607 GND.n440 GND.n439 185
R10608 GND.n443 GND.n442 185
R10609 GND.n427 GND.n426 185
R10610 GND.n425 GND.n424 185
R10611 GND.n404 GND.n403 185
R10612 GND.n419 GND.n418 185
R10613 GND.n417 GND.n416 185
R10614 GND.n408 GND.n407 185
R10615 GND.n411 GND.n410 185
R10616 GND.n395 GND.n394 185
R10617 GND.n393 GND.n392 185
R10618 GND.n372 GND.n371 185
R10619 GND.n387 GND.n386 185
R10620 GND.n385 GND.n384 185
R10621 GND.n376 GND.n375 185
R10622 GND.n379 GND.n378 185
R10623 GND.n364 GND.n363 185
R10624 GND.n362 GND.n361 185
R10625 GND.n341 GND.n340 185
R10626 GND.n356 GND.n355 185
R10627 GND.n354 GND.n353 185
R10628 GND.n345 GND.n344 185
R10629 GND.n348 GND.n347 185
R10630 GND.n3313 GND.t36 178.987
R10631 GND.n3724 GND.t61 178.987
R10632 GND.n712 GND.t65 178.987
R10633 GND.n3319 GND.t76 178.987
R10634 GND.n2001 GND.t92 178.987
R10635 GND.n768 GND.t89 178.987
R10636 GND.n795 GND.t74 178.987
R10637 GND.n1551 GND.t86 178.987
R10638 GND.n1577 GND.t68 178.987
R10639 GND.n1619 GND.t45 178.987
R10640 GND.n2822 GND.t56 178.987
R10641 GND.n2098 GND.t112 178.987
R10642 GND.n3254 GND.t104 178.987
R10643 GND.n2007 GND.t26 178.987
R10644 GND.n2119 GND.t100 178.987
R10645 GND.n1396 GND.t53 178.987
R10646 GND.n1416 GND.t40 178.987
R10647 GND.n4265 GND.t47 178.987
R10648 GND.n5367 GND.n5366 164.363
R10649 GND.n5368 GND.n5367 164.363
R10650 GND.n5368 GND.n978 164.363
R10651 GND.n5376 GND.n978 164.363
R10652 GND.n5377 GND.n5376 164.363
R10653 GND.n5378 GND.n5377 164.363
R10654 GND.n5378 GND.n972 164.363
R10655 GND.n5386 GND.n972 164.363
R10656 GND.n5387 GND.n5386 164.363
R10657 GND.n5388 GND.n5387 164.363
R10658 GND.n5388 GND.n966 164.363
R10659 GND.n5396 GND.n966 164.363
R10660 GND.n5397 GND.n5396 164.363
R10661 GND.n5398 GND.n5397 164.363
R10662 GND.n5398 GND.n960 164.363
R10663 GND.n5406 GND.n960 164.363
R10664 GND.n5407 GND.n5406 164.363
R10665 GND.n5408 GND.n5407 164.363
R10666 GND.n5408 GND.n954 164.363
R10667 GND.n5416 GND.n954 164.363
R10668 GND.n5417 GND.n5416 164.363
R10669 GND.n5418 GND.n5417 164.363
R10670 GND.n5418 GND.n948 164.363
R10671 GND.n5426 GND.n948 164.363
R10672 GND.n5427 GND.n5426 164.363
R10673 GND.n5428 GND.n5427 164.363
R10674 GND.n5428 GND.n942 164.363
R10675 GND.n5436 GND.n942 164.363
R10676 GND.n5437 GND.n5436 164.363
R10677 GND.n5438 GND.n5437 164.363
R10678 GND.n5438 GND.n936 164.363
R10679 GND.n5446 GND.n936 164.363
R10680 GND.n5447 GND.n5446 164.363
R10681 GND.n5448 GND.n5447 164.363
R10682 GND.n5448 GND.n930 164.363
R10683 GND.n5456 GND.n930 164.363
R10684 GND.n5457 GND.n5456 164.363
R10685 GND.n5458 GND.n5457 164.363
R10686 GND.n5458 GND.n924 164.363
R10687 GND.n5466 GND.n924 164.363
R10688 GND.n5467 GND.n5466 164.363
R10689 GND.n5468 GND.n5467 164.363
R10690 GND.n5468 GND.n918 164.363
R10691 GND.n5476 GND.n918 164.363
R10692 GND.n5477 GND.n5476 164.363
R10693 GND.n5478 GND.n5477 164.363
R10694 GND.n5478 GND.n912 164.363
R10695 GND.n5486 GND.n912 164.363
R10696 GND.n5487 GND.n5486 164.363
R10697 GND.n5488 GND.n5487 164.363
R10698 GND.n5488 GND.n906 164.363
R10699 GND.n5496 GND.n906 164.363
R10700 GND.n5497 GND.n5496 164.363
R10701 GND.n5498 GND.n5497 164.363
R10702 GND.n5498 GND.n900 164.363
R10703 GND.n5506 GND.n900 164.363
R10704 GND.n5507 GND.n5506 164.363
R10705 GND.n5508 GND.n5507 164.363
R10706 GND.n5508 GND.n894 164.363
R10707 GND.n5517 GND.n894 164.363
R10708 GND.n5518 GND.n5517 164.363
R10709 GND.n5519 GND.n5518 164.363
R10710 GND.n5519 GND.n724 164.363
R10711 GND.n4372 GND.n1968 163.367
R10712 GND.n4369 GND.n1999 163.367
R10713 GND.n4365 GND.n4364 163.367
R10714 GND.n4361 GND.n4360 163.367
R10715 GND.n4357 GND.n4356 163.367
R10716 GND.n4353 GND.n4352 163.367
R10717 GND.n4349 GND.n4348 163.367
R10718 GND.n4345 GND.n4344 163.367
R10719 GND.n4341 GND.n4340 163.367
R10720 GND.n4337 GND.n4336 163.367
R10721 GND.n4333 GND.n4332 163.367
R10722 GND.n4329 GND.n4328 163.367
R10723 GND.n4325 GND.n4324 163.367
R10724 GND.n4320 GND.n4319 163.367
R10725 GND.n4316 GND.n4315 163.367
R10726 GND.n3727 GND.n3726 163.367
R10727 GND.n3731 GND.n3730 163.367
R10728 GND.n3735 GND.n3734 163.367
R10729 GND.n3739 GND.n3738 163.367
R10730 GND.n3743 GND.n3742 163.367
R10731 GND.n3747 GND.n3746 163.367
R10732 GND.n3751 GND.n3750 163.367
R10733 GND.n3755 GND.n3754 163.367
R10734 GND.n3759 GND.n3758 163.367
R10735 GND.n3763 GND.n3762 163.367
R10736 GND.n3767 GND.n3766 163.367
R10737 GND.n3771 GND.n3770 163.367
R10738 GND.n3775 GND.n3774 163.367
R10739 GND.n3779 GND.n3778 163.367
R10740 GND.n3478 GND.n3298 163.367
R10741 GND.n3478 GND.n1748 163.367
R10742 GND.n3490 GND.n1748 163.367
R10743 GND.n3490 GND.n1756 163.367
R10744 GND.n3494 GND.n1756 163.367
R10745 GND.n3495 GND.n3494 163.367
R10746 GND.n3496 GND.n3495 163.367
R10747 GND.n3496 GND.n1768 163.367
R10748 GND.n3502 GND.n1768 163.367
R10749 GND.n3502 GND.n1776 163.367
R10750 GND.n2537 GND.n1776 163.367
R10751 GND.n3541 GND.n2537 163.367
R10752 GND.n3542 GND.n3541 163.367
R10753 GND.n3542 GND.n1788 163.367
R10754 GND.n3548 GND.n1788 163.367
R10755 GND.n3548 GND.n1796 163.367
R10756 GND.n2530 GND.n1796 163.367
R10757 GND.n3573 GND.n2530 163.367
R10758 GND.n3574 GND.n3573 163.367
R10759 GND.n3574 GND.n1808 163.367
R10760 GND.n3580 GND.n1808 163.367
R10761 GND.n3580 GND.n1815 163.367
R10762 GND.n2521 GND.n1815 163.367
R10763 GND.n3605 GND.n2521 163.367
R10764 GND.n3606 GND.n3605 163.367
R10765 GND.n3606 GND.n1826 163.367
R10766 GND.n3610 GND.n1826 163.367
R10767 GND.n3610 GND.n1834 163.367
R10768 GND.n3625 GND.n1834 163.367
R10769 GND.n3625 GND.n2513 163.367
R10770 GND.n3639 GND.n2513 163.367
R10771 GND.n3639 GND.n2514 163.367
R10772 GND.n2514 GND.n2507 163.367
R10773 GND.n3634 GND.n2507 163.367
R10774 GND.n3634 GND.n1855 163.367
R10775 GND.n3630 GND.n1855 163.367
R10776 GND.n3630 GND.n1863 163.367
R10777 GND.n2500 GND.n1863 163.367
R10778 GND.n3663 GND.n2500 163.367
R10779 GND.n3663 GND.n1880 163.367
R10780 GND.n3667 GND.n1880 163.367
R10781 GND.n3667 GND.n1889 163.367
R10782 GND.n2497 GND.n1889 163.367
R10783 GND.n3675 GND.n2497 163.367
R10784 GND.n3675 GND.n2498 163.367
R10785 GND.n3671 GND.n2498 163.367
R10786 GND.n3671 GND.n2481 163.367
R10787 GND.n3708 GND.n2481 163.367
R10788 GND.n3708 GND.n1919 163.367
R10789 GND.n3712 GND.n1919 163.367
R10790 GND.n3712 GND.n1927 163.367
R10791 GND.n3716 GND.n1927 163.367
R10792 GND.n3720 GND.n3716 163.367
R10793 GND.n3720 GND.n1943 163.367
R10794 GND.n3783 GND.n1943 163.367
R10795 GND.n3358 GND.n3331 163.367
R10796 GND.n3362 GND.n3331 163.367
R10797 GND.n3366 GND.n3364 163.367
R10798 GND.n3370 GND.n3329 163.367
R10799 GND.n3374 GND.n3372 163.367
R10800 GND.n3378 GND.n3327 163.367
R10801 GND.n3382 GND.n3380 163.367
R10802 GND.n3386 GND.n3325 163.367
R10803 GND.n3390 GND.n3388 163.367
R10804 GND.n3394 GND.n3323 163.367
R10805 GND.n3398 GND.n3396 163.367
R10806 GND.n3402 GND.n3321 163.367
R10807 GND.n3406 GND.n3404 163.367
R10808 GND.n3411 GND.n3317 163.367
R10809 GND.n3414 GND.n3413 163.367
R10810 GND.n3421 GND.n3418 163.367
R10811 GND.n3425 GND.n3423 163.367
R10812 GND.n3429 GND.n3311 163.367
R10813 GND.n3433 GND.n3431 163.367
R10814 GND.n3437 GND.n3309 163.367
R10815 GND.n3441 GND.n3439 163.367
R10816 GND.n3445 GND.n3307 163.367
R10817 GND.n3449 GND.n3447 163.367
R10818 GND.n3453 GND.n3305 163.367
R10819 GND.n3457 GND.n3455 163.367
R10820 GND.n3461 GND.n3303 163.367
R10821 GND.n3465 GND.n3463 163.367
R10822 GND.n3469 GND.n3301 163.367
R10823 GND.n3472 GND.n3471 163.367
R10824 GND.n3355 GND.n1750 163.367
R10825 GND.n4502 GND.n1750 163.367
R10826 GND.n4502 GND.n1751 163.367
R10827 GND.n4498 GND.n1751 163.367
R10828 GND.n4498 GND.n1754 163.367
R10829 GND.n2562 GND.n1754 163.367
R10830 GND.n2562 GND.n1770 163.367
R10831 GND.n4488 GND.n1770 163.367
R10832 GND.n4488 GND.n1771 163.367
R10833 GND.n4484 GND.n1771 163.367
R10834 GND.n4484 GND.n1774 163.367
R10835 GND.n3539 GND.n1774 163.367
R10836 GND.n3539 GND.n1790 163.367
R10837 GND.n4474 GND.n1790 163.367
R10838 GND.n4474 GND.n1791 163.367
R10839 GND.n4470 GND.n1791 163.367
R10840 GND.n4470 GND.n1794 163.367
R10841 GND.n3571 GND.n1794 163.367
R10842 GND.n3571 GND.n1809 163.367
R10843 GND.n4460 GND.n1809 163.367
R10844 GND.n4460 GND.n1810 163.367
R10845 GND.n4456 GND.n1810 163.367
R10846 GND.n4456 GND.n1813 163.367
R10847 GND.n3603 GND.n1813 163.367
R10848 GND.n3603 GND.n1828 163.367
R10849 GND.n4446 GND.n1828 163.367
R10850 GND.n4446 GND.n1829 163.367
R10851 GND.n4442 GND.n1829 163.367
R10852 GND.n4442 GND.n1832 163.367
R10853 GND.n2511 GND.n1832 163.367
R10854 GND.n3641 GND.n2511 163.367
R10855 GND.n3641 GND.n2509 163.367
R10856 GND.n3645 GND.n2509 163.367
R10857 GND.n3645 GND.n1857 163.367
R10858 GND.n4425 GND.n1857 163.367
R10859 GND.n4425 GND.n1858 163.367
R10860 GND.n4421 GND.n1858 163.367
R10861 GND.n4421 GND.n1861 163.367
R10862 GND.n1883 GND.n1861 163.367
R10863 GND.n4412 GND.n1883 163.367
R10864 GND.n4412 GND.n1884 163.367
R10865 GND.n4408 GND.n1884 163.367
R10866 GND.n4408 GND.n1887 163.367
R10867 GND.n3683 GND.n1887 163.367
R10868 GND.n3683 GND.n3676 163.367
R10869 GND.n3679 GND.n3676 163.367
R10870 GND.n3679 GND.n3678 163.367
R10871 GND.n3678 GND.n1921 163.367
R10872 GND.n4391 GND.n1921 163.367
R10873 GND.n4391 GND.n1922 163.367
R10874 GND.n4387 GND.n1922 163.367
R10875 GND.n4387 GND.n1925 163.367
R10876 GND.n1945 GND.n1925 163.367
R10877 GND.n4377 GND.n1945 163.367
R10878 GND.n4377 GND.n1946 163.367
R10879 GND.n1966 GND.n1965 156.462
R10880 GND.n272 GND.n240 153.042
R10881 GND.n336 GND.n335 152.079
R10882 GND.n304 GND.n303 152.079
R10883 GND.n272 GND.n271 152.079
R10884 GND.n3345 GND.n3344 152
R10885 GND.n3346 GND.n3335 152
R10886 GND.n3348 GND.n3347 152
R10887 GND.n3350 GND.n3333 152
R10888 GND.n3352 GND.n3351 152
R10889 GND.n1964 GND.n1948 152
R10890 GND.n1956 GND.n1949 152
R10891 GND.n1955 GND.n1954 152
R10892 GND.n1953 GND.n1950 152
R10893 GND.n1951 GND.t106 150.546
R10894 GND.t126 GND.n78 147.661
R10895 GND.t147 GND.n115 147.661
R10896 GND.t178 GND.n147 147.661
R10897 GND.t137 GND.n184 147.661
R10898 GND.t169 GND.n9 147.661
R10899 GND.t167 GND.n46 147.661
R10900 GND.t170 GND.n511 147.661
R10901 GND.t150 GND.n474 147.661
R10902 GND.t159 GND.n580 147.661
R10903 GND.t141 GND.n543 147.661
R10904 GND.t168 GND.n650 147.661
R10905 GND.t172 GND.n613 147.661
R10906 GND.t15 GND.n314 147.661
R10907 GND.t10 GND.n282 147.661
R10908 GND.t13 GND.n250 147.661
R10909 GND.t1 GND.n219 147.661
R10910 GND.t18 GND.n441 147.661
R10911 GND.t3 GND.n409 147.661
R10912 GND.t23 GND.n377 147.661
R10913 GND.t21 GND.n346 147.661
R10914 GND.n4313 GND.n1985 143.351
R10915 GND.n4313 GND.n1984 143.351
R10916 GND.n3416 GND.n3415 143.351
R10917 GND.n3417 GND.n3416 143.351
R10918 GND.n3342 GND.t28 130.484
R10919 GND.n3351 GND.t81 126.766
R10920 GND.n3349 GND.t93 126.766
R10921 GND.n3335 GND.t69 126.766
R10922 GND.n3343 GND.t113 126.766
R10923 GND.n1952 GND.t49 126.766
R10924 GND.n1954 GND.t31 126.766
R10925 GND.n1963 GND.t78 126.766
R10926 GND.n1965 GND.t96 126.766
R10927 GND.n4660 GND.n1554 110.912
R10928 GND.n4314 GND.n4312 110.912
R10929 GND.n95 GND.n94 104.615
R10930 GND.n94 GND.n72 104.615
R10931 GND.n87 GND.n72 104.615
R10932 GND.n87 GND.n86 104.615
R10933 GND.n86 GND.n76 104.615
R10934 GND.n79 GND.n76 104.615
R10935 GND.n132 GND.n131 104.615
R10936 GND.n131 GND.n109 104.615
R10937 GND.n124 GND.n109 104.615
R10938 GND.n124 GND.n123 104.615
R10939 GND.n123 GND.n113 104.615
R10940 GND.n116 GND.n113 104.615
R10941 GND.n164 GND.n163 104.615
R10942 GND.n163 GND.n141 104.615
R10943 GND.n156 GND.n141 104.615
R10944 GND.n156 GND.n155 104.615
R10945 GND.n155 GND.n145 104.615
R10946 GND.n148 GND.n145 104.615
R10947 GND.n201 GND.n200 104.615
R10948 GND.n200 GND.n178 104.615
R10949 GND.n193 GND.n178 104.615
R10950 GND.n193 GND.n192 104.615
R10951 GND.n192 GND.n182 104.615
R10952 GND.n185 GND.n182 104.615
R10953 GND.n26 GND.n25 104.615
R10954 GND.n25 GND.n3 104.615
R10955 GND.n18 GND.n3 104.615
R10956 GND.n18 GND.n17 104.615
R10957 GND.n17 GND.n7 104.615
R10958 GND.n10 GND.n7 104.615
R10959 GND.n63 GND.n62 104.615
R10960 GND.n62 GND.n40 104.615
R10961 GND.n55 GND.n40 104.615
R10962 GND.n55 GND.n54 104.615
R10963 GND.n54 GND.n44 104.615
R10964 GND.n47 GND.n44 104.615
R10965 GND.n528 GND.n527 104.615
R10966 GND.n527 GND.n505 104.615
R10967 GND.n520 GND.n505 104.615
R10968 GND.n520 GND.n519 104.615
R10969 GND.n519 GND.n509 104.615
R10970 GND.n512 GND.n509 104.615
R10971 GND.n491 GND.n490 104.615
R10972 GND.n490 GND.n468 104.615
R10973 GND.n483 GND.n468 104.615
R10974 GND.n483 GND.n482 104.615
R10975 GND.n482 GND.n472 104.615
R10976 GND.n475 GND.n472 104.615
R10977 GND.n597 GND.n596 104.615
R10978 GND.n596 GND.n574 104.615
R10979 GND.n589 GND.n574 104.615
R10980 GND.n589 GND.n588 104.615
R10981 GND.n588 GND.n578 104.615
R10982 GND.n581 GND.n578 104.615
R10983 GND.n560 GND.n559 104.615
R10984 GND.n559 GND.n537 104.615
R10985 GND.n552 GND.n537 104.615
R10986 GND.n552 GND.n551 104.615
R10987 GND.n551 GND.n541 104.615
R10988 GND.n544 GND.n541 104.615
R10989 GND.n667 GND.n666 104.615
R10990 GND.n666 GND.n644 104.615
R10991 GND.n659 GND.n644 104.615
R10992 GND.n659 GND.n658 104.615
R10993 GND.n658 GND.n648 104.615
R10994 GND.n651 GND.n648 104.615
R10995 GND.n630 GND.n629 104.615
R10996 GND.n629 GND.n607 104.615
R10997 GND.n622 GND.n607 104.615
R10998 GND.n622 GND.n621 104.615
R10999 GND.n621 GND.n611 104.615
R11000 GND.n614 GND.n611 104.615
R11001 GND.n331 GND.n330 104.615
R11002 GND.n330 GND.n308 104.615
R11003 GND.n323 GND.n308 104.615
R11004 GND.n323 GND.n322 104.615
R11005 GND.n322 GND.n312 104.615
R11006 GND.n315 GND.n312 104.615
R11007 GND.n299 GND.n298 104.615
R11008 GND.n298 GND.n276 104.615
R11009 GND.n291 GND.n276 104.615
R11010 GND.n291 GND.n290 104.615
R11011 GND.n290 GND.n280 104.615
R11012 GND.n283 GND.n280 104.615
R11013 GND.n267 GND.n266 104.615
R11014 GND.n266 GND.n244 104.615
R11015 GND.n259 GND.n244 104.615
R11016 GND.n259 GND.n258 104.615
R11017 GND.n258 GND.n248 104.615
R11018 GND.n251 GND.n248 104.615
R11019 GND.n236 GND.n235 104.615
R11020 GND.n235 GND.n213 104.615
R11021 GND.n228 GND.n213 104.615
R11022 GND.n228 GND.n227 104.615
R11023 GND.n227 GND.n217 104.615
R11024 GND.n220 GND.n217 104.615
R11025 GND.n458 GND.n457 104.615
R11026 GND.n457 GND.n435 104.615
R11027 GND.n450 GND.n435 104.615
R11028 GND.n450 GND.n449 104.615
R11029 GND.n449 GND.n439 104.615
R11030 GND.n442 GND.n439 104.615
R11031 GND.n426 GND.n425 104.615
R11032 GND.n425 GND.n403 104.615
R11033 GND.n418 GND.n403 104.615
R11034 GND.n418 GND.n417 104.615
R11035 GND.n417 GND.n407 104.615
R11036 GND.n410 GND.n407 104.615
R11037 GND.n394 GND.n393 104.615
R11038 GND.n393 GND.n371 104.615
R11039 GND.n386 GND.n371 104.615
R11040 GND.n386 GND.n385 104.615
R11041 GND.n385 GND.n375 104.615
R11042 GND.n378 GND.n375 104.615
R11043 GND.n363 GND.n362 104.615
R11044 GND.n362 GND.n340 104.615
R11045 GND.n355 GND.n340 104.615
R11046 GND.n355 GND.n354 104.615
R11047 GND.n354 GND.n344 104.615
R11048 GND.n347 GND.n344 104.615
R11049 GND.n747 GND.n741 99.6594
R11050 GND.n749 GND.n740 99.6594
R11051 GND.n753 GND.n739 99.6594
R11052 GND.n755 GND.n738 99.6594
R11053 GND.n759 GND.n737 99.6594
R11054 GND.n761 GND.n736 99.6594
R11055 GND.n765 GND.n735 99.6594
R11056 GND.n769 GND.n734 99.6594
R11057 GND.n773 GND.n733 99.6594
R11058 GND.n775 GND.n732 99.6594
R11059 GND.n779 GND.n731 99.6594
R11060 GND.n781 GND.n730 99.6594
R11061 GND.n785 GND.n729 99.6594
R11062 GND.n787 GND.n728 99.6594
R11063 GND.n791 GND.n727 99.6594
R11064 GND.n793 GND.n726 99.6594
R11065 GND.n5657 GND.n725 99.6594
R11066 GND.n2411 GND.n2012 99.6594
R11067 GND.n2407 GND.n2013 99.6594
R11068 GND.n2403 GND.n2014 99.6594
R11069 GND.n2399 GND.n2015 99.6594
R11070 GND.n2395 GND.n2016 99.6594
R11071 GND.n2391 GND.n2017 99.6594
R11072 GND.n2387 GND.n2018 99.6594
R11073 GND.n2020 GND.n2004 99.6594
R11074 GND.n2021 GND.n2010 99.6594
R11075 GND.n2129 GND.n2022 99.6594
R11076 GND.n2137 GND.n2023 99.6594
R11077 GND.n2139 GND.n2024 99.6594
R11078 GND.n2147 GND.n2025 99.6594
R11079 GND.n2149 GND.n2026 99.6594
R11080 GND.n2157 GND.n2027 99.6594
R11081 GND.n2159 GND.n2028 99.6594
R11082 GND.n2116 GND.n2029 99.6594
R11083 GND.n4582 GND.n1535 99.6594
R11084 GND.n4581 GND.n1538 99.6594
R11085 GND.n4579 GND.n1540 99.6594
R11086 GND.n4578 GND.n1543 99.6594
R11087 GND.n4576 GND.n1545 99.6594
R11088 GND.n4575 GND.n1548 99.6594
R11089 GND.n4572 GND.n1555 99.6594
R11090 GND.n4571 GND.n1558 99.6594
R11091 GND.n4569 GND.n1560 99.6594
R11092 GND.n4568 GND.n1563 99.6594
R11093 GND.n4566 GND.n1565 99.6594
R11094 GND.n4565 GND.n1568 99.6594
R11095 GND.n4563 GND.n1570 99.6594
R11096 GND.n4562 GND.n1573 99.6594
R11097 GND.n4560 GND.n1575 99.6594
R11098 GND.n4559 GND.n1524 99.6594
R11099 GND.n4836 GND.n4835 99.6594
R11100 GND.n4830 GND.n1350 99.6594
R11101 GND.n4827 GND.n1351 99.6594
R11102 GND.n4823 GND.n1352 99.6594
R11103 GND.n4819 GND.n1353 99.6594
R11104 GND.n4815 GND.n1354 99.6594
R11105 GND.n4811 GND.n1355 99.6594
R11106 GND.n4807 GND.n1356 99.6594
R11107 GND.n4802 GND.n1357 99.6594
R11108 GND.n4798 GND.n1358 99.6594
R11109 GND.n4794 GND.n1359 99.6594
R11110 GND.n4790 GND.n1360 99.6594
R11111 GND.n4786 GND.n1361 99.6594
R11112 GND.n4782 GND.n1362 99.6594
R11113 GND.n4778 GND.n1363 99.6594
R11114 GND.n4774 GND.n1364 99.6594
R11115 GND.n1414 GND.n1365 99.6594
R11116 GND.n1628 GND.n1583 99.6594
R11117 GND.n1630 GND.n1592 99.6594
R11118 GND.n1632 GND.n1631 99.6594
R11119 GND.n1633 GND.n1601 99.6594
R11120 GND.n1635 GND.n1608 99.6594
R11121 GND.n1637 GND.n1636 99.6594
R11122 GND.n1638 GND.n1617 99.6594
R11123 GND.n4585 GND.n4584 99.6594
R11124 GND.n2839 GND.n1366 99.6594
R11125 GND.n2837 GND.n1367 99.6594
R11126 GND.n2847 GND.n1368 99.6594
R11127 GND.n2833 GND.n1369 99.6594
R11128 GND.n2855 GND.n1370 99.6594
R11129 GND.n2829 GND.n1371 99.6594
R11130 GND.n2863 GND.n1372 99.6594
R11131 GND.n2825 GND.n1373 99.6594
R11132 GND.n3901 GND.n3900 99.6594
R11133 GND.n3899 GND.n2055 99.6594
R11134 GND.n3898 GND.n2062 99.6594
R11135 GND.n3896 GND.n3895 99.6594
R11136 GND.n3894 GND.n2073 99.6594
R11137 GND.n3893 GND.n2080 99.6594
R11138 GND.n3891 GND.n3890 99.6594
R11139 GND.n3889 GND.n2087 99.6594
R11140 GND.n3888 GND.n3887 99.6594
R11141 GND.n3886 GND.n2093 99.6594
R11142 GND.n3885 GND.n3884 99.6594
R11143 GND.n3883 GND.n2101 99.6594
R11144 GND.n3882 GND.n2107 99.6594
R11145 GND.n4549 GND.n4548 99.6594
R11146 GND.n1649 GND.n1648 99.6594
R11147 GND.n1651 GND.n1597 99.6594
R11148 GND.n1652 GND.n1604 99.6594
R11149 GND.n1654 GND.n1653 99.6594
R11150 GND.n1656 GND.n1613 99.6594
R11151 GND.n1657 GND.n1622 99.6594
R11152 GND.n1659 GND.n1658 99.6594
R11153 GND.n3239 GND.n1660 99.6594
R11154 GND.n3241 GND.n1661 99.6594
R11155 GND.n3249 GND.n1662 99.6594
R11156 GND.n3251 GND.n1663 99.6594
R11157 GND.n3262 GND.n1664 99.6594
R11158 GND.n4549 GND.n1588 99.6594
R11159 GND.n1649 GND.n1596 99.6594
R11160 GND.n1651 GND.n1650 99.6594
R11161 GND.n1652 GND.n1605 99.6594
R11162 GND.n1654 GND.n1612 99.6594
R11163 GND.n1656 GND.n1655 99.6594
R11164 GND.n1657 GND.n1623 99.6594
R11165 GND.n3238 GND.n1659 99.6594
R11166 GND.n3242 GND.n1660 99.6594
R11167 GND.n3248 GND.n1661 99.6594
R11168 GND.n3252 GND.n1662 99.6594
R11169 GND.n3261 GND.n1663 99.6594
R11170 GND.n3264 GND.n1664 99.6594
R11171 GND.n3882 GND.n2102 99.6594
R11172 GND.n3883 GND.n2100 99.6594
R11173 GND.n3885 GND.n2094 99.6594
R11174 GND.n3886 GND.n2092 99.6594
R11175 GND.n3888 GND.n2088 99.6594
R11176 GND.n3889 GND.n2086 99.6594
R11177 GND.n3891 GND.n2081 99.6594
R11178 GND.n3893 GND.n3892 99.6594
R11179 GND.n3894 GND.n2072 99.6594
R11180 GND.n3896 GND.n2063 99.6594
R11181 GND.n3898 GND.n3897 99.6594
R11182 GND.n3899 GND.n2054 99.6594
R11183 GND.n3901 GND.n2045 99.6594
R11184 GND.n2836 GND.n1366 99.6594
R11185 GND.n2846 GND.n1367 99.6594
R11186 GND.n2832 GND.n1368 99.6594
R11187 GND.n2854 GND.n1369 99.6594
R11188 GND.n2828 GND.n1370 99.6594
R11189 GND.n2862 GND.n1371 99.6594
R11190 GND.n2824 GND.n1372 99.6594
R11191 GND.n2820 GND.n1373 99.6594
R11192 GND.n4584 GND.n1626 99.6594
R11193 GND.n1638 GND.n1616 99.6594
R11194 GND.n1637 GND.n1609 99.6594
R11195 GND.n1635 GND.n1634 99.6594
R11196 GND.n1633 GND.n1600 99.6594
R11197 GND.n1632 GND.n1593 99.6594
R11198 GND.n1630 GND.n1629 99.6594
R11199 GND.n1628 GND.n1582 99.6594
R11200 GND.n4836 GND.n1377 99.6594
R11201 GND.n4828 GND.n1350 99.6594
R11202 GND.n4824 GND.n1351 99.6594
R11203 GND.n4820 GND.n1352 99.6594
R11204 GND.n4816 GND.n1353 99.6594
R11205 GND.n4812 GND.n1354 99.6594
R11206 GND.n4808 GND.n1355 99.6594
R11207 GND.n4803 GND.n1356 99.6594
R11208 GND.n4799 GND.n1357 99.6594
R11209 GND.n4795 GND.n1358 99.6594
R11210 GND.n4791 GND.n1359 99.6594
R11211 GND.n4787 GND.n1360 99.6594
R11212 GND.n4783 GND.n1361 99.6594
R11213 GND.n4779 GND.n1362 99.6594
R11214 GND.n4775 GND.n1363 99.6594
R11215 GND.n1413 GND.n1364 99.6594
R11216 GND.n4767 GND.n1365 99.6594
R11217 GND.n4559 GND.n4558 99.6594
R11218 GND.n4560 GND.n1574 99.6594
R11219 GND.n4562 GND.n4561 99.6594
R11220 GND.n4563 GND.n1569 99.6594
R11221 GND.n4565 GND.n4564 99.6594
R11222 GND.n4566 GND.n1564 99.6594
R11223 GND.n4568 GND.n4567 99.6594
R11224 GND.n4569 GND.n1559 99.6594
R11225 GND.n4571 GND.n4570 99.6594
R11226 GND.n4573 GND.n1549 99.6594
R11227 GND.n4575 GND.n4574 99.6594
R11228 GND.n4576 GND.n1544 99.6594
R11229 GND.n4578 GND.n4577 99.6594
R11230 GND.n4579 GND.n1539 99.6594
R11231 GND.n4581 GND.n4580 99.6594
R11232 GND.n4582 GND.n1534 99.6594
R11233 GND.n2408 GND.n2012 99.6594
R11234 GND.n2404 GND.n2013 99.6594
R11235 GND.n2400 GND.n2014 99.6594
R11236 GND.n2396 GND.n2015 99.6594
R11237 GND.n2392 GND.n2016 99.6594
R11238 GND.n2388 GND.n2017 99.6594
R11239 GND.n2019 GND.n2018 99.6594
R11240 GND.n4310 GND.n4309 99.6594
R11241 GND.n2130 GND.n2021 99.6594
R11242 GND.n2136 GND.n2022 99.6594
R11243 GND.n2140 GND.n2023 99.6594
R11244 GND.n2146 GND.n2024 99.6594
R11245 GND.n2150 GND.n2025 99.6594
R11246 GND.n2156 GND.n2026 99.6594
R11247 GND.n2160 GND.n2027 99.6594
R11248 GND.n2121 GND.n2028 99.6594
R11249 GND.n2168 GND.n2029 99.6594
R11250 GND.n796 GND.n725 99.6594
R11251 GND.n792 GND.n726 99.6594
R11252 GND.n788 GND.n727 99.6594
R11253 GND.n786 GND.n728 99.6594
R11254 GND.n782 GND.n729 99.6594
R11255 GND.n780 GND.n730 99.6594
R11256 GND.n776 GND.n731 99.6594
R11257 GND.n774 GND.n732 99.6594
R11258 GND.n770 GND.n733 99.6594
R11259 GND.n766 GND.n734 99.6594
R11260 GND.n762 GND.n735 99.6594
R11261 GND.n760 GND.n736 99.6594
R11262 GND.n756 GND.n737 99.6594
R11263 GND.n754 GND.n738 99.6594
R11264 GND.n750 GND.n739 99.6594
R11265 GND.n748 GND.n740 99.6594
R11266 GND.n743 GND.n741 99.6594
R11267 GND.n2040 GND.n2030 99.6594
R11268 GND.n2049 GND.n2031 99.6594
R11269 GND.n2051 GND.n2032 99.6594
R11270 GND.n2059 GND.n2033 99.6594
R11271 GND.n2067 GND.n2034 99.6594
R11272 GND.n2069 GND.n2035 99.6594
R11273 GND.n2077 GND.n2036 99.6594
R11274 GND.n4263 GND.n2037 99.6594
R11275 GND.n2048 GND.n2030 99.6594
R11276 GND.n2050 GND.n2031 99.6594
R11277 GND.n2058 GND.n2032 99.6594
R11278 GND.n2066 GND.n2033 99.6594
R11279 GND.n2068 GND.n2034 99.6594
R11280 GND.n2076 GND.n2035 99.6594
R11281 GND.n4262 GND.n2036 99.6594
R11282 GND.n2084 GND.n2037 99.6594
R11283 GND.n5651 GND.n716 99.6594
R11284 GND.n5610 GND.n717 99.6594
R11285 GND.n5612 GND.n718 99.6594
R11286 GND.n5616 GND.n719 99.6594
R11287 GND.n5618 GND.n720 99.6594
R11288 GND.n5622 GND.n721 99.6594
R11289 GND.n5624 GND.n722 99.6594
R11290 GND.n5627 GND.n723 99.6594
R11291 GND.n723 GND.n714 99.6594
R11292 GND.n5626 GND.n722 99.6594
R11293 GND.n5623 GND.n721 99.6594
R11294 GND.n5621 GND.n720 99.6594
R11295 GND.n5617 GND.n719 99.6594
R11296 GND.n5615 GND.n718 99.6594
R11297 GND.n5611 GND.n717 99.6594
R11298 GND.n5609 GND.n716 99.6594
R11299 GND.n3342 GND.n3341 81.8399
R11300 GND.n3343 GND.n3336 72.8411
R11301 GND.n3349 GND.n3334 72.8411
R11302 GND.n1963 GND.n1962 72.8411
R11303 GND.n4370 GND.n4369 71.676
R11304 GND.n4365 GND.n1998 71.676
R11305 GND.n4361 GND.n1997 71.676
R11306 GND.n4357 GND.n1996 71.676
R11307 GND.n4353 GND.n1995 71.676
R11308 GND.n4349 GND.n1994 71.676
R11309 GND.n4345 GND.n1993 71.676
R11310 GND.n4341 GND.n1992 71.676
R11311 GND.n4337 GND.n1991 71.676
R11312 GND.n4333 GND.n1990 71.676
R11313 GND.n4329 GND.n1989 71.676
R11314 GND.n4325 GND.n1988 71.676
R11315 GND.n4320 GND.n1987 71.676
R11316 GND.n4316 GND.n1986 71.676
R11317 GND.n3726 GND.n1984 71.676
R11318 GND.n3730 GND.n1983 71.676
R11319 GND.n3734 GND.n1982 71.676
R11320 GND.n3738 GND.n1981 71.676
R11321 GND.n3742 GND.n1980 71.676
R11322 GND.n3746 GND.n1979 71.676
R11323 GND.n3750 GND.n1978 71.676
R11324 GND.n3754 GND.n1977 71.676
R11325 GND.n3758 GND.n1976 71.676
R11326 GND.n3762 GND.n1975 71.676
R11327 GND.n3766 GND.n1974 71.676
R11328 GND.n3770 GND.n1973 71.676
R11329 GND.n3774 GND.n1972 71.676
R11330 GND.n3778 GND.n1971 71.676
R11331 GND.n2479 GND.n1970 71.676
R11332 GND.n3357 GND.n3356 71.676
R11333 GND.n3363 GND.n3362 71.676
R11334 GND.n3366 GND.n3365 71.676
R11335 GND.n3371 GND.n3370 71.676
R11336 GND.n3374 GND.n3373 71.676
R11337 GND.n3379 GND.n3378 71.676
R11338 GND.n3382 GND.n3381 71.676
R11339 GND.n3387 GND.n3386 71.676
R11340 GND.n3390 GND.n3389 71.676
R11341 GND.n3395 GND.n3394 71.676
R11342 GND.n3398 GND.n3397 71.676
R11343 GND.n3403 GND.n3402 71.676
R11344 GND.n3406 GND.n3405 71.676
R11345 GND.n3412 GND.n3411 71.676
R11346 GND.n3415 GND.n3414 71.676
R11347 GND.n3422 GND.n3421 71.676
R11348 GND.n3425 GND.n3424 71.676
R11349 GND.n3430 GND.n3429 71.676
R11350 GND.n3433 GND.n3432 71.676
R11351 GND.n3438 GND.n3437 71.676
R11352 GND.n3441 GND.n3440 71.676
R11353 GND.n3446 GND.n3445 71.676
R11354 GND.n3449 GND.n3448 71.676
R11355 GND.n3454 GND.n3453 71.676
R11356 GND.n3457 GND.n3456 71.676
R11357 GND.n3462 GND.n3461 71.676
R11358 GND.n3465 GND.n3464 71.676
R11359 GND.n3470 GND.n3469 71.676
R11360 GND.n3473 GND.n3472 71.676
R11361 GND.n3358 GND.n3357 71.676
R11362 GND.n3364 GND.n3363 71.676
R11363 GND.n3365 GND.n3329 71.676
R11364 GND.n3372 GND.n3371 71.676
R11365 GND.n3373 GND.n3327 71.676
R11366 GND.n3380 GND.n3379 71.676
R11367 GND.n3381 GND.n3325 71.676
R11368 GND.n3388 GND.n3387 71.676
R11369 GND.n3389 GND.n3323 71.676
R11370 GND.n3396 GND.n3395 71.676
R11371 GND.n3397 GND.n3321 71.676
R11372 GND.n3404 GND.n3403 71.676
R11373 GND.n3405 GND.n3317 71.676
R11374 GND.n3413 GND.n3412 71.676
R11375 GND.n3418 GND.n3417 71.676
R11376 GND.n3423 GND.n3422 71.676
R11377 GND.n3424 GND.n3311 71.676
R11378 GND.n3431 GND.n3430 71.676
R11379 GND.n3432 GND.n3309 71.676
R11380 GND.n3439 GND.n3438 71.676
R11381 GND.n3440 GND.n3307 71.676
R11382 GND.n3447 GND.n3446 71.676
R11383 GND.n3448 GND.n3305 71.676
R11384 GND.n3455 GND.n3454 71.676
R11385 GND.n3456 GND.n3303 71.676
R11386 GND.n3463 GND.n3462 71.676
R11387 GND.n3464 GND.n3301 71.676
R11388 GND.n3471 GND.n3470 71.676
R11389 GND.n3474 GND.n3473 71.676
R11390 GND.n3779 GND.n1970 71.676
R11391 GND.n3775 GND.n1971 71.676
R11392 GND.n3771 GND.n1972 71.676
R11393 GND.n3767 GND.n1973 71.676
R11394 GND.n3763 GND.n1974 71.676
R11395 GND.n3759 GND.n1975 71.676
R11396 GND.n3755 GND.n1976 71.676
R11397 GND.n3751 GND.n1977 71.676
R11398 GND.n3747 GND.n1978 71.676
R11399 GND.n3743 GND.n1979 71.676
R11400 GND.n3739 GND.n1980 71.676
R11401 GND.n3735 GND.n1981 71.676
R11402 GND.n3731 GND.n1982 71.676
R11403 GND.n3727 GND.n1983 71.676
R11404 GND.n4315 GND.n1985 71.676
R11405 GND.n4319 GND.n1986 71.676
R11406 GND.n4324 GND.n1987 71.676
R11407 GND.n4328 GND.n1988 71.676
R11408 GND.n4332 GND.n1989 71.676
R11409 GND.n4336 GND.n1990 71.676
R11410 GND.n4340 GND.n1991 71.676
R11411 GND.n4344 GND.n1992 71.676
R11412 GND.n4348 GND.n1993 71.676
R11413 GND.n4352 GND.n1994 71.676
R11414 GND.n4356 GND.n1995 71.676
R11415 GND.n4360 GND.n1996 71.676
R11416 GND.n4364 GND.n1997 71.676
R11417 GND.n1999 GND.n1998 71.676
R11418 GND.n4370 GND.n1968 71.676
R11419 GND.n3314 GND.n3313 59.5399
R11420 GND.n3725 GND.n3724 59.5399
R11421 GND.n3408 GND.n3319 59.5399
R11422 GND.n4322 GND.n2001 59.5399
R11423 GND.n3353 GND.n3352 59.1804
R11424 GND.n5713 GND.n724 57.5546
R11425 GND.n101 GND.n100 56.1363
R11426 GND.n103 GND.n102 56.1363
R11427 GND.n105 GND.n104 56.1363
R11428 GND.n170 GND.n169 56.1363
R11429 GND.n172 GND.n171 56.1363
R11430 GND.n174 GND.n173 56.1363
R11431 GND.n32 GND.n31 56.1363
R11432 GND.n34 GND.n33 56.1363
R11433 GND.n36 GND.n35 56.1363
R11434 GND.n501 GND.n500 56.1363
R11435 GND.n499 GND.n498 56.1363
R11436 GND.n497 GND.n496 56.1363
R11437 GND.n570 GND.n569 56.1363
R11438 GND.n568 GND.n567 56.1363
R11439 GND.n566 GND.n565 56.1363
R11440 GND.n640 GND.n639 56.1363
R11441 GND.n638 GND.n637 56.1363
R11442 GND.n636 GND.n635 56.1363
R11443 GND.n4837 GND.n1375 54.8683
R11444 GND.n5713 GND.n715 54.8683
R11445 GND.n3340 GND.n3339 54.358
R11446 GND.n1960 GND.n1959 54.358
R11447 GND.n1951 GND.n1950 52.4801
R11448 GND.n79 GND.t126 52.3082
R11449 GND.n116 GND.t147 52.3082
R11450 GND.n148 GND.t178 52.3082
R11451 GND.n185 GND.t137 52.3082
R11452 GND.n10 GND.t169 52.3082
R11453 GND.n47 GND.t167 52.3082
R11454 GND.n512 GND.t170 52.3082
R11455 GND.n475 GND.t150 52.3082
R11456 GND.n581 GND.t159 52.3082
R11457 GND.n544 GND.t141 52.3082
R11458 GND.n651 GND.t168 52.3082
R11459 GND.n614 GND.t172 52.3082
R11460 GND.n315 GND.t15 52.3082
R11461 GND.n283 GND.t10 52.3082
R11462 GND.n251 GND.t13 52.3082
R11463 GND.n220 GND.t1 52.3082
R11464 GND.n442 GND.t18 52.3082
R11465 GND.n410 GND.t3 52.3082
R11466 GND.n378 GND.t23 52.3082
R11467 GND.n347 GND.t21 52.3082
R11468 GND.n399 GND.n367 51.4173
R11469 GND.n463 GND.n462 50.455
R11470 GND.n431 GND.n430 50.455
R11471 GND.n399 GND.n398 50.455
R11472 GND.n4965 GND.n1223 47.2007
R11473 GND.n4959 GND.n1223 47.2007
R11474 GND.n4959 GND.n4958 47.2007
R11475 GND.n4958 GND.n4957 47.2007
R11476 GND.n4957 GND.n1230 47.2007
R11477 GND.n4951 GND.n1230 47.2007
R11478 GND.n4951 GND.n4950 47.2007
R11479 GND.n4950 GND.n4949 47.2007
R11480 GND.n4949 GND.n1238 47.2007
R11481 GND.n4943 GND.n1238 47.2007
R11482 GND.n4943 GND.n4942 47.2007
R11483 GND.n4942 GND.n4941 47.2007
R11484 GND.n4941 GND.n1246 47.2007
R11485 GND.n4935 GND.n1246 47.2007
R11486 GND.n4935 GND.n4934 47.2007
R11487 GND.n4934 GND.n4933 47.2007
R11488 GND.n4933 GND.n1254 47.2007
R11489 GND.n4927 GND.n1254 47.2007
R11490 GND.n4927 GND.n4926 47.2007
R11491 GND.n4926 GND.n4925 47.2007
R11492 GND.n4925 GND.n1262 47.2007
R11493 GND.n4919 GND.n1262 47.2007
R11494 GND.n4919 GND.n4918 47.2007
R11495 GND.n4918 GND.n4917 47.2007
R11496 GND.n4917 GND.n1270 47.2007
R11497 GND.n4911 GND.n1270 47.2007
R11498 GND.n4911 GND.n4910 47.2007
R11499 GND.n4910 GND.n4909 47.2007
R11500 GND.n4909 GND.n1278 47.2007
R11501 GND.n4903 GND.n1278 47.2007
R11502 GND.n4903 GND.n4902 47.2007
R11503 GND.n4902 GND.n4901 47.2007
R11504 GND.n4901 GND.n1286 47.2007
R11505 GND.n4895 GND.n1286 47.2007
R11506 GND.n4895 GND.n4894 47.2007
R11507 GND.n4894 GND.n4893 47.2007
R11508 GND.n4893 GND.n1294 47.2007
R11509 GND.n4887 GND.n1294 47.2007
R11510 GND.n4887 GND.n4886 47.2007
R11511 GND.n4886 GND.n4885 47.2007
R11512 GND.n4885 GND.n1302 47.2007
R11513 GND.n4879 GND.n1302 47.2007
R11514 GND.n4879 GND.n4878 47.2007
R11515 GND.n4878 GND.n4877 47.2007
R11516 GND.n4877 GND.n1310 47.2007
R11517 GND.n4871 GND.n1310 47.2007
R11518 GND.n4871 GND.n4870 47.2007
R11519 GND.n4870 GND.n4869 47.2007
R11520 GND.n4869 GND.n1318 47.2007
R11521 GND.n4863 GND.n1318 47.2007
R11522 GND.n4863 GND.n4862 47.2007
R11523 GND.n4862 GND.n4861 47.2007
R11524 GND.n4861 GND.n1326 47.2007
R11525 GND.n4855 GND.n1326 47.2007
R11526 GND.n4855 GND.n4854 47.2007
R11527 GND.n4854 GND.n4853 47.2007
R11528 GND.n4853 GND.n1334 47.2007
R11529 GND.n4847 GND.n1334 47.2007
R11530 GND.n4847 GND.n4846 47.2007
R11531 GND.n4846 GND.n4845 47.2007
R11532 GND.n4845 GND.n1342 47.2007
R11533 GND.n4839 GND.n1342 47.2007
R11534 GND.n4839 GND.n4838 47.2007
R11535 GND.n712 GND.n711 45.1884
R11536 GND.n768 GND.n767 45.1884
R11537 GND.n795 GND.n794 45.1884
R11538 GND.n1551 GND.n1550 45.1884
R11539 GND.n1577 GND.n1576 45.1884
R11540 GND.n1619 GND.n1618 45.1884
R11541 GND.n2822 GND.n2821 45.1884
R11542 GND.n2098 GND.n2097 45.1884
R11543 GND.n3254 GND.n3253 45.1884
R11544 GND.n2007 GND.n2006 45.1884
R11545 GND.n2119 GND.n2118 45.1884
R11546 GND.n1396 GND.n1395 45.1884
R11547 GND.n1416 GND.n1415 45.1884
R11548 GND.n4265 GND.n4264 45.1884
R11549 GND.n4374 GND.n1966 44.3322
R11550 GND.n3343 GND.n3342 44.3189
R11551 GND.n713 GND.n712 42.2793
R11552 GND.n5687 GND.n768 42.2793
R11553 GND.n797 GND.n795 42.2793
R11554 GND.n1578 GND.n1577 42.2793
R11555 GND.n1620 GND.n1619 42.2793
R11556 GND.n2869 GND.n2822 42.2793
R11557 GND.n2099 GND.n2098 42.2793
R11558 GND.n3255 GND.n3254 42.2793
R11559 GND.n2166 GND.n2119 42.2793
R11560 GND.n4805 GND.n1396 42.2793
R11561 GND.n1417 GND.n1416 42.2793
R11562 GND.n4266 GND.n4265 42.2793
R11563 GND.n3341 GND.n3340 41.6274
R11564 GND.n1961 GND.n1960 41.6274
R11565 GND.n3350 GND.n3349 40.8975
R11566 GND.n1964 GND.n1963 40.8975
R11567 GND.n101 GND.n99 38.8139
R11568 GND.n170 GND.n168 38.8139
R11569 GND.n32 GND.n30 38.8139
R11570 GND.n497 GND.n495 38.8139
R11571 GND.n566 GND.n564 38.8139
R11572 GND.n636 GND.n634 38.8139
R11573 GND.n137 GND.n136 37.8096
R11574 GND.n206 GND.n205 37.8096
R11575 GND.n68 GND.n67 37.8096
R11576 GND.n533 GND.n532 37.8096
R11577 GND.n602 GND.n601 37.8096
R11578 GND.n672 GND.n671 37.8096
R11579 GND.n4660 GND.n1551 36.9518
R11580 GND.n4312 GND.n2007 36.9518
R11581 GND.n3349 GND.n3348 35.055
R11582 GND.n3344 GND.n3343 35.055
R11583 GND.n1953 GND.n1952 35.055
R11584 GND.n1963 GND.n1949 35.055
R11585 GND.n3782 GND.n3781 33.8737
R11586 GND.n3476 GND.n3475 33.8737
R11587 GND.n2814 GND.n1375 33.0534
R11588 GND.n2910 GND.n2814 33.0534
R11589 GND.n2915 GND.n2811 33.0534
R11590 GND.n2915 GND.n2804 33.0534
R11591 GND.n2923 GND.n2804 33.0534
R11592 GND.n2923 GND.n2798 33.0534
R11593 GND.n2928 GND.n2798 33.0534
R11594 GND.n2928 GND.n2801 33.0534
R11595 GND.n2936 GND.n2772 33.0534
R11596 GND.n2944 GND.n2772 33.0534
R11597 GND.n1627 GND.n1527 33.0534
R11598 GND.n4557 GND.n1639 33.0534
R11599 GND.n4551 GND.n1639 33.0534
R11600 GND.n1668 GND.n1665 33.0534
R11601 GND.n3881 GND.n2109 33.0534
R11602 GND.n3904 GND.n3903 33.0534
R11603 GND.n3903 GND.n2011 33.0534
R11604 GND.n3919 GND.n2038 33.0534
R11605 GND.n5561 GND.n846 33.0534
R11606 GND.n5561 GND.n849 33.0534
R11607 GND.n5569 GND.n827 33.0534
R11608 GND.n5578 GND.n827 33.0534
R11609 GND.n5578 GND.n820 33.0534
R11610 GND.n5586 GND.n820 33.0534
R11611 GND.n5586 GND.n810 33.0534
R11612 GND.n5596 GND.n810 33.0534
R11613 GND.n5605 GND.n804 33.0534
R11614 GND.n5605 GND.n715 33.0534
R11615 GND.n2941 GND.n2790 31.7313
R11616 GND.n2954 GND.n2762 31.7313
R11617 GND.n2977 GND.n2755 31.7313
R11618 GND.n2981 GND.n2749 31.7313
R11619 GND.n2752 GND.n2738 31.7313
R11620 GND.n2991 GND.n2990 31.7313
R11621 GND.n2965 GND.n2961 31.7313
R11622 GND.n2962 GND.n2730 31.7313
R11623 GND.n3004 GND.n3003 31.7313
R11624 GND.n3101 GND.n2692 31.7313
R11625 GND.n3096 GND.n2699 31.7313
R11626 GND.n2706 GND.n2705 31.7313
R11627 GND.n3089 GND.n3088 31.7313
R11628 GND.n3083 GND.n2708 31.7313
R11629 GND.n3079 GND.n3021 31.7313
R11630 GND.n3111 GND.n2676 31.7313
R11631 GND.n3070 GND.n2677 31.7313
R11632 GND.n3126 GND.n2665 31.7313
R11633 GND.n3123 GND.n2667 31.7313
R11634 GND.n3136 GND.n2656 31.7313
R11635 GND.n3061 GND.n2657 31.7313
R11636 GND.n3151 GND.n2646 31.7313
R11637 GND.n3147 GND.n2648 31.7313
R11638 GND.n3161 GND.n2636 31.7313
R11639 GND.n3040 GND.n2638 31.7313
R11640 GND.n3177 GND.n2625 31.7313
R11641 GND.n2627 GND.n2619 31.7313
R11642 GND.n3186 GND.n3185 31.7313
R11643 GND.n3214 GND.n2604 31.7313
R11644 GND.n3217 GND.n2599 31.7313
R11645 GND.n3206 GND.n2601 31.7313
R11646 GND.n3230 GND.n2592 31.7313
R11647 GND.n4685 GND.n1525 31.7313
R11648 GND.n3918 GND.n2413 31.7313
R11649 GND.n3982 GND.n3977 31.7313
R11650 GND.n3992 GND.n2364 31.7313
R11651 GND.n2367 GND.n2355 31.7313
R11652 GND.n4001 GND.n2350 31.7313
R11653 GND.n4007 GND.n2352 31.7313
R11654 GND.n4004 GND.n2340 31.7313
R11655 GND.n4017 GND.n2341 31.7313
R11656 GND.n4026 GND.n2327 31.7313
R11657 GND.n4031 GND.n2330 31.7313
R11658 GND.n4028 GND.n2316 31.7313
R11659 GND.n4041 GND.n2317 31.7313
R11660 GND.n4050 GND.n2304 31.7313
R11661 GND.n4056 GND.n2306 31.7313
R11662 GND.n4053 GND.n2290 31.7313
R11663 GND.n4067 GND.n2291 31.7313
R11664 GND.n4144 GND.n2265 31.7313
R11665 GND.n4143 GND.n2267 31.7313
R11666 GND.n4075 GND.n2275 31.7313
R11667 GND.n4133 GND.n4132 31.7313
R11668 GND.n4127 GND.n4084 31.7313
R11669 GND.n4126 GND.n4090 31.7313
R11670 GND.n4104 GND.n4102 31.7313
R11671 GND.n4116 GND.n4115 31.7313
R11672 GND.n4160 GND.n2252 31.7313
R11673 GND.n4162 GND.n2247 31.7313
R11674 GND.n4165 GND.n2250 31.7313
R11675 GND.n2249 GND.n2239 31.7313
R11676 GND.n4175 GND.n2240 31.7313
R11677 GND.n5535 GND.n881 31.7313
R11678 GND.n5536 GND.n868 31.7313
R11679 GND.n5528 GND.n860 31.7313
R11680 GND.n5552 GND.n861 31.7313
R11681 GND.n3071 GND.t148 31.4007
R11682 GND.t118 GND.n2295 31.4007
R11683 GND.n2910 GND.t39 28.0955
R11684 GND.n3225 GND.t43 28.0955
R11685 GND.n3978 GND.t25 28.0955
R11686 GND.t63 GND.n804 28.0955
R11687 GND.n3313 GND.n3312 25.7944
R11688 GND.n3724 GND.n3723 25.7944
R11689 GND.n3319 GND.n3318 25.7944
R11690 GND.n2001 GND.n2000 25.7944
R11691 GND.n2801 GND.t136 22.807
R11692 GND.n3173 GND.t125 22.807
R11693 GND.n2344 GND.t140 22.807
R11694 GND.n5569 GND.t158 22.807
R11695 GND.n3080 GND.t131 22.1459
R11696 GND.n4136 GND.t120 22.1459
R11697 GND.n2766 GND.t127 21.4849
R11698 GND.n5544 GND.t133 21.4849
R11699 GND.n3354 GND.n3353 21.0737
R11700 GND.n4375 GND.n4374 21.0737
R11701 GND.t116 GND.n2694 20.8238
R11702 GND.n4113 GND.t145 20.8238
R11703 GND.n4583 GND.n1627 20.4933
R11704 GND.n4308 GND.n2038 20.4933
R11705 GND.n3062 GND.t129 20.1628
R11706 GND.t122 GND.n2308 20.1628
R11707 GND.n3337 GND.t115 19.8005
R11708 GND.n3337 GND.t30 19.8005
R11709 GND.n3338 GND.t95 19.8005
R11710 GND.n3338 GND.t71 19.8005
R11711 GND.n1957 GND.t80 19.8005
R11712 GND.n1957 GND.t98 19.8005
R11713 GND.n1958 GND.t51 19.8005
R11714 GND.n1958 GND.t33 19.8005
R11715 GND.n3334 GND.n3333 19.5087
R11716 GND.n3347 GND.n3334 19.5087
R11717 GND.n3345 GND.n3336 19.5087
R11718 GND.n1962 GND.n1956 19.5087
R11719 GND.n5650 GND.n5607 19.3944
R11720 GND.n5646 GND.n5607 19.3944
R11721 GND.n5646 GND.n5645 19.3944
R11722 GND.n5645 GND.n5644 19.3944
R11723 GND.n5644 GND.n5613 19.3944
R11724 GND.n5640 GND.n5613 19.3944
R11725 GND.n5640 GND.n5639 19.3944
R11726 GND.n5639 GND.n5638 19.3944
R11727 GND.n5638 GND.n5619 19.3944
R11728 GND.n5634 GND.n5619 19.3944
R11729 GND.n5634 GND.n5633 19.3944
R11730 GND.n5633 GND.n5632 19.3944
R11731 GND.n5632 GND.n5625 19.3944
R11732 GND.n5628 GND.n5625 19.3944
R11733 GND.n3980 GND.n2114 19.3944
R11734 GND.n3980 GND.n2173 19.3944
R11735 GND.n2174 GND.n2173 19.3944
R11736 GND.n2175 GND.n2174 19.3944
R11737 GND.n2354 GND.n2175 19.3944
R11738 GND.n2354 GND.n2181 19.3944
R11739 GND.n2182 GND.n2181 19.3944
R11740 GND.n2183 GND.n2182 19.3944
R11741 GND.n2331 GND.n2183 19.3944
R11742 GND.n2331 GND.n2189 19.3944
R11743 GND.n2190 GND.n2189 19.3944
R11744 GND.n2191 GND.n2190 19.3944
R11745 GND.n2318 GND.n2191 19.3944
R11746 GND.n2318 GND.n2197 19.3944
R11747 GND.n2198 GND.n2197 19.3944
R11748 GND.n2199 GND.n2198 19.3944
R11749 GND.n4052 GND.n2199 19.3944
R11750 GND.n4052 GND.n2205 19.3944
R11751 GND.n2206 GND.n2205 19.3944
R11752 GND.n2207 GND.n2206 19.3944
R11753 GND.n2268 GND.n2207 19.3944
R11754 GND.n2268 GND.n2213 19.3944
R11755 GND.n2214 GND.n2213 19.3944
R11756 GND.n2215 GND.n2214 19.3944
R11757 GND.n2279 GND.n2215 19.3944
R11758 GND.n2279 GND.n2221 19.3944
R11759 GND.n2222 GND.n2221 19.3944
R11760 GND.n2223 GND.n2222 19.3944
R11761 GND.n4106 GND.n2223 19.3944
R11762 GND.n4106 GND.n2229 19.3944
R11763 GND.n2230 GND.n2229 19.3944
R11764 GND.n2231 GND.n2230 19.3944
R11765 GND.n2237 GND.n2231 19.3944
R11766 GND.n2237 GND.n2236 19.3944
R11767 GND.n4178 GND.n2236 19.3944
R11768 GND.n4178 GND.n873 19.3944
R11769 GND.n5542 GND.n873 19.3944
R11770 GND.n5542 GND.n874 19.3944
R11771 GND.n876 GND.n874 19.3944
R11772 GND.n876 GND.n852 19.3944
R11773 GND.n5559 GND.n852 19.3944
R11774 GND.n5559 GND.n853 19.3944
R11775 GND.n855 GND.n853 19.3944
R11776 GND.n855 GND.n832 19.3944
R11777 GND.n5576 GND.n832 19.3944
R11778 GND.n5576 GND.n833 19.3944
R11779 GND.n835 GND.n833 19.3944
R11780 GND.n835 GND.n814 19.3944
R11781 GND.n5594 GND.n814 19.3944
R11782 GND.n5594 GND.n815 19.3944
R11783 GND.n815 GND.n802 19.3944
R11784 GND.n5653 GND.n802 19.3944
R11785 GND.n4231 GND.n4230 19.3944
R11786 GND.n4230 GND.n4229 19.3944
R11787 GND.n4229 GND.n2172 19.3944
R11788 GND.n4225 GND.n2172 19.3944
R11789 GND.n4225 GND.n4224 19.3944
R11790 GND.n4224 GND.n4223 19.3944
R11791 GND.n4223 GND.n2180 19.3944
R11792 GND.n4219 GND.n2180 19.3944
R11793 GND.n4219 GND.n4218 19.3944
R11794 GND.n4218 GND.n4217 19.3944
R11795 GND.n4217 GND.n2188 19.3944
R11796 GND.n4213 GND.n2188 19.3944
R11797 GND.n4213 GND.n4212 19.3944
R11798 GND.n4212 GND.n4211 19.3944
R11799 GND.n4211 GND.n2196 19.3944
R11800 GND.n4207 GND.n2196 19.3944
R11801 GND.n4207 GND.n4206 19.3944
R11802 GND.n4206 GND.n4205 19.3944
R11803 GND.n4205 GND.n2204 19.3944
R11804 GND.n4201 GND.n2204 19.3944
R11805 GND.n4201 GND.n4200 19.3944
R11806 GND.n4200 GND.n4199 19.3944
R11807 GND.n4199 GND.n2212 19.3944
R11808 GND.n4195 GND.n2212 19.3944
R11809 GND.n4195 GND.n4194 19.3944
R11810 GND.n4194 GND.n4193 19.3944
R11811 GND.n4193 GND.n2220 19.3944
R11812 GND.n4189 GND.n2220 19.3944
R11813 GND.n4189 GND.n4188 19.3944
R11814 GND.n4188 GND.n4187 19.3944
R11815 GND.n4187 GND.n2228 19.3944
R11816 GND.n4183 GND.n2228 19.3944
R11817 GND.n4183 GND.n4182 19.3944
R11818 GND.n4182 GND.n4181 19.3944
R11819 GND.n4181 GND.n879 19.3944
R11820 GND.n5538 GND.n879 19.3944
R11821 GND.n5540 GND.n5538 19.3944
R11822 GND.n5540 GND.n5539 19.3944
R11823 GND.n5539 GND.n858 19.3944
R11824 GND.n5555 GND.n858 19.3944
R11825 GND.n5557 GND.n5555 19.3944
R11826 GND.n5557 GND.n5556 19.3944
R11827 GND.n5556 GND.n838 19.3944
R11828 GND.n5572 GND.n838 19.3944
R11829 GND.n5574 GND.n5572 19.3944
R11830 GND.n5574 GND.n5573 19.3944
R11831 GND.n5573 GND.n818 19.3944
R11832 GND.n5589 GND.n818 19.3944
R11833 GND.n5592 GND.n5589 19.3944
R11834 GND.n5592 GND.n5591 19.3944
R11835 GND.n5591 GND.n800 19.3944
R11836 GND.n5655 GND.n800 19.3944
R11837 GND.n5711 GND.n744 19.3944
R11838 GND.n5707 GND.n744 19.3944
R11839 GND.n5707 GND.n5706 19.3944
R11840 GND.n5706 GND.n5705 19.3944
R11841 GND.n5705 GND.n751 19.3944
R11842 GND.n5701 GND.n751 19.3944
R11843 GND.n5701 GND.n5700 19.3944
R11844 GND.n5700 GND.n5699 19.3944
R11845 GND.n5699 GND.n757 19.3944
R11846 GND.n5695 GND.n757 19.3944
R11847 GND.n5695 GND.n5694 19.3944
R11848 GND.n5694 GND.n5693 19.3944
R11849 GND.n5693 GND.n763 19.3944
R11850 GND.n5689 GND.n763 19.3944
R11851 GND.n5689 GND.n5688 19.3944
R11852 GND.n5686 GND.n771 19.3944
R11853 GND.n5682 GND.n771 19.3944
R11854 GND.n5682 GND.n5681 19.3944
R11855 GND.n5681 GND.n5680 19.3944
R11856 GND.n5680 GND.n777 19.3944
R11857 GND.n5676 GND.n777 19.3944
R11858 GND.n5676 GND.n5675 19.3944
R11859 GND.n5675 GND.n5674 19.3944
R11860 GND.n5674 GND.n783 19.3944
R11861 GND.n5670 GND.n783 19.3944
R11862 GND.n5670 GND.n5669 19.3944
R11863 GND.n5669 GND.n5668 19.3944
R11864 GND.n5668 GND.n789 19.3944
R11865 GND.n5664 GND.n789 19.3944
R11866 GND.n5664 GND.n5663 19.3944
R11867 GND.n5663 GND.n5662 19.3944
R11868 GND.n4765 GND.n1420 19.3944
R11869 GND.n4761 GND.n1420 19.3944
R11870 GND.n4761 GND.n4760 19.3944
R11871 GND.n4760 GND.n4759 19.3944
R11872 GND.n4759 GND.n1428 19.3944
R11873 GND.n4755 GND.n1428 19.3944
R11874 GND.n4755 GND.n4754 19.3944
R11875 GND.n4754 GND.n4753 19.3944
R11876 GND.n4753 GND.n1436 19.3944
R11877 GND.n4749 GND.n1436 19.3944
R11878 GND.n4749 GND.n4748 19.3944
R11879 GND.n4748 GND.n4747 19.3944
R11880 GND.n4747 GND.n1444 19.3944
R11881 GND.n4743 GND.n1444 19.3944
R11882 GND.n4743 GND.n4742 19.3944
R11883 GND.n4742 GND.n4741 19.3944
R11884 GND.n4741 GND.n1452 19.3944
R11885 GND.n4737 GND.n1452 19.3944
R11886 GND.n4737 GND.n4736 19.3944
R11887 GND.n4736 GND.n4735 19.3944
R11888 GND.n4735 GND.n1460 19.3944
R11889 GND.n4731 GND.n1460 19.3944
R11890 GND.n4731 GND.n4730 19.3944
R11891 GND.n4730 GND.n4729 19.3944
R11892 GND.n4729 GND.n1468 19.3944
R11893 GND.n4725 GND.n1468 19.3944
R11894 GND.n4725 GND.n4724 19.3944
R11895 GND.n4724 GND.n4723 19.3944
R11896 GND.n4723 GND.n1476 19.3944
R11897 GND.n4719 GND.n1476 19.3944
R11898 GND.n4719 GND.n4718 19.3944
R11899 GND.n4718 GND.n4717 19.3944
R11900 GND.n4717 GND.n1484 19.3944
R11901 GND.n4713 GND.n1484 19.3944
R11902 GND.n4713 GND.n4712 19.3944
R11903 GND.n4712 GND.n4711 19.3944
R11904 GND.n4711 GND.n1492 19.3944
R11905 GND.n4707 GND.n1492 19.3944
R11906 GND.n4707 GND.n4706 19.3944
R11907 GND.n4706 GND.n4705 19.3944
R11908 GND.n4705 GND.n1500 19.3944
R11909 GND.n4701 GND.n1500 19.3944
R11910 GND.n4701 GND.n4700 19.3944
R11911 GND.n4700 GND.n4699 19.3944
R11912 GND.n4699 GND.n1508 19.3944
R11913 GND.n4695 GND.n1508 19.3944
R11914 GND.n4695 GND.n4694 19.3944
R11915 GND.n4694 GND.n4693 19.3944
R11916 GND.n4693 GND.n1516 19.3944
R11917 GND.n4689 GND.n1516 19.3944
R11918 GND.n4689 GND.n4688 19.3944
R11919 GND.n4688 GND.n4687 19.3944
R11920 GND.n4680 GND.n4679 19.3944
R11921 GND.n4679 GND.n4678 19.3944
R11922 GND.n4678 GND.n1536 19.3944
R11923 GND.n4674 GND.n1536 19.3944
R11924 GND.n4674 GND.n4673 19.3944
R11925 GND.n4673 GND.n4672 19.3944
R11926 GND.n4672 GND.n1541 19.3944
R11927 GND.n4668 GND.n1541 19.3944
R11928 GND.n4668 GND.n4667 19.3944
R11929 GND.n4667 GND.n4666 19.3944
R11930 GND.n4666 GND.n1546 19.3944
R11931 GND.n4662 GND.n1546 19.3944
R11932 GND.n4662 GND.n4661 19.3944
R11933 GND.n4659 GND.n1556 19.3944
R11934 GND.n4655 GND.n1556 19.3944
R11935 GND.n4655 GND.n4654 19.3944
R11936 GND.n4654 GND.n4653 19.3944
R11937 GND.n4653 GND.n1561 19.3944
R11938 GND.n4649 GND.n1561 19.3944
R11939 GND.n4649 GND.n4648 19.3944
R11940 GND.n4648 GND.n4647 19.3944
R11941 GND.n4647 GND.n1566 19.3944
R11942 GND.n4643 GND.n1566 19.3944
R11943 GND.n4643 GND.n4642 19.3944
R11944 GND.n4642 GND.n4641 19.3944
R11945 GND.n4641 GND.n1571 19.3944
R11946 GND.n4637 GND.n1571 19.3944
R11947 GND.n4637 GND.n4636 19.3944
R11948 GND.n4636 GND.n4635 19.3944
R11949 GND.n2873 GND.n2817 19.3944
R11950 GND.n2900 GND.n2817 19.3944
R11951 GND.n2900 GND.n2818 19.3944
R11952 GND.n2896 GND.n2818 19.3944
R11953 GND.n2896 GND.n2895 19.3944
R11954 GND.n2895 GND.n2894 19.3944
R11955 GND.n2894 GND.n2879 19.3944
R11956 GND.n2890 GND.n2879 19.3944
R11957 GND.n2890 GND.n2889 19.3944
R11958 GND.n2889 GND.n2888 19.3944
R11959 GND.n2888 GND.n2883 19.3944
R11960 GND.n2884 GND.n2883 19.3944
R11961 GND.n2884 GND.n2760 19.3944
R11962 GND.n2956 GND.n2760 19.3944
R11963 GND.n2956 GND.n2757 19.3944
R11964 GND.n2975 GND.n2757 19.3944
R11965 GND.n2975 GND.n2758 19.3944
R11966 GND.n2971 GND.n2758 19.3944
R11967 GND.n2971 GND.n2970 19.3944
R11968 GND.n2970 GND.n2969 19.3944
R11969 GND.n2969 GND.n2727 19.3944
R11970 GND.n3006 GND.n2727 19.3944
R11971 GND.n3007 GND.n3006 19.3944
R11972 GND.n3007 GND.n2725 19.3944
R11973 GND.n3011 GND.n2725 19.3944
R11974 GND.n3014 GND.n3011 19.3944
R11975 GND.n3015 GND.n3014 19.3944
R11976 GND.n3015 GND.n2723 19.3944
R11977 GND.n3019 GND.n2723 19.3944
R11978 GND.n3019 GND.n2674 19.3944
R11979 GND.n3113 GND.n2674 19.3944
R11980 GND.n3113 GND.n2671 19.3944
R11981 GND.n3118 GND.n2671 19.3944
R11982 GND.n3118 GND.n2672 19.3944
R11983 GND.n2672 GND.n2654 19.3944
R11984 GND.n3138 GND.n2654 19.3944
R11985 GND.n3138 GND.n2651 19.3944
R11986 GND.n3143 GND.n2651 19.3944
R11987 GND.n3143 GND.n2652 19.3944
R11988 GND.n2652 GND.n2634 19.3944
R11989 GND.n3163 GND.n2634 19.3944
R11990 GND.n3163 GND.n2631 19.3944
R11991 GND.n3171 GND.n2631 19.3944
R11992 GND.n3171 GND.n2632 19.3944
R11993 GND.n3167 GND.n2632 19.3944
R11994 GND.n3167 GND.n2606 19.3944
R11995 GND.n3212 GND.n2606 19.3944
R11996 GND.n3212 GND.n2607 19.3944
R11997 GND.n3208 GND.n2607 19.3944
R11998 GND.n3208 GND.n2590 19.3944
R11999 GND.n3232 GND.n2590 19.3944
R12000 GND.n3233 GND.n3232 19.3944
R12001 GND.n4627 GND.n4626 19.3944
R12002 GND.n4626 GND.n4625 19.3944
R12003 GND.n4625 GND.n1584 19.3944
R12004 GND.n4618 GND.n1584 19.3944
R12005 GND.n4618 GND.n4617 19.3944
R12006 GND.n4617 GND.n1594 19.3944
R12007 GND.n4610 GND.n1594 19.3944
R12008 GND.n4610 GND.n4609 19.3944
R12009 GND.n4609 GND.n1602 19.3944
R12010 GND.n4602 GND.n1602 19.3944
R12011 GND.n4602 GND.n4601 19.3944
R12012 GND.n4601 GND.n1610 19.3944
R12013 GND.n4594 GND.n1610 19.3944
R12014 GND.n4594 GND.n4593 19.3944
R12015 GND.n2840 GND.n2835 19.3944
R12016 GND.n2844 GND.n2835 19.3944
R12017 GND.n2845 GND.n2844 19.3944
R12018 GND.n2848 GND.n2845 19.3944
R12019 GND.n2848 GND.n2831 19.3944
R12020 GND.n2852 GND.n2831 19.3944
R12021 GND.n2853 GND.n2852 19.3944
R12022 GND.n2856 GND.n2853 19.3944
R12023 GND.n2856 GND.n2827 19.3944
R12024 GND.n2860 GND.n2827 19.3944
R12025 GND.n2861 GND.n2860 19.3944
R12026 GND.n2864 GND.n2861 19.3944
R12027 GND.n2864 GND.n2823 19.3944
R12028 GND.n2868 GND.n2823 19.3944
R12029 GND.n1422 GND.n1421 19.3944
R12030 GND.n1423 GND.n1422 19.3944
R12031 GND.n2912 GND.n1423 19.3944
R12032 GND.n2912 GND.n1429 19.3944
R12033 GND.n1430 GND.n1429 19.3944
R12034 GND.n1431 GND.n1430 19.3944
R12035 GND.n2925 GND.n1431 19.3944
R12036 GND.n2925 GND.n1437 19.3944
R12037 GND.n1438 GND.n1437 19.3944
R12038 GND.n1439 GND.n1438 19.3944
R12039 GND.n2938 GND.n1439 19.3944
R12040 GND.n2938 GND.n1445 19.3944
R12041 GND.n1446 GND.n1445 19.3944
R12042 GND.n1447 GND.n1446 19.3944
R12043 GND.n2753 GND.n1447 19.3944
R12044 GND.n2753 GND.n1453 19.3944
R12045 GND.n1454 GND.n1453 19.3944
R12046 GND.n1455 GND.n1454 19.3944
R12047 GND.n2740 GND.n1455 19.3944
R12048 GND.n2740 GND.n1461 19.3944
R12049 GND.n1462 GND.n1461 19.3944
R12050 GND.n1463 GND.n1462 19.3944
R12051 GND.n3099 GND.n1463 19.3944
R12052 GND.n3099 GND.n1469 19.3944
R12053 GND.n1470 GND.n1469 19.3944
R12054 GND.n1471 GND.n1470 19.3944
R12055 GND.n2710 GND.n1471 19.3944
R12056 GND.n2710 GND.n1477 19.3944
R12057 GND.n1478 GND.n1477 19.3944
R12058 GND.n1479 GND.n1478 19.3944
R12059 GND.n2678 GND.n1479 19.3944
R12060 GND.n2678 GND.n1485 19.3944
R12061 GND.n1486 GND.n1485 19.3944
R12062 GND.n1487 GND.n1486 19.3944
R12063 GND.n3122 GND.n1487 19.3944
R12064 GND.n3122 GND.n1493 19.3944
R12065 GND.n1494 GND.n1493 19.3944
R12066 GND.n1495 GND.n1494 19.3944
R12067 GND.n3149 GND.n1495 19.3944
R12068 GND.n3149 GND.n1501 19.3944
R12069 GND.n1502 GND.n1501 19.3944
R12070 GND.n1503 GND.n1502 19.3944
R12071 GND.n2629 GND.n1503 19.3944
R12072 GND.n2629 GND.n1509 19.3944
R12073 GND.n1510 GND.n1509 19.3944
R12074 GND.n1511 GND.n1510 19.3944
R12075 GND.n2603 GND.n1511 19.3944
R12076 GND.n2603 GND.n1517 19.3944
R12077 GND.n1518 GND.n1517 19.3944
R12078 GND.n1519 GND.n1518 19.3944
R12079 GND.n3228 GND.n1519 19.3944
R12080 GND.n3228 GND.n3227 19.3944
R12081 GND.n3269 GND.n3268 19.3944
R12082 GND.n3274 GND.n3269 19.3944
R12083 GND.n3274 GND.n2580 19.3944
R12084 GND.n3278 GND.n2580 19.3944
R12085 GND.n3279 GND.n3278 19.3944
R12086 GND.n3282 GND.n3279 19.3944
R12087 GND.n3282 GND.n2578 19.3944
R12088 GND.n3286 GND.n2578 19.3944
R12089 GND.n3289 GND.n3286 19.3944
R12090 GND.n3290 GND.n3289 19.3944
R12091 GND.n3290 GND.n2572 19.3944
R12092 GND.n3294 GND.n2572 19.3944
R12093 GND.n3295 GND.n3294 19.3944
R12094 GND.n3482 GND.n3295 19.3944
R12095 GND.n3482 GND.n2570 19.3944
R12096 GND.n3486 GND.n2570 19.3944
R12097 GND.n3486 GND.n2564 19.3944
R12098 GND.n3513 GND.n2564 19.3944
R12099 GND.n3513 GND.n2565 19.3944
R12100 GND.n3509 GND.n2565 19.3944
R12101 GND.n3509 GND.n3508 19.3944
R12102 GND.n3508 GND.n3507 19.3944
R12103 GND.n3507 GND.n2535 19.3944
R12104 GND.n3551 GND.n2535 19.3944
R12105 GND.n3551 GND.n2532 19.3944
R12106 GND.n3566 GND.n2532 19.3944
R12107 GND.n3566 GND.n2533 19.3944
R12108 GND.n3562 GND.n2533 19.3944
R12109 GND.n3562 GND.n3561 19.3944
R12110 GND.n3561 GND.n3560 19.3944
R12111 GND.n3560 GND.n2519 19.3944
R12112 GND.n3614 GND.n2519 19.3944
R12113 GND.n3614 GND.n2516 19.3944
R12114 GND.n3620 GND.n2516 19.3944
R12115 GND.n3620 GND.n2517 19.3944
R12116 GND.n2517 GND.n2506 19.3944
R12117 GND.n2506 GND.n2505 19.3944
R12118 GND.n3651 GND.n2505 19.3944
R12119 GND.n3651 GND.n2502 19.3944
R12120 GND.n3659 GND.n2502 19.3944
R12121 GND.n3659 GND.n2503 19.3944
R12122 GND.n3655 GND.n2503 19.3944
R12123 GND.n3655 GND.n2487 19.3944
R12124 GND.n3687 GND.n2487 19.3944
R12125 GND.n3687 GND.n2484 19.3944
R12126 GND.n3704 GND.n2484 19.3944
R12127 GND.n3704 GND.n2485 19.3944
R12128 GND.n3700 GND.n2485 19.3944
R12129 GND.n3700 GND.n3699 19.3944
R12130 GND.n3699 GND.n3698 19.3944
R12131 GND.n3698 GND.n3695 19.3944
R12132 GND.n3695 GND.n2476 19.3944
R12133 GND.n3808 GND.n2476 19.3944
R12134 GND.n3808 GND.n2473 19.3944
R12135 GND.n3813 GND.n2473 19.3944
R12136 GND.n3813 GND.n2474 19.3944
R12137 GND.n2474 GND.n2449 19.3944
R12138 GND.n3840 GND.n2449 19.3944
R12139 GND.n3840 GND.n2446 19.3944
R12140 GND.n3850 GND.n2446 19.3944
R12141 GND.n3850 GND.n2447 19.3944
R12142 GND.n3846 GND.n2447 19.3944
R12143 GND.n3846 GND.n3845 19.3944
R12144 GND.n3845 GND.n2105 19.3944
R12145 GND.n4240 GND.n2105 19.3944
R12146 GND.n4302 GND.n4301 19.3944
R12147 GND.n4301 GND.n2046 19.3944
R12148 GND.n4294 GND.n2046 19.3944
R12149 GND.n4294 GND.n4293 19.3944
R12150 GND.n4293 GND.n2056 19.3944
R12151 GND.n4286 GND.n2056 19.3944
R12152 GND.n4286 GND.n4285 19.3944
R12153 GND.n4285 GND.n2064 19.3944
R12154 GND.n4278 GND.n2064 19.3944
R12155 GND.n4278 GND.n4277 19.3944
R12156 GND.n4277 GND.n2074 19.3944
R12157 GND.n4270 GND.n2074 19.3944
R12158 GND.n4270 GND.n4269 19.3944
R12159 GND.n4269 GND.n2082 19.3944
R12160 GND.n4258 GND.n2082 19.3944
R12161 GND.n4258 GND.n4257 19.3944
R12162 GND.n4257 GND.n4256 19.3944
R12163 GND.n4256 GND.n2089 19.3944
R12164 GND.n4252 GND.n2089 19.3944
R12165 GND.n4252 GND.n4251 19.3944
R12166 GND.n4251 GND.n4250 19.3944
R12167 GND.n4250 GND.n2095 19.3944
R12168 GND.n4246 GND.n4245 19.3944
R12169 GND.n4245 GND.n4244 19.3944
R12170 GND.n4244 GND.n2103 19.3944
R12171 GND.n3260 GND.n2585 19.3944
R12172 GND.n3263 GND.n3260 19.3944
R12173 GND.n3265 GND.n3263 19.3944
R12174 GND.n4622 GND.n1587 19.3944
R12175 GND.n4622 GND.n4621 19.3944
R12176 GND.n4621 GND.n1590 19.3944
R12177 GND.n4614 GND.n1590 19.3944
R12178 GND.n4614 GND.n4613 19.3944
R12179 GND.n4613 GND.n1598 19.3944
R12180 GND.n4606 GND.n1598 19.3944
R12181 GND.n4606 GND.n4605 19.3944
R12182 GND.n4605 GND.n1606 19.3944
R12183 GND.n4598 GND.n1606 19.3944
R12184 GND.n4598 GND.n4597 19.3944
R12185 GND.n4597 GND.n1614 19.3944
R12186 GND.n4590 GND.n1614 19.3944
R12187 GND.n4590 GND.n4589 19.3944
R12188 GND.n4589 GND.n1624 19.3944
R12189 GND.n3237 GND.n1624 19.3944
R12190 GND.n3240 GND.n3237 19.3944
R12191 GND.n3243 GND.n3240 19.3944
R12192 GND.n3243 GND.n2587 19.3944
R12193 GND.n3247 GND.n2587 19.3944
R12194 GND.n3250 GND.n3247 19.3944
R12195 GND.n3256 GND.n3250 19.3944
R12196 GND.n1686 GND.n1667 19.3944
R12197 GND.n1686 GND.n1685 19.3944
R12198 GND.n4536 GND.n1685 19.3944
R12199 GND.n4536 GND.n4535 19.3944
R12200 GND.n4535 GND.n4534 19.3944
R12201 GND.n4534 GND.n1692 19.3944
R12202 GND.n1713 GND.n1692 19.3944
R12203 GND.n4522 GND.n1713 19.3944
R12204 GND.n4522 GND.n4521 19.3944
R12205 GND.n4521 GND.n4520 19.3944
R12206 GND.n4520 GND.n1719 19.3944
R12207 GND.n1738 GND.n1719 19.3944
R12208 GND.n4508 GND.n1738 19.3944
R12209 GND.n4508 GND.n4507 19.3944
R12210 GND.n4507 GND.n4506 19.3944
R12211 GND.n4506 GND.n1744 19.3944
R12212 GND.n4494 GND.n1744 19.3944
R12213 GND.n4494 GND.n4493 19.3944
R12214 GND.n4493 GND.n4492 19.3944
R12215 GND.n4492 GND.n1764 19.3944
R12216 GND.n4480 GND.n1764 19.3944
R12217 GND.n4480 GND.n4479 19.3944
R12218 GND.n4479 GND.n4478 19.3944
R12219 GND.n4478 GND.n1784 19.3944
R12220 GND.n4466 GND.n1784 19.3944
R12221 GND.n4466 GND.n4465 19.3944
R12222 GND.n4465 GND.n4464 19.3944
R12223 GND.n4464 GND.n1804 19.3944
R12224 GND.n4452 GND.n1804 19.3944
R12225 GND.n4452 GND.n4451 19.3944
R12226 GND.n4451 GND.n4450 19.3944
R12227 GND.n4450 GND.n1822 19.3944
R12228 GND.n4438 GND.n1822 19.3944
R12229 GND.n4438 GND.n4437 19.3944
R12230 GND.n4437 GND.n4436 19.3944
R12231 GND.n4436 GND.n1842 19.3944
R12232 GND.n1871 GND.n1842 19.3944
R12233 GND.n1871 GND.n1868 19.3944
R12234 GND.n4417 GND.n1868 19.3944
R12235 GND.n4417 GND.n4416 19.3944
R12236 GND.n4416 GND.n4415 19.3944
R12237 GND.n4415 GND.n1877 19.3944
R12238 GND.n2493 GND.n1877 19.3944
R12239 GND.n2493 GND.n1911 19.3944
R12240 GND.n4397 GND.n1911 19.3944
R12241 GND.n4397 GND.n4396 19.3944
R12242 GND.n4396 GND.n4395 19.3944
R12243 GND.n4395 GND.n1915 19.3944
R12244 GND.n3794 GND.n1915 19.3944
R12245 GND.n3794 GND.n3791 19.3944
R12246 GND.n3798 GND.n3791 19.3944
R12247 GND.n3798 GND.n3789 19.3944
R12248 GND.n3804 GND.n3789 19.3944
R12249 GND.n3804 GND.n3803 19.3944
R12250 GND.n3803 GND.n2457 19.3944
R12251 GND.n3830 GND.n2457 19.3944
R12252 GND.n3830 GND.n2455 19.3944
R12253 GND.n3836 GND.n2455 19.3944
R12254 GND.n3836 GND.n3835 19.3944
R12255 GND.n3835 GND.n2433 19.3944
R12256 GND.n3864 GND.n2433 19.3944
R12257 GND.n3864 GND.n2431 19.3944
R12258 GND.n3868 GND.n2431 19.3944
R12259 GND.n3868 GND.n2111 19.3944
R12260 GND.n4236 GND.n2111 19.3944
R12261 GND.n5364 GND.n982 19.3944
R12262 GND.n5370 GND.n982 19.3944
R12263 GND.n5370 GND.n980 19.3944
R12264 GND.n5374 GND.n980 19.3944
R12265 GND.n5374 GND.n976 19.3944
R12266 GND.n5380 GND.n976 19.3944
R12267 GND.n5380 GND.n974 19.3944
R12268 GND.n5384 GND.n974 19.3944
R12269 GND.n5384 GND.n970 19.3944
R12270 GND.n5390 GND.n970 19.3944
R12271 GND.n5390 GND.n968 19.3944
R12272 GND.n5394 GND.n968 19.3944
R12273 GND.n5394 GND.n964 19.3944
R12274 GND.n5400 GND.n964 19.3944
R12275 GND.n5400 GND.n962 19.3944
R12276 GND.n5404 GND.n962 19.3944
R12277 GND.n5404 GND.n958 19.3944
R12278 GND.n5410 GND.n958 19.3944
R12279 GND.n5410 GND.n956 19.3944
R12280 GND.n5414 GND.n956 19.3944
R12281 GND.n5414 GND.n952 19.3944
R12282 GND.n5420 GND.n952 19.3944
R12283 GND.n5420 GND.n950 19.3944
R12284 GND.n5424 GND.n950 19.3944
R12285 GND.n5424 GND.n946 19.3944
R12286 GND.n5430 GND.n946 19.3944
R12287 GND.n5430 GND.n944 19.3944
R12288 GND.n5434 GND.n944 19.3944
R12289 GND.n5434 GND.n940 19.3944
R12290 GND.n5440 GND.n940 19.3944
R12291 GND.n5440 GND.n938 19.3944
R12292 GND.n5444 GND.n938 19.3944
R12293 GND.n5444 GND.n934 19.3944
R12294 GND.n5450 GND.n934 19.3944
R12295 GND.n5450 GND.n932 19.3944
R12296 GND.n5454 GND.n932 19.3944
R12297 GND.n5454 GND.n928 19.3944
R12298 GND.n5460 GND.n928 19.3944
R12299 GND.n5460 GND.n926 19.3944
R12300 GND.n5464 GND.n926 19.3944
R12301 GND.n5464 GND.n922 19.3944
R12302 GND.n5470 GND.n922 19.3944
R12303 GND.n5470 GND.n920 19.3944
R12304 GND.n5474 GND.n920 19.3944
R12305 GND.n5474 GND.n916 19.3944
R12306 GND.n5480 GND.n916 19.3944
R12307 GND.n5480 GND.n914 19.3944
R12308 GND.n5484 GND.n914 19.3944
R12309 GND.n5484 GND.n910 19.3944
R12310 GND.n5490 GND.n910 19.3944
R12311 GND.n5490 GND.n908 19.3944
R12312 GND.n5494 GND.n908 19.3944
R12313 GND.n5494 GND.n904 19.3944
R12314 GND.n5500 GND.n904 19.3944
R12315 GND.n5500 GND.n902 19.3944
R12316 GND.n5504 GND.n902 19.3944
R12317 GND.n5504 GND.n898 19.3944
R12318 GND.n5510 GND.n898 19.3944
R12319 GND.n5510 GND.n896 19.3944
R12320 GND.n5515 GND.n896 19.3944
R12321 GND.n5515 GND.n892 19.3944
R12322 GND.n5521 GND.n892 19.3944
R12323 GND.n5522 GND.n5521 19.3944
R12324 GND.n4969 GND.n1221 19.3944
R12325 GND.n4969 GND.n1219 19.3944
R12326 GND.n4973 GND.n1219 19.3944
R12327 GND.n4973 GND.n1215 19.3944
R12328 GND.n4979 GND.n1215 19.3944
R12329 GND.n4979 GND.n1213 19.3944
R12330 GND.n4983 GND.n1213 19.3944
R12331 GND.n4983 GND.n1209 19.3944
R12332 GND.n4989 GND.n1209 19.3944
R12333 GND.n4989 GND.n1207 19.3944
R12334 GND.n4993 GND.n1207 19.3944
R12335 GND.n4993 GND.n1203 19.3944
R12336 GND.n4999 GND.n1203 19.3944
R12337 GND.n4999 GND.n1201 19.3944
R12338 GND.n5003 GND.n1201 19.3944
R12339 GND.n5003 GND.n1197 19.3944
R12340 GND.n5009 GND.n1197 19.3944
R12341 GND.n5009 GND.n1195 19.3944
R12342 GND.n5013 GND.n1195 19.3944
R12343 GND.n5013 GND.n1191 19.3944
R12344 GND.n5019 GND.n1191 19.3944
R12345 GND.n5019 GND.n1189 19.3944
R12346 GND.n5023 GND.n1189 19.3944
R12347 GND.n5023 GND.n1185 19.3944
R12348 GND.n5029 GND.n1185 19.3944
R12349 GND.n5029 GND.n1183 19.3944
R12350 GND.n5033 GND.n1183 19.3944
R12351 GND.n5033 GND.n1179 19.3944
R12352 GND.n5039 GND.n1179 19.3944
R12353 GND.n5039 GND.n1177 19.3944
R12354 GND.n5043 GND.n1177 19.3944
R12355 GND.n5043 GND.n1173 19.3944
R12356 GND.n5049 GND.n1173 19.3944
R12357 GND.n5049 GND.n1171 19.3944
R12358 GND.n5053 GND.n1171 19.3944
R12359 GND.n5053 GND.n1167 19.3944
R12360 GND.n5059 GND.n1167 19.3944
R12361 GND.n5059 GND.n1165 19.3944
R12362 GND.n5063 GND.n1165 19.3944
R12363 GND.n5063 GND.n1161 19.3944
R12364 GND.n5069 GND.n1161 19.3944
R12365 GND.n5069 GND.n1159 19.3944
R12366 GND.n5073 GND.n1159 19.3944
R12367 GND.n5073 GND.n1155 19.3944
R12368 GND.n5079 GND.n1155 19.3944
R12369 GND.n5079 GND.n1153 19.3944
R12370 GND.n5083 GND.n1153 19.3944
R12371 GND.n5083 GND.n1149 19.3944
R12372 GND.n5089 GND.n1149 19.3944
R12373 GND.n5089 GND.n1147 19.3944
R12374 GND.n5093 GND.n1147 19.3944
R12375 GND.n5093 GND.n1143 19.3944
R12376 GND.n5099 GND.n1143 19.3944
R12377 GND.n5099 GND.n1141 19.3944
R12378 GND.n5103 GND.n1141 19.3944
R12379 GND.n5103 GND.n1137 19.3944
R12380 GND.n5109 GND.n1137 19.3944
R12381 GND.n5109 GND.n1135 19.3944
R12382 GND.n5113 GND.n1135 19.3944
R12383 GND.n5113 GND.n1131 19.3944
R12384 GND.n5119 GND.n1131 19.3944
R12385 GND.n5119 GND.n1129 19.3944
R12386 GND.n5123 GND.n1129 19.3944
R12387 GND.n5123 GND.n1125 19.3944
R12388 GND.n5129 GND.n1125 19.3944
R12389 GND.n5129 GND.n1123 19.3944
R12390 GND.n5133 GND.n1123 19.3944
R12391 GND.n5133 GND.n1119 19.3944
R12392 GND.n5139 GND.n1119 19.3944
R12393 GND.n5139 GND.n1117 19.3944
R12394 GND.n5143 GND.n1117 19.3944
R12395 GND.n5143 GND.n1113 19.3944
R12396 GND.n5149 GND.n1113 19.3944
R12397 GND.n5149 GND.n1111 19.3944
R12398 GND.n5153 GND.n1111 19.3944
R12399 GND.n5153 GND.n1107 19.3944
R12400 GND.n5159 GND.n1107 19.3944
R12401 GND.n5159 GND.n1105 19.3944
R12402 GND.n5163 GND.n1105 19.3944
R12403 GND.n5163 GND.n1101 19.3944
R12404 GND.n5169 GND.n1101 19.3944
R12405 GND.n5169 GND.n1099 19.3944
R12406 GND.n5173 GND.n1099 19.3944
R12407 GND.n5173 GND.n1095 19.3944
R12408 GND.n5179 GND.n1095 19.3944
R12409 GND.n5179 GND.n1093 19.3944
R12410 GND.n5183 GND.n1093 19.3944
R12411 GND.n5183 GND.n1089 19.3944
R12412 GND.n5189 GND.n1089 19.3944
R12413 GND.n5189 GND.n1087 19.3944
R12414 GND.n5193 GND.n1087 19.3944
R12415 GND.n5193 GND.n1083 19.3944
R12416 GND.n5199 GND.n1083 19.3944
R12417 GND.n5199 GND.n1081 19.3944
R12418 GND.n5203 GND.n1081 19.3944
R12419 GND.n5203 GND.n1077 19.3944
R12420 GND.n5209 GND.n1077 19.3944
R12421 GND.n5209 GND.n1075 19.3944
R12422 GND.n5213 GND.n1075 19.3944
R12423 GND.n5213 GND.n1071 19.3944
R12424 GND.n5219 GND.n1071 19.3944
R12425 GND.n5219 GND.n1069 19.3944
R12426 GND.n5223 GND.n1069 19.3944
R12427 GND.n5223 GND.n1065 19.3944
R12428 GND.n5229 GND.n1065 19.3944
R12429 GND.n5229 GND.n1063 19.3944
R12430 GND.n5233 GND.n1063 19.3944
R12431 GND.n5233 GND.n1059 19.3944
R12432 GND.n5239 GND.n1059 19.3944
R12433 GND.n5239 GND.n1057 19.3944
R12434 GND.n5243 GND.n1057 19.3944
R12435 GND.n5243 GND.n1053 19.3944
R12436 GND.n5249 GND.n1053 19.3944
R12437 GND.n5249 GND.n1051 19.3944
R12438 GND.n5253 GND.n1051 19.3944
R12439 GND.n5253 GND.n1047 19.3944
R12440 GND.n5259 GND.n1047 19.3944
R12441 GND.n5259 GND.n1045 19.3944
R12442 GND.n5263 GND.n1045 19.3944
R12443 GND.n5263 GND.n1041 19.3944
R12444 GND.n5269 GND.n1041 19.3944
R12445 GND.n5269 GND.n1039 19.3944
R12446 GND.n5273 GND.n1039 19.3944
R12447 GND.n5273 GND.n1035 19.3944
R12448 GND.n5279 GND.n1035 19.3944
R12449 GND.n5279 GND.n1033 19.3944
R12450 GND.n5283 GND.n1033 19.3944
R12451 GND.n5283 GND.n1029 19.3944
R12452 GND.n5289 GND.n1029 19.3944
R12453 GND.n5289 GND.n1027 19.3944
R12454 GND.n5293 GND.n1027 19.3944
R12455 GND.n5293 GND.n1023 19.3944
R12456 GND.n5299 GND.n1023 19.3944
R12457 GND.n5299 GND.n1021 19.3944
R12458 GND.n5303 GND.n1021 19.3944
R12459 GND.n5303 GND.n1017 19.3944
R12460 GND.n5309 GND.n1017 19.3944
R12461 GND.n5309 GND.n1015 19.3944
R12462 GND.n5313 GND.n1015 19.3944
R12463 GND.n5313 GND.n1011 19.3944
R12464 GND.n5319 GND.n1011 19.3944
R12465 GND.n5319 GND.n1009 19.3944
R12466 GND.n5323 GND.n1009 19.3944
R12467 GND.n5323 GND.n1005 19.3944
R12468 GND.n5329 GND.n1005 19.3944
R12469 GND.n5329 GND.n1003 19.3944
R12470 GND.n5333 GND.n1003 19.3944
R12471 GND.n5333 GND.n999 19.3944
R12472 GND.n5339 GND.n999 19.3944
R12473 GND.n5339 GND.n997 19.3944
R12474 GND.n5343 GND.n997 19.3944
R12475 GND.n5343 GND.n993 19.3944
R12476 GND.n5349 GND.n993 19.3944
R12477 GND.n5349 GND.n991 19.3944
R12478 GND.n5354 GND.n991 19.3944
R12479 GND.n5354 GND.n987 19.3944
R12480 GND.n5360 GND.n987 19.3944
R12481 GND.n5361 GND.n5360 19.3944
R12482 GND.n2410 GND.n2409 19.3944
R12483 GND.n2409 GND.n2406 19.3944
R12484 GND.n2406 GND.n2405 19.3944
R12485 GND.n2405 GND.n2402 19.3944
R12486 GND.n2402 GND.n2401 19.3944
R12487 GND.n2401 GND.n2398 19.3944
R12488 GND.n2398 GND.n2397 19.3944
R12489 GND.n2397 GND.n2394 19.3944
R12490 GND.n2394 GND.n2393 19.3944
R12491 GND.n2393 GND.n2390 19.3944
R12492 GND.n2390 GND.n2389 19.3944
R12493 GND.n2389 GND.n2386 19.3944
R12494 GND.n2386 GND.n2003 19.3944
R12495 GND.n4311 GND.n2009 19.3944
R12496 GND.n2131 GND.n2009 19.3944
R12497 GND.n2131 GND.n2127 19.3944
R12498 GND.n2135 GND.n2127 19.3944
R12499 GND.n2138 GND.n2135 19.3944
R12500 GND.n2141 GND.n2138 19.3944
R12501 GND.n2141 GND.n2125 19.3944
R12502 GND.n2145 GND.n2125 19.3944
R12503 GND.n2148 GND.n2145 19.3944
R12504 GND.n2151 GND.n2148 19.3944
R12505 GND.n2151 GND.n2123 19.3944
R12506 GND.n2155 GND.n2123 19.3944
R12507 GND.n2158 GND.n2155 19.3944
R12508 GND.n2161 GND.n2158 19.3944
R12509 GND.n2161 GND.n2120 19.3944
R12510 GND.n2165 GND.n2120 19.3944
R12511 GND.n3984 GND.n2371 19.3944
R12512 GND.n3984 GND.n2369 19.3944
R12513 GND.n3990 GND.n2369 19.3944
R12514 GND.n3990 GND.n3989 19.3944
R12515 GND.n3989 GND.n2348 19.3944
R12516 GND.n4009 GND.n2348 19.3944
R12517 GND.n4009 GND.n2346 19.3944
R12518 GND.n4015 GND.n2346 19.3944
R12519 GND.n4015 GND.n4014 19.3944
R12520 GND.n4014 GND.n2325 19.3944
R12521 GND.n4033 GND.n2325 19.3944
R12522 GND.n4033 GND.n2323 19.3944
R12523 GND.n4039 GND.n2323 19.3944
R12524 GND.n4039 GND.n4038 19.3944
R12525 GND.n4038 GND.n2302 19.3944
R12526 GND.n4058 GND.n2302 19.3944
R12527 GND.n4058 GND.n2300 19.3944
R12528 GND.n4065 GND.n2300 19.3944
R12529 GND.n4065 GND.n4064 19.3944
R12530 GND.n4064 GND.n2272 19.3944
R12531 GND.n4141 GND.n2272 19.3944
R12532 GND.n4139 GND.n4138 19.3944
R12533 GND.n4095 GND.n4094 19.3944
R12534 GND.n4124 GND.n4123 19.3944
R12535 GND.n4121 GND.n4097 19.3944
R12536 GND.n4099 GND.n2245 19.3944
R12537 GND.n4167 GND.n2245 19.3944
R12538 GND.n4167 GND.n2243 19.3944
R12539 GND.n4173 GND.n2243 19.3944
R12540 GND.n4173 GND.n4172 19.3944
R12541 GND.n4172 GND.n866 19.3944
R12542 GND.n5546 GND.n866 19.3944
R12543 GND.n5546 GND.n864 19.3944
R12544 GND.n5550 GND.n864 19.3944
R12545 GND.n5550 GND.n844 19.3944
R12546 GND.n5563 GND.n844 19.3944
R12547 GND.n5563 GND.n842 19.3944
R12548 GND.n5567 GND.n842 19.3944
R12549 GND.n5567 GND.n825 19.3944
R12550 GND.n5580 GND.n825 19.3944
R12551 GND.n5580 GND.n823 19.3944
R12552 GND.n5584 GND.n823 19.3944
R12553 GND.n5584 GND.n808 19.3944
R12554 GND.n5598 GND.n808 19.3944
R12555 GND.n5598 GND.n806 19.3944
R12556 GND.n5603 GND.n806 19.3944
R12557 GND.n5603 GND.n5602 19.3944
R12558 GND.n2788 GND.n2787 19.3944
R12559 GND.n2787 GND.n2786 19.3944
R12560 GND.n2786 GND.n2779 19.3944
R12561 GND.n2782 GND.n2779 19.3944
R12562 GND.n2782 GND.n2735 19.3944
R12563 GND.n2993 GND.n2735 19.3944
R12564 GND.n2993 GND.n2733 19.3944
R12565 GND.n2997 GND.n2733 19.3944
R12566 GND.n3001 GND.n2997 19.3944
R12567 GND.n2999 GND.n2998 19.3944
R12568 GND.n3094 GND.n3093 19.3944
R12569 GND.n3091 GND.n2703 19.3944
R12570 GND.n3077 GND.n3025 19.3944
R12571 GND.n3075 GND.n3074 19.3944
R12572 GND.n3074 GND.n3027 19.3944
R12573 GND.n3068 GND.n3027 19.3944
R12574 GND.n3068 GND.n3067 19.3944
R12575 GND.n3067 GND.n3066 19.3944
R12576 GND.n3066 GND.n3033 19.3944
R12577 GND.n3059 GND.n3033 19.3944
R12578 GND.n3059 GND.n3058 19.3944
R12579 GND.n3058 GND.n3057 19.3944
R12580 GND.n3057 GND.n3039 19.3944
R12581 GND.n3053 GND.n3039 19.3944
R12582 GND.n3053 GND.n3052 19.3944
R12583 GND.n3052 GND.n3051 19.3944
R12584 GND.n3051 GND.n3049 19.3944
R12585 GND.n3049 GND.n2617 19.3944
R12586 GND.n2617 GND.n2615 19.3944
R12587 GND.n3190 GND.n2615 19.3944
R12588 GND.n3190 GND.n2613 19.3944
R12589 GND.n3203 GND.n2613 19.3944
R12590 GND.n3203 GND.n3202 19.3944
R12591 GND.n3202 GND.n3201 19.3944
R12592 GND.n3201 GND.n3198 19.3944
R12593 GND.n3198 GND.n1642 19.3944
R12594 GND.n4555 GND.n1642 19.3944
R12595 GND.n4555 GND.n4554 19.3944
R12596 GND.n4554 GND.n4553 19.3944
R12597 GND.n4553 GND.n1646 19.3944
R12598 GND.n1673 GND.n1646 19.3944
R12599 GND.n4543 GND.n1673 19.3944
R12600 GND.n4543 GND.n4542 19.3944
R12601 GND.n4542 GND.n4541 19.3944
R12602 GND.n4541 GND.n1679 19.3944
R12603 GND.n1699 GND.n1679 19.3944
R12604 GND.n4529 GND.n1699 19.3944
R12605 GND.n4529 GND.n4528 19.3944
R12606 GND.n4528 GND.n4527 19.3944
R12607 GND.n4527 GND.n1705 19.3944
R12608 GND.n1726 GND.n1705 19.3944
R12609 GND.n4515 GND.n1726 19.3944
R12610 GND.n4515 GND.n4514 19.3944
R12611 GND.n4514 GND.n4513 19.3944
R12612 GND.n4513 GND.n1732 19.3944
R12613 GND.n2551 GND.n1732 19.3944
R12614 GND.n2551 GND.n2548 19.3944
R12615 GND.n2555 GND.n2548 19.3944
R12616 GND.n2555 GND.n2546 19.3944
R12617 GND.n2559 GND.n2546 19.3944
R12618 GND.n2559 GND.n2544 19.3944
R12619 GND.n3520 GND.n2544 19.3944
R12620 GND.n3520 GND.n2542 19.3944
R12621 GND.n3534 GND.n2542 19.3944
R12622 GND.n3534 GND.n3533 19.3944
R12623 GND.n3533 GND.n3532 19.3944
R12624 GND.n3532 GND.n3529 19.3944
R12625 GND.n3529 GND.n3528 19.3944
R12626 GND.n3528 GND.n2526 19.3944
R12627 GND.n3586 GND.n2526 19.3944
R12628 GND.n3586 GND.n2524 19.3944
R12629 GND.n3599 GND.n2524 19.3944
R12630 GND.n3599 GND.n3598 19.3944
R12631 GND.n3598 GND.n3597 19.3944
R12632 GND.n3597 GND.n3594 19.3944
R12633 GND.n3594 GND.n1848 19.3944
R12634 GND.n4431 GND.n1848 19.3944
R12635 GND.n4431 GND.n4430 19.3944
R12636 GND.n4430 GND.n4429 19.3944
R12637 GND.n4429 GND.n1852 19.3944
R12638 GND.n1895 GND.n1852 19.3944
R12639 GND.n1898 GND.n1895 19.3944
R12640 GND.n1898 GND.n1892 19.3944
R12641 GND.n4404 GND.n1892 19.3944
R12642 GND.n4404 GND.n4403 19.3944
R12643 GND.n4403 GND.n4402 19.3944
R12644 GND.n4402 GND.n1904 19.3944
R12645 GND.n1934 GND.n1904 19.3944
R12646 GND.n1934 GND.n1931 19.3944
R12647 GND.n4383 GND.n1931 19.3944
R12648 GND.n4383 GND.n4382 19.3944
R12649 GND.n4382 GND.n4381 19.3944
R12650 GND.n4381 GND.n1940 19.3944
R12651 GND.n2468 GND.n1940 19.3944
R12652 GND.n2468 GND.n2465 19.3944
R12653 GND.n3819 GND.n2465 19.3944
R12654 GND.n3819 GND.n2463 19.3944
R12655 GND.n3825 GND.n2463 19.3944
R12656 GND.n3825 GND.n3824 19.3944
R12657 GND.n3824 GND.n2442 19.3944
R12658 GND.n3855 GND.n2442 19.3944
R12659 GND.n3855 GND.n2440 19.3944
R12660 GND.n3859 GND.n2440 19.3944
R12661 GND.n3859 GND.n2427 19.3944
R12662 GND.n3874 GND.n2427 19.3944
R12663 GND.n3874 GND.n2425 19.3944
R12664 GND.n3878 GND.n2425 19.3944
R12665 GND.n3878 GND.n2423 19.3944
R12666 GND.n3906 GND.n2423 19.3944
R12667 GND.n3906 GND.n2421 19.3944
R12668 GND.n3910 GND.n2421 19.3944
R12669 GND.n3910 GND.n2419 19.3944
R12670 GND.n3921 GND.n2419 19.3944
R12671 GND.n3921 GND.n2417 19.3944
R12672 GND.n3975 GND.n2417 19.3944
R12673 GND.n3975 GND.n3974 19.3944
R12674 GND.n3974 GND.n3973 19.3944
R12675 GND.n3973 GND.n3927 19.3944
R12676 GND.n3969 GND.n3927 19.3944
R12677 GND.n3969 GND.n3968 19.3944
R12678 GND.n3968 GND.n3967 19.3944
R12679 GND.n3967 GND.n3933 19.3944
R12680 GND.n3963 GND.n3933 19.3944
R12681 GND.n3963 GND.n3962 19.3944
R12682 GND.n3962 GND.n3961 19.3944
R12683 GND.n3961 GND.n3939 19.3944
R12684 GND.n3957 GND.n3939 19.3944
R12685 GND.n3957 GND.n3956 19.3944
R12686 GND.n3956 GND.n3955 19.3944
R12687 GND.n3955 GND.n3945 19.3944
R12688 GND.n3951 GND.n3945 19.3944
R12689 GND.n3951 GND.n3950 19.3944
R12690 GND.n3950 GND.n2261 19.3944
R12691 GND.n4146 GND.n2261 19.3944
R12692 GND.n4146 GND.n2262 19.3944
R12693 GND.n4087 GND.n4086 19.3944
R12694 GND.n4130 GND.n4129 19.3944
R12695 GND.n4108 GND.n4107 19.3944
R12696 GND.n4111 GND.n4110 19.3944
R12697 GND.n4158 GND.n4157 19.3944
R12698 GND.n4157 GND.n4156 19.3944
R12699 GND.n4156 GND.n4153 19.3944
R12700 GND.n4153 GND.n884 19.3944
R12701 GND.n5533 GND.n884 19.3944
R12702 GND.n5533 GND.n5532 19.3944
R12703 GND.n5532 GND.n5531 19.3944
R12704 GND.n5531 GND.n888 19.3944
R12705 GND.n5525 GND.n888 19.3944
R12706 GND.n4834 GND.n4833 19.3944
R12707 GND.n4833 GND.n4832 19.3944
R12708 GND.n4832 GND.n4831 19.3944
R12709 GND.n4831 GND.n4829 19.3944
R12710 GND.n4829 GND.n4826 19.3944
R12711 GND.n4826 GND.n4825 19.3944
R12712 GND.n4825 GND.n4822 19.3944
R12713 GND.n4822 GND.n4821 19.3944
R12714 GND.n4821 GND.n4818 19.3944
R12715 GND.n4818 GND.n4817 19.3944
R12716 GND.n4817 GND.n4814 19.3944
R12717 GND.n4814 GND.n4813 19.3944
R12718 GND.n4813 GND.n4810 19.3944
R12719 GND.n4810 GND.n4809 19.3944
R12720 GND.n4809 GND.n4806 19.3944
R12721 GND.n4804 GND.n4801 19.3944
R12722 GND.n4801 GND.n4800 19.3944
R12723 GND.n4800 GND.n4797 19.3944
R12724 GND.n4797 GND.n4796 19.3944
R12725 GND.n4796 GND.n4793 19.3944
R12726 GND.n4793 GND.n4792 19.3944
R12727 GND.n4792 GND.n4789 19.3944
R12728 GND.n4789 GND.n4788 19.3944
R12729 GND.n4788 GND.n4785 19.3944
R12730 GND.n4785 GND.n4784 19.3944
R12731 GND.n4784 GND.n4781 19.3944
R12732 GND.n4781 GND.n4780 19.3944
R12733 GND.n4780 GND.n4777 19.3944
R12734 GND.n4777 GND.n4776 19.3944
R12735 GND.n4776 GND.n4773 19.3944
R12736 GND.n4773 GND.n4772 19.3944
R12737 GND.n2904 GND.n2903 19.3944
R12738 GND.n2908 GND.n2903 19.3944
R12739 GND.n2908 GND.n2809 19.3944
R12740 GND.n2917 GND.n2809 19.3944
R12741 GND.n2917 GND.n2807 19.3944
R12742 GND.n2921 GND.n2807 19.3944
R12743 GND.n2921 GND.n2796 19.3944
R12744 GND.n2930 GND.n2796 19.3944
R12745 GND.n2930 GND.n2794 19.3944
R12746 GND.n2934 GND.n2794 19.3944
R12747 GND.n2934 GND.n2770 19.3944
R12748 GND.n2946 GND.n2770 19.3944
R12749 GND.n2946 GND.n2768 19.3944
R12750 GND.n2952 GND.n2768 19.3944
R12751 GND.n2952 GND.n2951 19.3944
R12752 GND.n2951 GND.n2747 19.3944
R12753 GND.n2983 GND.n2747 19.3944
R12754 GND.n2983 GND.n2745 19.3944
R12755 GND.n2988 GND.n2745 19.3944
R12756 GND.n2988 GND.n2987 19.3944
R12757 GND.n2987 GND.n2689 19.3944
R12758 GND.n3104 GND.n3103 19.3944
R12759 GND.n2713 GND.n2712 19.3944
R12760 GND.n3086 GND.n3085 19.3944
R12761 GND.n2718 GND.n2717 19.3944
R12762 GND.n3109 GND.n2682 19.3944
R12763 GND.n3109 GND.n3108 19.3944
R12764 GND.n3108 GND.n2663 19.3944
R12765 GND.n3128 GND.n2663 19.3944
R12766 GND.n3128 GND.n2661 19.3944
R12767 GND.n3134 GND.n2661 19.3944
R12768 GND.n3134 GND.n3133 19.3944
R12769 GND.n3133 GND.n2644 19.3944
R12770 GND.n3153 GND.n2644 19.3944
R12771 GND.n3153 GND.n2642 19.3944
R12772 GND.n3159 GND.n2642 19.3944
R12773 GND.n3159 GND.n3158 19.3944
R12774 GND.n3158 GND.n2623 19.3944
R12775 GND.n3179 GND.n2623 19.3944
R12776 GND.n3179 GND.n2621 19.3944
R12777 GND.n3183 GND.n2621 19.3944
R12778 GND.n3183 GND.n2597 19.3944
R12779 GND.n3219 GND.n2597 19.3944
R12780 GND.n3219 GND.n2595 19.3944
R12781 GND.n3223 GND.n2595 19.3944
R12782 GND.n3223 GND.n1531 19.3944
R12783 GND.n4683 GND.n1531 19.3944
R12784 GND.n4963 GND.n4962 19.3944
R12785 GND.n4962 GND.n4961 19.3944
R12786 GND.n4961 GND.n1228 19.3944
R12787 GND.n4955 GND.n1228 19.3944
R12788 GND.n4955 GND.n4954 19.3944
R12789 GND.n4954 GND.n4953 19.3944
R12790 GND.n4953 GND.n1236 19.3944
R12791 GND.n4947 GND.n1236 19.3944
R12792 GND.n4947 GND.n4946 19.3944
R12793 GND.n4946 GND.n4945 19.3944
R12794 GND.n4945 GND.n1244 19.3944
R12795 GND.n4939 GND.n1244 19.3944
R12796 GND.n4939 GND.n4938 19.3944
R12797 GND.n4938 GND.n4937 19.3944
R12798 GND.n4937 GND.n1252 19.3944
R12799 GND.n4931 GND.n1252 19.3944
R12800 GND.n4931 GND.n4930 19.3944
R12801 GND.n4930 GND.n4929 19.3944
R12802 GND.n4929 GND.n1260 19.3944
R12803 GND.n4923 GND.n1260 19.3944
R12804 GND.n4923 GND.n4922 19.3944
R12805 GND.n4922 GND.n4921 19.3944
R12806 GND.n4921 GND.n1268 19.3944
R12807 GND.n4915 GND.n1268 19.3944
R12808 GND.n4915 GND.n4914 19.3944
R12809 GND.n4914 GND.n4913 19.3944
R12810 GND.n4913 GND.n1276 19.3944
R12811 GND.n4907 GND.n1276 19.3944
R12812 GND.n4907 GND.n4906 19.3944
R12813 GND.n4906 GND.n4905 19.3944
R12814 GND.n4905 GND.n1284 19.3944
R12815 GND.n4899 GND.n1284 19.3944
R12816 GND.n4899 GND.n4898 19.3944
R12817 GND.n4898 GND.n4897 19.3944
R12818 GND.n4897 GND.n1292 19.3944
R12819 GND.n4891 GND.n1292 19.3944
R12820 GND.n4891 GND.n4890 19.3944
R12821 GND.n4890 GND.n4889 19.3944
R12822 GND.n4889 GND.n1300 19.3944
R12823 GND.n4883 GND.n1300 19.3944
R12824 GND.n4883 GND.n4882 19.3944
R12825 GND.n4882 GND.n4881 19.3944
R12826 GND.n4881 GND.n1308 19.3944
R12827 GND.n4875 GND.n1308 19.3944
R12828 GND.n4875 GND.n4874 19.3944
R12829 GND.n4874 GND.n4873 19.3944
R12830 GND.n4873 GND.n1316 19.3944
R12831 GND.n4867 GND.n1316 19.3944
R12832 GND.n4867 GND.n4866 19.3944
R12833 GND.n4866 GND.n4865 19.3944
R12834 GND.n4865 GND.n1324 19.3944
R12835 GND.n4859 GND.n1324 19.3944
R12836 GND.n4859 GND.n4858 19.3944
R12837 GND.n4858 GND.n4857 19.3944
R12838 GND.n4857 GND.n1332 19.3944
R12839 GND.n4851 GND.n1332 19.3944
R12840 GND.n4851 GND.n4850 19.3944
R12841 GND.n4850 GND.n4849 19.3944
R12842 GND.n4849 GND.n1340 19.3944
R12843 GND.n4843 GND.n1340 19.3944
R12844 GND.n4843 GND.n4842 19.3944
R12845 GND.n4842 GND.n4841 19.3944
R12846 GND.n4841 GND.n1348 19.3944
R12847 GND.n4306 GND.n4305 19.3944
R12848 GND.n4305 GND.n2042 19.3944
R12849 GND.n4298 GND.n2042 19.3944
R12850 GND.n4298 GND.n4297 19.3944
R12851 GND.n4297 GND.n2052 19.3944
R12852 GND.n4290 GND.n2052 19.3944
R12853 GND.n4290 GND.n4289 19.3944
R12854 GND.n4289 GND.n2060 19.3944
R12855 GND.n4282 GND.n2060 19.3944
R12856 GND.n4282 GND.n4281 19.3944
R12857 GND.n4281 GND.n2070 19.3944
R12858 GND.n4274 GND.n2070 19.3944
R12859 GND.n4274 GND.n4273 19.3944
R12860 GND.n4273 GND.n2078 19.3944
R12861 GND.n3916 GND.n3913 19.3944
R12862 GND.n3913 GND.n2360 19.3944
R12863 GND.n3994 GND.n2360 19.3944
R12864 GND.n3994 GND.n2357 19.3944
R12865 GND.n3999 GND.n2357 19.3944
R12866 GND.n3999 GND.n2358 19.3944
R12867 GND.n2358 GND.n2338 19.3944
R12868 GND.n4019 GND.n2338 19.3944
R12869 GND.n4019 GND.n2335 19.3944
R12870 GND.n4024 GND.n2335 19.3944
R12871 GND.n4024 GND.n2336 19.3944
R12872 GND.n2336 GND.n2314 19.3944
R12873 GND.n4043 GND.n2314 19.3944
R12874 GND.n4043 GND.n2311 19.3944
R12875 GND.n4048 GND.n2311 19.3944
R12876 GND.n4048 GND.n2312 19.3944
R12877 GND.n2312 GND.n2287 19.3944
R12878 GND.n4069 GND.n2287 19.3944
R12879 GND.n4069 GND.n2284 19.3944
R12880 GND.n4073 GND.n2284 19.3944
R12881 GND.n4074 GND.n4073 19.3944
R12882 GND.n4077 GND.n4074 19.3944
R12883 GND.n4077 GND.n2282 19.3944
R12884 GND.n4081 GND.n2282 19.3944
R12885 GND.n4081 GND.n676 19.3944
R12886 GND.n5756 GND.n676 19.3944
R12887 GND.n5756 GND.n5755 19.3944
R12888 GND.n5755 GND.n5754 19.3944
R12889 GND.n5754 GND.n680 19.3944
R12890 GND.n5750 GND.n680 19.3944
R12891 GND.n5750 GND.n5749 19.3944
R12892 GND.n5749 GND.n5748 19.3944
R12893 GND.n5748 GND.n685 19.3944
R12894 GND.n5744 GND.n685 19.3944
R12895 GND.n5744 GND.n5743 19.3944
R12896 GND.n5743 GND.n5742 19.3944
R12897 GND.n5742 GND.n690 19.3944
R12898 GND.n5738 GND.n690 19.3944
R12899 GND.n5738 GND.n5737 19.3944
R12900 GND.n5737 GND.n5736 19.3944
R12901 GND.n5736 GND.n695 19.3944
R12902 GND.n5732 GND.n695 19.3944
R12903 GND.n5732 GND.n5731 19.3944
R12904 GND.n5731 GND.n5730 19.3944
R12905 GND.n5730 GND.n700 19.3944
R12906 GND.n5726 GND.n700 19.3944
R12907 GND.n5726 GND.n5725 19.3944
R12908 GND.n5725 GND.n5724 19.3944
R12909 GND.n5724 GND.n705 19.3944
R12910 GND.n5720 GND.n705 19.3944
R12911 GND.n5720 GND.n5719 19.3944
R12912 GND.n5719 GND.n5718 19.3944
R12913 GND.n4661 GND.n4660 18.4247
R12914 GND.n4312 GND.n2003 18.4247
R12915 GND.n5628 GND.n713 18.2308
R12916 GND.n4593 GND.n1620 18.2308
R12917 GND.n2869 GND.n2868 18.2308
R12918 GND.n4266 GND.n2078 18.2308
R12919 GND.n4550 GND.n1665 17.188
R12920 GND.n3902 GND.n3881 17.188
R12921 GND.n4546 GND.n1668 16.5269
R12922 GND.n4546 GND.n4545 16.5269
R12923 GND.n4545 GND.n1670 16.5269
R12924 GND.n3271 GND.n1670 16.5269
R12925 GND.n3272 GND.n3271 16.5269
R12926 GND.n4539 GND.n4538 16.5269
R12927 GND.n4538 GND.n1682 16.5269
R12928 GND.n2581 GND.n1682 16.5269
R12929 GND.n2581 GND.n1694 16.5269
R12930 GND.n4532 GND.n1694 16.5269
R12931 GND.n4532 GND.n4531 16.5269
R12932 GND.n4531 GND.n1696 16.5269
R12933 GND.n1707 GND.n1696 16.5269
R12934 GND.n1708 GND.n1707 16.5269
R12935 GND.n4525 GND.n1708 16.5269
R12936 GND.n4525 GND.n4524 16.5269
R12937 GND.n4524 GND.n1710 16.5269
R12938 GND.n3287 GND.n1710 16.5269
R12939 GND.n4518 GND.n1721 16.5269
R12940 GND.n4518 GND.n4517 16.5269
R12941 GND.n4517 GND.n1723 16.5269
R12942 GND.n2574 GND.n1723 16.5269
R12943 GND.n2575 GND.n2574 16.5269
R12944 GND.n4511 GND.n4510 16.5269
R12945 GND.n4504 GND.n1746 16.5269
R12946 GND.n3488 GND.n1755 16.5269
R12947 GND.n3549 GND.n1789 16.5269
R12948 GND.n3549 GND.n1795 16.5269
R12949 GND.n3568 GND.n2531 16.5269
R12950 GND.n3583 GND.n3582 16.5269
R12951 GND.n3557 GND.n3556 16.5269
R12952 GND.n3612 GND.n1827 16.5269
R12953 GND.n4440 GND.n1836 16.5269
R12954 GND.n4434 GND.n4433 16.5269
R12955 GND.n4427 GND.n1854 16.5269
R12956 GND.n4419 GND.n1865 16.5269
R12957 GND.n4413 GND.n1879 16.5269
R12958 GND.n4413 GND.n1882 16.5269
R12959 GND.n4400 GND.n4399 16.5269
R12960 GND.n4393 GND.n1917 16.5269
R12961 GND.n4385 GND.n1928 16.5269
R12962 GND.n4379 GND.n1942 16.5269
R12963 GND.n3786 GND.n3785 16.5269
R12964 GND.n3786 GND.n1969 16.5269
R12965 GND.n3806 GND.n2478 16.5269
R12966 GND.n2478 GND.n2471 16.5269
R12967 GND.n3817 GND.n2471 16.5269
R12968 GND.n3817 GND.n3816 16.5269
R12969 GND.n3816 GND.n3815 16.5269
R12970 GND.n3828 GND.n3827 16.5269
R12971 GND.n3827 GND.n2460 16.5269
R12972 GND.n2460 GND.n2451 16.5269
R12973 GND.n3838 GND.n2451 16.5269
R12974 GND.n3838 GND.n2452 16.5269
R12975 GND.n2452 GND.n2444 16.5269
R12976 GND.n3853 GND.n2444 16.5269
R12977 GND.n3853 GND.n3852 16.5269
R12978 GND.n3852 GND.n2435 16.5269
R12979 GND.n3862 GND.n2435 16.5269
R12980 GND.n3862 GND.n3861 16.5269
R12981 GND.n3861 GND.n2438 16.5269
R12982 GND.n2438 GND.n2437 16.5269
R12983 GND.n3872 GND.n3870 16.5269
R12984 GND.n3872 GND.n3871 16.5269
R12985 GND.n3871 GND.n2108 16.5269
R12986 GND.n4238 GND.n2108 16.5269
R12987 GND.n4238 GND.n2109 16.5269
R12988 GND.n3272 GND.t103 16.1964
R12989 GND.n3870 GND.t110 16.1964
R12990 GND.n4551 GND.n4550 15.8659
R12991 GND.n3480 GND.n3479 15.8659
R12992 GND.n4448 GND.n4447 15.8659
R12993 GND.n3624 GND.n3623 15.8659
R12994 GND.n4386 GND.n1926 15.8659
R12995 GND.n4378 GND.n1944 15.8659
R12996 GND.n3904 GND.n3902 15.8659
R12997 GND.n80 GND.n78 15.6674
R12998 GND.n117 GND.n115 15.6674
R12999 GND.n149 GND.n147 15.6674
R13000 GND.n186 GND.n184 15.6674
R13001 GND.n11 GND.n9 15.6674
R13002 GND.n48 GND.n46 15.6674
R13003 GND.n513 GND.n511 15.6674
R13004 GND.n476 GND.n474 15.6674
R13005 GND.n582 GND.n580 15.6674
R13006 GND.n545 GND.n543 15.6674
R13007 GND.n652 GND.n650 15.6674
R13008 GND.n615 GND.n613 15.6674
R13009 GND.n316 GND.n314 15.6674
R13010 GND.n284 GND.n282 15.6674
R13011 GND.n252 GND.n250 15.6674
R13012 GND.n221 GND.n219 15.6674
R13013 GND.n443 GND.n441 15.6674
R13014 GND.n411 GND.n409 15.6674
R13015 GND.n379 GND.n377 15.6674
R13016 GND.n348 GND.n346 15.6674
R13017 GND.n3540 GND.n2538 15.2048
R13018 GND.n3572 GND.n3569 15.2048
R13019 GND.n4420 GND.n1862 15.2048
R13020 GND.n2496 GND.n2489 15.2048
R13021 GND.n1952 GND.n1951 15.0827
R13022 GND.n3341 GND.n3336 15.0481
R13023 GND.n1962 GND.n1961 15.0481
R13024 GND.n2575 GND.n1734 14.8743
R13025 GND.n4510 GND.t82 14.5438
R13026 GND.n4490 GND.n1766 14.5438
R13027 GND.t114 GND.n3515 13.8827
R13028 GND.n3503 GND.n1769 13.8827
R13029 GND.t29 GND.n1775 13.8827
R13030 GND.n3581 GND.n1814 13.8827
R13031 GND.n3633 GND.n2508 13.8827
R13032 GND.n2482 GND.n1908 13.8827
R13033 GND.n5662 GND.n797 13.5763
R13034 GND.n4635 GND.n1578 13.5763
R13035 GND.n2166 GND.n2165 13.5763
R13036 GND.n4772 GND.n1417 13.5763
R13037 GND.n4483 GND.n4482 13.2217
R13038 GND.t19 GND.n3536 13.2217
R13039 GND.n4462 GND.n4461 13.2217
R13040 GND.n4426 GND.n1856 13.2217
R13041 GND.n4406 GND.t7 13.2217
R13042 GND.n3685 GND.n1906 13.2217
R13043 GND.n3352 GND.n3333 13.1884
R13044 GND.n3347 GND.n3346 13.1884
R13045 GND.n3346 GND.n3345 13.1884
R13046 GND.n1955 GND.n1950 13.1884
R13047 GND.n1956 GND.n1955 13.1884
R13048 GND.n3348 GND.n3335 13.146
R13049 GND.n3344 GND.n3335 13.146
R13050 GND.n1954 GND.n1953 13.146
R13051 GND.n1954 GND.n1949 13.146
R13052 GND.n81 GND.n77 12.8005
R13053 GND.n118 GND.n114 12.8005
R13054 GND.n150 GND.n146 12.8005
R13055 GND.n187 GND.n183 12.8005
R13056 GND.n12 GND.n8 12.8005
R13057 GND.n49 GND.n45 12.8005
R13058 GND.n514 GND.n510 12.8005
R13059 GND.n477 GND.n473 12.8005
R13060 GND.n583 GND.n579 12.8005
R13061 GND.n546 GND.n542 12.8005
R13062 GND.n653 GND.n649 12.8005
R13063 GND.n616 GND.n612 12.8005
R13064 GND.n3353 GND.n3332 12.8005
R13065 GND.n4374 GND.n4373 12.8005
R13066 GND.n317 GND.n313 12.8005
R13067 GND.n285 GND.n281 12.8005
R13068 GND.n253 GND.n249 12.8005
R13069 GND.n222 GND.n218 12.8005
R13070 GND.n444 GND.n440 12.8005
R13071 GND.n412 GND.n408 12.8005
R13072 GND.n380 GND.n376 12.8005
R13073 GND.n349 GND.n345 12.8005
R13074 GND.n4583 GND.n4557 12.5606
R13075 GND.n2563 GND.n2560 12.5606
R13076 GND.n3604 GND.n3601 12.5606
R13077 GND.n3640 GND.n2512 12.5606
R13078 GND.n3707 GND.t107 12.5606
R13079 GND.n4392 GND.n1920 12.5606
R13080 GND.n4308 GND.n2011 12.5606
R13081 GND.n5658 GND.n797 12.4126
R13082 GND.n4631 GND.n1578 12.4126
R13083 GND.n2167 GND.n2166 12.4126
R13084 GND.n4768 GND.n1417 12.4126
R13085 GND.n85 GND.n84 12.0247
R13086 GND.n122 GND.n121 12.0247
R13087 GND.n154 GND.n153 12.0247
R13088 GND.n191 GND.n190 12.0247
R13089 GND.n16 GND.n15 12.0247
R13090 GND.n53 GND.n52 12.0247
R13091 GND.n518 GND.n517 12.0247
R13092 GND.n481 GND.n480 12.0247
R13093 GND.n587 GND.n586 12.0247
R13094 GND.n550 GND.n549 12.0247
R13095 GND.n657 GND.n656 12.0247
R13096 GND.n620 GND.n619 12.0247
R13097 GND.n321 GND.n320 12.0247
R13098 GND.n289 GND.n288 12.0247
R13099 GND.n257 GND.n256 12.0247
R13100 GND.n226 GND.n225 12.0247
R13101 GND.n448 GND.n447 12.0247
R13102 GND.n416 GND.n415 12.0247
R13103 GND.n384 GND.n383 12.0247
R13104 GND.n353 GND.n352 12.0247
R13105 GND.n4476 GND.n1786 11.8995
R13106 GND.n4468 GND.n1798 11.8995
R13107 GND.n3661 GND.n2501 11.8995
R13108 GND.n4407 GND.n1888 11.8995
R13109 GND.n3145 GND.t129 11.569
R13110 GND.n2321 GND.t122 11.569
R13111 GND.n88 GND.n75 11.249
R13112 GND.n125 GND.n112 11.249
R13113 GND.n157 GND.n144 11.249
R13114 GND.n194 GND.n181 11.249
R13115 GND.n19 GND.n6 11.249
R13116 GND.n56 GND.n43 11.249
R13117 GND.n521 GND.n508 11.249
R13118 GND.n484 GND.n471 11.249
R13119 GND.n590 GND.n577 11.249
R13120 GND.n553 GND.n540 11.249
R13121 GND.n660 GND.n647 11.249
R13122 GND.n623 GND.n610 11.249
R13123 GND.n324 GND.n311 11.249
R13124 GND.n292 GND.n279 11.249
R13125 GND.n260 GND.n247 11.249
R13126 GND.n229 GND.n216 11.249
R13127 GND.n451 GND.n438 11.249
R13128 GND.n419 GND.n406 11.249
R13129 GND.n387 GND.n374 11.249
R13130 GND.n356 GND.n343 11.249
R13131 GND.n4503 GND.n1749 11.2385
R13132 GND.n3489 GND.n1749 11.2385
R13133 GND.n3611 GND.n1833 11.2385
R13134 GND.n4441 GND.n1833 11.2385
R13135 GND.n3719 GND.n3718 11.2385
R13136 GND.n3097 GND.t116 10.908
R13137 GND.n3287 GND.t0 10.908
R13138 GND.n3828 GND.t17 10.908
R13139 GND.n4119 GND.t145 10.908
R13140 GND.n3728 GND.n2002 10.6151
R13141 GND.n3729 GND.n3728 10.6151
R13142 GND.n3733 GND.n3732 10.6151
R13143 GND.n3736 GND.n3733 10.6151
R13144 GND.n3737 GND.n3736 10.6151
R13145 GND.n3740 GND.n3737 10.6151
R13146 GND.n3741 GND.n3740 10.6151
R13147 GND.n3744 GND.n3741 10.6151
R13148 GND.n3745 GND.n3744 10.6151
R13149 GND.n3748 GND.n3745 10.6151
R13150 GND.n3749 GND.n3748 10.6151
R13151 GND.n3752 GND.n3749 10.6151
R13152 GND.n3753 GND.n3752 10.6151
R13153 GND.n3756 GND.n3753 10.6151
R13154 GND.n3757 GND.n3756 10.6151
R13155 GND.n3760 GND.n3757 10.6151
R13156 GND.n3761 GND.n3760 10.6151
R13157 GND.n3764 GND.n3761 10.6151
R13158 GND.n3765 GND.n3764 10.6151
R13159 GND.n3768 GND.n3765 10.6151
R13160 GND.n3769 GND.n3768 10.6151
R13161 GND.n3772 GND.n3769 10.6151
R13162 GND.n3773 GND.n3772 10.6151
R13163 GND.n3776 GND.n3773 10.6151
R13164 GND.n3777 GND.n3776 10.6151
R13165 GND.n3780 GND.n3777 10.6151
R13166 GND.n3781 GND.n3780 10.6151
R13167 GND.n3477 GND.n3476 10.6151
R13168 GND.n3477 GND.n2569 10.6151
R13169 GND.n3491 GND.n2569 10.6151
R13170 GND.n3492 GND.n3491 10.6151
R13171 GND.n3493 GND.n3492 10.6151
R13172 GND.n3493 GND.n2568 10.6151
R13173 GND.n3497 GND.n2568 10.6151
R13174 GND.n3498 GND.n3497 10.6151
R13175 GND.n3501 GND.n3498 10.6151
R13176 GND.n3501 GND.n3500 10.6151
R13177 GND.n3500 GND.n3499 10.6151
R13178 GND.n3499 GND.n2536 10.6151
R13179 GND.n3543 GND.n2536 10.6151
R13180 GND.n3544 GND.n3543 10.6151
R13181 GND.n3547 GND.n3544 10.6151
R13182 GND.n3547 GND.n3546 10.6151
R13183 GND.n3546 GND.n3545 10.6151
R13184 GND.n3545 GND.n2529 10.6151
R13185 GND.n3575 GND.n2529 10.6151
R13186 GND.n3576 GND.n3575 10.6151
R13187 GND.n3579 GND.n3576 10.6151
R13188 GND.n3579 GND.n3578 10.6151
R13189 GND.n3578 GND.n3577 10.6151
R13190 GND.n3577 GND.n2520 10.6151
R13191 GND.n3607 GND.n2520 10.6151
R13192 GND.n3608 GND.n3607 10.6151
R13193 GND.n3609 GND.n3608 10.6151
R13194 GND.n3609 GND.n2515 10.6151
R13195 GND.n3626 GND.n2515 10.6151
R13196 GND.n3627 GND.n3626 10.6151
R13197 GND.n3638 GND.n3627 10.6151
R13198 GND.n3638 GND.n3637 10.6151
R13199 GND.n3637 GND.n3636 10.6151
R13200 GND.n3636 GND.n3635 10.6151
R13201 GND.n3635 GND.n3632 10.6151
R13202 GND.n3632 GND.n3631 10.6151
R13203 GND.n3631 GND.n3628 10.6151
R13204 GND.n3628 GND.n2499 10.6151
R13205 GND.n3664 GND.n2499 10.6151
R13206 GND.n3665 GND.n3664 10.6151
R13207 GND.n3668 GND.n3665 10.6151
R13208 GND.n3669 GND.n3668 10.6151
R13209 GND.n3670 GND.n3669 10.6151
R13210 GND.n3674 GND.n3670 10.6151
R13211 GND.n3674 GND.n3673 10.6151
R13212 GND.n3673 GND.n3672 10.6151
R13213 GND.n3672 GND.n2480 10.6151
R13214 GND.n3709 GND.n2480 10.6151
R13215 GND.n3710 GND.n3709 10.6151
R13216 GND.n3713 GND.n3710 10.6151
R13217 GND.n3714 GND.n3713 10.6151
R13218 GND.n3715 GND.n3714 10.6151
R13219 GND.n3721 GND.n3715 10.6151
R13220 GND.n3722 GND.n3721 10.6151
R13221 GND.n3782 GND.n3722 10.6151
R13222 GND.n3420 GND.n3419 10.6151
R13223 GND.n3420 GND.n3315 10.6151
R13224 GND.n3427 GND.n3426 10.6151
R13225 GND.n3428 GND.n3427 10.6151
R13226 GND.n3428 GND.n3310 10.6151
R13227 GND.n3434 GND.n3310 10.6151
R13228 GND.n3435 GND.n3434 10.6151
R13229 GND.n3436 GND.n3435 10.6151
R13230 GND.n3436 GND.n3308 10.6151
R13231 GND.n3442 GND.n3308 10.6151
R13232 GND.n3443 GND.n3442 10.6151
R13233 GND.n3444 GND.n3443 10.6151
R13234 GND.n3444 GND.n3306 10.6151
R13235 GND.n3450 GND.n3306 10.6151
R13236 GND.n3451 GND.n3450 10.6151
R13237 GND.n3452 GND.n3451 10.6151
R13238 GND.n3452 GND.n3304 10.6151
R13239 GND.n3458 GND.n3304 10.6151
R13240 GND.n3459 GND.n3458 10.6151
R13241 GND.n3460 GND.n3459 10.6151
R13242 GND.n3460 GND.n3302 10.6151
R13243 GND.n3466 GND.n3302 10.6151
R13244 GND.n3467 GND.n3466 10.6151
R13245 GND.n3468 GND.n3467 10.6151
R13246 GND.n3468 GND.n3300 10.6151
R13247 GND.n3300 GND.n3299 10.6151
R13248 GND.n3475 GND.n3299 10.6151
R13249 GND.n3359 GND.n3332 10.6151
R13250 GND.n3360 GND.n3359 10.6151
R13251 GND.n3361 GND.n3360 10.6151
R13252 GND.n3361 GND.n3330 10.6151
R13253 GND.n3367 GND.n3330 10.6151
R13254 GND.n3368 GND.n3367 10.6151
R13255 GND.n3369 GND.n3368 10.6151
R13256 GND.n3369 GND.n3328 10.6151
R13257 GND.n3375 GND.n3328 10.6151
R13258 GND.n3376 GND.n3375 10.6151
R13259 GND.n3377 GND.n3376 10.6151
R13260 GND.n3377 GND.n3326 10.6151
R13261 GND.n3383 GND.n3326 10.6151
R13262 GND.n3384 GND.n3383 10.6151
R13263 GND.n3385 GND.n3384 10.6151
R13264 GND.n3385 GND.n3324 10.6151
R13265 GND.n3391 GND.n3324 10.6151
R13266 GND.n3392 GND.n3391 10.6151
R13267 GND.n3393 GND.n3392 10.6151
R13268 GND.n3393 GND.n3322 10.6151
R13269 GND.n3399 GND.n3322 10.6151
R13270 GND.n3400 GND.n3399 10.6151
R13271 GND.n3401 GND.n3400 10.6151
R13272 GND.n3401 GND.n3320 10.6151
R13273 GND.n3407 GND.n3320 10.6151
R13274 GND.n3410 GND.n3409 10.6151
R13275 GND.n3410 GND.n3316 10.6151
R13276 GND.n4373 GND.n1967 10.6151
R13277 GND.n4368 GND.n1967 10.6151
R13278 GND.n4368 GND.n4367 10.6151
R13279 GND.n4367 GND.n4366 10.6151
R13280 GND.n4366 GND.n4363 10.6151
R13281 GND.n4363 GND.n4362 10.6151
R13282 GND.n4362 GND.n4359 10.6151
R13283 GND.n4359 GND.n4358 10.6151
R13284 GND.n4358 GND.n4355 10.6151
R13285 GND.n4355 GND.n4354 10.6151
R13286 GND.n4354 GND.n4351 10.6151
R13287 GND.n4351 GND.n4350 10.6151
R13288 GND.n4350 GND.n4347 10.6151
R13289 GND.n4347 GND.n4346 10.6151
R13290 GND.n4346 GND.n4343 10.6151
R13291 GND.n4343 GND.n4342 10.6151
R13292 GND.n4342 GND.n4339 10.6151
R13293 GND.n4339 GND.n4338 10.6151
R13294 GND.n4338 GND.n4335 10.6151
R13295 GND.n4335 GND.n4334 10.6151
R13296 GND.n4334 GND.n4331 10.6151
R13297 GND.n4331 GND.n4330 10.6151
R13298 GND.n4330 GND.n4327 10.6151
R13299 GND.n4327 GND.n4326 10.6151
R13300 GND.n4326 GND.n4323 10.6151
R13301 GND.n4321 GND.n4318 10.6151
R13302 GND.n4318 GND.n4317 10.6151
R13303 GND.n3354 GND.n1752 10.6151
R13304 GND.n4501 GND.n1752 10.6151
R13305 GND.n4501 GND.n4500 10.6151
R13306 GND.n4500 GND.n4499 10.6151
R13307 GND.n4499 GND.n1753 10.6151
R13308 GND.n2561 GND.n1753 10.6151
R13309 GND.n2561 GND.n1772 10.6151
R13310 GND.n4487 GND.n1772 10.6151
R13311 GND.n4487 GND.n4486 10.6151
R13312 GND.n4486 GND.n4485 10.6151
R13313 GND.n4485 GND.n1773 10.6151
R13314 GND.n3538 GND.n1773 10.6151
R13315 GND.n3538 GND.n1792 10.6151
R13316 GND.n4473 GND.n1792 10.6151
R13317 GND.n4473 GND.n4472 10.6151
R13318 GND.n4472 GND.n4471 10.6151
R13319 GND.n4471 GND.n1793 10.6151
R13320 GND.n3570 GND.n1793 10.6151
R13321 GND.n3570 GND.n1811 10.6151
R13322 GND.n4459 GND.n1811 10.6151
R13323 GND.n4459 GND.n4458 10.6151
R13324 GND.n4458 GND.n4457 10.6151
R13325 GND.n4457 GND.n1812 10.6151
R13326 GND.n3602 GND.n1812 10.6151
R13327 GND.n3602 GND.n1830 10.6151
R13328 GND.n4445 GND.n1830 10.6151
R13329 GND.n4445 GND.n4444 10.6151
R13330 GND.n4444 GND.n4443 10.6151
R13331 GND.n4443 GND.n1831 10.6151
R13332 GND.n2510 GND.n1831 10.6151
R13333 GND.n3642 GND.n2510 10.6151
R13334 GND.n3643 GND.n3642 10.6151
R13335 GND.n3644 GND.n3643 10.6151
R13336 GND.n3644 GND.n1859 10.6151
R13337 GND.n4424 GND.n1859 10.6151
R13338 GND.n4424 GND.n4423 10.6151
R13339 GND.n4423 GND.n4422 10.6151
R13340 GND.n4422 GND.n1860 10.6151
R13341 GND.n1885 GND.n1860 10.6151
R13342 GND.n4411 GND.n1885 10.6151
R13343 GND.n4411 GND.n4410 10.6151
R13344 GND.n4410 GND.n4409 10.6151
R13345 GND.n4409 GND.n1886 10.6151
R13346 GND.n3682 GND.n1886 10.6151
R13347 GND.n3682 GND.n3681 10.6151
R13348 GND.n3681 GND.n3680 10.6151
R13349 GND.n3680 GND.n3677 10.6151
R13350 GND.n3677 GND.n1923 10.6151
R13351 GND.n4390 GND.n1923 10.6151
R13352 GND.n4390 GND.n4389 10.6151
R13353 GND.n4389 GND.n4388 10.6151
R13354 GND.n4388 GND.n1924 10.6151
R13355 GND.n1947 GND.n1924 10.6151
R13356 GND.n4376 GND.n1947 10.6151
R13357 GND.n4376 GND.n4375 10.6151
R13358 GND.n4476 GND.n4475 10.5774
R13359 GND.n3666 GND.n1888 10.5774
R13360 GND.n89 GND.n73 10.4732
R13361 GND.n126 GND.n110 10.4732
R13362 GND.n158 GND.n142 10.4732
R13363 GND.n195 GND.n179 10.4732
R13364 GND.n20 GND.n4 10.4732
R13365 GND.n57 GND.n41 10.4732
R13366 GND.n522 GND.n506 10.4732
R13367 GND.n485 GND.n469 10.4732
R13368 GND.n591 GND.n575 10.4732
R13369 GND.n554 GND.n538 10.4732
R13370 GND.n661 GND.n645 10.4732
R13371 GND.n624 GND.n608 10.4732
R13372 GND.n325 GND.n309 10.4732
R13373 GND.n293 GND.n277 10.4732
R13374 GND.n261 GND.n245 10.4732
R13375 GND.n230 GND.n214 10.4732
R13376 GND.n452 GND.n436 10.4732
R13377 GND.n420 GND.n404 10.4732
R13378 GND.n388 GND.n372 10.4732
R13379 GND.n357 GND.n341 10.4732
R13380 GND.n2936 GND.t136 10.2469
R13381 GND.t127 GND.n2763 10.2469
R13382 GND.n5529 GND.t133 10.2469
R13383 GND.n849 GND.t158 10.2469
R13384 GND.n3297 GND.n3296 9.91636
R13385 GND.n3601 GND.n1824 9.91636
R13386 GND.n3622 GND.n2512 9.91636
R13387 GND.n3785 GND.n3784 9.91636
R13388 GND.n3806 GND.t97 9.91636
R13389 GND.n93 GND.n92 9.69747
R13390 GND.n130 GND.n129 9.69747
R13391 GND.n162 GND.n161 9.69747
R13392 GND.n199 GND.n198 9.69747
R13393 GND.n24 GND.n23 9.69747
R13394 GND.n61 GND.n60 9.69747
R13395 GND.n526 GND.n525 9.69747
R13396 GND.n489 GND.n488 9.69747
R13397 GND.n595 GND.n594 9.69747
R13398 GND.n558 GND.n557 9.69747
R13399 GND.n665 GND.n664 9.69747
R13400 GND.n628 GND.n627 9.69747
R13401 GND.n329 GND.n328 9.69747
R13402 GND.n297 GND.n296 9.69747
R13403 GND.n265 GND.n264 9.69747
R13404 GND.n234 GND.n233 9.69747
R13405 GND.n456 GND.n455 9.69747
R13406 GND.n424 GND.n423 9.69747
R13407 GND.n392 GND.n391 9.69747
R13408 GND.n361 GND.n360 9.69747
R13409 GND.t131 GND.n2720 9.58584
R13410 GND.n2281 GND.t120 9.58584
R13411 GND.n99 GND.n98 9.45567
R13412 GND.n136 GND.n135 9.45567
R13413 GND.n168 GND.n167 9.45567
R13414 GND.n205 GND.n204 9.45567
R13415 GND.n30 GND.n29 9.45567
R13416 GND.n67 GND.n66 9.45567
R13417 GND.n532 GND.n531 9.45567
R13418 GND.n495 GND.n494 9.45567
R13419 GND.n601 GND.n600 9.45567
R13420 GND.n564 GND.n563 9.45567
R13421 GND.n671 GND.n670 9.45567
R13422 GND.n634 GND.n633 9.45567
R13423 GND.n335 GND.n334 9.45567
R13424 GND.n303 GND.n302 9.45567
R13425 GND.n271 GND.n270 9.45567
R13426 GND.n240 GND.n239 9.45567
R13427 GND.n462 GND.n461 9.45567
R13428 GND.n430 GND.n429 9.45567
R13429 GND.n398 GND.n397 9.45567
R13430 GND.n367 GND.n366 9.45567
R13431 GND.n98 GND.n97 9.3005
R13432 GND.n71 GND.n70 9.3005
R13433 GND.n92 GND.n91 9.3005
R13434 GND.n90 GND.n89 9.3005
R13435 GND.n75 GND.n74 9.3005
R13436 GND.n84 GND.n83 9.3005
R13437 GND.n82 GND.n81 9.3005
R13438 GND.n135 GND.n134 9.3005
R13439 GND.n108 GND.n107 9.3005
R13440 GND.n129 GND.n128 9.3005
R13441 GND.n127 GND.n126 9.3005
R13442 GND.n112 GND.n111 9.3005
R13443 GND.n121 GND.n120 9.3005
R13444 GND.n119 GND.n118 9.3005
R13445 GND.n167 GND.n166 9.3005
R13446 GND.n140 GND.n139 9.3005
R13447 GND.n161 GND.n160 9.3005
R13448 GND.n159 GND.n158 9.3005
R13449 GND.n144 GND.n143 9.3005
R13450 GND.n153 GND.n152 9.3005
R13451 GND.n151 GND.n150 9.3005
R13452 GND.n204 GND.n203 9.3005
R13453 GND.n177 GND.n176 9.3005
R13454 GND.n198 GND.n197 9.3005
R13455 GND.n196 GND.n195 9.3005
R13456 GND.n181 GND.n180 9.3005
R13457 GND.n190 GND.n189 9.3005
R13458 GND.n188 GND.n187 9.3005
R13459 GND.n29 GND.n28 9.3005
R13460 GND.n2 GND.n1 9.3005
R13461 GND.n23 GND.n22 9.3005
R13462 GND.n21 GND.n20 9.3005
R13463 GND.n6 GND.n5 9.3005
R13464 GND.n15 GND.n14 9.3005
R13465 GND.n13 GND.n12 9.3005
R13466 GND.n66 GND.n65 9.3005
R13467 GND.n39 GND.n38 9.3005
R13468 GND.n60 GND.n59 9.3005
R13469 GND.n58 GND.n57 9.3005
R13470 GND.n43 GND.n42 9.3005
R13471 GND.n52 GND.n51 9.3005
R13472 GND.n50 GND.n49 9.3005
R13473 GND.n531 GND.n530 9.3005
R13474 GND.n504 GND.n503 9.3005
R13475 GND.n525 GND.n524 9.3005
R13476 GND.n523 GND.n522 9.3005
R13477 GND.n508 GND.n507 9.3005
R13478 GND.n517 GND.n516 9.3005
R13479 GND.n515 GND.n514 9.3005
R13480 GND.n494 GND.n493 9.3005
R13481 GND.n467 GND.n466 9.3005
R13482 GND.n488 GND.n487 9.3005
R13483 GND.n486 GND.n485 9.3005
R13484 GND.n471 GND.n470 9.3005
R13485 GND.n480 GND.n479 9.3005
R13486 GND.n478 GND.n477 9.3005
R13487 GND.n600 GND.n599 9.3005
R13488 GND.n573 GND.n572 9.3005
R13489 GND.n594 GND.n593 9.3005
R13490 GND.n592 GND.n591 9.3005
R13491 GND.n577 GND.n576 9.3005
R13492 GND.n586 GND.n585 9.3005
R13493 GND.n584 GND.n583 9.3005
R13494 GND.n563 GND.n562 9.3005
R13495 GND.n536 GND.n535 9.3005
R13496 GND.n557 GND.n556 9.3005
R13497 GND.n555 GND.n554 9.3005
R13498 GND.n540 GND.n539 9.3005
R13499 GND.n549 GND.n548 9.3005
R13500 GND.n547 GND.n546 9.3005
R13501 GND.n670 GND.n669 9.3005
R13502 GND.n643 GND.n642 9.3005
R13503 GND.n664 GND.n663 9.3005
R13504 GND.n662 GND.n661 9.3005
R13505 GND.n647 GND.n646 9.3005
R13506 GND.n656 GND.n655 9.3005
R13507 GND.n654 GND.n653 9.3005
R13508 GND.n633 GND.n632 9.3005
R13509 GND.n606 GND.n605 9.3005
R13510 GND.n627 GND.n626 9.3005
R13511 GND.n625 GND.n624 9.3005
R13512 GND.n610 GND.n609 9.3005
R13513 GND.n619 GND.n618 9.3005
R13514 GND.n617 GND.n616 9.3005
R13515 GND.n1687 GND.n1686 9.3005
R13516 GND.n1688 GND.n1685 9.3005
R13517 GND.n4536 GND.n1689 9.3005
R13518 GND.n4535 GND.n1690 9.3005
R13519 GND.n4534 GND.n1691 9.3005
R13520 GND.n1714 GND.n1692 9.3005
R13521 GND.n1715 GND.n1713 9.3005
R13522 GND.n4522 GND.n1716 9.3005
R13523 GND.n4521 GND.n1717 9.3005
R13524 GND.n4520 GND.n1718 9.3005
R13525 GND.n1739 GND.n1719 9.3005
R13526 GND.n1740 GND.n1738 9.3005
R13527 GND.n4508 GND.n1741 9.3005
R13528 GND.n4507 GND.n1742 9.3005
R13529 GND.n4506 GND.n1743 9.3005
R13530 GND.n1760 GND.n1744 9.3005
R13531 GND.n4494 GND.n1761 9.3005
R13532 GND.n4493 GND.n1762 9.3005
R13533 GND.n4492 GND.n1763 9.3005
R13534 GND.n1780 GND.n1764 9.3005
R13535 GND.n4480 GND.n1781 9.3005
R13536 GND.n4479 GND.n1782 9.3005
R13537 GND.n4478 GND.n1783 9.3005
R13538 GND.n1800 GND.n1784 9.3005
R13539 GND.n4466 GND.n1801 9.3005
R13540 GND.n4465 GND.n1802 9.3005
R13541 GND.n4464 GND.n1803 9.3005
R13542 GND.n1818 GND.n1804 9.3005
R13543 GND.n4452 GND.n1819 9.3005
R13544 GND.n4451 GND.n1820 9.3005
R13545 GND.n4450 GND.n1821 9.3005
R13546 GND.n1838 GND.n1822 9.3005
R13547 GND.n4438 GND.n1839 9.3005
R13548 GND.n4437 GND.n1840 9.3005
R13549 GND.n4436 GND.n1841 9.3005
R13550 GND.n1869 GND.n1842 9.3005
R13551 GND.n1872 GND.n1871 9.3005
R13552 GND.n1873 GND.n1868 9.3005
R13553 GND.n4417 GND.n1874 9.3005
R13554 GND.n4416 GND.n1875 9.3005
R13555 GND.n4415 GND.n1876 9.3005
R13556 GND.n2490 GND.n1877 9.3005
R13557 GND.n2493 GND.n2492 9.3005
R13558 GND.n2491 GND.n1911 9.3005
R13559 GND.n4397 GND.n1912 9.3005
R13560 GND.n4396 GND.n1913 9.3005
R13561 GND.n4395 GND.n1914 9.3005
R13562 GND.n3792 GND.n1915 9.3005
R13563 GND.n3794 GND.n3793 9.3005
R13564 GND.n3791 GND.n3790 9.3005
R13565 GND.n3799 GND.n3798 9.3005
R13566 GND.n3800 GND.n3789 9.3005
R13567 GND.n3804 GND.n3801 9.3005
R13568 GND.n3803 GND.n3802 9.3005
R13569 GND.n2457 GND.n2456 9.3005
R13570 GND.n3831 GND.n3830 9.3005
R13571 GND.n3832 GND.n2455 9.3005
R13572 GND.n3836 GND.n3833 9.3005
R13573 GND.n3835 GND.n3834 9.3005
R13574 GND.n2433 GND.n2432 9.3005
R13575 GND.n3865 GND.n3864 9.3005
R13576 GND.n3866 GND.n2431 9.3005
R13577 GND.n3868 GND.n3867 9.3005
R13578 GND.n2112 GND.n2111 9.3005
R13579 GND.n4236 GND.n4235 9.3005
R13580 GND.n1667 GND.n1579 9.3005
R13581 GND.n1221 GND.n1220 9.3005
R13582 GND.n4970 GND.n4969 9.3005
R13583 GND.n4971 GND.n1219 9.3005
R13584 GND.n4973 GND.n4972 9.3005
R13585 GND.n1215 GND.n1214 9.3005
R13586 GND.n4980 GND.n4979 9.3005
R13587 GND.n4981 GND.n1213 9.3005
R13588 GND.n4983 GND.n4982 9.3005
R13589 GND.n1209 GND.n1208 9.3005
R13590 GND.n4990 GND.n4989 9.3005
R13591 GND.n4991 GND.n1207 9.3005
R13592 GND.n4993 GND.n4992 9.3005
R13593 GND.n1203 GND.n1202 9.3005
R13594 GND.n5000 GND.n4999 9.3005
R13595 GND.n5001 GND.n1201 9.3005
R13596 GND.n5003 GND.n5002 9.3005
R13597 GND.n1197 GND.n1196 9.3005
R13598 GND.n5010 GND.n5009 9.3005
R13599 GND.n5011 GND.n1195 9.3005
R13600 GND.n5013 GND.n5012 9.3005
R13601 GND.n1191 GND.n1190 9.3005
R13602 GND.n5020 GND.n5019 9.3005
R13603 GND.n5021 GND.n1189 9.3005
R13604 GND.n5023 GND.n5022 9.3005
R13605 GND.n1185 GND.n1184 9.3005
R13606 GND.n5030 GND.n5029 9.3005
R13607 GND.n5031 GND.n1183 9.3005
R13608 GND.n5033 GND.n5032 9.3005
R13609 GND.n1179 GND.n1178 9.3005
R13610 GND.n5040 GND.n5039 9.3005
R13611 GND.n5041 GND.n1177 9.3005
R13612 GND.n5043 GND.n5042 9.3005
R13613 GND.n1173 GND.n1172 9.3005
R13614 GND.n5050 GND.n5049 9.3005
R13615 GND.n5051 GND.n1171 9.3005
R13616 GND.n5053 GND.n5052 9.3005
R13617 GND.n1167 GND.n1166 9.3005
R13618 GND.n5060 GND.n5059 9.3005
R13619 GND.n5061 GND.n1165 9.3005
R13620 GND.n5063 GND.n5062 9.3005
R13621 GND.n1161 GND.n1160 9.3005
R13622 GND.n5070 GND.n5069 9.3005
R13623 GND.n5071 GND.n1159 9.3005
R13624 GND.n5073 GND.n5072 9.3005
R13625 GND.n1155 GND.n1154 9.3005
R13626 GND.n5080 GND.n5079 9.3005
R13627 GND.n5081 GND.n1153 9.3005
R13628 GND.n5083 GND.n5082 9.3005
R13629 GND.n1149 GND.n1148 9.3005
R13630 GND.n5090 GND.n5089 9.3005
R13631 GND.n5091 GND.n1147 9.3005
R13632 GND.n5093 GND.n5092 9.3005
R13633 GND.n1143 GND.n1142 9.3005
R13634 GND.n5100 GND.n5099 9.3005
R13635 GND.n5101 GND.n1141 9.3005
R13636 GND.n5103 GND.n5102 9.3005
R13637 GND.n1137 GND.n1136 9.3005
R13638 GND.n5110 GND.n5109 9.3005
R13639 GND.n5111 GND.n1135 9.3005
R13640 GND.n5113 GND.n5112 9.3005
R13641 GND.n1131 GND.n1130 9.3005
R13642 GND.n5120 GND.n5119 9.3005
R13643 GND.n5121 GND.n1129 9.3005
R13644 GND.n5123 GND.n5122 9.3005
R13645 GND.n1125 GND.n1124 9.3005
R13646 GND.n5130 GND.n5129 9.3005
R13647 GND.n5131 GND.n1123 9.3005
R13648 GND.n5133 GND.n5132 9.3005
R13649 GND.n1119 GND.n1118 9.3005
R13650 GND.n5140 GND.n5139 9.3005
R13651 GND.n5141 GND.n1117 9.3005
R13652 GND.n5143 GND.n5142 9.3005
R13653 GND.n1113 GND.n1112 9.3005
R13654 GND.n5150 GND.n5149 9.3005
R13655 GND.n5151 GND.n1111 9.3005
R13656 GND.n5153 GND.n5152 9.3005
R13657 GND.n1107 GND.n1106 9.3005
R13658 GND.n5160 GND.n5159 9.3005
R13659 GND.n5161 GND.n1105 9.3005
R13660 GND.n5163 GND.n5162 9.3005
R13661 GND.n1101 GND.n1100 9.3005
R13662 GND.n5170 GND.n5169 9.3005
R13663 GND.n5171 GND.n1099 9.3005
R13664 GND.n5173 GND.n5172 9.3005
R13665 GND.n1095 GND.n1094 9.3005
R13666 GND.n5180 GND.n5179 9.3005
R13667 GND.n5181 GND.n1093 9.3005
R13668 GND.n5183 GND.n5182 9.3005
R13669 GND.n1089 GND.n1088 9.3005
R13670 GND.n5190 GND.n5189 9.3005
R13671 GND.n5191 GND.n1087 9.3005
R13672 GND.n5193 GND.n5192 9.3005
R13673 GND.n1083 GND.n1082 9.3005
R13674 GND.n5200 GND.n5199 9.3005
R13675 GND.n5201 GND.n1081 9.3005
R13676 GND.n5203 GND.n5202 9.3005
R13677 GND.n1077 GND.n1076 9.3005
R13678 GND.n5210 GND.n5209 9.3005
R13679 GND.n5211 GND.n1075 9.3005
R13680 GND.n5213 GND.n5212 9.3005
R13681 GND.n1071 GND.n1070 9.3005
R13682 GND.n5220 GND.n5219 9.3005
R13683 GND.n5221 GND.n1069 9.3005
R13684 GND.n5223 GND.n5222 9.3005
R13685 GND.n1065 GND.n1064 9.3005
R13686 GND.n5230 GND.n5229 9.3005
R13687 GND.n5231 GND.n1063 9.3005
R13688 GND.n5233 GND.n5232 9.3005
R13689 GND.n1059 GND.n1058 9.3005
R13690 GND.n5240 GND.n5239 9.3005
R13691 GND.n5241 GND.n1057 9.3005
R13692 GND.n5243 GND.n5242 9.3005
R13693 GND.n1053 GND.n1052 9.3005
R13694 GND.n5250 GND.n5249 9.3005
R13695 GND.n5251 GND.n1051 9.3005
R13696 GND.n5253 GND.n5252 9.3005
R13697 GND.n1047 GND.n1046 9.3005
R13698 GND.n5260 GND.n5259 9.3005
R13699 GND.n5261 GND.n1045 9.3005
R13700 GND.n5263 GND.n5262 9.3005
R13701 GND.n1041 GND.n1040 9.3005
R13702 GND.n5270 GND.n5269 9.3005
R13703 GND.n5271 GND.n1039 9.3005
R13704 GND.n5273 GND.n5272 9.3005
R13705 GND.n1035 GND.n1034 9.3005
R13706 GND.n5280 GND.n5279 9.3005
R13707 GND.n5281 GND.n1033 9.3005
R13708 GND.n5283 GND.n5282 9.3005
R13709 GND.n1029 GND.n1028 9.3005
R13710 GND.n5290 GND.n5289 9.3005
R13711 GND.n5291 GND.n1027 9.3005
R13712 GND.n5293 GND.n5292 9.3005
R13713 GND.n1023 GND.n1022 9.3005
R13714 GND.n5300 GND.n5299 9.3005
R13715 GND.n5301 GND.n1021 9.3005
R13716 GND.n5303 GND.n5302 9.3005
R13717 GND.n1017 GND.n1016 9.3005
R13718 GND.n5310 GND.n5309 9.3005
R13719 GND.n5311 GND.n1015 9.3005
R13720 GND.n5313 GND.n5312 9.3005
R13721 GND.n1011 GND.n1010 9.3005
R13722 GND.n5320 GND.n5319 9.3005
R13723 GND.n5321 GND.n1009 9.3005
R13724 GND.n5323 GND.n5322 9.3005
R13725 GND.n1005 GND.n1004 9.3005
R13726 GND.n5330 GND.n5329 9.3005
R13727 GND.n5331 GND.n1003 9.3005
R13728 GND.n5333 GND.n5332 9.3005
R13729 GND.n999 GND.n998 9.3005
R13730 GND.n5340 GND.n5339 9.3005
R13731 GND.n5341 GND.n997 9.3005
R13732 GND.n5343 GND.n5342 9.3005
R13733 GND.n993 GND.n992 9.3005
R13734 GND.n5350 GND.n5349 9.3005
R13735 GND.n5351 GND.n991 9.3005
R13736 GND.n5354 GND.n5353 9.3005
R13737 GND.n5352 GND.n987 9.3005
R13738 GND.n5360 GND.n986 9.3005
R13739 GND.n5362 GND.n5361 9.3005
R13740 GND.n982 GND.n981 9.3005
R13741 GND.n5371 GND.n5370 9.3005
R13742 GND.n5372 GND.n980 9.3005
R13743 GND.n5374 GND.n5373 9.3005
R13744 GND.n976 GND.n975 9.3005
R13745 GND.n5381 GND.n5380 9.3005
R13746 GND.n5382 GND.n974 9.3005
R13747 GND.n5384 GND.n5383 9.3005
R13748 GND.n970 GND.n969 9.3005
R13749 GND.n5391 GND.n5390 9.3005
R13750 GND.n5392 GND.n968 9.3005
R13751 GND.n5394 GND.n5393 9.3005
R13752 GND.n964 GND.n963 9.3005
R13753 GND.n5401 GND.n5400 9.3005
R13754 GND.n5402 GND.n962 9.3005
R13755 GND.n5404 GND.n5403 9.3005
R13756 GND.n958 GND.n957 9.3005
R13757 GND.n5411 GND.n5410 9.3005
R13758 GND.n5412 GND.n956 9.3005
R13759 GND.n5414 GND.n5413 9.3005
R13760 GND.n952 GND.n951 9.3005
R13761 GND.n5421 GND.n5420 9.3005
R13762 GND.n5422 GND.n950 9.3005
R13763 GND.n5424 GND.n5423 9.3005
R13764 GND.n946 GND.n945 9.3005
R13765 GND.n5431 GND.n5430 9.3005
R13766 GND.n5432 GND.n944 9.3005
R13767 GND.n5434 GND.n5433 9.3005
R13768 GND.n940 GND.n939 9.3005
R13769 GND.n5441 GND.n5440 9.3005
R13770 GND.n5442 GND.n938 9.3005
R13771 GND.n5444 GND.n5443 9.3005
R13772 GND.n934 GND.n933 9.3005
R13773 GND.n5451 GND.n5450 9.3005
R13774 GND.n5452 GND.n932 9.3005
R13775 GND.n5454 GND.n5453 9.3005
R13776 GND.n928 GND.n927 9.3005
R13777 GND.n5461 GND.n5460 9.3005
R13778 GND.n5462 GND.n926 9.3005
R13779 GND.n5464 GND.n5463 9.3005
R13780 GND.n922 GND.n921 9.3005
R13781 GND.n5471 GND.n5470 9.3005
R13782 GND.n5472 GND.n920 9.3005
R13783 GND.n5474 GND.n5473 9.3005
R13784 GND.n916 GND.n915 9.3005
R13785 GND.n5481 GND.n5480 9.3005
R13786 GND.n5482 GND.n914 9.3005
R13787 GND.n5484 GND.n5483 9.3005
R13788 GND.n910 GND.n909 9.3005
R13789 GND.n5491 GND.n5490 9.3005
R13790 GND.n5492 GND.n908 9.3005
R13791 GND.n5494 GND.n5493 9.3005
R13792 GND.n904 GND.n903 9.3005
R13793 GND.n5501 GND.n5500 9.3005
R13794 GND.n5502 GND.n902 9.3005
R13795 GND.n5504 GND.n5503 9.3005
R13796 GND.n898 GND.n897 9.3005
R13797 GND.n5511 GND.n5510 9.3005
R13798 GND.n5512 GND.n896 9.3005
R13799 GND.n5515 GND.n5514 9.3005
R13800 GND.n5513 GND.n892 9.3005
R13801 GND.n5521 GND.n891 9.3005
R13802 GND.n5523 GND.n5522 9.3005
R13803 GND.n5364 GND.n5363 9.3005
R13804 GND.n2165 GND.n2164 9.3005
R13805 GND.n2163 GND.n2120 9.3005
R13806 GND.n2162 GND.n2161 9.3005
R13807 GND.n2158 GND.n2122 9.3005
R13808 GND.n2155 GND.n2154 9.3005
R13809 GND.n2153 GND.n2123 9.3005
R13810 GND.n2152 GND.n2151 9.3005
R13811 GND.n2148 GND.n2124 9.3005
R13812 GND.n2145 GND.n2144 9.3005
R13813 GND.n2143 GND.n2125 9.3005
R13814 GND.n2142 GND.n2141 9.3005
R13815 GND.n2138 GND.n2126 9.3005
R13816 GND.n2135 GND.n2134 9.3005
R13817 GND.n2133 GND.n2127 9.3005
R13818 GND.n2132 GND.n2131 9.3005
R13819 GND.n2128 GND.n2009 9.3005
R13820 GND.n4311 GND.n2008 9.3005
R13821 GND.n2384 GND.n2003 9.3005
R13822 GND.n2386 GND.n2385 9.3005
R13823 GND.n2389 GND.n2383 9.3005
R13824 GND.n2390 GND.n2382 9.3005
R13825 GND.n2393 GND.n2381 9.3005
R13826 GND.n2394 GND.n2380 9.3005
R13827 GND.n2397 GND.n2379 9.3005
R13828 GND.n2398 GND.n2378 9.3005
R13829 GND.n2401 GND.n2377 9.3005
R13830 GND.n2402 GND.n2376 9.3005
R13831 GND.n2405 GND.n2375 9.3005
R13832 GND.n2406 GND.n2374 9.3005
R13833 GND.n2409 GND.n2373 9.3005
R13834 GND.n2410 GND.n2372 9.3005
R13835 GND.n2166 GND.n2117 9.3005
R13836 GND.n2167 GND.n2113 9.3005
R13837 GND.n3985 GND.n3984 9.3005
R13838 GND.n3986 GND.n2369 9.3005
R13839 GND.n3990 GND.n3987 9.3005
R13840 GND.n3989 GND.n3988 9.3005
R13841 GND.n2348 GND.n2347 9.3005
R13842 GND.n4010 GND.n4009 9.3005
R13843 GND.n4011 GND.n2346 9.3005
R13844 GND.n4015 GND.n4012 9.3005
R13845 GND.n4014 GND.n4013 9.3005
R13846 GND.n2325 GND.n2324 9.3005
R13847 GND.n4034 GND.n4033 9.3005
R13848 GND.n4035 GND.n2323 9.3005
R13849 GND.n4039 GND.n4036 9.3005
R13850 GND.n4038 GND.n4037 9.3005
R13851 GND.n2302 GND.n2301 9.3005
R13852 GND.n4059 GND.n4058 9.3005
R13853 GND.n4060 GND.n2300 9.3005
R13854 GND.n4065 GND.n4061 9.3005
R13855 GND.n4064 GND.n4063 9.3005
R13856 GND.n4062 GND.n2272 9.3005
R13857 GND.n4168 GND.n4167 9.3005
R13858 GND.n4169 GND.n2243 9.3005
R13859 GND.n4173 GND.n4170 9.3005
R13860 GND.n4172 GND.n4171 9.3005
R13861 GND.n866 GND.n865 9.3005
R13862 GND.n5547 GND.n5546 9.3005
R13863 GND.n5548 GND.n864 9.3005
R13864 GND.n5550 GND.n5549 9.3005
R13865 GND.n844 GND.n843 9.3005
R13866 GND.n5564 GND.n5563 9.3005
R13867 GND.n5565 GND.n842 9.3005
R13868 GND.n5567 GND.n5566 9.3005
R13869 GND.n825 GND.n824 9.3005
R13870 GND.n5581 GND.n5580 9.3005
R13871 GND.n5582 GND.n823 9.3005
R13872 GND.n5584 GND.n5583 9.3005
R13873 GND.n808 GND.n807 9.3005
R13874 GND.n5599 GND.n5598 9.3005
R13875 GND.n5600 GND.n806 9.3005
R13876 GND.n5603 GND.n5601 9.3005
R13877 GND.n5602 GND.n745 9.3005
R13878 GND.n2371 GND.n2370 9.3005
R13879 GND.n2245 GND.n2244 9.3005
R13880 GND.n3074 GND.n3026 9.3005
R13881 GND.n3029 GND.n3027 9.3005
R13882 GND.n3068 GND.n3030 9.3005
R13883 GND.n3067 GND.n3031 9.3005
R13884 GND.n3066 GND.n3032 9.3005
R13885 GND.n3035 GND.n3033 9.3005
R13886 GND.n3059 GND.n3036 9.3005
R13887 GND.n3058 GND.n3037 9.3005
R13888 GND.n3057 GND.n3038 9.3005
R13889 GND.n3043 GND.n3039 9.3005
R13890 GND.n3053 GND.n3044 9.3005
R13891 GND.n3052 GND.n3045 9.3005
R13892 GND.n3051 GND.n3046 9.3005
R13893 GND.n3049 GND.n3048 9.3005
R13894 GND.n3047 GND.n2617 9.3005
R13895 GND.n2615 GND.n2614 9.3005
R13896 GND.n3191 GND.n3190 9.3005
R13897 GND.n3192 GND.n2613 9.3005
R13898 GND.n3203 GND.n3193 9.3005
R13899 GND.n3202 GND.n3194 9.3005
R13900 GND.n3201 GND.n3195 9.3005
R13901 GND.n3198 GND.n3197 9.3005
R13902 GND.n3196 GND.n1642 9.3005
R13903 GND.n4555 GND.n1643 9.3005
R13904 GND.n4554 GND.n1644 9.3005
R13905 GND.n4553 GND.n1645 9.3005
R13906 GND.n1674 GND.n1646 9.3005
R13907 GND.n1675 GND.n1673 9.3005
R13908 GND.n4543 GND.n1676 9.3005
R13909 GND.n4542 GND.n1677 9.3005
R13910 GND.n4541 GND.n1678 9.3005
R13911 GND.n1700 GND.n1679 9.3005
R13912 GND.n1701 GND.n1699 9.3005
R13913 GND.n4529 GND.n1702 9.3005
R13914 GND.n4528 GND.n1703 9.3005
R13915 GND.n4527 GND.n1704 9.3005
R13916 GND.n1727 GND.n1705 9.3005
R13917 GND.n1728 GND.n1726 9.3005
R13918 GND.n4515 GND.n1729 9.3005
R13919 GND.n4514 GND.n1730 9.3005
R13920 GND.n4513 GND.n1731 9.3005
R13921 GND.n2549 GND.n1732 9.3005
R13922 GND.n2551 GND.n2550 9.3005
R13923 GND.n2548 GND.n2547 9.3005
R13924 GND.n2556 GND.n2555 9.3005
R13925 GND.n2557 GND.n2546 9.3005
R13926 GND.n2559 GND.n2558 9.3005
R13927 GND.n2544 GND.n2543 9.3005
R13928 GND.n3521 GND.n3520 9.3005
R13929 GND.n3522 GND.n2542 9.3005
R13930 GND.n3534 GND.n3523 9.3005
R13931 GND.n3533 GND.n3524 9.3005
R13932 GND.n3532 GND.n3525 9.3005
R13933 GND.n3529 GND.n3526 9.3005
R13934 GND.n3528 GND.n3527 9.3005
R13935 GND.n2526 GND.n2525 9.3005
R13936 GND.n3587 GND.n3586 9.3005
R13937 GND.n3588 GND.n2524 9.3005
R13938 GND.n3599 GND.n3589 9.3005
R13939 GND.n3598 GND.n3590 9.3005
R13940 GND.n3597 GND.n3591 9.3005
R13941 GND.n3594 GND.n3593 9.3005
R13942 GND.n3592 GND.n1848 9.3005
R13943 GND.n4431 GND.n1849 9.3005
R13944 GND.n4430 GND.n1850 9.3005
R13945 GND.n4429 GND.n1851 9.3005
R13946 GND.n1893 GND.n1852 9.3005
R13947 GND.n1895 GND.n1894 9.3005
R13948 GND.n1899 GND.n1898 9.3005
R13949 GND.n1900 GND.n1892 9.3005
R13950 GND.n4404 GND.n1901 9.3005
R13951 GND.n4403 GND.n1902 9.3005
R13952 GND.n4402 GND.n1903 9.3005
R13953 GND.n1932 GND.n1904 9.3005
R13954 GND.n1935 GND.n1934 9.3005
R13955 GND.n1936 GND.n1931 9.3005
R13956 GND.n4383 GND.n1937 9.3005
R13957 GND.n4382 GND.n1938 9.3005
R13958 GND.n4381 GND.n1939 9.3005
R13959 GND.n2466 GND.n1940 9.3005
R13960 GND.n2468 GND.n2467 9.3005
R13961 GND.n2465 GND.n2464 9.3005
R13962 GND.n3820 GND.n3819 9.3005
R13963 GND.n3821 GND.n2463 9.3005
R13964 GND.n3825 GND.n3822 9.3005
R13965 GND.n3824 GND.n3823 9.3005
R13966 GND.n2442 GND.n2441 9.3005
R13967 GND.n3856 GND.n3855 9.3005
R13968 GND.n3857 GND.n2440 9.3005
R13969 GND.n3859 GND.n3858 9.3005
R13970 GND.n2427 GND.n2426 9.3005
R13971 GND.n3875 GND.n3874 9.3005
R13972 GND.n3876 GND.n2425 9.3005
R13973 GND.n3878 GND.n3877 9.3005
R13974 GND.n2423 GND.n2422 9.3005
R13975 GND.n3907 GND.n3906 9.3005
R13976 GND.n3908 GND.n2421 9.3005
R13977 GND.n3910 GND.n3909 9.3005
R13978 GND.n2419 GND.n2418 9.3005
R13979 GND.n3922 GND.n3921 9.3005
R13980 GND.n3923 GND.n2417 9.3005
R13981 GND.n3975 GND.n3924 9.3005
R13982 GND.n3974 GND.n3925 9.3005
R13983 GND.n3973 GND.n3926 9.3005
R13984 GND.n3929 GND.n3927 9.3005
R13985 GND.n3969 GND.n3930 9.3005
R13986 GND.n3968 GND.n3931 9.3005
R13987 GND.n3967 GND.n3932 9.3005
R13988 GND.n3935 GND.n3933 9.3005
R13989 GND.n3963 GND.n3936 9.3005
R13990 GND.n3962 GND.n3937 9.3005
R13991 GND.n3961 GND.n3938 9.3005
R13992 GND.n3941 GND.n3939 9.3005
R13993 GND.n3957 GND.n3942 9.3005
R13994 GND.n3956 GND.n3943 9.3005
R13995 GND.n3955 GND.n3944 9.3005
R13996 GND.n3947 GND.n3945 9.3005
R13997 GND.n3951 GND.n3948 9.3005
R13998 GND.n3950 GND.n3949 9.3005
R13999 GND.n2261 GND.n2260 9.3005
R14000 GND.n4147 GND.n4146 9.3005
R14001 GND.n4157 GND.n4149 9.3005
R14002 GND.n4156 GND.n4150 9.3005
R14003 GND.n4153 GND.n4152 9.3005
R14004 GND.n4151 GND.n884 9.3005
R14005 GND.n5533 GND.n885 9.3005
R14006 GND.n5532 GND.n886 9.3005
R14007 GND.n5531 GND.n887 9.3005
R14008 GND.n890 GND.n888 9.3005
R14009 GND.n5525 GND.n5524 9.3005
R14010 GND.n4772 GND.n4771 9.3005
R14011 GND.n4773 GND.n1412 9.3005
R14012 GND.n4776 GND.n1411 9.3005
R14013 GND.n4777 GND.n1410 9.3005
R14014 GND.n4780 GND.n1409 9.3005
R14015 GND.n4781 GND.n1408 9.3005
R14016 GND.n4784 GND.n1407 9.3005
R14017 GND.n4785 GND.n1406 9.3005
R14018 GND.n4788 GND.n1405 9.3005
R14019 GND.n4789 GND.n1404 9.3005
R14020 GND.n4792 GND.n1403 9.3005
R14021 GND.n4793 GND.n1402 9.3005
R14022 GND.n4796 GND.n1401 9.3005
R14023 GND.n4797 GND.n1400 9.3005
R14024 GND.n4800 GND.n1399 9.3005
R14025 GND.n4801 GND.n1398 9.3005
R14026 GND.n4804 GND.n1397 9.3005
R14027 GND.n4806 GND.n1394 9.3005
R14028 GND.n4809 GND.n1393 9.3005
R14029 GND.n4810 GND.n1392 9.3005
R14030 GND.n4813 GND.n1391 9.3005
R14031 GND.n4814 GND.n1390 9.3005
R14032 GND.n4817 GND.n1389 9.3005
R14033 GND.n4818 GND.n1388 9.3005
R14034 GND.n4821 GND.n1387 9.3005
R14035 GND.n4822 GND.n1386 9.3005
R14036 GND.n4825 GND.n1385 9.3005
R14037 GND.n4826 GND.n1384 9.3005
R14038 GND.n4829 GND.n1383 9.3005
R14039 GND.n4831 GND.n1382 9.3005
R14040 GND.n4832 GND.n1381 9.3005
R14041 GND.n4833 GND.n1380 9.3005
R14042 GND.n4834 GND.n1379 9.3005
R14043 GND.n4770 GND.n1417 9.3005
R14044 GND.n4769 GND.n4768 9.3005
R14045 GND.n2906 GND.n2903 9.3005
R14046 GND.n2908 GND.n2907 9.3005
R14047 GND.n2809 GND.n2808 9.3005
R14048 GND.n2918 GND.n2917 9.3005
R14049 GND.n2919 GND.n2807 9.3005
R14050 GND.n2921 GND.n2920 9.3005
R14051 GND.n2796 GND.n2795 9.3005
R14052 GND.n2931 GND.n2930 9.3005
R14053 GND.n2932 GND.n2794 9.3005
R14054 GND.n2934 GND.n2933 9.3005
R14055 GND.n2770 GND.n2769 9.3005
R14056 GND.n2947 GND.n2946 9.3005
R14057 GND.n2948 GND.n2768 9.3005
R14058 GND.n2952 GND.n2949 9.3005
R14059 GND.n2951 GND.n2950 9.3005
R14060 GND.n2747 GND.n2746 9.3005
R14061 GND.n2984 GND.n2983 9.3005
R14062 GND.n2985 GND.n2745 9.3005
R14063 GND.n2988 GND.n2986 9.3005
R14064 GND.n2987 GND.n2683 9.3005
R14065 GND.n3108 GND.n3107 9.3005
R14066 GND.n2663 GND.n2662 9.3005
R14067 GND.n3129 GND.n3128 9.3005
R14068 GND.n3130 GND.n2661 9.3005
R14069 GND.n3134 GND.n3131 9.3005
R14070 GND.n3133 GND.n3132 9.3005
R14071 GND.n2644 GND.n2643 9.3005
R14072 GND.n3154 GND.n3153 9.3005
R14073 GND.n3155 GND.n2642 9.3005
R14074 GND.n3159 GND.n3156 9.3005
R14075 GND.n3158 GND.n3157 9.3005
R14076 GND.n2623 GND.n2622 9.3005
R14077 GND.n3180 GND.n3179 9.3005
R14078 GND.n3181 GND.n2621 9.3005
R14079 GND.n3183 GND.n3182 9.3005
R14080 GND.n2597 GND.n2596 9.3005
R14081 GND.n3220 GND.n3219 9.3005
R14082 GND.n3221 GND.n2595 9.3005
R14083 GND.n3223 GND.n3222 9.3005
R14084 GND.n1532 GND.n1531 9.3005
R14085 GND.n4683 GND.n4682 9.3005
R14086 GND.n2905 GND.n2904 9.3005
R14087 GND.n3109 GND.n3106 9.3005
R14088 GND.n2787 GND.n2777 9.3005
R14089 GND.n2786 GND.n2778 9.3005
R14090 GND.n2780 GND.n2779 9.3005
R14091 GND.n2782 GND.n2781 9.3005
R14092 GND.n2735 GND.n2734 9.3005
R14093 GND.n2994 GND.n2993 9.3005
R14094 GND.n2995 GND.n2733 9.3005
R14095 GND.n2997 GND.n2996 9.3005
R14096 GND.n2788 GND.n2776 9.3005
R14097 GND.n4841 GND.n1347 9.3005
R14098 GND.n4842 GND.n1346 9.3005
R14099 GND.n4843 GND.n1345 9.3005
R14100 GND.n1344 GND.n1340 9.3005
R14101 GND.n4849 GND.n1339 9.3005
R14102 GND.n4850 GND.n1338 9.3005
R14103 GND.n4851 GND.n1337 9.3005
R14104 GND.n1336 GND.n1332 9.3005
R14105 GND.n4857 GND.n1331 9.3005
R14106 GND.n4858 GND.n1330 9.3005
R14107 GND.n4859 GND.n1329 9.3005
R14108 GND.n1328 GND.n1324 9.3005
R14109 GND.n4865 GND.n1323 9.3005
R14110 GND.n4866 GND.n1322 9.3005
R14111 GND.n4867 GND.n1321 9.3005
R14112 GND.n1320 GND.n1316 9.3005
R14113 GND.n4873 GND.n1315 9.3005
R14114 GND.n4874 GND.n1314 9.3005
R14115 GND.n4875 GND.n1313 9.3005
R14116 GND.n1312 GND.n1308 9.3005
R14117 GND.n4881 GND.n1307 9.3005
R14118 GND.n4882 GND.n1306 9.3005
R14119 GND.n4883 GND.n1305 9.3005
R14120 GND.n1304 GND.n1300 9.3005
R14121 GND.n4889 GND.n1299 9.3005
R14122 GND.n4890 GND.n1298 9.3005
R14123 GND.n4891 GND.n1297 9.3005
R14124 GND.n1296 GND.n1292 9.3005
R14125 GND.n4897 GND.n1291 9.3005
R14126 GND.n4898 GND.n1290 9.3005
R14127 GND.n4899 GND.n1289 9.3005
R14128 GND.n1288 GND.n1284 9.3005
R14129 GND.n4905 GND.n1283 9.3005
R14130 GND.n4906 GND.n1282 9.3005
R14131 GND.n4907 GND.n1281 9.3005
R14132 GND.n1280 GND.n1276 9.3005
R14133 GND.n4913 GND.n1275 9.3005
R14134 GND.n4914 GND.n1274 9.3005
R14135 GND.n4915 GND.n1273 9.3005
R14136 GND.n1272 GND.n1268 9.3005
R14137 GND.n4921 GND.n1267 9.3005
R14138 GND.n4922 GND.n1266 9.3005
R14139 GND.n4923 GND.n1265 9.3005
R14140 GND.n1264 GND.n1260 9.3005
R14141 GND.n4929 GND.n1259 9.3005
R14142 GND.n4930 GND.n1258 9.3005
R14143 GND.n4931 GND.n1257 9.3005
R14144 GND.n1256 GND.n1252 9.3005
R14145 GND.n4937 GND.n1251 9.3005
R14146 GND.n4938 GND.n1250 9.3005
R14147 GND.n4939 GND.n1249 9.3005
R14148 GND.n1248 GND.n1244 9.3005
R14149 GND.n4945 GND.n1243 9.3005
R14150 GND.n4946 GND.n1242 9.3005
R14151 GND.n4947 GND.n1241 9.3005
R14152 GND.n1240 GND.n1236 9.3005
R14153 GND.n4953 GND.n1235 9.3005
R14154 GND.n4954 GND.n1234 9.3005
R14155 GND.n4955 GND.n1233 9.3005
R14156 GND.n1232 GND.n1228 9.3005
R14157 GND.n4961 GND.n1227 9.3005
R14158 GND.n4962 GND.n1226 9.3005
R14159 GND.n4963 GND.n1225 9.3005
R14160 GND.n2775 GND.n1348 9.3005
R14161 GND.n3914 GND.n3913 9.3005
R14162 GND.n2360 GND.n2359 9.3005
R14163 GND.n3995 GND.n3994 9.3005
R14164 GND.n3996 GND.n2357 9.3005
R14165 GND.n3999 GND.n3998 9.3005
R14166 GND.n3997 GND.n2358 9.3005
R14167 GND.n2338 GND.n2337 9.3005
R14168 GND.n4020 GND.n4019 9.3005
R14169 GND.n4021 GND.n2335 9.3005
R14170 GND.n4024 GND.n4023 9.3005
R14171 GND.n4022 GND.n2336 9.3005
R14172 GND.n2314 GND.n2313 9.3005
R14173 GND.n4044 GND.n4043 9.3005
R14174 GND.n4045 GND.n2311 9.3005
R14175 GND.n4048 GND.n4047 9.3005
R14176 GND.n4046 GND.n2312 9.3005
R14177 GND.n2287 GND.n2286 9.3005
R14178 GND.n4070 GND.n4069 9.3005
R14179 GND.n4071 GND.n2284 9.3005
R14180 GND.n4073 GND.n4072 9.3005
R14181 GND.n4074 GND.n2283 9.3005
R14182 GND.n4078 GND.n4077 9.3005
R14183 GND.n4079 GND.n2282 9.3005
R14184 GND.n4081 GND.n4080 9.3005
R14185 GND.n676 GND.n674 9.3005
R14186 GND.n3916 GND.n3915 9.3005
R14187 GND.n5757 GND.n5756 9.3005
R14188 GND.n5755 GND.n675 9.3005
R14189 GND.n5754 GND.n5753 9.3005
R14190 GND.n5752 GND.n680 9.3005
R14191 GND.n5751 GND.n5750 9.3005
R14192 GND.n5749 GND.n681 9.3005
R14193 GND.n5748 GND.n5747 9.3005
R14194 GND.n5746 GND.n685 9.3005
R14195 GND.n5745 GND.n5744 9.3005
R14196 GND.n5743 GND.n686 9.3005
R14197 GND.n5742 GND.n5741 9.3005
R14198 GND.n5740 GND.n690 9.3005
R14199 GND.n5739 GND.n5738 9.3005
R14200 GND.n5737 GND.n691 9.3005
R14201 GND.n5736 GND.n5735 9.3005
R14202 GND.n5734 GND.n695 9.3005
R14203 GND.n5733 GND.n5732 9.3005
R14204 GND.n5731 GND.n696 9.3005
R14205 GND.n5730 GND.n5729 9.3005
R14206 GND.n5728 GND.n700 9.3005
R14207 GND.n5727 GND.n5726 9.3005
R14208 GND.n5725 GND.n701 9.3005
R14209 GND.n5724 GND.n5723 9.3005
R14210 GND.n5722 GND.n705 9.3005
R14211 GND.n5721 GND.n5720 9.3005
R14212 GND.n5719 GND.n706 9.3005
R14213 GND.n5718 GND.n5717 9.3005
R14214 GND.n5648 GND.n5607 9.3005
R14215 GND.n5647 GND.n5646 9.3005
R14216 GND.n5645 GND.n5608 9.3005
R14217 GND.n5644 GND.n5643 9.3005
R14218 GND.n5642 GND.n5613 9.3005
R14219 GND.n5641 GND.n5640 9.3005
R14220 GND.n5639 GND.n5614 9.3005
R14221 GND.n5638 GND.n5637 9.3005
R14222 GND.n5636 GND.n5619 9.3005
R14223 GND.n5635 GND.n5634 9.3005
R14224 GND.n5633 GND.n5620 9.3005
R14225 GND.n5632 GND.n5631 9.3005
R14226 GND.n5630 GND.n5625 9.3005
R14227 GND.n5629 GND.n5628 9.3005
R14228 GND.n713 GND.n710 9.3005
R14229 GND.n5716 GND.n5715 9.3005
R14230 GND.n5650 GND.n5649 9.3005
R14231 GND.n5709 GND.n744 9.3005
R14232 GND.n5708 GND.n5707 9.3005
R14233 GND.n5706 GND.n746 9.3005
R14234 GND.n5705 GND.n5704 9.3005
R14235 GND.n5703 GND.n751 9.3005
R14236 GND.n5702 GND.n5701 9.3005
R14237 GND.n5700 GND.n752 9.3005
R14238 GND.n5699 GND.n5698 9.3005
R14239 GND.n5697 GND.n757 9.3005
R14240 GND.n5696 GND.n5695 9.3005
R14241 GND.n5694 GND.n758 9.3005
R14242 GND.n5693 GND.n5692 9.3005
R14243 GND.n5691 GND.n763 9.3005
R14244 GND.n5690 GND.n5689 9.3005
R14245 GND.n5688 GND.n764 9.3005
R14246 GND.n5686 GND.n5685 9.3005
R14247 GND.n5684 GND.n771 9.3005
R14248 GND.n5683 GND.n5682 9.3005
R14249 GND.n5681 GND.n772 9.3005
R14250 GND.n5680 GND.n5679 9.3005
R14251 GND.n5678 GND.n777 9.3005
R14252 GND.n5677 GND.n5676 9.3005
R14253 GND.n5675 GND.n778 9.3005
R14254 GND.n5674 GND.n5673 9.3005
R14255 GND.n5672 GND.n783 9.3005
R14256 GND.n5671 GND.n5670 9.3005
R14257 GND.n5669 GND.n784 9.3005
R14258 GND.n5668 GND.n5667 9.3005
R14259 GND.n5666 GND.n789 9.3005
R14260 GND.n5665 GND.n5664 9.3005
R14261 GND.n5663 GND.n790 9.3005
R14262 GND.n5662 GND.n5661 9.3005
R14263 GND.n5660 GND.n797 9.3005
R14264 GND.n5659 GND.n5658 9.3005
R14265 GND.n5711 GND.n5710 9.3005
R14266 GND.n3980 GND.n2115 9.3005
R14267 GND.n4228 GND.n2173 9.3005
R14268 GND.n4227 GND.n2174 9.3005
R14269 GND.n4226 GND.n2175 9.3005
R14270 GND.n2354 GND.n2176 9.3005
R14271 GND.n4222 GND.n2181 9.3005
R14272 GND.n4221 GND.n2182 9.3005
R14273 GND.n4220 GND.n2183 9.3005
R14274 GND.n2331 GND.n2184 9.3005
R14275 GND.n4216 GND.n2189 9.3005
R14276 GND.n4215 GND.n2190 9.3005
R14277 GND.n4214 GND.n2191 9.3005
R14278 GND.n2318 GND.n2192 9.3005
R14279 GND.n4210 GND.n2197 9.3005
R14280 GND.n4209 GND.n2198 9.3005
R14281 GND.n4208 GND.n2199 9.3005
R14282 GND.n4052 GND.n2200 9.3005
R14283 GND.n4204 GND.n2205 9.3005
R14284 GND.n4203 GND.n2206 9.3005
R14285 GND.n4202 GND.n2207 9.3005
R14286 GND.n2268 GND.n2208 9.3005
R14287 GND.n4198 GND.n2213 9.3005
R14288 GND.n4197 GND.n2214 9.3005
R14289 GND.n4196 GND.n2215 9.3005
R14290 GND.n2279 GND.n2216 9.3005
R14291 GND.n4192 GND.n2221 9.3005
R14292 GND.n4191 GND.n2222 9.3005
R14293 GND.n4190 GND.n2223 9.3005
R14294 GND.n4106 GND.n2224 9.3005
R14295 GND.n4186 GND.n2229 9.3005
R14296 GND.n4185 GND.n2230 9.3005
R14297 GND.n4184 GND.n2231 9.3005
R14298 GND.n2237 GND.n2232 9.3005
R14299 GND.n4180 GND.n2236 9.3005
R14300 GND.n4179 GND.n4178 9.3005
R14301 GND.n875 GND.n873 9.3005
R14302 GND.n5542 GND.n5541 9.3005
R14303 GND.n878 GND.n874 9.3005
R14304 GND.n877 GND.n876 9.3005
R14305 GND.n854 GND.n852 9.3005
R14306 GND.n5559 GND.n5558 9.3005
R14307 GND.n857 GND.n853 9.3005
R14308 GND.n856 GND.n855 9.3005
R14309 GND.n834 GND.n832 9.3005
R14310 GND.n5576 GND.n5575 9.3005
R14311 GND.n837 GND.n833 9.3005
R14312 GND.n836 GND.n835 9.3005
R14313 GND.n816 GND.n814 9.3005
R14314 GND.n5594 GND.n5593 9.3005
R14315 GND.n817 GND.n815 9.3005
R14316 GND.n802 GND.n801 9.3005
R14317 GND.n5654 GND.n5653 9.3005
R14318 GND.n4232 GND.n2114 9.3005
R14319 GND.n4230 GND.n2115 9.3005
R14320 GND.n4229 GND.n4228 9.3005
R14321 GND.n4227 GND.n2172 9.3005
R14322 GND.n4226 GND.n4225 9.3005
R14323 GND.n4224 GND.n2176 9.3005
R14324 GND.n4223 GND.n4222 9.3005
R14325 GND.n4221 GND.n2180 9.3005
R14326 GND.n4220 GND.n4219 9.3005
R14327 GND.n4218 GND.n2184 9.3005
R14328 GND.n4217 GND.n4216 9.3005
R14329 GND.n4215 GND.n2188 9.3005
R14330 GND.n4214 GND.n4213 9.3005
R14331 GND.n4212 GND.n2192 9.3005
R14332 GND.n4211 GND.n4210 9.3005
R14333 GND.n4209 GND.n2196 9.3005
R14334 GND.n4208 GND.n4207 9.3005
R14335 GND.n4206 GND.n2200 9.3005
R14336 GND.n4205 GND.n4204 9.3005
R14337 GND.n4203 GND.n2204 9.3005
R14338 GND.n4202 GND.n4201 9.3005
R14339 GND.n4200 GND.n2208 9.3005
R14340 GND.n4199 GND.n4198 9.3005
R14341 GND.n4197 GND.n2212 9.3005
R14342 GND.n4196 GND.n4195 9.3005
R14343 GND.n4194 GND.n2216 9.3005
R14344 GND.n4193 GND.n4192 9.3005
R14345 GND.n4191 GND.n2220 9.3005
R14346 GND.n4190 GND.n4189 9.3005
R14347 GND.n4188 GND.n2224 9.3005
R14348 GND.n4187 GND.n4186 9.3005
R14349 GND.n4185 GND.n2228 9.3005
R14350 GND.n4184 GND.n4183 9.3005
R14351 GND.n4182 GND.n2232 9.3005
R14352 GND.n4181 GND.n4180 9.3005
R14353 GND.n4179 GND.n879 9.3005
R14354 GND.n5538 GND.n875 9.3005
R14355 GND.n5541 GND.n5540 9.3005
R14356 GND.n5539 GND.n878 9.3005
R14357 GND.n877 GND.n858 9.3005
R14358 GND.n5555 GND.n854 9.3005
R14359 GND.n5558 GND.n5557 9.3005
R14360 GND.n5556 GND.n857 9.3005
R14361 GND.n856 GND.n838 9.3005
R14362 GND.n5572 GND.n834 9.3005
R14363 GND.n5575 GND.n5574 9.3005
R14364 GND.n5573 GND.n837 9.3005
R14365 GND.n836 GND.n818 9.3005
R14366 GND.n5589 GND.n816 9.3005
R14367 GND.n5593 GND.n5592 9.3005
R14368 GND.n5591 GND.n817 9.3005
R14369 GND.n801 GND.n800 9.3005
R14370 GND.n5655 GND.n5654 9.3005
R14371 GND.n4232 GND.n4231 9.3005
R14372 GND.n4301 GND.n4300 9.3005
R14373 GND.n2047 GND.n2046 9.3005
R14374 GND.n4295 GND.n4294 9.3005
R14375 GND.n4293 GND.n4292 9.3005
R14376 GND.n2057 GND.n2056 9.3005
R14377 GND.n4287 GND.n4286 9.3005
R14378 GND.n4285 GND.n4284 9.3005
R14379 GND.n2065 GND.n2064 9.3005
R14380 GND.n4279 GND.n4278 9.3005
R14381 GND.n4277 GND.n4276 9.3005
R14382 GND.n2075 GND.n2074 9.3005
R14383 GND.n4271 GND.n4270 9.3005
R14384 GND.n4269 GND.n4268 9.3005
R14385 GND.n2083 GND.n2082 9.3005
R14386 GND.n4259 GND.n4258 9.3005
R14387 GND.n4257 GND.n2085 9.3005
R14388 GND.n4303 GND.n4302 9.3005
R14389 GND.n2079 GND.n2078 9.3005
R14390 GND.n4273 GND.n4272 9.3005
R14391 GND.n4275 GND.n4274 9.3005
R14392 GND.n2071 GND.n2070 9.3005
R14393 GND.n4281 GND.n4280 9.3005
R14394 GND.n4283 GND.n4282 9.3005
R14395 GND.n2061 GND.n2060 9.3005
R14396 GND.n4289 GND.n4288 9.3005
R14397 GND.n4291 GND.n4290 9.3005
R14398 GND.n2053 GND.n2052 9.3005
R14399 GND.n4297 GND.n4296 9.3005
R14400 GND.n4299 GND.n4298 9.3005
R14401 GND.n2043 GND.n2042 9.3005
R14402 GND.n4305 GND.n4304 9.3005
R14403 GND.n4306 GND.n2041 9.3005
R14404 GND.n4267 GND.n4266 9.3005
R14405 GND.n4261 GND.n4260 9.3005
R14406 GND.n4256 GND.n4255 9.3005
R14407 GND.n4254 GND.n2089 9.3005
R14408 GND.n4253 GND.n4252 9.3005
R14409 GND.n4251 GND.n2091 9.3005
R14410 GND.n4250 GND.n4249 9.3005
R14411 GND.n4248 GND.n2095 9.3005
R14412 GND.n4247 GND.n4246 9.3005
R14413 GND.n4245 GND.n2096 9.3005
R14414 GND.n4244 GND.n4243 9.3005
R14415 GND.n4242 GND.n2103 9.3005
R14416 GND.n3269 GND.n2583 9.3005
R14417 GND.n3275 GND.n3274 9.3005
R14418 GND.n3276 GND.n2580 9.3005
R14419 GND.n3278 GND.n3277 9.3005
R14420 GND.n3279 GND.n2579 9.3005
R14421 GND.n3283 GND.n3282 9.3005
R14422 GND.n3284 GND.n2578 9.3005
R14423 GND.n3286 GND.n3285 9.3005
R14424 GND.n3289 GND.n2577 9.3005
R14425 GND.n3291 GND.n3290 9.3005
R14426 GND.n3292 GND.n2572 9.3005
R14427 GND.n3294 GND.n3293 9.3005
R14428 GND.n3295 GND.n2571 9.3005
R14429 GND.n3483 GND.n3482 9.3005
R14430 GND.n3484 GND.n2570 9.3005
R14431 GND.n3486 GND.n3485 9.3005
R14432 GND.n2566 GND.n2564 9.3005
R14433 GND.n3513 GND.n3512 9.3005
R14434 GND.n3511 GND.n2565 9.3005
R14435 GND.n3510 GND.n3509 9.3005
R14436 GND.n3508 GND.n2567 9.3005
R14437 GND.n3507 GND.n3506 9.3005
R14438 GND.n2535 GND.n2534 9.3005
R14439 GND.n3552 GND.n3551 9.3005
R14440 GND.n3553 GND.n2532 9.3005
R14441 GND.n3566 GND.n3565 9.3005
R14442 GND.n3564 GND.n2533 9.3005
R14443 GND.n3563 GND.n3562 9.3005
R14444 GND.n3561 GND.n3554 9.3005
R14445 GND.n3560 GND.n3559 9.3005
R14446 GND.n2519 GND.n2518 9.3005
R14447 GND.n3615 GND.n3614 9.3005
R14448 GND.n3616 GND.n2516 9.3005
R14449 GND.n3620 GND.n3619 9.3005
R14450 GND.n3618 GND.n2517 9.3005
R14451 GND.n3617 GND.n2506 9.3005
R14452 GND.n2505 GND.n2504 9.3005
R14453 GND.n3652 GND.n3651 9.3005
R14454 GND.n3653 GND.n2502 9.3005
R14455 GND.n3659 GND.n3658 9.3005
R14456 GND.n3657 GND.n2503 9.3005
R14457 GND.n3656 GND.n3655 9.3005
R14458 GND.n2487 GND.n2486 9.3005
R14459 GND.n3688 GND.n3687 9.3005
R14460 GND.n3689 GND.n2484 9.3005
R14461 GND.n3704 GND.n3703 9.3005
R14462 GND.n3702 GND.n2485 9.3005
R14463 GND.n3701 GND.n3700 9.3005
R14464 GND.n3699 GND.n3690 9.3005
R14465 GND.n3698 GND.n3697 9.3005
R14466 GND.n3696 GND.n3695 9.3005
R14467 GND.n2476 GND.n2475 9.3005
R14468 GND.n3809 GND.n3808 9.3005
R14469 GND.n3810 GND.n2473 9.3005
R14470 GND.n3813 GND.n3812 9.3005
R14471 GND.n3811 GND.n2474 9.3005
R14472 GND.n2449 GND.n2448 9.3005
R14473 GND.n3841 GND.n3840 9.3005
R14474 GND.n3842 GND.n2446 9.3005
R14475 GND.n3850 GND.n3849 9.3005
R14476 GND.n3848 GND.n2447 9.3005
R14477 GND.n3847 GND.n3846 9.3005
R14478 GND.n3845 GND.n3843 9.3005
R14479 GND.n2105 GND.n2104 9.3005
R14480 GND.n4241 GND.n4240 9.3005
R14481 GND.n3268 GND.n3267 9.3005
R14482 GND.n3263 GND.n2584 9.3005
R14483 GND.n3260 GND.n3259 9.3005
R14484 GND.n3258 GND.n2585 9.3005
R14485 GND.n3257 GND.n3256 9.3005
R14486 GND.n3250 GND.n2586 9.3005
R14487 GND.n3247 GND.n3246 9.3005
R14488 GND.n3245 GND.n2587 9.3005
R14489 GND.n3244 GND.n3243 9.3005
R14490 GND.n3240 GND.n2588 9.3005
R14491 GND.n3266 GND.n3265 9.3005
R14492 GND.n3016 GND.n3015 9.3005
R14493 GND.n3017 GND.n2723 9.3005
R14494 GND.n3019 GND.n3018 9.3005
R14495 GND.n2674 GND.n2673 9.3005
R14496 GND.n3114 GND.n3113 9.3005
R14497 GND.n3115 GND.n2671 9.3005
R14498 GND.n3118 GND.n3117 9.3005
R14499 GND.n3116 GND.n2672 9.3005
R14500 GND.n2654 GND.n2653 9.3005
R14501 GND.n3139 GND.n3138 9.3005
R14502 GND.n3140 GND.n2651 9.3005
R14503 GND.n3143 GND.n3142 9.3005
R14504 GND.n3141 GND.n2652 9.3005
R14505 GND.n2634 GND.n2633 9.3005
R14506 GND.n3164 GND.n3163 9.3005
R14507 GND.n3165 GND.n2631 9.3005
R14508 GND.n3171 GND.n3170 9.3005
R14509 GND.n3169 GND.n2632 9.3005
R14510 GND.n3168 GND.n3167 9.3005
R14511 GND.n2608 GND.n2606 9.3005
R14512 GND.n3212 GND.n3211 9.3005
R14513 GND.n3210 GND.n2607 9.3005
R14514 GND.n3209 GND.n3208 9.3005
R14515 GND.n2609 GND.n2590 9.3005
R14516 GND.n3232 GND.n2589 9.3005
R14517 GND.n3234 GND.n3233 9.3005
R14518 GND.n3237 GND.n3236 9.3005
R14519 GND.n1625 GND.n1624 9.3005
R14520 GND.n4589 GND.n4588 9.3005
R14521 GND.n4591 GND.n4590 9.3005
R14522 GND.n1615 GND.n1614 9.3005
R14523 GND.n4597 GND.n4596 9.3005
R14524 GND.n4599 GND.n4598 9.3005
R14525 GND.n1607 GND.n1606 9.3005
R14526 GND.n4605 GND.n4604 9.3005
R14527 GND.n4607 GND.n4606 9.3005
R14528 GND.n1599 GND.n1598 9.3005
R14529 GND.n4613 GND.n4612 9.3005
R14530 GND.n4615 GND.n4614 9.3005
R14531 GND.n1591 GND.n1590 9.3005
R14532 GND.n4621 GND.n4620 9.3005
R14533 GND.n4623 GND.n4622 9.3005
R14534 GND.n1587 GND.n1585 9.3005
R14535 GND.n4626 GND.n1580 9.3005
R14536 GND.n4625 GND.n4624 9.3005
R14537 GND.n1586 GND.n1584 9.3005
R14538 GND.n4619 GND.n4618 9.3005
R14539 GND.n4617 GND.n4616 9.3005
R14540 GND.n1595 GND.n1594 9.3005
R14541 GND.n4611 GND.n4610 9.3005
R14542 GND.n4609 GND.n4608 9.3005
R14543 GND.n1603 GND.n1602 9.3005
R14544 GND.n4603 GND.n4602 9.3005
R14545 GND.n4601 GND.n4600 9.3005
R14546 GND.n1611 GND.n1610 9.3005
R14547 GND.n4595 GND.n4594 9.3005
R14548 GND.n4593 GND.n4592 9.3005
R14549 GND.n1621 GND.n1620 9.3005
R14550 GND.n4587 GND.n4586 9.3005
R14551 GND.n4628 GND.n4627 9.3005
R14552 GND.n4661 GND.n1547 9.3005
R14553 GND.n4663 GND.n4662 9.3005
R14554 GND.n4664 GND.n1546 9.3005
R14555 GND.n4666 GND.n4665 9.3005
R14556 GND.n4667 GND.n1542 9.3005
R14557 GND.n4669 GND.n4668 9.3005
R14558 GND.n4670 GND.n1541 9.3005
R14559 GND.n4672 GND.n4671 9.3005
R14560 GND.n4673 GND.n1537 9.3005
R14561 GND.n4675 GND.n4674 9.3005
R14562 GND.n4676 GND.n1536 9.3005
R14563 GND.n4678 GND.n4677 9.3005
R14564 GND.n4679 GND.n1533 9.3005
R14565 GND.n4681 GND.n4680 9.3005
R14566 GND.n4657 GND.n1556 9.3005
R14567 GND.n4656 GND.n4655 9.3005
R14568 GND.n4654 GND.n1557 9.3005
R14569 GND.n4653 GND.n4652 9.3005
R14570 GND.n4651 GND.n1561 9.3005
R14571 GND.n4650 GND.n4649 9.3005
R14572 GND.n4648 GND.n1562 9.3005
R14573 GND.n4647 GND.n4646 9.3005
R14574 GND.n4645 GND.n1566 9.3005
R14575 GND.n4644 GND.n4643 9.3005
R14576 GND.n4642 GND.n1567 9.3005
R14577 GND.n4641 GND.n4640 9.3005
R14578 GND.n4639 GND.n1571 9.3005
R14579 GND.n4638 GND.n4637 9.3005
R14580 GND.n4636 GND.n1572 9.3005
R14581 GND.n4635 GND.n4634 9.3005
R14582 GND.n4633 GND.n1578 9.3005
R14583 GND.n4632 GND.n4631 9.3005
R14584 GND.n4659 GND.n4658 9.3005
R14585 GND.n4763 GND.n1422 9.3005
R14586 GND.n4762 GND.n1423 9.3005
R14587 GND.n2912 GND.n1424 9.3005
R14588 GND.n4758 GND.n1429 9.3005
R14589 GND.n4757 GND.n1430 9.3005
R14590 GND.n4756 GND.n1431 9.3005
R14591 GND.n2925 GND.n1432 9.3005
R14592 GND.n4752 GND.n1437 9.3005
R14593 GND.n4751 GND.n1438 9.3005
R14594 GND.n4750 GND.n1439 9.3005
R14595 GND.n2938 GND.n1440 9.3005
R14596 GND.n4746 GND.n1445 9.3005
R14597 GND.n4745 GND.n1446 9.3005
R14598 GND.n4744 GND.n1447 9.3005
R14599 GND.n2753 GND.n1448 9.3005
R14600 GND.n4740 GND.n1453 9.3005
R14601 GND.n4739 GND.n1454 9.3005
R14602 GND.n4738 GND.n1455 9.3005
R14603 GND.n2740 GND.n1456 9.3005
R14604 GND.n4734 GND.n1461 9.3005
R14605 GND.n4733 GND.n1462 9.3005
R14606 GND.n4732 GND.n1463 9.3005
R14607 GND.n3099 GND.n1464 9.3005
R14608 GND.n4728 GND.n1469 9.3005
R14609 GND.n4727 GND.n1470 9.3005
R14610 GND.n4726 GND.n1471 9.3005
R14611 GND.n2710 GND.n1472 9.3005
R14612 GND.n4722 GND.n1477 9.3005
R14613 GND.n4721 GND.n1478 9.3005
R14614 GND.n4720 GND.n1479 9.3005
R14615 GND.n2678 GND.n1480 9.3005
R14616 GND.n4716 GND.n1485 9.3005
R14617 GND.n4715 GND.n1486 9.3005
R14618 GND.n4714 GND.n1487 9.3005
R14619 GND.n3122 GND.n1488 9.3005
R14620 GND.n4710 GND.n1493 9.3005
R14621 GND.n4709 GND.n1494 9.3005
R14622 GND.n4708 GND.n1495 9.3005
R14623 GND.n3149 GND.n1496 9.3005
R14624 GND.n4704 GND.n1501 9.3005
R14625 GND.n4703 GND.n1502 9.3005
R14626 GND.n4702 GND.n1503 9.3005
R14627 GND.n2629 GND.n1504 9.3005
R14628 GND.n4698 GND.n1509 9.3005
R14629 GND.n4697 GND.n1510 9.3005
R14630 GND.n4696 GND.n1511 9.3005
R14631 GND.n2603 GND.n1512 9.3005
R14632 GND.n4692 GND.n1517 9.3005
R14633 GND.n4691 GND.n1518 9.3005
R14634 GND.n4690 GND.n1519 9.3005
R14635 GND.n3228 GND.n1520 9.3005
R14636 GND.n3227 GND.n1523 9.3005
R14637 GND.n4764 GND.n1421 9.3005
R14638 GND.n4763 GND.n1420 9.3005
R14639 GND.n4762 GND.n4761 9.3005
R14640 GND.n4760 GND.n1424 9.3005
R14641 GND.n4759 GND.n4758 9.3005
R14642 GND.n4757 GND.n1428 9.3005
R14643 GND.n4756 GND.n4755 9.3005
R14644 GND.n4754 GND.n1432 9.3005
R14645 GND.n4753 GND.n4752 9.3005
R14646 GND.n4751 GND.n1436 9.3005
R14647 GND.n4750 GND.n4749 9.3005
R14648 GND.n4748 GND.n1440 9.3005
R14649 GND.n4747 GND.n4746 9.3005
R14650 GND.n4745 GND.n1444 9.3005
R14651 GND.n4744 GND.n4743 9.3005
R14652 GND.n4742 GND.n1448 9.3005
R14653 GND.n4741 GND.n4740 9.3005
R14654 GND.n4739 GND.n1452 9.3005
R14655 GND.n4738 GND.n4737 9.3005
R14656 GND.n4736 GND.n1456 9.3005
R14657 GND.n4735 GND.n4734 9.3005
R14658 GND.n4733 GND.n1460 9.3005
R14659 GND.n4732 GND.n4731 9.3005
R14660 GND.n4730 GND.n1464 9.3005
R14661 GND.n4729 GND.n4728 9.3005
R14662 GND.n4727 GND.n1468 9.3005
R14663 GND.n4726 GND.n4725 9.3005
R14664 GND.n4724 GND.n1472 9.3005
R14665 GND.n4723 GND.n4722 9.3005
R14666 GND.n4721 GND.n1476 9.3005
R14667 GND.n4720 GND.n4719 9.3005
R14668 GND.n4718 GND.n1480 9.3005
R14669 GND.n4717 GND.n4716 9.3005
R14670 GND.n4715 GND.n1484 9.3005
R14671 GND.n4714 GND.n4713 9.3005
R14672 GND.n4712 GND.n1488 9.3005
R14673 GND.n4711 GND.n4710 9.3005
R14674 GND.n4709 GND.n1492 9.3005
R14675 GND.n4708 GND.n4707 9.3005
R14676 GND.n4706 GND.n1496 9.3005
R14677 GND.n4705 GND.n4704 9.3005
R14678 GND.n4703 GND.n1500 9.3005
R14679 GND.n4702 GND.n4701 9.3005
R14680 GND.n4700 GND.n1504 9.3005
R14681 GND.n4699 GND.n4698 9.3005
R14682 GND.n4697 GND.n1508 9.3005
R14683 GND.n4696 GND.n4695 9.3005
R14684 GND.n4694 GND.n1512 9.3005
R14685 GND.n4693 GND.n4692 9.3005
R14686 GND.n4691 GND.n1516 9.3005
R14687 GND.n4690 GND.n4689 9.3005
R14688 GND.n4688 GND.n1520 9.3005
R14689 GND.n4687 GND.n1523 9.3005
R14690 GND.n4765 GND.n4764 9.3005
R14691 GND.n2868 GND.n2867 9.3005
R14692 GND.n2866 GND.n2823 9.3005
R14693 GND.n2865 GND.n2864 9.3005
R14694 GND.n2861 GND.n2826 9.3005
R14695 GND.n2860 GND.n2859 9.3005
R14696 GND.n2858 GND.n2827 9.3005
R14697 GND.n2857 GND.n2856 9.3005
R14698 GND.n2853 GND.n2830 9.3005
R14699 GND.n2852 GND.n2851 9.3005
R14700 GND.n2850 GND.n2831 9.3005
R14701 GND.n2849 GND.n2848 9.3005
R14702 GND.n2845 GND.n2834 9.3005
R14703 GND.n2844 GND.n2843 9.3005
R14704 GND.n2842 GND.n2835 9.3005
R14705 GND.n2841 GND.n2840 9.3005
R14706 GND.n2869 GND.n2819 9.3005
R14707 GND.n2871 GND.n2870 9.3005
R14708 GND.n2875 GND.n2817 9.3005
R14709 GND.n2900 GND.n2899 9.3005
R14710 GND.n2898 GND.n2818 9.3005
R14711 GND.n2897 GND.n2896 9.3005
R14712 GND.n2895 GND.n2876 9.3005
R14713 GND.n2894 GND.n2893 9.3005
R14714 GND.n2892 GND.n2879 9.3005
R14715 GND.n2891 GND.n2890 9.3005
R14716 GND.n2889 GND.n2880 9.3005
R14717 GND.n2888 GND.n2887 9.3005
R14718 GND.n2886 GND.n2883 9.3005
R14719 GND.n2885 GND.n2884 9.3005
R14720 GND.n2760 GND.n2759 9.3005
R14721 GND.n2957 GND.n2956 9.3005
R14722 GND.n2958 GND.n2757 9.3005
R14723 GND.n2975 GND.n2974 9.3005
R14724 GND.n2973 GND.n2758 9.3005
R14725 GND.n2972 GND.n2971 9.3005
R14726 GND.n2970 GND.n2959 9.3005
R14727 GND.n2969 GND.n2968 9.3005
R14728 GND.n2967 GND.n2727 9.3005
R14729 GND.n3006 GND.n2726 9.3005
R14730 GND.n3008 GND.n3007 9.3005
R14731 GND.n3009 GND.n2725 9.3005
R14732 GND.n3011 GND.n3010 9.3005
R14733 GND.n2874 GND.n2873 9.3005
R14734 GND.n3014 GND.n2724 9.3005
R14735 GND.n334 GND.n333 9.3005
R14736 GND.n307 GND.n306 9.3005
R14737 GND.n328 GND.n327 9.3005
R14738 GND.n326 GND.n325 9.3005
R14739 GND.n311 GND.n310 9.3005
R14740 GND.n320 GND.n319 9.3005
R14741 GND.n318 GND.n317 9.3005
R14742 GND.n302 GND.n301 9.3005
R14743 GND.n275 GND.n274 9.3005
R14744 GND.n296 GND.n295 9.3005
R14745 GND.n294 GND.n293 9.3005
R14746 GND.n279 GND.n278 9.3005
R14747 GND.n288 GND.n287 9.3005
R14748 GND.n286 GND.n285 9.3005
R14749 GND.n270 GND.n269 9.3005
R14750 GND.n243 GND.n242 9.3005
R14751 GND.n264 GND.n263 9.3005
R14752 GND.n262 GND.n261 9.3005
R14753 GND.n247 GND.n246 9.3005
R14754 GND.n256 GND.n255 9.3005
R14755 GND.n254 GND.n253 9.3005
R14756 GND.n239 GND.n238 9.3005
R14757 GND.n212 GND.n211 9.3005
R14758 GND.n233 GND.n232 9.3005
R14759 GND.n231 GND.n230 9.3005
R14760 GND.n216 GND.n215 9.3005
R14761 GND.n225 GND.n224 9.3005
R14762 GND.n223 GND.n222 9.3005
R14763 GND.n461 GND.n460 9.3005
R14764 GND.n434 GND.n433 9.3005
R14765 GND.n455 GND.n454 9.3005
R14766 GND.n453 GND.n452 9.3005
R14767 GND.n438 GND.n437 9.3005
R14768 GND.n447 GND.n446 9.3005
R14769 GND.n445 GND.n444 9.3005
R14770 GND.n429 GND.n428 9.3005
R14771 GND.n402 GND.n401 9.3005
R14772 GND.n423 GND.n422 9.3005
R14773 GND.n421 GND.n420 9.3005
R14774 GND.n406 GND.n405 9.3005
R14775 GND.n415 GND.n414 9.3005
R14776 GND.n413 GND.n412 9.3005
R14777 GND.n397 GND.n396 9.3005
R14778 GND.n370 GND.n369 9.3005
R14779 GND.n391 GND.n390 9.3005
R14780 GND.n389 GND.n388 9.3005
R14781 GND.n374 GND.n373 9.3005
R14782 GND.n383 GND.n382 9.3005
R14783 GND.n381 GND.n380 9.3005
R14784 GND.n366 GND.n365 9.3005
R14785 GND.n339 GND.n338 9.3005
R14786 GND.n360 GND.n359 9.3005
R14787 GND.n358 GND.n357 9.3005
R14788 GND.n343 GND.n342 9.3005
R14789 GND.n352 GND.n351 9.3005
R14790 GND.n350 GND.n349 9.3005
R14791 GND.n4482 GND.n1778 9.25531
R14792 GND.n4462 GND.n1806 9.25531
R14793 GND.n3629 GND.n1856 9.25531
R14794 GND.n3685 GND.n3684 9.25531
R14795 GND.n3041 GND.t125 8.92478
R14796 GND.t140 GND.n2333 8.92478
R14797 GND.n96 GND.n71 8.92171
R14798 GND.n133 GND.n108 8.92171
R14799 GND.n165 GND.n140 8.92171
R14800 GND.n202 GND.n177 8.92171
R14801 GND.n27 GND.n2 8.92171
R14802 GND.n64 GND.n39 8.92171
R14803 GND.n529 GND.n504 8.92171
R14804 GND.n492 GND.n467 8.92171
R14805 GND.n598 GND.n573 8.92171
R14806 GND.n561 GND.n536 8.92171
R14807 GND.n668 GND.n643 8.92171
R14808 GND.n631 GND.n606 8.92171
R14809 GND.n332 GND.n307 8.92171
R14810 GND.n300 GND.n275 8.92171
R14811 GND.n268 GND.n243 8.92171
R14812 GND.n237 GND.n212 8.92171
R14813 GND.n459 GND.n434 8.92171
R14814 GND.n427 GND.n402 8.92171
R14815 GND.n395 GND.n370 8.92171
R14816 GND.n364 GND.n339 8.92171
R14817 GND.n1966 GND.n1948 8.72777
R14818 GND.n4489 GND.n1769 8.59425
R14819 GND.n4455 GND.n1814 8.59425
R14820 GND.n3646 GND.n2508 8.59425
R14821 GND.n2483 GND.n2482 8.59425
R14822 GND.n5758 GND.n5757 8.41206
R14823 GND.n2724 GND.n209 8.41206
R14824 GND.n3555 GND.t22 8.26372
R14825 GND.t9 GND.n1845 8.26372
R14826 GND.n97 GND.n69 8.14595
R14827 GND.n134 GND.n106 8.14595
R14828 GND.n166 GND.n138 8.14595
R14829 GND.n203 GND.n175 8.14595
R14830 GND.n28 GND.n0 8.14595
R14831 GND.n65 GND.n37 8.14595
R14832 GND.n530 GND.n502 8.14595
R14833 GND.n493 GND.n465 8.14595
R14834 GND.n599 GND.n571 8.14595
R14835 GND.n562 GND.n534 8.14595
R14836 GND.n669 GND.n641 8.14595
R14837 GND.n632 GND.n604 8.14595
R14838 GND.n333 GND.n305 8.14595
R14839 GND.n301 GND.n273 8.14595
R14840 GND.n269 GND.n241 8.14595
R14841 GND.n238 GND.n210 8.14595
R14842 GND.n460 GND.n432 8.14595
R14843 GND.n428 GND.n400 8.14595
R14844 GND.n396 GND.n368 8.14595
R14845 GND.n365 GND.n337 8.14595
R14846 GND.n4497 GND.t70 7.93319
R14847 GND.t70 GND.n4496 7.93319
R14848 GND.n2560 GND.t35 7.93319
R14849 GND.n4490 GND.n4489 7.93319
R14850 GND.t8 GND.n4468 7.93319
R14851 GND.n4455 GND.n4454 7.93319
R14852 GND.n3647 GND.n3646 7.93319
R14853 GND.t6 GND.n3661 7.93319
R14854 GND.n3706 GND.n2483 7.93319
R14855 GND.n5715 GND.n713 7.75808
R14856 GND.n4586 GND.n1620 7.75808
R14857 GND.n2870 GND.n2869 7.75808
R14858 GND.n4266 GND.n4261 7.75808
R14859 GND.n3351 GND.n3350 7.30353
R14860 GND.n1965 GND.n1964 7.30353
R14861 GND.n2538 GND.n1778 7.27213
R14862 GND.n3569 GND.n1806 7.27213
R14863 GND.n3629 GND.n1862 7.27213
R14864 GND.n3684 GND.n2489 7.27213
R14865 GND.t50 GND.n1920 7.27213
R14866 GND.t32 GND.n3717 7.27213
R14867 GND.n209 GND.n208 6.93127
R14868 GND.n5758 GND.n673 6.93127
R14869 GND.n207 GND.n137 6.61257
R14870 GND.n603 GND.n533 6.61257
R14871 GND.n3480 GND.n3297 6.61108
R14872 GND.n4496 GND.n1758 6.61108
R14873 GND.n4448 GND.n1824 6.61108
R14874 GND.n3623 GND.n3622 6.61108
R14875 GND.n3711 GND.n1926 6.61108
R14876 GND.n3729 GND.n3725 6.5566
R14877 GND.n3315 GND.n3314 6.5566
R14878 GND.n3409 GND.n3408 6.5566
R14879 GND.n4322 GND.n4321 6.5566
R14880 GND.n4454 GND.t22 6.28055
R14881 GND.n3647 GND.t9 6.28055
R14882 GND.n5687 GND.n5686 6.20656
R14883 GND.n4805 GND.n4804 6.20656
R14884 GND.n4475 GND.n1789 5.95002
R14885 GND.n4469 GND.n1795 5.95002
R14886 GND.n3662 GND.n1879 5.95002
R14887 GND.n3666 GND.n1882 5.95002
R14888 GND.n99 GND.n69 5.81868
R14889 GND.n136 GND.n106 5.81868
R14890 GND.n168 GND.n138 5.81868
R14891 GND.n205 GND.n175 5.81868
R14892 GND.n30 GND.n0 5.81868
R14893 GND.n67 GND.n37 5.81868
R14894 GND.n532 GND.n502 5.81868
R14895 GND.n495 GND.n465 5.81868
R14896 GND.n601 GND.n571 5.81868
R14897 GND.n564 GND.n534 5.81868
R14898 GND.n671 GND.n641 5.81868
R14899 GND.n634 GND.n604 5.81868
R14900 GND.n335 GND.n305 5.81868
R14901 GND.n303 GND.n273 5.81868
R14902 GND.n271 GND.n241 5.81868
R14903 GND.n240 GND.n210 5.81868
R14904 GND.n462 GND.n432 5.81868
R14905 GND.n430 GND.n400 5.81868
R14906 GND.n398 GND.n368 5.81868
R14907 GND.n367 GND.n337 5.81868
R14908 GND.n4314 GND.n2002 5.62001
R14909 GND.n3419 GND.n1554 5.62001
R14910 GND.n3316 GND.n1554 5.62001
R14911 GND.n4317 GND.n4314 5.62001
R14912 GND.t0 GND.n1721 5.61949
R14913 GND.n3815 GND.t17 5.61949
R14914 GND.n4246 GND.n2099 5.4308
R14915 GND.n3255 GND.n2585 5.4308
R14916 GND.n3612 GND.n3611 5.28896
R14917 GND.n4441 GND.n4440 5.28896
R14918 GND.n3719 GND.n1942 5.28896
R14919 GND.n3784 GND.t79 5.28896
R14920 GND.n97 GND.n96 5.04292
R14921 GND.n134 GND.n133 5.04292
R14922 GND.n166 GND.n165 5.04292
R14923 GND.n203 GND.n202 5.04292
R14924 GND.n28 GND.n27 5.04292
R14925 GND.n65 GND.n64 5.04292
R14926 GND.n530 GND.n529 5.04292
R14927 GND.n493 GND.n492 5.04292
R14928 GND.n599 GND.n598 5.04292
R14929 GND.n562 GND.n561 5.04292
R14930 GND.n669 GND.n668 5.04292
R14931 GND.n632 GND.n631 5.04292
R14932 GND.n333 GND.n332 5.04292
R14933 GND.n301 GND.n300 5.04292
R14934 GND.n269 GND.n268 5.04292
R14935 GND.n238 GND.n237 5.04292
R14936 GND.n460 GND.n459 5.04292
R14937 GND.n428 GND.n427 5.04292
R14938 GND.n396 GND.n395 5.04292
R14939 GND.n365 GND.n364 5.04292
R14940 GND.t39 GND.n2811 4.95843
R14941 GND.n4371 GND.t97 4.95843
R14942 GND.n5596 GND.t63 4.95843
R14943 GND.n208 GND.n68 4.7699
R14944 GND.n673 GND.n672 4.7699
R14945 GND.n4140 GND.n4139 4.74817
R14946 GND.n4094 GND.n2273 4.74817
R14947 GND.n4124 GND.n4096 4.74817
R14948 GND.n4122 GND.n4121 4.74817
R14949 GND.n4099 GND.n4098 4.74817
R14950 GND.n4141 GND.n4140 4.74817
R14951 GND.n4138 GND.n2273 4.74817
R14952 GND.n4096 GND.n4095 4.74817
R14953 GND.n4123 GND.n4122 4.74817
R14954 GND.n4098 GND.n4097 4.74817
R14955 GND.n3001 GND.n3000 4.74817
R14956 GND.n3094 GND.n2702 4.74817
R14957 GND.n3092 GND.n3091 4.74817
R14958 GND.n3025 GND.n3024 4.74817
R14959 GND.n3076 GND.n3075 4.74817
R14960 GND.n4086 GND.n2259 4.74817
R14961 GND.n4130 GND.n2258 4.74817
R14962 GND.n4107 GND.n2257 4.74817
R14963 GND.n4111 GND.n2256 4.74817
R14964 GND.n4158 GND.n2255 4.74817
R14965 GND.n2262 GND.n2259 4.74817
R14966 GND.n4087 GND.n2258 4.74817
R14967 GND.n4129 GND.n2257 4.74817
R14968 GND.n4108 GND.n2256 4.74817
R14969 GND.n4110 GND.n2255 4.74817
R14970 GND.n3105 GND.n3104 4.74817
R14971 GND.n2712 GND.n2688 4.74817
R14972 GND.n3085 GND.n2687 4.74817
R14973 GND.n2718 GND.n2686 4.74817
R14974 GND.n2685 GND.n2682 4.74817
R14975 GND.n3105 GND.n2689 4.74817
R14976 GND.n3103 GND.n2688 4.74817
R14977 GND.n2713 GND.n2687 4.74817
R14978 GND.n3086 GND.n2686 4.74817
R14979 GND.n2717 GND.n2685 4.74817
R14980 GND.n3000 GND.n2999 4.74817
R14981 GND.n2998 GND.n2702 4.74817
R14982 GND.n3093 GND.n3092 4.74817
R14983 GND.n3024 GND.n2703 4.74817
R14984 GND.n3077 GND.n3076 4.74817
R14985 GND.n207 GND.n206 4.7074
R14986 GND.n603 GND.n602 4.7074
R14987 GND.n2531 GND.n1798 4.6279
R14988 GND.n2501 GND.n1865 4.6279
R14989 GND.n4312 GND.n2005 4.6132
R14990 GND.n4660 GND.n1552 4.6132
R14991 GND.n1961 GND.n1948 4.46111
R14992 GND.n82 GND.n78 4.38594
R14993 GND.n119 GND.n115 4.38594
R14994 GND.n151 GND.n147 4.38594
R14995 GND.n188 GND.n184 4.38594
R14996 GND.n13 GND.n9 4.38594
R14997 GND.n50 GND.n46 4.38594
R14998 GND.n515 GND.n511 4.38594
R14999 GND.n478 GND.n474 4.38594
R15000 GND.n584 GND.n580 4.38594
R15001 GND.n547 GND.n543 4.38594
R15002 GND.n654 GND.n650 4.38594
R15003 GND.n617 GND.n613 4.38594
R15004 GND.n318 GND.n314 4.38594
R15005 GND.n286 GND.n282 4.38594
R15006 GND.n254 GND.n250 4.38594
R15007 GND.n223 GND.n219 4.38594
R15008 GND.n445 GND.n441 4.38594
R15009 GND.n413 GND.n409 4.38594
R15010 GND.n381 GND.n377 4.38594
R15011 GND.n350 GND.n346 4.38594
R15012 GND.n93 GND.n71 4.26717
R15013 GND.n130 GND.n108 4.26717
R15014 GND.n162 GND.n140 4.26717
R15015 GND.n199 GND.n177 4.26717
R15016 GND.n24 GND.n2 4.26717
R15017 GND.n61 GND.n39 4.26717
R15018 GND.n526 GND.n504 4.26717
R15019 GND.n489 GND.n467 4.26717
R15020 GND.n595 GND.n573 4.26717
R15021 GND.n558 GND.n536 4.26717
R15022 GND.n665 GND.n643 4.26717
R15023 GND.n628 GND.n606 4.26717
R15024 GND.n329 GND.n307 4.26717
R15025 GND.n297 GND.n275 4.26717
R15026 GND.n265 GND.n243 4.26717
R15027 GND.n234 GND.n212 4.26717
R15028 GND.n456 GND.n434 4.26717
R15029 GND.n424 GND.n402 4.26717
R15030 GND.n392 GND.n370 4.26717
R15031 GND.n361 GND.n339 4.26717
R15032 GND.n464 GND.n336 4.14478
R15033 GND.n3732 GND.n3725 4.05904
R15034 GND.n3426 GND.n3314 4.05904
R15035 GND.n3408 GND.n3407 4.05904
R15036 GND.n4323 GND.n4322 4.05904
R15037 GND.n3515 GND.n2563 3.96685
R15038 GND.n4393 GND.n4392 3.96685
R15039 GND.n3718 GND.t32 3.96685
R15040 GND.n3205 GND.t43 3.63632
R15041 GND.n3489 GND.t20 3.63632
R15042 GND.n3717 GND.t14 3.63632
R15043 GND.t25 GND.n2362 3.63632
R15044 GND.n464 GND.n463 3.60163
R15045 GND.n92 GND.n73 3.49141
R15046 GND.n129 GND.n110 3.49141
R15047 GND.n161 GND.n142 3.49141
R15048 GND.n198 GND.n179 3.49141
R15049 GND.n23 GND.n4 3.49141
R15050 GND.n60 GND.n41 3.49141
R15051 GND.n525 GND.n506 3.49141
R15052 GND.n488 GND.n469 3.49141
R15053 GND.n594 GND.n575 3.49141
R15054 GND.n557 GND.n538 3.49141
R15055 GND.n664 GND.n645 3.49141
R15056 GND.n627 GND.n608 3.49141
R15057 GND.n328 GND.n309 3.49141
R15058 GND.n296 GND.n277 3.49141
R15059 GND.n264 GND.n245 3.49141
R15060 GND.n233 GND.n214 3.49141
R15061 GND.n455 GND.n436 3.49141
R15062 GND.n423 GND.n404 3.49141
R15063 GND.n391 GND.n372 3.49141
R15064 GND.n360 GND.n341 3.49141
R15065 GND.n4504 GND.t94 3.30579
R15066 GND.n4483 GND.n1775 3.30579
R15067 GND.n3537 GND.t19 3.30579
R15068 GND.n2495 GND.t7 3.30579
R15069 GND.n4400 GND.n1906 3.30579
R15070 GND.n100 GND.t153 3.3005
R15071 GND.n100 GND.t142 3.3005
R15072 GND.n102 GND.t176 3.3005
R15073 GND.n102 GND.t139 3.3005
R15074 GND.n104 GND.t128 3.3005
R15075 GND.n104 GND.t155 3.3005
R15076 GND.n169 GND.t149 3.3005
R15077 GND.n169 GND.t130 3.3005
R15078 GND.n171 GND.t163 3.3005
R15079 GND.n171 GND.t132 3.3005
R15080 GND.n173 GND.t179 3.3005
R15081 GND.n173 GND.t161 3.3005
R15082 GND.n31 GND.t165 3.3005
R15083 GND.n31 GND.t135 3.3005
R15084 GND.n33 GND.t117 3.3005
R15085 GND.n33 GND.t164 3.3005
R15086 GND.n35 GND.t138 3.3005
R15087 GND.n35 GND.t160 3.3005
R15088 GND.n500 GND.t152 3.3005
R15089 GND.n500 GND.t173 3.3005
R15090 GND.n498 GND.t121 3.3005
R15091 GND.n498 GND.t156 3.3005
R15092 GND.n496 GND.t123 3.3005
R15093 GND.n496 GND.t119 3.3005
R15094 GND.n569 GND.t144 3.3005
R15095 GND.n569 GND.t162 3.3005
R15096 GND.n567 GND.t174 3.3005
R15097 GND.n567 GND.t146 3.3005
R15098 GND.n565 GND.t175 3.3005
R15099 GND.n565 GND.t171 3.3005
R15100 GND.n639 GND.t151 3.3005
R15101 GND.n639 GND.t134 3.3005
R15102 GND.n637 GND.t157 3.3005
R15103 GND.n637 GND.t177 3.3005
R15104 GND.n635 GND.t124 3.3005
R15105 GND.n635 GND.t166 3.3005
R15106 GND.n89 GND.n88 2.71565
R15107 GND.n126 GND.n125 2.71565
R15108 GND.n158 GND.n157 2.71565
R15109 GND.n195 GND.n194 2.71565
R15110 GND.n20 GND.n19 2.71565
R15111 GND.n57 GND.n56 2.71565
R15112 GND.n522 GND.n521 2.71565
R15113 GND.n485 GND.n484 2.71565
R15114 GND.n591 GND.n590 2.71565
R15115 GND.n554 GND.n553 2.71565
R15116 GND.n661 GND.n660 2.71565
R15117 GND.n624 GND.n623 2.71565
R15118 GND.n325 GND.n324 2.71565
R15119 GND.n293 GND.n292 2.71565
R15120 GND.n261 GND.n260 2.71565
R15121 GND.n230 GND.n229 2.71565
R15122 GND.n452 GND.n451 2.71565
R15123 GND.n420 GND.n419 2.71565
R15124 GND.n388 GND.n387 2.71565
R15125 GND.n357 GND.n356 2.71565
R15126 GND.n3516 GND.t114 2.64473
R15127 GND.n3504 GND.n3503 2.64473
R15128 GND.n3504 GND.t29 2.64473
R15129 GND.n4469 GND.t8 2.64473
R15130 GND.n3583 GND.t5 2.64473
R15131 GND.n3582 GND.n3581 2.64473
R15132 GND.n3557 GND.t11 2.64473
R15133 GND.n4434 GND.t4 2.64473
R15134 GND.n3633 GND.n1854 2.64473
R15135 GND.n4427 GND.t16 2.64473
R15136 GND.n3662 GND.t6 2.64473
R15137 GND.n4399 GND.n1908 2.64473
R15138 GND.n208 GND.n207 2.4477
R15139 GND.n673 GND.n603 2.4477
R15140 GND.n3536 GND.t12 2.3142
R15141 GND.t12 GND.n1786 2.3142
R15142 GND.n4407 GND.t2 2.3142
R15143 GND.t2 GND.n4406 2.3142
R15144 GND.n4140 GND.n2244 2.27742
R15145 GND.n2273 GND.n2244 2.27742
R15146 GND.n4096 GND.n2244 2.27742
R15147 GND.n4122 GND.n2244 2.27742
R15148 GND.n4098 GND.n2244 2.27742
R15149 GND.n4148 GND.n2259 2.27742
R15150 GND.n4148 GND.n2258 2.27742
R15151 GND.n4148 GND.n2257 2.27742
R15152 GND.n4148 GND.n2256 2.27742
R15153 GND.n4148 GND.n2255 2.27742
R15154 GND.n3106 GND.n3105 2.27742
R15155 GND.n3106 GND.n2688 2.27742
R15156 GND.n3106 GND.n2687 2.27742
R15157 GND.n3106 GND.n2686 2.27742
R15158 GND.n3106 GND.n2685 2.27742
R15159 GND.n3000 GND.n2684 2.27742
R15160 GND.n2702 GND.n2684 2.27742
R15161 GND.n3092 GND.n2684 2.27742
R15162 GND.n3024 GND.n2684 2.27742
R15163 GND.n3076 GND.n2684 2.27742
R15164 GND.n3296 GND.t82 1.98367
R15165 GND.t94 GND.n4503 1.98367
R15166 GND.t35 GND.n1758 1.98367
R15167 GND.n3516 GND.n1766 1.98367
R15168 GND.n3556 GND.n3555 1.98367
R15169 GND.n4433 GND.n1845 1.98367
R15170 GND.t107 GND.n3706 1.98367
R15171 GND.n3707 GND.n1917 1.98367
R15172 GND.n3711 GND.t59 1.98367
R15173 GND.n85 GND.n75 1.93989
R15174 GND.n122 GND.n112 1.93989
R15175 GND.n154 GND.n144 1.93989
R15176 GND.n191 GND.n181 1.93989
R15177 GND.n16 GND.n6 1.93989
R15178 GND.n53 GND.n43 1.93989
R15179 GND.n518 GND.n508 1.93989
R15180 GND.n481 GND.n471 1.93989
R15181 GND.n587 GND.n577 1.93989
R15182 GND.n550 GND.n540 1.93989
R15183 GND.n657 GND.n647 1.93989
R15184 GND.n620 GND.n610 1.93989
R15185 GND.n321 GND.n311 1.93989
R15186 GND.n289 GND.n279 1.93989
R15187 GND.n257 GND.n247 1.93989
R15188 GND.n226 GND.n216 1.93989
R15189 GND.n448 GND.n438 1.93989
R15190 GND.n416 GND.n406 1.93989
R15191 GND.n384 GND.n374 1.93989
R15192 GND.n353 GND.n343 1.93989
R15193 GND.n4511 GND.n1734 1.65314
R15194 GND.t20 GND.n3488 1.65314
R15195 GND.t14 GND.n1928 1.65314
R15196 GND.n4371 GND.n1969 1.65314
R15197 GND.n2944 GND.n2790 1.32262
R15198 GND.n2941 GND.n2762 1.32262
R15199 GND.n2954 GND.n2763 1.32262
R15200 GND.n2766 GND.n2755 1.32262
R15201 GND.n2977 GND.n2749 1.32262
R15202 GND.n2981 GND.n2752 1.32262
R15203 GND.n2991 GND.n2738 1.32262
R15204 GND.n2965 GND.n2962 1.32262
R15205 GND.n3003 GND.n2730 1.32262
R15206 GND.n3004 GND.n2692 1.32262
R15207 GND.n3101 GND.n2694 1.32262
R15208 GND.n3097 GND.n3096 1.32262
R15209 GND.n2705 GND.n2699 1.32262
R15210 GND.n3089 GND.n2706 1.32262
R15211 GND.n3088 GND.n2708 1.32262
R15212 GND.n3083 GND.n2720 1.32262
R15213 GND.n3080 GND.n3079 1.32262
R15214 GND.n3021 GND.n2676 1.32262
R15215 GND.n3111 GND.n2677 1.32262
R15216 GND.n3071 GND.n3070 1.32262
R15217 GND.n3120 GND.n2665 1.32262
R15218 GND.n3126 GND.n2667 1.32262
R15219 GND.n3123 GND.n2656 1.32262
R15220 GND.n3136 GND.n2657 1.32262
R15221 GND.n3062 GND.n3061 1.32262
R15222 GND.n3145 GND.n2646 1.32262
R15223 GND.n3151 GND.n2648 1.32262
R15224 GND.n3147 GND.n2636 1.32262
R15225 GND.n3161 GND.n2638 1.32262
R15226 GND.n3041 GND.n3040 1.32262
R15227 GND.n3173 GND.n2625 1.32262
R15228 GND.n3177 GND.n2627 1.32262
R15229 GND.n3186 GND.n2619 1.32262
R15230 GND.n3185 GND.n2604 1.32262
R15231 GND.n3214 GND.n2599 1.32262
R15232 GND.n3217 GND.n2601 1.32262
R15233 GND.n3206 GND.n3205 1.32262
R15234 GND.n3225 GND.n2592 1.32262
R15235 GND.n3230 GND.n1525 1.32262
R15236 GND.n4685 GND.n1527 1.32262
R15237 GND.n3540 GND.n3537 1.32262
R15238 GND.n3572 GND.n3568 1.32262
R15239 GND.n3604 GND.t11 1.32262
R15240 GND.n3640 GND.t4 1.32262
R15241 GND.n4420 GND.n4419 1.32262
R15242 GND.n2496 GND.n2495 1.32262
R15243 GND.t79 GND.n1944 1.32262
R15244 GND.n3919 GND.n3918 1.32262
R15245 GND.n3982 GND.n2413 1.32262
R15246 GND.n3978 GND.n3977 1.32262
R15247 GND.n3992 GND.n2362 1.32262
R15248 GND.n2367 GND.n2364 1.32262
R15249 GND.n4001 GND.n2355 1.32262
R15250 GND.n4007 GND.n2350 1.32262
R15251 GND.n4004 GND.n2352 1.32262
R15252 GND.n4017 GND.n2340 1.32262
R15253 GND.n2344 GND.n2341 1.32262
R15254 GND.n4026 GND.n2333 1.32262
R15255 GND.n4031 GND.n2327 1.32262
R15256 GND.n4028 GND.n2330 1.32262
R15257 GND.n4041 GND.n2316 1.32262
R15258 GND.n2321 GND.n2317 1.32262
R15259 GND.n4050 GND.n2308 1.32262
R15260 GND.n4056 GND.n2304 1.32262
R15261 GND.n4053 GND.n2306 1.32262
R15262 GND.n4067 GND.n2290 1.32262
R15263 GND.n2298 GND.n2291 1.32262
R15264 GND.n2295 GND.n2265 1.32262
R15265 GND.n4144 GND.n4143 1.32262
R15266 GND.n4075 GND.n2267 1.32262
R15267 GND.n4136 GND.n2275 1.32262
R15268 GND.n4133 GND.n2281 1.32262
R15269 GND.n4132 GND.n4084 1.32262
R15270 GND.n4127 GND.n4126 1.32262
R15271 GND.n4104 GND.n4090 1.32262
R15272 GND.n4119 GND.n4102 1.32262
R15273 GND.n4116 GND.n4113 1.32262
R15274 GND.n4115 GND.n2252 1.32262
R15275 GND.n4162 GND.n4160 1.32262
R15276 GND.n4165 GND.n2247 1.32262
R15277 GND.n4175 GND.n2239 1.32262
R15278 GND.n2240 GND.n881 1.32262
R15279 GND.n5536 GND.n5535 1.32262
R15280 GND.n5544 GND.n868 1.32262
R15281 GND.n5529 GND.n5528 1.32262
R15282 GND.n5552 GND.n860 1.32262
R15283 GND.n861 GND.n846 1.32262
R15284 GND.n84 GND.n77 1.16414
R15285 GND.n121 GND.n114 1.16414
R15286 GND.n153 GND.n146 1.16414
R15287 GND.n190 GND.n183 1.16414
R15288 GND.n15 GND.n8 1.16414
R15289 GND.n52 GND.n45 1.16414
R15290 GND.n517 GND.n510 1.16414
R15291 GND.n480 GND.n473 1.16414
R15292 GND.n586 GND.n579 1.16414
R15293 GND.n549 GND.n542 1.16414
R15294 GND.n656 GND.n649 1.16414
R15295 GND.n619 GND.n612 1.16414
R15296 GND.n2099 GND.n2095 1.16414
R15297 GND.n3256 GND.n3255 1.16414
R15298 GND.n320 GND.n313 1.16414
R15299 GND.n288 GND.n281 1.16414
R15300 GND.n256 GND.n249 1.16414
R15301 GND.n225 GND.n218 1.16414
R15302 GND.n447 GND.n440 1.16414
R15303 GND.n415 GND.n408 1.16414
R15304 GND.n383 GND.n376 1.16414
R15305 GND.n352 GND.n345 1.16414
R15306 GND.n137 GND.n105 1.00481
R15307 GND.n105 GND.n103 1.00481
R15308 GND.n103 GND.n101 1.00481
R15309 GND.n206 GND.n174 1.00481
R15310 GND.n174 GND.n172 1.00481
R15311 GND.n172 GND.n170 1.00481
R15312 GND.n68 GND.n36 1.00481
R15313 GND.n36 GND.n34 1.00481
R15314 GND.n34 GND.n32 1.00481
R15315 GND.n499 GND.n497 1.00481
R15316 GND.n501 GND.n499 1.00481
R15317 GND.n533 GND.n501 1.00481
R15318 GND.n568 GND.n566 1.00481
R15319 GND.n570 GND.n568 1.00481
R15320 GND.n602 GND.n570 1.00481
R15321 GND.n638 GND.n636 1.00481
R15322 GND.n640 GND.n638 1.00481
R15323 GND.n672 GND.n640 1.00481
R15324 GND GND.n209 0.99596
R15325 GND.n2961 GND.t154 0.992087
R15326 GND.n2250 GND.t143 0.992087
R15327 GND.n4660 GND.n4659 0.970197
R15328 GND.n4312 GND.n4311 0.970197
R15329 GND.n304 GND.n272 0.962709
R15330 GND.n336 GND.n304 0.962709
R15331 GND.n431 GND.n399 0.962709
R15332 GND.n463 GND.n431 0.962709
R15333 GND.n3479 GND.n1746 0.661558
R15334 GND.n4497 GND.n1755 0.661558
R15335 GND.n4461 GND.t5 0.661558
R15336 GND.n4447 GND.n1827 0.661558
R15337 GND.n3624 GND.n1836 0.661558
R15338 GND.t16 GND.n4426 0.661558
R15339 GND.t59 GND.t50 0.661558
R15340 GND.n4386 GND.n4385 0.661558
R15341 GND.n4379 GND.n4378 0.661558
R15342 GND.n5759 GND.n5758 0.57484
R15343 GND.n4148 GND.n2244 0.570125
R15344 GND.n3106 GND.n2684 0.570125
R15345 GND.n1225 GND.n1220 0.486781
R15346 GND.n5363 GND.n5362 0.486781
R15347 GND.n5524 GND.n5523 0.486781
R15348 GND.n2776 GND.n2775 0.486781
R15349 GND.n4242 GND.n4241 0.48678
R15350 GND.n3267 GND.n3266 0.48678
R15351 GND.n5717 GND.n5716 0.483732
R15352 GND.n2874 GND.n2871 0.483732
R15353 GND.n2372 GND.n2370 0.471537
R15354 GND.n2905 GND.n1379 0.471537
R15355 GND.n5710 GND.n745 0.471537
R15356 GND.n4682 GND.n4681 0.471537
R15357 GND.n81 GND.n80 0.388379
R15358 GND.n118 GND.n117 0.388379
R15359 GND.n150 GND.n149 0.388379
R15360 GND.n187 GND.n186 0.388379
R15361 GND.n12 GND.n11 0.388379
R15362 GND.n49 GND.n48 0.388379
R15363 GND.n514 GND.n513 0.388379
R15364 GND.n477 GND.n476 0.388379
R15365 GND.n583 GND.n582 0.388379
R15366 GND.n546 GND.n545 0.388379
R15367 GND.n653 GND.n652 0.388379
R15368 GND.n616 GND.n615 0.388379
R15369 GND.n5688 GND.n5687 0.388379
R15370 GND.n4806 GND.n4805 0.388379
R15371 GND.n317 GND.n316 0.388379
R15372 GND.n285 GND.n284 0.388379
R15373 GND.n253 GND.n252 0.388379
R15374 GND.n222 GND.n221 0.388379
R15375 GND.n444 GND.n443 0.388379
R15376 GND.n412 GND.n411 0.388379
R15377 GND.n380 GND.n379 0.388379
R15378 GND.n349 GND.n348 0.388379
R15379 GND.n5759 GND.n464 0.341877
R15380 GND.n2990 GND.t154 0.331029
R15381 GND.n3120 GND.t148 0.331029
R15382 GND.n4539 GND.t103 0.331029
R15383 GND.n2437 GND.t110 0.331029
R15384 GND.n2298 GND.t118 0.331029
R15385 GND.t143 GND.n2249 0.331029
R15386 GND.n5649 GND.n798 0.293183
R15387 GND.n2841 GND.n1418 0.293183
R15388 GND.n4233 GND.n2113 0.280988
R15389 GND.n4769 GND.n1418 0.280988
R15390 GND.n5659 GND.n798 0.280988
R15391 GND.n4632 GND.n4630 0.280988
R15392 GND.n3915 GND.n2090 0.253549
R15393 GND.n3235 GND.n3234 0.253549
R15394 GND.n4629 GND.n1579 0.245927
R15395 GND.n4235 GND.n4234 0.245927
R15396 GND.n2384 GND.n2005 0.229039
R15397 GND.n2008 GND.n2005 0.229039
R15398 GND.n1552 GND.n1547 0.229039
R15399 GND.n4658 GND.n1552 0.229039
R15400 GND GND.n5759 0.213018
R15401 GND.n4234 GND.n4233 0.207029
R15402 GND.n4630 GND.n4629 0.207029
R15403 GND.n98 GND.n70 0.155672
R15404 GND.n91 GND.n70 0.155672
R15405 GND.n91 GND.n90 0.155672
R15406 GND.n90 GND.n74 0.155672
R15407 GND.n83 GND.n74 0.155672
R15408 GND.n83 GND.n82 0.155672
R15409 GND.n135 GND.n107 0.155672
R15410 GND.n128 GND.n107 0.155672
R15411 GND.n128 GND.n127 0.155672
R15412 GND.n127 GND.n111 0.155672
R15413 GND.n120 GND.n111 0.155672
R15414 GND.n120 GND.n119 0.155672
R15415 GND.n167 GND.n139 0.155672
R15416 GND.n160 GND.n139 0.155672
R15417 GND.n160 GND.n159 0.155672
R15418 GND.n159 GND.n143 0.155672
R15419 GND.n152 GND.n143 0.155672
R15420 GND.n152 GND.n151 0.155672
R15421 GND.n204 GND.n176 0.155672
R15422 GND.n197 GND.n176 0.155672
R15423 GND.n197 GND.n196 0.155672
R15424 GND.n196 GND.n180 0.155672
R15425 GND.n189 GND.n180 0.155672
R15426 GND.n189 GND.n188 0.155672
R15427 GND.n29 GND.n1 0.155672
R15428 GND.n22 GND.n1 0.155672
R15429 GND.n22 GND.n21 0.155672
R15430 GND.n21 GND.n5 0.155672
R15431 GND.n14 GND.n5 0.155672
R15432 GND.n14 GND.n13 0.155672
R15433 GND.n66 GND.n38 0.155672
R15434 GND.n59 GND.n38 0.155672
R15435 GND.n59 GND.n58 0.155672
R15436 GND.n58 GND.n42 0.155672
R15437 GND.n51 GND.n42 0.155672
R15438 GND.n51 GND.n50 0.155672
R15439 GND.n531 GND.n503 0.155672
R15440 GND.n524 GND.n503 0.155672
R15441 GND.n524 GND.n523 0.155672
R15442 GND.n523 GND.n507 0.155672
R15443 GND.n516 GND.n507 0.155672
R15444 GND.n516 GND.n515 0.155672
R15445 GND.n494 GND.n466 0.155672
R15446 GND.n487 GND.n466 0.155672
R15447 GND.n487 GND.n486 0.155672
R15448 GND.n486 GND.n470 0.155672
R15449 GND.n479 GND.n470 0.155672
R15450 GND.n479 GND.n478 0.155672
R15451 GND.n600 GND.n572 0.155672
R15452 GND.n593 GND.n572 0.155672
R15453 GND.n593 GND.n592 0.155672
R15454 GND.n592 GND.n576 0.155672
R15455 GND.n585 GND.n576 0.155672
R15456 GND.n585 GND.n584 0.155672
R15457 GND.n563 GND.n535 0.155672
R15458 GND.n556 GND.n535 0.155672
R15459 GND.n556 GND.n555 0.155672
R15460 GND.n555 GND.n539 0.155672
R15461 GND.n548 GND.n539 0.155672
R15462 GND.n548 GND.n547 0.155672
R15463 GND.n670 GND.n642 0.155672
R15464 GND.n663 GND.n642 0.155672
R15465 GND.n663 GND.n662 0.155672
R15466 GND.n662 GND.n646 0.155672
R15467 GND.n655 GND.n646 0.155672
R15468 GND.n655 GND.n654 0.155672
R15469 GND.n633 GND.n605 0.155672
R15470 GND.n626 GND.n605 0.155672
R15471 GND.n626 GND.n625 0.155672
R15472 GND.n625 GND.n609 0.155672
R15473 GND.n618 GND.n609 0.155672
R15474 GND.n618 GND.n617 0.155672
R15475 GND.n334 GND.n306 0.155672
R15476 GND.n327 GND.n306 0.155672
R15477 GND.n327 GND.n326 0.155672
R15478 GND.n326 GND.n310 0.155672
R15479 GND.n319 GND.n310 0.155672
R15480 GND.n319 GND.n318 0.155672
R15481 GND.n302 GND.n274 0.155672
R15482 GND.n295 GND.n274 0.155672
R15483 GND.n295 GND.n294 0.155672
R15484 GND.n294 GND.n278 0.155672
R15485 GND.n287 GND.n278 0.155672
R15486 GND.n287 GND.n286 0.155672
R15487 GND.n270 GND.n242 0.155672
R15488 GND.n263 GND.n242 0.155672
R15489 GND.n263 GND.n262 0.155672
R15490 GND.n262 GND.n246 0.155672
R15491 GND.n255 GND.n246 0.155672
R15492 GND.n255 GND.n254 0.155672
R15493 GND.n239 GND.n211 0.155672
R15494 GND.n232 GND.n211 0.155672
R15495 GND.n232 GND.n231 0.155672
R15496 GND.n231 GND.n215 0.155672
R15497 GND.n224 GND.n215 0.155672
R15498 GND.n224 GND.n223 0.155672
R15499 GND.n461 GND.n433 0.155672
R15500 GND.n454 GND.n433 0.155672
R15501 GND.n454 GND.n453 0.155672
R15502 GND.n453 GND.n437 0.155672
R15503 GND.n446 GND.n437 0.155672
R15504 GND.n446 GND.n445 0.155672
R15505 GND.n429 GND.n401 0.155672
R15506 GND.n422 GND.n401 0.155672
R15507 GND.n422 GND.n421 0.155672
R15508 GND.n421 GND.n405 0.155672
R15509 GND.n414 GND.n405 0.155672
R15510 GND.n414 GND.n413 0.155672
R15511 GND.n397 GND.n369 0.155672
R15512 GND.n390 GND.n369 0.155672
R15513 GND.n390 GND.n389 0.155672
R15514 GND.n389 GND.n373 0.155672
R15515 GND.n382 GND.n373 0.155672
R15516 GND.n382 GND.n381 0.155672
R15517 GND.n366 GND.n338 0.155672
R15518 GND.n359 GND.n338 0.155672
R15519 GND.n359 GND.n358 0.155672
R15520 GND.n358 GND.n342 0.155672
R15521 GND.n351 GND.n342 0.155672
R15522 GND.n351 GND.n350 0.155672
R15523 GND.n1687 GND.n1579 0.152939
R15524 GND.n1688 GND.n1687 0.152939
R15525 GND.n1689 GND.n1688 0.152939
R15526 GND.n1690 GND.n1689 0.152939
R15527 GND.n1691 GND.n1690 0.152939
R15528 GND.n1714 GND.n1691 0.152939
R15529 GND.n1715 GND.n1714 0.152939
R15530 GND.n1716 GND.n1715 0.152939
R15531 GND.n1717 GND.n1716 0.152939
R15532 GND.n1718 GND.n1717 0.152939
R15533 GND.n1739 GND.n1718 0.152939
R15534 GND.n1740 GND.n1739 0.152939
R15535 GND.n1741 GND.n1740 0.152939
R15536 GND.n1742 GND.n1741 0.152939
R15537 GND.n1743 GND.n1742 0.152939
R15538 GND.n1760 GND.n1743 0.152939
R15539 GND.n1761 GND.n1760 0.152939
R15540 GND.n1762 GND.n1761 0.152939
R15541 GND.n1763 GND.n1762 0.152939
R15542 GND.n1780 GND.n1763 0.152939
R15543 GND.n1781 GND.n1780 0.152939
R15544 GND.n1782 GND.n1781 0.152939
R15545 GND.n1783 GND.n1782 0.152939
R15546 GND.n1800 GND.n1783 0.152939
R15547 GND.n1801 GND.n1800 0.152939
R15548 GND.n1802 GND.n1801 0.152939
R15549 GND.n1803 GND.n1802 0.152939
R15550 GND.n1818 GND.n1803 0.152939
R15551 GND.n1819 GND.n1818 0.152939
R15552 GND.n1820 GND.n1819 0.152939
R15553 GND.n1821 GND.n1820 0.152939
R15554 GND.n1838 GND.n1821 0.152939
R15555 GND.n1839 GND.n1838 0.152939
R15556 GND.n1840 GND.n1839 0.152939
R15557 GND.n1841 GND.n1840 0.152939
R15558 GND.n1869 GND.n1841 0.152939
R15559 GND.n1872 GND.n1869 0.152939
R15560 GND.n1873 GND.n1872 0.152939
R15561 GND.n1874 GND.n1873 0.152939
R15562 GND.n1875 GND.n1874 0.152939
R15563 GND.n1876 GND.n1875 0.152939
R15564 GND.n2490 GND.n1876 0.152939
R15565 GND.n2492 GND.n2490 0.152939
R15566 GND.n2492 GND.n2491 0.152939
R15567 GND.n2491 GND.n1912 0.152939
R15568 GND.n1913 GND.n1912 0.152939
R15569 GND.n1914 GND.n1913 0.152939
R15570 GND.n3792 GND.n1914 0.152939
R15571 GND.n3793 GND.n3792 0.152939
R15572 GND.n3793 GND.n3790 0.152939
R15573 GND.n3799 GND.n3790 0.152939
R15574 GND.n3800 GND.n3799 0.152939
R15575 GND.n3801 GND.n3800 0.152939
R15576 GND.n3802 GND.n3801 0.152939
R15577 GND.n3802 GND.n2456 0.152939
R15578 GND.n3831 GND.n2456 0.152939
R15579 GND.n3832 GND.n3831 0.152939
R15580 GND.n3833 GND.n3832 0.152939
R15581 GND.n3834 GND.n3833 0.152939
R15582 GND.n3834 GND.n2432 0.152939
R15583 GND.n3865 GND.n2432 0.152939
R15584 GND.n3866 GND.n3865 0.152939
R15585 GND.n3867 GND.n3866 0.152939
R15586 GND.n3867 GND.n2112 0.152939
R15587 GND.n4235 GND.n2112 0.152939
R15588 GND.n4970 GND.n1220 0.152939
R15589 GND.n4971 GND.n4970 0.152939
R15590 GND.n4972 GND.n4971 0.152939
R15591 GND.n4972 GND.n1214 0.152939
R15592 GND.n4980 GND.n1214 0.152939
R15593 GND.n4981 GND.n4980 0.152939
R15594 GND.n4982 GND.n4981 0.152939
R15595 GND.n4982 GND.n1208 0.152939
R15596 GND.n4990 GND.n1208 0.152939
R15597 GND.n4991 GND.n4990 0.152939
R15598 GND.n4992 GND.n4991 0.152939
R15599 GND.n4992 GND.n1202 0.152939
R15600 GND.n5000 GND.n1202 0.152939
R15601 GND.n5001 GND.n5000 0.152939
R15602 GND.n5002 GND.n5001 0.152939
R15603 GND.n5002 GND.n1196 0.152939
R15604 GND.n5010 GND.n1196 0.152939
R15605 GND.n5011 GND.n5010 0.152939
R15606 GND.n5012 GND.n5011 0.152939
R15607 GND.n5012 GND.n1190 0.152939
R15608 GND.n5020 GND.n1190 0.152939
R15609 GND.n5021 GND.n5020 0.152939
R15610 GND.n5022 GND.n5021 0.152939
R15611 GND.n5022 GND.n1184 0.152939
R15612 GND.n5030 GND.n1184 0.152939
R15613 GND.n5031 GND.n5030 0.152939
R15614 GND.n5032 GND.n5031 0.152939
R15615 GND.n5032 GND.n1178 0.152939
R15616 GND.n5040 GND.n1178 0.152939
R15617 GND.n5041 GND.n5040 0.152939
R15618 GND.n5042 GND.n5041 0.152939
R15619 GND.n5042 GND.n1172 0.152939
R15620 GND.n5050 GND.n1172 0.152939
R15621 GND.n5051 GND.n5050 0.152939
R15622 GND.n5052 GND.n5051 0.152939
R15623 GND.n5052 GND.n1166 0.152939
R15624 GND.n5060 GND.n1166 0.152939
R15625 GND.n5061 GND.n5060 0.152939
R15626 GND.n5062 GND.n5061 0.152939
R15627 GND.n5062 GND.n1160 0.152939
R15628 GND.n5070 GND.n1160 0.152939
R15629 GND.n5071 GND.n5070 0.152939
R15630 GND.n5072 GND.n5071 0.152939
R15631 GND.n5072 GND.n1154 0.152939
R15632 GND.n5080 GND.n1154 0.152939
R15633 GND.n5081 GND.n5080 0.152939
R15634 GND.n5082 GND.n5081 0.152939
R15635 GND.n5082 GND.n1148 0.152939
R15636 GND.n5090 GND.n1148 0.152939
R15637 GND.n5091 GND.n5090 0.152939
R15638 GND.n5092 GND.n5091 0.152939
R15639 GND.n5092 GND.n1142 0.152939
R15640 GND.n5100 GND.n1142 0.152939
R15641 GND.n5101 GND.n5100 0.152939
R15642 GND.n5102 GND.n5101 0.152939
R15643 GND.n5102 GND.n1136 0.152939
R15644 GND.n5110 GND.n1136 0.152939
R15645 GND.n5111 GND.n5110 0.152939
R15646 GND.n5112 GND.n5111 0.152939
R15647 GND.n5112 GND.n1130 0.152939
R15648 GND.n5120 GND.n1130 0.152939
R15649 GND.n5121 GND.n5120 0.152939
R15650 GND.n5122 GND.n5121 0.152939
R15651 GND.n5122 GND.n1124 0.152939
R15652 GND.n5130 GND.n1124 0.152939
R15653 GND.n5131 GND.n5130 0.152939
R15654 GND.n5132 GND.n5131 0.152939
R15655 GND.n5132 GND.n1118 0.152939
R15656 GND.n5140 GND.n1118 0.152939
R15657 GND.n5141 GND.n5140 0.152939
R15658 GND.n5142 GND.n5141 0.152939
R15659 GND.n5142 GND.n1112 0.152939
R15660 GND.n5150 GND.n1112 0.152939
R15661 GND.n5151 GND.n5150 0.152939
R15662 GND.n5152 GND.n5151 0.152939
R15663 GND.n5152 GND.n1106 0.152939
R15664 GND.n5160 GND.n1106 0.152939
R15665 GND.n5161 GND.n5160 0.152939
R15666 GND.n5162 GND.n5161 0.152939
R15667 GND.n5162 GND.n1100 0.152939
R15668 GND.n5170 GND.n1100 0.152939
R15669 GND.n5171 GND.n5170 0.152939
R15670 GND.n5172 GND.n5171 0.152939
R15671 GND.n5172 GND.n1094 0.152939
R15672 GND.n5180 GND.n1094 0.152939
R15673 GND.n5181 GND.n5180 0.152939
R15674 GND.n5182 GND.n5181 0.152939
R15675 GND.n5182 GND.n1088 0.152939
R15676 GND.n5190 GND.n1088 0.152939
R15677 GND.n5191 GND.n5190 0.152939
R15678 GND.n5192 GND.n5191 0.152939
R15679 GND.n5192 GND.n1082 0.152939
R15680 GND.n5200 GND.n1082 0.152939
R15681 GND.n5201 GND.n5200 0.152939
R15682 GND.n5202 GND.n5201 0.152939
R15683 GND.n5202 GND.n1076 0.152939
R15684 GND.n5210 GND.n1076 0.152939
R15685 GND.n5211 GND.n5210 0.152939
R15686 GND.n5212 GND.n5211 0.152939
R15687 GND.n5212 GND.n1070 0.152939
R15688 GND.n5220 GND.n1070 0.152939
R15689 GND.n5221 GND.n5220 0.152939
R15690 GND.n5222 GND.n5221 0.152939
R15691 GND.n5222 GND.n1064 0.152939
R15692 GND.n5230 GND.n1064 0.152939
R15693 GND.n5231 GND.n5230 0.152939
R15694 GND.n5232 GND.n5231 0.152939
R15695 GND.n5232 GND.n1058 0.152939
R15696 GND.n5240 GND.n1058 0.152939
R15697 GND.n5241 GND.n5240 0.152939
R15698 GND.n5242 GND.n5241 0.152939
R15699 GND.n5242 GND.n1052 0.152939
R15700 GND.n5250 GND.n1052 0.152939
R15701 GND.n5251 GND.n5250 0.152939
R15702 GND.n5252 GND.n5251 0.152939
R15703 GND.n5252 GND.n1046 0.152939
R15704 GND.n5260 GND.n1046 0.152939
R15705 GND.n5261 GND.n5260 0.152939
R15706 GND.n5262 GND.n5261 0.152939
R15707 GND.n5262 GND.n1040 0.152939
R15708 GND.n5270 GND.n1040 0.152939
R15709 GND.n5271 GND.n5270 0.152939
R15710 GND.n5272 GND.n5271 0.152939
R15711 GND.n5272 GND.n1034 0.152939
R15712 GND.n5280 GND.n1034 0.152939
R15713 GND.n5281 GND.n5280 0.152939
R15714 GND.n5282 GND.n5281 0.152939
R15715 GND.n5282 GND.n1028 0.152939
R15716 GND.n5290 GND.n1028 0.152939
R15717 GND.n5291 GND.n5290 0.152939
R15718 GND.n5292 GND.n5291 0.152939
R15719 GND.n5292 GND.n1022 0.152939
R15720 GND.n5300 GND.n1022 0.152939
R15721 GND.n5301 GND.n5300 0.152939
R15722 GND.n5302 GND.n5301 0.152939
R15723 GND.n5302 GND.n1016 0.152939
R15724 GND.n5310 GND.n1016 0.152939
R15725 GND.n5311 GND.n5310 0.152939
R15726 GND.n5312 GND.n5311 0.152939
R15727 GND.n5312 GND.n1010 0.152939
R15728 GND.n5320 GND.n1010 0.152939
R15729 GND.n5321 GND.n5320 0.152939
R15730 GND.n5322 GND.n5321 0.152939
R15731 GND.n5322 GND.n1004 0.152939
R15732 GND.n5330 GND.n1004 0.152939
R15733 GND.n5331 GND.n5330 0.152939
R15734 GND.n5332 GND.n5331 0.152939
R15735 GND.n5332 GND.n998 0.152939
R15736 GND.n5340 GND.n998 0.152939
R15737 GND.n5341 GND.n5340 0.152939
R15738 GND.n5342 GND.n5341 0.152939
R15739 GND.n5342 GND.n992 0.152939
R15740 GND.n5350 GND.n992 0.152939
R15741 GND.n5351 GND.n5350 0.152939
R15742 GND.n5353 GND.n5351 0.152939
R15743 GND.n5353 GND.n5352 0.152939
R15744 GND.n5352 GND.n986 0.152939
R15745 GND.n5362 GND.n986 0.152939
R15746 GND.n5363 GND.n981 0.152939
R15747 GND.n5371 GND.n981 0.152939
R15748 GND.n5372 GND.n5371 0.152939
R15749 GND.n5373 GND.n5372 0.152939
R15750 GND.n5373 GND.n975 0.152939
R15751 GND.n5381 GND.n975 0.152939
R15752 GND.n5382 GND.n5381 0.152939
R15753 GND.n5383 GND.n5382 0.152939
R15754 GND.n5383 GND.n969 0.152939
R15755 GND.n5391 GND.n969 0.152939
R15756 GND.n5392 GND.n5391 0.152939
R15757 GND.n5393 GND.n5392 0.152939
R15758 GND.n5393 GND.n963 0.152939
R15759 GND.n5401 GND.n963 0.152939
R15760 GND.n5402 GND.n5401 0.152939
R15761 GND.n5403 GND.n5402 0.152939
R15762 GND.n5403 GND.n957 0.152939
R15763 GND.n5411 GND.n957 0.152939
R15764 GND.n5412 GND.n5411 0.152939
R15765 GND.n5413 GND.n5412 0.152939
R15766 GND.n5413 GND.n951 0.152939
R15767 GND.n5421 GND.n951 0.152939
R15768 GND.n5422 GND.n5421 0.152939
R15769 GND.n5423 GND.n5422 0.152939
R15770 GND.n5423 GND.n945 0.152939
R15771 GND.n5431 GND.n945 0.152939
R15772 GND.n5432 GND.n5431 0.152939
R15773 GND.n5433 GND.n5432 0.152939
R15774 GND.n5433 GND.n939 0.152939
R15775 GND.n5441 GND.n939 0.152939
R15776 GND.n5442 GND.n5441 0.152939
R15777 GND.n5443 GND.n5442 0.152939
R15778 GND.n5443 GND.n933 0.152939
R15779 GND.n5451 GND.n933 0.152939
R15780 GND.n5452 GND.n5451 0.152939
R15781 GND.n5453 GND.n5452 0.152939
R15782 GND.n5453 GND.n927 0.152939
R15783 GND.n5461 GND.n927 0.152939
R15784 GND.n5462 GND.n5461 0.152939
R15785 GND.n5463 GND.n5462 0.152939
R15786 GND.n5463 GND.n921 0.152939
R15787 GND.n5471 GND.n921 0.152939
R15788 GND.n5472 GND.n5471 0.152939
R15789 GND.n5473 GND.n5472 0.152939
R15790 GND.n5473 GND.n915 0.152939
R15791 GND.n5481 GND.n915 0.152939
R15792 GND.n5482 GND.n5481 0.152939
R15793 GND.n5483 GND.n5482 0.152939
R15794 GND.n5483 GND.n909 0.152939
R15795 GND.n5491 GND.n909 0.152939
R15796 GND.n5492 GND.n5491 0.152939
R15797 GND.n5493 GND.n5492 0.152939
R15798 GND.n5493 GND.n903 0.152939
R15799 GND.n5501 GND.n903 0.152939
R15800 GND.n5502 GND.n5501 0.152939
R15801 GND.n5503 GND.n5502 0.152939
R15802 GND.n5503 GND.n897 0.152939
R15803 GND.n5511 GND.n897 0.152939
R15804 GND.n5512 GND.n5511 0.152939
R15805 GND.n5514 GND.n5512 0.152939
R15806 GND.n5514 GND.n5513 0.152939
R15807 GND.n5513 GND.n891 0.152939
R15808 GND.n5523 GND.n891 0.152939
R15809 GND.n4150 GND.n4149 0.152939
R15810 GND.n4152 GND.n4150 0.152939
R15811 GND.n4152 GND.n4151 0.152939
R15812 GND.n4151 GND.n885 0.152939
R15813 GND.n886 GND.n885 0.152939
R15814 GND.n887 GND.n886 0.152939
R15815 GND.n890 GND.n887 0.152939
R15816 GND.n5524 GND.n890 0.152939
R15817 GND.n4168 GND.n2244 0.152939
R15818 GND.n4169 GND.n4168 0.152939
R15819 GND.n4170 GND.n4169 0.152939
R15820 GND.n4171 GND.n4170 0.152939
R15821 GND.n4171 GND.n865 0.152939
R15822 GND.n5547 GND.n865 0.152939
R15823 GND.n5548 GND.n5547 0.152939
R15824 GND.n5549 GND.n5548 0.152939
R15825 GND.n5549 GND.n843 0.152939
R15826 GND.n5564 GND.n843 0.152939
R15827 GND.n5565 GND.n5564 0.152939
R15828 GND.n5566 GND.n5565 0.152939
R15829 GND.n5566 GND.n824 0.152939
R15830 GND.n5581 GND.n824 0.152939
R15831 GND.n5582 GND.n5581 0.152939
R15832 GND.n5583 GND.n5582 0.152939
R15833 GND.n5583 GND.n807 0.152939
R15834 GND.n5599 GND.n807 0.152939
R15835 GND.n5600 GND.n5599 0.152939
R15836 GND.n5601 GND.n5600 0.152939
R15837 GND.n5601 GND.n745 0.152939
R15838 GND.n2373 GND.n2372 0.152939
R15839 GND.n2374 GND.n2373 0.152939
R15840 GND.n2375 GND.n2374 0.152939
R15841 GND.n2376 GND.n2375 0.152939
R15842 GND.n2377 GND.n2376 0.152939
R15843 GND.n2378 GND.n2377 0.152939
R15844 GND.n2379 GND.n2378 0.152939
R15845 GND.n2380 GND.n2379 0.152939
R15846 GND.n2381 GND.n2380 0.152939
R15847 GND.n2382 GND.n2381 0.152939
R15848 GND.n2383 GND.n2382 0.152939
R15849 GND.n2385 GND.n2383 0.152939
R15850 GND.n2385 GND.n2384 0.152939
R15851 GND.n2128 GND.n2008 0.152939
R15852 GND.n2132 GND.n2128 0.152939
R15853 GND.n2133 GND.n2132 0.152939
R15854 GND.n2134 GND.n2133 0.152939
R15855 GND.n2134 GND.n2126 0.152939
R15856 GND.n2142 GND.n2126 0.152939
R15857 GND.n2143 GND.n2142 0.152939
R15858 GND.n2144 GND.n2143 0.152939
R15859 GND.n2144 GND.n2124 0.152939
R15860 GND.n2152 GND.n2124 0.152939
R15861 GND.n2153 GND.n2152 0.152939
R15862 GND.n2154 GND.n2153 0.152939
R15863 GND.n2154 GND.n2122 0.152939
R15864 GND.n2162 GND.n2122 0.152939
R15865 GND.n2163 GND.n2162 0.152939
R15866 GND.n2164 GND.n2163 0.152939
R15867 GND.n2164 GND.n2117 0.152939
R15868 GND.n2117 GND.n2113 0.152939
R15869 GND.n3985 GND.n2370 0.152939
R15870 GND.n3986 GND.n3985 0.152939
R15871 GND.n3987 GND.n3986 0.152939
R15872 GND.n3988 GND.n3987 0.152939
R15873 GND.n3988 GND.n2347 0.152939
R15874 GND.n4010 GND.n2347 0.152939
R15875 GND.n4011 GND.n4010 0.152939
R15876 GND.n4012 GND.n4011 0.152939
R15877 GND.n4013 GND.n4012 0.152939
R15878 GND.n4013 GND.n2324 0.152939
R15879 GND.n4034 GND.n2324 0.152939
R15880 GND.n4035 GND.n4034 0.152939
R15881 GND.n4036 GND.n4035 0.152939
R15882 GND.n4037 GND.n4036 0.152939
R15883 GND.n4037 GND.n2301 0.152939
R15884 GND.n4059 GND.n2301 0.152939
R15885 GND.n4060 GND.n4059 0.152939
R15886 GND.n4061 GND.n4060 0.152939
R15887 GND.n4063 GND.n4061 0.152939
R15888 GND.n4063 GND.n4062 0.152939
R15889 GND.n4062 GND.n2244 0.152939
R15890 GND.n3029 GND.n3026 0.152939
R15891 GND.n3030 GND.n3029 0.152939
R15892 GND.n3031 GND.n3030 0.152939
R15893 GND.n3032 GND.n3031 0.152939
R15894 GND.n3035 GND.n3032 0.152939
R15895 GND.n3036 GND.n3035 0.152939
R15896 GND.n3037 GND.n3036 0.152939
R15897 GND.n3038 GND.n3037 0.152939
R15898 GND.n3043 GND.n3038 0.152939
R15899 GND.n3044 GND.n3043 0.152939
R15900 GND.n3045 GND.n3044 0.152939
R15901 GND.n3046 GND.n3045 0.152939
R15902 GND.n3048 GND.n3046 0.152939
R15903 GND.n3048 GND.n3047 0.152939
R15904 GND.n3047 GND.n2614 0.152939
R15905 GND.n3191 GND.n2614 0.152939
R15906 GND.n3192 GND.n3191 0.152939
R15907 GND.n3193 GND.n3192 0.152939
R15908 GND.n3194 GND.n3193 0.152939
R15909 GND.n3195 GND.n3194 0.152939
R15910 GND.n3197 GND.n3195 0.152939
R15911 GND.n3197 GND.n3196 0.152939
R15912 GND.n3196 GND.n1643 0.152939
R15913 GND.n1644 GND.n1643 0.152939
R15914 GND.n1645 GND.n1644 0.152939
R15915 GND.n1674 GND.n1645 0.152939
R15916 GND.n1675 GND.n1674 0.152939
R15917 GND.n1676 GND.n1675 0.152939
R15918 GND.n1677 GND.n1676 0.152939
R15919 GND.n1678 GND.n1677 0.152939
R15920 GND.n1700 GND.n1678 0.152939
R15921 GND.n1701 GND.n1700 0.152939
R15922 GND.n1702 GND.n1701 0.152939
R15923 GND.n1703 GND.n1702 0.152939
R15924 GND.n1704 GND.n1703 0.152939
R15925 GND.n1727 GND.n1704 0.152939
R15926 GND.n1728 GND.n1727 0.152939
R15927 GND.n1729 GND.n1728 0.152939
R15928 GND.n1730 GND.n1729 0.152939
R15929 GND.n1731 GND.n1730 0.152939
R15930 GND.n2549 GND.n1731 0.152939
R15931 GND.n2550 GND.n2549 0.152939
R15932 GND.n2550 GND.n2547 0.152939
R15933 GND.n2556 GND.n2547 0.152939
R15934 GND.n2557 GND.n2556 0.152939
R15935 GND.n2558 GND.n2557 0.152939
R15936 GND.n2558 GND.n2543 0.152939
R15937 GND.n3521 GND.n2543 0.152939
R15938 GND.n3522 GND.n3521 0.152939
R15939 GND.n3523 GND.n3522 0.152939
R15940 GND.n3524 GND.n3523 0.152939
R15941 GND.n3525 GND.n3524 0.152939
R15942 GND.n3526 GND.n3525 0.152939
R15943 GND.n3527 GND.n3526 0.152939
R15944 GND.n3527 GND.n2525 0.152939
R15945 GND.n3587 GND.n2525 0.152939
R15946 GND.n3588 GND.n3587 0.152939
R15947 GND.n3589 GND.n3588 0.152939
R15948 GND.n3590 GND.n3589 0.152939
R15949 GND.n3591 GND.n3590 0.152939
R15950 GND.n3593 GND.n3591 0.152939
R15951 GND.n3593 GND.n3592 0.152939
R15952 GND.n3592 GND.n1849 0.152939
R15953 GND.n1850 GND.n1849 0.152939
R15954 GND.n1851 GND.n1850 0.152939
R15955 GND.n1893 GND.n1851 0.152939
R15956 GND.n1894 GND.n1893 0.152939
R15957 GND.n1899 GND.n1894 0.152939
R15958 GND.n1900 GND.n1899 0.152939
R15959 GND.n1901 GND.n1900 0.152939
R15960 GND.n1902 GND.n1901 0.152939
R15961 GND.n1903 GND.n1902 0.152939
R15962 GND.n1932 GND.n1903 0.152939
R15963 GND.n1935 GND.n1932 0.152939
R15964 GND.n1936 GND.n1935 0.152939
R15965 GND.n1937 GND.n1936 0.152939
R15966 GND.n1938 GND.n1937 0.152939
R15967 GND.n1939 GND.n1938 0.152939
R15968 GND.n2466 GND.n1939 0.152939
R15969 GND.n2467 GND.n2466 0.152939
R15970 GND.n2467 GND.n2464 0.152939
R15971 GND.n3820 GND.n2464 0.152939
R15972 GND.n3821 GND.n3820 0.152939
R15973 GND.n3822 GND.n3821 0.152939
R15974 GND.n3823 GND.n3822 0.152939
R15975 GND.n3823 GND.n2441 0.152939
R15976 GND.n3856 GND.n2441 0.152939
R15977 GND.n3857 GND.n3856 0.152939
R15978 GND.n3858 GND.n3857 0.152939
R15979 GND.n3858 GND.n2426 0.152939
R15980 GND.n3875 GND.n2426 0.152939
R15981 GND.n3876 GND.n3875 0.152939
R15982 GND.n3877 GND.n3876 0.152939
R15983 GND.n3877 GND.n2422 0.152939
R15984 GND.n3907 GND.n2422 0.152939
R15985 GND.n3908 GND.n3907 0.152939
R15986 GND.n3909 GND.n3908 0.152939
R15987 GND.n3909 GND.n2418 0.152939
R15988 GND.n3922 GND.n2418 0.152939
R15989 GND.n3923 GND.n3922 0.152939
R15990 GND.n3924 GND.n3923 0.152939
R15991 GND.n3925 GND.n3924 0.152939
R15992 GND.n3926 GND.n3925 0.152939
R15993 GND.n3929 GND.n3926 0.152939
R15994 GND.n3930 GND.n3929 0.152939
R15995 GND.n3931 GND.n3930 0.152939
R15996 GND.n3932 GND.n3931 0.152939
R15997 GND.n3935 GND.n3932 0.152939
R15998 GND.n3936 GND.n3935 0.152939
R15999 GND.n3937 GND.n3936 0.152939
R16000 GND.n3938 GND.n3937 0.152939
R16001 GND.n3941 GND.n3938 0.152939
R16002 GND.n3942 GND.n3941 0.152939
R16003 GND.n3943 GND.n3942 0.152939
R16004 GND.n3944 GND.n3943 0.152939
R16005 GND.n3947 GND.n3944 0.152939
R16006 GND.n3948 GND.n3947 0.152939
R16007 GND.n3949 GND.n3948 0.152939
R16008 GND.n3949 GND.n2260 0.152939
R16009 GND.n4147 GND.n2260 0.152939
R16010 GND.n3107 GND.n3106 0.152939
R16011 GND.n3107 GND.n2662 0.152939
R16012 GND.n3129 GND.n2662 0.152939
R16013 GND.n3130 GND.n3129 0.152939
R16014 GND.n3131 GND.n3130 0.152939
R16015 GND.n3132 GND.n3131 0.152939
R16016 GND.n3132 GND.n2643 0.152939
R16017 GND.n3154 GND.n2643 0.152939
R16018 GND.n3155 GND.n3154 0.152939
R16019 GND.n3156 GND.n3155 0.152939
R16020 GND.n3157 GND.n3156 0.152939
R16021 GND.n3157 GND.n2622 0.152939
R16022 GND.n3180 GND.n2622 0.152939
R16023 GND.n3181 GND.n3180 0.152939
R16024 GND.n3182 GND.n3181 0.152939
R16025 GND.n3182 GND.n2596 0.152939
R16026 GND.n3220 GND.n2596 0.152939
R16027 GND.n3221 GND.n3220 0.152939
R16028 GND.n3222 GND.n3221 0.152939
R16029 GND.n3222 GND.n1532 0.152939
R16030 GND.n4682 GND.n1532 0.152939
R16031 GND.n1380 GND.n1379 0.152939
R16032 GND.n1381 GND.n1380 0.152939
R16033 GND.n1382 GND.n1381 0.152939
R16034 GND.n1383 GND.n1382 0.152939
R16035 GND.n1384 GND.n1383 0.152939
R16036 GND.n1385 GND.n1384 0.152939
R16037 GND.n1386 GND.n1385 0.152939
R16038 GND.n1387 GND.n1386 0.152939
R16039 GND.n1388 GND.n1387 0.152939
R16040 GND.n1389 GND.n1388 0.152939
R16041 GND.n1390 GND.n1389 0.152939
R16042 GND.n1391 GND.n1390 0.152939
R16043 GND.n1392 GND.n1391 0.152939
R16044 GND.n1393 GND.n1392 0.152939
R16045 GND.n1394 GND.n1393 0.152939
R16046 GND.n1397 GND.n1394 0.152939
R16047 GND.n1398 GND.n1397 0.152939
R16048 GND.n1399 GND.n1398 0.152939
R16049 GND.n1400 GND.n1399 0.152939
R16050 GND.n1401 GND.n1400 0.152939
R16051 GND.n1402 GND.n1401 0.152939
R16052 GND.n1403 GND.n1402 0.152939
R16053 GND.n1404 GND.n1403 0.152939
R16054 GND.n1405 GND.n1404 0.152939
R16055 GND.n1406 GND.n1405 0.152939
R16056 GND.n1407 GND.n1406 0.152939
R16057 GND.n1408 GND.n1407 0.152939
R16058 GND.n1409 GND.n1408 0.152939
R16059 GND.n1410 GND.n1409 0.152939
R16060 GND.n1411 GND.n1410 0.152939
R16061 GND.n1412 GND.n1411 0.152939
R16062 GND.n4771 GND.n1412 0.152939
R16063 GND.n4771 GND.n4770 0.152939
R16064 GND.n4770 GND.n4769 0.152939
R16065 GND.n2906 GND.n2905 0.152939
R16066 GND.n2907 GND.n2906 0.152939
R16067 GND.n2907 GND.n2808 0.152939
R16068 GND.n2918 GND.n2808 0.152939
R16069 GND.n2919 GND.n2918 0.152939
R16070 GND.n2920 GND.n2919 0.152939
R16071 GND.n2920 GND.n2795 0.152939
R16072 GND.n2931 GND.n2795 0.152939
R16073 GND.n2932 GND.n2931 0.152939
R16074 GND.n2933 GND.n2932 0.152939
R16075 GND.n2933 GND.n2769 0.152939
R16076 GND.n2947 GND.n2769 0.152939
R16077 GND.n2948 GND.n2947 0.152939
R16078 GND.n2949 GND.n2948 0.152939
R16079 GND.n2950 GND.n2949 0.152939
R16080 GND.n2950 GND.n2746 0.152939
R16081 GND.n2984 GND.n2746 0.152939
R16082 GND.n2985 GND.n2984 0.152939
R16083 GND.n2986 GND.n2985 0.152939
R16084 GND.n2986 GND.n2683 0.152939
R16085 GND.n3106 GND.n2683 0.152939
R16086 GND.n2777 GND.n2776 0.152939
R16087 GND.n2778 GND.n2777 0.152939
R16088 GND.n2780 GND.n2778 0.152939
R16089 GND.n2781 GND.n2780 0.152939
R16090 GND.n2781 GND.n2734 0.152939
R16091 GND.n2994 GND.n2734 0.152939
R16092 GND.n2995 GND.n2994 0.152939
R16093 GND.n2996 GND.n2995 0.152939
R16094 GND.n1226 GND.n1225 0.152939
R16095 GND.n1227 GND.n1226 0.152939
R16096 GND.n1232 GND.n1227 0.152939
R16097 GND.n1233 GND.n1232 0.152939
R16098 GND.n1234 GND.n1233 0.152939
R16099 GND.n1235 GND.n1234 0.152939
R16100 GND.n1240 GND.n1235 0.152939
R16101 GND.n1241 GND.n1240 0.152939
R16102 GND.n1242 GND.n1241 0.152939
R16103 GND.n1243 GND.n1242 0.152939
R16104 GND.n1248 GND.n1243 0.152939
R16105 GND.n1249 GND.n1248 0.152939
R16106 GND.n1250 GND.n1249 0.152939
R16107 GND.n1251 GND.n1250 0.152939
R16108 GND.n1256 GND.n1251 0.152939
R16109 GND.n1257 GND.n1256 0.152939
R16110 GND.n1258 GND.n1257 0.152939
R16111 GND.n1259 GND.n1258 0.152939
R16112 GND.n1264 GND.n1259 0.152939
R16113 GND.n1265 GND.n1264 0.152939
R16114 GND.n1266 GND.n1265 0.152939
R16115 GND.n1267 GND.n1266 0.152939
R16116 GND.n1272 GND.n1267 0.152939
R16117 GND.n1273 GND.n1272 0.152939
R16118 GND.n1274 GND.n1273 0.152939
R16119 GND.n1275 GND.n1274 0.152939
R16120 GND.n1280 GND.n1275 0.152939
R16121 GND.n1281 GND.n1280 0.152939
R16122 GND.n1282 GND.n1281 0.152939
R16123 GND.n1283 GND.n1282 0.152939
R16124 GND.n1288 GND.n1283 0.152939
R16125 GND.n1289 GND.n1288 0.152939
R16126 GND.n1290 GND.n1289 0.152939
R16127 GND.n1291 GND.n1290 0.152939
R16128 GND.n1296 GND.n1291 0.152939
R16129 GND.n1297 GND.n1296 0.152939
R16130 GND.n1298 GND.n1297 0.152939
R16131 GND.n1299 GND.n1298 0.152939
R16132 GND.n1304 GND.n1299 0.152939
R16133 GND.n1305 GND.n1304 0.152939
R16134 GND.n1306 GND.n1305 0.152939
R16135 GND.n1307 GND.n1306 0.152939
R16136 GND.n1312 GND.n1307 0.152939
R16137 GND.n1313 GND.n1312 0.152939
R16138 GND.n1314 GND.n1313 0.152939
R16139 GND.n1315 GND.n1314 0.152939
R16140 GND.n1320 GND.n1315 0.152939
R16141 GND.n1321 GND.n1320 0.152939
R16142 GND.n1322 GND.n1321 0.152939
R16143 GND.n1323 GND.n1322 0.152939
R16144 GND.n1328 GND.n1323 0.152939
R16145 GND.n1329 GND.n1328 0.152939
R16146 GND.n1330 GND.n1329 0.152939
R16147 GND.n1331 GND.n1330 0.152939
R16148 GND.n1336 GND.n1331 0.152939
R16149 GND.n1337 GND.n1336 0.152939
R16150 GND.n1338 GND.n1337 0.152939
R16151 GND.n1339 GND.n1338 0.152939
R16152 GND.n1344 GND.n1339 0.152939
R16153 GND.n1345 GND.n1344 0.152939
R16154 GND.n1346 GND.n1345 0.152939
R16155 GND.n1347 GND.n1346 0.152939
R16156 GND.n2775 GND.n1347 0.152939
R16157 GND.n3915 GND.n3914 0.152939
R16158 GND.n3914 GND.n2359 0.152939
R16159 GND.n3995 GND.n2359 0.152939
R16160 GND.n3996 GND.n3995 0.152939
R16161 GND.n3998 GND.n3996 0.152939
R16162 GND.n3998 GND.n3997 0.152939
R16163 GND.n3997 GND.n2337 0.152939
R16164 GND.n4020 GND.n2337 0.152939
R16165 GND.n4021 GND.n4020 0.152939
R16166 GND.n4023 GND.n4021 0.152939
R16167 GND.n4023 GND.n4022 0.152939
R16168 GND.n4022 GND.n2313 0.152939
R16169 GND.n4044 GND.n2313 0.152939
R16170 GND.n4045 GND.n4044 0.152939
R16171 GND.n4047 GND.n4045 0.152939
R16172 GND.n4047 GND.n4046 0.152939
R16173 GND.n4046 GND.n2286 0.152939
R16174 GND.n4070 GND.n2286 0.152939
R16175 GND.n4071 GND.n4070 0.152939
R16176 GND.n4072 GND.n4071 0.152939
R16177 GND.n4072 GND.n2283 0.152939
R16178 GND.n4078 GND.n2283 0.152939
R16179 GND.n4079 GND.n4078 0.152939
R16180 GND.n4080 GND.n4079 0.152939
R16181 GND.n4080 GND.n674 0.152939
R16182 GND.n5753 GND.n675 0.152939
R16183 GND.n5753 GND.n5752 0.152939
R16184 GND.n5752 GND.n5751 0.152939
R16185 GND.n5751 GND.n681 0.152939
R16186 GND.n5747 GND.n681 0.152939
R16187 GND.n5747 GND.n5746 0.152939
R16188 GND.n5746 GND.n5745 0.152939
R16189 GND.n5745 GND.n686 0.152939
R16190 GND.n5741 GND.n686 0.152939
R16191 GND.n5741 GND.n5740 0.152939
R16192 GND.n5740 GND.n5739 0.152939
R16193 GND.n5739 GND.n691 0.152939
R16194 GND.n5735 GND.n691 0.152939
R16195 GND.n5735 GND.n5734 0.152939
R16196 GND.n5734 GND.n5733 0.152939
R16197 GND.n5733 GND.n696 0.152939
R16198 GND.n5729 GND.n696 0.152939
R16199 GND.n5729 GND.n5728 0.152939
R16200 GND.n5728 GND.n5727 0.152939
R16201 GND.n5727 GND.n701 0.152939
R16202 GND.n5723 GND.n701 0.152939
R16203 GND.n5723 GND.n5722 0.152939
R16204 GND.n5722 GND.n5721 0.152939
R16205 GND.n5721 GND.n706 0.152939
R16206 GND.n5717 GND.n706 0.152939
R16207 GND.n5649 GND.n5648 0.152939
R16208 GND.n5648 GND.n5647 0.152939
R16209 GND.n5647 GND.n5608 0.152939
R16210 GND.n5643 GND.n5608 0.152939
R16211 GND.n5643 GND.n5642 0.152939
R16212 GND.n5642 GND.n5641 0.152939
R16213 GND.n5641 GND.n5614 0.152939
R16214 GND.n5637 GND.n5614 0.152939
R16215 GND.n5637 GND.n5636 0.152939
R16216 GND.n5636 GND.n5635 0.152939
R16217 GND.n5635 GND.n5620 0.152939
R16218 GND.n5631 GND.n5620 0.152939
R16219 GND.n5631 GND.n5630 0.152939
R16220 GND.n5630 GND.n5629 0.152939
R16221 GND.n5629 GND.n710 0.152939
R16222 GND.n5716 GND.n710 0.152939
R16223 GND.n5710 GND.n5709 0.152939
R16224 GND.n5709 GND.n5708 0.152939
R16225 GND.n5708 GND.n746 0.152939
R16226 GND.n5704 GND.n746 0.152939
R16227 GND.n5704 GND.n5703 0.152939
R16228 GND.n5703 GND.n5702 0.152939
R16229 GND.n5702 GND.n752 0.152939
R16230 GND.n5698 GND.n752 0.152939
R16231 GND.n5698 GND.n5697 0.152939
R16232 GND.n5697 GND.n5696 0.152939
R16233 GND.n5696 GND.n758 0.152939
R16234 GND.n5692 GND.n758 0.152939
R16235 GND.n5692 GND.n5691 0.152939
R16236 GND.n5691 GND.n5690 0.152939
R16237 GND.n5690 GND.n764 0.152939
R16238 GND.n5685 GND.n764 0.152939
R16239 GND.n5685 GND.n5684 0.152939
R16240 GND.n5684 GND.n5683 0.152939
R16241 GND.n5683 GND.n772 0.152939
R16242 GND.n5679 GND.n772 0.152939
R16243 GND.n5679 GND.n5678 0.152939
R16244 GND.n5678 GND.n5677 0.152939
R16245 GND.n5677 GND.n778 0.152939
R16246 GND.n5673 GND.n778 0.152939
R16247 GND.n5673 GND.n5672 0.152939
R16248 GND.n5672 GND.n5671 0.152939
R16249 GND.n5671 GND.n784 0.152939
R16250 GND.n5667 GND.n784 0.152939
R16251 GND.n5667 GND.n5666 0.152939
R16252 GND.n5666 GND.n5665 0.152939
R16253 GND.n5665 GND.n790 0.152939
R16254 GND.n5661 GND.n790 0.152939
R16255 GND.n5661 GND.n5660 0.152939
R16256 GND.n5660 GND.n5659 0.152939
R16257 GND.n4255 GND.n4254 0.152939
R16258 GND.n4254 GND.n4253 0.152939
R16259 GND.n4253 GND.n2091 0.152939
R16260 GND.n4249 GND.n2091 0.152939
R16261 GND.n4249 GND.n4248 0.152939
R16262 GND.n4248 GND.n4247 0.152939
R16263 GND.n4247 GND.n2096 0.152939
R16264 GND.n4243 GND.n2096 0.152939
R16265 GND.n4243 GND.n4242 0.152939
R16266 GND.n3267 GND.n2583 0.152939
R16267 GND.n3275 GND.n2583 0.152939
R16268 GND.n3276 GND.n3275 0.152939
R16269 GND.n3277 GND.n3276 0.152939
R16270 GND.n3277 GND.n2579 0.152939
R16271 GND.n3283 GND.n2579 0.152939
R16272 GND.n3284 GND.n3283 0.152939
R16273 GND.n3285 GND.n3284 0.152939
R16274 GND.n3285 GND.n2577 0.152939
R16275 GND.n3291 GND.n2577 0.152939
R16276 GND.n3292 GND.n3291 0.152939
R16277 GND.n3293 GND.n3292 0.152939
R16278 GND.n3293 GND.n2571 0.152939
R16279 GND.n3483 GND.n2571 0.152939
R16280 GND.n3484 GND.n3483 0.152939
R16281 GND.n3485 GND.n3484 0.152939
R16282 GND.n3485 GND.n2566 0.152939
R16283 GND.n3512 GND.n2566 0.152939
R16284 GND.n3512 GND.n3511 0.152939
R16285 GND.n3511 GND.n3510 0.152939
R16286 GND.n3510 GND.n2567 0.152939
R16287 GND.n3506 GND.n2567 0.152939
R16288 GND.n3506 GND.n2534 0.152939
R16289 GND.n3552 GND.n2534 0.152939
R16290 GND.n3553 GND.n3552 0.152939
R16291 GND.n3565 GND.n3553 0.152939
R16292 GND.n3565 GND.n3564 0.152939
R16293 GND.n3564 GND.n3563 0.152939
R16294 GND.n3563 GND.n3554 0.152939
R16295 GND.n3559 GND.n3554 0.152939
R16296 GND.n3559 GND.n2518 0.152939
R16297 GND.n3615 GND.n2518 0.152939
R16298 GND.n3616 GND.n3615 0.152939
R16299 GND.n3619 GND.n3616 0.152939
R16300 GND.n3619 GND.n3618 0.152939
R16301 GND.n3618 GND.n3617 0.152939
R16302 GND.n3617 GND.n2504 0.152939
R16303 GND.n3652 GND.n2504 0.152939
R16304 GND.n3653 GND.n3652 0.152939
R16305 GND.n3658 GND.n3653 0.152939
R16306 GND.n3658 GND.n3657 0.152939
R16307 GND.n3657 GND.n3656 0.152939
R16308 GND.n3656 GND.n2486 0.152939
R16309 GND.n3688 GND.n2486 0.152939
R16310 GND.n3689 GND.n3688 0.152939
R16311 GND.n3703 GND.n3689 0.152939
R16312 GND.n3703 GND.n3702 0.152939
R16313 GND.n3702 GND.n3701 0.152939
R16314 GND.n3701 GND.n3690 0.152939
R16315 GND.n3697 GND.n3690 0.152939
R16316 GND.n3697 GND.n3696 0.152939
R16317 GND.n3696 GND.n2475 0.152939
R16318 GND.n3809 GND.n2475 0.152939
R16319 GND.n3810 GND.n3809 0.152939
R16320 GND.n3812 GND.n3810 0.152939
R16321 GND.n3812 GND.n3811 0.152939
R16322 GND.n3811 GND.n2448 0.152939
R16323 GND.n3841 GND.n2448 0.152939
R16324 GND.n3842 GND.n3841 0.152939
R16325 GND.n3849 GND.n3842 0.152939
R16326 GND.n3849 GND.n3848 0.152939
R16327 GND.n3848 GND.n3847 0.152939
R16328 GND.n3847 GND.n3843 0.152939
R16329 GND.n3843 GND.n2104 0.152939
R16330 GND.n4241 GND.n2104 0.152939
R16331 GND.n3244 GND.n2588 0.152939
R16332 GND.n3245 GND.n3244 0.152939
R16333 GND.n3246 GND.n3245 0.152939
R16334 GND.n3246 GND.n2586 0.152939
R16335 GND.n3257 GND.n2586 0.152939
R16336 GND.n3258 GND.n3257 0.152939
R16337 GND.n3259 GND.n3258 0.152939
R16338 GND.n3259 GND.n2584 0.152939
R16339 GND.n3266 GND.n2584 0.152939
R16340 GND.n3017 GND.n3016 0.152939
R16341 GND.n3018 GND.n3017 0.152939
R16342 GND.n3018 GND.n2673 0.152939
R16343 GND.n3114 GND.n2673 0.152939
R16344 GND.n3115 GND.n3114 0.152939
R16345 GND.n3117 GND.n3115 0.152939
R16346 GND.n3117 GND.n3116 0.152939
R16347 GND.n3116 GND.n2653 0.152939
R16348 GND.n3139 GND.n2653 0.152939
R16349 GND.n3140 GND.n3139 0.152939
R16350 GND.n3142 GND.n3140 0.152939
R16351 GND.n3142 GND.n3141 0.152939
R16352 GND.n3141 GND.n2633 0.152939
R16353 GND.n3164 GND.n2633 0.152939
R16354 GND.n3165 GND.n3164 0.152939
R16355 GND.n3170 GND.n3165 0.152939
R16356 GND.n3170 GND.n3169 0.152939
R16357 GND.n3169 GND.n3168 0.152939
R16358 GND.n3168 GND.n2608 0.152939
R16359 GND.n3211 GND.n2608 0.152939
R16360 GND.n3211 GND.n3210 0.152939
R16361 GND.n3210 GND.n3209 0.152939
R16362 GND.n3209 GND.n2609 0.152939
R16363 GND.n2609 GND.n2589 0.152939
R16364 GND.n3234 GND.n2589 0.152939
R16365 GND.n4681 GND.n1533 0.152939
R16366 GND.n4677 GND.n1533 0.152939
R16367 GND.n4677 GND.n4676 0.152939
R16368 GND.n4676 GND.n4675 0.152939
R16369 GND.n4675 GND.n1537 0.152939
R16370 GND.n4671 GND.n1537 0.152939
R16371 GND.n4671 GND.n4670 0.152939
R16372 GND.n4670 GND.n4669 0.152939
R16373 GND.n4669 GND.n1542 0.152939
R16374 GND.n4665 GND.n1542 0.152939
R16375 GND.n4665 GND.n4664 0.152939
R16376 GND.n4664 GND.n4663 0.152939
R16377 GND.n4663 GND.n1547 0.152939
R16378 GND.n4658 GND.n4657 0.152939
R16379 GND.n4657 GND.n4656 0.152939
R16380 GND.n4656 GND.n1557 0.152939
R16381 GND.n4652 GND.n1557 0.152939
R16382 GND.n4652 GND.n4651 0.152939
R16383 GND.n4651 GND.n4650 0.152939
R16384 GND.n4650 GND.n1562 0.152939
R16385 GND.n4646 GND.n1562 0.152939
R16386 GND.n4646 GND.n4645 0.152939
R16387 GND.n4645 GND.n4644 0.152939
R16388 GND.n4644 GND.n1567 0.152939
R16389 GND.n4640 GND.n1567 0.152939
R16390 GND.n4640 GND.n4639 0.152939
R16391 GND.n4639 GND.n4638 0.152939
R16392 GND.n4638 GND.n1572 0.152939
R16393 GND.n4634 GND.n1572 0.152939
R16394 GND.n4634 GND.n4633 0.152939
R16395 GND.n4633 GND.n4632 0.152939
R16396 GND.n2842 GND.n2841 0.152939
R16397 GND.n2843 GND.n2842 0.152939
R16398 GND.n2843 GND.n2834 0.152939
R16399 GND.n2849 GND.n2834 0.152939
R16400 GND.n2850 GND.n2849 0.152939
R16401 GND.n2851 GND.n2850 0.152939
R16402 GND.n2851 GND.n2830 0.152939
R16403 GND.n2857 GND.n2830 0.152939
R16404 GND.n2858 GND.n2857 0.152939
R16405 GND.n2859 GND.n2858 0.152939
R16406 GND.n2859 GND.n2826 0.152939
R16407 GND.n2865 GND.n2826 0.152939
R16408 GND.n2866 GND.n2865 0.152939
R16409 GND.n2867 GND.n2866 0.152939
R16410 GND.n2867 GND.n2819 0.152939
R16411 GND.n2871 GND.n2819 0.152939
R16412 GND.n2875 GND.n2874 0.152939
R16413 GND.n2899 GND.n2875 0.152939
R16414 GND.n2899 GND.n2898 0.152939
R16415 GND.n2898 GND.n2897 0.152939
R16416 GND.n2897 GND.n2876 0.152939
R16417 GND.n2893 GND.n2876 0.152939
R16418 GND.n2893 GND.n2892 0.152939
R16419 GND.n2892 GND.n2891 0.152939
R16420 GND.n2891 GND.n2880 0.152939
R16421 GND.n2887 GND.n2880 0.152939
R16422 GND.n2887 GND.n2886 0.152939
R16423 GND.n2886 GND.n2885 0.152939
R16424 GND.n2885 GND.n2759 0.152939
R16425 GND.n2957 GND.n2759 0.152939
R16426 GND.n2958 GND.n2957 0.152939
R16427 GND.n2974 GND.n2958 0.152939
R16428 GND.n2974 GND.n2973 0.152939
R16429 GND.n2973 GND.n2972 0.152939
R16430 GND.n2972 GND.n2959 0.152939
R16431 GND.n2968 GND.n2959 0.152939
R16432 GND.n2968 GND.n2967 0.152939
R16433 GND.n2967 GND.n2726 0.152939
R16434 GND.n3008 GND.n2726 0.152939
R16435 GND.n3009 GND.n3008 0.152939
R16436 GND.n3010 GND.n3009 0.152939
R16437 GND.n4149 GND.n4148 0.146841
R16438 GND.n2996 GND.n2684 0.146841
R16439 GND.n5757 GND.n674 0.145814
R16440 GND.n5757 GND.n675 0.145814
R16441 GND.n3016 GND.n2724 0.145814
R16442 GND.n3010 GND.n2724 0.145814
R16443 GND.n4255 GND.n2090 0.145317
R16444 GND.n3235 GND.n2588 0.145317
R16445 GND.n4233 GND.n4232 0.0429592
R16446 GND.n5654 GND.n798 0.0429592
R16447 GND.n4764 GND.n1418 0.0429592
R16448 GND.n4630 GND.n1523 0.0429592
R16449 GND.n4232 GND.n2115 0.0344674
R16450 GND.n4228 GND.n2115 0.0344674
R16451 GND.n4228 GND.n4227 0.0344674
R16452 GND.n4227 GND.n4226 0.0344674
R16453 GND.n4226 GND.n2176 0.0344674
R16454 GND.n4222 GND.n2176 0.0344674
R16455 GND.n4222 GND.n4221 0.0344674
R16456 GND.n4221 GND.n4220 0.0344674
R16457 GND.n4220 GND.n2184 0.0344674
R16458 GND.n4216 GND.n2184 0.0344674
R16459 GND.n4216 GND.n4215 0.0344674
R16460 GND.n4215 GND.n4214 0.0344674
R16461 GND.n4214 GND.n2192 0.0344674
R16462 GND.n4210 GND.n2192 0.0344674
R16463 GND.n4210 GND.n4209 0.0344674
R16464 GND.n4209 GND.n4208 0.0344674
R16465 GND.n4208 GND.n2200 0.0344674
R16466 GND.n4204 GND.n2200 0.0344674
R16467 GND.n4204 GND.n4203 0.0344674
R16468 GND.n4203 GND.n4202 0.0344674
R16469 GND.n4202 GND.n2208 0.0344674
R16470 GND.n4198 GND.n2208 0.0344674
R16471 GND.n4198 GND.n4197 0.0344674
R16472 GND.n4197 GND.n4196 0.0344674
R16473 GND.n4196 GND.n2216 0.0344674
R16474 GND.n4192 GND.n2216 0.0344674
R16475 GND.n4192 GND.n4191 0.0344674
R16476 GND.n4191 GND.n4190 0.0344674
R16477 GND.n4190 GND.n2224 0.0344674
R16478 GND.n4186 GND.n2224 0.0344674
R16479 GND.n4186 GND.n4185 0.0344674
R16480 GND.n4185 GND.n4184 0.0344674
R16481 GND.n4184 GND.n2232 0.0344674
R16482 GND.n4180 GND.n2232 0.0344674
R16483 GND.n4180 GND.n4179 0.0344674
R16484 GND.n4179 GND.n875 0.0344674
R16485 GND.n5541 GND.n875 0.0344674
R16486 GND.n5541 GND.n878 0.0344674
R16487 GND.n878 GND.n877 0.0344674
R16488 GND.n877 GND.n854 0.0344674
R16489 GND.n5558 GND.n854 0.0344674
R16490 GND.n5558 GND.n857 0.0344674
R16491 GND.n857 GND.n856 0.0344674
R16492 GND.n856 GND.n834 0.0344674
R16493 GND.n5575 GND.n834 0.0344674
R16494 GND.n5575 GND.n837 0.0344674
R16495 GND.n837 GND.n836 0.0344674
R16496 GND.n836 GND.n816 0.0344674
R16497 GND.n5593 GND.n816 0.0344674
R16498 GND.n5593 GND.n817 0.0344674
R16499 GND.n817 GND.n801 0.0344674
R16500 GND.n5654 GND.n801 0.0344674
R16501 GND.n4304 GND.n2041 0.0344674
R16502 GND.n4259 GND.n2085 0.0344674
R16503 GND.n4628 GND.n1580 0.0344674
R16504 GND.n3236 GND.n1625 0.0344674
R16505 GND.n4764 GND.n4763 0.0344674
R16506 GND.n4763 GND.n4762 0.0344674
R16507 GND.n4762 GND.n1424 0.0344674
R16508 GND.n4758 GND.n1424 0.0344674
R16509 GND.n4758 GND.n4757 0.0344674
R16510 GND.n4757 GND.n4756 0.0344674
R16511 GND.n4756 GND.n1432 0.0344674
R16512 GND.n4752 GND.n1432 0.0344674
R16513 GND.n4752 GND.n4751 0.0344674
R16514 GND.n4751 GND.n4750 0.0344674
R16515 GND.n4750 GND.n1440 0.0344674
R16516 GND.n4746 GND.n1440 0.0344674
R16517 GND.n4746 GND.n4745 0.0344674
R16518 GND.n4745 GND.n4744 0.0344674
R16519 GND.n4744 GND.n1448 0.0344674
R16520 GND.n4740 GND.n1448 0.0344674
R16521 GND.n4740 GND.n4739 0.0344674
R16522 GND.n4739 GND.n4738 0.0344674
R16523 GND.n4738 GND.n1456 0.0344674
R16524 GND.n4734 GND.n1456 0.0344674
R16525 GND.n4734 GND.n4733 0.0344674
R16526 GND.n4733 GND.n4732 0.0344674
R16527 GND.n4732 GND.n1464 0.0344674
R16528 GND.n4728 GND.n1464 0.0344674
R16529 GND.n4728 GND.n4727 0.0344674
R16530 GND.n4727 GND.n4726 0.0344674
R16531 GND.n4726 GND.n1472 0.0344674
R16532 GND.n4722 GND.n1472 0.0344674
R16533 GND.n4722 GND.n4721 0.0344674
R16534 GND.n4721 GND.n4720 0.0344674
R16535 GND.n4720 GND.n1480 0.0344674
R16536 GND.n4716 GND.n1480 0.0344674
R16537 GND.n4716 GND.n4715 0.0344674
R16538 GND.n4715 GND.n4714 0.0344674
R16539 GND.n4714 GND.n1488 0.0344674
R16540 GND.n4710 GND.n1488 0.0344674
R16541 GND.n4710 GND.n4709 0.0344674
R16542 GND.n4709 GND.n4708 0.0344674
R16543 GND.n4708 GND.n1496 0.0344674
R16544 GND.n4704 GND.n1496 0.0344674
R16545 GND.n4704 GND.n4703 0.0344674
R16546 GND.n4703 GND.n4702 0.0344674
R16547 GND.n4702 GND.n1504 0.0344674
R16548 GND.n4698 GND.n1504 0.0344674
R16549 GND.n4698 GND.n4697 0.0344674
R16550 GND.n4697 GND.n4696 0.0344674
R16551 GND.n4696 GND.n1512 0.0344674
R16552 GND.n4692 GND.n1512 0.0344674
R16553 GND.n4692 GND.n4691 0.0344674
R16554 GND.n4691 GND.n4690 0.0344674
R16555 GND.n4690 GND.n1520 0.0344674
R16556 GND.n1523 GND.n1520 0.0344674
R16557 GND.n4303 GND.n2043 0.0188424
R16558 GND.n4300 GND.n4299 0.0188424
R16559 GND.n4296 GND.n2047 0.0188424
R16560 GND.n4295 GND.n2053 0.0188424
R16561 GND.n4292 GND.n4291 0.0188424
R16562 GND.n4288 GND.n2057 0.0188424
R16563 GND.n4287 GND.n2061 0.0188424
R16564 GND.n4284 GND.n4283 0.0188424
R16565 GND.n4280 GND.n2065 0.0188424
R16566 GND.n4279 GND.n2071 0.0188424
R16567 GND.n4276 GND.n4275 0.0188424
R16568 GND.n4272 GND.n2075 0.0188424
R16569 GND.n4271 GND.n2079 0.0188424
R16570 GND.n4268 GND.n4267 0.0188424
R16571 GND.n4260 GND.n2083 0.0188424
R16572 GND.n4624 GND.n1585 0.0188424
R16573 GND.n4623 GND.n1586 0.0188424
R16574 GND.n4620 GND.n4619 0.0188424
R16575 GND.n4616 GND.n1591 0.0188424
R16576 GND.n4615 GND.n1595 0.0188424
R16577 GND.n4612 GND.n4611 0.0188424
R16578 GND.n4608 GND.n1599 0.0188424
R16579 GND.n4607 GND.n1603 0.0188424
R16580 GND.n4604 GND.n4603 0.0188424
R16581 GND.n4600 GND.n1607 0.0188424
R16582 GND.n4599 GND.n1611 0.0188424
R16583 GND.n4596 GND.n4595 0.0188424
R16584 GND.n4592 GND.n1615 0.0188424
R16585 GND.n4591 GND.n1621 0.0188424
R16586 GND.n4588 GND.n4587 0.0188424
R16587 GND.n4304 GND.n4303 0.016125
R16588 GND.n4300 GND.n2043 0.016125
R16589 GND.n4299 GND.n2047 0.016125
R16590 GND.n4296 GND.n4295 0.016125
R16591 GND.n4292 GND.n2053 0.016125
R16592 GND.n4291 GND.n2057 0.016125
R16593 GND.n4288 GND.n4287 0.016125
R16594 GND.n4284 GND.n2061 0.016125
R16595 GND.n4283 GND.n2065 0.016125
R16596 GND.n4280 GND.n4279 0.016125
R16597 GND.n4276 GND.n2071 0.016125
R16598 GND.n4275 GND.n2075 0.016125
R16599 GND.n4272 GND.n4271 0.016125
R16600 GND.n4268 GND.n2079 0.016125
R16601 GND.n4267 GND.n2083 0.016125
R16602 GND.n4260 GND.n4259 0.016125
R16603 GND.n1585 GND.n1580 0.016125
R16604 GND.n4624 GND.n4623 0.016125
R16605 GND.n4620 GND.n1586 0.016125
R16606 GND.n4619 GND.n1591 0.016125
R16607 GND.n4616 GND.n4615 0.016125
R16608 GND.n4612 GND.n1595 0.016125
R16609 GND.n4611 GND.n1599 0.016125
R16610 GND.n4608 GND.n4607 0.016125
R16611 GND.n4604 GND.n1603 0.016125
R16612 GND.n4603 GND.n1607 0.016125
R16613 GND.n4600 GND.n4599 0.016125
R16614 GND.n4596 GND.n1611 0.016125
R16615 GND.n4595 GND.n1615 0.016125
R16616 GND.n4592 GND.n4591 0.016125
R16617 GND.n4588 GND.n1621 0.016125
R16618 GND.n4587 GND.n1625 0.016125
R16619 GND.n3026 GND.n2684 0.00659756
R16620 GND.n4148 GND.n4147 0.00659756
R16621 GND.n4234 GND.n2041 0.00457609
R16622 GND.n4629 GND.n4628 0.00457609
R16623 GND.n2090 GND.n2085 0.00219837
R16624 GND.n3236 GND.n3235 0.00219837
R16625 VN.n28 VN.t0 243.97
R16626 VN.n28 VN.n27 223.454
R16627 VN.n30 VN.n29 223.454
R16628 VN.n15 VN.t7 199.144
R16629 VN.n2 VN.t5 199.144
R16630 VN.n24 VN.t10 183.883
R16631 VN.n11 VN.t9 183.883
R16632 VN.n23 VN.n13 161.3
R16633 VN.n21 VN.n20 161.3
R16634 VN.n19 VN.n14 161.3
R16635 VN.n18 VN.n17 161.3
R16636 VN.n5 VN.n4 161.3
R16637 VN.n6 VN.n1 161.3
R16638 VN.n8 VN.n7 161.3
R16639 VN.n10 VN.n0 161.3
R16640 VN.n16 VN.t6 144.601
R16641 VN.n22 VN.t11 144.601
R16642 VN.n9 VN.t8 144.601
R16643 VN.n3 VN.t12 144.601
R16644 VN.n25 VN.n24 80.6037
R16645 VN.n12 VN.n11 80.6037
R16646 VN.n24 VN.n23 56.3158
R16647 VN.n11 VN.n10 56.3158
R16648 VN.n16 VN.n15 46.9082
R16649 VN.n3 VN.n2 46.9082
R16650 VN.n18 VN.n15 43.8991
R16651 VN.n5 VN.n2 43.8991
R16652 VN.n17 VN.n14 40.577
R16653 VN.n21 VN.n14 40.577
R16654 VN.n8 VN.n1 40.577
R16655 VN.n4 VN.n1 40.577
R16656 VN.n26 VN.n25 27.893
R16657 VN.n27 VN.t1 19.8005
R16658 VN.n27 VN.t4 19.8005
R16659 VN.n29 VN.t2 19.8005
R16660 VN.n29 VN.t3 19.8005
R16661 VN.n23 VN.n22 16.477
R16662 VN.n10 VN.n9 16.477
R16663 VN VN.n31 13.8471
R16664 VN.n26 VN.n12 11.6998
R16665 VN.n17 VN.n16 8.11581
R16666 VN.n22 VN.n21 8.11581
R16667 VN.n9 VN.n8 8.11581
R16668 VN.n4 VN.n3 8.11581
R16669 VN.n31 VN.n30 5.40567
R16670 VN.n31 VN.n26 1.188
R16671 VN.n30 VN.n28 0.716017
R16672 VN.n25 VN.n13 0.285035
R16673 VN.n12 VN.n0 0.285035
R16674 VN.n19 VN.n18 0.189894
R16675 VN.n20 VN.n19 0.189894
R16676 VN.n20 VN.n13 0.189894
R16677 VN.n7 VN.n0 0.189894
R16678 VN.n7 VN.n6 0.189894
R16679 VN.n6 VN.n5 0.189894
R16680 a_n1455_n3628.n350 a_n1455_n3628.n330 289.615
R16681 a_n1455_n3628.n60 a_n1455_n3628.n40 289.615
R16682 a_n1455_n3628.n112 a_n1455_n3628.n92 289.615
R16683 a_n1455_n3628.n140 a_n1455_n3628.n120 289.615
R16684 a_n1455_n3628.n86 a_n1455_n3628.n66 289.615
R16685 a_n1455_n3628.n191 a_n1455_n3628.n171 289.615
R16686 a_n1455_n3628.n217 a_n1455_n3628.n197 289.615
R16687 a_n1455_n3628.n166 a_n1455_n3628.n146 289.615
R16688 a_n1455_n3628.n324 a_n1455_n3628.n304 289.615
R16689 a_n1455_n3628.n297 a_n1455_n3628.n277 289.615
R16690 a_n1455_n3628.n272 a_n1455_n3628.n252 289.615
R16691 a_n1455_n3628.n245 a_n1455_n3628.n225 289.615
R16692 a_n1455_n3628.n223 a_n1455_n3628.n170 196.838
R16693 a_n1455_n3628.n91 a_n1455_n3628.n90 196.298
R16694 a_n1455_n3628.n196 a_n1455_n3628.n195 196.298
R16695 a_n1455_n3628.n222 a_n1455_n3628.n221 196.298
R16696 a_n1455_n3628.n351 a_n1455_n3628.n350 185
R16697 a_n1455_n3628.n349 a_n1455_n3628.n348 185
R16698 a_n1455_n3628.n333 a_n1455_n3628.n332 185
R16699 a_n1455_n3628.n345 a_n1455_n3628.n344 185
R16700 a_n1455_n3628.n343 a_n1455_n3628.n342 185
R16701 a_n1455_n3628.n336 a_n1455_n3628.n335 185
R16702 a_n1455_n3628.n339 a_n1455_n3628.n338 185
R16703 a_n1455_n3628.n61 a_n1455_n3628.n60 185
R16704 a_n1455_n3628.n59 a_n1455_n3628.n58 185
R16705 a_n1455_n3628.n43 a_n1455_n3628.n42 185
R16706 a_n1455_n3628.n55 a_n1455_n3628.n54 185
R16707 a_n1455_n3628.n53 a_n1455_n3628.n52 185
R16708 a_n1455_n3628.n46 a_n1455_n3628.n45 185
R16709 a_n1455_n3628.n49 a_n1455_n3628.n48 185
R16710 a_n1455_n3628.n113 a_n1455_n3628.n112 185
R16711 a_n1455_n3628.n111 a_n1455_n3628.n110 185
R16712 a_n1455_n3628.n95 a_n1455_n3628.n94 185
R16713 a_n1455_n3628.n107 a_n1455_n3628.n106 185
R16714 a_n1455_n3628.n105 a_n1455_n3628.n104 185
R16715 a_n1455_n3628.n98 a_n1455_n3628.n97 185
R16716 a_n1455_n3628.n101 a_n1455_n3628.n100 185
R16717 a_n1455_n3628.n141 a_n1455_n3628.n140 185
R16718 a_n1455_n3628.n139 a_n1455_n3628.n138 185
R16719 a_n1455_n3628.n123 a_n1455_n3628.n122 185
R16720 a_n1455_n3628.n135 a_n1455_n3628.n134 185
R16721 a_n1455_n3628.n133 a_n1455_n3628.n132 185
R16722 a_n1455_n3628.n126 a_n1455_n3628.n125 185
R16723 a_n1455_n3628.n129 a_n1455_n3628.n128 185
R16724 a_n1455_n3628.n87 a_n1455_n3628.n86 185
R16725 a_n1455_n3628.n85 a_n1455_n3628.n84 185
R16726 a_n1455_n3628.n69 a_n1455_n3628.n68 185
R16727 a_n1455_n3628.n81 a_n1455_n3628.n80 185
R16728 a_n1455_n3628.n79 a_n1455_n3628.n78 185
R16729 a_n1455_n3628.n72 a_n1455_n3628.n71 185
R16730 a_n1455_n3628.n75 a_n1455_n3628.n74 185
R16731 a_n1455_n3628.n192 a_n1455_n3628.n191 185
R16732 a_n1455_n3628.n190 a_n1455_n3628.n189 185
R16733 a_n1455_n3628.n174 a_n1455_n3628.n173 185
R16734 a_n1455_n3628.n186 a_n1455_n3628.n185 185
R16735 a_n1455_n3628.n184 a_n1455_n3628.n183 185
R16736 a_n1455_n3628.n177 a_n1455_n3628.n176 185
R16737 a_n1455_n3628.n180 a_n1455_n3628.n179 185
R16738 a_n1455_n3628.n218 a_n1455_n3628.n217 185
R16739 a_n1455_n3628.n216 a_n1455_n3628.n215 185
R16740 a_n1455_n3628.n200 a_n1455_n3628.n199 185
R16741 a_n1455_n3628.n212 a_n1455_n3628.n211 185
R16742 a_n1455_n3628.n210 a_n1455_n3628.n209 185
R16743 a_n1455_n3628.n203 a_n1455_n3628.n202 185
R16744 a_n1455_n3628.n206 a_n1455_n3628.n205 185
R16745 a_n1455_n3628.n167 a_n1455_n3628.n166 185
R16746 a_n1455_n3628.n165 a_n1455_n3628.n164 185
R16747 a_n1455_n3628.n149 a_n1455_n3628.n148 185
R16748 a_n1455_n3628.n161 a_n1455_n3628.n160 185
R16749 a_n1455_n3628.n159 a_n1455_n3628.n158 185
R16750 a_n1455_n3628.n152 a_n1455_n3628.n151 185
R16751 a_n1455_n3628.n155 a_n1455_n3628.n154 185
R16752 a_n1455_n3628.n313 a_n1455_n3628.n312 185
R16753 a_n1455_n3628.n310 a_n1455_n3628.n309 185
R16754 a_n1455_n3628.n317 a_n1455_n3628.n316 185
R16755 a_n1455_n3628.n319 a_n1455_n3628.n318 185
R16756 a_n1455_n3628.n307 a_n1455_n3628.n306 185
R16757 a_n1455_n3628.n323 a_n1455_n3628.n322 185
R16758 a_n1455_n3628.n325 a_n1455_n3628.n324 185
R16759 a_n1455_n3628.n286 a_n1455_n3628.n285 185
R16760 a_n1455_n3628.n283 a_n1455_n3628.n282 185
R16761 a_n1455_n3628.n290 a_n1455_n3628.n289 185
R16762 a_n1455_n3628.n292 a_n1455_n3628.n291 185
R16763 a_n1455_n3628.n280 a_n1455_n3628.n279 185
R16764 a_n1455_n3628.n296 a_n1455_n3628.n295 185
R16765 a_n1455_n3628.n298 a_n1455_n3628.n297 185
R16766 a_n1455_n3628.n261 a_n1455_n3628.n260 185
R16767 a_n1455_n3628.n258 a_n1455_n3628.n257 185
R16768 a_n1455_n3628.n265 a_n1455_n3628.n264 185
R16769 a_n1455_n3628.n267 a_n1455_n3628.n266 185
R16770 a_n1455_n3628.n255 a_n1455_n3628.n254 185
R16771 a_n1455_n3628.n271 a_n1455_n3628.n270 185
R16772 a_n1455_n3628.n273 a_n1455_n3628.n272 185
R16773 a_n1455_n3628.n234 a_n1455_n3628.n233 185
R16774 a_n1455_n3628.n231 a_n1455_n3628.n230 185
R16775 a_n1455_n3628.n238 a_n1455_n3628.n237 185
R16776 a_n1455_n3628.n240 a_n1455_n3628.n239 185
R16777 a_n1455_n3628.n228 a_n1455_n3628.n227 185
R16778 a_n1455_n3628.n244 a_n1455_n3628.n243 185
R16779 a_n1455_n3628.n246 a_n1455_n3628.n245 185
R16780 a_n1455_n3628.t14 a_n1455_n3628.n337 147.661
R16781 a_n1455_n3628.t17 a_n1455_n3628.n47 147.661
R16782 a_n1455_n3628.t6 a_n1455_n3628.n99 147.661
R16783 a_n1455_n3628.t9 a_n1455_n3628.n127 147.661
R16784 a_n1455_n3628.t8 a_n1455_n3628.n73 147.661
R16785 a_n1455_n3628.t5 a_n1455_n3628.n178 147.661
R16786 a_n1455_n3628.t7 a_n1455_n3628.n204 147.661
R16787 a_n1455_n3628.t0 a_n1455_n3628.n153 147.661
R16788 a_n1455_n3628.t4 a_n1455_n3628.n311 147.661
R16789 a_n1455_n3628.t1 a_n1455_n3628.n284 147.661
R16790 a_n1455_n3628.t19 a_n1455_n3628.n259 147.661
R16791 a_n1455_n3628.t15 a_n1455_n3628.n232 147.661
R16792 a_n1455_n3628.n350 a_n1455_n3628.n349 104.615
R16793 a_n1455_n3628.n349 a_n1455_n3628.n332 104.615
R16794 a_n1455_n3628.n344 a_n1455_n3628.n332 104.615
R16795 a_n1455_n3628.n344 a_n1455_n3628.n343 104.615
R16796 a_n1455_n3628.n343 a_n1455_n3628.n335 104.615
R16797 a_n1455_n3628.n338 a_n1455_n3628.n335 104.615
R16798 a_n1455_n3628.n60 a_n1455_n3628.n59 104.615
R16799 a_n1455_n3628.n59 a_n1455_n3628.n42 104.615
R16800 a_n1455_n3628.n54 a_n1455_n3628.n42 104.615
R16801 a_n1455_n3628.n54 a_n1455_n3628.n53 104.615
R16802 a_n1455_n3628.n53 a_n1455_n3628.n45 104.615
R16803 a_n1455_n3628.n48 a_n1455_n3628.n45 104.615
R16804 a_n1455_n3628.n112 a_n1455_n3628.n111 104.615
R16805 a_n1455_n3628.n111 a_n1455_n3628.n94 104.615
R16806 a_n1455_n3628.n106 a_n1455_n3628.n94 104.615
R16807 a_n1455_n3628.n106 a_n1455_n3628.n105 104.615
R16808 a_n1455_n3628.n105 a_n1455_n3628.n97 104.615
R16809 a_n1455_n3628.n100 a_n1455_n3628.n97 104.615
R16810 a_n1455_n3628.n140 a_n1455_n3628.n139 104.615
R16811 a_n1455_n3628.n139 a_n1455_n3628.n122 104.615
R16812 a_n1455_n3628.n134 a_n1455_n3628.n122 104.615
R16813 a_n1455_n3628.n134 a_n1455_n3628.n133 104.615
R16814 a_n1455_n3628.n133 a_n1455_n3628.n125 104.615
R16815 a_n1455_n3628.n128 a_n1455_n3628.n125 104.615
R16816 a_n1455_n3628.n86 a_n1455_n3628.n85 104.615
R16817 a_n1455_n3628.n85 a_n1455_n3628.n68 104.615
R16818 a_n1455_n3628.n80 a_n1455_n3628.n68 104.615
R16819 a_n1455_n3628.n80 a_n1455_n3628.n79 104.615
R16820 a_n1455_n3628.n79 a_n1455_n3628.n71 104.615
R16821 a_n1455_n3628.n74 a_n1455_n3628.n71 104.615
R16822 a_n1455_n3628.n191 a_n1455_n3628.n190 104.615
R16823 a_n1455_n3628.n190 a_n1455_n3628.n173 104.615
R16824 a_n1455_n3628.n185 a_n1455_n3628.n173 104.615
R16825 a_n1455_n3628.n185 a_n1455_n3628.n184 104.615
R16826 a_n1455_n3628.n184 a_n1455_n3628.n176 104.615
R16827 a_n1455_n3628.n179 a_n1455_n3628.n176 104.615
R16828 a_n1455_n3628.n217 a_n1455_n3628.n216 104.615
R16829 a_n1455_n3628.n216 a_n1455_n3628.n199 104.615
R16830 a_n1455_n3628.n211 a_n1455_n3628.n199 104.615
R16831 a_n1455_n3628.n211 a_n1455_n3628.n210 104.615
R16832 a_n1455_n3628.n210 a_n1455_n3628.n202 104.615
R16833 a_n1455_n3628.n205 a_n1455_n3628.n202 104.615
R16834 a_n1455_n3628.n166 a_n1455_n3628.n165 104.615
R16835 a_n1455_n3628.n165 a_n1455_n3628.n148 104.615
R16836 a_n1455_n3628.n160 a_n1455_n3628.n148 104.615
R16837 a_n1455_n3628.n160 a_n1455_n3628.n159 104.615
R16838 a_n1455_n3628.n159 a_n1455_n3628.n151 104.615
R16839 a_n1455_n3628.n154 a_n1455_n3628.n151 104.615
R16840 a_n1455_n3628.n312 a_n1455_n3628.n309 104.615
R16841 a_n1455_n3628.n317 a_n1455_n3628.n309 104.615
R16842 a_n1455_n3628.n318 a_n1455_n3628.n317 104.615
R16843 a_n1455_n3628.n318 a_n1455_n3628.n306 104.615
R16844 a_n1455_n3628.n323 a_n1455_n3628.n306 104.615
R16845 a_n1455_n3628.n324 a_n1455_n3628.n323 104.615
R16846 a_n1455_n3628.n285 a_n1455_n3628.n282 104.615
R16847 a_n1455_n3628.n290 a_n1455_n3628.n282 104.615
R16848 a_n1455_n3628.n291 a_n1455_n3628.n290 104.615
R16849 a_n1455_n3628.n291 a_n1455_n3628.n279 104.615
R16850 a_n1455_n3628.n296 a_n1455_n3628.n279 104.615
R16851 a_n1455_n3628.n297 a_n1455_n3628.n296 104.615
R16852 a_n1455_n3628.n260 a_n1455_n3628.n257 104.615
R16853 a_n1455_n3628.n265 a_n1455_n3628.n257 104.615
R16854 a_n1455_n3628.n266 a_n1455_n3628.n265 104.615
R16855 a_n1455_n3628.n266 a_n1455_n3628.n254 104.615
R16856 a_n1455_n3628.n271 a_n1455_n3628.n254 104.615
R16857 a_n1455_n3628.n272 a_n1455_n3628.n271 104.615
R16858 a_n1455_n3628.n233 a_n1455_n3628.n230 104.615
R16859 a_n1455_n3628.n238 a_n1455_n3628.n230 104.615
R16860 a_n1455_n3628.n239 a_n1455_n3628.n238 104.615
R16861 a_n1455_n3628.n239 a_n1455_n3628.n227 104.615
R16862 a_n1455_n3628.n244 a_n1455_n3628.n227 104.615
R16863 a_n1455_n3628.n245 a_n1455_n3628.n244 104.615
R16864 a_n1455_n3628.n119 a_n1455_n3628.n118 56.1363
R16865 a_n1455_n3628.n357 a_n1455_n3628.n356 56.1363
R16866 a_n1455_n3628.n303 a_n1455_n3628.n302 56.1361
R16867 a_n1455_n3628.n251 a_n1455_n3628.n250 56.1361
R16868 a_n1455_n3628.n338 a_n1455_n3628.t14 52.3082
R16869 a_n1455_n3628.n48 a_n1455_n3628.t17 52.3082
R16870 a_n1455_n3628.n100 a_n1455_n3628.t6 52.3082
R16871 a_n1455_n3628.n128 a_n1455_n3628.t9 52.3082
R16872 a_n1455_n3628.n74 a_n1455_n3628.t8 52.3082
R16873 a_n1455_n3628.n179 a_n1455_n3628.t5 52.3082
R16874 a_n1455_n3628.n205 a_n1455_n3628.t7 52.3082
R16875 a_n1455_n3628.n154 a_n1455_n3628.t0 52.3082
R16876 a_n1455_n3628.n312 a_n1455_n3628.t4 52.3082
R16877 a_n1455_n3628.n285 a_n1455_n3628.t1 52.3082
R16878 a_n1455_n3628.n260 a_n1455_n3628.t19 52.3082
R16879 a_n1455_n3628.n233 a_n1455_n3628.t15 52.3082
R16880 a_n1455_n3628.n355 a_n1455_n3628.n354 37.8096
R16881 a_n1455_n3628.n65 a_n1455_n3628.n64 37.8096
R16882 a_n1455_n3628.n117 a_n1455_n3628.n116 37.8096
R16883 a_n1455_n3628.n145 a_n1455_n3628.n144 37.8096
R16884 a_n1455_n3628.n328 a_n1455_n3628.n327 37.8096
R16885 a_n1455_n3628.n301 a_n1455_n3628.n300 37.8096
R16886 a_n1455_n3628.n276 a_n1455_n3628.n275 37.8096
R16887 a_n1455_n3628.n249 a_n1455_n3628.n248 37.8096
R16888 a_n1455_n3628.n339 a_n1455_n3628.n337 15.6674
R16889 a_n1455_n3628.n49 a_n1455_n3628.n47 15.6674
R16890 a_n1455_n3628.n101 a_n1455_n3628.n99 15.6674
R16891 a_n1455_n3628.n129 a_n1455_n3628.n127 15.6674
R16892 a_n1455_n3628.n75 a_n1455_n3628.n73 15.6674
R16893 a_n1455_n3628.n180 a_n1455_n3628.n178 15.6674
R16894 a_n1455_n3628.n206 a_n1455_n3628.n204 15.6674
R16895 a_n1455_n3628.n155 a_n1455_n3628.n153 15.6674
R16896 a_n1455_n3628.n313 a_n1455_n3628.n311 15.6674
R16897 a_n1455_n3628.n286 a_n1455_n3628.n284 15.6674
R16898 a_n1455_n3628.n261 a_n1455_n3628.n259 15.6674
R16899 a_n1455_n3628.n234 a_n1455_n3628.n232 15.6674
R16900 a_n1455_n3628.n340 a_n1455_n3628.n336 12.8005
R16901 a_n1455_n3628.n50 a_n1455_n3628.n46 12.8005
R16902 a_n1455_n3628.n102 a_n1455_n3628.n98 12.8005
R16903 a_n1455_n3628.n130 a_n1455_n3628.n126 12.8005
R16904 a_n1455_n3628.n76 a_n1455_n3628.n72 12.8005
R16905 a_n1455_n3628.n181 a_n1455_n3628.n177 12.8005
R16906 a_n1455_n3628.n207 a_n1455_n3628.n203 12.8005
R16907 a_n1455_n3628.n156 a_n1455_n3628.n152 12.8005
R16908 a_n1455_n3628.n314 a_n1455_n3628.n310 12.8005
R16909 a_n1455_n3628.n287 a_n1455_n3628.n283 12.8005
R16910 a_n1455_n3628.n262 a_n1455_n3628.n258 12.8005
R16911 a_n1455_n3628.n235 a_n1455_n3628.n231 12.8005
R16912 a_n1455_n3628.n342 a_n1455_n3628.n341 12.0247
R16913 a_n1455_n3628.n52 a_n1455_n3628.n51 12.0247
R16914 a_n1455_n3628.n104 a_n1455_n3628.n103 12.0247
R16915 a_n1455_n3628.n132 a_n1455_n3628.n131 12.0247
R16916 a_n1455_n3628.n78 a_n1455_n3628.n77 12.0247
R16917 a_n1455_n3628.n183 a_n1455_n3628.n182 12.0247
R16918 a_n1455_n3628.n209 a_n1455_n3628.n208 12.0247
R16919 a_n1455_n3628.n158 a_n1455_n3628.n157 12.0247
R16920 a_n1455_n3628.n316 a_n1455_n3628.n315 12.0247
R16921 a_n1455_n3628.n289 a_n1455_n3628.n288 12.0247
R16922 a_n1455_n3628.n264 a_n1455_n3628.n263 12.0247
R16923 a_n1455_n3628.n237 a_n1455_n3628.n236 12.0247
R16924 a_n1455_n3628.n224 a_n1455_n3628.n145 11.5057
R16925 a_n1455_n3628.n355 a_n1455_n3628.n329 11.5057
R16926 a_n1455_n3628.n345 a_n1455_n3628.n334 11.249
R16927 a_n1455_n3628.n55 a_n1455_n3628.n44 11.249
R16928 a_n1455_n3628.n107 a_n1455_n3628.n96 11.249
R16929 a_n1455_n3628.n135 a_n1455_n3628.n124 11.249
R16930 a_n1455_n3628.n81 a_n1455_n3628.n70 11.249
R16931 a_n1455_n3628.n186 a_n1455_n3628.n175 11.249
R16932 a_n1455_n3628.n212 a_n1455_n3628.n201 11.249
R16933 a_n1455_n3628.n161 a_n1455_n3628.n150 11.249
R16934 a_n1455_n3628.n319 a_n1455_n3628.n308 11.249
R16935 a_n1455_n3628.n292 a_n1455_n3628.n281 11.249
R16936 a_n1455_n3628.n267 a_n1455_n3628.n256 11.249
R16937 a_n1455_n3628.n240 a_n1455_n3628.n229 11.249
R16938 a_n1455_n3628.n346 a_n1455_n3628.n333 10.4732
R16939 a_n1455_n3628.n56 a_n1455_n3628.n43 10.4732
R16940 a_n1455_n3628.n108 a_n1455_n3628.n95 10.4732
R16941 a_n1455_n3628.n136 a_n1455_n3628.n123 10.4732
R16942 a_n1455_n3628.n82 a_n1455_n3628.n69 10.4732
R16943 a_n1455_n3628.n187 a_n1455_n3628.n174 10.4732
R16944 a_n1455_n3628.n213 a_n1455_n3628.n200 10.4732
R16945 a_n1455_n3628.n162 a_n1455_n3628.n149 10.4732
R16946 a_n1455_n3628.n320 a_n1455_n3628.n307 10.4732
R16947 a_n1455_n3628.n293 a_n1455_n3628.n280 10.4732
R16948 a_n1455_n3628.n268 a_n1455_n3628.n255 10.4732
R16949 a_n1455_n3628.n241 a_n1455_n3628.n228 10.4732
R16950 a_n1455_n3628.n348 a_n1455_n3628.n347 9.69747
R16951 a_n1455_n3628.n58 a_n1455_n3628.n57 9.69747
R16952 a_n1455_n3628.n110 a_n1455_n3628.n109 9.69747
R16953 a_n1455_n3628.n138 a_n1455_n3628.n137 9.69747
R16954 a_n1455_n3628.n84 a_n1455_n3628.n83 9.69747
R16955 a_n1455_n3628.n189 a_n1455_n3628.n188 9.69747
R16956 a_n1455_n3628.n215 a_n1455_n3628.n214 9.69747
R16957 a_n1455_n3628.n164 a_n1455_n3628.n163 9.69747
R16958 a_n1455_n3628.n322 a_n1455_n3628.n321 9.69747
R16959 a_n1455_n3628.n295 a_n1455_n3628.n294 9.69747
R16960 a_n1455_n3628.n270 a_n1455_n3628.n269 9.69747
R16961 a_n1455_n3628.n243 a_n1455_n3628.n242 9.69747
R16962 a_n1455_n3628.n354 a_n1455_n3628.n353 9.45567
R16963 a_n1455_n3628.n64 a_n1455_n3628.n63 9.45567
R16964 a_n1455_n3628.n116 a_n1455_n3628.n115 9.45567
R16965 a_n1455_n3628.n144 a_n1455_n3628.n143 9.45567
R16966 a_n1455_n3628.n90 a_n1455_n3628.n89 9.45567
R16967 a_n1455_n3628.n195 a_n1455_n3628.n194 9.45567
R16968 a_n1455_n3628.n221 a_n1455_n3628.n220 9.45567
R16969 a_n1455_n3628.n170 a_n1455_n3628.n169 9.45567
R16970 a_n1455_n3628.n327 a_n1455_n3628.n26 9.45567
R16971 a_n1455_n3628.n300 a_n1455_n3628.n30 9.45567
R16972 a_n1455_n3628.n275 a_n1455_n3628.n34 9.45567
R16973 a_n1455_n3628.n248 a_n1455_n3628.n38 9.45567
R16974 a_n1455_n3628.n353 a_n1455_n3628.n352 9.3005
R16975 a_n1455_n3628.n331 a_n1455_n3628.n1 9.3005
R16976 a_n1455_n3628.n347 a_n1455_n3628.n1 9.3005
R16977 a_n1455_n3628.n0 a_n1455_n3628.n346 9.3005
R16978 a_n1455_n3628.n334 a_n1455_n3628.n0 9.3005
R16979 a_n1455_n3628.n341 a_n1455_n3628.n2 9.3005
R16980 a_n1455_n3628.n2 a_n1455_n3628.n340 9.3005
R16981 a_n1455_n3628.n63 a_n1455_n3628.n62 9.3005
R16982 a_n1455_n3628.n41 a_n1455_n3628.n4 9.3005
R16983 a_n1455_n3628.n57 a_n1455_n3628.n4 9.3005
R16984 a_n1455_n3628.n3 a_n1455_n3628.n56 9.3005
R16985 a_n1455_n3628.n44 a_n1455_n3628.n3 9.3005
R16986 a_n1455_n3628.n51 a_n1455_n3628.n5 9.3005
R16987 a_n1455_n3628.n5 a_n1455_n3628.n50 9.3005
R16988 a_n1455_n3628.n115 a_n1455_n3628.n114 9.3005
R16989 a_n1455_n3628.n93 a_n1455_n3628.n7 9.3005
R16990 a_n1455_n3628.n109 a_n1455_n3628.n7 9.3005
R16991 a_n1455_n3628.n6 a_n1455_n3628.n108 9.3005
R16992 a_n1455_n3628.n96 a_n1455_n3628.n6 9.3005
R16993 a_n1455_n3628.n103 a_n1455_n3628.n8 9.3005
R16994 a_n1455_n3628.n8 a_n1455_n3628.n102 9.3005
R16995 a_n1455_n3628.n143 a_n1455_n3628.n142 9.3005
R16996 a_n1455_n3628.n121 a_n1455_n3628.n10 9.3005
R16997 a_n1455_n3628.n137 a_n1455_n3628.n10 9.3005
R16998 a_n1455_n3628.n9 a_n1455_n3628.n136 9.3005
R16999 a_n1455_n3628.n124 a_n1455_n3628.n9 9.3005
R17000 a_n1455_n3628.n131 a_n1455_n3628.n11 9.3005
R17001 a_n1455_n3628.n11 a_n1455_n3628.n130 9.3005
R17002 a_n1455_n3628.n89 a_n1455_n3628.n88 9.3005
R17003 a_n1455_n3628.n67 a_n1455_n3628.n13 9.3005
R17004 a_n1455_n3628.n83 a_n1455_n3628.n13 9.3005
R17005 a_n1455_n3628.n12 a_n1455_n3628.n82 9.3005
R17006 a_n1455_n3628.n70 a_n1455_n3628.n12 9.3005
R17007 a_n1455_n3628.n77 a_n1455_n3628.n14 9.3005
R17008 a_n1455_n3628.n14 a_n1455_n3628.n76 9.3005
R17009 a_n1455_n3628.n194 a_n1455_n3628.n193 9.3005
R17010 a_n1455_n3628.n172 a_n1455_n3628.n16 9.3005
R17011 a_n1455_n3628.n188 a_n1455_n3628.n16 9.3005
R17012 a_n1455_n3628.n15 a_n1455_n3628.n187 9.3005
R17013 a_n1455_n3628.n175 a_n1455_n3628.n15 9.3005
R17014 a_n1455_n3628.n182 a_n1455_n3628.n17 9.3005
R17015 a_n1455_n3628.n17 a_n1455_n3628.n181 9.3005
R17016 a_n1455_n3628.n220 a_n1455_n3628.n219 9.3005
R17017 a_n1455_n3628.n198 a_n1455_n3628.n19 9.3005
R17018 a_n1455_n3628.n214 a_n1455_n3628.n19 9.3005
R17019 a_n1455_n3628.n18 a_n1455_n3628.n213 9.3005
R17020 a_n1455_n3628.n201 a_n1455_n3628.n18 9.3005
R17021 a_n1455_n3628.n208 a_n1455_n3628.n20 9.3005
R17022 a_n1455_n3628.n20 a_n1455_n3628.n207 9.3005
R17023 a_n1455_n3628.n169 a_n1455_n3628.n168 9.3005
R17024 a_n1455_n3628.n147 a_n1455_n3628.n22 9.3005
R17025 a_n1455_n3628.n163 a_n1455_n3628.n22 9.3005
R17026 a_n1455_n3628.n21 a_n1455_n3628.n162 9.3005
R17027 a_n1455_n3628.n150 a_n1455_n3628.n21 9.3005
R17028 a_n1455_n3628.n157 a_n1455_n3628.n23 9.3005
R17029 a_n1455_n3628.n23 a_n1455_n3628.n156 9.3005
R17030 a_n1455_n3628.n26 a_n1455_n3628.n326 9.3005
R17031 a_n1455_n3628.n305 a_n1455_n3628.n26 9.3005
R17032 a_n1455_n3628.n321 a_n1455_n3628.n27 9.3005
R17033 a_n1455_n3628.n27 a_n1455_n3628.n320 9.3005
R17034 a_n1455_n3628.n308 a_n1455_n3628.n25 9.3005
R17035 a_n1455_n3628.n315 a_n1455_n3628.n25 9.3005
R17036 a_n1455_n3628.n24 a_n1455_n3628.n314 9.3005
R17037 a_n1455_n3628.n30 a_n1455_n3628.n299 9.3005
R17038 a_n1455_n3628.n278 a_n1455_n3628.n30 9.3005
R17039 a_n1455_n3628.n294 a_n1455_n3628.n31 9.3005
R17040 a_n1455_n3628.n31 a_n1455_n3628.n293 9.3005
R17041 a_n1455_n3628.n281 a_n1455_n3628.n29 9.3005
R17042 a_n1455_n3628.n288 a_n1455_n3628.n29 9.3005
R17043 a_n1455_n3628.n28 a_n1455_n3628.n287 9.3005
R17044 a_n1455_n3628.n34 a_n1455_n3628.n274 9.3005
R17045 a_n1455_n3628.n253 a_n1455_n3628.n34 9.3005
R17046 a_n1455_n3628.n269 a_n1455_n3628.n35 9.3005
R17047 a_n1455_n3628.n35 a_n1455_n3628.n268 9.3005
R17048 a_n1455_n3628.n256 a_n1455_n3628.n33 9.3005
R17049 a_n1455_n3628.n263 a_n1455_n3628.n33 9.3005
R17050 a_n1455_n3628.n32 a_n1455_n3628.n262 9.3005
R17051 a_n1455_n3628.n38 a_n1455_n3628.n247 9.3005
R17052 a_n1455_n3628.n226 a_n1455_n3628.n38 9.3005
R17053 a_n1455_n3628.n242 a_n1455_n3628.n39 9.3005
R17054 a_n1455_n3628.n39 a_n1455_n3628.n241 9.3005
R17055 a_n1455_n3628.n229 a_n1455_n3628.n37 9.3005
R17056 a_n1455_n3628.n236 a_n1455_n3628.n37 9.3005
R17057 a_n1455_n3628.n36 a_n1455_n3628.n235 9.3005
R17058 a_n1455_n3628.n351 a_n1455_n3628.n331 8.92171
R17059 a_n1455_n3628.n61 a_n1455_n3628.n41 8.92171
R17060 a_n1455_n3628.n113 a_n1455_n3628.n93 8.92171
R17061 a_n1455_n3628.n141 a_n1455_n3628.n121 8.92171
R17062 a_n1455_n3628.n87 a_n1455_n3628.n67 8.92171
R17063 a_n1455_n3628.n192 a_n1455_n3628.n172 8.92171
R17064 a_n1455_n3628.n218 a_n1455_n3628.n198 8.92171
R17065 a_n1455_n3628.n167 a_n1455_n3628.n147 8.92171
R17066 a_n1455_n3628.n325 a_n1455_n3628.n305 8.92171
R17067 a_n1455_n3628.n298 a_n1455_n3628.n278 8.92171
R17068 a_n1455_n3628.n273 a_n1455_n3628.n253 8.92171
R17069 a_n1455_n3628.n246 a_n1455_n3628.n226 8.92171
R17070 a_n1455_n3628.n352 a_n1455_n3628.n330 8.14595
R17071 a_n1455_n3628.n62 a_n1455_n3628.n40 8.14595
R17072 a_n1455_n3628.n114 a_n1455_n3628.n92 8.14595
R17073 a_n1455_n3628.n142 a_n1455_n3628.n120 8.14595
R17074 a_n1455_n3628.n88 a_n1455_n3628.n66 8.14595
R17075 a_n1455_n3628.n193 a_n1455_n3628.n171 8.14595
R17076 a_n1455_n3628.n219 a_n1455_n3628.n197 8.14595
R17077 a_n1455_n3628.n168 a_n1455_n3628.n146 8.14595
R17078 a_n1455_n3628.n326 a_n1455_n3628.n304 8.14595
R17079 a_n1455_n3628.n299 a_n1455_n3628.n277 8.14595
R17080 a_n1455_n3628.n274 a_n1455_n3628.n252 8.14595
R17081 a_n1455_n3628.n247 a_n1455_n3628.n225 8.14595
R17082 a_n1455_n3628.n354 a_n1455_n3628.n330 5.81868
R17083 a_n1455_n3628.n64 a_n1455_n3628.n40 5.81868
R17084 a_n1455_n3628.n116 a_n1455_n3628.n92 5.81868
R17085 a_n1455_n3628.n144 a_n1455_n3628.n120 5.81868
R17086 a_n1455_n3628.n90 a_n1455_n3628.n66 5.81868
R17087 a_n1455_n3628.n195 a_n1455_n3628.n171 5.81868
R17088 a_n1455_n3628.n221 a_n1455_n3628.n197 5.81868
R17089 a_n1455_n3628.n170 a_n1455_n3628.n146 5.81868
R17090 a_n1455_n3628.n327 a_n1455_n3628.n304 5.81868
R17091 a_n1455_n3628.n300 a_n1455_n3628.n277 5.81868
R17092 a_n1455_n3628.n275 a_n1455_n3628.n252 5.81868
R17093 a_n1455_n3628.n248 a_n1455_n3628.n225 5.81868
R17094 a_n1455_n3628.n249 a_n1455_n3628.n224 5.18369
R17095 a_n1455_n3628.n329 a_n1455_n3628.n328 5.18369
R17096 a_n1455_n3628.n352 a_n1455_n3628.n351 5.04292
R17097 a_n1455_n3628.n62 a_n1455_n3628.n61 5.04292
R17098 a_n1455_n3628.n114 a_n1455_n3628.n113 5.04292
R17099 a_n1455_n3628.n142 a_n1455_n3628.n141 5.04292
R17100 a_n1455_n3628.n88 a_n1455_n3628.n87 5.04292
R17101 a_n1455_n3628.n193 a_n1455_n3628.n192 5.04292
R17102 a_n1455_n3628.n219 a_n1455_n3628.n218 5.04292
R17103 a_n1455_n3628.n168 a_n1455_n3628.n167 5.04292
R17104 a_n1455_n3628.n326 a_n1455_n3628.n325 5.04292
R17105 a_n1455_n3628.n299 a_n1455_n3628.n298 5.04292
R17106 a_n1455_n3628.n274 a_n1455_n3628.n273 5.04292
R17107 a_n1455_n3628.n247 a_n1455_n3628.n246 5.04292
R17108 a_n1455_n3628.n2 a_n1455_n3628.n337 4.38594
R17109 a_n1455_n3628.n5 a_n1455_n3628.n47 4.38594
R17110 a_n1455_n3628.n8 a_n1455_n3628.n99 4.38594
R17111 a_n1455_n3628.n11 a_n1455_n3628.n127 4.38594
R17112 a_n1455_n3628.n14 a_n1455_n3628.n73 4.38594
R17113 a_n1455_n3628.n17 a_n1455_n3628.n178 4.38594
R17114 a_n1455_n3628.n20 a_n1455_n3628.n204 4.38594
R17115 a_n1455_n3628.n23 a_n1455_n3628.n153 4.38594
R17116 a_n1455_n3628.n24 a_n1455_n3628.n311 4.38594
R17117 a_n1455_n3628.n28 a_n1455_n3628.n284 4.38594
R17118 a_n1455_n3628.n32 a_n1455_n3628.n259 4.38594
R17119 a_n1455_n3628.n36 a_n1455_n3628.n232 4.38594
R17120 a_n1455_n3628.n348 a_n1455_n3628.n331 4.26717
R17121 a_n1455_n3628.n58 a_n1455_n3628.n41 4.26717
R17122 a_n1455_n3628.n110 a_n1455_n3628.n93 4.26717
R17123 a_n1455_n3628.n138 a_n1455_n3628.n121 4.26717
R17124 a_n1455_n3628.n84 a_n1455_n3628.n67 4.26717
R17125 a_n1455_n3628.n189 a_n1455_n3628.n172 4.26717
R17126 a_n1455_n3628.n215 a_n1455_n3628.n198 4.26717
R17127 a_n1455_n3628.n164 a_n1455_n3628.n147 4.26717
R17128 a_n1455_n3628.n322 a_n1455_n3628.n305 4.26717
R17129 a_n1455_n3628.n295 a_n1455_n3628.n278 4.26717
R17130 a_n1455_n3628.n270 a_n1455_n3628.n253 4.26717
R17131 a_n1455_n3628.n243 a_n1455_n3628.n226 4.26717
R17132 a_n1455_n3628.n347 a_n1455_n3628.n333 3.49141
R17133 a_n1455_n3628.n57 a_n1455_n3628.n43 3.49141
R17134 a_n1455_n3628.n109 a_n1455_n3628.n95 3.49141
R17135 a_n1455_n3628.n137 a_n1455_n3628.n123 3.49141
R17136 a_n1455_n3628.n83 a_n1455_n3628.n69 3.49141
R17137 a_n1455_n3628.n188 a_n1455_n3628.n174 3.49141
R17138 a_n1455_n3628.n214 a_n1455_n3628.n200 3.49141
R17139 a_n1455_n3628.n163 a_n1455_n3628.n149 3.49141
R17140 a_n1455_n3628.n321 a_n1455_n3628.n307 3.49141
R17141 a_n1455_n3628.n294 a_n1455_n3628.n280 3.49141
R17142 a_n1455_n3628.n269 a_n1455_n3628.n255 3.49141
R17143 a_n1455_n3628.n242 a_n1455_n3628.n228 3.49141
R17144 a_n1455_n3628.n118 a_n1455_n3628.t10 3.3005
R17145 a_n1455_n3628.n118 a_n1455_n3628.t2 3.3005
R17146 a_n1455_n3628.n302 a_n1455_n3628.t11 3.3005
R17147 a_n1455_n3628.n302 a_n1455_n3628.t3 3.3005
R17148 a_n1455_n3628.n250 a_n1455_n3628.t16 3.3005
R17149 a_n1455_n3628.n250 a_n1455_n3628.t12 3.3005
R17150 a_n1455_n3628.t18 a_n1455_n3628.n357 3.3005
R17151 a_n1455_n3628.n357 a_n1455_n3628.t13 3.3005
R17152 a_n1455_n3628.n346 a_n1455_n3628.n345 2.71565
R17153 a_n1455_n3628.n56 a_n1455_n3628.n55 2.71565
R17154 a_n1455_n3628.n108 a_n1455_n3628.n107 2.71565
R17155 a_n1455_n3628.n136 a_n1455_n3628.n135 2.71565
R17156 a_n1455_n3628.n82 a_n1455_n3628.n81 2.71565
R17157 a_n1455_n3628.n187 a_n1455_n3628.n186 2.71565
R17158 a_n1455_n3628.n213 a_n1455_n3628.n212 2.71565
R17159 a_n1455_n3628.n162 a_n1455_n3628.n161 2.71565
R17160 a_n1455_n3628.n320 a_n1455_n3628.n319 2.71565
R17161 a_n1455_n3628.n293 a_n1455_n3628.n292 2.71565
R17162 a_n1455_n3628.n268 a_n1455_n3628.n267 2.71565
R17163 a_n1455_n3628.n241 a_n1455_n3628.n240 2.71565
R17164 a_n1455_n3628.n329 a_n1455_n3628.n91 2.23674
R17165 a_n1455_n3628.n224 a_n1455_n3628.n223 1.95694
R17166 a_n1455_n3628.n342 a_n1455_n3628.n334 1.93989
R17167 a_n1455_n3628.n52 a_n1455_n3628.n44 1.93989
R17168 a_n1455_n3628.n104 a_n1455_n3628.n96 1.93989
R17169 a_n1455_n3628.n132 a_n1455_n3628.n124 1.93989
R17170 a_n1455_n3628.n78 a_n1455_n3628.n70 1.93989
R17171 a_n1455_n3628.n183 a_n1455_n3628.n175 1.93989
R17172 a_n1455_n3628.n209 a_n1455_n3628.n201 1.93989
R17173 a_n1455_n3628.n158 a_n1455_n3628.n150 1.93989
R17174 a_n1455_n3628.n316 a_n1455_n3628.n308 1.93989
R17175 a_n1455_n3628.n289 a_n1455_n3628.n281 1.93989
R17176 a_n1455_n3628.n264 a_n1455_n3628.n256 1.93989
R17177 a_n1455_n3628.n237 a_n1455_n3628.n229 1.93989
R17178 a_n1455_n3628.n341 a_n1455_n3628.n336 1.16414
R17179 a_n1455_n3628.n51 a_n1455_n3628.n46 1.16414
R17180 a_n1455_n3628.n103 a_n1455_n3628.n98 1.16414
R17181 a_n1455_n3628.n131 a_n1455_n3628.n126 1.16414
R17182 a_n1455_n3628.n77 a_n1455_n3628.n72 1.16414
R17183 a_n1455_n3628.n182 a_n1455_n3628.n177 1.16414
R17184 a_n1455_n3628.n208 a_n1455_n3628.n203 1.16414
R17185 a_n1455_n3628.n157 a_n1455_n3628.n152 1.16414
R17186 a_n1455_n3628.n315 a_n1455_n3628.n310 1.16414
R17187 a_n1455_n3628.n288 a_n1455_n3628.n283 1.16414
R17188 a_n1455_n3628.n263 a_n1455_n3628.n258 1.16414
R17189 a_n1455_n3628.n236 a_n1455_n3628.n231 1.16414
R17190 a_n1455_n3628.n222 a_n1455_n3628.n196 0.962709
R17191 a_n1455_n3628.n196 a_n1455_n3628.n91 0.962709
R17192 a_n1455_n3628.n251 a_n1455_n3628.n249 0.573776
R17193 a_n1455_n3628.n276 a_n1455_n3628.n251 0.573776
R17194 a_n1455_n3628.n303 a_n1455_n3628.n301 0.573776
R17195 a_n1455_n3628.n328 a_n1455_n3628.n303 0.573776
R17196 a_n1455_n3628.n145 a_n1455_n3628.n119 0.573776
R17197 a_n1455_n3628.n119 a_n1455_n3628.n117 0.573776
R17198 a_n1455_n3628.n356 a_n1455_n3628.n65 0.573776
R17199 a_n1455_n3628.n356 a_n1455_n3628.n355 0.573776
R17200 a_n1455_n3628.n223 a_n1455_n3628.n222 0.422738
R17201 a_n1455_n3628.n340 a_n1455_n3628.n339 0.388379
R17202 a_n1455_n3628.n50 a_n1455_n3628.n49 0.388379
R17203 a_n1455_n3628.n102 a_n1455_n3628.n101 0.388379
R17204 a_n1455_n3628.n130 a_n1455_n3628.n129 0.388379
R17205 a_n1455_n3628.n76 a_n1455_n3628.n75 0.388379
R17206 a_n1455_n3628.n181 a_n1455_n3628.n180 0.388379
R17207 a_n1455_n3628.n207 a_n1455_n3628.n206 0.388379
R17208 a_n1455_n3628.n156 a_n1455_n3628.n155 0.388379
R17209 a_n1455_n3628.n314 a_n1455_n3628.n313 0.388379
R17210 a_n1455_n3628.n287 a_n1455_n3628.n286 0.388379
R17211 a_n1455_n3628.n262 a_n1455_n3628.n261 0.388379
R17212 a_n1455_n3628.n235 a_n1455_n3628.n234 0.388379
R17213 a_n1455_n3628.n39 a_n1455_n3628.n38 0.310845
R17214 a_n1455_n3628.n39 a_n1455_n3628.n37 0.310845
R17215 a_n1455_n3628.n37 a_n1455_n3628.n36 0.310845
R17216 a_n1455_n3628.n35 a_n1455_n3628.n34 0.310845
R17217 a_n1455_n3628.n35 a_n1455_n3628.n33 0.310845
R17218 a_n1455_n3628.n33 a_n1455_n3628.n32 0.310845
R17219 a_n1455_n3628.n31 a_n1455_n3628.n30 0.310845
R17220 a_n1455_n3628.n31 a_n1455_n3628.n29 0.310845
R17221 a_n1455_n3628.n29 a_n1455_n3628.n28 0.310845
R17222 a_n1455_n3628.n27 a_n1455_n3628.n26 0.310845
R17223 a_n1455_n3628.n27 a_n1455_n3628.n25 0.310845
R17224 a_n1455_n3628.n25 a_n1455_n3628.n24 0.310845
R17225 a_n1455_n3628.n23 a_n1455_n3628.n21 0.310845
R17226 a_n1455_n3628.n22 a_n1455_n3628.n21 0.310845
R17227 a_n1455_n3628.n169 a_n1455_n3628.n22 0.310845
R17228 a_n1455_n3628.n20 a_n1455_n3628.n18 0.310845
R17229 a_n1455_n3628.n19 a_n1455_n3628.n18 0.310845
R17230 a_n1455_n3628.n220 a_n1455_n3628.n19 0.310845
R17231 a_n1455_n3628.n17 a_n1455_n3628.n15 0.310845
R17232 a_n1455_n3628.n16 a_n1455_n3628.n15 0.310845
R17233 a_n1455_n3628.n194 a_n1455_n3628.n16 0.310845
R17234 a_n1455_n3628.n14 a_n1455_n3628.n12 0.310845
R17235 a_n1455_n3628.n13 a_n1455_n3628.n12 0.310845
R17236 a_n1455_n3628.n89 a_n1455_n3628.n13 0.310845
R17237 a_n1455_n3628.n11 a_n1455_n3628.n9 0.310845
R17238 a_n1455_n3628.n10 a_n1455_n3628.n9 0.310845
R17239 a_n1455_n3628.n143 a_n1455_n3628.n10 0.310845
R17240 a_n1455_n3628.n8 a_n1455_n3628.n6 0.310845
R17241 a_n1455_n3628.n7 a_n1455_n3628.n6 0.310845
R17242 a_n1455_n3628.n115 a_n1455_n3628.n7 0.310845
R17243 a_n1455_n3628.n5 a_n1455_n3628.n3 0.310845
R17244 a_n1455_n3628.n4 a_n1455_n3628.n3 0.310845
R17245 a_n1455_n3628.n63 a_n1455_n3628.n4 0.310845
R17246 a_n1455_n3628.n2 a_n1455_n3628.n0 0.310845
R17247 a_n1455_n3628.n1 a_n1455_n3628.n0 0.310845
R17248 a_n1455_n3628.n353 a_n1455_n3628.n1 0.310845
R17249 a_n1455_n3628.n301 a_n1455_n3628.n276 0.235414
R17250 a_n1455_n3628.n117 a_n1455_n3628.n65 0.235414
R17251 a_n2433_10060.n0 a_n2433_10060.n1 39.6373
R17252 a_n2433_10060.n2 a_n2433_10060.n3 39.6373
R17253 a_n2433_10060.n4 a_n2433_10060.n5 39.6373
R17254 a_n2433_10060.n6 a_n2433_10060.n7 39.6373
R17255 a_n2433_10060.n35 a_n2433_10060.n8 161.3
R17256 a_n2433_10060.n6 a_n2433_10060.n36 71.6402
R17257 a_n2433_10060.n10 a_n2433_10060.n9 39.6373
R17258 a_n2433_10060.n37 a_n2433_10060.n31 161.3
R17259 a_n2433_10060.n9 a_n2433_10060.n38 71.6402
R17260 a_n2433_10060.n12 a_n2433_10060.n46 161.3
R17261 a_n2433_10060.n13 a_n2433_10060.n39 71.6402
R17262 a_n2433_10060.n33 a_n2433_10060.t7 175.006
R17263 a_n2433_10060.n30 a_n2433_10060.t36 175.006
R17264 a_n2433_10060.n28 a_n2433_10060.t29 175.006
R17265 a_n2433_10060.n26 a_n2433_10060.t44 175.006
R17266 a_n2433_10060.n24 a_n2433_10060.t46 175.006
R17267 a_n2433_10060.n19 a_n2433_10060.t19 175.006
R17268 a_n2433_10060.n17 a_n2433_10060.t39 175.006
R17269 a_n2433_10060.n22 a_n2433_10060.t37 175.006
R17270 a_n2433_10060.n47 a_n2433_10060.t9 120.501
R17271 a_n2433_10060.n45 a_n2433_10060.t21 120.501
R17272 a_n2433_10060.n55 a_n2433_10060.t25 120.501
R17273 a_n2433_10060.n56 a_n2433_10060.t40 120.501
R17274 a_n2433_10060.n53 a_n2433_10060.t38 120.501
R17275 a_n2433_10060.n54 a_n2433_10060.t35 120.501
R17276 a_n2433_10060.n51 a_n2433_10060.t31 120.501
R17277 a_n2433_10060.n52 a_n2433_10060.t34 120.501
R17278 a_n2433_10060.n49 a_n2433_10060.t33 120.501
R17279 a_n2433_10060.n50 a_n2433_10060.t45 120.501
R17280 a_n2433_10060.n42 a_n2433_10060.t15 120.501
R17281 a_n2433_10060.n41 a_n2433_10060.t17 120.501
R17282 a_n2433_10060.n44 a_n2433_10060.t47 120.501
R17283 a_n2433_10060.n43 a_n2433_10060.t30 120.501
R17284 a_n2433_10060.n59 a_n2433_10060.t42 120.501
R17285 a_n2433_10060.n58 a_n2433_10060.t41 120.501
R17286 a_n2433_10060.n14 a_n2433_10060.t20 98.012
R17287 a_n2433_10060.n15 a_n2433_10060.t14 98.012
R17288 a_n2433_10060.n15 a_n2433_10060.t8 97.4387
R17289 a_n2433_10060.n14 a_n2433_10060.t12 97.4386
R17290 a_n2433_10060.n14 a_n2433_10060.n40 90.9378
R17291 a_n2433_10060.n15 a_n2433_10060.n48 90.9378
R17292 a_n2433_10060.n64 a_n2433_10060.n63 84.3504
R17293 a_n2433_10060.n16 a_n2433_10060.n60 84.3502
R17294 a_n2433_10060.n63 a_n2433_10060.n62 84.35
R17295 a_n2433_10060.n16 a_n2433_10060.n61 84.0635
R17296 a_n2433_10060.n18 a_n2433_10060.n0 43.5975
R17297 a_n2433_10060.n0 a_n2433_10060.n17 43.5975
R17298 a_n2433_10060.n21 a_n2433_10060.n2 43.5975
R17299 a_n2433_10060.n2 a_n2433_10060.n19 43.5975
R17300 a_n2433_10060.n23 a_n2433_10060.n4 43.5975
R17301 a_n2433_10060.n4 a_n2433_10060.n22 43.5975
R17302 a_n2433_10060.n6 a_n2433_10060.n25 43.5975
R17303 a_n2433_10060.n24 a_n2433_10060.n6 43.5975
R17304 a_n2433_10060.n8 a_n2433_10060.n27 43.5975
R17305 a_n2433_10060.n26 a_n2433_10060.n6 43.5975
R17306 a_n2433_10060.n9 a_n2433_10060.n29 43.5975
R17307 a_n2433_10060.n28 a_n2433_10060.n9 43.5975
R17308 a_n2433_10060.n31 a_n2433_10060.n32 43.5975
R17309 a_n2433_10060.n30 a_n2433_10060.n9 43.5975
R17310 a_n2433_10060.n34 a_n2433_10060.n12 43.5975
R17311 a_n2433_10060.n13 a_n2433_10060.n33 43.5975
R17312 a_n2433_10060.n34 a_n2433_10060.t13 175.006
R17313 a_n2433_10060.t28 a_n2433_10060.n32 175.006
R17314 a_n2433_10060.t24 a_n2433_10060.n29 175.006
R17315 a_n2433_10060.t26 a_n2433_10060.n27 175.006
R17316 a_n2433_10060.t27 a_n2433_10060.n25 175.006
R17317 a_n2433_10060.n21 a_n2433_10060.t11 175.006
R17318 a_n2433_10060.n18 a_n2433_10060.t43 175.006
R17319 a_n2433_10060.n23 a_n2433_10060.t32 175.006
R17320 a_n2433_10060.n39 a_n2433_10060.n46 58.5991
R17321 a_n2433_10060.n38 a_n2433_10060.n37 58.5991
R17322 a_n2433_10060.n10 a_n2433_10060.n54 40.5373
R17323 a_n2433_10060.n36 a_n2433_10060.n35 58.5991
R17324 a_n2433_10060.n49 a_n2433_10060.n7 40.5378
R17325 a_n2433_10060.n3 a_n2433_10060.n41 40.5373
R17326 a_n2433_10060.n44 a_n2433_10060.n1 40.5378
R17327 a_n2433_10060.n5 a_n2433_10060.n58 40.5373
R17328 a_n2433_10060.n63 a_n2433_10060.n16 29.8404
R17329 a_n2433_10060.n33 a_n2433_10060.n47 46.9373
R17330 a_n2433_10060.n45 a_n2433_10060.n34 46.9373
R17331 a_n2433_10060.n55 a_n2433_10060.n30 46.9373
R17332 a_n2433_10060.n32 a_n2433_10060.n56 46.9373
R17333 a_n2433_10060.n53 a_n2433_10060.n28 46.9373
R17334 a_n2433_10060.n29 a_n2433_10060.n54 46.9373
R17335 a_n2433_10060.n51 a_n2433_10060.n26 46.9373
R17336 a_n2433_10060.n27 a_n2433_10060.n52 46.9373
R17337 a_n2433_10060.n49 a_n2433_10060.n24 46.9373
R17338 a_n2433_10060.n25 a_n2433_10060.n50 46.9373
R17339 a_n2433_10060.n19 a_n2433_10060.n42 46.9373
R17340 a_n2433_10060.n41 a_n2433_10060.n21 46.9373
R17341 a_n2433_10060.n17 a_n2433_10060.n44 46.9373
R17342 a_n2433_10060.n43 a_n2433_10060.n18 46.9373
R17343 a_n2433_10060.n22 a_n2433_10060.n59 46.9373
R17344 a_n2433_10060.n58 a_n2433_10060.n23 46.9373
R17345 a_n2433_10060.n11 a_n2433_10060.n0 10.41
R17346 a_n2433_10060.n4 a_n2433_10060.n57 10.2055
R17347 a_n2433_10060.n11 a_n2433_10060.n13 8.90057
R17348 a_n2433_10060.n47 a_n2433_10060.n39 26.1378
R17349 a_n2433_10060.n46 a_n2433_10060.n45 8.11581
R17350 a_n2433_10060.n38 a_n2433_10060.n55 26.1378
R17351 a_n2433_10060.n56 a_n2433_10060.n37 8.11581
R17352 a_n2433_10060.n10 a_n2433_10060.n53 40.5378
R17353 a_n2433_10060.n36 a_n2433_10060.n51 26.1378
R17354 a_n2433_10060.n52 a_n2433_10060.n35 8.11581
R17355 a_n2433_10060.n50 a_n2433_10060.n7 40.5373
R17356 a_n2433_10060.n42 a_n2433_10060.n3 40.5378
R17357 a_n2433_10060.n1 a_n2433_10060.n43 40.5373
R17358 a_n2433_10060.n59 a_n2433_10060.n5 40.5378
R17359 a_n2433_10060.n16 a_n2433_10060.n12 24.257
R17360 a_n2433_10060.n20 a_n2433_10060.n14 8.39986
R17361 a_n2433_10060.n0 a_n2433_10060.n2 7.30241
R17362 a_n2433_10060.n6 a_n2433_10060.n11 7.20928
R17363 a_n2433_10060.n2 a_n2433_10060.n20 6.58049
R17364 a_n2433_10060.n40 a_n2433_10060.t16 6.5015
R17365 a_n2433_10060.n40 a_n2433_10060.t18 6.5015
R17366 a_n2433_10060.n48 a_n2433_10060.t10 6.5015
R17367 a_n2433_10060.n48 a_n2433_10060.t22 6.5015
R17368 a_n2433_10060.n11 a_n2433_10060.n15 6.07162
R17369 a_n2433_10060.n57 a_n2433_10060.n31 5.90435
R17370 a_n2433_10060.n12 a_n2433_10060.n4 4.84653
R17371 a_n2433_10060.n57 a_n2433_10060.n20 3.83005
R17372 a_n2433_10060.n8 a_n2433_10060.n6 3.6168
R17373 a_n2433_10060.n62 a_n2433_10060.t2 3.3005
R17374 a_n2433_10060.n62 a_n2433_10060.t3 3.3005
R17375 a_n2433_10060.n60 a_n2433_10060.t1 3.3005
R17376 a_n2433_10060.n60 a_n2433_10060.t4 3.3005
R17377 a_n2433_10060.n61 a_n2433_10060.t5 3.3005
R17378 a_n2433_10060.n61 a_n2433_10060.t6 3.3005
R17379 a_n2433_10060.t0 a_n2433_10060.n64 3.3005
R17380 a_n2433_10060.n64 a_n2433_10060.t23 3.3005
R17381 a_n2433_10060.n9 a_n2433_10060.n8 2.75228
R17382 a_n2433_10060.n13 a_n2433_10060.n12 2.4185
R17383 a_n2433_10060.n31 a_n2433_10060.n9 2.29016
R17384 a_n2511_10256.n5 a_n2511_10256.n3 119.439
R17385 a_n2511_10256.n8 a_n2511_10256.n6 119.1
R17386 a_n2511_10256.n8 a_n2511_10256.n7 118.865
R17387 a_n2511_10256.n5 a_n2511_10256.n4 118.865
R17388 a_n2511_10256.n2 a_n2511_10256.t4 98.012
R17389 a_n2511_10256.n10 a_n2511_10256.t5 97.4387
R17390 a_n2511_10256.n0 a_n2511_10256.t2 97.4387
R17391 a_n2511_10256.t7 a_n2511_10256.n0 97.4387
R17392 a_n2511_10256.n12 a_n2511_10256.n11 90.9378
R17393 a_n2511_10256.n2 a_n2511_10256.n1 90.9378
R17394 a_n2511_10256.n9 a_n2511_10256.n8 12.2276
R17395 a_n2511_10256.n9 a_n2511_10256.n5 10.0093
R17396 a_n2511_10256.n11 a_n2511_10256.t6 6.5015
R17397 a_n2511_10256.n11 a_n2511_10256.t0 6.5015
R17398 a_n2511_10256.n1 a_n2511_10256.t1 6.5015
R17399 a_n2511_10256.n1 a_n2511_10256.t3 6.5015
R17400 a_n2511_10256.n4 a_n2511_10256.t13 6.5015
R17401 a_n2511_10256.n4 a_n2511_10256.t10 6.5015
R17402 a_n2511_10256.n3 a_n2511_10256.t8 6.5015
R17403 a_n2511_10256.n3 a_n2511_10256.t12 6.5015
R17404 a_n2511_10256.n7 a_n2511_10256.t9 6.5015
R17405 a_n2511_10256.n7 a_n2511_10256.t11 6.5015
R17406 a_n2511_10256.n6 a_n2511_10256.t14 6.5015
R17407 a_n2511_10256.n6 a_n2511_10256.t15 6.5015
R17408 a_n2511_10256.n10 a_n2511_10256.n9 5.29253
R17409 a_n2511_10256.n0 a_n2511_10256.n2 0.728948
R17410 a_n2511_10256.n0 a_n2511_10256.n12 0.573776
R17411 a_n2511_10256.n12 a_n2511_10256.n10 0.573776
R17412 VP.n30 VP.t3 243.255
R17413 VP.n29 VP.n27 224.169
R17414 VP.n29 VP.n28 223.454
R17415 VP.n15 VP.t9 199.144
R17416 VP.n2 VP.t11 199.144
R17417 VP.n24 VP.t7 183.883
R17418 VP.n11 VP.t5 183.883
R17419 VP.n18 VP.n17 161.3
R17420 VP.n19 VP.n14 161.3
R17421 VP.n21 VP.n20 161.3
R17422 VP.n23 VP.n13 161.3
R17423 VP.n10 VP.n0 161.3
R17424 VP.n8 VP.n7 161.3
R17425 VP.n6 VP.n1 161.3
R17426 VP.n5 VP.n4 161.3
R17427 VP.n22 VP.t12 144.601
R17428 VP.n16 VP.t8 144.601
R17429 VP.n3 VP.t10 144.601
R17430 VP.n9 VP.t6 144.601
R17431 VP.n25 VP.n24 80.6037
R17432 VP.n12 VP.n11 80.6037
R17433 VP.n24 VP.n23 56.3158
R17434 VP.n11 VP.n10 56.3158
R17435 VP.n16 VP.n15 46.9082
R17436 VP.n3 VP.n2 46.9082
R17437 VP.n5 VP.n2 43.8991
R17438 VP.n18 VP.n15 43.8991
R17439 VP.n21 VP.n14 40.577
R17440 VP.n17 VP.n14 40.577
R17441 VP.n4 VP.n1 40.577
R17442 VP.n8 VP.n1 40.577
R17443 VP.n26 VP.n25 28.1089
R17444 VP.n28 VP.t0 19.8005
R17445 VP.n28 VP.t2 19.8005
R17446 VP.n27 VP.t4 19.8005
R17447 VP.n27 VP.t1 19.8005
R17448 VP.n23 VP.n22 16.477
R17449 VP.n10 VP.n9 16.477
R17450 VP.n26 VP.n12 11.9157
R17451 VP VP.n31 11.5274
R17452 VP.n22 VP.n21 8.11581
R17453 VP.n17 VP.n16 8.11581
R17454 VP.n4 VP.n3 8.11581
R17455 VP.n9 VP.n8 8.11581
R17456 VP.n31 VP.n30 4.80222
R17457 VP.n31 VP.n26 0.972091
R17458 VP.n30 VP.n29 0.716017
R17459 VP.n25 VP.n13 0.285035
R17460 VP.n12 VP.n0 0.285035
R17461 VP.n20 VP.n13 0.189894
R17462 VP.n20 VP.n19 0.189894
R17463 VP.n19 VP.n18 0.189894
R17464 VP.n6 VP.n5 0.189894
R17465 VP.n7 VP.n6 0.189894
R17466 VP.n7 VP.n0 0.189894
R17467 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n1 289.615
R17468 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n32 289.615
R17469 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n64 289.615
R17470 DIFFPAIR_BIAS.n122 DIFFPAIR_BIAS.n96 289.615
R17471 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n27 185
R17472 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n25 185
R17473 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 185
R17474 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n19 185
R17475 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n17 185
R17476 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 185
R17477 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 185
R17478 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n58 185
R17479 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n56 185
R17480 DIFFPAIR_BIAS.n36 DIFFPAIR_BIAS.n35 185
R17481 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n50 185
R17482 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n48 185
R17483 DIFFPAIR_BIAS.n40 DIFFPAIR_BIAS.n39 185
R17484 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n42 185
R17485 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n90 185
R17486 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n88 185
R17487 DIFFPAIR_BIAS.n68 DIFFPAIR_BIAS.n67 185
R17488 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n82 185
R17489 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n80 185
R17490 DIFFPAIR_BIAS.n72 DIFFPAIR_BIAS.n71 185
R17491 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n74 185
R17492 DIFFPAIR_BIAS.n123 DIFFPAIR_BIAS.n122 185
R17493 DIFFPAIR_BIAS.n121 DIFFPAIR_BIAS.n120 185
R17494 DIFFPAIR_BIAS.n100 DIFFPAIR_BIAS.n99 185
R17495 DIFFPAIR_BIAS.n115 DIFFPAIR_BIAS.n114 185
R17496 DIFFPAIR_BIAS.n113 DIFFPAIR_BIAS.n112 185
R17497 DIFFPAIR_BIAS.n104 DIFFPAIR_BIAS.n103 185
R17498 DIFFPAIR_BIAS.n107 DIFFPAIR_BIAS.n106 185
R17499 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t9 178.945
R17500 DIFFPAIR_BIAS.n133 DIFFPAIR_BIAS.t10 177.018
R17501 DIFFPAIR_BIAS.n132 DIFFPAIR_BIAS.t11 177.018
R17502 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t8 177.018
R17503 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.n10 147.661
R17504 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.n41 147.661
R17505 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.n73 147.661
R17506 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.n105 147.661
R17507 DIFFPAIR_BIAS.n128 DIFFPAIR_BIAS.t0 132.363
R17508 DIFFPAIR_BIAS.n128 DIFFPAIR_BIAS.t2 130.436
R17509 DIFFPAIR_BIAS.n129 DIFFPAIR_BIAS.t4 130.436
R17510 DIFFPAIR_BIAS.n130 DIFFPAIR_BIAS.t6 130.436
R17511 DIFFPAIR_BIAS.n27 DIFFPAIR_BIAS.n26 104.615
R17512 DIFFPAIR_BIAS.n26 DIFFPAIR_BIAS.n4 104.615
R17513 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n4 104.615
R17514 DIFFPAIR_BIAS.n19 DIFFPAIR_BIAS.n18 104.615
R17515 DIFFPAIR_BIAS.n18 DIFFPAIR_BIAS.n8 104.615
R17516 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n8 104.615
R17517 DIFFPAIR_BIAS.n58 DIFFPAIR_BIAS.n57 104.615
R17518 DIFFPAIR_BIAS.n57 DIFFPAIR_BIAS.n35 104.615
R17519 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n35 104.615
R17520 DIFFPAIR_BIAS.n50 DIFFPAIR_BIAS.n49 104.615
R17521 DIFFPAIR_BIAS.n49 DIFFPAIR_BIAS.n39 104.615
R17522 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.n39 104.615
R17523 DIFFPAIR_BIAS.n90 DIFFPAIR_BIAS.n89 104.615
R17524 DIFFPAIR_BIAS.n89 DIFFPAIR_BIAS.n67 104.615
R17525 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n67 104.615
R17526 DIFFPAIR_BIAS.n82 DIFFPAIR_BIAS.n81 104.615
R17527 DIFFPAIR_BIAS.n81 DIFFPAIR_BIAS.n71 104.615
R17528 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.n71 104.615
R17529 DIFFPAIR_BIAS.n122 DIFFPAIR_BIAS.n121 104.615
R17530 DIFFPAIR_BIAS.n121 DIFFPAIR_BIAS.n99 104.615
R17531 DIFFPAIR_BIAS.n114 DIFFPAIR_BIAS.n99 104.615
R17532 DIFFPAIR_BIAS.n114 DIFFPAIR_BIAS.n113 104.615
R17533 DIFFPAIR_BIAS.n113 DIFFPAIR_BIAS.n103 104.615
R17534 DIFFPAIR_BIAS.n106 DIFFPAIR_BIAS.n103 104.615
R17535 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n31 95.6354
R17536 DIFFPAIR_BIAS.n63 DIFFPAIR_BIAS.n62 94.6732
R17537 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.n94 94.6732
R17538 DIFFPAIR_BIAS.n127 DIFFPAIR_BIAS.n126 94.6732
R17539 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.t1 52.3082
R17540 DIFFPAIR_BIAS.n42 DIFFPAIR_BIAS.t3 52.3082
R17541 DIFFPAIR_BIAS.n74 DIFFPAIR_BIAS.t5 52.3082
R17542 DIFFPAIR_BIAS.n106 DIFFPAIR_BIAS.t7 52.3082
R17543 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n10 15.6674
R17544 DIFFPAIR_BIAS.n43 DIFFPAIR_BIAS.n41 15.6674
R17545 DIFFPAIR_BIAS.n75 DIFFPAIR_BIAS.n73 15.6674
R17546 DIFFPAIR_BIAS.n107 DIFFPAIR_BIAS.n105 15.6674
R17547 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n9 12.8005
R17548 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n40 12.8005
R17549 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n72 12.8005
R17550 DIFFPAIR_BIAS.n108 DIFFPAIR_BIAS.n104 12.8005
R17551 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n16 12.0247
R17552 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n47 12.0247
R17553 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n79 12.0247
R17554 DIFFPAIR_BIAS.n112 DIFFPAIR_BIAS.n111 12.0247
R17555 DIFFPAIR_BIAS.n20 DIFFPAIR_BIAS.n7 11.249
R17556 DIFFPAIR_BIAS.n51 DIFFPAIR_BIAS.n38 11.249
R17557 DIFFPAIR_BIAS.n83 DIFFPAIR_BIAS.n70 11.249
R17558 DIFFPAIR_BIAS.n115 DIFFPAIR_BIAS.n102 11.249
R17559 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n5 10.4732
R17560 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n36 10.4732
R17561 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n68 10.4732
R17562 DIFFPAIR_BIAS.n116 DIFFPAIR_BIAS.n100 10.4732
R17563 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n24 9.69747
R17564 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n55 9.69747
R17565 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n87 9.69747
R17566 DIFFPAIR_BIAS.n120 DIFFPAIR_BIAS.n119 9.69747
R17567 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n30 9.45567
R17568 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n61 9.45567
R17569 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n93 9.45567
R17570 DIFFPAIR_BIAS.n126 DIFFPAIR_BIAS.n125 9.45567
R17571 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n29 9.3005
R17572 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 9.3005
R17573 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n23 9.3005
R17574 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n21 9.3005
R17575 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 9.3005
R17576 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n15 9.3005
R17577 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n13 9.3005
R17578 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n60 9.3005
R17579 DIFFPAIR_BIAS.n34 DIFFPAIR_BIAS.n33 9.3005
R17580 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n54 9.3005
R17581 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n52 9.3005
R17582 DIFFPAIR_BIAS.n38 DIFFPAIR_BIAS.n37 9.3005
R17583 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n46 9.3005
R17584 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n44 9.3005
R17585 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n92 9.3005
R17586 DIFFPAIR_BIAS.n66 DIFFPAIR_BIAS.n65 9.3005
R17587 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n86 9.3005
R17588 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n84 9.3005
R17589 DIFFPAIR_BIAS.n70 DIFFPAIR_BIAS.n69 9.3005
R17590 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n78 9.3005
R17591 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n76 9.3005
R17592 DIFFPAIR_BIAS.n125 DIFFPAIR_BIAS.n124 9.3005
R17593 DIFFPAIR_BIAS.n98 DIFFPAIR_BIAS.n97 9.3005
R17594 DIFFPAIR_BIAS.n119 DIFFPAIR_BIAS.n118 9.3005
R17595 DIFFPAIR_BIAS.n117 DIFFPAIR_BIAS.n116 9.3005
R17596 DIFFPAIR_BIAS.n102 DIFFPAIR_BIAS.n101 9.3005
R17597 DIFFPAIR_BIAS.n111 DIFFPAIR_BIAS.n110 9.3005
R17598 DIFFPAIR_BIAS.n109 DIFFPAIR_BIAS.n108 9.3005
R17599 DIFFPAIR_BIAS.n28 DIFFPAIR_BIAS.n3 8.92171
R17600 DIFFPAIR_BIAS.n59 DIFFPAIR_BIAS.n34 8.92171
R17601 DIFFPAIR_BIAS.n91 DIFFPAIR_BIAS.n66 8.92171
R17602 DIFFPAIR_BIAS.n123 DIFFPAIR_BIAS.n98 8.92171
R17603 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n1 8.14595
R17604 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n32 8.14595
R17605 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n64 8.14595
R17606 DIFFPAIR_BIAS.n124 DIFFPAIR_BIAS.n96 8.14595
R17607 DIFFPAIR_BIAS.n31 DIFFPAIR_BIAS.n1 5.81868
R17608 DIFFPAIR_BIAS.n62 DIFFPAIR_BIAS.n32 5.81868
R17609 DIFFPAIR_BIAS.n94 DIFFPAIR_BIAS.n64 5.81868
R17610 DIFFPAIR_BIAS.n126 DIFFPAIR_BIAS.n96 5.81868
R17611 DIFFPAIR_BIAS.n131 DIFFPAIR_BIAS.n130 5.20947
R17612 DIFFPAIR_BIAS.n29 DIFFPAIR_BIAS.n28 5.04292
R17613 DIFFPAIR_BIAS.n60 DIFFPAIR_BIAS.n59 5.04292
R17614 DIFFPAIR_BIAS.n92 DIFFPAIR_BIAS.n91 5.04292
R17615 DIFFPAIR_BIAS.n124 DIFFPAIR_BIAS.n123 5.04292
R17616 DIFFPAIR_BIAS.n131 DIFFPAIR_BIAS.n127 4.42209
R17617 DIFFPAIR_BIAS.n14 DIFFPAIR_BIAS.n10 4.38594
R17618 DIFFPAIR_BIAS.n45 DIFFPAIR_BIAS.n41 4.38594
R17619 DIFFPAIR_BIAS.n77 DIFFPAIR_BIAS.n73 4.38594
R17620 DIFFPAIR_BIAS.n109 DIFFPAIR_BIAS.n105 4.38594
R17621 DIFFPAIR_BIAS.n132 DIFFPAIR_BIAS.n131 4.28454
R17622 DIFFPAIR_BIAS.n25 DIFFPAIR_BIAS.n3 4.26717
R17623 DIFFPAIR_BIAS.n56 DIFFPAIR_BIAS.n34 4.26717
R17624 DIFFPAIR_BIAS.n88 DIFFPAIR_BIAS.n66 4.26717
R17625 DIFFPAIR_BIAS.n120 DIFFPAIR_BIAS.n98 4.26717
R17626 DIFFPAIR_BIAS.n24 DIFFPAIR_BIAS.n5 3.49141
R17627 DIFFPAIR_BIAS.n55 DIFFPAIR_BIAS.n36 3.49141
R17628 DIFFPAIR_BIAS.n87 DIFFPAIR_BIAS.n68 3.49141
R17629 DIFFPAIR_BIAS.n119 DIFFPAIR_BIAS.n100 3.49141
R17630 DIFFPAIR_BIAS.n21 DIFFPAIR_BIAS.n20 2.71565
R17631 DIFFPAIR_BIAS.n52 DIFFPAIR_BIAS.n51 2.71565
R17632 DIFFPAIR_BIAS.n84 DIFFPAIR_BIAS.n83 2.71565
R17633 DIFFPAIR_BIAS.n116 DIFFPAIR_BIAS.n115 2.71565
R17634 DIFFPAIR_BIAS.n17 DIFFPAIR_BIAS.n7 1.93989
R17635 DIFFPAIR_BIAS.n48 DIFFPAIR_BIAS.n38 1.93989
R17636 DIFFPAIR_BIAS.n80 DIFFPAIR_BIAS.n70 1.93989
R17637 DIFFPAIR_BIAS.n112 DIFFPAIR_BIAS.n102 1.93989
R17638 DIFFPAIR_BIAS.n130 DIFFPAIR_BIAS.n129 1.9266
R17639 DIFFPAIR_BIAS.n129 DIFFPAIR_BIAS.n128 1.9266
R17640 DIFFPAIR_BIAS.n133 DIFFPAIR_BIAS.n132 1.92658
R17641 DIFFPAIR_BIAS.n134 DIFFPAIR_BIAS.n133 1.29913
R17642 DIFFPAIR_BIAS.n16 DIFFPAIR_BIAS.n9 1.16414
R17643 DIFFPAIR_BIAS.n47 DIFFPAIR_BIAS.n40 1.16414
R17644 DIFFPAIR_BIAS.n79 DIFFPAIR_BIAS.n72 1.16414
R17645 DIFFPAIR_BIAS.n111 DIFFPAIR_BIAS.n104 1.16414
R17646 DIFFPAIR_BIAS.n127 DIFFPAIR_BIAS.n95 0.962709
R17647 DIFFPAIR_BIAS.n95 DIFFPAIR_BIAS.n63 0.962709
R17648 DIFFPAIR_BIAS DIFFPAIR_BIAS.n134 0.684875
R17649 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 0.388379
R17650 DIFFPAIR_BIAS.n44 DIFFPAIR_BIAS.n43 0.388379
R17651 DIFFPAIR_BIAS.n76 DIFFPAIR_BIAS.n75 0.388379
R17652 DIFFPAIR_BIAS.n108 DIFFPAIR_BIAS.n107 0.388379
R17653 DIFFPAIR_BIAS.n134 DIFFPAIR_BIAS.n0 0.337251
R17654 DIFFPAIR_BIAS.n30 DIFFPAIR_BIAS.n2 0.155672
R17655 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n2 0.155672
R17656 DIFFPAIR_BIAS.n23 DIFFPAIR_BIAS.n22 0.155672
R17657 DIFFPAIR_BIAS.n22 DIFFPAIR_BIAS.n6 0.155672
R17658 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n6 0.155672
R17659 DIFFPAIR_BIAS.n15 DIFFPAIR_BIAS.n14 0.155672
R17660 DIFFPAIR_BIAS.n61 DIFFPAIR_BIAS.n33 0.155672
R17661 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n33 0.155672
R17662 DIFFPAIR_BIAS.n54 DIFFPAIR_BIAS.n53 0.155672
R17663 DIFFPAIR_BIAS.n53 DIFFPAIR_BIAS.n37 0.155672
R17664 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n37 0.155672
R17665 DIFFPAIR_BIAS.n46 DIFFPAIR_BIAS.n45 0.155672
R17666 DIFFPAIR_BIAS.n93 DIFFPAIR_BIAS.n65 0.155672
R17667 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n65 0.155672
R17668 DIFFPAIR_BIAS.n86 DIFFPAIR_BIAS.n85 0.155672
R17669 DIFFPAIR_BIAS.n85 DIFFPAIR_BIAS.n69 0.155672
R17670 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n69 0.155672
R17671 DIFFPAIR_BIAS.n78 DIFFPAIR_BIAS.n77 0.155672
R17672 DIFFPAIR_BIAS.n125 DIFFPAIR_BIAS.n97 0.155672
R17673 DIFFPAIR_BIAS.n118 DIFFPAIR_BIAS.n97 0.155672
R17674 DIFFPAIR_BIAS.n118 DIFFPAIR_BIAS.n117 0.155672
R17675 DIFFPAIR_BIAS.n117 DIFFPAIR_BIAS.n101 0.155672
R17676 DIFFPAIR_BIAS.n110 DIFFPAIR_BIAS.n101 0.155672
R17677 DIFFPAIR_BIAS.n110 DIFFPAIR_BIAS.n109 0.155672
R17678 a_n2154_8322.n6 a_n2154_8322.t14 98.012
R17679 a_n2154_8322.t7 a_n2154_8322.n13 98.012
R17680 a_n2154_8322.n2 a_n2154_8322.t9 98.0119
R17681 a_n2154_8322.n0 a_n2154_8322.t2 97.4387
R17682 a_n2154_8322.n0 a_n2154_8322.t6 97.4387
R17683 a_n2154_8322.n9 a_n2154_8322.t0 97.4387
R17684 a_n2154_8322.n3 a_n2154_8322.t12 97.4387
R17685 a_n2154_8322.n7 a_n2154_8322.t13 97.4387
R17686 a_n2154_8322.n13 a_n2154_8322.n12 90.9378
R17687 a_n2154_8322.n11 a_n2154_8322.n10 90.9378
R17688 a_n2154_8322.n2 a_n2154_8322.n1 90.9378
R17689 a_n2154_8322.n6 a_n2154_8322.n5 90.9378
R17690 a_n2154_8322.n8 a_n2154_8322.n7 21.3698
R17691 a_n2154_8322.n4 a_n2154_8322.t16 8.84949
R17692 a_n2154_8322.n12 a_n2154_8322.t5 6.5015
R17693 a_n2154_8322.n12 a_n2154_8322.t3 6.5015
R17694 a_n2154_8322.n10 a_n2154_8322.t4 6.5015
R17695 a_n2154_8322.n10 a_n2154_8322.t1 6.5015
R17696 a_n2154_8322.n1 a_n2154_8322.t8 6.5015
R17697 a_n2154_8322.n1 a_n2154_8322.t15 6.5015
R17698 a_n2154_8322.n5 a_n2154_8322.t10 6.5015
R17699 a_n2154_8322.n5 a_n2154_8322.t11 6.5015
R17700 a_n2154_8322.n4 a_n2154_8322.n3 5.67722
R17701 a_n2154_8322.n9 a_n2154_8322.n8 5.29253
R17702 a_n2154_8322.n8 a_n2154_8322.n4 3.83005
R17703 a_n2154_8322.n13 a_n2154_8322.n0 0.728948
R17704 a_n2154_8322.n3 a_n2154_8322.n2 0.573776
R17705 a_n2154_8322.n7 a_n2154_8322.n6 0.573776
R17706 a_n2154_8322.n11 a_n2154_8322.n9 0.573776
R17707 a_n2154_8322.n0 a_n2154_8322.n11 0.573776
C0 VN DIFFPAIR_BIAS 2.16e-19
C1 CS_BIAS DIFFPAIR_BIAS 0.008433f
C2 VDD VOUT 54.2099f
C3 VDD VN 0.059349f
C4 VOUT VP 2.74686f
C5 VOUT VN 0.804612f
C6 VOUT CS_BIAS 23.0378f
C7 VP VN 7.84338f
C8 VP CS_BIAS 0.306594f
C9 VN CS_BIAS 0.266289f
C10 VP DIFFPAIR_BIAS 2.16e-19
C11 DIFFPAIR_BIAS GND 32.760902f
C12 CS_BIAS GND 0.11115p
C13 VN GND 25.75502f
C14 VP GND 22.45488f
C15 VOUT GND 62.252483f
C16 VDD GND 0.299201p
C17 a_n2154_8322.n0 GND 0.546541f
C18 a_n2154_8322.t16 GND 94.200096f
C19 a_n2154_8322.t9 GND 0.315967f
C20 a_n2154_8322.t8 GND 0.03909f
C21 a_n2154_8322.t15 GND 0.03909f
C22 a_n2154_8322.n1 GND 0.227514f
C23 a_n2154_8322.n2 GND 0.566827f
C24 a_n2154_8322.t12 GND 0.314439f
C25 a_n2154_8322.n3 GND 0.531848f
C26 a_n2154_8322.n4 GND 1.28703f
C27 a_n2154_8322.t14 GND 0.315969f
C28 a_n2154_8322.t10 GND 0.03909f
C29 a_n2154_8322.t11 GND 0.03909f
C30 a_n2154_8322.n5 GND 0.227514f
C31 a_n2154_8322.n6 GND 0.566825f
C32 a_n2154_8322.t13 GND 0.314439f
C33 a_n2154_8322.n7 GND 0.994496f
C34 a_n2154_8322.n8 GND 1.03933f
C35 a_n2154_8322.t0 GND 0.314439f
C36 a_n2154_8322.n9 GND 0.450407f
C37 a_n2154_8322.t4 GND 0.03909f
C38 a_n2154_8322.t1 GND 0.03909f
C39 a_n2154_8322.n10 GND 0.227514f
C40 a_n2154_8322.n11 GND 0.306901f
C41 a_n2154_8322.t6 GND 0.314439f
C42 a_n2154_8322.t2 GND 0.314439f
C43 a_n2154_8322.t5 GND 0.03909f
C44 a_n2154_8322.t3 GND 0.03909f
C45 a_n2154_8322.n12 GND 0.227514f
C46 a_n2154_8322.n13 GND 0.566825f
C47 a_n2154_8322.t7 GND 0.315969f
C48 DIFFPAIR_BIAS.t8 GND 0.108432f
C49 DIFFPAIR_BIAS.t9 GND 0.109185f
C50 DIFFPAIR_BIAS.n0 GND 0.122922f
C51 DIFFPAIR_BIAS.n1 GND 0.001296f
C52 DIFFPAIR_BIAS.n2 GND 9.22e-19
C53 DIFFPAIR_BIAS.n3 GND 4.95e-19
C54 DIFFPAIR_BIAS.n4 GND 0.001171f
C55 DIFFPAIR_BIAS.n5 GND 5.25e-19
C56 DIFFPAIR_BIAS.n6 GND 9.22e-19
C57 DIFFPAIR_BIAS.n7 GND 4.95e-19
C58 DIFFPAIR_BIAS.n8 GND 0.001171f
C59 DIFFPAIR_BIAS.n9 GND 5.25e-19
C60 DIFFPAIR_BIAS.n10 GND 0.003945f
C61 DIFFPAIR_BIAS.t1 GND 0.001909f
C62 DIFFPAIR_BIAS.n11 GND 8.78e-19
C63 DIFFPAIR_BIAS.n12 GND 6.92e-19
C64 DIFFPAIR_BIAS.n13 GND 4.95e-19
C65 DIFFPAIR_BIAS.n14 GND 0.021937f
C66 DIFFPAIR_BIAS.n15 GND 9.22e-19
C67 DIFFPAIR_BIAS.n16 GND 4.95e-19
C68 DIFFPAIR_BIAS.n17 GND 5.25e-19
C69 DIFFPAIR_BIAS.n18 GND 0.001171f
C70 DIFFPAIR_BIAS.n19 GND 0.001171f
C71 DIFFPAIR_BIAS.n20 GND 5.25e-19
C72 DIFFPAIR_BIAS.n21 GND 4.95e-19
C73 DIFFPAIR_BIAS.n22 GND 9.22e-19
C74 DIFFPAIR_BIAS.n23 GND 9.22e-19
C75 DIFFPAIR_BIAS.n24 GND 4.95e-19
C76 DIFFPAIR_BIAS.n25 GND 5.25e-19
C77 DIFFPAIR_BIAS.n26 GND 0.001171f
C78 DIFFPAIR_BIAS.n27 GND 0.002535f
C79 DIFFPAIR_BIAS.n28 GND 5.25e-19
C80 DIFFPAIR_BIAS.n29 GND 4.95e-19
C81 DIFFPAIR_BIAS.n30 GND 0.002131f
C82 DIFFPAIR_BIAS.n31 GND 0.005461f
C83 DIFFPAIR_BIAS.n32 GND 0.001296f
C84 DIFFPAIR_BIAS.n33 GND 9.22e-19
C85 DIFFPAIR_BIAS.n34 GND 4.95e-19
C86 DIFFPAIR_BIAS.n35 GND 0.001171f
C87 DIFFPAIR_BIAS.n36 GND 5.25e-19
C88 DIFFPAIR_BIAS.n37 GND 9.22e-19
C89 DIFFPAIR_BIAS.n38 GND 4.95e-19
C90 DIFFPAIR_BIAS.n39 GND 0.001171f
C91 DIFFPAIR_BIAS.n40 GND 5.25e-19
C92 DIFFPAIR_BIAS.n41 GND 0.003945f
C93 DIFFPAIR_BIAS.t3 GND 0.001909f
C94 DIFFPAIR_BIAS.n42 GND 8.78e-19
C95 DIFFPAIR_BIAS.n43 GND 6.92e-19
C96 DIFFPAIR_BIAS.n44 GND 4.95e-19
C97 DIFFPAIR_BIAS.n45 GND 0.021937f
C98 DIFFPAIR_BIAS.n46 GND 9.22e-19
C99 DIFFPAIR_BIAS.n47 GND 4.95e-19
C100 DIFFPAIR_BIAS.n48 GND 5.25e-19
C101 DIFFPAIR_BIAS.n49 GND 0.001171f
C102 DIFFPAIR_BIAS.n50 GND 0.001171f
C103 DIFFPAIR_BIAS.n51 GND 5.25e-19
C104 DIFFPAIR_BIAS.n52 GND 4.95e-19
C105 DIFFPAIR_BIAS.n53 GND 9.22e-19
C106 DIFFPAIR_BIAS.n54 GND 9.22e-19
C107 DIFFPAIR_BIAS.n55 GND 4.95e-19
C108 DIFFPAIR_BIAS.n56 GND 5.25e-19
C109 DIFFPAIR_BIAS.n57 GND 0.001171f
C110 DIFFPAIR_BIAS.n58 GND 0.002535f
C111 DIFFPAIR_BIAS.n59 GND 5.25e-19
C112 DIFFPAIR_BIAS.n60 GND 4.95e-19
C113 DIFFPAIR_BIAS.n61 GND 0.002131f
C114 DIFFPAIR_BIAS.n62 GND 0.00491f
C115 DIFFPAIR_BIAS.n63 GND 0.11516f
C116 DIFFPAIR_BIAS.n64 GND 0.001296f
C117 DIFFPAIR_BIAS.n65 GND 9.22e-19
C118 DIFFPAIR_BIAS.n66 GND 4.95e-19
C119 DIFFPAIR_BIAS.n67 GND 0.001171f
C120 DIFFPAIR_BIAS.n68 GND 5.25e-19
C121 DIFFPAIR_BIAS.n69 GND 9.22e-19
C122 DIFFPAIR_BIAS.n70 GND 4.95e-19
C123 DIFFPAIR_BIAS.n71 GND 0.001171f
C124 DIFFPAIR_BIAS.n72 GND 5.25e-19
C125 DIFFPAIR_BIAS.n73 GND 0.003945f
C126 DIFFPAIR_BIAS.t5 GND 0.001909f
C127 DIFFPAIR_BIAS.n74 GND 8.78e-19
C128 DIFFPAIR_BIAS.n75 GND 6.92e-19
C129 DIFFPAIR_BIAS.n76 GND 4.95e-19
C130 DIFFPAIR_BIAS.n77 GND 0.021937f
C131 DIFFPAIR_BIAS.n78 GND 9.22e-19
C132 DIFFPAIR_BIAS.n79 GND 4.95e-19
C133 DIFFPAIR_BIAS.n80 GND 5.25e-19
C134 DIFFPAIR_BIAS.n81 GND 0.001171f
C135 DIFFPAIR_BIAS.n82 GND 0.001171f
C136 DIFFPAIR_BIAS.n83 GND 5.25e-19
C137 DIFFPAIR_BIAS.n84 GND 4.95e-19
C138 DIFFPAIR_BIAS.n85 GND 9.22e-19
C139 DIFFPAIR_BIAS.n86 GND 9.22e-19
C140 DIFFPAIR_BIAS.n87 GND 4.95e-19
C141 DIFFPAIR_BIAS.n88 GND 5.25e-19
C142 DIFFPAIR_BIAS.n89 GND 0.001171f
C143 DIFFPAIR_BIAS.n90 GND 0.002535f
C144 DIFFPAIR_BIAS.n91 GND 5.25e-19
C145 DIFFPAIR_BIAS.n92 GND 4.95e-19
C146 DIFFPAIR_BIAS.n93 GND 0.002131f
C147 DIFFPAIR_BIAS.n94 GND 0.00491f
C148 DIFFPAIR_BIAS.n95 GND 0.06095f
C149 DIFFPAIR_BIAS.n96 GND 0.001296f
C150 DIFFPAIR_BIAS.n97 GND 9.22e-19
C151 DIFFPAIR_BIAS.n98 GND 4.95e-19
C152 DIFFPAIR_BIAS.n99 GND 0.001171f
C153 DIFFPAIR_BIAS.n100 GND 5.25e-19
C154 DIFFPAIR_BIAS.n101 GND 9.22e-19
C155 DIFFPAIR_BIAS.n102 GND 4.95e-19
C156 DIFFPAIR_BIAS.n103 GND 0.001171f
C157 DIFFPAIR_BIAS.n104 GND 5.25e-19
C158 DIFFPAIR_BIAS.n105 GND 0.003945f
C159 DIFFPAIR_BIAS.t7 GND 0.001909f
C160 DIFFPAIR_BIAS.n106 GND 8.78e-19
C161 DIFFPAIR_BIAS.n107 GND 6.92e-19
C162 DIFFPAIR_BIAS.n108 GND 4.95e-19
C163 DIFFPAIR_BIAS.n109 GND 0.021937f
C164 DIFFPAIR_BIAS.n110 GND 9.22e-19
C165 DIFFPAIR_BIAS.n111 GND 4.95e-19
C166 DIFFPAIR_BIAS.n112 GND 5.25e-19
C167 DIFFPAIR_BIAS.n113 GND 0.001171f
C168 DIFFPAIR_BIAS.n114 GND 0.001171f
C169 DIFFPAIR_BIAS.n115 GND 5.25e-19
C170 DIFFPAIR_BIAS.n116 GND 4.95e-19
C171 DIFFPAIR_BIAS.n117 GND 9.22e-19
C172 DIFFPAIR_BIAS.n118 GND 9.22e-19
C173 DIFFPAIR_BIAS.n119 GND 4.95e-19
C174 DIFFPAIR_BIAS.n120 GND 5.25e-19
C175 DIFFPAIR_BIAS.n121 GND 0.001171f
C176 DIFFPAIR_BIAS.n122 GND 0.002535f
C177 DIFFPAIR_BIAS.n123 GND 5.25e-19
C178 DIFFPAIR_BIAS.n124 GND 4.95e-19
C179 DIFFPAIR_BIAS.n125 GND 0.002131f
C180 DIFFPAIR_BIAS.n126 GND 0.00491f
C181 DIFFPAIR_BIAS.n127 GND 0.08013f
C182 DIFFPAIR_BIAS.t6 GND 0.102337f
C183 DIFFPAIR_BIAS.t4 GND 0.102337f
C184 DIFFPAIR_BIAS.t2 GND 0.102337f
C185 DIFFPAIR_BIAS.t0 GND 0.103205f
C186 DIFFPAIR_BIAS.n128 GND 0.127236f
C187 DIFFPAIR_BIAS.n129 GND 0.068439f
C188 DIFFPAIR_BIAS.n130 GND 0.07541f
C189 DIFFPAIR_BIAS.n131 GND 0.155794f
C190 DIFFPAIR_BIAS.t11 GND 0.108432f
C191 DIFFPAIR_BIAS.n132 GND 0.063754f
C192 DIFFPAIR_BIAS.t10 GND 0.108432f
C193 DIFFPAIR_BIAS.n133 GND 0.061519f
C194 DIFFPAIR_BIAS.n134 GND 0.040079f
C195 VP.n0 GND 0.037196f
C196 VP.t6 GND 0.442682f
C197 VP.n1 GND 0.022514f
C198 VP.t11 GND 0.502376f
C199 VP.n2 GND 0.221655f
C200 VP.t10 GND 0.442682f
C201 VP.n3 GND 0.206565f
C202 VP.n4 GND 0.038013f
C203 VP.n5 GND 0.119334f
C204 VP.n6 GND 0.027876f
C205 VP.n7 GND 0.027876f
C206 VP.n8 GND 0.038013f
C207 VP.n9 GND 0.18176f
C208 VP.n10 GND 0.038235f
C209 VP.t5 GND 0.485128f
C210 VP.n11 GND 0.224883f
C211 VP.n12 GND 0.333286f
C212 VP.n13 GND 0.037196f
C213 VP.t7 GND 0.485128f
C214 VP.t12 GND 0.442682f
C215 VP.n14 GND 0.022514f
C216 VP.t9 GND 0.502376f
C217 VP.n15 GND 0.221655f
C218 VP.t8 GND 0.442682f
C219 VP.n16 GND 0.206565f
C220 VP.n17 GND 0.038013f
C221 VP.n18 GND 0.119335f
C222 VP.n19 GND 0.027876f
C223 VP.n20 GND 0.027876f
C224 VP.n21 GND 0.038013f
C225 VP.n22 GND 0.18176f
C226 VP.n23 GND 0.038235f
C227 VP.n24 GND 0.224883f
C228 VP.n25 GND 0.737721f
C229 VP.n26 GND 1.10137f
C230 VP.t4 GND 0.008593f
C231 VP.t1 GND 0.008593f
C232 VP.n27 GND 0.028257f
C233 VP.t0 GND 0.008593f
C234 VP.t2 GND 0.008593f
C235 VP.n28 GND 0.027869f
C236 VP.n29 GND 0.237852f
C237 VP.t3 GND 0.047829f
C238 VP.n30 GND 0.129794f
C239 VP.n31 GND 1.74358f
C240 a_n2511_10256.n0 GND 1.36544f
C241 a_n2511_10256.t4 GND 0.789396f
C242 a_n2511_10256.t1 GND 0.097661f
C243 a_n2511_10256.t3 GND 0.097661f
C244 a_n2511_10256.n1 GND 0.568406f
C245 a_n2511_10256.n2 GND 1.41612f
C246 a_n2511_10256.t8 GND 0.097661f
C247 a_n2511_10256.t12 GND 0.097661f
C248 a_n2511_10256.n3 GND 0.67573f
C249 a_n2511_10256.t13 GND 0.097661f
C250 a_n2511_10256.t10 GND 0.097661f
C251 a_n2511_10256.n4 GND 0.67218f
C252 a_n2511_10256.n5 GND 2.33544f
C253 a_n2511_10256.t14 GND 0.097661f
C254 a_n2511_10256.t15 GND 0.097661f
C255 a_n2511_10256.n6 GND 0.674733f
C256 a_n2511_10256.t9 GND 0.097661f
C257 a_n2511_10256.t11 GND 0.097661f
C258 a_n2511_10256.n7 GND 0.672183f
C259 a_n2511_10256.n8 GND 5.00954f
C260 a_n2511_10256.n9 GND 1.93174f
C261 a_n2511_10256.t5 GND 0.785576f
C262 a_n2511_10256.n10 GND 1.12527f
C263 a_n2511_10256.t6 GND 0.097661f
C264 a_n2511_10256.t0 GND 0.097661f
C265 a_n2511_10256.n11 GND 0.568406f
C266 a_n2511_10256.n12 GND 0.766742f
C267 a_n2511_10256.t2 GND 0.785576f
C268 a_n2511_10256.t7 GND 0.785576f
C269 a_n2433_10060.n0 GND 1.19248f
C270 a_n2433_10060.n1 GND 0.047166f
C271 a_n2433_10060.n2 GND 1.05335f
C272 a_n2433_10060.n3 GND 0.047166f
C273 a_n2433_10060.n4 GND 1.09055f
C274 a_n2433_10060.n5 GND 0.047166f
C275 a_n2433_10060.n6 GND 0.970179f
C276 a_n2433_10060.n7 GND 0.047166f
C277 a_n2433_10060.n8 GND 0.281203f
C278 a_n2433_10060.n9 GND 0.868055f
C279 a_n2433_10060.n10 GND 0.047166f
C280 a_n2433_10060.n11 GND 1.21315f
C281 a_n2433_10060.n12 GND 3.19451f
C282 a_n2433_10060.n13 GND 0.580374f
C283 a_n2433_10060.n14 GND 2.13457f
C284 a_n2433_10060.n15 GND 2.05918f
C285 a_n2433_10060.n16 GND 5.25575f
C286 a_n2433_10060.n17 GND 0.344956f
C287 a_n2433_10060.n18 GND 0.344956f
C288 a_n2433_10060.n19 GND 0.344956f
C289 a_n2433_10060.n20 GND 0.731826f
C290 a_n2433_10060.n21 GND 0.344956f
C291 a_n2433_10060.n22 GND 0.344956f
C292 a_n2433_10060.n23 GND 0.344956f
C293 a_n2433_10060.n24 GND 0.344956f
C294 a_n2433_10060.n25 GND 0.344956f
C295 a_n2433_10060.n26 GND 0.344956f
C296 a_n2433_10060.n27 GND 0.344956f
C297 a_n2433_10060.n28 GND 0.344956f
C298 a_n2433_10060.n29 GND 0.344956f
C299 a_n2433_10060.n30 GND 0.344956f
C300 a_n2433_10060.n31 GND 0.383328f
C301 a_n2433_10060.n32 GND 0.344956f
C302 a_n2433_10060.n33 GND 0.344956f
C303 a_n2433_10060.n34 GND 0.344956f
C304 a_n2433_10060.n35 GND 0.079506f
C305 a_n2433_10060.n36 GND 0.048465f
C306 a_n2433_10060.n37 GND 0.079506f
C307 a_n2433_10060.n38 GND 0.048465f
C308 a_n2433_10060.n39 GND 0.048465f
C309 a_n2433_10060.t37 GND 0.750708f
C310 a_n2433_10060.t42 GND 0.645011f
C311 a_n2433_10060.t41 GND 0.645011f
C312 a_n2433_10060.t32 GND 0.750708f
C313 a_n2433_10060.t20 GND 0.614465f
C314 a_n2433_10060.t16 GND 0.076019f
C315 a_n2433_10060.t18 GND 0.076019f
C316 a_n2433_10060.n40 GND 0.442447f
C317 a_n2433_10060.t12 GND 0.611488f
C318 a_n2433_10060.t40 GND 0.645011f
C319 a_n2433_10060.t25 GND 0.645011f
C320 a_n2433_10060.t36 GND 0.750708f
C321 a_n2433_10060.t35 GND 0.645011f
C322 a_n2433_10060.t38 GND 0.645011f
C323 a_n2433_10060.t29 GND 0.750708f
C324 a_n2433_10060.t34 GND 0.645011f
C325 a_n2433_10060.t31 GND 0.645011f
C326 a_n2433_10060.t44 GND 0.750708f
C327 a_n2433_10060.t45 GND 0.645011f
C328 a_n2433_10060.t33 GND 0.645011f
C329 a_n2433_10060.t46 GND 0.750708f
C330 a_n2433_10060.t39 GND 0.750708f
C331 a_n2433_10060.t47 GND 0.645011f
C332 a_n2433_10060.t30 GND 0.645011f
C333 a_n2433_10060.t43 GND 0.750708f
C334 a_n2433_10060.t19 GND 0.750708f
C335 a_n2433_10060.t15 GND 0.645011f
C336 a_n2433_10060.t17 GND 0.645011f
C337 a_n2433_10060.t11 GND 0.750708f
C338 a_n2433_10060.n41 GND 0.383003f
C339 a_n2433_10060.n42 GND 0.383003f
C340 a_n2433_10060.n43 GND 0.383003f
C341 a_n2433_10060.n44 GND 0.383003f
C342 a_n2433_10060.t7 GND 0.750708f
C343 a_n2433_10060.t9 GND 0.645011f
C344 a_n2433_10060.t21 GND 0.645011f
C345 a_n2433_10060.t13 GND 0.750708f
C346 a_n2433_10060.n45 GND 0.319413f
C347 a_n2433_10060.n46 GND 0.079506f
C348 a_n2433_10060.n47 GND 0.365787f
C349 a_n2433_10060.t14 GND 0.614465f
C350 a_n2433_10060.t10 GND 0.076019f
C351 a_n2433_10060.t22 GND 0.076019f
C352 a_n2433_10060.n48 GND 0.442447f
C353 a_n2433_10060.t8 GND 0.611491f
C354 a_n2433_10060.n49 GND 0.383003f
C355 a_n2433_10060.n50 GND 0.383003f
C356 a_n2433_10060.t27 GND 0.750708f
C357 a_n2433_10060.n51 GND 0.365787f
C358 a_n2433_10060.n52 GND 0.319413f
C359 a_n2433_10060.t26 GND 0.750708f
C360 a_n2433_10060.n53 GND 0.383003f
C361 a_n2433_10060.n54 GND 0.383003f
C362 a_n2433_10060.t24 GND 0.750708f
C363 a_n2433_10060.n55 GND 0.365787f
C364 a_n2433_10060.n56 GND 0.319413f
C365 a_n2433_10060.t28 GND 0.750708f
C366 a_n2433_10060.n57 GND 0.864586f
C367 a_n2433_10060.n58 GND 0.383003f
C368 a_n2433_10060.n59 GND 0.383003f
C369 a_n2433_10060.t1 GND 0.091223f
C370 a_n2433_10060.t4 GND 0.091223f
C371 a_n2433_10060.n60 GND 0.797966f
C372 a_n2433_10060.t5 GND 0.091223f
C373 a_n2433_10060.t6 GND 0.091223f
C374 a_n2433_10060.n61 GND 0.79669f
C375 a_n2433_10060.t2 GND 0.091223f
C376 a_n2433_10060.t3 GND 0.091223f
C377 a_n2433_10060.n62 GND 0.797963f
C378 a_n2433_10060.n63 GND 2.30949f
C379 a_n2433_10060.t23 GND 0.091223f
C380 a_n2433_10060.n64 GND 0.797963f
C381 a_n2433_10060.t0 GND 0.091223f
C382 a_n1455_n3628.n0 GND 0.029433f
C383 a_n1455_n3628.n1 GND 0.029433f
C384 a_n1455_n3628.n2 GND 0.364885f
C385 a_n1455_n3628.n3 GND 0.029433f
C386 a_n1455_n3628.n4 GND 0.029433f
C387 a_n1455_n3628.n5 GND 0.364885f
C388 a_n1455_n3628.n6 GND 0.029433f
C389 a_n1455_n3628.n7 GND 0.029433f
C390 a_n1455_n3628.n8 GND 0.364885f
C391 a_n1455_n3628.n9 GND 0.029433f
C392 a_n1455_n3628.n10 GND 0.029433f
C393 a_n1455_n3628.n11 GND 0.364885f
C394 a_n1455_n3628.n12 GND 0.029433f
C395 a_n1455_n3628.n13 GND 0.029433f
C396 a_n1455_n3628.n14 GND 0.364885f
C397 a_n1455_n3628.n15 GND 0.029433f
C398 a_n1455_n3628.n16 GND 0.029433f
C399 a_n1455_n3628.n17 GND 0.364885f
C400 a_n1455_n3628.n18 GND 0.029433f
C401 a_n1455_n3628.n19 GND 0.029433f
C402 a_n1455_n3628.n20 GND 0.364885f
C403 a_n1455_n3628.n21 GND 0.029433f
C404 a_n1455_n3628.n22 GND 0.029433f
C405 a_n1455_n3628.n23 GND 0.364885f
C406 a_n1455_n3628.n24 GND 0.350169f
C407 a_n1455_n3628.n25 GND 0.029433f
C408 a_n1455_n3628.n26 GND 0.048734f
C409 a_n1455_n3628.n27 GND 0.029433f
C410 a_n1455_n3628.n28 GND 0.350169f
C411 a_n1455_n3628.n29 GND 0.029433f
C412 a_n1455_n3628.n30 GND 0.048734f
C413 a_n1455_n3628.n31 GND 0.029433f
C414 a_n1455_n3628.n32 GND 0.350169f
C415 a_n1455_n3628.n33 GND 0.029433f
C416 a_n1455_n3628.n34 GND 0.048734f
C417 a_n1455_n3628.n35 GND 0.029433f
C418 a_n1455_n3628.n36 GND 0.350169f
C419 a_n1455_n3628.n37 GND 0.029433f
C420 a_n1455_n3628.n38 GND 0.048734f
C421 a_n1455_n3628.n39 GND 0.029433f
C422 a_n1455_n3628.n40 GND 0.020686f
C423 a_n1455_n3628.n41 GND 0.007908f
C424 a_n1455_n3628.n42 GND 0.018692f
C425 a_n1455_n3628.n43 GND 0.008373f
C426 a_n1455_n3628.n44 GND 0.007908f
C427 a_n1455_n3628.n45 GND 0.018692f
C428 a_n1455_n3628.n46 GND 0.008373f
C429 a_n1455_n3628.n47 GND 0.062977f
C430 a_n1455_n3628.t17 GND 0.030465f
C431 a_n1455_n3628.n48 GND 0.014019f
C432 a_n1455_n3628.n49 GND 0.011041f
C433 a_n1455_n3628.n50 GND 0.007908f
C434 a_n1455_n3628.n51 GND 0.007908f
C435 a_n1455_n3628.n52 GND 0.008373f
C436 a_n1455_n3628.n53 GND 0.018692f
C437 a_n1455_n3628.n54 GND 0.018692f
C438 a_n1455_n3628.n55 GND 0.008373f
C439 a_n1455_n3628.n56 GND 0.007908f
C440 a_n1455_n3628.n57 GND 0.007908f
C441 a_n1455_n3628.n58 GND 0.008373f
C442 a_n1455_n3628.n59 GND 0.018692f
C443 a_n1455_n3628.n60 GND 0.040465f
C444 a_n1455_n3628.n61 GND 0.008373f
C445 a_n1455_n3628.n62 GND 0.007908f
C446 a_n1455_n3628.n63 GND 0.034017f
C447 a_n1455_n3628.n64 GND 0.026084f
C448 a_n1455_n3628.n65 GND 0.16917f
C449 a_n1455_n3628.n66 GND 0.020686f
C450 a_n1455_n3628.n67 GND 0.007908f
C451 a_n1455_n3628.n68 GND 0.018692f
C452 a_n1455_n3628.n69 GND 0.008373f
C453 a_n1455_n3628.n70 GND 0.007908f
C454 a_n1455_n3628.n71 GND 0.018692f
C455 a_n1455_n3628.n72 GND 0.008373f
C456 a_n1455_n3628.n73 GND 0.062977f
C457 a_n1455_n3628.t8 GND 0.030465f
C458 a_n1455_n3628.n74 GND 0.014019f
C459 a_n1455_n3628.n75 GND 0.011041f
C460 a_n1455_n3628.n76 GND 0.007908f
C461 a_n1455_n3628.n77 GND 0.007908f
C462 a_n1455_n3628.n78 GND 0.008373f
C463 a_n1455_n3628.n79 GND 0.018692f
C464 a_n1455_n3628.n80 GND 0.018692f
C465 a_n1455_n3628.n81 GND 0.008373f
C466 a_n1455_n3628.n82 GND 0.007908f
C467 a_n1455_n3628.n83 GND 0.007908f
C468 a_n1455_n3628.n84 GND 0.008373f
C469 a_n1455_n3628.n85 GND 0.018692f
C470 a_n1455_n3628.n86 GND 0.040465f
C471 a_n1455_n3628.n87 GND 0.008373f
C472 a_n1455_n3628.n88 GND 0.007908f
C473 a_n1455_n3628.n89 GND 0.034017f
C474 a_n1455_n3628.n90 GND 0.121814f
C475 a_n1455_n3628.n91 GND 1.26754f
C476 a_n1455_n3628.n92 GND 0.020686f
C477 a_n1455_n3628.n93 GND 0.007908f
C478 a_n1455_n3628.n94 GND 0.018692f
C479 a_n1455_n3628.n95 GND 0.008373f
C480 a_n1455_n3628.n96 GND 0.007908f
C481 a_n1455_n3628.n97 GND 0.018692f
C482 a_n1455_n3628.n98 GND 0.008373f
C483 a_n1455_n3628.n99 GND 0.062977f
C484 a_n1455_n3628.t6 GND 0.030465f
C485 a_n1455_n3628.n100 GND 0.014019f
C486 a_n1455_n3628.n101 GND 0.011041f
C487 a_n1455_n3628.n102 GND 0.007908f
C488 a_n1455_n3628.n103 GND 0.007908f
C489 a_n1455_n3628.n104 GND 0.008373f
C490 a_n1455_n3628.n105 GND 0.018692f
C491 a_n1455_n3628.n106 GND 0.018692f
C492 a_n1455_n3628.n107 GND 0.008373f
C493 a_n1455_n3628.n108 GND 0.007908f
C494 a_n1455_n3628.n109 GND 0.007908f
C495 a_n1455_n3628.n110 GND 0.008373f
C496 a_n1455_n3628.n111 GND 0.018692f
C497 a_n1455_n3628.n112 GND 0.040465f
C498 a_n1455_n3628.n113 GND 0.008373f
C499 a_n1455_n3628.n114 GND 0.007908f
C500 a_n1455_n3628.n115 GND 0.034017f
C501 a_n1455_n3628.n116 GND 0.026084f
C502 a_n1455_n3628.n117 GND 0.16917f
C503 a_n1455_n3628.t10 GND 0.069777f
C504 a_n1455_n3628.t2 GND 0.069777f
C505 a_n1455_n3628.n118 GND 0.558312f
C506 a_n1455_n3628.n119 GND 0.347298f
C507 a_n1455_n3628.n120 GND 0.020686f
C508 a_n1455_n3628.n121 GND 0.007908f
C509 a_n1455_n3628.n122 GND 0.018692f
C510 a_n1455_n3628.n123 GND 0.008373f
C511 a_n1455_n3628.n124 GND 0.007908f
C512 a_n1455_n3628.n125 GND 0.018692f
C513 a_n1455_n3628.n126 GND 0.008373f
C514 a_n1455_n3628.n127 GND 0.062977f
C515 a_n1455_n3628.t9 GND 0.030465f
C516 a_n1455_n3628.n128 GND 0.014019f
C517 a_n1455_n3628.n129 GND 0.011041f
C518 a_n1455_n3628.n130 GND 0.007908f
C519 a_n1455_n3628.n131 GND 0.007908f
C520 a_n1455_n3628.n132 GND 0.008373f
C521 a_n1455_n3628.n133 GND 0.018692f
C522 a_n1455_n3628.n134 GND 0.018692f
C523 a_n1455_n3628.n135 GND 0.008373f
C524 a_n1455_n3628.n136 GND 0.007908f
C525 a_n1455_n3628.n137 GND 0.007908f
C526 a_n1455_n3628.n138 GND 0.008373f
C527 a_n1455_n3628.n139 GND 0.018692f
C528 a_n1455_n3628.n140 GND 0.040465f
C529 a_n1455_n3628.n141 GND 0.008373f
C530 a_n1455_n3628.n142 GND 0.007908f
C531 a_n1455_n3628.n143 GND 0.034017f
C532 a_n1455_n3628.n144 GND 0.026084f
C533 a_n1455_n3628.n145 GND 0.610154f
C534 a_n1455_n3628.n146 GND 0.020686f
C535 a_n1455_n3628.n147 GND 0.007908f
C536 a_n1455_n3628.n148 GND 0.018692f
C537 a_n1455_n3628.n149 GND 0.008373f
C538 a_n1455_n3628.n150 GND 0.007908f
C539 a_n1455_n3628.n151 GND 0.018692f
C540 a_n1455_n3628.n152 GND 0.008373f
C541 a_n1455_n3628.n153 GND 0.062977f
C542 a_n1455_n3628.t0 GND 0.030465f
C543 a_n1455_n3628.n154 GND 0.014019f
C544 a_n1455_n3628.n155 GND 0.011041f
C545 a_n1455_n3628.n156 GND 0.007908f
C546 a_n1455_n3628.n157 GND 0.007908f
C547 a_n1455_n3628.n158 GND 0.008373f
C548 a_n1455_n3628.n159 GND 0.018692f
C549 a_n1455_n3628.n160 GND 0.018692f
C550 a_n1455_n3628.n161 GND 0.008373f
C551 a_n1455_n3628.n162 GND 0.007908f
C552 a_n1455_n3628.n163 GND 0.007908f
C553 a_n1455_n3628.n164 GND 0.008373f
C554 a_n1455_n3628.n165 GND 0.018692f
C555 a_n1455_n3628.n166 GND 0.040465f
C556 a_n1455_n3628.n167 GND 0.008373f
C557 a_n1455_n3628.n168 GND 0.007908f
C558 a_n1455_n3628.n169 GND 0.034017f
C559 a_n1455_n3628.n170 GND 0.122845f
C560 a_n1455_n3628.n171 GND 0.020686f
C561 a_n1455_n3628.n172 GND 0.007908f
C562 a_n1455_n3628.n173 GND 0.018692f
C563 a_n1455_n3628.n174 GND 0.008373f
C564 a_n1455_n3628.n175 GND 0.007908f
C565 a_n1455_n3628.n176 GND 0.018692f
C566 a_n1455_n3628.n177 GND 0.008373f
C567 a_n1455_n3628.n178 GND 0.062977f
C568 a_n1455_n3628.t5 GND 0.030465f
C569 a_n1455_n3628.n179 GND 0.014019f
C570 a_n1455_n3628.n180 GND 0.011041f
C571 a_n1455_n3628.n181 GND 0.007908f
C572 a_n1455_n3628.n182 GND 0.007908f
C573 a_n1455_n3628.n183 GND 0.008373f
C574 a_n1455_n3628.n184 GND 0.018692f
C575 a_n1455_n3628.n185 GND 0.018692f
C576 a_n1455_n3628.n186 GND 0.008373f
C577 a_n1455_n3628.n187 GND 0.007908f
C578 a_n1455_n3628.n188 GND 0.007908f
C579 a_n1455_n3628.n189 GND 0.008373f
C580 a_n1455_n3628.n190 GND 0.018692f
C581 a_n1455_n3628.n191 GND 0.040465f
C582 a_n1455_n3628.n192 GND 0.008373f
C583 a_n1455_n3628.n193 GND 0.007908f
C584 a_n1455_n3628.n194 GND 0.034017f
C585 a_n1455_n3628.n195 GND 0.121814f
C586 a_n1455_n3628.n196 GND 0.933421f
C587 a_n1455_n3628.n197 GND 0.020686f
C588 a_n1455_n3628.n198 GND 0.007908f
C589 a_n1455_n3628.n199 GND 0.018692f
C590 a_n1455_n3628.n200 GND 0.008373f
C591 a_n1455_n3628.n201 GND 0.007908f
C592 a_n1455_n3628.n202 GND 0.018692f
C593 a_n1455_n3628.n203 GND 0.008373f
C594 a_n1455_n3628.n204 GND 0.062977f
C595 a_n1455_n3628.t7 GND 0.030465f
C596 a_n1455_n3628.n205 GND 0.014019f
C597 a_n1455_n3628.n206 GND 0.011041f
C598 a_n1455_n3628.n207 GND 0.007908f
C599 a_n1455_n3628.n208 GND 0.007908f
C600 a_n1455_n3628.n209 GND 0.008373f
C601 a_n1455_n3628.n210 GND 0.018692f
C602 a_n1455_n3628.n211 GND 0.018692f
C603 a_n1455_n3628.n212 GND 0.008373f
C604 a_n1455_n3628.n213 GND 0.007908f
C605 a_n1455_n3628.n214 GND 0.007908f
C606 a_n1455_n3628.n215 GND 0.008373f
C607 a_n1455_n3628.n216 GND 0.018692f
C608 a_n1455_n3628.n217 GND 0.040465f
C609 a_n1455_n3628.n218 GND 0.008373f
C610 a_n1455_n3628.n219 GND 0.007908f
C611 a_n1455_n3628.n220 GND 0.034017f
C612 a_n1455_n3628.n221 GND 0.121814f
C613 a_n1455_n3628.n222 GND 0.708238f
C614 a_n1455_n3628.n223 GND 0.89644f
C615 a_n1455_n3628.n224 GND 0.714807f
C616 a_n1455_n3628.n225 GND 0.020686f
C617 a_n1455_n3628.n226 GND 0.007908f
C618 a_n1455_n3628.n227 GND 0.018692f
C619 a_n1455_n3628.n228 GND 0.008373f
C620 a_n1455_n3628.n229 GND 0.007908f
C621 a_n1455_n3628.n230 GND 0.018692f
C622 a_n1455_n3628.n231 GND 0.008373f
C623 a_n1455_n3628.n232 GND 0.062977f
C624 a_n1455_n3628.t15 GND 0.030465f
C625 a_n1455_n3628.n233 GND 0.014019f
C626 a_n1455_n3628.n234 GND 0.011041f
C627 a_n1455_n3628.n235 GND 0.007908f
C628 a_n1455_n3628.n236 GND 0.007908f
C629 a_n1455_n3628.n237 GND 0.008373f
C630 a_n1455_n3628.n238 GND 0.018692f
C631 a_n1455_n3628.n239 GND 0.018692f
C632 a_n1455_n3628.n240 GND 0.008373f
C633 a_n1455_n3628.n241 GND 0.007908f
C634 a_n1455_n3628.n242 GND 0.007908f
C635 a_n1455_n3628.n243 GND 0.008373f
C636 a_n1455_n3628.n244 GND 0.018692f
C637 a_n1455_n3628.n245 GND 0.040465f
C638 a_n1455_n3628.n246 GND 0.008373f
C639 a_n1455_n3628.n247 GND 0.007908f
C640 a_n1455_n3628.n248 GND 0.026084f
C641 a_n1455_n3628.n249 GND 0.381969f
C642 a_n1455_n3628.t16 GND 0.069777f
C643 a_n1455_n3628.t12 GND 0.069777f
C644 a_n1455_n3628.n250 GND 0.558309f
C645 a_n1455_n3628.n251 GND 0.347302f
C646 a_n1455_n3628.n252 GND 0.020686f
C647 a_n1455_n3628.n253 GND 0.007908f
C648 a_n1455_n3628.n254 GND 0.018692f
C649 a_n1455_n3628.n255 GND 0.008373f
C650 a_n1455_n3628.n256 GND 0.007908f
C651 a_n1455_n3628.n257 GND 0.018692f
C652 a_n1455_n3628.n258 GND 0.008373f
C653 a_n1455_n3628.n259 GND 0.062977f
C654 a_n1455_n3628.t19 GND 0.030465f
C655 a_n1455_n3628.n260 GND 0.014019f
C656 a_n1455_n3628.n261 GND 0.011041f
C657 a_n1455_n3628.n262 GND 0.007908f
C658 a_n1455_n3628.n263 GND 0.007908f
C659 a_n1455_n3628.n264 GND 0.008373f
C660 a_n1455_n3628.n265 GND 0.018692f
C661 a_n1455_n3628.n266 GND 0.018692f
C662 a_n1455_n3628.n267 GND 0.008373f
C663 a_n1455_n3628.n268 GND 0.007908f
C664 a_n1455_n3628.n269 GND 0.007908f
C665 a_n1455_n3628.n270 GND 0.008373f
C666 a_n1455_n3628.n271 GND 0.018692f
C667 a_n1455_n3628.n272 GND 0.040465f
C668 a_n1455_n3628.n273 GND 0.008373f
C669 a_n1455_n3628.n274 GND 0.007908f
C670 a_n1455_n3628.n275 GND 0.026084f
C671 a_n1455_n3628.n276 GND 0.16917f
C672 a_n1455_n3628.n277 GND 0.020686f
C673 a_n1455_n3628.n278 GND 0.007908f
C674 a_n1455_n3628.n279 GND 0.018692f
C675 a_n1455_n3628.n280 GND 0.008373f
C676 a_n1455_n3628.n281 GND 0.007908f
C677 a_n1455_n3628.n282 GND 0.018692f
C678 a_n1455_n3628.n283 GND 0.008373f
C679 a_n1455_n3628.n284 GND 0.062977f
C680 a_n1455_n3628.t1 GND 0.030465f
C681 a_n1455_n3628.n285 GND 0.014019f
C682 a_n1455_n3628.n286 GND 0.011041f
C683 a_n1455_n3628.n287 GND 0.007908f
C684 a_n1455_n3628.n288 GND 0.007908f
C685 a_n1455_n3628.n289 GND 0.008373f
C686 a_n1455_n3628.n290 GND 0.018692f
C687 a_n1455_n3628.n291 GND 0.018692f
C688 a_n1455_n3628.n292 GND 0.008373f
C689 a_n1455_n3628.n293 GND 0.007908f
C690 a_n1455_n3628.n294 GND 0.007908f
C691 a_n1455_n3628.n295 GND 0.008373f
C692 a_n1455_n3628.n296 GND 0.018692f
C693 a_n1455_n3628.n297 GND 0.040465f
C694 a_n1455_n3628.n298 GND 0.008373f
C695 a_n1455_n3628.n299 GND 0.007908f
C696 a_n1455_n3628.n300 GND 0.026084f
C697 a_n1455_n3628.n301 GND 0.16917f
C698 a_n1455_n3628.t11 GND 0.069777f
C699 a_n1455_n3628.t3 GND 0.069777f
C700 a_n1455_n3628.n302 GND 0.558309f
C701 a_n1455_n3628.n303 GND 0.347302f
C702 a_n1455_n3628.n304 GND 0.020686f
C703 a_n1455_n3628.n305 GND 0.007908f
C704 a_n1455_n3628.n306 GND 0.018692f
C705 a_n1455_n3628.n307 GND 0.008373f
C706 a_n1455_n3628.n308 GND 0.007908f
C707 a_n1455_n3628.n309 GND 0.018692f
C708 a_n1455_n3628.n310 GND 0.008373f
C709 a_n1455_n3628.n311 GND 0.062977f
C710 a_n1455_n3628.t4 GND 0.030465f
C711 a_n1455_n3628.n312 GND 0.014019f
C712 a_n1455_n3628.n313 GND 0.011041f
C713 a_n1455_n3628.n314 GND 0.007908f
C714 a_n1455_n3628.n315 GND 0.007908f
C715 a_n1455_n3628.n316 GND 0.008373f
C716 a_n1455_n3628.n317 GND 0.018692f
C717 a_n1455_n3628.n318 GND 0.018692f
C718 a_n1455_n3628.n319 GND 0.008373f
C719 a_n1455_n3628.n320 GND 0.007908f
C720 a_n1455_n3628.n321 GND 0.007908f
C721 a_n1455_n3628.n322 GND 0.008373f
C722 a_n1455_n3628.n323 GND 0.018692f
C723 a_n1455_n3628.n324 GND 0.040465f
C724 a_n1455_n3628.n325 GND 0.008373f
C725 a_n1455_n3628.n326 GND 0.007908f
C726 a_n1455_n3628.n327 GND 0.026084f
C727 a_n1455_n3628.n328 GND 0.381969f
C728 a_n1455_n3628.n329 GND 0.80329f
C729 a_n1455_n3628.n330 GND 0.020686f
C730 a_n1455_n3628.n331 GND 0.007908f
C731 a_n1455_n3628.n332 GND 0.018692f
C732 a_n1455_n3628.n333 GND 0.008373f
C733 a_n1455_n3628.n334 GND 0.007908f
C734 a_n1455_n3628.n335 GND 0.018692f
C735 a_n1455_n3628.n336 GND 0.008373f
C736 a_n1455_n3628.n337 GND 0.062977f
C737 a_n1455_n3628.t14 GND 0.030465f
C738 a_n1455_n3628.n338 GND 0.014019f
C739 a_n1455_n3628.n339 GND 0.011041f
C740 a_n1455_n3628.n340 GND 0.007908f
C741 a_n1455_n3628.n341 GND 0.007908f
C742 a_n1455_n3628.n342 GND 0.008373f
C743 a_n1455_n3628.n343 GND 0.018692f
C744 a_n1455_n3628.n344 GND 0.018692f
C745 a_n1455_n3628.n345 GND 0.008373f
C746 a_n1455_n3628.n346 GND 0.007908f
C747 a_n1455_n3628.n347 GND 0.007908f
C748 a_n1455_n3628.n348 GND 0.008373f
C749 a_n1455_n3628.n349 GND 0.018692f
C750 a_n1455_n3628.n350 GND 0.040465f
C751 a_n1455_n3628.n351 GND 0.008373f
C752 a_n1455_n3628.n352 GND 0.007908f
C753 a_n1455_n3628.n353 GND 0.034017f
C754 a_n1455_n3628.n354 GND 0.026084f
C755 a_n1455_n3628.n355 GND 0.610154f
C756 a_n1455_n3628.n356 GND 0.347298f
C757 a_n1455_n3628.t13 GND 0.069777f
C758 a_n1455_n3628.n357 GND 0.558312f
C759 a_n1455_n3628.t18 GND 0.069777f
C760 VN.n0 GND 0.026025f
C761 VN.t9 GND 0.339432f
C762 VN.t8 GND 0.309734f
C763 VN.n1 GND 0.015753f
C764 VN.t5 GND 0.351499f
C765 VN.n2 GND 0.155086f
C766 VN.t12 GND 0.309734f
C767 VN.n3 GND 0.144528f
C768 VN.n4 GND 0.026597f
C769 VN.n5 GND 0.083495f
C770 VN.n6 GND 0.019504f
C771 VN.n7 GND 0.019504f
C772 VN.n8 GND 0.026597f
C773 VN.n9 GND 0.127173f
C774 VN.n10 GND 0.026752f
C775 VN.n11 GND 0.157345f
C776 VN.n12 GND 0.228308f
C777 VN.n13 GND 0.026025f
C778 VN.t11 GND 0.309734f
C779 VN.n14 GND 0.015753f
C780 VN.t7 GND 0.351499f
C781 VN.n15 GND 0.155086f
C782 VN.t6 GND 0.309734f
C783 VN.n16 GND 0.144528f
C784 VN.n17 GND 0.026597f
C785 VN.n18 GND 0.083495f
C786 VN.n19 GND 0.019504f
C787 VN.n20 GND 0.019504f
C788 VN.n21 GND 0.026597f
C789 VN.n22 GND 0.127173f
C790 VN.n23 GND 0.026752f
C791 VN.t10 GND 0.339432f
C792 VN.n24 GND 0.157345f
C793 VN.n25 GND 0.508348f
C794 VN.n26 GND 0.762742f
C795 VN.t0 GND 0.033669f
C796 VN.t1 GND 0.006012f
C797 VN.t4 GND 0.006012f
C798 VN.n27 GND 0.019499f
C799 VN.n28 GND 0.151376f
C800 VN.t2 GND 0.006012f
C801 VN.t3 GND 0.006012f
C802 VN.n29 GND 0.019499f
C803 VN.n30 GND 0.113626f
C804 VN.n31 GND 1.86465f
C805 CS_BIAS.n0 GND 0.007684f
C806 CS_BIAS.t55 GND 0.185122f
C807 CS_BIAS.n1 GND 0.008311f
C808 CS_BIAS.n2 GND 0.005829f
C809 CS_BIAS.t35 GND 0.185122f
C810 CS_BIAS.n3 GND 0.005338f
C811 CS_BIAS.n4 GND 0.005829f
C812 CS_BIAS.t39 GND 0.185122f
C813 CS_BIAS.n5 GND 0.010861f
C814 CS_BIAS.n6 GND 0.005829f
C815 CS_BIAS.t36 GND 0.185122f
C816 CS_BIAS.n7 GND 0.070673f
C817 CS_BIAS.n8 GND 0.005092f
C818 CS_BIAS.n9 GND 0.009901f
C819 CS_BIAS.n10 GND 0.007684f
C820 CS_BIAS.t6 GND 0.185122f
C821 CS_BIAS.n11 GND 0.008311f
C822 CS_BIAS.n12 GND 0.005829f
C823 CS_BIAS.t30 GND 0.185122f
C824 CS_BIAS.n13 GND 0.005338f
C825 CS_BIAS.n14 GND 0.005829f
C826 CS_BIAS.t22 GND 0.185122f
C827 CS_BIAS.n15 GND 0.010861f
C828 CS_BIAS.n16 GND 0.005829f
C829 CS_BIAS.t18 GND 0.185122f
C830 CS_BIAS.n17 GND 0.070673f
C831 CS_BIAS.n18 GND 0.005829f
C832 CS_BIAS.n19 GND 0.009901f
C833 CS_BIAS.n20 GND 0.005829f
C834 CS_BIAS.t0 GND 0.185122f
C835 CS_BIAS.n21 GND 0.070673f
C836 CS_BIAS.n22 GND 0.010861f
C837 CS_BIAS.n23 GND 0.005829f
C838 CS_BIAS.t16 GND 0.185122f
C839 CS_BIAS.n24 GND 0.005338f
C840 CS_BIAS.n25 GND 0.043632f
C841 CS_BIAS.t2 GND 0.185122f
C842 CS_BIAS.t26 GND 0.214423f
C843 CS_BIAS.n26 GND 0.084881f
C844 CS_BIAS.n27 GND 0.082798f
C845 CS_BIAS.n28 GND 0.006273f
C846 CS_BIAS.n29 GND 0.01166f
C847 CS_BIAS.n30 GND 0.005829f
C848 CS_BIAS.n31 GND 0.005829f
C849 CS_BIAS.n32 GND 0.005829f
C850 CS_BIAS.n33 GND 0.010755f
C851 CS_BIAS.n34 GND 0.008194f
C852 CS_BIAS.n35 GND 0.070673f
C853 CS_BIAS.n36 GND 0.008087f
C854 CS_BIAS.n37 GND 0.005829f
C855 CS_BIAS.n38 GND 0.005829f
C856 CS_BIAS.n39 GND 0.005829f
C857 CS_BIAS.n40 GND 0.005201f
C858 CS_BIAS.n41 GND 0.011692f
C859 CS_BIAS.n42 GND 0.00638f
C860 CS_BIAS.n43 GND 0.005829f
C861 CS_BIAS.n44 GND 0.005829f
C862 CS_BIAS.n45 GND 0.005829f
C863 CS_BIAS.n46 GND 0.008473f
C864 CS_BIAS.n47 GND 0.008473f
C865 CS_BIAS.n48 GND 0.009901f
C866 CS_BIAS.n49 GND 0.005829f
C867 CS_BIAS.n50 GND 0.005829f
C868 CS_BIAS.n51 GND 0.00638f
C869 CS_BIAS.n52 GND 0.011692f
C870 CS_BIAS.n53 GND 0.005201f
C871 CS_BIAS.n54 GND 0.005829f
C872 CS_BIAS.n55 GND 0.005829f
C873 CS_BIAS.n56 GND 0.005829f
C874 CS_BIAS.n57 GND 0.008087f
C875 CS_BIAS.n58 GND 0.070673f
C876 CS_BIAS.n59 GND 0.008194f
C877 CS_BIAS.n60 GND 0.010755f
C878 CS_BIAS.n61 GND 0.005829f
C879 CS_BIAS.n62 GND 0.005829f
C880 CS_BIAS.n63 GND 0.005829f
C881 CS_BIAS.n64 GND 0.01166f
C882 CS_BIAS.n65 GND 0.006273f
C883 CS_BIAS.n66 GND 0.070673f
C884 CS_BIAS.n67 GND 0.010008f
C885 CS_BIAS.n68 GND 0.005829f
C886 CS_BIAS.n69 GND 0.005829f
C887 CS_BIAS.n70 GND 0.005829f
C888 CS_BIAS.n71 GND 0.008634f
C889 CS_BIAS.n72 GND 0.009795f
C890 CS_BIAS.n73 GND 0.088447f
C891 CS_BIAS.n74 GND 0.058541f
C892 CS_BIAS.t7 GND 0.010781f
C893 CS_BIAS.t31 GND 0.010781f
C894 CS_BIAS.n75 GND 0.094152f
C895 CS_BIAS.n76 GND 0.1167f
C896 CS_BIAS.t23 GND 0.010781f
C897 CS_BIAS.t19 GND 0.010781f
C898 CS_BIAS.n77 GND 0.094152f
C899 CS_BIAS.n78 GND 0.061488f
C900 CS_BIAS.t3 GND 0.010781f
C901 CS_BIAS.t27 GND 0.010781f
C902 CS_BIAS.n79 GND 0.095073f
C903 CS_BIAS.t1 GND 0.010781f
C904 CS_BIAS.t17 GND 0.010781f
C905 CS_BIAS.n80 GND 0.094152f
C906 CS_BIAS.n81 GND 0.138602f
C907 CS_BIAS.n82 GND 0.064277f
C908 CS_BIAS.n83 GND 0.037722f
C909 CS_BIAS.n84 GND 0.005829f
C910 CS_BIAS.t51 GND 0.185122f
C911 CS_BIAS.n85 GND 0.070673f
C912 CS_BIAS.n86 GND 0.010861f
C913 CS_BIAS.n87 GND 0.005829f
C914 CS_BIAS.t52 GND 0.185122f
C915 CS_BIAS.n88 GND 0.005338f
C916 CS_BIAS.n89 GND 0.043632f
C917 CS_BIAS.t42 GND 0.185122f
C918 CS_BIAS.t44 GND 0.214423f
C919 CS_BIAS.n90 GND 0.084881f
C920 CS_BIAS.n91 GND 0.082798f
C921 CS_BIAS.n92 GND 0.006273f
C922 CS_BIAS.n93 GND 0.01166f
C923 CS_BIAS.n94 GND 0.005829f
C924 CS_BIAS.n95 GND 0.005829f
C925 CS_BIAS.n96 GND 0.005829f
C926 CS_BIAS.n97 GND 0.010755f
C927 CS_BIAS.n98 GND 0.008194f
C928 CS_BIAS.n99 GND 0.070673f
C929 CS_BIAS.n100 GND 0.008087f
C930 CS_BIAS.n101 GND 0.005829f
C931 CS_BIAS.n102 GND 0.005829f
C932 CS_BIAS.n103 GND 0.005829f
C933 CS_BIAS.n104 GND 0.005201f
C934 CS_BIAS.n105 GND 0.011692f
C935 CS_BIAS.n106 GND 0.00638f
C936 CS_BIAS.n107 GND 0.005829f
C937 CS_BIAS.n108 GND 0.005829f
C938 CS_BIAS.n109 GND 0.005092f
C939 CS_BIAS.n110 GND 0.008473f
C940 CS_BIAS.n111 GND 0.008473f
C941 CS_BIAS.n112 GND 0.009901f
C942 CS_BIAS.n113 GND 0.005829f
C943 CS_BIAS.n114 GND 0.005829f
C944 CS_BIAS.n115 GND 0.00638f
C945 CS_BIAS.n116 GND 0.011692f
C946 CS_BIAS.n117 GND 0.005201f
C947 CS_BIAS.n118 GND 0.005829f
C948 CS_BIAS.n119 GND 0.005829f
C949 CS_BIAS.n120 GND 0.005829f
C950 CS_BIAS.n121 GND 0.008087f
C951 CS_BIAS.n122 GND 0.070673f
C952 CS_BIAS.n123 GND 0.008194f
C953 CS_BIAS.n124 GND 0.010755f
C954 CS_BIAS.n125 GND 0.005829f
C955 CS_BIAS.n126 GND 0.005829f
C956 CS_BIAS.n127 GND 0.005829f
C957 CS_BIAS.n128 GND 0.01166f
C958 CS_BIAS.n129 GND 0.006273f
C959 CS_BIAS.n130 GND 0.070673f
C960 CS_BIAS.n131 GND 0.010008f
C961 CS_BIAS.n132 GND 0.005829f
C962 CS_BIAS.n133 GND 0.005829f
C963 CS_BIAS.n134 GND 0.005829f
C964 CS_BIAS.n135 GND 0.008634f
C965 CS_BIAS.n136 GND 0.009795f
C966 CS_BIAS.n137 GND 0.088447f
C967 CS_BIAS.n138 GND 0.035075f
C968 CS_BIAS.n139 GND 0.007684f
C969 CS_BIAS.t48 GND 0.185122f
C970 CS_BIAS.n140 GND 0.008311f
C971 CS_BIAS.n141 GND 0.005829f
C972 CS_BIAS.t61 GND 0.185122f
C973 CS_BIAS.n142 GND 0.005338f
C974 CS_BIAS.n143 GND 0.005829f
C975 CS_BIAS.t63 GND 0.185122f
C976 CS_BIAS.n144 GND 0.010861f
C977 CS_BIAS.n145 GND 0.005829f
C978 CS_BIAS.t62 GND 0.185122f
C979 CS_BIAS.n146 GND 0.070673f
C980 CS_BIAS.n147 GND 0.005829f
C981 CS_BIAS.n148 GND 0.009901f
C982 CS_BIAS.n149 GND 0.005829f
C983 CS_BIAS.t46 GND 0.185122f
C984 CS_BIAS.n150 GND 0.070673f
C985 CS_BIAS.n151 GND 0.010861f
C986 CS_BIAS.n152 GND 0.005829f
C987 CS_BIAS.t47 GND 0.185122f
C988 CS_BIAS.n153 GND 0.005338f
C989 CS_BIAS.n154 GND 0.043632f
C990 CS_BIAS.t37 GND 0.185122f
C991 CS_BIAS.t40 GND 0.214423f
C992 CS_BIAS.n155 GND 0.084881f
C993 CS_BIAS.n156 GND 0.082798f
C994 CS_BIAS.n157 GND 0.006273f
C995 CS_BIAS.n158 GND 0.01166f
C996 CS_BIAS.n159 GND 0.005829f
C997 CS_BIAS.n160 GND 0.005829f
C998 CS_BIAS.n161 GND 0.005829f
C999 CS_BIAS.n162 GND 0.010755f
C1000 CS_BIAS.n163 GND 0.008194f
C1001 CS_BIAS.n164 GND 0.070673f
C1002 CS_BIAS.n165 GND 0.008087f
C1003 CS_BIAS.n166 GND 0.005829f
C1004 CS_BIAS.n167 GND 0.005829f
C1005 CS_BIAS.n168 GND 0.005829f
C1006 CS_BIAS.n169 GND 0.005201f
C1007 CS_BIAS.n170 GND 0.011692f
C1008 CS_BIAS.n171 GND 0.00638f
C1009 CS_BIAS.n172 GND 0.005829f
C1010 CS_BIAS.n173 GND 0.005829f
C1011 CS_BIAS.n174 GND 0.005829f
C1012 CS_BIAS.n175 GND 0.008473f
C1013 CS_BIAS.n176 GND 0.008473f
C1014 CS_BIAS.n177 GND 0.009901f
C1015 CS_BIAS.n178 GND 0.005829f
C1016 CS_BIAS.n179 GND 0.005829f
C1017 CS_BIAS.n180 GND 0.00638f
C1018 CS_BIAS.n181 GND 0.011692f
C1019 CS_BIAS.n182 GND 0.005201f
C1020 CS_BIAS.n183 GND 0.005829f
C1021 CS_BIAS.n184 GND 0.005829f
C1022 CS_BIAS.n185 GND 0.005829f
C1023 CS_BIAS.n186 GND 0.008087f
C1024 CS_BIAS.n187 GND 0.070673f
C1025 CS_BIAS.n188 GND 0.008194f
C1026 CS_BIAS.n189 GND 0.010755f
C1027 CS_BIAS.n190 GND 0.005829f
C1028 CS_BIAS.n191 GND 0.005829f
C1029 CS_BIAS.n192 GND 0.005829f
C1030 CS_BIAS.n193 GND 0.01166f
C1031 CS_BIAS.n194 GND 0.006273f
C1032 CS_BIAS.n195 GND 0.070673f
C1033 CS_BIAS.n196 GND 0.010008f
C1034 CS_BIAS.n197 GND 0.005829f
C1035 CS_BIAS.n198 GND 0.005829f
C1036 CS_BIAS.n199 GND 0.005829f
C1037 CS_BIAS.n200 GND 0.008634f
C1038 CS_BIAS.n201 GND 0.009795f
C1039 CS_BIAS.n202 GND 0.088447f
C1040 CS_BIAS.n203 GND 0.021125f
C1041 CS_BIAS.n204 GND 0.263448f
C1042 CS_BIAS.n205 GND 0.007684f
C1043 CS_BIAS.t33 GND 0.185122f
C1044 CS_BIAS.n206 GND 0.008311f
C1045 CS_BIAS.n207 GND 0.005829f
C1046 CS_BIAS.t58 GND 0.185122f
C1047 CS_BIAS.n208 GND 0.005338f
C1048 CS_BIAS.n209 GND 0.005829f
C1049 CS_BIAS.t49 GND 0.185122f
C1050 CS_BIAS.n210 GND 0.010861f
C1051 CS_BIAS.n211 GND 0.005829f
C1052 CS_BIAS.t57 GND 0.185122f
C1053 CS_BIAS.n212 GND 0.070673f
C1054 CS_BIAS.n213 GND 0.005092f
C1055 CS_BIAS.n214 GND 0.009901f
C1056 CS_BIAS.n215 GND 0.005829f
C1057 CS_BIAS.n216 GND 0.010861f
C1058 CS_BIAS.n217 GND 0.005829f
C1059 CS_BIAS.t43 GND 0.185122f
C1060 CS_BIAS.n218 GND 0.005338f
C1061 CS_BIAS.n219 GND 0.043632f
C1062 CS_BIAS.t32 GND 0.185122f
C1063 CS_BIAS.t56 GND 0.214423f
C1064 CS_BIAS.n220 GND 0.084881f
C1065 CS_BIAS.n221 GND 0.082798f
C1066 CS_BIAS.n222 GND 0.006273f
C1067 CS_BIAS.n223 GND 0.01166f
C1068 CS_BIAS.n224 GND 0.005829f
C1069 CS_BIAS.n225 GND 0.005829f
C1070 CS_BIAS.n226 GND 0.005829f
C1071 CS_BIAS.n227 GND 0.010755f
C1072 CS_BIAS.n228 GND 0.008194f
C1073 CS_BIAS.n229 GND 0.070673f
C1074 CS_BIAS.n230 GND 0.008087f
C1075 CS_BIAS.n231 GND 0.005829f
C1076 CS_BIAS.n232 GND 0.005829f
C1077 CS_BIAS.n233 GND 0.005829f
C1078 CS_BIAS.n234 GND 0.005201f
C1079 CS_BIAS.n235 GND 0.011692f
C1080 CS_BIAS.t41 GND 0.185122f
C1081 CS_BIAS.n236 GND 0.070673f
C1082 CS_BIAS.n237 GND 0.00638f
C1083 CS_BIAS.n238 GND 0.005829f
C1084 CS_BIAS.n239 GND 0.005829f
C1085 CS_BIAS.t25 GND 0.010781f
C1086 CS_BIAS.t15 GND 0.010781f
C1087 CS_BIAS.n240 GND 0.095073f
C1088 CS_BIAS.t21 GND 0.010781f
C1089 CS_BIAS.t13 GND 0.010781f
C1090 CS_BIAS.n241 GND 0.094152f
C1091 CS_BIAS.n242 GND 0.138602f
C1092 CS_BIAS.n243 GND 0.007684f
C1093 CS_BIAS.t28 GND 0.185122f
C1094 CS_BIAS.n244 GND 0.008311f
C1095 CS_BIAS.n245 GND 0.005829f
C1096 CS_BIAS.t4 GND 0.185122f
C1097 CS_BIAS.n246 GND 0.005338f
C1098 CS_BIAS.n247 GND 0.005829f
C1099 CS_BIAS.t10 GND 0.185122f
C1100 CS_BIAS.n248 GND 0.010861f
C1101 CS_BIAS.n249 GND 0.005829f
C1102 CS_BIAS.t8 GND 0.185122f
C1103 CS_BIAS.n250 GND 0.070673f
C1104 CS_BIAS.n251 GND 0.005829f
C1105 CS_BIAS.n252 GND 0.009901f
C1106 CS_BIAS.n253 GND 0.005829f
C1107 CS_BIAS.n254 GND 0.010861f
C1108 CS_BIAS.n255 GND 0.005829f
C1109 CS_BIAS.t20 GND 0.185122f
C1110 CS_BIAS.n256 GND 0.005338f
C1111 CS_BIAS.n257 GND 0.043632f
C1112 CS_BIAS.t14 GND 0.185122f
C1113 CS_BIAS.t24 GND 0.214423f
C1114 CS_BIAS.n258 GND 0.084881f
C1115 CS_BIAS.n259 GND 0.082798f
C1116 CS_BIAS.n260 GND 0.006273f
C1117 CS_BIAS.n261 GND 0.01166f
C1118 CS_BIAS.n262 GND 0.005829f
C1119 CS_BIAS.n263 GND 0.005829f
C1120 CS_BIAS.n264 GND 0.005829f
C1121 CS_BIAS.n265 GND 0.010755f
C1122 CS_BIAS.n266 GND 0.008194f
C1123 CS_BIAS.n267 GND 0.070673f
C1124 CS_BIAS.n268 GND 0.008087f
C1125 CS_BIAS.n269 GND 0.005829f
C1126 CS_BIAS.n270 GND 0.005829f
C1127 CS_BIAS.n271 GND 0.005829f
C1128 CS_BIAS.n272 GND 0.005201f
C1129 CS_BIAS.n273 GND 0.011692f
C1130 CS_BIAS.t12 GND 0.185122f
C1131 CS_BIAS.n274 GND 0.070673f
C1132 CS_BIAS.n275 GND 0.00638f
C1133 CS_BIAS.n276 GND 0.005829f
C1134 CS_BIAS.n277 GND 0.005829f
C1135 CS_BIAS.n278 GND 0.005829f
C1136 CS_BIAS.n279 GND 0.008473f
C1137 CS_BIAS.n280 GND 0.008473f
C1138 CS_BIAS.n281 GND 0.009901f
C1139 CS_BIAS.n282 GND 0.005829f
C1140 CS_BIAS.n283 GND 0.005829f
C1141 CS_BIAS.n284 GND 0.00638f
C1142 CS_BIAS.n285 GND 0.011692f
C1143 CS_BIAS.n286 GND 0.005201f
C1144 CS_BIAS.n287 GND 0.005829f
C1145 CS_BIAS.n288 GND 0.005829f
C1146 CS_BIAS.n289 GND 0.005829f
C1147 CS_BIAS.n290 GND 0.008087f
C1148 CS_BIAS.n291 GND 0.070673f
C1149 CS_BIAS.n292 GND 0.008194f
C1150 CS_BIAS.n293 GND 0.010755f
C1151 CS_BIAS.n294 GND 0.005829f
C1152 CS_BIAS.n295 GND 0.005829f
C1153 CS_BIAS.n296 GND 0.005829f
C1154 CS_BIAS.n297 GND 0.01166f
C1155 CS_BIAS.n298 GND 0.006273f
C1156 CS_BIAS.n299 GND 0.070673f
C1157 CS_BIAS.n300 GND 0.010008f
C1158 CS_BIAS.n301 GND 0.005829f
C1159 CS_BIAS.n302 GND 0.005829f
C1160 CS_BIAS.n303 GND 0.005829f
C1161 CS_BIAS.n304 GND 0.008634f
C1162 CS_BIAS.n305 GND 0.009795f
C1163 CS_BIAS.n306 GND 0.088447f
C1164 CS_BIAS.n307 GND 0.058541f
C1165 CS_BIAS.t5 GND 0.010781f
C1166 CS_BIAS.t29 GND 0.010781f
C1167 CS_BIAS.n308 GND 0.094152f
C1168 CS_BIAS.n309 GND 0.1167f
C1169 CS_BIAS.t9 GND 0.010781f
C1170 CS_BIAS.t11 GND 0.010781f
C1171 CS_BIAS.n310 GND 0.094152f
C1172 CS_BIAS.n311 GND 0.061488f
C1173 CS_BIAS.n312 GND 0.064277f
C1174 CS_BIAS.n313 GND 0.037722f
C1175 CS_BIAS.n314 GND 0.005092f
C1176 CS_BIAS.n315 GND 0.008473f
C1177 CS_BIAS.n316 GND 0.008473f
C1178 CS_BIAS.n317 GND 0.009901f
C1179 CS_BIAS.n318 GND 0.005829f
C1180 CS_BIAS.n319 GND 0.005829f
C1181 CS_BIAS.n320 GND 0.00638f
C1182 CS_BIAS.n321 GND 0.011692f
C1183 CS_BIAS.n322 GND 0.005201f
C1184 CS_BIAS.n323 GND 0.005829f
C1185 CS_BIAS.n324 GND 0.005829f
C1186 CS_BIAS.n325 GND 0.005829f
C1187 CS_BIAS.n326 GND 0.008087f
C1188 CS_BIAS.n327 GND 0.070673f
C1189 CS_BIAS.n328 GND 0.008194f
C1190 CS_BIAS.n329 GND 0.010755f
C1191 CS_BIAS.n330 GND 0.005829f
C1192 CS_BIAS.n331 GND 0.005829f
C1193 CS_BIAS.n332 GND 0.005829f
C1194 CS_BIAS.n333 GND 0.01166f
C1195 CS_BIAS.n334 GND 0.006273f
C1196 CS_BIAS.n335 GND 0.070673f
C1197 CS_BIAS.n336 GND 0.010008f
C1198 CS_BIAS.n337 GND 0.005829f
C1199 CS_BIAS.n338 GND 0.005829f
C1200 CS_BIAS.n339 GND 0.005829f
C1201 CS_BIAS.n340 GND 0.008634f
C1202 CS_BIAS.n341 GND 0.009795f
C1203 CS_BIAS.n342 GND 0.088447f
C1204 CS_BIAS.n343 GND 0.035075f
C1205 CS_BIAS.n344 GND 0.007684f
C1206 CS_BIAS.t60 GND 0.185122f
C1207 CS_BIAS.n345 GND 0.008311f
C1208 CS_BIAS.n346 GND 0.005829f
C1209 CS_BIAS.t54 GND 0.185122f
C1210 CS_BIAS.n347 GND 0.005338f
C1211 CS_BIAS.n348 GND 0.005829f
C1212 CS_BIAS.t45 GND 0.185122f
C1213 CS_BIAS.n349 GND 0.010861f
C1214 CS_BIAS.n350 GND 0.005829f
C1215 CS_BIAS.t53 GND 0.185122f
C1216 CS_BIAS.n351 GND 0.070673f
C1217 CS_BIAS.n352 GND 0.005829f
C1218 CS_BIAS.n353 GND 0.009901f
C1219 CS_BIAS.n354 GND 0.005829f
C1220 CS_BIAS.n355 GND 0.010861f
C1221 CS_BIAS.n356 GND 0.005829f
C1222 CS_BIAS.t38 GND 0.185122f
C1223 CS_BIAS.n357 GND 0.005338f
C1224 CS_BIAS.n358 GND 0.043632f
C1225 CS_BIAS.t59 GND 0.185122f
C1226 CS_BIAS.t50 GND 0.214423f
C1227 CS_BIAS.n359 GND 0.084881f
C1228 CS_BIAS.n360 GND 0.082798f
C1229 CS_BIAS.n361 GND 0.006273f
C1230 CS_BIAS.n362 GND 0.01166f
C1231 CS_BIAS.n363 GND 0.005829f
C1232 CS_BIAS.n364 GND 0.005829f
C1233 CS_BIAS.n365 GND 0.005829f
C1234 CS_BIAS.n366 GND 0.010755f
C1235 CS_BIAS.n367 GND 0.008194f
C1236 CS_BIAS.n368 GND 0.070673f
C1237 CS_BIAS.n369 GND 0.008087f
C1238 CS_BIAS.n370 GND 0.005829f
C1239 CS_BIAS.n371 GND 0.005829f
C1240 CS_BIAS.n372 GND 0.005829f
C1241 CS_BIAS.n373 GND 0.005201f
C1242 CS_BIAS.n374 GND 0.011692f
C1243 CS_BIAS.t34 GND 0.185122f
C1244 CS_BIAS.n375 GND 0.070673f
C1245 CS_BIAS.n376 GND 0.00638f
C1246 CS_BIAS.n377 GND 0.005829f
C1247 CS_BIAS.n378 GND 0.005829f
C1248 CS_BIAS.n379 GND 0.005829f
C1249 CS_BIAS.n380 GND 0.008473f
C1250 CS_BIAS.n381 GND 0.008473f
C1251 CS_BIAS.n382 GND 0.009901f
C1252 CS_BIAS.n383 GND 0.005829f
C1253 CS_BIAS.n384 GND 0.005829f
C1254 CS_BIAS.n385 GND 0.00638f
C1255 CS_BIAS.n386 GND 0.011692f
C1256 CS_BIAS.n387 GND 0.005201f
C1257 CS_BIAS.n388 GND 0.005829f
C1258 CS_BIAS.n389 GND 0.005829f
C1259 CS_BIAS.n390 GND 0.005829f
C1260 CS_BIAS.n391 GND 0.008087f
C1261 CS_BIAS.n392 GND 0.070673f
C1262 CS_BIAS.n393 GND 0.008194f
C1263 CS_BIAS.n394 GND 0.010755f
C1264 CS_BIAS.n395 GND 0.005829f
C1265 CS_BIAS.n396 GND 0.005829f
C1266 CS_BIAS.n397 GND 0.005829f
C1267 CS_BIAS.n398 GND 0.01166f
C1268 CS_BIAS.n399 GND 0.006273f
C1269 CS_BIAS.n400 GND 0.070673f
C1270 CS_BIAS.n401 GND 0.010008f
C1271 CS_BIAS.n402 GND 0.005829f
C1272 CS_BIAS.n403 GND 0.005829f
C1273 CS_BIAS.n404 GND 0.005829f
C1274 CS_BIAS.n405 GND 0.008634f
C1275 CS_BIAS.n406 GND 0.009795f
C1276 CS_BIAS.n407 GND 0.088447f
C1277 CS_BIAS.n408 GND 0.021125f
C1278 CS_BIAS.n409 GND 0.154927f
C1279 CS_BIAS.n410 GND 2.87933f
C1280 VOUT.t48 GND 0.03946f
C1281 VOUT.t58 GND 0.03946f
C1282 VOUT.n0 GND 0.294307f
C1283 VOUT.t65 GND 0.03946f
C1284 VOUT.t76 GND 0.03946f
C1285 VOUT.n1 GND 0.29307f
C1286 VOUT.n2 GND 0.436055f
C1287 VOUT.t42 GND 0.03946f
C1288 VOUT.t53 GND 0.03946f
C1289 VOUT.n3 GND 0.29307f
C1290 VOUT.n4 GND 0.215773f
C1291 VOUT.t57 GND 0.03946f
C1292 VOUT.t72 GND 0.03946f
C1293 VOUT.n5 GND 0.29307f
C1294 VOUT.n6 GND 0.215773f
C1295 VOUT.t38 GND 0.03946f
C1296 VOUT.t47 GND 0.03946f
C1297 VOUT.n7 GND 0.29307f
C1298 VOUT.n8 GND 0.360556f
C1299 VOUT.t49 GND 0.03946f
C1300 VOUT.t84 GND 0.03946f
C1301 VOUT.n9 GND 0.294307f
C1302 VOUT.t39 GND 0.03946f
C1303 VOUT.t77 GND 0.03946f
C1304 VOUT.n10 GND 0.29307f
C1305 VOUT.n11 GND 0.436055f
C1306 VOUT.t25 GND 0.03946f
C1307 VOUT.t64 GND 0.03946f
C1308 VOUT.n12 GND 0.29307f
C1309 VOUT.n13 GND 0.215773f
C1310 VOUT.t79 GND 0.03946f
C1311 VOUT.t56 GND 0.03946f
C1312 VOUT.n14 GND 0.29307f
C1313 VOUT.n15 GND 0.215773f
C1314 VOUT.t66 GND 0.03946f
C1315 VOUT.t40 GND 0.03946f
C1316 VOUT.n16 GND 0.29307f
C1317 VOUT.n17 GND 0.298771f
C1318 VOUT.n18 GND 0.554227f
C1319 VOUT.t80 GND 0.03946f
C1320 VOUT.t52 GND 0.03946f
C1321 VOUT.n19 GND 0.294307f
C1322 VOUT.t68 GND 0.03946f
C1323 VOUT.t44 GND 0.03946f
C1324 VOUT.n20 GND 0.29307f
C1325 VOUT.n21 GND 0.436055f
C1326 VOUT.t54 GND 0.03946f
C1327 VOUT.t34 GND 0.03946f
C1328 VOUT.n22 GND 0.29307f
C1329 VOUT.n23 GND 0.215773f
C1330 VOUT.t46 GND 0.03946f
C1331 VOUT.t28 GND 0.03946f
C1332 VOUT.n24 GND 0.29307f
C1333 VOUT.n25 GND 0.215773f
C1334 VOUT.t35 GND 0.03946f
C1335 VOUT.t70 GND 0.03946f
C1336 VOUT.n26 GND 0.29307f
C1337 VOUT.n27 GND 0.298771f
C1338 VOUT.n28 GND 0.524897f
C1339 VOUT.n29 GND 5.96249f
C1340 VOUT.n31 GND 0.639555f
C1341 VOUT.n32 GND 0.479666f
C1342 VOUT.n33 GND 0.639555f
C1343 VOUT.n34 GND 0.639555f
C1344 VOUT.n35 GND 1.72188f
C1345 VOUT.n36 GND 0.639555f
C1346 VOUT.n37 GND 0.639555f
C1347 VOUT.t93 GND 0.799444f
C1348 VOUT.n38 GND 0.639555f
C1349 VOUT.n39 GND 0.639555f
C1350 VOUT.n43 GND 0.639555f
C1351 VOUT.n47 GND 0.639555f
C1352 VOUT.n48 GND 0.639555f
C1353 VOUT.n50 GND 0.639555f
C1354 VOUT.n55 GND 0.639555f
C1355 VOUT.n57 GND 0.639555f
C1356 VOUT.n58 GND 0.639555f
C1357 VOUT.n60 GND 0.639555f
C1358 VOUT.n61 GND 0.639555f
C1359 VOUT.n63 GND 0.639555f
C1360 VOUT.t96 GND 10.6869f
C1361 VOUT.n65 GND 0.639555f
C1362 VOUT.n66 GND 0.479666f
C1363 VOUT.n67 GND 0.639555f
C1364 VOUT.n68 GND 0.639555f
C1365 VOUT.n69 GND 1.72188f
C1366 VOUT.n70 GND 0.639555f
C1367 VOUT.n71 GND 0.639555f
C1368 VOUT.t94 GND 0.799444f
C1369 VOUT.n72 GND 0.639555f
C1370 VOUT.n73 GND 0.639555f
C1371 VOUT.n77 GND 0.639555f
C1372 VOUT.n81 GND 0.639555f
C1373 VOUT.n82 GND 0.639555f
C1374 VOUT.n84 GND 0.639555f
C1375 VOUT.n89 GND 0.639555f
C1376 VOUT.n91 GND 0.639555f
C1377 VOUT.n92 GND 0.639555f
C1378 VOUT.n94 GND 0.639555f
C1379 VOUT.n95 GND 0.639555f
C1380 VOUT.n97 GND 0.639555f
C1381 VOUT.n98 GND 0.479666f
C1382 VOUT.n100 GND 0.639555f
C1383 VOUT.n101 GND 0.479666f
C1384 VOUT.n102 GND 0.639555f
C1385 VOUT.n103 GND 0.639555f
C1386 VOUT.n104 GND 1.72188f
C1387 VOUT.n105 GND 0.639555f
C1388 VOUT.n106 GND 0.639555f
C1389 VOUT.t92 GND 0.799444f
C1390 VOUT.n107 GND 0.639555f
C1391 VOUT.n108 GND 1.72188f
C1392 VOUT.n110 GND 0.639555f
C1393 VOUT.n111 GND 0.639555f
C1394 VOUT.n113 GND 0.639555f
C1395 VOUT.n114 GND 0.639555f
C1396 VOUT.t95 GND 10.5127f
C1397 VOUT.t97 GND 10.6869f
C1398 VOUT.n120 GND 2.00638f
C1399 VOUT.n121 GND 8.173249f
C1400 VOUT.n122 GND 8.51525f
C1401 VOUT.n127 GND 2.17345f
C1402 VOUT.n133 GND 0.639555f
C1403 VOUT.n135 GND 0.639555f
C1404 VOUT.n137 GND 0.639555f
C1405 VOUT.n139 GND 0.639555f
C1406 VOUT.n141 GND 0.639555f
C1407 VOUT.n147 GND 0.639555f
C1408 VOUT.n154 GND 1.17334f
C1409 VOUT.n155 GND 1.17334f
C1410 VOUT.n156 GND 0.639555f
C1411 VOUT.n157 GND 0.639555f
C1412 VOUT.n159 GND 0.479666f
C1413 VOUT.n160 GND 0.410791f
C1414 VOUT.n162 GND 0.479666f
C1415 VOUT.n163 GND 0.410791f
C1416 VOUT.n164 GND 0.479666f
C1417 VOUT.n166 GND 0.639555f
C1418 VOUT.n168 GND 1.72188f
C1419 VOUT.n169 GND 2.00638f
C1420 VOUT.n170 GND 7.51729f
C1421 VOUT.n172 GND 0.479666f
C1422 VOUT.n173 GND 1.23421f
C1423 VOUT.n174 GND 0.479666f
C1424 VOUT.n176 GND 0.639555f
C1425 VOUT.n178 GND 1.72188f
C1426 VOUT.n179 GND 3.25722f
C1427 VOUT.n180 GND 2.19028f
C1428 VOUT.t73 GND 0.03946f
C1429 VOUT.t63 GND 0.03946f
C1430 VOUT.n181 GND 0.294307f
C1431 VOUT.t30 GND 0.03946f
C1432 VOUT.t81 GND 0.03946f
C1433 VOUT.n182 GND 0.29307f
C1434 VOUT.n183 GND 0.436055f
C1435 VOUT.t69 GND 0.03946f
C1436 VOUT.t37 GND 0.03946f
C1437 VOUT.n184 GND 0.29307f
C1438 VOUT.n185 GND 0.215773f
C1439 VOUT.t27 GND 0.03946f
C1440 VOUT.t74 GND 0.03946f
C1441 VOUT.n186 GND 0.29307f
C1442 VOUT.n187 GND 0.215773f
C1443 VOUT.t61 GND 0.03946f
C1444 VOUT.t31 GND 0.03946f
C1445 VOUT.n188 GND 0.29307f
C1446 VOUT.n189 GND 0.360556f
C1447 VOUT.t67 GND 0.03946f
C1448 VOUT.t33 GND 0.03946f
C1449 VOUT.n190 GND 0.294307f
C1450 VOUT.t59 GND 0.03946f
C1451 VOUT.t82 GND 0.03946f
C1452 VOUT.n191 GND 0.29307f
C1453 VOUT.n192 GND 0.436055f
C1454 VOUT.t45 GND 0.03946f
C1455 VOUT.t75 GND 0.03946f
C1456 VOUT.n193 GND 0.29307f
C1457 VOUT.n194 GND 0.215773f
C1458 VOUT.t41 GND 0.03946f
C1459 VOUT.t60 GND 0.03946f
C1460 VOUT.n195 GND 0.29307f
C1461 VOUT.n196 GND 0.215773f
C1462 VOUT.t83 GND 0.03946f
C1463 VOUT.t55 GND 0.03946f
C1464 VOUT.n197 GND 0.29307f
C1465 VOUT.n198 GND 0.298771f
C1466 VOUT.n199 GND 0.554227f
C1467 VOUT.t36 GND 0.03946f
C1468 VOUT.t62 GND 0.03946f
C1469 VOUT.n200 GND 0.294307f
C1470 VOUT.t29 GND 0.03946f
C1471 VOUT.t50 GND 0.03946f
C1472 VOUT.n201 GND 0.29307f
C1473 VOUT.n202 GND 0.436055f
C1474 VOUT.t78 GND 0.03946f
C1475 VOUT.t43 GND 0.03946f
C1476 VOUT.n203 GND 0.29307f
C1477 VOUT.n204 GND 0.215773f
C1478 VOUT.t71 GND 0.03946f
C1479 VOUT.t32 GND 0.03946f
C1480 VOUT.n205 GND 0.29307f
C1481 VOUT.n206 GND 0.215773f
C1482 VOUT.t51 GND 0.03946f
C1483 VOUT.t26 GND 0.03946f
C1484 VOUT.n207 GND 0.293069f
C1485 VOUT.n208 GND 0.298772f
C1486 VOUT.n209 GND 0.524897f
C1487 VOUT.n210 GND 8.53831f
C1488 VOUT.t7 GND 0.033823f
C1489 VOUT.t2 GND 0.033823f
C1490 VOUT.n211 GND 0.298278f
C1491 VOUT.t11 GND 0.033823f
C1492 VOUT.t19 GND 0.033823f
C1493 VOUT.n212 GND 0.295388f
C1494 VOUT.n213 GND 0.481012f
C1495 VOUT.t12 GND 0.033823f
C1496 VOUT.t87 GND 0.033823f
C1497 VOUT.n214 GND 0.295388f
C1498 VOUT.n215 GND 0.239078f
C1499 VOUT.t20 GND 0.033823f
C1500 VOUT.t5 GND 0.033823f
C1501 VOUT.n216 GND 0.295388f
C1502 VOUT.n217 GND 0.367871f
C1503 VOUT.t3 GND 0.033823f
C1504 VOUT.t86 GND 0.033823f
C1505 VOUT.n218 GND 0.298278f
C1506 VOUT.t24 GND 0.033823f
C1507 VOUT.t16 GND 0.033823f
C1508 VOUT.n219 GND 0.295388f
C1509 VOUT.n220 GND 0.481012f
C1510 VOUT.t90 GND 0.033823f
C1511 VOUT.t9 GND 0.033823f
C1512 VOUT.n221 GND 0.295388f
C1513 VOUT.n222 GND 0.239078f
C1514 VOUT.t0 GND 0.033823f
C1515 VOUT.t8 GND 0.033823f
C1516 VOUT.n223 GND 0.295388f
C1517 VOUT.n224 GND 0.315946f
C1518 VOUT.n225 GND 0.79475f
C1519 VOUT.n226 GND 8.79295f
C1520 VOUT.t4 GND 0.033823f
C1521 VOUT.t85 GND 0.033823f
C1522 VOUT.n227 GND 0.298278f
C1523 VOUT.t22 GND 0.033823f
C1524 VOUT.t89 GND 0.033823f
C1525 VOUT.n228 GND 0.295388f
C1526 VOUT.n229 GND 0.481012f
C1527 VOUT.t91 GND 0.033823f
C1528 VOUT.t21 GND 0.033823f
C1529 VOUT.n230 GND 0.295388f
C1530 VOUT.n231 GND 0.239078f
C1531 VOUT.t23 GND 0.033823f
C1532 VOUT.t14 GND 0.033823f
C1533 VOUT.n232 GND 0.295388f
C1534 VOUT.n233 GND 0.367871f
C1535 VOUT.t6 GND 0.033823f
C1536 VOUT.t15 GND 0.033823f
C1537 VOUT.n234 GND 0.298278f
C1538 VOUT.t88 GND 0.033823f
C1539 VOUT.t18 GND 0.033823f
C1540 VOUT.n235 GND 0.295388f
C1541 VOUT.n236 GND 0.481012f
C1542 VOUT.t17 GND 0.033823f
C1543 VOUT.t1 GND 0.033823f
C1544 VOUT.n237 GND 0.295388f
C1545 VOUT.n238 GND 0.239078f
C1546 VOUT.t10 GND 0.033823f
C1547 VOUT.t13 GND 0.033823f
C1548 VOUT.n239 GND 0.295388f
C1549 VOUT.n240 GND 0.315946f
C1550 VOUT.n241 GND 0.79475f
C1551 VOUT.n242 GND 5.30444f
C1552 VOUT.n243 GND 6.19757f
C1553 VDD.t189 GND 0.018235f
C1554 VDD.t11 GND 0.018235f
C1555 VDD.n0 GND 0.126171f
C1556 VDD.t98 GND 0.018235f
C1557 VDD.t8 GND 0.018235f
C1558 VDD.n1 GND 0.125509f
C1559 VDD.n2 GND 0.280867f
C1560 VDD.t195 GND 0.018235f
C1561 VDD.t100 GND 0.018235f
C1562 VDD.n3 GND 0.125509f
C1563 VDD.n4 GND 0.143521f
C1564 VDD.t6 GND 0.018235f
C1565 VDD.t13 GND 0.018235f
C1566 VDD.n5 GND 0.125509f
C1567 VDD.n6 GND 0.129676f
C1568 VDD.t20 GND 0.018235f
C1569 VDD.t106 GND 0.018235f
C1570 VDD.n7 GND 0.126171f
C1571 VDD.t16 GND 0.018235f
C1572 VDD.t2 GND 0.018235f
C1573 VDD.n8 GND 0.125509f
C1574 VDD.n9 GND 0.280867f
C1575 VDD.t104 GND 0.018235f
C1576 VDD.t191 GND 0.018235f
C1577 VDD.n10 GND 0.125509f
C1578 VDD.n11 GND 0.143521f
C1579 VDD.t193 GND 0.018235f
C1580 VDD.t4 GND 0.018235f
C1581 VDD.n12 GND 0.125509f
C1582 VDD.n13 GND 0.129676f
C1583 VDD.n14 GND 0.087702f
C1584 VDD.n15 GND 2.11138f
C1585 VDD.t176 GND 0.222206f
C1586 VDD.t165 GND 0.025529f
C1587 VDD.t118 GND 0.025529f
C1588 VDD.n16 GND 0.163847f
C1589 VDD.n17 GND 0.290589f
C1590 VDD.t184 GND 0.025529f
C1591 VDD.t173 GND 0.025529f
C1592 VDD.n18 GND 0.163847f
C1593 VDD.n19 GND 0.154853f
C1594 VDD.t132 GND 0.025529f
C1595 VDD.t113 GND 0.025529f
C1596 VDD.n20 GND 0.163847f
C1597 VDD.n21 GND 0.154853f
C1598 VDD.t177 GND 0.025529f
C1599 VDD.t166 GND 0.025529f
C1600 VDD.n22 GND 0.163847f
C1601 VDD.n23 GND 0.154853f
C1602 VDD.t121 GND 0.221218f
C1603 VDD.n24 GND 0.203521f
C1604 VDD.t171 GND 0.222206f
C1605 VDD.t123 GND 0.025529f
C1606 VDD.t163 GND 0.025529f
C1607 VDD.n25 GND 0.163847f
C1608 VDD.n26 GND 0.290589f
C1609 VDD.t185 GND 0.025529f
C1610 VDD.t143 GND 0.025529f
C1611 VDD.n27 GND 0.163847f
C1612 VDD.n28 GND 0.154853f
C1613 VDD.t178 GND 0.025529f
C1614 VDD.t137 GND 0.025529f
C1615 VDD.n29 GND 0.163847f
C1616 VDD.n30 GND 0.154853f
C1617 VDD.t164 GND 0.025529f
C1618 VDD.t186 GND 0.025529f
C1619 VDD.n31 GND 0.163847f
C1620 VDD.n32 GND 0.154853f
C1621 VDD.t158 GND 0.221218f
C1622 VDD.n33 GND 0.162349f
C1623 VDD.n34 GND 0.344539f
C1624 VDD.t129 GND 0.222206f
C1625 VDD.t167 GND 0.025529f
C1626 VDD.t117 GND 0.025529f
C1627 VDD.n35 GND 0.163847f
C1628 VDD.n36 GND 0.290589f
C1629 VDD.t151 GND 0.025529f
C1630 VDD.t181 GND 0.025529f
C1631 VDD.n37 GND 0.163847f
C1632 VDD.n38 GND 0.154853f
C1633 VDD.t139 GND 0.025529f
C1634 VDD.t159 GND 0.025529f
C1635 VDD.n39 GND 0.163847f
C1636 VDD.n40 GND 0.154853f
C1637 VDD.t120 GND 0.025529f
C1638 VDD.t153 GND 0.025529f
C1639 VDD.n41 GND 0.163847f
C1640 VDD.n42 GND 0.154853f
C1641 VDD.t111 GND 0.221218f
C1642 VDD.n43 GND 0.162349f
C1643 VDD.n44 GND 0.303846f
C1644 VDD.n45 GND 0.006965f
C1645 VDD.n46 GND 0.009062f
C1646 VDD.n47 GND 0.007294f
C1647 VDD.n48 GND 0.007294f
C1648 VDD.n49 GND 0.009062f
C1649 VDD.n50 GND 0.009062f
C1650 VDD.n51 GND 0.643537f
C1651 VDD.n52 GND 0.009062f
C1652 VDD.n53 GND 0.009062f
C1653 VDD.n54 GND 0.009062f
C1654 VDD.n55 GND 0.523973f
C1655 VDD.n56 GND 0.009062f
C1656 VDD.n57 GND 0.009062f
C1657 VDD.n58 GND 0.009062f
C1658 VDD.n59 GND 0.009062f
C1659 VDD.n60 GND 0.007294f
C1660 VDD.n61 GND 0.009062f
C1661 VDD.t112 GND 0.35166f
C1662 VDD.n62 GND 0.009062f
C1663 VDD.n63 GND 0.009062f
C1664 VDD.n64 GND 0.009062f
C1665 VDD.t119 GND 0.35166f
C1666 VDD.n65 GND 0.009062f
C1667 VDD.n66 GND 0.009062f
C1668 VDD.n67 GND 0.009062f
C1669 VDD.n68 GND 0.009062f
C1670 VDD.n69 GND 0.009062f
C1671 VDD.n70 GND 0.007294f
C1672 VDD.n71 GND 0.009062f
C1673 VDD.n72 GND 0.65057f
C1674 VDD.n73 GND 0.009062f
C1675 VDD.n74 GND 0.009062f
C1676 VDD.n75 GND 0.009062f
C1677 VDD.n76 GND 0.51694f
C1678 VDD.n77 GND 0.009062f
C1679 VDD.n78 GND 0.009062f
C1680 VDD.n79 GND 0.009062f
C1681 VDD.n80 GND 0.009062f
C1682 VDD.n81 GND 0.009062f
C1683 VDD.n82 GND 0.007294f
C1684 VDD.n83 GND 0.009062f
C1685 VDD.t110 GND 0.35166f
C1686 VDD.n84 GND 0.009062f
C1687 VDD.n85 GND 0.009062f
C1688 VDD.n86 GND 0.009062f
C1689 VDD.n87 GND 0.703319f
C1690 VDD.n88 GND 0.009062f
C1691 VDD.n89 GND 0.009062f
C1692 VDD.n90 GND 0.009062f
C1693 VDD.n91 GND 0.009062f
C1694 VDD.n92 GND 0.009062f
C1695 VDD.n93 GND 0.007294f
C1696 VDD.n94 GND 0.009062f
C1697 VDD.n95 GND 0.009062f
C1698 VDD.n96 GND 0.009062f
C1699 VDD.n97 GND 0.02036f
C1700 VDD.n98 GND 1.52972f
C1701 VDD.n99 GND 0.02042f
C1702 VDD.n100 GND 0.009062f
C1703 VDD.n101 GND 0.009062f
C1704 VDD.n103 GND 0.009062f
C1705 VDD.n104 GND 0.009062f
C1706 VDD.n105 GND 0.007294f
C1707 VDD.n106 GND 0.007294f
C1708 VDD.n107 GND 0.009062f
C1709 VDD.n108 GND 0.009062f
C1710 VDD.n109 GND 0.009062f
C1711 VDD.n110 GND 0.009062f
C1712 VDD.n111 GND 0.009062f
C1713 VDD.n112 GND 0.009062f
C1714 VDD.n113 GND 0.007294f
C1715 VDD.n115 GND 0.009062f
C1716 VDD.n116 GND 0.009062f
C1717 VDD.n117 GND 0.009062f
C1718 VDD.n118 GND 0.009062f
C1719 VDD.n119 GND 0.009062f
C1720 VDD.n120 GND 0.007294f
C1721 VDD.n122 GND 0.009062f
C1722 VDD.n123 GND 0.009062f
C1723 VDD.n124 GND 0.009062f
C1724 VDD.n125 GND 0.009062f
C1725 VDD.n126 GND 0.009062f
C1726 VDD.n127 GND 0.00609f
C1727 VDD.n129 GND 0.009062f
C1728 VDD.n130 GND 0.00609f
C1729 VDD.t53 GND 0.18563f
C1730 VDD.t52 GND 0.194533f
C1731 VDD.t50 GND 0.271204f
C1732 VDD.n131 GND 0.091924f
C1733 VDD.n132 GND 0.052705f
C1734 VDD.n133 GND 0.009062f
C1735 VDD.n134 GND 0.009062f
C1736 VDD.n135 GND 0.007294f
C1737 VDD.n137 GND 0.009062f
C1738 VDD.n138 GND 0.009062f
C1739 VDD.n139 GND 0.009062f
C1740 VDD.n140 GND 0.009062f
C1741 VDD.n141 GND 0.007294f
C1742 VDD.n143 GND 0.009062f
C1743 VDD.n144 GND 0.009062f
C1744 VDD.n145 GND 0.009062f
C1745 VDD.n146 GND 0.009062f
C1746 VDD.n147 GND 0.009062f
C1747 VDD.n148 GND 0.007294f
C1748 VDD.n150 GND 0.009062f
C1749 VDD.n151 GND 0.009062f
C1750 VDD.n152 GND 0.009062f
C1751 VDD.n153 GND 0.009062f
C1752 VDD.n154 GND 0.009062f
C1753 VDD.n155 GND 0.007294f
C1754 VDD.n157 GND 0.009062f
C1755 VDD.n158 GND 0.009062f
C1756 VDD.n159 GND 0.009062f
C1757 VDD.n160 GND 0.009062f
C1758 VDD.n161 GND 0.009062f
C1759 VDD.n162 GND 0.00496f
C1760 VDD.n164 GND 0.009062f
C1761 VDD.n165 GND 0.007221f
C1762 VDD.t90 GND 0.18563f
C1763 VDD.t89 GND 0.194533f
C1764 VDD.t88 GND 0.271204f
C1765 VDD.n166 GND 0.091924f
C1766 VDD.n167 GND 0.052705f
C1767 VDD.n168 GND 0.009062f
C1768 VDD.n169 GND 0.009062f
C1769 VDD.n170 GND 0.007294f
C1770 VDD.n172 GND 0.009062f
C1771 VDD.n173 GND 0.009062f
C1772 VDD.n174 GND 0.009062f
C1773 VDD.n175 GND 0.009062f
C1774 VDD.n176 GND 0.007294f
C1775 VDD.n178 GND 0.009062f
C1776 VDD.n179 GND 0.009062f
C1777 VDD.n180 GND 0.009062f
C1778 VDD.n181 GND 0.009062f
C1779 VDD.n182 GND 0.009062f
C1780 VDD.n183 GND 0.007294f
C1781 VDD.n185 GND 0.009062f
C1782 VDD.n186 GND 0.009062f
C1783 VDD.n187 GND 0.009062f
C1784 VDD.n188 GND 0.009062f
C1785 VDD.n189 GND 0.009062f
C1786 VDD.n190 GND 0.007294f
C1787 VDD.n192 GND 0.009062f
C1788 VDD.n193 GND 0.009062f
C1789 VDD.n194 GND 0.009062f
C1790 VDD.n195 GND 0.009062f
C1791 VDD.n196 GND 0.009062f
C1792 VDD.n197 GND 0.003829f
C1793 VDD.t59 GND 0.18563f
C1794 VDD.t58 GND 0.194533f
C1795 VDD.t57 GND 0.271204f
C1796 VDD.n199 GND 0.091924f
C1797 VDD.n200 GND 0.052705f
C1798 VDD.n201 GND 0.011269f
C1799 VDD.n202 GND 0.009062f
C1800 VDD.n203 GND 0.009062f
C1801 VDD.n204 GND 0.009062f
C1802 VDD.n205 GND 0.007294f
C1803 VDD.n206 GND 0.009062f
C1804 VDD.n207 GND 0.009062f
C1805 VDD.n208 GND 0.007294f
C1806 VDD.n209 GND 0.009062f
C1807 VDD.n210 GND 0.009062f
C1808 VDD.n211 GND 0.007294f
C1809 VDD.n212 GND 0.009062f
C1810 VDD.n213 GND 0.009062f
C1811 VDD.n214 GND 0.007294f
C1812 VDD.n215 GND 0.009062f
C1813 VDD.n216 GND 0.007294f
C1814 VDD.n217 GND 0.009062f
C1815 VDD.n218 GND 0.007294f
C1816 VDD.n219 GND 0.009062f
C1817 VDD.n220 GND 0.009062f
C1818 VDD.n221 GND 0.703319f
C1819 VDD.t142 GND 0.35166f
C1820 VDD.n222 GND 0.009062f
C1821 VDD.n223 GND 0.007294f
C1822 VDD.n224 GND 0.009062f
C1823 VDD.n225 GND 0.007294f
C1824 VDD.n226 GND 0.009062f
C1825 VDD.t150 GND 0.35166f
C1826 VDD.n227 GND 0.009062f
C1827 VDD.n228 GND 0.007294f
C1828 VDD.n229 GND 0.009062f
C1829 VDD.n230 GND 0.007294f
C1830 VDD.n231 GND 0.009062f
C1831 VDD.n232 GND 0.404409f
C1832 VDD.n233 GND 0.531006f
C1833 VDD.n234 GND 0.009062f
C1834 VDD.n235 GND 0.007294f
C1835 VDD.n236 GND 0.009062f
C1836 VDD.n237 GND 0.007294f
C1837 VDD.n238 GND 0.009062f
C1838 VDD.n239 GND 0.636504f
C1839 VDD.n240 GND 0.009062f
C1840 VDD.n241 GND 0.007294f
C1841 VDD.n242 GND 0.009062f
C1842 VDD.n243 GND 0.007294f
C1843 VDD.n244 GND 0.009062f
C1844 VDD.n245 GND 0.703319f
C1845 VDD.t122 GND 0.35166f
C1846 VDD.n246 GND 0.009062f
C1847 VDD.n247 GND 0.007294f
C1848 VDD.n248 GND 0.009062f
C1849 VDD.n249 GND 0.007294f
C1850 VDD.n250 GND 0.009062f
C1851 VDD.t128 GND 0.35166f
C1852 VDD.n251 GND 0.009062f
C1853 VDD.n252 GND 0.007294f
C1854 VDD.n253 GND 0.009062f
C1855 VDD.n254 GND 0.007294f
C1856 VDD.n255 GND 0.009062f
C1857 VDD.n256 GND 0.703319f
C1858 VDD.n257 GND 0.538039f
C1859 VDD.n258 GND 0.009062f
C1860 VDD.n259 GND 0.007294f
C1861 VDD.n260 GND 0.009062f
C1862 VDD.n261 GND 0.007294f
C1863 VDD.n262 GND 0.009062f
C1864 VDD.n263 GND 0.460674f
C1865 VDD.n264 GND 0.009062f
C1866 VDD.n265 GND 0.007294f
C1867 VDD.n266 GND 0.02036f
C1868 VDD.n267 GND 0.006054f
C1869 VDD.n268 GND 0.02036f
C1870 VDD.n269 GND 0.903766f
C1871 VDD.t44 GND 0.35166f
C1872 VDD.n270 GND 0.02036f
C1873 VDD.n271 GND 0.006054f
C1874 VDD.n272 GND 0.009062f
C1875 VDD.n273 GND 0.007294f
C1876 VDD.n274 GND 0.009062f
C1877 VDD.t82 GND 3.52363f
C1878 VDD.n302 GND 0.02042f
C1879 VDD.n303 GND 0.009062f
C1880 VDD.n304 GND 0.009062f
C1881 VDD.n305 GND 0.009062f
C1882 VDD.n306 GND 0.009062f
C1883 VDD.n307 GND 0.009062f
C1884 VDD.n308 GND 0.007794f
C1885 VDD.n309 GND 0.007294f
C1886 VDD.n310 GND 0.0058f
C1887 VDD.n311 GND 0.011006f
C1888 VDD.n312 GND 0.009062f
C1889 VDD.n313 GND 0.009062f
C1890 VDD.n314 GND 0.007294f
C1891 VDD.n315 GND 0.009062f
C1892 VDD.n316 GND 0.009062f
C1893 VDD.n317 GND 0.009062f
C1894 VDD.n318 GND 0.009062f
C1895 VDD.n319 GND 0.009062f
C1896 VDD.n320 GND 0.009062f
C1897 VDD.n321 GND 0.00609f
C1898 VDD.n322 GND 0.009062f
C1899 VDD.n323 GND 0.009062f
C1900 VDD.n324 GND 0.009062f
C1901 VDD.n325 GND 0.009062f
C1902 VDD.n326 GND 0.009062f
C1903 VDD.n327 GND 0.009062f
C1904 VDD.n328 GND 0.009062f
C1905 VDD.n329 GND 0.009062f
C1906 VDD.n330 GND 0.009062f
C1907 VDD.n331 GND 0.009062f
C1908 VDD.n332 GND 0.009062f
C1909 VDD.n333 GND 0.009062f
C1910 VDD.n334 GND 0.009062f
C1911 VDD.n335 GND 0.009062f
C1912 VDD.n336 GND 0.009062f
C1913 VDD.n337 GND 0.009062f
C1914 VDD.n338 GND 0.009062f
C1915 VDD.n339 GND 0.007221f
C1916 VDD.t45 GND 0.18563f
C1917 VDD.t46 GND 0.194533f
C1918 VDD.t43 GND 0.271204f
C1919 VDD.n340 GND 0.091924f
C1920 VDD.n341 GND 0.052705f
C1921 VDD.n342 GND 0.009062f
C1922 VDD.n343 GND 0.009062f
C1923 VDD.n344 GND 0.009062f
C1924 VDD.n345 GND 0.009062f
C1925 VDD.n346 GND 0.009062f
C1926 VDD.n347 GND 0.009062f
C1927 VDD.n348 GND 0.0058f
C1928 VDD.n349 GND 0.007294f
C1929 VDD.n350 GND 0.007794f
C1930 VDD.n351 GND 0.006162f
C1931 VDD.n352 GND 0.006162f
C1932 VDD.n353 GND 0.006162f
C1933 VDD.n354 GND 0.534523f
C1934 VDD.n355 GND 0.006162f
C1935 VDD.n356 GND 0.006162f
C1936 VDD.n357 GND 0.006162f
C1937 VDD.n359 GND 0.006162f
C1938 VDD.t39 GND 0.122823f
C1939 VDD.t38 GND 0.131225f
C1940 VDD.t36 GND 0.198505f
C1941 VDD.n360 GND 0.075862f
C1942 VDD.n361 GND 0.050543f
C1943 VDD.n362 GND 0.006162f
C1944 VDD.n364 GND 0.014027f
C1945 VDD.n365 GND 0.006162f
C1946 VDD.n366 GND 0.006162f
C1947 VDD.n367 GND 0.478257f
C1948 VDD.n368 GND 0.006162f
C1949 VDD.n369 GND 0.68222f
C1950 VDD.n370 GND 0.006162f
C1951 VDD.n371 GND 0.006162f
C1952 VDD.n372 GND 0.014027f
C1953 VDD.n373 GND 0.006162f
C1954 VDD.n374 GND 0.006162f
C1955 VDD.n375 GND 0.006162f
C1956 VDD.n376 GND 0.006162f
C1957 VDD.n378 GND 0.006162f
C1958 VDD.n379 GND 0.006162f
C1959 VDD.n381 GND 0.006162f
C1960 VDD.n382 GND 0.006162f
C1961 VDD.n384 GND 0.006162f
C1962 VDD.n385 GND 0.004848f
C1963 VDD.n387 GND 0.006162f
C1964 VDD.t49 GND 0.122823f
C1965 VDD.t48 GND 0.131225f
C1966 VDD.t47 GND 0.198505f
C1967 VDD.n388 GND 0.075862f
C1968 VDD.n389 GND 0.050543f
C1969 VDD.n390 GND 0.008807f
C1970 VDD.n391 GND 0.006162f
C1971 VDD.n392 GND 0.006162f
C1972 VDD.t37 GND 0.239129f
C1973 VDD.n393 GND 0.006162f
C1974 VDD.n394 GND 0.006162f
C1975 VDD.n395 GND 0.006162f
C1976 VDD.n396 GND 0.006162f
C1977 VDD.n397 GND 0.006162f
C1978 VDD.n398 GND 0.478257f
C1979 VDD.n399 GND 0.006162f
C1980 VDD.n400 GND 0.006162f
C1981 VDD.t105 GND 0.239129f
C1982 VDD.n401 GND 0.006162f
C1983 VDD.n402 GND 0.006162f
C1984 VDD.n403 GND 0.006162f
C1985 VDD.n404 GND 0.006162f
C1986 VDD.n405 GND 0.429025f
C1987 VDD.n406 GND 0.006162f
C1988 VDD.n407 GND 0.006162f
C1989 VDD.n408 GND 0.006162f
C1990 VDD.n409 GND 0.006162f
C1991 VDD.n410 GND 0.006162f
C1992 VDD.n411 GND 0.270778f
C1993 VDD.n412 GND 0.006162f
C1994 VDD.n413 GND 0.006162f
C1995 VDD.t19 GND 0.239129f
C1996 VDD.n414 GND 0.006162f
C1997 VDD.n415 GND 0.006162f
C1998 VDD.n416 GND 0.006162f
C1999 VDD.n417 GND 0.407925f
C2000 VDD.n418 GND 0.006162f
C2001 VDD.n419 GND 0.006162f
C2002 VDD.t107 GND 0.239129f
C2003 VDD.n420 GND 0.006162f
C2004 VDD.n421 GND 0.006162f
C2005 VDD.n422 GND 0.006162f
C2006 VDD.n423 GND 0.249678f
C2007 VDD.n424 GND 0.006162f
C2008 VDD.n425 GND 0.006162f
C2009 VDD.t1 GND 0.239129f
C2010 VDD.n426 GND 0.006162f
C2011 VDD.n427 GND 0.006162f
C2012 VDD.n428 GND 0.006162f
C2013 VDD.n429 GND 0.386826f
C2014 VDD.n430 GND 0.006162f
C2015 VDD.n431 GND 0.006162f
C2016 VDD.t18 GND 0.239129f
C2017 VDD.n432 GND 0.006162f
C2018 VDD.n433 GND 0.006162f
C2019 VDD.n434 GND 0.006162f
C2020 VDD.t101 GND 0.239129f
C2021 VDD.n435 GND 0.006162f
C2022 VDD.n436 GND 0.006162f
C2023 VDD.t15 GND 0.239129f
C2024 VDD.n437 GND 0.006162f
C2025 VDD.n438 GND 0.006162f
C2026 VDD.n439 GND 0.006162f
C2027 VDD.n440 GND 0.478257f
C2028 VDD.n441 GND 0.006162f
C2029 VDD.n442 GND 0.006162f
C2030 VDD.n443 GND 0.249678f
C2031 VDD.n444 GND 0.006162f
C2032 VDD.n445 GND 0.006162f
C2033 VDD.n446 GND 0.006162f
C2034 VDD.t9 GND 0.239129f
C2035 VDD.n447 GND 0.006162f
C2036 VDD.n448 GND 0.006162f
C2037 VDD.n449 GND 0.006162f
C2038 VDD.n450 GND 0.006162f
C2039 VDD.n451 GND 0.006162f
C2040 VDD.n452 GND 0.478257f
C2041 VDD.n453 GND 0.006162f
C2042 VDD.n454 GND 0.006162f
C2043 VDD.t190 GND 0.239129f
C2044 VDD.n455 GND 0.006162f
C2045 VDD.n456 GND 0.006162f
C2046 VDD.n457 GND 0.006162f
C2047 VDD.n458 GND 0.372759f
C2048 VDD.n459 GND 0.006162f
C2049 VDD.n460 GND 0.006162f
C2050 VDD.n461 GND 0.006162f
C2051 VDD.n462 GND 0.006162f
C2052 VDD.n463 GND 0.006162f
C2053 VDD.n464 GND 0.474741f
C2054 VDD.n465 GND 0.006162f
C2055 VDD.n466 GND 0.006162f
C2056 VDD.t103 GND 0.239129f
C2057 VDD.n467 GND 0.006162f
C2058 VDD.n468 GND 0.006162f
C2059 VDD.n469 GND 0.006162f
C2060 VDD.n470 GND 0.35166f
C2061 VDD.n471 GND 0.006162f
C2062 VDD.n472 GND 0.006162f
C2063 VDD.t78 GND 0.239129f
C2064 VDD.n473 GND 0.006162f
C2065 VDD.n474 GND 0.014027f
C2066 VDD.n475 GND 0.014027f
C2067 VDD.n476 GND 0.68222f
C2068 VDD.n477 GND 0.006162f
C2069 VDD.n478 GND 0.006162f
C2070 VDD.t3 GND 0.239129f
C2071 VDD.n479 GND 0.014027f
C2072 VDD.n480 GND 0.006162f
C2073 VDD.n481 GND 0.006162f
C2074 VDD.n482 GND 0.68222f
C2075 VDD.n494 GND 0.014791f
C2076 VDD.n506 GND 0.014027f
C2077 VDD.n507 GND 0.006162f
C2078 VDD.n508 GND 0.014027f
C2079 VDD.t93 GND 0.122823f
C2080 VDD.t92 GND 0.131225f
C2081 VDD.t91 GND 0.198505f
C2082 VDD.n509 GND 0.075862f
C2083 VDD.n510 GND 0.050543f
C2084 VDD.n511 GND 0.014756f
C2085 VDD.n512 GND 0.006162f
C2086 VDD.n513 GND 0.006162f
C2087 VDD.t5 GND 0.239129f
C2088 VDD.n514 GND 0.006162f
C2089 VDD.n515 GND 0.006162f
C2090 VDD.n516 GND 0.006162f
C2091 VDD.n517 GND 0.006162f
C2092 VDD.n518 GND 0.006162f
C2093 VDD.t64 GND 0.239129f
C2094 VDD.n519 GND 0.006162f
C2095 VDD.n520 GND 0.006162f
C2096 VDD.n521 GND 0.35166f
C2097 VDD.n522 GND 0.006162f
C2098 VDD.n523 GND 0.006162f
C2099 VDD.n524 GND 0.006162f
C2100 VDD.t66 GND 0.122823f
C2101 VDD.t65 GND 0.131225f
C2102 VDD.t63 GND 0.198505f
C2103 VDD.n525 GND 0.075862f
C2104 VDD.n526 GND 0.050543f
C2105 VDD.n527 GND 0.008807f
C2106 VDD.n528 GND 0.006162f
C2107 VDD.n529 GND 0.006162f
C2108 VDD.n530 GND 0.344627f
C2109 VDD.n531 GND 0.006162f
C2110 VDD.n532 GND 0.006162f
C2111 VDD.n533 GND 0.006162f
C2112 VDD.n534 GND 0.478257f
C2113 VDD.n535 GND 0.006162f
C2114 VDD.t99 GND 0.239129f
C2115 VDD.n536 GND 0.006162f
C2116 VDD.n537 GND 0.006162f
C2117 VDD.n538 GND 0.006162f
C2118 VDD.n539 GND 0.006162f
C2119 VDD.n540 GND 0.006162f
C2120 VDD.n541 GND 0.323527f
C2121 VDD.n542 GND 0.006162f
C2122 VDD.n543 GND 0.006162f
C2123 VDD.n544 GND 0.006162f
C2124 VDD.n545 GND 0.006162f
C2125 VDD.n546 GND 0.006162f
C2126 VDD.n547 GND 0.006162f
C2127 VDD.t14 GND 0.239129f
C2128 VDD.n548 GND 0.006162f
C2129 VDD.n549 GND 0.006162f
C2130 VDD.t194 GND 0.239129f
C2131 VDD.n550 GND 0.006162f
C2132 VDD.n551 GND 0.006162f
C2133 VDD.n552 GND 0.006162f
C2134 VDD.n553 GND 0.478257f
C2135 VDD.n554 GND 0.006162f
C2136 VDD.n555 GND 0.006162f
C2137 VDD.n556 GND 0.446608f
C2138 VDD.n557 GND 0.006162f
C2139 VDD.n558 GND 0.006162f
C2140 VDD.n559 GND 0.006162f
C2141 VDD.t17 GND 0.239129f
C2142 VDD.n560 GND 0.006162f
C2143 VDD.n561 GND 0.006162f
C2144 VDD.n562 GND 0.006162f
C2145 VDD.n563 GND 0.006162f
C2146 VDD.n564 GND 0.006162f
C2147 VDD.n565 GND 0.467707f
C2148 VDD.n566 GND 0.006162f
C2149 VDD.n567 GND 0.006162f
C2150 VDD.t7 GND 0.239129f
C2151 VDD.n568 GND 0.006162f
C2152 VDD.n569 GND 0.006162f
C2153 VDD.n570 GND 0.006162f
C2154 VDD.n571 GND 0.309461f
C2155 VDD.n572 GND 0.006162f
C2156 VDD.n573 GND 0.006162f
C2157 VDD.t0 GND 0.239129f
C2158 VDD.n574 GND 0.006162f
C2159 VDD.n575 GND 0.006162f
C2160 VDD.n576 GND 0.006162f
C2161 VDD.n577 GND 0.446608f
C2162 VDD.n578 GND 0.006162f
C2163 VDD.n579 GND 0.006162f
C2164 VDD.t97 GND 0.239129f
C2165 VDD.n580 GND 0.006162f
C2166 VDD.n581 GND 0.006162f
C2167 VDD.n582 GND 0.006162f
C2168 VDD.n583 GND 0.288361f
C2169 VDD.n584 GND 0.006162f
C2170 VDD.n585 GND 0.006162f
C2171 VDD.t102 GND 0.239129f
C2172 VDD.n586 GND 0.006162f
C2173 VDD.n587 GND 0.006162f
C2174 VDD.n588 GND 0.006162f
C2175 VDD.n589 GND 0.478257f
C2176 VDD.n590 GND 0.006162f
C2177 VDD.n591 GND 0.006162f
C2178 VDD.t10 GND 0.239129f
C2179 VDD.n592 GND 0.006162f
C2180 VDD.n593 GND 0.006162f
C2181 VDD.n594 GND 0.006162f
C2182 VDD.n595 GND 0.267261f
C2183 VDD.n596 GND 0.006162f
C2184 VDD.n597 GND 0.006162f
C2185 VDD.n598 GND 0.006162f
C2186 VDD.n599 GND 0.006162f
C2187 VDD.n600 GND 0.006162f
C2188 VDD.t71 GND 0.239129f
C2189 VDD.n601 GND 0.006162f
C2190 VDD.n602 GND 0.006162f
C2191 VDD.t188 GND 0.239129f
C2192 VDD.n603 GND 0.006162f
C2193 VDD.n604 GND 0.006162f
C2194 VDD.n605 GND 0.006162f
C2195 VDD.n606 GND 0.478257f
C2196 VDD.n607 GND 0.006162f
C2197 VDD.n608 GND 0.006162f
C2198 VDD.n609 GND 0.242645f
C2199 VDD.n610 GND 0.006162f
C2200 VDD.n611 GND 0.014791f
C2201 VDD.n612 GND 0.014791f
C2202 VDD.n613 GND 0.534523f
C2203 VDD.n614 GND 0.014027f
C2204 VDD.n615 GND 0.014027f
C2205 VDD.n616 GND 0.014791f
C2206 VDD.t27 GND 0.131225f
C2207 VDD.t25 GND 0.198505f
C2208 VDD.t28 GND 0.131225f
C2209 VDD.n617 GND 0.130384f
C2210 VDD.n618 GND 0.006162f
C2211 VDD.n619 GND 0.006162f
C2212 VDD.n620 GND 0.006162f
C2213 VDD.n621 GND 0.006162f
C2214 VDD.n622 GND 0.006162f
C2215 VDD.n623 GND 0.006162f
C2216 VDD.n624 GND 0.006162f
C2217 VDD.n625 GND 0.0058f
C2218 VDD.n628 GND 0.009062f
C2219 VDD.n629 GND 0.007294f
C2220 VDD.n630 GND 0.009062f
C2221 VDD.n631 GND 0.009062f
C2222 VDD.n632 GND 0.009062f
C2223 VDD.n633 GND 0.007294f
C2224 VDD.n634 GND 0.009062f
C2225 VDD.n635 GND 0.009062f
C2226 VDD.n636 GND 0.009062f
C2227 VDD.n637 GND 0.02042f
C2228 VDD.n638 GND 0.009062f
C2229 VDD.n639 GND 0.007294f
C2230 VDD.n640 GND 0.009062f
C2231 VDD.n641 GND 0.594305f
C2232 VDD.n643 GND 0.009062f
C2233 VDD.t26 GND 3.52363f
C2234 VDD.n646 GND 3.9843f
C2235 VDD.n647 GND 0.009062f
C2236 VDD.n648 GND 0.02042f
C2237 VDD.n649 GND 0.007294f
C2238 VDD.n650 GND 0.009062f
C2239 VDD.n651 GND 0.007294f
C2240 VDD.n652 GND 0.009062f
C2241 VDD.n653 GND 0.703319f
C2242 VDD.n654 GND 0.009062f
C2243 VDD.n655 GND 0.007294f
C2244 VDD.n656 GND 0.009062f
C2245 VDD.n657 GND 0.007294f
C2246 VDD.n658 GND 0.009062f
C2247 VDD.n659 GND 0.703319f
C2248 VDD.n660 GND 0.009062f
C2249 VDD.n661 GND 0.007294f
C2250 VDD.n662 GND 0.009062f
C2251 VDD.n663 GND 0.007294f
C2252 VDD.n664 GND 0.009062f
C2253 VDD.t154 GND 0.35166f
C2254 VDD.n665 GND 0.009062f
C2255 VDD.n666 GND 0.007294f
C2256 VDD.n667 GND 0.009062f
C2257 VDD.n668 GND 0.007294f
C2258 VDD.n669 GND 0.009062f
C2259 VDD.n670 GND 0.418475f
C2260 VDD.n671 GND 0.51694f
C2261 VDD.n672 GND 0.009062f
C2262 VDD.n673 GND 0.007294f
C2263 VDD.n674 GND 0.009062f
C2264 VDD.n675 GND 0.007294f
C2265 VDD.n676 GND 0.009062f
C2266 VDD.n677 GND 0.65057f
C2267 VDD.n678 GND 0.009062f
C2268 VDD.n679 GND 0.007294f
C2269 VDD.n680 GND 0.009062f
C2270 VDD.n681 GND 0.007294f
C2271 VDD.n682 GND 0.009062f
C2272 VDD.n683 GND 0.703319f
C2273 VDD.t140 GND 0.35166f
C2274 VDD.n684 GND 0.009062f
C2275 VDD.n685 GND 0.007294f
C2276 VDD.n686 GND 0.009062f
C2277 VDD.n687 GND 0.007294f
C2278 VDD.n688 GND 0.009062f
C2279 VDD.t133 GND 0.35166f
C2280 VDD.n689 GND 0.009062f
C2281 VDD.n690 GND 0.007294f
C2282 VDD.n691 GND 0.009062f
C2283 VDD.n692 GND 0.007294f
C2284 VDD.n693 GND 0.009062f
C2285 VDD.n694 GND 0.411442f
C2286 VDD.n695 GND 0.523973f
C2287 VDD.n696 GND 0.009062f
C2288 VDD.n697 GND 0.007294f
C2289 VDD.t162 GND 0.222206f
C2290 VDD.t179 GND 0.025529f
C2291 VDD.t148 GND 0.025529f
C2292 VDD.n698 GND 0.163847f
C2293 VDD.n699 GND 0.290589f
C2294 VDD.t156 GND 0.025529f
C2295 VDD.t169 GND 0.025529f
C2296 VDD.n700 GND 0.163847f
C2297 VDD.n701 GND 0.154853f
C2298 VDD.t175 GND 0.025529f
C2299 VDD.t138 GND 0.025529f
C2300 VDD.n702 GND 0.163847f
C2301 VDD.n703 GND 0.154853f
C2302 VDD.t144 GND 0.025529f
C2303 VDD.t161 GND 0.025529f
C2304 VDD.n704 GND 0.163847f
C2305 VDD.n705 GND 0.154853f
C2306 VDD.t130 GND 0.221218f
C2307 VDD.n706 GND 0.203521f
C2308 VDD.t187 GND 0.222206f
C2309 VDD.t180 GND 0.025529f
C2310 VDD.t149 GND 0.025529f
C2311 VDD.n707 GND 0.163847f
C2312 VDD.n708 GND 0.290589f
C2313 VDD.t168 GND 0.025529f
C2314 VDD.t134 GND 0.025529f
C2315 VDD.n709 GND 0.163847f
C2316 VDD.n710 GND 0.154853f
C2317 VDD.t160 GND 0.025529f
C2318 VDD.t109 GND 0.025529f
C2319 VDD.n711 GND 0.163847f
C2320 VDD.n712 GND 0.154853f
C2321 VDD.t136 GND 0.025529f
C2322 VDD.t182 GND 0.025529f
C2323 VDD.n713 GND 0.163847f
C2324 VDD.n714 GND 0.154853f
C2325 VDD.t170 GND 0.221218f
C2326 VDD.n715 GND 0.162349f
C2327 VDD.n716 GND 0.344539f
C2328 VDD.t155 GND 0.222206f
C2329 VDD.t141 GND 0.025529f
C2330 VDD.t183 GND 0.025529f
C2331 VDD.n717 GND 0.163847f
C2332 VDD.n718 GND 0.290589f
C2333 VDD.t125 GND 0.025529f
C2334 VDD.t172 GND 0.025529f
C2335 VDD.n719 GND 0.163847f
C2336 VDD.n720 GND 0.154853f
C2337 VDD.t115 GND 0.025529f
C2338 VDD.t157 GND 0.025529f
C2339 VDD.n721 GND 0.163847f
C2340 VDD.n722 GND 0.154853f
C2341 VDD.t174 GND 0.025529f
C2342 VDD.t146 GND 0.025529f
C2343 VDD.n723 GND 0.163847f
C2344 VDD.n724 GND 0.154853f
C2345 VDD.t127 GND 0.221218f
C2346 VDD.n725 GND 0.162349f
C2347 VDD.n726 GND 0.303846f
C2348 VDD.n727 GND 1.71178f
C2349 VDD.n728 GND 0.19573f
C2350 VDD.n729 GND 0.007294f
C2351 VDD.n730 GND 0.009062f
C2352 VDD.n731 GND 0.643537f
C2353 VDD.n732 GND 0.009062f
C2354 VDD.n733 GND 0.007294f
C2355 VDD.n734 GND 0.009062f
C2356 VDD.n735 GND 0.007294f
C2357 VDD.n736 GND 0.009062f
C2358 VDD.n737 GND 0.703319f
C2359 VDD.t108 GND 0.35166f
C2360 VDD.n738 GND 0.009062f
C2361 VDD.n739 GND 0.007294f
C2362 VDD.n740 GND 0.009062f
C2363 VDD.n741 GND 0.007294f
C2364 VDD.n742 GND 0.009062f
C2365 VDD.t114 GND 0.35166f
C2366 VDD.n743 GND 0.009062f
C2367 VDD.n744 GND 0.007294f
C2368 VDD.n745 GND 0.009062f
C2369 VDD.n746 GND 0.007294f
C2370 VDD.n747 GND 0.009062f
C2371 VDD.n748 GND 0.404409f
C2372 VDD.n749 GND 0.531006f
C2373 VDD.n750 GND 0.009062f
C2374 VDD.n751 GND 0.007294f
C2375 VDD.n752 GND 0.009062f
C2376 VDD.n753 GND 0.007294f
C2377 VDD.n754 GND 0.009062f
C2378 VDD.n755 GND 0.636504f
C2379 VDD.n756 GND 0.009062f
C2380 VDD.n757 GND 0.007294f
C2381 VDD.n758 GND 0.009062f
C2382 VDD.n759 GND 0.007294f
C2383 VDD.n760 GND 0.009062f
C2384 VDD.n761 GND 0.703319f
C2385 VDD.t135 GND 0.35166f
C2386 VDD.n762 GND 0.009062f
C2387 VDD.n763 GND 0.007294f
C2388 VDD.n764 GND 0.009062f
C2389 VDD.n765 GND 0.007294f
C2390 VDD.n766 GND 0.009062f
C2391 VDD.t126 GND 0.35166f
C2392 VDD.n767 GND 0.009062f
C2393 VDD.n768 GND 0.007294f
C2394 VDD.n769 GND 0.009062f
C2395 VDD.n770 GND 0.007294f
C2396 VDD.n771 GND 0.009062f
C2397 VDD.n772 GND 0.703319f
C2398 VDD.n773 GND 0.538039f
C2399 VDD.n774 GND 0.009062f
C2400 VDD.n775 GND 0.007294f
C2401 VDD.n776 GND 0.009062f
C2402 VDD.n777 GND 0.007294f
C2403 VDD.n778 GND 0.009062f
C2404 VDD.n779 GND 0.460674f
C2405 VDD.n780 GND 0.009062f
C2406 VDD.n781 GND 0.007294f
C2407 VDD.n782 GND 0.02036f
C2408 VDD.n783 GND 0.006054f
C2409 VDD.n784 GND 0.02036f
C2410 VDD.n785 GND 0.903766f
C2411 VDD.t33 GND 0.35166f
C2412 VDD.n786 GND 0.02036f
C2413 VDD.n787 GND 0.006054f
C2414 VDD.n788 GND 0.009062f
C2415 VDD.n789 GND 0.007294f
C2416 VDD.n790 GND 0.009062f
C2417 VDD.n818 GND 0.02042f
C2418 VDD.n819 GND 0.009062f
C2419 VDD.n820 GND 0.007294f
C2420 VDD.n821 GND 0.009062f
C2421 VDD.n822 GND 0.009062f
C2422 VDD.n823 GND 0.009062f
C2423 VDD.n824 GND 0.009062f
C2424 VDD.n825 GND 0.009062f
C2425 VDD.n826 GND 0.007294f
C2426 VDD.n827 GND 0.009062f
C2427 VDD.n828 GND 0.009062f
C2428 VDD.n829 GND 0.009062f
C2429 VDD.n830 GND 0.009062f
C2430 VDD.n831 GND 0.009062f
C2431 VDD.n832 GND 0.007294f
C2432 VDD.n833 GND 0.009062f
C2433 VDD.n834 GND 0.009062f
C2434 VDD.n835 GND 0.009062f
C2435 VDD.n836 GND 0.009062f
C2436 VDD.n837 GND 0.009062f
C2437 VDD.n838 GND 0.007294f
C2438 VDD.n839 GND 0.009062f
C2439 VDD.n840 GND 0.009062f
C2440 VDD.n841 GND 0.009062f
C2441 VDD.n842 GND 0.009062f
C2442 VDD.n843 GND 0.007294f
C2443 VDD.n844 GND 0.009062f
C2444 VDD.n845 GND 0.009062f
C2445 VDD.n846 GND 0.009062f
C2446 VDD.n847 GND 0.009062f
C2447 VDD.n848 GND 0.009062f
C2448 VDD.n849 GND 0.007294f
C2449 VDD.n850 GND 0.009062f
C2450 VDD.n851 GND 0.009062f
C2451 VDD.n852 GND 0.009062f
C2452 VDD.n853 GND 0.009062f
C2453 VDD.n854 GND 0.009062f
C2454 VDD.n855 GND 0.007294f
C2455 VDD.n856 GND 0.009062f
C2456 VDD.n857 GND 0.009062f
C2457 VDD.n858 GND 0.009062f
C2458 VDD.n859 GND 0.009062f
C2459 VDD.n860 GND 0.009062f
C2460 VDD.n861 GND 0.007294f
C2461 VDD.n862 GND 0.009062f
C2462 VDD.n863 GND 0.009062f
C2463 VDD.n864 GND 0.009062f
C2464 VDD.n865 GND 0.009062f
C2465 VDD.n866 GND 0.009062f
C2466 VDD.n867 GND 0.007294f
C2467 VDD.n868 GND 0.009062f
C2468 VDD.n869 GND 0.009062f
C2469 VDD.n870 GND 0.009062f
C2470 VDD.n871 GND 0.009062f
C2471 VDD.n872 GND 0.007294f
C2472 VDD.n873 GND 0.009062f
C2473 VDD.n874 GND 0.009062f
C2474 VDD.n875 GND 0.009062f
C2475 VDD.n876 GND 0.009062f
C2476 VDD.n877 GND 0.009062f
C2477 VDD.n878 GND 0.007294f
C2478 VDD.n879 GND 0.009062f
C2479 VDD.n880 GND 0.009062f
C2480 VDD.n881 GND 0.009062f
C2481 VDD.n882 GND 0.009062f
C2482 VDD.n883 GND 0.009062f
C2483 VDD.n884 GND 0.007294f
C2484 VDD.n885 GND 0.009062f
C2485 VDD.n886 GND 0.009062f
C2486 VDD.n887 GND 0.009062f
C2487 VDD.n888 GND 0.009062f
C2488 VDD.n889 GND 0.009062f
C2489 VDD.n890 GND 0.007294f
C2490 VDD.n891 GND 0.009062f
C2491 VDD.n892 GND 0.009062f
C2492 VDD.n893 GND 0.009062f
C2493 VDD.n894 GND 0.009062f
C2494 VDD.n895 GND 0.009062f
C2495 VDD.n896 GND 0.007294f
C2496 VDD.n897 GND 0.02042f
C2497 VDD.n898 GND 0.009062f
C2498 VDD.n899 GND 0.003465f
C2499 VDD.t41 GND 0.18563f
C2500 VDD.t42 GND 0.194533f
C2501 VDD.t40 GND 0.271204f
C2502 VDD.n900 GND 0.091924f
C2503 VDD.n901 GND 0.052705f
C2504 VDD.n902 GND 0.011269f
C2505 VDD.n903 GND 0.003829f
C2506 VDD.n904 GND 0.009062f
C2507 VDD.n905 GND 0.009062f
C2508 VDD.n906 GND 0.009062f
C2509 VDD.n907 GND 0.007294f
C2510 VDD.n908 GND 0.007294f
C2511 VDD.n909 GND 0.007294f
C2512 VDD.n910 GND 0.009062f
C2513 VDD.n911 GND 0.009062f
C2514 VDD.n912 GND 0.009062f
C2515 VDD.n913 GND 0.007294f
C2516 VDD.n914 GND 0.007294f
C2517 VDD.n915 GND 0.007294f
C2518 VDD.n916 GND 0.009062f
C2519 VDD.n917 GND 0.009062f
C2520 VDD.n918 GND 0.009062f
C2521 VDD.n919 GND 0.007294f
C2522 VDD.n920 GND 0.007294f
C2523 VDD.n921 GND 0.007294f
C2524 VDD.n922 GND 0.009062f
C2525 VDD.n923 GND 0.009062f
C2526 VDD.n924 GND 0.009062f
C2527 VDD.n925 GND 0.007294f
C2528 VDD.n926 GND 0.007294f
C2529 VDD.n927 GND 0.007294f
C2530 VDD.n928 GND 0.009062f
C2531 VDD.n929 GND 0.009062f
C2532 VDD.n930 GND 0.009062f
C2533 VDD.n931 GND 0.007221f
C2534 VDD.n932 GND 0.009062f
C2535 VDD.t34 GND 0.18563f
C2536 VDD.t35 GND 0.194533f
C2537 VDD.t32 GND 0.271204f
C2538 VDD.n933 GND 0.091924f
C2539 VDD.n934 GND 0.052705f
C2540 VDD.n935 GND 0.014916f
C2541 VDD.n936 GND 0.00496f
C2542 VDD.n937 GND 0.009062f
C2543 VDD.n938 GND 0.009062f
C2544 VDD.n939 GND 0.009062f
C2545 VDD.n940 GND 0.007294f
C2546 VDD.n941 GND 0.007294f
C2547 VDD.n942 GND 0.007294f
C2548 VDD.n943 GND 0.009062f
C2549 VDD.n944 GND 0.009062f
C2550 VDD.n945 GND 0.009062f
C2551 VDD.n946 GND 0.007294f
C2552 VDD.n947 GND 0.007294f
C2553 VDD.n948 GND 0.007294f
C2554 VDD.n949 GND 0.009062f
C2555 VDD.n950 GND 0.009062f
C2556 VDD.n951 GND 0.009062f
C2557 VDD.n952 GND 0.007294f
C2558 VDD.n953 GND 0.007294f
C2559 VDD.n954 GND 0.007294f
C2560 VDD.n955 GND 0.009062f
C2561 VDD.n956 GND 0.009062f
C2562 VDD.n957 GND 0.009062f
C2563 VDD.n958 GND 0.007294f
C2564 VDD.n959 GND 0.007294f
C2565 VDD.n960 GND 0.007294f
C2566 VDD.n961 GND 0.009062f
C2567 VDD.n962 GND 0.009062f
C2568 VDD.n963 GND 0.009062f
C2569 VDD.n964 GND 0.00609f
C2570 VDD.n965 GND 0.009062f
C2571 VDD.t68 GND 0.18563f
C2572 VDD.t69 GND 0.194533f
C2573 VDD.t67 GND 0.271204f
C2574 VDD.n966 GND 0.091924f
C2575 VDD.n967 GND 0.052705f
C2576 VDD.n968 GND 0.014916f
C2577 VDD.n969 GND 0.00609f
C2578 VDD.n970 GND 0.009062f
C2579 VDD.n971 GND 0.009062f
C2580 VDD.n972 GND 0.009062f
C2581 VDD.n973 GND 0.007294f
C2582 VDD.n974 GND 0.007294f
C2583 VDD.n975 GND 0.007294f
C2584 VDD.n976 GND 0.009062f
C2585 VDD.n977 GND 0.009062f
C2586 VDD.n978 GND 0.009062f
C2587 VDD.n979 GND 0.007294f
C2588 VDD.n980 GND 0.007294f
C2589 VDD.n981 GND 0.007294f
C2590 VDD.n982 GND 0.009062f
C2591 VDD.n983 GND 0.009062f
C2592 VDD.n984 GND 0.009062f
C2593 VDD.n985 GND 0.007294f
C2594 VDD.n986 GND 0.007294f
C2595 VDD.n987 GND 0.007294f
C2596 VDD.n988 GND 0.009062f
C2597 VDD.n989 GND 0.009062f
C2598 VDD.n990 GND 0.009062f
C2599 VDD.n991 GND 0.007294f
C2600 VDD.n992 GND 0.009062f
C2601 VDD.n993 GND 1.52972f
C2602 VDD.n995 GND 0.02042f
C2603 VDD.n996 GND 0.006054f
C2604 VDD.n997 GND 0.02042f
C2605 VDD.n998 GND 0.02036f
C2606 VDD.n999 GND 0.009062f
C2607 VDD.n1000 GND 0.007294f
C2608 VDD.n1001 GND 0.009062f
C2609 VDD.n1002 GND 0.594305f
C2610 VDD.n1003 GND 0.009062f
C2611 VDD.n1004 GND 0.007294f
C2612 VDD.n1005 GND 0.009062f
C2613 VDD.n1006 GND 0.009062f
C2614 VDD.n1007 GND 0.009062f
C2615 VDD.n1008 GND 0.007294f
C2616 VDD.n1009 GND 0.009062f
C2617 VDD.n1010 GND 0.703319f
C2618 VDD.n1011 GND 0.009062f
C2619 VDD.n1012 GND 0.007294f
C2620 VDD.n1013 GND 0.009062f
C2621 VDD.n1014 GND 0.009062f
C2622 VDD.n1015 GND 0.009062f
C2623 VDD.n1016 GND 0.007294f
C2624 VDD.n1017 GND 0.009062f
C2625 VDD.n1018 GND 0.703319f
C2626 VDD.n1019 GND 0.009062f
C2627 VDD.n1020 GND 0.007294f
C2628 VDD.n1021 GND 0.009062f
C2629 VDD.n1022 GND 0.009062f
C2630 VDD.n1023 GND 0.009062f
C2631 VDD.n1024 GND 0.007294f
C2632 VDD.n1025 GND 0.009062f
C2633 VDD.n1026 GND 0.51694f
C2634 VDD.n1027 GND 0.009062f
C2635 VDD.n1028 GND 0.007294f
C2636 VDD.n1029 GND 0.009062f
C2637 VDD.n1030 GND 0.009062f
C2638 VDD.n1031 GND 0.009062f
C2639 VDD.n1032 GND 0.007294f
C2640 VDD.n1033 GND 0.009062f
C2641 VDD.n1034 GND 0.418475f
C2642 VDD.n1035 GND 0.009062f
C2643 VDD.n1036 GND 0.007294f
C2644 VDD.n1037 GND 0.009062f
C2645 VDD.n1038 GND 0.009062f
C2646 VDD.n1039 GND 0.009062f
C2647 VDD.n1040 GND 0.007294f
C2648 VDD.n1041 GND 0.009062f
C2649 VDD.t145 GND 0.35166f
C2650 VDD.n1042 GND 0.65057f
C2651 VDD.n1043 GND 0.009062f
C2652 VDD.n1044 GND 0.007294f
C2653 VDD.n1045 GND 0.009062f
C2654 VDD.n1046 GND 0.009062f
C2655 VDD.n1047 GND 0.009062f
C2656 VDD.n1048 GND 0.007294f
C2657 VDD.n1049 GND 0.009062f
C2658 VDD.n1050 GND 0.703319f
C2659 VDD.n1051 GND 0.009062f
C2660 VDD.n1052 GND 0.007294f
C2661 VDD.n1053 GND 0.009062f
C2662 VDD.n1054 GND 0.009062f
C2663 VDD.n1055 GND 0.009062f
C2664 VDD.n1056 GND 0.007294f
C2665 VDD.n1057 GND 0.009062f
C2666 VDD.n1058 GND 0.523973f
C2667 VDD.n1059 GND 0.009062f
C2668 VDD.n1060 GND 0.007294f
C2669 VDD.n1061 GND 0.009062f
C2670 VDD.n1062 GND 0.009062f
C2671 VDD.n1063 GND 0.006965f
C2672 VDD.n1064 GND 0.009062f
C2673 VDD.n1065 GND 0.007294f
C2674 VDD.n1066 GND 0.009062f
C2675 VDD.n1067 GND 0.411442f
C2676 VDD.n1068 GND 0.009062f
C2677 VDD.n1069 GND 0.007294f
C2678 VDD.n1070 GND 0.009062f
C2679 VDD.n1071 GND 0.009062f
C2680 VDD.n1072 GND 0.009062f
C2681 VDD.n1073 GND 0.007294f
C2682 VDD.n1074 GND 0.009062f
C2683 VDD.t124 GND 0.35166f
C2684 VDD.n1075 GND 0.643537f
C2685 VDD.n1076 GND 0.009062f
C2686 VDD.n1077 GND 0.007294f
C2687 VDD.n1078 GND 0.006965f
C2688 VDD.n1079 GND 0.009062f
C2689 VDD.n1080 GND 0.009062f
C2690 VDD.n1081 GND 0.007294f
C2691 VDD.n1082 GND 0.009062f
C2692 VDD.n1083 GND 0.703319f
C2693 VDD.n1084 GND 0.009062f
C2694 VDD.n1085 GND 0.007294f
C2695 VDD.n1086 GND 0.009062f
C2696 VDD.n1087 GND 0.009062f
C2697 VDD.n1088 GND 0.009062f
C2698 VDD.n1089 GND 0.007294f
C2699 VDD.n1090 GND 0.009062f
C2700 VDD.n1091 GND 0.531006f
C2701 VDD.n1092 GND 0.009062f
C2702 VDD.n1093 GND 0.007294f
C2703 VDD.n1094 GND 0.009062f
C2704 VDD.n1095 GND 0.009062f
C2705 VDD.n1096 GND 0.009062f
C2706 VDD.n1097 GND 0.007294f
C2707 VDD.n1098 GND 0.009062f
C2708 VDD.n1099 GND 0.404409f
C2709 VDD.n1100 GND 0.009062f
C2710 VDD.n1101 GND 0.007294f
C2711 VDD.n1102 GND 0.009062f
C2712 VDD.n1103 GND 0.009062f
C2713 VDD.n1104 GND 0.009062f
C2714 VDD.n1105 GND 0.007294f
C2715 VDD.n1106 GND 0.009062f
C2716 VDD.t147 GND 0.35166f
C2717 VDD.n1107 GND 0.636504f
C2718 VDD.n1108 GND 0.009062f
C2719 VDD.n1109 GND 0.007294f
C2720 VDD.n1110 GND 0.009062f
C2721 VDD.n1111 GND 0.009062f
C2722 VDD.n1112 GND 0.009062f
C2723 VDD.n1113 GND 0.007294f
C2724 VDD.n1114 GND 0.009062f
C2725 VDD.n1115 GND 0.703319f
C2726 VDD.n1116 GND 0.009062f
C2727 VDD.n1117 GND 0.007294f
C2728 VDD.n1118 GND 0.009062f
C2729 VDD.n1119 GND 0.009062f
C2730 VDD.n1120 GND 0.009062f
C2731 VDD.n1121 GND 0.007294f
C2732 VDD.n1122 GND 0.009062f
C2733 VDD.n1123 GND 0.538039f
C2734 VDD.n1124 GND 0.009062f
C2735 VDD.n1125 GND 0.007294f
C2736 VDD.n1126 GND 0.009062f
C2737 VDD.n1127 GND 0.009062f
C2738 VDD.n1128 GND 0.009062f
C2739 VDD.n1129 GND 0.007294f
C2740 VDD.n1130 GND 0.009062f
C2741 VDD.n1131 GND 0.703319f
C2742 VDD.n1132 GND 0.009062f
C2743 VDD.n1133 GND 0.007294f
C2744 VDD.n1134 GND 0.009062f
C2745 VDD.n1135 GND 0.009062f
C2746 VDD.n1136 GND 0.009062f
C2747 VDD.n1137 GND 0.007294f
C2748 VDD.n1138 GND 0.009062f
C2749 VDD.t22 GND 0.35166f
C2750 VDD.n1139 GND 0.460674f
C2751 VDD.n1140 GND 0.009062f
C2752 VDD.n1141 GND 0.007294f
C2753 VDD.n1142 GND 0.009062f
C2754 VDD.n1143 GND 0.009062f
C2755 VDD.n1144 GND 0.009062f
C2756 VDD.n1145 GND 0.007294f
C2757 VDD.n1147 GND 0.009062f
C2758 VDD.n1148 GND 0.009062f
C2759 VDD.n1149 GND 0.009062f
C2760 VDD.n1150 GND 0.009062f
C2761 VDD.n1151 GND 0.009062f
C2762 VDD.n1152 GND 0.007294f
C2763 VDD.n1154 GND 0.009062f
C2764 VDD.n1155 GND 0.007294f
C2765 VDD.n1156 GND 0.007794f
C2766 VDD.n1157 GND 0.0058f
C2767 VDD.n1158 GND 0.007294f
C2768 VDD.n1159 GND 0.007294f
C2769 VDD.n1161 GND 0.009062f
C2770 VDD.n1162 GND 0.007294f
C2771 VDD.n1163 GND 0.009062f
C2772 VDD.n1164 GND 0.009062f
C2773 VDD.n1165 GND 0.009062f
C2774 VDD.n1166 GND 0.009062f
C2775 VDD.n1167 GND 0.009062f
C2776 VDD.n1168 GND 0.00609f
C2777 VDD.n1170 GND 0.009062f
C2778 VDD.n1171 GND 0.00609f
C2779 VDD.t24 GND 0.18563f
C2780 VDD.t23 GND 0.194533f
C2781 VDD.t21 GND 0.271204f
C2782 VDD.n1172 GND 0.091924f
C2783 VDD.n1173 GND 0.052705f
C2784 VDD.n1174 GND 0.009062f
C2785 VDD.n1175 GND 0.009062f
C2786 VDD.n1176 GND 0.007294f
C2787 VDD.n1178 GND 0.009062f
C2788 VDD.n1179 GND 0.009062f
C2789 VDD.n1180 GND 0.009062f
C2790 VDD.n1181 GND 0.009062f
C2791 VDD.n1182 GND 0.007294f
C2792 VDD.n1184 GND 0.009062f
C2793 VDD.n1185 GND 0.009062f
C2794 VDD.n1186 GND 0.009062f
C2795 VDD.n1187 GND 0.009062f
C2796 VDD.n1188 GND 0.009062f
C2797 VDD.n1189 GND 0.007294f
C2798 VDD.n1191 GND 0.009062f
C2799 VDD.n1192 GND 0.009062f
C2800 VDD.n1193 GND 0.009062f
C2801 VDD.n1194 GND 0.009062f
C2802 VDD.n1195 GND 0.009062f
C2803 VDD.n1196 GND 0.007294f
C2804 VDD.n1198 GND 0.009062f
C2805 VDD.n1199 GND 0.009062f
C2806 VDD.n1200 GND 0.009062f
C2807 VDD.n1201 GND 0.009062f
C2808 VDD.n1202 GND 0.009062f
C2809 VDD.n1203 GND 0.00496f
C2810 VDD.n1205 GND 0.009062f
C2811 VDD.n1206 GND 0.007221f
C2812 VDD.t62 GND 0.18563f
C2813 VDD.t61 GND 0.194533f
C2814 VDD.t60 GND 0.271204f
C2815 VDD.n1207 GND 0.091924f
C2816 VDD.n1208 GND 0.052705f
C2817 VDD.n1209 GND 0.009062f
C2818 VDD.n1210 GND 0.009062f
C2819 VDD.n1211 GND 0.007294f
C2820 VDD.n1213 GND 0.009062f
C2821 VDD.n1214 GND 0.009062f
C2822 VDD.n1215 GND 0.009062f
C2823 VDD.n1216 GND 0.009062f
C2824 VDD.n1217 GND 0.007294f
C2825 VDD.n1219 GND 0.009062f
C2826 VDD.n1220 GND 0.009062f
C2827 VDD.n1221 GND 0.009062f
C2828 VDD.n1223 GND 0.007294f
C2829 VDD.n1225 GND 0.009062f
C2830 VDD.n1226 GND 0.007294f
C2831 VDD.n1227 GND 0.009062f
C2832 VDD.n1229 GND 0.009062f
C2833 VDD.n1230 GND 0.009062f
C2834 VDD.n1231 GND 0.007294f
C2835 VDD.n1232 GND 0.007294f
C2836 VDD.n1233 GND 0.007294f
C2837 VDD.n1234 GND 0.009062f
C2838 VDD.n1236 GND 0.009062f
C2839 VDD.n1237 GND 0.009062f
C2840 VDD.n1238 GND 0.007294f
C2841 VDD.n1239 GND 0.007294f
C2842 VDD.n1240 GND 0.007294f
C2843 VDD.n1241 GND 0.009062f
C2844 VDD.n1243 GND 0.009062f
C2845 VDD.n1244 GND 0.009062f
C2846 VDD.n1245 GND 0.007294f
C2847 VDD.n1246 GND 0.009062f
C2848 VDD.n1247 GND 0.009062f
C2849 VDD.n1248 GND 0.009062f
C2850 VDD.n1249 GND 0.014916f
C2851 VDD.n1250 GND 0.009062f
C2852 VDD.n1252 GND 0.009062f
C2853 VDD.n1253 GND 0.009062f
C2854 VDD.n1254 GND 0.007294f
C2855 VDD.n1255 GND 0.007294f
C2856 VDD.n1256 GND 0.007294f
C2857 VDD.n1257 GND 0.009062f
C2858 VDD.n1259 GND 0.009062f
C2859 VDD.n1260 GND 0.009062f
C2860 VDD.n1261 GND 0.007294f
C2861 VDD.n1262 GND 0.007294f
C2862 VDD.n1263 GND 0.007294f
C2863 VDD.n1264 GND 0.009062f
C2864 VDD.n1266 GND 0.009062f
C2865 VDD.n1267 GND 0.009062f
C2866 VDD.n1268 GND 0.007294f
C2867 VDD.n1269 GND 0.007294f
C2868 VDD.n1270 GND 0.007294f
C2869 VDD.n1271 GND 0.009062f
C2870 VDD.n1273 GND 0.009062f
C2871 VDD.n1274 GND 0.009062f
C2872 VDD.n1275 GND 0.007294f
C2873 VDD.n1276 GND 0.007294f
C2874 VDD.n1277 GND 0.007294f
C2875 VDD.n1278 GND 0.009062f
C2876 VDD.n1280 GND 0.009062f
C2877 VDD.n1281 GND 0.009062f
C2878 VDD.n1282 GND 0.007294f
C2879 VDD.n1283 GND 0.009062f
C2880 VDD.n1284 GND 0.009062f
C2881 VDD.n1285 GND 0.009062f
C2882 VDD.n1286 GND 0.014916f
C2883 VDD.n1287 GND 0.009062f
C2884 VDD.n1289 GND 0.009062f
C2885 VDD.n1290 GND 0.009062f
C2886 VDD.n1291 GND 0.007294f
C2887 VDD.n1292 GND 0.007294f
C2888 VDD.n1293 GND 0.007294f
C2889 VDD.n1294 GND 0.009062f
C2890 VDD.n1296 GND 0.009062f
C2891 VDD.n1297 GND 0.009062f
C2892 VDD.n1299 GND 0.009062f
C2893 VDD.n1300 GND 0.007294f
C2894 VDD.n1302 GND 0.006162f
C2895 VDD.n1303 GND 0.006162f
C2896 VDD.n1304 GND 0.006162f
C2897 VDD.n1305 GND 0.006162f
C2898 VDD.n1306 GND 0.006162f
C2899 VDD.n1307 GND 0.006162f
C2900 VDD.n1308 GND 0.006162f
C2901 VDD.n1310 GND 0.006162f
C2902 VDD.n1311 GND 0.006162f
C2903 VDD.n1313 GND 0.006162f
C2904 VDD.n1314 GND 0.006162f
C2905 VDD.n1315 GND 0.006162f
C2906 VDD.n1316 GND 0.006162f
C2907 VDD.n1317 GND 0.006162f
C2908 VDD.n1319 GND 0.006162f
C2909 VDD.n1321 GND 0.006162f
C2910 VDD.n1322 GND 0.006162f
C2911 VDD.n1323 GND 0.006162f
C2912 VDD.n1324 GND 0.006162f
C2913 VDD.n1325 GND 0.006162f
C2914 VDD.n1327 GND 0.006162f
C2915 VDD.n1329 GND 0.006162f
C2916 VDD.n1330 GND 0.006162f
C2917 VDD.n1331 GND 0.004848f
C2918 VDD.n1332 GND 0.006162f
C2919 VDD.t95 GND 0.122823f
C2920 VDD.t96 GND 0.131225f
C2921 VDD.t94 GND 0.198505f
C2922 VDD.n1333 GND 0.075862f
C2923 VDD.n1334 GND 0.050543f
C2924 VDD.n1335 GND 0.008807f
C2925 VDD.n1336 GND 0.006162f
C2926 VDD.n1337 GND 0.006162f
C2927 VDD.n1338 GND 0.006162f
C2928 VDD.n1339 GND 0.006162f
C2929 VDD.n1340 GND 0.006162f
C2930 VDD.n1341 GND 0.006162f
C2931 VDD.n1342 GND 0.006162f
C2932 VDD.n1343 GND 0.006162f
C2933 VDD.n1344 GND 0.006162f
C2934 VDD.n1345 GND 0.006162f
C2935 VDD.n1346 GND 0.006162f
C2936 VDD.n1347 GND 0.006162f
C2937 VDD.t72 GND 0.122823f
C2938 VDD.t73 GND 0.131225f
C2939 VDD.t70 GND 0.198505f
C2940 VDD.n1348 GND 0.075862f
C2941 VDD.n1349 GND 0.050543f
C2942 VDD.n1350 GND 0.006162f
C2943 VDD.n1351 GND 0.006162f
C2944 VDD.n1352 GND 0.006162f
C2945 VDD.n1354 GND 0.006162f
C2946 VDD.n1356 GND 0.006162f
C2947 VDD.n1357 GND 0.006162f
C2948 VDD.n1358 GND 0.006162f
C2949 VDD.n1359 GND 0.006162f
C2950 VDD.n1360 GND 0.006162f
C2951 VDD.n1362 GND 0.006162f
C2952 VDD.n1364 GND 0.006162f
C2953 VDD.n1365 GND 0.006162f
C2954 VDD.n1366 GND 0.004848f
C2955 VDD.n1367 GND 0.008807f
C2956 VDD.n1368 GND 0.004395f
C2957 VDD.n1369 GND 0.006162f
C2958 VDD.n1371 GND 0.006162f
C2959 VDD.n1372 GND 0.014791f
C2960 VDD.n1373 GND 0.014791f
C2961 VDD.n1374 GND 0.014027f
C2962 VDD.n1375 GND 0.006162f
C2963 VDD.n1376 GND 0.006162f
C2964 VDD.n1377 GND 0.006162f
C2965 VDD.n1378 GND 0.006162f
C2966 VDD.n1379 GND 0.006162f
C2967 VDD.n1380 GND 0.006162f
C2968 VDD.n1381 GND 0.006162f
C2969 VDD.n1382 GND 0.006162f
C2970 VDD.n1383 GND 0.006162f
C2971 VDD.n1384 GND 0.006162f
C2972 VDD.n1385 GND 0.006162f
C2973 VDD.n1386 GND 0.006162f
C2974 VDD.n1387 GND 0.006162f
C2975 VDD.n1388 GND 0.006162f
C2976 VDD.n1389 GND 0.006162f
C2977 VDD.n1390 GND 0.006162f
C2978 VDD.n1391 GND 0.006162f
C2979 VDD.n1392 GND 0.006162f
C2980 VDD.n1393 GND 0.006162f
C2981 VDD.n1394 GND 0.006162f
C2982 VDD.n1395 GND 0.006162f
C2983 VDD.n1396 GND 0.006162f
C2984 VDD.n1397 GND 0.006162f
C2985 VDD.n1398 GND 0.006162f
C2986 VDD.n1399 GND 0.006162f
C2987 VDD.n1400 GND 0.006162f
C2988 VDD.n1401 GND 0.006162f
C2989 VDD.n1402 GND 0.006162f
C2990 VDD.n1403 GND 0.006162f
C2991 VDD.n1404 GND 0.006162f
C2992 VDD.n1405 GND 0.006162f
C2993 VDD.n1406 GND 0.006162f
C2994 VDD.n1407 GND 0.006162f
C2995 VDD.n1408 GND 0.006162f
C2996 VDD.n1409 GND 0.006162f
C2997 VDD.n1410 GND 0.006162f
C2998 VDD.n1411 GND 0.006162f
C2999 VDD.n1412 GND 0.006162f
C3000 VDD.n1413 GND 0.006162f
C3001 VDD.n1414 GND 0.32001f
C3002 VDD.n1415 GND 0.006162f
C3003 VDD.n1416 GND 0.006162f
C3004 VDD.n1417 GND 0.006162f
C3005 VDD.n1418 GND 0.006162f
C3006 VDD.n1419 GND 0.006162f
C3007 VDD.n1420 GND 0.006162f
C3008 VDD.n1421 GND 0.006162f
C3009 VDD.n1422 GND 0.006162f
C3010 VDD.n1423 GND 0.006162f
C3011 VDD.n1424 GND 0.006162f
C3012 VDD.n1425 GND 0.006162f
C3013 VDD.n1426 GND 0.006162f
C3014 VDD.n1427 GND 0.006162f
C3015 VDD.n1428 GND 0.006162f
C3016 VDD.n1429 GND 0.006162f
C3017 VDD.n1430 GND 0.006162f
C3018 VDD.n1431 GND 0.006162f
C3019 VDD.n1432 GND 0.006162f
C3020 VDD.n1433 GND 0.006162f
C3021 VDD.n1434 GND 0.006162f
C3022 VDD.n1435 GND 0.006162f
C3023 VDD.n1436 GND 0.006162f
C3024 VDD.n1437 GND 0.006162f
C3025 VDD.n1438 GND 0.006162f
C3026 VDD.n1439 GND 0.006162f
C3027 VDD.n1440 GND 0.006162f
C3028 VDD.n1441 GND 0.014027f
C3029 VDD.n1443 GND 0.014791f
C3030 VDD.n1444 GND 0.014791f
C3031 VDD.n1445 GND 0.006162f
C3032 VDD.n1446 GND 0.004395f
C3033 VDD.n1447 GND 0.006162f
C3034 VDD.n1449 GND 0.006162f
C3035 VDD.n1451 GND 0.006162f
C3036 VDD.n1452 GND 0.006162f
C3037 VDD.n1453 GND 0.006162f
C3038 VDD.n1454 GND 0.006162f
C3039 VDD.n1455 GND 0.006162f
C3040 VDD.n1457 GND 0.006162f
C3041 VDD.n1458 GND 0.006162f
C3042 VDD.n1459 GND 0.006162f
C3043 VDD.n1460 GND 0.006162f
C3044 VDD.n1461 GND 0.006162f
C3045 VDD.n1462 GND 0.006162f
C3046 VDD.n1464 GND 0.006162f
C3047 VDD.n1465 GND 0.014608f
C3048 VDD.n1466 GND 0.439031f
C3049 VDD.n1468 GND 0.007294f
C3050 VDD.n1469 GND 0.009062f
C3051 VDD.n1471 GND 0.009062f
C3052 VDD.n1472 GND 0.009062f
C3053 VDD.n1473 GND 0.007294f
C3054 VDD.n1474 GND 0.007294f
C3055 VDD.n1475 GND 0.007294f
C3056 VDD.n1476 GND 0.009062f
C3057 VDD.n1478 GND 0.009062f
C3058 VDD.n1479 GND 0.009062f
C3059 VDD.n1480 GND 0.007294f
C3060 VDD.n1481 GND 0.006054f
C3061 VDD.n1482 GND 0.02042f
C3062 VDD.n1483 GND 0.02036f
C3063 VDD.n1484 GND 0.006054f
C3064 VDD.n1485 GND 0.02036f
C3065 VDD.n1486 GND 0.903766f
C3066 VDD.n1487 GND 0.02036f
C3067 VDD.n1488 GND 0.006054f
C3068 VDD.n1489 GND 0.02036f
C3069 VDD.n1490 GND 0.02042f
C3070 VDD.n1491 GND 0.003465f
C3071 VDD.t31 GND 0.18563f
C3072 VDD.t30 GND 0.194533f
C3073 VDD.t29 GND 0.271204f
C3074 VDD.n1492 GND 0.091924f
C3075 VDD.n1493 GND 0.052705f
C3076 VDD.n1494 GND 0.011269f
C3077 VDD.n1495 GND 0.003829f
C3078 VDD.n1496 GND 0.007294f
C3079 VDD.n1497 GND 0.009062f
C3080 VDD.n1498 GND 0.009062f
C3081 VDD.n1499 GND 0.009062f
C3082 VDD.n1500 GND 0.007294f
C3083 VDD.n1501 GND 0.007294f
C3084 VDD.n1502 GND 0.007294f
C3085 VDD.n1503 GND 0.007794f
C3086 VDD.n1504 GND 0.439031f
C3087 VDD.n1505 GND 0.014608f
C3088 VDD.n1506 GND 0.006162f
C3089 VDD.n1508 GND 0.006162f
C3090 VDD.n1510 GND 0.006162f
C3091 VDD.n1511 GND 0.006162f
C3092 VDD.n1512 GND 0.006162f
C3093 VDD.n1513 GND 0.006162f
C3094 VDD.n1514 GND 0.006162f
C3095 VDD.n1516 GND 0.006162f
C3096 VDD.n1518 GND 0.006162f
C3097 VDD.n1519 GND 0.006162f
C3098 VDD.n1520 GND 0.006162f
C3099 VDD.n1521 GND 0.006162f
C3100 VDD.n1522 GND 0.006162f
C3101 VDD.n1524 GND 0.006162f
C3102 VDD.n1526 GND 0.006162f
C3103 VDD.n1527 GND 0.006162f
C3104 VDD.n1528 GND 0.006842f
C3105 VDD.n1529 GND 0.028657f
C3106 VDD.n1530 GND 0.00879f
C3107 VDD.n1531 GND 0.014027f
C3108 VDD.n1532 GND 0.68222f
C3109 VDD.n1533 GND 0.014027f
C3110 VDD.n1534 GND 0.014027f
C3111 VDD.n1535 GND 0.006162f
C3112 VDD.n1536 GND 0.006162f
C3113 VDD.n1537 GND 0.006162f
C3114 VDD.n1538 GND 0.478257f
C3115 VDD.n1539 GND 0.006162f
C3116 VDD.n1540 GND 0.006162f
C3117 VDD.n1541 GND 0.006162f
C3118 VDD.n1542 GND 0.006162f
C3119 VDD.n1543 GND 0.006162f
C3120 VDD.n1544 GND 0.446608f
C3121 VDD.n1545 GND 0.006162f
C3122 VDD.n1546 GND 0.006162f
C3123 VDD.n1547 GND 0.006162f
C3124 VDD.n1548 GND 0.006162f
C3125 VDD.n1549 GND 0.006162f
C3126 VDD.n1550 GND 0.478257f
C3127 VDD.n1551 GND 0.006162f
C3128 VDD.n1552 GND 0.006162f
C3129 VDD.n1553 GND 0.006162f
C3130 VDD.n1554 GND 0.006162f
C3131 VDD.n1555 GND 0.006162f
C3132 VDD.n1556 GND 0.429025f
C3133 VDD.n1557 GND 0.006162f
C3134 VDD.n1558 GND 0.006162f
C3135 VDD.n1559 GND 0.006162f
C3136 VDD.n1560 GND 0.006162f
C3137 VDD.n1561 GND 0.006162f
C3138 VDD.n1562 GND 0.270778f
C3139 VDD.n1563 GND 0.006162f
C3140 VDD.n1564 GND 0.006162f
C3141 VDD.n1565 GND 0.006162f
C3142 VDD.n1566 GND 0.006162f
C3143 VDD.n1567 GND 0.006162f
C3144 VDD.n1568 GND 0.407925f
C3145 VDD.n1569 GND 0.006162f
C3146 VDD.n1570 GND 0.006162f
C3147 VDD.n1571 GND 0.006162f
C3148 VDD.n1572 GND 0.006162f
C3149 VDD.n1573 GND 0.006162f
C3150 VDD.n1574 GND 0.249678f
C3151 VDD.n1575 GND 0.006162f
C3152 VDD.n1576 GND 0.006162f
C3153 VDD.n1577 GND 0.006162f
C3154 VDD.n1578 GND 0.006162f
C3155 VDD.n1579 GND 0.006162f
C3156 VDD.n1580 GND 0.386826f
C3157 VDD.n1581 GND 0.006162f
C3158 VDD.n1582 GND 0.006162f
C3159 VDD.n1583 GND 0.006162f
C3160 VDD.n1584 GND 0.006162f
C3161 VDD.n1585 GND 0.006162f
C3162 VDD.n1586 GND 0.249678f
C3163 VDD.n1587 GND 0.006162f
C3164 VDD.n1588 GND 0.006162f
C3165 VDD.n1589 GND 0.006162f
C3166 VDD.n1590 GND 0.006162f
C3167 VDD.n1591 GND 0.006162f
C3168 VDD.n1592 GND 0.478257f
C3169 VDD.n1593 GND 0.006162f
C3170 VDD.n1594 GND 0.006162f
C3171 VDD.n1595 GND 0.006162f
C3172 VDD.n1596 GND 0.006162f
C3173 VDD.n1597 GND 0.006162f
C3174 VDD.n1598 GND 0.18638f
C3175 VDD.n1599 GND 0.006162f
C3176 VDD.n1600 GND 0.006162f
C3177 VDD.n1601 GND 0.006162f
C3178 VDD.n1602 GND 0.006162f
C3179 VDD.n1603 GND 0.006162f
C3180 VDD.n1604 GND 0.006162f
C3181 VDD.n1605 GND 0.006162f
C3182 VDD.n1606 GND 0.006162f
C3183 VDD.n1607 GND 0.006162f
C3184 VDD.n1608 GND 0.478257f
C3185 VDD.n1609 GND 0.006162f
C3186 VDD.n1610 GND 0.006162f
C3187 VDD.n1611 GND 0.006162f
C3188 VDD.n1612 GND 0.006162f
C3189 VDD.n1613 GND 0.006162f
C3190 VDD.n1614 GND 0.006162f
C3191 VDD.n1615 GND 0.372759f
C3192 VDD.n1616 GND 0.006162f
C3193 VDD.n1617 GND 0.006162f
C3194 VDD.n1618 GND 0.006162f
C3195 VDD.n1619 GND 0.006162f
C3196 VDD.n1620 GND 0.006162f
C3197 VDD.n1621 GND 0.006162f
C3198 VDD.n1622 GND 0.006162f
C3199 VDD.n1623 GND 0.474741f
C3200 VDD.n1624 GND 0.006162f
C3201 VDD.n1625 GND 0.006162f
C3202 VDD.n1626 GND 0.006162f
C3203 VDD.n1627 GND 0.006162f
C3204 VDD.n1628 GND 0.006162f
C3205 VDD.n1629 GND 0.006162f
C3206 VDD.n1630 GND 0.014027f
C3207 VDD.n1631 GND 0.014756f
C3208 VDD.n1632 GND 0.014062f
C3209 VDD.n1633 GND 0.006162f
C3210 VDD.n1634 GND 0.006162f
C3211 VDD.n1635 GND 0.004395f
C3212 VDD.n1636 GND 0.006162f
C3213 VDD.n1637 GND 0.006162f
C3214 VDD.n1638 GND 0.004848f
C3215 VDD.n1639 GND 0.006162f
C3216 VDD.n1640 GND 0.006162f
C3217 VDD.n1641 GND 0.006162f
C3218 VDD.n1642 GND 0.006162f
C3219 VDD.n1643 GND 0.006162f
C3220 VDD.n1644 GND 0.006162f
C3221 VDD.n1645 GND 0.006162f
C3222 VDD.n1646 GND 0.006162f
C3223 VDD.n1647 GND 0.006162f
C3224 VDD.n1648 GND 0.006162f
C3225 VDD.n1649 GND 0.006162f
C3226 VDD.n1650 GND 0.006162f
C3227 VDD.n1651 GND 0.006162f
C3228 VDD.n1652 GND 0.006162f
C3229 VDD.n1653 GND 0.006162f
C3230 VDD.n1654 GND 0.006162f
C3231 VDD.n1655 GND 0.006162f
C3232 VDD.n1656 GND 0.006162f
C3233 VDD.n1657 GND 0.006162f
C3234 VDD.n1658 GND 0.006162f
C3235 VDD.n1659 GND 0.006162f
C3236 VDD.n1660 GND 0.006162f
C3237 VDD.n1661 GND 0.006162f
C3238 VDD.n1662 GND 0.006162f
C3239 VDD.n1663 GND 0.006162f
C3240 VDD.n1664 GND 0.006162f
C3241 VDD.n1665 GND 0.006162f
C3242 VDD.n1666 GND 0.006162f
C3243 VDD.n1667 GND 0.006162f
C3244 VDD.n1668 GND 0.006162f
C3245 VDD.n1669 GND 0.006162f
C3246 VDD.n1670 GND 0.006162f
C3247 VDD.n1671 GND 0.006162f
C3248 VDD.n1672 GND 0.006162f
C3249 VDD.n1673 GND 0.006162f
C3250 VDD.n1674 GND 0.006162f
C3251 VDD.n1675 GND 0.014791f
C3252 VDD.n1676 GND 0.014791f
C3253 VDD.n1677 GND 0.014027f
C3254 VDD.n1678 GND 0.014027f
C3255 VDD.n1679 GND 0.006162f
C3256 VDD.n1680 GND 0.006162f
C3257 VDD.n1681 GND 0.006162f
C3258 VDD.n1682 GND 0.006162f
C3259 VDD.n1683 GND 0.242645f
C3260 VDD.n1684 GND 0.006162f
C3261 VDD.n1685 GND 0.006162f
C3262 VDD.n1686 GND 0.006162f
C3263 VDD.n1687 GND 0.006162f
C3264 VDD.n1688 GND 0.006162f
C3265 VDD.n1689 GND 0.365726f
C3266 VDD.n1690 GND 0.006162f
C3267 VDD.n1691 GND 0.014027f
C3268 VDD.n1692 GND 0.014791f
C3269 VDD.n1693 GND 0.014062f
C3270 VDD.n1694 GND 0.006162f
C3271 VDD.n1695 GND 0.006162f
C3272 VDD.n1696 GND 0.006162f
C3273 VDD.n1697 GND 0.004395f
C3274 VDD.n1698 GND 0.008807f
C3275 VDD.n1699 GND 0.004848f
C3276 VDD.n1700 GND 0.006162f
C3277 VDD.n1701 GND 0.006162f
C3278 VDD.n1702 GND 0.006162f
C3279 VDD.n1703 GND 0.006162f
C3280 VDD.n1704 GND 0.006162f
C3281 VDD.n1705 GND 0.006162f
C3282 VDD.n1706 GND 0.006162f
C3283 VDD.n1707 GND 0.006162f
C3284 VDD.n1708 GND 0.006162f
C3285 VDD.n1709 GND 0.006162f
C3286 VDD.n1710 GND 0.006162f
C3287 VDD.n1711 GND 0.006162f
C3288 VDD.n1712 GND 0.006162f
C3289 VDD.n1713 GND 0.006162f
C3290 VDD.n1714 GND 0.006162f
C3291 VDD.n1715 GND 0.006162f
C3292 VDD.n1716 GND 0.006162f
C3293 VDD.n1717 GND 0.006162f
C3294 VDD.n1718 GND 0.006162f
C3295 VDD.n1719 GND 0.006162f
C3296 VDD.n1720 GND 0.006162f
C3297 VDD.n1721 GND 0.006162f
C3298 VDD.n1722 GND 0.006162f
C3299 VDD.n1723 GND 0.006162f
C3300 VDD.n1724 GND 0.006162f
C3301 VDD.n1725 GND 0.006162f
C3302 VDD.n1726 GND 0.006162f
C3303 VDD.n1727 GND 0.006162f
C3304 VDD.n1728 GND 0.006162f
C3305 VDD.n1729 GND 0.006162f
C3306 VDD.n1730 GND 0.006162f
C3307 VDD.n1731 GND 0.006162f
C3308 VDD.n1732 GND 0.006162f
C3309 VDD.n1733 GND 0.006162f
C3310 VDD.n1734 GND 0.006162f
C3311 VDD.n1735 GND 0.006162f
C3312 VDD.n1736 GND 0.014791f
C3313 VDD.n1737 GND 0.014791f
C3314 VDD.n1738 GND 0.569689f
C3315 VDD.t12 GND 2.42645f
C3316 VDD.t192 GND 2.42645f
C3317 VDD.n1760 GND 0.014791f
C3318 VDD.n1761 GND 0.006162f
C3319 VDD.t79 GND 0.122823f
C3320 VDD.t80 GND 0.131225f
C3321 VDD.t77 GND 0.198505f
C3322 VDD.n1762 GND 0.075862f
C3323 VDD.n1763 GND 0.050543f
C3324 VDD.n1764 GND 0.006162f
C3325 VDD.n1765 GND 0.006162f
C3326 VDD.n1766 GND 0.006162f
C3327 VDD.n1767 GND 0.006162f
C3328 VDD.n1768 GND 0.006162f
C3329 VDD.n1769 GND 0.006162f
C3330 VDD.n1770 GND 0.006162f
C3331 VDD.n1771 GND 0.006162f
C3332 VDD.n1772 GND 0.006162f
C3333 VDD.n1773 GND 0.006162f
C3334 VDD.n1774 GND 0.006162f
C3335 VDD.n1775 GND 0.006162f
C3336 VDD.n1776 GND 0.006162f
C3337 VDD.n1777 GND 0.006162f
C3338 VDD.n1778 GND 0.006162f
C3339 VDD.n1779 GND 0.006162f
C3340 VDD.n1780 GND 0.006162f
C3341 VDD.n1781 GND 0.006162f
C3342 VDD.n1782 GND 0.006162f
C3343 VDD.n1783 GND 0.006162f
C3344 VDD.n1784 GND 0.006162f
C3345 VDD.n1785 GND 0.006162f
C3346 VDD.n1786 GND 0.006162f
C3347 VDD.n1787 GND 0.006162f
C3348 VDD.n1788 GND 0.006162f
C3349 VDD.n1789 GND 0.006162f
C3350 VDD.t86 GND 0.122823f
C3351 VDD.t87 GND 0.131225f
C3352 VDD.t85 GND 0.198505f
C3353 VDD.n1790 GND 0.075862f
C3354 VDD.n1791 GND 0.050543f
C3355 VDD.n1792 GND 0.008807f
C3356 VDD.n1793 GND 0.014791f
C3357 VDD.n1794 GND 0.014791f
C3358 VDD.n1795 GND 0.006162f
C3359 VDD.n1796 GND 0.006162f
C3360 VDD.n1797 GND 0.006162f
C3361 VDD.n1798 GND 0.006162f
C3362 VDD.n1799 GND 0.006162f
C3363 VDD.n1800 GND 0.006162f
C3364 VDD.n1801 GND 0.006162f
C3365 VDD.n1802 GND 0.006162f
C3366 VDD.n1803 GND 0.006162f
C3367 VDD.n1804 GND 0.006162f
C3368 VDD.n1805 GND 0.006162f
C3369 VDD.n1806 GND 0.006162f
C3370 VDD.n1807 GND 0.006162f
C3371 VDD.n1808 GND 0.006162f
C3372 VDD.n1809 GND 0.006162f
C3373 VDD.n1810 GND 0.006162f
C3374 VDD.n1811 GND 0.006162f
C3375 VDD.n1812 GND 0.006162f
C3376 VDD.n1813 GND 0.006162f
C3377 VDD.n1814 GND 0.006162f
C3378 VDD.n1815 GND 0.006162f
C3379 VDD.n1816 GND 0.006162f
C3380 VDD.n1817 GND 0.006162f
C3381 VDD.n1818 GND 0.006162f
C3382 VDD.n1819 GND 0.006162f
C3383 VDD.n1820 GND 0.006162f
C3384 VDD.n1821 GND 0.006162f
C3385 VDD.n1822 GND 0.006162f
C3386 VDD.n1823 GND 0.006162f
C3387 VDD.n1824 GND 0.006162f
C3388 VDD.n1825 GND 0.006162f
C3389 VDD.n1826 GND 0.006162f
C3390 VDD.n1827 GND 0.006162f
C3391 VDD.n1828 GND 0.006162f
C3392 VDD.n1829 GND 0.006162f
C3393 VDD.n1830 GND 0.006162f
C3394 VDD.n1831 GND 0.004848f
C3395 VDD.n1832 GND 0.006162f
C3396 VDD.n1833 GND 0.006162f
C3397 VDD.n1834 GND 0.004395f
C3398 VDD.n1835 GND 0.006162f
C3399 VDD.n1836 GND 0.006162f
C3400 VDD.n1837 GND 0.014791f
C3401 VDD.n1838 GND 0.014027f
C3402 VDD.n1839 GND 0.014027f
C3403 VDD.n1840 GND 0.006162f
C3404 VDD.n1841 GND 0.006162f
C3405 VDD.n1842 GND 0.006162f
C3406 VDD.n1843 GND 0.006162f
C3407 VDD.n1844 GND 0.006162f
C3408 VDD.n1845 GND 0.006162f
C3409 VDD.n1846 GND 0.006162f
C3410 VDD.n1847 GND 0.006162f
C3411 VDD.n1848 GND 0.006162f
C3412 VDD.n1849 GND 0.006162f
C3413 VDD.n1850 GND 0.006162f
C3414 VDD.n1851 GND 0.006162f
C3415 VDD.n1852 GND 0.006162f
C3416 VDD.n1853 GND 0.006162f
C3417 VDD.n1854 GND 0.446608f
C3418 VDD.n1855 GND 0.006162f
C3419 VDD.n1856 GND 0.006162f
C3420 VDD.n1857 GND 0.006162f
C3421 VDD.n1858 GND 0.006162f
C3422 VDD.n1859 GND 0.006162f
C3423 VDD.n1860 GND 0.006162f
C3424 VDD.n1861 GND 0.006162f
C3425 VDD.n1862 GND 0.006162f
C3426 VDD.n1863 GND 0.006162f
C3427 VDD.n1864 GND 0.006162f
C3428 VDD.n1865 GND 0.006162f
C3429 VDD.n1866 GND 0.006162f
C3430 VDD.n1867 GND 0.006162f
C3431 VDD.n1868 GND 0.006162f
C3432 VDD.n1869 GND 0.006162f
C3433 VDD.n1870 GND 0.006162f
C3434 VDD.n1871 GND 0.006162f
C3435 VDD.n1872 GND 0.006162f
C3436 VDD.n1873 GND 0.006162f
C3437 VDD.n1874 GND 0.006162f
C3438 VDD.n1875 GND 0.006162f
C3439 VDD.n1876 GND 0.006162f
C3440 VDD.n1877 GND 0.006162f
C3441 VDD.n1878 GND 0.006162f
C3442 VDD.n1879 GND 0.006162f
C3443 VDD.n1880 GND 0.006162f
C3444 VDD.n1881 GND 0.006162f
C3445 VDD.n1882 GND 0.006162f
C3446 VDD.n1883 GND 0.006162f
C3447 VDD.n1884 GND 0.18638f
C3448 VDD.n1885 GND 0.006162f
C3449 VDD.n1886 GND 0.006162f
C3450 VDD.n1887 GND 0.006162f
C3451 VDD.n1888 GND 0.006162f
C3452 VDD.n1889 GND 0.006162f
C3453 VDD.n1890 GND 0.006162f
C3454 VDD.n1891 GND 0.006162f
C3455 VDD.n1892 GND 0.006162f
C3456 VDD.n1893 GND 0.006162f
C3457 VDD.n1894 GND 0.006162f
C3458 VDD.n1895 GND 0.006162f
C3459 VDD.n1896 GND 0.006162f
C3460 VDD.n1897 GND 0.006162f
C3461 VDD.n1898 GND 0.006162f
C3462 VDD.n1899 GND 0.006162f
C3463 VDD.n1900 GND 0.014027f
C3464 VDD.n1901 GND 0.014027f
C3465 VDD.n1902 GND 0.014791f
C3466 VDD.n1903 GND 0.014791f
C3467 VDD.n1904 GND 0.006162f
C3468 VDD.n1905 GND 0.006162f
C3469 VDD.n1906 GND 0.006162f
C3470 VDD.n1907 GND 0.004395f
C3471 VDD.n1908 GND 0.008807f
C3472 VDD.n1909 GND 0.004848f
C3473 VDD.n1910 GND 0.006162f
C3474 VDD.n1911 GND 0.006162f
C3475 VDD.n1912 GND 0.006162f
C3476 VDD.n1913 GND 0.006162f
C3477 VDD.n1914 GND 0.006162f
C3478 VDD.n1915 GND 0.006162f
C3479 VDD.n1916 GND 0.006162f
C3480 VDD.n1917 GND 0.006162f
C3481 VDD.n1918 GND 0.006162f
C3482 VDD.n1919 GND 0.006162f
C3483 VDD.n1920 GND 0.006162f
C3484 VDD.n1921 GND 0.006162f
C3485 VDD.n1922 GND 0.006162f
C3486 VDD.n1923 GND 0.006162f
C3487 VDD.n1924 GND 0.006162f
C3488 VDD.n1925 GND 0.006162f
C3489 VDD.n1926 GND 0.006162f
C3490 VDD.n1927 GND 0.006162f
C3491 VDD.n1928 GND 0.006162f
C3492 VDD.n1929 GND 0.006162f
C3493 VDD.n1930 GND 0.006162f
C3494 VDD.n1931 GND 0.006162f
C3495 VDD.n1932 GND 0.006162f
C3496 VDD.n1933 GND 0.006162f
C3497 VDD.n1934 GND 0.006162f
C3498 VDD.n1935 GND 0.006162f
C3499 VDD.n1936 GND 0.006162f
C3500 VDD.n1937 GND 0.006162f
C3501 VDD.n1938 GND 0.006162f
C3502 VDD.n1939 GND 0.006162f
C3503 VDD.n1940 GND 0.006162f
C3504 VDD.n1941 GND 0.006162f
C3505 VDD.n1942 GND 0.006162f
C3506 VDD.n1943 GND 0.006162f
C3507 VDD.n1944 GND 0.569689f
C3508 VDD.n1946 GND 0.014791f
C3509 VDD.n1947 GND 0.014791f
C3510 VDD.n1948 GND 0.014027f
C3511 VDD.n1949 GND 0.006162f
C3512 VDD.n1950 GND 0.006162f
C3513 VDD.n1951 GND 0.365726f
C3514 VDD.n1952 GND 0.006162f
C3515 VDD.n1953 GND 0.006162f
C3516 VDD.n1954 GND 0.006162f
C3517 VDD.n1955 GND 0.006162f
C3518 VDD.n1956 GND 0.006162f
C3519 VDD.n1957 GND 0.242645f
C3520 VDD.n1958 GND 0.006162f
C3521 VDD.n1959 GND 0.006162f
C3522 VDD.n1960 GND 0.006162f
C3523 VDD.n1961 GND 0.006162f
C3524 VDD.n1962 GND 0.006162f
C3525 VDD.n1963 GND 0.344627f
C3526 VDD.n1964 GND 0.006162f
C3527 VDD.n1965 GND 0.006162f
C3528 VDD.n1966 GND 0.006162f
C3529 VDD.n1967 GND 0.006162f
C3530 VDD.n1968 GND 0.006162f
C3531 VDD.n1969 GND 0.478257f
C3532 VDD.n1970 GND 0.006162f
C3533 VDD.n1971 GND 0.006162f
C3534 VDD.n1972 GND 0.006162f
C3535 VDD.n1973 GND 0.006162f
C3536 VDD.n1974 GND 0.006162f
C3537 VDD.n1975 GND 0.323527f
C3538 VDD.n1976 GND 0.006162f
C3539 VDD.n1977 GND 0.006162f
C3540 VDD.n1978 GND 0.006162f
C3541 VDD.n1979 GND 0.006162f
C3542 VDD.n1980 GND 0.006162f
C3543 VDD.n1981 GND 0.446608f
C3544 VDD.n1982 GND 0.006162f
C3545 VDD.n1983 GND 0.006162f
C3546 VDD.n1984 GND 0.006162f
C3547 VDD.n1985 GND 0.006162f
C3548 VDD.n1986 GND 0.006162f
C3549 VDD.n1987 GND 0.478257f
C3550 VDD.n1988 GND 0.006162f
C3551 VDD.n1989 GND 0.006162f
C3552 VDD.n1990 GND 0.006162f
C3553 VDD.n1991 GND 0.006162f
C3554 VDD.n1992 GND 0.006162f
C3555 VDD.n1993 GND 0.32001f
C3556 VDD.n1994 GND 0.006162f
C3557 VDD.n1995 GND 0.006162f
C3558 VDD.n1996 GND 0.006162f
C3559 VDD.n1997 GND 0.006162f
C3560 VDD.n1998 GND 0.006162f
C3561 VDD.n1999 GND 0.467707f
C3562 VDD.n2000 GND 0.006162f
C3563 VDD.n2001 GND 0.006162f
C3564 VDD.n2002 GND 0.006162f
C3565 VDD.n2003 GND 0.006162f
C3566 VDD.n2004 GND 0.006162f
C3567 VDD.n2005 GND 0.309461f
C3568 VDD.n2006 GND 0.006162f
C3569 VDD.n2007 GND 0.006162f
C3570 VDD.n2008 GND 0.006162f
C3571 VDD.n2009 GND 0.006162f
C3572 VDD.n2010 GND 0.006162f
C3573 VDD.n2011 GND 0.446608f
C3574 VDD.n2012 GND 0.006162f
C3575 VDD.n2013 GND 0.006162f
C3576 VDD.n2014 GND 0.006162f
C3577 VDD.n2015 GND 0.006162f
C3578 VDD.n2016 GND 0.006162f
C3579 VDD.n2017 GND 0.288361f
C3580 VDD.n2018 GND 0.006162f
C3581 VDD.n2019 GND 0.006162f
C3582 VDD.n2020 GND 0.006162f
C3583 VDD.n2021 GND 0.006162f
C3584 VDD.n2022 GND 0.006162f
C3585 VDD.n2023 GND 0.478257f
C3586 VDD.n2024 GND 0.006162f
C3587 VDD.n2025 GND 0.006162f
C3588 VDD.n2026 GND 0.006162f
C3589 VDD.t83 GND 0.131225f
C3590 VDD.t81 GND 0.198505f
C3591 VDD.t84 GND 0.131225f
C3592 VDD.n2027 GND 0.130384f
C3593 VDD.n2028 GND 0.028657f
C3594 VDD.n2029 GND 0.006162f
C3595 VDD.n2030 GND 0.006162f
C3596 VDD.n2032 GND 0.006162f
C3597 VDD.n2033 GND 0.006162f
C3598 VDD.n2036 GND 0.006162f
C3599 VDD.n2037 GND 0.006162f
C3600 VDD.n2038 GND 0.006162f
C3601 VDD.n2039 GND 0.006162f
C3602 VDD.n2041 GND 0.006162f
C3603 VDD.n2042 GND 0.006162f
C3604 VDD.n2043 GND 0.006162f
C3605 VDD.n2044 GND 0.006162f
C3606 VDD.n2045 GND 0.006162f
C3607 VDD.n2046 GND 0.006162f
C3608 VDD.n2048 GND 0.006162f
C3609 VDD.n2049 GND 0.006162f
C3610 VDD.n2050 GND 0.006162f
C3611 VDD.n2051 GND 0.006162f
C3612 VDD.n2052 GND 0.006842f
C3613 VDD.n2053 GND 0.014791f
C3614 VDD.n2054 GND 0.014027f
C3615 VDD.n2055 GND 0.00879f
C3616 VDD.n2056 GND 0.006162f
C3617 VDD.n2057 GND 0.006162f
C3618 VDD.n2058 GND 0.006162f
C3619 VDD.n2059 GND 0.006162f
C3620 VDD.n2060 GND 0.006162f
C3621 VDD.n2061 GND 0.006162f
C3622 VDD.n2062 GND 0.006162f
C3623 VDD.n2063 GND 0.267261f
C3624 VDD.n2064 GND 0.006162f
C3625 VDD.n2065 GND 0.006162f
C3626 VDD.n2066 GND 0.006162f
C3627 VDD.n2067 GND 0.006162f
C3628 VDD.n2068 GND 0.006162f
C3629 VDD.n2069 GND 0.242645f
C3630 VDD.n2070 GND 0.006162f
C3631 VDD.n2071 GND 0.006162f
C3632 VDD.n2072 GND 0.006162f
C3633 VDD.n2073 GND 0.006162f
C3634 VDD.n2074 GND 0.014756f
C3635 VDD.n2076 GND 0.014027f
C3636 VDD.n2077 GND 0.014791f
C3637 VDD.n2078 GND 0.014062f
C3638 VDD.n2079 GND 0.006162f
C3639 VDD.n2080 GND 0.004395f
C3640 VDD.n2081 GND 0.006162f
C3641 VDD.n2083 GND 0.006162f
C3642 VDD.n2084 GND 0.006162f
C3643 VDD.n2085 GND 0.006162f
C3644 VDD.n2086 GND 0.006162f
C3645 VDD.n2087 GND 0.006162f
C3646 VDD.n2088 GND 0.006162f
C3647 VDD.n2090 GND 0.006162f
C3648 VDD.n2091 GND 0.006162f
C3649 VDD.n2092 GND 0.006162f
C3650 VDD.n2093 GND 0.006162f
C3651 VDD.n2094 GND 0.006162f
C3652 VDD.n2095 GND 0.006162f
C3653 VDD.n2097 GND 0.006162f
C3654 VDD.n2098 GND 0.006162f
C3655 VDD.n2099 GND 0.006162f
C3656 VDD.n2101 GND 0.006162f
C3657 VDD.n2102 GND 0.006162f
C3658 VDD.n2103 GND 0.006162f
C3659 VDD.n2104 GND 0.006162f
C3660 VDD.n2105 GND 0.006162f
C3661 VDD.n2106 GND 0.006162f
C3662 VDD.n2108 GND 0.006162f
C3663 VDD.n2109 GND 0.006162f
C3664 VDD.n2110 GND 0.006162f
C3665 VDD.n2111 GND 0.006162f
C3666 VDD.n2112 GND 0.006162f
C3667 VDD.n2113 GND 0.006162f
C3668 VDD.n2115 GND 0.006162f
C3669 VDD.n2116 GND 0.014791f
C3670 VDD.n2117 GND 0.014791f
C3671 VDD.n2118 GND 0.014027f
C3672 VDD.n2119 GND 0.006162f
C3673 VDD.n2120 GND 0.006162f
C3674 VDD.n2121 GND 0.478257f
C3675 VDD.n2122 GND 0.006162f
C3676 VDD.n2123 GND 0.006162f
C3677 VDD.n2124 GND 0.014756f
C3678 VDD.n2125 GND 0.014062f
C3679 VDD.n2126 GND 0.014791f
C3680 VDD.n2128 GND 0.006162f
C3681 VDD.n2129 GND 0.006162f
C3682 VDD.n2130 GND 0.004395f
C3683 VDD.n2131 GND 0.008807f
C3684 VDD.n2132 GND 0.004848f
C3685 VDD.n2133 GND 0.006162f
C3686 VDD.n2134 GND 0.006162f
C3687 VDD.n2136 GND 0.006162f
C3688 VDD.n2137 GND 0.006162f
C3689 VDD.n2138 GND 0.006162f
C3690 VDD.n2139 GND 0.006162f
C3691 VDD.n2140 GND 0.006162f
C3692 VDD.n2141 GND 0.006162f
C3693 VDD.n2143 GND 0.006162f
C3694 VDD.n2144 GND 0.006162f
C3695 VDD.n2146 GND 0.006162f
C3696 VDD.n2147 GND 0.011006f
C3697 VDD.n2148 GND 0.009062f
C3698 VDD.n2149 GND 0.009062f
C3699 VDD.n2150 GND 0.007294f
C3700 VDD.n2151 GND 0.009062f
C3701 VDD.n2152 GND 0.009062f
C3702 VDD.n2153 GND 0.009062f
C3703 VDD.n2154 GND 0.009062f
C3704 VDD.n2155 GND 0.009062f
C3705 VDD.n2156 GND 0.009062f
C3706 VDD.n2157 GND 0.02042f
C3707 VDD.n2158 GND 0.003465f
C3708 VDD.t55 GND 0.18563f
C3709 VDD.t56 GND 0.194533f
C3710 VDD.t54 GND 0.271204f
C3711 VDD.n2159 GND 0.091924f
C3712 VDD.n2160 GND 0.052705f
C3713 VDD.n2161 GND 0.011269f
C3714 VDD.n2162 GND 0.009062f
C3715 VDD.n2163 GND 0.003829f
C3716 VDD.n2164 GND 0.007294f
C3717 VDD.n2165 GND 0.009062f
C3718 VDD.n2166 GND 0.009062f
C3719 VDD.n2167 GND 0.007294f
C3720 VDD.n2168 GND 0.007294f
C3721 VDD.n2169 GND 0.009062f
C3722 VDD.n2170 GND 0.009062f
C3723 VDD.n2171 GND 0.007294f
C3724 VDD.n2172 GND 0.009062f
C3725 VDD.n2173 GND 0.007294f
C3726 VDD.n2174 GND 0.007294f
C3727 VDD.n2176 GND 0.442633f
C3728 VDD.n2178 GND 0.007294f
C3729 VDD.n2179 GND 0.009062f
C3730 VDD.n2180 GND 0.009062f
C3731 VDD.n2181 GND 0.007294f
C3732 VDD.n2182 GND 0.007294f
C3733 VDD.n2183 GND 0.009062f
C3734 VDD.n2184 GND 0.009062f
C3735 VDD.n2185 GND 0.007294f
C3736 VDD.n2186 GND 0.007294f
C3737 VDD.n2187 GND 0.009062f
C3738 VDD.n2188 GND 0.009062f
C3739 VDD.n2189 GND 0.007294f
C3740 VDD.n2190 GND 0.007294f
C3741 VDD.n2191 GND 0.009062f
C3742 VDD.n2192 GND 0.009062f
C3743 VDD.n2193 GND 0.007294f
C3744 VDD.n2194 GND 0.009062f
C3745 VDD.n2195 GND 0.009062f
C3746 VDD.n2196 GND 0.007294f
C3747 VDD.n2197 GND 0.009062f
C3748 VDD.n2198 GND 0.009062f
C3749 VDD.n2199 GND 0.009062f
C3750 VDD.n2200 GND 0.014916f
C3751 VDD.n2201 GND 0.009062f
C3752 VDD.n2202 GND 0.009062f
C3753 VDD.n2203 GND 0.00496f
C3754 VDD.n2204 GND 0.007294f
C3755 VDD.n2205 GND 0.009062f
C3756 VDD.n2206 GND 0.009062f
C3757 VDD.n2207 GND 0.007294f
C3758 VDD.n2208 GND 0.007294f
C3759 VDD.n2209 GND 0.009062f
C3760 VDD.n2210 GND 0.009062f
C3761 VDD.n2211 GND 0.007294f
C3762 VDD.n2212 GND 0.007294f
C3763 VDD.n2213 GND 0.009062f
C3764 VDD.n2214 GND 0.009062f
C3765 VDD.n2215 GND 0.007294f
C3766 VDD.n2216 GND 0.007294f
C3767 VDD.n2217 GND 0.009062f
C3768 VDD.n2218 GND 0.009062f
C3769 VDD.n2219 GND 0.007294f
C3770 VDD.n2220 GND 0.007294f
C3771 VDD.n2221 GND 0.009062f
C3772 VDD.n2222 GND 0.009062f
C3773 VDD.n2223 GND 0.007294f
C3774 VDD.n2224 GND 0.007294f
C3775 VDD.n2225 GND 0.009062f
C3776 VDD.n2226 GND 0.009062f
C3777 VDD.n2227 GND 0.007294f
C3778 VDD.n2228 GND 0.007294f
C3779 VDD.n2229 GND 0.009062f
C3780 VDD.n2230 GND 0.009062f
C3781 VDD.n2231 GND 0.007294f
C3782 VDD.n2232 GND 0.007294f
C3783 VDD.n2233 GND 0.009062f
C3784 VDD.n2234 GND 0.009062f
C3785 VDD.n2235 GND 0.007294f
C3786 VDD.n2236 GND 0.009062f
C3787 VDD.n2237 GND 0.009062f
C3788 VDD.n2238 GND 0.007294f
C3789 VDD.n2239 GND 0.009062f
C3790 VDD.n2240 GND 0.009062f
C3791 VDD.n2241 GND 0.009062f
C3792 VDD.t75 GND 0.18563f
C3793 VDD.t76 GND 0.194533f
C3794 VDD.t74 GND 0.271204f
C3795 VDD.n2242 GND 0.091924f
C3796 VDD.n2243 GND 0.052705f
C3797 VDD.n2244 GND 0.014916f
C3798 VDD.n2245 GND 0.009062f
C3799 VDD.n2246 GND 0.009062f
C3800 VDD.n2247 GND 0.00609f
C3801 VDD.n2248 GND 0.007294f
C3802 VDD.n2249 GND 0.009062f
C3803 VDD.n2250 GND 0.009062f
C3804 VDD.n2251 GND 0.007294f
C3805 VDD.n2252 GND 0.007294f
C3806 VDD.n2253 GND 0.009062f
C3807 VDD.n2254 GND 0.009062f
C3808 VDD.n2255 GND 0.007294f
C3809 VDD.n2256 GND 0.009062f
C3810 VDD.n2257 GND 0.007294f
C3811 VDD.n2258 GND 0.007294f
C3812 VDD.n2260 GND 0.442633f
C3813 VDD.n2262 GND 0.007294f
C3814 VDD.n2263 GND 0.009062f
C3815 VDD.n2264 GND 0.009062f
C3816 VDD.n2265 GND 0.007294f
C3817 VDD.n2266 GND 0.007294f
C3818 VDD.n2267 GND 0.009062f
C3819 VDD.n2268 GND 0.009062f
C3820 VDD.n2269 GND 0.007294f
C3821 VDD.n2270 GND 0.007294f
C3822 VDD.n2271 GND 0.007294f
C3823 VDD.n2272 GND 0.009062f
C3824 VDD.n2273 GND 3.9843f
C3825 VDD.n2275 GND 0.02042f
C3826 VDD.n2276 GND 0.006054f
C3827 VDD.n2277 GND 0.02042f
C3828 VDD.n2278 GND 0.02036f
C3829 VDD.n2279 GND 0.009062f
C3830 VDD.n2280 GND 0.007294f
C3831 VDD.n2281 GND 0.009062f
C3832 VDD.n2282 GND 0.594305f
C3833 VDD.n2283 GND 0.009062f
C3834 VDD.n2284 GND 0.007294f
C3835 VDD.n2285 GND 0.009062f
C3836 VDD.n2286 GND 0.009062f
C3837 VDD.n2287 GND 0.009062f
C3838 VDD.n2288 GND 0.007294f
C3839 VDD.n2289 GND 0.009062f
C3840 VDD.n2290 GND 0.703319f
C3841 VDD.n2291 GND 0.009062f
C3842 VDD.n2292 GND 0.007294f
C3843 VDD.n2293 GND 0.009062f
C3844 VDD.n2294 GND 0.009062f
C3845 VDD.n2295 GND 0.009062f
C3846 VDD.n2296 GND 0.007294f
C3847 VDD.n2297 GND 0.009062f
C3848 VDD.n2298 GND 0.703319f
C3849 VDD.n2299 GND 0.009062f
C3850 VDD.n2300 GND 0.007294f
C3851 VDD.n2301 GND 0.009062f
C3852 VDD.n2302 GND 0.009062f
C3853 VDD.n2303 GND 0.009062f
C3854 VDD.n2304 GND 0.007294f
C3855 VDD.n2305 GND 0.009062f
C3856 VDD.n2306 GND 0.51694f
C3857 VDD.n2307 GND 0.009062f
C3858 VDD.n2308 GND 0.007294f
C3859 VDD.n2309 GND 0.009062f
C3860 VDD.n2310 GND 0.009062f
C3861 VDD.n2311 GND 0.009062f
C3862 VDD.n2312 GND 0.007294f
C3863 VDD.n2313 GND 0.009062f
C3864 VDD.n2314 GND 0.418475f
C3865 VDD.n2315 GND 0.009062f
C3866 VDD.n2316 GND 0.007294f
C3867 VDD.n2317 GND 0.009062f
C3868 VDD.n2318 GND 0.009062f
C3869 VDD.n2319 GND 0.009062f
C3870 VDD.n2320 GND 0.007294f
C3871 VDD.n2321 GND 0.009062f
C3872 VDD.t116 GND 0.35166f
C3873 VDD.n2322 GND 0.65057f
C3874 VDD.n2323 GND 0.009062f
C3875 VDD.n2324 GND 0.007294f
C3876 VDD.n2325 GND 0.009062f
C3877 VDD.n2326 GND 0.009062f
C3878 VDD.n2327 GND 0.009062f
C3879 VDD.n2328 GND 0.007294f
C3880 VDD.n2329 GND 0.009062f
C3881 VDD.n2330 GND 0.703319f
C3882 VDD.n2331 GND 0.009062f
C3883 VDD.n2332 GND 0.007294f
C3884 VDD.n2333 GND 0.009062f
C3885 VDD.n2334 GND 0.009062f
C3886 VDD.n2335 GND 0.009062f
C3887 VDD.n2336 GND 0.007294f
C3888 VDD.n2337 GND 0.009062f
C3889 VDD.n2338 GND 0.523973f
C3890 VDD.n2339 GND 0.009062f
C3891 VDD.n2340 GND 0.007294f
C3892 VDD.n2341 GND 0.009062f
C3893 VDD.n2342 GND 0.009062f
C3894 VDD.n2343 GND 0.009062f
C3895 VDD.n2344 GND 0.007294f
C3896 VDD.n2345 GND 0.009062f
C3897 VDD.n2346 GND 0.411442f
C3898 VDD.n2347 GND 0.009062f
C3899 VDD.n2348 GND 0.007294f
C3900 VDD.n2349 GND 0.009062f
C3901 VDD.n2350 GND 0.009062f
C3902 VDD.n2351 GND 0.009062f
C3903 VDD.n2352 GND 0.007294f
C3904 VDD.n2353 GND 0.007294f
C3905 VDD.n2354 GND 0.007294f
C3906 VDD.n2355 GND 0.009062f
C3907 VDD.n2356 GND 0.009062f
C3908 VDD.n2357 GND 0.009062f
C3909 VDD.n2358 GND 0.007294f
C3910 VDD.n2359 GND 0.007294f
C3911 VDD.n2360 GND 0.007294f
C3912 VDD.n2361 GND 0.009062f
C3913 VDD.n2362 GND 0.009062f
C3914 VDD.n2363 GND 0.009062f
C3915 VDD.n2364 GND 0.007294f
C3916 VDD.n2365 GND 0.007294f
C3917 VDD.n2366 GND 0.007294f
C3918 VDD.n2367 GND 0.009062f
C3919 VDD.n2368 GND 0.009062f
C3920 VDD.n2369 GND 0.009062f
C3921 VDD.n2370 GND 0.007294f
C3922 VDD.n2371 GND 0.007294f
C3923 VDD.n2372 GND 0.007294f
C3924 VDD.n2373 GND 0.009062f
C3925 VDD.n2374 GND 0.009062f
C3926 VDD.n2375 GND 0.009062f
C3927 VDD.n2376 GND 0.007294f
C3928 VDD.n2377 GND 0.007294f
C3929 VDD.n2378 GND 0.006054f
C3930 VDD.n2379 GND 0.02036f
C3931 VDD.n2380 GND 0.02042f
C3932 VDD.n2381 GND 0.003465f
C3933 VDD.n2382 GND 0.02042f
C3934 VDD.n2384 GND 0.009062f
C3935 VDD.n2385 GND 0.009062f
C3936 VDD.n2386 GND 0.007294f
C3937 VDD.n2387 GND 0.007294f
C3938 VDD.n2388 GND 0.007294f
C3939 VDD.n2389 GND 0.009062f
C3940 VDD.n2391 GND 0.009062f
C3941 VDD.n2392 GND 0.009062f
C3942 VDD.n2393 GND 0.007294f
C3943 VDD.n2394 GND 0.007294f
C3944 VDD.n2395 GND 0.007294f
C3945 VDD.n2396 GND 0.009062f
C3946 VDD.n2398 GND 0.009062f
C3947 VDD.n2399 GND 0.009062f
C3948 VDD.n2400 GND 0.007294f
C3949 VDD.n2401 GND 0.007294f
C3950 VDD.n2402 GND 0.007294f
C3951 VDD.n2403 GND 0.009062f
C3952 VDD.n2405 GND 0.009062f
C3953 VDD.n2406 GND 0.009062f
C3954 VDD.n2407 GND 0.007294f
C3955 VDD.n2408 GND 0.007294f
C3956 VDD.n2409 GND 0.007294f
C3957 VDD.n2410 GND 0.009062f
C3958 VDD.n2412 GND 0.009062f
C3959 VDD.n2413 GND 0.009062f
C3960 VDD.n2414 GND 0.007294f
C3961 VDD.n2415 GND 0.009062f
C3962 VDD.n2416 GND 0.009062f
C3963 VDD.n2417 GND 0.009062f
C3964 VDD.n2418 GND 0.014916f
C3965 VDD.n2419 GND 0.009062f
C3966 VDD.n2421 GND 0.009062f
C3967 VDD.n2422 GND 0.009062f
C3968 VDD.n2423 GND 0.007294f
C3969 VDD.n2424 GND 0.007294f
C3970 VDD.n2425 GND 0.007294f
C3971 VDD.n2426 GND 0.009062f
C3972 VDD.n2428 GND 0.009062f
C3973 VDD.n2429 GND 0.009062f
C3974 VDD.n2430 GND 0.007294f
C3975 VDD.n2431 GND 0.007294f
C3976 VDD.n2432 GND 0.007294f
C3977 VDD.n2433 GND 0.009062f
C3978 VDD.n2435 GND 0.009062f
C3979 VDD.n2436 GND 0.009062f
C3980 VDD.n2437 GND 0.007294f
C3981 VDD.n2438 GND 0.007294f
C3982 VDD.n2439 GND 0.007294f
C3983 VDD.n2440 GND 0.009062f
C3984 VDD.n2442 GND 0.009062f
C3985 VDD.n2443 GND 0.009062f
C3986 VDD.n2444 GND 0.007294f
C3987 VDD.n2445 GND 0.007294f
C3988 VDD.n2446 GND 0.007294f
C3989 VDD.n2447 GND 0.009062f
C3990 VDD.n2449 GND 0.009062f
C3991 VDD.n2450 GND 0.009062f
C3992 VDD.n2451 GND 0.007294f
C3993 VDD.n2452 GND 0.009062f
C3994 VDD.n2453 GND 0.009062f
C3995 VDD.n2454 GND 0.009062f
C3996 VDD.n2455 GND 0.014916f
C3997 VDD.n2456 GND 0.009062f
C3998 VDD.n2458 GND 0.009062f
C3999 VDD.n2459 GND 0.009062f
C4000 VDD.n2460 GND 0.007294f
C4001 VDD.n2461 GND 0.007294f
C4002 VDD.n2462 GND 0.007294f
C4003 VDD.n2463 GND 0.009062f
C4004 VDD.n2465 GND 0.009062f
C4005 VDD.n2466 GND 0.009062f
C4006 VDD.n2467 GND 0.007294f
C4007 VDD.n2468 GND 0.007294f
C4008 VDD.n2469 GND 0.007294f
C4009 VDD.n2470 GND 0.009062f
C4010 VDD.n2472 GND 0.009062f
C4011 VDD.n2473 GND 0.009062f
C4012 VDD.n2474 GND 0.007294f
C4013 VDD.n2475 GND 0.007294f
C4014 VDD.n2476 GND 0.007294f
C4015 VDD.n2477 GND 0.009062f
C4016 VDD.n2479 GND 0.009062f
C4017 VDD.n2480 GND 0.009062f
C4018 VDD.n2482 GND 0.009062f
C4019 VDD.n2483 GND 0.007294f
C4020 VDD.n2484 GND 0.007294f
C4021 VDD.n2485 GND 0.006054f
C4022 VDD.n2486 GND 0.02042f
C4023 VDD.n2487 GND 0.02036f
C4024 VDD.n2488 GND 0.006054f
C4025 VDD.n2489 GND 0.02036f
C4026 VDD.n2490 GND 0.903766f
C4027 VDD.n2491 GND 0.594305f
C4028 VDD.t51 GND 0.35166f
C4029 VDD.n2492 GND 0.460674f
C4030 VDD.n2493 GND 0.009062f
C4031 VDD.n2494 GND 0.007294f
C4032 VDD.n2495 GND 0.007294f
C4033 VDD.n2496 GND 0.007294f
C4034 VDD.n2497 GND 0.009062f
C4035 VDD.n2498 GND 0.703319f
C4036 VDD.n2499 GND 0.703319f
C4037 VDD.n2500 GND 0.538039f
C4038 VDD.n2501 GND 0.009062f
C4039 VDD.n2502 GND 0.007294f
C4040 VDD.n2503 GND 0.007294f
C4041 VDD.n2504 GND 0.007294f
C4042 VDD.n2505 GND 0.009062f
C4043 VDD.n2506 GND 0.703319f
C4044 VDD.n2507 GND 0.418475f
C4045 VDD.t152 GND 0.35166f
C4046 VDD.n2508 GND 0.636504f
C4047 VDD.n2509 GND 0.009062f
C4048 VDD.n2510 GND 0.007294f
C4049 VDD.n2511 GND 0.007294f
C4050 VDD.n2512 GND 0.007294f
C4051 VDD.n2513 GND 0.009062f
C4052 VDD.n2514 GND 0.404409f
C4053 VDD.n2515 GND 0.703319f
C4054 VDD.n2516 GND 0.531006f
C4055 VDD.n2517 GND 0.009062f
C4056 VDD.n2518 GND 0.007294f
C4057 VDD.n2519 GND 0.007294f
C4058 VDD.n2520 GND 0.007294f
C4059 VDD.n2521 GND 0.009062f
C4060 VDD.n2522 GND 0.703319f
C4061 VDD.n2523 GND 0.411442f
C4062 VDD.t131 GND 0.35166f
C4063 VDD.n2524 GND 0.643537f
C4064 VDD.n2525 GND 0.009062f
C4065 VDD.n2526 GND 0.007294f
C4066 VDD.n2527 GND 0.006965f
C4067 VDD.n2528 GND 0.19573f
C4068 VDD.n2529 GND 1.70151f
C4069 a_n7097_7899.n0 GND 0.653304f
C4070 a_n7097_7899.n1 GND 0.49431f
C4071 a_n7097_7899.n2 GND 0.653304f
C4072 a_n7097_7899.n3 GND 0.49431f
C4073 a_n7097_7899.n4 GND 0.871171f
C4074 a_n7097_7899.n5 GND 0.038759f
C4075 a_n7097_7899.n6 GND 0.038759f
C4076 a_n7097_7899.n7 GND 0.085574f
C4077 a_n7097_7899.n8 GND 0.050196f
C4078 a_n7097_7899.n9 GND 0.379714f
C4079 a_n7097_7899.n10 GND 0.379714f
C4080 a_n7097_7899.n11 GND 0.379714f
C4081 a_n7097_7899.n12 GND 0.040918f
C4082 a_n7097_7899.n13 GND 0.038759f
C4083 a_n7097_7899.n14 GND 0.04091f
C4084 a_n7097_7899.n15 GND 0.040911f
C4085 a_n7097_7899.n16 GND 0.040918f
C4086 a_n7097_7899.n17 GND 0.038759f
C4087 a_n7097_7899.n18 GND 0.04091f
C4088 a_n7097_7899.n19 GND 0.040911f
C4089 a_n7097_7899.n20 GND 0.040918f
C4090 a_n7097_7899.n21 GND 0.038759f
C4091 a_n7097_7899.n22 GND 0.04091f
C4092 a_n7097_7899.n23 GND 0.385101f
C4093 a_n7097_7899.n24 GND 0.04354f
C4094 a_n7097_7899.n25 GND 0.385101f
C4095 a_n7097_7899.n26 GND 0.04354f
C4096 a_n7097_7899.n27 GND 0.385101f
C4097 a_n7097_7899.n28 GND 0.04354f
C4098 a_n7097_7899.n29 GND 0.050196f
C4099 a_n7097_7899.n30 GND 0.050196f
C4100 a_n7097_7899.n31 GND 0.050196f
C4101 a_n7097_7899.n32 GND 0.043015f
C4102 a_n7097_7899.n33 GND 0.225434f
C4103 a_n7097_7899.n34 GND 0.085574f
C4104 a_n7097_7899.n35 GND 0.041787f
C4105 a_n7097_7899.n36 GND 0.225434f
C4106 a_n7097_7899.n37 GND 0.041787f
C4107 a_n7097_7899.n38 GND 0.085574f
C4108 a_n7097_7899.n39 GND 0.085574f
C4109 a_n7097_7899.n40 GND 0.043015f
C4110 a_n7097_7899.n41 GND 0.085574f
C4111 a_n7097_7899.n42 GND 0.050196f
C4112 a_n7097_7899.n43 GND 0.068975f
C4113 a_n7097_7899.n44 GND 0.042045f
C4114 a_n7097_7899.n45 GND 0.085574f
C4115 a_n7097_7899.n46 GND 0.085574f
C4116 a_n7097_7899.n47 GND 0.085574f
C4117 a_n7097_7899.n48 GND 0.085574f
C4118 a_n7097_7899.n49 GND 0.04974f
C4119 a_n7097_7899.n50 GND 0.06894f
C4120 a_n7097_7899.n51 GND 0.042331f
C4121 a_n7097_7899.n52 GND 0.085574f
C4122 a_n7097_7899.n53 GND 0.099881f
C4123 a_n7097_7899.n54 GND 0.225434f
C4124 a_n7097_7899.n55 GND 0.041787f
C4125 a_n7097_7899.n56 GND 0.085574f
C4126 a_n7097_7899.n57 GND 0.085574f
C4127 a_n7097_7899.n58 GND 0.043015f
C4128 a_n7097_7899.n59 GND 0.085574f
C4129 a_n7097_7899.n60 GND 0.050196f
C4130 a_n7097_7899.n61 GND 0.068975f
C4131 a_n7097_7899.n62 GND 0.042045f
C4132 a_n7097_7899.n63 GND 0.085574f
C4133 a_n7097_7899.n64 GND 0.085574f
C4134 a_n7097_7899.n65 GND 0.085574f
C4135 a_n7097_7899.n66 GND 0.085574f
C4136 a_n7097_7899.n67 GND 0.04974f
C4137 a_n7097_7899.n68 GND 0.06894f
C4138 a_n7097_7899.n69 GND 0.042331f
C4139 a_n7097_7899.n70 GND 0.085574f
C4140 a_n7097_7899.n71 GND 0.099881f
C4141 a_n7097_7899.n72 GND 0.225434f
C4142 a_n7097_7899.n73 GND 0.041787f
C4143 a_n7097_7899.n74 GND 0.085574f
C4144 a_n7097_7899.n75 GND 0.085574f
C4145 a_n7097_7899.n76 GND 0.043015f
C4146 a_n7097_7899.n77 GND 0.085574f
C4147 a_n7097_7899.n78 GND 0.050196f
C4148 a_n7097_7899.n79 GND 0.068975f
C4149 a_n7097_7899.n80 GND 0.042045f
C4150 a_n7097_7899.n81 GND 0.085574f
C4151 a_n7097_7899.n82 GND 0.085574f
C4152 a_n7097_7899.n83 GND 0.085574f
C4153 a_n7097_7899.n84 GND 0.085574f
C4154 a_n7097_7899.n85 GND 0.04974f
C4155 a_n7097_7899.n86 GND 0.06894f
C4156 a_n7097_7899.n87 GND 0.042331f
C4157 a_n7097_7899.n88 GND 0.085574f
C4158 a_n7097_7899.n89 GND 0.099881f
C4159 a_n7097_7899.t15 GND 0.07914f
C4160 a_n7097_7899.t4 GND 0.06595f
C4161 a_n7097_7899.t13 GND 0.06595f
C4162 a_n7097_7899.n90 GND 0.456317f
C4163 a_n7097_7899.t14 GND 0.06595f
C4164 a_n7097_7899.t0 GND 0.06595f
C4165 a_n7097_7899.n91 GND 0.453923f
C4166 a_n7097_7899.n92 GND 2.57517f
C4167 a_n7097_7899.t2 GND 0.06595f
C4168 a_n7097_7899.t12 GND 0.06595f
C4169 a_n7097_7899.n93 GND 0.456319f
C4170 a_n7097_7899.t5 GND 0.06595f
C4171 a_n7097_7899.t11 GND 0.06595f
C4172 a_n7097_7899.n94 GND 0.453923f
C4173 a_n7097_7899.n95 GND 1.93472f
C4174 a_n7097_7899.n96 GND 4.27688f
C4175 a_n7097_7899.t20 GND 0.799395f
C4176 a_n7097_7899.t56 GND 0.799395f
C4177 a_n7097_7899.t66 GND 0.799395f
C4178 a_n7097_7899.t46 GND 0.799395f
C4179 a_n7097_7899.t72 GND 0.799395f
C4180 a_n7097_7899.n97 GND 0.385425f
C4181 a_n7097_7899.t54 GND 0.799395f
C4182 a_n7097_7899.n98 GND 0.318958f
C4183 a_n7097_7899.t30 GND 0.799395f
C4184 a_n7097_7899.n99 GND 0.396682f
C4185 a_n7097_7899.t65 GND 0.890701f
C4186 a_n7097_7899.n100 GND 0.380544f
C4187 a_n7097_7899.n101 GND 0.068995f
C4188 a_n7097_7899.n102 GND 0.067784f
C4189 a_n7097_7899.n103 GND 0.394056f
C4190 a_n7097_7899.n104 GND 0.318958f
C4191 a_n7097_7899.n105 GND 0.067537f
C4192 a_n7097_7899.t32 GND 0.799395f
C4193 a_n7097_7899.n106 GND 0.394308f
C4194 a_n7097_7899.n107 GND 0.318958f
C4195 a_n7097_7899.n108 GND 0.058175f
C4196 a_n7097_7899.t48 GND 0.864545f
C4197 a_n7097_7899.n109 GND 0.384879f
C4198 a_n7097_7899.n110 GND 0.257846f
C4199 a_n7097_7899.t51 GND 0.799395f
C4200 a_n7097_7899.t23 GND 0.799395f
C4201 a_n7097_7899.t36 GND 0.799395f
C4202 a_n7097_7899.t75 GND 0.799395f
C4203 a_n7097_7899.t44 GND 0.799395f
C4204 a_n7097_7899.n111 GND 0.385425f
C4205 a_n7097_7899.t21 GND 0.799395f
C4206 a_n7097_7899.n112 GND 0.318958f
C4207 a_n7097_7899.t60 GND 0.799395f
C4208 a_n7097_7899.n113 GND 0.396682f
C4209 a_n7097_7899.t34 GND 0.890701f
C4210 a_n7097_7899.n114 GND 0.380544f
C4211 a_n7097_7899.n115 GND 0.068995f
C4212 a_n7097_7899.n116 GND 0.067784f
C4213 a_n7097_7899.n117 GND 0.394056f
C4214 a_n7097_7899.n118 GND 0.318958f
C4215 a_n7097_7899.n119 GND 0.067537f
C4216 a_n7097_7899.t61 GND 0.799395f
C4217 a_n7097_7899.n120 GND 0.394308f
C4218 a_n7097_7899.n121 GND 0.318958f
C4219 a_n7097_7899.n122 GND 0.058175f
C4220 a_n7097_7899.t16 GND 0.864545f
C4221 a_n7097_7899.n123 GND 0.384879f
C4222 a_n7097_7899.n124 GND 0.137707f
C4223 a_n7097_7899.n125 GND 0.69844f
C4224 a_n7097_7899.t52 GND 0.799395f
C4225 a_n7097_7899.t24 GND 0.799395f
C4226 a_n7097_7899.t47 GND 0.799395f
C4227 a_n7097_7899.t58 GND 0.799395f
C4228 a_n7097_7899.t28 GND 0.799395f
C4229 a_n7097_7899.n126 GND 0.385425f
C4230 a_n7097_7899.t43 GND 0.799395f
C4231 a_n7097_7899.n127 GND 0.318958f
C4232 a_n7097_7899.t53 GND 0.799395f
C4233 a_n7097_7899.n128 GND 0.396682f
C4234 a_n7097_7899.t62 GND 0.890701f
C4235 a_n7097_7899.n129 GND 0.380544f
C4236 a_n7097_7899.n130 GND 0.068995f
C4237 a_n7097_7899.n131 GND 0.067784f
C4238 a_n7097_7899.n132 GND 0.394056f
C4239 a_n7097_7899.n133 GND 0.318958f
C4240 a_n7097_7899.n134 GND 0.067537f
C4241 a_n7097_7899.t35 GND 0.799395f
C4242 a_n7097_7899.n135 GND 0.394308f
C4243 a_n7097_7899.n136 GND 0.318958f
C4244 a_n7097_7899.n137 GND 0.058175f
C4245 a_n7097_7899.t42 GND 0.864545f
C4246 a_n7097_7899.n138 GND 0.384879f
C4247 a_n7097_7899.n139 GND 0.137707f
C4248 a_n7097_7899.n140 GND 1.13839f
C4249 a_n7097_7899.t64 GND 0.890619f
C4250 a_n7097_7899.t38 GND 0.799395f
C4251 a_n7097_7899.t71 GND 0.799395f
C4252 a_n7097_7899.t50 GND 0.799395f
C4253 a_n7097_7899.n141 GND 0.410546f
C4254 a_n7097_7899.t22 GND 0.799395f
C4255 a_n7097_7899.t57 GND 0.799395f
C4256 a_n7097_7899.t29 GND 0.799395f
C4257 a_n7097_7899.n142 GND 0.385425f
C4258 a_n7097_7899.t68 GND 0.799395f
C4259 a_n7097_7899.n143 GND 0.318958f
C4260 a_n7097_7899.t49 GND 0.799395f
C4261 a_n7097_7899.n144 GND 0.396682f
C4262 a_n7097_7899.t74 GND 0.890701f
C4263 a_n7097_7899.n145 GND 0.380543f
C4264 a_n7097_7899.n146 GND 0.068995f
C4265 a_n7097_7899.n147 GND 0.067784f
C4266 a_n7097_7899.n148 GND 0.408992f
C4267 a_n7097_7899.n149 GND 0.408992f
C4268 a_n7097_7899.n150 GND 0.420482f
C4269 a_n7097_7899.n151 GND 0.411962f
C4270 a_n7097_7899.t33 GND 0.890619f
C4271 a_n7097_7899.t67 GND 0.799395f
C4272 a_n7097_7899.t41 GND 0.799395f
C4273 a_n7097_7899.t18 GND 0.799395f
C4274 a_n7097_7899.n152 GND 0.384531f
C4275 a_n7097_7899.t55 GND 0.799395f
C4276 a_n7097_7899.t25 GND 0.799395f
C4277 a_n7097_7899.t59 GND 0.799395f
C4278 a_n7097_7899.n153 GND 0.410545f
C4279 a_n7097_7899.t40 GND 0.799395f
C4280 a_n7097_7899.n154 GND 0.420482f
C4281 a_n7097_7899.t17 GND 0.799395f
C4282 a_n7097_7899.n155 GND 0.41195f
C4283 a_n7097_7899.t45 GND 0.890701f
C4284 a_n7097_7899.n156 GND 0.380543f
C4285 a_n7097_7899.n157 GND 0.408992f
C4286 a_n7097_7899.n158 GND 0.374125f
C4287 a_n7097_7899.n159 GND 0.058742f
C4288 a_n7097_7899.n160 GND 0.052335f
C4289 a_n7097_7899.n161 GND 0.420482f
C4290 a_n7097_7899.n162 GND 0.411962f
C4291 a_n7097_7899.n163 GND 0.69844f
C4292 a_n7097_7899.t27 GND 0.890619f
C4293 a_n7097_7899.t37 GND 0.799395f
C4294 a_n7097_7899.t70 GND 0.799395f
C4295 a_n7097_7899.t19 GND 0.799395f
C4296 a_n7097_7899.n164 GND 0.384531f
C4297 a_n7097_7899.t31 GND 0.799395f
C4298 a_n7097_7899.t63 GND 0.799395f
C4299 a_n7097_7899.t73 GND 0.799395f
C4300 a_n7097_7899.n165 GND 0.410545f
C4301 a_n7097_7899.t26 GND 0.799395f
C4302 a_n7097_7899.n166 GND 0.420482f
C4303 a_n7097_7899.t39 GND 0.799395f
C4304 a_n7097_7899.n167 GND 0.41195f
C4305 a_n7097_7899.t69 GND 0.890701f
C4306 a_n7097_7899.n168 GND 0.380543f
C4307 a_n7097_7899.n169 GND 0.408992f
C4308 a_n7097_7899.n170 GND 0.374125f
C4309 a_n7097_7899.n171 GND 0.058742f
C4310 a_n7097_7899.n172 GND 0.052335f
C4311 a_n7097_7899.n173 GND 0.420482f
C4312 a_n7097_7899.n174 GND 0.411962f
C4313 a_n7097_7899.n175 GND 0.946967f
C4314 a_n7097_7899.n176 GND 9.981219f
C4315 a_n7097_7899.n177 GND 3.8081f
C4316 a_n7097_7899.t9 GND 0.07914f
C4317 a_n7097_7899.t3 GND 0.07914f
C4318 a_n7097_7899.n178 GND 0.692272f
C4319 a_n7097_7899.n179 GND 0.750678f
C4320 a_n7097_7899.t7 GND 0.07914f
C4321 a_n7097_7899.t6 GND 0.07914f
C4322 a_n7097_7899.n180 GND 0.691165f
C4323 a_n7097_7899.n181 GND 1.92166f
C4324 a_n7097_7899.t8 GND 0.07914f
C4325 a_n7097_7899.t10 GND 0.07914f
C4326 a_n7097_7899.n182 GND 0.692269f
C4327 a_n7097_7899.n183 GND 2.04622f
C4328 a_n7097_7899.n184 GND 0.692269f
C4329 a_n7097_7899.t1 GND 0.07914f
.ends

