* NGSPICE file created from diff_pair_sample_0450.ext - technology: sky130A

.subckt diff_pair_sample_0450 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=0 ps=0 w=9.87 l=1.24
X1 B.t8 B.t6 B.t7 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=0 ps=0 w=9.87 l=1.24
X2 VTAIL.t15 VP.t0 VDD1.t5 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=1.62855 ps=10.2 w=9.87 l=1.24
X3 VTAIL.t7 VN.t0 VDD2.t7 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=1.62855 ps=10.2 w=9.87 l=1.24
X4 VTAIL.t1 VN.t1 VDD2.t6 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=1.62855 ps=10.2 w=9.87 l=1.24
X5 VTAIL.t14 VP.t1 VDD1.t6 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X6 VDD2.t5 VN.t2 VTAIL.t2 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=3.8493 ps=20.52 w=9.87 l=1.24
X7 B.t5 B.t3 B.t4 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=0 ps=0 w=9.87 l=1.24
X8 VDD1.t0 VP.t2 VTAIL.t13 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=3.8493 ps=20.52 w=9.87 l=1.24
X9 VDD2.t4 VN.t3 VTAIL.t6 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X10 B.t2 B.t0 B.t1 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=0 ps=0 w=9.87 l=1.24
X11 VDD2.t3 VN.t4 VTAIL.t5 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X12 VTAIL.t12 VP.t3 VDD1.t2 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X13 VDD1.t4 VP.t4 VTAIL.t11 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X14 VTAIL.t0 VN.t5 VDD2.t2 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X15 VDD2.t1 VN.t6 VTAIL.t4 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=3.8493 ps=20.52 w=9.87 l=1.24
X16 VTAIL.t10 VP.t5 VDD1.t7 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=3.8493 pd=20.52 as=1.62855 ps=10.2 w=9.87 l=1.24
X17 VDD1.t1 VP.t6 VTAIL.t9 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=3.8493 ps=20.52 w=9.87 l=1.24
X18 VDD1.t3 VP.t7 VTAIL.t8 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
X19 VTAIL.t3 VN.t7 VDD2.t0 w_n2540_n2942# sky130_fd_pr__pfet_01v8 ad=1.62855 pd=10.2 as=1.62855 ps=10.2 w=9.87 l=1.24
R0 B.n415 B.n414 585
R1 B.n416 B.n61 585
R2 B.n418 B.n417 585
R3 B.n419 B.n60 585
R4 B.n421 B.n420 585
R5 B.n422 B.n59 585
R6 B.n424 B.n423 585
R7 B.n425 B.n58 585
R8 B.n427 B.n426 585
R9 B.n428 B.n57 585
R10 B.n430 B.n429 585
R11 B.n431 B.n56 585
R12 B.n433 B.n432 585
R13 B.n434 B.n55 585
R14 B.n436 B.n435 585
R15 B.n437 B.n54 585
R16 B.n439 B.n438 585
R17 B.n440 B.n53 585
R18 B.n442 B.n441 585
R19 B.n443 B.n52 585
R20 B.n445 B.n444 585
R21 B.n446 B.n51 585
R22 B.n448 B.n447 585
R23 B.n449 B.n50 585
R24 B.n451 B.n450 585
R25 B.n452 B.n49 585
R26 B.n454 B.n453 585
R27 B.n455 B.n48 585
R28 B.n457 B.n456 585
R29 B.n458 B.n47 585
R30 B.n460 B.n459 585
R31 B.n461 B.n46 585
R32 B.n463 B.n462 585
R33 B.n464 B.n45 585
R34 B.n466 B.n465 585
R35 B.n468 B.n467 585
R36 B.n469 B.n41 585
R37 B.n471 B.n470 585
R38 B.n472 B.n40 585
R39 B.n474 B.n473 585
R40 B.n475 B.n39 585
R41 B.n477 B.n476 585
R42 B.n478 B.n38 585
R43 B.n480 B.n479 585
R44 B.n481 B.n35 585
R45 B.n484 B.n483 585
R46 B.n485 B.n34 585
R47 B.n487 B.n486 585
R48 B.n488 B.n33 585
R49 B.n490 B.n489 585
R50 B.n491 B.n32 585
R51 B.n493 B.n492 585
R52 B.n494 B.n31 585
R53 B.n496 B.n495 585
R54 B.n497 B.n30 585
R55 B.n499 B.n498 585
R56 B.n500 B.n29 585
R57 B.n502 B.n501 585
R58 B.n503 B.n28 585
R59 B.n505 B.n504 585
R60 B.n506 B.n27 585
R61 B.n508 B.n507 585
R62 B.n509 B.n26 585
R63 B.n511 B.n510 585
R64 B.n512 B.n25 585
R65 B.n514 B.n513 585
R66 B.n515 B.n24 585
R67 B.n517 B.n516 585
R68 B.n518 B.n23 585
R69 B.n520 B.n519 585
R70 B.n521 B.n22 585
R71 B.n523 B.n522 585
R72 B.n524 B.n21 585
R73 B.n526 B.n525 585
R74 B.n527 B.n20 585
R75 B.n529 B.n528 585
R76 B.n530 B.n19 585
R77 B.n532 B.n531 585
R78 B.n533 B.n18 585
R79 B.n535 B.n534 585
R80 B.n413 B.n62 585
R81 B.n412 B.n411 585
R82 B.n410 B.n63 585
R83 B.n409 B.n408 585
R84 B.n407 B.n64 585
R85 B.n406 B.n405 585
R86 B.n404 B.n65 585
R87 B.n403 B.n402 585
R88 B.n401 B.n66 585
R89 B.n400 B.n399 585
R90 B.n398 B.n67 585
R91 B.n397 B.n396 585
R92 B.n395 B.n68 585
R93 B.n394 B.n393 585
R94 B.n392 B.n69 585
R95 B.n391 B.n390 585
R96 B.n389 B.n70 585
R97 B.n388 B.n387 585
R98 B.n386 B.n71 585
R99 B.n385 B.n384 585
R100 B.n383 B.n72 585
R101 B.n382 B.n381 585
R102 B.n380 B.n73 585
R103 B.n379 B.n378 585
R104 B.n377 B.n74 585
R105 B.n376 B.n375 585
R106 B.n374 B.n75 585
R107 B.n373 B.n372 585
R108 B.n371 B.n76 585
R109 B.n370 B.n369 585
R110 B.n368 B.n77 585
R111 B.n367 B.n366 585
R112 B.n365 B.n78 585
R113 B.n364 B.n363 585
R114 B.n362 B.n79 585
R115 B.n361 B.n360 585
R116 B.n359 B.n80 585
R117 B.n358 B.n357 585
R118 B.n356 B.n81 585
R119 B.n355 B.n354 585
R120 B.n353 B.n82 585
R121 B.n352 B.n351 585
R122 B.n350 B.n83 585
R123 B.n349 B.n348 585
R124 B.n347 B.n84 585
R125 B.n346 B.n345 585
R126 B.n344 B.n85 585
R127 B.n343 B.n342 585
R128 B.n341 B.n86 585
R129 B.n340 B.n339 585
R130 B.n338 B.n87 585
R131 B.n337 B.n336 585
R132 B.n335 B.n88 585
R133 B.n334 B.n333 585
R134 B.n332 B.n89 585
R135 B.n331 B.n330 585
R136 B.n329 B.n90 585
R137 B.n328 B.n327 585
R138 B.n326 B.n91 585
R139 B.n325 B.n324 585
R140 B.n323 B.n92 585
R141 B.n322 B.n321 585
R142 B.n320 B.n93 585
R143 B.n199 B.n198 585
R144 B.n200 B.n137 585
R145 B.n202 B.n201 585
R146 B.n203 B.n136 585
R147 B.n205 B.n204 585
R148 B.n206 B.n135 585
R149 B.n208 B.n207 585
R150 B.n209 B.n134 585
R151 B.n211 B.n210 585
R152 B.n212 B.n133 585
R153 B.n214 B.n213 585
R154 B.n215 B.n132 585
R155 B.n217 B.n216 585
R156 B.n218 B.n131 585
R157 B.n220 B.n219 585
R158 B.n221 B.n130 585
R159 B.n223 B.n222 585
R160 B.n224 B.n129 585
R161 B.n226 B.n225 585
R162 B.n227 B.n128 585
R163 B.n229 B.n228 585
R164 B.n230 B.n127 585
R165 B.n232 B.n231 585
R166 B.n233 B.n126 585
R167 B.n235 B.n234 585
R168 B.n236 B.n125 585
R169 B.n238 B.n237 585
R170 B.n239 B.n124 585
R171 B.n241 B.n240 585
R172 B.n242 B.n123 585
R173 B.n244 B.n243 585
R174 B.n245 B.n122 585
R175 B.n247 B.n246 585
R176 B.n248 B.n121 585
R177 B.n250 B.n249 585
R178 B.n252 B.n251 585
R179 B.n253 B.n117 585
R180 B.n255 B.n254 585
R181 B.n256 B.n116 585
R182 B.n258 B.n257 585
R183 B.n259 B.n115 585
R184 B.n261 B.n260 585
R185 B.n262 B.n114 585
R186 B.n264 B.n263 585
R187 B.n265 B.n111 585
R188 B.n268 B.n267 585
R189 B.n269 B.n110 585
R190 B.n271 B.n270 585
R191 B.n272 B.n109 585
R192 B.n274 B.n273 585
R193 B.n275 B.n108 585
R194 B.n277 B.n276 585
R195 B.n278 B.n107 585
R196 B.n280 B.n279 585
R197 B.n281 B.n106 585
R198 B.n283 B.n282 585
R199 B.n284 B.n105 585
R200 B.n286 B.n285 585
R201 B.n287 B.n104 585
R202 B.n289 B.n288 585
R203 B.n290 B.n103 585
R204 B.n292 B.n291 585
R205 B.n293 B.n102 585
R206 B.n295 B.n294 585
R207 B.n296 B.n101 585
R208 B.n298 B.n297 585
R209 B.n299 B.n100 585
R210 B.n301 B.n300 585
R211 B.n302 B.n99 585
R212 B.n304 B.n303 585
R213 B.n305 B.n98 585
R214 B.n307 B.n306 585
R215 B.n308 B.n97 585
R216 B.n310 B.n309 585
R217 B.n311 B.n96 585
R218 B.n313 B.n312 585
R219 B.n314 B.n95 585
R220 B.n316 B.n315 585
R221 B.n317 B.n94 585
R222 B.n319 B.n318 585
R223 B.n197 B.n138 585
R224 B.n196 B.n195 585
R225 B.n194 B.n139 585
R226 B.n193 B.n192 585
R227 B.n191 B.n140 585
R228 B.n190 B.n189 585
R229 B.n188 B.n141 585
R230 B.n187 B.n186 585
R231 B.n185 B.n142 585
R232 B.n184 B.n183 585
R233 B.n182 B.n143 585
R234 B.n181 B.n180 585
R235 B.n179 B.n144 585
R236 B.n178 B.n177 585
R237 B.n176 B.n145 585
R238 B.n175 B.n174 585
R239 B.n173 B.n146 585
R240 B.n172 B.n171 585
R241 B.n170 B.n147 585
R242 B.n169 B.n168 585
R243 B.n167 B.n148 585
R244 B.n166 B.n165 585
R245 B.n164 B.n149 585
R246 B.n163 B.n162 585
R247 B.n161 B.n150 585
R248 B.n160 B.n159 585
R249 B.n158 B.n151 585
R250 B.n157 B.n156 585
R251 B.n155 B.n152 585
R252 B.n154 B.n153 585
R253 B.n2 B.n0 585
R254 B.n581 B.n1 585
R255 B.n580 B.n579 585
R256 B.n578 B.n3 585
R257 B.n577 B.n576 585
R258 B.n575 B.n4 585
R259 B.n574 B.n573 585
R260 B.n572 B.n5 585
R261 B.n571 B.n570 585
R262 B.n569 B.n6 585
R263 B.n568 B.n567 585
R264 B.n566 B.n7 585
R265 B.n565 B.n564 585
R266 B.n563 B.n8 585
R267 B.n562 B.n561 585
R268 B.n560 B.n9 585
R269 B.n559 B.n558 585
R270 B.n557 B.n10 585
R271 B.n556 B.n555 585
R272 B.n554 B.n11 585
R273 B.n553 B.n552 585
R274 B.n551 B.n12 585
R275 B.n550 B.n549 585
R276 B.n548 B.n13 585
R277 B.n547 B.n546 585
R278 B.n545 B.n14 585
R279 B.n544 B.n543 585
R280 B.n542 B.n15 585
R281 B.n541 B.n540 585
R282 B.n539 B.n16 585
R283 B.n538 B.n537 585
R284 B.n536 B.n17 585
R285 B.n583 B.n582 585
R286 B.n198 B.n197 554.963
R287 B.n534 B.n17 554.963
R288 B.n318 B.n93 554.963
R289 B.n414 B.n413 554.963
R290 B.n112 B.t3 396.149
R291 B.n118 B.t0 396.149
R292 B.n36 B.t9 396.149
R293 B.n42 B.t6 396.149
R294 B.n112 B.t5 367.503
R295 B.n42 B.t7 367.503
R296 B.n118 B.t2 367.503
R297 B.n36 B.t10 367.503
R298 B.n113 B.t4 337.055
R299 B.n43 B.t8 337.055
R300 B.n119 B.t1 337.055
R301 B.n37 B.t11 337.055
R302 B.n197 B.n196 163.367
R303 B.n196 B.n139 163.367
R304 B.n192 B.n139 163.367
R305 B.n192 B.n191 163.367
R306 B.n191 B.n190 163.367
R307 B.n190 B.n141 163.367
R308 B.n186 B.n141 163.367
R309 B.n186 B.n185 163.367
R310 B.n185 B.n184 163.367
R311 B.n184 B.n143 163.367
R312 B.n180 B.n143 163.367
R313 B.n180 B.n179 163.367
R314 B.n179 B.n178 163.367
R315 B.n178 B.n145 163.367
R316 B.n174 B.n145 163.367
R317 B.n174 B.n173 163.367
R318 B.n173 B.n172 163.367
R319 B.n172 B.n147 163.367
R320 B.n168 B.n147 163.367
R321 B.n168 B.n167 163.367
R322 B.n167 B.n166 163.367
R323 B.n166 B.n149 163.367
R324 B.n162 B.n149 163.367
R325 B.n162 B.n161 163.367
R326 B.n161 B.n160 163.367
R327 B.n160 B.n151 163.367
R328 B.n156 B.n151 163.367
R329 B.n156 B.n155 163.367
R330 B.n155 B.n154 163.367
R331 B.n154 B.n2 163.367
R332 B.n582 B.n2 163.367
R333 B.n582 B.n581 163.367
R334 B.n581 B.n580 163.367
R335 B.n580 B.n3 163.367
R336 B.n576 B.n3 163.367
R337 B.n576 B.n575 163.367
R338 B.n575 B.n574 163.367
R339 B.n574 B.n5 163.367
R340 B.n570 B.n5 163.367
R341 B.n570 B.n569 163.367
R342 B.n569 B.n568 163.367
R343 B.n568 B.n7 163.367
R344 B.n564 B.n7 163.367
R345 B.n564 B.n563 163.367
R346 B.n563 B.n562 163.367
R347 B.n562 B.n9 163.367
R348 B.n558 B.n9 163.367
R349 B.n558 B.n557 163.367
R350 B.n557 B.n556 163.367
R351 B.n556 B.n11 163.367
R352 B.n552 B.n11 163.367
R353 B.n552 B.n551 163.367
R354 B.n551 B.n550 163.367
R355 B.n550 B.n13 163.367
R356 B.n546 B.n13 163.367
R357 B.n546 B.n545 163.367
R358 B.n545 B.n544 163.367
R359 B.n544 B.n15 163.367
R360 B.n540 B.n15 163.367
R361 B.n540 B.n539 163.367
R362 B.n539 B.n538 163.367
R363 B.n538 B.n17 163.367
R364 B.n198 B.n137 163.367
R365 B.n202 B.n137 163.367
R366 B.n203 B.n202 163.367
R367 B.n204 B.n203 163.367
R368 B.n204 B.n135 163.367
R369 B.n208 B.n135 163.367
R370 B.n209 B.n208 163.367
R371 B.n210 B.n209 163.367
R372 B.n210 B.n133 163.367
R373 B.n214 B.n133 163.367
R374 B.n215 B.n214 163.367
R375 B.n216 B.n215 163.367
R376 B.n216 B.n131 163.367
R377 B.n220 B.n131 163.367
R378 B.n221 B.n220 163.367
R379 B.n222 B.n221 163.367
R380 B.n222 B.n129 163.367
R381 B.n226 B.n129 163.367
R382 B.n227 B.n226 163.367
R383 B.n228 B.n227 163.367
R384 B.n228 B.n127 163.367
R385 B.n232 B.n127 163.367
R386 B.n233 B.n232 163.367
R387 B.n234 B.n233 163.367
R388 B.n234 B.n125 163.367
R389 B.n238 B.n125 163.367
R390 B.n239 B.n238 163.367
R391 B.n240 B.n239 163.367
R392 B.n240 B.n123 163.367
R393 B.n244 B.n123 163.367
R394 B.n245 B.n244 163.367
R395 B.n246 B.n245 163.367
R396 B.n246 B.n121 163.367
R397 B.n250 B.n121 163.367
R398 B.n251 B.n250 163.367
R399 B.n251 B.n117 163.367
R400 B.n255 B.n117 163.367
R401 B.n256 B.n255 163.367
R402 B.n257 B.n256 163.367
R403 B.n257 B.n115 163.367
R404 B.n261 B.n115 163.367
R405 B.n262 B.n261 163.367
R406 B.n263 B.n262 163.367
R407 B.n263 B.n111 163.367
R408 B.n268 B.n111 163.367
R409 B.n269 B.n268 163.367
R410 B.n270 B.n269 163.367
R411 B.n270 B.n109 163.367
R412 B.n274 B.n109 163.367
R413 B.n275 B.n274 163.367
R414 B.n276 B.n275 163.367
R415 B.n276 B.n107 163.367
R416 B.n280 B.n107 163.367
R417 B.n281 B.n280 163.367
R418 B.n282 B.n281 163.367
R419 B.n282 B.n105 163.367
R420 B.n286 B.n105 163.367
R421 B.n287 B.n286 163.367
R422 B.n288 B.n287 163.367
R423 B.n288 B.n103 163.367
R424 B.n292 B.n103 163.367
R425 B.n293 B.n292 163.367
R426 B.n294 B.n293 163.367
R427 B.n294 B.n101 163.367
R428 B.n298 B.n101 163.367
R429 B.n299 B.n298 163.367
R430 B.n300 B.n299 163.367
R431 B.n300 B.n99 163.367
R432 B.n304 B.n99 163.367
R433 B.n305 B.n304 163.367
R434 B.n306 B.n305 163.367
R435 B.n306 B.n97 163.367
R436 B.n310 B.n97 163.367
R437 B.n311 B.n310 163.367
R438 B.n312 B.n311 163.367
R439 B.n312 B.n95 163.367
R440 B.n316 B.n95 163.367
R441 B.n317 B.n316 163.367
R442 B.n318 B.n317 163.367
R443 B.n322 B.n93 163.367
R444 B.n323 B.n322 163.367
R445 B.n324 B.n323 163.367
R446 B.n324 B.n91 163.367
R447 B.n328 B.n91 163.367
R448 B.n329 B.n328 163.367
R449 B.n330 B.n329 163.367
R450 B.n330 B.n89 163.367
R451 B.n334 B.n89 163.367
R452 B.n335 B.n334 163.367
R453 B.n336 B.n335 163.367
R454 B.n336 B.n87 163.367
R455 B.n340 B.n87 163.367
R456 B.n341 B.n340 163.367
R457 B.n342 B.n341 163.367
R458 B.n342 B.n85 163.367
R459 B.n346 B.n85 163.367
R460 B.n347 B.n346 163.367
R461 B.n348 B.n347 163.367
R462 B.n348 B.n83 163.367
R463 B.n352 B.n83 163.367
R464 B.n353 B.n352 163.367
R465 B.n354 B.n353 163.367
R466 B.n354 B.n81 163.367
R467 B.n358 B.n81 163.367
R468 B.n359 B.n358 163.367
R469 B.n360 B.n359 163.367
R470 B.n360 B.n79 163.367
R471 B.n364 B.n79 163.367
R472 B.n365 B.n364 163.367
R473 B.n366 B.n365 163.367
R474 B.n366 B.n77 163.367
R475 B.n370 B.n77 163.367
R476 B.n371 B.n370 163.367
R477 B.n372 B.n371 163.367
R478 B.n372 B.n75 163.367
R479 B.n376 B.n75 163.367
R480 B.n377 B.n376 163.367
R481 B.n378 B.n377 163.367
R482 B.n378 B.n73 163.367
R483 B.n382 B.n73 163.367
R484 B.n383 B.n382 163.367
R485 B.n384 B.n383 163.367
R486 B.n384 B.n71 163.367
R487 B.n388 B.n71 163.367
R488 B.n389 B.n388 163.367
R489 B.n390 B.n389 163.367
R490 B.n390 B.n69 163.367
R491 B.n394 B.n69 163.367
R492 B.n395 B.n394 163.367
R493 B.n396 B.n395 163.367
R494 B.n396 B.n67 163.367
R495 B.n400 B.n67 163.367
R496 B.n401 B.n400 163.367
R497 B.n402 B.n401 163.367
R498 B.n402 B.n65 163.367
R499 B.n406 B.n65 163.367
R500 B.n407 B.n406 163.367
R501 B.n408 B.n407 163.367
R502 B.n408 B.n63 163.367
R503 B.n412 B.n63 163.367
R504 B.n413 B.n412 163.367
R505 B.n534 B.n533 163.367
R506 B.n533 B.n532 163.367
R507 B.n532 B.n19 163.367
R508 B.n528 B.n19 163.367
R509 B.n528 B.n527 163.367
R510 B.n527 B.n526 163.367
R511 B.n526 B.n21 163.367
R512 B.n522 B.n21 163.367
R513 B.n522 B.n521 163.367
R514 B.n521 B.n520 163.367
R515 B.n520 B.n23 163.367
R516 B.n516 B.n23 163.367
R517 B.n516 B.n515 163.367
R518 B.n515 B.n514 163.367
R519 B.n514 B.n25 163.367
R520 B.n510 B.n25 163.367
R521 B.n510 B.n509 163.367
R522 B.n509 B.n508 163.367
R523 B.n508 B.n27 163.367
R524 B.n504 B.n27 163.367
R525 B.n504 B.n503 163.367
R526 B.n503 B.n502 163.367
R527 B.n502 B.n29 163.367
R528 B.n498 B.n29 163.367
R529 B.n498 B.n497 163.367
R530 B.n497 B.n496 163.367
R531 B.n496 B.n31 163.367
R532 B.n492 B.n31 163.367
R533 B.n492 B.n491 163.367
R534 B.n491 B.n490 163.367
R535 B.n490 B.n33 163.367
R536 B.n486 B.n33 163.367
R537 B.n486 B.n485 163.367
R538 B.n485 B.n484 163.367
R539 B.n484 B.n35 163.367
R540 B.n479 B.n35 163.367
R541 B.n479 B.n478 163.367
R542 B.n478 B.n477 163.367
R543 B.n477 B.n39 163.367
R544 B.n473 B.n39 163.367
R545 B.n473 B.n472 163.367
R546 B.n472 B.n471 163.367
R547 B.n471 B.n41 163.367
R548 B.n467 B.n41 163.367
R549 B.n467 B.n466 163.367
R550 B.n466 B.n45 163.367
R551 B.n462 B.n45 163.367
R552 B.n462 B.n461 163.367
R553 B.n461 B.n460 163.367
R554 B.n460 B.n47 163.367
R555 B.n456 B.n47 163.367
R556 B.n456 B.n455 163.367
R557 B.n455 B.n454 163.367
R558 B.n454 B.n49 163.367
R559 B.n450 B.n49 163.367
R560 B.n450 B.n449 163.367
R561 B.n449 B.n448 163.367
R562 B.n448 B.n51 163.367
R563 B.n444 B.n51 163.367
R564 B.n444 B.n443 163.367
R565 B.n443 B.n442 163.367
R566 B.n442 B.n53 163.367
R567 B.n438 B.n53 163.367
R568 B.n438 B.n437 163.367
R569 B.n437 B.n436 163.367
R570 B.n436 B.n55 163.367
R571 B.n432 B.n55 163.367
R572 B.n432 B.n431 163.367
R573 B.n431 B.n430 163.367
R574 B.n430 B.n57 163.367
R575 B.n426 B.n57 163.367
R576 B.n426 B.n425 163.367
R577 B.n425 B.n424 163.367
R578 B.n424 B.n59 163.367
R579 B.n420 B.n59 163.367
R580 B.n420 B.n419 163.367
R581 B.n419 B.n418 163.367
R582 B.n418 B.n61 163.367
R583 B.n414 B.n61 163.367
R584 B.n266 B.n113 59.5399
R585 B.n120 B.n119 59.5399
R586 B.n482 B.n37 59.5399
R587 B.n44 B.n43 59.5399
R588 B.n536 B.n535 36.059
R589 B.n415 B.n62 36.059
R590 B.n320 B.n319 36.059
R591 B.n199 B.n138 36.059
R592 B.n113 B.n112 30.449
R593 B.n119 B.n118 30.449
R594 B.n37 B.n36 30.449
R595 B.n43 B.n42 30.449
R596 B B.n583 18.0485
R597 B.n535 B.n18 10.6151
R598 B.n531 B.n18 10.6151
R599 B.n531 B.n530 10.6151
R600 B.n530 B.n529 10.6151
R601 B.n529 B.n20 10.6151
R602 B.n525 B.n20 10.6151
R603 B.n525 B.n524 10.6151
R604 B.n524 B.n523 10.6151
R605 B.n523 B.n22 10.6151
R606 B.n519 B.n22 10.6151
R607 B.n519 B.n518 10.6151
R608 B.n518 B.n517 10.6151
R609 B.n517 B.n24 10.6151
R610 B.n513 B.n24 10.6151
R611 B.n513 B.n512 10.6151
R612 B.n512 B.n511 10.6151
R613 B.n511 B.n26 10.6151
R614 B.n507 B.n26 10.6151
R615 B.n507 B.n506 10.6151
R616 B.n506 B.n505 10.6151
R617 B.n505 B.n28 10.6151
R618 B.n501 B.n28 10.6151
R619 B.n501 B.n500 10.6151
R620 B.n500 B.n499 10.6151
R621 B.n499 B.n30 10.6151
R622 B.n495 B.n30 10.6151
R623 B.n495 B.n494 10.6151
R624 B.n494 B.n493 10.6151
R625 B.n493 B.n32 10.6151
R626 B.n489 B.n32 10.6151
R627 B.n489 B.n488 10.6151
R628 B.n488 B.n487 10.6151
R629 B.n487 B.n34 10.6151
R630 B.n483 B.n34 10.6151
R631 B.n481 B.n480 10.6151
R632 B.n480 B.n38 10.6151
R633 B.n476 B.n38 10.6151
R634 B.n476 B.n475 10.6151
R635 B.n475 B.n474 10.6151
R636 B.n474 B.n40 10.6151
R637 B.n470 B.n40 10.6151
R638 B.n470 B.n469 10.6151
R639 B.n469 B.n468 10.6151
R640 B.n465 B.n464 10.6151
R641 B.n464 B.n463 10.6151
R642 B.n463 B.n46 10.6151
R643 B.n459 B.n46 10.6151
R644 B.n459 B.n458 10.6151
R645 B.n458 B.n457 10.6151
R646 B.n457 B.n48 10.6151
R647 B.n453 B.n48 10.6151
R648 B.n453 B.n452 10.6151
R649 B.n452 B.n451 10.6151
R650 B.n451 B.n50 10.6151
R651 B.n447 B.n50 10.6151
R652 B.n447 B.n446 10.6151
R653 B.n446 B.n445 10.6151
R654 B.n445 B.n52 10.6151
R655 B.n441 B.n52 10.6151
R656 B.n441 B.n440 10.6151
R657 B.n440 B.n439 10.6151
R658 B.n439 B.n54 10.6151
R659 B.n435 B.n54 10.6151
R660 B.n435 B.n434 10.6151
R661 B.n434 B.n433 10.6151
R662 B.n433 B.n56 10.6151
R663 B.n429 B.n56 10.6151
R664 B.n429 B.n428 10.6151
R665 B.n428 B.n427 10.6151
R666 B.n427 B.n58 10.6151
R667 B.n423 B.n58 10.6151
R668 B.n423 B.n422 10.6151
R669 B.n422 B.n421 10.6151
R670 B.n421 B.n60 10.6151
R671 B.n417 B.n60 10.6151
R672 B.n417 B.n416 10.6151
R673 B.n416 B.n415 10.6151
R674 B.n321 B.n320 10.6151
R675 B.n321 B.n92 10.6151
R676 B.n325 B.n92 10.6151
R677 B.n326 B.n325 10.6151
R678 B.n327 B.n326 10.6151
R679 B.n327 B.n90 10.6151
R680 B.n331 B.n90 10.6151
R681 B.n332 B.n331 10.6151
R682 B.n333 B.n332 10.6151
R683 B.n333 B.n88 10.6151
R684 B.n337 B.n88 10.6151
R685 B.n338 B.n337 10.6151
R686 B.n339 B.n338 10.6151
R687 B.n339 B.n86 10.6151
R688 B.n343 B.n86 10.6151
R689 B.n344 B.n343 10.6151
R690 B.n345 B.n344 10.6151
R691 B.n345 B.n84 10.6151
R692 B.n349 B.n84 10.6151
R693 B.n350 B.n349 10.6151
R694 B.n351 B.n350 10.6151
R695 B.n351 B.n82 10.6151
R696 B.n355 B.n82 10.6151
R697 B.n356 B.n355 10.6151
R698 B.n357 B.n356 10.6151
R699 B.n357 B.n80 10.6151
R700 B.n361 B.n80 10.6151
R701 B.n362 B.n361 10.6151
R702 B.n363 B.n362 10.6151
R703 B.n363 B.n78 10.6151
R704 B.n367 B.n78 10.6151
R705 B.n368 B.n367 10.6151
R706 B.n369 B.n368 10.6151
R707 B.n369 B.n76 10.6151
R708 B.n373 B.n76 10.6151
R709 B.n374 B.n373 10.6151
R710 B.n375 B.n374 10.6151
R711 B.n375 B.n74 10.6151
R712 B.n379 B.n74 10.6151
R713 B.n380 B.n379 10.6151
R714 B.n381 B.n380 10.6151
R715 B.n381 B.n72 10.6151
R716 B.n385 B.n72 10.6151
R717 B.n386 B.n385 10.6151
R718 B.n387 B.n386 10.6151
R719 B.n387 B.n70 10.6151
R720 B.n391 B.n70 10.6151
R721 B.n392 B.n391 10.6151
R722 B.n393 B.n392 10.6151
R723 B.n393 B.n68 10.6151
R724 B.n397 B.n68 10.6151
R725 B.n398 B.n397 10.6151
R726 B.n399 B.n398 10.6151
R727 B.n399 B.n66 10.6151
R728 B.n403 B.n66 10.6151
R729 B.n404 B.n403 10.6151
R730 B.n405 B.n404 10.6151
R731 B.n405 B.n64 10.6151
R732 B.n409 B.n64 10.6151
R733 B.n410 B.n409 10.6151
R734 B.n411 B.n410 10.6151
R735 B.n411 B.n62 10.6151
R736 B.n200 B.n199 10.6151
R737 B.n201 B.n200 10.6151
R738 B.n201 B.n136 10.6151
R739 B.n205 B.n136 10.6151
R740 B.n206 B.n205 10.6151
R741 B.n207 B.n206 10.6151
R742 B.n207 B.n134 10.6151
R743 B.n211 B.n134 10.6151
R744 B.n212 B.n211 10.6151
R745 B.n213 B.n212 10.6151
R746 B.n213 B.n132 10.6151
R747 B.n217 B.n132 10.6151
R748 B.n218 B.n217 10.6151
R749 B.n219 B.n218 10.6151
R750 B.n219 B.n130 10.6151
R751 B.n223 B.n130 10.6151
R752 B.n224 B.n223 10.6151
R753 B.n225 B.n224 10.6151
R754 B.n225 B.n128 10.6151
R755 B.n229 B.n128 10.6151
R756 B.n230 B.n229 10.6151
R757 B.n231 B.n230 10.6151
R758 B.n231 B.n126 10.6151
R759 B.n235 B.n126 10.6151
R760 B.n236 B.n235 10.6151
R761 B.n237 B.n236 10.6151
R762 B.n237 B.n124 10.6151
R763 B.n241 B.n124 10.6151
R764 B.n242 B.n241 10.6151
R765 B.n243 B.n242 10.6151
R766 B.n243 B.n122 10.6151
R767 B.n247 B.n122 10.6151
R768 B.n248 B.n247 10.6151
R769 B.n249 B.n248 10.6151
R770 B.n253 B.n252 10.6151
R771 B.n254 B.n253 10.6151
R772 B.n254 B.n116 10.6151
R773 B.n258 B.n116 10.6151
R774 B.n259 B.n258 10.6151
R775 B.n260 B.n259 10.6151
R776 B.n260 B.n114 10.6151
R777 B.n264 B.n114 10.6151
R778 B.n265 B.n264 10.6151
R779 B.n267 B.n110 10.6151
R780 B.n271 B.n110 10.6151
R781 B.n272 B.n271 10.6151
R782 B.n273 B.n272 10.6151
R783 B.n273 B.n108 10.6151
R784 B.n277 B.n108 10.6151
R785 B.n278 B.n277 10.6151
R786 B.n279 B.n278 10.6151
R787 B.n279 B.n106 10.6151
R788 B.n283 B.n106 10.6151
R789 B.n284 B.n283 10.6151
R790 B.n285 B.n284 10.6151
R791 B.n285 B.n104 10.6151
R792 B.n289 B.n104 10.6151
R793 B.n290 B.n289 10.6151
R794 B.n291 B.n290 10.6151
R795 B.n291 B.n102 10.6151
R796 B.n295 B.n102 10.6151
R797 B.n296 B.n295 10.6151
R798 B.n297 B.n296 10.6151
R799 B.n297 B.n100 10.6151
R800 B.n301 B.n100 10.6151
R801 B.n302 B.n301 10.6151
R802 B.n303 B.n302 10.6151
R803 B.n303 B.n98 10.6151
R804 B.n307 B.n98 10.6151
R805 B.n308 B.n307 10.6151
R806 B.n309 B.n308 10.6151
R807 B.n309 B.n96 10.6151
R808 B.n313 B.n96 10.6151
R809 B.n314 B.n313 10.6151
R810 B.n315 B.n314 10.6151
R811 B.n315 B.n94 10.6151
R812 B.n319 B.n94 10.6151
R813 B.n195 B.n138 10.6151
R814 B.n195 B.n194 10.6151
R815 B.n194 B.n193 10.6151
R816 B.n193 B.n140 10.6151
R817 B.n189 B.n140 10.6151
R818 B.n189 B.n188 10.6151
R819 B.n188 B.n187 10.6151
R820 B.n187 B.n142 10.6151
R821 B.n183 B.n142 10.6151
R822 B.n183 B.n182 10.6151
R823 B.n182 B.n181 10.6151
R824 B.n181 B.n144 10.6151
R825 B.n177 B.n144 10.6151
R826 B.n177 B.n176 10.6151
R827 B.n176 B.n175 10.6151
R828 B.n175 B.n146 10.6151
R829 B.n171 B.n146 10.6151
R830 B.n171 B.n170 10.6151
R831 B.n170 B.n169 10.6151
R832 B.n169 B.n148 10.6151
R833 B.n165 B.n148 10.6151
R834 B.n165 B.n164 10.6151
R835 B.n164 B.n163 10.6151
R836 B.n163 B.n150 10.6151
R837 B.n159 B.n150 10.6151
R838 B.n159 B.n158 10.6151
R839 B.n158 B.n157 10.6151
R840 B.n157 B.n152 10.6151
R841 B.n153 B.n152 10.6151
R842 B.n153 B.n0 10.6151
R843 B.n579 B.n1 10.6151
R844 B.n579 B.n578 10.6151
R845 B.n578 B.n577 10.6151
R846 B.n577 B.n4 10.6151
R847 B.n573 B.n4 10.6151
R848 B.n573 B.n572 10.6151
R849 B.n572 B.n571 10.6151
R850 B.n571 B.n6 10.6151
R851 B.n567 B.n6 10.6151
R852 B.n567 B.n566 10.6151
R853 B.n566 B.n565 10.6151
R854 B.n565 B.n8 10.6151
R855 B.n561 B.n8 10.6151
R856 B.n561 B.n560 10.6151
R857 B.n560 B.n559 10.6151
R858 B.n559 B.n10 10.6151
R859 B.n555 B.n10 10.6151
R860 B.n555 B.n554 10.6151
R861 B.n554 B.n553 10.6151
R862 B.n553 B.n12 10.6151
R863 B.n549 B.n12 10.6151
R864 B.n549 B.n548 10.6151
R865 B.n548 B.n547 10.6151
R866 B.n547 B.n14 10.6151
R867 B.n543 B.n14 10.6151
R868 B.n543 B.n542 10.6151
R869 B.n542 B.n541 10.6151
R870 B.n541 B.n16 10.6151
R871 B.n537 B.n16 10.6151
R872 B.n537 B.n536 10.6151
R873 B.n483 B.n482 9.36635
R874 B.n465 B.n44 9.36635
R875 B.n249 B.n120 9.36635
R876 B.n267 B.n266 9.36635
R877 B.n583 B.n0 2.81026
R878 B.n583 B.n1 2.81026
R879 B.n482 B.n481 1.24928
R880 B.n468 B.n44 1.24928
R881 B.n252 B.n120 1.24928
R882 B.n266 B.n265 1.24928
R883 VP.n9 VP.t0 243.444
R884 VP.n21 VP.t5 223.702
R885 VP.n33 VP.t2 223.702
R886 VP.n18 VP.t6 223.702
R887 VP.n3 VP.t4 191.828
R888 VP.n1 VP.t3 191.828
R889 VP.n6 VP.t1 191.828
R890 VP.n8 VP.t7 191.828
R891 VP.n11 VP.n10 161.3
R892 VP.n12 VP.n7 161.3
R893 VP.n14 VP.n13 161.3
R894 VP.n16 VP.n15 161.3
R895 VP.n17 VP.n5 161.3
R896 VP.n32 VP.n0 161.3
R897 VP.n31 VP.n30 161.3
R898 VP.n29 VP.n28 161.3
R899 VP.n27 VP.n2 161.3
R900 VP.n26 VP.n25 161.3
R901 VP.n24 VP.n23 161.3
R902 VP.n22 VP.n4 161.3
R903 VP.n19 VP.n18 80.6037
R904 VP.n34 VP.n33 80.6037
R905 VP.n21 VP.n20 80.6037
R906 VP.n9 VP.n8 43.5433
R907 VP.n20 VP.n19 43.0847
R908 VP.n27 VP.n26 40.4934
R909 VP.n28 VP.n27 40.4934
R910 VP.n13 VP.n12 40.4934
R911 VP.n12 VP.n11 40.4934
R912 VP.n22 VP.n21 34.3247
R913 VP.n33 VP.n32 34.3247
R914 VP.n18 VP.n17 34.3247
R915 VP.n23 VP.n22 33.6945
R916 VP.n32 VP.n31 33.6945
R917 VP.n17 VP.n16 33.6945
R918 VP.n10 VP.n9 29.3131
R919 VP.n26 VP.n3 13.9467
R920 VP.n28 VP.n1 13.9467
R921 VP.n13 VP.n6 13.9467
R922 VP.n11 VP.n8 13.9467
R923 VP.n23 VP.n3 10.5213
R924 VP.n31 VP.n1 10.5213
R925 VP.n16 VP.n6 10.5213
R926 VP.n19 VP.n5 0.285035
R927 VP.n20 VP.n4 0.285035
R928 VP.n34 VP.n0 0.285035
R929 VP.n10 VP.n7 0.189894
R930 VP.n14 VP.n7 0.189894
R931 VP.n15 VP.n14 0.189894
R932 VP.n15 VP.n5 0.189894
R933 VP.n24 VP.n4 0.189894
R934 VP.n25 VP.n24 0.189894
R935 VP.n25 VP.n2 0.189894
R936 VP.n29 VP.n2 0.189894
R937 VP.n30 VP.n29 0.189894
R938 VP.n30 VP.n0 0.189894
R939 VP VP.n34 0.146778
R940 VDD1 VDD1.n0 76.1084
R941 VDD1.n3 VDD1.n2 75.9947
R942 VDD1.n3 VDD1.n1 75.9947
R943 VDD1.n5 VDD1.n4 75.3733
R944 VDD1.n5 VDD1.n3 38.8974
R945 VDD1.n4 VDD1.t6 3.29381
R946 VDD1.n4 VDD1.t1 3.29381
R947 VDD1.n0 VDD1.t5 3.29381
R948 VDD1.n0 VDD1.t3 3.29381
R949 VDD1.n2 VDD1.t2 3.29381
R950 VDD1.n2 VDD1.t0 3.29381
R951 VDD1.n1 VDD1.t7 3.29381
R952 VDD1.n1 VDD1.t4 3.29381
R953 VDD1 VDD1.n5 0.619035
R954 VTAIL.n434 VTAIL.n386 756.745
R955 VTAIL.n50 VTAIL.n2 756.745
R956 VTAIL.n104 VTAIL.n56 756.745
R957 VTAIL.n160 VTAIL.n112 756.745
R958 VTAIL.n380 VTAIL.n332 756.745
R959 VTAIL.n324 VTAIL.n276 756.745
R960 VTAIL.n270 VTAIL.n222 756.745
R961 VTAIL.n214 VTAIL.n166 756.745
R962 VTAIL.n402 VTAIL.n401 585
R963 VTAIL.n407 VTAIL.n406 585
R964 VTAIL.n409 VTAIL.n408 585
R965 VTAIL.n398 VTAIL.n397 585
R966 VTAIL.n415 VTAIL.n414 585
R967 VTAIL.n417 VTAIL.n416 585
R968 VTAIL.n394 VTAIL.n393 585
R969 VTAIL.n424 VTAIL.n423 585
R970 VTAIL.n425 VTAIL.n392 585
R971 VTAIL.n427 VTAIL.n426 585
R972 VTAIL.n390 VTAIL.n389 585
R973 VTAIL.n433 VTAIL.n432 585
R974 VTAIL.n435 VTAIL.n434 585
R975 VTAIL.n18 VTAIL.n17 585
R976 VTAIL.n23 VTAIL.n22 585
R977 VTAIL.n25 VTAIL.n24 585
R978 VTAIL.n14 VTAIL.n13 585
R979 VTAIL.n31 VTAIL.n30 585
R980 VTAIL.n33 VTAIL.n32 585
R981 VTAIL.n10 VTAIL.n9 585
R982 VTAIL.n40 VTAIL.n39 585
R983 VTAIL.n41 VTAIL.n8 585
R984 VTAIL.n43 VTAIL.n42 585
R985 VTAIL.n6 VTAIL.n5 585
R986 VTAIL.n49 VTAIL.n48 585
R987 VTAIL.n51 VTAIL.n50 585
R988 VTAIL.n72 VTAIL.n71 585
R989 VTAIL.n77 VTAIL.n76 585
R990 VTAIL.n79 VTAIL.n78 585
R991 VTAIL.n68 VTAIL.n67 585
R992 VTAIL.n85 VTAIL.n84 585
R993 VTAIL.n87 VTAIL.n86 585
R994 VTAIL.n64 VTAIL.n63 585
R995 VTAIL.n94 VTAIL.n93 585
R996 VTAIL.n95 VTAIL.n62 585
R997 VTAIL.n97 VTAIL.n96 585
R998 VTAIL.n60 VTAIL.n59 585
R999 VTAIL.n103 VTAIL.n102 585
R1000 VTAIL.n105 VTAIL.n104 585
R1001 VTAIL.n128 VTAIL.n127 585
R1002 VTAIL.n133 VTAIL.n132 585
R1003 VTAIL.n135 VTAIL.n134 585
R1004 VTAIL.n124 VTAIL.n123 585
R1005 VTAIL.n141 VTAIL.n140 585
R1006 VTAIL.n143 VTAIL.n142 585
R1007 VTAIL.n120 VTAIL.n119 585
R1008 VTAIL.n150 VTAIL.n149 585
R1009 VTAIL.n151 VTAIL.n118 585
R1010 VTAIL.n153 VTAIL.n152 585
R1011 VTAIL.n116 VTAIL.n115 585
R1012 VTAIL.n159 VTAIL.n158 585
R1013 VTAIL.n161 VTAIL.n160 585
R1014 VTAIL.n381 VTAIL.n380 585
R1015 VTAIL.n379 VTAIL.n378 585
R1016 VTAIL.n336 VTAIL.n335 585
R1017 VTAIL.n373 VTAIL.n372 585
R1018 VTAIL.n371 VTAIL.n338 585
R1019 VTAIL.n370 VTAIL.n369 585
R1020 VTAIL.n341 VTAIL.n339 585
R1021 VTAIL.n364 VTAIL.n363 585
R1022 VTAIL.n362 VTAIL.n361 585
R1023 VTAIL.n345 VTAIL.n344 585
R1024 VTAIL.n356 VTAIL.n355 585
R1025 VTAIL.n354 VTAIL.n353 585
R1026 VTAIL.n349 VTAIL.n348 585
R1027 VTAIL.n325 VTAIL.n324 585
R1028 VTAIL.n323 VTAIL.n322 585
R1029 VTAIL.n280 VTAIL.n279 585
R1030 VTAIL.n317 VTAIL.n316 585
R1031 VTAIL.n315 VTAIL.n282 585
R1032 VTAIL.n314 VTAIL.n313 585
R1033 VTAIL.n285 VTAIL.n283 585
R1034 VTAIL.n308 VTAIL.n307 585
R1035 VTAIL.n306 VTAIL.n305 585
R1036 VTAIL.n289 VTAIL.n288 585
R1037 VTAIL.n300 VTAIL.n299 585
R1038 VTAIL.n298 VTAIL.n297 585
R1039 VTAIL.n293 VTAIL.n292 585
R1040 VTAIL.n271 VTAIL.n270 585
R1041 VTAIL.n269 VTAIL.n268 585
R1042 VTAIL.n226 VTAIL.n225 585
R1043 VTAIL.n263 VTAIL.n262 585
R1044 VTAIL.n261 VTAIL.n228 585
R1045 VTAIL.n260 VTAIL.n259 585
R1046 VTAIL.n231 VTAIL.n229 585
R1047 VTAIL.n254 VTAIL.n253 585
R1048 VTAIL.n252 VTAIL.n251 585
R1049 VTAIL.n235 VTAIL.n234 585
R1050 VTAIL.n246 VTAIL.n245 585
R1051 VTAIL.n244 VTAIL.n243 585
R1052 VTAIL.n239 VTAIL.n238 585
R1053 VTAIL.n215 VTAIL.n214 585
R1054 VTAIL.n213 VTAIL.n212 585
R1055 VTAIL.n170 VTAIL.n169 585
R1056 VTAIL.n207 VTAIL.n206 585
R1057 VTAIL.n205 VTAIL.n172 585
R1058 VTAIL.n204 VTAIL.n203 585
R1059 VTAIL.n175 VTAIL.n173 585
R1060 VTAIL.n198 VTAIL.n197 585
R1061 VTAIL.n196 VTAIL.n195 585
R1062 VTAIL.n179 VTAIL.n178 585
R1063 VTAIL.n190 VTAIL.n189 585
R1064 VTAIL.n188 VTAIL.n187 585
R1065 VTAIL.n183 VTAIL.n182 585
R1066 VTAIL.n403 VTAIL.t4 329.038
R1067 VTAIL.n19 VTAIL.t1 329.038
R1068 VTAIL.n73 VTAIL.t13 329.038
R1069 VTAIL.n129 VTAIL.t10 329.038
R1070 VTAIL.n350 VTAIL.t9 329.038
R1071 VTAIL.n294 VTAIL.t15 329.038
R1072 VTAIL.n240 VTAIL.t2 329.038
R1073 VTAIL.n184 VTAIL.t7 329.038
R1074 VTAIL.n407 VTAIL.n401 171.744
R1075 VTAIL.n408 VTAIL.n407 171.744
R1076 VTAIL.n408 VTAIL.n397 171.744
R1077 VTAIL.n415 VTAIL.n397 171.744
R1078 VTAIL.n416 VTAIL.n415 171.744
R1079 VTAIL.n416 VTAIL.n393 171.744
R1080 VTAIL.n424 VTAIL.n393 171.744
R1081 VTAIL.n425 VTAIL.n424 171.744
R1082 VTAIL.n426 VTAIL.n425 171.744
R1083 VTAIL.n426 VTAIL.n389 171.744
R1084 VTAIL.n433 VTAIL.n389 171.744
R1085 VTAIL.n434 VTAIL.n433 171.744
R1086 VTAIL.n23 VTAIL.n17 171.744
R1087 VTAIL.n24 VTAIL.n23 171.744
R1088 VTAIL.n24 VTAIL.n13 171.744
R1089 VTAIL.n31 VTAIL.n13 171.744
R1090 VTAIL.n32 VTAIL.n31 171.744
R1091 VTAIL.n32 VTAIL.n9 171.744
R1092 VTAIL.n40 VTAIL.n9 171.744
R1093 VTAIL.n41 VTAIL.n40 171.744
R1094 VTAIL.n42 VTAIL.n41 171.744
R1095 VTAIL.n42 VTAIL.n5 171.744
R1096 VTAIL.n49 VTAIL.n5 171.744
R1097 VTAIL.n50 VTAIL.n49 171.744
R1098 VTAIL.n77 VTAIL.n71 171.744
R1099 VTAIL.n78 VTAIL.n77 171.744
R1100 VTAIL.n78 VTAIL.n67 171.744
R1101 VTAIL.n85 VTAIL.n67 171.744
R1102 VTAIL.n86 VTAIL.n85 171.744
R1103 VTAIL.n86 VTAIL.n63 171.744
R1104 VTAIL.n94 VTAIL.n63 171.744
R1105 VTAIL.n95 VTAIL.n94 171.744
R1106 VTAIL.n96 VTAIL.n95 171.744
R1107 VTAIL.n96 VTAIL.n59 171.744
R1108 VTAIL.n103 VTAIL.n59 171.744
R1109 VTAIL.n104 VTAIL.n103 171.744
R1110 VTAIL.n133 VTAIL.n127 171.744
R1111 VTAIL.n134 VTAIL.n133 171.744
R1112 VTAIL.n134 VTAIL.n123 171.744
R1113 VTAIL.n141 VTAIL.n123 171.744
R1114 VTAIL.n142 VTAIL.n141 171.744
R1115 VTAIL.n142 VTAIL.n119 171.744
R1116 VTAIL.n150 VTAIL.n119 171.744
R1117 VTAIL.n151 VTAIL.n150 171.744
R1118 VTAIL.n152 VTAIL.n151 171.744
R1119 VTAIL.n152 VTAIL.n115 171.744
R1120 VTAIL.n159 VTAIL.n115 171.744
R1121 VTAIL.n160 VTAIL.n159 171.744
R1122 VTAIL.n380 VTAIL.n379 171.744
R1123 VTAIL.n379 VTAIL.n335 171.744
R1124 VTAIL.n372 VTAIL.n335 171.744
R1125 VTAIL.n372 VTAIL.n371 171.744
R1126 VTAIL.n371 VTAIL.n370 171.744
R1127 VTAIL.n370 VTAIL.n339 171.744
R1128 VTAIL.n363 VTAIL.n339 171.744
R1129 VTAIL.n363 VTAIL.n362 171.744
R1130 VTAIL.n362 VTAIL.n344 171.744
R1131 VTAIL.n355 VTAIL.n344 171.744
R1132 VTAIL.n355 VTAIL.n354 171.744
R1133 VTAIL.n354 VTAIL.n348 171.744
R1134 VTAIL.n324 VTAIL.n323 171.744
R1135 VTAIL.n323 VTAIL.n279 171.744
R1136 VTAIL.n316 VTAIL.n279 171.744
R1137 VTAIL.n316 VTAIL.n315 171.744
R1138 VTAIL.n315 VTAIL.n314 171.744
R1139 VTAIL.n314 VTAIL.n283 171.744
R1140 VTAIL.n307 VTAIL.n283 171.744
R1141 VTAIL.n307 VTAIL.n306 171.744
R1142 VTAIL.n306 VTAIL.n288 171.744
R1143 VTAIL.n299 VTAIL.n288 171.744
R1144 VTAIL.n299 VTAIL.n298 171.744
R1145 VTAIL.n298 VTAIL.n292 171.744
R1146 VTAIL.n270 VTAIL.n269 171.744
R1147 VTAIL.n269 VTAIL.n225 171.744
R1148 VTAIL.n262 VTAIL.n225 171.744
R1149 VTAIL.n262 VTAIL.n261 171.744
R1150 VTAIL.n261 VTAIL.n260 171.744
R1151 VTAIL.n260 VTAIL.n229 171.744
R1152 VTAIL.n253 VTAIL.n229 171.744
R1153 VTAIL.n253 VTAIL.n252 171.744
R1154 VTAIL.n252 VTAIL.n234 171.744
R1155 VTAIL.n245 VTAIL.n234 171.744
R1156 VTAIL.n245 VTAIL.n244 171.744
R1157 VTAIL.n244 VTAIL.n238 171.744
R1158 VTAIL.n214 VTAIL.n213 171.744
R1159 VTAIL.n213 VTAIL.n169 171.744
R1160 VTAIL.n206 VTAIL.n169 171.744
R1161 VTAIL.n206 VTAIL.n205 171.744
R1162 VTAIL.n205 VTAIL.n204 171.744
R1163 VTAIL.n204 VTAIL.n173 171.744
R1164 VTAIL.n197 VTAIL.n173 171.744
R1165 VTAIL.n197 VTAIL.n196 171.744
R1166 VTAIL.n196 VTAIL.n178 171.744
R1167 VTAIL.n189 VTAIL.n178 171.744
R1168 VTAIL.n189 VTAIL.n188 171.744
R1169 VTAIL.n188 VTAIL.n182 171.744
R1170 VTAIL.t4 VTAIL.n401 85.8723
R1171 VTAIL.t1 VTAIL.n17 85.8723
R1172 VTAIL.t13 VTAIL.n71 85.8723
R1173 VTAIL.t10 VTAIL.n127 85.8723
R1174 VTAIL.t9 VTAIL.n348 85.8723
R1175 VTAIL.t15 VTAIL.n292 85.8723
R1176 VTAIL.t2 VTAIL.n238 85.8723
R1177 VTAIL.t7 VTAIL.n182 85.8723
R1178 VTAIL.n331 VTAIL.n330 58.6947
R1179 VTAIL.n221 VTAIL.n220 58.6947
R1180 VTAIL.n1 VTAIL.n0 58.6945
R1181 VTAIL.n111 VTAIL.n110 58.6945
R1182 VTAIL.n439 VTAIL.n438 30.4399
R1183 VTAIL.n55 VTAIL.n54 30.4399
R1184 VTAIL.n109 VTAIL.n108 30.4399
R1185 VTAIL.n165 VTAIL.n164 30.4399
R1186 VTAIL.n385 VTAIL.n384 30.4399
R1187 VTAIL.n329 VTAIL.n328 30.4399
R1188 VTAIL.n275 VTAIL.n274 30.4399
R1189 VTAIL.n219 VTAIL.n218 30.4399
R1190 VTAIL.n439 VTAIL.n385 22.2289
R1191 VTAIL.n219 VTAIL.n165 22.2289
R1192 VTAIL.n427 VTAIL.n392 13.1884
R1193 VTAIL.n43 VTAIL.n8 13.1884
R1194 VTAIL.n97 VTAIL.n62 13.1884
R1195 VTAIL.n153 VTAIL.n118 13.1884
R1196 VTAIL.n373 VTAIL.n338 13.1884
R1197 VTAIL.n317 VTAIL.n282 13.1884
R1198 VTAIL.n263 VTAIL.n228 13.1884
R1199 VTAIL.n207 VTAIL.n172 13.1884
R1200 VTAIL.n423 VTAIL.n422 12.8005
R1201 VTAIL.n428 VTAIL.n390 12.8005
R1202 VTAIL.n39 VTAIL.n38 12.8005
R1203 VTAIL.n44 VTAIL.n6 12.8005
R1204 VTAIL.n93 VTAIL.n92 12.8005
R1205 VTAIL.n98 VTAIL.n60 12.8005
R1206 VTAIL.n149 VTAIL.n148 12.8005
R1207 VTAIL.n154 VTAIL.n116 12.8005
R1208 VTAIL.n374 VTAIL.n336 12.8005
R1209 VTAIL.n369 VTAIL.n340 12.8005
R1210 VTAIL.n318 VTAIL.n280 12.8005
R1211 VTAIL.n313 VTAIL.n284 12.8005
R1212 VTAIL.n264 VTAIL.n226 12.8005
R1213 VTAIL.n259 VTAIL.n230 12.8005
R1214 VTAIL.n208 VTAIL.n170 12.8005
R1215 VTAIL.n203 VTAIL.n174 12.8005
R1216 VTAIL.n421 VTAIL.n394 12.0247
R1217 VTAIL.n432 VTAIL.n431 12.0247
R1218 VTAIL.n37 VTAIL.n10 12.0247
R1219 VTAIL.n48 VTAIL.n47 12.0247
R1220 VTAIL.n91 VTAIL.n64 12.0247
R1221 VTAIL.n102 VTAIL.n101 12.0247
R1222 VTAIL.n147 VTAIL.n120 12.0247
R1223 VTAIL.n158 VTAIL.n157 12.0247
R1224 VTAIL.n378 VTAIL.n377 12.0247
R1225 VTAIL.n368 VTAIL.n341 12.0247
R1226 VTAIL.n322 VTAIL.n321 12.0247
R1227 VTAIL.n312 VTAIL.n285 12.0247
R1228 VTAIL.n268 VTAIL.n267 12.0247
R1229 VTAIL.n258 VTAIL.n231 12.0247
R1230 VTAIL.n212 VTAIL.n211 12.0247
R1231 VTAIL.n202 VTAIL.n175 12.0247
R1232 VTAIL.n418 VTAIL.n417 11.249
R1233 VTAIL.n435 VTAIL.n388 11.249
R1234 VTAIL.n34 VTAIL.n33 11.249
R1235 VTAIL.n51 VTAIL.n4 11.249
R1236 VTAIL.n88 VTAIL.n87 11.249
R1237 VTAIL.n105 VTAIL.n58 11.249
R1238 VTAIL.n144 VTAIL.n143 11.249
R1239 VTAIL.n161 VTAIL.n114 11.249
R1240 VTAIL.n381 VTAIL.n334 11.249
R1241 VTAIL.n365 VTAIL.n364 11.249
R1242 VTAIL.n325 VTAIL.n278 11.249
R1243 VTAIL.n309 VTAIL.n308 11.249
R1244 VTAIL.n271 VTAIL.n224 11.249
R1245 VTAIL.n255 VTAIL.n254 11.249
R1246 VTAIL.n215 VTAIL.n168 11.249
R1247 VTAIL.n199 VTAIL.n198 11.249
R1248 VTAIL.n403 VTAIL.n402 10.7239
R1249 VTAIL.n19 VTAIL.n18 10.7239
R1250 VTAIL.n73 VTAIL.n72 10.7239
R1251 VTAIL.n129 VTAIL.n128 10.7239
R1252 VTAIL.n350 VTAIL.n349 10.7239
R1253 VTAIL.n294 VTAIL.n293 10.7239
R1254 VTAIL.n240 VTAIL.n239 10.7239
R1255 VTAIL.n184 VTAIL.n183 10.7239
R1256 VTAIL.n414 VTAIL.n396 10.4732
R1257 VTAIL.n436 VTAIL.n386 10.4732
R1258 VTAIL.n30 VTAIL.n12 10.4732
R1259 VTAIL.n52 VTAIL.n2 10.4732
R1260 VTAIL.n84 VTAIL.n66 10.4732
R1261 VTAIL.n106 VTAIL.n56 10.4732
R1262 VTAIL.n140 VTAIL.n122 10.4732
R1263 VTAIL.n162 VTAIL.n112 10.4732
R1264 VTAIL.n382 VTAIL.n332 10.4732
R1265 VTAIL.n361 VTAIL.n343 10.4732
R1266 VTAIL.n326 VTAIL.n276 10.4732
R1267 VTAIL.n305 VTAIL.n287 10.4732
R1268 VTAIL.n272 VTAIL.n222 10.4732
R1269 VTAIL.n251 VTAIL.n233 10.4732
R1270 VTAIL.n216 VTAIL.n166 10.4732
R1271 VTAIL.n195 VTAIL.n177 10.4732
R1272 VTAIL.n413 VTAIL.n398 9.69747
R1273 VTAIL.n29 VTAIL.n14 9.69747
R1274 VTAIL.n83 VTAIL.n68 9.69747
R1275 VTAIL.n139 VTAIL.n124 9.69747
R1276 VTAIL.n360 VTAIL.n345 9.69747
R1277 VTAIL.n304 VTAIL.n289 9.69747
R1278 VTAIL.n250 VTAIL.n235 9.69747
R1279 VTAIL.n194 VTAIL.n179 9.69747
R1280 VTAIL.n438 VTAIL.n437 9.45567
R1281 VTAIL.n54 VTAIL.n53 9.45567
R1282 VTAIL.n108 VTAIL.n107 9.45567
R1283 VTAIL.n164 VTAIL.n163 9.45567
R1284 VTAIL.n384 VTAIL.n383 9.45567
R1285 VTAIL.n328 VTAIL.n327 9.45567
R1286 VTAIL.n274 VTAIL.n273 9.45567
R1287 VTAIL.n218 VTAIL.n217 9.45567
R1288 VTAIL.n437 VTAIL.n436 9.3005
R1289 VTAIL.n388 VTAIL.n387 9.3005
R1290 VTAIL.n431 VTAIL.n430 9.3005
R1291 VTAIL.n429 VTAIL.n428 9.3005
R1292 VTAIL.n405 VTAIL.n404 9.3005
R1293 VTAIL.n400 VTAIL.n399 9.3005
R1294 VTAIL.n411 VTAIL.n410 9.3005
R1295 VTAIL.n413 VTAIL.n412 9.3005
R1296 VTAIL.n396 VTAIL.n395 9.3005
R1297 VTAIL.n419 VTAIL.n418 9.3005
R1298 VTAIL.n421 VTAIL.n420 9.3005
R1299 VTAIL.n422 VTAIL.n391 9.3005
R1300 VTAIL.n53 VTAIL.n52 9.3005
R1301 VTAIL.n4 VTAIL.n3 9.3005
R1302 VTAIL.n47 VTAIL.n46 9.3005
R1303 VTAIL.n45 VTAIL.n44 9.3005
R1304 VTAIL.n21 VTAIL.n20 9.3005
R1305 VTAIL.n16 VTAIL.n15 9.3005
R1306 VTAIL.n27 VTAIL.n26 9.3005
R1307 VTAIL.n29 VTAIL.n28 9.3005
R1308 VTAIL.n12 VTAIL.n11 9.3005
R1309 VTAIL.n35 VTAIL.n34 9.3005
R1310 VTAIL.n37 VTAIL.n36 9.3005
R1311 VTAIL.n38 VTAIL.n7 9.3005
R1312 VTAIL.n107 VTAIL.n106 9.3005
R1313 VTAIL.n58 VTAIL.n57 9.3005
R1314 VTAIL.n101 VTAIL.n100 9.3005
R1315 VTAIL.n99 VTAIL.n98 9.3005
R1316 VTAIL.n75 VTAIL.n74 9.3005
R1317 VTAIL.n70 VTAIL.n69 9.3005
R1318 VTAIL.n81 VTAIL.n80 9.3005
R1319 VTAIL.n83 VTAIL.n82 9.3005
R1320 VTAIL.n66 VTAIL.n65 9.3005
R1321 VTAIL.n89 VTAIL.n88 9.3005
R1322 VTAIL.n91 VTAIL.n90 9.3005
R1323 VTAIL.n92 VTAIL.n61 9.3005
R1324 VTAIL.n163 VTAIL.n162 9.3005
R1325 VTAIL.n114 VTAIL.n113 9.3005
R1326 VTAIL.n157 VTAIL.n156 9.3005
R1327 VTAIL.n155 VTAIL.n154 9.3005
R1328 VTAIL.n131 VTAIL.n130 9.3005
R1329 VTAIL.n126 VTAIL.n125 9.3005
R1330 VTAIL.n137 VTAIL.n136 9.3005
R1331 VTAIL.n139 VTAIL.n138 9.3005
R1332 VTAIL.n122 VTAIL.n121 9.3005
R1333 VTAIL.n145 VTAIL.n144 9.3005
R1334 VTAIL.n147 VTAIL.n146 9.3005
R1335 VTAIL.n148 VTAIL.n117 9.3005
R1336 VTAIL.n352 VTAIL.n351 9.3005
R1337 VTAIL.n347 VTAIL.n346 9.3005
R1338 VTAIL.n358 VTAIL.n357 9.3005
R1339 VTAIL.n360 VTAIL.n359 9.3005
R1340 VTAIL.n343 VTAIL.n342 9.3005
R1341 VTAIL.n366 VTAIL.n365 9.3005
R1342 VTAIL.n368 VTAIL.n367 9.3005
R1343 VTAIL.n340 VTAIL.n337 9.3005
R1344 VTAIL.n383 VTAIL.n382 9.3005
R1345 VTAIL.n334 VTAIL.n333 9.3005
R1346 VTAIL.n377 VTAIL.n376 9.3005
R1347 VTAIL.n375 VTAIL.n374 9.3005
R1348 VTAIL.n296 VTAIL.n295 9.3005
R1349 VTAIL.n291 VTAIL.n290 9.3005
R1350 VTAIL.n302 VTAIL.n301 9.3005
R1351 VTAIL.n304 VTAIL.n303 9.3005
R1352 VTAIL.n287 VTAIL.n286 9.3005
R1353 VTAIL.n310 VTAIL.n309 9.3005
R1354 VTAIL.n312 VTAIL.n311 9.3005
R1355 VTAIL.n284 VTAIL.n281 9.3005
R1356 VTAIL.n327 VTAIL.n326 9.3005
R1357 VTAIL.n278 VTAIL.n277 9.3005
R1358 VTAIL.n321 VTAIL.n320 9.3005
R1359 VTAIL.n319 VTAIL.n318 9.3005
R1360 VTAIL.n242 VTAIL.n241 9.3005
R1361 VTAIL.n237 VTAIL.n236 9.3005
R1362 VTAIL.n248 VTAIL.n247 9.3005
R1363 VTAIL.n250 VTAIL.n249 9.3005
R1364 VTAIL.n233 VTAIL.n232 9.3005
R1365 VTAIL.n256 VTAIL.n255 9.3005
R1366 VTAIL.n258 VTAIL.n257 9.3005
R1367 VTAIL.n230 VTAIL.n227 9.3005
R1368 VTAIL.n273 VTAIL.n272 9.3005
R1369 VTAIL.n224 VTAIL.n223 9.3005
R1370 VTAIL.n267 VTAIL.n266 9.3005
R1371 VTAIL.n265 VTAIL.n264 9.3005
R1372 VTAIL.n186 VTAIL.n185 9.3005
R1373 VTAIL.n181 VTAIL.n180 9.3005
R1374 VTAIL.n192 VTAIL.n191 9.3005
R1375 VTAIL.n194 VTAIL.n193 9.3005
R1376 VTAIL.n177 VTAIL.n176 9.3005
R1377 VTAIL.n200 VTAIL.n199 9.3005
R1378 VTAIL.n202 VTAIL.n201 9.3005
R1379 VTAIL.n174 VTAIL.n171 9.3005
R1380 VTAIL.n217 VTAIL.n216 9.3005
R1381 VTAIL.n168 VTAIL.n167 9.3005
R1382 VTAIL.n211 VTAIL.n210 9.3005
R1383 VTAIL.n209 VTAIL.n208 9.3005
R1384 VTAIL.n410 VTAIL.n409 8.92171
R1385 VTAIL.n26 VTAIL.n25 8.92171
R1386 VTAIL.n80 VTAIL.n79 8.92171
R1387 VTAIL.n136 VTAIL.n135 8.92171
R1388 VTAIL.n357 VTAIL.n356 8.92171
R1389 VTAIL.n301 VTAIL.n300 8.92171
R1390 VTAIL.n247 VTAIL.n246 8.92171
R1391 VTAIL.n191 VTAIL.n190 8.92171
R1392 VTAIL.n406 VTAIL.n400 8.14595
R1393 VTAIL.n22 VTAIL.n16 8.14595
R1394 VTAIL.n76 VTAIL.n70 8.14595
R1395 VTAIL.n132 VTAIL.n126 8.14595
R1396 VTAIL.n353 VTAIL.n347 8.14595
R1397 VTAIL.n297 VTAIL.n291 8.14595
R1398 VTAIL.n243 VTAIL.n237 8.14595
R1399 VTAIL.n187 VTAIL.n181 8.14595
R1400 VTAIL.n405 VTAIL.n402 7.3702
R1401 VTAIL.n21 VTAIL.n18 7.3702
R1402 VTAIL.n75 VTAIL.n72 7.3702
R1403 VTAIL.n131 VTAIL.n128 7.3702
R1404 VTAIL.n352 VTAIL.n349 7.3702
R1405 VTAIL.n296 VTAIL.n293 7.3702
R1406 VTAIL.n242 VTAIL.n239 7.3702
R1407 VTAIL.n186 VTAIL.n183 7.3702
R1408 VTAIL.n406 VTAIL.n405 5.81868
R1409 VTAIL.n22 VTAIL.n21 5.81868
R1410 VTAIL.n76 VTAIL.n75 5.81868
R1411 VTAIL.n132 VTAIL.n131 5.81868
R1412 VTAIL.n353 VTAIL.n352 5.81868
R1413 VTAIL.n297 VTAIL.n296 5.81868
R1414 VTAIL.n243 VTAIL.n242 5.81868
R1415 VTAIL.n187 VTAIL.n186 5.81868
R1416 VTAIL.n409 VTAIL.n400 5.04292
R1417 VTAIL.n25 VTAIL.n16 5.04292
R1418 VTAIL.n79 VTAIL.n70 5.04292
R1419 VTAIL.n135 VTAIL.n126 5.04292
R1420 VTAIL.n356 VTAIL.n347 5.04292
R1421 VTAIL.n300 VTAIL.n291 5.04292
R1422 VTAIL.n246 VTAIL.n237 5.04292
R1423 VTAIL.n190 VTAIL.n181 5.04292
R1424 VTAIL.n410 VTAIL.n398 4.26717
R1425 VTAIL.n26 VTAIL.n14 4.26717
R1426 VTAIL.n80 VTAIL.n68 4.26717
R1427 VTAIL.n136 VTAIL.n124 4.26717
R1428 VTAIL.n357 VTAIL.n345 4.26717
R1429 VTAIL.n301 VTAIL.n289 4.26717
R1430 VTAIL.n247 VTAIL.n235 4.26717
R1431 VTAIL.n191 VTAIL.n179 4.26717
R1432 VTAIL.n414 VTAIL.n413 3.49141
R1433 VTAIL.n438 VTAIL.n386 3.49141
R1434 VTAIL.n30 VTAIL.n29 3.49141
R1435 VTAIL.n54 VTAIL.n2 3.49141
R1436 VTAIL.n84 VTAIL.n83 3.49141
R1437 VTAIL.n108 VTAIL.n56 3.49141
R1438 VTAIL.n140 VTAIL.n139 3.49141
R1439 VTAIL.n164 VTAIL.n112 3.49141
R1440 VTAIL.n384 VTAIL.n332 3.49141
R1441 VTAIL.n361 VTAIL.n360 3.49141
R1442 VTAIL.n328 VTAIL.n276 3.49141
R1443 VTAIL.n305 VTAIL.n304 3.49141
R1444 VTAIL.n274 VTAIL.n222 3.49141
R1445 VTAIL.n251 VTAIL.n250 3.49141
R1446 VTAIL.n218 VTAIL.n166 3.49141
R1447 VTAIL.n195 VTAIL.n194 3.49141
R1448 VTAIL.n0 VTAIL.t5 3.29381
R1449 VTAIL.n0 VTAIL.t0 3.29381
R1450 VTAIL.n110 VTAIL.t11 3.29381
R1451 VTAIL.n110 VTAIL.t12 3.29381
R1452 VTAIL.n330 VTAIL.t8 3.29381
R1453 VTAIL.n330 VTAIL.t14 3.29381
R1454 VTAIL.n220 VTAIL.t6 3.29381
R1455 VTAIL.n220 VTAIL.t3 3.29381
R1456 VTAIL.n417 VTAIL.n396 2.71565
R1457 VTAIL.n436 VTAIL.n435 2.71565
R1458 VTAIL.n33 VTAIL.n12 2.71565
R1459 VTAIL.n52 VTAIL.n51 2.71565
R1460 VTAIL.n87 VTAIL.n66 2.71565
R1461 VTAIL.n106 VTAIL.n105 2.71565
R1462 VTAIL.n143 VTAIL.n122 2.71565
R1463 VTAIL.n162 VTAIL.n161 2.71565
R1464 VTAIL.n382 VTAIL.n381 2.71565
R1465 VTAIL.n364 VTAIL.n343 2.71565
R1466 VTAIL.n326 VTAIL.n325 2.71565
R1467 VTAIL.n308 VTAIL.n287 2.71565
R1468 VTAIL.n272 VTAIL.n271 2.71565
R1469 VTAIL.n254 VTAIL.n233 2.71565
R1470 VTAIL.n216 VTAIL.n215 2.71565
R1471 VTAIL.n198 VTAIL.n177 2.71565
R1472 VTAIL.n404 VTAIL.n403 2.41283
R1473 VTAIL.n20 VTAIL.n19 2.41283
R1474 VTAIL.n74 VTAIL.n73 2.41283
R1475 VTAIL.n130 VTAIL.n129 2.41283
R1476 VTAIL.n351 VTAIL.n350 2.41283
R1477 VTAIL.n295 VTAIL.n294 2.41283
R1478 VTAIL.n241 VTAIL.n240 2.41283
R1479 VTAIL.n185 VTAIL.n184 2.41283
R1480 VTAIL.n418 VTAIL.n394 1.93989
R1481 VTAIL.n432 VTAIL.n388 1.93989
R1482 VTAIL.n34 VTAIL.n10 1.93989
R1483 VTAIL.n48 VTAIL.n4 1.93989
R1484 VTAIL.n88 VTAIL.n64 1.93989
R1485 VTAIL.n102 VTAIL.n58 1.93989
R1486 VTAIL.n144 VTAIL.n120 1.93989
R1487 VTAIL.n158 VTAIL.n114 1.93989
R1488 VTAIL.n378 VTAIL.n334 1.93989
R1489 VTAIL.n365 VTAIL.n341 1.93989
R1490 VTAIL.n322 VTAIL.n278 1.93989
R1491 VTAIL.n309 VTAIL.n285 1.93989
R1492 VTAIL.n268 VTAIL.n224 1.93989
R1493 VTAIL.n255 VTAIL.n231 1.93989
R1494 VTAIL.n212 VTAIL.n168 1.93989
R1495 VTAIL.n199 VTAIL.n175 1.93989
R1496 VTAIL.n221 VTAIL.n219 1.35395
R1497 VTAIL.n275 VTAIL.n221 1.35395
R1498 VTAIL.n331 VTAIL.n329 1.35395
R1499 VTAIL.n385 VTAIL.n331 1.35395
R1500 VTAIL.n165 VTAIL.n111 1.35395
R1501 VTAIL.n111 VTAIL.n109 1.35395
R1502 VTAIL.n55 VTAIL.n1 1.35395
R1503 VTAIL VTAIL.n439 1.29576
R1504 VTAIL.n423 VTAIL.n421 1.16414
R1505 VTAIL.n431 VTAIL.n390 1.16414
R1506 VTAIL.n39 VTAIL.n37 1.16414
R1507 VTAIL.n47 VTAIL.n6 1.16414
R1508 VTAIL.n93 VTAIL.n91 1.16414
R1509 VTAIL.n101 VTAIL.n60 1.16414
R1510 VTAIL.n149 VTAIL.n147 1.16414
R1511 VTAIL.n157 VTAIL.n116 1.16414
R1512 VTAIL.n377 VTAIL.n336 1.16414
R1513 VTAIL.n369 VTAIL.n368 1.16414
R1514 VTAIL.n321 VTAIL.n280 1.16414
R1515 VTAIL.n313 VTAIL.n312 1.16414
R1516 VTAIL.n267 VTAIL.n226 1.16414
R1517 VTAIL.n259 VTAIL.n258 1.16414
R1518 VTAIL.n211 VTAIL.n170 1.16414
R1519 VTAIL.n203 VTAIL.n202 1.16414
R1520 VTAIL.n329 VTAIL.n275 0.470328
R1521 VTAIL.n109 VTAIL.n55 0.470328
R1522 VTAIL.n422 VTAIL.n392 0.388379
R1523 VTAIL.n428 VTAIL.n427 0.388379
R1524 VTAIL.n38 VTAIL.n8 0.388379
R1525 VTAIL.n44 VTAIL.n43 0.388379
R1526 VTAIL.n92 VTAIL.n62 0.388379
R1527 VTAIL.n98 VTAIL.n97 0.388379
R1528 VTAIL.n148 VTAIL.n118 0.388379
R1529 VTAIL.n154 VTAIL.n153 0.388379
R1530 VTAIL.n374 VTAIL.n373 0.388379
R1531 VTAIL.n340 VTAIL.n338 0.388379
R1532 VTAIL.n318 VTAIL.n317 0.388379
R1533 VTAIL.n284 VTAIL.n282 0.388379
R1534 VTAIL.n264 VTAIL.n263 0.388379
R1535 VTAIL.n230 VTAIL.n228 0.388379
R1536 VTAIL.n208 VTAIL.n207 0.388379
R1537 VTAIL.n174 VTAIL.n172 0.388379
R1538 VTAIL.n404 VTAIL.n399 0.155672
R1539 VTAIL.n411 VTAIL.n399 0.155672
R1540 VTAIL.n412 VTAIL.n411 0.155672
R1541 VTAIL.n412 VTAIL.n395 0.155672
R1542 VTAIL.n419 VTAIL.n395 0.155672
R1543 VTAIL.n420 VTAIL.n419 0.155672
R1544 VTAIL.n420 VTAIL.n391 0.155672
R1545 VTAIL.n429 VTAIL.n391 0.155672
R1546 VTAIL.n430 VTAIL.n429 0.155672
R1547 VTAIL.n430 VTAIL.n387 0.155672
R1548 VTAIL.n437 VTAIL.n387 0.155672
R1549 VTAIL.n20 VTAIL.n15 0.155672
R1550 VTAIL.n27 VTAIL.n15 0.155672
R1551 VTAIL.n28 VTAIL.n27 0.155672
R1552 VTAIL.n28 VTAIL.n11 0.155672
R1553 VTAIL.n35 VTAIL.n11 0.155672
R1554 VTAIL.n36 VTAIL.n35 0.155672
R1555 VTAIL.n36 VTAIL.n7 0.155672
R1556 VTAIL.n45 VTAIL.n7 0.155672
R1557 VTAIL.n46 VTAIL.n45 0.155672
R1558 VTAIL.n46 VTAIL.n3 0.155672
R1559 VTAIL.n53 VTAIL.n3 0.155672
R1560 VTAIL.n74 VTAIL.n69 0.155672
R1561 VTAIL.n81 VTAIL.n69 0.155672
R1562 VTAIL.n82 VTAIL.n81 0.155672
R1563 VTAIL.n82 VTAIL.n65 0.155672
R1564 VTAIL.n89 VTAIL.n65 0.155672
R1565 VTAIL.n90 VTAIL.n89 0.155672
R1566 VTAIL.n90 VTAIL.n61 0.155672
R1567 VTAIL.n99 VTAIL.n61 0.155672
R1568 VTAIL.n100 VTAIL.n99 0.155672
R1569 VTAIL.n100 VTAIL.n57 0.155672
R1570 VTAIL.n107 VTAIL.n57 0.155672
R1571 VTAIL.n130 VTAIL.n125 0.155672
R1572 VTAIL.n137 VTAIL.n125 0.155672
R1573 VTAIL.n138 VTAIL.n137 0.155672
R1574 VTAIL.n138 VTAIL.n121 0.155672
R1575 VTAIL.n145 VTAIL.n121 0.155672
R1576 VTAIL.n146 VTAIL.n145 0.155672
R1577 VTAIL.n146 VTAIL.n117 0.155672
R1578 VTAIL.n155 VTAIL.n117 0.155672
R1579 VTAIL.n156 VTAIL.n155 0.155672
R1580 VTAIL.n156 VTAIL.n113 0.155672
R1581 VTAIL.n163 VTAIL.n113 0.155672
R1582 VTAIL.n383 VTAIL.n333 0.155672
R1583 VTAIL.n376 VTAIL.n333 0.155672
R1584 VTAIL.n376 VTAIL.n375 0.155672
R1585 VTAIL.n375 VTAIL.n337 0.155672
R1586 VTAIL.n367 VTAIL.n337 0.155672
R1587 VTAIL.n367 VTAIL.n366 0.155672
R1588 VTAIL.n366 VTAIL.n342 0.155672
R1589 VTAIL.n359 VTAIL.n342 0.155672
R1590 VTAIL.n359 VTAIL.n358 0.155672
R1591 VTAIL.n358 VTAIL.n346 0.155672
R1592 VTAIL.n351 VTAIL.n346 0.155672
R1593 VTAIL.n327 VTAIL.n277 0.155672
R1594 VTAIL.n320 VTAIL.n277 0.155672
R1595 VTAIL.n320 VTAIL.n319 0.155672
R1596 VTAIL.n319 VTAIL.n281 0.155672
R1597 VTAIL.n311 VTAIL.n281 0.155672
R1598 VTAIL.n311 VTAIL.n310 0.155672
R1599 VTAIL.n310 VTAIL.n286 0.155672
R1600 VTAIL.n303 VTAIL.n286 0.155672
R1601 VTAIL.n303 VTAIL.n302 0.155672
R1602 VTAIL.n302 VTAIL.n290 0.155672
R1603 VTAIL.n295 VTAIL.n290 0.155672
R1604 VTAIL.n273 VTAIL.n223 0.155672
R1605 VTAIL.n266 VTAIL.n223 0.155672
R1606 VTAIL.n266 VTAIL.n265 0.155672
R1607 VTAIL.n265 VTAIL.n227 0.155672
R1608 VTAIL.n257 VTAIL.n227 0.155672
R1609 VTAIL.n257 VTAIL.n256 0.155672
R1610 VTAIL.n256 VTAIL.n232 0.155672
R1611 VTAIL.n249 VTAIL.n232 0.155672
R1612 VTAIL.n249 VTAIL.n248 0.155672
R1613 VTAIL.n248 VTAIL.n236 0.155672
R1614 VTAIL.n241 VTAIL.n236 0.155672
R1615 VTAIL.n217 VTAIL.n167 0.155672
R1616 VTAIL.n210 VTAIL.n167 0.155672
R1617 VTAIL.n210 VTAIL.n209 0.155672
R1618 VTAIL.n209 VTAIL.n171 0.155672
R1619 VTAIL.n201 VTAIL.n171 0.155672
R1620 VTAIL.n201 VTAIL.n200 0.155672
R1621 VTAIL.n200 VTAIL.n176 0.155672
R1622 VTAIL.n193 VTAIL.n176 0.155672
R1623 VTAIL.n193 VTAIL.n192 0.155672
R1624 VTAIL.n192 VTAIL.n180 0.155672
R1625 VTAIL.n185 VTAIL.n180 0.155672
R1626 VTAIL VTAIL.n1 0.0586897
R1627 VN.n4 VN.t1 243.444
R1628 VN.n19 VN.t2 243.444
R1629 VN.n13 VN.t6 223.702
R1630 VN.n28 VN.t0 223.702
R1631 VN.n3 VN.t4 191.828
R1632 VN.n1 VN.t5 191.828
R1633 VN.n18 VN.t7 191.828
R1634 VN.n16 VN.t3 191.828
R1635 VN.n27 VN.n15 161.3
R1636 VN.n26 VN.n25 161.3
R1637 VN.n24 VN.n23 161.3
R1638 VN.n22 VN.n17 161.3
R1639 VN.n21 VN.n20 161.3
R1640 VN.n12 VN.n0 161.3
R1641 VN.n11 VN.n10 161.3
R1642 VN.n9 VN.n8 161.3
R1643 VN.n7 VN.n2 161.3
R1644 VN.n6 VN.n5 161.3
R1645 VN.n29 VN.n28 80.6037
R1646 VN.n14 VN.n13 80.6037
R1647 VN.n4 VN.n3 43.5433
R1648 VN.n19 VN.n18 43.5433
R1649 VN VN.n29 43.3703
R1650 VN.n7 VN.n6 40.4934
R1651 VN.n8 VN.n7 40.4934
R1652 VN.n22 VN.n21 40.4934
R1653 VN.n23 VN.n22 40.4934
R1654 VN.n13 VN.n12 34.3247
R1655 VN.n28 VN.n27 34.3247
R1656 VN.n12 VN.n11 33.6945
R1657 VN.n27 VN.n26 33.6945
R1658 VN.n20 VN.n19 29.3131
R1659 VN.n5 VN.n4 29.3131
R1660 VN.n6 VN.n3 13.9467
R1661 VN.n8 VN.n1 13.9467
R1662 VN.n21 VN.n18 13.9467
R1663 VN.n23 VN.n16 13.9467
R1664 VN.n11 VN.n1 10.5213
R1665 VN.n26 VN.n16 10.5213
R1666 VN.n29 VN.n15 0.285035
R1667 VN.n14 VN.n0 0.285035
R1668 VN.n25 VN.n15 0.189894
R1669 VN.n25 VN.n24 0.189894
R1670 VN.n24 VN.n17 0.189894
R1671 VN.n20 VN.n17 0.189894
R1672 VN.n5 VN.n2 0.189894
R1673 VN.n9 VN.n2 0.189894
R1674 VN.n10 VN.n9 0.189894
R1675 VN.n10 VN.n0 0.189894
R1676 VN VN.n14 0.146778
R1677 VDD2.n2 VDD2.n1 75.9947
R1678 VDD2.n2 VDD2.n0 75.9947
R1679 VDD2 VDD2.n5 75.9919
R1680 VDD2.n4 VDD2.n3 75.3735
R1681 VDD2.n4 VDD2.n2 38.3144
R1682 VDD2.n5 VDD2.t0 3.29381
R1683 VDD2.n5 VDD2.t5 3.29381
R1684 VDD2.n3 VDD2.t7 3.29381
R1685 VDD2.n3 VDD2.t4 3.29381
R1686 VDD2.n1 VDD2.t2 3.29381
R1687 VDD2.n1 VDD2.t1 3.29381
R1688 VDD2.n0 VDD2.t6 3.29381
R1689 VDD2.n0 VDD2.t3 3.29381
R1690 VDD2 VDD2.n4 0.735414
C0 w_n2540_n2942# VP 5.07712f
C1 VN w_n2540_n2942# 4.75138f
C2 B VDD1 1.17768f
C3 B VP 1.42203f
C4 VN B 0.883237f
C5 VP VDD1 6.13172f
C6 VN VDD1 0.148976f
C7 VN VP 5.60373f
C8 VDD2 VTAIL 7.83996f
C9 VTAIL w_n2540_n2942# 3.64003f
C10 VDD2 w_n2540_n2942# 1.49655f
C11 VTAIL B 3.61478f
C12 VDD2 B 1.23108f
C13 VTAIL VDD1 7.79467f
C14 VDD2 VDD1 1.09481f
C15 VTAIL VP 5.9614f
C16 VTAIL VN 5.9473f
C17 VDD2 VP 0.374659f
C18 VDD2 VN 5.90674f
C19 B w_n2540_n2942# 7.43608f
C20 w_n2540_n2942# VDD1 1.43901f
C21 VDD2 VSUBS 1.364389f
C22 VDD1 VSUBS 1.769464f
C23 VTAIL VSUBS 0.965238f
C24 VN VSUBS 5.02754f
C25 VP VSUBS 2.13127f
C26 B VSUBS 3.306795f
C27 w_n2540_n2942# VSUBS 92.3239f
C28 VDD2.t6 VSUBS 0.196813f
C29 VDD2.t3 VSUBS 0.196813f
C30 VDD2.n0 VSUBS 1.48187f
C31 VDD2.t2 VSUBS 0.196813f
C32 VDD2.t1 VSUBS 0.196813f
C33 VDD2.n1 VSUBS 1.48187f
C34 VDD2.n2 VSUBS 2.88106f
C35 VDD2.t7 VSUBS 0.196813f
C36 VDD2.t4 VSUBS 0.196813f
C37 VDD2.n3 VSUBS 1.47671f
C38 VDD2.n4 VSUBS 2.58651f
C39 VDD2.t0 VSUBS 0.196813f
C40 VDD2.t5 VSUBS 0.196813f
C41 VDD2.n5 VSUBS 1.48184f
C42 VN.n0 VSUBS 0.058737f
C43 VN.t5 VSUBS 1.45878f
C44 VN.n1 VSUBS 0.543757f
C45 VN.n2 VSUBS 0.044018f
C46 VN.t4 VSUBS 1.45878f
C47 VN.n3 VSUBS 0.602383f
C48 VN.t1 VSUBS 1.59423f
C49 VN.n4 VSUBS 0.61724f
C50 VN.n5 VSUBS 0.230216f
C51 VN.n6 VSUBS 0.070067f
C52 VN.n7 VSUBS 0.035585f
C53 VN.n8 VSUBS 0.070067f
C54 VN.n9 VSUBS 0.044018f
C55 VN.n10 VSUBS 0.044018f
C56 VN.n11 VSUBS 0.065824f
C57 VN.n12 VSUBS 0.030801f
C58 VN.t6 VSUBS 1.54241f
C59 VN.n13 VSUBS 0.628975f
C60 VN.n14 VSUBS 0.041225f
C61 VN.n15 VSUBS 0.058737f
C62 VN.t3 VSUBS 1.45878f
C63 VN.n16 VSUBS 0.543757f
C64 VN.n17 VSUBS 0.044018f
C65 VN.t7 VSUBS 1.45878f
C66 VN.n18 VSUBS 0.602383f
C67 VN.t2 VSUBS 1.59423f
C68 VN.n19 VSUBS 0.61724f
C69 VN.n20 VSUBS 0.230216f
C70 VN.n21 VSUBS 0.070067f
C71 VN.n22 VSUBS 0.035585f
C72 VN.n23 VSUBS 0.070067f
C73 VN.n24 VSUBS 0.044018f
C74 VN.n25 VSUBS 0.044018f
C75 VN.n26 VSUBS 0.065824f
C76 VN.n27 VSUBS 0.030801f
C77 VN.t0 VSUBS 1.54241f
C78 VN.n28 VSUBS 0.628975f
C79 VN.n29 VSUBS 1.93538f
C80 VTAIL.t5 VSUBS 0.194061f
C81 VTAIL.t0 VSUBS 0.194061f
C82 VTAIL.n0 VSUBS 1.32845f
C83 VTAIL.n1 VSUBS 0.660728f
C84 VTAIL.n2 VSUBS 0.02502f
C85 VTAIL.n3 VSUBS 0.024881f
C86 VTAIL.n4 VSUBS 0.01337f
C87 VTAIL.n5 VSUBS 0.031602f
C88 VTAIL.n6 VSUBS 0.014156f
C89 VTAIL.n7 VSUBS 0.024881f
C90 VTAIL.n8 VSUBS 0.013763f
C91 VTAIL.n9 VSUBS 0.031602f
C92 VTAIL.n10 VSUBS 0.014156f
C93 VTAIL.n11 VSUBS 0.024881f
C94 VTAIL.n12 VSUBS 0.01337f
C95 VTAIL.n13 VSUBS 0.031602f
C96 VTAIL.n14 VSUBS 0.014156f
C97 VTAIL.n15 VSUBS 0.024881f
C98 VTAIL.n16 VSUBS 0.01337f
C99 VTAIL.n17 VSUBS 0.023701f
C100 VTAIL.n18 VSUBS 0.023772f
C101 VTAIL.t1 VSUBS 0.06793f
C102 VTAIL.n19 VSUBS 0.171999f
C103 VTAIL.n20 VSUBS 0.990248f
C104 VTAIL.n21 VSUBS 0.01337f
C105 VTAIL.n22 VSUBS 0.014156f
C106 VTAIL.n23 VSUBS 0.031602f
C107 VTAIL.n24 VSUBS 0.031602f
C108 VTAIL.n25 VSUBS 0.014156f
C109 VTAIL.n26 VSUBS 0.01337f
C110 VTAIL.n27 VSUBS 0.024881f
C111 VTAIL.n28 VSUBS 0.024881f
C112 VTAIL.n29 VSUBS 0.01337f
C113 VTAIL.n30 VSUBS 0.014156f
C114 VTAIL.n31 VSUBS 0.031602f
C115 VTAIL.n32 VSUBS 0.031602f
C116 VTAIL.n33 VSUBS 0.014156f
C117 VTAIL.n34 VSUBS 0.01337f
C118 VTAIL.n35 VSUBS 0.024881f
C119 VTAIL.n36 VSUBS 0.024881f
C120 VTAIL.n37 VSUBS 0.01337f
C121 VTAIL.n38 VSUBS 0.01337f
C122 VTAIL.n39 VSUBS 0.014156f
C123 VTAIL.n40 VSUBS 0.031602f
C124 VTAIL.n41 VSUBS 0.031602f
C125 VTAIL.n42 VSUBS 0.031602f
C126 VTAIL.n43 VSUBS 0.013763f
C127 VTAIL.n44 VSUBS 0.01337f
C128 VTAIL.n45 VSUBS 0.024881f
C129 VTAIL.n46 VSUBS 0.024881f
C130 VTAIL.n47 VSUBS 0.01337f
C131 VTAIL.n48 VSUBS 0.014156f
C132 VTAIL.n49 VSUBS 0.031602f
C133 VTAIL.n50 VSUBS 0.068605f
C134 VTAIL.n51 VSUBS 0.014156f
C135 VTAIL.n52 VSUBS 0.01337f
C136 VTAIL.n53 VSUBS 0.054452f
C137 VTAIL.n54 VSUBS 0.034054f
C138 VTAIL.n55 VSUBS 0.165702f
C139 VTAIL.n56 VSUBS 0.02502f
C140 VTAIL.n57 VSUBS 0.024881f
C141 VTAIL.n58 VSUBS 0.01337f
C142 VTAIL.n59 VSUBS 0.031602f
C143 VTAIL.n60 VSUBS 0.014156f
C144 VTAIL.n61 VSUBS 0.024881f
C145 VTAIL.n62 VSUBS 0.013763f
C146 VTAIL.n63 VSUBS 0.031602f
C147 VTAIL.n64 VSUBS 0.014156f
C148 VTAIL.n65 VSUBS 0.024881f
C149 VTAIL.n66 VSUBS 0.01337f
C150 VTAIL.n67 VSUBS 0.031602f
C151 VTAIL.n68 VSUBS 0.014156f
C152 VTAIL.n69 VSUBS 0.024881f
C153 VTAIL.n70 VSUBS 0.01337f
C154 VTAIL.n71 VSUBS 0.023701f
C155 VTAIL.n72 VSUBS 0.023772f
C156 VTAIL.t13 VSUBS 0.06793f
C157 VTAIL.n73 VSUBS 0.171999f
C158 VTAIL.n74 VSUBS 0.990248f
C159 VTAIL.n75 VSUBS 0.01337f
C160 VTAIL.n76 VSUBS 0.014156f
C161 VTAIL.n77 VSUBS 0.031602f
C162 VTAIL.n78 VSUBS 0.031602f
C163 VTAIL.n79 VSUBS 0.014156f
C164 VTAIL.n80 VSUBS 0.01337f
C165 VTAIL.n81 VSUBS 0.024881f
C166 VTAIL.n82 VSUBS 0.024881f
C167 VTAIL.n83 VSUBS 0.01337f
C168 VTAIL.n84 VSUBS 0.014156f
C169 VTAIL.n85 VSUBS 0.031602f
C170 VTAIL.n86 VSUBS 0.031602f
C171 VTAIL.n87 VSUBS 0.014156f
C172 VTAIL.n88 VSUBS 0.01337f
C173 VTAIL.n89 VSUBS 0.024881f
C174 VTAIL.n90 VSUBS 0.024881f
C175 VTAIL.n91 VSUBS 0.01337f
C176 VTAIL.n92 VSUBS 0.01337f
C177 VTAIL.n93 VSUBS 0.014156f
C178 VTAIL.n94 VSUBS 0.031602f
C179 VTAIL.n95 VSUBS 0.031602f
C180 VTAIL.n96 VSUBS 0.031602f
C181 VTAIL.n97 VSUBS 0.013763f
C182 VTAIL.n98 VSUBS 0.01337f
C183 VTAIL.n99 VSUBS 0.024881f
C184 VTAIL.n100 VSUBS 0.024881f
C185 VTAIL.n101 VSUBS 0.01337f
C186 VTAIL.n102 VSUBS 0.014156f
C187 VTAIL.n103 VSUBS 0.031602f
C188 VTAIL.n104 VSUBS 0.068605f
C189 VTAIL.n105 VSUBS 0.014156f
C190 VTAIL.n106 VSUBS 0.01337f
C191 VTAIL.n107 VSUBS 0.054452f
C192 VTAIL.n108 VSUBS 0.034054f
C193 VTAIL.n109 VSUBS 0.165702f
C194 VTAIL.t11 VSUBS 0.194061f
C195 VTAIL.t12 VSUBS 0.194061f
C196 VTAIL.n110 VSUBS 1.32845f
C197 VTAIL.n111 VSUBS 0.764571f
C198 VTAIL.n112 VSUBS 0.02502f
C199 VTAIL.n113 VSUBS 0.024881f
C200 VTAIL.n114 VSUBS 0.01337f
C201 VTAIL.n115 VSUBS 0.031602f
C202 VTAIL.n116 VSUBS 0.014156f
C203 VTAIL.n117 VSUBS 0.024881f
C204 VTAIL.n118 VSUBS 0.013763f
C205 VTAIL.n119 VSUBS 0.031602f
C206 VTAIL.n120 VSUBS 0.014156f
C207 VTAIL.n121 VSUBS 0.024881f
C208 VTAIL.n122 VSUBS 0.01337f
C209 VTAIL.n123 VSUBS 0.031602f
C210 VTAIL.n124 VSUBS 0.014156f
C211 VTAIL.n125 VSUBS 0.024881f
C212 VTAIL.n126 VSUBS 0.01337f
C213 VTAIL.n127 VSUBS 0.023701f
C214 VTAIL.n128 VSUBS 0.023772f
C215 VTAIL.t10 VSUBS 0.06793f
C216 VTAIL.n129 VSUBS 0.171999f
C217 VTAIL.n130 VSUBS 0.990248f
C218 VTAIL.n131 VSUBS 0.01337f
C219 VTAIL.n132 VSUBS 0.014156f
C220 VTAIL.n133 VSUBS 0.031602f
C221 VTAIL.n134 VSUBS 0.031602f
C222 VTAIL.n135 VSUBS 0.014156f
C223 VTAIL.n136 VSUBS 0.01337f
C224 VTAIL.n137 VSUBS 0.024881f
C225 VTAIL.n138 VSUBS 0.024881f
C226 VTAIL.n139 VSUBS 0.01337f
C227 VTAIL.n140 VSUBS 0.014156f
C228 VTAIL.n141 VSUBS 0.031602f
C229 VTAIL.n142 VSUBS 0.031602f
C230 VTAIL.n143 VSUBS 0.014156f
C231 VTAIL.n144 VSUBS 0.01337f
C232 VTAIL.n145 VSUBS 0.024881f
C233 VTAIL.n146 VSUBS 0.024881f
C234 VTAIL.n147 VSUBS 0.01337f
C235 VTAIL.n148 VSUBS 0.01337f
C236 VTAIL.n149 VSUBS 0.014156f
C237 VTAIL.n150 VSUBS 0.031602f
C238 VTAIL.n151 VSUBS 0.031602f
C239 VTAIL.n152 VSUBS 0.031602f
C240 VTAIL.n153 VSUBS 0.013763f
C241 VTAIL.n154 VSUBS 0.01337f
C242 VTAIL.n155 VSUBS 0.024881f
C243 VTAIL.n156 VSUBS 0.024881f
C244 VTAIL.n157 VSUBS 0.01337f
C245 VTAIL.n158 VSUBS 0.014156f
C246 VTAIL.n159 VSUBS 0.031602f
C247 VTAIL.n160 VSUBS 0.068605f
C248 VTAIL.n161 VSUBS 0.014156f
C249 VTAIL.n162 VSUBS 0.01337f
C250 VTAIL.n163 VSUBS 0.054452f
C251 VTAIL.n164 VSUBS 0.034054f
C252 VTAIL.n165 VSUBS 1.25667f
C253 VTAIL.n166 VSUBS 0.02502f
C254 VTAIL.n167 VSUBS 0.024881f
C255 VTAIL.n168 VSUBS 0.01337f
C256 VTAIL.n169 VSUBS 0.031602f
C257 VTAIL.n170 VSUBS 0.014156f
C258 VTAIL.n171 VSUBS 0.024881f
C259 VTAIL.n172 VSUBS 0.013763f
C260 VTAIL.n173 VSUBS 0.031602f
C261 VTAIL.n174 VSUBS 0.01337f
C262 VTAIL.n175 VSUBS 0.014156f
C263 VTAIL.n176 VSUBS 0.024881f
C264 VTAIL.n177 VSUBS 0.01337f
C265 VTAIL.n178 VSUBS 0.031602f
C266 VTAIL.n179 VSUBS 0.014156f
C267 VTAIL.n180 VSUBS 0.024881f
C268 VTAIL.n181 VSUBS 0.01337f
C269 VTAIL.n182 VSUBS 0.023701f
C270 VTAIL.n183 VSUBS 0.023772f
C271 VTAIL.t7 VSUBS 0.06793f
C272 VTAIL.n184 VSUBS 0.171999f
C273 VTAIL.n185 VSUBS 0.990248f
C274 VTAIL.n186 VSUBS 0.01337f
C275 VTAIL.n187 VSUBS 0.014156f
C276 VTAIL.n188 VSUBS 0.031602f
C277 VTAIL.n189 VSUBS 0.031602f
C278 VTAIL.n190 VSUBS 0.014156f
C279 VTAIL.n191 VSUBS 0.01337f
C280 VTAIL.n192 VSUBS 0.024881f
C281 VTAIL.n193 VSUBS 0.024881f
C282 VTAIL.n194 VSUBS 0.01337f
C283 VTAIL.n195 VSUBS 0.014156f
C284 VTAIL.n196 VSUBS 0.031602f
C285 VTAIL.n197 VSUBS 0.031602f
C286 VTAIL.n198 VSUBS 0.014156f
C287 VTAIL.n199 VSUBS 0.01337f
C288 VTAIL.n200 VSUBS 0.024881f
C289 VTAIL.n201 VSUBS 0.024881f
C290 VTAIL.n202 VSUBS 0.01337f
C291 VTAIL.n203 VSUBS 0.014156f
C292 VTAIL.n204 VSUBS 0.031602f
C293 VTAIL.n205 VSUBS 0.031602f
C294 VTAIL.n206 VSUBS 0.031602f
C295 VTAIL.n207 VSUBS 0.013763f
C296 VTAIL.n208 VSUBS 0.01337f
C297 VTAIL.n209 VSUBS 0.024881f
C298 VTAIL.n210 VSUBS 0.024881f
C299 VTAIL.n211 VSUBS 0.01337f
C300 VTAIL.n212 VSUBS 0.014156f
C301 VTAIL.n213 VSUBS 0.031602f
C302 VTAIL.n214 VSUBS 0.068605f
C303 VTAIL.n215 VSUBS 0.014156f
C304 VTAIL.n216 VSUBS 0.01337f
C305 VTAIL.n217 VSUBS 0.054452f
C306 VTAIL.n218 VSUBS 0.034054f
C307 VTAIL.n219 VSUBS 1.25667f
C308 VTAIL.t6 VSUBS 0.194061f
C309 VTAIL.t3 VSUBS 0.194061f
C310 VTAIL.n220 VSUBS 1.32846f
C311 VTAIL.n221 VSUBS 0.764561f
C312 VTAIL.n222 VSUBS 0.02502f
C313 VTAIL.n223 VSUBS 0.024881f
C314 VTAIL.n224 VSUBS 0.01337f
C315 VTAIL.n225 VSUBS 0.031602f
C316 VTAIL.n226 VSUBS 0.014156f
C317 VTAIL.n227 VSUBS 0.024881f
C318 VTAIL.n228 VSUBS 0.013763f
C319 VTAIL.n229 VSUBS 0.031602f
C320 VTAIL.n230 VSUBS 0.01337f
C321 VTAIL.n231 VSUBS 0.014156f
C322 VTAIL.n232 VSUBS 0.024881f
C323 VTAIL.n233 VSUBS 0.01337f
C324 VTAIL.n234 VSUBS 0.031602f
C325 VTAIL.n235 VSUBS 0.014156f
C326 VTAIL.n236 VSUBS 0.024881f
C327 VTAIL.n237 VSUBS 0.01337f
C328 VTAIL.n238 VSUBS 0.023701f
C329 VTAIL.n239 VSUBS 0.023772f
C330 VTAIL.t2 VSUBS 0.06793f
C331 VTAIL.n240 VSUBS 0.171999f
C332 VTAIL.n241 VSUBS 0.990248f
C333 VTAIL.n242 VSUBS 0.01337f
C334 VTAIL.n243 VSUBS 0.014156f
C335 VTAIL.n244 VSUBS 0.031602f
C336 VTAIL.n245 VSUBS 0.031602f
C337 VTAIL.n246 VSUBS 0.014156f
C338 VTAIL.n247 VSUBS 0.01337f
C339 VTAIL.n248 VSUBS 0.024881f
C340 VTAIL.n249 VSUBS 0.024881f
C341 VTAIL.n250 VSUBS 0.01337f
C342 VTAIL.n251 VSUBS 0.014156f
C343 VTAIL.n252 VSUBS 0.031602f
C344 VTAIL.n253 VSUBS 0.031602f
C345 VTAIL.n254 VSUBS 0.014156f
C346 VTAIL.n255 VSUBS 0.01337f
C347 VTAIL.n256 VSUBS 0.024881f
C348 VTAIL.n257 VSUBS 0.024881f
C349 VTAIL.n258 VSUBS 0.01337f
C350 VTAIL.n259 VSUBS 0.014156f
C351 VTAIL.n260 VSUBS 0.031602f
C352 VTAIL.n261 VSUBS 0.031602f
C353 VTAIL.n262 VSUBS 0.031602f
C354 VTAIL.n263 VSUBS 0.013763f
C355 VTAIL.n264 VSUBS 0.01337f
C356 VTAIL.n265 VSUBS 0.024881f
C357 VTAIL.n266 VSUBS 0.024881f
C358 VTAIL.n267 VSUBS 0.01337f
C359 VTAIL.n268 VSUBS 0.014156f
C360 VTAIL.n269 VSUBS 0.031602f
C361 VTAIL.n270 VSUBS 0.068605f
C362 VTAIL.n271 VSUBS 0.014156f
C363 VTAIL.n272 VSUBS 0.01337f
C364 VTAIL.n273 VSUBS 0.054452f
C365 VTAIL.n274 VSUBS 0.034054f
C366 VTAIL.n275 VSUBS 0.165702f
C367 VTAIL.n276 VSUBS 0.02502f
C368 VTAIL.n277 VSUBS 0.024881f
C369 VTAIL.n278 VSUBS 0.01337f
C370 VTAIL.n279 VSUBS 0.031602f
C371 VTAIL.n280 VSUBS 0.014156f
C372 VTAIL.n281 VSUBS 0.024881f
C373 VTAIL.n282 VSUBS 0.013763f
C374 VTAIL.n283 VSUBS 0.031602f
C375 VTAIL.n284 VSUBS 0.01337f
C376 VTAIL.n285 VSUBS 0.014156f
C377 VTAIL.n286 VSUBS 0.024881f
C378 VTAIL.n287 VSUBS 0.01337f
C379 VTAIL.n288 VSUBS 0.031602f
C380 VTAIL.n289 VSUBS 0.014156f
C381 VTAIL.n290 VSUBS 0.024881f
C382 VTAIL.n291 VSUBS 0.01337f
C383 VTAIL.n292 VSUBS 0.023701f
C384 VTAIL.n293 VSUBS 0.023772f
C385 VTAIL.t15 VSUBS 0.06793f
C386 VTAIL.n294 VSUBS 0.171999f
C387 VTAIL.n295 VSUBS 0.990248f
C388 VTAIL.n296 VSUBS 0.01337f
C389 VTAIL.n297 VSUBS 0.014156f
C390 VTAIL.n298 VSUBS 0.031602f
C391 VTAIL.n299 VSUBS 0.031602f
C392 VTAIL.n300 VSUBS 0.014156f
C393 VTAIL.n301 VSUBS 0.01337f
C394 VTAIL.n302 VSUBS 0.024881f
C395 VTAIL.n303 VSUBS 0.024881f
C396 VTAIL.n304 VSUBS 0.01337f
C397 VTAIL.n305 VSUBS 0.014156f
C398 VTAIL.n306 VSUBS 0.031602f
C399 VTAIL.n307 VSUBS 0.031602f
C400 VTAIL.n308 VSUBS 0.014156f
C401 VTAIL.n309 VSUBS 0.01337f
C402 VTAIL.n310 VSUBS 0.024881f
C403 VTAIL.n311 VSUBS 0.024881f
C404 VTAIL.n312 VSUBS 0.01337f
C405 VTAIL.n313 VSUBS 0.014156f
C406 VTAIL.n314 VSUBS 0.031602f
C407 VTAIL.n315 VSUBS 0.031602f
C408 VTAIL.n316 VSUBS 0.031602f
C409 VTAIL.n317 VSUBS 0.013763f
C410 VTAIL.n318 VSUBS 0.01337f
C411 VTAIL.n319 VSUBS 0.024881f
C412 VTAIL.n320 VSUBS 0.024881f
C413 VTAIL.n321 VSUBS 0.01337f
C414 VTAIL.n322 VSUBS 0.014156f
C415 VTAIL.n323 VSUBS 0.031602f
C416 VTAIL.n324 VSUBS 0.068605f
C417 VTAIL.n325 VSUBS 0.014156f
C418 VTAIL.n326 VSUBS 0.01337f
C419 VTAIL.n327 VSUBS 0.054452f
C420 VTAIL.n328 VSUBS 0.034054f
C421 VTAIL.n329 VSUBS 0.165702f
C422 VTAIL.t8 VSUBS 0.194061f
C423 VTAIL.t14 VSUBS 0.194061f
C424 VTAIL.n330 VSUBS 1.32846f
C425 VTAIL.n331 VSUBS 0.764561f
C426 VTAIL.n332 VSUBS 0.02502f
C427 VTAIL.n333 VSUBS 0.024881f
C428 VTAIL.n334 VSUBS 0.01337f
C429 VTAIL.n335 VSUBS 0.031602f
C430 VTAIL.n336 VSUBS 0.014156f
C431 VTAIL.n337 VSUBS 0.024881f
C432 VTAIL.n338 VSUBS 0.013763f
C433 VTAIL.n339 VSUBS 0.031602f
C434 VTAIL.n340 VSUBS 0.01337f
C435 VTAIL.n341 VSUBS 0.014156f
C436 VTAIL.n342 VSUBS 0.024881f
C437 VTAIL.n343 VSUBS 0.01337f
C438 VTAIL.n344 VSUBS 0.031602f
C439 VTAIL.n345 VSUBS 0.014156f
C440 VTAIL.n346 VSUBS 0.024881f
C441 VTAIL.n347 VSUBS 0.01337f
C442 VTAIL.n348 VSUBS 0.023701f
C443 VTAIL.n349 VSUBS 0.023772f
C444 VTAIL.t9 VSUBS 0.06793f
C445 VTAIL.n350 VSUBS 0.171999f
C446 VTAIL.n351 VSUBS 0.990248f
C447 VTAIL.n352 VSUBS 0.01337f
C448 VTAIL.n353 VSUBS 0.014156f
C449 VTAIL.n354 VSUBS 0.031602f
C450 VTAIL.n355 VSUBS 0.031602f
C451 VTAIL.n356 VSUBS 0.014156f
C452 VTAIL.n357 VSUBS 0.01337f
C453 VTAIL.n358 VSUBS 0.024881f
C454 VTAIL.n359 VSUBS 0.024881f
C455 VTAIL.n360 VSUBS 0.01337f
C456 VTAIL.n361 VSUBS 0.014156f
C457 VTAIL.n362 VSUBS 0.031602f
C458 VTAIL.n363 VSUBS 0.031602f
C459 VTAIL.n364 VSUBS 0.014156f
C460 VTAIL.n365 VSUBS 0.01337f
C461 VTAIL.n366 VSUBS 0.024881f
C462 VTAIL.n367 VSUBS 0.024881f
C463 VTAIL.n368 VSUBS 0.01337f
C464 VTAIL.n369 VSUBS 0.014156f
C465 VTAIL.n370 VSUBS 0.031602f
C466 VTAIL.n371 VSUBS 0.031602f
C467 VTAIL.n372 VSUBS 0.031602f
C468 VTAIL.n373 VSUBS 0.013763f
C469 VTAIL.n374 VSUBS 0.01337f
C470 VTAIL.n375 VSUBS 0.024881f
C471 VTAIL.n376 VSUBS 0.024881f
C472 VTAIL.n377 VSUBS 0.01337f
C473 VTAIL.n378 VSUBS 0.014156f
C474 VTAIL.n379 VSUBS 0.031602f
C475 VTAIL.n380 VSUBS 0.068605f
C476 VTAIL.n381 VSUBS 0.014156f
C477 VTAIL.n382 VSUBS 0.01337f
C478 VTAIL.n383 VSUBS 0.054452f
C479 VTAIL.n384 VSUBS 0.034054f
C480 VTAIL.n385 VSUBS 1.25667f
C481 VTAIL.n386 VSUBS 0.02502f
C482 VTAIL.n387 VSUBS 0.024881f
C483 VTAIL.n388 VSUBS 0.01337f
C484 VTAIL.n389 VSUBS 0.031602f
C485 VTAIL.n390 VSUBS 0.014156f
C486 VTAIL.n391 VSUBS 0.024881f
C487 VTAIL.n392 VSUBS 0.013763f
C488 VTAIL.n393 VSUBS 0.031602f
C489 VTAIL.n394 VSUBS 0.014156f
C490 VTAIL.n395 VSUBS 0.024881f
C491 VTAIL.n396 VSUBS 0.01337f
C492 VTAIL.n397 VSUBS 0.031602f
C493 VTAIL.n398 VSUBS 0.014156f
C494 VTAIL.n399 VSUBS 0.024881f
C495 VTAIL.n400 VSUBS 0.01337f
C496 VTAIL.n401 VSUBS 0.023701f
C497 VTAIL.n402 VSUBS 0.023772f
C498 VTAIL.t4 VSUBS 0.06793f
C499 VTAIL.n403 VSUBS 0.171999f
C500 VTAIL.n404 VSUBS 0.990248f
C501 VTAIL.n405 VSUBS 0.01337f
C502 VTAIL.n406 VSUBS 0.014156f
C503 VTAIL.n407 VSUBS 0.031602f
C504 VTAIL.n408 VSUBS 0.031602f
C505 VTAIL.n409 VSUBS 0.014156f
C506 VTAIL.n410 VSUBS 0.01337f
C507 VTAIL.n411 VSUBS 0.024881f
C508 VTAIL.n412 VSUBS 0.024881f
C509 VTAIL.n413 VSUBS 0.01337f
C510 VTAIL.n414 VSUBS 0.014156f
C511 VTAIL.n415 VSUBS 0.031602f
C512 VTAIL.n416 VSUBS 0.031602f
C513 VTAIL.n417 VSUBS 0.014156f
C514 VTAIL.n418 VSUBS 0.01337f
C515 VTAIL.n419 VSUBS 0.024881f
C516 VTAIL.n420 VSUBS 0.024881f
C517 VTAIL.n421 VSUBS 0.01337f
C518 VTAIL.n422 VSUBS 0.01337f
C519 VTAIL.n423 VSUBS 0.014156f
C520 VTAIL.n424 VSUBS 0.031602f
C521 VTAIL.n425 VSUBS 0.031602f
C522 VTAIL.n426 VSUBS 0.031602f
C523 VTAIL.n427 VSUBS 0.013763f
C524 VTAIL.n428 VSUBS 0.01337f
C525 VTAIL.n429 VSUBS 0.024881f
C526 VTAIL.n430 VSUBS 0.024881f
C527 VTAIL.n431 VSUBS 0.01337f
C528 VTAIL.n432 VSUBS 0.014156f
C529 VTAIL.n433 VSUBS 0.031602f
C530 VTAIL.n434 VSUBS 0.068605f
C531 VTAIL.n435 VSUBS 0.014156f
C532 VTAIL.n436 VSUBS 0.01337f
C533 VTAIL.n437 VSUBS 0.054452f
C534 VTAIL.n438 VSUBS 0.034054f
C535 VTAIL.n439 VSUBS 1.25201f
C536 VDD1.t5 VSUBS 0.198337f
C537 VDD1.t3 VSUBS 0.198337f
C538 VDD1.n0 VSUBS 1.49438f
C539 VDD1.t7 VSUBS 0.198337f
C540 VDD1.t4 VSUBS 0.198337f
C541 VDD1.n1 VSUBS 1.49335f
C542 VDD1.t2 VSUBS 0.198337f
C543 VDD1.t0 VSUBS 0.198337f
C544 VDD1.n2 VSUBS 1.49335f
C545 VDD1.n3 VSUBS 2.95731f
C546 VDD1.t6 VSUBS 0.198337f
C547 VDD1.t1 VSUBS 0.198337f
C548 VDD1.n4 VSUBS 1.48814f
C549 VDD1.n5 VSUBS 2.63698f
C550 VP.n0 VSUBS 0.060493f
C551 VP.t3 VSUBS 1.5024f
C552 VP.n1 VSUBS 0.560014f
C553 VP.n2 VSUBS 0.045334f
C554 VP.t4 VSUBS 1.5024f
C555 VP.n3 VSUBS 0.560014f
C556 VP.n4 VSUBS 0.060493f
C557 VP.n5 VSUBS 0.060493f
C558 VP.t6 VSUBS 1.58852f
C559 VP.t1 VSUBS 1.5024f
C560 VP.n6 VSUBS 0.560014f
C561 VP.n7 VSUBS 0.045334f
C562 VP.t7 VSUBS 1.5024f
C563 VP.n8 VSUBS 0.620393f
C564 VP.t0 VSUBS 1.64189f
C565 VP.n9 VSUBS 0.635694f
C566 VP.n10 VSUBS 0.237099f
C567 VP.n11 VSUBS 0.072162f
C568 VP.n12 VSUBS 0.036648f
C569 VP.n13 VSUBS 0.072162f
C570 VP.n14 VSUBS 0.045334f
C571 VP.n15 VSUBS 0.045334f
C572 VP.n16 VSUBS 0.067792f
C573 VP.n17 VSUBS 0.031722f
C574 VP.n18 VSUBS 0.64778f
C575 VP.n19 VSUBS 1.96792f
C576 VP.n20 VSUBS 2.00574f
C577 VP.t5 VSUBS 1.58852f
C578 VP.n21 VSUBS 0.64778f
C579 VP.n22 VSUBS 0.031722f
C580 VP.n23 VSUBS 0.067792f
C581 VP.n24 VSUBS 0.045334f
C582 VP.n25 VSUBS 0.045334f
C583 VP.n26 VSUBS 0.072162f
C584 VP.n27 VSUBS 0.036648f
C585 VP.n28 VSUBS 0.072162f
C586 VP.n29 VSUBS 0.045334f
C587 VP.n30 VSUBS 0.045334f
C588 VP.n31 VSUBS 0.067792f
C589 VP.n32 VSUBS 0.031722f
C590 VP.t2 VSUBS 1.58852f
C591 VP.n33 VSUBS 0.64778f
C592 VP.n34 VSUBS 0.042457f
C593 B.n0 VSUBS 0.004984f
C594 B.n1 VSUBS 0.004984f
C595 B.n2 VSUBS 0.007882f
C596 B.n3 VSUBS 0.007882f
C597 B.n4 VSUBS 0.007882f
C598 B.n5 VSUBS 0.007882f
C599 B.n6 VSUBS 0.007882f
C600 B.n7 VSUBS 0.007882f
C601 B.n8 VSUBS 0.007882f
C602 B.n9 VSUBS 0.007882f
C603 B.n10 VSUBS 0.007882f
C604 B.n11 VSUBS 0.007882f
C605 B.n12 VSUBS 0.007882f
C606 B.n13 VSUBS 0.007882f
C607 B.n14 VSUBS 0.007882f
C608 B.n15 VSUBS 0.007882f
C609 B.n16 VSUBS 0.007882f
C610 B.n17 VSUBS 0.019262f
C611 B.n18 VSUBS 0.007882f
C612 B.n19 VSUBS 0.007882f
C613 B.n20 VSUBS 0.007882f
C614 B.n21 VSUBS 0.007882f
C615 B.n22 VSUBS 0.007882f
C616 B.n23 VSUBS 0.007882f
C617 B.n24 VSUBS 0.007882f
C618 B.n25 VSUBS 0.007882f
C619 B.n26 VSUBS 0.007882f
C620 B.n27 VSUBS 0.007882f
C621 B.n28 VSUBS 0.007882f
C622 B.n29 VSUBS 0.007882f
C623 B.n30 VSUBS 0.007882f
C624 B.n31 VSUBS 0.007882f
C625 B.n32 VSUBS 0.007882f
C626 B.n33 VSUBS 0.007882f
C627 B.n34 VSUBS 0.007882f
C628 B.n35 VSUBS 0.007882f
C629 B.t11 VSUBS 0.185256f
C630 B.t10 VSUBS 0.204445f
C631 B.t9 VSUBS 0.601963f
C632 B.n36 VSUBS 0.32325f
C633 B.n37 VSUBS 0.242852f
C634 B.n38 VSUBS 0.007882f
C635 B.n39 VSUBS 0.007882f
C636 B.n40 VSUBS 0.007882f
C637 B.n41 VSUBS 0.007882f
C638 B.t8 VSUBS 0.185259f
C639 B.t7 VSUBS 0.204448f
C640 B.t6 VSUBS 0.601963f
C641 B.n42 VSUBS 0.323247f
C642 B.n43 VSUBS 0.242849f
C643 B.n44 VSUBS 0.018261f
C644 B.n45 VSUBS 0.007882f
C645 B.n46 VSUBS 0.007882f
C646 B.n47 VSUBS 0.007882f
C647 B.n48 VSUBS 0.007882f
C648 B.n49 VSUBS 0.007882f
C649 B.n50 VSUBS 0.007882f
C650 B.n51 VSUBS 0.007882f
C651 B.n52 VSUBS 0.007882f
C652 B.n53 VSUBS 0.007882f
C653 B.n54 VSUBS 0.007882f
C654 B.n55 VSUBS 0.007882f
C655 B.n56 VSUBS 0.007882f
C656 B.n57 VSUBS 0.007882f
C657 B.n58 VSUBS 0.007882f
C658 B.n59 VSUBS 0.007882f
C659 B.n60 VSUBS 0.007882f
C660 B.n61 VSUBS 0.007882f
C661 B.n62 VSUBS 0.020105f
C662 B.n63 VSUBS 0.007882f
C663 B.n64 VSUBS 0.007882f
C664 B.n65 VSUBS 0.007882f
C665 B.n66 VSUBS 0.007882f
C666 B.n67 VSUBS 0.007882f
C667 B.n68 VSUBS 0.007882f
C668 B.n69 VSUBS 0.007882f
C669 B.n70 VSUBS 0.007882f
C670 B.n71 VSUBS 0.007882f
C671 B.n72 VSUBS 0.007882f
C672 B.n73 VSUBS 0.007882f
C673 B.n74 VSUBS 0.007882f
C674 B.n75 VSUBS 0.007882f
C675 B.n76 VSUBS 0.007882f
C676 B.n77 VSUBS 0.007882f
C677 B.n78 VSUBS 0.007882f
C678 B.n79 VSUBS 0.007882f
C679 B.n80 VSUBS 0.007882f
C680 B.n81 VSUBS 0.007882f
C681 B.n82 VSUBS 0.007882f
C682 B.n83 VSUBS 0.007882f
C683 B.n84 VSUBS 0.007882f
C684 B.n85 VSUBS 0.007882f
C685 B.n86 VSUBS 0.007882f
C686 B.n87 VSUBS 0.007882f
C687 B.n88 VSUBS 0.007882f
C688 B.n89 VSUBS 0.007882f
C689 B.n90 VSUBS 0.007882f
C690 B.n91 VSUBS 0.007882f
C691 B.n92 VSUBS 0.007882f
C692 B.n93 VSUBS 0.019262f
C693 B.n94 VSUBS 0.007882f
C694 B.n95 VSUBS 0.007882f
C695 B.n96 VSUBS 0.007882f
C696 B.n97 VSUBS 0.007882f
C697 B.n98 VSUBS 0.007882f
C698 B.n99 VSUBS 0.007882f
C699 B.n100 VSUBS 0.007882f
C700 B.n101 VSUBS 0.007882f
C701 B.n102 VSUBS 0.007882f
C702 B.n103 VSUBS 0.007882f
C703 B.n104 VSUBS 0.007882f
C704 B.n105 VSUBS 0.007882f
C705 B.n106 VSUBS 0.007882f
C706 B.n107 VSUBS 0.007882f
C707 B.n108 VSUBS 0.007882f
C708 B.n109 VSUBS 0.007882f
C709 B.n110 VSUBS 0.007882f
C710 B.n111 VSUBS 0.007882f
C711 B.t4 VSUBS 0.185259f
C712 B.t5 VSUBS 0.204448f
C713 B.t3 VSUBS 0.601963f
C714 B.n112 VSUBS 0.323247f
C715 B.n113 VSUBS 0.242849f
C716 B.n114 VSUBS 0.007882f
C717 B.n115 VSUBS 0.007882f
C718 B.n116 VSUBS 0.007882f
C719 B.n117 VSUBS 0.007882f
C720 B.t1 VSUBS 0.185256f
C721 B.t2 VSUBS 0.204445f
C722 B.t0 VSUBS 0.601963f
C723 B.n118 VSUBS 0.32325f
C724 B.n119 VSUBS 0.242852f
C725 B.n120 VSUBS 0.018261f
C726 B.n121 VSUBS 0.007882f
C727 B.n122 VSUBS 0.007882f
C728 B.n123 VSUBS 0.007882f
C729 B.n124 VSUBS 0.007882f
C730 B.n125 VSUBS 0.007882f
C731 B.n126 VSUBS 0.007882f
C732 B.n127 VSUBS 0.007882f
C733 B.n128 VSUBS 0.007882f
C734 B.n129 VSUBS 0.007882f
C735 B.n130 VSUBS 0.007882f
C736 B.n131 VSUBS 0.007882f
C737 B.n132 VSUBS 0.007882f
C738 B.n133 VSUBS 0.007882f
C739 B.n134 VSUBS 0.007882f
C740 B.n135 VSUBS 0.007882f
C741 B.n136 VSUBS 0.007882f
C742 B.n137 VSUBS 0.007882f
C743 B.n138 VSUBS 0.019262f
C744 B.n139 VSUBS 0.007882f
C745 B.n140 VSUBS 0.007882f
C746 B.n141 VSUBS 0.007882f
C747 B.n142 VSUBS 0.007882f
C748 B.n143 VSUBS 0.007882f
C749 B.n144 VSUBS 0.007882f
C750 B.n145 VSUBS 0.007882f
C751 B.n146 VSUBS 0.007882f
C752 B.n147 VSUBS 0.007882f
C753 B.n148 VSUBS 0.007882f
C754 B.n149 VSUBS 0.007882f
C755 B.n150 VSUBS 0.007882f
C756 B.n151 VSUBS 0.007882f
C757 B.n152 VSUBS 0.007882f
C758 B.n153 VSUBS 0.007882f
C759 B.n154 VSUBS 0.007882f
C760 B.n155 VSUBS 0.007882f
C761 B.n156 VSUBS 0.007882f
C762 B.n157 VSUBS 0.007882f
C763 B.n158 VSUBS 0.007882f
C764 B.n159 VSUBS 0.007882f
C765 B.n160 VSUBS 0.007882f
C766 B.n161 VSUBS 0.007882f
C767 B.n162 VSUBS 0.007882f
C768 B.n163 VSUBS 0.007882f
C769 B.n164 VSUBS 0.007882f
C770 B.n165 VSUBS 0.007882f
C771 B.n166 VSUBS 0.007882f
C772 B.n167 VSUBS 0.007882f
C773 B.n168 VSUBS 0.007882f
C774 B.n169 VSUBS 0.007882f
C775 B.n170 VSUBS 0.007882f
C776 B.n171 VSUBS 0.007882f
C777 B.n172 VSUBS 0.007882f
C778 B.n173 VSUBS 0.007882f
C779 B.n174 VSUBS 0.007882f
C780 B.n175 VSUBS 0.007882f
C781 B.n176 VSUBS 0.007882f
C782 B.n177 VSUBS 0.007882f
C783 B.n178 VSUBS 0.007882f
C784 B.n179 VSUBS 0.007882f
C785 B.n180 VSUBS 0.007882f
C786 B.n181 VSUBS 0.007882f
C787 B.n182 VSUBS 0.007882f
C788 B.n183 VSUBS 0.007882f
C789 B.n184 VSUBS 0.007882f
C790 B.n185 VSUBS 0.007882f
C791 B.n186 VSUBS 0.007882f
C792 B.n187 VSUBS 0.007882f
C793 B.n188 VSUBS 0.007882f
C794 B.n189 VSUBS 0.007882f
C795 B.n190 VSUBS 0.007882f
C796 B.n191 VSUBS 0.007882f
C797 B.n192 VSUBS 0.007882f
C798 B.n193 VSUBS 0.007882f
C799 B.n194 VSUBS 0.007882f
C800 B.n195 VSUBS 0.007882f
C801 B.n196 VSUBS 0.007882f
C802 B.n197 VSUBS 0.019262f
C803 B.n198 VSUBS 0.020147f
C804 B.n199 VSUBS 0.020147f
C805 B.n200 VSUBS 0.007882f
C806 B.n201 VSUBS 0.007882f
C807 B.n202 VSUBS 0.007882f
C808 B.n203 VSUBS 0.007882f
C809 B.n204 VSUBS 0.007882f
C810 B.n205 VSUBS 0.007882f
C811 B.n206 VSUBS 0.007882f
C812 B.n207 VSUBS 0.007882f
C813 B.n208 VSUBS 0.007882f
C814 B.n209 VSUBS 0.007882f
C815 B.n210 VSUBS 0.007882f
C816 B.n211 VSUBS 0.007882f
C817 B.n212 VSUBS 0.007882f
C818 B.n213 VSUBS 0.007882f
C819 B.n214 VSUBS 0.007882f
C820 B.n215 VSUBS 0.007882f
C821 B.n216 VSUBS 0.007882f
C822 B.n217 VSUBS 0.007882f
C823 B.n218 VSUBS 0.007882f
C824 B.n219 VSUBS 0.007882f
C825 B.n220 VSUBS 0.007882f
C826 B.n221 VSUBS 0.007882f
C827 B.n222 VSUBS 0.007882f
C828 B.n223 VSUBS 0.007882f
C829 B.n224 VSUBS 0.007882f
C830 B.n225 VSUBS 0.007882f
C831 B.n226 VSUBS 0.007882f
C832 B.n227 VSUBS 0.007882f
C833 B.n228 VSUBS 0.007882f
C834 B.n229 VSUBS 0.007882f
C835 B.n230 VSUBS 0.007882f
C836 B.n231 VSUBS 0.007882f
C837 B.n232 VSUBS 0.007882f
C838 B.n233 VSUBS 0.007882f
C839 B.n234 VSUBS 0.007882f
C840 B.n235 VSUBS 0.007882f
C841 B.n236 VSUBS 0.007882f
C842 B.n237 VSUBS 0.007882f
C843 B.n238 VSUBS 0.007882f
C844 B.n239 VSUBS 0.007882f
C845 B.n240 VSUBS 0.007882f
C846 B.n241 VSUBS 0.007882f
C847 B.n242 VSUBS 0.007882f
C848 B.n243 VSUBS 0.007882f
C849 B.n244 VSUBS 0.007882f
C850 B.n245 VSUBS 0.007882f
C851 B.n246 VSUBS 0.007882f
C852 B.n247 VSUBS 0.007882f
C853 B.n248 VSUBS 0.007882f
C854 B.n249 VSUBS 0.007418f
C855 B.n250 VSUBS 0.007882f
C856 B.n251 VSUBS 0.007882f
C857 B.n252 VSUBS 0.004405f
C858 B.n253 VSUBS 0.007882f
C859 B.n254 VSUBS 0.007882f
C860 B.n255 VSUBS 0.007882f
C861 B.n256 VSUBS 0.007882f
C862 B.n257 VSUBS 0.007882f
C863 B.n258 VSUBS 0.007882f
C864 B.n259 VSUBS 0.007882f
C865 B.n260 VSUBS 0.007882f
C866 B.n261 VSUBS 0.007882f
C867 B.n262 VSUBS 0.007882f
C868 B.n263 VSUBS 0.007882f
C869 B.n264 VSUBS 0.007882f
C870 B.n265 VSUBS 0.004405f
C871 B.n266 VSUBS 0.018261f
C872 B.n267 VSUBS 0.007418f
C873 B.n268 VSUBS 0.007882f
C874 B.n269 VSUBS 0.007882f
C875 B.n270 VSUBS 0.007882f
C876 B.n271 VSUBS 0.007882f
C877 B.n272 VSUBS 0.007882f
C878 B.n273 VSUBS 0.007882f
C879 B.n274 VSUBS 0.007882f
C880 B.n275 VSUBS 0.007882f
C881 B.n276 VSUBS 0.007882f
C882 B.n277 VSUBS 0.007882f
C883 B.n278 VSUBS 0.007882f
C884 B.n279 VSUBS 0.007882f
C885 B.n280 VSUBS 0.007882f
C886 B.n281 VSUBS 0.007882f
C887 B.n282 VSUBS 0.007882f
C888 B.n283 VSUBS 0.007882f
C889 B.n284 VSUBS 0.007882f
C890 B.n285 VSUBS 0.007882f
C891 B.n286 VSUBS 0.007882f
C892 B.n287 VSUBS 0.007882f
C893 B.n288 VSUBS 0.007882f
C894 B.n289 VSUBS 0.007882f
C895 B.n290 VSUBS 0.007882f
C896 B.n291 VSUBS 0.007882f
C897 B.n292 VSUBS 0.007882f
C898 B.n293 VSUBS 0.007882f
C899 B.n294 VSUBS 0.007882f
C900 B.n295 VSUBS 0.007882f
C901 B.n296 VSUBS 0.007882f
C902 B.n297 VSUBS 0.007882f
C903 B.n298 VSUBS 0.007882f
C904 B.n299 VSUBS 0.007882f
C905 B.n300 VSUBS 0.007882f
C906 B.n301 VSUBS 0.007882f
C907 B.n302 VSUBS 0.007882f
C908 B.n303 VSUBS 0.007882f
C909 B.n304 VSUBS 0.007882f
C910 B.n305 VSUBS 0.007882f
C911 B.n306 VSUBS 0.007882f
C912 B.n307 VSUBS 0.007882f
C913 B.n308 VSUBS 0.007882f
C914 B.n309 VSUBS 0.007882f
C915 B.n310 VSUBS 0.007882f
C916 B.n311 VSUBS 0.007882f
C917 B.n312 VSUBS 0.007882f
C918 B.n313 VSUBS 0.007882f
C919 B.n314 VSUBS 0.007882f
C920 B.n315 VSUBS 0.007882f
C921 B.n316 VSUBS 0.007882f
C922 B.n317 VSUBS 0.007882f
C923 B.n318 VSUBS 0.020147f
C924 B.n319 VSUBS 0.020147f
C925 B.n320 VSUBS 0.019262f
C926 B.n321 VSUBS 0.007882f
C927 B.n322 VSUBS 0.007882f
C928 B.n323 VSUBS 0.007882f
C929 B.n324 VSUBS 0.007882f
C930 B.n325 VSUBS 0.007882f
C931 B.n326 VSUBS 0.007882f
C932 B.n327 VSUBS 0.007882f
C933 B.n328 VSUBS 0.007882f
C934 B.n329 VSUBS 0.007882f
C935 B.n330 VSUBS 0.007882f
C936 B.n331 VSUBS 0.007882f
C937 B.n332 VSUBS 0.007882f
C938 B.n333 VSUBS 0.007882f
C939 B.n334 VSUBS 0.007882f
C940 B.n335 VSUBS 0.007882f
C941 B.n336 VSUBS 0.007882f
C942 B.n337 VSUBS 0.007882f
C943 B.n338 VSUBS 0.007882f
C944 B.n339 VSUBS 0.007882f
C945 B.n340 VSUBS 0.007882f
C946 B.n341 VSUBS 0.007882f
C947 B.n342 VSUBS 0.007882f
C948 B.n343 VSUBS 0.007882f
C949 B.n344 VSUBS 0.007882f
C950 B.n345 VSUBS 0.007882f
C951 B.n346 VSUBS 0.007882f
C952 B.n347 VSUBS 0.007882f
C953 B.n348 VSUBS 0.007882f
C954 B.n349 VSUBS 0.007882f
C955 B.n350 VSUBS 0.007882f
C956 B.n351 VSUBS 0.007882f
C957 B.n352 VSUBS 0.007882f
C958 B.n353 VSUBS 0.007882f
C959 B.n354 VSUBS 0.007882f
C960 B.n355 VSUBS 0.007882f
C961 B.n356 VSUBS 0.007882f
C962 B.n357 VSUBS 0.007882f
C963 B.n358 VSUBS 0.007882f
C964 B.n359 VSUBS 0.007882f
C965 B.n360 VSUBS 0.007882f
C966 B.n361 VSUBS 0.007882f
C967 B.n362 VSUBS 0.007882f
C968 B.n363 VSUBS 0.007882f
C969 B.n364 VSUBS 0.007882f
C970 B.n365 VSUBS 0.007882f
C971 B.n366 VSUBS 0.007882f
C972 B.n367 VSUBS 0.007882f
C973 B.n368 VSUBS 0.007882f
C974 B.n369 VSUBS 0.007882f
C975 B.n370 VSUBS 0.007882f
C976 B.n371 VSUBS 0.007882f
C977 B.n372 VSUBS 0.007882f
C978 B.n373 VSUBS 0.007882f
C979 B.n374 VSUBS 0.007882f
C980 B.n375 VSUBS 0.007882f
C981 B.n376 VSUBS 0.007882f
C982 B.n377 VSUBS 0.007882f
C983 B.n378 VSUBS 0.007882f
C984 B.n379 VSUBS 0.007882f
C985 B.n380 VSUBS 0.007882f
C986 B.n381 VSUBS 0.007882f
C987 B.n382 VSUBS 0.007882f
C988 B.n383 VSUBS 0.007882f
C989 B.n384 VSUBS 0.007882f
C990 B.n385 VSUBS 0.007882f
C991 B.n386 VSUBS 0.007882f
C992 B.n387 VSUBS 0.007882f
C993 B.n388 VSUBS 0.007882f
C994 B.n389 VSUBS 0.007882f
C995 B.n390 VSUBS 0.007882f
C996 B.n391 VSUBS 0.007882f
C997 B.n392 VSUBS 0.007882f
C998 B.n393 VSUBS 0.007882f
C999 B.n394 VSUBS 0.007882f
C1000 B.n395 VSUBS 0.007882f
C1001 B.n396 VSUBS 0.007882f
C1002 B.n397 VSUBS 0.007882f
C1003 B.n398 VSUBS 0.007882f
C1004 B.n399 VSUBS 0.007882f
C1005 B.n400 VSUBS 0.007882f
C1006 B.n401 VSUBS 0.007882f
C1007 B.n402 VSUBS 0.007882f
C1008 B.n403 VSUBS 0.007882f
C1009 B.n404 VSUBS 0.007882f
C1010 B.n405 VSUBS 0.007882f
C1011 B.n406 VSUBS 0.007882f
C1012 B.n407 VSUBS 0.007882f
C1013 B.n408 VSUBS 0.007882f
C1014 B.n409 VSUBS 0.007882f
C1015 B.n410 VSUBS 0.007882f
C1016 B.n411 VSUBS 0.007882f
C1017 B.n412 VSUBS 0.007882f
C1018 B.n413 VSUBS 0.019262f
C1019 B.n414 VSUBS 0.020147f
C1020 B.n415 VSUBS 0.019303f
C1021 B.n416 VSUBS 0.007882f
C1022 B.n417 VSUBS 0.007882f
C1023 B.n418 VSUBS 0.007882f
C1024 B.n419 VSUBS 0.007882f
C1025 B.n420 VSUBS 0.007882f
C1026 B.n421 VSUBS 0.007882f
C1027 B.n422 VSUBS 0.007882f
C1028 B.n423 VSUBS 0.007882f
C1029 B.n424 VSUBS 0.007882f
C1030 B.n425 VSUBS 0.007882f
C1031 B.n426 VSUBS 0.007882f
C1032 B.n427 VSUBS 0.007882f
C1033 B.n428 VSUBS 0.007882f
C1034 B.n429 VSUBS 0.007882f
C1035 B.n430 VSUBS 0.007882f
C1036 B.n431 VSUBS 0.007882f
C1037 B.n432 VSUBS 0.007882f
C1038 B.n433 VSUBS 0.007882f
C1039 B.n434 VSUBS 0.007882f
C1040 B.n435 VSUBS 0.007882f
C1041 B.n436 VSUBS 0.007882f
C1042 B.n437 VSUBS 0.007882f
C1043 B.n438 VSUBS 0.007882f
C1044 B.n439 VSUBS 0.007882f
C1045 B.n440 VSUBS 0.007882f
C1046 B.n441 VSUBS 0.007882f
C1047 B.n442 VSUBS 0.007882f
C1048 B.n443 VSUBS 0.007882f
C1049 B.n444 VSUBS 0.007882f
C1050 B.n445 VSUBS 0.007882f
C1051 B.n446 VSUBS 0.007882f
C1052 B.n447 VSUBS 0.007882f
C1053 B.n448 VSUBS 0.007882f
C1054 B.n449 VSUBS 0.007882f
C1055 B.n450 VSUBS 0.007882f
C1056 B.n451 VSUBS 0.007882f
C1057 B.n452 VSUBS 0.007882f
C1058 B.n453 VSUBS 0.007882f
C1059 B.n454 VSUBS 0.007882f
C1060 B.n455 VSUBS 0.007882f
C1061 B.n456 VSUBS 0.007882f
C1062 B.n457 VSUBS 0.007882f
C1063 B.n458 VSUBS 0.007882f
C1064 B.n459 VSUBS 0.007882f
C1065 B.n460 VSUBS 0.007882f
C1066 B.n461 VSUBS 0.007882f
C1067 B.n462 VSUBS 0.007882f
C1068 B.n463 VSUBS 0.007882f
C1069 B.n464 VSUBS 0.007882f
C1070 B.n465 VSUBS 0.007418f
C1071 B.n466 VSUBS 0.007882f
C1072 B.n467 VSUBS 0.007882f
C1073 B.n468 VSUBS 0.004405f
C1074 B.n469 VSUBS 0.007882f
C1075 B.n470 VSUBS 0.007882f
C1076 B.n471 VSUBS 0.007882f
C1077 B.n472 VSUBS 0.007882f
C1078 B.n473 VSUBS 0.007882f
C1079 B.n474 VSUBS 0.007882f
C1080 B.n475 VSUBS 0.007882f
C1081 B.n476 VSUBS 0.007882f
C1082 B.n477 VSUBS 0.007882f
C1083 B.n478 VSUBS 0.007882f
C1084 B.n479 VSUBS 0.007882f
C1085 B.n480 VSUBS 0.007882f
C1086 B.n481 VSUBS 0.004405f
C1087 B.n482 VSUBS 0.018261f
C1088 B.n483 VSUBS 0.007418f
C1089 B.n484 VSUBS 0.007882f
C1090 B.n485 VSUBS 0.007882f
C1091 B.n486 VSUBS 0.007882f
C1092 B.n487 VSUBS 0.007882f
C1093 B.n488 VSUBS 0.007882f
C1094 B.n489 VSUBS 0.007882f
C1095 B.n490 VSUBS 0.007882f
C1096 B.n491 VSUBS 0.007882f
C1097 B.n492 VSUBS 0.007882f
C1098 B.n493 VSUBS 0.007882f
C1099 B.n494 VSUBS 0.007882f
C1100 B.n495 VSUBS 0.007882f
C1101 B.n496 VSUBS 0.007882f
C1102 B.n497 VSUBS 0.007882f
C1103 B.n498 VSUBS 0.007882f
C1104 B.n499 VSUBS 0.007882f
C1105 B.n500 VSUBS 0.007882f
C1106 B.n501 VSUBS 0.007882f
C1107 B.n502 VSUBS 0.007882f
C1108 B.n503 VSUBS 0.007882f
C1109 B.n504 VSUBS 0.007882f
C1110 B.n505 VSUBS 0.007882f
C1111 B.n506 VSUBS 0.007882f
C1112 B.n507 VSUBS 0.007882f
C1113 B.n508 VSUBS 0.007882f
C1114 B.n509 VSUBS 0.007882f
C1115 B.n510 VSUBS 0.007882f
C1116 B.n511 VSUBS 0.007882f
C1117 B.n512 VSUBS 0.007882f
C1118 B.n513 VSUBS 0.007882f
C1119 B.n514 VSUBS 0.007882f
C1120 B.n515 VSUBS 0.007882f
C1121 B.n516 VSUBS 0.007882f
C1122 B.n517 VSUBS 0.007882f
C1123 B.n518 VSUBS 0.007882f
C1124 B.n519 VSUBS 0.007882f
C1125 B.n520 VSUBS 0.007882f
C1126 B.n521 VSUBS 0.007882f
C1127 B.n522 VSUBS 0.007882f
C1128 B.n523 VSUBS 0.007882f
C1129 B.n524 VSUBS 0.007882f
C1130 B.n525 VSUBS 0.007882f
C1131 B.n526 VSUBS 0.007882f
C1132 B.n527 VSUBS 0.007882f
C1133 B.n528 VSUBS 0.007882f
C1134 B.n529 VSUBS 0.007882f
C1135 B.n530 VSUBS 0.007882f
C1136 B.n531 VSUBS 0.007882f
C1137 B.n532 VSUBS 0.007882f
C1138 B.n533 VSUBS 0.007882f
C1139 B.n534 VSUBS 0.020147f
C1140 B.n535 VSUBS 0.020147f
C1141 B.n536 VSUBS 0.019262f
C1142 B.n537 VSUBS 0.007882f
C1143 B.n538 VSUBS 0.007882f
C1144 B.n539 VSUBS 0.007882f
C1145 B.n540 VSUBS 0.007882f
C1146 B.n541 VSUBS 0.007882f
C1147 B.n542 VSUBS 0.007882f
C1148 B.n543 VSUBS 0.007882f
C1149 B.n544 VSUBS 0.007882f
C1150 B.n545 VSUBS 0.007882f
C1151 B.n546 VSUBS 0.007882f
C1152 B.n547 VSUBS 0.007882f
C1153 B.n548 VSUBS 0.007882f
C1154 B.n549 VSUBS 0.007882f
C1155 B.n550 VSUBS 0.007882f
C1156 B.n551 VSUBS 0.007882f
C1157 B.n552 VSUBS 0.007882f
C1158 B.n553 VSUBS 0.007882f
C1159 B.n554 VSUBS 0.007882f
C1160 B.n555 VSUBS 0.007882f
C1161 B.n556 VSUBS 0.007882f
C1162 B.n557 VSUBS 0.007882f
C1163 B.n558 VSUBS 0.007882f
C1164 B.n559 VSUBS 0.007882f
C1165 B.n560 VSUBS 0.007882f
C1166 B.n561 VSUBS 0.007882f
C1167 B.n562 VSUBS 0.007882f
C1168 B.n563 VSUBS 0.007882f
C1169 B.n564 VSUBS 0.007882f
C1170 B.n565 VSUBS 0.007882f
C1171 B.n566 VSUBS 0.007882f
C1172 B.n567 VSUBS 0.007882f
C1173 B.n568 VSUBS 0.007882f
C1174 B.n569 VSUBS 0.007882f
C1175 B.n570 VSUBS 0.007882f
C1176 B.n571 VSUBS 0.007882f
C1177 B.n572 VSUBS 0.007882f
C1178 B.n573 VSUBS 0.007882f
C1179 B.n574 VSUBS 0.007882f
C1180 B.n575 VSUBS 0.007882f
C1181 B.n576 VSUBS 0.007882f
C1182 B.n577 VSUBS 0.007882f
C1183 B.n578 VSUBS 0.007882f
C1184 B.n579 VSUBS 0.007882f
C1185 B.n580 VSUBS 0.007882f
C1186 B.n581 VSUBS 0.007882f
C1187 B.n582 VSUBS 0.007882f
C1188 B.n583 VSUBS 0.017847f
.ends

