* NGSPICE file created from diff_pair_sample_0286.ext - technology: sky130A

.subckt diff_pair_sample_0286 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t13 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X1 VTAIL.t3 VP.t0 VDD1.t7 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X2 VTAIL.t9 VN.t1 VDD2.t6 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=1.3299 ps=8.39 w=8.06 l=3.52
X3 VDD2.t5 VN.t2 VTAIL.t10 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=3.1434 ps=16.9 w=8.06 l=3.52
X4 VDD1.t6 VP.t1 VTAIL.t1 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=3.1434 ps=16.9 w=8.06 l=3.52
X5 VDD1.t5 VP.t2 VTAIL.t2 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X6 VTAIL.t12 VN.t3 VDD2.t4 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X7 VDD1.t4 VP.t3 VTAIL.t5 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=3.1434 ps=16.9 w=8.06 l=3.52
X8 VTAIL.t7 VP.t4 VDD1.t3 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X9 VDD2.t3 VN.t4 VTAIL.t15 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=3.1434 ps=16.9 w=8.06 l=3.52
X10 B.t11 B.t9 B.t10 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=0 ps=0 w=8.06 l=3.52
X11 VTAIL.t0 VP.t5 VDD1.t2 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=1.3299 ps=8.39 w=8.06 l=3.52
X12 VDD2.t2 VN.t5 VTAIL.t14 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X13 VTAIL.t8 VN.t6 VDD2.t1 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=1.3299 ps=8.39 w=8.06 l=3.52
X14 VDD1.t1 VP.t6 VTAIL.t4 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X15 VTAIL.t11 VN.t7 VDD2.t0 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=1.3299 pd=8.39 as=1.3299 ps=8.39 w=8.06 l=3.52
X16 B.t8 B.t6 B.t7 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=0 ps=0 w=8.06 l=3.52
X17 B.t5 B.t3 B.t4 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=0 ps=0 w=8.06 l=3.52
X18 VTAIL.t6 VP.t7 VDD1.t0 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=1.3299 ps=8.39 w=8.06 l=3.52
X19 B.t2 B.t0 B.t1 w_n4820_n2580# sky130_fd_pr__pfet_01v8 ad=3.1434 pd=16.9 as=0 ps=0 w=8.06 l=3.52
R0 VN.n68 VN.n67 161.3
R1 VN.n66 VN.n36 161.3
R2 VN.n65 VN.n64 161.3
R3 VN.n63 VN.n37 161.3
R4 VN.n62 VN.n61 161.3
R5 VN.n60 VN.n38 161.3
R6 VN.n59 VN.n58 161.3
R7 VN.n57 VN.n39 161.3
R8 VN.n56 VN.n55 161.3
R9 VN.n54 VN.n40 161.3
R10 VN.n53 VN.n52 161.3
R11 VN.n51 VN.n42 161.3
R12 VN.n50 VN.n49 161.3
R13 VN.n48 VN.n43 161.3
R14 VN.n47 VN.n46 161.3
R15 VN.n33 VN.n32 161.3
R16 VN.n31 VN.n1 161.3
R17 VN.n30 VN.n29 161.3
R18 VN.n28 VN.n2 161.3
R19 VN.n27 VN.n26 161.3
R20 VN.n25 VN.n3 161.3
R21 VN.n24 VN.n23 161.3
R22 VN.n22 VN.n4 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n18 VN.n5 161.3
R25 VN.n17 VN.n16 161.3
R26 VN.n15 VN.n6 161.3
R27 VN.n14 VN.n13 161.3
R28 VN.n12 VN.n7 161.3
R29 VN.n11 VN.n10 161.3
R30 VN.n45 VN.t4 88.9805
R31 VN.n9 VN.t6 88.9805
R32 VN.n34 VN.n0 76.5021
R33 VN.n69 VN.n35 76.5021
R34 VN.n8 VN.t5 55.184
R35 VN.n19 VN.t3 55.184
R36 VN.n0 VN.t2 55.184
R37 VN.n44 VN.t7 55.184
R38 VN.n41 VN.t0 55.184
R39 VN.n35 VN.t1 55.184
R40 VN.n26 VN.n2 55.0167
R41 VN.n61 VN.n37 55.0167
R42 VN.n9 VN.n8 53.7745
R43 VN.n45 VN.n44 53.7745
R44 VN VN.n69 52.5282
R45 VN.n13 VN.n6 40.4106
R46 VN.n17 VN.n6 40.4106
R47 VN.n49 VN.n42 40.4106
R48 VN.n53 VN.n42 40.4106
R49 VN.n30 VN.n2 25.8045
R50 VN.n65 VN.n37 25.8045
R51 VN.n12 VN.n11 24.3439
R52 VN.n13 VN.n12 24.3439
R53 VN.n18 VN.n17 24.3439
R54 VN.n20 VN.n18 24.3439
R55 VN.n24 VN.n4 24.3439
R56 VN.n25 VN.n24 24.3439
R57 VN.n26 VN.n25 24.3439
R58 VN.n31 VN.n30 24.3439
R59 VN.n32 VN.n31 24.3439
R60 VN.n49 VN.n48 24.3439
R61 VN.n48 VN.n47 24.3439
R62 VN.n61 VN.n60 24.3439
R63 VN.n60 VN.n59 24.3439
R64 VN.n59 VN.n39 24.3439
R65 VN.n55 VN.n54 24.3439
R66 VN.n54 VN.n53 24.3439
R67 VN.n67 VN.n66 24.3439
R68 VN.n66 VN.n65 24.3439
R69 VN.n11 VN.n8 20.6924
R70 VN.n20 VN.n19 20.6924
R71 VN.n47 VN.n44 20.6924
R72 VN.n55 VN.n41 20.6924
R73 VN.n32 VN.n0 13.3894
R74 VN.n67 VN.n35 13.3894
R75 VN.n19 VN.n4 3.65202
R76 VN.n41 VN.n39 3.65202
R77 VN.n46 VN.n45 3.05397
R78 VN.n10 VN.n9 3.05397
R79 VN.n69 VN.n68 0.355081
R80 VN.n34 VN.n33 0.355081
R81 VN VN.n34 0.26685
R82 VN.n68 VN.n36 0.189894
R83 VN.n64 VN.n36 0.189894
R84 VN.n64 VN.n63 0.189894
R85 VN.n63 VN.n62 0.189894
R86 VN.n62 VN.n38 0.189894
R87 VN.n58 VN.n38 0.189894
R88 VN.n58 VN.n57 0.189894
R89 VN.n57 VN.n56 0.189894
R90 VN.n56 VN.n40 0.189894
R91 VN.n52 VN.n40 0.189894
R92 VN.n52 VN.n51 0.189894
R93 VN.n51 VN.n50 0.189894
R94 VN.n50 VN.n43 0.189894
R95 VN.n46 VN.n43 0.189894
R96 VN.n10 VN.n7 0.189894
R97 VN.n14 VN.n7 0.189894
R98 VN.n15 VN.n14 0.189894
R99 VN.n16 VN.n15 0.189894
R100 VN.n16 VN.n5 0.189894
R101 VN.n21 VN.n5 0.189894
R102 VN.n22 VN.n21 0.189894
R103 VN.n23 VN.n22 0.189894
R104 VN.n23 VN.n3 0.189894
R105 VN.n27 VN.n3 0.189894
R106 VN.n28 VN.n27 0.189894
R107 VN.n29 VN.n28 0.189894
R108 VN.n29 VN.n1 0.189894
R109 VN.n33 VN.n1 0.189894
R110 VTAIL.n354 VTAIL.n316 756.745
R111 VTAIL.n40 VTAIL.n2 756.745
R112 VTAIL.n84 VTAIL.n46 756.745
R113 VTAIL.n130 VTAIL.n92 756.745
R114 VTAIL.n310 VTAIL.n272 756.745
R115 VTAIL.n264 VTAIL.n226 756.745
R116 VTAIL.n220 VTAIL.n182 756.745
R117 VTAIL.n174 VTAIL.n136 756.745
R118 VTAIL.n331 VTAIL.n330 585
R119 VTAIL.n328 VTAIL.n327 585
R120 VTAIL.n337 VTAIL.n336 585
R121 VTAIL.n339 VTAIL.n338 585
R122 VTAIL.n324 VTAIL.n323 585
R123 VTAIL.n345 VTAIL.n344 585
R124 VTAIL.n347 VTAIL.n346 585
R125 VTAIL.n320 VTAIL.n319 585
R126 VTAIL.n353 VTAIL.n352 585
R127 VTAIL.n355 VTAIL.n354 585
R128 VTAIL.n17 VTAIL.n16 585
R129 VTAIL.n14 VTAIL.n13 585
R130 VTAIL.n23 VTAIL.n22 585
R131 VTAIL.n25 VTAIL.n24 585
R132 VTAIL.n10 VTAIL.n9 585
R133 VTAIL.n31 VTAIL.n30 585
R134 VTAIL.n33 VTAIL.n32 585
R135 VTAIL.n6 VTAIL.n5 585
R136 VTAIL.n39 VTAIL.n38 585
R137 VTAIL.n41 VTAIL.n40 585
R138 VTAIL.n61 VTAIL.n60 585
R139 VTAIL.n58 VTAIL.n57 585
R140 VTAIL.n67 VTAIL.n66 585
R141 VTAIL.n69 VTAIL.n68 585
R142 VTAIL.n54 VTAIL.n53 585
R143 VTAIL.n75 VTAIL.n74 585
R144 VTAIL.n77 VTAIL.n76 585
R145 VTAIL.n50 VTAIL.n49 585
R146 VTAIL.n83 VTAIL.n82 585
R147 VTAIL.n85 VTAIL.n84 585
R148 VTAIL.n107 VTAIL.n106 585
R149 VTAIL.n104 VTAIL.n103 585
R150 VTAIL.n113 VTAIL.n112 585
R151 VTAIL.n115 VTAIL.n114 585
R152 VTAIL.n100 VTAIL.n99 585
R153 VTAIL.n121 VTAIL.n120 585
R154 VTAIL.n123 VTAIL.n122 585
R155 VTAIL.n96 VTAIL.n95 585
R156 VTAIL.n129 VTAIL.n128 585
R157 VTAIL.n131 VTAIL.n130 585
R158 VTAIL.n311 VTAIL.n310 585
R159 VTAIL.n309 VTAIL.n308 585
R160 VTAIL.n276 VTAIL.n275 585
R161 VTAIL.n303 VTAIL.n302 585
R162 VTAIL.n301 VTAIL.n300 585
R163 VTAIL.n280 VTAIL.n279 585
R164 VTAIL.n295 VTAIL.n294 585
R165 VTAIL.n293 VTAIL.n292 585
R166 VTAIL.n284 VTAIL.n283 585
R167 VTAIL.n287 VTAIL.n286 585
R168 VTAIL.n265 VTAIL.n264 585
R169 VTAIL.n263 VTAIL.n262 585
R170 VTAIL.n230 VTAIL.n229 585
R171 VTAIL.n257 VTAIL.n256 585
R172 VTAIL.n255 VTAIL.n254 585
R173 VTAIL.n234 VTAIL.n233 585
R174 VTAIL.n249 VTAIL.n248 585
R175 VTAIL.n247 VTAIL.n246 585
R176 VTAIL.n238 VTAIL.n237 585
R177 VTAIL.n241 VTAIL.n240 585
R178 VTAIL.n221 VTAIL.n220 585
R179 VTAIL.n219 VTAIL.n218 585
R180 VTAIL.n186 VTAIL.n185 585
R181 VTAIL.n213 VTAIL.n212 585
R182 VTAIL.n211 VTAIL.n210 585
R183 VTAIL.n190 VTAIL.n189 585
R184 VTAIL.n205 VTAIL.n204 585
R185 VTAIL.n203 VTAIL.n202 585
R186 VTAIL.n194 VTAIL.n193 585
R187 VTAIL.n197 VTAIL.n196 585
R188 VTAIL.n175 VTAIL.n174 585
R189 VTAIL.n173 VTAIL.n172 585
R190 VTAIL.n140 VTAIL.n139 585
R191 VTAIL.n167 VTAIL.n166 585
R192 VTAIL.n165 VTAIL.n164 585
R193 VTAIL.n144 VTAIL.n143 585
R194 VTAIL.n159 VTAIL.n158 585
R195 VTAIL.n157 VTAIL.n156 585
R196 VTAIL.n148 VTAIL.n147 585
R197 VTAIL.n151 VTAIL.n150 585
R198 VTAIL.t10 VTAIL.n329 327.473
R199 VTAIL.t8 VTAIL.n15 327.473
R200 VTAIL.t5 VTAIL.n59 327.473
R201 VTAIL.t0 VTAIL.n105 327.473
R202 VTAIL.t1 VTAIL.n285 327.473
R203 VTAIL.t6 VTAIL.n239 327.473
R204 VTAIL.t15 VTAIL.n195 327.473
R205 VTAIL.t9 VTAIL.n149 327.473
R206 VTAIL.n330 VTAIL.n327 171.744
R207 VTAIL.n337 VTAIL.n327 171.744
R208 VTAIL.n338 VTAIL.n337 171.744
R209 VTAIL.n338 VTAIL.n323 171.744
R210 VTAIL.n345 VTAIL.n323 171.744
R211 VTAIL.n346 VTAIL.n345 171.744
R212 VTAIL.n346 VTAIL.n319 171.744
R213 VTAIL.n353 VTAIL.n319 171.744
R214 VTAIL.n354 VTAIL.n353 171.744
R215 VTAIL.n16 VTAIL.n13 171.744
R216 VTAIL.n23 VTAIL.n13 171.744
R217 VTAIL.n24 VTAIL.n23 171.744
R218 VTAIL.n24 VTAIL.n9 171.744
R219 VTAIL.n31 VTAIL.n9 171.744
R220 VTAIL.n32 VTAIL.n31 171.744
R221 VTAIL.n32 VTAIL.n5 171.744
R222 VTAIL.n39 VTAIL.n5 171.744
R223 VTAIL.n40 VTAIL.n39 171.744
R224 VTAIL.n60 VTAIL.n57 171.744
R225 VTAIL.n67 VTAIL.n57 171.744
R226 VTAIL.n68 VTAIL.n67 171.744
R227 VTAIL.n68 VTAIL.n53 171.744
R228 VTAIL.n75 VTAIL.n53 171.744
R229 VTAIL.n76 VTAIL.n75 171.744
R230 VTAIL.n76 VTAIL.n49 171.744
R231 VTAIL.n83 VTAIL.n49 171.744
R232 VTAIL.n84 VTAIL.n83 171.744
R233 VTAIL.n106 VTAIL.n103 171.744
R234 VTAIL.n113 VTAIL.n103 171.744
R235 VTAIL.n114 VTAIL.n113 171.744
R236 VTAIL.n114 VTAIL.n99 171.744
R237 VTAIL.n121 VTAIL.n99 171.744
R238 VTAIL.n122 VTAIL.n121 171.744
R239 VTAIL.n122 VTAIL.n95 171.744
R240 VTAIL.n129 VTAIL.n95 171.744
R241 VTAIL.n130 VTAIL.n129 171.744
R242 VTAIL.n310 VTAIL.n309 171.744
R243 VTAIL.n309 VTAIL.n275 171.744
R244 VTAIL.n302 VTAIL.n275 171.744
R245 VTAIL.n302 VTAIL.n301 171.744
R246 VTAIL.n301 VTAIL.n279 171.744
R247 VTAIL.n294 VTAIL.n279 171.744
R248 VTAIL.n294 VTAIL.n293 171.744
R249 VTAIL.n293 VTAIL.n283 171.744
R250 VTAIL.n286 VTAIL.n283 171.744
R251 VTAIL.n264 VTAIL.n263 171.744
R252 VTAIL.n263 VTAIL.n229 171.744
R253 VTAIL.n256 VTAIL.n229 171.744
R254 VTAIL.n256 VTAIL.n255 171.744
R255 VTAIL.n255 VTAIL.n233 171.744
R256 VTAIL.n248 VTAIL.n233 171.744
R257 VTAIL.n248 VTAIL.n247 171.744
R258 VTAIL.n247 VTAIL.n237 171.744
R259 VTAIL.n240 VTAIL.n237 171.744
R260 VTAIL.n220 VTAIL.n219 171.744
R261 VTAIL.n219 VTAIL.n185 171.744
R262 VTAIL.n212 VTAIL.n185 171.744
R263 VTAIL.n212 VTAIL.n211 171.744
R264 VTAIL.n211 VTAIL.n189 171.744
R265 VTAIL.n204 VTAIL.n189 171.744
R266 VTAIL.n204 VTAIL.n203 171.744
R267 VTAIL.n203 VTAIL.n193 171.744
R268 VTAIL.n196 VTAIL.n193 171.744
R269 VTAIL.n174 VTAIL.n173 171.744
R270 VTAIL.n173 VTAIL.n139 171.744
R271 VTAIL.n166 VTAIL.n139 171.744
R272 VTAIL.n166 VTAIL.n165 171.744
R273 VTAIL.n165 VTAIL.n143 171.744
R274 VTAIL.n158 VTAIL.n143 171.744
R275 VTAIL.n158 VTAIL.n157 171.744
R276 VTAIL.n157 VTAIL.n147 171.744
R277 VTAIL.n150 VTAIL.n147 171.744
R278 VTAIL.n330 VTAIL.t10 85.8723
R279 VTAIL.n16 VTAIL.t8 85.8723
R280 VTAIL.n60 VTAIL.t5 85.8723
R281 VTAIL.n106 VTAIL.t0 85.8723
R282 VTAIL.n286 VTAIL.t1 85.8723
R283 VTAIL.n240 VTAIL.t6 85.8723
R284 VTAIL.n196 VTAIL.t15 85.8723
R285 VTAIL.n150 VTAIL.t9 85.8723
R286 VTAIL.n271 VTAIL.n270 64.1688
R287 VTAIL.n181 VTAIL.n180 64.1688
R288 VTAIL.n1 VTAIL.n0 64.1686
R289 VTAIL.n91 VTAIL.n90 64.1686
R290 VTAIL.n359 VTAIL.n358 30.246
R291 VTAIL.n45 VTAIL.n44 30.246
R292 VTAIL.n89 VTAIL.n88 30.246
R293 VTAIL.n135 VTAIL.n134 30.246
R294 VTAIL.n315 VTAIL.n314 30.246
R295 VTAIL.n269 VTAIL.n268 30.246
R296 VTAIL.n225 VTAIL.n224 30.246
R297 VTAIL.n179 VTAIL.n178 30.246
R298 VTAIL.n359 VTAIL.n315 22.6341
R299 VTAIL.n179 VTAIL.n135 22.6341
R300 VTAIL.n331 VTAIL.n329 16.3894
R301 VTAIL.n17 VTAIL.n15 16.3894
R302 VTAIL.n61 VTAIL.n59 16.3894
R303 VTAIL.n107 VTAIL.n105 16.3894
R304 VTAIL.n287 VTAIL.n285 16.3894
R305 VTAIL.n241 VTAIL.n239 16.3894
R306 VTAIL.n197 VTAIL.n195 16.3894
R307 VTAIL.n151 VTAIL.n149 16.3894
R308 VTAIL.n332 VTAIL.n328 12.8005
R309 VTAIL.n18 VTAIL.n14 12.8005
R310 VTAIL.n62 VTAIL.n58 12.8005
R311 VTAIL.n108 VTAIL.n104 12.8005
R312 VTAIL.n288 VTAIL.n284 12.8005
R313 VTAIL.n242 VTAIL.n238 12.8005
R314 VTAIL.n198 VTAIL.n194 12.8005
R315 VTAIL.n152 VTAIL.n148 12.8005
R316 VTAIL.n336 VTAIL.n335 12.0247
R317 VTAIL.n22 VTAIL.n21 12.0247
R318 VTAIL.n66 VTAIL.n65 12.0247
R319 VTAIL.n112 VTAIL.n111 12.0247
R320 VTAIL.n292 VTAIL.n291 12.0247
R321 VTAIL.n246 VTAIL.n245 12.0247
R322 VTAIL.n202 VTAIL.n201 12.0247
R323 VTAIL.n156 VTAIL.n155 12.0247
R324 VTAIL.n339 VTAIL.n326 11.249
R325 VTAIL.n25 VTAIL.n12 11.249
R326 VTAIL.n69 VTAIL.n56 11.249
R327 VTAIL.n115 VTAIL.n102 11.249
R328 VTAIL.n295 VTAIL.n282 11.249
R329 VTAIL.n249 VTAIL.n236 11.249
R330 VTAIL.n205 VTAIL.n192 11.249
R331 VTAIL.n159 VTAIL.n146 11.249
R332 VTAIL.n340 VTAIL.n324 10.4732
R333 VTAIL.n26 VTAIL.n10 10.4732
R334 VTAIL.n70 VTAIL.n54 10.4732
R335 VTAIL.n116 VTAIL.n100 10.4732
R336 VTAIL.n296 VTAIL.n280 10.4732
R337 VTAIL.n250 VTAIL.n234 10.4732
R338 VTAIL.n206 VTAIL.n190 10.4732
R339 VTAIL.n160 VTAIL.n144 10.4732
R340 VTAIL.n344 VTAIL.n343 9.69747
R341 VTAIL.n30 VTAIL.n29 9.69747
R342 VTAIL.n74 VTAIL.n73 9.69747
R343 VTAIL.n120 VTAIL.n119 9.69747
R344 VTAIL.n300 VTAIL.n299 9.69747
R345 VTAIL.n254 VTAIL.n253 9.69747
R346 VTAIL.n210 VTAIL.n209 9.69747
R347 VTAIL.n164 VTAIL.n163 9.69747
R348 VTAIL.n358 VTAIL.n357 9.45567
R349 VTAIL.n44 VTAIL.n43 9.45567
R350 VTAIL.n88 VTAIL.n87 9.45567
R351 VTAIL.n134 VTAIL.n133 9.45567
R352 VTAIL.n314 VTAIL.n313 9.45567
R353 VTAIL.n268 VTAIL.n267 9.45567
R354 VTAIL.n224 VTAIL.n223 9.45567
R355 VTAIL.n178 VTAIL.n177 9.45567
R356 VTAIL.n318 VTAIL.n317 9.3005
R357 VTAIL.n357 VTAIL.n356 9.3005
R358 VTAIL.n349 VTAIL.n348 9.3005
R359 VTAIL.n322 VTAIL.n321 9.3005
R360 VTAIL.n343 VTAIL.n342 9.3005
R361 VTAIL.n341 VTAIL.n340 9.3005
R362 VTAIL.n326 VTAIL.n325 9.3005
R363 VTAIL.n335 VTAIL.n334 9.3005
R364 VTAIL.n333 VTAIL.n332 9.3005
R365 VTAIL.n351 VTAIL.n350 9.3005
R366 VTAIL.n4 VTAIL.n3 9.3005
R367 VTAIL.n43 VTAIL.n42 9.3005
R368 VTAIL.n35 VTAIL.n34 9.3005
R369 VTAIL.n8 VTAIL.n7 9.3005
R370 VTAIL.n29 VTAIL.n28 9.3005
R371 VTAIL.n27 VTAIL.n26 9.3005
R372 VTAIL.n12 VTAIL.n11 9.3005
R373 VTAIL.n21 VTAIL.n20 9.3005
R374 VTAIL.n19 VTAIL.n18 9.3005
R375 VTAIL.n37 VTAIL.n36 9.3005
R376 VTAIL.n48 VTAIL.n47 9.3005
R377 VTAIL.n87 VTAIL.n86 9.3005
R378 VTAIL.n79 VTAIL.n78 9.3005
R379 VTAIL.n52 VTAIL.n51 9.3005
R380 VTAIL.n73 VTAIL.n72 9.3005
R381 VTAIL.n71 VTAIL.n70 9.3005
R382 VTAIL.n56 VTAIL.n55 9.3005
R383 VTAIL.n65 VTAIL.n64 9.3005
R384 VTAIL.n63 VTAIL.n62 9.3005
R385 VTAIL.n81 VTAIL.n80 9.3005
R386 VTAIL.n94 VTAIL.n93 9.3005
R387 VTAIL.n133 VTAIL.n132 9.3005
R388 VTAIL.n125 VTAIL.n124 9.3005
R389 VTAIL.n98 VTAIL.n97 9.3005
R390 VTAIL.n119 VTAIL.n118 9.3005
R391 VTAIL.n117 VTAIL.n116 9.3005
R392 VTAIL.n102 VTAIL.n101 9.3005
R393 VTAIL.n111 VTAIL.n110 9.3005
R394 VTAIL.n109 VTAIL.n108 9.3005
R395 VTAIL.n127 VTAIL.n126 9.3005
R396 VTAIL.n274 VTAIL.n273 9.3005
R397 VTAIL.n307 VTAIL.n306 9.3005
R398 VTAIL.n305 VTAIL.n304 9.3005
R399 VTAIL.n278 VTAIL.n277 9.3005
R400 VTAIL.n299 VTAIL.n298 9.3005
R401 VTAIL.n297 VTAIL.n296 9.3005
R402 VTAIL.n282 VTAIL.n281 9.3005
R403 VTAIL.n291 VTAIL.n290 9.3005
R404 VTAIL.n289 VTAIL.n288 9.3005
R405 VTAIL.n313 VTAIL.n312 9.3005
R406 VTAIL.n267 VTAIL.n266 9.3005
R407 VTAIL.n228 VTAIL.n227 9.3005
R408 VTAIL.n261 VTAIL.n260 9.3005
R409 VTAIL.n259 VTAIL.n258 9.3005
R410 VTAIL.n232 VTAIL.n231 9.3005
R411 VTAIL.n253 VTAIL.n252 9.3005
R412 VTAIL.n251 VTAIL.n250 9.3005
R413 VTAIL.n236 VTAIL.n235 9.3005
R414 VTAIL.n245 VTAIL.n244 9.3005
R415 VTAIL.n243 VTAIL.n242 9.3005
R416 VTAIL.n223 VTAIL.n222 9.3005
R417 VTAIL.n184 VTAIL.n183 9.3005
R418 VTAIL.n217 VTAIL.n216 9.3005
R419 VTAIL.n215 VTAIL.n214 9.3005
R420 VTAIL.n188 VTAIL.n187 9.3005
R421 VTAIL.n209 VTAIL.n208 9.3005
R422 VTAIL.n207 VTAIL.n206 9.3005
R423 VTAIL.n192 VTAIL.n191 9.3005
R424 VTAIL.n201 VTAIL.n200 9.3005
R425 VTAIL.n199 VTAIL.n198 9.3005
R426 VTAIL.n177 VTAIL.n176 9.3005
R427 VTAIL.n138 VTAIL.n137 9.3005
R428 VTAIL.n171 VTAIL.n170 9.3005
R429 VTAIL.n169 VTAIL.n168 9.3005
R430 VTAIL.n142 VTAIL.n141 9.3005
R431 VTAIL.n163 VTAIL.n162 9.3005
R432 VTAIL.n161 VTAIL.n160 9.3005
R433 VTAIL.n146 VTAIL.n145 9.3005
R434 VTAIL.n155 VTAIL.n154 9.3005
R435 VTAIL.n153 VTAIL.n152 9.3005
R436 VTAIL.n347 VTAIL.n322 8.92171
R437 VTAIL.n33 VTAIL.n8 8.92171
R438 VTAIL.n77 VTAIL.n52 8.92171
R439 VTAIL.n123 VTAIL.n98 8.92171
R440 VTAIL.n303 VTAIL.n278 8.92171
R441 VTAIL.n257 VTAIL.n232 8.92171
R442 VTAIL.n213 VTAIL.n188 8.92171
R443 VTAIL.n167 VTAIL.n142 8.92171
R444 VTAIL.n348 VTAIL.n320 8.14595
R445 VTAIL.n358 VTAIL.n316 8.14595
R446 VTAIL.n34 VTAIL.n6 8.14595
R447 VTAIL.n44 VTAIL.n2 8.14595
R448 VTAIL.n78 VTAIL.n50 8.14595
R449 VTAIL.n88 VTAIL.n46 8.14595
R450 VTAIL.n124 VTAIL.n96 8.14595
R451 VTAIL.n134 VTAIL.n92 8.14595
R452 VTAIL.n314 VTAIL.n272 8.14595
R453 VTAIL.n304 VTAIL.n276 8.14595
R454 VTAIL.n268 VTAIL.n226 8.14595
R455 VTAIL.n258 VTAIL.n230 8.14595
R456 VTAIL.n224 VTAIL.n182 8.14595
R457 VTAIL.n214 VTAIL.n186 8.14595
R458 VTAIL.n178 VTAIL.n136 8.14595
R459 VTAIL.n168 VTAIL.n140 8.14595
R460 VTAIL.n352 VTAIL.n351 7.3702
R461 VTAIL.n356 VTAIL.n355 7.3702
R462 VTAIL.n38 VTAIL.n37 7.3702
R463 VTAIL.n42 VTAIL.n41 7.3702
R464 VTAIL.n82 VTAIL.n81 7.3702
R465 VTAIL.n86 VTAIL.n85 7.3702
R466 VTAIL.n128 VTAIL.n127 7.3702
R467 VTAIL.n132 VTAIL.n131 7.3702
R468 VTAIL.n312 VTAIL.n311 7.3702
R469 VTAIL.n308 VTAIL.n307 7.3702
R470 VTAIL.n266 VTAIL.n265 7.3702
R471 VTAIL.n262 VTAIL.n261 7.3702
R472 VTAIL.n222 VTAIL.n221 7.3702
R473 VTAIL.n218 VTAIL.n217 7.3702
R474 VTAIL.n176 VTAIL.n175 7.3702
R475 VTAIL.n172 VTAIL.n171 7.3702
R476 VTAIL.n352 VTAIL.n318 6.59444
R477 VTAIL.n355 VTAIL.n318 6.59444
R478 VTAIL.n38 VTAIL.n4 6.59444
R479 VTAIL.n41 VTAIL.n4 6.59444
R480 VTAIL.n82 VTAIL.n48 6.59444
R481 VTAIL.n85 VTAIL.n48 6.59444
R482 VTAIL.n128 VTAIL.n94 6.59444
R483 VTAIL.n131 VTAIL.n94 6.59444
R484 VTAIL.n311 VTAIL.n274 6.59444
R485 VTAIL.n308 VTAIL.n274 6.59444
R486 VTAIL.n265 VTAIL.n228 6.59444
R487 VTAIL.n262 VTAIL.n228 6.59444
R488 VTAIL.n221 VTAIL.n184 6.59444
R489 VTAIL.n218 VTAIL.n184 6.59444
R490 VTAIL.n175 VTAIL.n138 6.59444
R491 VTAIL.n172 VTAIL.n138 6.59444
R492 VTAIL.n351 VTAIL.n320 5.81868
R493 VTAIL.n356 VTAIL.n316 5.81868
R494 VTAIL.n37 VTAIL.n6 5.81868
R495 VTAIL.n42 VTAIL.n2 5.81868
R496 VTAIL.n81 VTAIL.n50 5.81868
R497 VTAIL.n86 VTAIL.n46 5.81868
R498 VTAIL.n127 VTAIL.n96 5.81868
R499 VTAIL.n132 VTAIL.n92 5.81868
R500 VTAIL.n312 VTAIL.n272 5.81868
R501 VTAIL.n307 VTAIL.n276 5.81868
R502 VTAIL.n266 VTAIL.n226 5.81868
R503 VTAIL.n261 VTAIL.n230 5.81868
R504 VTAIL.n222 VTAIL.n182 5.81868
R505 VTAIL.n217 VTAIL.n186 5.81868
R506 VTAIL.n176 VTAIL.n136 5.81868
R507 VTAIL.n171 VTAIL.n140 5.81868
R508 VTAIL.n348 VTAIL.n347 5.04292
R509 VTAIL.n34 VTAIL.n33 5.04292
R510 VTAIL.n78 VTAIL.n77 5.04292
R511 VTAIL.n124 VTAIL.n123 5.04292
R512 VTAIL.n304 VTAIL.n303 5.04292
R513 VTAIL.n258 VTAIL.n257 5.04292
R514 VTAIL.n214 VTAIL.n213 5.04292
R515 VTAIL.n168 VTAIL.n167 5.04292
R516 VTAIL.n344 VTAIL.n322 4.26717
R517 VTAIL.n30 VTAIL.n8 4.26717
R518 VTAIL.n74 VTAIL.n52 4.26717
R519 VTAIL.n120 VTAIL.n98 4.26717
R520 VTAIL.n300 VTAIL.n278 4.26717
R521 VTAIL.n254 VTAIL.n232 4.26717
R522 VTAIL.n210 VTAIL.n188 4.26717
R523 VTAIL.n164 VTAIL.n142 4.26717
R524 VTAIL.n0 VTAIL.t14 4.03338
R525 VTAIL.n0 VTAIL.t12 4.03338
R526 VTAIL.n90 VTAIL.t4 4.03338
R527 VTAIL.n90 VTAIL.t7 4.03338
R528 VTAIL.n270 VTAIL.t2 4.03338
R529 VTAIL.n270 VTAIL.t3 4.03338
R530 VTAIL.n180 VTAIL.t13 4.03338
R531 VTAIL.n180 VTAIL.t11 4.03338
R532 VTAIL.n333 VTAIL.n329 3.70995
R533 VTAIL.n19 VTAIL.n15 3.70995
R534 VTAIL.n63 VTAIL.n59 3.70995
R535 VTAIL.n109 VTAIL.n105 3.70995
R536 VTAIL.n243 VTAIL.n239 3.70995
R537 VTAIL.n199 VTAIL.n195 3.70995
R538 VTAIL.n153 VTAIL.n149 3.70995
R539 VTAIL.n289 VTAIL.n285 3.70995
R540 VTAIL.n343 VTAIL.n324 3.49141
R541 VTAIL.n29 VTAIL.n10 3.49141
R542 VTAIL.n73 VTAIL.n54 3.49141
R543 VTAIL.n119 VTAIL.n100 3.49141
R544 VTAIL.n299 VTAIL.n280 3.49141
R545 VTAIL.n253 VTAIL.n234 3.49141
R546 VTAIL.n209 VTAIL.n190 3.49141
R547 VTAIL.n163 VTAIL.n144 3.49141
R548 VTAIL.n181 VTAIL.n179 3.31947
R549 VTAIL.n225 VTAIL.n181 3.31947
R550 VTAIL.n271 VTAIL.n269 3.31947
R551 VTAIL.n315 VTAIL.n271 3.31947
R552 VTAIL.n135 VTAIL.n91 3.31947
R553 VTAIL.n91 VTAIL.n89 3.31947
R554 VTAIL.n45 VTAIL.n1 3.31947
R555 VTAIL VTAIL.n359 3.26128
R556 VTAIL.n340 VTAIL.n339 2.71565
R557 VTAIL.n26 VTAIL.n25 2.71565
R558 VTAIL.n70 VTAIL.n69 2.71565
R559 VTAIL.n116 VTAIL.n115 2.71565
R560 VTAIL.n296 VTAIL.n295 2.71565
R561 VTAIL.n250 VTAIL.n249 2.71565
R562 VTAIL.n206 VTAIL.n205 2.71565
R563 VTAIL.n160 VTAIL.n159 2.71565
R564 VTAIL.n336 VTAIL.n326 1.93989
R565 VTAIL.n22 VTAIL.n12 1.93989
R566 VTAIL.n66 VTAIL.n56 1.93989
R567 VTAIL.n112 VTAIL.n102 1.93989
R568 VTAIL.n292 VTAIL.n282 1.93989
R569 VTAIL.n246 VTAIL.n236 1.93989
R570 VTAIL.n202 VTAIL.n192 1.93989
R571 VTAIL.n156 VTAIL.n146 1.93989
R572 VTAIL.n335 VTAIL.n328 1.16414
R573 VTAIL.n21 VTAIL.n14 1.16414
R574 VTAIL.n65 VTAIL.n58 1.16414
R575 VTAIL.n111 VTAIL.n104 1.16414
R576 VTAIL.n291 VTAIL.n284 1.16414
R577 VTAIL.n245 VTAIL.n238 1.16414
R578 VTAIL.n201 VTAIL.n194 1.16414
R579 VTAIL.n155 VTAIL.n148 1.16414
R580 VTAIL.n269 VTAIL.n225 0.470328
R581 VTAIL.n89 VTAIL.n45 0.470328
R582 VTAIL.n332 VTAIL.n331 0.388379
R583 VTAIL.n18 VTAIL.n17 0.388379
R584 VTAIL.n62 VTAIL.n61 0.388379
R585 VTAIL.n108 VTAIL.n107 0.388379
R586 VTAIL.n288 VTAIL.n287 0.388379
R587 VTAIL.n242 VTAIL.n241 0.388379
R588 VTAIL.n198 VTAIL.n197 0.388379
R589 VTAIL.n152 VTAIL.n151 0.388379
R590 VTAIL.n334 VTAIL.n333 0.155672
R591 VTAIL.n334 VTAIL.n325 0.155672
R592 VTAIL.n341 VTAIL.n325 0.155672
R593 VTAIL.n342 VTAIL.n341 0.155672
R594 VTAIL.n342 VTAIL.n321 0.155672
R595 VTAIL.n349 VTAIL.n321 0.155672
R596 VTAIL.n350 VTAIL.n349 0.155672
R597 VTAIL.n350 VTAIL.n317 0.155672
R598 VTAIL.n357 VTAIL.n317 0.155672
R599 VTAIL.n20 VTAIL.n19 0.155672
R600 VTAIL.n20 VTAIL.n11 0.155672
R601 VTAIL.n27 VTAIL.n11 0.155672
R602 VTAIL.n28 VTAIL.n27 0.155672
R603 VTAIL.n28 VTAIL.n7 0.155672
R604 VTAIL.n35 VTAIL.n7 0.155672
R605 VTAIL.n36 VTAIL.n35 0.155672
R606 VTAIL.n36 VTAIL.n3 0.155672
R607 VTAIL.n43 VTAIL.n3 0.155672
R608 VTAIL.n64 VTAIL.n63 0.155672
R609 VTAIL.n64 VTAIL.n55 0.155672
R610 VTAIL.n71 VTAIL.n55 0.155672
R611 VTAIL.n72 VTAIL.n71 0.155672
R612 VTAIL.n72 VTAIL.n51 0.155672
R613 VTAIL.n79 VTAIL.n51 0.155672
R614 VTAIL.n80 VTAIL.n79 0.155672
R615 VTAIL.n80 VTAIL.n47 0.155672
R616 VTAIL.n87 VTAIL.n47 0.155672
R617 VTAIL.n110 VTAIL.n109 0.155672
R618 VTAIL.n110 VTAIL.n101 0.155672
R619 VTAIL.n117 VTAIL.n101 0.155672
R620 VTAIL.n118 VTAIL.n117 0.155672
R621 VTAIL.n118 VTAIL.n97 0.155672
R622 VTAIL.n125 VTAIL.n97 0.155672
R623 VTAIL.n126 VTAIL.n125 0.155672
R624 VTAIL.n126 VTAIL.n93 0.155672
R625 VTAIL.n133 VTAIL.n93 0.155672
R626 VTAIL.n313 VTAIL.n273 0.155672
R627 VTAIL.n306 VTAIL.n273 0.155672
R628 VTAIL.n306 VTAIL.n305 0.155672
R629 VTAIL.n305 VTAIL.n277 0.155672
R630 VTAIL.n298 VTAIL.n277 0.155672
R631 VTAIL.n298 VTAIL.n297 0.155672
R632 VTAIL.n297 VTAIL.n281 0.155672
R633 VTAIL.n290 VTAIL.n281 0.155672
R634 VTAIL.n290 VTAIL.n289 0.155672
R635 VTAIL.n267 VTAIL.n227 0.155672
R636 VTAIL.n260 VTAIL.n227 0.155672
R637 VTAIL.n260 VTAIL.n259 0.155672
R638 VTAIL.n259 VTAIL.n231 0.155672
R639 VTAIL.n252 VTAIL.n231 0.155672
R640 VTAIL.n252 VTAIL.n251 0.155672
R641 VTAIL.n251 VTAIL.n235 0.155672
R642 VTAIL.n244 VTAIL.n235 0.155672
R643 VTAIL.n244 VTAIL.n243 0.155672
R644 VTAIL.n223 VTAIL.n183 0.155672
R645 VTAIL.n216 VTAIL.n183 0.155672
R646 VTAIL.n216 VTAIL.n215 0.155672
R647 VTAIL.n215 VTAIL.n187 0.155672
R648 VTAIL.n208 VTAIL.n187 0.155672
R649 VTAIL.n208 VTAIL.n207 0.155672
R650 VTAIL.n207 VTAIL.n191 0.155672
R651 VTAIL.n200 VTAIL.n191 0.155672
R652 VTAIL.n200 VTAIL.n199 0.155672
R653 VTAIL.n177 VTAIL.n137 0.155672
R654 VTAIL.n170 VTAIL.n137 0.155672
R655 VTAIL.n170 VTAIL.n169 0.155672
R656 VTAIL.n169 VTAIL.n141 0.155672
R657 VTAIL.n162 VTAIL.n141 0.155672
R658 VTAIL.n162 VTAIL.n161 0.155672
R659 VTAIL.n161 VTAIL.n145 0.155672
R660 VTAIL.n154 VTAIL.n145 0.155672
R661 VTAIL.n154 VTAIL.n153 0.155672
R662 VTAIL VTAIL.n1 0.0586897
R663 VDD2.n2 VDD2.n1 82.4515
R664 VDD2.n2 VDD2.n0 82.4515
R665 VDD2 VDD2.n5 82.4489
R666 VDD2.n4 VDD2.n3 80.8476
R667 VDD2.n4 VDD2.n2 45.5989
R668 VDD2.n5 VDD2.t0 4.03338
R669 VDD2.n5 VDD2.t3 4.03338
R670 VDD2.n3 VDD2.t6 4.03338
R671 VDD2.n3 VDD2.t7 4.03338
R672 VDD2.n1 VDD2.t4 4.03338
R673 VDD2.n1 VDD2.t5 4.03338
R674 VDD2.n0 VDD2.t1 4.03338
R675 VDD2.n0 VDD2.t2 4.03338
R676 VDD2 VDD2.n4 1.71817
R677 VP.n24 VP.n23 161.3
R678 VP.n25 VP.n20 161.3
R679 VP.n27 VP.n26 161.3
R680 VP.n28 VP.n19 161.3
R681 VP.n30 VP.n29 161.3
R682 VP.n31 VP.n18 161.3
R683 VP.n34 VP.n33 161.3
R684 VP.n35 VP.n17 161.3
R685 VP.n37 VP.n36 161.3
R686 VP.n38 VP.n16 161.3
R687 VP.n40 VP.n39 161.3
R688 VP.n41 VP.n15 161.3
R689 VP.n43 VP.n42 161.3
R690 VP.n44 VP.n14 161.3
R691 VP.n46 VP.n45 161.3
R692 VP.n85 VP.n84 161.3
R693 VP.n83 VP.n1 161.3
R694 VP.n82 VP.n81 161.3
R695 VP.n80 VP.n2 161.3
R696 VP.n79 VP.n78 161.3
R697 VP.n77 VP.n3 161.3
R698 VP.n76 VP.n75 161.3
R699 VP.n74 VP.n4 161.3
R700 VP.n73 VP.n72 161.3
R701 VP.n70 VP.n5 161.3
R702 VP.n69 VP.n68 161.3
R703 VP.n67 VP.n6 161.3
R704 VP.n66 VP.n65 161.3
R705 VP.n64 VP.n7 161.3
R706 VP.n63 VP.n62 161.3
R707 VP.n61 VP.n60 161.3
R708 VP.n59 VP.n9 161.3
R709 VP.n58 VP.n57 161.3
R710 VP.n56 VP.n10 161.3
R711 VP.n55 VP.n54 161.3
R712 VP.n53 VP.n11 161.3
R713 VP.n52 VP.n51 161.3
R714 VP.n50 VP.n12 161.3
R715 VP.n22 VP.t7 88.9803
R716 VP.n49 VP.n48 76.5021
R717 VP.n86 VP.n0 76.5021
R718 VP.n47 VP.n13 76.5021
R719 VP.n48 VP.t5 55.184
R720 VP.n8 VP.t6 55.184
R721 VP.n71 VP.t4 55.184
R722 VP.n0 VP.t3 55.184
R723 VP.n13 VP.t1 55.184
R724 VP.n32 VP.t0 55.184
R725 VP.n21 VP.t2 55.184
R726 VP.n54 VP.n10 55.0167
R727 VP.n78 VP.n2 55.0167
R728 VP.n39 VP.n15 55.0167
R729 VP.n22 VP.n21 53.7745
R730 VP.n49 VP.n47 52.3627
R731 VP.n65 VP.n6 40.4106
R732 VP.n69 VP.n6 40.4106
R733 VP.n30 VP.n19 40.4106
R734 VP.n26 VP.n19 40.4106
R735 VP.n54 VP.n53 25.8045
R736 VP.n82 VP.n2 25.8045
R737 VP.n43 VP.n15 25.8045
R738 VP.n52 VP.n12 24.3439
R739 VP.n53 VP.n52 24.3439
R740 VP.n58 VP.n10 24.3439
R741 VP.n59 VP.n58 24.3439
R742 VP.n60 VP.n59 24.3439
R743 VP.n64 VP.n63 24.3439
R744 VP.n65 VP.n64 24.3439
R745 VP.n70 VP.n69 24.3439
R746 VP.n72 VP.n70 24.3439
R747 VP.n76 VP.n4 24.3439
R748 VP.n77 VP.n76 24.3439
R749 VP.n78 VP.n77 24.3439
R750 VP.n83 VP.n82 24.3439
R751 VP.n84 VP.n83 24.3439
R752 VP.n44 VP.n43 24.3439
R753 VP.n45 VP.n44 24.3439
R754 VP.n31 VP.n30 24.3439
R755 VP.n33 VP.n31 24.3439
R756 VP.n37 VP.n17 24.3439
R757 VP.n38 VP.n37 24.3439
R758 VP.n39 VP.n38 24.3439
R759 VP.n25 VP.n24 24.3439
R760 VP.n26 VP.n25 24.3439
R761 VP.n63 VP.n8 20.6924
R762 VP.n72 VP.n71 20.6924
R763 VP.n33 VP.n32 20.6924
R764 VP.n24 VP.n21 20.6924
R765 VP.n48 VP.n12 13.3894
R766 VP.n84 VP.n0 13.3894
R767 VP.n45 VP.n13 13.3894
R768 VP.n60 VP.n8 3.65202
R769 VP.n71 VP.n4 3.65202
R770 VP.n32 VP.n17 3.65202
R771 VP.n23 VP.n22 3.05396
R772 VP.n47 VP.n46 0.355081
R773 VP.n50 VP.n49 0.355081
R774 VP.n86 VP.n85 0.355081
R775 VP VP.n86 0.26685
R776 VP.n23 VP.n20 0.189894
R777 VP.n27 VP.n20 0.189894
R778 VP.n28 VP.n27 0.189894
R779 VP.n29 VP.n28 0.189894
R780 VP.n29 VP.n18 0.189894
R781 VP.n34 VP.n18 0.189894
R782 VP.n35 VP.n34 0.189894
R783 VP.n36 VP.n35 0.189894
R784 VP.n36 VP.n16 0.189894
R785 VP.n40 VP.n16 0.189894
R786 VP.n41 VP.n40 0.189894
R787 VP.n42 VP.n41 0.189894
R788 VP.n42 VP.n14 0.189894
R789 VP.n46 VP.n14 0.189894
R790 VP.n51 VP.n50 0.189894
R791 VP.n51 VP.n11 0.189894
R792 VP.n55 VP.n11 0.189894
R793 VP.n56 VP.n55 0.189894
R794 VP.n57 VP.n56 0.189894
R795 VP.n57 VP.n9 0.189894
R796 VP.n61 VP.n9 0.189894
R797 VP.n62 VP.n61 0.189894
R798 VP.n62 VP.n7 0.189894
R799 VP.n66 VP.n7 0.189894
R800 VP.n67 VP.n66 0.189894
R801 VP.n68 VP.n67 0.189894
R802 VP.n68 VP.n5 0.189894
R803 VP.n73 VP.n5 0.189894
R804 VP.n74 VP.n73 0.189894
R805 VP.n75 VP.n74 0.189894
R806 VP.n75 VP.n3 0.189894
R807 VP.n79 VP.n3 0.189894
R808 VP.n80 VP.n79 0.189894
R809 VP.n81 VP.n80 0.189894
R810 VP.n81 VP.n1 0.189894
R811 VP.n85 VP.n1 0.189894
R812 VDD1 VDD1.n0 82.5652
R813 VDD1.n3 VDD1.n2 82.4515
R814 VDD1.n3 VDD1.n1 82.4515
R815 VDD1.n5 VDD1.n4 80.8476
R816 VDD1.n5 VDD1.n3 46.1819
R817 VDD1.n4 VDD1.t7 4.03338
R818 VDD1.n4 VDD1.t6 4.03338
R819 VDD1.n0 VDD1.t0 4.03338
R820 VDD1.n0 VDD1.t5 4.03338
R821 VDD1.n2 VDD1.t3 4.03338
R822 VDD1.n2 VDD1.t4 4.03338
R823 VDD1.n1 VDD1.t2 4.03338
R824 VDD1.n1 VDD1.t1 4.03338
R825 VDD1 VDD1.n5 1.60179
R826 B.n410 B.n409 585
R827 B.n408 B.n139 585
R828 B.n407 B.n406 585
R829 B.n405 B.n140 585
R830 B.n404 B.n403 585
R831 B.n402 B.n141 585
R832 B.n401 B.n400 585
R833 B.n399 B.n142 585
R834 B.n398 B.n397 585
R835 B.n396 B.n143 585
R836 B.n395 B.n394 585
R837 B.n393 B.n144 585
R838 B.n392 B.n391 585
R839 B.n390 B.n145 585
R840 B.n389 B.n388 585
R841 B.n387 B.n146 585
R842 B.n386 B.n385 585
R843 B.n384 B.n147 585
R844 B.n383 B.n382 585
R845 B.n381 B.n148 585
R846 B.n380 B.n379 585
R847 B.n378 B.n149 585
R848 B.n377 B.n376 585
R849 B.n375 B.n150 585
R850 B.n374 B.n373 585
R851 B.n372 B.n151 585
R852 B.n371 B.n370 585
R853 B.n369 B.n152 585
R854 B.n368 B.n367 585
R855 B.n366 B.n153 585
R856 B.n364 B.n363 585
R857 B.n362 B.n156 585
R858 B.n361 B.n360 585
R859 B.n359 B.n157 585
R860 B.n358 B.n357 585
R861 B.n356 B.n158 585
R862 B.n355 B.n354 585
R863 B.n353 B.n159 585
R864 B.n352 B.n351 585
R865 B.n350 B.n160 585
R866 B.n349 B.n348 585
R867 B.n344 B.n161 585
R868 B.n343 B.n342 585
R869 B.n341 B.n162 585
R870 B.n340 B.n339 585
R871 B.n338 B.n163 585
R872 B.n337 B.n336 585
R873 B.n335 B.n164 585
R874 B.n334 B.n333 585
R875 B.n332 B.n165 585
R876 B.n331 B.n330 585
R877 B.n329 B.n166 585
R878 B.n328 B.n327 585
R879 B.n326 B.n167 585
R880 B.n325 B.n324 585
R881 B.n323 B.n168 585
R882 B.n322 B.n321 585
R883 B.n320 B.n169 585
R884 B.n319 B.n318 585
R885 B.n317 B.n170 585
R886 B.n316 B.n315 585
R887 B.n314 B.n171 585
R888 B.n313 B.n312 585
R889 B.n311 B.n172 585
R890 B.n310 B.n309 585
R891 B.n308 B.n173 585
R892 B.n307 B.n306 585
R893 B.n305 B.n174 585
R894 B.n304 B.n303 585
R895 B.n302 B.n175 585
R896 B.n411 B.n138 585
R897 B.n413 B.n412 585
R898 B.n414 B.n137 585
R899 B.n416 B.n415 585
R900 B.n417 B.n136 585
R901 B.n419 B.n418 585
R902 B.n420 B.n135 585
R903 B.n422 B.n421 585
R904 B.n423 B.n134 585
R905 B.n425 B.n424 585
R906 B.n426 B.n133 585
R907 B.n428 B.n427 585
R908 B.n429 B.n132 585
R909 B.n431 B.n430 585
R910 B.n432 B.n131 585
R911 B.n434 B.n433 585
R912 B.n435 B.n130 585
R913 B.n437 B.n436 585
R914 B.n438 B.n129 585
R915 B.n440 B.n439 585
R916 B.n441 B.n128 585
R917 B.n443 B.n442 585
R918 B.n444 B.n127 585
R919 B.n446 B.n445 585
R920 B.n447 B.n126 585
R921 B.n449 B.n448 585
R922 B.n450 B.n125 585
R923 B.n452 B.n451 585
R924 B.n453 B.n124 585
R925 B.n455 B.n454 585
R926 B.n456 B.n123 585
R927 B.n458 B.n457 585
R928 B.n459 B.n122 585
R929 B.n461 B.n460 585
R930 B.n462 B.n121 585
R931 B.n464 B.n463 585
R932 B.n465 B.n120 585
R933 B.n467 B.n466 585
R934 B.n468 B.n119 585
R935 B.n470 B.n469 585
R936 B.n471 B.n118 585
R937 B.n473 B.n472 585
R938 B.n474 B.n117 585
R939 B.n476 B.n475 585
R940 B.n477 B.n116 585
R941 B.n479 B.n478 585
R942 B.n480 B.n115 585
R943 B.n482 B.n481 585
R944 B.n483 B.n114 585
R945 B.n485 B.n484 585
R946 B.n486 B.n113 585
R947 B.n488 B.n487 585
R948 B.n489 B.n112 585
R949 B.n491 B.n490 585
R950 B.n492 B.n111 585
R951 B.n494 B.n493 585
R952 B.n495 B.n110 585
R953 B.n497 B.n496 585
R954 B.n498 B.n109 585
R955 B.n500 B.n499 585
R956 B.n501 B.n108 585
R957 B.n503 B.n502 585
R958 B.n504 B.n107 585
R959 B.n506 B.n505 585
R960 B.n507 B.n106 585
R961 B.n509 B.n508 585
R962 B.n510 B.n105 585
R963 B.n512 B.n511 585
R964 B.n513 B.n104 585
R965 B.n515 B.n514 585
R966 B.n516 B.n103 585
R967 B.n518 B.n517 585
R968 B.n519 B.n102 585
R969 B.n521 B.n520 585
R970 B.n522 B.n101 585
R971 B.n524 B.n523 585
R972 B.n525 B.n100 585
R973 B.n527 B.n526 585
R974 B.n528 B.n99 585
R975 B.n530 B.n529 585
R976 B.n531 B.n98 585
R977 B.n533 B.n532 585
R978 B.n534 B.n97 585
R979 B.n536 B.n535 585
R980 B.n537 B.n96 585
R981 B.n539 B.n538 585
R982 B.n540 B.n95 585
R983 B.n542 B.n541 585
R984 B.n543 B.n94 585
R985 B.n545 B.n544 585
R986 B.n546 B.n93 585
R987 B.n548 B.n547 585
R988 B.n549 B.n92 585
R989 B.n551 B.n550 585
R990 B.n552 B.n91 585
R991 B.n554 B.n553 585
R992 B.n555 B.n90 585
R993 B.n557 B.n556 585
R994 B.n558 B.n89 585
R995 B.n560 B.n559 585
R996 B.n561 B.n88 585
R997 B.n563 B.n562 585
R998 B.n564 B.n87 585
R999 B.n566 B.n565 585
R1000 B.n567 B.n86 585
R1001 B.n569 B.n568 585
R1002 B.n570 B.n85 585
R1003 B.n572 B.n571 585
R1004 B.n573 B.n84 585
R1005 B.n575 B.n574 585
R1006 B.n576 B.n83 585
R1007 B.n578 B.n577 585
R1008 B.n579 B.n82 585
R1009 B.n581 B.n580 585
R1010 B.n582 B.n81 585
R1011 B.n584 B.n583 585
R1012 B.n585 B.n80 585
R1013 B.n587 B.n586 585
R1014 B.n588 B.n79 585
R1015 B.n590 B.n589 585
R1016 B.n591 B.n78 585
R1017 B.n593 B.n592 585
R1018 B.n594 B.n77 585
R1019 B.n596 B.n595 585
R1020 B.n597 B.n76 585
R1021 B.n599 B.n598 585
R1022 B.n600 B.n75 585
R1023 B.n602 B.n601 585
R1024 B.n603 B.n74 585
R1025 B.n605 B.n604 585
R1026 B.n711 B.n34 585
R1027 B.n710 B.n709 585
R1028 B.n708 B.n35 585
R1029 B.n707 B.n706 585
R1030 B.n705 B.n36 585
R1031 B.n704 B.n703 585
R1032 B.n702 B.n37 585
R1033 B.n701 B.n700 585
R1034 B.n699 B.n38 585
R1035 B.n698 B.n697 585
R1036 B.n696 B.n39 585
R1037 B.n695 B.n694 585
R1038 B.n693 B.n40 585
R1039 B.n692 B.n691 585
R1040 B.n690 B.n41 585
R1041 B.n689 B.n688 585
R1042 B.n687 B.n42 585
R1043 B.n686 B.n685 585
R1044 B.n684 B.n43 585
R1045 B.n683 B.n682 585
R1046 B.n681 B.n44 585
R1047 B.n680 B.n679 585
R1048 B.n678 B.n45 585
R1049 B.n677 B.n676 585
R1050 B.n675 B.n46 585
R1051 B.n674 B.n673 585
R1052 B.n672 B.n47 585
R1053 B.n671 B.n670 585
R1054 B.n669 B.n48 585
R1055 B.n668 B.n667 585
R1056 B.n665 B.n49 585
R1057 B.n664 B.n663 585
R1058 B.n662 B.n52 585
R1059 B.n661 B.n660 585
R1060 B.n659 B.n53 585
R1061 B.n658 B.n657 585
R1062 B.n656 B.n54 585
R1063 B.n655 B.n654 585
R1064 B.n653 B.n55 585
R1065 B.n652 B.n651 585
R1066 B.n650 B.n649 585
R1067 B.n648 B.n59 585
R1068 B.n647 B.n646 585
R1069 B.n645 B.n60 585
R1070 B.n644 B.n643 585
R1071 B.n642 B.n61 585
R1072 B.n641 B.n640 585
R1073 B.n639 B.n62 585
R1074 B.n638 B.n637 585
R1075 B.n636 B.n63 585
R1076 B.n635 B.n634 585
R1077 B.n633 B.n64 585
R1078 B.n632 B.n631 585
R1079 B.n630 B.n65 585
R1080 B.n629 B.n628 585
R1081 B.n627 B.n66 585
R1082 B.n626 B.n625 585
R1083 B.n624 B.n67 585
R1084 B.n623 B.n622 585
R1085 B.n621 B.n68 585
R1086 B.n620 B.n619 585
R1087 B.n618 B.n69 585
R1088 B.n617 B.n616 585
R1089 B.n615 B.n70 585
R1090 B.n614 B.n613 585
R1091 B.n612 B.n71 585
R1092 B.n611 B.n610 585
R1093 B.n609 B.n72 585
R1094 B.n608 B.n607 585
R1095 B.n606 B.n73 585
R1096 B.n713 B.n712 585
R1097 B.n714 B.n33 585
R1098 B.n716 B.n715 585
R1099 B.n717 B.n32 585
R1100 B.n719 B.n718 585
R1101 B.n720 B.n31 585
R1102 B.n722 B.n721 585
R1103 B.n723 B.n30 585
R1104 B.n725 B.n724 585
R1105 B.n726 B.n29 585
R1106 B.n728 B.n727 585
R1107 B.n729 B.n28 585
R1108 B.n731 B.n730 585
R1109 B.n732 B.n27 585
R1110 B.n734 B.n733 585
R1111 B.n735 B.n26 585
R1112 B.n737 B.n736 585
R1113 B.n738 B.n25 585
R1114 B.n740 B.n739 585
R1115 B.n741 B.n24 585
R1116 B.n743 B.n742 585
R1117 B.n744 B.n23 585
R1118 B.n746 B.n745 585
R1119 B.n747 B.n22 585
R1120 B.n749 B.n748 585
R1121 B.n750 B.n21 585
R1122 B.n752 B.n751 585
R1123 B.n753 B.n20 585
R1124 B.n755 B.n754 585
R1125 B.n756 B.n19 585
R1126 B.n758 B.n757 585
R1127 B.n759 B.n18 585
R1128 B.n761 B.n760 585
R1129 B.n762 B.n17 585
R1130 B.n764 B.n763 585
R1131 B.n765 B.n16 585
R1132 B.n767 B.n766 585
R1133 B.n768 B.n15 585
R1134 B.n770 B.n769 585
R1135 B.n771 B.n14 585
R1136 B.n773 B.n772 585
R1137 B.n774 B.n13 585
R1138 B.n776 B.n775 585
R1139 B.n777 B.n12 585
R1140 B.n779 B.n778 585
R1141 B.n780 B.n11 585
R1142 B.n782 B.n781 585
R1143 B.n783 B.n10 585
R1144 B.n785 B.n784 585
R1145 B.n786 B.n9 585
R1146 B.n788 B.n787 585
R1147 B.n789 B.n8 585
R1148 B.n791 B.n790 585
R1149 B.n792 B.n7 585
R1150 B.n794 B.n793 585
R1151 B.n795 B.n6 585
R1152 B.n797 B.n796 585
R1153 B.n798 B.n5 585
R1154 B.n800 B.n799 585
R1155 B.n801 B.n4 585
R1156 B.n803 B.n802 585
R1157 B.n804 B.n3 585
R1158 B.n806 B.n805 585
R1159 B.n807 B.n0 585
R1160 B.n2 B.n1 585
R1161 B.n208 B.n207 585
R1162 B.n209 B.n206 585
R1163 B.n211 B.n210 585
R1164 B.n212 B.n205 585
R1165 B.n214 B.n213 585
R1166 B.n215 B.n204 585
R1167 B.n217 B.n216 585
R1168 B.n218 B.n203 585
R1169 B.n220 B.n219 585
R1170 B.n221 B.n202 585
R1171 B.n223 B.n222 585
R1172 B.n224 B.n201 585
R1173 B.n226 B.n225 585
R1174 B.n227 B.n200 585
R1175 B.n229 B.n228 585
R1176 B.n230 B.n199 585
R1177 B.n232 B.n231 585
R1178 B.n233 B.n198 585
R1179 B.n235 B.n234 585
R1180 B.n236 B.n197 585
R1181 B.n238 B.n237 585
R1182 B.n239 B.n196 585
R1183 B.n241 B.n240 585
R1184 B.n242 B.n195 585
R1185 B.n244 B.n243 585
R1186 B.n245 B.n194 585
R1187 B.n247 B.n246 585
R1188 B.n248 B.n193 585
R1189 B.n250 B.n249 585
R1190 B.n251 B.n192 585
R1191 B.n253 B.n252 585
R1192 B.n254 B.n191 585
R1193 B.n256 B.n255 585
R1194 B.n257 B.n190 585
R1195 B.n259 B.n258 585
R1196 B.n260 B.n189 585
R1197 B.n262 B.n261 585
R1198 B.n263 B.n188 585
R1199 B.n265 B.n264 585
R1200 B.n266 B.n187 585
R1201 B.n268 B.n267 585
R1202 B.n269 B.n186 585
R1203 B.n271 B.n270 585
R1204 B.n272 B.n185 585
R1205 B.n274 B.n273 585
R1206 B.n275 B.n184 585
R1207 B.n277 B.n276 585
R1208 B.n278 B.n183 585
R1209 B.n280 B.n279 585
R1210 B.n281 B.n182 585
R1211 B.n283 B.n282 585
R1212 B.n284 B.n181 585
R1213 B.n286 B.n285 585
R1214 B.n287 B.n180 585
R1215 B.n289 B.n288 585
R1216 B.n290 B.n179 585
R1217 B.n292 B.n291 585
R1218 B.n293 B.n178 585
R1219 B.n295 B.n294 585
R1220 B.n296 B.n177 585
R1221 B.n298 B.n297 585
R1222 B.n299 B.n176 585
R1223 B.n301 B.n300 585
R1224 B.n300 B.n175 506.916
R1225 B.n411 B.n410 506.916
R1226 B.n604 B.n73 506.916
R1227 B.n712 B.n711 506.916
R1228 B.n154 B.t1 379.521
R1229 B.n56 B.t11 379.521
R1230 B.n345 B.t4 379.521
R1231 B.n50 B.t8 379.521
R1232 B.n155 B.t2 304.853
R1233 B.n57 B.t10 304.853
R1234 B.n346 B.t5 304.853
R1235 B.n51 B.t7 304.853
R1236 B.n345 B.t3 264.296
R1237 B.n154 B.t0 264.296
R1238 B.n56 B.t9 264.296
R1239 B.n50 B.t6 264.296
R1240 B.n809 B.n808 256.663
R1241 B.n808 B.n807 235.042
R1242 B.n808 B.n2 235.042
R1243 B.n304 B.n175 163.367
R1244 B.n305 B.n304 163.367
R1245 B.n306 B.n305 163.367
R1246 B.n306 B.n173 163.367
R1247 B.n310 B.n173 163.367
R1248 B.n311 B.n310 163.367
R1249 B.n312 B.n311 163.367
R1250 B.n312 B.n171 163.367
R1251 B.n316 B.n171 163.367
R1252 B.n317 B.n316 163.367
R1253 B.n318 B.n317 163.367
R1254 B.n318 B.n169 163.367
R1255 B.n322 B.n169 163.367
R1256 B.n323 B.n322 163.367
R1257 B.n324 B.n323 163.367
R1258 B.n324 B.n167 163.367
R1259 B.n328 B.n167 163.367
R1260 B.n329 B.n328 163.367
R1261 B.n330 B.n329 163.367
R1262 B.n330 B.n165 163.367
R1263 B.n334 B.n165 163.367
R1264 B.n335 B.n334 163.367
R1265 B.n336 B.n335 163.367
R1266 B.n336 B.n163 163.367
R1267 B.n340 B.n163 163.367
R1268 B.n341 B.n340 163.367
R1269 B.n342 B.n341 163.367
R1270 B.n342 B.n161 163.367
R1271 B.n349 B.n161 163.367
R1272 B.n350 B.n349 163.367
R1273 B.n351 B.n350 163.367
R1274 B.n351 B.n159 163.367
R1275 B.n355 B.n159 163.367
R1276 B.n356 B.n355 163.367
R1277 B.n357 B.n356 163.367
R1278 B.n357 B.n157 163.367
R1279 B.n361 B.n157 163.367
R1280 B.n362 B.n361 163.367
R1281 B.n363 B.n362 163.367
R1282 B.n363 B.n153 163.367
R1283 B.n368 B.n153 163.367
R1284 B.n369 B.n368 163.367
R1285 B.n370 B.n369 163.367
R1286 B.n370 B.n151 163.367
R1287 B.n374 B.n151 163.367
R1288 B.n375 B.n374 163.367
R1289 B.n376 B.n375 163.367
R1290 B.n376 B.n149 163.367
R1291 B.n380 B.n149 163.367
R1292 B.n381 B.n380 163.367
R1293 B.n382 B.n381 163.367
R1294 B.n382 B.n147 163.367
R1295 B.n386 B.n147 163.367
R1296 B.n387 B.n386 163.367
R1297 B.n388 B.n387 163.367
R1298 B.n388 B.n145 163.367
R1299 B.n392 B.n145 163.367
R1300 B.n393 B.n392 163.367
R1301 B.n394 B.n393 163.367
R1302 B.n394 B.n143 163.367
R1303 B.n398 B.n143 163.367
R1304 B.n399 B.n398 163.367
R1305 B.n400 B.n399 163.367
R1306 B.n400 B.n141 163.367
R1307 B.n404 B.n141 163.367
R1308 B.n405 B.n404 163.367
R1309 B.n406 B.n405 163.367
R1310 B.n406 B.n139 163.367
R1311 B.n410 B.n139 163.367
R1312 B.n604 B.n603 163.367
R1313 B.n603 B.n602 163.367
R1314 B.n602 B.n75 163.367
R1315 B.n598 B.n75 163.367
R1316 B.n598 B.n597 163.367
R1317 B.n597 B.n596 163.367
R1318 B.n596 B.n77 163.367
R1319 B.n592 B.n77 163.367
R1320 B.n592 B.n591 163.367
R1321 B.n591 B.n590 163.367
R1322 B.n590 B.n79 163.367
R1323 B.n586 B.n79 163.367
R1324 B.n586 B.n585 163.367
R1325 B.n585 B.n584 163.367
R1326 B.n584 B.n81 163.367
R1327 B.n580 B.n81 163.367
R1328 B.n580 B.n579 163.367
R1329 B.n579 B.n578 163.367
R1330 B.n578 B.n83 163.367
R1331 B.n574 B.n83 163.367
R1332 B.n574 B.n573 163.367
R1333 B.n573 B.n572 163.367
R1334 B.n572 B.n85 163.367
R1335 B.n568 B.n85 163.367
R1336 B.n568 B.n567 163.367
R1337 B.n567 B.n566 163.367
R1338 B.n566 B.n87 163.367
R1339 B.n562 B.n87 163.367
R1340 B.n562 B.n561 163.367
R1341 B.n561 B.n560 163.367
R1342 B.n560 B.n89 163.367
R1343 B.n556 B.n89 163.367
R1344 B.n556 B.n555 163.367
R1345 B.n555 B.n554 163.367
R1346 B.n554 B.n91 163.367
R1347 B.n550 B.n91 163.367
R1348 B.n550 B.n549 163.367
R1349 B.n549 B.n548 163.367
R1350 B.n548 B.n93 163.367
R1351 B.n544 B.n93 163.367
R1352 B.n544 B.n543 163.367
R1353 B.n543 B.n542 163.367
R1354 B.n542 B.n95 163.367
R1355 B.n538 B.n95 163.367
R1356 B.n538 B.n537 163.367
R1357 B.n537 B.n536 163.367
R1358 B.n536 B.n97 163.367
R1359 B.n532 B.n97 163.367
R1360 B.n532 B.n531 163.367
R1361 B.n531 B.n530 163.367
R1362 B.n530 B.n99 163.367
R1363 B.n526 B.n99 163.367
R1364 B.n526 B.n525 163.367
R1365 B.n525 B.n524 163.367
R1366 B.n524 B.n101 163.367
R1367 B.n520 B.n101 163.367
R1368 B.n520 B.n519 163.367
R1369 B.n519 B.n518 163.367
R1370 B.n518 B.n103 163.367
R1371 B.n514 B.n103 163.367
R1372 B.n514 B.n513 163.367
R1373 B.n513 B.n512 163.367
R1374 B.n512 B.n105 163.367
R1375 B.n508 B.n105 163.367
R1376 B.n508 B.n507 163.367
R1377 B.n507 B.n506 163.367
R1378 B.n506 B.n107 163.367
R1379 B.n502 B.n107 163.367
R1380 B.n502 B.n501 163.367
R1381 B.n501 B.n500 163.367
R1382 B.n500 B.n109 163.367
R1383 B.n496 B.n109 163.367
R1384 B.n496 B.n495 163.367
R1385 B.n495 B.n494 163.367
R1386 B.n494 B.n111 163.367
R1387 B.n490 B.n111 163.367
R1388 B.n490 B.n489 163.367
R1389 B.n489 B.n488 163.367
R1390 B.n488 B.n113 163.367
R1391 B.n484 B.n113 163.367
R1392 B.n484 B.n483 163.367
R1393 B.n483 B.n482 163.367
R1394 B.n482 B.n115 163.367
R1395 B.n478 B.n115 163.367
R1396 B.n478 B.n477 163.367
R1397 B.n477 B.n476 163.367
R1398 B.n476 B.n117 163.367
R1399 B.n472 B.n117 163.367
R1400 B.n472 B.n471 163.367
R1401 B.n471 B.n470 163.367
R1402 B.n470 B.n119 163.367
R1403 B.n466 B.n119 163.367
R1404 B.n466 B.n465 163.367
R1405 B.n465 B.n464 163.367
R1406 B.n464 B.n121 163.367
R1407 B.n460 B.n121 163.367
R1408 B.n460 B.n459 163.367
R1409 B.n459 B.n458 163.367
R1410 B.n458 B.n123 163.367
R1411 B.n454 B.n123 163.367
R1412 B.n454 B.n453 163.367
R1413 B.n453 B.n452 163.367
R1414 B.n452 B.n125 163.367
R1415 B.n448 B.n125 163.367
R1416 B.n448 B.n447 163.367
R1417 B.n447 B.n446 163.367
R1418 B.n446 B.n127 163.367
R1419 B.n442 B.n127 163.367
R1420 B.n442 B.n441 163.367
R1421 B.n441 B.n440 163.367
R1422 B.n440 B.n129 163.367
R1423 B.n436 B.n129 163.367
R1424 B.n436 B.n435 163.367
R1425 B.n435 B.n434 163.367
R1426 B.n434 B.n131 163.367
R1427 B.n430 B.n131 163.367
R1428 B.n430 B.n429 163.367
R1429 B.n429 B.n428 163.367
R1430 B.n428 B.n133 163.367
R1431 B.n424 B.n133 163.367
R1432 B.n424 B.n423 163.367
R1433 B.n423 B.n422 163.367
R1434 B.n422 B.n135 163.367
R1435 B.n418 B.n135 163.367
R1436 B.n418 B.n417 163.367
R1437 B.n417 B.n416 163.367
R1438 B.n416 B.n137 163.367
R1439 B.n412 B.n137 163.367
R1440 B.n412 B.n411 163.367
R1441 B.n711 B.n710 163.367
R1442 B.n710 B.n35 163.367
R1443 B.n706 B.n35 163.367
R1444 B.n706 B.n705 163.367
R1445 B.n705 B.n704 163.367
R1446 B.n704 B.n37 163.367
R1447 B.n700 B.n37 163.367
R1448 B.n700 B.n699 163.367
R1449 B.n699 B.n698 163.367
R1450 B.n698 B.n39 163.367
R1451 B.n694 B.n39 163.367
R1452 B.n694 B.n693 163.367
R1453 B.n693 B.n692 163.367
R1454 B.n692 B.n41 163.367
R1455 B.n688 B.n41 163.367
R1456 B.n688 B.n687 163.367
R1457 B.n687 B.n686 163.367
R1458 B.n686 B.n43 163.367
R1459 B.n682 B.n43 163.367
R1460 B.n682 B.n681 163.367
R1461 B.n681 B.n680 163.367
R1462 B.n680 B.n45 163.367
R1463 B.n676 B.n45 163.367
R1464 B.n676 B.n675 163.367
R1465 B.n675 B.n674 163.367
R1466 B.n674 B.n47 163.367
R1467 B.n670 B.n47 163.367
R1468 B.n670 B.n669 163.367
R1469 B.n669 B.n668 163.367
R1470 B.n668 B.n49 163.367
R1471 B.n663 B.n49 163.367
R1472 B.n663 B.n662 163.367
R1473 B.n662 B.n661 163.367
R1474 B.n661 B.n53 163.367
R1475 B.n657 B.n53 163.367
R1476 B.n657 B.n656 163.367
R1477 B.n656 B.n655 163.367
R1478 B.n655 B.n55 163.367
R1479 B.n651 B.n55 163.367
R1480 B.n651 B.n650 163.367
R1481 B.n650 B.n59 163.367
R1482 B.n646 B.n59 163.367
R1483 B.n646 B.n645 163.367
R1484 B.n645 B.n644 163.367
R1485 B.n644 B.n61 163.367
R1486 B.n640 B.n61 163.367
R1487 B.n640 B.n639 163.367
R1488 B.n639 B.n638 163.367
R1489 B.n638 B.n63 163.367
R1490 B.n634 B.n63 163.367
R1491 B.n634 B.n633 163.367
R1492 B.n633 B.n632 163.367
R1493 B.n632 B.n65 163.367
R1494 B.n628 B.n65 163.367
R1495 B.n628 B.n627 163.367
R1496 B.n627 B.n626 163.367
R1497 B.n626 B.n67 163.367
R1498 B.n622 B.n67 163.367
R1499 B.n622 B.n621 163.367
R1500 B.n621 B.n620 163.367
R1501 B.n620 B.n69 163.367
R1502 B.n616 B.n69 163.367
R1503 B.n616 B.n615 163.367
R1504 B.n615 B.n614 163.367
R1505 B.n614 B.n71 163.367
R1506 B.n610 B.n71 163.367
R1507 B.n610 B.n609 163.367
R1508 B.n609 B.n608 163.367
R1509 B.n608 B.n73 163.367
R1510 B.n712 B.n33 163.367
R1511 B.n716 B.n33 163.367
R1512 B.n717 B.n716 163.367
R1513 B.n718 B.n717 163.367
R1514 B.n718 B.n31 163.367
R1515 B.n722 B.n31 163.367
R1516 B.n723 B.n722 163.367
R1517 B.n724 B.n723 163.367
R1518 B.n724 B.n29 163.367
R1519 B.n728 B.n29 163.367
R1520 B.n729 B.n728 163.367
R1521 B.n730 B.n729 163.367
R1522 B.n730 B.n27 163.367
R1523 B.n734 B.n27 163.367
R1524 B.n735 B.n734 163.367
R1525 B.n736 B.n735 163.367
R1526 B.n736 B.n25 163.367
R1527 B.n740 B.n25 163.367
R1528 B.n741 B.n740 163.367
R1529 B.n742 B.n741 163.367
R1530 B.n742 B.n23 163.367
R1531 B.n746 B.n23 163.367
R1532 B.n747 B.n746 163.367
R1533 B.n748 B.n747 163.367
R1534 B.n748 B.n21 163.367
R1535 B.n752 B.n21 163.367
R1536 B.n753 B.n752 163.367
R1537 B.n754 B.n753 163.367
R1538 B.n754 B.n19 163.367
R1539 B.n758 B.n19 163.367
R1540 B.n759 B.n758 163.367
R1541 B.n760 B.n759 163.367
R1542 B.n760 B.n17 163.367
R1543 B.n764 B.n17 163.367
R1544 B.n765 B.n764 163.367
R1545 B.n766 B.n765 163.367
R1546 B.n766 B.n15 163.367
R1547 B.n770 B.n15 163.367
R1548 B.n771 B.n770 163.367
R1549 B.n772 B.n771 163.367
R1550 B.n772 B.n13 163.367
R1551 B.n776 B.n13 163.367
R1552 B.n777 B.n776 163.367
R1553 B.n778 B.n777 163.367
R1554 B.n778 B.n11 163.367
R1555 B.n782 B.n11 163.367
R1556 B.n783 B.n782 163.367
R1557 B.n784 B.n783 163.367
R1558 B.n784 B.n9 163.367
R1559 B.n788 B.n9 163.367
R1560 B.n789 B.n788 163.367
R1561 B.n790 B.n789 163.367
R1562 B.n790 B.n7 163.367
R1563 B.n794 B.n7 163.367
R1564 B.n795 B.n794 163.367
R1565 B.n796 B.n795 163.367
R1566 B.n796 B.n5 163.367
R1567 B.n800 B.n5 163.367
R1568 B.n801 B.n800 163.367
R1569 B.n802 B.n801 163.367
R1570 B.n802 B.n3 163.367
R1571 B.n806 B.n3 163.367
R1572 B.n807 B.n806 163.367
R1573 B.n208 B.n2 163.367
R1574 B.n209 B.n208 163.367
R1575 B.n210 B.n209 163.367
R1576 B.n210 B.n205 163.367
R1577 B.n214 B.n205 163.367
R1578 B.n215 B.n214 163.367
R1579 B.n216 B.n215 163.367
R1580 B.n216 B.n203 163.367
R1581 B.n220 B.n203 163.367
R1582 B.n221 B.n220 163.367
R1583 B.n222 B.n221 163.367
R1584 B.n222 B.n201 163.367
R1585 B.n226 B.n201 163.367
R1586 B.n227 B.n226 163.367
R1587 B.n228 B.n227 163.367
R1588 B.n228 B.n199 163.367
R1589 B.n232 B.n199 163.367
R1590 B.n233 B.n232 163.367
R1591 B.n234 B.n233 163.367
R1592 B.n234 B.n197 163.367
R1593 B.n238 B.n197 163.367
R1594 B.n239 B.n238 163.367
R1595 B.n240 B.n239 163.367
R1596 B.n240 B.n195 163.367
R1597 B.n244 B.n195 163.367
R1598 B.n245 B.n244 163.367
R1599 B.n246 B.n245 163.367
R1600 B.n246 B.n193 163.367
R1601 B.n250 B.n193 163.367
R1602 B.n251 B.n250 163.367
R1603 B.n252 B.n251 163.367
R1604 B.n252 B.n191 163.367
R1605 B.n256 B.n191 163.367
R1606 B.n257 B.n256 163.367
R1607 B.n258 B.n257 163.367
R1608 B.n258 B.n189 163.367
R1609 B.n262 B.n189 163.367
R1610 B.n263 B.n262 163.367
R1611 B.n264 B.n263 163.367
R1612 B.n264 B.n187 163.367
R1613 B.n268 B.n187 163.367
R1614 B.n269 B.n268 163.367
R1615 B.n270 B.n269 163.367
R1616 B.n270 B.n185 163.367
R1617 B.n274 B.n185 163.367
R1618 B.n275 B.n274 163.367
R1619 B.n276 B.n275 163.367
R1620 B.n276 B.n183 163.367
R1621 B.n280 B.n183 163.367
R1622 B.n281 B.n280 163.367
R1623 B.n282 B.n281 163.367
R1624 B.n282 B.n181 163.367
R1625 B.n286 B.n181 163.367
R1626 B.n287 B.n286 163.367
R1627 B.n288 B.n287 163.367
R1628 B.n288 B.n179 163.367
R1629 B.n292 B.n179 163.367
R1630 B.n293 B.n292 163.367
R1631 B.n294 B.n293 163.367
R1632 B.n294 B.n177 163.367
R1633 B.n298 B.n177 163.367
R1634 B.n299 B.n298 163.367
R1635 B.n300 B.n299 163.367
R1636 B.n346 B.n345 74.6672
R1637 B.n155 B.n154 74.6672
R1638 B.n57 B.n56 74.6672
R1639 B.n51 B.n50 74.6672
R1640 B.n347 B.n346 59.5399
R1641 B.n365 B.n155 59.5399
R1642 B.n58 B.n57 59.5399
R1643 B.n666 B.n51 59.5399
R1644 B.n713 B.n34 32.9371
R1645 B.n606 B.n605 32.9371
R1646 B.n409 B.n138 32.9371
R1647 B.n302 B.n301 32.9371
R1648 B B.n809 18.0485
R1649 B.n714 B.n713 10.6151
R1650 B.n715 B.n714 10.6151
R1651 B.n715 B.n32 10.6151
R1652 B.n719 B.n32 10.6151
R1653 B.n720 B.n719 10.6151
R1654 B.n721 B.n720 10.6151
R1655 B.n721 B.n30 10.6151
R1656 B.n725 B.n30 10.6151
R1657 B.n726 B.n725 10.6151
R1658 B.n727 B.n726 10.6151
R1659 B.n727 B.n28 10.6151
R1660 B.n731 B.n28 10.6151
R1661 B.n732 B.n731 10.6151
R1662 B.n733 B.n732 10.6151
R1663 B.n733 B.n26 10.6151
R1664 B.n737 B.n26 10.6151
R1665 B.n738 B.n737 10.6151
R1666 B.n739 B.n738 10.6151
R1667 B.n739 B.n24 10.6151
R1668 B.n743 B.n24 10.6151
R1669 B.n744 B.n743 10.6151
R1670 B.n745 B.n744 10.6151
R1671 B.n745 B.n22 10.6151
R1672 B.n749 B.n22 10.6151
R1673 B.n750 B.n749 10.6151
R1674 B.n751 B.n750 10.6151
R1675 B.n751 B.n20 10.6151
R1676 B.n755 B.n20 10.6151
R1677 B.n756 B.n755 10.6151
R1678 B.n757 B.n756 10.6151
R1679 B.n757 B.n18 10.6151
R1680 B.n761 B.n18 10.6151
R1681 B.n762 B.n761 10.6151
R1682 B.n763 B.n762 10.6151
R1683 B.n763 B.n16 10.6151
R1684 B.n767 B.n16 10.6151
R1685 B.n768 B.n767 10.6151
R1686 B.n769 B.n768 10.6151
R1687 B.n769 B.n14 10.6151
R1688 B.n773 B.n14 10.6151
R1689 B.n774 B.n773 10.6151
R1690 B.n775 B.n774 10.6151
R1691 B.n775 B.n12 10.6151
R1692 B.n779 B.n12 10.6151
R1693 B.n780 B.n779 10.6151
R1694 B.n781 B.n780 10.6151
R1695 B.n781 B.n10 10.6151
R1696 B.n785 B.n10 10.6151
R1697 B.n786 B.n785 10.6151
R1698 B.n787 B.n786 10.6151
R1699 B.n787 B.n8 10.6151
R1700 B.n791 B.n8 10.6151
R1701 B.n792 B.n791 10.6151
R1702 B.n793 B.n792 10.6151
R1703 B.n793 B.n6 10.6151
R1704 B.n797 B.n6 10.6151
R1705 B.n798 B.n797 10.6151
R1706 B.n799 B.n798 10.6151
R1707 B.n799 B.n4 10.6151
R1708 B.n803 B.n4 10.6151
R1709 B.n804 B.n803 10.6151
R1710 B.n805 B.n804 10.6151
R1711 B.n805 B.n0 10.6151
R1712 B.n709 B.n34 10.6151
R1713 B.n709 B.n708 10.6151
R1714 B.n708 B.n707 10.6151
R1715 B.n707 B.n36 10.6151
R1716 B.n703 B.n36 10.6151
R1717 B.n703 B.n702 10.6151
R1718 B.n702 B.n701 10.6151
R1719 B.n701 B.n38 10.6151
R1720 B.n697 B.n38 10.6151
R1721 B.n697 B.n696 10.6151
R1722 B.n696 B.n695 10.6151
R1723 B.n695 B.n40 10.6151
R1724 B.n691 B.n40 10.6151
R1725 B.n691 B.n690 10.6151
R1726 B.n690 B.n689 10.6151
R1727 B.n689 B.n42 10.6151
R1728 B.n685 B.n42 10.6151
R1729 B.n685 B.n684 10.6151
R1730 B.n684 B.n683 10.6151
R1731 B.n683 B.n44 10.6151
R1732 B.n679 B.n44 10.6151
R1733 B.n679 B.n678 10.6151
R1734 B.n678 B.n677 10.6151
R1735 B.n677 B.n46 10.6151
R1736 B.n673 B.n46 10.6151
R1737 B.n673 B.n672 10.6151
R1738 B.n672 B.n671 10.6151
R1739 B.n671 B.n48 10.6151
R1740 B.n667 B.n48 10.6151
R1741 B.n665 B.n664 10.6151
R1742 B.n664 B.n52 10.6151
R1743 B.n660 B.n52 10.6151
R1744 B.n660 B.n659 10.6151
R1745 B.n659 B.n658 10.6151
R1746 B.n658 B.n54 10.6151
R1747 B.n654 B.n54 10.6151
R1748 B.n654 B.n653 10.6151
R1749 B.n653 B.n652 10.6151
R1750 B.n649 B.n648 10.6151
R1751 B.n648 B.n647 10.6151
R1752 B.n647 B.n60 10.6151
R1753 B.n643 B.n60 10.6151
R1754 B.n643 B.n642 10.6151
R1755 B.n642 B.n641 10.6151
R1756 B.n641 B.n62 10.6151
R1757 B.n637 B.n62 10.6151
R1758 B.n637 B.n636 10.6151
R1759 B.n636 B.n635 10.6151
R1760 B.n635 B.n64 10.6151
R1761 B.n631 B.n64 10.6151
R1762 B.n631 B.n630 10.6151
R1763 B.n630 B.n629 10.6151
R1764 B.n629 B.n66 10.6151
R1765 B.n625 B.n66 10.6151
R1766 B.n625 B.n624 10.6151
R1767 B.n624 B.n623 10.6151
R1768 B.n623 B.n68 10.6151
R1769 B.n619 B.n68 10.6151
R1770 B.n619 B.n618 10.6151
R1771 B.n618 B.n617 10.6151
R1772 B.n617 B.n70 10.6151
R1773 B.n613 B.n70 10.6151
R1774 B.n613 B.n612 10.6151
R1775 B.n612 B.n611 10.6151
R1776 B.n611 B.n72 10.6151
R1777 B.n607 B.n72 10.6151
R1778 B.n607 B.n606 10.6151
R1779 B.n605 B.n74 10.6151
R1780 B.n601 B.n74 10.6151
R1781 B.n601 B.n600 10.6151
R1782 B.n600 B.n599 10.6151
R1783 B.n599 B.n76 10.6151
R1784 B.n595 B.n76 10.6151
R1785 B.n595 B.n594 10.6151
R1786 B.n594 B.n593 10.6151
R1787 B.n593 B.n78 10.6151
R1788 B.n589 B.n78 10.6151
R1789 B.n589 B.n588 10.6151
R1790 B.n588 B.n587 10.6151
R1791 B.n587 B.n80 10.6151
R1792 B.n583 B.n80 10.6151
R1793 B.n583 B.n582 10.6151
R1794 B.n582 B.n581 10.6151
R1795 B.n581 B.n82 10.6151
R1796 B.n577 B.n82 10.6151
R1797 B.n577 B.n576 10.6151
R1798 B.n576 B.n575 10.6151
R1799 B.n575 B.n84 10.6151
R1800 B.n571 B.n84 10.6151
R1801 B.n571 B.n570 10.6151
R1802 B.n570 B.n569 10.6151
R1803 B.n569 B.n86 10.6151
R1804 B.n565 B.n86 10.6151
R1805 B.n565 B.n564 10.6151
R1806 B.n564 B.n563 10.6151
R1807 B.n563 B.n88 10.6151
R1808 B.n559 B.n88 10.6151
R1809 B.n559 B.n558 10.6151
R1810 B.n558 B.n557 10.6151
R1811 B.n557 B.n90 10.6151
R1812 B.n553 B.n90 10.6151
R1813 B.n553 B.n552 10.6151
R1814 B.n552 B.n551 10.6151
R1815 B.n551 B.n92 10.6151
R1816 B.n547 B.n92 10.6151
R1817 B.n547 B.n546 10.6151
R1818 B.n546 B.n545 10.6151
R1819 B.n545 B.n94 10.6151
R1820 B.n541 B.n94 10.6151
R1821 B.n541 B.n540 10.6151
R1822 B.n540 B.n539 10.6151
R1823 B.n539 B.n96 10.6151
R1824 B.n535 B.n96 10.6151
R1825 B.n535 B.n534 10.6151
R1826 B.n534 B.n533 10.6151
R1827 B.n533 B.n98 10.6151
R1828 B.n529 B.n98 10.6151
R1829 B.n529 B.n528 10.6151
R1830 B.n528 B.n527 10.6151
R1831 B.n527 B.n100 10.6151
R1832 B.n523 B.n100 10.6151
R1833 B.n523 B.n522 10.6151
R1834 B.n522 B.n521 10.6151
R1835 B.n521 B.n102 10.6151
R1836 B.n517 B.n102 10.6151
R1837 B.n517 B.n516 10.6151
R1838 B.n516 B.n515 10.6151
R1839 B.n515 B.n104 10.6151
R1840 B.n511 B.n104 10.6151
R1841 B.n511 B.n510 10.6151
R1842 B.n510 B.n509 10.6151
R1843 B.n509 B.n106 10.6151
R1844 B.n505 B.n106 10.6151
R1845 B.n505 B.n504 10.6151
R1846 B.n504 B.n503 10.6151
R1847 B.n503 B.n108 10.6151
R1848 B.n499 B.n108 10.6151
R1849 B.n499 B.n498 10.6151
R1850 B.n498 B.n497 10.6151
R1851 B.n497 B.n110 10.6151
R1852 B.n493 B.n110 10.6151
R1853 B.n493 B.n492 10.6151
R1854 B.n492 B.n491 10.6151
R1855 B.n491 B.n112 10.6151
R1856 B.n487 B.n112 10.6151
R1857 B.n487 B.n486 10.6151
R1858 B.n486 B.n485 10.6151
R1859 B.n485 B.n114 10.6151
R1860 B.n481 B.n114 10.6151
R1861 B.n481 B.n480 10.6151
R1862 B.n480 B.n479 10.6151
R1863 B.n479 B.n116 10.6151
R1864 B.n475 B.n116 10.6151
R1865 B.n475 B.n474 10.6151
R1866 B.n474 B.n473 10.6151
R1867 B.n473 B.n118 10.6151
R1868 B.n469 B.n118 10.6151
R1869 B.n469 B.n468 10.6151
R1870 B.n468 B.n467 10.6151
R1871 B.n467 B.n120 10.6151
R1872 B.n463 B.n120 10.6151
R1873 B.n463 B.n462 10.6151
R1874 B.n462 B.n461 10.6151
R1875 B.n461 B.n122 10.6151
R1876 B.n457 B.n122 10.6151
R1877 B.n457 B.n456 10.6151
R1878 B.n456 B.n455 10.6151
R1879 B.n455 B.n124 10.6151
R1880 B.n451 B.n124 10.6151
R1881 B.n451 B.n450 10.6151
R1882 B.n450 B.n449 10.6151
R1883 B.n449 B.n126 10.6151
R1884 B.n445 B.n126 10.6151
R1885 B.n445 B.n444 10.6151
R1886 B.n444 B.n443 10.6151
R1887 B.n443 B.n128 10.6151
R1888 B.n439 B.n128 10.6151
R1889 B.n439 B.n438 10.6151
R1890 B.n438 B.n437 10.6151
R1891 B.n437 B.n130 10.6151
R1892 B.n433 B.n130 10.6151
R1893 B.n433 B.n432 10.6151
R1894 B.n432 B.n431 10.6151
R1895 B.n431 B.n132 10.6151
R1896 B.n427 B.n132 10.6151
R1897 B.n427 B.n426 10.6151
R1898 B.n426 B.n425 10.6151
R1899 B.n425 B.n134 10.6151
R1900 B.n421 B.n134 10.6151
R1901 B.n421 B.n420 10.6151
R1902 B.n420 B.n419 10.6151
R1903 B.n419 B.n136 10.6151
R1904 B.n415 B.n136 10.6151
R1905 B.n415 B.n414 10.6151
R1906 B.n414 B.n413 10.6151
R1907 B.n413 B.n138 10.6151
R1908 B.n207 B.n1 10.6151
R1909 B.n207 B.n206 10.6151
R1910 B.n211 B.n206 10.6151
R1911 B.n212 B.n211 10.6151
R1912 B.n213 B.n212 10.6151
R1913 B.n213 B.n204 10.6151
R1914 B.n217 B.n204 10.6151
R1915 B.n218 B.n217 10.6151
R1916 B.n219 B.n218 10.6151
R1917 B.n219 B.n202 10.6151
R1918 B.n223 B.n202 10.6151
R1919 B.n224 B.n223 10.6151
R1920 B.n225 B.n224 10.6151
R1921 B.n225 B.n200 10.6151
R1922 B.n229 B.n200 10.6151
R1923 B.n230 B.n229 10.6151
R1924 B.n231 B.n230 10.6151
R1925 B.n231 B.n198 10.6151
R1926 B.n235 B.n198 10.6151
R1927 B.n236 B.n235 10.6151
R1928 B.n237 B.n236 10.6151
R1929 B.n237 B.n196 10.6151
R1930 B.n241 B.n196 10.6151
R1931 B.n242 B.n241 10.6151
R1932 B.n243 B.n242 10.6151
R1933 B.n243 B.n194 10.6151
R1934 B.n247 B.n194 10.6151
R1935 B.n248 B.n247 10.6151
R1936 B.n249 B.n248 10.6151
R1937 B.n249 B.n192 10.6151
R1938 B.n253 B.n192 10.6151
R1939 B.n254 B.n253 10.6151
R1940 B.n255 B.n254 10.6151
R1941 B.n255 B.n190 10.6151
R1942 B.n259 B.n190 10.6151
R1943 B.n260 B.n259 10.6151
R1944 B.n261 B.n260 10.6151
R1945 B.n261 B.n188 10.6151
R1946 B.n265 B.n188 10.6151
R1947 B.n266 B.n265 10.6151
R1948 B.n267 B.n266 10.6151
R1949 B.n267 B.n186 10.6151
R1950 B.n271 B.n186 10.6151
R1951 B.n272 B.n271 10.6151
R1952 B.n273 B.n272 10.6151
R1953 B.n273 B.n184 10.6151
R1954 B.n277 B.n184 10.6151
R1955 B.n278 B.n277 10.6151
R1956 B.n279 B.n278 10.6151
R1957 B.n279 B.n182 10.6151
R1958 B.n283 B.n182 10.6151
R1959 B.n284 B.n283 10.6151
R1960 B.n285 B.n284 10.6151
R1961 B.n285 B.n180 10.6151
R1962 B.n289 B.n180 10.6151
R1963 B.n290 B.n289 10.6151
R1964 B.n291 B.n290 10.6151
R1965 B.n291 B.n178 10.6151
R1966 B.n295 B.n178 10.6151
R1967 B.n296 B.n295 10.6151
R1968 B.n297 B.n296 10.6151
R1969 B.n297 B.n176 10.6151
R1970 B.n301 B.n176 10.6151
R1971 B.n303 B.n302 10.6151
R1972 B.n303 B.n174 10.6151
R1973 B.n307 B.n174 10.6151
R1974 B.n308 B.n307 10.6151
R1975 B.n309 B.n308 10.6151
R1976 B.n309 B.n172 10.6151
R1977 B.n313 B.n172 10.6151
R1978 B.n314 B.n313 10.6151
R1979 B.n315 B.n314 10.6151
R1980 B.n315 B.n170 10.6151
R1981 B.n319 B.n170 10.6151
R1982 B.n320 B.n319 10.6151
R1983 B.n321 B.n320 10.6151
R1984 B.n321 B.n168 10.6151
R1985 B.n325 B.n168 10.6151
R1986 B.n326 B.n325 10.6151
R1987 B.n327 B.n326 10.6151
R1988 B.n327 B.n166 10.6151
R1989 B.n331 B.n166 10.6151
R1990 B.n332 B.n331 10.6151
R1991 B.n333 B.n332 10.6151
R1992 B.n333 B.n164 10.6151
R1993 B.n337 B.n164 10.6151
R1994 B.n338 B.n337 10.6151
R1995 B.n339 B.n338 10.6151
R1996 B.n339 B.n162 10.6151
R1997 B.n343 B.n162 10.6151
R1998 B.n344 B.n343 10.6151
R1999 B.n348 B.n344 10.6151
R2000 B.n352 B.n160 10.6151
R2001 B.n353 B.n352 10.6151
R2002 B.n354 B.n353 10.6151
R2003 B.n354 B.n158 10.6151
R2004 B.n358 B.n158 10.6151
R2005 B.n359 B.n358 10.6151
R2006 B.n360 B.n359 10.6151
R2007 B.n360 B.n156 10.6151
R2008 B.n364 B.n156 10.6151
R2009 B.n367 B.n366 10.6151
R2010 B.n367 B.n152 10.6151
R2011 B.n371 B.n152 10.6151
R2012 B.n372 B.n371 10.6151
R2013 B.n373 B.n372 10.6151
R2014 B.n373 B.n150 10.6151
R2015 B.n377 B.n150 10.6151
R2016 B.n378 B.n377 10.6151
R2017 B.n379 B.n378 10.6151
R2018 B.n379 B.n148 10.6151
R2019 B.n383 B.n148 10.6151
R2020 B.n384 B.n383 10.6151
R2021 B.n385 B.n384 10.6151
R2022 B.n385 B.n146 10.6151
R2023 B.n389 B.n146 10.6151
R2024 B.n390 B.n389 10.6151
R2025 B.n391 B.n390 10.6151
R2026 B.n391 B.n144 10.6151
R2027 B.n395 B.n144 10.6151
R2028 B.n396 B.n395 10.6151
R2029 B.n397 B.n396 10.6151
R2030 B.n397 B.n142 10.6151
R2031 B.n401 B.n142 10.6151
R2032 B.n402 B.n401 10.6151
R2033 B.n403 B.n402 10.6151
R2034 B.n403 B.n140 10.6151
R2035 B.n407 B.n140 10.6151
R2036 B.n408 B.n407 10.6151
R2037 B.n409 B.n408 10.6151
R2038 B.n667 B.n666 9.36635
R2039 B.n649 B.n58 9.36635
R2040 B.n348 B.n347 9.36635
R2041 B.n366 B.n365 9.36635
R2042 B.n809 B.n0 8.11757
R2043 B.n809 B.n1 8.11757
R2044 B.n666 B.n665 1.24928
R2045 B.n652 B.n58 1.24928
R2046 B.n347 B.n160 1.24928
R2047 B.n365 B.n364 1.24928
C0 VTAIL VDD2 7.367759f
C1 VDD1 B 1.82404f
C2 VP B 2.44694f
C3 VTAIL w_n4820_n2580# 3.4254f
C4 VDD1 VP 6.76221f
C5 VTAIL VN 7.19667f
C6 w_n4820_n2580# VDD2 2.29987f
C7 VDD2 VN 6.29989f
C8 w_n4820_n2580# VN 9.99991f
C9 VTAIL B 4.0158f
C10 VTAIL VDD1 7.30718f
C11 VTAIL VP 7.21078f
C12 VDD2 B 1.94901f
C13 VDD1 VDD2 2.25466f
C14 VP VDD2 0.617303f
C15 w_n4820_n2580# B 10.419f
C16 VDD1 w_n4820_n2580# 2.14657f
C17 VP w_n4820_n2580# 10.6284f
C18 B VN 1.38854f
C19 VDD1 VN 0.153126f
C20 VP VN 8.0638f
C21 VDD2 VSUBS 2.261012f
C22 VDD1 VSUBS 3.07082f
C23 VTAIL VSUBS 1.346313f
C24 VN VSUBS 7.940609f
C25 VP VSUBS 4.397891f
C26 B VSUBS 5.696528f
C27 w_n4820_n2580# VSUBS 0.154259p
C28 B.n0 VSUBS 0.007299f
C29 B.n1 VSUBS 0.007299f
C30 B.n2 VSUBS 0.010794f
C31 B.n3 VSUBS 0.008272f
C32 B.n4 VSUBS 0.008272f
C33 B.n5 VSUBS 0.008272f
C34 B.n6 VSUBS 0.008272f
C35 B.n7 VSUBS 0.008272f
C36 B.n8 VSUBS 0.008272f
C37 B.n9 VSUBS 0.008272f
C38 B.n10 VSUBS 0.008272f
C39 B.n11 VSUBS 0.008272f
C40 B.n12 VSUBS 0.008272f
C41 B.n13 VSUBS 0.008272f
C42 B.n14 VSUBS 0.008272f
C43 B.n15 VSUBS 0.008272f
C44 B.n16 VSUBS 0.008272f
C45 B.n17 VSUBS 0.008272f
C46 B.n18 VSUBS 0.008272f
C47 B.n19 VSUBS 0.008272f
C48 B.n20 VSUBS 0.008272f
C49 B.n21 VSUBS 0.008272f
C50 B.n22 VSUBS 0.008272f
C51 B.n23 VSUBS 0.008272f
C52 B.n24 VSUBS 0.008272f
C53 B.n25 VSUBS 0.008272f
C54 B.n26 VSUBS 0.008272f
C55 B.n27 VSUBS 0.008272f
C56 B.n28 VSUBS 0.008272f
C57 B.n29 VSUBS 0.008272f
C58 B.n30 VSUBS 0.008272f
C59 B.n31 VSUBS 0.008272f
C60 B.n32 VSUBS 0.008272f
C61 B.n33 VSUBS 0.008272f
C62 B.n34 VSUBS 0.020255f
C63 B.n35 VSUBS 0.008272f
C64 B.n36 VSUBS 0.008272f
C65 B.n37 VSUBS 0.008272f
C66 B.n38 VSUBS 0.008272f
C67 B.n39 VSUBS 0.008272f
C68 B.n40 VSUBS 0.008272f
C69 B.n41 VSUBS 0.008272f
C70 B.n42 VSUBS 0.008272f
C71 B.n43 VSUBS 0.008272f
C72 B.n44 VSUBS 0.008272f
C73 B.n45 VSUBS 0.008272f
C74 B.n46 VSUBS 0.008272f
C75 B.n47 VSUBS 0.008272f
C76 B.n48 VSUBS 0.008272f
C77 B.n49 VSUBS 0.008272f
C78 B.t7 VSUBS 0.151176f
C79 B.t8 VSUBS 0.194489f
C80 B.t6 VSUBS 1.58765f
C81 B.n50 VSUBS 0.316864f
C82 B.n51 VSUBS 0.231951f
C83 B.n52 VSUBS 0.008272f
C84 B.n53 VSUBS 0.008272f
C85 B.n54 VSUBS 0.008272f
C86 B.n55 VSUBS 0.008272f
C87 B.t10 VSUBS 0.151179f
C88 B.t11 VSUBS 0.194491f
C89 B.t9 VSUBS 1.58765f
C90 B.n56 VSUBS 0.316862f
C91 B.n57 VSUBS 0.231949f
C92 B.n58 VSUBS 0.019165f
C93 B.n59 VSUBS 0.008272f
C94 B.n60 VSUBS 0.008272f
C95 B.n61 VSUBS 0.008272f
C96 B.n62 VSUBS 0.008272f
C97 B.n63 VSUBS 0.008272f
C98 B.n64 VSUBS 0.008272f
C99 B.n65 VSUBS 0.008272f
C100 B.n66 VSUBS 0.008272f
C101 B.n67 VSUBS 0.008272f
C102 B.n68 VSUBS 0.008272f
C103 B.n69 VSUBS 0.008272f
C104 B.n70 VSUBS 0.008272f
C105 B.n71 VSUBS 0.008272f
C106 B.n72 VSUBS 0.008272f
C107 B.n73 VSUBS 0.020255f
C108 B.n74 VSUBS 0.008272f
C109 B.n75 VSUBS 0.008272f
C110 B.n76 VSUBS 0.008272f
C111 B.n77 VSUBS 0.008272f
C112 B.n78 VSUBS 0.008272f
C113 B.n79 VSUBS 0.008272f
C114 B.n80 VSUBS 0.008272f
C115 B.n81 VSUBS 0.008272f
C116 B.n82 VSUBS 0.008272f
C117 B.n83 VSUBS 0.008272f
C118 B.n84 VSUBS 0.008272f
C119 B.n85 VSUBS 0.008272f
C120 B.n86 VSUBS 0.008272f
C121 B.n87 VSUBS 0.008272f
C122 B.n88 VSUBS 0.008272f
C123 B.n89 VSUBS 0.008272f
C124 B.n90 VSUBS 0.008272f
C125 B.n91 VSUBS 0.008272f
C126 B.n92 VSUBS 0.008272f
C127 B.n93 VSUBS 0.008272f
C128 B.n94 VSUBS 0.008272f
C129 B.n95 VSUBS 0.008272f
C130 B.n96 VSUBS 0.008272f
C131 B.n97 VSUBS 0.008272f
C132 B.n98 VSUBS 0.008272f
C133 B.n99 VSUBS 0.008272f
C134 B.n100 VSUBS 0.008272f
C135 B.n101 VSUBS 0.008272f
C136 B.n102 VSUBS 0.008272f
C137 B.n103 VSUBS 0.008272f
C138 B.n104 VSUBS 0.008272f
C139 B.n105 VSUBS 0.008272f
C140 B.n106 VSUBS 0.008272f
C141 B.n107 VSUBS 0.008272f
C142 B.n108 VSUBS 0.008272f
C143 B.n109 VSUBS 0.008272f
C144 B.n110 VSUBS 0.008272f
C145 B.n111 VSUBS 0.008272f
C146 B.n112 VSUBS 0.008272f
C147 B.n113 VSUBS 0.008272f
C148 B.n114 VSUBS 0.008272f
C149 B.n115 VSUBS 0.008272f
C150 B.n116 VSUBS 0.008272f
C151 B.n117 VSUBS 0.008272f
C152 B.n118 VSUBS 0.008272f
C153 B.n119 VSUBS 0.008272f
C154 B.n120 VSUBS 0.008272f
C155 B.n121 VSUBS 0.008272f
C156 B.n122 VSUBS 0.008272f
C157 B.n123 VSUBS 0.008272f
C158 B.n124 VSUBS 0.008272f
C159 B.n125 VSUBS 0.008272f
C160 B.n126 VSUBS 0.008272f
C161 B.n127 VSUBS 0.008272f
C162 B.n128 VSUBS 0.008272f
C163 B.n129 VSUBS 0.008272f
C164 B.n130 VSUBS 0.008272f
C165 B.n131 VSUBS 0.008272f
C166 B.n132 VSUBS 0.008272f
C167 B.n133 VSUBS 0.008272f
C168 B.n134 VSUBS 0.008272f
C169 B.n135 VSUBS 0.008272f
C170 B.n136 VSUBS 0.008272f
C171 B.n137 VSUBS 0.008272f
C172 B.n138 VSUBS 0.01964f
C173 B.n139 VSUBS 0.008272f
C174 B.n140 VSUBS 0.008272f
C175 B.n141 VSUBS 0.008272f
C176 B.n142 VSUBS 0.008272f
C177 B.n143 VSUBS 0.008272f
C178 B.n144 VSUBS 0.008272f
C179 B.n145 VSUBS 0.008272f
C180 B.n146 VSUBS 0.008272f
C181 B.n147 VSUBS 0.008272f
C182 B.n148 VSUBS 0.008272f
C183 B.n149 VSUBS 0.008272f
C184 B.n150 VSUBS 0.008272f
C185 B.n151 VSUBS 0.008272f
C186 B.n152 VSUBS 0.008272f
C187 B.n153 VSUBS 0.008272f
C188 B.t2 VSUBS 0.151179f
C189 B.t1 VSUBS 0.194491f
C190 B.t0 VSUBS 1.58765f
C191 B.n154 VSUBS 0.316862f
C192 B.n155 VSUBS 0.231949f
C193 B.n156 VSUBS 0.008272f
C194 B.n157 VSUBS 0.008272f
C195 B.n158 VSUBS 0.008272f
C196 B.n159 VSUBS 0.008272f
C197 B.n160 VSUBS 0.004622f
C198 B.n161 VSUBS 0.008272f
C199 B.n162 VSUBS 0.008272f
C200 B.n163 VSUBS 0.008272f
C201 B.n164 VSUBS 0.008272f
C202 B.n165 VSUBS 0.008272f
C203 B.n166 VSUBS 0.008272f
C204 B.n167 VSUBS 0.008272f
C205 B.n168 VSUBS 0.008272f
C206 B.n169 VSUBS 0.008272f
C207 B.n170 VSUBS 0.008272f
C208 B.n171 VSUBS 0.008272f
C209 B.n172 VSUBS 0.008272f
C210 B.n173 VSUBS 0.008272f
C211 B.n174 VSUBS 0.008272f
C212 B.n175 VSUBS 0.020255f
C213 B.n176 VSUBS 0.008272f
C214 B.n177 VSUBS 0.008272f
C215 B.n178 VSUBS 0.008272f
C216 B.n179 VSUBS 0.008272f
C217 B.n180 VSUBS 0.008272f
C218 B.n181 VSUBS 0.008272f
C219 B.n182 VSUBS 0.008272f
C220 B.n183 VSUBS 0.008272f
C221 B.n184 VSUBS 0.008272f
C222 B.n185 VSUBS 0.008272f
C223 B.n186 VSUBS 0.008272f
C224 B.n187 VSUBS 0.008272f
C225 B.n188 VSUBS 0.008272f
C226 B.n189 VSUBS 0.008272f
C227 B.n190 VSUBS 0.008272f
C228 B.n191 VSUBS 0.008272f
C229 B.n192 VSUBS 0.008272f
C230 B.n193 VSUBS 0.008272f
C231 B.n194 VSUBS 0.008272f
C232 B.n195 VSUBS 0.008272f
C233 B.n196 VSUBS 0.008272f
C234 B.n197 VSUBS 0.008272f
C235 B.n198 VSUBS 0.008272f
C236 B.n199 VSUBS 0.008272f
C237 B.n200 VSUBS 0.008272f
C238 B.n201 VSUBS 0.008272f
C239 B.n202 VSUBS 0.008272f
C240 B.n203 VSUBS 0.008272f
C241 B.n204 VSUBS 0.008272f
C242 B.n205 VSUBS 0.008272f
C243 B.n206 VSUBS 0.008272f
C244 B.n207 VSUBS 0.008272f
C245 B.n208 VSUBS 0.008272f
C246 B.n209 VSUBS 0.008272f
C247 B.n210 VSUBS 0.008272f
C248 B.n211 VSUBS 0.008272f
C249 B.n212 VSUBS 0.008272f
C250 B.n213 VSUBS 0.008272f
C251 B.n214 VSUBS 0.008272f
C252 B.n215 VSUBS 0.008272f
C253 B.n216 VSUBS 0.008272f
C254 B.n217 VSUBS 0.008272f
C255 B.n218 VSUBS 0.008272f
C256 B.n219 VSUBS 0.008272f
C257 B.n220 VSUBS 0.008272f
C258 B.n221 VSUBS 0.008272f
C259 B.n222 VSUBS 0.008272f
C260 B.n223 VSUBS 0.008272f
C261 B.n224 VSUBS 0.008272f
C262 B.n225 VSUBS 0.008272f
C263 B.n226 VSUBS 0.008272f
C264 B.n227 VSUBS 0.008272f
C265 B.n228 VSUBS 0.008272f
C266 B.n229 VSUBS 0.008272f
C267 B.n230 VSUBS 0.008272f
C268 B.n231 VSUBS 0.008272f
C269 B.n232 VSUBS 0.008272f
C270 B.n233 VSUBS 0.008272f
C271 B.n234 VSUBS 0.008272f
C272 B.n235 VSUBS 0.008272f
C273 B.n236 VSUBS 0.008272f
C274 B.n237 VSUBS 0.008272f
C275 B.n238 VSUBS 0.008272f
C276 B.n239 VSUBS 0.008272f
C277 B.n240 VSUBS 0.008272f
C278 B.n241 VSUBS 0.008272f
C279 B.n242 VSUBS 0.008272f
C280 B.n243 VSUBS 0.008272f
C281 B.n244 VSUBS 0.008272f
C282 B.n245 VSUBS 0.008272f
C283 B.n246 VSUBS 0.008272f
C284 B.n247 VSUBS 0.008272f
C285 B.n248 VSUBS 0.008272f
C286 B.n249 VSUBS 0.008272f
C287 B.n250 VSUBS 0.008272f
C288 B.n251 VSUBS 0.008272f
C289 B.n252 VSUBS 0.008272f
C290 B.n253 VSUBS 0.008272f
C291 B.n254 VSUBS 0.008272f
C292 B.n255 VSUBS 0.008272f
C293 B.n256 VSUBS 0.008272f
C294 B.n257 VSUBS 0.008272f
C295 B.n258 VSUBS 0.008272f
C296 B.n259 VSUBS 0.008272f
C297 B.n260 VSUBS 0.008272f
C298 B.n261 VSUBS 0.008272f
C299 B.n262 VSUBS 0.008272f
C300 B.n263 VSUBS 0.008272f
C301 B.n264 VSUBS 0.008272f
C302 B.n265 VSUBS 0.008272f
C303 B.n266 VSUBS 0.008272f
C304 B.n267 VSUBS 0.008272f
C305 B.n268 VSUBS 0.008272f
C306 B.n269 VSUBS 0.008272f
C307 B.n270 VSUBS 0.008272f
C308 B.n271 VSUBS 0.008272f
C309 B.n272 VSUBS 0.008272f
C310 B.n273 VSUBS 0.008272f
C311 B.n274 VSUBS 0.008272f
C312 B.n275 VSUBS 0.008272f
C313 B.n276 VSUBS 0.008272f
C314 B.n277 VSUBS 0.008272f
C315 B.n278 VSUBS 0.008272f
C316 B.n279 VSUBS 0.008272f
C317 B.n280 VSUBS 0.008272f
C318 B.n281 VSUBS 0.008272f
C319 B.n282 VSUBS 0.008272f
C320 B.n283 VSUBS 0.008272f
C321 B.n284 VSUBS 0.008272f
C322 B.n285 VSUBS 0.008272f
C323 B.n286 VSUBS 0.008272f
C324 B.n287 VSUBS 0.008272f
C325 B.n288 VSUBS 0.008272f
C326 B.n289 VSUBS 0.008272f
C327 B.n290 VSUBS 0.008272f
C328 B.n291 VSUBS 0.008272f
C329 B.n292 VSUBS 0.008272f
C330 B.n293 VSUBS 0.008272f
C331 B.n294 VSUBS 0.008272f
C332 B.n295 VSUBS 0.008272f
C333 B.n296 VSUBS 0.008272f
C334 B.n297 VSUBS 0.008272f
C335 B.n298 VSUBS 0.008272f
C336 B.n299 VSUBS 0.008272f
C337 B.n300 VSUBS 0.018671f
C338 B.n301 VSUBS 0.018671f
C339 B.n302 VSUBS 0.020255f
C340 B.n303 VSUBS 0.008272f
C341 B.n304 VSUBS 0.008272f
C342 B.n305 VSUBS 0.008272f
C343 B.n306 VSUBS 0.008272f
C344 B.n307 VSUBS 0.008272f
C345 B.n308 VSUBS 0.008272f
C346 B.n309 VSUBS 0.008272f
C347 B.n310 VSUBS 0.008272f
C348 B.n311 VSUBS 0.008272f
C349 B.n312 VSUBS 0.008272f
C350 B.n313 VSUBS 0.008272f
C351 B.n314 VSUBS 0.008272f
C352 B.n315 VSUBS 0.008272f
C353 B.n316 VSUBS 0.008272f
C354 B.n317 VSUBS 0.008272f
C355 B.n318 VSUBS 0.008272f
C356 B.n319 VSUBS 0.008272f
C357 B.n320 VSUBS 0.008272f
C358 B.n321 VSUBS 0.008272f
C359 B.n322 VSUBS 0.008272f
C360 B.n323 VSUBS 0.008272f
C361 B.n324 VSUBS 0.008272f
C362 B.n325 VSUBS 0.008272f
C363 B.n326 VSUBS 0.008272f
C364 B.n327 VSUBS 0.008272f
C365 B.n328 VSUBS 0.008272f
C366 B.n329 VSUBS 0.008272f
C367 B.n330 VSUBS 0.008272f
C368 B.n331 VSUBS 0.008272f
C369 B.n332 VSUBS 0.008272f
C370 B.n333 VSUBS 0.008272f
C371 B.n334 VSUBS 0.008272f
C372 B.n335 VSUBS 0.008272f
C373 B.n336 VSUBS 0.008272f
C374 B.n337 VSUBS 0.008272f
C375 B.n338 VSUBS 0.008272f
C376 B.n339 VSUBS 0.008272f
C377 B.n340 VSUBS 0.008272f
C378 B.n341 VSUBS 0.008272f
C379 B.n342 VSUBS 0.008272f
C380 B.n343 VSUBS 0.008272f
C381 B.n344 VSUBS 0.008272f
C382 B.t5 VSUBS 0.151176f
C383 B.t4 VSUBS 0.194489f
C384 B.t3 VSUBS 1.58765f
C385 B.n345 VSUBS 0.316864f
C386 B.n346 VSUBS 0.231951f
C387 B.n347 VSUBS 0.019165f
C388 B.n348 VSUBS 0.007785f
C389 B.n349 VSUBS 0.008272f
C390 B.n350 VSUBS 0.008272f
C391 B.n351 VSUBS 0.008272f
C392 B.n352 VSUBS 0.008272f
C393 B.n353 VSUBS 0.008272f
C394 B.n354 VSUBS 0.008272f
C395 B.n355 VSUBS 0.008272f
C396 B.n356 VSUBS 0.008272f
C397 B.n357 VSUBS 0.008272f
C398 B.n358 VSUBS 0.008272f
C399 B.n359 VSUBS 0.008272f
C400 B.n360 VSUBS 0.008272f
C401 B.n361 VSUBS 0.008272f
C402 B.n362 VSUBS 0.008272f
C403 B.n363 VSUBS 0.008272f
C404 B.n364 VSUBS 0.004622f
C405 B.n365 VSUBS 0.019165f
C406 B.n366 VSUBS 0.007785f
C407 B.n367 VSUBS 0.008272f
C408 B.n368 VSUBS 0.008272f
C409 B.n369 VSUBS 0.008272f
C410 B.n370 VSUBS 0.008272f
C411 B.n371 VSUBS 0.008272f
C412 B.n372 VSUBS 0.008272f
C413 B.n373 VSUBS 0.008272f
C414 B.n374 VSUBS 0.008272f
C415 B.n375 VSUBS 0.008272f
C416 B.n376 VSUBS 0.008272f
C417 B.n377 VSUBS 0.008272f
C418 B.n378 VSUBS 0.008272f
C419 B.n379 VSUBS 0.008272f
C420 B.n380 VSUBS 0.008272f
C421 B.n381 VSUBS 0.008272f
C422 B.n382 VSUBS 0.008272f
C423 B.n383 VSUBS 0.008272f
C424 B.n384 VSUBS 0.008272f
C425 B.n385 VSUBS 0.008272f
C426 B.n386 VSUBS 0.008272f
C427 B.n387 VSUBS 0.008272f
C428 B.n388 VSUBS 0.008272f
C429 B.n389 VSUBS 0.008272f
C430 B.n390 VSUBS 0.008272f
C431 B.n391 VSUBS 0.008272f
C432 B.n392 VSUBS 0.008272f
C433 B.n393 VSUBS 0.008272f
C434 B.n394 VSUBS 0.008272f
C435 B.n395 VSUBS 0.008272f
C436 B.n396 VSUBS 0.008272f
C437 B.n397 VSUBS 0.008272f
C438 B.n398 VSUBS 0.008272f
C439 B.n399 VSUBS 0.008272f
C440 B.n400 VSUBS 0.008272f
C441 B.n401 VSUBS 0.008272f
C442 B.n402 VSUBS 0.008272f
C443 B.n403 VSUBS 0.008272f
C444 B.n404 VSUBS 0.008272f
C445 B.n405 VSUBS 0.008272f
C446 B.n406 VSUBS 0.008272f
C447 B.n407 VSUBS 0.008272f
C448 B.n408 VSUBS 0.008272f
C449 B.n409 VSUBS 0.019286f
C450 B.n410 VSUBS 0.020255f
C451 B.n411 VSUBS 0.018671f
C452 B.n412 VSUBS 0.008272f
C453 B.n413 VSUBS 0.008272f
C454 B.n414 VSUBS 0.008272f
C455 B.n415 VSUBS 0.008272f
C456 B.n416 VSUBS 0.008272f
C457 B.n417 VSUBS 0.008272f
C458 B.n418 VSUBS 0.008272f
C459 B.n419 VSUBS 0.008272f
C460 B.n420 VSUBS 0.008272f
C461 B.n421 VSUBS 0.008272f
C462 B.n422 VSUBS 0.008272f
C463 B.n423 VSUBS 0.008272f
C464 B.n424 VSUBS 0.008272f
C465 B.n425 VSUBS 0.008272f
C466 B.n426 VSUBS 0.008272f
C467 B.n427 VSUBS 0.008272f
C468 B.n428 VSUBS 0.008272f
C469 B.n429 VSUBS 0.008272f
C470 B.n430 VSUBS 0.008272f
C471 B.n431 VSUBS 0.008272f
C472 B.n432 VSUBS 0.008272f
C473 B.n433 VSUBS 0.008272f
C474 B.n434 VSUBS 0.008272f
C475 B.n435 VSUBS 0.008272f
C476 B.n436 VSUBS 0.008272f
C477 B.n437 VSUBS 0.008272f
C478 B.n438 VSUBS 0.008272f
C479 B.n439 VSUBS 0.008272f
C480 B.n440 VSUBS 0.008272f
C481 B.n441 VSUBS 0.008272f
C482 B.n442 VSUBS 0.008272f
C483 B.n443 VSUBS 0.008272f
C484 B.n444 VSUBS 0.008272f
C485 B.n445 VSUBS 0.008272f
C486 B.n446 VSUBS 0.008272f
C487 B.n447 VSUBS 0.008272f
C488 B.n448 VSUBS 0.008272f
C489 B.n449 VSUBS 0.008272f
C490 B.n450 VSUBS 0.008272f
C491 B.n451 VSUBS 0.008272f
C492 B.n452 VSUBS 0.008272f
C493 B.n453 VSUBS 0.008272f
C494 B.n454 VSUBS 0.008272f
C495 B.n455 VSUBS 0.008272f
C496 B.n456 VSUBS 0.008272f
C497 B.n457 VSUBS 0.008272f
C498 B.n458 VSUBS 0.008272f
C499 B.n459 VSUBS 0.008272f
C500 B.n460 VSUBS 0.008272f
C501 B.n461 VSUBS 0.008272f
C502 B.n462 VSUBS 0.008272f
C503 B.n463 VSUBS 0.008272f
C504 B.n464 VSUBS 0.008272f
C505 B.n465 VSUBS 0.008272f
C506 B.n466 VSUBS 0.008272f
C507 B.n467 VSUBS 0.008272f
C508 B.n468 VSUBS 0.008272f
C509 B.n469 VSUBS 0.008272f
C510 B.n470 VSUBS 0.008272f
C511 B.n471 VSUBS 0.008272f
C512 B.n472 VSUBS 0.008272f
C513 B.n473 VSUBS 0.008272f
C514 B.n474 VSUBS 0.008272f
C515 B.n475 VSUBS 0.008272f
C516 B.n476 VSUBS 0.008272f
C517 B.n477 VSUBS 0.008272f
C518 B.n478 VSUBS 0.008272f
C519 B.n479 VSUBS 0.008272f
C520 B.n480 VSUBS 0.008272f
C521 B.n481 VSUBS 0.008272f
C522 B.n482 VSUBS 0.008272f
C523 B.n483 VSUBS 0.008272f
C524 B.n484 VSUBS 0.008272f
C525 B.n485 VSUBS 0.008272f
C526 B.n486 VSUBS 0.008272f
C527 B.n487 VSUBS 0.008272f
C528 B.n488 VSUBS 0.008272f
C529 B.n489 VSUBS 0.008272f
C530 B.n490 VSUBS 0.008272f
C531 B.n491 VSUBS 0.008272f
C532 B.n492 VSUBS 0.008272f
C533 B.n493 VSUBS 0.008272f
C534 B.n494 VSUBS 0.008272f
C535 B.n495 VSUBS 0.008272f
C536 B.n496 VSUBS 0.008272f
C537 B.n497 VSUBS 0.008272f
C538 B.n498 VSUBS 0.008272f
C539 B.n499 VSUBS 0.008272f
C540 B.n500 VSUBS 0.008272f
C541 B.n501 VSUBS 0.008272f
C542 B.n502 VSUBS 0.008272f
C543 B.n503 VSUBS 0.008272f
C544 B.n504 VSUBS 0.008272f
C545 B.n505 VSUBS 0.008272f
C546 B.n506 VSUBS 0.008272f
C547 B.n507 VSUBS 0.008272f
C548 B.n508 VSUBS 0.008272f
C549 B.n509 VSUBS 0.008272f
C550 B.n510 VSUBS 0.008272f
C551 B.n511 VSUBS 0.008272f
C552 B.n512 VSUBS 0.008272f
C553 B.n513 VSUBS 0.008272f
C554 B.n514 VSUBS 0.008272f
C555 B.n515 VSUBS 0.008272f
C556 B.n516 VSUBS 0.008272f
C557 B.n517 VSUBS 0.008272f
C558 B.n518 VSUBS 0.008272f
C559 B.n519 VSUBS 0.008272f
C560 B.n520 VSUBS 0.008272f
C561 B.n521 VSUBS 0.008272f
C562 B.n522 VSUBS 0.008272f
C563 B.n523 VSUBS 0.008272f
C564 B.n524 VSUBS 0.008272f
C565 B.n525 VSUBS 0.008272f
C566 B.n526 VSUBS 0.008272f
C567 B.n527 VSUBS 0.008272f
C568 B.n528 VSUBS 0.008272f
C569 B.n529 VSUBS 0.008272f
C570 B.n530 VSUBS 0.008272f
C571 B.n531 VSUBS 0.008272f
C572 B.n532 VSUBS 0.008272f
C573 B.n533 VSUBS 0.008272f
C574 B.n534 VSUBS 0.008272f
C575 B.n535 VSUBS 0.008272f
C576 B.n536 VSUBS 0.008272f
C577 B.n537 VSUBS 0.008272f
C578 B.n538 VSUBS 0.008272f
C579 B.n539 VSUBS 0.008272f
C580 B.n540 VSUBS 0.008272f
C581 B.n541 VSUBS 0.008272f
C582 B.n542 VSUBS 0.008272f
C583 B.n543 VSUBS 0.008272f
C584 B.n544 VSUBS 0.008272f
C585 B.n545 VSUBS 0.008272f
C586 B.n546 VSUBS 0.008272f
C587 B.n547 VSUBS 0.008272f
C588 B.n548 VSUBS 0.008272f
C589 B.n549 VSUBS 0.008272f
C590 B.n550 VSUBS 0.008272f
C591 B.n551 VSUBS 0.008272f
C592 B.n552 VSUBS 0.008272f
C593 B.n553 VSUBS 0.008272f
C594 B.n554 VSUBS 0.008272f
C595 B.n555 VSUBS 0.008272f
C596 B.n556 VSUBS 0.008272f
C597 B.n557 VSUBS 0.008272f
C598 B.n558 VSUBS 0.008272f
C599 B.n559 VSUBS 0.008272f
C600 B.n560 VSUBS 0.008272f
C601 B.n561 VSUBS 0.008272f
C602 B.n562 VSUBS 0.008272f
C603 B.n563 VSUBS 0.008272f
C604 B.n564 VSUBS 0.008272f
C605 B.n565 VSUBS 0.008272f
C606 B.n566 VSUBS 0.008272f
C607 B.n567 VSUBS 0.008272f
C608 B.n568 VSUBS 0.008272f
C609 B.n569 VSUBS 0.008272f
C610 B.n570 VSUBS 0.008272f
C611 B.n571 VSUBS 0.008272f
C612 B.n572 VSUBS 0.008272f
C613 B.n573 VSUBS 0.008272f
C614 B.n574 VSUBS 0.008272f
C615 B.n575 VSUBS 0.008272f
C616 B.n576 VSUBS 0.008272f
C617 B.n577 VSUBS 0.008272f
C618 B.n578 VSUBS 0.008272f
C619 B.n579 VSUBS 0.008272f
C620 B.n580 VSUBS 0.008272f
C621 B.n581 VSUBS 0.008272f
C622 B.n582 VSUBS 0.008272f
C623 B.n583 VSUBS 0.008272f
C624 B.n584 VSUBS 0.008272f
C625 B.n585 VSUBS 0.008272f
C626 B.n586 VSUBS 0.008272f
C627 B.n587 VSUBS 0.008272f
C628 B.n588 VSUBS 0.008272f
C629 B.n589 VSUBS 0.008272f
C630 B.n590 VSUBS 0.008272f
C631 B.n591 VSUBS 0.008272f
C632 B.n592 VSUBS 0.008272f
C633 B.n593 VSUBS 0.008272f
C634 B.n594 VSUBS 0.008272f
C635 B.n595 VSUBS 0.008272f
C636 B.n596 VSUBS 0.008272f
C637 B.n597 VSUBS 0.008272f
C638 B.n598 VSUBS 0.008272f
C639 B.n599 VSUBS 0.008272f
C640 B.n600 VSUBS 0.008272f
C641 B.n601 VSUBS 0.008272f
C642 B.n602 VSUBS 0.008272f
C643 B.n603 VSUBS 0.008272f
C644 B.n604 VSUBS 0.018671f
C645 B.n605 VSUBS 0.018671f
C646 B.n606 VSUBS 0.020255f
C647 B.n607 VSUBS 0.008272f
C648 B.n608 VSUBS 0.008272f
C649 B.n609 VSUBS 0.008272f
C650 B.n610 VSUBS 0.008272f
C651 B.n611 VSUBS 0.008272f
C652 B.n612 VSUBS 0.008272f
C653 B.n613 VSUBS 0.008272f
C654 B.n614 VSUBS 0.008272f
C655 B.n615 VSUBS 0.008272f
C656 B.n616 VSUBS 0.008272f
C657 B.n617 VSUBS 0.008272f
C658 B.n618 VSUBS 0.008272f
C659 B.n619 VSUBS 0.008272f
C660 B.n620 VSUBS 0.008272f
C661 B.n621 VSUBS 0.008272f
C662 B.n622 VSUBS 0.008272f
C663 B.n623 VSUBS 0.008272f
C664 B.n624 VSUBS 0.008272f
C665 B.n625 VSUBS 0.008272f
C666 B.n626 VSUBS 0.008272f
C667 B.n627 VSUBS 0.008272f
C668 B.n628 VSUBS 0.008272f
C669 B.n629 VSUBS 0.008272f
C670 B.n630 VSUBS 0.008272f
C671 B.n631 VSUBS 0.008272f
C672 B.n632 VSUBS 0.008272f
C673 B.n633 VSUBS 0.008272f
C674 B.n634 VSUBS 0.008272f
C675 B.n635 VSUBS 0.008272f
C676 B.n636 VSUBS 0.008272f
C677 B.n637 VSUBS 0.008272f
C678 B.n638 VSUBS 0.008272f
C679 B.n639 VSUBS 0.008272f
C680 B.n640 VSUBS 0.008272f
C681 B.n641 VSUBS 0.008272f
C682 B.n642 VSUBS 0.008272f
C683 B.n643 VSUBS 0.008272f
C684 B.n644 VSUBS 0.008272f
C685 B.n645 VSUBS 0.008272f
C686 B.n646 VSUBS 0.008272f
C687 B.n647 VSUBS 0.008272f
C688 B.n648 VSUBS 0.008272f
C689 B.n649 VSUBS 0.007785f
C690 B.n650 VSUBS 0.008272f
C691 B.n651 VSUBS 0.008272f
C692 B.n652 VSUBS 0.004622f
C693 B.n653 VSUBS 0.008272f
C694 B.n654 VSUBS 0.008272f
C695 B.n655 VSUBS 0.008272f
C696 B.n656 VSUBS 0.008272f
C697 B.n657 VSUBS 0.008272f
C698 B.n658 VSUBS 0.008272f
C699 B.n659 VSUBS 0.008272f
C700 B.n660 VSUBS 0.008272f
C701 B.n661 VSUBS 0.008272f
C702 B.n662 VSUBS 0.008272f
C703 B.n663 VSUBS 0.008272f
C704 B.n664 VSUBS 0.008272f
C705 B.n665 VSUBS 0.004622f
C706 B.n666 VSUBS 0.019165f
C707 B.n667 VSUBS 0.007785f
C708 B.n668 VSUBS 0.008272f
C709 B.n669 VSUBS 0.008272f
C710 B.n670 VSUBS 0.008272f
C711 B.n671 VSUBS 0.008272f
C712 B.n672 VSUBS 0.008272f
C713 B.n673 VSUBS 0.008272f
C714 B.n674 VSUBS 0.008272f
C715 B.n675 VSUBS 0.008272f
C716 B.n676 VSUBS 0.008272f
C717 B.n677 VSUBS 0.008272f
C718 B.n678 VSUBS 0.008272f
C719 B.n679 VSUBS 0.008272f
C720 B.n680 VSUBS 0.008272f
C721 B.n681 VSUBS 0.008272f
C722 B.n682 VSUBS 0.008272f
C723 B.n683 VSUBS 0.008272f
C724 B.n684 VSUBS 0.008272f
C725 B.n685 VSUBS 0.008272f
C726 B.n686 VSUBS 0.008272f
C727 B.n687 VSUBS 0.008272f
C728 B.n688 VSUBS 0.008272f
C729 B.n689 VSUBS 0.008272f
C730 B.n690 VSUBS 0.008272f
C731 B.n691 VSUBS 0.008272f
C732 B.n692 VSUBS 0.008272f
C733 B.n693 VSUBS 0.008272f
C734 B.n694 VSUBS 0.008272f
C735 B.n695 VSUBS 0.008272f
C736 B.n696 VSUBS 0.008272f
C737 B.n697 VSUBS 0.008272f
C738 B.n698 VSUBS 0.008272f
C739 B.n699 VSUBS 0.008272f
C740 B.n700 VSUBS 0.008272f
C741 B.n701 VSUBS 0.008272f
C742 B.n702 VSUBS 0.008272f
C743 B.n703 VSUBS 0.008272f
C744 B.n704 VSUBS 0.008272f
C745 B.n705 VSUBS 0.008272f
C746 B.n706 VSUBS 0.008272f
C747 B.n707 VSUBS 0.008272f
C748 B.n708 VSUBS 0.008272f
C749 B.n709 VSUBS 0.008272f
C750 B.n710 VSUBS 0.008272f
C751 B.n711 VSUBS 0.020255f
C752 B.n712 VSUBS 0.018671f
C753 B.n713 VSUBS 0.018671f
C754 B.n714 VSUBS 0.008272f
C755 B.n715 VSUBS 0.008272f
C756 B.n716 VSUBS 0.008272f
C757 B.n717 VSUBS 0.008272f
C758 B.n718 VSUBS 0.008272f
C759 B.n719 VSUBS 0.008272f
C760 B.n720 VSUBS 0.008272f
C761 B.n721 VSUBS 0.008272f
C762 B.n722 VSUBS 0.008272f
C763 B.n723 VSUBS 0.008272f
C764 B.n724 VSUBS 0.008272f
C765 B.n725 VSUBS 0.008272f
C766 B.n726 VSUBS 0.008272f
C767 B.n727 VSUBS 0.008272f
C768 B.n728 VSUBS 0.008272f
C769 B.n729 VSUBS 0.008272f
C770 B.n730 VSUBS 0.008272f
C771 B.n731 VSUBS 0.008272f
C772 B.n732 VSUBS 0.008272f
C773 B.n733 VSUBS 0.008272f
C774 B.n734 VSUBS 0.008272f
C775 B.n735 VSUBS 0.008272f
C776 B.n736 VSUBS 0.008272f
C777 B.n737 VSUBS 0.008272f
C778 B.n738 VSUBS 0.008272f
C779 B.n739 VSUBS 0.008272f
C780 B.n740 VSUBS 0.008272f
C781 B.n741 VSUBS 0.008272f
C782 B.n742 VSUBS 0.008272f
C783 B.n743 VSUBS 0.008272f
C784 B.n744 VSUBS 0.008272f
C785 B.n745 VSUBS 0.008272f
C786 B.n746 VSUBS 0.008272f
C787 B.n747 VSUBS 0.008272f
C788 B.n748 VSUBS 0.008272f
C789 B.n749 VSUBS 0.008272f
C790 B.n750 VSUBS 0.008272f
C791 B.n751 VSUBS 0.008272f
C792 B.n752 VSUBS 0.008272f
C793 B.n753 VSUBS 0.008272f
C794 B.n754 VSUBS 0.008272f
C795 B.n755 VSUBS 0.008272f
C796 B.n756 VSUBS 0.008272f
C797 B.n757 VSUBS 0.008272f
C798 B.n758 VSUBS 0.008272f
C799 B.n759 VSUBS 0.008272f
C800 B.n760 VSUBS 0.008272f
C801 B.n761 VSUBS 0.008272f
C802 B.n762 VSUBS 0.008272f
C803 B.n763 VSUBS 0.008272f
C804 B.n764 VSUBS 0.008272f
C805 B.n765 VSUBS 0.008272f
C806 B.n766 VSUBS 0.008272f
C807 B.n767 VSUBS 0.008272f
C808 B.n768 VSUBS 0.008272f
C809 B.n769 VSUBS 0.008272f
C810 B.n770 VSUBS 0.008272f
C811 B.n771 VSUBS 0.008272f
C812 B.n772 VSUBS 0.008272f
C813 B.n773 VSUBS 0.008272f
C814 B.n774 VSUBS 0.008272f
C815 B.n775 VSUBS 0.008272f
C816 B.n776 VSUBS 0.008272f
C817 B.n777 VSUBS 0.008272f
C818 B.n778 VSUBS 0.008272f
C819 B.n779 VSUBS 0.008272f
C820 B.n780 VSUBS 0.008272f
C821 B.n781 VSUBS 0.008272f
C822 B.n782 VSUBS 0.008272f
C823 B.n783 VSUBS 0.008272f
C824 B.n784 VSUBS 0.008272f
C825 B.n785 VSUBS 0.008272f
C826 B.n786 VSUBS 0.008272f
C827 B.n787 VSUBS 0.008272f
C828 B.n788 VSUBS 0.008272f
C829 B.n789 VSUBS 0.008272f
C830 B.n790 VSUBS 0.008272f
C831 B.n791 VSUBS 0.008272f
C832 B.n792 VSUBS 0.008272f
C833 B.n793 VSUBS 0.008272f
C834 B.n794 VSUBS 0.008272f
C835 B.n795 VSUBS 0.008272f
C836 B.n796 VSUBS 0.008272f
C837 B.n797 VSUBS 0.008272f
C838 B.n798 VSUBS 0.008272f
C839 B.n799 VSUBS 0.008272f
C840 B.n800 VSUBS 0.008272f
C841 B.n801 VSUBS 0.008272f
C842 B.n802 VSUBS 0.008272f
C843 B.n803 VSUBS 0.008272f
C844 B.n804 VSUBS 0.008272f
C845 B.n805 VSUBS 0.008272f
C846 B.n806 VSUBS 0.008272f
C847 B.n807 VSUBS 0.010794f
C848 B.n808 VSUBS 0.011499f
C849 B.n809 VSUBS 0.022866f
C850 VDD1.t0 VSUBS 0.205994f
C851 VDD1.t5 VSUBS 0.205994f
C852 VDD1.n0 VSUBS 1.48879f
C853 VDD1.t2 VSUBS 0.205994f
C854 VDD1.t1 VSUBS 0.205994f
C855 VDD1.n1 VSUBS 1.48706f
C856 VDD1.t3 VSUBS 0.205994f
C857 VDD1.t4 VSUBS 0.205994f
C858 VDD1.n2 VSUBS 1.48706f
C859 VDD1.n3 VSUBS 5.294641f
C860 VDD1.t7 VSUBS 0.205994f
C861 VDD1.t6 VSUBS 0.205994f
C862 VDD1.n4 VSUBS 1.4656f
C863 VDD1.n5 VSUBS 4.19152f
C864 VP.t3 VSUBS 2.42726f
C865 VP.n0 VSUBS 1.00466f
C866 VP.n1 VSUBS 0.031845f
C867 VP.n2 VSUBS 0.036434f
C868 VP.n3 VSUBS 0.031845f
C869 VP.n4 VSUBS 0.034616f
C870 VP.n5 VSUBS 0.031845f
C871 VP.n6 VSUBS 0.02577f
C872 VP.n7 VSUBS 0.031845f
C873 VP.t6 VSUBS 2.42726f
C874 VP.n8 VSUBS 0.873443f
C875 VP.n9 VSUBS 0.031845f
C876 VP.n10 VSUBS 0.055379f
C877 VP.n11 VSUBS 0.031845f
C878 VP.n12 VSUBS 0.046396f
C879 VP.t1 VSUBS 2.42726f
C880 VP.n13 VSUBS 1.00466f
C881 VP.n14 VSUBS 0.031845f
C882 VP.n15 VSUBS 0.036434f
C883 VP.n16 VSUBS 0.031845f
C884 VP.n17 VSUBS 0.034616f
C885 VP.n18 VSUBS 0.031845f
C886 VP.n19 VSUBS 0.02577f
C887 VP.n20 VSUBS 0.031845f
C888 VP.t2 VSUBS 2.42726f
C889 VP.n21 VSUBS 0.995785f
C890 VP.t7 VSUBS 2.85185f
C891 VP.n22 VSUBS 0.936972f
C892 VP.n23 VSUBS 0.392181f
C893 VP.n24 VSUBS 0.055231f
C894 VP.n25 VSUBS 0.059649f
C895 VP.n26 VSUBS 0.06363f
C896 VP.n27 VSUBS 0.031845f
C897 VP.n28 VSUBS 0.031845f
C898 VP.n29 VSUBS 0.031845f
C899 VP.n30 VSUBS 0.06363f
C900 VP.n31 VSUBS 0.059649f
C901 VP.t0 VSUBS 2.42726f
C902 VP.n32 VSUBS 0.873443f
C903 VP.n33 VSUBS 0.055231f
C904 VP.n34 VSUBS 0.031845f
C905 VP.n35 VSUBS 0.031845f
C906 VP.n36 VSUBS 0.031845f
C907 VP.n37 VSUBS 0.059649f
C908 VP.n38 VSUBS 0.059649f
C909 VP.n39 VSUBS 0.055379f
C910 VP.n40 VSUBS 0.031845f
C911 VP.n41 VSUBS 0.031845f
C912 VP.n42 VSUBS 0.031845f
C913 VP.n43 VSUBS 0.061216f
C914 VP.n44 VSUBS 0.059649f
C915 VP.n45 VSUBS 0.046396f
C916 VP.n46 VSUBS 0.051405f
C917 VP.n47 VSUBS 1.94126f
C918 VP.t5 VSUBS 2.42726f
C919 VP.n48 VSUBS 1.00466f
C920 VP.n49 VSUBS 1.96305f
C921 VP.n50 VSUBS 0.051405f
C922 VP.n51 VSUBS 0.031845f
C923 VP.n52 VSUBS 0.059649f
C924 VP.n53 VSUBS 0.061216f
C925 VP.n54 VSUBS 0.036434f
C926 VP.n55 VSUBS 0.031845f
C927 VP.n56 VSUBS 0.031845f
C928 VP.n57 VSUBS 0.031845f
C929 VP.n58 VSUBS 0.059649f
C930 VP.n59 VSUBS 0.059649f
C931 VP.n60 VSUBS 0.034616f
C932 VP.n61 VSUBS 0.031845f
C933 VP.n62 VSUBS 0.031845f
C934 VP.n63 VSUBS 0.055231f
C935 VP.n64 VSUBS 0.059649f
C936 VP.n65 VSUBS 0.06363f
C937 VP.n66 VSUBS 0.031845f
C938 VP.n67 VSUBS 0.031845f
C939 VP.n68 VSUBS 0.031845f
C940 VP.n69 VSUBS 0.06363f
C941 VP.n70 VSUBS 0.059649f
C942 VP.t4 VSUBS 2.42726f
C943 VP.n71 VSUBS 0.873443f
C944 VP.n72 VSUBS 0.055231f
C945 VP.n73 VSUBS 0.031845f
C946 VP.n74 VSUBS 0.031845f
C947 VP.n75 VSUBS 0.031845f
C948 VP.n76 VSUBS 0.059649f
C949 VP.n77 VSUBS 0.059649f
C950 VP.n78 VSUBS 0.055379f
C951 VP.n79 VSUBS 0.031845f
C952 VP.n80 VSUBS 0.031845f
C953 VP.n81 VSUBS 0.031845f
C954 VP.n82 VSUBS 0.061216f
C955 VP.n83 VSUBS 0.059649f
C956 VP.n84 VSUBS 0.046396f
C957 VP.n85 VSUBS 0.051405f
C958 VP.n86 VSUBS 0.081674f
C959 VDD2.t1 VSUBS 0.205092f
C960 VDD2.t2 VSUBS 0.205092f
C961 VDD2.n0 VSUBS 1.48055f
C962 VDD2.t4 VSUBS 0.205092f
C963 VDD2.t5 VSUBS 0.205092f
C964 VDD2.n1 VSUBS 1.48055f
C965 VDD2.n2 VSUBS 5.20485f
C966 VDD2.t6 VSUBS 0.205092f
C967 VDD2.t7 VSUBS 0.205092f
C968 VDD2.n3 VSUBS 1.45918f
C969 VDD2.n4 VSUBS 4.13289f
C970 VDD2.t0 VSUBS 0.205092f
C971 VDD2.t3 VSUBS 0.205092f
C972 VDD2.n5 VSUBS 1.4805f
C973 VTAIL.t14 VSUBS 0.179487f
C974 VTAIL.t12 VSUBS 0.179487f
C975 VTAIL.n0 VSUBS 1.14778f
C976 VTAIL.n1 VSUBS 0.900133f
C977 VTAIL.n2 VSUBS 0.031085f
C978 VTAIL.n3 VSUBS 0.02818f
C979 VTAIL.n4 VSUBS 0.015143f
C980 VTAIL.n5 VSUBS 0.035792f
C981 VTAIL.n6 VSUBS 0.016034f
C982 VTAIL.n7 VSUBS 0.02818f
C983 VTAIL.n8 VSUBS 0.015143f
C984 VTAIL.n9 VSUBS 0.035792f
C985 VTAIL.n10 VSUBS 0.016034f
C986 VTAIL.n11 VSUBS 0.02818f
C987 VTAIL.n12 VSUBS 0.015143f
C988 VTAIL.n13 VSUBS 0.035792f
C989 VTAIL.n14 VSUBS 0.016034f
C990 VTAIL.n15 VSUBS 0.141134f
C991 VTAIL.t8 VSUBS 0.076313f
C992 VTAIL.n16 VSUBS 0.026844f
C993 VTAIL.n17 VSUBS 0.022769f
C994 VTAIL.n18 VSUBS 0.015143f
C995 VTAIL.n19 VSUBS 0.911181f
C996 VTAIL.n20 VSUBS 0.02818f
C997 VTAIL.n21 VSUBS 0.015143f
C998 VTAIL.n22 VSUBS 0.016034f
C999 VTAIL.n23 VSUBS 0.035792f
C1000 VTAIL.n24 VSUBS 0.035792f
C1001 VTAIL.n25 VSUBS 0.016034f
C1002 VTAIL.n26 VSUBS 0.015143f
C1003 VTAIL.n27 VSUBS 0.02818f
C1004 VTAIL.n28 VSUBS 0.02818f
C1005 VTAIL.n29 VSUBS 0.015143f
C1006 VTAIL.n30 VSUBS 0.016034f
C1007 VTAIL.n31 VSUBS 0.035792f
C1008 VTAIL.n32 VSUBS 0.035792f
C1009 VTAIL.n33 VSUBS 0.016034f
C1010 VTAIL.n34 VSUBS 0.015143f
C1011 VTAIL.n35 VSUBS 0.02818f
C1012 VTAIL.n36 VSUBS 0.02818f
C1013 VTAIL.n37 VSUBS 0.015143f
C1014 VTAIL.n38 VSUBS 0.016034f
C1015 VTAIL.n39 VSUBS 0.035792f
C1016 VTAIL.n40 VSUBS 0.087062f
C1017 VTAIL.n41 VSUBS 0.016034f
C1018 VTAIL.n42 VSUBS 0.015143f
C1019 VTAIL.n43 VSUBS 0.061288f
C1020 VTAIL.n44 VSUBS 0.043679f
C1021 VTAIL.n45 VSUBS 0.365933f
C1022 VTAIL.n46 VSUBS 0.031085f
C1023 VTAIL.n47 VSUBS 0.02818f
C1024 VTAIL.n48 VSUBS 0.015143f
C1025 VTAIL.n49 VSUBS 0.035792f
C1026 VTAIL.n50 VSUBS 0.016034f
C1027 VTAIL.n51 VSUBS 0.02818f
C1028 VTAIL.n52 VSUBS 0.015143f
C1029 VTAIL.n53 VSUBS 0.035792f
C1030 VTAIL.n54 VSUBS 0.016034f
C1031 VTAIL.n55 VSUBS 0.02818f
C1032 VTAIL.n56 VSUBS 0.015143f
C1033 VTAIL.n57 VSUBS 0.035792f
C1034 VTAIL.n58 VSUBS 0.016034f
C1035 VTAIL.n59 VSUBS 0.141134f
C1036 VTAIL.t5 VSUBS 0.076313f
C1037 VTAIL.n60 VSUBS 0.026844f
C1038 VTAIL.n61 VSUBS 0.022769f
C1039 VTAIL.n62 VSUBS 0.015143f
C1040 VTAIL.n63 VSUBS 0.911181f
C1041 VTAIL.n64 VSUBS 0.02818f
C1042 VTAIL.n65 VSUBS 0.015143f
C1043 VTAIL.n66 VSUBS 0.016034f
C1044 VTAIL.n67 VSUBS 0.035792f
C1045 VTAIL.n68 VSUBS 0.035792f
C1046 VTAIL.n69 VSUBS 0.016034f
C1047 VTAIL.n70 VSUBS 0.015143f
C1048 VTAIL.n71 VSUBS 0.02818f
C1049 VTAIL.n72 VSUBS 0.02818f
C1050 VTAIL.n73 VSUBS 0.015143f
C1051 VTAIL.n74 VSUBS 0.016034f
C1052 VTAIL.n75 VSUBS 0.035792f
C1053 VTAIL.n76 VSUBS 0.035792f
C1054 VTAIL.n77 VSUBS 0.016034f
C1055 VTAIL.n78 VSUBS 0.015143f
C1056 VTAIL.n79 VSUBS 0.02818f
C1057 VTAIL.n80 VSUBS 0.02818f
C1058 VTAIL.n81 VSUBS 0.015143f
C1059 VTAIL.n82 VSUBS 0.016034f
C1060 VTAIL.n83 VSUBS 0.035792f
C1061 VTAIL.n84 VSUBS 0.087062f
C1062 VTAIL.n85 VSUBS 0.016034f
C1063 VTAIL.n86 VSUBS 0.015143f
C1064 VTAIL.n87 VSUBS 0.061288f
C1065 VTAIL.n88 VSUBS 0.043679f
C1066 VTAIL.n89 VSUBS 0.365933f
C1067 VTAIL.t4 VSUBS 0.179487f
C1068 VTAIL.t7 VSUBS 0.179487f
C1069 VTAIL.n90 VSUBS 1.14778f
C1070 VTAIL.n91 VSUBS 1.19622f
C1071 VTAIL.n92 VSUBS 0.031085f
C1072 VTAIL.n93 VSUBS 0.02818f
C1073 VTAIL.n94 VSUBS 0.015143f
C1074 VTAIL.n95 VSUBS 0.035792f
C1075 VTAIL.n96 VSUBS 0.016034f
C1076 VTAIL.n97 VSUBS 0.02818f
C1077 VTAIL.n98 VSUBS 0.015143f
C1078 VTAIL.n99 VSUBS 0.035792f
C1079 VTAIL.n100 VSUBS 0.016034f
C1080 VTAIL.n101 VSUBS 0.02818f
C1081 VTAIL.n102 VSUBS 0.015143f
C1082 VTAIL.n103 VSUBS 0.035792f
C1083 VTAIL.n104 VSUBS 0.016034f
C1084 VTAIL.n105 VSUBS 0.141134f
C1085 VTAIL.t0 VSUBS 0.076313f
C1086 VTAIL.n106 VSUBS 0.026844f
C1087 VTAIL.n107 VSUBS 0.022769f
C1088 VTAIL.n108 VSUBS 0.015143f
C1089 VTAIL.n109 VSUBS 0.911181f
C1090 VTAIL.n110 VSUBS 0.02818f
C1091 VTAIL.n111 VSUBS 0.015143f
C1092 VTAIL.n112 VSUBS 0.016034f
C1093 VTAIL.n113 VSUBS 0.035792f
C1094 VTAIL.n114 VSUBS 0.035792f
C1095 VTAIL.n115 VSUBS 0.016034f
C1096 VTAIL.n116 VSUBS 0.015143f
C1097 VTAIL.n117 VSUBS 0.02818f
C1098 VTAIL.n118 VSUBS 0.02818f
C1099 VTAIL.n119 VSUBS 0.015143f
C1100 VTAIL.n120 VSUBS 0.016034f
C1101 VTAIL.n121 VSUBS 0.035792f
C1102 VTAIL.n122 VSUBS 0.035792f
C1103 VTAIL.n123 VSUBS 0.016034f
C1104 VTAIL.n124 VSUBS 0.015143f
C1105 VTAIL.n125 VSUBS 0.02818f
C1106 VTAIL.n126 VSUBS 0.02818f
C1107 VTAIL.n127 VSUBS 0.015143f
C1108 VTAIL.n128 VSUBS 0.016034f
C1109 VTAIL.n129 VSUBS 0.035792f
C1110 VTAIL.n130 VSUBS 0.087062f
C1111 VTAIL.n131 VSUBS 0.016034f
C1112 VTAIL.n132 VSUBS 0.015143f
C1113 VTAIL.n133 VSUBS 0.061288f
C1114 VTAIL.n134 VSUBS 0.043679f
C1115 VTAIL.n135 VSUBS 1.63836f
C1116 VTAIL.n136 VSUBS 0.031085f
C1117 VTAIL.n137 VSUBS 0.02818f
C1118 VTAIL.n138 VSUBS 0.015143f
C1119 VTAIL.n139 VSUBS 0.035792f
C1120 VTAIL.n140 VSUBS 0.016034f
C1121 VTAIL.n141 VSUBS 0.02818f
C1122 VTAIL.n142 VSUBS 0.015143f
C1123 VTAIL.n143 VSUBS 0.035792f
C1124 VTAIL.n144 VSUBS 0.016034f
C1125 VTAIL.n145 VSUBS 0.02818f
C1126 VTAIL.n146 VSUBS 0.015143f
C1127 VTAIL.n147 VSUBS 0.035792f
C1128 VTAIL.n148 VSUBS 0.016034f
C1129 VTAIL.n149 VSUBS 0.141134f
C1130 VTAIL.t9 VSUBS 0.076313f
C1131 VTAIL.n150 VSUBS 0.026844f
C1132 VTAIL.n151 VSUBS 0.022769f
C1133 VTAIL.n152 VSUBS 0.015143f
C1134 VTAIL.n153 VSUBS 0.911181f
C1135 VTAIL.n154 VSUBS 0.02818f
C1136 VTAIL.n155 VSUBS 0.015143f
C1137 VTAIL.n156 VSUBS 0.016034f
C1138 VTAIL.n157 VSUBS 0.035792f
C1139 VTAIL.n158 VSUBS 0.035792f
C1140 VTAIL.n159 VSUBS 0.016034f
C1141 VTAIL.n160 VSUBS 0.015143f
C1142 VTAIL.n161 VSUBS 0.02818f
C1143 VTAIL.n162 VSUBS 0.02818f
C1144 VTAIL.n163 VSUBS 0.015143f
C1145 VTAIL.n164 VSUBS 0.016034f
C1146 VTAIL.n165 VSUBS 0.035792f
C1147 VTAIL.n166 VSUBS 0.035792f
C1148 VTAIL.n167 VSUBS 0.016034f
C1149 VTAIL.n168 VSUBS 0.015143f
C1150 VTAIL.n169 VSUBS 0.02818f
C1151 VTAIL.n170 VSUBS 0.02818f
C1152 VTAIL.n171 VSUBS 0.015143f
C1153 VTAIL.n172 VSUBS 0.016034f
C1154 VTAIL.n173 VSUBS 0.035792f
C1155 VTAIL.n174 VSUBS 0.087062f
C1156 VTAIL.n175 VSUBS 0.016034f
C1157 VTAIL.n176 VSUBS 0.015143f
C1158 VTAIL.n177 VSUBS 0.061288f
C1159 VTAIL.n178 VSUBS 0.043679f
C1160 VTAIL.n179 VSUBS 1.63837f
C1161 VTAIL.t13 VSUBS 0.179487f
C1162 VTAIL.t11 VSUBS 0.179487f
C1163 VTAIL.n180 VSUBS 1.14778f
C1164 VTAIL.n181 VSUBS 1.19621f
C1165 VTAIL.n182 VSUBS 0.031085f
C1166 VTAIL.n183 VSUBS 0.02818f
C1167 VTAIL.n184 VSUBS 0.015143f
C1168 VTAIL.n185 VSUBS 0.035792f
C1169 VTAIL.n186 VSUBS 0.016034f
C1170 VTAIL.n187 VSUBS 0.02818f
C1171 VTAIL.n188 VSUBS 0.015143f
C1172 VTAIL.n189 VSUBS 0.035792f
C1173 VTAIL.n190 VSUBS 0.016034f
C1174 VTAIL.n191 VSUBS 0.02818f
C1175 VTAIL.n192 VSUBS 0.015143f
C1176 VTAIL.n193 VSUBS 0.035792f
C1177 VTAIL.n194 VSUBS 0.016034f
C1178 VTAIL.n195 VSUBS 0.141134f
C1179 VTAIL.t15 VSUBS 0.076313f
C1180 VTAIL.n196 VSUBS 0.026844f
C1181 VTAIL.n197 VSUBS 0.022769f
C1182 VTAIL.n198 VSUBS 0.015143f
C1183 VTAIL.n199 VSUBS 0.911181f
C1184 VTAIL.n200 VSUBS 0.02818f
C1185 VTAIL.n201 VSUBS 0.015143f
C1186 VTAIL.n202 VSUBS 0.016034f
C1187 VTAIL.n203 VSUBS 0.035792f
C1188 VTAIL.n204 VSUBS 0.035792f
C1189 VTAIL.n205 VSUBS 0.016034f
C1190 VTAIL.n206 VSUBS 0.015143f
C1191 VTAIL.n207 VSUBS 0.02818f
C1192 VTAIL.n208 VSUBS 0.02818f
C1193 VTAIL.n209 VSUBS 0.015143f
C1194 VTAIL.n210 VSUBS 0.016034f
C1195 VTAIL.n211 VSUBS 0.035792f
C1196 VTAIL.n212 VSUBS 0.035792f
C1197 VTAIL.n213 VSUBS 0.016034f
C1198 VTAIL.n214 VSUBS 0.015143f
C1199 VTAIL.n215 VSUBS 0.02818f
C1200 VTAIL.n216 VSUBS 0.02818f
C1201 VTAIL.n217 VSUBS 0.015143f
C1202 VTAIL.n218 VSUBS 0.016034f
C1203 VTAIL.n219 VSUBS 0.035792f
C1204 VTAIL.n220 VSUBS 0.087062f
C1205 VTAIL.n221 VSUBS 0.016034f
C1206 VTAIL.n222 VSUBS 0.015143f
C1207 VTAIL.n223 VSUBS 0.061288f
C1208 VTAIL.n224 VSUBS 0.043679f
C1209 VTAIL.n225 VSUBS 0.365933f
C1210 VTAIL.n226 VSUBS 0.031085f
C1211 VTAIL.n227 VSUBS 0.02818f
C1212 VTAIL.n228 VSUBS 0.015143f
C1213 VTAIL.n229 VSUBS 0.035792f
C1214 VTAIL.n230 VSUBS 0.016034f
C1215 VTAIL.n231 VSUBS 0.02818f
C1216 VTAIL.n232 VSUBS 0.015143f
C1217 VTAIL.n233 VSUBS 0.035792f
C1218 VTAIL.n234 VSUBS 0.016034f
C1219 VTAIL.n235 VSUBS 0.02818f
C1220 VTAIL.n236 VSUBS 0.015143f
C1221 VTAIL.n237 VSUBS 0.035792f
C1222 VTAIL.n238 VSUBS 0.016034f
C1223 VTAIL.n239 VSUBS 0.141134f
C1224 VTAIL.t6 VSUBS 0.076313f
C1225 VTAIL.n240 VSUBS 0.026844f
C1226 VTAIL.n241 VSUBS 0.022769f
C1227 VTAIL.n242 VSUBS 0.015143f
C1228 VTAIL.n243 VSUBS 0.911181f
C1229 VTAIL.n244 VSUBS 0.02818f
C1230 VTAIL.n245 VSUBS 0.015143f
C1231 VTAIL.n246 VSUBS 0.016034f
C1232 VTAIL.n247 VSUBS 0.035792f
C1233 VTAIL.n248 VSUBS 0.035792f
C1234 VTAIL.n249 VSUBS 0.016034f
C1235 VTAIL.n250 VSUBS 0.015143f
C1236 VTAIL.n251 VSUBS 0.02818f
C1237 VTAIL.n252 VSUBS 0.02818f
C1238 VTAIL.n253 VSUBS 0.015143f
C1239 VTAIL.n254 VSUBS 0.016034f
C1240 VTAIL.n255 VSUBS 0.035792f
C1241 VTAIL.n256 VSUBS 0.035792f
C1242 VTAIL.n257 VSUBS 0.016034f
C1243 VTAIL.n258 VSUBS 0.015143f
C1244 VTAIL.n259 VSUBS 0.02818f
C1245 VTAIL.n260 VSUBS 0.02818f
C1246 VTAIL.n261 VSUBS 0.015143f
C1247 VTAIL.n262 VSUBS 0.016034f
C1248 VTAIL.n263 VSUBS 0.035792f
C1249 VTAIL.n264 VSUBS 0.087062f
C1250 VTAIL.n265 VSUBS 0.016034f
C1251 VTAIL.n266 VSUBS 0.015143f
C1252 VTAIL.n267 VSUBS 0.061288f
C1253 VTAIL.n268 VSUBS 0.043679f
C1254 VTAIL.n269 VSUBS 0.365933f
C1255 VTAIL.t2 VSUBS 0.179487f
C1256 VTAIL.t3 VSUBS 0.179487f
C1257 VTAIL.n270 VSUBS 1.14778f
C1258 VTAIL.n271 VSUBS 1.19621f
C1259 VTAIL.n272 VSUBS 0.031085f
C1260 VTAIL.n273 VSUBS 0.02818f
C1261 VTAIL.n274 VSUBS 0.015143f
C1262 VTAIL.n275 VSUBS 0.035792f
C1263 VTAIL.n276 VSUBS 0.016034f
C1264 VTAIL.n277 VSUBS 0.02818f
C1265 VTAIL.n278 VSUBS 0.015143f
C1266 VTAIL.n279 VSUBS 0.035792f
C1267 VTAIL.n280 VSUBS 0.016034f
C1268 VTAIL.n281 VSUBS 0.02818f
C1269 VTAIL.n282 VSUBS 0.015143f
C1270 VTAIL.n283 VSUBS 0.035792f
C1271 VTAIL.n284 VSUBS 0.016034f
C1272 VTAIL.n285 VSUBS 0.141134f
C1273 VTAIL.t1 VSUBS 0.076313f
C1274 VTAIL.n286 VSUBS 0.026844f
C1275 VTAIL.n287 VSUBS 0.022769f
C1276 VTAIL.n288 VSUBS 0.015143f
C1277 VTAIL.n289 VSUBS 0.911182f
C1278 VTAIL.n290 VSUBS 0.02818f
C1279 VTAIL.n291 VSUBS 0.015143f
C1280 VTAIL.n292 VSUBS 0.016034f
C1281 VTAIL.n293 VSUBS 0.035792f
C1282 VTAIL.n294 VSUBS 0.035792f
C1283 VTAIL.n295 VSUBS 0.016034f
C1284 VTAIL.n296 VSUBS 0.015143f
C1285 VTAIL.n297 VSUBS 0.02818f
C1286 VTAIL.n298 VSUBS 0.02818f
C1287 VTAIL.n299 VSUBS 0.015143f
C1288 VTAIL.n300 VSUBS 0.016034f
C1289 VTAIL.n301 VSUBS 0.035792f
C1290 VTAIL.n302 VSUBS 0.035792f
C1291 VTAIL.n303 VSUBS 0.016034f
C1292 VTAIL.n304 VSUBS 0.015143f
C1293 VTAIL.n305 VSUBS 0.02818f
C1294 VTAIL.n306 VSUBS 0.02818f
C1295 VTAIL.n307 VSUBS 0.015143f
C1296 VTAIL.n308 VSUBS 0.016034f
C1297 VTAIL.n309 VSUBS 0.035792f
C1298 VTAIL.n310 VSUBS 0.087062f
C1299 VTAIL.n311 VSUBS 0.016034f
C1300 VTAIL.n312 VSUBS 0.015143f
C1301 VTAIL.n313 VSUBS 0.061288f
C1302 VTAIL.n314 VSUBS 0.043679f
C1303 VTAIL.n315 VSUBS 1.63837f
C1304 VTAIL.n316 VSUBS 0.031085f
C1305 VTAIL.n317 VSUBS 0.02818f
C1306 VTAIL.n318 VSUBS 0.015143f
C1307 VTAIL.n319 VSUBS 0.035792f
C1308 VTAIL.n320 VSUBS 0.016034f
C1309 VTAIL.n321 VSUBS 0.02818f
C1310 VTAIL.n322 VSUBS 0.015143f
C1311 VTAIL.n323 VSUBS 0.035792f
C1312 VTAIL.n324 VSUBS 0.016034f
C1313 VTAIL.n325 VSUBS 0.02818f
C1314 VTAIL.n326 VSUBS 0.015143f
C1315 VTAIL.n327 VSUBS 0.035792f
C1316 VTAIL.n328 VSUBS 0.016034f
C1317 VTAIL.n329 VSUBS 0.141134f
C1318 VTAIL.t10 VSUBS 0.076313f
C1319 VTAIL.n330 VSUBS 0.026844f
C1320 VTAIL.n331 VSUBS 0.022769f
C1321 VTAIL.n332 VSUBS 0.015143f
C1322 VTAIL.n333 VSUBS 0.911181f
C1323 VTAIL.n334 VSUBS 0.02818f
C1324 VTAIL.n335 VSUBS 0.015143f
C1325 VTAIL.n336 VSUBS 0.016034f
C1326 VTAIL.n337 VSUBS 0.035792f
C1327 VTAIL.n338 VSUBS 0.035792f
C1328 VTAIL.n339 VSUBS 0.016034f
C1329 VTAIL.n340 VSUBS 0.015143f
C1330 VTAIL.n341 VSUBS 0.02818f
C1331 VTAIL.n342 VSUBS 0.02818f
C1332 VTAIL.n343 VSUBS 0.015143f
C1333 VTAIL.n344 VSUBS 0.016034f
C1334 VTAIL.n345 VSUBS 0.035792f
C1335 VTAIL.n346 VSUBS 0.035792f
C1336 VTAIL.n347 VSUBS 0.016034f
C1337 VTAIL.n348 VSUBS 0.015143f
C1338 VTAIL.n349 VSUBS 0.02818f
C1339 VTAIL.n350 VSUBS 0.02818f
C1340 VTAIL.n351 VSUBS 0.015143f
C1341 VTAIL.n352 VSUBS 0.016034f
C1342 VTAIL.n353 VSUBS 0.035792f
C1343 VTAIL.n354 VSUBS 0.087062f
C1344 VTAIL.n355 VSUBS 0.016034f
C1345 VTAIL.n356 VSUBS 0.015143f
C1346 VTAIL.n357 VSUBS 0.061288f
C1347 VTAIL.n358 VSUBS 0.043679f
C1348 VTAIL.n359 VSUBS 1.63308f
C1349 VN.t2 VSUBS 2.18245f
C1350 VN.n0 VSUBS 0.903325f
C1351 VN.n1 VSUBS 0.028633f
C1352 VN.n2 VSUBS 0.032759f
C1353 VN.n3 VSUBS 0.028633f
C1354 VN.n4 VSUBS 0.031124f
C1355 VN.n5 VSUBS 0.028633f
C1356 VN.n6 VSUBS 0.02317f
C1357 VN.n7 VSUBS 0.028633f
C1358 VN.t5 VSUBS 2.18245f
C1359 VN.n8 VSUBS 0.895348f
C1360 VN.t6 VSUBS 2.56421f
C1361 VN.n9 VSUBS 0.842466f
C1362 VN.n10 VSUBS 0.352625f
C1363 VN.n11 VSUBS 0.04966f
C1364 VN.n12 VSUBS 0.053632f
C1365 VN.n13 VSUBS 0.057212f
C1366 VN.n14 VSUBS 0.028633f
C1367 VN.n15 VSUBS 0.028633f
C1368 VN.n16 VSUBS 0.028633f
C1369 VN.n17 VSUBS 0.057212f
C1370 VN.n18 VSUBS 0.053632f
C1371 VN.t3 VSUBS 2.18245f
C1372 VN.n19 VSUBS 0.785346f
C1373 VN.n20 VSUBS 0.04966f
C1374 VN.n21 VSUBS 0.028633f
C1375 VN.n22 VSUBS 0.028633f
C1376 VN.n23 VSUBS 0.028633f
C1377 VN.n24 VSUBS 0.053632f
C1378 VN.n25 VSUBS 0.053632f
C1379 VN.n26 VSUBS 0.049794f
C1380 VN.n27 VSUBS 0.028633f
C1381 VN.n28 VSUBS 0.028633f
C1382 VN.n29 VSUBS 0.028633f
C1383 VN.n30 VSUBS 0.055041f
C1384 VN.n31 VSUBS 0.053632f
C1385 VN.n32 VSUBS 0.041716f
C1386 VN.n33 VSUBS 0.04622f
C1387 VN.n34 VSUBS 0.073436f
C1388 VN.t1 VSUBS 2.18245f
C1389 VN.n35 VSUBS 0.903325f
C1390 VN.n36 VSUBS 0.028633f
C1391 VN.n37 VSUBS 0.032759f
C1392 VN.n38 VSUBS 0.028633f
C1393 VN.n39 VSUBS 0.031124f
C1394 VN.n40 VSUBS 0.028633f
C1395 VN.t0 VSUBS 2.18245f
C1396 VN.n41 VSUBS 0.785346f
C1397 VN.n42 VSUBS 0.02317f
C1398 VN.n43 VSUBS 0.028633f
C1399 VN.t7 VSUBS 2.18245f
C1400 VN.n44 VSUBS 0.895348f
C1401 VN.t4 VSUBS 2.56421f
C1402 VN.n45 VSUBS 0.842466f
C1403 VN.n46 VSUBS 0.352625f
C1404 VN.n47 VSUBS 0.04966f
C1405 VN.n48 VSUBS 0.053632f
C1406 VN.n49 VSUBS 0.057212f
C1407 VN.n50 VSUBS 0.028633f
C1408 VN.n51 VSUBS 0.028633f
C1409 VN.n52 VSUBS 0.028633f
C1410 VN.n53 VSUBS 0.057212f
C1411 VN.n54 VSUBS 0.053632f
C1412 VN.n55 VSUBS 0.04966f
C1413 VN.n56 VSUBS 0.028633f
C1414 VN.n57 VSUBS 0.028633f
C1415 VN.n58 VSUBS 0.028633f
C1416 VN.n59 VSUBS 0.053632f
C1417 VN.n60 VSUBS 0.053632f
C1418 VN.n61 VSUBS 0.049794f
C1419 VN.n62 VSUBS 0.028633f
C1420 VN.n63 VSUBS 0.028633f
C1421 VN.n64 VSUBS 0.028633f
C1422 VN.n65 VSUBS 0.055041f
C1423 VN.n66 VSUBS 0.053632f
C1424 VN.n67 VSUBS 0.041716f
C1425 VN.n68 VSUBS 0.04622f
C1426 VN.n69 VSUBS 1.75698f
.ends

