* NGSPICE file created from diff_pair_sample_0106.ext - technology: sky130A

.subckt diff_pair_sample_0106 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X1 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X2 VTAIL.t19 VN.t1 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X3 VDD1.t8 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X4 VTAIL.t17 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X5 VDD2.t6 VN.t3 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=2.61
X6 VDD1.t7 VP.t2 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=2.61
X7 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=2.61
X8 VDD2.t5 VN.t4 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=2.61
X9 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=2.61
X10 VTAIL.t6 VP.t3 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X11 VTAIL.t14 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X12 VDD1.t5 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=2.61
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=2.61
X14 VDD2.t3 VN.t6 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=2.61
X15 VDD2.t2 VN.t7 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=2.61
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=0 ps=0 w=6.3 l=2.61
X17 VDD1.t4 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=2.457 ps=13.38 w=6.3 l=2.61
X18 VTAIL.t11 VN.t8 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X19 VTAIL.t2 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X20 VDD1.t2 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.457 pd=13.38 as=1.0395 ps=6.63 w=6.3 l=2.61
X21 VTAIL.t0 VP.t8 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X22 VTAIL.t8 VP.t9 VDD1.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
X23 VDD2.t0 VN.t9 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0395 pd=6.63 as=1.0395 ps=6.63 w=6.3 l=2.61
R0 VN.n81 VN.n42 161.3
R1 VN.n80 VN.n79 161.3
R2 VN.n78 VN.n43 161.3
R3 VN.n77 VN.n76 161.3
R4 VN.n75 VN.n44 161.3
R5 VN.n74 VN.n73 161.3
R6 VN.n72 VN.n71 161.3
R7 VN.n70 VN.n46 161.3
R8 VN.n69 VN.n68 161.3
R9 VN.n67 VN.n47 161.3
R10 VN.n66 VN.n65 161.3
R11 VN.n64 VN.n48 161.3
R12 VN.n62 VN.n61 161.3
R13 VN.n60 VN.n49 161.3
R14 VN.n59 VN.n58 161.3
R15 VN.n57 VN.n50 161.3
R16 VN.n56 VN.n55 161.3
R17 VN.n54 VN.n51 161.3
R18 VN.n39 VN.n0 161.3
R19 VN.n38 VN.n37 161.3
R20 VN.n36 VN.n1 161.3
R21 VN.n35 VN.n34 161.3
R22 VN.n33 VN.n2 161.3
R23 VN.n32 VN.n31 161.3
R24 VN.n30 VN.n29 161.3
R25 VN.n28 VN.n4 161.3
R26 VN.n27 VN.n26 161.3
R27 VN.n25 VN.n5 161.3
R28 VN.n24 VN.n23 161.3
R29 VN.n22 VN.n6 161.3
R30 VN.n20 VN.n19 161.3
R31 VN.n18 VN.n7 161.3
R32 VN.n17 VN.n16 161.3
R33 VN.n15 VN.n8 161.3
R34 VN.n14 VN.n13 161.3
R35 VN.n12 VN.n9 161.3
R36 VN.n41 VN.n40 104.514
R37 VN.n83 VN.n82 104.514
R38 VN.n11 VN.t3 90.7511
R39 VN.n53 VN.t6 90.7511
R40 VN.n11 VN.n10 63.1649
R41 VN.n53 VN.n52 63.1649
R42 VN.n10 VN.t5 58.1729
R43 VN.n21 VN.t0 58.1729
R44 VN.n3 VN.t2 58.1729
R45 VN.n40 VN.t4 58.1729
R46 VN.n52 VN.t8 58.1729
R47 VN.n63 VN.t9 58.1729
R48 VN.n45 VN.t1 58.1729
R49 VN.n82 VN.t7 58.1729
R50 VN.n16 VN.n15 56.5617
R51 VN.n27 VN.n5 56.5617
R52 VN.n58 VN.n57 56.5617
R53 VN.n69 VN.n47 56.5617
R54 VN.n34 VN.n1 56.0773
R55 VN.n76 VN.n43 56.0773
R56 VN VN.n83 49.0967
R57 VN.n34 VN.n33 25.0767
R58 VN.n76 VN.n75 25.0767
R59 VN.n14 VN.n9 24.5923
R60 VN.n15 VN.n14 24.5923
R61 VN.n16 VN.n7 24.5923
R62 VN.n20 VN.n7 24.5923
R63 VN.n23 VN.n22 24.5923
R64 VN.n23 VN.n5 24.5923
R65 VN.n28 VN.n27 24.5923
R66 VN.n29 VN.n28 24.5923
R67 VN.n33 VN.n32 24.5923
R68 VN.n38 VN.n1 24.5923
R69 VN.n39 VN.n38 24.5923
R70 VN.n57 VN.n56 24.5923
R71 VN.n56 VN.n51 24.5923
R72 VN.n65 VN.n47 24.5923
R73 VN.n65 VN.n64 24.5923
R74 VN.n62 VN.n49 24.5923
R75 VN.n58 VN.n49 24.5923
R76 VN.n75 VN.n74 24.5923
R77 VN.n71 VN.n70 24.5923
R78 VN.n70 VN.n69 24.5923
R79 VN.n81 VN.n80 24.5923
R80 VN.n80 VN.n43 24.5923
R81 VN.n32 VN.n3 15.2474
R82 VN.n74 VN.n45 15.2474
R83 VN.n21 VN.n20 12.2964
R84 VN.n22 VN.n21 12.2964
R85 VN.n64 VN.n63 12.2964
R86 VN.n63 VN.n62 12.2964
R87 VN.n10 VN.n9 9.3454
R88 VN.n29 VN.n3 9.3454
R89 VN.n52 VN.n51 9.3454
R90 VN.n71 VN.n45 9.3454
R91 VN.n54 VN.n53 7.05922
R92 VN.n12 VN.n11 7.05922
R93 VN.n40 VN.n39 6.39438
R94 VN.n82 VN.n81 6.39438
R95 VN.n83 VN.n42 0.278335
R96 VN.n41 VN.n0 0.278335
R97 VN.n79 VN.n42 0.189894
R98 VN.n79 VN.n78 0.189894
R99 VN.n78 VN.n77 0.189894
R100 VN.n77 VN.n44 0.189894
R101 VN.n73 VN.n44 0.189894
R102 VN.n73 VN.n72 0.189894
R103 VN.n72 VN.n46 0.189894
R104 VN.n68 VN.n46 0.189894
R105 VN.n68 VN.n67 0.189894
R106 VN.n67 VN.n66 0.189894
R107 VN.n66 VN.n48 0.189894
R108 VN.n61 VN.n48 0.189894
R109 VN.n61 VN.n60 0.189894
R110 VN.n60 VN.n59 0.189894
R111 VN.n59 VN.n50 0.189894
R112 VN.n55 VN.n50 0.189894
R113 VN.n55 VN.n54 0.189894
R114 VN.n13 VN.n12 0.189894
R115 VN.n13 VN.n8 0.189894
R116 VN.n17 VN.n8 0.189894
R117 VN.n18 VN.n17 0.189894
R118 VN.n19 VN.n18 0.189894
R119 VN.n19 VN.n6 0.189894
R120 VN.n24 VN.n6 0.189894
R121 VN.n25 VN.n24 0.189894
R122 VN.n26 VN.n25 0.189894
R123 VN.n26 VN.n4 0.189894
R124 VN.n30 VN.n4 0.189894
R125 VN.n31 VN.n30 0.189894
R126 VN.n31 VN.n2 0.189894
R127 VN.n35 VN.n2 0.189894
R128 VN.n36 VN.n35 0.189894
R129 VN.n37 VN.n36 0.189894
R130 VN.n37 VN.n0 0.189894
R131 VN VN.n41 0.153485
R132 VTAIL.n11 VTAIL.t13 51.8964
R133 VTAIL.n16 VTAIL.t1 51.8963
R134 VTAIL.n17 VTAIL.t10 51.8963
R135 VTAIL.n2 VTAIL.t3 51.8963
R136 VTAIL.n15 VTAIL.n14 48.7536
R137 VTAIL.n13 VTAIL.n12 48.7536
R138 VTAIL.n10 VTAIL.n9 48.7536
R139 VTAIL.n8 VTAIL.n7 48.7536
R140 VTAIL.n19 VTAIL.n18 48.7534
R141 VTAIL.n1 VTAIL.n0 48.7534
R142 VTAIL.n4 VTAIL.n3 48.7534
R143 VTAIL.n6 VTAIL.n5 48.7534
R144 VTAIL.n8 VTAIL.n6 22.8669
R145 VTAIL.n17 VTAIL.n16 20.3324
R146 VTAIL.n18 VTAIL.t12 3.14336
R147 VTAIL.n18 VTAIL.t17 3.14336
R148 VTAIL.n0 VTAIL.t18 3.14336
R149 VTAIL.n0 VTAIL.t14 3.14336
R150 VTAIL.n3 VTAIL.t4 3.14336
R151 VTAIL.n3 VTAIL.t2 3.14336
R152 VTAIL.n5 VTAIL.t9 3.14336
R153 VTAIL.n5 VTAIL.t6 3.14336
R154 VTAIL.n14 VTAIL.t7 3.14336
R155 VTAIL.n14 VTAIL.t0 3.14336
R156 VTAIL.n12 VTAIL.t5 3.14336
R157 VTAIL.n12 VTAIL.t8 3.14336
R158 VTAIL.n9 VTAIL.t16 3.14336
R159 VTAIL.n9 VTAIL.t11 3.14336
R160 VTAIL.n7 VTAIL.t15 3.14336
R161 VTAIL.n7 VTAIL.t19 3.14336
R162 VTAIL.n10 VTAIL.n8 2.53498
R163 VTAIL.n11 VTAIL.n10 2.53498
R164 VTAIL.n15 VTAIL.n13 2.53498
R165 VTAIL.n16 VTAIL.n15 2.53498
R166 VTAIL.n6 VTAIL.n4 2.53498
R167 VTAIL.n4 VTAIL.n2 2.53498
R168 VTAIL.n19 VTAIL.n17 2.53498
R169 VTAIL VTAIL.n1 1.95955
R170 VTAIL.n13 VTAIL.n11 1.73757
R171 VTAIL.n2 VTAIL.n1 1.73757
R172 VTAIL VTAIL.n19 0.575931
R173 VDD2.n1 VDD2.t6 71.1096
R174 VDD2.n4 VDD2.t2 68.5752
R175 VDD2.n3 VDD2.n2 67.2777
R176 VDD2 VDD2.n7 67.2749
R177 VDD2.n6 VDD2.n5 65.4324
R178 VDD2.n1 VDD2.n0 65.4322
R179 VDD2.n4 VDD2.n3 41.1851
R180 VDD2.n7 VDD2.t1 3.14336
R181 VDD2.n7 VDD2.t3 3.14336
R182 VDD2.n5 VDD2.t8 3.14336
R183 VDD2.n5 VDD2.t0 3.14336
R184 VDD2.n2 VDD2.t7 3.14336
R185 VDD2.n2 VDD2.t5 3.14336
R186 VDD2.n0 VDD2.t4 3.14336
R187 VDD2.n0 VDD2.t9 3.14336
R188 VDD2.n6 VDD2.n4 2.53498
R189 VDD2 VDD2.n6 0.69231
R190 VDD2.n3 VDD2.n1 0.578775
R191 B.n788 B.n787 585
R192 B.n789 B.n788 585
R193 B.n259 B.n140 585
R194 B.n258 B.n257 585
R195 B.n256 B.n255 585
R196 B.n254 B.n253 585
R197 B.n252 B.n251 585
R198 B.n250 B.n249 585
R199 B.n248 B.n247 585
R200 B.n246 B.n245 585
R201 B.n244 B.n243 585
R202 B.n242 B.n241 585
R203 B.n240 B.n239 585
R204 B.n238 B.n237 585
R205 B.n236 B.n235 585
R206 B.n234 B.n233 585
R207 B.n232 B.n231 585
R208 B.n230 B.n229 585
R209 B.n228 B.n227 585
R210 B.n226 B.n225 585
R211 B.n224 B.n223 585
R212 B.n222 B.n221 585
R213 B.n220 B.n219 585
R214 B.n218 B.n217 585
R215 B.n216 B.n215 585
R216 B.n214 B.n213 585
R217 B.n212 B.n211 585
R218 B.n210 B.n209 585
R219 B.n208 B.n207 585
R220 B.n206 B.n205 585
R221 B.n204 B.n203 585
R222 B.n202 B.n201 585
R223 B.n200 B.n199 585
R224 B.n198 B.n197 585
R225 B.n196 B.n195 585
R226 B.n193 B.n192 585
R227 B.n191 B.n190 585
R228 B.n189 B.n188 585
R229 B.n187 B.n186 585
R230 B.n185 B.n184 585
R231 B.n183 B.n182 585
R232 B.n181 B.n180 585
R233 B.n179 B.n178 585
R234 B.n177 B.n176 585
R235 B.n175 B.n174 585
R236 B.n173 B.n172 585
R237 B.n171 B.n170 585
R238 B.n169 B.n168 585
R239 B.n167 B.n166 585
R240 B.n165 B.n164 585
R241 B.n163 B.n162 585
R242 B.n161 B.n160 585
R243 B.n159 B.n158 585
R244 B.n157 B.n156 585
R245 B.n155 B.n154 585
R246 B.n153 B.n152 585
R247 B.n151 B.n150 585
R248 B.n149 B.n148 585
R249 B.n147 B.n146 585
R250 B.n109 B.n108 585
R251 B.n786 B.n110 585
R252 B.n790 B.n110 585
R253 B.n785 B.n784 585
R254 B.n784 B.n106 585
R255 B.n783 B.n105 585
R256 B.n796 B.n105 585
R257 B.n782 B.n104 585
R258 B.n797 B.n104 585
R259 B.n781 B.n103 585
R260 B.n798 B.n103 585
R261 B.n780 B.n779 585
R262 B.n779 B.n99 585
R263 B.n778 B.n98 585
R264 B.n804 B.n98 585
R265 B.n777 B.n97 585
R266 B.n805 B.n97 585
R267 B.n776 B.n96 585
R268 B.n806 B.n96 585
R269 B.n775 B.n774 585
R270 B.n774 B.n92 585
R271 B.n773 B.n91 585
R272 B.n812 B.n91 585
R273 B.n772 B.n90 585
R274 B.n813 B.n90 585
R275 B.n771 B.n89 585
R276 B.n814 B.n89 585
R277 B.n770 B.n769 585
R278 B.n769 B.n85 585
R279 B.n768 B.n84 585
R280 B.n820 B.n84 585
R281 B.n767 B.n83 585
R282 B.n821 B.n83 585
R283 B.n766 B.n82 585
R284 B.n822 B.n82 585
R285 B.n765 B.n764 585
R286 B.n764 B.n78 585
R287 B.n763 B.n77 585
R288 B.n828 B.n77 585
R289 B.n762 B.n76 585
R290 B.n829 B.n76 585
R291 B.n761 B.n75 585
R292 B.n830 B.n75 585
R293 B.n760 B.n759 585
R294 B.n759 B.n71 585
R295 B.n758 B.n70 585
R296 B.n836 B.n70 585
R297 B.n757 B.n69 585
R298 B.n837 B.n69 585
R299 B.n756 B.n68 585
R300 B.n838 B.n68 585
R301 B.n755 B.n754 585
R302 B.n754 B.n64 585
R303 B.n753 B.n63 585
R304 B.n844 B.n63 585
R305 B.n752 B.n62 585
R306 B.n845 B.n62 585
R307 B.n751 B.n61 585
R308 B.n846 B.n61 585
R309 B.n750 B.n749 585
R310 B.n749 B.n57 585
R311 B.n748 B.n56 585
R312 B.n852 B.n56 585
R313 B.n747 B.n55 585
R314 B.n853 B.n55 585
R315 B.n746 B.n54 585
R316 B.n854 B.n54 585
R317 B.n745 B.n744 585
R318 B.n744 B.n50 585
R319 B.n743 B.n49 585
R320 B.n860 B.n49 585
R321 B.n742 B.n48 585
R322 B.n861 B.n48 585
R323 B.n741 B.n47 585
R324 B.n862 B.n47 585
R325 B.n740 B.n739 585
R326 B.n739 B.n43 585
R327 B.n738 B.n42 585
R328 B.n868 B.n42 585
R329 B.n737 B.n41 585
R330 B.n869 B.n41 585
R331 B.n736 B.n40 585
R332 B.n870 B.n40 585
R333 B.n735 B.n734 585
R334 B.n734 B.n36 585
R335 B.n733 B.n35 585
R336 B.n876 B.n35 585
R337 B.n732 B.n34 585
R338 B.n877 B.n34 585
R339 B.n731 B.n33 585
R340 B.n878 B.n33 585
R341 B.n730 B.n729 585
R342 B.n729 B.n32 585
R343 B.n728 B.n28 585
R344 B.n884 B.n28 585
R345 B.n727 B.n27 585
R346 B.n885 B.n27 585
R347 B.n726 B.n26 585
R348 B.n886 B.n26 585
R349 B.n725 B.n724 585
R350 B.n724 B.n22 585
R351 B.n723 B.n21 585
R352 B.n892 B.n21 585
R353 B.n722 B.n20 585
R354 B.n893 B.n20 585
R355 B.n721 B.n19 585
R356 B.n894 B.n19 585
R357 B.n720 B.n719 585
R358 B.n719 B.n15 585
R359 B.n718 B.n14 585
R360 B.n900 B.n14 585
R361 B.n717 B.n13 585
R362 B.n901 B.n13 585
R363 B.n716 B.n12 585
R364 B.n902 B.n12 585
R365 B.n715 B.n714 585
R366 B.n714 B.n8 585
R367 B.n713 B.n7 585
R368 B.n908 B.n7 585
R369 B.n712 B.n6 585
R370 B.n909 B.n6 585
R371 B.n711 B.n5 585
R372 B.n910 B.n5 585
R373 B.n710 B.n709 585
R374 B.n709 B.n4 585
R375 B.n708 B.n260 585
R376 B.n708 B.n707 585
R377 B.n698 B.n261 585
R378 B.n262 B.n261 585
R379 B.n700 B.n699 585
R380 B.n701 B.n700 585
R381 B.n697 B.n267 585
R382 B.n267 B.n266 585
R383 B.n696 B.n695 585
R384 B.n695 B.n694 585
R385 B.n269 B.n268 585
R386 B.n270 B.n269 585
R387 B.n687 B.n686 585
R388 B.n688 B.n687 585
R389 B.n685 B.n275 585
R390 B.n275 B.n274 585
R391 B.n684 B.n683 585
R392 B.n683 B.n682 585
R393 B.n277 B.n276 585
R394 B.n278 B.n277 585
R395 B.n675 B.n674 585
R396 B.n676 B.n675 585
R397 B.n673 B.n283 585
R398 B.n283 B.n282 585
R399 B.n672 B.n671 585
R400 B.n671 B.n670 585
R401 B.n285 B.n284 585
R402 B.n663 B.n285 585
R403 B.n662 B.n661 585
R404 B.n664 B.n662 585
R405 B.n660 B.n290 585
R406 B.n290 B.n289 585
R407 B.n659 B.n658 585
R408 B.n658 B.n657 585
R409 B.n292 B.n291 585
R410 B.n293 B.n292 585
R411 B.n650 B.n649 585
R412 B.n651 B.n650 585
R413 B.n648 B.n298 585
R414 B.n298 B.n297 585
R415 B.n647 B.n646 585
R416 B.n646 B.n645 585
R417 B.n300 B.n299 585
R418 B.n301 B.n300 585
R419 B.n638 B.n637 585
R420 B.n639 B.n638 585
R421 B.n636 B.n306 585
R422 B.n306 B.n305 585
R423 B.n635 B.n634 585
R424 B.n634 B.n633 585
R425 B.n308 B.n307 585
R426 B.n309 B.n308 585
R427 B.n626 B.n625 585
R428 B.n627 B.n626 585
R429 B.n624 B.n314 585
R430 B.n314 B.n313 585
R431 B.n623 B.n622 585
R432 B.n622 B.n621 585
R433 B.n316 B.n315 585
R434 B.n317 B.n316 585
R435 B.n614 B.n613 585
R436 B.n615 B.n614 585
R437 B.n612 B.n322 585
R438 B.n322 B.n321 585
R439 B.n611 B.n610 585
R440 B.n610 B.n609 585
R441 B.n324 B.n323 585
R442 B.n325 B.n324 585
R443 B.n602 B.n601 585
R444 B.n603 B.n602 585
R445 B.n600 B.n330 585
R446 B.n330 B.n329 585
R447 B.n599 B.n598 585
R448 B.n598 B.n597 585
R449 B.n332 B.n331 585
R450 B.n333 B.n332 585
R451 B.n590 B.n589 585
R452 B.n591 B.n590 585
R453 B.n588 B.n337 585
R454 B.n341 B.n337 585
R455 B.n587 B.n586 585
R456 B.n586 B.n585 585
R457 B.n339 B.n338 585
R458 B.n340 B.n339 585
R459 B.n578 B.n577 585
R460 B.n579 B.n578 585
R461 B.n576 B.n346 585
R462 B.n346 B.n345 585
R463 B.n575 B.n574 585
R464 B.n574 B.n573 585
R465 B.n348 B.n347 585
R466 B.n349 B.n348 585
R467 B.n566 B.n565 585
R468 B.n567 B.n566 585
R469 B.n564 B.n354 585
R470 B.n354 B.n353 585
R471 B.n563 B.n562 585
R472 B.n562 B.n561 585
R473 B.n356 B.n355 585
R474 B.n357 B.n356 585
R475 B.n554 B.n553 585
R476 B.n555 B.n554 585
R477 B.n552 B.n361 585
R478 B.n365 B.n361 585
R479 B.n551 B.n550 585
R480 B.n550 B.n549 585
R481 B.n363 B.n362 585
R482 B.n364 B.n363 585
R483 B.n542 B.n541 585
R484 B.n543 B.n542 585
R485 B.n540 B.n370 585
R486 B.n370 B.n369 585
R487 B.n539 B.n538 585
R488 B.n538 B.n537 585
R489 B.n372 B.n371 585
R490 B.n373 B.n372 585
R491 B.n530 B.n529 585
R492 B.n531 B.n530 585
R493 B.n376 B.n375 585
R494 B.n414 B.n413 585
R495 B.n415 B.n411 585
R496 B.n411 B.n377 585
R497 B.n417 B.n416 585
R498 B.n419 B.n410 585
R499 B.n422 B.n421 585
R500 B.n423 B.n409 585
R501 B.n425 B.n424 585
R502 B.n427 B.n408 585
R503 B.n430 B.n429 585
R504 B.n431 B.n407 585
R505 B.n433 B.n432 585
R506 B.n435 B.n406 585
R507 B.n438 B.n437 585
R508 B.n439 B.n405 585
R509 B.n441 B.n440 585
R510 B.n443 B.n404 585
R511 B.n446 B.n445 585
R512 B.n447 B.n403 585
R513 B.n449 B.n448 585
R514 B.n451 B.n402 585
R515 B.n454 B.n453 585
R516 B.n455 B.n401 585
R517 B.n457 B.n456 585
R518 B.n459 B.n400 585
R519 B.n462 B.n461 585
R520 B.n463 B.n396 585
R521 B.n465 B.n464 585
R522 B.n467 B.n395 585
R523 B.n470 B.n469 585
R524 B.n471 B.n394 585
R525 B.n473 B.n472 585
R526 B.n475 B.n393 585
R527 B.n478 B.n477 585
R528 B.n480 B.n390 585
R529 B.n482 B.n481 585
R530 B.n484 B.n389 585
R531 B.n487 B.n486 585
R532 B.n488 B.n388 585
R533 B.n490 B.n489 585
R534 B.n492 B.n387 585
R535 B.n495 B.n494 585
R536 B.n496 B.n386 585
R537 B.n498 B.n497 585
R538 B.n500 B.n385 585
R539 B.n503 B.n502 585
R540 B.n504 B.n384 585
R541 B.n506 B.n505 585
R542 B.n508 B.n383 585
R543 B.n511 B.n510 585
R544 B.n512 B.n382 585
R545 B.n514 B.n513 585
R546 B.n516 B.n381 585
R547 B.n519 B.n518 585
R548 B.n520 B.n380 585
R549 B.n522 B.n521 585
R550 B.n524 B.n379 585
R551 B.n527 B.n526 585
R552 B.n528 B.n378 585
R553 B.n533 B.n532 585
R554 B.n532 B.n531 585
R555 B.n534 B.n374 585
R556 B.n374 B.n373 585
R557 B.n536 B.n535 585
R558 B.n537 B.n536 585
R559 B.n368 B.n367 585
R560 B.n369 B.n368 585
R561 B.n545 B.n544 585
R562 B.n544 B.n543 585
R563 B.n546 B.n366 585
R564 B.n366 B.n364 585
R565 B.n548 B.n547 585
R566 B.n549 B.n548 585
R567 B.n360 B.n359 585
R568 B.n365 B.n360 585
R569 B.n557 B.n556 585
R570 B.n556 B.n555 585
R571 B.n558 B.n358 585
R572 B.n358 B.n357 585
R573 B.n560 B.n559 585
R574 B.n561 B.n560 585
R575 B.n352 B.n351 585
R576 B.n353 B.n352 585
R577 B.n569 B.n568 585
R578 B.n568 B.n567 585
R579 B.n570 B.n350 585
R580 B.n350 B.n349 585
R581 B.n572 B.n571 585
R582 B.n573 B.n572 585
R583 B.n344 B.n343 585
R584 B.n345 B.n344 585
R585 B.n581 B.n580 585
R586 B.n580 B.n579 585
R587 B.n582 B.n342 585
R588 B.n342 B.n340 585
R589 B.n584 B.n583 585
R590 B.n585 B.n584 585
R591 B.n336 B.n335 585
R592 B.n341 B.n336 585
R593 B.n593 B.n592 585
R594 B.n592 B.n591 585
R595 B.n594 B.n334 585
R596 B.n334 B.n333 585
R597 B.n596 B.n595 585
R598 B.n597 B.n596 585
R599 B.n328 B.n327 585
R600 B.n329 B.n328 585
R601 B.n605 B.n604 585
R602 B.n604 B.n603 585
R603 B.n606 B.n326 585
R604 B.n326 B.n325 585
R605 B.n608 B.n607 585
R606 B.n609 B.n608 585
R607 B.n320 B.n319 585
R608 B.n321 B.n320 585
R609 B.n617 B.n616 585
R610 B.n616 B.n615 585
R611 B.n618 B.n318 585
R612 B.n318 B.n317 585
R613 B.n620 B.n619 585
R614 B.n621 B.n620 585
R615 B.n312 B.n311 585
R616 B.n313 B.n312 585
R617 B.n629 B.n628 585
R618 B.n628 B.n627 585
R619 B.n630 B.n310 585
R620 B.n310 B.n309 585
R621 B.n632 B.n631 585
R622 B.n633 B.n632 585
R623 B.n304 B.n303 585
R624 B.n305 B.n304 585
R625 B.n641 B.n640 585
R626 B.n640 B.n639 585
R627 B.n642 B.n302 585
R628 B.n302 B.n301 585
R629 B.n644 B.n643 585
R630 B.n645 B.n644 585
R631 B.n296 B.n295 585
R632 B.n297 B.n296 585
R633 B.n653 B.n652 585
R634 B.n652 B.n651 585
R635 B.n654 B.n294 585
R636 B.n294 B.n293 585
R637 B.n656 B.n655 585
R638 B.n657 B.n656 585
R639 B.n288 B.n287 585
R640 B.n289 B.n288 585
R641 B.n666 B.n665 585
R642 B.n665 B.n664 585
R643 B.n667 B.n286 585
R644 B.n663 B.n286 585
R645 B.n669 B.n668 585
R646 B.n670 B.n669 585
R647 B.n281 B.n280 585
R648 B.n282 B.n281 585
R649 B.n678 B.n677 585
R650 B.n677 B.n676 585
R651 B.n679 B.n279 585
R652 B.n279 B.n278 585
R653 B.n681 B.n680 585
R654 B.n682 B.n681 585
R655 B.n273 B.n272 585
R656 B.n274 B.n273 585
R657 B.n690 B.n689 585
R658 B.n689 B.n688 585
R659 B.n691 B.n271 585
R660 B.n271 B.n270 585
R661 B.n693 B.n692 585
R662 B.n694 B.n693 585
R663 B.n265 B.n264 585
R664 B.n266 B.n265 585
R665 B.n703 B.n702 585
R666 B.n702 B.n701 585
R667 B.n704 B.n263 585
R668 B.n263 B.n262 585
R669 B.n706 B.n705 585
R670 B.n707 B.n706 585
R671 B.n2 B.n0 585
R672 B.n4 B.n2 585
R673 B.n3 B.n1 585
R674 B.n909 B.n3 585
R675 B.n907 B.n906 585
R676 B.n908 B.n907 585
R677 B.n905 B.n9 585
R678 B.n9 B.n8 585
R679 B.n904 B.n903 585
R680 B.n903 B.n902 585
R681 B.n11 B.n10 585
R682 B.n901 B.n11 585
R683 B.n899 B.n898 585
R684 B.n900 B.n899 585
R685 B.n897 B.n16 585
R686 B.n16 B.n15 585
R687 B.n896 B.n895 585
R688 B.n895 B.n894 585
R689 B.n18 B.n17 585
R690 B.n893 B.n18 585
R691 B.n891 B.n890 585
R692 B.n892 B.n891 585
R693 B.n889 B.n23 585
R694 B.n23 B.n22 585
R695 B.n888 B.n887 585
R696 B.n887 B.n886 585
R697 B.n25 B.n24 585
R698 B.n885 B.n25 585
R699 B.n883 B.n882 585
R700 B.n884 B.n883 585
R701 B.n881 B.n29 585
R702 B.n32 B.n29 585
R703 B.n880 B.n879 585
R704 B.n879 B.n878 585
R705 B.n31 B.n30 585
R706 B.n877 B.n31 585
R707 B.n875 B.n874 585
R708 B.n876 B.n875 585
R709 B.n873 B.n37 585
R710 B.n37 B.n36 585
R711 B.n872 B.n871 585
R712 B.n871 B.n870 585
R713 B.n39 B.n38 585
R714 B.n869 B.n39 585
R715 B.n867 B.n866 585
R716 B.n868 B.n867 585
R717 B.n865 B.n44 585
R718 B.n44 B.n43 585
R719 B.n864 B.n863 585
R720 B.n863 B.n862 585
R721 B.n46 B.n45 585
R722 B.n861 B.n46 585
R723 B.n859 B.n858 585
R724 B.n860 B.n859 585
R725 B.n857 B.n51 585
R726 B.n51 B.n50 585
R727 B.n856 B.n855 585
R728 B.n855 B.n854 585
R729 B.n53 B.n52 585
R730 B.n853 B.n53 585
R731 B.n851 B.n850 585
R732 B.n852 B.n851 585
R733 B.n849 B.n58 585
R734 B.n58 B.n57 585
R735 B.n848 B.n847 585
R736 B.n847 B.n846 585
R737 B.n60 B.n59 585
R738 B.n845 B.n60 585
R739 B.n843 B.n842 585
R740 B.n844 B.n843 585
R741 B.n841 B.n65 585
R742 B.n65 B.n64 585
R743 B.n840 B.n839 585
R744 B.n839 B.n838 585
R745 B.n67 B.n66 585
R746 B.n837 B.n67 585
R747 B.n835 B.n834 585
R748 B.n836 B.n835 585
R749 B.n833 B.n72 585
R750 B.n72 B.n71 585
R751 B.n832 B.n831 585
R752 B.n831 B.n830 585
R753 B.n74 B.n73 585
R754 B.n829 B.n74 585
R755 B.n827 B.n826 585
R756 B.n828 B.n827 585
R757 B.n825 B.n79 585
R758 B.n79 B.n78 585
R759 B.n824 B.n823 585
R760 B.n823 B.n822 585
R761 B.n81 B.n80 585
R762 B.n821 B.n81 585
R763 B.n819 B.n818 585
R764 B.n820 B.n819 585
R765 B.n817 B.n86 585
R766 B.n86 B.n85 585
R767 B.n816 B.n815 585
R768 B.n815 B.n814 585
R769 B.n88 B.n87 585
R770 B.n813 B.n88 585
R771 B.n811 B.n810 585
R772 B.n812 B.n811 585
R773 B.n809 B.n93 585
R774 B.n93 B.n92 585
R775 B.n808 B.n807 585
R776 B.n807 B.n806 585
R777 B.n95 B.n94 585
R778 B.n805 B.n95 585
R779 B.n803 B.n802 585
R780 B.n804 B.n803 585
R781 B.n801 B.n100 585
R782 B.n100 B.n99 585
R783 B.n800 B.n799 585
R784 B.n799 B.n798 585
R785 B.n102 B.n101 585
R786 B.n797 B.n102 585
R787 B.n795 B.n794 585
R788 B.n796 B.n795 585
R789 B.n793 B.n107 585
R790 B.n107 B.n106 585
R791 B.n792 B.n791 585
R792 B.n791 B.n790 585
R793 B.n912 B.n911 585
R794 B.n911 B.n910 585
R795 B.n532 B.n376 521.33
R796 B.n791 B.n109 521.33
R797 B.n530 B.n378 521.33
R798 B.n788 B.n110 521.33
R799 B.n391 B.t10 266.235
R800 B.n397 B.t21 266.235
R801 B.n144 B.t18 266.235
R802 B.n141 B.t14 266.235
R803 B.n789 B.n139 256.663
R804 B.n789 B.n138 256.663
R805 B.n789 B.n137 256.663
R806 B.n789 B.n136 256.663
R807 B.n789 B.n135 256.663
R808 B.n789 B.n134 256.663
R809 B.n789 B.n133 256.663
R810 B.n789 B.n132 256.663
R811 B.n789 B.n131 256.663
R812 B.n789 B.n130 256.663
R813 B.n789 B.n129 256.663
R814 B.n789 B.n128 256.663
R815 B.n789 B.n127 256.663
R816 B.n789 B.n126 256.663
R817 B.n789 B.n125 256.663
R818 B.n789 B.n124 256.663
R819 B.n789 B.n123 256.663
R820 B.n789 B.n122 256.663
R821 B.n789 B.n121 256.663
R822 B.n789 B.n120 256.663
R823 B.n789 B.n119 256.663
R824 B.n789 B.n118 256.663
R825 B.n789 B.n117 256.663
R826 B.n789 B.n116 256.663
R827 B.n789 B.n115 256.663
R828 B.n789 B.n114 256.663
R829 B.n789 B.n113 256.663
R830 B.n789 B.n112 256.663
R831 B.n789 B.n111 256.663
R832 B.n412 B.n377 256.663
R833 B.n418 B.n377 256.663
R834 B.n420 B.n377 256.663
R835 B.n426 B.n377 256.663
R836 B.n428 B.n377 256.663
R837 B.n434 B.n377 256.663
R838 B.n436 B.n377 256.663
R839 B.n442 B.n377 256.663
R840 B.n444 B.n377 256.663
R841 B.n450 B.n377 256.663
R842 B.n452 B.n377 256.663
R843 B.n458 B.n377 256.663
R844 B.n460 B.n377 256.663
R845 B.n466 B.n377 256.663
R846 B.n468 B.n377 256.663
R847 B.n474 B.n377 256.663
R848 B.n476 B.n377 256.663
R849 B.n483 B.n377 256.663
R850 B.n485 B.n377 256.663
R851 B.n491 B.n377 256.663
R852 B.n493 B.n377 256.663
R853 B.n499 B.n377 256.663
R854 B.n501 B.n377 256.663
R855 B.n507 B.n377 256.663
R856 B.n509 B.n377 256.663
R857 B.n515 B.n377 256.663
R858 B.n517 B.n377 256.663
R859 B.n523 B.n377 256.663
R860 B.n525 B.n377 256.663
R861 B.n532 B.n374 163.367
R862 B.n536 B.n374 163.367
R863 B.n536 B.n368 163.367
R864 B.n544 B.n368 163.367
R865 B.n544 B.n366 163.367
R866 B.n548 B.n366 163.367
R867 B.n548 B.n360 163.367
R868 B.n556 B.n360 163.367
R869 B.n556 B.n358 163.367
R870 B.n560 B.n358 163.367
R871 B.n560 B.n352 163.367
R872 B.n568 B.n352 163.367
R873 B.n568 B.n350 163.367
R874 B.n572 B.n350 163.367
R875 B.n572 B.n344 163.367
R876 B.n580 B.n344 163.367
R877 B.n580 B.n342 163.367
R878 B.n584 B.n342 163.367
R879 B.n584 B.n336 163.367
R880 B.n592 B.n336 163.367
R881 B.n592 B.n334 163.367
R882 B.n596 B.n334 163.367
R883 B.n596 B.n328 163.367
R884 B.n604 B.n328 163.367
R885 B.n604 B.n326 163.367
R886 B.n608 B.n326 163.367
R887 B.n608 B.n320 163.367
R888 B.n616 B.n320 163.367
R889 B.n616 B.n318 163.367
R890 B.n620 B.n318 163.367
R891 B.n620 B.n312 163.367
R892 B.n628 B.n312 163.367
R893 B.n628 B.n310 163.367
R894 B.n632 B.n310 163.367
R895 B.n632 B.n304 163.367
R896 B.n640 B.n304 163.367
R897 B.n640 B.n302 163.367
R898 B.n644 B.n302 163.367
R899 B.n644 B.n296 163.367
R900 B.n652 B.n296 163.367
R901 B.n652 B.n294 163.367
R902 B.n656 B.n294 163.367
R903 B.n656 B.n288 163.367
R904 B.n665 B.n288 163.367
R905 B.n665 B.n286 163.367
R906 B.n669 B.n286 163.367
R907 B.n669 B.n281 163.367
R908 B.n677 B.n281 163.367
R909 B.n677 B.n279 163.367
R910 B.n681 B.n279 163.367
R911 B.n681 B.n273 163.367
R912 B.n689 B.n273 163.367
R913 B.n689 B.n271 163.367
R914 B.n693 B.n271 163.367
R915 B.n693 B.n265 163.367
R916 B.n702 B.n265 163.367
R917 B.n702 B.n263 163.367
R918 B.n706 B.n263 163.367
R919 B.n706 B.n2 163.367
R920 B.n911 B.n2 163.367
R921 B.n911 B.n3 163.367
R922 B.n907 B.n3 163.367
R923 B.n907 B.n9 163.367
R924 B.n903 B.n9 163.367
R925 B.n903 B.n11 163.367
R926 B.n899 B.n11 163.367
R927 B.n899 B.n16 163.367
R928 B.n895 B.n16 163.367
R929 B.n895 B.n18 163.367
R930 B.n891 B.n18 163.367
R931 B.n891 B.n23 163.367
R932 B.n887 B.n23 163.367
R933 B.n887 B.n25 163.367
R934 B.n883 B.n25 163.367
R935 B.n883 B.n29 163.367
R936 B.n879 B.n29 163.367
R937 B.n879 B.n31 163.367
R938 B.n875 B.n31 163.367
R939 B.n875 B.n37 163.367
R940 B.n871 B.n37 163.367
R941 B.n871 B.n39 163.367
R942 B.n867 B.n39 163.367
R943 B.n867 B.n44 163.367
R944 B.n863 B.n44 163.367
R945 B.n863 B.n46 163.367
R946 B.n859 B.n46 163.367
R947 B.n859 B.n51 163.367
R948 B.n855 B.n51 163.367
R949 B.n855 B.n53 163.367
R950 B.n851 B.n53 163.367
R951 B.n851 B.n58 163.367
R952 B.n847 B.n58 163.367
R953 B.n847 B.n60 163.367
R954 B.n843 B.n60 163.367
R955 B.n843 B.n65 163.367
R956 B.n839 B.n65 163.367
R957 B.n839 B.n67 163.367
R958 B.n835 B.n67 163.367
R959 B.n835 B.n72 163.367
R960 B.n831 B.n72 163.367
R961 B.n831 B.n74 163.367
R962 B.n827 B.n74 163.367
R963 B.n827 B.n79 163.367
R964 B.n823 B.n79 163.367
R965 B.n823 B.n81 163.367
R966 B.n819 B.n81 163.367
R967 B.n819 B.n86 163.367
R968 B.n815 B.n86 163.367
R969 B.n815 B.n88 163.367
R970 B.n811 B.n88 163.367
R971 B.n811 B.n93 163.367
R972 B.n807 B.n93 163.367
R973 B.n807 B.n95 163.367
R974 B.n803 B.n95 163.367
R975 B.n803 B.n100 163.367
R976 B.n799 B.n100 163.367
R977 B.n799 B.n102 163.367
R978 B.n795 B.n102 163.367
R979 B.n795 B.n107 163.367
R980 B.n791 B.n107 163.367
R981 B.n413 B.n411 163.367
R982 B.n417 B.n411 163.367
R983 B.n421 B.n419 163.367
R984 B.n425 B.n409 163.367
R985 B.n429 B.n427 163.367
R986 B.n433 B.n407 163.367
R987 B.n437 B.n435 163.367
R988 B.n441 B.n405 163.367
R989 B.n445 B.n443 163.367
R990 B.n449 B.n403 163.367
R991 B.n453 B.n451 163.367
R992 B.n457 B.n401 163.367
R993 B.n461 B.n459 163.367
R994 B.n465 B.n396 163.367
R995 B.n469 B.n467 163.367
R996 B.n473 B.n394 163.367
R997 B.n477 B.n475 163.367
R998 B.n482 B.n390 163.367
R999 B.n486 B.n484 163.367
R1000 B.n490 B.n388 163.367
R1001 B.n494 B.n492 163.367
R1002 B.n498 B.n386 163.367
R1003 B.n502 B.n500 163.367
R1004 B.n506 B.n384 163.367
R1005 B.n510 B.n508 163.367
R1006 B.n514 B.n382 163.367
R1007 B.n518 B.n516 163.367
R1008 B.n522 B.n380 163.367
R1009 B.n526 B.n524 163.367
R1010 B.n530 B.n372 163.367
R1011 B.n538 B.n372 163.367
R1012 B.n538 B.n370 163.367
R1013 B.n542 B.n370 163.367
R1014 B.n542 B.n363 163.367
R1015 B.n550 B.n363 163.367
R1016 B.n550 B.n361 163.367
R1017 B.n554 B.n361 163.367
R1018 B.n554 B.n356 163.367
R1019 B.n562 B.n356 163.367
R1020 B.n562 B.n354 163.367
R1021 B.n566 B.n354 163.367
R1022 B.n566 B.n348 163.367
R1023 B.n574 B.n348 163.367
R1024 B.n574 B.n346 163.367
R1025 B.n578 B.n346 163.367
R1026 B.n578 B.n339 163.367
R1027 B.n586 B.n339 163.367
R1028 B.n586 B.n337 163.367
R1029 B.n590 B.n337 163.367
R1030 B.n590 B.n332 163.367
R1031 B.n598 B.n332 163.367
R1032 B.n598 B.n330 163.367
R1033 B.n602 B.n330 163.367
R1034 B.n602 B.n324 163.367
R1035 B.n610 B.n324 163.367
R1036 B.n610 B.n322 163.367
R1037 B.n614 B.n322 163.367
R1038 B.n614 B.n316 163.367
R1039 B.n622 B.n316 163.367
R1040 B.n622 B.n314 163.367
R1041 B.n626 B.n314 163.367
R1042 B.n626 B.n308 163.367
R1043 B.n634 B.n308 163.367
R1044 B.n634 B.n306 163.367
R1045 B.n638 B.n306 163.367
R1046 B.n638 B.n300 163.367
R1047 B.n646 B.n300 163.367
R1048 B.n646 B.n298 163.367
R1049 B.n650 B.n298 163.367
R1050 B.n650 B.n292 163.367
R1051 B.n658 B.n292 163.367
R1052 B.n658 B.n290 163.367
R1053 B.n662 B.n290 163.367
R1054 B.n662 B.n285 163.367
R1055 B.n671 B.n285 163.367
R1056 B.n671 B.n283 163.367
R1057 B.n675 B.n283 163.367
R1058 B.n675 B.n277 163.367
R1059 B.n683 B.n277 163.367
R1060 B.n683 B.n275 163.367
R1061 B.n687 B.n275 163.367
R1062 B.n687 B.n269 163.367
R1063 B.n695 B.n269 163.367
R1064 B.n695 B.n267 163.367
R1065 B.n700 B.n267 163.367
R1066 B.n700 B.n261 163.367
R1067 B.n708 B.n261 163.367
R1068 B.n709 B.n708 163.367
R1069 B.n709 B.n5 163.367
R1070 B.n6 B.n5 163.367
R1071 B.n7 B.n6 163.367
R1072 B.n714 B.n7 163.367
R1073 B.n714 B.n12 163.367
R1074 B.n13 B.n12 163.367
R1075 B.n14 B.n13 163.367
R1076 B.n719 B.n14 163.367
R1077 B.n719 B.n19 163.367
R1078 B.n20 B.n19 163.367
R1079 B.n21 B.n20 163.367
R1080 B.n724 B.n21 163.367
R1081 B.n724 B.n26 163.367
R1082 B.n27 B.n26 163.367
R1083 B.n28 B.n27 163.367
R1084 B.n729 B.n28 163.367
R1085 B.n729 B.n33 163.367
R1086 B.n34 B.n33 163.367
R1087 B.n35 B.n34 163.367
R1088 B.n734 B.n35 163.367
R1089 B.n734 B.n40 163.367
R1090 B.n41 B.n40 163.367
R1091 B.n42 B.n41 163.367
R1092 B.n739 B.n42 163.367
R1093 B.n739 B.n47 163.367
R1094 B.n48 B.n47 163.367
R1095 B.n49 B.n48 163.367
R1096 B.n744 B.n49 163.367
R1097 B.n744 B.n54 163.367
R1098 B.n55 B.n54 163.367
R1099 B.n56 B.n55 163.367
R1100 B.n749 B.n56 163.367
R1101 B.n749 B.n61 163.367
R1102 B.n62 B.n61 163.367
R1103 B.n63 B.n62 163.367
R1104 B.n754 B.n63 163.367
R1105 B.n754 B.n68 163.367
R1106 B.n69 B.n68 163.367
R1107 B.n70 B.n69 163.367
R1108 B.n759 B.n70 163.367
R1109 B.n759 B.n75 163.367
R1110 B.n76 B.n75 163.367
R1111 B.n77 B.n76 163.367
R1112 B.n764 B.n77 163.367
R1113 B.n764 B.n82 163.367
R1114 B.n83 B.n82 163.367
R1115 B.n84 B.n83 163.367
R1116 B.n769 B.n84 163.367
R1117 B.n769 B.n89 163.367
R1118 B.n90 B.n89 163.367
R1119 B.n91 B.n90 163.367
R1120 B.n774 B.n91 163.367
R1121 B.n774 B.n96 163.367
R1122 B.n97 B.n96 163.367
R1123 B.n98 B.n97 163.367
R1124 B.n779 B.n98 163.367
R1125 B.n779 B.n103 163.367
R1126 B.n104 B.n103 163.367
R1127 B.n105 B.n104 163.367
R1128 B.n784 B.n105 163.367
R1129 B.n784 B.n110 163.367
R1130 B.n148 B.n147 163.367
R1131 B.n152 B.n151 163.367
R1132 B.n156 B.n155 163.367
R1133 B.n160 B.n159 163.367
R1134 B.n164 B.n163 163.367
R1135 B.n168 B.n167 163.367
R1136 B.n172 B.n171 163.367
R1137 B.n176 B.n175 163.367
R1138 B.n180 B.n179 163.367
R1139 B.n184 B.n183 163.367
R1140 B.n188 B.n187 163.367
R1141 B.n192 B.n191 163.367
R1142 B.n197 B.n196 163.367
R1143 B.n201 B.n200 163.367
R1144 B.n205 B.n204 163.367
R1145 B.n209 B.n208 163.367
R1146 B.n213 B.n212 163.367
R1147 B.n217 B.n216 163.367
R1148 B.n221 B.n220 163.367
R1149 B.n225 B.n224 163.367
R1150 B.n229 B.n228 163.367
R1151 B.n233 B.n232 163.367
R1152 B.n237 B.n236 163.367
R1153 B.n241 B.n240 163.367
R1154 B.n245 B.n244 163.367
R1155 B.n249 B.n248 163.367
R1156 B.n253 B.n252 163.367
R1157 B.n257 B.n256 163.367
R1158 B.n788 B.n140 163.367
R1159 B.n391 B.t13 129.796
R1160 B.n141 B.t16 129.796
R1161 B.n397 B.t23 129.788
R1162 B.n144 B.t19 129.788
R1163 B.n531 B.n377 116.891
R1164 B.n790 B.n789 116.891
R1165 B.n392 B.t12 72.7769
R1166 B.n142 B.t17 72.7769
R1167 B.n398 B.t22 72.7701
R1168 B.n145 B.t20 72.7701
R1169 B.n412 B.n376 71.676
R1170 B.n418 B.n417 71.676
R1171 B.n421 B.n420 71.676
R1172 B.n426 B.n425 71.676
R1173 B.n429 B.n428 71.676
R1174 B.n434 B.n433 71.676
R1175 B.n437 B.n436 71.676
R1176 B.n442 B.n441 71.676
R1177 B.n445 B.n444 71.676
R1178 B.n450 B.n449 71.676
R1179 B.n453 B.n452 71.676
R1180 B.n458 B.n457 71.676
R1181 B.n461 B.n460 71.676
R1182 B.n466 B.n465 71.676
R1183 B.n469 B.n468 71.676
R1184 B.n474 B.n473 71.676
R1185 B.n477 B.n476 71.676
R1186 B.n483 B.n482 71.676
R1187 B.n486 B.n485 71.676
R1188 B.n491 B.n490 71.676
R1189 B.n494 B.n493 71.676
R1190 B.n499 B.n498 71.676
R1191 B.n502 B.n501 71.676
R1192 B.n507 B.n506 71.676
R1193 B.n510 B.n509 71.676
R1194 B.n515 B.n514 71.676
R1195 B.n518 B.n517 71.676
R1196 B.n523 B.n522 71.676
R1197 B.n526 B.n525 71.676
R1198 B.n111 B.n109 71.676
R1199 B.n148 B.n112 71.676
R1200 B.n152 B.n113 71.676
R1201 B.n156 B.n114 71.676
R1202 B.n160 B.n115 71.676
R1203 B.n164 B.n116 71.676
R1204 B.n168 B.n117 71.676
R1205 B.n172 B.n118 71.676
R1206 B.n176 B.n119 71.676
R1207 B.n180 B.n120 71.676
R1208 B.n184 B.n121 71.676
R1209 B.n188 B.n122 71.676
R1210 B.n192 B.n123 71.676
R1211 B.n197 B.n124 71.676
R1212 B.n201 B.n125 71.676
R1213 B.n205 B.n126 71.676
R1214 B.n209 B.n127 71.676
R1215 B.n213 B.n128 71.676
R1216 B.n217 B.n129 71.676
R1217 B.n221 B.n130 71.676
R1218 B.n225 B.n131 71.676
R1219 B.n229 B.n132 71.676
R1220 B.n233 B.n133 71.676
R1221 B.n237 B.n134 71.676
R1222 B.n241 B.n135 71.676
R1223 B.n245 B.n136 71.676
R1224 B.n249 B.n137 71.676
R1225 B.n253 B.n138 71.676
R1226 B.n257 B.n139 71.676
R1227 B.n140 B.n139 71.676
R1228 B.n256 B.n138 71.676
R1229 B.n252 B.n137 71.676
R1230 B.n248 B.n136 71.676
R1231 B.n244 B.n135 71.676
R1232 B.n240 B.n134 71.676
R1233 B.n236 B.n133 71.676
R1234 B.n232 B.n132 71.676
R1235 B.n228 B.n131 71.676
R1236 B.n224 B.n130 71.676
R1237 B.n220 B.n129 71.676
R1238 B.n216 B.n128 71.676
R1239 B.n212 B.n127 71.676
R1240 B.n208 B.n126 71.676
R1241 B.n204 B.n125 71.676
R1242 B.n200 B.n124 71.676
R1243 B.n196 B.n123 71.676
R1244 B.n191 B.n122 71.676
R1245 B.n187 B.n121 71.676
R1246 B.n183 B.n120 71.676
R1247 B.n179 B.n119 71.676
R1248 B.n175 B.n118 71.676
R1249 B.n171 B.n117 71.676
R1250 B.n167 B.n116 71.676
R1251 B.n163 B.n115 71.676
R1252 B.n159 B.n114 71.676
R1253 B.n155 B.n113 71.676
R1254 B.n151 B.n112 71.676
R1255 B.n147 B.n111 71.676
R1256 B.n413 B.n412 71.676
R1257 B.n419 B.n418 71.676
R1258 B.n420 B.n409 71.676
R1259 B.n427 B.n426 71.676
R1260 B.n428 B.n407 71.676
R1261 B.n435 B.n434 71.676
R1262 B.n436 B.n405 71.676
R1263 B.n443 B.n442 71.676
R1264 B.n444 B.n403 71.676
R1265 B.n451 B.n450 71.676
R1266 B.n452 B.n401 71.676
R1267 B.n459 B.n458 71.676
R1268 B.n460 B.n396 71.676
R1269 B.n467 B.n466 71.676
R1270 B.n468 B.n394 71.676
R1271 B.n475 B.n474 71.676
R1272 B.n476 B.n390 71.676
R1273 B.n484 B.n483 71.676
R1274 B.n485 B.n388 71.676
R1275 B.n492 B.n491 71.676
R1276 B.n493 B.n386 71.676
R1277 B.n500 B.n499 71.676
R1278 B.n501 B.n384 71.676
R1279 B.n508 B.n507 71.676
R1280 B.n509 B.n382 71.676
R1281 B.n516 B.n515 71.676
R1282 B.n517 B.n380 71.676
R1283 B.n524 B.n523 71.676
R1284 B.n525 B.n378 71.676
R1285 B.n531 B.n373 64.6225
R1286 B.n537 B.n373 64.6225
R1287 B.n537 B.n369 64.6225
R1288 B.n543 B.n369 64.6225
R1289 B.n543 B.n364 64.6225
R1290 B.n549 B.n364 64.6225
R1291 B.n549 B.n365 64.6225
R1292 B.n555 B.n357 64.6225
R1293 B.n561 B.n357 64.6225
R1294 B.n561 B.n353 64.6225
R1295 B.n567 B.n353 64.6225
R1296 B.n567 B.n349 64.6225
R1297 B.n573 B.n349 64.6225
R1298 B.n573 B.n345 64.6225
R1299 B.n579 B.n345 64.6225
R1300 B.n579 B.n340 64.6225
R1301 B.n585 B.n340 64.6225
R1302 B.n585 B.n341 64.6225
R1303 B.n591 B.n333 64.6225
R1304 B.n597 B.n333 64.6225
R1305 B.n597 B.n329 64.6225
R1306 B.n603 B.n329 64.6225
R1307 B.n603 B.n325 64.6225
R1308 B.n609 B.n325 64.6225
R1309 B.n609 B.n321 64.6225
R1310 B.n615 B.n321 64.6225
R1311 B.n621 B.n317 64.6225
R1312 B.n621 B.n313 64.6225
R1313 B.n627 B.n313 64.6225
R1314 B.n627 B.n309 64.6225
R1315 B.n633 B.n309 64.6225
R1316 B.n633 B.n305 64.6225
R1317 B.n639 B.n305 64.6225
R1318 B.n645 B.n301 64.6225
R1319 B.n645 B.n297 64.6225
R1320 B.n651 B.n297 64.6225
R1321 B.n651 B.n293 64.6225
R1322 B.n657 B.n293 64.6225
R1323 B.n657 B.n289 64.6225
R1324 B.n664 B.n289 64.6225
R1325 B.n664 B.n663 64.6225
R1326 B.n670 B.n282 64.6225
R1327 B.n676 B.n282 64.6225
R1328 B.n676 B.n278 64.6225
R1329 B.n682 B.n278 64.6225
R1330 B.n682 B.n274 64.6225
R1331 B.n688 B.n274 64.6225
R1332 B.n688 B.n270 64.6225
R1333 B.n694 B.n270 64.6225
R1334 B.n701 B.n266 64.6225
R1335 B.n701 B.n262 64.6225
R1336 B.n707 B.n262 64.6225
R1337 B.n707 B.n4 64.6225
R1338 B.n910 B.n4 64.6225
R1339 B.n910 B.n909 64.6225
R1340 B.n909 B.n908 64.6225
R1341 B.n908 B.n8 64.6225
R1342 B.n902 B.n8 64.6225
R1343 B.n902 B.n901 64.6225
R1344 B.n900 B.n15 64.6225
R1345 B.n894 B.n15 64.6225
R1346 B.n894 B.n893 64.6225
R1347 B.n893 B.n892 64.6225
R1348 B.n892 B.n22 64.6225
R1349 B.n886 B.n22 64.6225
R1350 B.n886 B.n885 64.6225
R1351 B.n885 B.n884 64.6225
R1352 B.n878 B.n32 64.6225
R1353 B.n878 B.n877 64.6225
R1354 B.n877 B.n876 64.6225
R1355 B.n876 B.n36 64.6225
R1356 B.n870 B.n36 64.6225
R1357 B.n870 B.n869 64.6225
R1358 B.n869 B.n868 64.6225
R1359 B.n868 B.n43 64.6225
R1360 B.n862 B.n861 64.6225
R1361 B.n861 B.n860 64.6225
R1362 B.n860 B.n50 64.6225
R1363 B.n854 B.n50 64.6225
R1364 B.n854 B.n853 64.6225
R1365 B.n853 B.n852 64.6225
R1366 B.n852 B.n57 64.6225
R1367 B.n846 B.n845 64.6225
R1368 B.n845 B.n844 64.6225
R1369 B.n844 B.n64 64.6225
R1370 B.n838 B.n64 64.6225
R1371 B.n838 B.n837 64.6225
R1372 B.n837 B.n836 64.6225
R1373 B.n836 B.n71 64.6225
R1374 B.n830 B.n71 64.6225
R1375 B.n829 B.n828 64.6225
R1376 B.n828 B.n78 64.6225
R1377 B.n822 B.n78 64.6225
R1378 B.n822 B.n821 64.6225
R1379 B.n821 B.n820 64.6225
R1380 B.n820 B.n85 64.6225
R1381 B.n814 B.n85 64.6225
R1382 B.n814 B.n813 64.6225
R1383 B.n813 B.n812 64.6225
R1384 B.n812 B.n92 64.6225
R1385 B.n806 B.n92 64.6225
R1386 B.n805 B.n804 64.6225
R1387 B.n804 B.n99 64.6225
R1388 B.n798 B.n99 64.6225
R1389 B.n798 B.n797 64.6225
R1390 B.n797 B.n796 64.6225
R1391 B.n796 B.n106 64.6225
R1392 B.n790 B.n106 64.6225
R1393 B.t3 B.n266 59.8709
R1394 B.n901 B.t5 59.8709
R1395 B.n479 B.n392 59.5399
R1396 B.n399 B.n398 59.5399
R1397 B.n194 B.n145 59.5399
R1398 B.n143 B.n142 59.5399
R1399 B.n392 B.n391 57.0187
R1400 B.n398 B.n397 57.0187
R1401 B.n145 B.n144 57.0187
R1402 B.n142 B.n141 57.0187
R1403 B.t6 B.n317 56.0696
R1404 B.t0 B.n57 56.0696
R1405 B.n639 B.t4 50.3677
R1406 B.n862 B.t7 50.3677
R1407 B.n365 B.t11 40.8644
R1408 B.t15 B.n805 40.8644
R1409 B.n670 B.t2 37.0631
R1410 B.n884 B.t8 37.0631
R1411 B.n792 B.n108 33.8737
R1412 B.n787 B.n786 33.8737
R1413 B.n529 B.n528 33.8737
R1414 B.n533 B.n375 33.8737
R1415 B.n591 B.t9 33.2618
R1416 B.n830 B.t1 33.2618
R1417 B.n341 B.t9 31.3612
R1418 B.t1 B.n829 31.3612
R1419 B.n663 B.t2 27.5599
R1420 B.n32 B.t8 27.5599
R1421 B.n555 B.t11 23.7586
R1422 B.n806 B.t15 23.7586
R1423 B B.n912 18.0485
R1424 B.t4 B.n301 14.2554
R1425 B.t7 B.n43 14.2554
R1426 B.n146 B.n108 10.6151
R1427 B.n149 B.n146 10.6151
R1428 B.n150 B.n149 10.6151
R1429 B.n153 B.n150 10.6151
R1430 B.n154 B.n153 10.6151
R1431 B.n157 B.n154 10.6151
R1432 B.n158 B.n157 10.6151
R1433 B.n161 B.n158 10.6151
R1434 B.n162 B.n161 10.6151
R1435 B.n165 B.n162 10.6151
R1436 B.n166 B.n165 10.6151
R1437 B.n169 B.n166 10.6151
R1438 B.n170 B.n169 10.6151
R1439 B.n173 B.n170 10.6151
R1440 B.n174 B.n173 10.6151
R1441 B.n177 B.n174 10.6151
R1442 B.n178 B.n177 10.6151
R1443 B.n181 B.n178 10.6151
R1444 B.n182 B.n181 10.6151
R1445 B.n185 B.n182 10.6151
R1446 B.n186 B.n185 10.6151
R1447 B.n189 B.n186 10.6151
R1448 B.n190 B.n189 10.6151
R1449 B.n193 B.n190 10.6151
R1450 B.n198 B.n195 10.6151
R1451 B.n199 B.n198 10.6151
R1452 B.n202 B.n199 10.6151
R1453 B.n203 B.n202 10.6151
R1454 B.n206 B.n203 10.6151
R1455 B.n207 B.n206 10.6151
R1456 B.n210 B.n207 10.6151
R1457 B.n211 B.n210 10.6151
R1458 B.n215 B.n214 10.6151
R1459 B.n218 B.n215 10.6151
R1460 B.n219 B.n218 10.6151
R1461 B.n222 B.n219 10.6151
R1462 B.n223 B.n222 10.6151
R1463 B.n226 B.n223 10.6151
R1464 B.n227 B.n226 10.6151
R1465 B.n230 B.n227 10.6151
R1466 B.n231 B.n230 10.6151
R1467 B.n234 B.n231 10.6151
R1468 B.n235 B.n234 10.6151
R1469 B.n238 B.n235 10.6151
R1470 B.n239 B.n238 10.6151
R1471 B.n242 B.n239 10.6151
R1472 B.n243 B.n242 10.6151
R1473 B.n246 B.n243 10.6151
R1474 B.n247 B.n246 10.6151
R1475 B.n250 B.n247 10.6151
R1476 B.n251 B.n250 10.6151
R1477 B.n254 B.n251 10.6151
R1478 B.n255 B.n254 10.6151
R1479 B.n258 B.n255 10.6151
R1480 B.n259 B.n258 10.6151
R1481 B.n787 B.n259 10.6151
R1482 B.n529 B.n371 10.6151
R1483 B.n539 B.n371 10.6151
R1484 B.n540 B.n539 10.6151
R1485 B.n541 B.n540 10.6151
R1486 B.n541 B.n362 10.6151
R1487 B.n551 B.n362 10.6151
R1488 B.n552 B.n551 10.6151
R1489 B.n553 B.n552 10.6151
R1490 B.n553 B.n355 10.6151
R1491 B.n563 B.n355 10.6151
R1492 B.n564 B.n563 10.6151
R1493 B.n565 B.n564 10.6151
R1494 B.n565 B.n347 10.6151
R1495 B.n575 B.n347 10.6151
R1496 B.n576 B.n575 10.6151
R1497 B.n577 B.n576 10.6151
R1498 B.n577 B.n338 10.6151
R1499 B.n587 B.n338 10.6151
R1500 B.n588 B.n587 10.6151
R1501 B.n589 B.n588 10.6151
R1502 B.n589 B.n331 10.6151
R1503 B.n599 B.n331 10.6151
R1504 B.n600 B.n599 10.6151
R1505 B.n601 B.n600 10.6151
R1506 B.n601 B.n323 10.6151
R1507 B.n611 B.n323 10.6151
R1508 B.n612 B.n611 10.6151
R1509 B.n613 B.n612 10.6151
R1510 B.n613 B.n315 10.6151
R1511 B.n623 B.n315 10.6151
R1512 B.n624 B.n623 10.6151
R1513 B.n625 B.n624 10.6151
R1514 B.n625 B.n307 10.6151
R1515 B.n635 B.n307 10.6151
R1516 B.n636 B.n635 10.6151
R1517 B.n637 B.n636 10.6151
R1518 B.n637 B.n299 10.6151
R1519 B.n647 B.n299 10.6151
R1520 B.n648 B.n647 10.6151
R1521 B.n649 B.n648 10.6151
R1522 B.n649 B.n291 10.6151
R1523 B.n659 B.n291 10.6151
R1524 B.n660 B.n659 10.6151
R1525 B.n661 B.n660 10.6151
R1526 B.n661 B.n284 10.6151
R1527 B.n672 B.n284 10.6151
R1528 B.n673 B.n672 10.6151
R1529 B.n674 B.n673 10.6151
R1530 B.n674 B.n276 10.6151
R1531 B.n684 B.n276 10.6151
R1532 B.n685 B.n684 10.6151
R1533 B.n686 B.n685 10.6151
R1534 B.n686 B.n268 10.6151
R1535 B.n696 B.n268 10.6151
R1536 B.n697 B.n696 10.6151
R1537 B.n699 B.n697 10.6151
R1538 B.n699 B.n698 10.6151
R1539 B.n698 B.n260 10.6151
R1540 B.n710 B.n260 10.6151
R1541 B.n711 B.n710 10.6151
R1542 B.n712 B.n711 10.6151
R1543 B.n713 B.n712 10.6151
R1544 B.n715 B.n713 10.6151
R1545 B.n716 B.n715 10.6151
R1546 B.n717 B.n716 10.6151
R1547 B.n718 B.n717 10.6151
R1548 B.n720 B.n718 10.6151
R1549 B.n721 B.n720 10.6151
R1550 B.n722 B.n721 10.6151
R1551 B.n723 B.n722 10.6151
R1552 B.n725 B.n723 10.6151
R1553 B.n726 B.n725 10.6151
R1554 B.n727 B.n726 10.6151
R1555 B.n728 B.n727 10.6151
R1556 B.n730 B.n728 10.6151
R1557 B.n731 B.n730 10.6151
R1558 B.n732 B.n731 10.6151
R1559 B.n733 B.n732 10.6151
R1560 B.n735 B.n733 10.6151
R1561 B.n736 B.n735 10.6151
R1562 B.n737 B.n736 10.6151
R1563 B.n738 B.n737 10.6151
R1564 B.n740 B.n738 10.6151
R1565 B.n741 B.n740 10.6151
R1566 B.n742 B.n741 10.6151
R1567 B.n743 B.n742 10.6151
R1568 B.n745 B.n743 10.6151
R1569 B.n746 B.n745 10.6151
R1570 B.n747 B.n746 10.6151
R1571 B.n748 B.n747 10.6151
R1572 B.n750 B.n748 10.6151
R1573 B.n751 B.n750 10.6151
R1574 B.n752 B.n751 10.6151
R1575 B.n753 B.n752 10.6151
R1576 B.n755 B.n753 10.6151
R1577 B.n756 B.n755 10.6151
R1578 B.n757 B.n756 10.6151
R1579 B.n758 B.n757 10.6151
R1580 B.n760 B.n758 10.6151
R1581 B.n761 B.n760 10.6151
R1582 B.n762 B.n761 10.6151
R1583 B.n763 B.n762 10.6151
R1584 B.n765 B.n763 10.6151
R1585 B.n766 B.n765 10.6151
R1586 B.n767 B.n766 10.6151
R1587 B.n768 B.n767 10.6151
R1588 B.n770 B.n768 10.6151
R1589 B.n771 B.n770 10.6151
R1590 B.n772 B.n771 10.6151
R1591 B.n773 B.n772 10.6151
R1592 B.n775 B.n773 10.6151
R1593 B.n776 B.n775 10.6151
R1594 B.n777 B.n776 10.6151
R1595 B.n778 B.n777 10.6151
R1596 B.n780 B.n778 10.6151
R1597 B.n781 B.n780 10.6151
R1598 B.n782 B.n781 10.6151
R1599 B.n783 B.n782 10.6151
R1600 B.n785 B.n783 10.6151
R1601 B.n786 B.n785 10.6151
R1602 B.n414 B.n375 10.6151
R1603 B.n415 B.n414 10.6151
R1604 B.n416 B.n415 10.6151
R1605 B.n416 B.n410 10.6151
R1606 B.n422 B.n410 10.6151
R1607 B.n423 B.n422 10.6151
R1608 B.n424 B.n423 10.6151
R1609 B.n424 B.n408 10.6151
R1610 B.n430 B.n408 10.6151
R1611 B.n431 B.n430 10.6151
R1612 B.n432 B.n431 10.6151
R1613 B.n432 B.n406 10.6151
R1614 B.n438 B.n406 10.6151
R1615 B.n439 B.n438 10.6151
R1616 B.n440 B.n439 10.6151
R1617 B.n440 B.n404 10.6151
R1618 B.n446 B.n404 10.6151
R1619 B.n447 B.n446 10.6151
R1620 B.n448 B.n447 10.6151
R1621 B.n448 B.n402 10.6151
R1622 B.n454 B.n402 10.6151
R1623 B.n455 B.n454 10.6151
R1624 B.n456 B.n455 10.6151
R1625 B.n456 B.n400 10.6151
R1626 B.n463 B.n462 10.6151
R1627 B.n464 B.n463 10.6151
R1628 B.n464 B.n395 10.6151
R1629 B.n470 B.n395 10.6151
R1630 B.n471 B.n470 10.6151
R1631 B.n472 B.n471 10.6151
R1632 B.n472 B.n393 10.6151
R1633 B.n478 B.n393 10.6151
R1634 B.n481 B.n480 10.6151
R1635 B.n481 B.n389 10.6151
R1636 B.n487 B.n389 10.6151
R1637 B.n488 B.n487 10.6151
R1638 B.n489 B.n488 10.6151
R1639 B.n489 B.n387 10.6151
R1640 B.n495 B.n387 10.6151
R1641 B.n496 B.n495 10.6151
R1642 B.n497 B.n496 10.6151
R1643 B.n497 B.n385 10.6151
R1644 B.n503 B.n385 10.6151
R1645 B.n504 B.n503 10.6151
R1646 B.n505 B.n504 10.6151
R1647 B.n505 B.n383 10.6151
R1648 B.n511 B.n383 10.6151
R1649 B.n512 B.n511 10.6151
R1650 B.n513 B.n512 10.6151
R1651 B.n513 B.n381 10.6151
R1652 B.n519 B.n381 10.6151
R1653 B.n520 B.n519 10.6151
R1654 B.n521 B.n520 10.6151
R1655 B.n521 B.n379 10.6151
R1656 B.n527 B.n379 10.6151
R1657 B.n528 B.n527 10.6151
R1658 B.n534 B.n533 10.6151
R1659 B.n535 B.n534 10.6151
R1660 B.n535 B.n367 10.6151
R1661 B.n545 B.n367 10.6151
R1662 B.n546 B.n545 10.6151
R1663 B.n547 B.n546 10.6151
R1664 B.n547 B.n359 10.6151
R1665 B.n557 B.n359 10.6151
R1666 B.n558 B.n557 10.6151
R1667 B.n559 B.n558 10.6151
R1668 B.n559 B.n351 10.6151
R1669 B.n569 B.n351 10.6151
R1670 B.n570 B.n569 10.6151
R1671 B.n571 B.n570 10.6151
R1672 B.n571 B.n343 10.6151
R1673 B.n581 B.n343 10.6151
R1674 B.n582 B.n581 10.6151
R1675 B.n583 B.n582 10.6151
R1676 B.n583 B.n335 10.6151
R1677 B.n593 B.n335 10.6151
R1678 B.n594 B.n593 10.6151
R1679 B.n595 B.n594 10.6151
R1680 B.n595 B.n327 10.6151
R1681 B.n605 B.n327 10.6151
R1682 B.n606 B.n605 10.6151
R1683 B.n607 B.n606 10.6151
R1684 B.n607 B.n319 10.6151
R1685 B.n617 B.n319 10.6151
R1686 B.n618 B.n617 10.6151
R1687 B.n619 B.n618 10.6151
R1688 B.n619 B.n311 10.6151
R1689 B.n629 B.n311 10.6151
R1690 B.n630 B.n629 10.6151
R1691 B.n631 B.n630 10.6151
R1692 B.n631 B.n303 10.6151
R1693 B.n641 B.n303 10.6151
R1694 B.n642 B.n641 10.6151
R1695 B.n643 B.n642 10.6151
R1696 B.n643 B.n295 10.6151
R1697 B.n653 B.n295 10.6151
R1698 B.n654 B.n653 10.6151
R1699 B.n655 B.n654 10.6151
R1700 B.n655 B.n287 10.6151
R1701 B.n666 B.n287 10.6151
R1702 B.n667 B.n666 10.6151
R1703 B.n668 B.n667 10.6151
R1704 B.n668 B.n280 10.6151
R1705 B.n678 B.n280 10.6151
R1706 B.n679 B.n678 10.6151
R1707 B.n680 B.n679 10.6151
R1708 B.n680 B.n272 10.6151
R1709 B.n690 B.n272 10.6151
R1710 B.n691 B.n690 10.6151
R1711 B.n692 B.n691 10.6151
R1712 B.n692 B.n264 10.6151
R1713 B.n703 B.n264 10.6151
R1714 B.n704 B.n703 10.6151
R1715 B.n705 B.n704 10.6151
R1716 B.n705 B.n0 10.6151
R1717 B.n906 B.n1 10.6151
R1718 B.n906 B.n905 10.6151
R1719 B.n905 B.n904 10.6151
R1720 B.n904 B.n10 10.6151
R1721 B.n898 B.n10 10.6151
R1722 B.n898 B.n897 10.6151
R1723 B.n897 B.n896 10.6151
R1724 B.n896 B.n17 10.6151
R1725 B.n890 B.n17 10.6151
R1726 B.n890 B.n889 10.6151
R1727 B.n889 B.n888 10.6151
R1728 B.n888 B.n24 10.6151
R1729 B.n882 B.n24 10.6151
R1730 B.n882 B.n881 10.6151
R1731 B.n881 B.n880 10.6151
R1732 B.n880 B.n30 10.6151
R1733 B.n874 B.n30 10.6151
R1734 B.n874 B.n873 10.6151
R1735 B.n873 B.n872 10.6151
R1736 B.n872 B.n38 10.6151
R1737 B.n866 B.n38 10.6151
R1738 B.n866 B.n865 10.6151
R1739 B.n865 B.n864 10.6151
R1740 B.n864 B.n45 10.6151
R1741 B.n858 B.n45 10.6151
R1742 B.n858 B.n857 10.6151
R1743 B.n857 B.n856 10.6151
R1744 B.n856 B.n52 10.6151
R1745 B.n850 B.n52 10.6151
R1746 B.n850 B.n849 10.6151
R1747 B.n849 B.n848 10.6151
R1748 B.n848 B.n59 10.6151
R1749 B.n842 B.n59 10.6151
R1750 B.n842 B.n841 10.6151
R1751 B.n841 B.n840 10.6151
R1752 B.n840 B.n66 10.6151
R1753 B.n834 B.n66 10.6151
R1754 B.n834 B.n833 10.6151
R1755 B.n833 B.n832 10.6151
R1756 B.n832 B.n73 10.6151
R1757 B.n826 B.n73 10.6151
R1758 B.n826 B.n825 10.6151
R1759 B.n825 B.n824 10.6151
R1760 B.n824 B.n80 10.6151
R1761 B.n818 B.n80 10.6151
R1762 B.n818 B.n817 10.6151
R1763 B.n817 B.n816 10.6151
R1764 B.n816 B.n87 10.6151
R1765 B.n810 B.n87 10.6151
R1766 B.n810 B.n809 10.6151
R1767 B.n809 B.n808 10.6151
R1768 B.n808 B.n94 10.6151
R1769 B.n802 B.n94 10.6151
R1770 B.n802 B.n801 10.6151
R1771 B.n801 B.n800 10.6151
R1772 B.n800 B.n101 10.6151
R1773 B.n794 B.n101 10.6151
R1774 B.n794 B.n793 10.6151
R1775 B.n793 B.n792 10.6151
R1776 B.n615 B.t6 8.55342
R1777 B.n846 B.t0 8.55342
R1778 B.n195 B.n194 6.5566
R1779 B.n211 B.n143 6.5566
R1780 B.n462 B.n399 6.5566
R1781 B.n479 B.n478 6.5566
R1782 B.n694 B.t3 4.75212
R1783 B.t5 B.n900 4.75212
R1784 B.n194 B.n193 4.05904
R1785 B.n214 B.n143 4.05904
R1786 B.n400 B.n399 4.05904
R1787 B.n480 B.n479 4.05904
R1788 B.n912 B.n0 2.81026
R1789 B.n912 B.n1 2.81026
R1790 VP.n25 VP.n22 161.3
R1791 VP.n27 VP.n26 161.3
R1792 VP.n28 VP.n21 161.3
R1793 VP.n30 VP.n29 161.3
R1794 VP.n31 VP.n20 161.3
R1795 VP.n33 VP.n32 161.3
R1796 VP.n35 VP.n19 161.3
R1797 VP.n37 VP.n36 161.3
R1798 VP.n38 VP.n18 161.3
R1799 VP.n40 VP.n39 161.3
R1800 VP.n41 VP.n17 161.3
R1801 VP.n43 VP.n42 161.3
R1802 VP.n45 VP.n44 161.3
R1803 VP.n46 VP.n15 161.3
R1804 VP.n48 VP.n47 161.3
R1805 VP.n49 VP.n14 161.3
R1806 VP.n51 VP.n50 161.3
R1807 VP.n52 VP.n13 161.3
R1808 VP.n94 VP.n0 161.3
R1809 VP.n93 VP.n92 161.3
R1810 VP.n91 VP.n1 161.3
R1811 VP.n90 VP.n89 161.3
R1812 VP.n88 VP.n2 161.3
R1813 VP.n87 VP.n86 161.3
R1814 VP.n85 VP.n84 161.3
R1815 VP.n83 VP.n4 161.3
R1816 VP.n82 VP.n81 161.3
R1817 VP.n80 VP.n5 161.3
R1818 VP.n79 VP.n78 161.3
R1819 VP.n77 VP.n6 161.3
R1820 VP.n75 VP.n74 161.3
R1821 VP.n73 VP.n7 161.3
R1822 VP.n72 VP.n71 161.3
R1823 VP.n70 VP.n8 161.3
R1824 VP.n69 VP.n68 161.3
R1825 VP.n67 VP.n9 161.3
R1826 VP.n66 VP.n65 161.3
R1827 VP.n63 VP.n10 161.3
R1828 VP.n62 VP.n61 161.3
R1829 VP.n60 VP.n11 161.3
R1830 VP.n59 VP.n58 161.3
R1831 VP.n57 VP.n12 161.3
R1832 VP.n56 VP.n55 104.514
R1833 VP.n96 VP.n95 104.514
R1834 VP.n54 VP.n53 104.514
R1835 VP.n24 VP.t7 90.7511
R1836 VP.n24 VP.n23 63.1649
R1837 VP.n56 VP.t2 58.1729
R1838 VP.n64 VP.t3 58.1729
R1839 VP.n76 VP.t1 58.1729
R1840 VP.n3 VP.t6 58.1729
R1841 VP.n95 VP.t4 58.1729
R1842 VP.n53 VP.t5 58.1729
R1843 VP.n16 VP.t8 58.1729
R1844 VP.n34 VP.t0 58.1729
R1845 VP.n23 VP.t9 58.1729
R1846 VP.n71 VP.n70 56.5617
R1847 VP.n82 VP.n5 56.5617
R1848 VP.n40 VP.n18 56.5617
R1849 VP.n29 VP.n28 56.5617
R1850 VP.n62 VP.n11 56.0773
R1851 VP.n89 VP.n1 56.0773
R1852 VP.n47 VP.n14 56.0773
R1853 VP.n55 VP.n54 48.8178
R1854 VP.n63 VP.n62 25.0767
R1855 VP.n89 VP.n88 25.0767
R1856 VP.n47 VP.n46 25.0767
R1857 VP.n58 VP.n57 24.5923
R1858 VP.n58 VP.n11 24.5923
R1859 VP.n65 VP.n63 24.5923
R1860 VP.n69 VP.n9 24.5923
R1861 VP.n70 VP.n69 24.5923
R1862 VP.n71 VP.n7 24.5923
R1863 VP.n75 VP.n7 24.5923
R1864 VP.n78 VP.n77 24.5923
R1865 VP.n78 VP.n5 24.5923
R1866 VP.n83 VP.n82 24.5923
R1867 VP.n84 VP.n83 24.5923
R1868 VP.n88 VP.n87 24.5923
R1869 VP.n93 VP.n1 24.5923
R1870 VP.n94 VP.n93 24.5923
R1871 VP.n51 VP.n14 24.5923
R1872 VP.n52 VP.n51 24.5923
R1873 VP.n41 VP.n40 24.5923
R1874 VP.n42 VP.n41 24.5923
R1875 VP.n46 VP.n45 24.5923
R1876 VP.n29 VP.n20 24.5923
R1877 VP.n33 VP.n20 24.5923
R1878 VP.n36 VP.n35 24.5923
R1879 VP.n36 VP.n18 24.5923
R1880 VP.n27 VP.n22 24.5923
R1881 VP.n28 VP.n27 24.5923
R1882 VP.n65 VP.n64 15.2474
R1883 VP.n87 VP.n3 15.2474
R1884 VP.n45 VP.n16 15.2474
R1885 VP.n76 VP.n75 12.2964
R1886 VP.n77 VP.n76 12.2964
R1887 VP.n34 VP.n33 12.2964
R1888 VP.n35 VP.n34 12.2964
R1889 VP.n64 VP.n9 9.3454
R1890 VP.n84 VP.n3 9.3454
R1891 VP.n42 VP.n16 9.3454
R1892 VP.n23 VP.n22 9.3454
R1893 VP.n25 VP.n24 7.05922
R1894 VP.n57 VP.n56 6.39438
R1895 VP.n95 VP.n94 6.39438
R1896 VP.n53 VP.n52 6.39438
R1897 VP.n54 VP.n13 0.278335
R1898 VP.n55 VP.n12 0.278335
R1899 VP.n96 VP.n0 0.278335
R1900 VP.n26 VP.n25 0.189894
R1901 VP.n26 VP.n21 0.189894
R1902 VP.n30 VP.n21 0.189894
R1903 VP.n31 VP.n30 0.189894
R1904 VP.n32 VP.n31 0.189894
R1905 VP.n32 VP.n19 0.189894
R1906 VP.n37 VP.n19 0.189894
R1907 VP.n38 VP.n37 0.189894
R1908 VP.n39 VP.n38 0.189894
R1909 VP.n39 VP.n17 0.189894
R1910 VP.n43 VP.n17 0.189894
R1911 VP.n44 VP.n43 0.189894
R1912 VP.n44 VP.n15 0.189894
R1913 VP.n48 VP.n15 0.189894
R1914 VP.n49 VP.n48 0.189894
R1915 VP.n50 VP.n49 0.189894
R1916 VP.n50 VP.n13 0.189894
R1917 VP.n59 VP.n12 0.189894
R1918 VP.n60 VP.n59 0.189894
R1919 VP.n61 VP.n60 0.189894
R1920 VP.n61 VP.n10 0.189894
R1921 VP.n66 VP.n10 0.189894
R1922 VP.n67 VP.n66 0.189894
R1923 VP.n68 VP.n67 0.189894
R1924 VP.n68 VP.n8 0.189894
R1925 VP.n72 VP.n8 0.189894
R1926 VP.n73 VP.n72 0.189894
R1927 VP.n74 VP.n73 0.189894
R1928 VP.n74 VP.n6 0.189894
R1929 VP.n79 VP.n6 0.189894
R1930 VP.n80 VP.n79 0.189894
R1931 VP.n81 VP.n80 0.189894
R1932 VP.n81 VP.n4 0.189894
R1933 VP.n85 VP.n4 0.189894
R1934 VP.n86 VP.n85 0.189894
R1935 VP.n86 VP.n2 0.189894
R1936 VP.n90 VP.n2 0.189894
R1937 VP.n91 VP.n90 0.189894
R1938 VP.n92 VP.n91 0.189894
R1939 VP.n92 VP.n0 0.189894
R1940 VP VP.n96 0.153485
R1941 VDD1.n1 VDD1.t2 71.1097
R1942 VDD1.n3 VDD1.t7 71.1096
R1943 VDD1.n5 VDD1.n4 67.2777
R1944 VDD1.n1 VDD1.n0 65.4324
R1945 VDD1.n7 VDD1.n6 65.4322
R1946 VDD1.n3 VDD1.n2 65.4322
R1947 VDD1.n7 VDD1.n5 43.0354
R1948 VDD1.n6 VDD1.t1 3.14336
R1949 VDD1.n6 VDD1.t4 3.14336
R1950 VDD1.n0 VDD1.t0 3.14336
R1951 VDD1.n0 VDD1.t9 3.14336
R1952 VDD1.n4 VDD1.t3 3.14336
R1953 VDD1.n4 VDD1.t5 3.14336
R1954 VDD1.n2 VDD1.t6 3.14336
R1955 VDD1.n2 VDD1.t8 3.14336
R1956 VDD1 VDD1.n7 1.84317
R1957 VDD1 VDD1.n1 0.69231
R1958 VDD1.n5 VDD1.n3 0.578775
C0 VTAIL VN 6.94837f
C1 VDD1 VDD2 2.18124f
C2 VP VDD2 0.584875f
C3 VN VDD2 5.84919f
C4 VP VDD1 6.27735f
C5 VN VDD1 0.153857f
C6 VN VP 7.35189f
C7 VTAIL VDD2 7.82366f
C8 VTAIL VDD1 7.77132f
C9 VTAIL VP 6.96257f
C10 VDD2 B 6.269975f
C11 VDD1 B 6.19837f
C12 VTAIL B 5.513348f
C13 VN B 17.53378f
C14 VP B 16.098946f
C15 VDD1.t2 B 1.42696f
C16 VDD1.t0 B 0.132316f
C17 VDD1.t9 B 0.132316f
C18 VDD1.n0 B 1.10937f
C19 VDD1.n1 B 0.981852f
C20 VDD1.t7 B 1.42695f
C21 VDD1.t6 B 0.132316f
C22 VDD1.t8 B 0.132316f
C23 VDD1.n2 B 1.10936f
C24 VDD1.n3 B 0.973205f
C25 VDD1.t3 B 0.132316f
C26 VDD1.t5 B 0.132316f
C27 VDD1.n4 B 1.12591f
C28 VDD1.n5 B 2.85248f
C29 VDD1.t1 B 0.132316f
C30 VDD1.t4 B 0.132316f
C31 VDD1.n6 B 1.10936f
C32 VDD1.n7 B 2.90898f
C33 VP.n0 B 0.032121f
C34 VP.t4 B 1.06337f
C35 VP.n1 B 0.041426f
C36 VP.n2 B 0.024365f
C37 VP.t6 B 1.06337f
C38 VP.n3 B 0.396563f
C39 VP.n4 B 0.024365f
C40 VP.n5 B 0.033396f
C41 VP.n6 B 0.024365f
C42 VP.t1 B 1.06337f
C43 VP.n7 B 0.045183f
C44 VP.n8 B 0.024365f
C45 VP.n9 B 0.031353f
C46 VP.n10 B 0.024365f
C47 VP.n11 B 0.041426f
C48 VP.n12 B 0.032121f
C49 VP.t2 B 1.06337f
C50 VP.n13 B 0.032121f
C51 VP.t5 B 1.06337f
C52 VP.n14 B 0.041426f
C53 VP.n15 B 0.024365f
C54 VP.t8 B 1.06337f
C55 VP.n16 B 0.396563f
C56 VP.n17 B 0.024365f
C57 VP.n18 B 0.033396f
C58 VP.n19 B 0.024365f
C59 VP.t0 B 1.06337f
C60 VP.n20 B 0.045183f
C61 VP.n21 B 0.024365f
C62 VP.n22 B 0.031353f
C63 VP.t7 B 1.2592f
C64 VP.t9 B 1.06337f
C65 VP.n23 B 0.463926f
C66 VP.n24 B 0.450314f
C67 VP.n25 B 0.235554f
C68 VP.n26 B 0.024365f
C69 VP.n27 B 0.045183f
C70 VP.n28 B 0.037441f
C71 VP.n29 B 0.033396f
C72 VP.n30 B 0.024365f
C73 VP.n31 B 0.024365f
C74 VP.n32 B 0.024365f
C75 VP.n33 B 0.03403f
C76 VP.n34 B 0.396563f
C77 VP.n35 B 0.03403f
C78 VP.n36 B 0.045183f
C79 VP.n37 B 0.024365f
C80 VP.n38 B 0.024365f
C81 VP.n39 B 0.024365f
C82 VP.n40 B 0.037441f
C83 VP.n41 B 0.045183f
C84 VP.n42 B 0.031353f
C85 VP.n43 B 0.024365f
C86 VP.n44 B 0.024365f
C87 VP.n45 B 0.036707f
C88 VP.n46 B 0.045605f
C89 VP.n47 B 0.028989f
C90 VP.n48 B 0.024365f
C91 VP.n49 B 0.024365f
C92 VP.n50 B 0.024365f
C93 VP.n51 B 0.045183f
C94 VP.n52 B 0.028677f
C95 VP.n53 B 0.473297f
C96 VP.n54 B 1.3104f
C97 VP.n55 B 1.3284f
C98 VP.n56 B 0.473297f
C99 VP.n57 B 0.028677f
C100 VP.n58 B 0.045183f
C101 VP.n59 B 0.024365f
C102 VP.n60 B 0.024365f
C103 VP.n61 B 0.024365f
C104 VP.n62 B 0.028989f
C105 VP.n63 B 0.045605f
C106 VP.t3 B 1.06337f
C107 VP.n64 B 0.396563f
C108 VP.n65 B 0.036707f
C109 VP.n66 B 0.024365f
C110 VP.n67 B 0.024365f
C111 VP.n68 B 0.024365f
C112 VP.n69 B 0.045183f
C113 VP.n70 B 0.037441f
C114 VP.n71 B 0.033396f
C115 VP.n72 B 0.024365f
C116 VP.n73 B 0.024365f
C117 VP.n74 B 0.024365f
C118 VP.n75 B 0.03403f
C119 VP.n76 B 0.396563f
C120 VP.n77 B 0.03403f
C121 VP.n78 B 0.045183f
C122 VP.n79 B 0.024365f
C123 VP.n80 B 0.024365f
C124 VP.n81 B 0.024365f
C125 VP.n82 B 0.037441f
C126 VP.n83 B 0.045183f
C127 VP.n84 B 0.031353f
C128 VP.n85 B 0.024365f
C129 VP.n86 B 0.024365f
C130 VP.n87 B 0.036707f
C131 VP.n88 B 0.045605f
C132 VP.n89 B 0.028989f
C133 VP.n90 B 0.024365f
C134 VP.n91 B 0.024365f
C135 VP.n92 B 0.024365f
C136 VP.n93 B 0.045183f
C137 VP.n94 B 0.028677f
C138 VP.n95 B 0.473297f
C139 VP.n96 B 0.041826f
C140 VDD2.t6 B 1.39156f
C141 VDD2.t4 B 0.129034f
C142 VDD2.t9 B 0.129034f
C143 VDD2.n0 B 1.08185f
C144 VDD2.n1 B 0.949068f
C145 VDD2.t7 B 0.129034f
C146 VDD2.t5 B 0.129034f
C147 VDD2.n2 B 1.09799f
C148 VDD2.n3 B 2.65656f
C149 VDD2.t2 B 1.37397f
C150 VDD2.n4 B 2.77218f
C151 VDD2.t8 B 0.129034f
C152 VDD2.t0 B 0.129034f
C153 VDD2.n5 B 1.08185f
C154 VDD2.n6 B 0.481321f
C155 VDD2.t1 B 0.129034f
C156 VDD2.t3 B 0.129034f
C157 VDD2.n7 B 1.09795f
C158 VTAIL.t18 B 0.140806f
C159 VTAIL.t14 B 0.140806f
C160 VTAIL.n0 B 1.10329f
C161 VTAIL.n1 B 0.606867f
C162 VTAIL.t3 B 1.40576f
C163 VTAIL.n2 B 0.740855f
C164 VTAIL.t4 B 0.140806f
C165 VTAIL.t2 B 0.140806f
C166 VTAIL.n3 B 1.10329f
C167 VTAIL.n4 B 0.731981f
C168 VTAIL.t9 B 0.140806f
C169 VTAIL.t6 B 0.140806f
C170 VTAIL.n5 B 1.10329f
C171 VTAIL.n6 B 1.8421f
C172 VTAIL.t15 B 0.140806f
C173 VTAIL.t19 B 0.140806f
C174 VTAIL.n7 B 1.10329f
C175 VTAIL.n8 B 1.8421f
C176 VTAIL.t16 B 0.140806f
C177 VTAIL.t11 B 0.140806f
C178 VTAIL.n9 B 1.10329f
C179 VTAIL.n10 B 0.731974f
C180 VTAIL.t13 B 1.40576f
C181 VTAIL.n11 B 0.740846f
C182 VTAIL.t5 B 0.140806f
C183 VTAIL.t8 B 0.140806f
C184 VTAIL.n12 B 1.10329f
C185 VTAIL.n13 B 0.659303f
C186 VTAIL.t7 B 0.140806f
C187 VTAIL.t0 B 0.140806f
C188 VTAIL.n14 B 1.10329f
C189 VTAIL.n15 B 0.731974f
C190 VTAIL.t1 B 1.40576f
C191 VTAIL.n16 B 1.69267f
C192 VTAIL.t10 B 1.40576f
C193 VTAIL.n17 B 1.69267f
C194 VTAIL.t12 B 0.140806f
C195 VTAIL.t17 B 0.140806f
C196 VTAIL.n18 B 1.10329f
C197 VTAIL.n19 B 0.553444f
C198 VN.n0 B 0.031139f
C199 VN.t4 B 1.03084f
C200 VN.n1 B 0.040159f
C201 VN.n2 B 0.02362f
C202 VN.t2 B 1.03084f
C203 VN.n3 B 0.384432f
C204 VN.n4 B 0.02362f
C205 VN.n5 B 0.032375f
C206 VN.n6 B 0.02362f
C207 VN.t0 B 1.03084f
C208 VN.n7 B 0.043801f
C209 VN.n8 B 0.02362f
C210 VN.n9 B 0.030394f
C211 VN.t3 B 1.22068f
C212 VN.t5 B 1.03084f
C213 VN.n10 B 0.449735f
C214 VN.n11 B 0.436539f
C215 VN.n12 B 0.228349f
C216 VN.n13 B 0.02362f
C217 VN.n14 B 0.043801f
C218 VN.n15 B 0.036296f
C219 VN.n16 B 0.032375f
C220 VN.n17 B 0.02362f
C221 VN.n18 B 0.02362f
C222 VN.n19 B 0.02362f
C223 VN.n20 B 0.032989f
C224 VN.n21 B 0.384432f
C225 VN.n22 B 0.032989f
C226 VN.n23 B 0.043801f
C227 VN.n24 B 0.02362f
C228 VN.n25 B 0.02362f
C229 VN.n26 B 0.02362f
C230 VN.n27 B 0.036296f
C231 VN.n28 B 0.043801f
C232 VN.n29 B 0.030394f
C233 VN.n30 B 0.02362f
C234 VN.n31 B 0.02362f
C235 VN.n32 B 0.035584f
C236 VN.n33 B 0.04421f
C237 VN.n34 B 0.028102f
C238 VN.n35 B 0.02362f
C239 VN.n36 B 0.02362f
C240 VN.n37 B 0.02362f
C241 VN.n38 B 0.043801f
C242 VN.n39 B 0.0278f
C243 VN.n40 B 0.458819f
C244 VN.n41 B 0.040547f
C245 VN.n42 B 0.031139f
C246 VN.t7 B 1.03084f
C247 VN.n43 B 0.040159f
C248 VN.n44 B 0.02362f
C249 VN.t1 B 1.03084f
C250 VN.n45 B 0.384432f
C251 VN.n46 B 0.02362f
C252 VN.n47 B 0.032375f
C253 VN.n48 B 0.02362f
C254 VN.t9 B 1.03084f
C255 VN.n49 B 0.043801f
C256 VN.n50 B 0.02362f
C257 VN.n51 B 0.030394f
C258 VN.t6 B 1.22068f
C259 VN.t8 B 1.03084f
C260 VN.n52 B 0.449735f
C261 VN.n53 B 0.436539f
C262 VN.n54 B 0.228349f
C263 VN.n55 B 0.02362f
C264 VN.n56 B 0.043801f
C265 VN.n57 B 0.036296f
C266 VN.n58 B 0.032375f
C267 VN.n59 B 0.02362f
C268 VN.n60 B 0.02362f
C269 VN.n61 B 0.02362f
C270 VN.n62 B 0.032989f
C271 VN.n63 B 0.384432f
C272 VN.n64 B 0.032989f
C273 VN.n65 B 0.043801f
C274 VN.n66 B 0.02362f
C275 VN.n67 B 0.02362f
C276 VN.n68 B 0.02362f
C277 VN.n69 B 0.036296f
C278 VN.n70 B 0.043801f
C279 VN.n71 B 0.030394f
C280 VN.n72 B 0.02362f
C281 VN.n73 B 0.02362f
C282 VN.n74 B 0.035584f
C283 VN.n75 B 0.04421f
C284 VN.n76 B 0.028102f
C285 VN.n77 B 0.02362f
C286 VN.n78 B 0.02362f
C287 VN.n79 B 0.02362f
C288 VN.n80 B 0.043801f
C289 VN.n81 B 0.0278f
C290 VN.n82 B 0.458819f
C291 VN.n83 B 1.28306f
.ends

