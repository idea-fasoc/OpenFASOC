* NGSPICE file created from diff_pair_sample_1625.ext - technology: sky130A

.subckt diff_pair_sample_1625 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t17 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X1 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X2 VDD1.t8 VP.t1 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X3 VDD2.t8 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X4 VDD1.t7 VP.t2 VTAIL.t16 B.t0 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.62
X5 VDD2.t7 VN.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.62
X6 VDD1.t6 VP.t3 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.62
X7 B.t22 B.t20 B.t21 B.t10 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.62
X8 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.62
X9 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.62
X10 VTAIL.t9 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X11 VDD2.t6 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X12 VTAIL.t7 VN.t4 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X13 VTAIL.t13 VP.t5 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X14 VTAIL.t8 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X15 VDD1.t3 VP.t6 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.62
X16 VTAIL.t15 VP.t7 VDD1.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X17 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.62
X18 VDD2.t2 VN.t7 VTAIL.t19 B.t23 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.62
X19 VTAIL.t2 VN.t8 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X20 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=0 ps=0 w=11.11 l=3.62
X21 VTAIL.t10 VP.t8 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=1.83315 ps=11.44 w=11.11 l=3.62
X22 VDD1.t0 VP.t9 VTAIL.t14 B.t23 sky130_fd_pr__nfet_01v8 ad=4.3329 pd=23 as=1.83315 ps=11.44 w=11.11 l=3.62
X23 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.83315 pd=11.44 as=4.3329 ps=23 w=11.11 l=3.62
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n31 VP.t6 106.894
R57 VP.n72 VP.n71 82.7273
R58 VP.n124 VP.n0 82.7273
R59 VP.n70 VP.n17 82.7273
R60 VP.n71 VP.t9 73.9649
R61 VP.n83 VP.t5 73.9649
R62 VP.n96 VP.t1 73.9649
R63 VP.n109 VP.t8 73.9649
R64 VP.n0 VP.t3 73.9649
R65 VP.n17 VP.t2 73.9649
R66 VP.n55 VP.t7 73.9649
R67 VP.n42 VP.t0 73.9649
R68 VP.n30 VP.t4 73.9649
R69 VP.n31 VP.n30 64.7311
R70 VP.n72 VP.n70 58.0637
R71 VP.n77 VP.n14 56.5193
R72 VP.n90 VP.n10 56.5193
R73 VP.n103 VP.n6 56.5193
R74 VP.n116 VP.n2 56.5193
R75 VP.n62 VP.n19 56.5193
R76 VP.n49 VP.n23 56.5193
R77 VP.n36 VP.n27 56.5193
R78 VP.n75 VP.n16 24.4675
R79 VP.n76 VP.n75 24.4675
R80 VP.n77 VP.n76 24.4675
R81 VP.n81 VP.n14 24.4675
R82 VP.n82 VP.n81 24.4675
R83 VP.n84 VP.n82 24.4675
R84 VP.n88 VP.n12 24.4675
R85 VP.n89 VP.n88 24.4675
R86 VP.n90 VP.n89 24.4675
R87 VP.n94 VP.n10 24.4675
R88 VP.n95 VP.n94 24.4675
R89 VP.n97 VP.n95 24.4675
R90 VP.n101 VP.n8 24.4675
R91 VP.n102 VP.n101 24.4675
R92 VP.n103 VP.n102 24.4675
R93 VP.n107 VP.n6 24.4675
R94 VP.n108 VP.n107 24.4675
R95 VP.n110 VP.n108 24.4675
R96 VP.n114 VP.n4 24.4675
R97 VP.n115 VP.n114 24.4675
R98 VP.n116 VP.n115 24.4675
R99 VP.n120 VP.n2 24.4675
R100 VP.n121 VP.n120 24.4675
R101 VP.n122 VP.n121 24.4675
R102 VP.n66 VP.n19 24.4675
R103 VP.n67 VP.n66 24.4675
R104 VP.n68 VP.n67 24.4675
R105 VP.n53 VP.n23 24.4675
R106 VP.n54 VP.n53 24.4675
R107 VP.n56 VP.n54 24.4675
R108 VP.n60 VP.n21 24.4675
R109 VP.n61 VP.n60 24.4675
R110 VP.n62 VP.n61 24.4675
R111 VP.n40 VP.n27 24.4675
R112 VP.n41 VP.n40 24.4675
R113 VP.n43 VP.n41 24.4675
R114 VP.n47 VP.n25 24.4675
R115 VP.n48 VP.n47 24.4675
R116 VP.n49 VP.n48 24.4675
R117 VP.n34 VP.n29 24.4675
R118 VP.n35 VP.n34 24.4675
R119 VP.n36 VP.n35 24.4675
R120 VP.n84 VP.n83 14.6807
R121 VP.n109 VP.n4 14.6807
R122 VP.n55 VP.n21 14.6807
R123 VP.n97 VP.n96 12.234
R124 VP.n96 VP.n8 12.234
R125 VP.n43 VP.n42 12.234
R126 VP.n42 VP.n25 12.234
R127 VP.n83 VP.n12 9.7873
R128 VP.n110 VP.n109 9.7873
R129 VP.n56 VP.n55 9.7873
R130 VP.n30 VP.n29 9.7873
R131 VP.n71 VP.n16 7.3406
R132 VP.n122 VP.n0 7.3406
R133 VP.n68 VP.n17 7.3406
R134 VP.n32 VP.n31 3.24374
R135 VP.n70 VP.n69 0.354971
R136 VP.n73 VP.n72 0.354971
R137 VP.n124 VP.n123 0.354971
R138 VP VP.n124 0.26696
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VTAIL.n11 VTAIL.t6 48.67
R194 VTAIL.n17 VTAIL.t0 48.6699
R195 VTAIL.n2 VTAIL.t11 48.6699
R196 VTAIL.n16 VTAIL.t16 48.6699
R197 VTAIL.n15 VTAIL.n14 46.8879
R198 VTAIL.n13 VTAIL.n12 46.8879
R199 VTAIL.n10 VTAIL.n9 46.8879
R200 VTAIL.n8 VTAIL.n7 46.8879
R201 VTAIL.n19 VTAIL.n18 46.8877
R202 VTAIL.n1 VTAIL.n0 46.8877
R203 VTAIL.n4 VTAIL.n3 46.8877
R204 VTAIL.n6 VTAIL.n5 46.8877
R205 VTAIL.n8 VTAIL.n6 28.7548
R206 VTAIL.n17 VTAIL.n16 25.3496
R207 VTAIL.n10 VTAIL.n8 3.40567
R208 VTAIL.n11 VTAIL.n10 3.40567
R209 VTAIL.n15 VTAIL.n13 3.40567
R210 VTAIL.n16 VTAIL.n15 3.40567
R211 VTAIL.n6 VTAIL.n4 3.40567
R212 VTAIL.n4 VTAIL.n2 3.40567
R213 VTAIL.n19 VTAIL.n17 3.40567
R214 VTAIL VTAIL.n1 2.61257
R215 VTAIL.n13 VTAIL.n11 2.17291
R216 VTAIL.n2 VTAIL.n1 2.17291
R217 VTAIL.n18 VTAIL.t3 1.78268
R218 VTAIL.n18 VTAIL.t8 1.78268
R219 VTAIL.n0 VTAIL.t4 1.78268
R220 VTAIL.n0 VTAIL.t2 1.78268
R221 VTAIL.n3 VTAIL.t18 1.78268
R222 VTAIL.n3 VTAIL.t10 1.78268
R223 VTAIL.n5 VTAIL.t14 1.78268
R224 VTAIL.n5 VTAIL.t13 1.78268
R225 VTAIL.n14 VTAIL.t17 1.78268
R226 VTAIL.n14 VTAIL.t15 1.78268
R227 VTAIL.n12 VTAIL.t12 1.78268
R228 VTAIL.n12 VTAIL.t9 1.78268
R229 VTAIL.n9 VTAIL.t1 1.78268
R230 VTAIL.n9 VTAIL.t7 1.78268
R231 VTAIL.n7 VTAIL.t19 1.78268
R232 VTAIL.n7 VTAIL.t5 1.78268
R233 VTAIL VTAIL.n19 0.793603
R234 VDD1.n1 VDD1.t3 68.754
R235 VDD1.n3 VDD1.t0 68.7539
R236 VDD1.n5 VDD1.n4 66.065
R237 VDD1.n1 VDD1.n0 63.5667
R238 VDD1.n7 VDD1.n6 63.5665
R239 VDD1.n3 VDD1.n2 63.5665
R240 VDD1.n7 VDD1.n5 51.753
R241 VDD1 VDD1.n7 2.49619
R242 VDD1.n6 VDD1.t2 1.78268
R243 VDD1.n6 VDD1.t7 1.78268
R244 VDD1.n0 VDD1.t5 1.78268
R245 VDD1.n0 VDD1.t9 1.78268
R246 VDD1.n4 VDD1.t1 1.78268
R247 VDD1.n4 VDD1.t6 1.78268
R248 VDD1.n2 VDD1.t4 1.78268
R249 VDD1.n2 VDD1.t8 1.78268
R250 VDD1 VDD1.n1 0.909983
R251 VDD1.n5 VDD1.n3 0.796447
R252 B.n903 B.n902 585
R253 B.n905 B.n190 585
R254 B.n908 B.n907 585
R255 B.n909 B.n189 585
R256 B.n911 B.n910 585
R257 B.n913 B.n188 585
R258 B.n916 B.n915 585
R259 B.n917 B.n187 585
R260 B.n919 B.n918 585
R261 B.n921 B.n186 585
R262 B.n924 B.n923 585
R263 B.n925 B.n185 585
R264 B.n927 B.n926 585
R265 B.n929 B.n184 585
R266 B.n932 B.n931 585
R267 B.n933 B.n183 585
R268 B.n935 B.n934 585
R269 B.n937 B.n182 585
R270 B.n940 B.n939 585
R271 B.n941 B.n181 585
R272 B.n943 B.n942 585
R273 B.n945 B.n180 585
R274 B.n948 B.n947 585
R275 B.n949 B.n179 585
R276 B.n951 B.n950 585
R277 B.n953 B.n178 585
R278 B.n956 B.n955 585
R279 B.n957 B.n177 585
R280 B.n959 B.n958 585
R281 B.n961 B.n176 585
R282 B.n964 B.n963 585
R283 B.n965 B.n175 585
R284 B.n967 B.n966 585
R285 B.n969 B.n174 585
R286 B.n972 B.n971 585
R287 B.n973 B.n173 585
R288 B.n975 B.n974 585
R289 B.n977 B.n172 585
R290 B.n980 B.n979 585
R291 B.n982 B.n169 585
R292 B.n984 B.n983 585
R293 B.n986 B.n168 585
R294 B.n989 B.n988 585
R295 B.n990 B.n167 585
R296 B.n992 B.n991 585
R297 B.n994 B.n166 585
R298 B.n997 B.n996 585
R299 B.n998 B.n162 585
R300 B.n1000 B.n999 585
R301 B.n1002 B.n161 585
R302 B.n1005 B.n1004 585
R303 B.n1006 B.n160 585
R304 B.n1008 B.n1007 585
R305 B.n1010 B.n159 585
R306 B.n1013 B.n1012 585
R307 B.n1014 B.n158 585
R308 B.n1016 B.n1015 585
R309 B.n1018 B.n157 585
R310 B.n1021 B.n1020 585
R311 B.n1022 B.n156 585
R312 B.n1024 B.n1023 585
R313 B.n1026 B.n155 585
R314 B.n1029 B.n1028 585
R315 B.n1030 B.n154 585
R316 B.n1032 B.n1031 585
R317 B.n1034 B.n153 585
R318 B.n1037 B.n1036 585
R319 B.n1038 B.n152 585
R320 B.n1040 B.n1039 585
R321 B.n1042 B.n151 585
R322 B.n1045 B.n1044 585
R323 B.n1046 B.n150 585
R324 B.n1048 B.n1047 585
R325 B.n1050 B.n149 585
R326 B.n1053 B.n1052 585
R327 B.n1054 B.n148 585
R328 B.n1056 B.n1055 585
R329 B.n1058 B.n147 585
R330 B.n1061 B.n1060 585
R331 B.n1062 B.n146 585
R332 B.n1064 B.n1063 585
R333 B.n1066 B.n145 585
R334 B.n1069 B.n1068 585
R335 B.n1070 B.n144 585
R336 B.n1072 B.n1071 585
R337 B.n1074 B.n143 585
R338 B.n1077 B.n1076 585
R339 B.n1078 B.n142 585
R340 B.n901 B.n140 585
R341 B.n1081 B.n140 585
R342 B.n900 B.n139 585
R343 B.n1082 B.n139 585
R344 B.n899 B.n138 585
R345 B.n1083 B.n138 585
R346 B.n898 B.n897 585
R347 B.n897 B.n134 585
R348 B.n896 B.n133 585
R349 B.n1089 B.n133 585
R350 B.n895 B.n132 585
R351 B.n1090 B.n132 585
R352 B.n894 B.n131 585
R353 B.n1091 B.n131 585
R354 B.n893 B.n892 585
R355 B.n892 B.n127 585
R356 B.n891 B.n126 585
R357 B.n1097 B.n126 585
R358 B.n890 B.n125 585
R359 B.n1098 B.n125 585
R360 B.n889 B.n124 585
R361 B.n1099 B.n124 585
R362 B.n888 B.n887 585
R363 B.n887 B.n120 585
R364 B.n886 B.n119 585
R365 B.n1105 B.n119 585
R366 B.n885 B.n118 585
R367 B.n1106 B.n118 585
R368 B.n884 B.n117 585
R369 B.n1107 B.n117 585
R370 B.n883 B.n882 585
R371 B.n882 B.n113 585
R372 B.n881 B.n112 585
R373 B.n1113 B.n112 585
R374 B.n880 B.n111 585
R375 B.n1114 B.n111 585
R376 B.n879 B.n110 585
R377 B.n1115 B.n110 585
R378 B.n878 B.n877 585
R379 B.n877 B.n106 585
R380 B.n876 B.n105 585
R381 B.n1121 B.n105 585
R382 B.n875 B.n104 585
R383 B.n1122 B.n104 585
R384 B.n874 B.n103 585
R385 B.n1123 B.n103 585
R386 B.n873 B.n872 585
R387 B.n872 B.n99 585
R388 B.n871 B.n98 585
R389 B.n1129 B.n98 585
R390 B.n870 B.n97 585
R391 B.n1130 B.n97 585
R392 B.n869 B.n96 585
R393 B.n1131 B.n96 585
R394 B.n868 B.n867 585
R395 B.n867 B.n92 585
R396 B.n866 B.n91 585
R397 B.n1137 B.n91 585
R398 B.n865 B.n90 585
R399 B.n1138 B.n90 585
R400 B.n864 B.n89 585
R401 B.n1139 B.n89 585
R402 B.n863 B.n862 585
R403 B.n862 B.n85 585
R404 B.n861 B.n84 585
R405 B.n1145 B.n84 585
R406 B.n860 B.n83 585
R407 B.n1146 B.n83 585
R408 B.n859 B.n82 585
R409 B.n1147 B.n82 585
R410 B.n858 B.n857 585
R411 B.n857 B.n81 585
R412 B.n856 B.n77 585
R413 B.n1153 B.n77 585
R414 B.n855 B.n76 585
R415 B.n1154 B.n76 585
R416 B.n854 B.n75 585
R417 B.n1155 B.n75 585
R418 B.n853 B.n852 585
R419 B.n852 B.n71 585
R420 B.n851 B.n70 585
R421 B.n1161 B.n70 585
R422 B.n850 B.n69 585
R423 B.n1162 B.n69 585
R424 B.n849 B.n68 585
R425 B.n1163 B.n68 585
R426 B.n848 B.n847 585
R427 B.n847 B.n64 585
R428 B.n846 B.n63 585
R429 B.n1169 B.n63 585
R430 B.n845 B.n62 585
R431 B.n1170 B.n62 585
R432 B.n844 B.n61 585
R433 B.n1171 B.n61 585
R434 B.n843 B.n842 585
R435 B.n842 B.n60 585
R436 B.n841 B.n56 585
R437 B.n1177 B.n56 585
R438 B.n840 B.n55 585
R439 B.n1178 B.n55 585
R440 B.n839 B.n54 585
R441 B.n1179 B.n54 585
R442 B.n838 B.n837 585
R443 B.n837 B.n50 585
R444 B.n836 B.n49 585
R445 B.n1185 B.n49 585
R446 B.n835 B.n48 585
R447 B.n1186 B.n48 585
R448 B.n834 B.n47 585
R449 B.n1187 B.n47 585
R450 B.n833 B.n832 585
R451 B.n832 B.n43 585
R452 B.n831 B.n42 585
R453 B.n1193 B.n42 585
R454 B.n830 B.n41 585
R455 B.n1194 B.n41 585
R456 B.n829 B.n40 585
R457 B.n1195 B.n40 585
R458 B.n828 B.n827 585
R459 B.n827 B.n36 585
R460 B.n826 B.n35 585
R461 B.n1201 B.n35 585
R462 B.n825 B.n34 585
R463 B.n1202 B.n34 585
R464 B.n824 B.n33 585
R465 B.n1203 B.n33 585
R466 B.n823 B.n822 585
R467 B.n822 B.n29 585
R468 B.n821 B.n28 585
R469 B.n1209 B.n28 585
R470 B.n820 B.n27 585
R471 B.n1210 B.n27 585
R472 B.n819 B.n26 585
R473 B.n1211 B.n26 585
R474 B.n818 B.n817 585
R475 B.n817 B.n22 585
R476 B.n816 B.n21 585
R477 B.n1217 B.n21 585
R478 B.n815 B.n20 585
R479 B.n1218 B.n20 585
R480 B.n814 B.n19 585
R481 B.n1219 B.n19 585
R482 B.n813 B.n812 585
R483 B.n812 B.n15 585
R484 B.n811 B.n14 585
R485 B.n1225 B.n14 585
R486 B.n810 B.n13 585
R487 B.n1226 B.n13 585
R488 B.n809 B.n12 585
R489 B.n1227 B.n12 585
R490 B.n808 B.n807 585
R491 B.n807 B.n8 585
R492 B.n806 B.n7 585
R493 B.n1233 B.n7 585
R494 B.n805 B.n6 585
R495 B.n1234 B.n6 585
R496 B.n804 B.n5 585
R497 B.n1235 B.n5 585
R498 B.n803 B.n802 585
R499 B.n802 B.n4 585
R500 B.n801 B.n191 585
R501 B.n801 B.n800 585
R502 B.n791 B.n192 585
R503 B.n193 B.n192 585
R504 B.n793 B.n792 585
R505 B.n794 B.n793 585
R506 B.n790 B.n198 585
R507 B.n198 B.n197 585
R508 B.n789 B.n788 585
R509 B.n788 B.n787 585
R510 B.n200 B.n199 585
R511 B.n201 B.n200 585
R512 B.n780 B.n779 585
R513 B.n781 B.n780 585
R514 B.n778 B.n206 585
R515 B.n206 B.n205 585
R516 B.n777 B.n776 585
R517 B.n776 B.n775 585
R518 B.n208 B.n207 585
R519 B.n209 B.n208 585
R520 B.n768 B.n767 585
R521 B.n769 B.n768 585
R522 B.n766 B.n214 585
R523 B.n214 B.n213 585
R524 B.n765 B.n764 585
R525 B.n764 B.n763 585
R526 B.n216 B.n215 585
R527 B.n217 B.n216 585
R528 B.n756 B.n755 585
R529 B.n757 B.n756 585
R530 B.n754 B.n222 585
R531 B.n222 B.n221 585
R532 B.n753 B.n752 585
R533 B.n752 B.n751 585
R534 B.n224 B.n223 585
R535 B.n225 B.n224 585
R536 B.n744 B.n743 585
R537 B.n745 B.n744 585
R538 B.n742 B.n230 585
R539 B.n230 B.n229 585
R540 B.n741 B.n740 585
R541 B.n740 B.n739 585
R542 B.n232 B.n231 585
R543 B.n233 B.n232 585
R544 B.n732 B.n731 585
R545 B.n733 B.n732 585
R546 B.n730 B.n238 585
R547 B.n238 B.n237 585
R548 B.n729 B.n728 585
R549 B.n728 B.n727 585
R550 B.n240 B.n239 585
R551 B.n241 B.n240 585
R552 B.n720 B.n719 585
R553 B.n721 B.n720 585
R554 B.n718 B.n246 585
R555 B.n246 B.n245 585
R556 B.n717 B.n716 585
R557 B.n716 B.n715 585
R558 B.n248 B.n247 585
R559 B.n708 B.n248 585
R560 B.n707 B.n706 585
R561 B.n709 B.n707 585
R562 B.n705 B.n253 585
R563 B.n253 B.n252 585
R564 B.n704 B.n703 585
R565 B.n703 B.n702 585
R566 B.n255 B.n254 585
R567 B.n256 B.n255 585
R568 B.n695 B.n694 585
R569 B.n696 B.n695 585
R570 B.n693 B.n261 585
R571 B.n261 B.n260 585
R572 B.n692 B.n691 585
R573 B.n691 B.n690 585
R574 B.n263 B.n262 585
R575 B.n264 B.n263 585
R576 B.n683 B.n682 585
R577 B.n684 B.n683 585
R578 B.n681 B.n269 585
R579 B.n269 B.n268 585
R580 B.n680 B.n679 585
R581 B.n679 B.n678 585
R582 B.n271 B.n270 585
R583 B.n671 B.n271 585
R584 B.n670 B.n669 585
R585 B.n672 B.n670 585
R586 B.n668 B.n276 585
R587 B.n276 B.n275 585
R588 B.n667 B.n666 585
R589 B.n666 B.n665 585
R590 B.n278 B.n277 585
R591 B.n279 B.n278 585
R592 B.n658 B.n657 585
R593 B.n659 B.n658 585
R594 B.n656 B.n284 585
R595 B.n284 B.n283 585
R596 B.n655 B.n654 585
R597 B.n654 B.n653 585
R598 B.n286 B.n285 585
R599 B.n287 B.n286 585
R600 B.n646 B.n645 585
R601 B.n647 B.n646 585
R602 B.n644 B.n292 585
R603 B.n292 B.n291 585
R604 B.n643 B.n642 585
R605 B.n642 B.n641 585
R606 B.n294 B.n293 585
R607 B.n295 B.n294 585
R608 B.n634 B.n633 585
R609 B.n635 B.n634 585
R610 B.n632 B.n300 585
R611 B.n300 B.n299 585
R612 B.n631 B.n630 585
R613 B.n630 B.n629 585
R614 B.n302 B.n301 585
R615 B.n303 B.n302 585
R616 B.n622 B.n621 585
R617 B.n623 B.n622 585
R618 B.n620 B.n308 585
R619 B.n308 B.n307 585
R620 B.n619 B.n618 585
R621 B.n618 B.n617 585
R622 B.n310 B.n309 585
R623 B.n311 B.n310 585
R624 B.n610 B.n609 585
R625 B.n611 B.n610 585
R626 B.n608 B.n316 585
R627 B.n316 B.n315 585
R628 B.n607 B.n606 585
R629 B.n606 B.n605 585
R630 B.n318 B.n317 585
R631 B.n319 B.n318 585
R632 B.n598 B.n597 585
R633 B.n599 B.n598 585
R634 B.n596 B.n323 585
R635 B.n327 B.n323 585
R636 B.n595 B.n594 585
R637 B.n594 B.n593 585
R638 B.n325 B.n324 585
R639 B.n326 B.n325 585
R640 B.n586 B.n585 585
R641 B.n587 B.n586 585
R642 B.n584 B.n332 585
R643 B.n332 B.n331 585
R644 B.n583 B.n582 585
R645 B.n582 B.n581 585
R646 B.n334 B.n333 585
R647 B.n335 B.n334 585
R648 B.n574 B.n573 585
R649 B.n575 B.n574 585
R650 B.n572 B.n340 585
R651 B.n340 B.n339 585
R652 B.n571 B.n570 585
R653 B.n570 B.n569 585
R654 B.n566 B.n344 585
R655 B.n565 B.n564 585
R656 B.n562 B.n345 585
R657 B.n562 B.n343 585
R658 B.n561 B.n560 585
R659 B.n559 B.n558 585
R660 B.n557 B.n347 585
R661 B.n555 B.n554 585
R662 B.n553 B.n348 585
R663 B.n552 B.n551 585
R664 B.n549 B.n349 585
R665 B.n547 B.n546 585
R666 B.n545 B.n350 585
R667 B.n544 B.n543 585
R668 B.n541 B.n351 585
R669 B.n539 B.n538 585
R670 B.n537 B.n352 585
R671 B.n536 B.n535 585
R672 B.n533 B.n353 585
R673 B.n531 B.n530 585
R674 B.n529 B.n354 585
R675 B.n528 B.n527 585
R676 B.n525 B.n355 585
R677 B.n523 B.n522 585
R678 B.n521 B.n356 585
R679 B.n520 B.n519 585
R680 B.n517 B.n357 585
R681 B.n515 B.n514 585
R682 B.n513 B.n358 585
R683 B.n512 B.n511 585
R684 B.n509 B.n359 585
R685 B.n507 B.n506 585
R686 B.n505 B.n360 585
R687 B.n504 B.n503 585
R688 B.n501 B.n361 585
R689 B.n499 B.n498 585
R690 B.n497 B.n362 585
R691 B.n496 B.n495 585
R692 B.n493 B.n363 585
R693 B.n491 B.n490 585
R694 B.n488 B.n364 585
R695 B.n487 B.n486 585
R696 B.n484 B.n367 585
R697 B.n482 B.n481 585
R698 B.n480 B.n368 585
R699 B.n479 B.n478 585
R700 B.n476 B.n369 585
R701 B.n474 B.n473 585
R702 B.n472 B.n370 585
R703 B.n471 B.n470 585
R704 B.n468 B.n467 585
R705 B.n466 B.n465 585
R706 B.n464 B.n375 585
R707 B.n462 B.n461 585
R708 B.n460 B.n376 585
R709 B.n459 B.n458 585
R710 B.n456 B.n377 585
R711 B.n454 B.n453 585
R712 B.n452 B.n378 585
R713 B.n451 B.n450 585
R714 B.n448 B.n379 585
R715 B.n446 B.n445 585
R716 B.n444 B.n380 585
R717 B.n443 B.n442 585
R718 B.n440 B.n381 585
R719 B.n438 B.n437 585
R720 B.n436 B.n382 585
R721 B.n435 B.n434 585
R722 B.n432 B.n383 585
R723 B.n430 B.n429 585
R724 B.n428 B.n384 585
R725 B.n427 B.n426 585
R726 B.n424 B.n385 585
R727 B.n422 B.n421 585
R728 B.n420 B.n386 585
R729 B.n419 B.n418 585
R730 B.n416 B.n387 585
R731 B.n414 B.n413 585
R732 B.n412 B.n388 585
R733 B.n411 B.n410 585
R734 B.n408 B.n389 585
R735 B.n406 B.n405 585
R736 B.n404 B.n390 585
R737 B.n403 B.n402 585
R738 B.n400 B.n391 585
R739 B.n398 B.n397 585
R740 B.n396 B.n392 585
R741 B.n395 B.n394 585
R742 B.n342 B.n341 585
R743 B.n343 B.n342 585
R744 B.n568 B.n567 585
R745 B.n569 B.n568 585
R746 B.n338 B.n337 585
R747 B.n339 B.n338 585
R748 B.n577 B.n576 585
R749 B.n576 B.n575 585
R750 B.n578 B.n336 585
R751 B.n336 B.n335 585
R752 B.n580 B.n579 585
R753 B.n581 B.n580 585
R754 B.n330 B.n329 585
R755 B.n331 B.n330 585
R756 B.n589 B.n588 585
R757 B.n588 B.n587 585
R758 B.n590 B.n328 585
R759 B.n328 B.n326 585
R760 B.n592 B.n591 585
R761 B.n593 B.n592 585
R762 B.n322 B.n321 585
R763 B.n327 B.n322 585
R764 B.n601 B.n600 585
R765 B.n600 B.n599 585
R766 B.n602 B.n320 585
R767 B.n320 B.n319 585
R768 B.n604 B.n603 585
R769 B.n605 B.n604 585
R770 B.n314 B.n313 585
R771 B.n315 B.n314 585
R772 B.n613 B.n612 585
R773 B.n612 B.n611 585
R774 B.n614 B.n312 585
R775 B.n312 B.n311 585
R776 B.n616 B.n615 585
R777 B.n617 B.n616 585
R778 B.n306 B.n305 585
R779 B.n307 B.n306 585
R780 B.n625 B.n624 585
R781 B.n624 B.n623 585
R782 B.n626 B.n304 585
R783 B.n304 B.n303 585
R784 B.n628 B.n627 585
R785 B.n629 B.n628 585
R786 B.n298 B.n297 585
R787 B.n299 B.n298 585
R788 B.n637 B.n636 585
R789 B.n636 B.n635 585
R790 B.n638 B.n296 585
R791 B.n296 B.n295 585
R792 B.n640 B.n639 585
R793 B.n641 B.n640 585
R794 B.n290 B.n289 585
R795 B.n291 B.n290 585
R796 B.n649 B.n648 585
R797 B.n648 B.n647 585
R798 B.n650 B.n288 585
R799 B.n288 B.n287 585
R800 B.n652 B.n651 585
R801 B.n653 B.n652 585
R802 B.n282 B.n281 585
R803 B.n283 B.n282 585
R804 B.n661 B.n660 585
R805 B.n660 B.n659 585
R806 B.n662 B.n280 585
R807 B.n280 B.n279 585
R808 B.n664 B.n663 585
R809 B.n665 B.n664 585
R810 B.n274 B.n273 585
R811 B.n275 B.n274 585
R812 B.n674 B.n673 585
R813 B.n673 B.n672 585
R814 B.n675 B.n272 585
R815 B.n671 B.n272 585
R816 B.n677 B.n676 585
R817 B.n678 B.n677 585
R818 B.n267 B.n266 585
R819 B.n268 B.n267 585
R820 B.n686 B.n685 585
R821 B.n685 B.n684 585
R822 B.n687 B.n265 585
R823 B.n265 B.n264 585
R824 B.n689 B.n688 585
R825 B.n690 B.n689 585
R826 B.n259 B.n258 585
R827 B.n260 B.n259 585
R828 B.n698 B.n697 585
R829 B.n697 B.n696 585
R830 B.n699 B.n257 585
R831 B.n257 B.n256 585
R832 B.n701 B.n700 585
R833 B.n702 B.n701 585
R834 B.n251 B.n250 585
R835 B.n252 B.n251 585
R836 B.n711 B.n710 585
R837 B.n710 B.n709 585
R838 B.n712 B.n249 585
R839 B.n708 B.n249 585
R840 B.n714 B.n713 585
R841 B.n715 B.n714 585
R842 B.n244 B.n243 585
R843 B.n245 B.n244 585
R844 B.n723 B.n722 585
R845 B.n722 B.n721 585
R846 B.n724 B.n242 585
R847 B.n242 B.n241 585
R848 B.n726 B.n725 585
R849 B.n727 B.n726 585
R850 B.n236 B.n235 585
R851 B.n237 B.n236 585
R852 B.n735 B.n734 585
R853 B.n734 B.n733 585
R854 B.n736 B.n234 585
R855 B.n234 B.n233 585
R856 B.n738 B.n737 585
R857 B.n739 B.n738 585
R858 B.n228 B.n227 585
R859 B.n229 B.n228 585
R860 B.n747 B.n746 585
R861 B.n746 B.n745 585
R862 B.n748 B.n226 585
R863 B.n226 B.n225 585
R864 B.n750 B.n749 585
R865 B.n751 B.n750 585
R866 B.n220 B.n219 585
R867 B.n221 B.n220 585
R868 B.n759 B.n758 585
R869 B.n758 B.n757 585
R870 B.n760 B.n218 585
R871 B.n218 B.n217 585
R872 B.n762 B.n761 585
R873 B.n763 B.n762 585
R874 B.n212 B.n211 585
R875 B.n213 B.n212 585
R876 B.n771 B.n770 585
R877 B.n770 B.n769 585
R878 B.n772 B.n210 585
R879 B.n210 B.n209 585
R880 B.n774 B.n773 585
R881 B.n775 B.n774 585
R882 B.n204 B.n203 585
R883 B.n205 B.n204 585
R884 B.n783 B.n782 585
R885 B.n782 B.n781 585
R886 B.n784 B.n202 585
R887 B.n202 B.n201 585
R888 B.n786 B.n785 585
R889 B.n787 B.n786 585
R890 B.n196 B.n195 585
R891 B.n197 B.n196 585
R892 B.n796 B.n795 585
R893 B.n795 B.n794 585
R894 B.n797 B.n194 585
R895 B.n194 B.n193 585
R896 B.n799 B.n798 585
R897 B.n800 B.n799 585
R898 B.n2 B.n0 585
R899 B.n4 B.n2 585
R900 B.n3 B.n1 585
R901 B.n1234 B.n3 585
R902 B.n1232 B.n1231 585
R903 B.n1233 B.n1232 585
R904 B.n1230 B.n9 585
R905 B.n9 B.n8 585
R906 B.n1229 B.n1228 585
R907 B.n1228 B.n1227 585
R908 B.n11 B.n10 585
R909 B.n1226 B.n11 585
R910 B.n1224 B.n1223 585
R911 B.n1225 B.n1224 585
R912 B.n1222 B.n16 585
R913 B.n16 B.n15 585
R914 B.n1221 B.n1220 585
R915 B.n1220 B.n1219 585
R916 B.n18 B.n17 585
R917 B.n1218 B.n18 585
R918 B.n1216 B.n1215 585
R919 B.n1217 B.n1216 585
R920 B.n1214 B.n23 585
R921 B.n23 B.n22 585
R922 B.n1213 B.n1212 585
R923 B.n1212 B.n1211 585
R924 B.n25 B.n24 585
R925 B.n1210 B.n25 585
R926 B.n1208 B.n1207 585
R927 B.n1209 B.n1208 585
R928 B.n1206 B.n30 585
R929 B.n30 B.n29 585
R930 B.n1205 B.n1204 585
R931 B.n1204 B.n1203 585
R932 B.n32 B.n31 585
R933 B.n1202 B.n32 585
R934 B.n1200 B.n1199 585
R935 B.n1201 B.n1200 585
R936 B.n1198 B.n37 585
R937 B.n37 B.n36 585
R938 B.n1197 B.n1196 585
R939 B.n1196 B.n1195 585
R940 B.n39 B.n38 585
R941 B.n1194 B.n39 585
R942 B.n1192 B.n1191 585
R943 B.n1193 B.n1192 585
R944 B.n1190 B.n44 585
R945 B.n44 B.n43 585
R946 B.n1189 B.n1188 585
R947 B.n1188 B.n1187 585
R948 B.n46 B.n45 585
R949 B.n1186 B.n46 585
R950 B.n1184 B.n1183 585
R951 B.n1185 B.n1184 585
R952 B.n1182 B.n51 585
R953 B.n51 B.n50 585
R954 B.n1181 B.n1180 585
R955 B.n1180 B.n1179 585
R956 B.n53 B.n52 585
R957 B.n1178 B.n53 585
R958 B.n1176 B.n1175 585
R959 B.n1177 B.n1176 585
R960 B.n1174 B.n57 585
R961 B.n60 B.n57 585
R962 B.n1173 B.n1172 585
R963 B.n1172 B.n1171 585
R964 B.n59 B.n58 585
R965 B.n1170 B.n59 585
R966 B.n1168 B.n1167 585
R967 B.n1169 B.n1168 585
R968 B.n1166 B.n65 585
R969 B.n65 B.n64 585
R970 B.n1165 B.n1164 585
R971 B.n1164 B.n1163 585
R972 B.n67 B.n66 585
R973 B.n1162 B.n67 585
R974 B.n1160 B.n1159 585
R975 B.n1161 B.n1160 585
R976 B.n1158 B.n72 585
R977 B.n72 B.n71 585
R978 B.n1157 B.n1156 585
R979 B.n1156 B.n1155 585
R980 B.n74 B.n73 585
R981 B.n1154 B.n74 585
R982 B.n1152 B.n1151 585
R983 B.n1153 B.n1152 585
R984 B.n1150 B.n78 585
R985 B.n81 B.n78 585
R986 B.n1149 B.n1148 585
R987 B.n1148 B.n1147 585
R988 B.n80 B.n79 585
R989 B.n1146 B.n80 585
R990 B.n1144 B.n1143 585
R991 B.n1145 B.n1144 585
R992 B.n1142 B.n86 585
R993 B.n86 B.n85 585
R994 B.n1141 B.n1140 585
R995 B.n1140 B.n1139 585
R996 B.n88 B.n87 585
R997 B.n1138 B.n88 585
R998 B.n1136 B.n1135 585
R999 B.n1137 B.n1136 585
R1000 B.n1134 B.n93 585
R1001 B.n93 B.n92 585
R1002 B.n1133 B.n1132 585
R1003 B.n1132 B.n1131 585
R1004 B.n95 B.n94 585
R1005 B.n1130 B.n95 585
R1006 B.n1128 B.n1127 585
R1007 B.n1129 B.n1128 585
R1008 B.n1126 B.n100 585
R1009 B.n100 B.n99 585
R1010 B.n1125 B.n1124 585
R1011 B.n1124 B.n1123 585
R1012 B.n102 B.n101 585
R1013 B.n1122 B.n102 585
R1014 B.n1120 B.n1119 585
R1015 B.n1121 B.n1120 585
R1016 B.n1118 B.n107 585
R1017 B.n107 B.n106 585
R1018 B.n1117 B.n1116 585
R1019 B.n1116 B.n1115 585
R1020 B.n109 B.n108 585
R1021 B.n1114 B.n109 585
R1022 B.n1112 B.n1111 585
R1023 B.n1113 B.n1112 585
R1024 B.n1110 B.n114 585
R1025 B.n114 B.n113 585
R1026 B.n1109 B.n1108 585
R1027 B.n1108 B.n1107 585
R1028 B.n116 B.n115 585
R1029 B.n1106 B.n116 585
R1030 B.n1104 B.n1103 585
R1031 B.n1105 B.n1104 585
R1032 B.n1102 B.n121 585
R1033 B.n121 B.n120 585
R1034 B.n1101 B.n1100 585
R1035 B.n1100 B.n1099 585
R1036 B.n123 B.n122 585
R1037 B.n1098 B.n123 585
R1038 B.n1096 B.n1095 585
R1039 B.n1097 B.n1096 585
R1040 B.n1094 B.n128 585
R1041 B.n128 B.n127 585
R1042 B.n1093 B.n1092 585
R1043 B.n1092 B.n1091 585
R1044 B.n130 B.n129 585
R1045 B.n1090 B.n130 585
R1046 B.n1088 B.n1087 585
R1047 B.n1089 B.n1088 585
R1048 B.n1086 B.n135 585
R1049 B.n135 B.n134 585
R1050 B.n1085 B.n1084 585
R1051 B.n1084 B.n1083 585
R1052 B.n137 B.n136 585
R1053 B.n1082 B.n137 585
R1054 B.n1080 B.n1079 585
R1055 B.n1081 B.n1080 585
R1056 B.n1237 B.n1236 585
R1057 B.n1236 B.n1235 585
R1058 B.n568 B.n344 434.841
R1059 B.n1080 B.n142 434.841
R1060 B.n570 B.n342 434.841
R1061 B.n903 B.n140 434.841
R1062 B.n371 B.t20 283.163
R1063 B.n365 B.t9 283.163
R1064 B.n163 B.t13 283.163
R1065 B.n170 B.t17 283.163
R1066 B.n904 B.n141 256.663
R1067 B.n906 B.n141 256.663
R1068 B.n912 B.n141 256.663
R1069 B.n914 B.n141 256.663
R1070 B.n920 B.n141 256.663
R1071 B.n922 B.n141 256.663
R1072 B.n928 B.n141 256.663
R1073 B.n930 B.n141 256.663
R1074 B.n936 B.n141 256.663
R1075 B.n938 B.n141 256.663
R1076 B.n944 B.n141 256.663
R1077 B.n946 B.n141 256.663
R1078 B.n952 B.n141 256.663
R1079 B.n954 B.n141 256.663
R1080 B.n960 B.n141 256.663
R1081 B.n962 B.n141 256.663
R1082 B.n968 B.n141 256.663
R1083 B.n970 B.n141 256.663
R1084 B.n976 B.n141 256.663
R1085 B.n978 B.n141 256.663
R1086 B.n985 B.n141 256.663
R1087 B.n987 B.n141 256.663
R1088 B.n993 B.n141 256.663
R1089 B.n995 B.n141 256.663
R1090 B.n1001 B.n141 256.663
R1091 B.n1003 B.n141 256.663
R1092 B.n1009 B.n141 256.663
R1093 B.n1011 B.n141 256.663
R1094 B.n1017 B.n141 256.663
R1095 B.n1019 B.n141 256.663
R1096 B.n1025 B.n141 256.663
R1097 B.n1027 B.n141 256.663
R1098 B.n1033 B.n141 256.663
R1099 B.n1035 B.n141 256.663
R1100 B.n1041 B.n141 256.663
R1101 B.n1043 B.n141 256.663
R1102 B.n1049 B.n141 256.663
R1103 B.n1051 B.n141 256.663
R1104 B.n1057 B.n141 256.663
R1105 B.n1059 B.n141 256.663
R1106 B.n1065 B.n141 256.663
R1107 B.n1067 B.n141 256.663
R1108 B.n1073 B.n141 256.663
R1109 B.n1075 B.n141 256.663
R1110 B.n563 B.n343 256.663
R1111 B.n346 B.n343 256.663
R1112 B.n556 B.n343 256.663
R1113 B.n550 B.n343 256.663
R1114 B.n548 B.n343 256.663
R1115 B.n542 B.n343 256.663
R1116 B.n540 B.n343 256.663
R1117 B.n534 B.n343 256.663
R1118 B.n532 B.n343 256.663
R1119 B.n526 B.n343 256.663
R1120 B.n524 B.n343 256.663
R1121 B.n518 B.n343 256.663
R1122 B.n516 B.n343 256.663
R1123 B.n510 B.n343 256.663
R1124 B.n508 B.n343 256.663
R1125 B.n502 B.n343 256.663
R1126 B.n500 B.n343 256.663
R1127 B.n494 B.n343 256.663
R1128 B.n492 B.n343 256.663
R1129 B.n485 B.n343 256.663
R1130 B.n483 B.n343 256.663
R1131 B.n477 B.n343 256.663
R1132 B.n475 B.n343 256.663
R1133 B.n469 B.n343 256.663
R1134 B.n374 B.n343 256.663
R1135 B.n463 B.n343 256.663
R1136 B.n457 B.n343 256.663
R1137 B.n455 B.n343 256.663
R1138 B.n449 B.n343 256.663
R1139 B.n447 B.n343 256.663
R1140 B.n441 B.n343 256.663
R1141 B.n439 B.n343 256.663
R1142 B.n433 B.n343 256.663
R1143 B.n431 B.n343 256.663
R1144 B.n425 B.n343 256.663
R1145 B.n423 B.n343 256.663
R1146 B.n417 B.n343 256.663
R1147 B.n415 B.n343 256.663
R1148 B.n409 B.n343 256.663
R1149 B.n407 B.n343 256.663
R1150 B.n401 B.n343 256.663
R1151 B.n399 B.n343 256.663
R1152 B.n393 B.n343 256.663
R1153 B.n568 B.n338 163.367
R1154 B.n576 B.n338 163.367
R1155 B.n576 B.n336 163.367
R1156 B.n580 B.n336 163.367
R1157 B.n580 B.n330 163.367
R1158 B.n588 B.n330 163.367
R1159 B.n588 B.n328 163.367
R1160 B.n592 B.n328 163.367
R1161 B.n592 B.n322 163.367
R1162 B.n600 B.n322 163.367
R1163 B.n600 B.n320 163.367
R1164 B.n604 B.n320 163.367
R1165 B.n604 B.n314 163.367
R1166 B.n612 B.n314 163.367
R1167 B.n612 B.n312 163.367
R1168 B.n616 B.n312 163.367
R1169 B.n616 B.n306 163.367
R1170 B.n624 B.n306 163.367
R1171 B.n624 B.n304 163.367
R1172 B.n628 B.n304 163.367
R1173 B.n628 B.n298 163.367
R1174 B.n636 B.n298 163.367
R1175 B.n636 B.n296 163.367
R1176 B.n640 B.n296 163.367
R1177 B.n640 B.n290 163.367
R1178 B.n648 B.n290 163.367
R1179 B.n648 B.n288 163.367
R1180 B.n652 B.n288 163.367
R1181 B.n652 B.n282 163.367
R1182 B.n660 B.n282 163.367
R1183 B.n660 B.n280 163.367
R1184 B.n664 B.n280 163.367
R1185 B.n664 B.n274 163.367
R1186 B.n673 B.n274 163.367
R1187 B.n673 B.n272 163.367
R1188 B.n677 B.n272 163.367
R1189 B.n677 B.n267 163.367
R1190 B.n685 B.n267 163.367
R1191 B.n685 B.n265 163.367
R1192 B.n689 B.n265 163.367
R1193 B.n689 B.n259 163.367
R1194 B.n697 B.n259 163.367
R1195 B.n697 B.n257 163.367
R1196 B.n701 B.n257 163.367
R1197 B.n701 B.n251 163.367
R1198 B.n710 B.n251 163.367
R1199 B.n710 B.n249 163.367
R1200 B.n714 B.n249 163.367
R1201 B.n714 B.n244 163.367
R1202 B.n722 B.n244 163.367
R1203 B.n722 B.n242 163.367
R1204 B.n726 B.n242 163.367
R1205 B.n726 B.n236 163.367
R1206 B.n734 B.n236 163.367
R1207 B.n734 B.n234 163.367
R1208 B.n738 B.n234 163.367
R1209 B.n738 B.n228 163.367
R1210 B.n746 B.n228 163.367
R1211 B.n746 B.n226 163.367
R1212 B.n750 B.n226 163.367
R1213 B.n750 B.n220 163.367
R1214 B.n758 B.n220 163.367
R1215 B.n758 B.n218 163.367
R1216 B.n762 B.n218 163.367
R1217 B.n762 B.n212 163.367
R1218 B.n770 B.n212 163.367
R1219 B.n770 B.n210 163.367
R1220 B.n774 B.n210 163.367
R1221 B.n774 B.n204 163.367
R1222 B.n782 B.n204 163.367
R1223 B.n782 B.n202 163.367
R1224 B.n786 B.n202 163.367
R1225 B.n786 B.n196 163.367
R1226 B.n795 B.n196 163.367
R1227 B.n795 B.n194 163.367
R1228 B.n799 B.n194 163.367
R1229 B.n799 B.n2 163.367
R1230 B.n1236 B.n2 163.367
R1231 B.n1236 B.n3 163.367
R1232 B.n1232 B.n3 163.367
R1233 B.n1232 B.n9 163.367
R1234 B.n1228 B.n9 163.367
R1235 B.n1228 B.n11 163.367
R1236 B.n1224 B.n11 163.367
R1237 B.n1224 B.n16 163.367
R1238 B.n1220 B.n16 163.367
R1239 B.n1220 B.n18 163.367
R1240 B.n1216 B.n18 163.367
R1241 B.n1216 B.n23 163.367
R1242 B.n1212 B.n23 163.367
R1243 B.n1212 B.n25 163.367
R1244 B.n1208 B.n25 163.367
R1245 B.n1208 B.n30 163.367
R1246 B.n1204 B.n30 163.367
R1247 B.n1204 B.n32 163.367
R1248 B.n1200 B.n32 163.367
R1249 B.n1200 B.n37 163.367
R1250 B.n1196 B.n37 163.367
R1251 B.n1196 B.n39 163.367
R1252 B.n1192 B.n39 163.367
R1253 B.n1192 B.n44 163.367
R1254 B.n1188 B.n44 163.367
R1255 B.n1188 B.n46 163.367
R1256 B.n1184 B.n46 163.367
R1257 B.n1184 B.n51 163.367
R1258 B.n1180 B.n51 163.367
R1259 B.n1180 B.n53 163.367
R1260 B.n1176 B.n53 163.367
R1261 B.n1176 B.n57 163.367
R1262 B.n1172 B.n57 163.367
R1263 B.n1172 B.n59 163.367
R1264 B.n1168 B.n59 163.367
R1265 B.n1168 B.n65 163.367
R1266 B.n1164 B.n65 163.367
R1267 B.n1164 B.n67 163.367
R1268 B.n1160 B.n67 163.367
R1269 B.n1160 B.n72 163.367
R1270 B.n1156 B.n72 163.367
R1271 B.n1156 B.n74 163.367
R1272 B.n1152 B.n74 163.367
R1273 B.n1152 B.n78 163.367
R1274 B.n1148 B.n78 163.367
R1275 B.n1148 B.n80 163.367
R1276 B.n1144 B.n80 163.367
R1277 B.n1144 B.n86 163.367
R1278 B.n1140 B.n86 163.367
R1279 B.n1140 B.n88 163.367
R1280 B.n1136 B.n88 163.367
R1281 B.n1136 B.n93 163.367
R1282 B.n1132 B.n93 163.367
R1283 B.n1132 B.n95 163.367
R1284 B.n1128 B.n95 163.367
R1285 B.n1128 B.n100 163.367
R1286 B.n1124 B.n100 163.367
R1287 B.n1124 B.n102 163.367
R1288 B.n1120 B.n102 163.367
R1289 B.n1120 B.n107 163.367
R1290 B.n1116 B.n107 163.367
R1291 B.n1116 B.n109 163.367
R1292 B.n1112 B.n109 163.367
R1293 B.n1112 B.n114 163.367
R1294 B.n1108 B.n114 163.367
R1295 B.n1108 B.n116 163.367
R1296 B.n1104 B.n116 163.367
R1297 B.n1104 B.n121 163.367
R1298 B.n1100 B.n121 163.367
R1299 B.n1100 B.n123 163.367
R1300 B.n1096 B.n123 163.367
R1301 B.n1096 B.n128 163.367
R1302 B.n1092 B.n128 163.367
R1303 B.n1092 B.n130 163.367
R1304 B.n1088 B.n130 163.367
R1305 B.n1088 B.n135 163.367
R1306 B.n1084 B.n135 163.367
R1307 B.n1084 B.n137 163.367
R1308 B.n1080 B.n137 163.367
R1309 B.n564 B.n562 163.367
R1310 B.n562 B.n561 163.367
R1311 B.n558 B.n557 163.367
R1312 B.n555 B.n348 163.367
R1313 B.n551 B.n549 163.367
R1314 B.n547 B.n350 163.367
R1315 B.n543 B.n541 163.367
R1316 B.n539 B.n352 163.367
R1317 B.n535 B.n533 163.367
R1318 B.n531 B.n354 163.367
R1319 B.n527 B.n525 163.367
R1320 B.n523 B.n356 163.367
R1321 B.n519 B.n517 163.367
R1322 B.n515 B.n358 163.367
R1323 B.n511 B.n509 163.367
R1324 B.n507 B.n360 163.367
R1325 B.n503 B.n501 163.367
R1326 B.n499 B.n362 163.367
R1327 B.n495 B.n493 163.367
R1328 B.n491 B.n364 163.367
R1329 B.n486 B.n484 163.367
R1330 B.n482 B.n368 163.367
R1331 B.n478 B.n476 163.367
R1332 B.n474 B.n370 163.367
R1333 B.n470 B.n468 163.367
R1334 B.n465 B.n464 163.367
R1335 B.n462 B.n376 163.367
R1336 B.n458 B.n456 163.367
R1337 B.n454 B.n378 163.367
R1338 B.n450 B.n448 163.367
R1339 B.n446 B.n380 163.367
R1340 B.n442 B.n440 163.367
R1341 B.n438 B.n382 163.367
R1342 B.n434 B.n432 163.367
R1343 B.n430 B.n384 163.367
R1344 B.n426 B.n424 163.367
R1345 B.n422 B.n386 163.367
R1346 B.n418 B.n416 163.367
R1347 B.n414 B.n388 163.367
R1348 B.n410 B.n408 163.367
R1349 B.n406 B.n390 163.367
R1350 B.n402 B.n400 163.367
R1351 B.n398 B.n392 163.367
R1352 B.n394 B.n342 163.367
R1353 B.n570 B.n340 163.367
R1354 B.n574 B.n340 163.367
R1355 B.n574 B.n334 163.367
R1356 B.n582 B.n334 163.367
R1357 B.n582 B.n332 163.367
R1358 B.n586 B.n332 163.367
R1359 B.n586 B.n325 163.367
R1360 B.n594 B.n325 163.367
R1361 B.n594 B.n323 163.367
R1362 B.n598 B.n323 163.367
R1363 B.n598 B.n318 163.367
R1364 B.n606 B.n318 163.367
R1365 B.n606 B.n316 163.367
R1366 B.n610 B.n316 163.367
R1367 B.n610 B.n310 163.367
R1368 B.n618 B.n310 163.367
R1369 B.n618 B.n308 163.367
R1370 B.n622 B.n308 163.367
R1371 B.n622 B.n302 163.367
R1372 B.n630 B.n302 163.367
R1373 B.n630 B.n300 163.367
R1374 B.n634 B.n300 163.367
R1375 B.n634 B.n294 163.367
R1376 B.n642 B.n294 163.367
R1377 B.n642 B.n292 163.367
R1378 B.n646 B.n292 163.367
R1379 B.n646 B.n286 163.367
R1380 B.n654 B.n286 163.367
R1381 B.n654 B.n284 163.367
R1382 B.n658 B.n284 163.367
R1383 B.n658 B.n278 163.367
R1384 B.n666 B.n278 163.367
R1385 B.n666 B.n276 163.367
R1386 B.n670 B.n276 163.367
R1387 B.n670 B.n271 163.367
R1388 B.n679 B.n271 163.367
R1389 B.n679 B.n269 163.367
R1390 B.n683 B.n269 163.367
R1391 B.n683 B.n263 163.367
R1392 B.n691 B.n263 163.367
R1393 B.n691 B.n261 163.367
R1394 B.n695 B.n261 163.367
R1395 B.n695 B.n255 163.367
R1396 B.n703 B.n255 163.367
R1397 B.n703 B.n253 163.367
R1398 B.n707 B.n253 163.367
R1399 B.n707 B.n248 163.367
R1400 B.n716 B.n248 163.367
R1401 B.n716 B.n246 163.367
R1402 B.n720 B.n246 163.367
R1403 B.n720 B.n240 163.367
R1404 B.n728 B.n240 163.367
R1405 B.n728 B.n238 163.367
R1406 B.n732 B.n238 163.367
R1407 B.n732 B.n232 163.367
R1408 B.n740 B.n232 163.367
R1409 B.n740 B.n230 163.367
R1410 B.n744 B.n230 163.367
R1411 B.n744 B.n224 163.367
R1412 B.n752 B.n224 163.367
R1413 B.n752 B.n222 163.367
R1414 B.n756 B.n222 163.367
R1415 B.n756 B.n216 163.367
R1416 B.n764 B.n216 163.367
R1417 B.n764 B.n214 163.367
R1418 B.n768 B.n214 163.367
R1419 B.n768 B.n208 163.367
R1420 B.n776 B.n208 163.367
R1421 B.n776 B.n206 163.367
R1422 B.n780 B.n206 163.367
R1423 B.n780 B.n200 163.367
R1424 B.n788 B.n200 163.367
R1425 B.n788 B.n198 163.367
R1426 B.n793 B.n198 163.367
R1427 B.n793 B.n192 163.367
R1428 B.n801 B.n192 163.367
R1429 B.n802 B.n801 163.367
R1430 B.n802 B.n5 163.367
R1431 B.n6 B.n5 163.367
R1432 B.n7 B.n6 163.367
R1433 B.n807 B.n7 163.367
R1434 B.n807 B.n12 163.367
R1435 B.n13 B.n12 163.367
R1436 B.n14 B.n13 163.367
R1437 B.n812 B.n14 163.367
R1438 B.n812 B.n19 163.367
R1439 B.n20 B.n19 163.367
R1440 B.n21 B.n20 163.367
R1441 B.n817 B.n21 163.367
R1442 B.n817 B.n26 163.367
R1443 B.n27 B.n26 163.367
R1444 B.n28 B.n27 163.367
R1445 B.n822 B.n28 163.367
R1446 B.n822 B.n33 163.367
R1447 B.n34 B.n33 163.367
R1448 B.n35 B.n34 163.367
R1449 B.n827 B.n35 163.367
R1450 B.n827 B.n40 163.367
R1451 B.n41 B.n40 163.367
R1452 B.n42 B.n41 163.367
R1453 B.n832 B.n42 163.367
R1454 B.n832 B.n47 163.367
R1455 B.n48 B.n47 163.367
R1456 B.n49 B.n48 163.367
R1457 B.n837 B.n49 163.367
R1458 B.n837 B.n54 163.367
R1459 B.n55 B.n54 163.367
R1460 B.n56 B.n55 163.367
R1461 B.n842 B.n56 163.367
R1462 B.n842 B.n61 163.367
R1463 B.n62 B.n61 163.367
R1464 B.n63 B.n62 163.367
R1465 B.n847 B.n63 163.367
R1466 B.n847 B.n68 163.367
R1467 B.n69 B.n68 163.367
R1468 B.n70 B.n69 163.367
R1469 B.n852 B.n70 163.367
R1470 B.n852 B.n75 163.367
R1471 B.n76 B.n75 163.367
R1472 B.n77 B.n76 163.367
R1473 B.n857 B.n77 163.367
R1474 B.n857 B.n82 163.367
R1475 B.n83 B.n82 163.367
R1476 B.n84 B.n83 163.367
R1477 B.n862 B.n84 163.367
R1478 B.n862 B.n89 163.367
R1479 B.n90 B.n89 163.367
R1480 B.n91 B.n90 163.367
R1481 B.n867 B.n91 163.367
R1482 B.n867 B.n96 163.367
R1483 B.n97 B.n96 163.367
R1484 B.n98 B.n97 163.367
R1485 B.n872 B.n98 163.367
R1486 B.n872 B.n103 163.367
R1487 B.n104 B.n103 163.367
R1488 B.n105 B.n104 163.367
R1489 B.n877 B.n105 163.367
R1490 B.n877 B.n110 163.367
R1491 B.n111 B.n110 163.367
R1492 B.n112 B.n111 163.367
R1493 B.n882 B.n112 163.367
R1494 B.n882 B.n117 163.367
R1495 B.n118 B.n117 163.367
R1496 B.n119 B.n118 163.367
R1497 B.n887 B.n119 163.367
R1498 B.n887 B.n124 163.367
R1499 B.n125 B.n124 163.367
R1500 B.n126 B.n125 163.367
R1501 B.n892 B.n126 163.367
R1502 B.n892 B.n131 163.367
R1503 B.n132 B.n131 163.367
R1504 B.n133 B.n132 163.367
R1505 B.n897 B.n133 163.367
R1506 B.n897 B.n138 163.367
R1507 B.n139 B.n138 163.367
R1508 B.n140 B.n139 163.367
R1509 B.n1076 B.n1074 163.367
R1510 B.n1072 B.n144 163.367
R1511 B.n1068 B.n1066 163.367
R1512 B.n1064 B.n146 163.367
R1513 B.n1060 B.n1058 163.367
R1514 B.n1056 B.n148 163.367
R1515 B.n1052 B.n1050 163.367
R1516 B.n1048 B.n150 163.367
R1517 B.n1044 B.n1042 163.367
R1518 B.n1040 B.n152 163.367
R1519 B.n1036 B.n1034 163.367
R1520 B.n1032 B.n154 163.367
R1521 B.n1028 B.n1026 163.367
R1522 B.n1024 B.n156 163.367
R1523 B.n1020 B.n1018 163.367
R1524 B.n1016 B.n158 163.367
R1525 B.n1012 B.n1010 163.367
R1526 B.n1008 B.n160 163.367
R1527 B.n1004 B.n1002 163.367
R1528 B.n1000 B.n162 163.367
R1529 B.n996 B.n994 163.367
R1530 B.n992 B.n167 163.367
R1531 B.n988 B.n986 163.367
R1532 B.n984 B.n169 163.367
R1533 B.n979 B.n977 163.367
R1534 B.n975 B.n173 163.367
R1535 B.n971 B.n969 163.367
R1536 B.n967 B.n175 163.367
R1537 B.n963 B.n961 163.367
R1538 B.n959 B.n177 163.367
R1539 B.n955 B.n953 163.367
R1540 B.n951 B.n179 163.367
R1541 B.n947 B.n945 163.367
R1542 B.n943 B.n181 163.367
R1543 B.n939 B.n937 163.367
R1544 B.n935 B.n183 163.367
R1545 B.n931 B.n929 163.367
R1546 B.n927 B.n185 163.367
R1547 B.n923 B.n921 163.367
R1548 B.n919 B.n187 163.367
R1549 B.n915 B.n913 163.367
R1550 B.n911 B.n189 163.367
R1551 B.n907 B.n905 163.367
R1552 B.n371 B.t22 148.988
R1553 B.n170 B.t18 148.988
R1554 B.n365 B.t12 148.974
R1555 B.n163 B.t15 148.974
R1556 B.n372 B.n371 76.6066
R1557 B.n366 B.n365 76.6066
R1558 B.n164 B.n163 76.6066
R1559 B.n171 B.n170 76.6066
R1560 B.n569 B.n343 74.5199
R1561 B.n1081 B.n141 74.5199
R1562 B.n372 B.t21 72.3812
R1563 B.n171 B.t19 72.3812
R1564 B.n366 B.t11 72.3675
R1565 B.n164 B.t16 72.3675
R1566 B.n563 B.n344 71.676
R1567 B.n561 B.n346 71.676
R1568 B.n557 B.n556 71.676
R1569 B.n550 B.n348 71.676
R1570 B.n549 B.n548 71.676
R1571 B.n542 B.n350 71.676
R1572 B.n541 B.n540 71.676
R1573 B.n534 B.n352 71.676
R1574 B.n533 B.n532 71.676
R1575 B.n526 B.n354 71.676
R1576 B.n525 B.n524 71.676
R1577 B.n518 B.n356 71.676
R1578 B.n517 B.n516 71.676
R1579 B.n510 B.n358 71.676
R1580 B.n509 B.n508 71.676
R1581 B.n502 B.n360 71.676
R1582 B.n501 B.n500 71.676
R1583 B.n494 B.n362 71.676
R1584 B.n493 B.n492 71.676
R1585 B.n485 B.n364 71.676
R1586 B.n484 B.n483 71.676
R1587 B.n477 B.n368 71.676
R1588 B.n476 B.n475 71.676
R1589 B.n469 B.n370 71.676
R1590 B.n468 B.n374 71.676
R1591 B.n464 B.n463 71.676
R1592 B.n457 B.n376 71.676
R1593 B.n456 B.n455 71.676
R1594 B.n449 B.n378 71.676
R1595 B.n448 B.n447 71.676
R1596 B.n441 B.n380 71.676
R1597 B.n440 B.n439 71.676
R1598 B.n433 B.n382 71.676
R1599 B.n432 B.n431 71.676
R1600 B.n425 B.n384 71.676
R1601 B.n424 B.n423 71.676
R1602 B.n417 B.n386 71.676
R1603 B.n416 B.n415 71.676
R1604 B.n409 B.n388 71.676
R1605 B.n408 B.n407 71.676
R1606 B.n401 B.n390 71.676
R1607 B.n400 B.n399 71.676
R1608 B.n393 B.n392 71.676
R1609 B.n1075 B.n142 71.676
R1610 B.n1074 B.n1073 71.676
R1611 B.n1067 B.n144 71.676
R1612 B.n1066 B.n1065 71.676
R1613 B.n1059 B.n146 71.676
R1614 B.n1058 B.n1057 71.676
R1615 B.n1051 B.n148 71.676
R1616 B.n1050 B.n1049 71.676
R1617 B.n1043 B.n150 71.676
R1618 B.n1042 B.n1041 71.676
R1619 B.n1035 B.n152 71.676
R1620 B.n1034 B.n1033 71.676
R1621 B.n1027 B.n154 71.676
R1622 B.n1026 B.n1025 71.676
R1623 B.n1019 B.n156 71.676
R1624 B.n1018 B.n1017 71.676
R1625 B.n1011 B.n158 71.676
R1626 B.n1010 B.n1009 71.676
R1627 B.n1003 B.n160 71.676
R1628 B.n1002 B.n1001 71.676
R1629 B.n995 B.n162 71.676
R1630 B.n994 B.n993 71.676
R1631 B.n987 B.n167 71.676
R1632 B.n986 B.n985 71.676
R1633 B.n978 B.n169 71.676
R1634 B.n977 B.n976 71.676
R1635 B.n970 B.n173 71.676
R1636 B.n969 B.n968 71.676
R1637 B.n962 B.n175 71.676
R1638 B.n961 B.n960 71.676
R1639 B.n954 B.n177 71.676
R1640 B.n953 B.n952 71.676
R1641 B.n946 B.n179 71.676
R1642 B.n945 B.n944 71.676
R1643 B.n938 B.n181 71.676
R1644 B.n937 B.n936 71.676
R1645 B.n930 B.n183 71.676
R1646 B.n929 B.n928 71.676
R1647 B.n922 B.n185 71.676
R1648 B.n921 B.n920 71.676
R1649 B.n914 B.n187 71.676
R1650 B.n913 B.n912 71.676
R1651 B.n906 B.n189 71.676
R1652 B.n905 B.n904 71.676
R1653 B.n904 B.n903 71.676
R1654 B.n907 B.n906 71.676
R1655 B.n912 B.n911 71.676
R1656 B.n915 B.n914 71.676
R1657 B.n920 B.n919 71.676
R1658 B.n923 B.n922 71.676
R1659 B.n928 B.n927 71.676
R1660 B.n931 B.n930 71.676
R1661 B.n936 B.n935 71.676
R1662 B.n939 B.n938 71.676
R1663 B.n944 B.n943 71.676
R1664 B.n947 B.n946 71.676
R1665 B.n952 B.n951 71.676
R1666 B.n955 B.n954 71.676
R1667 B.n960 B.n959 71.676
R1668 B.n963 B.n962 71.676
R1669 B.n968 B.n967 71.676
R1670 B.n971 B.n970 71.676
R1671 B.n976 B.n975 71.676
R1672 B.n979 B.n978 71.676
R1673 B.n985 B.n984 71.676
R1674 B.n988 B.n987 71.676
R1675 B.n993 B.n992 71.676
R1676 B.n996 B.n995 71.676
R1677 B.n1001 B.n1000 71.676
R1678 B.n1004 B.n1003 71.676
R1679 B.n1009 B.n1008 71.676
R1680 B.n1012 B.n1011 71.676
R1681 B.n1017 B.n1016 71.676
R1682 B.n1020 B.n1019 71.676
R1683 B.n1025 B.n1024 71.676
R1684 B.n1028 B.n1027 71.676
R1685 B.n1033 B.n1032 71.676
R1686 B.n1036 B.n1035 71.676
R1687 B.n1041 B.n1040 71.676
R1688 B.n1044 B.n1043 71.676
R1689 B.n1049 B.n1048 71.676
R1690 B.n1052 B.n1051 71.676
R1691 B.n1057 B.n1056 71.676
R1692 B.n1060 B.n1059 71.676
R1693 B.n1065 B.n1064 71.676
R1694 B.n1068 B.n1067 71.676
R1695 B.n1073 B.n1072 71.676
R1696 B.n1076 B.n1075 71.676
R1697 B.n564 B.n563 71.676
R1698 B.n558 B.n346 71.676
R1699 B.n556 B.n555 71.676
R1700 B.n551 B.n550 71.676
R1701 B.n548 B.n547 71.676
R1702 B.n543 B.n542 71.676
R1703 B.n540 B.n539 71.676
R1704 B.n535 B.n534 71.676
R1705 B.n532 B.n531 71.676
R1706 B.n527 B.n526 71.676
R1707 B.n524 B.n523 71.676
R1708 B.n519 B.n518 71.676
R1709 B.n516 B.n515 71.676
R1710 B.n511 B.n510 71.676
R1711 B.n508 B.n507 71.676
R1712 B.n503 B.n502 71.676
R1713 B.n500 B.n499 71.676
R1714 B.n495 B.n494 71.676
R1715 B.n492 B.n491 71.676
R1716 B.n486 B.n485 71.676
R1717 B.n483 B.n482 71.676
R1718 B.n478 B.n477 71.676
R1719 B.n475 B.n474 71.676
R1720 B.n470 B.n469 71.676
R1721 B.n465 B.n374 71.676
R1722 B.n463 B.n462 71.676
R1723 B.n458 B.n457 71.676
R1724 B.n455 B.n454 71.676
R1725 B.n450 B.n449 71.676
R1726 B.n447 B.n446 71.676
R1727 B.n442 B.n441 71.676
R1728 B.n439 B.n438 71.676
R1729 B.n434 B.n433 71.676
R1730 B.n431 B.n430 71.676
R1731 B.n426 B.n425 71.676
R1732 B.n423 B.n422 71.676
R1733 B.n418 B.n417 71.676
R1734 B.n415 B.n414 71.676
R1735 B.n410 B.n409 71.676
R1736 B.n407 B.n406 71.676
R1737 B.n402 B.n401 71.676
R1738 B.n399 B.n398 71.676
R1739 B.n394 B.n393 71.676
R1740 B.n373 B.n372 59.5399
R1741 B.n489 B.n366 59.5399
R1742 B.n165 B.n164 59.5399
R1743 B.n981 B.n171 59.5399
R1744 B.n569 B.n339 45.652
R1745 B.n575 B.n339 45.652
R1746 B.n575 B.n335 45.652
R1747 B.n581 B.n335 45.652
R1748 B.n581 B.n331 45.652
R1749 B.n587 B.n331 45.652
R1750 B.n587 B.n326 45.652
R1751 B.n593 B.n326 45.652
R1752 B.n593 B.n327 45.652
R1753 B.n599 B.n319 45.652
R1754 B.n605 B.n319 45.652
R1755 B.n605 B.n315 45.652
R1756 B.n611 B.n315 45.652
R1757 B.n611 B.n311 45.652
R1758 B.n617 B.n311 45.652
R1759 B.n617 B.n307 45.652
R1760 B.n623 B.n307 45.652
R1761 B.n623 B.n303 45.652
R1762 B.n629 B.n303 45.652
R1763 B.n629 B.n299 45.652
R1764 B.n635 B.n299 45.652
R1765 B.n635 B.n295 45.652
R1766 B.n641 B.n295 45.652
R1767 B.n647 B.n291 45.652
R1768 B.n647 B.n287 45.652
R1769 B.n653 B.n287 45.652
R1770 B.n653 B.n283 45.652
R1771 B.n659 B.n283 45.652
R1772 B.n659 B.n279 45.652
R1773 B.n665 B.n279 45.652
R1774 B.n665 B.n275 45.652
R1775 B.n672 B.n275 45.652
R1776 B.n672 B.n671 45.652
R1777 B.n678 B.n268 45.652
R1778 B.n684 B.n268 45.652
R1779 B.n684 B.n264 45.652
R1780 B.n690 B.n264 45.652
R1781 B.n690 B.n260 45.652
R1782 B.n696 B.n260 45.652
R1783 B.n696 B.n256 45.652
R1784 B.n702 B.n256 45.652
R1785 B.n702 B.n252 45.652
R1786 B.n709 B.n252 45.652
R1787 B.n709 B.n708 45.652
R1788 B.n715 B.n245 45.652
R1789 B.n721 B.n245 45.652
R1790 B.n721 B.n241 45.652
R1791 B.n727 B.n241 45.652
R1792 B.n727 B.n237 45.652
R1793 B.n733 B.n237 45.652
R1794 B.n733 B.n233 45.652
R1795 B.n739 B.n233 45.652
R1796 B.n739 B.n229 45.652
R1797 B.n745 B.n229 45.652
R1798 B.n751 B.n225 45.652
R1799 B.n751 B.n221 45.652
R1800 B.n757 B.n221 45.652
R1801 B.n757 B.n217 45.652
R1802 B.n763 B.n217 45.652
R1803 B.n763 B.n213 45.652
R1804 B.n769 B.n213 45.652
R1805 B.n769 B.n209 45.652
R1806 B.n775 B.n209 45.652
R1807 B.n775 B.n205 45.652
R1808 B.n781 B.n205 45.652
R1809 B.n787 B.n201 45.652
R1810 B.n787 B.n197 45.652
R1811 B.n794 B.n197 45.652
R1812 B.n794 B.n193 45.652
R1813 B.n800 B.n193 45.652
R1814 B.n800 B.n4 45.652
R1815 B.n1235 B.n4 45.652
R1816 B.n1235 B.n1234 45.652
R1817 B.n1234 B.n1233 45.652
R1818 B.n1233 B.n8 45.652
R1819 B.n1227 B.n8 45.652
R1820 B.n1227 B.n1226 45.652
R1821 B.n1226 B.n1225 45.652
R1822 B.n1225 B.n15 45.652
R1823 B.n1219 B.n1218 45.652
R1824 B.n1218 B.n1217 45.652
R1825 B.n1217 B.n22 45.652
R1826 B.n1211 B.n22 45.652
R1827 B.n1211 B.n1210 45.652
R1828 B.n1210 B.n1209 45.652
R1829 B.n1209 B.n29 45.652
R1830 B.n1203 B.n29 45.652
R1831 B.n1203 B.n1202 45.652
R1832 B.n1202 B.n1201 45.652
R1833 B.n1201 B.n36 45.652
R1834 B.n1195 B.n1194 45.652
R1835 B.n1194 B.n1193 45.652
R1836 B.n1193 B.n43 45.652
R1837 B.n1187 B.n43 45.652
R1838 B.n1187 B.n1186 45.652
R1839 B.n1186 B.n1185 45.652
R1840 B.n1185 B.n50 45.652
R1841 B.n1179 B.n50 45.652
R1842 B.n1179 B.n1178 45.652
R1843 B.n1178 B.n1177 45.652
R1844 B.n1171 B.n60 45.652
R1845 B.n1171 B.n1170 45.652
R1846 B.n1170 B.n1169 45.652
R1847 B.n1169 B.n64 45.652
R1848 B.n1163 B.n64 45.652
R1849 B.n1163 B.n1162 45.652
R1850 B.n1162 B.n1161 45.652
R1851 B.n1161 B.n71 45.652
R1852 B.n1155 B.n71 45.652
R1853 B.n1155 B.n1154 45.652
R1854 B.n1154 B.n1153 45.652
R1855 B.n1147 B.n81 45.652
R1856 B.n1147 B.n1146 45.652
R1857 B.n1146 B.n1145 45.652
R1858 B.n1145 B.n85 45.652
R1859 B.n1139 B.n85 45.652
R1860 B.n1139 B.n1138 45.652
R1861 B.n1138 B.n1137 45.652
R1862 B.n1137 B.n92 45.652
R1863 B.n1131 B.n92 45.652
R1864 B.n1131 B.n1130 45.652
R1865 B.n1129 B.n99 45.652
R1866 B.n1123 B.n99 45.652
R1867 B.n1123 B.n1122 45.652
R1868 B.n1122 B.n1121 45.652
R1869 B.n1121 B.n106 45.652
R1870 B.n1115 B.n106 45.652
R1871 B.n1115 B.n1114 45.652
R1872 B.n1114 B.n1113 45.652
R1873 B.n1113 B.n113 45.652
R1874 B.n1107 B.n113 45.652
R1875 B.n1107 B.n1106 45.652
R1876 B.n1106 B.n1105 45.652
R1877 B.n1105 B.n120 45.652
R1878 B.n1099 B.n120 45.652
R1879 B.n1098 B.n1097 45.652
R1880 B.n1097 B.n127 45.652
R1881 B.n1091 B.n127 45.652
R1882 B.n1091 B.n1090 45.652
R1883 B.n1090 B.n1089 45.652
R1884 B.n1089 B.n134 45.652
R1885 B.n1083 B.n134 45.652
R1886 B.n1083 B.n1082 45.652
R1887 B.n1082 B.n1081 45.652
R1888 B.n745 B.t7 44.3093
R1889 B.n1195 B.t2 44.3093
R1890 B.t23 B.n291 40.2812
R1891 B.n1130 B.t0 40.2812
R1892 B.n671 B.t5 33.5678
R1893 B.n81 B.t8 33.5678
R1894 B.n599 B.t10 32.2251
R1895 B.n1099 B.t14 32.2251
R1896 B.n715 B.t1 29.5397
R1897 B.n1177 B.t3 29.5397
R1898 B.n1079 B.n1078 28.2542
R1899 B.n902 B.n901 28.2542
R1900 B.n571 B.n341 28.2542
R1901 B.n567 B.n566 28.2542
R1902 B.n781 B.t6 26.8543
R1903 B.n1219 B.t4 26.8543
R1904 B.t6 B.n201 18.7982
R1905 B.t4 B.n15 18.7982
R1906 B B.n1237 18.0485
R1907 B.n708 B.t1 16.1128
R1908 B.n60 B.t3 16.1128
R1909 B.n327 B.t10 13.4274
R1910 B.t14 B.n1098 13.4274
R1911 B.n678 B.t5 12.0847
R1912 B.n1153 B.t8 12.0847
R1913 B.n1078 B.n1077 10.6151
R1914 B.n1077 B.n143 10.6151
R1915 B.n1071 B.n143 10.6151
R1916 B.n1071 B.n1070 10.6151
R1917 B.n1070 B.n1069 10.6151
R1918 B.n1069 B.n145 10.6151
R1919 B.n1063 B.n145 10.6151
R1920 B.n1063 B.n1062 10.6151
R1921 B.n1062 B.n1061 10.6151
R1922 B.n1061 B.n147 10.6151
R1923 B.n1055 B.n147 10.6151
R1924 B.n1055 B.n1054 10.6151
R1925 B.n1054 B.n1053 10.6151
R1926 B.n1053 B.n149 10.6151
R1927 B.n1047 B.n149 10.6151
R1928 B.n1047 B.n1046 10.6151
R1929 B.n1046 B.n1045 10.6151
R1930 B.n1045 B.n151 10.6151
R1931 B.n1039 B.n151 10.6151
R1932 B.n1039 B.n1038 10.6151
R1933 B.n1038 B.n1037 10.6151
R1934 B.n1037 B.n153 10.6151
R1935 B.n1031 B.n153 10.6151
R1936 B.n1031 B.n1030 10.6151
R1937 B.n1030 B.n1029 10.6151
R1938 B.n1029 B.n155 10.6151
R1939 B.n1023 B.n155 10.6151
R1940 B.n1023 B.n1022 10.6151
R1941 B.n1022 B.n1021 10.6151
R1942 B.n1021 B.n157 10.6151
R1943 B.n1015 B.n157 10.6151
R1944 B.n1015 B.n1014 10.6151
R1945 B.n1014 B.n1013 10.6151
R1946 B.n1013 B.n159 10.6151
R1947 B.n1007 B.n159 10.6151
R1948 B.n1007 B.n1006 10.6151
R1949 B.n1006 B.n1005 10.6151
R1950 B.n1005 B.n161 10.6151
R1951 B.n999 B.n998 10.6151
R1952 B.n998 B.n997 10.6151
R1953 B.n997 B.n166 10.6151
R1954 B.n991 B.n166 10.6151
R1955 B.n991 B.n990 10.6151
R1956 B.n990 B.n989 10.6151
R1957 B.n989 B.n168 10.6151
R1958 B.n983 B.n168 10.6151
R1959 B.n983 B.n982 10.6151
R1960 B.n980 B.n172 10.6151
R1961 B.n974 B.n172 10.6151
R1962 B.n974 B.n973 10.6151
R1963 B.n973 B.n972 10.6151
R1964 B.n972 B.n174 10.6151
R1965 B.n966 B.n174 10.6151
R1966 B.n966 B.n965 10.6151
R1967 B.n965 B.n964 10.6151
R1968 B.n964 B.n176 10.6151
R1969 B.n958 B.n176 10.6151
R1970 B.n958 B.n957 10.6151
R1971 B.n957 B.n956 10.6151
R1972 B.n956 B.n178 10.6151
R1973 B.n950 B.n178 10.6151
R1974 B.n950 B.n949 10.6151
R1975 B.n949 B.n948 10.6151
R1976 B.n948 B.n180 10.6151
R1977 B.n942 B.n180 10.6151
R1978 B.n942 B.n941 10.6151
R1979 B.n941 B.n940 10.6151
R1980 B.n940 B.n182 10.6151
R1981 B.n934 B.n182 10.6151
R1982 B.n934 B.n933 10.6151
R1983 B.n933 B.n932 10.6151
R1984 B.n932 B.n184 10.6151
R1985 B.n926 B.n184 10.6151
R1986 B.n926 B.n925 10.6151
R1987 B.n925 B.n924 10.6151
R1988 B.n924 B.n186 10.6151
R1989 B.n918 B.n186 10.6151
R1990 B.n918 B.n917 10.6151
R1991 B.n917 B.n916 10.6151
R1992 B.n916 B.n188 10.6151
R1993 B.n910 B.n188 10.6151
R1994 B.n910 B.n909 10.6151
R1995 B.n909 B.n908 10.6151
R1996 B.n908 B.n190 10.6151
R1997 B.n902 B.n190 10.6151
R1998 B.n572 B.n571 10.6151
R1999 B.n573 B.n572 10.6151
R2000 B.n573 B.n333 10.6151
R2001 B.n583 B.n333 10.6151
R2002 B.n584 B.n583 10.6151
R2003 B.n585 B.n584 10.6151
R2004 B.n585 B.n324 10.6151
R2005 B.n595 B.n324 10.6151
R2006 B.n596 B.n595 10.6151
R2007 B.n597 B.n596 10.6151
R2008 B.n597 B.n317 10.6151
R2009 B.n607 B.n317 10.6151
R2010 B.n608 B.n607 10.6151
R2011 B.n609 B.n608 10.6151
R2012 B.n609 B.n309 10.6151
R2013 B.n619 B.n309 10.6151
R2014 B.n620 B.n619 10.6151
R2015 B.n621 B.n620 10.6151
R2016 B.n621 B.n301 10.6151
R2017 B.n631 B.n301 10.6151
R2018 B.n632 B.n631 10.6151
R2019 B.n633 B.n632 10.6151
R2020 B.n633 B.n293 10.6151
R2021 B.n643 B.n293 10.6151
R2022 B.n644 B.n643 10.6151
R2023 B.n645 B.n644 10.6151
R2024 B.n645 B.n285 10.6151
R2025 B.n655 B.n285 10.6151
R2026 B.n656 B.n655 10.6151
R2027 B.n657 B.n656 10.6151
R2028 B.n657 B.n277 10.6151
R2029 B.n667 B.n277 10.6151
R2030 B.n668 B.n667 10.6151
R2031 B.n669 B.n668 10.6151
R2032 B.n669 B.n270 10.6151
R2033 B.n680 B.n270 10.6151
R2034 B.n681 B.n680 10.6151
R2035 B.n682 B.n681 10.6151
R2036 B.n682 B.n262 10.6151
R2037 B.n692 B.n262 10.6151
R2038 B.n693 B.n692 10.6151
R2039 B.n694 B.n693 10.6151
R2040 B.n694 B.n254 10.6151
R2041 B.n704 B.n254 10.6151
R2042 B.n705 B.n704 10.6151
R2043 B.n706 B.n705 10.6151
R2044 B.n706 B.n247 10.6151
R2045 B.n717 B.n247 10.6151
R2046 B.n718 B.n717 10.6151
R2047 B.n719 B.n718 10.6151
R2048 B.n719 B.n239 10.6151
R2049 B.n729 B.n239 10.6151
R2050 B.n730 B.n729 10.6151
R2051 B.n731 B.n730 10.6151
R2052 B.n731 B.n231 10.6151
R2053 B.n741 B.n231 10.6151
R2054 B.n742 B.n741 10.6151
R2055 B.n743 B.n742 10.6151
R2056 B.n743 B.n223 10.6151
R2057 B.n753 B.n223 10.6151
R2058 B.n754 B.n753 10.6151
R2059 B.n755 B.n754 10.6151
R2060 B.n755 B.n215 10.6151
R2061 B.n765 B.n215 10.6151
R2062 B.n766 B.n765 10.6151
R2063 B.n767 B.n766 10.6151
R2064 B.n767 B.n207 10.6151
R2065 B.n777 B.n207 10.6151
R2066 B.n778 B.n777 10.6151
R2067 B.n779 B.n778 10.6151
R2068 B.n779 B.n199 10.6151
R2069 B.n789 B.n199 10.6151
R2070 B.n790 B.n789 10.6151
R2071 B.n792 B.n790 10.6151
R2072 B.n792 B.n791 10.6151
R2073 B.n791 B.n191 10.6151
R2074 B.n803 B.n191 10.6151
R2075 B.n804 B.n803 10.6151
R2076 B.n805 B.n804 10.6151
R2077 B.n806 B.n805 10.6151
R2078 B.n808 B.n806 10.6151
R2079 B.n809 B.n808 10.6151
R2080 B.n810 B.n809 10.6151
R2081 B.n811 B.n810 10.6151
R2082 B.n813 B.n811 10.6151
R2083 B.n814 B.n813 10.6151
R2084 B.n815 B.n814 10.6151
R2085 B.n816 B.n815 10.6151
R2086 B.n818 B.n816 10.6151
R2087 B.n819 B.n818 10.6151
R2088 B.n820 B.n819 10.6151
R2089 B.n821 B.n820 10.6151
R2090 B.n823 B.n821 10.6151
R2091 B.n824 B.n823 10.6151
R2092 B.n825 B.n824 10.6151
R2093 B.n826 B.n825 10.6151
R2094 B.n828 B.n826 10.6151
R2095 B.n829 B.n828 10.6151
R2096 B.n830 B.n829 10.6151
R2097 B.n831 B.n830 10.6151
R2098 B.n833 B.n831 10.6151
R2099 B.n834 B.n833 10.6151
R2100 B.n835 B.n834 10.6151
R2101 B.n836 B.n835 10.6151
R2102 B.n838 B.n836 10.6151
R2103 B.n839 B.n838 10.6151
R2104 B.n840 B.n839 10.6151
R2105 B.n841 B.n840 10.6151
R2106 B.n843 B.n841 10.6151
R2107 B.n844 B.n843 10.6151
R2108 B.n845 B.n844 10.6151
R2109 B.n846 B.n845 10.6151
R2110 B.n848 B.n846 10.6151
R2111 B.n849 B.n848 10.6151
R2112 B.n850 B.n849 10.6151
R2113 B.n851 B.n850 10.6151
R2114 B.n853 B.n851 10.6151
R2115 B.n854 B.n853 10.6151
R2116 B.n855 B.n854 10.6151
R2117 B.n856 B.n855 10.6151
R2118 B.n858 B.n856 10.6151
R2119 B.n859 B.n858 10.6151
R2120 B.n860 B.n859 10.6151
R2121 B.n861 B.n860 10.6151
R2122 B.n863 B.n861 10.6151
R2123 B.n864 B.n863 10.6151
R2124 B.n865 B.n864 10.6151
R2125 B.n866 B.n865 10.6151
R2126 B.n868 B.n866 10.6151
R2127 B.n869 B.n868 10.6151
R2128 B.n870 B.n869 10.6151
R2129 B.n871 B.n870 10.6151
R2130 B.n873 B.n871 10.6151
R2131 B.n874 B.n873 10.6151
R2132 B.n875 B.n874 10.6151
R2133 B.n876 B.n875 10.6151
R2134 B.n878 B.n876 10.6151
R2135 B.n879 B.n878 10.6151
R2136 B.n880 B.n879 10.6151
R2137 B.n881 B.n880 10.6151
R2138 B.n883 B.n881 10.6151
R2139 B.n884 B.n883 10.6151
R2140 B.n885 B.n884 10.6151
R2141 B.n886 B.n885 10.6151
R2142 B.n888 B.n886 10.6151
R2143 B.n889 B.n888 10.6151
R2144 B.n890 B.n889 10.6151
R2145 B.n891 B.n890 10.6151
R2146 B.n893 B.n891 10.6151
R2147 B.n894 B.n893 10.6151
R2148 B.n895 B.n894 10.6151
R2149 B.n896 B.n895 10.6151
R2150 B.n898 B.n896 10.6151
R2151 B.n899 B.n898 10.6151
R2152 B.n900 B.n899 10.6151
R2153 B.n901 B.n900 10.6151
R2154 B.n566 B.n565 10.6151
R2155 B.n565 B.n345 10.6151
R2156 B.n560 B.n345 10.6151
R2157 B.n560 B.n559 10.6151
R2158 B.n559 B.n347 10.6151
R2159 B.n554 B.n347 10.6151
R2160 B.n554 B.n553 10.6151
R2161 B.n553 B.n552 10.6151
R2162 B.n552 B.n349 10.6151
R2163 B.n546 B.n349 10.6151
R2164 B.n546 B.n545 10.6151
R2165 B.n545 B.n544 10.6151
R2166 B.n544 B.n351 10.6151
R2167 B.n538 B.n351 10.6151
R2168 B.n538 B.n537 10.6151
R2169 B.n537 B.n536 10.6151
R2170 B.n536 B.n353 10.6151
R2171 B.n530 B.n353 10.6151
R2172 B.n530 B.n529 10.6151
R2173 B.n529 B.n528 10.6151
R2174 B.n528 B.n355 10.6151
R2175 B.n522 B.n355 10.6151
R2176 B.n522 B.n521 10.6151
R2177 B.n521 B.n520 10.6151
R2178 B.n520 B.n357 10.6151
R2179 B.n514 B.n357 10.6151
R2180 B.n514 B.n513 10.6151
R2181 B.n513 B.n512 10.6151
R2182 B.n512 B.n359 10.6151
R2183 B.n506 B.n359 10.6151
R2184 B.n506 B.n505 10.6151
R2185 B.n505 B.n504 10.6151
R2186 B.n504 B.n361 10.6151
R2187 B.n498 B.n361 10.6151
R2188 B.n498 B.n497 10.6151
R2189 B.n497 B.n496 10.6151
R2190 B.n496 B.n363 10.6151
R2191 B.n490 B.n363 10.6151
R2192 B.n488 B.n487 10.6151
R2193 B.n487 B.n367 10.6151
R2194 B.n481 B.n367 10.6151
R2195 B.n481 B.n480 10.6151
R2196 B.n480 B.n479 10.6151
R2197 B.n479 B.n369 10.6151
R2198 B.n473 B.n369 10.6151
R2199 B.n473 B.n472 10.6151
R2200 B.n472 B.n471 10.6151
R2201 B.n467 B.n466 10.6151
R2202 B.n466 B.n375 10.6151
R2203 B.n461 B.n375 10.6151
R2204 B.n461 B.n460 10.6151
R2205 B.n460 B.n459 10.6151
R2206 B.n459 B.n377 10.6151
R2207 B.n453 B.n377 10.6151
R2208 B.n453 B.n452 10.6151
R2209 B.n452 B.n451 10.6151
R2210 B.n451 B.n379 10.6151
R2211 B.n445 B.n379 10.6151
R2212 B.n445 B.n444 10.6151
R2213 B.n444 B.n443 10.6151
R2214 B.n443 B.n381 10.6151
R2215 B.n437 B.n381 10.6151
R2216 B.n437 B.n436 10.6151
R2217 B.n436 B.n435 10.6151
R2218 B.n435 B.n383 10.6151
R2219 B.n429 B.n383 10.6151
R2220 B.n429 B.n428 10.6151
R2221 B.n428 B.n427 10.6151
R2222 B.n427 B.n385 10.6151
R2223 B.n421 B.n385 10.6151
R2224 B.n421 B.n420 10.6151
R2225 B.n420 B.n419 10.6151
R2226 B.n419 B.n387 10.6151
R2227 B.n413 B.n387 10.6151
R2228 B.n413 B.n412 10.6151
R2229 B.n412 B.n411 10.6151
R2230 B.n411 B.n389 10.6151
R2231 B.n405 B.n389 10.6151
R2232 B.n405 B.n404 10.6151
R2233 B.n404 B.n403 10.6151
R2234 B.n403 B.n391 10.6151
R2235 B.n397 B.n391 10.6151
R2236 B.n397 B.n396 10.6151
R2237 B.n396 B.n395 10.6151
R2238 B.n395 B.n341 10.6151
R2239 B.n567 B.n337 10.6151
R2240 B.n577 B.n337 10.6151
R2241 B.n578 B.n577 10.6151
R2242 B.n579 B.n578 10.6151
R2243 B.n579 B.n329 10.6151
R2244 B.n589 B.n329 10.6151
R2245 B.n590 B.n589 10.6151
R2246 B.n591 B.n590 10.6151
R2247 B.n591 B.n321 10.6151
R2248 B.n601 B.n321 10.6151
R2249 B.n602 B.n601 10.6151
R2250 B.n603 B.n602 10.6151
R2251 B.n603 B.n313 10.6151
R2252 B.n613 B.n313 10.6151
R2253 B.n614 B.n613 10.6151
R2254 B.n615 B.n614 10.6151
R2255 B.n615 B.n305 10.6151
R2256 B.n625 B.n305 10.6151
R2257 B.n626 B.n625 10.6151
R2258 B.n627 B.n626 10.6151
R2259 B.n627 B.n297 10.6151
R2260 B.n637 B.n297 10.6151
R2261 B.n638 B.n637 10.6151
R2262 B.n639 B.n638 10.6151
R2263 B.n639 B.n289 10.6151
R2264 B.n649 B.n289 10.6151
R2265 B.n650 B.n649 10.6151
R2266 B.n651 B.n650 10.6151
R2267 B.n651 B.n281 10.6151
R2268 B.n661 B.n281 10.6151
R2269 B.n662 B.n661 10.6151
R2270 B.n663 B.n662 10.6151
R2271 B.n663 B.n273 10.6151
R2272 B.n674 B.n273 10.6151
R2273 B.n675 B.n674 10.6151
R2274 B.n676 B.n675 10.6151
R2275 B.n676 B.n266 10.6151
R2276 B.n686 B.n266 10.6151
R2277 B.n687 B.n686 10.6151
R2278 B.n688 B.n687 10.6151
R2279 B.n688 B.n258 10.6151
R2280 B.n698 B.n258 10.6151
R2281 B.n699 B.n698 10.6151
R2282 B.n700 B.n699 10.6151
R2283 B.n700 B.n250 10.6151
R2284 B.n711 B.n250 10.6151
R2285 B.n712 B.n711 10.6151
R2286 B.n713 B.n712 10.6151
R2287 B.n713 B.n243 10.6151
R2288 B.n723 B.n243 10.6151
R2289 B.n724 B.n723 10.6151
R2290 B.n725 B.n724 10.6151
R2291 B.n725 B.n235 10.6151
R2292 B.n735 B.n235 10.6151
R2293 B.n736 B.n735 10.6151
R2294 B.n737 B.n736 10.6151
R2295 B.n737 B.n227 10.6151
R2296 B.n747 B.n227 10.6151
R2297 B.n748 B.n747 10.6151
R2298 B.n749 B.n748 10.6151
R2299 B.n749 B.n219 10.6151
R2300 B.n759 B.n219 10.6151
R2301 B.n760 B.n759 10.6151
R2302 B.n761 B.n760 10.6151
R2303 B.n761 B.n211 10.6151
R2304 B.n771 B.n211 10.6151
R2305 B.n772 B.n771 10.6151
R2306 B.n773 B.n772 10.6151
R2307 B.n773 B.n203 10.6151
R2308 B.n783 B.n203 10.6151
R2309 B.n784 B.n783 10.6151
R2310 B.n785 B.n784 10.6151
R2311 B.n785 B.n195 10.6151
R2312 B.n796 B.n195 10.6151
R2313 B.n797 B.n796 10.6151
R2314 B.n798 B.n797 10.6151
R2315 B.n798 B.n0 10.6151
R2316 B.n1231 B.n1 10.6151
R2317 B.n1231 B.n1230 10.6151
R2318 B.n1230 B.n1229 10.6151
R2319 B.n1229 B.n10 10.6151
R2320 B.n1223 B.n10 10.6151
R2321 B.n1223 B.n1222 10.6151
R2322 B.n1222 B.n1221 10.6151
R2323 B.n1221 B.n17 10.6151
R2324 B.n1215 B.n17 10.6151
R2325 B.n1215 B.n1214 10.6151
R2326 B.n1214 B.n1213 10.6151
R2327 B.n1213 B.n24 10.6151
R2328 B.n1207 B.n24 10.6151
R2329 B.n1207 B.n1206 10.6151
R2330 B.n1206 B.n1205 10.6151
R2331 B.n1205 B.n31 10.6151
R2332 B.n1199 B.n31 10.6151
R2333 B.n1199 B.n1198 10.6151
R2334 B.n1198 B.n1197 10.6151
R2335 B.n1197 B.n38 10.6151
R2336 B.n1191 B.n38 10.6151
R2337 B.n1191 B.n1190 10.6151
R2338 B.n1190 B.n1189 10.6151
R2339 B.n1189 B.n45 10.6151
R2340 B.n1183 B.n45 10.6151
R2341 B.n1183 B.n1182 10.6151
R2342 B.n1182 B.n1181 10.6151
R2343 B.n1181 B.n52 10.6151
R2344 B.n1175 B.n52 10.6151
R2345 B.n1175 B.n1174 10.6151
R2346 B.n1174 B.n1173 10.6151
R2347 B.n1173 B.n58 10.6151
R2348 B.n1167 B.n58 10.6151
R2349 B.n1167 B.n1166 10.6151
R2350 B.n1166 B.n1165 10.6151
R2351 B.n1165 B.n66 10.6151
R2352 B.n1159 B.n66 10.6151
R2353 B.n1159 B.n1158 10.6151
R2354 B.n1158 B.n1157 10.6151
R2355 B.n1157 B.n73 10.6151
R2356 B.n1151 B.n73 10.6151
R2357 B.n1151 B.n1150 10.6151
R2358 B.n1150 B.n1149 10.6151
R2359 B.n1149 B.n79 10.6151
R2360 B.n1143 B.n79 10.6151
R2361 B.n1143 B.n1142 10.6151
R2362 B.n1142 B.n1141 10.6151
R2363 B.n1141 B.n87 10.6151
R2364 B.n1135 B.n87 10.6151
R2365 B.n1135 B.n1134 10.6151
R2366 B.n1134 B.n1133 10.6151
R2367 B.n1133 B.n94 10.6151
R2368 B.n1127 B.n94 10.6151
R2369 B.n1127 B.n1126 10.6151
R2370 B.n1126 B.n1125 10.6151
R2371 B.n1125 B.n101 10.6151
R2372 B.n1119 B.n101 10.6151
R2373 B.n1119 B.n1118 10.6151
R2374 B.n1118 B.n1117 10.6151
R2375 B.n1117 B.n108 10.6151
R2376 B.n1111 B.n108 10.6151
R2377 B.n1111 B.n1110 10.6151
R2378 B.n1110 B.n1109 10.6151
R2379 B.n1109 B.n115 10.6151
R2380 B.n1103 B.n115 10.6151
R2381 B.n1103 B.n1102 10.6151
R2382 B.n1102 B.n1101 10.6151
R2383 B.n1101 B.n122 10.6151
R2384 B.n1095 B.n122 10.6151
R2385 B.n1095 B.n1094 10.6151
R2386 B.n1094 B.n1093 10.6151
R2387 B.n1093 B.n129 10.6151
R2388 B.n1087 B.n129 10.6151
R2389 B.n1087 B.n1086 10.6151
R2390 B.n1086 B.n1085 10.6151
R2391 B.n1085 B.n136 10.6151
R2392 B.n1079 B.n136 10.6151
R2393 B.n165 B.n161 9.36635
R2394 B.n981 B.n980 9.36635
R2395 B.n490 B.n489 9.36635
R2396 B.n467 B.n373 9.36635
R2397 B.n641 B.t23 5.37127
R2398 B.t0 B.n1129 5.37127
R2399 B.n1237 B.n0 2.81026
R2400 B.n1237 B.n1 2.81026
R2401 B.t7 B.n225 1.34319
R2402 B.t2 B.n36 1.34319
R2403 B.n999 B.n165 1.24928
R2404 B.n982 B.n981 1.24928
R2405 B.n489 B.n488 1.24928
R2406 B.n471 B.n373 1.24928
R2407 VN.n106 VN.n105 161.3
R2408 VN.n104 VN.n55 161.3
R2409 VN.n103 VN.n102 161.3
R2410 VN.n101 VN.n56 161.3
R2411 VN.n100 VN.n99 161.3
R2412 VN.n98 VN.n57 161.3
R2413 VN.n97 VN.n96 161.3
R2414 VN.n95 VN.n58 161.3
R2415 VN.n94 VN.n93 161.3
R2416 VN.n92 VN.n59 161.3
R2417 VN.n91 VN.n90 161.3
R2418 VN.n89 VN.n61 161.3
R2419 VN.n88 VN.n87 161.3
R2420 VN.n86 VN.n62 161.3
R2421 VN.n85 VN.n84 161.3
R2422 VN.n83 VN.n63 161.3
R2423 VN.n82 VN.n81 161.3
R2424 VN.n80 VN.n64 161.3
R2425 VN.n79 VN.n78 161.3
R2426 VN.n77 VN.n66 161.3
R2427 VN.n76 VN.n75 161.3
R2428 VN.n74 VN.n67 161.3
R2429 VN.n73 VN.n72 161.3
R2430 VN.n71 VN.n68 161.3
R2431 VN.n52 VN.n51 161.3
R2432 VN.n50 VN.n1 161.3
R2433 VN.n49 VN.n48 161.3
R2434 VN.n47 VN.n2 161.3
R2435 VN.n46 VN.n45 161.3
R2436 VN.n44 VN.n3 161.3
R2437 VN.n43 VN.n42 161.3
R2438 VN.n41 VN.n4 161.3
R2439 VN.n40 VN.n39 161.3
R2440 VN.n37 VN.n5 161.3
R2441 VN.n36 VN.n35 161.3
R2442 VN.n34 VN.n6 161.3
R2443 VN.n33 VN.n32 161.3
R2444 VN.n31 VN.n7 161.3
R2445 VN.n30 VN.n29 161.3
R2446 VN.n28 VN.n8 161.3
R2447 VN.n27 VN.n26 161.3
R2448 VN.n24 VN.n9 161.3
R2449 VN.n23 VN.n22 161.3
R2450 VN.n21 VN.n10 161.3
R2451 VN.n20 VN.n19 161.3
R2452 VN.n18 VN.n11 161.3
R2453 VN.n17 VN.n16 161.3
R2454 VN.n15 VN.n12 161.3
R2455 VN.n70 VN.t6 106.894
R2456 VN.n14 VN.t2 106.894
R2457 VN.n53 VN.n0 82.7273
R2458 VN.n107 VN.n54 82.7273
R2459 VN.n13 VN.t8 73.9649
R2460 VN.n25 VN.t1 73.9649
R2461 VN.n38 VN.t5 73.9649
R2462 VN.n0 VN.t9 73.9649
R2463 VN.n69 VN.t4 73.9649
R2464 VN.n65 VN.t3 73.9649
R2465 VN.n60 VN.t0 73.9649
R2466 VN.n54 VN.t7 73.9649
R2467 VN.n70 VN.n69 64.731
R2468 VN.n14 VN.n13 64.731
R2469 VN VN.n107 58.2291
R2470 VN.n19 VN.n10 56.5193
R2471 VN.n32 VN.n6 56.5193
R2472 VN.n45 VN.n2 56.5193
R2473 VN.n75 VN.n66 56.5193
R2474 VN.n87 VN.n61 56.5193
R2475 VN.n99 VN.n56 56.5193
R2476 VN.n17 VN.n12 24.4675
R2477 VN.n18 VN.n17 24.4675
R2478 VN.n19 VN.n18 24.4675
R2479 VN.n23 VN.n10 24.4675
R2480 VN.n24 VN.n23 24.4675
R2481 VN.n26 VN.n24 24.4675
R2482 VN.n30 VN.n8 24.4675
R2483 VN.n31 VN.n30 24.4675
R2484 VN.n32 VN.n31 24.4675
R2485 VN.n36 VN.n6 24.4675
R2486 VN.n37 VN.n36 24.4675
R2487 VN.n39 VN.n37 24.4675
R2488 VN.n43 VN.n4 24.4675
R2489 VN.n44 VN.n43 24.4675
R2490 VN.n45 VN.n44 24.4675
R2491 VN.n49 VN.n2 24.4675
R2492 VN.n50 VN.n49 24.4675
R2493 VN.n51 VN.n50 24.4675
R2494 VN.n75 VN.n74 24.4675
R2495 VN.n74 VN.n73 24.4675
R2496 VN.n73 VN.n68 24.4675
R2497 VN.n87 VN.n86 24.4675
R2498 VN.n86 VN.n85 24.4675
R2499 VN.n85 VN.n63 24.4675
R2500 VN.n81 VN.n80 24.4675
R2501 VN.n80 VN.n79 24.4675
R2502 VN.n79 VN.n66 24.4675
R2503 VN.n99 VN.n98 24.4675
R2504 VN.n98 VN.n97 24.4675
R2505 VN.n97 VN.n58 24.4675
R2506 VN.n93 VN.n92 24.4675
R2507 VN.n92 VN.n91 24.4675
R2508 VN.n91 VN.n61 24.4675
R2509 VN.n105 VN.n104 24.4675
R2510 VN.n104 VN.n103 24.4675
R2511 VN.n103 VN.n56 24.4675
R2512 VN.n38 VN.n4 14.6807
R2513 VN.n60 VN.n58 14.6807
R2514 VN.n26 VN.n25 12.234
R2515 VN.n25 VN.n8 12.234
R2516 VN.n65 VN.n63 12.234
R2517 VN.n81 VN.n65 12.234
R2518 VN.n13 VN.n12 9.7873
R2519 VN.n39 VN.n38 9.7873
R2520 VN.n69 VN.n68 9.7873
R2521 VN.n93 VN.n60 9.7873
R2522 VN.n51 VN.n0 7.3406
R2523 VN.n105 VN.n54 7.3406
R2524 VN.n71 VN.n70 3.24375
R2525 VN.n15 VN.n14 3.24375
R2526 VN.n107 VN.n106 0.354971
R2527 VN.n53 VN.n52 0.354971
R2528 VN VN.n53 0.26696
R2529 VN.n106 VN.n55 0.189894
R2530 VN.n102 VN.n55 0.189894
R2531 VN.n102 VN.n101 0.189894
R2532 VN.n101 VN.n100 0.189894
R2533 VN.n100 VN.n57 0.189894
R2534 VN.n96 VN.n57 0.189894
R2535 VN.n96 VN.n95 0.189894
R2536 VN.n95 VN.n94 0.189894
R2537 VN.n94 VN.n59 0.189894
R2538 VN.n90 VN.n59 0.189894
R2539 VN.n90 VN.n89 0.189894
R2540 VN.n89 VN.n88 0.189894
R2541 VN.n88 VN.n62 0.189894
R2542 VN.n84 VN.n62 0.189894
R2543 VN.n84 VN.n83 0.189894
R2544 VN.n83 VN.n82 0.189894
R2545 VN.n82 VN.n64 0.189894
R2546 VN.n78 VN.n64 0.189894
R2547 VN.n78 VN.n77 0.189894
R2548 VN.n77 VN.n76 0.189894
R2549 VN.n76 VN.n67 0.189894
R2550 VN.n72 VN.n67 0.189894
R2551 VN.n72 VN.n71 0.189894
R2552 VN.n16 VN.n15 0.189894
R2553 VN.n16 VN.n11 0.189894
R2554 VN.n20 VN.n11 0.189894
R2555 VN.n21 VN.n20 0.189894
R2556 VN.n22 VN.n21 0.189894
R2557 VN.n22 VN.n9 0.189894
R2558 VN.n27 VN.n9 0.189894
R2559 VN.n28 VN.n27 0.189894
R2560 VN.n29 VN.n28 0.189894
R2561 VN.n29 VN.n7 0.189894
R2562 VN.n33 VN.n7 0.189894
R2563 VN.n34 VN.n33 0.189894
R2564 VN.n35 VN.n34 0.189894
R2565 VN.n35 VN.n5 0.189894
R2566 VN.n40 VN.n5 0.189894
R2567 VN.n41 VN.n40 0.189894
R2568 VN.n42 VN.n41 0.189894
R2569 VN.n42 VN.n3 0.189894
R2570 VN.n46 VN.n3 0.189894
R2571 VN.n47 VN.n46 0.189894
R2572 VN.n48 VN.n47 0.189894
R2573 VN.n48 VN.n1 0.189894
R2574 VN.n52 VN.n1 0.189894
R2575 VDD2.n1 VDD2.t7 68.7539
R2576 VDD2.n3 VDD2.n2 66.065
R2577 VDD2 VDD2.n7 66.0622
R2578 VDD2.n4 VDD2.t2 65.3488
R2579 VDD2.n6 VDD2.n5 63.5667
R2580 VDD2.n1 VDD2.n0 63.5665
R2581 VDD2.n4 VDD2.n3 49.4674
R2582 VDD2.n6 VDD2.n4 3.40567
R2583 VDD2.n7 VDD2.t5 1.78268
R2584 VDD2.n7 VDD2.t3 1.78268
R2585 VDD2.n5 VDD2.t9 1.78268
R2586 VDD2.n5 VDD2.t6 1.78268
R2587 VDD2.n2 VDD2.t4 1.78268
R2588 VDD2.n2 VDD2.t0 1.78268
R2589 VDD2.n0 VDD2.t1 1.78268
R2590 VDD2.n0 VDD2.t8 1.78268
R2591 VDD2 VDD2.n6 0.909983
R2592 VDD2.n3 VDD2.n1 0.796447
C0 VTAIL VDD1 10.531f
C1 VDD1 VP 11.045599f
C2 VDD2 VDD1 2.84008f
C3 VDD1 VN 0.155869f
C4 VTAIL VP 11.6275f
C5 VDD2 VTAIL 10.5898f
C6 VTAIL VN 11.6132f
C7 VDD2 VP 0.713736f
C8 VP VN 9.73832f
C9 VDD2 VN 10.4915f
C10 VDD2 B 8.250154f
C11 VDD1 B 8.215906f
C12 VTAIL B 8.623637f
C13 VN B 22.941929f
C14 VP B 21.531853f
C15 VDD2.t7 B 2.50177f
C16 VDD2.t1 B 0.218759f
C17 VDD2.t8 B 0.218759f
C18 VDD2.n0 B 1.94114f
C19 VDD2.n1 B 1.06503f
C20 VDD2.t4 B 0.218759f
C21 VDD2.t0 B 0.218759f
C22 VDD2.n2 B 1.96716f
C23 VDD2.n3 B 3.36856f
C24 VDD2.t2 B 2.47452f
C25 VDD2.n4 B 3.43827f
C26 VDD2.t9 B 0.218759f
C27 VDD2.t6 B 0.218759f
C28 VDD2.n5 B 1.94114f
C29 VDD2.n6 B 0.550205f
C30 VDD2.t5 B 0.218759f
C31 VDD2.t3 B 0.218759f
C32 VDD2.n7 B 1.96711f
C33 VN.t9 B 1.91289f
C34 VN.n0 B 0.740373f
C35 VN.n1 B 0.017497f
C36 VN.n2 B 0.0292f
C37 VN.n3 B 0.017497f
C38 VN.n4 B 0.02617f
C39 VN.n5 B 0.017497f
C40 VN.n6 B 0.026763f
C41 VN.n7 B 0.017497f
C42 VN.n8 B 0.02456f
C43 VN.n9 B 0.017497f
C44 VN.n10 B 0.024325f
C45 VN.n11 B 0.017497f
C46 VN.n12 B 0.02295f
C47 VN.t8 B 1.91289f
C48 VN.n13 B 0.732753f
C49 VN.t2 B 2.16126f
C50 VN.n14 B 0.696328f
C51 VN.n15 B 0.219501f
C52 VN.n16 B 0.017497f
C53 VN.n17 B 0.032609f
C54 VN.n18 B 0.032609f
C55 VN.n19 B 0.026763f
C56 VN.n20 B 0.017497f
C57 VN.n21 B 0.017497f
C58 VN.n22 B 0.017497f
C59 VN.n23 B 0.032609f
C60 VN.n24 B 0.032609f
C61 VN.t1 B 1.91289f
C62 VN.n25 B 0.673452f
C63 VN.n26 B 0.02456f
C64 VN.n27 B 0.017497f
C65 VN.n28 B 0.017497f
C66 VN.n29 B 0.017497f
C67 VN.n30 B 0.032609f
C68 VN.n31 B 0.032609f
C69 VN.n32 B 0.024325f
C70 VN.n33 B 0.017497f
C71 VN.n34 B 0.017497f
C72 VN.n35 B 0.017497f
C73 VN.n36 B 0.032609f
C74 VN.n37 B 0.032609f
C75 VN.t5 B 1.91289f
C76 VN.n38 B 0.673452f
C77 VN.n39 B 0.02295f
C78 VN.n40 B 0.017497f
C79 VN.n41 B 0.017497f
C80 VN.n42 B 0.017497f
C81 VN.n43 B 0.032609f
C82 VN.n44 B 0.032609f
C83 VN.n45 B 0.021887f
C84 VN.n46 B 0.017497f
C85 VN.n47 B 0.017497f
C86 VN.n48 B 0.017497f
C87 VN.n49 B 0.032609f
C88 VN.n50 B 0.032609f
C89 VN.n51 B 0.02134f
C90 VN.n52 B 0.028239f
C91 VN.n53 B 0.049625f
C92 VN.t7 B 1.91289f
C93 VN.n54 B 0.740373f
C94 VN.n55 B 0.017497f
C95 VN.n56 B 0.0292f
C96 VN.n57 B 0.017497f
C97 VN.n58 B 0.02617f
C98 VN.n59 B 0.017497f
C99 VN.t0 B 1.91289f
C100 VN.n60 B 0.673452f
C101 VN.n61 B 0.026763f
C102 VN.n62 B 0.017497f
C103 VN.n63 B 0.02456f
C104 VN.n64 B 0.017497f
C105 VN.t3 B 1.91289f
C106 VN.n65 B 0.673452f
C107 VN.n66 B 0.024325f
C108 VN.n67 B 0.017497f
C109 VN.n68 B 0.02295f
C110 VN.t6 B 2.16126f
C111 VN.t4 B 1.91289f
C112 VN.n69 B 0.732753f
C113 VN.n70 B 0.696327f
C114 VN.n71 B 0.219501f
C115 VN.n72 B 0.017497f
C116 VN.n73 B 0.032609f
C117 VN.n74 B 0.032609f
C118 VN.n75 B 0.026763f
C119 VN.n76 B 0.017497f
C120 VN.n77 B 0.017497f
C121 VN.n78 B 0.017497f
C122 VN.n79 B 0.032609f
C123 VN.n80 B 0.032609f
C124 VN.n81 B 0.02456f
C125 VN.n82 B 0.017497f
C126 VN.n83 B 0.017497f
C127 VN.n84 B 0.017497f
C128 VN.n85 B 0.032609f
C129 VN.n86 B 0.032609f
C130 VN.n87 B 0.024325f
C131 VN.n88 B 0.017497f
C132 VN.n89 B 0.017497f
C133 VN.n90 B 0.017497f
C134 VN.n91 B 0.032609f
C135 VN.n92 B 0.032609f
C136 VN.n93 B 0.02295f
C137 VN.n94 B 0.017497f
C138 VN.n95 B 0.017497f
C139 VN.n96 B 0.017497f
C140 VN.n97 B 0.032609f
C141 VN.n98 B 0.032609f
C142 VN.n99 B 0.021887f
C143 VN.n100 B 0.017497f
C144 VN.n101 B 0.017497f
C145 VN.n102 B 0.017497f
C146 VN.n103 B 0.032609f
C147 VN.n104 B 0.032609f
C148 VN.n105 B 0.02134f
C149 VN.n106 B 0.028239f
C150 VN.n107 B 1.24016f
C151 VDD1.t3 B 2.5339f
C152 VDD1.t5 B 0.221567f
C153 VDD1.t9 B 0.221567f
C154 VDD1.n0 B 1.96606f
C155 VDD1.n1 B 1.08718f
C156 VDD1.t0 B 2.53388f
C157 VDD1.t4 B 0.221567f
C158 VDD1.t8 B 0.221567f
C159 VDD1.n2 B 1.96606f
C160 VDD1.n3 B 1.0787f
C161 VDD1.t1 B 0.221567f
C162 VDD1.t6 B 0.221567f
C163 VDD1.n4 B 1.99241f
C164 VDD1.n5 B 3.56565f
C165 VDD1.t2 B 0.221567f
C166 VDD1.t7 B 0.221567f
C167 VDD1.n6 B 1.96605f
C168 VDD1.n7 B 3.56067f
C169 VTAIL.t4 B 0.22877f
C170 VTAIL.t2 B 0.22877f
C171 VTAIL.n0 B 1.95592f
C172 VTAIL.n1 B 0.653463f
C173 VTAIL.t11 B 2.49374f
C174 VTAIL.n2 B 0.806151f
C175 VTAIL.t18 B 0.22877f
C176 VTAIL.t10 B 0.22877f
C177 VTAIL.n3 B 1.95592f
C178 VTAIL.n4 B 0.82356f
C179 VTAIL.t14 B 0.22877f
C180 VTAIL.t13 B 0.22877f
C181 VTAIL.n5 B 1.95592f
C182 VTAIL.n6 B 2.26759f
C183 VTAIL.t19 B 0.22877f
C184 VTAIL.t5 B 0.22877f
C185 VTAIL.n7 B 1.95593f
C186 VTAIL.n8 B 2.26758f
C187 VTAIL.t1 B 0.22877f
C188 VTAIL.t7 B 0.22877f
C189 VTAIL.n9 B 1.95593f
C190 VTAIL.n10 B 0.823554f
C191 VTAIL.t6 B 2.49376f
C192 VTAIL.n11 B 0.806135f
C193 VTAIL.t12 B 0.22877f
C194 VTAIL.t9 B 0.22877f
C195 VTAIL.n12 B 1.95593f
C196 VTAIL.n13 B 0.720048f
C197 VTAIL.t17 B 0.22877f
C198 VTAIL.t15 B 0.22877f
C199 VTAIL.n14 B 1.95593f
C200 VTAIL.n15 B 0.823554f
C201 VTAIL.t16 B 2.49374f
C202 VTAIL.n16 B 2.06778f
C203 VTAIL.t0 B 2.49374f
C204 VTAIL.n17 B 2.06778f
C205 VTAIL.t3 B 0.22877f
C206 VTAIL.t8 B 0.22877f
C207 VTAIL.n18 B 1.95592f
C208 VTAIL.n19 B 0.604244f
C209 VP.t3 B 1.94447f
C210 VP.n0 B 0.752596f
C211 VP.n1 B 0.017786f
C212 VP.n2 B 0.029682f
C213 VP.n3 B 0.017786f
C214 VP.n4 B 0.026602f
C215 VP.n5 B 0.017786f
C216 VP.n6 B 0.027204f
C217 VP.n7 B 0.017786f
C218 VP.n8 B 0.024965f
C219 VP.n9 B 0.017786f
C220 VP.n10 B 0.024726f
C221 VP.n11 B 0.017786f
C222 VP.n12 B 0.023329f
C223 VP.n13 B 0.017786f
C224 VP.n14 B 0.022248f
C225 VP.n15 B 0.017786f
C226 VP.n16 B 0.021692f
C227 VP.t2 B 1.94447f
C228 VP.n17 B 0.752596f
C229 VP.n18 B 0.017786f
C230 VP.n19 B 0.029682f
C231 VP.n20 B 0.017786f
C232 VP.n21 B 0.026602f
C233 VP.n22 B 0.017786f
C234 VP.n23 B 0.027204f
C235 VP.n24 B 0.017786f
C236 VP.n25 B 0.024965f
C237 VP.n26 B 0.017786f
C238 VP.n27 B 0.024726f
C239 VP.n28 B 0.017786f
C240 VP.n29 B 0.023329f
C241 VP.t6 B 2.19694f
C242 VP.t4 B 1.94447f
C243 VP.n30 B 0.74485f
C244 VP.n31 B 0.707824f
C245 VP.n32 B 0.223125f
C246 VP.n33 B 0.017786f
C247 VP.n34 B 0.033148f
C248 VP.n35 B 0.033148f
C249 VP.n36 B 0.027204f
C250 VP.n37 B 0.017786f
C251 VP.n38 B 0.017786f
C252 VP.n39 B 0.017786f
C253 VP.n40 B 0.033148f
C254 VP.n41 B 0.033148f
C255 VP.t0 B 1.94447f
C256 VP.n42 B 0.68457f
C257 VP.n43 B 0.024965f
C258 VP.n44 B 0.017786f
C259 VP.n45 B 0.017786f
C260 VP.n46 B 0.017786f
C261 VP.n47 B 0.033148f
C262 VP.n48 B 0.033148f
C263 VP.n49 B 0.024726f
C264 VP.n50 B 0.017786f
C265 VP.n51 B 0.017786f
C266 VP.n52 B 0.017786f
C267 VP.n53 B 0.033148f
C268 VP.n54 B 0.033148f
C269 VP.t7 B 1.94447f
C270 VP.n55 B 0.68457f
C271 VP.n56 B 0.023329f
C272 VP.n57 B 0.017786f
C273 VP.n58 B 0.017786f
C274 VP.n59 B 0.017786f
C275 VP.n60 B 0.033148f
C276 VP.n61 B 0.033148f
C277 VP.n62 B 0.022248f
C278 VP.n63 B 0.017786f
C279 VP.n64 B 0.017786f
C280 VP.n65 B 0.017786f
C281 VP.n66 B 0.033148f
C282 VP.n67 B 0.033148f
C283 VP.n68 B 0.021692f
C284 VP.n69 B 0.028706f
C285 VP.n70 B 1.25371f
C286 VP.t9 B 1.94447f
C287 VP.n71 B 0.752596f
C288 VP.n72 B 1.26472f
C289 VP.n73 B 0.028706f
C290 VP.n74 B 0.017786f
C291 VP.n75 B 0.033148f
C292 VP.n76 B 0.033148f
C293 VP.n77 B 0.029682f
C294 VP.n78 B 0.017786f
C295 VP.n79 B 0.017786f
C296 VP.n80 B 0.017786f
C297 VP.n81 B 0.033148f
C298 VP.n82 B 0.033148f
C299 VP.t5 B 1.94447f
C300 VP.n83 B 0.68457f
C301 VP.n84 B 0.026602f
C302 VP.n85 B 0.017786f
C303 VP.n86 B 0.017786f
C304 VP.n87 B 0.017786f
C305 VP.n88 B 0.033148f
C306 VP.n89 B 0.033148f
C307 VP.n90 B 0.027204f
C308 VP.n91 B 0.017786f
C309 VP.n92 B 0.017786f
C310 VP.n93 B 0.017786f
C311 VP.n94 B 0.033148f
C312 VP.n95 B 0.033148f
C313 VP.t1 B 1.94447f
C314 VP.n96 B 0.68457f
C315 VP.n97 B 0.024965f
C316 VP.n98 B 0.017786f
C317 VP.n99 B 0.017786f
C318 VP.n100 B 0.017786f
C319 VP.n101 B 0.033148f
C320 VP.n102 B 0.033148f
C321 VP.n103 B 0.024726f
C322 VP.n104 B 0.017786f
C323 VP.n105 B 0.017786f
C324 VP.n106 B 0.017786f
C325 VP.n107 B 0.033148f
C326 VP.n108 B 0.033148f
C327 VP.t8 B 1.94447f
C328 VP.n109 B 0.68457f
C329 VP.n110 B 0.023329f
C330 VP.n111 B 0.017786f
C331 VP.n112 B 0.017786f
C332 VP.n113 B 0.017786f
C333 VP.n114 B 0.033148f
C334 VP.n115 B 0.033148f
C335 VP.n116 B 0.022248f
C336 VP.n117 B 0.017786f
C337 VP.n118 B 0.017786f
C338 VP.n119 B 0.017786f
C339 VP.n120 B 0.033148f
C340 VP.n121 B 0.033148f
C341 VP.n122 B 0.021692f
C342 VP.n123 B 0.028706f
C343 VP.n124 B 0.050445f
.ends

