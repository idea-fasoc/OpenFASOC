* NGSPICE file created from diff_pair_sample_1331.ext - technology: sky130A

.subckt diff_pair_sample_1331 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t3 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=0.73095 ps=4.76 w=4.43 l=0.44
X1 B.t11 B.t9 B.t10 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0 ps=0 w=4.43 l=0.44
X2 VDD1.t1 VP.t1 VTAIL.t10 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=1.7277 ps=9.64 w=4.43 l=0.44
X3 VDD1.t0 VP.t2 VTAIL.t9 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0.73095 ps=4.76 w=4.43 l=0.44
X4 B.t8 B.t6 B.t7 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0 ps=0 w=4.43 l=0.44
X5 B.t5 B.t3 B.t4 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0 ps=0 w=4.43 l=0.44
X6 VDD2.t5 VN.t0 VTAIL.t1 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=1.7277 ps=9.64 w=4.43 l=0.44
X7 VDD1.t5 VP.t3 VTAIL.t8 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=1.7277 ps=9.64 w=4.43 l=0.44
X8 VDD2.t4 VN.t1 VTAIL.t0 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0.73095 ps=4.76 w=4.43 l=0.44
X9 VTAIL.t5 VN.t2 VDD2.t3 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=0.73095 ps=4.76 w=4.43 l=0.44
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=1.7277 ps=9.64 w=4.43 l=0.44
X11 VTAIL.t7 VP.t4 VDD1.t4 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=0.73095 ps=4.76 w=4.43 l=0.44
X12 VTAIL.t3 VN.t4 VDD2.t1 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=0.73095 pd=4.76 as=0.73095 ps=4.76 w=4.43 l=0.44
X13 B.t2 B.t0 B.t1 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0 ps=0 w=4.43 l=0.44
X14 VDD2.t0 VN.t5 VTAIL.t2 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0.73095 ps=4.76 w=4.43 l=0.44
X15 VDD1.t2 VP.t5 VTAIL.t6 w_n1586_n1854# sky130_fd_pr__pfet_01v8 ad=1.7277 pd=9.64 as=0.73095 ps=4.76 w=4.43 l=0.44
R0 VP.n1 VP.t5 357.935
R1 VP.n8 VP.t1 339.774
R2 VP.n6 VP.t2 339.774
R3 VP.n3 VP.t3 339.774
R4 VP.n7 VP.t4 332.471
R5 VP.n2 VP.t0 332.471
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n7 VP.n0 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n4 VP.n1 71.8132
R11 VP.n7 VP.n6 40.8975
R12 VP.n8 VP.n7 40.8975
R13 VP.n3 VP.n2 40.8975
R14 VP.n5 VP.n4 34.5649
R15 VP.n2 VP.n1 18.1394
R16 VP.n5 VP.n0 0.189894
R17 VP.n9 VP.n0 0.189894
R18 VP VP.n9 0.0516364
R19 VDD1.n20 VDD1.n19 756.745
R20 VDD1.n41 VDD1.n40 756.745
R21 VDD1.n19 VDD1.n18 585
R22 VDD1.n2 VDD1.n1 585
R23 VDD1.n13 VDD1.n12 585
R24 VDD1.n11 VDD1.n10 585
R25 VDD1.n6 VDD1.n5 585
R26 VDD1.n27 VDD1.n26 585
R27 VDD1.n32 VDD1.n31 585
R28 VDD1.n34 VDD1.n33 585
R29 VDD1.n23 VDD1.n22 585
R30 VDD1.n40 VDD1.n39 585
R31 VDD1.n28 VDD1.t0 330.188
R32 VDD1.n7 VDD1.t2 330.188
R33 VDD1.n19 VDD1.n1 171.744
R34 VDD1.n12 VDD1.n1 171.744
R35 VDD1.n12 VDD1.n11 171.744
R36 VDD1.n11 VDD1.n5 171.744
R37 VDD1.n32 VDD1.n26 171.744
R38 VDD1.n33 VDD1.n32 171.744
R39 VDD1.n33 VDD1.n22 171.744
R40 VDD1.n40 VDD1.n22 171.744
R41 VDD1.n43 VDD1.n42 107.617
R42 VDD1.n45 VDD1.n44 107.504
R43 VDD1.t2 VDD1.n5 85.8723
R44 VDD1.t0 VDD1.n26 85.8723
R45 VDD1 VDD1.n20 51.1656
R46 VDD1.n43 VDD1.n41 51.0521
R47 VDD1.n45 VDD1.n43 30.6065
R48 VDD1.n7 VDD1.n6 10.7082
R49 VDD1.n28 VDD1.n27 10.7082
R50 VDD1.n18 VDD1.n0 10.4732
R51 VDD1.n39 VDD1.n21 10.4732
R52 VDD1.n17 VDD1.n2 9.69747
R53 VDD1.n38 VDD1.n23 9.69747
R54 VDD1.n16 VDD1.n0 9.45567
R55 VDD1.n37 VDD1.n21 9.45567
R56 VDD1.n4 VDD1.n3 9.3005
R57 VDD1.n15 VDD1.n14 9.3005
R58 VDD1.n17 VDD1.n16 9.3005
R59 VDD1.n9 VDD1.n8 9.3005
R60 VDD1.n30 VDD1.n29 9.3005
R61 VDD1.n25 VDD1.n24 9.3005
R62 VDD1.n36 VDD1.n35 9.3005
R63 VDD1.n38 VDD1.n37 9.3005
R64 VDD1.n14 VDD1.n13 8.92171
R65 VDD1.n35 VDD1.n34 8.92171
R66 VDD1.n10 VDD1.n4 8.14595
R67 VDD1.n31 VDD1.n25 8.14595
R68 VDD1.n9 VDD1.n6 7.3702
R69 VDD1.n30 VDD1.n27 7.3702
R70 VDD1.n44 VDD1.t3 7.33797
R71 VDD1.n44 VDD1.t5 7.33797
R72 VDD1.n42 VDD1.t4 7.33797
R73 VDD1.n42 VDD1.t1 7.33797
R74 VDD1.n10 VDD1.n9 5.81868
R75 VDD1.n31 VDD1.n30 5.81868
R76 VDD1.n13 VDD1.n4 5.04292
R77 VDD1.n34 VDD1.n25 5.04292
R78 VDD1.n14 VDD1.n2 4.26717
R79 VDD1.n35 VDD1.n23 4.26717
R80 VDD1.n18 VDD1.n17 3.49141
R81 VDD1.n39 VDD1.n38 3.49141
R82 VDD1.n20 VDD1.n0 2.71565
R83 VDD1.n41 VDD1.n21 2.71565
R84 VDD1.n8 VDD1.n7 2.42873
R85 VDD1.n29 VDD1.n28 2.42873
R86 VDD1.n16 VDD1.n15 0.155672
R87 VDD1.n15 VDD1.n3 0.155672
R88 VDD1.n8 VDD1.n3 0.155672
R89 VDD1.n29 VDD1.n24 0.155672
R90 VDD1.n36 VDD1.n24 0.155672
R91 VDD1.n37 VDD1.n36 0.155672
R92 VDD1 VDD1.n45 0.108259
R93 VTAIL.n94 VTAIL.n93 756.745
R94 VTAIL.n22 VTAIL.n21 756.745
R95 VTAIL.n72 VTAIL.n71 756.745
R96 VTAIL.n48 VTAIL.n47 756.745
R97 VTAIL.n80 VTAIL.n79 585
R98 VTAIL.n85 VTAIL.n84 585
R99 VTAIL.n87 VTAIL.n86 585
R100 VTAIL.n76 VTAIL.n75 585
R101 VTAIL.n93 VTAIL.n92 585
R102 VTAIL.n8 VTAIL.n7 585
R103 VTAIL.n13 VTAIL.n12 585
R104 VTAIL.n15 VTAIL.n14 585
R105 VTAIL.n4 VTAIL.n3 585
R106 VTAIL.n21 VTAIL.n20 585
R107 VTAIL.n71 VTAIL.n70 585
R108 VTAIL.n54 VTAIL.n53 585
R109 VTAIL.n65 VTAIL.n64 585
R110 VTAIL.n63 VTAIL.n62 585
R111 VTAIL.n58 VTAIL.n57 585
R112 VTAIL.n47 VTAIL.n46 585
R113 VTAIL.n30 VTAIL.n29 585
R114 VTAIL.n41 VTAIL.n40 585
R115 VTAIL.n39 VTAIL.n38 585
R116 VTAIL.n34 VTAIL.n33 585
R117 VTAIL.n81 VTAIL.t4 330.188
R118 VTAIL.n9 VTAIL.t10 330.188
R119 VTAIL.n59 VTAIL.t8 330.188
R120 VTAIL.n35 VTAIL.t1 330.188
R121 VTAIL.n85 VTAIL.n79 171.744
R122 VTAIL.n86 VTAIL.n85 171.744
R123 VTAIL.n86 VTAIL.n75 171.744
R124 VTAIL.n93 VTAIL.n75 171.744
R125 VTAIL.n13 VTAIL.n7 171.744
R126 VTAIL.n14 VTAIL.n13 171.744
R127 VTAIL.n14 VTAIL.n3 171.744
R128 VTAIL.n21 VTAIL.n3 171.744
R129 VTAIL.n71 VTAIL.n53 171.744
R130 VTAIL.n64 VTAIL.n53 171.744
R131 VTAIL.n64 VTAIL.n63 171.744
R132 VTAIL.n63 VTAIL.n57 171.744
R133 VTAIL.n47 VTAIL.n29 171.744
R134 VTAIL.n40 VTAIL.n29 171.744
R135 VTAIL.n40 VTAIL.n39 171.744
R136 VTAIL.n39 VTAIL.n33 171.744
R137 VTAIL.n51 VTAIL.n50 90.8271
R138 VTAIL.n27 VTAIL.n26 90.8271
R139 VTAIL.n1 VTAIL.n0 90.827
R140 VTAIL.n25 VTAIL.n24 90.827
R141 VTAIL.t4 VTAIL.n79 85.8723
R142 VTAIL.t10 VTAIL.n7 85.8723
R143 VTAIL.t8 VTAIL.n57 85.8723
R144 VTAIL.t1 VTAIL.n33 85.8723
R145 VTAIL.n95 VTAIL.n94 33.9308
R146 VTAIL.n23 VTAIL.n22 33.9308
R147 VTAIL.n73 VTAIL.n72 33.9308
R148 VTAIL.n49 VTAIL.n48 33.9308
R149 VTAIL.n27 VTAIL.n25 17.5134
R150 VTAIL.n95 VTAIL.n73 16.8496
R151 VTAIL.n81 VTAIL.n80 10.7082
R152 VTAIL.n9 VTAIL.n8 10.7082
R153 VTAIL.n59 VTAIL.n58 10.7082
R154 VTAIL.n35 VTAIL.n34 10.7082
R155 VTAIL.n92 VTAIL.n74 10.4732
R156 VTAIL.n20 VTAIL.n2 10.4732
R157 VTAIL.n70 VTAIL.n52 10.4732
R158 VTAIL.n46 VTAIL.n28 10.4732
R159 VTAIL.n91 VTAIL.n76 9.69747
R160 VTAIL.n19 VTAIL.n4 9.69747
R161 VTAIL.n69 VTAIL.n54 9.69747
R162 VTAIL.n45 VTAIL.n30 9.69747
R163 VTAIL.n90 VTAIL.n74 9.45567
R164 VTAIL.n18 VTAIL.n2 9.45567
R165 VTAIL.n68 VTAIL.n52 9.45567
R166 VTAIL.n44 VTAIL.n28 9.45567
R167 VTAIL.n83 VTAIL.n82 9.3005
R168 VTAIL.n78 VTAIL.n77 9.3005
R169 VTAIL.n89 VTAIL.n88 9.3005
R170 VTAIL.n91 VTAIL.n90 9.3005
R171 VTAIL.n11 VTAIL.n10 9.3005
R172 VTAIL.n6 VTAIL.n5 9.3005
R173 VTAIL.n17 VTAIL.n16 9.3005
R174 VTAIL.n19 VTAIL.n18 9.3005
R175 VTAIL.n69 VTAIL.n68 9.3005
R176 VTAIL.n67 VTAIL.n66 9.3005
R177 VTAIL.n56 VTAIL.n55 9.3005
R178 VTAIL.n61 VTAIL.n60 9.3005
R179 VTAIL.n32 VTAIL.n31 9.3005
R180 VTAIL.n43 VTAIL.n42 9.3005
R181 VTAIL.n45 VTAIL.n44 9.3005
R182 VTAIL.n37 VTAIL.n36 9.3005
R183 VTAIL.n88 VTAIL.n87 8.92171
R184 VTAIL.n16 VTAIL.n15 8.92171
R185 VTAIL.n66 VTAIL.n65 8.92171
R186 VTAIL.n42 VTAIL.n41 8.92171
R187 VTAIL.n84 VTAIL.n78 8.14595
R188 VTAIL.n12 VTAIL.n6 8.14595
R189 VTAIL.n62 VTAIL.n56 8.14595
R190 VTAIL.n38 VTAIL.n32 8.14595
R191 VTAIL.n83 VTAIL.n80 7.3702
R192 VTAIL.n11 VTAIL.n8 7.3702
R193 VTAIL.n61 VTAIL.n58 7.3702
R194 VTAIL.n37 VTAIL.n34 7.3702
R195 VTAIL.n0 VTAIL.t0 7.33797
R196 VTAIL.n0 VTAIL.t3 7.33797
R197 VTAIL.n24 VTAIL.t9 7.33797
R198 VTAIL.n24 VTAIL.t7 7.33797
R199 VTAIL.n50 VTAIL.t6 7.33797
R200 VTAIL.n50 VTAIL.t11 7.33797
R201 VTAIL.n26 VTAIL.t2 7.33797
R202 VTAIL.n26 VTAIL.t5 7.33797
R203 VTAIL.n84 VTAIL.n83 5.81868
R204 VTAIL.n12 VTAIL.n11 5.81868
R205 VTAIL.n62 VTAIL.n61 5.81868
R206 VTAIL.n38 VTAIL.n37 5.81868
R207 VTAIL.n87 VTAIL.n78 5.04292
R208 VTAIL.n15 VTAIL.n6 5.04292
R209 VTAIL.n65 VTAIL.n56 5.04292
R210 VTAIL.n41 VTAIL.n32 5.04292
R211 VTAIL.n88 VTAIL.n76 4.26717
R212 VTAIL.n16 VTAIL.n4 4.26717
R213 VTAIL.n66 VTAIL.n54 4.26717
R214 VTAIL.n42 VTAIL.n30 4.26717
R215 VTAIL.n92 VTAIL.n91 3.49141
R216 VTAIL.n20 VTAIL.n19 3.49141
R217 VTAIL.n70 VTAIL.n69 3.49141
R218 VTAIL.n46 VTAIL.n45 3.49141
R219 VTAIL.n94 VTAIL.n74 2.71565
R220 VTAIL.n22 VTAIL.n2 2.71565
R221 VTAIL.n72 VTAIL.n52 2.71565
R222 VTAIL.n48 VTAIL.n28 2.71565
R223 VTAIL.n60 VTAIL.n59 2.42873
R224 VTAIL.n82 VTAIL.n81 2.42873
R225 VTAIL.n10 VTAIL.n9 2.42873
R226 VTAIL.n36 VTAIL.n35 2.42873
R227 VTAIL.n51 VTAIL.n49 0.802224
R228 VTAIL.n23 VTAIL.n1 0.802224
R229 VTAIL.n49 VTAIL.n27 0.664293
R230 VTAIL.n73 VTAIL.n51 0.664293
R231 VTAIL.n25 VTAIL.n23 0.664293
R232 VTAIL VTAIL.n95 0.440155
R233 VTAIL VTAIL.n1 0.224638
R234 VTAIL.n82 VTAIL.n77 0.155672
R235 VTAIL.n89 VTAIL.n77 0.155672
R236 VTAIL.n90 VTAIL.n89 0.155672
R237 VTAIL.n10 VTAIL.n5 0.155672
R238 VTAIL.n17 VTAIL.n5 0.155672
R239 VTAIL.n18 VTAIL.n17 0.155672
R240 VTAIL.n68 VTAIL.n67 0.155672
R241 VTAIL.n67 VTAIL.n55 0.155672
R242 VTAIL.n60 VTAIL.n55 0.155672
R243 VTAIL.n44 VTAIL.n43 0.155672
R244 VTAIL.n43 VTAIL.n31 0.155672
R245 VTAIL.n36 VTAIL.n31 0.155672
R246 B.n244 B.n243 585
R247 B.n245 B.n38 585
R248 B.n247 B.n246 585
R249 B.n248 B.n37 585
R250 B.n250 B.n249 585
R251 B.n251 B.n36 585
R252 B.n253 B.n252 585
R253 B.n254 B.n35 585
R254 B.n256 B.n255 585
R255 B.n257 B.n34 585
R256 B.n259 B.n258 585
R257 B.n260 B.n33 585
R258 B.n262 B.n261 585
R259 B.n263 B.n32 585
R260 B.n265 B.n264 585
R261 B.n266 B.n31 585
R262 B.n268 B.n267 585
R263 B.n269 B.n30 585
R264 B.n271 B.n270 585
R265 B.n273 B.n27 585
R266 B.n275 B.n274 585
R267 B.n276 B.n26 585
R268 B.n278 B.n277 585
R269 B.n279 B.n25 585
R270 B.n281 B.n280 585
R271 B.n282 B.n24 585
R272 B.n284 B.n283 585
R273 B.n285 B.n23 585
R274 B.n287 B.n286 585
R275 B.n289 B.n288 585
R276 B.n290 B.n19 585
R277 B.n292 B.n291 585
R278 B.n293 B.n18 585
R279 B.n295 B.n294 585
R280 B.n296 B.n17 585
R281 B.n298 B.n297 585
R282 B.n299 B.n16 585
R283 B.n301 B.n300 585
R284 B.n302 B.n15 585
R285 B.n304 B.n303 585
R286 B.n305 B.n14 585
R287 B.n307 B.n306 585
R288 B.n308 B.n13 585
R289 B.n310 B.n309 585
R290 B.n311 B.n12 585
R291 B.n313 B.n312 585
R292 B.n314 B.n11 585
R293 B.n316 B.n315 585
R294 B.n242 B.n39 585
R295 B.n241 B.n240 585
R296 B.n239 B.n40 585
R297 B.n238 B.n237 585
R298 B.n236 B.n41 585
R299 B.n235 B.n234 585
R300 B.n233 B.n42 585
R301 B.n232 B.n231 585
R302 B.n230 B.n43 585
R303 B.n229 B.n228 585
R304 B.n227 B.n44 585
R305 B.n226 B.n225 585
R306 B.n224 B.n45 585
R307 B.n223 B.n222 585
R308 B.n221 B.n46 585
R309 B.n220 B.n219 585
R310 B.n218 B.n47 585
R311 B.n217 B.n216 585
R312 B.n215 B.n48 585
R313 B.n214 B.n213 585
R314 B.n212 B.n49 585
R315 B.n211 B.n210 585
R316 B.n209 B.n50 585
R317 B.n208 B.n207 585
R318 B.n206 B.n51 585
R319 B.n205 B.n204 585
R320 B.n203 B.n52 585
R321 B.n202 B.n201 585
R322 B.n200 B.n53 585
R323 B.n199 B.n198 585
R324 B.n197 B.n54 585
R325 B.n196 B.n195 585
R326 B.n194 B.n55 585
R327 B.n193 B.n192 585
R328 B.n191 B.n56 585
R329 B.n118 B.n117 585
R330 B.n119 B.n84 585
R331 B.n121 B.n120 585
R332 B.n122 B.n83 585
R333 B.n124 B.n123 585
R334 B.n125 B.n82 585
R335 B.n127 B.n126 585
R336 B.n128 B.n81 585
R337 B.n130 B.n129 585
R338 B.n131 B.n80 585
R339 B.n133 B.n132 585
R340 B.n134 B.n79 585
R341 B.n136 B.n135 585
R342 B.n137 B.n78 585
R343 B.n139 B.n138 585
R344 B.n140 B.n77 585
R345 B.n142 B.n141 585
R346 B.n143 B.n76 585
R347 B.n145 B.n144 585
R348 B.n147 B.n73 585
R349 B.n149 B.n148 585
R350 B.n150 B.n72 585
R351 B.n152 B.n151 585
R352 B.n153 B.n71 585
R353 B.n155 B.n154 585
R354 B.n156 B.n70 585
R355 B.n158 B.n157 585
R356 B.n159 B.n69 585
R357 B.n161 B.n160 585
R358 B.n163 B.n162 585
R359 B.n164 B.n65 585
R360 B.n166 B.n165 585
R361 B.n167 B.n64 585
R362 B.n169 B.n168 585
R363 B.n170 B.n63 585
R364 B.n172 B.n171 585
R365 B.n173 B.n62 585
R366 B.n175 B.n174 585
R367 B.n176 B.n61 585
R368 B.n178 B.n177 585
R369 B.n179 B.n60 585
R370 B.n181 B.n180 585
R371 B.n182 B.n59 585
R372 B.n184 B.n183 585
R373 B.n185 B.n58 585
R374 B.n187 B.n186 585
R375 B.n188 B.n57 585
R376 B.n190 B.n189 585
R377 B.n116 B.n85 585
R378 B.n115 B.n114 585
R379 B.n113 B.n86 585
R380 B.n112 B.n111 585
R381 B.n110 B.n87 585
R382 B.n109 B.n108 585
R383 B.n107 B.n88 585
R384 B.n106 B.n105 585
R385 B.n104 B.n89 585
R386 B.n103 B.n102 585
R387 B.n101 B.n90 585
R388 B.n100 B.n99 585
R389 B.n98 B.n91 585
R390 B.n97 B.n96 585
R391 B.n95 B.n92 585
R392 B.n94 B.n93 585
R393 B.n2 B.n0 585
R394 B.n341 B.n1 585
R395 B.n340 B.n339 585
R396 B.n338 B.n3 585
R397 B.n337 B.n336 585
R398 B.n335 B.n4 585
R399 B.n334 B.n333 585
R400 B.n332 B.n5 585
R401 B.n331 B.n330 585
R402 B.n329 B.n6 585
R403 B.n328 B.n327 585
R404 B.n326 B.n7 585
R405 B.n325 B.n324 585
R406 B.n323 B.n8 585
R407 B.n322 B.n321 585
R408 B.n320 B.n9 585
R409 B.n319 B.n318 585
R410 B.n317 B.n10 585
R411 B.n343 B.n342 585
R412 B.n118 B.n85 550.159
R413 B.n317 B.n316 550.159
R414 B.n191 B.n190 550.159
R415 B.n244 B.n39 550.159
R416 B.n66 B.t9 450.695
R417 B.n74 B.t0 450.695
R418 B.n20 B.t3 450.695
R419 B.n28 B.t6 450.695
R420 B.n66 B.t11 255.982
R421 B.n28 B.t7 255.982
R422 B.n74 B.t2 255.981
R423 B.n20 B.t4 255.981
R424 B.n67 B.t10 241.048
R425 B.n29 B.t8 241.048
R426 B.n75 B.t1 241.048
R427 B.n21 B.t5 241.048
R428 B.n114 B.n85 163.367
R429 B.n114 B.n113 163.367
R430 B.n113 B.n112 163.367
R431 B.n112 B.n87 163.367
R432 B.n108 B.n87 163.367
R433 B.n108 B.n107 163.367
R434 B.n107 B.n106 163.367
R435 B.n106 B.n89 163.367
R436 B.n102 B.n89 163.367
R437 B.n102 B.n101 163.367
R438 B.n101 B.n100 163.367
R439 B.n100 B.n91 163.367
R440 B.n96 B.n91 163.367
R441 B.n96 B.n95 163.367
R442 B.n95 B.n94 163.367
R443 B.n94 B.n2 163.367
R444 B.n342 B.n2 163.367
R445 B.n342 B.n341 163.367
R446 B.n341 B.n340 163.367
R447 B.n340 B.n3 163.367
R448 B.n336 B.n3 163.367
R449 B.n336 B.n335 163.367
R450 B.n335 B.n334 163.367
R451 B.n334 B.n5 163.367
R452 B.n330 B.n5 163.367
R453 B.n330 B.n329 163.367
R454 B.n329 B.n328 163.367
R455 B.n328 B.n7 163.367
R456 B.n324 B.n7 163.367
R457 B.n324 B.n323 163.367
R458 B.n323 B.n322 163.367
R459 B.n322 B.n9 163.367
R460 B.n318 B.n9 163.367
R461 B.n318 B.n317 163.367
R462 B.n119 B.n118 163.367
R463 B.n120 B.n119 163.367
R464 B.n120 B.n83 163.367
R465 B.n124 B.n83 163.367
R466 B.n125 B.n124 163.367
R467 B.n126 B.n125 163.367
R468 B.n126 B.n81 163.367
R469 B.n130 B.n81 163.367
R470 B.n131 B.n130 163.367
R471 B.n132 B.n131 163.367
R472 B.n132 B.n79 163.367
R473 B.n136 B.n79 163.367
R474 B.n137 B.n136 163.367
R475 B.n138 B.n137 163.367
R476 B.n138 B.n77 163.367
R477 B.n142 B.n77 163.367
R478 B.n143 B.n142 163.367
R479 B.n144 B.n143 163.367
R480 B.n144 B.n73 163.367
R481 B.n149 B.n73 163.367
R482 B.n150 B.n149 163.367
R483 B.n151 B.n150 163.367
R484 B.n151 B.n71 163.367
R485 B.n155 B.n71 163.367
R486 B.n156 B.n155 163.367
R487 B.n157 B.n156 163.367
R488 B.n157 B.n69 163.367
R489 B.n161 B.n69 163.367
R490 B.n162 B.n161 163.367
R491 B.n162 B.n65 163.367
R492 B.n166 B.n65 163.367
R493 B.n167 B.n166 163.367
R494 B.n168 B.n167 163.367
R495 B.n168 B.n63 163.367
R496 B.n172 B.n63 163.367
R497 B.n173 B.n172 163.367
R498 B.n174 B.n173 163.367
R499 B.n174 B.n61 163.367
R500 B.n178 B.n61 163.367
R501 B.n179 B.n178 163.367
R502 B.n180 B.n179 163.367
R503 B.n180 B.n59 163.367
R504 B.n184 B.n59 163.367
R505 B.n185 B.n184 163.367
R506 B.n186 B.n185 163.367
R507 B.n186 B.n57 163.367
R508 B.n190 B.n57 163.367
R509 B.n192 B.n191 163.367
R510 B.n192 B.n55 163.367
R511 B.n196 B.n55 163.367
R512 B.n197 B.n196 163.367
R513 B.n198 B.n197 163.367
R514 B.n198 B.n53 163.367
R515 B.n202 B.n53 163.367
R516 B.n203 B.n202 163.367
R517 B.n204 B.n203 163.367
R518 B.n204 B.n51 163.367
R519 B.n208 B.n51 163.367
R520 B.n209 B.n208 163.367
R521 B.n210 B.n209 163.367
R522 B.n210 B.n49 163.367
R523 B.n214 B.n49 163.367
R524 B.n215 B.n214 163.367
R525 B.n216 B.n215 163.367
R526 B.n216 B.n47 163.367
R527 B.n220 B.n47 163.367
R528 B.n221 B.n220 163.367
R529 B.n222 B.n221 163.367
R530 B.n222 B.n45 163.367
R531 B.n226 B.n45 163.367
R532 B.n227 B.n226 163.367
R533 B.n228 B.n227 163.367
R534 B.n228 B.n43 163.367
R535 B.n232 B.n43 163.367
R536 B.n233 B.n232 163.367
R537 B.n234 B.n233 163.367
R538 B.n234 B.n41 163.367
R539 B.n238 B.n41 163.367
R540 B.n239 B.n238 163.367
R541 B.n240 B.n239 163.367
R542 B.n240 B.n39 163.367
R543 B.n316 B.n11 163.367
R544 B.n312 B.n11 163.367
R545 B.n312 B.n311 163.367
R546 B.n311 B.n310 163.367
R547 B.n310 B.n13 163.367
R548 B.n306 B.n13 163.367
R549 B.n306 B.n305 163.367
R550 B.n305 B.n304 163.367
R551 B.n304 B.n15 163.367
R552 B.n300 B.n15 163.367
R553 B.n300 B.n299 163.367
R554 B.n299 B.n298 163.367
R555 B.n298 B.n17 163.367
R556 B.n294 B.n17 163.367
R557 B.n294 B.n293 163.367
R558 B.n293 B.n292 163.367
R559 B.n292 B.n19 163.367
R560 B.n288 B.n19 163.367
R561 B.n288 B.n287 163.367
R562 B.n287 B.n23 163.367
R563 B.n283 B.n23 163.367
R564 B.n283 B.n282 163.367
R565 B.n282 B.n281 163.367
R566 B.n281 B.n25 163.367
R567 B.n277 B.n25 163.367
R568 B.n277 B.n276 163.367
R569 B.n276 B.n275 163.367
R570 B.n275 B.n27 163.367
R571 B.n270 B.n27 163.367
R572 B.n270 B.n269 163.367
R573 B.n269 B.n268 163.367
R574 B.n268 B.n31 163.367
R575 B.n264 B.n31 163.367
R576 B.n264 B.n263 163.367
R577 B.n263 B.n262 163.367
R578 B.n262 B.n33 163.367
R579 B.n258 B.n33 163.367
R580 B.n258 B.n257 163.367
R581 B.n257 B.n256 163.367
R582 B.n256 B.n35 163.367
R583 B.n252 B.n35 163.367
R584 B.n252 B.n251 163.367
R585 B.n251 B.n250 163.367
R586 B.n250 B.n37 163.367
R587 B.n246 B.n37 163.367
R588 B.n246 B.n245 163.367
R589 B.n245 B.n244 163.367
R590 B.n68 B.n67 59.5399
R591 B.n146 B.n75 59.5399
R592 B.n22 B.n21 59.5399
R593 B.n272 B.n29 59.5399
R594 B.n315 B.n10 35.7468
R595 B.n243 B.n242 35.7468
R596 B.n189 B.n56 35.7468
R597 B.n117 B.n116 35.7468
R598 B B.n343 18.0485
R599 B.n67 B.n66 14.9338
R600 B.n75 B.n74 14.9338
R601 B.n21 B.n20 14.9338
R602 B.n29 B.n28 14.9338
R603 B.n315 B.n314 10.6151
R604 B.n314 B.n313 10.6151
R605 B.n313 B.n12 10.6151
R606 B.n309 B.n12 10.6151
R607 B.n309 B.n308 10.6151
R608 B.n308 B.n307 10.6151
R609 B.n307 B.n14 10.6151
R610 B.n303 B.n14 10.6151
R611 B.n303 B.n302 10.6151
R612 B.n302 B.n301 10.6151
R613 B.n301 B.n16 10.6151
R614 B.n297 B.n16 10.6151
R615 B.n297 B.n296 10.6151
R616 B.n296 B.n295 10.6151
R617 B.n295 B.n18 10.6151
R618 B.n291 B.n18 10.6151
R619 B.n291 B.n290 10.6151
R620 B.n290 B.n289 10.6151
R621 B.n286 B.n285 10.6151
R622 B.n285 B.n284 10.6151
R623 B.n284 B.n24 10.6151
R624 B.n280 B.n24 10.6151
R625 B.n280 B.n279 10.6151
R626 B.n279 B.n278 10.6151
R627 B.n278 B.n26 10.6151
R628 B.n274 B.n26 10.6151
R629 B.n274 B.n273 10.6151
R630 B.n271 B.n30 10.6151
R631 B.n267 B.n30 10.6151
R632 B.n267 B.n266 10.6151
R633 B.n266 B.n265 10.6151
R634 B.n265 B.n32 10.6151
R635 B.n261 B.n32 10.6151
R636 B.n261 B.n260 10.6151
R637 B.n260 B.n259 10.6151
R638 B.n259 B.n34 10.6151
R639 B.n255 B.n34 10.6151
R640 B.n255 B.n254 10.6151
R641 B.n254 B.n253 10.6151
R642 B.n253 B.n36 10.6151
R643 B.n249 B.n36 10.6151
R644 B.n249 B.n248 10.6151
R645 B.n248 B.n247 10.6151
R646 B.n247 B.n38 10.6151
R647 B.n243 B.n38 10.6151
R648 B.n193 B.n56 10.6151
R649 B.n194 B.n193 10.6151
R650 B.n195 B.n194 10.6151
R651 B.n195 B.n54 10.6151
R652 B.n199 B.n54 10.6151
R653 B.n200 B.n199 10.6151
R654 B.n201 B.n200 10.6151
R655 B.n201 B.n52 10.6151
R656 B.n205 B.n52 10.6151
R657 B.n206 B.n205 10.6151
R658 B.n207 B.n206 10.6151
R659 B.n207 B.n50 10.6151
R660 B.n211 B.n50 10.6151
R661 B.n212 B.n211 10.6151
R662 B.n213 B.n212 10.6151
R663 B.n213 B.n48 10.6151
R664 B.n217 B.n48 10.6151
R665 B.n218 B.n217 10.6151
R666 B.n219 B.n218 10.6151
R667 B.n219 B.n46 10.6151
R668 B.n223 B.n46 10.6151
R669 B.n224 B.n223 10.6151
R670 B.n225 B.n224 10.6151
R671 B.n225 B.n44 10.6151
R672 B.n229 B.n44 10.6151
R673 B.n230 B.n229 10.6151
R674 B.n231 B.n230 10.6151
R675 B.n231 B.n42 10.6151
R676 B.n235 B.n42 10.6151
R677 B.n236 B.n235 10.6151
R678 B.n237 B.n236 10.6151
R679 B.n237 B.n40 10.6151
R680 B.n241 B.n40 10.6151
R681 B.n242 B.n241 10.6151
R682 B.n117 B.n84 10.6151
R683 B.n121 B.n84 10.6151
R684 B.n122 B.n121 10.6151
R685 B.n123 B.n122 10.6151
R686 B.n123 B.n82 10.6151
R687 B.n127 B.n82 10.6151
R688 B.n128 B.n127 10.6151
R689 B.n129 B.n128 10.6151
R690 B.n129 B.n80 10.6151
R691 B.n133 B.n80 10.6151
R692 B.n134 B.n133 10.6151
R693 B.n135 B.n134 10.6151
R694 B.n135 B.n78 10.6151
R695 B.n139 B.n78 10.6151
R696 B.n140 B.n139 10.6151
R697 B.n141 B.n140 10.6151
R698 B.n141 B.n76 10.6151
R699 B.n145 B.n76 10.6151
R700 B.n148 B.n147 10.6151
R701 B.n148 B.n72 10.6151
R702 B.n152 B.n72 10.6151
R703 B.n153 B.n152 10.6151
R704 B.n154 B.n153 10.6151
R705 B.n154 B.n70 10.6151
R706 B.n158 B.n70 10.6151
R707 B.n159 B.n158 10.6151
R708 B.n160 B.n159 10.6151
R709 B.n164 B.n163 10.6151
R710 B.n165 B.n164 10.6151
R711 B.n165 B.n64 10.6151
R712 B.n169 B.n64 10.6151
R713 B.n170 B.n169 10.6151
R714 B.n171 B.n170 10.6151
R715 B.n171 B.n62 10.6151
R716 B.n175 B.n62 10.6151
R717 B.n176 B.n175 10.6151
R718 B.n177 B.n176 10.6151
R719 B.n177 B.n60 10.6151
R720 B.n181 B.n60 10.6151
R721 B.n182 B.n181 10.6151
R722 B.n183 B.n182 10.6151
R723 B.n183 B.n58 10.6151
R724 B.n187 B.n58 10.6151
R725 B.n188 B.n187 10.6151
R726 B.n189 B.n188 10.6151
R727 B.n116 B.n115 10.6151
R728 B.n115 B.n86 10.6151
R729 B.n111 B.n86 10.6151
R730 B.n111 B.n110 10.6151
R731 B.n110 B.n109 10.6151
R732 B.n109 B.n88 10.6151
R733 B.n105 B.n88 10.6151
R734 B.n105 B.n104 10.6151
R735 B.n104 B.n103 10.6151
R736 B.n103 B.n90 10.6151
R737 B.n99 B.n90 10.6151
R738 B.n99 B.n98 10.6151
R739 B.n98 B.n97 10.6151
R740 B.n97 B.n92 10.6151
R741 B.n93 B.n92 10.6151
R742 B.n93 B.n0 10.6151
R743 B.n339 B.n1 10.6151
R744 B.n339 B.n338 10.6151
R745 B.n338 B.n337 10.6151
R746 B.n337 B.n4 10.6151
R747 B.n333 B.n4 10.6151
R748 B.n333 B.n332 10.6151
R749 B.n332 B.n331 10.6151
R750 B.n331 B.n6 10.6151
R751 B.n327 B.n6 10.6151
R752 B.n327 B.n326 10.6151
R753 B.n326 B.n325 10.6151
R754 B.n325 B.n8 10.6151
R755 B.n321 B.n8 10.6151
R756 B.n321 B.n320 10.6151
R757 B.n320 B.n319 10.6151
R758 B.n319 B.n10 10.6151
R759 B.n289 B.n22 9.36635
R760 B.n272 B.n271 9.36635
R761 B.n146 B.n145 9.36635
R762 B.n163 B.n68 9.36635
R763 B.n343 B.n0 2.81026
R764 B.n343 B.n1 2.81026
R765 B.n286 B.n22 1.24928
R766 B.n273 B.n272 1.24928
R767 B.n147 B.n146 1.24928
R768 B.n160 B.n68 1.24928
R769 VN.n0 VN.t1 357.935
R770 VN.n4 VN.t0 357.935
R771 VN.n2 VN.t3 339.774
R772 VN.n6 VN.t5 339.774
R773 VN.n1 VN.t4 332.471
R774 VN.n5 VN.t2 332.471
R775 VN.n3 VN.n2 161.3
R776 VN.n7 VN.n6 161.3
R777 VN.n7 VN.n4 71.8132
R778 VN.n3 VN.n0 71.8132
R779 VN.n2 VN.n1 40.8975
R780 VN.n6 VN.n5 40.8975
R781 VN VN.n7 34.9456
R782 VN.n5 VN.n4 18.1394
R783 VN.n1 VN.n0 18.1394
R784 VN VN.n3 0.0516364
R785 VDD2.n43 VDD2.n42 756.745
R786 VDD2.n20 VDD2.n19 756.745
R787 VDD2.n42 VDD2.n41 585
R788 VDD2.n25 VDD2.n24 585
R789 VDD2.n36 VDD2.n35 585
R790 VDD2.n34 VDD2.n33 585
R791 VDD2.n29 VDD2.n28 585
R792 VDD2.n6 VDD2.n5 585
R793 VDD2.n11 VDD2.n10 585
R794 VDD2.n13 VDD2.n12 585
R795 VDD2.n2 VDD2.n1 585
R796 VDD2.n19 VDD2.n18 585
R797 VDD2.n7 VDD2.t4 330.188
R798 VDD2.n30 VDD2.t0 330.188
R799 VDD2.n42 VDD2.n24 171.744
R800 VDD2.n35 VDD2.n24 171.744
R801 VDD2.n35 VDD2.n34 171.744
R802 VDD2.n34 VDD2.n28 171.744
R803 VDD2.n11 VDD2.n5 171.744
R804 VDD2.n12 VDD2.n11 171.744
R805 VDD2.n12 VDD2.n1 171.744
R806 VDD2.n19 VDD2.n1 171.744
R807 VDD2.n22 VDD2.n21 107.617
R808 VDD2 VDD2.n45 107.612
R809 VDD2.t0 VDD2.n28 85.8723
R810 VDD2.t4 VDD2.n5 85.8723
R811 VDD2.n22 VDD2.n20 51.0521
R812 VDD2.n44 VDD2.n43 50.6096
R813 VDD2.n44 VDD2.n22 29.6916
R814 VDD2.n30 VDD2.n29 10.7082
R815 VDD2.n7 VDD2.n6 10.7082
R816 VDD2.n41 VDD2.n23 10.4732
R817 VDD2.n18 VDD2.n0 10.4732
R818 VDD2.n40 VDD2.n25 9.69747
R819 VDD2.n17 VDD2.n2 9.69747
R820 VDD2.n39 VDD2.n23 9.45567
R821 VDD2.n16 VDD2.n0 9.45567
R822 VDD2.n27 VDD2.n26 9.3005
R823 VDD2.n38 VDD2.n37 9.3005
R824 VDD2.n40 VDD2.n39 9.3005
R825 VDD2.n32 VDD2.n31 9.3005
R826 VDD2.n9 VDD2.n8 9.3005
R827 VDD2.n4 VDD2.n3 9.3005
R828 VDD2.n15 VDD2.n14 9.3005
R829 VDD2.n17 VDD2.n16 9.3005
R830 VDD2.n37 VDD2.n36 8.92171
R831 VDD2.n14 VDD2.n13 8.92171
R832 VDD2.n33 VDD2.n27 8.14595
R833 VDD2.n10 VDD2.n4 8.14595
R834 VDD2.n32 VDD2.n29 7.3702
R835 VDD2.n9 VDD2.n6 7.3702
R836 VDD2.n45 VDD2.t3 7.33797
R837 VDD2.n45 VDD2.t5 7.33797
R838 VDD2.n21 VDD2.t1 7.33797
R839 VDD2.n21 VDD2.t2 7.33797
R840 VDD2.n33 VDD2.n32 5.81868
R841 VDD2.n10 VDD2.n9 5.81868
R842 VDD2.n36 VDD2.n27 5.04292
R843 VDD2.n13 VDD2.n4 5.04292
R844 VDD2.n37 VDD2.n25 4.26717
R845 VDD2.n14 VDD2.n2 4.26717
R846 VDD2.n41 VDD2.n40 3.49141
R847 VDD2.n18 VDD2.n17 3.49141
R848 VDD2.n43 VDD2.n23 2.71565
R849 VDD2.n20 VDD2.n0 2.71565
R850 VDD2.n31 VDD2.n30 2.42873
R851 VDD2.n8 VDD2.n7 2.42873
R852 VDD2 VDD2.n44 0.556535
R853 VDD2.n39 VDD2.n38 0.155672
R854 VDD2.n38 VDD2.n26 0.155672
R855 VDD2.n31 VDD2.n26 0.155672
R856 VDD2.n8 VDD2.n3 0.155672
R857 VDD2.n15 VDD2.n3 0.155672
R858 VDD2.n16 VDD2.n15 0.155672
C0 VP w_n1586_n1854# 2.52467f
C1 VDD1 VTAIL 5.46742f
C2 VDD1 B 0.938441f
C3 VN VTAIL 1.41836f
C4 VN B 0.618198f
C5 VDD2 VDD1 0.615841f
C6 VP VTAIL 1.43269f
C7 VDD2 VN 1.45255f
C8 w_n1586_n1854# VTAIL 1.71195f
C9 VP B 0.939502f
C10 w_n1586_n1854# B 4.5709f
C11 VP VDD2 0.278747f
C12 VDD2 w_n1586_n1854# 1.18497f
C13 VTAIL B 1.24242f
C14 VDD2 VTAIL 5.50352f
C15 VDD2 B 0.96156f
C16 VN VDD1 0.151789f
C17 VP VDD1 1.57721f
C18 VDD1 w_n1586_n1854# 1.16911f
C19 VP VN 3.42901f
C20 VN w_n1586_n1854# 2.32596f
C21 VDD2 VSUBS 0.829328f
C22 VDD1 VSUBS 0.768237f
C23 VTAIL VSUBS 0.340681f
C24 VN VSUBS 2.97085f
C25 VP VSUBS 0.905321f
C26 B VSUBS 1.773754f
C27 w_n1586_n1854# VSUBS 36.9411f
C28 VDD2.n0 VSUBS 0.011219f
C29 VDD2.n1 VSUBS 0.025242f
C30 VDD2.n2 VSUBS 0.011308f
C31 VDD2.n3 VSUBS 0.019874f
C32 VDD2.n4 VSUBS 0.01068f
C33 VDD2.n5 VSUBS 0.018932f
C34 VDD2.n6 VSUBS 0.018922f
C35 VDD2.t4 VSUBS 0.054833f
C36 VDD2.n7 VSUBS 0.08924f
C37 VDD2.n8 VSUBS 0.315649f
C38 VDD2.n9 VSUBS 0.01068f
C39 VDD2.n10 VSUBS 0.011308f
C40 VDD2.n11 VSUBS 0.025242f
C41 VDD2.n12 VSUBS 0.025242f
C42 VDD2.n13 VSUBS 0.011308f
C43 VDD2.n14 VSUBS 0.01068f
C44 VDD2.n15 VSUBS 0.019874f
C45 VDD2.n16 VSUBS 0.052182f
C46 VDD2.n17 VSUBS 0.01068f
C47 VDD2.n18 VSUBS 0.011308f
C48 VDD2.n19 VSUBS 0.0548f
C49 VDD2.n20 VSUBS 0.052055f
C50 VDD2.t1 VSUBS 0.069574f
C51 VDD2.t2 VSUBS 0.069574f
C52 VDD2.n21 VSUBS 0.43348f
C53 VDD2.n22 VSUBS 1.14619f
C54 VDD2.n23 VSUBS 0.011219f
C55 VDD2.n24 VSUBS 0.025242f
C56 VDD2.n25 VSUBS 0.011308f
C57 VDD2.n26 VSUBS 0.019874f
C58 VDD2.n27 VSUBS 0.01068f
C59 VDD2.n28 VSUBS 0.018932f
C60 VDD2.n29 VSUBS 0.018922f
C61 VDD2.t0 VSUBS 0.054833f
C62 VDD2.n30 VSUBS 0.08924f
C63 VDD2.n31 VSUBS 0.315649f
C64 VDD2.n32 VSUBS 0.01068f
C65 VDD2.n33 VSUBS 0.011308f
C66 VDD2.n34 VSUBS 0.025242f
C67 VDD2.n35 VSUBS 0.025242f
C68 VDD2.n36 VSUBS 0.011308f
C69 VDD2.n37 VSUBS 0.01068f
C70 VDD2.n38 VSUBS 0.019874f
C71 VDD2.n39 VSUBS 0.052182f
C72 VDD2.n40 VSUBS 0.01068f
C73 VDD2.n41 VSUBS 0.011308f
C74 VDD2.n42 VSUBS 0.0548f
C75 VDD2.n43 VSUBS 0.051456f
C76 VDD2.n44 VSUBS 1.08762f
C77 VDD2.t3 VSUBS 0.069574f
C78 VDD2.t5 VSUBS 0.069574f
C79 VDD2.n45 VSUBS 0.433466f
C80 VN.t1 VSUBS 0.286936f
C81 VN.n0 VSUBS 0.136356f
C82 VN.t4 VSUBS 0.276758f
C83 VN.n1 VSUBS 0.151533f
C84 VN.t3 VSUBS 0.279664f
C85 VN.n2 VSUBS 0.143263f
C86 VN.n3 VSUBS 0.148071f
C87 VN.t0 VSUBS 0.286936f
C88 VN.n4 VSUBS 0.136356f
C89 VN.t5 VSUBS 0.279664f
C90 VN.t2 VSUBS 0.276758f
C91 VN.n5 VSUBS 0.151533f
C92 VN.n6 VSUBS 0.143263f
C93 VN.n7 VSUBS 1.54854f
C94 B.n0 VSUBS 0.004633f
C95 B.n1 VSUBS 0.004633f
C96 B.n2 VSUBS 0.007327f
C97 B.n3 VSUBS 0.007327f
C98 B.n4 VSUBS 0.007327f
C99 B.n5 VSUBS 0.007327f
C100 B.n6 VSUBS 0.007327f
C101 B.n7 VSUBS 0.007327f
C102 B.n8 VSUBS 0.007327f
C103 B.n9 VSUBS 0.007327f
C104 B.n10 VSUBS 0.017815f
C105 B.n11 VSUBS 0.007327f
C106 B.n12 VSUBS 0.007327f
C107 B.n13 VSUBS 0.007327f
C108 B.n14 VSUBS 0.007327f
C109 B.n15 VSUBS 0.007327f
C110 B.n16 VSUBS 0.007327f
C111 B.n17 VSUBS 0.007327f
C112 B.n18 VSUBS 0.007327f
C113 B.n19 VSUBS 0.007327f
C114 B.t5 VSUBS 0.066486f
C115 B.t4 VSUBS 0.073003f
C116 B.t3 VSUBS 0.087384f
C117 B.n20 VSUBS 0.132664f
C118 B.n21 VSUBS 0.12216f
C119 B.n22 VSUBS 0.016977f
C120 B.n23 VSUBS 0.007327f
C121 B.n24 VSUBS 0.007327f
C122 B.n25 VSUBS 0.007327f
C123 B.n26 VSUBS 0.007327f
C124 B.n27 VSUBS 0.007327f
C125 B.t8 VSUBS 0.066487f
C126 B.t7 VSUBS 0.073004f
C127 B.t6 VSUBS 0.087384f
C128 B.n28 VSUBS 0.132663f
C129 B.n29 VSUBS 0.122158f
C130 B.n30 VSUBS 0.007327f
C131 B.n31 VSUBS 0.007327f
C132 B.n32 VSUBS 0.007327f
C133 B.n33 VSUBS 0.007327f
C134 B.n34 VSUBS 0.007327f
C135 B.n35 VSUBS 0.007327f
C136 B.n36 VSUBS 0.007327f
C137 B.n37 VSUBS 0.007327f
C138 B.n38 VSUBS 0.007327f
C139 B.n39 VSUBS 0.017815f
C140 B.n40 VSUBS 0.007327f
C141 B.n41 VSUBS 0.007327f
C142 B.n42 VSUBS 0.007327f
C143 B.n43 VSUBS 0.007327f
C144 B.n44 VSUBS 0.007327f
C145 B.n45 VSUBS 0.007327f
C146 B.n46 VSUBS 0.007327f
C147 B.n47 VSUBS 0.007327f
C148 B.n48 VSUBS 0.007327f
C149 B.n49 VSUBS 0.007327f
C150 B.n50 VSUBS 0.007327f
C151 B.n51 VSUBS 0.007327f
C152 B.n52 VSUBS 0.007327f
C153 B.n53 VSUBS 0.007327f
C154 B.n54 VSUBS 0.007327f
C155 B.n55 VSUBS 0.007327f
C156 B.n56 VSUBS 0.017815f
C157 B.n57 VSUBS 0.007327f
C158 B.n58 VSUBS 0.007327f
C159 B.n59 VSUBS 0.007327f
C160 B.n60 VSUBS 0.007327f
C161 B.n61 VSUBS 0.007327f
C162 B.n62 VSUBS 0.007327f
C163 B.n63 VSUBS 0.007327f
C164 B.n64 VSUBS 0.007327f
C165 B.n65 VSUBS 0.007327f
C166 B.t10 VSUBS 0.066487f
C167 B.t11 VSUBS 0.073004f
C168 B.t9 VSUBS 0.087384f
C169 B.n66 VSUBS 0.132663f
C170 B.n67 VSUBS 0.122158f
C171 B.n68 VSUBS 0.016977f
C172 B.n69 VSUBS 0.007327f
C173 B.n70 VSUBS 0.007327f
C174 B.n71 VSUBS 0.007327f
C175 B.n72 VSUBS 0.007327f
C176 B.n73 VSUBS 0.007327f
C177 B.t1 VSUBS 0.066486f
C178 B.t2 VSUBS 0.073003f
C179 B.t0 VSUBS 0.087384f
C180 B.n74 VSUBS 0.132664f
C181 B.n75 VSUBS 0.12216f
C182 B.n76 VSUBS 0.007327f
C183 B.n77 VSUBS 0.007327f
C184 B.n78 VSUBS 0.007327f
C185 B.n79 VSUBS 0.007327f
C186 B.n80 VSUBS 0.007327f
C187 B.n81 VSUBS 0.007327f
C188 B.n82 VSUBS 0.007327f
C189 B.n83 VSUBS 0.007327f
C190 B.n84 VSUBS 0.007327f
C191 B.n85 VSUBS 0.017815f
C192 B.n86 VSUBS 0.007327f
C193 B.n87 VSUBS 0.007327f
C194 B.n88 VSUBS 0.007327f
C195 B.n89 VSUBS 0.007327f
C196 B.n90 VSUBS 0.007327f
C197 B.n91 VSUBS 0.007327f
C198 B.n92 VSUBS 0.007327f
C199 B.n93 VSUBS 0.007327f
C200 B.n94 VSUBS 0.007327f
C201 B.n95 VSUBS 0.007327f
C202 B.n96 VSUBS 0.007327f
C203 B.n97 VSUBS 0.007327f
C204 B.n98 VSUBS 0.007327f
C205 B.n99 VSUBS 0.007327f
C206 B.n100 VSUBS 0.007327f
C207 B.n101 VSUBS 0.007327f
C208 B.n102 VSUBS 0.007327f
C209 B.n103 VSUBS 0.007327f
C210 B.n104 VSUBS 0.007327f
C211 B.n105 VSUBS 0.007327f
C212 B.n106 VSUBS 0.007327f
C213 B.n107 VSUBS 0.007327f
C214 B.n108 VSUBS 0.007327f
C215 B.n109 VSUBS 0.007327f
C216 B.n110 VSUBS 0.007327f
C217 B.n111 VSUBS 0.007327f
C218 B.n112 VSUBS 0.007327f
C219 B.n113 VSUBS 0.007327f
C220 B.n114 VSUBS 0.007327f
C221 B.n115 VSUBS 0.007327f
C222 B.n116 VSUBS 0.017815f
C223 B.n117 VSUBS 0.018606f
C224 B.n118 VSUBS 0.018606f
C225 B.n119 VSUBS 0.007327f
C226 B.n120 VSUBS 0.007327f
C227 B.n121 VSUBS 0.007327f
C228 B.n122 VSUBS 0.007327f
C229 B.n123 VSUBS 0.007327f
C230 B.n124 VSUBS 0.007327f
C231 B.n125 VSUBS 0.007327f
C232 B.n126 VSUBS 0.007327f
C233 B.n127 VSUBS 0.007327f
C234 B.n128 VSUBS 0.007327f
C235 B.n129 VSUBS 0.007327f
C236 B.n130 VSUBS 0.007327f
C237 B.n131 VSUBS 0.007327f
C238 B.n132 VSUBS 0.007327f
C239 B.n133 VSUBS 0.007327f
C240 B.n134 VSUBS 0.007327f
C241 B.n135 VSUBS 0.007327f
C242 B.n136 VSUBS 0.007327f
C243 B.n137 VSUBS 0.007327f
C244 B.n138 VSUBS 0.007327f
C245 B.n139 VSUBS 0.007327f
C246 B.n140 VSUBS 0.007327f
C247 B.n141 VSUBS 0.007327f
C248 B.n142 VSUBS 0.007327f
C249 B.n143 VSUBS 0.007327f
C250 B.n144 VSUBS 0.007327f
C251 B.n145 VSUBS 0.006896f
C252 B.n146 VSUBS 0.016977f
C253 B.n147 VSUBS 0.004095f
C254 B.n148 VSUBS 0.007327f
C255 B.n149 VSUBS 0.007327f
C256 B.n150 VSUBS 0.007327f
C257 B.n151 VSUBS 0.007327f
C258 B.n152 VSUBS 0.007327f
C259 B.n153 VSUBS 0.007327f
C260 B.n154 VSUBS 0.007327f
C261 B.n155 VSUBS 0.007327f
C262 B.n156 VSUBS 0.007327f
C263 B.n157 VSUBS 0.007327f
C264 B.n158 VSUBS 0.007327f
C265 B.n159 VSUBS 0.007327f
C266 B.n160 VSUBS 0.004095f
C267 B.n161 VSUBS 0.007327f
C268 B.n162 VSUBS 0.007327f
C269 B.n163 VSUBS 0.006896f
C270 B.n164 VSUBS 0.007327f
C271 B.n165 VSUBS 0.007327f
C272 B.n166 VSUBS 0.007327f
C273 B.n167 VSUBS 0.007327f
C274 B.n168 VSUBS 0.007327f
C275 B.n169 VSUBS 0.007327f
C276 B.n170 VSUBS 0.007327f
C277 B.n171 VSUBS 0.007327f
C278 B.n172 VSUBS 0.007327f
C279 B.n173 VSUBS 0.007327f
C280 B.n174 VSUBS 0.007327f
C281 B.n175 VSUBS 0.007327f
C282 B.n176 VSUBS 0.007327f
C283 B.n177 VSUBS 0.007327f
C284 B.n178 VSUBS 0.007327f
C285 B.n179 VSUBS 0.007327f
C286 B.n180 VSUBS 0.007327f
C287 B.n181 VSUBS 0.007327f
C288 B.n182 VSUBS 0.007327f
C289 B.n183 VSUBS 0.007327f
C290 B.n184 VSUBS 0.007327f
C291 B.n185 VSUBS 0.007327f
C292 B.n186 VSUBS 0.007327f
C293 B.n187 VSUBS 0.007327f
C294 B.n188 VSUBS 0.007327f
C295 B.n189 VSUBS 0.018606f
C296 B.n190 VSUBS 0.018606f
C297 B.n191 VSUBS 0.017815f
C298 B.n192 VSUBS 0.007327f
C299 B.n193 VSUBS 0.007327f
C300 B.n194 VSUBS 0.007327f
C301 B.n195 VSUBS 0.007327f
C302 B.n196 VSUBS 0.007327f
C303 B.n197 VSUBS 0.007327f
C304 B.n198 VSUBS 0.007327f
C305 B.n199 VSUBS 0.007327f
C306 B.n200 VSUBS 0.007327f
C307 B.n201 VSUBS 0.007327f
C308 B.n202 VSUBS 0.007327f
C309 B.n203 VSUBS 0.007327f
C310 B.n204 VSUBS 0.007327f
C311 B.n205 VSUBS 0.007327f
C312 B.n206 VSUBS 0.007327f
C313 B.n207 VSUBS 0.007327f
C314 B.n208 VSUBS 0.007327f
C315 B.n209 VSUBS 0.007327f
C316 B.n210 VSUBS 0.007327f
C317 B.n211 VSUBS 0.007327f
C318 B.n212 VSUBS 0.007327f
C319 B.n213 VSUBS 0.007327f
C320 B.n214 VSUBS 0.007327f
C321 B.n215 VSUBS 0.007327f
C322 B.n216 VSUBS 0.007327f
C323 B.n217 VSUBS 0.007327f
C324 B.n218 VSUBS 0.007327f
C325 B.n219 VSUBS 0.007327f
C326 B.n220 VSUBS 0.007327f
C327 B.n221 VSUBS 0.007327f
C328 B.n222 VSUBS 0.007327f
C329 B.n223 VSUBS 0.007327f
C330 B.n224 VSUBS 0.007327f
C331 B.n225 VSUBS 0.007327f
C332 B.n226 VSUBS 0.007327f
C333 B.n227 VSUBS 0.007327f
C334 B.n228 VSUBS 0.007327f
C335 B.n229 VSUBS 0.007327f
C336 B.n230 VSUBS 0.007327f
C337 B.n231 VSUBS 0.007327f
C338 B.n232 VSUBS 0.007327f
C339 B.n233 VSUBS 0.007327f
C340 B.n234 VSUBS 0.007327f
C341 B.n235 VSUBS 0.007327f
C342 B.n236 VSUBS 0.007327f
C343 B.n237 VSUBS 0.007327f
C344 B.n238 VSUBS 0.007327f
C345 B.n239 VSUBS 0.007327f
C346 B.n240 VSUBS 0.007327f
C347 B.n241 VSUBS 0.007327f
C348 B.n242 VSUBS 0.018606f
C349 B.n243 VSUBS 0.017815f
C350 B.n244 VSUBS 0.018606f
C351 B.n245 VSUBS 0.007327f
C352 B.n246 VSUBS 0.007327f
C353 B.n247 VSUBS 0.007327f
C354 B.n248 VSUBS 0.007327f
C355 B.n249 VSUBS 0.007327f
C356 B.n250 VSUBS 0.007327f
C357 B.n251 VSUBS 0.007327f
C358 B.n252 VSUBS 0.007327f
C359 B.n253 VSUBS 0.007327f
C360 B.n254 VSUBS 0.007327f
C361 B.n255 VSUBS 0.007327f
C362 B.n256 VSUBS 0.007327f
C363 B.n257 VSUBS 0.007327f
C364 B.n258 VSUBS 0.007327f
C365 B.n259 VSUBS 0.007327f
C366 B.n260 VSUBS 0.007327f
C367 B.n261 VSUBS 0.007327f
C368 B.n262 VSUBS 0.007327f
C369 B.n263 VSUBS 0.007327f
C370 B.n264 VSUBS 0.007327f
C371 B.n265 VSUBS 0.007327f
C372 B.n266 VSUBS 0.007327f
C373 B.n267 VSUBS 0.007327f
C374 B.n268 VSUBS 0.007327f
C375 B.n269 VSUBS 0.007327f
C376 B.n270 VSUBS 0.007327f
C377 B.n271 VSUBS 0.006896f
C378 B.n272 VSUBS 0.016977f
C379 B.n273 VSUBS 0.004095f
C380 B.n274 VSUBS 0.007327f
C381 B.n275 VSUBS 0.007327f
C382 B.n276 VSUBS 0.007327f
C383 B.n277 VSUBS 0.007327f
C384 B.n278 VSUBS 0.007327f
C385 B.n279 VSUBS 0.007327f
C386 B.n280 VSUBS 0.007327f
C387 B.n281 VSUBS 0.007327f
C388 B.n282 VSUBS 0.007327f
C389 B.n283 VSUBS 0.007327f
C390 B.n284 VSUBS 0.007327f
C391 B.n285 VSUBS 0.007327f
C392 B.n286 VSUBS 0.004095f
C393 B.n287 VSUBS 0.007327f
C394 B.n288 VSUBS 0.007327f
C395 B.n289 VSUBS 0.006896f
C396 B.n290 VSUBS 0.007327f
C397 B.n291 VSUBS 0.007327f
C398 B.n292 VSUBS 0.007327f
C399 B.n293 VSUBS 0.007327f
C400 B.n294 VSUBS 0.007327f
C401 B.n295 VSUBS 0.007327f
C402 B.n296 VSUBS 0.007327f
C403 B.n297 VSUBS 0.007327f
C404 B.n298 VSUBS 0.007327f
C405 B.n299 VSUBS 0.007327f
C406 B.n300 VSUBS 0.007327f
C407 B.n301 VSUBS 0.007327f
C408 B.n302 VSUBS 0.007327f
C409 B.n303 VSUBS 0.007327f
C410 B.n304 VSUBS 0.007327f
C411 B.n305 VSUBS 0.007327f
C412 B.n306 VSUBS 0.007327f
C413 B.n307 VSUBS 0.007327f
C414 B.n308 VSUBS 0.007327f
C415 B.n309 VSUBS 0.007327f
C416 B.n310 VSUBS 0.007327f
C417 B.n311 VSUBS 0.007327f
C418 B.n312 VSUBS 0.007327f
C419 B.n313 VSUBS 0.007327f
C420 B.n314 VSUBS 0.007327f
C421 B.n315 VSUBS 0.018606f
C422 B.n316 VSUBS 0.018606f
C423 B.n317 VSUBS 0.017815f
C424 B.n318 VSUBS 0.007327f
C425 B.n319 VSUBS 0.007327f
C426 B.n320 VSUBS 0.007327f
C427 B.n321 VSUBS 0.007327f
C428 B.n322 VSUBS 0.007327f
C429 B.n323 VSUBS 0.007327f
C430 B.n324 VSUBS 0.007327f
C431 B.n325 VSUBS 0.007327f
C432 B.n326 VSUBS 0.007327f
C433 B.n327 VSUBS 0.007327f
C434 B.n328 VSUBS 0.007327f
C435 B.n329 VSUBS 0.007327f
C436 B.n330 VSUBS 0.007327f
C437 B.n331 VSUBS 0.007327f
C438 B.n332 VSUBS 0.007327f
C439 B.n333 VSUBS 0.007327f
C440 B.n334 VSUBS 0.007327f
C441 B.n335 VSUBS 0.007327f
C442 B.n336 VSUBS 0.007327f
C443 B.n337 VSUBS 0.007327f
C444 B.n338 VSUBS 0.007327f
C445 B.n339 VSUBS 0.007327f
C446 B.n340 VSUBS 0.007327f
C447 B.n341 VSUBS 0.007327f
C448 B.n342 VSUBS 0.007327f
C449 B.n343 VSUBS 0.016592f
C450 VTAIL.t0 VSUBS 0.079236f
C451 VTAIL.t3 VSUBS 0.079236f
C452 VTAIL.n0 VSUBS 0.435629f
C453 VTAIL.n1 VSUBS 0.419957f
C454 VTAIL.n2 VSUBS 0.012776f
C455 VTAIL.n3 VSUBS 0.028748f
C456 VTAIL.n4 VSUBS 0.012878f
C457 VTAIL.n5 VSUBS 0.022634f
C458 VTAIL.n6 VSUBS 0.012163f
C459 VTAIL.n7 VSUBS 0.021561f
C460 VTAIL.n8 VSUBS 0.02155f
C461 VTAIL.t10 VSUBS 0.062448f
C462 VTAIL.n9 VSUBS 0.101633f
C463 VTAIL.n10 VSUBS 0.359485f
C464 VTAIL.n11 VSUBS 0.012163f
C465 VTAIL.n12 VSUBS 0.012878f
C466 VTAIL.n13 VSUBS 0.028748f
C467 VTAIL.n14 VSUBS 0.028748f
C468 VTAIL.n15 VSUBS 0.012878f
C469 VTAIL.n16 VSUBS 0.012163f
C470 VTAIL.n17 VSUBS 0.022634f
C471 VTAIL.n18 VSUBS 0.059429f
C472 VTAIL.n19 VSUBS 0.012163f
C473 VTAIL.n20 VSUBS 0.012878f
C474 VTAIL.n21 VSUBS 0.06241f
C475 VTAIL.n22 VSUBS 0.042995f
C476 VTAIL.n23 VSUBS 0.127787f
C477 VTAIL.t9 VSUBS 0.079236f
C478 VTAIL.t7 VSUBS 0.079236f
C479 VTAIL.n24 VSUBS 0.435629f
C480 VTAIL.n25 VSUBS 1.07636f
C481 VTAIL.t2 VSUBS 0.079236f
C482 VTAIL.t5 VSUBS 0.079236f
C483 VTAIL.n26 VSUBS 0.435632f
C484 VTAIL.n27 VSUBS 1.07635f
C485 VTAIL.n28 VSUBS 0.012776f
C486 VTAIL.n29 VSUBS 0.028748f
C487 VTAIL.n30 VSUBS 0.012878f
C488 VTAIL.n31 VSUBS 0.022634f
C489 VTAIL.n32 VSUBS 0.012163f
C490 VTAIL.n33 VSUBS 0.021561f
C491 VTAIL.n34 VSUBS 0.02155f
C492 VTAIL.t1 VSUBS 0.062448f
C493 VTAIL.n35 VSUBS 0.101633f
C494 VTAIL.n36 VSUBS 0.359485f
C495 VTAIL.n37 VSUBS 0.012163f
C496 VTAIL.n38 VSUBS 0.012878f
C497 VTAIL.n39 VSUBS 0.028748f
C498 VTAIL.n40 VSUBS 0.028748f
C499 VTAIL.n41 VSUBS 0.012878f
C500 VTAIL.n42 VSUBS 0.012163f
C501 VTAIL.n43 VSUBS 0.022634f
C502 VTAIL.n44 VSUBS 0.059429f
C503 VTAIL.n45 VSUBS 0.012163f
C504 VTAIL.n46 VSUBS 0.012878f
C505 VTAIL.n47 VSUBS 0.06241f
C506 VTAIL.n48 VSUBS 0.042995f
C507 VTAIL.n49 VSUBS 0.127787f
C508 VTAIL.t6 VSUBS 0.079236f
C509 VTAIL.t11 VSUBS 0.079236f
C510 VTAIL.n50 VSUBS 0.435632f
C511 VTAIL.n51 VSUBS 0.45202f
C512 VTAIL.n52 VSUBS 0.012776f
C513 VTAIL.n53 VSUBS 0.028748f
C514 VTAIL.n54 VSUBS 0.012878f
C515 VTAIL.n55 VSUBS 0.022634f
C516 VTAIL.n56 VSUBS 0.012163f
C517 VTAIL.n57 VSUBS 0.021561f
C518 VTAIL.n58 VSUBS 0.02155f
C519 VTAIL.t8 VSUBS 0.062448f
C520 VTAIL.n59 VSUBS 0.101633f
C521 VTAIL.n60 VSUBS 0.359485f
C522 VTAIL.n61 VSUBS 0.012163f
C523 VTAIL.n62 VSUBS 0.012878f
C524 VTAIL.n63 VSUBS 0.028748f
C525 VTAIL.n64 VSUBS 0.028748f
C526 VTAIL.n65 VSUBS 0.012878f
C527 VTAIL.n66 VSUBS 0.012163f
C528 VTAIL.n67 VSUBS 0.022634f
C529 VTAIL.n68 VSUBS 0.059429f
C530 VTAIL.n69 VSUBS 0.012163f
C531 VTAIL.n70 VSUBS 0.012878f
C532 VTAIL.n71 VSUBS 0.06241f
C533 VTAIL.n72 VSUBS 0.042995f
C534 VTAIL.n73 VSUBS 0.70371f
C535 VTAIL.n74 VSUBS 0.012776f
C536 VTAIL.n75 VSUBS 0.028748f
C537 VTAIL.n76 VSUBS 0.012878f
C538 VTAIL.n77 VSUBS 0.022634f
C539 VTAIL.n78 VSUBS 0.012163f
C540 VTAIL.n79 VSUBS 0.021561f
C541 VTAIL.n80 VSUBS 0.02155f
C542 VTAIL.t4 VSUBS 0.062448f
C543 VTAIL.n81 VSUBS 0.101633f
C544 VTAIL.n82 VSUBS 0.359485f
C545 VTAIL.n83 VSUBS 0.012163f
C546 VTAIL.n84 VSUBS 0.012878f
C547 VTAIL.n85 VSUBS 0.028748f
C548 VTAIL.n86 VSUBS 0.028748f
C549 VTAIL.n87 VSUBS 0.012878f
C550 VTAIL.n88 VSUBS 0.012163f
C551 VTAIL.n89 VSUBS 0.022634f
C552 VTAIL.n90 VSUBS 0.059429f
C553 VTAIL.n91 VSUBS 0.012163f
C554 VTAIL.n92 VSUBS 0.012878f
C555 VTAIL.n93 VSUBS 0.06241f
C556 VTAIL.n94 VSUBS 0.042995f
C557 VTAIL.n95 VSUBS 0.687363f
C558 VDD1.n0 VSUBS 0.011071f
C559 VDD1.n1 VSUBS 0.02491f
C560 VDD1.n2 VSUBS 0.011159f
C561 VDD1.n3 VSUBS 0.019612f
C562 VDD1.n4 VSUBS 0.010539f
C563 VDD1.n5 VSUBS 0.018683f
C564 VDD1.n6 VSUBS 0.018673f
C565 VDD1.t2 VSUBS 0.054111f
C566 VDD1.n7 VSUBS 0.088064f
C567 VDD1.n8 VSUBS 0.311492f
C568 VDD1.n9 VSUBS 0.010539f
C569 VDD1.n10 VSUBS 0.011159f
C570 VDD1.n11 VSUBS 0.02491f
C571 VDD1.n12 VSUBS 0.02491f
C572 VDD1.n13 VSUBS 0.011159f
C573 VDD1.n14 VSUBS 0.010539f
C574 VDD1.n15 VSUBS 0.019612f
C575 VDD1.n16 VSUBS 0.051495f
C576 VDD1.n17 VSUBS 0.010539f
C577 VDD1.n18 VSUBS 0.011159f
C578 VDD1.n19 VSUBS 0.054078f
C579 VDD1.n20 VSUBS 0.051586f
C580 VDD1.n21 VSUBS 0.011071f
C581 VDD1.n22 VSUBS 0.02491f
C582 VDD1.n23 VSUBS 0.011159f
C583 VDD1.n24 VSUBS 0.019612f
C584 VDD1.n25 VSUBS 0.010539f
C585 VDD1.n26 VSUBS 0.018683f
C586 VDD1.n27 VSUBS 0.018673f
C587 VDD1.t0 VSUBS 0.054111f
C588 VDD1.n28 VSUBS 0.088064f
C589 VDD1.n29 VSUBS 0.311492f
C590 VDD1.n30 VSUBS 0.010539f
C591 VDD1.n31 VSUBS 0.011159f
C592 VDD1.n32 VSUBS 0.02491f
C593 VDD1.n33 VSUBS 0.02491f
C594 VDD1.n34 VSUBS 0.011159f
C595 VDD1.n35 VSUBS 0.010539f
C596 VDD1.n36 VSUBS 0.019612f
C597 VDD1.n37 VSUBS 0.051495f
C598 VDD1.n38 VSUBS 0.010539f
C599 VDD1.n39 VSUBS 0.011159f
C600 VDD1.n40 VSUBS 0.054078f
C601 VDD1.n41 VSUBS 0.051369f
C602 VDD1.t4 VSUBS 0.068657f
C603 VDD1.t1 VSUBS 0.068657f
C604 VDD1.n42 VSUBS 0.427771f
C605 VDD1.n43 VSUBS 1.18484f
C606 VDD1.t3 VSUBS 0.068657f
C607 VDD1.t5 VSUBS 0.068657f
C608 VDD1.n44 VSUBS 0.427424f
C609 VDD1.n45 VSUBS 1.35013f
C610 VP.n0 VSUBS 0.050636f
C611 VP.t2 VSUBS 0.292969f
C612 VP.t5 VSUBS 0.300587f
C613 VP.n1 VSUBS 0.142843f
C614 VP.t0 VSUBS 0.289924f
C615 VP.n2 VSUBS 0.158742f
C616 VP.t3 VSUBS 0.292969f
C617 VP.n3 VSUBS 0.150078f
C618 VP.n4 VSUBS 1.58853f
C619 VP.n5 VSUBS 1.52531f
C620 VP.n6 VSUBS 0.150078f
C621 VP.t4 VSUBS 0.289924f
C622 VP.n7 VSUBS 0.158742f
C623 VP.t1 VSUBS 0.292969f
C624 VP.n8 VSUBS 0.150078f
C625 VP.n9 VSUBS 0.039241f
.ends

