* NGSPICE file created from diff_pair_sample_1294.ext - technology: sky130A

.subckt diff_pair_sample_1294 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=0 ps=0 w=15.12 l=1.16
X1 VDD1.t9 VP.t0 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X2 VDD2.t9 VN.t0 VTAIL.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X3 VDD2.t8 VN.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=5.8968 ps=31.02 w=15.12 l=1.16
X4 VTAIL.t15 VP.t1 VDD1.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X5 VDD1.t7 VP.t2 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=2.4948 ps=15.45 w=15.12 l=1.16
X6 VTAIL.t14 VP.t3 VDD1.t6 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X7 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=0 ps=0 w=15.12 l=1.16
X8 VTAIL.t3 VN.t2 VDD2.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X9 VDD1.t5 VP.t4 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=5.8968 ps=31.02 w=15.12 l=1.16
X10 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=0 ps=0 w=15.12 l=1.16
X11 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=0 ps=0 w=15.12 l=1.16
X12 VDD1.t4 VP.t5 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=2.4948 ps=15.45 w=15.12 l=1.16
X13 VDD2.t6 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X14 VDD2.t5 VN.t4 VTAIL.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=5.8968 ps=31.02 w=15.12 l=1.16
X15 VDD2.t4 VN.t5 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=2.4948 ps=15.45 w=15.12 l=1.16
X16 VTAIL.t9 VP.t6 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X17 VDD2.t3 VN.t6 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.8968 pd=31.02 as=2.4948 ps=15.45 w=15.12 l=1.16
X18 VDD1.t2 VP.t7 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X19 VTAIL.t4 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X20 VDD1.t1 VP.t8 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=5.8968 ps=31.02 w=15.12 l=1.16
X21 VTAIL.t18 VP.t9 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X22 VTAIL.t1 VN.t8 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
X23 VTAIL.t19 VN.t9 VDD2.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=2.4948 pd=15.45 as=2.4948 ps=15.45 w=15.12 l=1.16
R0 B.n623 B.n622 585
R1 B.n623 B.n64 585
R2 B.n626 B.n625 585
R3 B.n627 B.n124 585
R4 B.n629 B.n628 585
R5 B.n631 B.n123 585
R6 B.n634 B.n633 585
R7 B.n635 B.n122 585
R8 B.n637 B.n636 585
R9 B.n639 B.n121 585
R10 B.n642 B.n641 585
R11 B.n643 B.n120 585
R12 B.n645 B.n644 585
R13 B.n647 B.n119 585
R14 B.n650 B.n649 585
R15 B.n651 B.n118 585
R16 B.n653 B.n652 585
R17 B.n655 B.n117 585
R18 B.n658 B.n657 585
R19 B.n659 B.n116 585
R20 B.n661 B.n660 585
R21 B.n663 B.n115 585
R22 B.n666 B.n665 585
R23 B.n667 B.n114 585
R24 B.n669 B.n668 585
R25 B.n671 B.n113 585
R26 B.n674 B.n673 585
R27 B.n675 B.n112 585
R28 B.n677 B.n676 585
R29 B.n679 B.n111 585
R30 B.n682 B.n681 585
R31 B.n683 B.n110 585
R32 B.n685 B.n684 585
R33 B.n687 B.n109 585
R34 B.n690 B.n689 585
R35 B.n691 B.n108 585
R36 B.n693 B.n692 585
R37 B.n695 B.n107 585
R38 B.n698 B.n697 585
R39 B.n699 B.n106 585
R40 B.n701 B.n700 585
R41 B.n703 B.n105 585
R42 B.n706 B.n705 585
R43 B.n707 B.n104 585
R44 B.n709 B.n708 585
R45 B.n711 B.n103 585
R46 B.n714 B.n713 585
R47 B.n715 B.n102 585
R48 B.n717 B.n716 585
R49 B.n719 B.n101 585
R50 B.n722 B.n721 585
R51 B.n723 B.n98 585
R52 B.n726 B.n725 585
R53 B.n728 B.n97 585
R54 B.n731 B.n730 585
R55 B.n732 B.n96 585
R56 B.n734 B.n733 585
R57 B.n736 B.n95 585
R58 B.n739 B.n738 585
R59 B.n740 B.n91 585
R60 B.n742 B.n741 585
R61 B.n744 B.n90 585
R62 B.n747 B.n746 585
R63 B.n748 B.n89 585
R64 B.n750 B.n749 585
R65 B.n752 B.n88 585
R66 B.n755 B.n754 585
R67 B.n756 B.n87 585
R68 B.n758 B.n757 585
R69 B.n760 B.n86 585
R70 B.n763 B.n762 585
R71 B.n764 B.n85 585
R72 B.n766 B.n765 585
R73 B.n768 B.n84 585
R74 B.n771 B.n770 585
R75 B.n772 B.n83 585
R76 B.n774 B.n773 585
R77 B.n776 B.n82 585
R78 B.n779 B.n778 585
R79 B.n780 B.n81 585
R80 B.n782 B.n781 585
R81 B.n784 B.n80 585
R82 B.n787 B.n786 585
R83 B.n788 B.n79 585
R84 B.n790 B.n789 585
R85 B.n792 B.n78 585
R86 B.n795 B.n794 585
R87 B.n796 B.n77 585
R88 B.n798 B.n797 585
R89 B.n800 B.n76 585
R90 B.n803 B.n802 585
R91 B.n804 B.n75 585
R92 B.n806 B.n805 585
R93 B.n808 B.n74 585
R94 B.n811 B.n810 585
R95 B.n812 B.n73 585
R96 B.n814 B.n813 585
R97 B.n816 B.n72 585
R98 B.n819 B.n818 585
R99 B.n820 B.n71 585
R100 B.n822 B.n821 585
R101 B.n824 B.n70 585
R102 B.n827 B.n826 585
R103 B.n828 B.n69 585
R104 B.n830 B.n829 585
R105 B.n832 B.n68 585
R106 B.n835 B.n834 585
R107 B.n836 B.n67 585
R108 B.n838 B.n837 585
R109 B.n840 B.n66 585
R110 B.n843 B.n842 585
R111 B.n844 B.n65 585
R112 B.n621 B.n63 585
R113 B.n847 B.n63 585
R114 B.n620 B.n62 585
R115 B.n848 B.n62 585
R116 B.n619 B.n61 585
R117 B.n849 B.n61 585
R118 B.n618 B.n617 585
R119 B.n617 B.n57 585
R120 B.n616 B.n56 585
R121 B.n855 B.n56 585
R122 B.n615 B.n55 585
R123 B.n856 B.n55 585
R124 B.n614 B.n54 585
R125 B.n857 B.n54 585
R126 B.n613 B.n612 585
R127 B.n612 B.n50 585
R128 B.n611 B.n49 585
R129 B.n863 B.n49 585
R130 B.n610 B.n48 585
R131 B.n864 B.n48 585
R132 B.n609 B.n47 585
R133 B.n865 B.n47 585
R134 B.n608 B.n607 585
R135 B.n607 B.n43 585
R136 B.n606 B.n42 585
R137 B.n871 B.n42 585
R138 B.n605 B.n41 585
R139 B.n872 B.n41 585
R140 B.n604 B.n40 585
R141 B.n873 B.n40 585
R142 B.n603 B.n602 585
R143 B.n602 B.n36 585
R144 B.n601 B.n35 585
R145 B.n879 B.n35 585
R146 B.n600 B.n34 585
R147 B.n880 B.n34 585
R148 B.n599 B.n33 585
R149 B.n881 B.n33 585
R150 B.n598 B.n597 585
R151 B.n597 B.n29 585
R152 B.n596 B.n28 585
R153 B.n887 B.n28 585
R154 B.n595 B.n27 585
R155 B.n888 B.n27 585
R156 B.n594 B.n26 585
R157 B.n889 B.n26 585
R158 B.n593 B.n592 585
R159 B.n592 B.n22 585
R160 B.n591 B.n21 585
R161 B.n895 B.n21 585
R162 B.n590 B.n20 585
R163 B.n896 B.n20 585
R164 B.n589 B.n19 585
R165 B.n897 B.n19 585
R166 B.n588 B.n587 585
R167 B.n587 B.n15 585
R168 B.n586 B.n14 585
R169 B.n903 B.n14 585
R170 B.n585 B.n13 585
R171 B.n904 B.n13 585
R172 B.n584 B.n12 585
R173 B.n905 B.n12 585
R174 B.n583 B.n582 585
R175 B.n582 B.n581 585
R176 B.n580 B.n579 585
R177 B.n580 B.n8 585
R178 B.n578 B.n7 585
R179 B.n912 B.n7 585
R180 B.n577 B.n6 585
R181 B.n913 B.n6 585
R182 B.n576 B.n5 585
R183 B.n914 B.n5 585
R184 B.n575 B.n574 585
R185 B.n574 B.n4 585
R186 B.n573 B.n125 585
R187 B.n573 B.n572 585
R188 B.n563 B.n126 585
R189 B.n127 B.n126 585
R190 B.n565 B.n564 585
R191 B.n566 B.n565 585
R192 B.n562 B.n132 585
R193 B.n132 B.n131 585
R194 B.n561 B.n560 585
R195 B.n560 B.n559 585
R196 B.n134 B.n133 585
R197 B.n135 B.n134 585
R198 B.n552 B.n551 585
R199 B.n553 B.n552 585
R200 B.n550 B.n140 585
R201 B.n140 B.n139 585
R202 B.n549 B.n548 585
R203 B.n548 B.n547 585
R204 B.n142 B.n141 585
R205 B.n143 B.n142 585
R206 B.n540 B.n539 585
R207 B.n541 B.n540 585
R208 B.n538 B.n147 585
R209 B.n151 B.n147 585
R210 B.n537 B.n536 585
R211 B.n536 B.n535 585
R212 B.n149 B.n148 585
R213 B.n150 B.n149 585
R214 B.n528 B.n527 585
R215 B.n529 B.n528 585
R216 B.n526 B.n155 585
R217 B.n159 B.n155 585
R218 B.n525 B.n524 585
R219 B.n524 B.n523 585
R220 B.n157 B.n156 585
R221 B.n158 B.n157 585
R222 B.n516 B.n515 585
R223 B.n517 B.n516 585
R224 B.n514 B.n163 585
R225 B.n167 B.n163 585
R226 B.n513 B.n512 585
R227 B.n512 B.n511 585
R228 B.n165 B.n164 585
R229 B.n166 B.n165 585
R230 B.n504 B.n503 585
R231 B.n505 B.n504 585
R232 B.n502 B.n172 585
R233 B.n172 B.n171 585
R234 B.n501 B.n500 585
R235 B.n500 B.n499 585
R236 B.n174 B.n173 585
R237 B.n175 B.n174 585
R238 B.n492 B.n491 585
R239 B.n493 B.n492 585
R240 B.n490 B.n179 585
R241 B.n183 B.n179 585
R242 B.n489 B.n488 585
R243 B.n488 B.n487 585
R244 B.n181 B.n180 585
R245 B.n182 B.n181 585
R246 B.n480 B.n479 585
R247 B.n481 B.n480 585
R248 B.n478 B.n188 585
R249 B.n188 B.n187 585
R250 B.n477 B.n476 585
R251 B.n476 B.n475 585
R252 B.n472 B.n192 585
R253 B.n471 B.n470 585
R254 B.n468 B.n193 585
R255 B.n468 B.n191 585
R256 B.n467 B.n466 585
R257 B.n465 B.n464 585
R258 B.n463 B.n195 585
R259 B.n461 B.n460 585
R260 B.n459 B.n196 585
R261 B.n458 B.n457 585
R262 B.n455 B.n197 585
R263 B.n453 B.n452 585
R264 B.n451 B.n198 585
R265 B.n450 B.n449 585
R266 B.n447 B.n199 585
R267 B.n445 B.n444 585
R268 B.n443 B.n200 585
R269 B.n442 B.n441 585
R270 B.n439 B.n201 585
R271 B.n437 B.n436 585
R272 B.n435 B.n202 585
R273 B.n434 B.n433 585
R274 B.n431 B.n203 585
R275 B.n429 B.n428 585
R276 B.n427 B.n204 585
R277 B.n426 B.n425 585
R278 B.n423 B.n205 585
R279 B.n421 B.n420 585
R280 B.n419 B.n206 585
R281 B.n418 B.n417 585
R282 B.n415 B.n207 585
R283 B.n413 B.n412 585
R284 B.n411 B.n208 585
R285 B.n410 B.n409 585
R286 B.n407 B.n209 585
R287 B.n405 B.n404 585
R288 B.n403 B.n210 585
R289 B.n402 B.n401 585
R290 B.n399 B.n211 585
R291 B.n397 B.n396 585
R292 B.n395 B.n212 585
R293 B.n394 B.n393 585
R294 B.n391 B.n213 585
R295 B.n389 B.n388 585
R296 B.n387 B.n214 585
R297 B.n386 B.n385 585
R298 B.n383 B.n215 585
R299 B.n381 B.n380 585
R300 B.n379 B.n216 585
R301 B.n378 B.n377 585
R302 B.n375 B.n217 585
R303 B.n373 B.n372 585
R304 B.n370 B.n218 585
R305 B.n369 B.n368 585
R306 B.n366 B.n221 585
R307 B.n364 B.n363 585
R308 B.n362 B.n222 585
R309 B.n361 B.n360 585
R310 B.n358 B.n223 585
R311 B.n356 B.n355 585
R312 B.n354 B.n224 585
R313 B.n352 B.n351 585
R314 B.n349 B.n227 585
R315 B.n347 B.n346 585
R316 B.n345 B.n228 585
R317 B.n344 B.n343 585
R318 B.n341 B.n229 585
R319 B.n339 B.n338 585
R320 B.n337 B.n230 585
R321 B.n336 B.n335 585
R322 B.n333 B.n231 585
R323 B.n331 B.n330 585
R324 B.n329 B.n232 585
R325 B.n328 B.n327 585
R326 B.n325 B.n233 585
R327 B.n323 B.n322 585
R328 B.n321 B.n234 585
R329 B.n320 B.n319 585
R330 B.n317 B.n235 585
R331 B.n315 B.n314 585
R332 B.n313 B.n236 585
R333 B.n312 B.n311 585
R334 B.n309 B.n237 585
R335 B.n307 B.n306 585
R336 B.n305 B.n238 585
R337 B.n304 B.n303 585
R338 B.n301 B.n239 585
R339 B.n299 B.n298 585
R340 B.n297 B.n240 585
R341 B.n296 B.n295 585
R342 B.n293 B.n241 585
R343 B.n291 B.n290 585
R344 B.n289 B.n242 585
R345 B.n288 B.n287 585
R346 B.n285 B.n243 585
R347 B.n283 B.n282 585
R348 B.n281 B.n244 585
R349 B.n280 B.n279 585
R350 B.n277 B.n245 585
R351 B.n275 B.n274 585
R352 B.n273 B.n246 585
R353 B.n272 B.n271 585
R354 B.n269 B.n247 585
R355 B.n267 B.n266 585
R356 B.n265 B.n248 585
R357 B.n264 B.n263 585
R358 B.n261 B.n249 585
R359 B.n259 B.n258 585
R360 B.n257 B.n250 585
R361 B.n256 B.n255 585
R362 B.n253 B.n251 585
R363 B.n190 B.n189 585
R364 B.n474 B.n473 585
R365 B.n475 B.n474 585
R366 B.n186 B.n185 585
R367 B.n187 B.n186 585
R368 B.n483 B.n482 585
R369 B.n482 B.n481 585
R370 B.n484 B.n184 585
R371 B.n184 B.n182 585
R372 B.n486 B.n485 585
R373 B.n487 B.n486 585
R374 B.n178 B.n177 585
R375 B.n183 B.n178 585
R376 B.n495 B.n494 585
R377 B.n494 B.n493 585
R378 B.n496 B.n176 585
R379 B.n176 B.n175 585
R380 B.n498 B.n497 585
R381 B.n499 B.n498 585
R382 B.n170 B.n169 585
R383 B.n171 B.n170 585
R384 B.n507 B.n506 585
R385 B.n506 B.n505 585
R386 B.n508 B.n168 585
R387 B.n168 B.n166 585
R388 B.n510 B.n509 585
R389 B.n511 B.n510 585
R390 B.n162 B.n161 585
R391 B.n167 B.n162 585
R392 B.n519 B.n518 585
R393 B.n518 B.n517 585
R394 B.n520 B.n160 585
R395 B.n160 B.n158 585
R396 B.n522 B.n521 585
R397 B.n523 B.n522 585
R398 B.n154 B.n153 585
R399 B.n159 B.n154 585
R400 B.n531 B.n530 585
R401 B.n530 B.n529 585
R402 B.n532 B.n152 585
R403 B.n152 B.n150 585
R404 B.n534 B.n533 585
R405 B.n535 B.n534 585
R406 B.n146 B.n145 585
R407 B.n151 B.n146 585
R408 B.n543 B.n542 585
R409 B.n542 B.n541 585
R410 B.n544 B.n144 585
R411 B.n144 B.n143 585
R412 B.n546 B.n545 585
R413 B.n547 B.n546 585
R414 B.n138 B.n137 585
R415 B.n139 B.n138 585
R416 B.n555 B.n554 585
R417 B.n554 B.n553 585
R418 B.n556 B.n136 585
R419 B.n136 B.n135 585
R420 B.n558 B.n557 585
R421 B.n559 B.n558 585
R422 B.n130 B.n129 585
R423 B.n131 B.n130 585
R424 B.n568 B.n567 585
R425 B.n567 B.n566 585
R426 B.n569 B.n128 585
R427 B.n128 B.n127 585
R428 B.n571 B.n570 585
R429 B.n572 B.n571 585
R430 B.n3 B.n0 585
R431 B.n4 B.n3 585
R432 B.n911 B.n1 585
R433 B.n912 B.n911 585
R434 B.n910 B.n909 585
R435 B.n910 B.n8 585
R436 B.n908 B.n9 585
R437 B.n581 B.n9 585
R438 B.n907 B.n906 585
R439 B.n906 B.n905 585
R440 B.n11 B.n10 585
R441 B.n904 B.n11 585
R442 B.n902 B.n901 585
R443 B.n903 B.n902 585
R444 B.n900 B.n16 585
R445 B.n16 B.n15 585
R446 B.n899 B.n898 585
R447 B.n898 B.n897 585
R448 B.n18 B.n17 585
R449 B.n896 B.n18 585
R450 B.n894 B.n893 585
R451 B.n895 B.n894 585
R452 B.n892 B.n23 585
R453 B.n23 B.n22 585
R454 B.n891 B.n890 585
R455 B.n890 B.n889 585
R456 B.n25 B.n24 585
R457 B.n888 B.n25 585
R458 B.n886 B.n885 585
R459 B.n887 B.n886 585
R460 B.n884 B.n30 585
R461 B.n30 B.n29 585
R462 B.n883 B.n882 585
R463 B.n882 B.n881 585
R464 B.n32 B.n31 585
R465 B.n880 B.n32 585
R466 B.n878 B.n877 585
R467 B.n879 B.n878 585
R468 B.n876 B.n37 585
R469 B.n37 B.n36 585
R470 B.n875 B.n874 585
R471 B.n874 B.n873 585
R472 B.n39 B.n38 585
R473 B.n872 B.n39 585
R474 B.n870 B.n869 585
R475 B.n871 B.n870 585
R476 B.n868 B.n44 585
R477 B.n44 B.n43 585
R478 B.n867 B.n866 585
R479 B.n866 B.n865 585
R480 B.n46 B.n45 585
R481 B.n864 B.n46 585
R482 B.n862 B.n861 585
R483 B.n863 B.n862 585
R484 B.n860 B.n51 585
R485 B.n51 B.n50 585
R486 B.n859 B.n858 585
R487 B.n858 B.n857 585
R488 B.n53 B.n52 585
R489 B.n856 B.n53 585
R490 B.n854 B.n853 585
R491 B.n855 B.n854 585
R492 B.n852 B.n58 585
R493 B.n58 B.n57 585
R494 B.n851 B.n850 585
R495 B.n850 B.n849 585
R496 B.n60 B.n59 585
R497 B.n848 B.n60 585
R498 B.n846 B.n845 585
R499 B.n847 B.n846 585
R500 B.n915 B.n914 585
R501 B.n913 B.n2 585
R502 B.n92 B.t14 518.034
R503 B.n99 B.t18 518.034
R504 B.n225 B.t10 518.034
R505 B.n219 B.t21 518.034
R506 B.n846 B.n65 497.305
R507 B.n623 B.n63 497.305
R508 B.n476 B.n190 497.305
R509 B.n474 B.n192 497.305
R510 B.n624 B.n64 256.663
R511 B.n630 B.n64 256.663
R512 B.n632 B.n64 256.663
R513 B.n638 B.n64 256.663
R514 B.n640 B.n64 256.663
R515 B.n646 B.n64 256.663
R516 B.n648 B.n64 256.663
R517 B.n654 B.n64 256.663
R518 B.n656 B.n64 256.663
R519 B.n662 B.n64 256.663
R520 B.n664 B.n64 256.663
R521 B.n670 B.n64 256.663
R522 B.n672 B.n64 256.663
R523 B.n678 B.n64 256.663
R524 B.n680 B.n64 256.663
R525 B.n686 B.n64 256.663
R526 B.n688 B.n64 256.663
R527 B.n694 B.n64 256.663
R528 B.n696 B.n64 256.663
R529 B.n702 B.n64 256.663
R530 B.n704 B.n64 256.663
R531 B.n710 B.n64 256.663
R532 B.n712 B.n64 256.663
R533 B.n718 B.n64 256.663
R534 B.n720 B.n64 256.663
R535 B.n727 B.n64 256.663
R536 B.n729 B.n64 256.663
R537 B.n735 B.n64 256.663
R538 B.n737 B.n64 256.663
R539 B.n743 B.n64 256.663
R540 B.n745 B.n64 256.663
R541 B.n751 B.n64 256.663
R542 B.n753 B.n64 256.663
R543 B.n759 B.n64 256.663
R544 B.n761 B.n64 256.663
R545 B.n767 B.n64 256.663
R546 B.n769 B.n64 256.663
R547 B.n775 B.n64 256.663
R548 B.n777 B.n64 256.663
R549 B.n783 B.n64 256.663
R550 B.n785 B.n64 256.663
R551 B.n791 B.n64 256.663
R552 B.n793 B.n64 256.663
R553 B.n799 B.n64 256.663
R554 B.n801 B.n64 256.663
R555 B.n807 B.n64 256.663
R556 B.n809 B.n64 256.663
R557 B.n815 B.n64 256.663
R558 B.n817 B.n64 256.663
R559 B.n823 B.n64 256.663
R560 B.n825 B.n64 256.663
R561 B.n831 B.n64 256.663
R562 B.n833 B.n64 256.663
R563 B.n839 B.n64 256.663
R564 B.n841 B.n64 256.663
R565 B.n469 B.n191 256.663
R566 B.n194 B.n191 256.663
R567 B.n462 B.n191 256.663
R568 B.n456 B.n191 256.663
R569 B.n454 B.n191 256.663
R570 B.n448 B.n191 256.663
R571 B.n446 B.n191 256.663
R572 B.n440 B.n191 256.663
R573 B.n438 B.n191 256.663
R574 B.n432 B.n191 256.663
R575 B.n430 B.n191 256.663
R576 B.n424 B.n191 256.663
R577 B.n422 B.n191 256.663
R578 B.n416 B.n191 256.663
R579 B.n414 B.n191 256.663
R580 B.n408 B.n191 256.663
R581 B.n406 B.n191 256.663
R582 B.n400 B.n191 256.663
R583 B.n398 B.n191 256.663
R584 B.n392 B.n191 256.663
R585 B.n390 B.n191 256.663
R586 B.n384 B.n191 256.663
R587 B.n382 B.n191 256.663
R588 B.n376 B.n191 256.663
R589 B.n374 B.n191 256.663
R590 B.n367 B.n191 256.663
R591 B.n365 B.n191 256.663
R592 B.n359 B.n191 256.663
R593 B.n357 B.n191 256.663
R594 B.n350 B.n191 256.663
R595 B.n348 B.n191 256.663
R596 B.n342 B.n191 256.663
R597 B.n340 B.n191 256.663
R598 B.n334 B.n191 256.663
R599 B.n332 B.n191 256.663
R600 B.n326 B.n191 256.663
R601 B.n324 B.n191 256.663
R602 B.n318 B.n191 256.663
R603 B.n316 B.n191 256.663
R604 B.n310 B.n191 256.663
R605 B.n308 B.n191 256.663
R606 B.n302 B.n191 256.663
R607 B.n300 B.n191 256.663
R608 B.n294 B.n191 256.663
R609 B.n292 B.n191 256.663
R610 B.n286 B.n191 256.663
R611 B.n284 B.n191 256.663
R612 B.n278 B.n191 256.663
R613 B.n276 B.n191 256.663
R614 B.n270 B.n191 256.663
R615 B.n268 B.n191 256.663
R616 B.n262 B.n191 256.663
R617 B.n260 B.n191 256.663
R618 B.n254 B.n191 256.663
R619 B.n252 B.n191 256.663
R620 B.n917 B.n916 256.663
R621 B.n842 B.n840 163.367
R622 B.n838 B.n67 163.367
R623 B.n834 B.n832 163.367
R624 B.n830 B.n69 163.367
R625 B.n826 B.n824 163.367
R626 B.n822 B.n71 163.367
R627 B.n818 B.n816 163.367
R628 B.n814 B.n73 163.367
R629 B.n810 B.n808 163.367
R630 B.n806 B.n75 163.367
R631 B.n802 B.n800 163.367
R632 B.n798 B.n77 163.367
R633 B.n794 B.n792 163.367
R634 B.n790 B.n79 163.367
R635 B.n786 B.n784 163.367
R636 B.n782 B.n81 163.367
R637 B.n778 B.n776 163.367
R638 B.n774 B.n83 163.367
R639 B.n770 B.n768 163.367
R640 B.n766 B.n85 163.367
R641 B.n762 B.n760 163.367
R642 B.n758 B.n87 163.367
R643 B.n754 B.n752 163.367
R644 B.n750 B.n89 163.367
R645 B.n746 B.n744 163.367
R646 B.n742 B.n91 163.367
R647 B.n738 B.n736 163.367
R648 B.n734 B.n96 163.367
R649 B.n730 B.n728 163.367
R650 B.n726 B.n98 163.367
R651 B.n721 B.n719 163.367
R652 B.n717 B.n102 163.367
R653 B.n713 B.n711 163.367
R654 B.n709 B.n104 163.367
R655 B.n705 B.n703 163.367
R656 B.n701 B.n106 163.367
R657 B.n697 B.n695 163.367
R658 B.n693 B.n108 163.367
R659 B.n689 B.n687 163.367
R660 B.n685 B.n110 163.367
R661 B.n681 B.n679 163.367
R662 B.n677 B.n112 163.367
R663 B.n673 B.n671 163.367
R664 B.n669 B.n114 163.367
R665 B.n665 B.n663 163.367
R666 B.n661 B.n116 163.367
R667 B.n657 B.n655 163.367
R668 B.n653 B.n118 163.367
R669 B.n649 B.n647 163.367
R670 B.n645 B.n120 163.367
R671 B.n641 B.n639 163.367
R672 B.n637 B.n122 163.367
R673 B.n633 B.n631 163.367
R674 B.n629 B.n124 163.367
R675 B.n625 B.n623 163.367
R676 B.n476 B.n188 163.367
R677 B.n480 B.n188 163.367
R678 B.n480 B.n181 163.367
R679 B.n488 B.n181 163.367
R680 B.n488 B.n179 163.367
R681 B.n492 B.n179 163.367
R682 B.n492 B.n174 163.367
R683 B.n500 B.n174 163.367
R684 B.n500 B.n172 163.367
R685 B.n504 B.n172 163.367
R686 B.n504 B.n165 163.367
R687 B.n512 B.n165 163.367
R688 B.n512 B.n163 163.367
R689 B.n516 B.n163 163.367
R690 B.n516 B.n157 163.367
R691 B.n524 B.n157 163.367
R692 B.n524 B.n155 163.367
R693 B.n528 B.n155 163.367
R694 B.n528 B.n149 163.367
R695 B.n536 B.n149 163.367
R696 B.n536 B.n147 163.367
R697 B.n540 B.n147 163.367
R698 B.n540 B.n142 163.367
R699 B.n548 B.n142 163.367
R700 B.n548 B.n140 163.367
R701 B.n552 B.n140 163.367
R702 B.n552 B.n134 163.367
R703 B.n560 B.n134 163.367
R704 B.n560 B.n132 163.367
R705 B.n565 B.n132 163.367
R706 B.n565 B.n126 163.367
R707 B.n573 B.n126 163.367
R708 B.n574 B.n573 163.367
R709 B.n574 B.n5 163.367
R710 B.n6 B.n5 163.367
R711 B.n7 B.n6 163.367
R712 B.n580 B.n7 163.367
R713 B.n582 B.n580 163.367
R714 B.n582 B.n12 163.367
R715 B.n13 B.n12 163.367
R716 B.n14 B.n13 163.367
R717 B.n587 B.n14 163.367
R718 B.n587 B.n19 163.367
R719 B.n20 B.n19 163.367
R720 B.n21 B.n20 163.367
R721 B.n592 B.n21 163.367
R722 B.n592 B.n26 163.367
R723 B.n27 B.n26 163.367
R724 B.n28 B.n27 163.367
R725 B.n597 B.n28 163.367
R726 B.n597 B.n33 163.367
R727 B.n34 B.n33 163.367
R728 B.n35 B.n34 163.367
R729 B.n602 B.n35 163.367
R730 B.n602 B.n40 163.367
R731 B.n41 B.n40 163.367
R732 B.n42 B.n41 163.367
R733 B.n607 B.n42 163.367
R734 B.n607 B.n47 163.367
R735 B.n48 B.n47 163.367
R736 B.n49 B.n48 163.367
R737 B.n612 B.n49 163.367
R738 B.n612 B.n54 163.367
R739 B.n55 B.n54 163.367
R740 B.n56 B.n55 163.367
R741 B.n617 B.n56 163.367
R742 B.n617 B.n61 163.367
R743 B.n62 B.n61 163.367
R744 B.n63 B.n62 163.367
R745 B.n470 B.n468 163.367
R746 B.n468 B.n467 163.367
R747 B.n464 B.n463 163.367
R748 B.n461 B.n196 163.367
R749 B.n457 B.n455 163.367
R750 B.n453 B.n198 163.367
R751 B.n449 B.n447 163.367
R752 B.n445 B.n200 163.367
R753 B.n441 B.n439 163.367
R754 B.n437 B.n202 163.367
R755 B.n433 B.n431 163.367
R756 B.n429 B.n204 163.367
R757 B.n425 B.n423 163.367
R758 B.n421 B.n206 163.367
R759 B.n417 B.n415 163.367
R760 B.n413 B.n208 163.367
R761 B.n409 B.n407 163.367
R762 B.n405 B.n210 163.367
R763 B.n401 B.n399 163.367
R764 B.n397 B.n212 163.367
R765 B.n393 B.n391 163.367
R766 B.n389 B.n214 163.367
R767 B.n385 B.n383 163.367
R768 B.n381 B.n216 163.367
R769 B.n377 B.n375 163.367
R770 B.n373 B.n218 163.367
R771 B.n368 B.n366 163.367
R772 B.n364 B.n222 163.367
R773 B.n360 B.n358 163.367
R774 B.n356 B.n224 163.367
R775 B.n351 B.n349 163.367
R776 B.n347 B.n228 163.367
R777 B.n343 B.n341 163.367
R778 B.n339 B.n230 163.367
R779 B.n335 B.n333 163.367
R780 B.n331 B.n232 163.367
R781 B.n327 B.n325 163.367
R782 B.n323 B.n234 163.367
R783 B.n319 B.n317 163.367
R784 B.n315 B.n236 163.367
R785 B.n311 B.n309 163.367
R786 B.n307 B.n238 163.367
R787 B.n303 B.n301 163.367
R788 B.n299 B.n240 163.367
R789 B.n295 B.n293 163.367
R790 B.n291 B.n242 163.367
R791 B.n287 B.n285 163.367
R792 B.n283 B.n244 163.367
R793 B.n279 B.n277 163.367
R794 B.n275 B.n246 163.367
R795 B.n271 B.n269 163.367
R796 B.n267 B.n248 163.367
R797 B.n263 B.n261 163.367
R798 B.n259 B.n250 163.367
R799 B.n255 B.n253 163.367
R800 B.n474 B.n186 163.367
R801 B.n482 B.n186 163.367
R802 B.n482 B.n184 163.367
R803 B.n486 B.n184 163.367
R804 B.n486 B.n178 163.367
R805 B.n494 B.n178 163.367
R806 B.n494 B.n176 163.367
R807 B.n498 B.n176 163.367
R808 B.n498 B.n170 163.367
R809 B.n506 B.n170 163.367
R810 B.n506 B.n168 163.367
R811 B.n510 B.n168 163.367
R812 B.n510 B.n162 163.367
R813 B.n518 B.n162 163.367
R814 B.n518 B.n160 163.367
R815 B.n522 B.n160 163.367
R816 B.n522 B.n154 163.367
R817 B.n530 B.n154 163.367
R818 B.n530 B.n152 163.367
R819 B.n534 B.n152 163.367
R820 B.n534 B.n146 163.367
R821 B.n542 B.n146 163.367
R822 B.n542 B.n144 163.367
R823 B.n546 B.n144 163.367
R824 B.n546 B.n138 163.367
R825 B.n554 B.n138 163.367
R826 B.n554 B.n136 163.367
R827 B.n558 B.n136 163.367
R828 B.n558 B.n130 163.367
R829 B.n567 B.n130 163.367
R830 B.n567 B.n128 163.367
R831 B.n571 B.n128 163.367
R832 B.n571 B.n3 163.367
R833 B.n915 B.n3 163.367
R834 B.n911 B.n2 163.367
R835 B.n911 B.n910 163.367
R836 B.n910 B.n9 163.367
R837 B.n906 B.n9 163.367
R838 B.n906 B.n11 163.367
R839 B.n902 B.n11 163.367
R840 B.n902 B.n16 163.367
R841 B.n898 B.n16 163.367
R842 B.n898 B.n18 163.367
R843 B.n894 B.n18 163.367
R844 B.n894 B.n23 163.367
R845 B.n890 B.n23 163.367
R846 B.n890 B.n25 163.367
R847 B.n886 B.n25 163.367
R848 B.n886 B.n30 163.367
R849 B.n882 B.n30 163.367
R850 B.n882 B.n32 163.367
R851 B.n878 B.n32 163.367
R852 B.n878 B.n37 163.367
R853 B.n874 B.n37 163.367
R854 B.n874 B.n39 163.367
R855 B.n870 B.n39 163.367
R856 B.n870 B.n44 163.367
R857 B.n866 B.n44 163.367
R858 B.n866 B.n46 163.367
R859 B.n862 B.n46 163.367
R860 B.n862 B.n51 163.367
R861 B.n858 B.n51 163.367
R862 B.n858 B.n53 163.367
R863 B.n854 B.n53 163.367
R864 B.n854 B.n58 163.367
R865 B.n850 B.n58 163.367
R866 B.n850 B.n60 163.367
R867 B.n846 B.n60 163.367
R868 B.n99 B.t19 99.4539
R869 B.n225 B.t13 99.4539
R870 B.n92 B.t16 99.4342
R871 B.n219 B.t23 99.4342
R872 B.n841 B.n65 71.676
R873 B.n840 B.n839 71.676
R874 B.n833 B.n67 71.676
R875 B.n832 B.n831 71.676
R876 B.n825 B.n69 71.676
R877 B.n824 B.n823 71.676
R878 B.n817 B.n71 71.676
R879 B.n816 B.n815 71.676
R880 B.n809 B.n73 71.676
R881 B.n808 B.n807 71.676
R882 B.n801 B.n75 71.676
R883 B.n800 B.n799 71.676
R884 B.n793 B.n77 71.676
R885 B.n792 B.n791 71.676
R886 B.n785 B.n79 71.676
R887 B.n784 B.n783 71.676
R888 B.n777 B.n81 71.676
R889 B.n776 B.n775 71.676
R890 B.n769 B.n83 71.676
R891 B.n768 B.n767 71.676
R892 B.n761 B.n85 71.676
R893 B.n760 B.n759 71.676
R894 B.n753 B.n87 71.676
R895 B.n752 B.n751 71.676
R896 B.n745 B.n89 71.676
R897 B.n744 B.n743 71.676
R898 B.n737 B.n91 71.676
R899 B.n736 B.n735 71.676
R900 B.n729 B.n96 71.676
R901 B.n728 B.n727 71.676
R902 B.n720 B.n98 71.676
R903 B.n719 B.n718 71.676
R904 B.n712 B.n102 71.676
R905 B.n711 B.n710 71.676
R906 B.n704 B.n104 71.676
R907 B.n703 B.n702 71.676
R908 B.n696 B.n106 71.676
R909 B.n695 B.n694 71.676
R910 B.n688 B.n108 71.676
R911 B.n687 B.n686 71.676
R912 B.n680 B.n110 71.676
R913 B.n679 B.n678 71.676
R914 B.n672 B.n112 71.676
R915 B.n671 B.n670 71.676
R916 B.n664 B.n114 71.676
R917 B.n663 B.n662 71.676
R918 B.n656 B.n116 71.676
R919 B.n655 B.n654 71.676
R920 B.n648 B.n118 71.676
R921 B.n647 B.n646 71.676
R922 B.n640 B.n120 71.676
R923 B.n639 B.n638 71.676
R924 B.n632 B.n122 71.676
R925 B.n631 B.n630 71.676
R926 B.n624 B.n124 71.676
R927 B.n625 B.n624 71.676
R928 B.n630 B.n629 71.676
R929 B.n633 B.n632 71.676
R930 B.n638 B.n637 71.676
R931 B.n641 B.n640 71.676
R932 B.n646 B.n645 71.676
R933 B.n649 B.n648 71.676
R934 B.n654 B.n653 71.676
R935 B.n657 B.n656 71.676
R936 B.n662 B.n661 71.676
R937 B.n665 B.n664 71.676
R938 B.n670 B.n669 71.676
R939 B.n673 B.n672 71.676
R940 B.n678 B.n677 71.676
R941 B.n681 B.n680 71.676
R942 B.n686 B.n685 71.676
R943 B.n689 B.n688 71.676
R944 B.n694 B.n693 71.676
R945 B.n697 B.n696 71.676
R946 B.n702 B.n701 71.676
R947 B.n705 B.n704 71.676
R948 B.n710 B.n709 71.676
R949 B.n713 B.n712 71.676
R950 B.n718 B.n717 71.676
R951 B.n721 B.n720 71.676
R952 B.n727 B.n726 71.676
R953 B.n730 B.n729 71.676
R954 B.n735 B.n734 71.676
R955 B.n738 B.n737 71.676
R956 B.n743 B.n742 71.676
R957 B.n746 B.n745 71.676
R958 B.n751 B.n750 71.676
R959 B.n754 B.n753 71.676
R960 B.n759 B.n758 71.676
R961 B.n762 B.n761 71.676
R962 B.n767 B.n766 71.676
R963 B.n770 B.n769 71.676
R964 B.n775 B.n774 71.676
R965 B.n778 B.n777 71.676
R966 B.n783 B.n782 71.676
R967 B.n786 B.n785 71.676
R968 B.n791 B.n790 71.676
R969 B.n794 B.n793 71.676
R970 B.n799 B.n798 71.676
R971 B.n802 B.n801 71.676
R972 B.n807 B.n806 71.676
R973 B.n810 B.n809 71.676
R974 B.n815 B.n814 71.676
R975 B.n818 B.n817 71.676
R976 B.n823 B.n822 71.676
R977 B.n826 B.n825 71.676
R978 B.n831 B.n830 71.676
R979 B.n834 B.n833 71.676
R980 B.n839 B.n838 71.676
R981 B.n842 B.n841 71.676
R982 B.n469 B.n192 71.676
R983 B.n467 B.n194 71.676
R984 B.n463 B.n462 71.676
R985 B.n456 B.n196 71.676
R986 B.n455 B.n454 71.676
R987 B.n448 B.n198 71.676
R988 B.n447 B.n446 71.676
R989 B.n440 B.n200 71.676
R990 B.n439 B.n438 71.676
R991 B.n432 B.n202 71.676
R992 B.n431 B.n430 71.676
R993 B.n424 B.n204 71.676
R994 B.n423 B.n422 71.676
R995 B.n416 B.n206 71.676
R996 B.n415 B.n414 71.676
R997 B.n408 B.n208 71.676
R998 B.n407 B.n406 71.676
R999 B.n400 B.n210 71.676
R1000 B.n399 B.n398 71.676
R1001 B.n392 B.n212 71.676
R1002 B.n391 B.n390 71.676
R1003 B.n384 B.n214 71.676
R1004 B.n383 B.n382 71.676
R1005 B.n376 B.n216 71.676
R1006 B.n375 B.n374 71.676
R1007 B.n367 B.n218 71.676
R1008 B.n366 B.n365 71.676
R1009 B.n359 B.n222 71.676
R1010 B.n358 B.n357 71.676
R1011 B.n350 B.n224 71.676
R1012 B.n349 B.n348 71.676
R1013 B.n342 B.n228 71.676
R1014 B.n341 B.n340 71.676
R1015 B.n334 B.n230 71.676
R1016 B.n333 B.n332 71.676
R1017 B.n326 B.n232 71.676
R1018 B.n325 B.n324 71.676
R1019 B.n318 B.n234 71.676
R1020 B.n317 B.n316 71.676
R1021 B.n310 B.n236 71.676
R1022 B.n309 B.n308 71.676
R1023 B.n302 B.n238 71.676
R1024 B.n301 B.n300 71.676
R1025 B.n294 B.n240 71.676
R1026 B.n293 B.n292 71.676
R1027 B.n286 B.n242 71.676
R1028 B.n285 B.n284 71.676
R1029 B.n278 B.n244 71.676
R1030 B.n277 B.n276 71.676
R1031 B.n270 B.n246 71.676
R1032 B.n269 B.n268 71.676
R1033 B.n262 B.n248 71.676
R1034 B.n261 B.n260 71.676
R1035 B.n254 B.n250 71.676
R1036 B.n253 B.n252 71.676
R1037 B.n470 B.n469 71.676
R1038 B.n464 B.n194 71.676
R1039 B.n462 B.n461 71.676
R1040 B.n457 B.n456 71.676
R1041 B.n454 B.n453 71.676
R1042 B.n449 B.n448 71.676
R1043 B.n446 B.n445 71.676
R1044 B.n441 B.n440 71.676
R1045 B.n438 B.n437 71.676
R1046 B.n433 B.n432 71.676
R1047 B.n430 B.n429 71.676
R1048 B.n425 B.n424 71.676
R1049 B.n422 B.n421 71.676
R1050 B.n417 B.n416 71.676
R1051 B.n414 B.n413 71.676
R1052 B.n409 B.n408 71.676
R1053 B.n406 B.n405 71.676
R1054 B.n401 B.n400 71.676
R1055 B.n398 B.n397 71.676
R1056 B.n393 B.n392 71.676
R1057 B.n390 B.n389 71.676
R1058 B.n385 B.n384 71.676
R1059 B.n382 B.n381 71.676
R1060 B.n377 B.n376 71.676
R1061 B.n374 B.n373 71.676
R1062 B.n368 B.n367 71.676
R1063 B.n365 B.n364 71.676
R1064 B.n360 B.n359 71.676
R1065 B.n357 B.n356 71.676
R1066 B.n351 B.n350 71.676
R1067 B.n348 B.n347 71.676
R1068 B.n343 B.n342 71.676
R1069 B.n340 B.n339 71.676
R1070 B.n335 B.n334 71.676
R1071 B.n332 B.n331 71.676
R1072 B.n327 B.n326 71.676
R1073 B.n324 B.n323 71.676
R1074 B.n319 B.n318 71.676
R1075 B.n316 B.n315 71.676
R1076 B.n311 B.n310 71.676
R1077 B.n308 B.n307 71.676
R1078 B.n303 B.n302 71.676
R1079 B.n300 B.n299 71.676
R1080 B.n295 B.n294 71.676
R1081 B.n292 B.n291 71.676
R1082 B.n287 B.n286 71.676
R1083 B.n284 B.n283 71.676
R1084 B.n279 B.n278 71.676
R1085 B.n276 B.n275 71.676
R1086 B.n271 B.n270 71.676
R1087 B.n268 B.n267 71.676
R1088 B.n263 B.n262 71.676
R1089 B.n260 B.n259 71.676
R1090 B.n255 B.n254 71.676
R1091 B.n252 B.n190 71.676
R1092 B.n916 B.n915 71.676
R1093 B.n916 B.n2 71.676
R1094 B.n100 B.t20 70.5569
R1095 B.n226 B.t12 70.5569
R1096 B.n93 B.t17 70.5372
R1097 B.n220 B.t22 70.5372
R1098 B.n475 B.n191 63.1042
R1099 B.n847 B.n64 63.1042
R1100 B.n94 B.n93 59.5399
R1101 B.n724 B.n100 59.5399
R1102 B.n353 B.n226 59.5399
R1103 B.n371 B.n220 59.5399
R1104 B.n475 B.n187 36.6762
R1105 B.n481 B.n187 36.6762
R1106 B.n481 B.n182 36.6762
R1107 B.n487 B.n182 36.6762
R1108 B.n487 B.n183 36.6762
R1109 B.n493 B.n175 36.6762
R1110 B.n499 B.n175 36.6762
R1111 B.n499 B.n171 36.6762
R1112 B.n505 B.n171 36.6762
R1113 B.n505 B.n166 36.6762
R1114 B.n511 B.n166 36.6762
R1115 B.n511 B.n167 36.6762
R1116 B.n517 B.n158 36.6762
R1117 B.n523 B.n158 36.6762
R1118 B.n523 B.n159 36.6762
R1119 B.n529 B.n150 36.6762
R1120 B.n535 B.n150 36.6762
R1121 B.n535 B.n151 36.6762
R1122 B.n541 B.n143 36.6762
R1123 B.n547 B.n143 36.6762
R1124 B.n547 B.n139 36.6762
R1125 B.n553 B.n139 36.6762
R1126 B.n559 B.n135 36.6762
R1127 B.n559 B.n131 36.6762
R1128 B.n566 B.n131 36.6762
R1129 B.n572 B.n127 36.6762
R1130 B.n572 B.n4 36.6762
R1131 B.n914 B.n4 36.6762
R1132 B.n914 B.n913 36.6762
R1133 B.n913 B.n912 36.6762
R1134 B.n912 B.n8 36.6762
R1135 B.n581 B.n8 36.6762
R1136 B.n905 B.n904 36.6762
R1137 B.n904 B.n903 36.6762
R1138 B.n903 B.n15 36.6762
R1139 B.n897 B.n896 36.6762
R1140 B.n896 B.n895 36.6762
R1141 B.n895 B.n22 36.6762
R1142 B.n889 B.n22 36.6762
R1143 B.n888 B.n887 36.6762
R1144 B.n887 B.n29 36.6762
R1145 B.n881 B.n29 36.6762
R1146 B.n880 B.n879 36.6762
R1147 B.n879 B.n36 36.6762
R1148 B.n873 B.n36 36.6762
R1149 B.n872 B.n871 36.6762
R1150 B.n871 B.n43 36.6762
R1151 B.n865 B.n43 36.6762
R1152 B.n865 B.n864 36.6762
R1153 B.n864 B.n863 36.6762
R1154 B.n863 B.n50 36.6762
R1155 B.n857 B.n50 36.6762
R1156 B.n856 B.n855 36.6762
R1157 B.n855 B.n57 36.6762
R1158 B.n849 B.n57 36.6762
R1159 B.n849 B.n848 36.6762
R1160 B.n848 B.n847 36.6762
R1161 B.n151 B.t6 34.5188
R1162 B.t2 B.n888 34.5188
R1163 B.n473 B.n472 32.3127
R1164 B.n477 B.n189 32.3127
R1165 B.n622 B.n621 32.3127
R1166 B.n845 B.n844 32.3127
R1167 B.n517 B.t1 30.204
R1168 B.n873 B.t4 30.204
R1169 B.n93 B.n92 28.8975
R1170 B.n100 B.n99 28.8975
R1171 B.n226 B.n225 28.8975
R1172 B.n220 B.n219 28.8975
R1173 B.n566 B.t8 25.8892
R1174 B.n905 B.t5 25.8892
R1175 B.t0 B.n135 24.8105
R1176 B.t9 B.n15 24.8105
R1177 B.n183 B.t11 21.5744
R1178 B.t15 B.n856 21.5744
R1179 B.n159 B.t3 20.4957
R1180 B.t7 B.n880 20.4957
R1181 B B.n917 18.0485
R1182 B.n529 B.t3 16.1809
R1183 B.n881 B.t7 16.1809
R1184 B.n493 B.t11 15.1022
R1185 B.n857 B.t15 15.1022
R1186 B.n553 B.t0 11.8662
R1187 B.n897 B.t9 11.8662
R1188 B.t8 B.n127 10.7875
R1189 B.n581 B.t5 10.7875
R1190 B.n473 B.n185 10.6151
R1191 B.n483 B.n185 10.6151
R1192 B.n484 B.n483 10.6151
R1193 B.n485 B.n484 10.6151
R1194 B.n485 B.n177 10.6151
R1195 B.n495 B.n177 10.6151
R1196 B.n496 B.n495 10.6151
R1197 B.n497 B.n496 10.6151
R1198 B.n497 B.n169 10.6151
R1199 B.n507 B.n169 10.6151
R1200 B.n508 B.n507 10.6151
R1201 B.n509 B.n508 10.6151
R1202 B.n509 B.n161 10.6151
R1203 B.n519 B.n161 10.6151
R1204 B.n520 B.n519 10.6151
R1205 B.n521 B.n520 10.6151
R1206 B.n521 B.n153 10.6151
R1207 B.n531 B.n153 10.6151
R1208 B.n532 B.n531 10.6151
R1209 B.n533 B.n532 10.6151
R1210 B.n533 B.n145 10.6151
R1211 B.n543 B.n145 10.6151
R1212 B.n544 B.n543 10.6151
R1213 B.n545 B.n544 10.6151
R1214 B.n545 B.n137 10.6151
R1215 B.n555 B.n137 10.6151
R1216 B.n556 B.n555 10.6151
R1217 B.n557 B.n556 10.6151
R1218 B.n557 B.n129 10.6151
R1219 B.n568 B.n129 10.6151
R1220 B.n569 B.n568 10.6151
R1221 B.n570 B.n569 10.6151
R1222 B.n570 B.n0 10.6151
R1223 B.n472 B.n471 10.6151
R1224 B.n471 B.n193 10.6151
R1225 B.n466 B.n193 10.6151
R1226 B.n466 B.n465 10.6151
R1227 B.n465 B.n195 10.6151
R1228 B.n460 B.n195 10.6151
R1229 B.n460 B.n459 10.6151
R1230 B.n459 B.n458 10.6151
R1231 B.n458 B.n197 10.6151
R1232 B.n452 B.n197 10.6151
R1233 B.n452 B.n451 10.6151
R1234 B.n451 B.n450 10.6151
R1235 B.n450 B.n199 10.6151
R1236 B.n444 B.n199 10.6151
R1237 B.n444 B.n443 10.6151
R1238 B.n443 B.n442 10.6151
R1239 B.n442 B.n201 10.6151
R1240 B.n436 B.n201 10.6151
R1241 B.n436 B.n435 10.6151
R1242 B.n435 B.n434 10.6151
R1243 B.n434 B.n203 10.6151
R1244 B.n428 B.n203 10.6151
R1245 B.n428 B.n427 10.6151
R1246 B.n427 B.n426 10.6151
R1247 B.n426 B.n205 10.6151
R1248 B.n420 B.n205 10.6151
R1249 B.n420 B.n419 10.6151
R1250 B.n419 B.n418 10.6151
R1251 B.n418 B.n207 10.6151
R1252 B.n412 B.n207 10.6151
R1253 B.n412 B.n411 10.6151
R1254 B.n411 B.n410 10.6151
R1255 B.n410 B.n209 10.6151
R1256 B.n404 B.n209 10.6151
R1257 B.n404 B.n403 10.6151
R1258 B.n403 B.n402 10.6151
R1259 B.n402 B.n211 10.6151
R1260 B.n396 B.n211 10.6151
R1261 B.n396 B.n395 10.6151
R1262 B.n395 B.n394 10.6151
R1263 B.n394 B.n213 10.6151
R1264 B.n388 B.n213 10.6151
R1265 B.n388 B.n387 10.6151
R1266 B.n387 B.n386 10.6151
R1267 B.n386 B.n215 10.6151
R1268 B.n380 B.n215 10.6151
R1269 B.n380 B.n379 10.6151
R1270 B.n379 B.n378 10.6151
R1271 B.n378 B.n217 10.6151
R1272 B.n372 B.n217 10.6151
R1273 B.n370 B.n369 10.6151
R1274 B.n369 B.n221 10.6151
R1275 B.n363 B.n221 10.6151
R1276 B.n363 B.n362 10.6151
R1277 B.n362 B.n361 10.6151
R1278 B.n361 B.n223 10.6151
R1279 B.n355 B.n223 10.6151
R1280 B.n355 B.n354 10.6151
R1281 B.n352 B.n227 10.6151
R1282 B.n346 B.n227 10.6151
R1283 B.n346 B.n345 10.6151
R1284 B.n345 B.n344 10.6151
R1285 B.n344 B.n229 10.6151
R1286 B.n338 B.n229 10.6151
R1287 B.n338 B.n337 10.6151
R1288 B.n337 B.n336 10.6151
R1289 B.n336 B.n231 10.6151
R1290 B.n330 B.n231 10.6151
R1291 B.n330 B.n329 10.6151
R1292 B.n329 B.n328 10.6151
R1293 B.n328 B.n233 10.6151
R1294 B.n322 B.n233 10.6151
R1295 B.n322 B.n321 10.6151
R1296 B.n321 B.n320 10.6151
R1297 B.n320 B.n235 10.6151
R1298 B.n314 B.n235 10.6151
R1299 B.n314 B.n313 10.6151
R1300 B.n313 B.n312 10.6151
R1301 B.n312 B.n237 10.6151
R1302 B.n306 B.n237 10.6151
R1303 B.n306 B.n305 10.6151
R1304 B.n305 B.n304 10.6151
R1305 B.n304 B.n239 10.6151
R1306 B.n298 B.n239 10.6151
R1307 B.n298 B.n297 10.6151
R1308 B.n297 B.n296 10.6151
R1309 B.n296 B.n241 10.6151
R1310 B.n290 B.n241 10.6151
R1311 B.n290 B.n289 10.6151
R1312 B.n289 B.n288 10.6151
R1313 B.n288 B.n243 10.6151
R1314 B.n282 B.n243 10.6151
R1315 B.n282 B.n281 10.6151
R1316 B.n281 B.n280 10.6151
R1317 B.n280 B.n245 10.6151
R1318 B.n274 B.n245 10.6151
R1319 B.n274 B.n273 10.6151
R1320 B.n273 B.n272 10.6151
R1321 B.n272 B.n247 10.6151
R1322 B.n266 B.n247 10.6151
R1323 B.n266 B.n265 10.6151
R1324 B.n265 B.n264 10.6151
R1325 B.n264 B.n249 10.6151
R1326 B.n258 B.n249 10.6151
R1327 B.n258 B.n257 10.6151
R1328 B.n257 B.n256 10.6151
R1329 B.n256 B.n251 10.6151
R1330 B.n251 B.n189 10.6151
R1331 B.n478 B.n477 10.6151
R1332 B.n479 B.n478 10.6151
R1333 B.n479 B.n180 10.6151
R1334 B.n489 B.n180 10.6151
R1335 B.n490 B.n489 10.6151
R1336 B.n491 B.n490 10.6151
R1337 B.n491 B.n173 10.6151
R1338 B.n501 B.n173 10.6151
R1339 B.n502 B.n501 10.6151
R1340 B.n503 B.n502 10.6151
R1341 B.n503 B.n164 10.6151
R1342 B.n513 B.n164 10.6151
R1343 B.n514 B.n513 10.6151
R1344 B.n515 B.n514 10.6151
R1345 B.n515 B.n156 10.6151
R1346 B.n525 B.n156 10.6151
R1347 B.n526 B.n525 10.6151
R1348 B.n527 B.n526 10.6151
R1349 B.n527 B.n148 10.6151
R1350 B.n537 B.n148 10.6151
R1351 B.n538 B.n537 10.6151
R1352 B.n539 B.n538 10.6151
R1353 B.n539 B.n141 10.6151
R1354 B.n549 B.n141 10.6151
R1355 B.n550 B.n549 10.6151
R1356 B.n551 B.n550 10.6151
R1357 B.n551 B.n133 10.6151
R1358 B.n561 B.n133 10.6151
R1359 B.n562 B.n561 10.6151
R1360 B.n564 B.n562 10.6151
R1361 B.n564 B.n563 10.6151
R1362 B.n563 B.n125 10.6151
R1363 B.n575 B.n125 10.6151
R1364 B.n576 B.n575 10.6151
R1365 B.n577 B.n576 10.6151
R1366 B.n578 B.n577 10.6151
R1367 B.n579 B.n578 10.6151
R1368 B.n583 B.n579 10.6151
R1369 B.n584 B.n583 10.6151
R1370 B.n585 B.n584 10.6151
R1371 B.n586 B.n585 10.6151
R1372 B.n588 B.n586 10.6151
R1373 B.n589 B.n588 10.6151
R1374 B.n590 B.n589 10.6151
R1375 B.n591 B.n590 10.6151
R1376 B.n593 B.n591 10.6151
R1377 B.n594 B.n593 10.6151
R1378 B.n595 B.n594 10.6151
R1379 B.n596 B.n595 10.6151
R1380 B.n598 B.n596 10.6151
R1381 B.n599 B.n598 10.6151
R1382 B.n600 B.n599 10.6151
R1383 B.n601 B.n600 10.6151
R1384 B.n603 B.n601 10.6151
R1385 B.n604 B.n603 10.6151
R1386 B.n605 B.n604 10.6151
R1387 B.n606 B.n605 10.6151
R1388 B.n608 B.n606 10.6151
R1389 B.n609 B.n608 10.6151
R1390 B.n610 B.n609 10.6151
R1391 B.n611 B.n610 10.6151
R1392 B.n613 B.n611 10.6151
R1393 B.n614 B.n613 10.6151
R1394 B.n615 B.n614 10.6151
R1395 B.n616 B.n615 10.6151
R1396 B.n618 B.n616 10.6151
R1397 B.n619 B.n618 10.6151
R1398 B.n620 B.n619 10.6151
R1399 B.n621 B.n620 10.6151
R1400 B.n909 B.n1 10.6151
R1401 B.n909 B.n908 10.6151
R1402 B.n908 B.n907 10.6151
R1403 B.n907 B.n10 10.6151
R1404 B.n901 B.n10 10.6151
R1405 B.n901 B.n900 10.6151
R1406 B.n900 B.n899 10.6151
R1407 B.n899 B.n17 10.6151
R1408 B.n893 B.n17 10.6151
R1409 B.n893 B.n892 10.6151
R1410 B.n892 B.n891 10.6151
R1411 B.n891 B.n24 10.6151
R1412 B.n885 B.n24 10.6151
R1413 B.n885 B.n884 10.6151
R1414 B.n884 B.n883 10.6151
R1415 B.n883 B.n31 10.6151
R1416 B.n877 B.n31 10.6151
R1417 B.n877 B.n876 10.6151
R1418 B.n876 B.n875 10.6151
R1419 B.n875 B.n38 10.6151
R1420 B.n869 B.n38 10.6151
R1421 B.n869 B.n868 10.6151
R1422 B.n868 B.n867 10.6151
R1423 B.n867 B.n45 10.6151
R1424 B.n861 B.n45 10.6151
R1425 B.n861 B.n860 10.6151
R1426 B.n860 B.n859 10.6151
R1427 B.n859 B.n52 10.6151
R1428 B.n853 B.n52 10.6151
R1429 B.n853 B.n852 10.6151
R1430 B.n852 B.n851 10.6151
R1431 B.n851 B.n59 10.6151
R1432 B.n845 B.n59 10.6151
R1433 B.n844 B.n843 10.6151
R1434 B.n843 B.n66 10.6151
R1435 B.n837 B.n66 10.6151
R1436 B.n837 B.n836 10.6151
R1437 B.n836 B.n835 10.6151
R1438 B.n835 B.n68 10.6151
R1439 B.n829 B.n68 10.6151
R1440 B.n829 B.n828 10.6151
R1441 B.n828 B.n827 10.6151
R1442 B.n827 B.n70 10.6151
R1443 B.n821 B.n70 10.6151
R1444 B.n821 B.n820 10.6151
R1445 B.n820 B.n819 10.6151
R1446 B.n819 B.n72 10.6151
R1447 B.n813 B.n72 10.6151
R1448 B.n813 B.n812 10.6151
R1449 B.n812 B.n811 10.6151
R1450 B.n811 B.n74 10.6151
R1451 B.n805 B.n74 10.6151
R1452 B.n805 B.n804 10.6151
R1453 B.n804 B.n803 10.6151
R1454 B.n803 B.n76 10.6151
R1455 B.n797 B.n76 10.6151
R1456 B.n797 B.n796 10.6151
R1457 B.n796 B.n795 10.6151
R1458 B.n795 B.n78 10.6151
R1459 B.n789 B.n78 10.6151
R1460 B.n789 B.n788 10.6151
R1461 B.n788 B.n787 10.6151
R1462 B.n787 B.n80 10.6151
R1463 B.n781 B.n80 10.6151
R1464 B.n781 B.n780 10.6151
R1465 B.n780 B.n779 10.6151
R1466 B.n779 B.n82 10.6151
R1467 B.n773 B.n82 10.6151
R1468 B.n773 B.n772 10.6151
R1469 B.n772 B.n771 10.6151
R1470 B.n771 B.n84 10.6151
R1471 B.n765 B.n84 10.6151
R1472 B.n765 B.n764 10.6151
R1473 B.n764 B.n763 10.6151
R1474 B.n763 B.n86 10.6151
R1475 B.n757 B.n86 10.6151
R1476 B.n757 B.n756 10.6151
R1477 B.n756 B.n755 10.6151
R1478 B.n755 B.n88 10.6151
R1479 B.n749 B.n88 10.6151
R1480 B.n749 B.n748 10.6151
R1481 B.n748 B.n747 10.6151
R1482 B.n747 B.n90 10.6151
R1483 B.n741 B.n740 10.6151
R1484 B.n740 B.n739 10.6151
R1485 B.n739 B.n95 10.6151
R1486 B.n733 B.n95 10.6151
R1487 B.n733 B.n732 10.6151
R1488 B.n732 B.n731 10.6151
R1489 B.n731 B.n97 10.6151
R1490 B.n725 B.n97 10.6151
R1491 B.n723 B.n722 10.6151
R1492 B.n722 B.n101 10.6151
R1493 B.n716 B.n101 10.6151
R1494 B.n716 B.n715 10.6151
R1495 B.n715 B.n714 10.6151
R1496 B.n714 B.n103 10.6151
R1497 B.n708 B.n103 10.6151
R1498 B.n708 B.n707 10.6151
R1499 B.n707 B.n706 10.6151
R1500 B.n706 B.n105 10.6151
R1501 B.n700 B.n105 10.6151
R1502 B.n700 B.n699 10.6151
R1503 B.n699 B.n698 10.6151
R1504 B.n698 B.n107 10.6151
R1505 B.n692 B.n107 10.6151
R1506 B.n692 B.n691 10.6151
R1507 B.n691 B.n690 10.6151
R1508 B.n690 B.n109 10.6151
R1509 B.n684 B.n109 10.6151
R1510 B.n684 B.n683 10.6151
R1511 B.n683 B.n682 10.6151
R1512 B.n682 B.n111 10.6151
R1513 B.n676 B.n111 10.6151
R1514 B.n676 B.n675 10.6151
R1515 B.n675 B.n674 10.6151
R1516 B.n674 B.n113 10.6151
R1517 B.n668 B.n113 10.6151
R1518 B.n668 B.n667 10.6151
R1519 B.n667 B.n666 10.6151
R1520 B.n666 B.n115 10.6151
R1521 B.n660 B.n115 10.6151
R1522 B.n660 B.n659 10.6151
R1523 B.n659 B.n658 10.6151
R1524 B.n658 B.n117 10.6151
R1525 B.n652 B.n117 10.6151
R1526 B.n652 B.n651 10.6151
R1527 B.n651 B.n650 10.6151
R1528 B.n650 B.n119 10.6151
R1529 B.n644 B.n119 10.6151
R1530 B.n644 B.n643 10.6151
R1531 B.n643 B.n642 10.6151
R1532 B.n642 B.n121 10.6151
R1533 B.n636 B.n121 10.6151
R1534 B.n636 B.n635 10.6151
R1535 B.n635 B.n634 10.6151
R1536 B.n634 B.n123 10.6151
R1537 B.n628 B.n123 10.6151
R1538 B.n628 B.n627 10.6151
R1539 B.n627 B.n626 10.6151
R1540 B.n626 B.n622 10.6151
R1541 B.n917 B.n0 8.11757
R1542 B.n917 B.n1 8.11757
R1543 B.n371 B.n370 6.5566
R1544 B.n354 B.n353 6.5566
R1545 B.n741 B.n94 6.5566
R1546 B.n725 B.n724 6.5566
R1547 B.n167 B.t1 6.47267
R1548 B.t4 B.n872 6.47267
R1549 B.n372 B.n371 4.05904
R1550 B.n353 B.n352 4.05904
R1551 B.n94 B.n90 4.05904
R1552 B.n724 B.n723 4.05904
R1553 B.n541 B.t6 2.15789
R1554 B.n889 B.t2 2.15789
R1555 VP.n14 VP.t5 343.613
R1556 VP.n7 VP.t2 314.132
R1557 VP.n5 VP.t9 314.132
R1558 VP.n3 VP.t7 314.132
R1559 VP.n46 VP.t1 314.132
R1560 VP.n53 VP.t8 314.132
R1561 VP.n30 VP.t4 314.132
R1562 VP.n23 VP.t6 314.132
R1563 VP.n11 VP.t0 314.132
R1564 VP.n13 VP.t3 314.132
R1565 VP.n32 VP.n7 174.581
R1566 VP.n54 VP.n53 174.581
R1567 VP.n31 VP.n30 174.581
R1568 VP.n16 VP.n15 161.3
R1569 VP.n17 VP.n12 161.3
R1570 VP.n19 VP.n18 161.3
R1571 VP.n21 VP.n20 161.3
R1572 VP.n22 VP.n10 161.3
R1573 VP.n25 VP.n24 161.3
R1574 VP.n26 VP.n9 161.3
R1575 VP.n28 VP.n27 161.3
R1576 VP.n29 VP.n8 161.3
R1577 VP.n52 VP.n0 161.3
R1578 VP.n51 VP.n50 161.3
R1579 VP.n49 VP.n1 161.3
R1580 VP.n48 VP.n47 161.3
R1581 VP.n45 VP.n2 161.3
R1582 VP.n44 VP.n43 161.3
R1583 VP.n42 VP.n41 161.3
R1584 VP.n40 VP.n4 161.3
R1585 VP.n39 VP.n38 161.3
R1586 VP.n37 VP.n36 161.3
R1587 VP.n35 VP.n6 161.3
R1588 VP.n34 VP.n33 161.3
R1589 VP.n14 VP.n13 52.1879
R1590 VP.n32 VP.n31 47.5119
R1591 VP.n36 VP.n35 42.0302
R1592 VP.n51 VP.n1 42.0302
R1593 VP.n28 VP.n9 42.0302
R1594 VP.n41 VP.n40 41.0614
R1595 VP.n45 VP.n44 41.0614
R1596 VP.n22 VP.n21 41.0614
R1597 VP.n18 VP.n17 41.0614
R1598 VP.n40 VP.n39 40.0926
R1599 VP.n47 VP.n45 40.0926
R1600 VP.n24 VP.n22 40.0926
R1601 VP.n17 VP.n16 40.0926
R1602 VP.n35 VP.n34 39.1239
R1603 VP.n52 VP.n51 39.1239
R1604 VP.n29 VP.n28 39.1239
R1605 VP.n15 VP.n14 27.1955
R1606 VP.n36 VP.n5 12.7883
R1607 VP.n46 VP.n1 12.7883
R1608 VP.n23 VP.n9 12.7883
R1609 VP.n41 VP.n3 12.2964
R1610 VP.n44 VP.n3 12.2964
R1611 VP.n18 VP.n11 12.2964
R1612 VP.n21 VP.n11 12.2964
R1613 VP.n39 VP.n5 11.8046
R1614 VP.n47 VP.n46 11.8046
R1615 VP.n24 VP.n23 11.8046
R1616 VP.n16 VP.n13 11.8046
R1617 VP.n34 VP.n7 11.3127
R1618 VP.n53 VP.n52 11.3127
R1619 VP.n30 VP.n29 11.3127
R1620 VP.n15 VP.n12 0.189894
R1621 VP.n19 VP.n12 0.189894
R1622 VP.n20 VP.n19 0.189894
R1623 VP.n20 VP.n10 0.189894
R1624 VP.n25 VP.n10 0.189894
R1625 VP.n26 VP.n25 0.189894
R1626 VP.n27 VP.n26 0.189894
R1627 VP.n27 VP.n8 0.189894
R1628 VP.n31 VP.n8 0.189894
R1629 VP.n33 VP.n32 0.189894
R1630 VP.n33 VP.n6 0.189894
R1631 VP.n37 VP.n6 0.189894
R1632 VP.n38 VP.n37 0.189894
R1633 VP.n38 VP.n4 0.189894
R1634 VP.n42 VP.n4 0.189894
R1635 VP.n43 VP.n42 0.189894
R1636 VP.n43 VP.n2 0.189894
R1637 VP.n48 VP.n2 0.189894
R1638 VP.n49 VP.n48 0.189894
R1639 VP.n50 VP.n49 0.189894
R1640 VP.n50 VP.n0 0.189894
R1641 VP.n54 VP.n0 0.189894
R1642 VP VP.n54 0.0516364
R1643 VTAIL.n11 VTAIL.t5 47.8378
R1644 VTAIL.n17 VTAIL.t8 47.8376
R1645 VTAIL.n2 VTAIL.t13 47.8376
R1646 VTAIL.n16 VTAIL.t12 47.8376
R1647 VTAIL.n15 VTAIL.n14 46.5283
R1648 VTAIL.n13 VTAIL.n12 46.5283
R1649 VTAIL.n10 VTAIL.n9 46.5283
R1650 VTAIL.n8 VTAIL.n7 46.5283
R1651 VTAIL.n19 VTAIL.n18 46.528
R1652 VTAIL.n1 VTAIL.n0 46.528
R1653 VTAIL.n4 VTAIL.n3 46.528
R1654 VTAIL.n6 VTAIL.n5 46.528
R1655 VTAIL.n8 VTAIL.n6 27.9703
R1656 VTAIL.n17 VTAIL.n16 26.6858
R1657 VTAIL.n18 VTAIL.t6 1.31002
R1658 VTAIL.n18 VTAIL.t4 1.31002
R1659 VTAIL.n0 VTAIL.t7 1.31002
R1660 VTAIL.n0 VTAIL.t19 1.31002
R1661 VTAIL.n3 VTAIL.t16 1.31002
R1662 VTAIL.n3 VTAIL.t15 1.31002
R1663 VTAIL.n5 VTAIL.t11 1.31002
R1664 VTAIL.n5 VTAIL.t18 1.31002
R1665 VTAIL.n14 VTAIL.t17 1.31002
R1666 VTAIL.n14 VTAIL.t9 1.31002
R1667 VTAIL.n12 VTAIL.t10 1.31002
R1668 VTAIL.n12 VTAIL.t14 1.31002
R1669 VTAIL.n9 VTAIL.t2 1.31002
R1670 VTAIL.n9 VTAIL.t3 1.31002
R1671 VTAIL.n7 VTAIL.t0 1.31002
R1672 VTAIL.n7 VTAIL.t1 1.31002
R1673 VTAIL.n10 VTAIL.n8 1.28498
R1674 VTAIL.n11 VTAIL.n10 1.28498
R1675 VTAIL.n15 VTAIL.n13 1.28498
R1676 VTAIL.n16 VTAIL.n15 1.28498
R1677 VTAIL.n6 VTAIL.n4 1.28498
R1678 VTAIL.n4 VTAIL.n2 1.28498
R1679 VTAIL.n19 VTAIL.n17 1.28498
R1680 VTAIL.n13 VTAIL.n11 1.11257
R1681 VTAIL.n2 VTAIL.n1 1.11257
R1682 VTAIL VTAIL.n1 1.02205
R1683 VTAIL VTAIL.n19 0.263431
R1684 VDD1.n1 VDD1.t4 65.8011
R1685 VDD1.n3 VDD1.t7 65.8008
R1686 VDD1.n5 VDD1.n4 64.1148
R1687 VDD1.n1 VDD1.n0 63.2071
R1688 VDD1.n7 VDD1.n6 63.2069
R1689 VDD1.n3 VDD1.n2 63.2068
R1690 VDD1.n7 VDD1.n5 44.0763
R1691 VDD1.n6 VDD1.t3 1.31002
R1692 VDD1.n6 VDD1.t5 1.31002
R1693 VDD1.n0 VDD1.t6 1.31002
R1694 VDD1.n0 VDD1.t9 1.31002
R1695 VDD1.n4 VDD1.t8 1.31002
R1696 VDD1.n4 VDD1.t1 1.31002
R1697 VDD1.n2 VDD1.t0 1.31002
R1698 VDD1.n2 VDD1.t2 1.31002
R1699 VDD1 VDD1.n7 0.905672
R1700 VDD1 VDD1.n1 0.37981
R1701 VDD1.n5 VDD1.n3 0.266275
R1702 VN.n6 VN.t5 343.613
R1703 VN.n31 VN.t4 343.613
R1704 VN.n5 VN.t9 314.132
R1705 VN.n3 VN.t3 314.132
R1706 VN.n15 VN.t7 314.132
R1707 VN.n22 VN.t1 314.132
R1708 VN.n30 VN.t2 314.132
R1709 VN.n28 VN.t0 314.132
R1710 VN.n27 VN.t8 314.132
R1711 VN.n46 VN.t6 314.132
R1712 VN.n23 VN.n22 174.581
R1713 VN.n47 VN.n46 174.581
R1714 VN.n45 VN.n24 161.3
R1715 VN.n44 VN.n43 161.3
R1716 VN.n42 VN.n25 161.3
R1717 VN.n41 VN.n40 161.3
R1718 VN.n39 VN.n26 161.3
R1719 VN.n38 VN.n37 161.3
R1720 VN.n36 VN.n35 161.3
R1721 VN.n34 VN.n29 161.3
R1722 VN.n33 VN.n32 161.3
R1723 VN.n21 VN.n0 161.3
R1724 VN.n20 VN.n19 161.3
R1725 VN.n18 VN.n1 161.3
R1726 VN.n17 VN.n16 161.3
R1727 VN.n14 VN.n2 161.3
R1728 VN.n13 VN.n12 161.3
R1729 VN.n11 VN.n10 161.3
R1730 VN.n9 VN.n4 161.3
R1731 VN.n8 VN.n7 161.3
R1732 VN.n6 VN.n5 52.1879
R1733 VN.n31 VN.n30 52.1879
R1734 VN VN.n47 47.8925
R1735 VN.n20 VN.n1 42.0302
R1736 VN.n44 VN.n25 42.0302
R1737 VN.n10 VN.n9 41.0614
R1738 VN.n14 VN.n13 41.0614
R1739 VN.n35 VN.n34 41.0614
R1740 VN.n39 VN.n38 41.0614
R1741 VN.n9 VN.n8 40.0926
R1742 VN.n16 VN.n14 40.0926
R1743 VN.n34 VN.n33 40.0926
R1744 VN.n40 VN.n39 40.0926
R1745 VN.n21 VN.n20 39.1239
R1746 VN.n45 VN.n44 39.1239
R1747 VN.n32 VN.n31 27.1955
R1748 VN.n7 VN.n6 27.1955
R1749 VN.n15 VN.n1 12.7883
R1750 VN.n27 VN.n25 12.7883
R1751 VN.n10 VN.n3 12.2964
R1752 VN.n13 VN.n3 12.2964
R1753 VN.n38 VN.n28 12.2964
R1754 VN.n35 VN.n28 12.2964
R1755 VN.n8 VN.n5 11.8046
R1756 VN.n16 VN.n15 11.8046
R1757 VN.n33 VN.n30 11.8046
R1758 VN.n40 VN.n27 11.8046
R1759 VN.n22 VN.n21 11.3127
R1760 VN.n46 VN.n45 11.3127
R1761 VN.n47 VN.n24 0.189894
R1762 VN.n43 VN.n24 0.189894
R1763 VN.n43 VN.n42 0.189894
R1764 VN.n42 VN.n41 0.189894
R1765 VN.n41 VN.n26 0.189894
R1766 VN.n37 VN.n26 0.189894
R1767 VN.n37 VN.n36 0.189894
R1768 VN.n36 VN.n29 0.189894
R1769 VN.n32 VN.n29 0.189894
R1770 VN.n7 VN.n4 0.189894
R1771 VN.n11 VN.n4 0.189894
R1772 VN.n12 VN.n11 0.189894
R1773 VN.n12 VN.n2 0.189894
R1774 VN.n17 VN.n2 0.189894
R1775 VN.n18 VN.n17 0.189894
R1776 VN.n19 VN.n18 0.189894
R1777 VN.n19 VN.n0 0.189894
R1778 VN.n23 VN.n0 0.189894
R1779 VN VN.n23 0.0516364
R1780 VDD2.n1 VDD2.t4 65.8008
R1781 VDD2.n4 VDD2.t3 64.5166
R1782 VDD2.n3 VDD2.n2 64.1148
R1783 VDD2 VDD2.n7 64.1121
R1784 VDD2.n6 VDD2.n5 63.2071
R1785 VDD2.n1 VDD2.n0 63.2068
R1786 VDD2.n4 VDD2.n3 42.8511
R1787 VDD2.n7 VDD2.t7 1.31002
R1788 VDD2.n7 VDD2.t5 1.31002
R1789 VDD2.n5 VDD2.t1 1.31002
R1790 VDD2.n5 VDD2.t9 1.31002
R1791 VDD2.n2 VDD2.t2 1.31002
R1792 VDD2.n2 VDD2.t8 1.31002
R1793 VDD2.n0 VDD2.t0 1.31002
R1794 VDD2.n0 VDD2.t6 1.31002
R1795 VDD2.n6 VDD2.n4 1.28498
R1796 VDD2 VDD2.n6 0.37981
R1797 VDD2.n3 VDD2.n1 0.266275
C0 VN VDD1 0.149971f
C1 VTAIL VDD1 13.955701f
C2 VDD1 VP 10.7769f
C3 VTAIL VN 10.4487f
C4 VDD2 VDD1 1.25209f
C5 VN VP 6.85325f
C6 VTAIL VP 10.4633f
C7 VDD2 VN 10.5317f
C8 VDD2 VTAIL 13.993099f
C9 VDD2 VP 0.400383f
C10 VDD2 B 6.058437f
C11 VDD1 B 6.018214f
C12 VTAIL B 8.137722f
C13 VN B 11.79635f
C14 VP B 9.935272f
C15 VDD2.t4 B 3.16405f
C16 VDD2.t0 B 0.273135f
C17 VDD2.t6 B 0.273135f
C18 VDD2.n0 B 2.47209f
C19 VDD2.n1 B 0.642956f
C20 VDD2.t2 B 0.273135f
C21 VDD2.t8 B 0.273135f
C22 VDD2.n2 B 2.47713f
C23 VDD2.n3 B 2.13701f
C24 VDD2.t3 B 3.15725f
C25 VDD2.n4 B 2.5626f
C26 VDD2.t1 B 0.273135f
C27 VDD2.t9 B 0.273135f
C28 VDD2.n5 B 2.47209f
C29 VDD2.n6 B 0.307552f
C30 VDD2.t7 B 0.273135f
C31 VDD2.t5 B 0.273135f
C32 VDD2.n7 B 2.4771f
C33 VN.n0 B 0.033909f
C34 VN.t1 B 1.63f
C35 VN.n1 B 0.051587f
C36 VN.n2 B 0.033909f
C37 VN.t3 B 1.63f
C38 VN.n3 B 0.586625f
C39 VN.n4 B 0.033909f
C40 VN.t9 B 1.63f
C41 VN.n5 B 0.634987f
C42 VN.t5 B 1.68859f
C43 VN.n6 B 0.662918f
C44 VN.n7 B 0.174667f
C45 VN.n8 B 0.05106f
C46 VN.n9 B 0.027398f
C47 VN.n10 B 0.051344f
C48 VN.n11 B 0.033909f
C49 VN.n12 B 0.033909f
C50 VN.n13 B 0.051344f
C51 VN.n14 B 0.027398f
C52 VN.t7 B 1.63f
C53 VN.n15 B 0.586625f
C54 VN.n16 B 0.05106f
C55 VN.n17 B 0.033909f
C56 VN.n18 B 0.033909f
C57 VN.n19 B 0.033909f
C58 VN.n20 B 0.027485f
C59 VN.n21 B 0.050731f
C60 VN.n22 B 0.638413f
C61 VN.n23 B 0.030542f
C62 VN.n24 B 0.033909f
C63 VN.t6 B 1.63f
C64 VN.n25 B 0.051587f
C65 VN.n26 B 0.033909f
C66 VN.t8 B 1.63f
C67 VN.n27 B 0.586625f
C68 VN.t0 B 1.63f
C69 VN.n28 B 0.586625f
C70 VN.n29 B 0.033909f
C71 VN.t2 B 1.63f
C72 VN.n30 B 0.634987f
C73 VN.t4 B 1.68859f
C74 VN.n31 B 0.662918f
C75 VN.n32 B 0.174667f
C76 VN.n33 B 0.05106f
C77 VN.n34 B 0.027398f
C78 VN.n35 B 0.051344f
C79 VN.n36 B 0.033909f
C80 VN.n37 B 0.033909f
C81 VN.n38 B 0.051344f
C82 VN.n39 B 0.027398f
C83 VN.n40 B 0.05106f
C84 VN.n41 B 0.033909f
C85 VN.n42 B 0.033909f
C86 VN.n43 B 0.033909f
C87 VN.n44 B 0.027485f
C88 VN.n45 B 0.050731f
C89 VN.n46 B 0.638413f
C90 VN.n47 B 1.7319f
C91 VDD1.t4 B 3.1918f
C92 VDD1.t6 B 0.27553f
C93 VDD1.t9 B 0.27553f
C94 VDD1.n0 B 2.49377f
C95 VDD1.n1 B 0.655014f
C96 VDD1.t7 B 3.1918f
C97 VDD1.t0 B 0.27553f
C98 VDD1.t2 B 0.27553f
C99 VDD1.n2 B 2.49376f
C100 VDD1.n3 B 0.648594f
C101 VDD1.t8 B 0.27553f
C102 VDD1.t1 B 0.27553f
C103 VDD1.n4 B 2.49885f
C104 VDD1.n5 B 2.23807f
C105 VDD1.t3 B 0.27553f
C106 VDD1.t5 B 0.27553f
C107 VDD1.n6 B 2.49376f
C108 VDD1.n7 B 2.59491f
C109 VTAIL.t7 B 0.288139f
C110 VTAIL.t19 B 0.288139f
C111 VTAIL.n0 B 2.53957f
C112 VTAIL.n1 B 0.396493f
C113 VTAIL.t13 B 3.24226f
C114 VTAIL.n2 B 0.500068f
C115 VTAIL.t16 B 0.288139f
C116 VTAIL.t15 B 0.288139f
C117 VTAIL.n3 B 2.53957f
C118 VTAIL.n4 B 0.430322f
C119 VTAIL.t11 B 0.288139f
C120 VTAIL.t18 B 0.288139f
C121 VTAIL.n5 B 2.53957f
C122 VTAIL.n6 B 1.87057f
C123 VTAIL.t0 B 0.288139f
C124 VTAIL.t1 B 0.288139f
C125 VTAIL.n7 B 2.53957f
C126 VTAIL.n8 B 1.87056f
C127 VTAIL.t2 B 0.288139f
C128 VTAIL.t3 B 0.288139f
C129 VTAIL.n9 B 2.53957f
C130 VTAIL.n10 B 0.430319f
C131 VTAIL.t5 B 3.24226f
C132 VTAIL.n11 B 0.500065f
C133 VTAIL.t10 B 0.288139f
C134 VTAIL.t14 B 0.288139f
C135 VTAIL.n12 B 2.53957f
C136 VTAIL.n13 B 0.416921f
C137 VTAIL.t17 B 0.288139f
C138 VTAIL.t9 B 0.288139f
C139 VTAIL.n14 B 2.53957f
C140 VTAIL.n15 B 0.430319f
C141 VTAIL.t12 B 3.24226f
C142 VTAIL.n16 B 1.8539f
C143 VTAIL.t8 B 3.24226f
C144 VTAIL.n17 B 1.8539f
C145 VTAIL.t6 B 0.288139f
C146 VTAIL.t4 B 0.288139f
C147 VTAIL.n18 B 2.53957f
C148 VTAIL.n19 B 0.350942f
C149 VP.n0 B 0.034456f
C150 VP.t8 B 1.65629f
C151 VP.n1 B 0.052419f
C152 VP.n2 B 0.034456f
C153 VP.t7 B 1.65629f
C154 VP.n3 B 0.596087f
C155 VP.n4 B 0.034456f
C156 VP.t9 B 1.65629f
C157 VP.n5 B 0.596087f
C158 VP.n6 B 0.034456f
C159 VP.t2 B 1.65629f
C160 VP.n7 B 0.648711f
C161 VP.n8 B 0.034456f
C162 VP.t4 B 1.65629f
C163 VP.n9 B 0.052419f
C164 VP.n10 B 0.034456f
C165 VP.t0 B 1.65629f
C166 VP.n11 B 0.596087f
C167 VP.n12 B 0.034456f
C168 VP.t3 B 1.65629f
C169 VP.n13 B 0.64523f
C170 VP.t5 B 1.71583f
C171 VP.n14 B 0.673611f
C172 VP.n15 B 0.177485f
C173 VP.n16 B 0.051883f
C174 VP.n17 B 0.02784f
C175 VP.n18 B 0.052173f
C176 VP.n19 B 0.034456f
C177 VP.n20 B 0.034456f
C178 VP.n21 B 0.052173f
C179 VP.n22 B 0.02784f
C180 VP.t6 B 1.65629f
C181 VP.n23 B 0.596087f
C182 VP.n24 B 0.051883f
C183 VP.n25 B 0.034456f
C184 VP.n26 B 0.034456f
C185 VP.n27 B 0.034456f
C186 VP.n28 B 0.027928f
C187 VP.n29 B 0.051549f
C188 VP.n30 B 0.648711f
C189 VP.n31 B 1.73738f
C190 VP.n32 B 1.76352f
C191 VP.n33 B 0.034456f
C192 VP.n34 B 0.051549f
C193 VP.n35 B 0.027928f
C194 VP.n36 B 0.052419f
C195 VP.n37 B 0.034456f
C196 VP.n38 B 0.034456f
C197 VP.n39 B 0.051883f
C198 VP.n40 B 0.02784f
C199 VP.n41 B 0.052173f
C200 VP.n42 B 0.034456f
C201 VP.n43 B 0.034456f
C202 VP.n44 B 0.052173f
C203 VP.n45 B 0.02784f
C204 VP.t1 B 1.65629f
C205 VP.n46 B 0.596087f
C206 VP.n47 B 0.051883f
C207 VP.n48 B 0.034456f
C208 VP.n49 B 0.034456f
C209 VP.n50 B 0.034456f
C210 VP.n51 B 0.027928f
C211 VP.n52 B 0.051549f
C212 VP.n53 B 0.648711f
C213 VP.n54 B 0.031035f
.ends

