* NGSPICE file created from diff_pair_sample_1514.ext - technology: sky130A

.subckt diff_pair_sample_1514 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=0 ps=0 w=18.44 l=2.23
X1 VTAIL.t14 VN.t0 VDD2.t7 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X2 VTAIL.t13 VN.t1 VDD2.t1 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X3 VTAIL.t2 VP.t0 VDD1.t7 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X4 VTAIL.t6 VP.t1 VDD1.t6 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=3.0426 ps=18.77 w=18.44 l=2.23
X5 B.t8 B.t6 B.t7 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=0 ps=0 w=18.44 l=2.23
X6 B.t5 B.t3 B.t4 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=0 ps=0 w=18.44 l=2.23
X7 VDD2.t2 VN.t2 VTAIL.t12 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X8 VTAIL.t1 VP.t2 VDD1.t5 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=3.0426 ps=18.77 w=18.44 l=2.23
X9 VTAIL.t11 VN.t3 VDD2.t4 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=3.0426 ps=18.77 w=18.44 l=2.23
X10 VDD1.t4 VP.t3 VTAIL.t5 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=7.1916 ps=37.66 w=18.44 l=2.23
X11 VDD2.t6 VN.t4 VTAIL.t10 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=7.1916 ps=37.66 w=18.44 l=2.23
X12 B.t2 B.t0 B.t1 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=0 ps=0 w=18.44 l=2.23
X13 VTAIL.t15 VP.t4 VDD1.t3 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X14 VTAIL.t9 VN.t5 VDD2.t3 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=7.1916 pd=37.66 as=3.0426 ps=18.77 w=18.44 l=2.23
X15 VDD2.t5 VN.t6 VTAIL.t8 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=7.1916 ps=37.66 w=18.44 l=2.23
X16 VDD1.t2 VP.t5 VTAIL.t4 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X17 VDD1.t1 VP.t6 VTAIL.t0 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X18 VDD2.t0 VN.t7 VTAIL.t7 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=3.0426 ps=18.77 w=18.44 l=2.23
X19 VDD1.t0 VP.t7 VTAIL.t3 w_n3530_n4656# sky130_fd_pr__pfet_01v8 ad=3.0426 pd=18.77 as=7.1916 ps=37.66 w=18.44 l=2.23
R0 B.n495 B.n140 585
R1 B.n494 B.n493 585
R2 B.n492 B.n141 585
R3 B.n491 B.n490 585
R4 B.n489 B.n142 585
R5 B.n488 B.n487 585
R6 B.n486 B.n143 585
R7 B.n485 B.n484 585
R8 B.n483 B.n144 585
R9 B.n482 B.n481 585
R10 B.n480 B.n145 585
R11 B.n479 B.n478 585
R12 B.n477 B.n146 585
R13 B.n476 B.n475 585
R14 B.n474 B.n147 585
R15 B.n473 B.n472 585
R16 B.n471 B.n148 585
R17 B.n470 B.n469 585
R18 B.n468 B.n149 585
R19 B.n467 B.n466 585
R20 B.n465 B.n150 585
R21 B.n464 B.n463 585
R22 B.n462 B.n151 585
R23 B.n461 B.n460 585
R24 B.n459 B.n152 585
R25 B.n458 B.n457 585
R26 B.n456 B.n153 585
R27 B.n455 B.n454 585
R28 B.n453 B.n154 585
R29 B.n452 B.n451 585
R30 B.n450 B.n155 585
R31 B.n449 B.n448 585
R32 B.n447 B.n156 585
R33 B.n446 B.n445 585
R34 B.n444 B.n157 585
R35 B.n443 B.n442 585
R36 B.n441 B.n158 585
R37 B.n440 B.n439 585
R38 B.n438 B.n159 585
R39 B.n437 B.n436 585
R40 B.n435 B.n160 585
R41 B.n434 B.n433 585
R42 B.n432 B.n161 585
R43 B.n431 B.n430 585
R44 B.n429 B.n162 585
R45 B.n428 B.n427 585
R46 B.n426 B.n163 585
R47 B.n425 B.n424 585
R48 B.n423 B.n164 585
R49 B.n422 B.n421 585
R50 B.n420 B.n165 585
R51 B.n419 B.n418 585
R52 B.n417 B.n166 585
R53 B.n416 B.n415 585
R54 B.n414 B.n167 585
R55 B.n413 B.n412 585
R56 B.n411 B.n168 585
R57 B.n410 B.n409 585
R58 B.n408 B.n169 585
R59 B.n407 B.n406 585
R60 B.n405 B.n170 585
R61 B.n404 B.n403 585
R62 B.n399 B.n171 585
R63 B.n398 B.n397 585
R64 B.n396 B.n172 585
R65 B.n395 B.n394 585
R66 B.n393 B.n173 585
R67 B.n392 B.n391 585
R68 B.n390 B.n174 585
R69 B.n389 B.n388 585
R70 B.n386 B.n175 585
R71 B.n385 B.n384 585
R72 B.n383 B.n178 585
R73 B.n382 B.n381 585
R74 B.n380 B.n179 585
R75 B.n379 B.n378 585
R76 B.n377 B.n180 585
R77 B.n376 B.n375 585
R78 B.n374 B.n181 585
R79 B.n373 B.n372 585
R80 B.n371 B.n182 585
R81 B.n370 B.n369 585
R82 B.n368 B.n183 585
R83 B.n367 B.n366 585
R84 B.n365 B.n184 585
R85 B.n364 B.n363 585
R86 B.n362 B.n185 585
R87 B.n361 B.n360 585
R88 B.n359 B.n186 585
R89 B.n358 B.n357 585
R90 B.n356 B.n187 585
R91 B.n355 B.n354 585
R92 B.n353 B.n188 585
R93 B.n352 B.n351 585
R94 B.n350 B.n189 585
R95 B.n349 B.n348 585
R96 B.n347 B.n190 585
R97 B.n346 B.n345 585
R98 B.n344 B.n191 585
R99 B.n343 B.n342 585
R100 B.n341 B.n192 585
R101 B.n340 B.n339 585
R102 B.n338 B.n193 585
R103 B.n337 B.n336 585
R104 B.n335 B.n194 585
R105 B.n334 B.n333 585
R106 B.n332 B.n195 585
R107 B.n331 B.n330 585
R108 B.n329 B.n196 585
R109 B.n328 B.n327 585
R110 B.n326 B.n197 585
R111 B.n325 B.n324 585
R112 B.n323 B.n198 585
R113 B.n322 B.n321 585
R114 B.n320 B.n199 585
R115 B.n319 B.n318 585
R116 B.n317 B.n200 585
R117 B.n316 B.n315 585
R118 B.n314 B.n201 585
R119 B.n313 B.n312 585
R120 B.n311 B.n202 585
R121 B.n310 B.n309 585
R122 B.n308 B.n203 585
R123 B.n307 B.n306 585
R124 B.n305 B.n204 585
R125 B.n304 B.n303 585
R126 B.n302 B.n205 585
R127 B.n301 B.n300 585
R128 B.n299 B.n206 585
R129 B.n298 B.n297 585
R130 B.n296 B.n207 585
R131 B.n497 B.n496 585
R132 B.n498 B.n139 585
R133 B.n500 B.n499 585
R134 B.n501 B.n138 585
R135 B.n503 B.n502 585
R136 B.n504 B.n137 585
R137 B.n506 B.n505 585
R138 B.n507 B.n136 585
R139 B.n509 B.n508 585
R140 B.n510 B.n135 585
R141 B.n512 B.n511 585
R142 B.n513 B.n134 585
R143 B.n515 B.n514 585
R144 B.n516 B.n133 585
R145 B.n518 B.n517 585
R146 B.n519 B.n132 585
R147 B.n521 B.n520 585
R148 B.n522 B.n131 585
R149 B.n524 B.n523 585
R150 B.n525 B.n130 585
R151 B.n527 B.n526 585
R152 B.n528 B.n129 585
R153 B.n530 B.n529 585
R154 B.n531 B.n128 585
R155 B.n533 B.n532 585
R156 B.n534 B.n127 585
R157 B.n536 B.n535 585
R158 B.n537 B.n126 585
R159 B.n539 B.n538 585
R160 B.n540 B.n125 585
R161 B.n542 B.n541 585
R162 B.n543 B.n124 585
R163 B.n545 B.n544 585
R164 B.n546 B.n123 585
R165 B.n548 B.n547 585
R166 B.n549 B.n122 585
R167 B.n551 B.n550 585
R168 B.n552 B.n121 585
R169 B.n554 B.n553 585
R170 B.n555 B.n120 585
R171 B.n557 B.n556 585
R172 B.n558 B.n119 585
R173 B.n560 B.n559 585
R174 B.n561 B.n118 585
R175 B.n563 B.n562 585
R176 B.n564 B.n117 585
R177 B.n566 B.n565 585
R178 B.n567 B.n116 585
R179 B.n569 B.n568 585
R180 B.n570 B.n115 585
R181 B.n572 B.n571 585
R182 B.n573 B.n114 585
R183 B.n575 B.n574 585
R184 B.n576 B.n113 585
R185 B.n578 B.n577 585
R186 B.n579 B.n112 585
R187 B.n581 B.n580 585
R188 B.n582 B.n111 585
R189 B.n584 B.n583 585
R190 B.n585 B.n110 585
R191 B.n587 B.n586 585
R192 B.n588 B.n109 585
R193 B.n590 B.n589 585
R194 B.n591 B.n108 585
R195 B.n593 B.n592 585
R196 B.n594 B.n107 585
R197 B.n596 B.n595 585
R198 B.n597 B.n106 585
R199 B.n599 B.n598 585
R200 B.n600 B.n105 585
R201 B.n602 B.n601 585
R202 B.n603 B.n104 585
R203 B.n605 B.n604 585
R204 B.n606 B.n103 585
R205 B.n608 B.n607 585
R206 B.n609 B.n102 585
R207 B.n611 B.n610 585
R208 B.n612 B.n101 585
R209 B.n614 B.n613 585
R210 B.n615 B.n100 585
R211 B.n617 B.n616 585
R212 B.n618 B.n99 585
R213 B.n620 B.n619 585
R214 B.n621 B.n98 585
R215 B.n623 B.n622 585
R216 B.n624 B.n97 585
R217 B.n626 B.n625 585
R218 B.n627 B.n96 585
R219 B.n629 B.n628 585
R220 B.n630 B.n95 585
R221 B.n632 B.n631 585
R222 B.n633 B.n94 585
R223 B.n832 B.n831 585
R224 B.n830 B.n25 585
R225 B.n829 B.n828 585
R226 B.n827 B.n26 585
R227 B.n826 B.n825 585
R228 B.n824 B.n27 585
R229 B.n823 B.n822 585
R230 B.n821 B.n28 585
R231 B.n820 B.n819 585
R232 B.n818 B.n29 585
R233 B.n817 B.n816 585
R234 B.n815 B.n30 585
R235 B.n814 B.n813 585
R236 B.n812 B.n31 585
R237 B.n811 B.n810 585
R238 B.n809 B.n32 585
R239 B.n808 B.n807 585
R240 B.n806 B.n33 585
R241 B.n805 B.n804 585
R242 B.n803 B.n34 585
R243 B.n802 B.n801 585
R244 B.n800 B.n35 585
R245 B.n799 B.n798 585
R246 B.n797 B.n36 585
R247 B.n796 B.n795 585
R248 B.n794 B.n37 585
R249 B.n793 B.n792 585
R250 B.n791 B.n38 585
R251 B.n790 B.n789 585
R252 B.n788 B.n39 585
R253 B.n787 B.n786 585
R254 B.n785 B.n40 585
R255 B.n784 B.n783 585
R256 B.n782 B.n41 585
R257 B.n781 B.n780 585
R258 B.n779 B.n42 585
R259 B.n778 B.n777 585
R260 B.n776 B.n43 585
R261 B.n775 B.n774 585
R262 B.n773 B.n44 585
R263 B.n772 B.n771 585
R264 B.n770 B.n45 585
R265 B.n769 B.n768 585
R266 B.n767 B.n46 585
R267 B.n766 B.n765 585
R268 B.n764 B.n47 585
R269 B.n763 B.n762 585
R270 B.n761 B.n48 585
R271 B.n760 B.n759 585
R272 B.n758 B.n49 585
R273 B.n757 B.n756 585
R274 B.n755 B.n50 585
R275 B.n754 B.n753 585
R276 B.n752 B.n51 585
R277 B.n751 B.n750 585
R278 B.n749 B.n52 585
R279 B.n748 B.n747 585
R280 B.n746 B.n53 585
R281 B.n745 B.n744 585
R282 B.n743 B.n54 585
R283 B.n742 B.n741 585
R284 B.n739 B.n55 585
R285 B.n738 B.n737 585
R286 B.n736 B.n58 585
R287 B.n735 B.n734 585
R288 B.n733 B.n59 585
R289 B.n732 B.n731 585
R290 B.n730 B.n60 585
R291 B.n729 B.n728 585
R292 B.n727 B.n61 585
R293 B.n725 B.n724 585
R294 B.n723 B.n64 585
R295 B.n722 B.n721 585
R296 B.n720 B.n65 585
R297 B.n719 B.n718 585
R298 B.n717 B.n66 585
R299 B.n716 B.n715 585
R300 B.n714 B.n67 585
R301 B.n713 B.n712 585
R302 B.n711 B.n68 585
R303 B.n710 B.n709 585
R304 B.n708 B.n69 585
R305 B.n707 B.n706 585
R306 B.n705 B.n70 585
R307 B.n704 B.n703 585
R308 B.n702 B.n71 585
R309 B.n701 B.n700 585
R310 B.n699 B.n72 585
R311 B.n698 B.n697 585
R312 B.n696 B.n73 585
R313 B.n695 B.n694 585
R314 B.n693 B.n74 585
R315 B.n692 B.n691 585
R316 B.n690 B.n75 585
R317 B.n689 B.n688 585
R318 B.n687 B.n76 585
R319 B.n686 B.n685 585
R320 B.n684 B.n77 585
R321 B.n683 B.n682 585
R322 B.n681 B.n78 585
R323 B.n680 B.n679 585
R324 B.n678 B.n79 585
R325 B.n677 B.n676 585
R326 B.n675 B.n80 585
R327 B.n674 B.n673 585
R328 B.n672 B.n81 585
R329 B.n671 B.n670 585
R330 B.n669 B.n82 585
R331 B.n668 B.n667 585
R332 B.n666 B.n83 585
R333 B.n665 B.n664 585
R334 B.n663 B.n84 585
R335 B.n662 B.n661 585
R336 B.n660 B.n85 585
R337 B.n659 B.n658 585
R338 B.n657 B.n86 585
R339 B.n656 B.n655 585
R340 B.n654 B.n87 585
R341 B.n653 B.n652 585
R342 B.n651 B.n88 585
R343 B.n650 B.n649 585
R344 B.n648 B.n89 585
R345 B.n647 B.n646 585
R346 B.n645 B.n90 585
R347 B.n644 B.n643 585
R348 B.n642 B.n91 585
R349 B.n641 B.n640 585
R350 B.n639 B.n92 585
R351 B.n638 B.n637 585
R352 B.n636 B.n93 585
R353 B.n635 B.n634 585
R354 B.n833 B.n24 585
R355 B.n835 B.n834 585
R356 B.n836 B.n23 585
R357 B.n838 B.n837 585
R358 B.n839 B.n22 585
R359 B.n841 B.n840 585
R360 B.n842 B.n21 585
R361 B.n844 B.n843 585
R362 B.n845 B.n20 585
R363 B.n847 B.n846 585
R364 B.n848 B.n19 585
R365 B.n850 B.n849 585
R366 B.n851 B.n18 585
R367 B.n853 B.n852 585
R368 B.n854 B.n17 585
R369 B.n856 B.n855 585
R370 B.n857 B.n16 585
R371 B.n859 B.n858 585
R372 B.n860 B.n15 585
R373 B.n862 B.n861 585
R374 B.n863 B.n14 585
R375 B.n865 B.n864 585
R376 B.n866 B.n13 585
R377 B.n868 B.n867 585
R378 B.n869 B.n12 585
R379 B.n871 B.n870 585
R380 B.n872 B.n11 585
R381 B.n874 B.n873 585
R382 B.n875 B.n10 585
R383 B.n877 B.n876 585
R384 B.n878 B.n9 585
R385 B.n880 B.n879 585
R386 B.n881 B.n8 585
R387 B.n883 B.n882 585
R388 B.n884 B.n7 585
R389 B.n886 B.n885 585
R390 B.n887 B.n6 585
R391 B.n889 B.n888 585
R392 B.n890 B.n5 585
R393 B.n892 B.n891 585
R394 B.n893 B.n4 585
R395 B.n895 B.n894 585
R396 B.n896 B.n3 585
R397 B.n898 B.n897 585
R398 B.n899 B.n0 585
R399 B.n2 B.n1 585
R400 B.n230 B.n229 585
R401 B.n232 B.n231 585
R402 B.n233 B.n228 585
R403 B.n235 B.n234 585
R404 B.n236 B.n227 585
R405 B.n238 B.n237 585
R406 B.n239 B.n226 585
R407 B.n241 B.n240 585
R408 B.n242 B.n225 585
R409 B.n244 B.n243 585
R410 B.n245 B.n224 585
R411 B.n247 B.n246 585
R412 B.n248 B.n223 585
R413 B.n250 B.n249 585
R414 B.n251 B.n222 585
R415 B.n253 B.n252 585
R416 B.n254 B.n221 585
R417 B.n256 B.n255 585
R418 B.n257 B.n220 585
R419 B.n259 B.n258 585
R420 B.n260 B.n219 585
R421 B.n262 B.n261 585
R422 B.n263 B.n218 585
R423 B.n265 B.n264 585
R424 B.n266 B.n217 585
R425 B.n268 B.n267 585
R426 B.n269 B.n216 585
R427 B.n271 B.n270 585
R428 B.n272 B.n215 585
R429 B.n274 B.n273 585
R430 B.n275 B.n214 585
R431 B.n277 B.n276 585
R432 B.n278 B.n213 585
R433 B.n280 B.n279 585
R434 B.n281 B.n212 585
R435 B.n283 B.n282 585
R436 B.n284 B.n211 585
R437 B.n286 B.n285 585
R438 B.n287 B.n210 585
R439 B.n289 B.n288 585
R440 B.n290 B.n209 585
R441 B.n292 B.n291 585
R442 B.n293 B.n208 585
R443 B.n295 B.n294 585
R444 B.n294 B.n207 516.524
R445 B.n496 B.n495 516.524
R446 B.n634 B.n633 516.524
R447 B.n833 B.n832 516.524
R448 B.n176 B.t9 406.695
R449 B.n400 B.t3 406.695
R450 B.n62 B.t6 406.695
R451 B.n56 B.t0 406.695
R452 B.n901 B.n900 256.663
R453 B.n900 B.n899 235.042
R454 B.n900 B.n2 235.042
R455 B.n298 B.n207 163.367
R456 B.n299 B.n298 163.367
R457 B.n300 B.n299 163.367
R458 B.n300 B.n205 163.367
R459 B.n304 B.n205 163.367
R460 B.n305 B.n304 163.367
R461 B.n306 B.n305 163.367
R462 B.n306 B.n203 163.367
R463 B.n310 B.n203 163.367
R464 B.n311 B.n310 163.367
R465 B.n312 B.n311 163.367
R466 B.n312 B.n201 163.367
R467 B.n316 B.n201 163.367
R468 B.n317 B.n316 163.367
R469 B.n318 B.n317 163.367
R470 B.n318 B.n199 163.367
R471 B.n322 B.n199 163.367
R472 B.n323 B.n322 163.367
R473 B.n324 B.n323 163.367
R474 B.n324 B.n197 163.367
R475 B.n328 B.n197 163.367
R476 B.n329 B.n328 163.367
R477 B.n330 B.n329 163.367
R478 B.n330 B.n195 163.367
R479 B.n334 B.n195 163.367
R480 B.n335 B.n334 163.367
R481 B.n336 B.n335 163.367
R482 B.n336 B.n193 163.367
R483 B.n340 B.n193 163.367
R484 B.n341 B.n340 163.367
R485 B.n342 B.n341 163.367
R486 B.n342 B.n191 163.367
R487 B.n346 B.n191 163.367
R488 B.n347 B.n346 163.367
R489 B.n348 B.n347 163.367
R490 B.n348 B.n189 163.367
R491 B.n352 B.n189 163.367
R492 B.n353 B.n352 163.367
R493 B.n354 B.n353 163.367
R494 B.n354 B.n187 163.367
R495 B.n358 B.n187 163.367
R496 B.n359 B.n358 163.367
R497 B.n360 B.n359 163.367
R498 B.n360 B.n185 163.367
R499 B.n364 B.n185 163.367
R500 B.n365 B.n364 163.367
R501 B.n366 B.n365 163.367
R502 B.n366 B.n183 163.367
R503 B.n370 B.n183 163.367
R504 B.n371 B.n370 163.367
R505 B.n372 B.n371 163.367
R506 B.n372 B.n181 163.367
R507 B.n376 B.n181 163.367
R508 B.n377 B.n376 163.367
R509 B.n378 B.n377 163.367
R510 B.n378 B.n179 163.367
R511 B.n382 B.n179 163.367
R512 B.n383 B.n382 163.367
R513 B.n384 B.n383 163.367
R514 B.n384 B.n175 163.367
R515 B.n389 B.n175 163.367
R516 B.n390 B.n389 163.367
R517 B.n391 B.n390 163.367
R518 B.n391 B.n173 163.367
R519 B.n395 B.n173 163.367
R520 B.n396 B.n395 163.367
R521 B.n397 B.n396 163.367
R522 B.n397 B.n171 163.367
R523 B.n404 B.n171 163.367
R524 B.n405 B.n404 163.367
R525 B.n406 B.n405 163.367
R526 B.n406 B.n169 163.367
R527 B.n410 B.n169 163.367
R528 B.n411 B.n410 163.367
R529 B.n412 B.n411 163.367
R530 B.n412 B.n167 163.367
R531 B.n416 B.n167 163.367
R532 B.n417 B.n416 163.367
R533 B.n418 B.n417 163.367
R534 B.n418 B.n165 163.367
R535 B.n422 B.n165 163.367
R536 B.n423 B.n422 163.367
R537 B.n424 B.n423 163.367
R538 B.n424 B.n163 163.367
R539 B.n428 B.n163 163.367
R540 B.n429 B.n428 163.367
R541 B.n430 B.n429 163.367
R542 B.n430 B.n161 163.367
R543 B.n434 B.n161 163.367
R544 B.n435 B.n434 163.367
R545 B.n436 B.n435 163.367
R546 B.n436 B.n159 163.367
R547 B.n440 B.n159 163.367
R548 B.n441 B.n440 163.367
R549 B.n442 B.n441 163.367
R550 B.n442 B.n157 163.367
R551 B.n446 B.n157 163.367
R552 B.n447 B.n446 163.367
R553 B.n448 B.n447 163.367
R554 B.n448 B.n155 163.367
R555 B.n452 B.n155 163.367
R556 B.n453 B.n452 163.367
R557 B.n454 B.n453 163.367
R558 B.n454 B.n153 163.367
R559 B.n458 B.n153 163.367
R560 B.n459 B.n458 163.367
R561 B.n460 B.n459 163.367
R562 B.n460 B.n151 163.367
R563 B.n464 B.n151 163.367
R564 B.n465 B.n464 163.367
R565 B.n466 B.n465 163.367
R566 B.n466 B.n149 163.367
R567 B.n470 B.n149 163.367
R568 B.n471 B.n470 163.367
R569 B.n472 B.n471 163.367
R570 B.n472 B.n147 163.367
R571 B.n476 B.n147 163.367
R572 B.n477 B.n476 163.367
R573 B.n478 B.n477 163.367
R574 B.n478 B.n145 163.367
R575 B.n482 B.n145 163.367
R576 B.n483 B.n482 163.367
R577 B.n484 B.n483 163.367
R578 B.n484 B.n143 163.367
R579 B.n488 B.n143 163.367
R580 B.n489 B.n488 163.367
R581 B.n490 B.n489 163.367
R582 B.n490 B.n141 163.367
R583 B.n494 B.n141 163.367
R584 B.n495 B.n494 163.367
R585 B.n633 B.n632 163.367
R586 B.n632 B.n95 163.367
R587 B.n628 B.n95 163.367
R588 B.n628 B.n627 163.367
R589 B.n627 B.n626 163.367
R590 B.n626 B.n97 163.367
R591 B.n622 B.n97 163.367
R592 B.n622 B.n621 163.367
R593 B.n621 B.n620 163.367
R594 B.n620 B.n99 163.367
R595 B.n616 B.n99 163.367
R596 B.n616 B.n615 163.367
R597 B.n615 B.n614 163.367
R598 B.n614 B.n101 163.367
R599 B.n610 B.n101 163.367
R600 B.n610 B.n609 163.367
R601 B.n609 B.n608 163.367
R602 B.n608 B.n103 163.367
R603 B.n604 B.n103 163.367
R604 B.n604 B.n603 163.367
R605 B.n603 B.n602 163.367
R606 B.n602 B.n105 163.367
R607 B.n598 B.n105 163.367
R608 B.n598 B.n597 163.367
R609 B.n597 B.n596 163.367
R610 B.n596 B.n107 163.367
R611 B.n592 B.n107 163.367
R612 B.n592 B.n591 163.367
R613 B.n591 B.n590 163.367
R614 B.n590 B.n109 163.367
R615 B.n586 B.n109 163.367
R616 B.n586 B.n585 163.367
R617 B.n585 B.n584 163.367
R618 B.n584 B.n111 163.367
R619 B.n580 B.n111 163.367
R620 B.n580 B.n579 163.367
R621 B.n579 B.n578 163.367
R622 B.n578 B.n113 163.367
R623 B.n574 B.n113 163.367
R624 B.n574 B.n573 163.367
R625 B.n573 B.n572 163.367
R626 B.n572 B.n115 163.367
R627 B.n568 B.n115 163.367
R628 B.n568 B.n567 163.367
R629 B.n567 B.n566 163.367
R630 B.n566 B.n117 163.367
R631 B.n562 B.n117 163.367
R632 B.n562 B.n561 163.367
R633 B.n561 B.n560 163.367
R634 B.n560 B.n119 163.367
R635 B.n556 B.n119 163.367
R636 B.n556 B.n555 163.367
R637 B.n555 B.n554 163.367
R638 B.n554 B.n121 163.367
R639 B.n550 B.n121 163.367
R640 B.n550 B.n549 163.367
R641 B.n549 B.n548 163.367
R642 B.n548 B.n123 163.367
R643 B.n544 B.n123 163.367
R644 B.n544 B.n543 163.367
R645 B.n543 B.n542 163.367
R646 B.n542 B.n125 163.367
R647 B.n538 B.n125 163.367
R648 B.n538 B.n537 163.367
R649 B.n537 B.n536 163.367
R650 B.n536 B.n127 163.367
R651 B.n532 B.n127 163.367
R652 B.n532 B.n531 163.367
R653 B.n531 B.n530 163.367
R654 B.n530 B.n129 163.367
R655 B.n526 B.n129 163.367
R656 B.n526 B.n525 163.367
R657 B.n525 B.n524 163.367
R658 B.n524 B.n131 163.367
R659 B.n520 B.n131 163.367
R660 B.n520 B.n519 163.367
R661 B.n519 B.n518 163.367
R662 B.n518 B.n133 163.367
R663 B.n514 B.n133 163.367
R664 B.n514 B.n513 163.367
R665 B.n513 B.n512 163.367
R666 B.n512 B.n135 163.367
R667 B.n508 B.n135 163.367
R668 B.n508 B.n507 163.367
R669 B.n507 B.n506 163.367
R670 B.n506 B.n137 163.367
R671 B.n502 B.n137 163.367
R672 B.n502 B.n501 163.367
R673 B.n501 B.n500 163.367
R674 B.n500 B.n139 163.367
R675 B.n496 B.n139 163.367
R676 B.n832 B.n25 163.367
R677 B.n828 B.n25 163.367
R678 B.n828 B.n827 163.367
R679 B.n827 B.n826 163.367
R680 B.n826 B.n27 163.367
R681 B.n822 B.n27 163.367
R682 B.n822 B.n821 163.367
R683 B.n821 B.n820 163.367
R684 B.n820 B.n29 163.367
R685 B.n816 B.n29 163.367
R686 B.n816 B.n815 163.367
R687 B.n815 B.n814 163.367
R688 B.n814 B.n31 163.367
R689 B.n810 B.n31 163.367
R690 B.n810 B.n809 163.367
R691 B.n809 B.n808 163.367
R692 B.n808 B.n33 163.367
R693 B.n804 B.n33 163.367
R694 B.n804 B.n803 163.367
R695 B.n803 B.n802 163.367
R696 B.n802 B.n35 163.367
R697 B.n798 B.n35 163.367
R698 B.n798 B.n797 163.367
R699 B.n797 B.n796 163.367
R700 B.n796 B.n37 163.367
R701 B.n792 B.n37 163.367
R702 B.n792 B.n791 163.367
R703 B.n791 B.n790 163.367
R704 B.n790 B.n39 163.367
R705 B.n786 B.n39 163.367
R706 B.n786 B.n785 163.367
R707 B.n785 B.n784 163.367
R708 B.n784 B.n41 163.367
R709 B.n780 B.n41 163.367
R710 B.n780 B.n779 163.367
R711 B.n779 B.n778 163.367
R712 B.n778 B.n43 163.367
R713 B.n774 B.n43 163.367
R714 B.n774 B.n773 163.367
R715 B.n773 B.n772 163.367
R716 B.n772 B.n45 163.367
R717 B.n768 B.n45 163.367
R718 B.n768 B.n767 163.367
R719 B.n767 B.n766 163.367
R720 B.n766 B.n47 163.367
R721 B.n762 B.n47 163.367
R722 B.n762 B.n761 163.367
R723 B.n761 B.n760 163.367
R724 B.n760 B.n49 163.367
R725 B.n756 B.n49 163.367
R726 B.n756 B.n755 163.367
R727 B.n755 B.n754 163.367
R728 B.n754 B.n51 163.367
R729 B.n750 B.n51 163.367
R730 B.n750 B.n749 163.367
R731 B.n749 B.n748 163.367
R732 B.n748 B.n53 163.367
R733 B.n744 B.n53 163.367
R734 B.n744 B.n743 163.367
R735 B.n743 B.n742 163.367
R736 B.n742 B.n55 163.367
R737 B.n737 B.n55 163.367
R738 B.n737 B.n736 163.367
R739 B.n736 B.n735 163.367
R740 B.n735 B.n59 163.367
R741 B.n731 B.n59 163.367
R742 B.n731 B.n730 163.367
R743 B.n730 B.n729 163.367
R744 B.n729 B.n61 163.367
R745 B.n724 B.n61 163.367
R746 B.n724 B.n723 163.367
R747 B.n723 B.n722 163.367
R748 B.n722 B.n65 163.367
R749 B.n718 B.n65 163.367
R750 B.n718 B.n717 163.367
R751 B.n717 B.n716 163.367
R752 B.n716 B.n67 163.367
R753 B.n712 B.n67 163.367
R754 B.n712 B.n711 163.367
R755 B.n711 B.n710 163.367
R756 B.n710 B.n69 163.367
R757 B.n706 B.n69 163.367
R758 B.n706 B.n705 163.367
R759 B.n705 B.n704 163.367
R760 B.n704 B.n71 163.367
R761 B.n700 B.n71 163.367
R762 B.n700 B.n699 163.367
R763 B.n699 B.n698 163.367
R764 B.n698 B.n73 163.367
R765 B.n694 B.n73 163.367
R766 B.n694 B.n693 163.367
R767 B.n693 B.n692 163.367
R768 B.n692 B.n75 163.367
R769 B.n688 B.n75 163.367
R770 B.n688 B.n687 163.367
R771 B.n687 B.n686 163.367
R772 B.n686 B.n77 163.367
R773 B.n682 B.n77 163.367
R774 B.n682 B.n681 163.367
R775 B.n681 B.n680 163.367
R776 B.n680 B.n79 163.367
R777 B.n676 B.n79 163.367
R778 B.n676 B.n675 163.367
R779 B.n675 B.n674 163.367
R780 B.n674 B.n81 163.367
R781 B.n670 B.n81 163.367
R782 B.n670 B.n669 163.367
R783 B.n669 B.n668 163.367
R784 B.n668 B.n83 163.367
R785 B.n664 B.n83 163.367
R786 B.n664 B.n663 163.367
R787 B.n663 B.n662 163.367
R788 B.n662 B.n85 163.367
R789 B.n658 B.n85 163.367
R790 B.n658 B.n657 163.367
R791 B.n657 B.n656 163.367
R792 B.n656 B.n87 163.367
R793 B.n652 B.n87 163.367
R794 B.n652 B.n651 163.367
R795 B.n651 B.n650 163.367
R796 B.n650 B.n89 163.367
R797 B.n646 B.n89 163.367
R798 B.n646 B.n645 163.367
R799 B.n645 B.n644 163.367
R800 B.n644 B.n91 163.367
R801 B.n640 B.n91 163.367
R802 B.n640 B.n639 163.367
R803 B.n639 B.n638 163.367
R804 B.n638 B.n93 163.367
R805 B.n634 B.n93 163.367
R806 B.n834 B.n833 163.367
R807 B.n834 B.n23 163.367
R808 B.n838 B.n23 163.367
R809 B.n839 B.n838 163.367
R810 B.n840 B.n839 163.367
R811 B.n840 B.n21 163.367
R812 B.n844 B.n21 163.367
R813 B.n845 B.n844 163.367
R814 B.n846 B.n845 163.367
R815 B.n846 B.n19 163.367
R816 B.n850 B.n19 163.367
R817 B.n851 B.n850 163.367
R818 B.n852 B.n851 163.367
R819 B.n852 B.n17 163.367
R820 B.n856 B.n17 163.367
R821 B.n857 B.n856 163.367
R822 B.n858 B.n857 163.367
R823 B.n858 B.n15 163.367
R824 B.n862 B.n15 163.367
R825 B.n863 B.n862 163.367
R826 B.n864 B.n863 163.367
R827 B.n864 B.n13 163.367
R828 B.n868 B.n13 163.367
R829 B.n869 B.n868 163.367
R830 B.n870 B.n869 163.367
R831 B.n870 B.n11 163.367
R832 B.n874 B.n11 163.367
R833 B.n875 B.n874 163.367
R834 B.n876 B.n875 163.367
R835 B.n876 B.n9 163.367
R836 B.n880 B.n9 163.367
R837 B.n881 B.n880 163.367
R838 B.n882 B.n881 163.367
R839 B.n882 B.n7 163.367
R840 B.n886 B.n7 163.367
R841 B.n887 B.n886 163.367
R842 B.n888 B.n887 163.367
R843 B.n888 B.n5 163.367
R844 B.n892 B.n5 163.367
R845 B.n893 B.n892 163.367
R846 B.n894 B.n893 163.367
R847 B.n894 B.n3 163.367
R848 B.n898 B.n3 163.367
R849 B.n899 B.n898 163.367
R850 B.n229 B.n2 163.367
R851 B.n232 B.n229 163.367
R852 B.n233 B.n232 163.367
R853 B.n234 B.n233 163.367
R854 B.n234 B.n227 163.367
R855 B.n238 B.n227 163.367
R856 B.n239 B.n238 163.367
R857 B.n240 B.n239 163.367
R858 B.n240 B.n225 163.367
R859 B.n244 B.n225 163.367
R860 B.n245 B.n244 163.367
R861 B.n246 B.n245 163.367
R862 B.n246 B.n223 163.367
R863 B.n250 B.n223 163.367
R864 B.n251 B.n250 163.367
R865 B.n252 B.n251 163.367
R866 B.n252 B.n221 163.367
R867 B.n256 B.n221 163.367
R868 B.n257 B.n256 163.367
R869 B.n258 B.n257 163.367
R870 B.n258 B.n219 163.367
R871 B.n262 B.n219 163.367
R872 B.n263 B.n262 163.367
R873 B.n264 B.n263 163.367
R874 B.n264 B.n217 163.367
R875 B.n268 B.n217 163.367
R876 B.n269 B.n268 163.367
R877 B.n270 B.n269 163.367
R878 B.n270 B.n215 163.367
R879 B.n274 B.n215 163.367
R880 B.n275 B.n274 163.367
R881 B.n276 B.n275 163.367
R882 B.n276 B.n213 163.367
R883 B.n280 B.n213 163.367
R884 B.n281 B.n280 163.367
R885 B.n282 B.n281 163.367
R886 B.n282 B.n211 163.367
R887 B.n286 B.n211 163.367
R888 B.n287 B.n286 163.367
R889 B.n288 B.n287 163.367
R890 B.n288 B.n209 163.367
R891 B.n292 B.n209 163.367
R892 B.n293 B.n292 163.367
R893 B.n294 B.n293 163.367
R894 B.n400 B.t4 157.362
R895 B.n62 B.t8 157.362
R896 B.n176 B.t10 157.338
R897 B.n56 B.t2 157.338
R898 B.n401 B.t5 107.713
R899 B.n63 B.t7 107.713
R900 B.n177 B.t11 107.689
R901 B.n57 B.t1 107.689
R902 B.n387 B.n177 59.5399
R903 B.n402 B.n401 59.5399
R904 B.n726 B.n63 59.5399
R905 B.n740 B.n57 59.5399
R906 B.n177 B.n176 49.649
R907 B.n401 B.n400 49.649
R908 B.n63 B.n62 49.649
R909 B.n57 B.n56 49.649
R910 B.n831 B.n24 33.5615
R911 B.n635 B.n94 33.5615
R912 B.n497 B.n140 33.5615
R913 B.n296 B.n295 33.5615
R914 B B.n901 18.0485
R915 B.n835 B.n24 10.6151
R916 B.n836 B.n835 10.6151
R917 B.n837 B.n836 10.6151
R918 B.n837 B.n22 10.6151
R919 B.n841 B.n22 10.6151
R920 B.n842 B.n841 10.6151
R921 B.n843 B.n842 10.6151
R922 B.n843 B.n20 10.6151
R923 B.n847 B.n20 10.6151
R924 B.n848 B.n847 10.6151
R925 B.n849 B.n848 10.6151
R926 B.n849 B.n18 10.6151
R927 B.n853 B.n18 10.6151
R928 B.n854 B.n853 10.6151
R929 B.n855 B.n854 10.6151
R930 B.n855 B.n16 10.6151
R931 B.n859 B.n16 10.6151
R932 B.n860 B.n859 10.6151
R933 B.n861 B.n860 10.6151
R934 B.n861 B.n14 10.6151
R935 B.n865 B.n14 10.6151
R936 B.n866 B.n865 10.6151
R937 B.n867 B.n866 10.6151
R938 B.n867 B.n12 10.6151
R939 B.n871 B.n12 10.6151
R940 B.n872 B.n871 10.6151
R941 B.n873 B.n872 10.6151
R942 B.n873 B.n10 10.6151
R943 B.n877 B.n10 10.6151
R944 B.n878 B.n877 10.6151
R945 B.n879 B.n878 10.6151
R946 B.n879 B.n8 10.6151
R947 B.n883 B.n8 10.6151
R948 B.n884 B.n883 10.6151
R949 B.n885 B.n884 10.6151
R950 B.n885 B.n6 10.6151
R951 B.n889 B.n6 10.6151
R952 B.n890 B.n889 10.6151
R953 B.n891 B.n890 10.6151
R954 B.n891 B.n4 10.6151
R955 B.n895 B.n4 10.6151
R956 B.n896 B.n895 10.6151
R957 B.n897 B.n896 10.6151
R958 B.n897 B.n0 10.6151
R959 B.n831 B.n830 10.6151
R960 B.n830 B.n829 10.6151
R961 B.n829 B.n26 10.6151
R962 B.n825 B.n26 10.6151
R963 B.n825 B.n824 10.6151
R964 B.n824 B.n823 10.6151
R965 B.n823 B.n28 10.6151
R966 B.n819 B.n28 10.6151
R967 B.n819 B.n818 10.6151
R968 B.n818 B.n817 10.6151
R969 B.n817 B.n30 10.6151
R970 B.n813 B.n30 10.6151
R971 B.n813 B.n812 10.6151
R972 B.n812 B.n811 10.6151
R973 B.n811 B.n32 10.6151
R974 B.n807 B.n32 10.6151
R975 B.n807 B.n806 10.6151
R976 B.n806 B.n805 10.6151
R977 B.n805 B.n34 10.6151
R978 B.n801 B.n34 10.6151
R979 B.n801 B.n800 10.6151
R980 B.n800 B.n799 10.6151
R981 B.n799 B.n36 10.6151
R982 B.n795 B.n36 10.6151
R983 B.n795 B.n794 10.6151
R984 B.n794 B.n793 10.6151
R985 B.n793 B.n38 10.6151
R986 B.n789 B.n38 10.6151
R987 B.n789 B.n788 10.6151
R988 B.n788 B.n787 10.6151
R989 B.n787 B.n40 10.6151
R990 B.n783 B.n40 10.6151
R991 B.n783 B.n782 10.6151
R992 B.n782 B.n781 10.6151
R993 B.n781 B.n42 10.6151
R994 B.n777 B.n42 10.6151
R995 B.n777 B.n776 10.6151
R996 B.n776 B.n775 10.6151
R997 B.n775 B.n44 10.6151
R998 B.n771 B.n44 10.6151
R999 B.n771 B.n770 10.6151
R1000 B.n770 B.n769 10.6151
R1001 B.n769 B.n46 10.6151
R1002 B.n765 B.n46 10.6151
R1003 B.n765 B.n764 10.6151
R1004 B.n764 B.n763 10.6151
R1005 B.n763 B.n48 10.6151
R1006 B.n759 B.n48 10.6151
R1007 B.n759 B.n758 10.6151
R1008 B.n758 B.n757 10.6151
R1009 B.n757 B.n50 10.6151
R1010 B.n753 B.n50 10.6151
R1011 B.n753 B.n752 10.6151
R1012 B.n752 B.n751 10.6151
R1013 B.n751 B.n52 10.6151
R1014 B.n747 B.n52 10.6151
R1015 B.n747 B.n746 10.6151
R1016 B.n746 B.n745 10.6151
R1017 B.n745 B.n54 10.6151
R1018 B.n741 B.n54 10.6151
R1019 B.n739 B.n738 10.6151
R1020 B.n738 B.n58 10.6151
R1021 B.n734 B.n58 10.6151
R1022 B.n734 B.n733 10.6151
R1023 B.n733 B.n732 10.6151
R1024 B.n732 B.n60 10.6151
R1025 B.n728 B.n60 10.6151
R1026 B.n728 B.n727 10.6151
R1027 B.n725 B.n64 10.6151
R1028 B.n721 B.n64 10.6151
R1029 B.n721 B.n720 10.6151
R1030 B.n720 B.n719 10.6151
R1031 B.n719 B.n66 10.6151
R1032 B.n715 B.n66 10.6151
R1033 B.n715 B.n714 10.6151
R1034 B.n714 B.n713 10.6151
R1035 B.n713 B.n68 10.6151
R1036 B.n709 B.n68 10.6151
R1037 B.n709 B.n708 10.6151
R1038 B.n708 B.n707 10.6151
R1039 B.n707 B.n70 10.6151
R1040 B.n703 B.n70 10.6151
R1041 B.n703 B.n702 10.6151
R1042 B.n702 B.n701 10.6151
R1043 B.n701 B.n72 10.6151
R1044 B.n697 B.n72 10.6151
R1045 B.n697 B.n696 10.6151
R1046 B.n696 B.n695 10.6151
R1047 B.n695 B.n74 10.6151
R1048 B.n691 B.n74 10.6151
R1049 B.n691 B.n690 10.6151
R1050 B.n690 B.n689 10.6151
R1051 B.n689 B.n76 10.6151
R1052 B.n685 B.n76 10.6151
R1053 B.n685 B.n684 10.6151
R1054 B.n684 B.n683 10.6151
R1055 B.n683 B.n78 10.6151
R1056 B.n679 B.n78 10.6151
R1057 B.n679 B.n678 10.6151
R1058 B.n678 B.n677 10.6151
R1059 B.n677 B.n80 10.6151
R1060 B.n673 B.n80 10.6151
R1061 B.n673 B.n672 10.6151
R1062 B.n672 B.n671 10.6151
R1063 B.n671 B.n82 10.6151
R1064 B.n667 B.n82 10.6151
R1065 B.n667 B.n666 10.6151
R1066 B.n666 B.n665 10.6151
R1067 B.n665 B.n84 10.6151
R1068 B.n661 B.n84 10.6151
R1069 B.n661 B.n660 10.6151
R1070 B.n660 B.n659 10.6151
R1071 B.n659 B.n86 10.6151
R1072 B.n655 B.n86 10.6151
R1073 B.n655 B.n654 10.6151
R1074 B.n654 B.n653 10.6151
R1075 B.n653 B.n88 10.6151
R1076 B.n649 B.n88 10.6151
R1077 B.n649 B.n648 10.6151
R1078 B.n648 B.n647 10.6151
R1079 B.n647 B.n90 10.6151
R1080 B.n643 B.n90 10.6151
R1081 B.n643 B.n642 10.6151
R1082 B.n642 B.n641 10.6151
R1083 B.n641 B.n92 10.6151
R1084 B.n637 B.n92 10.6151
R1085 B.n637 B.n636 10.6151
R1086 B.n636 B.n635 10.6151
R1087 B.n631 B.n94 10.6151
R1088 B.n631 B.n630 10.6151
R1089 B.n630 B.n629 10.6151
R1090 B.n629 B.n96 10.6151
R1091 B.n625 B.n96 10.6151
R1092 B.n625 B.n624 10.6151
R1093 B.n624 B.n623 10.6151
R1094 B.n623 B.n98 10.6151
R1095 B.n619 B.n98 10.6151
R1096 B.n619 B.n618 10.6151
R1097 B.n618 B.n617 10.6151
R1098 B.n617 B.n100 10.6151
R1099 B.n613 B.n100 10.6151
R1100 B.n613 B.n612 10.6151
R1101 B.n612 B.n611 10.6151
R1102 B.n611 B.n102 10.6151
R1103 B.n607 B.n102 10.6151
R1104 B.n607 B.n606 10.6151
R1105 B.n606 B.n605 10.6151
R1106 B.n605 B.n104 10.6151
R1107 B.n601 B.n104 10.6151
R1108 B.n601 B.n600 10.6151
R1109 B.n600 B.n599 10.6151
R1110 B.n599 B.n106 10.6151
R1111 B.n595 B.n106 10.6151
R1112 B.n595 B.n594 10.6151
R1113 B.n594 B.n593 10.6151
R1114 B.n593 B.n108 10.6151
R1115 B.n589 B.n108 10.6151
R1116 B.n589 B.n588 10.6151
R1117 B.n588 B.n587 10.6151
R1118 B.n587 B.n110 10.6151
R1119 B.n583 B.n110 10.6151
R1120 B.n583 B.n582 10.6151
R1121 B.n582 B.n581 10.6151
R1122 B.n581 B.n112 10.6151
R1123 B.n577 B.n112 10.6151
R1124 B.n577 B.n576 10.6151
R1125 B.n576 B.n575 10.6151
R1126 B.n575 B.n114 10.6151
R1127 B.n571 B.n114 10.6151
R1128 B.n571 B.n570 10.6151
R1129 B.n570 B.n569 10.6151
R1130 B.n569 B.n116 10.6151
R1131 B.n565 B.n116 10.6151
R1132 B.n565 B.n564 10.6151
R1133 B.n564 B.n563 10.6151
R1134 B.n563 B.n118 10.6151
R1135 B.n559 B.n118 10.6151
R1136 B.n559 B.n558 10.6151
R1137 B.n558 B.n557 10.6151
R1138 B.n557 B.n120 10.6151
R1139 B.n553 B.n120 10.6151
R1140 B.n553 B.n552 10.6151
R1141 B.n552 B.n551 10.6151
R1142 B.n551 B.n122 10.6151
R1143 B.n547 B.n122 10.6151
R1144 B.n547 B.n546 10.6151
R1145 B.n546 B.n545 10.6151
R1146 B.n545 B.n124 10.6151
R1147 B.n541 B.n124 10.6151
R1148 B.n541 B.n540 10.6151
R1149 B.n540 B.n539 10.6151
R1150 B.n539 B.n126 10.6151
R1151 B.n535 B.n126 10.6151
R1152 B.n535 B.n534 10.6151
R1153 B.n534 B.n533 10.6151
R1154 B.n533 B.n128 10.6151
R1155 B.n529 B.n128 10.6151
R1156 B.n529 B.n528 10.6151
R1157 B.n528 B.n527 10.6151
R1158 B.n527 B.n130 10.6151
R1159 B.n523 B.n130 10.6151
R1160 B.n523 B.n522 10.6151
R1161 B.n522 B.n521 10.6151
R1162 B.n521 B.n132 10.6151
R1163 B.n517 B.n132 10.6151
R1164 B.n517 B.n516 10.6151
R1165 B.n516 B.n515 10.6151
R1166 B.n515 B.n134 10.6151
R1167 B.n511 B.n134 10.6151
R1168 B.n511 B.n510 10.6151
R1169 B.n510 B.n509 10.6151
R1170 B.n509 B.n136 10.6151
R1171 B.n505 B.n136 10.6151
R1172 B.n505 B.n504 10.6151
R1173 B.n504 B.n503 10.6151
R1174 B.n503 B.n138 10.6151
R1175 B.n499 B.n138 10.6151
R1176 B.n499 B.n498 10.6151
R1177 B.n498 B.n497 10.6151
R1178 B.n230 B.n1 10.6151
R1179 B.n231 B.n230 10.6151
R1180 B.n231 B.n228 10.6151
R1181 B.n235 B.n228 10.6151
R1182 B.n236 B.n235 10.6151
R1183 B.n237 B.n236 10.6151
R1184 B.n237 B.n226 10.6151
R1185 B.n241 B.n226 10.6151
R1186 B.n242 B.n241 10.6151
R1187 B.n243 B.n242 10.6151
R1188 B.n243 B.n224 10.6151
R1189 B.n247 B.n224 10.6151
R1190 B.n248 B.n247 10.6151
R1191 B.n249 B.n248 10.6151
R1192 B.n249 B.n222 10.6151
R1193 B.n253 B.n222 10.6151
R1194 B.n254 B.n253 10.6151
R1195 B.n255 B.n254 10.6151
R1196 B.n255 B.n220 10.6151
R1197 B.n259 B.n220 10.6151
R1198 B.n260 B.n259 10.6151
R1199 B.n261 B.n260 10.6151
R1200 B.n261 B.n218 10.6151
R1201 B.n265 B.n218 10.6151
R1202 B.n266 B.n265 10.6151
R1203 B.n267 B.n266 10.6151
R1204 B.n267 B.n216 10.6151
R1205 B.n271 B.n216 10.6151
R1206 B.n272 B.n271 10.6151
R1207 B.n273 B.n272 10.6151
R1208 B.n273 B.n214 10.6151
R1209 B.n277 B.n214 10.6151
R1210 B.n278 B.n277 10.6151
R1211 B.n279 B.n278 10.6151
R1212 B.n279 B.n212 10.6151
R1213 B.n283 B.n212 10.6151
R1214 B.n284 B.n283 10.6151
R1215 B.n285 B.n284 10.6151
R1216 B.n285 B.n210 10.6151
R1217 B.n289 B.n210 10.6151
R1218 B.n290 B.n289 10.6151
R1219 B.n291 B.n290 10.6151
R1220 B.n291 B.n208 10.6151
R1221 B.n295 B.n208 10.6151
R1222 B.n297 B.n296 10.6151
R1223 B.n297 B.n206 10.6151
R1224 B.n301 B.n206 10.6151
R1225 B.n302 B.n301 10.6151
R1226 B.n303 B.n302 10.6151
R1227 B.n303 B.n204 10.6151
R1228 B.n307 B.n204 10.6151
R1229 B.n308 B.n307 10.6151
R1230 B.n309 B.n308 10.6151
R1231 B.n309 B.n202 10.6151
R1232 B.n313 B.n202 10.6151
R1233 B.n314 B.n313 10.6151
R1234 B.n315 B.n314 10.6151
R1235 B.n315 B.n200 10.6151
R1236 B.n319 B.n200 10.6151
R1237 B.n320 B.n319 10.6151
R1238 B.n321 B.n320 10.6151
R1239 B.n321 B.n198 10.6151
R1240 B.n325 B.n198 10.6151
R1241 B.n326 B.n325 10.6151
R1242 B.n327 B.n326 10.6151
R1243 B.n327 B.n196 10.6151
R1244 B.n331 B.n196 10.6151
R1245 B.n332 B.n331 10.6151
R1246 B.n333 B.n332 10.6151
R1247 B.n333 B.n194 10.6151
R1248 B.n337 B.n194 10.6151
R1249 B.n338 B.n337 10.6151
R1250 B.n339 B.n338 10.6151
R1251 B.n339 B.n192 10.6151
R1252 B.n343 B.n192 10.6151
R1253 B.n344 B.n343 10.6151
R1254 B.n345 B.n344 10.6151
R1255 B.n345 B.n190 10.6151
R1256 B.n349 B.n190 10.6151
R1257 B.n350 B.n349 10.6151
R1258 B.n351 B.n350 10.6151
R1259 B.n351 B.n188 10.6151
R1260 B.n355 B.n188 10.6151
R1261 B.n356 B.n355 10.6151
R1262 B.n357 B.n356 10.6151
R1263 B.n357 B.n186 10.6151
R1264 B.n361 B.n186 10.6151
R1265 B.n362 B.n361 10.6151
R1266 B.n363 B.n362 10.6151
R1267 B.n363 B.n184 10.6151
R1268 B.n367 B.n184 10.6151
R1269 B.n368 B.n367 10.6151
R1270 B.n369 B.n368 10.6151
R1271 B.n369 B.n182 10.6151
R1272 B.n373 B.n182 10.6151
R1273 B.n374 B.n373 10.6151
R1274 B.n375 B.n374 10.6151
R1275 B.n375 B.n180 10.6151
R1276 B.n379 B.n180 10.6151
R1277 B.n380 B.n379 10.6151
R1278 B.n381 B.n380 10.6151
R1279 B.n381 B.n178 10.6151
R1280 B.n385 B.n178 10.6151
R1281 B.n386 B.n385 10.6151
R1282 B.n388 B.n174 10.6151
R1283 B.n392 B.n174 10.6151
R1284 B.n393 B.n392 10.6151
R1285 B.n394 B.n393 10.6151
R1286 B.n394 B.n172 10.6151
R1287 B.n398 B.n172 10.6151
R1288 B.n399 B.n398 10.6151
R1289 B.n403 B.n399 10.6151
R1290 B.n407 B.n170 10.6151
R1291 B.n408 B.n407 10.6151
R1292 B.n409 B.n408 10.6151
R1293 B.n409 B.n168 10.6151
R1294 B.n413 B.n168 10.6151
R1295 B.n414 B.n413 10.6151
R1296 B.n415 B.n414 10.6151
R1297 B.n415 B.n166 10.6151
R1298 B.n419 B.n166 10.6151
R1299 B.n420 B.n419 10.6151
R1300 B.n421 B.n420 10.6151
R1301 B.n421 B.n164 10.6151
R1302 B.n425 B.n164 10.6151
R1303 B.n426 B.n425 10.6151
R1304 B.n427 B.n426 10.6151
R1305 B.n427 B.n162 10.6151
R1306 B.n431 B.n162 10.6151
R1307 B.n432 B.n431 10.6151
R1308 B.n433 B.n432 10.6151
R1309 B.n433 B.n160 10.6151
R1310 B.n437 B.n160 10.6151
R1311 B.n438 B.n437 10.6151
R1312 B.n439 B.n438 10.6151
R1313 B.n439 B.n158 10.6151
R1314 B.n443 B.n158 10.6151
R1315 B.n444 B.n443 10.6151
R1316 B.n445 B.n444 10.6151
R1317 B.n445 B.n156 10.6151
R1318 B.n449 B.n156 10.6151
R1319 B.n450 B.n449 10.6151
R1320 B.n451 B.n450 10.6151
R1321 B.n451 B.n154 10.6151
R1322 B.n455 B.n154 10.6151
R1323 B.n456 B.n455 10.6151
R1324 B.n457 B.n456 10.6151
R1325 B.n457 B.n152 10.6151
R1326 B.n461 B.n152 10.6151
R1327 B.n462 B.n461 10.6151
R1328 B.n463 B.n462 10.6151
R1329 B.n463 B.n150 10.6151
R1330 B.n467 B.n150 10.6151
R1331 B.n468 B.n467 10.6151
R1332 B.n469 B.n468 10.6151
R1333 B.n469 B.n148 10.6151
R1334 B.n473 B.n148 10.6151
R1335 B.n474 B.n473 10.6151
R1336 B.n475 B.n474 10.6151
R1337 B.n475 B.n146 10.6151
R1338 B.n479 B.n146 10.6151
R1339 B.n480 B.n479 10.6151
R1340 B.n481 B.n480 10.6151
R1341 B.n481 B.n144 10.6151
R1342 B.n485 B.n144 10.6151
R1343 B.n486 B.n485 10.6151
R1344 B.n487 B.n486 10.6151
R1345 B.n487 B.n142 10.6151
R1346 B.n491 B.n142 10.6151
R1347 B.n492 B.n491 10.6151
R1348 B.n493 B.n492 10.6151
R1349 B.n493 B.n140 10.6151
R1350 B.n901 B.n0 8.11757
R1351 B.n901 B.n1 8.11757
R1352 B.n740 B.n739 6.5566
R1353 B.n727 B.n726 6.5566
R1354 B.n388 B.n387 6.5566
R1355 B.n403 B.n402 6.5566
R1356 B.n741 B.n740 4.05904
R1357 B.n726 B.n725 4.05904
R1358 B.n387 B.n386 4.05904
R1359 B.n402 B.n170 4.05904
R1360 VN.n6 VN.t5 232.452
R1361 VN.n31 VN.t4 232.452
R1362 VN.n5 VN.t2 199.285
R1363 VN.n15 VN.t0 199.285
R1364 VN.n23 VN.t6 199.285
R1365 VN.n30 VN.t1 199.285
R1366 VN.n40 VN.t7 199.285
R1367 VN.n48 VN.t3 199.285
R1368 VN.n47 VN.n25 161.3
R1369 VN.n46 VN.n45 161.3
R1370 VN.n44 VN.n26 161.3
R1371 VN.n43 VN.n42 161.3
R1372 VN.n41 VN.n27 161.3
R1373 VN.n39 VN.n38 161.3
R1374 VN.n37 VN.n28 161.3
R1375 VN.n36 VN.n35 161.3
R1376 VN.n34 VN.n29 161.3
R1377 VN.n33 VN.n32 161.3
R1378 VN.n22 VN.n0 161.3
R1379 VN.n21 VN.n20 161.3
R1380 VN.n19 VN.n1 161.3
R1381 VN.n18 VN.n17 161.3
R1382 VN.n16 VN.n2 161.3
R1383 VN.n14 VN.n13 161.3
R1384 VN.n12 VN.n3 161.3
R1385 VN.n11 VN.n10 161.3
R1386 VN.n9 VN.n4 161.3
R1387 VN.n8 VN.n7 161.3
R1388 VN.n24 VN.n23 94.0526
R1389 VN.n49 VN.n48 94.0526
R1390 VN.n6 VN.n5 57.4839
R1391 VN.n31 VN.n30 57.4839
R1392 VN VN.n49 54.3542
R1393 VN.n21 VN.n1 46.253
R1394 VN.n46 VN.n26 46.253
R1395 VN.n10 VN.n9 40.4106
R1396 VN.n10 VN.n3 40.4106
R1397 VN.n35 VN.n34 40.4106
R1398 VN.n35 VN.n28 40.4106
R1399 VN.n17 VN.n1 34.5682
R1400 VN.n42 VN.n26 34.5682
R1401 VN.n9 VN.n8 24.3439
R1402 VN.n14 VN.n3 24.3439
R1403 VN.n17 VN.n16 24.3439
R1404 VN.n22 VN.n21 24.3439
R1405 VN.n34 VN.n33 24.3439
R1406 VN.n42 VN.n41 24.3439
R1407 VN.n39 VN.n28 24.3439
R1408 VN.n47 VN.n46 24.3439
R1409 VN.n23 VN.n22 16.554
R1410 VN.n48 VN.n47 16.554
R1411 VN.n8 VN.n5 13.6328
R1412 VN.n15 VN.n14 13.6328
R1413 VN.n33 VN.n30 13.6328
R1414 VN.n40 VN.n39 13.6328
R1415 VN.n16 VN.n15 10.7116
R1416 VN.n41 VN.n40 10.7116
R1417 VN.n32 VN.n31 9.31384
R1418 VN.n7 VN.n6 9.31384
R1419 VN.n49 VN.n25 0.278398
R1420 VN.n24 VN.n0 0.278398
R1421 VN.n45 VN.n25 0.189894
R1422 VN.n45 VN.n44 0.189894
R1423 VN.n44 VN.n43 0.189894
R1424 VN.n43 VN.n27 0.189894
R1425 VN.n38 VN.n27 0.189894
R1426 VN.n38 VN.n37 0.189894
R1427 VN.n37 VN.n36 0.189894
R1428 VN.n36 VN.n29 0.189894
R1429 VN.n32 VN.n29 0.189894
R1430 VN.n7 VN.n4 0.189894
R1431 VN.n11 VN.n4 0.189894
R1432 VN.n12 VN.n11 0.189894
R1433 VN.n13 VN.n12 0.189894
R1434 VN.n13 VN.n2 0.189894
R1435 VN.n18 VN.n2 0.189894
R1436 VN.n19 VN.n18 0.189894
R1437 VN.n20 VN.n19 0.189894
R1438 VN.n20 VN.n0 0.189894
R1439 VN VN.n24 0.153422
R1440 VDD2.n2 VDD2.n1 73.1364
R1441 VDD2.n2 VDD2.n0 73.1364
R1442 VDD2 VDD2.n5 73.1327
R1443 VDD2.n4 VDD2.n3 72.0886
R1444 VDD2.n4 VDD2.n2 49.5429
R1445 VDD2.n5 VDD2.t1 1.76324
R1446 VDD2.n5 VDD2.t6 1.76324
R1447 VDD2.n3 VDD2.t4 1.76324
R1448 VDD2.n3 VDD2.t0 1.76324
R1449 VDD2.n1 VDD2.t7 1.76324
R1450 VDD2.n1 VDD2.t5 1.76324
R1451 VDD2.n0 VDD2.t3 1.76324
R1452 VDD2.n0 VDD2.t2 1.76324
R1453 VDD2 VDD2.n4 1.16214
R1454 VTAIL.n11 VTAIL.t6 57.1725
R1455 VTAIL.n10 VTAIL.t10 57.1725
R1456 VTAIL.n7 VTAIL.t11 57.1725
R1457 VTAIL.n15 VTAIL.t8 57.1715
R1458 VTAIL.n2 VTAIL.t9 57.1715
R1459 VTAIL.n3 VTAIL.t5 57.1715
R1460 VTAIL.n6 VTAIL.t1 57.1715
R1461 VTAIL.n14 VTAIL.t3 57.1714
R1462 VTAIL.n13 VTAIL.n12 55.4098
R1463 VTAIL.n9 VTAIL.n8 55.4098
R1464 VTAIL.n1 VTAIL.n0 55.4096
R1465 VTAIL.n5 VTAIL.n4 55.4096
R1466 VTAIL.n15 VTAIL.n14 30.4703
R1467 VTAIL.n7 VTAIL.n6 30.4703
R1468 VTAIL.n9 VTAIL.n7 2.2074
R1469 VTAIL.n10 VTAIL.n9 2.2074
R1470 VTAIL.n13 VTAIL.n11 2.2074
R1471 VTAIL.n14 VTAIL.n13 2.2074
R1472 VTAIL.n6 VTAIL.n5 2.2074
R1473 VTAIL.n5 VTAIL.n3 2.2074
R1474 VTAIL.n2 VTAIL.n1 2.2074
R1475 VTAIL VTAIL.n15 2.14921
R1476 VTAIL.n0 VTAIL.t12 1.76324
R1477 VTAIL.n0 VTAIL.t14 1.76324
R1478 VTAIL.n4 VTAIL.t4 1.76324
R1479 VTAIL.n4 VTAIL.t2 1.76324
R1480 VTAIL.n12 VTAIL.t0 1.76324
R1481 VTAIL.n12 VTAIL.t15 1.76324
R1482 VTAIL.n8 VTAIL.t7 1.76324
R1483 VTAIL.n8 VTAIL.t13 1.76324
R1484 VTAIL.n11 VTAIL.n10 0.470328
R1485 VTAIL.n3 VTAIL.n2 0.470328
R1486 VTAIL VTAIL.n1 0.0586897
R1487 VP.n14 VP.t1 232.452
R1488 VP.n34 VP.t2 199.285
R1489 VP.n5 VP.t5 199.285
R1490 VP.n51 VP.t0 199.285
R1491 VP.n59 VP.t3 199.285
R1492 VP.n31 VP.t7 199.285
R1493 VP.n23 VP.t4 199.285
R1494 VP.n13 VP.t6 199.285
R1495 VP.n16 VP.n15 161.3
R1496 VP.n17 VP.n12 161.3
R1497 VP.n19 VP.n18 161.3
R1498 VP.n20 VP.n11 161.3
R1499 VP.n22 VP.n21 161.3
R1500 VP.n24 VP.n10 161.3
R1501 VP.n26 VP.n25 161.3
R1502 VP.n27 VP.n9 161.3
R1503 VP.n29 VP.n28 161.3
R1504 VP.n30 VP.n8 161.3
R1505 VP.n58 VP.n0 161.3
R1506 VP.n57 VP.n56 161.3
R1507 VP.n55 VP.n1 161.3
R1508 VP.n54 VP.n53 161.3
R1509 VP.n52 VP.n2 161.3
R1510 VP.n50 VP.n49 161.3
R1511 VP.n48 VP.n3 161.3
R1512 VP.n47 VP.n46 161.3
R1513 VP.n45 VP.n4 161.3
R1514 VP.n44 VP.n43 161.3
R1515 VP.n42 VP.n41 161.3
R1516 VP.n40 VP.n6 161.3
R1517 VP.n39 VP.n38 161.3
R1518 VP.n37 VP.n7 161.3
R1519 VP.n36 VP.n35 161.3
R1520 VP.n34 VP.n33 94.0526
R1521 VP.n60 VP.n59 94.0526
R1522 VP.n32 VP.n31 94.0526
R1523 VP.n14 VP.n13 57.4839
R1524 VP.n33 VP.n32 54.0753
R1525 VP.n39 VP.n7 46.253
R1526 VP.n57 VP.n1 46.253
R1527 VP.n29 VP.n9 46.253
R1528 VP.n46 VP.n45 40.4106
R1529 VP.n46 VP.n3 40.4106
R1530 VP.n18 VP.n11 40.4106
R1531 VP.n18 VP.n17 40.4106
R1532 VP.n40 VP.n39 34.5682
R1533 VP.n53 VP.n1 34.5682
R1534 VP.n25 VP.n9 34.5682
R1535 VP.n35 VP.n7 24.3439
R1536 VP.n41 VP.n40 24.3439
R1537 VP.n45 VP.n44 24.3439
R1538 VP.n50 VP.n3 24.3439
R1539 VP.n53 VP.n52 24.3439
R1540 VP.n58 VP.n57 24.3439
R1541 VP.n30 VP.n29 24.3439
R1542 VP.n22 VP.n11 24.3439
R1543 VP.n25 VP.n24 24.3439
R1544 VP.n17 VP.n16 24.3439
R1545 VP.n35 VP.n34 16.554
R1546 VP.n59 VP.n58 16.554
R1547 VP.n31 VP.n30 16.554
R1548 VP.n44 VP.n5 13.6328
R1549 VP.n51 VP.n50 13.6328
R1550 VP.n23 VP.n22 13.6328
R1551 VP.n16 VP.n13 13.6328
R1552 VP.n41 VP.n5 10.7116
R1553 VP.n52 VP.n51 10.7116
R1554 VP.n24 VP.n23 10.7116
R1555 VP.n15 VP.n14 9.31384
R1556 VP.n32 VP.n8 0.278398
R1557 VP.n36 VP.n33 0.278398
R1558 VP.n60 VP.n0 0.278398
R1559 VP.n15 VP.n12 0.189894
R1560 VP.n19 VP.n12 0.189894
R1561 VP.n20 VP.n19 0.189894
R1562 VP.n21 VP.n20 0.189894
R1563 VP.n21 VP.n10 0.189894
R1564 VP.n26 VP.n10 0.189894
R1565 VP.n27 VP.n26 0.189894
R1566 VP.n28 VP.n27 0.189894
R1567 VP.n28 VP.n8 0.189894
R1568 VP.n37 VP.n36 0.189894
R1569 VP.n38 VP.n37 0.189894
R1570 VP.n38 VP.n6 0.189894
R1571 VP.n42 VP.n6 0.189894
R1572 VP.n43 VP.n42 0.189894
R1573 VP.n43 VP.n4 0.189894
R1574 VP.n47 VP.n4 0.189894
R1575 VP.n48 VP.n47 0.189894
R1576 VP.n49 VP.n48 0.189894
R1577 VP.n49 VP.n2 0.189894
R1578 VP.n54 VP.n2 0.189894
R1579 VP.n55 VP.n54 0.189894
R1580 VP.n56 VP.n55 0.189894
R1581 VP.n56 VP.n0 0.189894
R1582 VP VP.n60 0.153422
R1583 VDD1 VDD1.n0 73.2502
R1584 VDD1.n3 VDD1.n2 73.1364
R1585 VDD1.n3 VDD1.n1 73.1364
R1586 VDD1.n5 VDD1.n4 72.0874
R1587 VDD1.n5 VDD1.n3 50.1259
R1588 VDD1.n4 VDD1.t3 1.76324
R1589 VDD1.n4 VDD1.t0 1.76324
R1590 VDD1.n0 VDD1.t6 1.76324
R1591 VDD1.n0 VDD1.t1 1.76324
R1592 VDD1.n2 VDD1.t7 1.76324
R1593 VDD1.n2 VDD1.t4 1.76324
R1594 VDD1.n1 VDD1.t5 1.76324
R1595 VDD1.n1 VDD1.t2 1.76324
R1596 VDD1 VDD1.n5 1.04576
C0 VTAIL B 6.87061f
C1 B w_n3530_n4656# 11.3547f
C2 B VN 1.2113f
C3 VDD2 VP 0.479669f
C4 VDD1 VP 13.0321f
C5 VTAIL w_n3530_n4656# 5.64599f
C6 VTAIL VN 12.7024f
C7 w_n3530_n4656# VN 7.21488f
C8 B VP 1.97572f
C9 VDD1 VDD2 1.58276f
C10 VTAIL VP 12.716499f
C11 VDD2 B 1.79556f
C12 w_n3530_n4656# VP 7.67206f
C13 VN VP 8.40828f
C14 VDD1 B 1.71117f
C15 VTAIL VDD2 10.466701f
C16 VDD2 w_n3530_n4656# 2.10226f
C17 VDD2 VN 12.7041f
C18 VDD1 VTAIL 10.4148f
C19 VDD1 w_n3530_n4656# 2.00307f
C20 VDD1 VN 0.150429f
C21 VDD2 VSUBS 1.92525f
C22 VDD1 VSUBS 2.499494f
C23 VTAIL VSUBS 1.571591f
C24 VN VSUBS 6.56353f
C25 VP VSUBS 3.443419f
C26 B VSUBS 5.130712f
C27 w_n3530_n4656# VSUBS 0.200913p
C28 VDD1.t6 VSUBS 0.389539f
C29 VDD1.t1 VSUBS 0.389539f
C30 VDD1.n0 VSUBS 3.28456f
C31 VDD1.t5 VSUBS 0.389539f
C32 VDD1.t2 VSUBS 0.389539f
C33 VDD1.n1 VSUBS 3.2832f
C34 VDD1.t7 VSUBS 0.389539f
C35 VDD1.t4 VSUBS 0.389539f
C36 VDD1.n2 VSUBS 3.2832f
C37 VDD1.n3 VSUBS 4.32512f
C38 VDD1.t3 VSUBS 0.389539f
C39 VDD1.t0 VSUBS 0.389539f
C40 VDD1.n4 VSUBS 3.2718f
C41 VDD1.n5 VSUBS 3.85481f
C42 VP.n0 VSUBS 0.03826f
C43 VP.t3 VSUBS 3.28367f
C44 VP.n1 VSUBS 0.024863f
C45 VP.n2 VSUBS 0.029018f
C46 VP.t0 VSUBS 3.28367f
C47 VP.n3 VSUBS 0.057982f
C48 VP.n4 VSUBS 0.029018f
C49 VP.t5 VSUBS 3.28367f
C50 VP.n5 VSUBS 1.14154f
C51 VP.n6 VSUBS 0.029018f
C52 VP.n7 VSUBS 0.055626f
C53 VP.n8 VSUBS 0.03826f
C54 VP.t7 VSUBS 3.28367f
C55 VP.n9 VSUBS 0.024863f
C56 VP.n10 VSUBS 0.029018f
C57 VP.t4 VSUBS 3.28367f
C58 VP.n11 VSUBS 0.057982f
C59 VP.n12 VSUBS 0.029018f
C60 VP.t6 VSUBS 3.28367f
C61 VP.n13 VSUBS 1.21894f
C62 VP.t1 VSUBS 3.4695f
C63 VP.n14 VSUBS 1.20683f
C64 VP.n15 VSUBS 0.247972f
C65 VP.n16 VSUBS 0.042546f
C66 VP.n17 VSUBS 0.057982f
C67 VP.n18 VSUBS 0.023482f
C68 VP.n19 VSUBS 0.029018f
C69 VP.n20 VSUBS 0.029018f
C70 VP.n21 VSUBS 0.029018f
C71 VP.n22 VSUBS 0.042546f
C72 VP.n23 VSUBS 1.14154f
C73 VP.n24 VSUBS 0.039326f
C74 VP.n25 VSUBS 0.058958f
C75 VP.n26 VSUBS 0.029018f
C76 VP.n27 VSUBS 0.029018f
C77 VP.n28 VSUBS 0.029018f
C78 VP.n29 VSUBS 0.055626f
C79 VP.n30 VSUBS 0.045766f
C80 VP.n31 VSUBS 1.23551f
C81 VP.n32 VSUBS 1.7996f
C82 VP.n33 VSUBS 1.81884f
C83 VP.t2 VSUBS 3.28367f
C84 VP.n34 VSUBS 1.23551f
C85 VP.n35 VSUBS 0.045766f
C86 VP.n36 VSUBS 0.03826f
C87 VP.n37 VSUBS 0.029018f
C88 VP.n38 VSUBS 0.029018f
C89 VP.n39 VSUBS 0.024863f
C90 VP.n40 VSUBS 0.058958f
C91 VP.n41 VSUBS 0.039326f
C92 VP.n42 VSUBS 0.029018f
C93 VP.n43 VSUBS 0.029018f
C94 VP.n44 VSUBS 0.042546f
C95 VP.n45 VSUBS 0.057982f
C96 VP.n46 VSUBS 0.023482f
C97 VP.n47 VSUBS 0.029018f
C98 VP.n48 VSUBS 0.029018f
C99 VP.n49 VSUBS 0.029018f
C100 VP.n50 VSUBS 0.042546f
C101 VP.n51 VSUBS 1.14154f
C102 VP.n52 VSUBS 0.039326f
C103 VP.n53 VSUBS 0.058958f
C104 VP.n54 VSUBS 0.029018f
C105 VP.n55 VSUBS 0.029018f
C106 VP.n56 VSUBS 0.029018f
C107 VP.n57 VSUBS 0.055626f
C108 VP.n58 VSUBS 0.045766f
C109 VP.n59 VSUBS 1.23551f
C110 VP.n60 VSUBS 0.039131f
C111 VTAIL.t12 VSUBS 0.34f
C112 VTAIL.t14 VSUBS 0.34f
C113 VTAIL.n0 VSUBS 2.72498f
C114 VTAIL.n1 VSUBS 0.708128f
C115 VTAIL.t9 VSUBS 3.55013f
C116 VTAIL.n2 VSUBS 0.841192f
C117 VTAIL.t5 VSUBS 3.55013f
C118 VTAIL.n3 VSUBS 0.841192f
C119 VTAIL.t4 VSUBS 0.34f
C120 VTAIL.t2 VSUBS 0.34f
C121 VTAIL.n4 VSUBS 2.72498f
C122 VTAIL.n5 VSUBS 0.869675f
C123 VTAIL.t1 VSUBS 3.55013f
C124 VTAIL.n6 VSUBS 2.48389f
C125 VTAIL.t11 VSUBS 3.55013f
C126 VTAIL.n7 VSUBS 2.48389f
C127 VTAIL.t7 VSUBS 0.34f
C128 VTAIL.t13 VSUBS 0.34f
C129 VTAIL.n8 VSUBS 2.72498f
C130 VTAIL.n9 VSUBS 0.869668f
C131 VTAIL.t10 VSUBS 3.55013f
C132 VTAIL.n10 VSUBS 0.841195f
C133 VTAIL.t6 VSUBS 3.55013f
C134 VTAIL.n11 VSUBS 0.841195f
C135 VTAIL.t0 VSUBS 0.34f
C136 VTAIL.t15 VSUBS 0.34f
C137 VTAIL.n12 VSUBS 2.72498f
C138 VTAIL.n13 VSUBS 0.869668f
C139 VTAIL.t3 VSUBS 3.55012f
C140 VTAIL.n14 VSUBS 2.4839f
C141 VTAIL.t8 VSUBS 3.55013f
C142 VTAIL.n15 VSUBS 2.47951f
C143 VDD2.t3 VSUBS 0.389519f
C144 VDD2.t2 VSUBS 0.389519f
C145 VDD2.n0 VSUBS 3.28303f
C146 VDD2.t7 VSUBS 0.389519f
C147 VDD2.t5 VSUBS 0.389519f
C148 VDD2.n1 VSUBS 3.28303f
C149 VDD2.n2 VSUBS 4.2693f
C150 VDD2.t4 VSUBS 0.389519f
C151 VDD2.t0 VSUBS 0.389519f
C152 VDD2.n3 VSUBS 3.27165f
C153 VDD2.n4 VSUBS 3.8215f
C154 VDD2.t1 VSUBS 0.389519f
C155 VDD2.t6 VSUBS 0.389519f
C156 VDD2.n5 VSUBS 3.28298f
C157 VN.n0 VSUBS 0.037491f
C158 VN.t6 VSUBS 3.21768f
C159 VN.n1 VSUBS 0.024363f
C160 VN.n2 VSUBS 0.028435f
C161 VN.t0 VSUBS 3.21768f
C162 VN.n3 VSUBS 0.056817f
C163 VN.n4 VSUBS 0.028435f
C164 VN.t2 VSUBS 3.21768f
C165 VN.n5 VSUBS 1.19444f
C166 VN.t5 VSUBS 3.39978f
C167 VN.n6 VSUBS 1.18258f
C168 VN.n7 VSUBS 0.242989f
C169 VN.n8 VSUBS 0.041691f
C170 VN.n9 VSUBS 0.056817f
C171 VN.n10 VSUBS 0.02301f
C172 VN.n11 VSUBS 0.028435f
C173 VN.n12 VSUBS 0.028435f
C174 VN.n13 VSUBS 0.028435f
C175 VN.n14 VSUBS 0.041691f
C176 VN.n15 VSUBS 1.1186f
C177 VN.n16 VSUBS 0.038535f
C178 VN.n17 VSUBS 0.057773f
C179 VN.n18 VSUBS 0.028435f
C180 VN.n19 VSUBS 0.028435f
C181 VN.n20 VSUBS 0.028435f
C182 VN.n21 VSUBS 0.054508f
C183 VN.n22 VSUBS 0.044847f
C184 VN.n23 VSUBS 1.21068f
C185 VN.n24 VSUBS 0.038344f
C186 VN.n25 VSUBS 0.037491f
C187 VN.t3 VSUBS 3.21768f
C188 VN.n26 VSUBS 0.024363f
C189 VN.n27 VSUBS 0.028435f
C190 VN.t7 VSUBS 3.21768f
C191 VN.n28 VSUBS 0.056817f
C192 VN.n29 VSUBS 0.028435f
C193 VN.t1 VSUBS 3.21768f
C194 VN.n30 VSUBS 1.19444f
C195 VN.t4 VSUBS 3.39978f
C196 VN.n31 VSUBS 1.18258f
C197 VN.n32 VSUBS 0.242989f
C198 VN.n33 VSUBS 0.041691f
C199 VN.n34 VSUBS 0.056817f
C200 VN.n35 VSUBS 0.02301f
C201 VN.n36 VSUBS 0.028435f
C202 VN.n37 VSUBS 0.028435f
C203 VN.n38 VSUBS 0.028435f
C204 VN.n39 VSUBS 0.041691f
C205 VN.n40 VSUBS 1.1186f
C206 VN.n41 VSUBS 0.038535f
C207 VN.n42 VSUBS 0.057773f
C208 VN.n43 VSUBS 0.028435f
C209 VN.n44 VSUBS 0.028435f
C210 VN.n45 VSUBS 0.028435f
C211 VN.n46 VSUBS 0.054508f
C212 VN.n47 VSUBS 0.044847f
C213 VN.n48 VSUBS 1.21068f
C214 VN.n49 VSUBS 1.77854f
C215 B.n0 VSUBS 0.005556f
C216 B.n1 VSUBS 0.005556f
C217 B.n2 VSUBS 0.008218f
C218 B.n3 VSUBS 0.006297f
C219 B.n4 VSUBS 0.006297f
C220 B.n5 VSUBS 0.006297f
C221 B.n6 VSUBS 0.006297f
C222 B.n7 VSUBS 0.006297f
C223 B.n8 VSUBS 0.006297f
C224 B.n9 VSUBS 0.006297f
C225 B.n10 VSUBS 0.006297f
C226 B.n11 VSUBS 0.006297f
C227 B.n12 VSUBS 0.006297f
C228 B.n13 VSUBS 0.006297f
C229 B.n14 VSUBS 0.006297f
C230 B.n15 VSUBS 0.006297f
C231 B.n16 VSUBS 0.006297f
C232 B.n17 VSUBS 0.006297f
C233 B.n18 VSUBS 0.006297f
C234 B.n19 VSUBS 0.006297f
C235 B.n20 VSUBS 0.006297f
C236 B.n21 VSUBS 0.006297f
C237 B.n22 VSUBS 0.006297f
C238 B.n23 VSUBS 0.006297f
C239 B.n24 VSUBS 0.014411f
C240 B.n25 VSUBS 0.006297f
C241 B.n26 VSUBS 0.006297f
C242 B.n27 VSUBS 0.006297f
C243 B.n28 VSUBS 0.006297f
C244 B.n29 VSUBS 0.006297f
C245 B.n30 VSUBS 0.006297f
C246 B.n31 VSUBS 0.006297f
C247 B.n32 VSUBS 0.006297f
C248 B.n33 VSUBS 0.006297f
C249 B.n34 VSUBS 0.006297f
C250 B.n35 VSUBS 0.006297f
C251 B.n36 VSUBS 0.006297f
C252 B.n37 VSUBS 0.006297f
C253 B.n38 VSUBS 0.006297f
C254 B.n39 VSUBS 0.006297f
C255 B.n40 VSUBS 0.006297f
C256 B.n41 VSUBS 0.006297f
C257 B.n42 VSUBS 0.006297f
C258 B.n43 VSUBS 0.006297f
C259 B.n44 VSUBS 0.006297f
C260 B.n45 VSUBS 0.006297f
C261 B.n46 VSUBS 0.006297f
C262 B.n47 VSUBS 0.006297f
C263 B.n48 VSUBS 0.006297f
C264 B.n49 VSUBS 0.006297f
C265 B.n50 VSUBS 0.006297f
C266 B.n51 VSUBS 0.006297f
C267 B.n52 VSUBS 0.006297f
C268 B.n53 VSUBS 0.006297f
C269 B.n54 VSUBS 0.006297f
C270 B.n55 VSUBS 0.006297f
C271 B.t1 VSUBS 0.560955f
C272 B.t2 VSUBS 0.578167f
C273 B.t0 VSUBS 1.61933f
C274 B.n56 VSUBS 0.299631f
C275 B.n57 VSUBS 0.063527f
C276 B.n58 VSUBS 0.006297f
C277 B.n59 VSUBS 0.006297f
C278 B.n60 VSUBS 0.006297f
C279 B.n61 VSUBS 0.006297f
C280 B.t7 VSUBS 0.560933f
C281 B.t8 VSUBS 0.578149f
C282 B.t6 VSUBS 1.61933f
C283 B.n62 VSUBS 0.299649f
C284 B.n63 VSUBS 0.063549f
C285 B.n64 VSUBS 0.006297f
C286 B.n65 VSUBS 0.006297f
C287 B.n66 VSUBS 0.006297f
C288 B.n67 VSUBS 0.006297f
C289 B.n68 VSUBS 0.006297f
C290 B.n69 VSUBS 0.006297f
C291 B.n70 VSUBS 0.006297f
C292 B.n71 VSUBS 0.006297f
C293 B.n72 VSUBS 0.006297f
C294 B.n73 VSUBS 0.006297f
C295 B.n74 VSUBS 0.006297f
C296 B.n75 VSUBS 0.006297f
C297 B.n76 VSUBS 0.006297f
C298 B.n77 VSUBS 0.006297f
C299 B.n78 VSUBS 0.006297f
C300 B.n79 VSUBS 0.006297f
C301 B.n80 VSUBS 0.006297f
C302 B.n81 VSUBS 0.006297f
C303 B.n82 VSUBS 0.006297f
C304 B.n83 VSUBS 0.006297f
C305 B.n84 VSUBS 0.006297f
C306 B.n85 VSUBS 0.006297f
C307 B.n86 VSUBS 0.006297f
C308 B.n87 VSUBS 0.006297f
C309 B.n88 VSUBS 0.006297f
C310 B.n89 VSUBS 0.006297f
C311 B.n90 VSUBS 0.006297f
C312 B.n91 VSUBS 0.006297f
C313 B.n92 VSUBS 0.006297f
C314 B.n93 VSUBS 0.006297f
C315 B.n94 VSUBS 0.014411f
C316 B.n95 VSUBS 0.006297f
C317 B.n96 VSUBS 0.006297f
C318 B.n97 VSUBS 0.006297f
C319 B.n98 VSUBS 0.006297f
C320 B.n99 VSUBS 0.006297f
C321 B.n100 VSUBS 0.006297f
C322 B.n101 VSUBS 0.006297f
C323 B.n102 VSUBS 0.006297f
C324 B.n103 VSUBS 0.006297f
C325 B.n104 VSUBS 0.006297f
C326 B.n105 VSUBS 0.006297f
C327 B.n106 VSUBS 0.006297f
C328 B.n107 VSUBS 0.006297f
C329 B.n108 VSUBS 0.006297f
C330 B.n109 VSUBS 0.006297f
C331 B.n110 VSUBS 0.006297f
C332 B.n111 VSUBS 0.006297f
C333 B.n112 VSUBS 0.006297f
C334 B.n113 VSUBS 0.006297f
C335 B.n114 VSUBS 0.006297f
C336 B.n115 VSUBS 0.006297f
C337 B.n116 VSUBS 0.006297f
C338 B.n117 VSUBS 0.006297f
C339 B.n118 VSUBS 0.006297f
C340 B.n119 VSUBS 0.006297f
C341 B.n120 VSUBS 0.006297f
C342 B.n121 VSUBS 0.006297f
C343 B.n122 VSUBS 0.006297f
C344 B.n123 VSUBS 0.006297f
C345 B.n124 VSUBS 0.006297f
C346 B.n125 VSUBS 0.006297f
C347 B.n126 VSUBS 0.006297f
C348 B.n127 VSUBS 0.006297f
C349 B.n128 VSUBS 0.006297f
C350 B.n129 VSUBS 0.006297f
C351 B.n130 VSUBS 0.006297f
C352 B.n131 VSUBS 0.006297f
C353 B.n132 VSUBS 0.006297f
C354 B.n133 VSUBS 0.006297f
C355 B.n134 VSUBS 0.006297f
C356 B.n135 VSUBS 0.006297f
C357 B.n136 VSUBS 0.006297f
C358 B.n137 VSUBS 0.006297f
C359 B.n138 VSUBS 0.006297f
C360 B.n139 VSUBS 0.006297f
C361 B.n140 VSUBS 0.01487f
C362 B.n141 VSUBS 0.006297f
C363 B.n142 VSUBS 0.006297f
C364 B.n143 VSUBS 0.006297f
C365 B.n144 VSUBS 0.006297f
C366 B.n145 VSUBS 0.006297f
C367 B.n146 VSUBS 0.006297f
C368 B.n147 VSUBS 0.006297f
C369 B.n148 VSUBS 0.006297f
C370 B.n149 VSUBS 0.006297f
C371 B.n150 VSUBS 0.006297f
C372 B.n151 VSUBS 0.006297f
C373 B.n152 VSUBS 0.006297f
C374 B.n153 VSUBS 0.006297f
C375 B.n154 VSUBS 0.006297f
C376 B.n155 VSUBS 0.006297f
C377 B.n156 VSUBS 0.006297f
C378 B.n157 VSUBS 0.006297f
C379 B.n158 VSUBS 0.006297f
C380 B.n159 VSUBS 0.006297f
C381 B.n160 VSUBS 0.006297f
C382 B.n161 VSUBS 0.006297f
C383 B.n162 VSUBS 0.006297f
C384 B.n163 VSUBS 0.006297f
C385 B.n164 VSUBS 0.006297f
C386 B.n165 VSUBS 0.006297f
C387 B.n166 VSUBS 0.006297f
C388 B.n167 VSUBS 0.006297f
C389 B.n168 VSUBS 0.006297f
C390 B.n169 VSUBS 0.006297f
C391 B.n170 VSUBS 0.004353f
C392 B.n171 VSUBS 0.006297f
C393 B.n172 VSUBS 0.006297f
C394 B.n173 VSUBS 0.006297f
C395 B.n174 VSUBS 0.006297f
C396 B.n175 VSUBS 0.006297f
C397 B.t11 VSUBS 0.560955f
C398 B.t10 VSUBS 0.578167f
C399 B.t9 VSUBS 1.61933f
C400 B.n176 VSUBS 0.299631f
C401 B.n177 VSUBS 0.063527f
C402 B.n178 VSUBS 0.006297f
C403 B.n179 VSUBS 0.006297f
C404 B.n180 VSUBS 0.006297f
C405 B.n181 VSUBS 0.006297f
C406 B.n182 VSUBS 0.006297f
C407 B.n183 VSUBS 0.006297f
C408 B.n184 VSUBS 0.006297f
C409 B.n185 VSUBS 0.006297f
C410 B.n186 VSUBS 0.006297f
C411 B.n187 VSUBS 0.006297f
C412 B.n188 VSUBS 0.006297f
C413 B.n189 VSUBS 0.006297f
C414 B.n190 VSUBS 0.006297f
C415 B.n191 VSUBS 0.006297f
C416 B.n192 VSUBS 0.006297f
C417 B.n193 VSUBS 0.006297f
C418 B.n194 VSUBS 0.006297f
C419 B.n195 VSUBS 0.006297f
C420 B.n196 VSUBS 0.006297f
C421 B.n197 VSUBS 0.006297f
C422 B.n198 VSUBS 0.006297f
C423 B.n199 VSUBS 0.006297f
C424 B.n200 VSUBS 0.006297f
C425 B.n201 VSUBS 0.006297f
C426 B.n202 VSUBS 0.006297f
C427 B.n203 VSUBS 0.006297f
C428 B.n204 VSUBS 0.006297f
C429 B.n205 VSUBS 0.006297f
C430 B.n206 VSUBS 0.006297f
C431 B.n207 VSUBS 0.015594f
C432 B.n208 VSUBS 0.006297f
C433 B.n209 VSUBS 0.006297f
C434 B.n210 VSUBS 0.006297f
C435 B.n211 VSUBS 0.006297f
C436 B.n212 VSUBS 0.006297f
C437 B.n213 VSUBS 0.006297f
C438 B.n214 VSUBS 0.006297f
C439 B.n215 VSUBS 0.006297f
C440 B.n216 VSUBS 0.006297f
C441 B.n217 VSUBS 0.006297f
C442 B.n218 VSUBS 0.006297f
C443 B.n219 VSUBS 0.006297f
C444 B.n220 VSUBS 0.006297f
C445 B.n221 VSUBS 0.006297f
C446 B.n222 VSUBS 0.006297f
C447 B.n223 VSUBS 0.006297f
C448 B.n224 VSUBS 0.006297f
C449 B.n225 VSUBS 0.006297f
C450 B.n226 VSUBS 0.006297f
C451 B.n227 VSUBS 0.006297f
C452 B.n228 VSUBS 0.006297f
C453 B.n229 VSUBS 0.006297f
C454 B.n230 VSUBS 0.006297f
C455 B.n231 VSUBS 0.006297f
C456 B.n232 VSUBS 0.006297f
C457 B.n233 VSUBS 0.006297f
C458 B.n234 VSUBS 0.006297f
C459 B.n235 VSUBS 0.006297f
C460 B.n236 VSUBS 0.006297f
C461 B.n237 VSUBS 0.006297f
C462 B.n238 VSUBS 0.006297f
C463 B.n239 VSUBS 0.006297f
C464 B.n240 VSUBS 0.006297f
C465 B.n241 VSUBS 0.006297f
C466 B.n242 VSUBS 0.006297f
C467 B.n243 VSUBS 0.006297f
C468 B.n244 VSUBS 0.006297f
C469 B.n245 VSUBS 0.006297f
C470 B.n246 VSUBS 0.006297f
C471 B.n247 VSUBS 0.006297f
C472 B.n248 VSUBS 0.006297f
C473 B.n249 VSUBS 0.006297f
C474 B.n250 VSUBS 0.006297f
C475 B.n251 VSUBS 0.006297f
C476 B.n252 VSUBS 0.006297f
C477 B.n253 VSUBS 0.006297f
C478 B.n254 VSUBS 0.006297f
C479 B.n255 VSUBS 0.006297f
C480 B.n256 VSUBS 0.006297f
C481 B.n257 VSUBS 0.006297f
C482 B.n258 VSUBS 0.006297f
C483 B.n259 VSUBS 0.006297f
C484 B.n260 VSUBS 0.006297f
C485 B.n261 VSUBS 0.006297f
C486 B.n262 VSUBS 0.006297f
C487 B.n263 VSUBS 0.006297f
C488 B.n264 VSUBS 0.006297f
C489 B.n265 VSUBS 0.006297f
C490 B.n266 VSUBS 0.006297f
C491 B.n267 VSUBS 0.006297f
C492 B.n268 VSUBS 0.006297f
C493 B.n269 VSUBS 0.006297f
C494 B.n270 VSUBS 0.006297f
C495 B.n271 VSUBS 0.006297f
C496 B.n272 VSUBS 0.006297f
C497 B.n273 VSUBS 0.006297f
C498 B.n274 VSUBS 0.006297f
C499 B.n275 VSUBS 0.006297f
C500 B.n276 VSUBS 0.006297f
C501 B.n277 VSUBS 0.006297f
C502 B.n278 VSUBS 0.006297f
C503 B.n279 VSUBS 0.006297f
C504 B.n280 VSUBS 0.006297f
C505 B.n281 VSUBS 0.006297f
C506 B.n282 VSUBS 0.006297f
C507 B.n283 VSUBS 0.006297f
C508 B.n284 VSUBS 0.006297f
C509 B.n285 VSUBS 0.006297f
C510 B.n286 VSUBS 0.006297f
C511 B.n287 VSUBS 0.006297f
C512 B.n288 VSUBS 0.006297f
C513 B.n289 VSUBS 0.006297f
C514 B.n290 VSUBS 0.006297f
C515 B.n291 VSUBS 0.006297f
C516 B.n292 VSUBS 0.006297f
C517 B.n293 VSUBS 0.006297f
C518 B.n294 VSUBS 0.014411f
C519 B.n295 VSUBS 0.014411f
C520 B.n296 VSUBS 0.015594f
C521 B.n297 VSUBS 0.006297f
C522 B.n298 VSUBS 0.006297f
C523 B.n299 VSUBS 0.006297f
C524 B.n300 VSUBS 0.006297f
C525 B.n301 VSUBS 0.006297f
C526 B.n302 VSUBS 0.006297f
C527 B.n303 VSUBS 0.006297f
C528 B.n304 VSUBS 0.006297f
C529 B.n305 VSUBS 0.006297f
C530 B.n306 VSUBS 0.006297f
C531 B.n307 VSUBS 0.006297f
C532 B.n308 VSUBS 0.006297f
C533 B.n309 VSUBS 0.006297f
C534 B.n310 VSUBS 0.006297f
C535 B.n311 VSUBS 0.006297f
C536 B.n312 VSUBS 0.006297f
C537 B.n313 VSUBS 0.006297f
C538 B.n314 VSUBS 0.006297f
C539 B.n315 VSUBS 0.006297f
C540 B.n316 VSUBS 0.006297f
C541 B.n317 VSUBS 0.006297f
C542 B.n318 VSUBS 0.006297f
C543 B.n319 VSUBS 0.006297f
C544 B.n320 VSUBS 0.006297f
C545 B.n321 VSUBS 0.006297f
C546 B.n322 VSUBS 0.006297f
C547 B.n323 VSUBS 0.006297f
C548 B.n324 VSUBS 0.006297f
C549 B.n325 VSUBS 0.006297f
C550 B.n326 VSUBS 0.006297f
C551 B.n327 VSUBS 0.006297f
C552 B.n328 VSUBS 0.006297f
C553 B.n329 VSUBS 0.006297f
C554 B.n330 VSUBS 0.006297f
C555 B.n331 VSUBS 0.006297f
C556 B.n332 VSUBS 0.006297f
C557 B.n333 VSUBS 0.006297f
C558 B.n334 VSUBS 0.006297f
C559 B.n335 VSUBS 0.006297f
C560 B.n336 VSUBS 0.006297f
C561 B.n337 VSUBS 0.006297f
C562 B.n338 VSUBS 0.006297f
C563 B.n339 VSUBS 0.006297f
C564 B.n340 VSUBS 0.006297f
C565 B.n341 VSUBS 0.006297f
C566 B.n342 VSUBS 0.006297f
C567 B.n343 VSUBS 0.006297f
C568 B.n344 VSUBS 0.006297f
C569 B.n345 VSUBS 0.006297f
C570 B.n346 VSUBS 0.006297f
C571 B.n347 VSUBS 0.006297f
C572 B.n348 VSUBS 0.006297f
C573 B.n349 VSUBS 0.006297f
C574 B.n350 VSUBS 0.006297f
C575 B.n351 VSUBS 0.006297f
C576 B.n352 VSUBS 0.006297f
C577 B.n353 VSUBS 0.006297f
C578 B.n354 VSUBS 0.006297f
C579 B.n355 VSUBS 0.006297f
C580 B.n356 VSUBS 0.006297f
C581 B.n357 VSUBS 0.006297f
C582 B.n358 VSUBS 0.006297f
C583 B.n359 VSUBS 0.006297f
C584 B.n360 VSUBS 0.006297f
C585 B.n361 VSUBS 0.006297f
C586 B.n362 VSUBS 0.006297f
C587 B.n363 VSUBS 0.006297f
C588 B.n364 VSUBS 0.006297f
C589 B.n365 VSUBS 0.006297f
C590 B.n366 VSUBS 0.006297f
C591 B.n367 VSUBS 0.006297f
C592 B.n368 VSUBS 0.006297f
C593 B.n369 VSUBS 0.006297f
C594 B.n370 VSUBS 0.006297f
C595 B.n371 VSUBS 0.006297f
C596 B.n372 VSUBS 0.006297f
C597 B.n373 VSUBS 0.006297f
C598 B.n374 VSUBS 0.006297f
C599 B.n375 VSUBS 0.006297f
C600 B.n376 VSUBS 0.006297f
C601 B.n377 VSUBS 0.006297f
C602 B.n378 VSUBS 0.006297f
C603 B.n379 VSUBS 0.006297f
C604 B.n380 VSUBS 0.006297f
C605 B.n381 VSUBS 0.006297f
C606 B.n382 VSUBS 0.006297f
C607 B.n383 VSUBS 0.006297f
C608 B.n384 VSUBS 0.006297f
C609 B.n385 VSUBS 0.006297f
C610 B.n386 VSUBS 0.004353f
C611 B.n387 VSUBS 0.01459f
C612 B.n388 VSUBS 0.005093f
C613 B.n389 VSUBS 0.006297f
C614 B.n390 VSUBS 0.006297f
C615 B.n391 VSUBS 0.006297f
C616 B.n392 VSUBS 0.006297f
C617 B.n393 VSUBS 0.006297f
C618 B.n394 VSUBS 0.006297f
C619 B.n395 VSUBS 0.006297f
C620 B.n396 VSUBS 0.006297f
C621 B.n397 VSUBS 0.006297f
C622 B.n398 VSUBS 0.006297f
C623 B.n399 VSUBS 0.006297f
C624 B.t5 VSUBS 0.560933f
C625 B.t4 VSUBS 0.578149f
C626 B.t3 VSUBS 1.61933f
C627 B.n400 VSUBS 0.299649f
C628 B.n401 VSUBS 0.063549f
C629 B.n402 VSUBS 0.01459f
C630 B.n403 VSUBS 0.005093f
C631 B.n404 VSUBS 0.006297f
C632 B.n405 VSUBS 0.006297f
C633 B.n406 VSUBS 0.006297f
C634 B.n407 VSUBS 0.006297f
C635 B.n408 VSUBS 0.006297f
C636 B.n409 VSUBS 0.006297f
C637 B.n410 VSUBS 0.006297f
C638 B.n411 VSUBS 0.006297f
C639 B.n412 VSUBS 0.006297f
C640 B.n413 VSUBS 0.006297f
C641 B.n414 VSUBS 0.006297f
C642 B.n415 VSUBS 0.006297f
C643 B.n416 VSUBS 0.006297f
C644 B.n417 VSUBS 0.006297f
C645 B.n418 VSUBS 0.006297f
C646 B.n419 VSUBS 0.006297f
C647 B.n420 VSUBS 0.006297f
C648 B.n421 VSUBS 0.006297f
C649 B.n422 VSUBS 0.006297f
C650 B.n423 VSUBS 0.006297f
C651 B.n424 VSUBS 0.006297f
C652 B.n425 VSUBS 0.006297f
C653 B.n426 VSUBS 0.006297f
C654 B.n427 VSUBS 0.006297f
C655 B.n428 VSUBS 0.006297f
C656 B.n429 VSUBS 0.006297f
C657 B.n430 VSUBS 0.006297f
C658 B.n431 VSUBS 0.006297f
C659 B.n432 VSUBS 0.006297f
C660 B.n433 VSUBS 0.006297f
C661 B.n434 VSUBS 0.006297f
C662 B.n435 VSUBS 0.006297f
C663 B.n436 VSUBS 0.006297f
C664 B.n437 VSUBS 0.006297f
C665 B.n438 VSUBS 0.006297f
C666 B.n439 VSUBS 0.006297f
C667 B.n440 VSUBS 0.006297f
C668 B.n441 VSUBS 0.006297f
C669 B.n442 VSUBS 0.006297f
C670 B.n443 VSUBS 0.006297f
C671 B.n444 VSUBS 0.006297f
C672 B.n445 VSUBS 0.006297f
C673 B.n446 VSUBS 0.006297f
C674 B.n447 VSUBS 0.006297f
C675 B.n448 VSUBS 0.006297f
C676 B.n449 VSUBS 0.006297f
C677 B.n450 VSUBS 0.006297f
C678 B.n451 VSUBS 0.006297f
C679 B.n452 VSUBS 0.006297f
C680 B.n453 VSUBS 0.006297f
C681 B.n454 VSUBS 0.006297f
C682 B.n455 VSUBS 0.006297f
C683 B.n456 VSUBS 0.006297f
C684 B.n457 VSUBS 0.006297f
C685 B.n458 VSUBS 0.006297f
C686 B.n459 VSUBS 0.006297f
C687 B.n460 VSUBS 0.006297f
C688 B.n461 VSUBS 0.006297f
C689 B.n462 VSUBS 0.006297f
C690 B.n463 VSUBS 0.006297f
C691 B.n464 VSUBS 0.006297f
C692 B.n465 VSUBS 0.006297f
C693 B.n466 VSUBS 0.006297f
C694 B.n467 VSUBS 0.006297f
C695 B.n468 VSUBS 0.006297f
C696 B.n469 VSUBS 0.006297f
C697 B.n470 VSUBS 0.006297f
C698 B.n471 VSUBS 0.006297f
C699 B.n472 VSUBS 0.006297f
C700 B.n473 VSUBS 0.006297f
C701 B.n474 VSUBS 0.006297f
C702 B.n475 VSUBS 0.006297f
C703 B.n476 VSUBS 0.006297f
C704 B.n477 VSUBS 0.006297f
C705 B.n478 VSUBS 0.006297f
C706 B.n479 VSUBS 0.006297f
C707 B.n480 VSUBS 0.006297f
C708 B.n481 VSUBS 0.006297f
C709 B.n482 VSUBS 0.006297f
C710 B.n483 VSUBS 0.006297f
C711 B.n484 VSUBS 0.006297f
C712 B.n485 VSUBS 0.006297f
C713 B.n486 VSUBS 0.006297f
C714 B.n487 VSUBS 0.006297f
C715 B.n488 VSUBS 0.006297f
C716 B.n489 VSUBS 0.006297f
C717 B.n490 VSUBS 0.006297f
C718 B.n491 VSUBS 0.006297f
C719 B.n492 VSUBS 0.006297f
C720 B.n493 VSUBS 0.006297f
C721 B.n494 VSUBS 0.006297f
C722 B.n495 VSUBS 0.015594f
C723 B.n496 VSUBS 0.014411f
C724 B.n497 VSUBS 0.015135f
C725 B.n498 VSUBS 0.006297f
C726 B.n499 VSUBS 0.006297f
C727 B.n500 VSUBS 0.006297f
C728 B.n501 VSUBS 0.006297f
C729 B.n502 VSUBS 0.006297f
C730 B.n503 VSUBS 0.006297f
C731 B.n504 VSUBS 0.006297f
C732 B.n505 VSUBS 0.006297f
C733 B.n506 VSUBS 0.006297f
C734 B.n507 VSUBS 0.006297f
C735 B.n508 VSUBS 0.006297f
C736 B.n509 VSUBS 0.006297f
C737 B.n510 VSUBS 0.006297f
C738 B.n511 VSUBS 0.006297f
C739 B.n512 VSUBS 0.006297f
C740 B.n513 VSUBS 0.006297f
C741 B.n514 VSUBS 0.006297f
C742 B.n515 VSUBS 0.006297f
C743 B.n516 VSUBS 0.006297f
C744 B.n517 VSUBS 0.006297f
C745 B.n518 VSUBS 0.006297f
C746 B.n519 VSUBS 0.006297f
C747 B.n520 VSUBS 0.006297f
C748 B.n521 VSUBS 0.006297f
C749 B.n522 VSUBS 0.006297f
C750 B.n523 VSUBS 0.006297f
C751 B.n524 VSUBS 0.006297f
C752 B.n525 VSUBS 0.006297f
C753 B.n526 VSUBS 0.006297f
C754 B.n527 VSUBS 0.006297f
C755 B.n528 VSUBS 0.006297f
C756 B.n529 VSUBS 0.006297f
C757 B.n530 VSUBS 0.006297f
C758 B.n531 VSUBS 0.006297f
C759 B.n532 VSUBS 0.006297f
C760 B.n533 VSUBS 0.006297f
C761 B.n534 VSUBS 0.006297f
C762 B.n535 VSUBS 0.006297f
C763 B.n536 VSUBS 0.006297f
C764 B.n537 VSUBS 0.006297f
C765 B.n538 VSUBS 0.006297f
C766 B.n539 VSUBS 0.006297f
C767 B.n540 VSUBS 0.006297f
C768 B.n541 VSUBS 0.006297f
C769 B.n542 VSUBS 0.006297f
C770 B.n543 VSUBS 0.006297f
C771 B.n544 VSUBS 0.006297f
C772 B.n545 VSUBS 0.006297f
C773 B.n546 VSUBS 0.006297f
C774 B.n547 VSUBS 0.006297f
C775 B.n548 VSUBS 0.006297f
C776 B.n549 VSUBS 0.006297f
C777 B.n550 VSUBS 0.006297f
C778 B.n551 VSUBS 0.006297f
C779 B.n552 VSUBS 0.006297f
C780 B.n553 VSUBS 0.006297f
C781 B.n554 VSUBS 0.006297f
C782 B.n555 VSUBS 0.006297f
C783 B.n556 VSUBS 0.006297f
C784 B.n557 VSUBS 0.006297f
C785 B.n558 VSUBS 0.006297f
C786 B.n559 VSUBS 0.006297f
C787 B.n560 VSUBS 0.006297f
C788 B.n561 VSUBS 0.006297f
C789 B.n562 VSUBS 0.006297f
C790 B.n563 VSUBS 0.006297f
C791 B.n564 VSUBS 0.006297f
C792 B.n565 VSUBS 0.006297f
C793 B.n566 VSUBS 0.006297f
C794 B.n567 VSUBS 0.006297f
C795 B.n568 VSUBS 0.006297f
C796 B.n569 VSUBS 0.006297f
C797 B.n570 VSUBS 0.006297f
C798 B.n571 VSUBS 0.006297f
C799 B.n572 VSUBS 0.006297f
C800 B.n573 VSUBS 0.006297f
C801 B.n574 VSUBS 0.006297f
C802 B.n575 VSUBS 0.006297f
C803 B.n576 VSUBS 0.006297f
C804 B.n577 VSUBS 0.006297f
C805 B.n578 VSUBS 0.006297f
C806 B.n579 VSUBS 0.006297f
C807 B.n580 VSUBS 0.006297f
C808 B.n581 VSUBS 0.006297f
C809 B.n582 VSUBS 0.006297f
C810 B.n583 VSUBS 0.006297f
C811 B.n584 VSUBS 0.006297f
C812 B.n585 VSUBS 0.006297f
C813 B.n586 VSUBS 0.006297f
C814 B.n587 VSUBS 0.006297f
C815 B.n588 VSUBS 0.006297f
C816 B.n589 VSUBS 0.006297f
C817 B.n590 VSUBS 0.006297f
C818 B.n591 VSUBS 0.006297f
C819 B.n592 VSUBS 0.006297f
C820 B.n593 VSUBS 0.006297f
C821 B.n594 VSUBS 0.006297f
C822 B.n595 VSUBS 0.006297f
C823 B.n596 VSUBS 0.006297f
C824 B.n597 VSUBS 0.006297f
C825 B.n598 VSUBS 0.006297f
C826 B.n599 VSUBS 0.006297f
C827 B.n600 VSUBS 0.006297f
C828 B.n601 VSUBS 0.006297f
C829 B.n602 VSUBS 0.006297f
C830 B.n603 VSUBS 0.006297f
C831 B.n604 VSUBS 0.006297f
C832 B.n605 VSUBS 0.006297f
C833 B.n606 VSUBS 0.006297f
C834 B.n607 VSUBS 0.006297f
C835 B.n608 VSUBS 0.006297f
C836 B.n609 VSUBS 0.006297f
C837 B.n610 VSUBS 0.006297f
C838 B.n611 VSUBS 0.006297f
C839 B.n612 VSUBS 0.006297f
C840 B.n613 VSUBS 0.006297f
C841 B.n614 VSUBS 0.006297f
C842 B.n615 VSUBS 0.006297f
C843 B.n616 VSUBS 0.006297f
C844 B.n617 VSUBS 0.006297f
C845 B.n618 VSUBS 0.006297f
C846 B.n619 VSUBS 0.006297f
C847 B.n620 VSUBS 0.006297f
C848 B.n621 VSUBS 0.006297f
C849 B.n622 VSUBS 0.006297f
C850 B.n623 VSUBS 0.006297f
C851 B.n624 VSUBS 0.006297f
C852 B.n625 VSUBS 0.006297f
C853 B.n626 VSUBS 0.006297f
C854 B.n627 VSUBS 0.006297f
C855 B.n628 VSUBS 0.006297f
C856 B.n629 VSUBS 0.006297f
C857 B.n630 VSUBS 0.006297f
C858 B.n631 VSUBS 0.006297f
C859 B.n632 VSUBS 0.006297f
C860 B.n633 VSUBS 0.014411f
C861 B.n634 VSUBS 0.015594f
C862 B.n635 VSUBS 0.015594f
C863 B.n636 VSUBS 0.006297f
C864 B.n637 VSUBS 0.006297f
C865 B.n638 VSUBS 0.006297f
C866 B.n639 VSUBS 0.006297f
C867 B.n640 VSUBS 0.006297f
C868 B.n641 VSUBS 0.006297f
C869 B.n642 VSUBS 0.006297f
C870 B.n643 VSUBS 0.006297f
C871 B.n644 VSUBS 0.006297f
C872 B.n645 VSUBS 0.006297f
C873 B.n646 VSUBS 0.006297f
C874 B.n647 VSUBS 0.006297f
C875 B.n648 VSUBS 0.006297f
C876 B.n649 VSUBS 0.006297f
C877 B.n650 VSUBS 0.006297f
C878 B.n651 VSUBS 0.006297f
C879 B.n652 VSUBS 0.006297f
C880 B.n653 VSUBS 0.006297f
C881 B.n654 VSUBS 0.006297f
C882 B.n655 VSUBS 0.006297f
C883 B.n656 VSUBS 0.006297f
C884 B.n657 VSUBS 0.006297f
C885 B.n658 VSUBS 0.006297f
C886 B.n659 VSUBS 0.006297f
C887 B.n660 VSUBS 0.006297f
C888 B.n661 VSUBS 0.006297f
C889 B.n662 VSUBS 0.006297f
C890 B.n663 VSUBS 0.006297f
C891 B.n664 VSUBS 0.006297f
C892 B.n665 VSUBS 0.006297f
C893 B.n666 VSUBS 0.006297f
C894 B.n667 VSUBS 0.006297f
C895 B.n668 VSUBS 0.006297f
C896 B.n669 VSUBS 0.006297f
C897 B.n670 VSUBS 0.006297f
C898 B.n671 VSUBS 0.006297f
C899 B.n672 VSUBS 0.006297f
C900 B.n673 VSUBS 0.006297f
C901 B.n674 VSUBS 0.006297f
C902 B.n675 VSUBS 0.006297f
C903 B.n676 VSUBS 0.006297f
C904 B.n677 VSUBS 0.006297f
C905 B.n678 VSUBS 0.006297f
C906 B.n679 VSUBS 0.006297f
C907 B.n680 VSUBS 0.006297f
C908 B.n681 VSUBS 0.006297f
C909 B.n682 VSUBS 0.006297f
C910 B.n683 VSUBS 0.006297f
C911 B.n684 VSUBS 0.006297f
C912 B.n685 VSUBS 0.006297f
C913 B.n686 VSUBS 0.006297f
C914 B.n687 VSUBS 0.006297f
C915 B.n688 VSUBS 0.006297f
C916 B.n689 VSUBS 0.006297f
C917 B.n690 VSUBS 0.006297f
C918 B.n691 VSUBS 0.006297f
C919 B.n692 VSUBS 0.006297f
C920 B.n693 VSUBS 0.006297f
C921 B.n694 VSUBS 0.006297f
C922 B.n695 VSUBS 0.006297f
C923 B.n696 VSUBS 0.006297f
C924 B.n697 VSUBS 0.006297f
C925 B.n698 VSUBS 0.006297f
C926 B.n699 VSUBS 0.006297f
C927 B.n700 VSUBS 0.006297f
C928 B.n701 VSUBS 0.006297f
C929 B.n702 VSUBS 0.006297f
C930 B.n703 VSUBS 0.006297f
C931 B.n704 VSUBS 0.006297f
C932 B.n705 VSUBS 0.006297f
C933 B.n706 VSUBS 0.006297f
C934 B.n707 VSUBS 0.006297f
C935 B.n708 VSUBS 0.006297f
C936 B.n709 VSUBS 0.006297f
C937 B.n710 VSUBS 0.006297f
C938 B.n711 VSUBS 0.006297f
C939 B.n712 VSUBS 0.006297f
C940 B.n713 VSUBS 0.006297f
C941 B.n714 VSUBS 0.006297f
C942 B.n715 VSUBS 0.006297f
C943 B.n716 VSUBS 0.006297f
C944 B.n717 VSUBS 0.006297f
C945 B.n718 VSUBS 0.006297f
C946 B.n719 VSUBS 0.006297f
C947 B.n720 VSUBS 0.006297f
C948 B.n721 VSUBS 0.006297f
C949 B.n722 VSUBS 0.006297f
C950 B.n723 VSUBS 0.006297f
C951 B.n724 VSUBS 0.006297f
C952 B.n725 VSUBS 0.004353f
C953 B.n726 VSUBS 0.01459f
C954 B.n727 VSUBS 0.005093f
C955 B.n728 VSUBS 0.006297f
C956 B.n729 VSUBS 0.006297f
C957 B.n730 VSUBS 0.006297f
C958 B.n731 VSUBS 0.006297f
C959 B.n732 VSUBS 0.006297f
C960 B.n733 VSUBS 0.006297f
C961 B.n734 VSUBS 0.006297f
C962 B.n735 VSUBS 0.006297f
C963 B.n736 VSUBS 0.006297f
C964 B.n737 VSUBS 0.006297f
C965 B.n738 VSUBS 0.006297f
C966 B.n739 VSUBS 0.005093f
C967 B.n740 VSUBS 0.01459f
C968 B.n741 VSUBS 0.004353f
C969 B.n742 VSUBS 0.006297f
C970 B.n743 VSUBS 0.006297f
C971 B.n744 VSUBS 0.006297f
C972 B.n745 VSUBS 0.006297f
C973 B.n746 VSUBS 0.006297f
C974 B.n747 VSUBS 0.006297f
C975 B.n748 VSUBS 0.006297f
C976 B.n749 VSUBS 0.006297f
C977 B.n750 VSUBS 0.006297f
C978 B.n751 VSUBS 0.006297f
C979 B.n752 VSUBS 0.006297f
C980 B.n753 VSUBS 0.006297f
C981 B.n754 VSUBS 0.006297f
C982 B.n755 VSUBS 0.006297f
C983 B.n756 VSUBS 0.006297f
C984 B.n757 VSUBS 0.006297f
C985 B.n758 VSUBS 0.006297f
C986 B.n759 VSUBS 0.006297f
C987 B.n760 VSUBS 0.006297f
C988 B.n761 VSUBS 0.006297f
C989 B.n762 VSUBS 0.006297f
C990 B.n763 VSUBS 0.006297f
C991 B.n764 VSUBS 0.006297f
C992 B.n765 VSUBS 0.006297f
C993 B.n766 VSUBS 0.006297f
C994 B.n767 VSUBS 0.006297f
C995 B.n768 VSUBS 0.006297f
C996 B.n769 VSUBS 0.006297f
C997 B.n770 VSUBS 0.006297f
C998 B.n771 VSUBS 0.006297f
C999 B.n772 VSUBS 0.006297f
C1000 B.n773 VSUBS 0.006297f
C1001 B.n774 VSUBS 0.006297f
C1002 B.n775 VSUBS 0.006297f
C1003 B.n776 VSUBS 0.006297f
C1004 B.n777 VSUBS 0.006297f
C1005 B.n778 VSUBS 0.006297f
C1006 B.n779 VSUBS 0.006297f
C1007 B.n780 VSUBS 0.006297f
C1008 B.n781 VSUBS 0.006297f
C1009 B.n782 VSUBS 0.006297f
C1010 B.n783 VSUBS 0.006297f
C1011 B.n784 VSUBS 0.006297f
C1012 B.n785 VSUBS 0.006297f
C1013 B.n786 VSUBS 0.006297f
C1014 B.n787 VSUBS 0.006297f
C1015 B.n788 VSUBS 0.006297f
C1016 B.n789 VSUBS 0.006297f
C1017 B.n790 VSUBS 0.006297f
C1018 B.n791 VSUBS 0.006297f
C1019 B.n792 VSUBS 0.006297f
C1020 B.n793 VSUBS 0.006297f
C1021 B.n794 VSUBS 0.006297f
C1022 B.n795 VSUBS 0.006297f
C1023 B.n796 VSUBS 0.006297f
C1024 B.n797 VSUBS 0.006297f
C1025 B.n798 VSUBS 0.006297f
C1026 B.n799 VSUBS 0.006297f
C1027 B.n800 VSUBS 0.006297f
C1028 B.n801 VSUBS 0.006297f
C1029 B.n802 VSUBS 0.006297f
C1030 B.n803 VSUBS 0.006297f
C1031 B.n804 VSUBS 0.006297f
C1032 B.n805 VSUBS 0.006297f
C1033 B.n806 VSUBS 0.006297f
C1034 B.n807 VSUBS 0.006297f
C1035 B.n808 VSUBS 0.006297f
C1036 B.n809 VSUBS 0.006297f
C1037 B.n810 VSUBS 0.006297f
C1038 B.n811 VSUBS 0.006297f
C1039 B.n812 VSUBS 0.006297f
C1040 B.n813 VSUBS 0.006297f
C1041 B.n814 VSUBS 0.006297f
C1042 B.n815 VSUBS 0.006297f
C1043 B.n816 VSUBS 0.006297f
C1044 B.n817 VSUBS 0.006297f
C1045 B.n818 VSUBS 0.006297f
C1046 B.n819 VSUBS 0.006297f
C1047 B.n820 VSUBS 0.006297f
C1048 B.n821 VSUBS 0.006297f
C1049 B.n822 VSUBS 0.006297f
C1050 B.n823 VSUBS 0.006297f
C1051 B.n824 VSUBS 0.006297f
C1052 B.n825 VSUBS 0.006297f
C1053 B.n826 VSUBS 0.006297f
C1054 B.n827 VSUBS 0.006297f
C1055 B.n828 VSUBS 0.006297f
C1056 B.n829 VSUBS 0.006297f
C1057 B.n830 VSUBS 0.006297f
C1058 B.n831 VSUBS 0.015594f
C1059 B.n832 VSUBS 0.015594f
C1060 B.n833 VSUBS 0.014411f
C1061 B.n834 VSUBS 0.006297f
C1062 B.n835 VSUBS 0.006297f
C1063 B.n836 VSUBS 0.006297f
C1064 B.n837 VSUBS 0.006297f
C1065 B.n838 VSUBS 0.006297f
C1066 B.n839 VSUBS 0.006297f
C1067 B.n840 VSUBS 0.006297f
C1068 B.n841 VSUBS 0.006297f
C1069 B.n842 VSUBS 0.006297f
C1070 B.n843 VSUBS 0.006297f
C1071 B.n844 VSUBS 0.006297f
C1072 B.n845 VSUBS 0.006297f
C1073 B.n846 VSUBS 0.006297f
C1074 B.n847 VSUBS 0.006297f
C1075 B.n848 VSUBS 0.006297f
C1076 B.n849 VSUBS 0.006297f
C1077 B.n850 VSUBS 0.006297f
C1078 B.n851 VSUBS 0.006297f
C1079 B.n852 VSUBS 0.006297f
C1080 B.n853 VSUBS 0.006297f
C1081 B.n854 VSUBS 0.006297f
C1082 B.n855 VSUBS 0.006297f
C1083 B.n856 VSUBS 0.006297f
C1084 B.n857 VSUBS 0.006297f
C1085 B.n858 VSUBS 0.006297f
C1086 B.n859 VSUBS 0.006297f
C1087 B.n860 VSUBS 0.006297f
C1088 B.n861 VSUBS 0.006297f
C1089 B.n862 VSUBS 0.006297f
C1090 B.n863 VSUBS 0.006297f
C1091 B.n864 VSUBS 0.006297f
C1092 B.n865 VSUBS 0.006297f
C1093 B.n866 VSUBS 0.006297f
C1094 B.n867 VSUBS 0.006297f
C1095 B.n868 VSUBS 0.006297f
C1096 B.n869 VSUBS 0.006297f
C1097 B.n870 VSUBS 0.006297f
C1098 B.n871 VSUBS 0.006297f
C1099 B.n872 VSUBS 0.006297f
C1100 B.n873 VSUBS 0.006297f
C1101 B.n874 VSUBS 0.006297f
C1102 B.n875 VSUBS 0.006297f
C1103 B.n876 VSUBS 0.006297f
C1104 B.n877 VSUBS 0.006297f
C1105 B.n878 VSUBS 0.006297f
C1106 B.n879 VSUBS 0.006297f
C1107 B.n880 VSUBS 0.006297f
C1108 B.n881 VSUBS 0.006297f
C1109 B.n882 VSUBS 0.006297f
C1110 B.n883 VSUBS 0.006297f
C1111 B.n884 VSUBS 0.006297f
C1112 B.n885 VSUBS 0.006297f
C1113 B.n886 VSUBS 0.006297f
C1114 B.n887 VSUBS 0.006297f
C1115 B.n888 VSUBS 0.006297f
C1116 B.n889 VSUBS 0.006297f
C1117 B.n890 VSUBS 0.006297f
C1118 B.n891 VSUBS 0.006297f
C1119 B.n892 VSUBS 0.006297f
C1120 B.n893 VSUBS 0.006297f
C1121 B.n894 VSUBS 0.006297f
C1122 B.n895 VSUBS 0.006297f
C1123 B.n896 VSUBS 0.006297f
C1124 B.n897 VSUBS 0.006297f
C1125 B.n898 VSUBS 0.006297f
C1126 B.n899 VSUBS 0.008218f
C1127 B.n900 VSUBS 0.008754f
C1128 B.n901 VSUBS 0.017408f
.ends

