* NGSPICE file created from diff_pair_sample_0617.ext - technology: sky130A

.subckt diff_pair_sample_0617 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=2.84
X1 B.t11 B.t9 B.t10 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=2.84
X2 VDD1.t2 VP.t1 VTAIL.t4 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=2.84
X3 VDD2.t3 VN.t0 VTAIL.t1 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=2.84
X4 B.t8 B.t6 B.t7 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=2.84
X5 B.t5 B.t3 B.t4 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=2.84
X6 VTAIL.t0 VN.t1 VDD2.t2 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=2.84
X7 B.t2 B.t0 B.t1 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=0 ps=0 w=19.19 l=2.84
X8 VTAIL.t3 VN.t2 VDD2.t1 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=2.84
X9 VTAIL.t7 VP.t2 VDD1.t1 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=2.84
X10 VDD2.t0 VN.t3 VTAIL.t2 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=3.16635 pd=19.52 as=7.4841 ps=39.16 w=19.19 l=2.84
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n2872_n4806# sky130_fd_pr__pfet_01v8 ad=7.4841 pd=39.16 as=3.16635 ps=19.52 w=19.19 l=2.84
R0 VP.n4 VP.t3 198.16
R1 VP.n4 VP.t0 197.263
R2 VP.n5 VP.t2 162.845
R3 VP.n17 VP.t1 162.845
R4 VP.n16 VP.n0 161.3
R5 VP.n15 VP.n14 161.3
R6 VP.n13 VP.n1 161.3
R7 VP.n12 VP.n11 161.3
R8 VP.n10 VP.n2 161.3
R9 VP.n9 VP.n8 161.3
R10 VP.n7 VP.n3 161.3
R11 VP.n6 VP.n5 106.597
R12 VP.n18 VP.n17 106.597
R13 VP.n6 VP.n4 55.9485
R14 VP.n11 VP.n10 40.4934
R15 VP.n11 VP.n1 40.4934
R16 VP.n9 VP.n3 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n1 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n5 VP.n3 4.15989
R21 VP.n17 VP.n16 4.15989
R22 VP.n7 VP.n6 0.278367
R23 VP.n18 VP.n0 0.278367
R24 VP.n8 VP.n7 0.189894
R25 VP.n8 VP.n2 0.189894
R26 VP.n12 VP.n2 0.189894
R27 VP.n13 VP.n12 0.189894
R28 VP.n14 VP.n13 0.189894
R29 VP.n14 VP.n0 0.189894
R30 VP VP.n18 0.153454
R31 VTAIL.n5 VTAIL.t6 57.4456
R32 VTAIL.n4 VTAIL.t1 57.4456
R33 VTAIL.n3 VTAIL.t0 57.4456
R34 VTAIL.n6 VTAIL.t5 57.4455
R35 VTAIL.n7 VTAIL.t2 57.4455
R36 VTAIL.n0 VTAIL.t3 57.4455
R37 VTAIL.n1 VTAIL.t4 57.4455
R38 VTAIL.n2 VTAIL.t7 57.4455
R39 VTAIL.n7 VTAIL.n6 31.6427
R40 VTAIL.n3 VTAIL.n2 31.6427
R41 VTAIL.n4 VTAIL.n3 2.73326
R42 VTAIL.n6 VTAIL.n5 2.73326
R43 VTAIL.n2 VTAIL.n1 2.73326
R44 VTAIL VTAIL.n0 1.42507
R45 VTAIL VTAIL.n7 1.30869
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 VDD1 VDD1.n1 121.41
R49 VDD1 VDD1.n0 72.4886
R50 VDD1.n0 VDD1.t0 1.69435
R51 VDD1.n0 VDD1.t3 1.69435
R52 VDD1.n1 VDD1.t1 1.69435
R53 VDD1.n1 VDD1.t2 1.69435
R54 B.n585 B.n584 585
R55 B.n586 B.n91 585
R56 B.n588 B.n587 585
R57 B.n589 B.n90 585
R58 B.n591 B.n590 585
R59 B.n592 B.n89 585
R60 B.n594 B.n593 585
R61 B.n595 B.n88 585
R62 B.n597 B.n596 585
R63 B.n598 B.n87 585
R64 B.n600 B.n599 585
R65 B.n601 B.n86 585
R66 B.n603 B.n602 585
R67 B.n604 B.n85 585
R68 B.n606 B.n605 585
R69 B.n607 B.n84 585
R70 B.n609 B.n608 585
R71 B.n610 B.n83 585
R72 B.n612 B.n611 585
R73 B.n613 B.n82 585
R74 B.n615 B.n614 585
R75 B.n616 B.n81 585
R76 B.n618 B.n617 585
R77 B.n619 B.n80 585
R78 B.n621 B.n620 585
R79 B.n622 B.n79 585
R80 B.n624 B.n623 585
R81 B.n625 B.n78 585
R82 B.n627 B.n626 585
R83 B.n628 B.n77 585
R84 B.n630 B.n629 585
R85 B.n631 B.n76 585
R86 B.n633 B.n632 585
R87 B.n634 B.n75 585
R88 B.n636 B.n635 585
R89 B.n637 B.n74 585
R90 B.n639 B.n638 585
R91 B.n640 B.n73 585
R92 B.n642 B.n641 585
R93 B.n643 B.n72 585
R94 B.n645 B.n644 585
R95 B.n646 B.n71 585
R96 B.n648 B.n647 585
R97 B.n649 B.n70 585
R98 B.n651 B.n650 585
R99 B.n652 B.n69 585
R100 B.n654 B.n653 585
R101 B.n655 B.n68 585
R102 B.n657 B.n656 585
R103 B.n658 B.n67 585
R104 B.n660 B.n659 585
R105 B.n661 B.n66 585
R106 B.n663 B.n662 585
R107 B.n664 B.n65 585
R108 B.n666 B.n665 585
R109 B.n667 B.n64 585
R110 B.n669 B.n668 585
R111 B.n670 B.n63 585
R112 B.n672 B.n671 585
R113 B.n673 B.n62 585
R114 B.n675 B.n674 585
R115 B.n676 B.n61 585
R116 B.n678 B.n677 585
R117 B.n680 B.n679 585
R118 B.n681 B.n57 585
R119 B.n683 B.n682 585
R120 B.n684 B.n56 585
R121 B.n686 B.n685 585
R122 B.n687 B.n55 585
R123 B.n689 B.n688 585
R124 B.n690 B.n54 585
R125 B.n692 B.n691 585
R126 B.n694 B.n51 585
R127 B.n696 B.n695 585
R128 B.n697 B.n50 585
R129 B.n699 B.n698 585
R130 B.n700 B.n49 585
R131 B.n702 B.n701 585
R132 B.n703 B.n48 585
R133 B.n705 B.n704 585
R134 B.n706 B.n47 585
R135 B.n708 B.n707 585
R136 B.n709 B.n46 585
R137 B.n711 B.n710 585
R138 B.n712 B.n45 585
R139 B.n714 B.n713 585
R140 B.n715 B.n44 585
R141 B.n717 B.n716 585
R142 B.n718 B.n43 585
R143 B.n720 B.n719 585
R144 B.n721 B.n42 585
R145 B.n723 B.n722 585
R146 B.n724 B.n41 585
R147 B.n726 B.n725 585
R148 B.n727 B.n40 585
R149 B.n729 B.n728 585
R150 B.n730 B.n39 585
R151 B.n732 B.n731 585
R152 B.n733 B.n38 585
R153 B.n735 B.n734 585
R154 B.n736 B.n37 585
R155 B.n738 B.n737 585
R156 B.n739 B.n36 585
R157 B.n741 B.n740 585
R158 B.n742 B.n35 585
R159 B.n744 B.n743 585
R160 B.n745 B.n34 585
R161 B.n747 B.n746 585
R162 B.n748 B.n33 585
R163 B.n750 B.n749 585
R164 B.n751 B.n32 585
R165 B.n753 B.n752 585
R166 B.n754 B.n31 585
R167 B.n756 B.n755 585
R168 B.n757 B.n30 585
R169 B.n759 B.n758 585
R170 B.n760 B.n29 585
R171 B.n762 B.n761 585
R172 B.n763 B.n28 585
R173 B.n765 B.n764 585
R174 B.n766 B.n27 585
R175 B.n768 B.n767 585
R176 B.n769 B.n26 585
R177 B.n771 B.n770 585
R178 B.n772 B.n25 585
R179 B.n774 B.n773 585
R180 B.n775 B.n24 585
R181 B.n777 B.n776 585
R182 B.n778 B.n23 585
R183 B.n780 B.n779 585
R184 B.n781 B.n22 585
R185 B.n783 B.n782 585
R186 B.n784 B.n21 585
R187 B.n786 B.n785 585
R188 B.n787 B.n20 585
R189 B.n583 B.n92 585
R190 B.n582 B.n581 585
R191 B.n580 B.n93 585
R192 B.n579 B.n578 585
R193 B.n577 B.n94 585
R194 B.n576 B.n575 585
R195 B.n574 B.n95 585
R196 B.n573 B.n572 585
R197 B.n571 B.n96 585
R198 B.n570 B.n569 585
R199 B.n568 B.n97 585
R200 B.n567 B.n566 585
R201 B.n565 B.n98 585
R202 B.n564 B.n563 585
R203 B.n562 B.n99 585
R204 B.n561 B.n560 585
R205 B.n559 B.n100 585
R206 B.n558 B.n557 585
R207 B.n556 B.n101 585
R208 B.n555 B.n554 585
R209 B.n553 B.n102 585
R210 B.n552 B.n551 585
R211 B.n550 B.n103 585
R212 B.n549 B.n548 585
R213 B.n547 B.n104 585
R214 B.n546 B.n545 585
R215 B.n544 B.n105 585
R216 B.n543 B.n542 585
R217 B.n541 B.n106 585
R218 B.n540 B.n539 585
R219 B.n538 B.n107 585
R220 B.n537 B.n536 585
R221 B.n535 B.n108 585
R222 B.n534 B.n533 585
R223 B.n532 B.n109 585
R224 B.n531 B.n530 585
R225 B.n529 B.n110 585
R226 B.n528 B.n527 585
R227 B.n526 B.n111 585
R228 B.n525 B.n524 585
R229 B.n523 B.n112 585
R230 B.n522 B.n521 585
R231 B.n520 B.n113 585
R232 B.n519 B.n518 585
R233 B.n517 B.n114 585
R234 B.n516 B.n515 585
R235 B.n514 B.n115 585
R236 B.n513 B.n512 585
R237 B.n511 B.n116 585
R238 B.n510 B.n509 585
R239 B.n508 B.n117 585
R240 B.n507 B.n506 585
R241 B.n505 B.n118 585
R242 B.n504 B.n503 585
R243 B.n502 B.n119 585
R244 B.n501 B.n500 585
R245 B.n499 B.n120 585
R246 B.n498 B.n497 585
R247 B.n496 B.n121 585
R248 B.n495 B.n494 585
R249 B.n493 B.n122 585
R250 B.n492 B.n491 585
R251 B.n490 B.n123 585
R252 B.n489 B.n488 585
R253 B.n487 B.n124 585
R254 B.n486 B.n485 585
R255 B.n484 B.n125 585
R256 B.n483 B.n482 585
R257 B.n481 B.n126 585
R258 B.n480 B.n479 585
R259 B.n478 B.n127 585
R260 B.n477 B.n476 585
R261 B.n475 B.n128 585
R262 B.n271 B.n200 585
R263 B.n273 B.n272 585
R264 B.n274 B.n199 585
R265 B.n276 B.n275 585
R266 B.n277 B.n198 585
R267 B.n279 B.n278 585
R268 B.n280 B.n197 585
R269 B.n282 B.n281 585
R270 B.n283 B.n196 585
R271 B.n285 B.n284 585
R272 B.n286 B.n195 585
R273 B.n288 B.n287 585
R274 B.n289 B.n194 585
R275 B.n291 B.n290 585
R276 B.n292 B.n193 585
R277 B.n294 B.n293 585
R278 B.n295 B.n192 585
R279 B.n297 B.n296 585
R280 B.n298 B.n191 585
R281 B.n300 B.n299 585
R282 B.n301 B.n190 585
R283 B.n303 B.n302 585
R284 B.n304 B.n189 585
R285 B.n306 B.n305 585
R286 B.n307 B.n188 585
R287 B.n309 B.n308 585
R288 B.n310 B.n187 585
R289 B.n312 B.n311 585
R290 B.n313 B.n186 585
R291 B.n315 B.n314 585
R292 B.n316 B.n185 585
R293 B.n318 B.n317 585
R294 B.n319 B.n184 585
R295 B.n321 B.n320 585
R296 B.n322 B.n183 585
R297 B.n324 B.n323 585
R298 B.n325 B.n182 585
R299 B.n327 B.n326 585
R300 B.n328 B.n181 585
R301 B.n330 B.n329 585
R302 B.n331 B.n180 585
R303 B.n333 B.n332 585
R304 B.n334 B.n179 585
R305 B.n336 B.n335 585
R306 B.n337 B.n178 585
R307 B.n339 B.n338 585
R308 B.n340 B.n177 585
R309 B.n342 B.n341 585
R310 B.n343 B.n176 585
R311 B.n345 B.n344 585
R312 B.n346 B.n175 585
R313 B.n348 B.n347 585
R314 B.n349 B.n174 585
R315 B.n351 B.n350 585
R316 B.n352 B.n173 585
R317 B.n354 B.n353 585
R318 B.n355 B.n172 585
R319 B.n357 B.n356 585
R320 B.n358 B.n171 585
R321 B.n360 B.n359 585
R322 B.n361 B.n170 585
R323 B.n363 B.n362 585
R324 B.n364 B.n167 585
R325 B.n367 B.n366 585
R326 B.n368 B.n166 585
R327 B.n370 B.n369 585
R328 B.n371 B.n165 585
R329 B.n373 B.n372 585
R330 B.n374 B.n164 585
R331 B.n376 B.n375 585
R332 B.n377 B.n163 585
R333 B.n379 B.n378 585
R334 B.n381 B.n380 585
R335 B.n382 B.n159 585
R336 B.n384 B.n383 585
R337 B.n385 B.n158 585
R338 B.n387 B.n386 585
R339 B.n388 B.n157 585
R340 B.n390 B.n389 585
R341 B.n391 B.n156 585
R342 B.n393 B.n392 585
R343 B.n394 B.n155 585
R344 B.n396 B.n395 585
R345 B.n397 B.n154 585
R346 B.n399 B.n398 585
R347 B.n400 B.n153 585
R348 B.n402 B.n401 585
R349 B.n403 B.n152 585
R350 B.n405 B.n404 585
R351 B.n406 B.n151 585
R352 B.n408 B.n407 585
R353 B.n409 B.n150 585
R354 B.n411 B.n410 585
R355 B.n412 B.n149 585
R356 B.n414 B.n413 585
R357 B.n415 B.n148 585
R358 B.n417 B.n416 585
R359 B.n418 B.n147 585
R360 B.n420 B.n419 585
R361 B.n421 B.n146 585
R362 B.n423 B.n422 585
R363 B.n424 B.n145 585
R364 B.n426 B.n425 585
R365 B.n427 B.n144 585
R366 B.n429 B.n428 585
R367 B.n430 B.n143 585
R368 B.n432 B.n431 585
R369 B.n433 B.n142 585
R370 B.n435 B.n434 585
R371 B.n436 B.n141 585
R372 B.n438 B.n437 585
R373 B.n439 B.n140 585
R374 B.n441 B.n440 585
R375 B.n442 B.n139 585
R376 B.n444 B.n443 585
R377 B.n445 B.n138 585
R378 B.n447 B.n446 585
R379 B.n448 B.n137 585
R380 B.n450 B.n449 585
R381 B.n451 B.n136 585
R382 B.n453 B.n452 585
R383 B.n454 B.n135 585
R384 B.n456 B.n455 585
R385 B.n457 B.n134 585
R386 B.n459 B.n458 585
R387 B.n460 B.n133 585
R388 B.n462 B.n461 585
R389 B.n463 B.n132 585
R390 B.n465 B.n464 585
R391 B.n466 B.n131 585
R392 B.n468 B.n467 585
R393 B.n469 B.n130 585
R394 B.n471 B.n470 585
R395 B.n472 B.n129 585
R396 B.n474 B.n473 585
R397 B.n270 B.n269 585
R398 B.n268 B.n201 585
R399 B.n267 B.n266 585
R400 B.n265 B.n202 585
R401 B.n264 B.n263 585
R402 B.n262 B.n203 585
R403 B.n261 B.n260 585
R404 B.n259 B.n204 585
R405 B.n258 B.n257 585
R406 B.n256 B.n205 585
R407 B.n255 B.n254 585
R408 B.n253 B.n206 585
R409 B.n252 B.n251 585
R410 B.n250 B.n207 585
R411 B.n249 B.n248 585
R412 B.n247 B.n208 585
R413 B.n246 B.n245 585
R414 B.n244 B.n209 585
R415 B.n243 B.n242 585
R416 B.n241 B.n210 585
R417 B.n240 B.n239 585
R418 B.n238 B.n211 585
R419 B.n237 B.n236 585
R420 B.n235 B.n212 585
R421 B.n234 B.n233 585
R422 B.n232 B.n213 585
R423 B.n231 B.n230 585
R424 B.n229 B.n214 585
R425 B.n228 B.n227 585
R426 B.n226 B.n215 585
R427 B.n225 B.n224 585
R428 B.n223 B.n216 585
R429 B.n222 B.n221 585
R430 B.n220 B.n217 585
R431 B.n219 B.n218 585
R432 B.n2 B.n0 585
R433 B.n841 B.n1 585
R434 B.n840 B.n839 585
R435 B.n838 B.n3 585
R436 B.n837 B.n836 585
R437 B.n835 B.n4 585
R438 B.n834 B.n833 585
R439 B.n832 B.n5 585
R440 B.n831 B.n830 585
R441 B.n829 B.n6 585
R442 B.n828 B.n827 585
R443 B.n826 B.n7 585
R444 B.n825 B.n824 585
R445 B.n823 B.n8 585
R446 B.n822 B.n821 585
R447 B.n820 B.n9 585
R448 B.n819 B.n818 585
R449 B.n817 B.n10 585
R450 B.n816 B.n815 585
R451 B.n814 B.n11 585
R452 B.n813 B.n812 585
R453 B.n811 B.n12 585
R454 B.n810 B.n809 585
R455 B.n808 B.n13 585
R456 B.n807 B.n806 585
R457 B.n805 B.n14 585
R458 B.n804 B.n803 585
R459 B.n802 B.n15 585
R460 B.n801 B.n800 585
R461 B.n799 B.n16 585
R462 B.n798 B.n797 585
R463 B.n796 B.n17 585
R464 B.n795 B.n794 585
R465 B.n793 B.n18 585
R466 B.n792 B.n791 585
R467 B.n790 B.n19 585
R468 B.n789 B.n788 585
R469 B.n843 B.n842 585
R470 B.n271 B.n270 521.33
R471 B.n788 B.n787 521.33
R472 B.n475 B.n474 521.33
R473 B.n584 B.n583 521.33
R474 B.n160 B.t3 371.228
R475 B.n168 B.t0 371.228
R476 B.n52 B.t6 371.228
R477 B.n58 B.t9 371.228
R478 B.n160 B.t5 170.482
R479 B.n58 B.t10 170.482
R480 B.n168 B.t2 170.457
R481 B.n52 B.t7 170.457
R482 B.n270 B.n201 163.367
R483 B.n266 B.n201 163.367
R484 B.n266 B.n265 163.367
R485 B.n265 B.n264 163.367
R486 B.n264 B.n203 163.367
R487 B.n260 B.n203 163.367
R488 B.n260 B.n259 163.367
R489 B.n259 B.n258 163.367
R490 B.n258 B.n205 163.367
R491 B.n254 B.n205 163.367
R492 B.n254 B.n253 163.367
R493 B.n253 B.n252 163.367
R494 B.n252 B.n207 163.367
R495 B.n248 B.n207 163.367
R496 B.n248 B.n247 163.367
R497 B.n247 B.n246 163.367
R498 B.n246 B.n209 163.367
R499 B.n242 B.n209 163.367
R500 B.n242 B.n241 163.367
R501 B.n241 B.n240 163.367
R502 B.n240 B.n211 163.367
R503 B.n236 B.n211 163.367
R504 B.n236 B.n235 163.367
R505 B.n235 B.n234 163.367
R506 B.n234 B.n213 163.367
R507 B.n230 B.n213 163.367
R508 B.n230 B.n229 163.367
R509 B.n229 B.n228 163.367
R510 B.n228 B.n215 163.367
R511 B.n224 B.n215 163.367
R512 B.n224 B.n223 163.367
R513 B.n223 B.n222 163.367
R514 B.n222 B.n217 163.367
R515 B.n218 B.n217 163.367
R516 B.n218 B.n2 163.367
R517 B.n842 B.n2 163.367
R518 B.n842 B.n841 163.367
R519 B.n841 B.n840 163.367
R520 B.n840 B.n3 163.367
R521 B.n836 B.n3 163.367
R522 B.n836 B.n835 163.367
R523 B.n835 B.n834 163.367
R524 B.n834 B.n5 163.367
R525 B.n830 B.n5 163.367
R526 B.n830 B.n829 163.367
R527 B.n829 B.n828 163.367
R528 B.n828 B.n7 163.367
R529 B.n824 B.n7 163.367
R530 B.n824 B.n823 163.367
R531 B.n823 B.n822 163.367
R532 B.n822 B.n9 163.367
R533 B.n818 B.n9 163.367
R534 B.n818 B.n817 163.367
R535 B.n817 B.n816 163.367
R536 B.n816 B.n11 163.367
R537 B.n812 B.n11 163.367
R538 B.n812 B.n811 163.367
R539 B.n811 B.n810 163.367
R540 B.n810 B.n13 163.367
R541 B.n806 B.n13 163.367
R542 B.n806 B.n805 163.367
R543 B.n805 B.n804 163.367
R544 B.n804 B.n15 163.367
R545 B.n800 B.n15 163.367
R546 B.n800 B.n799 163.367
R547 B.n799 B.n798 163.367
R548 B.n798 B.n17 163.367
R549 B.n794 B.n17 163.367
R550 B.n794 B.n793 163.367
R551 B.n793 B.n792 163.367
R552 B.n792 B.n19 163.367
R553 B.n788 B.n19 163.367
R554 B.n272 B.n271 163.367
R555 B.n272 B.n199 163.367
R556 B.n276 B.n199 163.367
R557 B.n277 B.n276 163.367
R558 B.n278 B.n277 163.367
R559 B.n278 B.n197 163.367
R560 B.n282 B.n197 163.367
R561 B.n283 B.n282 163.367
R562 B.n284 B.n283 163.367
R563 B.n284 B.n195 163.367
R564 B.n288 B.n195 163.367
R565 B.n289 B.n288 163.367
R566 B.n290 B.n289 163.367
R567 B.n290 B.n193 163.367
R568 B.n294 B.n193 163.367
R569 B.n295 B.n294 163.367
R570 B.n296 B.n295 163.367
R571 B.n296 B.n191 163.367
R572 B.n300 B.n191 163.367
R573 B.n301 B.n300 163.367
R574 B.n302 B.n301 163.367
R575 B.n302 B.n189 163.367
R576 B.n306 B.n189 163.367
R577 B.n307 B.n306 163.367
R578 B.n308 B.n307 163.367
R579 B.n308 B.n187 163.367
R580 B.n312 B.n187 163.367
R581 B.n313 B.n312 163.367
R582 B.n314 B.n313 163.367
R583 B.n314 B.n185 163.367
R584 B.n318 B.n185 163.367
R585 B.n319 B.n318 163.367
R586 B.n320 B.n319 163.367
R587 B.n320 B.n183 163.367
R588 B.n324 B.n183 163.367
R589 B.n325 B.n324 163.367
R590 B.n326 B.n325 163.367
R591 B.n326 B.n181 163.367
R592 B.n330 B.n181 163.367
R593 B.n331 B.n330 163.367
R594 B.n332 B.n331 163.367
R595 B.n332 B.n179 163.367
R596 B.n336 B.n179 163.367
R597 B.n337 B.n336 163.367
R598 B.n338 B.n337 163.367
R599 B.n338 B.n177 163.367
R600 B.n342 B.n177 163.367
R601 B.n343 B.n342 163.367
R602 B.n344 B.n343 163.367
R603 B.n344 B.n175 163.367
R604 B.n348 B.n175 163.367
R605 B.n349 B.n348 163.367
R606 B.n350 B.n349 163.367
R607 B.n350 B.n173 163.367
R608 B.n354 B.n173 163.367
R609 B.n355 B.n354 163.367
R610 B.n356 B.n355 163.367
R611 B.n356 B.n171 163.367
R612 B.n360 B.n171 163.367
R613 B.n361 B.n360 163.367
R614 B.n362 B.n361 163.367
R615 B.n362 B.n167 163.367
R616 B.n367 B.n167 163.367
R617 B.n368 B.n367 163.367
R618 B.n369 B.n368 163.367
R619 B.n369 B.n165 163.367
R620 B.n373 B.n165 163.367
R621 B.n374 B.n373 163.367
R622 B.n375 B.n374 163.367
R623 B.n375 B.n163 163.367
R624 B.n379 B.n163 163.367
R625 B.n380 B.n379 163.367
R626 B.n380 B.n159 163.367
R627 B.n384 B.n159 163.367
R628 B.n385 B.n384 163.367
R629 B.n386 B.n385 163.367
R630 B.n386 B.n157 163.367
R631 B.n390 B.n157 163.367
R632 B.n391 B.n390 163.367
R633 B.n392 B.n391 163.367
R634 B.n392 B.n155 163.367
R635 B.n396 B.n155 163.367
R636 B.n397 B.n396 163.367
R637 B.n398 B.n397 163.367
R638 B.n398 B.n153 163.367
R639 B.n402 B.n153 163.367
R640 B.n403 B.n402 163.367
R641 B.n404 B.n403 163.367
R642 B.n404 B.n151 163.367
R643 B.n408 B.n151 163.367
R644 B.n409 B.n408 163.367
R645 B.n410 B.n409 163.367
R646 B.n410 B.n149 163.367
R647 B.n414 B.n149 163.367
R648 B.n415 B.n414 163.367
R649 B.n416 B.n415 163.367
R650 B.n416 B.n147 163.367
R651 B.n420 B.n147 163.367
R652 B.n421 B.n420 163.367
R653 B.n422 B.n421 163.367
R654 B.n422 B.n145 163.367
R655 B.n426 B.n145 163.367
R656 B.n427 B.n426 163.367
R657 B.n428 B.n427 163.367
R658 B.n428 B.n143 163.367
R659 B.n432 B.n143 163.367
R660 B.n433 B.n432 163.367
R661 B.n434 B.n433 163.367
R662 B.n434 B.n141 163.367
R663 B.n438 B.n141 163.367
R664 B.n439 B.n438 163.367
R665 B.n440 B.n439 163.367
R666 B.n440 B.n139 163.367
R667 B.n444 B.n139 163.367
R668 B.n445 B.n444 163.367
R669 B.n446 B.n445 163.367
R670 B.n446 B.n137 163.367
R671 B.n450 B.n137 163.367
R672 B.n451 B.n450 163.367
R673 B.n452 B.n451 163.367
R674 B.n452 B.n135 163.367
R675 B.n456 B.n135 163.367
R676 B.n457 B.n456 163.367
R677 B.n458 B.n457 163.367
R678 B.n458 B.n133 163.367
R679 B.n462 B.n133 163.367
R680 B.n463 B.n462 163.367
R681 B.n464 B.n463 163.367
R682 B.n464 B.n131 163.367
R683 B.n468 B.n131 163.367
R684 B.n469 B.n468 163.367
R685 B.n470 B.n469 163.367
R686 B.n470 B.n129 163.367
R687 B.n474 B.n129 163.367
R688 B.n476 B.n475 163.367
R689 B.n476 B.n127 163.367
R690 B.n480 B.n127 163.367
R691 B.n481 B.n480 163.367
R692 B.n482 B.n481 163.367
R693 B.n482 B.n125 163.367
R694 B.n486 B.n125 163.367
R695 B.n487 B.n486 163.367
R696 B.n488 B.n487 163.367
R697 B.n488 B.n123 163.367
R698 B.n492 B.n123 163.367
R699 B.n493 B.n492 163.367
R700 B.n494 B.n493 163.367
R701 B.n494 B.n121 163.367
R702 B.n498 B.n121 163.367
R703 B.n499 B.n498 163.367
R704 B.n500 B.n499 163.367
R705 B.n500 B.n119 163.367
R706 B.n504 B.n119 163.367
R707 B.n505 B.n504 163.367
R708 B.n506 B.n505 163.367
R709 B.n506 B.n117 163.367
R710 B.n510 B.n117 163.367
R711 B.n511 B.n510 163.367
R712 B.n512 B.n511 163.367
R713 B.n512 B.n115 163.367
R714 B.n516 B.n115 163.367
R715 B.n517 B.n516 163.367
R716 B.n518 B.n517 163.367
R717 B.n518 B.n113 163.367
R718 B.n522 B.n113 163.367
R719 B.n523 B.n522 163.367
R720 B.n524 B.n523 163.367
R721 B.n524 B.n111 163.367
R722 B.n528 B.n111 163.367
R723 B.n529 B.n528 163.367
R724 B.n530 B.n529 163.367
R725 B.n530 B.n109 163.367
R726 B.n534 B.n109 163.367
R727 B.n535 B.n534 163.367
R728 B.n536 B.n535 163.367
R729 B.n536 B.n107 163.367
R730 B.n540 B.n107 163.367
R731 B.n541 B.n540 163.367
R732 B.n542 B.n541 163.367
R733 B.n542 B.n105 163.367
R734 B.n546 B.n105 163.367
R735 B.n547 B.n546 163.367
R736 B.n548 B.n547 163.367
R737 B.n548 B.n103 163.367
R738 B.n552 B.n103 163.367
R739 B.n553 B.n552 163.367
R740 B.n554 B.n553 163.367
R741 B.n554 B.n101 163.367
R742 B.n558 B.n101 163.367
R743 B.n559 B.n558 163.367
R744 B.n560 B.n559 163.367
R745 B.n560 B.n99 163.367
R746 B.n564 B.n99 163.367
R747 B.n565 B.n564 163.367
R748 B.n566 B.n565 163.367
R749 B.n566 B.n97 163.367
R750 B.n570 B.n97 163.367
R751 B.n571 B.n570 163.367
R752 B.n572 B.n571 163.367
R753 B.n572 B.n95 163.367
R754 B.n576 B.n95 163.367
R755 B.n577 B.n576 163.367
R756 B.n578 B.n577 163.367
R757 B.n578 B.n93 163.367
R758 B.n582 B.n93 163.367
R759 B.n583 B.n582 163.367
R760 B.n787 B.n786 163.367
R761 B.n786 B.n21 163.367
R762 B.n782 B.n21 163.367
R763 B.n782 B.n781 163.367
R764 B.n781 B.n780 163.367
R765 B.n780 B.n23 163.367
R766 B.n776 B.n23 163.367
R767 B.n776 B.n775 163.367
R768 B.n775 B.n774 163.367
R769 B.n774 B.n25 163.367
R770 B.n770 B.n25 163.367
R771 B.n770 B.n769 163.367
R772 B.n769 B.n768 163.367
R773 B.n768 B.n27 163.367
R774 B.n764 B.n27 163.367
R775 B.n764 B.n763 163.367
R776 B.n763 B.n762 163.367
R777 B.n762 B.n29 163.367
R778 B.n758 B.n29 163.367
R779 B.n758 B.n757 163.367
R780 B.n757 B.n756 163.367
R781 B.n756 B.n31 163.367
R782 B.n752 B.n31 163.367
R783 B.n752 B.n751 163.367
R784 B.n751 B.n750 163.367
R785 B.n750 B.n33 163.367
R786 B.n746 B.n33 163.367
R787 B.n746 B.n745 163.367
R788 B.n745 B.n744 163.367
R789 B.n744 B.n35 163.367
R790 B.n740 B.n35 163.367
R791 B.n740 B.n739 163.367
R792 B.n739 B.n738 163.367
R793 B.n738 B.n37 163.367
R794 B.n734 B.n37 163.367
R795 B.n734 B.n733 163.367
R796 B.n733 B.n732 163.367
R797 B.n732 B.n39 163.367
R798 B.n728 B.n39 163.367
R799 B.n728 B.n727 163.367
R800 B.n727 B.n726 163.367
R801 B.n726 B.n41 163.367
R802 B.n722 B.n41 163.367
R803 B.n722 B.n721 163.367
R804 B.n721 B.n720 163.367
R805 B.n720 B.n43 163.367
R806 B.n716 B.n43 163.367
R807 B.n716 B.n715 163.367
R808 B.n715 B.n714 163.367
R809 B.n714 B.n45 163.367
R810 B.n710 B.n45 163.367
R811 B.n710 B.n709 163.367
R812 B.n709 B.n708 163.367
R813 B.n708 B.n47 163.367
R814 B.n704 B.n47 163.367
R815 B.n704 B.n703 163.367
R816 B.n703 B.n702 163.367
R817 B.n702 B.n49 163.367
R818 B.n698 B.n49 163.367
R819 B.n698 B.n697 163.367
R820 B.n697 B.n696 163.367
R821 B.n696 B.n51 163.367
R822 B.n691 B.n51 163.367
R823 B.n691 B.n690 163.367
R824 B.n690 B.n689 163.367
R825 B.n689 B.n55 163.367
R826 B.n685 B.n55 163.367
R827 B.n685 B.n684 163.367
R828 B.n684 B.n683 163.367
R829 B.n683 B.n57 163.367
R830 B.n679 B.n57 163.367
R831 B.n679 B.n678 163.367
R832 B.n678 B.n61 163.367
R833 B.n674 B.n61 163.367
R834 B.n674 B.n673 163.367
R835 B.n673 B.n672 163.367
R836 B.n672 B.n63 163.367
R837 B.n668 B.n63 163.367
R838 B.n668 B.n667 163.367
R839 B.n667 B.n666 163.367
R840 B.n666 B.n65 163.367
R841 B.n662 B.n65 163.367
R842 B.n662 B.n661 163.367
R843 B.n661 B.n660 163.367
R844 B.n660 B.n67 163.367
R845 B.n656 B.n67 163.367
R846 B.n656 B.n655 163.367
R847 B.n655 B.n654 163.367
R848 B.n654 B.n69 163.367
R849 B.n650 B.n69 163.367
R850 B.n650 B.n649 163.367
R851 B.n649 B.n648 163.367
R852 B.n648 B.n71 163.367
R853 B.n644 B.n71 163.367
R854 B.n644 B.n643 163.367
R855 B.n643 B.n642 163.367
R856 B.n642 B.n73 163.367
R857 B.n638 B.n73 163.367
R858 B.n638 B.n637 163.367
R859 B.n637 B.n636 163.367
R860 B.n636 B.n75 163.367
R861 B.n632 B.n75 163.367
R862 B.n632 B.n631 163.367
R863 B.n631 B.n630 163.367
R864 B.n630 B.n77 163.367
R865 B.n626 B.n77 163.367
R866 B.n626 B.n625 163.367
R867 B.n625 B.n624 163.367
R868 B.n624 B.n79 163.367
R869 B.n620 B.n79 163.367
R870 B.n620 B.n619 163.367
R871 B.n619 B.n618 163.367
R872 B.n618 B.n81 163.367
R873 B.n614 B.n81 163.367
R874 B.n614 B.n613 163.367
R875 B.n613 B.n612 163.367
R876 B.n612 B.n83 163.367
R877 B.n608 B.n83 163.367
R878 B.n608 B.n607 163.367
R879 B.n607 B.n606 163.367
R880 B.n606 B.n85 163.367
R881 B.n602 B.n85 163.367
R882 B.n602 B.n601 163.367
R883 B.n601 B.n600 163.367
R884 B.n600 B.n87 163.367
R885 B.n596 B.n87 163.367
R886 B.n596 B.n595 163.367
R887 B.n595 B.n594 163.367
R888 B.n594 B.n89 163.367
R889 B.n590 B.n89 163.367
R890 B.n590 B.n589 163.367
R891 B.n589 B.n588 163.367
R892 B.n588 B.n91 163.367
R893 B.n584 B.n91 163.367
R894 B.n161 B.t4 109.002
R895 B.n59 B.t11 109.002
R896 B.n169 B.t1 108.978
R897 B.n53 B.t8 108.978
R898 B.n161 B.n160 61.4793
R899 B.n169 B.n168 61.4793
R900 B.n53 B.n52 61.4793
R901 B.n59 B.n58 61.4793
R902 B.n162 B.n161 59.5399
R903 B.n365 B.n169 59.5399
R904 B.n693 B.n53 59.5399
R905 B.n60 B.n59 59.5399
R906 B.n789 B.n20 33.8737
R907 B.n585 B.n92 33.8737
R908 B.n473 B.n128 33.8737
R909 B.n269 B.n200 33.8737
R910 B B.n843 18.0485
R911 B.n785 B.n20 10.6151
R912 B.n785 B.n784 10.6151
R913 B.n784 B.n783 10.6151
R914 B.n783 B.n22 10.6151
R915 B.n779 B.n22 10.6151
R916 B.n779 B.n778 10.6151
R917 B.n778 B.n777 10.6151
R918 B.n777 B.n24 10.6151
R919 B.n773 B.n24 10.6151
R920 B.n773 B.n772 10.6151
R921 B.n772 B.n771 10.6151
R922 B.n771 B.n26 10.6151
R923 B.n767 B.n26 10.6151
R924 B.n767 B.n766 10.6151
R925 B.n766 B.n765 10.6151
R926 B.n765 B.n28 10.6151
R927 B.n761 B.n28 10.6151
R928 B.n761 B.n760 10.6151
R929 B.n760 B.n759 10.6151
R930 B.n759 B.n30 10.6151
R931 B.n755 B.n30 10.6151
R932 B.n755 B.n754 10.6151
R933 B.n754 B.n753 10.6151
R934 B.n753 B.n32 10.6151
R935 B.n749 B.n32 10.6151
R936 B.n749 B.n748 10.6151
R937 B.n748 B.n747 10.6151
R938 B.n747 B.n34 10.6151
R939 B.n743 B.n34 10.6151
R940 B.n743 B.n742 10.6151
R941 B.n742 B.n741 10.6151
R942 B.n741 B.n36 10.6151
R943 B.n737 B.n36 10.6151
R944 B.n737 B.n736 10.6151
R945 B.n736 B.n735 10.6151
R946 B.n735 B.n38 10.6151
R947 B.n731 B.n38 10.6151
R948 B.n731 B.n730 10.6151
R949 B.n730 B.n729 10.6151
R950 B.n729 B.n40 10.6151
R951 B.n725 B.n40 10.6151
R952 B.n725 B.n724 10.6151
R953 B.n724 B.n723 10.6151
R954 B.n723 B.n42 10.6151
R955 B.n719 B.n42 10.6151
R956 B.n719 B.n718 10.6151
R957 B.n718 B.n717 10.6151
R958 B.n717 B.n44 10.6151
R959 B.n713 B.n44 10.6151
R960 B.n713 B.n712 10.6151
R961 B.n712 B.n711 10.6151
R962 B.n711 B.n46 10.6151
R963 B.n707 B.n46 10.6151
R964 B.n707 B.n706 10.6151
R965 B.n706 B.n705 10.6151
R966 B.n705 B.n48 10.6151
R967 B.n701 B.n48 10.6151
R968 B.n701 B.n700 10.6151
R969 B.n700 B.n699 10.6151
R970 B.n699 B.n50 10.6151
R971 B.n695 B.n50 10.6151
R972 B.n695 B.n694 10.6151
R973 B.n692 B.n54 10.6151
R974 B.n688 B.n54 10.6151
R975 B.n688 B.n687 10.6151
R976 B.n687 B.n686 10.6151
R977 B.n686 B.n56 10.6151
R978 B.n682 B.n56 10.6151
R979 B.n682 B.n681 10.6151
R980 B.n681 B.n680 10.6151
R981 B.n677 B.n676 10.6151
R982 B.n676 B.n675 10.6151
R983 B.n675 B.n62 10.6151
R984 B.n671 B.n62 10.6151
R985 B.n671 B.n670 10.6151
R986 B.n670 B.n669 10.6151
R987 B.n669 B.n64 10.6151
R988 B.n665 B.n64 10.6151
R989 B.n665 B.n664 10.6151
R990 B.n664 B.n663 10.6151
R991 B.n663 B.n66 10.6151
R992 B.n659 B.n66 10.6151
R993 B.n659 B.n658 10.6151
R994 B.n658 B.n657 10.6151
R995 B.n657 B.n68 10.6151
R996 B.n653 B.n68 10.6151
R997 B.n653 B.n652 10.6151
R998 B.n652 B.n651 10.6151
R999 B.n651 B.n70 10.6151
R1000 B.n647 B.n70 10.6151
R1001 B.n647 B.n646 10.6151
R1002 B.n646 B.n645 10.6151
R1003 B.n645 B.n72 10.6151
R1004 B.n641 B.n72 10.6151
R1005 B.n641 B.n640 10.6151
R1006 B.n640 B.n639 10.6151
R1007 B.n639 B.n74 10.6151
R1008 B.n635 B.n74 10.6151
R1009 B.n635 B.n634 10.6151
R1010 B.n634 B.n633 10.6151
R1011 B.n633 B.n76 10.6151
R1012 B.n629 B.n76 10.6151
R1013 B.n629 B.n628 10.6151
R1014 B.n628 B.n627 10.6151
R1015 B.n627 B.n78 10.6151
R1016 B.n623 B.n78 10.6151
R1017 B.n623 B.n622 10.6151
R1018 B.n622 B.n621 10.6151
R1019 B.n621 B.n80 10.6151
R1020 B.n617 B.n80 10.6151
R1021 B.n617 B.n616 10.6151
R1022 B.n616 B.n615 10.6151
R1023 B.n615 B.n82 10.6151
R1024 B.n611 B.n82 10.6151
R1025 B.n611 B.n610 10.6151
R1026 B.n610 B.n609 10.6151
R1027 B.n609 B.n84 10.6151
R1028 B.n605 B.n84 10.6151
R1029 B.n605 B.n604 10.6151
R1030 B.n604 B.n603 10.6151
R1031 B.n603 B.n86 10.6151
R1032 B.n599 B.n86 10.6151
R1033 B.n599 B.n598 10.6151
R1034 B.n598 B.n597 10.6151
R1035 B.n597 B.n88 10.6151
R1036 B.n593 B.n88 10.6151
R1037 B.n593 B.n592 10.6151
R1038 B.n592 B.n591 10.6151
R1039 B.n591 B.n90 10.6151
R1040 B.n587 B.n90 10.6151
R1041 B.n587 B.n586 10.6151
R1042 B.n586 B.n585 10.6151
R1043 B.n477 B.n128 10.6151
R1044 B.n478 B.n477 10.6151
R1045 B.n479 B.n478 10.6151
R1046 B.n479 B.n126 10.6151
R1047 B.n483 B.n126 10.6151
R1048 B.n484 B.n483 10.6151
R1049 B.n485 B.n484 10.6151
R1050 B.n485 B.n124 10.6151
R1051 B.n489 B.n124 10.6151
R1052 B.n490 B.n489 10.6151
R1053 B.n491 B.n490 10.6151
R1054 B.n491 B.n122 10.6151
R1055 B.n495 B.n122 10.6151
R1056 B.n496 B.n495 10.6151
R1057 B.n497 B.n496 10.6151
R1058 B.n497 B.n120 10.6151
R1059 B.n501 B.n120 10.6151
R1060 B.n502 B.n501 10.6151
R1061 B.n503 B.n502 10.6151
R1062 B.n503 B.n118 10.6151
R1063 B.n507 B.n118 10.6151
R1064 B.n508 B.n507 10.6151
R1065 B.n509 B.n508 10.6151
R1066 B.n509 B.n116 10.6151
R1067 B.n513 B.n116 10.6151
R1068 B.n514 B.n513 10.6151
R1069 B.n515 B.n514 10.6151
R1070 B.n515 B.n114 10.6151
R1071 B.n519 B.n114 10.6151
R1072 B.n520 B.n519 10.6151
R1073 B.n521 B.n520 10.6151
R1074 B.n521 B.n112 10.6151
R1075 B.n525 B.n112 10.6151
R1076 B.n526 B.n525 10.6151
R1077 B.n527 B.n526 10.6151
R1078 B.n527 B.n110 10.6151
R1079 B.n531 B.n110 10.6151
R1080 B.n532 B.n531 10.6151
R1081 B.n533 B.n532 10.6151
R1082 B.n533 B.n108 10.6151
R1083 B.n537 B.n108 10.6151
R1084 B.n538 B.n537 10.6151
R1085 B.n539 B.n538 10.6151
R1086 B.n539 B.n106 10.6151
R1087 B.n543 B.n106 10.6151
R1088 B.n544 B.n543 10.6151
R1089 B.n545 B.n544 10.6151
R1090 B.n545 B.n104 10.6151
R1091 B.n549 B.n104 10.6151
R1092 B.n550 B.n549 10.6151
R1093 B.n551 B.n550 10.6151
R1094 B.n551 B.n102 10.6151
R1095 B.n555 B.n102 10.6151
R1096 B.n556 B.n555 10.6151
R1097 B.n557 B.n556 10.6151
R1098 B.n557 B.n100 10.6151
R1099 B.n561 B.n100 10.6151
R1100 B.n562 B.n561 10.6151
R1101 B.n563 B.n562 10.6151
R1102 B.n563 B.n98 10.6151
R1103 B.n567 B.n98 10.6151
R1104 B.n568 B.n567 10.6151
R1105 B.n569 B.n568 10.6151
R1106 B.n569 B.n96 10.6151
R1107 B.n573 B.n96 10.6151
R1108 B.n574 B.n573 10.6151
R1109 B.n575 B.n574 10.6151
R1110 B.n575 B.n94 10.6151
R1111 B.n579 B.n94 10.6151
R1112 B.n580 B.n579 10.6151
R1113 B.n581 B.n580 10.6151
R1114 B.n581 B.n92 10.6151
R1115 B.n273 B.n200 10.6151
R1116 B.n274 B.n273 10.6151
R1117 B.n275 B.n274 10.6151
R1118 B.n275 B.n198 10.6151
R1119 B.n279 B.n198 10.6151
R1120 B.n280 B.n279 10.6151
R1121 B.n281 B.n280 10.6151
R1122 B.n281 B.n196 10.6151
R1123 B.n285 B.n196 10.6151
R1124 B.n286 B.n285 10.6151
R1125 B.n287 B.n286 10.6151
R1126 B.n287 B.n194 10.6151
R1127 B.n291 B.n194 10.6151
R1128 B.n292 B.n291 10.6151
R1129 B.n293 B.n292 10.6151
R1130 B.n293 B.n192 10.6151
R1131 B.n297 B.n192 10.6151
R1132 B.n298 B.n297 10.6151
R1133 B.n299 B.n298 10.6151
R1134 B.n299 B.n190 10.6151
R1135 B.n303 B.n190 10.6151
R1136 B.n304 B.n303 10.6151
R1137 B.n305 B.n304 10.6151
R1138 B.n305 B.n188 10.6151
R1139 B.n309 B.n188 10.6151
R1140 B.n310 B.n309 10.6151
R1141 B.n311 B.n310 10.6151
R1142 B.n311 B.n186 10.6151
R1143 B.n315 B.n186 10.6151
R1144 B.n316 B.n315 10.6151
R1145 B.n317 B.n316 10.6151
R1146 B.n317 B.n184 10.6151
R1147 B.n321 B.n184 10.6151
R1148 B.n322 B.n321 10.6151
R1149 B.n323 B.n322 10.6151
R1150 B.n323 B.n182 10.6151
R1151 B.n327 B.n182 10.6151
R1152 B.n328 B.n327 10.6151
R1153 B.n329 B.n328 10.6151
R1154 B.n329 B.n180 10.6151
R1155 B.n333 B.n180 10.6151
R1156 B.n334 B.n333 10.6151
R1157 B.n335 B.n334 10.6151
R1158 B.n335 B.n178 10.6151
R1159 B.n339 B.n178 10.6151
R1160 B.n340 B.n339 10.6151
R1161 B.n341 B.n340 10.6151
R1162 B.n341 B.n176 10.6151
R1163 B.n345 B.n176 10.6151
R1164 B.n346 B.n345 10.6151
R1165 B.n347 B.n346 10.6151
R1166 B.n347 B.n174 10.6151
R1167 B.n351 B.n174 10.6151
R1168 B.n352 B.n351 10.6151
R1169 B.n353 B.n352 10.6151
R1170 B.n353 B.n172 10.6151
R1171 B.n357 B.n172 10.6151
R1172 B.n358 B.n357 10.6151
R1173 B.n359 B.n358 10.6151
R1174 B.n359 B.n170 10.6151
R1175 B.n363 B.n170 10.6151
R1176 B.n364 B.n363 10.6151
R1177 B.n366 B.n166 10.6151
R1178 B.n370 B.n166 10.6151
R1179 B.n371 B.n370 10.6151
R1180 B.n372 B.n371 10.6151
R1181 B.n372 B.n164 10.6151
R1182 B.n376 B.n164 10.6151
R1183 B.n377 B.n376 10.6151
R1184 B.n378 B.n377 10.6151
R1185 B.n382 B.n381 10.6151
R1186 B.n383 B.n382 10.6151
R1187 B.n383 B.n158 10.6151
R1188 B.n387 B.n158 10.6151
R1189 B.n388 B.n387 10.6151
R1190 B.n389 B.n388 10.6151
R1191 B.n389 B.n156 10.6151
R1192 B.n393 B.n156 10.6151
R1193 B.n394 B.n393 10.6151
R1194 B.n395 B.n394 10.6151
R1195 B.n395 B.n154 10.6151
R1196 B.n399 B.n154 10.6151
R1197 B.n400 B.n399 10.6151
R1198 B.n401 B.n400 10.6151
R1199 B.n401 B.n152 10.6151
R1200 B.n405 B.n152 10.6151
R1201 B.n406 B.n405 10.6151
R1202 B.n407 B.n406 10.6151
R1203 B.n407 B.n150 10.6151
R1204 B.n411 B.n150 10.6151
R1205 B.n412 B.n411 10.6151
R1206 B.n413 B.n412 10.6151
R1207 B.n413 B.n148 10.6151
R1208 B.n417 B.n148 10.6151
R1209 B.n418 B.n417 10.6151
R1210 B.n419 B.n418 10.6151
R1211 B.n419 B.n146 10.6151
R1212 B.n423 B.n146 10.6151
R1213 B.n424 B.n423 10.6151
R1214 B.n425 B.n424 10.6151
R1215 B.n425 B.n144 10.6151
R1216 B.n429 B.n144 10.6151
R1217 B.n430 B.n429 10.6151
R1218 B.n431 B.n430 10.6151
R1219 B.n431 B.n142 10.6151
R1220 B.n435 B.n142 10.6151
R1221 B.n436 B.n435 10.6151
R1222 B.n437 B.n436 10.6151
R1223 B.n437 B.n140 10.6151
R1224 B.n441 B.n140 10.6151
R1225 B.n442 B.n441 10.6151
R1226 B.n443 B.n442 10.6151
R1227 B.n443 B.n138 10.6151
R1228 B.n447 B.n138 10.6151
R1229 B.n448 B.n447 10.6151
R1230 B.n449 B.n448 10.6151
R1231 B.n449 B.n136 10.6151
R1232 B.n453 B.n136 10.6151
R1233 B.n454 B.n453 10.6151
R1234 B.n455 B.n454 10.6151
R1235 B.n455 B.n134 10.6151
R1236 B.n459 B.n134 10.6151
R1237 B.n460 B.n459 10.6151
R1238 B.n461 B.n460 10.6151
R1239 B.n461 B.n132 10.6151
R1240 B.n465 B.n132 10.6151
R1241 B.n466 B.n465 10.6151
R1242 B.n467 B.n466 10.6151
R1243 B.n467 B.n130 10.6151
R1244 B.n471 B.n130 10.6151
R1245 B.n472 B.n471 10.6151
R1246 B.n473 B.n472 10.6151
R1247 B.n269 B.n268 10.6151
R1248 B.n268 B.n267 10.6151
R1249 B.n267 B.n202 10.6151
R1250 B.n263 B.n202 10.6151
R1251 B.n263 B.n262 10.6151
R1252 B.n262 B.n261 10.6151
R1253 B.n261 B.n204 10.6151
R1254 B.n257 B.n204 10.6151
R1255 B.n257 B.n256 10.6151
R1256 B.n256 B.n255 10.6151
R1257 B.n255 B.n206 10.6151
R1258 B.n251 B.n206 10.6151
R1259 B.n251 B.n250 10.6151
R1260 B.n250 B.n249 10.6151
R1261 B.n249 B.n208 10.6151
R1262 B.n245 B.n208 10.6151
R1263 B.n245 B.n244 10.6151
R1264 B.n244 B.n243 10.6151
R1265 B.n243 B.n210 10.6151
R1266 B.n239 B.n210 10.6151
R1267 B.n239 B.n238 10.6151
R1268 B.n238 B.n237 10.6151
R1269 B.n237 B.n212 10.6151
R1270 B.n233 B.n212 10.6151
R1271 B.n233 B.n232 10.6151
R1272 B.n232 B.n231 10.6151
R1273 B.n231 B.n214 10.6151
R1274 B.n227 B.n214 10.6151
R1275 B.n227 B.n226 10.6151
R1276 B.n226 B.n225 10.6151
R1277 B.n225 B.n216 10.6151
R1278 B.n221 B.n216 10.6151
R1279 B.n221 B.n220 10.6151
R1280 B.n220 B.n219 10.6151
R1281 B.n219 B.n0 10.6151
R1282 B.n839 B.n1 10.6151
R1283 B.n839 B.n838 10.6151
R1284 B.n838 B.n837 10.6151
R1285 B.n837 B.n4 10.6151
R1286 B.n833 B.n4 10.6151
R1287 B.n833 B.n832 10.6151
R1288 B.n832 B.n831 10.6151
R1289 B.n831 B.n6 10.6151
R1290 B.n827 B.n6 10.6151
R1291 B.n827 B.n826 10.6151
R1292 B.n826 B.n825 10.6151
R1293 B.n825 B.n8 10.6151
R1294 B.n821 B.n8 10.6151
R1295 B.n821 B.n820 10.6151
R1296 B.n820 B.n819 10.6151
R1297 B.n819 B.n10 10.6151
R1298 B.n815 B.n10 10.6151
R1299 B.n815 B.n814 10.6151
R1300 B.n814 B.n813 10.6151
R1301 B.n813 B.n12 10.6151
R1302 B.n809 B.n12 10.6151
R1303 B.n809 B.n808 10.6151
R1304 B.n808 B.n807 10.6151
R1305 B.n807 B.n14 10.6151
R1306 B.n803 B.n14 10.6151
R1307 B.n803 B.n802 10.6151
R1308 B.n802 B.n801 10.6151
R1309 B.n801 B.n16 10.6151
R1310 B.n797 B.n16 10.6151
R1311 B.n797 B.n796 10.6151
R1312 B.n796 B.n795 10.6151
R1313 B.n795 B.n18 10.6151
R1314 B.n791 B.n18 10.6151
R1315 B.n791 B.n790 10.6151
R1316 B.n790 B.n789 10.6151
R1317 B.n693 B.n692 6.5566
R1318 B.n680 B.n60 6.5566
R1319 B.n366 B.n365 6.5566
R1320 B.n378 B.n162 6.5566
R1321 B.n694 B.n693 4.05904
R1322 B.n677 B.n60 4.05904
R1323 B.n365 B.n364 4.05904
R1324 B.n381 B.n162 4.05904
R1325 B.n843 B.n0 2.81026
R1326 B.n843 B.n1 2.81026
R1327 VN.n0 VN.t2 198.16
R1328 VN.n1 VN.t0 198.16
R1329 VN.n0 VN.t3 197.263
R1330 VN.n1 VN.t1 197.263
R1331 VN VN.n1 56.2274
R1332 VN VN.n0 3.45085
R1333 VDD2.n2 VDD2.n0 120.885
R1334 VDD2.n2 VDD2.n1 72.4304
R1335 VDD2.n1 VDD2.t2 1.69435
R1336 VDD2.n1 VDD2.t3 1.69435
R1337 VDD2.n0 VDD2.t1 1.69435
R1338 VDD2.n0 VDD2.t0 1.69435
R1339 VDD2 VDD2.n2 0.0586897
C0 B VP 1.8535f
C1 w_n2872_n4806# VP 5.41111f
C2 VDD2 VTAIL 7.16118f
C3 VDD2 VDD1 1.08002f
C4 VDD1 VTAIL 7.10536f
C5 VDD2 B 1.55334f
C6 VDD2 w_n2872_n4806# 1.75053f
C7 B VTAIL 7.44333f
C8 w_n2872_n4806# VTAIL 5.58346f
C9 B VDD1 1.49721f
C10 w_n2872_n4806# VDD1 1.68909f
C11 VN VP 7.69416f
C12 w_n2872_n4806# B 11.556901f
C13 VDD2 VN 7.52769f
C14 VN VTAIL 7.146221f
C15 VN VDD1 0.149055f
C16 VDD2 VP 0.409415f
C17 VP VTAIL 7.16032f
C18 VN B 1.2387f
C19 VDD1 VP 7.78725f
C20 VN w_n2872_n4806# 5.0413f
C21 VDD2 VSUBS 1.15987f
C22 VDD1 VSUBS 6.76466f
C23 VTAIL VSUBS 1.581894f
C24 VN VSUBS 5.83522f
C25 VP VSUBS 2.66672f
C26 B VSUBS 5.090873f
C27 w_n2872_n4806# VSUBS 0.168632p
C28 VDD2.t1 VSUBS 0.401924f
C29 VDD2.t0 VSUBS 0.401924f
C30 VDD2.n0 VSUBS 4.36793f
C31 VDD2.t2 VSUBS 0.401924f
C32 VDD2.t3 VSUBS 0.401924f
C33 VDD2.n1 VSUBS 3.39279f
C34 VDD2.n2 VSUBS 5.09249f
C35 VN.t2 VSUBS 4.44306f
C36 VN.t3 VSUBS 4.4359f
C37 VN.n0 VSUBS 2.82245f
C38 VN.t0 VSUBS 4.44306f
C39 VN.t1 VSUBS 4.4359f
C40 VN.n1 VSUBS 4.64263f
C41 B.n0 VSUBS 0.003678f
C42 B.n1 VSUBS 0.003678f
C43 B.n2 VSUBS 0.005816f
C44 B.n3 VSUBS 0.005816f
C45 B.n4 VSUBS 0.005816f
C46 B.n5 VSUBS 0.005816f
C47 B.n6 VSUBS 0.005816f
C48 B.n7 VSUBS 0.005816f
C49 B.n8 VSUBS 0.005816f
C50 B.n9 VSUBS 0.005816f
C51 B.n10 VSUBS 0.005816f
C52 B.n11 VSUBS 0.005816f
C53 B.n12 VSUBS 0.005816f
C54 B.n13 VSUBS 0.005816f
C55 B.n14 VSUBS 0.005816f
C56 B.n15 VSUBS 0.005816f
C57 B.n16 VSUBS 0.005816f
C58 B.n17 VSUBS 0.005816f
C59 B.n18 VSUBS 0.005816f
C60 B.n19 VSUBS 0.005816f
C61 B.n20 VSUBS 0.014272f
C62 B.n21 VSUBS 0.005816f
C63 B.n22 VSUBS 0.005816f
C64 B.n23 VSUBS 0.005816f
C65 B.n24 VSUBS 0.005816f
C66 B.n25 VSUBS 0.005816f
C67 B.n26 VSUBS 0.005816f
C68 B.n27 VSUBS 0.005816f
C69 B.n28 VSUBS 0.005816f
C70 B.n29 VSUBS 0.005816f
C71 B.n30 VSUBS 0.005816f
C72 B.n31 VSUBS 0.005816f
C73 B.n32 VSUBS 0.005816f
C74 B.n33 VSUBS 0.005816f
C75 B.n34 VSUBS 0.005816f
C76 B.n35 VSUBS 0.005816f
C77 B.n36 VSUBS 0.005816f
C78 B.n37 VSUBS 0.005816f
C79 B.n38 VSUBS 0.005816f
C80 B.n39 VSUBS 0.005816f
C81 B.n40 VSUBS 0.005816f
C82 B.n41 VSUBS 0.005816f
C83 B.n42 VSUBS 0.005816f
C84 B.n43 VSUBS 0.005816f
C85 B.n44 VSUBS 0.005816f
C86 B.n45 VSUBS 0.005816f
C87 B.n46 VSUBS 0.005816f
C88 B.n47 VSUBS 0.005816f
C89 B.n48 VSUBS 0.005816f
C90 B.n49 VSUBS 0.005816f
C91 B.n50 VSUBS 0.005816f
C92 B.n51 VSUBS 0.005816f
C93 B.t8 VSUBS 0.540599f
C94 B.t7 VSUBS 0.559527f
C95 B.t6 VSUBS 2.01298f
C96 B.n52 VSUBS 0.320723f
C97 B.n53 VSUBS 0.060775f
C98 B.n54 VSUBS 0.005816f
C99 B.n55 VSUBS 0.005816f
C100 B.n56 VSUBS 0.005816f
C101 B.n57 VSUBS 0.005816f
C102 B.t11 VSUBS 0.540577f
C103 B.t10 VSUBS 0.55951f
C104 B.t9 VSUBS 2.01298f
C105 B.n58 VSUBS 0.32074f
C106 B.n59 VSUBS 0.060797f
C107 B.n60 VSUBS 0.013475f
C108 B.n61 VSUBS 0.005816f
C109 B.n62 VSUBS 0.005816f
C110 B.n63 VSUBS 0.005816f
C111 B.n64 VSUBS 0.005816f
C112 B.n65 VSUBS 0.005816f
C113 B.n66 VSUBS 0.005816f
C114 B.n67 VSUBS 0.005816f
C115 B.n68 VSUBS 0.005816f
C116 B.n69 VSUBS 0.005816f
C117 B.n70 VSUBS 0.005816f
C118 B.n71 VSUBS 0.005816f
C119 B.n72 VSUBS 0.005816f
C120 B.n73 VSUBS 0.005816f
C121 B.n74 VSUBS 0.005816f
C122 B.n75 VSUBS 0.005816f
C123 B.n76 VSUBS 0.005816f
C124 B.n77 VSUBS 0.005816f
C125 B.n78 VSUBS 0.005816f
C126 B.n79 VSUBS 0.005816f
C127 B.n80 VSUBS 0.005816f
C128 B.n81 VSUBS 0.005816f
C129 B.n82 VSUBS 0.005816f
C130 B.n83 VSUBS 0.005816f
C131 B.n84 VSUBS 0.005816f
C132 B.n85 VSUBS 0.005816f
C133 B.n86 VSUBS 0.005816f
C134 B.n87 VSUBS 0.005816f
C135 B.n88 VSUBS 0.005816f
C136 B.n89 VSUBS 0.005816f
C137 B.n90 VSUBS 0.005816f
C138 B.n91 VSUBS 0.005816f
C139 B.n92 VSUBS 0.014272f
C140 B.n93 VSUBS 0.005816f
C141 B.n94 VSUBS 0.005816f
C142 B.n95 VSUBS 0.005816f
C143 B.n96 VSUBS 0.005816f
C144 B.n97 VSUBS 0.005816f
C145 B.n98 VSUBS 0.005816f
C146 B.n99 VSUBS 0.005816f
C147 B.n100 VSUBS 0.005816f
C148 B.n101 VSUBS 0.005816f
C149 B.n102 VSUBS 0.005816f
C150 B.n103 VSUBS 0.005816f
C151 B.n104 VSUBS 0.005816f
C152 B.n105 VSUBS 0.005816f
C153 B.n106 VSUBS 0.005816f
C154 B.n107 VSUBS 0.005816f
C155 B.n108 VSUBS 0.005816f
C156 B.n109 VSUBS 0.005816f
C157 B.n110 VSUBS 0.005816f
C158 B.n111 VSUBS 0.005816f
C159 B.n112 VSUBS 0.005816f
C160 B.n113 VSUBS 0.005816f
C161 B.n114 VSUBS 0.005816f
C162 B.n115 VSUBS 0.005816f
C163 B.n116 VSUBS 0.005816f
C164 B.n117 VSUBS 0.005816f
C165 B.n118 VSUBS 0.005816f
C166 B.n119 VSUBS 0.005816f
C167 B.n120 VSUBS 0.005816f
C168 B.n121 VSUBS 0.005816f
C169 B.n122 VSUBS 0.005816f
C170 B.n123 VSUBS 0.005816f
C171 B.n124 VSUBS 0.005816f
C172 B.n125 VSUBS 0.005816f
C173 B.n126 VSUBS 0.005816f
C174 B.n127 VSUBS 0.005816f
C175 B.n128 VSUBS 0.01361f
C176 B.n129 VSUBS 0.005816f
C177 B.n130 VSUBS 0.005816f
C178 B.n131 VSUBS 0.005816f
C179 B.n132 VSUBS 0.005816f
C180 B.n133 VSUBS 0.005816f
C181 B.n134 VSUBS 0.005816f
C182 B.n135 VSUBS 0.005816f
C183 B.n136 VSUBS 0.005816f
C184 B.n137 VSUBS 0.005816f
C185 B.n138 VSUBS 0.005816f
C186 B.n139 VSUBS 0.005816f
C187 B.n140 VSUBS 0.005816f
C188 B.n141 VSUBS 0.005816f
C189 B.n142 VSUBS 0.005816f
C190 B.n143 VSUBS 0.005816f
C191 B.n144 VSUBS 0.005816f
C192 B.n145 VSUBS 0.005816f
C193 B.n146 VSUBS 0.005816f
C194 B.n147 VSUBS 0.005816f
C195 B.n148 VSUBS 0.005816f
C196 B.n149 VSUBS 0.005816f
C197 B.n150 VSUBS 0.005816f
C198 B.n151 VSUBS 0.005816f
C199 B.n152 VSUBS 0.005816f
C200 B.n153 VSUBS 0.005816f
C201 B.n154 VSUBS 0.005816f
C202 B.n155 VSUBS 0.005816f
C203 B.n156 VSUBS 0.005816f
C204 B.n157 VSUBS 0.005816f
C205 B.n158 VSUBS 0.005816f
C206 B.n159 VSUBS 0.005816f
C207 B.t4 VSUBS 0.540577f
C208 B.t5 VSUBS 0.55951f
C209 B.t3 VSUBS 2.01298f
C210 B.n160 VSUBS 0.32074f
C211 B.n161 VSUBS 0.060797f
C212 B.n162 VSUBS 0.013475f
C213 B.n163 VSUBS 0.005816f
C214 B.n164 VSUBS 0.005816f
C215 B.n165 VSUBS 0.005816f
C216 B.n166 VSUBS 0.005816f
C217 B.n167 VSUBS 0.005816f
C218 B.t1 VSUBS 0.540599f
C219 B.t2 VSUBS 0.559527f
C220 B.t0 VSUBS 2.01298f
C221 B.n168 VSUBS 0.320723f
C222 B.n169 VSUBS 0.060775f
C223 B.n170 VSUBS 0.005816f
C224 B.n171 VSUBS 0.005816f
C225 B.n172 VSUBS 0.005816f
C226 B.n173 VSUBS 0.005816f
C227 B.n174 VSUBS 0.005816f
C228 B.n175 VSUBS 0.005816f
C229 B.n176 VSUBS 0.005816f
C230 B.n177 VSUBS 0.005816f
C231 B.n178 VSUBS 0.005816f
C232 B.n179 VSUBS 0.005816f
C233 B.n180 VSUBS 0.005816f
C234 B.n181 VSUBS 0.005816f
C235 B.n182 VSUBS 0.005816f
C236 B.n183 VSUBS 0.005816f
C237 B.n184 VSUBS 0.005816f
C238 B.n185 VSUBS 0.005816f
C239 B.n186 VSUBS 0.005816f
C240 B.n187 VSUBS 0.005816f
C241 B.n188 VSUBS 0.005816f
C242 B.n189 VSUBS 0.005816f
C243 B.n190 VSUBS 0.005816f
C244 B.n191 VSUBS 0.005816f
C245 B.n192 VSUBS 0.005816f
C246 B.n193 VSUBS 0.005816f
C247 B.n194 VSUBS 0.005816f
C248 B.n195 VSUBS 0.005816f
C249 B.n196 VSUBS 0.005816f
C250 B.n197 VSUBS 0.005816f
C251 B.n198 VSUBS 0.005816f
C252 B.n199 VSUBS 0.005816f
C253 B.n200 VSUBS 0.014272f
C254 B.n201 VSUBS 0.005816f
C255 B.n202 VSUBS 0.005816f
C256 B.n203 VSUBS 0.005816f
C257 B.n204 VSUBS 0.005816f
C258 B.n205 VSUBS 0.005816f
C259 B.n206 VSUBS 0.005816f
C260 B.n207 VSUBS 0.005816f
C261 B.n208 VSUBS 0.005816f
C262 B.n209 VSUBS 0.005816f
C263 B.n210 VSUBS 0.005816f
C264 B.n211 VSUBS 0.005816f
C265 B.n212 VSUBS 0.005816f
C266 B.n213 VSUBS 0.005816f
C267 B.n214 VSUBS 0.005816f
C268 B.n215 VSUBS 0.005816f
C269 B.n216 VSUBS 0.005816f
C270 B.n217 VSUBS 0.005816f
C271 B.n218 VSUBS 0.005816f
C272 B.n219 VSUBS 0.005816f
C273 B.n220 VSUBS 0.005816f
C274 B.n221 VSUBS 0.005816f
C275 B.n222 VSUBS 0.005816f
C276 B.n223 VSUBS 0.005816f
C277 B.n224 VSUBS 0.005816f
C278 B.n225 VSUBS 0.005816f
C279 B.n226 VSUBS 0.005816f
C280 B.n227 VSUBS 0.005816f
C281 B.n228 VSUBS 0.005816f
C282 B.n229 VSUBS 0.005816f
C283 B.n230 VSUBS 0.005816f
C284 B.n231 VSUBS 0.005816f
C285 B.n232 VSUBS 0.005816f
C286 B.n233 VSUBS 0.005816f
C287 B.n234 VSUBS 0.005816f
C288 B.n235 VSUBS 0.005816f
C289 B.n236 VSUBS 0.005816f
C290 B.n237 VSUBS 0.005816f
C291 B.n238 VSUBS 0.005816f
C292 B.n239 VSUBS 0.005816f
C293 B.n240 VSUBS 0.005816f
C294 B.n241 VSUBS 0.005816f
C295 B.n242 VSUBS 0.005816f
C296 B.n243 VSUBS 0.005816f
C297 B.n244 VSUBS 0.005816f
C298 B.n245 VSUBS 0.005816f
C299 B.n246 VSUBS 0.005816f
C300 B.n247 VSUBS 0.005816f
C301 B.n248 VSUBS 0.005816f
C302 B.n249 VSUBS 0.005816f
C303 B.n250 VSUBS 0.005816f
C304 B.n251 VSUBS 0.005816f
C305 B.n252 VSUBS 0.005816f
C306 B.n253 VSUBS 0.005816f
C307 B.n254 VSUBS 0.005816f
C308 B.n255 VSUBS 0.005816f
C309 B.n256 VSUBS 0.005816f
C310 B.n257 VSUBS 0.005816f
C311 B.n258 VSUBS 0.005816f
C312 B.n259 VSUBS 0.005816f
C313 B.n260 VSUBS 0.005816f
C314 B.n261 VSUBS 0.005816f
C315 B.n262 VSUBS 0.005816f
C316 B.n263 VSUBS 0.005816f
C317 B.n264 VSUBS 0.005816f
C318 B.n265 VSUBS 0.005816f
C319 B.n266 VSUBS 0.005816f
C320 B.n267 VSUBS 0.005816f
C321 B.n268 VSUBS 0.005816f
C322 B.n269 VSUBS 0.01361f
C323 B.n270 VSUBS 0.01361f
C324 B.n271 VSUBS 0.014272f
C325 B.n272 VSUBS 0.005816f
C326 B.n273 VSUBS 0.005816f
C327 B.n274 VSUBS 0.005816f
C328 B.n275 VSUBS 0.005816f
C329 B.n276 VSUBS 0.005816f
C330 B.n277 VSUBS 0.005816f
C331 B.n278 VSUBS 0.005816f
C332 B.n279 VSUBS 0.005816f
C333 B.n280 VSUBS 0.005816f
C334 B.n281 VSUBS 0.005816f
C335 B.n282 VSUBS 0.005816f
C336 B.n283 VSUBS 0.005816f
C337 B.n284 VSUBS 0.005816f
C338 B.n285 VSUBS 0.005816f
C339 B.n286 VSUBS 0.005816f
C340 B.n287 VSUBS 0.005816f
C341 B.n288 VSUBS 0.005816f
C342 B.n289 VSUBS 0.005816f
C343 B.n290 VSUBS 0.005816f
C344 B.n291 VSUBS 0.005816f
C345 B.n292 VSUBS 0.005816f
C346 B.n293 VSUBS 0.005816f
C347 B.n294 VSUBS 0.005816f
C348 B.n295 VSUBS 0.005816f
C349 B.n296 VSUBS 0.005816f
C350 B.n297 VSUBS 0.005816f
C351 B.n298 VSUBS 0.005816f
C352 B.n299 VSUBS 0.005816f
C353 B.n300 VSUBS 0.005816f
C354 B.n301 VSUBS 0.005816f
C355 B.n302 VSUBS 0.005816f
C356 B.n303 VSUBS 0.005816f
C357 B.n304 VSUBS 0.005816f
C358 B.n305 VSUBS 0.005816f
C359 B.n306 VSUBS 0.005816f
C360 B.n307 VSUBS 0.005816f
C361 B.n308 VSUBS 0.005816f
C362 B.n309 VSUBS 0.005816f
C363 B.n310 VSUBS 0.005816f
C364 B.n311 VSUBS 0.005816f
C365 B.n312 VSUBS 0.005816f
C366 B.n313 VSUBS 0.005816f
C367 B.n314 VSUBS 0.005816f
C368 B.n315 VSUBS 0.005816f
C369 B.n316 VSUBS 0.005816f
C370 B.n317 VSUBS 0.005816f
C371 B.n318 VSUBS 0.005816f
C372 B.n319 VSUBS 0.005816f
C373 B.n320 VSUBS 0.005816f
C374 B.n321 VSUBS 0.005816f
C375 B.n322 VSUBS 0.005816f
C376 B.n323 VSUBS 0.005816f
C377 B.n324 VSUBS 0.005816f
C378 B.n325 VSUBS 0.005816f
C379 B.n326 VSUBS 0.005816f
C380 B.n327 VSUBS 0.005816f
C381 B.n328 VSUBS 0.005816f
C382 B.n329 VSUBS 0.005816f
C383 B.n330 VSUBS 0.005816f
C384 B.n331 VSUBS 0.005816f
C385 B.n332 VSUBS 0.005816f
C386 B.n333 VSUBS 0.005816f
C387 B.n334 VSUBS 0.005816f
C388 B.n335 VSUBS 0.005816f
C389 B.n336 VSUBS 0.005816f
C390 B.n337 VSUBS 0.005816f
C391 B.n338 VSUBS 0.005816f
C392 B.n339 VSUBS 0.005816f
C393 B.n340 VSUBS 0.005816f
C394 B.n341 VSUBS 0.005816f
C395 B.n342 VSUBS 0.005816f
C396 B.n343 VSUBS 0.005816f
C397 B.n344 VSUBS 0.005816f
C398 B.n345 VSUBS 0.005816f
C399 B.n346 VSUBS 0.005816f
C400 B.n347 VSUBS 0.005816f
C401 B.n348 VSUBS 0.005816f
C402 B.n349 VSUBS 0.005816f
C403 B.n350 VSUBS 0.005816f
C404 B.n351 VSUBS 0.005816f
C405 B.n352 VSUBS 0.005816f
C406 B.n353 VSUBS 0.005816f
C407 B.n354 VSUBS 0.005816f
C408 B.n355 VSUBS 0.005816f
C409 B.n356 VSUBS 0.005816f
C410 B.n357 VSUBS 0.005816f
C411 B.n358 VSUBS 0.005816f
C412 B.n359 VSUBS 0.005816f
C413 B.n360 VSUBS 0.005816f
C414 B.n361 VSUBS 0.005816f
C415 B.n362 VSUBS 0.005816f
C416 B.n363 VSUBS 0.005816f
C417 B.n364 VSUBS 0.00402f
C418 B.n365 VSUBS 0.013475f
C419 B.n366 VSUBS 0.004704f
C420 B.n367 VSUBS 0.005816f
C421 B.n368 VSUBS 0.005816f
C422 B.n369 VSUBS 0.005816f
C423 B.n370 VSUBS 0.005816f
C424 B.n371 VSUBS 0.005816f
C425 B.n372 VSUBS 0.005816f
C426 B.n373 VSUBS 0.005816f
C427 B.n374 VSUBS 0.005816f
C428 B.n375 VSUBS 0.005816f
C429 B.n376 VSUBS 0.005816f
C430 B.n377 VSUBS 0.005816f
C431 B.n378 VSUBS 0.004704f
C432 B.n379 VSUBS 0.005816f
C433 B.n380 VSUBS 0.005816f
C434 B.n381 VSUBS 0.00402f
C435 B.n382 VSUBS 0.005816f
C436 B.n383 VSUBS 0.005816f
C437 B.n384 VSUBS 0.005816f
C438 B.n385 VSUBS 0.005816f
C439 B.n386 VSUBS 0.005816f
C440 B.n387 VSUBS 0.005816f
C441 B.n388 VSUBS 0.005816f
C442 B.n389 VSUBS 0.005816f
C443 B.n390 VSUBS 0.005816f
C444 B.n391 VSUBS 0.005816f
C445 B.n392 VSUBS 0.005816f
C446 B.n393 VSUBS 0.005816f
C447 B.n394 VSUBS 0.005816f
C448 B.n395 VSUBS 0.005816f
C449 B.n396 VSUBS 0.005816f
C450 B.n397 VSUBS 0.005816f
C451 B.n398 VSUBS 0.005816f
C452 B.n399 VSUBS 0.005816f
C453 B.n400 VSUBS 0.005816f
C454 B.n401 VSUBS 0.005816f
C455 B.n402 VSUBS 0.005816f
C456 B.n403 VSUBS 0.005816f
C457 B.n404 VSUBS 0.005816f
C458 B.n405 VSUBS 0.005816f
C459 B.n406 VSUBS 0.005816f
C460 B.n407 VSUBS 0.005816f
C461 B.n408 VSUBS 0.005816f
C462 B.n409 VSUBS 0.005816f
C463 B.n410 VSUBS 0.005816f
C464 B.n411 VSUBS 0.005816f
C465 B.n412 VSUBS 0.005816f
C466 B.n413 VSUBS 0.005816f
C467 B.n414 VSUBS 0.005816f
C468 B.n415 VSUBS 0.005816f
C469 B.n416 VSUBS 0.005816f
C470 B.n417 VSUBS 0.005816f
C471 B.n418 VSUBS 0.005816f
C472 B.n419 VSUBS 0.005816f
C473 B.n420 VSUBS 0.005816f
C474 B.n421 VSUBS 0.005816f
C475 B.n422 VSUBS 0.005816f
C476 B.n423 VSUBS 0.005816f
C477 B.n424 VSUBS 0.005816f
C478 B.n425 VSUBS 0.005816f
C479 B.n426 VSUBS 0.005816f
C480 B.n427 VSUBS 0.005816f
C481 B.n428 VSUBS 0.005816f
C482 B.n429 VSUBS 0.005816f
C483 B.n430 VSUBS 0.005816f
C484 B.n431 VSUBS 0.005816f
C485 B.n432 VSUBS 0.005816f
C486 B.n433 VSUBS 0.005816f
C487 B.n434 VSUBS 0.005816f
C488 B.n435 VSUBS 0.005816f
C489 B.n436 VSUBS 0.005816f
C490 B.n437 VSUBS 0.005816f
C491 B.n438 VSUBS 0.005816f
C492 B.n439 VSUBS 0.005816f
C493 B.n440 VSUBS 0.005816f
C494 B.n441 VSUBS 0.005816f
C495 B.n442 VSUBS 0.005816f
C496 B.n443 VSUBS 0.005816f
C497 B.n444 VSUBS 0.005816f
C498 B.n445 VSUBS 0.005816f
C499 B.n446 VSUBS 0.005816f
C500 B.n447 VSUBS 0.005816f
C501 B.n448 VSUBS 0.005816f
C502 B.n449 VSUBS 0.005816f
C503 B.n450 VSUBS 0.005816f
C504 B.n451 VSUBS 0.005816f
C505 B.n452 VSUBS 0.005816f
C506 B.n453 VSUBS 0.005816f
C507 B.n454 VSUBS 0.005816f
C508 B.n455 VSUBS 0.005816f
C509 B.n456 VSUBS 0.005816f
C510 B.n457 VSUBS 0.005816f
C511 B.n458 VSUBS 0.005816f
C512 B.n459 VSUBS 0.005816f
C513 B.n460 VSUBS 0.005816f
C514 B.n461 VSUBS 0.005816f
C515 B.n462 VSUBS 0.005816f
C516 B.n463 VSUBS 0.005816f
C517 B.n464 VSUBS 0.005816f
C518 B.n465 VSUBS 0.005816f
C519 B.n466 VSUBS 0.005816f
C520 B.n467 VSUBS 0.005816f
C521 B.n468 VSUBS 0.005816f
C522 B.n469 VSUBS 0.005816f
C523 B.n470 VSUBS 0.005816f
C524 B.n471 VSUBS 0.005816f
C525 B.n472 VSUBS 0.005816f
C526 B.n473 VSUBS 0.014272f
C527 B.n474 VSUBS 0.014272f
C528 B.n475 VSUBS 0.01361f
C529 B.n476 VSUBS 0.005816f
C530 B.n477 VSUBS 0.005816f
C531 B.n478 VSUBS 0.005816f
C532 B.n479 VSUBS 0.005816f
C533 B.n480 VSUBS 0.005816f
C534 B.n481 VSUBS 0.005816f
C535 B.n482 VSUBS 0.005816f
C536 B.n483 VSUBS 0.005816f
C537 B.n484 VSUBS 0.005816f
C538 B.n485 VSUBS 0.005816f
C539 B.n486 VSUBS 0.005816f
C540 B.n487 VSUBS 0.005816f
C541 B.n488 VSUBS 0.005816f
C542 B.n489 VSUBS 0.005816f
C543 B.n490 VSUBS 0.005816f
C544 B.n491 VSUBS 0.005816f
C545 B.n492 VSUBS 0.005816f
C546 B.n493 VSUBS 0.005816f
C547 B.n494 VSUBS 0.005816f
C548 B.n495 VSUBS 0.005816f
C549 B.n496 VSUBS 0.005816f
C550 B.n497 VSUBS 0.005816f
C551 B.n498 VSUBS 0.005816f
C552 B.n499 VSUBS 0.005816f
C553 B.n500 VSUBS 0.005816f
C554 B.n501 VSUBS 0.005816f
C555 B.n502 VSUBS 0.005816f
C556 B.n503 VSUBS 0.005816f
C557 B.n504 VSUBS 0.005816f
C558 B.n505 VSUBS 0.005816f
C559 B.n506 VSUBS 0.005816f
C560 B.n507 VSUBS 0.005816f
C561 B.n508 VSUBS 0.005816f
C562 B.n509 VSUBS 0.005816f
C563 B.n510 VSUBS 0.005816f
C564 B.n511 VSUBS 0.005816f
C565 B.n512 VSUBS 0.005816f
C566 B.n513 VSUBS 0.005816f
C567 B.n514 VSUBS 0.005816f
C568 B.n515 VSUBS 0.005816f
C569 B.n516 VSUBS 0.005816f
C570 B.n517 VSUBS 0.005816f
C571 B.n518 VSUBS 0.005816f
C572 B.n519 VSUBS 0.005816f
C573 B.n520 VSUBS 0.005816f
C574 B.n521 VSUBS 0.005816f
C575 B.n522 VSUBS 0.005816f
C576 B.n523 VSUBS 0.005816f
C577 B.n524 VSUBS 0.005816f
C578 B.n525 VSUBS 0.005816f
C579 B.n526 VSUBS 0.005816f
C580 B.n527 VSUBS 0.005816f
C581 B.n528 VSUBS 0.005816f
C582 B.n529 VSUBS 0.005816f
C583 B.n530 VSUBS 0.005816f
C584 B.n531 VSUBS 0.005816f
C585 B.n532 VSUBS 0.005816f
C586 B.n533 VSUBS 0.005816f
C587 B.n534 VSUBS 0.005816f
C588 B.n535 VSUBS 0.005816f
C589 B.n536 VSUBS 0.005816f
C590 B.n537 VSUBS 0.005816f
C591 B.n538 VSUBS 0.005816f
C592 B.n539 VSUBS 0.005816f
C593 B.n540 VSUBS 0.005816f
C594 B.n541 VSUBS 0.005816f
C595 B.n542 VSUBS 0.005816f
C596 B.n543 VSUBS 0.005816f
C597 B.n544 VSUBS 0.005816f
C598 B.n545 VSUBS 0.005816f
C599 B.n546 VSUBS 0.005816f
C600 B.n547 VSUBS 0.005816f
C601 B.n548 VSUBS 0.005816f
C602 B.n549 VSUBS 0.005816f
C603 B.n550 VSUBS 0.005816f
C604 B.n551 VSUBS 0.005816f
C605 B.n552 VSUBS 0.005816f
C606 B.n553 VSUBS 0.005816f
C607 B.n554 VSUBS 0.005816f
C608 B.n555 VSUBS 0.005816f
C609 B.n556 VSUBS 0.005816f
C610 B.n557 VSUBS 0.005816f
C611 B.n558 VSUBS 0.005816f
C612 B.n559 VSUBS 0.005816f
C613 B.n560 VSUBS 0.005816f
C614 B.n561 VSUBS 0.005816f
C615 B.n562 VSUBS 0.005816f
C616 B.n563 VSUBS 0.005816f
C617 B.n564 VSUBS 0.005816f
C618 B.n565 VSUBS 0.005816f
C619 B.n566 VSUBS 0.005816f
C620 B.n567 VSUBS 0.005816f
C621 B.n568 VSUBS 0.005816f
C622 B.n569 VSUBS 0.005816f
C623 B.n570 VSUBS 0.005816f
C624 B.n571 VSUBS 0.005816f
C625 B.n572 VSUBS 0.005816f
C626 B.n573 VSUBS 0.005816f
C627 B.n574 VSUBS 0.005816f
C628 B.n575 VSUBS 0.005816f
C629 B.n576 VSUBS 0.005816f
C630 B.n577 VSUBS 0.005816f
C631 B.n578 VSUBS 0.005816f
C632 B.n579 VSUBS 0.005816f
C633 B.n580 VSUBS 0.005816f
C634 B.n581 VSUBS 0.005816f
C635 B.n582 VSUBS 0.005816f
C636 B.n583 VSUBS 0.01361f
C637 B.n584 VSUBS 0.014272f
C638 B.n585 VSUBS 0.01361f
C639 B.n586 VSUBS 0.005816f
C640 B.n587 VSUBS 0.005816f
C641 B.n588 VSUBS 0.005816f
C642 B.n589 VSUBS 0.005816f
C643 B.n590 VSUBS 0.005816f
C644 B.n591 VSUBS 0.005816f
C645 B.n592 VSUBS 0.005816f
C646 B.n593 VSUBS 0.005816f
C647 B.n594 VSUBS 0.005816f
C648 B.n595 VSUBS 0.005816f
C649 B.n596 VSUBS 0.005816f
C650 B.n597 VSUBS 0.005816f
C651 B.n598 VSUBS 0.005816f
C652 B.n599 VSUBS 0.005816f
C653 B.n600 VSUBS 0.005816f
C654 B.n601 VSUBS 0.005816f
C655 B.n602 VSUBS 0.005816f
C656 B.n603 VSUBS 0.005816f
C657 B.n604 VSUBS 0.005816f
C658 B.n605 VSUBS 0.005816f
C659 B.n606 VSUBS 0.005816f
C660 B.n607 VSUBS 0.005816f
C661 B.n608 VSUBS 0.005816f
C662 B.n609 VSUBS 0.005816f
C663 B.n610 VSUBS 0.005816f
C664 B.n611 VSUBS 0.005816f
C665 B.n612 VSUBS 0.005816f
C666 B.n613 VSUBS 0.005816f
C667 B.n614 VSUBS 0.005816f
C668 B.n615 VSUBS 0.005816f
C669 B.n616 VSUBS 0.005816f
C670 B.n617 VSUBS 0.005816f
C671 B.n618 VSUBS 0.005816f
C672 B.n619 VSUBS 0.005816f
C673 B.n620 VSUBS 0.005816f
C674 B.n621 VSUBS 0.005816f
C675 B.n622 VSUBS 0.005816f
C676 B.n623 VSUBS 0.005816f
C677 B.n624 VSUBS 0.005816f
C678 B.n625 VSUBS 0.005816f
C679 B.n626 VSUBS 0.005816f
C680 B.n627 VSUBS 0.005816f
C681 B.n628 VSUBS 0.005816f
C682 B.n629 VSUBS 0.005816f
C683 B.n630 VSUBS 0.005816f
C684 B.n631 VSUBS 0.005816f
C685 B.n632 VSUBS 0.005816f
C686 B.n633 VSUBS 0.005816f
C687 B.n634 VSUBS 0.005816f
C688 B.n635 VSUBS 0.005816f
C689 B.n636 VSUBS 0.005816f
C690 B.n637 VSUBS 0.005816f
C691 B.n638 VSUBS 0.005816f
C692 B.n639 VSUBS 0.005816f
C693 B.n640 VSUBS 0.005816f
C694 B.n641 VSUBS 0.005816f
C695 B.n642 VSUBS 0.005816f
C696 B.n643 VSUBS 0.005816f
C697 B.n644 VSUBS 0.005816f
C698 B.n645 VSUBS 0.005816f
C699 B.n646 VSUBS 0.005816f
C700 B.n647 VSUBS 0.005816f
C701 B.n648 VSUBS 0.005816f
C702 B.n649 VSUBS 0.005816f
C703 B.n650 VSUBS 0.005816f
C704 B.n651 VSUBS 0.005816f
C705 B.n652 VSUBS 0.005816f
C706 B.n653 VSUBS 0.005816f
C707 B.n654 VSUBS 0.005816f
C708 B.n655 VSUBS 0.005816f
C709 B.n656 VSUBS 0.005816f
C710 B.n657 VSUBS 0.005816f
C711 B.n658 VSUBS 0.005816f
C712 B.n659 VSUBS 0.005816f
C713 B.n660 VSUBS 0.005816f
C714 B.n661 VSUBS 0.005816f
C715 B.n662 VSUBS 0.005816f
C716 B.n663 VSUBS 0.005816f
C717 B.n664 VSUBS 0.005816f
C718 B.n665 VSUBS 0.005816f
C719 B.n666 VSUBS 0.005816f
C720 B.n667 VSUBS 0.005816f
C721 B.n668 VSUBS 0.005816f
C722 B.n669 VSUBS 0.005816f
C723 B.n670 VSUBS 0.005816f
C724 B.n671 VSUBS 0.005816f
C725 B.n672 VSUBS 0.005816f
C726 B.n673 VSUBS 0.005816f
C727 B.n674 VSUBS 0.005816f
C728 B.n675 VSUBS 0.005816f
C729 B.n676 VSUBS 0.005816f
C730 B.n677 VSUBS 0.00402f
C731 B.n678 VSUBS 0.005816f
C732 B.n679 VSUBS 0.005816f
C733 B.n680 VSUBS 0.004704f
C734 B.n681 VSUBS 0.005816f
C735 B.n682 VSUBS 0.005816f
C736 B.n683 VSUBS 0.005816f
C737 B.n684 VSUBS 0.005816f
C738 B.n685 VSUBS 0.005816f
C739 B.n686 VSUBS 0.005816f
C740 B.n687 VSUBS 0.005816f
C741 B.n688 VSUBS 0.005816f
C742 B.n689 VSUBS 0.005816f
C743 B.n690 VSUBS 0.005816f
C744 B.n691 VSUBS 0.005816f
C745 B.n692 VSUBS 0.004704f
C746 B.n693 VSUBS 0.013475f
C747 B.n694 VSUBS 0.00402f
C748 B.n695 VSUBS 0.005816f
C749 B.n696 VSUBS 0.005816f
C750 B.n697 VSUBS 0.005816f
C751 B.n698 VSUBS 0.005816f
C752 B.n699 VSUBS 0.005816f
C753 B.n700 VSUBS 0.005816f
C754 B.n701 VSUBS 0.005816f
C755 B.n702 VSUBS 0.005816f
C756 B.n703 VSUBS 0.005816f
C757 B.n704 VSUBS 0.005816f
C758 B.n705 VSUBS 0.005816f
C759 B.n706 VSUBS 0.005816f
C760 B.n707 VSUBS 0.005816f
C761 B.n708 VSUBS 0.005816f
C762 B.n709 VSUBS 0.005816f
C763 B.n710 VSUBS 0.005816f
C764 B.n711 VSUBS 0.005816f
C765 B.n712 VSUBS 0.005816f
C766 B.n713 VSUBS 0.005816f
C767 B.n714 VSUBS 0.005816f
C768 B.n715 VSUBS 0.005816f
C769 B.n716 VSUBS 0.005816f
C770 B.n717 VSUBS 0.005816f
C771 B.n718 VSUBS 0.005816f
C772 B.n719 VSUBS 0.005816f
C773 B.n720 VSUBS 0.005816f
C774 B.n721 VSUBS 0.005816f
C775 B.n722 VSUBS 0.005816f
C776 B.n723 VSUBS 0.005816f
C777 B.n724 VSUBS 0.005816f
C778 B.n725 VSUBS 0.005816f
C779 B.n726 VSUBS 0.005816f
C780 B.n727 VSUBS 0.005816f
C781 B.n728 VSUBS 0.005816f
C782 B.n729 VSUBS 0.005816f
C783 B.n730 VSUBS 0.005816f
C784 B.n731 VSUBS 0.005816f
C785 B.n732 VSUBS 0.005816f
C786 B.n733 VSUBS 0.005816f
C787 B.n734 VSUBS 0.005816f
C788 B.n735 VSUBS 0.005816f
C789 B.n736 VSUBS 0.005816f
C790 B.n737 VSUBS 0.005816f
C791 B.n738 VSUBS 0.005816f
C792 B.n739 VSUBS 0.005816f
C793 B.n740 VSUBS 0.005816f
C794 B.n741 VSUBS 0.005816f
C795 B.n742 VSUBS 0.005816f
C796 B.n743 VSUBS 0.005816f
C797 B.n744 VSUBS 0.005816f
C798 B.n745 VSUBS 0.005816f
C799 B.n746 VSUBS 0.005816f
C800 B.n747 VSUBS 0.005816f
C801 B.n748 VSUBS 0.005816f
C802 B.n749 VSUBS 0.005816f
C803 B.n750 VSUBS 0.005816f
C804 B.n751 VSUBS 0.005816f
C805 B.n752 VSUBS 0.005816f
C806 B.n753 VSUBS 0.005816f
C807 B.n754 VSUBS 0.005816f
C808 B.n755 VSUBS 0.005816f
C809 B.n756 VSUBS 0.005816f
C810 B.n757 VSUBS 0.005816f
C811 B.n758 VSUBS 0.005816f
C812 B.n759 VSUBS 0.005816f
C813 B.n760 VSUBS 0.005816f
C814 B.n761 VSUBS 0.005816f
C815 B.n762 VSUBS 0.005816f
C816 B.n763 VSUBS 0.005816f
C817 B.n764 VSUBS 0.005816f
C818 B.n765 VSUBS 0.005816f
C819 B.n766 VSUBS 0.005816f
C820 B.n767 VSUBS 0.005816f
C821 B.n768 VSUBS 0.005816f
C822 B.n769 VSUBS 0.005816f
C823 B.n770 VSUBS 0.005816f
C824 B.n771 VSUBS 0.005816f
C825 B.n772 VSUBS 0.005816f
C826 B.n773 VSUBS 0.005816f
C827 B.n774 VSUBS 0.005816f
C828 B.n775 VSUBS 0.005816f
C829 B.n776 VSUBS 0.005816f
C830 B.n777 VSUBS 0.005816f
C831 B.n778 VSUBS 0.005816f
C832 B.n779 VSUBS 0.005816f
C833 B.n780 VSUBS 0.005816f
C834 B.n781 VSUBS 0.005816f
C835 B.n782 VSUBS 0.005816f
C836 B.n783 VSUBS 0.005816f
C837 B.n784 VSUBS 0.005816f
C838 B.n785 VSUBS 0.005816f
C839 B.n786 VSUBS 0.005816f
C840 B.n787 VSUBS 0.014272f
C841 B.n788 VSUBS 0.01361f
C842 B.n789 VSUBS 0.01361f
C843 B.n790 VSUBS 0.005816f
C844 B.n791 VSUBS 0.005816f
C845 B.n792 VSUBS 0.005816f
C846 B.n793 VSUBS 0.005816f
C847 B.n794 VSUBS 0.005816f
C848 B.n795 VSUBS 0.005816f
C849 B.n796 VSUBS 0.005816f
C850 B.n797 VSUBS 0.005816f
C851 B.n798 VSUBS 0.005816f
C852 B.n799 VSUBS 0.005816f
C853 B.n800 VSUBS 0.005816f
C854 B.n801 VSUBS 0.005816f
C855 B.n802 VSUBS 0.005816f
C856 B.n803 VSUBS 0.005816f
C857 B.n804 VSUBS 0.005816f
C858 B.n805 VSUBS 0.005816f
C859 B.n806 VSUBS 0.005816f
C860 B.n807 VSUBS 0.005816f
C861 B.n808 VSUBS 0.005816f
C862 B.n809 VSUBS 0.005816f
C863 B.n810 VSUBS 0.005816f
C864 B.n811 VSUBS 0.005816f
C865 B.n812 VSUBS 0.005816f
C866 B.n813 VSUBS 0.005816f
C867 B.n814 VSUBS 0.005816f
C868 B.n815 VSUBS 0.005816f
C869 B.n816 VSUBS 0.005816f
C870 B.n817 VSUBS 0.005816f
C871 B.n818 VSUBS 0.005816f
C872 B.n819 VSUBS 0.005816f
C873 B.n820 VSUBS 0.005816f
C874 B.n821 VSUBS 0.005816f
C875 B.n822 VSUBS 0.005816f
C876 B.n823 VSUBS 0.005816f
C877 B.n824 VSUBS 0.005816f
C878 B.n825 VSUBS 0.005816f
C879 B.n826 VSUBS 0.005816f
C880 B.n827 VSUBS 0.005816f
C881 B.n828 VSUBS 0.005816f
C882 B.n829 VSUBS 0.005816f
C883 B.n830 VSUBS 0.005816f
C884 B.n831 VSUBS 0.005816f
C885 B.n832 VSUBS 0.005816f
C886 B.n833 VSUBS 0.005816f
C887 B.n834 VSUBS 0.005816f
C888 B.n835 VSUBS 0.005816f
C889 B.n836 VSUBS 0.005816f
C890 B.n837 VSUBS 0.005816f
C891 B.n838 VSUBS 0.005816f
C892 B.n839 VSUBS 0.005816f
C893 B.n840 VSUBS 0.005816f
C894 B.n841 VSUBS 0.005816f
C895 B.n842 VSUBS 0.005816f
C896 B.n843 VSUBS 0.013169f
C897 VDD1.t0 VSUBS 0.404697f
C898 VDD1.t3 VSUBS 0.404697f
C899 VDD1.n0 VSUBS 3.41681f
C900 VDD1.t1 VSUBS 0.404697f
C901 VDD1.t2 VSUBS 0.404697f
C902 VDD1.n1 VSUBS 4.42549f
C903 VTAIL.t3 VSUBS 3.53871f
C904 VTAIL.n0 VSUBS 0.744345f
C905 VTAIL.t4 VSUBS 3.53871f
C906 VTAIL.n1 VSUBS 0.83792f
C907 VTAIL.t7 VSUBS 3.53871f
C908 VTAIL.n2 VSUBS 2.48466f
C909 VTAIL.t0 VSUBS 3.53874f
C910 VTAIL.n3 VSUBS 2.48463f
C911 VTAIL.t1 VSUBS 3.53874f
C912 VTAIL.n4 VSUBS 0.837888f
C913 VTAIL.t6 VSUBS 3.53874f
C914 VTAIL.n5 VSUBS 0.837888f
C915 VTAIL.t5 VSUBS 3.53871f
C916 VTAIL.n6 VSUBS 2.48466f
C917 VTAIL.t2 VSUBS 3.53871f
C918 VTAIL.n7 VSUBS 2.38276f
C919 VP.n0 VSUBS 0.037605f
C920 VP.t1 VSUBS 4.28081f
C921 VP.n1 VSUBS 0.05669f
C922 VP.n2 VSUBS 0.028523f
C923 VP.n3 VSUBS 0.031375f
C924 VP.t0 VSUBS 4.5724f
C925 VP.t3 VSUBS 4.57978f
C926 VP.n4 VSUBS 4.7706f
C927 VP.t2 VSUBS 4.28081f
C928 VP.n5 VSUBS 1.574f
C929 VP.n6 VSUBS 1.8543f
C930 VP.n7 VSUBS 0.037605f
C931 VP.n8 VSUBS 0.028523f
C932 VP.n9 VSUBS 0.05316f
C933 VP.n10 VSUBS 0.05669f
C934 VP.n11 VSUBS 0.023059f
C935 VP.n12 VSUBS 0.028523f
C936 VP.n13 VSUBS 0.028523f
C937 VP.n14 VSUBS 0.028523f
C938 VP.n15 VSUBS 0.05316f
C939 VP.n16 VSUBS 0.031375f
C940 VP.n17 VSUBS 1.574f
C941 VP.n18 VSUBS 0.052851f
.ends

