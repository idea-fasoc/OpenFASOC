* NGSPICE file created from diff_pair_sample_1664.ext - technology: sky130A

.subckt diff_pair_sample_1664 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=2.244 ps=13.93 w=13.6 l=3.33
X1 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=5.304 ps=27.98 w=13.6 l=3.33
X2 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=5.304 ps=27.98 w=13.6 l=3.33
X3 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=0 ps=0 w=13.6 l=3.33
X4 VTAIL.t3 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=2.244 ps=13.93 w=13.6 l=3.33
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=0 ps=0 w=13.6 l=3.33
X6 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=2.244 ps=13.93 w=13.6 l=3.33
X7 VDD1.t1 VP.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=2.244 ps=13.93 w=13.6 l=3.33
X8 VDD2.t0 VN.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=5.304 ps=27.98 w=13.6 l=3.33
X9 VDD2.t2 VN.t2 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=5.304 ps=27.98 w=13.6 l=3.33
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=0 ps=0 w=13.6 l=3.33
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=0 ps=0 w=13.6 l=3.33
X12 VTAIL.t5 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=2.244 ps=13.93 w=13.6 l=3.33
X13 VDD2.t5 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=2.244 ps=13.93 w=13.6 l=3.33
X14 VDD2.t1 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=5.304 pd=27.98 as=2.244 ps=13.93 w=13.6 l=3.33
X15 VTAIL.t6 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.244 pd=13.93 as=2.244 ps=13.93 w=13.6 l=3.33
R0 VN.n34 VN.n33 161.3
R1 VN.n32 VN.n19 161.3
R2 VN.n31 VN.n30 161.3
R3 VN.n29 VN.n20 161.3
R4 VN.n28 VN.n27 161.3
R5 VN.n26 VN.n21 161.3
R6 VN.n25 VN.n24 161.3
R7 VN.n16 VN.n15 161.3
R8 VN.n14 VN.n1 161.3
R9 VN.n13 VN.n12 161.3
R10 VN.n11 VN.n2 161.3
R11 VN.n10 VN.n9 161.3
R12 VN.n8 VN.n3 161.3
R13 VN.n7 VN.n6 161.3
R14 VN.n23 VN.t1 131.531
R15 VN.n5 VN.t4 131.531
R16 VN.n4 VN.t5 98.4269
R17 VN.n0 VN.t2 98.4269
R18 VN.n22 VN.t0 98.4269
R19 VN.n18 VN.t3 98.4269
R20 VN.n17 VN.n0 82.3762
R21 VN.n35 VN.n18 82.3762
R22 VN.n9 VN.n2 56.5617
R23 VN.n27 VN.n20 56.5617
R24 VN VN.n35 52.93
R25 VN.n5 VN.n4 50.1747
R26 VN.n23 VN.n22 50.1747
R27 VN.n7 VN.n4 24.5923
R28 VN.n8 VN.n7 24.5923
R29 VN.n9 VN.n8 24.5923
R30 VN.n13 VN.n2 24.5923
R31 VN.n14 VN.n13 24.5923
R32 VN.n15 VN.n14 24.5923
R33 VN.n27 VN.n26 24.5923
R34 VN.n26 VN.n25 24.5923
R35 VN.n25 VN.n22 24.5923
R36 VN.n33 VN.n32 24.5923
R37 VN.n32 VN.n31 24.5923
R38 VN.n31 VN.n20 24.5923
R39 VN.n15 VN.n0 7.86989
R40 VN.n33 VN.n18 7.86989
R41 VN.n6 VN.n5 3.21487
R42 VN.n24 VN.n23 3.21487
R43 VN.n35 VN.n34 0.354861
R44 VN.n17 VN.n16 0.354861
R45 VN VN.n17 0.267071
R46 VN.n34 VN.n19 0.189894
R47 VN.n30 VN.n19 0.189894
R48 VN.n30 VN.n29 0.189894
R49 VN.n29 VN.n28 0.189894
R50 VN.n28 VN.n21 0.189894
R51 VN.n24 VN.n21 0.189894
R52 VN.n6 VN.n3 0.189894
R53 VN.n10 VN.n3 0.189894
R54 VN.n11 VN.n10 0.189894
R55 VN.n12 VN.n11 0.189894
R56 VN.n12 VN.n1 0.189894
R57 VN.n16 VN.n1 0.189894
R58 VDD2.n143 VDD2.n75 289.615
R59 VDD2.n68 VDD2.n0 289.615
R60 VDD2.n144 VDD2.n143 185
R61 VDD2.n142 VDD2.n141 185
R62 VDD2.n79 VDD2.n78 185
R63 VDD2.n136 VDD2.n135 185
R64 VDD2.n134 VDD2.n133 185
R65 VDD2.n83 VDD2.n82 185
R66 VDD2.n128 VDD2.n127 185
R67 VDD2.n126 VDD2.n125 185
R68 VDD2.n87 VDD2.n86 185
R69 VDD2.n91 VDD2.n89 185
R70 VDD2.n120 VDD2.n119 185
R71 VDD2.n118 VDD2.n117 185
R72 VDD2.n93 VDD2.n92 185
R73 VDD2.n112 VDD2.n111 185
R74 VDD2.n110 VDD2.n109 185
R75 VDD2.n97 VDD2.n96 185
R76 VDD2.n104 VDD2.n103 185
R77 VDD2.n102 VDD2.n101 185
R78 VDD2.n25 VDD2.n24 185
R79 VDD2.n27 VDD2.n26 185
R80 VDD2.n20 VDD2.n19 185
R81 VDD2.n33 VDD2.n32 185
R82 VDD2.n35 VDD2.n34 185
R83 VDD2.n16 VDD2.n15 185
R84 VDD2.n42 VDD2.n41 185
R85 VDD2.n43 VDD2.n14 185
R86 VDD2.n45 VDD2.n44 185
R87 VDD2.n12 VDD2.n11 185
R88 VDD2.n51 VDD2.n50 185
R89 VDD2.n53 VDD2.n52 185
R90 VDD2.n8 VDD2.n7 185
R91 VDD2.n59 VDD2.n58 185
R92 VDD2.n61 VDD2.n60 185
R93 VDD2.n4 VDD2.n3 185
R94 VDD2.n67 VDD2.n66 185
R95 VDD2.n69 VDD2.n68 185
R96 VDD2.n100 VDD2.t5 149.524
R97 VDD2.n23 VDD2.t1 149.524
R98 VDD2.n143 VDD2.n142 104.615
R99 VDD2.n142 VDD2.n78 104.615
R100 VDD2.n135 VDD2.n78 104.615
R101 VDD2.n135 VDD2.n134 104.615
R102 VDD2.n134 VDD2.n82 104.615
R103 VDD2.n127 VDD2.n82 104.615
R104 VDD2.n127 VDD2.n126 104.615
R105 VDD2.n126 VDD2.n86 104.615
R106 VDD2.n91 VDD2.n86 104.615
R107 VDD2.n119 VDD2.n91 104.615
R108 VDD2.n119 VDD2.n118 104.615
R109 VDD2.n118 VDD2.n92 104.615
R110 VDD2.n111 VDD2.n92 104.615
R111 VDD2.n111 VDD2.n110 104.615
R112 VDD2.n110 VDD2.n96 104.615
R113 VDD2.n103 VDD2.n96 104.615
R114 VDD2.n103 VDD2.n102 104.615
R115 VDD2.n26 VDD2.n25 104.615
R116 VDD2.n26 VDD2.n19 104.615
R117 VDD2.n33 VDD2.n19 104.615
R118 VDD2.n34 VDD2.n33 104.615
R119 VDD2.n34 VDD2.n15 104.615
R120 VDD2.n42 VDD2.n15 104.615
R121 VDD2.n43 VDD2.n42 104.615
R122 VDD2.n44 VDD2.n43 104.615
R123 VDD2.n44 VDD2.n11 104.615
R124 VDD2.n51 VDD2.n11 104.615
R125 VDD2.n52 VDD2.n51 104.615
R126 VDD2.n52 VDD2.n7 104.615
R127 VDD2.n59 VDD2.n7 104.615
R128 VDD2.n60 VDD2.n59 104.615
R129 VDD2.n60 VDD2.n3 104.615
R130 VDD2.n67 VDD2.n3 104.615
R131 VDD2.n68 VDD2.n67 104.615
R132 VDD2.n74 VDD2.n73 63.0632
R133 VDD2 VDD2.n149 63.0604
R134 VDD2.n102 VDD2.t5 52.3082
R135 VDD2.n25 VDD2.t1 52.3082
R136 VDD2.n74 VDD2.n72 51.9509
R137 VDD2.n148 VDD2.n147 49.6399
R138 VDD2.n148 VDD2.n74 45.6937
R139 VDD2.n89 VDD2.n87 13.1884
R140 VDD2.n45 VDD2.n12 13.1884
R141 VDD2.n125 VDD2.n124 12.8005
R142 VDD2.n121 VDD2.n120 12.8005
R143 VDD2.n46 VDD2.n14 12.8005
R144 VDD2.n50 VDD2.n49 12.8005
R145 VDD2.n128 VDD2.n85 12.0247
R146 VDD2.n117 VDD2.n90 12.0247
R147 VDD2.n41 VDD2.n40 12.0247
R148 VDD2.n53 VDD2.n10 12.0247
R149 VDD2.n129 VDD2.n83 11.249
R150 VDD2.n116 VDD2.n93 11.249
R151 VDD2.n39 VDD2.n16 11.249
R152 VDD2.n54 VDD2.n8 11.249
R153 VDD2.n133 VDD2.n132 10.4732
R154 VDD2.n113 VDD2.n112 10.4732
R155 VDD2.n36 VDD2.n35 10.4732
R156 VDD2.n58 VDD2.n57 10.4732
R157 VDD2.n101 VDD2.n100 10.2747
R158 VDD2.n24 VDD2.n23 10.2747
R159 VDD2.n136 VDD2.n81 9.69747
R160 VDD2.n109 VDD2.n95 9.69747
R161 VDD2.n32 VDD2.n18 9.69747
R162 VDD2.n61 VDD2.n6 9.69747
R163 VDD2.n147 VDD2.n146 9.45567
R164 VDD2.n72 VDD2.n71 9.45567
R165 VDD2.n99 VDD2.n98 9.3005
R166 VDD2.n106 VDD2.n105 9.3005
R167 VDD2.n108 VDD2.n107 9.3005
R168 VDD2.n95 VDD2.n94 9.3005
R169 VDD2.n114 VDD2.n113 9.3005
R170 VDD2.n116 VDD2.n115 9.3005
R171 VDD2.n90 VDD2.n88 9.3005
R172 VDD2.n122 VDD2.n121 9.3005
R173 VDD2.n146 VDD2.n145 9.3005
R174 VDD2.n77 VDD2.n76 9.3005
R175 VDD2.n140 VDD2.n139 9.3005
R176 VDD2.n138 VDD2.n137 9.3005
R177 VDD2.n81 VDD2.n80 9.3005
R178 VDD2.n132 VDD2.n131 9.3005
R179 VDD2.n130 VDD2.n129 9.3005
R180 VDD2.n85 VDD2.n84 9.3005
R181 VDD2.n124 VDD2.n123 9.3005
R182 VDD2.n71 VDD2.n70 9.3005
R183 VDD2.n65 VDD2.n64 9.3005
R184 VDD2.n63 VDD2.n62 9.3005
R185 VDD2.n6 VDD2.n5 9.3005
R186 VDD2.n57 VDD2.n56 9.3005
R187 VDD2.n55 VDD2.n54 9.3005
R188 VDD2.n10 VDD2.n9 9.3005
R189 VDD2.n49 VDD2.n48 9.3005
R190 VDD2.n22 VDD2.n21 9.3005
R191 VDD2.n29 VDD2.n28 9.3005
R192 VDD2.n31 VDD2.n30 9.3005
R193 VDD2.n18 VDD2.n17 9.3005
R194 VDD2.n37 VDD2.n36 9.3005
R195 VDD2.n39 VDD2.n38 9.3005
R196 VDD2.n40 VDD2.n13 9.3005
R197 VDD2.n47 VDD2.n46 9.3005
R198 VDD2.n2 VDD2.n1 9.3005
R199 VDD2.n137 VDD2.n79 8.92171
R200 VDD2.n108 VDD2.n97 8.92171
R201 VDD2.n31 VDD2.n20 8.92171
R202 VDD2.n62 VDD2.n4 8.92171
R203 VDD2.n141 VDD2.n140 8.14595
R204 VDD2.n105 VDD2.n104 8.14595
R205 VDD2.n28 VDD2.n27 8.14595
R206 VDD2.n66 VDD2.n65 8.14595
R207 VDD2.n147 VDD2.n75 7.3702
R208 VDD2.n144 VDD2.n77 7.3702
R209 VDD2.n101 VDD2.n99 7.3702
R210 VDD2.n24 VDD2.n22 7.3702
R211 VDD2.n69 VDD2.n2 7.3702
R212 VDD2.n72 VDD2.n0 7.3702
R213 VDD2.n145 VDD2.n75 6.59444
R214 VDD2.n145 VDD2.n144 6.59444
R215 VDD2.n70 VDD2.n69 6.59444
R216 VDD2.n70 VDD2.n0 6.59444
R217 VDD2.n141 VDD2.n77 5.81868
R218 VDD2.n104 VDD2.n99 5.81868
R219 VDD2.n27 VDD2.n22 5.81868
R220 VDD2.n66 VDD2.n2 5.81868
R221 VDD2.n140 VDD2.n79 5.04292
R222 VDD2.n105 VDD2.n97 5.04292
R223 VDD2.n28 VDD2.n20 5.04292
R224 VDD2.n65 VDD2.n4 5.04292
R225 VDD2.n137 VDD2.n136 4.26717
R226 VDD2.n109 VDD2.n108 4.26717
R227 VDD2.n32 VDD2.n31 4.26717
R228 VDD2.n62 VDD2.n61 4.26717
R229 VDD2.n133 VDD2.n81 3.49141
R230 VDD2.n112 VDD2.n95 3.49141
R231 VDD2.n35 VDD2.n18 3.49141
R232 VDD2.n58 VDD2.n6 3.49141
R233 VDD2.n100 VDD2.n98 2.84303
R234 VDD2.n23 VDD2.n21 2.84303
R235 VDD2.n132 VDD2.n83 2.71565
R236 VDD2.n113 VDD2.n93 2.71565
R237 VDD2.n36 VDD2.n16 2.71565
R238 VDD2.n57 VDD2.n8 2.71565
R239 VDD2 VDD2.n148 2.42507
R240 VDD2.n129 VDD2.n128 1.93989
R241 VDD2.n117 VDD2.n116 1.93989
R242 VDD2.n41 VDD2.n39 1.93989
R243 VDD2.n54 VDD2.n53 1.93989
R244 VDD2.n149 VDD2.t3 1.45638
R245 VDD2.n149 VDD2.t0 1.45638
R246 VDD2.n73 VDD2.t4 1.45638
R247 VDD2.n73 VDD2.t2 1.45638
R248 VDD2.n125 VDD2.n85 1.16414
R249 VDD2.n120 VDD2.n90 1.16414
R250 VDD2.n40 VDD2.n14 1.16414
R251 VDD2.n50 VDD2.n10 1.16414
R252 VDD2.n124 VDD2.n87 0.388379
R253 VDD2.n121 VDD2.n89 0.388379
R254 VDD2.n46 VDD2.n45 0.388379
R255 VDD2.n49 VDD2.n12 0.388379
R256 VDD2.n146 VDD2.n76 0.155672
R257 VDD2.n139 VDD2.n76 0.155672
R258 VDD2.n139 VDD2.n138 0.155672
R259 VDD2.n138 VDD2.n80 0.155672
R260 VDD2.n131 VDD2.n80 0.155672
R261 VDD2.n131 VDD2.n130 0.155672
R262 VDD2.n130 VDD2.n84 0.155672
R263 VDD2.n123 VDD2.n84 0.155672
R264 VDD2.n123 VDD2.n122 0.155672
R265 VDD2.n122 VDD2.n88 0.155672
R266 VDD2.n115 VDD2.n88 0.155672
R267 VDD2.n115 VDD2.n114 0.155672
R268 VDD2.n114 VDD2.n94 0.155672
R269 VDD2.n107 VDD2.n94 0.155672
R270 VDD2.n107 VDD2.n106 0.155672
R271 VDD2.n106 VDD2.n98 0.155672
R272 VDD2.n29 VDD2.n21 0.155672
R273 VDD2.n30 VDD2.n29 0.155672
R274 VDD2.n30 VDD2.n17 0.155672
R275 VDD2.n37 VDD2.n17 0.155672
R276 VDD2.n38 VDD2.n37 0.155672
R277 VDD2.n38 VDD2.n13 0.155672
R278 VDD2.n47 VDD2.n13 0.155672
R279 VDD2.n48 VDD2.n47 0.155672
R280 VDD2.n48 VDD2.n9 0.155672
R281 VDD2.n55 VDD2.n9 0.155672
R282 VDD2.n56 VDD2.n55 0.155672
R283 VDD2.n56 VDD2.n5 0.155672
R284 VDD2.n63 VDD2.n5 0.155672
R285 VDD2.n64 VDD2.n63 0.155672
R286 VDD2.n64 VDD2.n1 0.155672
R287 VDD2.n71 VDD2.n1 0.155672
R288 VTAIL.n298 VTAIL.n230 289.615
R289 VTAIL.n70 VTAIL.n2 289.615
R290 VTAIL.n224 VTAIL.n156 289.615
R291 VTAIL.n148 VTAIL.n80 289.615
R292 VTAIL.n255 VTAIL.n254 185
R293 VTAIL.n257 VTAIL.n256 185
R294 VTAIL.n250 VTAIL.n249 185
R295 VTAIL.n263 VTAIL.n262 185
R296 VTAIL.n265 VTAIL.n264 185
R297 VTAIL.n246 VTAIL.n245 185
R298 VTAIL.n272 VTAIL.n271 185
R299 VTAIL.n273 VTAIL.n244 185
R300 VTAIL.n275 VTAIL.n274 185
R301 VTAIL.n242 VTAIL.n241 185
R302 VTAIL.n281 VTAIL.n280 185
R303 VTAIL.n283 VTAIL.n282 185
R304 VTAIL.n238 VTAIL.n237 185
R305 VTAIL.n289 VTAIL.n288 185
R306 VTAIL.n291 VTAIL.n290 185
R307 VTAIL.n234 VTAIL.n233 185
R308 VTAIL.n297 VTAIL.n296 185
R309 VTAIL.n299 VTAIL.n298 185
R310 VTAIL.n27 VTAIL.n26 185
R311 VTAIL.n29 VTAIL.n28 185
R312 VTAIL.n22 VTAIL.n21 185
R313 VTAIL.n35 VTAIL.n34 185
R314 VTAIL.n37 VTAIL.n36 185
R315 VTAIL.n18 VTAIL.n17 185
R316 VTAIL.n44 VTAIL.n43 185
R317 VTAIL.n45 VTAIL.n16 185
R318 VTAIL.n47 VTAIL.n46 185
R319 VTAIL.n14 VTAIL.n13 185
R320 VTAIL.n53 VTAIL.n52 185
R321 VTAIL.n55 VTAIL.n54 185
R322 VTAIL.n10 VTAIL.n9 185
R323 VTAIL.n61 VTAIL.n60 185
R324 VTAIL.n63 VTAIL.n62 185
R325 VTAIL.n6 VTAIL.n5 185
R326 VTAIL.n69 VTAIL.n68 185
R327 VTAIL.n71 VTAIL.n70 185
R328 VTAIL.n225 VTAIL.n224 185
R329 VTAIL.n223 VTAIL.n222 185
R330 VTAIL.n160 VTAIL.n159 185
R331 VTAIL.n217 VTAIL.n216 185
R332 VTAIL.n215 VTAIL.n214 185
R333 VTAIL.n164 VTAIL.n163 185
R334 VTAIL.n209 VTAIL.n208 185
R335 VTAIL.n207 VTAIL.n206 185
R336 VTAIL.n168 VTAIL.n167 185
R337 VTAIL.n172 VTAIL.n170 185
R338 VTAIL.n201 VTAIL.n200 185
R339 VTAIL.n199 VTAIL.n198 185
R340 VTAIL.n174 VTAIL.n173 185
R341 VTAIL.n193 VTAIL.n192 185
R342 VTAIL.n191 VTAIL.n190 185
R343 VTAIL.n178 VTAIL.n177 185
R344 VTAIL.n185 VTAIL.n184 185
R345 VTAIL.n183 VTAIL.n182 185
R346 VTAIL.n149 VTAIL.n148 185
R347 VTAIL.n147 VTAIL.n146 185
R348 VTAIL.n84 VTAIL.n83 185
R349 VTAIL.n141 VTAIL.n140 185
R350 VTAIL.n139 VTAIL.n138 185
R351 VTAIL.n88 VTAIL.n87 185
R352 VTAIL.n133 VTAIL.n132 185
R353 VTAIL.n131 VTAIL.n130 185
R354 VTAIL.n92 VTAIL.n91 185
R355 VTAIL.n96 VTAIL.n94 185
R356 VTAIL.n125 VTAIL.n124 185
R357 VTAIL.n123 VTAIL.n122 185
R358 VTAIL.n98 VTAIL.n97 185
R359 VTAIL.n117 VTAIL.n116 185
R360 VTAIL.n115 VTAIL.n114 185
R361 VTAIL.n102 VTAIL.n101 185
R362 VTAIL.n109 VTAIL.n108 185
R363 VTAIL.n107 VTAIL.n106 185
R364 VTAIL.n253 VTAIL.t9 149.524
R365 VTAIL.n25 VTAIL.t0 149.524
R366 VTAIL.n181 VTAIL.t2 149.524
R367 VTAIL.n105 VTAIL.t10 149.524
R368 VTAIL.n256 VTAIL.n255 104.615
R369 VTAIL.n256 VTAIL.n249 104.615
R370 VTAIL.n263 VTAIL.n249 104.615
R371 VTAIL.n264 VTAIL.n263 104.615
R372 VTAIL.n264 VTAIL.n245 104.615
R373 VTAIL.n272 VTAIL.n245 104.615
R374 VTAIL.n273 VTAIL.n272 104.615
R375 VTAIL.n274 VTAIL.n273 104.615
R376 VTAIL.n274 VTAIL.n241 104.615
R377 VTAIL.n281 VTAIL.n241 104.615
R378 VTAIL.n282 VTAIL.n281 104.615
R379 VTAIL.n282 VTAIL.n237 104.615
R380 VTAIL.n289 VTAIL.n237 104.615
R381 VTAIL.n290 VTAIL.n289 104.615
R382 VTAIL.n290 VTAIL.n233 104.615
R383 VTAIL.n297 VTAIL.n233 104.615
R384 VTAIL.n298 VTAIL.n297 104.615
R385 VTAIL.n28 VTAIL.n27 104.615
R386 VTAIL.n28 VTAIL.n21 104.615
R387 VTAIL.n35 VTAIL.n21 104.615
R388 VTAIL.n36 VTAIL.n35 104.615
R389 VTAIL.n36 VTAIL.n17 104.615
R390 VTAIL.n44 VTAIL.n17 104.615
R391 VTAIL.n45 VTAIL.n44 104.615
R392 VTAIL.n46 VTAIL.n45 104.615
R393 VTAIL.n46 VTAIL.n13 104.615
R394 VTAIL.n53 VTAIL.n13 104.615
R395 VTAIL.n54 VTAIL.n53 104.615
R396 VTAIL.n54 VTAIL.n9 104.615
R397 VTAIL.n61 VTAIL.n9 104.615
R398 VTAIL.n62 VTAIL.n61 104.615
R399 VTAIL.n62 VTAIL.n5 104.615
R400 VTAIL.n69 VTAIL.n5 104.615
R401 VTAIL.n70 VTAIL.n69 104.615
R402 VTAIL.n224 VTAIL.n223 104.615
R403 VTAIL.n223 VTAIL.n159 104.615
R404 VTAIL.n216 VTAIL.n159 104.615
R405 VTAIL.n216 VTAIL.n215 104.615
R406 VTAIL.n215 VTAIL.n163 104.615
R407 VTAIL.n208 VTAIL.n163 104.615
R408 VTAIL.n208 VTAIL.n207 104.615
R409 VTAIL.n207 VTAIL.n167 104.615
R410 VTAIL.n172 VTAIL.n167 104.615
R411 VTAIL.n200 VTAIL.n172 104.615
R412 VTAIL.n200 VTAIL.n199 104.615
R413 VTAIL.n199 VTAIL.n173 104.615
R414 VTAIL.n192 VTAIL.n173 104.615
R415 VTAIL.n192 VTAIL.n191 104.615
R416 VTAIL.n191 VTAIL.n177 104.615
R417 VTAIL.n184 VTAIL.n177 104.615
R418 VTAIL.n184 VTAIL.n183 104.615
R419 VTAIL.n148 VTAIL.n147 104.615
R420 VTAIL.n147 VTAIL.n83 104.615
R421 VTAIL.n140 VTAIL.n83 104.615
R422 VTAIL.n140 VTAIL.n139 104.615
R423 VTAIL.n139 VTAIL.n87 104.615
R424 VTAIL.n132 VTAIL.n87 104.615
R425 VTAIL.n132 VTAIL.n131 104.615
R426 VTAIL.n131 VTAIL.n91 104.615
R427 VTAIL.n96 VTAIL.n91 104.615
R428 VTAIL.n124 VTAIL.n96 104.615
R429 VTAIL.n124 VTAIL.n123 104.615
R430 VTAIL.n123 VTAIL.n97 104.615
R431 VTAIL.n116 VTAIL.n97 104.615
R432 VTAIL.n116 VTAIL.n115 104.615
R433 VTAIL.n115 VTAIL.n101 104.615
R434 VTAIL.n108 VTAIL.n101 104.615
R435 VTAIL.n108 VTAIL.n107 104.615
R436 VTAIL.n255 VTAIL.t9 52.3082
R437 VTAIL.n27 VTAIL.t0 52.3082
R438 VTAIL.n183 VTAIL.t2 52.3082
R439 VTAIL.n107 VTAIL.t10 52.3082
R440 VTAIL.n155 VTAIL.n154 45.6511
R441 VTAIL.n79 VTAIL.n78 45.6511
R442 VTAIL.n1 VTAIL.n0 45.651
R443 VTAIL.n77 VTAIL.n76 45.651
R444 VTAIL.n303 VTAIL.n302 32.9611
R445 VTAIL.n75 VTAIL.n74 32.9611
R446 VTAIL.n229 VTAIL.n228 32.9611
R447 VTAIL.n153 VTAIL.n152 32.9611
R448 VTAIL.n79 VTAIL.n77 30.4014
R449 VTAIL.n303 VTAIL.n229 27.2462
R450 VTAIL.n275 VTAIL.n242 13.1884
R451 VTAIL.n47 VTAIL.n14 13.1884
R452 VTAIL.n170 VTAIL.n168 13.1884
R453 VTAIL.n94 VTAIL.n92 13.1884
R454 VTAIL.n276 VTAIL.n244 12.8005
R455 VTAIL.n280 VTAIL.n279 12.8005
R456 VTAIL.n48 VTAIL.n16 12.8005
R457 VTAIL.n52 VTAIL.n51 12.8005
R458 VTAIL.n206 VTAIL.n205 12.8005
R459 VTAIL.n202 VTAIL.n201 12.8005
R460 VTAIL.n130 VTAIL.n129 12.8005
R461 VTAIL.n126 VTAIL.n125 12.8005
R462 VTAIL.n271 VTAIL.n270 12.0247
R463 VTAIL.n283 VTAIL.n240 12.0247
R464 VTAIL.n43 VTAIL.n42 12.0247
R465 VTAIL.n55 VTAIL.n12 12.0247
R466 VTAIL.n209 VTAIL.n166 12.0247
R467 VTAIL.n198 VTAIL.n171 12.0247
R468 VTAIL.n133 VTAIL.n90 12.0247
R469 VTAIL.n122 VTAIL.n95 12.0247
R470 VTAIL.n269 VTAIL.n246 11.249
R471 VTAIL.n284 VTAIL.n238 11.249
R472 VTAIL.n41 VTAIL.n18 11.249
R473 VTAIL.n56 VTAIL.n10 11.249
R474 VTAIL.n210 VTAIL.n164 11.249
R475 VTAIL.n197 VTAIL.n174 11.249
R476 VTAIL.n134 VTAIL.n88 11.249
R477 VTAIL.n121 VTAIL.n98 11.249
R478 VTAIL.n266 VTAIL.n265 10.4732
R479 VTAIL.n288 VTAIL.n287 10.4732
R480 VTAIL.n38 VTAIL.n37 10.4732
R481 VTAIL.n60 VTAIL.n59 10.4732
R482 VTAIL.n214 VTAIL.n213 10.4732
R483 VTAIL.n194 VTAIL.n193 10.4732
R484 VTAIL.n138 VTAIL.n137 10.4732
R485 VTAIL.n118 VTAIL.n117 10.4732
R486 VTAIL.n254 VTAIL.n253 10.2747
R487 VTAIL.n26 VTAIL.n25 10.2747
R488 VTAIL.n182 VTAIL.n181 10.2747
R489 VTAIL.n106 VTAIL.n105 10.2747
R490 VTAIL.n262 VTAIL.n248 9.69747
R491 VTAIL.n291 VTAIL.n236 9.69747
R492 VTAIL.n34 VTAIL.n20 9.69747
R493 VTAIL.n63 VTAIL.n8 9.69747
R494 VTAIL.n217 VTAIL.n162 9.69747
R495 VTAIL.n190 VTAIL.n176 9.69747
R496 VTAIL.n141 VTAIL.n86 9.69747
R497 VTAIL.n114 VTAIL.n100 9.69747
R498 VTAIL.n302 VTAIL.n301 9.45567
R499 VTAIL.n74 VTAIL.n73 9.45567
R500 VTAIL.n228 VTAIL.n227 9.45567
R501 VTAIL.n152 VTAIL.n151 9.45567
R502 VTAIL.n301 VTAIL.n300 9.3005
R503 VTAIL.n295 VTAIL.n294 9.3005
R504 VTAIL.n293 VTAIL.n292 9.3005
R505 VTAIL.n236 VTAIL.n235 9.3005
R506 VTAIL.n287 VTAIL.n286 9.3005
R507 VTAIL.n285 VTAIL.n284 9.3005
R508 VTAIL.n240 VTAIL.n239 9.3005
R509 VTAIL.n279 VTAIL.n278 9.3005
R510 VTAIL.n252 VTAIL.n251 9.3005
R511 VTAIL.n259 VTAIL.n258 9.3005
R512 VTAIL.n261 VTAIL.n260 9.3005
R513 VTAIL.n248 VTAIL.n247 9.3005
R514 VTAIL.n267 VTAIL.n266 9.3005
R515 VTAIL.n269 VTAIL.n268 9.3005
R516 VTAIL.n270 VTAIL.n243 9.3005
R517 VTAIL.n277 VTAIL.n276 9.3005
R518 VTAIL.n232 VTAIL.n231 9.3005
R519 VTAIL.n73 VTAIL.n72 9.3005
R520 VTAIL.n67 VTAIL.n66 9.3005
R521 VTAIL.n65 VTAIL.n64 9.3005
R522 VTAIL.n8 VTAIL.n7 9.3005
R523 VTAIL.n59 VTAIL.n58 9.3005
R524 VTAIL.n57 VTAIL.n56 9.3005
R525 VTAIL.n12 VTAIL.n11 9.3005
R526 VTAIL.n51 VTAIL.n50 9.3005
R527 VTAIL.n24 VTAIL.n23 9.3005
R528 VTAIL.n31 VTAIL.n30 9.3005
R529 VTAIL.n33 VTAIL.n32 9.3005
R530 VTAIL.n20 VTAIL.n19 9.3005
R531 VTAIL.n39 VTAIL.n38 9.3005
R532 VTAIL.n41 VTAIL.n40 9.3005
R533 VTAIL.n42 VTAIL.n15 9.3005
R534 VTAIL.n49 VTAIL.n48 9.3005
R535 VTAIL.n4 VTAIL.n3 9.3005
R536 VTAIL.n180 VTAIL.n179 9.3005
R537 VTAIL.n187 VTAIL.n186 9.3005
R538 VTAIL.n189 VTAIL.n188 9.3005
R539 VTAIL.n176 VTAIL.n175 9.3005
R540 VTAIL.n195 VTAIL.n194 9.3005
R541 VTAIL.n197 VTAIL.n196 9.3005
R542 VTAIL.n171 VTAIL.n169 9.3005
R543 VTAIL.n203 VTAIL.n202 9.3005
R544 VTAIL.n227 VTAIL.n226 9.3005
R545 VTAIL.n158 VTAIL.n157 9.3005
R546 VTAIL.n221 VTAIL.n220 9.3005
R547 VTAIL.n219 VTAIL.n218 9.3005
R548 VTAIL.n162 VTAIL.n161 9.3005
R549 VTAIL.n213 VTAIL.n212 9.3005
R550 VTAIL.n211 VTAIL.n210 9.3005
R551 VTAIL.n166 VTAIL.n165 9.3005
R552 VTAIL.n205 VTAIL.n204 9.3005
R553 VTAIL.n104 VTAIL.n103 9.3005
R554 VTAIL.n111 VTAIL.n110 9.3005
R555 VTAIL.n113 VTAIL.n112 9.3005
R556 VTAIL.n100 VTAIL.n99 9.3005
R557 VTAIL.n119 VTAIL.n118 9.3005
R558 VTAIL.n121 VTAIL.n120 9.3005
R559 VTAIL.n95 VTAIL.n93 9.3005
R560 VTAIL.n127 VTAIL.n126 9.3005
R561 VTAIL.n151 VTAIL.n150 9.3005
R562 VTAIL.n82 VTAIL.n81 9.3005
R563 VTAIL.n145 VTAIL.n144 9.3005
R564 VTAIL.n143 VTAIL.n142 9.3005
R565 VTAIL.n86 VTAIL.n85 9.3005
R566 VTAIL.n137 VTAIL.n136 9.3005
R567 VTAIL.n135 VTAIL.n134 9.3005
R568 VTAIL.n90 VTAIL.n89 9.3005
R569 VTAIL.n129 VTAIL.n128 9.3005
R570 VTAIL.n261 VTAIL.n250 8.92171
R571 VTAIL.n292 VTAIL.n234 8.92171
R572 VTAIL.n33 VTAIL.n22 8.92171
R573 VTAIL.n64 VTAIL.n6 8.92171
R574 VTAIL.n218 VTAIL.n160 8.92171
R575 VTAIL.n189 VTAIL.n178 8.92171
R576 VTAIL.n142 VTAIL.n84 8.92171
R577 VTAIL.n113 VTAIL.n102 8.92171
R578 VTAIL.n258 VTAIL.n257 8.14595
R579 VTAIL.n296 VTAIL.n295 8.14595
R580 VTAIL.n30 VTAIL.n29 8.14595
R581 VTAIL.n68 VTAIL.n67 8.14595
R582 VTAIL.n222 VTAIL.n221 8.14595
R583 VTAIL.n186 VTAIL.n185 8.14595
R584 VTAIL.n146 VTAIL.n145 8.14595
R585 VTAIL.n110 VTAIL.n109 8.14595
R586 VTAIL.n254 VTAIL.n252 7.3702
R587 VTAIL.n299 VTAIL.n232 7.3702
R588 VTAIL.n302 VTAIL.n230 7.3702
R589 VTAIL.n26 VTAIL.n24 7.3702
R590 VTAIL.n71 VTAIL.n4 7.3702
R591 VTAIL.n74 VTAIL.n2 7.3702
R592 VTAIL.n228 VTAIL.n156 7.3702
R593 VTAIL.n225 VTAIL.n158 7.3702
R594 VTAIL.n182 VTAIL.n180 7.3702
R595 VTAIL.n152 VTAIL.n80 7.3702
R596 VTAIL.n149 VTAIL.n82 7.3702
R597 VTAIL.n106 VTAIL.n104 7.3702
R598 VTAIL.n300 VTAIL.n299 6.59444
R599 VTAIL.n300 VTAIL.n230 6.59444
R600 VTAIL.n72 VTAIL.n71 6.59444
R601 VTAIL.n72 VTAIL.n2 6.59444
R602 VTAIL.n226 VTAIL.n156 6.59444
R603 VTAIL.n226 VTAIL.n225 6.59444
R604 VTAIL.n150 VTAIL.n80 6.59444
R605 VTAIL.n150 VTAIL.n149 6.59444
R606 VTAIL.n257 VTAIL.n252 5.81868
R607 VTAIL.n296 VTAIL.n232 5.81868
R608 VTAIL.n29 VTAIL.n24 5.81868
R609 VTAIL.n68 VTAIL.n4 5.81868
R610 VTAIL.n222 VTAIL.n158 5.81868
R611 VTAIL.n185 VTAIL.n180 5.81868
R612 VTAIL.n146 VTAIL.n82 5.81868
R613 VTAIL.n109 VTAIL.n104 5.81868
R614 VTAIL.n258 VTAIL.n250 5.04292
R615 VTAIL.n295 VTAIL.n234 5.04292
R616 VTAIL.n30 VTAIL.n22 5.04292
R617 VTAIL.n67 VTAIL.n6 5.04292
R618 VTAIL.n221 VTAIL.n160 5.04292
R619 VTAIL.n186 VTAIL.n178 5.04292
R620 VTAIL.n145 VTAIL.n84 5.04292
R621 VTAIL.n110 VTAIL.n102 5.04292
R622 VTAIL.n262 VTAIL.n261 4.26717
R623 VTAIL.n292 VTAIL.n291 4.26717
R624 VTAIL.n34 VTAIL.n33 4.26717
R625 VTAIL.n64 VTAIL.n63 4.26717
R626 VTAIL.n218 VTAIL.n217 4.26717
R627 VTAIL.n190 VTAIL.n189 4.26717
R628 VTAIL.n142 VTAIL.n141 4.26717
R629 VTAIL.n114 VTAIL.n113 4.26717
R630 VTAIL.n265 VTAIL.n248 3.49141
R631 VTAIL.n288 VTAIL.n236 3.49141
R632 VTAIL.n37 VTAIL.n20 3.49141
R633 VTAIL.n60 VTAIL.n8 3.49141
R634 VTAIL.n214 VTAIL.n162 3.49141
R635 VTAIL.n193 VTAIL.n176 3.49141
R636 VTAIL.n138 VTAIL.n86 3.49141
R637 VTAIL.n117 VTAIL.n100 3.49141
R638 VTAIL.n153 VTAIL.n79 3.15567
R639 VTAIL.n229 VTAIL.n155 3.15567
R640 VTAIL.n77 VTAIL.n75 3.15567
R641 VTAIL.n253 VTAIL.n251 2.84303
R642 VTAIL.n25 VTAIL.n23 2.84303
R643 VTAIL.n181 VTAIL.n179 2.84303
R644 VTAIL.n105 VTAIL.n103 2.84303
R645 VTAIL.n266 VTAIL.n246 2.71565
R646 VTAIL.n287 VTAIL.n238 2.71565
R647 VTAIL.n38 VTAIL.n18 2.71565
R648 VTAIL.n59 VTAIL.n10 2.71565
R649 VTAIL.n213 VTAIL.n164 2.71565
R650 VTAIL.n194 VTAIL.n174 2.71565
R651 VTAIL.n137 VTAIL.n88 2.71565
R652 VTAIL.n118 VTAIL.n98 2.71565
R653 VTAIL VTAIL.n303 2.30869
R654 VTAIL.n155 VTAIL.n153 2.04791
R655 VTAIL.n75 VTAIL.n1 2.04791
R656 VTAIL.n271 VTAIL.n269 1.93989
R657 VTAIL.n284 VTAIL.n283 1.93989
R658 VTAIL.n43 VTAIL.n41 1.93989
R659 VTAIL.n56 VTAIL.n55 1.93989
R660 VTAIL.n210 VTAIL.n209 1.93989
R661 VTAIL.n198 VTAIL.n197 1.93989
R662 VTAIL.n134 VTAIL.n133 1.93989
R663 VTAIL.n122 VTAIL.n121 1.93989
R664 VTAIL.n0 VTAIL.t7 1.45638
R665 VTAIL.n0 VTAIL.t6 1.45638
R666 VTAIL.n76 VTAIL.t4 1.45638
R667 VTAIL.n76 VTAIL.t3 1.45638
R668 VTAIL.n154 VTAIL.t1 1.45638
R669 VTAIL.n154 VTAIL.t5 1.45638
R670 VTAIL.n78 VTAIL.t8 1.45638
R671 VTAIL.n78 VTAIL.t11 1.45638
R672 VTAIL.n270 VTAIL.n244 1.16414
R673 VTAIL.n280 VTAIL.n240 1.16414
R674 VTAIL.n42 VTAIL.n16 1.16414
R675 VTAIL.n52 VTAIL.n12 1.16414
R676 VTAIL.n206 VTAIL.n166 1.16414
R677 VTAIL.n201 VTAIL.n171 1.16414
R678 VTAIL.n130 VTAIL.n90 1.16414
R679 VTAIL.n125 VTAIL.n95 1.16414
R680 VTAIL VTAIL.n1 0.847483
R681 VTAIL.n276 VTAIL.n275 0.388379
R682 VTAIL.n279 VTAIL.n242 0.388379
R683 VTAIL.n48 VTAIL.n47 0.388379
R684 VTAIL.n51 VTAIL.n14 0.388379
R685 VTAIL.n205 VTAIL.n168 0.388379
R686 VTAIL.n202 VTAIL.n170 0.388379
R687 VTAIL.n129 VTAIL.n92 0.388379
R688 VTAIL.n126 VTAIL.n94 0.388379
R689 VTAIL.n259 VTAIL.n251 0.155672
R690 VTAIL.n260 VTAIL.n259 0.155672
R691 VTAIL.n260 VTAIL.n247 0.155672
R692 VTAIL.n267 VTAIL.n247 0.155672
R693 VTAIL.n268 VTAIL.n267 0.155672
R694 VTAIL.n268 VTAIL.n243 0.155672
R695 VTAIL.n277 VTAIL.n243 0.155672
R696 VTAIL.n278 VTAIL.n277 0.155672
R697 VTAIL.n278 VTAIL.n239 0.155672
R698 VTAIL.n285 VTAIL.n239 0.155672
R699 VTAIL.n286 VTAIL.n285 0.155672
R700 VTAIL.n286 VTAIL.n235 0.155672
R701 VTAIL.n293 VTAIL.n235 0.155672
R702 VTAIL.n294 VTAIL.n293 0.155672
R703 VTAIL.n294 VTAIL.n231 0.155672
R704 VTAIL.n301 VTAIL.n231 0.155672
R705 VTAIL.n31 VTAIL.n23 0.155672
R706 VTAIL.n32 VTAIL.n31 0.155672
R707 VTAIL.n32 VTAIL.n19 0.155672
R708 VTAIL.n39 VTAIL.n19 0.155672
R709 VTAIL.n40 VTAIL.n39 0.155672
R710 VTAIL.n40 VTAIL.n15 0.155672
R711 VTAIL.n49 VTAIL.n15 0.155672
R712 VTAIL.n50 VTAIL.n49 0.155672
R713 VTAIL.n50 VTAIL.n11 0.155672
R714 VTAIL.n57 VTAIL.n11 0.155672
R715 VTAIL.n58 VTAIL.n57 0.155672
R716 VTAIL.n58 VTAIL.n7 0.155672
R717 VTAIL.n65 VTAIL.n7 0.155672
R718 VTAIL.n66 VTAIL.n65 0.155672
R719 VTAIL.n66 VTAIL.n3 0.155672
R720 VTAIL.n73 VTAIL.n3 0.155672
R721 VTAIL.n227 VTAIL.n157 0.155672
R722 VTAIL.n220 VTAIL.n157 0.155672
R723 VTAIL.n220 VTAIL.n219 0.155672
R724 VTAIL.n219 VTAIL.n161 0.155672
R725 VTAIL.n212 VTAIL.n161 0.155672
R726 VTAIL.n212 VTAIL.n211 0.155672
R727 VTAIL.n211 VTAIL.n165 0.155672
R728 VTAIL.n204 VTAIL.n165 0.155672
R729 VTAIL.n204 VTAIL.n203 0.155672
R730 VTAIL.n203 VTAIL.n169 0.155672
R731 VTAIL.n196 VTAIL.n169 0.155672
R732 VTAIL.n196 VTAIL.n195 0.155672
R733 VTAIL.n195 VTAIL.n175 0.155672
R734 VTAIL.n188 VTAIL.n175 0.155672
R735 VTAIL.n188 VTAIL.n187 0.155672
R736 VTAIL.n187 VTAIL.n179 0.155672
R737 VTAIL.n151 VTAIL.n81 0.155672
R738 VTAIL.n144 VTAIL.n81 0.155672
R739 VTAIL.n144 VTAIL.n143 0.155672
R740 VTAIL.n143 VTAIL.n85 0.155672
R741 VTAIL.n136 VTAIL.n85 0.155672
R742 VTAIL.n136 VTAIL.n135 0.155672
R743 VTAIL.n135 VTAIL.n89 0.155672
R744 VTAIL.n128 VTAIL.n89 0.155672
R745 VTAIL.n128 VTAIL.n127 0.155672
R746 VTAIL.n127 VTAIL.n93 0.155672
R747 VTAIL.n120 VTAIL.n93 0.155672
R748 VTAIL.n120 VTAIL.n119 0.155672
R749 VTAIL.n119 VTAIL.n99 0.155672
R750 VTAIL.n112 VTAIL.n99 0.155672
R751 VTAIL.n112 VTAIL.n111 0.155672
R752 VTAIL.n111 VTAIL.n103 0.155672
R753 B.n928 B.n927 585
R754 B.n349 B.n145 585
R755 B.n348 B.n347 585
R756 B.n346 B.n345 585
R757 B.n344 B.n343 585
R758 B.n342 B.n341 585
R759 B.n340 B.n339 585
R760 B.n338 B.n337 585
R761 B.n336 B.n335 585
R762 B.n334 B.n333 585
R763 B.n332 B.n331 585
R764 B.n330 B.n329 585
R765 B.n328 B.n327 585
R766 B.n326 B.n325 585
R767 B.n324 B.n323 585
R768 B.n322 B.n321 585
R769 B.n320 B.n319 585
R770 B.n318 B.n317 585
R771 B.n316 B.n315 585
R772 B.n314 B.n313 585
R773 B.n312 B.n311 585
R774 B.n310 B.n309 585
R775 B.n308 B.n307 585
R776 B.n306 B.n305 585
R777 B.n304 B.n303 585
R778 B.n302 B.n301 585
R779 B.n300 B.n299 585
R780 B.n298 B.n297 585
R781 B.n296 B.n295 585
R782 B.n294 B.n293 585
R783 B.n292 B.n291 585
R784 B.n290 B.n289 585
R785 B.n288 B.n287 585
R786 B.n286 B.n285 585
R787 B.n284 B.n283 585
R788 B.n282 B.n281 585
R789 B.n280 B.n279 585
R790 B.n278 B.n277 585
R791 B.n276 B.n275 585
R792 B.n274 B.n273 585
R793 B.n272 B.n271 585
R794 B.n270 B.n269 585
R795 B.n268 B.n267 585
R796 B.n266 B.n265 585
R797 B.n264 B.n263 585
R798 B.n262 B.n261 585
R799 B.n260 B.n259 585
R800 B.n258 B.n257 585
R801 B.n256 B.n255 585
R802 B.n254 B.n253 585
R803 B.n252 B.n251 585
R804 B.n250 B.n249 585
R805 B.n248 B.n247 585
R806 B.n246 B.n245 585
R807 B.n244 B.n243 585
R808 B.n242 B.n241 585
R809 B.n240 B.n239 585
R810 B.n238 B.n237 585
R811 B.n236 B.n235 585
R812 B.n234 B.n233 585
R813 B.n232 B.n231 585
R814 B.n230 B.n229 585
R815 B.n228 B.n227 585
R816 B.n226 B.n225 585
R817 B.n224 B.n223 585
R818 B.n222 B.n221 585
R819 B.n220 B.n219 585
R820 B.n218 B.n217 585
R821 B.n216 B.n215 585
R822 B.n214 B.n213 585
R823 B.n212 B.n211 585
R824 B.n210 B.n209 585
R825 B.n208 B.n207 585
R826 B.n206 B.n205 585
R827 B.n204 B.n203 585
R828 B.n202 B.n201 585
R829 B.n200 B.n199 585
R830 B.n198 B.n197 585
R831 B.n196 B.n195 585
R832 B.n194 B.n193 585
R833 B.n192 B.n191 585
R834 B.n190 B.n189 585
R835 B.n188 B.n187 585
R836 B.n186 B.n185 585
R837 B.n184 B.n183 585
R838 B.n182 B.n181 585
R839 B.n180 B.n179 585
R840 B.n178 B.n177 585
R841 B.n176 B.n175 585
R842 B.n174 B.n173 585
R843 B.n172 B.n171 585
R844 B.n170 B.n169 585
R845 B.n168 B.n167 585
R846 B.n166 B.n165 585
R847 B.n164 B.n163 585
R848 B.n162 B.n161 585
R849 B.n160 B.n159 585
R850 B.n158 B.n157 585
R851 B.n156 B.n155 585
R852 B.n154 B.n153 585
R853 B.n95 B.n94 585
R854 B.n933 B.n932 585
R855 B.n926 B.n146 585
R856 B.n146 B.n92 585
R857 B.n925 B.n91 585
R858 B.n937 B.n91 585
R859 B.n924 B.n90 585
R860 B.n938 B.n90 585
R861 B.n923 B.n89 585
R862 B.n939 B.n89 585
R863 B.n922 B.n921 585
R864 B.n921 B.n85 585
R865 B.n920 B.n84 585
R866 B.n945 B.n84 585
R867 B.n919 B.n83 585
R868 B.n946 B.n83 585
R869 B.n918 B.n82 585
R870 B.n947 B.n82 585
R871 B.n917 B.n916 585
R872 B.n916 B.n81 585
R873 B.n915 B.n77 585
R874 B.n953 B.n77 585
R875 B.n914 B.n76 585
R876 B.n954 B.n76 585
R877 B.n913 B.n75 585
R878 B.n955 B.n75 585
R879 B.n912 B.n911 585
R880 B.n911 B.n71 585
R881 B.n910 B.n70 585
R882 B.n961 B.n70 585
R883 B.n909 B.n69 585
R884 B.n962 B.n69 585
R885 B.n908 B.n68 585
R886 B.n963 B.n68 585
R887 B.n907 B.n906 585
R888 B.n906 B.n64 585
R889 B.n905 B.n63 585
R890 B.n969 B.n63 585
R891 B.n904 B.n62 585
R892 B.n970 B.n62 585
R893 B.n903 B.n61 585
R894 B.n971 B.n61 585
R895 B.n902 B.n901 585
R896 B.n901 B.n57 585
R897 B.n900 B.n56 585
R898 B.n977 B.n56 585
R899 B.n899 B.n55 585
R900 B.n978 B.n55 585
R901 B.n898 B.n54 585
R902 B.n979 B.n54 585
R903 B.n897 B.n896 585
R904 B.n896 B.n50 585
R905 B.n895 B.n49 585
R906 B.n985 B.n49 585
R907 B.n894 B.n48 585
R908 B.n986 B.n48 585
R909 B.n893 B.n47 585
R910 B.n987 B.n47 585
R911 B.n892 B.n891 585
R912 B.n891 B.n43 585
R913 B.n890 B.n42 585
R914 B.n993 B.n42 585
R915 B.n889 B.n41 585
R916 B.n994 B.n41 585
R917 B.n888 B.n40 585
R918 B.n995 B.n40 585
R919 B.n887 B.n886 585
R920 B.n886 B.n36 585
R921 B.n885 B.n35 585
R922 B.n1001 B.n35 585
R923 B.n884 B.n34 585
R924 B.n1002 B.n34 585
R925 B.n883 B.n33 585
R926 B.n1003 B.n33 585
R927 B.n882 B.n881 585
R928 B.n881 B.n29 585
R929 B.n880 B.n28 585
R930 B.n1009 B.n28 585
R931 B.n879 B.n27 585
R932 B.n1010 B.n27 585
R933 B.n878 B.n26 585
R934 B.n1011 B.n26 585
R935 B.n877 B.n876 585
R936 B.n876 B.n22 585
R937 B.n875 B.n21 585
R938 B.n1017 B.n21 585
R939 B.n874 B.n20 585
R940 B.n1018 B.n20 585
R941 B.n873 B.n19 585
R942 B.n1019 B.n19 585
R943 B.n872 B.n871 585
R944 B.n871 B.n18 585
R945 B.n870 B.n14 585
R946 B.n1025 B.n14 585
R947 B.n869 B.n13 585
R948 B.n1026 B.n13 585
R949 B.n868 B.n12 585
R950 B.n1027 B.n12 585
R951 B.n867 B.n866 585
R952 B.n866 B.n8 585
R953 B.n865 B.n7 585
R954 B.n1033 B.n7 585
R955 B.n864 B.n6 585
R956 B.n1034 B.n6 585
R957 B.n863 B.n5 585
R958 B.n1035 B.n5 585
R959 B.n862 B.n861 585
R960 B.n861 B.n4 585
R961 B.n860 B.n350 585
R962 B.n860 B.n859 585
R963 B.n850 B.n351 585
R964 B.n352 B.n351 585
R965 B.n852 B.n851 585
R966 B.n853 B.n852 585
R967 B.n849 B.n357 585
R968 B.n357 B.n356 585
R969 B.n848 B.n847 585
R970 B.n847 B.n846 585
R971 B.n359 B.n358 585
R972 B.n839 B.n359 585
R973 B.n838 B.n837 585
R974 B.n840 B.n838 585
R975 B.n836 B.n364 585
R976 B.n364 B.n363 585
R977 B.n835 B.n834 585
R978 B.n834 B.n833 585
R979 B.n366 B.n365 585
R980 B.n367 B.n366 585
R981 B.n826 B.n825 585
R982 B.n827 B.n826 585
R983 B.n824 B.n372 585
R984 B.n372 B.n371 585
R985 B.n823 B.n822 585
R986 B.n822 B.n821 585
R987 B.n374 B.n373 585
R988 B.n375 B.n374 585
R989 B.n814 B.n813 585
R990 B.n815 B.n814 585
R991 B.n812 B.n380 585
R992 B.n380 B.n379 585
R993 B.n811 B.n810 585
R994 B.n810 B.n809 585
R995 B.n382 B.n381 585
R996 B.n383 B.n382 585
R997 B.n802 B.n801 585
R998 B.n803 B.n802 585
R999 B.n800 B.n388 585
R1000 B.n388 B.n387 585
R1001 B.n799 B.n798 585
R1002 B.n798 B.n797 585
R1003 B.n390 B.n389 585
R1004 B.n391 B.n390 585
R1005 B.n790 B.n789 585
R1006 B.n791 B.n790 585
R1007 B.n788 B.n396 585
R1008 B.n396 B.n395 585
R1009 B.n787 B.n786 585
R1010 B.n786 B.n785 585
R1011 B.n398 B.n397 585
R1012 B.n399 B.n398 585
R1013 B.n778 B.n777 585
R1014 B.n779 B.n778 585
R1015 B.n776 B.n403 585
R1016 B.n407 B.n403 585
R1017 B.n775 B.n774 585
R1018 B.n774 B.n773 585
R1019 B.n405 B.n404 585
R1020 B.n406 B.n405 585
R1021 B.n766 B.n765 585
R1022 B.n767 B.n766 585
R1023 B.n764 B.n412 585
R1024 B.n412 B.n411 585
R1025 B.n763 B.n762 585
R1026 B.n762 B.n761 585
R1027 B.n414 B.n413 585
R1028 B.n415 B.n414 585
R1029 B.n754 B.n753 585
R1030 B.n755 B.n754 585
R1031 B.n752 B.n420 585
R1032 B.n420 B.n419 585
R1033 B.n751 B.n750 585
R1034 B.n750 B.n749 585
R1035 B.n422 B.n421 585
R1036 B.n423 B.n422 585
R1037 B.n742 B.n741 585
R1038 B.n743 B.n742 585
R1039 B.n740 B.n428 585
R1040 B.n428 B.n427 585
R1041 B.n739 B.n738 585
R1042 B.n738 B.n737 585
R1043 B.n430 B.n429 585
R1044 B.n730 B.n430 585
R1045 B.n729 B.n728 585
R1046 B.n731 B.n729 585
R1047 B.n727 B.n435 585
R1048 B.n435 B.n434 585
R1049 B.n726 B.n725 585
R1050 B.n725 B.n724 585
R1051 B.n437 B.n436 585
R1052 B.n438 B.n437 585
R1053 B.n717 B.n716 585
R1054 B.n718 B.n717 585
R1055 B.n715 B.n443 585
R1056 B.n443 B.n442 585
R1057 B.n714 B.n713 585
R1058 B.n713 B.n712 585
R1059 B.n445 B.n444 585
R1060 B.n446 B.n445 585
R1061 B.n708 B.n707 585
R1062 B.n449 B.n448 585
R1063 B.n704 B.n703 585
R1064 B.n705 B.n704 585
R1065 B.n702 B.n500 585
R1066 B.n701 B.n700 585
R1067 B.n699 B.n698 585
R1068 B.n697 B.n696 585
R1069 B.n695 B.n694 585
R1070 B.n693 B.n692 585
R1071 B.n691 B.n690 585
R1072 B.n689 B.n688 585
R1073 B.n687 B.n686 585
R1074 B.n685 B.n684 585
R1075 B.n683 B.n682 585
R1076 B.n681 B.n680 585
R1077 B.n679 B.n678 585
R1078 B.n677 B.n676 585
R1079 B.n675 B.n674 585
R1080 B.n673 B.n672 585
R1081 B.n671 B.n670 585
R1082 B.n669 B.n668 585
R1083 B.n667 B.n666 585
R1084 B.n665 B.n664 585
R1085 B.n663 B.n662 585
R1086 B.n661 B.n660 585
R1087 B.n659 B.n658 585
R1088 B.n657 B.n656 585
R1089 B.n655 B.n654 585
R1090 B.n653 B.n652 585
R1091 B.n651 B.n650 585
R1092 B.n649 B.n648 585
R1093 B.n647 B.n646 585
R1094 B.n645 B.n644 585
R1095 B.n643 B.n642 585
R1096 B.n641 B.n640 585
R1097 B.n639 B.n638 585
R1098 B.n637 B.n636 585
R1099 B.n635 B.n634 585
R1100 B.n633 B.n632 585
R1101 B.n631 B.n630 585
R1102 B.n629 B.n628 585
R1103 B.n627 B.n626 585
R1104 B.n625 B.n624 585
R1105 B.n623 B.n622 585
R1106 B.n621 B.n620 585
R1107 B.n619 B.n618 585
R1108 B.n616 B.n615 585
R1109 B.n614 B.n613 585
R1110 B.n612 B.n611 585
R1111 B.n610 B.n609 585
R1112 B.n608 B.n607 585
R1113 B.n606 B.n605 585
R1114 B.n604 B.n603 585
R1115 B.n602 B.n601 585
R1116 B.n600 B.n599 585
R1117 B.n598 B.n597 585
R1118 B.n595 B.n594 585
R1119 B.n593 B.n592 585
R1120 B.n591 B.n590 585
R1121 B.n589 B.n588 585
R1122 B.n587 B.n586 585
R1123 B.n585 B.n584 585
R1124 B.n583 B.n582 585
R1125 B.n581 B.n580 585
R1126 B.n579 B.n578 585
R1127 B.n577 B.n576 585
R1128 B.n575 B.n574 585
R1129 B.n573 B.n572 585
R1130 B.n571 B.n570 585
R1131 B.n569 B.n568 585
R1132 B.n567 B.n566 585
R1133 B.n565 B.n564 585
R1134 B.n563 B.n562 585
R1135 B.n561 B.n560 585
R1136 B.n559 B.n558 585
R1137 B.n557 B.n556 585
R1138 B.n555 B.n554 585
R1139 B.n553 B.n552 585
R1140 B.n551 B.n550 585
R1141 B.n549 B.n548 585
R1142 B.n547 B.n546 585
R1143 B.n545 B.n544 585
R1144 B.n543 B.n542 585
R1145 B.n541 B.n540 585
R1146 B.n539 B.n538 585
R1147 B.n537 B.n536 585
R1148 B.n535 B.n534 585
R1149 B.n533 B.n532 585
R1150 B.n531 B.n530 585
R1151 B.n529 B.n528 585
R1152 B.n527 B.n526 585
R1153 B.n525 B.n524 585
R1154 B.n523 B.n522 585
R1155 B.n521 B.n520 585
R1156 B.n519 B.n518 585
R1157 B.n517 B.n516 585
R1158 B.n515 B.n514 585
R1159 B.n513 B.n512 585
R1160 B.n511 B.n510 585
R1161 B.n509 B.n508 585
R1162 B.n507 B.n506 585
R1163 B.n505 B.n499 585
R1164 B.n705 B.n499 585
R1165 B.n709 B.n447 585
R1166 B.n447 B.n446 585
R1167 B.n711 B.n710 585
R1168 B.n712 B.n711 585
R1169 B.n441 B.n440 585
R1170 B.n442 B.n441 585
R1171 B.n720 B.n719 585
R1172 B.n719 B.n718 585
R1173 B.n721 B.n439 585
R1174 B.n439 B.n438 585
R1175 B.n723 B.n722 585
R1176 B.n724 B.n723 585
R1177 B.n433 B.n432 585
R1178 B.n434 B.n433 585
R1179 B.n733 B.n732 585
R1180 B.n732 B.n731 585
R1181 B.n734 B.n431 585
R1182 B.n730 B.n431 585
R1183 B.n736 B.n735 585
R1184 B.n737 B.n736 585
R1185 B.n426 B.n425 585
R1186 B.n427 B.n426 585
R1187 B.n745 B.n744 585
R1188 B.n744 B.n743 585
R1189 B.n746 B.n424 585
R1190 B.n424 B.n423 585
R1191 B.n748 B.n747 585
R1192 B.n749 B.n748 585
R1193 B.n418 B.n417 585
R1194 B.n419 B.n418 585
R1195 B.n757 B.n756 585
R1196 B.n756 B.n755 585
R1197 B.n758 B.n416 585
R1198 B.n416 B.n415 585
R1199 B.n760 B.n759 585
R1200 B.n761 B.n760 585
R1201 B.n410 B.n409 585
R1202 B.n411 B.n410 585
R1203 B.n769 B.n768 585
R1204 B.n768 B.n767 585
R1205 B.n770 B.n408 585
R1206 B.n408 B.n406 585
R1207 B.n772 B.n771 585
R1208 B.n773 B.n772 585
R1209 B.n402 B.n401 585
R1210 B.n407 B.n402 585
R1211 B.n781 B.n780 585
R1212 B.n780 B.n779 585
R1213 B.n782 B.n400 585
R1214 B.n400 B.n399 585
R1215 B.n784 B.n783 585
R1216 B.n785 B.n784 585
R1217 B.n394 B.n393 585
R1218 B.n395 B.n394 585
R1219 B.n793 B.n792 585
R1220 B.n792 B.n791 585
R1221 B.n794 B.n392 585
R1222 B.n392 B.n391 585
R1223 B.n796 B.n795 585
R1224 B.n797 B.n796 585
R1225 B.n386 B.n385 585
R1226 B.n387 B.n386 585
R1227 B.n805 B.n804 585
R1228 B.n804 B.n803 585
R1229 B.n806 B.n384 585
R1230 B.n384 B.n383 585
R1231 B.n808 B.n807 585
R1232 B.n809 B.n808 585
R1233 B.n378 B.n377 585
R1234 B.n379 B.n378 585
R1235 B.n817 B.n816 585
R1236 B.n816 B.n815 585
R1237 B.n818 B.n376 585
R1238 B.n376 B.n375 585
R1239 B.n820 B.n819 585
R1240 B.n821 B.n820 585
R1241 B.n370 B.n369 585
R1242 B.n371 B.n370 585
R1243 B.n829 B.n828 585
R1244 B.n828 B.n827 585
R1245 B.n830 B.n368 585
R1246 B.n368 B.n367 585
R1247 B.n832 B.n831 585
R1248 B.n833 B.n832 585
R1249 B.n362 B.n361 585
R1250 B.n363 B.n362 585
R1251 B.n842 B.n841 585
R1252 B.n841 B.n840 585
R1253 B.n843 B.n360 585
R1254 B.n839 B.n360 585
R1255 B.n845 B.n844 585
R1256 B.n846 B.n845 585
R1257 B.n355 B.n354 585
R1258 B.n356 B.n355 585
R1259 B.n855 B.n854 585
R1260 B.n854 B.n853 585
R1261 B.n856 B.n353 585
R1262 B.n353 B.n352 585
R1263 B.n858 B.n857 585
R1264 B.n859 B.n858 585
R1265 B.n2 B.n0 585
R1266 B.n4 B.n2 585
R1267 B.n3 B.n1 585
R1268 B.n1034 B.n3 585
R1269 B.n1032 B.n1031 585
R1270 B.n1033 B.n1032 585
R1271 B.n1030 B.n9 585
R1272 B.n9 B.n8 585
R1273 B.n1029 B.n1028 585
R1274 B.n1028 B.n1027 585
R1275 B.n11 B.n10 585
R1276 B.n1026 B.n11 585
R1277 B.n1024 B.n1023 585
R1278 B.n1025 B.n1024 585
R1279 B.n1022 B.n15 585
R1280 B.n18 B.n15 585
R1281 B.n1021 B.n1020 585
R1282 B.n1020 B.n1019 585
R1283 B.n17 B.n16 585
R1284 B.n1018 B.n17 585
R1285 B.n1016 B.n1015 585
R1286 B.n1017 B.n1016 585
R1287 B.n1014 B.n23 585
R1288 B.n23 B.n22 585
R1289 B.n1013 B.n1012 585
R1290 B.n1012 B.n1011 585
R1291 B.n25 B.n24 585
R1292 B.n1010 B.n25 585
R1293 B.n1008 B.n1007 585
R1294 B.n1009 B.n1008 585
R1295 B.n1006 B.n30 585
R1296 B.n30 B.n29 585
R1297 B.n1005 B.n1004 585
R1298 B.n1004 B.n1003 585
R1299 B.n32 B.n31 585
R1300 B.n1002 B.n32 585
R1301 B.n1000 B.n999 585
R1302 B.n1001 B.n1000 585
R1303 B.n998 B.n37 585
R1304 B.n37 B.n36 585
R1305 B.n997 B.n996 585
R1306 B.n996 B.n995 585
R1307 B.n39 B.n38 585
R1308 B.n994 B.n39 585
R1309 B.n992 B.n991 585
R1310 B.n993 B.n992 585
R1311 B.n990 B.n44 585
R1312 B.n44 B.n43 585
R1313 B.n989 B.n988 585
R1314 B.n988 B.n987 585
R1315 B.n46 B.n45 585
R1316 B.n986 B.n46 585
R1317 B.n984 B.n983 585
R1318 B.n985 B.n984 585
R1319 B.n982 B.n51 585
R1320 B.n51 B.n50 585
R1321 B.n981 B.n980 585
R1322 B.n980 B.n979 585
R1323 B.n53 B.n52 585
R1324 B.n978 B.n53 585
R1325 B.n976 B.n975 585
R1326 B.n977 B.n976 585
R1327 B.n974 B.n58 585
R1328 B.n58 B.n57 585
R1329 B.n973 B.n972 585
R1330 B.n972 B.n971 585
R1331 B.n60 B.n59 585
R1332 B.n970 B.n60 585
R1333 B.n968 B.n967 585
R1334 B.n969 B.n968 585
R1335 B.n966 B.n65 585
R1336 B.n65 B.n64 585
R1337 B.n965 B.n964 585
R1338 B.n964 B.n963 585
R1339 B.n67 B.n66 585
R1340 B.n962 B.n67 585
R1341 B.n960 B.n959 585
R1342 B.n961 B.n960 585
R1343 B.n958 B.n72 585
R1344 B.n72 B.n71 585
R1345 B.n957 B.n956 585
R1346 B.n956 B.n955 585
R1347 B.n74 B.n73 585
R1348 B.n954 B.n74 585
R1349 B.n952 B.n951 585
R1350 B.n953 B.n952 585
R1351 B.n950 B.n78 585
R1352 B.n81 B.n78 585
R1353 B.n949 B.n948 585
R1354 B.n948 B.n947 585
R1355 B.n80 B.n79 585
R1356 B.n946 B.n80 585
R1357 B.n944 B.n943 585
R1358 B.n945 B.n944 585
R1359 B.n942 B.n86 585
R1360 B.n86 B.n85 585
R1361 B.n941 B.n940 585
R1362 B.n940 B.n939 585
R1363 B.n88 B.n87 585
R1364 B.n938 B.n88 585
R1365 B.n936 B.n935 585
R1366 B.n937 B.n936 585
R1367 B.n934 B.n93 585
R1368 B.n93 B.n92 585
R1369 B.n1037 B.n1036 585
R1370 B.n1036 B.n1035 585
R1371 B.n707 B.n447 545.355
R1372 B.n932 B.n93 545.355
R1373 B.n499 B.n445 545.355
R1374 B.n928 B.n146 545.355
R1375 B.n503 B.t16 381.07
R1376 B.n147 B.t8 381.07
R1377 B.n501 B.t13 381.07
R1378 B.n150 B.t18 381.07
R1379 B.n504 B.t15 310.087
R1380 B.n148 B.t9 310.087
R1381 B.n502 B.t12 310.087
R1382 B.n151 B.t19 310.087
R1383 B.n503 B.t14 307.361
R1384 B.n501 B.t10 307.361
R1385 B.n150 B.t17 307.361
R1386 B.n147 B.t6 307.361
R1387 B.n930 B.n929 256.663
R1388 B.n930 B.n144 256.663
R1389 B.n930 B.n143 256.663
R1390 B.n930 B.n142 256.663
R1391 B.n930 B.n141 256.663
R1392 B.n930 B.n140 256.663
R1393 B.n930 B.n139 256.663
R1394 B.n930 B.n138 256.663
R1395 B.n930 B.n137 256.663
R1396 B.n930 B.n136 256.663
R1397 B.n930 B.n135 256.663
R1398 B.n930 B.n134 256.663
R1399 B.n930 B.n133 256.663
R1400 B.n930 B.n132 256.663
R1401 B.n930 B.n131 256.663
R1402 B.n930 B.n130 256.663
R1403 B.n930 B.n129 256.663
R1404 B.n930 B.n128 256.663
R1405 B.n930 B.n127 256.663
R1406 B.n930 B.n126 256.663
R1407 B.n930 B.n125 256.663
R1408 B.n930 B.n124 256.663
R1409 B.n930 B.n123 256.663
R1410 B.n930 B.n122 256.663
R1411 B.n930 B.n121 256.663
R1412 B.n930 B.n120 256.663
R1413 B.n930 B.n119 256.663
R1414 B.n930 B.n118 256.663
R1415 B.n930 B.n117 256.663
R1416 B.n930 B.n116 256.663
R1417 B.n930 B.n115 256.663
R1418 B.n930 B.n114 256.663
R1419 B.n930 B.n113 256.663
R1420 B.n930 B.n112 256.663
R1421 B.n930 B.n111 256.663
R1422 B.n930 B.n110 256.663
R1423 B.n930 B.n109 256.663
R1424 B.n930 B.n108 256.663
R1425 B.n930 B.n107 256.663
R1426 B.n930 B.n106 256.663
R1427 B.n930 B.n105 256.663
R1428 B.n930 B.n104 256.663
R1429 B.n930 B.n103 256.663
R1430 B.n930 B.n102 256.663
R1431 B.n930 B.n101 256.663
R1432 B.n930 B.n100 256.663
R1433 B.n930 B.n99 256.663
R1434 B.n930 B.n98 256.663
R1435 B.n930 B.n97 256.663
R1436 B.n930 B.n96 256.663
R1437 B.n931 B.n930 256.663
R1438 B.n706 B.n705 256.663
R1439 B.n705 B.n450 256.663
R1440 B.n705 B.n451 256.663
R1441 B.n705 B.n452 256.663
R1442 B.n705 B.n453 256.663
R1443 B.n705 B.n454 256.663
R1444 B.n705 B.n455 256.663
R1445 B.n705 B.n456 256.663
R1446 B.n705 B.n457 256.663
R1447 B.n705 B.n458 256.663
R1448 B.n705 B.n459 256.663
R1449 B.n705 B.n460 256.663
R1450 B.n705 B.n461 256.663
R1451 B.n705 B.n462 256.663
R1452 B.n705 B.n463 256.663
R1453 B.n705 B.n464 256.663
R1454 B.n705 B.n465 256.663
R1455 B.n705 B.n466 256.663
R1456 B.n705 B.n467 256.663
R1457 B.n705 B.n468 256.663
R1458 B.n705 B.n469 256.663
R1459 B.n705 B.n470 256.663
R1460 B.n705 B.n471 256.663
R1461 B.n705 B.n472 256.663
R1462 B.n705 B.n473 256.663
R1463 B.n705 B.n474 256.663
R1464 B.n705 B.n475 256.663
R1465 B.n705 B.n476 256.663
R1466 B.n705 B.n477 256.663
R1467 B.n705 B.n478 256.663
R1468 B.n705 B.n479 256.663
R1469 B.n705 B.n480 256.663
R1470 B.n705 B.n481 256.663
R1471 B.n705 B.n482 256.663
R1472 B.n705 B.n483 256.663
R1473 B.n705 B.n484 256.663
R1474 B.n705 B.n485 256.663
R1475 B.n705 B.n486 256.663
R1476 B.n705 B.n487 256.663
R1477 B.n705 B.n488 256.663
R1478 B.n705 B.n489 256.663
R1479 B.n705 B.n490 256.663
R1480 B.n705 B.n491 256.663
R1481 B.n705 B.n492 256.663
R1482 B.n705 B.n493 256.663
R1483 B.n705 B.n494 256.663
R1484 B.n705 B.n495 256.663
R1485 B.n705 B.n496 256.663
R1486 B.n705 B.n497 256.663
R1487 B.n705 B.n498 256.663
R1488 B.n711 B.n447 163.367
R1489 B.n711 B.n441 163.367
R1490 B.n719 B.n441 163.367
R1491 B.n719 B.n439 163.367
R1492 B.n723 B.n439 163.367
R1493 B.n723 B.n433 163.367
R1494 B.n732 B.n433 163.367
R1495 B.n732 B.n431 163.367
R1496 B.n736 B.n431 163.367
R1497 B.n736 B.n426 163.367
R1498 B.n744 B.n426 163.367
R1499 B.n744 B.n424 163.367
R1500 B.n748 B.n424 163.367
R1501 B.n748 B.n418 163.367
R1502 B.n756 B.n418 163.367
R1503 B.n756 B.n416 163.367
R1504 B.n760 B.n416 163.367
R1505 B.n760 B.n410 163.367
R1506 B.n768 B.n410 163.367
R1507 B.n768 B.n408 163.367
R1508 B.n772 B.n408 163.367
R1509 B.n772 B.n402 163.367
R1510 B.n780 B.n402 163.367
R1511 B.n780 B.n400 163.367
R1512 B.n784 B.n400 163.367
R1513 B.n784 B.n394 163.367
R1514 B.n792 B.n394 163.367
R1515 B.n792 B.n392 163.367
R1516 B.n796 B.n392 163.367
R1517 B.n796 B.n386 163.367
R1518 B.n804 B.n386 163.367
R1519 B.n804 B.n384 163.367
R1520 B.n808 B.n384 163.367
R1521 B.n808 B.n378 163.367
R1522 B.n816 B.n378 163.367
R1523 B.n816 B.n376 163.367
R1524 B.n820 B.n376 163.367
R1525 B.n820 B.n370 163.367
R1526 B.n828 B.n370 163.367
R1527 B.n828 B.n368 163.367
R1528 B.n832 B.n368 163.367
R1529 B.n832 B.n362 163.367
R1530 B.n841 B.n362 163.367
R1531 B.n841 B.n360 163.367
R1532 B.n845 B.n360 163.367
R1533 B.n845 B.n355 163.367
R1534 B.n854 B.n355 163.367
R1535 B.n854 B.n353 163.367
R1536 B.n858 B.n353 163.367
R1537 B.n858 B.n2 163.367
R1538 B.n1036 B.n2 163.367
R1539 B.n1036 B.n3 163.367
R1540 B.n1032 B.n3 163.367
R1541 B.n1032 B.n9 163.367
R1542 B.n1028 B.n9 163.367
R1543 B.n1028 B.n11 163.367
R1544 B.n1024 B.n11 163.367
R1545 B.n1024 B.n15 163.367
R1546 B.n1020 B.n15 163.367
R1547 B.n1020 B.n17 163.367
R1548 B.n1016 B.n17 163.367
R1549 B.n1016 B.n23 163.367
R1550 B.n1012 B.n23 163.367
R1551 B.n1012 B.n25 163.367
R1552 B.n1008 B.n25 163.367
R1553 B.n1008 B.n30 163.367
R1554 B.n1004 B.n30 163.367
R1555 B.n1004 B.n32 163.367
R1556 B.n1000 B.n32 163.367
R1557 B.n1000 B.n37 163.367
R1558 B.n996 B.n37 163.367
R1559 B.n996 B.n39 163.367
R1560 B.n992 B.n39 163.367
R1561 B.n992 B.n44 163.367
R1562 B.n988 B.n44 163.367
R1563 B.n988 B.n46 163.367
R1564 B.n984 B.n46 163.367
R1565 B.n984 B.n51 163.367
R1566 B.n980 B.n51 163.367
R1567 B.n980 B.n53 163.367
R1568 B.n976 B.n53 163.367
R1569 B.n976 B.n58 163.367
R1570 B.n972 B.n58 163.367
R1571 B.n972 B.n60 163.367
R1572 B.n968 B.n60 163.367
R1573 B.n968 B.n65 163.367
R1574 B.n964 B.n65 163.367
R1575 B.n964 B.n67 163.367
R1576 B.n960 B.n67 163.367
R1577 B.n960 B.n72 163.367
R1578 B.n956 B.n72 163.367
R1579 B.n956 B.n74 163.367
R1580 B.n952 B.n74 163.367
R1581 B.n952 B.n78 163.367
R1582 B.n948 B.n78 163.367
R1583 B.n948 B.n80 163.367
R1584 B.n944 B.n80 163.367
R1585 B.n944 B.n86 163.367
R1586 B.n940 B.n86 163.367
R1587 B.n940 B.n88 163.367
R1588 B.n936 B.n88 163.367
R1589 B.n936 B.n93 163.367
R1590 B.n704 B.n449 163.367
R1591 B.n704 B.n500 163.367
R1592 B.n700 B.n699 163.367
R1593 B.n696 B.n695 163.367
R1594 B.n692 B.n691 163.367
R1595 B.n688 B.n687 163.367
R1596 B.n684 B.n683 163.367
R1597 B.n680 B.n679 163.367
R1598 B.n676 B.n675 163.367
R1599 B.n672 B.n671 163.367
R1600 B.n668 B.n667 163.367
R1601 B.n664 B.n663 163.367
R1602 B.n660 B.n659 163.367
R1603 B.n656 B.n655 163.367
R1604 B.n652 B.n651 163.367
R1605 B.n648 B.n647 163.367
R1606 B.n644 B.n643 163.367
R1607 B.n640 B.n639 163.367
R1608 B.n636 B.n635 163.367
R1609 B.n632 B.n631 163.367
R1610 B.n628 B.n627 163.367
R1611 B.n624 B.n623 163.367
R1612 B.n620 B.n619 163.367
R1613 B.n615 B.n614 163.367
R1614 B.n611 B.n610 163.367
R1615 B.n607 B.n606 163.367
R1616 B.n603 B.n602 163.367
R1617 B.n599 B.n598 163.367
R1618 B.n594 B.n593 163.367
R1619 B.n590 B.n589 163.367
R1620 B.n586 B.n585 163.367
R1621 B.n582 B.n581 163.367
R1622 B.n578 B.n577 163.367
R1623 B.n574 B.n573 163.367
R1624 B.n570 B.n569 163.367
R1625 B.n566 B.n565 163.367
R1626 B.n562 B.n561 163.367
R1627 B.n558 B.n557 163.367
R1628 B.n554 B.n553 163.367
R1629 B.n550 B.n549 163.367
R1630 B.n546 B.n545 163.367
R1631 B.n542 B.n541 163.367
R1632 B.n538 B.n537 163.367
R1633 B.n534 B.n533 163.367
R1634 B.n530 B.n529 163.367
R1635 B.n526 B.n525 163.367
R1636 B.n522 B.n521 163.367
R1637 B.n518 B.n517 163.367
R1638 B.n514 B.n513 163.367
R1639 B.n510 B.n509 163.367
R1640 B.n506 B.n499 163.367
R1641 B.n713 B.n445 163.367
R1642 B.n713 B.n443 163.367
R1643 B.n717 B.n443 163.367
R1644 B.n717 B.n437 163.367
R1645 B.n725 B.n437 163.367
R1646 B.n725 B.n435 163.367
R1647 B.n729 B.n435 163.367
R1648 B.n729 B.n430 163.367
R1649 B.n738 B.n430 163.367
R1650 B.n738 B.n428 163.367
R1651 B.n742 B.n428 163.367
R1652 B.n742 B.n422 163.367
R1653 B.n750 B.n422 163.367
R1654 B.n750 B.n420 163.367
R1655 B.n754 B.n420 163.367
R1656 B.n754 B.n414 163.367
R1657 B.n762 B.n414 163.367
R1658 B.n762 B.n412 163.367
R1659 B.n766 B.n412 163.367
R1660 B.n766 B.n405 163.367
R1661 B.n774 B.n405 163.367
R1662 B.n774 B.n403 163.367
R1663 B.n778 B.n403 163.367
R1664 B.n778 B.n398 163.367
R1665 B.n786 B.n398 163.367
R1666 B.n786 B.n396 163.367
R1667 B.n790 B.n396 163.367
R1668 B.n790 B.n390 163.367
R1669 B.n798 B.n390 163.367
R1670 B.n798 B.n388 163.367
R1671 B.n802 B.n388 163.367
R1672 B.n802 B.n382 163.367
R1673 B.n810 B.n382 163.367
R1674 B.n810 B.n380 163.367
R1675 B.n814 B.n380 163.367
R1676 B.n814 B.n374 163.367
R1677 B.n822 B.n374 163.367
R1678 B.n822 B.n372 163.367
R1679 B.n826 B.n372 163.367
R1680 B.n826 B.n366 163.367
R1681 B.n834 B.n366 163.367
R1682 B.n834 B.n364 163.367
R1683 B.n838 B.n364 163.367
R1684 B.n838 B.n359 163.367
R1685 B.n847 B.n359 163.367
R1686 B.n847 B.n357 163.367
R1687 B.n852 B.n357 163.367
R1688 B.n852 B.n351 163.367
R1689 B.n860 B.n351 163.367
R1690 B.n861 B.n860 163.367
R1691 B.n861 B.n5 163.367
R1692 B.n6 B.n5 163.367
R1693 B.n7 B.n6 163.367
R1694 B.n866 B.n7 163.367
R1695 B.n866 B.n12 163.367
R1696 B.n13 B.n12 163.367
R1697 B.n14 B.n13 163.367
R1698 B.n871 B.n14 163.367
R1699 B.n871 B.n19 163.367
R1700 B.n20 B.n19 163.367
R1701 B.n21 B.n20 163.367
R1702 B.n876 B.n21 163.367
R1703 B.n876 B.n26 163.367
R1704 B.n27 B.n26 163.367
R1705 B.n28 B.n27 163.367
R1706 B.n881 B.n28 163.367
R1707 B.n881 B.n33 163.367
R1708 B.n34 B.n33 163.367
R1709 B.n35 B.n34 163.367
R1710 B.n886 B.n35 163.367
R1711 B.n886 B.n40 163.367
R1712 B.n41 B.n40 163.367
R1713 B.n42 B.n41 163.367
R1714 B.n891 B.n42 163.367
R1715 B.n891 B.n47 163.367
R1716 B.n48 B.n47 163.367
R1717 B.n49 B.n48 163.367
R1718 B.n896 B.n49 163.367
R1719 B.n896 B.n54 163.367
R1720 B.n55 B.n54 163.367
R1721 B.n56 B.n55 163.367
R1722 B.n901 B.n56 163.367
R1723 B.n901 B.n61 163.367
R1724 B.n62 B.n61 163.367
R1725 B.n63 B.n62 163.367
R1726 B.n906 B.n63 163.367
R1727 B.n906 B.n68 163.367
R1728 B.n69 B.n68 163.367
R1729 B.n70 B.n69 163.367
R1730 B.n911 B.n70 163.367
R1731 B.n911 B.n75 163.367
R1732 B.n76 B.n75 163.367
R1733 B.n77 B.n76 163.367
R1734 B.n916 B.n77 163.367
R1735 B.n916 B.n82 163.367
R1736 B.n83 B.n82 163.367
R1737 B.n84 B.n83 163.367
R1738 B.n921 B.n84 163.367
R1739 B.n921 B.n89 163.367
R1740 B.n90 B.n89 163.367
R1741 B.n91 B.n90 163.367
R1742 B.n146 B.n91 163.367
R1743 B.n153 B.n95 163.367
R1744 B.n157 B.n156 163.367
R1745 B.n161 B.n160 163.367
R1746 B.n165 B.n164 163.367
R1747 B.n169 B.n168 163.367
R1748 B.n173 B.n172 163.367
R1749 B.n177 B.n176 163.367
R1750 B.n181 B.n180 163.367
R1751 B.n185 B.n184 163.367
R1752 B.n189 B.n188 163.367
R1753 B.n193 B.n192 163.367
R1754 B.n197 B.n196 163.367
R1755 B.n201 B.n200 163.367
R1756 B.n205 B.n204 163.367
R1757 B.n209 B.n208 163.367
R1758 B.n213 B.n212 163.367
R1759 B.n217 B.n216 163.367
R1760 B.n221 B.n220 163.367
R1761 B.n225 B.n224 163.367
R1762 B.n229 B.n228 163.367
R1763 B.n233 B.n232 163.367
R1764 B.n237 B.n236 163.367
R1765 B.n241 B.n240 163.367
R1766 B.n245 B.n244 163.367
R1767 B.n249 B.n248 163.367
R1768 B.n253 B.n252 163.367
R1769 B.n257 B.n256 163.367
R1770 B.n261 B.n260 163.367
R1771 B.n265 B.n264 163.367
R1772 B.n269 B.n268 163.367
R1773 B.n273 B.n272 163.367
R1774 B.n277 B.n276 163.367
R1775 B.n281 B.n280 163.367
R1776 B.n285 B.n284 163.367
R1777 B.n289 B.n288 163.367
R1778 B.n293 B.n292 163.367
R1779 B.n297 B.n296 163.367
R1780 B.n301 B.n300 163.367
R1781 B.n305 B.n304 163.367
R1782 B.n309 B.n308 163.367
R1783 B.n313 B.n312 163.367
R1784 B.n317 B.n316 163.367
R1785 B.n321 B.n320 163.367
R1786 B.n325 B.n324 163.367
R1787 B.n329 B.n328 163.367
R1788 B.n333 B.n332 163.367
R1789 B.n337 B.n336 163.367
R1790 B.n341 B.n340 163.367
R1791 B.n345 B.n344 163.367
R1792 B.n347 B.n145 163.367
R1793 B.n705 B.n446 78.676
R1794 B.n930 B.n92 78.676
R1795 B.n707 B.n706 71.676
R1796 B.n500 B.n450 71.676
R1797 B.n699 B.n451 71.676
R1798 B.n695 B.n452 71.676
R1799 B.n691 B.n453 71.676
R1800 B.n687 B.n454 71.676
R1801 B.n683 B.n455 71.676
R1802 B.n679 B.n456 71.676
R1803 B.n675 B.n457 71.676
R1804 B.n671 B.n458 71.676
R1805 B.n667 B.n459 71.676
R1806 B.n663 B.n460 71.676
R1807 B.n659 B.n461 71.676
R1808 B.n655 B.n462 71.676
R1809 B.n651 B.n463 71.676
R1810 B.n647 B.n464 71.676
R1811 B.n643 B.n465 71.676
R1812 B.n639 B.n466 71.676
R1813 B.n635 B.n467 71.676
R1814 B.n631 B.n468 71.676
R1815 B.n627 B.n469 71.676
R1816 B.n623 B.n470 71.676
R1817 B.n619 B.n471 71.676
R1818 B.n614 B.n472 71.676
R1819 B.n610 B.n473 71.676
R1820 B.n606 B.n474 71.676
R1821 B.n602 B.n475 71.676
R1822 B.n598 B.n476 71.676
R1823 B.n593 B.n477 71.676
R1824 B.n589 B.n478 71.676
R1825 B.n585 B.n479 71.676
R1826 B.n581 B.n480 71.676
R1827 B.n577 B.n481 71.676
R1828 B.n573 B.n482 71.676
R1829 B.n569 B.n483 71.676
R1830 B.n565 B.n484 71.676
R1831 B.n561 B.n485 71.676
R1832 B.n557 B.n486 71.676
R1833 B.n553 B.n487 71.676
R1834 B.n549 B.n488 71.676
R1835 B.n545 B.n489 71.676
R1836 B.n541 B.n490 71.676
R1837 B.n537 B.n491 71.676
R1838 B.n533 B.n492 71.676
R1839 B.n529 B.n493 71.676
R1840 B.n525 B.n494 71.676
R1841 B.n521 B.n495 71.676
R1842 B.n517 B.n496 71.676
R1843 B.n513 B.n497 71.676
R1844 B.n509 B.n498 71.676
R1845 B.n932 B.n931 71.676
R1846 B.n153 B.n96 71.676
R1847 B.n157 B.n97 71.676
R1848 B.n161 B.n98 71.676
R1849 B.n165 B.n99 71.676
R1850 B.n169 B.n100 71.676
R1851 B.n173 B.n101 71.676
R1852 B.n177 B.n102 71.676
R1853 B.n181 B.n103 71.676
R1854 B.n185 B.n104 71.676
R1855 B.n189 B.n105 71.676
R1856 B.n193 B.n106 71.676
R1857 B.n197 B.n107 71.676
R1858 B.n201 B.n108 71.676
R1859 B.n205 B.n109 71.676
R1860 B.n209 B.n110 71.676
R1861 B.n213 B.n111 71.676
R1862 B.n217 B.n112 71.676
R1863 B.n221 B.n113 71.676
R1864 B.n225 B.n114 71.676
R1865 B.n229 B.n115 71.676
R1866 B.n233 B.n116 71.676
R1867 B.n237 B.n117 71.676
R1868 B.n241 B.n118 71.676
R1869 B.n245 B.n119 71.676
R1870 B.n249 B.n120 71.676
R1871 B.n253 B.n121 71.676
R1872 B.n257 B.n122 71.676
R1873 B.n261 B.n123 71.676
R1874 B.n265 B.n124 71.676
R1875 B.n269 B.n125 71.676
R1876 B.n273 B.n126 71.676
R1877 B.n277 B.n127 71.676
R1878 B.n281 B.n128 71.676
R1879 B.n285 B.n129 71.676
R1880 B.n289 B.n130 71.676
R1881 B.n293 B.n131 71.676
R1882 B.n297 B.n132 71.676
R1883 B.n301 B.n133 71.676
R1884 B.n305 B.n134 71.676
R1885 B.n309 B.n135 71.676
R1886 B.n313 B.n136 71.676
R1887 B.n317 B.n137 71.676
R1888 B.n321 B.n138 71.676
R1889 B.n325 B.n139 71.676
R1890 B.n329 B.n140 71.676
R1891 B.n333 B.n141 71.676
R1892 B.n337 B.n142 71.676
R1893 B.n341 B.n143 71.676
R1894 B.n345 B.n144 71.676
R1895 B.n929 B.n145 71.676
R1896 B.n929 B.n928 71.676
R1897 B.n347 B.n144 71.676
R1898 B.n344 B.n143 71.676
R1899 B.n340 B.n142 71.676
R1900 B.n336 B.n141 71.676
R1901 B.n332 B.n140 71.676
R1902 B.n328 B.n139 71.676
R1903 B.n324 B.n138 71.676
R1904 B.n320 B.n137 71.676
R1905 B.n316 B.n136 71.676
R1906 B.n312 B.n135 71.676
R1907 B.n308 B.n134 71.676
R1908 B.n304 B.n133 71.676
R1909 B.n300 B.n132 71.676
R1910 B.n296 B.n131 71.676
R1911 B.n292 B.n130 71.676
R1912 B.n288 B.n129 71.676
R1913 B.n284 B.n128 71.676
R1914 B.n280 B.n127 71.676
R1915 B.n276 B.n126 71.676
R1916 B.n272 B.n125 71.676
R1917 B.n268 B.n124 71.676
R1918 B.n264 B.n123 71.676
R1919 B.n260 B.n122 71.676
R1920 B.n256 B.n121 71.676
R1921 B.n252 B.n120 71.676
R1922 B.n248 B.n119 71.676
R1923 B.n244 B.n118 71.676
R1924 B.n240 B.n117 71.676
R1925 B.n236 B.n116 71.676
R1926 B.n232 B.n115 71.676
R1927 B.n228 B.n114 71.676
R1928 B.n224 B.n113 71.676
R1929 B.n220 B.n112 71.676
R1930 B.n216 B.n111 71.676
R1931 B.n212 B.n110 71.676
R1932 B.n208 B.n109 71.676
R1933 B.n204 B.n108 71.676
R1934 B.n200 B.n107 71.676
R1935 B.n196 B.n106 71.676
R1936 B.n192 B.n105 71.676
R1937 B.n188 B.n104 71.676
R1938 B.n184 B.n103 71.676
R1939 B.n180 B.n102 71.676
R1940 B.n176 B.n101 71.676
R1941 B.n172 B.n100 71.676
R1942 B.n168 B.n99 71.676
R1943 B.n164 B.n98 71.676
R1944 B.n160 B.n97 71.676
R1945 B.n156 B.n96 71.676
R1946 B.n931 B.n95 71.676
R1947 B.n706 B.n449 71.676
R1948 B.n700 B.n450 71.676
R1949 B.n696 B.n451 71.676
R1950 B.n692 B.n452 71.676
R1951 B.n688 B.n453 71.676
R1952 B.n684 B.n454 71.676
R1953 B.n680 B.n455 71.676
R1954 B.n676 B.n456 71.676
R1955 B.n672 B.n457 71.676
R1956 B.n668 B.n458 71.676
R1957 B.n664 B.n459 71.676
R1958 B.n660 B.n460 71.676
R1959 B.n656 B.n461 71.676
R1960 B.n652 B.n462 71.676
R1961 B.n648 B.n463 71.676
R1962 B.n644 B.n464 71.676
R1963 B.n640 B.n465 71.676
R1964 B.n636 B.n466 71.676
R1965 B.n632 B.n467 71.676
R1966 B.n628 B.n468 71.676
R1967 B.n624 B.n469 71.676
R1968 B.n620 B.n470 71.676
R1969 B.n615 B.n471 71.676
R1970 B.n611 B.n472 71.676
R1971 B.n607 B.n473 71.676
R1972 B.n603 B.n474 71.676
R1973 B.n599 B.n475 71.676
R1974 B.n594 B.n476 71.676
R1975 B.n590 B.n477 71.676
R1976 B.n586 B.n478 71.676
R1977 B.n582 B.n479 71.676
R1978 B.n578 B.n480 71.676
R1979 B.n574 B.n481 71.676
R1980 B.n570 B.n482 71.676
R1981 B.n566 B.n483 71.676
R1982 B.n562 B.n484 71.676
R1983 B.n558 B.n485 71.676
R1984 B.n554 B.n486 71.676
R1985 B.n550 B.n487 71.676
R1986 B.n546 B.n488 71.676
R1987 B.n542 B.n489 71.676
R1988 B.n538 B.n490 71.676
R1989 B.n534 B.n491 71.676
R1990 B.n530 B.n492 71.676
R1991 B.n526 B.n493 71.676
R1992 B.n522 B.n494 71.676
R1993 B.n518 B.n495 71.676
R1994 B.n514 B.n496 71.676
R1995 B.n510 B.n497 71.676
R1996 B.n506 B.n498 71.676
R1997 B.n504 B.n503 70.9823
R1998 B.n502 B.n501 70.9823
R1999 B.n151 B.n150 70.9823
R2000 B.n148 B.n147 70.9823
R2001 B.n596 B.n504 59.5399
R2002 B.n617 B.n502 59.5399
R2003 B.n152 B.n151 59.5399
R2004 B.n149 B.n148 59.5399
R2005 B.n712 B.n446 39.6296
R2006 B.n712 B.n442 39.6296
R2007 B.n718 B.n442 39.6296
R2008 B.n718 B.n438 39.6296
R2009 B.n724 B.n438 39.6296
R2010 B.n724 B.n434 39.6296
R2011 B.n731 B.n434 39.6296
R2012 B.n731 B.n730 39.6296
R2013 B.n737 B.n427 39.6296
R2014 B.n743 B.n427 39.6296
R2015 B.n743 B.n423 39.6296
R2016 B.n749 B.n423 39.6296
R2017 B.n749 B.n419 39.6296
R2018 B.n755 B.n419 39.6296
R2019 B.n755 B.n415 39.6296
R2020 B.n761 B.n415 39.6296
R2021 B.n761 B.n411 39.6296
R2022 B.n767 B.n411 39.6296
R2023 B.n767 B.n406 39.6296
R2024 B.n773 B.n406 39.6296
R2025 B.n773 B.n407 39.6296
R2026 B.n779 B.n399 39.6296
R2027 B.n785 B.n399 39.6296
R2028 B.n785 B.n395 39.6296
R2029 B.n791 B.n395 39.6296
R2030 B.n791 B.n391 39.6296
R2031 B.n797 B.n391 39.6296
R2032 B.n797 B.n387 39.6296
R2033 B.n803 B.n387 39.6296
R2034 B.n803 B.n383 39.6296
R2035 B.n809 B.n383 39.6296
R2036 B.n815 B.n379 39.6296
R2037 B.n815 B.n375 39.6296
R2038 B.n821 B.n375 39.6296
R2039 B.n821 B.n371 39.6296
R2040 B.n827 B.n371 39.6296
R2041 B.n827 B.n367 39.6296
R2042 B.n833 B.n367 39.6296
R2043 B.n833 B.n363 39.6296
R2044 B.n840 B.n363 39.6296
R2045 B.n840 B.n839 39.6296
R2046 B.n846 B.n356 39.6296
R2047 B.n853 B.n356 39.6296
R2048 B.n853 B.n352 39.6296
R2049 B.n859 B.n352 39.6296
R2050 B.n859 B.n4 39.6296
R2051 B.n1035 B.n4 39.6296
R2052 B.n1035 B.n1034 39.6296
R2053 B.n1034 B.n1033 39.6296
R2054 B.n1033 B.n8 39.6296
R2055 B.n1027 B.n8 39.6296
R2056 B.n1027 B.n1026 39.6296
R2057 B.n1026 B.n1025 39.6296
R2058 B.n1019 B.n18 39.6296
R2059 B.n1019 B.n1018 39.6296
R2060 B.n1018 B.n1017 39.6296
R2061 B.n1017 B.n22 39.6296
R2062 B.n1011 B.n22 39.6296
R2063 B.n1011 B.n1010 39.6296
R2064 B.n1010 B.n1009 39.6296
R2065 B.n1009 B.n29 39.6296
R2066 B.n1003 B.n29 39.6296
R2067 B.n1003 B.n1002 39.6296
R2068 B.n1001 B.n36 39.6296
R2069 B.n995 B.n36 39.6296
R2070 B.n995 B.n994 39.6296
R2071 B.n994 B.n993 39.6296
R2072 B.n993 B.n43 39.6296
R2073 B.n987 B.n43 39.6296
R2074 B.n987 B.n986 39.6296
R2075 B.n986 B.n985 39.6296
R2076 B.n985 B.n50 39.6296
R2077 B.n979 B.n50 39.6296
R2078 B.n978 B.n977 39.6296
R2079 B.n977 B.n57 39.6296
R2080 B.n971 B.n57 39.6296
R2081 B.n971 B.n970 39.6296
R2082 B.n970 B.n969 39.6296
R2083 B.n969 B.n64 39.6296
R2084 B.n963 B.n64 39.6296
R2085 B.n963 B.n962 39.6296
R2086 B.n962 B.n961 39.6296
R2087 B.n961 B.n71 39.6296
R2088 B.n955 B.n71 39.6296
R2089 B.n955 B.n954 39.6296
R2090 B.n954 B.n953 39.6296
R2091 B.n947 B.n81 39.6296
R2092 B.n947 B.n946 39.6296
R2093 B.n946 B.n945 39.6296
R2094 B.n945 B.n85 39.6296
R2095 B.n939 B.n85 39.6296
R2096 B.n939 B.n938 39.6296
R2097 B.n938 B.n937 39.6296
R2098 B.n937 B.n92 39.6296
R2099 B.n846 B.t0 39.0469
R2100 B.n1025 B.t1 39.0469
R2101 B.n927 B.n926 35.4346
R2102 B.n934 B.n933 35.4346
R2103 B.n505 B.n444 35.4346
R2104 B.n709 B.n708 35.4346
R2105 B.t3 B.n379 29.7224
R2106 B.n1002 B.t5 29.7224
R2107 B.n730 B.t11 20.3979
R2108 B.n779 B.t4 20.3979
R2109 B.n979 B.t2 20.3979
R2110 B.n81 B.t7 20.3979
R2111 B.n737 B.t11 19.2323
R2112 B.n407 B.t4 19.2323
R2113 B.t2 B.n978 19.2323
R2114 B.n953 B.t7 19.2323
R2115 B B.n1037 18.0485
R2116 B.n933 B.n94 10.6151
R2117 B.n154 B.n94 10.6151
R2118 B.n155 B.n154 10.6151
R2119 B.n158 B.n155 10.6151
R2120 B.n159 B.n158 10.6151
R2121 B.n162 B.n159 10.6151
R2122 B.n163 B.n162 10.6151
R2123 B.n166 B.n163 10.6151
R2124 B.n167 B.n166 10.6151
R2125 B.n170 B.n167 10.6151
R2126 B.n171 B.n170 10.6151
R2127 B.n174 B.n171 10.6151
R2128 B.n175 B.n174 10.6151
R2129 B.n178 B.n175 10.6151
R2130 B.n179 B.n178 10.6151
R2131 B.n182 B.n179 10.6151
R2132 B.n183 B.n182 10.6151
R2133 B.n186 B.n183 10.6151
R2134 B.n187 B.n186 10.6151
R2135 B.n190 B.n187 10.6151
R2136 B.n191 B.n190 10.6151
R2137 B.n194 B.n191 10.6151
R2138 B.n195 B.n194 10.6151
R2139 B.n198 B.n195 10.6151
R2140 B.n199 B.n198 10.6151
R2141 B.n202 B.n199 10.6151
R2142 B.n203 B.n202 10.6151
R2143 B.n206 B.n203 10.6151
R2144 B.n207 B.n206 10.6151
R2145 B.n210 B.n207 10.6151
R2146 B.n211 B.n210 10.6151
R2147 B.n214 B.n211 10.6151
R2148 B.n215 B.n214 10.6151
R2149 B.n218 B.n215 10.6151
R2150 B.n219 B.n218 10.6151
R2151 B.n222 B.n219 10.6151
R2152 B.n223 B.n222 10.6151
R2153 B.n226 B.n223 10.6151
R2154 B.n227 B.n226 10.6151
R2155 B.n230 B.n227 10.6151
R2156 B.n231 B.n230 10.6151
R2157 B.n234 B.n231 10.6151
R2158 B.n235 B.n234 10.6151
R2159 B.n238 B.n235 10.6151
R2160 B.n239 B.n238 10.6151
R2161 B.n243 B.n242 10.6151
R2162 B.n246 B.n243 10.6151
R2163 B.n247 B.n246 10.6151
R2164 B.n250 B.n247 10.6151
R2165 B.n251 B.n250 10.6151
R2166 B.n254 B.n251 10.6151
R2167 B.n255 B.n254 10.6151
R2168 B.n258 B.n255 10.6151
R2169 B.n259 B.n258 10.6151
R2170 B.n263 B.n262 10.6151
R2171 B.n266 B.n263 10.6151
R2172 B.n267 B.n266 10.6151
R2173 B.n270 B.n267 10.6151
R2174 B.n271 B.n270 10.6151
R2175 B.n274 B.n271 10.6151
R2176 B.n275 B.n274 10.6151
R2177 B.n278 B.n275 10.6151
R2178 B.n279 B.n278 10.6151
R2179 B.n282 B.n279 10.6151
R2180 B.n283 B.n282 10.6151
R2181 B.n286 B.n283 10.6151
R2182 B.n287 B.n286 10.6151
R2183 B.n290 B.n287 10.6151
R2184 B.n291 B.n290 10.6151
R2185 B.n294 B.n291 10.6151
R2186 B.n295 B.n294 10.6151
R2187 B.n298 B.n295 10.6151
R2188 B.n299 B.n298 10.6151
R2189 B.n302 B.n299 10.6151
R2190 B.n303 B.n302 10.6151
R2191 B.n306 B.n303 10.6151
R2192 B.n307 B.n306 10.6151
R2193 B.n310 B.n307 10.6151
R2194 B.n311 B.n310 10.6151
R2195 B.n314 B.n311 10.6151
R2196 B.n315 B.n314 10.6151
R2197 B.n318 B.n315 10.6151
R2198 B.n319 B.n318 10.6151
R2199 B.n322 B.n319 10.6151
R2200 B.n323 B.n322 10.6151
R2201 B.n326 B.n323 10.6151
R2202 B.n327 B.n326 10.6151
R2203 B.n330 B.n327 10.6151
R2204 B.n331 B.n330 10.6151
R2205 B.n334 B.n331 10.6151
R2206 B.n335 B.n334 10.6151
R2207 B.n338 B.n335 10.6151
R2208 B.n339 B.n338 10.6151
R2209 B.n342 B.n339 10.6151
R2210 B.n343 B.n342 10.6151
R2211 B.n346 B.n343 10.6151
R2212 B.n348 B.n346 10.6151
R2213 B.n349 B.n348 10.6151
R2214 B.n927 B.n349 10.6151
R2215 B.n714 B.n444 10.6151
R2216 B.n715 B.n714 10.6151
R2217 B.n716 B.n715 10.6151
R2218 B.n716 B.n436 10.6151
R2219 B.n726 B.n436 10.6151
R2220 B.n727 B.n726 10.6151
R2221 B.n728 B.n727 10.6151
R2222 B.n728 B.n429 10.6151
R2223 B.n739 B.n429 10.6151
R2224 B.n740 B.n739 10.6151
R2225 B.n741 B.n740 10.6151
R2226 B.n741 B.n421 10.6151
R2227 B.n751 B.n421 10.6151
R2228 B.n752 B.n751 10.6151
R2229 B.n753 B.n752 10.6151
R2230 B.n753 B.n413 10.6151
R2231 B.n763 B.n413 10.6151
R2232 B.n764 B.n763 10.6151
R2233 B.n765 B.n764 10.6151
R2234 B.n765 B.n404 10.6151
R2235 B.n775 B.n404 10.6151
R2236 B.n776 B.n775 10.6151
R2237 B.n777 B.n776 10.6151
R2238 B.n777 B.n397 10.6151
R2239 B.n787 B.n397 10.6151
R2240 B.n788 B.n787 10.6151
R2241 B.n789 B.n788 10.6151
R2242 B.n789 B.n389 10.6151
R2243 B.n799 B.n389 10.6151
R2244 B.n800 B.n799 10.6151
R2245 B.n801 B.n800 10.6151
R2246 B.n801 B.n381 10.6151
R2247 B.n811 B.n381 10.6151
R2248 B.n812 B.n811 10.6151
R2249 B.n813 B.n812 10.6151
R2250 B.n813 B.n373 10.6151
R2251 B.n823 B.n373 10.6151
R2252 B.n824 B.n823 10.6151
R2253 B.n825 B.n824 10.6151
R2254 B.n825 B.n365 10.6151
R2255 B.n835 B.n365 10.6151
R2256 B.n836 B.n835 10.6151
R2257 B.n837 B.n836 10.6151
R2258 B.n837 B.n358 10.6151
R2259 B.n848 B.n358 10.6151
R2260 B.n849 B.n848 10.6151
R2261 B.n851 B.n849 10.6151
R2262 B.n851 B.n850 10.6151
R2263 B.n850 B.n350 10.6151
R2264 B.n862 B.n350 10.6151
R2265 B.n863 B.n862 10.6151
R2266 B.n864 B.n863 10.6151
R2267 B.n865 B.n864 10.6151
R2268 B.n867 B.n865 10.6151
R2269 B.n868 B.n867 10.6151
R2270 B.n869 B.n868 10.6151
R2271 B.n870 B.n869 10.6151
R2272 B.n872 B.n870 10.6151
R2273 B.n873 B.n872 10.6151
R2274 B.n874 B.n873 10.6151
R2275 B.n875 B.n874 10.6151
R2276 B.n877 B.n875 10.6151
R2277 B.n878 B.n877 10.6151
R2278 B.n879 B.n878 10.6151
R2279 B.n880 B.n879 10.6151
R2280 B.n882 B.n880 10.6151
R2281 B.n883 B.n882 10.6151
R2282 B.n884 B.n883 10.6151
R2283 B.n885 B.n884 10.6151
R2284 B.n887 B.n885 10.6151
R2285 B.n888 B.n887 10.6151
R2286 B.n889 B.n888 10.6151
R2287 B.n890 B.n889 10.6151
R2288 B.n892 B.n890 10.6151
R2289 B.n893 B.n892 10.6151
R2290 B.n894 B.n893 10.6151
R2291 B.n895 B.n894 10.6151
R2292 B.n897 B.n895 10.6151
R2293 B.n898 B.n897 10.6151
R2294 B.n899 B.n898 10.6151
R2295 B.n900 B.n899 10.6151
R2296 B.n902 B.n900 10.6151
R2297 B.n903 B.n902 10.6151
R2298 B.n904 B.n903 10.6151
R2299 B.n905 B.n904 10.6151
R2300 B.n907 B.n905 10.6151
R2301 B.n908 B.n907 10.6151
R2302 B.n909 B.n908 10.6151
R2303 B.n910 B.n909 10.6151
R2304 B.n912 B.n910 10.6151
R2305 B.n913 B.n912 10.6151
R2306 B.n914 B.n913 10.6151
R2307 B.n915 B.n914 10.6151
R2308 B.n917 B.n915 10.6151
R2309 B.n918 B.n917 10.6151
R2310 B.n919 B.n918 10.6151
R2311 B.n920 B.n919 10.6151
R2312 B.n922 B.n920 10.6151
R2313 B.n923 B.n922 10.6151
R2314 B.n924 B.n923 10.6151
R2315 B.n925 B.n924 10.6151
R2316 B.n926 B.n925 10.6151
R2317 B.n708 B.n448 10.6151
R2318 B.n703 B.n448 10.6151
R2319 B.n703 B.n702 10.6151
R2320 B.n702 B.n701 10.6151
R2321 B.n701 B.n698 10.6151
R2322 B.n698 B.n697 10.6151
R2323 B.n697 B.n694 10.6151
R2324 B.n694 B.n693 10.6151
R2325 B.n693 B.n690 10.6151
R2326 B.n690 B.n689 10.6151
R2327 B.n689 B.n686 10.6151
R2328 B.n686 B.n685 10.6151
R2329 B.n685 B.n682 10.6151
R2330 B.n682 B.n681 10.6151
R2331 B.n681 B.n678 10.6151
R2332 B.n678 B.n677 10.6151
R2333 B.n677 B.n674 10.6151
R2334 B.n674 B.n673 10.6151
R2335 B.n673 B.n670 10.6151
R2336 B.n670 B.n669 10.6151
R2337 B.n669 B.n666 10.6151
R2338 B.n666 B.n665 10.6151
R2339 B.n665 B.n662 10.6151
R2340 B.n662 B.n661 10.6151
R2341 B.n661 B.n658 10.6151
R2342 B.n658 B.n657 10.6151
R2343 B.n657 B.n654 10.6151
R2344 B.n654 B.n653 10.6151
R2345 B.n653 B.n650 10.6151
R2346 B.n650 B.n649 10.6151
R2347 B.n649 B.n646 10.6151
R2348 B.n646 B.n645 10.6151
R2349 B.n645 B.n642 10.6151
R2350 B.n642 B.n641 10.6151
R2351 B.n641 B.n638 10.6151
R2352 B.n638 B.n637 10.6151
R2353 B.n637 B.n634 10.6151
R2354 B.n634 B.n633 10.6151
R2355 B.n633 B.n630 10.6151
R2356 B.n630 B.n629 10.6151
R2357 B.n629 B.n626 10.6151
R2358 B.n626 B.n625 10.6151
R2359 B.n625 B.n622 10.6151
R2360 B.n622 B.n621 10.6151
R2361 B.n621 B.n618 10.6151
R2362 B.n616 B.n613 10.6151
R2363 B.n613 B.n612 10.6151
R2364 B.n612 B.n609 10.6151
R2365 B.n609 B.n608 10.6151
R2366 B.n608 B.n605 10.6151
R2367 B.n605 B.n604 10.6151
R2368 B.n604 B.n601 10.6151
R2369 B.n601 B.n600 10.6151
R2370 B.n600 B.n597 10.6151
R2371 B.n595 B.n592 10.6151
R2372 B.n592 B.n591 10.6151
R2373 B.n591 B.n588 10.6151
R2374 B.n588 B.n587 10.6151
R2375 B.n587 B.n584 10.6151
R2376 B.n584 B.n583 10.6151
R2377 B.n583 B.n580 10.6151
R2378 B.n580 B.n579 10.6151
R2379 B.n579 B.n576 10.6151
R2380 B.n576 B.n575 10.6151
R2381 B.n575 B.n572 10.6151
R2382 B.n572 B.n571 10.6151
R2383 B.n571 B.n568 10.6151
R2384 B.n568 B.n567 10.6151
R2385 B.n567 B.n564 10.6151
R2386 B.n564 B.n563 10.6151
R2387 B.n563 B.n560 10.6151
R2388 B.n560 B.n559 10.6151
R2389 B.n559 B.n556 10.6151
R2390 B.n556 B.n555 10.6151
R2391 B.n555 B.n552 10.6151
R2392 B.n552 B.n551 10.6151
R2393 B.n551 B.n548 10.6151
R2394 B.n548 B.n547 10.6151
R2395 B.n547 B.n544 10.6151
R2396 B.n544 B.n543 10.6151
R2397 B.n543 B.n540 10.6151
R2398 B.n540 B.n539 10.6151
R2399 B.n539 B.n536 10.6151
R2400 B.n536 B.n535 10.6151
R2401 B.n535 B.n532 10.6151
R2402 B.n532 B.n531 10.6151
R2403 B.n531 B.n528 10.6151
R2404 B.n528 B.n527 10.6151
R2405 B.n527 B.n524 10.6151
R2406 B.n524 B.n523 10.6151
R2407 B.n523 B.n520 10.6151
R2408 B.n520 B.n519 10.6151
R2409 B.n519 B.n516 10.6151
R2410 B.n516 B.n515 10.6151
R2411 B.n515 B.n512 10.6151
R2412 B.n512 B.n511 10.6151
R2413 B.n511 B.n508 10.6151
R2414 B.n508 B.n507 10.6151
R2415 B.n507 B.n505 10.6151
R2416 B.n710 B.n709 10.6151
R2417 B.n710 B.n440 10.6151
R2418 B.n720 B.n440 10.6151
R2419 B.n721 B.n720 10.6151
R2420 B.n722 B.n721 10.6151
R2421 B.n722 B.n432 10.6151
R2422 B.n733 B.n432 10.6151
R2423 B.n734 B.n733 10.6151
R2424 B.n735 B.n734 10.6151
R2425 B.n735 B.n425 10.6151
R2426 B.n745 B.n425 10.6151
R2427 B.n746 B.n745 10.6151
R2428 B.n747 B.n746 10.6151
R2429 B.n747 B.n417 10.6151
R2430 B.n757 B.n417 10.6151
R2431 B.n758 B.n757 10.6151
R2432 B.n759 B.n758 10.6151
R2433 B.n759 B.n409 10.6151
R2434 B.n769 B.n409 10.6151
R2435 B.n770 B.n769 10.6151
R2436 B.n771 B.n770 10.6151
R2437 B.n771 B.n401 10.6151
R2438 B.n781 B.n401 10.6151
R2439 B.n782 B.n781 10.6151
R2440 B.n783 B.n782 10.6151
R2441 B.n783 B.n393 10.6151
R2442 B.n793 B.n393 10.6151
R2443 B.n794 B.n793 10.6151
R2444 B.n795 B.n794 10.6151
R2445 B.n795 B.n385 10.6151
R2446 B.n805 B.n385 10.6151
R2447 B.n806 B.n805 10.6151
R2448 B.n807 B.n806 10.6151
R2449 B.n807 B.n377 10.6151
R2450 B.n817 B.n377 10.6151
R2451 B.n818 B.n817 10.6151
R2452 B.n819 B.n818 10.6151
R2453 B.n819 B.n369 10.6151
R2454 B.n829 B.n369 10.6151
R2455 B.n830 B.n829 10.6151
R2456 B.n831 B.n830 10.6151
R2457 B.n831 B.n361 10.6151
R2458 B.n842 B.n361 10.6151
R2459 B.n843 B.n842 10.6151
R2460 B.n844 B.n843 10.6151
R2461 B.n844 B.n354 10.6151
R2462 B.n855 B.n354 10.6151
R2463 B.n856 B.n855 10.6151
R2464 B.n857 B.n856 10.6151
R2465 B.n857 B.n0 10.6151
R2466 B.n1031 B.n1 10.6151
R2467 B.n1031 B.n1030 10.6151
R2468 B.n1030 B.n1029 10.6151
R2469 B.n1029 B.n10 10.6151
R2470 B.n1023 B.n10 10.6151
R2471 B.n1023 B.n1022 10.6151
R2472 B.n1022 B.n1021 10.6151
R2473 B.n1021 B.n16 10.6151
R2474 B.n1015 B.n16 10.6151
R2475 B.n1015 B.n1014 10.6151
R2476 B.n1014 B.n1013 10.6151
R2477 B.n1013 B.n24 10.6151
R2478 B.n1007 B.n24 10.6151
R2479 B.n1007 B.n1006 10.6151
R2480 B.n1006 B.n1005 10.6151
R2481 B.n1005 B.n31 10.6151
R2482 B.n999 B.n31 10.6151
R2483 B.n999 B.n998 10.6151
R2484 B.n998 B.n997 10.6151
R2485 B.n997 B.n38 10.6151
R2486 B.n991 B.n38 10.6151
R2487 B.n991 B.n990 10.6151
R2488 B.n990 B.n989 10.6151
R2489 B.n989 B.n45 10.6151
R2490 B.n983 B.n45 10.6151
R2491 B.n983 B.n982 10.6151
R2492 B.n982 B.n981 10.6151
R2493 B.n981 B.n52 10.6151
R2494 B.n975 B.n52 10.6151
R2495 B.n975 B.n974 10.6151
R2496 B.n974 B.n973 10.6151
R2497 B.n973 B.n59 10.6151
R2498 B.n967 B.n59 10.6151
R2499 B.n967 B.n966 10.6151
R2500 B.n966 B.n965 10.6151
R2501 B.n965 B.n66 10.6151
R2502 B.n959 B.n66 10.6151
R2503 B.n959 B.n958 10.6151
R2504 B.n958 B.n957 10.6151
R2505 B.n957 B.n73 10.6151
R2506 B.n951 B.n73 10.6151
R2507 B.n951 B.n950 10.6151
R2508 B.n950 B.n949 10.6151
R2509 B.n949 B.n79 10.6151
R2510 B.n943 B.n79 10.6151
R2511 B.n943 B.n942 10.6151
R2512 B.n942 B.n941 10.6151
R2513 B.n941 B.n87 10.6151
R2514 B.n935 B.n87 10.6151
R2515 B.n935 B.n934 10.6151
R2516 B.n809 B.t3 9.90778
R2517 B.t5 B.n1001 9.90778
R2518 B.n239 B.n152 9.36635
R2519 B.n262 B.n149 9.36635
R2520 B.n618 B.n617 9.36635
R2521 B.n596 B.n595 9.36635
R2522 B.n1037 B.n0 2.81026
R2523 B.n1037 B.n1 2.81026
R2524 B.n242 B.n152 1.24928
R2525 B.n259 B.n149 1.24928
R2526 B.n617 B.n616 1.24928
R2527 B.n597 B.n596 1.24928
R2528 B.n839 B.t0 0.583281
R2529 B.n18 B.t1 0.583281
R2530 VP.n16 VP.n15 161.3
R2531 VP.n17 VP.n12 161.3
R2532 VP.n19 VP.n18 161.3
R2533 VP.n20 VP.n11 161.3
R2534 VP.n22 VP.n21 161.3
R2535 VP.n23 VP.n10 161.3
R2536 VP.n25 VP.n24 161.3
R2537 VP.n50 VP.n49 161.3
R2538 VP.n48 VP.n1 161.3
R2539 VP.n47 VP.n46 161.3
R2540 VP.n45 VP.n2 161.3
R2541 VP.n44 VP.n43 161.3
R2542 VP.n42 VP.n3 161.3
R2543 VP.n41 VP.n40 161.3
R2544 VP.n39 VP.n4 161.3
R2545 VP.n38 VP.n37 161.3
R2546 VP.n36 VP.n5 161.3
R2547 VP.n35 VP.n34 161.3
R2548 VP.n33 VP.n6 161.3
R2549 VP.n32 VP.n31 161.3
R2550 VP.n30 VP.n7 161.3
R2551 VP.n29 VP.n28 161.3
R2552 VP.n14 VP.t4 131.531
R2553 VP.n4 VP.t2 98.4269
R2554 VP.n8 VP.t3 98.4269
R2555 VP.n0 VP.t1 98.4269
R2556 VP.n13 VP.t5 98.4269
R2557 VP.n9 VP.t0 98.4269
R2558 VP.n27 VP.n8 82.3762
R2559 VP.n51 VP.n0 82.3762
R2560 VP.n26 VP.n9 82.3762
R2561 VP.n35 VP.n6 56.5617
R2562 VP.n43 VP.n2 56.5617
R2563 VP.n18 VP.n11 56.5617
R2564 VP.n27 VP.n26 52.7647
R2565 VP.n14 VP.n13 50.1747
R2566 VP.n30 VP.n29 24.5923
R2567 VP.n31 VP.n30 24.5923
R2568 VP.n31 VP.n6 24.5923
R2569 VP.n36 VP.n35 24.5923
R2570 VP.n37 VP.n36 24.5923
R2571 VP.n37 VP.n4 24.5923
R2572 VP.n41 VP.n4 24.5923
R2573 VP.n42 VP.n41 24.5923
R2574 VP.n43 VP.n42 24.5923
R2575 VP.n47 VP.n2 24.5923
R2576 VP.n48 VP.n47 24.5923
R2577 VP.n49 VP.n48 24.5923
R2578 VP.n22 VP.n11 24.5923
R2579 VP.n23 VP.n22 24.5923
R2580 VP.n24 VP.n23 24.5923
R2581 VP.n16 VP.n13 24.5923
R2582 VP.n17 VP.n16 24.5923
R2583 VP.n18 VP.n17 24.5923
R2584 VP.n29 VP.n8 7.86989
R2585 VP.n49 VP.n0 7.86989
R2586 VP.n24 VP.n9 7.86989
R2587 VP.n15 VP.n14 3.21486
R2588 VP.n26 VP.n25 0.354861
R2589 VP.n28 VP.n27 0.354861
R2590 VP.n51 VP.n50 0.354861
R2591 VP VP.n51 0.267071
R2592 VP.n15 VP.n12 0.189894
R2593 VP.n19 VP.n12 0.189894
R2594 VP.n20 VP.n19 0.189894
R2595 VP.n21 VP.n20 0.189894
R2596 VP.n21 VP.n10 0.189894
R2597 VP.n25 VP.n10 0.189894
R2598 VP.n28 VP.n7 0.189894
R2599 VP.n32 VP.n7 0.189894
R2600 VP.n33 VP.n32 0.189894
R2601 VP.n34 VP.n33 0.189894
R2602 VP.n34 VP.n5 0.189894
R2603 VP.n38 VP.n5 0.189894
R2604 VP.n39 VP.n38 0.189894
R2605 VP.n40 VP.n39 0.189894
R2606 VP.n40 VP.n3 0.189894
R2607 VP.n44 VP.n3 0.189894
R2608 VP.n45 VP.n44 0.189894
R2609 VP.n46 VP.n45 0.189894
R2610 VP.n46 VP.n1 0.189894
R2611 VP.n50 VP.n1 0.189894
R2612 VDD1.n68 VDD1.n0 289.615
R2613 VDD1.n141 VDD1.n73 289.615
R2614 VDD1.n69 VDD1.n68 185
R2615 VDD1.n67 VDD1.n66 185
R2616 VDD1.n4 VDD1.n3 185
R2617 VDD1.n61 VDD1.n60 185
R2618 VDD1.n59 VDD1.n58 185
R2619 VDD1.n8 VDD1.n7 185
R2620 VDD1.n53 VDD1.n52 185
R2621 VDD1.n51 VDD1.n50 185
R2622 VDD1.n12 VDD1.n11 185
R2623 VDD1.n16 VDD1.n14 185
R2624 VDD1.n45 VDD1.n44 185
R2625 VDD1.n43 VDD1.n42 185
R2626 VDD1.n18 VDD1.n17 185
R2627 VDD1.n37 VDD1.n36 185
R2628 VDD1.n35 VDD1.n34 185
R2629 VDD1.n22 VDD1.n21 185
R2630 VDD1.n29 VDD1.n28 185
R2631 VDD1.n27 VDD1.n26 185
R2632 VDD1.n98 VDD1.n97 185
R2633 VDD1.n100 VDD1.n99 185
R2634 VDD1.n93 VDD1.n92 185
R2635 VDD1.n106 VDD1.n105 185
R2636 VDD1.n108 VDD1.n107 185
R2637 VDD1.n89 VDD1.n88 185
R2638 VDD1.n115 VDD1.n114 185
R2639 VDD1.n116 VDD1.n87 185
R2640 VDD1.n118 VDD1.n117 185
R2641 VDD1.n85 VDD1.n84 185
R2642 VDD1.n124 VDD1.n123 185
R2643 VDD1.n126 VDD1.n125 185
R2644 VDD1.n81 VDD1.n80 185
R2645 VDD1.n132 VDD1.n131 185
R2646 VDD1.n134 VDD1.n133 185
R2647 VDD1.n77 VDD1.n76 185
R2648 VDD1.n140 VDD1.n139 185
R2649 VDD1.n142 VDD1.n141 185
R2650 VDD1.n25 VDD1.t1 149.524
R2651 VDD1.n96 VDD1.t2 149.524
R2652 VDD1.n68 VDD1.n67 104.615
R2653 VDD1.n67 VDD1.n3 104.615
R2654 VDD1.n60 VDD1.n3 104.615
R2655 VDD1.n60 VDD1.n59 104.615
R2656 VDD1.n59 VDD1.n7 104.615
R2657 VDD1.n52 VDD1.n7 104.615
R2658 VDD1.n52 VDD1.n51 104.615
R2659 VDD1.n51 VDD1.n11 104.615
R2660 VDD1.n16 VDD1.n11 104.615
R2661 VDD1.n44 VDD1.n16 104.615
R2662 VDD1.n44 VDD1.n43 104.615
R2663 VDD1.n43 VDD1.n17 104.615
R2664 VDD1.n36 VDD1.n17 104.615
R2665 VDD1.n36 VDD1.n35 104.615
R2666 VDD1.n35 VDD1.n21 104.615
R2667 VDD1.n28 VDD1.n21 104.615
R2668 VDD1.n28 VDD1.n27 104.615
R2669 VDD1.n99 VDD1.n98 104.615
R2670 VDD1.n99 VDD1.n92 104.615
R2671 VDD1.n106 VDD1.n92 104.615
R2672 VDD1.n107 VDD1.n106 104.615
R2673 VDD1.n107 VDD1.n88 104.615
R2674 VDD1.n115 VDD1.n88 104.615
R2675 VDD1.n116 VDD1.n115 104.615
R2676 VDD1.n117 VDD1.n116 104.615
R2677 VDD1.n117 VDD1.n84 104.615
R2678 VDD1.n124 VDD1.n84 104.615
R2679 VDD1.n125 VDD1.n124 104.615
R2680 VDD1.n125 VDD1.n80 104.615
R2681 VDD1.n132 VDD1.n80 104.615
R2682 VDD1.n133 VDD1.n132 104.615
R2683 VDD1.n133 VDD1.n76 104.615
R2684 VDD1.n140 VDD1.n76 104.615
R2685 VDD1.n141 VDD1.n140 104.615
R2686 VDD1.n147 VDD1.n146 63.0632
R2687 VDD1.n149 VDD1.n148 62.3298
R2688 VDD1.n27 VDD1.t1 52.3082
R2689 VDD1.n98 VDD1.t2 52.3082
R2690 VDD1 VDD1.n72 52.0645
R2691 VDD1.n147 VDD1.n145 51.9509
R2692 VDD1.n149 VDD1.n147 47.8543
R2693 VDD1.n14 VDD1.n12 13.1884
R2694 VDD1.n118 VDD1.n85 13.1884
R2695 VDD1.n50 VDD1.n49 12.8005
R2696 VDD1.n46 VDD1.n45 12.8005
R2697 VDD1.n119 VDD1.n87 12.8005
R2698 VDD1.n123 VDD1.n122 12.8005
R2699 VDD1.n53 VDD1.n10 12.0247
R2700 VDD1.n42 VDD1.n15 12.0247
R2701 VDD1.n114 VDD1.n113 12.0247
R2702 VDD1.n126 VDD1.n83 12.0247
R2703 VDD1.n54 VDD1.n8 11.249
R2704 VDD1.n41 VDD1.n18 11.249
R2705 VDD1.n112 VDD1.n89 11.249
R2706 VDD1.n127 VDD1.n81 11.249
R2707 VDD1.n58 VDD1.n57 10.4732
R2708 VDD1.n38 VDD1.n37 10.4732
R2709 VDD1.n109 VDD1.n108 10.4732
R2710 VDD1.n131 VDD1.n130 10.4732
R2711 VDD1.n26 VDD1.n25 10.2747
R2712 VDD1.n97 VDD1.n96 10.2747
R2713 VDD1.n61 VDD1.n6 9.69747
R2714 VDD1.n34 VDD1.n20 9.69747
R2715 VDD1.n105 VDD1.n91 9.69747
R2716 VDD1.n134 VDD1.n79 9.69747
R2717 VDD1.n72 VDD1.n71 9.45567
R2718 VDD1.n145 VDD1.n144 9.45567
R2719 VDD1.n24 VDD1.n23 9.3005
R2720 VDD1.n31 VDD1.n30 9.3005
R2721 VDD1.n33 VDD1.n32 9.3005
R2722 VDD1.n20 VDD1.n19 9.3005
R2723 VDD1.n39 VDD1.n38 9.3005
R2724 VDD1.n41 VDD1.n40 9.3005
R2725 VDD1.n15 VDD1.n13 9.3005
R2726 VDD1.n47 VDD1.n46 9.3005
R2727 VDD1.n71 VDD1.n70 9.3005
R2728 VDD1.n2 VDD1.n1 9.3005
R2729 VDD1.n65 VDD1.n64 9.3005
R2730 VDD1.n63 VDD1.n62 9.3005
R2731 VDD1.n6 VDD1.n5 9.3005
R2732 VDD1.n57 VDD1.n56 9.3005
R2733 VDD1.n55 VDD1.n54 9.3005
R2734 VDD1.n10 VDD1.n9 9.3005
R2735 VDD1.n49 VDD1.n48 9.3005
R2736 VDD1.n144 VDD1.n143 9.3005
R2737 VDD1.n138 VDD1.n137 9.3005
R2738 VDD1.n136 VDD1.n135 9.3005
R2739 VDD1.n79 VDD1.n78 9.3005
R2740 VDD1.n130 VDD1.n129 9.3005
R2741 VDD1.n128 VDD1.n127 9.3005
R2742 VDD1.n83 VDD1.n82 9.3005
R2743 VDD1.n122 VDD1.n121 9.3005
R2744 VDD1.n95 VDD1.n94 9.3005
R2745 VDD1.n102 VDD1.n101 9.3005
R2746 VDD1.n104 VDD1.n103 9.3005
R2747 VDD1.n91 VDD1.n90 9.3005
R2748 VDD1.n110 VDD1.n109 9.3005
R2749 VDD1.n112 VDD1.n111 9.3005
R2750 VDD1.n113 VDD1.n86 9.3005
R2751 VDD1.n120 VDD1.n119 9.3005
R2752 VDD1.n75 VDD1.n74 9.3005
R2753 VDD1.n62 VDD1.n4 8.92171
R2754 VDD1.n33 VDD1.n22 8.92171
R2755 VDD1.n104 VDD1.n93 8.92171
R2756 VDD1.n135 VDD1.n77 8.92171
R2757 VDD1.n66 VDD1.n65 8.14595
R2758 VDD1.n30 VDD1.n29 8.14595
R2759 VDD1.n101 VDD1.n100 8.14595
R2760 VDD1.n139 VDD1.n138 8.14595
R2761 VDD1.n72 VDD1.n0 7.3702
R2762 VDD1.n69 VDD1.n2 7.3702
R2763 VDD1.n26 VDD1.n24 7.3702
R2764 VDD1.n97 VDD1.n95 7.3702
R2765 VDD1.n142 VDD1.n75 7.3702
R2766 VDD1.n145 VDD1.n73 7.3702
R2767 VDD1.n70 VDD1.n0 6.59444
R2768 VDD1.n70 VDD1.n69 6.59444
R2769 VDD1.n143 VDD1.n142 6.59444
R2770 VDD1.n143 VDD1.n73 6.59444
R2771 VDD1.n66 VDD1.n2 5.81868
R2772 VDD1.n29 VDD1.n24 5.81868
R2773 VDD1.n100 VDD1.n95 5.81868
R2774 VDD1.n139 VDD1.n75 5.81868
R2775 VDD1.n65 VDD1.n4 5.04292
R2776 VDD1.n30 VDD1.n22 5.04292
R2777 VDD1.n101 VDD1.n93 5.04292
R2778 VDD1.n138 VDD1.n77 5.04292
R2779 VDD1.n62 VDD1.n61 4.26717
R2780 VDD1.n34 VDD1.n33 4.26717
R2781 VDD1.n105 VDD1.n104 4.26717
R2782 VDD1.n135 VDD1.n134 4.26717
R2783 VDD1.n58 VDD1.n6 3.49141
R2784 VDD1.n37 VDD1.n20 3.49141
R2785 VDD1.n108 VDD1.n91 3.49141
R2786 VDD1.n131 VDD1.n79 3.49141
R2787 VDD1.n25 VDD1.n23 2.84303
R2788 VDD1.n96 VDD1.n94 2.84303
R2789 VDD1.n57 VDD1.n8 2.71565
R2790 VDD1.n38 VDD1.n18 2.71565
R2791 VDD1.n109 VDD1.n89 2.71565
R2792 VDD1.n130 VDD1.n81 2.71565
R2793 VDD1.n54 VDD1.n53 1.93989
R2794 VDD1.n42 VDD1.n41 1.93989
R2795 VDD1.n114 VDD1.n112 1.93989
R2796 VDD1.n127 VDD1.n126 1.93989
R2797 VDD1.n148 VDD1.t0 1.45638
R2798 VDD1.n148 VDD1.t5 1.45638
R2799 VDD1.n146 VDD1.t3 1.45638
R2800 VDD1.n146 VDD1.t4 1.45638
R2801 VDD1.n50 VDD1.n10 1.16414
R2802 VDD1.n45 VDD1.n15 1.16414
R2803 VDD1.n113 VDD1.n87 1.16414
R2804 VDD1.n123 VDD1.n83 1.16414
R2805 VDD1 VDD1.n149 0.731103
R2806 VDD1.n49 VDD1.n12 0.388379
R2807 VDD1.n46 VDD1.n14 0.388379
R2808 VDD1.n119 VDD1.n118 0.388379
R2809 VDD1.n122 VDD1.n85 0.388379
R2810 VDD1.n71 VDD1.n1 0.155672
R2811 VDD1.n64 VDD1.n1 0.155672
R2812 VDD1.n64 VDD1.n63 0.155672
R2813 VDD1.n63 VDD1.n5 0.155672
R2814 VDD1.n56 VDD1.n5 0.155672
R2815 VDD1.n56 VDD1.n55 0.155672
R2816 VDD1.n55 VDD1.n9 0.155672
R2817 VDD1.n48 VDD1.n9 0.155672
R2818 VDD1.n48 VDD1.n47 0.155672
R2819 VDD1.n47 VDD1.n13 0.155672
R2820 VDD1.n40 VDD1.n13 0.155672
R2821 VDD1.n40 VDD1.n39 0.155672
R2822 VDD1.n39 VDD1.n19 0.155672
R2823 VDD1.n32 VDD1.n19 0.155672
R2824 VDD1.n32 VDD1.n31 0.155672
R2825 VDD1.n31 VDD1.n23 0.155672
R2826 VDD1.n102 VDD1.n94 0.155672
R2827 VDD1.n103 VDD1.n102 0.155672
R2828 VDD1.n103 VDD1.n90 0.155672
R2829 VDD1.n110 VDD1.n90 0.155672
R2830 VDD1.n111 VDD1.n110 0.155672
R2831 VDD1.n111 VDD1.n86 0.155672
R2832 VDD1.n120 VDD1.n86 0.155672
R2833 VDD1.n121 VDD1.n120 0.155672
R2834 VDD1.n121 VDD1.n82 0.155672
R2835 VDD1.n128 VDD1.n82 0.155672
R2836 VDD1.n129 VDD1.n128 0.155672
R2837 VDD1.n129 VDD1.n78 0.155672
R2838 VDD1.n136 VDD1.n78 0.155672
R2839 VDD1.n137 VDD1.n136 0.155672
R2840 VDD1.n137 VDD1.n74 0.155672
R2841 VDD1.n144 VDD1.n74 0.155672
C0 VDD1 VDD2 1.69253f
C1 VTAIL VN 8.1542f
C2 VDD1 VN 0.152162f
C3 VP VDD2 0.52075f
C4 VTAIL VDD1 8.48026f
C5 VP VN 7.93174f
C6 VN VDD2 7.89362f
C7 VTAIL VP 8.16846f
C8 VDD1 VP 8.25891f
C9 VTAIL VDD2 8.536361f
C10 VDD2 B 6.826932f
C11 VDD1 B 6.991603f
C12 VTAIL B 8.940211f
C13 VN B 15.158879f
C14 VP B 13.836947f
C15 VDD1.n0 B 0.032181f
C16 VDD1.n1 B 0.021648f
C17 VDD1.n2 B 0.011633f
C18 VDD1.n3 B 0.027496f
C19 VDD1.n4 B 0.012317f
C20 VDD1.n5 B 0.021648f
C21 VDD1.n6 B 0.011633f
C22 VDD1.n7 B 0.027496f
C23 VDD1.n8 B 0.012317f
C24 VDD1.n9 B 0.021648f
C25 VDD1.n10 B 0.011633f
C26 VDD1.n11 B 0.027496f
C27 VDD1.n12 B 0.011975f
C28 VDD1.n13 B 0.021648f
C29 VDD1.n14 B 0.011975f
C30 VDD1.n15 B 0.011633f
C31 VDD1.n16 B 0.027496f
C32 VDD1.n17 B 0.027496f
C33 VDD1.n18 B 0.012317f
C34 VDD1.n19 B 0.021648f
C35 VDD1.n20 B 0.011633f
C36 VDD1.n21 B 0.027496f
C37 VDD1.n22 B 0.012317f
C38 VDD1.n23 B 1.24618f
C39 VDD1.n24 B 0.011633f
C40 VDD1.t1 B 0.046625f
C41 VDD1.n25 B 0.16938f
C42 VDD1.n26 B 0.019438f
C43 VDD1.n27 B 0.020622f
C44 VDD1.n28 B 0.027496f
C45 VDD1.n29 B 0.012317f
C46 VDD1.n30 B 0.011633f
C47 VDD1.n31 B 0.021648f
C48 VDD1.n32 B 0.021648f
C49 VDD1.n33 B 0.011633f
C50 VDD1.n34 B 0.012317f
C51 VDD1.n35 B 0.027496f
C52 VDD1.n36 B 0.027496f
C53 VDD1.n37 B 0.012317f
C54 VDD1.n38 B 0.011633f
C55 VDD1.n39 B 0.021648f
C56 VDD1.n40 B 0.021648f
C57 VDD1.n41 B 0.011633f
C58 VDD1.n42 B 0.012317f
C59 VDD1.n43 B 0.027496f
C60 VDD1.n44 B 0.027496f
C61 VDD1.n45 B 0.012317f
C62 VDD1.n46 B 0.011633f
C63 VDD1.n47 B 0.021648f
C64 VDD1.n48 B 0.021648f
C65 VDD1.n49 B 0.011633f
C66 VDD1.n50 B 0.012317f
C67 VDD1.n51 B 0.027496f
C68 VDD1.n52 B 0.027496f
C69 VDD1.n53 B 0.012317f
C70 VDD1.n54 B 0.011633f
C71 VDD1.n55 B 0.021648f
C72 VDD1.n56 B 0.021648f
C73 VDD1.n57 B 0.011633f
C74 VDD1.n58 B 0.012317f
C75 VDD1.n59 B 0.027496f
C76 VDD1.n60 B 0.027496f
C77 VDD1.n61 B 0.012317f
C78 VDD1.n62 B 0.011633f
C79 VDD1.n63 B 0.021648f
C80 VDD1.n64 B 0.021648f
C81 VDD1.n65 B 0.011633f
C82 VDD1.n66 B 0.012317f
C83 VDD1.n67 B 0.027496f
C84 VDD1.n68 B 0.062623f
C85 VDD1.n69 B 0.012317f
C86 VDD1.n70 B 0.011633f
C87 VDD1.n71 B 0.051222f
C88 VDD1.n72 B 0.060182f
C89 VDD1.n73 B 0.032181f
C90 VDD1.n74 B 0.021648f
C91 VDD1.n75 B 0.011633f
C92 VDD1.n76 B 0.027496f
C93 VDD1.n77 B 0.012317f
C94 VDD1.n78 B 0.021648f
C95 VDD1.n79 B 0.011633f
C96 VDD1.n80 B 0.027496f
C97 VDD1.n81 B 0.012317f
C98 VDD1.n82 B 0.021648f
C99 VDD1.n83 B 0.011633f
C100 VDD1.n84 B 0.027496f
C101 VDD1.n85 B 0.011975f
C102 VDD1.n86 B 0.021648f
C103 VDD1.n87 B 0.012317f
C104 VDD1.n88 B 0.027496f
C105 VDD1.n89 B 0.012317f
C106 VDD1.n90 B 0.021648f
C107 VDD1.n91 B 0.011633f
C108 VDD1.n92 B 0.027496f
C109 VDD1.n93 B 0.012317f
C110 VDD1.n94 B 1.24618f
C111 VDD1.n95 B 0.011633f
C112 VDD1.t2 B 0.046625f
C113 VDD1.n96 B 0.16938f
C114 VDD1.n97 B 0.019438f
C115 VDD1.n98 B 0.020622f
C116 VDD1.n99 B 0.027496f
C117 VDD1.n100 B 0.012317f
C118 VDD1.n101 B 0.011633f
C119 VDD1.n102 B 0.021648f
C120 VDD1.n103 B 0.021648f
C121 VDD1.n104 B 0.011633f
C122 VDD1.n105 B 0.012317f
C123 VDD1.n106 B 0.027496f
C124 VDD1.n107 B 0.027496f
C125 VDD1.n108 B 0.012317f
C126 VDD1.n109 B 0.011633f
C127 VDD1.n110 B 0.021648f
C128 VDD1.n111 B 0.021648f
C129 VDD1.n112 B 0.011633f
C130 VDD1.n113 B 0.011633f
C131 VDD1.n114 B 0.012317f
C132 VDD1.n115 B 0.027496f
C133 VDD1.n116 B 0.027496f
C134 VDD1.n117 B 0.027496f
C135 VDD1.n118 B 0.011975f
C136 VDD1.n119 B 0.011633f
C137 VDD1.n120 B 0.021648f
C138 VDD1.n121 B 0.021648f
C139 VDD1.n122 B 0.011633f
C140 VDD1.n123 B 0.012317f
C141 VDD1.n124 B 0.027496f
C142 VDD1.n125 B 0.027496f
C143 VDD1.n126 B 0.012317f
C144 VDD1.n127 B 0.011633f
C145 VDD1.n128 B 0.021648f
C146 VDD1.n129 B 0.021648f
C147 VDD1.n130 B 0.011633f
C148 VDD1.n131 B 0.012317f
C149 VDD1.n132 B 0.027496f
C150 VDD1.n133 B 0.027496f
C151 VDD1.n134 B 0.012317f
C152 VDD1.n135 B 0.011633f
C153 VDD1.n136 B 0.021648f
C154 VDD1.n137 B 0.021648f
C155 VDD1.n138 B 0.011633f
C156 VDD1.n139 B 0.012317f
C157 VDD1.n140 B 0.027496f
C158 VDD1.n141 B 0.062623f
C159 VDD1.n142 B 0.012317f
C160 VDD1.n143 B 0.011633f
C161 VDD1.n144 B 0.051222f
C162 VDD1.n145 B 0.059399f
C163 VDD1.t3 B 0.232657f
C164 VDD1.t4 B 0.232657f
C165 VDD1.n146 B 2.09383f
C166 VDD1.n147 B 2.80605f
C167 VDD1.t0 B 0.232657f
C168 VDD1.t5 B 0.232657f
C169 VDD1.n148 B 2.08847f
C170 VDD1.n149 B 2.70091f
C171 VP.t1 B 2.45663f
C172 VP.n0 B 0.927871f
C173 VP.n1 B 0.019842f
C174 VP.n2 B 0.024452f
C175 VP.n3 B 0.019842f
C176 VP.t2 B 2.45663f
C177 VP.n4 B 0.876247f
C178 VP.n5 B 0.019842f
C179 VP.n6 B 0.024452f
C180 VP.n7 B 0.019842f
C181 VP.t3 B 2.45663f
C182 VP.n8 B 0.927871f
C183 VP.t0 B 2.45663f
C184 VP.n9 B 0.927871f
C185 VP.n10 B 0.019842f
C186 VP.n11 B 0.024452f
C187 VP.n12 B 0.019842f
C188 VP.t5 B 2.45663f
C189 VP.n13 B 0.934853f
C190 VP.t4 B 2.70836f
C191 VP.n14 B 0.884955f
C192 VP.n15 B 0.241605f
C193 VP.n16 B 0.036796f
C194 VP.n17 B 0.036796f
C195 VP.n18 B 0.033236f
C196 VP.n19 B 0.019842f
C197 VP.n20 B 0.019842f
C198 VP.n21 B 0.019842f
C199 VP.n22 B 0.036796f
C200 VP.n23 B 0.036796f
C201 VP.n24 B 0.024443f
C202 VP.n25 B 0.03202f
C203 VP.n26 B 1.22177f
C204 VP.n27 B 1.23533f
C205 VP.n28 B 0.03202f
C206 VP.n29 B 0.024443f
C207 VP.n30 B 0.036796f
C208 VP.n31 B 0.036796f
C209 VP.n32 B 0.019842f
C210 VP.n33 B 0.019842f
C211 VP.n34 B 0.019842f
C212 VP.n35 B 0.033236f
C213 VP.n36 B 0.036796f
C214 VP.n37 B 0.036796f
C215 VP.n38 B 0.019842f
C216 VP.n39 B 0.019842f
C217 VP.n40 B 0.019842f
C218 VP.n41 B 0.036796f
C219 VP.n42 B 0.036796f
C220 VP.n43 B 0.033236f
C221 VP.n44 B 0.019842f
C222 VP.n45 B 0.019842f
C223 VP.n46 B 0.019842f
C224 VP.n47 B 0.036796f
C225 VP.n48 B 0.036796f
C226 VP.n49 B 0.024443f
C227 VP.n50 B 0.03202f
C228 VP.n51 B 0.053007f
C229 VTAIL.t7 B 0.255492f
C230 VTAIL.t6 B 0.255492f
C231 VTAIL.n0 B 2.22272f
C232 VTAIL.n1 B 0.458215f
C233 VTAIL.n2 B 0.03534f
C234 VTAIL.n3 B 0.023773f
C235 VTAIL.n4 B 0.012775f
C236 VTAIL.n5 B 0.030195f
C237 VTAIL.n6 B 0.013526f
C238 VTAIL.n7 B 0.023773f
C239 VTAIL.n8 B 0.012775f
C240 VTAIL.n9 B 0.030195f
C241 VTAIL.n10 B 0.013526f
C242 VTAIL.n11 B 0.023773f
C243 VTAIL.n12 B 0.012775f
C244 VTAIL.n13 B 0.030195f
C245 VTAIL.n14 B 0.01315f
C246 VTAIL.n15 B 0.023773f
C247 VTAIL.n16 B 0.013526f
C248 VTAIL.n17 B 0.030195f
C249 VTAIL.n18 B 0.013526f
C250 VTAIL.n19 B 0.023773f
C251 VTAIL.n20 B 0.012775f
C252 VTAIL.n21 B 0.030195f
C253 VTAIL.n22 B 0.013526f
C254 VTAIL.n23 B 1.36849f
C255 VTAIL.n24 B 0.012775f
C256 VTAIL.t0 B 0.051201f
C257 VTAIL.n25 B 0.186003f
C258 VTAIL.n26 B 0.021345f
C259 VTAIL.n27 B 0.022646f
C260 VTAIL.n28 B 0.030195f
C261 VTAIL.n29 B 0.013526f
C262 VTAIL.n30 B 0.012775f
C263 VTAIL.n31 B 0.023773f
C264 VTAIL.n32 B 0.023773f
C265 VTAIL.n33 B 0.012775f
C266 VTAIL.n34 B 0.013526f
C267 VTAIL.n35 B 0.030195f
C268 VTAIL.n36 B 0.030195f
C269 VTAIL.n37 B 0.013526f
C270 VTAIL.n38 B 0.012775f
C271 VTAIL.n39 B 0.023773f
C272 VTAIL.n40 B 0.023773f
C273 VTAIL.n41 B 0.012775f
C274 VTAIL.n42 B 0.012775f
C275 VTAIL.n43 B 0.013526f
C276 VTAIL.n44 B 0.030195f
C277 VTAIL.n45 B 0.030195f
C278 VTAIL.n46 B 0.030195f
C279 VTAIL.n47 B 0.01315f
C280 VTAIL.n48 B 0.012775f
C281 VTAIL.n49 B 0.023773f
C282 VTAIL.n50 B 0.023773f
C283 VTAIL.n51 B 0.012775f
C284 VTAIL.n52 B 0.013526f
C285 VTAIL.n53 B 0.030195f
C286 VTAIL.n54 B 0.030195f
C287 VTAIL.n55 B 0.013526f
C288 VTAIL.n56 B 0.012775f
C289 VTAIL.n57 B 0.023773f
C290 VTAIL.n58 B 0.023773f
C291 VTAIL.n59 B 0.012775f
C292 VTAIL.n60 B 0.013526f
C293 VTAIL.n61 B 0.030195f
C294 VTAIL.n62 B 0.030195f
C295 VTAIL.n63 B 0.013526f
C296 VTAIL.n64 B 0.012775f
C297 VTAIL.n65 B 0.023773f
C298 VTAIL.n66 B 0.023773f
C299 VTAIL.n67 B 0.012775f
C300 VTAIL.n68 B 0.013526f
C301 VTAIL.n69 B 0.030195f
C302 VTAIL.n70 B 0.06877f
C303 VTAIL.n71 B 0.013526f
C304 VTAIL.n72 B 0.012775f
C305 VTAIL.n73 B 0.056249f
C306 VTAIL.n74 B 0.038869f
C307 VTAIL.n75 B 0.419566f
C308 VTAIL.t4 B 0.255492f
C309 VTAIL.t3 B 0.255492f
C310 VTAIL.n76 B 2.22272f
C311 VTAIL.n77 B 2.1826f
C312 VTAIL.t8 B 0.255492f
C313 VTAIL.t11 B 0.255492f
C314 VTAIL.n78 B 2.22273f
C315 VTAIL.n79 B 2.18258f
C316 VTAIL.n80 B 0.03534f
C317 VTAIL.n81 B 0.023773f
C318 VTAIL.n82 B 0.012775f
C319 VTAIL.n83 B 0.030195f
C320 VTAIL.n84 B 0.013526f
C321 VTAIL.n85 B 0.023773f
C322 VTAIL.n86 B 0.012775f
C323 VTAIL.n87 B 0.030195f
C324 VTAIL.n88 B 0.013526f
C325 VTAIL.n89 B 0.023773f
C326 VTAIL.n90 B 0.012775f
C327 VTAIL.n91 B 0.030195f
C328 VTAIL.n92 B 0.01315f
C329 VTAIL.n93 B 0.023773f
C330 VTAIL.n94 B 0.01315f
C331 VTAIL.n95 B 0.012775f
C332 VTAIL.n96 B 0.030195f
C333 VTAIL.n97 B 0.030195f
C334 VTAIL.n98 B 0.013526f
C335 VTAIL.n99 B 0.023773f
C336 VTAIL.n100 B 0.012775f
C337 VTAIL.n101 B 0.030195f
C338 VTAIL.n102 B 0.013526f
C339 VTAIL.n103 B 1.36849f
C340 VTAIL.n104 B 0.012775f
C341 VTAIL.t10 B 0.051201f
C342 VTAIL.n105 B 0.186004f
C343 VTAIL.n106 B 0.021345f
C344 VTAIL.n107 B 0.022646f
C345 VTAIL.n108 B 0.030195f
C346 VTAIL.n109 B 0.013526f
C347 VTAIL.n110 B 0.012775f
C348 VTAIL.n111 B 0.023773f
C349 VTAIL.n112 B 0.023773f
C350 VTAIL.n113 B 0.012775f
C351 VTAIL.n114 B 0.013526f
C352 VTAIL.n115 B 0.030195f
C353 VTAIL.n116 B 0.030195f
C354 VTAIL.n117 B 0.013526f
C355 VTAIL.n118 B 0.012775f
C356 VTAIL.n119 B 0.023773f
C357 VTAIL.n120 B 0.023773f
C358 VTAIL.n121 B 0.012775f
C359 VTAIL.n122 B 0.013526f
C360 VTAIL.n123 B 0.030195f
C361 VTAIL.n124 B 0.030195f
C362 VTAIL.n125 B 0.013526f
C363 VTAIL.n126 B 0.012775f
C364 VTAIL.n127 B 0.023773f
C365 VTAIL.n128 B 0.023773f
C366 VTAIL.n129 B 0.012775f
C367 VTAIL.n130 B 0.013526f
C368 VTAIL.n131 B 0.030195f
C369 VTAIL.n132 B 0.030195f
C370 VTAIL.n133 B 0.013526f
C371 VTAIL.n134 B 0.012775f
C372 VTAIL.n135 B 0.023773f
C373 VTAIL.n136 B 0.023773f
C374 VTAIL.n137 B 0.012775f
C375 VTAIL.n138 B 0.013526f
C376 VTAIL.n139 B 0.030195f
C377 VTAIL.n140 B 0.030195f
C378 VTAIL.n141 B 0.013526f
C379 VTAIL.n142 B 0.012775f
C380 VTAIL.n143 B 0.023773f
C381 VTAIL.n144 B 0.023773f
C382 VTAIL.n145 B 0.012775f
C383 VTAIL.n146 B 0.013526f
C384 VTAIL.n147 B 0.030195f
C385 VTAIL.n148 B 0.06877f
C386 VTAIL.n149 B 0.013526f
C387 VTAIL.n150 B 0.012775f
C388 VTAIL.n151 B 0.056249f
C389 VTAIL.n152 B 0.038869f
C390 VTAIL.n153 B 0.419566f
C391 VTAIL.t1 B 0.255492f
C392 VTAIL.t5 B 0.255492f
C393 VTAIL.n154 B 2.22273f
C394 VTAIL.n155 B 0.635015f
C395 VTAIL.n156 B 0.03534f
C396 VTAIL.n157 B 0.023773f
C397 VTAIL.n158 B 0.012775f
C398 VTAIL.n159 B 0.030195f
C399 VTAIL.n160 B 0.013526f
C400 VTAIL.n161 B 0.023773f
C401 VTAIL.n162 B 0.012775f
C402 VTAIL.n163 B 0.030195f
C403 VTAIL.n164 B 0.013526f
C404 VTAIL.n165 B 0.023773f
C405 VTAIL.n166 B 0.012775f
C406 VTAIL.n167 B 0.030195f
C407 VTAIL.n168 B 0.01315f
C408 VTAIL.n169 B 0.023773f
C409 VTAIL.n170 B 0.01315f
C410 VTAIL.n171 B 0.012775f
C411 VTAIL.n172 B 0.030195f
C412 VTAIL.n173 B 0.030195f
C413 VTAIL.n174 B 0.013526f
C414 VTAIL.n175 B 0.023773f
C415 VTAIL.n176 B 0.012775f
C416 VTAIL.n177 B 0.030195f
C417 VTAIL.n178 B 0.013526f
C418 VTAIL.n179 B 1.36849f
C419 VTAIL.n180 B 0.012775f
C420 VTAIL.t2 B 0.051201f
C421 VTAIL.n181 B 0.186004f
C422 VTAIL.n182 B 0.021345f
C423 VTAIL.n183 B 0.022646f
C424 VTAIL.n184 B 0.030195f
C425 VTAIL.n185 B 0.013526f
C426 VTAIL.n186 B 0.012775f
C427 VTAIL.n187 B 0.023773f
C428 VTAIL.n188 B 0.023773f
C429 VTAIL.n189 B 0.012775f
C430 VTAIL.n190 B 0.013526f
C431 VTAIL.n191 B 0.030195f
C432 VTAIL.n192 B 0.030195f
C433 VTAIL.n193 B 0.013526f
C434 VTAIL.n194 B 0.012775f
C435 VTAIL.n195 B 0.023773f
C436 VTAIL.n196 B 0.023773f
C437 VTAIL.n197 B 0.012775f
C438 VTAIL.n198 B 0.013526f
C439 VTAIL.n199 B 0.030195f
C440 VTAIL.n200 B 0.030195f
C441 VTAIL.n201 B 0.013526f
C442 VTAIL.n202 B 0.012775f
C443 VTAIL.n203 B 0.023773f
C444 VTAIL.n204 B 0.023773f
C445 VTAIL.n205 B 0.012775f
C446 VTAIL.n206 B 0.013526f
C447 VTAIL.n207 B 0.030195f
C448 VTAIL.n208 B 0.030195f
C449 VTAIL.n209 B 0.013526f
C450 VTAIL.n210 B 0.012775f
C451 VTAIL.n211 B 0.023773f
C452 VTAIL.n212 B 0.023773f
C453 VTAIL.n213 B 0.012775f
C454 VTAIL.n214 B 0.013526f
C455 VTAIL.n215 B 0.030195f
C456 VTAIL.n216 B 0.030195f
C457 VTAIL.n217 B 0.013526f
C458 VTAIL.n218 B 0.012775f
C459 VTAIL.n219 B 0.023773f
C460 VTAIL.n220 B 0.023773f
C461 VTAIL.n221 B 0.012775f
C462 VTAIL.n222 B 0.013526f
C463 VTAIL.n223 B 0.030195f
C464 VTAIL.n224 B 0.06877f
C465 VTAIL.n225 B 0.013526f
C466 VTAIL.n226 B 0.012775f
C467 VTAIL.n227 B 0.056249f
C468 VTAIL.n228 B 0.038869f
C469 VTAIL.n229 B 1.72544f
C470 VTAIL.n230 B 0.03534f
C471 VTAIL.n231 B 0.023773f
C472 VTAIL.n232 B 0.012775f
C473 VTAIL.n233 B 0.030195f
C474 VTAIL.n234 B 0.013526f
C475 VTAIL.n235 B 0.023773f
C476 VTAIL.n236 B 0.012775f
C477 VTAIL.n237 B 0.030195f
C478 VTAIL.n238 B 0.013526f
C479 VTAIL.n239 B 0.023773f
C480 VTAIL.n240 B 0.012775f
C481 VTAIL.n241 B 0.030195f
C482 VTAIL.n242 B 0.01315f
C483 VTAIL.n243 B 0.023773f
C484 VTAIL.n244 B 0.013526f
C485 VTAIL.n245 B 0.030195f
C486 VTAIL.n246 B 0.013526f
C487 VTAIL.n247 B 0.023773f
C488 VTAIL.n248 B 0.012775f
C489 VTAIL.n249 B 0.030195f
C490 VTAIL.n250 B 0.013526f
C491 VTAIL.n251 B 1.36849f
C492 VTAIL.n252 B 0.012775f
C493 VTAIL.t9 B 0.051201f
C494 VTAIL.n253 B 0.186003f
C495 VTAIL.n254 B 0.021345f
C496 VTAIL.n255 B 0.022646f
C497 VTAIL.n256 B 0.030195f
C498 VTAIL.n257 B 0.013526f
C499 VTAIL.n258 B 0.012775f
C500 VTAIL.n259 B 0.023773f
C501 VTAIL.n260 B 0.023773f
C502 VTAIL.n261 B 0.012775f
C503 VTAIL.n262 B 0.013526f
C504 VTAIL.n263 B 0.030195f
C505 VTAIL.n264 B 0.030195f
C506 VTAIL.n265 B 0.013526f
C507 VTAIL.n266 B 0.012775f
C508 VTAIL.n267 B 0.023773f
C509 VTAIL.n268 B 0.023773f
C510 VTAIL.n269 B 0.012775f
C511 VTAIL.n270 B 0.012775f
C512 VTAIL.n271 B 0.013526f
C513 VTAIL.n272 B 0.030195f
C514 VTAIL.n273 B 0.030195f
C515 VTAIL.n274 B 0.030195f
C516 VTAIL.n275 B 0.01315f
C517 VTAIL.n276 B 0.012775f
C518 VTAIL.n277 B 0.023773f
C519 VTAIL.n278 B 0.023773f
C520 VTAIL.n279 B 0.012775f
C521 VTAIL.n280 B 0.013526f
C522 VTAIL.n281 B 0.030195f
C523 VTAIL.n282 B 0.030195f
C524 VTAIL.n283 B 0.013526f
C525 VTAIL.n284 B 0.012775f
C526 VTAIL.n285 B 0.023773f
C527 VTAIL.n286 B 0.023773f
C528 VTAIL.n287 B 0.012775f
C529 VTAIL.n288 B 0.013526f
C530 VTAIL.n289 B 0.030195f
C531 VTAIL.n290 B 0.030195f
C532 VTAIL.n291 B 0.013526f
C533 VTAIL.n292 B 0.012775f
C534 VTAIL.n293 B 0.023773f
C535 VTAIL.n294 B 0.023773f
C536 VTAIL.n295 B 0.012775f
C537 VTAIL.n296 B 0.013526f
C538 VTAIL.n297 B 0.030195f
C539 VTAIL.n298 B 0.06877f
C540 VTAIL.n299 B 0.013526f
C541 VTAIL.n300 B 0.012775f
C542 VTAIL.n301 B 0.056249f
C543 VTAIL.n302 B 0.038869f
C544 VTAIL.n303 B 1.66056f
C545 VDD2.n0 B 0.031565f
C546 VDD2.n1 B 0.021234f
C547 VDD2.n2 B 0.01141f
C548 VDD2.n3 B 0.02697f
C549 VDD2.n4 B 0.012081f
C550 VDD2.n5 B 0.021234f
C551 VDD2.n6 B 0.01141f
C552 VDD2.n7 B 0.02697f
C553 VDD2.n8 B 0.012081f
C554 VDD2.n9 B 0.021234f
C555 VDD2.n10 B 0.01141f
C556 VDD2.n11 B 0.02697f
C557 VDD2.n12 B 0.011746f
C558 VDD2.n13 B 0.021234f
C559 VDD2.n14 B 0.012081f
C560 VDD2.n15 B 0.02697f
C561 VDD2.n16 B 0.012081f
C562 VDD2.n17 B 0.021234f
C563 VDD2.n18 B 0.01141f
C564 VDD2.n19 B 0.02697f
C565 VDD2.n20 B 0.012081f
C566 VDD2.n21 B 1.22233f
C567 VDD2.n22 B 0.01141f
C568 VDD2.t1 B 0.045733f
C569 VDD2.n23 B 0.166138f
C570 VDD2.n24 B 0.019065f
C571 VDD2.n25 B 0.020227f
C572 VDD2.n26 B 0.02697f
C573 VDD2.n27 B 0.012081f
C574 VDD2.n28 B 0.01141f
C575 VDD2.n29 B 0.021234f
C576 VDD2.n30 B 0.021234f
C577 VDD2.n31 B 0.01141f
C578 VDD2.n32 B 0.012081f
C579 VDD2.n33 B 0.02697f
C580 VDD2.n34 B 0.02697f
C581 VDD2.n35 B 0.012081f
C582 VDD2.n36 B 0.01141f
C583 VDD2.n37 B 0.021234f
C584 VDD2.n38 B 0.021234f
C585 VDD2.n39 B 0.01141f
C586 VDD2.n40 B 0.01141f
C587 VDD2.n41 B 0.012081f
C588 VDD2.n42 B 0.02697f
C589 VDD2.n43 B 0.02697f
C590 VDD2.n44 B 0.02697f
C591 VDD2.n45 B 0.011746f
C592 VDD2.n46 B 0.01141f
C593 VDD2.n47 B 0.021234f
C594 VDD2.n48 B 0.021234f
C595 VDD2.n49 B 0.01141f
C596 VDD2.n50 B 0.012081f
C597 VDD2.n51 B 0.02697f
C598 VDD2.n52 B 0.02697f
C599 VDD2.n53 B 0.012081f
C600 VDD2.n54 B 0.01141f
C601 VDD2.n55 B 0.021234f
C602 VDD2.n56 B 0.021234f
C603 VDD2.n57 B 0.01141f
C604 VDD2.n58 B 0.012081f
C605 VDD2.n59 B 0.02697f
C606 VDD2.n60 B 0.02697f
C607 VDD2.n61 B 0.012081f
C608 VDD2.n62 B 0.01141f
C609 VDD2.n63 B 0.021234f
C610 VDD2.n64 B 0.021234f
C611 VDD2.n65 B 0.01141f
C612 VDD2.n66 B 0.012081f
C613 VDD2.n67 B 0.02697f
C614 VDD2.n68 B 0.061425f
C615 VDD2.n69 B 0.012081f
C616 VDD2.n70 B 0.01141f
C617 VDD2.n71 B 0.050242f
C618 VDD2.n72 B 0.058262f
C619 VDD2.t4 B 0.228204f
C620 VDD2.t2 B 0.228204f
C621 VDD2.n73 B 2.05375f
C622 VDD2.n74 B 2.62934f
C623 VDD2.n75 B 0.031565f
C624 VDD2.n76 B 0.021234f
C625 VDD2.n77 B 0.01141f
C626 VDD2.n78 B 0.02697f
C627 VDD2.n79 B 0.012081f
C628 VDD2.n80 B 0.021234f
C629 VDD2.n81 B 0.01141f
C630 VDD2.n82 B 0.02697f
C631 VDD2.n83 B 0.012081f
C632 VDD2.n84 B 0.021234f
C633 VDD2.n85 B 0.01141f
C634 VDD2.n86 B 0.02697f
C635 VDD2.n87 B 0.011746f
C636 VDD2.n88 B 0.021234f
C637 VDD2.n89 B 0.011746f
C638 VDD2.n90 B 0.01141f
C639 VDD2.n91 B 0.02697f
C640 VDD2.n92 B 0.02697f
C641 VDD2.n93 B 0.012081f
C642 VDD2.n94 B 0.021234f
C643 VDD2.n95 B 0.01141f
C644 VDD2.n96 B 0.02697f
C645 VDD2.n97 B 0.012081f
C646 VDD2.n98 B 1.22233f
C647 VDD2.n99 B 0.01141f
C648 VDD2.t5 B 0.045733f
C649 VDD2.n100 B 0.166138f
C650 VDD2.n101 B 0.019065f
C651 VDD2.n102 B 0.020227f
C652 VDD2.n103 B 0.02697f
C653 VDD2.n104 B 0.012081f
C654 VDD2.n105 B 0.01141f
C655 VDD2.n106 B 0.021234f
C656 VDD2.n107 B 0.021234f
C657 VDD2.n108 B 0.01141f
C658 VDD2.n109 B 0.012081f
C659 VDD2.n110 B 0.02697f
C660 VDD2.n111 B 0.02697f
C661 VDD2.n112 B 0.012081f
C662 VDD2.n113 B 0.01141f
C663 VDD2.n114 B 0.021234f
C664 VDD2.n115 B 0.021234f
C665 VDD2.n116 B 0.01141f
C666 VDD2.n117 B 0.012081f
C667 VDD2.n118 B 0.02697f
C668 VDD2.n119 B 0.02697f
C669 VDD2.n120 B 0.012081f
C670 VDD2.n121 B 0.01141f
C671 VDD2.n122 B 0.021234f
C672 VDD2.n123 B 0.021234f
C673 VDD2.n124 B 0.01141f
C674 VDD2.n125 B 0.012081f
C675 VDD2.n126 B 0.02697f
C676 VDD2.n127 B 0.02697f
C677 VDD2.n128 B 0.012081f
C678 VDD2.n129 B 0.01141f
C679 VDD2.n130 B 0.021234f
C680 VDD2.n131 B 0.021234f
C681 VDD2.n132 B 0.01141f
C682 VDD2.n133 B 0.012081f
C683 VDD2.n134 B 0.02697f
C684 VDD2.n135 B 0.02697f
C685 VDD2.n136 B 0.012081f
C686 VDD2.n137 B 0.01141f
C687 VDD2.n138 B 0.021234f
C688 VDD2.n139 B 0.021234f
C689 VDD2.n140 B 0.01141f
C690 VDD2.n141 B 0.012081f
C691 VDD2.n142 B 0.02697f
C692 VDD2.n143 B 0.061425f
C693 VDD2.n144 B 0.012081f
C694 VDD2.n145 B 0.01141f
C695 VDD2.n146 B 0.050242f
C696 VDD2.n147 B 0.04937f
C697 VDD2.n148 B 2.44987f
C698 VDD2.t3 B 0.228204f
C699 VDD2.t0 B 0.228204f
C700 VDD2.n149 B 2.05372f
C701 VN.t2 B 2.4136f
C702 VN.n0 B 0.911617f
C703 VN.n1 B 0.019495f
C704 VN.n2 B 0.024024f
C705 VN.n3 B 0.019495f
C706 VN.t5 B 2.4136f
C707 VN.n4 B 0.918477f
C708 VN.t4 B 2.66092f
C709 VN.n5 B 0.869453f
C710 VN.n6 B 0.237372f
C711 VN.n7 B 0.036151f
C712 VN.n8 B 0.036151f
C713 VN.n9 B 0.032654f
C714 VN.n10 B 0.019495f
C715 VN.n11 B 0.019495f
C716 VN.n12 B 0.019495f
C717 VN.n13 B 0.036151f
C718 VN.n14 B 0.036151f
C719 VN.n15 B 0.024015f
C720 VN.n16 B 0.031459f
C721 VN.n17 B 0.052078f
C722 VN.t3 B 2.4136f
C723 VN.n18 B 0.911617f
C724 VN.n19 B 0.019495f
C725 VN.n20 B 0.024024f
C726 VN.n21 B 0.019495f
C727 VN.t0 B 2.4136f
C728 VN.n22 B 0.918477f
C729 VN.t1 B 2.66092f
C730 VN.n23 B 0.869453f
C731 VN.n24 B 0.237372f
C732 VN.n25 B 0.036151f
C733 VN.n26 B 0.036151f
C734 VN.n27 B 0.032654f
C735 VN.n28 B 0.019495f
C736 VN.n29 B 0.019495f
C737 VN.n30 B 0.019495f
C738 VN.n31 B 0.036151f
C739 VN.n32 B 0.036151f
C740 VN.n33 B 0.024015f
C741 VN.n34 B 0.031459f
C742 VN.n35 B 1.20821f
.ends

