* NGSPICE file created from diff_pair_sample_1129.ext - technology: sky130A

.subckt diff_pair_sample_1129 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=5.2494 ps=27.7 w=13.46 l=0.45
X1 VTAIL.t15 VN.t1 VDD2.t6 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X2 VDD2.t5 VN.t2 VTAIL.t9 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X3 B.t11 B.t9 B.t10 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=0 ps=0 w=13.46 l=0.45
X4 VTAIL.t14 VN.t3 VDD2.t4 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=2.2209 ps=13.79 w=13.46 l=0.45
X5 VTAIL.t6 VP.t0 VDD1.t7 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=2.2209 ps=13.79 w=13.46 l=0.45
X6 VTAIL.t13 VN.t4 VDD2.t3 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=2.2209 ps=13.79 w=13.46 l=0.45
X7 B.t8 B.t6 B.t7 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=0 ps=0 w=13.46 l=0.45
X8 VDD2.t2 VN.t5 VTAIL.t12 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=5.2494 ps=27.7 w=13.46 l=0.45
X9 VTAIL.t1 VP.t1 VDD1.t6 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X10 B.t5 B.t3 B.t4 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=0 ps=0 w=13.46 l=0.45
X11 VDD2.t1 VN.t6 VTAIL.t10 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X12 VTAIL.t5 VP.t2 VDD1.t5 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=2.2209 ps=13.79 w=13.46 l=0.45
X13 VTAIL.t4 VP.t3 VDD1.t4 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X14 VDD1.t3 VP.t4 VTAIL.t2 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X15 VDD1.t2 VP.t5 VTAIL.t3 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X16 VDD1.t1 VP.t6 VTAIL.t7 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=5.2494 ps=27.7 w=13.46 l=0.45
X17 B.t2 B.t0 B.t1 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=5.2494 pd=27.7 as=0 ps=0 w=13.46 l=0.45
X18 VTAIL.t8 VN.t7 VDD2.t0 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=2.2209 ps=13.79 w=13.46 l=0.45
X19 VDD1.t0 VP.t7 VTAIL.t0 w_n1750_n3660# sky130_fd_pr__pfet_01v8 ad=2.2209 pd=13.79 as=5.2494 ps=27.7 w=13.46 l=0.45
R0 VN.n2 VN.t3 830.207
R1 VN.n10 VN.t5 830.207
R2 VN.n1 VN.t2 809.225
R3 VN.n5 VN.t1 809.225
R4 VN.n6 VN.t0 809.225
R5 VN.n9 VN.t7 809.225
R6 VN.n13 VN.t6 809.225
R7 VN.n14 VN.t4 809.225
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n11 VN.n10 70.4033
R15 VN.n3 VN.n2 70.4033
R16 VN.n6 VN.n5 48.2005
R17 VN.n14 VN.n13 48.2005
R18 VN VN.n15 42.3433
R19 VN.n4 VN.n1 24.1005
R20 VN.n5 VN.n4 24.1005
R21 VN.n13 VN.n12 24.1005
R22 VN.n12 VN.n9 24.1005
R23 VN.n10 VN.n9 20.9576
R24 VN.n2 VN.n1 20.9576
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VTAIL.n594 VTAIL.n526 756.745
R31 VTAIL.n70 VTAIL.n2 756.745
R32 VTAIL.n144 VTAIL.n76 756.745
R33 VTAIL.n220 VTAIL.n152 756.745
R34 VTAIL.n520 VTAIL.n452 756.745
R35 VTAIL.n444 VTAIL.n376 756.745
R36 VTAIL.n370 VTAIL.n302 756.745
R37 VTAIL.n294 VTAIL.n226 756.745
R38 VTAIL.n551 VTAIL.n550 585
R39 VTAIL.n553 VTAIL.n552 585
R40 VTAIL.n546 VTAIL.n545 585
R41 VTAIL.n559 VTAIL.n558 585
R42 VTAIL.n561 VTAIL.n560 585
R43 VTAIL.n542 VTAIL.n541 585
R44 VTAIL.n568 VTAIL.n567 585
R45 VTAIL.n569 VTAIL.n540 585
R46 VTAIL.n571 VTAIL.n570 585
R47 VTAIL.n538 VTAIL.n537 585
R48 VTAIL.n577 VTAIL.n576 585
R49 VTAIL.n579 VTAIL.n578 585
R50 VTAIL.n534 VTAIL.n533 585
R51 VTAIL.n585 VTAIL.n584 585
R52 VTAIL.n587 VTAIL.n586 585
R53 VTAIL.n530 VTAIL.n529 585
R54 VTAIL.n593 VTAIL.n592 585
R55 VTAIL.n595 VTAIL.n594 585
R56 VTAIL.n27 VTAIL.n26 585
R57 VTAIL.n29 VTAIL.n28 585
R58 VTAIL.n22 VTAIL.n21 585
R59 VTAIL.n35 VTAIL.n34 585
R60 VTAIL.n37 VTAIL.n36 585
R61 VTAIL.n18 VTAIL.n17 585
R62 VTAIL.n44 VTAIL.n43 585
R63 VTAIL.n45 VTAIL.n16 585
R64 VTAIL.n47 VTAIL.n46 585
R65 VTAIL.n14 VTAIL.n13 585
R66 VTAIL.n53 VTAIL.n52 585
R67 VTAIL.n55 VTAIL.n54 585
R68 VTAIL.n10 VTAIL.n9 585
R69 VTAIL.n61 VTAIL.n60 585
R70 VTAIL.n63 VTAIL.n62 585
R71 VTAIL.n6 VTAIL.n5 585
R72 VTAIL.n69 VTAIL.n68 585
R73 VTAIL.n71 VTAIL.n70 585
R74 VTAIL.n101 VTAIL.n100 585
R75 VTAIL.n103 VTAIL.n102 585
R76 VTAIL.n96 VTAIL.n95 585
R77 VTAIL.n109 VTAIL.n108 585
R78 VTAIL.n111 VTAIL.n110 585
R79 VTAIL.n92 VTAIL.n91 585
R80 VTAIL.n118 VTAIL.n117 585
R81 VTAIL.n119 VTAIL.n90 585
R82 VTAIL.n121 VTAIL.n120 585
R83 VTAIL.n88 VTAIL.n87 585
R84 VTAIL.n127 VTAIL.n126 585
R85 VTAIL.n129 VTAIL.n128 585
R86 VTAIL.n84 VTAIL.n83 585
R87 VTAIL.n135 VTAIL.n134 585
R88 VTAIL.n137 VTAIL.n136 585
R89 VTAIL.n80 VTAIL.n79 585
R90 VTAIL.n143 VTAIL.n142 585
R91 VTAIL.n145 VTAIL.n144 585
R92 VTAIL.n177 VTAIL.n176 585
R93 VTAIL.n179 VTAIL.n178 585
R94 VTAIL.n172 VTAIL.n171 585
R95 VTAIL.n185 VTAIL.n184 585
R96 VTAIL.n187 VTAIL.n186 585
R97 VTAIL.n168 VTAIL.n167 585
R98 VTAIL.n194 VTAIL.n193 585
R99 VTAIL.n195 VTAIL.n166 585
R100 VTAIL.n197 VTAIL.n196 585
R101 VTAIL.n164 VTAIL.n163 585
R102 VTAIL.n203 VTAIL.n202 585
R103 VTAIL.n205 VTAIL.n204 585
R104 VTAIL.n160 VTAIL.n159 585
R105 VTAIL.n211 VTAIL.n210 585
R106 VTAIL.n213 VTAIL.n212 585
R107 VTAIL.n156 VTAIL.n155 585
R108 VTAIL.n219 VTAIL.n218 585
R109 VTAIL.n221 VTAIL.n220 585
R110 VTAIL.n521 VTAIL.n520 585
R111 VTAIL.n519 VTAIL.n518 585
R112 VTAIL.n456 VTAIL.n455 585
R113 VTAIL.n513 VTAIL.n512 585
R114 VTAIL.n511 VTAIL.n510 585
R115 VTAIL.n460 VTAIL.n459 585
R116 VTAIL.n505 VTAIL.n504 585
R117 VTAIL.n503 VTAIL.n502 585
R118 VTAIL.n464 VTAIL.n463 585
R119 VTAIL.n468 VTAIL.n466 585
R120 VTAIL.n497 VTAIL.n496 585
R121 VTAIL.n495 VTAIL.n494 585
R122 VTAIL.n470 VTAIL.n469 585
R123 VTAIL.n489 VTAIL.n488 585
R124 VTAIL.n487 VTAIL.n486 585
R125 VTAIL.n474 VTAIL.n473 585
R126 VTAIL.n481 VTAIL.n480 585
R127 VTAIL.n479 VTAIL.n478 585
R128 VTAIL.n445 VTAIL.n444 585
R129 VTAIL.n443 VTAIL.n442 585
R130 VTAIL.n380 VTAIL.n379 585
R131 VTAIL.n437 VTAIL.n436 585
R132 VTAIL.n435 VTAIL.n434 585
R133 VTAIL.n384 VTAIL.n383 585
R134 VTAIL.n429 VTAIL.n428 585
R135 VTAIL.n427 VTAIL.n426 585
R136 VTAIL.n388 VTAIL.n387 585
R137 VTAIL.n392 VTAIL.n390 585
R138 VTAIL.n421 VTAIL.n420 585
R139 VTAIL.n419 VTAIL.n418 585
R140 VTAIL.n394 VTAIL.n393 585
R141 VTAIL.n413 VTAIL.n412 585
R142 VTAIL.n411 VTAIL.n410 585
R143 VTAIL.n398 VTAIL.n397 585
R144 VTAIL.n405 VTAIL.n404 585
R145 VTAIL.n403 VTAIL.n402 585
R146 VTAIL.n371 VTAIL.n370 585
R147 VTAIL.n369 VTAIL.n368 585
R148 VTAIL.n306 VTAIL.n305 585
R149 VTAIL.n363 VTAIL.n362 585
R150 VTAIL.n361 VTAIL.n360 585
R151 VTAIL.n310 VTAIL.n309 585
R152 VTAIL.n355 VTAIL.n354 585
R153 VTAIL.n353 VTAIL.n352 585
R154 VTAIL.n314 VTAIL.n313 585
R155 VTAIL.n318 VTAIL.n316 585
R156 VTAIL.n347 VTAIL.n346 585
R157 VTAIL.n345 VTAIL.n344 585
R158 VTAIL.n320 VTAIL.n319 585
R159 VTAIL.n339 VTAIL.n338 585
R160 VTAIL.n337 VTAIL.n336 585
R161 VTAIL.n324 VTAIL.n323 585
R162 VTAIL.n331 VTAIL.n330 585
R163 VTAIL.n329 VTAIL.n328 585
R164 VTAIL.n295 VTAIL.n294 585
R165 VTAIL.n293 VTAIL.n292 585
R166 VTAIL.n230 VTAIL.n229 585
R167 VTAIL.n287 VTAIL.n286 585
R168 VTAIL.n285 VTAIL.n284 585
R169 VTAIL.n234 VTAIL.n233 585
R170 VTAIL.n279 VTAIL.n278 585
R171 VTAIL.n277 VTAIL.n276 585
R172 VTAIL.n238 VTAIL.n237 585
R173 VTAIL.n242 VTAIL.n240 585
R174 VTAIL.n271 VTAIL.n270 585
R175 VTAIL.n269 VTAIL.n268 585
R176 VTAIL.n244 VTAIL.n243 585
R177 VTAIL.n263 VTAIL.n262 585
R178 VTAIL.n261 VTAIL.n260 585
R179 VTAIL.n248 VTAIL.n247 585
R180 VTAIL.n255 VTAIL.n254 585
R181 VTAIL.n253 VTAIL.n252 585
R182 VTAIL.n549 VTAIL.t11 329.036
R183 VTAIL.n25 VTAIL.t14 329.036
R184 VTAIL.n99 VTAIL.t7 329.036
R185 VTAIL.n175 VTAIL.t5 329.036
R186 VTAIL.n477 VTAIL.t0 329.036
R187 VTAIL.n401 VTAIL.t6 329.036
R188 VTAIL.n327 VTAIL.t12 329.036
R189 VTAIL.n251 VTAIL.t13 329.036
R190 VTAIL.n552 VTAIL.n551 171.744
R191 VTAIL.n552 VTAIL.n545 171.744
R192 VTAIL.n559 VTAIL.n545 171.744
R193 VTAIL.n560 VTAIL.n559 171.744
R194 VTAIL.n560 VTAIL.n541 171.744
R195 VTAIL.n568 VTAIL.n541 171.744
R196 VTAIL.n569 VTAIL.n568 171.744
R197 VTAIL.n570 VTAIL.n569 171.744
R198 VTAIL.n570 VTAIL.n537 171.744
R199 VTAIL.n577 VTAIL.n537 171.744
R200 VTAIL.n578 VTAIL.n577 171.744
R201 VTAIL.n578 VTAIL.n533 171.744
R202 VTAIL.n585 VTAIL.n533 171.744
R203 VTAIL.n586 VTAIL.n585 171.744
R204 VTAIL.n586 VTAIL.n529 171.744
R205 VTAIL.n593 VTAIL.n529 171.744
R206 VTAIL.n594 VTAIL.n593 171.744
R207 VTAIL.n28 VTAIL.n27 171.744
R208 VTAIL.n28 VTAIL.n21 171.744
R209 VTAIL.n35 VTAIL.n21 171.744
R210 VTAIL.n36 VTAIL.n35 171.744
R211 VTAIL.n36 VTAIL.n17 171.744
R212 VTAIL.n44 VTAIL.n17 171.744
R213 VTAIL.n45 VTAIL.n44 171.744
R214 VTAIL.n46 VTAIL.n45 171.744
R215 VTAIL.n46 VTAIL.n13 171.744
R216 VTAIL.n53 VTAIL.n13 171.744
R217 VTAIL.n54 VTAIL.n53 171.744
R218 VTAIL.n54 VTAIL.n9 171.744
R219 VTAIL.n61 VTAIL.n9 171.744
R220 VTAIL.n62 VTAIL.n61 171.744
R221 VTAIL.n62 VTAIL.n5 171.744
R222 VTAIL.n69 VTAIL.n5 171.744
R223 VTAIL.n70 VTAIL.n69 171.744
R224 VTAIL.n102 VTAIL.n101 171.744
R225 VTAIL.n102 VTAIL.n95 171.744
R226 VTAIL.n109 VTAIL.n95 171.744
R227 VTAIL.n110 VTAIL.n109 171.744
R228 VTAIL.n110 VTAIL.n91 171.744
R229 VTAIL.n118 VTAIL.n91 171.744
R230 VTAIL.n119 VTAIL.n118 171.744
R231 VTAIL.n120 VTAIL.n119 171.744
R232 VTAIL.n120 VTAIL.n87 171.744
R233 VTAIL.n127 VTAIL.n87 171.744
R234 VTAIL.n128 VTAIL.n127 171.744
R235 VTAIL.n128 VTAIL.n83 171.744
R236 VTAIL.n135 VTAIL.n83 171.744
R237 VTAIL.n136 VTAIL.n135 171.744
R238 VTAIL.n136 VTAIL.n79 171.744
R239 VTAIL.n143 VTAIL.n79 171.744
R240 VTAIL.n144 VTAIL.n143 171.744
R241 VTAIL.n178 VTAIL.n177 171.744
R242 VTAIL.n178 VTAIL.n171 171.744
R243 VTAIL.n185 VTAIL.n171 171.744
R244 VTAIL.n186 VTAIL.n185 171.744
R245 VTAIL.n186 VTAIL.n167 171.744
R246 VTAIL.n194 VTAIL.n167 171.744
R247 VTAIL.n195 VTAIL.n194 171.744
R248 VTAIL.n196 VTAIL.n195 171.744
R249 VTAIL.n196 VTAIL.n163 171.744
R250 VTAIL.n203 VTAIL.n163 171.744
R251 VTAIL.n204 VTAIL.n203 171.744
R252 VTAIL.n204 VTAIL.n159 171.744
R253 VTAIL.n211 VTAIL.n159 171.744
R254 VTAIL.n212 VTAIL.n211 171.744
R255 VTAIL.n212 VTAIL.n155 171.744
R256 VTAIL.n219 VTAIL.n155 171.744
R257 VTAIL.n220 VTAIL.n219 171.744
R258 VTAIL.n520 VTAIL.n519 171.744
R259 VTAIL.n519 VTAIL.n455 171.744
R260 VTAIL.n512 VTAIL.n455 171.744
R261 VTAIL.n512 VTAIL.n511 171.744
R262 VTAIL.n511 VTAIL.n459 171.744
R263 VTAIL.n504 VTAIL.n459 171.744
R264 VTAIL.n504 VTAIL.n503 171.744
R265 VTAIL.n503 VTAIL.n463 171.744
R266 VTAIL.n468 VTAIL.n463 171.744
R267 VTAIL.n496 VTAIL.n468 171.744
R268 VTAIL.n496 VTAIL.n495 171.744
R269 VTAIL.n495 VTAIL.n469 171.744
R270 VTAIL.n488 VTAIL.n469 171.744
R271 VTAIL.n488 VTAIL.n487 171.744
R272 VTAIL.n487 VTAIL.n473 171.744
R273 VTAIL.n480 VTAIL.n473 171.744
R274 VTAIL.n480 VTAIL.n479 171.744
R275 VTAIL.n444 VTAIL.n443 171.744
R276 VTAIL.n443 VTAIL.n379 171.744
R277 VTAIL.n436 VTAIL.n379 171.744
R278 VTAIL.n436 VTAIL.n435 171.744
R279 VTAIL.n435 VTAIL.n383 171.744
R280 VTAIL.n428 VTAIL.n383 171.744
R281 VTAIL.n428 VTAIL.n427 171.744
R282 VTAIL.n427 VTAIL.n387 171.744
R283 VTAIL.n392 VTAIL.n387 171.744
R284 VTAIL.n420 VTAIL.n392 171.744
R285 VTAIL.n420 VTAIL.n419 171.744
R286 VTAIL.n419 VTAIL.n393 171.744
R287 VTAIL.n412 VTAIL.n393 171.744
R288 VTAIL.n412 VTAIL.n411 171.744
R289 VTAIL.n411 VTAIL.n397 171.744
R290 VTAIL.n404 VTAIL.n397 171.744
R291 VTAIL.n404 VTAIL.n403 171.744
R292 VTAIL.n370 VTAIL.n369 171.744
R293 VTAIL.n369 VTAIL.n305 171.744
R294 VTAIL.n362 VTAIL.n305 171.744
R295 VTAIL.n362 VTAIL.n361 171.744
R296 VTAIL.n361 VTAIL.n309 171.744
R297 VTAIL.n354 VTAIL.n309 171.744
R298 VTAIL.n354 VTAIL.n353 171.744
R299 VTAIL.n353 VTAIL.n313 171.744
R300 VTAIL.n318 VTAIL.n313 171.744
R301 VTAIL.n346 VTAIL.n318 171.744
R302 VTAIL.n346 VTAIL.n345 171.744
R303 VTAIL.n345 VTAIL.n319 171.744
R304 VTAIL.n338 VTAIL.n319 171.744
R305 VTAIL.n338 VTAIL.n337 171.744
R306 VTAIL.n337 VTAIL.n323 171.744
R307 VTAIL.n330 VTAIL.n323 171.744
R308 VTAIL.n330 VTAIL.n329 171.744
R309 VTAIL.n294 VTAIL.n293 171.744
R310 VTAIL.n293 VTAIL.n229 171.744
R311 VTAIL.n286 VTAIL.n229 171.744
R312 VTAIL.n286 VTAIL.n285 171.744
R313 VTAIL.n285 VTAIL.n233 171.744
R314 VTAIL.n278 VTAIL.n233 171.744
R315 VTAIL.n278 VTAIL.n277 171.744
R316 VTAIL.n277 VTAIL.n237 171.744
R317 VTAIL.n242 VTAIL.n237 171.744
R318 VTAIL.n270 VTAIL.n242 171.744
R319 VTAIL.n270 VTAIL.n269 171.744
R320 VTAIL.n269 VTAIL.n243 171.744
R321 VTAIL.n262 VTAIL.n243 171.744
R322 VTAIL.n262 VTAIL.n261 171.744
R323 VTAIL.n261 VTAIL.n247 171.744
R324 VTAIL.n254 VTAIL.n247 171.744
R325 VTAIL.n254 VTAIL.n253 171.744
R326 VTAIL.n551 VTAIL.t11 85.8723
R327 VTAIL.n27 VTAIL.t14 85.8723
R328 VTAIL.n101 VTAIL.t7 85.8723
R329 VTAIL.n177 VTAIL.t5 85.8723
R330 VTAIL.n479 VTAIL.t0 85.8723
R331 VTAIL.n403 VTAIL.t6 85.8723
R332 VTAIL.n329 VTAIL.t12 85.8723
R333 VTAIL.n253 VTAIL.t13 85.8723
R334 VTAIL.n451 VTAIL.n450 53.6627
R335 VTAIL.n301 VTAIL.n300 53.6627
R336 VTAIL.n1 VTAIL.n0 53.6625
R337 VTAIL.n151 VTAIL.n150 53.6625
R338 VTAIL.n599 VTAIL.n598 30.246
R339 VTAIL.n75 VTAIL.n74 30.246
R340 VTAIL.n149 VTAIL.n148 30.246
R341 VTAIL.n225 VTAIL.n224 30.246
R342 VTAIL.n525 VTAIL.n524 30.246
R343 VTAIL.n449 VTAIL.n448 30.246
R344 VTAIL.n375 VTAIL.n374 30.246
R345 VTAIL.n299 VTAIL.n298 30.246
R346 VTAIL.n599 VTAIL.n525 24.6427
R347 VTAIL.n299 VTAIL.n225 24.6427
R348 VTAIL.n571 VTAIL.n538 13.1884
R349 VTAIL.n47 VTAIL.n14 13.1884
R350 VTAIL.n121 VTAIL.n88 13.1884
R351 VTAIL.n197 VTAIL.n164 13.1884
R352 VTAIL.n466 VTAIL.n464 13.1884
R353 VTAIL.n390 VTAIL.n388 13.1884
R354 VTAIL.n316 VTAIL.n314 13.1884
R355 VTAIL.n240 VTAIL.n238 13.1884
R356 VTAIL.n572 VTAIL.n540 12.8005
R357 VTAIL.n576 VTAIL.n575 12.8005
R358 VTAIL.n48 VTAIL.n16 12.8005
R359 VTAIL.n52 VTAIL.n51 12.8005
R360 VTAIL.n122 VTAIL.n90 12.8005
R361 VTAIL.n126 VTAIL.n125 12.8005
R362 VTAIL.n198 VTAIL.n166 12.8005
R363 VTAIL.n202 VTAIL.n201 12.8005
R364 VTAIL.n502 VTAIL.n501 12.8005
R365 VTAIL.n498 VTAIL.n497 12.8005
R366 VTAIL.n426 VTAIL.n425 12.8005
R367 VTAIL.n422 VTAIL.n421 12.8005
R368 VTAIL.n352 VTAIL.n351 12.8005
R369 VTAIL.n348 VTAIL.n347 12.8005
R370 VTAIL.n276 VTAIL.n275 12.8005
R371 VTAIL.n272 VTAIL.n271 12.8005
R372 VTAIL.n567 VTAIL.n566 12.0247
R373 VTAIL.n579 VTAIL.n536 12.0247
R374 VTAIL.n43 VTAIL.n42 12.0247
R375 VTAIL.n55 VTAIL.n12 12.0247
R376 VTAIL.n117 VTAIL.n116 12.0247
R377 VTAIL.n129 VTAIL.n86 12.0247
R378 VTAIL.n193 VTAIL.n192 12.0247
R379 VTAIL.n205 VTAIL.n162 12.0247
R380 VTAIL.n505 VTAIL.n462 12.0247
R381 VTAIL.n494 VTAIL.n467 12.0247
R382 VTAIL.n429 VTAIL.n386 12.0247
R383 VTAIL.n418 VTAIL.n391 12.0247
R384 VTAIL.n355 VTAIL.n312 12.0247
R385 VTAIL.n344 VTAIL.n317 12.0247
R386 VTAIL.n279 VTAIL.n236 12.0247
R387 VTAIL.n268 VTAIL.n241 12.0247
R388 VTAIL.n565 VTAIL.n542 11.249
R389 VTAIL.n580 VTAIL.n534 11.249
R390 VTAIL.n41 VTAIL.n18 11.249
R391 VTAIL.n56 VTAIL.n10 11.249
R392 VTAIL.n115 VTAIL.n92 11.249
R393 VTAIL.n130 VTAIL.n84 11.249
R394 VTAIL.n191 VTAIL.n168 11.249
R395 VTAIL.n206 VTAIL.n160 11.249
R396 VTAIL.n506 VTAIL.n460 11.249
R397 VTAIL.n493 VTAIL.n470 11.249
R398 VTAIL.n430 VTAIL.n384 11.249
R399 VTAIL.n417 VTAIL.n394 11.249
R400 VTAIL.n356 VTAIL.n310 11.249
R401 VTAIL.n343 VTAIL.n320 11.249
R402 VTAIL.n280 VTAIL.n234 11.249
R403 VTAIL.n267 VTAIL.n244 11.249
R404 VTAIL.n550 VTAIL.n549 10.7239
R405 VTAIL.n26 VTAIL.n25 10.7239
R406 VTAIL.n100 VTAIL.n99 10.7239
R407 VTAIL.n176 VTAIL.n175 10.7239
R408 VTAIL.n478 VTAIL.n477 10.7239
R409 VTAIL.n402 VTAIL.n401 10.7239
R410 VTAIL.n328 VTAIL.n327 10.7239
R411 VTAIL.n252 VTAIL.n251 10.7239
R412 VTAIL.n562 VTAIL.n561 10.4732
R413 VTAIL.n584 VTAIL.n583 10.4732
R414 VTAIL.n38 VTAIL.n37 10.4732
R415 VTAIL.n60 VTAIL.n59 10.4732
R416 VTAIL.n112 VTAIL.n111 10.4732
R417 VTAIL.n134 VTAIL.n133 10.4732
R418 VTAIL.n188 VTAIL.n187 10.4732
R419 VTAIL.n210 VTAIL.n209 10.4732
R420 VTAIL.n510 VTAIL.n509 10.4732
R421 VTAIL.n490 VTAIL.n489 10.4732
R422 VTAIL.n434 VTAIL.n433 10.4732
R423 VTAIL.n414 VTAIL.n413 10.4732
R424 VTAIL.n360 VTAIL.n359 10.4732
R425 VTAIL.n340 VTAIL.n339 10.4732
R426 VTAIL.n284 VTAIL.n283 10.4732
R427 VTAIL.n264 VTAIL.n263 10.4732
R428 VTAIL.n558 VTAIL.n544 9.69747
R429 VTAIL.n587 VTAIL.n532 9.69747
R430 VTAIL.n34 VTAIL.n20 9.69747
R431 VTAIL.n63 VTAIL.n8 9.69747
R432 VTAIL.n108 VTAIL.n94 9.69747
R433 VTAIL.n137 VTAIL.n82 9.69747
R434 VTAIL.n184 VTAIL.n170 9.69747
R435 VTAIL.n213 VTAIL.n158 9.69747
R436 VTAIL.n513 VTAIL.n458 9.69747
R437 VTAIL.n486 VTAIL.n472 9.69747
R438 VTAIL.n437 VTAIL.n382 9.69747
R439 VTAIL.n410 VTAIL.n396 9.69747
R440 VTAIL.n363 VTAIL.n308 9.69747
R441 VTAIL.n336 VTAIL.n322 9.69747
R442 VTAIL.n287 VTAIL.n232 9.69747
R443 VTAIL.n260 VTAIL.n246 9.69747
R444 VTAIL.n598 VTAIL.n597 9.45567
R445 VTAIL.n74 VTAIL.n73 9.45567
R446 VTAIL.n148 VTAIL.n147 9.45567
R447 VTAIL.n224 VTAIL.n223 9.45567
R448 VTAIL.n524 VTAIL.n523 9.45567
R449 VTAIL.n448 VTAIL.n447 9.45567
R450 VTAIL.n374 VTAIL.n373 9.45567
R451 VTAIL.n298 VTAIL.n297 9.45567
R452 VTAIL.n597 VTAIL.n596 9.3005
R453 VTAIL.n591 VTAIL.n590 9.3005
R454 VTAIL.n589 VTAIL.n588 9.3005
R455 VTAIL.n532 VTAIL.n531 9.3005
R456 VTAIL.n583 VTAIL.n582 9.3005
R457 VTAIL.n581 VTAIL.n580 9.3005
R458 VTAIL.n536 VTAIL.n535 9.3005
R459 VTAIL.n575 VTAIL.n574 9.3005
R460 VTAIL.n548 VTAIL.n547 9.3005
R461 VTAIL.n555 VTAIL.n554 9.3005
R462 VTAIL.n557 VTAIL.n556 9.3005
R463 VTAIL.n544 VTAIL.n543 9.3005
R464 VTAIL.n563 VTAIL.n562 9.3005
R465 VTAIL.n565 VTAIL.n564 9.3005
R466 VTAIL.n566 VTAIL.n539 9.3005
R467 VTAIL.n573 VTAIL.n572 9.3005
R468 VTAIL.n528 VTAIL.n527 9.3005
R469 VTAIL.n73 VTAIL.n72 9.3005
R470 VTAIL.n67 VTAIL.n66 9.3005
R471 VTAIL.n65 VTAIL.n64 9.3005
R472 VTAIL.n8 VTAIL.n7 9.3005
R473 VTAIL.n59 VTAIL.n58 9.3005
R474 VTAIL.n57 VTAIL.n56 9.3005
R475 VTAIL.n12 VTAIL.n11 9.3005
R476 VTAIL.n51 VTAIL.n50 9.3005
R477 VTAIL.n24 VTAIL.n23 9.3005
R478 VTAIL.n31 VTAIL.n30 9.3005
R479 VTAIL.n33 VTAIL.n32 9.3005
R480 VTAIL.n20 VTAIL.n19 9.3005
R481 VTAIL.n39 VTAIL.n38 9.3005
R482 VTAIL.n41 VTAIL.n40 9.3005
R483 VTAIL.n42 VTAIL.n15 9.3005
R484 VTAIL.n49 VTAIL.n48 9.3005
R485 VTAIL.n4 VTAIL.n3 9.3005
R486 VTAIL.n147 VTAIL.n146 9.3005
R487 VTAIL.n141 VTAIL.n140 9.3005
R488 VTAIL.n139 VTAIL.n138 9.3005
R489 VTAIL.n82 VTAIL.n81 9.3005
R490 VTAIL.n133 VTAIL.n132 9.3005
R491 VTAIL.n131 VTAIL.n130 9.3005
R492 VTAIL.n86 VTAIL.n85 9.3005
R493 VTAIL.n125 VTAIL.n124 9.3005
R494 VTAIL.n98 VTAIL.n97 9.3005
R495 VTAIL.n105 VTAIL.n104 9.3005
R496 VTAIL.n107 VTAIL.n106 9.3005
R497 VTAIL.n94 VTAIL.n93 9.3005
R498 VTAIL.n113 VTAIL.n112 9.3005
R499 VTAIL.n115 VTAIL.n114 9.3005
R500 VTAIL.n116 VTAIL.n89 9.3005
R501 VTAIL.n123 VTAIL.n122 9.3005
R502 VTAIL.n78 VTAIL.n77 9.3005
R503 VTAIL.n223 VTAIL.n222 9.3005
R504 VTAIL.n217 VTAIL.n216 9.3005
R505 VTAIL.n215 VTAIL.n214 9.3005
R506 VTAIL.n158 VTAIL.n157 9.3005
R507 VTAIL.n209 VTAIL.n208 9.3005
R508 VTAIL.n207 VTAIL.n206 9.3005
R509 VTAIL.n162 VTAIL.n161 9.3005
R510 VTAIL.n201 VTAIL.n200 9.3005
R511 VTAIL.n174 VTAIL.n173 9.3005
R512 VTAIL.n181 VTAIL.n180 9.3005
R513 VTAIL.n183 VTAIL.n182 9.3005
R514 VTAIL.n170 VTAIL.n169 9.3005
R515 VTAIL.n189 VTAIL.n188 9.3005
R516 VTAIL.n191 VTAIL.n190 9.3005
R517 VTAIL.n192 VTAIL.n165 9.3005
R518 VTAIL.n199 VTAIL.n198 9.3005
R519 VTAIL.n154 VTAIL.n153 9.3005
R520 VTAIL.n476 VTAIL.n475 9.3005
R521 VTAIL.n483 VTAIL.n482 9.3005
R522 VTAIL.n485 VTAIL.n484 9.3005
R523 VTAIL.n472 VTAIL.n471 9.3005
R524 VTAIL.n491 VTAIL.n490 9.3005
R525 VTAIL.n493 VTAIL.n492 9.3005
R526 VTAIL.n467 VTAIL.n465 9.3005
R527 VTAIL.n499 VTAIL.n498 9.3005
R528 VTAIL.n523 VTAIL.n522 9.3005
R529 VTAIL.n454 VTAIL.n453 9.3005
R530 VTAIL.n517 VTAIL.n516 9.3005
R531 VTAIL.n515 VTAIL.n514 9.3005
R532 VTAIL.n458 VTAIL.n457 9.3005
R533 VTAIL.n509 VTAIL.n508 9.3005
R534 VTAIL.n507 VTAIL.n506 9.3005
R535 VTAIL.n462 VTAIL.n461 9.3005
R536 VTAIL.n501 VTAIL.n500 9.3005
R537 VTAIL.n400 VTAIL.n399 9.3005
R538 VTAIL.n407 VTAIL.n406 9.3005
R539 VTAIL.n409 VTAIL.n408 9.3005
R540 VTAIL.n396 VTAIL.n395 9.3005
R541 VTAIL.n415 VTAIL.n414 9.3005
R542 VTAIL.n417 VTAIL.n416 9.3005
R543 VTAIL.n391 VTAIL.n389 9.3005
R544 VTAIL.n423 VTAIL.n422 9.3005
R545 VTAIL.n447 VTAIL.n446 9.3005
R546 VTAIL.n378 VTAIL.n377 9.3005
R547 VTAIL.n441 VTAIL.n440 9.3005
R548 VTAIL.n439 VTAIL.n438 9.3005
R549 VTAIL.n382 VTAIL.n381 9.3005
R550 VTAIL.n433 VTAIL.n432 9.3005
R551 VTAIL.n431 VTAIL.n430 9.3005
R552 VTAIL.n386 VTAIL.n385 9.3005
R553 VTAIL.n425 VTAIL.n424 9.3005
R554 VTAIL.n326 VTAIL.n325 9.3005
R555 VTAIL.n333 VTAIL.n332 9.3005
R556 VTAIL.n335 VTAIL.n334 9.3005
R557 VTAIL.n322 VTAIL.n321 9.3005
R558 VTAIL.n341 VTAIL.n340 9.3005
R559 VTAIL.n343 VTAIL.n342 9.3005
R560 VTAIL.n317 VTAIL.n315 9.3005
R561 VTAIL.n349 VTAIL.n348 9.3005
R562 VTAIL.n373 VTAIL.n372 9.3005
R563 VTAIL.n304 VTAIL.n303 9.3005
R564 VTAIL.n367 VTAIL.n366 9.3005
R565 VTAIL.n365 VTAIL.n364 9.3005
R566 VTAIL.n308 VTAIL.n307 9.3005
R567 VTAIL.n359 VTAIL.n358 9.3005
R568 VTAIL.n357 VTAIL.n356 9.3005
R569 VTAIL.n312 VTAIL.n311 9.3005
R570 VTAIL.n351 VTAIL.n350 9.3005
R571 VTAIL.n250 VTAIL.n249 9.3005
R572 VTAIL.n257 VTAIL.n256 9.3005
R573 VTAIL.n259 VTAIL.n258 9.3005
R574 VTAIL.n246 VTAIL.n245 9.3005
R575 VTAIL.n265 VTAIL.n264 9.3005
R576 VTAIL.n267 VTAIL.n266 9.3005
R577 VTAIL.n241 VTAIL.n239 9.3005
R578 VTAIL.n273 VTAIL.n272 9.3005
R579 VTAIL.n297 VTAIL.n296 9.3005
R580 VTAIL.n228 VTAIL.n227 9.3005
R581 VTAIL.n291 VTAIL.n290 9.3005
R582 VTAIL.n289 VTAIL.n288 9.3005
R583 VTAIL.n232 VTAIL.n231 9.3005
R584 VTAIL.n283 VTAIL.n282 9.3005
R585 VTAIL.n281 VTAIL.n280 9.3005
R586 VTAIL.n236 VTAIL.n235 9.3005
R587 VTAIL.n275 VTAIL.n274 9.3005
R588 VTAIL.n557 VTAIL.n546 8.92171
R589 VTAIL.n588 VTAIL.n530 8.92171
R590 VTAIL.n33 VTAIL.n22 8.92171
R591 VTAIL.n64 VTAIL.n6 8.92171
R592 VTAIL.n107 VTAIL.n96 8.92171
R593 VTAIL.n138 VTAIL.n80 8.92171
R594 VTAIL.n183 VTAIL.n172 8.92171
R595 VTAIL.n214 VTAIL.n156 8.92171
R596 VTAIL.n514 VTAIL.n456 8.92171
R597 VTAIL.n485 VTAIL.n474 8.92171
R598 VTAIL.n438 VTAIL.n380 8.92171
R599 VTAIL.n409 VTAIL.n398 8.92171
R600 VTAIL.n364 VTAIL.n306 8.92171
R601 VTAIL.n335 VTAIL.n324 8.92171
R602 VTAIL.n288 VTAIL.n230 8.92171
R603 VTAIL.n259 VTAIL.n248 8.92171
R604 VTAIL.n554 VTAIL.n553 8.14595
R605 VTAIL.n592 VTAIL.n591 8.14595
R606 VTAIL.n30 VTAIL.n29 8.14595
R607 VTAIL.n68 VTAIL.n67 8.14595
R608 VTAIL.n104 VTAIL.n103 8.14595
R609 VTAIL.n142 VTAIL.n141 8.14595
R610 VTAIL.n180 VTAIL.n179 8.14595
R611 VTAIL.n218 VTAIL.n217 8.14595
R612 VTAIL.n518 VTAIL.n517 8.14595
R613 VTAIL.n482 VTAIL.n481 8.14595
R614 VTAIL.n442 VTAIL.n441 8.14595
R615 VTAIL.n406 VTAIL.n405 8.14595
R616 VTAIL.n368 VTAIL.n367 8.14595
R617 VTAIL.n332 VTAIL.n331 8.14595
R618 VTAIL.n292 VTAIL.n291 8.14595
R619 VTAIL.n256 VTAIL.n255 8.14595
R620 VTAIL.n550 VTAIL.n548 7.3702
R621 VTAIL.n595 VTAIL.n528 7.3702
R622 VTAIL.n598 VTAIL.n526 7.3702
R623 VTAIL.n26 VTAIL.n24 7.3702
R624 VTAIL.n71 VTAIL.n4 7.3702
R625 VTAIL.n74 VTAIL.n2 7.3702
R626 VTAIL.n100 VTAIL.n98 7.3702
R627 VTAIL.n145 VTAIL.n78 7.3702
R628 VTAIL.n148 VTAIL.n76 7.3702
R629 VTAIL.n176 VTAIL.n174 7.3702
R630 VTAIL.n221 VTAIL.n154 7.3702
R631 VTAIL.n224 VTAIL.n152 7.3702
R632 VTAIL.n524 VTAIL.n452 7.3702
R633 VTAIL.n521 VTAIL.n454 7.3702
R634 VTAIL.n478 VTAIL.n476 7.3702
R635 VTAIL.n448 VTAIL.n376 7.3702
R636 VTAIL.n445 VTAIL.n378 7.3702
R637 VTAIL.n402 VTAIL.n400 7.3702
R638 VTAIL.n374 VTAIL.n302 7.3702
R639 VTAIL.n371 VTAIL.n304 7.3702
R640 VTAIL.n328 VTAIL.n326 7.3702
R641 VTAIL.n298 VTAIL.n226 7.3702
R642 VTAIL.n295 VTAIL.n228 7.3702
R643 VTAIL.n252 VTAIL.n250 7.3702
R644 VTAIL.n596 VTAIL.n595 6.59444
R645 VTAIL.n596 VTAIL.n526 6.59444
R646 VTAIL.n72 VTAIL.n71 6.59444
R647 VTAIL.n72 VTAIL.n2 6.59444
R648 VTAIL.n146 VTAIL.n145 6.59444
R649 VTAIL.n146 VTAIL.n76 6.59444
R650 VTAIL.n222 VTAIL.n221 6.59444
R651 VTAIL.n222 VTAIL.n152 6.59444
R652 VTAIL.n522 VTAIL.n452 6.59444
R653 VTAIL.n522 VTAIL.n521 6.59444
R654 VTAIL.n446 VTAIL.n376 6.59444
R655 VTAIL.n446 VTAIL.n445 6.59444
R656 VTAIL.n372 VTAIL.n302 6.59444
R657 VTAIL.n372 VTAIL.n371 6.59444
R658 VTAIL.n296 VTAIL.n226 6.59444
R659 VTAIL.n296 VTAIL.n295 6.59444
R660 VTAIL.n553 VTAIL.n548 5.81868
R661 VTAIL.n592 VTAIL.n528 5.81868
R662 VTAIL.n29 VTAIL.n24 5.81868
R663 VTAIL.n68 VTAIL.n4 5.81868
R664 VTAIL.n103 VTAIL.n98 5.81868
R665 VTAIL.n142 VTAIL.n78 5.81868
R666 VTAIL.n179 VTAIL.n174 5.81868
R667 VTAIL.n218 VTAIL.n154 5.81868
R668 VTAIL.n518 VTAIL.n454 5.81868
R669 VTAIL.n481 VTAIL.n476 5.81868
R670 VTAIL.n442 VTAIL.n378 5.81868
R671 VTAIL.n405 VTAIL.n400 5.81868
R672 VTAIL.n368 VTAIL.n304 5.81868
R673 VTAIL.n331 VTAIL.n326 5.81868
R674 VTAIL.n292 VTAIL.n228 5.81868
R675 VTAIL.n255 VTAIL.n250 5.81868
R676 VTAIL.n554 VTAIL.n546 5.04292
R677 VTAIL.n591 VTAIL.n530 5.04292
R678 VTAIL.n30 VTAIL.n22 5.04292
R679 VTAIL.n67 VTAIL.n6 5.04292
R680 VTAIL.n104 VTAIL.n96 5.04292
R681 VTAIL.n141 VTAIL.n80 5.04292
R682 VTAIL.n180 VTAIL.n172 5.04292
R683 VTAIL.n217 VTAIL.n156 5.04292
R684 VTAIL.n517 VTAIL.n456 5.04292
R685 VTAIL.n482 VTAIL.n474 5.04292
R686 VTAIL.n441 VTAIL.n380 5.04292
R687 VTAIL.n406 VTAIL.n398 5.04292
R688 VTAIL.n367 VTAIL.n306 5.04292
R689 VTAIL.n332 VTAIL.n324 5.04292
R690 VTAIL.n291 VTAIL.n230 5.04292
R691 VTAIL.n256 VTAIL.n248 5.04292
R692 VTAIL.n558 VTAIL.n557 4.26717
R693 VTAIL.n588 VTAIL.n587 4.26717
R694 VTAIL.n34 VTAIL.n33 4.26717
R695 VTAIL.n64 VTAIL.n63 4.26717
R696 VTAIL.n108 VTAIL.n107 4.26717
R697 VTAIL.n138 VTAIL.n137 4.26717
R698 VTAIL.n184 VTAIL.n183 4.26717
R699 VTAIL.n214 VTAIL.n213 4.26717
R700 VTAIL.n514 VTAIL.n513 4.26717
R701 VTAIL.n486 VTAIL.n485 4.26717
R702 VTAIL.n438 VTAIL.n437 4.26717
R703 VTAIL.n410 VTAIL.n409 4.26717
R704 VTAIL.n364 VTAIL.n363 4.26717
R705 VTAIL.n336 VTAIL.n335 4.26717
R706 VTAIL.n288 VTAIL.n287 4.26717
R707 VTAIL.n260 VTAIL.n259 4.26717
R708 VTAIL.n561 VTAIL.n544 3.49141
R709 VTAIL.n584 VTAIL.n532 3.49141
R710 VTAIL.n37 VTAIL.n20 3.49141
R711 VTAIL.n60 VTAIL.n8 3.49141
R712 VTAIL.n111 VTAIL.n94 3.49141
R713 VTAIL.n134 VTAIL.n82 3.49141
R714 VTAIL.n187 VTAIL.n170 3.49141
R715 VTAIL.n210 VTAIL.n158 3.49141
R716 VTAIL.n510 VTAIL.n458 3.49141
R717 VTAIL.n489 VTAIL.n472 3.49141
R718 VTAIL.n434 VTAIL.n382 3.49141
R719 VTAIL.n413 VTAIL.n396 3.49141
R720 VTAIL.n360 VTAIL.n308 3.49141
R721 VTAIL.n339 VTAIL.n322 3.49141
R722 VTAIL.n284 VTAIL.n232 3.49141
R723 VTAIL.n263 VTAIL.n246 3.49141
R724 VTAIL.n562 VTAIL.n542 2.71565
R725 VTAIL.n583 VTAIL.n534 2.71565
R726 VTAIL.n38 VTAIL.n18 2.71565
R727 VTAIL.n59 VTAIL.n10 2.71565
R728 VTAIL.n112 VTAIL.n92 2.71565
R729 VTAIL.n133 VTAIL.n84 2.71565
R730 VTAIL.n188 VTAIL.n168 2.71565
R731 VTAIL.n209 VTAIL.n160 2.71565
R732 VTAIL.n509 VTAIL.n460 2.71565
R733 VTAIL.n490 VTAIL.n470 2.71565
R734 VTAIL.n433 VTAIL.n384 2.71565
R735 VTAIL.n414 VTAIL.n394 2.71565
R736 VTAIL.n359 VTAIL.n310 2.71565
R737 VTAIL.n340 VTAIL.n320 2.71565
R738 VTAIL.n283 VTAIL.n234 2.71565
R739 VTAIL.n264 VTAIL.n244 2.71565
R740 VTAIL.n0 VTAIL.t9 2.41543
R741 VTAIL.n0 VTAIL.t15 2.41543
R742 VTAIL.n150 VTAIL.t2 2.41543
R743 VTAIL.n150 VTAIL.t4 2.41543
R744 VTAIL.n450 VTAIL.t3 2.41543
R745 VTAIL.n450 VTAIL.t1 2.41543
R746 VTAIL.n300 VTAIL.t10 2.41543
R747 VTAIL.n300 VTAIL.t8 2.41543
R748 VTAIL.n549 VTAIL.n547 2.41282
R749 VTAIL.n25 VTAIL.n23 2.41282
R750 VTAIL.n99 VTAIL.n97 2.41282
R751 VTAIL.n175 VTAIL.n173 2.41282
R752 VTAIL.n477 VTAIL.n475 2.41282
R753 VTAIL.n401 VTAIL.n399 2.41282
R754 VTAIL.n327 VTAIL.n325 2.41282
R755 VTAIL.n251 VTAIL.n249 2.41282
R756 VTAIL.n567 VTAIL.n565 1.93989
R757 VTAIL.n580 VTAIL.n579 1.93989
R758 VTAIL.n43 VTAIL.n41 1.93989
R759 VTAIL.n56 VTAIL.n55 1.93989
R760 VTAIL.n117 VTAIL.n115 1.93989
R761 VTAIL.n130 VTAIL.n129 1.93989
R762 VTAIL.n193 VTAIL.n191 1.93989
R763 VTAIL.n206 VTAIL.n205 1.93989
R764 VTAIL.n506 VTAIL.n505 1.93989
R765 VTAIL.n494 VTAIL.n493 1.93989
R766 VTAIL.n430 VTAIL.n429 1.93989
R767 VTAIL.n418 VTAIL.n417 1.93989
R768 VTAIL.n356 VTAIL.n355 1.93989
R769 VTAIL.n344 VTAIL.n343 1.93989
R770 VTAIL.n280 VTAIL.n279 1.93989
R771 VTAIL.n268 VTAIL.n267 1.93989
R772 VTAIL.n566 VTAIL.n540 1.16414
R773 VTAIL.n576 VTAIL.n536 1.16414
R774 VTAIL.n42 VTAIL.n16 1.16414
R775 VTAIL.n52 VTAIL.n12 1.16414
R776 VTAIL.n116 VTAIL.n90 1.16414
R777 VTAIL.n126 VTAIL.n86 1.16414
R778 VTAIL.n192 VTAIL.n166 1.16414
R779 VTAIL.n202 VTAIL.n162 1.16414
R780 VTAIL.n502 VTAIL.n462 1.16414
R781 VTAIL.n497 VTAIL.n467 1.16414
R782 VTAIL.n426 VTAIL.n386 1.16414
R783 VTAIL.n421 VTAIL.n391 1.16414
R784 VTAIL.n352 VTAIL.n312 1.16414
R785 VTAIL.n347 VTAIL.n317 1.16414
R786 VTAIL.n276 VTAIL.n236 1.16414
R787 VTAIL.n271 VTAIL.n241 1.16414
R788 VTAIL.n301 VTAIL.n299 0.672914
R789 VTAIL.n375 VTAIL.n301 0.672914
R790 VTAIL.n451 VTAIL.n449 0.672914
R791 VTAIL.n525 VTAIL.n451 0.672914
R792 VTAIL.n225 VTAIL.n151 0.672914
R793 VTAIL.n151 VTAIL.n149 0.672914
R794 VTAIL.n75 VTAIL.n1 0.672914
R795 VTAIL VTAIL.n599 0.614724
R796 VTAIL.n449 VTAIL.n375 0.470328
R797 VTAIL.n149 VTAIL.n75 0.470328
R798 VTAIL.n572 VTAIL.n571 0.388379
R799 VTAIL.n575 VTAIL.n538 0.388379
R800 VTAIL.n48 VTAIL.n47 0.388379
R801 VTAIL.n51 VTAIL.n14 0.388379
R802 VTAIL.n122 VTAIL.n121 0.388379
R803 VTAIL.n125 VTAIL.n88 0.388379
R804 VTAIL.n198 VTAIL.n197 0.388379
R805 VTAIL.n201 VTAIL.n164 0.388379
R806 VTAIL.n501 VTAIL.n464 0.388379
R807 VTAIL.n498 VTAIL.n466 0.388379
R808 VTAIL.n425 VTAIL.n388 0.388379
R809 VTAIL.n422 VTAIL.n390 0.388379
R810 VTAIL.n351 VTAIL.n314 0.388379
R811 VTAIL.n348 VTAIL.n316 0.388379
R812 VTAIL.n275 VTAIL.n238 0.388379
R813 VTAIL.n272 VTAIL.n240 0.388379
R814 VTAIL.n555 VTAIL.n547 0.155672
R815 VTAIL.n556 VTAIL.n555 0.155672
R816 VTAIL.n556 VTAIL.n543 0.155672
R817 VTAIL.n563 VTAIL.n543 0.155672
R818 VTAIL.n564 VTAIL.n563 0.155672
R819 VTAIL.n564 VTAIL.n539 0.155672
R820 VTAIL.n573 VTAIL.n539 0.155672
R821 VTAIL.n574 VTAIL.n573 0.155672
R822 VTAIL.n574 VTAIL.n535 0.155672
R823 VTAIL.n581 VTAIL.n535 0.155672
R824 VTAIL.n582 VTAIL.n581 0.155672
R825 VTAIL.n582 VTAIL.n531 0.155672
R826 VTAIL.n589 VTAIL.n531 0.155672
R827 VTAIL.n590 VTAIL.n589 0.155672
R828 VTAIL.n590 VTAIL.n527 0.155672
R829 VTAIL.n597 VTAIL.n527 0.155672
R830 VTAIL.n31 VTAIL.n23 0.155672
R831 VTAIL.n32 VTAIL.n31 0.155672
R832 VTAIL.n32 VTAIL.n19 0.155672
R833 VTAIL.n39 VTAIL.n19 0.155672
R834 VTAIL.n40 VTAIL.n39 0.155672
R835 VTAIL.n40 VTAIL.n15 0.155672
R836 VTAIL.n49 VTAIL.n15 0.155672
R837 VTAIL.n50 VTAIL.n49 0.155672
R838 VTAIL.n50 VTAIL.n11 0.155672
R839 VTAIL.n57 VTAIL.n11 0.155672
R840 VTAIL.n58 VTAIL.n57 0.155672
R841 VTAIL.n58 VTAIL.n7 0.155672
R842 VTAIL.n65 VTAIL.n7 0.155672
R843 VTAIL.n66 VTAIL.n65 0.155672
R844 VTAIL.n66 VTAIL.n3 0.155672
R845 VTAIL.n73 VTAIL.n3 0.155672
R846 VTAIL.n105 VTAIL.n97 0.155672
R847 VTAIL.n106 VTAIL.n105 0.155672
R848 VTAIL.n106 VTAIL.n93 0.155672
R849 VTAIL.n113 VTAIL.n93 0.155672
R850 VTAIL.n114 VTAIL.n113 0.155672
R851 VTAIL.n114 VTAIL.n89 0.155672
R852 VTAIL.n123 VTAIL.n89 0.155672
R853 VTAIL.n124 VTAIL.n123 0.155672
R854 VTAIL.n124 VTAIL.n85 0.155672
R855 VTAIL.n131 VTAIL.n85 0.155672
R856 VTAIL.n132 VTAIL.n131 0.155672
R857 VTAIL.n132 VTAIL.n81 0.155672
R858 VTAIL.n139 VTAIL.n81 0.155672
R859 VTAIL.n140 VTAIL.n139 0.155672
R860 VTAIL.n140 VTAIL.n77 0.155672
R861 VTAIL.n147 VTAIL.n77 0.155672
R862 VTAIL.n181 VTAIL.n173 0.155672
R863 VTAIL.n182 VTAIL.n181 0.155672
R864 VTAIL.n182 VTAIL.n169 0.155672
R865 VTAIL.n189 VTAIL.n169 0.155672
R866 VTAIL.n190 VTAIL.n189 0.155672
R867 VTAIL.n190 VTAIL.n165 0.155672
R868 VTAIL.n199 VTAIL.n165 0.155672
R869 VTAIL.n200 VTAIL.n199 0.155672
R870 VTAIL.n200 VTAIL.n161 0.155672
R871 VTAIL.n207 VTAIL.n161 0.155672
R872 VTAIL.n208 VTAIL.n207 0.155672
R873 VTAIL.n208 VTAIL.n157 0.155672
R874 VTAIL.n215 VTAIL.n157 0.155672
R875 VTAIL.n216 VTAIL.n215 0.155672
R876 VTAIL.n216 VTAIL.n153 0.155672
R877 VTAIL.n223 VTAIL.n153 0.155672
R878 VTAIL.n523 VTAIL.n453 0.155672
R879 VTAIL.n516 VTAIL.n453 0.155672
R880 VTAIL.n516 VTAIL.n515 0.155672
R881 VTAIL.n515 VTAIL.n457 0.155672
R882 VTAIL.n508 VTAIL.n457 0.155672
R883 VTAIL.n508 VTAIL.n507 0.155672
R884 VTAIL.n507 VTAIL.n461 0.155672
R885 VTAIL.n500 VTAIL.n461 0.155672
R886 VTAIL.n500 VTAIL.n499 0.155672
R887 VTAIL.n499 VTAIL.n465 0.155672
R888 VTAIL.n492 VTAIL.n465 0.155672
R889 VTAIL.n492 VTAIL.n491 0.155672
R890 VTAIL.n491 VTAIL.n471 0.155672
R891 VTAIL.n484 VTAIL.n471 0.155672
R892 VTAIL.n484 VTAIL.n483 0.155672
R893 VTAIL.n483 VTAIL.n475 0.155672
R894 VTAIL.n447 VTAIL.n377 0.155672
R895 VTAIL.n440 VTAIL.n377 0.155672
R896 VTAIL.n440 VTAIL.n439 0.155672
R897 VTAIL.n439 VTAIL.n381 0.155672
R898 VTAIL.n432 VTAIL.n381 0.155672
R899 VTAIL.n432 VTAIL.n431 0.155672
R900 VTAIL.n431 VTAIL.n385 0.155672
R901 VTAIL.n424 VTAIL.n385 0.155672
R902 VTAIL.n424 VTAIL.n423 0.155672
R903 VTAIL.n423 VTAIL.n389 0.155672
R904 VTAIL.n416 VTAIL.n389 0.155672
R905 VTAIL.n416 VTAIL.n415 0.155672
R906 VTAIL.n415 VTAIL.n395 0.155672
R907 VTAIL.n408 VTAIL.n395 0.155672
R908 VTAIL.n408 VTAIL.n407 0.155672
R909 VTAIL.n407 VTAIL.n399 0.155672
R910 VTAIL.n373 VTAIL.n303 0.155672
R911 VTAIL.n366 VTAIL.n303 0.155672
R912 VTAIL.n366 VTAIL.n365 0.155672
R913 VTAIL.n365 VTAIL.n307 0.155672
R914 VTAIL.n358 VTAIL.n307 0.155672
R915 VTAIL.n358 VTAIL.n357 0.155672
R916 VTAIL.n357 VTAIL.n311 0.155672
R917 VTAIL.n350 VTAIL.n311 0.155672
R918 VTAIL.n350 VTAIL.n349 0.155672
R919 VTAIL.n349 VTAIL.n315 0.155672
R920 VTAIL.n342 VTAIL.n315 0.155672
R921 VTAIL.n342 VTAIL.n341 0.155672
R922 VTAIL.n341 VTAIL.n321 0.155672
R923 VTAIL.n334 VTAIL.n321 0.155672
R924 VTAIL.n334 VTAIL.n333 0.155672
R925 VTAIL.n333 VTAIL.n325 0.155672
R926 VTAIL.n297 VTAIL.n227 0.155672
R927 VTAIL.n290 VTAIL.n227 0.155672
R928 VTAIL.n290 VTAIL.n289 0.155672
R929 VTAIL.n289 VTAIL.n231 0.155672
R930 VTAIL.n282 VTAIL.n231 0.155672
R931 VTAIL.n282 VTAIL.n281 0.155672
R932 VTAIL.n281 VTAIL.n235 0.155672
R933 VTAIL.n274 VTAIL.n235 0.155672
R934 VTAIL.n274 VTAIL.n273 0.155672
R935 VTAIL.n273 VTAIL.n239 0.155672
R936 VTAIL.n266 VTAIL.n239 0.155672
R937 VTAIL.n266 VTAIL.n265 0.155672
R938 VTAIL.n265 VTAIL.n245 0.155672
R939 VTAIL.n258 VTAIL.n245 0.155672
R940 VTAIL.n258 VTAIL.n257 0.155672
R941 VTAIL.n257 VTAIL.n249 0.155672
R942 VTAIL VTAIL.n1 0.0586897
R943 VDD2.n2 VDD2.n1 70.6222
R944 VDD2.n2 VDD2.n0 70.6222
R945 VDD2 VDD2.n5 70.6193
R946 VDD2.n4 VDD2.n3 70.3415
R947 VDD2.n4 VDD2.n2 38.3446
R948 VDD2.n5 VDD2.t0 2.41543
R949 VDD2.n5 VDD2.t2 2.41543
R950 VDD2.n3 VDD2.t3 2.41543
R951 VDD2.n3 VDD2.t1 2.41543
R952 VDD2.n1 VDD2.t6 2.41543
R953 VDD2.n1 VDD2.t7 2.41543
R954 VDD2.n0 VDD2.t4 2.41543
R955 VDD2.n0 VDD2.t5 2.41543
R956 VDD2 VDD2.n4 0.394897
R957 B.n117 B.t9 928.605
R958 B.n111 B.t0 928.605
R959 B.n43 B.t3 928.605
R960 B.n36 B.t6 928.605
R961 B.n330 B.n87 585
R962 B.n329 B.n328 585
R963 B.n327 B.n88 585
R964 B.n326 B.n325 585
R965 B.n324 B.n89 585
R966 B.n323 B.n322 585
R967 B.n321 B.n90 585
R968 B.n320 B.n319 585
R969 B.n318 B.n91 585
R970 B.n317 B.n316 585
R971 B.n315 B.n92 585
R972 B.n314 B.n313 585
R973 B.n312 B.n93 585
R974 B.n311 B.n310 585
R975 B.n309 B.n94 585
R976 B.n308 B.n307 585
R977 B.n306 B.n95 585
R978 B.n305 B.n304 585
R979 B.n303 B.n96 585
R980 B.n302 B.n301 585
R981 B.n300 B.n97 585
R982 B.n299 B.n298 585
R983 B.n297 B.n98 585
R984 B.n296 B.n295 585
R985 B.n294 B.n99 585
R986 B.n293 B.n292 585
R987 B.n291 B.n100 585
R988 B.n290 B.n289 585
R989 B.n288 B.n101 585
R990 B.n287 B.n286 585
R991 B.n285 B.n102 585
R992 B.n284 B.n283 585
R993 B.n282 B.n103 585
R994 B.n281 B.n280 585
R995 B.n279 B.n104 585
R996 B.n278 B.n277 585
R997 B.n276 B.n105 585
R998 B.n275 B.n274 585
R999 B.n273 B.n106 585
R1000 B.n272 B.n271 585
R1001 B.n270 B.n107 585
R1002 B.n269 B.n268 585
R1003 B.n267 B.n108 585
R1004 B.n266 B.n265 585
R1005 B.n264 B.n109 585
R1006 B.n263 B.n262 585
R1007 B.n260 B.n110 585
R1008 B.n259 B.n258 585
R1009 B.n257 B.n113 585
R1010 B.n256 B.n255 585
R1011 B.n254 B.n114 585
R1012 B.n253 B.n252 585
R1013 B.n251 B.n115 585
R1014 B.n250 B.n249 585
R1015 B.n248 B.n116 585
R1016 B.n246 B.n245 585
R1017 B.n244 B.n119 585
R1018 B.n243 B.n242 585
R1019 B.n241 B.n120 585
R1020 B.n240 B.n239 585
R1021 B.n238 B.n121 585
R1022 B.n237 B.n236 585
R1023 B.n235 B.n122 585
R1024 B.n234 B.n233 585
R1025 B.n232 B.n123 585
R1026 B.n231 B.n230 585
R1027 B.n229 B.n124 585
R1028 B.n228 B.n227 585
R1029 B.n226 B.n125 585
R1030 B.n225 B.n224 585
R1031 B.n223 B.n126 585
R1032 B.n222 B.n221 585
R1033 B.n220 B.n127 585
R1034 B.n219 B.n218 585
R1035 B.n217 B.n128 585
R1036 B.n216 B.n215 585
R1037 B.n214 B.n129 585
R1038 B.n213 B.n212 585
R1039 B.n211 B.n130 585
R1040 B.n210 B.n209 585
R1041 B.n208 B.n131 585
R1042 B.n207 B.n206 585
R1043 B.n205 B.n132 585
R1044 B.n204 B.n203 585
R1045 B.n202 B.n133 585
R1046 B.n201 B.n200 585
R1047 B.n199 B.n134 585
R1048 B.n198 B.n197 585
R1049 B.n196 B.n135 585
R1050 B.n195 B.n194 585
R1051 B.n193 B.n136 585
R1052 B.n192 B.n191 585
R1053 B.n190 B.n137 585
R1054 B.n189 B.n188 585
R1055 B.n187 B.n138 585
R1056 B.n186 B.n185 585
R1057 B.n184 B.n139 585
R1058 B.n183 B.n182 585
R1059 B.n181 B.n140 585
R1060 B.n180 B.n179 585
R1061 B.n178 B.n141 585
R1062 B.n332 B.n331 585
R1063 B.n333 B.n86 585
R1064 B.n335 B.n334 585
R1065 B.n336 B.n85 585
R1066 B.n338 B.n337 585
R1067 B.n339 B.n84 585
R1068 B.n341 B.n340 585
R1069 B.n342 B.n83 585
R1070 B.n344 B.n343 585
R1071 B.n345 B.n82 585
R1072 B.n347 B.n346 585
R1073 B.n348 B.n81 585
R1074 B.n350 B.n349 585
R1075 B.n351 B.n80 585
R1076 B.n353 B.n352 585
R1077 B.n354 B.n79 585
R1078 B.n356 B.n355 585
R1079 B.n357 B.n78 585
R1080 B.n359 B.n358 585
R1081 B.n360 B.n77 585
R1082 B.n362 B.n361 585
R1083 B.n363 B.n76 585
R1084 B.n365 B.n364 585
R1085 B.n366 B.n75 585
R1086 B.n368 B.n367 585
R1087 B.n369 B.n74 585
R1088 B.n371 B.n370 585
R1089 B.n372 B.n73 585
R1090 B.n374 B.n373 585
R1091 B.n375 B.n72 585
R1092 B.n377 B.n376 585
R1093 B.n378 B.n71 585
R1094 B.n380 B.n379 585
R1095 B.n381 B.n70 585
R1096 B.n383 B.n382 585
R1097 B.n384 B.n69 585
R1098 B.n386 B.n385 585
R1099 B.n387 B.n68 585
R1100 B.n389 B.n388 585
R1101 B.n390 B.n67 585
R1102 B.n543 B.n542 585
R1103 B.n541 B.n12 585
R1104 B.n540 B.n539 585
R1105 B.n538 B.n13 585
R1106 B.n537 B.n536 585
R1107 B.n535 B.n14 585
R1108 B.n534 B.n533 585
R1109 B.n532 B.n15 585
R1110 B.n531 B.n530 585
R1111 B.n529 B.n16 585
R1112 B.n528 B.n527 585
R1113 B.n526 B.n17 585
R1114 B.n525 B.n524 585
R1115 B.n523 B.n18 585
R1116 B.n522 B.n521 585
R1117 B.n520 B.n19 585
R1118 B.n519 B.n518 585
R1119 B.n517 B.n20 585
R1120 B.n516 B.n515 585
R1121 B.n514 B.n21 585
R1122 B.n513 B.n512 585
R1123 B.n511 B.n22 585
R1124 B.n510 B.n509 585
R1125 B.n508 B.n23 585
R1126 B.n507 B.n506 585
R1127 B.n505 B.n24 585
R1128 B.n504 B.n503 585
R1129 B.n502 B.n25 585
R1130 B.n501 B.n500 585
R1131 B.n499 B.n26 585
R1132 B.n498 B.n497 585
R1133 B.n496 B.n27 585
R1134 B.n495 B.n494 585
R1135 B.n493 B.n28 585
R1136 B.n492 B.n491 585
R1137 B.n490 B.n29 585
R1138 B.n489 B.n488 585
R1139 B.n487 B.n30 585
R1140 B.n486 B.n485 585
R1141 B.n484 B.n31 585
R1142 B.n483 B.n482 585
R1143 B.n481 B.n32 585
R1144 B.n480 B.n479 585
R1145 B.n478 B.n33 585
R1146 B.n477 B.n476 585
R1147 B.n475 B.n34 585
R1148 B.n474 B.n473 585
R1149 B.n472 B.n35 585
R1150 B.n471 B.n470 585
R1151 B.n469 B.n39 585
R1152 B.n468 B.n467 585
R1153 B.n466 B.n40 585
R1154 B.n465 B.n464 585
R1155 B.n463 B.n41 585
R1156 B.n462 B.n461 585
R1157 B.n459 B.n42 585
R1158 B.n458 B.n457 585
R1159 B.n456 B.n45 585
R1160 B.n455 B.n454 585
R1161 B.n453 B.n46 585
R1162 B.n452 B.n451 585
R1163 B.n450 B.n47 585
R1164 B.n449 B.n448 585
R1165 B.n447 B.n48 585
R1166 B.n446 B.n445 585
R1167 B.n444 B.n49 585
R1168 B.n443 B.n442 585
R1169 B.n441 B.n50 585
R1170 B.n440 B.n439 585
R1171 B.n438 B.n51 585
R1172 B.n437 B.n436 585
R1173 B.n435 B.n52 585
R1174 B.n434 B.n433 585
R1175 B.n432 B.n53 585
R1176 B.n431 B.n430 585
R1177 B.n429 B.n54 585
R1178 B.n428 B.n427 585
R1179 B.n426 B.n55 585
R1180 B.n425 B.n424 585
R1181 B.n423 B.n56 585
R1182 B.n422 B.n421 585
R1183 B.n420 B.n57 585
R1184 B.n419 B.n418 585
R1185 B.n417 B.n58 585
R1186 B.n416 B.n415 585
R1187 B.n414 B.n59 585
R1188 B.n413 B.n412 585
R1189 B.n411 B.n60 585
R1190 B.n410 B.n409 585
R1191 B.n408 B.n61 585
R1192 B.n407 B.n406 585
R1193 B.n405 B.n62 585
R1194 B.n404 B.n403 585
R1195 B.n402 B.n63 585
R1196 B.n401 B.n400 585
R1197 B.n399 B.n64 585
R1198 B.n398 B.n397 585
R1199 B.n396 B.n65 585
R1200 B.n395 B.n394 585
R1201 B.n393 B.n66 585
R1202 B.n392 B.n391 585
R1203 B.n544 B.n11 585
R1204 B.n546 B.n545 585
R1205 B.n547 B.n10 585
R1206 B.n549 B.n548 585
R1207 B.n550 B.n9 585
R1208 B.n552 B.n551 585
R1209 B.n553 B.n8 585
R1210 B.n555 B.n554 585
R1211 B.n556 B.n7 585
R1212 B.n558 B.n557 585
R1213 B.n559 B.n6 585
R1214 B.n561 B.n560 585
R1215 B.n562 B.n5 585
R1216 B.n564 B.n563 585
R1217 B.n565 B.n4 585
R1218 B.n567 B.n566 585
R1219 B.n568 B.n3 585
R1220 B.n570 B.n569 585
R1221 B.n571 B.n0 585
R1222 B.n2 B.n1 585
R1223 B.n151 B.n150 585
R1224 B.n153 B.n152 585
R1225 B.n154 B.n149 585
R1226 B.n156 B.n155 585
R1227 B.n157 B.n148 585
R1228 B.n159 B.n158 585
R1229 B.n160 B.n147 585
R1230 B.n162 B.n161 585
R1231 B.n163 B.n146 585
R1232 B.n165 B.n164 585
R1233 B.n166 B.n145 585
R1234 B.n168 B.n167 585
R1235 B.n169 B.n144 585
R1236 B.n171 B.n170 585
R1237 B.n172 B.n143 585
R1238 B.n174 B.n173 585
R1239 B.n175 B.n142 585
R1240 B.n177 B.n176 585
R1241 B.n178 B.n177 545.355
R1242 B.n331 B.n330 545.355
R1243 B.n391 B.n390 545.355
R1244 B.n542 B.n11 545.355
R1245 B.n111 B.t1 417.091
R1246 B.n43 B.t5 417.091
R1247 B.n117 B.t10 417.091
R1248 B.n36 B.t8 417.091
R1249 B.n112 B.t2 401.964
R1250 B.n44 B.t4 401.964
R1251 B.n118 B.t11 401.964
R1252 B.n37 B.t7 401.964
R1253 B.n573 B.n572 256.663
R1254 B.n572 B.n571 235.042
R1255 B.n572 B.n2 235.042
R1256 B.n179 B.n178 163.367
R1257 B.n179 B.n140 163.367
R1258 B.n183 B.n140 163.367
R1259 B.n184 B.n183 163.367
R1260 B.n185 B.n184 163.367
R1261 B.n185 B.n138 163.367
R1262 B.n189 B.n138 163.367
R1263 B.n190 B.n189 163.367
R1264 B.n191 B.n190 163.367
R1265 B.n191 B.n136 163.367
R1266 B.n195 B.n136 163.367
R1267 B.n196 B.n195 163.367
R1268 B.n197 B.n196 163.367
R1269 B.n197 B.n134 163.367
R1270 B.n201 B.n134 163.367
R1271 B.n202 B.n201 163.367
R1272 B.n203 B.n202 163.367
R1273 B.n203 B.n132 163.367
R1274 B.n207 B.n132 163.367
R1275 B.n208 B.n207 163.367
R1276 B.n209 B.n208 163.367
R1277 B.n209 B.n130 163.367
R1278 B.n213 B.n130 163.367
R1279 B.n214 B.n213 163.367
R1280 B.n215 B.n214 163.367
R1281 B.n215 B.n128 163.367
R1282 B.n219 B.n128 163.367
R1283 B.n220 B.n219 163.367
R1284 B.n221 B.n220 163.367
R1285 B.n221 B.n126 163.367
R1286 B.n225 B.n126 163.367
R1287 B.n226 B.n225 163.367
R1288 B.n227 B.n226 163.367
R1289 B.n227 B.n124 163.367
R1290 B.n231 B.n124 163.367
R1291 B.n232 B.n231 163.367
R1292 B.n233 B.n232 163.367
R1293 B.n233 B.n122 163.367
R1294 B.n237 B.n122 163.367
R1295 B.n238 B.n237 163.367
R1296 B.n239 B.n238 163.367
R1297 B.n239 B.n120 163.367
R1298 B.n243 B.n120 163.367
R1299 B.n244 B.n243 163.367
R1300 B.n245 B.n244 163.367
R1301 B.n245 B.n116 163.367
R1302 B.n250 B.n116 163.367
R1303 B.n251 B.n250 163.367
R1304 B.n252 B.n251 163.367
R1305 B.n252 B.n114 163.367
R1306 B.n256 B.n114 163.367
R1307 B.n257 B.n256 163.367
R1308 B.n258 B.n257 163.367
R1309 B.n258 B.n110 163.367
R1310 B.n263 B.n110 163.367
R1311 B.n264 B.n263 163.367
R1312 B.n265 B.n264 163.367
R1313 B.n265 B.n108 163.367
R1314 B.n269 B.n108 163.367
R1315 B.n270 B.n269 163.367
R1316 B.n271 B.n270 163.367
R1317 B.n271 B.n106 163.367
R1318 B.n275 B.n106 163.367
R1319 B.n276 B.n275 163.367
R1320 B.n277 B.n276 163.367
R1321 B.n277 B.n104 163.367
R1322 B.n281 B.n104 163.367
R1323 B.n282 B.n281 163.367
R1324 B.n283 B.n282 163.367
R1325 B.n283 B.n102 163.367
R1326 B.n287 B.n102 163.367
R1327 B.n288 B.n287 163.367
R1328 B.n289 B.n288 163.367
R1329 B.n289 B.n100 163.367
R1330 B.n293 B.n100 163.367
R1331 B.n294 B.n293 163.367
R1332 B.n295 B.n294 163.367
R1333 B.n295 B.n98 163.367
R1334 B.n299 B.n98 163.367
R1335 B.n300 B.n299 163.367
R1336 B.n301 B.n300 163.367
R1337 B.n301 B.n96 163.367
R1338 B.n305 B.n96 163.367
R1339 B.n306 B.n305 163.367
R1340 B.n307 B.n306 163.367
R1341 B.n307 B.n94 163.367
R1342 B.n311 B.n94 163.367
R1343 B.n312 B.n311 163.367
R1344 B.n313 B.n312 163.367
R1345 B.n313 B.n92 163.367
R1346 B.n317 B.n92 163.367
R1347 B.n318 B.n317 163.367
R1348 B.n319 B.n318 163.367
R1349 B.n319 B.n90 163.367
R1350 B.n323 B.n90 163.367
R1351 B.n324 B.n323 163.367
R1352 B.n325 B.n324 163.367
R1353 B.n325 B.n88 163.367
R1354 B.n329 B.n88 163.367
R1355 B.n330 B.n329 163.367
R1356 B.n390 B.n389 163.367
R1357 B.n389 B.n68 163.367
R1358 B.n385 B.n68 163.367
R1359 B.n385 B.n384 163.367
R1360 B.n384 B.n383 163.367
R1361 B.n383 B.n70 163.367
R1362 B.n379 B.n70 163.367
R1363 B.n379 B.n378 163.367
R1364 B.n378 B.n377 163.367
R1365 B.n377 B.n72 163.367
R1366 B.n373 B.n72 163.367
R1367 B.n373 B.n372 163.367
R1368 B.n372 B.n371 163.367
R1369 B.n371 B.n74 163.367
R1370 B.n367 B.n74 163.367
R1371 B.n367 B.n366 163.367
R1372 B.n366 B.n365 163.367
R1373 B.n365 B.n76 163.367
R1374 B.n361 B.n76 163.367
R1375 B.n361 B.n360 163.367
R1376 B.n360 B.n359 163.367
R1377 B.n359 B.n78 163.367
R1378 B.n355 B.n78 163.367
R1379 B.n355 B.n354 163.367
R1380 B.n354 B.n353 163.367
R1381 B.n353 B.n80 163.367
R1382 B.n349 B.n80 163.367
R1383 B.n349 B.n348 163.367
R1384 B.n348 B.n347 163.367
R1385 B.n347 B.n82 163.367
R1386 B.n343 B.n82 163.367
R1387 B.n343 B.n342 163.367
R1388 B.n342 B.n341 163.367
R1389 B.n341 B.n84 163.367
R1390 B.n337 B.n84 163.367
R1391 B.n337 B.n336 163.367
R1392 B.n336 B.n335 163.367
R1393 B.n335 B.n86 163.367
R1394 B.n331 B.n86 163.367
R1395 B.n542 B.n541 163.367
R1396 B.n541 B.n540 163.367
R1397 B.n540 B.n13 163.367
R1398 B.n536 B.n13 163.367
R1399 B.n536 B.n535 163.367
R1400 B.n535 B.n534 163.367
R1401 B.n534 B.n15 163.367
R1402 B.n530 B.n15 163.367
R1403 B.n530 B.n529 163.367
R1404 B.n529 B.n528 163.367
R1405 B.n528 B.n17 163.367
R1406 B.n524 B.n17 163.367
R1407 B.n524 B.n523 163.367
R1408 B.n523 B.n522 163.367
R1409 B.n522 B.n19 163.367
R1410 B.n518 B.n19 163.367
R1411 B.n518 B.n517 163.367
R1412 B.n517 B.n516 163.367
R1413 B.n516 B.n21 163.367
R1414 B.n512 B.n21 163.367
R1415 B.n512 B.n511 163.367
R1416 B.n511 B.n510 163.367
R1417 B.n510 B.n23 163.367
R1418 B.n506 B.n23 163.367
R1419 B.n506 B.n505 163.367
R1420 B.n505 B.n504 163.367
R1421 B.n504 B.n25 163.367
R1422 B.n500 B.n25 163.367
R1423 B.n500 B.n499 163.367
R1424 B.n499 B.n498 163.367
R1425 B.n498 B.n27 163.367
R1426 B.n494 B.n27 163.367
R1427 B.n494 B.n493 163.367
R1428 B.n493 B.n492 163.367
R1429 B.n492 B.n29 163.367
R1430 B.n488 B.n29 163.367
R1431 B.n488 B.n487 163.367
R1432 B.n487 B.n486 163.367
R1433 B.n486 B.n31 163.367
R1434 B.n482 B.n31 163.367
R1435 B.n482 B.n481 163.367
R1436 B.n481 B.n480 163.367
R1437 B.n480 B.n33 163.367
R1438 B.n476 B.n33 163.367
R1439 B.n476 B.n475 163.367
R1440 B.n475 B.n474 163.367
R1441 B.n474 B.n35 163.367
R1442 B.n470 B.n35 163.367
R1443 B.n470 B.n469 163.367
R1444 B.n469 B.n468 163.367
R1445 B.n468 B.n40 163.367
R1446 B.n464 B.n40 163.367
R1447 B.n464 B.n463 163.367
R1448 B.n463 B.n462 163.367
R1449 B.n462 B.n42 163.367
R1450 B.n457 B.n42 163.367
R1451 B.n457 B.n456 163.367
R1452 B.n456 B.n455 163.367
R1453 B.n455 B.n46 163.367
R1454 B.n451 B.n46 163.367
R1455 B.n451 B.n450 163.367
R1456 B.n450 B.n449 163.367
R1457 B.n449 B.n48 163.367
R1458 B.n445 B.n48 163.367
R1459 B.n445 B.n444 163.367
R1460 B.n444 B.n443 163.367
R1461 B.n443 B.n50 163.367
R1462 B.n439 B.n50 163.367
R1463 B.n439 B.n438 163.367
R1464 B.n438 B.n437 163.367
R1465 B.n437 B.n52 163.367
R1466 B.n433 B.n52 163.367
R1467 B.n433 B.n432 163.367
R1468 B.n432 B.n431 163.367
R1469 B.n431 B.n54 163.367
R1470 B.n427 B.n54 163.367
R1471 B.n427 B.n426 163.367
R1472 B.n426 B.n425 163.367
R1473 B.n425 B.n56 163.367
R1474 B.n421 B.n56 163.367
R1475 B.n421 B.n420 163.367
R1476 B.n420 B.n419 163.367
R1477 B.n419 B.n58 163.367
R1478 B.n415 B.n58 163.367
R1479 B.n415 B.n414 163.367
R1480 B.n414 B.n413 163.367
R1481 B.n413 B.n60 163.367
R1482 B.n409 B.n60 163.367
R1483 B.n409 B.n408 163.367
R1484 B.n408 B.n407 163.367
R1485 B.n407 B.n62 163.367
R1486 B.n403 B.n62 163.367
R1487 B.n403 B.n402 163.367
R1488 B.n402 B.n401 163.367
R1489 B.n401 B.n64 163.367
R1490 B.n397 B.n64 163.367
R1491 B.n397 B.n396 163.367
R1492 B.n396 B.n395 163.367
R1493 B.n395 B.n66 163.367
R1494 B.n391 B.n66 163.367
R1495 B.n546 B.n11 163.367
R1496 B.n547 B.n546 163.367
R1497 B.n548 B.n547 163.367
R1498 B.n548 B.n9 163.367
R1499 B.n552 B.n9 163.367
R1500 B.n553 B.n552 163.367
R1501 B.n554 B.n553 163.367
R1502 B.n554 B.n7 163.367
R1503 B.n558 B.n7 163.367
R1504 B.n559 B.n558 163.367
R1505 B.n560 B.n559 163.367
R1506 B.n560 B.n5 163.367
R1507 B.n564 B.n5 163.367
R1508 B.n565 B.n564 163.367
R1509 B.n566 B.n565 163.367
R1510 B.n566 B.n3 163.367
R1511 B.n570 B.n3 163.367
R1512 B.n571 B.n570 163.367
R1513 B.n150 B.n2 163.367
R1514 B.n153 B.n150 163.367
R1515 B.n154 B.n153 163.367
R1516 B.n155 B.n154 163.367
R1517 B.n155 B.n148 163.367
R1518 B.n159 B.n148 163.367
R1519 B.n160 B.n159 163.367
R1520 B.n161 B.n160 163.367
R1521 B.n161 B.n146 163.367
R1522 B.n165 B.n146 163.367
R1523 B.n166 B.n165 163.367
R1524 B.n167 B.n166 163.367
R1525 B.n167 B.n144 163.367
R1526 B.n171 B.n144 163.367
R1527 B.n172 B.n171 163.367
R1528 B.n173 B.n172 163.367
R1529 B.n173 B.n142 163.367
R1530 B.n177 B.n142 163.367
R1531 B.n247 B.n118 59.5399
R1532 B.n261 B.n112 59.5399
R1533 B.n460 B.n44 59.5399
R1534 B.n38 B.n37 59.5399
R1535 B.n544 B.n543 35.4346
R1536 B.n392 B.n67 35.4346
R1537 B.n176 B.n141 35.4346
R1538 B.n332 B.n87 35.4346
R1539 B B.n573 18.0485
R1540 B.n118 B.n117 15.1278
R1541 B.n112 B.n111 15.1278
R1542 B.n44 B.n43 15.1278
R1543 B.n37 B.n36 15.1278
R1544 B.n545 B.n544 10.6151
R1545 B.n545 B.n10 10.6151
R1546 B.n549 B.n10 10.6151
R1547 B.n550 B.n549 10.6151
R1548 B.n551 B.n550 10.6151
R1549 B.n551 B.n8 10.6151
R1550 B.n555 B.n8 10.6151
R1551 B.n556 B.n555 10.6151
R1552 B.n557 B.n556 10.6151
R1553 B.n557 B.n6 10.6151
R1554 B.n561 B.n6 10.6151
R1555 B.n562 B.n561 10.6151
R1556 B.n563 B.n562 10.6151
R1557 B.n563 B.n4 10.6151
R1558 B.n567 B.n4 10.6151
R1559 B.n568 B.n567 10.6151
R1560 B.n569 B.n568 10.6151
R1561 B.n569 B.n0 10.6151
R1562 B.n543 B.n12 10.6151
R1563 B.n539 B.n12 10.6151
R1564 B.n539 B.n538 10.6151
R1565 B.n538 B.n537 10.6151
R1566 B.n537 B.n14 10.6151
R1567 B.n533 B.n14 10.6151
R1568 B.n533 B.n532 10.6151
R1569 B.n532 B.n531 10.6151
R1570 B.n531 B.n16 10.6151
R1571 B.n527 B.n16 10.6151
R1572 B.n527 B.n526 10.6151
R1573 B.n526 B.n525 10.6151
R1574 B.n525 B.n18 10.6151
R1575 B.n521 B.n18 10.6151
R1576 B.n521 B.n520 10.6151
R1577 B.n520 B.n519 10.6151
R1578 B.n519 B.n20 10.6151
R1579 B.n515 B.n20 10.6151
R1580 B.n515 B.n514 10.6151
R1581 B.n514 B.n513 10.6151
R1582 B.n513 B.n22 10.6151
R1583 B.n509 B.n22 10.6151
R1584 B.n509 B.n508 10.6151
R1585 B.n508 B.n507 10.6151
R1586 B.n507 B.n24 10.6151
R1587 B.n503 B.n24 10.6151
R1588 B.n503 B.n502 10.6151
R1589 B.n502 B.n501 10.6151
R1590 B.n501 B.n26 10.6151
R1591 B.n497 B.n26 10.6151
R1592 B.n497 B.n496 10.6151
R1593 B.n496 B.n495 10.6151
R1594 B.n495 B.n28 10.6151
R1595 B.n491 B.n28 10.6151
R1596 B.n491 B.n490 10.6151
R1597 B.n490 B.n489 10.6151
R1598 B.n489 B.n30 10.6151
R1599 B.n485 B.n30 10.6151
R1600 B.n485 B.n484 10.6151
R1601 B.n484 B.n483 10.6151
R1602 B.n483 B.n32 10.6151
R1603 B.n479 B.n32 10.6151
R1604 B.n479 B.n478 10.6151
R1605 B.n478 B.n477 10.6151
R1606 B.n477 B.n34 10.6151
R1607 B.n473 B.n472 10.6151
R1608 B.n472 B.n471 10.6151
R1609 B.n471 B.n39 10.6151
R1610 B.n467 B.n39 10.6151
R1611 B.n467 B.n466 10.6151
R1612 B.n466 B.n465 10.6151
R1613 B.n465 B.n41 10.6151
R1614 B.n461 B.n41 10.6151
R1615 B.n459 B.n458 10.6151
R1616 B.n458 B.n45 10.6151
R1617 B.n454 B.n45 10.6151
R1618 B.n454 B.n453 10.6151
R1619 B.n453 B.n452 10.6151
R1620 B.n452 B.n47 10.6151
R1621 B.n448 B.n47 10.6151
R1622 B.n448 B.n447 10.6151
R1623 B.n447 B.n446 10.6151
R1624 B.n446 B.n49 10.6151
R1625 B.n442 B.n49 10.6151
R1626 B.n442 B.n441 10.6151
R1627 B.n441 B.n440 10.6151
R1628 B.n440 B.n51 10.6151
R1629 B.n436 B.n51 10.6151
R1630 B.n436 B.n435 10.6151
R1631 B.n435 B.n434 10.6151
R1632 B.n434 B.n53 10.6151
R1633 B.n430 B.n53 10.6151
R1634 B.n430 B.n429 10.6151
R1635 B.n429 B.n428 10.6151
R1636 B.n428 B.n55 10.6151
R1637 B.n424 B.n55 10.6151
R1638 B.n424 B.n423 10.6151
R1639 B.n423 B.n422 10.6151
R1640 B.n422 B.n57 10.6151
R1641 B.n418 B.n57 10.6151
R1642 B.n418 B.n417 10.6151
R1643 B.n417 B.n416 10.6151
R1644 B.n416 B.n59 10.6151
R1645 B.n412 B.n59 10.6151
R1646 B.n412 B.n411 10.6151
R1647 B.n411 B.n410 10.6151
R1648 B.n410 B.n61 10.6151
R1649 B.n406 B.n61 10.6151
R1650 B.n406 B.n405 10.6151
R1651 B.n405 B.n404 10.6151
R1652 B.n404 B.n63 10.6151
R1653 B.n400 B.n63 10.6151
R1654 B.n400 B.n399 10.6151
R1655 B.n399 B.n398 10.6151
R1656 B.n398 B.n65 10.6151
R1657 B.n394 B.n65 10.6151
R1658 B.n394 B.n393 10.6151
R1659 B.n393 B.n392 10.6151
R1660 B.n388 B.n67 10.6151
R1661 B.n388 B.n387 10.6151
R1662 B.n387 B.n386 10.6151
R1663 B.n386 B.n69 10.6151
R1664 B.n382 B.n69 10.6151
R1665 B.n382 B.n381 10.6151
R1666 B.n381 B.n380 10.6151
R1667 B.n380 B.n71 10.6151
R1668 B.n376 B.n71 10.6151
R1669 B.n376 B.n375 10.6151
R1670 B.n375 B.n374 10.6151
R1671 B.n374 B.n73 10.6151
R1672 B.n370 B.n73 10.6151
R1673 B.n370 B.n369 10.6151
R1674 B.n369 B.n368 10.6151
R1675 B.n368 B.n75 10.6151
R1676 B.n364 B.n75 10.6151
R1677 B.n364 B.n363 10.6151
R1678 B.n363 B.n362 10.6151
R1679 B.n362 B.n77 10.6151
R1680 B.n358 B.n77 10.6151
R1681 B.n358 B.n357 10.6151
R1682 B.n357 B.n356 10.6151
R1683 B.n356 B.n79 10.6151
R1684 B.n352 B.n79 10.6151
R1685 B.n352 B.n351 10.6151
R1686 B.n351 B.n350 10.6151
R1687 B.n350 B.n81 10.6151
R1688 B.n346 B.n81 10.6151
R1689 B.n346 B.n345 10.6151
R1690 B.n345 B.n344 10.6151
R1691 B.n344 B.n83 10.6151
R1692 B.n340 B.n83 10.6151
R1693 B.n340 B.n339 10.6151
R1694 B.n339 B.n338 10.6151
R1695 B.n338 B.n85 10.6151
R1696 B.n334 B.n85 10.6151
R1697 B.n334 B.n333 10.6151
R1698 B.n333 B.n332 10.6151
R1699 B.n151 B.n1 10.6151
R1700 B.n152 B.n151 10.6151
R1701 B.n152 B.n149 10.6151
R1702 B.n156 B.n149 10.6151
R1703 B.n157 B.n156 10.6151
R1704 B.n158 B.n157 10.6151
R1705 B.n158 B.n147 10.6151
R1706 B.n162 B.n147 10.6151
R1707 B.n163 B.n162 10.6151
R1708 B.n164 B.n163 10.6151
R1709 B.n164 B.n145 10.6151
R1710 B.n168 B.n145 10.6151
R1711 B.n169 B.n168 10.6151
R1712 B.n170 B.n169 10.6151
R1713 B.n170 B.n143 10.6151
R1714 B.n174 B.n143 10.6151
R1715 B.n175 B.n174 10.6151
R1716 B.n176 B.n175 10.6151
R1717 B.n180 B.n141 10.6151
R1718 B.n181 B.n180 10.6151
R1719 B.n182 B.n181 10.6151
R1720 B.n182 B.n139 10.6151
R1721 B.n186 B.n139 10.6151
R1722 B.n187 B.n186 10.6151
R1723 B.n188 B.n187 10.6151
R1724 B.n188 B.n137 10.6151
R1725 B.n192 B.n137 10.6151
R1726 B.n193 B.n192 10.6151
R1727 B.n194 B.n193 10.6151
R1728 B.n194 B.n135 10.6151
R1729 B.n198 B.n135 10.6151
R1730 B.n199 B.n198 10.6151
R1731 B.n200 B.n199 10.6151
R1732 B.n200 B.n133 10.6151
R1733 B.n204 B.n133 10.6151
R1734 B.n205 B.n204 10.6151
R1735 B.n206 B.n205 10.6151
R1736 B.n206 B.n131 10.6151
R1737 B.n210 B.n131 10.6151
R1738 B.n211 B.n210 10.6151
R1739 B.n212 B.n211 10.6151
R1740 B.n212 B.n129 10.6151
R1741 B.n216 B.n129 10.6151
R1742 B.n217 B.n216 10.6151
R1743 B.n218 B.n217 10.6151
R1744 B.n218 B.n127 10.6151
R1745 B.n222 B.n127 10.6151
R1746 B.n223 B.n222 10.6151
R1747 B.n224 B.n223 10.6151
R1748 B.n224 B.n125 10.6151
R1749 B.n228 B.n125 10.6151
R1750 B.n229 B.n228 10.6151
R1751 B.n230 B.n229 10.6151
R1752 B.n230 B.n123 10.6151
R1753 B.n234 B.n123 10.6151
R1754 B.n235 B.n234 10.6151
R1755 B.n236 B.n235 10.6151
R1756 B.n236 B.n121 10.6151
R1757 B.n240 B.n121 10.6151
R1758 B.n241 B.n240 10.6151
R1759 B.n242 B.n241 10.6151
R1760 B.n242 B.n119 10.6151
R1761 B.n246 B.n119 10.6151
R1762 B.n249 B.n248 10.6151
R1763 B.n249 B.n115 10.6151
R1764 B.n253 B.n115 10.6151
R1765 B.n254 B.n253 10.6151
R1766 B.n255 B.n254 10.6151
R1767 B.n255 B.n113 10.6151
R1768 B.n259 B.n113 10.6151
R1769 B.n260 B.n259 10.6151
R1770 B.n262 B.n109 10.6151
R1771 B.n266 B.n109 10.6151
R1772 B.n267 B.n266 10.6151
R1773 B.n268 B.n267 10.6151
R1774 B.n268 B.n107 10.6151
R1775 B.n272 B.n107 10.6151
R1776 B.n273 B.n272 10.6151
R1777 B.n274 B.n273 10.6151
R1778 B.n274 B.n105 10.6151
R1779 B.n278 B.n105 10.6151
R1780 B.n279 B.n278 10.6151
R1781 B.n280 B.n279 10.6151
R1782 B.n280 B.n103 10.6151
R1783 B.n284 B.n103 10.6151
R1784 B.n285 B.n284 10.6151
R1785 B.n286 B.n285 10.6151
R1786 B.n286 B.n101 10.6151
R1787 B.n290 B.n101 10.6151
R1788 B.n291 B.n290 10.6151
R1789 B.n292 B.n291 10.6151
R1790 B.n292 B.n99 10.6151
R1791 B.n296 B.n99 10.6151
R1792 B.n297 B.n296 10.6151
R1793 B.n298 B.n297 10.6151
R1794 B.n298 B.n97 10.6151
R1795 B.n302 B.n97 10.6151
R1796 B.n303 B.n302 10.6151
R1797 B.n304 B.n303 10.6151
R1798 B.n304 B.n95 10.6151
R1799 B.n308 B.n95 10.6151
R1800 B.n309 B.n308 10.6151
R1801 B.n310 B.n309 10.6151
R1802 B.n310 B.n93 10.6151
R1803 B.n314 B.n93 10.6151
R1804 B.n315 B.n314 10.6151
R1805 B.n316 B.n315 10.6151
R1806 B.n316 B.n91 10.6151
R1807 B.n320 B.n91 10.6151
R1808 B.n321 B.n320 10.6151
R1809 B.n322 B.n321 10.6151
R1810 B.n322 B.n89 10.6151
R1811 B.n326 B.n89 10.6151
R1812 B.n327 B.n326 10.6151
R1813 B.n328 B.n327 10.6151
R1814 B.n328 B.n87 10.6151
R1815 B.n573 B.n0 8.11757
R1816 B.n573 B.n1 8.11757
R1817 B.n473 B.n38 6.5566
R1818 B.n461 B.n460 6.5566
R1819 B.n248 B.n247 6.5566
R1820 B.n261 B.n260 6.5566
R1821 B.n38 B.n34 4.05904
R1822 B.n460 B.n459 4.05904
R1823 B.n247 B.n246 4.05904
R1824 B.n262 B.n261 4.05904
R1825 VP.n4 VP.t0 830.207
R1826 VP.n10 VP.t2 809.225
R1827 VP.n1 VP.t4 809.225
R1828 VP.n15 VP.t3 809.225
R1829 VP.n16 VP.t6 809.225
R1830 VP.n8 VP.t7 809.225
R1831 VP.n7 VP.t1 809.225
R1832 VP.n3 VP.t5 809.225
R1833 VP.n17 VP.n16 161.3
R1834 VP.n6 VP.n5 161.3
R1835 VP.n7 VP.n2 161.3
R1836 VP.n9 VP.n8 161.3
R1837 VP.n15 VP.n0 161.3
R1838 VP.n14 VP.n13 161.3
R1839 VP.n12 VP.n1 161.3
R1840 VP.n11 VP.n10 161.3
R1841 VP.n5 VP.n4 70.4033
R1842 VP.n10 VP.n1 48.2005
R1843 VP.n16 VP.n15 48.2005
R1844 VP.n8 VP.n7 48.2005
R1845 VP.n11 VP.n9 41.9626
R1846 VP.n14 VP.n1 24.1005
R1847 VP.n15 VP.n14 24.1005
R1848 VP.n6 VP.n3 24.1005
R1849 VP.n7 VP.n6 24.1005
R1850 VP.n4 VP.n3 20.9576
R1851 VP.n5 VP.n2 0.189894
R1852 VP.n9 VP.n2 0.189894
R1853 VP.n12 VP.n11 0.189894
R1854 VP.n13 VP.n12 0.189894
R1855 VP.n13 VP.n0 0.189894
R1856 VP.n17 VP.n0 0.189894
R1857 VP VP.n17 0.0516364
R1858 VDD1 VDD1.n0 70.7359
R1859 VDD1.n3 VDD1.n2 70.6222
R1860 VDD1.n3 VDD1.n1 70.6222
R1861 VDD1.n5 VDD1.n4 70.3413
R1862 VDD1.n5 VDD1.n3 38.9276
R1863 VDD1.n4 VDD1.t6 2.41543
R1864 VDD1.n4 VDD1.t0 2.41543
R1865 VDD1.n0 VDD1.t7 2.41543
R1866 VDD1.n0 VDD1.t2 2.41543
R1867 VDD1.n2 VDD1.t4 2.41543
R1868 VDD1.n2 VDD1.t1 2.41543
R1869 VDD1.n1 VDD1.t5 2.41543
R1870 VDD1.n1 VDD1.t3 2.41543
R1871 VDD1 VDD1.n5 0.278517
C0 VTAIL VP 4.38846f
C1 w_n1750_n3660# VDD1 1.24059f
C2 w_n1750_n3660# VDD2 1.26507f
C3 VN VP 5.30727f
C4 B VP 1.09585f
C5 VDD1 VP 4.91494f
C6 VN VTAIL 4.37436f
C7 VTAIL B 4.00434f
C8 VDD2 VP 0.290591f
C9 VTAIL VDD1 15.022f
C10 VN B 0.737095f
C11 VTAIL VDD2 15.061999f
C12 VN VDD1 0.147544f
C13 VDD1 B 1.03301f
C14 VN VDD2 4.7722f
C15 VDD2 B 1.06196f
C16 w_n1750_n3660# VP 3.2144f
C17 VDD1 VDD2 0.704224f
C18 w_n1750_n3660# VTAIL 4.61445f
C19 w_n1750_n3660# VN 2.99355f
C20 w_n1750_n3660# B 7.23626f
C21 VDD2 VSUBS 1.396926f
C22 VDD1 VSUBS 1.654983f
C23 VTAIL VSUBS 0.862452f
C24 VN VSUBS 4.67674f
C25 VP VSUBS 1.447582f
C26 B VSUBS 2.724325f
C27 w_n1750_n3660# VSUBS 78.687004f
C28 VDD1.t7 VSUBS 0.31968f
C29 VDD1.t2 VSUBS 0.31968f
C30 VDD1.n0 VSUBS 2.53546f
C31 VDD1.t5 VSUBS 0.31968f
C32 VDD1.t3 VSUBS 0.31968f
C33 VDD1.n1 VSUBS 2.53429f
C34 VDD1.t4 VSUBS 0.31968f
C35 VDD1.t1 VSUBS 0.31968f
C36 VDD1.n2 VSUBS 2.53429f
C37 VDD1.n3 VSUBS 3.28351f
C38 VDD1.t6 VSUBS 0.31968f
C39 VDD1.t0 VSUBS 0.31968f
C40 VDD1.n4 VSUBS 2.53153f
C41 VDD1.n5 VSUBS 3.16012f
C42 VP.n0 VSUBS 0.062382f
C43 VP.t4 VSUBS 1.07595f
C44 VP.n1 VSUBS 0.434048f
C45 VP.n2 VSUBS 0.062382f
C46 VP.t7 VSUBS 1.07595f
C47 VP.t1 VSUBS 1.07595f
C48 VP.t5 VSUBS 1.07595f
C49 VP.n3 VSUBS 0.434048f
C50 VP.t0 VSUBS 1.08677f
C51 VP.n4 VSUBS 0.417342f
C52 VP.n5 VSUBS 0.197849f
C53 VP.n6 VSUBS 0.014156f
C54 VP.n7 VSUBS 0.434048f
C55 VP.n8 VSUBS 0.427702f
C56 VP.n9 VSUBS 2.5712f
C57 VP.t2 VSUBS 1.07595f
C58 VP.n10 VSUBS 0.427702f
C59 VP.n11 VSUBS 2.62449f
C60 VP.n12 VSUBS 0.062382f
C61 VP.n13 VSUBS 0.062382f
C62 VP.n14 VSUBS 0.014156f
C63 VP.t3 VSUBS 1.07595f
C64 VP.n15 VSUBS 0.434048f
C65 VP.t6 VSUBS 1.07595f
C66 VP.n16 VSUBS 0.427702f
C67 VP.n17 VSUBS 0.048344f
C68 B.n0 VSUBS 0.007317f
C69 B.n1 VSUBS 0.007317f
C70 B.n2 VSUBS 0.010821f
C71 B.n3 VSUBS 0.008292f
C72 B.n4 VSUBS 0.008292f
C73 B.n5 VSUBS 0.008292f
C74 B.n6 VSUBS 0.008292f
C75 B.n7 VSUBS 0.008292f
C76 B.n8 VSUBS 0.008292f
C77 B.n9 VSUBS 0.008292f
C78 B.n10 VSUBS 0.008292f
C79 B.n11 VSUBS 0.020146f
C80 B.n12 VSUBS 0.008292f
C81 B.n13 VSUBS 0.008292f
C82 B.n14 VSUBS 0.008292f
C83 B.n15 VSUBS 0.008292f
C84 B.n16 VSUBS 0.008292f
C85 B.n17 VSUBS 0.008292f
C86 B.n18 VSUBS 0.008292f
C87 B.n19 VSUBS 0.008292f
C88 B.n20 VSUBS 0.008292f
C89 B.n21 VSUBS 0.008292f
C90 B.n22 VSUBS 0.008292f
C91 B.n23 VSUBS 0.008292f
C92 B.n24 VSUBS 0.008292f
C93 B.n25 VSUBS 0.008292f
C94 B.n26 VSUBS 0.008292f
C95 B.n27 VSUBS 0.008292f
C96 B.n28 VSUBS 0.008292f
C97 B.n29 VSUBS 0.008292f
C98 B.n30 VSUBS 0.008292f
C99 B.n31 VSUBS 0.008292f
C100 B.n32 VSUBS 0.008292f
C101 B.n33 VSUBS 0.008292f
C102 B.n34 VSUBS 0.005732f
C103 B.n35 VSUBS 0.008292f
C104 B.t7 VSUBS 0.289074f
C105 B.t8 VSUBS 0.299933f
C106 B.t6 VSUBS 0.286195f
C107 B.n36 VSUBS 0.376784f
C108 B.n37 VSUBS 0.311222f
C109 B.n38 VSUBS 0.019213f
C110 B.n39 VSUBS 0.008292f
C111 B.n40 VSUBS 0.008292f
C112 B.n41 VSUBS 0.008292f
C113 B.n42 VSUBS 0.008292f
C114 B.t4 VSUBS 0.289078f
C115 B.t5 VSUBS 0.299937f
C116 B.t3 VSUBS 0.286195f
C117 B.n43 VSUBS 0.376781f
C118 B.n44 VSUBS 0.311218f
C119 B.n45 VSUBS 0.008292f
C120 B.n46 VSUBS 0.008292f
C121 B.n47 VSUBS 0.008292f
C122 B.n48 VSUBS 0.008292f
C123 B.n49 VSUBS 0.008292f
C124 B.n50 VSUBS 0.008292f
C125 B.n51 VSUBS 0.008292f
C126 B.n52 VSUBS 0.008292f
C127 B.n53 VSUBS 0.008292f
C128 B.n54 VSUBS 0.008292f
C129 B.n55 VSUBS 0.008292f
C130 B.n56 VSUBS 0.008292f
C131 B.n57 VSUBS 0.008292f
C132 B.n58 VSUBS 0.008292f
C133 B.n59 VSUBS 0.008292f
C134 B.n60 VSUBS 0.008292f
C135 B.n61 VSUBS 0.008292f
C136 B.n62 VSUBS 0.008292f
C137 B.n63 VSUBS 0.008292f
C138 B.n64 VSUBS 0.008292f
C139 B.n65 VSUBS 0.008292f
C140 B.n66 VSUBS 0.008292f
C141 B.n67 VSUBS 0.020146f
C142 B.n68 VSUBS 0.008292f
C143 B.n69 VSUBS 0.008292f
C144 B.n70 VSUBS 0.008292f
C145 B.n71 VSUBS 0.008292f
C146 B.n72 VSUBS 0.008292f
C147 B.n73 VSUBS 0.008292f
C148 B.n74 VSUBS 0.008292f
C149 B.n75 VSUBS 0.008292f
C150 B.n76 VSUBS 0.008292f
C151 B.n77 VSUBS 0.008292f
C152 B.n78 VSUBS 0.008292f
C153 B.n79 VSUBS 0.008292f
C154 B.n80 VSUBS 0.008292f
C155 B.n81 VSUBS 0.008292f
C156 B.n82 VSUBS 0.008292f
C157 B.n83 VSUBS 0.008292f
C158 B.n84 VSUBS 0.008292f
C159 B.n85 VSUBS 0.008292f
C160 B.n86 VSUBS 0.008292f
C161 B.n87 VSUBS 0.019925f
C162 B.n88 VSUBS 0.008292f
C163 B.n89 VSUBS 0.008292f
C164 B.n90 VSUBS 0.008292f
C165 B.n91 VSUBS 0.008292f
C166 B.n92 VSUBS 0.008292f
C167 B.n93 VSUBS 0.008292f
C168 B.n94 VSUBS 0.008292f
C169 B.n95 VSUBS 0.008292f
C170 B.n96 VSUBS 0.008292f
C171 B.n97 VSUBS 0.008292f
C172 B.n98 VSUBS 0.008292f
C173 B.n99 VSUBS 0.008292f
C174 B.n100 VSUBS 0.008292f
C175 B.n101 VSUBS 0.008292f
C176 B.n102 VSUBS 0.008292f
C177 B.n103 VSUBS 0.008292f
C178 B.n104 VSUBS 0.008292f
C179 B.n105 VSUBS 0.008292f
C180 B.n106 VSUBS 0.008292f
C181 B.n107 VSUBS 0.008292f
C182 B.n108 VSUBS 0.008292f
C183 B.n109 VSUBS 0.008292f
C184 B.n110 VSUBS 0.008292f
C185 B.t2 VSUBS 0.289078f
C186 B.t1 VSUBS 0.299937f
C187 B.t0 VSUBS 0.286195f
C188 B.n111 VSUBS 0.376781f
C189 B.n112 VSUBS 0.311218f
C190 B.n113 VSUBS 0.008292f
C191 B.n114 VSUBS 0.008292f
C192 B.n115 VSUBS 0.008292f
C193 B.n116 VSUBS 0.008292f
C194 B.t11 VSUBS 0.289074f
C195 B.t10 VSUBS 0.299933f
C196 B.t9 VSUBS 0.286195f
C197 B.n117 VSUBS 0.376784f
C198 B.n118 VSUBS 0.311222f
C199 B.n119 VSUBS 0.008292f
C200 B.n120 VSUBS 0.008292f
C201 B.n121 VSUBS 0.008292f
C202 B.n122 VSUBS 0.008292f
C203 B.n123 VSUBS 0.008292f
C204 B.n124 VSUBS 0.008292f
C205 B.n125 VSUBS 0.008292f
C206 B.n126 VSUBS 0.008292f
C207 B.n127 VSUBS 0.008292f
C208 B.n128 VSUBS 0.008292f
C209 B.n129 VSUBS 0.008292f
C210 B.n130 VSUBS 0.008292f
C211 B.n131 VSUBS 0.008292f
C212 B.n132 VSUBS 0.008292f
C213 B.n133 VSUBS 0.008292f
C214 B.n134 VSUBS 0.008292f
C215 B.n135 VSUBS 0.008292f
C216 B.n136 VSUBS 0.008292f
C217 B.n137 VSUBS 0.008292f
C218 B.n138 VSUBS 0.008292f
C219 B.n139 VSUBS 0.008292f
C220 B.n140 VSUBS 0.008292f
C221 B.n141 VSUBS 0.020829f
C222 B.n142 VSUBS 0.008292f
C223 B.n143 VSUBS 0.008292f
C224 B.n144 VSUBS 0.008292f
C225 B.n145 VSUBS 0.008292f
C226 B.n146 VSUBS 0.008292f
C227 B.n147 VSUBS 0.008292f
C228 B.n148 VSUBS 0.008292f
C229 B.n149 VSUBS 0.008292f
C230 B.n150 VSUBS 0.008292f
C231 B.n151 VSUBS 0.008292f
C232 B.n152 VSUBS 0.008292f
C233 B.n153 VSUBS 0.008292f
C234 B.n154 VSUBS 0.008292f
C235 B.n155 VSUBS 0.008292f
C236 B.n156 VSUBS 0.008292f
C237 B.n157 VSUBS 0.008292f
C238 B.n158 VSUBS 0.008292f
C239 B.n159 VSUBS 0.008292f
C240 B.n160 VSUBS 0.008292f
C241 B.n161 VSUBS 0.008292f
C242 B.n162 VSUBS 0.008292f
C243 B.n163 VSUBS 0.008292f
C244 B.n164 VSUBS 0.008292f
C245 B.n165 VSUBS 0.008292f
C246 B.n166 VSUBS 0.008292f
C247 B.n167 VSUBS 0.008292f
C248 B.n168 VSUBS 0.008292f
C249 B.n169 VSUBS 0.008292f
C250 B.n170 VSUBS 0.008292f
C251 B.n171 VSUBS 0.008292f
C252 B.n172 VSUBS 0.008292f
C253 B.n173 VSUBS 0.008292f
C254 B.n174 VSUBS 0.008292f
C255 B.n175 VSUBS 0.008292f
C256 B.n176 VSUBS 0.020146f
C257 B.n177 VSUBS 0.020146f
C258 B.n178 VSUBS 0.020829f
C259 B.n179 VSUBS 0.008292f
C260 B.n180 VSUBS 0.008292f
C261 B.n181 VSUBS 0.008292f
C262 B.n182 VSUBS 0.008292f
C263 B.n183 VSUBS 0.008292f
C264 B.n184 VSUBS 0.008292f
C265 B.n185 VSUBS 0.008292f
C266 B.n186 VSUBS 0.008292f
C267 B.n187 VSUBS 0.008292f
C268 B.n188 VSUBS 0.008292f
C269 B.n189 VSUBS 0.008292f
C270 B.n190 VSUBS 0.008292f
C271 B.n191 VSUBS 0.008292f
C272 B.n192 VSUBS 0.008292f
C273 B.n193 VSUBS 0.008292f
C274 B.n194 VSUBS 0.008292f
C275 B.n195 VSUBS 0.008292f
C276 B.n196 VSUBS 0.008292f
C277 B.n197 VSUBS 0.008292f
C278 B.n198 VSUBS 0.008292f
C279 B.n199 VSUBS 0.008292f
C280 B.n200 VSUBS 0.008292f
C281 B.n201 VSUBS 0.008292f
C282 B.n202 VSUBS 0.008292f
C283 B.n203 VSUBS 0.008292f
C284 B.n204 VSUBS 0.008292f
C285 B.n205 VSUBS 0.008292f
C286 B.n206 VSUBS 0.008292f
C287 B.n207 VSUBS 0.008292f
C288 B.n208 VSUBS 0.008292f
C289 B.n209 VSUBS 0.008292f
C290 B.n210 VSUBS 0.008292f
C291 B.n211 VSUBS 0.008292f
C292 B.n212 VSUBS 0.008292f
C293 B.n213 VSUBS 0.008292f
C294 B.n214 VSUBS 0.008292f
C295 B.n215 VSUBS 0.008292f
C296 B.n216 VSUBS 0.008292f
C297 B.n217 VSUBS 0.008292f
C298 B.n218 VSUBS 0.008292f
C299 B.n219 VSUBS 0.008292f
C300 B.n220 VSUBS 0.008292f
C301 B.n221 VSUBS 0.008292f
C302 B.n222 VSUBS 0.008292f
C303 B.n223 VSUBS 0.008292f
C304 B.n224 VSUBS 0.008292f
C305 B.n225 VSUBS 0.008292f
C306 B.n226 VSUBS 0.008292f
C307 B.n227 VSUBS 0.008292f
C308 B.n228 VSUBS 0.008292f
C309 B.n229 VSUBS 0.008292f
C310 B.n230 VSUBS 0.008292f
C311 B.n231 VSUBS 0.008292f
C312 B.n232 VSUBS 0.008292f
C313 B.n233 VSUBS 0.008292f
C314 B.n234 VSUBS 0.008292f
C315 B.n235 VSUBS 0.008292f
C316 B.n236 VSUBS 0.008292f
C317 B.n237 VSUBS 0.008292f
C318 B.n238 VSUBS 0.008292f
C319 B.n239 VSUBS 0.008292f
C320 B.n240 VSUBS 0.008292f
C321 B.n241 VSUBS 0.008292f
C322 B.n242 VSUBS 0.008292f
C323 B.n243 VSUBS 0.008292f
C324 B.n244 VSUBS 0.008292f
C325 B.n245 VSUBS 0.008292f
C326 B.n246 VSUBS 0.005732f
C327 B.n247 VSUBS 0.019213f
C328 B.n248 VSUBS 0.006707f
C329 B.n249 VSUBS 0.008292f
C330 B.n250 VSUBS 0.008292f
C331 B.n251 VSUBS 0.008292f
C332 B.n252 VSUBS 0.008292f
C333 B.n253 VSUBS 0.008292f
C334 B.n254 VSUBS 0.008292f
C335 B.n255 VSUBS 0.008292f
C336 B.n256 VSUBS 0.008292f
C337 B.n257 VSUBS 0.008292f
C338 B.n258 VSUBS 0.008292f
C339 B.n259 VSUBS 0.008292f
C340 B.n260 VSUBS 0.006707f
C341 B.n261 VSUBS 0.019213f
C342 B.n262 VSUBS 0.005732f
C343 B.n263 VSUBS 0.008292f
C344 B.n264 VSUBS 0.008292f
C345 B.n265 VSUBS 0.008292f
C346 B.n266 VSUBS 0.008292f
C347 B.n267 VSUBS 0.008292f
C348 B.n268 VSUBS 0.008292f
C349 B.n269 VSUBS 0.008292f
C350 B.n270 VSUBS 0.008292f
C351 B.n271 VSUBS 0.008292f
C352 B.n272 VSUBS 0.008292f
C353 B.n273 VSUBS 0.008292f
C354 B.n274 VSUBS 0.008292f
C355 B.n275 VSUBS 0.008292f
C356 B.n276 VSUBS 0.008292f
C357 B.n277 VSUBS 0.008292f
C358 B.n278 VSUBS 0.008292f
C359 B.n279 VSUBS 0.008292f
C360 B.n280 VSUBS 0.008292f
C361 B.n281 VSUBS 0.008292f
C362 B.n282 VSUBS 0.008292f
C363 B.n283 VSUBS 0.008292f
C364 B.n284 VSUBS 0.008292f
C365 B.n285 VSUBS 0.008292f
C366 B.n286 VSUBS 0.008292f
C367 B.n287 VSUBS 0.008292f
C368 B.n288 VSUBS 0.008292f
C369 B.n289 VSUBS 0.008292f
C370 B.n290 VSUBS 0.008292f
C371 B.n291 VSUBS 0.008292f
C372 B.n292 VSUBS 0.008292f
C373 B.n293 VSUBS 0.008292f
C374 B.n294 VSUBS 0.008292f
C375 B.n295 VSUBS 0.008292f
C376 B.n296 VSUBS 0.008292f
C377 B.n297 VSUBS 0.008292f
C378 B.n298 VSUBS 0.008292f
C379 B.n299 VSUBS 0.008292f
C380 B.n300 VSUBS 0.008292f
C381 B.n301 VSUBS 0.008292f
C382 B.n302 VSUBS 0.008292f
C383 B.n303 VSUBS 0.008292f
C384 B.n304 VSUBS 0.008292f
C385 B.n305 VSUBS 0.008292f
C386 B.n306 VSUBS 0.008292f
C387 B.n307 VSUBS 0.008292f
C388 B.n308 VSUBS 0.008292f
C389 B.n309 VSUBS 0.008292f
C390 B.n310 VSUBS 0.008292f
C391 B.n311 VSUBS 0.008292f
C392 B.n312 VSUBS 0.008292f
C393 B.n313 VSUBS 0.008292f
C394 B.n314 VSUBS 0.008292f
C395 B.n315 VSUBS 0.008292f
C396 B.n316 VSUBS 0.008292f
C397 B.n317 VSUBS 0.008292f
C398 B.n318 VSUBS 0.008292f
C399 B.n319 VSUBS 0.008292f
C400 B.n320 VSUBS 0.008292f
C401 B.n321 VSUBS 0.008292f
C402 B.n322 VSUBS 0.008292f
C403 B.n323 VSUBS 0.008292f
C404 B.n324 VSUBS 0.008292f
C405 B.n325 VSUBS 0.008292f
C406 B.n326 VSUBS 0.008292f
C407 B.n327 VSUBS 0.008292f
C408 B.n328 VSUBS 0.008292f
C409 B.n329 VSUBS 0.008292f
C410 B.n330 VSUBS 0.020829f
C411 B.n331 VSUBS 0.020146f
C412 B.n332 VSUBS 0.021049f
C413 B.n333 VSUBS 0.008292f
C414 B.n334 VSUBS 0.008292f
C415 B.n335 VSUBS 0.008292f
C416 B.n336 VSUBS 0.008292f
C417 B.n337 VSUBS 0.008292f
C418 B.n338 VSUBS 0.008292f
C419 B.n339 VSUBS 0.008292f
C420 B.n340 VSUBS 0.008292f
C421 B.n341 VSUBS 0.008292f
C422 B.n342 VSUBS 0.008292f
C423 B.n343 VSUBS 0.008292f
C424 B.n344 VSUBS 0.008292f
C425 B.n345 VSUBS 0.008292f
C426 B.n346 VSUBS 0.008292f
C427 B.n347 VSUBS 0.008292f
C428 B.n348 VSUBS 0.008292f
C429 B.n349 VSUBS 0.008292f
C430 B.n350 VSUBS 0.008292f
C431 B.n351 VSUBS 0.008292f
C432 B.n352 VSUBS 0.008292f
C433 B.n353 VSUBS 0.008292f
C434 B.n354 VSUBS 0.008292f
C435 B.n355 VSUBS 0.008292f
C436 B.n356 VSUBS 0.008292f
C437 B.n357 VSUBS 0.008292f
C438 B.n358 VSUBS 0.008292f
C439 B.n359 VSUBS 0.008292f
C440 B.n360 VSUBS 0.008292f
C441 B.n361 VSUBS 0.008292f
C442 B.n362 VSUBS 0.008292f
C443 B.n363 VSUBS 0.008292f
C444 B.n364 VSUBS 0.008292f
C445 B.n365 VSUBS 0.008292f
C446 B.n366 VSUBS 0.008292f
C447 B.n367 VSUBS 0.008292f
C448 B.n368 VSUBS 0.008292f
C449 B.n369 VSUBS 0.008292f
C450 B.n370 VSUBS 0.008292f
C451 B.n371 VSUBS 0.008292f
C452 B.n372 VSUBS 0.008292f
C453 B.n373 VSUBS 0.008292f
C454 B.n374 VSUBS 0.008292f
C455 B.n375 VSUBS 0.008292f
C456 B.n376 VSUBS 0.008292f
C457 B.n377 VSUBS 0.008292f
C458 B.n378 VSUBS 0.008292f
C459 B.n379 VSUBS 0.008292f
C460 B.n380 VSUBS 0.008292f
C461 B.n381 VSUBS 0.008292f
C462 B.n382 VSUBS 0.008292f
C463 B.n383 VSUBS 0.008292f
C464 B.n384 VSUBS 0.008292f
C465 B.n385 VSUBS 0.008292f
C466 B.n386 VSUBS 0.008292f
C467 B.n387 VSUBS 0.008292f
C468 B.n388 VSUBS 0.008292f
C469 B.n389 VSUBS 0.008292f
C470 B.n390 VSUBS 0.020146f
C471 B.n391 VSUBS 0.020829f
C472 B.n392 VSUBS 0.020829f
C473 B.n393 VSUBS 0.008292f
C474 B.n394 VSUBS 0.008292f
C475 B.n395 VSUBS 0.008292f
C476 B.n396 VSUBS 0.008292f
C477 B.n397 VSUBS 0.008292f
C478 B.n398 VSUBS 0.008292f
C479 B.n399 VSUBS 0.008292f
C480 B.n400 VSUBS 0.008292f
C481 B.n401 VSUBS 0.008292f
C482 B.n402 VSUBS 0.008292f
C483 B.n403 VSUBS 0.008292f
C484 B.n404 VSUBS 0.008292f
C485 B.n405 VSUBS 0.008292f
C486 B.n406 VSUBS 0.008292f
C487 B.n407 VSUBS 0.008292f
C488 B.n408 VSUBS 0.008292f
C489 B.n409 VSUBS 0.008292f
C490 B.n410 VSUBS 0.008292f
C491 B.n411 VSUBS 0.008292f
C492 B.n412 VSUBS 0.008292f
C493 B.n413 VSUBS 0.008292f
C494 B.n414 VSUBS 0.008292f
C495 B.n415 VSUBS 0.008292f
C496 B.n416 VSUBS 0.008292f
C497 B.n417 VSUBS 0.008292f
C498 B.n418 VSUBS 0.008292f
C499 B.n419 VSUBS 0.008292f
C500 B.n420 VSUBS 0.008292f
C501 B.n421 VSUBS 0.008292f
C502 B.n422 VSUBS 0.008292f
C503 B.n423 VSUBS 0.008292f
C504 B.n424 VSUBS 0.008292f
C505 B.n425 VSUBS 0.008292f
C506 B.n426 VSUBS 0.008292f
C507 B.n427 VSUBS 0.008292f
C508 B.n428 VSUBS 0.008292f
C509 B.n429 VSUBS 0.008292f
C510 B.n430 VSUBS 0.008292f
C511 B.n431 VSUBS 0.008292f
C512 B.n432 VSUBS 0.008292f
C513 B.n433 VSUBS 0.008292f
C514 B.n434 VSUBS 0.008292f
C515 B.n435 VSUBS 0.008292f
C516 B.n436 VSUBS 0.008292f
C517 B.n437 VSUBS 0.008292f
C518 B.n438 VSUBS 0.008292f
C519 B.n439 VSUBS 0.008292f
C520 B.n440 VSUBS 0.008292f
C521 B.n441 VSUBS 0.008292f
C522 B.n442 VSUBS 0.008292f
C523 B.n443 VSUBS 0.008292f
C524 B.n444 VSUBS 0.008292f
C525 B.n445 VSUBS 0.008292f
C526 B.n446 VSUBS 0.008292f
C527 B.n447 VSUBS 0.008292f
C528 B.n448 VSUBS 0.008292f
C529 B.n449 VSUBS 0.008292f
C530 B.n450 VSUBS 0.008292f
C531 B.n451 VSUBS 0.008292f
C532 B.n452 VSUBS 0.008292f
C533 B.n453 VSUBS 0.008292f
C534 B.n454 VSUBS 0.008292f
C535 B.n455 VSUBS 0.008292f
C536 B.n456 VSUBS 0.008292f
C537 B.n457 VSUBS 0.008292f
C538 B.n458 VSUBS 0.008292f
C539 B.n459 VSUBS 0.005732f
C540 B.n460 VSUBS 0.019213f
C541 B.n461 VSUBS 0.006707f
C542 B.n462 VSUBS 0.008292f
C543 B.n463 VSUBS 0.008292f
C544 B.n464 VSUBS 0.008292f
C545 B.n465 VSUBS 0.008292f
C546 B.n466 VSUBS 0.008292f
C547 B.n467 VSUBS 0.008292f
C548 B.n468 VSUBS 0.008292f
C549 B.n469 VSUBS 0.008292f
C550 B.n470 VSUBS 0.008292f
C551 B.n471 VSUBS 0.008292f
C552 B.n472 VSUBS 0.008292f
C553 B.n473 VSUBS 0.006707f
C554 B.n474 VSUBS 0.008292f
C555 B.n475 VSUBS 0.008292f
C556 B.n476 VSUBS 0.008292f
C557 B.n477 VSUBS 0.008292f
C558 B.n478 VSUBS 0.008292f
C559 B.n479 VSUBS 0.008292f
C560 B.n480 VSUBS 0.008292f
C561 B.n481 VSUBS 0.008292f
C562 B.n482 VSUBS 0.008292f
C563 B.n483 VSUBS 0.008292f
C564 B.n484 VSUBS 0.008292f
C565 B.n485 VSUBS 0.008292f
C566 B.n486 VSUBS 0.008292f
C567 B.n487 VSUBS 0.008292f
C568 B.n488 VSUBS 0.008292f
C569 B.n489 VSUBS 0.008292f
C570 B.n490 VSUBS 0.008292f
C571 B.n491 VSUBS 0.008292f
C572 B.n492 VSUBS 0.008292f
C573 B.n493 VSUBS 0.008292f
C574 B.n494 VSUBS 0.008292f
C575 B.n495 VSUBS 0.008292f
C576 B.n496 VSUBS 0.008292f
C577 B.n497 VSUBS 0.008292f
C578 B.n498 VSUBS 0.008292f
C579 B.n499 VSUBS 0.008292f
C580 B.n500 VSUBS 0.008292f
C581 B.n501 VSUBS 0.008292f
C582 B.n502 VSUBS 0.008292f
C583 B.n503 VSUBS 0.008292f
C584 B.n504 VSUBS 0.008292f
C585 B.n505 VSUBS 0.008292f
C586 B.n506 VSUBS 0.008292f
C587 B.n507 VSUBS 0.008292f
C588 B.n508 VSUBS 0.008292f
C589 B.n509 VSUBS 0.008292f
C590 B.n510 VSUBS 0.008292f
C591 B.n511 VSUBS 0.008292f
C592 B.n512 VSUBS 0.008292f
C593 B.n513 VSUBS 0.008292f
C594 B.n514 VSUBS 0.008292f
C595 B.n515 VSUBS 0.008292f
C596 B.n516 VSUBS 0.008292f
C597 B.n517 VSUBS 0.008292f
C598 B.n518 VSUBS 0.008292f
C599 B.n519 VSUBS 0.008292f
C600 B.n520 VSUBS 0.008292f
C601 B.n521 VSUBS 0.008292f
C602 B.n522 VSUBS 0.008292f
C603 B.n523 VSUBS 0.008292f
C604 B.n524 VSUBS 0.008292f
C605 B.n525 VSUBS 0.008292f
C606 B.n526 VSUBS 0.008292f
C607 B.n527 VSUBS 0.008292f
C608 B.n528 VSUBS 0.008292f
C609 B.n529 VSUBS 0.008292f
C610 B.n530 VSUBS 0.008292f
C611 B.n531 VSUBS 0.008292f
C612 B.n532 VSUBS 0.008292f
C613 B.n533 VSUBS 0.008292f
C614 B.n534 VSUBS 0.008292f
C615 B.n535 VSUBS 0.008292f
C616 B.n536 VSUBS 0.008292f
C617 B.n537 VSUBS 0.008292f
C618 B.n538 VSUBS 0.008292f
C619 B.n539 VSUBS 0.008292f
C620 B.n540 VSUBS 0.008292f
C621 B.n541 VSUBS 0.008292f
C622 B.n542 VSUBS 0.020829f
C623 B.n543 VSUBS 0.020829f
C624 B.n544 VSUBS 0.020146f
C625 B.n545 VSUBS 0.008292f
C626 B.n546 VSUBS 0.008292f
C627 B.n547 VSUBS 0.008292f
C628 B.n548 VSUBS 0.008292f
C629 B.n549 VSUBS 0.008292f
C630 B.n550 VSUBS 0.008292f
C631 B.n551 VSUBS 0.008292f
C632 B.n552 VSUBS 0.008292f
C633 B.n553 VSUBS 0.008292f
C634 B.n554 VSUBS 0.008292f
C635 B.n555 VSUBS 0.008292f
C636 B.n556 VSUBS 0.008292f
C637 B.n557 VSUBS 0.008292f
C638 B.n558 VSUBS 0.008292f
C639 B.n559 VSUBS 0.008292f
C640 B.n560 VSUBS 0.008292f
C641 B.n561 VSUBS 0.008292f
C642 B.n562 VSUBS 0.008292f
C643 B.n563 VSUBS 0.008292f
C644 B.n564 VSUBS 0.008292f
C645 B.n565 VSUBS 0.008292f
C646 B.n566 VSUBS 0.008292f
C647 B.n567 VSUBS 0.008292f
C648 B.n568 VSUBS 0.008292f
C649 B.n569 VSUBS 0.008292f
C650 B.n570 VSUBS 0.008292f
C651 B.n571 VSUBS 0.010821f
C652 B.n572 VSUBS 0.011527f
C653 B.n573 VSUBS 0.022923f
C654 VDD2.t4 VSUBS 0.321473f
C655 VDD2.t5 VSUBS 0.321473f
C656 VDD2.n0 VSUBS 2.54851f
C657 VDD2.t6 VSUBS 0.321473f
C658 VDD2.t7 VSUBS 0.321473f
C659 VDD2.n1 VSUBS 2.54851f
C660 VDD2.n2 VSUBS 3.23728f
C661 VDD2.t3 VSUBS 0.321473f
C662 VDD2.t1 VSUBS 0.321473f
C663 VDD2.n3 VSUBS 2.54575f
C664 VDD2.n4 VSUBS 3.14218f
C665 VDD2.t0 VSUBS 0.321473f
C666 VDD2.t2 VSUBS 0.321473f
C667 VDD2.n5 VSUBS 2.54847f
C668 VTAIL.t9 VSUBS 0.280817f
C669 VTAIL.t15 VSUBS 0.280817f
C670 VTAIL.n0 VSUBS 2.06514f
C671 VTAIL.n1 VSUBS 0.700322f
C672 VTAIL.n2 VSUBS 0.028675f
C673 VTAIL.n3 VSUBS 0.026401f
C674 VTAIL.n4 VSUBS 0.014187f
C675 VTAIL.n5 VSUBS 0.033533f
C676 VTAIL.n6 VSUBS 0.015021f
C677 VTAIL.n7 VSUBS 0.026401f
C678 VTAIL.n8 VSUBS 0.014187f
C679 VTAIL.n9 VSUBS 0.033533f
C680 VTAIL.n10 VSUBS 0.015021f
C681 VTAIL.n11 VSUBS 0.026401f
C682 VTAIL.n12 VSUBS 0.014187f
C683 VTAIL.n13 VSUBS 0.033533f
C684 VTAIL.n14 VSUBS 0.014604f
C685 VTAIL.n15 VSUBS 0.026401f
C686 VTAIL.n16 VSUBS 0.015021f
C687 VTAIL.n17 VSUBS 0.033533f
C688 VTAIL.n18 VSUBS 0.015021f
C689 VTAIL.n19 VSUBS 0.026401f
C690 VTAIL.n20 VSUBS 0.014187f
C691 VTAIL.n21 VSUBS 0.033533f
C692 VTAIL.n22 VSUBS 0.015021f
C693 VTAIL.n23 VSUBS 1.46607f
C694 VTAIL.n24 VSUBS 0.014187f
C695 VTAIL.t14 VSUBS 0.072386f
C696 VTAIL.n25 VSUBS 0.225351f
C697 VTAIL.n26 VSUBS 0.025225f
C698 VTAIL.n27 VSUBS 0.025149f
C699 VTAIL.n28 VSUBS 0.033533f
C700 VTAIL.n29 VSUBS 0.015021f
C701 VTAIL.n30 VSUBS 0.014187f
C702 VTAIL.n31 VSUBS 0.026401f
C703 VTAIL.n32 VSUBS 0.026401f
C704 VTAIL.n33 VSUBS 0.014187f
C705 VTAIL.n34 VSUBS 0.015021f
C706 VTAIL.n35 VSUBS 0.033533f
C707 VTAIL.n36 VSUBS 0.033533f
C708 VTAIL.n37 VSUBS 0.015021f
C709 VTAIL.n38 VSUBS 0.014187f
C710 VTAIL.n39 VSUBS 0.026401f
C711 VTAIL.n40 VSUBS 0.026401f
C712 VTAIL.n41 VSUBS 0.014187f
C713 VTAIL.n42 VSUBS 0.014187f
C714 VTAIL.n43 VSUBS 0.015021f
C715 VTAIL.n44 VSUBS 0.033533f
C716 VTAIL.n45 VSUBS 0.033533f
C717 VTAIL.n46 VSUBS 0.033533f
C718 VTAIL.n47 VSUBS 0.014604f
C719 VTAIL.n48 VSUBS 0.014187f
C720 VTAIL.n49 VSUBS 0.026401f
C721 VTAIL.n50 VSUBS 0.026401f
C722 VTAIL.n51 VSUBS 0.014187f
C723 VTAIL.n52 VSUBS 0.015021f
C724 VTAIL.n53 VSUBS 0.033533f
C725 VTAIL.n54 VSUBS 0.033533f
C726 VTAIL.n55 VSUBS 0.015021f
C727 VTAIL.n56 VSUBS 0.014187f
C728 VTAIL.n57 VSUBS 0.026401f
C729 VTAIL.n58 VSUBS 0.026401f
C730 VTAIL.n59 VSUBS 0.014187f
C731 VTAIL.n60 VSUBS 0.015021f
C732 VTAIL.n61 VSUBS 0.033533f
C733 VTAIL.n62 VSUBS 0.033533f
C734 VTAIL.n63 VSUBS 0.015021f
C735 VTAIL.n64 VSUBS 0.014187f
C736 VTAIL.n65 VSUBS 0.026401f
C737 VTAIL.n66 VSUBS 0.026401f
C738 VTAIL.n67 VSUBS 0.014187f
C739 VTAIL.n68 VSUBS 0.015021f
C740 VTAIL.n69 VSUBS 0.033533f
C741 VTAIL.n70 VSUBS 0.08004f
C742 VTAIL.n71 VSUBS 0.015021f
C743 VTAIL.n72 VSUBS 0.014187f
C744 VTAIL.n73 VSUBS 0.057418f
C745 VTAIL.n74 VSUBS 0.040087f
C746 VTAIL.n75 VSUBS 0.117687f
C747 VTAIL.n76 VSUBS 0.028675f
C748 VTAIL.n77 VSUBS 0.026401f
C749 VTAIL.n78 VSUBS 0.014187f
C750 VTAIL.n79 VSUBS 0.033533f
C751 VTAIL.n80 VSUBS 0.015021f
C752 VTAIL.n81 VSUBS 0.026401f
C753 VTAIL.n82 VSUBS 0.014187f
C754 VTAIL.n83 VSUBS 0.033533f
C755 VTAIL.n84 VSUBS 0.015021f
C756 VTAIL.n85 VSUBS 0.026401f
C757 VTAIL.n86 VSUBS 0.014187f
C758 VTAIL.n87 VSUBS 0.033533f
C759 VTAIL.n88 VSUBS 0.014604f
C760 VTAIL.n89 VSUBS 0.026401f
C761 VTAIL.n90 VSUBS 0.015021f
C762 VTAIL.n91 VSUBS 0.033533f
C763 VTAIL.n92 VSUBS 0.015021f
C764 VTAIL.n93 VSUBS 0.026401f
C765 VTAIL.n94 VSUBS 0.014187f
C766 VTAIL.n95 VSUBS 0.033533f
C767 VTAIL.n96 VSUBS 0.015021f
C768 VTAIL.n97 VSUBS 1.46607f
C769 VTAIL.n98 VSUBS 0.014187f
C770 VTAIL.t7 VSUBS 0.072386f
C771 VTAIL.n99 VSUBS 0.225351f
C772 VTAIL.n100 VSUBS 0.025225f
C773 VTAIL.n101 VSUBS 0.025149f
C774 VTAIL.n102 VSUBS 0.033533f
C775 VTAIL.n103 VSUBS 0.015021f
C776 VTAIL.n104 VSUBS 0.014187f
C777 VTAIL.n105 VSUBS 0.026401f
C778 VTAIL.n106 VSUBS 0.026401f
C779 VTAIL.n107 VSUBS 0.014187f
C780 VTAIL.n108 VSUBS 0.015021f
C781 VTAIL.n109 VSUBS 0.033533f
C782 VTAIL.n110 VSUBS 0.033533f
C783 VTAIL.n111 VSUBS 0.015021f
C784 VTAIL.n112 VSUBS 0.014187f
C785 VTAIL.n113 VSUBS 0.026401f
C786 VTAIL.n114 VSUBS 0.026401f
C787 VTAIL.n115 VSUBS 0.014187f
C788 VTAIL.n116 VSUBS 0.014187f
C789 VTAIL.n117 VSUBS 0.015021f
C790 VTAIL.n118 VSUBS 0.033533f
C791 VTAIL.n119 VSUBS 0.033533f
C792 VTAIL.n120 VSUBS 0.033533f
C793 VTAIL.n121 VSUBS 0.014604f
C794 VTAIL.n122 VSUBS 0.014187f
C795 VTAIL.n123 VSUBS 0.026401f
C796 VTAIL.n124 VSUBS 0.026401f
C797 VTAIL.n125 VSUBS 0.014187f
C798 VTAIL.n126 VSUBS 0.015021f
C799 VTAIL.n127 VSUBS 0.033533f
C800 VTAIL.n128 VSUBS 0.033533f
C801 VTAIL.n129 VSUBS 0.015021f
C802 VTAIL.n130 VSUBS 0.014187f
C803 VTAIL.n131 VSUBS 0.026401f
C804 VTAIL.n132 VSUBS 0.026401f
C805 VTAIL.n133 VSUBS 0.014187f
C806 VTAIL.n134 VSUBS 0.015021f
C807 VTAIL.n135 VSUBS 0.033533f
C808 VTAIL.n136 VSUBS 0.033533f
C809 VTAIL.n137 VSUBS 0.015021f
C810 VTAIL.n138 VSUBS 0.014187f
C811 VTAIL.n139 VSUBS 0.026401f
C812 VTAIL.n140 VSUBS 0.026401f
C813 VTAIL.n141 VSUBS 0.014187f
C814 VTAIL.n142 VSUBS 0.015021f
C815 VTAIL.n143 VSUBS 0.033533f
C816 VTAIL.n144 VSUBS 0.08004f
C817 VTAIL.n145 VSUBS 0.015021f
C818 VTAIL.n146 VSUBS 0.014187f
C819 VTAIL.n147 VSUBS 0.057418f
C820 VTAIL.n148 VSUBS 0.040087f
C821 VTAIL.n149 VSUBS 0.117687f
C822 VTAIL.t2 VSUBS 0.280817f
C823 VTAIL.t4 VSUBS 0.280817f
C824 VTAIL.n150 VSUBS 2.06514f
C825 VTAIL.n151 VSUBS 0.752575f
C826 VTAIL.n152 VSUBS 0.028675f
C827 VTAIL.n153 VSUBS 0.026401f
C828 VTAIL.n154 VSUBS 0.014187f
C829 VTAIL.n155 VSUBS 0.033533f
C830 VTAIL.n156 VSUBS 0.015021f
C831 VTAIL.n157 VSUBS 0.026401f
C832 VTAIL.n158 VSUBS 0.014187f
C833 VTAIL.n159 VSUBS 0.033533f
C834 VTAIL.n160 VSUBS 0.015021f
C835 VTAIL.n161 VSUBS 0.026401f
C836 VTAIL.n162 VSUBS 0.014187f
C837 VTAIL.n163 VSUBS 0.033533f
C838 VTAIL.n164 VSUBS 0.014604f
C839 VTAIL.n165 VSUBS 0.026401f
C840 VTAIL.n166 VSUBS 0.015021f
C841 VTAIL.n167 VSUBS 0.033533f
C842 VTAIL.n168 VSUBS 0.015021f
C843 VTAIL.n169 VSUBS 0.026401f
C844 VTAIL.n170 VSUBS 0.014187f
C845 VTAIL.n171 VSUBS 0.033533f
C846 VTAIL.n172 VSUBS 0.015021f
C847 VTAIL.n173 VSUBS 1.46607f
C848 VTAIL.n174 VSUBS 0.014187f
C849 VTAIL.t5 VSUBS 0.072386f
C850 VTAIL.n175 VSUBS 0.225351f
C851 VTAIL.n176 VSUBS 0.025225f
C852 VTAIL.n177 VSUBS 0.025149f
C853 VTAIL.n178 VSUBS 0.033533f
C854 VTAIL.n179 VSUBS 0.015021f
C855 VTAIL.n180 VSUBS 0.014187f
C856 VTAIL.n181 VSUBS 0.026401f
C857 VTAIL.n182 VSUBS 0.026401f
C858 VTAIL.n183 VSUBS 0.014187f
C859 VTAIL.n184 VSUBS 0.015021f
C860 VTAIL.n185 VSUBS 0.033533f
C861 VTAIL.n186 VSUBS 0.033533f
C862 VTAIL.n187 VSUBS 0.015021f
C863 VTAIL.n188 VSUBS 0.014187f
C864 VTAIL.n189 VSUBS 0.026401f
C865 VTAIL.n190 VSUBS 0.026401f
C866 VTAIL.n191 VSUBS 0.014187f
C867 VTAIL.n192 VSUBS 0.014187f
C868 VTAIL.n193 VSUBS 0.015021f
C869 VTAIL.n194 VSUBS 0.033533f
C870 VTAIL.n195 VSUBS 0.033533f
C871 VTAIL.n196 VSUBS 0.033533f
C872 VTAIL.n197 VSUBS 0.014604f
C873 VTAIL.n198 VSUBS 0.014187f
C874 VTAIL.n199 VSUBS 0.026401f
C875 VTAIL.n200 VSUBS 0.026401f
C876 VTAIL.n201 VSUBS 0.014187f
C877 VTAIL.n202 VSUBS 0.015021f
C878 VTAIL.n203 VSUBS 0.033533f
C879 VTAIL.n204 VSUBS 0.033533f
C880 VTAIL.n205 VSUBS 0.015021f
C881 VTAIL.n206 VSUBS 0.014187f
C882 VTAIL.n207 VSUBS 0.026401f
C883 VTAIL.n208 VSUBS 0.026401f
C884 VTAIL.n209 VSUBS 0.014187f
C885 VTAIL.n210 VSUBS 0.015021f
C886 VTAIL.n211 VSUBS 0.033533f
C887 VTAIL.n212 VSUBS 0.033533f
C888 VTAIL.n213 VSUBS 0.015021f
C889 VTAIL.n214 VSUBS 0.014187f
C890 VTAIL.n215 VSUBS 0.026401f
C891 VTAIL.n216 VSUBS 0.026401f
C892 VTAIL.n217 VSUBS 0.014187f
C893 VTAIL.n218 VSUBS 0.015021f
C894 VTAIL.n219 VSUBS 0.033533f
C895 VTAIL.n220 VSUBS 0.08004f
C896 VTAIL.n221 VSUBS 0.015021f
C897 VTAIL.n222 VSUBS 0.014187f
C898 VTAIL.n223 VSUBS 0.057418f
C899 VTAIL.n224 VSUBS 0.040087f
C900 VTAIL.n225 VSUBS 1.48066f
C901 VTAIL.n226 VSUBS 0.028675f
C902 VTAIL.n227 VSUBS 0.026401f
C903 VTAIL.n228 VSUBS 0.014187f
C904 VTAIL.n229 VSUBS 0.033533f
C905 VTAIL.n230 VSUBS 0.015021f
C906 VTAIL.n231 VSUBS 0.026401f
C907 VTAIL.n232 VSUBS 0.014187f
C908 VTAIL.n233 VSUBS 0.033533f
C909 VTAIL.n234 VSUBS 0.015021f
C910 VTAIL.n235 VSUBS 0.026401f
C911 VTAIL.n236 VSUBS 0.014187f
C912 VTAIL.n237 VSUBS 0.033533f
C913 VTAIL.n238 VSUBS 0.014604f
C914 VTAIL.n239 VSUBS 0.026401f
C915 VTAIL.n240 VSUBS 0.014604f
C916 VTAIL.n241 VSUBS 0.014187f
C917 VTAIL.n242 VSUBS 0.033533f
C918 VTAIL.n243 VSUBS 0.033533f
C919 VTAIL.n244 VSUBS 0.015021f
C920 VTAIL.n245 VSUBS 0.026401f
C921 VTAIL.n246 VSUBS 0.014187f
C922 VTAIL.n247 VSUBS 0.033533f
C923 VTAIL.n248 VSUBS 0.015021f
C924 VTAIL.n249 VSUBS 1.46607f
C925 VTAIL.n250 VSUBS 0.014187f
C926 VTAIL.t13 VSUBS 0.072386f
C927 VTAIL.n251 VSUBS 0.225351f
C928 VTAIL.n252 VSUBS 0.025225f
C929 VTAIL.n253 VSUBS 0.025149f
C930 VTAIL.n254 VSUBS 0.033533f
C931 VTAIL.n255 VSUBS 0.015021f
C932 VTAIL.n256 VSUBS 0.014187f
C933 VTAIL.n257 VSUBS 0.026401f
C934 VTAIL.n258 VSUBS 0.026401f
C935 VTAIL.n259 VSUBS 0.014187f
C936 VTAIL.n260 VSUBS 0.015021f
C937 VTAIL.n261 VSUBS 0.033533f
C938 VTAIL.n262 VSUBS 0.033533f
C939 VTAIL.n263 VSUBS 0.015021f
C940 VTAIL.n264 VSUBS 0.014187f
C941 VTAIL.n265 VSUBS 0.026401f
C942 VTAIL.n266 VSUBS 0.026401f
C943 VTAIL.n267 VSUBS 0.014187f
C944 VTAIL.n268 VSUBS 0.015021f
C945 VTAIL.n269 VSUBS 0.033533f
C946 VTAIL.n270 VSUBS 0.033533f
C947 VTAIL.n271 VSUBS 0.015021f
C948 VTAIL.n272 VSUBS 0.014187f
C949 VTAIL.n273 VSUBS 0.026401f
C950 VTAIL.n274 VSUBS 0.026401f
C951 VTAIL.n275 VSUBS 0.014187f
C952 VTAIL.n276 VSUBS 0.015021f
C953 VTAIL.n277 VSUBS 0.033533f
C954 VTAIL.n278 VSUBS 0.033533f
C955 VTAIL.n279 VSUBS 0.015021f
C956 VTAIL.n280 VSUBS 0.014187f
C957 VTAIL.n281 VSUBS 0.026401f
C958 VTAIL.n282 VSUBS 0.026401f
C959 VTAIL.n283 VSUBS 0.014187f
C960 VTAIL.n284 VSUBS 0.015021f
C961 VTAIL.n285 VSUBS 0.033533f
C962 VTAIL.n286 VSUBS 0.033533f
C963 VTAIL.n287 VSUBS 0.015021f
C964 VTAIL.n288 VSUBS 0.014187f
C965 VTAIL.n289 VSUBS 0.026401f
C966 VTAIL.n290 VSUBS 0.026401f
C967 VTAIL.n291 VSUBS 0.014187f
C968 VTAIL.n292 VSUBS 0.015021f
C969 VTAIL.n293 VSUBS 0.033533f
C970 VTAIL.n294 VSUBS 0.08004f
C971 VTAIL.n295 VSUBS 0.015021f
C972 VTAIL.n296 VSUBS 0.014187f
C973 VTAIL.n297 VSUBS 0.057418f
C974 VTAIL.n298 VSUBS 0.040087f
C975 VTAIL.n299 VSUBS 1.48066f
C976 VTAIL.t10 VSUBS 0.280817f
C977 VTAIL.t8 VSUBS 0.280817f
C978 VTAIL.n300 VSUBS 2.06515f
C979 VTAIL.n301 VSUBS 0.75256f
C980 VTAIL.n302 VSUBS 0.028675f
C981 VTAIL.n303 VSUBS 0.026401f
C982 VTAIL.n304 VSUBS 0.014187f
C983 VTAIL.n305 VSUBS 0.033533f
C984 VTAIL.n306 VSUBS 0.015021f
C985 VTAIL.n307 VSUBS 0.026401f
C986 VTAIL.n308 VSUBS 0.014187f
C987 VTAIL.n309 VSUBS 0.033533f
C988 VTAIL.n310 VSUBS 0.015021f
C989 VTAIL.n311 VSUBS 0.026401f
C990 VTAIL.n312 VSUBS 0.014187f
C991 VTAIL.n313 VSUBS 0.033533f
C992 VTAIL.n314 VSUBS 0.014604f
C993 VTAIL.n315 VSUBS 0.026401f
C994 VTAIL.n316 VSUBS 0.014604f
C995 VTAIL.n317 VSUBS 0.014187f
C996 VTAIL.n318 VSUBS 0.033533f
C997 VTAIL.n319 VSUBS 0.033533f
C998 VTAIL.n320 VSUBS 0.015021f
C999 VTAIL.n321 VSUBS 0.026401f
C1000 VTAIL.n322 VSUBS 0.014187f
C1001 VTAIL.n323 VSUBS 0.033533f
C1002 VTAIL.n324 VSUBS 0.015021f
C1003 VTAIL.n325 VSUBS 1.46607f
C1004 VTAIL.n326 VSUBS 0.014187f
C1005 VTAIL.t12 VSUBS 0.072386f
C1006 VTAIL.n327 VSUBS 0.225351f
C1007 VTAIL.n328 VSUBS 0.025225f
C1008 VTAIL.n329 VSUBS 0.025149f
C1009 VTAIL.n330 VSUBS 0.033533f
C1010 VTAIL.n331 VSUBS 0.015021f
C1011 VTAIL.n332 VSUBS 0.014187f
C1012 VTAIL.n333 VSUBS 0.026401f
C1013 VTAIL.n334 VSUBS 0.026401f
C1014 VTAIL.n335 VSUBS 0.014187f
C1015 VTAIL.n336 VSUBS 0.015021f
C1016 VTAIL.n337 VSUBS 0.033533f
C1017 VTAIL.n338 VSUBS 0.033533f
C1018 VTAIL.n339 VSUBS 0.015021f
C1019 VTAIL.n340 VSUBS 0.014187f
C1020 VTAIL.n341 VSUBS 0.026401f
C1021 VTAIL.n342 VSUBS 0.026401f
C1022 VTAIL.n343 VSUBS 0.014187f
C1023 VTAIL.n344 VSUBS 0.015021f
C1024 VTAIL.n345 VSUBS 0.033533f
C1025 VTAIL.n346 VSUBS 0.033533f
C1026 VTAIL.n347 VSUBS 0.015021f
C1027 VTAIL.n348 VSUBS 0.014187f
C1028 VTAIL.n349 VSUBS 0.026401f
C1029 VTAIL.n350 VSUBS 0.026401f
C1030 VTAIL.n351 VSUBS 0.014187f
C1031 VTAIL.n352 VSUBS 0.015021f
C1032 VTAIL.n353 VSUBS 0.033533f
C1033 VTAIL.n354 VSUBS 0.033533f
C1034 VTAIL.n355 VSUBS 0.015021f
C1035 VTAIL.n356 VSUBS 0.014187f
C1036 VTAIL.n357 VSUBS 0.026401f
C1037 VTAIL.n358 VSUBS 0.026401f
C1038 VTAIL.n359 VSUBS 0.014187f
C1039 VTAIL.n360 VSUBS 0.015021f
C1040 VTAIL.n361 VSUBS 0.033533f
C1041 VTAIL.n362 VSUBS 0.033533f
C1042 VTAIL.n363 VSUBS 0.015021f
C1043 VTAIL.n364 VSUBS 0.014187f
C1044 VTAIL.n365 VSUBS 0.026401f
C1045 VTAIL.n366 VSUBS 0.026401f
C1046 VTAIL.n367 VSUBS 0.014187f
C1047 VTAIL.n368 VSUBS 0.015021f
C1048 VTAIL.n369 VSUBS 0.033533f
C1049 VTAIL.n370 VSUBS 0.08004f
C1050 VTAIL.n371 VSUBS 0.015021f
C1051 VTAIL.n372 VSUBS 0.014187f
C1052 VTAIL.n373 VSUBS 0.057418f
C1053 VTAIL.n374 VSUBS 0.040087f
C1054 VTAIL.n375 VSUBS 0.117687f
C1055 VTAIL.n376 VSUBS 0.028675f
C1056 VTAIL.n377 VSUBS 0.026401f
C1057 VTAIL.n378 VSUBS 0.014187f
C1058 VTAIL.n379 VSUBS 0.033533f
C1059 VTAIL.n380 VSUBS 0.015021f
C1060 VTAIL.n381 VSUBS 0.026401f
C1061 VTAIL.n382 VSUBS 0.014187f
C1062 VTAIL.n383 VSUBS 0.033533f
C1063 VTAIL.n384 VSUBS 0.015021f
C1064 VTAIL.n385 VSUBS 0.026401f
C1065 VTAIL.n386 VSUBS 0.014187f
C1066 VTAIL.n387 VSUBS 0.033533f
C1067 VTAIL.n388 VSUBS 0.014604f
C1068 VTAIL.n389 VSUBS 0.026401f
C1069 VTAIL.n390 VSUBS 0.014604f
C1070 VTAIL.n391 VSUBS 0.014187f
C1071 VTAIL.n392 VSUBS 0.033533f
C1072 VTAIL.n393 VSUBS 0.033533f
C1073 VTAIL.n394 VSUBS 0.015021f
C1074 VTAIL.n395 VSUBS 0.026401f
C1075 VTAIL.n396 VSUBS 0.014187f
C1076 VTAIL.n397 VSUBS 0.033533f
C1077 VTAIL.n398 VSUBS 0.015021f
C1078 VTAIL.n399 VSUBS 1.46607f
C1079 VTAIL.n400 VSUBS 0.014187f
C1080 VTAIL.t6 VSUBS 0.072386f
C1081 VTAIL.n401 VSUBS 0.225351f
C1082 VTAIL.n402 VSUBS 0.025225f
C1083 VTAIL.n403 VSUBS 0.025149f
C1084 VTAIL.n404 VSUBS 0.033533f
C1085 VTAIL.n405 VSUBS 0.015021f
C1086 VTAIL.n406 VSUBS 0.014187f
C1087 VTAIL.n407 VSUBS 0.026401f
C1088 VTAIL.n408 VSUBS 0.026401f
C1089 VTAIL.n409 VSUBS 0.014187f
C1090 VTAIL.n410 VSUBS 0.015021f
C1091 VTAIL.n411 VSUBS 0.033533f
C1092 VTAIL.n412 VSUBS 0.033533f
C1093 VTAIL.n413 VSUBS 0.015021f
C1094 VTAIL.n414 VSUBS 0.014187f
C1095 VTAIL.n415 VSUBS 0.026401f
C1096 VTAIL.n416 VSUBS 0.026401f
C1097 VTAIL.n417 VSUBS 0.014187f
C1098 VTAIL.n418 VSUBS 0.015021f
C1099 VTAIL.n419 VSUBS 0.033533f
C1100 VTAIL.n420 VSUBS 0.033533f
C1101 VTAIL.n421 VSUBS 0.015021f
C1102 VTAIL.n422 VSUBS 0.014187f
C1103 VTAIL.n423 VSUBS 0.026401f
C1104 VTAIL.n424 VSUBS 0.026401f
C1105 VTAIL.n425 VSUBS 0.014187f
C1106 VTAIL.n426 VSUBS 0.015021f
C1107 VTAIL.n427 VSUBS 0.033533f
C1108 VTAIL.n428 VSUBS 0.033533f
C1109 VTAIL.n429 VSUBS 0.015021f
C1110 VTAIL.n430 VSUBS 0.014187f
C1111 VTAIL.n431 VSUBS 0.026401f
C1112 VTAIL.n432 VSUBS 0.026401f
C1113 VTAIL.n433 VSUBS 0.014187f
C1114 VTAIL.n434 VSUBS 0.015021f
C1115 VTAIL.n435 VSUBS 0.033533f
C1116 VTAIL.n436 VSUBS 0.033533f
C1117 VTAIL.n437 VSUBS 0.015021f
C1118 VTAIL.n438 VSUBS 0.014187f
C1119 VTAIL.n439 VSUBS 0.026401f
C1120 VTAIL.n440 VSUBS 0.026401f
C1121 VTAIL.n441 VSUBS 0.014187f
C1122 VTAIL.n442 VSUBS 0.015021f
C1123 VTAIL.n443 VSUBS 0.033533f
C1124 VTAIL.n444 VSUBS 0.08004f
C1125 VTAIL.n445 VSUBS 0.015021f
C1126 VTAIL.n446 VSUBS 0.014187f
C1127 VTAIL.n447 VSUBS 0.057418f
C1128 VTAIL.n448 VSUBS 0.040087f
C1129 VTAIL.n449 VSUBS 0.117687f
C1130 VTAIL.t3 VSUBS 0.280817f
C1131 VTAIL.t1 VSUBS 0.280817f
C1132 VTAIL.n450 VSUBS 2.06515f
C1133 VTAIL.n451 VSUBS 0.75256f
C1134 VTAIL.n452 VSUBS 0.028675f
C1135 VTAIL.n453 VSUBS 0.026401f
C1136 VTAIL.n454 VSUBS 0.014187f
C1137 VTAIL.n455 VSUBS 0.033533f
C1138 VTAIL.n456 VSUBS 0.015021f
C1139 VTAIL.n457 VSUBS 0.026401f
C1140 VTAIL.n458 VSUBS 0.014187f
C1141 VTAIL.n459 VSUBS 0.033533f
C1142 VTAIL.n460 VSUBS 0.015021f
C1143 VTAIL.n461 VSUBS 0.026401f
C1144 VTAIL.n462 VSUBS 0.014187f
C1145 VTAIL.n463 VSUBS 0.033533f
C1146 VTAIL.n464 VSUBS 0.014604f
C1147 VTAIL.n465 VSUBS 0.026401f
C1148 VTAIL.n466 VSUBS 0.014604f
C1149 VTAIL.n467 VSUBS 0.014187f
C1150 VTAIL.n468 VSUBS 0.033533f
C1151 VTAIL.n469 VSUBS 0.033533f
C1152 VTAIL.n470 VSUBS 0.015021f
C1153 VTAIL.n471 VSUBS 0.026401f
C1154 VTAIL.n472 VSUBS 0.014187f
C1155 VTAIL.n473 VSUBS 0.033533f
C1156 VTAIL.n474 VSUBS 0.015021f
C1157 VTAIL.n475 VSUBS 1.46607f
C1158 VTAIL.n476 VSUBS 0.014187f
C1159 VTAIL.t0 VSUBS 0.072386f
C1160 VTAIL.n477 VSUBS 0.225351f
C1161 VTAIL.n478 VSUBS 0.025225f
C1162 VTAIL.n479 VSUBS 0.025149f
C1163 VTAIL.n480 VSUBS 0.033533f
C1164 VTAIL.n481 VSUBS 0.015021f
C1165 VTAIL.n482 VSUBS 0.014187f
C1166 VTAIL.n483 VSUBS 0.026401f
C1167 VTAIL.n484 VSUBS 0.026401f
C1168 VTAIL.n485 VSUBS 0.014187f
C1169 VTAIL.n486 VSUBS 0.015021f
C1170 VTAIL.n487 VSUBS 0.033533f
C1171 VTAIL.n488 VSUBS 0.033533f
C1172 VTAIL.n489 VSUBS 0.015021f
C1173 VTAIL.n490 VSUBS 0.014187f
C1174 VTAIL.n491 VSUBS 0.026401f
C1175 VTAIL.n492 VSUBS 0.026401f
C1176 VTAIL.n493 VSUBS 0.014187f
C1177 VTAIL.n494 VSUBS 0.015021f
C1178 VTAIL.n495 VSUBS 0.033533f
C1179 VTAIL.n496 VSUBS 0.033533f
C1180 VTAIL.n497 VSUBS 0.015021f
C1181 VTAIL.n498 VSUBS 0.014187f
C1182 VTAIL.n499 VSUBS 0.026401f
C1183 VTAIL.n500 VSUBS 0.026401f
C1184 VTAIL.n501 VSUBS 0.014187f
C1185 VTAIL.n502 VSUBS 0.015021f
C1186 VTAIL.n503 VSUBS 0.033533f
C1187 VTAIL.n504 VSUBS 0.033533f
C1188 VTAIL.n505 VSUBS 0.015021f
C1189 VTAIL.n506 VSUBS 0.014187f
C1190 VTAIL.n507 VSUBS 0.026401f
C1191 VTAIL.n508 VSUBS 0.026401f
C1192 VTAIL.n509 VSUBS 0.014187f
C1193 VTAIL.n510 VSUBS 0.015021f
C1194 VTAIL.n511 VSUBS 0.033533f
C1195 VTAIL.n512 VSUBS 0.033533f
C1196 VTAIL.n513 VSUBS 0.015021f
C1197 VTAIL.n514 VSUBS 0.014187f
C1198 VTAIL.n515 VSUBS 0.026401f
C1199 VTAIL.n516 VSUBS 0.026401f
C1200 VTAIL.n517 VSUBS 0.014187f
C1201 VTAIL.n518 VSUBS 0.015021f
C1202 VTAIL.n519 VSUBS 0.033533f
C1203 VTAIL.n520 VSUBS 0.08004f
C1204 VTAIL.n521 VSUBS 0.015021f
C1205 VTAIL.n522 VSUBS 0.014187f
C1206 VTAIL.n523 VSUBS 0.057418f
C1207 VTAIL.n524 VSUBS 0.040087f
C1208 VTAIL.n525 VSUBS 1.48066f
C1209 VTAIL.n526 VSUBS 0.028675f
C1210 VTAIL.n527 VSUBS 0.026401f
C1211 VTAIL.n528 VSUBS 0.014187f
C1212 VTAIL.n529 VSUBS 0.033533f
C1213 VTAIL.n530 VSUBS 0.015021f
C1214 VTAIL.n531 VSUBS 0.026401f
C1215 VTAIL.n532 VSUBS 0.014187f
C1216 VTAIL.n533 VSUBS 0.033533f
C1217 VTAIL.n534 VSUBS 0.015021f
C1218 VTAIL.n535 VSUBS 0.026401f
C1219 VTAIL.n536 VSUBS 0.014187f
C1220 VTAIL.n537 VSUBS 0.033533f
C1221 VTAIL.n538 VSUBS 0.014604f
C1222 VTAIL.n539 VSUBS 0.026401f
C1223 VTAIL.n540 VSUBS 0.015021f
C1224 VTAIL.n541 VSUBS 0.033533f
C1225 VTAIL.n542 VSUBS 0.015021f
C1226 VTAIL.n543 VSUBS 0.026401f
C1227 VTAIL.n544 VSUBS 0.014187f
C1228 VTAIL.n545 VSUBS 0.033533f
C1229 VTAIL.n546 VSUBS 0.015021f
C1230 VTAIL.n547 VSUBS 1.46607f
C1231 VTAIL.n548 VSUBS 0.014187f
C1232 VTAIL.t11 VSUBS 0.072386f
C1233 VTAIL.n549 VSUBS 0.225351f
C1234 VTAIL.n550 VSUBS 0.025225f
C1235 VTAIL.n551 VSUBS 0.025149f
C1236 VTAIL.n552 VSUBS 0.033533f
C1237 VTAIL.n553 VSUBS 0.015021f
C1238 VTAIL.n554 VSUBS 0.014187f
C1239 VTAIL.n555 VSUBS 0.026401f
C1240 VTAIL.n556 VSUBS 0.026401f
C1241 VTAIL.n557 VSUBS 0.014187f
C1242 VTAIL.n558 VSUBS 0.015021f
C1243 VTAIL.n559 VSUBS 0.033533f
C1244 VTAIL.n560 VSUBS 0.033533f
C1245 VTAIL.n561 VSUBS 0.015021f
C1246 VTAIL.n562 VSUBS 0.014187f
C1247 VTAIL.n563 VSUBS 0.026401f
C1248 VTAIL.n564 VSUBS 0.026401f
C1249 VTAIL.n565 VSUBS 0.014187f
C1250 VTAIL.n566 VSUBS 0.014187f
C1251 VTAIL.n567 VSUBS 0.015021f
C1252 VTAIL.n568 VSUBS 0.033533f
C1253 VTAIL.n569 VSUBS 0.033533f
C1254 VTAIL.n570 VSUBS 0.033533f
C1255 VTAIL.n571 VSUBS 0.014604f
C1256 VTAIL.n572 VSUBS 0.014187f
C1257 VTAIL.n573 VSUBS 0.026401f
C1258 VTAIL.n574 VSUBS 0.026401f
C1259 VTAIL.n575 VSUBS 0.014187f
C1260 VTAIL.n576 VSUBS 0.015021f
C1261 VTAIL.n577 VSUBS 0.033533f
C1262 VTAIL.n578 VSUBS 0.033533f
C1263 VTAIL.n579 VSUBS 0.015021f
C1264 VTAIL.n580 VSUBS 0.014187f
C1265 VTAIL.n581 VSUBS 0.026401f
C1266 VTAIL.n582 VSUBS 0.026401f
C1267 VTAIL.n583 VSUBS 0.014187f
C1268 VTAIL.n584 VSUBS 0.015021f
C1269 VTAIL.n585 VSUBS 0.033533f
C1270 VTAIL.n586 VSUBS 0.033533f
C1271 VTAIL.n587 VSUBS 0.015021f
C1272 VTAIL.n588 VSUBS 0.014187f
C1273 VTAIL.n589 VSUBS 0.026401f
C1274 VTAIL.n590 VSUBS 0.026401f
C1275 VTAIL.n591 VSUBS 0.014187f
C1276 VTAIL.n592 VSUBS 0.015021f
C1277 VTAIL.n593 VSUBS 0.033533f
C1278 VTAIL.n594 VSUBS 0.08004f
C1279 VTAIL.n595 VSUBS 0.015021f
C1280 VTAIL.n596 VSUBS 0.014187f
C1281 VTAIL.n597 VSUBS 0.057418f
C1282 VTAIL.n598 VSUBS 0.040087f
C1283 VTAIL.n599 VSUBS 1.47571f
C1284 VN.n0 VSUBS 0.06103f
C1285 VN.t2 VSUBS 1.05263f
C1286 VN.n1 VSUBS 0.424641f
C1287 VN.t3 VSUBS 1.06321f
C1288 VN.n2 VSUBS 0.408297f
C1289 VN.n3 VSUBS 0.19356f
C1290 VN.n4 VSUBS 0.013849f
C1291 VN.t1 VSUBS 1.05263f
C1292 VN.n5 VSUBS 0.424641f
C1293 VN.t0 VSUBS 1.05263f
C1294 VN.n6 VSUBS 0.418432f
C1295 VN.n7 VSUBS 0.047296f
C1296 VN.n8 VSUBS 0.06103f
C1297 VN.t7 VSUBS 1.05263f
C1298 VN.n9 VSUBS 0.424641f
C1299 VN.t5 VSUBS 1.06321f
C1300 VN.n10 VSUBS 0.408297f
C1301 VN.n11 VSUBS 0.19356f
C1302 VN.n12 VSUBS 0.013849f
C1303 VN.t6 VSUBS 1.05263f
C1304 VN.n13 VSUBS 0.424641f
C1305 VN.t4 VSUBS 1.05263f
C1306 VN.n14 VSUBS 0.418432f
C1307 VN.n15 VSUBS 2.55554f
.ends

