* NGSPICE file created from diff_pair_sample_1078.ext - technology: sky130A

.subckt diff_pair_sample_1078 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t5 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=0.56595 pd=3.76 as=1.3377 ps=7.64 w=3.43 l=2.33
X1 VTAIL.t3 VP.t0 VDD1.t3 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0.56595 ps=3.76 w=3.43 l=2.33
X2 B.t11 B.t9 B.t10 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0 ps=0 w=3.43 l=2.33
X3 B.t8 B.t6 B.t7 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0 ps=0 w=3.43 l=2.33
X4 VDD2.t2 VN.t1 VTAIL.t7 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=0.56595 pd=3.76 as=1.3377 ps=7.64 w=3.43 l=2.33
X5 VTAIL.t6 VN.t2 VDD2.t1 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0.56595 ps=3.76 w=3.43 l=2.33
X6 B.t5 B.t3 B.t4 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0 ps=0 w=3.43 l=2.33
X7 B.t2 B.t0 B.t1 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0 ps=0 w=3.43 l=2.33
X8 VTAIL.t4 VN.t3 VDD2.t0 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0.56595 ps=3.76 w=3.43 l=2.33
X9 VDD1.t2 VP.t1 VTAIL.t2 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=0.56595 pd=3.76 as=1.3377 ps=7.64 w=3.43 l=2.33
X10 VTAIL.t1 VP.t2 VDD1.t1 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=1.3377 pd=7.64 as=0.56595 ps=3.76 w=3.43 l=2.33
X11 VDD1.t0 VP.t3 VTAIL.t0 w_n2566_n1654# sky130_fd_pr__pfet_01v8 ad=0.56595 pd=3.76 as=1.3377 ps=7.64 w=3.43 l=2.33
R0 VN.n0 VN.t3 72.0047
R1 VN.n1 VN.t1 72.0047
R2 VN.n0 VN.t0 71.3464
R3 VN.n1 VN.t2 71.3464
R4 VN VN.n1 44.7715
R5 VN VN.n0 5.4874
R6 VTAIL.n5 VTAIL.t1 111.737
R7 VTAIL.n4 VTAIL.t7 111.737
R8 VTAIL.n3 VTAIL.t6 111.737
R9 VTAIL.n7 VTAIL.t5 111.737
R10 VTAIL.n0 VTAIL.t4 111.737
R11 VTAIL.n1 VTAIL.t2 111.737
R12 VTAIL.n2 VTAIL.t3 111.737
R13 VTAIL.n6 VTAIL.t0 111.737
R14 VTAIL.n7 VTAIL.n6 17.6169
R15 VTAIL.n3 VTAIL.n2 17.6169
R16 VTAIL.n4 VTAIL.n3 2.2936
R17 VTAIL.n6 VTAIL.n5 2.2936
R18 VTAIL.n2 VTAIL.n1 2.2936
R19 VTAIL VTAIL.n0 1.20524
R20 VTAIL VTAIL.n7 1.08886
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 152.489
R24 VDD2.n2 VDD2.n1 118.939
R25 VDD2.n1 VDD2.t1 9.47718
R26 VDD2.n1 VDD2.t2 9.47718
R27 VDD2.n0 VDD2.t0 9.47718
R28 VDD2.n0 VDD2.t3 9.47718
R29 VDD2 VDD2.n2 0.0586897
R30 VP.n12 VP.n0 161.3
R31 VP.n11 VP.n10 161.3
R32 VP.n9 VP.n1 161.3
R33 VP.n8 VP.n7 161.3
R34 VP.n6 VP.n2 161.3
R35 VP.n5 VP.n4 94.6082
R36 VP.n14 VP.n13 94.6082
R37 VP.n3 VP.t2 72.0047
R38 VP.n3 VP.t3 71.3464
R39 VP.n4 VP.n3 44.4926
R40 VP.n7 VP.n1 40.4934
R41 VP.n11 VP.n1 40.4934
R42 VP.n5 VP.t0 35.4782
R43 VP.n13 VP.t1 35.4782
R44 VP.n7 VP.n6 24.4675
R45 VP.n12 VP.n11 24.4675
R46 VP.n6 VP.n5 16.1487
R47 VP.n13 VP.n12 16.1487
R48 VP.n4 VP.n2 0.278367
R49 VP.n14 VP.n0 0.278367
R50 VP.n8 VP.n2 0.189894
R51 VP.n9 VP.n8 0.189894
R52 VP.n10 VP.n9 0.189894
R53 VP.n10 VP.n0 0.189894
R54 VP VP.n14 0.153454
R55 VDD1 VDD1.n1 153.014
R56 VDD1 VDD1.n0 118.996
R57 VDD1.n0 VDD1.t1 9.47718
R58 VDD1.n0 VDD1.t0 9.47718
R59 VDD1.n1 VDD1.t3 9.47718
R60 VDD1.n1 VDD1.t2 9.47718
R61 B.n225 B.n224 585
R62 B.n223 B.n76 585
R63 B.n222 B.n221 585
R64 B.n220 B.n77 585
R65 B.n219 B.n218 585
R66 B.n217 B.n78 585
R67 B.n216 B.n215 585
R68 B.n214 B.n79 585
R69 B.n213 B.n212 585
R70 B.n211 B.n80 585
R71 B.n210 B.n209 585
R72 B.n208 B.n81 585
R73 B.n207 B.n206 585
R74 B.n205 B.n82 585
R75 B.n204 B.n203 585
R76 B.n202 B.n83 585
R77 B.n201 B.n200 585
R78 B.n196 B.n84 585
R79 B.n195 B.n194 585
R80 B.n193 B.n85 585
R81 B.n192 B.n191 585
R82 B.n190 B.n86 585
R83 B.n189 B.n188 585
R84 B.n187 B.n87 585
R85 B.n186 B.n185 585
R86 B.n184 B.n88 585
R87 B.n182 B.n181 585
R88 B.n180 B.n91 585
R89 B.n179 B.n178 585
R90 B.n177 B.n92 585
R91 B.n176 B.n175 585
R92 B.n174 B.n93 585
R93 B.n173 B.n172 585
R94 B.n171 B.n94 585
R95 B.n170 B.n169 585
R96 B.n168 B.n95 585
R97 B.n167 B.n166 585
R98 B.n165 B.n96 585
R99 B.n164 B.n163 585
R100 B.n162 B.n97 585
R101 B.n161 B.n160 585
R102 B.n159 B.n98 585
R103 B.n226 B.n75 585
R104 B.n228 B.n227 585
R105 B.n229 B.n74 585
R106 B.n231 B.n230 585
R107 B.n232 B.n73 585
R108 B.n234 B.n233 585
R109 B.n235 B.n72 585
R110 B.n237 B.n236 585
R111 B.n238 B.n71 585
R112 B.n240 B.n239 585
R113 B.n241 B.n70 585
R114 B.n243 B.n242 585
R115 B.n244 B.n69 585
R116 B.n246 B.n245 585
R117 B.n247 B.n68 585
R118 B.n249 B.n248 585
R119 B.n250 B.n67 585
R120 B.n252 B.n251 585
R121 B.n253 B.n66 585
R122 B.n255 B.n254 585
R123 B.n256 B.n65 585
R124 B.n258 B.n257 585
R125 B.n259 B.n64 585
R126 B.n261 B.n260 585
R127 B.n262 B.n63 585
R128 B.n264 B.n263 585
R129 B.n265 B.n62 585
R130 B.n267 B.n266 585
R131 B.n268 B.n61 585
R132 B.n270 B.n269 585
R133 B.n271 B.n60 585
R134 B.n273 B.n272 585
R135 B.n274 B.n59 585
R136 B.n276 B.n275 585
R137 B.n277 B.n58 585
R138 B.n279 B.n278 585
R139 B.n280 B.n57 585
R140 B.n282 B.n281 585
R141 B.n283 B.n56 585
R142 B.n285 B.n284 585
R143 B.n286 B.n55 585
R144 B.n288 B.n287 585
R145 B.n289 B.n54 585
R146 B.n291 B.n290 585
R147 B.n292 B.n53 585
R148 B.n294 B.n293 585
R149 B.n295 B.n52 585
R150 B.n297 B.n296 585
R151 B.n298 B.n51 585
R152 B.n300 B.n299 585
R153 B.n301 B.n50 585
R154 B.n303 B.n302 585
R155 B.n304 B.n49 585
R156 B.n306 B.n305 585
R157 B.n307 B.n48 585
R158 B.n309 B.n308 585
R159 B.n310 B.n47 585
R160 B.n312 B.n311 585
R161 B.n313 B.n46 585
R162 B.n315 B.n314 585
R163 B.n316 B.n45 585
R164 B.n318 B.n317 585
R165 B.n319 B.n44 585
R166 B.n321 B.n320 585
R167 B.n385 B.n384 585
R168 B.n383 B.n18 585
R169 B.n382 B.n381 585
R170 B.n380 B.n19 585
R171 B.n379 B.n378 585
R172 B.n377 B.n20 585
R173 B.n376 B.n375 585
R174 B.n374 B.n21 585
R175 B.n373 B.n372 585
R176 B.n371 B.n22 585
R177 B.n370 B.n369 585
R178 B.n368 B.n23 585
R179 B.n367 B.n366 585
R180 B.n365 B.n24 585
R181 B.n364 B.n363 585
R182 B.n362 B.n25 585
R183 B.n360 B.n359 585
R184 B.n358 B.n28 585
R185 B.n357 B.n356 585
R186 B.n355 B.n29 585
R187 B.n354 B.n353 585
R188 B.n352 B.n30 585
R189 B.n351 B.n350 585
R190 B.n349 B.n31 585
R191 B.n348 B.n347 585
R192 B.n346 B.n32 585
R193 B.n345 B.n344 585
R194 B.n343 B.n33 585
R195 B.n342 B.n341 585
R196 B.n340 B.n37 585
R197 B.n339 B.n338 585
R198 B.n337 B.n38 585
R199 B.n336 B.n335 585
R200 B.n334 B.n39 585
R201 B.n333 B.n332 585
R202 B.n331 B.n40 585
R203 B.n330 B.n329 585
R204 B.n328 B.n41 585
R205 B.n327 B.n326 585
R206 B.n325 B.n42 585
R207 B.n324 B.n323 585
R208 B.n322 B.n43 585
R209 B.n386 B.n17 585
R210 B.n388 B.n387 585
R211 B.n389 B.n16 585
R212 B.n391 B.n390 585
R213 B.n392 B.n15 585
R214 B.n394 B.n393 585
R215 B.n395 B.n14 585
R216 B.n397 B.n396 585
R217 B.n398 B.n13 585
R218 B.n400 B.n399 585
R219 B.n401 B.n12 585
R220 B.n403 B.n402 585
R221 B.n404 B.n11 585
R222 B.n406 B.n405 585
R223 B.n407 B.n10 585
R224 B.n409 B.n408 585
R225 B.n410 B.n9 585
R226 B.n412 B.n411 585
R227 B.n413 B.n8 585
R228 B.n415 B.n414 585
R229 B.n416 B.n7 585
R230 B.n418 B.n417 585
R231 B.n419 B.n6 585
R232 B.n421 B.n420 585
R233 B.n422 B.n5 585
R234 B.n424 B.n423 585
R235 B.n425 B.n4 585
R236 B.n427 B.n426 585
R237 B.n428 B.n3 585
R238 B.n430 B.n429 585
R239 B.n431 B.n0 585
R240 B.n2 B.n1 585
R241 B.n114 B.n113 585
R242 B.n116 B.n115 585
R243 B.n117 B.n112 585
R244 B.n119 B.n118 585
R245 B.n120 B.n111 585
R246 B.n122 B.n121 585
R247 B.n123 B.n110 585
R248 B.n125 B.n124 585
R249 B.n126 B.n109 585
R250 B.n128 B.n127 585
R251 B.n129 B.n108 585
R252 B.n131 B.n130 585
R253 B.n132 B.n107 585
R254 B.n134 B.n133 585
R255 B.n135 B.n106 585
R256 B.n137 B.n136 585
R257 B.n138 B.n105 585
R258 B.n140 B.n139 585
R259 B.n141 B.n104 585
R260 B.n143 B.n142 585
R261 B.n144 B.n103 585
R262 B.n146 B.n145 585
R263 B.n147 B.n102 585
R264 B.n149 B.n148 585
R265 B.n150 B.n101 585
R266 B.n152 B.n151 585
R267 B.n153 B.n100 585
R268 B.n155 B.n154 585
R269 B.n156 B.n99 585
R270 B.n158 B.n157 585
R271 B.n157 B.n98 545.355
R272 B.n226 B.n225 545.355
R273 B.n322 B.n321 545.355
R274 B.n384 B.n17 545.355
R275 B.n433 B.n432 256.663
R276 B.n89 B.t0 243.077
R277 B.n197 B.t9 243.077
R278 B.n34 B.t6 243.077
R279 B.n26 B.t3 243.077
R280 B.n432 B.n431 235.042
R281 B.n432 B.n2 235.042
R282 B.n197 B.t10 178.714
R283 B.n34 B.t8 178.714
R284 B.n89 B.t1 178.713
R285 B.n26 B.t5 178.713
R286 B.n161 B.n98 163.367
R287 B.n162 B.n161 163.367
R288 B.n163 B.n162 163.367
R289 B.n163 B.n96 163.367
R290 B.n167 B.n96 163.367
R291 B.n168 B.n167 163.367
R292 B.n169 B.n168 163.367
R293 B.n169 B.n94 163.367
R294 B.n173 B.n94 163.367
R295 B.n174 B.n173 163.367
R296 B.n175 B.n174 163.367
R297 B.n175 B.n92 163.367
R298 B.n179 B.n92 163.367
R299 B.n180 B.n179 163.367
R300 B.n181 B.n180 163.367
R301 B.n181 B.n88 163.367
R302 B.n186 B.n88 163.367
R303 B.n187 B.n186 163.367
R304 B.n188 B.n187 163.367
R305 B.n188 B.n86 163.367
R306 B.n192 B.n86 163.367
R307 B.n193 B.n192 163.367
R308 B.n194 B.n193 163.367
R309 B.n194 B.n84 163.367
R310 B.n201 B.n84 163.367
R311 B.n202 B.n201 163.367
R312 B.n203 B.n202 163.367
R313 B.n203 B.n82 163.367
R314 B.n207 B.n82 163.367
R315 B.n208 B.n207 163.367
R316 B.n209 B.n208 163.367
R317 B.n209 B.n80 163.367
R318 B.n213 B.n80 163.367
R319 B.n214 B.n213 163.367
R320 B.n215 B.n214 163.367
R321 B.n215 B.n78 163.367
R322 B.n219 B.n78 163.367
R323 B.n220 B.n219 163.367
R324 B.n221 B.n220 163.367
R325 B.n221 B.n76 163.367
R326 B.n225 B.n76 163.367
R327 B.n321 B.n44 163.367
R328 B.n317 B.n44 163.367
R329 B.n317 B.n316 163.367
R330 B.n316 B.n315 163.367
R331 B.n315 B.n46 163.367
R332 B.n311 B.n46 163.367
R333 B.n311 B.n310 163.367
R334 B.n310 B.n309 163.367
R335 B.n309 B.n48 163.367
R336 B.n305 B.n48 163.367
R337 B.n305 B.n304 163.367
R338 B.n304 B.n303 163.367
R339 B.n303 B.n50 163.367
R340 B.n299 B.n50 163.367
R341 B.n299 B.n298 163.367
R342 B.n298 B.n297 163.367
R343 B.n297 B.n52 163.367
R344 B.n293 B.n52 163.367
R345 B.n293 B.n292 163.367
R346 B.n292 B.n291 163.367
R347 B.n291 B.n54 163.367
R348 B.n287 B.n54 163.367
R349 B.n287 B.n286 163.367
R350 B.n286 B.n285 163.367
R351 B.n285 B.n56 163.367
R352 B.n281 B.n56 163.367
R353 B.n281 B.n280 163.367
R354 B.n280 B.n279 163.367
R355 B.n279 B.n58 163.367
R356 B.n275 B.n58 163.367
R357 B.n275 B.n274 163.367
R358 B.n274 B.n273 163.367
R359 B.n273 B.n60 163.367
R360 B.n269 B.n60 163.367
R361 B.n269 B.n268 163.367
R362 B.n268 B.n267 163.367
R363 B.n267 B.n62 163.367
R364 B.n263 B.n62 163.367
R365 B.n263 B.n262 163.367
R366 B.n262 B.n261 163.367
R367 B.n261 B.n64 163.367
R368 B.n257 B.n64 163.367
R369 B.n257 B.n256 163.367
R370 B.n256 B.n255 163.367
R371 B.n255 B.n66 163.367
R372 B.n251 B.n66 163.367
R373 B.n251 B.n250 163.367
R374 B.n250 B.n249 163.367
R375 B.n249 B.n68 163.367
R376 B.n245 B.n68 163.367
R377 B.n245 B.n244 163.367
R378 B.n244 B.n243 163.367
R379 B.n243 B.n70 163.367
R380 B.n239 B.n70 163.367
R381 B.n239 B.n238 163.367
R382 B.n238 B.n237 163.367
R383 B.n237 B.n72 163.367
R384 B.n233 B.n72 163.367
R385 B.n233 B.n232 163.367
R386 B.n232 B.n231 163.367
R387 B.n231 B.n74 163.367
R388 B.n227 B.n74 163.367
R389 B.n227 B.n226 163.367
R390 B.n384 B.n383 163.367
R391 B.n383 B.n382 163.367
R392 B.n382 B.n19 163.367
R393 B.n378 B.n19 163.367
R394 B.n378 B.n377 163.367
R395 B.n377 B.n376 163.367
R396 B.n376 B.n21 163.367
R397 B.n372 B.n21 163.367
R398 B.n372 B.n371 163.367
R399 B.n371 B.n370 163.367
R400 B.n370 B.n23 163.367
R401 B.n366 B.n23 163.367
R402 B.n366 B.n365 163.367
R403 B.n365 B.n364 163.367
R404 B.n364 B.n25 163.367
R405 B.n359 B.n25 163.367
R406 B.n359 B.n358 163.367
R407 B.n358 B.n357 163.367
R408 B.n357 B.n29 163.367
R409 B.n353 B.n29 163.367
R410 B.n353 B.n352 163.367
R411 B.n352 B.n351 163.367
R412 B.n351 B.n31 163.367
R413 B.n347 B.n31 163.367
R414 B.n347 B.n346 163.367
R415 B.n346 B.n345 163.367
R416 B.n345 B.n33 163.367
R417 B.n341 B.n33 163.367
R418 B.n341 B.n340 163.367
R419 B.n340 B.n339 163.367
R420 B.n339 B.n38 163.367
R421 B.n335 B.n38 163.367
R422 B.n335 B.n334 163.367
R423 B.n334 B.n333 163.367
R424 B.n333 B.n40 163.367
R425 B.n329 B.n40 163.367
R426 B.n329 B.n328 163.367
R427 B.n328 B.n327 163.367
R428 B.n327 B.n42 163.367
R429 B.n323 B.n42 163.367
R430 B.n323 B.n322 163.367
R431 B.n388 B.n17 163.367
R432 B.n389 B.n388 163.367
R433 B.n390 B.n389 163.367
R434 B.n390 B.n15 163.367
R435 B.n394 B.n15 163.367
R436 B.n395 B.n394 163.367
R437 B.n396 B.n395 163.367
R438 B.n396 B.n13 163.367
R439 B.n400 B.n13 163.367
R440 B.n401 B.n400 163.367
R441 B.n402 B.n401 163.367
R442 B.n402 B.n11 163.367
R443 B.n406 B.n11 163.367
R444 B.n407 B.n406 163.367
R445 B.n408 B.n407 163.367
R446 B.n408 B.n9 163.367
R447 B.n412 B.n9 163.367
R448 B.n413 B.n412 163.367
R449 B.n414 B.n413 163.367
R450 B.n414 B.n7 163.367
R451 B.n418 B.n7 163.367
R452 B.n419 B.n418 163.367
R453 B.n420 B.n419 163.367
R454 B.n420 B.n5 163.367
R455 B.n424 B.n5 163.367
R456 B.n425 B.n424 163.367
R457 B.n426 B.n425 163.367
R458 B.n426 B.n3 163.367
R459 B.n430 B.n3 163.367
R460 B.n431 B.n430 163.367
R461 B.n114 B.n2 163.367
R462 B.n115 B.n114 163.367
R463 B.n115 B.n112 163.367
R464 B.n119 B.n112 163.367
R465 B.n120 B.n119 163.367
R466 B.n121 B.n120 163.367
R467 B.n121 B.n110 163.367
R468 B.n125 B.n110 163.367
R469 B.n126 B.n125 163.367
R470 B.n127 B.n126 163.367
R471 B.n127 B.n108 163.367
R472 B.n131 B.n108 163.367
R473 B.n132 B.n131 163.367
R474 B.n133 B.n132 163.367
R475 B.n133 B.n106 163.367
R476 B.n137 B.n106 163.367
R477 B.n138 B.n137 163.367
R478 B.n139 B.n138 163.367
R479 B.n139 B.n104 163.367
R480 B.n143 B.n104 163.367
R481 B.n144 B.n143 163.367
R482 B.n145 B.n144 163.367
R483 B.n145 B.n102 163.367
R484 B.n149 B.n102 163.367
R485 B.n150 B.n149 163.367
R486 B.n151 B.n150 163.367
R487 B.n151 B.n100 163.367
R488 B.n155 B.n100 163.367
R489 B.n156 B.n155 163.367
R490 B.n157 B.n156 163.367
R491 B.n198 B.t11 127.127
R492 B.n35 B.t7 127.127
R493 B.n90 B.t2 127.124
R494 B.n27 B.t4 127.124
R495 B.n183 B.n90 59.5399
R496 B.n199 B.n198 59.5399
R497 B.n36 B.n35 59.5399
R498 B.n361 B.n27 59.5399
R499 B.n90 B.n89 51.5884
R500 B.n198 B.n197 51.5884
R501 B.n35 B.n34 51.5884
R502 B.n27 B.n26 51.5884
R503 B.n386 B.n385 35.4346
R504 B.n320 B.n43 35.4346
R505 B.n159 B.n158 35.4346
R506 B.n224 B.n75 35.4346
R507 B B.n433 18.0485
R508 B.n387 B.n386 10.6151
R509 B.n387 B.n16 10.6151
R510 B.n391 B.n16 10.6151
R511 B.n392 B.n391 10.6151
R512 B.n393 B.n392 10.6151
R513 B.n393 B.n14 10.6151
R514 B.n397 B.n14 10.6151
R515 B.n398 B.n397 10.6151
R516 B.n399 B.n398 10.6151
R517 B.n399 B.n12 10.6151
R518 B.n403 B.n12 10.6151
R519 B.n404 B.n403 10.6151
R520 B.n405 B.n404 10.6151
R521 B.n405 B.n10 10.6151
R522 B.n409 B.n10 10.6151
R523 B.n410 B.n409 10.6151
R524 B.n411 B.n410 10.6151
R525 B.n411 B.n8 10.6151
R526 B.n415 B.n8 10.6151
R527 B.n416 B.n415 10.6151
R528 B.n417 B.n416 10.6151
R529 B.n417 B.n6 10.6151
R530 B.n421 B.n6 10.6151
R531 B.n422 B.n421 10.6151
R532 B.n423 B.n422 10.6151
R533 B.n423 B.n4 10.6151
R534 B.n427 B.n4 10.6151
R535 B.n428 B.n427 10.6151
R536 B.n429 B.n428 10.6151
R537 B.n429 B.n0 10.6151
R538 B.n385 B.n18 10.6151
R539 B.n381 B.n18 10.6151
R540 B.n381 B.n380 10.6151
R541 B.n380 B.n379 10.6151
R542 B.n379 B.n20 10.6151
R543 B.n375 B.n20 10.6151
R544 B.n375 B.n374 10.6151
R545 B.n374 B.n373 10.6151
R546 B.n373 B.n22 10.6151
R547 B.n369 B.n22 10.6151
R548 B.n369 B.n368 10.6151
R549 B.n368 B.n367 10.6151
R550 B.n367 B.n24 10.6151
R551 B.n363 B.n24 10.6151
R552 B.n363 B.n362 10.6151
R553 B.n360 B.n28 10.6151
R554 B.n356 B.n28 10.6151
R555 B.n356 B.n355 10.6151
R556 B.n355 B.n354 10.6151
R557 B.n354 B.n30 10.6151
R558 B.n350 B.n30 10.6151
R559 B.n350 B.n349 10.6151
R560 B.n349 B.n348 10.6151
R561 B.n348 B.n32 10.6151
R562 B.n344 B.n343 10.6151
R563 B.n343 B.n342 10.6151
R564 B.n342 B.n37 10.6151
R565 B.n338 B.n37 10.6151
R566 B.n338 B.n337 10.6151
R567 B.n337 B.n336 10.6151
R568 B.n336 B.n39 10.6151
R569 B.n332 B.n39 10.6151
R570 B.n332 B.n331 10.6151
R571 B.n331 B.n330 10.6151
R572 B.n330 B.n41 10.6151
R573 B.n326 B.n41 10.6151
R574 B.n326 B.n325 10.6151
R575 B.n325 B.n324 10.6151
R576 B.n324 B.n43 10.6151
R577 B.n320 B.n319 10.6151
R578 B.n319 B.n318 10.6151
R579 B.n318 B.n45 10.6151
R580 B.n314 B.n45 10.6151
R581 B.n314 B.n313 10.6151
R582 B.n313 B.n312 10.6151
R583 B.n312 B.n47 10.6151
R584 B.n308 B.n47 10.6151
R585 B.n308 B.n307 10.6151
R586 B.n307 B.n306 10.6151
R587 B.n306 B.n49 10.6151
R588 B.n302 B.n49 10.6151
R589 B.n302 B.n301 10.6151
R590 B.n301 B.n300 10.6151
R591 B.n300 B.n51 10.6151
R592 B.n296 B.n51 10.6151
R593 B.n296 B.n295 10.6151
R594 B.n295 B.n294 10.6151
R595 B.n294 B.n53 10.6151
R596 B.n290 B.n53 10.6151
R597 B.n290 B.n289 10.6151
R598 B.n289 B.n288 10.6151
R599 B.n288 B.n55 10.6151
R600 B.n284 B.n55 10.6151
R601 B.n284 B.n283 10.6151
R602 B.n283 B.n282 10.6151
R603 B.n282 B.n57 10.6151
R604 B.n278 B.n57 10.6151
R605 B.n278 B.n277 10.6151
R606 B.n277 B.n276 10.6151
R607 B.n276 B.n59 10.6151
R608 B.n272 B.n59 10.6151
R609 B.n272 B.n271 10.6151
R610 B.n271 B.n270 10.6151
R611 B.n270 B.n61 10.6151
R612 B.n266 B.n61 10.6151
R613 B.n266 B.n265 10.6151
R614 B.n265 B.n264 10.6151
R615 B.n264 B.n63 10.6151
R616 B.n260 B.n63 10.6151
R617 B.n260 B.n259 10.6151
R618 B.n259 B.n258 10.6151
R619 B.n258 B.n65 10.6151
R620 B.n254 B.n65 10.6151
R621 B.n254 B.n253 10.6151
R622 B.n253 B.n252 10.6151
R623 B.n252 B.n67 10.6151
R624 B.n248 B.n67 10.6151
R625 B.n248 B.n247 10.6151
R626 B.n247 B.n246 10.6151
R627 B.n246 B.n69 10.6151
R628 B.n242 B.n69 10.6151
R629 B.n242 B.n241 10.6151
R630 B.n241 B.n240 10.6151
R631 B.n240 B.n71 10.6151
R632 B.n236 B.n71 10.6151
R633 B.n236 B.n235 10.6151
R634 B.n235 B.n234 10.6151
R635 B.n234 B.n73 10.6151
R636 B.n230 B.n73 10.6151
R637 B.n230 B.n229 10.6151
R638 B.n229 B.n228 10.6151
R639 B.n228 B.n75 10.6151
R640 B.n113 B.n1 10.6151
R641 B.n116 B.n113 10.6151
R642 B.n117 B.n116 10.6151
R643 B.n118 B.n117 10.6151
R644 B.n118 B.n111 10.6151
R645 B.n122 B.n111 10.6151
R646 B.n123 B.n122 10.6151
R647 B.n124 B.n123 10.6151
R648 B.n124 B.n109 10.6151
R649 B.n128 B.n109 10.6151
R650 B.n129 B.n128 10.6151
R651 B.n130 B.n129 10.6151
R652 B.n130 B.n107 10.6151
R653 B.n134 B.n107 10.6151
R654 B.n135 B.n134 10.6151
R655 B.n136 B.n135 10.6151
R656 B.n136 B.n105 10.6151
R657 B.n140 B.n105 10.6151
R658 B.n141 B.n140 10.6151
R659 B.n142 B.n141 10.6151
R660 B.n142 B.n103 10.6151
R661 B.n146 B.n103 10.6151
R662 B.n147 B.n146 10.6151
R663 B.n148 B.n147 10.6151
R664 B.n148 B.n101 10.6151
R665 B.n152 B.n101 10.6151
R666 B.n153 B.n152 10.6151
R667 B.n154 B.n153 10.6151
R668 B.n154 B.n99 10.6151
R669 B.n158 B.n99 10.6151
R670 B.n160 B.n159 10.6151
R671 B.n160 B.n97 10.6151
R672 B.n164 B.n97 10.6151
R673 B.n165 B.n164 10.6151
R674 B.n166 B.n165 10.6151
R675 B.n166 B.n95 10.6151
R676 B.n170 B.n95 10.6151
R677 B.n171 B.n170 10.6151
R678 B.n172 B.n171 10.6151
R679 B.n172 B.n93 10.6151
R680 B.n176 B.n93 10.6151
R681 B.n177 B.n176 10.6151
R682 B.n178 B.n177 10.6151
R683 B.n178 B.n91 10.6151
R684 B.n182 B.n91 10.6151
R685 B.n185 B.n184 10.6151
R686 B.n185 B.n87 10.6151
R687 B.n189 B.n87 10.6151
R688 B.n190 B.n189 10.6151
R689 B.n191 B.n190 10.6151
R690 B.n191 B.n85 10.6151
R691 B.n195 B.n85 10.6151
R692 B.n196 B.n195 10.6151
R693 B.n200 B.n196 10.6151
R694 B.n204 B.n83 10.6151
R695 B.n205 B.n204 10.6151
R696 B.n206 B.n205 10.6151
R697 B.n206 B.n81 10.6151
R698 B.n210 B.n81 10.6151
R699 B.n211 B.n210 10.6151
R700 B.n212 B.n211 10.6151
R701 B.n212 B.n79 10.6151
R702 B.n216 B.n79 10.6151
R703 B.n217 B.n216 10.6151
R704 B.n218 B.n217 10.6151
R705 B.n218 B.n77 10.6151
R706 B.n222 B.n77 10.6151
R707 B.n223 B.n222 10.6151
R708 B.n224 B.n223 10.6151
R709 B.n362 B.n361 9.36635
R710 B.n344 B.n36 9.36635
R711 B.n183 B.n182 9.36635
R712 B.n199 B.n83 9.36635
R713 B.n433 B.n0 8.11757
R714 B.n433 B.n1 8.11757
R715 B.n361 B.n360 1.24928
R716 B.n36 B.n32 1.24928
R717 B.n184 B.n183 1.24928
R718 B.n200 B.n199 1.24928
C0 w_n2566_n1654# VP 4.4549f
C1 w_n2566_n1654# VN 4.12738f
C2 w_n2566_n1654# VDD1 1.1663f
C3 w_n2566_n1654# VTAIL 2.00208f
C4 w_n2566_n1654# B 6.52836f
C5 VP VDD2 0.382075f
C6 VN VDD2 1.56209f
C7 VDD2 VDD1 0.964595f
C8 VN VP 4.41419f
C9 VDD2 VTAIL 3.30079f
C10 VDD2 B 1.03201f
C11 VP VDD1 1.78974f
C12 VN VDD1 0.153197f
C13 VP VTAIL 1.95864f
C14 VP B 1.49722f
C15 VN VTAIL 1.94453f
C16 VN B 0.952524f
C17 VTAIL VDD1 3.24839f
C18 B VDD1 0.984141f
C19 B VTAIL 2.01039f
C20 w_n2566_n1654# VDD2 1.21595f
C21 VDD2 VSUBS 0.62093f
C22 VDD1 VSUBS 3.100759f
C23 VTAIL VSUBS 0.518523f
C24 VN VSUBS 4.51499f
C25 VP VSUBS 1.665149f
C26 B VSUBS 3.14204f
C27 w_n2566_n1654# VSUBS 53.6089f
C28 B.n0 VSUBS 0.008625f
C29 B.n1 VSUBS 0.008625f
C30 B.n2 VSUBS 0.012757f
C31 B.n3 VSUBS 0.009776f
C32 B.n4 VSUBS 0.009776f
C33 B.n5 VSUBS 0.009776f
C34 B.n6 VSUBS 0.009776f
C35 B.n7 VSUBS 0.009776f
C36 B.n8 VSUBS 0.009776f
C37 B.n9 VSUBS 0.009776f
C38 B.n10 VSUBS 0.009776f
C39 B.n11 VSUBS 0.009776f
C40 B.n12 VSUBS 0.009776f
C41 B.n13 VSUBS 0.009776f
C42 B.n14 VSUBS 0.009776f
C43 B.n15 VSUBS 0.009776f
C44 B.n16 VSUBS 0.009776f
C45 B.n17 VSUBS 0.023749f
C46 B.n18 VSUBS 0.009776f
C47 B.n19 VSUBS 0.009776f
C48 B.n20 VSUBS 0.009776f
C49 B.n21 VSUBS 0.009776f
C50 B.n22 VSUBS 0.009776f
C51 B.n23 VSUBS 0.009776f
C52 B.n24 VSUBS 0.009776f
C53 B.n25 VSUBS 0.009776f
C54 B.t4 VSUBS 0.120499f
C55 B.t5 VSUBS 0.142922f
C56 B.t3 VSUBS 0.538169f
C57 B.n26 VSUBS 0.115938f
C58 B.n27 VSUBS 0.091619f
C59 B.n28 VSUBS 0.009776f
C60 B.n29 VSUBS 0.009776f
C61 B.n30 VSUBS 0.009776f
C62 B.n31 VSUBS 0.009776f
C63 B.n32 VSUBS 0.005463f
C64 B.n33 VSUBS 0.009776f
C65 B.t7 VSUBS 0.120499f
C66 B.t8 VSUBS 0.142921f
C67 B.t6 VSUBS 0.538169f
C68 B.n34 VSUBS 0.115938f
C69 B.n35 VSUBS 0.091619f
C70 B.n36 VSUBS 0.022649f
C71 B.n37 VSUBS 0.009776f
C72 B.n38 VSUBS 0.009776f
C73 B.n39 VSUBS 0.009776f
C74 B.n40 VSUBS 0.009776f
C75 B.n41 VSUBS 0.009776f
C76 B.n42 VSUBS 0.009776f
C77 B.n43 VSUBS 0.024554f
C78 B.n44 VSUBS 0.009776f
C79 B.n45 VSUBS 0.009776f
C80 B.n46 VSUBS 0.009776f
C81 B.n47 VSUBS 0.009776f
C82 B.n48 VSUBS 0.009776f
C83 B.n49 VSUBS 0.009776f
C84 B.n50 VSUBS 0.009776f
C85 B.n51 VSUBS 0.009776f
C86 B.n52 VSUBS 0.009776f
C87 B.n53 VSUBS 0.009776f
C88 B.n54 VSUBS 0.009776f
C89 B.n55 VSUBS 0.009776f
C90 B.n56 VSUBS 0.009776f
C91 B.n57 VSUBS 0.009776f
C92 B.n58 VSUBS 0.009776f
C93 B.n59 VSUBS 0.009776f
C94 B.n60 VSUBS 0.009776f
C95 B.n61 VSUBS 0.009776f
C96 B.n62 VSUBS 0.009776f
C97 B.n63 VSUBS 0.009776f
C98 B.n64 VSUBS 0.009776f
C99 B.n65 VSUBS 0.009776f
C100 B.n66 VSUBS 0.009776f
C101 B.n67 VSUBS 0.009776f
C102 B.n68 VSUBS 0.009776f
C103 B.n69 VSUBS 0.009776f
C104 B.n70 VSUBS 0.009776f
C105 B.n71 VSUBS 0.009776f
C106 B.n72 VSUBS 0.009776f
C107 B.n73 VSUBS 0.009776f
C108 B.n74 VSUBS 0.009776f
C109 B.n75 VSUBS 0.024813f
C110 B.n76 VSUBS 0.009776f
C111 B.n77 VSUBS 0.009776f
C112 B.n78 VSUBS 0.009776f
C113 B.n79 VSUBS 0.009776f
C114 B.n80 VSUBS 0.009776f
C115 B.n81 VSUBS 0.009776f
C116 B.n82 VSUBS 0.009776f
C117 B.n83 VSUBS 0.0092f
C118 B.n84 VSUBS 0.009776f
C119 B.n85 VSUBS 0.009776f
C120 B.n86 VSUBS 0.009776f
C121 B.n87 VSUBS 0.009776f
C122 B.n88 VSUBS 0.009776f
C123 B.t2 VSUBS 0.120499f
C124 B.t1 VSUBS 0.142922f
C125 B.t0 VSUBS 0.538169f
C126 B.n89 VSUBS 0.115938f
C127 B.n90 VSUBS 0.091619f
C128 B.n91 VSUBS 0.009776f
C129 B.n92 VSUBS 0.009776f
C130 B.n93 VSUBS 0.009776f
C131 B.n94 VSUBS 0.009776f
C132 B.n95 VSUBS 0.009776f
C133 B.n96 VSUBS 0.009776f
C134 B.n97 VSUBS 0.009776f
C135 B.n98 VSUBS 0.024554f
C136 B.n99 VSUBS 0.009776f
C137 B.n100 VSUBS 0.009776f
C138 B.n101 VSUBS 0.009776f
C139 B.n102 VSUBS 0.009776f
C140 B.n103 VSUBS 0.009776f
C141 B.n104 VSUBS 0.009776f
C142 B.n105 VSUBS 0.009776f
C143 B.n106 VSUBS 0.009776f
C144 B.n107 VSUBS 0.009776f
C145 B.n108 VSUBS 0.009776f
C146 B.n109 VSUBS 0.009776f
C147 B.n110 VSUBS 0.009776f
C148 B.n111 VSUBS 0.009776f
C149 B.n112 VSUBS 0.009776f
C150 B.n113 VSUBS 0.009776f
C151 B.n114 VSUBS 0.009776f
C152 B.n115 VSUBS 0.009776f
C153 B.n116 VSUBS 0.009776f
C154 B.n117 VSUBS 0.009776f
C155 B.n118 VSUBS 0.009776f
C156 B.n119 VSUBS 0.009776f
C157 B.n120 VSUBS 0.009776f
C158 B.n121 VSUBS 0.009776f
C159 B.n122 VSUBS 0.009776f
C160 B.n123 VSUBS 0.009776f
C161 B.n124 VSUBS 0.009776f
C162 B.n125 VSUBS 0.009776f
C163 B.n126 VSUBS 0.009776f
C164 B.n127 VSUBS 0.009776f
C165 B.n128 VSUBS 0.009776f
C166 B.n129 VSUBS 0.009776f
C167 B.n130 VSUBS 0.009776f
C168 B.n131 VSUBS 0.009776f
C169 B.n132 VSUBS 0.009776f
C170 B.n133 VSUBS 0.009776f
C171 B.n134 VSUBS 0.009776f
C172 B.n135 VSUBS 0.009776f
C173 B.n136 VSUBS 0.009776f
C174 B.n137 VSUBS 0.009776f
C175 B.n138 VSUBS 0.009776f
C176 B.n139 VSUBS 0.009776f
C177 B.n140 VSUBS 0.009776f
C178 B.n141 VSUBS 0.009776f
C179 B.n142 VSUBS 0.009776f
C180 B.n143 VSUBS 0.009776f
C181 B.n144 VSUBS 0.009776f
C182 B.n145 VSUBS 0.009776f
C183 B.n146 VSUBS 0.009776f
C184 B.n147 VSUBS 0.009776f
C185 B.n148 VSUBS 0.009776f
C186 B.n149 VSUBS 0.009776f
C187 B.n150 VSUBS 0.009776f
C188 B.n151 VSUBS 0.009776f
C189 B.n152 VSUBS 0.009776f
C190 B.n153 VSUBS 0.009776f
C191 B.n154 VSUBS 0.009776f
C192 B.n155 VSUBS 0.009776f
C193 B.n156 VSUBS 0.009776f
C194 B.n157 VSUBS 0.023749f
C195 B.n158 VSUBS 0.023749f
C196 B.n159 VSUBS 0.024554f
C197 B.n160 VSUBS 0.009776f
C198 B.n161 VSUBS 0.009776f
C199 B.n162 VSUBS 0.009776f
C200 B.n163 VSUBS 0.009776f
C201 B.n164 VSUBS 0.009776f
C202 B.n165 VSUBS 0.009776f
C203 B.n166 VSUBS 0.009776f
C204 B.n167 VSUBS 0.009776f
C205 B.n168 VSUBS 0.009776f
C206 B.n169 VSUBS 0.009776f
C207 B.n170 VSUBS 0.009776f
C208 B.n171 VSUBS 0.009776f
C209 B.n172 VSUBS 0.009776f
C210 B.n173 VSUBS 0.009776f
C211 B.n174 VSUBS 0.009776f
C212 B.n175 VSUBS 0.009776f
C213 B.n176 VSUBS 0.009776f
C214 B.n177 VSUBS 0.009776f
C215 B.n178 VSUBS 0.009776f
C216 B.n179 VSUBS 0.009776f
C217 B.n180 VSUBS 0.009776f
C218 B.n181 VSUBS 0.009776f
C219 B.n182 VSUBS 0.0092f
C220 B.n183 VSUBS 0.022649f
C221 B.n184 VSUBS 0.005463f
C222 B.n185 VSUBS 0.009776f
C223 B.n186 VSUBS 0.009776f
C224 B.n187 VSUBS 0.009776f
C225 B.n188 VSUBS 0.009776f
C226 B.n189 VSUBS 0.009776f
C227 B.n190 VSUBS 0.009776f
C228 B.n191 VSUBS 0.009776f
C229 B.n192 VSUBS 0.009776f
C230 B.n193 VSUBS 0.009776f
C231 B.n194 VSUBS 0.009776f
C232 B.n195 VSUBS 0.009776f
C233 B.n196 VSUBS 0.009776f
C234 B.t11 VSUBS 0.120499f
C235 B.t10 VSUBS 0.142921f
C236 B.t9 VSUBS 0.538169f
C237 B.n197 VSUBS 0.115938f
C238 B.n198 VSUBS 0.091619f
C239 B.n199 VSUBS 0.022649f
C240 B.n200 VSUBS 0.005463f
C241 B.n201 VSUBS 0.009776f
C242 B.n202 VSUBS 0.009776f
C243 B.n203 VSUBS 0.009776f
C244 B.n204 VSUBS 0.009776f
C245 B.n205 VSUBS 0.009776f
C246 B.n206 VSUBS 0.009776f
C247 B.n207 VSUBS 0.009776f
C248 B.n208 VSUBS 0.009776f
C249 B.n209 VSUBS 0.009776f
C250 B.n210 VSUBS 0.009776f
C251 B.n211 VSUBS 0.009776f
C252 B.n212 VSUBS 0.009776f
C253 B.n213 VSUBS 0.009776f
C254 B.n214 VSUBS 0.009776f
C255 B.n215 VSUBS 0.009776f
C256 B.n216 VSUBS 0.009776f
C257 B.n217 VSUBS 0.009776f
C258 B.n218 VSUBS 0.009776f
C259 B.n219 VSUBS 0.009776f
C260 B.n220 VSUBS 0.009776f
C261 B.n221 VSUBS 0.009776f
C262 B.n222 VSUBS 0.009776f
C263 B.n223 VSUBS 0.009776f
C264 B.n224 VSUBS 0.023489f
C265 B.n225 VSUBS 0.024554f
C266 B.n226 VSUBS 0.023749f
C267 B.n227 VSUBS 0.009776f
C268 B.n228 VSUBS 0.009776f
C269 B.n229 VSUBS 0.009776f
C270 B.n230 VSUBS 0.009776f
C271 B.n231 VSUBS 0.009776f
C272 B.n232 VSUBS 0.009776f
C273 B.n233 VSUBS 0.009776f
C274 B.n234 VSUBS 0.009776f
C275 B.n235 VSUBS 0.009776f
C276 B.n236 VSUBS 0.009776f
C277 B.n237 VSUBS 0.009776f
C278 B.n238 VSUBS 0.009776f
C279 B.n239 VSUBS 0.009776f
C280 B.n240 VSUBS 0.009776f
C281 B.n241 VSUBS 0.009776f
C282 B.n242 VSUBS 0.009776f
C283 B.n243 VSUBS 0.009776f
C284 B.n244 VSUBS 0.009776f
C285 B.n245 VSUBS 0.009776f
C286 B.n246 VSUBS 0.009776f
C287 B.n247 VSUBS 0.009776f
C288 B.n248 VSUBS 0.009776f
C289 B.n249 VSUBS 0.009776f
C290 B.n250 VSUBS 0.009776f
C291 B.n251 VSUBS 0.009776f
C292 B.n252 VSUBS 0.009776f
C293 B.n253 VSUBS 0.009776f
C294 B.n254 VSUBS 0.009776f
C295 B.n255 VSUBS 0.009776f
C296 B.n256 VSUBS 0.009776f
C297 B.n257 VSUBS 0.009776f
C298 B.n258 VSUBS 0.009776f
C299 B.n259 VSUBS 0.009776f
C300 B.n260 VSUBS 0.009776f
C301 B.n261 VSUBS 0.009776f
C302 B.n262 VSUBS 0.009776f
C303 B.n263 VSUBS 0.009776f
C304 B.n264 VSUBS 0.009776f
C305 B.n265 VSUBS 0.009776f
C306 B.n266 VSUBS 0.009776f
C307 B.n267 VSUBS 0.009776f
C308 B.n268 VSUBS 0.009776f
C309 B.n269 VSUBS 0.009776f
C310 B.n270 VSUBS 0.009776f
C311 B.n271 VSUBS 0.009776f
C312 B.n272 VSUBS 0.009776f
C313 B.n273 VSUBS 0.009776f
C314 B.n274 VSUBS 0.009776f
C315 B.n275 VSUBS 0.009776f
C316 B.n276 VSUBS 0.009776f
C317 B.n277 VSUBS 0.009776f
C318 B.n278 VSUBS 0.009776f
C319 B.n279 VSUBS 0.009776f
C320 B.n280 VSUBS 0.009776f
C321 B.n281 VSUBS 0.009776f
C322 B.n282 VSUBS 0.009776f
C323 B.n283 VSUBS 0.009776f
C324 B.n284 VSUBS 0.009776f
C325 B.n285 VSUBS 0.009776f
C326 B.n286 VSUBS 0.009776f
C327 B.n287 VSUBS 0.009776f
C328 B.n288 VSUBS 0.009776f
C329 B.n289 VSUBS 0.009776f
C330 B.n290 VSUBS 0.009776f
C331 B.n291 VSUBS 0.009776f
C332 B.n292 VSUBS 0.009776f
C333 B.n293 VSUBS 0.009776f
C334 B.n294 VSUBS 0.009776f
C335 B.n295 VSUBS 0.009776f
C336 B.n296 VSUBS 0.009776f
C337 B.n297 VSUBS 0.009776f
C338 B.n298 VSUBS 0.009776f
C339 B.n299 VSUBS 0.009776f
C340 B.n300 VSUBS 0.009776f
C341 B.n301 VSUBS 0.009776f
C342 B.n302 VSUBS 0.009776f
C343 B.n303 VSUBS 0.009776f
C344 B.n304 VSUBS 0.009776f
C345 B.n305 VSUBS 0.009776f
C346 B.n306 VSUBS 0.009776f
C347 B.n307 VSUBS 0.009776f
C348 B.n308 VSUBS 0.009776f
C349 B.n309 VSUBS 0.009776f
C350 B.n310 VSUBS 0.009776f
C351 B.n311 VSUBS 0.009776f
C352 B.n312 VSUBS 0.009776f
C353 B.n313 VSUBS 0.009776f
C354 B.n314 VSUBS 0.009776f
C355 B.n315 VSUBS 0.009776f
C356 B.n316 VSUBS 0.009776f
C357 B.n317 VSUBS 0.009776f
C358 B.n318 VSUBS 0.009776f
C359 B.n319 VSUBS 0.009776f
C360 B.n320 VSUBS 0.023749f
C361 B.n321 VSUBS 0.023749f
C362 B.n322 VSUBS 0.024554f
C363 B.n323 VSUBS 0.009776f
C364 B.n324 VSUBS 0.009776f
C365 B.n325 VSUBS 0.009776f
C366 B.n326 VSUBS 0.009776f
C367 B.n327 VSUBS 0.009776f
C368 B.n328 VSUBS 0.009776f
C369 B.n329 VSUBS 0.009776f
C370 B.n330 VSUBS 0.009776f
C371 B.n331 VSUBS 0.009776f
C372 B.n332 VSUBS 0.009776f
C373 B.n333 VSUBS 0.009776f
C374 B.n334 VSUBS 0.009776f
C375 B.n335 VSUBS 0.009776f
C376 B.n336 VSUBS 0.009776f
C377 B.n337 VSUBS 0.009776f
C378 B.n338 VSUBS 0.009776f
C379 B.n339 VSUBS 0.009776f
C380 B.n340 VSUBS 0.009776f
C381 B.n341 VSUBS 0.009776f
C382 B.n342 VSUBS 0.009776f
C383 B.n343 VSUBS 0.009776f
C384 B.n344 VSUBS 0.0092f
C385 B.n345 VSUBS 0.009776f
C386 B.n346 VSUBS 0.009776f
C387 B.n347 VSUBS 0.009776f
C388 B.n348 VSUBS 0.009776f
C389 B.n349 VSUBS 0.009776f
C390 B.n350 VSUBS 0.009776f
C391 B.n351 VSUBS 0.009776f
C392 B.n352 VSUBS 0.009776f
C393 B.n353 VSUBS 0.009776f
C394 B.n354 VSUBS 0.009776f
C395 B.n355 VSUBS 0.009776f
C396 B.n356 VSUBS 0.009776f
C397 B.n357 VSUBS 0.009776f
C398 B.n358 VSUBS 0.009776f
C399 B.n359 VSUBS 0.009776f
C400 B.n360 VSUBS 0.005463f
C401 B.n361 VSUBS 0.022649f
C402 B.n362 VSUBS 0.0092f
C403 B.n363 VSUBS 0.009776f
C404 B.n364 VSUBS 0.009776f
C405 B.n365 VSUBS 0.009776f
C406 B.n366 VSUBS 0.009776f
C407 B.n367 VSUBS 0.009776f
C408 B.n368 VSUBS 0.009776f
C409 B.n369 VSUBS 0.009776f
C410 B.n370 VSUBS 0.009776f
C411 B.n371 VSUBS 0.009776f
C412 B.n372 VSUBS 0.009776f
C413 B.n373 VSUBS 0.009776f
C414 B.n374 VSUBS 0.009776f
C415 B.n375 VSUBS 0.009776f
C416 B.n376 VSUBS 0.009776f
C417 B.n377 VSUBS 0.009776f
C418 B.n378 VSUBS 0.009776f
C419 B.n379 VSUBS 0.009776f
C420 B.n380 VSUBS 0.009776f
C421 B.n381 VSUBS 0.009776f
C422 B.n382 VSUBS 0.009776f
C423 B.n383 VSUBS 0.009776f
C424 B.n384 VSUBS 0.024554f
C425 B.n385 VSUBS 0.024554f
C426 B.n386 VSUBS 0.023749f
C427 B.n387 VSUBS 0.009776f
C428 B.n388 VSUBS 0.009776f
C429 B.n389 VSUBS 0.009776f
C430 B.n390 VSUBS 0.009776f
C431 B.n391 VSUBS 0.009776f
C432 B.n392 VSUBS 0.009776f
C433 B.n393 VSUBS 0.009776f
C434 B.n394 VSUBS 0.009776f
C435 B.n395 VSUBS 0.009776f
C436 B.n396 VSUBS 0.009776f
C437 B.n397 VSUBS 0.009776f
C438 B.n398 VSUBS 0.009776f
C439 B.n399 VSUBS 0.009776f
C440 B.n400 VSUBS 0.009776f
C441 B.n401 VSUBS 0.009776f
C442 B.n402 VSUBS 0.009776f
C443 B.n403 VSUBS 0.009776f
C444 B.n404 VSUBS 0.009776f
C445 B.n405 VSUBS 0.009776f
C446 B.n406 VSUBS 0.009776f
C447 B.n407 VSUBS 0.009776f
C448 B.n408 VSUBS 0.009776f
C449 B.n409 VSUBS 0.009776f
C450 B.n410 VSUBS 0.009776f
C451 B.n411 VSUBS 0.009776f
C452 B.n412 VSUBS 0.009776f
C453 B.n413 VSUBS 0.009776f
C454 B.n414 VSUBS 0.009776f
C455 B.n415 VSUBS 0.009776f
C456 B.n416 VSUBS 0.009776f
C457 B.n417 VSUBS 0.009776f
C458 B.n418 VSUBS 0.009776f
C459 B.n419 VSUBS 0.009776f
C460 B.n420 VSUBS 0.009776f
C461 B.n421 VSUBS 0.009776f
C462 B.n422 VSUBS 0.009776f
C463 B.n423 VSUBS 0.009776f
C464 B.n424 VSUBS 0.009776f
C465 B.n425 VSUBS 0.009776f
C466 B.n426 VSUBS 0.009776f
C467 B.n427 VSUBS 0.009776f
C468 B.n428 VSUBS 0.009776f
C469 B.n429 VSUBS 0.009776f
C470 B.n430 VSUBS 0.009776f
C471 B.n431 VSUBS 0.012757f
C472 B.n432 VSUBS 0.013589f
C473 B.n433 VSUBS 0.027023f
C474 VDD1.t1 VSUBS 0.049041f
C475 VDD1.t0 VSUBS 0.049041f
C476 VDD1.n0 VSUBS 0.272066f
C477 VDD1.t3 VSUBS 0.049041f
C478 VDD1.t2 VSUBS 0.049041f
C479 VDD1.n1 VSUBS 0.465168f
C480 VP.n0 VSUBS 0.049638f
C481 VP.t1 VSUBS 0.76131f
C482 VP.n1 VSUBS 0.030437f
C483 VP.n2 VSUBS 0.049638f
C484 VP.t0 VSUBS 0.76131f
C485 VP.t3 VSUBS 1.03133f
C486 VP.t2 VSUBS 1.03613f
C487 VP.n3 VSUBS 2.15973f
C488 VP.n4 VSUBS 1.65791f
C489 VP.n5 VSUBS 0.441335f
C490 VP.n6 VSUBS 0.058392f
C491 VP.n7 VSUBS 0.07483f
C492 VP.n8 VSUBS 0.037651f
C493 VP.n9 VSUBS 0.037651f
C494 VP.n10 VSUBS 0.037651f
C495 VP.n11 VSUBS 0.07483f
C496 VP.n12 VSUBS 0.058392f
C497 VP.n13 VSUBS 0.441335f
C498 VP.n14 VSUBS 0.052111f
C499 VDD2.t0 VSUBS 0.051652f
C500 VDD2.t3 VSUBS 0.051652f
C501 VDD2.n0 VSUBS 0.478987f
C502 VDD2.t1 VSUBS 0.051652f
C503 VDD2.t2 VSUBS 0.051652f
C504 VDD2.n1 VSUBS 0.286354f
C505 VDD2.n2 VSUBS 2.18314f
C506 VTAIL.t4 VSUBS 0.42692f
C507 VTAIL.n0 VSUBS 0.476585f
C508 VTAIL.t2 VSUBS 0.42692f
C509 VTAIL.n1 VSUBS 0.556269f
C510 VTAIL.t3 VSUBS 0.42692f
C511 VTAIL.n2 VSUBS 1.21489f
C512 VTAIL.t6 VSUBS 0.426922f
C513 VTAIL.n3 VSUBS 1.21489f
C514 VTAIL.t7 VSUBS 0.426922f
C515 VTAIL.n4 VSUBS 0.556267f
C516 VTAIL.t1 VSUBS 0.426922f
C517 VTAIL.n5 VSUBS 0.556267f
C518 VTAIL.t0 VSUBS 0.42692f
C519 VTAIL.n6 VSUBS 1.21489f
C520 VTAIL.t5 VSUBS 0.42692f
C521 VTAIL.n7 VSUBS 1.12669f
C522 VN.t3 VSUBS 0.983709f
C523 VN.t0 VSUBS 0.979152f
C524 VN.n0 VSUBS 0.627129f
C525 VN.t1 VSUBS 0.983709f
C526 VN.t2 VSUBS 0.979152f
C527 VN.n1 VSUBS 2.06935f
.ends

