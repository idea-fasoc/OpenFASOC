* NGSPICE file created from diff_pair_sample_0534.ext - technology: sky130A

.subckt diff_pair_sample_0534 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=1.0098 ps=6.45 w=6.12 l=3.08
X1 VDD2.t4 VN.t1 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=2.3868 ps=13.02 w=6.12 l=3.08
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=0 ps=0 w=6.12 l=3.08
X3 VTAIL.t2 VP.t0 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=1.0098 ps=6.45 w=6.12 l=3.08
X4 VDD2.t3 VN.t2 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=1.0098 ps=6.45 w=6.12 l=3.08
X5 VTAIL.t8 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=1.0098 ps=6.45 w=6.12 l=3.08
X6 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=0 ps=0 w=6.12 l=3.08
X7 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=2.3868 ps=13.02 w=6.12 l=3.08
X8 VTAIL.t9 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=1.0098 ps=6.45 w=6.12 l=3.08
X9 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=1.0098 ps=6.45 w=6.12 l=3.08
X10 VTAIL.t5 VP.t3 VDD1.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=1.0098 ps=6.45 w=6.12 l=3.08
X11 VDD2.t0 VN.t5 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=2.3868 ps=13.02 w=6.12 l=3.08
X12 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=1.0098 ps=6.45 w=6.12 l=3.08
X13 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=0 ps=0 w=6.12 l=3.08
X14 VDD1.t0 VP.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0098 pd=6.45 as=2.3868 ps=13.02 w=6.12 l=3.08
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3868 pd=13.02 as=0 ps=0 w=6.12 l=3.08
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t5 81.3682
R13 VN.n4 VN.t0 81.3682
R14 VN.n15 VN.n0 70.0803
R15 VN.n31 VN.n16 70.0803
R16 VN.n11 VN.n2 56.5617
R17 VN.n27 VN.n18 56.5617
R18 VN.n5 VN.n4 49.5116
R19 VN.n21 VN.n20 49.5116
R20 VN.n5 VN.t3 47.8875
R21 VN.n0 VN.t1 47.8875
R22 VN.n21 VN.t4 47.8875
R23 VN.n16 VN.t2 47.8875
R24 VN VN.n31 46.411
R25 VN.n6 VN.n5 24.5923
R26 VN.n7 VN.n6 24.5923
R27 VN.n7 VN.n2 24.5923
R28 VN.n12 VN.n11 24.5923
R29 VN.n13 VN.n12 24.5923
R30 VN.n23 VN.n18 24.5923
R31 VN.n23 VN.n22 24.5923
R32 VN.n22 VN.n21 24.5923
R33 VN.n29 VN.n28 24.5923
R34 VN.n28 VN.n27 24.5923
R35 VN.n13 VN.n0 20.1658
R36 VN.n29 VN.n16 20.1658
R37 VN.n20 VN.n19 3.89686
R38 VN.n4 VN.n3 3.89686
R39 VN.n31 VN.n30 0.354861
R40 VN.n15 VN.n14 0.354861
R41 VN VN.n15 0.267071
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n7 VTAIL.t10 54.7458
R53 VTAIL.n10 VTAIL.t0 54.7449
R54 VTAIL.n11 VTAIL.t7 54.7448
R55 VTAIL.n2 VTAIL.t1 54.7448
R56 VTAIL.n9 VTAIL.n8 51.5105
R57 VTAIL.n6 VTAIL.n5 51.5105
R58 VTAIL.n1 VTAIL.n0 51.5104
R59 VTAIL.n4 VTAIL.n3 51.5104
R60 VTAIL.n6 VTAIL.n4 23.5221
R61 VTAIL.n11 VTAIL.n10 20.5824
R62 VTAIL.n0 VTAIL.t6 3.23579
R63 VTAIL.n0 VTAIL.t8 3.23579
R64 VTAIL.n3 VTAIL.t4 3.23579
R65 VTAIL.n3 VTAIL.t5 3.23579
R66 VTAIL.n8 VTAIL.t3 3.23579
R67 VTAIL.n8 VTAIL.t2 3.23579
R68 VTAIL.n5 VTAIL.t11 3.23579
R69 VTAIL.n5 VTAIL.t9 3.23579
R70 VTAIL.n7 VTAIL.n6 2.94016
R71 VTAIL.n10 VTAIL.n9 2.94016
R72 VTAIL.n4 VTAIL.n2 2.94016
R73 VTAIL VTAIL.n11 2.14705
R74 VTAIL.n9 VTAIL.n7 1.94016
R75 VTAIL.n2 VTAIL.n1 1.94016
R76 VTAIL VTAIL.n1 0.793603
R77 VDD2.n1 VDD2.t5 73.573
R78 VDD2.n2 VDD2.t3 71.4246
R79 VDD2.n1 VDD2.n0 68.8688
R80 VDD2 VDD2.n3 68.8651
R81 VDD2.n2 VDD2.n1 38.545
R82 VDD2.n3 VDD2.t1 3.23579
R83 VDD2.n3 VDD2.t0 3.23579
R84 VDD2.n0 VDD2.t2 3.23579
R85 VDD2.n0 VDD2.t4 3.23579
R86 VDD2 VDD2.n2 2.26343
R87 B.n686 B.n685 585
R88 B.n235 B.n118 585
R89 B.n234 B.n233 585
R90 B.n232 B.n231 585
R91 B.n230 B.n229 585
R92 B.n228 B.n227 585
R93 B.n226 B.n225 585
R94 B.n224 B.n223 585
R95 B.n222 B.n221 585
R96 B.n220 B.n219 585
R97 B.n218 B.n217 585
R98 B.n216 B.n215 585
R99 B.n214 B.n213 585
R100 B.n212 B.n211 585
R101 B.n210 B.n209 585
R102 B.n208 B.n207 585
R103 B.n206 B.n205 585
R104 B.n204 B.n203 585
R105 B.n202 B.n201 585
R106 B.n200 B.n199 585
R107 B.n198 B.n197 585
R108 B.n196 B.n195 585
R109 B.n194 B.n193 585
R110 B.n192 B.n191 585
R111 B.n190 B.n189 585
R112 B.n188 B.n187 585
R113 B.n186 B.n185 585
R114 B.n184 B.n183 585
R115 B.n182 B.n181 585
R116 B.n180 B.n179 585
R117 B.n178 B.n177 585
R118 B.n176 B.n175 585
R119 B.n174 B.n173 585
R120 B.n172 B.n171 585
R121 B.n170 B.n169 585
R122 B.n168 B.n167 585
R123 B.n166 B.n165 585
R124 B.n164 B.n163 585
R125 B.n162 B.n161 585
R126 B.n160 B.n159 585
R127 B.n158 B.n157 585
R128 B.n156 B.n155 585
R129 B.n154 B.n153 585
R130 B.n152 B.n151 585
R131 B.n150 B.n149 585
R132 B.n148 B.n147 585
R133 B.n146 B.n145 585
R134 B.n144 B.n143 585
R135 B.n142 B.n141 585
R136 B.n140 B.n139 585
R137 B.n138 B.n137 585
R138 B.n136 B.n135 585
R139 B.n134 B.n133 585
R140 B.n132 B.n131 585
R141 B.n130 B.n129 585
R142 B.n128 B.n127 585
R143 B.n126 B.n125 585
R144 B.n88 B.n87 585
R145 B.n684 B.n89 585
R146 B.n689 B.n89 585
R147 B.n683 B.n682 585
R148 B.n682 B.n85 585
R149 B.n681 B.n84 585
R150 B.n695 B.n84 585
R151 B.n680 B.n83 585
R152 B.n696 B.n83 585
R153 B.n679 B.n82 585
R154 B.n697 B.n82 585
R155 B.n678 B.n677 585
R156 B.n677 B.n78 585
R157 B.n676 B.n77 585
R158 B.n703 B.n77 585
R159 B.n675 B.n76 585
R160 B.n704 B.n76 585
R161 B.n674 B.n75 585
R162 B.n705 B.n75 585
R163 B.n673 B.n672 585
R164 B.n672 B.n71 585
R165 B.n671 B.n70 585
R166 B.n711 B.n70 585
R167 B.n670 B.n69 585
R168 B.n712 B.n69 585
R169 B.n669 B.n68 585
R170 B.n713 B.n68 585
R171 B.n668 B.n667 585
R172 B.n667 B.n64 585
R173 B.n666 B.n63 585
R174 B.n719 B.n63 585
R175 B.n665 B.n62 585
R176 B.n720 B.n62 585
R177 B.n664 B.n61 585
R178 B.n721 B.n61 585
R179 B.n663 B.n662 585
R180 B.n662 B.n57 585
R181 B.n661 B.n56 585
R182 B.n727 B.n56 585
R183 B.n660 B.n55 585
R184 B.n728 B.n55 585
R185 B.n659 B.n54 585
R186 B.n729 B.n54 585
R187 B.n658 B.n657 585
R188 B.n657 B.n53 585
R189 B.n656 B.n49 585
R190 B.n735 B.n49 585
R191 B.n655 B.n48 585
R192 B.n736 B.n48 585
R193 B.n654 B.n47 585
R194 B.n737 B.n47 585
R195 B.n653 B.n652 585
R196 B.n652 B.n43 585
R197 B.n651 B.n42 585
R198 B.n743 B.n42 585
R199 B.n650 B.n41 585
R200 B.n744 B.n41 585
R201 B.n649 B.n40 585
R202 B.n745 B.n40 585
R203 B.n648 B.n647 585
R204 B.n647 B.n36 585
R205 B.n646 B.n35 585
R206 B.n751 B.n35 585
R207 B.n645 B.n34 585
R208 B.n752 B.n34 585
R209 B.n644 B.n33 585
R210 B.n753 B.n33 585
R211 B.n643 B.n642 585
R212 B.n642 B.n29 585
R213 B.n641 B.n28 585
R214 B.n759 B.n28 585
R215 B.n640 B.n27 585
R216 B.n760 B.n27 585
R217 B.n639 B.n26 585
R218 B.n761 B.n26 585
R219 B.n638 B.n637 585
R220 B.n637 B.n22 585
R221 B.n636 B.n21 585
R222 B.n767 B.n21 585
R223 B.n635 B.n20 585
R224 B.n768 B.n20 585
R225 B.n634 B.n19 585
R226 B.n769 B.n19 585
R227 B.n633 B.n632 585
R228 B.n632 B.n18 585
R229 B.n631 B.n14 585
R230 B.n775 B.n14 585
R231 B.n630 B.n13 585
R232 B.n776 B.n13 585
R233 B.n629 B.n12 585
R234 B.n777 B.n12 585
R235 B.n628 B.n627 585
R236 B.n627 B.n8 585
R237 B.n626 B.n7 585
R238 B.n783 B.n7 585
R239 B.n625 B.n6 585
R240 B.n784 B.n6 585
R241 B.n624 B.n5 585
R242 B.n785 B.n5 585
R243 B.n623 B.n622 585
R244 B.n622 B.n4 585
R245 B.n621 B.n236 585
R246 B.n621 B.n620 585
R247 B.n611 B.n237 585
R248 B.n238 B.n237 585
R249 B.n613 B.n612 585
R250 B.n614 B.n613 585
R251 B.n610 B.n243 585
R252 B.n243 B.n242 585
R253 B.n609 B.n608 585
R254 B.n608 B.n607 585
R255 B.n245 B.n244 585
R256 B.n600 B.n245 585
R257 B.n599 B.n598 585
R258 B.n601 B.n599 585
R259 B.n597 B.n250 585
R260 B.n250 B.n249 585
R261 B.n596 B.n595 585
R262 B.n595 B.n594 585
R263 B.n252 B.n251 585
R264 B.n253 B.n252 585
R265 B.n587 B.n586 585
R266 B.n588 B.n587 585
R267 B.n585 B.n258 585
R268 B.n258 B.n257 585
R269 B.n584 B.n583 585
R270 B.n583 B.n582 585
R271 B.n260 B.n259 585
R272 B.n261 B.n260 585
R273 B.n575 B.n574 585
R274 B.n576 B.n575 585
R275 B.n573 B.n265 585
R276 B.n269 B.n265 585
R277 B.n572 B.n571 585
R278 B.n571 B.n570 585
R279 B.n267 B.n266 585
R280 B.n268 B.n267 585
R281 B.n563 B.n562 585
R282 B.n564 B.n563 585
R283 B.n561 B.n274 585
R284 B.n274 B.n273 585
R285 B.n560 B.n559 585
R286 B.n559 B.n558 585
R287 B.n276 B.n275 585
R288 B.n277 B.n276 585
R289 B.n551 B.n550 585
R290 B.n552 B.n551 585
R291 B.n549 B.n282 585
R292 B.n282 B.n281 585
R293 B.n548 B.n547 585
R294 B.n547 B.n546 585
R295 B.n284 B.n283 585
R296 B.n539 B.n284 585
R297 B.n538 B.n537 585
R298 B.n540 B.n538 585
R299 B.n536 B.n289 585
R300 B.n289 B.n288 585
R301 B.n535 B.n534 585
R302 B.n534 B.n533 585
R303 B.n291 B.n290 585
R304 B.n292 B.n291 585
R305 B.n526 B.n525 585
R306 B.n527 B.n526 585
R307 B.n524 B.n297 585
R308 B.n297 B.n296 585
R309 B.n523 B.n522 585
R310 B.n522 B.n521 585
R311 B.n299 B.n298 585
R312 B.n300 B.n299 585
R313 B.n514 B.n513 585
R314 B.n515 B.n514 585
R315 B.n512 B.n305 585
R316 B.n305 B.n304 585
R317 B.n511 B.n510 585
R318 B.n510 B.n509 585
R319 B.n307 B.n306 585
R320 B.n308 B.n307 585
R321 B.n502 B.n501 585
R322 B.n503 B.n502 585
R323 B.n500 B.n313 585
R324 B.n313 B.n312 585
R325 B.n499 B.n498 585
R326 B.n498 B.n497 585
R327 B.n315 B.n314 585
R328 B.n316 B.n315 585
R329 B.n490 B.n489 585
R330 B.n491 B.n490 585
R331 B.n488 B.n321 585
R332 B.n321 B.n320 585
R333 B.n487 B.n486 585
R334 B.n486 B.n485 585
R335 B.n323 B.n322 585
R336 B.n324 B.n323 585
R337 B.n478 B.n477 585
R338 B.n479 B.n478 585
R339 B.n327 B.n326 585
R340 B.n362 B.n360 585
R341 B.n363 B.n359 585
R342 B.n363 B.n328 585
R343 B.n366 B.n365 585
R344 B.n367 B.n358 585
R345 B.n369 B.n368 585
R346 B.n371 B.n357 585
R347 B.n374 B.n373 585
R348 B.n375 B.n356 585
R349 B.n377 B.n376 585
R350 B.n379 B.n355 585
R351 B.n382 B.n381 585
R352 B.n383 B.n354 585
R353 B.n385 B.n384 585
R354 B.n387 B.n353 585
R355 B.n390 B.n389 585
R356 B.n391 B.n352 585
R357 B.n393 B.n392 585
R358 B.n395 B.n351 585
R359 B.n398 B.n397 585
R360 B.n399 B.n350 585
R361 B.n401 B.n400 585
R362 B.n403 B.n349 585
R363 B.n406 B.n405 585
R364 B.n408 B.n346 585
R365 B.n410 B.n409 585
R366 B.n412 B.n345 585
R367 B.n415 B.n414 585
R368 B.n416 B.n344 585
R369 B.n418 B.n417 585
R370 B.n420 B.n343 585
R371 B.n423 B.n422 585
R372 B.n424 B.n342 585
R373 B.n429 B.n428 585
R374 B.n431 B.n341 585
R375 B.n434 B.n433 585
R376 B.n435 B.n340 585
R377 B.n437 B.n436 585
R378 B.n439 B.n339 585
R379 B.n442 B.n441 585
R380 B.n443 B.n338 585
R381 B.n445 B.n444 585
R382 B.n447 B.n337 585
R383 B.n450 B.n449 585
R384 B.n451 B.n336 585
R385 B.n453 B.n452 585
R386 B.n455 B.n335 585
R387 B.n458 B.n457 585
R388 B.n459 B.n334 585
R389 B.n461 B.n460 585
R390 B.n463 B.n333 585
R391 B.n466 B.n465 585
R392 B.n467 B.n332 585
R393 B.n469 B.n468 585
R394 B.n471 B.n331 585
R395 B.n472 B.n330 585
R396 B.n475 B.n474 585
R397 B.n476 B.n329 585
R398 B.n329 B.n328 585
R399 B.n481 B.n480 585
R400 B.n480 B.n479 585
R401 B.n482 B.n325 585
R402 B.n325 B.n324 585
R403 B.n484 B.n483 585
R404 B.n485 B.n484 585
R405 B.n319 B.n318 585
R406 B.n320 B.n319 585
R407 B.n493 B.n492 585
R408 B.n492 B.n491 585
R409 B.n494 B.n317 585
R410 B.n317 B.n316 585
R411 B.n496 B.n495 585
R412 B.n497 B.n496 585
R413 B.n311 B.n310 585
R414 B.n312 B.n311 585
R415 B.n505 B.n504 585
R416 B.n504 B.n503 585
R417 B.n506 B.n309 585
R418 B.n309 B.n308 585
R419 B.n508 B.n507 585
R420 B.n509 B.n508 585
R421 B.n303 B.n302 585
R422 B.n304 B.n303 585
R423 B.n517 B.n516 585
R424 B.n516 B.n515 585
R425 B.n518 B.n301 585
R426 B.n301 B.n300 585
R427 B.n520 B.n519 585
R428 B.n521 B.n520 585
R429 B.n295 B.n294 585
R430 B.n296 B.n295 585
R431 B.n529 B.n528 585
R432 B.n528 B.n527 585
R433 B.n530 B.n293 585
R434 B.n293 B.n292 585
R435 B.n532 B.n531 585
R436 B.n533 B.n532 585
R437 B.n287 B.n286 585
R438 B.n288 B.n287 585
R439 B.n542 B.n541 585
R440 B.n541 B.n540 585
R441 B.n543 B.n285 585
R442 B.n539 B.n285 585
R443 B.n545 B.n544 585
R444 B.n546 B.n545 585
R445 B.n280 B.n279 585
R446 B.n281 B.n280 585
R447 B.n554 B.n553 585
R448 B.n553 B.n552 585
R449 B.n555 B.n278 585
R450 B.n278 B.n277 585
R451 B.n557 B.n556 585
R452 B.n558 B.n557 585
R453 B.n272 B.n271 585
R454 B.n273 B.n272 585
R455 B.n566 B.n565 585
R456 B.n565 B.n564 585
R457 B.n567 B.n270 585
R458 B.n270 B.n268 585
R459 B.n569 B.n568 585
R460 B.n570 B.n569 585
R461 B.n264 B.n263 585
R462 B.n269 B.n264 585
R463 B.n578 B.n577 585
R464 B.n577 B.n576 585
R465 B.n579 B.n262 585
R466 B.n262 B.n261 585
R467 B.n581 B.n580 585
R468 B.n582 B.n581 585
R469 B.n256 B.n255 585
R470 B.n257 B.n256 585
R471 B.n590 B.n589 585
R472 B.n589 B.n588 585
R473 B.n591 B.n254 585
R474 B.n254 B.n253 585
R475 B.n593 B.n592 585
R476 B.n594 B.n593 585
R477 B.n248 B.n247 585
R478 B.n249 B.n248 585
R479 B.n603 B.n602 585
R480 B.n602 B.n601 585
R481 B.n604 B.n246 585
R482 B.n600 B.n246 585
R483 B.n606 B.n605 585
R484 B.n607 B.n606 585
R485 B.n241 B.n240 585
R486 B.n242 B.n241 585
R487 B.n616 B.n615 585
R488 B.n615 B.n614 585
R489 B.n617 B.n239 585
R490 B.n239 B.n238 585
R491 B.n619 B.n618 585
R492 B.n620 B.n619 585
R493 B.n2 B.n0 585
R494 B.n4 B.n2 585
R495 B.n3 B.n1 585
R496 B.n784 B.n3 585
R497 B.n782 B.n781 585
R498 B.n783 B.n782 585
R499 B.n780 B.n9 585
R500 B.n9 B.n8 585
R501 B.n779 B.n778 585
R502 B.n778 B.n777 585
R503 B.n11 B.n10 585
R504 B.n776 B.n11 585
R505 B.n774 B.n773 585
R506 B.n775 B.n774 585
R507 B.n772 B.n15 585
R508 B.n18 B.n15 585
R509 B.n771 B.n770 585
R510 B.n770 B.n769 585
R511 B.n17 B.n16 585
R512 B.n768 B.n17 585
R513 B.n766 B.n765 585
R514 B.n767 B.n766 585
R515 B.n764 B.n23 585
R516 B.n23 B.n22 585
R517 B.n763 B.n762 585
R518 B.n762 B.n761 585
R519 B.n25 B.n24 585
R520 B.n760 B.n25 585
R521 B.n758 B.n757 585
R522 B.n759 B.n758 585
R523 B.n756 B.n30 585
R524 B.n30 B.n29 585
R525 B.n755 B.n754 585
R526 B.n754 B.n753 585
R527 B.n32 B.n31 585
R528 B.n752 B.n32 585
R529 B.n750 B.n749 585
R530 B.n751 B.n750 585
R531 B.n748 B.n37 585
R532 B.n37 B.n36 585
R533 B.n747 B.n746 585
R534 B.n746 B.n745 585
R535 B.n39 B.n38 585
R536 B.n744 B.n39 585
R537 B.n742 B.n741 585
R538 B.n743 B.n742 585
R539 B.n740 B.n44 585
R540 B.n44 B.n43 585
R541 B.n739 B.n738 585
R542 B.n738 B.n737 585
R543 B.n46 B.n45 585
R544 B.n736 B.n46 585
R545 B.n734 B.n733 585
R546 B.n735 B.n734 585
R547 B.n732 B.n50 585
R548 B.n53 B.n50 585
R549 B.n731 B.n730 585
R550 B.n730 B.n729 585
R551 B.n52 B.n51 585
R552 B.n728 B.n52 585
R553 B.n726 B.n725 585
R554 B.n727 B.n726 585
R555 B.n724 B.n58 585
R556 B.n58 B.n57 585
R557 B.n723 B.n722 585
R558 B.n722 B.n721 585
R559 B.n60 B.n59 585
R560 B.n720 B.n60 585
R561 B.n718 B.n717 585
R562 B.n719 B.n718 585
R563 B.n716 B.n65 585
R564 B.n65 B.n64 585
R565 B.n715 B.n714 585
R566 B.n714 B.n713 585
R567 B.n67 B.n66 585
R568 B.n712 B.n67 585
R569 B.n710 B.n709 585
R570 B.n711 B.n710 585
R571 B.n708 B.n72 585
R572 B.n72 B.n71 585
R573 B.n707 B.n706 585
R574 B.n706 B.n705 585
R575 B.n74 B.n73 585
R576 B.n704 B.n74 585
R577 B.n702 B.n701 585
R578 B.n703 B.n702 585
R579 B.n700 B.n79 585
R580 B.n79 B.n78 585
R581 B.n699 B.n698 585
R582 B.n698 B.n697 585
R583 B.n81 B.n80 585
R584 B.n696 B.n81 585
R585 B.n694 B.n693 585
R586 B.n695 B.n694 585
R587 B.n692 B.n86 585
R588 B.n86 B.n85 585
R589 B.n691 B.n690 585
R590 B.n690 B.n689 585
R591 B.n787 B.n786 585
R592 B.n786 B.n785 585
R593 B.n480 B.n327 554.963
R594 B.n690 B.n88 554.963
R595 B.n478 B.n329 554.963
R596 B.n686 B.n89 554.963
R597 B.n688 B.n687 256.663
R598 B.n688 B.n117 256.663
R599 B.n688 B.n116 256.663
R600 B.n688 B.n115 256.663
R601 B.n688 B.n114 256.663
R602 B.n688 B.n113 256.663
R603 B.n688 B.n112 256.663
R604 B.n688 B.n111 256.663
R605 B.n688 B.n110 256.663
R606 B.n688 B.n109 256.663
R607 B.n688 B.n108 256.663
R608 B.n688 B.n107 256.663
R609 B.n688 B.n106 256.663
R610 B.n688 B.n105 256.663
R611 B.n688 B.n104 256.663
R612 B.n688 B.n103 256.663
R613 B.n688 B.n102 256.663
R614 B.n688 B.n101 256.663
R615 B.n688 B.n100 256.663
R616 B.n688 B.n99 256.663
R617 B.n688 B.n98 256.663
R618 B.n688 B.n97 256.663
R619 B.n688 B.n96 256.663
R620 B.n688 B.n95 256.663
R621 B.n688 B.n94 256.663
R622 B.n688 B.n93 256.663
R623 B.n688 B.n92 256.663
R624 B.n688 B.n91 256.663
R625 B.n688 B.n90 256.663
R626 B.n361 B.n328 256.663
R627 B.n364 B.n328 256.663
R628 B.n370 B.n328 256.663
R629 B.n372 B.n328 256.663
R630 B.n378 B.n328 256.663
R631 B.n380 B.n328 256.663
R632 B.n386 B.n328 256.663
R633 B.n388 B.n328 256.663
R634 B.n394 B.n328 256.663
R635 B.n396 B.n328 256.663
R636 B.n402 B.n328 256.663
R637 B.n404 B.n328 256.663
R638 B.n411 B.n328 256.663
R639 B.n413 B.n328 256.663
R640 B.n419 B.n328 256.663
R641 B.n421 B.n328 256.663
R642 B.n430 B.n328 256.663
R643 B.n432 B.n328 256.663
R644 B.n438 B.n328 256.663
R645 B.n440 B.n328 256.663
R646 B.n446 B.n328 256.663
R647 B.n448 B.n328 256.663
R648 B.n454 B.n328 256.663
R649 B.n456 B.n328 256.663
R650 B.n462 B.n328 256.663
R651 B.n464 B.n328 256.663
R652 B.n470 B.n328 256.663
R653 B.n473 B.n328 256.663
R654 B.n425 B.t10 256.56
R655 B.n347 B.t14 256.56
R656 B.n122 B.t6 256.56
R657 B.n119 B.t17 256.56
R658 B.n480 B.n325 163.367
R659 B.n484 B.n325 163.367
R660 B.n484 B.n319 163.367
R661 B.n492 B.n319 163.367
R662 B.n492 B.n317 163.367
R663 B.n496 B.n317 163.367
R664 B.n496 B.n311 163.367
R665 B.n504 B.n311 163.367
R666 B.n504 B.n309 163.367
R667 B.n508 B.n309 163.367
R668 B.n508 B.n303 163.367
R669 B.n516 B.n303 163.367
R670 B.n516 B.n301 163.367
R671 B.n520 B.n301 163.367
R672 B.n520 B.n295 163.367
R673 B.n528 B.n295 163.367
R674 B.n528 B.n293 163.367
R675 B.n532 B.n293 163.367
R676 B.n532 B.n287 163.367
R677 B.n541 B.n287 163.367
R678 B.n541 B.n285 163.367
R679 B.n545 B.n285 163.367
R680 B.n545 B.n280 163.367
R681 B.n553 B.n280 163.367
R682 B.n553 B.n278 163.367
R683 B.n557 B.n278 163.367
R684 B.n557 B.n272 163.367
R685 B.n565 B.n272 163.367
R686 B.n565 B.n270 163.367
R687 B.n569 B.n270 163.367
R688 B.n569 B.n264 163.367
R689 B.n577 B.n264 163.367
R690 B.n577 B.n262 163.367
R691 B.n581 B.n262 163.367
R692 B.n581 B.n256 163.367
R693 B.n589 B.n256 163.367
R694 B.n589 B.n254 163.367
R695 B.n593 B.n254 163.367
R696 B.n593 B.n248 163.367
R697 B.n602 B.n248 163.367
R698 B.n602 B.n246 163.367
R699 B.n606 B.n246 163.367
R700 B.n606 B.n241 163.367
R701 B.n615 B.n241 163.367
R702 B.n615 B.n239 163.367
R703 B.n619 B.n239 163.367
R704 B.n619 B.n2 163.367
R705 B.n786 B.n2 163.367
R706 B.n786 B.n3 163.367
R707 B.n782 B.n3 163.367
R708 B.n782 B.n9 163.367
R709 B.n778 B.n9 163.367
R710 B.n778 B.n11 163.367
R711 B.n774 B.n11 163.367
R712 B.n774 B.n15 163.367
R713 B.n770 B.n15 163.367
R714 B.n770 B.n17 163.367
R715 B.n766 B.n17 163.367
R716 B.n766 B.n23 163.367
R717 B.n762 B.n23 163.367
R718 B.n762 B.n25 163.367
R719 B.n758 B.n25 163.367
R720 B.n758 B.n30 163.367
R721 B.n754 B.n30 163.367
R722 B.n754 B.n32 163.367
R723 B.n750 B.n32 163.367
R724 B.n750 B.n37 163.367
R725 B.n746 B.n37 163.367
R726 B.n746 B.n39 163.367
R727 B.n742 B.n39 163.367
R728 B.n742 B.n44 163.367
R729 B.n738 B.n44 163.367
R730 B.n738 B.n46 163.367
R731 B.n734 B.n46 163.367
R732 B.n734 B.n50 163.367
R733 B.n730 B.n50 163.367
R734 B.n730 B.n52 163.367
R735 B.n726 B.n52 163.367
R736 B.n726 B.n58 163.367
R737 B.n722 B.n58 163.367
R738 B.n722 B.n60 163.367
R739 B.n718 B.n60 163.367
R740 B.n718 B.n65 163.367
R741 B.n714 B.n65 163.367
R742 B.n714 B.n67 163.367
R743 B.n710 B.n67 163.367
R744 B.n710 B.n72 163.367
R745 B.n706 B.n72 163.367
R746 B.n706 B.n74 163.367
R747 B.n702 B.n74 163.367
R748 B.n702 B.n79 163.367
R749 B.n698 B.n79 163.367
R750 B.n698 B.n81 163.367
R751 B.n694 B.n81 163.367
R752 B.n694 B.n86 163.367
R753 B.n690 B.n86 163.367
R754 B.n363 B.n362 163.367
R755 B.n365 B.n363 163.367
R756 B.n369 B.n358 163.367
R757 B.n373 B.n371 163.367
R758 B.n377 B.n356 163.367
R759 B.n381 B.n379 163.367
R760 B.n385 B.n354 163.367
R761 B.n389 B.n387 163.367
R762 B.n393 B.n352 163.367
R763 B.n397 B.n395 163.367
R764 B.n401 B.n350 163.367
R765 B.n405 B.n403 163.367
R766 B.n410 B.n346 163.367
R767 B.n414 B.n412 163.367
R768 B.n418 B.n344 163.367
R769 B.n422 B.n420 163.367
R770 B.n429 B.n342 163.367
R771 B.n433 B.n431 163.367
R772 B.n437 B.n340 163.367
R773 B.n441 B.n439 163.367
R774 B.n445 B.n338 163.367
R775 B.n449 B.n447 163.367
R776 B.n453 B.n336 163.367
R777 B.n457 B.n455 163.367
R778 B.n461 B.n334 163.367
R779 B.n465 B.n463 163.367
R780 B.n469 B.n332 163.367
R781 B.n472 B.n471 163.367
R782 B.n474 B.n329 163.367
R783 B.n478 B.n323 163.367
R784 B.n486 B.n323 163.367
R785 B.n486 B.n321 163.367
R786 B.n490 B.n321 163.367
R787 B.n490 B.n315 163.367
R788 B.n498 B.n315 163.367
R789 B.n498 B.n313 163.367
R790 B.n502 B.n313 163.367
R791 B.n502 B.n307 163.367
R792 B.n510 B.n307 163.367
R793 B.n510 B.n305 163.367
R794 B.n514 B.n305 163.367
R795 B.n514 B.n299 163.367
R796 B.n522 B.n299 163.367
R797 B.n522 B.n297 163.367
R798 B.n526 B.n297 163.367
R799 B.n526 B.n291 163.367
R800 B.n534 B.n291 163.367
R801 B.n534 B.n289 163.367
R802 B.n538 B.n289 163.367
R803 B.n538 B.n284 163.367
R804 B.n547 B.n284 163.367
R805 B.n547 B.n282 163.367
R806 B.n551 B.n282 163.367
R807 B.n551 B.n276 163.367
R808 B.n559 B.n276 163.367
R809 B.n559 B.n274 163.367
R810 B.n563 B.n274 163.367
R811 B.n563 B.n267 163.367
R812 B.n571 B.n267 163.367
R813 B.n571 B.n265 163.367
R814 B.n575 B.n265 163.367
R815 B.n575 B.n260 163.367
R816 B.n583 B.n260 163.367
R817 B.n583 B.n258 163.367
R818 B.n587 B.n258 163.367
R819 B.n587 B.n252 163.367
R820 B.n595 B.n252 163.367
R821 B.n595 B.n250 163.367
R822 B.n599 B.n250 163.367
R823 B.n599 B.n245 163.367
R824 B.n608 B.n245 163.367
R825 B.n608 B.n243 163.367
R826 B.n613 B.n243 163.367
R827 B.n613 B.n237 163.367
R828 B.n621 B.n237 163.367
R829 B.n622 B.n621 163.367
R830 B.n622 B.n5 163.367
R831 B.n6 B.n5 163.367
R832 B.n7 B.n6 163.367
R833 B.n627 B.n7 163.367
R834 B.n627 B.n12 163.367
R835 B.n13 B.n12 163.367
R836 B.n14 B.n13 163.367
R837 B.n632 B.n14 163.367
R838 B.n632 B.n19 163.367
R839 B.n20 B.n19 163.367
R840 B.n21 B.n20 163.367
R841 B.n637 B.n21 163.367
R842 B.n637 B.n26 163.367
R843 B.n27 B.n26 163.367
R844 B.n28 B.n27 163.367
R845 B.n642 B.n28 163.367
R846 B.n642 B.n33 163.367
R847 B.n34 B.n33 163.367
R848 B.n35 B.n34 163.367
R849 B.n647 B.n35 163.367
R850 B.n647 B.n40 163.367
R851 B.n41 B.n40 163.367
R852 B.n42 B.n41 163.367
R853 B.n652 B.n42 163.367
R854 B.n652 B.n47 163.367
R855 B.n48 B.n47 163.367
R856 B.n49 B.n48 163.367
R857 B.n657 B.n49 163.367
R858 B.n657 B.n54 163.367
R859 B.n55 B.n54 163.367
R860 B.n56 B.n55 163.367
R861 B.n662 B.n56 163.367
R862 B.n662 B.n61 163.367
R863 B.n62 B.n61 163.367
R864 B.n63 B.n62 163.367
R865 B.n667 B.n63 163.367
R866 B.n667 B.n68 163.367
R867 B.n69 B.n68 163.367
R868 B.n70 B.n69 163.367
R869 B.n672 B.n70 163.367
R870 B.n672 B.n75 163.367
R871 B.n76 B.n75 163.367
R872 B.n77 B.n76 163.367
R873 B.n677 B.n77 163.367
R874 B.n677 B.n82 163.367
R875 B.n83 B.n82 163.367
R876 B.n84 B.n83 163.367
R877 B.n682 B.n84 163.367
R878 B.n682 B.n89 163.367
R879 B.n127 B.n126 163.367
R880 B.n131 B.n130 163.367
R881 B.n135 B.n134 163.367
R882 B.n139 B.n138 163.367
R883 B.n143 B.n142 163.367
R884 B.n147 B.n146 163.367
R885 B.n151 B.n150 163.367
R886 B.n155 B.n154 163.367
R887 B.n159 B.n158 163.367
R888 B.n163 B.n162 163.367
R889 B.n167 B.n166 163.367
R890 B.n171 B.n170 163.367
R891 B.n175 B.n174 163.367
R892 B.n179 B.n178 163.367
R893 B.n183 B.n182 163.367
R894 B.n187 B.n186 163.367
R895 B.n191 B.n190 163.367
R896 B.n195 B.n194 163.367
R897 B.n199 B.n198 163.367
R898 B.n203 B.n202 163.367
R899 B.n207 B.n206 163.367
R900 B.n211 B.n210 163.367
R901 B.n215 B.n214 163.367
R902 B.n219 B.n218 163.367
R903 B.n223 B.n222 163.367
R904 B.n227 B.n226 163.367
R905 B.n231 B.n230 163.367
R906 B.n233 B.n118 163.367
R907 B.n425 B.t13 135.512
R908 B.n119 B.t18 135.512
R909 B.n347 B.t16 135.505
R910 B.n122 B.t8 135.505
R911 B.n479 B.n328 134.183
R912 B.n689 B.n688 134.183
R913 B.n361 B.n327 71.676
R914 B.n365 B.n364 71.676
R915 B.n370 B.n369 71.676
R916 B.n373 B.n372 71.676
R917 B.n378 B.n377 71.676
R918 B.n381 B.n380 71.676
R919 B.n386 B.n385 71.676
R920 B.n389 B.n388 71.676
R921 B.n394 B.n393 71.676
R922 B.n397 B.n396 71.676
R923 B.n402 B.n401 71.676
R924 B.n405 B.n404 71.676
R925 B.n411 B.n410 71.676
R926 B.n414 B.n413 71.676
R927 B.n419 B.n418 71.676
R928 B.n422 B.n421 71.676
R929 B.n430 B.n429 71.676
R930 B.n433 B.n432 71.676
R931 B.n438 B.n437 71.676
R932 B.n441 B.n440 71.676
R933 B.n446 B.n445 71.676
R934 B.n449 B.n448 71.676
R935 B.n454 B.n453 71.676
R936 B.n457 B.n456 71.676
R937 B.n462 B.n461 71.676
R938 B.n465 B.n464 71.676
R939 B.n470 B.n469 71.676
R940 B.n473 B.n472 71.676
R941 B.n90 B.n88 71.676
R942 B.n127 B.n91 71.676
R943 B.n131 B.n92 71.676
R944 B.n135 B.n93 71.676
R945 B.n139 B.n94 71.676
R946 B.n143 B.n95 71.676
R947 B.n147 B.n96 71.676
R948 B.n151 B.n97 71.676
R949 B.n155 B.n98 71.676
R950 B.n159 B.n99 71.676
R951 B.n163 B.n100 71.676
R952 B.n167 B.n101 71.676
R953 B.n171 B.n102 71.676
R954 B.n175 B.n103 71.676
R955 B.n179 B.n104 71.676
R956 B.n183 B.n105 71.676
R957 B.n187 B.n106 71.676
R958 B.n191 B.n107 71.676
R959 B.n195 B.n108 71.676
R960 B.n199 B.n109 71.676
R961 B.n203 B.n110 71.676
R962 B.n207 B.n111 71.676
R963 B.n211 B.n112 71.676
R964 B.n215 B.n113 71.676
R965 B.n219 B.n114 71.676
R966 B.n223 B.n115 71.676
R967 B.n227 B.n116 71.676
R968 B.n231 B.n117 71.676
R969 B.n687 B.n118 71.676
R970 B.n687 B.n686 71.676
R971 B.n233 B.n117 71.676
R972 B.n230 B.n116 71.676
R973 B.n226 B.n115 71.676
R974 B.n222 B.n114 71.676
R975 B.n218 B.n113 71.676
R976 B.n214 B.n112 71.676
R977 B.n210 B.n111 71.676
R978 B.n206 B.n110 71.676
R979 B.n202 B.n109 71.676
R980 B.n198 B.n108 71.676
R981 B.n194 B.n107 71.676
R982 B.n190 B.n106 71.676
R983 B.n186 B.n105 71.676
R984 B.n182 B.n104 71.676
R985 B.n178 B.n103 71.676
R986 B.n174 B.n102 71.676
R987 B.n170 B.n101 71.676
R988 B.n166 B.n100 71.676
R989 B.n162 B.n99 71.676
R990 B.n158 B.n98 71.676
R991 B.n154 B.n97 71.676
R992 B.n150 B.n96 71.676
R993 B.n146 B.n95 71.676
R994 B.n142 B.n94 71.676
R995 B.n138 B.n93 71.676
R996 B.n134 B.n92 71.676
R997 B.n130 B.n91 71.676
R998 B.n126 B.n90 71.676
R999 B.n362 B.n361 71.676
R1000 B.n364 B.n358 71.676
R1001 B.n371 B.n370 71.676
R1002 B.n372 B.n356 71.676
R1003 B.n379 B.n378 71.676
R1004 B.n380 B.n354 71.676
R1005 B.n387 B.n386 71.676
R1006 B.n388 B.n352 71.676
R1007 B.n395 B.n394 71.676
R1008 B.n396 B.n350 71.676
R1009 B.n403 B.n402 71.676
R1010 B.n404 B.n346 71.676
R1011 B.n412 B.n411 71.676
R1012 B.n413 B.n344 71.676
R1013 B.n420 B.n419 71.676
R1014 B.n421 B.n342 71.676
R1015 B.n431 B.n430 71.676
R1016 B.n432 B.n340 71.676
R1017 B.n439 B.n438 71.676
R1018 B.n440 B.n338 71.676
R1019 B.n447 B.n446 71.676
R1020 B.n448 B.n336 71.676
R1021 B.n455 B.n454 71.676
R1022 B.n456 B.n334 71.676
R1023 B.n463 B.n462 71.676
R1024 B.n464 B.n332 71.676
R1025 B.n471 B.n470 71.676
R1026 B.n474 B.n473 71.676
R1027 B.n426 B.t12 69.3784
R1028 B.n120 B.t19 69.3784
R1029 B.n348 B.t15 69.3716
R1030 B.n123 B.t9 69.3716
R1031 B.n426 B.n425 66.1338
R1032 B.n348 B.n347 66.1338
R1033 B.n123 B.n122 66.1338
R1034 B.n120 B.n119 66.1338
R1035 B.n479 B.n324 65.6433
R1036 B.n485 B.n324 65.6433
R1037 B.n485 B.n320 65.6433
R1038 B.n491 B.n320 65.6433
R1039 B.n491 B.n316 65.6433
R1040 B.n497 B.n316 65.6433
R1041 B.n497 B.n312 65.6433
R1042 B.n503 B.n312 65.6433
R1043 B.n509 B.n308 65.6433
R1044 B.n509 B.n304 65.6433
R1045 B.n515 B.n304 65.6433
R1046 B.n515 B.n300 65.6433
R1047 B.n521 B.n300 65.6433
R1048 B.n521 B.n296 65.6433
R1049 B.n527 B.n296 65.6433
R1050 B.n527 B.n292 65.6433
R1051 B.n533 B.n292 65.6433
R1052 B.n533 B.n288 65.6433
R1053 B.n540 B.n288 65.6433
R1054 B.n540 B.n539 65.6433
R1055 B.n546 B.n281 65.6433
R1056 B.n552 B.n281 65.6433
R1057 B.n552 B.n277 65.6433
R1058 B.n558 B.n277 65.6433
R1059 B.n558 B.n273 65.6433
R1060 B.n564 B.n273 65.6433
R1061 B.n564 B.n268 65.6433
R1062 B.n570 B.n268 65.6433
R1063 B.n570 B.n269 65.6433
R1064 B.n576 B.n261 65.6433
R1065 B.n582 B.n261 65.6433
R1066 B.n582 B.n257 65.6433
R1067 B.n588 B.n257 65.6433
R1068 B.n588 B.n253 65.6433
R1069 B.n594 B.n253 65.6433
R1070 B.n594 B.n249 65.6433
R1071 B.n601 B.n249 65.6433
R1072 B.n601 B.n600 65.6433
R1073 B.n607 B.n242 65.6433
R1074 B.n614 B.n242 65.6433
R1075 B.n614 B.n238 65.6433
R1076 B.n620 B.n238 65.6433
R1077 B.n620 B.n4 65.6433
R1078 B.n785 B.n4 65.6433
R1079 B.n785 B.n784 65.6433
R1080 B.n784 B.n783 65.6433
R1081 B.n783 B.n8 65.6433
R1082 B.n777 B.n8 65.6433
R1083 B.n777 B.n776 65.6433
R1084 B.n776 B.n775 65.6433
R1085 B.n769 B.n18 65.6433
R1086 B.n769 B.n768 65.6433
R1087 B.n768 B.n767 65.6433
R1088 B.n767 B.n22 65.6433
R1089 B.n761 B.n22 65.6433
R1090 B.n761 B.n760 65.6433
R1091 B.n760 B.n759 65.6433
R1092 B.n759 B.n29 65.6433
R1093 B.n753 B.n29 65.6433
R1094 B.n752 B.n751 65.6433
R1095 B.n751 B.n36 65.6433
R1096 B.n745 B.n36 65.6433
R1097 B.n745 B.n744 65.6433
R1098 B.n744 B.n743 65.6433
R1099 B.n743 B.n43 65.6433
R1100 B.n737 B.n43 65.6433
R1101 B.n737 B.n736 65.6433
R1102 B.n736 B.n735 65.6433
R1103 B.n729 B.n53 65.6433
R1104 B.n729 B.n728 65.6433
R1105 B.n728 B.n727 65.6433
R1106 B.n727 B.n57 65.6433
R1107 B.n721 B.n57 65.6433
R1108 B.n721 B.n720 65.6433
R1109 B.n720 B.n719 65.6433
R1110 B.n719 B.n64 65.6433
R1111 B.n713 B.n64 65.6433
R1112 B.n713 B.n712 65.6433
R1113 B.n712 B.n711 65.6433
R1114 B.n711 B.n71 65.6433
R1115 B.n705 B.n704 65.6433
R1116 B.n704 B.n703 65.6433
R1117 B.n703 B.n78 65.6433
R1118 B.n697 B.n78 65.6433
R1119 B.n697 B.n696 65.6433
R1120 B.n696 B.n695 65.6433
R1121 B.n695 B.n85 65.6433
R1122 B.n689 B.n85 65.6433
R1123 B.t11 B.n308 59.8513
R1124 B.t7 B.n71 59.8513
R1125 B.n427 B.n426 59.5399
R1126 B.n407 B.n348 59.5399
R1127 B.n124 B.n123 59.5399
R1128 B.n121 B.n120 59.5399
R1129 B.n546 B.t4 44.4059
R1130 B.n735 B.t0 44.4059
R1131 B.n576 B.t5 42.4753
R1132 B.n753 B.t2 42.4753
R1133 B.n607 B.t1 40.5446
R1134 B.n775 B.t3 40.5446
R1135 B.n685 B.n684 36.059
R1136 B.n691 B.n87 36.059
R1137 B.n477 B.n476 36.059
R1138 B.n481 B.n326 36.059
R1139 B.n600 B.t1 25.0992
R1140 B.n18 B.t3 25.0992
R1141 B.n269 B.t5 23.1686
R1142 B.t2 B.n752 23.1686
R1143 B.n539 B.t4 21.2379
R1144 B.n53 B.t0 21.2379
R1145 B B.n787 18.0485
R1146 B.n125 B.n87 10.6151
R1147 B.n128 B.n125 10.6151
R1148 B.n129 B.n128 10.6151
R1149 B.n132 B.n129 10.6151
R1150 B.n133 B.n132 10.6151
R1151 B.n136 B.n133 10.6151
R1152 B.n137 B.n136 10.6151
R1153 B.n140 B.n137 10.6151
R1154 B.n141 B.n140 10.6151
R1155 B.n144 B.n141 10.6151
R1156 B.n145 B.n144 10.6151
R1157 B.n148 B.n145 10.6151
R1158 B.n149 B.n148 10.6151
R1159 B.n152 B.n149 10.6151
R1160 B.n153 B.n152 10.6151
R1161 B.n156 B.n153 10.6151
R1162 B.n157 B.n156 10.6151
R1163 B.n160 B.n157 10.6151
R1164 B.n161 B.n160 10.6151
R1165 B.n164 B.n161 10.6151
R1166 B.n165 B.n164 10.6151
R1167 B.n168 B.n165 10.6151
R1168 B.n169 B.n168 10.6151
R1169 B.n173 B.n172 10.6151
R1170 B.n176 B.n173 10.6151
R1171 B.n177 B.n176 10.6151
R1172 B.n180 B.n177 10.6151
R1173 B.n181 B.n180 10.6151
R1174 B.n184 B.n181 10.6151
R1175 B.n185 B.n184 10.6151
R1176 B.n188 B.n185 10.6151
R1177 B.n189 B.n188 10.6151
R1178 B.n193 B.n192 10.6151
R1179 B.n196 B.n193 10.6151
R1180 B.n197 B.n196 10.6151
R1181 B.n200 B.n197 10.6151
R1182 B.n201 B.n200 10.6151
R1183 B.n204 B.n201 10.6151
R1184 B.n205 B.n204 10.6151
R1185 B.n208 B.n205 10.6151
R1186 B.n209 B.n208 10.6151
R1187 B.n212 B.n209 10.6151
R1188 B.n213 B.n212 10.6151
R1189 B.n216 B.n213 10.6151
R1190 B.n217 B.n216 10.6151
R1191 B.n220 B.n217 10.6151
R1192 B.n221 B.n220 10.6151
R1193 B.n224 B.n221 10.6151
R1194 B.n225 B.n224 10.6151
R1195 B.n228 B.n225 10.6151
R1196 B.n229 B.n228 10.6151
R1197 B.n232 B.n229 10.6151
R1198 B.n234 B.n232 10.6151
R1199 B.n235 B.n234 10.6151
R1200 B.n685 B.n235 10.6151
R1201 B.n477 B.n322 10.6151
R1202 B.n487 B.n322 10.6151
R1203 B.n488 B.n487 10.6151
R1204 B.n489 B.n488 10.6151
R1205 B.n489 B.n314 10.6151
R1206 B.n499 B.n314 10.6151
R1207 B.n500 B.n499 10.6151
R1208 B.n501 B.n500 10.6151
R1209 B.n501 B.n306 10.6151
R1210 B.n511 B.n306 10.6151
R1211 B.n512 B.n511 10.6151
R1212 B.n513 B.n512 10.6151
R1213 B.n513 B.n298 10.6151
R1214 B.n523 B.n298 10.6151
R1215 B.n524 B.n523 10.6151
R1216 B.n525 B.n524 10.6151
R1217 B.n525 B.n290 10.6151
R1218 B.n535 B.n290 10.6151
R1219 B.n536 B.n535 10.6151
R1220 B.n537 B.n536 10.6151
R1221 B.n537 B.n283 10.6151
R1222 B.n548 B.n283 10.6151
R1223 B.n549 B.n548 10.6151
R1224 B.n550 B.n549 10.6151
R1225 B.n550 B.n275 10.6151
R1226 B.n560 B.n275 10.6151
R1227 B.n561 B.n560 10.6151
R1228 B.n562 B.n561 10.6151
R1229 B.n562 B.n266 10.6151
R1230 B.n572 B.n266 10.6151
R1231 B.n573 B.n572 10.6151
R1232 B.n574 B.n573 10.6151
R1233 B.n574 B.n259 10.6151
R1234 B.n584 B.n259 10.6151
R1235 B.n585 B.n584 10.6151
R1236 B.n586 B.n585 10.6151
R1237 B.n586 B.n251 10.6151
R1238 B.n596 B.n251 10.6151
R1239 B.n597 B.n596 10.6151
R1240 B.n598 B.n597 10.6151
R1241 B.n598 B.n244 10.6151
R1242 B.n609 B.n244 10.6151
R1243 B.n610 B.n609 10.6151
R1244 B.n612 B.n610 10.6151
R1245 B.n612 B.n611 10.6151
R1246 B.n611 B.n236 10.6151
R1247 B.n623 B.n236 10.6151
R1248 B.n624 B.n623 10.6151
R1249 B.n625 B.n624 10.6151
R1250 B.n626 B.n625 10.6151
R1251 B.n628 B.n626 10.6151
R1252 B.n629 B.n628 10.6151
R1253 B.n630 B.n629 10.6151
R1254 B.n631 B.n630 10.6151
R1255 B.n633 B.n631 10.6151
R1256 B.n634 B.n633 10.6151
R1257 B.n635 B.n634 10.6151
R1258 B.n636 B.n635 10.6151
R1259 B.n638 B.n636 10.6151
R1260 B.n639 B.n638 10.6151
R1261 B.n640 B.n639 10.6151
R1262 B.n641 B.n640 10.6151
R1263 B.n643 B.n641 10.6151
R1264 B.n644 B.n643 10.6151
R1265 B.n645 B.n644 10.6151
R1266 B.n646 B.n645 10.6151
R1267 B.n648 B.n646 10.6151
R1268 B.n649 B.n648 10.6151
R1269 B.n650 B.n649 10.6151
R1270 B.n651 B.n650 10.6151
R1271 B.n653 B.n651 10.6151
R1272 B.n654 B.n653 10.6151
R1273 B.n655 B.n654 10.6151
R1274 B.n656 B.n655 10.6151
R1275 B.n658 B.n656 10.6151
R1276 B.n659 B.n658 10.6151
R1277 B.n660 B.n659 10.6151
R1278 B.n661 B.n660 10.6151
R1279 B.n663 B.n661 10.6151
R1280 B.n664 B.n663 10.6151
R1281 B.n665 B.n664 10.6151
R1282 B.n666 B.n665 10.6151
R1283 B.n668 B.n666 10.6151
R1284 B.n669 B.n668 10.6151
R1285 B.n670 B.n669 10.6151
R1286 B.n671 B.n670 10.6151
R1287 B.n673 B.n671 10.6151
R1288 B.n674 B.n673 10.6151
R1289 B.n675 B.n674 10.6151
R1290 B.n676 B.n675 10.6151
R1291 B.n678 B.n676 10.6151
R1292 B.n679 B.n678 10.6151
R1293 B.n680 B.n679 10.6151
R1294 B.n681 B.n680 10.6151
R1295 B.n683 B.n681 10.6151
R1296 B.n684 B.n683 10.6151
R1297 B.n360 B.n326 10.6151
R1298 B.n360 B.n359 10.6151
R1299 B.n366 B.n359 10.6151
R1300 B.n367 B.n366 10.6151
R1301 B.n368 B.n367 10.6151
R1302 B.n368 B.n357 10.6151
R1303 B.n374 B.n357 10.6151
R1304 B.n375 B.n374 10.6151
R1305 B.n376 B.n375 10.6151
R1306 B.n376 B.n355 10.6151
R1307 B.n382 B.n355 10.6151
R1308 B.n383 B.n382 10.6151
R1309 B.n384 B.n383 10.6151
R1310 B.n384 B.n353 10.6151
R1311 B.n390 B.n353 10.6151
R1312 B.n391 B.n390 10.6151
R1313 B.n392 B.n391 10.6151
R1314 B.n392 B.n351 10.6151
R1315 B.n398 B.n351 10.6151
R1316 B.n399 B.n398 10.6151
R1317 B.n400 B.n399 10.6151
R1318 B.n400 B.n349 10.6151
R1319 B.n406 B.n349 10.6151
R1320 B.n409 B.n408 10.6151
R1321 B.n409 B.n345 10.6151
R1322 B.n415 B.n345 10.6151
R1323 B.n416 B.n415 10.6151
R1324 B.n417 B.n416 10.6151
R1325 B.n417 B.n343 10.6151
R1326 B.n423 B.n343 10.6151
R1327 B.n424 B.n423 10.6151
R1328 B.n428 B.n424 10.6151
R1329 B.n434 B.n341 10.6151
R1330 B.n435 B.n434 10.6151
R1331 B.n436 B.n435 10.6151
R1332 B.n436 B.n339 10.6151
R1333 B.n442 B.n339 10.6151
R1334 B.n443 B.n442 10.6151
R1335 B.n444 B.n443 10.6151
R1336 B.n444 B.n337 10.6151
R1337 B.n450 B.n337 10.6151
R1338 B.n451 B.n450 10.6151
R1339 B.n452 B.n451 10.6151
R1340 B.n452 B.n335 10.6151
R1341 B.n458 B.n335 10.6151
R1342 B.n459 B.n458 10.6151
R1343 B.n460 B.n459 10.6151
R1344 B.n460 B.n333 10.6151
R1345 B.n466 B.n333 10.6151
R1346 B.n467 B.n466 10.6151
R1347 B.n468 B.n467 10.6151
R1348 B.n468 B.n331 10.6151
R1349 B.n331 B.n330 10.6151
R1350 B.n475 B.n330 10.6151
R1351 B.n476 B.n475 10.6151
R1352 B.n482 B.n481 10.6151
R1353 B.n483 B.n482 10.6151
R1354 B.n483 B.n318 10.6151
R1355 B.n493 B.n318 10.6151
R1356 B.n494 B.n493 10.6151
R1357 B.n495 B.n494 10.6151
R1358 B.n495 B.n310 10.6151
R1359 B.n505 B.n310 10.6151
R1360 B.n506 B.n505 10.6151
R1361 B.n507 B.n506 10.6151
R1362 B.n507 B.n302 10.6151
R1363 B.n517 B.n302 10.6151
R1364 B.n518 B.n517 10.6151
R1365 B.n519 B.n518 10.6151
R1366 B.n519 B.n294 10.6151
R1367 B.n529 B.n294 10.6151
R1368 B.n530 B.n529 10.6151
R1369 B.n531 B.n530 10.6151
R1370 B.n531 B.n286 10.6151
R1371 B.n542 B.n286 10.6151
R1372 B.n543 B.n542 10.6151
R1373 B.n544 B.n543 10.6151
R1374 B.n544 B.n279 10.6151
R1375 B.n554 B.n279 10.6151
R1376 B.n555 B.n554 10.6151
R1377 B.n556 B.n555 10.6151
R1378 B.n556 B.n271 10.6151
R1379 B.n566 B.n271 10.6151
R1380 B.n567 B.n566 10.6151
R1381 B.n568 B.n567 10.6151
R1382 B.n568 B.n263 10.6151
R1383 B.n578 B.n263 10.6151
R1384 B.n579 B.n578 10.6151
R1385 B.n580 B.n579 10.6151
R1386 B.n580 B.n255 10.6151
R1387 B.n590 B.n255 10.6151
R1388 B.n591 B.n590 10.6151
R1389 B.n592 B.n591 10.6151
R1390 B.n592 B.n247 10.6151
R1391 B.n603 B.n247 10.6151
R1392 B.n604 B.n603 10.6151
R1393 B.n605 B.n604 10.6151
R1394 B.n605 B.n240 10.6151
R1395 B.n616 B.n240 10.6151
R1396 B.n617 B.n616 10.6151
R1397 B.n618 B.n617 10.6151
R1398 B.n618 B.n0 10.6151
R1399 B.n781 B.n1 10.6151
R1400 B.n781 B.n780 10.6151
R1401 B.n780 B.n779 10.6151
R1402 B.n779 B.n10 10.6151
R1403 B.n773 B.n10 10.6151
R1404 B.n773 B.n772 10.6151
R1405 B.n772 B.n771 10.6151
R1406 B.n771 B.n16 10.6151
R1407 B.n765 B.n16 10.6151
R1408 B.n765 B.n764 10.6151
R1409 B.n764 B.n763 10.6151
R1410 B.n763 B.n24 10.6151
R1411 B.n757 B.n24 10.6151
R1412 B.n757 B.n756 10.6151
R1413 B.n756 B.n755 10.6151
R1414 B.n755 B.n31 10.6151
R1415 B.n749 B.n31 10.6151
R1416 B.n749 B.n748 10.6151
R1417 B.n748 B.n747 10.6151
R1418 B.n747 B.n38 10.6151
R1419 B.n741 B.n38 10.6151
R1420 B.n741 B.n740 10.6151
R1421 B.n740 B.n739 10.6151
R1422 B.n739 B.n45 10.6151
R1423 B.n733 B.n45 10.6151
R1424 B.n733 B.n732 10.6151
R1425 B.n732 B.n731 10.6151
R1426 B.n731 B.n51 10.6151
R1427 B.n725 B.n51 10.6151
R1428 B.n725 B.n724 10.6151
R1429 B.n724 B.n723 10.6151
R1430 B.n723 B.n59 10.6151
R1431 B.n717 B.n59 10.6151
R1432 B.n717 B.n716 10.6151
R1433 B.n716 B.n715 10.6151
R1434 B.n715 B.n66 10.6151
R1435 B.n709 B.n66 10.6151
R1436 B.n709 B.n708 10.6151
R1437 B.n708 B.n707 10.6151
R1438 B.n707 B.n73 10.6151
R1439 B.n701 B.n73 10.6151
R1440 B.n701 B.n700 10.6151
R1441 B.n700 B.n699 10.6151
R1442 B.n699 B.n80 10.6151
R1443 B.n693 B.n80 10.6151
R1444 B.n693 B.n692 10.6151
R1445 B.n692 B.n691 10.6151
R1446 B.n169 B.n124 9.36635
R1447 B.n192 B.n121 9.36635
R1448 B.n407 B.n406 9.36635
R1449 B.n427 B.n341 9.36635
R1450 B.n503 B.t11 5.79251
R1451 B.n705 B.t7 5.79251
R1452 B.n787 B.n0 2.81026
R1453 B.n787 B.n1 2.81026
R1454 B.n172 B.n124 1.24928
R1455 B.n189 B.n121 1.24928
R1456 B.n408 B.n407 1.24928
R1457 B.n428 B.n427 1.24928
R1458 VP.n13 VP.n10 161.3
R1459 VP.n15 VP.n14 161.3
R1460 VP.n16 VP.n9 161.3
R1461 VP.n18 VP.n17 161.3
R1462 VP.n19 VP.n8 161.3
R1463 VP.n21 VP.n20 161.3
R1464 VP.n44 VP.n43 161.3
R1465 VP.n42 VP.n1 161.3
R1466 VP.n41 VP.n40 161.3
R1467 VP.n39 VP.n2 161.3
R1468 VP.n38 VP.n37 161.3
R1469 VP.n36 VP.n3 161.3
R1470 VP.n35 VP.n34 161.3
R1471 VP.n33 VP.n4 161.3
R1472 VP.n32 VP.n31 161.3
R1473 VP.n30 VP.n5 161.3
R1474 VP.n29 VP.n28 161.3
R1475 VP.n27 VP.n6 161.3
R1476 VP.n26 VP.n25 161.3
R1477 VP.n11 VP.t2 81.3679
R1478 VP.n24 VP.n23 70.0803
R1479 VP.n45 VP.n0 70.0803
R1480 VP.n22 VP.n7 70.0803
R1481 VP.n30 VP.n29 56.5617
R1482 VP.n41 VP.n2 56.5617
R1483 VP.n18 VP.n9 56.5617
R1484 VP.n12 VP.n11 49.5116
R1485 VP.n35 VP.t3 47.8875
R1486 VP.n24 VP.t4 47.8875
R1487 VP.n0 VP.t1 47.8875
R1488 VP.n12 VP.t0 47.8875
R1489 VP.n7 VP.t5 47.8875
R1490 VP.n23 VP.n22 46.2458
R1491 VP.n25 VP.n6 24.5923
R1492 VP.n29 VP.n6 24.5923
R1493 VP.n31 VP.n30 24.5923
R1494 VP.n31 VP.n4 24.5923
R1495 VP.n35 VP.n4 24.5923
R1496 VP.n36 VP.n35 24.5923
R1497 VP.n37 VP.n36 24.5923
R1498 VP.n37 VP.n2 24.5923
R1499 VP.n42 VP.n41 24.5923
R1500 VP.n43 VP.n42 24.5923
R1501 VP.n19 VP.n18 24.5923
R1502 VP.n20 VP.n19 24.5923
R1503 VP.n13 VP.n12 24.5923
R1504 VP.n14 VP.n13 24.5923
R1505 VP.n14 VP.n9 24.5923
R1506 VP.n25 VP.n24 20.1658
R1507 VP.n43 VP.n0 20.1658
R1508 VP.n20 VP.n7 20.1658
R1509 VP.n11 VP.n10 3.89684
R1510 VP.n22 VP.n21 0.354861
R1511 VP.n26 VP.n23 0.354861
R1512 VP.n45 VP.n44 0.354861
R1513 VP VP.n45 0.267071
R1514 VP.n15 VP.n10 0.189894
R1515 VP.n16 VP.n15 0.189894
R1516 VP.n17 VP.n16 0.189894
R1517 VP.n17 VP.n8 0.189894
R1518 VP.n21 VP.n8 0.189894
R1519 VP.n27 VP.n26 0.189894
R1520 VP.n28 VP.n27 0.189894
R1521 VP.n28 VP.n5 0.189894
R1522 VP.n32 VP.n5 0.189894
R1523 VP.n33 VP.n32 0.189894
R1524 VP.n34 VP.n33 0.189894
R1525 VP.n34 VP.n3 0.189894
R1526 VP.n38 VP.n3 0.189894
R1527 VP.n39 VP.n38 0.189894
R1528 VP.n40 VP.n39 0.189894
R1529 VP.n40 VP.n1 0.189894
R1530 VP.n44 VP.n1 0.189894
R1531 VDD1 VDD1.t3 73.6876
R1532 VDD1.n1 VDD1.t1 73.573
R1533 VDD1.n1 VDD1.n0 68.8688
R1534 VDD1.n3 VDD1.n2 68.1884
R1535 VDD1.n3 VDD1.n1 40.5979
R1536 VDD1.n2 VDD1.t5 3.23579
R1537 VDD1.n2 VDD1.t0 3.23579
R1538 VDD1.n0 VDD1.t2 3.23579
R1539 VDD1.n0 VDD1.t4 3.23579
R1540 VDD1 VDD1.n3 0.677224
C0 VDD1 VN 0.151817f
C1 VN VDD2 3.72593f
C2 VTAIL VP 4.449399f
C3 VDD1 VP 4.07093f
C4 VDD1 VTAIL 5.85031f
C5 VDD2 VP 0.499027f
C6 VTAIL VDD2 5.90597f
C7 VN VP 6.29968f
C8 VTAIL VN 4.43522f
C9 VDD1 VDD2 1.59422f
C10 VDD2 B 5.300449f
C11 VDD1 B 5.650989f
C12 VTAIL B 5.398242f
C13 VN B 13.69681f
C14 VP B 12.392368f
C15 VDD1.t3 B 1.17647f
C16 VDD1.t1 B 1.17565f
C17 VDD1.t2 B 0.108692f
C18 VDD1.t4 B 0.108692f
C19 VDD1.n0 B 0.922342f
C20 VDD1.n1 B 2.56504f
C21 VDD1.t5 B 0.108692f
C22 VDD1.t0 B 0.108692f
C23 VDD1.n2 B 0.917948f
C24 VDD1.n3 B 2.21061f
C25 VP.t1 B 1.21614f
C26 VP.n0 B 0.548964f
C27 VP.n1 B 0.024348f
C28 VP.n2 B 0.032362f
C29 VP.n3 B 0.024348f
C30 VP.t3 B 1.21614f
C31 VP.n4 B 0.045151f
C32 VP.n5 B 0.024348f
C33 VP.n6 B 0.045151f
C34 VP.t5 B 1.21614f
C35 VP.n7 B 0.548964f
C36 VP.n8 B 0.024348f
C37 VP.n9 B 0.032362f
C38 VP.n10 B 0.276941f
C39 VP.t0 B 1.21614f
C40 VP.t2 B 1.47229f
C41 VP.n11 B 0.506243f
C42 VP.n12 B 0.541791f
C43 VP.n13 B 0.045151f
C44 VP.n14 B 0.045151f
C45 VP.n15 B 0.024348f
C46 VP.n16 B 0.024348f
C47 VP.n17 B 0.024348f
C48 VP.n18 B 0.038425f
C49 VP.n19 B 0.045151f
C50 VP.n20 B 0.041139f
C51 VP.n21 B 0.039291f
C52 VP.n22 B 1.22794f
C53 VP.n23 B 1.24692f
C54 VP.t4 B 1.21614f
C55 VP.n24 B 0.548964f
C56 VP.n25 B 0.041139f
C57 VP.n26 B 0.039291f
C58 VP.n27 B 0.024348f
C59 VP.n28 B 0.024348f
C60 VP.n29 B 0.038425f
C61 VP.n30 B 0.032362f
C62 VP.n31 B 0.045151f
C63 VP.n32 B 0.024348f
C64 VP.n33 B 0.024348f
C65 VP.n34 B 0.024348f
C66 VP.n35 B 0.473882f
C67 VP.n36 B 0.045151f
C68 VP.n37 B 0.045151f
C69 VP.n38 B 0.024348f
C70 VP.n39 B 0.024348f
C71 VP.n40 B 0.024348f
C72 VP.n41 B 0.038425f
C73 VP.n42 B 0.045151f
C74 VP.n43 B 0.041139f
C75 VP.n44 B 0.039291f
C76 VP.n45 B 0.051202f
C77 VDD2.t5 B 1.13807f
C78 VDD2.t2 B 0.105218f
C79 VDD2.t4 B 0.105218f
C80 VDD2.n0 B 0.89286f
C81 VDD2.n1 B 2.36919f
C82 VDD2.t3 B 1.12708f
C83 VDD2.n2 B 2.12705f
C84 VDD2.t1 B 0.105218f
C85 VDD2.t0 B 0.105218f
C86 VDD2.n3 B 0.892834f
C87 VTAIL.t6 B 0.133009f
C88 VTAIL.t8 B 0.133009f
C89 VTAIL.n0 B 1.05628f
C90 VTAIL.n1 B 0.484098f
C91 VTAIL.t1 B 1.34304f
C92 VTAIL.n2 B 0.750321f
C93 VTAIL.t4 B 0.133009f
C94 VTAIL.t5 B 0.133009f
C95 VTAIL.n3 B 1.05628f
C96 VTAIL.n4 B 1.8646f
C97 VTAIL.t11 B 0.133009f
C98 VTAIL.t9 B 0.133009f
C99 VTAIL.n5 B 1.05629f
C100 VTAIL.n6 B 1.86459f
C101 VTAIL.t10 B 1.34304f
C102 VTAIL.n7 B 0.750321f
C103 VTAIL.t3 B 0.133009f
C104 VTAIL.t2 B 0.133009f
C105 VTAIL.n8 B 1.05629f
C106 VTAIL.n9 B 0.67432f
C107 VTAIL.t0 B 1.34303f
C108 VTAIL.n10 B 1.68009f
C109 VTAIL.t7 B 1.34304f
C110 VTAIL.n11 B 1.6098f
C111 VN.t1 B 1.18054f
C112 VN.n0 B 0.532894f
C113 VN.n1 B 0.023635f
C114 VN.n2 B 0.031415f
C115 VN.n3 B 0.268834f
C116 VN.t3 B 1.18054f
C117 VN.t0 B 1.42919f
C118 VN.n4 B 0.491423f
C119 VN.n5 B 0.525932f
C120 VN.n6 B 0.043829f
C121 VN.n7 B 0.043829f
C122 VN.n8 B 0.023635f
C123 VN.n9 B 0.023635f
C124 VN.n10 B 0.023635f
C125 VN.n11 B 0.0373f
C126 VN.n12 B 0.043829f
C127 VN.n13 B 0.039935f
C128 VN.n14 B 0.038141f
C129 VN.n15 B 0.049704f
C130 VN.t2 B 1.18054f
C131 VN.n16 B 0.532894f
C132 VN.n17 B 0.023635f
C133 VN.n18 B 0.031415f
C134 VN.n19 B 0.268834f
C135 VN.t4 B 1.18054f
C136 VN.t5 B 1.42919f
C137 VN.n20 B 0.491423f
C138 VN.n21 B 0.525932f
C139 VN.n22 B 0.043829f
C140 VN.n23 B 0.043829f
C141 VN.n24 B 0.023635f
C142 VN.n25 B 0.023635f
C143 VN.n26 B 0.023635f
C144 VN.n27 B 0.0373f
C145 VN.n28 B 0.043829f
C146 VN.n29 B 0.039935f
C147 VN.n30 B 0.038141f
C148 VN.n31 B 1.20194f
.ends

