* NGSPICE file created from diff_pair_sample_0411.ext - technology: sky130A

.subckt diff_pair_sample_0411 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t14 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=2.14
X1 VTAIL.t2 VP.t0 VDD1.t9 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X2 VDD1.t8 VP.t1 VTAIL.t16 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=2.14
X3 B.t11 B.t9 B.t10 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=2.14
X4 B.t8 B.t6 B.t7 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=2.14
X5 VDD2.t8 VN.t1 VTAIL.t7 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=2.14
X6 VTAIL.t12 VN.t2 VDD2.t7 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X7 B.t5 B.t3 B.t4 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=2.14
X8 B.t2 B.t0 B.t1 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=0 ps=0 w=13.23 l=2.14
X9 VTAIL.t19 VP.t2 VDD1.t7 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X10 VTAIL.t9 VN.t3 VDD2.t6 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X11 VTAIL.t15 VP.t3 VDD1.t6 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X12 VDD2.t5 VN.t4 VTAIL.t8 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=2.14
X13 VDD2.t4 VN.t5 VTAIL.t5 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X14 VDD1.t5 VP.t4 VTAIL.t17 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=2.14
X15 VTAIL.t18 VP.t5 VDD1.t4 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X16 VDD1.t3 VP.t6 VTAIL.t4 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X17 VDD2.t3 VN.t6 VTAIL.t6 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=2.14
X18 VDD1.t2 VP.t7 VTAIL.t3 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=5.1597 pd=27.24 as=2.18295 ps=13.56 w=13.23 l=2.14
X19 VDD1.t1 VP.t8 VTAIL.t1 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X20 VTAIL.t11 VN.t7 VDD2.t2 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X21 VTAIL.t10 VN.t8 VDD2.t1 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X22 VDD2.t0 VN.t9 VTAIL.t13 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=2.18295 ps=13.56 w=13.23 l=2.14
X23 VDD1.t0 VP.t9 VTAIL.t0 w_n3934_n3614# sky130_fd_pr__pfet_01v8 ad=2.18295 pd=13.56 as=5.1597 ps=27.24 w=13.23 l=2.14
R0 VN.n8 VN.t0 183.385
R1 VN.n41 VN.t4 183.385
R2 VN.n63 VN.n33 161.3
R3 VN.n62 VN.n61 161.3
R4 VN.n60 VN.n34 161.3
R5 VN.n59 VN.n58 161.3
R6 VN.n57 VN.n35 161.3
R7 VN.n55 VN.n54 161.3
R8 VN.n53 VN.n36 161.3
R9 VN.n52 VN.n51 161.3
R10 VN.n50 VN.n37 161.3
R11 VN.n49 VN.n48 161.3
R12 VN.n47 VN.n38 161.3
R13 VN.n46 VN.n45 161.3
R14 VN.n44 VN.n39 161.3
R15 VN.n43 VN.n42 161.3
R16 VN.n30 VN.n0 161.3
R17 VN.n29 VN.n28 161.3
R18 VN.n27 VN.n1 161.3
R19 VN.n26 VN.n25 161.3
R20 VN.n24 VN.n2 161.3
R21 VN.n22 VN.n21 161.3
R22 VN.n20 VN.n3 161.3
R23 VN.n19 VN.n18 161.3
R24 VN.n17 VN.n4 161.3
R25 VN.n16 VN.n15 161.3
R26 VN.n14 VN.n5 161.3
R27 VN.n13 VN.n12 161.3
R28 VN.n11 VN.n6 161.3
R29 VN.n10 VN.n9 161.3
R30 VN.n16 VN.t9 148.993
R31 VN.n7 VN.t3 148.993
R32 VN.n23 VN.t2 148.993
R33 VN.n31 VN.t6 148.993
R34 VN.n49 VN.t5 148.993
R35 VN.n40 VN.t8 148.993
R36 VN.n56 VN.t7 148.993
R37 VN.n64 VN.t1 148.993
R38 VN.n32 VN.n31 89.2255
R39 VN.n65 VN.n64 89.2255
R40 VN.n12 VN.n11 56.5193
R41 VN.n18 VN.n3 56.5193
R42 VN.n29 VN.n1 56.5193
R43 VN.n45 VN.n44 56.5193
R44 VN.n51 VN.n36 56.5193
R45 VN.n62 VN.n34 56.5193
R46 VN VN.n65 51.911
R47 VN.n8 VN.n7 47.6808
R48 VN.n41 VN.n40 47.6808
R49 VN.n11 VN.n10 24.4675
R50 VN.n12 VN.n5 24.4675
R51 VN.n16 VN.n5 24.4675
R52 VN.n17 VN.n16 24.4675
R53 VN.n18 VN.n17 24.4675
R54 VN.n22 VN.n3 24.4675
R55 VN.n25 VN.n24 24.4675
R56 VN.n25 VN.n1 24.4675
R57 VN.n30 VN.n29 24.4675
R58 VN.n44 VN.n43 24.4675
R59 VN.n51 VN.n50 24.4675
R60 VN.n50 VN.n49 24.4675
R61 VN.n49 VN.n38 24.4675
R62 VN.n45 VN.n38 24.4675
R63 VN.n58 VN.n34 24.4675
R64 VN.n58 VN.n57 24.4675
R65 VN.n55 VN.n36 24.4675
R66 VN.n63 VN.n62 24.4675
R67 VN.n10 VN.n7 22.9995
R68 VN.n23 VN.n22 22.9995
R69 VN.n43 VN.n40 22.9995
R70 VN.n56 VN.n55 22.9995
R71 VN.n31 VN.n30 21.5315
R72 VN.n64 VN.n63 21.5315
R73 VN.n42 VN.n41 8.82758
R74 VN.n9 VN.n8 8.82758
R75 VN.n24 VN.n23 1.46852
R76 VN.n57 VN.n56 1.46852
R77 VN.n65 VN.n33 0.278367
R78 VN.n32 VN.n0 0.278367
R79 VN.n61 VN.n33 0.189894
R80 VN.n61 VN.n60 0.189894
R81 VN.n60 VN.n59 0.189894
R82 VN.n59 VN.n35 0.189894
R83 VN.n54 VN.n35 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n52 0.189894
R86 VN.n52 VN.n37 0.189894
R87 VN.n48 VN.n37 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n46 0.189894
R90 VN.n46 VN.n39 0.189894
R91 VN.n42 VN.n39 0.189894
R92 VN.n9 VN.n6 0.189894
R93 VN.n13 VN.n6 0.189894
R94 VN.n14 VN.n13 0.189894
R95 VN.n15 VN.n14 0.189894
R96 VN.n15 VN.n4 0.189894
R97 VN.n19 VN.n4 0.189894
R98 VN.n20 VN.n19 0.189894
R99 VN.n21 VN.n20 0.189894
R100 VN.n21 VN.n2 0.189894
R101 VN.n26 VN.n2 0.189894
R102 VN.n27 VN.n26 0.189894
R103 VN.n28 VN.n27 0.189894
R104 VN.n28 VN.n0 0.189894
R105 VN VN.n32 0.153454
R106 VTAIL.n11 VTAIL.t8 58.9946
R107 VTAIL.n17 VTAIL.t6 58.9944
R108 VTAIL.n2 VTAIL.t0 58.9944
R109 VTAIL.n16 VTAIL.t17 58.9944
R110 VTAIL.n15 VTAIL.n14 56.5377
R111 VTAIL.n13 VTAIL.n12 56.5377
R112 VTAIL.n10 VTAIL.n9 56.5377
R113 VTAIL.n8 VTAIL.n7 56.5377
R114 VTAIL.n19 VTAIL.n18 56.5377
R115 VTAIL.n1 VTAIL.n0 56.5377
R116 VTAIL.n4 VTAIL.n3 56.5377
R117 VTAIL.n6 VTAIL.n5 56.5377
R118 VTAIL.n8 VTAIL.n6 28.0307
R119 VTAIL.n17 VTAIL.n16 25.9014
R120 VTAIL.n18 VTAIL.t13 2.45742
R121 VTAIL.n18 VTAIL.t12 2.45742
R122 VTAIL.n0 VTAIL.t14 2.45742
R123 VTAIL.n0 VTAIL.t9 2.45742
R124 VTAIL.n3 VTAIL.t4 2.45742
R125 VTAIL.n3 VTAIL.t18 2.45742
R126 VTAIL.n5 VTAIL.t3 2.45742
R127 VTAIL.n5 VTAIL.t19 2.45742
R128 VTAIL.n14 VTAIL.t1 2.45742
R129 VTAIL.n14 VTAIL.t2 2.45742
R130 VTAIL.n12 VTAIL.t16 2.45742
R131 VTAIL.n12 VTAIL.t15 2.45742
R132 VTAIL.n9 VTAIL.t5 2.45742
R133 VTAIL.n9 VTAIL.t10 2.45742
R134 VTAIL.n7 VTAIL.t7 2.45742
R135 VTAIL.n7 VTAIL.t11 2.45742
R136 VTAIL.n10 VTAIL.n8 2.12981
R137 VTAIL.n11 VTAIL.n10 2.12981
R138 VTAIL.n15 VTAIL.n13 2.12981
R139 VTAIL.n16 VTAIL.n15 2.12981
R140 VTAIL.n6 VTAIL.n4 2.12981
R141 VTAIL.n4 VTAIL.n2 2.12981
R142 VTAIL.n19 VTAIL.n17 2.12981
R143 VTAIL VTAIL.n1 1.65567
R144 VTAIL.n13 VTAIL.n11 1.53498
R145 VTAIL.n2 VTAIL.n1 1.53498
R146 VTAIL VTAIL.n19 0.474638
R147 VDD2.n1 VDD2.t9 77.8025
R148 VDD2.n4 VDD2.t8 75.6734
R149 VDD2.n3 VDD2.n2 74.7581
R150 VDD2 VDD2.n7 74.7551
R151 VDD2.n6 VDD2.n5 73.2165
R152 VDD2.n1 VDD2.n0 73.2164
R153 VDD2.n4 VDD2.n3 45.2347
R154 VDD2.n7 VDD2.t1 2.45742
R155 VDD2.n7 VDD2.t5 2.45742
R156 VDD2.n5 VDD2.t2 2.45742
R157 VDD2.n5 VDD2.t4 2.45742
R158 VDD2.n2 VDD2.t7 2.45742
R159 VDD2.n2 VDD2.t3 2.45742
R160 VDD2.n0 VDD2.t6 2.45742
R161 VDD2.n0 VDD2.t0 2.45742
R162 VDD2.n6 VDD2.n4 2.12981
R163 VDD2 VDD2.n6 0.591017
R164 VDD2.n3 VDD2.n1 0.477482
R165 VP.n18 VP.t1 183.385
R166 VP.n20 VP.n19 161.3
R167 VP.n21 VP.n16 161.3
R168 VP.n23 VP.n22 161.3
R169 VP.n24 VP.n15 161.3
R170 VP.n26 VP.n25 161.3
R171 VP.n27 VP.n14 161.3
R172 VP.n29 VP.n28 161.3
R173 VP.n30 VP.n13 161.3
R174 VP.n32 VP.n31 161.3
R175 VP.n34 VP.n12 161.3
R176 VP.n36 VP.n35 161.3
R177 VP.n37 VP.n11 161.3
R178 VP.n39 VP.n38 161.3
R179 VP.n40 VP.n10 161.3
R180 VP.n74 VP.n0 161.3
R181 VP.n73 VP.n72 161.3
R182 VP.n71 VP.n1 161.3
R183 VP.n70 VP.n69 161.3
R184 VP.n68 VP.n2 161.3
R185 VP.n66 VP.n65 161.3
R186 VP.n64 VP.n3 161.3
R187 VP.n63 VP.n62 161.3
R188 VP.n61 VP.n4 161.3
R189 VP.n60 VP.n59 161.3
R190 VP.n58 VP.n5 161.3
R191 VP.n57 VP.n56 161.3
R192 VP.n55 VP.n6 161.3
R193 VP.n54 VP.n53 161.3
R194 VP.n52 VP.n51 161.3
R195 VP.n50 VP.n8 161.3
R196 VP.n49 VP.n48 161.3
R197 VP.n47 VP.n9 161.3
R198 VP.n46 VP.n45 161.3
R199 VP.n60 VP.t6 148.993
R200 VP.n44 VP.t7 148.993
R201 VP.n7 VP.t2 148.993
R202 VP.n67 VP.t5 148.993
R203 VP.n75 VP.t9 148.993
R204 VP.n26 VP.t8 148.993
R205 VP.n41 VP.t4 148.993
R206 VP.n33 VP.t0 148.993
R207 VP.n17 VP.t3 148.993
R208 VP.n44 VP.n43 89.2255
R209 VP.n76 VP.n75 89.2255
R210 VP.n42 VP.n41 89.2255
R211 VP.n49 VP.n9 56.5193
R212 VP.n56 VP.n55 56.5193
R213 VP.n62 VP.n3 56.5193
R214 VP.n73 VP.n1 56.5193
R215 VP.n39 VP.n11 56.5193
R216 VP.n28 VP.n13 56.5193
R217 VP.n22 VP.n21 56.5193
R218 VP.n43 VP.n42 51.6322
R219 VP.n18 VP.n17 47.6808
R220 VP.n45 VP.n9 24.4675
R221 VP.n50 VP.n49 24.4675
R222 VP.n51 VP.n50 24.4675
R223 VP.n55 VP.n54 24.4675
R224 VP.n56 VP.n5 24.4675
R225 VP.n60 VP.n5 24.4675
R226 VP.n61 VP.n60 24.4675
R227 VP.n62 VP.n61 24.4675
R228 VP.n66 VP.n3 24.4675
R229 VP.n69 VP.n68 24.4675
R230 VP.n69 VP.n1 24.4675
R231 VP.n74 VP.n73 24.4675
R232 VP.n40 VP.n39 24.4675
R233 VP.n32 VP.n13 24.4675
R234 VP.n35 VP.n34 24.4675
R235 VP.n35 VP.n11 24.4675
R236 VP.n22 VP.n15 24.4675
R237 VP.n26 VP.n15 24.4675
R238 VP.n27 VP.n26 24.4675
R239 VP.n28 VP.n27 24.4675
R240 VP.n21 VP.n20 24.4675
R241 VP.n54 VP.n7 22.9995
R242 VP.n67 VP.n66 22.9995
R243 VP.n33 VP.n32 22.9995
R244 VP.n20 VP.n17 22.9995
R245 VP.n45 VP.n44 21.5315
R246 VP.n75 VP.n74 21.5315
R247 VP.n41 VP.n40 21.5315
R248 VP.n19 VP.n18 8.82758
R249 VP.n51 VP.n7 1.46852
R250 VP.n68 VP.n67 1.46852
R251 VP.n34 VP.n33 1.46852
R252 VP.n42 VP.n10 0.278367
R253 VP.n46 VP.n43 0.278367
R254 VP.n76 VP.n0 0.278367
R255 VP.n19 VP.n16 0.189894
R256 VP.n23 VP.n16 0.189894
R257 VP.n24 VP.n23 0.189894
R258 VP.n25 VP.n24 0.189894
R259 VP.n25 VP.n14 0.189894
R260 VP.n29 VP.n14 0.189894
R261 VP.n30 VP.n29 0.189894
R262 VP.n31 VP.n30 0.189894
R263 VP.n31 VP.n12 0.189894
R264 VP.n36 VP.n12 0.189894
R265 VP.n37 VP.n36 0.189894
R266 VP.n38 VP.n37 0.189894
R267 VP.n38 VP.n10 0.189894
R268 VP.n47 VP.n46 0.189894
R269 VP.n48 VP.n47 0.189894
R270 VP.n48 VP.n8 0.189894
R271 VP.n52 VP.n8 0.189894
R272 VP.n53 VP.n52 0.189894
R273 VP.n53 VP.n6 0.189894
R274 VP.n57 VP.n6 0.189894
R275 VP.n58 VP.n57 0.189894
R276 VP.n59 VP.n58 0.189894
R277 VP.n59 VP.n4 0.189894
R278 VP.n63 VP.n4 0.189894
R279 VP.n64 VP.n63 0.189894
R280 VP.n65 VP.n64 0.189894
R281 VP.n65 VP.n2 0.189894
R282 VP.n70 VP.n2 0.189894
R283 VP.n71 VP.n70 0.189894
R284 VP.n72 VP.n71 0.189894
R285 VP.n72 VP.n0 0.189894
R286 VP VP.n76 0.153454
R287 VDD1.n1 VDD1.t8 77.8027
R288 VDD1.n3 VDD1.t2 77.8025
R289 VDD1.n5 VDD1.n4 74.7581
R290 VDD1.n1 VDD1.n0 73.2165
R291 VDD1.n3 VDD1.n2 73.2164
R292 VDD1.n7 VDD1.n6 73.2163
R293 VDD1.n7 VDD1.n5 46.8824
R294 VDD1.n6 VDD1.t9 2.45742
R295 VDD1.n6 VDD1.t5 2.45742
R296 VDD1.n0 VDD1.t6 2.45742
R297 VDD1.n0 VDD1.t1 2.45742
R298 VDD1.n4 VDD1.t4 2.45742
R299 VDD1.n4 VDD1.t0 2.45742
R300 VDD1.n2 VDD1.t7 2.45742
R301 VDD1.n2 VDD1.t3 2.45742
R302 VDD1 VDD1.n7 1.53929
R303 VDD1 VDD1.n1 0.591017
R304 VDD1.n5 VDD1.n3 0.477482
R305 B.n439 B.n134 585
R306 B.n438 B.n437 585
R307 B.n436 B.n135 585
R308 B.n435 B.n434 585
R309 B.n433 B.n136 585
R310 B.n432 B.n431 585
R311 B.n430 B.n137 585
R312 B.n429 B.n428 585
R313 B.n427 B.n138 585
R314 B.n426 B.n425 585
R315 B.n424 B.n139 585
R316 B.n423 B.n422 585
R317 B.n421 B.n140 585
R318 B.n420 B.n419 585
R319 B.n418 B.n141 585
R320 B.n417 B.n416 585
R321 B.n415 B.n142 585
R322 B.n414 B.n413 585
R323 B.n412 B.n143 585
R324 B.n411 B.n410 585
R325 B.n409 B.n144 585
R326 B.n408 B.n407 585
R327 B.n406 B.n145 585
R328 B.n405 B.n404 585
R329 B.n403 B.n146 585
R330 B.n402 B.n401 585
R331 B.n400 B.n147 585
R332 B.n399 B.n398 585
R333 B.n397 B.n148 585
R334 B.n396 B.n395 585
R335 B.n394 B.n149 585
R336 B.n393 B.n392 585
R337 B.n391 B.n150 585
R338 B.n390 B.n389 585
R339 B.n388 B.n151 585
R340 B.n387 B.n386 585
R341 B.n385 B.n152 585
R342 B.n384 B.n383 585
R343 B.n382 B.n153 585
R344 B.n381 B.n380 585
R345 B.n379 B.n154 585
R346 B.n378 B.n377 585
R347 B.n376 B.n155 585
R348 B.n375 B.n374 585
R349 B.n373 B.n156 585
R350 B.n372 B.n371 585
R351 B.n367 B.n157 585
R352 B.n366 B.n365 585
R353 B.n364 B.n158 585
R354 B.n363 B.n362 585
R355 B.n361 B.n159 585
R356 B.n360 B.n359 585
R357 B.n358 B.n160 585
R358 B.n357 B.n356 585
R359 B.n355 B.n161 585
R360 B.n353 B.n352 585
R361 B.n351 B.n164 585
R362 B.n350 B.n349 585
R363 B.n348 B.n165 585
R364 B.n347 B.n346 585
R365 B.n345 B.n166 585
R366 B.n344 B.n343 585
R367 B.n342 B.n167 585
R368 B.n341 B.n340 585
R369 B.n339 B.n168 585
R370 B.n338 B.n337 585
R371 B.n336 B.n169 585
R372 B.n335 B.n334 585
R373 B.n333 B.n170 585
R374 B.n332 B.n331 585
R375 B.n330 B.n171 585
R376 B.n329 B.n328 585
R377 B.n327 B.n172 585
R378 B.n326 B.n325 585
R379 B.n324 B.n173 585
R380 B.n323 B.n322 585
R381 B.n321 B.n174 585
R382 B.n320 B.n319 585
R383 B.n318 B.n175 585
R384 B.n317 B.n316 585
R385 B.n315 B.n176 585
R386 B.n314 B.n313 585
R387 B.n312 B.n177 585
R388 B.n311 B.n310 585
R389 B.n309 B.n178 585
R390 B.n308 B.n307 585
R391 B.n306 B.n179 585
R392 B.n305 B.n304 585
R393 B.n303 B.n180 585
R394 B.n302 B.n301 585
R395 B.n300 B.n181 585
R396 B.n299 B.n298 585
R397 B.n297 B.n182 585
R398 B.n296 B.n295 585
R399 B.n294 B.n183 585
R400 B.n293 B.n292 585
R401 B.n291 B.n184 585
R402 B.n290 B.n289 585
R403 B.n288 B.n185 585
R404 B.n287 B.n286 585
R405 B.n441 B.n440 585
R406 B.n442 B.n133 585
R407 B.n444 B.n443 585
R408 B.n445 B.n132 585
R409 B.n447 B.n446 585
R410 B.n448 B.n131 585
R411 B.n450 B.n449 585
R412 B.n451 B.n130 585
R413 B.n453 B.n452 585
R414 B.n454 B.n129 585
R415 B.n456 B.n455 585
R416 B.n457 B.n128 585
R417 B.n459 B.n458 585
R418 B.n460 B.n127 585
R419 B.n462 B.n461 585
R420 B.n463 B.n126 585
R421 B.n465 B.n464 585
R422 B.n466 B.n125 585
R423 B.n468 B.n467 585
R424 B.n469 B.n124 585
R425 B.n471 B.n470 585
R426 B.n472 B.n123 585
R427 B.n474 B.n473 585
R428 B.n475 B.n122 585
R429 B.n477 B.n476 585
R430 B.n478 B.n121 585
R431 B.n480 B.n479 585
R432 B.n481 B.n120 585
R433 B.n483 B.n482 585
R434 B.n484 B.n119 585
R435 B.n486 B.n485 585
R436 B.n487 B.n118 585
R437 B.n489 B.n488 585
R438 B.n490 B.n117 585
R439 B.n492 B.n491 585
R440 B.n493 B.n116 585
R441 B.n495 B.n494 585
R442 B.n496 B.n115 585
R443 B.n498 B.n497 585
R444 B.n499 B.n114 585
R445 B.n501 B.n500 585
R446 B.n502 B.n113 585
R447 B.n504 B.n503 585
R448 B.n505 B.n112 585
R449 B.n507 B.n506 585
R450 B.n508 B.n111 585
R451 B.n510 B.n509 585
R452 B.n511 B.n110 585
R453 B.n513 B.n512 585
R454 B.n514 B.n109 585
R455 B.n516 B.n515 585
R456 B.n517 B.n108 585
R457 B.n519 B.n518 585
R458 B.n520 B.n107 585
R459 B.n522 B.n521 585
R460 B.n523 B.n106 585
R461 B.n525 B.n524 585
R462 B.n526 B.n105 585
R463 B.n528 B.n527 585
R464 B.n529 B.n104 585
R465 B.n531 B.n530 585
R466 B.n532 B.n103 585
R467 B.n534 B.n533 585
R468 B.n535 B.n102 585
R469 B.n537 B.n536 585
R470 B.n538 B.n101 585
R471 B.n540 B.n539 585
R472 B.n541 B.n100 585
R473 B.n543 B.n542 585
R474 B.n544 B.n99 585
R475 B.n546 B.n545 585
R476 B.n547 B.n98 585
R477 B.n549 B.n548 585
R478 B.n550 B.n97 585
R479 B.n552 B.n551 585
R480 B.n553 B.n96 585
R481 B.n555 B.n554 585
R482 B.n556 B.n95 585
R483 B.n558 B.n557 585
R484 B.n559 B.n94 585
R485 B.n561 B.n560 585
R486 B.n562 B.n93 585
R487 B.n564 B.n563 585
R488 B.n565 B.n92 585
R489 B.n567 B.n566 585
R490 B.n568 B.n91 585
R491 B.n570 B.n569 585
R492 B.n571 B.n90 585
R493 B.n573 B.n572 585
R494 B.n574 B.n89 585
R495 B.n576 B.n575 585
R496 B.n577 B.n88 585
R497 B.n579 B.n578 585
R498 B.n580 B.n87 585
R499 B.n582 B.n581 585
R500 B.n583 B.n86 585
R501 B.n585 B.n584 585
R502 B.n586 B.n85 585
R503 B.n588 B.n587 585
R504 B.n589 B.n84 585
R505 B.n591 B.n590 585
R506 B.n592 B.n83 585
R507 B.n594 B.n593 585
R508 B.n595 B.n82 585
R509 B.n747 B.n746 585
R510 B.n745 B.n28 585
R511 B.n744 B.n743 585
R512 B.n742 B.n29 585
R513 B.n741 B.n740 585
R514 B.n739 B.n30 585
R515 B.n738 B.n737 585
R516 B.n736 B.n31 585
R517 B.n735 B.n734 585
R518 B.n733 B.n32 585
R519 B.n732 B.n731 585
R520 B.n730 B.n33 585
R521 B.n729 B.n728 585
R522 B.n727 B.n34 585
R523 B.n726 B.n725 585
R524 B.n724 B.n35 585
R525 B.n723 B.n722 585
R526 B.n721 B.n36 585
R527 B.n720 B.n719 585
R528 B.n718 B.n37 585
R529 B.n717 B.n716 585
R530 B.n715 B.n38 585
R531 B.n714 B.n713 585
R532 B.n712 B.n39 585
R533 B.n711 B.n710 585
R534 B.n709 B.n40 585
R535 B.n708 B.n707 585
R536 B.n706 B.n41 585
R537 B.n705 B.n704 585
R538 B.n703 B.n42 585
R539 B.n702 B.n701 585
R540 B.n700 B.n43 585
R541 B.n699 B.n698 585
R542 B.n697 B.n44 585
R543 B.n696 B.n695 585
R544 B.n694 B.n45 585
R545 B.n693 B.n692 585
R546 B.n691 B.n46 585
R547 B.n690 B.n689 585
R548 B.n688 B.n47 585
R549 B.n687 B.n686 585
R550 B.n685 B.n48 585
R551 B.n684 B.n683 585
R552 B.n682 B.n49 585
R553 B.n681 B.n680 585
R554 B.n679 B.n678 585
R555 B.n677 B.n53 585
R556 B.n676 B.n675 585
R557 B.n674 B.n54 585
R558 B.n673 B.n672 585
R559 B.n671 B.n55 585
R560 B.n670 B.n669 585
R561 B.n668 B.n56 585
R562 B.n667 B.n666 585
R563 B.n665 B.n57 585
R564 B.n663 B.n662 585
R565 B.n661 B.n60 585
R566 B.n660 B.n659 585
R567 B.n658 B.n61 585
R568 B.n657 B.n656 585
R569 B.n655 B.n62 585
R570 B.n654 B.n653 585
R571 B.n652 B.n63 585
R572 B.n651 B.n650 585
R573 B.n649 B.n64 585
R574 B.n648 B.n647 585
R575 B.n646 B.n65 585
R576 B.n645 B.n644 585
R577 B.n643 B.n66 585
R578 B.n642 B.n641 585
R579 B.n640 B.n67 585
R580 B.n639 B.n638 585
R581 B.n637 B.n68 585
R582 B.n636 B.n635 585
R583 B.n634 B.n69 585
R584 B.n633 B.n632 585
R585 B.n631 B.n70 585
R586 B.n630 B.n629 585
R587 B.n628 B.n71 585
R588 B.n627 B.n626 585
R589 B.n625 B.n72 585
R590 B.n624 B.n623 585
R591 B.n622 B.n73 585
R592 B.n621 B.n620 585
R593 B.n619 B.n74 585
R594 B.n618 B.n617 585
R595 B.n616 B.n75 585
R596 B.n615 B.n614 585
R597 B.n613 B.n76 585
R598 B.n612 B.n611 585
R599 B.n610 B.n77 585
R600 B.n609 B.n608 585
R601 B.n607 B.n78 585
R602 B.n606 B.n605 585
R603 B.n604 B.n79 585
R604 B.n603 B.n602 585
R605 B.n601 B.n80 585
R606 B.n600 B.n599 585
R607 B.n598 B.n81 585
R608 B.n597 B.n596 585
R609 B.n748 B.n27 585
R610 B.n750 B.n749 585
R611 B.n751 B.n26 585
R612 B.n753 B.n752 585
R613 B.n754 B.n25 585
R614 B.n756 B.n755 585
R615 B.n757 B.n24 585
R616 B.n759 B.n758 585
R617 B.n760 B.n23 585
R618 B.n762 B.n761 585
R619 B.n763 B.n22 585
R620 B.n765 B.n764 585
R621 B.n766 B.n21 585
R622 B.n768 B.n767 585
R623 B.n769 B.n20 585
R624 B.n771 B.n770 585
R625 B.n772 B.n19 585
R626 B.n774 B.n773 585
R627 B.n775 B.n18 585
R628 B.n777 B.n776 585
R629 B.n778 B.n17 585
R630 B.n780 B.n779 585
R631 B.n781 B.n16 585
R632 B.n783 B.n782 585
R633 B.n784 B.n15 585
R634 B.n786 B.n785 585
R635 B.n787 B.n14 585
R636 B.n789 B.n788 585
R637 B.n790 B.n13 585
R638 B.n792 B.n791 585
R639 B.n793 B.n12 585
R640 B.n795 B.n794 585
R641 B.n796 B.n11 585
R642 B.n798 B.n797 585
R643 B.n799 B.n10 585
R644 B.n801 B.n800 585
R645 B.n802 B.n9 585
R646 B.n804 B.n803 585
R647 B.n805 B.n8 585
R648 B.n807 B.n806 585
R649 B.n808 B.n7 585
R650 B.n810 B.n809 585
R651 B.n811 B.n6 585
R652 B.n813 B.n812 585
R653 B.n814 B.n5 585
R654 B.n816 B.n815 585
R655 B.n817 B.n4 585
R656 B.n819 B.n818 585
R657 B.n820 B.n3 585
R658 B.n822 B.n821 585
R659 B.n823 B.n0 585
R660 B.n2 B.n1 585
R661 B.n212 B.n211 585
R662 B.n213 B.n210 585
R663 B.n215 B.n214 585
R664 B.n216 B.n209 585
R665 B.n218 B.n217 585
R666 B.n219 B.n208 585
R667 B.n221 B.n220 585
R668 B.n222 B.n207 585
R669 B.n224 B.n223 585
R670 B.n225 B.n206 585
R671 B.n227 B.n226 585
R672 B.n228 B.n205 585
R673 B.n230 B.n229 585
R674 B.n231 B.n204 585
R675 B.n233 B.n232 585
R676 B.n234 B.n203 585
R677 B.n236 B.n235 585
R678 B.n237 B.n202 585
R679 B.n239 B.n238 585
R680 B.n240 B.n201 585
R681 B.n242 B.n241 585
R682 B.n243 B.n200 585
R683 B.n245 B.n244 585
R684 B.n246 B.n199 585
R685 B.n248 B.n247 585
R686 B.n249 B.n198 585
R687 B.n251 B.n250 585
R688 B.n252 B.n197 585
R689 B.n254 B.n253 585
R690 B.n255 B.n196 585
R691 B.n257 B.n256 585
R692 B.n258 B.n195 585
R693 B.n260 B.n259 585
R694 B.n261 B.n194 585
R695 B.n263 B.n262 585
R696 B.n264 B.n193 585
R697 B.n266 B.n265 585
R698 B.n267 B.n192 585
R699 B.n269 B.n268 585
R700 B.n270 B.n191 585
R701 B.n272 B.n271 585
R702 B.n273 B.n190 585
R703 B.n275 B.n274 585
R704 B.n276 B.n189 585
R705 B.n278 B.n277 585
R706 B.n279 B.n188 585
R707 B.n281 B.n280 585
R708 B.n282 B.n187 585
R709 B.n284 B.n283 585
R710 B.n285 B.n186 585
R711 B.n286 B.n285 535.745
R712 B.n440 B.n439 535.745
R713 B.n596 B.n595 535.745
R714 B.n746 B.n27 535.745
R715 B.n162 B.t0 356.221
R716 B.n368 B.t3 356.221
R717 B.n58 B.t9 356.221
R718 B.n50 B.t6 356.221
R719 B.n825 B.n824 256.663
R720 B.n824 B.n823 235.042
R721 B.n824 B.n2 235.042
R722 B.n286 B.n185 163.367
R723 B.n290 B.n185 163.367
R724 B.n291 B.n290 163.367
R725 B.n292 B.n291 163.367
R726 B.n292 B.n183 163.367
R727 B.n296 B.n183 163.367
R728 B.n297 B.n296 163.367
R729 B.n298 B.n297 163.367
R730 B.n298 B.n181 163.367
R731 B.n302 B.n181 163.367
R732 B.n303 B.n302 163.367
R733 B.n304 B.n303 163.367
R734 B.n304 B.n179 163.367
R735 B.n308 B.n179 163.367
R736 B.n309 B.n308 163.367
R737 B.n310 B.n309 163.367
R738 B.n310 B.n177 163.367
R739 B.n314 B.n177 163.367
R740 B.n315 B.n314 163.367
R741 B.n316 B.n315 163.367
R742 B.n316 B.n175 163.367
R743 B.n320 B.n175 163.367
R744 B.n321 B.n320 163.367
R745 B.n322 B.n321 163.367
R746 B.n322 B.n173 163.367
R747 B.n326 B.n173 163.367
R748 B.n327 B.n326 163.367
R749 B.n328 B.n327 163.367
R750 B.n328 B.n171 163.367
R751 B.n332 B.n171 163.367
R752 B.n333 B.n332 163.367
R753 B.n334 B.n333 163.367
R754 B.n334 B.n169 163.367
R755 B.n338 B.n169 163.367
R756 B.n339 B.n338 163.367
R757 B.n340 B.n339 163.367
R758 B.n340 B.n167 163.367
R759 B.n344 B.n167 163.367
R760 B.n345 B.n344 163.367
R761 B.n346 B.n345 163.367
R762 B.n346 B.n165 163.367
R763 B.n350 B.n165 163.367
R764 B.n351 B.n350 163.367
R765 B.n352 B.n351 163.367
R766 B.n352 B.n161 163.367
R767 B.n357 B.n161 163.367
R768 B.n358 B.n357 163.367
R769 B.n359 B.n358 163.367
R770 B.n359 B.n159 163.367
R771 B.n363 B.n159 163.367
R772 B.n364 B.n363 163.367
R773 B.n365 B.n364 163.367
R774 B.n365 B.n157 163.367
R775 B.n372 B.n157 163.367
R776 B.n373 B.n372 163.367
R777 B.n374 B.n373 163.367
R778 B.n374 B.n155 163.367
R779 B.n378 B.n155 163.367
R780 B.n379 B.n378 163.367
R781 B.n380 B.n379 163.367
R782 B.n380 B.n153 163.367
R783 B.n384 B.n153 163.367
R784 B.n385 B.n384 163.367
R785 B.n386 B.n385 163.367
R786 B.n386 B.n151 163.367
R787 B.n390 B.n151 163.367
R788 B.n391 B.n390 163.367
R789 B.n392 B.n391 163.367
R790 B.n392 B.n149 163.367
R791 B.n396 B.n149 163.367
R792 B.n397 B.n396 163.367
R793 B.n398 B.n397 163.367
R794 B.n398 B.n147 163.367
R795 B.n402 B.n147 163.367
R796 B.n403 B.n402 163.367
R797 B.n404 B.n403 163.367
R798 B.n404 B.n145 163.367
R799 B.n408 B.n145 163.367
R800 B.n409 B.n408 163.367
R801 B.n410 B.n409 163.367
R802 B.n410 B.n143 163.367
R803 B.n414 B.n143 163.367
R804 B.n415 B.n414 163.367
R805 B.n416 B.n415 163.367
R806 B.n416 B.n141 163.367
R807 B.n420 B.n141 163.367
R808 B.n421 B.n420 163.367
R809 B.n422 B.n421 163.367
R810 B.n422 B.n139 163.367
R811 B.n426 B.n139 163.367
R812 B.n427 B.n426 163.367
R813 B.n428 B.n427 163.367
R814 B.n428 B.n137 163.367
R815 B.n432 B.n137 163.367
R816 B.n433 B.n432 163.367
R817 B.n434 B.n433 163.367
R818 B.n434 B.n135 163.367
R819 B.n438 B.n135 163.367
R820 B.n439 B.n438 163.367
R821 B.n595 B.n594 163.367
R822 B.n594 B.n83 163.367
R823 B.n590 B.n83 163.367
R824 B.n590 B.n589 163.367
R825 B.n589 B.n588 163.367
R826 B.n588 B.n85 163.367
R827 B.n584 B.n85 163.367
R828 B.n584 B.n583 163.367
R829 B.n583 B.n582 163.367
R830 B.n582 B.n87 163.367
R831 B.n578 B.n87 163.367
R832 B.n578 B.n577 163.367
R833 B.n577 B.n576 163.367
R834 B.n576 B.n89 163.367
R835 B.n572 B.n89 163.367
R836 B.n572 B.n571 163.367
R837 B.n571 B.n570 163.367
R838 B.n570 B.n91 163.367
R839 B.n566 B.n91 163.367
R840 B.n566 B.n565 163.367
R841 B.n565 B.n564 163.367
R842 B.n564 B.n93 163.367
R843 B.n560 B.n93 163.367
R844 B.n560 B.n559 163.367
R845 B.n559 B.n558 163.367
R846 B.n558 B.n95 163.367
R847 B.n554 B.n95 163.367
R848 B.n554 B.n553 163.367
R849 B.n553 B.n552 163.367
R850 B.n552 B.n97 163.367
R851 B.n548 B.n97 163.367
R852 B.n548 B.n547 163.367
R853 B.n547 B.n546 163.367
R854 B.n546 B.n99 163.367
R855 B.n542 B.n99 163.367
R856 B.n542 B.n541 163.367
R857 B.n541 B.n540 163.367
R858 B.n540 B.n101 163.367
R859 B.n536 B.n101 163.367
R860 B.n536 B.n535 163.367
R861 B.n535 B.n534 163.367
R862 B.n534 B.n103 163.367
R863 B.n530 B.n103 163.367
R864 B.n530 B.n529 163.367
R865 B.n529 B.n528 163.367
R866 B.n528 B.n105 163.367
R867 B.n524 B.n105 163.367
R868 B.n524 B.n523 163.367
R869 B.n523 B.n522 163.367
R870 B.n522 B.n107 163.367
R871 B.n518 B.n107 163.367
R872 B.n518 B.n517 163.367
R873 B.n517 B.n516 163.367
R874 B.n516 B.n109 163.367
R875 B.n512 B.n109 163.367
R876 B.n512 B.n511 163.367
R877 B.n511 B.n510 163.367
R878 B.n510 B.n111 163.367
R879 B.n506 B.n111 163.367
R880 B.n506 B.n505 163.367
R881 B.n505 B.n504 163.367
R882 B.n504 B.n113 163.367
R883 B.n500 B.n113 163.367
R884 B.n500 B.n499 163.367
R885 B.n499 B.n498 163.367
R886 B.n498 B.n115 163.367
R887 B.n494 B.n115 163.367
R888 B.n494 B.n493 163.367
R889 B.n493 B.n492 163.367
R890 B.n492 B.n117 163.367
R891 B.n488 B.n117 163.367
R892 B.n488 B.n487 163.367
R893 B.n487 B.n486 163.367
R894 B.n486 B.n119 163.367
R895 B.n482 B.n119 163.367
R896 B.n482 B.n481 163.367
R897 B.n481 B.n480 163.367
R898 B.n480 B.n121 163.367
R899 B.n476 B.n121 163.367
R900 B.n476 B.n475 163.367
R901 B.n475 B.n474 163.367
R902 B.n474 B.n123 163.367
R903 B.n470 B.n123 163.367
R904 B.n470 B.n469 163.367
R905 B.n469 B.n468 163.367
R906 B.n468 B.n125 163.367
R907 B.n464 B.n125 163.367
R908 B.n464 B.n463 163.367
R909 B.n463 B.n462 163.367
R910 B.n462 B.n127 163.367
R911 B.n458 B.n127 163.367
R912 B.n458 B.n457 163.367
R913 B.n457 B.n456 163.367
R914 B.n456 B.n129 163.367
R915 B.n452 B.n129 163.367
R916 B.n452 B.n451 163.367
R917 B.n451 B.n450 163.367
R918 B.n450 B.n131 163.367
R919 B.n446 B.n131 163.367
R920 B.n446 B.n445 163.367
R921 B.n445 B.n444 163.367
R922 B.n444 B.n133 163.367
R923 B.n440 B.n133 163.367
R924 B.n746 B.n745 163.367
R925 B.n745 B.n744 163.367
R926 B.n744 B.n29 163.367
R927 B.n740 B.n29 163.367
R928 B.n740 B.n739 163.367
R929 B.n739 B.n738 163.367
R930 B.n738 B.n31 163.367
R931 B.n734 B.n31 163.367
R932 B.n734 B.n733 163.367
R933 B.n733 B.n732 163.367
R934 B.n732 B.n33 163.367
R935 B.n728 B.n33 163.367
R936 B.n728 B.n727 163.367
R937 B.n727 B.n726 163.367
R938 B.n726 B.n35 163.367
R939 B.n722 B.n35 163.367
R940 B.n722 B.n721 163.367
R941 B.n721 B.n720 163.367
R942 B.n720 B.n37 163.367
R943 B.n716 B.n37 163.367
R944 B.n716 B.n715 163.367
R945 B.n715 B.n714 163.367
R946 B.n714 B.n39 163.367
R947 B.n710 B.n39 163.367
R948 B.n710 B.n709 163.367
R949 B.n709 B.n708 163.367
R950 B.n708 B.n41 163.367
R951 B.n704 B.n41 163.367
R952 B.n704 B.n703 163.367
R953 B.n703 B.n702 163.367
R954 B.n702 B.n43 163.367
R955 B.n698 B.n43 163.367
R956 B.n698 B.n697 163.367
R957 B.n697 B.n696 163.367
R958 B.n696 B.n45 163.367
R959 B.n692 B.n45 163.367
R960 B.n692 B.n691 163.367
R961 B.n691 B.n690 163.367
R962 B.n690 B.n47 163.367
R963 B.n686 B.n47 163.367
R964 B.n686 B.n685 163.367
R965 B.n685 B.n684 163.367
R966 B.n684 B.n49 163.367
R967 B.n680 B.n49 163.367
R968 B.n680 B.n679 163.367
R969 B.n679 B.n53 163.367
R970 B.n675 B.n53 163.367
R971 B.n675 B.n674 163.367
R972 B.n674 B.n673 163.367
R973 B.n673 B.n55 163.367
R974 B.n669 B.n55 163.367
R975 B.n669 B.n668 163.367
R976 B.n668 B.n667 163.367
R977 B.n667 B.n57 163.367
R978 B.n662 B.n57 163.367
R979 B.n662 B.n661 163.367
R980 B.n661 B.n660 163.367
R981 B.n660 B.n61 163.367
R982 B.n656 B.n61 163.367
R983 B.n656 B.n655 163.367
R984 B.n655 B.n654 163.367
R985 B.n654 B.n63 163.367
R986 B.n650 B.n63 163.367
R987 B.n650 B.n649 163.367
R988 B.n649 B.n648 163.367
R989 B.n648 B.n65 163.367
R990 B.n644 B.n65 163.367
R991 B.n644 B.n643 163.367
R992 B.n643 B.n642 163.367
R993 B.n642 B.n67 163.367
R994 B.n638 B.n67 163.367
R995 B.n638 B.n637 163.367
R996 B.n637 B.n636 163.367
R997 B.n636 B.n69 163.367
R998 B.n632 B.n69 163.367
R999 B.n632 B.n631 163.367
R1000 B.n631 B.n630 163.367
R1001 B.n630 B.n71 163.367
R1002 B.n626 B.n71 163.367
R1003 B.n626 B.n625 163.367
R1004 B.n625 B.n624 163.367
R1005 B.n624 B.n73 163.367
R1006 B.n620 B.n73 163.367
R1007 B.n620 B.n619 163.367
R1008 B.n619 B.n618 163.367
R1009 B.n618 B.n75 163.367
R1010 B.n614 B.n75 163.367
R1011 B.n614 B.n613 163.367
R1012 B.n613 B.n612 163.367
R1013 B.n612 B.n77 163.367
R1014 B.n608 B.n77 163.367
R1015 B.n608 B.n607 163.367
R1016 B.n607 B.n606 163.367
R1017 B.n606 B.n79 163.367
R1018 B.n602 B.n79 163.367
R1019 B.n602 B.n601 163.367
R1020 B.n601 B.n600 163.367
R1021 B.n600 B.n81 163.367
R1022 B.n596 B.n81 163.367
R1023 B.n750 B.n27 163.367
R1024 B.n751 B.n750 163.367
R1025 B.n752 B.n751 163.367
R1026 B.n752 B.n25 163.367
R1027 B.n756 B.n25 163.367
R1028 B.n757 B.n756 163.367
R1029 B.n758 B.n757 163.367
R1030 B.n758 B.n23 163.367
R1031 B.n762 B.n23 163.367
R1032 B.n763 B.n762 163.367
R1033 B.n764 B.n763 163.367
R1034 B.n764 B.n21 163.367
R1035 B.n768 B.n21 163.367
R1036 B.n769 B.n768 163.367
R1037 B.n770 B.n769 163.367
R1038 B.n770 B.n19 163.367
R1039 B.n774 B.n19 163.367
R1040 B.n775 B.n774 163.367
R1041 B.n776 B.n775 163.367
R1042 B.n776 B.n17 163.367
R1043 B.n780 B.n17 163.367
R1044 B.n781 B.n780 163.367
R1045 B.n782 B.n781 163.367
R1046 B.n782 B.n15 163.367
R1047 B.n786 B.n15 163.367
R1048 B.n787 B.n786 163.367
R1049 B.n788 B.n787 163.367
R1050 B.n788 B.n13 163.367
R1051 B.n792 B.n13 163.367
R1052 B.n793 B.n792 163.367
R1053 B.n794 B.n793 163.367
R1054 B.n794 B.n11 163.367
R1055 B.n798 B.n11 163.367
R1056 B.n799 B.n798 163.367
R1057 B.n800 B.n799 163.367
R1058 B.n800 B.n9 163.367
R1059 B.n804 B.n9 163.367
R1060 B.n805 B.n804 163.367
R1061 B.n806 B.n805 163.367
R1062 B.n806 B.n7 163.367
R1063 B.n810 B.n7 163.367
R1064 B.n811 B.n810 163.367
R1065 B.n812 B.n811 163.367
R1066 B.n812 B.n5 163.367
R1067 B.n816 B.n5 163.367
R1068 B.n817 B.n816 163.367
R1069 B.n818 B.n817 163.367
R1070 B.n818 B.n3 163.367
R1071 B.n822 B.n3 163.367
R1072 B.n823 B.n822 163.367
R1073 B.n212 B.n2 163.367
R1074 B.n213 B.n212 163.367
R1075 B.n214 B.n213 163.367
R1076 B.n214 B.n209 163.367
R1077 B.n218 B.n209 163.367
R1078 B.n219 B.n218 163.367
R1079 B.n220 B.n219 163.367
R1080 B.n220 B.n207 163.367
R1081 B.n224 B.n207 163.367
R1082 B.n225 B.n224 163.367
R1083 B.n226 B.n225 163.367
R1084 B.n226 B.n205 163.367
R1085 B.n230 B.n205 163.367
R1086 B.n231 B.n230 163.367
R1087 B.n232 B.n231 163.367
R1088 B.n232 B.n203 163.367
R1089 B.n236 B.n203 163.367
R1090 B.n237 B.n236 163.367
R1091 B.n238 B.n237 163.367
R1092 B.n238 B.n201 163.367
R1093 B.n242 B.n201 163.367
R1094 B.n243 B.n242 163.367
R1095 B.n244 B.n243 163.367
R1096 B.n244 B.n199 163.367
R1097 B.n248 B.n199 163.367
R1098 B.n249 B.n248 163.367
R1099 B.n250 B.n249 163.367
R1100 B.n250 B.n197 163.367
R1101 B.n254 B.n197 163.367
R1102 B.n255 B.n254 163.367
R1103 B.n256 B.n255 163.367
R1104 B.n256 B.n195 163.367
R1105 B.n260 B.n195 163.367
R1106 B.n261 B.n260 163.367
R1107 B.n262 B.n261 163.367
R1108 B.n262 B.n193 163.367
R1109 B.n266 B.n193 163.367
R1110 B.n267 B.n266 163.367
R1111 B.n268 B.n267 163.367
R1112 B.n268 B.n191 163.367
R1113 B.n272 B.n191 163.367
R1114 B.n273 B.n272 163.367
R1115 B.n274 B.n273 163.367
R1116 B.n274 B.n189 163.367
R1117 B.n278 B.n189 163.367
R1118 B.n279 B.n278 163.367
R1119 B.n280 B.n279 163.367
R1120 B.n280 B.n187 163.367
R1121 B.n284 B.n187 163.367
R1122 B.n285 B.n284 163.367
R1123 B.n368 B.t4 160.766
R1124 B.n58 B.t11 160.766
R1125 B.n162 B.t1 160.75
R1126 B.n50 B.t8 160.75
R1127 B.n369 B.t5 112.862
R1128 B.n59 B.t10 112.862
R1129 B.n163 B.t2 112.847
R1130 B.n51 B.t7 112.847
R1131 B.n354 B.n163 59.5399
R1132 B.n370 B.n369 59.5399
R1133 B.n664 B.n59 59.5399
R1134 B.n52 B.n51 59.5399
R1135 B.n163 B.n162 47.9035
R1136 B.n369 B.n368 47.9035
R1137 B.n59 B.n58 47.9035
R1138 B.n51 B.n50 47.9035
R1139 B.n748 B.n747 34.8103
R1140 B.n597 B.n82 34.8103
R1141 B.n441 B.n134 34.8103
R1142 B.n287 B.n186 34.8103
R1143 B B.n825 18.0485
R1144 B.n749 B.n748 10.6151
R1145 B.n749 B.n26 10.6151
R1146 B.n753 B.n26 10.6151
R1147 B.n754 B.n753 10.6151
R1148 B.n755 B.n754 10.6151
R1149 B.n755 B.n24 10.6151
R1150 B.n759 B.n24 10.6151
R1151 B.n760 B.n759 10.6151
R1152 B.n761 B.n760 10.6151
R1153 B.n761 B.n22 10.6151
R1154 B.n765 B.n22 10.6151
R1155 B.n766 B.n765 10.6151
R1156 B.n767 B.n766 10.6151
R1157 B.n767 B.n20 10.6151
R1158 B.n771 B.n20 10.6151
R1159 B.n772 B.n771 10.6151
R1160 B.n773 B.n772 10.6151
R1161 B.n773 B.n18 10.6151
R1162 B.n777 B.n18 10.6151
R1163 B.n778 B.n777 10.6151
R1164 B.n779 B.n778 10.6151
R1165 B.n779 B.n16 10.6151
R1166 B.n783 B.n16 10.6151
R1167 B.n784 B.n783 10.6151
R1168 B.n785 B.n784 10.6151
R1169 B.n785 B.n14 10.6151
R1170 B.n789 B.n14 10.6151
R1171 B.n790 B.n789 10.6151
R1172 B.n791 B.n790 10.6151
R1173 B.n791 B.n12 10.6151
R1174 B.n795 B.n12 10.6151
R1175 B.n796 B.n795 10.6151
R1176 B.n797 B.n796 10.6151
R1177 B.n797 B.n10 10.6151
R1178 B.n801 B.n10 10.6151
R1179 B.n802 B.n801 10.6151
R1180 B.n803 B.n802 10.6151
R1181 B.n803 B.n8 10.6151
R1182 B.n807 B.n8 10.6151
R1183 B.n808 B.n807 10.6151
R1184 B.n809 B.n808 10.6151
R1185 B.n809 B.n6 10.6151
R1186 B.n813 B.n6 10.6151
R1187 B.n814 B.n813 10.6151
R1188 B.n815 B.n814 10.6151
R1189 B.n815 B.n4 10.6151
R1190 B.n819 B.n4 10.6151
R1191 B.n820 B.n819 10.6151
R1192 B.n821 B.n820 10.6151
R1193 B.n821 B.n0 10.6151
R1194 B.n747 B.n28 10.6151
R1195 B.n743 B.n28 10.6151
R1196 B.n743 B.n742 10.6151
R1197 B.n742 B.n741 10.6151
R1198 B.n741 B.n30 10.6151
R1199 B.n737 B.n30 10.6151
R1200 B.n737 B.n736 10.6151
R1201 B.n736 B.n735 10.6151
R1202 B.n735 B.n32 10.6151
R1203 B.n731 B.n32 10.6151
R1204 B.n731 B.n730 10.6151
R1205 B.n730 B.n729 10.6151
R1206 B.n729 B.n34 10.6151
R1207 B.n725 B.n34 10.6151
R1208 B.n725 B.n724 10.6151
R1209 B.n724 B.n723 10.6151
R1210 B.n723 B.n36 10.6151
R1211 B.n719 B.n36 10.6151
R1212 B.n719 B.n718 10.6151
R1213 B.n718 B.n717 10.6151
R1214 B.n717 B.n38 10.6151
R1215 B.n713 B.n38 10.6151
R1216 B.n713 B.n712 10.6151
R1217 B.n712 B.n711 10.6151
R1218 B.n711 B.n40 10.6151
R1219 B.n707 B.n40 10.6151
R1220 B.n707 B.n706 10.6151
R1221 B.n706 B.n705 10.6151
R1222 B.n705 B.n42 10.6151
R1223 B.n701 B.n42 10.6151
R1224 B.n701 B.n700 10.6151
R1225 B.n700 B.n699 10.6151
R1226 B.n699 B.n44 10.6151
R1227 B.n695 B.n44 10.6151
R1228 B.n695 B.n694 10.6151
R1229 B.n694 B.n693 10.6151
R1230 B.n693 B.n46 10.6151
R1231 B.n689 B.n46 10.6151
R1232 B.n689 B.n688 10.6151
R1233 B.n688 B.n687 10.6151
R1234 B.n687 B.n48 10.6151
R1235 B.n683 B.n48 10.6151
R1236 B.n683 B.n682 10.6151
R1237 B.n682 B.n681 10.6151
R1238 B.n678 B.n677 10.6151
R1239 B.n677 B.n676 10.6151
R1240 B.n676 B.n54 10.6151
R1241 B.n672 B.n54 10.6151
R1242 B.n672 B.n671 10.6151
R1243 B.n671 B.n670 10.6151
R1244 B.n670 B.n56 10.6151
R1245 B.n666 B.n56 10.6151
R1246 B.n666 B.n665 10.6151
R1247 B.n663 B.n60 10.6151
R1248 B.n659 B.n60 10.6151
R1249 B.n659 B.n658 10.6151
R1250 B.n658 B.n657 10.6151
R1251 B.n657 B.n62 10.6151
R1252 B.n653 B.n62 10.6151
R1253 B.n653 B.n652 10.6151
R1254 B.n652 B.n651 10.6151
R1255 B.n651 B.n64 10.6151
R1256 B.n647 B.n64 10.6151
R1257 B.n647 B.n646 10.6151
R1258 B.n646 B.n645 10.6151
R1259 B.n645 B.n66 10.6151
R1260 B.n641 B.n66 10.6151
R1261 B.n641 B.n640 10.6151
R1262 B.n640 B.n639 10.6151
R1263 B.n639 B.n68 10.6151
R1264 B.n635 B.n68 10.6151
R1265 B.n635 B.n634 10.6151
R1266 B.n634 B.n633 10.6151
R1267 B.n633 B.n70 10.6151
R1268 B.n629 B.n70 10.6151
R1269 B.n629 B.n628 10.6151
R1270 B.n628 B.n627 10.6151
R1271 B.n627 B.n72 10.6151
R1272 B.n623 B.n72 10.6151
R1273 B.n623 B.n622 10.6151
R1274 B.n622 B.n621 10.6151
R1275 B.n621 B.n74 10.6151
R1276 B.n617 B.n74 10.6151
R1277 B.n617 B.n616 10.6151
R1278 B.n616 B.n615 10.6151
R1279 B.n615 B.n76 10.6151
R1280 B.n611 B.n76 10.6151
R1281 B.n611 B.n610 10.6151
R1282 B.n610 B.n609 10.6151
R1283 B.n609 B.n78 10.6151
R1284 B.n605 B.n78 10.6151
R1285 B.n605 B.n604 10.6151
R1286 B.n604 B.n603 10.6151
R1287 B.n603 B.n80 10.6151
R1288 B.n599 B.n80 10.6151
R1289 B.n599 B.n598 10.6151
R1290 B.n598 B.n597 10.6151
R1291 B.n593 B.n82 10.6151
R1292 B.n593 B.n592 10.6151
R1293 B.n592 B.n591 10.6151
R1294 B.n591 B.n84 10.6151
R1295 B.n587 B.n84 10.6151
R1296 B.n587 B.n586 10.6151
R1297 B.n586 B.n585 10.6151
R1298 B.n585 B.n86 10.6151
R1299 B.n581 B.n86 10.6151
R1300 B.n581 B.n580 10.6151
R1301 B.n580 B.n579 10.6151
R1302 B.n579 B.n88 10.6151
R1303 B.n575 B.n88 10.6151
R1304 B.n575 B.n574 10.6151
R1305 B.n574 B.n573 10.6151
R1306 B.n573 B.n90 10.6151
R1307 B.n569 B.n90 10.6151
R1308 B.n569 B.n568 10.6151
R1309 B.n568 B.n567 10.6151
R1310 B.n567 B.n92 10.6151
R1311 B.n563 B.n92 10.6151
R1312 B.n563 B.n562 10.6151
R1313 B.n562 B.n561 10.6151
R1314 B.n561 B.n94 10.6151
R1315 B.n557 B.n94 10.6151
R1316 B.n557 B.n556 10.6151
R1317 B.n556 B.n555 10.6151
R1318 B.n555 B.n96 10.6151
R1319 B.n551 B.n96 10.6151
R1320 B.n551 B.n550 10.6151
R1321 B.n550 B.n549 10.6151
R1322 B.n549 B.n98 10.6151
R1323 B.n545 B.n98 10.6151
R1324 B.n545 B.n544 10.6151
R1325 B.n544 B.n543 10.6151
R1326 B.n543 B.n100 10.6151
R1327 B.n539 B.n100 10.6151
R1328 B.n539 B.n538 10.6151
R1329 B.n538 B.n537 10.6151
R1330 B.n537 B.n102 10.6151
R1331 B.n533 B.n102 10.6151
R1332 B.n533 B.n532 10.6151
R1333 B.n532 B.n531 10.6151
R1334 B.n531 B.n104 10.6151
R1335 B.n527 B.n104 10.6151
R1336 B.n527 B.n526 10.6151
R1337 B.n526 B.n525 10.6151
R1338 B.n525 B.n106 10.6151
R1339 B.n521 B.n106 10.6151
R1340 B.n521 B.n520 10.6151
R1341 B.n520 B.n519 10.6151
R1342 B.n519 B.n108 10.6151
R1343 B.n515 B.n108 10.6151
R1344 B.n515 B.n514 10.6151
R1345 B.n514 B.n513 10.6151
R1346 B.n513 B.n110 10.6151
R1347 B.n509 B.n110 10.6151
R1348 B.n509 B.n508 10.6151
R1349 B.n508 B.n507 10.6151
R1350 B.n507 B.n112 10.6151
R1351 B.n503 B.n112 10.6151
R1352 B.n503 B.n502 10.6151
R1353 B.n502 B.n501 10.6151
R1354 B.n501 B.n114 10.6151
R1355 B.n497 B.n114 10.6151
R1356 B.n497 B.n496 10.6151
R1357 B.n496 B.n495 10.6151
R1358 B.n495 B.n116 10.6151
R1359 B.n491 B.n116 10.6151
R1360 B.n491 B.n490 10.6151
R1361 B.n490 B.n489 10.6151
R1362 B.n489 B.n118 10.6151
R1363 B.n485 B.n118 10.6151
R1364 B.n485 B.n484 10.6151
R1365 B.n484 B.n483 10.6151
R1366 B.n483 B.n120 10.6151
R1367 B.n479 B.n120 10.6151
R1368 B.n479 B.n478 10.6151
R1369 B.n478 B.n477 10.6151
R1370 B.n477 B.n122 10.6151
R1371 B.n473 B.n122 10.6151
R1372 B.n473 B.n472 10.6151
R1373 B.n472 B.n471 10.6151
R1374 B.n471 B.n124 10.6151
R1375 B.n467 B.n124 10.6151
R1376 B.n467 B.n466 10.6151
R1377 B.n466 B.n465 10.6151
R1378 B.n465 B.n126 10.6151
R1379 B.n461 B.n126 10.6151
R1380 B.n461 B.n460 10.6151
R1381 B.n460 B.n459 10.6151
R1382 B.n459 B.n128 10.6151
R1383 B.n455 B.n128 10.6151
R1384 B.n455 B.n454 10.6151
R1385 B.n454 B.n453 10.6151
R1386 B.n453 B.n130 10.6151
R1387 B.n449 B.n130 10.6151
R1388 B.n449 B.n448 10.6151
R1389 B.n448 B.n447 10.6151
R1390 B.n447 B.n132 10.6151
R1391 B.n443 B.n132 10.6151
R1392 B.n443 B.n442 10.6151
R1393 B.n442 B.n441 10.6151
R1394 B.n211 B.n1 10.6151
R1395 B.n211 B.n210 10.6151
R1396 B.n215 B.n210 10.6151
R1397 B.n216 B.n215 10.6151
R1398 B.n217 B.n216 10.6151
R1399 B.n217 B.n208 10.6151
R1400 B.n221 B.n208 10.6151
R1401 B.n222 B.n221 10.6151
R1402 B.n223 B.n222 10.6151
R1403 B.n223 B.n206 10.6151
R1404 B.n227 B.n206 10.6151
R1405 B.n228 B.n227 10.6151
R1406 B.n229 B.n228 10.6151
R1407 B.n229 B.n204 10.6151
R1408 B.n233 B.n204 10.6151
R1409 B.n234 B.n233 10.6151
R1410 B.n235 B.n234 10.6151
R1411 B.n235 B.n202 10.6151
R1412 B.n239 B.n202 10.6151
R1413 B.n240 B.n239 10.6151
R1414 B.n241 B.n240 10.6151
R1415 B.n241 B.n200 10.6151
R1416 B.n245 B.n200 10.6151
R1417 B.n246 B.n245 10.6151
R1418 B.n247 B.n246 10.6151
R1419 B.n247 B.n198 10.6151
R1420 B.n251 B.n198 10.6151
R1421 B.n252 B.n251 10.6151
R1422 B.n253 B.n252 10.6151
R1423 B.n253 B.n196 10.6151
R1424 B.n257 B.n196 10.6151
R1425 B.n258 B.n257 10.6151
R1426 B.n259 B.n258 10.6151
R1427 B.n259 B.n194 10.6151
R1428 B.n263 B.n194 10.6151
R1429 B.n264 B.n263 10.6151
R1430 B.n265 B.n264 10.6151
R1431 B.n265 B.n192 10.6151
R1432 B.n269 B.n192 10.6151
R1433 B.n270 B.n269 10.6151
R1434 B.n271 B.n270 10.6151
R1435 B.n271 B.n190 10.6151
R1436 B.n275 B.n190 10.6151
R1437 B.n276 B.n275 10.6151
R1438 B.n277 B.n276 10.6151
R1439 B.n277 B.n188 10.6151
R1440 B.n281 B.n188 10.6151
R1441 B.n282 B.n281 10.6151
R1442 B.n283 B.n282 10.6151
R1443 B.n283 B.n186 10.6151
R1444 B.n288 B.n287 10.6151
R1445 B.n289 B.n288 10.6151
R1446 B.n289 B.n184 10.6151
R1447 B.n293 B.n184 10.6151
R1448 B.n294 B.n293 10.6151
R1449 B.n295 B.n294 10.6151
R1450 B.n295 B.n182 10.6151
R1451 B.n299 B.n182 10.6151
R1452 B.n300 B.n299 10.6151
R1453 B.n301 B.n300 10.6151
R1454 B.n301 B.n180 10.6151
R1455 B.n305 B.n180 10.6151
R1456 B.n306 B.n305 10.6151
R1457 B.n307 B.n306 10.6151
R1458 B.n307 B.n178 10.6151
R1459 B.n311 B.n178 10.6151
R1460 B.n312 B.n311 10.6151
R1461 B.n313 B.n312 10.6151
R1462 B.n313 B.n176 10.6151
R1463 B.n317 B.n176 10.6151
R1464 B.n318 B.n317 10.6151
R1465 B.n319 B.n318 10.6151
R1466 B.n319 B.n174 10.6151
R1467 B.n323 B.n174 10.6151
R1468 B.n324 B.n323 10.6151
R1469 B.n325 B.n324 10.6151
R1470 B.n325 B.n172 10.6151
R1471 B.n329 B.n172 10.6151
R1472 B.n330 B.n329 10.6151
R1473 B.n331 B.n330 10.6151
R1474 B.n331 B.n170 10.6151
R1475 B.n335 B.n170 10.6151
R1476 B.n336 B.n335 10.6151
R1477 B.n337 B.n336 10.6151
R1478 B.n337 B.n168 10.6151
R1479 B.n341 B.n168 10.6151
R1480 B.n342 B.n341 10.6151
R1481 B.n343 B.n342 10.6151
R1482 B.n343 B.n166 10.6151
R1483 B.n347 B.n166 10.6151
R1484 B.n348 B.n347 10.6151
R1485 B.n349 B.n348 10.6151
R1486 B.n349 B.n164 10.6151
R1487 B.n353 B.n164 10.6151
R1488 B.n356 B.n355 10.6151
R1489 B.n356 B.n160 10.6151
R1490 B.n360 B.n160 10.6151
R1491 B.n361 B.n360 10.6151
R1492 B.n362 B.n361 10.6151
R1493 B.n362 B.n158 10.6151
R1494 B.n366 B.n158 10.6151
R1495 B.n367 B.n366 10.6151
R1496 B.n371 B.n367 10.6151
R1497 B.n375 B.n156 10.6151
R1498 B.n376 B.n375 10.6151
R1499 B.n377 B.n376 10.6151
R1500 B.n377 B.n154 10.6151
R1501 B.n381 B.n154 10.6151
R1502 B.n382 B.n381 10.6151
R1503 B.n383 B.n382 10.6151
R1504 B.n383 B.n152 10.6151
R1505 B.n387 B.n152 10.6151
R1506 B.n388 B.n387 10.6151
R1507 B.n389 B.n388 10.6151
R1508 B.n389 B.n150 10.6151
R1509 B.n393 B.n150 10.6151
R1510 B.n394 B.n393 10.6151
R1511 B.n395 B.n394 10.6151
R1512 B.n395 B.n148 10.6151
R1513 B.n399 B.n148 10.6151
R1514 B.n400 B.n399 10.6151
R1515 B.n401 B.n400 10.6151
R1516 B.n401 B.n146 10.6151
R1517 B.n405 B.n146 10.6151
R1518 B.n406 B.n405 10.6151
R1519 B.n407 B.n406 10.6151
R1520 B.n407 B.n144 10.6151
R1521 B.n411 B.n144 10.6151
R1522 B.n412 B.n411 10.6151
R1523 B.n413 B.n412 10.6151
R1524 B.n413 B.n142 10.6151
R1525 B.n417 B.n142 10.6151
R1526 B.n418 B.n417 10.6151
R1527 B.n419 B.n418 10.6151
R1528 B.n419 B.n140 10.6151
R1529 B.n423 B.n140 10.6151
R1530 B.n424 B.n423 10.6151
R1531 B.n425 B.n424 10.6151
R1532 B.n425 B.n138 10.6151
R1533 B.n429 B.n138 10.6151
R1534 B.n430 B.n429 10.6151
R1535 B.n431 B.n430 10.6151
R1536 B.n431 B.n136 10.6151
R1537 B.n435 B.n136 10.6151
R1538 B.n436 B.n435 10.6151
R1539 B.n437 B.n436 10.6151
R1540 B.n437 B.n134 10.6151
R1541 B.n681 B.n52 9.36635
R1542 B.n664 B.n663 9.36635
R1543 B.n354 B.n353 9.36635
R1544 B.n370 B.n156 9.36635
R1545 B.n825 B.n0 8.11757
R1546 B.n825 B.n1 8.11757
R1547 B.n678 B.n52 1.24928
R1548 B.n665 B.n664 1.24928
R1549 B.n355 B.n354 1.24928
R1550 B.n371 B.n370 1.24928
C0 VN VTAIL 11.612401f
C1 VP w_n3934_n3614# 8.79832f
C2 B VP 2.03716f
C3 VN VDD2 11.2148f
C4 VTAIL w_n3934_n3614# 3.33131f
C5 VDD1 VN 0.15246f
C6 B VTAIL 3.79675f
C7 VTAIL VP 11.6267f
C8 VDD2 w_n3934_n3614# 2.82267f
C9 VDD1 w_n3934_n3614# 2.70294f
C10 B VDD2 2.49563f
C11 VDD1 B 2.39563f
C12 VDD2 VP 0.525185f
C13 VDD1 VP 11.5834f
C14 VDD2 VTAIL 11.0703f
C15 VN w_n3934_n3614# 8.28755f
C16 VDD1 VTAIL 11.0234f
C17 VN B 1.18081f
C18 VN VP 7.9464f
C19 VDD1 VDD2 1.87634f
C20 B w_n3934_n3614# 10.1181f
C21 VDD2 VSUBS 1.975756f
C22 VDD1 VSUBS 1.791936f
C23 VTAIL VSUBS 1.232821f
C24 VN VSUBS 6.98157f
C25 VP VSUBS 3.705671f
C26 B VSUBS 4.899343f
C27 w_n3934_n3614# VSUBS 0.174717p
C28 B.n0 VSUBS 0.008167f
C29 B.n1 VSUBS 0.008167f
C30 B.n2 VSUBS 0.012078f
C31 B.n3 VSUBS 0.009256f
C32 B.n4 VSUBS 0.009256f
C33 B.n5 VSUBS 0.009256f
C34 B.n6 VSUBS 0.009256f
C35 B.n7 VSUBS 0.009256f
C36 B.n8 VSUBS 0.009256f
C37 B.n9 VSUBS 0.009256f
C38 B.n10 VSUBS 0.009256f
C39 B.n11 VSUBS 0.009256f
C40 B.n12 VSUBS 0.009256f
C41 B.n13 VSUBS 0.009256f
C42 B.n14 VSUBS 0.009256f
C43 B.n15 VSUBS 0.009256f
C44 B.n16 VSUBS 0.009256f
C45 B.n17 VSUBS 0.009256f
C46 B.n18 VSUBS 0.009256f
C47 B.n19 VSUBS 0.009256f
C48 B.n20 VSUBS 0.009256f
C49 B.n21 VSUBS 0.009256f
C50 B.n22 VSUBS 0.009256f
C51 B.n23 VSUBS 0.009256f
C52 B.n24 VSUBS 0.009256f
C53 B.n25 VSUBS 0.009256f
C54 B.n26 VSUBS 0.009256f
C55 B.n27 VSUBS 0.021957f
C56 B.n28 VSUBS 0.009256f
C57 B.n29 VSUBS 0.009256f
C58 B.n30 VSUBS 0.009256f
C59 B.n31 VSUBS 0.009256f
C60 B.n32 VSUBS 0.009256f
C61 B.n33 VSUBS 0.009256f
C62 B.n34 VSUBS 0.009256f
C63 B.n35 VSUBS 0.009256f
C64 B.n36 VSUBS 0.009256f
C65 B.n37 VSUBS 0.009256f
C66 B.n38 VSUBS 0.009256f
C67 B.n39 VSUBS 0.009256f
C68 B.n40 VSUBS 0.009256f
C69 B.n41 VSUBS 0.009256f
C70 B.n42 VSUBS 0.009256f
C71 B.n43 VSUBS 0.009256f
C72 B.n44 VSUBS 0.009256f
C73 B.n45 VSUBS 0.009256f
C74 B.n46 VSUBS 0.009256f
C75 B.n47 VSUBS 0.009256f
C76 B.n48 VSUBS 0.009256f
C77 B.n49 VSUBS 0.009256f
C78 B.t7 VSUBS 0.575784f
C79 B.t8 VSUBS 0.599417f
C80 B.t6 VSUBS 1.67113f
C81 B.n50 VSUBS 0.29867f
C82 B.n51 VSUBS 0.09251f
C83 B.n52 VSUBS 0.021444f
C84 B.n53 VSUBS 0.009256f
C85 B.n54 VSUBS 0.009256f
C86 B.n55 VSUBS 0.009256f
C87 B.n56 VSUBS 0.009256f
C88 B.n57 VSUBS 0.009256f
C89 B.t10 VSUBS 0.575771f
C90 B.t11 VSUBS 0.599406f
C91 B.t9 VSUBS 1.67113f
C92 B.n58 VSUBS 0.298681f
C93 B.n59 VSUBS 0.092522f
C94 B.n60 VSUBS 0.009256f
C95 B.n61 VSUBS 0.009256f
C96 B.n62 VSUBS 0.009256f
C97 B.n63 VSUBS 0.009256f
C98 B.n64 VSUBS 0.009256f
C99 B.n65 VSUBS 0.009256f
C100 B.n66 VSUBS 0.009256f
C101 B.n67 VSUBS 0.009256f
C102 B.n68 VSUBS 0.009256f
C103 B.n69 VSUBS 0.009256f
C104 B.n70 VSUBS 0.009256f
C105 B.n71 VSUBS 0.009256f
C106 B.n72 VSUBS 0.009256f
C107 B.n73 VSUBS 0.009256f
C108 B.n74 VSUBS 0.009256f
C109 B.n75 VSUBS 0.009256f
C110 B.n76 VSUBS 0.009256f
C111 B.n77 VSUBS 0.009256f
C112 B.n78 VSUBS 0.009256f
C113 B.n79 VSUBS 0.009256f
C114 B.n80 VSUBS 0.009256f
C115 B.n81 VSUBS 0.009256f
C116 B.n82 VSUBS 0.021957f
C117 B.n83 VSUBS 0.009256f
C118 B.n84 VSUBS 0.009256f
C119 B.n85 VSUBS 0.009256f
C120 B.n86 VSUBS 0.009256f
C121 B.n87 VSUBS 0.009256f
C122 B.n88 VSUBS 0.009256f
C123 B.n89 VSUBS 0.009256f
C124 B.n90 VSUBS 0.009256f
C125 B.n91 VSUBS 0.009256f
C126 B.n92 VSUBS 0.009256f
C127 B.n93 VSUBS 0.009256f
C128 B.n94 VSUBS 0.009256f
C129 B.n95 VSUBS 0.009256f
C130 B.n96 VSUBS 0.009256f
C131 B.n97 VSUBS 0.009256f
C132 B.n98 VSUBS 0.009256f
C133 B.n99 VSUBS 0.009256f
C134 B.n100 VSUBS 0.009256f
C135 B.n101 VSUBS 0.009256f
C136 B.n102 VSUBS 0.009256f
C137 B.n103 VSUBS 0.009256f
C138 B.n104 VSUBS 0.009256f
C139 B.n105 VSUBS 0.009256f
C140 B.n106 VSUBS 0.009256f
C141 B.n107 VSUBS 0.009256f
C142 B.n108 VSUBS 0.009256f
C143 B.n109 VSUBS 0.009256f
C144 B.n110 VSUBS 0.009256f
C145 B.n111 VSUBS 0.009256f
C146 B.n112 VSUBS 0.009256f
C147 B.n113 VSUBS 0.009256f
C148 B.n114 VSUBS 0.009256f
C149 B.n115 VSUBS 0.009256f
C150 B.n116 VSUBS 0.009256f
C151 B.n117 VSUBS 0.009256f
C152 B.n118 VSUBS 0.009256f
C153 B.n119 VSUBS 0.009256f
C154 B.n120 VSUBS 0.009256f
C155 B.n121 VSUBS 0.009256f
C156 B.n122 VSUBS 0.009256f
C157 B.n123 VSUBS 0.009256f
C158 B.n124 VSUBS 0.009256f
C159 B.n125 VSUBS 0.009256f
C160 B.n126 VSUBS 0.009256f
C161 B.n127 VSUBS 0.009256f
C162 B.n128 VSUBS 0.009256f
C163 B.n129 VSUBS 0.009256f
C164 B.n130 VSUBS 0.009256f
C165 B.n131 VSUBS 0.009256f
C166 B.n132 VSUBS 0.009256f
C167 B.n133 VSUBS 0.009256f
C168 B.n134 VSUBS 0.022207f
C169 B.n135 VSUBS 0.009256f
C170 B.n136 VSUBS 0.009256f
C171 B.n137 VSUBS 0.009256f
C172 B.n138 VSUBS 0.009256f
C173 B.n139 VSUBS 0.009256f
C174 B.n140 VSUBS 0.009256f
C175 B.n141 VSUBS 0.009256f
C176 B.n142 VSUBS 0.009256f
C177 B.n143 VSUBS 0.009256f
C178 B.n144 VSUBS 0.009256f
C179 B.n145 VSUBS 0.009256f
C180 B.n146 VSUBS 0.009256f
C181 B.n147 VSUBS 0.009256f
C182 B.n148 VSUBS 0.009256f
C183 B.n149 VSUBS 0.009256f
C184 B.n150 VSUBS 0.009256f
C185 B.n151 VSUBS 0.009256f
C186 B.n152 VSUBS 0.009256f
C187 B.n153 VSUBS 0.009256f
C188 B.n154 VSUBS 0.009256f
C189 B.n155 VSUBS 0.009256f
C190 B.n156 VSUBS 0.008711f
C191 B.n157 VSUBS 0.009256f
C192 B.n158 VSUBS 0.009256f
C193 B.n159 VSUBS 0.009256f
C194 B.n160 VSUBS 0.009256f
C195 B.n161 VSUBS 0.009256f
C196 B.t2 VSUBS 0.575784f
C197 B.t1 VSUBS 0.599417f
C198 B.t0 VSUBS 1.67113f
C199 B.n162 VSUBS 0.29867f
C200 B.n163 VSUBS 0.09251f
C201 B.n164 VSUBS 0.009256f
C202 B.n165 VSUBS 0.009256f
C203 B.n166 VSUBS 0.009256f
C204 B.n167 VSUBS 0.009256f
C205 B.n168 VSUBS 0.009256f
C206 B.n169 VSUBS 0.009256f
C207 B.n170 VSUBS 0.009256f
C208 B.n171 VSUBS 0.009256f
C209 B.n172 VSUBS 0.009256f
C210 B.n173 VSUBS 0.009256f
C211 B.n174 VSUBS 0.009256f
C212 B.n175 VSUBS 0.009256f
C213 B.n176 VSUBS 0.009256f
C214 B.n177 VSUBS 0.009256f
C215 B.n178 VSUBS 0.009256f
C216 B.n179 VSUBS 0.009256f
C217 B.n180 VSUBS 0.009256f
C218 B.n181 VSUBS 0.009256f
C219 B.n182 VSUBS 0.009256f
C220 B.n183 VSUBS 0.009256f
C221 B.n184 VSUBS 0.009256f
C222 B.n185 VSUBS 0.009256f
C223 B.n186 VSUBS 0.021957f
C224 B.n187 VSUBS 0.009256f
C225 B.n188 VSUBS 0.009256f
C226 B.n189 VSUBS 0.009256f
C227 B.n190 VSUBS 0.009256f
C228 B.n191 VSUBS 0.009256f
C229 B.n192 VSUBS 0.009256f
C230 B.n193 VSUBS 0.009256f
C231 B.n194 VSUBS 0.009256f
C232 B.n195 VSUBS 0.009256f
C233 B.n196 VSUBS 0.009256f
C234 B.n197 VSUBS 0.009256f
C235 B.n198 VSUBS 0.009256f
C236 B.n199 VSUBS 0.009256f
C237 B.n200 VSUBS 0.009256f
C238 B.n201 VSUBS 0.009256f
C239 B.n202 VSUBS 0.009256f
C240 B.n203 VSUBS 0.009256f
C241 B.n204 VSUBS 0.009256f
C242 B.n205 VSUBS 0.009256f
C243 B.n206 VSUBS 0.009256f
C244 B.n207 VSUBS 0.009256f
C245 B.n208 VSUBS 0.009256f
C246 B.n209 VSUBS 0.009256f
C247 B.n210 VSUBS 0.009256f
C248 B.n211 VSUBS 0.009256f
C249 B.n212 VSUBS 0.009256f
C250 B.n213 VSUBS 0.009256f
C251 B.n214 VSUBS 0.009256f
C252 B.n215 VSUBS 0.009256f
C253 B.n216 VSUBS 0.009256f
C254 B.n217 VSUBS 0.009256f
C255 B.n218 VSUBS 0.009256f
C256 B.n219 VSUBS 0.009256f
C257 B.n220 VSUBS 0.009256f
C258 B.n221 VSUBS 0.009256f
C259 B.n222 VSUBS 0.009256f
C260 B.n223 VSUBS 0.009256f
C261 B.n224 VSUBS 0.009256f
C262 B.n225 VSUBS 0.009256f
C263 B.n226 VSUBS 0.009256f
C264 B.n227 VSUBS 0.009256f
C265 B.n228 VSUBS 0.009256f
C266 B.n229 VSUBS 0.009256f
C267 B.n230 VSUBS 0.009256f
C268 B.n231 VSUBS 0.009256f
C269 B.n232 VSUBS 0.009256f
C270 B.n233 VSUBS 0.009256f
C271 B.n234 VSUBS 0.009256f
C272 B.n235 VSUBS 0.009256f
C273 B.n236 VSUBS 0.009256f
C274 B.n237 VSUBS 0.009256f
C275 B.n238 VSUBS 0.009256f
C276 B.n239 VSUBS 0.009256f
C277 B.n240 VSUBS 0.009256f
C278 B.n241 VSUBS 0.009256f
C279 B.n242 VSUBS 0.009256f
C280 B.n243 VSUBS 0.009256f
C281 B.n244 VSUBS 0.009256f
C282 B.n245 VSUBS 0.009256f
C283 B.n246 VSUBS 0.009256f
C284 B.n247 VSUBS 0.009256f
C285 B.n248 VSUBS 0.009256f
C286 B.n249 VSUBS 0.009256f
C287 B.n250 VSUBS 0.009256f
C288 B.n251 VSUBS 0.009256f
C289 B.n252 VSUBS 0.009256f
C290 B.n253 VSUBS 0.009256f
C291 B.n254 VSUBS 0.009256f
C292 B.n255 VSUBS 0.009256f
C293 B.n256 VSUBS 0.009256f
C294 B.n257 VSUBS 0.009256f
C295 B.n258 VSUBS 0.009256f
C296 B.n259 VSUBS 0.009256f
C297 B.n260 VSUBS 0.009256f
C298 B.n261 VSUBS 0.009256f
C299 B.n262 VSUBS 0.009256f
C300 B.n263 VSUBS 0.009256f
C301 B.n264 VSUBS 0.009256f
C302 B.n265 VSUBS 0.009256f
C303 B.n266 VSUBS 0.009256f
C304 B.n267 VSUBS 0.009256f
C305 B.n268 VSUBS 0.009256f
C306 B.n269 VSUBS 0.009256f
C307 B.n270 VSUBS 0.009256f
C308 B.n271 VSUBS 0.009256f
C309 B.n272 VSUBS 0.009256f
C310 B.n273 VSUBS 0.009256f
C311 B.n274 VSUBS 0.009256f
C312 B.n275 VSUBS 0.009256f
C313 B.n276 VSUBS 0.009256f
C314 B.n277 VSUBS 0.009256f
C315 B.n278 VSUBS 0.009256f
C316 B.n279 VSUBS 0.009256f
C317 B.n280 VSUBS 0.009256f
C318 B.n281 VSUBS 0.009256f
C319 B.n282 VSUBS 0.009256f
C320 B.n283 VSUBS 0.009256f
C321 B.n284 VSUBS 0.009256f
C322 B.n285 VSUBS 0.021957f
C323 B.n286 VSUBS 0.023233f
C324 B.n287 VSUBS 0.023233f
C325 B.n288 VSUBS 0.009256f
C326 B.n289 VSUBS 0.009256f
C327 B.n290 VSUBS 0.009256f
C328 B.n291 VSUBS 0.009256f
C329 B.n292 VSUBS 0.009256f
C330 B.n293 VSUBS 0.009256f
C331 B.n294 VSUBS 0.009256f
C332 B.n295 VSUBS 0.009256f
C333 B.n296 VSUBS 0.009256f
C334 B.n297 VSUBS 0.009256f
C335 B.n298 VSUBS 0.009256f
C336 B.n299 VSUBS 0.009256f
C337 B.n300 VSUBS 0.009256f
C338 B.n301 VSUBS 0.009256f
C339 B.n302 VSUBS 0.009256f
C340 B.n303 VSUBS 0.009256f
C341 B.n304 VSUBS 0.009256f
C342 B.n305 VSUBS 0.009256f
C343 B.n306 VSUBS 0.009256f
C344 B.n307 VSUBS 0.009256f
C345 B.n308 VSUBS 0.009256f
C346 B.n309 VSUBS 0.009256f
C347 B.n310 VSUBS 0.009256f
C348 B.n311 VSUBS 0.009256f
C349 B.n312 VSUBS 0.009256f
C350 B.n313 VSUBS 0.009256f
C351 B.n314 VSUBS 0.009256f
C352 B.n315 VSUBS 0.009256f
C353 B.n316 VSUBS 0.009256f
C354 B.n317 VSUBS 0.009256f
C355 B.n318 VSUBS 0.009256f
C356 B.n319 VSUBS 0.009256f
C357 B.n320 VSUBS 0.009256f
C358 B.n321 VSUBS 0.009256f
C359 B.n322 VSUBS 0.009256f
C360 B.n323 VSUBS 0.009256f
C361 B.n324 VSUBS 0.009256f
C362 B.n325 VSUBS 0.009256f
C363 B.n326 VSUBS 0.009256f
C364 B.n327 VSUBS 0.009256f
C365 B.n328 VSUBS 0.009256f
C366 B.n329 VSUBS 0.009256f
C367 B.n330 VSUBS 0.009256f
C368 B.n331 VSUBS 0.009256f
C369 B.n332 VSUBS 0.009256f
C370 B.n333 VSUBS 0.009256f
C371 B.n334 VSUBS 0.009256f
C372 B.n335 VSUBS 0.009256f
C373 B.n336 VSUBS 0.009256f
C374 B.n337 VSUBS 0.009256f
C375 B.n338 VSUBS 0.009256f
C376 B.n339 VSUBS 0.009256f
C377 B.n340 VSUBS 0.009256f
C378 B.n341 VSUBS 0.009256f
C379 B.n342 VSUBS 0.009256f
C380 B.n343 VSUBS 0.009256f
C381 B.n344 VSUBS 0.009256f
C382 B.n345 VSUBS 0.009256f
C383 B.n346 VSUBS 0.009256f
C384 B.n347 VSUBS 0.009256f
C385 B.n348 VSUBS 0.009256f
C386 B.n349 VSUBS 0.009256f
C387 B.n350 VSUBS 0.009256f
C388 B.n351 VSUBS 0.009256f
C389 B.n352 VSUBS 0.009256f
C390 B.n353 VSUBS 0.008711f
C391 B.n354 VSUBS 0.021444f
C392 B.n355 VSUBS 0.005172f
C393 B.n356 VSUBS 0.009256f
C394 B.n357 VSUBS 0.009256f
C395 B.n358 VSUBS 0.009256f
C396 B.n359 VSUBS 0.009256f
C397 B.n360 VSUBS 0.009256f
C398 B.n361 VSUBS 0.009256f
C399 B.n362 VSUBS 0.009256f
C400 B.n363 VSUBS 0.009256f
C401 B.n364 VSUBS 0.009256f
C402 B.n365 VSUBS 0.009256f
C403 B.n366 VSUBS 0.009256f
C404 B.n367 VSUBS 0.009256f
C405 B.t5 VSUBS 0.575771f
C406 B.t4 VSUBS 0.599406f
C407 B.t3 VSUBS 1.67113f
C408 B.n368 VSUBS 0.298681f
C409 B.n369 VSUBS 0.092522f
C410 B.n370 VSUBS 0.021444f
C411 B.n371 VSUBS 0.005172f
C412 B.n372 VSUBS 0.009256f
C413 B.n373 VSUBS 0.009256f
C414 B.n374 VSUBS 0.009256f
C415 B.n375 VSUBS 0.009256f
C416 B.n376 VSUBS 0.009256f
C417 B.n377 VSUBS 0.009256f
C418 B.n378 VSUBS 0.009256f
C419 B.n379 VSUBS 0.009256f
C420 B.n380 VSUBS 0.009256f
C421 B.n381 VSUBS 0.009256f
C422 B.n382 VSUBS 0.009256f
C423 B.n383 VSUBS 0.009256f
C424 B.n384 VSUBS 0.009256f
C425 B.n385 VSUBS 0.009256f
C426 B.n386 VSUBS 0.009256f
C427 B.n387 VSUBS 0.009256f
C428 B.n388 VSUBS 0.009256f
C429 B.n389 VSUBS 0.009256f
C430 B.n390 VSUBS 0.009256f
C431 B.n391 VSUBS 0.009256f
C432 B.n392 VSUBS 0.009256f
C433 B.n393 VSUBS 0.009256f
C434 B.n394 VSUBS 0.009256f
C435 B.n395 VSUBS 0.009256f
C436 B.n396 VSUBS 0.009256f
C437 B.n397 VSUBS 0.009256f
C438 B.n398 VSUBS 0.009256f
C439 B.n399 VSUBS 0.009256f
C440 B.n400 VSUBS 0.009256f
C441 B.n401 VSUBS 0.009256f
C442 B.n402 VSUBS 0.009256f
C443 B.n403 VSUBS 0.009256f
C444 B.n404 VSUBS 0.009256f
C445 B.n405 VSUBS 0.009256f
C446 B.n406 VSUBS 0.009256f
C447 B.n407 VSUBS 0.009256f
C448 B.n408 VSUBS 0.009256f
C449 B.n409 VSUBS 0.009256f
C450 B.n410 VSUBS 0.009256f
C451 B.n411 VSUBS 0.009256f
C452 B.n412 VSUBS 0.009256f
C453 B.n413 VSUBS 0.009256f
C454 B.n414 VSUBS 0.009256f
C455 B.n415 VSUBS 0.009256f
C456 B.n416 VSUBS 0.009256f
C457 B.n417 VSUBS 0.009256f
C458 B.n418 VSUBS 0.009256f
C459 B.n419 VSUBS 0.009256f
C460 B.n420 VSUBS 0.009256f
C461 B.n421 VSUBS 0.009256f
C462 B.n422 VSUBS 0.009256f
C463 B.n423 VSUBS 0.009256f
C464 B.n424 VSUBS 0.009256f
C465 B.n425 VSUBS 0.009256f
C466 B.n426 VSUBS 0.009256f
C467 B.n427 VSUBS 0.009256f
C468 B.n428 VSUBS 0.009256f
C469 B.n429 VSUBS 0.009256f
C470 B.n430 VSUBS 0.009256f
C471 B.n431 VSUBS 0.009256f
C472 B.n432 VSUBS 0.009256f
C473 B.n433 VSUBS 0.009256f
C474 B.n434 VSUBS 0.009256f
C475 B.n435 VSUBS 0.009256f
C476 B.n436 VSUBS 0.009256f
C477 B.n437 VSUBS 0.009256f
C478 B.n438 VSUBS 0.009256f
C479 B.n439 VSUBS 0.023233f
C480 B.n440 VSUBS 0.021957f
C481 B.n441 VSUBS 0.022983f
C482 B.n442 VSUBS 0.009256f
C483 B.n443 VSUBS 0.009256f
C484 B.n444 VSUBS 0.009256f
C485 B.n445 VSUBS 0.009256f
C486 B.n446 VSUBS 0.009256f
C487 B.n447 VSUBS 0.009256f
C488 B.n448 VSUBS 0.009256f
C489 B.n449 VSUBS 0.009256f
C490 B.n450 VSUBS 0.009256f
C491 B.n451 VSUBS 0.009256f
C492 B.n452 VSUBS 0.009256f
C493 B.n453 VSUBS 0.009256f
C494 B.n454 VSUBS 0.009256f
C495 B.n455 VSUBS 0.009256f
C496 B.n456 VSUBS 0.009256f
C497 B.n457 VSUBS 0.009256f
C498 B.n458 VSUBS 0.009256f
C499 B.n459 VSUBS 0.009256f
C500 B.n460 VSUBS 0.009256f
C501 B.n461 VSUBS 0.009256f
C502 B.n462 VSUBS 0.009256f
C503 B.n463 VSUBS 0.009256f
C504 B.n464 VSUBS 0.009256f
C505 B.n465 VSUBS 0.009256f
C506 B.n466 VSUBS 0.009256f
C507 B.n467 VSUBS 0.009256f
C508 B.n468 VSUBS 0.009256f
C509 B.n469 VSUBS 0.009256f
C510 B.n470 VSUBS 0.009256f
C511 B.n471 VSUBS 0.009256f
C512 B.n472 VSUBS 0.009256f
C513 B.n473 VSUBS 0.009256f
C514 B.n474 VSUBS 0.009256f
C515 B.n475 VSUBS 0.009256f
C516 B.n476 VSUBS 0.009256f
C517 B.n477 VSUBS 0.009256f
C518 B.n478 VSUBS 0.009256f
C519 B.n479 VSUBS 0.009256f
C520 B.n480 VSUBS 0.009256f
C521 B.n481 VSUBS 0.009256f
C522 B.n482 VSUBS 0.009256f
C523 B.n483 VSUBS 0.009256f
C524 B.n484 VSUBS 0.009256f
C525 B.n485 VSUBS 0.009256f
C526 B.n486 VSUBS 0.009256f
C527 B.n487 VSUBS 0.009256f
C528 B.n488 VSUBS 0.009256f
C529 B.n489 VSUBS 0.009256f
C530 B.n490 VSUBS 0.009256f
C531 B.n491 VSUBS 0.009256f
C532 B.n492 VSUBS 0.009256f
C533 B.n493 VSUBS 0.009256f
C534 B.n494 VSUBS 0.009256f
C535 B.n495 VSUBS 0.009256f
C536 B.n496 VSUBS 0.009256f
C537 B.n497 VSUBS 0.009256f
C538 B.n498 VSUBS 0.009256f
C539 B.n499 VSUBS 0.009256f
C540 B.n500 VSUBS 0.009256f
C541 B.n501 VSUBS 0.009256f
C542 B.n502 VSUBS 0.009256f
C543 B.n503 VSUBS 0.009256f
C544 B.n504 VSUBS 0.009256f
C545 B.n505 VSUBS 0.009256f
C546 B.n506 VSUBS 0.009256f
C547 B.n507 VSUBS 0.009256f
C548 B.n508 VSUBS 0.009256f
C549 B.n509 VSUBS 0.009256f
C550 B.n510 VSUBS 0.009256f
C551 B.n511 VSUBS 0.009256f
C552 B.n512 VSUBS 0.009256f
C553 B.n513 VSUBS 0.009256f
C554 B.n514 VSUBS 0.009256f
C555 B.n515 VSUBS 0.009256f
C556 B.n516 VSUBS 0.009256f
C557 B.n517 VSUBS 0.009256f
C558 B.n518 VSUBS 0.009256f
C559 B.n519 VSUBS 0.009256f
C560 B.n520 VSUBS 0.009256f
C561 B.n521 VSUBS 0.009256f
C562 B.n522 VSUBS 0.009256f
C563 B.n523 VSUBS 0.009256f
C564 B.n524 VSUBS 0.009256f
C565 B.n525 VSUBS 0.009256f
C566 B.n526 VSUBS 0.009256f
C567 B.n527 VSUBS 0.009256f
C568 B.n528 VSUBS 0.009256f
C569 B.n529 VSUBS 0.009256f
C570 B.n530 VSUBS 0.009256f
C571 B.n531 VSUBS 0.009256f
C572 B.n532 VSUBS 0.009256f
C573 B.n533 VSUBS 0.009256f
C574 B.n534 VSUBS 0.009256f
C575 B.n535 VSUBS 0.009256f
C576 B.n536 VSUBS 0.009256f
C577 B.n537 VSUBS 0.009256f
C578 B.n538 VSUBS 0.009256f
C579 B.n539 VSUBS 0.009256f
C580 B.n540 VSUBS 0.009256f
C581 B.n541 VSUBS 0.009256f
C582 B.n542 VSUBS 0.009256f
C583 B.n543 VSUBS 0.009256f
C584 B.n544 VSUBS 0.009256f
C585 B.n545 VSUBS 0.009256f
C586 B.n546 VSUBS 0.009256f
C587 B.n547 VSUBS 0.009256f
C588 B.n548 VSUBS 0.009256f
C589 B.n549 VSUBS 0.009256f
C590 B.n550 VSUBS 0.009256f
C591 B.n551 VSUBS 0.009256f
C592 B.n552 VSUBS 0.009256f
C593 B.n553 VSUBS 0.009256f
C594 B.n554 VSUBS 0.009256f
C595 B.n555 VSUBS 0.009256f
C596 B.n556 VSUBS 0.009256f
C597 B.n557 VSUBS 0.009256f
C598 B.n558 VSUBS 0.009256f
C599 B.n559 VSUBS 0.009256f
C600 B.n560 VSUBS 0.009256f
C601 B.n561 VSUBS 0.009256f
C602 B.n562 VSUBS 0.009256f
C603 B.n563 VSUBS 0.009256f
C604 B.n564 VSUBS 0.009256f
C605 B.n565 VSUBS 0.009256f
C606 B.n566 VSUBS 0.009256f
C607 B.n567 VSUBS 0.009256f
C608 B.n568 VSUBS 0.009256f
C609 B.n569 VSUBS 0.009256f
C610 B.n570 VSUBS 0.009256f
C611 B.n571 VSUBS 0.009256f
C612 B.n572 VSUBS 0.009256f
C613 B.n573 VSUBS 0.009256f
C614 B.n574 VSUBS 0.009256f
C615 B.n575 VSUBS 0.009256f
C616 B.n576 VSUBS 0.009256f
C617 B.n577 VSUBS 0.009256f
C618 B.n578 VSUBS 0.009256f
C619 B.n579 VSUBS 0.009256f
C620 B.n580 VSUBS 0.009256f
C621 B.n581 VSUBS 0.009256f
C622 B.n582 VSUBS 0.009256f
C623 B.n583 VSUBS 0.009256f
C624 B.n584 VSUBS 0.009256f
C625 B.n585 VSUBS 0.009256f
C626 B.n586 VSUBS 0.009256f
C627 B.n587 VSUBS 0.009256f
C628 B.n588 VSUBS 0.009256f
C629 B.n589 VSUBS 0.009256f
C630 B.n590 VSUBS 0.009256f
C631 B.n591 VSUBS 0.009256f
C632 B.n592 VSUBS 0.009256f
C633 B.n593 VSUBS 0.009256f
C634 B.n594 VSUBS 0.009256f
C635 B.n595 VSUBS 0.021957f
C636 B.n596 VSUBS 0.023233f
C637 B.n597 VSUBS 0.023233f
C638 B.n598 VSUBS 0.009256f
C639 B.n599 VSUBS 0.009256f
C640 B.n600 VSUBS 0.009256f
C641 B.n601 VSUBS 0.009256f
C642 B.n602 VSUBS 0.009256f
C643 B.n603 VSUBS 0.009256f
C644 B.n604 VSUBS 0.009256f
C645 B.n605 VSUBS 0.009256f
C646 B.n606 VSUBS 0.009256f
C647 B.n607 VSUBS 0.009256f
C648 B.n608 VSUBS 0.009256f
C649 B.n609 VSUBS 0.009256f
C650 B.n610 VSUBS 0.009256f
C651 B.n611 VSUBS 0.009256f
C652 B.n612 VSUBS 0.009256f
C653 B.n613 VSUBS 0.009256f
C654 B.n614 VSUBS 0.009256f
C655 B.n615 VSUBS 0.009256f
C656 B.n616 VSUBS 0.009256f
C657 B.n617 VSUBS 0.009256f
C658 B.n618 VSUBS 0.009256f
C659 B.n619 VSUBS 0.009256f
C660 B.n620 VSUBS 0.009256f
C661 B.n621 VSUBS 0.009256f
C662 B.n622 VSUBS 0.009256f
C663 B.n623 VSUBS 0.009256f
C664 B.n624 VSUBS 0.009256f
C665 B.n625 VSUBS 0.009256f
C666 B.n626 VSUBS 0.009256f
C667 B.n627 VSUBS 0.009256f
C668 B.n628 VSUBS 0.009256f
C669 B.n629 VSUBS 0.009256f
C670 B.n630 VSUBS 0.009256f
C671 B.n631 VSUBS 0.009256f
C672 B.n632 VSUBS 0.009256f
C673 B.n633 VSUBS 0.009256f
C674 B.n634 VSUBS 0.009256f
C675 B.n635 VSUBS 0.009256f
C676 B.n636 VSUBS 0.009256f
C677 B.n637 VSUBS 0.009256f
C678 B.n638 VSUBS 0.009256f
C679 B.n639 VSUBS 0.009256f
C680 B.n640 VSUBS 0.009256f
C681 B.n641 VSUBS 0.009256f
C682 B.n642 VSUBS 0.009256f
C683 B.n643 VSUBS 0.009256f
C684 B.n644 VSUBS 0.009256f
C685 B.n645 VSUBS 0.009256f
C686 B.n646 VSUBS 0.009256f
C687 B.n647 VSUBS 0.009256f
C688 B.n648 VSUBS 0.009256f
C689 B.n649 VSUBS 0.009256f
C690 B.n650 VSUBS 0.009256f
C691 B.n651 VSUBS 0.009256f
C692 B.n652 VSUBS 0.009256f
C693 B.n653 VSUBS 0.009256f
C694 B.n654 VSUBS 0.009256f
C695 B.n655 VSUBS 0.009256f
C696 B.n656 VSUBS 0.009256f
C697 B.n657 VSUBS 0.009256f
C698 B.n658 VSUBS 0.009256f
C699 B.n659 VSUBS 0.009256f
C700 B.n660 VSUBS 0.009256f
C701 B.n661 VSUBS 0.009256f
C702 B.n662 VSUBS 0.009256f
C703 B.n663 VSUBS 0.008711f
C704 B.n664 VSUBS 0.021444f
C705 B.n665 VSUBS 0.005172f
C706 B.n666 VSUBS 0.009256f
C707 B.n667 VSUBS 0.009256f
C708 B.n668 VSUBS 0.009256f
C709 B.n669 VSUBS 0.009256f
C710 B.n670 VSUBS 0.009256f
C711 B.n671 VSUBS 0.009256f
C712 B.n672 VSUBS 0.009256f
C713 B.n673 VSUBS 0.009256f
C714 B.n674 VSUBS 0.009256f
C715 B.n675 VSUBS 0.009256f
C716 B.n676 VSUBS 0.009256f
C717 B.n677 VSUBS 0.009256f
C718 B.n678 VSUBS 0.005172f
C719 B.n679 VSUBS 0.009256f
C720 B.n680 VSUBS 0.009256f
C721 B.n681 VSUBS 0.008711f
C722 B.n682 VSUBS 0.009256f
C723 B.n683 VSUBS 0.009256f
C724 B.n684 VSUBS 0.009256f
C725 B.n685 VSUBS 0.009256f
C726 B.n686 VSUBS 0.009256f
C727 B.n687 VSUBS 0.009256f
C728 B.n688 VSUBS 0.009256f
C729 B.n689 VSUBS 0.009256f
C730 B.n690 VSUBS 0.009256f
C731 B.n691 VSUBS 0.009256f
C732 B.n692 VSUBS 0.009256f
C733 B.n693 VSUBS 0.009256f
C734 B.n694 VSUBS 0.009256f
C735 B.n695 VSUBS 0.009256f
C736 B.n696 VSUBS 0.009256f
C737 B.n697 VSUBS 0.009256f
C738 B.n698 VSUBS 0.009256f
C739 B.n699 VSUBS 0.009256f
C740 B.n700 VSUBS 0.009256f
C741 B.n701 VSUBS 0.009256f
C742 B.n702 VSUBS 0.009256f
C743 B.n703 VSUBS 0.009256f
C744 B.n704 VSUBS 0.009256f
C745 B.n705 VSUBS 0.009256f
C746 B.n706 VSUBS 0.009256f
C747 B.n707 VSUBS 0.009256f
C748 B.n708 VSUBS 0.009256f
C749 B.n709 VSUBS 0.009256f
C750 B.n710 VSUBS 0.009256f
C751 B.n711 VSUBS 0.009256f
C752 B.n712 VSUBS 0.009256f
C753 B.n713 VSUBS 0.009256f
C754 B.n714 VSUBS 0.009256f
C755 B.n715 VSUBS 0.009256f
C756 B.n716 VSUBS 0.009256f
C757 B.n717 VSUBS 0.009256f
C758 B.n718 VSUBS 0.009256f
C759 B.n719 VSUBS 0.009256f
C760 B.n720 VSUBS 0.009256f
C761 B.n721 VSUBS 0.009256f
C762 B.n722 VSUBS 0.009256f
C763 B.n723 VSUBS 0.009256f
C764 B.n724 VSUBS 0.009256f
C765 B.n725 VSUBS 0.009256f
C766 B.n726 VSUBS 0.009256f
C767 B.n727 VSUBS 0.009256f
C768 B.n728 VSUBS 0.009256f
C769 B.n729 VSUBS 0.009256f
C770 B.n730 VSUBS 0.009256f
C771 B.n731 VSUBS 0.009256f
C772 B.n732 VSUBS 0.009256f
C773 B.n733 VSUBS 0.009256f
C774 B.n734 VSUBS 0.009256f
C775 B.n735 VSUBS 0.009256f
C776 B.n736 VSUBS 0.009256f
C777 B.n737 VSUBS 0.009256f
C778 B.n738 VSUBS 0.009256f
C779 B.n739 VSUBS 0.009256f
C780 B.n740 VSUBS 0.009256f
C781 B.n741 VSUBS 0.009256f
C782 B.n742 VSUBS 0.009256f
C783 B.n743 VSUBS 0.009256f
C784 B.n744 VSUBS 0.009256f
C785 B.n745 VSUBS 0.009256f
C786 B.n746 VSUBS 0.023233f
C787 B.n747 VSUBS 0.023233f
C788 B.n748 VSUBS 0.021957f
C789 B.n749 VSUBS 0.009256f
C790 B.n750 VSUBS 0.009256f
C791 B.n751 VSUBS 0.009256f
C792 B.n752 VSUBS 0.009256f
C793 B.n753 VSUBS 0.009256f
C794 B.n754 VSUBS 0.009256f
C795 B.n755 VSUBS 0.009256f
C796 B.n756 VSUBS 0.009256f
C797 B.n757 VSUBS 0.009256f
C798 B.n758 VSUBS 0.009256f
C799 B.n759 VSUBS 0.009256f
C800 B.n760 VSUBS 0.009256f
C801 B.n761 VSUBS 0.009256f
C802 B.n762 VSUBS 0.009256f
C803 B.n763 VSUBS 0.009256f
C804 B.n764 VSUBS 0.009256f
C805 B.n765 VSUBS 0.009256f
C806 B.n766 VSUBS 0.009256f
C807 B.n767 VSUBS 0.009256f
C808 B.n768 VSUBS 0.009256f
C809 B.n769 VSUBS 0.009256f
C810 B.n770 VSUBS 0.009256f
C811 B.n771 VSUBS 0.009256f
C812 B.n772 VSUBS 0.009256f
C813 B.n773 VSUBS 0.009256f
C814 B.n774 VSUBS 0.009256f
C815 B.n775 VSUBS 0.009256f
C816 B.n776 VSUBS 0.009256f
C817 B.n777 VSUBS 0.009256f
C818 B.n778 VSUBS 0.009256f
C819 B.n779 VSUBS 0.009256f
C820 B.n780 VSUBS 0.009256f
C821 B.n781 VSUBS 0.009256f
C822 B.n782 VSUBS 0.009256f
C823 B.n783 VSUBS 0.009256f
C824 B.n784 VSUBS 0.009256f
C825 B.n785 VSUBS 0.009256f
C826 B.n786 VSUBS 0.009256f
C827 B.n787 VSUBS 0.009256f
C828 B.n788 VSUBS 0.009256f
C829 B.n789 VSUBS 0.009256f
C830 B.n790 VSUBS 0.009256f
C831 B.n791 VSUBS 0.009256f
C832 B.n792 VSUBS 0.009256f
C833 B.n793 VSUBS 0.009256f
C834 B.n794 VSUBS 0.009256f
C835 B.n795 VSUBS 0.009256f
C836 B.n796 VSUBS 0.009256f
C837 B.n797 VSUBS 0.009256f
C838 B.n798 VSUBS 0.009256f
C839 B.n799 VSUBS 0.009256f
C840 B.n800 VSUBS 0.009256f
C841 B.n801 VSUBS 0.009256f
C842 B.n802 VSUBS 0.009256f
C843 B.n803 VSUBS 0.009256f
C844 B.n804 VSUBS 0.009256f
C845 B.n805 VSUBS 0.009256f
C846 B.n806 VSUBS 0.009256f
C847 B.n807 VSUBS 0.009256f
C848 B.n808 VSUBS 0.009256f
C849 B.n809 VSUBS 0.009256f
C850 B.n810 VSUBS 0.009256f
C851 B.n811 VSUBS 0.009256f
C852 B.n812 VSUBS 0.009256f
C853 B.n813 VSUBS 0.009256f
C854 B.n814 VSUBS 0.009256f
C855 B.n815 VSUBS 0.009256f
C856 B.n816 VSUBS 0.009256f
C857 B.n817 VSUBS 0.009256f
C858 B.n818 VSUBS 0.009256f
C859 B.n819 VSUBS 0.009256f
C860 B.n820 VSUBS 0.009256f
C861 B.n821 VSUBS 0.009256f
C862 B.n822 VSUBS 0.009256f
C863 B.n823 VSUBS 0.012078f
C864 B.n824 VSUBS 0.012866f
C865 B.n825 VSUBS 0.025586f
C866 VDD1.t8 VSUBS 2.9817f
C867 VDD1.t6 VSUBS 0.285974f
C868 VDD1.t1 VSUBS 0.285974f
C869 VDD1.n0 VSUBS 2.26933f
C870 VDD1.n1 VSUBS 1.54869f
C871 VDD1.t2 VSUBS 2.9817f
C872 VDD1.t7 VSUBS 0.285974f
C873 VDD1.t3 VSUBS 0.285974f
C874 VDD1.n2 VSUBS 2.26932f
C875 VDD1.n3 VSUBS 1.54003f
C876 VDD1.t4 VSUBS 0.285974f
C877 VDD1.t0 VSUBS 0.285974f
C878 VDD1.n4 VSUBS 2.28698f
C879 VDD1.n5 VSUBS 3.41503f
C880 VDD1.t9 VSUBS 0.285974f
C881 VDD1.t5 VSUBS 0.285974f
C882 VDD1.n6 VSUBS 2.26932f
C883 VDD1.n7 VSUBS 3.66243f
C884 VP.n0 VSUBS 0.043165f
C885 VP.t9 VSUBS 2.53229f
C886 VP.n1 VSUBS 0.043692f
C887 VP.n2 VSUBS 0.03274f
C888 VP.t5 VSUBS 2.53229f
C889 VP.n3 VSUBS 0.049166f
C890 VP.n4 VSUBS 0.03274f
C891 VP.t6 VSUBS 2.53229f
C892 VP.n5 VSUBS 0.061019f
C893 VP.n6 VSUBS 0.03274f
C894 VP.t2 VSUBS 2.53229f
C895 VP.n7 VSUBS 0.896039f
C896 VP.n8 VSUBS 0.03274f
C897 VP.n9 VSUBS 0.051903f
C898 VP.n10 VSUBS 0.043165f
C899 VP.t4 VSUBS 2.53229f
C900 VP.n11 VSUBS 0.043692f
C901 VP.n12 VSUBS 0.03274f
C902 VP.t0 VSUBS 2.53229f
C903 VP.n13 VSUBS 0.049166f
C904 VP.n14 VSUBS 0.03274f
C905 VP.t8 VSUBS 2.53229f
C906 VP.n15 VSUBS 0.061019f
C907 VP.n16 VSUBS 0.03274f
C908 VP.t3 VSUBS 2.53229f
C909 VP.n17 VSUBS 0.993131f
C910 VP.t1 VSUBS 2.73434f
C911 VP.n18 VSUBS 0.966386f
C912 VP.n19 VSUBS 0.276506f
C913 VP.n20 VSUBS 0.059212f
C914 VP.n21 VSUBS 0.049166f
C915 VP.n22 VSUBS 0.046429f
C916 VP.n23 VSUBS 0.03274f
C917 VP.n24 VSUBS 0.03274f
C918 VP.n25 VSUBS 0.03274f
C919 VP.n26 VSUBS 0.926932f
C920 VP.n27 VSUBS 0.061019f
C921 VP.n28 VSUBS 0.046429f
C922 VP.n29 VSUBS 0.03274f
C923 VP.n30 VSUBS 0.03274f
C924 VP.n31 VSUBS 0.03274f
C925 VP.n32 VSUBS 0.059212f
C926 VP.n33 VSUBS 0.896039f
C927 VP.n34 VSUBS 0.032701f
C928 VP.n35 VSUBS 0.061019f
C929 VP.n36 VSUBS 0.03274f
C930 VP.n37 VSUBS 0.03274f
C931 VP.n38 VSUBS 0.03274f
C932 VP.n39 VSUBS 0.051903f
C933 VP.n40 VSUBS 0.057404f
C934 VP.n41 VSUBS 1.00696f
C935 VP.n42 VSUBS 1.89473f
C936 VP.n43 VSUBS 1.91752f
C937 VP.t7 VSUBS 2.53229f
C938 VP.n44 VSUBS 1.00696f
C939 VP.n45 VSUBS 0.057404f
C940 VP.n46 VSUBS 0.043165f
C941 VP.n47 VSUBS 0.03274f
C942 VP.n48 VSUBS 0.03274f
C943 VP.n49 VSUBS 0.043692f
C944 VP.n50 VSUBS 0.061019f
C945 VP.n51 VSUBS 0.032701f
C946 VP.n52 VSUBS 0.03274f
C947 VP.n53 VSUBS 0.03274f
C948 VP.n54 VSUBS 0.059212f
C949 VP.n55 VSUBS 0.049166f
C950 VP.n56 VSUBS 0.046429f
C951 VP.n57 VSUBS 0.03274f
C952 VP.n58 VSUBS 0.03274f
C953 VP.n59 VSUBS 0.03274f
C954 VP.n60 VSUBS 0.926932f
C955 VP.n61 VSUBS 0.061019f
C956 VP.n62 VSUBS 0.046429f
C957 VP.n63 VSUBS 0.03274f
C958 VP.n64 VSUBS 0.03274f
C959 VP.n65 VSUBS 0.03274f
C960 VP.n66 VSUBS 0.059212f
C961 VP.n67 VSUBS 0.896039f
C962 VP.n68 VSUBS 0.032701f
C963 VP.n69 VSUBS 0.061019f
C964 VP.n70 VSUBS 0.03274f
C965 VP.n71 VSUBS 0.03274f
C966 VP.n72 VSUBS 0.03274f
C967 VP.n73 VSUBS 0.051903f
C968 VP.n74 VSUBS 0.057404f
C969 VP.n75 VSUBS 1.00696f
C970 VP.n76 VSUBS 0.038639f
C971 VDD2.t9 VSUBS 2.98181f
C972 VDD2.t6 VSUBS 0.285985f
C973 VDD2.t0 VSUBS 0.285985f
C974 VDD2.n0 VSUBS 2.26941f
C975 VDD2.n1 VSUBS 1.54008f
C976 VDD2.t7 VSUBS 0.285985f
C977 VDD2.t3 VSUBS 0.285985f
C978 VDD2.n2 VSUBS 2.28707f
C979 VDD2.n3 VSUBS 3.29085f
C980 VDD2.t8 VSUBS 2.95965f
C981 VDD2.n4 VSUBS 3.63992f
C982 VDD2.t2 VSUBS 0.285985f
C983 VDD2.t4 VSUBS 0.285985f
C984 VDD2.n5 VSUBS 2.26941f
C985 VDD2.n6 VSUBS 0.761113f
C986 VDD2.t1 VSUBS 0.285985f
C987 VDD2.t5 VSUBS 0.285985f
C988 VDD2.n7 VSUBS 2.28702f
C989 VTAIL.t14 VSUBS 0.294318f
C990 VTAIL.t9 VSUBS 0.294318f
C991 VTAIL.n0 VSUBS 2.17882f
C992 VTAIL.n1 VSUBS 0.94436f
C993 VTAIL.t0 VSUBS 2.86959f
C994 VTAIL.n2 VSUBS 1.09929f
C995 VTAIL.t4 VSUBS 0.294318f
C996 VTAIL.t18 VSUBS 0.294318f
C997 VTAIL.n3 VSUBS 2.17882f
C998 VTAIL.n4 VSUBS 1.04133f
C999 VTAIL.t3 VSUBS 0.294318f
C1000 VTAIL.t19 VSUBS 0.294318f
C1001 VTAIL.n5 VSUBS 2.17882f
C1002 VTAIL.n6 VSUBS 2.65146f
C1003 VTAIL.t7 VSUBS 0.294318f
C1004 VTAIL.t11 VSUBS 0.294318f
C1005 VTAIL.n7 VSUBS 2.17883f
C1006 VTAIL.n8 VSUBS 2.65145f
C1007 VTAIL.t5 VSUBS 0.294318f
C1008 VTAIL.t10 VSUBS 0.294318f
C1009 VTAIL.n9 VSUBS 2.17883f
C1010 VTAIL.n10 VSUBS 1.04132f
C1011 VTAIL.t8 VSUBS 2.8696f
C1012 VTAIL.n11 VSUBS 1.09928f
C1013 VTAIL.t16 VSUBS 0.294318f
C1014 VTAIL.t15 VSUBS 0.294318f
C1015 VTAIL.n12 VSUBS 2.17883f
C1016 VTAIL.n13 VSUBS 0.987365f
C1017 VTAIL.t1 VSUBS 0.294318f
C1018 VTAIL.t2 VSUBS 0.294318f
C1019 VTAIL.n14 VSUBS 2.17883f
C1020 VTAIL.n15 VSUBS 1.04132f
C1021 VTAIL.t17 VSUBS 2.86959f
C1022 VTAIL.n16 VSUBS 2.57022f
C1023 VTAIL.t6 VSUBS 2.86959f
C1024 VTAIL.n17 VSUBS 2.57022f
C1025 VTAIL.t13 VSUBS 0.294318f
C1026 VTAIL.t12 VSUBS 0.294318f
C1027 VTAIL.n18 VSUBS 2.17882f
C1028 VTAIL.n19 VSUBS 0.891185f
C1029 VN.n0 VSUBS 0.040133f
C1030 VN.t6 VSUBS 2.35444f
C1031 VN.n1 VSUBS 0.040624f
C1032 VN.n2 VSUBS 0.030441f
C1033 VN.t2 VSUBS 2.35444f
C1034 VN.n3 VSUBS 0.045713f
C1035 VN.n4 VSUBS 0.030441f
C1036 VN.t9 VSUBS 2.35444f
C1037 VN.n5 VSUBS 0.056734f
C1038 VN.n6 VSUBS 0.030441f
C1039 VN.t3 VSUBS 2.35444f
C1040 VN.n7 VSUBS 0.92338f
C1041 VN.t0 VSUBS 2.5423f
C1042 VN.n8 VSUBS 0.898513f
C1043 VN.n9 VSUBS 0.257086f
C1044 VN.n10 VSUBS 0.055053f
C1045 VN.n11 VSUBS 0.045713f
C1046 VN.n12 VSUBS 0.043168f
C1047 VN.n13 VSUBS 0.030441f
C1048 VN.n14 VSUBS 0.030441f
C1049 VN.n15 VSUBS 0.030441f
C1050 VN.n16 VSUBS 0.861831f
C1051 VN.n17 VSUBS 0.056734f
C1052 VN.n18 VSUBS 0.043168f
C1053 VN.n19 VSUBS 0.030441f
C1054 VN.n20 VSUBS 0.030441f
C1055 VN.n21 VSUBS 0.030441f
C1056 VN.n22 VSUBS 0.055053f
C1057 VN.n23 VSUBS 0.833107f
C1058 VN.n24 VSUBS 0.030405f
C1059 VN.n25 VSUBS 0.056734f
C1060 VN.n26 VSUBS 0.030441f
C1061 VN.n27 VSUBS 0.030441f
C1062 VN.n28 VSUBS 0.030441f
C1063 VN.n29 VSUBS 0.048258f
C1064 VN.n30 VSUBS 0.053373f
C1065 VN.n31 VSUBS 0.936238f
C1066 VN.n32 VSUBS 0.035925f
C1067 VN.n33 VSUBS 0.040133f
C1068 VN.t1 VSUBS 2.35444f
C1069 VN.n34 VSUBS 0.040624f
C1070 VN.n35 VSUBS 0.030441f
C1071 VN.t7 VSUBS 2.35444f
C1072 VN.n36 VSUBS 0.045713f
C1073 VN.n37 VSUBS 0.030441f
C1074 VN.t5 VSUBS 2.35444f
C1075 VN.n38 VSUBS 0.056734f
C1076 VN.n39 VSUBS 0.030441f
C1077 VN.t8 VSUBS 2.35444f
C1078 VN.n40 VSUBS 0.92338f
C1079 VN.t4 VSUBS 2.5423f
C1080 VN.n41 VSUBS 0.898513f
C1081 VN.n42 VSUBS 0.257086f
C1082 VN.n43 VSUBS 0.055053f
C1083 VN.n44 VSUBS 0.045713f
C1084 VN.n45 VSUBS 0.043168f
C1085 VN.n46 VSUBS 0.030441f
C1086 VN.n47 VSUBS 0.030441f
C1087 VN.n48 VSUBS 0.030441f
C1088 VN.n49 VSUBS 0.861831f
C1089 VN.n50 VSUBS 0.056734f
C1090 VN.n51 VSUBS 0.043168f
C1091 VN.n52 VSUBS 0.030441f
C1092 VN.n53 VSUBS 0.030441f
C1093 VN.n54 VSUBS 0.030441f
C1094 VN.n55 VSUBS 0.055053f
C1095 VN.n56 VSUBS 0.833107f
C1096 VN.n57 VSUBS 0.030405f
C1097 VN.n58 VSUBS 0.056734f
C1098 VN.n59 VSUBS 0.030441f
C1099 VN.n60 VSUBS 0.030441f
C1100 VN.n61 VSUBS 0.030441f
C1101 VN.n62 VSUBS 0.048258f
C1102 VN.n63 VSUBS 0.053373f
C1103 VN.n64 VSUBS 0.936238f
C1104 VN.n65 VSUBS 1.77793f
.ends

