* NGSPICE file created from diff_pair_sample_0793.ext - technology: sky130A

.subckt diff_pair_sample_0793 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X1 VTAIL.t6 VP.t0 VDD1.t9 B.t20 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X2 VTAIL.t18 VN.t1 VDD2.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X3 B.t18 B.t16 B.t17 B.t10 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=0 ps=0 w=14.31 l=2.34
X4 VDD1.t8 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=5.5809 ps=29.4 w=14.31 l=2.34
X5 VDD1.t7 VP.t2 VTAIL.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X6 VTAIL.t17 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X7 VDD1.t6 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=5.5809 ps=29.4 w=14.31 l=2.34
X8 VTAIL.t16 VN.t3 VDD2.t0 B.t20 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X9 B.t15 B.t13 B.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=0 ps=0 w=14.31 l=2.34
X10 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=0 ps=0 w=14.31 l=2.34
X11 VDD1.t5 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X12 VDD1.t4 VP.t5 VTAIL.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=2.36115 ps=14.64 w=14.31 l=2.34
X13 VDD2.t9 VN.t4 VTAIL.t15 B.t22 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=2.36115 ps=14.64 w=14.31 l=2.34
X14 VDD1.t3 VP.t6 VTAIL.t8 B.t22 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=2.36115 ps=14.64 w=14.31 l=2.34
X15 VDD2.t8 VN.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=5.5809 ps=29.4 w=14.31 l=2.34
X16 VTAIL.t3 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X17 VDD2.t5 VN.t6 VTAIL.t13 B.t19 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X18 VDD2.t4 VN.t7 VTAIL.t12 B.t23 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=2.36115 ps=14.64 w=14.31 l=2.34
X19 VTAIL.t2 VP.t8 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X20 VDD2.t7 VN.t8 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
X21 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.5809 pd=29.4 as=0 ps=0 w=14.31 l=2.34
X22 VDD2.t6 VN.t9 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=5.5809 ps=29.4 w=14.31 l=2.34
X23 VTAIL.t7 VP.t9 VDD1.t0 B.t21 sky130_fd_pr__nfet_01v8 ad=2.36115 pd=14.64 as=2.36115 ps=14.64 w=14.31 l=2.34
R0 VN.n8 VN.t7 180.448
R1 VN.n45 VN.t5 180.448
R2 VN.n71 VN.n37 161.3
R3 VN.n70 VN.n69 161.3
R4 VN.n68 VN.n38 161.3
R5 VN.n67 VN.n66 161.3
R6 VN.n65 VN.n39 161.3
R7 VN.n63 VN.n62 161.3
R8 VN.n61 VN.n40 161.3
R9 VN.n60 VN.n59 161.3
R10 VN.n58 VN.n41 161.3
R11 VN.n57 VN.n56 161.3
R12 VN.n55 VN.n42 161.3
R13 VN.n54 VN.n53 161.3
R14 VN.n52 VN.n43 161.3
R15 VN.n51 VN.n50 161.3
R16 VN.n49 VN.n44 161.3
R17 VN.n48 VN.n47 161.3
R18 VN.n34 VN.n0 161.3
R19 VN.n33 VN.n32 161.3
R20 VN.n31 VN.n1 161.3
R21 VN.n30 VN.n29 161.3
R22 VN.n28 VN.n2 161.3
R23 VN.n26 VN.n25 161.3
R24 VN.n24 VN.n3 161.3
R25 VN.n23 VN.n22 161.3
R26 VN.n21 VN.n4 161.3
R27 VN.n20 VN.n19 161.3
R28 VN.n18 VN.n5 161.3
R29 VN.n17 VN.n16 161.3
R30 VN.n15 VN.n6 161.3
R31 VN.n14 VN.n13 161.3
R32 VN.n12 VN.n7 161.3
R33 VN.n11 VN.n10 161.3
R34 VN.n5 VN.t6 147.381
R35 VN.n9 VN.t0 147.381
R36 VN.n27 VN.t2 147.381
R37 VN.n35 VN.t9 147.381
R38 VN.n42 VN.t8 147.381
R39 VN.n46 VN.t1 147.381
R40 VN.n64 VN.t3 147.381
R41 VN.n72 VN.t4 147.381
R42 VN.n36 VN.n35 94.1189
R43 VN.n73 VN.n72 94.1189
R44 VN.n9 VN.n8 63.5395
R45 VN.n46 VN.n45 63.5395
R46 VN.n15 VN.n14 56.5193
R47 VN.n22 VN.n21 56.5193
R48 VN.n52 VN.n51 56.5193
R49 VN.n59 VN.n58 56.5193
R50 VN VN.n73 53.7898
R51 VN.n33 VN.n1 40.979
R52 VN.n70 VN.n38 40.979
R53 VN.n29 VN.n1 40.0078
R54 VN.n66 VN.n38 40.0078
R55 VN.n10 VN.n7 24.4675
R56 VN.n14 VN.n7 24.4675
R57 VN.n16 VN.n15 24.4675
R58 VN.n16 VN.n5 24.4675
R59 VN.n20 VN.n5 24.4675
R60 VN.n21 VN.n20 24.4675
R61 VN.n22 VN.n3 24.4675
R62 VN.n26 VN.n3 24.4675
R63 VN.n29 VN.n28 24.4675
R64 VN.n34 VN.n33 24.4675
R65 VN.n51 VN.n44 24.4675
R66 VN.n47 VN.n44 24.4675
R67 VN.n58 VN.n57 24.4675
R68 VN.n57 VN.n42 24.4675
R69 VN.n53 VN.n42 24.4675
R70 VN.n53 VN.n52 24.4675
R71 VN.n66 VN.n65 24.4675
R72 VN.n63 VN.n40 24.4675
R73 VN.n59 VN.n40 24.4675
R74 VN.n71 VN.n70 24.4675
R75 VN.n35 VN.n34 16.6381
R76 VN.n72 VN.n71 16.6381
R77 VN.n28 VN.n27 16.1487
R78 VN.n65 VN.n64 16.1487
R79 VN.n48 VN.n45 9.31187
R80 VN.n11 VN.n8 9.31187
R81 VN.n10 VN.n9 8.31928
R82 VN.n27 VN.n26 8.31928
R83 VN.n47 VN.n46 8.31928
R84 VN.n64 VN.n63 8.31928
R85 VN.n73 VN.n37 0.278367
R86 VN.n36 VN.n0 0.278367
R87 VN.n69 VN.n37 0.189894
R88 VN.n69 VN.n68 0.189894
R89 VN.n68 VN.n67 0.189894
R90 VN.n67 VN.n39 0.189894
R91 VN.n62 VN.n39 0.189894
R92 VN.n62 VN.n61 0.189894
R93 VN.n61 VN.n60 0.189894
R94 VN.n60 VN.n41 0.189894
R95 VN.n56 VN.n41 0.189894
R96 VN.n56 VN.n55 0.189894
R97 VN.n55 VN.n54 0.189894
R98 VN.n54 VN.n43 0.189894
R99 VN.n50 VN.n43 0.189894
R100 VN.n50 VN.n49 0.189894
R101 VN.n49 VN.n48 0.189894
R102 VN.n12 VN.n11 0.189894
R103 VN.n13 VN.n12 0.189894
R104 VN.n13 VN.n6 0.189894
R105 VN.n17 VN.n6 0.189894
R106 VN.n18 VN.n17 0.189894
R107 VN.n19 VN.n18 0.189894
R108 VN.n19 VN.n4 0.189894
R109 VN.n23 VN.n4 0.189894
R110 VN.n24 VN.n23 0.189894
R111 VN.n25 VN.n24 0.189894
R112 VN.n25 VN.n2 0.189894
R113 VN.n30 VN.n2 0.189894
R114 VN.n31 VN.n30 0.189894
R115 VN.n32 VN.n31 0.189894
R116 VN.n32 VN.n0 0.189894
R117 VN VN.n36 0.153454
R118 VDD2.n1 VDD2.t4 65.2329
R119 VDD2.n3 VDD2.n2 63.2184
R120 VDD2 VDD2.n7 63.2156
R121 VDD2.n4 VDD2.t9 62.9313
R122 VDD2.n6 VDD2.n5 61.5477
R123 VDD2.n1 VDD2.n0 61.5475
R124 VDD2.n4 VDD2.n3 46.9847
R125 VDD2.n6 VDD2.n4 2.30222
R126 VDD2.n7 VDD2.t2 1.38415
R127 VDD2.n7 VDD2.t8 1.38415
R128 VDD2.n5 VDD2.t0 1.38415
R129 VDD2.n5 VDD2.t7 1.38415
R130 VDD2.n2 VDD2.t1 1.38415
R131 VDD2.n2 VDD2.t6 1.38415
R132 VDD2.n0 VDD2.t3 1.38415
R133 VDD2.n0 VDD2.t5 1.38415
R134 VDD2 VDD2.n6 0.634121
R135 VDD2.n3 VDD2.n1 0.520585
R136 VTAIL.n11 VTAIL.t14 46.2525
R137 VTAIL.n17 VTAIL.t10 46.2524
R138 VTAIL.n2 VTAIL.t1 46.2524
R139 VTAIL.n16 VTAIL.t0 46.2524
R140 VTAIL.n15 VTAIL.n14 44.8689
R141 VTAIL.n13 VTAIL.n12 44.8689
R142 VTAIL.n10 VTAIL.n9 44.8689
R143 VTAIL.n8 VTAIL.n7 44.8689
R144 VTAIL.n19 VTAIL.n18 44.8687
R145 VTAIL.n1 VTAIL.n0 44.8687
R146 VTAIL.n4 VTAIL.n3 44.8687
R147 VTAIL.n6 VTAIL.n5 44.8687
R148 VTAIL.n8 VTAIL.n6 29.3065
R149 VTAIL.n17 VTAIL.n16 27.0048
R150 VTAIL.n10 VTAIL.n8 2.30222
R151 VTAIL.n11 VTAIL.n10 2.30222
R152 VTAIL.n15 VTAIL.n13 2.30222
R153 VTAIL.n16 VTAIL.n15 2.30222
R154 VTAIL.n6 VTAIL.n4 2.30222
R155 VTAIL.n4 VTAIL.n2 2.30222
R156 VTAIL.n19 VTAIL.n17 2.30222
R157 VTAIL VTAIL.n1 1.78498
R158 VTAIL.n13 VTAIL.n11 1.62119
R159 VTAIL.n2 VTAIL.n1 1.62119
R160 VTAIL.n18 VTAIL.t13 1.38415
R161 VTAIL.n18 VTAIL.t17 1.38415
R162 VTAIL.n0 VTAIL.t12 1.38415
R163 VTAIL.n0 VTAIL.t19 1.38415
R164 VTAIL.n3 VTAIL.t4 1.38415
R165 VTAIL.n3 VTAIL.t7 1.38415
R166 VTAIL.n5 VTAIL.t8 1.38415
R167 VTAIL.n5 VTAIL.t6 1.38415
R168 VTAIL.n14 VTAIL.t5 1.38415
R169 VTAIL.n14 VTAIL.t3 1.38415
R170 VTAIL.n12 VTAIL.t9 1.38415
R171 VTAIL.n12 VTAIL.t2 1.38415
R172 VTAIL.n9 VTAIL.t11 1.38415
R173 VTAIL.n9 VTAIL.t18 1.38415
R174 VTAIL.n7 VTAIL.t15 1.38415
R175 VTAIL.n7 VTAIL.t16 1.38415
R176 VTAIL VTAIL.n19 0.517741
R177 B.n979 B.n978 585
R178 B.n366 B.n154 585
R179 B.n365 B.n364 585
R180 B.n363 B.n362 585
R181 B.n361 B.n360 585
R182 B.n359 B.n358 585
R183 B.n357 B.n356 585
R184 B.n355 B.n354 585
R185 B.n353 B.n352 585
R186 B.n351 B.n350 585
R187 B.n349 B.n348 585
R188 B.n347 B.n346 585
R189 B.n345 B.n344 585
R190 B.n343 B.n342 585
R191 B.n341 B.n340 585
R192 B.n339 B.n338 585
R193 B.n337 B.n336 585
R194 B.n335 B.n334 585
R195 B.n333 B.n332 585
R196 B.n331 B.n330 585
R197 B.n329 B.n328 585
R198 B.n327 B.n326 585
R199 B.n325 B.n324 585
R200 B.n323 B.n322 585
R201 B.n321 B.n320 585
R202 B.n319 B.n318 585
R203 B.n317 B.n316 585
R204 B.n315 B.n314 585
R205 B.n313 B.n312 585
R206 B.n311 B.n310 585
R207 B.n309 B.n308 585
R208 B.n307 B.n306 585
R209 B.n305 B.n304 585
R210 B.n303 B.n302 585
R211 B.n301 B.n300 585
R212 B.n299 B.n298 585
R213 B.n297 B.n296 585
R214 B.n295 B.n294 585
R215 B.n293 B.n292 585
R216 B.n291 B.n290 585
R217 B.n289 B.n288 585
R218 B.n287 B.n286 585
R219 B.n285 B.n284 585
R220 B.n283 B.n282 585
R221 B.n281 B.n280 585
R222 B.n279 B.n278 585
R223 B.n277 B.n276 585
R224 B.n275 B.n274 585
R225 B.n273 B.n272 585
R226 B.n271 B.n270 585
R227 B.n269 B.n268 585
R228 B.n267 B.n266 585
R229 B.n265 B.n264 585
R230 B.n263 B.n262 585
R231 B.n261 B.n260 585
R232 B.n259 B.n258 585
R233 B.n257 B.n256 585
R234 B.n255 B.n254 585
R235 B.n253 B.n252 585
R236 B.n251 B.n250 585
R237 B.n249 B.n248 585
R238 B.n247 B.n246 585
R239 B.n245 B.n244 585
R240 B.n243 B.n242 585
R241 B.n241 B.n240 585
R242 B.n239 B.n238 585
R243 B.n237 B.n236 585
R244 B.n235 B.n234 585
R245 B.n233 B.n232 585
R246 B.n231 B.n230 585
R247 B.n229 B.n228 585
R248 B.n227 B.n226 585
R249 B.n225 B.n224 585
R250 B.n223 B.n222 585
R251 B.n221 B.n220 585
R252 B.n219 B.n218 585
R253 B.n217 B.n216 585
R254 B.n215 B.n214 585
R255 B.n213 B.n212 585
R256 B.n211 B.n210 585
R257 B.n209 B.n208 585
R258 B.n207 B.n206 585
R259 B.n205 B.n204 585
R260 B.n203 B.n202 585
R261 B.n201 B.n200 585
R262 B.n199 B.n198 585
R263 B.n197 B.n196 585
R264 B.n195 B.n194 585
R265 B.n193 B.n192 585
R266 B.n191 B.n190 585
R267 B.n189 B.n188 585
R268 B.n187 B.n186 585
R269 B.n185 B.n184 585
R270 B.n183 B.n182 585
R271 B.n181 B.n180 585
R272 B.n179 B.n178 585
R273 B.n177 B.n176 585
R274 B.n175 B.n174 585
R275 B.n173 B.n172 585
R276 B.n171 B.n170 585
R277 B.n169 B.n168 585
R278 B.n167 B.n166 585
R279 B.n165 B.n164 585
R280 B.n163 B.n162 585
R281 B.n102 B.n101 585
R282 B.n984 B.n983 585
R283 B.n977 B.n155 585
R284 B.n155 B.n99 585
R285 B.n976 B.n98 585
R286 B.n988 B.n98 585
R287 B.n975 B.n97 585
R288 B.n989 B.n97 585
R289 B.n974 B.n96 585
R290 B.n990 B.n96 585
R291 B.n973 B.n972 585
R292 B.n972 B.n92 585
R293 B.n971 B.n91 585
R294 B.n996 B.n91 585
R295 B.n970 B.n90 585
R296 B.n997 B.n90 585
R297 B.n969 B.n89 585
R298 B.t6 B.n89 585
R299 B.n968 B.n967 585
R300 B.n967 B.n85 585
R301 B.n966 B.n84 585
R302 B.n1003 B.n84 585
R303 B.n965 B.n83 585
R304 B.n1004 B.n83 585
R305 B.n964 B.n82 585
R306 B.n1005 B.n82 585
R307 B.n963 B.n962 585
R308 B.n962 B.n78 585
R309 B.n961 B.n77 585
R310 B.n1011 B.n77 585
R311 B.n960 B.n76 585
R312 B.n1012 B.n76 585
R313 B.n959 B.n75 585
R314 B.n1013 B.n75 585
R315 B.n958 B.n957 585
R316 B.n957 B.n71 585
R317 B.n956 B.n70 585
R318 B.n1019 B.n70 585
R319 B.n955 B.n69 585
R320 B.n1020 B.n69 585
R321 B.n954 B.n68 585
R322 B.n1021 B.n68 585
R323 B.n953 B.n952 585
R324 B.n952 B.n64 585
R325 B.n951 B.n63 585
R326 B.n1027 B.n63 585
R327 B.n950 B.n62 585
R328 B.n1028 B.n62 585
R329 B.n949 B.n61 585
R330 B.n1029 B.n61 585
R331 B.n948 B.n947 585
R332 B.n947 B.n57 585
R333 B.n946 B.n56 585
R334 B.n1035 B.n56 585
R335 B.n945 B.n55 585
R336 B.n1036 B.n55 585
R337 B.n944 B.n54 585
R338 B.n1037 B.n54 585
R339 B.n943 B.n942 585
R340 B.n942 B.n50 585
R341 B.n941 B.n49 585
R342 B.n1043 B.n49 585
R343 B.n940 B.n48 585
R344 B.n1044 B.n48 585
R345 B.n939 B.n47 585
R346 B.n1045 B.n47 585
R347 B.n938 B.n937 585
R348 B.n937 B.n43 585
R349 B.n936 B.n42 585
R350 B.n1051 B.n42 585
R351 B.n935 B.n41 585
R352 B.n1052 B.n41 585
R353 B.n934 B.n40 585
R354 B.n1053 B.n40 585
R355 B.n933 B.n932 585
R356 B.n932 B.n36 585
R357 B.n931 B.n35 585
R358 B.n1059 B.n35 585
R359 B.n930 B.n34 585
R360 B.n1060 B.n34 585
R361 B.n929 B.n33 585
R362 B.n1061 B.n33 585
R363 B.n928 B.n927 585
R364 B.n927 B.n29 585
R365 B.n926 B.n28 585
R366 B.n1067 B.n28 585
R367 B.n925 B.n27 585
R368 B.n1068 B.n27 585
R369 B.n924 B.n26 585
R370 B.n1069 B.n26 585
R371 B.n923 B.n922 585
R372 B.n922 B.n22 585
R373 B.n921 B.n21 585
R374 B.n1075 B.n21 585
R375 B.n920 B.n20 585
R376 B.n1076 B.n20 585
R377 B.n919 B.n19 585
R378 B.n1077 B.n19 585
R379 B.n918 B.n917 585
R380 B.n917 B.n15 585
R381 B.n916 B.n14 585
R382 B.n1083 B.n14 585
R383 B.n915 B.n13 585
R384 B.n1084 B.n13 585
R385 B.n914 B.n12 585
R386 B.n1085 B.n12 585
R387 B.n913 B.n912 585
R388 B.n912 B.n8 585
R389 B.n911 B.n7 585
R390 B.n1091 B.n7 585
R391 B.n910 B.n6 585
R392 B.n1092 B.n6 585
R393 B.n909 B.n5 585
R394 B.n1093 B.n5 585
R395 B.n908 B.n907 585
R396 B.n907 B.n4 585
R397 B.n906 B.n367 585
R398 B.n906 B.n905 585
R399 B.n896 B.n368 585
R400 B.n369 B.n368 585
R401 B.n898 B.n897 585
R402 B.n899 B.n898 585
R403 B.n895 B.n374 585
R404 B.n374 B.n373 585
R405 B.n894 B.n893 585
R406 B.n893 B.n892 585
R407 B.n376 B.n375 585
R408 B.n377 B.n376 585
R409 B.n885 B.n884 585
R410 B.n886 B.n885 585
R411 B.n883 B.n382 585
R412 B.n382 B.n381 585
R413 B.n882 B.n881 585
R414 B.n881 B.n880 585
R415 B.n384 B.n383 585
R416 B.n385 B.n384 585
R417 B.n873 B.n872 585
R418 B.n874 B.n873 585
R419 B.n871 B.n390 585
R420 B.n390 B.n389 585
R421 B.n870 B.n869 585
R422 B.n869 B.n868 585
R423 B.n392 B.n391 585
R424 B.n393 B.n392 585
R425 B.n861 B.n860 585
R426 B.n862 B.n861 585
R427 B.n859 B.n398 585
R428 B.n398 B.n397 585
R429 B.n858 B.n857 585
R430 B.n857 B.n856 585
R431 B.n400 B.n399 585
R432 B.n401 B.n400 585
R433 B.n849 B.n848 585
R434 B.n850 B.n849 585
R435 B.n847 B.n406 585
R436 B.n406 B.n405 585
R437 B.n846 B.n845 585
R438 B.n845 B.n844 585
R439 B.n408 B.n407 585
R440 B.n409 B.n408 585
R441 B.n837 B.n836 585
R442 B.n838 B.n837 585
R443 B.n835 B.n414 585
R444 B.n414 B.n413 585
R445 B.n834 B.n833 585
R446 B.n833 B.n832 585
R447 B.n416 B.n415 585
R448 B.n417 B.n416 585
R449 B.n825 B.n824 585
R450 B.n826 B.n825 585
R451 B.n823 B.n422 585
R452 B.n422 B.n421 585
R453 B.n822 B.n821 585
R454 B.n821 B.n820 585
R455 B.n424 B.n423 585
R456 B.n425 B.n424 585
R457 B.n813 B.n812 585
R458 B.n814 B.n813 585
R459 B.n811 B.n430 585
R460 B.n430 B.n429 585
R461 B.n810 B.n809 585
R462 B.n809 B.n808 585
R463 B.n432 B.n431 585
R464 B.n433 B.n432 585
R465 B.n801 B.n800 585
R466 B.n802 B.n801 585
R467 B.n799 B.n437 585
R468 B.n441 B.n437 585
R469 B.n798 B.n797 585
R470 B.n797 B.n796 585
R471 B.n439 B.n438 585
R472 B.n440 B.n439 585
R473 B.n789 B.n788 585
R474 B.n790 B.n789 585
R475 B.n787 B.n446 585
R476 B.n446 B.n445 585
R477 B.n786 B.n785 585
R478 B.n785 B.n784 585
R479 B.n448 B.n447 585
R480 B.n449 B.n448 585
R481 B.n777 B.n776 585
R482 B.n778 B.n777 585
R483 B.n775 B.n454 585
R484 B.n454 B.n453 585
R485 B.n774 B.n773 585
R486 B.n773 B.n772 585
R487 B.n456 B.n455 585
R488 B.n457 B.n456 585
R489 B.n766 B.n765 585
R490 B.t10 B.n766 585
R491 B.n764 B.n462 585
R492 B.n462 B.n461 585
R493 B.n763 B.n762 585
R494 B.n762 B.n761 585
R495 B.n464 B.n463 585
R496 B.n465 B.n464 585
R497 B.n754 B.n753 585
R498 B.n755 B.n754 585
R499 B.n752 B.n470 585
R500 B.n470 B.n469 585
R501 B.n751 B.n750 585
R502 B.n750 B.n749 585
R503 B.n472 B.n471 585
R504 B.n473 B.n472 585
R505 B.n745 B.n744 585
R506 B.n476 B.n475 585
R507 B.n741 B.n740 585
R508 B.n742 B.n741 585
R509 B.n739 B.n529 585
R510 B.n738 B.n737 585
R511 B.n736 B.n735 585
R512 B.n734 B.n733 585
R513 B.n732 B.n731 585
R514 B.n730 B.n729 585
R515 B.n728 B.n727 585
R516 B.n726 B.n725 585
R517 B.n724 B.n723 585
R518 B.n722 B.n721 585
R519 B.n720 B.n719 585
R520 B.n718 B.n717 585
R521 B.n716 B.n715 585
R522 B.n714 B.n713 585
R523 B.n712 B.n711 585
R524 B.n710 B.n709 585
R525 B.n708 B.n707 585
R526 B.n706 B.n705 585
R527 B.n704 B.n703 585
R528 B.n702 B.n701 585
R529 B.n700 B.n699 585
R530 B.n698 B.n697 585
R531 B.n696 B.n695 585
R532 B.n694 B.n693 585
R533 B.n692 B.n691 585
R534 B.n690 B.n689 585
R535 B.n688 B.n687 585
R536 B.n686 B.n685 585
R537 B.n684 B.n683 585
R538 B.n682 B.n681 585
R539 B.n680 B.n679 585
R540 B.n678 B.n677 585
R541 B.n676 B.n675 585
R542 B.n674 B.n673 585
R543 B.n672 B.n671 585
R544 B.n670 B.n669 585
R545 B.n668 B.n667 585
R546 B.n666 B.n665 585
R547 B.n664 B.n663 585
R548 B.n662 B.n661 585
R549 B.n660 B.n659 585
R550 B.n658 B.n657 585
R551 B.n656 B.n655 585
R552 B.n654 B.n653 585
R553 B.n652 B.n651 585
R554 B.n649 B.n648 585
R555 B.n647 B.n646 585
R556 B.n645 B.n644 585
R557 B.n643 B.n642 585
R558 B.n641 B.n640 585
R559 B.n639 B.n638 585
R560 B.n637 B.n636 585
R561 B.n635 B.n634 585
R562 B.n633 B.n632 585
R563 B.n631 B.n630 585
R564 B.n628 B.n627 585
R565 B.n626 B.n625 585
R566 B.n624 B.n623 585
R567 B.n622 B.n621 585
R568 B.n620 B.n619 585
R569 B.n618 B.n617 585
R570 B.n616 B.n615 585
R571 B.n614 B.n613 585
R572 B.n612 B.n611 585
R573 B.n610 B.n609 585
R574 B.n608 B.n607 585
R575 B.n606 B.n605 585
R576 B.n604 B.n603 585
R577 B.n602 B.n601 585
R578 B.n600 B.n599 585
R579 B.n598 B.n597 585
R580 B.n596 B.n595 585
R581 B.n594 B.n593 585
R582 B.n592 B.n591 585
R583 B.n590 B.n589 585
R584 B.n588 B.n587 585
R585 B.n586 B.n585 585
R586 B.n584 B.n583 585
R587 B.n582 B.n581 585
R588 B.n580 B.n579 585
R589 B.n578 B.n577 585
R590 B.n576 B.n575 585
R591 B.n574 B.n573 585
R592 B.n572 B.n571 585
R593 B.n570 B.n569 585
R594 B.n568 B.n567 585
R595 B.n566 B.n565 585
R596 B.n564 B.n563 585
R597 B.n562 B.n561 585
R598 B.n560 B.n559 585
R599 B.n558 B.n557 585
R600 B.n556 B.n555 585
R601 B.n554 B.n553 585
R602 B.n552 B.n551 585
R603 B.n550 B.n549 585
R604 B.n548 B.n547 585
R605 B.n546 B.n545 585
R606 B.n544 B.n543 585
R607 B.n542 B.n541 585
R608 B.n540 B.n539 585
R609 B.n538 B.n537 585
R610 B.n536 B.n535 585
R611 B.n534 B.n528 585
R612 B.n742 B.n528 585
R613 B.n746 B.n474 585
R614 B.n474 B.n473 585
R615 B.n748 B.n747 585
R616 B.n749 B.n748 585
R617 B.n468 B.n467 585
R618 B.n469 B.n468 585
R619 B.n757 B.n756 585
R620 B.n756 B.n755 585
R621 B.n758 B.n466 585
R622 B.n466 B.n465 585
R623 B.n760 B.n759 585
R624 B.n761 B.n760 585
R625 B.n460 B.n459 585
R626 B.n461 B.n460 585
R627 B.n768 B.n767 585
R628 B.n767 B.t10 585
R629 B.n769 B.n458 585
R630 B.n458 B.n457 585
R631 B.n771 B.n770 585
R632 B.n772 B.n771 585
R633 B.n452 B.n451 585
R634 B.n453 B.n452 585
R635 B.n780 B.n779 585
R636 B.n779 B.n778 585
R637 B.n781 B.n450 585
R638 B.n450 B.n449 585
R639 B.n783 B.n782 585
R640 B.n784 B.n783 585
R641 B.n444 B.n443 585
R642 B.n445 B.n444 585
R643 B.n792 B.n791 585
R644 B.n791 B.n790 585
R645 B.n793 B.n442 585
R646 B.n442 B.n440 585
R647 B.n795 B.n794 585
R648 B.n796 B.n795 585
R649 B.n436 B.n435 585
R650 B.n441 B.n436 585
R651 B.n804 B.n803 585
R652 B.n803 B.n802 585
R653 B.n805 B.n434 585
R654 B.n434 B.n433 585
R655 B.n807 B.n806 585
R656 B.n808 B.n807 585
R657 B.n428 B.n427 585
R658 B.n429 B.n428 585
R659 B.n816 B.n815 585
R660 B.n815 B.n814 585
R661 B.n817 B.n426 585
R662 B.n426 B.n425 585
R663 B.n819 B.n818 585
R664 B.n820 B.n819 585
R665 B.n420 B.n419 585
R666 B.n421 B.n420 585
R667 B.n828 B.n827 585
R668 B.n827 B.n826 585
R669 B.n829 B.n418 585
R670 B.n418 B.n417 585
R671 B.n831 B.n830 585
R672 B.n832 B.n831 585
R673 B.n412 B.n411 585
R674 B.n413 B.n412 585
R675 B.n840 B.n839 585
R676 B.n839 B.n838 585
R677 B.n841 B.n410 585
R678 B.n410 B.n409 585
R679 B.n843 B.n842 585
R680 B.n844 B.n843 585
R681 B.n404 B.n403 585
R682 B.n405 B.n404 585
R683 B.n852 B.n851 585
R684 B.n851 B.n850 585
R685 B.n853 B.n402 585
R686 B.n402 B.n401 585
R687 B.n855 B.n854 585
R688 B.n856 B.n855 585
R689 B.n396 B.n395 585
R690 B.n397 B.n396 585
R691 B.n864 B.n863 585
R692 B.n863 B.n862 585
R693 B.n865 B.n394 585
R694 B.n394 B.n393 585
R695 B.n867 B.n866 585
R696 B.n868 B.n867 585
R697 B.n388 B.n387 585
R698 B.n389 B.n388 585
R699 B.n876 B.n875 585
R700 B.n875 B.n874 585
R701 B.n877 B.n386 585
R702 B.n386 B.n385 585
R703 B.n879 B.n878 585
R704 B.n880 B.n879 585
R705 B.n380 B.n379 585
R706 B.n381 B.n380 585
R707 B.n888 B.n887 585
R708 B.n887 B.n886 585
R709 B.n889 B.n378 585
R710 B.n378 B.n377 585
R711 B.n891 B.n890 585
R712 B.n892 B.n891 585
R713 B.n372 B.n371 585
R714 B.n373 B.n372 585
R715 B.n901 B.n900 585
R716 B.n900 B.n899 585
R717 B.n902 B.n370 585
R718 B.n370 B.n369 585
R719 B.n904 B.n903 585
R720 B.n905 B.n904 585
R721 B.n2 B.n0 585
R722 B.n4 B.n2 585
R723 B.n3 B.n1 585
R724 B.n1092 B.n3 585
R725 B.n1090 B.n1089 585
R726 B.n1091 B.n1090 585
R727 B.n1088 B.n9 585
R728 B.n9 B.n8 585
R729 B.n1087 B.n1086 585
R730 B.n1086 B.n1085 585
R731 B.n11 B.n10 585
R732 B.n1084 B.n11 585
R733 B.n1082 B.n1081 585
R734 B.n1083 B.n1082 585
R735 B.n1080 B.n16 585
R736 B.n16 B.n15 585
R737 B.n1079 B.n1078 585
R738 B.n1078 B.n1077 585
R739 B.n18 B.n17 585
R740 B.n1076 B.n18 585
R741 B.n1074 B.n1073 585
R742 B.n1075 B.n1074 585
R743 B.n1072 B.n23 585
R744 B.n23 B.n22 585
R745 B.n1071 B.n1070 585
R746 B.n1070 B.n1069 585
R747 B.n25 B.n24 585
R748 B.n1068 B.n25 585
R749 B.n1066 B.n1065 585
R750 B.n1067 B.n1066 585
R751 B.n1064 B.n30 585
R752 B.n30 B.n29 585
R753 B.n1063 B.n1062 585
R754 B.n1062 B.n1061 585
R755 B.n32 B.n31 585
R756 B.n1060 B.n32 585
R757 B.n1058 B.n1057 585
R758 B.n1059 B.n1058 585
R759 B.n1056 B.n37 585
R760 B.n37 B.n36 585
R761 B.n1055 B.n1054 585
R762 B.n1054 B.n1053 585
R763 B.n39 B.n38 585
R764 B.n1052 B.n39 585
R765 B.n1050 B.n1049 585
R766 B.n1051 B.n1050 585
R767 B.n1048 B.n44 585
R768 B.n44 B.n43 585
R769 B.n1047 B.n1046 585
R770 B.n1046 B.n1045 585
R771 B.n46 B.n45 585
R772 B.n1044 B.n46 585
R773 B.n1042 B.n1041 585
R774 B.n1043 B.n1042 585
R775 B.n1040 B.n51 585
R776 B.n51 B.n50 585
R777 B.n1039 B.n1038 585
R778 B.n1038 B.n1037 585
R779 B.n53 B.n52 585
R780 B.n1036 B.n53 585
R781 B.n1034 B.n1033 585
R782 B.n1035 B.n1034 585
R783 B.n1032 B.n58 585
R784 B.n58 B.n57 585
R785 B.n1031 B.n1030 585
R786 B.n1030 B.n1029 585
R787 B.n60 B.n59 585
R788 B.n1028 B.n60 585
R789 B.n1026 B.n1025 585
R790 B.n1027 B.n1026 585
R791 B.n1024 B.n65 585
R792 B.n65 B.n64 585
R793 B.n1023 B.n1022 585
R794 B.n1022 B.n1021 585
R795 B.n67 B.n66 585
R796 B.n1020 B.n67 585
R797 B.n1018 B.n1017 585
R798 B.n1019 B.n1018 585
R799 B.n1016 B.n72 585
R800 B.n72 B.n71 585
R801 B.n1015 B.n1014 585
R802 B.n1014 B.n1013 585
R803 B.n74 B.n73 585
R804 B.n1012 B.n74 585
R805 B.n1010 B.n1009 585
R806 B.n1011 B.n1010 585
R807 B.n1008 B.n79 585
R808 B.n79 B.n78 585
R809 B.n1007 B.n1006 585
R810 B.n1006 B.n1005 585
R811 B.n81 B.n80 585
R812 B.n1004 B.n81 585
R813 B.n1002 B.n1001 585
R814 B.n1003 B.n1002 585
R815 B.n1000 B.n86 585
R816 B.n86 B.n85 585
R817 B.n999 B.n998 585
R818 B.n998 B.t6 585
R819 B.n88 B.n87 585
R820 B.n997 B.n88 585
R821 B.n995 B.n994 585
R822 B.n996 B.n995 585
R823 B.n993 B.n93 585
R824 B.n93 B.n92 585
R825 B.n992 B.n991 585
R826 B.n991 B.n990 585
R827 B.n95 B.n94 585
R828 B.n989 B.n95 585
R829 B.n987 B.n986 585
R830 B.n988 B.n987 585
R831 B.n985 B.n100 585
R832 B.n100 B.n99 585
R833 B.n1095 B.n1094 585
R834 B.n1094 B.n1093 585
R835 B.n744 B.n474 569.379
R836 B.n983 B.n100 569.379
R837 B.n528 B.n472 569.379
R838 B.n979 B.n155 569.379
R839 B.n532 B.t16 354.998
R840 B.n530 B.t9 354.998
R841 B.n159 B.t5 354.998
R842 B.n156 B.t13 354.998
R843 B.n981 B.n980 256.663
R844 B.n981 B.n153 256.663
R845 B.n981 B.n152 256.663
R846 B.n981 B.n151 256.663
R847 B.n981 B.n150 256.663
R848 B.n981 B.n149 256.663
R849 B.n981 B.n148 256.663
R850 B.n981 B.n147 256.663
R851 B.n981 B.n146 256.663
R852 B.n981 B.n145 256.663
R853 B.n981 B.n144 256.663
R854 B.n981 B.n143 256.663
R855 B.n981 B.n142 256.663
R856 B.n981 B.n141 256.663
R857 B.n981 B.n140 256.663
R858 B.n981 B.n139 256.663
R859 B.n981 B.n138 256.663
R860 B.n981 B.n137 256.663
R861 B.n981 B.n136 256.663
R862 B.n981 B.n135 256.663
R863 B.n981 B.n134 256.663
R864 B.n981 B.n133 256.663
R865 B.n981 B.n132 256.663
R866 B.n981 B.n131 256.663
R867 B.n981 B.n130 256.663
R868 B.n981 B.n129 256.663
R869 B.n981 B.n128 256.663
R870 B.n981 B.n127 256.663
R871 B.n981 B.n126 256.663
R872 B.n981 B.n125 256.663
R873 B.n981 B.n124 256.663
R874 B.n981 B.n123 256.663
R875 B.n981 B.n122 256.663
R876 B.n981 B.n121 256.663
R877 B.n981 B.n120 256.663
R878 B.n981 B.n119 256.663
R879 B.n981 B.n118 256.663
R880 B.n981 B.n117 256.663
R881 B.n981 B.n116 256.663
R882 B.n981 B.n115 256.663
R883 B.n981 B.n114 256.663
R884 B.n981 B.n113 256.663
R885 B.n981 B.n112 256.663
R886 B.n981 B.n111 256.663
R887 B.n981 B.n110 256.663
R888 B.n981 B.n109 256.663
R889 B.n981 B.n108 256.663
R890 B.n981 B.n107 256.663
R891 B.n981 B.n106 256.663
R892 B.n981 B.n105 256.663
R893 B.n981 B.n104 256.663
R894 B.n981 B.n103 256.663
R895 B.n982 B.n981 256.663
R896 B.n743 B.n742 256.663
R897 B.n742 B.n477 256.663
R898 B.n742 B.n478 256.663
R899 B.n742 B.n479 256.663
R900 B.n742 B.n480 256.663
R901 B.n742 B.n481 256.663
R902 B.n742 B.n482 256.663
R903 B.n742 B.n483 256.663
R904 B.n742 B.n484 256.663
R905 B.n742 B.n485 256.663
R906 B.n742 B.n486 256.663
R907 B.n742 B.n487 256.663
R908 B.n742 B.n488 256.663
R909 B.n742 B.n489 256.663
R910 B.n742 B.n490 256.663
R911 B.n742 B.n491 256.663
R912 B.n742 B.n492 256.663
R913 B.n742 B.n493 256.663
R914 B.n742 B.n494 256.663
R915 B.n742 B.n495 256.663
R916 B.n742 B.n496 256.663
R917 B.n742 B.n497 256.663
R918 B.n742 B.n498 256.663
R919 B.n742 B.n499 256.663
R920 B.n742 B.n500 256.663
R921 B.n742 B.n501 256.663
R922 B.n742 B.n502 256.663
R923 B.n742 B.n503 256.663
R924 B.n742 B.n504 256.663
R925 B.n742 B.n505 256.663
R926 B.n742 B.n506 256.663
R927 B.n742 B.n507 256.663
R928 B.n742 B.n508 256.663
R929 B.n742 B.n509 256.663
R930 B.n742 B.n510 256.663
R931 B.n742 B.n511 256.663
R932 B.n742 B.n512 256.663
R933 B.n742 B.n513 256.663
R934 B.n742 B.n514 256.663
R935 B.n742 B.n515 256.663
R936 B.n742 B.n516 256.663
R937 B.n742 B.n517 256.663
R938 B.n742 B.n518 256.663
R939 B.n742 B.n519 256.663
R940 B.n742 B.n520 256.663
R941 B.n742 B.n521 256.663
R942 B.n742 B.n522 256.663
R943 B.n742 B.n523 256.663
R944 B.n742 B.n524 256.663
R945 B.n742 B.n525 256.663
R946 B.n742 B.n526 256.663
R947 B.n742 B.n527 256.663
R948 B.n748 B.n474 163.367
R949 B.n748 B.n468 163.367
R950 B.n756 B.n468 163.367
R951 B.n756 B.n466 163.367
R952 B.n760 B.n466 163.367
R953 B.n760 B.n460 163.367
R954 B.n767 B.n460 163.367
R955 B.n767 B.n458 163.367
R956 B.n771 B.n458 163.367
R957 B.n771 B.n452 163.367
R958 B.n779 B.n452 163.367
R959 B.n779 B.n450 163.367
R960 B.n783 B.n450 163.367
R961 B.n783 B.n444 163.367
R962 B.n791 B.n444 163.367
R963 B.n791 B.n442 163.367
R964 B.n795 B.n442 163.367
R965 B.n795 B.n436 163.367
R966 B.n803 B.n436 163.367
R967 B.n803 B.n434 163.367
R968 B.n807 B.n434 163.367
R969 B.n807 B.n428 163.367
R970 B.n815 B.n428 163.367
R971 B.n815 B.n426 163.367
R972 B.n819 B.n426 163.367
R973 B.n819 B.n420 163.367
R974 B.n827 B.n420 163.367
R975 B.n827 B.n418 163.367
R976 B.n831 B.n418 163.367
R977 B.n831 B.n412 163.367
R978 B.n839 B.n412 163.367
R979 B.n839 B.n410 163.367
R980 B.n843 B.n410 163.367
R981 B.n843 B.n404 163.367
R982 B.n851 B.n404 163.367
R983 B.n851 B.n402 163.367
R984 B.n855 B.n402 163.367
R985 B.n855 B.n396 163.367
R986 B.n863 B.n396 163.367
R987 B.n863 B.n394 163.367
R988 B.n867 B.n394 163.367
R989 B.n867 B.n388 163.367
R990 B.n875 B.n388 163.367
R991 B.n875 B.n386 163.367
R992 B.n879 B.n386 163.367
R993 B.n879 B.n380 163.367
R994 B.n887 B.n380 163.367
R995 B.n887 B.n378 163.367
R996 B.n891 B.n378 163.367
R997 B.n891 B.n372 163.367
R998 B.n900 B.n372 163.367
R999 B.n900 B.n370 163.367
R1000 B.n904 B.n370 163.367
R1001 B.n904 B.n2 163.367
R1002 B.n1094 B.n2 163.367
R1003 B.n1094 B.n3 163.367
R1004 B.n1090 B.n3 163.367
R1005 B.n1090 B.n9 163.367
R1006 B.n1086 B.n9 163.367
R1007 B.n1086 B.n11 163.367
R1008 B.n1082 B.n11 163.367
R1009 B.n1082 B.n16 163.367
R1010 B.n1078 B.n16 163.367
R1011 B.n1078 B.n18 163.367
R1012 B.n1074 B.n18 163.367
R1013 B.n1074 B.n23 163.367
R1014 B.n1070 B.n23 163.367
R1015 B.n1070 B.n25 163.367
R1016 B.n1066 B.n25 163.367
R1017 B.n1066 B.n30 163.367
R1018 B.n1062 B.n30 163.367
R1019 B.n1062 B.n32 163.367
R1020 B.n1058 B.n32 163.367
R1021 B.n1058 B.n37 163.367
R1022 B.n1054 B.n37 163.367
R1023 B.n1054 B.n39 163.367
R1024 B.n1050 B.n39 163.367
R1025 B.n1050 B.n44 163.367
R1026 B.n1046 B.n44 163.367
R1027 B.n1046 B.n46 163.367
R1028 B.n1042 B.n46 163.367
R1029 B.n1042 B.n51 163.367
R1030 B.n1038 B.n51 163.367
R1031 B.n1038 B.n53 163.367
R1032 B.n1034 B.n53 163.367
R1033 B.n1034 B.n58 163.367
R1034 B.n1030 B.n58 163.367
R1035 B.n1030 B.n60 163.367
R1036 B.n1026 B.n60 163.367
R1037 B.n1026 B.n65 163.367
R1038 B.n1022 B.n65 163.367
R1039 B.n1022 B.n67 163.367
R1040 B.n1018 B.n67 163.367
R1041 B.n1018 B.n72 163.367
R1042 B.n1014 B.n72 163.367
R1043 B.n1014 B.n74 163.367
R1044 B.n1010 B.n74 163.367
R1045 B.n1010 B.n79 163.367
R1046 B.n1006 B.n79 163.367
R1047 B.n1006 B.n81 163.367
R1048 B.n1002 B.n81 163.367
R1049 B.n1002 B.n86 163.367
R1050 B.n998 B.n86 163.367
R1051 B.n998 B.n88 163.367
R1052 B.n995 B.n88 163.367
R1053 B.n995 B.n93 163.367
R1054 B.n991 B.n93 163.367
R1055 B.n991 B.n95 163.367
R1056 B.n987 B.n95 163.367
R1057 B.n987 B.n100 163.367
R1058 B.n741 B.n476 163.367
R1059 B.n741 B.n529 163.367
R1060 B.n737 B.n736 163.367
R1061 B.n733 B.n732 163.367
R1062 B.n729 B.n728 163.367
R1063 B.n725 B.n724 163.367
R1064 B.n721 B.n720 163.367
R1065 B.n717 B.n716 163.367
R1066 B.n713 B.n712 163.367
R1067 B.n709 B.n708 163.367
R1068 B.n705 B.n704 163.367
R1069 B.n701 B.n700 163.367
R1070 B.n697 B.n696 163.367
R1071 B.n693 B.n692 163.367
R1072 B.n689 B.n688 163.367
R1073 B.n685 B.n684 163.367
R1074 B.n681 B.n680 163.367
R1075 B.n677 B.n676 163.367
R1076 B.n673 B.n672 163.367
R1077 B.n669 B.n668 163.367
R1078 B.n665 B.n664 163.367
R1079 B.n661 B.n660 163.367
R1080 B.n657 B.n656 163.367
R1081 B.n653 B.n652 163.367
R1082 B.n648 B.n647 163.367
R1083 B.n644 B.n643 163.367
R1084 B.n640 B.n639 163.367
R1085 B.n636 B.n635 163.367
R1086 B.n632 B.n631 163.367
R1087 B.n627 B.n626 163.367
R1088 B.n623 B.n622 163.367
R1089 B.n619 B.n618 163.367
R1090 B.n615 B.n614 163.367
R1091 B.n611 B.n610 163.367
R1092 B.n607 B.n606 163.367
R1093 B.n603 B.n602 163.367
R1094 B.n599 B.n598 163.367
R1095 B.n595 B.n594 163.367
R1096 B.n591 B.n590 163.367
R1097 B.n587 B.n586 163.367
R1098 B.n583 B.n582 163.367
R1099 B.n579 B.n578 163.367
R1100 B.n575 B.n574 163.367
R1101 B.n571 B.n570 163.367
R1102 B.n567 B.n566 163.367
R1103 B.n563 B.n562 163.367
R1104 B.n559 B.n558 163.367
R1105 B.n555 B.n554 163.367
R1106 B.n551 B.n550 163.367
R1107 B.n547 B.n546 163.367
R1108 B.n543 B.n542 163.367
R1109 B.n539 B.n538 163.367
R1110 B.n535 B.n528 163.367
R1111 B.n750 B.n472 163.367
R1112 B.n750 B.n470 163.367
R1113 B.n754 B.n470 163.367
R1114 B.n754 B.n464 163.367
R1115 B.n762 B.n464 163.367
R1116 B.n762 B.n462 163.367
R1117 B.n766 B.n462 163.367
R1118 B.n766 B.n456 163.367
R1119 B.n773 B.n456 163.367
R1120 B.n773 B.n454 163.367
R1121 B.n777 B.n454 163.367
R1122 B.n777 B.n448 163.367
R1123 B.n785 B.n448 163.367
R1124 B.n785 B.n446 163.367
R1125 B.n789 B.n446 163.367
R1126 B.n789 B.n439 163.367
R1127 B.n797 B.n439 163.367
R1128 B.n797 B.n437 163.367
R1129 B.n801 B.n437 163.367
R1130 B.n801 B.n432 163.367
R1131 B.n809 B.n432 163.367
R1132 B.n809 B.n430 163.367
R1133 B.n813 B.n430 163.367
R1134 B.n813 B.n424 163.367
R1135 B.n821 B.n424 163.367
R1136 B.n821 B.n422 163.367
R1137 B.n825 B.n422 163.367
R1138 B.n825 B.n416 163.367
R1139 B.n833 B.n416 163.367
R1140 B.n833 B.n414 163.367
R1141 B.n837 B.n414 163.367
R1142 B.n837 B.n408 163.367
R1143 B.n845 B.n408 163.367
R1144 B.n845 B.n406 163.367
R1145 B.n849 B.n406 163.367
R1146 B.n849 B.n400 163.367
R1147 B.n857 B.n400 163.367
R1148 B.n857 B.n398 163.367
R1149 B.n861 B.n398 163.367
R1150 B.n861 B.n392 163.367
R1151 B.n869 B.n392 163.367
R1152 B.n869 B.n390 163.367
R1153 B.n873 B.n390 163.367
R1154 B.n873 B.n384 163.367
R1155 B.n881 B.n384 163.367
R1156 B.n881 B.n382 163.367
R1157 B.n885 B.n382 163.367
R1158 B.n885 B.n376 163.367
R1159 B.n893 B.n376 163.367
R1160 B.n893 B.n374 163.367
R1161 B.n898 B.n374 163.367
R1162 B.n898 B.n368 163.367
R1163 B.n906 B.n368 163.367
R1164 B.n907 B.n906 163.367
R1165 B.n907 B.n5 163.367
R1166 B.n6 B.n5 163.367
R1167 B.n7 B.n6 163.367
R1168 B.n912 B.n7 163.367
R1169 B.n912 B.n12 163.367
R1170 B.n13 B.n12 163.367
R1171 B.n14 B.n13 163.367
R1172 B.n917 B.n14 163.367
R1173 B.n917 B.n19 163.367
R1174 B.n20 B.n19 163.367
R1175 B.n21 B.n20 163.367
R1176 B.n922 B.n21 163.367
R1177 B.n922 B.n26 163.367
R1178 B.n27 B.n26 163.367
R1179 B.n28 B.n27 163.367
R1180 B.n927 B.n28 163.367
R1181 B.n927 B.n33 163.367
R1182 B.n34 B.n33 163.367
R1183 B.n35 B.n34 163.367
R1184 B.n932 B.n35 163.367
R1185 B.n932 B.n40 163.367
R1186 B.n41 B.n40 163.367
R1187 B.n42 B.n41 163.367
R1188 B.n937 B.n42 163.367
R1189 B.n937 B.n47 163.367
R1190 B.n48 B.n47 163.367
R1191 B.n49 B.n48 163.367
R1192 B.n942 B.n49 163.367
R1193 B.n942 B.n54 163.367
R1194 B.n55 B.n54 163.367
R1195 B.n56 B.n55 163.367
R1196 B.n947 B.n56 163.367
R1197 B.n947 B.n61 163.367
R1198 B.n62 B.n61 163.367
R1199 B.n63 B.n62 163.367
R1200 B.n952 B.n63 163.367
R1201 B.n952 B.n68 163.367
R1202 B.n69 B.n68 163.367
R1203 B.n70 B.n69 163.367
R1204 B.n957 B.n70 163.367
R1205 B.n957 B.n75 163.367
R1206 B.n76 B.n75 163.367
R1207 B.n77 B.n76 163.367
R1208 B.n962 B.n77 163.367
R1209 B.n962 B.n82 163.367
R1210 B.n83 B.n82 163.367
R1211 B.n84 B.n83 163.367
R1212 B.n967 B.n84 163.367
R1213 B.n967 B.n89 163.367
R1214 B.n90 B.n89 163.367
R1215 B.n91 B.n90 163.367
R1216 B.n972 B.n91 163.367
R1217 B.n972 B.n96 163.367
R1218 B.n97 B.n96 163.367
R1219 B.n98 B.n97 163.367
R1220 B.n155 B.n98 163.367
R1221 B.n162 B.n102 163.367
R1222 B.n166 B.n165 163.367
R1223 B.n170 B.n169 163.367
R1224 B.n174 B.n173 163.367
R1225 B.n178 B.n177 163.367
R1226 B.n182 B.n181 163.367
R1227 B.n186 B.n185 163.367
R1228 B.n190 B.n189 163.367
R1229 B.n194 B.n193 163.367
R1230 B.n198 B.n197 163.367
R1231 B.n202 B.n201 163.367
R1232 B.n206 B.n205 163.367
R1233 B.n210 B.n209 163.367
R1234 B.n214 B.n213 163.367
R1235 B.n218 B.n217 163.367
R1236 B.n222 B.n221 163.367
R1237 B.n226 B.n225 163.367
R1238 B.n230 B.n229 163.367
R1239 B.n234 B.n233 163.367
R1240 B.n238 B.n237 163.367
R1241 B.n242 B.n241 163.367
R1242 B.n246 B.n245 163.367
R1243 B.n250 B.n249 163.367
R1244 B.n254 B.n253 163.367
R1245 B.n258 B.n257 163.367
R1246 B.n262 B.n261 163.367
R1247 B.n266 B.n265 163.367
R1248 B.n270 B.n269 163.367
R1249 B.n274 B.n273 163.367
R1250 B.n278 B.n277 163.367
R1251 B.n282 B.n281 163.367
R1252 B.n286 B.n285 163.367
R1253 B.n290 B.n289 163.367
R1254 B.n294 B.n293 163.367
R1255 B.n298 B.n297 163.367
R1256 B.n302 B.n301 163.367
R1257 B.n306 B.n305 163.367
R1258 B.n310 B.n309 163.367
R1259 B.n314 B.n313 163.367
R1260 B.n318 B.n317 163.367
R1261 B.n322 B.n321 163.367
R1262 B.n326 B.n325 163.367
R1263 B.n330 B.n329 163.367
R1264 B.n334 B.n333 163.367
R1265 B.n338 B.n337 163.367
R1266 B.n342 B.n341 163.367
R1267 B.n346 B.n345 163.367
R1268 B.n350 B.n349 163.367
R1269 B.n354 B.n353 163.367
R1270 B.n358 B.n357 163.367
R1271 B.n362 B.n361 163.367
R1272 B.n364 B.n154 163.367
R1273 B.n532 B.t18 119.891
R1274 B.n156 B.t14 119.891
R1275 B.n530 B.t12 119.871
R1276 B.n159 B.t7 119.871
R1277 B.n742 B.n473 78.0705
R1278 B.n981 B.n99 78.0705
R1279 B.n744 B.n743 71.676
R1280 B.n529 B.n477 71.676
R1281 B.n736 B.n478 71.676
R1282 B.n732 B.n479 71.676
R1283 B.n728 B.n480 71.676
R1284 B.n724 B.n481 71.676
R1285 B.n720 B.n482 71.676
R1286 B.n716 B.n483 71.676
R1287 B.n712 B.n484 71.676
R1288 B.n708 B.n485 71.676
R1289 B.n704 B.n486 71.676
R1290 B.n700 B.n487 71.676
R1291 B.n696 B.n488 71.676
R1292 B.n692 B.n489 71.676
R1293 B.n688 B.n490 71.676
R1294 B.n684 B.n491 71.676
R1295 B.n680 B.n492 71.676
R1296 B.n676 B.n493 71.676
R1297 B.n672 B.n494 71.676
R1298 B.n668 B.n495 71.676
R1299 B.n664 B.n496 71.676
R1300 B.n660 B.n497 71.676
R1301 B.n656 B.n498 71.676
R1302 B.n652 B.n499 71.676
R1303 B.n647 B.n500 71.676
R1304 B.n643 B.n501 71.676
R1305 B.n639 B.n502 71.676
R1306 B.n635 B.n503 71.676
R1307 B.n631 B.n504 71.676
R1308 B.n626 B.n505 71.676
R1309 B.n622 B.n506 71.676
R1310 B.n618 B.n507 71.676
R1311 B.n614 B.n508 71.676
R1312 B.n610 B.n509 71.676
R1313 B.n606 B.n510 71.676
R1314 B.n602 B.n511 71.676
R1315 B.n598 B.n512 71.676
R1316 B.n594 B.n513 71.676
R1317 B.n590 B.n514 71.676
R1318 B.n586 B.n515 71.676
R1319 B.n582 B.n516 71.676
R1320 B.n578 B.n517 71.676
R1321 B.n574 B.n518 71.676
R1322 B.n570 B.n519 71.676
R1323 B.n566 B.n520 71.676
R1324 B.n562 B.n521 71.676
R1325 B.n558 B.n522 71.676
R1326 B.n554 B.n523 71.676
R1327 B.n550 B.n524 71.676
R1328 B.n546 B.n525 71.676
R1329 B.n542 B.n526 71.676
R1330 B.n538 B.n527 71.676
R1331 B.n983 B.n982 71.676
R1332 B.n162 B.n103 71.676
R1333 B.n166 B.n104 71.676
R1334 B.n170 B.n105 71.676
R1335 B.n174 B.n106 71.676
R1336 B.n178 B.n107 71.676
R1337 B.n182 B.n108 71.676
R1338 B.n186 B.n109 71.676
R1339 B.n190 B.n110 71.676
R1340 B.n194 B.n111 71.676
R1341 B.n198 B.n112 71.676
R1342 B.n202 B.n113 71.676
R1343 B.n206 B.n114 71.676
R1344 B.n210 B.n115 71.676
R1345 B.n214 B.n116 71.676
R1346 B.n218 B.n117 71.676
R1347 B.n222 B.n118 71.676
R1348 B.n226 B.n119 71.676
R1349 B.n230 B.n120 71.676
R1350 B.n234 B.n121 71.676
R1351 B.n238 B.n122 71.676
R1352 B.n242 B.n123 71.676
R1353 B.n246 B.n124 71.676
R1354 B.n250 B.n125 71.676
R1355 B.n254 B.n126 71.676
R1356 B.n258 B.n127 71.676
R1357 B.n262 B.n128 71.676
R1358 B.n266 B.n129 71.676
R1359 B.n270 B.n130 71.676
R1360 B.n274 B.n131 71.676
R1361 B.n278 B.n132 71.676
R1362 B.n282 B.n133 71.676
R1363 B.n286 B.n134 71.676
R1364 B.n290 B.n135 71.676
R1365 B.n294 B.n136 71.676
R1366 B.n298 B.n137 71.676
R1367 B.n302 B.n138 71.676
R1368 B.n306 B.n139 71.676
R1369 B.n310 B.n140 71.676
R1370 B.n314 B.n141 71.676
R1371 B.n318 B.n142 71.676
R1372 B.n322 B.n143 71.676
R1373 B.n326 B.n144 71.676
R1374 B.n330 B.n145 71.676
R1375 B.n334 B.n146 71.676
R1376 B.n338 B.n147 71.676
R1377 B.n342 B.n148 71.676
R1378 B.n346 B.n149 71.676
R1379 B.n350 B.n150 71.676
R1380 B.n354 B.n151 71.676
R1381 B.n358 B.n152 71.676
R1382 B.n362 B.n153 71.676
R1383 B.n980 B.n154 71.676
R1384 B.n980 B.n979 71.676
R1385 B.n364 B.n153 71.676
R1386 B.n361 B.n152 71.676
R1387 B.n357 B.n151 71.676
R1388 B.n353 B.n150 71.676
R1389 B.n349 B.n149 71.676
R1390 B.n345 B.n148 71.676
R1391 B.n341 B.n147 71.676
R1392 B.n337 B.n146 71.676
R1393 B.n333 B.n145 71.676
R1394 B.n329 B.n144 71.676
R1395 B.n325 B.n143 71.676
R1396 B.n321 B.n142 71.676
R1397 B.n317 B.n141 71.676
R1398 B.n313 B.n140 71.676
R1399 B.n309 B.n139 71.676
R1400 B.n305 B.n138 71.676
R1401 B.n301 B.n137 71.676
R1402 B.n297 B.n136 71.676
R1403 B.n293 B.n135 71.676
R1404 B.n289 B.n134 71.676
R1405 B.n285 B.n133 71.676
R1406 B.n281 B.n132 71.676
R1407 B.n277 B.n131 71.676
R1408 B.n273 B.n130 71.676
R1409 B.n269 B.n129 71.676
R1410 B.n265 B.n128 71.676
R1411 B.n261 B.n127 71.676
R1412 B.n257 B.n126 71.676
R1413 B.n253 B.n125 71.676
R1414 B.n249 B.n124 71.676
R1415 B.n245 B.n123 71.676
R1416 B.n241 B.n122 71.676
R1417 B.n237 B.n121 71.676
R1418 B.n233 B.n120 71.676
R1419 B.n229 B.n119 71.676
R1420 B.n225 B.n118 71.676
R1421 B.n221 B.n117 71.676
R1422 B.n217 B.n116 71.676
R1423 B.n213 B.n115 71.676
R1424 B.n209 B.n114 71.676
R1425 B.n205 B.n113 71.676
R1426 B.n201 B.n112 71.676
R1427 B.n197 B.n111 71.676
R1428 B.n193 B.n110 71.676
R1429 B.n189 B.n109 71.676
R1430 B.n185 B.n108 71.676
R1431 B.n181 B.n107 71.676
R1432 B.n177 B.n106 71.676
R1433 B.n173 B.n105 71.676
R1434 B.n169 B.n104 71.676
R1435 B.n165 B.n103 71.676
R1436 B.n982 B.n102 71.676
R1437 B.n743 B.n476 71.676
R1438 B.n737 B.n477 71.676
R1439 B.n733 B.n478 71.676
R1440 B.n729 B.n479 71.676
R1441 B.n725 B.n480 71.676
R1442 B.n721 B.n481 71.676
R1443 B.n717 B.n482 71.676
R1444 B.n713 B.n483 71.676
R1445 B.n709 B.n484 71.676
R1446 B.n705 B.n485 71.676
R1447 B.n701 B.n486 71.676
R1448 B.n697 B.n487 71.676
R1449 B.n693 B.n488 71.676
R1450 B.n689 B.n489 71.676
R1451 B.n685 B.n490 71.676
R1452 B.n681 B.n491 71.676
R1453 B.n677 B.n492 71.676
R1454 B.n673 B.n493 71.676
R1455 B.n669 B.n494 71.676
R1456 B.n665 B.n495 71.676
R1457 B.n661 B.n496 71.676
R1458 B.n657 B.n497 71.676
R1459 B.n653 B.n498 71.676
R1460 B.n648 B.n499 71.676
R1461 B.n644 B.n500 71.676
R1462 B.n640 B.n501 71.676
R1463 B.n636 B.n502 71.676
R1464 B.n632 B.n503 71.676
R1465 B.n627 B.n504 71.676
R1466 B.n623 B.n505 71.676
R1467 B.n619 B.n506 71.676
R1468 B.n615 B.n507 71.676
R1469 B.n611 B.n508 71.676
R1470 B.n607 B.n509 71.676
R1471 B.n603 B.n510 71.676
R1472 B.n599 B.n511 71.676
R1473 B.n595 B.n512 71.676
R1474 B.n591 B.n513 71.676
R1475 B.n587 B.n514 71.676
R1476 B.n583 B.n515 71.676
R1477 B.n579 B.n516 71.676
R1478 B.n575 B.n517 71.676
R1479 B.n571 B.n518 71.676
R1480 B.n567 B.n519 71.676
R1481 B.n563 B.n520 71.676
R1482 B.n559 B.n521 71.676
R1483 B.n555 B.n522 71.676
R1484 B.n551 B.n523 71.676
R1485 B.n547 B.n524 71.676
R1486 B.n543 B.n525 71.676
R1487 B.n539 B.n526 71.676
R1488 B.n535 B.n527 71.676
R1489 B.n533 B.t17 68.1089
R1490 B.n157 B.t15 68.1089
R1491 B.n531 B.t11 68.0901
R1492 B.n160 B.t8 68.0901
R1493 B.n629 B.n533 59.5399
R1494 B.n650 B.n531 59.5399
R1495 B.n161 B.n160 59.5399
R1496 B.n158 B.n157 59.5399
R1497 B.n533 B.n532 51.7823
R1498 B.n531 B.n530 51.7823
R1499 B.n160 B.n159 51.7823
R1500 B.n157 B.n156 51.7823
R1501 B.n749 B.n473 38.193
R1502 B.n749 B.n469 38.193
R1503 B.n755 B.n469 38.193
R1504 B.n755 B.n465 38.193
R1505 B.n761 B.n465 38.193
R1506 B.n761 B.n461 38.193
R1507 B.t10 B.n461 38.193
R1508 B.t10 B.n457 38.193
R1509 B.n772 B.n457 38.193
R1510 B.n772 B.n453 38.193
R1511 B.n778 B.n453 38.193
R1512 B.n778 B.n449 38.193
R1513 B.n784 B.n449 38.193
R1514 B.n784 B.n445 38.193
R1515 B.n790 B.n445 38.193
R1516 B.n790 B.n440 38.193
R1517 B.n796 B.n440 38.193
R1518 B.n796 B.n441 38.193
R1519 B.n802 B.n433 38.193
R1520 B.n808 B.n433 38.193
R1521 B.n808 B.n429 38.193
R1522 B.n814 B.n429 38.193
R1523 B.n814 B.n425 38.193
R1524 B.n820 B.n425 38.193
R1525 B.n826 B.n421 38.193
R1526 B.n826 B.n417 38.193
R1527 B.n832 B.n417 38.193
R1528 B.n832 B.n413 38.193
R1529 B.n838 B.n413 38.193
R1530 B.n838 B.n409 38.193
R1531 B.n844 B.n409 38.193
R1532 B.n850 B.n405 38.193
R1533 B.n850 B.n401 38.193
R1534 B.n856 B.n401 38.193
R1535 B.n856 B.n397 38.193
R1536 B.n862 B.n397 38.193
R1537 B.n862 B.n393 38.193
R1538 B.n868 B.n393 38.193
R1539 B.n874 B.n389 38.193
R1540 B.n874 B.n385 38.193
R1541 B.n880 B.n385 38.193
R1542 B.n880 B.n381 38.193
R1543 B.n886 B.n381 38.193
R1544 B.n886 B.n377 38.193
R1545 B.n892 B.n377 38.193
R1546 B.n899 B.n373 38.193
R1547 B.n899 B.n369 38.193
R1548 B.n905 B.n369 38.193
R1549 B.n905 B.n4 38.193
R1550 B.n1093 B.n4 38.193
R1551 B.n1093 B.n1092 38.193
R1552 B.n1092 B.n1091 38.193
R1553 B.n1091 B.n8 38.193
R1554 B.n1085 B.n8 38.193
R1555 B.n1085 B.n1084 38.193
R1556 B.n1083 B.n15 38.193
R1557 B.n1077 B.n15 38.193
R1558 B.n1077 B.n1076 38.193
R1559 B.n1076 B.n1075 38.193
R1560 B.n1075 B.n22 38.193
R1561 B.n1069 B.n22 38.193
R1562 B.n1069 B.n1068 38.193
R1563 B.n1067 B.n29 38.193
R1564 B.n1061 B.n29 38.193
R1565 B.n1061 B.n1060 38.193
R1566 B.n1060 B.n1059 38.193
R1567 B.n1059 B.n36 38.193
R1568 B.n1053 B.n36 38.193
R1569 B.n1053 B.n1052 38.193
R1570 B.n1051 B.n43 38.193
R1571 B.n1045 B.n43 38.193
R1572 B.n1045 B.n1044 38.193
R1573 B.n1044 B.n1043 38.193
R1574 B.n1043 B.n50 38.193
R1575 B.n1037 B.n50 38.193
R1576 B.n1037 B.n1036 38.193
R1577 B.n1035 B.n57 38.193
R1578 B.n1029 B.n57 38.193
R1579 B.n1029 B.n1028 38.193
R1580 B.n1028 B.n1027 38.193
R1581 B.n1027 B.n64 38.193
R1582 B.n1021 B.n64 38.193
R1583 B.n1020 B.n1019 38.193
R1584 B.n1019 B.n71 38.193
R1585 B.n1013 B.n71 38.193
R1586 B.n1013 B.n1012 38.193
R1587 B.n1012 B.n1011 38.193
R1588 B.n1011 B.n78 38.193
R1589 B.n1005 B.n78 38.193
R1590 B.n1005 B.n1004 38.193
R1591 B.n1004 B.n1003 38.193
R1592 B.n1003 B.n85 38.193
R1593 B.t6 B.n85 38.193
R1594 B.t6 B.n997 38.193
R1595 B.n997 B.n996 38.193
R1596 B.n996 B.n92 38.193
R1597 B.n990 B.n92 38.193
R1598 B.n990 B.n989 38.193
R1599 B.n989 B.n988 38.193
R1600 B.n988 B.n99 38.193
R1601 B.n985 B.n984 36.9956
R1602 B.n978 B.n977 36.9956
R1603 B.n534 B.n471 36.9956
R1604 B.n746 B.n745 36.9956
R1605 B.n802 B.t22 35.9464
R1606 B.n1021 B.t0 35.9464
R1607 B.n820 B.t20 34.8231
R1608 B.t3 B.n1035 34.8231
R1609 B.n844 B.t4 29.2065
R1610 B.t19 B.n1051 29.2065
R1611 B.n868 B.t21 23.59
R1612 B.t2 B.n1067 23.59
R1613 B.t1 B.n373 20.2201
R1614 B.n1084 B.t23 20.2201
R1615 B B.n1095 18.0485
R1616 B.n892 B.t1 17.9734
R1617 B.t23 B.n1083 17.9734
R1618 B.t21 B.n389 14.6035
R1619 B.n1068 B.t2 14.6035
R1620 B.n984 B.n101 10.6151
R1621 B.n163 B.n101 10.6151
R1622 B.n164 B.n163 10.6151
R1623 B.n167 B.n164 10.6151
R1624 B.n168 B.n167 10.6151
R1625 B.n171 B.n168 10.6151
R1626 B.n172 B.n171 10.6151
R1627 B.n175 B.n172 10.6151
R1628 B.n176 B.n175 10.6151
R1629 B.n179 B.n176 10.6151
R1630 B.n180 B.n179 10.6151
R1631 B.n183 B.n180 10.6151
R1632 B.n184 B.n183 10.6151
R1633 B.n187 B.n184 10.6151
R1634 B.n188 B.n187 10.6151
R1635 B.n191 B.n188 10.6151
R1636 B.n192 B.n191 10.6151
R1637 B.n195 B.n192 10.6151
R1638 B.n196 B.n195 10.6151
R1639 B.n199 B.n196 10.6151
R1640 B.n200 B.n199 10.6151
R1641 B.n203 B.n200 10.6151
R1642 B.n204 B.n203 10.6151
R1643 B.n207 B.n204 10.6151
R1644 B.n208 B.n207 10.6151
R1645 B.n211 B.n208 10.6151
R1646 B.n212 B.n211 10.6151
R1647 B.n215 B.n212 10.6151
R1648 B.n216 B.n215 10.6151
R1649 B.n219 B.n216 10.6151
R1650 B.n220 B.n219 10.6151
R1651 B.n223 B.n220 10.6151
R1652 B.n224 B.n223 10.6151
R1653 B.n227 B.n224 10.6151
R1654 B.n228 B.n227 10.6151
R1655 B.n231 B.n228 10.6151
R1656 B.n232 B.n231 10.6151
R1657 B.n235 B.n232 10.6151
R1658 B.n236 B.n235 10.6151
R1659 B.n239 B.n236 10.6151
R1660 B.n240 B.n239 10.6151
R1661 B.n243 B.n240 10.6151
R1662 B.n244 B.n243 10.6151
R1663 B.n247 B.n244 10.6151
R1664 B.n248 B.n247 10.6151
R1665 B.n251 B.n248 10.6151
R1666 B.n252 B.n251 10.6151
R1667 B.n256 B.n255 10.6151
R1668 B.n259 B.n256 10.6151
R1669 B.n260 B.n259 10.6151
R1670 B.n263 B.n260 10.6151
R1671 B.n264 B.n263 10.6151
R1672 B.n267 B.n264 10.6151
R1673 B.n268 B.n267 10.6151
R1674 B.n271 B.n268 10.6151
R1675 B.n272 B.n271 10.6151
R1676 B.n276 B.n275 10.6151
R1677 B.n279 B.n276 10.6151
R1678 B.n280 B.n279 10.6151
R1679 B.n283 B.n280 10.6151
R1680 B.n284 B.n283 10.6151
R1681 B.n287 B.n284 10.6151
R1682 B.n288 B.n287 10.6151
R1683 B.n291 B.n288 10.6151
R1684 B.n292 B.n291 10.6151
R1685 B.n295 B.n292 10.6151
R1686 B.n296 B.n295 10.6151
R1687 B.n299 B.n296 10.6151
R1688 B.n300 B.n299 10.6151
R1689 B.n303 B.n300 10.6151
R1690 B.n304 B.n303 10.6151
R1691 B.n307 B.n304 10.6151
R1692 B.n308 B.n307 10.6151
R1693 B.n311 B.n308 10.6151
R1694 B.n312 B.n311 10.6151
R1695 B.n315 B.n312 10.6151
R1696 B.n316 B.n315 10.6151
R1697 B.n319 B.n316 10.6151
R1698 B.n320 B.n319 10.6151
R1699 B.n323 B.n320 10.6151
R1700 B.n324 B.n323 10.6151
R1701 B.n327 B.n324 10.6151
R1702 B.n328 B.n327 10.6151
R1703 B.n331 B.n328 10.6151
R1704 B.n332 B.n331 10.6151
R1705 B.n335 B.n332 10.6151
R1706 B.n336 B.n335 10.6151
R1707 B.n339 B.n336 10.6151
R1708 B.n340 B.n339 10.6151
R1709 B.n343 B.n340 10.6151
R1710 B.n344 B.n343 10.6151
R1711 B.n347 B.n344 10.6151
R1712 B.n348 B.n347 10.6151
R1713 B.n351 B.n348 10.6151
R1714 B.n352 B.n351 10.6151
R1715 B.n355 B.n352 10.6151
R1716 B.n356 B.n355 10.6151
R1717 B.n359 B.n356 10.6151
R1718 B.n360 B.n359 10.6151
R1719 B.n363 B.n360 10.6151
R1720 B.n365 B.n363 10.6151
R1721 B.n366 B.n365 10.6151
R1722 B.n978 B.n366 10.6151
R1723 B.n751 B.n471 10.6151
R1724 B.n752 B.n751 10.6151
R1725 B.n753 B.n752 10.6151
R1726 B.n753 B.n463 10.6151
R1727 B.n763 B.n463 10.6151
R1728 B.n764 B.n763 10.6151
R1729 B.n765 B.n764 10.6151
R1730 B.n765 B.n455 10.6151
R1731 B.n774 B.n455 10.6151
R1732 B.n775 B.n774 10.6151
R1733 B.n776 B.n775 10.6151
R1734 B.n776 B.n447 10.6151
R1735 B.n786 B.n447 10.6151
R1736 B.n787 B.n786 10.6151
R1737 B.n788 B.n787 10.6151
R1738 B.n788 B.n438 10.6151
R1739 B.n798 B.n438 10.6151
R1740 B.n799 B.n798 10.6151
R1741 B.n800 B.n799 10.6151
R1742 B.n800 B.n431 10.6151
R1743 B.n810 B.n431 10.6151
R1744 B.n811 B.n810 10.6151
R1745 B.n812 B.n811 10.6151
R1746 B.n812 B.n423 10.6151
R1747 B.n822 B.n423 10.6151
R1748 B.n823 B.n822 10.6151
R1749 B.n824 B.n823 10.6151
R1750 B.n824 B.n415 10.6151
R1751 B.n834 B.n415 10.6151
R1752 B.n835 B.n834 10.6151
R1753 B.n836 B.n835 10.6151
R1754 B.n836 B.n407 10.6151
R1755 B.n846 B.n407 10.6151
R1756 B.n847 B.n846 10.6151
R1757 B.n848 B.n847 10.6151
R1758 B.n848 B.n399 10.6151
R1759 B.n858 B.n399 10.6151
R1760 B.n859 B.n858 10.6151
R1761 B.n860 B.n859 10.6151
R1762 B.n860 B.n391 10.6151
R1763 B.n870 B.n391 10.6151
R1764 B.n871 B.n870 10.6151
R1765 B.n872 B.n871 10.6151
R1766 B.n872 B.n383 10.6151
R1767 B.n882 B.n383 10.6151
R1768 B.n883 B.n882 10.6151
R1769 B.n884 B.n883 10.6151
R1770 B.n884 B.n375 10.6151
R1771 B.n894 B.n375 10.6151
R1772 B.n895 B.n894 10.6151
R1773 B.n897 B.n895 10.6151
R1774 B.n897 B.n896 10.6151
R1775 B.n896 B.n367 10.6151
R1776 B.n908 B.n367 10.6151
R1777 B.n909 B.n908 10.6151
R1778 B.n910 B.n909 10.6151
R1779 B.n911 B.n910 10.6151
R1780 B.n913 B.n911 10.6151
R1781 B.n914 B.n913 10.6151
R1782 B.n915 B.n914 10.6151
R1783 B.n916 B.n915 10.6151
R1784 B.n918 B.n916 10.6151
R1785 B.n919 B.n918 10.6151
R1786 B.n920 B.n919 10.6151
R1787 B.n921 B.n920 10.6151
R1788 B.n923 B.n921 10.6151
R1789 B.n924 B.n923 10.6151
R1790 B.n925 B.n924 10.6151
R1791 B.n926 B.n925 10.6151
R1792 B.n928 B.n926 10.6151
R1793 B.n929 B.n928 10.6151
R1794 B.n930 B.n929 10.6151
R1795 B.n931 B.n930 10.6151
R1796 B.n933 B.n931 10.6151
R1797 B.n934 B.n933 10.6151
R1798 B.n935 B.n934 10.6151
R1799 B.n936 B.n935 10.6151
R1800 B.n938 B.n936 10.6151
R1801 B.n939 B.n938 10.6151
R1802 B.n940 B.n939 10.6151
R1803 B.n941 B.n940 10.6151
R1804 B.n943 B.n941 10.6151
R1805 B.n944 B.n943 10.6151
R1806 B.n945 B.n944 10.6151
R1807 B.n946 B.n945 10.6151
R1808 B.n948 B.n946 10.6151
R1809 B.n949 B.n948 10.6151
R1810 B.n950 B.n949 10.6151
R1811 B.n951 B.n950 10.6151
R1812 B.n953 B.n951 10.6151
R1813 B.n954 B.n953 10.6151
R1814 B.n955 B.n954 10.6151
R1815 B.n956 B.n955 10.6151
R1816 B.n958 B.n956 10.6151
R1817 B.n959 B.n958 10.6151
R1818 B.n960 B.n959 10.6151
R1819 B.n961 B.n960 10.6151
R1820 B.n963 B.n961 10.6151
R1821 B.n964 B.n963 10.6151
R1822 B.n965 B.n964 10.6151
R1823 B.n966 B.n965 10.6151
R1824 B.n968 B.n966 10.6151
R1825 B.n969 B.n968 10.6151
R1826 B.n970 B.n969 10.6151
R1827 B.n971 B.n970 10.6151
R1828 B.n973 B.n971 10.6151
R1829 B.n974 B.n973 10.6151
R1830 B.n975 B.n974 10.6151
R1831 B.n976 B.n975 10.6151
R1832 B.n977 B.n976 10.6151
R1833 B.n745 B.n475 10.6151
R1834 B.n740 B.n475 10.6151
R1835 B.n740 B.n739 10.6151
R1836 B.n739 B.n738 10.6151
R1837 B.n738 B.n735 10.6151
R1838 B.n735 B.n734 10.6151
R1839 B.n734 B.n731 10.6151
R1840 B.n731 B.n730 10.6151
R1841 B.n730 B.n727 10.6151
R1842 B.n727 B.n726 10.6151
R1843 B.n726 B.n723 10.6151
R1844 B.n723 B.n722 10.6151
R1845 B.n722 B.n719 10.6151
R1846 B.n719 B.n718 10.6151
R1847 B.n718 B.n715 10.6151
R1848 B.n715 B.n714 10.6151
R1849 B.n714 B.n711 10.6151
R1850 B.n711 B.n710 10.6151
R1851 B.n710 B.n707 10.6151
R1852 B.n707 B.n706 10.6151
R1853 B.n706 B.n703 10.6151
R1854 B.n703 B.n702 10.6151
R1855 B.n702 B.n699 10.6151
R1856 B.n699 B.n698 10.6151
R1857 B.n698 B.n695 10.6151
R1858 B.n695 B.n694 10.6151
R1859 B.n694 B.n691 10.6151
R1860 B.n691 B.n690 10.6151
R1861 B.n690 B.n687 10.6151
R1862 B.n687 B.n686 10.6151
R1863 B.n686 B.n683 10.6151
R1864 B.n683 B.n682 10.6151
R1865 B.n682 B.n679 10.6151
R1866 B.n679 B.n678 10.6151
R1867 B.n678 B.n675 10.6151
R1868 B.n675 B.n674 10.6151
R1869 B.n674 B.n671 10.6151
R1870 B.n671 B.n670 10.6151
R1871 B.n670 B.n667 10.6151
R1872 B.n667 B.n666 10.6151
R1873 B.n666 B.n663 10.6151
R1874 B.n663 B.n662 10.6151
R1875 B.n662 B.n659 10.6151
R1876 B.n659 B.n658 10.6151
R1877 B.n658 B.n655 10.6151
R1878 B.n655 B.n654 10.6151
R1879 B.n654 B.n651 10.6151
R1880 B.n649 B.n646 10.6151
R1881 B.n646 B.n645 10.6151
R1882 B.n645 B.n642 10.6151
R1883 B.n642 B.n641 10.6151
R1884 B.n641 B.n638 10.6151
R1885 B.n638 B.n637 10.6151
R1886 B.n637 B.n634 10.6151
R1887 B.n634 B.n633 10.6151
R1888 B.n633 B.n630 10.6151
R1889 B.n628 B.n625 10.6151
R1890 B.n625 B.n624 10.6151
R1891 B.n624 B.n621 10.6151
R1892 B.n621 B.n620 10.6151
R1893 B.n620 B.n617 10.6151
R1894 B.n617 B.n616 10.6151
R1895 B.n616 B.n613 10.6151
R1896 B.n613 B.n612 10.6151
R1897 B.n612 B.n609 10.6151
R1898 B.n609 B.n608 10.6151
R1899 B.n608 B.n605 10.6151
R1900 B.n605 B.n604 10.6151
R1901 B.n604 B.n601 10.6151
R1902 B.n601 B.n600 10.6151
R1903 B.n600 B.n597 10.6151
R1904 B.n597 B.n596 10.6151
R1905 B.n596 B.n593 10.6151
R1906 B.n593 B.n592 10.6151
R1907 B.n592 B.n589 10.6151
R1908 B.n589 B.n588 10.6151
R1909 B.n588 B.n585 10.6151
R1910 B.n585 B.n584 10.6151
R1911 B.n584 B.n581 10.6151
R1912 B.n581 B.n580 10.6151
R1913 B.n580 B.n577 10.6151
R1914 B.n577 B.n576 10.6151
R1915 B.n576 B.n573 10.6151
R1916 B.n573 B.n572 10.6151
R1917 B.n572 B.n569 10.6151
R1918 B.n569 B.n568 10.6151
R1919 B.n568 B.n565 10.6151
R1920 B.n565 B.n564 10.6151
R1921 B.n564 B.n561 10.6151
R1922 B.n561 B.n560 10.6151
R1923 B.n560 B.n557 10.6151
R1924 B.n557 B.n556 10.6151
R1925 B.n556 B.n553 10.6151
R1926 B.n553 B.n552 10.6151
R1927 B.n552 B.n549 10.6151
R1928 B.n549 B.n548 10.6151
R1929 B.n548 B.n545 10.6151
R1930 B.n545 B.n544 10.6151
R1931 B.n544 B.n541 10.6151
R1932 B.n541 B.n540 10.6151
R1933 B.n540 B.n537 10.6151
R1934 B.n537 B.n536 10.6151
R1935 B.n536 B.n534 10.6151
R1936 B.n747 B.n746 10.6151
R1937 B.n747 B.n467 10.6151
R1938 B.n757 B.n467 10.6151
R1939 B.n758 B.n757 10.6151
R1940 B.n759 B.n758 10.6151
R1941 B.n759 B.n459 10.6151
R1942 B.n768 B.n459 10.6151
R1943 B.n769 B.n768 10.6151
R1944 B.n770 B.n769 10.6151
R1945 B.n770 B.n451 10.6151
R1946 B.n780 B.n451 10.6151
R1947 B.n781 B.n780 10.6151
R1948 B.n782 B.n781 10.6151
R1949 B.n782 B.n443 10.6151
R1950 B.n792 B.n443 10.6151
R1951 B.n793 B.n792 10.6151
R1952 B.n794 B.n793 10.6151
R1953 B.n794 B.n435 10.6151
R1954 B.n804 B.n435 10.6151
R1955 B.n805 B.n804 10.6151
R1956 B.n806 B.n805 10.6151
R1957 B.n806 B.n427 10.6151
R1958 B.n816 B.n427 10.6151
R1959 B.n817 B.n816 10.6151
R1960 B.n818 B.n817 10.6151
R1961 B.n818 B.n419 10.6151
R1962 B.n828 B.n419 10.6151
R1963 B.n829 B.n828 10.6151
R1964 B.n830 B.n829 10.6151
R1965 B.n830 B.n411 10.6151
R1966 B.n840 B.n411 10.6151
R1967 B.n841 B.n840 10.6151
R1968 B.n842 B.n841 10.6151
R1969 B.n842 B.n403 10.6151
R1970 B.n852 B.n403 10.6151
R1971 B.n853 B.n852 10.6151
R1972 B.n854 B.n853 10.6151
R1973 B.n854 B.n395 10.6151
R1974 B.n864 B.n395 10.6151
R1975 B.n865 B.n864 10.6151
R1976 B.n866 B.n865 10.6151
R1977 B.n866 B.n387 10.6151
R1978 B.n876 B.n387 10.6151
R1979 B.n877 B.n876 10.6151
R1980 B.n878 B.n877 10.6151
R1981 B.n878 B.n379 10.6151
R1982 B.n888 B.n379 10.6151
R1983 B.n889 B.n888 10.6151
R1984 B.n890 B.n889 10.6151
R1985 B.n890 B.n371 10.6151
R1986 B.n901 B.n371 10.6151
R1987 B.n902 B.n901 10.6151
R1988 B.n903 B.n902 10.6151
R1989 B.n903 B.n0 10.6151
R1990 B.n1089 B.n1 10.6151
R1991 B.n1089 B.n1088 10.6151
R1992 B.n1088 B.n1087 10.6151
R1993 B.n1087 B.n10 10.6151
R1994 B.n1081 B.n10 10.6151
R1995 B.n1081 B.n1080 10.6151
R1996 B.n1080 B.n1079 10.6151
R1997 B.n1079 B.n17 10.6151
R1998 B.n1073 B.n17 10.6151
R1999 B.n1073 B.n1072 10.6151
R2000 B.n1072 B.n1071 10.6151
R2001 B.n1071 B.n24 10.6151
R2002 B.n1065 B.n24 10.6151
R2003 B.n1065 B.n1064 10.6151
R2004 B.n1064 B.n1063 10.6151
R2005 B.n1063 B.n31 10.6151
R2006 B.n1057 B.n31 10.6151
R2007 B.n1057 B.n1056 10.6151
R2008 B.n1056 B.n1055 10.6151
R2009 B.n1055 B.n38 10.6151
R2010 B.n1049 B.n38 10.6151
R2011 B.n1049 B.n1048 10.6151
R2012 B.n1048 B.n1047 10.6151
R2013 B.n1047 B.n45 10.6151
R2014 B.n1041 B.n45 10.6151
R2015 B.n1041 B.n1040 10.6151
R2016 B.n1040 B.n1039 10.6151
R2017 B.n1039 B.n52 10.6151
R2018 B.n1033 B.n52 10.6151
R2019 B.n1033 B.n1032 10.6151
R2020 B.n1032 B.n1031 10.6151
R2021 B.n1031 B.n59 10.6151
R2022 B.n1025 B.n59 10.6151
R2023 B.n1025 B.n1024 10.6151
R2024 B.n1024 B.n1023 10.6151
R2025 B.n1023 B.n66 10.6151
R2026 B.n1017 B.n66 10.6151
R2027 B.n1017 B.n1016 10.6151
R2028 B.n1016 B.n1015 10.6151
R2029 B.n1015 B.n73 10.6151
R2030 B.n1009 B.n73 10.6151
R2031 B.n1009 B.n1008 10.6151
R2032 B.n1008 B.n1007 10.6151
R2033 B.n1007 B.n80 10.6151
R2034 B.n1001 B.n80 10.6151
R2035 B.n1001 B.n1000 10.6151
R2036 B.n1000 B.n999 10.6151
R2037 B.n999 B.n87 10.6151
R2038 B.n994 B.n87 10.6151
R2039 B.n994 B.n993 10.6151
R2040 B.n993 B.n992 10.6151
R2041 B.n992 B.n94 10.6151
R2042 B.n986 B.n94 10.6151
R2043 B.n986 B.n985 10.6151
R2044 B.n252 B.n161 9.36635
R2045 B.n275 B.n158 9.36635
R2046 B.n651 B.n650 9.36635
R2047 B.n629 B.n628 9.36635
R2048 B.t4 B.n405 8.98697
R2049 B.n1052 B.t19 8.98697
R2050 B.t20 B.n421 3.37043
R2051 B.n1036 B.t3 3.37043
R2052 B.n1095 B.n0 2.81026
R2053 B.n1095 B.n1 2.81026
R2054 B.n441 B.t22 2.24712
R2055 B.t0 B.n1020 2.24712
R2056 B.n255 B.n161 1.24928
R2057 B.n272 B.n158 1.24928
R2058 B.n650 B.n649 1.24928
R2059 B.n630 B.n629 1.24928
R2060 VP.n19 VP.t5 180.448
R2061 VP.n22 VP.n21 161.3
R2062 VP.n23 VP.n18 161.3
R2063 VP.n25 VP.n24 161.3
R2064 VP.n26 VP.n17 161.3
R2065 VP.n28 VP.n27 161.3
R2066 VP.n29 VP.n16 161.3
R2067 VP.n31 VP.n30 161.3
R2068 VP.n32 VP.n15 161.3
R2069 VP.n34 VP.n33 161.3
R2070 VP.n35 VP.n14 161.3
R2071 VP.n37 VP.n36 161.3
R2072 VP.n39 VP.n13 161.3
R2073 VP.n41 VP.n40 161.3
R2074 VP.n42 VP.n12 161.3
R2075 VP.n44 VP.n43 161.3
R2076 VP.n45 VP.n11 161.3
R2077 VP.n82 VP.n0 161.3
R2078 VP.n81 VP.n80 161.3
R2079 VP.n79 VP.n1 161.3
R2080 VP.n78 VP.n77 161.3
R2081 VP.n76 VP.n2 161.3
R2082 VP.n74 VP.n73 161.3
R2083 VP.n72 VP.n3 161.3
R2084 VP.n71 VP.n70 161.3
R2085 VP.n69 VP.n4 161.3
R2086 VP.n68 VP.n67 161.3
R2087 VP.n66 VP.n5 161.3
R2088 VP.n65 VP.n64 161.3
R2089 VP.n63 VP.n6 161.3
R2090 VP.n62 VP.n61 161.3
R2091 VP.n60 VP.n7 161.3
R2092 VP.n59 VP.n58 161.3
R2093 VP.n56 VP.n8 161.3
R2094 VP.n55 VP.n54 161.3
R2095 VP.n53 VP.n9 161.3
R2096 VP.n52 VP.n51 161.3
R2097 VP.n50 VP.n10 161.3
R2098 VP.n5 VP.t4 147.381
R2099 VP.n49 VP.t6 147.381
R2100 VP.n57 VP.t0 147.381
R2101 VP.n75 VP.t9 147.381
R2102 VP.n83 VP.t3 147.381
R2103 VP.n16 VP.t2 147.381
R2104 VP.n46 VP.t1 147.381
R2105 VP.n38 VP.t7 147.381
R2106 VP.n20 VP.t8 147.381
R2107 VP.n49 VP.n48 94.1189
R2108 VP.n84 VP.n83 94.1189
R2109 VP.n47 VP.n46 94.1189
R2110 VP.n20 VP.n19 63.5395
R2111 VP.n63 VP.n62 56.5193
R2112 VP.n70 VP.n69 56.5193
R2113 VP.n33 VP.n32 56.5193
R2114 VP.n26 VP.n25 56.5193
R2115 VP.n48 VP.n47 53.511
R2116 VP.n51 VP.n9 40.979
R2117 VP.n81 VP.n1 40.979
R2118 VP.n44 VP.n12 40.979
R2119 VP.n55 VP.n9 40.0078
R2120 VP.n77 VP.n1 40.0078
R2121 VP.n40 VP.n12 40.0078
R2122 VP.n51 VP.n50 24.4675
R2123 VP.n56 VP.n55 24.4675
R2124 VP.n58 VP.n7 24.4675
R2125 VP.n62 VP.n7 24.4675
R2126 VP.n64 VP.n63 24.4675
R2127 VP.n64 VP.n5 24.4675
R2128 VP.n68 VP.n5 24.4675
R2129 VP.n69 VP.n68 24.4675
R2130 VP.n70 VP.n3 24.4675
R2131 VP.n74 VP.n3 24.4675
R2132 VP.n77 VP.n76 24.4675
R2133 VP.n82 VP.n81 24.4675
R2134 VP.n45 VP.n44 24.4675
R2135 VP.n33 VP.n14 24.4675
R2136 VP.n37 VP.n14 24.4675
R2137 VP.n40 VP.n39 24.4675
R2138 VP.n27 VP.n26 24.4675
R2139 VP.n27 VP.n16 24.4675
R2140 VP.n31 VP.n16 24.4675
R2141 VP.n32 VP.n31 24.4675
R2142 VP.n21 VP.n18 24.4675
R2143 VP.n25 VP.n18 24.4675
R2144 VP.n50 VP.n49 16.6381
R2145 VP.n83 VP.n82 16.6381
R2146 VP.n46 VP.n45 16.6381
R2147 VP.n57 VP.n56 16.1487
R2148 VP.n76 VP.n75 16.1487
R2149 VP.n39 VP.n38 16.1487
R2150 VP.n22 VP.n19 9.31187
R2151 VP.n58 VP.n57 8.31928
R2152 VP.n75 VP.n74 8.31928
R2153 VP.n38 VP.n37 8.31928
R2154 VP.n21 VP.n20 8.31928
R2155 VP.n47 VP.n11 0.278367
R2156 VP.n48 VP.n10 0.278367
R2157 VP.n84 VP.n0 0.278367
R2158 VP.n23 VP.n22 0.189894
R2159 VP.n24 VP.n23 0.189894
R2160 VP.n24 VP.n17 0.189894
R2161 VP.n28 VP.n17 0.189894
R2162 VP.n29 VP.n28 0.189894
R2163 VP.n30 VP.n29 0.189894
R2164 VP.n30 VP.n15 0.189894
R2165 VP.n34 VP.n15 0.189894
R2166 VP.n35 VP.n34 0.189894
R2167 VP.n36 VP.n35 0.189894
R2168 VP.n36 VP.n13 0.189894
R2169 VP.n41 VP.n13 0.189894
R2170 VP.n42 VP.n41 0.189894
R2171 VP.n43 VP.n42 0.189894
R2172 VP.n43 VP.n11 0.189894
R2173 VP.n52 VP.n10 0.189894
R2174 VP.n53 VP.n52 0.189894
R2175 VP.n54 VP.n53 0.189894
R2176 VP.n54 VP.n8 0.189894
R2177 VP.n59 VP.n8 0.189894
R2178 VP.n60 VP.n59 0.189894
R2179 VP.n61 VP.n60 0.189894
R2180 VP.n61 VP.n6 0.189894
R2181 VP.n65 VP.n6 0.189894
R2182 VP.n66 VP.n65 0.189894
R2183 VP.n67 VP.n66 0.189894
R2184 VP.n67 VP.n4 0.189894
R2185 VP.n71 VP.n4 0.189894
R2186 VP.n72 VP.n71 0.189894
R2187 VP.n73 VP.n72 0.189894
R2188 VP.n73 VP.n2 0.189894
R2189 VP.n78 VP.n2 0.189894
R2190 VP.n79 VP.n78 0.189894
R2191 VP.n80 VP.n79 0.189894
R2192 VP.n80 VP.n0 0.189894
R2193 VP VP.n84 0.153454
R2194 VDD1.n1 VDD1.t4 65.233
R2195 VDD1.n3 VDD1.t3 65.2329
R2196 VDD1.n5 VDD1.n4 63.2184
R2197 VDD1.n1 VDD1.n0 61.5477
R2198 VDD1.n7 VDD1.n6 61.5475
R2199 VDD1.n3 VDD1.n2 61.5475
R2200 VDD1.n7 VDD1.n5 48.7186
R2201 VDD1 VDD1.n7 1.6686
R2202 VDD1.n6 VDD1.t2 1.38415
R2203 VDD1.n6 VDD1.t8 1.38415
R2204 VDD1.n0 VDD1.t1 1.38415
R2205 VDD1.n0 VDD1.t7 1.38415
R2206 VDD1.n4 VDD1.t0 1.38415
R2207 VDD1.n4 VDD1.t6 1.38415
R2208 VDD1.n2 VDD1.t9 1.38415
R2209 VDD1.n2 VDD1.t5 1.38415
R2210 VDD1 VDD1.n1 0.634121
R2211 VDD1.n5 VDD1.n3 0.520585
C0 VDD1 VDD2 2.00449f
C1 VTAIL VP 12.7946f
C2 VN VDD2 12.348599f
C3 VDD1 VN 0.15262f
C4 VP VDD2 0.550474f
C5 VDD1 VP 12.7421f
C6 VP VN 8.44139f
C7 VTAIL VDD2 11.541f
C8 VDD1 VTAIL 11.492701f
C9 VTAIL VN 12.7802f
C10 VDD2 B 7.317884f
C11 VDD1 B 7.28688f
C12 VTAIL B 8.912727f
C13 VN B 17.10482f
C14 VP B 15.570601f
C15 VDD1.t4 B 3.14577f
C16 VDD1.t1 B 0.271885f
C17 VDD1.t7 B 0.271885f
C18 VDD1.n0 B 2.45272f
C19 VDD1.n1 B 0.85483f
C20 VDD1.t3 B 3.14576f
C21 VDD1.t9 B 0.271885f
C22 VDD1.t5 B 0.271885f
C23 VDD1.n2 B 2.45272f
C24 VDD1.n3 B 0.847122f
C25 VDD1.t0 B 0.271885f
C26 VDD1.t6 B 0.271885f
C27 VDD1.n4 B 2.46628f
C28 VDD1.n5 B 2.91373f
C29 VDD1.t2 B 0.271885f
C30 VDD1.t8 B 0.271885f
C31 VDD1.n6 B 2.45271f
C32 VDD1.n7 B 3.11495f
C33 VP.n0 B 0.03002f
C34 VP.t3 B 2.08703f
C35 VP.n1 B 0.018416f
C36 VP.n2 B 0.02277f
C37 VP.t9 B 2.08703f
C38 VP.n3 B 0.042438f
C39 VP.n4 B 0.02277f
C40 VP.t4 B 2.08703f
C41 VP.n5 B 0.754708f
C42 VP.n6 B 0.02277f
C43 VP.n7 B 0.042438f
C44 VP.n8 B 0.02277f
C45 VP.t0 B 2.08703f
C46 VP.n9 B 0.018416f
C47 VP.n10 B 0.03002f
C48 VP.t6 B 2.08703f
C49 VP.n11 B 0.03002f
C50 VP.t1 B 2.08703f
C51 VP.n12 B 0.018416f
C52 VP.n13 B 0.02277f
C53 VP.t7 B 2.08703f
C54 VP.n14 B 0.042438f
C55 VP.n15 B 0.02277f
C56 VP.t2 B 2.08703f
C57 VP.n16 B 0.754708f
C58 VP.n17 B 0.02277f
C59 VP.n18 B 0.042438f
C60 VP.t5 B 2.24519f
C61 VP.n19 B 0.781896f
C62 VP.t8 B 2.08703f
C63 VP.n20 B 0.791291f
C64 VP.n21 B 0.02861f
C65 VP.n22 B 0.196953f
C66 VP.n23 B 0.02277f
C67 VP.n24 B 0.02277f
C68 VP.n25 B 0.027849f
C69 VP.n26 B 0.038636f
C70 VP.n27 B 0.042438f
C71 VP.n28 B 0.02277f
C72 VP.n29 B 0.02277f
C73 VP.n30 B 0.02277f
C74 VP.n31 B 0.042438f
C75 VP.n32 B 0.038636f
C76 VP.n33 B 0.027849f
C77 VP.n34 B 0.02277f
C78 VP.n35 B 0.02277f
C79 VP.n36 B 0.02277f
C80 VP.n37 B 0.02861f
C81 VP.n38 B 0.733222f
C82 VP.n39 B 0.035314f
C83 VP.n40 B 0.045368f
C84 VP.n41 B 0.02277f
C85 VP.n42 B 0.02277f
C86 VP.n43 B 0.02277f
C87 VP.n44 B 0.04514f
C88 VP.n45 B 0.035734f
C89 VP.n46 B 0.810197f
C90 VP.n47 B 1.39203f
C91 VP.n48 B 1.40733f
C92 VP.n49 B 0.810197f
C93 VP.n50 B 0.035734f
C94 VP.n51 B 0.04514f
C95 VP.n52 B 0.02277f
C96 VP.n53 B 0.02277f
C97 VP.n54 B 0.02277f
C98 VP.n55 B 0.045368f
C99 VP.n56 B 0.035314f
C100 VP.n57 B 0.733222f
C101 VP.n58 B 0.02861f
C102 VP.n59 B 0.02277f
C103 VP.n60 B 0.02277f
C104 VP.n61 B 0.02277f
C105 VP.n62 B 0.027849f
C106 VP.n63 B 0.038636f
C107 VP.n64 B 0.042438f
C108 VP.n65 B 0.02277f
C109 VP.n66 B 0.02277f
C110 VP.n67 B 0.02277f
C111 VP.n68 B 0.042438f
C112 VP.n69 B 0.038636f
C113 VP.n70 B 0.027849f
C114 VP.n71 B 0.02277f
C115 VP.n72 B 0.02277f
C116 VP.n73 B 0.02277f
C117 VP.n74 B 0.02861f
C118 VP.n75 B 0.733222f
C119 VP.n76 B 0.035314f
C120 VP.n77 B 0.045368f
C121 VP.n78 B 0.02277f
C122 VP.n79 B 0.02277f
C123 VP.n80 B 0.02277f
C124 VP.n81 B 0.04514f
C125 VP.n82 B 0.035734f
C126 VP.n83 B 0.810197f
C127 VP.n84 B 0.031232f
C128 VTAIL.t12 B 0.273817f
C129 VTAIL.t19 B 0.273817f
C130 VTAIL.n0 B 2.39868f
C131 VTAIL.n1 B 0.501117f
C132 VTAIL.t1 B 3.05954f
C133 VTAIL.n2 B 0.62739f
C134 VTAIL.t4 B 0.273817f
C135 VTAIL.t7 B 0.273817f
C136 VTAIL.n3 B 2.39868f
C137 VTAIL.n4 B 0.594611f
C138 VTAIL.t8 B 0.273817f
C139 VTAIL.t6 B 0.273817f
C140 VTAIL.n5 B 2.39868f
C141 VTAIL.n6 B 2.06563f
C142 VTAIL.t15 B 0.273817f
C143 VTAIL.t16 B 0.273817f
C144 VTAIL.n7 B 2.39868f
C145 VTAIL.n8 B 2.06562f
C146 VTAIL.t11 B 0.273817f
C147 VTAIL.t18 B 0.273817f
C148 VTAIL.n9 B 2.39868f
C149 VTAIL.n10 B 0.594607f
C150 VTAIL.t14 B 3.05956f
C151 VTAIL.n11 B 0.627368f
C152 VTAIL.t9 B 0.273817f
C153 VTAIL.t2 B 0.273817f
C154 VTAIL.n12 B 2.39868f
C155 VTAIL.n13 B 0.541471f
C156 VTAIL.t5 B 0.273817f
C157 VTAIL.t3 B 0.273817f
C158 VTAIL.n14 B 2.39868f
C159 VTAIL.n15 B 0.594607f
C160 VTAIL.t0 B 3.05954f
C161 VTAIL.n16 B 1.97195f
C162 VTAIL.t10 B 3.05954f
C163 VTAIL.n17 B 1.97195f
C164 VTAIL.t13 B 0.273817f
C165 VTAIL.t17 B 0.273817f
C166 VTAIL.n18 B 2.39868f
C167 VTAIL.n19 B 0.45538f
C168 VDD2.t4 B 3.10827f
C169 VDD2.t3 B 0.268644f
C170 VDD2.t5 B 0.268644f
C171 VDD2.n0 B 2.42349f
C172 VDD2.n1 B 0.837026f
C173 VDD2.t1 B 0.268644f
C174 VDD2.t6 B 0.268644f
C175 VDD2.n2 B 2.43689f
C176 VDD2.n3 B 2.7654f
C177 VDD2.t9 B 3.09267f
C178 VDD2.n4 B 3.03947f
C179 VDD2.t0 B 0.268644f
C180 VDD2.t7 B 0.268644f
C181 VDD2.n5 B 2.42349f
C182 VDD2.n6 B 0.417853f
C183 VDD2.t2 B 0.268644f
C184 VDD2.t8 B 0.268644f
C185 VDD2.n7 B 2.43685f
C186 VN.n0 B 0.029638f
C187 VN.t9 B 2.06046f
C188 VN.n1 B 0.018181f
C189 VN.n2 B 0.02248f
C190 VN.t2 B 2.06046f
C191 VN.n3 B 0.041898f
C192 VN.n4 B 0.02248f
C193 VN.t6 B 2.06046f
C194 VN.n5 B 0.745099f
C195 VN.n6 B 0.02248f
C196 VN.n7 B 0.041898f
C197 VN.t7 B 2.21661f
C198 VN.n8 B 0.771941f
C199 VN.t0 B 2.06046f
C200 VN.n9 B 0.781216f
C201 VN.n10 B 0.028246f
C202 VN.n11 B 0.194446f
C203 VN.n12 B 0.02248f
C204 VN.n13 B 0.02248f
C205 VN.n14 B 0.027495f
C206 VN.n15 B 0.038144f
C207 VN.n16 B 0.041898f
C208 VN.n17 B 0.02248f
C209 VN.n18 B 0.02248f
C210 VN.n19 B 0.02248f
C211 VN.n20 B 0.041898f
C212 VN.n21 B 0.038144f
C213 VN.n22 B 0.027495f
C214 VN.n23 B 0.02248f
C215 VN.n24 B 0.02248f
C216 VN.n25 B 0.02248f
C217 VN.n26 B 0.028246f
C218 VN.n27 B 0.723887f
C219 VN.n28 B 0.034865f
C220 VN.n29 B 0.04479f
C221 VN.n30 B 0.02248f
C222 VN.n31 B 0.02248f
C223 VN.n32 B 0.02248f
C224 VN.n33 B 0.044565f
C225 VN.n34 B 0.035279f
C226 VN.n35 B 0.799882f
C227 VN.n36 B 0.030835f
C228 VN.n37 B 0.029638f
C229 VN.t4 B 2.06046f
C230 VN.n38 B 0.018181f
C231 VN.n39 B 0.02248f
C232 VN.t3 B 2.06046f
C233 VN.n40 B 0.041898f
C234 VN.n41 B 0.02248f
C235 VN.t8 B 2.06046f
C236 VN.n42 B 0.745099f
C237 VN.n43 B 0.02248f
C238 VN.n44 B 0.041898f
C239 VN.t5 B 2.21661f
C240 VN.n45 B 0.771941f
C241 VN.t1 B 2.06046f
C242 VN.n46 B 0.781216f
C243 VN.n47 B 0.028246f
C244 VN.n48 B 0.194446f
C245 VN.n49 B 0.02248f
C246 VN.n50 B 0.02248f
C247 VN.n51 B 0.027495f
C248 VN.n52 B 0.038144f
C249 VN.n53 B 0.041898f
C250 VN.n54 B 0.02248f
C251 VN.n55 B 0.02248f
C252 VN.n56 B 0.02248f
C253 VN.n57 B 0.041898f
C254 VN.n58 B 0.038144f
C255 VN.n59 B 0.027495f
C256 VN.n60 B 0.02248f
C257 VN.n61 B 0.02248f
C258 VN.n62 B 0.02248f
C259 VN.n63 B 0.028246f
C260 VN.n64 B 0.723887f
C261 VN.n65 B 0.034865f
C262 VN.n66 B 0.04479f
C263 VN.n67 B 0.02248f
C264 VN.n68 B 0.02248f
C265 VN.n69 B 0.02248f
C266 VN.n70 B 0.044565f
C267 VN.n71 B 0.035279f
C268 VN.n72 B 0.799882f
C269 VN.n73 B 1.38626f
.ends

