* NGSPICE file created from diff_pair_sample_0472.ext - technology: sky130A

.subckt diff_pair_sample_0472 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=2.04725 ps=9.57 w=4.31 l=0.16
X1 VDD1.t4 VP.t1 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=1.0775 ps=4.81 w=4.31 l=0.16
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=0 ps=0 w=4.31 l=0.16
X3 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=0 ps=0 w=4.31 l=0.16
X4 VDD2.t5 VN.t0 VTAIL.t11 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=2.04725 ps=9.57 w=4.31 l=0.16
X5 VDD1.t3 VP.t2 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=1.0775 ps=4.81 w=4.31 l=0.16
X6 VTAIL.t6 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=1.0775 ps=4.81 w=4.31 l=0.16
X7 VDD2.t4 VN.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=1.0775 ps=4.81 w=4.31 l=0.16
X8 VTAIL.t7 VP.t4 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=1.0775 ps=4.81 w=4.31 l=0.16
X9 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=2.04725 ps=9.57 w=4.31 l=0.16
X10 VTAIL.t10 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=1.0775 ps=4.81 w=4.31 l=0.16
X11 VDD2.t1 VN.t4 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=1.0775 ps=4.81 w=4.31 l=0.16
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=0 ps=0 w=4.31 l=0.16
X13 VTAIL.t0 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=1.0775 ps=4.81 w=4.31 l=0.16
X14 VDD1.t0 VP.t5 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0775 pd=4.81 as=2.04725 ps=9.57 w=4.31 l=0.16
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.04725 pd=9.57 as=0 ps=0 w=4.31 l=0.16
R0 VP.n7 VP.t0 906.398
R1 VP.n5 VP.t2 906.398
R2 VP.n0 VP.t1 906.398
R3 VP.n2 VP.t5 906.398
R4 VP.n6 VP.t3 846.514
R5 VP.n1 VP.t4 846.514
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n6 VP.n5 36.5157
R11 VP.n7 VP.n6 36.5157
R12 VP.n1 VP.n0 36.5157
R13 VP.n2 VP.n1 36.5157
R14 VP.n4 VP.n3 34.1217
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VTAIL.n7 VTAIL.t1 64.3335
R18 VTAIL.n10 VTAIL.t3 64.3333
R19 VTAIL.n11 VTAIL.t11 64.3333
R20 VTAIL.n2 VTAIL.t2 64.3333
R21 VTAIL.n9 VTAIL.n8 57.373
R22 VTAIL.n6 VTAIL.n5 57.373
R23 VTAIL.n1 VTAIL.n0 57.3728
R24 VTAIL.n4 VTAIL.n3 57.3728
R25 VTAIL.n6 VTAIL.n4 17.2203
R26 VTAIL.n11 VTAIL.n10 16.6514
R27 VTAIL.n0 VTAIL.t9 6.96106
R28 VTAIL.n0 VTAIL.t10 6.96106
R29 VTAIL.n3 VTAIL.t5 6.96106
R30 VTAIL.n3 VTAIL.t6 6.96106
R31 VTAIL.n8 VTAIL.t4 6.96106
R32 VTAIL.n8 VTAIL.t7 6.96106
R33 VTAIL.n5 VTAIL.t8 6.96106
R34 VTAIL.n5 VTAIL.t0 6.96106
R35 VTAIL.n9 VTAIL.n7 0.75481
R36 VTAIL.n2 VTAIL.n1 0.75481
R37 VTAIL.n7 VTAIL.n6 0.569465
R38 VTAIL.n10 VTAIL.n9 0.569465
R39 VTAIL.n4 VTAIL.n2 0.569465
R40 VTAIL VTAIL.n11 0.369034
R41 VTAIL VTAIL.n1 0.200931
R42 VDD1 VDD1.t4 81.4972
R43 VDD1.n1 VDD1.t3 81.3835
R44 VDD1.n1 VDD1.n0 74.1384
R45 VDD1.n3 VDD1.n2 74.0516
R46 VDD1.n3 VDD1.n1 30.1474
R47 VDD1.n2 VDD1.t1 6.96106
R48 VDD1.n2 VDD1.t0 6.96106
R49 VDD1.n0 VDD1.t2 6.96106
R50 VDD1.n0 VDD1.t5 6.96106
R51 VDD1 VDD1.n3 0.0845517
R52 B.n194 B.t10 900.606
R53 B.n203 B.t14 900.606
R54 B.n60 B.t6 900.606
R55 B.n58 B.t17 900.606
R56 B.n380 B.n379 585
R57 B.n154 B.n57 585
R58 B.n153 B.n152 585
R59 B.n151 B.n150 585
R60 B.n149 B.n148 585
R61 B.n147 B.n146 585
R62 B.n145 B.n144 585
R63 B.n143 B.n142 585
R64 B.n141 B.n140 585
R65 B.n139 B.n138 585
R66 B.n137 B.n136 585
R67 B.n135 B.n134 585
R68 B.n133 B.n132 585
R69 B.n131 B.n130 585
R70 B.n129 B.n128 585
R71 B.n127 B.n126 585
R72 B.n125 B.n124 585
R73 B.n123 B.n122 585
R74 B.n121 B.n120 585
R75 B.n118 B.n117 585
R76 B.n116 B.n115 585
R77 B.n114 B.n113 585
R78 B.n112 B.n111 585
R79 B.n110 B.n109 585
R80 B.n108 B.n107 585
R81 B.n106 B.n105 585
R82 B.n104 B.n103 585
R83 B.n102 B.n101 585
R84 B.n100 B.n99 585
R85 B.n97 B.n96 585
R86 B.n95 B.n94 585
R87 B.n93 B.n92 585
R88 B.n91 B.n90 585
R89 B.n89 B.n88 585
R90 B.n87 B.n86 585
R91 B.n85 B.n84 585
R92 B.n83 B.n82 585
R93 B.n81 B.n80 585
R94 B.n79 B.n78 585
R95 B.n77 B.n76 585
R96 B.n75 B.n74 585
R97 B.n73 B.n72 585
R98 B.n71 B.n70 585
R99 B.n69 B.n68 585
R100 B.n67 B.n66 585
R101 B.n65 B.n64 585
R102 B.n63 B.n62 585
R103 B.n32 B.n31 585
R104 B.n378 B.n33 585
R105 B.n383 B.n33 585
R106 B.n377 B.n376 585
R107 B.n376 B.n29 585
R108 B.n375 B.n28 585
R109 B.n389 B.n28 585
R110 B.n374 B.n27 585
R111 B.n390 B.n27 585
R112 B.n373 B.n26 585
R113 B.n391 B.n26 585
R114 B.n372 B.n371 585
R115 B.n371 B.n22 585
R116 B.n370 B.n21 585
R117 B.n397 B.n21 585
R118 B.n369 B.n20 585
R119 B.n398 B.n20 585
R120 B.n368 B.n19 585
R121 B.n399 B.n19 585
R122 B.n367 B.n366 585
R123 B.n366 B.n18 585
R124 B.n365 B.n14 585
R125 B.n405 B.n14 585
R126 B.n364 B.n13 585
R127 B.n406 B.n13 585
R128 B.n363 B.n12 585
R129 B.n407 B.n12 585
R130 B.n362 B.n361 585
R131 B.n361 B.n11 585
R132 B.n360 B.n7 585
R133 B.n413 B.n7 585
R134 B.n359 B.n6 585
R135 B.n414 B.n6 585
R136 B.n358 B.n5 585
R137 B.n415 B.n5 585
R138 B.n357 B.n356 585
R139 B.n356 B.n4 585
R140 B.n355 B.n155 585
R141 B.n355 B.n354 585
R142 B.n344 B.n156 585
R143 B.n347 B.n156 585
R144 B.n346 B.n345 585
R145 B.n348 B.n346 585
R146 B.n343 B.n160 585
R147 B.n163 B.n160 585
R148 B.n342 B.n341 585
R149 B.n341 B.n340 585
R150 B.n162 B.n161 585
R151 B.n333 B.n162 585
R152 B.n332 B.n331 585
R153 B.n334 B.n332 585
R154 B.n330 B.n168 585
R155 B.n168 B.n167 585
R156 B.n329 B.n328 585
R157 B.n328 B.n327 585
R158 B.n170 B.n169 585
R159 B.n171 B.n170 585
R160 B.n320 B.n319 585
R161 B.n321 B.n320 585
R162 B.n318 B.n176 585
R163 B.n176 B.n175 585
R164 B.n317 B.n316 585
R165 B.n316 B.n315 585
R166 B.n178 B.n177 585
R167 B.n179 B.n178 585
R168 B.n308 B.n307 585
R169 B.n309 B.n308 585
R170 B.n182 B.n181 585
R171 B.n215 B.n214 585
R172 B.n216 B.n212 585
R173 B.n212 B.n183 585
R174 B.n218 B.n217 585
R175 B.n220 B.n211 585
R176 B.n223 B.n222 585
R177 B.n224 B.n210 585
R178 B.n226 B.n225 585
R179 B.n228 B.n209 585
R180 B.n231 B.n230 585
R181 B.n232 B.n208 585
R182 B.n234 B.n233 585
R183 B.n236 B.n207 585
R184 B.n239 B.n238 585
R185 B.n240 B.n206 585
R186 B.n242 B.n241 585
R187 B.n244 B.n205 585
R188 B.n247 B.n246 585
R189 B.n248 B.n202 585
R190 B.n251 B.n250 585
R191 B.n253 B.n201 585
R192 B.n256 B.n255 585
R193 B.n257 B.n200 585
R194 B.n259 B.n258 585
R195 B.n261 B.n199 585
R196 B.n264 B.n263 585
R197 B.n265 B.n198 585
R198 B.n267 B.n266 585
R199 B.n269 B.n197 585
R200 B.n272 B.n271 585
R201 B.n273 B.n193 585
R202 B.n275 B.n274 585
R203 B.n277 B.n192 585
R204 B.n280 B.n279 585
R205 B.n281 B.n191 585
R206 B.n283 B.n282 585
R207 B.n285 B.n190 585
R208 B.n288 B.n287 585
R209 B.n289 B.n189 585
R210 B.n291 B.n290 585
R211 B.n293 B.n188 585
R212 B.n296 B.n295 585
R213 B.n297 B.n187 585
R214 B.n299 B.n298 585
R215 B.n301 B.n186 585
R216 B.n302 B.n185 585
R217 B.n305 B.n304 585
R218 B.n306 B.n184 585
R219 B.n184 B.n183 585
R220 B.n311 B.n310 585
R221 B.n310 B.n309 585
R222 B.n312 B.n180 585
R223 B.n180 B.n179 585
R224 B.n314 B.n313 585
R225 B.n315 B.n314 585
R226 B.n174 B.n173 585
R227 B.n175 B.n174 585
R228 B.n323 B.n322 585
R229 B.n322 B.n321 585
R230 B.n324 B.n172 585
R231 B.n172 B.n171 585
R232 B.n326 B.n325 585
R233 B.n327 B.n326 585
R234 B.n166 B.n165 585
R235 B.n167 B.n166 585
R236 B.n336 B.n335 585
R237 B.n335 B.n334 585
R238 B.n337 B.n164 585
R239 B.n333 B.n164 585
R240 B.n339 B.n338 585
R241 B.n340 B.n339 585
R242 B.n159 B.n158 585
R243 B.n163 B.n159 585
R244 B.n350 B.n349 585
R245 B.n349 B.n348 585
R246 B.n351 B.n157 585
R247 B.n347 B.n157 585
R248 B.n353 B.n352 585
R249 B.n354 B.n353 585
R250 B.n2 B.n0 585
R251 B.n4 B.n2 585
R252 B.n3 B.n1 585
R253 B.n414 B.n3 585
R254 B.n412 B.n411 585
R255 B.n413 B.n412 585
R256 B.n410 B.n8 585
R257 B.n11 B.n8 585
R258 B.n409 B.n408 585
R259 B.n408 B.n407 585
R260 B.n10 B.n9 585
R261 B.n406 B.n10 585
R262 B.n404 B.n403 585
R263 B.n405 B.n404 585
R264 B.n402 B.n15 585
R265 B.n18 B.n15 585
R266 B.n401 B.n400 585
R267 B.n400 B.n399 585
R268 B.n17 B.n16 585
R269 B.n398 B.n17 585
R270 B.n396 B.n395 585
R271 B.n397 B.n396 585
R272 B.n394 B.n23 585
R273 B.n23 B.n22 585
R274 B.n393 B.n392 585
R275 B.n392 B.n391 585
R276 B.n25 B.n24 585
R277 B.n390 B.n25 585
R278 B.n388 B.n387 585
R279 B.n389 B.n388 585
R280 B.n386 B.n30 585
R281 B.n30 B.n29 585
R282 B.n385 B.n384 585
R283 B.n384 B.n383 585
R284 B.n417 B.n416 585
R285 B.n416 B.n415 585
R286 B.n310 B.n182 444.452
R287 B.n384 B.n32 444.452
R288 B.n308 B.n184 444.452
R289 B.n380 B.n33 444.452
R290 B.n382 B.n381 256.663
R291 B.n382 B.n56 256.663
R292 B.n382 B.n55 256.663
R293 B.n382 B.n54 256.663
R294 B.n382 B.n53 256.663
R295 B.n382 B.n52 256.663
R296 B.n382 B.n51 256.663
R297 B.n382 B.n50 256.663
R298 B.n382 B.n49 256.663
R299 B.n382 B.n48 256.663
R300 B.n382 B.n47 256.663
R301 B.n382 B.n46 256.663
R302 B.n382 B.n45 256.663
R303 B.n382 B.n44 256.663
R304 B.n382 B.n43 256.663
R305 B.n382 B.n42 256.663
R306 B.n382 B.n41 256.663
R307 B.n382 B.n40 256.663
R308 B.n382 B.n39 256.663
R309 B.n382 B.n38 256.663
R310 B.n382 B.n37 256.663
R311 B.n382 B.n36 256.663
R312 B.n382 B.n35 256.663
R313 B.n382 B.n34 256.663
R314 B.n213 B.n183 256.663
R315 B.n219 B.n183 256.663
R316 B.n221 B.n183 256.663
R317 B.n227 B.n183 256.663
R318 B.n229 B.n183 256.663
R319 B.n235 B.n183 256.663
R320 B.n237 B.n183 256.663
R321 B.n243 B.n183 256.663
R322 B.n245 B.n183 256.663
R323 B.n252 B.n183 256.663
R324 B.n254 B.n183 256.663
R325 B.n260 B.n183 256.663
R326 B.n262 B.n183 256.663
R327 B.n268 B.n183 256.663
R328 B.n270 B.n183 256.663
R329 B.n276 B.n183 256.663
R330 B.n278 B.n183 256.663
R331 B.n284 B.n183 256.663
R332 B.n286 B.n183 256.663
R333 B.n292 B.n183 256.663
R334 B.n294 B.n183 256.663
R335 B.n300 B.n183 256.663
R336 B.n303 B.n183 256.663
R337 B.n310 B.n180 163.367
R338 B.n314 B.n180 163.367
R339 B.n314 B.n174 163.367
R340 B.n322 B.n174 163.367
R341 B.n322 B.n172 163.367
R342 B.n326 B.n172 163.367
R343 B.n326 B.n166 163.367
R344 B.n335 B.n166 163.367
R345 B.n335 B.n164 163.367
R346 B.n339 B.n164 163.367
R347 B.n339 B.n159 163.367
R348 B.n349 B.n159 163.367
R349 B.n349 B.n157 163.367
R350 B.n353 B.n157 163.367
R351 B.n353 B.n2 163.367
R352 B.n416 B.n2 163.367
R353 B.n416 B.n3 163.367
R354 B.n412 B.n3 163.367
R355 B.n412 B.n8 163.367
R356 B.n408 B.n8 163.367
R357 B.n408 B.n10 163.367
R358 B.n404 B.n10 163.367
R359 B.n404 B.n15 163.367
R360 B.n400 B.n15 163.367
R361 B.n400 B.n17 163.367
R362 B.n396 B.n17 163.367
R363 B.n396 B.n23 163.367
R364 B.n392 B.n23 163.367
R365 B.n392 B.n25 163.367
R366 B.n388 B.n25 163.367
R367 B.n388 B.n30 163.367
R368 B.n384 B.n30 163.367
R369 B.n214 B.n212 163.367
R370 B.n218 B.n212 163.367
R371 B.n222 B.n220 163.367
R372 B.n226 B.n210 163.367
R373 B.n230 B.n228 163.367
R374 B.n234 B.n208 163.367
R375 B.n238 B.n236 163.367
R376 B.n242 B.n206 163.367
R377 B.n246 B.n244 163.367
R378 B.n251 B.n202 163.367
R379 B.n255 B.n253 163.367
R380 B.n259 B.n200 163.367
R381 B.n263 B.n261 163.367
R382 B.n267 B.n198 163.367
R383 B.n271 B.n269 163.367
R384 B.n275 B.n193 163.367
R385 B.n279 B.n277 163.367
R386 B.n283 B.n191 163.367
R387 B.n287 B.n285 163.367
R388 B.n291 B.n189 163.367
R389 B.n295 B.n293 163.367
R390 B.n299 B.n187 163.367
R391 B.n302 B.n301 163.367
R392 B.n304 B.n184 163.367
R393 B.n308 B.n178 163.367
R394 B.n316 B.n178 163.367
R395 B.n316 B.n176 163.367
R396 B.n320 B.n176 163.367
R397 B.n320 B.n170 163.367
R398 B.n328 B.n170 163.367
R399 B.n328 B.n168 163.367
R400 B.n332 B.n168 163.367
R401 B.n332 B.n162 163.367
R402 B.n341 B.n162 163.367
R403 B.n341 B.n160 163.367
R404 B.n346 B.n160 163.367
R405 B.n346 B.n156 163.367
R406 B.n355 B.n156 163.367
R407 B.n356 B.n355 163.367
R408 B.n356 B.n5 163.367
R409 B.n6 B.n5 163.367
R410 B.n7 B.n6 163.367
R411 B.n361 B.n7 163.367
R412 B.n361 B.n12 163.367
R413 B.n13 B.n12 163.367
R414 B.n14 B.n13 163.367
R415 B.n366 B.n14 163.367
R416 B.n366 B.n19 163.367
R417 B.n20 B.n19 163.367
R418 B.n21 B.n20 163.367
R419 B.n371 B.n21 163.367
R420 B.n371 B.n26 163.367
R421 B.n27 B.n26 163.367
R422 B.n28 B.n27 163.367
R423 B.n376 B.n28 163.367
R424 B.n376 B.n33 163.367
R425 B.n64 B.n63 163.367
R426 B.n68 B.n67 163.367
R427 B.n72 B.n71 163.367
R428 B.n76 B.n75 163.367
R429 B.n80 B.n79 163.367
R430 B.n84 B.n83 163.367
R431 B.n88 B.n87 163.367
R432 B.n92 B.n91 163.367
R433 B.n96 B.n95 163.367
R434 B.n101 B.n100 163.367
R435 B.n105 B.n104 163.367
R436 B.n109 B.n108 163.367
R437 B.n113 B.n112 163.367
R438 B.n117 B.n116 163.367
R439 B.n122 B.n121 163.367
R440 B.n126 B.n125 163.367
R441 B.n130 B.n129 163.367
R442 B.n134 B.n133 163.367
R443 B.n138 B.n137 163.367
R444 B.n142 B.n141 163.367
R445 B.n146 B.n145 163.367
R446 B.n150 B.n149 163.367
R447 B.n152 B.n57 163.367
R448 B.n309 B.n183 131.977
R449 B.n383 B.n382 131.977
R450 B.n194 B.t13 90.6357
R451 B.n58 B.t18 90.6357
R452 B.n203 B.t16 90.6318
R453 B.n60 B.t8 90.6318
R454 B.n309 B.n179 78.0391
R455 B.n315 B.n179 78.0391
R456 B.n315 B.n175 78.0391
R457 B.n321 B.n175 78.0391
R458 B.n327 B.n171 78.0391
R459 B.n327 B.n167 78.0391
R460 B.n334 B.n167 78.0391
R461 B.n334 B.n333 78.0391
R462 B.n340 B.n163 78.0391
R463 B.n348 B.n347 78.0391
R464 B.n354 B.n4 78.0391
R465 B.n415 B.n4 78.0391
R466 B.n415 B.n414 78.0391
R467 B.n414 B.n413 78.0391
R468 B.n407 B.n11 78.0391
R469 B.n406 B.n405 78.0391
R470 B.n399 B.n18 78.0391
R471 B.n399 B.n398 78.0391
R472 B.n398 B.n397 78.0391
R473 B.n397 B.n22 78.0391
R474 B.n391 B.n390 78.0391
R475 B.n390 B.n389 78.0391
R476 B.n389 B.n29 78.0391
R477 B.n383 B.n29 78.0391
R478 B.n195 B.t12 77.8357
R479 B.n59 B.t19 77.8357
R480 B.n204 B.t15 77.8318
R481 B.n61 B.t9 77.8318
R482 B.n213 B.n182 71.676
R483 B.n219 B.n218 71.676
R484 B.n222 B.n221 71.676
R485 B.n227 B.n226 71.676
R486 B.n230 B.n229 71.676
R487 B.n235 B.n234 71.676
R488 B.n238 B.n237 71.676
R489 B.n243 B.n242 71.676
R490 B.n246 B.n245 71.676
R491 B.n252 B.n251 71.676
R492 B.n255 B.n254 71.676
R493 B.n260 B.n259 71.676
R494 B.n263 B.n262 71.676
R495 B.n268 B.n267 71.676
R496 B.n271 B.n270 71.676
R497 B.n276 B.n275 71.676
R498 B.n279 B.n278 71.676
R499 B.n284 B.n283 71.676
R500 B.n287 B.n286 71.676
R501 B.n292 B.n291 71.676
R502 B.n295 B.n294 71.676
R503 B.n300 B.n299 71.676
R504 B.n303 B.n302 71.676
R505 B.n34 B.n32 71.676
R506 B.n64 B.n35 71.676
R507 B.n68 B.n36 71.676
R508 B.n72 B.n37 71.676
R509 B.n76 B.n38 71.676
R510 B.n80 B.n39 71.676
R511 B.n84 B.n40 71.676
R512 B.n88 B.n41 71.676
R513 B.n92 B.n42 71.676
R514 B.n96 B.n43 71.676
R515 B.n101 B.n44 71.676
R516 B.n105 B.n45 71.676
R517 B.n109 B.n46 71.676
R518 B.n113 B.n47 71.676
R519 B.n117 B.n48 71.676
R520 B.n122 B.n49 71.676
R521 B.n126 B.n50 71.676
R522 B.n130 B.n51 71.676
R523 B.n134 B.n52 71.676
R524 B.n138 B.n53 71.676
R525 B.n142 B.n54 71.676
R526 B.n146 B.n55 71.676
R527 B.n150 B.n56 71.676
R528 B.n381 B.n57 71.676
R529 B.n381 B.n380 71.676
R530 B.n152 B.n56 71.676
R531 B.n149 B.n55 71.676
R532 B.n145 B.n54 71.676
R533 B.n141 B.n53 71.676
R534 B.n137 B.n52 71.676
R535 B.n133 B.n51 71.676
R536 B.n129 B.n50 71.676
R537 B.n125 B.n49 71.676
R538 B.n121 B.n48 71.676
R539 B.n116 B.n47 71.676
R540 B.n112 B.n46 71.676
R541 B.n108 B.n45 71.676
R542 B.n104 B.n44 71.676
R543 B.n100 B.n43 71.676
R544 B.n95 B.n42 71.676
R545 B.n91 B.n41 71.676
R546 B.n87 B.n40 71.676
R547 B.n83 B.n39 71.676
R548 B.n79 B.n38 71.676
R549 B.n75 B.n37 71.676
R550 B.n71 B.n36 71.676
R551 B.n67 B.n35 71.676
R552 B.n63 B.n34 71.676
R553 B.n214 B.n213 71.676
R554 B.n220 B.n219 71.676
R555 B.n221 B.n210 71.676
R556 B.n228 B.n227 71.676
R557 B.n229 B.n208 71.676
R558 B.n236 B.n235 71.676
R559 B.n237 B.n206 71.676
R560 B.n244 B.n243 71.676
R561 B.n245 B.n202 71.676
R562 B.n253 B.n252 71.676
R563 B.n254 B.n200 71.676
R564 B.n261 B.n260 71.676
R565 B.n262 B.n198 71.676
R566 B.n269 B.n268 71.676
R567 B.n270 B.n193 71.676
R568 B.n277 B.n276 71.676
R569 B.n278 B.n191 71.676
R570 B.n285 B.n284 71.676
R571 B.n286 B.n189 71.676
R572 B.n293 B.n292 71.676
R573 B.n294 B.n187 71.676
R574 B.n301 B.n300 71.676
R575 B.n304 B.n303 71.676
R576 B.n196 B.n195 59.5399
R577 B.n249 B.n204 59.5399
R578 B.n98 B.n61 59.5399
R579 B.n119 B.n59 59.5399
R580 B.t11 B.n171 47.0532
R581 B.t7 B.n22 47.0532
R582 B.n354 B.t1 44.7579
R583 B.n413 B.t5 44.7579
R584 B.n333 B.t4 42.4627
R585 B.n18 B.t2 42.4627
R586 B.n348 B.t0 40.1674
R587 B.n407 B.t3 40.1674
R588 B.n163 B.t0 37.8722
R589 B.t3 B.n406 37.8722
R590 B.n340 B.t4 35.5769
R591 B.n405 B.t2 35.5769
R592 B.n347 B.t1 33.2817
R593 B.n11 B.t5 33.2817
R594 B.n321 B.t11 30.9864
R595 B.n391 B.t7 30.9864
R596 B.n379 B.n378 28.8785
R597 B.n385 B.n31 28.8785
R598 B.n307 B.n306 28.8785
R599 B.n311 B.n181 28.8785
R600 B B.n417 18.0485
R601 B.n195 B.n194 12.8005
R602 B.n204 B.n203 12.8005
R603 B.n61 B.n60 12.8005
R604 B.n59 B.n58 12.8005
R605 B.n62 B.n31 10.6151
R606 B.n65 B.n62 10.6151
R607 B.n66 B.n65 10.6151
R608 B.n69 B.n66 10.6151
R609 B.n70 B.n69 10.6151
R610 B.n73 B.n70 10.6151
R611 B.n74 B.n73 10.6151
R612 B.n77 B.n74 10.6151
R613 B.n78 B.n77 10.6151
R614 B.n81 B.n78 10.6151
R615 B.n82 B.n81 10.6151
R616 B.n85 B.n82 10.6151
R617 B.n86 B.n85 10.6151
R618 B.n89 B.n86 10.6151
R619 B.n90 B.n89 10.6151
R620 B.n93 B.n90 10.6151
R621 B.n94 B.n93 10.6151
R622 B.n97 B.n94 10.6151
R623 B.n102 B.n99 10.6151
R624 B.n103 B.n102 10.6151
R625 B.n106 B.n103 10.6151
R626 B.n107 B.n106 10.6151
R627 B.n110 B.n107 10.6151
R628 B.n111 B.n110 10.6151
R629 B.n114 B.n111 10.6151
R630 B.n115 B.n114 10.6151
R631 B.n118 B.n115 10.6151
R632 B.n123 B.n120 10.6151
R633 B.n124 B.n123 10.6151
R634 B.n127 B.n124 10.6151
R635 B.n128 B.n127 10.6151
R636 B.n131 B.n128 10.6151
R637 B.n132 B.n131 10.6151
R638 B.n135 B.n132 10.6151
R639 B.n136 B.n135 10.6151
R640 B.n139 B.n136 10.6151
R641 B.n140 B.n139 10.6151
R642 B.n143 B.n140 10.6151
R643 B.n144 B.n143 10.6151
R644 B.n147 B.n144 10.6151
R645 B.n148 B.n147 10.6151
R646 B.n151 B.n148 10.6151
R647 B.n153 B.n151 10.6151
R648 B.n154 B.n153 10.6151
R649 B.n379 B.n154 10.6151
R650 B.n307 B.n177 10.6151
R651 B.n317 B.n177 10.6151
R652 B.n318 B.n317 10.6151
R653 B.n319 B.n318 10.6151
R654 B.n319 B.n169 10.6151
R655 B.n329 B.n169 10.6151
R656 B.n330 B.n329 10.6151
R657 B.n331 B.n330 10.6151
R658 B.n331 B.n161 10.6151
R659 B.n342 B.n161 10.6151
R660 B.n343 B.n342 10.6151
R661 B.n345 B.n343 10.6151
R662 B.n345 B.n344 10.6151
R663 B.n344 B.n155 10.6151
R664 B.n357 B.n155 10.6151
R665 B.n358 B.n357 10.6151
R666 B.n359 B.n358 10.6151
R667 B.n360 B.n359 10.6151
R668 B.n362 B.n360 10.6151
R669 B.n363 B.n362 10.6151
R670 B.n364 B.n363 10.6151
R671 B.n365 B.n364 10.6151
R672 B.n367 B.n365 10.6151
R673 B.n368 B.n367 10.6151
R674 B.n369 B.n368 10.6151
R675 B.n370 B.n369 10.6151
R676 B.n372 B.n370 10.6151
R677 B.n373 B.n372 10.6151
R678 B.n374 B.n373 10.6151
R679 B.n375 B.n374 10.6151
R680 B.n377 B.n375 10.6151
R681 B.n378 B.n377 10.6151
R682 B.n215 B.n181 10.6151
R683 B.n216 B.n215 10.6151
R684 B.n217 B.n216 10.6151
R685 B.n217 B.n211 10.6151
R686 B.n223 B.n211 10.6151
R687 B.n224 B.n223 10.6151
R688 B.n225 B.n224 10.6151
R689 B.n225 B.n209 10.6151
R690 B.n231 B.n209 10.6151
R691 B.n232 B.n231 10.6151
R692 B.n233 B.n232 10.6151
R693 B.n233 B.n207 10.6151
R694 B.n239 B.n207 10.6151
R695 B.n240 B.n239 10.6151
R696 B.n241 B.n240 10.6151
R697 B.n241 B.n205 10.6151
R698 B.n247 B.n205 10.6151
R699 B.n248 B.n247 10.6151
R700 B.n250 B.n201 10.6151
R701 B.n256 B.n201 10.6151
R702 B.n257 B.n256 10.6151
R703 B.n258 B.n257 10.6151
R704 B.n258 B.n199 10.6151
R705 B.n264 B.n199 10.6151
R706 B.n265 B.n264 10.6151
R707 B.n266 B.n265 10.6151
R708 B.n266 B.n197 10.6151
R709 B.n273 B.n272 10.6151
R710 B.n274 B.n273 10.6151
R711 B.n274 B.n192 10.6151
R712 B.n280 B.n192 10.6151
R713 B.n281 B.n280 10.6151
R714 B.n282 B.n281 10.6151
R715 B.n282 B.n190 10.6151
R716 B.n288 B.n190 10.6151
R717 B.n289 B.n288 10.6151
R718 B.n290 B.n289 10.6151
R719 B.n290 B.n188 10.6151
R720 B.n296 B.n188 10.6151
R721 B.n297 B.n296 10.6151
R722 B.n298 B.n297 10.6151
R723 B.n298 B.n186 10.6151
R724 B.n186 B.n185 10.6151
R725 B.n305 B.n185 10.6151
R726 B.n306 B.n305 10.6151
R727 B.n312 B.n311 10.6151
R728 B.n313 B.n312 10.6151
R729 B.n313 B.n173 10.6151
R730 B.n323 B.n173 10.6151
R731 B.n324 B.n323 10.6151
R732 B.n325 B.n324 10.6151
R733 B.n325 B.n165 10.6151
R734 B.n336 B.n165 10.6151
R735 B.n337 B.n336 10.6151
R736 B.n338 B.n337 10.6151
R737 B.n338 B.n158 10.6151
R738 B.n350 B.n158 10.6151
R739 B.n351 B.n350 10.6151
R740 B.n352 B.n351 10.6151
R741 B.n352 B.n0 10.6151
R742 B.n411 B.n1 10.6151
R743 B.n411 B.n410 10.6151
R744 B.n410 B.n409 10.6151
R745 B.n409 B.n9 10.6151
R746 B.n403 B.n9 10.6151
R747 B.n403 B.n402 10.6151
R748 B.n402 B.n401 10.6151
R749 B.n401 B.n16 10.6151
R750 B.n395 B.n16 10.6151
R751 B.n395 B.n394 10.6151
R752 B.n394 B.n393 10.6151
R753 B.n393 B.n24 10.6151
R754 B.n387 B.n24 10.6151
R755 B.n387 B.n386 10.6151
R756 B.n386 B.n385 10.6151
R757 B.n98 B.n97 9.36635
R758 B.n120 B.n119 9.36635
R759 B.n249 B.n248 9.36635
R760 B.n272 B.n196 9.36635
R761 B.n417 B.n0 2.81026
R762 B.n417 B.n1 2.81026
R763 B.n99 B.n98 1.24928
R764 B.n119 B.n118 1.24928
R765 B.n250 B.n249 1.24928
R766 B.n197 B.n196 1.24928
R767 VN.n2 VN.t0 906.398
R768 VN.n0 VN.t4 906.398
R769 VN.n6 VN.t1 906.398
R770 VN.n4 VN.t2 906.398
R771 VN.n1 VN.t3 846.514
R772 VN.n5 VN.t5 846.514
R773 VN.n7 VN.n4 161.489
R774 VN.n3 VN.n0 161.489
R775 VN.n3 VN.n2 161.3
R776 VN.n7 VN.n6 161.3
R777 VN.n1 VN.n0 36.5157
R778 VN.n2 VN.n1 36.5157
R779 VN.n6 VN.n5 36.5157
R780 VN.n5 VN.n4 36.5157
R781 VN VN.n7 34.5024
R782 VN VN.n3 0.0516364
R783 VDD2.n1 VDD2.t1 81.3835
R784 VDD2.n2 VDD2.t4 81.0123
R785 VDD2.n1 VDD2.n0 74.1384
R786 VDD2 VDD2.n3 74.1357
R787 VDD2.n2 VDD2.n1 29.2799
R788 VDD2.n3 VDD2.t0 6.96106
R789 VDD2.n3 VDD2.t3 6.96106
R790 VDD2.n0 VDD2.t2 6.96106
R791 VDD2.n0 VDD2.t5 6.96106
R792 VDD2 VDD2.n2 0.485414
C0 VN VDD1 0.151379f
C1 VDD1 VTAIL 6.08304f
C2 VN VDD2 0.868904f
C3 VN VP 3.28524f
C4 VTAIL VDD2 6.11832f
C5 VP VTAIL 0.743532f
C6 VDD1 VDD2 0.577295f
C7 VP VDD1 0.984519f
C8 VN VTAIL 0.729196f
C9 VP VDD2 0.269097f
C10 VDD2 B 2.759663f
C11 VDD1 B 2.960594f
C12 VTAIL B 3.217461f
C13 VN B 5.08612f
C14 VP B 3.816312f
C15 VDD2.t1 B 0.780934f
C16 VDD2.t2 B 0.108996f
C17 VDD2.t5 B 0.108996f
C18 VDD2.n0 B 0.646846f
C19 VDD2.n1 B 1.23559f
C20 VDD2.t4 B 0.779732f
C21 VDD2.n2 B 1.31688f
C22 VDD2.t0 B 0.108996f
C23 VDD2.t3 B 0.108996f
C24 VDD2.n3 B 0.64683f
C25 VN.t4 B 0.082387f
C26 VN.n0 B 0.061846f
C27 VN.t3 B 0.079235f
C28 VN.n1 B 0.045976f
C29 VN.t0 B 0.082387f
C30 VN.n2 B 0.061785f
C31 VN.n3 B 0.082858f
C32 VN.t2 B 0.082387f
C33 VN.n4 B 0.061846f
C34 VN.t1 B 0.082387f
C35 VN.t5 B 0.079235f
C36 VN.n5 B 0.045976f
C37 VN.n6 B 0.061785f
C38 VN.n7 B 1.21382f
C39 VDD1.t4 B 0.771474f
C40 VDD1.t3 B 0.771073f
C41 VDD1.t2 B 0.10762f
C42 VDD1.t5 B 0.10762f
C43 VDD1.n0 B 0.638678f
C44 VDD1.n1 B 1.27532f
C45 VDD1.t1 B 0.10762f
C46 VDD1.t0 B 0.10762f
C47 VDD1.n2 B 0.638418f
C48 VDD1.n3 B 1.27099f
C49 VTAIL.t9 B 0.122756f
C50 VTAIL.t10 B 0.122756f
C51 VTAIL.n0 B 0.675243f
C52 VTAIL.n1 B 0.280513f
C53 VTAIL.t2 B 0.812519f
C54 VTAIL.n2 B 0.392445f
C55 VTAIL.t5 B 0.122756f
C56 VTAIL.t6 B 0.122756f
C57 VTAIL.n3 B 0.675243f
C58 VTAIL.n4 B 0.946087f
C59 VTAIL.t8 B 0.122756f
C60 VTAIL.t0 B 0.122756f
C61 VTAIL.n5 B 0.675246f
C62 VTAIL.n6 B 0.946084f
C63 VTAIL.t1 B 0.812522f
C64 VTAIL.n7 B 0.392442f
C65 VTAIL.t4 B 0.122756f
C66 VTAIL.t7 B 0.122756f
C67 VTAIL.n8 B 0.675246f
C68 VTAIL.n9 B 0.308758f
C69 VTAIL.t3 B 0.812519f
C70 VTAIL.n10 B 0.98616f
C71 VTAIL.t11 B 0.812519f
C72 VTAIL.n11 B 0.970797f
C73 VP.t1 B 0.083817f
C74 VP.n0 B 0.062919f
C75 VP.t4 B 0.08061f
C76 VP.n1 B 0.046774f
C77 VP.t5 B 0.083817f
C78 VP.n2 B 0.062857f
C79 VP.n3 B 1.20775f
C80 VP.n4 B 1.19794f
C81 VP.t3 B 0.08061f
C82 VP.t2 B 0.083817f
C83 VP.n5 B 0.062857f
C84 VP.n6 B 0.046774f
C85 VP.t0 B 0.083817f
C86 VP.n7 B 0.062857f
C87 VP.n8 B 0.031568f
.ends

