* NGSPICE file created from diff_pair_sample_1241.ext - technology: sky130A

.subckt diff_pair_sample_1241 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X1 VTAIL.t2 VN.t0 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X2 VTAIL.t1 VN.t1 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X3 VDD1.t0 VP.t1 VTAIL.t14 B.t9 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=0.56
X4 VTAIL.t3 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=0.56
X6 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=0.56
X7 VDD1.t3 VP.t2 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=0.56
X8 VDD1.t2 VP.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=0.56
X9 VTAIL.t5 VN.t3 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X10 VDD2.t5 VN.t4 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=0.56
X11 VDD1.t7 VP.t4 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X12 VDD2.t4 VN.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X13 VDD2.t3 VN.t6 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X14 VDD1.t6 VP.t5 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=0.56
X15 VDD2.t2 VN.t7 VTAIL.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=0.56
X16 VDD2.t1 VN.t8 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=3.14325 ps=19.38 w=19.05 l=0.56
X17 VTAIL.t9 VP.t6 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X18 VTAIL.t8 VP.t7 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X19 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=0.56
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.4295 pd=38.88 as=0 ps=0 w=19.05 l=0.56
X21 VDD1.t9 VP.t8 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X22 VTAIL.t6 VP.t9 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=3.14325 ps=19.38 w=19.05 l=0.56
X23 VDD2.t0 VN.t9 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=3.14325 pd=19.38 as=7.4295 ps=38.88 w=19.05 l=0.56
R0 VP.n6 VP.t3 914.61
R1 VP.n14 VP.t5 890.409
R2 VP.n16 VP.t6 890.409
R3 VP.n1 VP.t8 890.409
R4 VP.n20 VP.t0 890.409
R5 VP.n22 VP.t1 890.409
R6 VP.n11 VP.t2 890.409
R7 VP.n9 VP.t7 890.409
R8 VP.n8 VP.t4 890.409
R9 VP.n7 VP.t9 890.409
R10 VP.n23 VP.n22 161.3
R11 VP.n9 VP.n4 161.3
R12 VP.n10 VP.n3 161.3
R13 VP.n12 VP.n11 161.3
R14 VP.n21 VP.n0 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n15 VP.n2 161.3
R18 VP.n14 VP.n13 161.3
R19 VP.n8 VP.n5 80.6037
R20 VP.n18 VP.n1 80.6037
R21 VP.n16 VP.n1 48.2005
R22 VP.n20 VP.n1 48.2005
R23 VP.n9 VP.n8 48.2005
R24 VP.n8 VP.n7 48.2005
R25 VP.n13 VP.n12 47.3073
R26 VP.n6 VP.n5 45.0238
R27 VP.n15 VP.n14 36.5157
R28 VP.n22 VP.n21 36.5157
R29 VP.n11 VP.n10 36.5157
R30 VP.n7 VP.n6 17.2829
R31 VP.n16 VP.n15 11.6853
R32 VP.n21 VP.n20 11.6853
R33 VP.n10 VP.n9 11.6853
R34 VP.n5 VP.n4 0.285035
R35 VP.n18 VP.n17 0.285035
R36 VP.n19 VP.n18 0.285035
R37 VP.n4 VP.n3 0.189894
R38 VP.n12 VP.n3 0.189894
R39 VP.n13 VP.n2 0.189894
R40 VP.n17 VP.n2 0.189894
R41 VP.n19 VP.n0 0.189894
R42 VP.n23 VP.n0 0.189894
R43 VP VP.n23 0.0516364
R44 VDD1.n1 VDD1.t2 63.7516
R45 VDD1.n3 VDD1.t6 63.7515
R46 VDD1.n5 VDD1.n4 62.4639
R47 VDD1.n1 VDD1.n0 61.945
R48 VDD1.n7 VDD1.n6 61.9448
R49 VDD1.n3 VDD1.n2 61.9438
R50 VDD1.n7 VDD1.n5 44.7487
R51 VDD1.n6 VDD1.t4 1.03987
R52 VDD1.n6 VDD1.t3 1.03987
R53 VDD1.n0 VDD1.t8 1.03987
R54 VDD1.n0 VDD1.t7 1.03987
R55 VDD1.n4 VDD1.t1 1.03987
R56 VDD1.n4 VDD1.t0 1.03987
R57 VDD1.n2 VDD1.t5 1.03987
R58 VDD1.n2 VDD1.t9 1.03987
R59 VDD1 VDD1.n7 0.517741
R60 VDD1 VDD1.n1 0.2505
R61 VDD1.n5 VDD1.n3 0.136964
R62 VTAIL.n11 VTAIL.t16 46.3055
R63 VTAIL.n17 VTAIL.t19 46.3054
R64 VTAIL.n2 VTAIL.t14 46.3054
R65 VTAIL.n16 VTAIL.t13 46.3054
R66 VTAIL.n15 VTAIL.n14 45.2662
R67 VTAIL.n13 VTAIL.n12 45.2662
R68 VTAIL.n10 VTAIL.n9 45.2662
R69 VTAIL.n8 VTAIL.n7 45.2662
R70 VTAIL.n19 VTAIL.n18 45.265
R71 VTAIL.n1 VTAIL.n0 45.265
R72 VTAIL.n4 VTAIL.n3 45.265
R73 VTAIL.n6 VTAIL.n5 45.265
R74 VTAIL.n8 VTAIL.n6 30.3238
R75 VTAIL.n17 VTAIL.n16 29.5565
R76 VTAIL.n18 VTAIL.t18 1.03987
R77 VTAIL.n18 VTAIL.t1 1.03987
R78 VTAIL.n0 VTAIL.t17 1.03987
R79 VTAIL.n0 VTAIL.t5 1.03987
R80 VTAIL.n3 VTAIL.t7 1.03987
R81 VTAIL.n3 VTAIL.t15 1.03987
R82 VTAIL.n5 VTAIL.t10 1.03987
R83 VTAIL.n5 VTAIL.t9 1.03987
R84 VTAIL.n14 VTAIL.t11 1.03987
R85 VTAIL.n14 VTAIL.t8 1.03987
R86 VTAIL.n12 VTAIL.t12 1.03987
R87 VTAIL.n12 VTAIL.t6 1.03987
R88 VTAIL.n9 VTAIL.t4 1.03987
R89 VTAIL.n9 VTAIL.t3 1.03987
R90 VTAIL.n7 VTAIL.t0 1.03987
R91 VTAIL.n7 VTAIL.t2 1.03987
R92 VTAIL.n13 VTAIL.n11 0.853948
R93 VTAIL.n2 VTAIL.n1 0.853948
R94 VTAIL.n10 VTAIL.n8 0.767741
R95 VTAIL.n11 VTAIL.n10 0.767741
R96 VTAIL.n15 VTAIL.n13 0.767741
R97 VTAIL.n16 VTAIL.n15 0.767741
R98 VTAIL.n6 VTAIL.n4 0.767741
R99 VTAIL.n4 VTAIL.n2 0.767741
R100 VTAIL.n19 VTAIL.n17 0.767741
R101 VTAIL VTAIL.n1 0.634121
R102 VTAIL VTAIL.n19 0.134121
R103 B.n461 B.t21 1024.95
R104 B.n618 B.t14 1024.95
R105 B.n118 B.t18 1024.95
R106 B.n115 B.t10 1024.95
R107 B.n874 B.n873 585
R108 B.n383 B.n114 585
R109 B.n382 B.n381 585
R110 B.n380 B.n379 585
R111 B.n378 B.n377 585
R112 B.n376 B.n375 585
R113 B.n374 B.n373 585
R114 B.n372 B.n371 585
R115 B.n370 B.n369 585
R116 B.n368 B.n367 585
R117 B.n366 B.n365 585
R118 B.n364 B.n363 585
R119 B.n362 B.n361 585
R120 B.n360 B.n359 585
R121 B.n358 B.n357 585
R122 B.n356 B.n355 585
R123 B.n354 B.n353 585
R124 B.n352 B.n351 585
R125 B.n350 B.n349 585
R126 B.n348 B.n347 585
R127 B.n346 B.n345 585
R128 B.n344 B.n343 585
R129 B.n342 B.n341 585
R130 B.n340 B.n339 585
R131 B.n338 B.n337 585
R132 B.n336 B.n335 585
R133 B.n334 B.n333 585
R134 B.n332 B.n331 585
R135 B.n330 B.n329 585
R136 B.n328 B.n327 585
R137 B.n326 B.n325 585
R138 B.n324 B.n323 585
R139 B.n322 B.n321 585
R140 B.n320 B.n319 585
R141 B.n318 B.n317 585
R142 B.n316 B.n315 585
R143 B.n314 B.n313 585
R144 B.n312 B.n311 585
R145 B.n310 B.n309 585
R146 B.n308 B.n307 585
R147 B.n306 B.n305 585
R148 B.n304 B.n303 585
R149 B.n302 B.n301 585
R150 B.n300 B.n299 585
R151 B.n298 B.n297 585
R152 B.n296 B.n295 585
R153 B.n294 B.n293 585
R154 B.n292 B.n291 585
R155 B.n290 B.n289 585
R156 B.n288 B.n287 585
R157 B.n286 B.n285 585
R158 B.n284 B.n283 585
R159 B.n282 B.n281 585
R160 B.n280 B.n279 585
R161 B.n278 B.n277 585
R162 B.n276 B.n275 585
R163 B.n274 B.n273 585
R164 B.n272 B.n271 585
R165 B.n270 B.n269 585
R166 B.n268 B.n267 585
R167 B.n266 B.n265 585
R168 B.n264 B.n263 585
R169 B.n262 B.n261 585
R170 B.n260 B.n259 585
R171 B.n258 B.n257 585
R172 B.n256 B.n255 585
R173 B.n254 B.n253 585
R174 B.n252 B.n251 585
R175 B.n250 B.n249 585
R176 B.n248 B.n247 585
R177 B.n246 B.n245 585
R178 B.n244 B.n243 585
R179 B.n242 B.n241 585
R180 B.n240 B.n239 585
R181 B.n238 B.n237 585
R182 B.n236 B.n235 585
R183 B.n234 B.n233 585
R184 B.n232 B.n231 585
R185 B.n230 B.n229 585
R186 B.n228 B.n227 585
R187 B.n226 B.n225 585
R188 B.n224 B.n223 585
R189 B.n222 B.n221 585
R190 B.n220 B.n219 585
R191 B.n218 B.n217 585
R192 B.n216 B.n215 585
R193 B.n214 B.n213 585
R194 B.n212 B.n211 585
R195 B.n210 B.n209 585
R196 B.n208 B.n207 585
R197 B.n206 B.n205 585
R198 B.n204 B.n203 585
R199 B.n202 B.n201 585
R200 B.n200 B.n199 585
R201 B.n198 B.n197 585
R202 B.n196 B.n195 585
R203 B.n194 B.n193 585
R204 B.n192 B.n191 585
R205 B.n190 B.n189 585
R206 B.n188 B.n187 585
R207 B.n186 B.n185 585
R208 B.n184 B.n183 585
R209 B.n182 B.n181 585
R210 B.n180 B.n179 585
R211 B.n178 B.n177 585
R212 B.n176 B.n175 585
R213 B.n174 B.n173 585
R214 B.n172 B.n171 585
R215 B.n170 B.n169 585
R216 B.n168 B.n167 585
R217 B.n166 B.n165 585
R218 B.n164 B.n163 585
R219 B.n162 B.n161 585
R220 B.n160 B.n159 585
R221 B.n158 B.n157 585
R222 B.n156 B.n155 585
R223 B.n154 B.n153 585
R224 B.n152 B.n151 585
R225 B.n150 B.n149 585
R226 B.n148 B.n147 585
R227 B.n146 B.n145 585
R228 B.n144 B.n143 585
R229 B.n142 B.n141 585
R230 B.n140 B.n139 585
R231 B.n138 B.n137 585
R232 B.n136 B.n135 585
R233 B.n134 B.n133 585
R234 B.n132 B.n131 585
R235 B.n130 B.n129 585
R236 B.n128 B.n127 585
R237 B.n126 B.n125 585
R238 B.n124 B.n123 585
R239 B.n122 B.n121 585
R240 B.n46 B.n45 585
R241 B.n872 B.n47 585
R242 B.n877 B.n47 585
R243 B.n871 B.n870 585
R244 B.n870 B.n43 585
R245 B.n869 B.n42 585
R246 B.n883 B.n42 585
R247 B.n868 B.n41 585
R248 B.n884 B.n41 585
R249 B.n867 B.n40 585
R250 B.n885 B.n40 585
R251 B.n866 B.n865 585
R252 B.n865 B.n36 585
R253 B.n864 B.n35 585
R254 B.n891 B.n35 585
R255 B.n863 B.n34 585
R256 B.n892 B.n34 585
R257 B.n862 B.n33 585
R258 B.n893 B.n33 585
R259 B.n861 B.n860 585
R260 B.n860 B.n29 585
R261 B.n859 B.n28 585
R262 B.n899 B.n28 585
R263 B.n858 B.n27 585
R264 B.n900 B.n27 585
R265 B.n857 B.n26 585
R266 B.n901 B.n26 585
R267 B.n856 B.n855 585
R268 B.n855 B.n25 585
R269 B.n854 B.n21 585
R270 B.n907 B.n21 585
R271 B.n853 B.n20 585
R272 B.n908 B.n20 585
R273 B.n852 B.n19 585
R274 B.n909 B.n19 585
R275 B.n851 B.n850 585
R276 B.n850 B.n15 585
R277 B.n849 B.n14 585
R278 B.n915 B.n14 585
R279 B.n848 B.n13 585
R280 B.n916 B.n13 585
R281 B.n847 B.n12 585
R282 B.n917 B.n12 585
R283 B.n846 B.n845 585
R284 B.n845 B.n11 585
R285 B.n844 B.n7 585
R286 B.n923 B.n7 585
R287 B.n843 B.n6 585
R288 B.n924 B.n6 585
R289 B.n842 B.n5 585
R290 B.n925 B.n5 585
R291 B.n841 B.n840 585
R292 B.n840 B.n4 585
R293 B.n839 B.n384 585
R294 B.n839 B.n838 585
R295 B.n828 B.n385 585
R296 B.n831 B.n385 585
R297 B.n830 B.n829 585
R298 B.n832 B.n830 585
R299 B.n827 B.n390 585
R300 B.n390 B.n389 585
R301 B.n826 B.n825 585
R302 B.n825 B.n824 585
R303 B.n392 B.n391 585
R304 B.n393 B.n392 585
R305 B.n817 B.n816 585
R306 B.n818 B.n817 585
R307 B.n815 B.n397 585
R308 B.n400 B.n397 585
R309 B.n814 B.n813 585
R310 B.n813 B.n812 585
R311 B.n399 B.n398 585
R312 B.n805 B.n399 585
R313 B.n804 B.n803 585
R314 B.n806 B.n804 585
R315 B.n802 B.n405 585
R316 B.n405 B.n404 585
R317 B.n801 B.n800 585
R318 B.n800 B.n799 585
R319 B.n407 B.n406 585
R320 B.n408 B.n407 585
R321 B.n792 B.n791 585
R322 B.n793 B.n792 585
R323 B.n790 B.n413 585
R324 B.n413 B.n412 585
R325 B.n789 B.n788 585
R326 B.n788 B.n787 585
R327 B.n415 B.n414 585
R328 B.n416 B.n415 585
R329 B.n780 B.n779 585
R330 B.n781 B.n780 585
R331 B.n778 B.n421 585
R332 B.n421 B.n420 585
R333 B.n777 B.n776 585
R334 B.n776 B.n775 585
R335 B.n423 B.n422 585
R336 B.n424 B.n423 585
R337 B.n768 B.n767 585
R338 B.n769 B.n768 585
R339 B.n427 B.n426 585
R340 B.n500 B.n498 585
R341 B.n501 B.n497 585
R342 B.n501 B.n428 585
R343 B.n504 B.n503 585
R344 B.n505 B.n496 585
R345 B.n507 B.n506 585
R346 B.n509 B.n495 585
R347 B.n512 B.n511 585
R348 B.n513 B.n494 585
R349 B.n515 B.n514 585
R350 B.n517 B.n493 585
R351 B.n520 B.n519 585
R352 B.n521 B.n492 585
R353 B.n523 B.n522 585
R354 B.n525 B.n491 585
R355 B.n528 B.n527 585
R356 B.n529 B.n490 585
R357 B.n531 B.n530 585
R358 B.n533 B.n489 585
R359 B.n536 B.n535 585
R360 B.n537 B.n488 585
R361 B.n539 B.n538 585
R362 B.n541 B.n487 585
R363 B.n544 B.n543 585
R364 B.n545 B.n486 585
R365 B.n547 B.n546 585
R366 B.n549 B.n485 585
R367 B.n552 B.n551 585
R368 B.n553 B.n484 585
R369 B.n555 B.n554 585
R370 B.n557 B.n483 585
R371 B.n560 B.n559 585
R372 B.n561 B.n482 585
R373 B.n563 B.n562 585
R374 B.n565 B.n481 585
R375 B.n568 B.n567 585
R376 B.n569 B.n480 585
R377 B.n571 B.n570 585
R378 B.n573 B.n479 585
R379 B.n576 B.n575 585
R380 B.n577 B.n478 585
R381 B.n579 B.n578 585
R382 B.n581 B.n477 585
R383 B.n584 B.n583 585
R384 B.n585 B.n476 585
R385 B.n587 B.n586 585
R386 B.n589 B.n475 585
R387 B.n592 B.n591 585
R388 B.n593 B.n474 585
R389 B.n595 B.n594 585
R390 B.n597 B.n473 585
R391 B.n600 B.n599 585
R392 B.n601 B.n472 585
R393 B.n603 B.n602 585
R394 B.n605 B.n471 585
R395 B.n608 B.n607 585
R396 B.n609 B.n470 585
R397 B.n611 B.n610 585
R398 B.n613 B.n469 585
R399 B.n616 B.n615 585
R400 B.n617 B.n468 585
R401 B.n622 B.n621 585
R402 B.n624 B.n467 585
R403 B.n627 B.n626 585
R404 B.n628 B.n466 585
R405 B.n630 B.n629 585
R406 B.n632 B.n465 585
R407 B.n635 B.n634 585
R408 B.n636 B.n464 585
R409 B.n638 B.n637 585
R410 B.n640 B.n463 585
R411 B.n643 B.n642 585
R412 B.n645 B.n460 585
R413 B.n647 B.n646 585
R414 B.n649 B.n459 585
R415 B.n652 B.n651 585
R416 B.n653 B.n458 585
R417 B.n655 B.n654 585
R418 B.n657 B.n457 585
R419 B.n660 B.n659 585
R420 B.n661 B.n456 585
R421 B.n663 B.n662 585
R422 B.n665 B.n455 585
R423 B.n668 B.n667 585
R424 B.n669 B.n454 585
R425 B.n671 B.n670 585
R426 B.n673 B.n453 585
R427 B.n676 B.n675 585
R428 B.n677 B.n452 585
R429 B.n679 B.n678 585
R430 B.n681 B.n451 585
R431 B.n684 B.n683 585
R432 B.n685 B.n450 585
R433 B.n687 B.n686 585
R434 B.n689 B.n449 585
R435 B.n692 B.n691 585
R436 B.n693 B.n448 585
R437 B.n695 B.n694 585
R438 B.n697 B.n447 585
R439 B.n700 B.n699 585
R440 B.n701 B.n446 585
R441 B.n703 B.n702 585
R442 B.n705 B.n445 585
R443 B.n708 B.n707 585
R444 B.n709 B.n444 585
R445 B.n711 B.n710 585
R446 B.n713 B.n443 585
R447 B.n716 B.n715 585
R448 B.n717 B.n442 585
R449 B.n719 B.n718 585
R450 B.n721 B.n441 585
R451 B.n724 B.n723 585
R452 B.n725 B.n440 585
R453 B.n727 B.n726 585
R454 B.n729 B.n439 585
R455 B.n732 B.n731 585
R456 B.n733 B.n438 585
R457 B.n735 B.n734 585
R458 B.n737 B.n437 585
R459 B.n740 B.n739 585
R460 B.n741 B.n436 585
R461 B.n743 B.n742 585
R462 B.n745 B.n435 585
R463 B.n748 B.n747 585
R464 B.n749 B.n434 585
R465 B.n751 B.n750 585
R466 B.n753 B.n433 585
R467 B.n756 B.n755 585
R468 B.n757 B.n432 585
R469 B.n759 B.n758 585
R470 B.n761 B.n431 585
R471 B.n762 B.n430 585
R472 B.n765 B.n764 585
R473 B.n766 B.n429 585
R474 B.n429 B.n428 585
R475 B.n771 B.n770 585
R476 B.n770 B.n769 585
R477 B.n772 B.n425 585
R478 B.n425 B.n424 585
R479 B.n774 B.n773 585
R480 B.n775 B.n774 585
R481 B.n419 B.n418 585
R482 B.n420 B.n419 585
R483 B.n783 B.n782 585
R484 B.n782 B.n781 585
R485 B.n784 B.n417 585
R486 B.n417 B.n416 585
R487 B.n786 B.n785 585
R488 B.n787 B.n786 585
R489 B.n411 B.n410 585
R490 B.n412 B.n411 585
R491 B.n795 B.n794 585
R492 B.n794 B.n793 585
R493 B.n796 B.n409 585
R494 B.n409 B.n408 585
R495 B.n798 B.n797 585
R496 B.n799 B.n798 585
R497 B.n403 B.n402 585
R498 B.n404 B.n403 585
R499 B.n808 B.n807 585
R500 B.n807 B.n806 585
R501 B.n809 B.n401 585
R502 B.n805 B.n401 585
R503 B.n811 B.n810 585
R504 B.n812 B.n811 585
R505 B.n396 B.n395 585
R506 B.n400 B.n396 585
R507 B.n820 B.n819 585
R508 B.n819 B.n818 585
R509 B.n821 B.n394 585
R510 B.n394 B.n393 585
R511 B.n823 B.n822 585
R512 B.n824 B.n823 585
R513 B.n388 B.n387 585
R514 B.n389 B.n388 585
R515 B.n834 B.n833 585
R516 B.n833 B.n832 585
R517 B.n835 B.n386 585
R518 B.n831 B.n386 585
R519 B.n837 B.n836 585
R520 B.n838 B.n837 585
R521 B.n2 B.n0 585
R522 B.n4 B.n2 585
R523 B.n3 B.n1 585
R524 B.n924 B.n3 585
R525 B.n922 B.n921 585
R526 B.n923 B.n922 585
R527 B.n920 B.n8 585
R528 B.n11 B.n8 585
R529 B.n919 B.n918 585
R530 B.n918 B.n917 585
R531 B.n10 B.n9 585
R532 B.n916 B.n10 585
R533 B.n914 B.n913 585
R534 B.n915 B.n914 585
R535 B.n912 B.n16 585
R536 B.n16 B.n15 585
R537 B.n911 B.n910 585
R538 B.n910 B.n909 585
R539 B.n18 B.n17 585
R540 B.n908 B.n18 585
R541 B.n906 B.n905 585
R542 B.n907 B.n906 585
R543 B.n904 B.n22 585
R544 B.n25 B.n22 585
R545 B.n903 B.n902 585
R546 B.n902 B.n901 585
R547 B.n24 B.n23 585
R548 B.n900 B.n24 585
R549 B.n898 B.n897 585
R550 B.n899 B.n898 585
R551 B.n896 B.n30 585
R552 B.n30 B.n29 585
R553 B.n895 B.n894 585
R554 B.n894 B.n893 585
R555 B.n32 B.n31 585
R556 B.n892 B.n32 585
R557 B.n890 B.n889 585
R558 B.n891 B.n890 585
R559 B.n888 B.n37 585
R560 B.n37 B.n36 585
R561 B.n887 B.n886 585
R562 B.n886 B.n885 585
R563 B.n39 B.n38 585
R564 B.n884 B.n39 585
R565 B.n882 B.n881 585
R566 B.n883 B.n882 585
R567 B.n880 B.n44 585
R568 B.n44 B.n43 585
R569 B.n879 B.n878 585
R570 B.n878 B.n877 585
R571 B.n927 B.n926 585
R572 B.n926 B.n925 585
R573 B.n770 B.n427 492.5
R574 B.n878 B.n46 492.5
R575 B.n768 B.n429 492.5
R576 B.n874 B.n47 492.5
R577 B.n876 B.n875 256.663
R578 B.n876 B.n113 256.663
R579 B.n876 B.n112 256.663
R580 B.n876 B.n111 256.663
R581 B.n876 B.n110 256.663
R582 B.n876 B.n109 256.663
R583 B.n876 B.n108 256.663
R584 B.n876 B.n107 256.663
R585 B.n876 B.n106 256.663
R586 B.n876 B.n105 256.663
R587 B.n876 B.n104 256.663
R588 B.n876 B.n103 256.663
R589 B.n876 B.n102 256.663
R590 B.n876 B.n101 256.663
R591 B.n876 B.n100 256.663
R592 B.n876 B.n99 256.663
R593 B.n876 B.n98 256.663
R594 B.n876 B.n97 256.663
R595 B.n876 B.n96 256.663
R596 B.n876 B.n95 256.663
R597 B.n876 B.n94 256.663
R598 B.n876 B.n93 256.663
R599 B.n876 B.n92 256.663
R600 B.n876 B.n91 256.663
R601 B.n876 B.n90 256.663
R602 B.n876 B.n89 256.663
R603 B.n876 B.n88 256.663
R604 B.n876 B.n87 256.663
R605 B.n876 B.n86 256.663
R606 B.n876 B.n85 256.663
R607 B.n876 B.n84 256.663
R608 B.n876 B.n83 256.663
R609 B.n876 B.n82 256.663
R610 B.n876 B.n81 256.663
R611 B.n876 B.n80 256.663
R612 B.n876 B.n79 256.663
R613 B.n876 B.n78 256.663
R614 B.n876 B.n77 256.663
R615 B.n876 B.n76 256.663
R616 B.n876 B.n75 256.663
R617 B.n876 B.n74 256.663
R618 B.n876 B.n73 256.663
R619 B.n876 B.n72 256.663
R620 B.n876 B.n71 256.663
R621 B.n876 B.n70 256.663
R622 B.n876 B.n69 256.663
R623 B.n876 B.n68 256.663
R624 B.n876 B.n67 256.663
R625 B.n876 B.n66 256.663
R626 B.n876 B.n65 256.663
R627 B.n876 B.n64 256.663
R628 B.n876 B.n63 256.663
R629 B.n876 B.n62 256.663
R630 B.n876 B.n61 256.663
R631 B.n876 B.n60 256.663
R632 B.n876 B.n59 256.663
R633 B.n876 B.n58 256.663
R634 B.n876 B.n57 256.663
R635 B.n876 B.n56 256.663
R636 B.n876 B.n55 256.663
R637 B.n876 B.n54 256.663
R638 B.n876 B.n53 256.663
R639 B.n876 B.n52 256.663
R640 B.n876 B.n51 256.663
R641 B.n876 B.n50 256.663
R642 B.n876 B.n49 256.663
R643 B.n876 B.n48 256.663
R644 B.n499 B.n428 256.663
R645 B.n502 B.n428 256.663
R646 B.n508 B.n428 256.663
R647 B.n510 B.n428 256.663
R648 B.n516 B.n428 256.663
R649 B.n518 B.n428 256.663
R650 B.n524 B.n428 256.663
R651 B.n526 B.n428 256.663
R652 B.n532 B.n428 256.663
R653 B.n534 B.n428 256.663
R654 B.n540 B.n428 256.663
R655 B.n542 B.n428 256.663
R656 B.n548 B.n428 256.663
R657 B.n550 B.n428 256.663
R658 B.n556 B.n428 256.663
R659 B.n558 B.n428 256.663
R660 B.n564 B.n428 256.663
R661 B.n566 B.n428 256.663
R662 B.n572 B.n428 256.663
R663 B.n574 B.n428 256.663
R664 B.n580 B.n428 256.663
R665 B.n582 B.n428 256.663
R666 B.n588 B.n428 256.663
R667 B.n590 B.n428 256.663
R668 B.n596 B.n428 256.663
R669 B.n598 B.n428 256.663
R670 B.n604 B.n428 256.663
R671 B.n606 B.n428 256.663
R672 B.n612 B.n428 256.663
R673 B.n614 B.n428 256.663
R674 B.n623 B.n428 256.663
R675 B.n625 B.n428 256.663
R676 B.n631 B.n428 256.663
R677 B.n633 B.n428 256.663
R678 B.n639 B.n428 256.663
R679 B.n641 B.n428 256.663
R680 B.n648 B.n428 256.663
R681 B.n650 B.n428 256.663
R682 B.n656 B.n428 256.663
R683 B.n658 B.n428 256.663
R684 B.n664 B.n428 256.663
R685 B.n666 B.n428 256.663
R686 B.n672 B.n428 256.663
R687 B.n674 B.n428 256.663
R688 B.n680 B.n428 256.663
R689 B.n682 B.n428 256.663
R690 B.n688 B.n428 256.663
R691 B.n690 B.n428 256.663
R692 B.n696 B.n428 256.663
R693 B.n698 B.n428 256.663
R694 B.n704 B.n428 256.663
R695 B.n706 B.n428 256.663
R696 B.n712 B.n428 256.663
R697 B.n714 B.n428 256.663
R698 B.n720 B.n428 256.663
R699 B.n722 B.n428 256.663
R700 B.n728 B.n428 256.663
R701 B.n730 B.n428 256.663
R702 B.n736 B.n428 256.663
R703 B.n738 B.n428 256.663
R704 B.n744 B.n428 256.663
R705 B.n746 B.n428 256.663
R706 B.n752 B.n428 256.663
R707 B.n754 B.n428 256.663
R708 B.n760 B.n428 256.663
R709 B.n763 B.n428 256.663
R710 B.n770 B.n425 163.367
R711 B.n774 B.n425 163.367
R712 B.n774 B.n419 163.367
R713 B.n782 B.n419 163.367
R714 B.n782 B.n417 163.367
R715 B.n786 B.n417 163.367
R716 B.n786 B.n411 163.367
R717 B.n794 B.n411 163.367
R718 B.n794 B.n409 163.367
R719 B.n798 B.n409 163.367
R720 B.n798 B.n403 163.367
R721 B.n807 B.n403 163.367
R722 B.n807 B.n401 163.367
R723 B.n811 B.n401 163.367
R724 B.n811 B.n396 163.367
R725 B.n819 B.n396 163.367
R726 B.n819 B.n394 163.367
R727 B.n823 B.n394 163.367
R728 B.n823 B.n388 163.367
R729 B.n833 B.n388 163.367
R730 B.n833 B.n386 163.367
R731 B.n837 B.n386 163.367
R732 B.n837 B.n2 163.367
R733 B.n926 B.n2 163.367
R734 B.n926 B.n3 163.367
R735 B.n922 B.n3 163.367
R736 B.n922 B.n8 163.367
R737 B.n918 B.n8 163.367
R738 B.n918 B.n10 163.367
R739 B.n914 B.n10 163.367
R740 B.n914 B.n16 163.367
R741 B.n910 B.n16 163.367
R742 B.n910 B.n18 163.367
R743 B.n906 B.n18 163.367
R744 B.n906 B.n22 163.367
R745 B.n902 B.n22 163.367
R746 B.n902 B.n24 163.367
R747 B.n898 B.n24 163.367
R748 B.n898 B.n30 163.367
R749 B.n894 B.n30 163.367
R750 B.n894 B.n32 163.367
R751 B.n890 B.n32 163.367
R752 B.n890 B.n37 163.367
R753 B.n886 B.n37 163.367
R754 B.n886 B.n39 163.367
R755 B.n882 B.n39 163.367
R756 B.n882 B.n44 163.367
R757 B.n878 B.n44 163.367
R758 B.n501 B.n500 163.367
R759 B.n503 B.n501 163.367
R760 B.n507 B.n496 163.367
R761 B.n511 B.n509 163.367
R762 B.n515 B.n494 163.367
R763 B.n519 B.n517 163.367
R764 B.n523 B.n492 163.367
R765 B.n527 B.n525 163.367
R766 B.n531 B.n490 163.367
R767 B.n535 B.n533 163.367
R768 B.n539 B.n488 163.367
R769 B.n543 B.n541 163.367
R770 B.n547 B.n486 163.367
R771 B.n551 B.n549 163.367
R772 B.n555 B.n484 163.367
R773 B.n559 B.n557 163.367
R774 B.n563 B.n482 163.367
R775 B.n567 B.n565 163.367
R776 B.n571 B.n480 163.367
R777 B.n575 B.n573 163.367
R778 B.n579 B.n478 163.367
R779 B.n583 B.n581 163.367
R780 B.n587 B.n476 163.367
R781 B.n591 B.n589 163.367
R782 B.n595 B.n474 163.367
R783 B.n599 B.n597 163.367
R784 B.n603 B.n472 163.367
R785 B.n607 B.n605 163.367
R786 B.n611 B.n470 163.367
R787 B.n615 B.n613 163.367
R788 B.n622 B.n468 163.367
R789 B.n626 B.n624 163.367
R790 B.n630 B.n466 163.367
R791 B.n634 B.n632 163.367
R792 B.n638 B.n464 163.367
R793 B.n642 B.n640 163.367
R794 B.n647 B.n460 163.367
R795 B.n651 B.n649 163.367
R796 B.n655 B.n458 163.367
R797 B.n659 B.n657 163.367
R798 B.n663 B.n456 163.367
R799 B.n667 B.n665 163.367
R800 B.n671 B.n454 163.367
R801 B.n675 B.n673 163.367
R802 B.n679 B.n452 163.367
R803 B.n683 B.n681 163.367
R804 B.n687 B.n450 163.367
R805 B.n691 B.n689 163.367
R806 B.n695 B.n448 163.367
R807 B.n699 B.n697 163.367
R808 B.n703 B.n446 163.367
R809 B.n707 B.n705 163.367
R810 B.n711 B.n444 163.367
R811 B.n715 B.n713 163.367
R812 B.n719 B.n442 163.367
R813 B.n723 B.n721 163.367
R814 B.n727 B.n440 163.367
R815 B.n731 B.n729 163.367
R816 B.n735 B.n438 163.367
R817 B.n739 B.n737 163.367
R818 B.n743 B.n436 163.367
R819 B.n747 B.n745 163.367
R820 B.n751 B.n434 163.367
R821 B.n755 B.n753 163.367
R822 B.n759 B.n432 163.367
R823 B.n762 B.n761 163.367
R824 B.n764 B.n429 163.367
R825 B.n768 B.n423 163.367
R826 B.n776 B.n423 163.367
R827 B.n776 B.n421 163.367
R828 B.n780 B.n421 163.367
R829 B.n780 B.n415 163.367
R830 B.n788 B.n415 163.367
R831 B.n788 B.n413 163.367
R832 B.n792 B.n413 163.367
R833 B.n792 B.n407 163.367
R834 B.n800 B.n407 163.367
R835 B.n800 B.n405 163.367
R836 B.n804 B.n405 163.367
R837 B.n804 B.n399 163.367
R838 B.n813 B.n399 163.367
R839 B.n813 B.n397 163.367
R840 B.n817 B.n397 163.367
R841 B.n817 B.n392 163.367
R842 B.n825 B.n392 163.367
R843 B.n825 B.n390 163.367
R844 B.n830 B.n390 163.367
R845 B.n830 B.n385 163.367
R846 B.n839 B.n385 163.367
R847 B.n840 B.n839 163.367
R848 B.n840 B.n5 163.367
R849 B.n6 B.n5 163.367
R850 B.n7 B.n6 163.367
R851 B.n845 B.n7 163.367
R852 B.n845 B.n12 163.367
R853 B.n13 B.n12 163.367
R854 B.n14 B.n13 163.367
R855 B.n850 B.n14 163.367
R856 B.n850 B.n19 163.367
R857 B.n20 B.n19 163.367
R858 B.n21 B.n20 163.367
R859 B.n855 B.n21 163.367
R860 B.n855 B.n26 163.367
R861 B.n27 B.n26 163.367
R862 B.n28 B.n27 163.367
R863 B.n860 B.n28 163.367
R864 B.n860 B.n33 163.367
R865 B.n34 B.n33 163.367
R866 B.n35 B.n34 163.367
R867 B.n865 B.n35 163.367
R868 B.n865 B.n40 163.367
R869 B.n41 B.n40 163.367
R870 B.n42 B.n41 163.367
R871 B.n870 B.n42 163.367
R872 B.n870 B.n47 163.367
R873 B.n123 B.n122 163.367
R874 B.n127 B.n126 163.367
R875 B.n131 B.n130 163.367
R876 B.n135 B.n134 163.367
R877 B.n139 B.n138 163.367
R878 B.n143 B.n142 163.367
R879 B.n147 B.n146 163.367
R880 B.n151 B.n150 163.367
R881 B.n155 B.n154 163.367
R882 B.n159 B.n158 163.367
R883 B.n163 B.n162 163.367
R884 B.n167 B.n166 163.367
R885 B.n171 B.n170 163.367
R886 B.n175 B.n174 163.367
R887 B.n179 B.n178 163.367
R888 B.n183 B.n182 163.367
R889 B.n187 B.n186 163.367
R890 B.n191 B.n190 163.367
R891 B.n195 B.n194 163.367
R892 B.n199 B.n198 163.367
R893 B.n203 B.n202 163.367
R894 B.n207 B.n206 163.367
R895 B.n211 B.n210 163.367
R896 B.n215 B.n214 163.367
R897 B.n219 B.n218 163.367
R898 B.n223 B.n222 163.367
R899 B.n227 B.n226 163.367
R900 B.n231 B.n230 163.367
R901 B.n235 B.n234 163.367
R902 B.n239 B.n238 163.367
R903 B.n243 B.n242 163.367
R904 B.n247 B.n246 163.367
R905 B.n251 B.n250 163.367
R906 B.n255 B.n254 163.367
R907 B.n259 B.n258 163.367
R908 B.n263 B.n262 163.367
R909 B.n267 B.n266 163.367
R910 B.n271 B.n270 163.367
R911 B.n275 B.n274 163.367
R912 B.n279 B.n278 163.367
R913 B.n283 B.n282 163.367
R914 B.n287 B.n286 163.367
R915 B.n291 B.n290 163.367
R916 B.n295 B.n294 163.367
R917 B.n299 B.n298 163.367
R918 B.n303 B.n302 163.367
R919 B.n307 B.n306 163.367
R920 B.n311 B.n310 163.367
R921 B.n315 B.n314 163.367
R922 B.n319 B.n318 163.367
R923 B.n323 B.n322 163.367
R924 B.n327 B.n326 163.367
R925 B.n331 B.n330 163.367
R926 B.n335 B.n334 163.367
R927 B.n339 B.n338 163.367
R928 B.n343 B.n342 163.367
R929 B.n347 B.n346 163.367
R930 B.n351 B.n350 163.367
R931 B.n355 B.n354 163.367
R932 B.n359 B.n358 163.367
R933 B.n363 B.n362 163.367
R934 B.n367 B.n366 163.367
R935 B.n371 B.n370 163.367
R936 B.n375 B.n374 163.367
R937 B.n379 B.n378 163.367
R938 B.n381 B.n114 163.367
R939 B.n461 B.t23 84.6443
R940 B.n115 B.t12 84.6443
R941 B.n618 B.t17 84.6186
R942 B.n118 B.t19 84.6186
R943 B.n499 B.n427 71.676
R944 B.n503 B.n502 71.676
R945 B.n508 B.n507 71.676
R946 B.n511 B.n510 71.676
R947 B.n516 B.n515 71.676
R948 B.n519 B.n518 71.676
R949 B.n524 B.n523 71.676
R950 B.n527 B.n526 71.676
R951 B.n532 B.n531 71.676
R952 B.n535 B.n534 71.676
R953 B.n540 B.n539 71.676
R954 B.n543 B.n542 71.676
R955 B.n548 B.n547 71.676
R956 B.n551 B.n550 71.676
R957 B.n556 B.n555 71.676
R958 B.n559 B.n558 71.676
R959 B.n564 B.n563 71.676
R960 B.n567 B.n566 71.676
R961 B.n572 B.n571 71.676
R962 B.n575 B.n574 71.676
R963 B.n580 B.n579 71.676
R964 B.n583 B.n582 71.676
R965 B.n588 B.n587 71.676
R966 B.n591 B.n590 71.676
R967 B.n596 B.n595 71.676
R968 B.n599 B.n598 71.676
R969 B.n604 B.n603 71.676
R970 B.n607 B.n606 71.676
R971 B.n612 B.n611 71.676
R972 B.n615 B.n614 71.676
R973 B.n623 B.n622 71.676
R974 B.n626 B.n625 71.676
R975 B.n631 B.n630 71.676
R976 B.n634 B.n633 71.676
R977 B.n639 B.n638 71.676
R978 B.n642 B.n641 71.676
R979 B.n648 B.n647 71.676
R980 B.n651 B.n650 71.676
R981 B.n656 B.n655 71.676
R982 B.n659 B.n658 71.676
R983 B.n664 B.n663 71.676
R984 B.n667 B.n666 71.676
R985 B.n672 B.n671 71.676
R986 B.n675 B.n674 71.676
R987 B.n680 B.n679 71.676
R988 B.n683 B.n682 71.676
R989 B.n688 B.n687 71.676
R990 B.n691 B.n690 71.676
R991 B.n696 B.n695 71.676
R992 B.n699 B.n698 71.676
R993 B.n704 B.n703 71.676
R994 B.n707 B.n706 71.676
R995 B.n712 B.n711 71.676
R996 B.n715 B.n714 71.676
R997 B.n720 B.n719 71.676
R998 B.n723 B.n722 71.676
R999 B.n728 B.n727 71.676
R1000 B.n731 B.n730 71.676
R1001 B.n736 B.n735 71.676
R1002 B.n739 B.n738 71.676
R1003 B.n744 B.n743 71.676
R1004 B.n747 B.n746 71.676
R1005 B.n752 B.n751 71.676
R1006 B.n755 B.n754 71.676
R1007 B.n760 B.n759 71.676
R1008 B.n763 B.n762 71.676
R1009 B.n48 B.n46 71.676
R1010 B.n123 B.n49 71.676
R1011 B.n127 B.n50 71.676
R1012 B.n131 B.n51 71.676
R1013 B.n135 B.n52 71.676
R1014 B.n139 B.n53 71.676
R1015 B.n143 B.n54 71.676
R1016 B.n147 B.n55 71.676
R1017 B.n151 B.n56 71.676
R1018 B.n155 B.n57 71.676
R1019 B.n159 B.n58 71.676
R1020 B.n163 B.n59 71.676
R1021 B.n167 B.n60 71.676
R1022 B.n171 B.n61 71.676
R1023 B.n175 B.n62 71.676
R1024 B.n179 B.n63 71.676
R1025 B.n183 B.n64 71.676
R1026 B.n187 B.n65 71.676
R1027 B.n191 B.n66 71.676
R1028 B.n195 B.n67 71.676
R1029 B.n199 B.n68 71.676
R1030 B.n203 B.n69 71.676
R1031 B.n207 B.n70 71.676
R1032 B.n211 B.n71 71.676
R1033 B.n215 B.n72 71.676
R1034 B.n219 B.n73 71.676
R1035 B.n223 B.n74 71.676
R1036 B.n227 B.n75 71.676
R1037 B.n231 B.n76 71.676
R1038 B.n235 B.n77 71.676
R1039 B.n239 B.n78 71.676
R1040 B.n243 B.n79 71.676
R1041 B.n247 B.n80 71.676
R1042 B.n251 B.n81 71.676
R1043 B.n255 B.n82 71.676
R1044 B.n259 B.n83 71.676
R1045 B.n263 B.n84 71.676
R1046 B.n267 B.n85 71.676
R1047 B.n271 B.n86 71.676
R1048 B.n275 B.n87 71.676
R1049 B.n279 B.n88 71.676
R1050 B.n283 B.n89 71.676
R1051 B.n287 B.n90 71.676
R1052 B.n291 B.n91 71.676
R1053 B.n295 B.n92 71.676
R1054 B.n299 B.n93 71.676
R1055 B.n303 B.n94 71.676
R1056 B.n307 B.n95 71.676
R1057 B.n311 B.n96 71.676
R1058 B.n315 B.n97 71.676
R1059 B.n319 B.n98 71.676
R1060 B.n323 B.n99 71.676
R1061 B.n327 B.n100 71.676
R1062 B.n331 B.n101 71.676
R1063 B.n335 B.n102 71.676
R1064 B.n339 B.n103 71.676
R1065 B.n343 B.n104 71.676
R1066 B.n347 B.n105 71.676
R1067 B.n351 B.n106 71.676
R1068 B.n355 B.n107 71.676
R1069 B.n359 B.n108 71.676
R1070 B.n363 B.n109 71.676
R1071 B.n367 B.n110 71.676
R1072 B.n371 B.n111 71.676
R1073 B.n375 B.n112 71.676
R1074 B.n379 B.n113 71.676
R1075 B.n875 B.n114 71.676
R1076 B.n875 B.n874 71.676
R1077 B.n381 B.n113 71.676
R1078 B.n378 B.n112 71.676
R1079 B.n374 B.n111 71.676
R1080 B.n370 B.n110 71.676
R1081 B.n366 B.n109 71.676
R1082 B.n362 B.n108 71.676
R1083 B.n358 B.n107 71.676
R1084 B.n354 B.n106 71.676
R1085 B.n350 B.n105 71.676
R1086 B.n346 B.n104 71.676
R1087 B.n342 B.n103 71.676
R1088 B.n338 B.n102 71.676
R1089 B.n334 B.n101 71.676
R1090 B.n330 B.n100 71.676
R1091 B.n326 B.n99 71.676
R1092 B.n322 B.n98 71.676
R1093 B.n318 B.n97 71.676
R1094 B.n314 B.n96 71.676
R1095 B.n310 B.n95 71.676
R1096 B.n306 B.n94 71.676
R1097 B.n302 B.n93 71.676
R1098 B.n298 B.n92 71.676
R1099 B.n294 B.n91 71.676
R1100 B.n290 B.n90 71.676
R1101 B.n286 B.n89 71.676
R1102 B.n282 B.n88 71.676
R1103 B.n278 B.n87 71.676
R1104 B.n274 B.n86 71.676
R1105 B.n270 B.n85 71.676
R1106 B.n266 B.n84 71.676
R1107 B.n262 B.n83 71.676
R1108 B.n258 B.n82 71.676
R1109 B.n254 B.n81 71.676
R1110 B.n250 B.n80 71.676
R1111 B.n246 B.n79 71.676
R1112 B.n242 B.n78 71.676
R1113 B.n238 B.n77 71.676
R1114 B.n234 B.n76 71.676
R1115 B.n230 B.n75 71.676
R1116 B.n226 B.n74 71.676
R1117 B.n222 B.n73 71.676
R1118 B.n218 B.n72 71.676
R1119 B.n214 B.n71 71.676
R1120 B.n210 B.n70 71.676
R1121 B.n206 B.n69 71.676
R1122 B.n202 B.n68 71.676
R1123 B.n198 B.n67 71.676
R1124 B.n194 B.n66 71.676
R1125 B.n190 B.n65 71.676
R1126 B.n186 B.n64 71.676
R1127 B.n182 B.n63 71.676
R1128 B.n178 B.n62 71.676
R1129 B.n174 B.n61 71.676
R1130 B.n170 B.n60 71.676
R1131 B.n166 B.n59 71.676
R1132 B.n162 B.n58 71.676
R1133 B.n158 B.n57 71.676
R1134 B.n154 B.n56 71.676
R1135 B.n150 B.n55 71.676
R1136 B.n146 B.n54 71.676
R1137 B.n142 B.n53 71.676
R1138 B.n138 B.n52 71.676
R1139 B.n134 B.n51 71.676
R1140 B.n130 B.n50 71.676
R1141 B.n126 B.n49 71.676
R1142 B.n122 B.n48 71.676
R1143 B.n500 B.n499 71.676
R1144 B.n502 B.n496 71.676
R1145 B.n509 B.n508 71.676
R1146 B.n510 B.n494 71.676
R1147 B.n517 B.n516 71.676
R1148 B.n518 B.n492 71.676
R1149 B.n525 B.n524 71.676
R1150 B.n526 B.n490 71.676
R1151 B.n533 B.n532 71.676
R1152 B.n534 B.n488 71.676
R1153 B.n541 B.n540 71.676
R1154 B.n542 B.n486 71.676
R1155 B.n549 B.n548 71.676
R1156 B.n550 B.n484 71.676
R1157 B.n557 B.n556 71.676
R1158 B.n558 B.n482 71.676
R1159 B.n565 B.n564 71.676
R1160 B.n566 B.n480 71.676
R1161 B.n573 B.n572 71.676
R1162 B.n574 B.n478 71.676
R1163 B.n581 B.n580 71.676
R1164 B.n582 B.n476 71.676
R1165 B.n589 B.n588 71.676
R1166 B.n590 B.n474 71.676
R1167 B.n597 B.n596 71.676
R1168 B.n598 B.n472 71.676
R1169 B.n605 B.n604 71.676
R1170 B.n606 B.n470 71.676
R1171 B.n613 B.n612 71.676
R1172 B.n614 B.n468 71.676
R1173 B.n624 B.n623 71.676
R1174 B.n625 B.n466 71.676
R1175 B.n632 B.n631 71.676
R1176 B.n633 B.n464 71.676
R1177 B.n640 B.n639 71.676
R1178 B.n641 B.n460 71.676
R1179 B.n649 B.n648 71.676
R1180 B.n650 B.n458 71.676
R1181 B.n657 B.n656 71.676
R1182 B.n658 B.n456 71.676
R1183 B.n665 B.n664 71.676
R1184 B.n666 B.n454 71.676
R1185 B.n673 B.n672 71.676
R1186 B.n674 B.n452 71.676
R1187 B.n681 B.n680 71.676
R1188 B.n682 B.n450 71.676
R1189 B.n689 B.n688 71.676
R1190 B.n690 B.n448 71.676
R1191 B.n697 B.n696 71.676
R1192 B.n698 B.n446 71.676
R1193 B.n705 B.n704 71.676
R1194 B.n706 B.n444 71.676
R1195 B.n713 B.n712 71.676
R1196 B.n714 B.n442 71.676
R1197 B.n721 B.n720 71.676
R1198 B.n722 B.n440 71.676
R1199 B.n729 B.n728 71.676
R1200 B.n730 B.n438 71.676
R1201 B.n737 B.n736 71.676
R1202 B.n738 B.n436 71.676
R1203 B.n745 B.n744 71.676
R1204 B.n746 B.n434 71.676
R1205 B.n753 B.n752 71.676
R1206 B.n754 B.n432 71.676
R1207 B.n761 B.n760 71.676
R1208 B.n764 B.n763 71.676
R1209 B.n462 B.t22 67.3837
R1210 B.n116 B.t13 67.3837
R1211 B.n619 B.t16 67.358
R1212 B.n119 B.t20 67.358
R1213 B.n644 B.n462 59.5399
R1214 B.n620 B.n619 59.5399
R1215 B.n120 B.n119 59.5399
R1216 B.n117 B.n116 59.5399
R1217 B.n769 B.n428 50.1958
R1218 B.n877 B.n876 50.1958
R1219 B.n879 B.n45 32.0005
R1220 B.n873 B.n872 32.0005
R1221 B.n767 B.n766 32.0005
R1222 B.n771 B.n426 32.0005
R1223 B.n769 B.n424 30.7508
R1224 B.n775 B.n424 30.7508
R1225 B.n775 B.n420 30.7508
R1226 B.n781 B.n420 30.7508
R1227 B.n787 B.n416 30.7508
R1228 B.n787 B.n412 30.7508
R1229 B.n793 B.n412 30.7508
R1230 B.n793 B.n408 30.7508
R1231 B.n799 B.n408 30.7508
R1232 B.n806 B.n404 30.7508
R1233 B.n806 B.n805 30.7508
R1234 B.n812 B.n400 30.7508
R1235 B.n818 B.n393 30.7508
R1236 B.n824 B.n393 30.7508
R1237 B.n832 B.n389 30.7508
R1238 B.n832 B.n831 30.7508
R1239 B.n838 B.n4 30.7508
R1240 B.n925 B.n4 30.7508
R1241 B.n925 B.n924 30.7508
R1242 B.n924 B.n923 30.7508
R1243 B.n917 B.n11 30.7508
R1244 B.n917 B.n916 30.7508
R1245 B.n915 B.n15 30.7508
R1246 B.n909 B.n15 30.7508
R1247 B.n908 B.n907 30.7508
R1248 B.n901 B.n25 30.7508
R1249 B.n901 B.n900 30.7508
R1250 B.n899 B.n29 30.7508
R1251 B.n893 B.n29 30.7508
R1252 B.n893 B.n892 30.7508
R1253 B.n892 B.n891 30.7508
R1254 B.n891 B.n36 30.7508
R1255 B.n885 B.n884 30.7508
R1256 B.n884 B.n883 30.7508
R1257 B.n883 B.n43 30.7508
R1258 B.n877 B.n43 30.7508
R1259 B.n838 B.t9 28.0375
R1260 B.n923 B.t7 28.0375
R1261 B.n400 B.t4 26.2287
R1262 B.t6 B.n908 26.2287
R1263 B.n781 B.t15 24.4198
R1264 B.n885 B.t11 24.4198
R1265 B.n812 B.t2 23.5154
R1266 B.n907 B.t1 23.5154
R1267 B.n799 B.t0 18.9933
R1268 B.t8 B.n899 18.9933
R1269 B B.n927 18.0485
R1270 B.n462 B.n461 17.2611
R1271 B.n619 B.n618 17.2611
R1272 B.n119 B.n118 17.2611
R1273 B.n116 B.n115 17.2611
R1274 B.t3 B.n389 16.28
R1275 B.n916 B.t5 16.28
R1276 B.n824 B.t3 14.4712
R1277 B.t5 B.n915 14.4712
R1278 B.t0 B.n404 11.758
R1279 B.n900 B.t8 11.758
R1280 B.n121 B.n45 10.6151
R1281 B.n124 B.n121 10.6151
R1282 B.n125 B.n124 10.6151
R1283 B.n128 B.n125 10.6151
R1284 B.n129 B.n128 10.6151
R1285 B.n132 B.n129 10.6151
R1286 B.n133 B.n132 10.6151
R1287 B.n136 B.n133 10.6151
R1288 B.n137 B.n136 10.6151
R1289 B.n140 B.n137 10.6151
R1290 B.n141 B.n140 10.6151
R1291 B.n144 B.n141 10.6151
R1292 B.n145 B.n144 10.6151
R1293 B.n148 B.n145 10.6151
R1294 B.n149 B.n148 10.6151
R1295 B.n152 B.n149 10.6151
R1296 B.n153 B.n152 10.6151
R1297 B.n156 B.n153 10.6151
R1298 B.n157 B.n156 10.6151
R1299 B.n160 B.n157 10.6151
R1300 B.n161 B.n160 10.6151
R1301 B.n164 B.n161 10.6151
R1302 B.n165 B.n164 10.6151
R1303 B.n168 B.n165 10.6151
R1304 B.n169 B.n168 10.6151
R1305 B.n172 B.n169 10.6151
R1306 B.n173 B.n172 10.6151
R1307 B.n176 B.n173 10.6151
R1308 B.n177 B.n176 10.6151
R1309 B.n180 B.n177 10.6151
R1310 B.n181 B.n180 10.6151
R1311 B.n184 B.n181 10.6151
R1312 B.n185 B.n184 10.6151
R1313 B.n188 B.n185 10.6151
R1314 B.n189 B.n188 10.6151
R1315 B.n192 B.n189 10.6151
R1316 B.n193 B.n192 10.6151
R1317 B.n196 B.n193 10.6151
R1318 B.n197 B.n196 10.6151
R1319 B.n200 B.n197 10.6151
R1320 B.n201 B.n200 10.6151
R1321 B.n204 B.n201 10.6151
R1322 B.n205 B.n204 10.6151
R1323 B.n208 B.n205 10.6151
R1324 B.n209 B.n208 10.6151
R1325 B.n212 B.n209 10.6151
R1326 B.n213 B.n212 10.6151
R1327 B.n216 B.n213 10.6151
R1328 B.n217 B.n216 10.6151
R1329 B.n220 B.n217 10.6151
R1330 B.n221 B.n220 10.6151
R1331 B.n224 B.n221 10.6151
R1332 B.n225 B.n224 10.6151
R1333 B.n228 B.n225 10.6151
R1334 B.n229 B.n228 10.6151
R1335 B.n232 B.n229 10.6151
R1336 B.n233 B.n232 10.6151
R1337 B.n236 B.n233 10.6151
R1338 B.n237 B.n236 10.6151
R1339 B.n240 B.n237 10.6151
R1340 B.n241 B.n240 10.6151
R1341 B.n245 B.n244 10.6151
R1342 B.n248 B.n245 10.6151
R1343 B.n249 B.n248 10.6151
R1344 B.n252 B.n249 10.6151
R1345 B.n253 B.n252 10.6151
R1346 B.n256 B.n253 10.6151
R1347 B.n257 B.n256 10.6151
R1348 B.n260 B.n257 10.6151
R1349 B.n261 B.n260 10.6151
R1350 B.n265 B.n264 10.6151
R1351 B.n268 B.n265 10.6151
R1352 B.n269 B.n268 10.6151
R1353 B.n272 B.n269 10.6151
R1354 B.n273 B.n272 10.6151
R1355 B.n276 B.n273 10.6151
R1356 B.n277 B.n276 10.6151
R1357 B.n280 B.n277 10.6151
R1358 B.n281 B.n280 10.6151
R1359 B.n284 B.n281 10.6151
R1360 B.n285 B.n284 10.6151
R1361 B.n288 B.n285 10.6151
R1362 B.n289 B.n288 10.6151
R1363 B.n292 B.n289 10.6151
R1364 B.n293 B.n292 10.6151
R1365 B.n296 B.n293 10.6151
R1366 B.n297 B.n296 10.6151
R1367 B.n300 B.n297 10.6151
R1368 B.n301 B.n300 10.6151
R1369 B.n304 B.n301 10.6151
R1370 B.n305 B.n304 10.6151
R1371 B.n308 B.n305 10.6151
R1372 B.n309 B.n308 10.6151
R1373 B.n312 B.n309 10.6151
R1374 B.n313 B.n312 10.6151
R1375 B.n316 B.n313 10.6151
R1376 B.n317 B.n316 10.6151
R1377 B.n320 B.n317 10.6151
R1378 B.n321 B.n320 10.6151
R1379 B.n324 B.n321 10.6151
R1380 B.n325 B.n324 10.6151
R1381 B.n328 B.n325 10.6151
R1382 B.n329 B.n328 10.6151
R1383 B.n332 B.n329 10.6151
R1384 B.n333 B.n332 10.6151
R1385 B.n336 B.n333 10.6151
R1386 B.n337 B.n336 10.6151
R1387 B.n340 B.n337 10.6151
R1388 B.n341 B.n340 10.6151
R1389 B.n344 B.n341 10.6151
R1390 B.n345 B.n344 10.6151
R1391 B.n348 B.n345 10.6151
R1392 B.n349 B.n348 10.6151
R1393 B.n352 B.n349 10.6151
R1394 B.n353 B.n352 10.6151
R1395 B.n356 B.n353 10.6151
R1396 B.n357 B.n356 10.6151
R1397 B.n360 B.n357 10.6151
R1398 B.n361 B.n360 10.6151
R1399 B.n364 B.n361 10.6151
R1400 B.n365 B.n364 10.6151
R1401 B.n368 B.n365 10.6151
R1402 B.n369 B.n368 10.6151
R1403 B.n372 B.n369 10.6151
R1404 B.n373 B.n372 10.6151
R1405 B.n376 B.n373 10.6151
R1406 B.n377 B.n376 10.6151
R1407 B.n380 B.n377 10.6151
R1408 B.n382 B.n380 10.6151
R1409 B.n383 B.n382 10.6151
R1410 B.n873 B.n383 10.6151
R1411 B.n767 B.n422 10.6151
R1412 B.n777 B.n422 10.6151
R1413 B.n778 B.n777 10.6151
R1414 B.n779 B.n778 10.6151
R1415 B.n779 B.n414 10.6151
R1416 B.n789 B.n414 10.6151
R1417 B.n790 B.n789 10.6151
R1418 B.n791 B.n790 10.6151
R1419 B.n791 B.n406 10.6151
R1420 B.n801 B.n406 10.6151
R1421 B.n802 B.n801 10.6151
R1422 B.n803 B.n802 10.6151
R1423 B.n803 B.n398 10.6151
R1424 B.n814 B.n398 10.6151
R1425 B.n815 B.n814 10.6151
R1426 B.n816 B.n815 10.6151
R1427 B.n816 B.n391 10.6151
R1428 B.n826 B.n391 10.6151
R1429 B.n827 B.n826 10.6151
R1430 B.n829 B.n827 10.6151
R1431 B.n829 B.n828 10.6151
R1432 B.n828 B.n384 10.6151
R1433 B.n841 B.n384 10.6151
R1434 B.n842 B.n841 10.6151
R1435 B.n843 B.n842 10.6151
R1436 B.n844 B.n843 10.6151
R1437 B.n846 B.n844 10.6151
R1438 B.n847 B.n846 10.6151
R1439 B.n848 B.n847 10.6151
R1440 B.n849 B.n848 10.6151
R1441 B.n851 B.n849 10.6151
R1442 B.n852 B.n851 10.6151
R1443 B.n853 B.n852 10.6151
R1444 B.n854 B.n853 10.6151
R1445 B.n856 B.n854 10.6151
R1446 B.n857 B.n856 10.6151
R1447 B.n858 B.n857 10.6151
R1448 B.n859 B.n858 10.6151
R1449 B.n861 B.n859 10.6151
R1450 B.n862 B.n861 10.6151
R1451 B.n863 B.n862 10.6151
R1452 B.n864 B.n863 10.6151
R1453 B.n866 B.n864 10.6151
R1454 B.n867 B.n866 10.6151
R1455 B.n868 B.n867 10.6151
R1456 B.n869 B.n868 10.6151
R1457 B.n871 B.n869 10.6151
R1458 B.n872 B.n871 10.6151
R1459 B.n498 B.n426 10.6151
R1460 B.n498 B.n497 10.6151
R1461 B.n504 B.n497 10.6151
R1462 B.n505 B.n504 10.6151
R1463 B.n506 B.n505 10.6151
R1464 B.n506 B.n495 10.6151
R1465 B.n512 B.n495 10.6151
R1466 B.n513 B.n512 10.6151
R1467 B.n514 B.n513 10.6151
R1468 B.n514 B.n493 10.6151
R1469 B.n520 B.n493 10.6151
R1470 B.n521 B.n520 10.6151
R1471 B.n522 B.n521 10.6151
R1472 B.n522 B.n491 10.6151
R1473 B.n528 B.n491 10.6151
R1474 B.n529 B.n528 10.6151
R1475 B.n530 B.n529 10.6151
R1476 B.n530 B.n489 10.6151
R1477 B.n536 B.n489 10.6151
R1478 B.n537 B.n536 10.6151
R1479 B.n538 B.n537 10.6151
R1480 B.n538 B.n487 10.6151
R1481 B.n544 B.n487 10.6151
R1482 B.n545 B.n544 10.6151
R1483 B.n546 B.n545 10.6151
R1484 B.n546 B.n485 10.6151
R1485 B.n552 B.n485 10.6151
R1486 B.n553 B.n552 10.6151
R1487 B.n554 B.n553 10.6151
R1488 B.n554 B.n483 10.6151
R1489 B.n560 B.n483 10.6151
R1490 B.n561 B.n560 10.6151
R1491 B.n562 B.n561 10.6151
R1492 B.n562 B.n481 10.6151
R1493 B.n568 B.n481 10.6151
R1494 B.n569 B.n568 10.6151
R1495 B.n570 B.n569 10.6151
R1496 B.n570 B.n479 10.6151
R1497 B.n576 B.n479 10.6151
R1498 B.n577 B.n576 10.6151
R1499 B.n578 B.n577 10.6151
R1500 B.n578 B.n477 10.6151
R1501 B.n584 B.n477 10.6151
R1502 B.n585 B.n584 10.6151
R1503 B.n586 B.n585 10.6151
R1504 B.n586 B.n475 10.6151
R1505 B.n592 B.n475 10.6151
R1506 B.n593 B.n592 10.6151
R1507 B.n594 B.n593 10.6151
R1508 B.n594 B.n473 10.6151
R1509 B.n600 B.n473 10.6151
R1510 B.n601 B.n600 10.6151
R1511 B.n602 B.n601 10.6151
R1512 B.n602 B.n471 10.6151
R1513 B.n608 B.n471 10.6151
R1514 B.n609 B.n608 10.6151
R1515 B.n610 B.n609 10.6151
R1516 B.n610 B.n469 10.6151
R1517 B.n616 B.n469 10.6151
R1518 B.n617 B.n616 10.6151
R1519 B.n621 B.n617 10.6151
R1520 B.n627 B.n467 10.6151
R1521 B.n628 B.n627 10.6151
R1522 B.n629 B.n628 10.6151
R1523 B.n629 B.n465 10.6151
R1524 B.n635 B.n465 10.6151
R1525 B.n636 B.n635 10.6151
R1526 B.n637 B.n636 10.6151
R1527 B.n637 B.n463 10.6151
R1528 B.n643 B.n463 10.6151
R1529 B.n646 B.n645 10.6151
R1530 B.n646 B.n459 10.6151
R1531 B.n652 B.n459 10.6151
R1532 B.n653 B.n652 10.6151
R1533 B.n654 B.n653 10.6151
R1534 B.n654 B.n457 10.6151
R1535 B.n660 B.n457 10.6151
R1536 B.n661 B.n660 10.6151
R1537 B.n662 B.n661 10.6151
R1538 B.n662 B.n455 10.6151
R1539 B.n668 B.n455 10.6151
R1540 B.n669 B.n668 10.6151
R1541 B.n670 B.n669 10.6151
R1542 B.n670 B.n453 10.6151
R1543 B.n676 B.n453 10.6151
R1544 B.n677 B.n676 10.6151
R1545 B.n678 B.n677 10.6151
R1546 B.n678 B.n451 10.6151
R1547 B.n684 B.n451 10.6151
R1548 B.n685 B.n684 10.6151
R1549 B.n686 B.n685 10.6151
R1550 B.n686 B.n449 10.6151
R1551 B.n692 B.n449 10.6151
R1552 B.n693 B.n692 10.6151
R1553 B.n694 B.n693 10.6151
R1554 B.n694 B.n447 10.6151
R1555 B.n700 B.n447 10.6151
R1556 B.n701 B.n700 10.6151
R1557 B.n702 B.n701 10.6151
R1558 B.n702 B.n445 10.6151
R1559 B.n708 B.n445 10.6151
R1560 B.n709 B.n708 10.6151
R1561 B.n710 B.n709 10.6151
R1562 B.n710 B.n443 10.6151
R1563 B.n716 B.n443 10.6151
R1564 B.n717 B.n716 10.6151
R1565 B.n718 B.n717 10.6151
R1566 B.n718 B.n441 10.6151
R1567 B.n724 B.n441 10.6151
R1568 B.n725 B.n724 10.6151
R1569 B.n726 B.n725 10.6151
R1570 B.n726 B.n439 10.6151
R1571 B.n732 B.n439 10.6151
R1572 B.n733 B.n732 10.6151
R1573 B.n734 B.n733 10.6151
R1574 B.n734 B.n437 10.6151
R1575 B.n740 B.n437 10.6151
R1576 B.n741 B.n740 10.6151
R1577 B.n742 B.n741 10.6151
R1578 B.n742 B.n435 10.6151
R1579 B.n748 B.n435 10.6151
R1580 B.n749 B.n748 10.6151
R1581 B.n750 B.n749 10.6151
R1582 B.n750 B.n433 10.6151
R1583 B.n756 B.n433 10.6151
R1584 B.n757 B.n756 10.6151
R1585 B.n758 B.n757 10.6151
R1586 B.n758 B.n431 10.6151
R1587 B.n431 B.n430 10.6151
R1588 B.n765 B.n430 10.6151
R1589 B.n766 B.n765 10.6151
R1590 B.n772 B.n771 10.6151
R1591 B.n773 B.n772 10.6151
R1592 B.n773 B.n418 10.6151
R1593 B.n783 B.n418 10.6151
R1594 B.n784 B.n783 10.6151
R1595 B.n785 B.n784 10.6151
R1596 B.n785 B.n410 10.6151
R1597 B.n795 B.n410 10.6151
R1598 B.n796 B.n795 10.6151
R1599 B.n797 B.n796 10.6151
R1600 B.n797 B.n402 10.6151
R1601 B.n808 B.n402 10.6151
R1602 B.n809 B.n808 10.6151
R1603 B.n810 B.n809 10.6151
R1604 B.n810 B.n395 10.6151
R1605 B.n820 B.n395 10.6151
R1606 B.n821 B.n820 10.6151
R1607 B.n822 B.n821 10.6151
R1608 B.n822 B.n387 10.6151
R1609 B.n834 B.n387 10.6151
R1610 B.n835 B.n834 10.6151
R1611 B.n836 B.n835 10.6151
R1612 B.n836 B.n0 10.6151
R1613 B.n921 B.n1 10.6151
R1614 B.n921 B.n920 10.6151
R1615 B.n920 B.n919 10.6151
R1616 B.n919 B.n9 10.6151
R1617 B.n913 B.n9 10.6151
R1618 B.n913 B.n912 10.6151
R1619 B.n912 B.n911 10.6151
R1620 B.n911 B.n17 10.6151
R1621 B.n905 B.n17 10.6151
R1622 B.n905 B.n904 10.6151
R1623 B.n904 B.n903 10.6151
R1624 B.n903 B.n23 10.6151
R1625 B.n897 B.n23 10.6151
R1626 B.n897 B.n896 10.6151
R1627 B.n896 B.n895 10.6151
R1628 B.n895 B.n31 10.6151
R1629 B.n889 B.n31 10.6151
R1630 B.n889 B.n888 10.6151
R1631 B.n888 B.n887 10.6151
R1632 B.n887 B.n38 10.6151
R1633 B.n881 B.n38 10.6151
R1634 B.n881 B.n880 10.6151
R1635 B.n880 B.n879 10.6151
R1636 B.n241 B.n120 9.36635
R1637 B.n264 B.n117 9.36635
R1638 B.n621 B.n620 9.36635
R1639 B.n645 B.n644 9.36635
R1640 B.n805 B.t2 7.23585
R1641 B.n25 B.t1 7.23585
R1642 B.t15 B.n416 6.33144
R1643 B.t11 B.n36 6.33144
R1644 B.n818 B.t4 4.5226
R1645 B.n909 B.t6 4.5226
R1646 B.n927 B.n0 2.81026
R1647 B.n927 B.n1 2.81026
R1648 B.n831 B.t9 2.71376
R1649 B.n11 B.t7 2.71376
R1650 B.n244 B.n120 1.24928
R1651 B.n261 B.n117 1.24928
R1652 B.n620 B.n467 1.24928
R1653 B.n644 B.n643 1.24928
R1654 VN.n3 VN.t4 914.61
R1655 VN.n13 VN.t7 914.61
R1656 VN.n2 VN.t3 890.409
R1657 VN.n1 VN.t6 890.409
R1658 VN.n6 VN.t1 890.409
R1659 VN.n8 VN.t9 890.409
R1660 VN.n12 VN.t2 890.409
R1661 VN.n11 VN.t5 890.409
R1662 VN.n16 VN.t0 890.409
R1663 VN.n18 VN.t8 890.409
R1664 VN.n9 VN.n8 161.3
R1665 VN.n19 VN.n18 161.3
R1666 VN.n17 VN.n10 161.3
R1667 VN.n16 VN.n15 161.3
R1668 VN.n7 VN.n0 161.3
R1669 VN.n6 VN.n5 161.3
R1670 VN.n14 VN.n11 80.6037
R1671 VN.n4 VN.n1 80.6037
R1672 VN.n2 VN.n1 48.2005
R1673 VN.n6 VN.n1 48.2005
R1674 VN.n12 VN.n11 48.2005
R1675 VN.n16 VN.n11 48.2005
R1676 VN VN.n19 47.688
R1677 VN.n14 VN.n13 45.0238
R1678 VN.n4 VN.n3 45.0238
R1679 VN.n8 VN.n7 36.5157
R1680 VN.n18 VN.n17 36.5157
R1681 VN.n3 VN.n2 17.2829
R1682 VN.n13 VN.n12 17.2829
R1683 VN.n7 VN.n6 11.6853
R1684 VN.n17 VN.n16 11.6853
R1685 VN.n15 VN.n14 0.285035
R1686 VN.n5 VN.n4 0.285035
R1687 VN.n19 VN.n10 0.189894
R1688 VN.n15 VN.n10 0.189894
R1689 VN.n5 VN.n0 0.189894
R1690 VN.n9 VN.n0 0.189894
R1691 VN VN.n9 0.0516364
R1692 VDD2.n1 VDD2.t5 63.7515
R1693 VDD2.n4 VDD2.t1 62.9843
R1694 VDD2.n3 VDD2.n2 62.4639
R1695 VDD2 VDD2.n7 62.4621
R1696 VDD2.n6 VDD2.n5 61.945
R1697 VDD2.n1 VDD2.n0 61.9438
R1698 VDD2.n4 VDD2.n3 43.7821
R1699 VDD2.n7 VDD2.t7 1.03987
R1700 VDD2.n7 VDD2.t2 1.03987
R1701 VDD2.n5 VDD2.t9 1.03987
R1702 VDD2.n5 VDD2.t4 1.03987
R1703 VDD2.n2 VDD2.t8 1.03987
R1704 VDD2.n2 VDD2.t0 1.03987
R1705 VDD2.n0 VDD2.t6 1.03987
R1706 VDD2.n0 VDD2.t3 1.03987
R1707 VDD2.n6 VDD2.n4 0.767741
R1708 VDD2 VDD2.n6 0.2505
R1709 VDD2.n3 VDD2.n1 0.136964
C0 VN VP 6.70038f
C1 VDD2 VTAIL 23.5723f
C2 VDD2 VDD1 0.887319f
C3 VDD2 VN 9.13098f
C4 VDD1 VTAIL 23.543901f
C5 VDD2 VP 0.324899f
C6 VTAIL VN 8.61095f
C7 VTAIL VP 8.62593f
C8 VDD1 VN 0.148673f
C9 VDD1 VP 9.29974f
C10 VDD2 B 6.068377f
C11 VDD1 B 5.98175f
C12 VTAIL B 8.910639f
C13 VN B 9.728089f
C14 VP B 7.306675f
C15 VDD2.t5 B 4.50184f
C16 VDD2.t6 B 0.384528f
C17 VDD2.t3 B 0.384528f
C18 VDD2.n0 B 3.51796f
C19 VDD2.n1 B 0.628753f
C20 VDD2.t8 B 0.384528f
C21 VDD2.t0 B 0.384528f
C22 VDD2.n2 B 3.52065f
C23 VDD2.n3 B 2.30981f
C24 VDD2.t1 B 4.49767f
C25 VDD2.n4 B 2.93652f
C26 VDD2.t9 B 0.384528f
C27 VDD2.t4 B 0.384528f
C28 VDD2.n5 B 3.51797f
C29 VDD2.n6 B 0.289599f
C30 VDD2.t7 B 0.384528f
C31 VDD2.t2 B 0.384528f
C32 VDD2.n7 B 3.52061f
C33 VN.n0 B 0.045704f
C34 VN.t6 B 1.38169f
C35 VN.n1 B 0.531196f
C36 VN.t4 B 1.39545f
C37 VN.t3 B 1.38169f
C38 VN.n2 B 0.529134f
C39 VN.n3 B 0.510412f
C40 VN.n4 B 0.215331f
C41 VN.n5 B 0.060986f
C42 VN.t1 B 1.38169f
C43 VN.n6 B 0.523079f
C44 VN.n7 B 0.010371f
C45 VN.t9 B 1.38169f
C46 VN.n8 B 0.51857f
C47 VN.n9 B 0.035419f
C48 VN.n10 B 0.045704f
C49 VN.t5 B 1.38169f
C50 VN.n11 B 0.531196f
C51 VN.t0 B 1.38169f
C52 VN.t7 B 1.39545f
C53 VN.t2 B 1.38169f
C54 VN.n12 B 0.529134f
C55 VN.n13 B 0.510412f
C56 VN.n14 B 0.215331f
C57 VN.n15 B 0.060986f
C58 VN.n16 B 0.523079f
C59 VN.n17 B 0.010371f
C60 VN.t8 B 1.38169f
C61 VN.n18 B 0.51857f
C62 VN.n19 B 2.31331f
C63 VTAIL.t17 B 0.391955f
C64 VTAIL.t5 B 0.391955f
C65 VTAIL.n0 B 3.51041f
C66 VTAIL.n1 B 0.374726f
C67 VTAIL.t14 B 4.48537f
C68 VTAIL.n2 B 0.479945f
C69 VTAIL.t7 B 0.391955f
C70 VTAIL.t15 B 0.391955f
C71 VTAIL.n3 B 3.51041f
C72 VTAIL.n4 B 0.378704f
C73 VTAIL.t10 B 0.391955f
C74 VTAIL.t9 B 0.391955f
C75 VTAIL.n5 B 3.51041f
C76 VTAIL.n6 B 2.17453f
C77 VTAIL.t0 B 0.391955f
C78 VTAIL.t2 B 0.391955f
C79 VTAIL.n7 B 3.51042f
C80 VTAIL.n8 B 2.17452f
C81 VTAIL.t4 B 0.391955f
C82 VTAIL.t3 B 0.391955f
C83 VTAIL.n9 B 3.51042f
C84 VTAIL.n10 B 0.378693f
C85 VTAIL.t16 B 4.4854f
C86 VTAIL.n11 B 0.479912f
C87 VTAIL.t12 B 0.391955f
C88 VTAIL.t6 B 0.391955f
C89 VTAIL.n12 B 3.51042f
C90 VTAIL.n13 B 0.385926f
C91 VTAIL.t11 B 0.391955f
C92 VTAIL.t8 B 0.391955f
C93 VTAIL.n14 B 3.51042f
C94 VTAIL.n15 B 0.378693f
C95 VTAIL.t13 B 4.48537f
C96 VTAIL.n16 B 2.20417f
C97 VTAIL.t19 B 4.48537f
C98 VTAIL.n17 B 2.20417f
C99 VTAIL.t18 B 0.391955f
C100 VTAIL.t1 B 0.391955f
C101 VTAIL.n18 B 3.51041f
C102 VTAIL.n19 B 0.325545f
C103 VDD1.t2 B 4.50264f
C104 VDD1.t8 B 0.384595f
C105 VDD1.t7 B 0.384595f
C106 VDD1.n0 B 3.51857f
C107 VDD1.n1 B 0.633837f
C108 VDD1.t6 B 4.50261f
C109 VDD1.t5 B 0.384595f
C110 VDD1.t9 B 0.384595f
C111 VDD1.n2 B 3.51857f
C112 VDD1.n3 B 0.628861f
C113 VDD1.t1 B 0.384595f
C114 VDD1.t0 B 0.384595f
C115 VDD1.n4 B 3.52126f
C116 VDD1.n5 B 2.38708f
C117 VDD1.t4 B 0.384595f
C118 VDD1.t3 B 0.384595f
C119 VDD1.n6 B 3.51855f
C120 VDD1.n7 B 2.92809f
C121 VP.n0 B 0.0462f
C122 VP.t8 B 1.39669f
C123 VP.n1 B 0.536963f
C124 VP.n2 B 0.0462f
C125 VP.n3 B 0.0462f
C126 VP.t2 B 1.39669f
C127 VP.t7 B 1.39669f
C128 VP.n4 B 0.061648f
C129 VP.t4 B 1.39669f
C130 VP.n5 B 0.217669f
C131 VP.t9 B 1.39669f
C132 VP.t3 B 1.4106f
C133 VP.n6 B 0.515954f
C134 VP.n7 B 0.534879f
C135 VP.n8 B 0.536963f
C136 VP.n9 B 0.528758f
C137 VP.n10 B 0.010484f
C138 VP.n11 B 0.524201f
C139 VP.n12 B 2.30831f
C140 VP.n13 B 2.34341f
C141 VP.t5 B 1.39669f
C142 VP.n14 B 0.524201f
C143 VP.n15 B 0.010484f
C144 VP.t6 B 1.39669f
C145 VP.n16 B 0.528758f
C146 VP.n17 B 0.061648f
C147 VP.n18 B 0.061504f
C148 VP.n19 B 0.061648f
C149 VP.t0 B 1.39669f
C150 VP.n20 B 0.528758f
C151 VP.n21 B 0.010484f
C152 VP.t1 B 1.39669f
C153 VP.n22 B 0.524201f
C154 VP.n23 B 0.035803f
.ends

