* NGSPICE file created from diff_pair_sample_0796.ext - technology: sky130A

.subckt diff_pair_sample_0796 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=1.47
X1 VTAIL.t11 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=1.47
X2 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=1.47
X3 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=1.47
X4 VDD2.t4 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=1.47
X5 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=1.47
X6 VDD2.t3 VN.t2 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=1.47
X7 VTAIL.t9 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=1.47
X8 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=1.47
X9 VDD1.t2 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=1.47
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=1.47
X11 VDD2.t1 VN.t4 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=1.47
X12 VTAIL.t8 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=1.47
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=1.47
X14 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=1.47
X15 VTAIL.t3 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=1.47
R0 VN.n3 VN.t2 363.995
R1 VN.n13 VN.t4 363.995
R2 VN.n2 VN.t5 327.072
R3 VN.n8 VN.t1 327.072
R4 VN.n12 VN.t3 327.072
R5 VN.n18 VN.t0 327.072
R6 VN.n9 VN.n8 171.088
R7 VN.n19 VN.n18 171.088
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN VN.n19 50.6388
R15 VN.n6 VN.n1 50.2061
R16 VN.n16 VN.n11 50.2061
R17 VN.n3 VN.n2 41.8683
R18 VN.n13 VN.n12 41.8683
R19 VN.n7 VN.n6 30.7807
R20 VN.n17 VN.n16 30.7807
R21 VN.n2 VN.n1 24.4675
R22 VN.n12 VN.n11 24.4675
R23 VN.n14 VN.n13 17.2768
R24 VN.n4 VN.n3 17.2768
R25 VN.n8 VN.n7 14.6807
R26 VN.n18 VN.n17 14.6807
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VTAIL.n10 VTAIL.t4 43.1624
R35 VTAIL.n7 VTAIL.t7 43.1624
R36 VTAIL.n11 VTAIL.t10 43.1623
R37 VTAIL.n2 VTAIL.t0 43.1623
R38 VTAIL.n9 VTAIL.n8 42.17
R39 VTAIL.n6 VTAIL.n5 42.17
R40 VTAIL.n1 VTAIL.n0 42.1699
R41 VTAIL.n4 VTAIL.n3 42.1699
R42 VTAIL.n6 VTAIL.n4 32.6686
R43 VTAIL.n11 VTAIL.n10 31.1169
R44 VTAIL.n7 VTAIL.n6 1.55222
R45 VTAIL.n10 VTAIL.n9 1.55222
R46 VTAIL.n4 VTAIL.n2 1.55222
R47 VTAIL.n9 VTAIL.n7 1.24619
R48 VTAIL.n2 VTAIL.n1 1.24619
R49 VTAIL VTAIL.n11 1.1061
R50 VTAIL.n0 VTAIL.t6 0.992981
R51 VTAIL.n0 VTAIL.t8 0.992981
R52 VTAIL.n3 VTAIL.t2 0.992981
R53 VTAIL.n3 VTAIL.t3 0.992981
R54 VTAIL.n8 VTAIL.t1 0.992981
R55 VTAIL.n8 VTAIL.t11 0.992981
R56 VTAIL.n5 VTAIL.t5 0.992981
R57 VTAIL.n5 VTAIL.t9 0.992981
R58 VTAIL VTAIL.n1 0.446621
R59 VDD2.n1 VDD2.t3 60.9495
R60 VDD2.n2 VDD2.t5 59.8412
R61 VDD2.n1 VDD2.n0 59.1813
R62 VDD2 VDD2.n3 59.1785
R63 VDD2.n2 VDD2.n1 45.9567
R64 VDD2 VDD2.n2 1.22248
R65 VDD2.n3 VDD2.t2 0.992981
R66 VDD2.n3 VDD2.t1 0.992981
R67 VDD2.n0 VDD2.t0 0.992981
R68 VDD2.n0 VDD2.t4 0.992981
R69 B.n945 B.n944 585
R70 B.n408 B.n125 585
R71 B.n407 B.n406 585
R72 B.n405 B.n404 585
R73 B.n403 B.n402 585
R74 B.n401 B.n400 585
R75 B.n399 B.n398 585
R76 B.n397 B.n396 585
R77 B.n395 B.n394 585
R78 B.n393 B.n392 585
R79 B.n391 B.n390 585
R80 B.n389 B.n388 585
R81 B.n387 B.n386 585
R82 B.n385 B.n384 585
R83 B.n383 B.n382 585
R84 B.n381 B.n380 585
R85 B.n379 B.n378 585
R86 B.n377 B.n376 585
R87 B.n375 B.n374 585
R88 B.n373 B.n372 585
R89 B.n371 B.n370 585
R90 B.n369 B.n368 585
R91 B.n367 B.n366 585
R92 B.n365 B.n364 585
R93 B.n363 B.n362 585
R94 B.n361 B.n360 585
R95 B.n359 B.n358 585
R96 B.n357 B.n356 585
R97 B.n355 B.n354 585
R98 B.n353 B.n352 585
R99 B.n351 B.n350 585
R100 B.n349 B.n348 585
R101 B.n347 B.n346 585
R102 B.n345 B.n344 585
R103 B.n343 B.n342 585
R104 B.n341 B.n340 585
R105 B.n339 B.n338 585
R106 B.n337 B.n336 585
R107 B.n335 B.n334 585
R108 B.n333 B.n332 585
R109 B.n331 B.n330 585
R110 B.n329 B.n328 585
R111 B.n327 B.n326 585
R112 B.n325 B.n324 585
R113 B.n323 B.n322 585
R114 B.n321 B.n320 585
R115 B.n319 B.n318 585
R116 B.n317 B.n316 585
R117 B.n315 B.n314 585
R118 B.n313 B.n312 585
R119 B.n311 B.n310 585
R120 B.n309 B.n308 585
R121 B.n307 B.n306 585
R122 B.n305 B.n304 585
R123 B.n303 B.n302 585
R124 B.n301 B.n300 585
R125 B.n299 B.n298 585
R126 B.n297 B.n296 585
R127 B.n295 B.n294 585
R128 B.n293 B.n292 585
R129 B.n291 B.n290 585
R130 B.n289 B.n288 585
R131 B.n287 B.n286 585
R132 B.n285 B.n284 585
R133 B.n283 B.n282 585
R134 B.n280 B.n279 585
R135 B.n278 B.n277 585
R136 B.n276 B.n275 585
R137 B.n274 B.n273 585
R138 B.n272 B.n271 585
R139 B.n270 B.n269 585
R140 B.n268 B.n267 585
R141 B.n266 B.n265 585
R142 B.n264 B.n263 585
R143 B.n262 B.n261 585
R144 B.n259 B.n258 585
R145 B.n257 B.n256 585
R146 B.n255 B.n254 585
R147 B.n253 B.n252 585
R148 B.n251 B.n250 585
R149 B.n249 B.n248 585
R150 B.n247 B.n246 585
R151 B.n245 B.n244 585
R152 B.n243 B.n242 585
R153 B.n241 B.n240 585
R154 B.n239 B.n238 585
R155 B.n237 B.n236 585
R156 B.n235 B.n234 585
R157 B.n233 B.n232 585
R158 B.n231 B.n230 585
R159 B.n229 B.n228 585
R160 B.n227 B.n226 585
R161 B.n225 B.n224 585
R162 B.n223 B.n222 585
R163 B.n221 B.n220 585
R164 B.n219 B.n218 585
R165 B.n217 B.n216 585
R166 B.n215 B.n214 585
R167 B.n213 B.n212 585
R168 B.n211 B.n210 585
R169 B.n209 B.n208 585
R170 B.n207 B.n206 585
R171 B.n205 B.n204 585
R172 B.n203 B.n202 585
R173 B.n201 B.n200 585
R174 B.n199 B.n198 585
R175 B.n197 B.n196 585
R176 B.n195 B.n194 585
R177 B.n193 B.n192 585
R178 B.n191 B.n190 585
R179 B.n189 B.n188 585
R180 B.n187 B.n186 585
R181 B.n185 B.n184 585
R182 B.n183 B.n182 585
R183 B.n181 B.n180 585
R184 B.n179 B.n178 585
R185 B.n177 B.n176 585
R186 B.n175 B.n174 585
R187 B.n173 B.n172 585
R188 B.n171 B.n170 585
R189 B.n169 B.n168 585
R190 B.n167 B.n166 585
R191 B.n165 B.n164 585
R192 B.n163 B.n162 585
R193 B.n161 B.n160 585
R194 B.n159 B.n158 585
R195 B.n157 B.n156 585
R196 B.n155 B.n154 585
R197 B.n153 B.n152 585
R198 B.n151 B.n150 585
R199 B.n149 B.n148 585
R200 B.n147 B.n146 585
R201 B.n145 B.n144 585
R202 B.n143 B.n142 585
R203 B.n141 B.n140 585
R204 B.n139 B.n138 585
R205 B.n137 B.n136 585
R206 B.n135 B.n134 585
R207 B.n133 B.n132 585
R208 B.n131 B.n130 585
R209 B.n943 B.n55 585
R210 B.n948 B.n55 585
R211 B.n942 B.n54 585
R212 B.n949 B.n54 585
R213 B.n941 B.n940 585
R214 B.n940 B.n50 585
R215 B.n939 B.n49 585
R216 B.n955 B.n49 585
R217 B.n938 B.n48 585
R218 B.n956 B.n48 585
R219 B.n937 B.n47 585
R220 B.n957 B.n47 585
R221 B.n936 B.n935 585
R222 B.n935 B.n43 585
R223 B.n934 B.n42 585
R224 B.n963 B.n42 585
R225 B.n933 B.n41 585
R226 B.n964 B.n41 585
R227 B.n932 B.n40 585
R228 B.n965 B.n40 585
R229 B.n931 B.n930 585
R230 B.n930 B.n36 585
R231 B.n929 B.n35 585
R232 B.n971 B.n35 585
R233 B.n928 B.n34 585
R234 B.n972 B.n34 585
R235 B.n927 B.n33 585
R236 B.n973 B.n33 585
R237 B.n926 B.n925 585
R238 B.n925 B.n32 585
R239 B.n924 B.n28 585
R240 B.n979 B.n28 585
R241 B.n923 B.n27 585
R242 B.n980 B.n27 585
R243 B.n922 B.n26 585
R244 B.n981 B.n26 585
R245 B.n921 B.n920 585
R246 B.n920 B.n22 585
R247 B.n919 B.n21 585
R248 B.n987 B.n21 585
R249 B.n918 B.n20 585
R250 B.n988 B.n20 585
R251 B.n917 B.n19 585
R252 B.n989 B.n19 585
R253 B.n916 B.n915 585
R254 B.n915 B.n15 585
R255 B.n914 B.n14 585
R256 B.n995 B.n14 585
R257 B.n913 B.n13 585
R258 B.n996 B.n13 585
R259 B.n912 B.n12 585
R260 B.n997 B.n12 585
R261 B.n911 B.n910 585
R262 B.n910 B.n8 585
R263 B.n909 B.n7 585
R264 B.n1003 B.n7 585
R265 B.n908 B.n6 585
R266 B.n1004 B.n6 585
R267 B.n907 B.n5 585
R268 B.n1005 B.n5 585
R269 B.n906 B.n905 585
R270 B.n905 B.n4 585
R271 B.n904 B.n409 585
R272 B.n904 B.n903 585
R273 B.n894 B.n410 585
R274 B.n411 B.n410 585
R275 B.n896 B.n895 585
R276 B.n897 B.n896 585
R277 B.n893 B.n415 585
R278 B.n419 B.n415 585
R279 B.n892 B.n891 585
R280 B.n891 B.n890 585
R281 B.n417 B.n416 585
R282 B.n418 B.n417 585
R283 B.n883 B.n882 585
R284 B.n884 B.n883 585
R285 B.n881 B.n424 585
R286 B.n424 B.n423 585
R287 B.n880 B.n879 585
R288 B.n879 B.n878 585
R289 B.n426 B.n425 585
R290 B.n427 B.n426 585
R291 B.n871 B.n870 585
R292 B.n872 B.n871 585
R293 B.n869 B.n432 585
R294 B.n432 B.n431 585
R295 B.n868 B.n867 585
R296 B.n867 B.n866 585
R297 B.n434 B.n433 585
R298 B.n859 B.n434 585
R299 B.n858 B.n857 585
R300 B.n860 B.n858 585
R301 B.n856 B.n439 585
R302 B.n439 B.n438 585
R303 B.n855 B.n854 585
R304 B.n854 B.n853 585
R305 B.n441 B.n440 585
R306 B.n442 B.n441 585
R307 B.n846 B.n845 585
R308 B.n847 B.n846 585
R309 B.n844 B.n447 585
R310 B.n447 B.n446 585
R311 B.n843 B.n842 585
R312 B.n842 B.n841 585
R313 B.n449 B.n448 585
R314 B.n450 B.n449 585
R315 B.n834 B.n833 585
R316 B.n835 B.n834 585
R317 B.n832 B.n455 585
R318 B.n455 B.n454 585
R319 B.n831 B.n830 585
R320 B.n830 B.n829 585
R321 B.n457 B.n456 585
R322 B.n458 B.n457 585
R323 B.n822 B.n821 585
R324 B.n823 B.n822 585
R325 B.n820 B.n463 585
R326 B.n463 B.n462 585
R327 B.n815 B.n814 585
R328 B.n813 B.n535 585
R329 B.n812 B.n534 585
R330 B.n817 B.n534 585
R331 B.n811 B.n810 585
R332 B.n809 B.n808 585
R333 B.n807 B.n806 585
R334 B.n805 B.n804 585
R335 B.n803 B.n802 585
R336 B.n801 B.n800 585
R337 B.n799 B.n798 585
R338 B.n797 B.n796 585
R339 B.n795 B.n794 585
R340 B.n793 B.n792 585
R341 B.n791 B.n790 585
R342 B.n789 B.n788 585
R343 B.n787 B.n786 585
R344 B.n785 B.n784 585
R345 B.n783 B.n782 585
R346 B.n781 B.n780 585
R347 B.n779 B.n778 585
R348 B.n777 B.n776 585
R349 B.n775 B.n774 585
R350 B.n773 B.n772 585
R351 B.n771 B.n770 585
R352 B.n769 B.n768 585
R353 B.n767 B.n766 585
R354 B.n765 B.n764 585
R355 B.n763 B.n762 585
R356 B.n761 B.n760 585
R357 B.n759 B.n758 585
R358 B.n757 B.n756 585
R359 B.n755 B.n754 585
R360 B.n753 B.n752 585
R361 B.n751 B.n750 585
R362 B.n749 B.n748 585
R363 B.n747 B.n746 585
R364 B.n745 B.n744 585
R365 B.n743 B.n742 585
R366 B.n741 B.n740 585
R367 B.n739 B.n738 585
R368 B.n737 B.n736 585
R369 B.n735 B.n734 585
R370 B.n733 B.n732 585
R371 B.n731 B.n730 585
R372 B.n729 B.n728 585
R373 B.n727 B.n726 585
R374 B.n725 B.n724 585
R375 B.n723 B.n722 585
R376 B.n721 B.n720 585
R377 B.n719 B.n718 585
R378 B.n717 B.n716 585
R379 B.n715 B.n714 585
R380 B.n713 B.n712 585
R381 B.n711 B.n710 585
R382 B.n709 B.n708 585
R383 B.n707 B.n706 585
R384 B.n705 B.n704 585
R385 B.n703 B.n702 585
R386 B.n701 B.n700 585
R387 B.n699 B.n698 585
R388 B.n697 B.n696 585
R389 B.n695 B.n694 585
R390 B.n693 B.n692 585
R391 B.n691 B.n690 585
R392 B.n689 B.n688 585
R393 B.n687 B.n686 585
R394 B.n685 B.n684 585
R395 B.n683 B.n682 585
R396 B.n681 B.n680 585
R397 B.n679 B.n678 585
R398 B.n677 B.n676 585
R399 B.n675 B.n674 585
R400 B.n673 B.n672 585
R401 B.n671 B.n670 585
R402 B.n669 B.n668 585
R403 B.n667 B.n666 585
R404 B.n665 B.n664 585
R405 B.n663 B.n662 585
R406 B.n661 B.n660 585
R407 B.n659 B.n658 585
R408 B.n657 B.n656 585
R409 B.n655 B.n654 585
R410 B.n653 B.n652 585
R411 B.n651 B.n650 585
R412 B.n649 B.n648 585
R413 B.n647 B.n646 585
R414 B.n645 B.n644 585
R415 B.n643 B.n642 585
R416 B.n641 B.n640 585
R417 B.n639 B.n638 585
R418 B.n637 B.n636 585
R419 B.n635 B.n634 585
R420 B.n633 B.n632 585
R421 B.n631 B.n630 585
R422 B.n629 B.n628 585
R423 B.n627 B.n626 585
R424 B.n625 B.n624 585
R425 B.n623 B.n622 585
R426 B.n621 B.n620 585
R427 B.n619 B.n618 585
R428 B.n617 B.n616 585
R429 B.n615 B.n614 585
R430 B.n613 B.n612 585
R431 B.n611 B.n610 585
R432 B.n609 B.n608 585
R433 B.n607 B.n606 585
R434 B.n605 B.n604 585
R435 B.n603 B.n602 585
R436 B.n601 B.n600 585
R437 B.n599 B.n598 585
R438 B.n597 B.n596 585
R439 B.n595 B.n594 585
R440 B.n593 B.n592 585
R441 B.n591 B.n590 585
R442 B.n589 B.n588 585
R443 B.n587 B.n586 585
R444 B.n585 B.n584 585
R445 B.n583 B.n582 585
R446 B.n581 B.n580 585
R447 B.n579 B.n578 585
R448 B.n577 B.n576 585
R449 B.n575 B.n574 585
R450 B.n573 B.n572 585
R451 B.n571 B.n570 585
R452 B.n569 B.n568 585
R453 B.n567 B.n566 585
R454 B.n565 B.n564 585
R455 B.n563 B.n562 585
R456 B.n561 B.n560 585
R457 B.n559 B.n558 585
R458 B.n557 B.n556 585
R459 B.n555 B.n554 585
R460 B.n553 B.n552 585
R461 B.n551 B.n550 585
R462 B.n549 B.n548 585
R463 B.n547 B.n546 585
R464 B.n545 B.n544 585
R465 B.n543 B.n542 585
R466 B.n465 B.n464 585
R467 B.n819 B.n818 585
R468 B.n818 B.n817 585
R469 B.n461 B.n460 585
R470 B.n462 B.n461 585
R471 B.n825 B.n824 585
R472 B.n824 B.n823 585
R473 B.n826 B.n459 585
R474 B.n459 B.n458 585
R475 B.n828 B.n827 585
R476 B.n829 B.n828 585
R477 B.n453 B.n452 585
R478 B.n454 B.n453 585
R479 B.n837 B.n836 585
R480 B.n836 B.n835 585
R481 B.n838 B.n451 585
R482 B.n451 B.n450 585
R483 B.n840 B.n839 585
R484 B.n841 B.n840 585
R485 B.n445 B.n444 585
R486 B.n446 B.n445 585
R487 B.n849 B.n848 585
R488 B.n848 B.n847 585
R489 B.n850 B.n443 585
R490 B.n443 B.n442 585
R491 B.n852 B.n851 585
R492 B.n853 B.n852 585
R493 B.n437 B.n436 585
R494 B.n438 B.n437 585
R495 B.n862 B.n861 585
R496 B.n861 B.n860 585
R497 B.n863 B.n435 585
R498 B.n859 B.n435 585
R499 B.n865 B.n864 585
R500 B.n866 B.n865 585
R501 B.n430 B.n429 585
R502 B.n431 B.n430 585
R503 B.n874 B.n873 585
R504 B.n873 B.n872 585
R505 B.n875 B.n428 585
R506 B.n428 B.n427 585
R507 B.n877 B.n876 585
R508 B.n878 B.n877 585
R509 B.n422 B.n421 585
R510 B.n423 B.n422 585
R511 B.n886 B.n885 585
R512 B.n885 B.n884 585
R513 B.n887 B.n420 585
R514 B.n420 B.n418 585
R515 B.n889 B.n888 585
R516 B.n890 B.n889 585
R517 B.n414 B.n413 585
R518 B.n419 B.n414 585
R519 B.n899 B.n898 585
R520 B.n898 B.n897 585
R521 B.n900 B.n412 585
R522 B.n412 B.n411 585
R523 B.n902 B.n901 585
R524 B.n903 B.n902 585
R525 B.n2 B.n0 585
R526 B.n4 B.n2 585
R527 B.n3 B.n1 585
R528 B.n1004 B.n3 585
R529 B.n1002 B.n1001 585
R530 B.n1003 B.n1002 585
R531 B.n1000 B.n9 585
R532 B.n9 B.n8 585
R533 B.n999 B.n998 585
R534 B.n998 B.n997 585
R535 B.n11 B.n10 585
R536 B.n996 B.n11 585
R537 B.n994 B.n993 585
R538 B.n995 B.n994 585
R539 B.n992 B.n16 585
R540 B.n16 B.n15 585
R541 B.n991 B.n990 585
R542 B.n990 B.n989 585
R543 B.n18 B.n17 585
R544 B.n988 B.n18 585
R545 B.n986 B.n985 585
R546 B.n987 B.n986 585
R547 B.n984 B.n23 585
R548 B.n23 B.n22 585
R549 B.n983 B.n982 585
R550 B.n982 B.n981 585
R551 B.n25 B.n24 585
R552 B.n980 B.n25 585
R553 B.n978 B.n977 585
R554 B.n979 B.n978 585
R555 B.n976 B.n29 585
R556 B.n32 B.n29 585
R557 B.n975 B.n974 585
R558 B.n974 B.n973 585
R559 B.n31 B.n30 585
R560 B.n972 B.n31 585
R561 B.n970 B.n969 585
R562 B.n971 B.n970 585
R563 B.n968 B.n37 585
R564 B.n37 B.n36 585
R565 B.n967 B.n966 585
R566 B.n966 B.n965 585
R567 B.n39 B.n38 585
R568 B.n964 B.n39 585
R569 B.n962 B.n961 585
R570 B.n963 B.n962 585
R571 B.n960 B.n44 585
R572 B.n44 B.n43 585
R573 B.n959 B.n958 585
R574 B.n958 B.n957 585
R575 B.n46 B.n45 585
R576 B.n956 B.n46 585
R577 B.n954 B.n953 585
R578 B.n955 B.n954 585
R579 B.n952 B.n51 585
R580 B.n51 B.n50 585
R581 B.n951 B.n950 585
R582 B.n950 B.n949 585
R583 B.n53 B.n52 585
R584 B.n948 B.n53 585
R585 B.n1007 B.n1006 585
R586 B.n1006 B.n1005 585
R587 B.n539 B.t10 532.399
R588 B.n536 B.t14 532.399
R589 B.n128 B.t17 532.399
R590 B.n126 B.t6 532.399
R591 B.n815 B.n461 511.721
R592 B.n130 B.n53 511.721
R593 B.n818 B.n463 511.721
R594 B.n945 B.n55 511.721
R595 B.n947 B.n946 256.663
R596 B.n947 B.n124 256.663
R597 B.n947 B.n123 256.663
R598 B.n947 B.n122 256.663
R599 B.n947 B.n121 256.663
R600 B.n947 B.n120 256.663
R601 B.n947 B.n119 256.663
R602 B.n947 B.n118 256.663
R603 B.n947 B.n117 256.663
R604 B.n947 B.n116 256.663
R605 B.n947 B.n115 256.663
R606 B.n947 B.n114 256.663
R607 B.n947 B.n113 256.663
R608 B.n947 B.n112 256.663
R609 B.n947 B.n111 256.663
R610 B.n947 B.n110 256.663
R611 B.n947 B.n109 256.663
R612 B.n947 B.n108 256.663
R613 B.n947 B.n107 256.663
R614 B.n947 B.n106 256.663
R615 B.n947 B.n105 256.663
R616 B.n947 B.n104 256.663
R617 B.n947 B.n103 256.663
R618 B.n947 B.n102 256.663
R619 B.n947 B.n101 256.663
R620 B.n947 B.n100 256.663
R621 B.n947 B.n99 256.663
R622 B.n947 B.n98 256.663
R623 B.n947 B.n97 256.663
R624 B.n947 B.n96 256.663
R625 B.n947 B.n95 256.663
R626 B.n947 B.n94 256.663
R627 B.n947 B.n93 256.663
R628 B.n947 B.n92 256.663
R629 B.n947 B.n91 256.663
R630 B.n947 B.n90 256.663
R631 B.n947 B.n89 256.663
R632 B.n947 B.n88 256.663
R633 B.n947 B.n87 256.663
R634 B.n947 B.n86 256.663
R635 B.n947 B.n85 256.663
R636 B.n947 B.n84 256.663
R637 B.n947 B.n83 256.663
R638 B.n947 B.n82 256.663
R639 B.n947 B.n81 256.663
R640 B.n947 B.n80 256.663
R641 B.n947 B.n79 256.663
R642 B.n947 B.n78 256.663
R643 B.n947 B.n77 256.663
R644 B.n947 B.n76 256.663
R645 B.n947 B.n75 256.663
R646 B.n947 B.n74 256.663
R647 B.n947 B.n73 256.663
R648 B.n947 B.n72 256.663
R649 B.n947 B.n71 256.663
R650 B.n947 B.n70 256.663
R651 B.n947 B.n69 256.663
R652 B.n947 B.n68 256.663
R653 B.n947 B.n67 256.663
R654 B.n947 B.n66 256.663
R655 B.n947 B.n65 256.663
R656 B.n947 B.n64 256.663
R657 B.n947 B.n63 256.663
R658 B.n947 B.n62 256.663
R659 B.n947 B.n61 256.663
R660 B.n947 B.n60 256.663
R661 B.n947 B.n59 256.663
R662 B.n947 B.n58 256.663
R663 B.n947 B.n57 256.663
R664 B.n947 B.n56 256.663
R665 B.n817 B.n816 256.663
R666 B.n817 B.n466 256.663
R667 B.n817 B.n467 256.663
R668 B.n817 B.n468 256.663
R669 B.n817 B.n469 256.663
R670 B.n817 B.n470 256.663
R671 B.n817 B.n471 256.663
R672 B.n817 B.n472 256.663
R673 B.n817 B.n473 256.663
R674 B.n817 B.n474 256.663
R675 B.n817 B.n475 256.663
R676 B.n817 B.n476 256.663
R677 B.n817 B.n477 256.663
R678 B.n817 B.n478 256.663
R679 B.n817 B.n479 256.663
R680 B.n817 B.n480 256.663
R681 B.n817 B.n481 256.663
R682 B.n817 B.n482 256.663
R683 B.n817 B.n483 256.663
R684 B.n817 B.n484 256.663
R685 B.n817 B.n485 256.663
R686 B.n817 B.n486 256.663
R687 B.n817 B.n487 256.663
R688 B.n817 B.n488 256.663
R689 B.n817 B.n489 256.663
R690 B.n817 B.n490 256.663
R691 B.n817 B.n491 256.663
R692 B.n817 B.n492 256.663
R693 B.n817 B.n493 256.663
R694 B.n817 B.n494 256.663
R695 B.n817 B.n495 256.663
R696 B.n817 B.n496 256.663
R697 B.n817 B.n497 256.663
R698 B.n817 B.n498 256.663
R699 B.n817 B.n499 256.663
R700 B.n817 B.n500 256.663
R701 B.n817 B.n501 256.663
R702 B.n817 B.n502 256.663
R703 B.n817 B.n503 256.663
R704 B.n817 B.n504 256.663
R705 B.n817 B.n505 256.663
R706 B.n817 B.n506 256.663
R707 B.n817 B.n507 256.663
R708 B.n817 B.n508 256.663
R709 B.n817 B.n509 256.663
R710 B.n817 B.n510 256.663
R711 B.n817 B.n511 256.663
R712 B.n817 B.n512 256.663
R713 B.n817 B.n513 256.663
R714 B.n817 B.n514 256.663
R715 B.n817 B.n515 256.663
R716 B.n817 B.n516 256.663
R717 B.n817 B.n517 256.663
R718 B.n817 B.n518 256.663
R719 B.n817 B.n519 256.663
R720 B.n817 B.n520 256.663
R721 B.n817 B.n521 256.663
R722 B.n817 B.n522 256.663
R723 B.n817 B.n523 256.663
R724 B.n817 B.n524 256.663
R725 B.n817 B.n525 256.663
R726 B.n817 B.n526 256.663
R727 B.n817 B.n527 256.663
R728 B.n817 B.n528 256.663
R729 B.n817 B.n529 256.663
R730 B.n817 B.n530 256.663
R731 B.n817 B.n531 256.663
R732 B.n817 B.n532 256.663
R733 B.n817 B.n533 256.663
R734 B.n824 B.n461 163.367
R735 B.n824 B.n459 163.367
R736 B.n828 B.n459 163.367
R737 B.n828 B.n453 163.367
R738 B.n836 B.n453 163.367
R739 B.n836 B.n451 163.367
R740 B.n840 B.n451 163.367
R741 B.n840 B.n445 163.367
R742 B.n848 B.n445 163.367
R743 B.n848 B.n443 163.367
R744 B.n852 B.n443 163.367
R745 B.n852 B.n437 163.367
R746 B.n861 B.n437 163.367
R747 B.n861 B.n435 163.367
R748 B.n865 B.n435 163.367
R749 B.n865 B.n430 163.367
R750 B.n873 B.n430 163.367
R751 B.n873 B.n428 163.367
R752 B.n877 B.n428 163.367
R753 B.n877 B.n422 163.367
R754 B.n885 B.n422 163.367
R755 B.n885 B.n420 163.367
R756 B.n889 B.n420 163.367
R757 B.n889 B.n414 163.367
R758 B.n898 B.n414 163.367
R759 B.n898 B.n412 163.367
R760 B.n902 B.n412 163.367
R761 B.n902 B.n2 163.367
R762 B.n1006 B.n2 163.367
R763 B.n1006 B.n3 163.367
R764 B.n1002 B.n3 163.367
R765 B.n1002 B.n9 163.367
R766 B.n998 B.n9 163.367
R767 B.n998 B.n11 163.367
R768 B.n994 B.n11 163.367
R769 B.n994 B.n16 163.367
R770 B.n990 B.n16 163.367
R771 B.n990 B.n18 163.367
R772 B.n986 B.n18 163.367
R773 B.n986 B.n23 163.367
R774 B.n982 B.n23 163.367
R775 B.n982 B.n25 163.367
R776 B.n978 B.n25 163.367
R777 B.n978 B.n29 163.367
R778 B.n974 B.n29 163.367
R779 B.n974 B.n31 163.367
R780 B.n970 B.n31 163.367
R781 B.n970 B.n37 163.367
R782 B.n966 B.n37 163.367
R783 B.n966 B.n39 163.367
R784 B.n962 B.n39 163.367
R785 B.n962 B.n44 163.367
R786 B.n958 B.n44 163.367
R787 B.n958 B.n46 163.367
R788 B.n954 B.n46 163.367
R789 B.n954 B.n51 163.367
R790 B.n950 B.n51 163.367
R791 B.n950 B.n53 163.367
R792 B.n535 B.n534 163.367
R793 B.n810 B.n534 163.367
R794 B.n808 B.n807 163.367
R795 B.n804 B.n803 163.367
R796 B.n800 B.n799 163.367
R797 B.n796 B.n795 163.367
R798 B.n792 B.n791 163.367
R799 B.n788 B.n787 163.367
R800 B.n784 B.n783 163.367
R801 B.n780 B.n779 163.367
R802 B.n776 B.n775 163.367
R803 B.n772 B.n771 163.367
R804 B.n768 B.n767 163.367
R805 B.n764 B.n763 163.367
R806 B.n760 B.n759 163.367
R807 B.n756 B.n755 163.367
R808 B.n752 B.n751 163.367
R809 B.n748 B.n747 163.367
R810 B.n744 B.n743 163.367
R811 B.n740 B.n739 163.367
R812 B.n736 B.n735 163.367
R813 B.n732 B.n731 163.367
R814 B.n728 B.n727 163.367
R815 B.n724 B.n723 163.367
R816 B.n720 B.n719 163.367
R817 B.n716 B.n715 163.367
R818 B.n712 B.n711 163.367
R819 B.n708 B.n707 163.367
R820 B.n704 B.n703 163.367
R821 B.n700 B.n699 163.367
R822 B.n696 B.n695 163.367
R823 B.n692 B.n691 163.367
R824 B.n688 B.n687 163.367
R825 B.n684 B.n683 163.367
R826 B.n680 B.n679 163.367
R827 B.n676 B.n675 163.367
R828 B.n672 B.n671 163.367
R829 B.n668 B.n667 163.367
R830 B.n664 B.n663 163.367
R831 B.n660 B.n659 163.367
R832 B.n656 B.n655 163.367
R833 B.n652 B.n651 163.367
R834 B.n648 B.n647 163.367
R835 B.n644 B.n643 163.367
R836 B.n640 B.n639 163.367
R837 B.n636 B.n635 163.367
R838 B.n632 B.n631 163.367
R839 B.n628 B.n627 163.367
R840 B.n624 B.n623 163.367
R841 B.n620 B.n619 163.367
R842 B.n616 B.n615 163.367
R843 B.n612 B.n611 163.367
R844 B.n608 B.n607 163.367
R845 B.n604 B.n603 163.367
R846 B.n600 B.n599 163.367
R847 B.n596 B.n595 163.367
R848 B.n592 B.n591 163.367
R849 B.n588 B.n587 163.367
R850 B.n584 B.n583 163.367
R851 B.n580 B.n579 163.367
R852 B.n576 B.n575 163.367
R853 B.n572 B.n571 163.367
R854 B.n568 B.n567 163.367
R855 B.n564 B.n563 163.367
R856 B.n560 B.n559 163.367
R857 B.n556 B.n555 163.367
R858 B.n552 B.n551 163.367
R859 B.n548 B.n547 163.367
R860 B.n544 B.n543 163.367
R861 B.n818 B.n465 163.367
R862 B.n822 B.n463 163.367
R863 B.n822 B.n457 163.367
R864 B.n830 B.n457 163.367
R865 B.n830 B.n455 163.367
R866 B.n834 B.n455 163.367
R867 B.n834 B.n449 163.367
R868 B.n842 B.n449 163.367
R869 B.n842 B.n447 163.367
R870 B.n846 B.n447 163.367
R871 B.n846 B.n441 163.367
R872 B.n854 B.n441 163.367
R873 B.n854 B.n439 163.367
R874 B.n858 B.n439 163.367
R875 B.n858 B.n434 163.367
R876 B.n867 B.n434 163.367
R877 B.n867 B.n432 163.367
R878 B.n871 B.n432 163.367
R879 B.n871 B.n426 163.367
R880 B.n879 B.n426 163.367
R881 B.n879 B.n424 163.367
R882 B.n883 B.n424 163.367
R883 B.n883 B.n417 163.367
R884 B.n891 B.n417 163.367
R885 B.n891 B.n415 163.367
R886 B.n896 B.n415 163.367
R887 B.n896 B.n410 163.367
R888 B.n904 B.n410 163.367
R889 B.n905 B.n904 163.367
R890 B.n905 B.n5 163.367
R891 B.n6 B.n5 163.367
R892 B.n7 B.n6 163.367
R893 B.n910 B.n7 163.367
R894 B.n910 B.n12 163.367
R895 B.n13 B.n12 163.367
R896 B.n14 B.n13 163.367
R897 B.n915 B.n14 163.367
R898 B.n915 B.n19 163.367
R899 B.n20 B.n19 163.367
R900 B.n21 B.n20 163.367
R901 B.n920 B.n21 163.367
R902 B.n920 B.n26 163.367
R903 B.n27 B.n26 163.367
R904 B.n28 B.n27 163.367
R905 B.n925 B.n28 163.367
R906 B.n925 B.n33 163.367
R907 B.n34 B.n33 163.367
R908 B.n35 B.n34 163.367
R909 B.n930 B.n35 163.367
R910 B.n930 B.n40 163.367
R911 B.n41 B.n40 163.367
R912 B.n42 B.n41 163.367
R913 B.n935 B.n42 163.367
R914 B.n935 B.n47 163.367
R915 B.n48 B.n47 163.367
R916 B.n49 B.n48 163.367
R917 B.n940 B.n49 163.367
R918 B.n940 B.n54 163.367
R919 B.n55 B.n54 163.367
R920 B.n134 B.n133 163.367
R921 B.n138 B.n137 163.367
R922 B.n142 B.n141 163.367
R923 B.n146 B.n145 163.367
R924 B.n150 B.n149 163.367
R925 B.n154 B.n153 163.367
R926 B.n158 B.n157 163.367
R927 B.n162 B.n161 163.367
R928 B.n166 B.n165 163.367
R929 B.n170 B.n169 163.367
R930 B.n174 B.n173 163.367
R931 B.n178 B.n177 163.367
R932 B.n182 B.n181 163.367
R933 B.n186 B.n185 163.367
R934 B.n190 B.n189 163.367
R935 B.n194 B.n193 163.367
R936 B.n198 B.n197 163.367
R937 B.n202 B.n201 163.367
R938 B.n206 B.n205 163.367
R939 B.n210 B.n209 163.367
R940 B.n214 B.n213 163.367
R941 B.n218 B.n217 163.367
R942 B.n222 B.n221 163.367
R943 B.n226 B.n225 163.367
R944 B.n230 B.n229 163.367
R945 B.n234 B.n233 163.367
R946 B.n238 B.n237 163.367
R947 B.n242 B.n241 163.367
R948 B.n246 B.n245 163.367
R949 B.n250 B.n249 163.367
R950 B.n254 B.n253 163.367
R951 B.n258 B.n257 163.367
R952 B.n263 B.n262 163.367
R953 B.n267 B.n266 163.367
R954 B.n271 B.n270 163.367
R955 B.n275 B.n274 163.367
R956 B.n279 B.n278 163.367
R957 B.n284 B.n283 163.367
R958 B.n288 B.n287 163.367
R959 B.n292 B.n291 163.367
R960 B.n296 B.n295 163.367
R961 B.n300 B.n299 163.367
R962 B.n304 B.n303 163.367
R963 B.n308 B.n307 163.367
R964 B.n312 B.n311 163.367
R965 B.n316 B.n315 163.367
R966 B.n320 B.n319 163.367
R967 B.n324 B.n323 163.367
R968 B.n328 B.n327 163.367
R969 B.n332 B.n331 163.367
R970 B.n336 B.n335 163.367
R971 B.n340 B.n339 163.367
R972 B.n344 B.n343 163.367
R973 B.n348 B.n347 163.367
R974 B.n352 B.n351 163.367
R975 B.n356 B.n355 163.367
R976 B.n360 B.n359 163.367
R977 B.n364 B.n363 163.367
R978 B.n368 B.n367 163.367
R979 B.n372 B.n371 163.367
R980 B.n376 B.n375 163.367
R981 B.n380 B.n379 163.367
R982 B.n384 B.n383 163.367
R983 B.n388 B.n387 163.367
R984 B.n392 B.n391 163.367
R985 B.n396 B.n395 163.367
R986 B.n400 B.n399 163.367
R987 B.n404 B.n403 163.367
R988 B.n406 B.n125 163.367
R989 B.n539 B.t13 106.513
R990 B.n126 B.t8 106.513
R991 B.n536 B.t16 106.487
R992 B.n128 B.t18 106.487
R993 B.n816 B.n815 71.676
R994 B.n810 B.n466 71.676
R995 B.n807 B.n467 71.676
R996 B.n803 B.n468 71.676
R997 B.n799 B.n469 71.676
R998 B.n795 B.n470 71.676
R999 B.n791 B.n471 71.676
R1000 B.n787 B.n472 71.676
R1001 B.n783 B.n473 71.676
R1002 B.n779 B.n474 71.676
R1003 B.n775 B.n475 71.676
R1004 B.n771 B.n476 71.676
R1005 B.n767 B.n477 71.676
R1006 B.n763 B.n478 71.676
R1007 B.n759 B.n479 71.676
R1008 B.n755 B.n480 71.676
R1009 B.n751 B.n481 71.676
R1010 B.n747 B.n482 71.676
R1011 B.n743 B.n483 71.676
R1012 B.n739 B.n484 71.676
R1013 B.n735 B.n485 71.676
R1014 B.n731 B.n486 71.676
R1015 B.n727 B.n487 71.676
R1016 B.n723 B.n488 71.676
R1017 B.n719 B.n489 71.676
R1018 B.n715 B.n490 71.676
R1019 B.n711 B.n491 71.676
R1020 B.n707 B.n492 71.676
R1021 B.n703 B.n493 71.676
R1022 B.n699 B.n494 71.676
R1023 B.n695 B.n495 71.676
R1024 B.n691 B.n496 71.676
R1025 B.n687 B.n497 71.676
R1026 B.n683 B.n498 71.676
R1027 B.n679 B.n499 71.676
R1028 B.n675 B.n500 71.676
R1029 B.n671 B.n501 71.676
R1030 B.n667 B.n502 71.676
R1031 B.n663 B.n503 71.676
R1032 B.n659 B.n504 71.676
R1033 B.n655 B.n505 71.676
R1034 B.n651 B.n506 71.676
R1035 B.n647 B.n507 71.676
R1036 B.n643 B.n508 71.676
R1037 B.n639 B.n509 71.676
R1038 B.n635 B.n510 71.676
R1039 B.n631 B.n511 71.676
R1040 B.n627 B.n512 71.676
R1041 B.n623 B.n513 71.676
R1042 B.n619 B.n514 71.676
R1043 B.n615 B.n515 71.676
R1044 B.n611 B.n516 71.676
R1045 B.n607 B.n517 71.676
R1046 B.n603 B.n518 71.676
R1047 B.n599 B.n519 71.676
R1048 B.n595 B.n520 71.676
R1049 B.n591 B.n521 71.676
R1050 B.n587 B.n522 71.676
R1051 B.n583 B.n523 71.676
R1052 B.n579 B.n524 71.676
R1053 B.n575 B.n525 71.676
R1054 B.n571 B.n526 71.676
R1055 B.n567 B.n527 71.676
R1056 B.n563 B.n528 71.676
R1057 B.n559 B.n529 71.676
R1058 B.n555 B.n530 71.676
R1059 B.n551 B.n531 71.676
R1060 B.n547 B.n532 71.676
R1061 B.n543 B.n533 71.676
R1062 B.n130 B.n56 71.676
R1063 B.n134 B.n57 71.676
R1064 B.n138 B.n58 71.676
R1065 B.n142 B.n59 71.676
R1066 B.n146 B.n60 71.676
R1067 B.n150 B.n61 71.676
R1068 B.n154 B.n62 71.676
R1069 B.n158 B.n63 71.676
R1070 B.n162 B.n64 71.676
R1071 B.n166 B.n65 71.676
R1072 B.n170 B.n66 71.676
R1073 B.n174 B.n67 71.676
R1074 B.n178 B.n68 71.676
R1075 B.n182 B.n69 71.676
R1076 B.n186 B.n70 71.676
R1077 B.n190 B.n71 71.676
R1078 B.n194 B.n72 71.676
R1079 B.n198 B.n73 71.676
R1080 B.n202 B.n74 71.676
R1081 B.n206 B.n75 71.676
R1082 B.n210 B.n76 71.676
R1083 B.n214 B.n77 71.676
R1084 B.n218 B.n78 71.676
R1085 B.n222 B.n79 71.676
R1086 B.n226 B.n80 71.676
R1087 B.n230 B.n81 71.676
R1088 B.n234 B.n82 71.676
R1089 B.n238 B.n83 71.676
R1090 B.n242 B.n84 71.676
R1091 B.n246 B.n85 71.676
R1092 B.n250 B.n86 71.676
R1093 B.n254 B.n87 71.676
R1094 B.n258 B.n88 71.676
R1095 B.n263 B.n89 71.676
R1096 B.n267 B.n90 71.676
R1097 B.n271 B.n91 71.676
R1098 B.n275 B.n92 71.676
R1099 B.n279 B.n93 71.676
R1100 B.n284 B.n94 71.676
R1101 B.n288 B.n95 71.676
R1102 B.n292 B.n96 71.676
R1103 B.n296 B.n97 71.676
R1104 B.n300 B.n98 71.676
R1105 B.n304 B.n99 71.676
R1106 B.n308 B.n100 71.676
R1107 B.n312 B.n101 71.676
R1108 B.n316 B.n102 71.676
R1109 B.n320 B.n103 71.676
R1110 B.n324 B.n104 71.676
R1111 B.n328 B.n105 71.676
R1112 B.n332 B.n106 71.676
R1113 B.n336 B.n107 71.676
R1114 B.n340 B.n108 71.676
R1115 B.n344 B.n109 71.676
R1116 B.n348 B.n110 71.676
R1117 B.n352 B.n111 71.676
R1118 B.n356 B.n112 71.676
R1119 B.n360 B.n113 71.676
R1120 B.n364 B.n114 71.676
R1121 B.n368 B.n115 71.676
R1122 B.n372 B.n116 71.676
R1123 B.n376 B.n117 71.676
R1124 B.n380 B.n118 71.676
R1125 B.n384 B.n119 71.676
R1126 B.n388 B.n120 71.676
R1127 B.n392 B.n121 71.676
R1128 B.n396 B.n122 71.676
R1129 B.n400 B.n123 71.676
R1130 B.n404 B.n124 71.676
R1131 B.n946 B.n125 71.676
R1132 B.n946 B.n945 71.676
R1133 B.n406 B.n124 71.676
R1134 B.n403 B.n123 71.676
R1135 B.n399 B.n122 71.676
R1136 B.n395 B.n121 71.676
R1137 B.n391 B.n120 71.676
R1138 B.n387 B.n119 71.676
R1139 B.n383 B.n118 71.676
R1140 B.n379 B.n117 71.676
R1141 B.n375 B.n116 71.676
R1142 B.n371 B.n115 71.676
R1143 B.n367 B.n114 71.676
R1144 B.n363 B.n113 71.676
R1145 B.n359 B.n112 71.676
R1146 B.n355 B.n111 71.676
R1147 B.n351 B.n110 71.676
R1148 B.n347 B.n109 71.676
R1149 B.n343 B.n108 71.676
R1150 B.n339 B.n107 71.676
R1151 B.n335 B.n106 71.676
R1152 B.n331 B.n105 71.676
R1153 B.n327 B.n104 71.676
R1154 B.n323 B.n103 71.676
R1155 B.n319 B.n102 71.676
R1156 B.n315 B.n101 71.676
R1157 B.n311 B.n100 71.676
R1158 B.n307 B.n99 71.676
R1159 B.n303 B.n98 71.676
R1160 B.n299 B.n97 71.676
R1161 B.n295 B.n96 71.676
R1162 B.n291 B.n95 71.676
R1163 B.n287 B.n94 71.676
R1164 B.n283 B.n93 71.676
R1165 B.n278 B.n92 71.676
R1166 B.n274 B.n91 71.676
R1167 B.n270 B.n90 71.676
R1168 B.n266 B.n89 71.676
R1169 B.n262 B.n88 71.676
R1170 B.n257 B.n87 71.676
R1171 B.n253 B.n86 71.676
R1172 B.n249 B.n85 71.676
R1173 B.n245 B.n84 71.676
R1174 B.n241 B.n83 71.676
R1175 B.n237 B.n82 71.676
R1176 B.n233 B.n81 71.676
R1177 B.n229 B.n80 71.676
R1178 B.n225 B.n79 71.676
R1179 B.n221 B.n78 71.676
R1180 B.n217 B.n77 71.676
R1181 B.n213 B.n76 71.676
R1182 B.n209 B.n75 71.676
R1183 B.n205 B.n74 71.676
R1184 B.n201 B.n73 71.676
R1185 B.n197 B.n72 71.676
R1186 B.n193 B.n71 71.676
R1187 B.n189 B.n70 71.676
R1188 B.n185 B.n69 71.676
R1189 B.n181 B.n68 71.676
R1190 B.n177 B.n67 71.676
R1191 B.n173 B.n66 71.676
R1192 B.n169 B.n65 71.676
R1193 B.n165 B.n64 71.676
R1194 B.n161 B.n63 71.676
R1195 B.n157 B.n62 71.676
R1196 B.n153 B.n61 71.676
R1197 B.n149 B.n60 71.676
R1198 B.n145 B.n59 71.676
R1199 B.n141 B.n58 71.676
R1200 B.n137 B.n57 71.676
R1201 B.n133 B.n56 71.676
R1202 B.n816 B.n535 71.676
R1203 B.n808 B.n466 71.676
R1204 B.n804 B.n467 71.676
R1205 B.n800 B.n468 71.676
R1206 B.n796 B.n469 71.676
R1207 B.n792 B.n470 71.676
R1208 B.n788 B.n471 71.676
R1209 B.n784 B.n472 71.676
R1210 B.n780 B.n473 71.676
R1211 B.n776 B.n474 71.676
R1212 B.n772 B.n475 71.676
R1213 B.n768 B.n476 71.676
R1214 B.n764 B.n477 71.676
R1215 B.n760 B.n478 71.676
R1216 B.n756 B.n479 71.676
R1217 B.n752 B.n480 71.676
R1218 B.n748 B.n481 71.676
R1219 B.n744 B.n482 71.676
R1220 B.n740 B.n483 71.676
R1221 B.n736 B.n484 71.676
R1222 B.n732 B.n485 71.676
R1223 B.n728 B.n486 71.676
R1224 B.n724 B.n487 71.676
R1225 B.n720 B.n488 71.676
R1226 B.n716 B.n489 71.676
R1227 B.n712 B.n490 71.676
R1228 B.n708 B.n491 71.676
R1229 B.n704 B.n492 71.676
R1230 B.n700 B.n493 71.676
R1231 B.n696 B.n494 71.676
R1232 B.n692 B.n495 71.676
R1233 B.n688 B.n496 71.676
R1234 B.n684 B.n497 71.676
R1235 B.n680 B.n498 71.676
R1236 B.n676 B.n499 71.676
R1237 B.n672 B.n500 71.676
R1238 B.n668 B.n501 71.676
R1239 B.n664 B.n502 71.676
R1240 B.n660 B.n503 71.676
R1241 B.n656 B.n504 71.676
R1242 B.n652 B.n505 71.676
R1243 B.n648 B.n506 71.676
R1244 B.n644 B.n507 71.676
R1245 B.n640 B.n508 71.676
R1246 B.n636 B.n509 71.676
R1247 B.n632 B.n510 71.676
R1248 B.n628 B.n511 71.676
R1249 B.n624 B.n512 71.676
R1250 B.n620 B.n513 71.676
R1251 B.n616 B.n514 71.676
R1252 B.n612 B.n515 71.676
R1253 B.n608 B.n516 71.676
R1254 B.n604 B.n517 71.676
R1255 B.n600 B.n518 71.676
R1256 B.n596 B.n519 71.676
R1257 B.n592 B.n520 71.676
R1258 B.n588 B.n521 71.676
R1259 B.n584 B.n522 71.676
R1260 B.n580 B.n523 71.676
R1261 B.n576 B.n524 71.676
R1262 B.n572 B.n525 71.676
R1263 B.n568 B.n526 71.676
R1264 B.n564 B.n527 71.676
R1265 B.n560 B.n528 71.676
R1266 B.n556 B.n529 71.676
R1267 B.n552 B.n530 71.676
R1268 B.n548 B.n531 71.676
R1269 B.n544 B.n532 71.676
R1270 B.n533 B.n465 71.676
R1271 B.n540 B.t12 71.6045
R1272 B.n127 B.t9 71.6045
R1273 B.n537 B.t15 71.5777
R1274 B.n129 B.t19 71.5777
R1275 B.n817 B.n462 62.3593
R1276 B.n948 B.n947 62.3593
R1277 B.n541 B.n540 59.5399
R1278 B.n538 B.n537 59.5399
R1279 B.n260 B.n129 59.5399
R1280 B.n281 B.n127 59.5399
R1281 B.n540 B.n539 34.9096
R1282 B.n537 B.n536 34.9096
R1283 B.n129 B.n128 34.9096
R1284 B.n127 B.n126 34.9096
R1285 B.n131 B.n52 33.2493
R1286 B.n944 B.n943 33.2493
R1287 B.n820 B.n819 33.2493
R1288 B.n814 B.n460 33.2493
R1289 B.n823 B.n462 29.6536
R1290 B.n823 B.n458 29.6536
R1291 B.n829 B.n458 29.6536
R1292 B.n829 B.n454 29.6536
R1293 B.n835 B.n454 29.6536
R1294 B.n841 B.n450 29.6536
R1295 B.n841 B.n446 29.6536
R1296 B.n847 B.n446 29.6536
R1297 B.n847 B.n442 29.6536
R1298 B.n853 B.n442 29.6536
R1299 B.n853 B.n438 29.6536
R1300 B.n860 B.n438 29.6536
R1301 B.n860 B.n859 29.6536
R1302 B.n866 B.n431 29.6536
R1303 B.n872 B.n431 29.6536
R1304 B.n872 B.n427 29.6536
R1305 B.n878 B.n427 29.6536
R1306 B.n884 B.n423 29.6536
R1307 B.n884 B.n418 29.6536
R1308 B.n890 B.n418 29.6536
R1309 B.n890 B.n419 29.6536
R1310 B.n897 B.n411 29.6536
R1311 B.n903 B.n411 29.6536
R1312 B.n903 B.n4 29.6536
R1313 B.n1005 B.n4 29.6536
R1314 B.n1005 B.n1004 29.6536
R1315 B.n1004 B.n1003 29.6536
R1316 B.n1003 B.n8 29.6536
R1317 B.n997 B.n8 29.6536
R1318 B.n996 B.n995 29.6536
R1319 B.n995 B.n15 29.6536
R1320 B.n989 B.n15 29.6536
R1321 B.n989 B.n988 29.6536
R1322 B.n987 B.n22 29.6536
R1323 B.n981 B.n22 29.6536
R1324 B.n981 B.n980 29.6536
R1325 B.n980 B.n979 29.6536
R1326 B.n973 B.n32 29.6536
R1327 B.n973 B.n972 29.6536
R1328 B.n972 B.n971 29.6536
R1329 B.n971 B.n36 29.6536
R1330 B.n965 B.n36 29.6536
R1331 B.n965 B.n964 29.6536
R1332 B.n964 B.n963 29.6536
R1333 B.n963 B.n43 29.6536
R1334 B.n957 B.n956 29.6536
R1335 B.n956 B.n955 29.6536
R1336 B.n955 B.n50 29.6536
R1337 B.n949 B.n50 29.6536
R1338 B.n949 B.n948 29.6536
R1339 B.n866 B.t2 24.8568
R1340 B.n979 B.t4 24.8568
R1341 B.n419 B.t0 22.2403
R1342 B.t1 B.n996 22.2403
R1343 B.n835 B.t11 19.6239
R1344 B.n957 B.t7 19.6239
R1345 B B.n1007 18.0485
R1346 B.t3 B.n423 16.1353
R1347 B.n988 B.t5 16.1353
R1348 B.n878 B.t3 13.5188
R1349 B.t5 B.n987 13.5188
R1350 B.n132 B.n131 10.6151
R1351 B.n135 B.n132 10.6151
R1352 B.n136 B.n135 10.6151
R1353 B.n139 B.n136 10.6151
R1354 B.n140 B.n139 10.6151
R1355 B.n143 B.n140 10.6151
R1356 B.n144 B.n143 10.6151
R1357 B.n147 B.n144 10.6151
R1358 B.n148 B.n147 10.6151
R1359 B.n151 B.n148 10.6151
R1360 B.n152 B.n151 10.6151
R1361 B.n155 B.n152 10.6151
R1362 B.n156 B.n155 10.6151
R1363 B.n159 B.n156 10.6151
R1364 B.n160 B.n159 10.6151
R1365 B.n163 B.n160 10.6151
R1366 B.n164 B.n163 10.6151
R1367 B.n167 B.n164 10.6151
R1368 B.n168 B.n167 10.6151
R1369 B.n171 B.n168 10.6151
R1370 B.n172 B.n171 10.6151
R1371 B.n175 B.n172 10.6151
R1372 B.n176 B.n175 10.6151
R1373 B.n179 B.n176 10.6151
R1374 B.n180 B.n179 10.6151
R1375 B.n183 B.n180 10.6151
R1376 B.n184 B.n183 10.6151
R1377 B.n187 B.n184 10.6151
R1378 B.n188 B.n187 10.6151
R1379 B.n191 B.n188 10.6151
R1380 B.n192 B.n191 10.6151
R1381 B.n195 B.n192 10.6151
R1382 B.n196 B.n195 10.6151
R1383 B.n199 B.n196 10.6151
R1384 B.n200 B.n199 10.6151
R1385 B.n203 B.n200 10.6151
R1386 B.n204 B.n203 10.6151
R1387 B.n207 B.n204 10.6151
R1388 B.n208 B.n207 10.6151
R1389 B.n211 B.n208 10.6151
R1390 B.n212 B.n211 10.6151
R1391 B.n215 B.n212 10.6151
R1392 B.n216 B.n215 10.6151
R1393 B.n219 B.n216 10.6151
R1394 B.n220 B.n219 10.6151
R1395 B.n223 B.n220 10.6151
R1396 B.n224 B.n223 10.6151
R1397 B.n227 B.n224 10.6151
R1398 B.n228 B.n227 10.6151
R1399 B.n231 B.n228 10.6151
R1400 B.n232 B.n231 10.6151
R1401 B.n235 B.n232 10.6151
R1402 B.n236 B.n235 10.6151
R1403 B.n239 B.n236 10.6151
R1404 B.n240 B.n239 10.6151
R1405 B.n243 B.n240 10.6151
R1406 B.n244 B.n243 10.6151
R1407 B.n247 B.n244 10.6151
R1408 B.n248 B.n247 10.6151
R1409 B.n251 B.n248 10.6151
R1410 B.n252 B.n251 10.6151
R1411 B.n255 B.n252 10.6151
R1412 B.n256 B.n255 10.6151
R1413 B.n259 B.n256 10.6151
R1414 B.n264 B.n261 10.6151
R1415 B.n265 B.n264 10.6151
R1416 B.n268 B.n265 10.6151
R1417 B.n269 B.n268 10.6151
R1418 B.n272 B.n269 10.6151
R1419 B.n273 B.n272 10.6151
R1420 B.n276 B.n273 10.6151
R1421 B.n277 B.n276 10.6151
R1422 B.n280 B.n277 10.6151
R1423 B.n285 B.n282 10.6151
R1424 B.n286 B.n285 10.6151
R1425 B.n289 B.n286 10.6151
R1426 B.n290 B.n289 10.6151
R1427 B.n293 B.n290 10.6151
R1428 B.n294 B.n293 10.6151
R1429 B.n297 B.n294 10.6151
R1430 B.n298 B.n297 10.6151
R1431 B.n301 B.n298 10.6151
R1432 B.n302 B.n301 10.6151
R1433 B.n305 B.n302 10.6151
R1434 B.n306 B.n305 10.6151
R1435 B.n309 B.n306 10.6151
R1436 B.n310 B.n309 10.6151
R1437 B.n313 B.n310 10.6151
R1438 B.n314 B.n313 10.6151
R1439 B.n317 B.n314 10.6151
R1440 B.n318 B.n317 10.6151
R1441 B.n321 B.n318 10.6151
R1442 B.n322 B.n321 10.6151
R1443 B.n325 B.n322 10.6151
R1444 B.n326 B.n325 10.6151
R1445 B.n329 B.n326 10.6151
R1446 B.n330 B.n329 10.6151
R1447 B.n333 B.n330 10.6151
R1448 B.n334 B.n333 10.6151
R1449 B.n337 B.n334 10.6151
R1450 B.n338 B.n337 10.6151
R1451 B.n341 B.n338 10.6151
R1452 B.n342 B.n341 10.6151
R1453 B.n345 B.n342 10.6151
R1454 B.n346 B.n345 10.6151
R1455 B.n349 B.n346 10.6151
R1456 B.n350 B.n349 10.6151
R1457 B.n353 B.n350 10.6151
R1458 B.n354 B.n353 10.6151
R1459 B.n357 B.n354 10.6151
R1460 B.n358 B.n357 10.6151
R1461 B.n361 B.n358 10.6151
R1462 B.n362 B.n361 10.6151
R1463 B.n365 B.n362 10.6151
R1464 B.n366 B.n365 10.6151
R1465 B.n369 B.n366 10.6151
R1466 B.n370 B.n369 10.6151
R1467 B.n373 B.n370 10.6151
R1468 B.n374 B.n373 10.6151
R1469 B.n377 B.n374 10.6151
R1470 B.n378 B.n377 10.6151
R1471 B.n381 B.n378 10.6151
R1472 B.n382 B.n381 10.6151
R1473 B.n385 B.n382 10.6151
R1474 B.n386 B.n385 10.6151
R1475 B.n389 B.n386 10.6151
R1476 B.n390 B.n389 10.6151
R1477 B.n393 B.n390 10.6151
R1478 B.n394 B.n393 10.6151
R1479 B.n397 B.n394 10.6151
R1480 B.n398 B.n397 10.6151
R1481 B.n401 B.n398 10.6151
R1482 B.n402 B.n401 10.6151
R1483 B.n405 B.n402 10.6151
R1484 B.n407 B.n405 10.6151
R1485 B.n408 B.n407 10.6151
R1486 B.n944 B.n408 10.6151
R1487 B.n821 B.n820 10.6151
R1488 B.n821 B.n456 10.6151
R1489 B.n831 B.n456 10.6151
R1490 B.n832 B.n831 10.6151
R1491 B.n833 B.n832 10.6151
R1492 B.n833 B.n448 10.6151
R1493 B.n843 B.n448 10.6151
R1494 B.n844 B.n843 10.6151
R1495 B.n845 B.n844 10.6151
R1496 B.n845 B.n440 10.6151
R1497 B.n855 B.n440 10.6151
R1498 B.n856 B.n855 10.6151
R1499 B.n857 B.n856 10.6151
R1500 B.n857 B.n433 10.6151
R1501 B.n868 B.n433 10.6151
R1502 B.n869 B.n868 10.6151
R1503 B.n870 B.n869 10.6151
R1504 B.n870 B.n425 10.6151
R1505 B.n880 B.n425 10.6151
R1506 B.n881 B.n880 10.6151
R1507 B.n882 B.n881 10.6151
R1508 B.n882 B.n416 10.6151
R1509 B.n892 B.n416 10.6151
R1510 B.n893 B.n892 10.6151
R1511 B.n895 B.n893 10.6151
R1512 B.n895 B.n894 10.6151
R1513 B.n894 B.n409 10.6151
R1514 B.n906 B.n409 10.6151
R1515 B.n907 B.n906 10.6151
R1516 B.n908 B.n907 10.6151
R1517 B.n909 B.n908 10.6151
R1518 B.n911 B.n909 10.6151
R1519 B.n912 B.n911 10.6151
R1520 B.n913 B.n912 10.6151
R1521 B.n914 B.n913 10.6151
R1522 B.n916 B.n914 10.6151
R1523 B.n917 B.n916 10.6151
R1524 B.n918 B.n917 10.6151
R1525 B.n919 B.n918 10.6151
R1526 B.n921 B.n919 10.6151
R1527 B.n922 B.n921 10.6151
R1528 B.n923 B.n922 10.6151
R1529 B.n924 B.n923 10.6151
R1530 B.n926 B.n924 10.6151
R1531 B.n927 B.n926 10.6151
R1532 B.n928 B.n927 10.6151
R1533 B.n929 B.n928 10.6151
R1534 B.n931 B.n929 10.6151
R1535 B.n932 B.n931 10.6151
R1536 B.n933 B.n932 10.6151
R1537 B.n934 B.n933 10.6151
R1538 B.n936 B.n934 10.6151
R1539 B.n937 B.n936 10.6151
R1540 B.n938 B.n937 10.6151
R1541 B.n939 B.n938 10.6151
R1542 B.n941 B.n939 10.6151
R1543 B.n942 B.n941 10.6151
R1544 B.n943 B.n942 10.6151
R1545 B.n814 B.n813 10.6151
R1546 B.n813 B.n812 10.6151
R1547 B.n812 B.n811 10.6151
R1548 B.n811 B.n809 10.6151
R1549 B.n809 B.n806 10.6151
R1550 B.n806 B.n805 10.6151
R1551 B.n805 B.n802 10.6151
R1552 B.n802 B.n801 10.6151
R1553 B.n801 B.n798 10.6151
R1554 B.n798 B.n797 10.6151
R1555 B.n797 B.n794 10.6151
R1556 B.n794 B.n793 10.6151
R1557 B.n793 B.n790 10.6151
R1558 B.n790 B.n789 10.6151
R1559 B.n789 B.n786 10.6151
R1560 B.n786 B.n785 10.6151
R1561 B.n785 B.n782 10.6151
R1562 B.n782 B.n781 10.6151
R1563 B.n781 B.n778 10.6151
R1564 B.n778 B.n777 10.6151
R1565 B.n777 B.n774 10.6151
R1566 B.n774 B.n773 10.6151
R1567 B.n773 B.n770 10.6151
R1568 B.n770 B.n769 10.6151
R1569 B.n769 B.n766 10.6151
R1570 B.n766 B.n765 10.6151
R1571 B.n765 B.n762 10.6151
R1572 B.n762 B.n761 10.6151
R1573 B.n761 B.n758 10.6151
R1574 B.n758 B.n757 10.6151
R1575 B.n757 B.n754 10.6151
R1576 B.n754 B.n753 10.6151
R1577 B.n753 B.n750 10.6151
R1578 B.n750 B.n749 10.6151
R1579 B.n749 B.n746 10.6151
R1580 B.n746 B.n745 10.6151
R1581 B.n745 B.n742 10.6151
R1582 B.n742 B.n741 10.6151
R1583 B.n741 B.n738 10.6151
R1584 B.n738 B.n737 10.6151
R1585 B.n737 B.n734 10.6151
R1586 B.n734 B.n733 10.6151
R1587 B.n733 B.n730 10.6151
R1588 B.n730 B.n729 10.6151
R1589 B.n729 B.n726 10.6151
R1590 B.n726 B.n725 10.6151
R1591 B.n725 B.n722 10.6151
R1592 B.n722 B.n721 10.6151
R1593 B.n721 B.n718 10.6151
R1594 B.n718 B.n717 10.6151
R1595 B.n717 B.n714 10.6151
R1596 B.n714 B.n713 10.6151
R1597 B.n713 B.n710 10.6151
R1598 B.n710 B.n709 10.6151
R1599 B.n709 B.n706 10.6151
R1600 B.n706 B.n705 10.6151
R1601 B.n705 B.n702 10.6151
R1602 B.n702 B.n701 10.6151
R1603 B.n701 B.n698 10.6151
R1604 B.n698 B.n697 10.6151
R1605 B.n697 B.n694 10.6151
R1606 B.n694 B.n693 10.6151
R1607 B.n693 B.n690 10.6151
R1608 B.n690 B.n689 10.6151
R1609 B.n686 B.n685 10.6151
R1610 B.n685 B.n682 10.6151
R1611 B.n682 B.n681 10.6151
R1612 B.n681 B.n678 10.6151
R1613 B.n678 B.n677 10.6151
R1614 B.n677 B.n674 10.6151
R1615 B.n674 B.n673 10.6151
R1616 B.n673 B.n670 10.6151
R1617 B.n670 B.n669 10.6151
R1618 B.n666 B.n665 10.6151
R1619 B.n665 B.n662 10.6151
R1620 B.n662 B.n661 10.6151
R1621 B.n661 B.n658 10.6151
R1622 B.n658 B.n657 10.6151
R1623 B.n657 B.n654 10.6151
R1624 B.n654 B.n653 10.6151
R1625 B.n653 B.n650 10.6151
R1626 B.n650 B.n649 10.6151
R1627 B.n649 B.n646 10.6151
R1628 B.n646 B.n645 10.6151
R1629 B.n645 B.n642 10.6151
R1630 B.n642 B.n641 10.6151
R1631 B.n641 B.n638 10.6151
R1632 B.n638 B.n637 10.6151
R1633 B.n637 B.n634 10.6151
R1634 B.n634 B.n633 10.6151
R1635 B.n633 B.n630 10.6151
R1636 B.n630 B.n629 10.6151
R1637 B.n629 B.n626 10.6151
R1638 B.n626 B.n625 10.6151
R1639 B.n625 B.n622 10.6151
R1640 B.n622 B.n621 10.6151
R1641 B.n621 B.n618 10.6151
R1642 B.n618 B.n617 10.6151
R1643 B.n617 B.n614 10.6151
R1644 B.n614 B.n613 10.6151
R1645 B.n613 B.n610 10.6151
R1646 B.n610 B.n609 10.6151
R1647 B.n609 B.n606 10.6151
R1648 B.n606 B.n605 10.6151
R1649 B.n605 B.n602 10.6151
R1650 B.n602 B.n601 10.6151
R1651 B.n601 B.n598 10.6151
R1652 B.n598 B.n597 10.6151
R1653 B.n597 B.n594 10.6151
R1654 B.n594 B.n593 10.6151
R1655 B.n593 B.n590 10.6151
R1656 B.n590 B.n589 10.6151
R1657 B.n589 B.n586 10.6151
R1658 B.n586 B.n585 10.6151
R1659 B.n585 B.n582 10.6151
R1660 B.n582 B.n581 10.6151
R1661 B.n581 B.n578 10.6151
R1662 B.n578 B.n577 10.6151
R1663 B.n577 B.n574 10.6151
R1664 B.n574 B.n573 10.6151
R1665 B.n573 B.n570 10.6151
R1666 B.n570 B.n569 10.6151
R1667 B.n569 B.n566 10.6151
R1668 B.n566 B.n565 10.6151
R1669 B.n565 B.n562 10.6151
R1670 B.n562 B.n561 10.6151
R1671 B.n561 B.n558 10.6151
R1672 B.n558 B.n557 10.6151
R1673 B.n557 B.n554 10.6151
R1674 B.n554 B.n553 10.6151
R1675 B.n553 B.n550 10.6151
R1676 B.n550 B.n549 10.6151
R1677 B.n549 B.n546 10.6151
R1678 B.n546 B.n545 10.6151
R1679 B.n545 B.n542 10.6151
R1680 B.n542 B.n464 10.6151
R1681 B.n819 B.n464 10.6151
R1682 B.n825 B.n460 10.6151
R1683 B.n826 B.n825 10.6151
R1684 B.n827 B.n826 10.6151
R1685 B.n827 B.n452 10.6151
R1686 B.n837 B.n452 10.6151
R1687 B.n838 B.n837 10.6151
R1688 B.n839 B.n838 10.6151
R1689 B.n839 B.n444 10.6151
R1690 B.n849 B.n444 10.6151
R1691 B.n850 B.n849 10.6151
R1692 B.n851 B.n850 10.6151
R1693 B.n851 B.n436 10.6151
R1694 B.n862 B.n436 10.6151
R1695 B.n863 B.n862 10.6151
R1696 B.n864 B.n863 10.6151
R1697 B.n864 B.n429 10.6151
R1698 B.n874 B.n429 10.6151
R1699 B.n875 B.n874 10.6151
R1700 B.n876 B.n875 10.6151
R1701 B.n876 B.n421 10.6151
R1702 B.n886 B.n421 10.6151
R1703 B.n887 B.n886 10.6151
R1704 B.n888 B.n887 10.6151
R1705 B.n888 B.n413 10.6151
R1706 B.n899 B.n413 10.6151
R1707 B.n900 B.n899 10.6151
R1708 B.n901 B.n900 10.6151
R1709 B.n901 B.n0 10.6151
R1710 B.n1001 B.n1 10.6151
R1711 B.n1001 B.n1000 10.6151
R1712 B.n1000 B.n999 10.6151
R1713 B.n999 B.n10 10.6151
R1714 B.n993 B.n10 10.6151
R1715 B.n993 B.n992 10.6151
R1716 B.n992 B.n991 10.6151
R1717 B.n991 B.n17 10.6151
R1718 B.n985 B.n17 10.6151
R1719 B.n985 B.n984 10.6151
R1720 B.n984 B.n983 10.6151
R1721 B.n983 B.n24 10.6151
R1722 B.n977 B.n24 10.6151
R1723 B.n977 B.n976 10.6151
R1724 B.n976 B.n975 10.6151
R1725 B.n975 B.n30 10.6151
R1726 B.n969 B.n30 10.6151
R1727 B.n969 B.n968 10.6151
R1728 B.n968 B.n967 10.6151
R1729 B.n967 B.n38 10.6151
R1730 B.n961 B.n38 10.6151
R1731 B.n961 B.n960 10.6151
R1732 B.n960 B.n959 10.6151
R1733 B.n959 B.n45 10.6151
R1734 B.n953 B.n45 10.6151
R1735 B.n953 B.n952 10.6151
R1736 B.n952 B.n951 10.6151
R1737 B.n951 B.n52 10.6151
R1738 B.t11 B.n450 10.0302
R1739 B.t7 B.n43 10.0302
R1740 B.n260 B.n259 9.36635
R1741 B.n282 B.n281 9.36635
R1742 B.n689 B.n538 9.36635
R1743 B.n666 B.n541 9.36635
R1744 B.n897 B.t0 7.41378
R1745 B.n997 B.t1 7.41378
R1746 B.n859 B.t2 4.79733
R1747 B.n32 B.t4 4.79733
R1748 B.n1007 B.n0 2.81026
R1749 B.n1007 B.n1 2.81026
R1750 B.n261 B.n260 1.24928
R1751 B.n281 B.n280 1.24928
R1752 B.n686 B.n538 1.24928
R1753 B.n669 B.n541 1.24928
R1754 VP.n7 VP.t3 363.995
R1755 VP.n20 VP.t5 327.072
R1756 VP.n14 VP.t1 327.072
R1757 VP.n26 VP.t2 327.072
R1758 VP.n6 VP.t0 327.072
R1759 VP.n12 VP.t4 327.072
R1760 VP.n15 VP.n14 171.088
R1761 VP.n27 VP.n26 171.088
R1762 VP.n13 VP.n12 171.088
R1763 VP.n8 VP.n5 161.3
R1764 VP.n10 VP.n9 161.3
R1765 VP.n11 VP.n4 161.3
R1766 VP.n25 VP.n0 161.3
R1767 VP.n24 VP.n23 161.3
R1768 VP.n22 VP.n1 161.3
R1769 VP.n21 VP.n20 161.3
R1770 VP.n19 VP.n2 161.3
R1771 VP.n18 VP.n17 161.3
R1772 VP.n16 VP.n3 161.3
R1773 VP.n15 VP.n13 50.2581
R1774 VP.n19 VP.n18 50.2061
R1775 VP.n24 VP.n1 50.2061
R1776 VP.n10 VP.n5 50.2061
R1777 VP.n7 VP.n6 41.8683
R1778 VP.n18 VP.n3 30.7807
R1779 VP.n25 VP.n24 30.7807
R1780 VP.n11 VP.n10 30.7807
R1781 VP.n20 VP.n19 24.4675
R1782 VP.n20 VP.n1 24.4675
R1783 VP.n6 VP.n5 24.4675
R1784 VP.n8 VP.n7 17.2768
R1785 VP.n14 VP.n3 14.6807
R1786 VP.n26 VP.n25 14.6807
R1787 VP.n12 VP.n11 14.6807
R1788 VP.n9 VP.n8 0.189894
R1789 VP.n9 VP.n4 0.189894
R1790 VP.n13 VP.n4 0.189894
R1791 VP.n16 VP.n15 0.189894
R1792 VP.n17 VP.n16 0.189894
R1793 VP.n17 VP.n2 0.189894
R1794 VP.n21 VP.n2 0.189894
R1795 VP.n22 VP.n21 0.189894
R1796 VP.n23 VP.n22 0.189894
R1797 VP.n23 VP.n0 0.189894
R1798 VP.n27 VP.n0 0.189894
R1799 VP VP.n27 0.0516364
R1800 VDD1 VDD1.t2 61.0632
R1801 VDD1.n1 VDD1.t4 60.9495
R1802 VDD1.n1 VDD1.n0 59.1813
R1803 VDD1.n3 VDD1.n2 58.8488
R1804 VDD1.n3 VDD1.n1 47.3156
R1805 VDD1.n2 VDD1.t5 0.992981
R1806 VDD1.n2 VDD1.t1 0.992981
R1807 VDD1.n0 VDD1.t0 0.992981
R1808 VDD1.n0 VDD1.t3 0.992981
R1809 VDD1 VDD1.n3 0.330241
C0 VDD1 VDD2 0.996924f
C1 VN VTAIL 9.05233f
C2 VN VDD2 9.475441f
C3 VP VTAIL 9.066969f
C4 VP VDD2 0.363497f
C5 VDD1 VN 0.149137f
C6 VP VDD1 9.68405f
C7 VTAIL VDD2 11.7358f
C8 VP VN 7.297851f
C9 VDD1 VTAIL 11.697201f
C10 VDD2 B 6.515659f
C11 VDD1 B 6.788326f
C12 VTAIL B 10.069888f
C13 VN B 10.49814f
C14 VP B 8.617678f
C15 VDD1.t2 B 4.00834f
C16 VDD1.t4 B 4.00756f
C17 VDD1.t0 B 0.342453f
C18 VDD1.t3 B 0.342453f
C19 VDD1.n0 B 3.1311f
C20 VDD1.n1 B 2.63336f
C21 VDD1.t5 B 0.342453f
C22 VDD1.t1 B 0.342453f
C23 VDD1.n2 B 3.12926f
C24 VDD1.n3 B 2.67827f
C25 VP.n0 B 0.032192f
C26 VP.t2 B 2.60154f
C27 VP.n1 B 0.059084f
C28 VP.n2 B 0.032192f
C29 VP.t5 B 2.60154f
C30 VP.n3 B 0.052643f
C31 VP.n4 B 0.032192f
C32 VP.t4 B 2.60154f
C33 VP.n5 B 0.059084f
C34 VP.t3 B 2.70681f
C35 VP.t0 B 2.60154f
C36 VP.n6 B 0.986693f
C37 VP.n7 B 0.978904f
C38 VP.n8 B 0.205183f
C39 VP.n9 B 0.032192f
C40 VP.n10 B 0.030411f
C41 VP.n11 B 0.052643f
C42 VP.n12 B 0.983184f
C43 VP.n13 B 1.7681f
C44 VP.t1 B 2.60154f
C45 VP.n14 B 0.983184f
C46 VP.n15 B 1.79113f
C47 VP.n16 B 0.032192f
C48 VP.n17 B 0.032192f
C49 VP.n18 B 0.030411f
C50 VP.n19 B 0.059084f
C51 VP.n20 B 0.941914f
C52 VP.n21 B 0.032192f
C53 VP.n22 B 0.032192f
C54 VP.n23 B 0.032192f
C55 VP.n24 B 0.030411f
C56 VP.n25 B 0.052643f
C57 VP.n26 B 0.983184f
C58 VP.n27 B 0.029295f
C59 VDD2.t3 B 3.98505f
C60 VDD2.t0 B 0.340529f
C61 VDD2.t4 B 0.340529f
C62 VDD2.n0 B 3.11351f
C63 VDD2.n1 B 2.5331f
C64 VDD2.t5 B 3.97904f
C65 VDD2.n2 B 2.68437f
C66 VDD2.t2 B 0.340529f
C67 VDD2.t1 B 0.340529f
C68 VDD2.n3 B 3.11348f
C69 VTAIL.t6 B 0.350766f
C70 VTAIL.t8 B 0.350766f
C71 VTAIL.n0 B 3.13216f
C72 VTAIL.n1 B 0.353096f
C73 VTAIL.t0 B 4.00282f
C74 VTAIL.n2 B 0.518333f
C75 VTAIL.t2 B 0.350766f
C76 VTAIL.t3 B 0.350766f
C77 VTAIL.n3 B 3.13216f
C78 VTAIL.n4 B 2.10078f
C79 VTAIL.t5 B 0.350766f
C80 VTAIL.t9 B 0.350766f
C81 VTAIL.n5 B 3.13215f
C82 VTAIL.n6 B 2.10078f
C83 VTAIL.t7 B 4.00284f
C84 VTAIL.n7 B 0.518311f
C85 VTAIL.t1 B 0.350766f
C86 VTAIL.t11 B 0.350766f
C87 VTAIL.n8 B 3.13215f
C88 VTAIL.n9 B 0.432366f
C89 VTAIL.t4 B 4.00283f
C90 VTAIL.n10 B 2.07549f
C91 VTAIL.t10 B 4.00282f
C92 VTAIL.n11 B 2.04352f
C93 VN.n0 B 0.03189f
C94 VN.t1 B 2.57714f
C95 VN.n1 B 0.05853f
C96 VN.t2 B 2.68142f
C97 VN.t5 B 2.57714f
C98 VN.n2 B 0.977438f
C99 VN.n3 B 0.969721f
C100 VN.n4 B 0.203259f
C101 VN.n5 B 0.03189f
C102 VN.n6 B 0.030126f
C103 VN.n7 B 0.052149f
C104 VN.n8 B 0.973961f
C105 VN.n9 B 0.02902f
C106 VN.n10 B 0.03189f
C107 VN.t0 B 2.57714f
C108 VN.n11 B 0.05853f
C109 VN.t4 B 2.68142f
C110 VN.t3 B 2.57714f
C111 VN.n12 B 0.977438f
C112 VN.n13 B 0.969721f
C113 VN.n14 B 0.203259f
C114 VN.n15 B 0.03189f
C115 VN.n16 B 0.030126f
C116 VN.n17 B 0.052149f
C117 VN.n18 B 0.973961f
C118 VN.n19 B 1.77224f
.ends

