* NGSPICE file created from diff_pair_sample_1721.ext - technology: sky130A

.subckt diff_pair_sample_1721 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=2.9
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=2.9
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=2.9
X3 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=2.9
X4 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=2.9
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=2.9
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=1.1505 ps=6.68 w=2.95 l=2.9
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1505 pd=6.68 as=0 ps=0 w=2.95 l=2.9
R0 B.n426 B.n425 585
R1 B.n152 B.n72 585
R2 B.n151 B.n150 585
R3 B.n149 B.n148 585
R4 B.n147 B.n146 585
R5 B.n145 B.n144 585
R6 B.n143 B.n142 585
R7 B.n141 B.n140 585
R8 B.n139 B.n138 585
R9 B.n137 B.n136 585
R10 B.n135 B.n134 585
R11 B.n133 B.n132 585
R12 B.n131 B.n130 585
R13 B.n129 B.n128 585
R14 B.n127 B.n126 585
R15 B.n124 B.n123 585
R16 B.n122 B.n121 585
R17 B.n120 B.n119 585
R18 B.n118 B.n117 585
R19 B.n116 B.n115 585
R20 B.n114 B.n113 585
R21 B.n112 B.n111 585
R22 B.n110 B.n109 585
R23 B.n108 B.n107 585
R24 B.n106 B.n105 585
R25 B.n103 B.n102 585
R26 B.n101 B.n100 585
R27 B.n99 B.n98 585
R28 B.n97 B.n96 585
R29 B.n95 B.n94 585
R30 B.n93 B.n92 585
R31 B.n91 B.n90 585
R32 B.n89 B.n88 585
R33 B.n87 B.n86 585
R34 B.n85 B.n84 585
R35 B.n83 B.n82 585
R36 B.n81 B.n80 585
R37 B.n79 B.n78 585
R38 B.n53 B.n52 585
R39 B.n431 B.n430 585
R40 B.n424 B.n73 585
R41 B.n73 B.n50 585
R42 B.n423 B.n49 585
R43 B.n435 B.n49 585
R44 B.n422 B.n48 585
R45 B.n436 B.n48 585
R46 B.n421 B.n47 585
R47 B.n437 B.n47 585
R48 B.n420 B.n419 585
R49 B.n419 B.n43 585
R50 B.n418 B.n42 585
R51 B.n443 B.n42 585
R52 B.n417 B.n41 585
R53 B.n444 B.n41 585
R54 B.n416 B.n40 585
R55 B.n445 B.n40 585
R56 B.n415 B.n414 585
R57 B.n414 B.n36 585
R58 B.n413 B.n35 585
R59 B.n451 B.n35 585
R60 B.n412 B.n34 585
R61 B.n452 B.n34 585
R62 B.n411 B.n33 585
R63 B.n453 B.n33 585
R64 B.n410 B.n409 585
R65 B.n409 B.n29 585
R66 B.n408 B.n28 585
R67 B.n459 B.n28 585
R68 B.n407 B.n27 585
R69 B.n460 B.n27 585
R70 B.n406 B.n26 585
R71 B.n461 B.n26 585
R72 B.n405 B.n404 585
R73 B.n404 B.n22 585
R74 B.n403 B.n21 585
R75 B.n467 B.n21 585
R76 B.n402 B.n20 585
R77 B.n468 B.n20 585
R78 B.n401 B.n19 585
R79 B.n469 B.n19 585
R80 B.n400 B.n399 585
R81 B.n399 B.n18 585
R82 B.n398 B.n14 585
R83 B.n475 B.n14 585
R84 B.n397 B.n13 585
R85 B.n476 B.n13 585
R86 B.n396 B.n12 585
R87 B.n477 B.n12 585
R88 B.n395 B.n394 585
R89 B.n394 B.n8 585
R90 B.n393 B.n7 585
R91 B.n483 B.n7 585
R92 B.n392 B.n6 585
R93 B.n484 B.n6 585
R94 B.n391 B.n5 585
R95 B.n485 B.n5 585
R96 B.n390 B.n389 585
R97 B.n389 B.n4 585
R98 B.n388 B.n153 585
R99 B.n388 B.n387 585
R100 B.n378 B.n154 585
R101 B.n155 B.n154 585
R102 B.n380 B.n379 585
R103 B.n381 B.n380 585
R104 B.n377 B.n160 585
R105 B.n160 B.n159 585
R106 B.n376 B.n375 585
R107 B.n375 B.n374 585
R108 B.n162 B.n161 585
R109 B.n367 B.n162 585
R110 B.n366 B.n365 585
R111 B.n368 B.n366 585
R112 B.n364 B.n167 585
R113 B.n167 B.n166 585
R114 B.n363 B.n362 585
R115 B.n362 B.n361 585
R116 B.n169 B.n168 585
R117 B.n170 B.n169 585
R118 B.n354 B.n353 585
R119 B.n355 B.n354 585
R120 B.n352 B.n175 585
R121 B.n175 B.n174 585
R122 B.n351 B.n350 585
R123 B.n350 B.n349 585
R124 B.n177 B.n176 585
R125 B.n178 B.n177 585
R126 B.n342 B.n341 585
R127 B.n343 B.n342 585
R128 B.n340 B.n183 585
R129 B.n183 B.n182 585
R130 B.n339 B.n338 585
R131 B.n338 B.n337 585
R132 B.n185 B.n184 585
R133 B.n186 B.n185 585
R134 B.n330 B.n329 585
R135 B.n331 B.n330 585
R136 B.n328 B.n191 585
R137 B.n191 B.n190 585
R138 B.n327 B.n326 585
R139 B.n326 B.n325 585
R140 B.n193 B.n192 585
R141 B.n194 B.n193 585
R142 B.n318 B.n317 585
R143 B.n319 B.n318 585
R144 B.n316 B.n199 585
R145 B.n199 B.n198 585
R146 B.n315 B.n314 585
R147 B.n314 B.n313 585
R148 B.n201 B.n200 585
R149 B.n202 B.n201 585
R150 B.n309 B.n308 585
R151 B.n205 B.n204 585
R152 B.n305 B.n304 585
R153 B.n306 B.n305 585
R154 B.n303 B.n225 585
R155 B.n302 B.n301 585
R156 B.n300 B.n299 585
R157 B.n298 B.n297 585
R158 B.n296 B.n295 585
R159 B.n294 B.n293 585
R160 B.n292 B.n291 585
R161 B.n290 B.n289 585
R162 B.n288 B.n287 585
R163 B.n286 B.n285 585
R164 B.n284 B.n283 585
R165 B.n282 B.n281 585
R166 B.n280 B.n279 585
R167 B.n278 B.n277 585
R168 B.n276 B.n275 585
R169 B.n274 B.n273 585
R170 B.n272 B.n271 585
R171 B.n270 B.n269 585
R172 B.n268 B.n267 585
R173 B.n266 B.n265 585
R174 B.n264 B.n263 585
R175 B.n262 B.n261 585
R176 B.n260 B.n259 585
R177 B.n258 B.n257 585
R178 B.n256 B.n255 585
R179 B.n254 B.n253 585
R180 B.n252 B.n251 585
R181 B.n250 B.n249 585
R182 B.n248 B.n247 585
R183 B.n246 B.n245 585
R184 B.n244 B.n243 585
R185 B.n242 B.n241 585
R186 B.n240 B.n239 585
R187 B.n238 B.n237 585
R188 B.n236 B.n235 585
R189 B.n234 B.n233 585
R190 B.n232 B.n224 585
R191 B.n306 B.n224 585
R192 B.n310 B.n203 585
R193 B.n203 B.n202 585
R194 B.n312 B.n311 585
R195 B.n313 B.n312 585
R196 B.n197 B.n196 585
R197 B.n198 B.n197 585
R198 B.n321 B.n320 585
R199 B.n320 B.n319 585
R200 B.n322 B.n195 585
R201 B.n195 B.n194 585
R202 B.n324 B.n323 585
R203 B.n325 B.n324 585
R204 B.n189 B.n188 585
R205 B.n190 B.n189 585
R206 B.n333 B.n332 585
R207 B.n332 B.n331 585
R208 B.n334 B.n187 585
R209 B.n187 B.n186 585
R210 B.n336 B.n335 585
R211 B.n337 B.n336 585
R212 B.n181 B.n180 585
R213 B.n182 B.n181 585
R214 B.n345 B.n344 585
R215 B.n344 B.n343 585
R216 B.n346 B.n179 585
R217 B.n179 B.n178 585
R218 B.n348 B.n347 585
R219 B.n349 B.n348 585
R220 B.n173 B.n172 585
R221 B.n174 B.n173 585
R222 B.n357 B.n356 585
R223 B.n356 B.n355 585
R224 B.n358 B.n171 585
R225 B.n171 B.n170 585
R226 B.n360 B.n359 585
R227 B.n361 B.n360 585
R228 B.n165 B.n164 585
R229 B.n166 B.n165 585
R230 B.n370 B.n369 585
R231 B.n369 B.n368 585
R232 B.n371 B.n163 585
R233 B.n367 B.n163 585
R234 B.n373 B.n372 585
R235 B.n374 B.n373 585
R236 B.n158 B.n157 585
R237 B.n159 B.n158 585
R238 B.n383 B.n382 585
R239 B.n382 B.n381 585
R240 B.n384 B.n156 585
R241 B.n156 B.n155 585
R242 B.n386 B.n385 585
R243 B.n387 B.n386 585
R244 B.n2 B.n0 585
R245 B.n4 B.n2 585
R246 B.n3 B.n1 585
R247 B.n484 B.n3 585
R248 B.n482 B.n481 585
R249 B.n483 B.n482 585
R250 B.n480 B.n9 585
R251 B.n9 B.n8 585
R252 B.n479 B.n478 585
R253 B.n478 B.n477 585
R254 B.n11 B.n10 585
R255 B.n476 B.n11 585
R256 B.n474 B.n473 585
R257 B.n475 B.n474 585
R258 B.n472 B.n15 585
R259 B.n18 B.n15 585
R260 B.n471 B.n470 585
R261 B.n470 B.n469 585
R262 B.n17 B.n16 585
R263 B.n468 B.n17 585
R264 B.n466 B.n465 585
R265 B.n467 B.n466 585
R266 B.n464 B.n23 585
R267 B.n23 B.n22 585
R268 B.n463 B.n462 585
R269 B.n462 B.n461 585
R270 B.n25 B.n24 585
R271 B.n460 B.n25 585
R272 B.n458 B.n457 585
R273 B.n459 B.n458 585
R274 B.n456 B.n30 585
R275 B.n30 B.n29 585
R276 B.n455 B.n454 585
R277 B.n454 B.n453 585
R278 B.n32 B.n31 585
R279 B.n452 B.n32 585
R280 B.n450 B.n449 585
R281 B.n451 B.n450 585
R282 B.n448 B.n37 585
R283 B.n37 B.n36 585
R284 B.n447 B.n446 585
R285 B.n446 B.n445 585
R286 B.n39 B.n38 585
R287 B.n444 B.n39 585
R288 B.n442 B.n441 585
R289 B.n443 B.n442 585
R290 B.n440 B.n44 585
R291 B.n44 B.n43 585
R292 B.n439 B.n438 585
R293 B.n438 B.n437 585
R294 B.n46 B.n45 585
R295 B.n436 B.n46 585
R296 B.n434 B.n433 585
R297 B.n435 B.n434 585
R298 B.n432 B.n51 585
R299 B.n51 B.n50 585
R300 B.n487 B.n486 585
R301 B.n486 B.n485 585
R302 B.n308 B.n203 482.89
R303 B.n430 B.n51 482.89
R304 B.n224 B.n201 482.89
R305 B.n426 B.n73 482.89
R306 B.n428 B.n427 256.663
R307 B.n428 B.n71 256.663
R308 B.n428 B.n70 256.663
R309 B.n428 B.n69 256.663
R310 B.n428 B.n68 256.663
R311 B.n428 B.n67 256.663
R312 B.n428 B.n66 256.663
R313 B.n428 B.n65 256.663
R314 B.n428 B.n64 256.663
R315 B.n428 B.n63 256.663
R316 B.n428 B.n62 256.663
R317 B.n428 B.n61 256.663
R318 B.n428 B.n60 256.663
R319 B.n428 B.n59 256.663
R320 B.n428 B.n58 256.663
R321 B.n428 B.n57 256.663
R322 B.n428 B.n56 256.663
R323 B.n428 B.n55 256.663
R324 B.n428 B.n54 256.663
R325 B.n429 B.n428 256.663
R326 B.n307 B.n306 256.663
R327 B.n306 B.n206 256.663
R328 B.n306 B.n207 256.663
R329 B.n306 B.n208 256.663
R330 B.n306 B.n209 256.663
R331 B.n306 B.n210 256.663
R332 B.n306 B.n211 256.663
R333 B.n306 B.n212 256.663
R334 B.n306 B.n213 256.663
R335 B.n306 B.n214 256.663
R336 B.n306 B.n215 256.663
R337 B.n306 B.n216 256.663
R338 B.n306 B.n217 256.663
R339 B.n306 B.n218 256.663
R340 B.n306 B.n219 256.663
R341 B.n306 B.n220 256.663
R342 B.n306 B.n221 256.663
R343 B.n306 B.n222 256.663
R344 B.n306 B.n223 256.663
R345 B.n229 B.t10 232.975
R346 B.n226 B.t6 232.975
R347 B.n76 B.t2 232.975
R348 B.n74 B.t13 232.975
R349 B.n306 B.n202 175.198
R350 B.n428 B.n50 175.198
R351 B.n312 B.n203 163.367
R352 B.n312 B.n197 163.367
R353 B.n320 B.n197 163.367
R354 B.n320 B.n195 163.367
R355 B.n324 B.n195 163.367
R356 B.n324 B.n189 163.367
R357 B.n332 B.n189 163.367
R358 B.n332 B.n187 163.367
R359 B.n336 B.n187 163.367
R360 B.n336 B.n181 163.367
R361 B.n344 B.n181 163.367
R362 B.n344 B.n179 163.367
R363 B.n348 B.n179 163.367
R364 B.n348 B.n173 163.367
R365 B.n356 B.n173 163.367
R366 B.n356 B.n171 163.367
R367 B.n360 B.n171 163.367
R368 B.n360 B.n165 163.367
R369 B.n369 B.n165 163.367
R370 B.n369 B.n163 163.367
R371 B.n373 B.n163 163.367
R372 B.n373 B.n158 163.367
R373 B.n382 B.n158 163.367
R374 B.n382 B.n156 163.367
R375 B.n386 B.n156 163.367
R376 B.n386 B.n2 163.367
R377 B.n486 B.n2 163.367
R378 B.n486 B.n3 163.367
R379 B.n482 B.n3 163.367
R380 B.n482 B.n9 163.367
R381 B.n478 B.n9 163.367
R382 B.n478 B.n11 163.367
R383 B.n474 B.n11 163.367
R384 B.n474 B.n15 163.367
R385 B.n470 B.n15 163.367
R386 B.n470 B.n17 163.367
R387 B.n466 B.n17 163.367
R388 B.n466 B.n23 163.367
R389 B.n462 B.n23 163.367
R390 B.n462 B.n25 163.367
R391 B.n458 B.n25 163.367
R392 B.n458 B.n30 163.367
R393 B.n454 B.n30 163.367
R394 B.n454 B.n32 163.367
R395 B.n450 B.n32 163.367
R396 B.n450 B.n37 163.367
R397 B.n446 B.n37 163.367
R398 B.n446 B.n39 163.367
R399 B.n442 B.n39 163.367
R400 B.n442 B.n44 163.367
R401 B.n438 B.n44 163.367
R402 B.n438 B.n46 163.367
R403 B.n434 B.n46 163.367
R404 B.n434 B.n51 163.367
R405 B.n305 B.n205 163.367
R406 B.n305 B.n225 163.367
R407 B.n301 B.n300 163.367
R408 B.n297 B.n296 163.367
R409 B.n293 B.n292 163.367
R410 B.n289 B.n288 163.367
R411 B.n285 B.n284 163.367
R412 B.n281 B.n280 163.367
R413 B.n277 B.n276 163.367
R414 B.n273 B.n272 163.367
R415 B.n269 B.n268 163.367
R416 B.n265 B.n264 163.367
R417 B.n261 B.n260 163.367
R418 B.n257 B.n256 163.367
R419 B.n253 B.n252 163.367
R420 B.n249 B.n248 163.367
R421 B.n245 B.n244 163.367
R422 B.n241 B.n240 163.367
R423 B.n237 B.n236 163.367
R424 B.n233 B.n224 163.367
R425 B.n314 B.n201 163.367
R426 B.n314 B.n199 163.367
R427 B.n318 B.n199 163.367
R428 B.n318 B.n193 163.367
R429 B.n326 B.n193 163.367
R430 B.n326 B.n191 163.367
R431 B.n330 B.n191 163.367
R432 B.n330 B.n185 163.367
R433 B.n338 B.n185 163.367
R434 B.n338 B.n183 163.367
R435 B.n342 B.n183 163.367
R436 B.n342 B.n177 163.367
R437 B.n350 B.n177 163.367
R438 B.n350 B.n175 163.367
R439 B.n354 B.n175 163.367
R440 B.n354 B.n169 163.367
R441 B.n362 B.n169 163.367
R442 B.n362 B.n167 163.367
R443 B.n366 B.n167 163.367
R444 B.n366 B.n162 163.367
R445 B.n375 B.n162 163.367
R446 B.n375 B.n160 163.367
R447 B.n380 B.n160 163.367
R448 B.n380 B.n154 163.367
R449 B.n388 B.n154 163.367
R450 B.n389 B.n388 163.367
R451 B.n389 B.n5 163.367
R452 B.n6 B.n5 163.367
R453 B.n7 B.n6 163.367
R454 B.n394 B.n7 163.367
R455 B.n394 B.n12 163.367
R456 B.n13 B.n12 163.367
R457 B.n14 B.n13 163.367
R458 B.n399 B.n14 163.367
R459 B.n399 B.n19 163.367
R460 B.n20 B.n19 163.367
R461 B.n21 B.n20 163.367
R462 B.n404 B.n21 163.367
R463 B.n404 B.n26 163.367
R464 B.n27 B.n26 163.367
R465 B.n28 B.n27 163.367
R466 B.n409 B.n28 163.367
R467 B.n409 B.n33 163.367
R468 B.n34 B.n33 163.367
R469 B.n35 B.n34 163.367
R470 B.n414 B.n35 163.367
R471 B.n414 B.n40 163.367
R472 B.n41 B.n40 163.367
R473 B.n42 B.n41 163.367
R474 B.n419 B.n42 163.367
R475 B.n419 B.n47 163.367
R476 B.n48 B.n47 163.367
R477 B.n49 B.n48 163.367
R478 B.n73 B.n49 163.367
R479 B.n78 B.n53 163.367
R480 B.n82 B.n81 163.367
R481 B.n86 B.n85 163.367
R482 B.n90 B.n89 163.367
R483 B.n94 B.n93 163.367
R484 B.n98 B.n97 163.367
R485 B.n102 B.n101 163.367
R486 B.n107 B.n106 163.367
R487 B.n111 B.n110 163.367
R488 B.n115 B.n114 163.367
R489 B.n119 B.n118 163.367
R490 B.n123 B.n122 163.367
R491 B.n128 B.n127 163.367
R492 B.n132 B.n131 163.367
R493 B.n136 B.n135 163.367
R494 B.n140 B.n139 163.367
R495 B.n144 B.n143 163.367
R496 B.n148 B.n147 163.367
R497 B.n150 B.n72 163.367
R498 B.n229 B.t12 142.399
R499 B.n74 B.t14 142.399
R500 B.n226 B.t9 142.398
R501 B.n76 B.t4 142.398
R502 B.n313 B.n202 90.9428
R503 B.n313 B.n198 90.9428
R504 B.n319 B.n198 90.9428
R505 B.n319 B.n194 90.9428
R506 B.n325 B.n194 90.9428
R507 B.n325 B.n190 90.9428
R508 B.n331 B.n190 90.9428
R509 B.n337 B.n186 90.9428
R510 B.n337 B.n182 90.9428
R511 B.n343 B.n182 90.9428
R512 B.n343 B.n178 90.9428
R513 B.n349 B.n178 90.9428
R514 B.n349 B.n174 90.9428
R515 B.n355 B.n174 90.9428
R516 B.n355 B.n170 90.9428
R517 B.n361 B.n170 90.9428
R518 B.n361 B.n166 90.9428
R519 B.n368 B.n166 90.9428
R520 B.n368 B.n367 90.9428
R521 B.n374 B.n159 90.9428
R522 B.n381 B.n159 90.9428
R523 B.n381 B.n155 90.9428
R524 B.n387 B.n155 90.9428
R525 B.n387 B.n4 90.9428
R526 B.n485 B.n4 90.9428
R527 B.n485 B.n484 90.9428
R528 B.n484 B.n483 90.9428
R529 B.n483 B.n8 90.9428
R530 B.n477 B.n8 90.9428
R531 B.n477 B.n476 90.9428
R532 B.n476 B.n475 90.9428
R533 B.n469 B.n18 90.9428
R534 B.n469 B.n468 90.9428
R535 B.n468 B.n467 90.9428
R536 B.n467 B.n22 90.9428
R537 B.n461 B.n22 90.9428
R538 B.n461 B.n460 90.9428
R539 B.n460 B.n459 90.9428
R540 B.n459 B.n29 90.9428
R541 B.n453 B.n29 90.9428
R542 B.n453 B.n452 90.9428
R543 B.n452 B.n451 90.9428
R544 B.n451 B.n36 90.9428
R545 B.n445 B.n444 90.9428
R546 B.n444 B.n443 90.9428
R547 B.n443 B.n43 90.9428
R548 B.n437 B.n43 90.9428
R549 B.n437 B.n436 90.9428
R550 B.n436 B.n435 90.9428
R551 B.n435 B.n50 90.9428
R552 B.n331 B.t7 85.5932
R553 B.n445 B.t3 85.5932
R554 B.n230 B.t11 79.757
R555 B.n75 B.t15 79.757
R556 B.n227 B.t8 79.7551
R557 B.n77 B.t5 79.7551
R558 B.n308 B.n307 71.676
R559 B.n225 B.n206 71.676
R560 B.n300 B.n207 71.676
R561 B.n296 B.n208 71.676
R562 B.n292 B.n209 71.676
R563 B.n288 B.n210 71.676
R564 B.n284 B.n211 71.676
R565 B.n280 B.n212 71.676
R566 B.n276 B.n213 71.676
R567 B.n272 B.n214 71.676
R568 B.n268 B.n215 71.676
R569 B.n264 B.n216 71.676
R570 B.n260 B.n217 71.676
R571 B.n256 B.n218 71.676
R572 B.n252 B.n219 71.676
R573 B.n248 B.n220 71.676
R574 B.n244 B.n221 71.676
R575 B.n240 B.n222 71.676
R576 B.n236 B.n223 71.676
R577 B.n430 B.n429 71.676
R578 B.n78 B.n54 71.676
R579 B.n82 B.n55 71.676
R580 B.n86 B.n56 71.676
R581 B.n90 B.n57 71.676
R582 B.n94 B.n58 71.676
R583 B.n98 B.n59 71.676
R584 B.n102 B.n60 71.676
R585 B.n107 B.n61 71.676
R586 B.n111 B.n62 71.676
R587 B.n115 B.n63 71.676
R588 B.n119 B.n64 71.676
R589 B.n123 B.n65 71.676
R590 B.n128 B.n66 71.676
R591 B.n132 B.n67 71.676
R592 B.n136 B.n68 71.676
R593 B.n140 B.n69 71.676
R594 B.n144 B.n70 71.676
R595 B.n148 B.n71 71.676
R596 B.n427 B.n72 71.676
R597 B.n427 B.n426 71.676
R598 B.n150 B.n71 71.676
R599 B.n147 B.n70 71.676
R600 B.n143 B.n69 71.676
R601 B.n139 B.n68 71.676
R602 B.n135 B.n67 71.676
R603 B.n131 B.n66 71.676
R604 B.n127 B.n65 71.676
R605 B.n122 B.n64 71.676
R606 B.n118 B.n63 71.676
R607 B.n114 B.n62 71.676
R608 B.n110 B.n61 71.676
R609 B.n106 B.n60 71.676
R610 B.n101 B.n59 71.676
R611 B.n97 B.n58 71.676
R612 B.n93 B.n57 71.676
R613 B.n89 B.n56 71.676
R614 B.n85 B.n55 71.676
R615 B.n81 B.n54 71.676
R616 B.n429 B.n53 71.676
R617 B.n307 B.n205 71.676
R618 B.n301 B.n206 71.676
R619 B.n297 B.n207 71.676
R620 B.n293 B.n208 71.676
R621 B.n289 B.n209 71.676
R622 B.n285 B.n210 71.676
R623 B.n281 B.n211 71.676
R624 B.n277 B.n212 71.676
R625 B.n273 B.n213 71.676
R626 B.n269 B.n214 71.676
R627 B.n265 B.n215 71.676
R628 B.n261 B.n216 71.676
R629 B.n257 B.n217 71.676
R630 B.n253 B.n218 71.676
R631 B.n249 B.n219 71.676
R632 B.n245 B.n220 71.676
R633 B.n241 B.n221 71.676
R634 B.n237 B.n222 71.676
R635 B.n233 B.n223 71.676
R636 B.n230 B.n229 62.6429
R637 B.n227 B.n226 62.6429
R638 B.n77 B.n76 62.6429
R639 B.n75 B.n74 62.6429
R640 B.n231 B.n230 59.5399
R641 B.n228 B.n227 59.5399
R642 B.n104 B.n77 59.5399
R643 B.n125 B.n75 59.5399
R644 B.n367 B.t1 58.8455
R645 B.n18 B.t0 58.8455
R646 B.n374 B.t1 32.0978
R647 B.n475 B.t0 32.0978
R648 B.n432 B.n431 31.3761
R649 B.n425 B.n424 31.3761
R650 B.n232 B.n200 31.3761
R651 B.n310 B.n309 31.3761
R652 B B.n487 18.0485
R653 B.n431 B.n52 10.6151
R654 B.n79 B.n52 10.6151
R655 B.n80 B.n79 10.6151
R656 B.n83 B.n80 10.6151
R657 B.n84 B.n83 10.6151
R658 B.n87 B.n84 10.6151
R659 B.n88 B.n87 10.6151
R660 B.n91 B.n88 10.6151
R661 B.n92 B.n91 10.6151
R662 B.n95 B.n92 10.6151
R663 B.n96 B.n95 10.6151
R664 B.n99 B.n96 10.6151
R665 B.n100 B.n99 10.6151
R666 B.n103 B.n100 10.6151
R667 B.n108 B.n105 10.6151
R668 B.n109 B.n108 10.6151
R669 B.n112 B.n109 10.6151
R670 B.n113 B.n112 10.6151
R671 B.n116 B.n113 10.6151
R672 B.n117 B.n116 10.6151
R673 B.n120 B.n117 10.6151
R674 B.n121 B.n120 10.6151
R675 B.n124 B.n121 10.6151
R676 B.n129 B.n126 10.6151
R677 B.n130 B.n129 10.6151
R678 B.n133 B.n130 10.6151
R679 B.n134 B.n133 10.6151
R680 B.n137 B.n134 10.6151
R681 B.n138 B.n137 10.6151
R682 B.n141 B.n138 10.6151
R683 B.n142 B.n141 10.6151
R684 B.n145 B.n142 10.6151
R685 B.n146 B.n145 10.6151
R686 B.n149 B.n146 10.6151
R687 B.n151 B.n149 10.6151
R688 B.n152 B.n151 10.6151
R689 B.n425 B.n152 10.6151
R690 B.n315 B.n200 10.6151
R691 B.n316 B.n315 10.6151
R692 B.n317 B.n316 10.6151
R693 B.n317 B.n192 10.6151
R694 B.n327 B.n192 10.6151
R695 B.n328 B.n327 10.6151
R696 B.n329 B.n328 10.6151
R697 B.n329 B.n184 10.6151
R698 B.n339 B.n184 10.6151
R699 B.n340 B.n339 10.6151
R700 B.n341 B.n340 10.6151
R701 B.n341 B.n176 10.6151
R702 B.n351 B.n176 10.6151
R703 B.n352 B.n351 10.6151
R704 B.n353 B.n352 10.6151
R705 B.n353 B.n168 10.6151
R706 B.n363 B.n168 10.6151
R707 B.n364 B.n363 10.6151
R708 B.n365 B.n364 10.6151
R709 B.n365 B.n161 10.6151
R710 B.n376 B.n161 10.6151
R711 B.n377 B.n376 10.6151
R712 B.n379 B.n377 10.6151
R713 B.n379 B.n378 10.6151
R714 B.n378 B.n153 10.6151
R715 B.n390 B.n153 10.6151
R716 B.n391 B.n390 10.6151
R717 B.n392 B.n391 10.6151
R718 B.n393 B.n392 10.6151
R719 B.n395 B.n393 10.6151
R720 B.n396 B.n395 10.6151
R721 B.n397 B.n396 10.6151
R722 B.n398 B.n397 10.6151
R723 B.n400 B.n398 10.6151
R724 B.n401 B.n400 10.6151
R725 B.n402 B.n401 10.6151
R726 B.n403 B.n402 10.6151
R727 B.n405 B.n403 10.6151
R728 B.n406 B.n405 10.6151
R729 B.n407 B.n406 10.6151
R730 B.n408 B.n407 10.6151
R731 B.n410 B.n408 10.6151
R732 B.n411 B.n410 10.6151
R733 B.n412 B.n411 10.6151
R734 B.n413 B.n412 10.6151
R735 B.n415 B.n413 10.6151
R736 B.n416 B.n415 10.6151
R737 B.n417 B.n416 10.6151
R738 B.n418 B.n417 10.6151
R739 B.n420 B.n418 10.6151
R740 B.n421 B.n420 10.6151
R741 B.n422 B.n421 10.6151
R742 B.n423 B.n422 10.6151
R743 B.n424 B.n423 10.6151
R744 B.n309 B.n204 10.6151
R745 B.n304 B.n204 10.6151
R746 B.n304 B.n303 10.6151
R747 B.n303 B.n302 10.6151
R748 B.n302 B.n299 10.6151
R749 B.n299 B.n298 10.6151
R750 B.n298 B.n295 10.6151
R751 B.n295 B.n294 10.6151
R752 B.n294 B.n291 10.6151
R753 B.n291 B.n290 10.6151
R754 B.n290 B.n287 10.6151
R755 B.n287 B.n286 10.6151
R756 B.n286 B.n283 10.6151
R757 B.n283 B.n282 10.6151
R758 B.n279 B.n278 10.6151
R759 B.n278 B.n275 10.6151
R760 B.n275 B.n274 10.6151
R761 B.n274 B.n271 10.6151
R762 B.n271 B.n270 10.6151
R763 B.n270 B.n267 10.6151
R764 B.n267 B.n266 10.6151
R765 B.n266 B.n263 10.6151
R766 B.n263 B.n262 10.6151
R767 B.n259 B.n258 10.6151
R768 B.n258 B.n255 10.6151
R769 B.n255 B.n254 10.6151
R770 B.n254 B.n251 10.6151
R771 B.n251 B.n250 10.6151
R772 B.n250 B.n247 10.6151
R773 B.n247 B.n246 10.6151
R774 B.n246 B.n243 10.6151
R775 B.n243 B.n242 10.6151
R776 B.n242 B.n239 10.6151
R777 B.n239 B.n238 10.6151
R778 B.n238 B.n235 10.6151
R779 B.n235 B.n234 10.6151
R780 B.n234 B.n232 10.6151
R781 B.n311 B.n310 10.6151
R782 B.n311 B.n196 10.6151
R783 B.n321 B.n196 10.6151
R784 B.n322 B.n321 10.6151
R785 B.n323 B.n322 10.6151
R786 B.n323 B.n188 10.6151
R787 B.n333 B.n188 10.6151
R788 B.n334 B.n333 10.6151
R789 B.n335 B.n334 10.6151
R790 B.n335 B.n180 10.6151
R791 B.n345 B.n180 10.6151
R792 B.n346 B.n345 10.6151
R793 B.n347 B.n346 10.6151
R794 B.n347 B.n172 10.6151
R795 B.n357 B.n172 10.6151
R796 B.n358 B.n357 10.6151
R797 B.n359 B.n358 10.6151
R798 B.n359 B.n164 10.6151
R799 B.n370 B.n164 10.6151
R800 B.n371 B.n370 10.6151
R801 B.n372 B.n371 10.6151
R802 B.n372 B.n157 10.6151
R803 B.n383 B.n157 10.6151
R804 B.n384 B.n383 10.6151
R805 B.n385 B.n384 10.6151
R806 B.n385 B.n0 10.6151
R807 B.n481 B.n1 10.6151
R808 B.n481 B.n480 10.6151
R809 B.n480 B.n479 10.6151
R810 B.n479 B.n10 10.6151
R811 B.n473 B.n10 10.6151
R812 B.n473 B.n472 10.6151
R813 B.n472 B.n471 10.6151
R814 B.n471 B.n16 10.6151
R815 B.n465 B.n16 10.6151
R816 B.n465 B.n464 10.6151
R817 B.n464 B.n463 10.6151
R818 B.n463 B.n24 10.6151
R819 B.n457 B.n24 10.6151
R820 B.n457 B.n456 10.6151
R821 B.n456 B.n455 10.6151
R822 B.n455 B.n31 10.6151
R823 B.n449 B.n31 10.6151
R824 B.n449 B.n448 10.6151
R825 B.n448 B.n447 10.6151
R826 B.n447 B.n38 10.6151
R827 B.n441 B.n38 10.6151
R828 B.n441 B.n440 10.6151
R829 B.n440 B.n439 10.6151
R830 B.n439 B.n45 10.6151
R831 B.n433 B.n45 10.6151
R832 B.n433 B.n432 10.6151
R833 B.n104 B.n103 9.36635
R834 B.n126 B.n125 9.36635
R835 B.n282 B.n228 9.36635
R836 B.n259 B.n231 9.36635
R837 B.t7 B.n186 5.35004
R838 B.t3 B.n36 5.35004
R839 B.n487 B.n0 2.81026
R840 B.n487 B.n1 2.81026
R841 B.n105 B.n104 1.24928
R842 B.n125 B.n124 1.24928
R843 B.n279 B.n228 1.24928
R844 B.n262 B.n231 1.24928
R845 VP.n0 VP.t0 104.209
R846 VP.n0 VP.t1 65.6117
R847 VP VP.n0 0.431811
R848 VTAIL.n1 VTAIL.t1 74.5465
R849 VTAIL.n3 VTAIL.t0 74.5463
R850 VTAIL.n0 VTAIL.t2 74.5463
R851 VTAIL.n2 VTAIL.t3 74.5463
R852 VTAIL.n1 VTAIL.n0 20.4789
R853 VTAIL.n3 VTAIL.n2 17.6945
R854 VTAIL.n2 VTAIL.n1 1.86257
R855 VTAIL VTAIL.n0 1.22464
R856 VTAIL VTAIL.n3 0.638431
R857 VDD1 VDD1.t0 124.218
R858 VDD1 VDD1.t1 91.9794
R859 VN VN.t0 104.21
R860 VN VN.t1 66.043
R861 VDD2.n0 VDD2.t0 122.996
R862 VDD2.n0 VDD2.t1 91.2251
R863 VDD2 VDD2.n0 0.75481
C0 VN VP 3.92696f
C1 VDD1 VN 0.153405f
C2 VTAIL VN 1.1353f
C3 VDD1 VP 1.08407f
C4 VDD2 VN 0.888315f
C5 VTAIL VP 1.14945f
C6 VDD1 VTAIL 2.76711f
C7 VDD2 VP 0.350686f
C8 VDD1 VDD2 0.71f
C9 VTAIL VDD2 2.82192f
C10 VDD2 B 2.870903f
C11 VDD1 B 4.82531f
C12 VTAIL B 3.515835f
C13 VN B 7.96756f
C14 VP B 5.966f
C15 VDD2.t0 B 0.574962f
C16 VDD2.t1 B 0.365514f
C17 VDD2.n0 B 1.74392f
C18 VN.t1 B 0.769342f
C19 VN.t0 B 1.19755f
C20 VDD1.t1 B 0.359258f
C21 VDD1.t0 B 0.582631f
C22 VTAIL.t2 B 0.393743f
C23 VTAIL.n0 B 1.05421f
C24 VTAIL.t1 B 0.393745f
C25 VTAIL.n1 B 1.09476f
C26 VTAIL.t3 B 0.393743f
C27 VTAIL.n2 B 0.91775f
C28 VTAIL.t0 B 0.393743f
C29 VTAIL.n3 B 0.839929f
C30 VP.t1 B 0.774366f
C31 VP.t0 B 1.20556f
C32 VP.n0 B 1.84928f
.ends

