* NGSPICE file created from diff_pair_sample_1534.ext - technology: sky130A

.subckt diff_pair_sample_1534 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=7.7493 ps=40.52 w=19.87 l=0.28
X1 B.t11 B.t9 B.t10 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=0 ps=0 w=19.87 l=0.28
X2 VDD1.t1 VP.t0 VTAIL.t0 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=7.7493 ps=40.52 w=19.87 l=0.28
X3 B.t8 B.t6 B.t7 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=0 ps=0 w=19.87 l=0.28
X4 VDD1.t0 VP.t1 VTAIL.t1 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=7.7493 ps=40.52 w=19.87 l=0.28
X5 B.t5 B.t3 B.t4 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=0 ps=0 w=19.87 l=0.28
X6 VDD2.t0 VN.t1 VTAIL.t2 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=7.7493 ps=40.52 w=19.87 l=0.28
X7 B.t2 B.t0 B.t1 w_n1214_n4946# sky130_fd_pr__pfet_01v8 ad=7.7493 pd=40.52 as=0 ps=0 w=19.87 l=0.28
R0 VN VN.t1 2053.25
R1 VN VN.t0 2008.44
R2 VTAIL.n1 VTAIL.t2 56.3641
R3 VTAIL.n3 VTAIL.t3 56.3639
R4 VTAIL.n0 VTAIL.t1 56.3639
R5 VTAIL.n2 VTAIL.t0 56.3639
R6 VTAIL.n1 VTAIL.n0 30.5652
R7 VTAIL.n3 VTAIL.n2 30.0393
R8 VTAIL.n2 VTAIL.n1 0.733259
R9 VTAIL VTAIL.n0 0.659983
R10 VTAIL VTAIL.n3 0.0737759
R11 VDD2.n0 VDD2.t1 114.9
R12 VDD2.n0 VDD2.t0 73.0427
R13 VDD2 VDD2.n0 0.190155
R14 B.n134 B.t3 1929.38
R15 B.n126 B.t9 1929.38
R16 B.n48 B.t6 1929.38
R17 B.n40 B.t0 1929.38
R18 B.n397 B.n396 585
R19 B.n395 B.n94 585
R20 B.n394 B.n393 585
R21 B.n392 B.n95 585
R22 B.n391 B.n390 585
R23 B.n389 B.n96 585
R24 B.n388 B.n387 585
R25 B.n386 B.n97 585
R26 B.n385 B.n384 585
R27 B.n383 B.n98 585
R28 B.n382 B.n381 585
R29 B.n380 B.n99 585
R30 B.n379 B.n378 585
R31 B.n377 B.n100 585
R32 B.n376 B.n375 585
R33 B.n374 B.n101 585
R34 B.n373 B.n372 585
R35 B.n371 B.n102 585
R36 B.n370 B.n369 585
R37 B.n368 B.n103 585
R38 B.n367 B.n366 585
R39 B.n365 B.n104 585
R40 B.n364 B.n363 585
R41 B.n362 B.n105 585
R42 B.n361 B.n360 585
R43 B.n359 B.n106 585
R44 B.n358 B.n357 585
R45 B.n356 B.n107 585
R46 B.n355 B.n354 585
R47 B.n353 B.n108 585
R48 B.n352 B.n351 585
R49 B.n350 B.n109 585
R50 B.n349 B.n348 585
R51 B.n347 B.n110 585
R52 B.n346 B.n345 585
R53 B.n344 B.n111 585
R54 B.n343 B.n342 585
R55 B.n341 B.n112 585
R56 B.n340 B.n339 585
R57 B.n338 B.n113 585
R58 B.n337 B.n336 585
R59 B.n335 B.n114 585
R60 B.n334 B.n333 585
R61 B.n332 B.n115 585
R62 B.n331 B.n330 585
R63 B.n329 B.n116 585
R64 B.n328 B.n327 585
R65 B.n326 B.n117 585
R66 B.n325 B.n324 585
R67 B.n323 B.n118 585
R68 B.n322 B.n321 585
R69 B.n320 B.n119 585
R70 B.n319 B.n318 585
R71 B.n317 B.n120 585
R72 B.n316 B.n315 585
R73 B.n314 B.n121 585
R74 B.n313 B.n312 585
R75 B.n311 B.n122 585
R76 B.n310 B.n309 585
R77 B.n308 B.n123 585
R78 B.n307 B.n306 585
R79 B.n305 B.n124 585
R80 B.n304 B.n303 585
R81 B.n302 B.n125 585
R82 B.n301 B.n300 585
R83 B.n299 B.n298 585
R84 B.n297 B.n129 585
R85 B.n296 B.n295 585
R86 B.n294 B.n130 585
R87 B.n293 B.n292 585
R88 B.n291 B.n131 585
R89 B.n290 B.n289 585
R90 B.n288 B.n132 585
R91 B.n287 B.n286 585
R92 B.n284 B.n133 585
R93 B.n283 B.n282 585
R94 B.n281 B.n136 585
R95 B.n280 B.n279 585
R96 B.n278 B.n137 585
R97 B.n277 B.n276 585
R98 B.n275 B.n138 585
R99 B.n274 B.n273 585
R100 B.n272 B.n139 585
R101 B.n271 B.n270 585
R102 B.n269 B.n140 585
R103 B.n268 B.n267 585
R104 B.n266 B.n141 585
R105 B.n265 B.n264 585
R106 B.n263 B.n142 585
R107 B.n262 B.n261 585
R108 B.n260 B.n143 585
R109 B.n259 B.n258 585
R110 B.n257 B.n144 585
R111 B.n256 B.n255 585
R112 B.n254 B.n145 585
R113 B.n253 B.n252 585
R114 B.n251 B.n146 585
R115 B.n250 B.n249 585
R116 B.n248 B.n147 585
R117 B.n247 B.n246 585
R118 B.n245 B.n148 585
R119 B.n244 B.n243 585
R120 B.n242 B.n149 585
R121 B.n241 B.n240 585
R122 B.n239 B.n150 585
R123 B.n238 B.n237 585
R124 B.n236 B.n151 585
R125 B.n235 B.n234 585
R126 B.n233 B.n152 585
R127 B.n232 B.n231 585
R128 B.n230 B.n153 585
R129 B.n229 B.n228 585
R130 B.n227 B.n154 585
R131 B.n226 B.n225 585
R132 B.n224 B.n155 585
R133 B.n223 B.n222 585
R134 B.n221 B.n156 585
R135 B.n220 B.n219 585
R136 B.n218 B.n157 585
R137 B.n217 B.n216 585
R138 B.n215 B.n158 585
R139 B.n214 B.n213 585
R140 B.n212 B.n159 585
R141 B.n211 B.n210 585
R142 B.n209 B.n160 585
R143 B.n208 B.n207 585
R144 B.n206 B.n161 585
R145 B.n205 B.n204 585
R146 B.n203 B.n162 585
R147 B.n202 B.n201 585
R148 B.n200 B.n163 585
R149 B.n199 B.n198 585
R150 B.n197 B.n164 585
R151 B.n196 B.n195 585
R152 B.n194 B.n165 585
R153 B.n193 B.n192 585
R154 B.n191 B.n166 585
R155 B.n190 B.n189 585
R156 B.n188 B.n167 585
R157 B.n398 B.n93 585
R158 B.n400 B.n399 585
R159 B.n401 B.n92 585
R160 B.n403 B.n402 585
R161 B.n404 B.n91 585
R162 B.n406 B.n405 585
R163 B.n407 B.n90 585
R164 B.n409 B.n408 585
R165 B.n410 B.n89 585
R166 B.n412 B.n411 585
R167 B.n413 B.n88 585
R168 B.n415 B.n414 585
R169 B.n416 B.n87 585
R170 B.n418 B.n417 585
R171 B.n419 B.n86 585
R172 B.n421 B.n420 585
R173 B.n422 B.n85 585
R174 B.n424 B.n423 585
R175 B.n425 B.n84 585
R176 B.n427 B.n426 585
R177 B.n428 B.n83 585
R178 B.n430 B.n429 585
R179 B.n431 B.n82 585
R180 B.n433 B.n432 585
R181 B.n643 B.n642 585
R182 B.n641 B.n8 585
R183 B.n640 B.n639 585
R184 B.n638 B.n9 585
R185 B.n637 B.n636 585
R186 B.n635 B.n10 585
R187 B.n634 B.n633 585
R188 B.n632 B.n11 585
R189 B.n631 B.n630 585
R190 B.n629 B.n12 585
R191 B.n628 B.n627 585
R192 B.n626 B.n13 585
R193 B.n625 B.n624 585
R194 B.n623 B.n14 585
R195 B.n622 B.n621 585
R196 B.n620 B.n15 585
R197 B.n619 B.n618 585
R198 B.n617 B.n16 585
R199 B.n616 B.n615 585
R200 B.n614 B.n17 585
R201 B.n613 B.n612 585
R202 B.n611 B.n18 585
R203 B.n610 B.n609 585
R204 B.n608 B.n19 585
R205 B.n607 B.n606 585
R206 B.n605 B.n20 585
R207 B.n604 B.n603 585
R208 B.n602 B.n21 585
R209 B.n601 B.n600 585
R210 B.n599 B.n22 585
R211 B.n598 B.n597 585
R212 B.n596 B.n23 585
R213 B.n595 B.n594 585
R214 B.n593 B.n24 585
R215 B.n592 B.n591 585
R216 B.n590 B.n25 585
R217 B.n589 B.n588 585
R218 B.n587 B.n26 585
R219 B.n586 B.n585 585
R220 B.n584 B.n27 585
R221 B.n583 B.n582 585
R222 B.n581 B.n28 585
R223 B.n580 B.n579 585
R224 B.n578 B.n29 585
R225 B.n577 B.n576 585
R226 B.n575 B.n30 585
R227 B.n574 B.n573 585
R228 B.n572 B.n31 585
R229 B.n571 B.n570 585
R230 B.n569 B.n32 585
R231 B.n568 B.n567 585
R232 B.n566 B.n33 585
R233 B.n565 B.n564 585
R234 B.n563 B.n34 585
R235 B.n562 B.n561 585
R236 B.n560 B.n35 585
R237 B.n559 B.n558 585
R238 B.n557 B.n36 585
R239 B.n556 B.n555 585
R240 B.n554 B.n37 585
R241 B.n553 B.n552 585
R242 B.n551 B.n38 585
R243 B.n550 B.n549 585
R244 B.n548 B.n39 585
R245 B.n547 B.n546 585
R246 B.n545 B.n544 585
R247 B.n543 B.n43 585
R248 B.n542 B.n541 585
R249 B.n540 B.n44 585
R250 B.n539 B.n538 585
R251 B.n537 B.n45 585
R252 B.n536 B.n535 585
R253 B.n534 B.n46 585
R254 B.n533 B.n532 585
R255 B.n530 B.n47 585
R256 B.n529 B.n528 585
R257 B.n527 B.n50 585
R258 B.n526 B.n525 585
R259 B.n524 B.n51 585
R260 B.n523 B.n522 585
R261 B.n521 B.n52 585
R262 B.n520 B.n519 585
R263 B.n518 B.n53 585
R264 B.n517 B.n516 585
R265 B.n515 B.n54 585
R266 B.n514 B.n513 585
R267 B.n512 B.n55 585
R268 B.n511 B.n510 585
R269 B.n509 B.n56 585
R270 B.n508 B.n507 585
R271 B.n506 B.n57 585
R272 B.n505 B.n504 585
R273 B.n503 B.n58 585
R274 B.n502 B.n501 585
R275 B.n500 B.n59 585
R276 B.n499 B.n498 585
R277 B.n497 B.n60 585
R278 B.n496 B.n495 585
R279 B.n494 B.n61 585
R280 B.n493 B.n492 585
R281 B.n491 B.n62 585
R282 B.n490 B.n489 585
R283 B.n488 B.n63 585
R284 B.n487 B.n486 585
R285 B.n485 B.n64 585
R286 B.n484 B.n483 585
R287 B.n482 B.n65 585
R288 B.n481 B.n480 585
R289 B.n479 B.n66 585
R290 B.n478 B.n477 585
R291 B.n476 B.n67 585
R292 B.n475 B.n474 585
R293 B.n473 B.n68 585
R294 B.n472 B.n471 585
R295 B.n470 B.n69 585
R296 B.n469 B.n468 585
R297 B.n467 B.n70 585
R298 B.n466 B.n465 585
R299 B.n464 B.n71 585
R300 B.n463 B.n462 585
R301 B.n461 B.n72 585
R302 B.n460 B.n459 585
R303 B.n458 B.n73 585
R304 B.n457 B.n456 585
R305 B.n455 B.n74 585
R306 B.n454 B.n453 585
R307 B.n452 B.n75 585
R308 B.n451 B.n450 585
R309 B.n449 B.n76 585
R310 B.n448 B.n447 585
R311 B.n446 B.n77 585
R312 B.n445 B.n444 585
R313 B.n443 B.n78 585
R314 B.n442 B.n441 585
R315 B.n440 B.n79 585
R316 B.n439 B.n438 585
R317 B.n437 B.n80 585
R318 B.n436 B.n435 585
R319 B.n434 B.n81 585
R320 B.n644 B.n7 585
R321 B.n646 B.n645 585
R322 B.n647 B.n6 585
R323 B.n649 B.n648 585
R324 B.n650 B.n5 585
R325 B.n652 B.n651 585
R326 B.n653 B.n4 585
R327 B.n655 B.n654 585
R328 B.n656 B.n3 585
R329 B.n658 B.n657 585
R330 B.n659 B.n0 585
R331 B.n2 B.n1 585
R332 B.n173 B.n172 585
R333 B.n175 B.n174 585
R334 B.n176 B.n171 585
R335 B.n178 B.n177 585
R336 B.n179 B.n170 585
R337 B.n181 B.n180 585
R338 B.n182 B.n169 585
R339 B.n184 B.n183 585
R340 B.n185 B.n168 585
R341 B.n187 B.n186 585
R342 B.n186 B.n167 550.159
R343 B.n396 B.n93 550.159
R344 B.n432 B.n81 550.159
R345 B.n642 B.n7 550.159
R346 B.n661 B.n660 256.663
R347 B.n660 B.n659 235.042
R348 B.n660 B.n2 235.042
R349 B.n190 B.n167 163.367
R350 B.n191 B.n190 163.367
R351 B.n192 B.n191 163.367
R352 B.n192 B.n165 163.367
R353 B.n196 B.n165 163.367
R354 B.n197 B.n196 163.367
R355 B.n198 B.n197 163.367
R356 B.n198 B.n163 163.367
R357 B.n202 B.n163 163.367
R358 B.n203 B.n202 163.367
R359 B.n204 B.n203 163.367
R360 B.n204 B.n161 163.367
R361 B.n208 B.n161 163.367
R362 B.n209 B.n208 163.367
R363 B.n210 B.n209 163.367
R364 B.n210 B.n159 163.367
R365 B.n214 B.n159 163.367
R366 B.n215 B.n214 163.367
R367 B.n216 B.n215 163.367
R368 B.n216 B.n157 163.367
R369 B.n220 B.n157 163.367
R370 B.n221 B.n220 163.367
R371 B.n222 B.n221 163.367
R372 B.n222 B.n155 163.367
R373 B.n226 B.n155 163.367
R374 B.n227 B.n226 163.367
R375 B.n228 B.n227 163.367
R376 B.n228 B.n153 163.367
R377 B.n232 B.n153 163.367
R378 B.n233 B.n232 163.367
R379 B.n234 B.n233 163.367
R380 B.n234 B.n151 163.367
R381 B.n238 B.n151 163.367
R382 B.n239 B.n238 163.367
R383 B.n240 B.n239 163.367
R384 B.n240 B.n149 163.367
R385 B.n244 B.n149 163.367
R386 B.n245 B.n244 163.367
R387 B.n246 B.n245 163.367
R388 B.n246 B.n147 163.367
R389 B.n250 B.n147 163.367
R390 B.n251 B.n250 163.367
R391 B.n252 B.n251 163.367
R392 B.n252 B.n145 163.367
R393 B.n256 B.n145 163.367
R394 B.n257 B.n256 163.367
R395 B.n258 B.n257 163.367
R396 B.n258 B.n143 163.367
R397 B.n262 B.n143 163.367
R398 B.n263 B.n262 163.367
R399 B.n264 B.n263 163.367
R400 B.n264 B.n141 163.367
R401 B.n268 B.n141 163.367
R402 B.n269 B.n268 163.367
R403 B.n270 B.n269 163.367
R404 B.n270 B.n139 163.367
R405 B.n274 B.n139 163.367
R406 B.n275 B.n274 163.367
R407 B.n276 B.n275 163.367
R408 B.n276 B.n137 163.367
R409 B.n280 B.n137 163.367
R410 B.n281 B.n280 163.367
R411 B.n282 B.n281 163.367
R412 B.n282 B.n133 163.367
R413 B.n287 B.n133 163.367
R414 B.n288 B.n287 163.367
R415 B.n289 B.n288 163.367
R416 B.n289 B.n131 163.367
R417 B.n293 B.n131 163.367
R418 B.n294 B.n293 163.367
R419 B.n295 B.n294 163.367
R420 B.n295 B.n129 163.367
R421 B.n299 B.n129 163.367
R422 B.n300 B.n299 163.367
R423 B.n300 B.n125 163.367
R424 B.n304 B.n125 163.367
R425 B.n305 B.n304 163.367
R426 B.n306 B.n305 163.367
R427 B.n306 B.n123 163.367
R428 B.n310 B.n123 163.367
R429 B.n311 B.n310 163.367
R430 B.n312 B.n311 163.367
R431 B.n312 B.n121 163.367
R432 B.n316 B.n121 163.367
R433 B.n317 B.n316 163.367
R434 B.n318 B.n317 163.367
R435 B.n318 B.n119 163.367
R436 B.n322 B.n119 163.367
R437 B.n323 B.n322 163.367
R438 B.n324 B.n323 163.367
R439 B.n324 B.n117 163.367
R440 B.n328 B.n117 163.367
R441 B.n329 B.n328 163.367
R442 B.n330 B.n329 163.367
R443 B.n330 B.n115 163.367
R444 B.n334 B.n115 163.367
R445 B.n335 B.n334 163.367
R446 B.n336 B.n335 163.367
R447 B.n336 B.n113 163.367
R448 B.n340 B.n113 163.367
R449 B.n341 B.n340 163.367
R450 B.n342 B.n341 163.367
R451 B.n342 B.n111 163.367
R452 B.n346 B.n111 163.367
R453 B.n347 B.n346 163.367
R454 B.n348 B.n347 163.367
R455 B.n348 B.n109 163.367
R456 B.n352 B.n109 163.367
R457 B.n353 B.n352 163.367
R458 B.n354 B.n353 163.367
R459 B.n354 B.n107 163.367
R460 B.n358 B.n107 163.367
R461 B.n359 B.n358 163.367
R462 B.n360 B.n359 163.367
R463 B.n360 B.n105 163.367
R464 B.n364 B.n105 163.367
R465 B.n365 B.n364 163.367
R466 B.n366 B.n365 163.367
R467 B.n366 B.n103 163.367
R468 B.n370 B.n103 163.367
R469 B.n371 B.n370 163.367
R470 B.n372 B.n371 163.367
R471 B.n372 B.n101 163.367
R472 B.n376 B.n101 163.367
R473 B.n377 B.n376 163.367
R474 B.n378 B.n377 163.367
R475 B.n378 B.n99 163.367
R476 B.n382 B.n99 163.367
R477 B.n383 B.n382 163.367
R478 B.n384 B.n383 163.367
R479 B.n384 B.n97 163.367
R480 B.n388 B.n97 163.367
R481 B.n389 B.n388 163.367
R482 B.n390 B.n389 163.367
R483 B.n390 B.n95 163.367
R484 B.n394 B.n95 163.367
R485 B.n395 B.n394 163.367
R486 B.n396 B.n395 163.367
R487 B.n432 B.n431 163.367
R488 B.n431 B.n430 163.367
R489 B.n430 B.n83 163.367
R490 B.n426 B.n83 163.367
R491 B.n426 B.n425 163.367
R492 B.n425 B.n424 163.367
R493 B.n424 B.n85 163.367
R494 B.n420 B.n85 163.367
R495 B.n420 B.n419 163.367
R496 B.n419 B.n418 163.367
R497 B.n418 B.n87 163.367
R498 B.n414 B.n87 163.367
R499 B.n414 B.n413 163.367
R500 B.n413 B.n412 163.367
R501 B.n412 B.n89 163.367
R502 B.n408 B.n89 163.367
R503 B.n408 B.n407 163.367
R504 B.n407 B.n406 163.367
R505 B.n406 B.n91 163.367
R506 B.n402 B.n91 163.367
R507 B.n402 B.n401 163.367
R508 B.n401 B.n400 163.367
R509 B.n400 B.n93 163.367
R510 B.n642 B.n641 163.367
R511 B.n641 B.n640 163.367
R512 B.n640 B.n9 163.367
R513 B.n636 B.n9 163.367
R514 B.n636 B.n635 163.367
R515 B.n635 B.n634 163.367
R516 B.n634 B.n11 163.367
R517 B.n630 B.n11 163.367
R518 B.n630 B.n629 163.367
R519 B.n629 B.n628 163.367
R520 B.n628 B.n13 163.367
R521 B.n624 B.n13 163.367
R522 B.n624 B.n623 163.367
R523 B.n623 B.n622 163.367
R524 B.n622 B.n15 163.367
R525 B.n618 B.n15 163.367
R526 B.n618 B.n617 163.367
R527 B.n617 B.n616 163.367
R528 B.n616 B.n17 163.367
R529 B.n612 B.n17 163.367
R530 B.n612 B.n611 163.367
R531 B.n611 B.n610 163.367
R532 B.n610 B.n19 163.367
R533 B.n606 B.n19 163.367
R534 B.n606 B.n605 163.367
R535 B.n605 B.n604 163.367
R536 B.n604 B.n21 163.367
R537 B.n600 B.n21 163.367
R538 B.n600 B.n599 163.367
R539 B.n599 B.n598 163.367
R540 B.n598 B.n23 163.367
R541 B.n594 B.n23 163.367
R542 B.n594 B.n593 163.367
R543 B.n593 B.n592 163.367
R544 B.n592 B.n25 163.367
R545 B.n588 B.n25 163.367
R546 B.n588 B.n587 163.367
R547 B.n587 B.n586 163.367
R548 B.n586 B.n27 163.367
R549 B.n582 B.n27 163.367
R550 B.n582 B.n581 163.367
R551 B.n581 B.n580 163.367
R552 B.n580 B.n29 163.367
R553 B.n576 B.n29 163.367
R554 B.n576 B.n575 163.367
R555 B.n575 B.n574 163.367
R556 B.n574 B.n31 163.367
R557 B.n570 B.n31 163.367
R558 B.n570 B.n569 163.367
R559 B.n569 B.n568 163.367
R560 B.n568 B.n33 163.367
R561 B.n564 B.n33 163.367
R562 B.n564 B.n563 163.367
R563 B.n563 B.n562 163.367
R564 B.n562 B.n35 163.367
R565 B.n558 B.n35 163.367
R566 B.n558 B.n557 163.367
R567 B.n557 B.n556 163.367
R568 B.n556 B.n37 163.367
R569 B.n552 B.n37 163.367
R570 B.n552 B.n551 163.367
R571 B.n551 B.n550 163.367
R572 B.n550 B.n39 163.367
R573 B.n546 B.n39 163.367
R574 B.n546 B.n545 163.367
R575 B.n545 B.n43 163.367
R576 B.n541 B.n43 163.367
R577 B.n541 B.n540 163.367
R578 B.n540 B.n539 163.367
R579 B.n539 B.n45 163.367
R580 B.n535 B.n45 163.367
R581 B.n535 B.n534 163.367
R582 B.n534 B.n533 163.367
R583 B.n533 B.n47 163.367
R584 B.n528 B.n47 163.367
R585 B.n528 B.n527 163.367
R586 B.n527 B.n526 163.367
R587 B.n526 B.n51 163.367
R588 B.n522 B.n51 163.367
R589 B.n522 B.n521 163.367
R590 B.n521 B.n520 163.367
R591 B.n520 B.n53 163.367
R592 B.n516 B.n53 163.367
R593 B.n516 B.n515 163.367
R594 B.n515 B.n514 163.367
R595 B.n514 B.n55 163.367
R596 B.n510 B.n55 163.367
R597 B.n510 B.n509 163.367
R598 B.n509 B.n508 163.367
R599 B.n508 B.n57 163.367
R600 B.n504 B.n57 163.367
R601 B.n504 B.n503 163.367
R602 B.n503 B.n502 163.367
R603 B.n502 B.n59 163.367
R604 B.n498 B.n59 163.367
R605 B.n498 B.n497 163.367
R606 B.n497 B.n496 163.367
R607 B.n496 B.n61 163.367
R608 B.n492 B.n61 163.367
R609 B.n492 B.n491 163.367
R610 B.n491 B.n490 163.367
R611 B.n490 B.n63 163.367
R612 B.n486 B.n63 163.367
R613 B.n486 B.n485 163.367
R614 B.n485 B.n484 163.367
R615 B.n484 B.n65 163.367
R616 B.n480 B.n65 163.367
R617 B.n480 B.n479 163.367
R618 B.n479 B.n478 163.367
R619 B.n478 B.n67 163.367
R620 B.n474 B.n67 163.367
R621 B.n474 B.n473 163.367
R622 B.n473 B.n472 163.367
R623 B.n472 B.n69 163.367
R624 B.n468 B.n69 163.367
R625 B.n468 B.n467 163.367
R626 B.n467 B.n466 163.367
R627 B.n466 B.n71 163.367
R628 B.n462 B.n71 163.367
R629 B.n462 B.n461 163.367
R630 B.n461 B.n460 163.367
R631 B.n460 B.n73 163.367
R632 B.n456 B.n73 163.367
R633 B.n456 B.n455 163.367
R634 B.n455 B.n454 163.367
R635 B.n454 B.n75 163.367
R636 B.n450 B.n75 163.367
R637 B.n450 B.n449 163.367
R638 B.n449 B.n448 163.367
R639 B.n448 B.n77 163.367
R640 B.n444 B.n77 163.367
R641 B.n444 B.n443 163.367
R642 B.n443 B.n442 163.367
R643 B.n442 B.n79 163.367
R644 B.n438 B.n79 163.367
R645 B.n438 B.n437 163.367
R646 B.n437 B.n436 163.367
R647 B.n436 B.n81 163.367
R648 B.n646 B.n7 163.367
R649 B.n647 B.n646 163.367
R650 B.n648 B.n647 163.367
R651 B.n648 B.n5 163.367
R652 B.n652 B.n5 163.367
R653 B.n653 B.n652 163.367
R654 B.n654 B.n653 163.367
R655 B.n654 B.n3 163.367
R656 B.n658 B.n3 163.367
R657 B.n659 B.n658 163.367
R658 B.n173 B.n2 163.367
R659 B.n174 B.n173 163.367
R660 B.n174 B.n171 163.367
R661 B.n178 B.n171 163.367
R662 B.n179 B.n178 163.367
R663 B.n180 B.n179 163.367
R664 B.n180 B.n169 163.367
R665 B.n184 B.n169 163.367
R666 B.n185 B.n184 163.367
R667 B.n186 B.n185 163.367
R668 B.n126 B.t10 120.776
R669 B.n48 B.t8 120.776
R670 B.n134 B.t4 120.751
R671 B.n40 B.t2 120.751
R672 B.n127 B.t11 108.945
R673 B.n49 B.t7 108.945
R674 B.n135 B.t5 108.919
R675 B.n41 B.t1 108.919
R676 B.n285 B.n135 59.5399
R677 B.n128 B.n127 59.5399
R678 B.n531 B.n49 59.5399
R679 B.n42 B.n41 59.5399
R680 B.n398 B.n397 35.7468
R681 B.n644 B.n643 35.7468
R682 B.n434 B.n433 35.7468
R683 B.n188 B.n187 35.7468
R684 B B.n661 18.0485
R685 B.n135 B.n134 11.8308
R686 B.n127 B.n126 11.8308
R687 B.n49 B.n48 11.8308
R688 B.n41 B.n40 11.8308
R689 B.n645 B.n644 10.6151
R690 B.n645 B.n6 10.6151
R691 B.n649 B.n6 10.6151
R692 B.n650 B.n649 10.6151
R693 B.n651 B.n650 10.6151
R694 B.n651 B.n4 10.6151
R695 B.n655 B.n4 10.6151
R696 B.n656 B.n655 10.6151
R697 B.n657 B.n656 10.6151
R698 B.n657 B.n0 10.6151
R699 B.n643 B.n8 10.6151
R700 B.n639 B.n8 10.6151
R701 B.n639 B.n638 10.6151
R702 B.n638 B.n637 10.6151
R703 B.n637 B.n10 10.6151
R704 B.n633 B.n10 10.6151
R705 B.n633 B.n632 10.6151
R706 B.n632 B.n631 10.6151
R707 B.n631 B.n12 10.6151
R708 B.n627 B.n12 10.6151
R709 B.n627 B.n626 10.6151
R710 B.n626 B.n625 10.6151
R711 B.n625 B.n14 10.6151
R712 B.n621 B.n14 10.6151
R713 B.n621 B.n620 10.6151
R714 B.n620 B.n619 10.6151
R715 B.n619 B.n16 10.6151
R716 B.n615 B.n16 10.6151
R717 B.n615 B.n614 10.6151
R718 B.n614 B.n613 10.6151
R719 B.n613 B.n18 10.6151
R720 B.n609 B.n18 10.6151
R721 B.n609 B.n608 10.6151
R722 B.n608 B.n607 10.6151
R723 B.n607 B.n20 10.6151
R724 B.n603 B.n20 10.6151
R725 B.n603 B.n602 10.6151
R726 B.n602 B.n601 10.6151
R727 B.n601 B.n22 10.6151
R728 B.n597 B.n22 10.6151
R729 B.n597 B.n596 10.6151
R730 B.n596 B.n595 10.6151
R731 B.n595 B.n24 10.6151
R732 B.n591 B.n24 10.6151
R733 B.n591 B.n590 10.6151
R734 B.n590 B.n589 10.6151
R735 B.n589 B.n26 10.6151
R736 B.n585 B.n26 10.6151
R737 B.n585 B.n584 10.6151
R738 B.n584 B.n583 10.6151
R739 B.n583 B.n28 10.6151
R740 B.n579 B.n28 10.6151
R741 B.n579 B.n578 10.6151
R742 B.n578 B.n577 10.6151
R743 B.n577 B.n30 10.6151
R744 B.n573 B.n30 10.6151
R745 B.n573 B.n572 10.6151
R746 B.n572 B.n571 10.6151
R747 B.n571 B.n32 10.6151
R748 B.n567 B.n32 10.6151
R749 B.n567 B.n566 10.6151
R750 B.n566 B.n565 10.6151
R751 B.n565 B.n34 10.6151
R752 B.n561 B.n34 10.6151
R753 B.n561 B.n560 10.6151
R754 B.n560 B.n559 10.6151
R755 B.n559 B.n36 10.6151
R756 B.n555 B.n36 10.6151
R757 B.n555 B.n554 10.6151
R758 B.n554 B.n553 10.6151
R759 B.n553 B.n38 10.6151
R760 B.n549 B.n38 10.6151
R761 B.n549 B.n548 10.6151
R762 B.n548 B.n547 10.6151
R763 B.n544 B.n543 10.6151
R764 B.n543 B.n542 10.6151
R765 B.n542 B.n44 10.6151
R766 B.n538 B.n44 10.6151
R767 B.n538 B.n537 10.6151
R768 B.n537 B.n536 10.6151
R769 B.n536 B.n46 10.6151
R770 B.n532 B.n46 10.6151
R771 B.n530 B.n529 10.6151
R772 B.n529 B.n50 10.6151
R773 B.n525 B.n50 10.6151
R774 B.n525 B.n524 10.6151
R775 B.n524 B.n523 10.6151
R776 B.n523 B.n52 10.6151
R777 B.n519 B.n52 10.6151
R778 B.n519 B.n518 10.6151
R779 B.n518 B.n517 10.6151
R780 B.n517 B.n54 10.6151
R781 B.n513 B.n54 10.6151
R782 B.n513 B.n512 10.6151
R783 B.n512 B.n511 10.6151
R784 B.n511 B.n56 10.6151
R785 B.n507 B.n56 10.6151
R786 B.n507 B.n506 10.6151
R787 B.n506 B.n505 10.6151
R788 B.n505 B.n58 10.6151
R789 B.n501 B.n58 10.6151
R790 B.n501 B.n500 10.6151
R791 B.n500 B.n499 10.6151
R792 B.n499 B.n60 10.6151
R793 B.n495 B.n60 10.6151
R794 B.n495 B.n494 10.6151
R795 B.n494 B.n493 10.6151
R796 B.n493 B.n62 10.6151
R797 B.n489 B.n62 10.6151
R798 B.n489 B.n488 10.6151
R799 B.n488 B.n487 10.6151
R800 B.n487 B.n64 10.6151
R801 B.n483 B.n64 10.6151
R802 B.n483 B.n482 10.6151
R803 B.n482 B.n481 10.6151
R804 B.n481 B.n66 10.6151
R805 B.n477 B.n66 10.6151
R806 B.n477 B.n476 10.6151
R807 B.n476 B.n475 10.6151
R808 B.n475 B.n68 10.6151
R809 B.n471 B.n68 10.6151
R810 B.n471 B.n470 10.6151
R811 B.n470 B.n469 10.6151
R812 B.n469 B.n70 10.6151
R813 B.n465 B.n70 10.6151
R814 B.n465 B.n464 10.6151
R815 B.n464 B.n463 10.6151
R816 B.n463 B.n72 10.6151
R817 B.n459 B.n72 10.6151
R818 B.n459 B.n458 10.6151
R819 B.n458 B.n457 10.6151
R820 B.n457 B.n74 10.6151
R821 B.n453 B.n74 10.6151
R822 B.n453 B.n452 10.6151
R823 B.n452 B.n451 10.6151
R824 B.n451 B.n76 10.6151
R825 B.n447 B.n76 10.6151
R826 B.n447 B.n446 10.6151
R827 B.n446 B.n445 10.6151
R828 B.n445 B.n78 10.6151
R829 B.n441 B.n78 10.6151
R830 B.n441 B.n440 10.6151
R831 B.n440 B.n439 10.6151
R832 B.n439 B.n80 10.6151
R833 B.n435 B.n80 10.6151
R834 B.n435 B.n434 10.6151
R835 B.n433 B.n82 10.6151
R836 B.n429 B.n82 10.6151
R837 B.n429 B.n428 10.6151
R838 B.n428 B.n427 10.6151
R839 B.n427 B.n84 10.6151
R840 B.n423 B.n84 10.6151
R841 B.n423 B.n422 10.6151
R842 B.n422 B.n421 10.6151
R843 B.n421 B.n86 10.6151
R844 B.n417 B.n86 10.6151
R845 B.n417 B.n416 10.6151
R846 B.n416 B.n415 10.6151
R847 B.n415 B.n88 10.6151
R848 B.n411 B.n88 10.6151
R849 B.n411 B.n410 10.6151
R850 B.n410 B.n409 10.6151
R851 B.n409 B.n90 10.6151
R852 B.n405 B.n90 10.6151
R853 B.n405 B.n404 10.6151
R854 B.n404 B.n403 10.6151
R855 B.n403 B.n92 10.6151
R856 B.n399 B.n92 10.6151
R857 B.n399 B.n398 10.6151
R858 B.n172 B.n1 10.6151
R859 B.n175 B.n172 10.6151
R860 B.n176 B.n175 10.6151
R861 B.n177 B.n176 10.6151
R862 B.n177 B.n170 10.6151
R863 B.n181 B.n170 10.6151
R864 B.n182 B.n181 10.6151
R865 B.n183 B.n182 10.6151
R866 B.n183 B.n168 10.6151
R867 B.n187 B.n168 10.6151
R868 B.n189 B.n188 10.6151
R869 B.n189 B.n166 10.6151
R870 B.n193 B.n166 10.6151
R871 B.n194 B.n193 10.6151
R872 B.n195 B.n194 10.6151
R873 B.n195 B.n164 10.6151
R874 B.n199 B.n164 10.6151
R875 B.n200 B.n199 10.6151
R876 B.n201 B.n200 10.6151
R877 B.n201 B.n162 10.6151
R878 B.n205 B.n162 10.6151
R879 B.n206 B.n205 10.6151
R880 B.n207 B.n206 10.6151
R881 B.n207 B.n160 10.6151
R882 B.n211 B.n160 10.6151
R883 B.n212 B.n211 10.6151
R884 B.n213 B.n212 10.6151
R885 B.n213 B.n158 10.6151
R886 B.n217 B.n158 10.6151
R887 B.n218 B.n217 10.6151
R888 B.n219 B.n218 10.6151
R889 B.n219 B.n156 10.6151
R890 B.n223 B.n156 10.6151
R891 B.n224 B.n223 10.6151
R892 B.n225 B.n224 10.6151
R893 B.n225 B.n154 10.6151
R894 B.n229 B.n154 10.6151
R895 B.n230 B.n229 10.6151
R896 B.n231 B.n230 10.6151
R897 B.n231 B.n152 10.6151
R898 B.n235 B.n152 10.6151
R899 B.n236 B.n235 10.6151
R900 B.n237 B.n236 10.6151
R901 B.n237 B.n150 10.6151
R902 B.n241 B.n150 10.6151
R903 B.n242 B.n241 10.6151
R904 B.n243 B.n242 10.6151
R905 B.n243 B.n148 10.6151
R906 B.n247 B.n148 10.6151
R907 B.n248 B.n247 10.6151
R908 B.n249 B.n248 10.6151
R909 B.n249 B.n146 10.6151
R910 B.n253 B.n146 10.6151
R911 B.n254 B.n253 10.6151
R912 B.n255 B.n254 10.6151
R913 B.n255 B.n144 10.6151
R914 B.n259 B.n144 10.6151
R915 B.n260 B.n259 10.6151
R916 B.n261 B.n260 10.6151
R917 B.n261 B.n142 10.6151
R918 B.n265 B.n142 10.6151
R919 B.n266 B.n265 10.6151
R920 B.n267 B.n266 10.6151
R921 B.n267 B.n140 10.6151
R922 B.n271 B.n140 10.6151
R923 B.n272 B.n271 10.6151
R924 B.n273 B.n272 10.6151
R925 B.n273 B.n138 10.6151
R926 B.n277 B.n138 10.6151
R927 B.n278 B.n277 10.6151
R928 B.n279 B.n278 10.6151
R929 B.n279 B.n136 10.6151
R930 B.n283 B.n136 10.6151
R931 B.n284 B.n283 10.6151
R932 B.n286 B.n132 10.6151
R933 B.n290 B.n132 10.6151
R934 B.n291 B.n290 10.6151
R935 B.n292 B.n291 10.6151
R936 B.n292 B.n130 10.6151
R937 B.n296 B.n130 10.6151
R938 B.n297 B.n296 10.6151
R939 B.n298 B.n297 10.6151
R940 B.n302 B.n301 10.6151
R941 B.n303 B.n302 10.6151
R942 B.n303 B.n124 10.6151
R943 B.n307 B.n124 10.6151
R944 B.n308 B.n307 10.6151
R945 B.n309 B.n308 10.6151
R946 B.n309 B.n122 10.6151
R947 B.n313 B.n122 10.6151
R948 B.n314 B.n313 10.6151
R949 B.n315 B.n314 10.6151
R950 B.n315 B.n120 10.6151
R951 B.n319 B.n120 10.6151
R952 B.n320 B.n319 10.6151
R953 B.n321 B.n320 10.6151
R954 B.n321 B.n118 10.6151
R955 B.n325 B.n118 10.6151
R956 B.n326 B.n325 10.6151
R957 B.n327 B.n326 10.6151
R958 B.n327 B.n116 10.6151
R959 B.n331 B.n116 10.6151
R960 B.n332 B.n331 10.6151
R961 B.n333 B.n332 10.6151
R962 B.n333 B.n114 10.6151
R963 B.n337 B.n114 10.6151
R964 B.n338 B.n337 10.6151
R965 B.n339 B.n338 10.6151
R966 B.n339 B.n112 10.6151
R967 B.n343 B.n112 10.6151
R968 B.n344 B.n343 10.6151
R969 B.n345 B.n344 10.6151
R970 B.n345 B.n110 10.6151
R971 B.n349 B.n110 10.6151
R972 B.n350 B.n349 10.6151
R973 B.n351 B.n350 10.6151
R974 B.n351 B.n108 10.6151
R975 B.n355 B.n108 10.6151
R976 B.n356 B.n355 10.6151
R977 B.n357 B.n356 10.6151
R978 B.n357 B.n106 10.6151
R979 B.n361 B.n106 10.6151
R980 B.n362 B.n361 10.6151
R981 B.n363 B.n362 10.6151
R982 B.n363 B.n104 10.6151
R983 B.n367 B.n104 10.6151
R984 B.n368 B.n367 10.6151
R985 B.n369 B.n368 10.6151
R986 B.n369 B.n102 10.6151
R987 B.n373 B.n102 10.6151
R988 B.n374 B.n373 10.6151
R989 B.n375 B.n374 10.6151
R990 B.n375 B.n100 10.6151
R991 B.n379 B.n100 10.6151
R992 B.n380 B.n379 10.6151
R993 B.n381 B.n380 10.6151
R994 B.n381 B.n98 10.6151
R995 B.n385 B.n98 10.6151
R996 B.n386 B.n385 10.6151
R997 B.n387 B.n386 10.6151
R998 B.n387 B.n96 10.6151
R999 B.n391 B.n96 10.6151
R1000 B.n392 B.n391 10.6151
R1001 B.n393 B.n392 10.6151
R1002 B.n393 B.n94 10.6151
R1003 B.n397 B.n94 10.6151
R1004 B.n661 B.n0 8.11757
R1005 B.n661 B.n1 8.11757
R1006 B.n544 B.n42 7.18099
R1007 B.n532 B.n531 7.18099
R1008 B.n286 B.n285 7.18099
R1009 B.n298 B.n128 7.18099
R1010 B.n547 B.n42 3.43465
R1011 B.n531 B.n530 3.43465
R1012 B.n285 B.n284 3.43465
R1013 B.n301 B.n128 3.43465
R1014 VP.n0 VP.t0 2052.87
R1015 VP.n0 VP.t1 2008.39
R1016 VP VP.n0 0.0516364
R1017 VDD1 VDD1.t0 115.556
R1018 VDD1 VDD1.t1 73.2324
C0 VDD1 VTAIL 11.0158f
C1 VTAIL VDD2 11.0392f
C2 B VTAIL 3.76246f
C3 VTAIL VN 1.22153f
C4 VDD1 VDD2 0.427852f
C5 w_n1214_n4946# VTAIL 4.39582f
C6 B VDD1 1.88655f
C7 B VDD2 1.89834f
C8 VDD1 VN 0.14839f
C9 VDD2 VN 2.18803f
C10 B VN 0.746858f
C11 VDD1 w_n1214_n4946# 2.1215f
C12 w_n1214_n4946# VDD2 2.12201f
C13 B w_n1214_n4946# 8.532559f
C14 w_n1214_n4946# VN 1.65422f
C15 VTAIL VP 1.23673f
C16 VDD1 VP 2.27031f
C17 VDD2 VP 0.239024f
C18 B VP 0.983562f
C19 VP VN 5.83194f
C20 w_n1214_n4946# VP 1.80386f
C21 VDD2 VSUBS 1.000367f
C22 VDD1 VSUBS 6.08157f
C23 VTAIL VSUBS 0.21987f
C24 VN VSUBS 7.78189f
C25 VP VSUBS 1.285757f
C26 B VSUBS 2.855293f
C27 w_n1214_n4946# VSUBS 73.3207f
C28 VDD1.t1 VSUBS 4.7303f
C29 VDD1.t0 VSUBS 5.67747f
C30 VP.t0 VSUBS 1.04242f
C31 VP.t1 VSUBS 0.976353f
C32 VP.n0 VSUBS 6.07399f
C33 B.n0 VSUBS 0.00643f
C34 B.n1 VSUBS 0.00643f
C35 B.n2 VSUBS 0.009509f
C36 B.n3 VSUBS 0.007287f
C37 B.n4 VSUBS 0.007287f
C38 B.n5 VSUBS 0.007287f
C39 B.n6 VSUBS 0.007287f
C40 B.n7 VSUBS 0.017678f
C41 B.n8 VSUBS 0.007287f
C42 B.n9 VSUBS 0.007287f
C43 B.n10 VSUBS 0.007287f
C44 B.n11 VSUBS 0.007287f
C45 B.n12 VSUBS 0.007287f
C46 B.n13 VSUBS 0.007287f
C47 B.n14 VSUBS 0.007287f
C48 B.n15 VSUBS 0.007287f
C49 B.n16 VSUBS 0.007287f
C50 B.n17 VSUBS 0.007287f
C51 B.n18 VSUBS 0.007287f
C52 B.n19 VSUBS 0.007287f
C53 B.n20 VSUBS 0.007287f
C54 B.n21 VSUBS 0.007287f
C55 B.n22 VSUBS 0.007287f
C56 B.n23 VSUBS 0.007287f
C57 B.n24 VSUBS 0.007287f
C58 B.n25 VSUBS 0.007287f
C59 B.n26 VSUBS 0.007287f
C60 B.n27 VSUBS 0.007287f
C61 B.n28 VSUBS 0.007287f
C62 B.n29 VSUBS 0.007287f
C63 B.n30 VSUBS 0.007287f
C64 B.n31 VSUBS 0.007287f
C65 B.n32 VSUBS 0.007287f
C66 B.n33 VSUBS 0.007287f
C67 B.n34 VSUBS 0.007287f
C68 B.n35 VSUBS 0.007287f
C69 B.n36 VSUBS 0.007287f
C70 B.n37 VSUBS 0.007287f
C71 B.n38 VSUBS 0.007287f
C72 B.n39 VSUBS 0.007287f
C73 B.t1 VSUBS 0.702896f
C74 B.t2 VSUBS 0.708258f
C75 B.t0 VSUBS 0.22356f
C76 B.n40 VSUBS 0.127594f
C77 B.n41 VSUBS 0.065129f
C78 B.n42 VSUBS 0.016883f
C79 B.n43 VSUBS 0.007287f
C80 B.n44 VSUBS 0.007287f
C81 B.n45 VSUBS 0.007287f
C82 B.n46 VSUBS 0.007287f
C83 B.n47 VSUBS 0.007287f
C84 B.t7 VSUBS 0.702866f
C85 B.t8 VSUBS 0.70823f
C86 B.t6 VSUBS 0.22356f
C87 B.n48 VSUBS 0.127622f
C88 B.n49 VSUBS 0.065159f
C89 B.n50 VSUBS 0.007287f
C90 B.n51 VSUBS 0.007287f
C91 B.n52 VSUBS 0.007287f
C92 B.n53 VSUBS 0.007287f
C93 B.n54 VSUBS 0.007287f
C94 B.n55 VSUBS 0.007287f
C95 B.n56 VSUBS 0.007287f
C96 B.n57 VSUBS 0.007287f
C97 B.n58 VSUBS 0.007287f
C98 B.n59 VSUBS 0.007287f
C99 B.n60 VSUBS 0.007287f
C100 B.n61 VSUBS 0.007287f
C101 B.n62 VSUBS 0.007287f
C102 B.n63 VSUBS 0.007287f
C103 B.n64 VSUBS 0.007287f
C104 B.n65 VSUBS 0.007287f
C105 B.n66 VSUBS 0.007287f
C106 B.n67 VSUBS 0.007287f
C107 B.n68 VSUBS 0.007287f
C108 B.n69 VSUBS 0.007287f
C109 B.n70 VSUBS 0.007287f
C110 B.n71 VSUBS 0.007287f
C111 B.n72 VSUBS 0.007287f
C112 B.n73 VSUBS 0.007287f
C113 B.n74 VSUBS 0.007287f
C114 B.n75 VSUBS 0.007287f
C115 B.n76 VSUBS 0.007287f
C116 B.n77 VSUBS 0.007287f
C117 B.n78 VSUBS 0.007287f
C118 B.n79 VSUBS 0.007287f
C119 B.n80 VSUBS 0.007287f
C120 B.n81 VSUBS 0.018542f
C121 B.n82 VSUBS 0.007287f
C122 B.n83 VSUBS 0.007287f
C123 B.n84 VSUBS 0.007287f
C124 B.n85 VSUBS 0.007287f
C125 B.n86 VSUBS 0.007287f
C126 B.n87 VSUBS 0.007287f
C127 B.n88 VSUBS 0.007287f
C128 B.n89 VSUBS 0.007287f
C129 B.n90 VSUBS 0.007287f
C130 B.n91 VSUBS 0.007287f
C131 B.n92 VSUBS 0.007287f
C132 B.n93 VSUBS 0.017678f
C133 B.n94 VSUBS 0.007287f
C134 B.n95 VSUBS 0.007287f
C135 B.n96 VSUBS 0.007287f
C136 B.n97 VSUBS 0.007287f
C137 B.n98 VSUBS 0.007287f
C138 B.n99 VSUBS 0.007287f
C139 B.n100 VSUBS 0.007287f
C140 B.n101 VSUBS 0.007287f
C141 B.n102 VSUBS 0.007287f
C142 B.n103 VSUBS 0.007287f
C143 B.n104 VSUBS 0.007287f
C144 B.n105 VSUBS 0.007287f
C145 B.n106 VSUBS 0.007287f
C146 B.n107 VSUBS 0.007287f
C147 B.n108 VSUBS 0.007287f
C148 B.n109 VSUBS 0.007287f
C149 B.n110 VSUBS 0.007287f
C150 B.n111 VSUBS 0.007287f
C151 B.n112 VSUBS 0.007287f
C152 B.n113 VSUBS 0.007287f
C153 B.n114 VSUBS 0.007287f
C154 B.n115 VSUBS 0.007287f
C155 B.n116 VSUBS 0.007287f
C156 B.n117 VSUBS 0.007287f
C157 B.n118 VSUBS 0.007287f
C158 B.n119 VSUBS 0.007287f
C159 B.n120 VSUBS 0.007287f
C160 B.n121 VSUBS 0.007287f
C161 B.n122 VSUBS 0.007287f
C162 B.n123 VSUBS 0.007287f
C163 B.n124 VSUBS 0.007287f
C164 B.n125 VSUBS 0.007287f
C165 B.t11 VSUBS 0.702866f
C166 B.t10 VSUBS 0.70823f
C167 B.t9 VSUBS 0.22356f
C168 B.n126 VSUBS 0.127622f
C169 B.n127 VSUBS 0.065159f
C170 B.n128 VSUBS 0.016883f
C171 B.n129 VSUBS 0.007287f
C172 B.n130 VSUBS 0.007287f
C173 B.n131 VSUBS 0.007287f
C174 B.n132 VSUBS 0.007287f
C175 B.n133 VSUBS 0.007287f
C176 B.t5 VSUBS 0.702896f
C177 B.t4 VSUBS 0.708258f
C178 B.t3 VSUBS 0.22356f
C179 B.n134 VSUBS 0.127594f
C180 B.n135 VSUBS 0.065129f
C181 B.n136 VSUBS 0.007287f
C182 B.n137 VSUBS 0.007287f
C183 B.n138 VSUBS 0.007287f
C184 B.n139 VSUBS 0.007287f
C185 B.n140 VSUBS 0.007287f
C186 B.n141 VSUBS 0.007287f
C187 B.n142 VSUBS 0.007287f
C188 B.n143 VSUBS 0.007287f
C189 B.n144 VSUBS 0.007287f
C190 B.n145 VSUBS 0.007287f
C191 B.n146 VSUBS 0.007287f
C192 B.n147 VSUBS 0.007287f
C193 B.n148 VSUBS 0.007287f
C194 B.n149 VSUBS 0.007287f
C195 B.n150 VSUBS 0.007287f
C196 B.n151 VSUBS 0.007287f
C197 B.n152 VSUBS 0.007287f
C198 B.n153 VSUBS 0.007287f
C199 B.n154 VSUBS 0.007287f
C200 B.n155 VSUBS 0.007287f
C201 B.n156 VSUBS 0.007287f
C202 B.n157 VSUBS 0.007287f
C203 B.n158 VSUBS 0.007287f
C204 B.n159 VSUBS 0.007287f
C205 B.n160 VSUBS 0.007287f
C206 B.n161 VSUBS 0.007287f
C207 B.n162 VSUBS 0.007287f
C208 B.n163 VSUBS 0.007287f
C209 B.n164 VSUBS 0.007287f
C210 B.n165 VSUBS 0.007287f
C211 B.n166 VSUBS 0.007287f
C212 B.n167 VSUBS 0.018542f
C213 B.n168 VSUBS 0.007287f
C214 B.n169 VSUBS 0.007287f
C215 B.n170 VSUBS 0.007287f
C216 B.n171 VSUBS 0.007287f
C217 B.n172 VSUBS 0.007287f
C218 B.n173 VSUBS 0.007287f
C219 B.n174 VSUBS 0.007287f
C220 B.n175 VSUBS 0.007287f
C221 B.n176 VSUBS 0.007287f
C222 B.n177 VSUBS 0.007287f
C223 B.n178 VSUBS 0.007287f
C224 B.n179 VSUBS 0.007287f
C225 B.n180 VSUBS 0.007287f
C226 B.n181 VSUBS 0.007287f
C227 B.n182 VSUBS 0.007287f
C228 B.n183 VSUBS 0.007287f
C229 B.n184 VSUBS 0.007287f
C230 B.n185 VSUBS 0.007287f
C231 B.n186 VSUBS 0.017678f
C232 B.n187 VSUBS 0.017678f
C233 B.n188 VSUBS 0.018542f
C234 B.n189 VSUBS 0.007287f
C235 B.n190 VSUBS 0.007287f
C236 B.n191 VSUBS 0.007287f
C237 B.n192 VSUBS 0.007287f
C238 B.n193 VSUBS 0.007287f
C239 B.n194 VSUBS 0.007287f
C240 B.n195 VSUBS 0.007287f
C241 B.n196 VSUBS 0.007287f
C242 B.n197 VSUBS 0.007287f
C243 B.n198 VSUBS 0.007287f
C244 B.n199 VSUBS 0.007287f
C245 B.n200 VSUBS 0.007287f
C246 B.n201 VSUBS 0.007287f
C247 B.n202 VSUBS 0.007287f
C248 B.n203 VSUBS 0.007287f
C249 B.n204 VSUBS 0.007287f
C250 B.n205 VSUBS 0.007287f
C251 B.n206 VSUBS 0.007287f
C252 B.n207 VSUBS 0.007287f
C253 B.n208 VSUBS 0.007287f
C254 B.n209 VSUBS 0.007287f
C255 B.n210 VSUBS 0.007287f
C256 B.n211 VSUBS 0.007287f
C257 B.n212 VSUBS 0.007287f
C258 B.n213 VSUBS 0.007287f
C259 B.n214 VSUBS 0.007287f
C260 B.n215 VSUBS 0.007287f
C261 B.n216 VSUBS 0.007287f
C262 B.n217 VSUBS 0.007287f
C263 B.n218 VSUBS 0.007287f
C264 B.n219 VSUBS 0.007287f
C265 B.n220 VSUBS 0.007287f
C266 B.n221 VSUBS 0.007287f
C267 B.n222 VSUBS 0.007287f
C268 B.n223 VSUBS 0.007287f
C269 B.n224 VSUBS 0.007287f
C270 B.n225 VSUBS 0.007287f
C271 B.n226 VSUBS 0.007287f
C272 B.n227 VSUBS 0.007287f
C273 B.n228 VSUBS 0.007287f
C274 B.n229 VSUBS 0.007287f
C275 B.n230 VSUBS 0.007287f
C276 B.n231 VSUBS 0.007287f
C277 B.n232 VSUBS 0.007287f
C278 B.n233 VSUBS 0.007287f
C279 B.n234 VSUBS 0.007287f
C280 B.n235 VSUBS 0.007287f
C281 B.n236 VSUBS 0.007287f
C282 B.n237 VSUBS 0.007287f
C283 B.n238 VSUBS 0.007287f
C284 B.n239 VSUBS 0.007287f
C285 B.n240 VSUBS 0.007287f
C286 B.n241 VSUBS 0.007287f
C287 B.n242 VSUBS 0.007287f
C288 B.n243 VSUBS 0.007287f
C289 B.n244 VSUBS 0.007287f
C290 B.n245 VSUBS 0.007287f
C291 B.n246 VSUBS 0.007287f
C292 B.n247 VSUBS 0.007287f
C293 B.n248 VSUBS 0.007287f
C294 B.n249 VSUBS 0.007287f
C295 B.n250 VSUBS 0.007287f
C296 B.n251 VSUBS 0.007287f
C297 B.n252 VSUBS 0.007287f
C298 B.n253 VSUBS 0.007287f
C299 B.n254 VSUBS 0.007287f
C300 B.n255 VSUBS 0.007287f
C301 B.n256 VSUBS 0.007287f
C302 B.n257 VSUBS 0.007287f
C303 B.n258 VSUBS 0.007287f
C304 B.n259 VSUBS 0.007287f
C305 B.n260 VSUBS 0.007287f
C306 B.n261 VSUBS 0.007287f
C307 B.n262 VSUBS 0.007287f
C308 B.n263 VSUBS 0.007287f
C309 B.n264 VSUBS 0.007287f
C310 B.n265 VSUBS 0.007287f
C311 B.n266 VSUBS 0.007287f
C312 B.n267 VSUBS 0.007287f
C313 B.n268 VSUBS 0.007287f
C314 B.n269 VSUBS 0.007287f
C315 B.n270 VSUBS 0.007287f
C316 B.n271 VSUBS 0.007287f
C317 B.n272 VSUBS 0.007287f
C318 B.n273 VSUBS 0.007287f
C319 B.n274 VSUBS 0.007287f
C320 B.n275 VSUBS 0.007287f
C321 B.n276 VSUBS 0.007287f
C322 B.n277 VSUBS 0.007287f
C323 B.n278 VSUBS 0.007287f
C324 B.n279 VSUBS 0.007287f
C325 B.n280 VSUBS 0.007287f
C326 B.n281 VSUBS 0.007287f
C327 B.n282 VSUBS 0.007287f
C328 B.n283 VSUBS 0.007287f
C329 B.n284 VSUBS 0.004822f
C330 B.n285 VSUBS 0.016883f
C331 B.n286 VSUBS 0.006108f
C332 B.n287 VSUBS 0.007287f
C333 B.n288 VSUBS 0.007287f
C334 B.n289 VSUBS 0.007287f
C335 B.n290 VSUBS 0.007287f
C336 B.n291 VSUBS 0.007287f
C337 B.n292 VSUBS 0.007287f
C338 B.n293 VSUBS 0.007287f
C339 B.n294 VSUBS 0.007287f
C340 B.n295 VSUBS 0.007287f
C341 B.n296 VSUBS 0.007287f
C342 B.n297 VSUBS 0.007287f
C343 B.n298 VSUBS 0.006108f
C344 B.n299 VSUBS 0.007287f
C345 B.n300 VSUBS 0.007287f
C346 B.n301 VSUBS 0.004822f
C347 B.n302 VSUBS 0.007287f
C348 B.n303 VSUBS 0.007287f
C349 B.n304 VSUBS 0.007287f
C350 B.n305 VSUBS 0.007287f
C351 B.n306 VSUBS 0.007287f
C352 B.n307 VSUBS 0.007287f
C353 B.n308 VSUBS 0.007287f
C354 B.n309 VSUBS 0.007287f
C355 B.n310 VSUBS 0.007287f
C356 B.n311 VSUBS 0.007287f
C357 B.n312 VSUBS 0.007287f
C358 B.n313 VSUBS 0.007287f
C359 B.n314 VSUBS 0.007287f
C360 B.n315 VSUBS 0.007287f
C361 B.n316 VSUBS 0.007287f
C362 B.n317 VSUBS 0.007287f
C363 B.n318 VSUBS 0.007287f
C364 B.n319 VSUBS 0.007287f
C365 B.n320 VSUBS 0.007287f
C366 B.n321 VSUBS 0.007287f
C367 B.n322 VSUBS 0.007287f
C368 B.n323 VSUBS 0.007287f
C369 B.n324 VSUBS 0.007287f
C370 B.n325 VSUBS 0.007287f
C371 B.n326 VSUBS 0.007287f
C372 B.n327 VSUBS 0.007287f
C373 B.n328 VSUBS 0.007287f
C374 B.n329 VSUBS 0.007287f
C375 B.n330 VSUBS 0.007287f
C376 B.n331 VSUBS 0.007287f
C377 B.n332 VSUBS 0.007287f
C378 B.n333 VSUBS 0.007287f
C379 B.n334 VSUBS 0.007287f
C380 B.n335 VSUBS 0.007287f
C381 B.n336 VSUBS 0.007287f
C382 B.n337 VSUBS 0.007287f
C383 B.n338 VSUBS 0.007287f
C384 B.n339 VSUBS 0.007287f
C385 B.n340 VSUBS 0.007287f
C386 B.n341 VSUBS 0.007287f
C387 B.n342 VSUBS 0.007287f
C388 B.n343 VSUBS 0.007287f
C389 B.n344 VSUBS 0.007287f
C390 B.n345 VSUBS 0.007287f
C391 B.n346 VSUBS 0.007287f
C392 B.n347 VSUBS 0.007287f
C393 B.n348 VSUBS 0.007287f
C394 B.n349 VSUBS 0.007287f
C395 B.n350 VSUBS 0.007287f
C396 B.n351 VSUBS 0.007287f
C397 B.n352 VSUBS 0.007287f
C398 B.n353 VSUBS 0.007287f
C399 B.n354 VSUBS 0.007287f
C400 B.n355 VSUBS 0.007287f
C401 B.n356 VSUBS 0.007287f
C402 B.n357 VSUBS 0.007287f
C403 B.n358 VSUBS 0.007287f
C404 B.n359 VSUBS 0.007287f
C405 B.n360 VSUBS 0.007287f
C406 B.n361 VSUBS 0.007287f
C407 B.n362 VSUBS 0.007287f
C408 B.n363 VSUBS 0.007287f
C409 B.n364 VSUBS 0.007287f
C410 B.n365 VSUBS 0.007287f
C411 B.n366 VSUBS 0.007287f
C412 B.n367 VSUBS 0.007287f
C413 B.n368 VSUBS 0.007287f
C414 B.n369 VSUBS 0.007287f
C415 B.n370 VSUBS 0.007287f
C416 B.n371 VSUBS 0.007287f
C417 B.n372 VSUBS 0.007287f
C418 B.n373 VSUBS 0.007287f
C419 B.n374 VSUBS 0.007287f
C420 B.n375 VSUBS 0.007287f
C421 B.n376 VSUBS 0.007287f
C422 B.n377 VSUBS 0.007287f
C423 B.n378 VSUBS 0.007287f
C424 B.n379 VSUBS 0.007287f
C425 B.n380 VSUBS 0.007287f
C426 B.n381 VSUBS 0.007287f
C427 B.n382 VSUBS 0.007287f
C428 B.n383 VSUBS 0.007287f
C429 B.n384 VSUBS 0.007287f
C430 B.n385 VSUBS 0.007287f
C431 B.n386 VSUBS 0.007287f
C432 B.n387 VSUBS 0.007287f
C433 B.n388 VSUBS 0.007287f
C434 B.n389 VSUBS 0.007287f
C435 B.n390 VSUBS 0.007287f
C436 B.n391 VSUBS 0.007287f
C437 B.n392 VSUBS 0.007287f
C438 B.n393 VSUBS 0.007287f
C439 B.n394 VSUBS 0.007287f
C440 B.n395 VSUBS 0.007287f
C441 B.n396 VSUBS 0.018542f
C442 B.n397 VSUBS 0.017755f
C443 B.n398 VSUBS 0.018465f
C444 B.n399 VSUBS 0.007287f
C445 B.n400 VSUBS 0.007287f
C446 B.n401 VSUBS 0.007287f
C447 B.n402 VSUBS 0.007287f
C448 B.n403 VSUBS 0.007287f
C449 B.n404 VSUBS 0.007287f
C450 B.n405 VSUBS 0.007287f
C451 B.n406 VSUBS 0.007287f
C452 B.n407 VSUBS 0.007287f
C453 B.n408 VSUBS 0.007287f
C454 B.n409 VSUBS 0.007287f
C455 B.n410 VSUBS 0.007287f
C456 B.n411 VSUBS 0.007287f
C457 B.n412 VSUBS 0.007287f
C458 B.n413 VSUBS 0.007287f
C459 B.n414 VSUBS 0.007287f
C460 B.n415 VSUBS 0.007287f
C461 B.n416 VSUBS 0.007287f
C462 B.n417 VSUBS 0.007287f
C463 B.n418 VSUBS 0.007287f
C464 B.n419 VSUBS 0.007287f
C465 B.n420 VSUBS 0.007287f
C466 B.n421 VSUBS 0.007287f
C467 B.n422 VSUBS 0.007287f
C468 B.n423 VSUBS 0.007287f
C469 B.n424 VSUBS 0.007287f
C470 B.n425 VSUBS 0.007287f
C471 B.n426 VSUBS 0.007287f
C472 B.n427 VSUBS 0.007287f
C473 B.n428 VSUBS 0.007287f
C474 B.n429 VSUBS 0.007287f
C475 B.n430 VSUBS 0.007287f
C476 B.n431 VSUBS 0.007287f
C477 B.n432 VSUBS 0.017678f
C478 B.n433 VSUBS 0.017678f
C479 B.n434 VSUBS 0.018542f
C480 B.n435 VSUBS 0.007287f
C481 B.n436 VSUBS 0.007287f
C482 B.n437 VSUBS 0.007287f
C483 B.n438 VSUBS 0.007287f
C484 B.n439 VSUBS 0.007287f
C485 B.n440 VSUBS 0.007287f
C486 B.n441 VSUBS 0.007287f
C487 B.n442 VSUBS 0.007287f
C488 B.n443 VSUBS 0.007287f
C489 B.n444 VSUBS 0.007287f
C490 B.n445 VSUBS 0.007287f
C491 B.n446 VSUBS 0.007287f
C492 B.n447 VSUBS 0.007287f
C493 B.n448 VSUBS 0.007287f
C494 B.n449 VSUBS 0.007287f
C495 B.n450 VSUBS 0.007287f
C496 B.n451 VSUBS 0.007287f
C497 B.n452 VSUBS 0.007287f
C498 B.n453 VSUBS 0.007287f
C499 B.n454 VSUBS 0.007287f
C500 B.n455 VSUBS 0.007287f
C501 B.n456 VSUBS 0.007287f
C502 B.n457 VSUBS 0.007287f
C503 B.n458 VSUBS 0.007287f
C504 B.n459 VSUBS 0.007287f
C505 B.n460 VSUBS 0.007287f
C506 B.n461 VSUBS 0.007287f
C507 B.n462 VSUBS 0.007287f
C508 B.n463 VSUBS 0.007287f
C509 B.n464 VSUBS 0.007287f
C510 B.n465 VSUBS 0.007287f
C511 B.n466 VSUBS 0.007287f
C512 B.n467 VSUBS 0.007287f
C513 B.n468 VSUBS 0.007287f
C514 B.n469 VSUBS 0.007287f
C515 B.n470 VSUBS 0.007287f
C516 B.n471 VSUBS 0.007287f
C517 B.n472 VSUBS 0.007287f
C518 B.n473 VSUBS 0.007287f
C519 B.n474 VSUBS 0.007287f
C520 B.n475 VSUBS 0.007287f
C521 B.n476 VSUBS 0.007287f
C522 B.n477 VSUBS 0.007287f
C523 B.n478 VSUBS 0.007287f
C524 B.n479 VSUBS 0.007287f
C525 B.n480 VSUBS 0.007287f
C526 B.n481 VSUBS 0.007287f
C527 B.n482 VSUBS 0.007287f
C528 B.n483 VSUBS 0.007287f
C529 B.n484 VSUBS 0.007287f
C530 B.n485 VSUBS 0.007287f
C531 B.n486 VSUBS 0.007287f
C532 B.n487 VSUBS 0.007287f
C533 B.n488 VSUBS 0.007287f
C534 B.n489 VSUBS 0.007287f
C535 B.n490 VSUBS 0.007287f
C536 B.n491 VSUBS 0.007287f
C537 B.n492 VSUBS 0.007287f
C538 B.n493 VSUBS 0.007287f
C539 B.n494 VSUBS 0.007287f
C540 B.n495 VSUBS 0.007287f
C541 B.n496 VSUBS 0.007287f
C542 B.n497 VSUBS 0.007287f
C543 B.n498 VSUBS 0.007287f
C544 B.n499 VSUBS 0.007287f
C545 B.n500 VSUBS 0.007287f
C546 B.n501 VSUBS 0.007287f
C547 B.n502 VSUBS 0.007287f
C548 B.n503 VSUBS 0.007287f
C549 B.n504 VSUBS 0.007287f
C550 B.n505 VSUBS 0.007287f
C551 B.n506 VSUBS 0.007287f
C552 B.n507 VSUBS 0.007287f
C553 B.n508 VSUBS 0.007287f
C554 B.n509 VSUBS 0.007287f
C555 B.n510 VSUBS 0.007287f
C556 B.n511 VSUBS 0.007287f
C557 B.n512 VSUBS 0.007287f
C558 B.n513 VSUBS 0.007287f
C559 B.n514 VSUBS 0.007287f
C560 B.n515 VSUBS 0.007287f
C561 B.n516 VSUBS 0.007287f
C562 B.n517 VSUBS 0.007287f
C563 B.n518 VSUBS 0.007287f
C564 B.n519 VSUBS 0.007287f
C565 B.n520 VSUBS 0.007287f
C566 B.n521 VSUBS 0.007287f
C567 B.n522 VSUBS 0.007287f
C568 B.n523 VSUBS 0.007287f
C569 B.n524 VSUBS 0.007287f
C570 B.n525 VSUBS 0.007287f
C571 B.n526 VSUBS 0.007287f
C572 B.n527 VSUBS 0.007287f
C573 B.n528 VSUBS 0.007287f
C574 B.n529 VSUBS 0.007287f
C575 B.n530 VSUBS 0.004822f
C576 B.n531 VSUBS 0.016883f
C577 B.n532 VSUBS 0.006108f
C578 B.n533 VSUBS 0.007287f
C579 B.n534 VSUBS 0.007287f
C580 B.n535 VSUBS 0.007287f
C581 B.n536 VSUBS 0.007287f
C582 B.n537 VSUBS 0.007287f
C583 B.n538 VSUBS 0.007287f
C584 B.n539 VSUBS 0.007287f
C585 B.n540 VSUBS 0.007287f
C586 B.n541 VSUBS 0.007287f
C587 B.n542 VSUBS 0.007287f
C588 B.n543 VSUBS 0.007287f
C589 B.n544 VSUBS 0.006108f
C590 B.n545 VSUBS 0.007287f
C591 B.n546 VSUBS 0.007287f
C592 B.n547 VSUBS 0.004822f
C593 B.n548 VSUBS 0.007287f
C594 B.n549 VSUBS 0.007287f
C595 B.n550 VSUBS 0.007287f
C596 B.n551 VSUBS 0.007287f
C597 B.n552 VSUBS 0.007287f
C598 B.n553 VSUBS 0.007287f
C599 B.n554 VSUBS 0.007287f
C600 B.n555 VSUBS 0.007287f
C601 B.n556 VSUBS 0.007287f
C602 B.n557 VSUBS 0.007287f
C603 B.n558 VSUBS 0.007287f
C604 B.n559 VSUBS 0.007287f
C605 B.n560 VSUBS 0.007287f
C606 B.n561 VSUBS 0.007287f
C607 B.n562 VSUBS 0.007287f
C608 B.n563 VSUBS 0.007287f
C609 B.n564 VSUBS 0.007287f
C610 B.n565 VSUBS 0.007287f
C611 B.n566 VSUBS 0.007287f
C612 B.n567 VSUBS 0.007287f
C613 B.n568 VSUBS 0.007287f
C614 B.n569 VSUBS 0.007287f
C615 B.n570 VSUBS 0.007287f
C616 B.n571 VSUBS 0.007287f
C617 B.n572 VSUBS 0.007287f
C618 B.n573 VSUBS 0.007287f
C619 B.n574 VSUBS 0.007287f
C620 B.n575 VSUBS 0.007287f
C621 B.n576 VSUBS 0.007287f
C622 B.n577 VSUBS 0.007287f
C623 B.n578 VSUBS 0.007287f
C624 B.n579 VSUBS 0.007287f
C625 B.n580 VSUBS 0.007287f
C626 B.n581 VSUBS 0.007287f
C627 B.n582 VSUBS 0.007287f
C628 B.n583 VSUBS 0.007287f
C629 B.n584 VSUBS 0.007287f
C630 B.n585 VSUBS 0.007287f
C631 B.n586 VSUBS 0.007287f
C632 B.n587 VSUBS 0.007287f
C633 B.n588 VSUBS 0.007287f
C634 B.n589 VSUBS 0.007287f
C635 B.n590 VSUBS 0.007287f
C636 B.n591 VSUBS 0.007287f
C637 B.n592 VSUBS 0.007287f
C638 B.n593 VSUBS 0.007287f
C639 B.n594 VSUBS 0.007287f
C640 B.n595 VSUBS 0.007287f
C641 B.n596 VSUBS 0.007287f
C642 B.n597 VSUBS 0.007287f
C643 B.n598 VSUBS 0.007287f
C644 B.n599 VSUBS 0.007287f
C645 B.n600 VSUBS 0.007287f
C646 B.n601 VSUBS 0.007287f
C647 B.n602 VSUBS 0.007287f
C648 B.n603 VSUBS 0.007287f
C649 B.n604 VSUBS 0.007287f
C650 B.n605 VSUBS 0.007287f
C651 B.n606 VSUBS 0.007287f
C652 B.n607 VSUBS 0.007287f
C653 B.n608 VSUBS 0.007287f
C654 B.n609 VSUBS 0.007287f
C655 B.n610 VSUBS 0.007287f
C656 B.n611 VSUBS 0.007287f
C657 B.n612 VSUBS 0.007287f
C658 B.n613 VSUBS 0.007287f
C659 B.n614 VSUBS 0.007287f
C660 B.n615 VSUBS 0.007287f
C661 B.n616 VSUBS 0.007287f
C662 B.n617 VSUBS 0.007287f
C663 B.n618 VSUBS 0.007287f
C664 B.n619 VSUBS 0.007287f
C665 B.n620 VSUBS 0.007287f
C666 B.n621 VSUBS 0.007287f
C667 B.n622 VSUBS 0.007287f
C668 B.n623 VSUBS 0.007287f
C669 B.n624 VSUBS 0.007287f
C670 B.n625 VSUBS 0.007287f
C671 B.n626 VSUBS 0.007287f
C672 B.n627 VSUBS 0.007287f
C673 B.n628 VSUBS 0.007287f
C674 B.n629 VSUBS 0.007287f
C675 B.n630 VSUBS 0.007287f
C676 B.n631 VSUBS 0.007287f
C677 B.n632 VSUBS 0.007287f
C678 B.n633 VSUBS 0.007287f
C679 B.n634 VSUBS 0.007287f
C680 B.n635 VSUBS 0.007287f
C681 B.n636 VSUBS 0.007287f
C682 B.n637 VSUBS 0.007287f
C683 B.n638 VSUBS 0.007287f
C684 B.n639 VSUBS 0.007287f
C685 B.n640 VSUBS 0.007287f
C686 B.n641 VSUBS 0.007287f
C687 B.n642 VSUBS 0.018542f
C688 B.n643 VSUBS 0.018542f
C689 B.n644 VSUBS 0.017678f
C690 B.n645 VSUBS 0.007287f
C691 B.n646 VSUBS 0.007287f
C692 B.n647 VSUBS 0.007287f
C693 B.n648 VSUBS 0.007287f
C694 B.n649 VSUBS 0.007287f
C695 B.n650 VSUBS 0.007287f
C696 B.n651 VSUBS 0.007287f
C697 B.n652 VSUBS 0.007287f
C698 B.n653 VSUBS 0.007287f
C699 B.n654 VSUBS 0.007287f
C700 B.n655 VSUBS 0.007287f
C701 B.n656 VSUBS 0.007287f
C702 B.n657 VSUBS 0.007287f
C703 B.n658 VSUBS 0.007287f
C704 B.n659 VSUBS 0.009509f
C705 B.n660 VSUBS 0.01013f
C706 B.n661 VSUBS 0.020143f
C707 VDD2.t1 VSUBS 5.64561f
C708 VDD2.t0 VSUBS 4.72907f
C709 VDD2.n0 VSUBS 4.88449f
C710 VTAIL.t1 VSUBS 4.67735f
C711 VTAIL.n0 VSUBS 2.88992f
C712 VTAIL.t2 VSUBS 4.67735f
C713 VTAIL.n1 VSUBS 2.89659f
C714 VTAIL.t0 VSUBS 4.67735f
C715 VTAIL.n2 VSUBS 2.84871f
C716 VTAIL.t3 VSUBS 4.67735f
C717 VTAIL.n3 VSUBS 2.78865f
C718 VN.t0 VSUBS 0.954339f
C719 VN.t1 VSUBS 1.02029f
.ends

