* NGSPICE file created from diff_pair_sample_1104.ext - technology: sky130A

.subckt diff_pair_sample_1104 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t1 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=2.4453 ps=15.15 w=14.82 l=3.05
X1 VTAIL.t5 VN.t0 VDD2.t5 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=2.4453 ps=15.15 w=14.82 l=3.05
X2 VDD1.t5 VP.t1 VTAIL.t10 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=2.4453 ps=15.15 w=14.82 l=3.05
X3 VDD2.t4 VN.t1 VTAIL.t4 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=2.4453 ps=15.15 w=14.82 l=3.05
X4 B.t11 B.t9 B.t10 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=0 ps=0 w=14.82 l=3.05
X5 VDD1.t3 VP.t2 VTAIL.t9 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=5.7798 ps=30.42 w=14.82 l=3.05
X6 B.t8 B.t6 B.t7 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=0 ps=0 w=14.82 l=3.05
X7 VDD2.t3 VN.t2 VTAIL.t2 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=5.7798 ps=30.42 w=14.82 l=3.05
X8 VDD2.t2 VN.t3 VTAIL.t3 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=5.7798 ps=30.42 w=14.82 l=3.05
X9 VTAIL.t0 VN.t4 VDD2.t1 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=2.4453 ps=15.15 w=14.82 l=3.05
X10 VDD1.t2 VP.t3 VTAIL.t8 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=2.4453 ps=15.15 w=14.82 l=3.05
X11 B.t5 B.t3 B.t4 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=0 ps=0 w=14.82 l=3.05
X12 VDD2.t0 VN.t5 VTAIL.t1 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=2.4453 ps=15.15 w=14.82 l=3.05
X13 B.t2 B.t0 B.t1 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=5.7798 pd=30.42 as=0 ps=0 w=14.82 l=3.05
X14 VDD1.t4 VP.t4 VTAIL.t7 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=5.7798 ps=30.42 w=14.82 l=3.05
X15 VTAIL.t6 VP.t5 VDD1.t0 w_n3674_n3932# sky130_fd_pr__pfet_01v8 ad=2.4453 pd=15.15 as=2.4453 ps=15.15 w=14.82 l=3.05
R0 VP.n13 VP.n10 161.3
R1 VP.n15 VP.n14 161.3
R2 VP.n16 VP.n9 161.3
R3 VP.n18 VP.n17 161.3
R4 VP.n19 VP.n8 161.3
R5 VP.n21 VP.n20 161.3
R6 VP.n44 VP.n43 161.3
R7 VP.n42 VP.n1 161.3
R8 VP.n41 VP.n40 161.3
R9 VP.n39 VP.n2 161.3
R10 VP.n38 VP.n37 161.3
R11 VP.n36 VP.n3 161.3
R12 VP.n35 VP.n34 161.3
R13 VP.n33 VP.n4 161.3
R14 VP.n32 VP.n31 161.3
R15 VP.n30 VP.n5 161.3
R16 VP.n29 VP.n28 161.3
R17 VP.n27 VP.n6 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n11 VP.t1 150.538
R20 VP.n35 VP.t0 117.103
R21 VP.n24 VP.t3 117.103
R22 VP.n0 VP.t4 117.103
R23 VP.n12 VP.t5 117.103
R24 VP.n7 VP.t2 117.103
R25 VP.n24 VP.n23 71.5558
R26 VP.n45 VP.n0 71.5558
R27 VP.n22 VP.n7 71.5558
R28 VP.n30 VP.n29 56.5617
R29 VP.n41 VP.n2 56.5617
R30 VP.n18 VP.n9 56.5617
R31 VP.n23 VP.n22 52.6889
R32 VP.n12 VP.n11 49.4409
R33 VP.n25 VP.n6 24.5923
R34 VP.n29 VP.n6 24.5923
R35 VP.n31 VP.n30 24.5923
R36 VP.n31 VP.n4 24.5923
R37 VP.n35 VP.n4 24.5923
R38 VP.n36 VP.n35 24.5923
R39 VP.n37 VP.n36 24.5923
R40 VP.n37 VP.n2 24.5923
R41 VP.n42 VP.n41 24.5923
R42 VP.n43 VP.n42 24.5923
R43 VP.n19 VP.n18 24.5923
R44 VP.n20 VP.n19 24.5923
R45 VP.n13 VP.n12 24.5923
R46 VP.n14 VP.n13 24.5923
R47 VP.n14 VP.n9 24.5923
R48 VP.n25 VP.n24 18.6903
R49 VP.n43 VP.n0 18.6903
R50 VP.n20 VP.n7 18.6903
R51 VP.n11 VP.n10 3.9675
R52 VP.n22 VP.n21 0.354861
R53 VP.n26 VP.n23 0.354861
R54 VP.n45 VP.n44 0.354861
R55 VP VP.n45 0.267071
R56 VP.n15 VP.n10 0.189894
R57 VP.n16 VP.n15 0.189894
R58 VP.n17 VP.n16 0.189894
R59 VP.n17 VP.n8 0.189894
R60 VP.n21 VP.n8 0.189894
R61 VP.n27 VP.n26 0.189894
R62 VP.n28 VP.n27 0.189894
R63 VP.n28 VP.n5 0.189894
R64 VP.n32 VP.n5 0.189894
R65 VP.n33 VP.n32 0.189894
R66 VP.n34 VP.n33 0.189894
R67 VP.n34 VP.n3 0.189894
R68 VP.n38 VP.n3 0.189894
R69 VP.n39 VP.n38 0.189894
R70 VP.n40 VP.n39 0.189894
R71 VP.n40 VP.n1 0.189894
R72 VP.n44 VP.n1 0.189894
R73 VDD1.n76 VDD1.n0 756.745
R74 VDD1.n157 VDD1.n81 756.745
R75 VDD1.n77 VDD1.n76 585
R76 VDD1.n75 VDD1.n74 585
R77 VDD1.n73 VDD1.n3 585
R78 VDD1.n7 VDD1.n4 585
R79 VDD1.n68 VDD1.n67 585
R80 VDD1.n66 VDD1.n65 585
R81 VDD1.n9 VDD1.n8 585
R82 VDD1.n60 VDD1.n59 585
R83 VDD1.n58 VDD1.n57 585
R84 VDD1.n13 VDD1.n12 585
R85 VDD1.n52 VDD1.n51 585
R86 VDD1.n50 VDD1.n49 585
R87 VDD1.n17 VDD1.n16 585
R88 VDD1.n44 VDD1.n43 585
R89 VDD1.n42 VDD1.n41 585
R90 VDD1.n21 VDD1.n20 585
R91 VDD1.n36 VDD1.n35 585
R92 VDD1.n34 VDD1.n33 585
R93 VDD1.n25 VDD1.n24 585
R94 VDD1.n28 VDD1.n27 585
R95 VDD1.n108 VDD1.n107 585
R96 VDD1.n105 VDD1.n104 585
R97 VDD1.n114 VDD1.n113 585
R98 VDD1.n116 VDD1.n115 585
R99 VDD1.n101 VDD1.n100 585
R100 VDD1.n122 VDD1.n121 585
R101 VDD1.n124 VDD1.n123 585
R102 VDD1.n97 VDD1.n96 585
R103 VDD1.n130 VDD1.n129 585
R104 VDD1.n132 VDD1.n131 585
R105 VDD1.n93 VDD1.n92 585
R106 VDD1.n138 VDD1.n137 585
R107 VDD1.n140 VDD1.n139 585
R108 VDD1.n89 VDD1.n88 585
R109 VDD1.n146 VDD1.n145 585
R110 VDD1.n149 VDD1.n148 585
R111 VDD1.n147 VDD1.n85 585
R112 VDD1.n154 VDD1.n84 585
R113 VDD1.n156 VDD1.n155 585
R114 VDD1.n158 VDD1.n157 585
R115 VDD1.t5 VDD1.n26 327.466
R116 VDD1.t2 VDD1.n106 327.466
R117 VDD1.n76 VDD1.n75 171.744
R118 VDD1.n75 VDD1.n3 171.744
R119 VDD1.n7 VDD1.n3 171.744
R120 VDD1.n67 VDD1.n7 171.744
R121 VDD1.n67 VDD1.n66 171.744
R122 VDD1.n66 VDD1.n8 171.744
R123 VDD1.n59 VDD1.n8 171.744
R124 VDD1.n59 VDD1.n58 171.744
R125 VDD1.n58 VDD1.n12 171.744
R126 VDD1.n51 VDD1.n12 171.744
R127 VDD1.n51 VDD1.n50 171.744
R128 VDD1.n50 VDD1.n16 171.744
R129 VDD1.n43 VDD1.n16 171.744
R130 VDD1.n43 VDD1.n42 171.744
R131 VDD1.n42 VDD1.n20 171.744
R132 VDD1.n35 VDD1.n20 171.744
R133 VDD1.n35 VDD1.n34 171.744
R134 VDD1.n34 VDD1.n24 171.744
R135 VDD1.n27 VDD1.n24 171.744
R136 VDD1.n107 VDD1.n104 171.744
R137 VDD1.n114 VDD1.n104 171.744
R138 VDD1.n115 VDD1.n114 171.744
R139 VDD1.n115 VDD1.n100 171.744
R140 VDD1.n122 VDD1.n100 171.744
R141 VDD1.n123 VDD1.n122 171.744
R142 VDD1.n123 VDD1.n96 171.744
R143 VDD1.n130 VDD1.n96 171.744
R144 VDD1.n131 VDD1.n130 171.744
R145 VDD1.n131 VDD1.n92 171.744
R146 VDD1.n138 VDD1.n92 171.744
R147 VDD1.n139 VDD1.n138 171.744
R148 VDD1.n139 VDD1.n88 171.744
R149 VDD1.n146 VDD1.n88 171.744
R150 VDD1.n148 VDD1.n146 171.744
R151 VDD1.n148 VDD1.n147 171.744
R152 VDD1.n147 VDD1.n84 171.744
R153 VDD1.n156 VDD1.n84 171.744
R154 VDD1.n157 VDD1.n156 171.744
R155 VDD1.n27 VDD1.t5 85.8723
R156 VDD1.n107 VDD1.t2 85.8723
R157 VDD1.n163 VDD1.n162 74.9304
R158 VDD1.n165 VDD1.n164 74.2573
R159 VDD1 VDD1.n80 54.5986
R160 VDD1.n163 VDD1.n161 54.485
R161 VDD1.n165 VDD1.n163 48.0009
R162 VDD1.n28 VDD1.n26 16.3895
R163 VDD1.n108 VDD1.n106 16.3895
R164 VDD1.n74 VDD1.n73 13.1884
R165 VDD1.n155 VDD1.n154 13.1884
R166 VDD1.n77 VDD1.n2 12.8005
R167 VDD1.n72 VDD1.n4 12.8005
R168 VDD1.n29 VDD1.n25 12.8005
R169 VDD1.n109 VDD1.n105 12.8005
R170 VDD1.n153 VDD1.n85 12.8005
R171 VDD1.n158 VDD1.n83 12.8005
R172 VDD1.n78 VDD1.n0 12.0247
R173 VDD1.n69 VDD1.n68 12.0247
R174 VDD1.n33 VDD1.n32 12.0247
R175 VDD1.n113 VDD1.n112 12.0247
R176 VDD1.n150 VDD1.n149 12.0247
R177 VDD1.n159 VDD1.n81 12.0247
R178 VDD1.n65 VDD1.n6 11.249
R179 VDD1.n36 VDD1.n23 11.249
R180 VDD1.n116 VDD1.n103 11.249
R181 VDD1.n145 VDD1.n87 11.249
R182 VDD1.n64 VDD1.n9 10.4732
R183 VDD1.n37 VDD1.n21 10.4732
R184 VDD1.n117 VDD1.n101 10.4732
R185 VDD1.n144 VDD1.n89 10.4732
R186 VDD1.n61 VDD1.n60 9.69747
R187 VDD1.n41 VDD1.n40 9.69747
R188 VDD1.n121 VDD1.n120 9.69747
R189 VDD1.n141 VDD1.n140 9.69747
R190 VDD1.n80 VDD1.n79 9.45567
R191 VDD1.n161 VDD1.n160 9.45567
R192 VDD1.n54 VDD1.n53 9.3005
R193 VDD1.n56 VDD1.n55 9.3005
R194 VDD1.n11 VDD1.n10 9.3005
R195 VDD1.n62 VDD1.n61 9.3005
R196 VDD1.n64 VDD1.n63 9.3005
R197 VDD1.n6 VDD1.n5 9.3005
R198 VDD1.n70 VDD1.n69 9.3005
R199 VDD1.n72 VDD1.n71 9.3005
R200 VDD1.n79 VDD1.n78 9.3005
R201 VDD1.n2 VDD1.n1 9.3005
R202 VDD1.n15 VDD1.n14 9.3005
R203 VDD1.n48 VDD1.n47 9.3005
R204 VDD1.n46 VDD1.n45 9.3005
R205 VDD1.n19 VDD1.n18 9.3005
R206 VDD1.n40 VDD1.n39 9.3005
R207 VDD1.n38 VDD1.n37 9.3005
R208 VDD1.n23 VDD1.n22 9.3005
R209 VDD1.n32 VDD1.n31 9.3005
R210 VDD1.n30 VDD1.n29 9.3005
R211 VDD1.n160 VDD1.n159 9.3005
R212 VDD1.n83 VDD1.n82 9.3005
R213 VDD1.n128 VDD1.n127 9.3005
R214 VDD1.n126 VDD1.n125 9.3005
R215 VDD1.n99 VDD1.n98 9.3005
R216 VDD1.n120 VDD1.n119 9.3005
R217 VDD1.n118 VDD1.n117 9.3005
R218 VDD1.n103 VDD1.n102 9.3005
R219 VDD1.n112 VDD1.n111 9.3005
R220 VDD1.n110 VDD1.n109 9.3005
R221 VDD1.n95 VDD1.n94 9.3005
R222 VDD1.n134 VDD1.n133 9.3005
R223 VDD1.n136 VDD1.n135 9.3005
R224 VDD1.n91 VDD1.n90 9.3005
R225 VDD1.n142 VDD1.n141 9.3005
R226 VDD1.n144 VDD1.n143 9.3005
R227 VDD1.n87 VDD1.n86 9.3005
R228 VDD1.n151 VDD1.n150 9.3005
R229 VDD1.n153 VDD1.n152 9.3005
R230 VDD1.n57 VDD1.n11 8.92171
R231 VDD1.n44 VDD1.n19 8.92171
R232 VDD1.n124 VDD1.n99 8.92171
R233 VDD1.n137 VDD1.n91 8.92171
R234 VDD1.n56 VDD1.n13 8.14595
R235 VDD1.n45 VDD1.n17 8.14595
R236 VDD1.n125 VDD1.n97 8.14595
R237 VDD1.n136 VDD1.n93 8.14595
R238 VDD1.n53 VDD1.n52 7.3702
R239 VDD1.n49 VDD1.n48 7.3702
R240 VDD1.n129 VDD1.n128 7.3702
R241 VDD1.n133 VDD1.n132 7.3702
R242 VDD1.n52 VDD1.n15 6.59444
R243 VDD1.n49 VDD1.n15 6.59444
R244 VDD1.n129 VDD1.n95 6.59444
R245 VDD1.n132 VDD1.n95 6.59444
R246 VDD1.n53 VDD1.n13 5.81868
R247 VDD1.n48 VDD1.n17 5.81868
R248 VDD1.n128 VDD1.n97 5.81868
R249 VDD1.n133 VDD1.n93 5.81868
R250 VDD1.n57 VDD1.n56 5.04292
R251 VDD1.n45 VDD1.n44 5.04292
R252 VDD1.n125 VDD1.n124 5.04292
R253 VDD1.n137 VDD1.n136 5.04292
R254 VDD1.n60 VDD1.n11 4.26717
R255 VDD1.n41 VDD1.n19 4.26717
R256 VDD1.n121 VDD1.n99 4.26717
R257 VDD1.n140 VDD1.n91 4.26717
R258 VDD1.n30 VDD1.n26 3.70982
R259 VDD1.n110 VDD1.n106 3.70982
R260 VDD1.n61 VDD1.n9 3.49141
R261 VDD1.n40 VDD1.n21 3.49141
R262 VDD1.n120 VDD1.n101 3.49141
R263 VDD1.n141 VDD1.n89 3.49141
R264 VDD1.n65 VDD1.n64 2.71565
R265 VDD1.n37 VDD1.n36 2.71565
R266 VDD1.n117 VDD1.n116 2.71565
R267 VDD1.n145 VDD1.n144 2.71565
R268 VDD1.n164 VDD1.t0 2.19382
R269 VDD1.n164 VDD1.t3 2.19382
R270 VDD1.n162 VDD1.t1 2.19382
R271 VDD1.n162 VDD1.t4 2.19382
R272 VDD1.n80 VDD1.n0 1.93989
R273 VDD1.n68 VDD1.n6 1.93989
R274 VDD1.n33 VDD1.n23 1.93989
R275 VDD1.n113 VDD1.n103 1.93989
R276 VDD1.n149 VDD1.n87 1.93989
R277 VDD1.n161 VDD1.n81 1.93989
R278 VDD1.n78 VDD1.n77 1.16414
R279 VDD1.n69 VDD1.n4 1.16414
R280 VDD1.n32 VDD1.n25 1.16414
R281 VDD1.n112 VDD1.n105 1.16414
R282 VDD1.n150 VDD1.n85 1.16414
R283 VDD1.n159 VDD1.n158 1.16414
R284 VDD1 VDD1.n165 0.670759
R285 VDD1.n74 VDD1.n2 0.388379
R286 VDD1.n73 VDD1.n72 0.388379
R287 VDD1.n29 VDD1.n28 0.388379
R288 VDD1.n109 VDD1.n108 0.388379
R289 VDD1.n154 VDD1.n153 0.388379
R290 VDD1.n155 VDD1.n83 0.388379
R291 VDD1.n79 VDD1.n1 0.155672
R292 VDD1.n71 VDD1.n1 0.155672
R293 VDD1.n71 VDD1.n70 0.155672
R294 VDD1.n70 VDD1.n5 0.155672
R295 VDD1.n63 VDD1.n5 0.155672
R296 VDD1.n63 VDD1.n62 0.155672
R297 VDD1.n62 VDD1.n10 0.155672
R298 VDD1.n55 VDD1.n10 0.155672
R299 VDD1.n55 VDD1.n54 0.155672
R300 VDD1.n54 VDD1.n14 0.155672
R301 VDD1.n47 VDD1.n14 0.155672
R302 VDD1.n47 VDD1.n46 0.155672
R303 VDD1.n46 VDD1.n18 0.155672
R304 VDD1.n39 VDD1.n18 0.155672
R305 VDD1.n39 VDD1.n38 0.155672
R306 VDD1.n38 VDD1.n22 0.155672
R307 VDD1.n31 VDD1.n22 0.155672
R308 VDD1.n31 VDD1.n30 0.155672
R309 VDD1.n111 VDD1.n110 0.155672
R310 VDD1.n111 VDD1.n102 0.155672
R311 VDD1.n118 VDD1.n102 0.155672
R312 VDD1.n119 VDD1.n118 0.155672
R313 VDD1.n119 VDD1.n98 0.155672
R314 VDD1.n126 VDD1.n98 0.155672
R315 VDD1.n127 VDD1.n126 0.155672
R316 VDD1.n127 VDD1.n94 0.155672
R317 VDD1.n134 VDD1.n94 0.155672
R318 VDD1.n135 VDD1.n134 0.155672
R319 VDD1.n135 VDD1.n90 0.155672
R320 VDD1.n142 VDD1.n90 0.155672
R321 VDD1.n143 VDD1.n142 0.155672
R322 VDD1.n143 VDD1.n86 0.155672
R323 VDD1.n151 VDD1.n86 0.155672
R324 VDD1.n152 VDD1.n151 0.155672
R325 VDD1.n152 VDD1.n82 0.155672
R326 VDD1.n160 VDD1.n82 0.155672
R327 VTAIL.n330 VTAIL.n254 756.745
R328 VTAIL.n78 VTAIL.n2 756.745
R329 VTAIL.n248 VTAIL.n172 756.745
R330 VTAIL.n164 VTAIL.n88 756.745
R331 VTAIL.n281 VTAIL.n280 585
R332 VTAIL.n278 VTAIL.n277 585
R333 VTAIL.n287 VTAIL.n286 585
R334 VTAIL.n289 VTAIL.n288 585
R335 VTAIL.n274 VTAIL.n273 585
R336 VTAIL.n295 VTAIL.n294 585
R337 VTAIL.n297 VTAIL.n296 585
R338 VTAIL.n270 VTAIL.n269 585
R339 VTAIL.n303 VTAIL.n302 585
R340 VTAIL.n305 VTAIL.n304 585
R341 VTAIL.n266 VTAIL.n265 585
R342 VTAIL.n311 VTAIL.n310 585
R343 VTAIL.n313 VTAIL.n312 585
R344 VTAIL.n262 VTAIL.n261 585
R345 VTAIL.n319 VTAIL.n318 585
R346 VTAIL.n322 VTAIL.n321 585
R347 VTAIL.n320 VTAIL.n258 585
R348 VTAIL.n327 VTAIL.n257 585
R349 VTAIL.n329 VTAIL.n328 585
R350 VTAIL.n331 VTAIL.n330 585
R351 VTAIL.n29 VTAIL.n28 585
R352 VTAIL.n26 VTAIL.n25 585
R353 VTAIL.n35 VTAIL.n34 585
R354 VTAIL.n37 VTAIL.n36 585
R355 VTAIL.n22 VTAIL.n21 585
R356 VTAIL.n43 VTAIL.n42 585
R357 VTAIL.n45 VTAIL.n44 585
R358 VTAIL.n18 VTAIL.n17 585
R359 VTAIL.n51 VTAIL.n50 585
R360 VTAIL.n53 VTAIL.n52 585
R361 VTAIL.n14 VTAIL.n13 585
R362 VTAIL.n59 VTAIL.n58 585
R363 VTAIL.n61 VTAIL.n60 585
R364 VTAIL.n10 VTAIL.n9 585
R365 VTAIL.n67 VTAIL.n66 585
R366 VTAIL.n70 VTAIL.n69 585
R367 VTAIL.n68 VTAIL.n6 585
R368 VTAIL.n75 VTAIL.n5 585
R369 VTAIL.n77 VTAIL.n76 585
R370 VTAIL.n79 VTAIL.n78 585
R371 VTAIL.n249 VTAIL.n248 585
R372 VTAIL.n247 VTAIL.n246 585
R373 VTAIL.n245 VTAIL.n175 585
R374 VTAIL.n179 VTAIL.n176 585
R375 VTAIL.n240 VTAIL.n239 585
R376 VTAIL.n238 VTAIL.n237 585
R377 VTAIL.n181 VTAIL.n180 585
R378 VTAIL.n232 VTAIL.n231 585
R379 VTAIL.n230 VTAIL.n229 585
R380 VTAIL.n185 VTAIL.n184 585
R381 VTAIL.n224 VTAIL.n223 585
R382 VTAIL.n222 VTAIL.n221 585
R383 VTAIL.n189 VTAIL.n188 585
R384 VTAIL.n216 VTAIL.n215 585
R385 VTAIL.n214 VTAIL.n213 585
R386 VTAIL.n193 VTAIL.n192 585
R387 VTAIL.n208 VTAIL.n207 585
R388 VTAIL.n206 VTAIL.n205 585
R389 VTAIL.n197 VTAIL.n196 585
R390 VTAIL.n200 VTAIL.n199 585
R391 VTAIL.n165 VTAIL.n164 585
R392 VTAIL.n163 VTAIL.n162 585
R393 VTAIL.n161 VTAIL.n91 585
R394 VTAIL.n95 VTAIL.n92 585
R395 VTAIL.n156 VTAIL.n155 585
R396 VTAIL.n154 VTAIL.n153 585
R397 VTAIL.n97 VTAIL.n96 585
R398 VTAIL.n148 VTAIL.n147 585
R399 VTAIL.n146 VTAIL.n145 585
R400 VTAIL.n101 VTAIL.n100 585
R401 VTAIL.n140 VTAIL.n139 585
R402 VTAIL.n138 VTAIL.n137 585
R403 VTAIL.n105 VTAIL.n104 585
R404 VTAIL.n132 VTAIL.n131 585
R405 VTAIL.n130 VTAIL.n129 585
R406 VTAIL.n109 VTAIL.n108 585
R407 VTAIL.n124 VTAIL.n123 585
R408 VTAIL.n122 VTAIL.n121 585
R409 VTAIL.n113 VTAIL.n112 585
R410 VTAIL.n116 VTAIL.n115 585
R411 VTAIL.t9 VTAIL.n198 327.466
R412 VTAIL.t2 VTAIL.n114 327.466
R413 VTAIL.t3 VTAIL.n279 327.466
R414 VTAIL.t7 VTAIL.n27 327.466
R415 VTAIL.n280 VTAIL.n277 171.744
R416 VTAIL.n287 VTAIL.n277 171.744
R417 VTAIL.n288 VTAIL.n287 171.744
R418 VTAIL.n288 VTAIL.n273 171.744
R419 VTAIL.n295 VTAIL.n273 171.744
R420 VTAIL.n296 VTAIL.n295 171.744
R421 VTAIL.n296 VTAIL.n269 171.744
R422 VTAIL.n303 VTAIL.n269 171.744
R423 VTAIL.n304 VTAIL.n303 171.744
R424 VTAIL.n304 VTAIL.n265 171.744
R425 VTAIL.n311 VTAIL.n265 171.744
R426 VTAIL.n312 VTAIL.n311 171.744
R427 VTAIL.n312 VTAIL.n261 171.744
R428 VTAIL.n319 VTAIL.n261 171.744
R429 VTAIL.n321 VTAIL.n319 171.744
R430 VTAIL.n321 VTAIL.n320 171.744
R431 VTAIL.n320 VTAIL.n257 171.744
R432 VTAIL.n329 VTAIL.n257 171.744
R433 VTAIL.n330 VTAIL.n329 171.744
R434 VTAIL.n28 VTAIL.n25 171.744
R435 VTAIL.n35 VTAIL.n25 171.744
R436 VTAIL.n36 VTAIL.n35 171.744
R437 VTAIL.n36 VTAIL.n21 171.744
R438 VTAIL.n43 VTAIL.n21 171.744
R439 VTAIL.n44 VTAIL.n43 171.744
R440 VTAIL.n44 VTAIL.n17 171.744
R441 VTAIL.n51 VTAIL.n17 171.744
R442 VTAIL.n52 VTAIL.n51 171.744
R443 VTAIL.n52 VTAIL.n13 171.744
R444 VTAIL.n59 VTAIL.n13 171.744
R445 VTAIL.n60 VTAIL.n59 171.744
R446 VTAIL.n60 VTAIL.n9 171.744
R447 VTAIL.n67 VTAIL.n9 171.744
R448 VTAIL.n69 VTAIL.n67 171.744
R449 VTAIL.n69 VTAIL.n68 171.744
R450 VTAIL.n68 VTAIL.n5 171.744
R451 VTAIL.n77 VTAIL.n5 171.744
R452 VTAIL.n78 VTAIL.n77 171.744
R453 VTAIL.n248 VTAIL.n247 171.744
R454 VTAIL.n247 VTAIL.n175 171.744
R455 VTAIL.n179 VTAIL.n175 171.744
R456 VTAIL.n239 VTAIL.n179 171.744
R457 VTAIL.n239 VTAIL.n238 171.744
R458 VTAIL.n238 VTAIL.n180 171.744
R459 VTAIL.n231 VTAIL.n180 171.744
R460 VTAIL.n231 VTAIL.n230 171.744
R461 VTAIL.n230 VTAIL.n184 171.744
R462 VTAIL.n223 VTAIL.n184 171.744
R463 VTAIL.n223 VTAIL.n222 171.744
R464 VTAIL.n222 VTAIL.n188 171.744
R465 VTAIL.n215 VTAIL.n188 171.744
R466 VTAIL.n215 VTAIL.n214 171.744
R467 VTAIL.n214 VTAIL.n192 171.744
R468 VTAIL.n207 VTAIL.n192 171.744
R469 VTAIL.n207 VTAIL.n206 171.744
R470 VTAIL.n206 VTAIL.n196 171.744
R471 VTAIL.n199 VTAIL.n196 171.744
R472 VTAIL.n164 VTAIL.n163 171.744
R473 VTAIL.n163 VTAIL.n91 171.744
R474 VTAIL.n95 VTAIL.n91 171.744
R475 VTAIL.n155 VTAIL.n95 171.744
R476 VTAIL.n155 VTAIL.n154 171.744
R477 VTAIL.n154 VTAIL.n96 171.744
R478 VTAIL.n147 VTAIL.n96 171.744
R479 VTAIL.n147 VTAIL.n146 171.744
R480 VTAIL.n146 VTAIL.n100 171.744
R481 VTAIL.n139 VTAIL.n100 171.744
R482 VTAIL.n139 VTAIL.n138 171.744
R483 VTAIL.n138 VTAIL.n104 171.744
R484 VTAIL.n131 VTAIL.n104 171.744
R485 VTAIL.n131 VTAIL.n130 171.744
R486 VTAIL.n130 VTAIL.n108 171.744
R487 VTAIL.n123 VTAIL.n108 171.744
R488 VTAIL.n123 VTAIL.n122 171.744
R489 VTAIL.n122 VTAIL.n112 171.744
R490 VTAIL.n115 VTAIL.n112 171.744
R491 VTAIL.n280 VTAIL.t3 85.8723
R492 VTAIL.n28 VTAIL.t7 85.8723
R493 VTAIL.n199 VTAIL.t9 85.8723
R494 VTAIL.n115 VTAIL.t2 85.8723
R495 VTAIL.n171 VTAIL.n170 57.5787
R496 VTAIL.n87 VTAIL.n86 57.5787
R497 VTAIL.n1 VTAIL.n0 57.5785
R498 VTAIL.n85 VTAIL.n84 57.5785
R499 VTAIL.n335 VTAIL.n334 35.6763
R500 VTAIL.n83 VTAIL.n82 35.6763
R501 VTAIL.n253 VTAIL.n252 35.6763
R502 VTAIL.n169 VTAIL.n168 35.6763
R503 VTAIL.n87 VTAIL.n85 30.9703
R504 VTAIL.n335 VTAIL.n253 28.0565
R505 VTAIL.n281 VTAIL.n279 16.3895
R506 VTAIL.n29 VTAIL.n27 16.3895
R507 VTAIL.n200 VTAIL.n198 16.3895
R508 VTAIL.n116 VTAIL.n114 16.3895
R509 VTAIL.n328 VTAIL.n327 13.1884
R510 VTAIL.n76 VTAIL.n75 13.1884
R511 VTAIL.n246 VTAIL.n245 13.1884
R512 VTAIL.n162 VTAIL.n161 13.1884
R513 VTAIL.n282 VTAIL.n278 12.8005
R514 VTAIL.n326 VTAIL.n258 12.8005
R515 VTAIL.n331 VTAIL.n256 12.8005
R516 VTAIL.n30 VTAIL.n26 12.8005
R517 VTAIL.n74 VTAIL.n6 12.8005
R518 VTAIL.n79 VTAIL.n4 12.8005
R519 VTAIL.n249 VTAIL.n174 12.8005
R520 VTAIL.n244 VTAIL.n176 12.8005
R521 VTAIL.n201 VTAIL.n197 12.8005
R522 VTAIL.n165 VTAIL.n90 12.8005
R523 VTAIL.n160 VTAIL.n92 12.8005
R524 VTAIL.n117 VTAIL.n113 12.8005
R525 VTAIL.n286 VTAIL.n285 12.0247
R526 VTAIL.n323 VTAIL.n322 12.0247
R527 VTAIL.n332 VTAIL.n254 12.0247
R528 VTAIL.n34 VTAIL.n33 12.0247
R529 VTAIL.n71 VTAIL.n70 12.0247
R530 VTAIL.n80 VTAIL.n2 12.0247
R531 VTAIL.n250 VTAIL.n172 12.0247
R532 VTAIL.n241 VTAIL.n240 12.0247
R533 VTAIL.n205 VTAIL.n204 12.0247
R534 VTAIL.n166 VTAIL.n88 12.0247
R535 VTAIL.n157 VTAIL.n156 12.0247
R536 VTAIL.n121 VTAIL.n120 12.0247
R537 VTAIL.n289 VTAIL.n276 11.249
R538 VTAIL.n318 VTAIL.n260 11.249
R539 VTAIL.n37 VTAIL.n24 11.249
R540 VTAIL.n66 VTAIL.n8 11.249
R541 VTAIL.n237 VTAIL.n178 11.249
R542 VTAIL.n208 VTAIL.n195 11.249
R543 VTAIL.n153 VTAIL.n94 11.249
R544 VTAIL.n124 VTAIL.n111 11.249
R545 VTAIL.n290 VTAIL.n274 10.4732
R546 VTAIL.n317 VTAIL.n262 10.4732
R547 VTAIL.n38 VTAIL.n22 10.4732
R548 VTAIL.n65 VTAIL.n10 10.4732
R549 VTAIL.n236 VTAIL.n181 10.4732
R550 VTAIL.n209 VTAIL.n193 10.4732
R551 VTAIL.n152 VTAIL.n97 10.4732
R552 VTAIL.n125 VTAIL.n109 10.4732
R553 VTAIL.n294 VTAIL.n293 9.69747
R554 VTAIL.n314 VTAIL.n313 9.69747
R555 VTAIL.n42 VTAIL.n41 9.69747
R556 VTAIL.n62 VTAIL.n61 9.69747
R557 VTAIL.n233 VTAIL.n232 9.69747
R558 VTAIL.n213 VTAIL.n212 9.69747
R559 VTAIL.n149 VTAIL.n148 9.69747
R560 VTAIL.n129 VTAIL.n128 9.69747
R561 VTAIL.n334 VTAIL.n333 9.45567
R562 VTAIL.n82 VTAIL.n81 9.45567
R563 VTAIL.n252 VTAIL.n251 9.45567
R564 VTAIL.n168 VTAIL.n167 9.45567
R565 VTAIL.n333 VTAIL.n332 9.3005
R566 VTAIL.n256 VTAIL.n255 9.3005
R567 VTAIL.n301 VTAIL.n300 9.3005
R568 VTAIL.n299 VTAIL.n298 9.3005
R569 VTAIL.n272 VTAIL.n271 9.3005
R570 VTAIL.n293 VTAIL.n292 9.3005
R571 VTAIL.n291 VTAIL.n290 9.3005
R572 VTAIL.n276 VTAIL.n275 9.3005
R573 VTAIL.n285 VTAIL.n284 9.3005
R574 VTAIL.n283 VTAIL.n282 9.3005
R575 VTAIL.n268 VTAIL.n267 9.3005
R576 VTAIL.n307 VTAIL.n306 9.3005
R577 VTAIL.n309 VTAIL.n308 9.3005
R578 VTAIL.n264 VTAIL.n263 9.3005
R579 VTAIL.n315 VTAIL.n314 9.3005
R580 VTAIL.n317 VTAIL.n316 9.3005
R581 VTAIL.n260 VTAIL.n259 9.3005
R582 VTAIL.n324 VTAIL.n323 9.3005
R583 VTAIL.n326 VTAIL.n325 9.3005
R584 VTAIL.n81 VTAIL.n80 9.3005
R585 VTAIL.n4 VTAIL.n3 9.3005
R586 VTAIL.n49 VTAIL.n48 9.3005
R587 VTAIL.n47 VTAIL.n46 9.3005
R588 VTAIL.n20 VTAIL.n19 9.3005
R589 VTAIL.n41 VTAIL.n40 9.3005
R590 VTAIL.n39 VTAIL.n38 9.3005
R591 VTAIL.n24 VTAIL.n23 9.3005
R592 VTAIL.n33 VTAIL.n32 9.3005
R593 VTAIL.n31 VTAIL.n30 9.3005
R594 VTAIL.n16 VTAIL.n15 9.3005
R595 VTAIL.n55 VTAIL.n54 9.3005
R596 VTAIL.n57 VTAIL.n56 9.3005
R597 VTAIL.n12 VTAIL.n11 9.3005
R598 VTAIL.n63 VTAIL.n62 9.3005
R599 VTAIL.n65 VTAIL.n64 9.3005
R600 VTAIL.n8 VTAIL.n7 9.3005
R601 VTAIL.n72 VTAIL.n71 9.3005
R602 VTAIL.n74 VTAIL.n73 9.3005
R603 VTAIL.n226 VTAIL.n225 9.3005
R604 VTAIL.n228 VTAIL.n227 9.3005
R605 VTAIL.n183 VTAIL.n182 9.3005
R606 VTAIL.n234 VTAIL.n233 9.3005
R607 VTAIL.n236 VTAIL.n235 9.3005
R608 VTAIL.n178 VTAIL.n177 9.3005
R609 VTAIL.n242 VTAIL.n241 9.3005
R610 VTAIL.n244 VTAIL.n243 9.3005
R611 VTAIL.n251 VTAIL.n250 9.3005
R612 VTAIL.n174 VTAIL.n173 9.3005
R613 VTAIL.n187 VTAIL.n186 9.3005
R614 VTAIL.n220 VTAIL.n219 9.3005
R615 VTAIL.n218 VTAIL.n217 9.3005
R616 VTAIL.n191 VTAIL.n190 9.3005
R617 VTAIL.n212 VTAIL.n211 9.3005
R618 VTAIL.n210 VTAIL.n209 9.3005
R619 VTAIL.n195 VTAIL.n194 9.3005
R620 VTAIL.n204 VTAIL.n203 9.3005
R621 VTAIL.n202 VTAIL.n201 9.3005
R622 VTAIL.n142 VTAIL.n141 9.3005
R623 VTAIL.n144 VTAIL.n143 9.3005
R624 VTAIL.n99 VTAIL.n98 9.3005
R625 VTAIL.n150 VTAIL.n149 9.3005
R626 VTAIL.n152 VTAIL.n151 9.3005
R627 VTAIL.n94 VTAIL.n93 9.3005
R628 VTAIL.n158 VTAIL.n157 9.3005
R629 VTAIL.n160 VTAIL.n159 9.3005
R630 VTAIL.n167 VTAIL.n166 9.3005
R631 VTAIL.n90 VTAIL.n89 9.3005
R632 VTAIL.n103 VTAIL.n102 9.3005
R633 VTAIL.n136 VTAIL.n135 9.3005
R634 VTAIL.n134 VTAIL.n133 9.3005
R635 VTAIL.n107 VTAIL.n106 9.3005
R636 VTAIL.n128 VTAIL.n127 9.3005
R637 VTAIL.n126 VTAIL.n125 9.3005
R638 VTAIL.n111 VTAIL.n110 9.3005
R639 VTAIL.n120 VTAIL.n119 9.3005
R640 VTAIL.n118 VTAIL.n117 9.3005
R641 VTAIL.n297 VTAIL.n272 8.92171
R642 VTAIL.n310 VTAIL.n264 8.92171
R643 VTAIL.n45 VTAIL.n20 8.92171
R644 VTAIL.n58 VTAIL.n12 8.92171
R645 VTAIL.n229 VTAIL.n183 8.92171
R646 VTAIL.n216 VTAIL.n191 8.92171
R647 VTAIL.n145 VTAIL.n99 8.92171
R648 VTAIL.n132 VTAIL.n107 8.92171
R649 VTAIL.n298 VTAIL.n270 8.14595
R650 VTAIL.n309 VTAIL.n266 8.14595
R651 VTAIL.n46 VTAIL.n18 8.14595
R652 VTAIL.n57 VTAIL.n14 8.14595
R653 VTAIL.n228 VTAIL.n185 8.14595
R654 VTAIL.n217 VTAIL.n189 8.14595
R655 VTAIL.n144 VTAIL.n101 8.14595
R656 VTAIL.n133 VTAIL.n105 8.14595
R657 VTAIL.n302 VTAIL.n301 7.3702
R658 VTAIL.n306 VTAIL.n305 7.3702
R659 VTAIL.n50 VTAIL.n49 7.3702
R660 VTAIL.n54 VTAIL.n53 7.3702
R661 VTAIL.n225 VTAIL.n224 7.3702
R662 VTAIL.n221 VTAIL.n220 7.3702
R663 VTAIL.n141 VTAIL.n140 7.3702
R664 VTAIL.n137 VTAIL.n136 7.3702
R665 VTAIL.n302 VTAIL.n268 6.59444
R666 VTAIL.n305 VTAIL.n268 6.59444
R667 VTAIL.n50 VTAIL.n16 6.59444
R668 VTAIL.n53 VTAIL.n16 6.59444
R669 VTAIL.n224 VTAIL.n187 6.59444
R670 VTAIL.n221 VTAIL.n187 6.59444
R671 VTAIL.n140 VTAIL.n103 6.59444
R672 VTAIL.n137 VTAIL.n103 6.59444
R673 VTAIL.n301 VTAIL.n270 5.81868
R674 VTAIL.n306 VTAIL.n266 5.81868
R675 VTAIL.n49 VTAIL.n18 5.81868
R676 VTAIL.n54 VTAIL.n14 5.81868
R677 VTAIL.n225 VTAIL.n185 5.81868
R678 VTAIL.n220 VTAIL.n189 5.81868
R679 VTAIL.n141 VTAIL.n101 5.81868
R680 VTAIL.n136 VTAIL.n105 5.81868
R681 VTAIL.n298 VTAIL.n297 5.04292
R682 VTAIL.n310 VTAIL.n309 5.04292
R683 VTAIL.n46 VTAIL.n45 5.04292
R684 VTAIL.n58 VTAIL.n57 5.04292
R685 VTAIL.n229 VTAIL.n228 5.04292
R686 VTAIL.n217 VTAIL.n216 5.04292
R687 VTAIL.n145 VTAIL.n144 5.04292
R688 VTAIL.n133 VTAIL.n132 5.04292
R689 VTAIL.n294 VTAIL.n272 4.26717
R690 VTAIL.n313 VTAIL.n264 4.26717
R691 VTAIL.n42 VTAIL.n20 4.26717
R692 VTAIL.n61 VTAIL.n12 4.26717
R693 VTAIL.n232 VTAIL.n183 4.26717
R694 VTAIL.n213 VTAIL.n191 4.26717
R695 VTAIL.n148 VTAIL.n99 4.26717
R696 VTAIL.n129 VTAIL.n107 4.26717
R697 VTAIL.n283 VTAIL.n279 3.70982
R698 VTAIL.n31 VTAIL.n27 3.70982
R699 VTAIL.n202 VTAIL.n198 3.70982
R700 VTAIL.n118 VTAIL.n114 3.70982
R701 VTAIL.n293 VTAIL.n274 3.49141
R702 VTAIL.n314 VTAIL.n262 3.49141
R703 VTAIL.n41 VTAIL.n22 3.49141
R704 VTAIL.n62 VTAIL.n10 3.49141
R705 VTAIL.n233 VTAIL.n181 3.49141
R706 VTAIL.n212 VTAIL.n193 3.49141
R707 VTAIL.n149 VTAIL.n97 3.49141
R708 VTAIL.n128 VTAIL.n109 3.49141
R709 VTAIL.n169 VTAIL.n87 2.91429
R710 VTAIL.n253 VTAIL.n171 2.91429
R711 VTAIL.n85 VTAIL.n83 2.91429
R712 VTAIL.n290 VTAIL.n289 2.71565
R713 VTAIL.n318 VTAIL.n317 2.71565
R714 VTAIL.n38 VTAIL.n37 2.71565
R715 VTAIL.n66 VTAIL.n65 2.71565
R716 VTAIL.n237 VTAIL.n236 2.71565
R717 VTAIL.n209 VTAIL.n208 2.71565
R718 VTAIL.n153 VTAIL.n152 2.71565
R719 VTAIL.n125 VTAIL.n124 2.71565
R720 VTAIL.n0 VTAIL.t4 2.19382
R721 VTAIL.n0 VTAIL.t0 2.19382
R722 VTAIL.n84 VTAIL.t8 2.19382
R723 VTAIL.n84 VTAIL.t11 2.19382
R724 VTAIL.n170 VTAIL.t10 2.19382
R725 VTAIL.n170 VTAIL.t6 2.19382
R726 VTAIL.n86 VTAIL.t1 2.19382
R727 VTAIL.n86 VTAIL.t5 2.19382
R728 VTAIL VTAIL.n335 2.12766
R729 VTAIL.n286 VTAIL.n276 1.93989
R730 VTAIL.n322 VTAIL.n260 1.93989
R731 VTAIL.n334 VTAIL.n254 1.93989
R732 VTAIL.n34 VTAIL.n24 1.93989
R733 VTAIL.n70 VTAIL.n8 1.93989
R734 VTAIL.n82 VTAIL.n2 1.93989
R735 VTAIL.n252 VTAIL.n172 1.93989
R736 VTAIL.n240 VTAIL.n178 1.93989
R737 VTAIL.n205 VTAIL.n195 1.93989
R738 VTAIL.n168 VTAIL.n88 1.93989
R739 VTAIL.n156 VTAIL.n94 1.93989
R740 VTAIL.n121 VTAIL.n111 1.93989
R741 VTAIL.n171 VTAIL.n169 1.92722
R742 VTAIL.n83 VTAIL.n1 1.92722
R743 VTAIL.n285 VTAIL.n278 1.16414
R744 VTAIL.n323 VTAIL.n258 1.16414
R745 VTAIL.n332 VTAIL.n331 1.16414
R746 VTAIL.n33 VTAIL.n26 1.16414
R747 VTAIL.n71 VTAIL.n6 1.16414
R748 VTAIL.n80 VTAIL.n79 1.16414
R749 VTAIL.n250 VTAIL.n249 1.16414
R750 VTAIL.n241 VTAIL.n176 1.16414
R751 VTAIL.n204 VTAIL.n197 1.16414
R752 VTAIL.n166 VTAIL.n165 1.16414
R753 VTAIL.n157 VTAIL.n92 1.16414
R754 VTAIL.n120 VTAIL.n113 1.16414
R755 VTAIL VTAIL.n1 0.787138
R756 VTAIL.n282 VTAIL.n281 0.388379
R757 VTAIL.n327 VTAIL.n326 0.388379
R758 VTAIL.n328 VTAIL.n256 0.388379
R759 VTAIL.n30 VTAIL.n29 0.388379
R760 VTAIL.n75 VTAIL.n74 0.388379
R761 VTAIL.n76 VTAIL.n4 0.388379
R762 VTAIL.n246 VTAIL.n174 0.388379
R763 VTAIL.n245 VTAIL.n244 0.388379
R764 VTAIL.n201 VTAIL.n200 0.388379
R765 VTAIL.n162 VTAIL.n90 0.388379
R766 VTAIL.n161 VTAIL.n160 0.388379
R767 VTAIL.n117 VTAIL.n116 0.388379
R768 VTAIL.n284 VTAIL.n283 0.155672
R769 VTAIL.n284 VTAIL.n275 0.155672
R770 VTAIL.n291 VTAIL.n275 0.155672
R771 VTAIL.n292 VTAIL.n291 0.155672
R772 VTAIL.n292 VTAIL.n271 0.155672
R773 VTAIL.n299 VTAIL.n271 0.155672
R774 VTAIL.n300 VTAIL.n299 0.155672
R775 VTAIL.n300 VTAIL.n267 0.155672
R776 VTAIL.n307 VTAIL.n267 0.155672
R777 VTAIL.n308 VTAIL.n307 0.155672
R778 VTAIL.n308 VTAIL.n263 0.155672
R779 VTAIL.n315 VTAIL.n263 0.155672
R780 VTAIL.n316 VTAIL.n315 0.155672
R781 VTAIL.n316 VTAIL.n259 0.155672
R782 VTAIL.n324 VTAIL.n259 0.155672
R783 VTAIL.n325 VTAIL.n324 0.155672
R784 VTAIL.n325 VTAIL.n255 0.155672
R785 VTAIL.n333 VTAIL.n255 0.155672
R786 VTAIL.n32 VTAIL.n31 0.155672
R787 VTAIL.n32 VTAIL.n23 0.155672
R788 VTAIL.n39 VTAIL.n23 0.155672
R789 VTAIL.n40 VTAIL.n39 0.155672
R790 VTAIL.n40 VTAIL.n19 0.155672
R791 VTAIL.n47 VTAIL.n19 0.155672
R792 VTAIL.n48 VTAIL.n47 0.155672
R793 VTAIL.n48 VTAIL.n15 0.155672
R794 VTAIL.n55 VTAIL.n15 0.155672
R795 VTAIL.n56 VTAIL.n55 0.155672
R796 VTAIL.n56 VTAIL.n11 0.155672
R797 VTAIL.n63 VTAIL.n11 0.155672
R798 VTAIL.n64 VTAIL.n63 0.155672
R799 VTAIL.n64 VTAIL.n7 0.155672
R800 VTAIL.n72 VTAIL.n7 0.155672
R801 VTAIL.n73 VTAIL.n72 0.155672
R802 VTAIL.n73 VTAIL.n3 0.155672
R803 VTAIL.n81 VTAIL.n3 0.155672
R804 VTAIL.n251 VTAIL.n173 0.155672
R805 VTAIL.n243 VTAIL.n173 0.155672
R806 VTAIL.n243 VTAIL.n242 0.155672
R807 VTAIL.n242 VTAIL.n177 0.155672
R808 VTAIL.n235 VTAIL.n177 0.155672
R809 VTAIL.n235 VTAIL.n234 0.155672
R810 VTAIL.n234 VTAIL.n182 0.155672
R811 VTAIL.n227 VTAIL.n182 0.155672
R812 VTAIL.n227 VTAIL.n226 0.155672
R813 VTAIL.n226 VTAIL.n186 0.155672
R814 VTAIL.n219 VTAIL.n186 0.155672
R815 VTAIL.n219 VTAIL.n218 0.155672
R816 VTAIL.n218 VTAIL.n190 0.155672
R817 VTAIL.n211 VTAIL.n190 0.155672
R818 VTAIL.n211 VTAIL.n210 0.155672
R819 VTAIL.n210 VTAIL.n194 0.155672
R820 VTAIL.n203 VTAIL.n194 0.155672
R821 VTAIL.n203 VTAIL.n202 0.155672
R822 VTAIL.n167 VTAIL.n89 0.155672
R823 VTAIL.n159 VTAIL.n89 0.155672
R824 VTAIL.n159 VTAIL.n158 0.155672
R825 VTAIL.n158 VTAIL.n93 0.155672
R826 VTAIL.n151 VTAIL.n93 0.155672
R827 VTAIL.n151 VTAIL.n150 0.155672
R828 VTAIL.n150 VTAIL.n98 0.155672
R829 VTAIL.n143 VTAIL.n98 0.155672
R830 VTAIL.n143 VTAIL.n142 0.155672
R831 VTAIL.n142 VTAIL.n102 0.155672
R832 VTAIL.n135 VTAIL.n102 0.155672
R833 VTAIL.n135 VTAIL.n134 0.155672
R834 VTAIL.n134 VTAIL.n106 0.155672
R835 VTAIL.n127 VTAIL.n106 0.155672
R836 VTAIL.n127 VTAIL.n126 0.155672
R837 VTAIL.n126 VTAIL.n110 0.155672
R838 VTAIL.n119 VTAIL.n110 0.155672
R839 VTAIL.n119 VTAIL.n118 0.155672
R840 VN.n30 VN.n29 161.3
R841 VN.n28 VN.n17 161.3
R842 VN.n27 VN.n26 161.3
R843 VN.n25 VN.n18 161.3
R844 VN.n24 VN.n23 161.3
R845 VN.n22 VN.n19 161.3
R846 VN.n14 VN.n13 161.3
R847 VN.n12 VN.n1 161.3
R848 VN.n11 VN.n10 161.3
R849 VN.n9 VN.n2 161.3
R850 VN.n8 VN.n7 161.3
R851 VN.n6 VN.n3 161.3
R852 VN.n20 VN.t2 150.538
R853 VN.n4 VN.t1 150.538
R854 VN.n5 VN.t4 117.103
R855 VN.n0 VN.t3 117.103
R856 VN.n21 VN.t0 117.103
R857 VN.n16 VN.t5 117.103
R858 VN.n15 VN.n0 71.5558
R859 VN.n31 VN.n16 71.5558
R860 VN.n11 VN.n2 56.5617
R861 VN.n27 VN.n18 56.5617
R862 VN VN.n31 52.8542
R863 VN.n5 VN.n4 49.4409
R864 VN.n21 VN.n20 49.4409
R865 VN.n6 VN.n5 24.5923
R866 VN.n7 VN.n6 24.5923
R867 VN.n7 VN.n2 24.5923
R868 VN.n12 VN.n11 24.5923
R869 VN.n13 VN.n12 24.5923
R870 VN.n23 VN.n18 24.5923
R871 VN.n23 VN.n22 24.5923
R872 VN.n22 VN.n21 24.5923
R873 VN.n29 VN.n28 24.5923
R874 VN.n28 VN.n27 24.5923
R875 VN.n13 VN.n0 18.6903
R876 VN.n29 VN.n16 18.6903
R877 VN.n4 VN.n3 3.96753
R878 VN.n20 VN.n19 3.96753
R879 VN.n31 VN.n30 0.354861
R880 VN.n15 VN.n14 0.354861
R881 VN VN.n15 0.267071
R882 VN.n30 VN.n17 0.189894
R883 VN.n26 VN.n17 0.189894
R884 VN.n26 VN.n25 0.189894
R885 VN.n25 VN.n24 0.189894
R886 VN.n24 VN.n19 0.189894
R887 VN.n8 VN.n3 0.189894
R888 VN.n9 VN.n8 0.189894
R889 VN.n10 VN.n9 0.189894
R890 VN.n10 VN.n1 0.189894
R891 VN.n14 VN.n1 0.189894
R892 VDD2.n159 VDD2.n83 756.745
R893 VDD2.n76 VDD2.n0 756.745
R894 VDD2.n160 VDD2.n159 585
R895 VDD2.n158 VDD2.n157 585
R896 VDD2.n156 VDD2.n86 585
R897 VDD2.n90 VDD2.n87 585
R898 VDD2.n151 VDD2.n150 585
R899 VDD2.n149 VDD2.n148 585
R900 VDD2.n92 VDD2.n91 585
R901 VDD2.n143 VDD2.n142 585
R902 VDD2.n141 VDD2.n140 585
R903 VDD2.n96 VDD2.n95 585
R904 VDD2.n135 VDD2.n134 585
R905 VDD2.n133 VDD2.n132 585
R906 VDD2.n100 VDD2.n99 585
R907 VDD2.n127 VDD2.n126 585
R908 VDD2.n125 VDD2.n124 585
R909 VDD2.n104 VDD2.n103 585
R910 VDD2.n119 VDD2.n118 585
R911 VDD2.n117 VDD2.n116 585
R912 VDD2.n108 VDD2.n107 585
R913 VDD2.n111 VDD2.n110 585
R914 VDD2.n27 VDD2.n26 585
R915 VDD2.n24 VDD2.n23 585
R916 VDD2.n33 VDD2.n32 585
R917 VDD2.n35 VDD2.n34 585
R918 VDD2.n20 VDD2.n19 585
R919 VDD2.n41 VDD2.n40 585
R920 VDD2.n43 VDD2.n42 585
R921 VDD2.n16 VDD2.n15 585
R922 VDD2.n49 VDD2.n48 585
R923 VDD2.n51 VDD2.n50 585
R924 VDD2.n12 VDD2.n11 585
R925 VDD2.n57 VDD2.n56 585
R926 VDD2.n59 VDD2.n58 585
R927 VDD2.n8 VDD2.n7 585
R928 VDD2.n65 VDD2.n64 585
R929 VDD2.n68 VDD2.n67 585
R930 VDD2.n66 VDD2.n4 585
R931 VDD2.n73 VDD2.n3 585
R932 VDD2.n75 VDD2.n74 585
R933 VDD2.n77 VDD2.n76 585
R934 VDD2.t0 VDD2.n109 327.466
R935 VDD2.t4 VDD2.n25 327.466
R936 VDD2.n159 VDD2.n158 171.744
R937 VDD2.n158 VDD2.n86 171.744
R938 VDD2.n90 VDD2.n86 171.744
R939 VDD2.n150 VDD2.n90 171.744
R940 VDD2.n150 VDD2.n149 171.744
R941 VDD2.n149 VDD2.n91 171.744
R942 VDD2.n142 VDD2.n91 171.744
R943 VDD2.n142 VDD2.n141 171.744
R944 VDD2.n141 VDD2.n95 171.744
R945 VDD2.n134 VDD2.n95 171.744
R946 VDD2.n134 VDD2.n133 171.744
R947 VDD2.n133 VDD2.n99 171.744
R948 VDD2.n126 VDD2.n99 171.744
R949 VDD2.n126 VDD2.n125 171.744
R950 VDD2.n125 VDD2.n103 171.744
R951 VDD2.n118 VDD2.n103 171.744
R952 VDD2.n118 VDD2.n117 171.744
R953 VDD2.n117 VDD2.n107 171.744
R954 VDD2.n110 VDD2.n107 171.744
R955 VDD2.n26 VDD2.n23 171.744
R956 VDD2.n33 VDD2.n23 171.744
R957 VDD2.n34 VDD2.n33 171.744
R958 VDD2.n34 VDD2.n19 171.744
R959 VDD2.n41 VDD2.n19 171.744
R960 VDD2.n42 VDD2.n41 171.744
R961 VDD2.n42 VDD2.n15 171.744
R962 VDD2.n49 VDD2.n15 171.744
R963 VDD2.n50 VDD2.n49 171.744
R964 VDD2.n50 VDD2.n11 171.744
R965 VDD2.n57 VDD2.n11 171.744
R966 VDD2.n58 VDD2.n57 171.744
R967 VDD2.n58 VDD2.n7 171.744
R968 VDD2.n65 VDD2.n7 171.744
R969 VDD2.n67 VDD2.n65 171.744
R970 VDD2.n67 VDD2.n66 171.744
R971 VDD2.n66 VDD2.n3 171.744
R972 VDD2.n75 VDD2.n3 171.744
R973 VDD2.n76 VDD2.n75 171.744
R974 VDD2.n110 VDD2.t0 85.8723
R975 VDD2.n26 VDD2.t4 85.8723
R976 VDD2.n82 VDD2.n81 74.9304
R977 VDD2 VDD2.n165 74.9275
R978 VDD2.n82 VDD2.n80 54.485
R979 VDD2.n164 VDD2.n163 52.355
R980 VDD2.n164 VDD2.n82 45.961
R981 VDD2.n111 VDD2.n109 16.3895
R982 VDD2.n27 VDD2.n25 16.3895
R983 VDD2.n157 VDD2.n156 13.1884
R984 VDD2.n74 VDD2.n73 13.1884
R985 VDD2.n160 VDD2.n85 12.8005
R986 VDD2.n155 VDD2.n87 12.8005
R987 VDD2.n112 VDD2.n108 12.8005
R988 VDD2.n28 VDD2.n24 12.8005
R989 VDD2.n72 VDD2.n4 12.8005
R990 VDD2.n77 VDD2.n2 12.8005
R991 VDD2.n161 VDD2.n83 12.0247
R992 VDD2.n152 VDD2.n151 12.0247
R993 VDD2.n116 VDD2.n115 12.0247
R994 VDD2.n32 VDD2.n31 12.0247
R995 VDD2.n69 VDD2.n68 12.0247
R996 VDD2.n78 VDD2.n0 12.0247
R997 VDD2.n148 VDD2.n89 11.249
R998 VDD2.n119 VDD2.n106 11.249
R999 VDD2.n35 VDD2.n22 11.249
R1000 VDD2.n64 VDD2.n6 11.249
R1001 VDD2.n147 VDD2.n92 10.4732
R1002 VDD2.n120 VDD2.n104 10.4732
R1003 VDD2.n36 VDD2.n20 10.4732
R1004 VDD2.n63 VDD2.n8 10.4732
R1005 VDD2.n144 VDD2.n143 9.69747
R1006 VDD2.n124 VDD2.n123 9.69747
R1007 VDD2.n40 VDD2.n39 9.69747
R1008 VDD2.n60 VDD2.n59 9.69747
R1009 VDD2.n163 VDD2.n162 9.45567
R1010 VDD2.n80 VDD2.n79 9.45567
R1011 VDD2.n137 VDD2.n136 9.3005
R1012 VDD2.n139 VDD2.n138 9.3005
R1013 VDD2.n94 VDD2.n93 9.3005
R1014 VDD2.n145 VDD2.n144 9.3005
R1015 VDD2.n147 VDD2.n146 9.3005
R1016 VDD2.n89 VDD2.n88 9.3005
R1017 VDD2.n153 VDD2.n152 9.3005
R1018 VDD2.n155 VDD2.n154 9.3005
R1019 VDD2.n162 VDD2.n161 9.3005
R1020 VDD2.n85 VDD2.n84 9.3005
R1021 VDD2.n98 VDD2.n97 9.3005
R1022 VDD2.n131 VDD2.n130 9.3005
R1023 VDD2.n129 VDD2.n128 9.3005
R1024 VDD2.n102 VDD2.n101 9.3005
R1025 VDD2.n123 VDD2.n122 9.3005
R1026 VDD2.n121 VDD2.n120 9.3005
R1027 VDD2.n106 VDD2.n105 9.3005
R1028 VDD2.n115 VDD2.n114 9.3005
R1029 VDD2.n113 VDD2.n112 9.3005
R1030 VDD2.n79 VDD2.n78 9.3005
R1031 VDD2.n2 VDD2.n1 9.3005
R1032 VDD2.n47 VDD2.n46 9.3005
R1033 VDD2.n45 VDD2.n44 9.3005
R1034 VDD2.n18 VDD2.n17 9.3005
R1035 VDD2.n39 VDD2.n38 9.3005
R1036 VDD2.n37 VDD2.n36 9.3005
R1037 VDD2.n22 VDD2.n21 9.3005
R1038 VDD2.n31 VDD2.n30 9.3005
R1039 VDD2.n29 VDD2.n28 9.3005
R1040 VDD2.n14 VDD2.n13 9.3005
R1041 VDD2.n53 VDD2.n52 9.3005
R1042 VDD2.n55 VDD2.n54 9.3005
R1043 VDD2.n10 VDD2.n9 9.3005
R1044 VDD2.n61 VDD2.n60 9.3005
R1045 VDD2.n63 VDD2.n62 9.3005
R1046 VDD2.n6 VDD2.n5 9.3005
R1047 VDD2.n70 VDD2.n69 9.3005
R1048 VDD2.n72 VDD2.n71 9.3005
R1049 VDD2.n140 VDD2.n94 8.92171
R1050 VDD2.n127 VDD2.n102 8.92171
R1051 VDD2.n43 VDD2.n18 8.92171
R1052 VDD2.n56 VDD2.n10 8.92171
R1053 VDD2.n139 VDD2.n96 8.14595
R1054 VDD2.n128 VDD2.n100 8.14595
R1055 VDD2.n44 VDD2.n16 8.14595
R1056 VDD2.n55 VDD2.n12 8.14595
R1057 VDD2.n136 VDD2.n135 7.3702
R1058 VDD2.n132 VDD2.n131 7.3702
R1059 VDD2.n48 VDD2.n47 7.3702
R1060 VDD2.n52 VDD2.n51 7.3702
R1061 VDD2.n135 VDD2.n98 6.59444
R1062 VDD2.n132 VDD2.n98 6.59444
R1063 VDD2.n48 VDD2.n14 6.59444
R1064 VDD2.n51 VDD2.n14 6.59444
R1065 VDD2.n136 VDD2.n96 5.81868
R1066 VDD2.n131 VDD2.n100 5.81868
R1067 VDD2.n47 VDD2.n16 5.81868
R1068 VDD2.n52 VDD2.n12 5.81868
R1069 VDD2.n140 VDD2.n139 5.04292
R1070 VDD2.n128 VDD2.n127 5.04292
R1071 VDD2.n44 VDD2.n43 5.04292
R1072 VDD2.n56 VDD2.n55 5.04292
R1073 VDD2.n143 VDD2.n94 4.26717
R1074 VDD2.n124 VDD2.n102 4.26717
R1075 VDD2.n40 VDD2.n18 4.26717
R1076 VDD2.n59 VDD2.n10 4.26717
R1077 VDD2.n113 VDD2.n109 3.70982
R1078 VDD2.n29 VDD2.n25 3.70982
R1079 VDD2.n144 VDD2.n92 3.49141
R1080 VDD2.n123 VDD2.n104 3.49141
R1081 VDD2.n39 VDD2.n20 3.49141
R1082 VDD2.n60 VDD2.n8 3.49141
R1083 VDD2.n148 VDD2.n147 2.71565
R1084 VDD2.n120 VDD2.n119 2.71565
R1085 VDD2.n36 VDD2.n35 2.71565
R1086 VDD2.n64 VDD2.n63 2.71565
R1087 VDD2 VDD2.n164 2.24403
R1088 VDD2.n165 VDD2.t5 2.19382
R1089 VDD2.n165 VDD2.t3 2.19382
R1090 VDD2.n81 VDD2.t1 2.19382
R1091 VDD2.n81 VDD2.t2 2.19382
R1092 VDD2.n163 VDD2.n83 1.93989
R1093 VDD2.n151 VDD2.n89 1.93989
R1094 VDD2.n116 VDD2.n106 1.93989
R1095 VDD2.n32 VDD2.n22 1.93989
R1096 VDD2.n68 VDD2.n6 1.93989
R1097 VDD2.n80 VDD2.n0 1.93989
R1098 VDD2.n161 VDD2.n160 1.16414
R1099 VDD2.n152 VDD2.n87 1.16414
R1100 VDD2.n115 VDD2.n108 1.16414
R1101 VDD2.n31 VDD2.n24 1.16414
R1102 VDD2.n69 VDD2.n4 1.16414
R1103 VDD2.n78 VDD2.n77 1.16414
R1104 VDD2.n157 VDD2.n85 0.388379
R1105 VDD2.n156 VDD2.n155 0.388379
R1106 VDD2.n112 VDD2.n111 0.388379
R1107 VDD2.n28 VDD2.n27 0.388379
R1108 VDD2.n73 VDD2.n72 0.388379
R1109 VDD2.n74 VDD2.n2 0.388379
R1110 VDD2.n162 VDD2.n84 0.155672
R1111 VDD2.n154 VDD2.n84 0.155672
R1112 VDD2.n154 VDD2.n153 0.155672
R1113 VDD2.n153 VDD2.n88 0.155672
R1114 VDD2.n146 VDD2.n88 0.155672
R1115 VDD2.n146 VDD2.n145 0.155672
R1116 VDD2.n145 VDD2.n93 0.155672
R1117 VDD2.n138 VDD2.n93 0.155672
R1118 VDD2.n138 VDD2.n137 0.155672
R1119 VDD2.n137 VDD2.n97 0.155672
R1120 VDD2.n130 VDD2.n97 0.155672
R1121 VDD2.n130 VDD2.n129 0.155672
R1122 VDD2.n129 VDD2.n101 0.155672
R1123 VDD2.n122 VDD2.n101 0.155672
R1124 VDD2.n122 VDD2.n121 0.155672
R1125 VDD2.n121 VDD2.n105 0.155672
R1126 VDD2.n114 VDD2.n105 0.155672
R1127 VDD2.n114 VDD2.n113 0.155672
R1128 VDD2.n30 VDD2.n29 0.155672
R1129 VDD2.n30 VDD2.n21 0.155672
R1130 VDD2.n37 VDD2.n21 0.155672
R1131 VDD2.n38 VDD2.n37 0.155672
R1132 VDD2.n38 VDD2.n17 0.155672
R1133 VDD2.n45 VDD2.n17 0.155672
R1134 VDD2.n46 VDD2.n45 0.155672
R1135 VDD2.n46 VDD2.n13 0.155672
R1136 VDD2.n53 VDD2.n13 0.155672
R1137 VDD2.n54 VDD2.n53 0.155672
R1138 VDD2.n54 VDD2.n9 0.155672
R1139 VDD2.n61 VDD2.n9 0.155672
R1140 VDD2.n62 VDD2.n61 0.155672
R1141 VDD2.n62 VDD2.n5 0.155672
R1142 VDD2.n70 VDD2.n5 0.155672
R1143 VDD2.n71 VDD2.n70 0.155672
R1144 VDD2.n71 VDD2.n1 0.155672
R1145 VDD2.n79 VDD2.n1 0.155672
R1146 B.n597 B.n84 585
R1147 B.n599 B.n598 585
R1148 B.n600 B.n83 585
R1149 B.n602 B.n601 585
R1150 B.n603 B.n82 585
R1151 B.n605 B.n604 585
R1152 B.n606 B.n81 585
R1153 B.n608 B.n607 585
R1154 B.n609 B.n80 585
R1155 B.n611 B.n610 585
R1156 B.n612 B.n79 585
R1157 B.n614 B.n613 585
R1158 B.n615 B.n78 585
R1159 B.n617 B.n616 585
R1160 B.n618 B.n77 585
R1161 B.n620 B.n619 585
R1162 B.n621 B.n76 585
R1163 B.n623 B.n622 585
R1164 B.n624 B.n75 585
R1165 B.n626 B.n625 585
R1166 B.n627 B.n74 585
R1167 B.n629 B.n628 585
R1168 B.n630 B.n73 585
R1169 B.n632 B.n631 585
R1170 B.n633 B.n72 585
R1171 B.n635 B.n634 585
R1172 B.n636 B.n71 585
R1173 B.n638 B.n637 585
R1174 B.n639 B.n70 585
R1175 B.n641 B.n640 585
R1176 B.n642 B.n69 585
R1177 B.n644 B.n643 585
R1178 B.n645 B.n68 585
R1179 B.n647 B.n646 585
R1180 B.n648 B.n67 585
R1181 B.n650 B.n649 585
R1182 B.n651 B.n66 585
R1183 B.n653 B.n652 585
R1184 B.n654 B.n65 585
R1185 B.n656 B.n655 585
R1186 B.n657 B.n64 585
R1187 B.n659 B.n658 585
R1188 B.n660 B.n63 585
R1189 B.n662 B.n661 585
R1190 B.n663 B.n62 585
R1191 B.n665 B.n664 585
R1192 B.n666 B.n61 585
R1193 B.n668 B.n667 585
R1194 B.n669 B.n60 585
R1195 B.n671 B.n670 585
R1196 B.n673 B.n57 585
R1197 B.n675 B.n674 585
R1198 B.n676 B.n56 585
R1199 B.n678 B.n677 585
R1200 B.n679 B.n55 585
R1201 B.n681 B.n680 585
R1202 B.n682 B.n54 585
R1203 B.n684 B.n683 585
R1204 B.n685 B.n51 585
R1205 B.n688 B.n687 585
R1206 B.n689 B.n50 585
R1207 B.n691 B.n690 585
R1208 B.n692 B.n49 585
R1209 B.n694 B.n693 585
R1210 B.n695 B.n48 585
R1211 B.n697 B.n696 585
R1212 B.n698 B.n47 585
R1213 B.n700 B.n699 585
R1214 B.n701 B.n46 585
R1215 B.n703 B.n702 585
R1216 B.n704 B.n45 585
R1217 B.n706 B.n705 585
R1218 B.n707 B.n44 585
R1219 B.n709 B.n708 585
R1220 B.n710 B.n43 585
R1221 B.n712 B.n711 585
R1222 B.n713 B.n42 585
R1223 B.n715 B.n714 585
R1224 B.n716 B.n41 585
R1225 B.n718 B.n717 585
R1226 B.n719 B.n40 585
R1227 B.n721 B.n720 585
R1228 B.n722 B.n39 585
R1229 B.n724 B.n723 585
R1230 B.n725 B.n38 585
R1231 B.n727 B.n726 585
R1232 B.n728 B.n37 585
R1233 B.n730 B.n729 585
R1234 B.n731 B.n36 585
R1235 B.n733 B.n732 585
R1236 B.n734 B.n35 585
R1237 B.n736 B.n735 585
R1238 B.n737 B.n34 585
R1239 B.n739 B.n738 585
R1240 B.n740 B.n33 585
R1241 B.n742 B.n741 585
R1242 B.n743 B.n32 585
R1243 B.n745 B.n744 585
R1244 B.n746 B.n31 585
R1245 B.n748 B.n747 585
R1246 B.n749 B.n30 585
R1247 B.n751 B.n750 585
R1248 B.n752 B.n29 585
R1249 B.n754 B.n753 585
R1250 B.n755 B.n28 585
R1251 B.n757 B.n756 585
R1252 B.n758 B.n27 585
R1253 B.n760 B.n759 585
R1254 B.n761 B.n26 585
R1255 B.n596 B.n595 585
R1256 B.n594 B.n85 585
R1257 B.n593 B.n592 585
R1258 B.n591 B.n86 585
R1259 B.n590 B.n589 585
R1260 B.n588 B.n87 585
R1261 B.n587 B.n586 585
R1262 B.n585 B.n88 585
R1263 B.n584 B.n583 585
R1264 B.n582 B.n89 585
R1265 B.n581 B.n580 585
R1266 B.n579 B.n90 585
R1267 B.n578 B.n577 585
R1268 B.n576 B.n91 585
R1269 B.n575 B.n574 585
R1270 B.n573 B.n92 585
R1271 B.n572 B.n571 585
R1272 B.n570 B.n93 585
R1273 B.n569 B.n568 585
R1274 B.n567 B.n94 585
R1275 B.n566 B.n565 585
R1276 B.n564 B.n95 585
R1277 B.n563 B.n562 585
R1278 B.n561 B.n96 585
R1279 B.n560 B.n559 585
R1280 B.n558 B.n97 585
R1281 B.n557 B.n556 585
R1282 B.n555 B.n98 585
R1283 B.n554 B.n553 585
R1284 B.n552 B.n99 585
R1285 B.n551 B.n550 585
R1286 B.n549 B.n100 585
R1287 B.n548 B.n547 585
R1288 B.n546 B.n101 585
R1289 B.n545 B.n544 585
R1290 B.n543 B.n102 585
R1291 B.n542 B.n541 585
R1292 B.n540 B.n103 585
R1293 B.n539 B.n538 585
R1294 B.n537 B.n104 585
R1295 B.n536 B.n535 585
R1296 B.n534 B.n105 585
R1297 B.n533 B.n532 585
R1298 B.n531 B.n106 585
R1299 B.n530 B.n529 585
R1300 B.n528 B.n107 585
R1301 B.n527 B.n526 585
R1302 B.n525 B.n108 585
R1303 B.n524 B.n523 585
R1304 B.n522 B.n109 585
R1305 B.n521 B.n520 585
R1306 B.n519 B.n110 585
R1307 B.n518 B.n517 585
R1308 B.n516 B.n111 585
R1309 B.n515 B.n514 585
R1310 B.n513 B.n112 585
R1311 B.n512 B.n511 585
R1312 B.n510 B.n113 585
R1313 B.n509 B.n508 585
R1314 B.n507 B.n114 585
R1315 B.n506 B.n505 585
R1316 B.n504 B.n115 585
R1317 B.n503 B.n502 585
R1318 B.n501 B.n116 585
R1319 B.n500 B.n499 585
R1320 B.n498 B.n117 585
R1321 B.n497 B.n496 585
R1322 B.n495 B.n118 585
R1323 B.n494 B.n493 585
R1324 B.n492 B.n119 585
R1325 B.n491 B.n490 585
R1326 B.n489 B.n120 585
R1327 B.n488 B.n487 585
R1328 B.n486 B.n121 585
R1329 B.n485 B.n484 585
R1330 B.n483 B.n122 585
R1331 B.n482 B.n481 585
R1332 B.n480 B.n123 585
R1333 B.n479 B.n478 585
R1334 B.n477 B.n124 585
R1335 B.n476 B.n475 585
R1336 B.n474 B.n125 585
R1337 B.n473 B.n472 585
R1338 B.n471 B.n126 585
R1339 B.n470 B.n469 585
R1340 B.n468 B.n127 585
R1341 B.n467 B.n466 585
R1342 B.n465 B.n128 585
R1343 B.n464 B.n463 585
R1344 B.n462 B.n129 585
R1345 B.n461 B.n460 585
R1346 B.n459 B.n130 585
R1347 B.n458 B.n457 585
R1348 B.n456 B.n131 585
R1349 B.n455 B.n454 585
R1350 B.n453 B.n132 585
R1351 B.n452 B.n451 585
R1352 B.n287 B.n286 585
R1353 B.n288 B.n191 585
R1354 B.n290 B.n289 585
R1355 B.n291 B.n190 585
R1356 B.n293 B.n292 585
R1357 B.n294 B.n189 585
R1358 B.n296 B.n295 585
R1359 B.n297 B.n188 585
R1360 B.n299 B.n298 585
R1361 B.n300 B.n187 585
R1362 B.n302 B.n301 585
R1363 B.n303 B.n186 585
R1364 B.n305 B.n304 585
R1365 B.n306 B.n185 585
R1366 B.n308 B.n307 585
R1367 B.n309 B.n184 585
R1368 B.n311 B.n310 585
R1369 B.n312 B.n183 585
R1370 B.n314 B.n313 585
R1371 B.n315 B.n182 585
R1372 B.n317 B.n316 585
R1373 B.n318 B.n181 585
R1374 B.n320 B.n319 585
R1375 B.n321 B.n180 585
R1376 B.n323 B.n322 585
R1377 B.n324 B.n179 585
R1378 B.n326 B.n325 585
R1379 B.n327 B.n178 585
R1380 B.n329 B.n328 585
R1381 B.n330 B.n177 585
R1382 B.n332 B.n331 585
R1383 B.n333 B.n176 585
R1384 B.n335 B.n334 585
R1385 B.n336 B.n175 585
R1386 B.n338 B.n337 585
R1387 B.n339 B.n174 585
R1388 B.n341 B.n340 585
R1389 B.n342 B.n173 585
R1390 B.n344 B.n343 585
R1391 B.n345 B.n172 585
R1392 B.n347 B.n346 585
R1393 B.n348 B.n171 585
R1394 B.n350 B.n349 585
R1395 B.n351 B.n170 585
R1396 B.n353 B.n352 585
R1397 B.n354 B.n169 585
R1398 B.n356 B.n355 585
R1399 B.n357 B.n168 585
R1400 B.n359 B.n358 585
R1401 B.n360 B.n165 585
R1402 B.n363 B.n362 585
R1403 B.n364 B.n164 585
R1404 B.n366 B.n365 585
R1405 B.n367 B.n163 585
R1406 B.n369 B.n368 585
R1407 B.n370 B.n162 585
R1408 B.n372 B.n371 585
R1409 B.n373 B.n161 585
R1410 B.n375 B.n374 585
R1411 B.n377 B.n376 585
R1412 B.n378 B.n157 585
R1413 B.n380 B.n379 585
R1414 B.n381 B.n156 585
R1415 B.n383 B.n382 585
R1416 B.n384 B.n155 585
R1417 B.n386 B.n385 585
R1418 B.n387 B.n154 585
R1419 B.n389 B.n388 585
R1420 B.n390 B.n153 585
R1421 B.n392 B.n391 585
R1422 B.n393 B.n152 585
R1423 B.n395 B.n394 585
R1424 B.n396 B.n151 585
R1425 B.n398 B.n397 585
R1426 B.n399 B.n150 585
R1427 B.n401 B.n400 585
R1428 B.n402 B.n149 585
R1429 B.n404 B.n403 585
R1430 B.n405 B.n148 585
R1431 B.n407 B.n406 585
R1432 B.n408 B.n147 585
R1433 B.n410 B.n409 585
R1434 B.n411 B.n146 585
R1435 B.n413 B.n412 585
R1436 B.n414 B.n145 585
R1437 B.n416 B.n415 585
R1438 B.n417 B.n144 585
R1439 B.n419 B.n418 585
R1440 B.n420 B.n143 585
R1441 B.n422 B.n421 585
R1442 B.n423 B.n142 585
R1443 B.n425 B.n424 585
R1444 B.n426 B.n141 585
R1445 B.n428 B.n427 585
R1446 B.n429 B.n140 585
R1447 B.n431 B.n430 585
R1448 B.n432 B.n139 585
R1449 B.n434 B.n433 585
R1450 B.n435 B.n138 585
R1451 B.n437 B.n436 585
R1452 B.n438 B.n137 585
R1453 B.n440 B.n439 585
R1454 B.n441 B.n136 585
R1455 B.n443 B.n442 585
R1456 B.n444 B.n135 585
R1457 B.n446 B.n445 585
R1458 B.n447 B.n134 585
R1459 B.n449 B.n448 585
R1460 B.n450 B.n133 585
R1461 B.n285 B.n192 585
R1462 B.n284 B.n283 585
R1463 B.n282 B.n193 585
R1464 B.n281 B.n280 585
R1465 B.n279 B.n194 585
R1466 B.n278 B.n277 585
R1467 B.n276 B.n195 585
R1468 B.n275 B.n274 585
R1469 B.n273 B.n196 585
R1470 B.n272 B.n271 585
R1471 B.n270 B.n197 585
R1472 B.n269 B.n268 585
R1473 B.n267 B.n198 585
R1474 B.n266 B.n265 585
R1475 B.n264 B.n199 585
R1476 B.n263 B.n262 585
R1477 B.n261 B.n200 585
R1478 B.n260 B.n259 585
R1479 B.n258 B.n201 585
R1480 B.n257 B.n256 585
R1481 B.n255 B.n202 585
R1482 B.n254 B.n253 585
R1483 B.n252 B.n203 585
R1484 B.n251 B.n250 585
R1485 B.n249 B.n204 585
R1486 B.n248 B.n247 585
R1487 B.n246 B.n205 585
R1488 B.n245 B.n244 585
R1489 B.n243 B.n206 585
R1490 B.n242 B.n241 585
R1491 B.n240 B.n207 585
R1492 B.n239 B.n238 585
R1493 B.n237 B.n208 585
R1494 B.n236 B.n235 585
R1495 B.n234 B.n209 585
R1496 B.n233 B.n232 585
R1497 B.n231 B.n210 585
R1498 B.n230 B.n229 585
R1499 B.n228 B.n211 585
R1500 B.n227 B.n226 585
R1501 B.n225 B.n212 585
R1502 B.n224 B.n223 585
R1503 B.n222 B.n213 585
R1504 B.n221 B.n220 585
R1505 B.n219 B.n214 585
R1506 B.n218 B.n217 585
R1507 B.n216 B.n215 585
R1508 B.n2 B.n0 585
R1509 B.n833 B.n1 585
R1510 B.n832 B.n831 585
R1511 B.n830 B.n3 585
R1512 B.n829 B.n828 585
R1513 B.n827 B.n4 585
R1514 B.n826 B.n825 585
R1515 B.n824 B.n5 585
R1516 B.n823 B.n822 585
R1517 B.n821 B.n6 585
R1518 B.n820 B.n819 585
R1519 B.n818 B.n7 585
R1520 B.n817 B.n816 585
R1521 B.n815 B.n8 585
R1522 B.n814 B.n813 585
R1523 B.n812 B.n9 585
R1524 B.n811 B.n810 585
R1525 B.n809 B.n10 585
R1526 B.n808 B.n807 585
R1527 B.n806 B.n11 585
R1528 B.n805 B.n804 585
R1529 B.n803 B.n12 585
R1530 B.n802 B.n801 585
R1531 B.n800 B.n13 585
R1532 B.n799 B.n798 585
R1533 B.n797 B.n14 585
R1534 B.n796 B.n795 585
R1535 B.n794 B.n15 585
R1536 B.n793 B.n792 585
R1537 B.n791 B.n16 585
R1538 B.n790 B.n789 585
R1539 B.n788 B.n17 585
R1540 B.n787 B.n786 585
R1541 B.n785 B.n18 585
R1542 B.n784 B.n783 585
R1543 B.n782 B.n19 585
R1544 B.n781 B.n780 585
R1545 B.n779 B.n20 585
R1546 B.n778 B.n777 585
R1547 B.n776 B.n21 585
R1548 B.n775 B.n774 585
R1549 B.n773 B.n22 585
R1550 B.n772 B.n771 585
R1551 B.n770 B.n23 585
R1552 B.n769 B.n768 585
R1553 B.n767 B.n24 585
R1554 B.n766 B.n765 585
R1555 B.n764 B.n25 585
R1556 B.n763 B.n762 585
R1557 B.n835 B.n834 585
R1558 B.n286 B.n285 511.721
R1559 B.n762 B.n761 511.721
R1560 B.n452 B.n133 511.721
R1561 B.n597 B.n596 511.721
R1562 B.n158 B.t5 492.012
R1563 B.n58 B.t10 492.012
R1564 B.n166 B.t2 492.012
R1565 B.n52 B.t7 492.012
R1566 B.n159 B.t4 426.459
R1567 B.n59 B.t11 426.459
R1568 B.n167 B.t1 426.459
R1569 B.n53 B.t8 426.459
R1570 B.n158 B.t3 325.74
R1571 B.n166 B.t0 325.74
R1572 B.n52 B.t6 325.74
R1573 B.n58 B.t9 325.74
R1574 B.n285 B.n284 163.367
R1575 B.n284 B.n193 163.367
R1576 B.n280 B.n193 163.367
R1577 B.n280 B.n279 163.367
R1578 B.n279 B.n278 163.367
R1579 B.n278 B.n195 163.367
R1580 B.n274 B.n195 163.367
R1581 B.n274 B.n273 163.367
R1582 B.n273 B.n272 163.367
R1583 B.n272 B.n197 163.367
R1584 B.n268 B.n197 163.367
R1585 B.n268 B.n267 163.367
R1586 B.n267 B.n266 163.367
R1587 B.n266 B.n199 163.367
R1588 B.n262 B.n199 163.367
R1589 B.n262 B.n261 163.367
R1590 B.n261 B.n260 163.367
R1591 B.n260 B.n201 163.367
R1592 B.n256 B.n201 163.367
R1593 B.n256 B.n255 163.367
R1594 B.n255 B.n254 163.367
R1595 B.n254 B.n203 163.367
R1596 B.n250 B.n203 163.367
R1597 B.n250 B.n249 163.367
R1598 B.n249 B.n248 163.367
R1599 B.n248 B.n205 163.367
R1600 B.n244 B.n205 163.367
R1601 B.n244 B.n243 163.367
R1602 B.n243 B.n242 163.367
R1603 B.n242 B.n207 163.367
R1604 B.n238 B.n207 163.367
R1605 B.n238 B.n237 163.367
R1606 B.n237 B.n236 163.367
R1607 B.n236 B.n209 163.367
R1608 B.n232 B.n209 163.367
R1609 B.n232 B.n231 163.367
R1610 B.n231 B.n230 163.367
R1611 B.n230 B.n211 163.367
R1612 B.n226 B.n211 163.367
R1613 B.n226 B.n225 163.367
R1614 B.n225 B.n224 163.367
R1615 B.n224 B.n213 163.367
R1616 B.n220 B.n213 163.367
R1617 B.n220 B.n219 163.367
R1618 B.n219 B.n218 163.367
R1619 B.n218 B.n215 163.367
R1620 B.n215 B.n2 163.367
R1621 B.n834 B.n2 163.367
R1622 B.n834 B.n833 163.367
R1623 B.n833 B.n832 163.367
R1624 B.n832 B.n3 163.367
R1625 B.n828 B.n3 163.367
R1626 B.n828 B.n827 163.367
R1627 B.n827 B.n826 163.367
R1628 B.n826 B.n5 163.367
R1629 B.n822 B.n5 163.367
R1630 B.n822 B.n821 163.367
R1631 B.n821 B.n820 163.367
R1632 B.n820 B.n7 163.367
R1633 B.n816 B.n7 163.367
R1634 B.n816 B.n815 163.367
R1635 B.n815 B.n814 163.367
R1636 B.n814 B.n9 163.367
R1637 B.n810 B.n9 163.367
R1638 B.n810 B.n809 163.367
R1639 B.n809 B.n808 163.367
R1640 B.n808 B.n11 163.367
R1641 B.n804 B.n11 163.367
R1642 B.n804 B.n803 163.367
R1643 B.n803 B.n802 163.367
R1644 B.n802 B.n13 163.367
R1645 B.n798 B.n13 163.367
R1646 B.n798 B.n797 163.367
R1647 B.n797 B.n796 163.367
R1648 B.n796 B.n15 163.367
R1649 B.n792 B.n15 163.367
R1650 B.n792 B.n791 163.367
R1651 B.n791 B.n790 163.367
R1652 B.n790 B.n17 163.367
R1653 B.n786 B.n17 163.367
R1654 B.n786 B.n785 163.367
R1655 B.n785 B.n784 163.367
R1656 B.n784 B.n19 163.367
R1657 B.n780 B.n19 163.367
R1658 B.n780 B.n779 163.367
R1659 B.n779 B.n778 163.367
R1660 B.n778 B.n21 163.367
R1661 B.n774 B.n21 163.367
R1662 B.n774 B.n773 163.367
R1663 B.n773 B.n772 163.367
R1664 B.n772 B.n23 163.367
R1665 B.n768 B.n23 163.367
R1666 B.n768 B.n767 163.367
R1667 B.n767 B.n766 163.367
R1668 B.n766 B.n25 163.367
R1669 B.n762 B.n25 163.367
R1670 B.n286 B.n191 163.367
R1671 B.n290 B.n191 163.367
R1672 B.n291 B.n290 163.367
R1673 B.n292 B.n291 163.367
R1674 B.n292 B.n189 163.367
R1675 B.n296 B.n189 163.367
R1676 B.n297 B.n296 163.367
R1677 B.n298 B.n297 163.367
R1678 B.n298 B.n187 163.367
R1679 B.n302 B.n187 163.367
R1680 B.n303 B.n302 163.367
R1681 B.n304 B.n303 163.367
R1682 B.n304 B.n185 163.367
R1683 B.n308 B.n185 163.367
R1684 B.n309 B.n308 163.367
R1685 B.n310 B.n309 163.367
R1686 B.n310 B.n183 163.367
R1687 B.n314 B.n183 163.367
R1688 B.n315 B.n314 163.367
R1689 B.n316 B.n315 163.367
R1690 B.n316 B.n181 163.367
R1691 B.n320 B.n181 163.367
R1692 B.n321 B.n320 163.367
R1693 B.n322 B.n321 163.367
R1694 B.n322 B.n179 163.367
R1695 B.n326 B.n179 163.367
R1696 B.n327 B.n326 163.367
R1697 B.n328 B.n327 163.367
R1698 B.n328 B.n177 163.367
R1699 B.n332 B.n177 163.367
R1700 B.n333 B.n332 163.367
R1701 B.n334 B.n333 163.367
R1702 B.n334 B.n175 163.367
R1703 B.n338 B.n175 163.367
R1704 B.n339 B.n338 163.367
R1705 B.n340 B.n339 163.367
R1706 B.n340 B.n173 163.367
R1707 B.n344 B.n173 163.367
R1708 B.n345 B.n344 163.367
R1709 B.n346 B.n345 163.367
R1710 B.n346 B.n171 163.367
R1711 B.n350 B.n171 163.367
R1712 B.n351 B.n350 163.367
R1713 B.n352 B.n351 163.367
R1714 B.n352 B.n169 163.367
R1715 B.n356 B.n169 163.367
R1716 B.n357 B.n356 163.367
R1717 B.n358 B.n357 163.367
R1718 B.n358 B.n165 163.367
R1719 B.n363 B.n165 163.367
R1720 B.n364 B.n363 163.367
R1721 B.n365 B.n364 163.367
R1722 B.n365 B.n163 163.367
R1723 B.n369 B.n163 163.367
R1724 B.n370 B.n369 163.367
R1725 B.n371 B.n370 163.367
R1726 B.n371 B.n161 163.367
R1727 B.n375 B.n161 163.367
R1728 B.n376 B.n375 163.367
R1729 B.n376 B.n157 163.367
R1730 B.n380 B.n157 163.367
R1731 B.n381 B.n380 163.367
R1732 B.n382 B.n381 163.367
R1733 B.n382 B.n155 163.367
R1734 B.n386 B.n155 163.367
R1735 B.n387 B.n386 163.367
R1736 B.n388 B.n387 163.367
R1737 B.n388 B.n153 163.367
R1738 B.n392 B.n153 163.367
R1739 B.n393 B.n392 163.367
R1740 B.n394 B.n393 163.367
R1741 B.n394 B.n151 163.367
R1742 B.n398 B.n151 163.367
R1743 B.n399 B.n398 163.367
R1744 B.n400 B.n399 163.367
R1745 B.n400 B.n149 163.367
R1746 B.n404 B.n149 163.367
R1747 B.n405 B.n404 163.367
R1748 B.n406 B.n405 163.367
R1749 B.n406 B.n147 163.367
R1750 B.n410 B.n147 163.367
R1751 B.n411 B.n410 163.367
R1752 B.n412 B.n411 163.367
R1753 B.n412 B.n145 163.367
R1754 B.n416 B.n145 163.367
R1755 B.n417 B.n416 163.367
R1756 B.n418 B.n417 163.367
R1757 B.n418 B.n143 163.367
R1758 B.n422 B.n143 163.367
R1759 B.n423 B.n422 163.367
R1760 B.n424 B.n423 163.367
R1761 B.n424 B.n141 163.367
R1762 B.n428 B.n141 163.367
R1763 B.n429 B.n428 163.367
R1764 B.n430 B.n429 163.367
R1765 B.n430 B.n139 163.367
R1766 B.n434 B.n139 163.367
R1767 B.n435 B.n434 163.367
R1768 B.n436 B.n435 163.367
R1769 B.n436 B.n137 163.367
R1770 B.n440 B.n137 163.367
R1771 B.n441 B.n440 163.367
R1772 B.n442 B.n441 163.367
R1773 B.n442 B.n135 163.367
R1774 B.n446 B.n135 163.367
R1775 B.n447 B.n446 163.367
R1776 B.n448 B.n447 163.367
R1777 B.n448 B.n133 163.367
R1778 B.n453 B.n452 163.367
R1779 B.n454 B.n453 163.367
R1780 B.n454 B.n131 163.367
R1781 B.n458 B.n131 163.367
R1782 B.n459 B.n458 163.367
R1783 B.n460 B.n459 163.367
R1784 B.n460 B.n129 163.367
R1785 B.n464 B.n129 163.367
R1786 B.n465 B.n464 163.367
R1787 B.n466 B.n465 163.367
R1788 B.n466 B.n127 163.367
R1789 B.n470 B.n127 163.367
R1790 B.n471 B.n470 163.367
R1791 B.n472 B.n471 163.367
R1792 B.n472 B.n125 163.367
R1793 B.n476 B.n125 163.367
R1794 B.n477 B.n476 163.367
R1795 B.n478 B.n477 163.367
R1796 B.n478 B.n123 163.367
R1797 B.n482 B.n123 163.367
R1798 B.n483 B.n482 163.367
R1799 B.n484 B.n483 163.367
R1800 B.n484 B.n121 163.367
R1801 B.n488 B.n121 163.367
R1802 B.n489 B.n488 163.367
R1803 B.n490 B.n489 163.367
R1804 B.n490 B.n119 163.367
R1805 B.n494 B.n119 163.367
R1806 B.n495 B.n494 163.367
R1807 B.n496 B.n495 163.367
R1808 B.n496 B.n117 163.367
R1809 B.n500 B.n117 163.367
R1810 B.n501 B.n500 163.367
R1811 B.n502 B.n501 163.367
R1812 B.n502 B.n115 163.367
R1813 B.n506 B.n115 163.367
R1814 B.n507 B.n506 163.367
R1815 B.n508 B.n507 163.367
R1816 B.n508 B.n113 163.367
R1817 B.n512 B.n113 163.367
R1818 B.n513 B.n512 163.367
R1819 B.n514 B.n513 163.367
R1820 B.n514 B.n111 163.367
R1821 B.n518 B.n111 163.367
R1822 B.n519 B.n518 163.367
R1823 B.n520 B.n519 163.367
R1824 B.n520 B.n109 163.367
R1825 B.n524 B.n109 163.367
R1826 B.n525 B.n524 163.367
R1827 B.n526 B.n525 163.367
R1828 B.n526 B.n107 163.367
R1829 B.n530 B.n107 163.367
R1830 B.n531 B.n530 163.367
R1831 B.n532 B.n531 163.367
R1832 B.n532 B.n105 163.367
R1833 B.n536 B.n105 163.367
R1834 B.n537 B.n536 163.367
R1835 B.n538 B.n537 163.367
R1836 B.n538 B.n103 163.367
R1837 B.n542 B.n103 163.367
R1838 B.n543 B.n542 163.367
R1839 B.n544 B.n543 163.367
R1840 B.n544 B.n101 163.367
R1841 B.n548 B.n101 163.367
R1842 B.n549 B.n548 163.367
R1843 B.n550 B.n549 163.367
R1844 B.n550 B.n99 163.367
R1845 B.n554 B.n99 163.367
R1846 B.n555 B.n554 163.367
R1847 B.n556 B.n555 163.367
R1848 B.n556 B.n97 163.367
R1849 B.n560 B.n97 163.367
R1850 B.n561 B.n560 163.367
R1851 B.n562 B.n561 163.367
R1852 B.n562 B.n95 163.367
R1853 B.n566 B.n95 163.367
R1854 B.n567 B.n566 163.367
R1855 B.n568 B.n567 163.367
R1856 B.n568 B.n93 163.367
R1857 B.n572 B.n93 163.367
R1858 B.n573 B.n572 163.367
R1859 B.n574 B.n573 163.367
R1860 B.n574 B.n91 163.367
R1861 B.n578 B.n91 163.367
R1862 B.n579 B.n578 163.367
R1863 B.n580 B.n579 163.367
R1864 B.n580 B.n89 163.367
R1865 B.n584 B.n89 163.367
R1866 B.n585 B.n584 163.367
R1867 B.n586 B.n585 163.367
R1868 B.n586 B.n87 163.367
R1869 B.n590 B.n87 163.367
R1870 B.n591 B.n590 163.367
R1871 B.n592 B.n591 163.367
R1872 B.n592 B.n85 163.367
R1873 B.n596 B.n85 163.367
R1874 B.n761 B.n760 163.367
R1875 B.n760 B.n27 163.367
R1876 B.n756 B.n27 163.367
R1877 B.n756 B.n755 163.367
R1878 B.n755 B.n754 163.367
R1879 B.n754 B.n29 163.367
R1880 B.n750 B.n29 163.367
R1881 B.n750 B.n749 163.367
R1882 B.n749 B.n748 163.367
R1883 B.n748 B.n31 163.367
R1884 B.n744 B.n31 163.367
R1885 B.n744 B.n743 163.367
R1886 B.n743 B.n742 163.367
R1887 B.n742 B.n33 163.367
R1888 B.n738 B.n33 163.367
R1889 B.n738 B.n737 163.367
R1890 B.n737 B.n736 163.367
R1891 B.n736 B.n35 163.367
R1892 B.n732 B.n35 163.367
R1893 B.n732 B.n731 163.367
R1894 B.n731 B.n730 163.367
R1895 B.n730 B.n37 163.367
R1896 B.n726 B.n37 163.367
R1897 B.n726 B.n725 163.367
R1898 B.n725 B.n724 163.367
R1899 B.n724 B.n39 163.367
R1900 B.n720 B.n39 163.367
R1901 B.n720 B.n719 163.367
R1902 B.n719 B.n718 163.367
R1903 B.n718 B.n41 163.367
R1904 B.n714 B.n41 163.367
R1905 B.n714 B.n713 163.367
R1906 B.n713 B.n712 163.367
R1907 B.n712 B.n43 163.367
R1908 B.n708 B.n43 163.367
R1909 B.n708 B.n707 163.367
R1910 B.n707 B.n706 163.367
R1911 B.n706 B.n45 163.367
R1912 B.n702 B.n45 163.367
R1913 B.n702 B.n701 163.367
R1914 B.n701 B.n700 163.367
R1915 B.n700 B.n47 163.367
R1916 B.n696 B.n47 163.367
R1917 B.n696 B.n695 163.367
R1918 B.n695 B.n694 163.367
R1919 B.n694 B.n49 163.367
R1920 B.n690 B.n49 163.367
R1921 B.n690 B.n689 163.367
R1922 B.n689 B.n688 163.367
R1923 B.n688 B.n51 163.367
R1924 B.n683 B.n51 163.367
R1925 B.n683 B.n682 163.367
R1926 B.n682 B.n681 163.367
R1927 B.n681 B.n55 163.367
R1928 B.n677 B.n55 163.367
R1929 B.n677 B.n676 163.367
R1930 B.n676 B.n675 163.367
R1931 B.n675 B.n57 163.367
R1932 B.n670 B.n57 163.367
R1933 B.n670 B.n669 163.367
R1934 B.n669 B.n668 163.367
R1935 B.n668 B.n61 163.367
R1936 B.n664 B.n61 163.367
R1937 B.n664 B.n663 163.367
R1938 B.n663 B.n662 163.367
R1939 B.n662 B.n63 163.367
R1940 B.n658 B.n63 163.367
R1941 B.n658 B.n657 163.367
R1942 B.n657 B.n656 163.367
R1943 B.n656 B.n65 163.367
R1944 B.n652 B.n65 163.367
R1945 B.n652 B.n651 163.367
R1946 B.n651 B.n650 163.367
R1947 B.n650 B.n67 163.367
R1948 B.n646 B.n67 163.367
R1949 B.n646 B.n645 163.367
R1950 B.n645 B.n644 163.367
R1951 B.n644 B.n69 163.367
R1952 B.n640 B.n69 163.367
R1953 B.n640 B.n639 163.367
R1954 B.n639 B.n638 163.367
R1955 B.n638 B.n71 163.367
R1956 B.n634 B.n71 163.367
R1957 B.n634 B.n633 163.367
R1958 B.n633 B.n632 163.367
R1959 B.n632 B.n73 163.367
R1960 B.n628 B.n73 163.367
R1961 B.n628 B.n627 163.367
R1962 B.n627 B.n626 163.367
R1963 B.n626 B.n75 163.367
R1964 B.n622 B.n75 163.367
R1965 B.n622 B.n621 163.367
R1966 B.n621 B.n620 163.367
R1967 B.n620 B.n77 163.367
R1968 B.n616 B.n77 163.367
R1969 B.n616 B.n615 163.367
R1970 B.n615 B.n614 163.367
R1971 B.n614 B.n79 163.367
R1972 B.n610 B.n79 163.367
R1973 B.n610 B.n609 163.367
R1974 B.n609 B.n608 163.367
R1975 B.n608 B.n81 163.367
R1976 B.n604 B.n81 163.367
R1977 B.n604 B.n603 163.367
R1978 B.n603 B.n602 163.367
R1979 B.n602 B.n83 163.367
R1980 B.n598 B.n83 163.367
R1981 B.n598 B.n597 163.367
R1982 B.n159 B.n158 65.552
R1983 B.n167 B.n166 65.552
R1984 B.n53 B.n52 65.552
R1985 B.n59 B.n58 65.552
R1986 B.n160 B.n159 59.5399
R1987 B.n361 B.n167 59.5399
R1988 B.n686 B.n53 59.5399
R1989 B.n672 B.n59 59.5399
R1990 B.n763 B.n26 33.2493
R1991 B.n595 B.n84 33.2493
R1992 B.n451 B.n450 33.2493
R1993 B.n287 B.n192 33.2493
R1994 B B.n835 18.0485
R1995 B.n759 B.n26 10.6151
R1996 B.n759 B.n758 10.6151
R1997 B.n758 B.n757 10.6151
R1998 B.n757 B.n28 10.6151
R1999 B.n753 B.n28 10.6151
R2000 B.n753 B.n752 10.6151
R2001 B.n752 B.n751 10.6151
R2002 B.n751 B.n30 10.6151
R2003 B.n747 B.n30 10.6151
R2004 B.n747 B.n746 10.6151
R2005 B.n746 B.n745 10.6151
R2006 B.n745 B.n32 10.6151
R2007 B.n741 B.n32 10.6151
R2008 B.n741 B.n740 10.6151
R2009 B.n740 B.n739 10.6151
R2010 B.n739 B.n34 10.6151
R2011 B.n735 B.n34 10.6151
R2012 B.n735 B.n734 10.6151
R2013 B.n734 B.n733 10.6151
R2014 B.n733 B.n36 10.6151
R2015 B.n729 B.n36 10.6151
R2016 B.n729 B.n728 10.6151
R2017 B.n728 B.n727 10.6151
R2018 B.n727 B.n38 10.6151
R2019 B.n723 B.n38 10.6151
R2020 B.n723 B.n722 10.6151
R2021 B.n722 B.n721 10.6151
R2022 B.n721 B.n40 10.6151
R2023 B.n717 B.n40 10.6151
R2024 B.n717 B.n716 10.6151
R2025 B.n716 B.n715 10.6151
R2026 B.n715 B.n42 10.6151
R2027 B.n711 B.n42 10.6151
R2028 B.n711 B.n710 10.6151
R2029 B.n710 B.n709 10.6151
R2030 B.n709 B.n44 10.6151
R2031 B.n705 B.n44 10.6151
R2032 B.n705 B.n704 10.6151
R2033 B.n704 B.n703 10.6151
R2034 B.n703 B.n46 10.6151
R2035 B.n699 B.n46 10.6151
R2036 B.n699 B.n698 10.6151
R2037 B.n698 B.n697 10.6151
R2038 B.n697 B.n48 10.6151
R2039 B.n693 B.n48 10.6151
R2040 B.n693 B.n692 10.6151
R2041 B.n692 B.n691 10.6151
R2042 B.n691 B.n50 10.6151
R2043 B.n687 B.n50 10.6151
R2044 B.n685 B.n684 10.6151
R2045 B.n684 B.n54 10.6151
R2046 B.n680 B.n54 10.6151
R2047 B.n680 B.n679 10.6151
R2048 B.n679 B.n678 10.6151
R2049 B.n678 B.n56 10.6151
R2050 B.n674 B.n56 10.6151
R2051 B.n674 B.n673 10.6151
R2052 B.n671 B.n60 10.6151
R2053 B.n667 B.n60 10.6151
R2054 B.n667 B.n666 10.6151
R2055 B.n666 B.n665 10.6151
R2056 B.n665 B.n62 10.6151
R2057 B.n661 B.n62 10.6151
R2058 B.n661 B.n660 10.6151
R2059 B.n660 B.n659 10.6151
R2060 B.n659 B.n64 10.6151
R2061 B.n655 B.n64 10.6151
R2062 B.n655 B.n654 10.6151
R2063 B.n654 B.n653 10.6151
R2064 B.n653 B.n66 10.6151
R2065 B.n649 B.n66 10.6151
R2066 B.n649 B.n648 10.6151
R2067 B.n648 B.n647 10.6151
R2068 B.n647 B.n68 10.6151
R2069 B.n643 B.n68 10.6151
R2070 B.n643 B.n642 10.6151
R2071 B.n642 B.n641 10.6151
R2072 B.n641 B.n70 10.6151
R2073 B.n637 B.n70 10.6151
R2074 B.n637 B.n636 10.6151
R2075 B.n636 B.n635 10.6151
R2076 B.n635 B.n72 10.6151
R2077 B.n631 B.n72 10.6151
R2078 B.n631 B.n630 10.6151
R2079 B.n630 B.n629 10.6151
R2080 B.n629 B.n74 10.6151
R2081 B.n625 B.n74 10.6151
R2082 B.n625 B.n624 10.6151
R2083 B.n624 B.n623 10.6151
R2084 B.n623 B.n76 10.6151
R2085 B.n619 B.n76 10.6151
R2086 B.n619 B.n618 10.6151
R2087 B.n618 B.n617 10.6151
R2088 B.n617 B.n78 10.6151
R2089 B.n613 B.n78 10.6151
R2090 B.n613 B.n612 10.6151
R2091 B.n612 B.n611 10.6151
R2092 B.n611 B.n80 10.6151
R2093 B.n607 B.n80 10.6151
R2094 B.n607 B.n606 10.6151
R2095 B.n606 B.n605 10.6151
R2096 B.n605 B.n82 10.6151
R2097 B.n601 B.n82 10.6151
R2098 B.n601 B.n600 10.6151
R2099 B.n600 B.n599 10.6151
R2100 B.n599 B.n84 10.6151
R2101 B.n451 B.n132 10.6151
R2102 B.n455 B.n132 10.6151
R2103 B.n456 B.n455 10.6151
R2104 B.n457 B.n456 10.6151
R2105 B.n457 B.n130 10.6151
R2106 B.n461 B.n130 10.6151
R2107 B.n462 B.n461 10.6151
R2108 B.n463 B.n462 10.6151
R2109 B.n463 B.n128 10.6151
R2110 B.n467 B.n128 10.6151
R2111 B.n468 B.n467 10.6151
R2112 B.n469 B.n468 10.6151
R2113 B.n469 B.n126 10.6151
R2114 B.n473 B.n126 10.6151
R2115 B.n474 B.n473 10.6151
R2116 B.n475 B.n474 10.6151
R2117 B.n475 B.n124 10.6151
R2118 B.n479 B.n124 10.6151
R2119 B.n480 B.n479 10.6151
R2120 B.n481 B.n480 10.6151
R2121 B.n481 B.n122 10.6151
R2122 B.n485 B.n122 10.6151
R2123 B.n486 B.n485 10.6151
R2124 B.n487 B.n486 10.6151
R2125 B.n487 B.n120 10.6151
R2126 B.n491 B.n120 10.6151
R2127 B.n492 B.n491 10.6151
R2128 B.n493 B.n492 10.6151
R2129 B.n493 B.n118 10.6151
R2130 B.n497 B.n118 10.6151
R2131 B.n498 B.n497 10.6151
R2132 B.n499 B.n498 10.6151
R2133 B.n499 B.n116 10.6151
R2134 B.n503 B.n116 10.6151
R2135 B.n504 B.n503 10.6151
R2136 B.n505 B.n504 10.6151
R2137 B.n505 B.n114 10.6151
R2138 B.n509 B.n114 10.6151
R2139 B.n510 B.n509 10.6151
R2140 B.n511 B.n510 10.6151
R2141 B.n511 B.n112 10.6151
R2142 B.n515 B.n112 10.6151
R2143 B.n516 B.n515 10.6151
R2144 B.n517 B.n516 10.6151
R2145 B.n517 B.n110 10.6151
R2146 B.n521 B.n110 10.6151
R2147 B.n522 B.n521 10.6151
R2148 B.n523 B.n522 10.6151
R2149 B.n523 B.n108 10.6151
R2150 B.n527 B.n108 10.6151
R2151 B.n528 B.n527 10.6151
R2152 B.n529 B.n528 10.6151
R2153 B.n529 B.n106 10.6151
R2154 B.n533 B.n106 10.6151
R2155 B.n534 B.n533 10.6151
R2156 B.n535 B.n534 10.6151
R2157 B.n535 B.n104 10.6151
R2158 B.n539 B.n104 10.6151
R2159 B.n540 B.n539 10.6151
R2160 B.n541 B.n540 10.6151
R2161 B.n541 B.n102 10.6151
R2162 B.n545 B.n102 10.6151
R2163 B.n546 B.n545 10.6151
R2164 B.n547 B.n546 10.6151
R2165 B.n547 B.n100 10.6151
R2166 B.n551 B.n100 10.6151
R2167 B.n552 B.n551 10.6151
R2168 B.n553 B.n552 10.6151
R2169 B.n553 B.n98 10.6151
R2170 B.n557 B.n98 10.6151
R2171 B.n558 B.n557 10.6151
R2172 B.n559 B.n558 10.6151
R2173 B.n559 B.n96 10.6151
R2174 B.n563 B.n96 10.6151
R2175 B.n564 B.n563 10.6151
R2176 B.n565 B.n564 10.6151
R2177 B.n565 B.n94 10.6151
R2178 B.n569 B.n94 10.6151
R2179 B.n570 B.n569 10.6151
R2180 B.n571 B.n570 10.6151
R2181 B.n571 B.n92 10.6151
R2182 B.n575 B.n92 10.6151
R2183 B.n576 B.n575 10.6151
R2184 B.n577 B.n576 10.6151
R2185 B.n577 B.n90 10.6151
R2186 B.n581 B.n90 10.6151
R2187 B.n582 B.n581 10.6151
R2188 B.n583 B.n582 10.6151
R2189 B.n583 B.n88 10.6151
R2190 B.n587 B.n88 10.6151
R2191 B.n588 B.n587 10.6151
R2192 B.n589 B.n588 10.6151
R2193 B.n589 B.n86 10.6151
R2194 B.n593 B.n86 10.6151
R2195 B.n594 B.n593 10.6151
R2196 B.n595 B.n594 10.6151
R2197 B.n288 B.n287 10.6151
R2198 B.n289 B.n288 10.6151
R2199 B.n289 B.n190 10.6151
R2200 B.n293 B.n190 10.6151
R2201 B.n294 B.n293 10.6151
R2202 B.n295 B.n294 10.6151
R2203 B.n295 B.n188 10.6151
R2204 B.n299 B.n188 10.6151
R2205 B.n300 B.n299 10.6151
R2206 B.n301 B.n300 10.6151
R2207 B.n301 B.n186 10.6151
R2208 B.n305 B.n186 10.6151
R2209 B.n306 B.n305 10.6151
R2210 B.n307 B.n306 10.6151
R2211 B.n307 B.n184 10.6151
R2212 B.n311 B.n184 10.6151
R2213 B.n312 B.n311 10.6151
R2214 B.n313 B.n312 10.6151
R2215 B.n313 B.n182 10.6151
R2216 B.n317 B.n182 10.6151
R2217 B.n318 B.n317 10.6151
R2218 B.n319 B.n318 10.6151
R2219 B.n319 B.n180 10.6151
R2220 B.n323 B.n180 10.6151
R2221 B.n324 B.n323 10.6151
R2222 B.n325 B.n324 10.6151
R2223 B.n325 B.n178 10.6151
R2224 B.n329 B.n178 10.6151
R2225 B.n330 B.n329 10.6151
R2226 B.n331 B.n330 10.6151
R2227 B.n331 B.n176 10.6151
R2228 B.n335 B.n176 10.6151
R2229 B.n336 B.n335 10.6151
R2230 B.n337 B.n336 10.6151
R2231 B.n337 B.n174 10.6151
R2232 B.n341 B.n174 10.6151
R2233 B.n342 B.n341 10.6151
R2234 B.n343 B.n342 10.6151
R2235 B.n343 B.n172 10.6151
R2236 B.n347 B.n172 10.6151
R2237 B.n348 B.n347 10.6151
R2238 B.n349 B.n348 10.6151
R2239 B.n349 B.n170 10.6151
R2240 B.n353 B.n170 10.6151
R2241 B.n354 B.n353 10.6151
R2242 B.n355 B.n354 10.6151
R2243 B.n355 B.n168 10.6151
R2244 B.n359 B.n168 10.6151
R2245 B.n360 B.n359 10.6151
R2246 B.n362 B.n164 10.6151
R2247 B.n366 B.n164 10.6151
R2248 B.n367 B.n366 10.6151
R2249 B.n368 B.n367 10.6151
R2250 B.n368 B.n162 10.6151
R2251 B.n372 B.n162 10.6151
R2252 B.n373 B.n372 10.6151
R2253 B.n374 B.n373 10.6151
R2254 B.n378 B.n377 10.6151
R2255 B.n379 B.n378 10.6151
R2256 B.n379 B.n156 10.6151
R2257 B.n383 B.n156 10.6151
R2258 B.n384 B.n383 10.6151
R2259 B.n385 B.n384 10.6151
R2260 B.n385 B.n154 10.6151
R2261 B.n389 B.n154 10.6151
R2262 B.n390 B.n389 10.6151
R2263 B.n391 B.n390 10.6151
R2264 B.n391 B.n152 10.6151
R2265 B.n395 B.n152 10.6151
R2266 B.n396 B.n395 10.6151
R2267 B.n397 B.n396 10.6151
R2268 B.n397 B.n150 10.6151
R2269 B.n401 B.n150 10.6151
R2270 B.n402 B.n401 10.6151
R2271 B.n403 B.n402 10.6151
R2272 B.n403 B.n148 10.6151
R2273 B.n407 B.n148 10.6151
R2274 B.n408 B.n407 10.6151
R2275 B.n409 B.n408 10.6151
R2276 B.n409 B.n146 10.6151
R2277 B.n413 B.n146 10.6151
R2278 B.n414 B.n413 10.6151
R2279 B.n415 B.n414 10.6151
R2280 B.n415 B.n144 10.6151
R2281 B.n419 B.n144 10.6151
R2282 B.n420 B.n419 10.6151
R2283 B.n421 B.n420 10.6151
R2284 B.n421 B.n142 10.6151
R2285 B.n425 B.n142 10.6151
R2286 B.n426 B.n425 10.6151
R2287 B.n427 B.n426 10.6151
R2288 B.n427 B.n140 10.6151
R2289 B.n431 B.n140 10.6151
R2290 B.n432 B.n431 10.6151
R2291 B.n433 B.n432 10.6151
R2292 B.n433 B.n138 10.6151
R2293 B.n437 B.n138 10.6151
R2294 B.n438 B.n437 10.6151
R2295 B.n439 B.n438 10.6151
R2296 B.n439 B.n136 10.6151
R2297 B.n443 B.n136 10.6151
R2298 B.n444 B.n443 10.6151
R2299 B.n445 B.n444 10.6151
R2300 B.n445 B.n134 10.6151
R2301 B.n449 B.n134 10.6151
R2302 B.n450 B.n449 10.6151
R2303 B.n283 B.n192 10.6151
R2304 B.n283 B.n282 10.6151
R2305 B.n282 B.n281 10.6151
R2306 B.n281 B.n194 10.6151
R2307 B.n277 B.n194 10.6151
R2308 B.n277 B.n276 10.6151
R2309 B.n276 B.n275 10.6151
R2310 B.n275 B.n196 10.6151
R2311 B.n271 B.n196 10.6151
R2312 B.n271 B.n270 10.6151
R2313 B.n270 B.n269 10.6151
R2314 B.n269 B.n198 10.6151
R2315 B.n265 B.n198 10.6151
R2316 B.n265 B.n264 10.6151
R2317 B.n264 B.n263 10.6151
R2318 B.n263 B.n200 10.6151
R2319 B.n259 B.n200 10.6151
R2320 B.n259 B.n258 10.6151
R2321 B.n258 B.n257 10.6151
R2322 B.n257 B.n202 10.6151
R2323 B.n253 B.n202 10.6151
R2324 B.n253 B.n252 10.6151
R2325 B.n252 B.n251 10.6151
R2326 B.n251 B.n204 10.6151
R2327 B.n247 B.n204 10.6151
R2328 B.n247 B.n246 10.6151
R2329 B.n246 B.n245 10.6151
R2330 B.n245 B.n206 10.6151
R2331 B.n241 B.n206 10.6151
R2332 B.n241 B.n240 10.6151
R2333 B.n240 B.n239 10.6151
R2334 B.n239 B.n208 10.6151
R2335 B.n235 B.n208 10.6151
R2336 B.n235 B.n234 10.6151
R2337 B.n234 B.n233 10.6151
R2338 B.n233 B.n210 10.6151
R2339 B.n229 B.n210 10.6151
R2340 B.n229 B.n228 10.6151
R2341 B.n228 B.n227 10.6151
R2342 B.n227 B.n212 10.6151
R2343 B.n223 B.n212 10.6151
R2344 B.n223 B.n222 10.6151
R2345 B.n222 B.n221 10.6151
R2346 B.n221 B.n214 10.6151
R2347 B.n217 B.n214 10.6151
R2348 B.n217 B.n216 10.6151
R2349 B.n216 B.n0 10.6151
R2350 B.n831 B.n1 10.6151
R2351 B.n831 B.n830 10.6151
R2352 B.n830 B.n829 10.6151
R2353 B.n829 B.n4 10.6151
R2354 B.n825 B.n4 10.6151
R2355 B.n825 B.n824 10.6151
R2356 B.n824 B.n823 10.6151
R2357 B.n823 B.n6 10.6151
R2358 B.n819 B.n6 10.6151
R2359 B.n819 B.n818 10.6151
R2360 B.n818 B.n817 10.6151
R2361 B.n817 B.n8 10.6151
R2362 B.n813 B.n8 10.6151
R2363 B.n813 B.n812 10.6151
R2364 B.n812 B.n811 10.6151
R2365 B.n811 B.n10 10.6151
R2366 B.n807 B.n10 10.6151
R2367 B.n807 B.n806 10.6151
R2368 B.n806 B.n805 10.6151
R2369 B.n805 B.n12 10.6151
R2370 B.n801 B.n12 10.6151
R2371 B.n801 B.n800 10.6151
R2372 B.n800 B.n799 10.6151
R2373 B.n799 B.n14 10.6151
R2374 B.n795 B.n14 10.6151
R2375 B.n795 B.n794 10.6151
R2376 B.n794 B.n793 10.6151
R2377 B.n793 B.n16 10.6151
R2378 B.n789 B.n16 10.6151
R2379 B.n789 B.n788 10.6151
R2380 B.n788 B.n787 10.6151
R2381 B.n787 B.n18 10.6151
R2382 B.n783 B.n18 10.6151
R2383 B.n783 B.n782 10.6151
R2384 B.n782 B.n781 10.6151
R2385 B.n781 B.n20 10.6151
R2386 B.n777 B.n20 10.6151
R2387 B.n777 B.n776 10.6151
R2388 B.n776 B.n775 10.6151
R2389 B.n775 B.n22 10.6151
R2390 B.n771 B.n22 10.6151
R2391 B.n771 B.n770 10.6151
R2392 B.n770 B.n769 10.6151
R2393 B.n769 B.n24 10.6151
R2394 B.n765 B.n24 10.6151
R2395 B.n765 B.n764 10.6151
R2396 B.n764 B.n763 10.6151
R2397 B.n686 B.n685 6.5566
R2398 B.n673 B.n672 6.5566
R2399 B.n362 B.n361 6.5566
R2400 B.n374 B.n160 6.5566
R2401 B.n687 B.n686 4.05904
R2402 B.n672 B.n671 4.05904
R2403 B.n361 B.n360 4.05904
R2404 B.n377 B.n160 4.05904
R2405 B.n835 B.n0 2.81026
R2406 B.n835 B.n1 2.81026
C0 VN VDD2 8.448429f
C1 VN VTAIL 8.58813f
C2 B w_n3674_n3932# 11.0885f
C3 VP w_n3674_n3932# 7.59178f
C4 VDD1 w_n3674_n3932# 2.59626f
C5 VDD2 w_n3674_n3932# 2.6957f
C6 B VP 2.09676f
C7 B VDD1 2.43591f
C8 VTAIL w_n3674_n3932# 3.40249f
C9 VP VDD1 8.79021f
C10 B VDD2 2.52079f
C11 VN w_n3674_n3932# 7.11553f
C12 VP VDD2 0.497091f
C13 VTAIL B 4.52026f
C14 VDD1 VDD2 1.58336f
C15 VTAIL VP 8.60242f
C16 VTAIL VDD1 8.80954f
C17 VN B 1.29934f
C18 VTAIL VDD2 8.86327f
C19 VN VP 7.88313f
C20 VN VDD1 0.151775f
C21 VDD2 VSUBS 2.085461f
C22 VDD1 VSUBS 2.063069f
C23 VTAIL VSUBS 1.383891f
C24 VN VSUBS 6.37229f
C25 VP VSUBS 3.398517f
C26 B VSUBS 5.321308f
C27 w_n3674_n3932# VSUBS 0.17719p
C28 B.n0 VSUBS 0.00508f
C29 B.n1 VSUBS 0.00508f
C30 B.n2 VSUBS 0.008034f
C31 B.n3 VSUBS 0.008034f
C32 B.n4 VSUBS 0.008034f
C33 B.n5 VSUBS 0.008034f
C34 B.n6 VSUBS 0.008034f
C35 B.n7 VSUBS 0.008034f
C36 B.n8 VSUBS 0.008034f
C37 B.n9 VSUBS 0.008034f
C38 B.n10 VSUBS 0.008034f
C39 B.n11 VSUBS 0.008034f
C40 B.n12 VSUBS 0.008034f
C41 B.n13 VSUBS 0.008034f
C42 B.n14 VSUBS 0.008034f
C43 B.n15 VSUBS 0.008034f
C44 B.n16 VSUBS 0.008034f
C45 B.n17 VSUBS 0.008034f
C46 B.n18 VSUBS 0.008034f
C47 B.n19 VSUBS 0.008034f
C48 B.n20 VSUBS 0.008034f
C49 B.n21 VSUBS 0.008034f
C50 B.n22 VSUBS 0.008034f
C51 B.n23 VSUBS 0.008034f
C52 B.n24 VSUBS 0.008034f
C53 B.n25 VSUBS 0.008034f
C54 B.n26 VSUBS 0.019215f
C55 B.n27 VSUBS 0.008034f
C56 B.n28 VSUBS 0.008034f
C57 B.n29 VSUBS 0.008034f
C58 B.n30 VSUBS 0.008034f
C59 B.n31 VSUBS 0.008034f
C60 B.n32 VSUBS 0.008034f
C61 B.n33 VSUBS 0.008034f
C62 B.n34 VSUBS 0.008034f
C63 B.n35 VSUBS 0.008034f
C64 B.n36 VSUBS 0.008034f
C65 B.n37 VSUBS 0.008034f
C66 B.n38 VSUBS 0.008034f
C67 B.n39 VSUBS 0.008034f
C68 B.n40 VSUBS 0.008034f
C69 B.n41 VSUBS 0.008034f
C70 B.n42 VSUBS 0.008034f
C71 B.n43 VSUBS 0.008034f
C72 B.n44 VSUBS 0.008034f
C73 B.n45 VSUBS 0.008034f
C74 B.n46 VSUBS 0.008034f
C75 B.n47 VSUBS 0.008034f
C76 B.n48 VSUBS 0.008034f
C77 B.n49 VSUBS 0.008034f
C78 B.n50 VSUBS 0.008034f
C79 B.n51 VSUBS 0.008034f
C80 B.t8 VSUBS 0.31615f
C81 B.t7 VSUBS 0.359155f
C82 B.t6 VSUBS 2.35755f
C83 B.n52 VSUBS 0.565733f
C84 B.n53 VSUBS 0.334244f
C85 B.n54 VSUBS 0.008034f
C86 B.n55 VSUBS 0.008034f
C87 B.n56 VSUBS 0.008034f
C88 B.n57 VSUBS 0.008034f
C89 B.t11 VSUBS 0.316153f
C90 B.t10 VSUBS 0.359158f
C91 B.t9 VSUBS 2.35755f
C92 B.n58 VSUBS 0.56573f
C93 B.n59 VSUBS 0.33424f
C94 B.n60 VSUBS 0.008034f
C95 B.n61 VSUBS 0.008034f
C96 B.n62 VSUBS 0.008034f
C97 B.n63 VSUBS 0.008034f
C98 B.n64 VSUBS 0.008034f
C99 B.n65 VSUBS 0.008034f
C100 B.n66 VSUBS 0.008034f
C101 B.n67 VSUBS 0.008034f
C102 B.n68 VSUBS 0.008034f
C103 B.n69 VSUBS 0.008034f
C104 B.n70 VSUBS 0.008034f
C105 B.n71 VSUBS 0.008034f
C106 B.n72 VSUBS 0.008034f
C107 B.n73 VSUBS 0.008034f
C108 B.n74 VSUBS 0.008034f
C109 B.n75 VSUBS 0.008034f
C110 B.n76 VSUBS 0.008034f
C111 B.n77 VSUBS 0.008034f
C112 B.n78 VSUBS 0.008034f
C113 B.n79 VSUBS 0.008034f
C114 B.n80 VSUBS 0.008034f
C115 B.n81 VSUBS 0.008034f
C116 B.n82 VSUBS 0.008034f
C117 B.n83 VSUBS 0.008034f
C118 B.n84 VSUBS 0.018283f
C119 B.n85 VSUBS 0.008034f
C120 B.n86 VSUBS 0.008034f
C121 B.n87 VSUBS 0.008034f
C122 B.n88 VSUBS 0.008034f
C123 B.n89 VSUBS 0.008034f
C124 B.n90 VSUBS 0.008034f
C125 B.n91 VSUBS 0.008034f
C126 B.n92 VSUBS 0.008034f
C127 B.n93 VSUBS 0.008034f
C128 B.n94 VSUBS 0.008034f
C129 B.n95 VSUBS 0.008034f
C130 B.n96 VSUBS 0.008034f
C131 B.n97 VSUBS 0.008034f
C132 B.n98 VSUBS 0.008034f
C133 B.n99 VSUBS 0.008034f
C134 B.n100 VSUBS 0.008034f
C135 B.n101 VSUBS 0.008034f
C136 B.n102 VSUBS 0.008034f
C137 B.n103 VSUBS 0.008034f
C138 B.n104 VSUBS 0.008034f
C139 B.n105 VSUBS 0.008034f
C140 B.n106 VSUBS 0.008034f
C141 B.n107 VSUBS 0.008034f
C142 B.n108 VSUBS 0.008034f
C143 B.n109 VSUBS 0.008034f
C144 B.n110 VSUBS 0.008034f
C145 B.n111 VSUBS 0.008034f
C146 B.n112 VSUBS 0.008034f
C147 B.n113 VSUBS 0.008034f
C148 B.n114 VSUBS 0.008034f
C149 B.n115 VSUBS 0.008034f
C150 B.n116 VSUBS 0.008034f
C151 B.n117 VSUBS 0.008034f
C152 B.n118 VSUBS 0.008034f
C153 B.n119 VSUBS 0.008034f
C154 B.n120 VSUBS 0.008034f
C155 B.n121 VSUBS 0.008034f
C156 B.n122 VSUBS 0.008034f
C157 B.n123 VSUBS 0.008034f
C158 B.n124 VSUBS 0.008034f
C159 B.n125 VSUBS 0.008034f
C160 B.n126 VSUBS 0.008034f
C161 B.n127 VSUBS 0.008034f
C162 B.n128 VSUBS 0.008034f
C163 B.n129 VSUBS 0.008034f
C164 B.n130 VSUBS 0.008034f
C165 B.n131 VSUBS 0.008034f
C166 B.n132 VSUBS 0.008034f
C167 B.n133 VSUBS 0.019215f
C168 B.n134 VSUBS 0.008034f
C169 B.n135 VSUBS 0.008034f
C170 B.n136 VSUBS 0.008034f
C171 B.n137 VSUBS 0.008034f
C172 B.n138 VSUBS 0.008034f
C173 B.n139 VSUBS 0.008034f
C174 B.n140 VSUBS 0.008034f
C175 B.n141 VSUBS 0.008034f
C176 B.n142 VSUBS 0.008034f
C177 B.n143 VSUBS 0.008034f
C178 B.n144 VSUBS 0.008034f
C179 B.n145 VSUBS 0.008034f
C180 B.n146 VSUBS 0.008034f
C181 B.n147 VSUBS 0.008034f
C182 B.n148 VSUBS 0.008034f
C183 B.n149 VSUBS 0.008034f
C184 B.n150 VSUBS 0.008034f
C185 B.n151 VSUBS 0.008034f
C186 B.n152 VSUBS 0.008034f
C187 B.n153 VSUBS 0.008034f
C188 B.n154 VSUBS 0.008034f
C189 B.n155 VSUBS 0.008034f
C190 B.n156 VSUBS 0.008034f
C191 B.n157 VSUBS 0.008034f
C192 B.t4 VSUBS 0.316153f
C193 B.t5 VSUBS 0.359158f
C194 B.t3 VSUBS 2.35755f
C195 B.n158 VSUBS 0.56573f
C196 B.n159 VSUBS 0.33424f
C197 B.n160 VSUBS 0.018614f
C198 B.n161 VSUBS 0.008034f
C199 B.n162 VSUBS 0.008034f
C200 B.n163 VSUBS 0.008034f
C201 B.n164 VSUBS 0.008034f
C202 B.n165 VSUBS 0.008034f
C203 B.t1 VSUBS 0.31615f
C204 B.t2 VSUBS 0.359155f
C205 B.t0 VSUBS 2.35755f
C206 B.n166 VSUBS 0.565733f
C207 B.n167 VSUBS 0.334244f
C208 B.n168 VSUBS 0.008034f
C209 B.n169 VSUBS 0.008034f
C210 B.n170 VSUBS 0.008034f
C211 B.n171 VSUBS 0.008034f
C212 B.n172 VSUBS 0.008034f
C213 B.n173 VSUBS 0.008034f
C214 B.n174 VSUBS 0.008034f
C215 B.n175 VSUBS 0.008034f
C216 B.n176 VSUBS 0.008034f
C217 B.n177 VSUBS 0.008034f
C218 B.n178 VSUBS 0.008034f
C219 B.n179 VSUBS 0.008034f
C220 B.n180 VSUBS 0.008034f
C221 B.n181 VSUBS 0.008034f
C222 B.n182 VSUBS 0.008034f
C223 B.n183 VSUBS 0.008034f
C224 B.n184 VSUBS 0.008034f
C225 B.n185 VSUBS 0.008034f
C226 B.n186 VSUBS 0.008034f
C227 B.n187 VSUBS 0.008034f
C228 B.n188 VSUBS 0.008034f
C229 B.n189 VSUBS 0.008034f
C230 B.n190 VSUBS 0.008034f
C231 B.n191 VSUBS 0.008034f
C232 B.n192 VSUBS 0.018829f
C233 B.n193 VSUBS 0.008034f
C234 B.n194 VSUBS 0.008034f
C235 B.n195 VSUBS 0.008034f
C236 B.n196 VSUBS 0.008034f
C237 B.n197 VSUBS 0.008034f
C238 B.n198 VSUBS 0.008034f
C239 B.n199 VSUBS 0.008034f
C240 B.n200 VSUBS 0.008034f
C241 B.n201 VSUBS 0.008034f
C242 B.n202 VSUBS 0.008034f
C243 B.n203 VSUBS 0.008034f
C244 B.n204 VSUBS 0.008034f
C245 B.n205 VSUBS 0.008034f
C246 B.n206 VSUBS 0.008034f
C247 B.n207 VSUBS 0.008034f
C248 B.n208 VSUBS 0.008034f
C249 B.n209 VSUBS 0.008034f
C250 B.n210 VSUBS 0.008034f
C251 B.n211 VSUBS 0.008034f
C252 B.n212 VSUBS 0.008034f
C253 B.n213 VSUBS 0.008034f
C254 B.n214 VSUBS 0.008034f
C255 B.n215 VSUBS 0.008034f
C256 B.n216 VSUBS 0.008034f
C257 B.n217 VSUBS 0.008034f
C258 B.n218 VSUBS 0.008034f
C259 B.n219 VSUBS 0.008034f
C260 B.n220 VSUBS 0.008034f
C261 B.n221 VSUBS 0.008034f
C262 B.n222 VSUBS 0.008034f
C263 B.n223 VSUBS 0.008034f
C264 B.n224 VSUBS 0.008034f
C265 B.n225 VSUBS 0.008034f
C266 B.n226 VSUBS 0.008034f
C267 B.n227 VSUBS 0.008034f
C268 B.n228 VSUBS 0.008034f
C269 B.n229 VSUBS 0.008034f
C270 B.n230 VSUBS 0.008034f
C271 B.n231 VSUBS 0.008034f
C272 B.n232 VSUBS 0.008034f
C273 B.n233 VSUBS 0.008034f
C274 B.n234 VSUBS 0.008034f
C275 B.n235 VSUBS 0.008034f
C276 B.n236 VSUBS 0.008034f
C277 B.n237 VSUBS 0.008034f
C278 B.n238 VSUBS 0.008034f
C279 B.n239 VSUBS 0.008034f
C280 B.n240 VSUBS 0.008034f
C281 B.n241 VSUBS 0.008034f
C282 B.n242 VSUBS 0.008034f
C283 B.n243 VSUBS 0.008034f
C284 B.n244 VSUBS 0.008034f
C285 B.n245 VSUBS 0.008034f
C286 B.n246 VSUBS 0.008034f
C287 B.n247 VSUBS 0.008034f
C288 B.n248 VSUBS 0.008034f
C289 B.n249 VSUBS 0.008034f
C290 B.n250 VSUBS 0.008034f
C291 B.n251 VSUBS 0.008034f
C292 B.n252 VSUBS 0.008034f
C293 B.n253 VSUBS 0.008034f
C294 B.n254 VSUBS 0.008034f
C295 B.n255 VSUBS 0.008034f
C296 B.n256 VSUBS 0.008034f
C297 B.n257 VSUBS 0.008034f
C298 B.n258 VSUBS 0.008034f
C299 B.n259 VSUBS 0.008034f
C300 B.n260 VSUBS 0.008034f
C301 B.n261 VSUBS 0.008034f
C302 B.n262 VSUBS 0.008034f
C303 B.n263 VSUBS 0.008034f
C304 B.n264 VSUBS 0.008034f
C305 B.n265 VSUBS 0.008034f
C306 B.n266 VSUBS 0.008034f
C307 B.n267 VSUBS 0.008034f
C308 B.n268 VSUBS 0.008034f
C309 B.n269 VSUBS 0.008034f
C310 B.n270 VSUBS 0.008034f
C311 B.n271 VSUBS 0.008034f
C312 B.n272 VSUBS 0.008034f
C313 B.n273 VSUBS 0.008034f
C314 B.n274 VSUBS 0.008034f
C315 B.n275 VSUBS 0.008034f
C316 B.n276 VSUBS 0.008034f
C317 B.n277 VSUBS 0.008034f
C318 B.n278 VSUBS 0.008034f
C319 B.n279 VSUBS 0.008034f
C320 B.n280 VSUBS 0.008034f
C321 B.n281 VSUBS 0.008034f
C322 B.n282 VSUBS 0.008034f
C323 B.n283 VSUBS 0.008034f
C324 B.n284 VSUBS 0.008034f
C325 B.n285 VSUBS 0.018829f
C326 B.n286 VSUBS 0.019215f
C327 B.n287 VSUBS 0.019215f
C328 B.n288 VSUBS 0.008034f
C329 B.n289 VSUBS 0.008034f
C330 B.n290 VSUBS 0.008034f
C331 B.n291 VSUBS 0.008034f
C332 B.n292 VSUBS 0.008034f
C333 B.n293 VSUBS 0.008034f
C334 B.n294 VSUBS 0.008034f
C335 B.n295 VSUBS 0.008034f
C336 B.n296 VSUBS 0.008034f
C337 B.n297 VSUBS 0.008034f
C338 B.n298 VSUBS 0.008034f
C339 B.n299 VSUBS 0.008034f
C340 B.n300 VSUBS 0.008034f
C341 B.n301 VSUBS 0.008034f
C342 B.n302 VSUBS 0.008034f
C343 B.n303 VSUBS 0.008034f
C344 B.n304 VSUBS 0.008034f
C345 B.n305 VSUBS 0.008034f
C346 B.n306 VSUBS 0.008034f
C347 B.n307 VSUBS 0.008034f
C348 B.n308 VSUBS 0.008034f
C349 B.n309 VSUBS 0.008034f
C350 B.n310 VSUBS 0.008034f
C351 B.n311 VSUBS 0.008034f
C352 B.n312 VSUBS 0.008034f
C353 B.n313 VSUBS 0.008034f
C354 B.n314 VSUBS 0.008034f
C355 B.n315 VSUBS 0.008034f
C356 B.n316 VSUBS 0.008034f
C357 B.n317 VSUBS 0.008034f
C358 B.n318 VSUBS 0.008034f
C359 B.n319 VSUBS 0.008034f
C360 B.n320 VSUBS 0.008034f
C361 B.n321 VSUBS 0.008034f
C362 B.n322 VSUBS 0.008034f
C363 B.n323 VSUBS 0.008034f
C364 B.n324 VSUBS 0.008034f
C365 B.n325 VSUBS 0.008034f
C366 B.n326 VSUBS 0.008034f
C367 B.n327 VSUBS 0.008034f
C368 B.n328 VSUBS 0.008034f
C369 B.n329 VSUBS 0.008034f
C370 B.n330 VSUBS 0.008034f
C371 B.n331 VSUBS 0.008034f
C372 B.n332 VSUBS 0.008034f
C373 B.n333 VSUBS 0.008034f
C374 B.n334 VSUBS 0.008034f
C375 B.n335 VSUBS 0.008034f
C376 B.n336 VSUBS 0.008034f
C377 B.n337 VSUBS 0.008034f
C378 B.n338 VSUBS 0.008034f
C379 B.n339 VSUBS 0.008034f
C380 B.n340 VSUBS 0.008034f
C381 B.n341 VSUBS 0.008034f
C382 B.n342 VSUBS 0.008034f
C383 B.n343 VSUBS 0.008034f
C384 B.n344 VSUBS 0.008034f
C385 B.n345 VSUBS 0.008034f
C386 B.n346 VSUBS 0.008034f
C387 B.n347 VSUBS 0.008034f
C388 B.n348 VSUBS 0.008034f
C389 B.n349 VSUBS 0.008034f
C390 B.n350 VSUBS 0.008034f
C391 B.n351 VSUBS 0.008034f
C392 B.n352 VSUBS 0.008034f
C393 B.n353 VSUBS 0.008034f
C394 B.n354 VSUBS 0.008034f
C395 B.n355 VSUBS 0.008034f
C396 B.n356 VSUBS 0.008034f
C397 B.n357 VSUBS 0.008034f
C398 B.n358 VSUBS 0.008034f
C399 B.n359 VSUBS 0.008034f
C400 B.n360 VSUBS 0.005553f
C401 B.n361 VSUBS 0.018614f
C402 B.n362 VSUBS 0.006498f
C403 B.n363 VSUBS 0.008034f
C404 B.n364 VSUBS 0.008034f
C405 B.n365 VSUBS 0.008034f
C406 B.n366 VSUBS 0.008034f
C407 B.n367 VSUBS 0.008034f
C408 B.n368 VSUBS 0.008034f
C409 B.n369 VSUBS 0.008034f
C410 B.n370 VSUBS 0.008034f
C411 B.n371 VSUBS 0.008034f
C412 B.n372 VSUBS 0.008034f
C413 B.n373 VSUBS 0.008034f
C414 B.n374 VSUBS 0.006498f
C415 B.n375 VSUBS 0.008034f
C416 B.n376 VSUBS 0.008034f
C417 B.n377 VSUBS 0.005553f
C418 B.n378 VSUBS 0.008034f
C419 B.n379 VSUBS 0.008034f
C420 B.n380 VSUBS 0.008034f
C421 B.n381 VSUBS 0.008034f
C422 B.n382 VSUBS 0.008034f
C423 B.n383 VSUBS 0.008034f
C424 B.n384 VSUBS 0.008034f
C425 B.n385 VSUBS 0.008034f
C426 B.n386 VSUBS 0.008034f
C427 B.n387 VSUBS 0.008034f
C428 B.n388 VSUBS 0.008034f
C429 B.n389 VSUBS 0.008034f
C430 B.n390 VSUBS 0.008034f
C431 B.n391 VSUBS 0.008034f
C432 B.n392 VSUBS 0.008034f
C433 B.n393 VSUBS 0.008034f
C434 B.n394 VSUBS 0.008034f
C435 B.n395 VSUBS 0.008034f
C436 B.n396 VSUBS 0.008034f
C437 B.n397 VSUBS 0.008034f
C438 B.n398 VSUBS 0.008034f
C439 B.n399 VSUBS 0.008034f
C440 B.n400 VSUBS 0.008034f
C441 B.n401 VSUBS 0.008034f
C442 B.n402 VSUBS 0.008034f
C443 B.n403 VSUBS 0.008034f
C444 B.n404 VSUBS 0.008034f
C445 B.n405 VSUBS 0.008034f
C446 B.n406 VSUBS 0.008034f
C447 B.n407 VSUBS 0.008034f
C448 B.n408 VSUBS 0.008034f
C449 B.n409 VSUBS 0.008034f
C450 B.n410 VSUBS 0.008034f
C451 B.n411 VSUBS 0.008034f
C452 B.n412 VSUBS 0.008034f
C453 B.n413 VSUBS 0.008034f
C454 B.n414 VSUBS 0.008034f
C455 B.n415 VSUBS 0.008034f
C456 B.n416 VSUBS 0.008034f
C457 B.n417 VSUBS 0.008034f
C458 B.n418 VSUBS 0.008034f
C459 B.n419 VSUBS 0.008034f
C460 B.n420 VSUBS 0.008034f
C461 B.n421 VSUBS 0.008034f
C462 B.n422 VSUBS 0.008034f
C463 B.n423 VSUBS 0.008034f
C464 B.n424 VSUBS 0.008034f
C465 B.n425 VSUBS 0.008034f
C466 B.n426 VSUBS 0.008034f
C467 B.n427 VSUBS 0.008034f
C468 B.n428 VSUBS 0.008034f
C469 B.n429 VSUBS 0.008034f
C470 B.n430 VSUBS 0.008034f
C471 B.n431 VSUBS 0.008034f
C472 B.n432 VSUBS 0.008034f
C473 B.n433 VSUBS 0.008034f
C474 B.n434 VSUBS 0.008034f
C475 B.n435 VSUBS 0.008034f
C476 B.n436 VSUBS 0.008034f
C477 B.n437 VSUBS 0.008034f
C478 B.n438 VSUBS 0.008034f
C479 B.n439 VSUBS 0.008034f
C480 B.n440 VSUBS 0.008034f
C481 B.n441 VSUBS 0.008034f
C482 B.n442 VSUBS 0.008034f
C483 B.n443 VSUBS 0.008034f
C484 B.n444 VSUBS 0.008034f
C485 B.n445 VSUBS 0.008034f
C486 B.n446 VSUBS 0.008034f
C487 B.n447 VSUBS 0.008034f
C488 B.n448 VSUBS 0.008034f
C489 B.n449 VSUBS 0.008034f
C490 B.n450 VSUBS 0.019215f
C491 B.n451 VSUBS 0.018829f
C492 B.n452 VSUBS 0.018829f
C493 B.n453 VSUBS 0.008034f
C494 B.n454 VSUBS 0.008034f
C495 B.n455 VSUBS 0.008034f
C496 B.n456 VSUBS 0.008034f
C497 B.n457 VSUBS 0.008034f
C498 B.n458 VSUBS 0.008034f
C499 B.n459 VSUBS 0.008034f
C500 B.n460 VSUBS 0.008034f
C501 B.n461 VSUBS 0.008034f
C502 B.n462 VSUBS 0.008034f
C503 B.n463 VSUBS 0.008034f
C504 B.n464 VSUBS 0.008034f
C505 B.n465 VSUBS 0.008034f
C506 B.n466 VSUBS 0.008034f
C507 B.n467 VSUBS 0.008034f
C508 B.n468 VSUBS 0.008034f
C509 B.n469 VSUBS 0.008034f
C510 B.n470 VSUBS 0.008034f
C511 B.n471 VSUBS 0.008034f
C512 B.n472 VSUBS 0.008034f
C513 B.n473 VSUBS 0.008034f
C514 B.n474 VSUBS 0.008034f
C515 B.n475 VSUBS 0.008034f
C516 B.n476 VSUBS 0.008034f
C517 B.n477 VSUBS 0.008034f
C518 B.n478 VSUBS 0.008034f
C519 B.n479 VSUBS 0.008034f
C520 B.n480 VSUBS 0.008034f
C521 B.n481 VSUBS 0.008034f
C522 B.n482 VSUBS 0.008034f
C523 B.n483 VSUBS 0.008034f
C524 B.n484 VSUBS 0.008034f
C525 B.n485 VSUBS 0.008034f
C526 B.n486 VSUBS 0.008034f
C527 B.n487 VSUBS 0.008034f
C528 B.n488 VSUBS 0.008034f
C529 B.n489 VSUBS 0.008034f
C530 B.n490 VSUBS 0.008034f
C531 B.n491 VSUBS 0.008034f
C532 B.n492 VSUBS 0.008034f
C533 B.n493 VSUBS 0.008034f
C534 B.n494 VSUBS 0.008034f
C535 B.n495 VSUBS 0.008034f
C536 B.n496 VSUBS 0.008034f
C537 B.n497 VSUBS 0.008034f
C538 B.n498 VSUBS 0.008034f
C539 B.n499 VSUBS 0.008034f
C540 B.n500 VSUBS 0.008034f
C541 B.n501 VSUBS 0.008034f
C542 B.n502 VSUBS 0.008034f
C543 B.n503 VSUBS 0.008034f
C544 B.n504 VSUBS 0.008034f
C545 B.n505 VSUBS 0.008034f
C546 B.n506 VSUBS 0.008034f
C547 B.n507 VSUBS 0.008034f
C548 B.n508 VSUBS 0.008034f
C549 B.n509 VSUBS 0.008034f
C550 B.n510 VSUBS 0.008034f
C551 B.n511 VSUBS 0.008034f
C552 B.n512 VSUBS 0.008034f
C553 B.n513 VSUBS 0.008034f
C554 B.n514 VSUBS 0.008034f
C555 B.n515 VSUBS 0.008034f
C556 B.n516 VSUBS 0.008034f
C557 B.n517 VSUBS 0.008034f
C558 B.n518 VSUBS 0.008034f
C559 B.n519 VSUBS 0.008034f
C560 B.n520 VSUBS 0.008034f
C561 B.n521 VSUBS 0.008034f
C562 B.n522 VSUBS 0.008034f
C563 B.n523 VSUBS 0.008034f
C564 B.n524 VSUBS 0.008034f
C565 B.n525 VSUBS 0.008034f
C566 B.n526 VSUBS 0.008034f
C567 B.n527 VSUBS 0.008034f
C568 B.n528 VSUBS 0.008034f
C569 B.n529 VSUBS 0.008034f
C570 B.n530 VSUBS 0.008034f
C571 B.n531 VSUBS 0.008034f
C572 B.n532 VSUBS 0.008034f
C573 B.n533 VSUBS 0.008034f
C574 B.n534 VSUBS 0.008034f
C575 B.n535 VSUBS 0.008034f
C576 B.n536 VSUBS 0.008034f
C577 B.n537 VSUBS 0.008034f
C578 B.n538 VSUBS 0.008034f
C579 B.n539 VSUBS 0.008034f
C580 B.n540 VSUBS 0.008034f
C581 B.n541 VSUBS 0.008034f
C582 B.n542 VSUBS 0.008034f
C583 B.n543 VSUBS 0.008034f
C584 B.n544 VSUBS 0.008034f
C585 B.n545 VSUBS 0.008034f
C586 B.n546 VSUBS 0.008034f
C587 B.n547 VSUBS 0.008034f
C588 B.n548 VSUBS 0.008034f
C589 B.n549 VSUBS 0.008034f
C590 B.n550 VSUBS 0.008034f
C591 B.n551 VSUBS 0.008034f
C592 B.n552 VSUBS 0.008034f
C593 B.n553 VSUBS 0.008034f
C594 B.n554 VSUBS 0.008034f
C595 B.n555 VSUBS 0.008034f
C596 B.n556 VSUBS 0.008034f
C597 B.n557 VSUBS 0.008034f
C598 B.n558 VSUBS 0.008034f
C599 B.n559 VSUBS 0.008034f
C600 B.n560 VSUBS 0.008034f
C601 B.n561 VSUBS 0.008034f
C602 B.n562 VSUBS 0.008034f
C603 B.n563 VSUBS 0.008034f
C604 B.n564 VSUBS 0.008034f
C605 B.n565 VSUBS 0.008034f
C606 B.n566 VSUBS 0.008034f
C607 B.n567 VSUBS 0.008034f
C608 B.n568 VSUBS 0.008034f
C609 B.n569 VSUBS 0.008034f
C610 B.n570 VSUBS 0.008034f
C611 B.n571 VSUBS 0.008034f
C612 B.n572 VSUBS 0.008034f
C613 B.n573 VSUBS 0.008034f
C614 B.n574 VSUBS 0.008034f
C615 B.n575 VSUBS 0.008034f
C616 B.n576 VSUBS 0.008034f
C617 B.n577 VSUBS 0.008034f
C618 B.n578 VSUBS 0.008034f
C619 B.n579 VSUBS 0.008034f
C620 B.n580 VSUBS 0.008034f
C621 B.n581 VSUBS 0.008034f
C622 B.n582 VSUBS 0.008034f
C623 B.n583 VSUBS 0.008034f
C624 B.n584 VSUBS 0.008034f
C625 B.n585 VSUBS 0.008034f
C626 B.n586 VSUBS 0.008034f
C627 B.n587 VSUBS 0.008034f
C628 B.n588 VSUBS 0.008034f
C629 B.n589 VSUBS 0.008034f
C630 B.n590 VSUBS 0.008034f
C631 B.n591 VSUBS 0.008034f
C632 B.n592 VSUBS 0.008034f
C633 B.n593 VSUBS 0.008034f
C634 B.n594 VSUBS 0.008034f
C635 B.n595 VSUBS 0.019761f
C636 B.n596 VSUBS 0.018829f
C637 B.n597 VSUBS 0.019215f
C638 B.n598 VSUBS 0.008034f
C639 B.n599 VSUBS 0.008034f
C640 B.n600 VSUBS 0.008034f
C641 B.n601 VSUBS 0.008034f
C642 B.n602 VSUBS 0.008034f
C643 B.n603 VSUBS 0.008034f
C644 B.n604 VSUBS 0.008034f
C645 B.n605 VSUBS 0.008034f
C646 B.n606 VSUBS 0.008034f
C647 B.n607 VSUBS 0.008034f
C648 B.n608 VSUBS 0.008034f
C649 B.n609 VSUBS 0.008034f
C650 B.n610 VSUBS 0.008034f
C651 B.n611 VSUBS 0.008034f
C652 B.n612 VSUBS 0.008034f
C653 B.n613 VSUBS 0.008034f
C654 B.n614 VSUBS 0.008034f
C655 B.n615 VSUBS 0.008034f
C656 B.n616 VSUBS 0.008034f
C657 B.n617 VSUBS 0.008034f
C658 B.n618 VSUBS 0.008034f
C659 B.n619 VSUBS 0.008034f
C660 B.n620 VSUBS 0.008034f
C661 B.n621 VSUBS 0.008034f
C662 B.n622 VSUBS 0.008034f
C663 B.n623 VSUBS 0.008034f
C664 B.n624 VSUBS 0.008034f
C665 B.n625 VSUBS 0.008034f
C666 B.n626 VSUBS 0.008034f
C667 B.n627 VSUBS 0.008034f
C668 B.n628 VSUBS 0.008034f
C669 B.n629 VSUBS 0.008034f
C670 B.n630 VSUBS 0.008034f
C671 B.n631 VSUBS 0.008034f
C672 B.n632 VSUBS 0.008034f
C673 B.n633 VSUBS 0.008034f
C674 B.n634 VSUBS 0.008034f
C675 B.n635 VSUBS 0.008034f
C676 B.n636 VSUBS 0.008034f
C677 B.n637 VSUBS 0.008034f
C678 B.n638 VSUBS 0.008034f
C679 B.n639 VSUBS 0.008034f
C680 B.n640 VSUBS 0.008034f
C681 B.n641 VSUBS 0.008034f
C682 B.n642 VSUBS 0.008034f
C683 B.n643 VSUBS 0.008034f
C684 B.n644 VSUBS 0.008034f
C685 B.n645 VSUBS 0.008034f
C686 B.n646 VSUBS 0.008034f
C687 B.n647 VSUBS 0.008034f
C688 B.n648 VSUBS 0.008034f
C689 B.n649 VSUBS 0.008034f
C690 B.n650 VSUBS 0.008034f
C691 B.n651 VSUBS 0.008034f
C692 B.n652 VSUBS 0.008034f
C693 B.n653 VSUBS 0.008034f
C694 B.n654 VSUBS 0.008034f
C695 B.n655 VSUBS 0.008034f
C696 B.n656 VSUBS 0.008034f
C697 B.n657 VSUBS 0.008034f
C698 B.n658 VSUBS 0.008034f
C699 B.n659 VSUBS 0.008034f
C700 B.n660 VSUBS 0.008034f
C701 B.n661 VSUBS 0.008034f
C702 B.n662 VSUBS 0.008034f
C703 B.n663 VSUBS 0.008034f
C704 B.n664 VSUBS 0.008034f
C705 B.n665 VSUBS 0.008034f
C706 B.n666 VSUBS 0.008034f
C707 B.n667 VSUBS 0.008034f
C708 B.n668 VSUBS 0.008034f
C709 B.n669 VSUBS 0.008034f
C710 B.n670 VSUBS 0.008034f
C711 B.n671 VSUBS 0.005553f
C712 B.n672 VSUBS 0.018614f
C713 B.n673 VSUBS 0.006498f
C714 B.n674 VSUBS 0.008034f
C715 B.n675 VSUBS 0.008034f
C716 B.n676 VSUBS 0.008034f
C717 B.n677 VSUBS 0.008034f
C718 B.n678 VSUBS 0.008034f
C719 B.n679 VSUBS 0.008034f
C720 B.n680 VSUBS 0.008034f
C721 B.n681 VSUBS 0.008034f
C722 B.n682 VSUBS 0.008034f
C723 B.n683 VSUBS 0.008034f
C724 B.n684 VSUBS 0.008034f
C725 B.n685 VSUBS 0.006498f
C726 B.n686 VSUBS 0.018614f
C727 B.n687 VSUBS 0.005553f
C728 B.n688 VSUBS 0.008034f
C729 B.n689 VSUBS 0.008034f
C730 B.n690 VSUBS 0.008034f
C731 B.n691 VSUBS 0.008034f
C732 B.n692 VSUBS 0.008034f
C733 B.n693 VSUBS 0.008034f
C734 B.n694 VSUBS 0.008034f
C735 B.n695 VSUBS 0.008034f
C736 B.n696 VSUBS 0.008034f
C737 B.n697 VSUBS 0.008034f
C738 B.n698 VSUBS 0.008034f
C739 B.n699 VSUBS 0.008034f
C740 B.n700 VSUBS 0.008034f
C741 B.n701 VSUBS 0.008034f
C742 B.n702 VSUBS 0.008034f
C743 B.n703 VSUBS 0.008034f
C744 B.n704 VSUBS 0.008034f
C745 B.n705 VSUBS 0.008034f
C746 B.n706 VSUBS 0.008034f
C747 B.n707 VSUBS 0.008034f
C748 B.n708 VSUBS 0.008034f
C749 B.n709 VSUBS 0.008034f
C750 B.n710 VSUBS 0.008034f
C751 B.n711 VSUBS 0.008034f
C752 B.n712 VSUBS 0.008034f
C753 B.n713 VSUBS 0.008034f
C754 B.n714 VSUBS 0.008034f
C755 B.n715 VSUBS 0.008034f
C756 B.n716 VSUBS 0.008034f
C757 B.n717 VSUBS 0.008034f
C758 B.n718 VSUBS 0.008034f
C759 B.n719 VSUBS 0.008034f
C760 B.n720 VSUBS 0.008034f
C761 B.n721 VSUBS 0.008034f
C762 B.n722 VSUBS 0.008034f
C763 B.n723 VSUBS 0.008034f
C764 B.n724 VSUBS 0.008034f
C765 B.n725 VSUBS 0.008034f
C766 B.n726 VSUBS 0.008034f
C767 B.n727 VSUBS 0.008034f
C768 B.n728 VSUBS 0.008034f
C769 B.n729 VSUBS 0.008034f
C770 B.n730 VSUBS 0.008034f
C771 B.n731 VSUBS 0.008034f
C772 B.n732 VSUBS 0.008034f
C773 B.n733 VSUBS 0.008034f
C774 B.n734 VSUBS 0.008034f
C775 B.n735 VSUBS 0.008034f
C776 B.n736 VSUBS 0.008034f
C777 B.n737 VSUBS 0.008034f
C778 B.n738 VSUBS 0.008034f
C779 B.n739 VSUBS 0.008034f
C780 B.n740 VSUBS 0.008034f
C781 B.n741 VSUBS 0.008034f
C782 B.n742 VSUBS 0.008034f
C783 B.n743 VSUBS 0.008034f
C784 B.n744 VSUBS 0.008034f
C785 B.n745 VSUBS 0.008034f
C786 B.n746 VSUBS 0.008034f
C787 B.n747 VSUBS 0.008034f
C788 B.n748 VSUBS 0.008034f
C789 B.n749 VSUBS 0.008034f
C790 B.n750 VSUBS 0.008034f
C791 B.n751 VSUBS 0.008034f
C792 B.n752 VSUBS 0.008034f
C793 B.n753 VSUBS 0.008034f
C794 B.n754 VSUBS 0.008034f
C795 B.n755 VSUBS 0.008034f
C796 B.n756 VSUBS 0.008034f
C797 B.n757 VSUBS 0.008034f
C798 B.n758 VSUBS 0.008034f
C799 B.n759 VSUBS 0.008034f
C800 B.n760 VSUBS 0.008034f
C801 B.n761 VSUBS 0.019215f
C802 B.n762 VSUBS 0.018829f
C803 B.n763 VSUBS 0.018829f
C804 B.n764 VSUBS 0.008034f
C805 B.n765 VSUBS 0.008034f
C806 B.n766 VSUBS 0.008034f
C807 B.n767 VSUBS 0.008034f
C808 B.n768 VSUBS 0.008034f
C809 B.n769 VSUBS 0.008034f
C810 B.n770 VSUBS 0.008034f
C811 B.n771 VSUBS 0.008034f
C812 B.n772 VSUBS 0.008034f
C813 B.n773 VSUBS 0.008034f
C814 B.n774 VSUBS 0.008034f
C815 B.n775 VSUBS 0.008034f
C816 B.n776 VSUBS 0.008034f
C817 B.n777 VSUBS 0.008034f
C818 B.n778 VSUBS 0.008034f
C819 B.n779 VSUBS 0.008034f
C820 B.n780 VSUBS 0.008034f
C821 B.n781 VSUBS 0.008034f
C822 B.n782 VSUBS 0.008034f
C823 B.n783 VSUBS 0.008034f
C824 B.n784 VSUBS 0.008034f
C825 B.n785 VSUBS 0.008034f
C826 B.n786 VSUBS 0.008034f
C827 B.n787 VSUBS 0.008034f
C828 B.n788 VSUBS 0.008034f
C829 B.n789 VSUBS 0.008034f
C830 B.n790 VSUBS 0.008034f
C831 B.n791 VSUBS 0.008034f
C832 B.n792 VSUBS 0.008034f
C833 B.n793 VSUBS 0.008034f
C834 B.n794 VSUBS 0.008034f
C835 B.n795 VSUBS 0.008034f
C836 B.n796 VSUBS 0.008034f
C837 B.n797 VSUBS 0.008034f
C838 B.n798 VSUBS 0.008034f
C839 B.n799 VSUBS 0.008034f
C840 B.n800 VSUBS 0.008034f
C841 B.n801 VSUBS 0.008034f
C842 B.n802 VSUBS 0.008034f
C843 B.n803 VSUBS 0.008034f
C844 B.n804 VSUBS 0.008034f
C845 B.n805 VSUBS 0.008034f
C846 B.n806 VSUBS 0.008034f
C847 B.n807 VSUBS 0.008034f
C848 B.n808 VSUBS 0.008034f
C849 B.n809 VSUBS 0.008034f
C850 B.n810 VSUBS 0.008034f
C851 B.n811 VSUBS 0.008034f
C852 B.n812 VSUBS 0.008034f
C853 B.n813 VSUBS 0.008034f
C854 B.n814 VSUBS 0.008034f
C855 B.n815 VSUBS 0.008034f
C856 B.n816 VSUBS 0.008034f
C857 B.n817 VSUBS 0.008034f
C858 B.n818 VSUBS 0.008034f
C859 B.n819 VSUBS 0.008034f
C860 B.n820 VSUBS 0.008034f
C861 B.n821 VSUBS 0.008034f
C862 B.n822 VSUBS 0.008034f
C863 B.n823 VSUBS 0.008034f
C864 B.n824 VSUBS 0.008034f
C865 B.n825 VSUBS 0.008034f
C866 B.n826 VSUBS 0.008034f
C867 B.n827 VSUBS 0.008034f
C868 B.n828 VSUBS 0.008034f
C869 B.n829 VSUBS 0.008034f
C870 B.n830 VSUBS 0.008034f
C871 B.n831 VSUBS 0.008034f
C872 B.n832 VSUBS 0.008034f
C873 B.n833 VSUBS 0.008034f
C874 B.n834 VSUBS 0.008034f
C875 B.n835 VSUBS 0.018192f
C876 VDD2.n0 VSUBS 0.029977f
C877 VDD2.n1 VSUBS 0.0276f
C878 VDD2.n2 VSUBS 0.014831f
C879 VDD2.n3 VSUBS 0.035055f
C880 VDD2.n4 VSUBS 0.015704f
C881 VDD2.n5 VSUBS 0.0276f
C882 VDD2.n6 VSUBS 0.014831f
C883 VDD2.n7 VSUBS 0.035055f
C884 VDD2.n8 VSUBS 0.015704f
C885 VDD2.n9 VSUBS 0.0276f
C886 VDD2.n10 VSUBS 0.014831f
C887 VDD2.n11 VSUBS 0.035055f
C888 VDD2.n12 VSUBS 0.015704f
C889 VDD2.n13 VSUBS 0.0276f
C890 VDD2.n14 VSUBS 0.014831f
C891 VDD2.n15 VSUBS 0.035055f
C892 VDD2.n16 VSUBS 0.015704f
C893 VDD2.n17 VSUBS 0.0276f
C894 VDD2.n18 VSUBS 0.014831f
C895 VDD2.n19 VSUBS 0.035055f
C896 VDD2.n20 VSUBS 0.015704f
C897 VDD2.n21 VSUBS 0.0276f
C898 VDD2.n22 VSUBS 0.014831f
C899 VDD2.n23 VSUBS 0.035055f
C900 VDD2.n24 VSUBS 0.015704f
C901 VDD2.n25 VSUBS 0.193092f
C902 VDD2.t4 VSUBS 0.075035f
C903 VDD2.n26 VSUBS 0.026292f
C904 VDD2.n27 VSUBS 0.022301f
C905 VDD2.n28 VSUBS 0.014831f
C906 VDD2.n29 VSUBS 1.73977f
C907 VDD2.n30 VSUBS 0.0276f
C908 VDD2.n31 VSUBS 0.014831f
C909 VDD2.n32 VSUBS 0.015704f
C910 VDD2.n33 VSUBS 0.035055f
C911 VDD2.n34 VSUBS 0.035055f
C912 VDD2.n35 VSUBS 0.015704f
C913 VDD2.n36 VSUBS 0.014831f
C914 VDD2.n37 VSUBS 0.0276f
C915 VDD2.n38 VSUBS 0.0276f
C916 VDD2.n39 VSUBS 0.014831f
C917 VDD2.n40 VSUBS 0.015704f
C918 VDD2.n41 VSUBS 0.035055f
C919 VDD2.n42 VSUBS 0.035055f
C920 VDD2.n43 VSUBS 0.015704f
C921 VDD2.n44 VSUBS 0.014831f
C922 VDD2.n45 VSUBS 0.0276f
C923 VDD2.n46 VSUBS 0.0276f
C924 VDD2.n47 VSUBS 0.014831f
C925 VDD2.n48 VSUBS 0.015704f
C926 VDD2.n49 VSUBS 0.035055f
C927 VDD2.n50 VSUBS 0.035055f
C928 VDD2.n51 VSUBS 0.015704f
C929 VDD2.n52 VSUBS 0.014831f
C930 VDD2.n53 VSUBS 0.0276f
C931 VDD2.n54 VSUBS 0.0276f
C932 VDD2.n55 VSUBS 0.014831f
C933 VDD2.n56 VSUBS 0.015704f
C934 VDD2.n57 VSUBS 0.035055f
C935 VDD2.n58 VSUBS 0.035055f
C936 VDD2.n59 VSUBS 0.015704f
C937 VDD2.n60 VSUBS 0.014831f
C938 VDD2.n61 VSUBS 0.0276f
C939 VDD2.n62 VSUBS 0.0276f
C940 VDD2.n63 VSUBS 0.014831f
C941 VDD2.n64 VSUBS 0.015704f
C942 VDD2.n65 VSUBS 0.035055f
C943 VDD2.n66 VSUBS 0.035055f
C944 VDD2.n67 VSUBS 0.035055f
C945 VDD2.n68 VSUBS 0.015704f
C946 VDD2.n69 VSUBS 0.014831f
C947 VDD2.n70 VSUBS 0.0276f
C948 VDD2.n71 VSUBS 0.0276f
C949 VDD2.n72 VSUBS 0.014831f
C950 VDD2.n73 VSUBS 0.015267f
C951 VDD2.n74 VSUBS 0.015267f
C952 VDD2.n75 VSUBS 0.035055f
C953 VDD2.n76 VSUBS 0.083675f
C954 VDD2.n77 VSUBS 0.015704f
C955 VDD2.n78 VSUBS 0.014831f
C956 VDD2.n79 VSUBS 0.070583f
C957 VDD2.n80 VSUBS 0.070883f
C958 VDD2.t1 VSUBS 0.323232f
C959 VDD2.t2 VSUBS 0.323232f
C960 VDD2.n81 VSUBS 2.63998f
C961 VDD2.n82 VSUBS 3.65369f
C962 VDD2.n83 VSUBS 0.029977f
C963 VDD2.n84 VSUBS 0.0276f
C964 VDD2.n85 VSUBS 0.014831f
C965 VDD2.n86 VSUBS 0.035055f
C966 VDD2.n87 VSUBS 0.015704f
C967 VDD2.n88 VSUBS 0.0276f
C968 VDD2.n89 VSUBS 0.014831f
C969 VDD2.n90 VSUBS 0.035055f
C970 VDD2.n91 VSUBS 0.035055f
C971 VDD2.n92 VSUBS 0.015704f
C972 VDD2.n93 VSUBS 0.0276f
C973 VDD2.n94 VSUBS 0.014831f
C974 VDD2.n95 VSUBS 0.035055f
C975 VDD2.n96 VSUBS 0.015704f
C976 VDD2.n97 VSUBS 0.0276f
C977 VDD2.n98 VSUBS 0.014831f
C978 VDD2.n99 VSUBS 0.035055f
C979 VDD2.n100 VSUBS 0.015704f
C980 VDD2.n101 VSUBS 0.0276f
C981 VDD2.n102 VSUBS 0.014831f
C982 VDD2.n103 VSUBS 0.035055f
C983 VDD2.n104 VSUBS 0.015704f
C984 VDD2.n105 VSUBS 0.0276f
C985 VDD2.n106 VSUBS 0.014831f
C986 VDD2.n107 VSUBS 0.035055f
C987 VDD2.n108 VSUBS 0.015704f
C988 VDD2.n109 VSUBS 0.193092f
C989 VDD2.t0 VSUBS 0.075035f
C990 VDD2.n110 VSUBS 0.026292f
C991 VDD2.n111 VSUBS 0.022301f
C992 VDD2.n112 VSUBS 0.014831f
C993 VDD2.n113 VSUBS 1.73977f
C994 VDD2.n114 VSUBS 0.0276f
C995 VDD2.n115 VSUBS 0.014831f
C996 VDD2.n116 VSUBS 0.015704f
C997 VDD2.n117 VSUBS 0.035055f
C998 VDD2.n118 VSUBS 0.035055f
C999 VDD2.n119 VSUBS 0.015704f
C1000 VDD2.n120 VSUBS 0.014831f
C1001 VDD2.n121 VSUBS 0.0276f
C1002 VDD2.n122 VSUBS 0.0276f
C1003 VDD2.n123 VSUBS 0.014831f
C1004 VDD2.n124 VSUBS 0.015704f
C1005 VDD2.n125 VSUBS 0.035055f
C1006 VDD2.n126 VSUBS 0.035055f
C1007 VDD2.n127 VSUBS 0.015704f
C1008 VDD2.n128 VSUBS 0.014831f
C1009 VDD2.n129 VSUBS 0.0276f
C1010 VDD2.n130 VSUBS 0.0276f
C1011 VDD2.n131 VSUBS 0.014831f
C1012 VDD2.n132 VSUBS 0.015704f
C1013 VDD2.n133 VSUBS 0.035055f
C1014 VDD2.n134 VSUBS 0.035055f
C1015 VDD2.n135 VSUBS 0.015704f
C1016 VDD2.n136 VSUBS 0.014831f
C1017 VDD2.n137 VSUBS 0.0276f
C1018 VDD2.n138 VSUBS 0.0276f
C1019 VDD2.n139 VSUBS 0.014831f
C1020 VDD2.n140 VSUBS 0.015704f
C1021 VDD2.n141 VSUBS 0.035055f
C1022 VDD2.n142 VSUBS 0.035055f
C1023 VDD2.n143 VSUBS 0.015704f
C1024 VDD2.n144 VSUBS 0.014831f
C1025 VDD2.n145 VSUBS 0.0276f
C1026 VDD2.n146 VSUBS 0.0276f
C1027 VDD2.n147 VSUBS 0.014831f
C1028 VDD2.n148 VSUBS 0.015704f
C1029 VDD2.n149 VSUBS 0.035055f
C1030 VDD2.n150 VSUBS 0.035055f
C1031 VDD2.n151 VSUBS 0.015704f
C1032 VDD2.n152 VSUBS 0.014831f
C1033 VDD2.n153 VSUBS 0.0276f
C1034 VDD2.n154 VSUBS 0.0276f
C1035 VDD2.n155 VSUBS 0.014831f
C1036 VDD2.n156 VSUBS 0.015267f
C1037 VDD2.n157 VSUBS 0.015267f
C1038 VDD2.n158 VSUBS 0.035055f
C1039 VDD2.n159 VSUBS 0.083675f
C1040 VDD2.n160 VSUBS 0.015704f
C1041 VDD2.n161 VSUBS 0.014831f
C1042 VDD2.n162 VSUBS 0.070583f
C1043 VDD2.n163 VSUBS 0.061236f
C1044 VDD2.n164 VSUBS 3.20603f
C1045 VDD2.t5 VSUBS 0.323232f
C1046 VDD2.t3 VSUBS 0.323232f
C1047 VDD2.n165 VSUBS 2.63994f
C1048 VN.t3 VSUBS 3.24675f
C1049 VN.n0 VSUBS 1.2331f
C1050 VN.n1 VSUBS 0.02622f
C1051 VN.n2 VSUBS 0.033763f
C1052 VN.n3 VSUBS 0.298194f
C1053 VN.t4 VSUBS 3.24675f
C1054 VN.t1 VSUBS 3.53839f
C1055 VN.n4 VSUBS 1.16961f
C1056 VN.n5 VSUBS 1.22839f
C1057 VN.n6 VSUBS 0.048623f
C1058 VN.n7 VSUBS 0.048623f
C1059 VN.n8 VSUBS 0.02622f
C1060 VN.n9 VSUBS 0.02622f
C1061 VN.n10 VSUBS 0.02622f
C1062 VN.n11 VSUBS 0.042468f
C1063 VN.n12 VSUBS 0.048623f
C1064 VN.n13 VSUBS 0.042862f
C1065 VN.n14 VSUBS 0.042312f
C1066 VN.n15 VSUBS 0.056606f
C1067 VN.t5 VSUBS 3.24675f
C1068 VN.n16 VSUBS 1.2331f
C1069 VN.n17 VSUBS 0.02622f
C1070 VN.n18 VSUBS 0.033763f
C1071 VN.n19 VSUBS 0.298194f
C1072 VN.t0 VSUBS 3.24675f
C1073 VN.t2 VSUBS 3.53839f
C1074 VN.n20 VSUBS 1.16961f
C1075 VN.n21 VSUBS 1.22839f
C1076 VN.n22 VSUBS 0.048623f
C1077 VN.n23 VSUBS 0.048623f
C1078 VN.n24 VSUBS 0.02622f
C1079 VN.n25 VSUBS 0.02622f
C1080 VN.n26 VSUBS 0.02622f
C1081 VN.n27 VSUBS 0.042468f
C1082 VN.n28 VSUBS 0.048623f
C1083 VN.n29 VSUBS 0.042862f
C1084 VN.n30 VSUBS 0.042312f
C1085 VN.n31 VSUBS 1.6098f
C1086 VTAIL.t4 VSUBS 0.334677f
C1087 VTAIL.t0 VSUBS 0.334677f
C1088 VTAIL.n0 VSUBS 2.57318f
C1089 VTAIL.n1 VSUBS 0.895047f
C1090 VTAIL.n2 VSUBS 0.031039f
C1091 VTAIL.n3 VSUBS 0.028577f
C1092 VTAIL.n4 VSUBS 0.015356f
C1093 VTAIL.n5 VSUBS 0.036297f
C1094 VTAIL.n6 VSUBS 0.01626f
C1095 VTAIL.n7 VSUBS 0.028577f
C1096 VTAIL.n8 VSUBS 0.015356f
C1097 VTAIL.n9 VSUBS 0.036297f
C1098 VTAIL.n10 VSUBS 0.01626f
C1099 VTAIL.n11 VSUBS 0.028577f
C1100 VTAIL.n12 VSUBS 0.015356f
C1101 VTAIL.n13 VSUBS 0.036297f
C1102 VTAIL.n14 VSUBS 0.01626f
C1103 VTAIL.n15 VSUBS 0.028577f
C1104 VTAIL.n16 VSUBS 0.015356f
C1105 VTAIL.n17 VSUBS 0.036297f
C1106 VTAIL.n18 VSUBS 0.01626f
C1107 VTAIL.n19 VSUBS 0.028577f
C1108 VTAIL.n20 VSUBS 0.015356f
C1109 VTAIL.n21 VSUBS 0.036297f
C1110 VTAIL.n22 VSUBS 0.01626f
C1111 VTAIL.n23 VSUBS 0.028577f
C1112 VTAIL.n24 VSUBS 0.015356f
C1113 VTAIL.n25 VSUBS 0.036297f
C1114 VTAIL.n26 VSUBS 0.01626f
C1115 VTAIL.n27 VSUBS 0.19993f
C1116 VTAIL.t7 VSUBS 0.077691f
C1117 VTAIL.n28 VSUBS 0.027222f
C1118 VTAIL.n29 VSUBS 0.02309f
C1119 VTAIL.n30 VSUBS 0.015356f
C1120 VTAIL.n31 VSUBS 1.80138f
C1121 VTAIL.n32 VSUBS 0.028577f
C1122 VTAIL.n33 VSUBS 0.015356f
C1123 VTAIL.n34 VSUBS 0.01626f
C1124 VTAIL.n35 VSUBS 0.036297f
C1125 VTAIL.n36 VSUBS 0.036297f
C1126 VTAIL.n37 VSUBS 0.01626f
C1127 VTAIL.n38 VSUBS 0.015356f
C1128 VTAIL.n39 VSUBS 0.028577f
C1129 VTAIL.n40 VSUBS 0.028577f
C1130 VTAIL.n41 VSUBS 0.015356f
C1131 VTAIL.n42 VSUBS 0.01626f
C1132 VTAIL.n43 VSUBS 0.036297f
C1133 VTAIL.n44 VSUBS 0.036297f
C1134 VTAIL.n45 VSUBS 0.01626f
C1135 VTAIL.n46 VSUBS 0.015356f
C1136 VTAIL.n47 VSUBS 0.028577f
C1137 VTAIL.n48 VSUBS 0.028577f
C1138 VTAIL.n49 VSUBS 0.015356f
C1139 VTAIL.n50 VSUBS 0.01626f
C1140 VTAIL.n51 VSUBS 0.036297f
C1141 VTAIL.n52 VSUBS 0.036297f
C1142 VTAIL.n53 VSUBS 0.01626f
C1143 VTAIL.n54 VSUBS 0.015356f
C1144 VTAIL.n55 VSUBS 0.028577f
C1145 VTAIL.n56 VSUBS 0.028577f
C1146 VTAIL.n57 VSUBS 0.015356f
C1147 VTAIL.n58 VSUBS 0.01626f
C1148 VTAIL.n59 VSUBS 0.036297f
C1149 VTAIL.n60 VSUBS 0.036297f
C1150 VTAIL.n61 VSUBS 0.01626f
C1151 VTAIL.n62 VSUBS 0.015356f
C1152 VTAIL.n63 VSUBS 0.028577f
C1153 VTAIL.n64 VSUBS 0.028577f
C1154 VTAIL.n65 VSUBS 0.015356f
C1155 VTAIL.n66 VSUBS 0.01626f
C1156 VTAIL.n67 VSUBS 0.036297f
C1157 VTAIL.n68 VSUBS 0.036297f
C1158 VTAIL.n69 VSUBS 0.036297f
C1159 VTAIL.n70 VSUBS 0.01626f
C1160 VTAIL.n71 VSUBS 0.015356f
C1161 VTAIL.n72 VSUBS 0.028577f
C1162 VTAIL.n73 VSUBS 0.028577f
C1163 VTAIL.n74 VSUBS 0.015356f
C1164 VTAIL.n75 VSUBS 0.015808f
C1165 VTAIL.n76 VSUBS 0.015808f
C1166 VTAIL.n77 VSUBS 0.036297f
C1167 VTAIL.n78 VSUBS 0.086638f
C1168 VTAIL.n79 VSUBS 0.01626f
C1169 VTAIL.n80 VSUBS 0.015356f
C1170 VTAIL.n81 VSUBS 0.073083f
C1171 VTAIL.n82 VSUBS 0.043721f
C1172 VTAIL.n83 VSUBS 0.474112f
C1173 VTAIL.t8 VSUBS 0.334677f
C1174 VTAIL.t11 VSUBS 0.334677f
C1175 VTAIL.n84 VSUBS 2.57318f
C1176 VTAIL.n85 VSUBS 3.01476f
C1177 VTAIL.t1 VSUBS 0.334677f
C1178 VTAIL.t5 VSUBS 0.334677f
C1179 VTAIL.n86 VSUBS 2.5732f
C1180 VTAIL.n87 VSUBS 3.01474f
C1181 VTAIL.n88 VSUBS 0.031039f
C1182 VTAIL.n89 VSUBS 0.028577f
C1183 VTAIL.n90 VSUBS 0.015356f
C1184 VTAIL.n91 VSUBS 0.036297f
C1185 VTAIL.n92 VSUBS 0.01626f
C1186 VTAIL.n93 VSUBS 0.028577f
C1187 VTAIL.n94 VSUBS 0.015356f
C1188 VTAIL.n95 VSUBS 0.036297f
C1189 VTAIL.n96 VSUBS 0.036297f
C1190 VTAIL.n97 VSUBS 0.01626f
C1191 VTAIL.n98 VSUBS 0.028577f
C1192 VTAIL.n99 VSUBS 0.015356f
C1193 VTAIL.n100 VSUBS 0.036297f
C1194 VTAIL.n101 VSUBS 0.01626f
C1195 VTAIL.n102 VSUBS 0.028577f
C1196 VTAIL.n103 VSUBS 0.015356f
C1197 VTAIL.n104 VSUBS 0.036297f
C1198 VTAIL.n105 VSUBS 0.01626f
C1199 VTAIL.n106 VSUBS 0.028577f
C1200 VTAIL.n107 VSUBS 0.015356f
C1201 VTAIL.n108 VSUBS 0.036297f
C1202 VTAIL.n109 VSUBS 0.01626f
C1203 VTAIL.n110 VSUBS 0.028577f
C1204 VTAIL.n111 VSUBS 0.015356f
C1205 VTAIL.n112 VSUBS 0.036297f
C1206 VTAIL.n113 VSUBS 0.01626f
C1207 VTAIL.n114 VSUBS 0.19993f
C1208 VTAIL.t2 VSUBS 0.077691f
C1209 VTAIL.n115 VSUBS 0.027222f
C1210 VTAIL.n116 VSUBS 0.02309f
C1211 VTAIL.n117 VSUBS 0.015356f
C1212 VTAIL.n118 VSUBS 1.80138f
C1213 VTAIL.n119 VSUBS 0.028577f
C1214 VTAIL.n120 VSUBS 0.015356f
C1215 VTAIL.n121 VSUBS 0.01626f
C1216 VTAIL.n122 VSUBS 0.036297f
C1217 VTAIL.n123 VSUBS 0.036297f
C1218 VTAIL.n124 VSUBS 0.01626f
C1219 VTAIL.n125 VSUBS 0.015356f
C1220 VTAIL.n126 VSUBS 0.028577f
C1221 VTAIL.n127 VSUBS 0.028577f
C1222 VTAIL.n128 VSUBS 0.015356f
C1223 VTAIL.n129 VSUBS 0.01626f
C1224 VTAIL.n130 VSUBS 0.036297f
C1225 VTAIL.n131 VSUBS 0.036297f
C1226 VTAIL.n132 VSUBS 0.01626f
C1227 VTAIL.n133 VSUBS 0.015356f
C1228 VTAIL.n134 VSUBS 0.028577f
C1229 VTAIL.n135 VSUBS 0.028577f
C1230 VTAIL.n136 VSUBS 0.015356f
C1231 VTAIL.n137 VSUBS 0.01626f
C1232 VTAIL.n138 VSUBS 0.036297f
C1233 VTAIL.n139 VSUBS 0.036297f
C1234 VTAIL.n140 VSUBS 0.01626f
C1235 VTAIL.n141 VSUBS 0.015356f
C1236 VTAIL.n142 VSUBS 0.028577f
C1237 VTAIL.n143 VSUBS 0.028577f
C1238 VTAIL.n144 VSUBS 0.015356f
C1239 VTAIL.n145 VSUBS 0.01626f
C1240 VTAIL.n146 VSUBS 0.036297f
C1241 VTAIL.n147 VSUBS 0.036297f
C1242 VTAIL.n148 VSUBS 0.01626f
C1243 VTAIL.n149 VSUBS 0.015356f
C1244 VTAIL.n150 VSUBS 0.028577f
C1245 VTAIL.n151 VSUBS 0.028577f
C1246 VTAIL.n152 VSUBS 0.015356f
C1247 VTAIL.n153 VSUBS 0.01626f
C1248 VTAIL.n154 VSUBS 0.036297f
C1249 VTAIL.n155 VSUBS 0.036297f
C1250 VTAIL.n156 VSUBS 0.01626f
C1251 VTAIL.n157 VSUBS 0.015356f
C1252 VTAIL.n158 VSUBS 0.028577f
C1253 VTAIL.n159 VSUBS 0.028577f
C1254 VTAIL.n160 VSUBS 0.015356f
C1255 VTAIL.n161 VSUBS 0.015808f
C1256 VTAIL.n162 VSUBS 0.015808f
C1257 VTAIL.n163 VSUBS 0.036297f
C1258 VTAIL.n164 VSUBS 0.086638f
C1259 VTAIL.n165 VSUBS 0.01626f
C1260 VTAIL.n166 VSUBS 0.015356f
C1261 VTAIL.n167 VSUBS 0.073083f
C1262 VTAIL.n168 VSUBS 0.043721f
C1263 VTAIL.n169 VSUBS 0.474112f
C1264 VTAIL.t10 VSUBS 0.334677f
C1265 VTAIL.t6 VSUBS 0.334677f
C1266 VTAIL.n170 VSUBS 2.5732f
C1267 VTAIL.n171 VSUBS 1.09091f
C1268 VTAIL.n172 VSUBS 0.031039f
C1269 VTAIL.n173 VSUBS 0.028577f
C1270 VTAIL.n174 VSUBS 0.015356f
C1271 VTAIL.n175 VSUBS 0.036297f
C1272 VTAIL.n176 VSUBS 0.01626f
C1273 VTAIL.n177 VSUBS 0.028577f
C1274 VTAIL.n178 VSUBS 0.015356f
C1275 VTAIL.n179 VSUBS 0.036297f
C1276 VTAIL.n180 VSUBS 0.036297f
C1277 VTAIL.n181 VSUBS 0.01626f
C1278 VTAIL.n182 VSUBS 0.028577f
C1279 VTAIL.n183 VSUBS 0.015356f
C1280 VTAIL.n184 VSUBS 0.036297f
C1281 VTAIL.n185 VSUBS 0.01626f
C1282 VTAIL.n186 VSUBS 0.028577f
C1283 VTAIL.n187 VSUBS 0.015356f
C1284 VTAIL.n188 VSUBS 0.036297f
C1285 VTAIL.n189 VSUBS 0.01626f
C1286 VTAIL.n190 VSUBS 0.028577f
C1287 VTAIL.n191 VSUBS 0.015356f
C1288 VTAIL.n192 VSUBS 0.036297f
C1289 VTAIL.n193 VSUBS 0.01626f
C1290 VTAIL.n194 VSUBS 0.028577f
C1291 VTAIL.n195 VSUBS 0.015356f
C1292 VTAIL.n196 VSUBS 0.036297f
C1293 VTAIL.n197 VSUBS 0.01626f
C1294 VTAIL.n198 VSUBS 0.19993f
C1295 VTAIL.t9 VSUBS 0.077691f
C1296 VTAIL.n199 VSUBS 0.027222f
C1297 VTAIL.n200 VSUBS 0.02309f
C1298 VTAIL.n201 VSUBS 0.015356f
C1299 VTAIL.n202 VSUBS 1.80138f
C1300 VTAIL.n203 VSUBS 0.028577f
C1301 VTAIL.n204 VSUBS 0.015356f
C1302 VTAIL.n205 VSUBS 0.01626f
C1303 VTAIL.n206 VSUBS 0.036297f
C1304 VTAIL.n207 VSUBS 0.036297f
C1305 VTAIL.n208 VSUBS 0.01626f
C1306 VTAIL.n209 VSUBS 0.015356f
C1307 VTAIL.n210 VSUBS 0.028577f
C1308 VTAIL.n211 VSUBS 0.028577f
C1309 VTAIL.n212 VSUBS 0.015356f
C1310 VTAIL.n213 VSUBS 0.01626f
C1311 VTAIL.n214 VSUBS 0.036297f
C1312 VTAIL.n215 VSUBS 0.036297f
C1313 VTAIL.n216 VSUBS 0.01626f
C1314 VTAIL.n217 VSUBS 0.015356f
C1315 VTAIL.n218 VSUBS 0.028577f
C1316 VTAIL.n219 VSUBS 0.028577f
C1317 VTAIL.n220 VSUBS 0.015356f
C1318 VTAIL.n221 VSUBS 0.01626f
C1319 VTAIL.n222 VSUBS 0.036297f
C1320 VTAIL.n223 VSUBS 0.036297f
C1321 VTAIL.n224 VSUBS 0.01626f
C1322 VTAIL.n225 VSUBS 0.015356f
C1323 VTAIL.n226 VSUBS 0.028577f
C1324 VTAIL.n227 VSUBS 0.028577f
C1325 VTAIL.n228 VSUBS 0.015356f
C1326 VTAIL.n229 VSUBS 0.01626f
C1327 VTAIL.n230 VSUBS 0.036297f
C1328 VTAIL.n231 VSUBS 0.036297f
C1329 VTAIL.n232 VSUBS 0.01626f
C1330 VTAIL.n233 VSUBS 0.015356f
C1331 VTAIL.n234 VSUBS 0.028577f
C1332 VTAIL.n235 VSUBS 0.028577f
C1333 VTAIL.n236 VSUBS 0.015356f
C1334 VTAIL.n237 VSUBS 0.01626f
C1335 VTAIL.n238 VSUBS 0.036297f
C1336 VTAIL.n239 VSUBS 0.036297f
C1337 VTAIL.n240 VSUBS 0.01626f
C1338 VTAIL.n241 VSUBS 0.015356f
C1339 VTAIL.n242 VSUBS 0.028577f
C1340 VTAIL.n243 VSUBS 0.028577f
C1341 VTAIL.n244 VSUBS 0.015356f
C1342 VTAIL.n245 VSUBS 0.015808f
C1343 VTAIL.n246 VSUBS 0.015808f
C1344 VTAIL.n247 VSUBS 0.036297f
C1345 VTAIL.n248 VSUBS 0.086638f
C1346 VTAIL.n249 VSUBS 0.01626f
C1347 VTAIL.n250 VSUBS 0.015356f
C1348 VTAIL.n251 VSUBS 0.073083f
C1349 VTAIL.n252 VSUBS 0.043721f
C1350 VTAIL.n253 VSUBS 2.12964f
C1351 VTAIL.n254 VSUBS 0.031039f
C1352 VTAIL.n255 VSUBS 0.028577f
C1353 VTAIL.n256 VSUBS 0.015356f
C1354 VTAIL.n257 VSUBS 0.036297f
C1355 VTAIL.n258 VSUBS 0.01626f
C1356 VTAIL.n259 VSUBS 0.028577f
C1357 VTAIL.n260 VSUBS 0.015356f
C1358 VTAIL.n261 VSUBS 0.036297f
C1359 VTAIL.n262 VSUBS 0.01626f
C1360 VTAIL.n263 VSUBS 0.028577f
C1361 VTAIL.n264 VSUBS 0.015356f
C1362 VTAIL.n265 VSUBS 0.036297f
C1363 VTAIL.n266 VSUBS 0.01626f
C1364 VTAIL.n267 VSUBS 0.028577f
C1365 VTAIL.n268 VSUBS 0.015356f
C1366 VTAIL.n269 VSUBS 0.036297f
C1367 VTAIL.n270 VSUBS 0.01626f
C1368 VTAIL.n271 VSUBS 0.028577f
C1369 VTAIL.n272 VSUBS 0.015356f
C1370 VTAIL.n273 VSUBS 0.036297f
C1371 VTAIL.n274 VSUBS 0.01626f
C1372 VTAIL.n275 VSUBS 0.028577f
C1373 VTAIL.n276 VSUBS 0.015356f
C1374 VTAIL.n277 VSUBS 0.036297f
C1375 VTAIL.n278 VSUBS 0.01626f
C1376 VTAIL.n279 VSUBS 0.19993f
C1377 VTAIL.t3 VSUBS 0.077691f
C1378 VTAIL.n280 VSUBS 0.027222f
C1379 VTAIL.n281 VSUBS 0.02309f
C1380 VTAIL.n282 VSUBS 0.015356f
C1381 VTAIL.n283 VSUBS 1.80138f
C1382 VTAIL.n284 VSUBS 0.028577f
C1383 VTAIL.n285 VSUBS 0.015356f
C1384 VTAIL.n286 VSUBS 0.01626f
C1385 VTAIL.n287 VSUBS 0.036297f
C1386 VTAIL.n288 VSUBS 0.036297f
C1387 VTAIL.n289 VSUBS 0.01626f
C1388 VTAIL.n290 VSUBS 0.015356f
C1389 VTAIL.n291 VSUBS 0.028577f
C1390 VTAIL.n292 VSUBS 0.028577f
C1391 VTAIL.n293 VSUBS 0.015356f
C1392 VTAIL.n294 VSUBS 0.01626f
C1393 VTAIL.n295 VSUBS 0.036297f
C1394 VTAIL.n296 VSUBS 0.036297f
C1395 VTAIL.n297 VSUBS 0.01626f
C1396 VTAIL.n298 VSUBS 0.015356f
C1397 VTAIL.n299 VSUBS 0.028577f
C1398 VTAIL.n300 VSUBS 0.028577f
C1399 VTAIL.n301 VSUBS 0.015356f
C1400 VTAIL.n302 VSUBS 0.01626f
C1401 VTAIL.n303 VSUBS 0.036297f
C1402 VTAIL.n304 VSUBS 0.036297f
C1403 VTAIL.n305 VSUBS 0.01626f
C1404 VTAIL.n306 VSUBS 0.015356f
C1405 VTAIL.n307 VSUBS 0.028577f
C1406 VTAIL.n308 VSUBS 0.028577f
C1407 VTAIL.n309 VSUBS 0.015356f
C1408 VTAIL.n310 VSUBS 0.01626f
C1409 VTAIL.n311 VSUBS 0.036297f
C1410 VTAIL.n312 VSUBS 0.036297f
C1411 VTAIL.n313 VSUBS 0.01626f
C1412 VTAIL.n314 VSUBS 0.015356f
C1413 VTAIL.n315 VSUBS 0.028577f
C1414 VTAIL.n316 VSUBS 0.028577f
C1415 VTAIL.n317 VSUBS 0.015356f
C1416 VTAIL.n318 VSUBS 0.01626f
C1417 VTAIL.n319 VSUBS 0.036297f
C1418 VTAIL.n320 VSUBS 0.036297f
C1419 VTAIL.n321 VSUBS 0.036297f
C1420 VTAIL.n322 VSUBS 0.01626f
C1421 VTAIL.n323 VSUBS 0.015356f
C1422 VTAIL.n324 VSUBS 0.028577f
C1423 VTAIL.n325 VSUBS 0.028577f
C1424 VTAIL.n326 VSUBS 0.015356f
C1425 VTAIL.n327 VSUBS 0.015808f
C1426 VTAIL.n328 VSUBS 0.015808f
C1427 VTAIL.n329 VSUBS 0.036297f
C1428 VTAIL.n330 VSUBS 0.086638f
C1429 VTAIL.n331 VSUBS 0.01626f
C1430 VTAIL.n332 VSUBS 0.015356f
C1431 VTAIL.n333 VSUBS 0.073083f
C1432 VTAIL.n334 VSUBS 0.043721f
C1433 VTAIL.n335 VSUBS 2.0572f
C1434 VDD1.n0 VSUBS 0.029975f
C1435 VDD1.n1 VSUBS 0.027598f
C1436 VDD1.n2 VSUBS 0.01483f
C1437 VDD1.n3 VSUBS 0.035052f
C1438 VDD1.n4 VSUBS 0.015702f
C1439 VDD1.n5 VSUBS 0.027598f
C1440 VDD1.n6 VSUBS 0.01483f
C1441 VDD1.n7 VSUBS 0.035052f
C1442 VDD1.n8 VSUBS 0.035052f
C1443 VDD1.n9 VSUBS 0.015702f
C1444 VDD1.n10 VSUBS 0.027598f
C1445 VDD1.n11 VSUBS 0.01483f
C1446 VDD1.n12 VSUBS 0.035052f
C1447 VDD1.n13 VSUBS 0.015702f
C1448 VDD1.n14 VSUBS 0.027598f
C1449 VDD1.n15 VSUBS 0.01483f
C1450 VDD1.n16 VSUBS 0.035052f
C1451 VDD1.n17 VSUBS 0.015702f
C1452 VDD1.n18 VSUBS 0.027598f
C1453 VDD1.n19 VSUBS 0.01483f
C1454 VDD1.n20 VSUBS 0.035052f
C1455 VDD1.n21 VSUBS 0.015702f
C1456 VDD1.n22 VSUBS 0.027598f
C1457 VDD1.n23 VSUBS 0.01483f
C1458 VDD1.n24 VSUBS 0.035052f
C1459 VDD1.n25 VSUBS 0.015702f
C1460 VDD1.n26 VSUBS 0.193076f
C1461 VDD1.t5 VSUBS 0.075028f
C1462 VDD1.n27 VSUBS 0.026289f
C1463 VDD1.n28 VSUBS 0.022299f
C1464 VDD1.n29 VSUBS 0.01483f
C1465 VDD1.n30 VSUBS 1.73962f
C1466 VDD1.n31 VSUBS 0.027598f
C1467 VDD1.n32 VSUBS 0.01483f
C1468 VDD1.n33 VSUBS 0.015702f
C1469 VDD1.n34 VSUBS 0.035052f
C1470 VDD1.n35 VSUBS 0.035052f
C1471 VDD1.n36 VSUBS 0.015702f
C1472 VDD1.n37 VSUBS 0.01483f
C1473 VDD1.n38 VSUBS 0.027598f
C1474 VDD1.n39 VSUBS 0.027598f
C1475 VDD1.n40 VSUBS 0.01483f
C1476 VDD1.n41 VSUBS 0.015702f
C1477 VDD1.n42 VSUBS 0.035052f
C1478 VDD1.n43 VSUBS 0.035052f
C1479 VDD1.n44 VSUBS 0.015702f
C1480 VDD1.n45 VSUBS 0.01483f
C1481 VDD1.n46 VSUBS 0.027598f
C1482 VDD1.n47 VSUBS 0.027598f
C1483 VDD1.n48 VSUBS 0.01483f
C1484 VDD1.n49 VSUBS 0.015702f
C1485 VDD1.n50 VSUBS 0.035052f
C1486 VDD1.n51 VSUBS 0.035052f
C1487 VDD1.n52 VSUBS 0.015702f
C1488 VDD1.n53 VSUBS 0.01483f
C1489 VDD1.n54 VSUBS 0.027598f
C1490 VDD1.n55 VSUBS 0.027598f
C1491 VDD1.n56 VSUBS 0.01483f
C1492 VDD1.n57 VSUBS 0.015702f
C1493 VDD1.n58 VSUBS 0.035052f
C1494 VDD1.n59 VSUBS 0.035052f
C1495 VDD1.n60 VSUBS 0.015702f
C1496 VDD1.n61 VSUBS 0.01483f
C1497 VDD1.n62 VSUBS 0.027598f
C1498 VDD1.n63 VSUBS 0.027598f
C1499 VDD1.n64 VSUBS 0.01483f
C1500 VDD1.n65 VSUBS 0.015702f
C1501 VDD1.n66 VSUBS 0.035052f
C1502 VDD1.n67 VSUBS 0.035052f
C1503 VDD1.n68 VSUBS 0.015702f
C1504 VDD1.n69 VSUBS 0.01483f
C1505 VDD1.n70 VSUBS 0.027598f
C1506 VDD1.n71 VSUBS 0.027598f
C1507 VDD1.n72 VSUBS 0.01483f
C1508 VDD1.n73 VSUBS 0.015266f
C1509 VDD1.n74 VSUBS 0.015266f
C1510 VDD1.n75 VSUBS 0.035052f
C1511 VDD1.n76 VSUBS 0.083668f
C1512 VDD1.n77 VSUBS 0.015702f
C1513 VDD1.n78 VSUBS 0.01483f
C1514 VDD1.n79 VSUBS 0.070577f
C1515 VDD1.n80 VSUBS 0.071772f
C1516 VDD1.n81 VSUBS 0.029975f
C1517 VDD1.n82 VSUBS 0.027598f
C1518 VDD1.n83 VSUBS 0.01483f
C1519 VDD1.n84 VSUBS 0.035052f
C1520 VDD1.n85 VSUBS 0.015702f
C1521 VDD1.n86 VSUBS 0.027598f
C1522 VDD1.n87 VSUBS 0.01483f
C1523 VDD1.n88 VSUBS 0.035052f
C1524 VDD1.n89 VSUBS 0.015702f
C1525 VDD1.n90 VSUBS 0.027598f
C1526 VDD1.n91 VSUBS 0.01483f
C1527 VDD1.n92 VSUBS 0.035052f
C1528 VDD1.n93 VSUBS 0.015702f
C1529 VDD1.n94 VSUBS 0.027598f
C1530 VDD1.n95 VSUBS 0.01483f
C1531 VDD1.n96 VSUBS 0.035052f
C1532 VDD1.n97 VSUBS 0.015702f
C1533 VDD1.n98 VSUBS 0.027598f
C1534 VDD1.n99 VSUBS 0.01483f
C1535 VDD1.n100 VSUBS 0.035052f
C1536 VDD1.n101 VSUBS 0.015702f
C1537 VDD1.n102 VSUBS 0.027598f
C1538 VDD1.n103 VSUBS 0.01483f
C1539 VDD1.n104 VSUBS 0.035052f
C1540 VDD1.n105 VSUBS 0.015702f
C1541 VDD1.n106 VSUBS 0.193076f
C1542 VDD1.t2 VSUBS 0.075028f
C1543 VDD1.n107 VSUBS 0.026289f
C1544 VDD1.n108 VSUBS 0.022299f
C1545 VDD1.n109 VSUBS 0.01483f
C1546 VDD1.n110 VSUBS 1.73962f
C1547 VDD1.n111 VSUBS 0.027598f
C1548 VDD1.n112 VSUBS 0.01483f
C1549 VDD1.n113 VSUBS 0.015702f
C1550 VDD1.n114 VSUBS 0.035052f
C1551 VDD1.n115 VSUBS 0.035052f
C1552 VDD1.n116 VSUBS 0.015702f
C1553 VDD1.n117 VSUBS 0.01483f
C1554 VDD1.n118 VSUBS 0.027598f
C1555 VDD1.n119 VSUBS 0.027598f
C1556 VDD1.n120 VSUBS 0.01483f
C1557 VDD1.n121 VSUBS 0.015702f
C1558 VDD1.n122 VSUBS 0.035052f
C1559 VDD1.n123 VSUBS 0.035052f
C1560 VDD1.n124 VSUBS 0.015702f
C1561 VDD1.n125 VSUBS 0.01483f
C1562 VDD1.n126 VSUBS 0.027598f
C1563 VDD1.n127 VSUBS 0.027598f
C1564 VDD1.n128 VSUBS 0.01483f
C1565 VDD1.n129 VSUBS 0.015702f
C1566 VDD1.n130 VSUBS 0.035052f
C1567 VDD1.n131 VSUBS 0.035052f
C1568 VDD1.n132 VSUBS 0.015702f
C1569 VDD1.n133 VSUBS 0.01483f
C1570 VDD1.n134 VSUBS 0.027598f
C1571 VDD1.n135 VSUBS 0.027598f
C1572 VDD1.n136 VSUBS 0.01483f
C1573 VDD1.n137 VSUBS 0.015702f
C1574 VDD1.n138 VSUBS 0.035052f
C1575 VDD1.n139 VSUBS 0.035052f
C1576 VDD1.n140 VSUBS 0.015702f
C1577 VDD1.n141 VSUBS 0.01483f
C1578 VDD1.n142 VSUBS 0.027598f
C1579 VDD1.n143 VSUBS 0.027598f
C1580 VDD1.n144 VSUBS 0.01483f
C1581 VDD1.n145 VSUBS 0.015702f
C1582 VDD1.n146 VSUBS 0.035052f
C1583 VDD1.n147 VSUBS 0.035052f
C1584 VDD1.n148 VSUBS 0.035052f
C1585 VDD1.n149 VSUBS 0.015702f
C1586 VDD1.n150 VSUBS 0.01483f
C1587 VDD1.n151 VSUBS 0.027598f
C1588 VDD1.n152 VSUBS 0.027598f
C1589 VDD1.n153 VSUBS 0.01483f
C1590 VDD1.n154 VSUBS 0.015266f
C1591 VDD1.n155 VSUBS 0.015266f
C1592 VDD1.n156 VSUBS 0.035052f
C1593 VDD1.n157 VSUBS 0.083668f
C1594 VDD1.n158 VSUBS 0.015702f
C1595 VDD1.n159 VSUBS 0.01483f
C1596 VDD1.n160 VSUBS 0.070577f
C1597 VDD1.n161 VSUBS 0.070877f
C1598 VDD1.t1 VSUBS 0.323204f
C1599 VDD1.t4 VSUBS 0.323204f
C1600 VDD1.n162 VSUBS 2.63975f
C1601 VDD1.n163 VSUBS 3.80592f
C1602 VDD1.t0 VSUBS 0.323204f
C1603 VDD1.t3 VSUBS 0.323204f
C1604 VDD1.n164 VSUBS 2.63217f
C1605 VDD1.n165 VSUBS 3.74183f
C1606 VP.t4 VSUBS 3.55523f
C1607 VP.n0 VSUBS 1.35026f
C1608 VP.n1 VSUBS 0.028712f
C1609 VP.n2 VSUBS 0.036971f
C1610 VP.n3 VSUBS 0.028712f
C1611 VP.t0 VSUBS 3.55523f
C1612 VP.n4 VSUBS 0.053243f
C1613 VP.n5 VSUBS 0.028712f
C1614 VP.n6 VSUBS 0.053243f
C1615 VP.t2 VSUBS 3.55523f
C1616 VP.n7 VSUBS 1.35026f
C1617 VP.n8 VSUBS 0.028712f
C1618 VP.n9 VSUBS 0.036971f
C1619 VP.n10 VSUBS 0.326526f
C1620 VP.t5 VSUBS 3.55523f
C1621 VP.t1 VSUBS 3.87458f
C1622 VP.n11 VSUBS 1.28073f
C1623 VP.n12 VSUBS 1.3451f
C1624 VP.n13 VSUBS 0.053243f
C1625 VP.n14 VSUBS 0.053243f
C1626 VP.n15 VSUBS 0.028712f
C1627 VP.n16 VSUBS 0.028712f
C1628 VP.n17 VSUBS 0.028712f
C1629 VP.n18 VSUBS 0.046503f
C1630 VP.n19 VSUBS 0.053243f
C1631 VP.n20 VSUBS 0.046935f
C1632 VP.n21 VSUBS 0.046333f
C1633 VP.n22 VSUBS 1.75121f
C1634 VP.n23 VSUBS 1.77085f
C1635 VP.t3 VSUBS 3.55523f
C1636 VP.n24 VSUBS 1.35026f
C1637 VP.n25 VSUBS 0.046935f
C1638 VP.n26 VSUBS 0.046333f
C1639 VP.n27 VSUBS 0.028712f
C1640 VP.n28 VSUBS 0.028712f
C1641 VP.n29 VSUBS 0.046503f
C1642 VP.n30 VSUBS 0.036971f
C1643 VP.n31 VSUBS 0.053243f
C1644 VP.n32 VSUBS 0.028712f
C1645 VP.n33 VSUBS 0.028712f
C1646 VP.n34 VSUBS 0.028712f
C1647 VP.n35 VSUBS 1.26559f
C1648 VP.n36 VSUBS 0.053243f
C1649 VP.n37 VSUBS 0.053243f
C1650 VP.n38 VSUBS 0.028712f
C1651 VP.n39 VSUBS 0.028712f
C1652 VP.n40 VSUBS 0.028712f
C1653 VP.n41 VSUBS 0.046503f
C1654 VP.n42 VSUBS 0.053243f
C1655 VP.n43 VSUBS 0.046935f
C1656 VP.n44 VSUBS 0.046333f
C1657 VP.n45 VSUBS 0.061985f
.ends

