* NGSPICE file created from diff_pair_sample_0850.ext - technology: sky130A

.subckt diff_pair_sample_0850 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=1.5939 ps=9.99 w=9.66 l=0.71
X1 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=3.7674 ps=20.1 w=9.66 l=0.71
X2 VDD1.t5 VP.t1 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=3.7674 ps=20.1 w=9.66 l=0.71
X3 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=1.5939 ps=9.99 w=9.66 l=0.71
X4 VTAIL.t7 VP.t2 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=1.5939 ps=9.99 w=9.66 l=0.71
X5 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=1.5939 ps=9.99 w=9.66 l=0.71
X6 VDD1.t1 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=1.5939 ps=9.99 w=9.66 l=0.71
X7 VDD1.t0 VP.t4 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=1.5939 ps=9.99 w=9.66 l=0.71
X8 VDD2.t2 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=1.5939 ps=9.99 w=9.66 l=0.71
X9 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=0 ps=0 w=9.66 l=0.71
X10 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=0 ps=0 w=9.66 l=0.71
X11 VDD2.t1 VN.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=3.7674 ps=20.1 w=9.66 l=0.71
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=0 ps=0 w=9.66 l=0.71
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.7674 pd=20.1 as=0 ps=0 w=9.66 l=0.71
X14 VTAIL.t10 VN.t5 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=1.5939 ps=9.99 w=9.66 l=0.71
X15 VDD1.t2 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.5939 pd=9.99 as=3.7674 ps=20.1 w=9.66 l=0.71
R0 VP.n3 VP.t4 405.014
R1 VP.n8 VP.t3 383.224
R2 VP.n12 VP.t0 383.224
R3 VP.n14 VP.t5 383.224
R4 VP.n6 VP.t1 383.224
R5 VP.n4 VP.t2 383.224
R6 VP.n15 VP.n14 161.3
R7 VP.n5 VP.n2 161.3
R8 VP.n7 VP.n6 161.3
R9 VP.n13 VP.n0 161.3
R10 VP.n12 VP.n11 161.3
R11 VP.n10 VP.n1 161.3
R12 VP.n9 VP.n8 161.3
R13 VP.n3 VP.n2 44.8565
R14 VP.n9 VP.n7 39.4778
R15 VP.n8 VP.n1 27.0217
R16 VP.n14 VP.n13 27.0217
R17 VP.n6 VP.n5 27.0217
R18 VP.n12 VP.n1 21.1793
R19 VP.n13 VP.n12 21.1793
R20 VP.n5 VP.n4 21.1793
R21 VP.n4 VP.n3 20.1275
R22 VP.n7 VP.n2 0.189894
R23 VP.n10 VP.n9 0.189894
R24 VP.n11 VP.n10 0.189894
R25 VP.n11 VP.n0 0.189894
R26 VP.n15 VP.n0 0.189894
R27 VP VP.n15 0.0516364
R28 VDD1 VDD1.t0 66.756
R29 VDD1.n1 VDD1.t1 66.6423
R30 VDD1.n1 VDD1.n0 64.1443
R31 VDD1.n3 VDD1.n2 63.9756
R32 VDD1.n3 VDD1.n1 35.988
R33 VDD1.n2 VDD1.t4 2.05019
R34 VDD1.n2 VDD1.t5 2.05019
R35 VDD1.n0 VDD1.t3 2.05019
R36 VDD1.n0 VDD1.t2 2.05019
R37 VDD1 VDD1.n3 0.166448
R38 VTAIL.n7 VTAIL.t11 49.3466
R39 VTAIL.n11 VTAIL.t3 49.3465
R40 VTAIL.n2 VTAIL.t4 49.3465
R41 VTAIL.n10 VTAIL.t8 49.3465
R42 VTAIL.n9 VTAIL.n8 47.297
R43 VTAIL.n6 VTAIL.n5 47.297
R44 VTAIL.n1 VTAIL.n0 47.2967
R45 VTAIL.n4 VTAIL.n3 47.2967
R46 VTAIL.n6 VTAIL.n4 22.4876
R47 VTAIL.n11 VTAIL.n10 21.591
R48 VTAIL.n0 VTAIL.t0 2.05019
R49 VTAIL.n0 VTAIL.t10 2.05019
R50 VTAIL.n3 VTAIL.t6 2.05019
R51 VTAIL.n3 VTAIL.t9 2.05019
R52 VTAIL.n8 VTAIL.t5 2.05019
R53 VTAIL.n8 VTAIL.t7 2.05019
R54 VTAIL.n5 VTAIL.t2 2.05019
R55 VTAIL.n5 VTAIL.t1 2.05019
R56 VTAIL.n9 VTAIL.n7 0.918603
R57 VTAIL.n2 VTAIL.n1 0.918603
R58 VTAIL.n7 VTAIL.n6 0.897052
R59 VTAIL.n10 VTAIL.n9 0.897052
R60 VTAIL.n4 VTAIL.n2 0.897052
R61 VTAIL VTAIL.n11 0.614724
R62 VTAIL VTAIL.n1 0.282828
R63 B.n571 B.n570 585
R64 B.n572 B.n571 585
R65 B.n240 B.n81 585
R66 B.n239 B.n238 585
R67 B.n237 B.n236 585
R68 B.n235 B.n234 585
R69 B.n233 B.n232 585
R70 B.n231 B.n230 585
R71 B.n229 B.n228 585
R72 B.n227 B.n226 585
R73 B.n225 B.n224 585
R74 B.n223 B.n222 585
R75 B.n221 B.n220 585
R76 B.n219 B.n218 585
R77 B.n217 B.n216 585
R78 B.n215 B.n214 585
R79 B.n213 B.n212 585
R80 B.n211 B.n210 585
R81 B.n209 B.n208 585
R82 B.n207 B.n206 585
R83 B.n205 B.n204 585
R84 B.n203 B.n202 585
R85 B.n201 B.n200 585
R86 B.n199 B.n198 585
R87 B.n197 B.n196 585
R88 B.n195 B.n194 585
R89 B.n193 B.n192 585
R90 B.n191 B.n190 585
R91 B.n189 B.n188 585
R92 B.n187 B.n186 585
R93 B.n185 B.n184 585
R94 B.n183 B.n182 585
R95 B.n181 B.n180 585
R96 B.n179 B.n178 585
R97 B.n177 B.n176 585
R98 B.n175 B.n174 585
R99 B.n173 B.n172 585
R100 B.n171 B.n170 585
R101 B.n169 B.n168 585
R102 B.n167 B.n166 585
R103 B.n165 B.n164 585
R104 B.n163 B.n162 585
R105 B.n161 B.n160 585
R106 B.n159 B.n158 585
R107 B.n157 B.n156 585
R108 B.n154 B.n153 585
R109 B.n152 B.n151 585
R110 B.n150 B.n149 585
R111 B.n148 B.n147 585
R112 B.n146 B.n145 585
R113 B.n144 B.n143 585
R114 B.n142 B.n141 585
R115 B.n140 B.n139 585
R116 B.n138 B.n137 585
R117 B.n136 B.n135 585
R118 B.n134 B.n133 585
R119 B.n132 B.n131 585
R120 B.n130 B.n129 585
R121 B.n128 B.n127 585
R122 B.n126 B.n125 585
R123 B.n124 B.n123 585
R124 B.n122 B.n121 585
R125 B.n120 B.n119 585
R126 B.n118 B.n117 585
R127 B.n116 B.n115 585
R128 B.n114 B.n113 585
R129 B.n112 B.n111 585
R130 B.n110 B.n109 585
R131 B.n108 B.n107 585
R132 B.n106 B.n105 585
R133 B.n104 B.n103 585
R134 B.n102 B.n101 585
R135 B.n100 B.n99 585
R136 B.n98 B.n97 585
R137 B.n96 B.n95 585
R138 B.n94 B.n93 585
R139 B.n92 B.n91 585
R140 B.n90 B.n89 585
R141 B.n88 B.n87 585
R142 B.n40 B.n39 585
R143 B.n569 B.n41 585
R144 B.n573 B.n41 585
R145 B.n568 B.n567 585
R146 B.n567 B.n37 585
R147 B.n566 B.n36 585
R148 B.n579 B.n36 585
R149 B.n565 B.n35 585
R150 B.n580 B.n35 585
R151 B.n564 B.n34 585
R152 B.n581 B.n34 585
R153 B.n563 B.n562 585
R154 B.n562 B.n30 585
R155 B.n561 B.n29 585
R156 B.n587 B.n29 585
R157 B.n560 B.n28 585
R158 B.n588 B.n28 585
R159 B.n559 B.n27 585
R160 B.n589 B.n27 585
R161 B.n558 B.n557 585
R162 B.n557 B.n23 585
R163 B.n556 B.n22 585
R164 B.n595 B.n22 585
R165 B.n555 B.n21 585
R166 B.n596 B.n21 585
R167 B.n554 B.n20 585
R168 B.n597 B.n20 585
R169 B.n553 B.n552 585
R170 B.n552 B.n16 585
R171 B.n551 B.n15 585
R172 B.n603 B.n15 585
R173 B.n550 B.n14 585
R174 B.n604 B.n14 585
R175 B.n549 B.n13 585
R176 B.n605 B.n13 585
R177 B.n548 B.n547 585
R178 B.n547 B.n12 585
R179 B.n546 B.n545 585
R180 B.n546 B.n8 585
R181 B.n544 B.n7 585
R182 B.n612 B.n7 585
R183 B.n543 B.n6 585
R184 B.n613 B.n6 585
R185 B.n542 B.n5 585
R186 B.n614 B.n5 585
R187 B.n541 B.n540 585
R188 B.n540 B.n4 585
R189 B.n539 B.n241 585
R190 B.n539 B.n538 585
R191 B.n528 B.n242 585
R192 B.n531 B.n242 585
R193 B.n530 B.n529 585
R194 B.n532 B.n530 585
R195 B.n527 B.n247 585
R196 B.n247 B.n246 585
R197 B.n526 B.n525 585
R198 B.n525 B.n524 585
R199 B.n249 B.n248 585
R200 B.n250 B.n249 585
R201 B.n517 B.n516 585
R202 B.n518 B.n517 585
R203 B.n515 B.n254 585
R204 B.n258 B.n254 585
R205 B.n514 B.n513 585
R206 B.n513 B.n512 585
R207 B.n256 B.n255 585
R208 B.n257 B.n256 585
R209 B.n505 B.n504 585
R210 B.n506 B.n505 585
R211 B.n503 B.n263 585
R212 B.n263 B.n262 585
R213 B.n502 B.n501 585
R214 B.n501 B.n500 585
R215 B.n265 B.n264 585
R216 B.n266 B.n265 585
R217 B.n493 B.n492 585
R218 B.n494 B.n493 585
R219 B.n491 B.n271 585
R220 B.n271 B.n270 585
R221 B.n490 B.n489 585
R222 B.n489 B.n488 585
R223 B.n273 B.n272 585
R224 B.n274 B.n273 585
R225 B.n481 B.n480 585
R226 B.n482 B.n481 585
R227 B.n277 B.n276 585
R228 B.n322 B.n321 585
R229 B.n323 B.n319 585
R230 B.n319 B.n278 585
R231 B.n325 B.n324 585
R232 B.n327 B.n318 585
R233 B.n330 B.n329 585
R234 B.n331 B.n317 585
R235 B.n333 B.n332 585
R236 B.n335 B.n316 585
R237 B.n338 B.n337 585
R238 B.n339 B.n315 585
R239 B.n341 B.n340 585
R240 B.n343 B.n314 585
R241 B.n346 B.n345 585
R242 B.n347 B.n313 585
R243 B.n349 B.n348 585
R244 B.n351 B.n312 585
R245 B.n354 B.n353 585
R246 B.n355 B.n311 585
R247 B.n357 B.n356 585
R248 B.n359 B.n310 585
R249 B.n362 B.n361 585
R250 B.n363 B.n309 585
R251 B.n365 B.n364 585
R252 B.n367 B.n308 585
R253 B.n370 B.n369 585
R254 B.n371 B.n307 585
R255 B.n373 B.n372 585
R256 B.n375 B.n306 585
R257 B.n378 B.n377 585
R258 B.n379 B.n305 585
R259 B.n381 B.n380 585
R260 B.n383 B.n304 585
R261 B.n386 B.n385 585
R262 B.n387 B.n301 585
R263 B.n390 B.n389 585
R264 B.n392 B.n300 585
R265 B.n395 B.n394 585
R266 B.n396 B.n299 585
R267 B.n398 B.n397 585
R268 B.n400 B.n298 585
R269 B.n403 B.n402 585
R270 B.n404 B.n297 585
R271 B.n409 B.n408 585
R272 B.n411 B.n296 585
R273 B.n414 B.n413 585
R274 B.n415 B.n295 585
R275 B.n417 B.n416 585
R276 B.n419 B.n294 585
R277 B.n422 B.n421 585
R278 B.n423 B.n293 585
R279 B.n425 B.n424 585
R280 B.n427 B.n292 585
R281 B.n430 B.n429 585
R282 B.n431 B.n291 585
R283 B.n433 B.n432 585
R284 B.n435 B.n290 585
R285 B.n438 B.n437 585
R286 B.n439 B.n289 585
R287 B.n441 B.n440 585
R288 B.n443 B.n288 585
R289 B.n446 B.n445 585
R290 B.n447 B.n287 585
R291 B.n449 B.n448 585
R292 B.n451 B.n286 585
R293 B.n454 B.n453 585
R294 B.n455 B.n285 585
R295 B.n457 B.n456 585
R296 B.n459 B.n284 585
R297 B.n462 B.n461 585
R298 B.n463 B.n283 585
R299 B.n465 B.n464 585
R300 B.n467 B.n282 585
R301 B.n470 B.n469 585
R302 B.n471 B.n281 585
R303 B.n473 B.n472 585
R304 B.n475 B.n280 585
R305 B.n478 B.n477 585
R306 B.n479 B.n279 585
R307 B.n484 B.n483 585
R308 B.n483 B.n482 585
R309 B.n485 B.n275 585
R310 B.n275 B.n274 585
R311 B.n487 B.n486 585
R312 B.n488 B.n487 585
R313 B.n269 B.n268 585
R314 B.n270 B.n269 585
R315 B.n496 B.n495 585
R316 B.n495 B.n494 585
R317 B.n497 B.n267 585
R318 B.n267 B.n266 585
R319 B.n499 B.n498 585
R320 B.n500 B.n499 585
R321 B.n261 B.n260 585
R322 B.n262 B.n261 585
R323 B.n508 B.n507 585
R324 B.n507 B.n506 585
R325 B.n509 B.n259 585
R326 B.n259 B.n257 585
R327 B.n511 B.n510 585
R328 B.n512 B.n511 585
R329 B.n253 B.n252 585
R330 B.n258 B.n253 585
R331 B.n520 B.n519 585
R332 B.n519 B.n518 585
R333 B.n521 B.n251 585
R334 B.n251 B.n250 585
R335 B.n523 B.n522 585
R336 B.n524 B.n523 585
R337 B.n245 B.n244 585
R338 B.n246 B.n245 585
R339 B.n534 B.n533 585
R340 B.n533 B.n532 585
R341 B.n535 B.n243 585
R342 B.n531 B.n243 585
R343 B.n537 B.n536 585
R344 B.n538 B.n537 585
R345 B.n3 B.n0 585
R346 B.n4 B.n3 585
R347 B.n611 B.n1 585
R348 B.n612 B.n611 585
R349 B.n610 B.n609 585
R350 B.n610 B.n8 585
R351 B.n608 B.n9 585
R352 B.n12 B.n9 585
R353 B.n607 B.n606 585
R354 B.n606 B.n605 585
R355 B.n11 B.n10 585
R356 B.n604 B.n11 585
R357 B.n602 B.n601 585
R358 B.n603 B.n602 585
R359 B.n600 B.n17 585
R360 B.n17 B.n16 585
R361 B.n599 B.n598 585
R362 B.n598 B.n597 585
R363 B.n19 B.n18 585
R364 B.n596 B.n19 585
R365 B.n594 B.n593 585
R366 B.n595 B.n594 585
R367 B.n592 B.n24 585
R368 B.n24 B.n23 585
R369 B.n591 B.n590 585
R370 B.n590 B.n589 585
R371 B.n26 B.n25 585
R372 B.n588 B.n26 585
R373 B.n586 B.n585 585
R374 B.n587 B.n586 585
R375 B.n584 B.n31 585
R376 B.n31 B.n30 585
R377 B.n583 B.n582 585
R378 B.n582 B.n581 585
R379 B.n33 B.n32 585
R380 B.n580 B.n33 585
R381 B.n578 B.n577 585
R382 B.n579 B.n578 585
R383 B.n576 B.n38 585
R384 B.n38 B.n37 585
R385 B.n575 B.n574 585
R386 B.n574 B.n573 585
R387 B.n615 B.n614 585
R388 B.n613 B.n2 585
R389 B.n85 B.t6 530.74
R390 B.n82 B.t14 530.74
R391 B.n405 B.t10 530.74
R392 B.n302 B.t17 530.74
R393 B.n574 B.n40 478.086
R394 B.n571 B.n41 478.086
R395 B.n481 B.n279 478.086
R396 B.n483 B.n277 478.086
R397 B.n572 B.n80 256.663
R398 B.n572 B.n79 256.663
R399 B.n572 B.n78 256.663
R400 B.n572 B.n77 256.663
R401 B.n572 B.n76 256.663
R402 B.n572 B.n75 256.663
R403 B.n572 B.n74 256.663
R404 B.n572 B.n73 256.663
R405 B.n572 B.n72 256.663
R406 B.n572 B.n71 256.663
R407 B.n572 B.n70 256.663
R408 B.n572 B.n69 256.663
R409 B.n572 B.n68 256.663
R410 B.n572 B.n67 256.663
R411 B.n572 B.n66 256.663
R412 B.n572 B.n65 256.663
R413 B.n572 B.n64 256.663
R414 B.n572 B.n63 256.663
R415 B.n572 B.n62 256.663
R416 B.n572 B.n61 256.663
R417 B.n572 B.n60 256.663
R418 B.n572 B.n59 256.663
R419 B.n572 B.n58 256.663
R420 B.n572 B.n57 256.663
R421 B.n572 B.n56 256.663
R422 B.n572 B.n55 256.663
R423 B.n572 B.n54 256.663
R424 B.n572 B.n53 256.663
R425 B.n572 B.n52 256.663
R426 B.n572 B.n51 256.663
R427 B.n572 B.n50 256.663
R428 B.n572 B.n49 256.663
R429 B.n572 B.n48 256.663
R430 B.n572 B.n47 256.663
R431 B.n572 B.n46 256.663
R432 B.n572 B.n45 256.663
R433 B.n572 B.n44 256.663
R434 B.n572 B.n43 256.663
R435 B.n572 B.n42 256.663
R436 B.n320 B.n278 256.663
R437 B.n326 B.n278 256.663
R438 B.n328 B.n278 256.663
R439 B.n334 B.n278 256.663
R440 B.n336 B.n278 256.663
R441 B.n342 B.n278 256.663
R442 B.n344 B.n278 256.663
R443 B.n350 B.n278 256.663
R444 B.n352 B.n278 256.663
R445 B.n358 B.n278 256.663
R446 B.n360 B.n278 256.663
R447 B.n366 B.n278 256.663
R448 B.n368 B.n278 256.663
R449 B.n374 B.n278 256.663
R450 B.n376 B.n278 256.663
R451 B.n382 B.n278 256.663
R452 B.n384 B.n278 256.663
R453 B.n391 B.n278 256.663
R454 B.n393 B.n278 256.663
R455 B.n399 B.n278 256.663
R456 B.n401 B.n278 256.663
R457 B.n410 B.n278 256.663
R458 B.n412 B.n278 256.663
R459 B.n418 B.n278 256.663
R460 B.n420 B.n278 256.663
R461 B.n426 B.n278 256.663
R462 B.n428 B.n278 256.663
R463 B.n434 B.n278 256.663
R464 B.n436 B.n278 256.663
R465 B.n442 B.n278 256.663
R466 B.n444 B.n278 256.663
R467 B.n450 B.n278 256.663
R468 B.n452 B.n278 256.663
R469 B.n458 B.n278 256.663
R470 B.n460 B.n278 256.663
R471 B.n466 B.n278 256.663
R472 B.n468 B.n278 256.663
R473 B.n474 B.n278 256.663
R474 B.n476 B.n278 256.663
R475 B.n617 B.n616 256.663
R476 B.n89 B.n88 163.367
R477 B.n93 B.n92 163.367
R478 B.n97 B.n96 163.367
R479 B.n101 B.n100 163.367
R480 B.n105 B.n104 163.367
R481 B.n109 B.n108 163.367
R482 B.n113 B.n112 163.367
R483 B.n117 B.n116 163.367
R484 B.n121 B.n120 163.367
R485 B.n125 B.n124 163.367
R486 B.n129 B.n128 163.367
R487 B.n133 B.n132 163.367
R488 B.n137 B.n136 163.367
R489 B.n141 B.n140 163.367
R490 B.n145 B.n144 163.367
R491 B.n149 B.n148 163.367
R492 B.n153 B.n152 163.367
R493 B.n158 B.n157 163.367
R494 B.n162 B.n161 163.367
R495 B.n166 B.n165 163.367
R496 B.n170 B.n169 163.367
R497 B.n174 B.n173 163.367
R498 B.n178 B.n177 163.367
R499 B.n182 B.n181 163.367
R500 B.n186 B.n185 163.367
R501 B.n190 B.n189 163.367
R502 B.n194 B.n193 163.367
R503 B.n198 B.n197 163.367
R504 B.n202 B.n201 163.367
R505 B.n206 B.n205 163.367
R506 B.n210 B.n209 163.367
R507 B.n214 B.n213 163.367
R508 B.n218 B.n217 163.367
R509 B.n222 B.n221 163.367
R510 B.n226 B.n225 163.367
R511 B.n230 B.n229 163.367
R512 B.n234 B.n233 163.367
R513 B.n238 B.n237 163.367
R514 B.n571 B.n81 163.367
R515 B.n481 B.n273 163.367
R516 B.n489 B.n273 163.367
R517 B.n489 B.n271 163.367
R518 B.n493 B.n271 163.367
R519 B.n493 B.n265 163.367
R520 B.n501 B.n265 163.367
R521 B.n501 B.n263 163.367
R522 B.n505 B.n263 163.367
R523 B.n505 B.n256 163.367
R524 B.n513 B.n256 163.367
R525 B.n513 B.n254 163.367
R526 B.n517 B.n254 163.367
R527 B.n517 B.n249 163.367
R528 B.n525 B.n249 163.367
R529 B.n525 B.n247 163.367
R530 B.n530 B.n247 163.367
R531 B.n530 B.n242 163.367
R532 B.n539 B.n242 163.367
R533 B.n540 B.n539 163.367
R534 B.n540 B.n5 163.367
R535 B.n6 B.n5 163.367
R536 B.n7 B.n6 163.367
R537 B.n546 B.n7 163.367
R538 B.n547 B.n546 163.367
R539 B.n547 B.n13 163.367
R540 B.n14 B.n13 163.367
R541 B.n15 B.n14 163.367
R542 B.n552 B.n15 163.367
R543 B.n552 B.n20 163.367
R544 B.n21 B.n20 163.367
R545 B.n22 B.n21 163.367
R546 B.n557 B.n22 163.367
R547 B.n557 B.n27 163.367
R548 B.n28 B.n27 163.367
R549 B.n29 B.n28 163.367
R550 B.n562 B.n29 163.367
R551 B.n562 B.n34 163.367
R552 B.n35 B.n34 163.367
R553 B.n36 B.n35 163.367
R554 B.n567 B.n36 163.367
R555 B.n567 B.n41 163.367
R556 B.n321 B.n319 163.367
R557 B.n325 B.n319 163.367
R558 B.n329 B.n327 163.367
R559 B.n333 B.n317 163.367
R560 B.n337 B.n335 163.367
R561 B.n341 B.n315 163.367
R562 B.n345 B.n343 163.367
R563 B.n349 B.n313 163.367
R564 B.n353 B.n351 163.367
R565 B.n357 B.n311 163.367
R566 B.n361 B.n359 163.367
R567 B.n365 B.n309 163.367
R568 B.n369 B.n367 163.367
R569 B.n373 B.n307 163.367
R570 B.n377 B.n375 163.367
R571 B.n381 B.n305 163.367
R572 B.n385 B.n383 163.367
R573 B.n390 B.n301 163.367
R574 B.n394 B.n392 163.367
R575 B.n398 B.n299 163.367
R576 B.n402 B.n400 163.367
R577 B.n409 B.n297 163.367
R578 B.n413 B.n411 163.367
R579 B.n417 B.n295 163.367
R580 B.n421 B.n419 163.367
R581 B.n425 B.n293 163.367
R582 B.n429 B.n427 163.367
R583 B.n433 B.n291 163.367
R584 B.n437 B.n435 163.367
R585 B.n441 B.n289 163.367
R586 B.n445 B.n443 163.367
R587 B.n449 B.n287 163.367
R588 B.n453 B.n451 163.367
R589 B.n457 B.n285 163.367
R590 B.n461 B.n459 163.367
R591 B.n465 B.n283 163.367
R592 B.n469 B.n467 163.367
R593 B.n473 B.n281 163.367
R594 B.n477 B.n475 163.367
R595 B.n483 B.n275 163.367
R596 B.n487 B.n275 163.367
R597 B.n487 B.n269 163.367
R598 B.n495 B.n269 163.367
R599 B.n495 B.n267 163.367
R600 B.n499 B.n267 163.367
R601 B.n499 B.n261 163.367
R602 B.n507 B.n261 163.367
R603 B.n507 B.n259 163.367
R604 B.n511 B.n259 163.367
R605 B.n511 B.n253 163.367
R606 B.n519 B.n253 163.367
R607 B.n519 B.n251 163.367
R608 B.n523 B.n251 163.367
R609 B.n523 B.n245 163.367
R610 B.n533 B.n245 163.367
R611 B.n533 B.n243 163.367
R612 B.n537 B.n243 163.367
R613 B.n537 B.n3 163.367
R614 B.n615 B.n3 163.367
R615 B.n611 B.n2 163.367
R616 B.n611 B.n610 163.367
R617 B.n610 B.n9 163.367
R618 B.n606 B.n9 163.367
R619 B.n606 B.n11 163.367
R620 B.n602 B.n11 163.367
R621 B.n602 B.n17 163.367
R622 B.n598 B.n17 163.367
R623 B.n598 B.n19 163.367
R624 B.n594 B.n19 163.367
R625 B.n594 B.n24 163.367
R626 B.n590 B.n24 163.367
R627 B.n590 B.n26 163.367
R628 B.n586 B.n26 163.367
R629 B.n586 B.n31 163.367
R630 B.n582 B.n31 163.367
R631 B.n582 B.n33 163.367
R632 B.n578 B.n33 163.367
R633 B.n578 B.n38 163.367
R634 B.n574 B.n38 163.367
R635 B.n82 B.t15 91.071
R636 B.n405 B.t13 91.071
R637 B.n85 B.t8 91.0592
R638 B.n302 B.t19 91.0592
R639 B.n482 B.n278 83.2278
R640 B.n573 B.n572 83.2278
R641 B.n42 B.n40 71.676
R642 B.n89 B.n43 71.676
R643 B.n93 B.n44 71.676
R644 B.n97 B.n45 71.676
R645 B.n101 B.n46 71.676
R646 B.n105 B.n47 71.676
R647 B.n109 B.n48 71.676
R648 B.n113 B.n49 71.676
R649 B.n117 B.n50 71.676
R650 B.n121 B.n51 71.676
R651 B.n125 B.n52 71.676
R652 B.n129 B.n53 71.676
R653 B.n133 B.n54 71.676
R654 B.n137 B.n55 71.676
R655 B.n141 B.n56 71.676
R656 B.n145 B.n57 71.676
R657 B.n149 B.n58 71.676
R658 B.n153 B.n59 71.676
R659 B.n158 B.n60 71.676
R660 B.n162 B.n61 71.676
R661 B.n166 B.n62 71.676
R662 B.n170 B.n63 71.676
R663 B.n174 B.n64 71.676
R664 B.n178 B.n65 71.676
R665 B.n182 B.n66 71.676
R666 B.n186 B.n67 71.676
R667 B.n190 B.n68 71.676
R668 B.n194 B.n69 71.676
R669 B.n198 B.n70 71.676
R670 B.n202 B.n71 71.676
R671 B.n206 B.n72 71.676
R672 B.n210 B.n73 71.676
R673 B.n214 B.n74 71.676
R674 B.n218 B.n75 71.676
R675 B.n222 B.n76 71.676
R676 B.n226 B.n77 71.676
R677 B.n230 B.n78 71.676
R678 B.n234 B.n79 71.676
R679 B.n238 B.n80 71.676
R680 B.n81 B.n80 71.676
R681 B.n237 B.n79 71.676
R682 B.n233 B.n78 71.676
R683 B.n229 B.n77 71.676
R684 B.n225 B.n76 71.676
R685 B.n221 B.n75 71.676
R686 B.n217 B.n74 71.676
R687 B.n213 B.n73 71.676
R688 B.n209 B.n72 71.676
R689 B.n205 B.n71 71.676
R690 B.n201 B.n70 71.676
R691 B.n197 B.n69 71.676
R692 B.n193 B.n68 71.676
R693 B.n189 B.n67 71.676
R694 B.n185 B.n66 71.676
R695 B.n181 B.n65 71.676
R696 B.n177 B.n64 71.676
R697 B.n173 B.n63 71.676
R698 B.n169 B.n62 71.676
R699 B.n165 B.n61 71.676
R700 B.n161 B.n60 71.676
R701 B.n157 B.n59 71.676
R702 B.n152 B.n58 71.676
R703 B.n148 B.n57 71.676
R704 B.n144 B.n56 71.676
R705 B.n140 B.n55 71.676
R706 B.n136 B.n54 71.676
R707 B.n132 B.n53 71.676
R708 B.n128 B.n52 71.676
R709 B.n124 B.n51 71.676
R710 B.n120 B.n50 71.676
R711 B.n116 B.n49 71.676
R712 B.n112 B.n48 71.676
R713 B.n108 B.n47 71.676
R714 B.n104 B.n46 71.676
R715 B.n100 B.n45 71.676
R716 B.n96 B.n44 71.676
R717 B.n92 B.n43 71.676
R718 B.n88 B.n42 71.676
R719 B.n320 B.n277 71.676
R720 B.n326 B.n325 71.676
R721 B.n329 B.n328 71.676
R722 B.n334 B.n333 71.676
R723 B.n337 B.n336 71.676
R724 B.n342 B.n341 71.676
R725 B.n345 B.n344 71.676
R726 B.n350 B.n349 71.676
R727 B.n353 B.n352 71.676
R728 B.n358 B.n357 71.676
R729 B.n361 B.n360 71.676
R730 B.n366 B.n365 71.676
R731 B.n369 B.n368 71.676
R732 B.n374 B.n373 71.676
R733 B.n377 B.n376 71.676
R734 B.n382 B.n381 71.676
R735 B.n385 B.n384 71.676
R736 B.n391 B.n390 71.676
R737 B.n394 B.n393 71.676
R738 B.n399 B.n398 71.676
R739 B.n402 B.n401 71.676
R740 B.n410 B.n409 71.676
R741 B.n413 B.n412 71.676
R742 B.n418 B.n417 71.676
R743 B.n421 B.n420 71.676
R744 B.n426 B.n425 71.676
R745 B.n429 B.n428 71.676
R746 B.n434 B.n433 71.676
R747 B.n437 B.n436 71.676
R748 B.n442 B.n441 71.676
R749 B.n445 B.n444 71.676
R750 B.n450 B.n449 71.676
R751 B.n453 B.n452 71.676
R752 B.n458 B.n457 71.676
R753 B.n461 B.n460 71.676
R754 B.n466 B.n465 71.676
R755 B.n469 B.n468 71.676
R756 B.n474 B.n473 71.676
R757 B.n477 B.n476 71.676
R758 B.n321 B.n320 71.676
R759 B.n327 B.n326 71.676
R760 B.n328 B.n317 71.676
R761 B.n335 B.n334 71.676
R762 B.n336 B.n315 71.676
R763 B.n343 B.n342 71.676
R764 B.n344 B.n313 71.676
R765 B.n351 B.n350 71.676
R766 B.n352 B.n311 71.676
R767 B.n359 B.n358 71.676
R768 B.n360 B.n309 71.676
R769 B.n367 B.n366 71.676
R770 B.n368 B.n307 71.676
R771 B.n375 B.n374 71.676
R772 B.n376 B.n305 71.676
R773 B.n383 B.n382 71.676
R774 B.n384 B.n301 71.676
R775 B.n392 B.n391 71.676
R776 B.n393 B.n299 71.676
R777 B.n400 B.n399 71.676
R778 B.n401 B.n297 71.676
R779 B.n411 B.n410 71.676
R780 B.n412 B.n295 71.676
R781 B.n419 B.n418 71.676
R782 B.n420 B.n293 71.676
R783 B.n427 B.n426 71.676
R784 B.n428 B.n291 71.676
R785 B.n435 B.n434 71.676
R786 B.n436 B.n289 71.676
R787 B.n443 B.n442 71.676
R788 B.n444 B.n287 71.676
R789 B.n451 B.n450 71.676
R790 B.n452 B.n285 71.676
R791 B.n459 B.n458 71.676
R792 B.n460 B.n283 71.676
R793 B.n467 B.n466 71.676
R794 B.n468 B.n281 71.676
R795 B.n475 B.n474 71.676
R796 B.n476 B.n279 71.676
R797 B.n616 B.n615 71.676
R798 B.n616 B.n2 71.676
R799 B.n83 B.t16 70.9013
R800 B.n406 B.t12 70.9013
R801 B.n86 B.t9 70.8896
R802 B.n303 B.t18 70.8896
R803 B.n155 B.n86 59.5399
R804 B.n84 B.n83 59.5399
R805 B.n407 B.n406 59.5399
R806 B.n388 B.n303 59.5399
R807 B.n482 B.n274 50.0842
R808 B.n488 B.n274 50.0842
R809 B.n488 B.n270 50.0842
R810 B.n494 B.n270 50.0842
R811 B.n500 B.n266 50.0842
R812 B.n500 B.n262 50.0842
R813 B.n506 B.n262 50.0842
R814 B.n506 B.n257 50.0842
R815 B.n512 B.n257 50.0842
R816 B.n512 B.n258 50.0842
R817 B.n518 B.n250 50.0842
R818 B.n524 B.n250 50.0842
R819 B.n532 B.n246 50.0842
R820 B.n532 B.n531 50.0842
R821 B.n538 B.n4 50.0842
R822 B.n614 B.n4 50.0842
R823 B.n614 B.n613 50.0842
R824 B.n613 B.n612 50.0842
R825 B.n612 B.n8 50.0842
R826 B.n605 B.n12 50.0842
R827 B.n605 B.n604 50.0842
R828 B.n603 B.n16 50.0842
R829 B.n597 B.n16 50.0842
R830 B.n596 B.n595 50.0842
R831 B.n595 B.n23 50.0842
R832 B.n589 B.n23 50.0842
R833 B.n589 B.n588 50.0842
R834 B.n588 B.n587 50.0842
R835 B.n587 B.n30 50.0842
R836 B.n581 B.n580 50.0842
R837 B.n580 B.n579 50.0842
R838 B.n579 B.n37 50.0842
R839 B.n573 B.n37 50.0842
R840 B.n494 B.t11 49.3477
R841 B.n581 B.t7 49.3477
R842 B.n518 B.t2 37.5633
R843 B.n597 B.t3 37.5633
R844 B.t1 B.n246 34.6172
R845 B.n604 B.t5 34.6172
R846 B.n538 B.t4 31.6711
R847 B.t0 B.n8 31.6711
R848 B.n484 B.n276 31.0639
R849 B.n480 B.n479 31.0639
R850 B.n570 B.n569 31.0639
R851 B.n575 B.n39 31.0639
R852 B.n86 B.n85 20.1702
R853 B.n83 B.n82 20.1702
R854 B.n406 B.n405 20.1702
R855 B.n303 B.n302 20.1702
R856 B.n531 B.t4 18.4136
R857 B.n12 B.t0 18.4136
R858 B B.n617 18.0485
R859 B.n524 B.t1 15.4675
R860 B.t5 B.n603 15.4675
R861 B.n258 B.t2 12.5214
R862 B.t3 B.n596 12.5214
R863 B.n485 B.n484 10.6151
R864 B.n486 B.n485 10.6151
R865 B.n486 B.n268 10.6151
R866 B.n496 B.n268 10.6151
R867 B.n497 B.n496 10.6151
R868 B.n498 B.n497 10.6151
R869 B.n498 B.n260 10.6151
R870 B.n508 B.n260 10.6151
R871 B.n509 B.n508 10.6151
R872 B.n510 B.n509 10.6151
R873 B.n510 B.n252 10.6151
R874 B.n520 B.n252 10.6151
R875 B.n521 B.n520 10.6151
R876 B.n522 B.n521 10.6151
R877 B.n522 B.n244 10.6151
R878 B.n534 B.n244 10.6151
R879 B.n535 B.n534 10.6151
R880 B.n536 B.n535 10.6151
R881 B.n536 B.n0 10.6151
R882 B.n322 B.n276 10.6151
R883 B.n323 B.n322 10.6151
R884 B.n324 B.n323 10.6151
R885 B.n324 B.n318 10.6151
R886 B.n330 B.n318 10.6151
R887 B.n331 B.n330 10.6151
R888 B.n332 B.n331 10.6151
R889 B.n332 B.n316 10.6151
R890 B.n338 B.n316 10.6151
R891 B.n339 B.n338 10.6151
R892 B.n340 B.n339 10.6151
R893 B.n340 B.n314 10.6151
R894 B.n346 B.n314 10.6151
R895 B.n347 B.n346 10.6151
R896 B.n348 B.n347 10.6151
R897 B.n348 B.n312 10.6151
R898 B.n354 B.n312 10.6151
R899 B.n355 B.n354 10.6151
R900 B.n356 B.n355 10.6151
R901 B.n356 B.n310 10.6151
R902 B.n362 B.n310 10.6151
R903 B.n363 B.n362 10.6151
R904 B.n364 B.n363 10.6151
R905 B.n364 B.n308 10.6151
R906 B.n370 B.n308 10.6151
R907 B.n371 B.n370 10.6151
R908 B.n372 B.n371 10.6151
R909 B.n372 B.n306 10.6151
R910 B.n378 B.n306 10.6151
R911 B.n379 B.n378 10.6151
R912 B.n380 B.n379 10.6151
R913 B.n380 B.n304 10.6151
R914 B.n386 B.n304 10.6151
R915 B.n387 B.n386 10.6151
R916 B.n389 B.n300 10.6151
R917 B.n395 B.n300 10.6151
R918 B.n396 B.n395 10.6151
R919 B.n397 B.n396 10.6151
R920 B.n397 B.n298 10.6151
R921 B.n403 B.n298 10.6151
R922 B.n404 B.n403 10.6151
R923 B.n408 B.n404 10.6151
R924 B.n414 B.n296 10.6151
R925 B.n415 B.n414 10.6151
R926 B.n416 B.n415 10.6151
R927 B.n416 B.n294 10.6151
R928 B.n422 B.n294 10.6151
R929 B.n423 B.n422 10.6151
R930 B.n424 B.n423 10.6151
R931 B.n424 B.n292 10.6151
R932 B.n430 B.n292 10.6151
R933 B.n431 B.n430 10.6151
R934 B.n432 B.n431 10.6151
R935 B.n432 B.n290 10.6151
R936 B.n438 B.n290 10.6151
R937 B.n439 B.n438 10.6151
R938 B.n440 B.n439 10.6151
R939 B.n440 B.n288 10.6151
R940 B.n446 B.n288 10.6151
R941 B.n447 B.n446 10.6151
R942 B.n448 B.n447 10.6151
R943 B.n448 B.n286 10.6151
R944 B.n454 B.n286 10.6151
R945 B.n455 B.n454 10.6151
R946 B.n456 B.n455 10.6151
R947 B.n456 B.n284 10.6151
R948 B.n462 B.n284 10.6151
R949 B.n463 B.n462 10.6151
R950 B.n464 B.n463 10.6151
R951 B.n464 B.n282 10.6151
R952 B.n470 B.n282 10.6151
R953 B.n471 B.n470 10.6151
R954 B.n472 B.n471 10.6151
R955 B.n472 B.n280 10.6151
R956 B.n478 B.n280 10.6151
R957 B.n479 B.n478 10.6151
R958 B.n480 B.n272 10.6151
R959 B.n490 B.n272 10.6151
R960 B.n491 B.n490 10.6151
R961 B.n492 B.n491 10.6151
R962 B.n492 B.n264 10.6151
R963 B.n502 B.n264 10.6151
R964 B.n503 B.n502 10.6151
R965 B.n504 B.n503 10.6151
R966 B.n504 B.n255 10.6151
R967 B.n514 B.n255 10.6151
R968 B.n515 B.n514 10.6151
R969 B.n516 B.n515 10.6151
R970 B.n516 B.n248 10.6151
R971 B.n526 B.n248 10.6151
R972 B.n527 B.n526 10.6151
R973 B.n529 B.n527 10.6151
R974 B.n529 B.n528 10.6151
R975 B.n528 B.n241 10.6151
R976 B.n541 B.n241 10.6151
R977 B.n542 B.n541 10.6151
R978 B.n543 B.n542 10.6151
R979 B.n544 B.n543 10.6151
R980 B.n545 B.n544 10.6151
R981 B.n548 B.n545 10.6151
R982 B.n549 B.n548 10.6151
R983 B.n550 B.n549 10.6151
R984 B.n551 B.n550 10.6151
R985 B.n553 B.n551 10.6151
R986 B.n554 B.n553 10.6151
R987 B.n555 B.n554 10.6151
R988 B.n556 B.n555 10.6151
R989 B.n558 B.n556 10.6151
R990 B.n559 B.n558 10.6151
R991 B.n560 B.n559 10.6151
R992 B.n561 B.n560 10.6151
R993 B.n563 B.n561 10.6151
R994 B.n564 B.n563 10.6151
R995 B.n565 B.n564 10.6151
R996 B.n566 B.n565 10.6151
R997 B.n568 B.n566 10.6151
R998 B.n569 B.n568 10.6151
R999 B.n609 B.n1 10.6151
R1000 B.n609 B.n608 10.6151
R1001 B.n608 B.n607 10.6151
R1002 B.n607 B.n10 10.6151
R1003 B.n601 B.n10 10.6151
R1004 B.n601 B.n600 10.6151
R1005 B.n600 B.n599 10.6151
R1006 B.n599 B.n18 10.6151
R1007 B.n593 B.n18 10.6151
R1008 B.n593 B.n592 10.6151
R1009 B.n592 B.n591 10.6151
R1010 B.n591 B.n25 10.6151
R1011 B.n585 B.n25 10.6151
R1012 B.n585 B.n584 10.6151
R1013 B.n584 B.n583 10.6151
R1014 B.n583 B.n32 10.6151
R1015 B.n577 B.n32 10.6151
R1016 B.n577 B.n576 10.6151
R1017 B.n576 B.n575 10.6151
R1018 B.n87 B.n39 10.6151
R1019 B.n90 B.n87 10.6151
R1020 B.n91 B.n90 10.6151
R1021 B.n94 B.n91 10.6151
R1022 B.n95 B.n94 10.6151
R1023 B.n98 B.n95 10.6151
R1024 B.n99 B.n98 10.6151
R1025 B.n102 B.n99 10.6151
R1026 B.n103 B.n102 10.6151
R1027 B.n106 B.n103 10.6151
R1028 B.n107 B.n106 10.6151
R1029 B.n110 B.n107 10.6151
R1030 B.n111 B.n110 10.6151
R1031 B.n114 B.n111 10.6151
R1032 B.n115 B.n114 10.6151
R1033 B.n118 B.n115 10.6151
R1034 B.n119 B.n118 10.6151
R1035 B.n122 B.n119 10.6151
R1036 B.n123 B.n122 10.6151
R1037 B.n126 B.n123 10.6151
R1038 B.n127 B.n126 10.6151
R1039 B.n130 B.n127 10.6151
R1040 B.n131 B.n130 10.6151
R1041 B.n134 B.n131 10.6151
R1042 B.n135 B.n134 10.6151
R1043 B.n138 B.n135 10.6151
R1044 B.n139 B.n138 10.6151
R1045 B.n142 B.n139 10.6151
R1046 B.n143 B.n142 10.6151
R1047 B.n146 B.n143 10.6151
R1048 B.n147 B.n146 10.6151
R1049 B.n150 B.n147 10.6151
R1050 B.n151 B.n150 10.6151
R1051 B.n154 B.n151 10.6151
R1052 B.n159 B.n156 10.6151
R1053 B.n160 B.n159 10.6151
R1054 B.n163 B.n160 10.6151
R1055 B.n164 B.n163 10.6151
R1056 B.n167 B.n164 10.6151
R1057 B.n168 B.n167 10.6151
R1058 B.n171 B.n168 10.6151
R1059 B.n172 B.n171 10.6151
R1060 B.n176 B.n175 10.6151
R1061 B.n179 B.n176 10.6151
R1062 B.n180 B.n179 10.6151
R1063 B.n183 B.n180 10.6151
R1064 B.n184 B.n183 10.6151
R1065 B.n187 B.n184 10.6151
R1066 B.n188 B.n187 10.6151
R1067 B.n191 B.n188 10.6151
R1068 B.n192 B.n191 10.6151
R1069 B.n195 B.n192 10.6151
R1070 B.n196 B.n195 10.6151
R1071 B.n199 B.n196 10.6151
R1072 B.n200 B.n199 10.6151
R1073 B.n203 B.n200 10.6151
R1074 B.n204 B.n203 10.6151
R1075 B.n207 B.n204 10.6151
R1076 B.n208 B.n207 10.6151
R1077 B.n211 B.n208 10.6151
R1078 B.n212 B.n211 10.6151
R1079 B.n215 B.n212 10.6151
R1080 B.n216 B.n215 10.6151
R1081 B.n219 B.n216 10.6151
R1082 B.n220 B.n219 10.6151
R1083 B.n223 B.n220 10.6151
R1084 B.n224 B.n223 10.6151
R1085 B.n227 B.n224 10.6151
R1086 B.n228 B.n227 10.6151
R1087 B.n231 B.n228 10.6151
R1088 B.n232 B.n231 10.6151
R1089 B.n235 B.n232 10.6151
R1090 B.n236 B.n235 10.6151
R1091 B.n239 B.n236 10.6151
R1092 B.n240 B.n239 10.6151
R1093 B.n570 B.n240 10.6151
R1094 B.n617 B.n0 8.11757
R1095 B.n617 B.n1 8.11757
R1096 B.n389 B.n388 6.5566
R1097 B.n408 B.n407 6.5566
R1098 B.n156 B.n155 6.5566
R1099 B.n172 B.n84 6.5566
R1100 B.n388 B.n387 4.05904
R1101 B.n407 B.n296 4.05904
R1102 B.n155 B.n154 4.05904
R1103 B.n175 B.n84 4.05904
R1104 B.t11 B.n266 0.737025
R1105 B.t7 B.n30 0.737025
R1106 VN.n1 VN.t3 405.014
R1107 VN.n7 VN.t4 405.014
R1108 VN.n2 VN.t5 383.224
R1109 VN.n4 VN.t0 383.224
R1110 VN.n8 VN.t2 383.224
R1111 VN.n10 VN.t1 383.224
R1112 VN.n5 VN.n4 161.3
R1113 VN.n11 VN.n10 161.3
R1114 VN.n9 VN.n6 161.3
R1115 VN.n3 VN.n0 161.3
R1116 VN.n7 VN.n6 44.8565
R1117 VN.n1 VN.n0 44.8565
R1118 VN VN.n11 39.8585
R1119 VN.n4 VN.n3 27.0217
R1120 VN.n10 VN.n9 27.0217
R1121 VN.n3 VN.n2 21.1793
R1122 VN.n9 VN.n8 21.1793
R1123 VN.n2 VN.n1 20.1275
R1124 VN.n8 VN.n7 20.1275
R1125 VN.n11 VN.n6 0.189894
R1126 VN.n5 VN.n0 0.189894
R1127 VN VN.n5 0.0516364
R1128 VDD2.n1 VDD2.t2 66.6423
R1129 VDD2.n2 VDD2.t4 66.0254
R1130 VDD2.n1 VDD2.n0 64.1443
R1131 VDD2 VDD2.n3 64.1415
R1132 VDD2.n2 VDD2.n1 34.9567
R1133 VDD2.n3 VDD2.t3 2.05019
R1134 VDD2.n3 VDD2.t1 2.05019
R1135 VDD2.n0 VDD2.t0 2.05019
R1136 VDD2.n0 VDD2.t5 2.05019
R1137 VDD2 VDD2.n2 0.731103
C0 VP VN 4.65512f
C1 VDD1 VTAIL 8.32172f
C2 VDD1 VDD2 0.712349f
C3 VTAIL VP 3.38057f
C4 VDD2 VP 0.298241f
C5 VDD1 VP 3.73034f
C6 VTAIL VN 3.36606f
C7 VDD2 VN 3.58408f
C8 VDD1 VN 0.148281f
C9 VTAIL VDD2 8.35719f
C10 VDD2 B 4.077812f
C11 VDD1 B 4.306287f
C12 VTAIL B 5.534708f
C13 VN B 7.49353f
C14 VP B 5.638089f
C15 VDD2.t2 B 2.0065f
C16 VDD2.t0 B 0.179071f
C17 VDD2.t5 B 0.179071f
C18 VDD2.n0 B 1.5745f
C19 VDD2.n1 B 1.81749f
C20 VDD2.t4 B 2.00368f
C21 VDD2.n2 B 1.96044f
C22 VDD2.t3 B 0.179071f
C23 VDD2.t1 B 0.179071f
C24 VDD2.n3 B 1.57447f
C25 VN.n0 B 0.19291f
C26 VN.t3 B 0.931321f
C27 VN.n1 B 0.361338f
C28 VN.t5 B 0.911035f
C29 VN.n2 B 0.380957f
C30 VN.n3 B 0.010527f
C31 VN.t0 B 0.911035f
C32 VN.n4 B 0.374055f
C33 VN.n5 B 0.03595f
C34 VN.n6 B 0.19291f
C35 VN.t4 B 0.931321f
C36 VN.n7 B 0.361338f
C37 VN.t2 B 0.911035f
C38 VN.n8 B 0.380957f
C39 VN.n9 B 0.010527f
C40 VN.t1 B 0.911035f
C41 VN.n10 B 0.374055f
C42 VN.n11 B 1.75361f
C43 VTAIL.t0 B 0.18906f
C44 VTAIL.t10 B 0.18906f
C45 VTAIL.n0 B 1.59253f
C46 VTAIL.n1 B 0.33156f
C47 VTAIL.t4 B 2.02843f
C48 VTAIL.n2 B 0.460295f
C49 VTAIL.t6 B 0.18906f
C50 VTAIL.t9 B 0.18906f
C51 VTAIL.n3 B 1.59253f
C52 VTAIL.n4 B 1.45141f
C53 VTAIL.t2 B 0.18906f
C54 VTAIL.t1 B 0.18906f
C55 VTAIL.n5 B 1.59253f
C56 VTAIL.n6 B 1.4514f
C57 VTAIL.t11 B 2.02844f
C58 VTAIL.n7 B 0.460281f
C59 VTAIL.t5 B 0.18906f
C60 VTAIL.t7 B 0.18906f
C61 VTAIL.n8 B 1.59253f
C62 VTAIL.n9 B 0.380573f
C63 VTAIL.t8 B 2.02843f
C64 VTAIL.n10 B 1.45958f
C65 VTAIL.t3 B 2.02843f
C66 VTAIL.n11 B 1.43704f
C67 VDD1.t0 B 1.99272f
C68 VDD1.t1 B 1.99211f
C69 VDD1.t3 B 0.177787f
C70 VDD1.t2 B 0.177787f
C71 VDD1.n0 B 1.56321f
C72 VDD1.n1 B 1.87573f
C73 VDD1.t4 B 0.177787f
C74 VDD1.t5 B 0.177787f
C75 VDD1.n2 B 1.56247f
C76 VDD1.n3 B 1.92802f
C77 VP.n0 B 0.047048f
C78 VP.n1 B 0.010676f
C79 VP.n2 B 0.19565f
C80 VP.t1 B 0.923971f
C81 VP.t2 B 0.923971f
C82 VP.t4 B 0.944546f
C83 VP.n3 B 0.366468f
C84 VP.n4 B 0.386367f
C85 VP.n5 B 0.010676f
C86 VP.n6 B 0.379366f
C87 VP.n7 B 1.7475f
C88 VP.t3 B 0.923971f
C89 VP.n8 B 0.379366f
C90 VP.n9 B 1.79047f
C91 VP.n10 B 0.047048f
C92 VP.n11 B 0.047048f
C93 VP.t0 B 0.923971f
C94 VP.n12 B 0.382412f
C95 VP.n13 B 0.010676f
C96 VP.t5 B 0.923971f
C97 VP.n14 B 0.379366f
C98 VP.n15 B 0.036461f
.ends

