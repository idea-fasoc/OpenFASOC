* NGSPICE file created from diff_pair_sample_1009.ext - technology: sky130A

.subckt diff_pair_sample_1009 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=0 ps=0 w=7.64 l=0.63
X1 B.t8 B.t6 B.t7 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=0 ps=0 w=7.64 l=0.63
X2 B.t5 B.t3 B.t4 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=0 ps=0 w=7.64 l=0.63
X3 B.t2 B.t0 B.t1 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=0 ps=0 w=7.64 l=0.63
X4 VDD2.t1 VN.t0 VTAIL.t3 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=2.9796 ps=16.06 w=7.64 l=0.63
X5 VDD2.t0 VN.t1 VTAIL.t2 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=2.9796 ps=16.06 w=7.64 l=0.63
X6 VDD1.t1 VP.t0 VTAIL.t1 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=2.9796 ps=16.06 w=7.64 l=0.63
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1354_n2500# sky130_fd_pr__pfet_01v8 ad=2.9796 pd=16.06 as=2.9796 ps=16.06 w=7.64 l=0.63
R0 B.n223 B.n60 585
R1 B.n222 B.n221 585
R2 B.n220 B.n61 585
R3 B.n219 B.n218 585
R4 B.n217 B.n62 585
R5 B.n216 B.n215 585
R6 B.n214 B.n63 585
R7 B.n213 B.n212 585
R8 B.n211 B.n64 585
R9 B.n210 B.n209 585
R10 B.n208 B.n65 585
R11 B.n207 B.n206 585
R12 B.n205 B.n66 585
R13 B.n204 B.n203 585
R14 B.n202 B.n67 585
R15 B.n201 B.n200 585
R16 B.n199 B.n68 585
R17 B.n198 B.n197 585
R18 B.n196 B.n69 585
R19 B.n195 B.n194 585
R20 B.n193 B.n70 585
R21 B.n192 B.n191 585
R22 B.n190 B.n71 585
R23 B.n189 B.n188 585
R24 B.n187 B.n72 585
R25 B.n186 B.n185 585
R26 B.n184 B.n73 585
R27 B.n183 B.n182 585
R28 B.n181 B.n74 585
R29 B.n180 B.n179 585
R30 B.n175 B.n75 585
R31 B.n174 B.n173 585
R32 B.n172 B.n76 585
R33 B.n171 B.n170 585
R34 B.n169 B.n77 585
R35 B.n168 B.n167 585
R36 B.n166 B.n78 585
R37 B.n165 B.n164 585
R38 B.n162 B.n79 585
R39 B.n161 B.n160 585
R40 B.n159 B.n82 585
R41 B.n158 B.n157 585
R42 B.n156 B.n83 585
R43 B.n155 B.n154 585
R44 B.n153 B.n84 585
R45 B.n152 B.n151 585
R46 B.n150 B.n85 585
R47 B.n149 B.n148 585
R48 B.n147 B.n86 585
R49 B.n146 B.n145 585
R50 B.n144 B.n87 585
R51 B.n143 B.n142 585
R52 B.n141 B.n88 585
R53 B.n140 B.n139 585
R54 B.n138 B.n89 585
R55 B.n137 B.n136 585
R56 B.n135 B.n90 585
R57 B.n134 B.n133 585
R58 B.n132 B.n91 585
R59 B.n131 B.n130 585
R60 B.n129 B.n92 585
R61 B.n128 B.n127 585
R62 B.n126 B.n93 585
R63 B.n125 B.n124 585
R64 B.n123 B.n94 585
R65 B.n122 B.n121 585
R66 B.n120 B.n95 585
R67 B.n225 B.n224 585
R68 B.n226 B.n59 585
R69 B.n228 B.n227 585
R70 B.n229 B.n58 585
R71 B.n231 B.n230 585
R72 B.n232 B.n57 585
R73 B.n234 B.n233 585
R74 B.n235 B.n56 585
R75 B.n237 B.n236 585
R76 B.n238 B.n55 585
R77 B.n240 B.n239 585
R78 B.n241 B.n54 585
R79 B.n243 B.n242 585
R80 B.n244 B.n53 585
R81 B.n246 B.n245 585
R82 B.n247 B.n52 585
R83 B.n249 B.n248 585
R84 B.n250 B.n51 585
R85 B.n252 B.n251 585
R86 B.n253 B.n50 585
R87 B.n255 B.n254 585
R88 B.n256 B.n49 585
R89 B.n258 B.n257 585
R90 B.n259 B.n48 585
R91 B.n261 B.n260 585
R92 B.n262 B.n47 585
R93 B.n264 B.n263 585
R94 B.n265 B.n46 585
R95 B.n368 B.n367 585
R96 B.n366 B.n9 585
R97 B.n365 B.n364 585
R98 B.n363 B.n10 585
R99 B.n362 B.n361 585
R100 B.n360 B.n11 585
R101 B.n359 B.n358 585
R102 B.n357 B.n12 585
R103 B.n356 B.n355 585
R104 B.n354 B.n13 585
R105 B.n353 B.n352 585
R106 B.n351 B.n14 585
R107 B.n350 B.n349 585
R108 B.n348 B.n15 585
R109 B.n347 B.n346 585
R110 B.n345 B.n16 585
R111 B.n344 B.n343 585
R112 B.n342 B.n17 585
R113 B.n341 B.n340 585
R114 B.n339 B.n18 585
R115 B.n338 B.n337 585
R116 B.n336 B.n19 585
R117 B.n335 B.n334 585
R118 B.n333 B.n20 585
R119 B.n332 B.n331 585
R120 B.n330 B.n21 585
R121 B.n329 B.n328 585
R122 B.n327 B.n22 585
R123 B.n326 B.n325 585
R124 B.n323 B.n23 585
R125 B.n322 B.n321 585
R126 B.n320 B.n26 585
R127 B.n319 B.n318 585
R128 B.n317 B.n27 585
R129 B.n316 B.n315 585
R130 B.n314 B.n28 585
R131 B.n313 B.n312 585
R132 B.n311 B.n29 585
R133 B.n309 B.n308 585
R134 B.n307 B.n32 585
R135 B.n306 B.n305 585
R136 B.n304 B.n33 585
R137 B.n303 B.n302 585
R138 B.n301 B.n34 585
R139 B.n300 B.n299 585
R140 B.n298 B.n35 585
R141 B.n297 B.n296 585
R142 B.n295 B.n36 585
R143 B.n294 B.n293 585
R144 B.n292 B.n37 585
R145 B.n291 B.n290 585
R146 B.n289 B.n38 585
R147 B.n288 B.n287 585
R148 B.n286 B.n39 585
R149 B.n285 B.n284 585
R150 B.n283 B.n40 585
R151 B.n282 B.n281 585
R152 B.n280 B.n41 585
R153 B.n279 B.n278 585
R154 B.n277 B.n42 585
R155 B.n276 B.n275 585
R156 B.n274 B.n43 585
R157 B.n273 B.n272 585
R158 B.n271 B.n44 585
R159 B.n270 B.n269 585
R160 B.n268 B.n45 585
R161 B.n267 B.n266 585
R162 B.n369 B.n8 585
R163 B.n371 B.n370 585
R164 B.n372 B.n7 585
R165 B.n374 B.n373 585
R166 B.n375 B.n6 585
R167 B.n377 B.n376 585
R168 B.n378 B.n5 585
R169 B.n380 B.n379 585
R170 B.n381 B.n4 585
R171 B.n383 B.n382 585
R172 B.n384 B.n3 585
R173 B.n386 B.n385 585
R174 B.n387 B.n0 585
R175 B.n2 B.n1 585
R176 B.n102 B.n101 585
R177 B.n104 B.n103 585
R178 B.n105 B.n100 585
R179 B.n107 B.n106 585
R180 B.n108 B.n99 585
R181 B.n110 B.n109 585
R182 B.n111 B.n98 585
R183 B.n113 B.n112 585
R184 B.n114 B.n97 585
R185 B.n116 B.n115 585
R186 B.n117 B.n96 585
R187 B.n119 B.n118 585
R188 B.n118 B.n95 564.573
R189 B.n224 B.n223 564.573
R190 B.n266 B.n265 564.573
R191 B.n369 B.n368 564.573
R192 B.n80 B.t0 496.182
R193 B.n176 B.t9 496.182
R194 B.n30 B.t6 496.182
R195 B.n24 B.t3 496.182
R196 B.n389 B.n388 256.663
R197 B.n388 B.n387 235.042
R198 B.n388 B.n2 235.042
R199 B.n122 B.n95 163.367
R200 B.n123 B.n122 163.367
R201 B.n124 B.n123 163.367
R202 B.n124 B.n93 163.367
R203 B.n128 B.n93 163.367
R204 B.n129 B.n128 163.367
R205 B.n130 B.n129 163.367
R206 B.n130 B.n91 163.367
R207 B.n134 B.n91 163.367
R208 B.n135 B.n134 163.367
R209 B.n136 B.n135 163.367
R210 B.n136 B.n89 163.367
R211 B.n140 B.n89 163.367
R212 B.n141 B.n140 163.367
R213 B.n142 B.n141 163.367
R214 B.n142 B.n87 163.367
R215 B.n146 B.n87 163.367
R216 B.n147 B.n146 163.367
R217 B.n148 B.n147 163.367
R218 B.n148 B.n85 163.367
R219 B.n152 B.n85 163.367
R220 B.n153 B.n152 163.367
R221 B.n154 B.n153 163.367
R222 B.n154 B.n83 163.367
R223 B.n158 B.n83 163.367
R224 B.n159 B.n158 163.367
R225 B.n160 B.n159 163.367
R226 B.n160 B.n79 163.367
R227 B.n165 B.n79 163.367
R228 B.n166 B.n165 163.367
R229 B.n167 B.n166 163.367
R230 B.n167 B.n77 163.367
R231 B.n171 B.n77 163.367
R232 B.n172 B.n171 163.367
R233 B.n173 B.n172 163.367
R234 B.n173 B.n75 163.367
R235 B.n180 B.n75 163.367
R236 B.n181 B.n180 163.367
R237 B.n182 B.n181 163.367
R238 B.n182 B.n73 163.367
R239 B.n186 B.n73 163.367
R240 B.n187 B.n186 163.367
R241 B.n188 B.n187 163.367
R242 B.n188 B.n71 163.367
R243 B.n192 B.n71 163.367
R244 B.n193 B.n192 163.367
R245 B.n194 B.n193 163.367
R246 B.n194 B.n69 163.367
R247 B.n198 B.n69 163.367
R248 B.n199 B.n198 163.367
R249 B.n200 B.n199 163.367
R250 B.n200 B.n67 163.367
R251 B.n204 B.n67 163.367
R252 B.n205 B.n204 163.367
R253 B.n206 B.n205 163.367
R254 B.n206 B.n65 163.367
R255 B.n210 B.n65 163.367
R256 B.n211 B.n210 163.367
R257 B.n212 B.n211 163.367
R258 B.n212 B.n63 163.367
R259 B.n216 B.n63 163.367
R260 B.n217 B.n216 163.367
R261 B.n218 B.n217 163.367
R262 B.n218 B.n61 163.367
R263 B.n222 B.n61 163.367
R264 B.n223 B.n222 163.367
R265 B.n265 B.n264 163.367
R266 B.n264 B.n47 163.367
R267 B.n260 B.n47 163.367
R268 B.n260 B.n259 163.367
R269 B.n259 B.n258 163.367
R270 B.n258 B.n49 163.367
R271 B.n254 B.n49 163.367
R272 B.n254 B.n253 163.367
R273 B.n253 B.n252 163.367
R274 B.n252 B.n51 163.367
R275 B.n248 B.n51 163.367
R276 B.n248 B.n247 163.367
R277 B.n247 B.n246 163.367
R278 B.n246 B.n53 163.367
R279 B.n242 B.n53 163.367
R280 B.n242 B.n241 163.367
R281 B.n241 B.n240 163.367
R282 B.n240 B.n55 163.367
R283 B.n236 B.n55 163.367
R284 B.n236 B.n235 163.367
R285 B.n235 B.n234 163.367
R286 B.n234 B.n57 163.367
R287 B.n230 B.n57 163.367
R288 B.n230 B.n229 163.367
R289 B.n229 B.n228 163.367
R290 B.n228 B.n59 163.367
R291 B.n224 B.n59 163.367
R292 B.n368 B.n9 163.367
R293 B.n364 B.n9 163.367
R294 B.n364 B.n363 163.367
R295 B.n363 B.n362 163.367
R296 B.n362 B.n11 163.367
R297 B.n358 B.n11 163.367
R298 B.n358 B.n357 163.367
R299 B.n357 B.n356 163.367
R300 B.n356 B.n13 163.367
R301 B.n352 B.n13 163.367
R302 B.n352 B.n351 163.367
R303 B.n351 B.n350 163.367
R304 B.n350 B.n15 163.367
R305 B.n346 B.n15 163.367
R306 B.n346 B.n345 163.367
R307 B.n345 B.n344 163.367
R308 B.n344 B.n17 163.367
R309 B.n340 B.n17 163.367
R310 B.n340 B.n339 163.367
R311 B.n339 B.n338 163.367
R312 B.n338 B.n19 163.367
R313 B.n334 B.n19 163.367
R314 B.n334 B.n333 163.367
R315 B.n333 B.n332 163.367
R316 B.n332 B.n21 163.367
R317 B.n328 B.n21 163.367
R318 B.n328 B.n327 163.367
R319 B.n327 B.n326 163.367
R320 B.n326 B.n23 163.367
R321 B.n321 B.n23 163.367
R322 B.n321 B.n320 163.367
R323 B.n320 B.n319 163.367
R324 B.n319 B.n27 163.367
R325 B.n315 B.n27 163.367
R326 B.n315 B.n314 163.367
R327 B.n314 B.n313 163.367
R328 B.n313 B.n29 163.367
R329 B.n308 B.n29 163.367
R330 B.n308 B.n307 163.367
R331 B.n307 B.n306 163.367
R332 B.n306 B.n33 163.367
R333 B.n302 B.n33 163.367
R334 B.n302 B.n301 163.367
R335 B.n301 B.n300 163.367
R336 B.n300 B.n35 163.367
R337 B.n296 B.n35 163.367
R338 B.n296 B.n295 163.367
R339 B.n295 B.n294 163.367
R340 B.n294 B.n37 163.367
R341 B.n290 B.n37 163.367
R342 B.n290 B.n289 163.367
R343 B.n289 B.n288 163.367
R344 B.n288 B.n39 163.367
R345 B.n284 B.n39 163.367
R346 B.n284 B.n283 163.367
R347 B.n283 B.n282 163.367
R348 B.n282 B.n41 163.367
R349 B.n278 B.n41 163.367
R350 B.n278 B.n277 163.367
R351 B.n277 B.n276 163.367
R352 B.n276 B.n43 163.367
R353 B.n272 B.n43 163.367
R354 B.n272 B.n271 163.367
R355 B.n271 B.n270 163.367
R356 B.n270 B.n45 163.367
R357 B.n266 B.n45 163.367
R358 B.n370 B.n369 163.367
R359 B.n370 B.n7 163.367
R360 B.n374 B.n7 163.367
R361 B.n375 B.n374 163.367
R362 B.n376 B.n375 163.367
R363 B.n376 B.n5 163.367
R364 B.n380 B.n5 163.367
R365 B.n381 B.n380 163.367
R366 B.n382 B.n381 163.367
R367 B.n382 B.n3 163.367
R368 B.n386 B.n3 163.367
R369 B.n387 B.n386 163.367
R370 B.n101 B.n2 163.367
R371 B.n104 B.n101 163.367
R372 B.n105 B.n104 163.367
R373 B.n106 B.n105 163.367
R374 B.n106 B.n99 163.367
R375 B.n110 B.n99 163.367
R376 B.n111 B.n110 163.367
R377 B.n112 B.n111 163.367
R378 B.n112 B.n97 163.367
R379 B.n116 B.n97 163.367
R380 B.n117 B.n116 163.367
R381 B.n118 B.n117 163.367
R382 B.n176 B.t10 130.683
R383 B.n30 B.t8 130.683
R384 B.n80 B.t1 130.674
R385 B.n24 B.t5 130.674
R386 B.n177 B.t11 112.064
R387 B.n31 B.t7 112.064
R388 B.n81 B.t2 112.056
R389 B.n25 B.t4 112.056
R390 B.n163 B.n81 59.5399
R391 B.n178 B.n177 59.5399
R392 B.n310 B.n31 59.5399
R393 B.n324 B.n25 59.5399
R394 B.n367 B.n8 36.6834
R395 B.n267 B.n46 36.6834
R396 B.n225 B.n60 36.6834
R397 B.n120 B.n119 36.6834
R398 B.n81 B.n80 18.6187
R399 B.n177 B.n176 18.6187
R400 B.n31 B.n30 18.6187
R401 B.n25 B.n24 18.6187
R402 B B.n389 18.0485
R403 B.n371 B.n8 10.6151
R404 B.n372 B.n371 10.6151
R405 B.n373 B.n372 10.6151
R406 B.n373 B.n6 10.6151
R407 B.n377 B.n6 10.6151
R408 B.n378 B.n377 10.6151
R409 B.n379 B.n378 10.6151
R410 B.n379 B.n4 10.6151
R411 B.n383 B.n4 10.6151
R412 B.n384 B.n383 10.6151
R413 B.n385 B.n384 10.6151
R414 B.n385 B.n0 10.6151
R415 B.n367 B.n366 10.6151
R416 B.n366 B.n365 10.6151
R417 B.n365 B.n10 10.6151
R418 B.n361 B.n10 10.6151
R419 B.n361 B.n360 10.6151
R420 B.n360 B.n359 10.6151
R421 B.n359 B.n12 10.6151
R422 B.n355 B.n12 10.6151
R423 B.n355 B.n354 10.6151
R424 B.n354 B.n353 10.6151
R425 B.n353 B.n14 10.6151
R426 B.n349 B.n14 10.6151
R427 B.n349 B.n348 10.6151
R428 B.n348 B.n347 10.6151
R429 B.n347 B.n16 10.6151
R430 B.n343 B.n16 10.6151
R431 B.n343 B.n342 10.6151
R432 B.n342 B.n341 10.6151
R433 B.n341 B.n18 10.6151
R434 B.n337 B.n18 10.6151
R435 B.n337 B.n336 10.6151
R436 B.n336 B.n335 10.6151
R437 B.n335 B.n20 10.6151
R438 B.n331 B.n20 10.6151
R439 B.n331 B.n330 10.6151
R440 B.n330 B.n329 10.6151
R441 B.n329 B.n22 10.6151
R442 B.n325 B.n22 10.6151
R443 B.n323 B.n322 10.6151
R444 B.n322 B.n26 10.6151
R445 B.n318 B.n26 10.6151
R446 B.n318 B.n317 10.6151
R447 B.n317 B.n316 10.6151
R448 B.n316 B.n28 10.6151
R449 B.n312 B.n28 10.6151
R450 B.n312 B.n311 10.6151
R451 B.n309 B.n32 10.6151
R452 B.n305 B.n32 10.6151
R453 B.n305 B.n304 10.6151
R454 B.n304 B.n303 10.6151
R455 B.n303 B.n34 10.6151
R456 B.n299 B.n34 10.6151
R457 B.n299 B.n298 10.6151
R458 B.n298 B.n297 10.6151
R459 B.n297 B.n36 10.6151
R460 B.n293 B.n36 10.6151
R461 B.n293 B.n292 10.6151
R462 B.n292 B.n291 10.6151
R463 B.n291 B.n38 10.6151
R464 B.n287 B.n38 10.6151
R465 B.n287 B.n286 10.6151
R466 B.n286 B.n285 10.6151
R467 B.n285 B.n40 10.6151
R468 B.n281 B.n40 10.6151
R469 B.n281 B.n280 10.6151
R470 B.n280 B.n279 10.6151
R471 B.n279 B.n42 10.6151
R472 B.n275 B.n42 10.6151
R473 B.n275 B.n274 10.6151
R474 B.n274 B.n273 10.6151
R475 B.n273 B.n44 10.6151
R476 B.n269 B.n44 10.6151
R477 B.n269 B.n268 10.6151
R478 B.n268 B.n267 10.6151
R479 B.n263 B.n46 10.6151
R480 B.n263 B.n262 10.6151
R481 B.n262 B.n261 10.6151
R482 B.n261 B.n48 10.6151
R483 B.n257 B.n48 10.6151
R484 B.n257 B.n256 10.6151
R485 B.n256 B.n255 10.6151
R486 B.n255 B.n50 10.6151
R487 B.n251 B.n50 10.6151
R488 B.n251 B.n250 10.6151
R489 B.n250 B.n249 10.6151
R490 B.n249 B.n52 10.6151
R491 B.n245 B.n52 10.6151
R492 B.n245 B.n244 10.6151
R493 B.n244 B.n243 10.6151
R494 B.n243 B.n54 10.6151
R495 B.n239 B.n54 10.6151
R496 B.n239 B.n238 10.6151
R497 B.n238 B.n237 10.6151
R498 B.n237 B.n56 10.6151
R499 B.n233 B.n56 10.6151
R500 B.n233 B.n232 10.6151
R501 B.n232 B.n231 10.6151
R502 B.n231 B.n58 10.6151
R503 B.n227 B.n58 10.6151
R504 B.n227 B.n226 10.6151
R505 B.n226 B.n225 10.6151
R506 B.n102 B.n1 10.6151
R507 B.n103 B.n102 10.6151
R508 B.n103 B.n100 10.6151
R509 B.n107 B.n100 10.6151
R510 B.n108 B.n107 10.6151
R511 B.n109 B.n108 10.6151
R512 B.n109 B.n98 10.6151
R513 B.n113 B.n98 10.6151
R514 B.n114 B.n113 10.6151
R515 B.n115 B.n114 10.6151
R516 B.n115 B.n96 10.6151
R517 B.n119 B.n96 10.6151
R518 B.n121 B.n120 10.6151
R519 B.n121 B.n94 10.6151
R520 B.n125 B.n94 10.6151
R521 B.n126 B.n125 10.6151
R522 B.n127 B.n126 10.6151
R523 B.n127 B.n92 10.6151
R524 B.n131 B.n92 10.6151
R525 B.n132 B.n131 10.6151
R526 B.n133 B.n132 10.6151
R527 B.n133 B.n90 10.6151
R528 B.n137 B.n90 10.6151
R529 B.n138 B.n137 10.6151
R530 B.n139 B.n138 10.6151
R531 B.n139 B.n88 10.6151
R532 B.n143 B.n88 10.6151
R533 B.n144 B.n143 10.6151
R534 B.n145 B.n144 10.6151
R535 B.n145 B.n86 10.6151
R536 B.n149 B.n86 10.6151
R537 B.n150 B.n149 10.6151
R538 B.n151 B.n150 10.6151
R539 B.n151 B.n84 10.6151
R540 B.n155 B.n84 10.6151
R541 B.n156 B.n155 10.6151
R542 B.n157 B.n156 10.6151
R543 B.n157 B.n82 10.6151
R544 B.n161 B.n82 10.6151
R545 B.n162 B.n161 10.6151
R546 B.n164 B.n78 10.6151
R547 B.n168 B.n78 10.6151
R548 B.n169 B.n168 10.6151
R549 B.n170 B.n169 10.6151
R550 B.n170 B.n76 10.6151
R551 B.n174 B.n76 10.6151
R552 B.n175 B.n174 10.6151
R553 B.n179 B.n175 10.6151
R554 B.n183 B.n74 10.6151
R555 B.n184 B.n183 10.6151
R556 B.n185 B.n184 10.6151
R557 B.n185 B.n72 10.6151
R558 B.n189 B.n72 10.6151
R559 B.n190 B.n189 10.6151
R560 B.n191 B.n190 10.6151
R561 B.n191 B.n70 10.6151
R562 B.n195 B.n70 10.6151
R563 B.n196 B.n195 10.6151
R564 B.n197 B.n196 10.6151
R565 B.n197 B.n68 10.6151
R566 B.n201 B.n68 10.6151
R567 B.n202 B.n201 10.6151
R568 B.n203 B.n202 10.6151
R569 B.n203 B.n66 10.6151
R570 B.n207 B.n66 10.6151
R571 B.n208 B.n207 10.6151
R572 B.n209 B.n208 10.6151
R573 B.n209 B.n64 10.6151
R574 B.n213 B.n64 10.6151
R575 B.n214 B.n213 10.6151
R576 B.n215 B.n214 10.6151
R577 B.n215 B.n62 10.6151
R578 B.n219 B.n62 10.6151
R579 B.n220 B.n219 10.6151
R580 B.n221 B.n220 10.6151
R581 B.n221 B.n60 10.6151
R582 B.n389 B.n0 8.11757
R583 B.n389 B.n1 8.11757
R584 B.n324 B.n323 7.18099
R585 B.n311 B.n310 7.18099
R586 B.n164 B.n163 7.18099
R587 B.n179 B.n178 7.18099
R588 B.n325 B.n324 3.43465
R589 B.n310 B.n309 3.43465
R590 B.n163 B.n162 3.43465
R591 B.n178 B.n74 3.43465
R592 VN VN.t1 553.205
R593 VN VN.t0 516.731
R594 VTAIL.n1 VTAIL.t2 74.9947
R595 VTAIL.n3 VTAIL.t3 74.9945
R596 VTAIL.n0 VTAIL.t1 74.9945
R597 VTAIL.n2 VTAIL.t0 74.9945
R598 VTAIL.n1 VTAIL.n0 20.6255
R599 VTAIL.n3 VTAIL.n2 19.7979
R600 VTAIL.n2 VTAIL.n1 0.884121
R601 VTAIL VTAIL.n0 0.735414
R602 VTAIL VTAIL.n3 0.149207
R603 VDD2.n0 VDD2.t1 123.591
R604 VDD2.n0 VDD2.t0 91.6733
R605 VDD2 VDD2.n0 0.265586
R606 VP.n0 VP.t1 552.823
R607 VP.n0 VP.t0 516.679
R608 VP VP.n0 0.0516364
R609 VDD1 VDD1.t1 124.323
R610 VDD1 VDD1.t0 91.9384
C0 VDD2 VTAIL 4.15729f
C1 w_n1354_n2500# VDD2 1.24583f
C2 VDD2 VDD1 0.454242f
C3 VN B 0.662005f
C4 VP B 0.930673f
C5 VN VP 3.72477f
C6 VTAIL B 1.91193f
C7 w_n1354_n2500# B 5.46162f
C8 VN VTAIL 0.978246f
C9 w_n1354_n2500# VN 1.62473f
C10 VP VTAIL 0.992686f
C11 VDD1 B 1.08724f
C12 w_n1354_n2500# VP 1.79295f
C13 VN VDD1 0.148223f
C14 VDD1 VP 1.40013f
C15 w_n1354_n2500# VTAIL 2.20117f
C16 VDD1 VTAIL 4.12167f
C17 w_n1354_n2500# VDD1 1.24189f
C18 VDD2 B 1.10127f
C19 VN VDD2 1.30019f
C20 VDD2 VP 0.251078f
C21 VDD2 VSUBS 0.587375f
C22 VDD1 VSUBS 2.73373f
C23 VTAIL VSUBS 0.586831f
C24 VN VSUBS 3.95718f
C25 VP VSUBS 0.922201f
C26 B VSUBS 2.074956f
C27 w_n1354_n2500# VSUBS 42.0336f
C28 VDD1.t0 VSUBS 0.904146f
C29 VDD1.t1 VSUBS 1.16024f
C30 VP.t1 VSUBS 0.642005f
C31 VP.t0 VSUBS 0.558749f
C32 VP.n0 VSUBS 2.48839f
C33 VDD2.t1 VSUBS 1.19087f
C34 VDD2.t0 VSUBS 0.938564f
C35 VDD2.n0 VSUBS 2.03433f
C36 VTAIL.t1 VSUBS 1.1949f
C37 VTAIL.n0 VSUBS 1.44929f
C38 VTAIL.t2 VSUBS 1.19491f
C39 VTAIL.n1 VSUBS 1.46006f
C40 VTAIL.t0 VSUBS 1.1949f
C41 VTAIL.n2 VSUBS 1.40013f
C42 VTAIL.t3 VSUBS 1.1949f
C43 VTAIL.n3 VSUBS 1.34691f
C44 VN.t0 VSUBS 0.551315f
C45 VN.t1 VSUBS 0.635789f
C46 B.n0 VSUBS 0.005434f
C47 B.n1 VSUBS 0.005434f
C48 B.n2 VSUBS 0.008036f
C49 B.n3 VSUBS 0.006158f
C50 B.n4 VSUBS 0.006158f
C51 B.n5 VSUBS 0.006158f
C52 B.n6 VSUBS 0.006158f
C53 B.n7 VSUBS 0.006158f
C54 B.n8 VSUBS 0.015206f
C55 B.n9 VSUBS 0.006158f
C56 B.n10 VSUBS 0.006158f
C57 B.n11 VSUBS 0.006158f
C58 B.n12 VSUBS 0.006158f
C59 B.n13 VSUBS 0.006158f
C60 B.n14 VSUBS 0.006158f
C61 B.n15 VSUBS 0.006158f
C62 B.n16 VSUBS 0.006158f
C63 B.n17 VSUBS 0.006158f
C64 B.n18 VSUBS 0.006158f
C65 B.n19 VSUBS 0.006158f
C66 B.n20 VSUBS 0.006158f
C67 B.n21 VSUBS 0.006158f
C68 B.n22 VSUBS 0.006158f
C69 B.n23 VSUBS 0.006158f
C70 B.t4 VSUBS 0.205768f
C71 B.t5 VSUBS 0.212435f
C72 B.t3 VSUBS 0.178621f
C73 B.n24 VSUBS 0.085943f
C74 B.n25 VSUBS 0.055573f
C75 B.n26 VSUBS 0.006158f
C76 B.n27 VSUBS 0.006158f
C77 B.n28 VSUBS 0.006158f
C78 B.n29 VSUBS 0.006158f
C79 B.t7 VSUBS 0.205767f
C80 B.t8 VSUBS 0.212433f
C81 B.t6 VSUBS 0.178621f
C82 B.n30 VSUBS 0.085945f
C83 B.n31 VSUBS 0.055574f
C84 B.n32 VSUBS 0.006158f
C85 B.n33 VSUBS 0.006158f
C86 B.n34 VSUBS 0.006158f
C87 B.n35 VSUBS 0.006158f
C88 B.n36 VSUBS 0.006158f
C89 B.n37 VSUBS 0.006158f
C90 B.n38 VSUBS 0.006158f
C91 B.n39 VSUBS 0.006158f
C92 B.n40 VSUBS 0.006158f
C93 B.n41 VSUBS 0.006158f
C94 B.n42 VSUBS 0.006158f
C95 B.n43 VSUBS 0.006158f
C96 B.n44 VSUBS 0.006158f
C97 B.n45 VSUBS 0.006158f
C98 B.n46 VSUBS 0.015206f
C99 B.n47 VSUBS 0.006158f
C100 B.n48 VSUBS 0.006158f
C101 B.n49 VSUBS 0.006158f
C102 B.n50 VSUBS 0.006158f
C103 B.n51 VSUBS 0.006158f
C104 B.n52 VSUBS 0.006158f
C105 B.n53 VSUBS 0.006158f
C106 B.n54 VSUBS 0.006158f
C107 B.n55 VSUBS 0.006158f
C108 B.n56 VSUBS 0.006158f
C109 B.n57 VSUBS 0.006158f
C110 B.n58 VSUBS 0.006158f
C111 B.n59 VSUBS 0.006158f
C112 B.n60 VSUBS 0.0153f
C113 B.n61 VSUBS 0.006158f
C114 B.n62 VSUBS 0.006158f
C115 B.n63 VSUBS 0.006158f
C116 B.n64 VSUBS 0.006158f
C117 B.n65 VSUBS 0.006158f
C118 B.n66 VSUBS 0.006158f
C119 B.n67 VSUBS 0.006158f
C120 B.n68 VSUBS 0.006158f
C121 B.n69 VSUBS 0.006158f
C122 B.n70 VSUBS 0.006158f
C123 B.n71 VSUBS 0.006158f
C124 B.n72 VSUBS 0.006158f
C125 B.n73 VSUBS 0.006158f
C126 B.n74 VSUBS 0.004075f
C127 B.n75 VSUBS 0.006158f
C128 B.n76 VSUBS 0.006158f
C129 B.n77 VSUBS 0.006158f
C130 B.n78 VSUBS 0.006158f
C131 B.n79 VSUBS 0.006158f
C132 B.t2 VSUBS 0.205768f
C133 B.t1 VSUBS 0.212435f
C134 B.t0 VSUBS 0.178621f
C135 B.n80 VSUBS 0.085943f
C136 B.n81 VSUBS 0.055573f
C137 B.n82 VSUBS 0.006158f
C138 B.n83 VSUBS 0.006158f
C139 B.n84 VSUBS 0.006158f
C140 B.n85 VSUBS 0.006158f
C141 B.n86 VSUBS 0.006158f
C142 B.n87 VSUBS 0.006158f
C143 B.n88 VSUBS 0.006158f
C144 B.n89 VSUBS 0.006158f
C145 B.n90 VSUBS 0.006158f
C146 B.n91 VSUBS 0.006158f
C147 B.n92 VSUBS 0.006158f
C148 B.n93 VSUBS 0.006158f
C149 B.n94 VSUBS 0.006158f
C150 B.n95 VSUBS 0.015948f
C151 B.n96 VSUBS 0.006158f
C152 B.n97 VSUBS 0.006158f
C153 B.n98 VSUBS 0.006158f
C154 B.n99 VSUBS 0.006158f
C155 B.n100 VSUBS 0.006158f
C156 B.n101 VSUBS 0.006158f
C157 B.n102 VSUBS 0.006158f
C158 B.n103 VSUBS 0.006158f
C159 B.n104 VSUBS 0.006158f
C160 B.n105 VSUBS 0.006158f
C161 B.n106 VSUBS 0.006158f
C162 B.n107 VSUBS 0.006158f
C163 B.n108 VSUBS 0.006158f
C164 B.n109 VSUBS 0.006158f
C165 B.n110 VSUBS 0.006158f
C166 B.n111 VSUBS 0.006158f
C167 B.n112 VSUBS 0.006158f
C168 B.n113 VSUBS 0.006158f
C169 B.n114 VSUBS 0.006158f
C170 B.n115 VSUBS 0.006158f
C171 B.n116 VSUBS 0.006158f
C172 B.n117 VSUBS 0.006158f
C173 B.n118 VSUBS 0.015206f
C174 B.n119 VSUBS 0.015206f
C175 B.n120 VSUBS 0.015948f
C176 B.n121 VSUBS 0.006158f
C177 B.n122 VSUBS 0.006158f
C178 B.n123 VSUBS 0.006158f
C179 B.n124 VSUBS 0.006158f
C180 B.n125 VSUBS 0.006158f
C181 B.n126 VSUBS 0.006158f
C182 B.n127 VSUBS 0.006158f
C183 B.n128 VSUBS 0.006158f
C184 B.n129 VSUBS 0.006158f
C185 B.n130 VSUBS 0.006158f
C186 B.n131 VSUBS 0.006158f
C187 B.n132 VSUBS 0.006158f
C188 B.n133 VSUBS 0.006158f
C189 B.n134 VSUBS 0.006158f
C190 B.n135 VSUBS 0.006158f
C191 B.n136 VSUBS 0.006158f
C192 B.n137 VSUBS 0.006158f
C193 B.n138 VSUBS 0.006158f
C194 B.n139 VSUBS 0.006158f
C195 B.n140 VSUBS 0.006158f
C196 B.n141 VSUBS 0.006158f
C197 B.n142 VSUBS 0.006158f
C198 B.n143 VSUBS 0.006158f
C199 B.n144 VSUBS 0.006158f
C200 B.n145 VSUBS 0.006158f
C201 B.n146 VSUBS 0.006158f
C202 B.n147 VSUBS 0.006158f
C203 B.n148 VSUBS 0.006158f
C204 B.n149 VSUBS 0.006158f
C205 B.n150 VSUBS 0.006158f
C206 B.n151 VSUBS 0.006158f
C207 B.n152 VSUBS 0.006158f
C208 B.n153 VSUBS 0.006158f
C209 B.n154 VSUBS 0.006158f
C210 B.n155 VSUBS 0.006158f
C211 B.n156 VSUBS 0.006158f
C212 B.n157 VSUBS 0.006158f
C213 B.n158 VSUBS 0.006158f
C214 B.n159 VSUBS 0.006158f
C215 B.n160 VSUBS 0.006158f
C216 B.n161 VSUBS 0.006158f
C217 B.n162 VSUBS 0.004075f
C218 B.n163 VSUBS 0.014268f
C219 B.n164 VSUBS 0.005162f
C220 B.n165 VSUBS 0.006158f
C221 B.n166 VSUBS 0.006158f
C222 B.n167 VSUBS 0.006158f
C223 B.n168 VSUBS 0.006158f
C224 B.n169 VSUBS 0.006158f
C225 B.n170 VSUBS 0.006158f
C226 B.n171 VSUBS 0.006158f
C227 B.n172 VSUBS 0.006158f
C228 B.n173 VSUBS 0.006158f
C229 B.n174 VSUBS 0.006158f
C230 B.n175 VSUBS 0.006158f
C231 B.t11 VSUBS 0.205767f
C232 B.t10 VSUBS 0.212433f
C233 B.t9 VSUBS 0.178621f
C234 B.n176 VSUBS 0.085945f
C235 B.n177 VSUBS 0.055574f
C236 B.n178 VSUBS 0.014268f
C237 B.n179 VSUBS 0.005162f
C238 B.n180 VSUBS 0.006158f
C239 B.n181 VSUBS 0.006158f
C240 B.n182 VSUBS 0.006158f
C241 B.n183 VSUBS 0.006158f
C242 B.n184 VSUBS 0.006158f
C243 B.n185 VSUBS 0.006158f
C244 B.n186 VSUBS 0.006158f
C245 B.n187 VSUBS 0.006158f
C246 B.n188 VSUBS 0.006158f
C247 B.n189 VSUBS 0.006158f
C248 B.n190 VSUBS 0.006158f
C249 B.n191 VSUBS 0.006158f
C250 B.n192 VSUBS 0.006158f
C251 B.n193 VSUBS 0.006158f
C252 B.n194 VSUBS 0.006158f
C253 B.n195 VSUBS 0.006158f
C254 B.n196 VSUBS 0.006158f
C255 B.n197 VSUBS 0.006158f
C256 B.n198 VSUBS 0.006158f
C257 B.n199 VSUBS 0.006158f
C258 B.n200 VSUBS 0.006158f
C259 B.n201 VSUBS 0.006158f
C260 B.n202 VSUBS 0.006158f
C261 B.n203 VSUBS 0.006158f
C262 B.n204 VSUBS 0.006158f
C263 B.n205 VSUBS 0.006158f
C264 B.n206 VSUBS 0.006158f
C265 B.n207 VSUBS 0.006158f
C266 B.n208 VSUBS 0.006158f
C267 B.n209 VSUBS 0.006158f
C268 B.n210 VSUBS 0.006158f
C269 B.n211 VSUBS 0.006158f
C270 B.n212 VSUBS 0.006158f
C271 B.n213 VSUBS 0.006158f
C272 B.n214 VSUBS 0.006158f
C273 B.n215 VSUBS 0.006158f
C274 B.n216 VSUBS 0.006158f
C275 B.n217 VSUBS 0.006158f
C276 B.n218 VSUBS 0.006158f
C277 B.n219 VSUBS 0.006158f
C278 B.n220 VSUBS 0.006158f
C279 B.n221 VSUBS 0.006158f
C280 B.n222 VSUBS 0.006158f
C281 B.n223 VSUBS 0.015948f
C282 B.n224 VSUBS 0.015206f
C283 B.n225 VSUBS 0.015853f
C284 B.n226 VSUBS 0.006158f
C285 B.n227 VSUBS 0.006158f
C286 B.n228 VSUBS 0.006158f
C287 B.n229 VSUBS 0.006158f
C288 B.n230 VSUBS 0.006158f
C289 B.n231 VSUBS 0.006158f
C290 B.n232 VSUBS 0.006158f
C291 B.n233 VSUBS 0.006158f
C292 B.n234 VSUBS 0.006158f
C293 B.n235 VSUBS 0.006158f
C294 B.n236 VSUBS 0.006158f
C295 B.n237 VSUBS 0.006158f
C296 B.n238 VSUBS 0.006158f
C297 B.n239 VSUBS 0.006158f
C298 B.n240 VSUBS 0.006158f
C299 B.n241 VSUBS 0.006158f
C300 B.n242 VSUBS 0.006158f
C301 B.n243 VSUBS 0.006158f
C302 B.n244 VSUBS 0.006158f
C303 B.n245 VSUBS 0.006158f
C304 B.n246 VSUBS 0.006158f
C305 B.n247 VSUBS 0.006158f
C306 B.n248 VSUBS 0.006158f
C307 B.n249 VSUBS 0.006158f
C308 B.n250 VSUBS 0.006158f
C309 B.n251 VSUBS 0.006158f
C310 B.n252 VSUBS 0.006158f
C311 B.n253 VSUBS 0.006158f
C312 B.n254 VSUBS 0.006158f
C313 B.n255 VSUBS 0.006158f
C314 B.n256 VSUBS 0.006158f
C315 B.n257 VSUBS 0.006158f
C316 B.n258 VSUBS 0.006158f
C317 B.n259 VSUBS 0.006158f
C318 B.n260 VSUBS 0.006158f
C319 B.n261 VSUBS 0.006158f
C320 B.n262 VSUBS 0.006158f
C321 B.n263 VSUBS 0.006158f
C322 B.n264 VSUBS 0.006158f
C323 B.n265 VSUBS 0.015206f
C324 B.n266 VSUBS 0.015948f
C325 B.n267 VSUBS 0.015948f
C326 B.n268 VSUBS 0.006158f
C327 B.n269 VSUBS 0.006158f
C328 B.n270 VSUBS 0.006158f
C329 B.n271 VSUBS 0.006158f
C330 B.n272 VSUBS 0.006158f
C331 B.n273 VSUBS 0.006158f
C332 B.n274 VSUBS 0.006158f
C333 B.n275 VSUBS 0.006158f
C334 B.n276 VSUBS 0.006158f
C335 B.n277 VSUBS 0.006158f
C336 B.n278 VSUBS 0.006158f
C337 B.n279 VSUBS 0.006158f
C338 B.n280 VSUBS 0.006158f
C339 B.n281 VSUBS 0.006158f
C340 B.n282 VSUBS 0.006158f
C341 B.n283 VSUBS 0.006158f
C342 B.n284 VSUBS 0.006158f
C343 B.n285 VSUBS 0.006158f
C344 B.n286 VSUBS 0.006158f
C345 B.n287 VSUBS 0.006158f
C346 B.n288 VSUBS 0.006158f
C347 B.n289 VSUBS 0.006158f
C348 B.n290 VSUBS 0.006158f
C349 B.n291 VSUBS 0.006158f
C350 B.n292 VSUBS 0.006158f
C351 B.n293 VSUBS 0.006158f
C352 B.n294 VSUBS 0.006158f
C353 B.n295 VSUBS 0.006158f
C354 B.n296 VSUBS 0.006158f
C355 B.n297 VSUBS 0.006158f
C356 B.n298 VSUBS 0.006158f
C357 B.n299 VSUBS 0.006158f
C358 B.n300 VSUBS 0.006158f
C359 B.n301 VSUBS 0.006158f
C360 B.n302 VSUBS 0.006158f
C361 B.n303 VSUBS 0.006158f
C362 B.n304 VSUBS 0.006158f
C363 B.n305 VSUBS 0.006158f
C364 B.n306 VSUBS 0.006158f
C365 B.n307 VSUBS 0.006158f
C366 B.n308 VSUBS 0.006158f
C367 B.n309 VSUBS 0.004075f
C368 B.n310 VSUBS 0.014268f
C369 B.n311 VSUBS 0.005162f
C370 B.n312 VSUBS 0.006158f
C371 B.n313 VSUBS 0.006158f
C372 B.n314 VSUBS 0.006158f
C373 B.n315 VSUBS 0.006158f
C374 B.n316 VSUBS 0.006158f
C375 B.n317 VSUBS 0.006158f
C376 B.n318 VSUBS 0.006158f
C377 B.n319 VSUBS 0.006158f
C378 B.n320 VSUBS 0.006158f
C379 B.n321 VSUBS 0.006158f
C380 B.n322 VSUBS 0.006158f
C381 B.n323 VSUBS 0.005162f
C382 B.n324 VSUBS 0.014268f
C383 B.n325 VSUBS 0.004075f
C384 B.n326 VSUBS 0.006158f
C385 B.n327 VSUBS 0.006158f
C386 B.n328 VSUBS 0.006158f
C387 B.n329 VSUBS 0.006158f
C388 B.n330 VSUBS 0.006158f
C389 B.n331 VSUBS 0.006158f
C390 B.n332 VSUBS 0.006158f
C391 B.n333 VSUBS 0.006158f
C392 B.n334 VSUBS 0.006158f
C393 B.n335 VSUBS 0.006158f
C394 B.n336 VSUBS 0.006158f
C395 B.n337 VSUBS 0.006158f
C396 B.n338 VSUBS 0.006158f
C397 B.n339 VSUBS 0.006158f
C398 B.n340 VSUBS 0.006158f
C399 B.n341 VSUBS 0.006158f
C400 B.n342 VSUBS 0.006158f
C401 B.n343 VSUBS 0.006158f
C402 B.n344 VSUBS 0.006158f
C403 B.n345 VSUBS 0.006158f
C404 B.n346 VSUBS 0.006158f
C405 B.n347 VSUBS 0.006158f
C406 B.n348 VSUBS 0.006158f
C407 B.n349 VSUBS 0.006158f
C408 B.n350 VSUBS 0.006158f
C409 B.n351 VSUBS 0.006158f
C410 B.n352 VSUBS 0.006158f
C411 B.n353 VSUBS 0.006158f
C412 B.n354 VSUBS 0.006158f
C413 B.n355 VSUBS 0.006158f
C414 B.n356 VSUBS 0.006158f
C415 B.n357 VSUBS 0.006158f
C416 B.n358 VSUBS 0.006158f
C417 B.n359 VSUBS 0.006158f
C418 B.n360 VSUBS 0.006158f
C419 B.n361 VSUBS 0.006158f
C420 B.n362 VSUBS 0.006158f
C421 B.n363 VSUBS 0.006158f
C422 B.n364 VSUBS 0.006158f
C423 B.n365 VSUBS 0.006158f
C424 B.n366 VSUBS 0.006158f
C425 B.n367 VSUBS 0.015948f
C426 B.n368 VSUBS 0.015948f
C427 B.n369 VSUBS 0.015206f
C428 B.n370 VSUBS 0.006158f
C429 B.n371 VSUBS 0.006158f
C430 B.n372 VSUBS 0.006158f
C431 B.n373 VSUBS 0.006158f
C432 B.n374 VSUBS 0.006158f
C433 B.n375 VSUBS 0.006158f
C434 B.n376 VSUBS 0.006158f
C435 B.n377 VSUBS 0.006158f
C436 B.n378 VSUBS 0.006158f
C437 B.n379 VSUBS 0.006158f
C438 B.n380 VSUBS 0.006158f
C439 B.n381 VSUBS 0.006158f
C440 B.n382 VSUBS 0.006158f
C441 B.n383 VSUBS 0.006158f
C442 B.n384 VSUBS 0.006158f
C443 B.n385 VSUBS 0.006158f
C444 B.n386 VSUBS 0.006158f
C445 B.n387 VSUBS 0.008036f
C446 B.n388 VSUBS 0.008561f
C447 B.n389 VSUBS 0.017024f
.ends

