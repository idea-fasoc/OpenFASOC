* NGSPICE file created from diff_pair_sample_0910.ext - technology: sky130A

.subckt diff_pair_sample_0910 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t17 VN.t0 VDD2.t9 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X1 VDD1.t9 VP.t0 VTAIL.t2 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X2 VDD1.t8 VP.t1 VTAIL.t6 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=3.06735 ps=18.92 w=18.59 l=3.7
X3 B.t11 B.t9 B.t10 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=0 ps=0 w=18.59 l=3.7
X4 VTAIL.t16 VN.t1 VDD2.t8 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X5 VDD1.t7 VP.t2 VTAIL.t5 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=7.2501 ps=37.96 w=18.59 l=3.7
X6 VDD1.t6 VP.t3 VTAIL.t19 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=3.06735 ps=18.92 w=18.59 l=3.7
X7 VDD1.t5 VP.t4 VTAIL.t7 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=7.2501 ps=37.96 w=18.59 l=3.7
X8 B.t8 B.t6 B.t7 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=0 ps=0 w=18.59 l=3.7
X9 VDD2.t5 VN.t2 VTAIL.t15 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=7.2501 ps=37.96 w=18.59 l=3.7
X10 VTAIL.t14 VN.t3 VDD2.t4 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X11 VDD2.t3 VN.t4 VTAIL.t13 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=7.2501 ps=37.96 w=18.59 l=3.7
X12 VDD2.t2 VN.t5 VTAIL.t12 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X13 B.t5 B.t3 B.t4 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=0 ps=0 w=18.59 l=3.7
X14 B.t2 B.t0 B.t1 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=0 ps=0 w=18.59 l=3.7
X15 VTAIL.t18 VP.t5 VDD1.t4 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X16 VDD2.t1 VN.t6 VTAIL.t11 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=3.06735 ps=18.92 w=18.59 l=3.7
X17 VTAIL.t0 VP.t6 VDD1.t3 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X18 VDD1.t2 VP.t7 VTAIL.t4 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X19 VTAIL.t3 VP.t8 VDD1.t1 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X20 VDD2.t0 VN.t7 VTAIL.t10 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X21 VTAIL.t9 VN.t8 VDD2.t7 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X22 VTAIL.t1 VP.t9 VDD1.t0 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=3.06735 pd=18.92 as=3.06735 ps=18.92 w=18.59 l=3.7
X23 VDD2.t6 VN.t9 VTAIL.t8 w_n5806_n4686# sky130_fd_pr__pfet_01v8 ad=7.2501 pd=37.96 as=3.06735 ps=18.92 w=18.59 l=3.7
R0 VN.n108 VN.n107 161.3
R1 VN.n106 VN.n56 161.3
R2 VN.n105 VN.n104 161.3
R3 VN.n103 VN.n57 161.3
R4 VN.n102 VN.n101 161.3
R5 VN.n100 VN.n58 161.3
R6 VN.n99 VN.n98 161.3
R7 VN.n97 VN.n59 161.3
R8 VN.n96 VN.n95 161.3
R9 VN.n94 VN.n60 161.3
R10 VN.n93 VN.n92 161.3
R11 VN.n91 VN.n62 161.3
R12 VN.n90 VN.n89 161.3
R13 VN.n88 VN.n63 161.3
R14 VN.n87 VN.n86 161.3
R15 VN.n85 VN.n64 161.3
R16 VN.n84 VN.n83 161.3
R17 VN.n82 VN.n65 161.3
R18 VN.n81 VN.n80 161.3
R19 VN.n79 VN.n66 161.3
R20 VN.n78 VN.n77 161.3
R21 VN.n76 VN.n67 161.3
R22 VN.n75 VN.n74 161.3
R23 VN.n73 VN.n68 161.3
R24 VN.n72 VN.n71 161.3
R25 VN.n53 VN.n52 161.3
R26 VN.n51 VN.n1 161.3
R27 VN.n50 VN.n49 161.3
R28 VN.n48 VN.n2 161.3
R29 VN.n47 VN.n46 161.3
R30 VN.n45 VN.n3 161.3
R31 VN.n44 VN.n43 161.3
R32 VN.n42 VN.n4 161.3
R33 VN.n41 VN.n40 161.3
R34 VN.n38 VN.n5 161.3
R35 VN.n37 VN.n36 161.3
R36 VN.n35 VN.n6 161.3
R37 VN.n34 VN.n33 161.3
R38 VN.n32 VN.n7 161.3
R39 VN.n31 VN.n30 161.3
R40 VN.n29 VN.n8 161.3
R41 VN.n28 VN.n27 161.3
R42 VN.n26 VN.n9 161.3
R43 VN.n25 VN.n24 161.3
R44 VN.n23 VN.n10 161.3
R45 VN.n22 VN.n21 161.3
R46 VN.n20 VN.n11 161.3
R47 VN.n19 VN.n18 161.3
R48 VN.n17 VN.n12 161.3
R49 VN.n16 VN.n15 161.3
R50 VN.n69 VN.t4 152.959
R51 VN.n13 VN.t9 152.959
R52 VN.n27 VN.t5 121.087
R53 VN.n14 VN.t3 121.087
R54 VN.n39 VN.t8 121.087
R55 VN.n0 VN.t2 121.087
R56 VN.n83 VN.t7 121.087
R57 VN.n70 VN.t0 121.087
R58 VN.n61 VN.t1 121.087
R59 VN.n55 VN.t6 121.087
R60 VN.n54 VN.n0 87.1314
R61 VN.n109 VN.n55 87.1314
R62 VN.n14 VN.n13 73.4859
R63 VN.n70 VN.n69 73.4859
R64 VN VN.n109 64.2821
R65 VN.n46 VN.n2 44.8641
R66 VN.n101 VN.n57 44.8641
R67 VN.n21 VN.n20 41.9503
R68 VN.n33 VN.n6 41.9503
R69 VN.n77 VN.n76 41.9503
R70 VN.n89 VN.n62 41.9503
R71 VN.n21 VN.n10 39.0365
R72 VN.n33 VN.n32 39.0365
R73 VN.n77 VN.n66 39.0365
R74 VN.n89 VN.n88 39.0365
R75 VN.n46 VN.n45 36.1227
R76 VN.n101 VN.n100 36.1227
R77 VN.n15 VN.n12 24.4675
R78 VN.n19 VN.n12 24.4675
R79 VN.n20 VN.n19 24.4675
R80 VN.n25 VN.n10 24.4675
R81 VN.n26 VN.n25 24.4675
R82 VN.n27 VN.n26 24.4675
R83 VN.n27 VN.n8 24.4675
R84 VN.n31 VN.n8 24.4675
R85 VN.n32 VN.n31 24.4675
R86 VN.n37 VN.n6 24.4675
R87 VN.n38 VN.n37 24.4675
R88 VN.n40 VN.n38 24.4675
R89 VN.n44 VN.n4 24.4675
R90 VN.n45 VN.n44 24.4675
R91 VN.n50 VN.n2 24.4675
R92 VN.n51 VN.n50 24.4675
R93 VN.n52 VN.n51 24.4675
R94 VN.n76 VN.n75 24.4675
R95 VN.n75 VN.n68 24.4675
R96 VN.n71 VN.n68 24.4675
R97 VN.n88 VN.n87 24.4675
R98 VN.n87 VN.n64 24.4675
R99 VN.n83 VN.n64 24.4675
R100 VN.n83 VN.n82 24.4675
R101 VN.n82 VN.n81 24.4675
R102 VN.n81 VN.n66 24.4675
R103 VN.n100 VN.n99 24.4675
R104 VN.n99 VN.n59 24.4675
R105 VN.n95 VN.n94 24.4675
R106 VN.n94 VN.n93 24.4675
R107 VN.n93 VN.n62 24.4675
R108 VN.n107 VN.n106 24.4675
R109 VN.n106 VN.n105 24.4675
R110 VN.n105 VN.n57 24.4675
R111 VN.n39 VN.n4 22.9995
R112 VN.n61 VN.n59 22.9995
R113 VN.n72 VN.n69 3.37703
R114 VN.n16 VN.n13 3.37703
R115 VN.n52 VN.n0 2.93654
R116 VN.n107 VN.n55 2.93654
R117 VN.n15 VN.n14 1.46852
R118 VN.n40 VN.n39 1.46852
R119 VN.n71 VN.n70 1.46852
R120 VN.n95 VN.n61 1.46852
R121 VN.n109 VN.n108 0.354971
R122 VN.n54 VN.n53 0.354971
R123 VN VN.n54 0.26696
R124 VN.n108 VN.n56 0.189894
R125 VN.n104 VN.n56 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n102 0.189894
R128 VN.n102 VN.n58 0.189894
R129 VN.n98 VN.n58 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n96 0.189894
R132 VN.n96 VN.n60 0.189894
R133 VN.n92 VN.n60 0.189894
R134 VN.n92 VN.n91 0.189894
R135 VN.n91 VN.n90 0.189894
R136 VN.n90 VN.n63 0.189894
R137 VN.n86 VN.n63 0.189894
R138 VN.n86 VN.n85 0.189894
R139 VN.n85 VN.n84 0.189894
R140 VN.n84 VN.n65 0.189894
R141 VN.n80 VN.n65 0.189894
R142 VN.n80 VN.n79 0.189894
R143 VN.n79 VN.n78 0.189894
R144 VN.n78 VN.n67 0.189894
R145 VN.n74 VN.n67 0.189894
R146 VN.n74 VN.n73 0.189894
R147 VN.n73 VN.n72 0.189894
R148 VN.n17 VN.n16 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n18 VN.n11 0.189894
R151 VN.n22 VN.n11 0.189894
R152 VN.n23 VN.n22 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n24 VN.n9 0.189894
R155 VN.n28 VN.n9 0.189894
R156 VN.n29 VN.n28 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n30 VN.n7 0.189894
R159 VN.n34 VN.n7 0.189894
R160 VN.n35 VN.n34 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n36 VN.n5 0.189894
R163 VN.n41 VN.n5 0.189894
R164 VN.n42 VN.n41 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n43 VN.n3 0.189894
R167 VN.n47 VN.n3 0.189894
R168 VN.n48 VN.n47 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n49 VN.n1 0.189894
R171 VN.n53 VN.n1 0.189894
R172 VDD2.n1 VDD2.t6 73.5611
R173 VDD2.n3 VDD2.n2 70.8886
R174 VDD2 VDD2.n7 70.8858
R175 VDD2.n4 VDD2.t1 70.0871
R176 VDD2.n6 VDD2.n5 68.3386
R177 VDD2.n1 VDD2.n0 68.3383
R178 VDD2.n4 VDD2.n3 56.2433
R179 VDD2.n6 VDD2.n4 3.47464
R180 VDD2.n7 VDD2.t9 1.74902
R181 VDD2.n7 VDD2.t3 1.74902
R182 VDD2.n5 VDD2.t8 1.74902
R183 VDD2.n5 VDD2.t0 1.74902
R184 VDD2.n2 VDD2.t7 1.74902
R185 VDD2.n2 VDD2.t5 1.74902
R186 VDD2.n0 VDD2.t4 1.74902
R187 VDD2.n0 VDD2.t2 1.74902
R188 VDD2 VDD2.n6 0.927224
R189 VDD2.n3 VDD2.n1 0.813688
R190 VTAIL.n11 VTAIL.t13 53.4083
R191 VTAIL.n16 VTAIL.t7 53.4081
R192 VTAIL.n17 VTAIL.t15 53.4081
R193 VTAIL.n2 VTAIL.t5 53.4081
R194 VTAIL.n15 VTAIL.n14 51.6598
R195 VTAIL.n13 VTAIL.n12 51.6598
R196 VTAIL.n10 VTAIL.n9 51.6598
R197 VTAIL.n8 VTAIL.n7 51.6598
R198 VTAIL.n19 VTAIL.n18 51.6596
R199 VTAIL.n1 VTAIL.n0 51.6596
R200 VTAIL.n4 VTAIL.n3 51.6596
R201 VTAIL.n6 VTAIL.n5 51.6596
R202 VTAIL.n8 VTAIL.n6 35.341
R203 VTAIL.n17 VTAIL.n16 31.8669
R204 VTAIL.n10 VTAIL.n8 3.47464
R205 VTAIL.n11 VTAIL.n10 3.47464
R206 VTAIL.n15 VTAIL.n13 3.47464
R207 VTAIL.n16 VTAIL.n15 3.47464
R208 VTAIL.n6 VTAIL.n4 3.47464
R209 VTAIL.n4 VTAIL.n2 3.47464
R210 VTAIL.n19 VTAIL.n17 3.47464
R211 VTAIL VTAIL.n1 2.66429
R212 VTAIL.n13 VTAIL.n11 2.2074
R213 VTAIL.n2 VTAIL.n1 2.2074
R214 VTAIL.n18 VTAIL.t12 1.74902
R215 VTAIL.n18 VTAIL.t9 1.74902
R216 VTAIL.n0 VTAIL.t8 1.74902
R217 VTAIL.n0 VTAIL.t14 1.74902
R218 VTAIL.n3 VTAIL.t4 1.74902
R219 VTAIL.n3 VTAIL.t0 1.74902
R220 VTAIL.n5 VTAIL.t19 1.74902
R221 VTAIL.n5 VTAIL.t1 1.74902
R222 VTAIL.n14 VTAIL.t2 1.74902
R223 VTAIL.n14 VTAIL.t18 1.74902
R224 VTAIL.n12 VTAIL.t6 1.74902
R225 VTAIL.n12 VTAIL.t3 1.74902
R226 VTAIL.n9 VTAIL.t10 1.74902
R227 VTAIL.n9 VTAIL.t17 1.74902
R228 VTAIL.n7 VTAIL.t11 1.74902
R229 VTAIL.n7 VTAIL.t16 1.74902
R230 VTAIL VTAIL.n19 0.810845
R231 VP.n33 VP.n32 161.3
R232 VP.n34 VP.n29 161.3
R233 VP.n36 VP.n35 161.3
R234 VP.n37 VP.n28 161.3
R235 VP.n39 VP.n38 161.3
R236 VP.n40 VP.n27 161.3
R237 VP.n42 VP.n41 161.3
R238 VP.n43 VP.n26 161.3
R239 VP.n45 VP.n44 161.3
R240 VP.n46 VP.n25 161.3
R241 VP.n48 VP.n47 161.3
R242 VP.n49 VP.n24 161.3
R243 VP.n51 VP.n50 161.3
R244 VP.n52 VP.n23 161.3
R245 VP.n54 VP.n53 161.3
R246 VP.n55 VP.n22 161.3
R247 VP.n58 VP.n57 161.3
R248 VP.n59 VP.n21 161.3
R249 VP.n61 VP.n60 161.3
R250 VP.n62 VP.n20 161.3
R251 VP.n64 VP.n63 161.3
R252 VP.n65 VP.n19 161.3
R253 VP.n67 VP.n66 161.3
R254 VP.n68 VP.n18 161.3
R255 VP.n70 VP.n69 161.3
R256 VP.n125 VP.n124 161.3
R257 VP.n123 VP.n1 161.3
R258 VP.n122 VP.n121 161.3
R259 VP.n120 VP.n2 161.3
R260 VP.n119 VP.n118 161.3
R261 VP.n117 VP.n3 161.3
R262 VP.n116 VP.n115 161.3
R263 VP.n114 VP.n4 161.3
R264 VP.n113 VP.n112 161.3
R265 VP.n110 VP.n5 161.3
R266 VP.n109 VP.n108 161.3
R267 VP.n107 VP.n6 161.3
R268 VP.n106 VP.n105 161.3
R269 VP.n104 VP.n7 161.3
R270 VP.n103 VP.n102 161.3
R271 VP.n101 VP.n8 161.3
R272 VP.n100 VP.n99 161.3
R273 VP.n98 VP.n9 161.3
R274 VP.n97 VP.n96 161.3
R275 VP.n95 VP.n10 161.3
R276 VP.n94 VP.n93 161.3
R277 VP.n92 VP.n11 161.3
R278 VP.n91 VP.n90 161.3
R279 VP.n89 VP.n12 161.3
R280 VP.n88 VP.n87 161.3
R281 VP.n85 VP.n13 161.3
R282 VP.n84 VP.n83 161.3
R283 VP.n82 VP.n14 161.3
R284 VP.n81 VP.n80 161.3
R285 VP.n79 VP.n15 161.3
R286 VP.n78 VP.n77 161.3
R287 VP.n76 VP.n16 161.3
R288 VP.n75 VP.n74 161.3
R289 VP.n30 VP.t1 152.959
R290 VP.n99 VP.t7 121.087
R291 VP.n73 VP.t3 121.087
R292 VP.n86 VP.t9 121.087
R293 VP.n111 VP.t6 121.087
R294 VP.n0 VP.t2 121.087
R295 VP.n44 VP.t0 121.087
R296 VP.n17 VP.t4 121.087
R297 VP.n56 VP.t5 121.087
R298 VP.n31 VP.t8 121.087
R299 VP.n73 VP.n72 87.1314
R300 VP.n126 VP.n0 87.1314
R301 VP.n71 VP.n17 87.1314
R302 VP.n31 VP.n30 73.4859
R303 VP.n72 VP.n71 64.1168
R304 VP.n80 VP.n79 44.8641
R305 VP.n118 VP.n2 44.8641
R306 VP.n63 VP.n19 44.8641
R307 VP.n93 VP.n92 41.9503
R308 VP.n105 VP.n6 41.9503
R309 VP.n50 VP.n23 41.9503
R310 VP.n38 VP.n37 41.9503
R311 VP.n93 VP.n10 39.0365
R312 VP.n105 VP.n104 39.0365
R313 VP.n50 VP.n49 39.0365
R314 VP.n38 VP.n27 39.0365
R315 VP.n80 VP.n14 36.1227
R316 VP.n118 VP.n117 36.1227
R317 VP.n63 VP.n62 36.1227
R318 VP.n74 VP.n16 24.4675
R319 VP.n78 VP.n16 24.4675
R320 VP.n79 VP.n78 24.4675
R321 VP.n84 VP.n14 24.4675
R322 VP.n85 VP.n84 24.4675
R323 VP.n87 VP.n12 24.4675
R324 VP.n91 VP.n12 24.4675
R325 VP.n92 VP.n91 24.4675
R326 VP.n97 VP.n10 24.4675
R327 VP.n98 VP.n97 24.4675
R328 VP.n99 VP.n98 24.4675
R329 VP.n99 VP.n8 24.4675
R330 VP.n103 VP.n8 24.4675
R331 VP.n104 VP.n103 24.4675
R332 VP.n109 VP.n6 24.4675
R333 VP.n110 VP.n109 24.4675
R334 VP.n112 VP.n110 24.4675
R335 VP.n116 VP.n4 24.4675
R336 VP.n117 VP.n116 24.4675
R337 VP.n122 VP.n2 24.4675
R338 VP.n123 VP.n122 24.4675
R339 VP.n124 VP.n123 24.4675
R340 VP.n67 VP.n19 24.4675
R341 VP.n68 VP.n67 24.4675
R342 VP.n69 VP.n68 24.4675
R343 VP.n54 VP.n23 24.4675
R344 VP.n55 VP.n54 24.4675
R345 VP.n57 VP.n55 24.4675
R346 VP.n61 VP.n21 24.4675
R347 VP.n62 VP.n61 24.4675
R348 VP.n42 VP.n27 24.4675
R349 VP.n43 VP.n42 24.4675
R350 VP.n44 VP.n43 24.4675
R351 VP.n44 VP.n25 24.4675
R352 VP.n48 VP.n25 24.4675
R353 VP.n49 VP.n48 24.4675
R354 VP.n32 VP.n29 24.4675
R355 VP.n36 VP.n29 24.4675
R356 VP.n37 VP.n36 24.4675
R357 VP.n86 VP.n85 22.9995
R358 VP.n111 VP.n4 22.9995
R359 VP.n56 VP.n21 22.9995
R360 VP.n33 VP.n30 3.37702
R361 VP.n74 VP.n73 2.93654
R362 VP.n124 VP.n0 2.93654
R363 VP.n69 VP.n17 2.93654
R364 VP.n87 VP.n86 1.46852
R365 VP.n112 VP.n111 1.46852
R366 VP.n57 VP.n56 1.46852
R367 VP.n32 VP.n31 1.46852
R368 VP.n71 VP.n70 0.354971
R369 VP.n75 VP.n72 0.354971
R370 VP.n126 VP.n125 0.354971
R371 VP VP.n126 0.26696
R372 VP.n34 VP.n33 0.189894
R373 VP.n35 VP.n34 0.189894
R374 VP.n35 VP.n28 0.189894
R375 VP.n39 VP.n28 0.189894
R376 VP.n40 VP.n39 0.189894
R377 VP.n41 VP.n40 0.189894
R378 VP.n41 VP.n26 0.189894
R379 VP.n45 VP.n26 0.189894
R380 VP.n46 VP.n45 0.189894
R381 VP.n47 VP.n46 0.189894
R382 VP.n47 VP.n24 0.189894
R383 VP.n51 VP.n24 0.189894
R384 VP.n52 VP.n51 0.189894
R385 VP.n53 VP.n52 0.189894
R386 VP.n53 VP.n22 0.189894
R387 VP.n58 VP.n22 0.189894
R388 VP.n59 VP.n58 0.189894
R389 VP.n60 VP.n59 0.189894
R390 VP.n60 VP.n20 0.189894
R391 VP.n64 VP.n20 0.189894
R392 VP.n65 VP.n64 0.189894
R393 VP.n66 VP.n65 0.189894
R394 VP.n66 VP.n18 0.189894
R395 VP.n70 VP.n18 0.189894
R396 VP.n76 VP.n75 0.189894
R397 VP.n77 VP.n76 0.189894
R398 VP.n77 VP.n15 0.189894
R399 VP.n81 VP.n15 0.189894
R400 VP.n82 VP.n81 0.189894
R401 VP.n83 VP.n82 0.189894
R402 VP.n83 VP.n13 0.189894
R403 VP.n88 VP.n13 0.189894
R404 VP.n89 VP.n88 0.189894
R405 VP.n90 VP.n89 0.189894
R406 VP.n90 VP.n11 0.189894
R407 VP.n94 VP.n11 0.189894
R408 VP.n95 VP.n94 0.189894
R409 VP.n96 VP.n95 0.189894
R410 VP.n96 VP.n9 0.189894
R411 VP.n100 VP.n9 0.189894
R412 VP.n101 VP.n100 0.189894
R413 VP.n102 VP.n101 0.189894
R414 VP.n102 VP.n7 0.189894
R415 VP.n106 VP.n7 0.189894
R416 VP.n107 VP.n106 0.189894
R417 VP.n108 VP.n107 0.189894
R418 VP.n108 VP.n5 0.189894
R419 VP.n113 VP.n5 0.189894
R420 VP.n114 VP.n113 0.189894
R421 VP.n115 VP.n114 0.189894
R422 VP.n115 VP.n3 0.189894
R423 VP.n119 VP.n3 0.189894
R424 VP.n120 VP.n119 0.189894
R425 VP.n121 VP.n120 0.189894
R426 VP.n121 VP.n1 0.189894
R427 VP.n125 VP.n1 0.189894
R428 VDD1.n1 VDD1.t8 73.5612
R429 VDD1.n3 VDD1.t6 73.5611
R430 VDD1.n5 VDD1.n4 70.8886
R431 VDD1.n1 VDD1.n0 68.3386
R432 VDD1.n7 VDD1.n6 68.3384
R433 VDD1.n3 VDD1.n2 68.3383
R434 VDD1.n7 VDD1.n5 58.5634
R435 VDD1 VDD1.n7 2.54791
R436 VDD1.n6 VDD1.t4 1.74902
R437 VDD1.n6 VDD1.t5 1.74902
R438 VDD1.n0 VDD1.t1 1.74902
R439 VDD1.n0 VDD1.t9 1.74902
R440 VDD1.n4 VDD1.t3 1.74902
R441 VDD1.n4 VDD1.t7 1.74902
R442 VDD1.n2 VDD1.t0 1.74902
R443 VDD1.n2 VDD1.t2 1.74902
R444 VDD1 VDD1.n1 0.927224
R445 VDD1.n5 VDD1.n3 0.813688
R446 B.n857 B.n856 585
R447 B.n858 B.n111 585
R448 B.n860 B.n859 585
R449 B.n861 B.n110 585
R450 B.n863 B.n862 585
R451 B.n864 B.n109 585
R452 B.n866 B.n865 585
R453 B.n867 B.n108 585
R454 B.n869 B.n868 585
R455 B.n870 B.n107 585
R456 B.n872 B.n871 585
R457 B.n873 B.n106 585
R458 B.n875 B.n874 585
R459 B.n876 B.n105 585
R460 B.n878 B.n877 585
R461 B.n879 B.n104 585
R462 B.n881 B.n880 585
R463 B.n882 B.n103 585
R464 B.n884 B.n883 585
R465 B.n885 B.n102 585
R466 B.n887 B.n886 585
R467 B.n888 B.n101 585
R468 B.n890 B.n889 585
R469 B.n891 B.n100 585
R470 B.n893 B.n892 585
R471 B.n894 B.n99 585
R472 B.n896 B.n895 585
R473 B.n897 B.n98 585
R474 B.n899 B.n898 585
R475 B.n900 B.n97 585
R476 B.n902 B.n901 585
R477 B.n903 B.n96 585
R478 B.n905 B.n904 585
R479 B.n906 B.n95 585
R480 B.n908 B.n907 585
R481 B.n909 B.n94 585
R482 B.n911 B.n910 585
R483 B.n912 B.n93 585
R484 B.n914 B.n913 585
R485 B.n915 B.n92 585
R486 B.n917 B.n916 585
R487 B.n918 B.n91 585
R488 B.n920 B.n919 585
R489 B.n921 B.n90 585
R490 B.n923 B.n922 585
R491 B.n924 B.n89 585
R492 B.n926 B.n925 585
R493 B.n927 B.n88 585
R494 B.n929 B.n928 585
R495 B.n930 B.n87 585
R496 B.n932 B.n931 585
R497 B.n933 B.n86 585
R498 B.n935 B.n934 585
R499 B.n936 B.n85 585
R500 B.n938 B.n937 585
R501 B.n939 B.n84 585
R502 B.n941 B.n940 585
R503 B.n942 B.n83 585
R504 B.n944 B.n943 585
R505 B.n945 B.n82 585
R506 B.n947 B.n946 585
R507 B.n949 B.n79 585
R508 B.n951 B.n950 585
R509 B.n952 B.n78 585
R510 B.n954 B.n953 585
R511 B.n955 B.n77 585
R512 B.n957 B.n956 585
R513 B.n958 B.n76 585
R514 B.n960 B.n959 585
R515 B.n961 B.n75 585
R516 B.n963 B.n962 585
R517 B.n965 B.n964 585
R518 B.n966 B.n71 585
R519 B.n968 B.n967 585
R520 B.n969 B.n70 585
R521 B.n971 B.n970 585
R522 B.n972 B.n69 585
R523 B.n974 B.n973 585
R524 B.n975 B.n68 585
R525 B.n977 B.n976 585
R526 B.n978 B.n67 585
R527 B.n980 B.n979 585
R528 B.n981 B.n66 585
R529 B.n983 B.n982 585
R530 B.n984 B.n65 585
R531 B.n986 B.n985 585
R532 B.n987 B.n64 585
R533 B.n989 B.n988 585
R534 B.n990 B.n63 585
R535 B.n992 B.n991 585
R536 B.n993 B.n62 585
R537 B.n995 B.n994 585
R538 B.n996 B.n61 585
R539 B.n998 B.n997 585
R540 B.n999 B.n60 585
R541 B.n1001 B.n1000 585
R542 B.n1002 B.n59 585
R543 B.n1004 B.n1003 585
R544 B.n1005 B.n58 585
R545 B.n1007 B.n1006 585
R546 B.n1008 B.n57 585
R547 B.n1010 B.n1009 585
R548 B.n1011 B.n56 585
R549 B.n1013 B.n1012 585
R550 B.n1014 B.n55 585
R551 B.n1016 B.n1015 585
R552 B.n1017 B.n54 585
R553 B.n1019 B.n1018 585
R554 B.n1020 B.n53 585
R555 B.n1022 B.n1021 585
R556 B.n1023 B.n52 585
R557 B.n1025 B.n1024 585
R558 B.n1026 B.n51 585
R559 B.n1028 B.n1027 585
R560 B.n1029 B.n50 585
R561 B.n1031 B.n1030 585
R562 B.n1032 B.n49 585
R563 B.n1034 B.n1033 585
R564 B.n1035 B.n48 585
R565 B.n1037 B.n1036 585
R566 B.n1038 B.n47 585
R567 B.n1040 B.n1039 585
R568 B.n1041 B.n46 585
R569 B.n1043 B.n1042 585
R570 B.n1044 B.n45 585
R571 B.n1046 B.n1045 585
R572 B.n1047 B.n44 585
R573 B.n1049 B.n1048 585
R574 B.n1050 B.n43 585
R575 B.n1052 B.n1051 585
R576 B.n1053 B.n42 585
R577 B.n1055 B.n1054 585
R578 B.n855 B.n112 585
R579 B.n854 B.n853 585
R580 B.n852 B.n113 585
R581 B.n851 B.n850 585
R582 B.n849 B.n114 585
R583 B.n848 B.n847 585
R584 B.n846 B.n115 585
R585 B.n845 B.n844 585
R586 B.n843 B.n116 585
R587 B.n842 B.n841 585
R588 B.n840 B.n117 585
R589 B.n839 B.n838 585
R590 B.n837 B.n118 585
R591 B.n836 B.n835 585
R592 B.n834 B.n119 585
R593 B.n833 B.n832 585
R594 B.n831 B.n120 585
R595 B.n830 B.n829 585
R596 B.n828 B.n121 585
R597 B.n827 B.n826 585
R598 B.n825 B.n122 585
R599 B.n824 B.n823 585
R600 B.n822 B.n123 585
R601 B.n821 B.n820 585
R602 B.n819 B.n124 585
R603 B.n818 B.n817 585
R604 B.n816 B.n125 585
R605 B.n815 B.n814 585
R606 B.n813 B.n126 585
R607 B.n812 B.n811 585
R608 B.n810 B.n127 585
R609 B.n809 B.n808 585
R610 B.n807 B.n128 585
R611 B.n806 B.n805 585
R612 B.n804 B.n129 585
R613 B.n803 B.n802 585
R614 B.n801 B.n130 585
R615 B.n800 B.n799 585
R616 B.n798 B.n131 585
R617 B.n797 B.n796 585
R618 B.n795 B.n132 585
R619 B.n794 B.n793 585
R620 B.n792 B.n133 585
R621 B.n791 B.n790 585
R622 B.n789 B.n134 585
R623 B.n788 B.n787 585
R624 B.n786 B.n135 585
R625 B.n785 B.n784 585
R626 B.n783 B.n136 585
R627 B.n782 B.n781 585
R628 B.n780 B.n137 585
R629 B.n779 B.n778 585
R630 B.n777 B.n138 585
R631 B.n776 B.n775 585
R632 B.n774 B.n139 585
R633 B.n773 B.n772 585
R634 B.n771 B.n140 585
R635 B.n770 B.n769 585
R636 B.n768 B.n141 585
R637 B.n767 B.n766 585
R638 B.n765 B.n142 585
R639 B.n764 B.n763 585
R640 B.n762 B.n143 585
R641 B.n761 B.n760 585
R642 B.n759 B.n144 585
R643 B.n758 B.n757 585
R644 B.n756 B.n145 585
R645 B.n755 B.n754 585
R646 B.n753 B.n146 585
R647 B.n752 B.n751 585
R648 B.n750 B.n147 585
R649 B.n749 B.n748 585
R650 B.n747 B.n148 585
R651 B.n746 B.n745 585
R652 B.n744 B.n149 585
R653 B.n743 B.n742 585
R654 B.n741 B.n150 585
R655 B.n740 B.n739 585
R656 B.n738 B.n151 585
R657 B.n737 B.n736 585
R658 B.n735 B.n152 585
R659 B.n734 B.n733 585
R660 B.n732 B.n153 585
R661 B.n731 B.n730 585
R662 B.n729 B.n154 585
R663 B.n728 B.n727 585
R664 B.n726 B.n155 585
R665 B.n725 B.n724 585
R666 B.n723 B.n156 585
R667 B.n722 B.n721 585
R668 B.n720 B.n157 585
R669 B.n719 B.n718 585
R670 B.n717 B.n158 585
R671 B.n716 B.n715 585
R672 B.n714 B.n159 585
R673 B.n713 B.n712 585
R674 B.n711 B.n160 585
R675 B.n710 B.n709 585
R676 B.n708 B.n161 585
R677 B.n707 B.n706 585
R678 B.n705 B.n162 585
R679 B.n704 B.n703 585
R680 B.n702 B.n163 585
R681 B.n701 B.n700 585
R682 B.n699 B.n164 585
R683 B.n698 B.n697 585
R684 B.n696 B.n165 585
R685 B.n695 B.n694 585
R686 B.n693 B.n166 585
R687 B.n692 B.n691 585
R688 B.n690 B.n167 585
R689 B.n689 B.n688 585
R690 B.n687 B.n168 585
R691 B.n686 B.n685 585
R692 B.n684 B.n169 585
R693 B.n683 B.n682 585
R694 B.n681 B.n170 585
R695 B.n680 B.n679 585
R696 B.n678 B.n171 585
R697 B.n677 B.n676 585
R698 B.n675 B.n172 585
R699 B.n674 B.n673 585
R700 B.n672 B.n173 585
R701 B.n671 B.n670 585
R702 B.n669 B.n174 585
R703 B.n668 B.n667 585
R704 B.n666 B.n175 585
R705 B.n665 B.n664 585
R706 B.n663 B.n176 585
R707 B.n662 B.n661 585
R708 B.n660 B.n177 585
R709 B.n659 B.n658 585
R710 B.n657 B.n178 585
R711 B.n656 B.n655 585
R712 B.n654 B.n179 585
R713 B.n653 B.n652 585
R714 B.n651 B.n180 585
R715 B.n650 B.n649 585
R716 B.n648 B.n181 585
R717 B.n647 B.n646 585
R718 B.n645 B.n182 585
R719 B.n644 B.n643 585
R720 B.n642 B.n183 585
R721 B.n641 B.n640 585
R722 B.n639 B.n184 585
R723 B.n638 B.n637 585
R724 B.n636 B.n185 585
R725 B.n635 B.n634 585
R726 B.n633 B.n186 585
R727 B.n632 B.n631 585
R728 B.n630 B.n187 585
R729 B.n629 B.n628 585
R730 B.n627 B.n188 585
R731 B.n626 B.n625 585
R732 B.n624 B.n189 585
R733 B.n623 B.n622 585
R734 B.n621 B.n190 585
R735 B.n620 B.n619 585
R736 B.n618 B.n191 585
R737 B.n419 B.n418 585
R738 B.n420 B.n261 585
R739 B.n422 B.n421 585
R740 B.n423 B.n260 585
R741 B.n425 B.n424 585
R742 B.n426 B.n259 585
R743 B.n428 B.n427 585
R744 B.n429 B.n258 585
R745 B.n431 B.n430 585
R746 B.n432 B.n257 585
R747 B.n434 B.n433 585
R748 B.n435 B.n256 585
R749 B.n437 B.n436 585
R750 B.n438 B.n255 585
R751 B.n440 B.n439 585
R752 B.n441 B.n254 585
R753 B.n443 B.n442 585
R754 B.n444 B.n253 585
R755 B.n446 B.n445 585
R756 B.n447 B.n252 585
R757 B.n449 B.n448 585
R758 B.n450 B.n251 585
R759 B.n452 B.n451 585
R760 B.n453 B.n250 585
R761 B.n455 B.n454 585
R762 B.n456 B.n249 585
R763 B.n458 B.n457 585
R764 B.n459 B.n248 585
R765 B.n461 B.n460 585
R766 B.n462 B.n247 585
R767 B.n464 B.n463 585
R768 B.n465 B.n246 585
R769 B.n467 B.n466 585
R770 B.n468 B.n245 585
R771 B.n470 B.n469 585
R772 B.n471 B.n244 585
R773 B.n473 B.n472 585
R774 B.n474 B.n243 585
R775 B.n476 B.n475 585
R776 B.n477 B.n242 585
R777 B.n479 B.n478 585
R778 B.n480 B.n241 585
R779 B.n482 B.n481 585
R780 B.n483 B.n240 585
R781 B.n485 B.n484 585
R782 B.n486 B.n239 585
R783 B.n488 B.n487 585
R784 B.n489 B.n238 585
R785 B.n491 B.n490 585
R786 B.n492 B.n237 585
R787 B.n494 B.n493 585
R788 B.n495 B.n236 585
R789 B.n497 B.n496 585
R790 B.n498 B.n235 585
R791 B.n500 B.n499 585
R792 B.n501 B.n234 585
R793 B.n503 B.n502 585
R794 B.n504 B.n233 585
R795 B.n506 B.n505 585
R796 B.n507 B.n232 585
R797 B.n509 B.n508 585
R798 B.n511 B.n229 585
R799 B.n513 B.n512 585
R800 B.n514 B.n228 585
R801 B.n516 B.n515 585
R802 B.n517 B.n227 585
R803 B.n519 B.n518 585
R804 B.n520 B.n226 585
R805 B.n522 B.n521 585
R806 B.n523 B.n225 585
R807 B.n525 B.n524 585
R808 B.n527 B.n526 585
R809 B.n528 B.n221 585
R810 B.n530 B.n529 585
R811 B.n531 B.n220 585
R812 B.n533 B.n532 585
R813 B.n534 B.n219 585
R814 B.n536 B.n535 585
R815 B.n537 B.n218 585
R816 B.n539 B.n538 585
R817 B.n540 B.n217 585
R818 B.n542 B.n541 585
R819 B.n543 B.n216 585
R820 B.n545 B.n544 585
R821 B.n546 B.n215 585
R822 B.n548 B.n547 585
R823 B.n549 B.n214 585
R824 B.n551 B.n550 585
R825 B.n552 B.n213 585
R826 B.n554 B.n553 585
R827 B.n555 B.n212 585
R828 B.n557 B.n556 585
R829 B.n558 B.n211 585
R830 B.n560 B.n559 585
R831 B.n561 B.n210 585
R832 B.n563 B.n562 585
R833 B.n564 B.n209 585
R834 B.n566 B.n565 585
R835 B.n567 B.n208 585
R836 B.n569 B.n568 585
R837 B.n570 B.n207 585
R838 B.n572 B.n571 585
R839 B.n573 B.n206 585
R840 B.n575 B.n574 585
R841 B.n576 B.n205 585
R842 B.n578 B.n577 585
R843 B.n579 B.n204 585
R844 B.n581 B.n580 585
R845 B.n582 B.n203 585
R846 B.n584 B.n583 585
R847 B.n585 B.n202 585
R848 B.n587 B.n586 585
R849 B.n588 B.n201 585
R850 B.n590 B.n589 585
R851 B.n591 B.n200 585
R852 B.n593 B.n592 585
R853 B.n594 B.n199 585
R854 B.n596 B.n595 585
R855 B.n597 B.n198 585
R856 B.n599 B.n598 585
R857 B.n600 B.n197 585
R858 B.n602 B.n601 585
R859 B.n603 B.n196 585
R860 B.n605 B.n604 585
R861 B.n606 B.n195 585
R862 B.n608 B.n607 585
R863 B.n609 B.n194 585
R864 B.n611 B.n610 585
R865 B.n612 B.n193 585
R866 B.n614 B.n613 585
R867 B.n615 B.n192 585
R868 B.n617 B.n616 585
R869 B.n417 B.n262 585
R870 B.n416 B.n415 585
R871 B.n414 B.n263 585
R872 B.n413 B.n412 585
R873 B.n411 B.n264 585
R874 B.n410 B.n409 585
R875 B.n408 B.n265 585
R876 B.n407 B.n406 585
R877 B.n405 B.n266 585
R878 B.n404 B.n403 585
R879 B.n402 B.n267 585
R880 B.n401 B.n400 585
R881 B.n399 B.n268 585
R882 B.n398 B.n397 585
R883 B.n396 B.n269 585
R884 B.n395 B.n394 585
R885 B.n393 B.n270 585
R886 B.n392 B.n391 585
R887 B.n390 B.n271 585
R888 B.n389 B.n388 585
R889 B.n387 B.n272 585
R890 B.n386 B.n385 585
R891 B.n384 B.n273 585
R892 B.n383 B.n382 585
R893 B.n381 B.n274 585
R894 B.n380 B.n379 585
R895 B.n378 B.n275 585
R896 B.n377 B.n376 585
R897 B.n375 B.n276 585
R898 B.n374 B.n373 585
R899 B.n372 B.n277 585
R900 B.n371 B.n370 585
R901 B.n369 B.n278 585
R902 B.n368 B.n367 585
R903 B.n366 B.n279 585
R904 B.n365 B.n364 585
R905 B.n363 B.n280 585
R906 B.n362 B.n361 585
R907 B.n360 B.n281 585
R908 B.n359 B.n358 585
R909 B.n357 B.n282 585
R910 B.n356 B.n355 585
R911 B.n354 B.n283 585
R912 B.n353 B.n352 585
R913 B.n351 B.n284 585
R914 B.n350 B.n349 585
R915 B.n348 B.n285 585
R916 B.n347 B.n346 585
R917 B.n345 B.n286 585
R918 B.n344 B.n343 585
R919 B.n342 B.n287 585
R920 B.n341 B.n340 585
R921 B.n339 B.n288 585
R922 B.n338 B.n337 585
R923 B.n336 B.n289 585
R924 B.n335 B.n334 585
R925 B.n333 B.n290 585
R926 B.n332 B.n331 585
R927 B.n330 B.n291 585
R928 B.n329 B.n328 585
R929 B.n327 B.n292 585
R930 B.n326 B.n325 585
R931 B.n324 B.n293 585
R932 B.n323 B.n322 585
R933 B.n321 B.n294 585
R934 B.n320 B.n319 585
R935 B.n318 B.n295 585
R936 B.n317 B.n316 585
R937 B.n315 B.n296 585
R938 B.n314 B.n313 585
R939 B.n312 B.n297 585
R940 B.n311 B.n310 585
R941 B.n309 B.n298 585
R942 B.n308 B.n307 585
R943 B.n306 B.n299 585
R944 B.n305 B.n304 585
R945 B.n303 B.n300 585
R946 B.n302 B.n301 585
R947 B.n2 B.n0 585
R948 B.n1173 B.n1 585
R949 B.n1172 B.n1171 585
R950 B.n1170 B.n3 585
R951 B.n1169 B.n1168 585
R952 B.n1167 B.n4 585
R953 B.n1166 B.n1165 585
R954 B.n1164 B.n5 585
R955 B.n1163 B.n1162 585
R956 B.n1161 B.n6 585
R957 B.n1160 B.n1159 585
R958 B.n1158 B.n7 585
R959 B.n1157 B.n1156 585
R960 B.n1155 B.n8 585
R961 B.n1154 B.n1153 585
R962 B.n1152 B.n9 585
R963 B.n1151 B.n1150 585
R964 B.n1149 B.n10 585
R965 B.n1148 B.n1147 585
R966 B.n1146 B.n11 585
R967 B.n1145 B.n1144 585
R968 B.n1143 B.n12 585
R969 B.n1142 B.n1141 585
R970 B.n1140 B.n13 585
R971 B.n1139 B.n1138 585
R972 B.n1137 B.n14 585
R973 B.n1136 B.n1135 585
R974 B.n1134 B.n15 585
R975 B.n1133 B.n1132 585
R976 B.n1131 B.n16 585
R977 B.n1130 B.n1129 585
R978 B.n1128 B.n17 585
R979 B.n1127 B.n1126 585
R980 B.n1125 B.n18 585
R981 B.n1124 B.n1123 585
R982 B.n1122 B.n19 585
R983 B.n1121 B.n1120 585
R984 B.n1119 B.n20 585
R985 B.n1118 B.n1117 585
R986 B.n1116 B.n21 585
R987 B.n1115 B.n1114 585
R988 B.n1113 B.n22 585
R989 B.n1112 B.n1111 585
R990 B.n1110 B.n23 585
R991 B.n1109 B.n1108 585
R992 B.n1107 B.n24 585
R993 B.n1106 B.n1105 585
R994 B.n1104 B.n25 585
R995 B.n1103 B.n1102 585
R996 B.n1101 B.n26 585
R997 B.n1100 B.n1099 585
R998 B.n1098 B.n27 585
R999 B.n1097 B.n1096 585
R1000 B.n1095 B.n28 585
R1001 B.n1094 B.n1093 585
R1002 B.n1092 B.n29 585
R1003 B.n1091 B.n1090 585
R1004 B.n1089 B.n30 585
R1005 B.n1088 B.n1087 585
R1006 B.n1086 B.n31 585
R1007 B.n1085 B.n1084 585
R1008 B.n1083 B.n32 585
R1009 B.n1082 B.n1081 585
R1010 B.n1080 B.n33 585
R1011 B.n1079 B.n1078 585
R1012 B.n1077 B.n34 585
R1013 B.n1076 B.n1075 585
R1014 B.n1074 B.n35 585
R1015 B.n1073 B.n1072 585
R1016 B.n1071 B.n36 585
R1017 B.n1070 B.n1069 585
R1018 B.n1068 B.n37 585
R1019 B.n1067 B.n1066 585
R1020 B.n1065 B.n38 585
R1021 B.n1064 B.n1063 585
R1022 B.n1062 B.n39 585
R1023 B.n1061 B.n1060 585
R1024 B.n1059 B.n40 585
R1025 B.n1058 B.n1057 585
R1026 B.n1056 B.n41 585
R1027 B.n1175 B.n1174 585
R1028 B.n418 B.n417 502.111
R1029 B.n1054 B.n41 502.111
R1030 B.n616 B.n191 502.111
R1031 B.n856 B.n855 502.111
R1032 B.n222 B.t6 330.351
R1033 B.n230 B.t3 330.351
R1034 B.n72 B.t9 330.351
R1035 B.n80 B.t0 330.351
R1036 B.n222 B.t8 188.766
R1037 B.n80 B.t1 188.766
R1038 B.n230 B.t5 188.742
R1039 B.n72 B.t10 188.742
R1040 B.n417 B.n416 163.367
R1041 B.n416 B.n263 163.367
R1042 B.n412 B.n263 163.367
R1043 B.n412 B.n411 163.367
R1044 B.n411 B.n410 163.367
R1045 B.n410 B.n265 163.367
R1046 B.n406 B.n265 163.367
R1047 B.n406 B.n405 163.367
R1048 B.n405 B.n404 163.367
R1049 B.n404 B.n267 163.367
R1050 B.n400 B.n267 163.367
R1051 B.n400 B.n399 163.367
R1052 B.n399 B.n398 163.367
R1053 B.n398 B.n269 163.367
R1054 B.n394 B.n269 163.367
R1055 B.n394 B.n393 163.367
R1056 B.n393 B.n392 163.367
R1057 B.n392 B.n271 163.367
R1058 B.n388 B.n271 163.367
R1059 B.n388 B.n387 163.367
R1060 B.n387 B.n386 163.367
R1061 B.n386 B.n273 163.367
R1062 B.n382 B.n273 163.367
R1063 B.n382 B.n381 163.367
R1064 B.n381 B.n380 163.367
R1065 B.n380 B.n275 163.367
R1066 B.n376 B.n275 163.367
R1067 B.n376 B.n375 163.367
R1068 B.n375 B.n374 163.367
R1069 B.n374 B.n277 163.367
R1070 B.n370 B.n277 163.367
R1071 B.n370 B.n369 163.367
R1072 B.n369 B.n368 163.367
R1073 B.n368 B.n279 163.367
R1074 B.n364 B.n279 163.367
R1075 B.n364 B.n363 163.367
R1076 B.n363 B.n362 163.367
R1077 B.n362 B.n281 163.367
R1078 B.n358 B.n281 163.367
R1079 B.n358 B.n357 163.367
R1080 B.n357 B.n356 163.367
R1081 B.n356 B.n283 163.367
R1082 B.n352 B.n283 163.367
R1083 B.n352 B.n351 163.367
R1084 B.n351 B.n350 163.367
R1085 B.n350 B.n285 163.367
R1086 B.n346 B.n285 163.367
R1087 B.n346 B.n345 163.367
R1088 B.n345 B.n344 163.367
R1089 B.n344 B.n287 163.367
R1090 B.n340 B.n287 163.367
R1091 B.n340 B.n339 163.367
R1092 B.n339 B.n338 163.367
R1093 B.n338 B.n289 163.367
R1094 B.n334 B.n289 163.367
R1095 B.n334 B.n333 163.367
R1096 B.n333 B.n332 163.367
R1097 B.n332 B.n291 163.367
R1098 B.n328 B.n291 163.367
R1099 B.n328 B.n327 163.367
R1100 B.n327 B.n326 163.367
R1101 B.n326 B.n293 163.367
R1102 B.n322 B.n293 163.367
R1103 B.n322 B.n321 163.367
R1104 B.n321 B.n320 163.367
R1105 B.n320 B.n295 163.367
R1106 B.n316 B.n295 163.367
R1107 B.n316 B.n315 163.367
R1108 B.n315 B.n314 163.367
R1109 B.n314 B.n297 163.367
R1110 B.n310 B.n297 163.367
R1111 B.n310 B.n309 163.367
R1112 B.n309 B.n308 163.367
R1113 B.n308 B.n299 163.367
R1114 B.n304 B.n299 163.367
R1115 B.n304 B.n303 163.367
R1116 B.n303 B.n302 163.367
R1117 B.n302 B.n2 163.367
R1118 B.n1174 B.n2 163.367
R1119 B.n1174 B.n1173 163.367
R1120 B.n1173 B.n1172 163.367
R1121 B.n1172 B.n3 163.367
R1122 B.n1168 B.n3 163.367
R1123 B.n1168 B.n1167 163.367
R1124 B.n1167 B.n1166 163.367
R1125 B.n1166 B.n5 163.367
R1126 B.n1162 B.n5 163.367
R1127 B.n1162 B.n1161 163.367
R1128 B.n1161 B.n1160 163.367
R1129 B.n1160 B.n7 163.367
R1130 B.n1156 B.n7 163.367
R1131 B.n1156 B.n1155 163.367
R1132 B.n1155 B.n1154 163.367
R1133 B.n1154 B.n9 163.367
R1134 B.n1150 B.n9 163.367
R1135 B.n1150 B.n1149 163.367
R1136 B.n1149 B.n1148 163.367
R1137 B.n1148 B.n11 163.367
R1138 B.n1144 B.n11 163.367
R1139 B.n1144 B.n1143 163.367
R1140 B.n1143 B.n1142 163.367
R1141 B.n1142 B.n13 163.367
R1142 B.n1138 B.n13 163.367
R1143 B.n1138 B.n1137 163.367
R1144 B.n1137 B.n1136 163.367
R1145 B.n1136 B.n15 163.367
R1146 B.n1132 B.n15 163.367
R1147 B.n1132 B.n1131 163.367
R1148 B.n1131 B.n1130 163.367
R1149 B.n1130 B.n17 163.367
R1150 B.n1126 B.n17 163.367
R1151 B.n1126 B.n1125 163.367
R1152 B.n1125 B.n1124 163.367
R1153 B.n1124 B.n19 163.367
R1154 B.n1120 B.n19 163.367
R1155 B.n1120 B.n1119 163.367
R1156 B.n1119 B.n1118 163.367
R1157 B.n1118 B.n21 163.367
R1158 B.n1114 B.n21 163.367
R1159 B.n1114 B.n1113 163.367
R1160 B.n1113 B.n1112 163.367
R1161 B.n1112 B.n23 163.367
R1162 B.n1108 B.n23 163.367
R1163 B.n1108 B.n1107 163.367
R1164 B.n1107 B.n1106 163.367
R1165 B.n1106 B.n25 163.367
R1166 B.n1102 B.n25 163.367
R1167 B.n1102 B.n1101 163.367
R1168 B.n1101 B.n1100 163.367
R1169 B.n1100 B.n27 163.367
R1170 B.n1096 B.n27 163.367
R1171 B.n1096 B.n1095 163.367
R1172 B.n1095 B.n1094 163.367
R1173 B.n1094 B.n29 163.367
R1174 B.n1090 B.n29 163.367
R1175 B.n1090 B.n1089 163.367
R1176 B.n1089 B.n1088 163.367
R1177 B.n1088 B.n31 163.367
R1178 B.n1084 B.n31 163.367
R1179 B.n1084 B.n1083 163.367
R1180 B.n1083 B.n1082 163.367
R1181 B.n1082 B.n33 163.367
R1182 B.n1078 B.n33 163.367
R1183 B.n1078 B.n1077 163.367
R1184 B.n1077 B.n1076 163.367
R1185 B.n1076 B.n35 163.367
R1186 B.n1072 B.n35 163.367
R1187 B.n1072 B.n1071 163.367
R1188 B.n1071 B.n1070 163.367
R1189 B.n1070 B.n37 163.367
R1190 B.n1066 B.n37 163.367
R1191 B.n1066 B.n1065 163.367
R1192 B.n1065 B.n1064 163.367
R1193 B.n1064 B.n39 163.367
R1194 B.n1060 B.n39 163.367
R1195 B.n1060 B.n1059 163.367
R1196 B.n1059 B.n1058 163.367
R1197 B.n1058 B.n41 163.367
R1198 B.n418 B.n261 163.367
R1199 B.n422 B.n261 163.367
R1200 B.n423 B.n422 163.367
R1201 B.n424 B.n423 163.367
R1202 B.n424 B.n259 163.367
R1203 B.n428 B.n259 163.367
R1204 B.n429 B.n428 163.367
R1205 B.n430 B.n429 163.367
R1206 B.n430 B.n257 163.367
R1207 B.n434 B.n257 163.367
R1208 B.n435 B.n434 163.367
R1209 B.n436 B.n435 163.367
R1210 B.n436 B.n255 163.367
R1211 B.n440 B.n255 163.367
R1212 B.n441 B.n440 163.367
R1213 B.n442 B.n441 163.367
R1214 B.n442 B.n253 163.367
R1215 B.n446 B.n253 163.367
R1216 B.n447 B.n446 163.367
R1217 B.n448 B.n447 163.367
R1218 B.n448 B.n251 163.367
R1219 B.n452 B.n251 163.367
R1220 B.n453 B.n452 163.367
R1221 B.n454 B.n453 163.367
R1222 B.n454 B.n249 163.367
R1223 B.n458 B.n249 163.367
R1224 B.n459 B.n458 163.367
R1225 B.n460 B.n459 163.367
R1226 B.n460 B.n247 163.367
R1227 B.n464 B.n247 163.367
R1228 B.n465 B.n464 163.367
R1229 B.n466 B.n465 163.367
R1230 B.n466 B.n245 163.367
R1231 B.n470 B.n245 163.367
R1232 B.n471 B.n470 163.367
R1233 B.n472 B.n471 163.367
R1234 B.n472 B.n243 163.367
R1235 B.n476 B.n243 163.367
R1236 B.n477 B.n476 163.367
R1237 B.n478 B.n477 163.367
R1238 B.n478 B.n241 163.367
R1239 B.n482 B.n241 163.367
R1240 B.n483 B.n482 163.367
R1241 B.n484 B.n483 163.367
R1242 B.n484 B.n239 163.367
R1243 B.n488 B.n239 163.367
R1244 B.n489 B.n488 163.367
R1245 B.n490 B.n489 163.367
R1246 B.n490 B.n237 163.367
R1247 B.n494 B.n237 163.367
R1248 B.n495 B.n494 163.367
R1249 B.n496 B.n495 163.367
R1250 B.n496 B.n235 163.367
R1251 B.n500 B.n235 163.367
R1252 B.n501 B.n500 163.367
R1253 B.n502 B.n501 163.367
R1254 B.n502 B.n233 163.367
R1255 B.n506 B.n233 163.367
R1256 B.n507 B.n506 163.367
R1257 B.n508 B.n507 163.367
R1258 B.n508 B.n229 163.367
R1259 B.n513 B.n229 163.367
R1260 B.n514 B.n513 163.367
R1261 B.n515 B.n514 163.367
R1262 B.n515 B.n227 163.367
R1263 B.n519 B.n227 163.367
R1264 B.n520 B.n519 163.367
R1265 B.n521 B.n520 163.367
R1266 B.n521 B.n225 163.367
R1267 B.n525 B.n225 163.367
R1268 B.n526 B.n525 163.367
R1269 B.n526 B.n221 163.367
R1270 B.n530 B.n221 163.367
R1271 B.n531 B.n530 163.367
R1272 B.n532 B.n531 163.367
R1273 B.n532 B.n219 163.367
R1274 B.n536 B.n219 163.367
R1275 B.n537 B.n536 163.367
R1276 B.n538 B.n537 163.367
R1277 B.n538 B.n217 163.367
R1278 B.n542 B.n217 163.367
R1279 B.n543 B.n542 163.367
R1280 B.n544 B.n543 163.367
R1281 B.n544 B.n215 163.367
R1282 B.n548 B.n215 163.367
R1283 B.n549 B.n548 163.367
R1284 B.n550 B.n549 163.367
R1285 B.n550 B.n213 163.367
R1286 B.n554 B.n213 163.367
R1287 B.n555 B.n554 163.367
R1288 B.n556 B.n555 163.367
R1289 B.n556 B.n211 163.367
R1290 B.n560 B.n211 163.367
R1291 B.n561 B.n560 163.367
R1292 B.n562 B.n561 163.367
R1293 B.n562 B.n209 163.367
R1294 B.n566 B.n209 163.367
R1295 B.n567 B.n566 163.367
R1296 B.n568 B.n567 163.367
R1297 B.n568 B.n207 163.367
R1298 B.n572 B.n207 163.367
R1299 B.n573 B.n572 163.367
R1300 B.n574 B.n573 163.367
R1301 B.n574 B.n205 163.367
R1302 B.n578 B.n205 163.367
R1303 B.n579 B.n578 163.367
R1304 B.n580 B.n579 163.367
R1305 B.n580 B.n203 163.367
R1306 B.n584 B.n203 163.367
R1307 B.n585 B.n584 163.367
R1308 B.n586 B.n585 163.367
R1309 B.n586 B.n201 163.367
R1310 B.n590 B.n201 163.367
R1311 B.n591 B.n590 163.367
R1312 B.n592 B.n591 163.367
R1313 B.n592 B.n199 163.367
R1314 B.n596 B.n199 163.367
R1315 B.n597 B.n596 163.367
R1316 B.n598 B.n597 163.367
R1317 B.n598 B.n197 163.367
R1318 B.n602 B.n197 163.367
R1319 B.n603 B.n602 163.367
R1320 B.n604 B.n603 163.367
R1321 B.n604 B.n195 163.367
R1322 B.n608 B.n195 163.367
R1323 B.n609 B.n608 163.367
R1324 B.n610 B.n609 163.367
R1325 B.n610 B.n193 163.367
R1326 B.n614 B.n193 163.367
R1327 B.n615 B.n614 163.367
R1328 B.n616 B.n615 163.367
R1329 B.n620 B.n191 163.367
R1330 B.n621 B.n620 163.367
R1331 B.n622 B.n621 163.367
R1332 B.n622 B.n189 163.367
R1333 B.n626 B.n189 163.367
R1334 B.n627 B.n626 163.367
R1335 B.n628 B.n627 163.367
R1336 B.n628 B.n187 163.367
R1337 B.n632 B.n187 163.367
R1338 B.n633 B.n632 163.367
R1339 B.n634 B.n633 163.367
R1340 B.n634 B.n185 163.367
R1341 B.n638 B.n185 163.367
R1342 B.n639 B.n638 163.367
R1343 B.n640 B.n639 163.367
R1344 B.n640 B.n183 163.367
R1345 B.n644 B.n183 163.367
R1346 B.n645 B.n644 163.367
R1347 B.n646 B.n645 163.367
R1348 B.n646 B.n181 163.367
R1349 B.n650 B.n181 163.367
R1350 B.n651 B.n650 163.367
R1351 B.n652 B.n651 163.367
R1352 B.n652 B.n179 163.367
R1353 B.n656 B.n179 163.367
R1354 B.n657 B.n656 163.367
R1355 B.n658 B.n657 163.367
R1356 B.n658 B.n177 163.367
R1357 B.n662 B.n177 163.367
R1358 B.n663 B.n662 163.367
R1359 B.n664 B.n663 163.367
R1360 B.n664 B.n175 163.367
R1361 B.n668 B.n175 163.367
R1362 B.n669 B.n668 163.367
R1363 B.n670 B.n669 163.367
R1364 B.n670 B.n173 163.367
R1365 B.n674 B.n173 163.367
R1366 B.n675 B.n674 163.367
R1367 B.n676 B.n675 163.367
R1368 B.n676 B.n171 163.367
R1369 B.n680 B.n171 163.367
R1370 B.n681 B.n680 163.367
R1371 B.n682 B.n681 163.367
R1372 B.n682 B.n169 163.367
R1373 B.n686 B.n169 163.367
R1374 B.n687 B.n686 163.367
R1375 B.n688 B.n687 163.367
R1376 B.n688 B.n167 163.367
R1377 B.n692 B.n167 163.367
R1378 B.n693 B.n692 163.367
R1379 B.n694 B.n693 163.367
R1380 B.n694 B.n165 163.367
R1381 B.n698 B.n165 163.367
R1382 B.n699 B.n698 163.367
R1383 B.n700 B.n699 163.367
R1384 B.n700 B.n163 163.367
R1385 B.n704 B.n163 163.367
R1386 B.n705 B.n704 163.367
R1387 B.n706 B.n705 163.367
R1388 B.n706 B.n161 163.367
R1389 B.n710 B.n161 163.367
R1390 B.n711 B.n710 163.367
R1391 B.n712 B.n711 163.367
R1392 B.n712 B.n159 163.367
R1393 B.n716 B.n159 163.367
R1394 B.n717 B.n716 163.367
R1395 B.n718 B.n717 163.367
R1396 B.n718 B.n157 163.367
R1397 B.n722 B.n157 163.367
R1398 B.n723 B.n722 163.367
R1399 B.n724 B.n723 163.367
R1400 B.n724 B.n155 163.367
R1401 B.n728 B.n155 163.367
R1402 B.n729 B.n728 163.367
R1403 B.n730 B.n729 163.367
R1404 B.n730 B.n153 163.367
R1405 B.n734 B.n153 163.367
R1406 B.n735 B.n734 163.367
R1407 B.n736 B.n735 163.367
R1408 B.n736 B.n151 163.367
R1409 B.n740 B.n151 163.367
R1410 B.n741 B.n740 163.367
R1411 B.n742 B.n741 163.367
R1412 B.n742 B.n149 163.367
R1413 B.n746 B.n149 163.367
R1414 B.n747 B.n746 163.367
R1415 B.n748 B.n747 163.367
R1416 B.n748 B.n147 163.367
R1417 B.n752 B.n147 163.367
R1418 B.n753 B.n752 163.367
R1419 B.n754 B.n753 163.367
R1420 B.n754 B.n145 163.367
R1421 B.n758 B.n145 163.367
R1422 B.n759 B.n758 163.367
R1423 B.n760 B.n759 163.367
R1424 B.n760 B.n143 163.367
R1425 B.n764 B.n143 163.367
R1426 B.n765 B.n764 163.367
R1427 B.n766 B.n765 163.367
R1428 B.n766 B.n141 163.367
R1429 B.n770 B.n141 163.367
R1430 B.n771 B.n770 163.367
R1431 B.n772 B.n771 163.367
R1432 B.n772 B.n139 163.367
R1433 B.n776 B.n139 163.367
R1434 B.n777 B.n776 163.367
R1435 B.n778 B.n777 163.367
R1436 B.n778 B.n137 163.367
R1437 B.n782 B.n137 163.367
R1438 B.n783 B.n782 163.367
R1439 B.n784 B.n783 163.367
R1440 B.n784 B.n135 163.367
R1441 B.n788 B.n135 163.367
R1442 B.n789 B.n788 163.367
R1443 B.n790 B.n789 163.367
R1444 B.n790 B.n133 163.367
R1445 B.n794 B.n133 163.367
R1446 B.n795 B.n794 163.367
R1447 B.n796 B.n795 163.367
R1448 B.n796 B.n131 163.367
R1449 B.n800 B.n131 163.367
R1450 B.n801 B.n800 163.367
R1451 B.n802 B.n801 163.367
R1452 B.n802 B.n129 163.367
R1453 B.n806 B.n129 163.367
R1454 B.n807 B.n806 163.367
R1455 B.n808 B.n807 163.367
R1456 B.n808 B.n127 163.367
R1457 B.n812 B.n127 163.367
R1458 B.n813 B.n812 163.367
R1459 B.n814 B.n813 163.367
R1460 B.n814 B.n125 163.367
R1461 B.n818 B.n125 163.367
R1462 B.n819 B.n818 163.367
R1463 B.n820 B.n819 163.367
R1464 B.n820 B.n123 163.367
R1465 B.n824 B.n123 163.367
R1466 B.n825 B.n824 163.367
R1467 B.n826 B.n825 163.367
R1468 B.n826 B.n121 163.367
R1469 B.n830 B.n121 163.367
R1470 B.n831 B.n830 163.367
R1471 B.n832 B.n831 163.367
R1472 B.n832 B.n119 163.367
R1473 B.n836 B.n119 163.367
R1474 B.n837 B.n836 163.367
R1475 B.n838 B.n837 163.367
R1476 B.n838 B.n117 163.367
R1477 B.n842 B.n117 163.367
R1478 B.n843 B.n842 163.367
R1479 B.n844 B.n843 163.367
R1480 B.n844 B.n115 163.367
R1481 B.n848 B.n115 163.367
R1482 B.n849 B.n848 163.367
R1483 B.n850 B.n849 163.367
R1484 B.n850 B.n113 163.367
R1485 B.n854 B.n113 163.367
R1486 B.n855 B.n854 163.367
R1487 B.n1054 B.n1053 163.367
R1488 B.n1053 B.n1052 163.367
R1489 B.n1052 B.n43 163.367
R1490 B.n1048 B.n43 163.367
R1491 B.n1048 B.n1047 163.367
R1492 B.n1047 B.n1046 163.367
R1493 B.n1046 B.n45 163.367
R1494 B.n1042 B.n45 163.367
R1495 B.n1042 B.n1041 163.367
R1496 B.n1041 B.n1040 163.367
R1497 B.n1040 B.n47 163.367
R1498 B.n1036 B.n47 163.367
R1499 B.n1036 B.n1035 163.367
R1500 B.n1035 B.n1034 163.367
R1501 B.n1034 B.n49 163.367
R1502 B.n1030 B.n49 163.367
R1503 B.n1030 B.n1029 163.367
R1504 B.n1029 B.n1028 163.367
R1505 B.n1028 B.n51 163.367
R1506 B.n1024 B.n51 163.367
R1507 B.n1024 B.n1023 163.367
R1508 B.n1023 B.n1022 163.367
R1509 B.n1022 B.n53 163.367
R1510 B.n1018 B.n53 163.367
R1511 B.n1018 B.n1017 163.367
R1512 B.n1017 B.n1016 163.367
R1513 B.n1016 B.n55 163.367
R1514 B.n1012 B.n55 163.367
R1515 B.n1012 B.n1011 163.367
R1516 B.n1011 B.n1010 163.367
R1517 B.n1010 B.n57 163.367
R1518 B.n1006 B.n57 163.367
R1519 B.n1006 B.n1005 163.367
R1520 B.n1005 B.n1004 163.367
R1521 B.n1004 B.n59 163.367
R1522 B.n1000 B.n59 163.367
R1523 B.n1000 B.n999 163.367
R1524 B.n999 B.n998 163.367
R1525 B.n998 B.n61 163.367
R1526 B.n994 B.n61 163.367
R1527 B.n994 B.n993 163.367
R1528 B.n993 B.n992 163.367
R1529 B.n992 B.n63 163.367
R1530 B.n988 B.n63 163.367
R1531 B.n988 B.n987 163.367
R1532 B.n987 B.n986 163.367
R1533 B.n986 B.n65 163.367
R1534 B.n982 B.n65 163.367
R1535 B.n982 B.n981 163.367
R1536 B.n981 B.n980 163.367
R1537 B.n980 B.n67 163.367
R1538 B.n976 B.n67 163.367
R1539 B.n976 B.n975 163.367
R1540 B.n975 B.n974 163.367
R1541 B.n974 B.n69 163.367
R1542 B.n970 B.n69 163.367
R1543 B.n970 B.n969 163.367
R1544 B.n969 B.n968 163.367
R1545 B.n968 B.n71 163.367
R1546 B.n964 B.n71 163.367
R1547 B.n964 B.n963 163.367
R1548 B.n963 B.n75 163.367
R1549 B.n959 B.n75 163.367
R1550 B.n959 B.n958 163.367
R1551 B.n958 B.n957 163.367
R1552 B.n957 B.n77 163.367
R1553 B.n953 B.n77 163.367
R1554 B.n953 B.n952 163.367
R1555 B.n952 B.n951 163.367
R1556 B.n951 B.n79 163.367
R1557 B.n946 B.n79 163.367
R1558 B.n946 B.n945 163.367
R1559 B.n945 B.n944 163.367
R1560 B.n944 B.n83 163.367
R1561 B.n940 B.n83 163.367
R1562 B.n940 B.n939 163.367
R1563 B.n939 B.n938 163.367
R1564 B.n938 B.n85 163.367
R1565 B.n934 B.n85 163.367
R1566 B.n934 B.n933 163.367
R1567 B.n933 B.n932 163.367
R1568 B.n932 B.n87 163.367
R1569 B.n928 B.n87 163.367
R1570 B.n928 B.n927 163.367
R1571 B.n927 B.n926 163.367
R1572 B.n926 B.n89 163.367
R1573 B.n922 B.n89 163.367
R1574 B.n922 B.n921 163.367
R1575 B.n921 B.n920 163.367
R1576 B.n920 B.n91 163.367
R1577 B.n916 B.n91 163.367
R1578 B.n916 B.n915 163.367
R1579 B.n915 B.n914 163.367
R1580 B.n914 B.n93 163.367
R1581 B.n910 B.n93 163.367
R1582 B.n910 B.n909 163.367
R1583 B.n909 B.n908 163.367
R1584 B.n908 B.n95 163.367
R1585 B.n904 B.n95 163.367
R1586 B.n904 B.n903 163.367
R1587 B.n903 B.n902 163.367
R1588 B.n902 B.n97 163.367
R1589 B.n898 B.n97 163.367
R1590 B.n898 B.n897 163.367
R1591 B.n897 B.n896 163.367
R1592 B.n896 B.n99 163.367
R1593 B.n892 B.n99 163.367
R1594 B.n892 B.n891 163.367
R1595 B.n891 B.n890 163.367
R1596 B.n890 B.n101 163.367
R1597 B.n886 B.n101 163.367
R1598 B.n886 B.n885 163.367
R1599 B.n885 B.n884 163.367
R1600 B.n884 B.n103 163.367
R1601 B.n880 B.n103 163.367
R1602 B.n880 B.n879 163.367
R1603 B.n879 B.n878 163.367
R1604 B.n878 B.n105 163.367
R1605 B.n874 B.n105 163.367
R1606 B.n874 B.n873 163.367
R1607 B.n873 B.n872 163.367
R1608 B.n872 B.n107 163.367
R1609 B.n868 B.n107 163.367
R1610 B.n868 B.n867 163.367
R1611 B.n867 B.n866 163.367
R1612 B.n866 B.n109 163.367
R1613 B.n862 B.n109 163.367
R1614 B.n862 B.n861 163.367
R1615 B.n861 B.n860 163.367
R1616 B.n860 B.n111 163.367
R1617 B.n856 B.n111 163.367
R1618 B.n223 B.t7 110.609
R1619 B.n81 B.t2 110.609
R1620 B.n231 B.t4 110.585
R1621 B.n73 B.t11 110.585
R1622 B.n223 B.n222 78.1581
R1623 B.n231 B.n230 78.1581
R1624 B.n73 B.n72 78.1581
R1625 B.n81 B.n80 78.1581
R1626 B.n224 B.n223 59.5399
R1627 B.n510 B.n231 59.5399
R1628 B.n74 B.n73 59.5399
R1629 B.n948 B.n81 59.5399
R1630 B.n1056 B.n1055 32.6249
R1631 B.n857 B.n112 32.6249
R1632 B.n618 B.n617 32.6249
R1633 B.n419 B.n262 32.6249
R1634 B B.n1175 18.0485
R1635 B.n1055 B.n42 10.6151
R1636 B.n1051 B.n42 10.6151
R1637 B.n1051 B.n1050 10.6151
R1638 B.n1050 B.n1049 10.6151
R1639 B.n1049 B.n44 10.6151
R1640 B.n1045 B.n44 10.6151
R1641 B.n1045 B.n1044 10.6151
R1642 B.n1044 B.n1043 10.6151
R1643 B.n1043 B.n46 10.6151
R1644 B.n1039 B.n46 10.6151
R1645 B.n1039 B.n1038 10.6151
R1646 B.n1038 B.n1037 10.6151
R1647 B.n1037 B.n48 10.6151
R1648 B.n1033 B.n48 10.6151
R1649 B.n1033 B.n1032 10.6151
R1650 B.n1032 B.n1031 10.6151
R1651 B.n1031 B.n50 10.6151
R1652 B.n1027 B.n50 10.6151
R1653 B.n1027 B.n1026 10.6151
R1654 B.n1026 B.n1025 10.6151
R1655 B.n1025 B.n52 10.6151
R1656 B.n1021 B.n52 10.6151
R1657 B.n1021 B.n1020 10.6151
R1658 B.n1020 B.n1019 10.6151
R1659 B.n1019 B.n54 10.6151
R1660 B.n1015 B.n54 10.6151
R1661 B.n1015 B.n1014 10.6151
R1662 B.n1014 B.n1013 10.6151
R1663 B.n1013 B.n56 10.6151
R1664 B.n1009 B.n56 10.6151
R1665 B.n1009 B.n1008 10.6151
R1666 B.n1008 B.n1007 10.6151
R1667 B.n1007 B.n58 10.6151
R1668 B.n1003 B.n58 10.6151
R1669 B.n1003 B.n1002 10.6151
R1670 B.n1002 B.n1001 10.6151
R1671 B.n1001 B.n60 10.6151
R1672 B.n997 B.n60 10.6151
R1673 B.n997 B.n996 10.6151
R1674 B.n996 B.n995 10.6151
R1675 B.n995 B.n62 10.6151
R1676 B.n991 B.n62 10.6151
R1677 B.n991 B.n990 10.6151
R1678 B.n990 B.n989 10.6151
R1679 B.n989 B.n64 10.6151
R1680 B.n985 B.n64 10.6151
R1681 B.n985 B.n984 10.6151
R1682 B.n984 B.n983 10.6151
R1683 B.n983 B.n66 10.6151
R1684 B.n979 B.n66 10.6151
R1685 B.n979 B.n978 10.6151
R1686 B.n978 B.n977 10.6151
R1687 B.n977 B.n68 10.6151
R1688 B.n973 B.n68 10.6151
R1689 B.n973 B.n972 10.6151
R1690 B.n972 B.n971 10.6151
R1691 B.n971 B.n70 10.6151
R1692 B.n967 B.n70 10.6151
R1693 B.n967 B.n966 10.6151
R1694 B.n966 B.n965 10.6151
R1695 B.n962 B.n961 10.6151
R1696 B.n961 B.n960 10.6151
R1697 B.n960 B.n76 10.6151
R1698 B.n956 B.n76 10.6151
R1699 B.n956 B.n955 10.6151
R1700 B.n955 B.n954 10.6151
R1701 B.n954 B.n78 10.6151
R1702 B.n950 B.n78 10.6151
R1703 B.n950 B.n949 10.6151
R1704 B.n947 B.n82 10.6151
R1705 B.n943 B.n82 10.6151
R1706 B.n943 B.n942 10.6151
R1707 B.n942 B.n941 10.6151
R1708 B.n941 B.n84 10.6151
R1709 B.n937 B.n84 10.6151
R1710 B.n937 B.n936 10.6151
R1711 B.n936 B.n935 10.6151
R1712 B.n935 B.n86 10.6151
R1713 B.n931 B.n86 10.6151
R1714 B.n931 B.n930 10.6151
R1715 B.n930 B.n929 10.6151
R1716 B.n929 B.n88 10.6151
R1717 B.n925 B.n88 10.6151
R1718 B.n925 B.n924 10.6151
R1719 B.n924 B.n923 10.6151
R1720 B.n923 B.n90 10.6151
R1721 B.n919 B.n90 10.6151
R1722 B.n919 B.n918 10.6151
R1723 B.n918 B.n917 10.6151
R1724 B.n917 B.n92 10.6151
R1725 B.n913 B.n92 10.6151
R1726 B.n913 B.n912 10.6151
R1727 B.n912 B.n911 10.6151
R1728 B.n911 B.n94 10.6151
R1729 B.n907 B.n94 10.6151
R1730 B.n907 B.n906 10.6151
R1731 B.n906 B.n905 10.6151
R1732 B.n905 B.n96 10.6151
R1733 B.n901 B.n96 10.6151
R1734 B.n901 B.n900 10.6151
R1735 B.n900 B.n899 10.6151
R1736 B.n899 B.n98 10.6151
R1737 B.n895 B.n98 10.6151
R1738 B.n895 B.n894 10.6151
R1739 B.n894 B.n893 10.6151
R1740 B.n893 B.n100 10.6151
R1741 B.n889 B.n100 10.6151
R1742 B.n889 B.n888 10.6151
R1743 B.n888 B.n887 10.6151
R1744 B.n887 B.n102 10.6151
R1745 B.n883 B.n102 10.6151
R1746 B.n883 B.n882 10.6151
R1747 B.n882 B.n881 10.6151
R1748 B.n881 B.n104 10.6151
R1749 B.n877 B.n104 10.6151
R1750 B.n877 B.n876 10.6151
R1751 B.n876 B.n875 10.6151
R1752 B.n875 B.n106 10.6151
R1753 B.n871 B.n106 10.6151
R1754 B.n871 B.n870 10.6151
R1755 B.n870 B.n869 10.6151
R1756 B.n869 B.n108 10.6151
R1757 B.n865 B.n108 10.6151
R1758 B.n865 B.n864 10.6151
R1759 B.n864 B.n863 10.6151
R1760 B.n863 B.n110 10.6151
R1761 B.n859 B.n110 10.6151
R1762 B.n859 B.n858 10.6151
R1763 B.n858 B.n857 10.6151
R1764 B.n619 B.n618 10.6151
R1765 B.n619 B.n190 10.6151
R1766 B.n623 B.n190 10.6151
R1767 B.n624 B.n623 10.6151
R1768 B.n625 B.n624 10.6151
R1769 B.n625 B.n188 10.6151
R1770 B.n629 B.n188 10.6151
R1771 B.n630 B.n629 10.6151
R1772 B.n631 B.n630 10.6151
R1773 B.n631 B.n186 10.6151
R1774 B.n635 B.n186 10.6151
R1775 B.n636 B.n635 10.6151
R1776 B.n637 B.n636 10.6151
R1777 B.n637 B.n184 10.6151
R1778 B.n641 B.n184 10.6151
R1779 B.n642 B.n641 10.6151
R1780 B.n643 B.n642 10.6151
R1781 B.n643 B.n182 10.6151
R1782 B.n647 B.n182 10.6151
R1783 B.n648 B.n647 10.6151
R1784 B.n649 B.n648 10.6151
R1785 B.n649 B.n180 10.6151
R1786 B.n653 B.n180 10.6151
R1787 B.n654 B.n653 10.6151
R1788 B.n655 B.n654 10.6151
R1789 B.n655 B.n178 10.6151
R1790 B.n659 B.n178 10.6151
R1791 B.n660 B.n659 10.6151
R1792 B.n661 B.n660 10.6151
R1793 B.n661 B.n176 10.6151
R1794 B.n665 B.n176 10.6151
R1795 B.n666 B.n665 10.6151
R1796 B.n667 B.n666 10.6151
R1797 B.n667 B.n174 10.6151
R1798 B.n671 B.n174 10.6151
R1799 B.n672 B.n671 10.6151
R1800 B.n673 B.n672 10.6151
R1801 B.n673 B.n172 10.6151
R1802 B.n677 B.n172 10.6151
R1803 B.n678 B.n677 10.6151
R1804 B.n679 B.n678 10.6151
R1805 B.n679 B.n170 10.6151
R1806 B.n683 B.n170 10.6151
R1807 B.n684 B.n683 10.6151
R1808 B.n685 B.n684 10.6151
R1809 B.n685 B.n168 10.6151
R1810 B.n689 B.n168 10.6151
R1811 B.n690 B.n689 10.6151
R1812 B.n691 B.n690 10.6151
R1813 B.n691 B.n166 10.6151
R1814 B.n695 B.n166 10.6151
R1815 B.n696 B.n695 10.6151
R1816 B.n697 B.n696 10.6151
R1817 B.n697 B.n164 10.6151
R1818 B.n701 B.n164 10.6151
R1819 B.n702 B.n701 10.6151
R1820 B.n703 B.n702 10.6151
R1821 B.n703 B.n162 10.6151
R1822 B.n707 B.n162 10.6151
R1823 B.n708 B.n707 10.6151
R1824 B.n709 B.n708 10.6151
R1825 B.n709 B.n160 10.6151
R1826 B.n713 B.n160 10.6151
R1827 B.n714 B.n713 10.6151
R1828 B.n715 B.n714 10.6151
R1829 B.n715 B.n158 10.6151
R1830 B.n719 B.n158 10.6151
R1831 B.n720 B.n719 10.6151
R1832 B.n721 B.n720 10.6151
R1833 B.n721 B.n156 10.6151
R1834 B.n725 B.n156 10.6151
R1835 B.n726 B.n725 10.6151
R1836 B.n727 B.n726 10.6151
R1837 B.n727 B.n154 10.6151
R1838 B.n731 B.n154 10.6151
R1839 B.n732 B.n731 10.6151
R1840 B.n733 B.n732 10.6151
R1841 B.n733 B.n152 10.6151
R1842 B.n737 B.n152 10.6151
R1843 B.n738 B.n737 10.6151
R1844 B.n739 B.n738 10.6151
R1845 B.n739 B.n150 10.6151
R1846 B.n743 B.n150 10.6151
R1847 B.n744 B.n743 10.6151
R1848 B.n745 B.n744 10.6151
R1849 B.n745 B.n148 10.6151
R1850 B.n749 B.n148 10.6151
R1851 B.n750 B.n749 10.6151
R1852 B.n751 B.n750 10.6151
R1853 B.n751 B.n146 10.6151
R1854 B.n755 B.n146 10.6151
R1855 B.n756 B.n755 10.6151
R1856 B.n757 B.n756 10.6151
R1857 B.n757 B.n144 10.6151
R1858 B.n761 B.n144 10.6151
R1859 B.n762 B.n761 10.6151
R1860 B.n763 B.n762 10.6151
R1861 B.n763 B.n142 10.6151
R1862 B.n767 B.n142 10.6151
R1863 B.n768 B.n767 10.6151
R1864 B.n769 B.n768 10.6151
R1865 B.n769 B.n140 10.6151
R1866 B.n773 B.n140 10.6151
R1867 B.n774 B.n773 10.6151
R1868 B.n775 B.n774 10.6151
R1869 B.n775 B.n138 10.6151
R1870 B.n779 B.n138 10.6151
R1871 B.n780 B.n779 10.6151
R1872 B.n781 B.n780 10.6151
R1873 B.n781 B.n136 10.6151
R1874 B.n785 B.n136 10.6151
R1875 B.n786 B.n785 10.6151
R1876 B.n787 B.n786 10.6151
R1877 B.n787 B.n134 10.6151
R1878 B.n791 B.n134 10.6151
R1879 B.n792 B.n791 10.6151
R1880 B.n793 B.n792 10.6151
R1881 B.n793 B.n132 10.6151
R1882 B.n797 B.n132 10.6151
R1883 B.n798 B.n797 10.6151
R1884 B.n799 B.n798 10.6151
R1885 B.n799 B.n130 10.6151
R1886 B.n803 B.n130 10.6151
R1887 B.n804 B.n803 10.6151
R1888 B.n805 B.n804 10.6151
R1889 B.n805 B.n128 10.6151
R1890 B.n809 B.n128 10.6151
R1891 B.n810 B.n809 10.6151
R1892 B.n811 B.n810 10.6151
R1893 B.n811 B.n126 10.6151
R1894 B.n815 B.n126 10.6151
R1895 B.n816 B.n815 10.6151
R1896 B.n817 B.n816 10.6151
R1897 B.n817 B.n124 10.6151
R1898 B.n821 B.n124 10.6151
R1899 B.n822 B.n821 10.6151
R1900 B.n823 B.n822 10.6151
R1901 B.n823 B.n122 10.6151
R1902 B.n827 B.n122 10.6151
R1903 B.n828 B.n827 10.6151
R1904 B.n829 B.n828 10.6151
R1905 B.n829 B.n120 10.6151
R1906 B.n833 B.n120 10.6151
R1907 B.n834 B.n833 10.6151
R1908 B.n835 B.n834 10.6151
R1909 B.n835 B.n118 10.6151
R1910 B.n839 B.n118 10.6151
R1911 B.n840 B.n839 10.6151
R1912 B.n841 B.n840 10.6151
R1913 B.n841 B.n116 10.6151
R1914 B.n845 B.n116 10.6151
R1915 B.n846 B.n845 10.6151
R1916 B.n847 B.n846 10.6151
R1917 B.n847 B.n114 10.6151
R1918 B.n851 B.n114 10.6151
R1919 B.n852 B.n851 10.6151
R1920 B.n853 B.n852 10.6151
R1921 B.n853 B.n112 10.6151
R1922 B.n420 B.n419 10.6151
R1923 B.n421 B.n420 10.6151
R1924 B.n421 B.n260 10.6151
R1925 B.n425 B.n260 10.6151
R1926 B.n426 B.n425 10.6151
R1927 B.n427 B.n426 10.6151
R1928 B.n427 B.n258 10.6151
R1929 B.n431 B.n258 10.6151
R1930 B.n432 B.n431 10.6151
R1931 B.n433 B.n432 10.6151
R1932 B.n433 B.n256 10.6151
R1933 B.n437 B.n256 10.6151
R1934 B.n438 B.n437 10.6151
R1935 B.n439 B.n438 10.6151
R1936 B.n439 B.n254 10.6151
R1937 B.n443 B.n254 10.6151
R1938 B.n444 B.n443 10.6151
R1939 B.n445 B.n444 10.6151
R1940 B.n445 B.n252 10.6151
R1941 B.n449 B.n252 10.6151
R1942 B.n450 B.n449 10.6151
R1943 B.n451 B.n450 10.6151
R1944 B.n451 B.n250 10.6151
R1945 B.n455 B.n250 10.6151
R1946 B.n456 B.n455 10.6151
R1947 B.n457 B.n456 10.6151
R1948 B.n457 B.n248 10.6151
R1949 B.n461 B.n248 10.6151
R1950 B.n462 B.n461 10.6151
R1951 B.n463 B.n462 10.6151
R1952 B.n463 B.n246 10.6151
R1953 B.n467 B.n246 10.6151
R1954 B.n468 B.n467 10.6151
R1955 B.n469 B.n468 10.6151
R1956 B.n469 B.n244 10.6151
R1957 B.n473 B.n244 10.6151
R1958 B.n474 B.n473 10.6151
R1959 B.n475 B.n474 10.6151
R1960 B.n475 B.n242 10.6151
R1961 B.n479 B.n242 10.6151
R1962 B.n480 B.n479 10.6151
R1963 B.n481 B.n480 10.6151
R1964 B.n481 B.n240 10.6151
R1965 B.n485 B.n240 10.6151
R1966 B.n486 B.n485 10.6151
R1967 B.n487 B.n486 10.6151
R1968 B.n487 B.n238 10.6151
R1969 B.n491 B.n238 10.6151
R1970 B.n492 B.n491 10.6151
R1971 B.n493 B.n492 10.6151
R1972 B.n493 B.n236 10.6151
R1973 B.n497 B.n236 10.6151
R1974 B.n498 B.n497 10.6151
R1975 B.n499 B.n498 10.6151
R1976 B.n499 B.n234 10.6151
R1977 B.n503 B.n234 10.6151
R1978 B.n504 B.n503 10.6151
R1979 B.n505 B.n504 10.6151
R1980 B.n505 B.n232 10.6151
R1981 B.n509 B.n232 10.6151
R1982 B.n512 B.n511 10.6151
R1983 B.n512 B.n228 10.6151
R1984 B.n516 B.n228 10.6151
R1985 B.n517 B.n516 10.6151
R1986 B.n518 B.n517 10.6151
R1987 B.n518 B.n226 10.6151
R1988 B.n522 B.n226 10.6151
R1989 B.n523 B.n522 10.6151
R1990 B.n524 B.n523 10.6151
R1991 B.n528 B.n527 10.6151
R1992 B.n529 B.n528 10.6151
R1993 B.n529 B.n220 10.6151
R1994 B.n533 B.n220 10.6151
R1995 B.n534 B.n533 10.6151
R1996 B.n535 B.n534 10.6151
R1997 B.n535 B.n218 10.6151
R1998 B.n539 B.n218 10.6151
R1999 B.n540 B.n539 10.6151
R2000 B.n541 B.n540 10.6151
R2001 B.n541 B.n216 10.6151
R2002 B.n545 B.n216 10.6151
R2003 B.n546 B.n545 10.6151
R2004 B.n547 B.n546 10.6151
R2005 B.n547 B.n214 10.6151
R2006 B.n551 B.n214 10.6151
R2007 B.n552 B.n551 10.6151
R2008 B.n553 B.n552 10.6151
R2009 B.n553 B.n212 10.6151
R2010 B.n557 B.n212 10.6151
R2011 B.n558 B.n557 10.6151
R2012 B.n559 B.n558 10.6151
R2013 B.n559 B.n210 10.6151
R2014 B.n563 B.n210 10.6151
R2015 B.n564 B.n563 10.6151
R2016 B.n565 B.n564 10.6151
R2017 B.n565 B.n208 10.6151
R2018 B.n569 B.n208 10.6151
R2019 B.n570 B.n569 10.6151
R2020 B.n571 B.n570 10.6151
R2021 B.n571 B.n206 10.6151
R2022 B.n575 B.n206 10.6151
R2023 B.n576 B.n575 10.6151
R2024 B.n577 B.n576 10.6151
R2025 B.n577 B.n204 10.6151
R2026 B.n581 B.n204 10.6151
R2027 B.n582 B.n581 10.6151
R2028 B.n583 B.n582 10.6151
R2029 B.n583 B.n202 10.6151
R2030 B.n587 B.n202 10.6151
R2031 B.n588 B.n587 10.6151
R2032 B.n589 B.n588 10.6151
R2033 B.n589 B.n200 10.6151
R2034 B.n593 B.n200 10.6151
R2035 B.n594 B.n593 10.6151
R2036 B.n595 B.n594 10.6151
R2037 B.n595 B.n198 10.6151
R2038 B.n599 B.n198 10.6151
R2039 B.n600 B.n599 10.6151
R2040 B.n601 B.n600 10.6151
R2041 B.n601 B.n196 10.6151
R2042 B.n605 B.n196 10.6151
R2043 B.n606 B.n605 10.6151
R2044 B.n607 B.n606 10.6151
R2045 B.n607 B.n194 10.6151
R2046 B.n611 B.n194 10.6151
R2047 B.n612 B.n611 10.6151
R2048 B.n613 B.n612 10.6151
R2049 B.n613 B.n192 10.6151
R2050 B.n617 B.n192 10.6151
R2051 B.n415 B.n262 10.6151
R2052 B.n415 B.n414 10.6151
R2053 B.n414 B.n413 10.6151
R2054 B.n413 B.n264 10.6151
R2055 B.n409 B.n264 10.6151
R2056 B.n409 B.n408 10.6151
R2057 B.n408 B.n407 10.6151
R2058 B.n407 B.n266 10.6151
R2059 B.n403 B.n266 10.6151
R2060 B.n403 B.n402 10.6151
R2061 B.n402 B.n401 10.6151
R2062 B.n401 B.n268 10.6151
R2063 B.n397 B.n268 10.6151
R2064 B.n397 B.n396 10.6151
R2065 B.n396 B.n395 10.6151
R2066 B.n395 B.n270 10.6151
R2067 B.n391 B.n270 10.6151
R2068 B.n391 B.n390 10.6151
R2069 B.n390 B.n389 10.6151
R2070 B.n389 B.n272 10.6151
R2071 B.n385 B.n272 10.6151
R2072 B.n385 B.n384 10.6151
R2073 B.n384 B.n383 10.6151
R2074 B.n383 B.n274 10.6151
R2075 B.n379 B.n274 10.6151
R2076 B.n379 B.n378 10.6151
R2077 B.n378 B.n377 10.6151
R2078 B.n377 B.n276 10.6151
R2079 B.n373 B.n276 10.6151
R2080 B.n373 B.n372 10.6151
R2081 B.n372 B.n371 10.6151
R2082 B.n371 B.n278 10.6151
R2083 B.n367 B.n278 10.6151
R2084 B.n367 B.n366 10.6151
R2085 B.n366 B.n365 10.6151
R2086 B.n365 B.n280 10.6151
R2087 B.n361 B.n280 10.6151
R2088 B.n361 B.n360 10.6151
R2089 B.n360 B.n359 10.6151
R2090 B.n359 B.n282 10.6151
R2091 B.n355 B.n282 10.6151
R2092 B.n355 B.n354 10.6151
R2093 B.n354 B.n353 10.6151
R2094 B.n353 B.n284 10.6151
R2095 B.n349 B.n284 10.6151
R2096 B.n349 B.n348 10.6151
R2097 B.n348 B.n347 10.6151
R2098 B.n347 B.n286 10.6151
R2099 B.n343 B.n286 10.6151
R2100 B.n343 B.n342 10.6151
R2101 B.n342 B.n341 10.6151
R2102 B.n341 B.n288 10.6151
R2103 B.n337 B.n288 10.6151
R2104 B.n337 B.n336 10.6151
R2105 B.n336 B.n335 10.6151
R2106 B.n335 B.n290 10.6151
R2107 B.n331 B.n290 10.6151
R2108 B.n331 B.n330 10.6151
R2109 B.n330 B.n329 10.6151
R2110 B.n329 B.n292 10.6151
R2111 B.n325 B.n292 10.6151
R2112 B.n325 B.n324 10.6151
R2113 B.n324 B.n323 10.6151
R2114 B.n323 B.n294 10.6151
R2115 B.n319 B.n294 10.6151
R2116 B.n319 B.n318 10.6151
R2117 B.n318 B.n317 10.6151
R2118 B.n317 B.n296 10.6151
R2119 B.n313 B.n296 10.6151
R2120 B.n313 B.n312 10.6151
R2121 B.n312 B.n311 10.6151
R2122 B.n311 B.n298 10.6151
R2123 B.n307 B.n298 10.6151
R2124 B.n307 B.n306 10.6151
R2125 B.n306 B.n305 10.6151
R2126 B.n305 B.n300 10.6151
R2127 B.n301 B.n300 10.6151
R2128 B.n301 B.n0 10.6151
R2129 B.n1171 B.n1 10.6151
R2130 B.n1171 B.n1170 10.6151
R2131 B.n1170 B.n1169 10.6151
R2132 B.n1169 B.n4 10.6151
R2133 B.n1165 B.n4 10.6151
R2134 B.n1165 B.n1164 10.6151
R2135 B.n1164 B.n1163 10.6151
R2136 B.n1163 B.n6 10.6151
R2137 B.n1159 B.n6 10.6151
R2138 B.n1159 B.n1158 10.6151
R2139 B.n1158 B.n1157 10.6151
R2140 B.n1157 B.n8 10.6151
R2141 B.n1153 B.n8 10.6151
R2142 B.n1153 B.n1152 10.6151
R2143 B.n1152 B.n1151 10.6151
R2144 B.n1151 B.n10 10.6151
R2145 B.n1147 B.n10 10.6151
R2146 B.n1147 B.n1146 10.6151
R2147 B.n1146 B.n1145 10.6151
R2148 B.n1145 B.n12 10.6151
R2149 B.n1141 B.n12 10.6151
R2150 B.n1141 B.n1140 10.6151
R2151 B.n1140 B.n1139 10.6151
R2152 B.n1139 B.n14 10.6151
R2153 B.n1135 B.n14 10.6151
R2154 B.n1135 B.n1134 10.6151
R2155 B.n1134 B.n1133 10.6151
R2156 B.n1133 B.n16 10.6151
R2157 B.n1129 B.n16 10.6151
R2158 B.n1129 B.n1128 10.6151
R2159 B.n1128 B.n1127 10.6151
R2160 B.n1127 B.n18 10.6151
R2161 B.n1123 B.n18 10.6151
R2162 B.n1123 B.n1122 10.6151
R2163 B.n1122 B.n1121 10.6151
R2164 B.n1121 B.n20 10.6151
R2165 B.n1117 B.n20 10.6151
R2166 B.n1117 B.n1116 10.6151
R2167 B.n1116 B.n1115 10.6151
R2168 B.n1115 B.n22 10.6151
R2169 B.n1111 B.n22 10.6151
R2170 B.n1111 B.n1110 10.6151
R2171 B.n1110 B.n1109 10.6151
R2172 B.n1109 B.n24 10.6151
R2173 B.n1105 B.n24 10.6151
R2174 B.n1105 B.n1104 10.6151
R2175 B.n1104 B.n1103 10.6151
R2176 B.n1103 B.n26 10.6151
R2177 B.n1099 B.n26 10.6151
R2178 B.n1099 B.n1098 10.6151
R2179 B.n1098 B.n1097 10.6151
R2180 B.n1097 B.n28 10.6151
R2181 B.n1093 B.n28 10.6151
R2182 B.n1093 B.n1092 10.6151
R2183 B.n1092 B.n1091 10.6151
R2184 B.n1091 B.n30 10.6151
R2185 B.n1087 B.n30 10.6151
R2186 B.n1087 B.n1086 10.6151
R2187 B.n1086 B.n1085 10.6151
R2188 B.n1085 B.n32 10.6151
R2189 B.n1081 B.n32 10.6151
R2190 B.n1081 B.n1080 10.6151
R2191 B.n1080 B.n1079 10.6151
R2192 B.n1079 B.n34 10.6151
R2193 B.n1075 B.n34 10.6151
R2194 B.n1075 B.n1074 10.6151
R2195 B.n1074 B.n1073 10.6151
R2196 B.n1073 B.n36 10.6151
R2197 B.n1069 B.n36 10.6151
R2198 B.n1069 B.n1068 10.6151
R2199 B.n1068 B.n1067 10.6151
R2200 B.n1067 B.n38 10.6151
R2201 B.n1063 B.n38 10.6151
R2202 B.n1063 B.n1062 10.6151
R2203 B.n1062 B.n1061 10.6151
R2204 B.n1061 B.n40 10.6151
R2205 B.n1057 B.n40 10.6151
R2206 B.n1057 B.n1056 10.6151
R2207 B.n965 B.n74 9.36635
R2208 B.n948 B.n947 9.36635
R2209 B.n510 B.n509 9.36635
R2210 B.n527 B.n224 9.36635
R2211 B.n1175 B.n0 2.81026
R2212 B.n1175 B.n1 2.81026
R2213 B.n962 B.n74 1.24928
R2214 B.n949 B.n948 1.24928
R2215 B.n511 B.n510 1.24928
R2216 B.n524 B.n224 1.24928
C0 VDD2 VTAIL 13.5782f
C1 VDD2 VP 0.72356f
C2 w_n5806_n4686# VDD1 3.64854f
C3 VDD2 VN 17.260199f
C4 VTAIL VDD1 13.52f
C5 w_n5806_n4686# VTAIL 4.24641f
C6 VDD1 VP 17.823801f
C7 w_n5806_n4686# VP 13.648f
C8 VDD1 VN 0.155558f
C9 w_n5806_n4686# VN 12.8887f
C10 VTAIL VP 18.073599f
C11 VTAIL VN 18.0589f
C12 VP VN 11.2432f
C13 B VDD2 3.59999f
C14 B VDD1 3.43924f
C15 w_n5806_n4686# B 14.243599f
C16 B VTAIL 5.71505f
C17 B VP 2.92345f
C18 VDD2 VDD1 2.88936f
C19 w_n5806_n4686# VDD2 3.84926f
C20 B VN 1.64056f
C21 VDD2 VSUBS 2.69265f
C22 VDD1 VSUBS 2.578737f
C23 VTAIL VSUBS 1.786101f
C24 VN VSUBS 9.726939f
C25 VP VSUBS 5.872422f
C26 B VSUBS 7.2858f
C27 w_n5806_n4686# VSUBS 0.332544p
C28 B.n0 VSUBS 0.004721f
C29 B.n1 VSUBS 0.004721f
C30 B.n2 VSUBS 0.007467f
C31 B.n3 VSUBS 0.007467f
C32 B.n4 VSUBS 0.007467f
C33 B.n5 VSUBS 0.007467f
C34 B.n6 VSUBS 0.007467f
C35 B.n7 VSUBS 0.007467f
C36 B.n8 VSUBS 0.007467f
C37 B.n9 VSUBS 0.007467f
C38 B.n10 VSUBS 0.007467f
C39 B.n11 VSUBS 0.007467f
C40 B.n12 VSUBS 0.007467f
C41 B.n13 VSUBS 0.007467f
C42 B.n14 VSUBS 0.007467f
C43 B.n15 VSUBS 0.007467f
C44 B.n16 VSUBS 0.007467f
C45 B.n17 VSUBS 0.007467f
C46 B.n18 VSUBS 0.007467f
C47 B.n19 VSUBS 0.007467f
C48 B.n20 VSUBS 0.007467f
C49 B.n21 VSUBS 0.007467f
C50 B.n22 VSUBS 0.007467f
C51 B.n23 VSUBS 0.007467f
C52 B.n24 VSUBS 0.007467f
C53 B.n25 VSUBS 0.007467f
C54 B.n26 VSUBS 0.007467f
C55 B.n27 VSUBS 0.007467f
C56 B.n28 VSUBS 0.007467f
C57 B.n29 VSUBS 0.007467f
C58 B.n30 VSUBS 0.007467f
C59 B.n31 VSUBS 0.007467f
C60 B.n32 VSUBS 0.007467f
C61 B.n33 VSUBS 0.007467f
C62 B.n34 VSUBS 0.007467f
C63 B.n35 VSUBS 0.007467f
C64 B.n36 VSUBS 0.007467f
C65 B.n37 VSUBS 0.007467f
C66 B.n38 VSUBS 0.007467f
C67 B.n39 VSUBS 0.007467f
C68 B.n40 VSUBS 0.007467f
C69 B.n41 VSUBS 0.016715f
C70 B.n42 VSUBS 0.007467f
C71 B.n43 VSUBS 0.007467f
C72 B.n44 VSUBS 0.007467f
C73 B.n45 VSUBS 0.007467f
C74 B.n46 VSUBS 0.007467f
C75 B.n47 VSUBS 0.007467f
C76 B.n48 VSUBS 0.007467f
C77 B.n49 VSUBS 0.007467f
C78 B.n50 VSUBS 0.007467f
C79 B.n51 VSUBS 0.007467f
C80 B.n52 VSUBS 0.007467f
C81 B.n53 VSUBS 0.007467f
C82 B.n54 VSUBS 0.007467f
C83 B.n55 VSUBS 0.007467f
C84 B.n56 VSUBS 0.007467f
C85 B.n57 VSUBS 0.007467f
C86 B.n58 VSUBS 0.007467f
C87 B.n59 VSUBS 0.007467f
C88 B.n60 VSUBS 0.007467f
C89 B.n61 VSUBS 0.007467f
C90 B.n62 VSUBS 0.007467f
C91 B.n63 VSUBS 0.007467f
C92 B.n64 VSUBS 0.007467f
C93 B.n65 VSUBS 0.007467f
C94 B.n66 VSUBS 0.007467f
C95 B.n67 VSUBS 0.007467f
C96 B.n68 VSUBS 0.007467f
C97 B.n69 VSUBS 0.007467f
C98 B.n70 VSUBS 0.007467f
C99 B.n71 VSUBS 0.007467f
C100 B.t11 VSUBS 0.670923f
C101 B.t10 VSUBS 0.70038f
C102 B.t9 VSUBS 3.33046f
C103 B.n72 VSUBS 0.436812f
C104 B.n73 VSUBS 0.081784f
C105 B.n74 VSUBS 0.017299f
C106 B.n75 VSUBS 0.007467f
C107 B.n76 VSUBS 0.007467f
C108 B.n77 VSUBS 0.007467f
C109 B.n78 VSUBS 0.007467f
C110 B.n79 VSUBS 0.007467f
C111 B.t2 VSUBS 0.670898f
C112 B.t1 VSUBS 0.700361f
C113 B.t0 VSUBS 3.33046f
C114 B.n80 VSUBS 0.436831f
C115 B.n81 VSUBS 0.08181f
C116 B.n82 VSUBS 0.007467f
C117 B.n83 VSUBS 0.007467f
C118 B.n84 VSUBS 0.007467f
C119 B.n85 VSUBS 0.007467f
C120 B.n86 VSUBS 0.007467f
C121 B.n87 VSUBS 0.007467f
C122 B.n88 VSUBS 0.007467f
C123 B.n89 VSUBS 0.007467f
C124 B.n90 VSUBS 0.007467f
C125 B.n91 VSUBS 0.007467f
C126 B.n92 VSUBS 0.007467f
C127 B.n93 VSUBS 0.007467f
C128 B.n94 VSUBS 0.007467f
C129 B.n95 VSUBS 0.007467f
C130 B.n96 VSUBS 0.007467f
C131 B.n97 VSUBS 0.007467f
C132 B.n98 VSUBS 0.007467f
C133 B.n99 VSUBS 0.007467f
C134 B.n100 VSUBS 0.007467f
C135 B.n101 VSUBS 0.007467f
C136 B.n102 VSUBS 0.007467f
C137 B.n103 VSUBS 0.007467f
C138 B.n104 VSUBS 0.007467f
C139 B.n105 VSUBS 0.007467f
C140 B.n106 VSUBS 0.007467f
C141 B.n107 VSUBS 0.007467f
C142 B.n108 VSUBS 0.007467f
C143 B.n109 VSUBS 0.007467f
C144 B.n110 VSUBS 0.007467f
C145 B.n111 VSUBS 0.007467f
C146 B.n112 VSUBS 0.017598f
C147 B.n113 VSUBS 0.007467f
C148 B.n114 VSUBS 0.007467f
C149 B.n115 VSUBS 0.007467f
C150 B.n116 VSUBS 0.007467f
C151 B.n117 VSUBS 0.007467f
C152 B.n118 VSUBS 0.007467f
C153 B.n119 VSUBS 0.007467f
C154 B.n120 VSUBS 0.007467f
C155 B.n121 VSUBS 0.007467f
C156 B.n122 VSUBS 0.007467f
C157 B.n123 VSUBS 0.007467f
C158 B.n124 VSUBS 0.007467f
C159 B.n125 VSUBS 0.007467f
C160 B.n126 VSUBS 0.007467f
C161 B.n127 VSUBS 0.007467f
C162 B.n128 VSUBS 0.007467f
C163 B.n129 VSUBS 0.007467f
C164 B.n130 VSUBS 0.007467f
C165 B.n131 VSUBS 0.007467f
C166 B.n132 VSUBS 0.007467f
C167 B.n133 VSUBS 0.007467f
C168 B.n134 VSUBS 0.007467f
C169 B.n135 VSUBS 0.007467f
C170 B.n136 VSUBS 0.007467f
C171 B.n137 VSUBS 0.007467f
C172 B.n138 VSUBS 0.007467f
C173 B.n139 VSUBS 0.007467f
C174 B.n140 VSUBS 0.007467f
C175 B.n141 VSUBS 0.007467f
C176 B.n142 VSUBS 0.007467f
C177 B.n143 VSUBS 0.007467f
C178 B.n144 VSUBS 0.007467f
C179 B.n145 VSUBS 0.007467f
C180 B.n146 VSUBS 0.007467f
C181 B.n147 VSUBS 0.007467f
C182 B.n148 VSUBS 0.007467f
C183 B.n149 VSUBS 0.007467f
C184 B.n150 VSUBS 0.007467f
C185 B.n151 VSUBS 0.007467f
C186 B.n152 VSUBS 0.007467f
C187 B.n153 VSUBS 0.007467f
C188 B.n154 VSUBS 0.007467f
C189 B.n155 VSUBS 0.007467f
C190 B.n156 VSUBS 0.007467f
C191 B.n157 VSUBS 0.007467f
C192 B.n158 VSUBS 0.007467f
C193 B.n159 VSUBS 0.007467f
C194 B.n160 VSUBS 0.007467f
C195 B.n161 VSUBS 0.007467f
C196 B.n162 VSUBS 0.007467f
C197 B.n163 VSUBS 0.007467f
C198 B.n164 VSUBS 0.007467f
C199 B.n165 VSUBS 0.007467f
C200 B.n166 VSUBS 0.007467f
C201 B.n167 VSUBS 0.007467f
C202 B.n168 VSUBS 0.007467f
C203 B.n169 VSUBS 0.007467f
C204 B.n170 VSUBS 0.007467f
C205 B.n171 VSUBS 0.007467f
C206 B.n172 VSUBS 0.007467f
C207 B.n173 VSUBS 0.007467f
C208 B.n174 VSUBS 0.007467f
C209 B.n175 VSUBS 0.007467f
C210 B.n176 VSUBS 0.007467f
C211 B.n177 VSUBS 0.007467f
C212 B.n178 VSUBS 0.007467f
C213 B.n179 VSUBS 0.007467f
C214 B.n180 VSUBS 0.007467f
C215 B.n181 VSUBS 0.007467f
C216 B.n182 VSUBS 0.007467f
C217 B.n183 VSUBS 0.007467f
C218 B.n184 VSUBS 0.007467f
C219 B.n185 VSUBS 0.007467f
C220 B.n186 VSUBS 0.007467f
C221 B.n187 VSUBS 0.007467f
C222 B.n188 VSUBS 0.007467f
C223 B.n189 VSUBS 0.007467f
C224 B.n190 VSUBS 0.007467f
C225 B.n191 VSUBS 0.016715f
C226 B.n192 VSUBS 0.007467f
C227 B.n193 VSUBS 0.007467f
C228 B.n194 VSUBS 0.007467f
C229 B.n195 VSUBS 0.007467f
C230 B.n196 VSUBS 0.007467f
C231 B.n197 VSUBS 0.007467f
C232 B.n198 VSUBS 0.007467f
C233 B.n199 VSUBS 0.007467f
C234 B.n200 VSUBS 0.007467f
C235 B.n201 VSUBS 0.007467f
C236 B.n202 VSUBS 0.007467f
C237 B.n203 VSUBS 0.007467f
C238 B.n204 VSUBS 0.007467f
C239 B.n205 VSUBS 0.007467f
C240 B.n206 VSUBS 0.007467f
C241 B.n207 VSUBS 0.007467f
C242 B.n208 VSUBS 0.007467f
C243 B.n209 VSUBS 0.007467f
C244 B.n210 VSUBS 0.007467f
C245 B.n211 VSUBS 0.007467f
C246 B.n212 VSUBS 0.007467f
C247 B.n213 VSUBS 0.007467f
C248 B.n214 VSUBS 0.007467f
C249 B.n215 VSUBS 0.007467f
C250 B.n216 VSUBS 0.007467f
C251 B.n217 VSUBS 0.007467f
C252 B.n218 VSUBS 0.007467f
C253 B.n219 VSUBS 0.007467f
C254 B.n220 VSUBS 0.007467f
C255 B.n221 VSUBS 0.007467f
C256 B.t7 VSUBS 0.670898f
C257 B.t8 VSUBS 0.700361f
C258 B.t6 VSUBS 3.33046f
C259 B.n222 VSUBS 0.436831f
C260 B.n223 VSUBS 0.08181f
C261 B.n224 VSUBS 0.017299f
C262 B.n225 VSUBS 0.007467f
C263 B.n226 VSUBS 0.007467f
C264 B.n227 VSUBS 0.007467f
C265 B.n228 VSUBS 0.007467f
C266 B.n229 VSUBS 0.007467f
C267 B.t4 VSUBS 0.670923f
C268 B.t5 VSUBS 0.70038f
C269 B.t3 VSUBS 3.33046f
C270 B.n230 VSUBS 0.436812f
C271 B.n231 VSUBS 0.081784f
C272 B.n232 VSUBS 0.007467f
C273 B.n233 VSUBS 0.007467f
C274 B.n234 VSUBS 0.007467f
C275 B.n235 VSUBS 0.007467f
C276 B.n236 VSUBS 0.007467f
C277 B.n237 VSUBS 0.007467f
C278 B.n238 VSUBS 0.007467f
C279 B.n239 VSUBS 0.007467f
C280 B.n240 VSUBS 0.007467f
C281 B.n241 VSUBS 0.007467f
C282 B.n242 VSUBS 0.007467f
C283 B.n243 VSUBS 0.007467f
C284 B.n244 VSUBS 0.007467f
C285 B.n245 VSUBS 0.007467f
C286 B.n246 VSUBS 0.007467f
C287 B.n247 VSUBS 0.007467f
C288 B.n248 VSUBS 0.007467f
C289 B.n249 VSUBS 0.007467f
C290 B.n250 VSUBS 0.007467f
C291 B.n251 VSUBS 0.007467f
C292 B.n252 VSUBS 0.007467f
C293 B.n253 VSUBS 0.007467f
C294 B.n254 VSUBS 0.007467f
C295 B.n255 VSUBS 0.007467f
C296 B.n256 VSUBS 0.007467f
C297 B.n257 VSUBS 0.007467f
C298 B.n258 VSUBS 0.007467f
C299 B.n259 VSUBS 0.007467f
C300 B.n260 VSUBS 0.007467f
C301 B.n261 VSUBS 0.007467f
C302 B.n262 VSUBS 0.016715f
C303 B.n263 VSUBS 0.007467f
C304 B.n264 VSUBS 0.007467f
C305 B.n265 VSUBS 0.007467f
C306 B.n266 VSUBS 0.007467f
C307 B.n267 VSUBS 0.007467f
C308 B.n268 VSUBS 0.007467f
C309 B.n269 VSUBS 0.007467f
C310 B.n270 VSUBS 0.007467f
C311 B.n271 VSUBS 0.007467f
C312 B.n272 VSUBS 0.007467f
C313 B.n273 VSUBS 0.007467f
C314 B.n274 VSUBS 0.007467f
C315 B.n275 VSUBS 0.007467f
C316 B.n276 VSUBS 0.007467f
C317 B.n277 VSUBS 0.007467f
C318 B.n278 VSUBS 0.007467f
C319 B.n279 VSUBS 0.007467f
C320 B.n280 VSUBS 0.007467f
C321 B.n281 VSUBS 0.007467f
C322 B.n282 VSUBS 0.007467f
C323 B.n283 VSUBS 0.007467f
C324 B.n284 VSUBS 0.007467f
C325 B.n285 VSUBS 0.007467f
C326 B.n286 VSUBS 0.007467f
C327 B.n287 VSUBS 0.007467f
C328 B.n288 VSUBS 0.007467f
C329 B.n289 VSUBS 0.007467f
C330 B.n290 VSUBS 0.007467f
C331 B.n291 VSUBS 0.007467f
C332 B.n292 VSUBS 0.007467f
C333 B.n293 VSUBS 0.007467f
C334 B.n294 VSUBS 0.007467f
C335 B.n295 VSUBS 0.007467f
C336 B.n296 VSUBS 0.007467f
C337 B.n297 VSUBS 0.007467f
C338 B.n298 VSUBS 0.007467f
C339 B.n299 VSUBS 0.007467f
C340 B.n300 VSUBS 0.007467f
C341 B.n301 VSUBS 0.007467f
C342 B.n302 VSUBS 0.007467f
C343 B.n303 VSUBS 0.007467f
C344 B.n304 VSUBS 0.007467f
C345 B.n305 VSUBS 0.007467f
C346 B.n306 VSUBS 0.007467f
C347 B.n307 VSUBS 0.007467f
C348 B.n308 VSUBS 0.007467f
C349 B.n309 VSUBS 0.007467f
C350 B.n310 VSUBS 0.007467f
C351 B.n311 VSUBS 0.007467f
C352 B.n312 VSUBS 0.007467f
C353 B.n313 VSUBS 0.007467f
C354 B.n314 VSUBS 0.007467f
C355 B.n315 VSUBS 0.007467f
C356 B.n316 VSUBS 0.007467f
C357 B.n317 VSUBS 0.007467f
C358 B.n318 VSUBS 0.007467f
C359 B.n319 VSUBS 0.007467f
C360 B.n320 VSUBS 0.007467f
C361 B.n321 VSUBS 0.007467f
C362 B.n322 VSUBS 0.007467f
C363 B.n323 VSUBS 0.007467f
C364 B.n324 VSUBS 0.007467f
C365 B.n325 VSUBS 0.007467f
C366 B.n326 VSUBS 0.007467f
C367 B.n327 VSUBS 0.007467f
C368 B.n328 VSUBS 0.007467f
C369 B.n329 VSUBS 0.007467f
C370 B.n330 VSUBS 0.007467f
C371 B.n331 VSUBS 0.007467f
C372 B.n332 VSUBS 0.007467f
C373 B.n333 VSUBS 0.007467f
C374 B.n334 VSUBS 0.007467f
C375 B.n335 VSUBS 0.007467f
C376 B.n336 VSUBS 0.007467f
C377 B.n337 VSUBS 0.007467f
C378 B.n338 VSUBS 0.007467f
C379 B.n339 VSUBS 0.007467f
C380 B.n340 VSUBS 0.007467f
C381 B.n341 VSUBS 0.007467f
C382 B.n342 VSUBS 0.007467f
C383 B.n343 VSUBS 0.007467f
C384 B.n344 VSUBS 0.007467f
C385 B.n345 VSUBS 0.007467f
C386 B.n346 VSUBS 0.007467f
C387 B.n347 VSUBS 0.007467f
C388 B.n348 VSUBS 0.007467f
C389 B.n349 VSUBS 0.007467f
C390 B.n350 VSUBS 0.007467f
C391 B.n351 VSUBS 0.007467f
C392 B.n352 VSUBS 0.007467f
C393 B.n353 VSUBS 0.007467f
C394 B.n354 VSUBS 0.007467f
C395 B.n355 VSUBS 0.007467f
C396 B.n356 VSUBS 0.007467f
C397 B.n357 VSUBS 0.007467f
C398 B.n358 VSUBS 0.007467f
C399 B.n359 VSUBS 0.007467f
C400 B.n360 VSUBS 0.007467f
C401 B.n361 VSUBS 0.007467f
C402 B.n362 VSUBS 0.007467f
C403 B.n363 VSUBS 0.007467f
C404 B.n364 VSUBS 0.007467f
C405 B.n365 VSUBS 0.007467f
C406 B.n366 VSUBS 0.007467f
C407 B.n367 VSUBS 0.007467f
C408 B.n368 VSUBS 0.007467f
C409 B.n369 VSUBS 0.007467f
C410 B.n370 VSUBS 0.007467f
C411 B.n371 VSUBS 0.007467f
C412 B.n372 VSUBS 0.007467f
C413 B.n373 VSUBS 0.007467f
C414 B.n374 VSUBS 0.007467f
C415 B.n375 VSUBS 0.007467f
C416 B.n376 VSUBS 0.007467f
C417 B.n377 VSUBS 0.007467f
C418 B.n378 VSUBS 0.007467f
C419 B.n379 VSUBS 0.007467f
C420 B.n380 VSUBS 0.007467f
C421 B.n381 VSUBS 0.007467f
C422 B.n382 VSUBS 0.007467f
C423 B.n383 VSUBS 0.007467f
C424 B.n384 VSUBS 0.007467f
C425 B.n385 VSUBS 0.007467f
C426 B.n386 VSUBS 0.007467f
C427 B.n387 VSUBS 0.007467f
C428 B.n388 VSUBS 0.007467f
C429 B.n389 VSUBS 0.007467f
C430 B.n390 VSUBS 0.007467f
C431 B.n391 VSUBS 0.007467f
C432 B.n392 VSUBS 0.007467f
C433 B.n393 VSUBS 0.007467f
C434 B.n394 VSUBS 0.007467f
C435 B.n395 VSUBS 0.007467f
C436 B.n396 VSUBS 0.007467f
C437 B.n397 VSUBS 0.007467f
C438 B.n398 VSUBS 0.007467f
C439 B.n399 VSUBS 0.007467f
C440 B.n400 VSUBS 0.007467f
C441 B.n401 VSUBS 0.007467f
C442 B.n402 VSUBS 0.007467f
C443 B.n403 VSUBS 0.007467f
C444 B.n404 VSUBS 0.007467f
C445 B.n405 VSUBS 0.007467f
C446 B.n406 VSUBS 0.007467f
C447 B.n407 VSUBS 0.007467f
C448 B.n408 VSUBS 0.007467f
C449 B.n409 VSUBS 0.007467f
C450 B.n410 VSUBS 0.007467f
C451 B.n411 VSUBS 0.007467f
C452 B.n412 VSUBS 0.007467f
C453 B.n413 VSUBS 0.007467f
C454 B.n414 VSUBS 0.007467f
C455 B.n415 VSUBS 0.007467f
C456 B.n416 VSUBS 0.007467f
C457 B.n417 VSUBS 0.016715f
C458 B.n418 VSUBS 0.018202f
C459 B.n419 VSUBS 0.018202f
C460 B.n420 VSUBS 0.007467f
C461 B.n421 VSUBS 0.007467f
C462 B.n422 VSUBS 0.007467f
C463 B.n423 VSUBS 0.007467f
C464 B.n424 VSUBS 0.007467f
C465 B.n425 VSUBS 0.007467f
C466 B.n426 VSUBS 0.007467f
C467 B.n427 VSUBS 0.007467f
C468 B.n428 VSUBS 0.007467f
C469 B.n429 VSUBS 0.007467f
C470 B.n430 VSUBS 0.007467f
C471 B.n431 VSUBS 0.007467f
C472 B.n432 VSUBS 0.007467f
C473 B.n433 VSUBS 0.007467f
C474 B.n434 VSUBS 0.007467f
C475 B.n435 VSUBS 0.007467f
C476 B.n436 VSUBS 0.007467f
C477 B.n437 VSUBS 0.007467f
C478 B.n438 VSUBS 0.007467f
C479 B.n439 VSUBS 0.007467f
C480 B.n440 VSUBS 0.007467f
C481 B.n441 VSUBS 0.007467f
C482 B.n442 VSUBS 0.007467f
C483 B.n443 VSUBS 0.007467f
C484 B.n444 VSUBS 0.007467f
C485 B.n445 VSUBS 0.007467f
C486 B.n446 VSUBS 0.007467f
C487 B.n447 VSUBS 0.007467f
C488 B.n448 VSUBS 0.007467f
C489 B.n449 VSUBS 0.007467f
C490 B.n450 VSUBS 0.007467f
C491 B.n451 VSUBS 0.007467f
C492 B.n452 VSUBS 0.007467f
C493 B.n453 VSUBS 0.007467f
C494 B.n454 VSUBS 0.007467f
C495 B.n455 VSUBS 0.007467f
C496 B.n456 VSUBS 0.007467f
C497 B.n457 VSUBS 0.007467f
C498 B.n458 VSUBS 0.007467f
C499 B.n459 VSUBS 0.007467f
C500 B.n460 VSUBS 0.007467f
C501 B.n461 VSUBS 0.007467f
C502 B.n462 VSUBS 0.007467f
C503 B.n463 VSUBS 0.007467f
C504 B.n464 VSUBS 0.007467f
C505 B.n465 VSUBS 0.007467f
C506 B.n466 VSUBS 0.007467f
C507 B.n467 VSUBS 0.007467f
C508 B.n468 VSUBS 0.007467f
C509 B.n469 VSUBS 0.007467f
C510 B.n470 VSUBS 0.007467f
C511 B.n471 VSUBS 0.007467f
C512 B.n472 VSUBS 0.007467f
C513 B.n473 VSUBS 0.007467f
C514 B.n474 VSUBS 0.007467f
C515 B.n475 VSUBS 0.007467f
C516 B.n476 VSUBS 0.007467f
C517 B.n477 VSUBS 0.007467f
C518 B.n478 VSUBS 0.007467f
C519 B.n479 VSUBS 0.007467f
C520 B.n480 VSUBS 0.007467f
C521 B.n481 VSUBS 0.007467f
C522 B.n482 VSUBS 0.007467f
C523 B.n483 VSUBS 0.007467f
C524 B.n484 VSUBS 0.007467f
C525 B.n485 VSUBS 0.007467f
C526 B.n486 VSUBS 0.007467f
C527 B.n487 VSUBS 0.007467f
C528 B.n488 VSUBS 0.007467f
C529 B.n489 VSUBS 0.007467f
C530 B.n490 VSUBS 0.007467f
C531 B.n491 VSUBS 0.007467f
C532 B.n492 VSUBS 0.007467f
C533 B.n493 VSUBS 0.007467f
C534 B.n494 VSUBS 0.007467f
C535 B.n495 VSUBS 0.007467f
C536 B.n496 VSUBS 0.007467f
C537 B.n497 VSUBS 0.007467f
C538 B.n498 VSUBS 0.007467f
C539 B.n499 VSUBS 0.007467f
C540 B.n500 VSUBS 0.007467f
C541 B.n501 VSUBS 0.007467f
C542 B.n502 VSUBS 0.007467f
C543 B.n503 VSUBS 0.007467f
C544 B.n504 VSUBS 0.007467f
C545 B.n505 VSUBS 0.007467f
C546 B.n506 VSUBS 0.007467f
C547 B.n507 VSUBS 0.007467f
C548 B.n508 VSUBS 0.007467f
C549 B.n509 VSUBS 0.007027f
C550 B.n510 VSUBS 0.017299f
C551 B.n511 VSUBS 0.004172f
C552 B.n512 VSUBS 0.007467f
C553 B.n513 VSUBS 0.007467f
C554 B.n514 VSUBS 0.007467f
C555 B.n515 VSUBS 0.007467f
C556 B.n516 VSUBS 0.007467f
C557 B.n517 VSUBS 0.007467f
C558 B.n518 VSUBS 0.007467f
C559 B.n519 VSUBS 0.007467f
C560 B.n520 VSUBS 0.007467f
C561 B.n521 VSUBS 0.007467f
C562 B.n522 VSUBS 0.007467f
C563 B.n523 VSUBS 0.007467f
C564 B.n524 VSUBS 0.004172f
C565 B.n525 VSUBS 0.007467f
C566 B.n526 VSUBS 0.007467f
C567 B.n527 VSUBS 0.007027f
C568 B.n528 VSUBS 0.007467f
C569 B.n529 VSUBS 0.007467f
C570 B.n530 VSUBS 0.007467f
C571 B.n531 VSUBS 0.007467f
C572 B.n532 VSUBS 0.007467f
C573 B.n533 VSUBS 0.007467f
C574 B.n534 VSUBS 0.007467f
C575 B.n535 VSUBS 0.007467f
C576 B.n536 VSUBS 0.007467f
C577 B.n537 VSUBS 0.007467f
C578 B.n538 VSUBS 0.007467f
C579 B.n539 VSUBS 0.007467f
C580 B.n540 VSUBS 0.007467f
C581 B.n541 VSUBS 0.007467f
C582 B.n542 VSUBS 0.007467f
C583 B.n543 VSUBS 0.007467f
C584 B.n544 VSUBS 0.007467f
C585 B.n545 VSUBS 0.007467f
C586 B.n546 VSUBS 0.007467f
C587 B.n547 VSUBS 0.007467f
C588 B.n548 VSUBS 0.007467f
C589 B.n549 VSUBS 0.007467f
C590 B.n550 VSUBS 0.007467f
C591 B.n551 VSUBS 0.007467f
C592 B.n552 VSUBS 0.007467f
C593 B.n553 VSUBS 0.007467f
C594 B.n554 VSUBS 0.007467f
C595 B.n555 VSUBS 0.007467f
C596 B.n556 VSUBS 0.007467f
C597 B.n557 VSUBS 0.007467f
C598 B.n558 VSUBS 0.007467f
C599 B.n559 VSUBS 0.007467f
C600 B.n560 VSUBS 0.007467f
C601 B.n561 VSUBS 0.007467f
C602 B.n562 VSUBS 0.007467f
C603 B.n563 VSUBS 0.007467f
C604 B.n564 VSUBS 0.007467f
C605 B.n565 VSUBS 0.007467f
C606 B.n566 VSUBS 0.007467f
C607 B.n567 VSUBS 0.007467f
C608 B.n568 VSUBS 0.007467f
C609 B.n569 VSUBS 0.007467f
C610 B.n570 VSUBS 0.007467f
C611 B.n571 VSUBS 0.007467f
C612 B.n572 VSUBS 0.007467f
C613 B.n573 VSUBS 0.007467f
C614 B.n574 VSUBS 0.007467f
C615 B.n575 VSUBS 0.007467f
C616 B.n576 VSUBS 0.007467f
C617 B.n577 VSUBS 0.007467f
C618 B.n578 VSUBS 0.007467f
C619 B.n579 VSUBS 0.007467f
C620 B.n580 VSUBS 0.007467f
C621 B.n581 VSUBS 0.007467f
C622 B.n582 VSUBS 0.007467f
C623 B.n583 VSUBS 0.007467f
C624 B.n584 VSUBS 0.007467f
C625 B.n585 VSUBS 0.007467f
C626 B.n586 VSUBS 0.007467f
C627 B.n587 VSUBS 0.007467f
C628 B.n588 VSUBS 0.007467f
C629 B.n589 VSUBS 0.007467f
C630 B.n590 VSUBS 0.007467f
C631 B.n591 VSUBS 0.007467f
C632 B.n592 VSUBS 0.007467f
C633 B.n593 VSUBS 0.007467f
C634 B.n594 VSUBS 0.007467f
C635 B.n595 VSUBS 0.007467f
C636 B.n596 VSUBS 0.007467f
C637 B.n597 VSUBS 0.007467f
C638 B.n598 VSUBS 0.007467f
C639 B.n599 VSUBS 0.007467f
C640 B.n600 VSUBS 0.007467f
C641 B.n601 VSUBS 0.007467f
C642 B.n602 VSUBS 0.007467f
C643 B.n603 VSUBS 0.007467f
C644 B.n604 VSUBS 0.007467f
C645 B.n605 VSUBS 0.007467f
C646 B.n606 VSUBS 0.007467f
C647 B.n607 VSUBS 0.007467f
C648 B.n608 VSUBS 0.007467f
C649 B.n609 VSUBS 0.007467f
C650 B.n610 VSUBS 0.007467f
C651 B.n611 VSUBS 0.007467f
C652 B.n612 VSUBS 0.007467f
C653 B.n613 VSUBS 0.007467f
C654 B.n614 VSUBS 0.007467f
C655 B.n615 VSUBS 0.007467f
C656 B.n616 VSUBS 0.018202f
C657 B.n617 VSUBS 0.018202f
C658 B.n618 VSUBS 0.016715f
C659 B.n619 VSUBS 0.007467f
C660 B.n620 VSUBS 0.007467f
C661 B.n621 VSUBS 0.007467f
C662 B.n622 VSUBS 0.007467f
C663 B.n623 VSUBS 0.007467f
C664 B.n624 VSUBS 0.007467f
C665 B.n625 VSUBS 0.007467f
C666 B.n626 VSUBS 0.007467f
C667 B.n627 VSUBS 0.007467f
C668 B.n628 VSUBS 0.007467f
C669 B.n629 VSUBS 0.007467f
C670 B.n630 VSUBS 0.007467f
C671 B.n631 VSUBS 0.007467f
C672 B.n632 VSUBS 0.007467f
C673 B.n633 VSUBS 0.007467f
C674 B.n634 VSUBS 0.007467f
C675 B.n635 VSUBS 0.007467f
C676 B.n636 VSUBS 0.007467f
C677 B.n637 VSUBS 0.007467f
C678 B.n638 VSUBS 0.007467f
C679 B.n639 VSUBS 0.007467f
C680 B.n640 VSUBS 0.007467f
C681 B.n641 VSUBS 0.007467f
C682 B.n642 VSUBS 0.007467f
C683 B.n643 VSUBS 0.007467f
C684 B.n644 VSUBS 0.007467f
C685 B.n645 VSUBS 0.007467f
C686 B.n646 VSUBS 0.007467f
C687 B.n647 VSUBS 0.007467f
C688 B.n648 VSUBS 0.007467f
C689 B.n649 VSUBS 0.007467f
C690 B.n650 VSUBS 0.007467f
C691 B.n651 VSUBS 0.007467f
C692 B.n652 VSUBS 0.007467f
C693 B.n653 VSUBS 0.007467f
C694 B.n654 VSUBS 0.007467f
C695 B.n655 VSUBS 0.007467f
C696 B.n656 VSUBS 0.007467f
C697 B.n657 VSUBS 0.007467f
C698 B.n658 VSUBS 0.007467f
C699 B.n659 VSUBS 0.007467f
C700 B.n660 VSUBS 0.007467f
C701 B.n661 VSUBS 0.007467f
C702 B.n662 VSUBS 0.007467f
C703 B.n663 VSUBS 0.007467f
C704 B.n664 VSUBS 0.007467f
C705 B.n665 VSUBS 0.007467f
C706 B.n666 VSUBS 0.007467f
C707 B.n667 VSUBS 0.007467f
C708 B.n668 VSUBS 0.007467f
C709 B.n669 VSUBS 0.007467f
C710 B.n670 VSUBS 0.007467f
C711 B.n671 VSUBS 0.007467f
C712 B.n672 VSUBS 0.007467f
C713 B.n673 VSUBS 0.007467f
C714 B.n674 VSUBS 0.007467f
C715 B.n675 VSUBS 0.007467f
C716 B.n676 VSUBS 0.007467f
C717 B.n677 VSUBS 0.007467f
C718 B.n678 VSUBS 0.007467f
C719 B.n679 VSUBS 0.007467f
C720 B.n680 VSUBS 0.007467f
C721 B.n681 VSUBS 0.007467f
C722 B.n682 VSUBS 0.007467f
C723 B.n683 VSUBS 0.007467f
C724 B.n684 VSUBS 0.007467f
C725 B.n685 VSUBS 0.007467f
C726 B.n686 VSUBS 0.007467f
C727 B.n687 VSUBS 0.007467f
C728 B.n688 VSUBS 0.007467f
C729 B.n689 VSUBS 0.007467f
C730 B.n690 VSUBS 0.007467f
C731 B.n691 VSUBS 0.007467f
C732 B.n692 VSUBS 0.007467f
C733 B.n693 VSUBS 0.007467f
C734 B.n694 VSUBS 0.007467f
C735 B.n695 VSUBS 0.007467f
C736 B.n696 VSUBS 0.007467f
C737 B.n697 VSUBS 0.007467f
C738 B.n698 VSUBS 0.007467f
C739 B.n699 VSUBS 0.007467f
C740 B.n700 VSUBS 0.007467f
C741 B.n701 VSUBS 0.007467f
C742 B.n702 VSUBS 0.007467f
C743 B.n703 VSUBS 0.007467f
C744 B.n704 VSUBS 0.007467f
C745 B.n705 VSUBS 0.007467f
C746 B.n706 VSUBS 0.007467f
C747 B.n707 VSUBS 0.007467f
C748 B.n708 VSUBS 0.007467f
C749 B.n709 VSUBS 0.007467f
C750 B.n710 VSUBS 0.007467f
C751 B.n711 VSUBS 0.007467f
C752 B.n712 VSUBS 0.007467f
C753 B.n713 VSUBS 0.007467f
C754 B.n714 VSUBS 0.007467f
C755 B.n715 VSUBS 0.007467f
C756 B.n716 VSUBS 0.007467f
C757 B.n717 VSUBS 0.007467f
C758 B.n718 VSUBS 0.007467f
C759 B.n719 VSUBS 0.007467f
C760 B.n720 VSUBS 0.007467f
C761 B.n721 VSUBS 0.007467f
C762 B.n722 VSUBS 0.007467f
C763 B.n723 VSUBS 0.007467f
C764 B.n724 VSUBS 0.007467f
C765 B.n725 VSUBS 0.007467f
C766 B.n726 VSUBS 0.007467f
C767 B.n727 VSUBS 0.007467f
C768 B.n728 VSUBS 0.007467f
C769 B.n729 VSUBS 0.007467f
C770 B.n730 VSUBS 0.007467f
C771 B.n731 VSUBS 0.007467f
C772 B.n732 VSUBS 0.007467f
C773 B.n733 VSUBS 0.007467f
C774 B.n734 VSUBS 0.007467f
C775 B.n735 VSUBS 0.007467f
C776 B.n736 VSUBS 0.007467f
C777 B.n737 VSUBS 0.007467f
C778 B.n738 VSUBS 0.007467f
C779 B.n739 VSUBS 0.007467f
C780 B.n740 VSUBS 0.007467f
C781 B.n741 VSUBS 0.007467f
C782 B.n742 VSUBS 0.007467f
C783 B.n743 VSUBS 0.007467f
C784 B.n744 VSUBS 0.007467f
C785 B.n745 VSUBS 0.007467f
C786 B.n746 VSUBS 0.007467f
C787 B.n747 VSUBS 0.007467f
C788 B.n748 VSUBS 0.007467f
C789 B.n749 VSUBS 0.007467f
C790 B.n750 VSUBS 0.007467f
C791 B.n751 VSUBS 0.007467f
C792 B.n752 VSUBS 0.007467f
C793 B.n753 VSUBS 0.007467f
C794 B.n754 VSUBS 0.007467f
C795 B.n755 VSUBS 0.007467f
C796 B.n756 VSUBS 0.007467f
C797 B.n757 VSUBS 0.007467f
C798 B.n758 VSUBS 0.007467f
C799 B.n759 VSUBS 0.007467f
C800 B.n760 VSUBS 0.007467f
C801 B.n761 VSUBS 0.007467f
C802 B.n762 VSUBS 0.007467f
C803 B.n763 VSUBS 0.007467f
C804 B.n764 VSUBS 0.007467f
C805 B.n765 VSUBS 0.007467f
C806 B.n766 VSUBS 0.007467f
C807 B.n767 VSUBS 0.007467f
C808 B.n768 VSUBS 0.007467f
C809 B.n769 VSUBS 0.007467f
C810 B.n770 VSUBS 0.007467f
C811 B.n771 VSUBS 0.007467f
C812 B.n772 VSUBS 0.007467f
C813 B.n773 VSUBS 0.007467f
C814 B.n774 VSUBS 0.007467f
C815 B.n775 VSUBS 0.007467f
C816 B.n776 VSUBS 0.007467f
C817 B.n777 VSUBS 0.007467f
C818 B.n778 VSUBS 0.007467f
C819 B.n779 VSUBS 0.007467f
C820 B.n780 VSUBS 0.007467f
C821 B.n781 VSUBS 0.007467f
C822 B.n782 VSUBS 0.007467f
C823 B.n783 VSUBS 0.007467f
C824 B.n784 VSUBS 0.007467f
C825 B.n785 VSUBS 0.007467f
C826 B.n786 VSUBS 0.007467f
C827 B.n787 VSUBS 0.007467f
C828 B.n788 VSUBS 0.007467f
C829 B.n789 VSUBS 0.007467f
C830 B.n790 VSUBS 0.007467f
C831 B.n791 VSUBS 0.007467f
C832 B.n792 VSUBS 0.007467f
C833 B.n793 VSUBS 0.007467f
C834 B.n794 VSUBS 0.007467f
C835 B.n795 VSUBS 0.007467f
C836 B.n796 VSUBS 0.007467f
C837 B.n797 VSUBS 0.007467f
C838 B.n798 VSUBS 0.007467f
C839 B.n799 VSUBS 0.007467f
C840 B.n800 VSUBS 0.007467f
C841 B.n801 VSUBS 0.007467f
C842 B.n802 VSUBS 0.007467f
C843 B.n803 VSUBS 0.007467f
C844 B.n804 VSUBS 0.007467f
C845 B.n805 VSUBS 0.007467f
C846 B.n806 VSUBS 0.007467f
C847 B.n807 VSUBS 0.007467f
C848 B.n808 VSUBS 0.007467f
C849 B.n809 VSUBS 0.007467f
C850 B.n810 VSUBS 0.007467f
C851 B.n811 VSUBS 0.007467f
C852 B.n812 VSUBS 0.007467f
C853 B.n813 VSUBS 0.007467f
C854 B.n814 VSUBS 0.007467f
C855 B.n815 VSUBS 0.007467f
C856 B.n816 VSUBS 0.007467f
C857 B.n817 VSUBS 0.007467f
C858 B.n818 VSUBS 0.007467f
C859 B.n819 VSUBS 0.007467f
C860 B.n820 VSUBS 0.007467f
C861 B.n821 VSUBS 0.007467f
C862 B.n822 VSUBS 0.007467f
C863 B.n823 VSUBS 0.007467f
C864 B.n824 VSUBS 0.007467f
C865 B.n825 VSUBS 0.007467f
C866 B.n826 VSUBS 0.007467f
C867 B.n827 VSUBS 0.007467f
C868 B.n828 VSUBS 0.007467f
C869 B.n829 VSUBS 0.007467f
C870 B.n830 VSUBS 0.007467f
C871 B.n831 VSUBS 0.007467f
C872 B.n832 VSUBS 0.007467f
C873 B.n833 VSUBS 0.007467f
C874 B.n834 VSUBS 0.007467f
C875 B.n835 VSUBS 0.007467f
C876 B.n836 VSUBS 0.007467f
C877 B.n837 VSUBS 0.007467f
C878 B.n838 VSUBS 0.007467f
C879 B.n839 VSUBS 0.007467f
C880 B.n840 VSUBS 0.007467f
C881 B.n841 VSUBS 0.007467f
C882 B.n842 VSUBS 0.007467f
C883 B.n843 VSUBS 0.007467f
C884 B.n844 VSUBS 0.007467f
C885 B.n845 VSUBS 0.007467f
C886 B.n846 VSUBS 0.007467f
C887 B.n847 VSUBS 0.007467f
C888 B.n848 VSUBS 0.007467f
C889 B.n849 VSUBS 0.007467f
C890 B.n850 VSUBS 0.007467f
C891 B.n851 VSUBS 0.007467f
C892 B.n852 VSUBS 0.007467f
C893 B.n853 VSUBS 0.007467f
C894 B.n854 VSUBS 0.007467f
C895 B.n855 VSUBS 0.016715f
C896 B.n856 VSUBS 0.018202f
C897 B.n857 VSUBS 0.017319f
C898 B.n858 VSUBS 0.007467f
C899 B.n859 VSUBS 0.007467f
C900 B.n860 VSUBS 0.007467f
C901 B.n861 VSUBS 0.007467f
C902 B.n862 VSUBS 0.007467f
C903 B.n863 VSUBS 0.007467f
C904 B.n864 VSUBS 0.007467f
C905 B.n865 VSUBS 0.007467f
C906 B.n866 VSUBS 0.007467f
C907 B.n867 VSUBS 0.007467f
C908 B.n868 VSUBS 0.007467f
C909 B.n869 VSUBS 0.007467f
C910 B.n870 VSUBS 0.007467f
C911 B.n871 VSUBS 0.007467f
C912 B.n872 VSUBS 0.007467f
C913 B.n873 VSUBS 0.007467f
C914 B.n874 VSUBS 0.007467f
C915 B.n875 VSUBS 0.007467f
C916 B.n876 VSUBS 0.007467f
C917 B.n877 VSUBS 0.007467f
C918 B.n878 VSUBS 0.007467f
C919 B.n879 VSUBS 0.007467f
C920 B.n880 VSUBS 0.007467f
C921 B.n881 VSUBS 0.007467f
C922 B.n882 VSUBS 0.007467f
C923 B.n883 VSUBS 0.007467f
C924 B.n884 VSUBS 0.007467f
C925 B.n885 VSUBS 0.007467f
C926 B.n886 VSUBS 0.007467f
C927 B.n887 VSUBS 0.007467f
C928 B.n888 VSUBS 0.007467f
C929 B.n889 VSUBS 0.007467f
C930 B.n890 VSUBS 0.007467f
C931 B.n891 VSUBS 0.007467f
C932 B.n892 VSUBS 0.007467f
C933 B.n893 VSUBS 0.007467f
C934 B.n894 VSUBS 0.007467f
C935 B.n895 VSUBS 0.007467f
C936 B.n896 VSUBS 0.007467f
C937 B.n897 VSUBS 0.007467f
C938 B.n898 VSUBS 0.007467f
C939 B.n899 VSUBS 0.007467f
C940 B.n900 VSUBS 0.007467f
C941 B.n901 VSUBS 0.007467f
C942 B.n902 VSUBS 0.007467f
C943 B.n903 VSUBS 0.007467f
C944 B.n904 VSUBS 0.007467f
C945 B.n905 VSUBS 0.007467f
C946 B.n906 VSUBS 0.007467f
C947 B.n907 VSUBS 0.007467f
C948 B.n908 VSUBS 0.007467f
C949 B.n909 VSUBS 0.007467f
C950 B.n910 VSUBS 0.007467f
C951 B.n911 VSUBS 0.007467f
C952 B.n912 VSUBS 0.007467f
C953 B.n913 VSUBS 0.007467f
C954 B.n914 VSUBS 0.007467f
C955 B.n915 VSUBS 0.007467f
C956 B.n916 VSUBS 0.007467f
C957 B.n917 VSUBS 0.007467f
C958 B.n918 VSUBS 0.007467f
C959 B.n919 VSUBS 0.007467f
C960 B.n920 VSUBS 0.007467f
C961 B.n921 VSUBS 0.007467f
C962 B.n922 VSUBS 0.007467f
C963 B.n923 VSUBS 0.007467f
C964 B.n924 VSUBS 0.007467f
C965 B.n925 VSUBS 0.007467f
C966 B.n926 VSUBS 0.007467f
C967 B.n927 VSUBS 0.007467f
C968 B.n928 VSUBS 0.007467f
C969 B.n929 VSUBS 0.007467f
C970 B.n930 VSUBS 0.007467f
C971 B.n931 VSUBS 0.007467f
C972 B.n932 VSUBS 0.007467f
C973 B.n933 VSUBS 0.007467f
C974 B.n934 VSUBS 0.007467f
C975 B.n935 VSUBS 0.007467f
C976 B.n936 VSUBS 0.007467f
C977 B.n937 VSUBS 0.007467f
C978 B.n938 VSUBS 0.007467f
C979 B.n939 VSUBS 0.007467f
C980 B.n940 VSUBS 0.007467f
C981 B.n941 VSUBS 0.007467f
C982 B.n942 VSUBS 0.007467f
C983 B.n943 VSUBS 0.007467f
C984 B.n944 VSUBS 0.007467f
C985 B.n945 VSUBS 0.007467f
C986 B.n946 VSUBS 0.007467f
C987 B.n947 VSUBS 0.007027f
C988 B.n948 VSUBS 0.017299f
C989 B.n949 VSUBS 0.004172f
C990 B.n950 VSUBS 0.007467f
C991 B.n951 VSUBS 0.007467f
C992 B.n952 VSUBS 0.007467f
C993 B.n953 VSUBS 0.007467f
C994 B.n954 VSUBS 0.007467f
C995 B.n955 VSUBS 0.007467f
C996 B.n956 VSUBS 0.007467f
C997 B.n957 VSUBS 0.007467f
C998 B.n958 VSUBS 0.007467f
C999 B.n959 VSUBS 0.007467f
C1000 B.n960 VSUBS 0.007467f
C1001 B.n961 VSUBS 0.007467f
C1002 B.n962 VSUBS 0.004172f
C1003 B.n963 VSUBS 0.007467f
C1004 B.n964 VSUBS 0.007467f
C1005 B.n965 VSUBS 0.007027f
C1006 B.n966 VSUBS 0.007467f
C1007 B.n967 VSUBS 0.007467f
C1008 B.n968 VSUBS 0.007467f
C1009 B.n969 VSUBS 0.007467f
C1010 B.n970 VSUBS 0.007467f
C1011 B.n971 VSUBS 0.007467f
C1012 B.n972 VSUBS 0.007467f
C1013 B.n973 VSUBS 0.007467f
C1014 B.n974 VSUBS 0.007467f
C1015 B.n975 VSUBS 0.007467f
C1016 B.n976 VSUBS 0.007467f
C1017 B.n977 VSUBS 0.007467f
C1018 B.n978 VSUBS 0.007467f
C1019 B.n979 VSUBS 0.007467f
C1020 B.n980 VSUBS 0.007467f
C1021 B.n981 VSUBS 0.007467f
C1022 B.n982 VSUBS 0.007467f
C1023 B.n983 VSUBS 0.007467f
C1024 B.n984 VSUBS 0.007467f
C1025 B.n985 VSUBS 0.007467f
C1026 B.n986 VSUBS 0.007467f
C1027 B.n987 VSUBS 0.007467f
C1028 B.n988 VSUBS 0.007467f
C1029 B.n989 VSUBS 0.007467f
C1030 B.n990 VSUBS 0.007467f
C1031 B.n991 VSUBS 0.007467f
C1032 B.n992 VSUBS 0.007467f
C1033 B.n993 VSUBS 0.007467f
C1034 B.n994 VSUBS 0.007467f
C1035 B.n995 VSUBS 0.007467f
C1036 B.n996 VSUBS 0.007467f
C1037 B.n997 VSUBS 0.007467f
C1038 B.n998 VSUBS 0.007467f
C1039 B.n999 VSUBS 0.007467f
C1040 B.n1000 VSUBS 0.007467f
C1041 B.n1001 VSUBS 0.007467f
C1042 B.n1002 VSUBS 0.007467f
C1043 B.n1003 VSUBS 0.007467f
C1044 B.n1004 VSUBS 0.007467f
C1045 B.n1005 VSUBS 0.007467f
C1046 B.n1006 VSUBS 0.007467f
C1047 B.n1007 VSUBS 0.007467f
C1048 B.n1008 VSUBS 0.007467f
C1049 B.n1009 VSUBS 0.007467f
C1050 B.n1010 VSUBS 0.007467f
C1051 B.n1011 VSUBS 0.007467f
C1052 B.n1012 VSUBS 0.007467f
C1053 B.n1013 VSUBS 0.007467f
C1054 B.n1014 VSUBS 0.007467f
C1055 B.n1015 VSUBS 0.007467f
C1056 B.n1016 VSUBS 0.007467f
C1057 B.n1017 VSUBS 0.007467f
C1058 B.n1018 VSUBS 0.007467f
C1059 B.n1019 VSUBS 0.007467f
C1060 B.n1020 VSUBS 0.007467f
C1061 B.n1021 VSUBS 0.007467f
C1062 B.n1022 VSUBS 0.007467f
C1063 B.n1023 VSUBS 0.007467f
C1064 B.n1024 VSUBS 0.007467f
C1065 B.n1025 VSUBS 0.007467f
C1066 B.n1026 VSUBS 0.007467f
C1067 B.n1027 VSUBS 0.007467f
C1068 B.n1028 VSUBS 0.007467f
C1069 B.n1029 VSUBS 0.007467f
C1070 B.n1030 VSUBS 0.007467f
C1071 B.n1031 VSUBS 0.007467f
C1072 B.n1032 VSUBS 0.007467f
C1073 B.n1033 VSUBS 0.007467f
C1074 B.n1034 VSUBS 0.007467f
C1075 B.n1035 VSUBS 0.007467f
C1076 B.n1036 VSUBS 0.007467f
C1077 B.n1037 VSUBS 0.007467f
C1078 B.n1038 VSUBS 0.007467f
C1079 B.n1039 VSUBS 0.007467f
C1080 B.n1040 VSUBS 0.007467f
C1081 B.n1041 VSUBS 0.007467f
C1082 B.n1042 VSUBS 0.007467f
C1083 B.n1043 VSUBS 0.007467f
C1084 B.n1044 VSUBS 0.007467f
C1085 B.n1045 VSUBS 0.007467f
C1086 B.n1046 VSUBS 0.007467f
C1087 B.n1047 VSUBS 0.007467f
C1088 B.n1048 VSUBS 0.007467f
C1089 B.n1049 VSUBS 0.007467f
C1090 B.n1050 VSUBS 0.007467f
C1091 B.n1051 VSUBS 0.007467f
C1092 B.n1052 VSUBS 0.007467f
C1093 B.n1053 VSUBS 0.007467f
C1094 B.n1054 VSUBS 0.018202f
C1095 B.n1055 VSUBS 0.018202f
C1096 B.n1056 VSUBS 0.016715f
C1097 B.n1057 VSUBS 0.007467f
C1098 B.n1058 VSUBS 0.007467f
C1099 B.n1059 VSUBS 0.007467f
C1100 B.n1060 VSUBS 0.007467f
C1101 B.n1061 VSUBS 0.007467f
C1102 B.n1062 VSUBS 0.007467f
C1103 B.n1063 VSUBS 0.007467f
C1104 B.n1064 VSUBS 0.007467f
C1105 B.n1065 VSUBS 0.007467f
C1106 B.n1066 VSUBS 0.007467f
C1107 B.n1067 VSUBS 0.007467f
C1108 B.n1068 VSUBS 0.007467f
C1109 B.n1069 VSUBS 0.007467f
C1110 B.n1070 VSUBS 0.007467f
C1111 B.n1071 VSUBS 0.007467f
C1112 B.n1072 VSUBS 0.007467f
C1113 B.n1073 VSUBS 0.007467f
C1114 B.n1074 VSUBS 0.007467f
C1115 B.n1075 VSUBS 0.007467f
C1116 B.n1076 VSUBS 0.007467f
C1117 B.n1077 VSUBS 0.007467f
C1118 B.n1078 VSUBS 0.007467f
C1119 B.n1079 VSUBS 0.007467f
C1120 B.n1080 VSUBS 0.007467f
C1121 B.n1081 VSUBS 0.007467f
C1122 B.n1082 VSUBS 0.007467f
C1123 B.n1083 VSUBS 0.007467f
C1124 B.n1084 VSUBS 0.007467f
C1125 B.n1085 VSUBS 0.007467f
C1126 B.n1086 VSUBS 0.007467f
C1127 B.n1087 VSUBS 0.007467f
C1128 B.n1088 VSUBS 0.007467f
C1129 B.n1089 VSUBS 0.007467f
C1130 B.n1090 VSUBS 0.007467f
C1131 B.n1091 VSUBS 0.007467f
C1132 B.n1092 VSUBS 0.007467f
C1133 B.n1093 VSUBS 0.007467f
C1134 B.n1094 VSUBS 0.007467f
C1135 B.n1095 VSUBS 0.007467f
C1136 B.n1096 VSUBS 0.007467f
C1137 B.n1097 VSUBS 0.007467f
C1138 B.n1098 VSUBS 0.007467f
C1139 B.n1099 VSUBS 0.007467f
C1140 B.n1100 VSUBS 0.007467f
C1141 B.n1101 VSUBS 0.007467f
C1142 B.n1102 VSUBS 0.007467f
C1143 B.n1103 VSUBS 0.007467f
C1144 B.n1104 VSUBS 0.007467f
C1145 B.n1105 VSUBS 0.007467f
C1146 B.n1106 VSUBS 0.007467f
C1147 B.n1107 VSUBS 0.007467f
C1148 B.n1108 VSUBS 0.007467f
C1149 B.n1109 VSUBS 0.007467f
C1150 B.n1110 VSUBS 0.007467f
C1151 B.n1111 VSUBS 0.007467f
C1152 B.n1112 VSUBS 0.007467f
C1153 B.n1113 VSUBS 0.007467f
C1154 B.n1114 VSUBS 0.007467f
C1155 B.n1115 VSUBS 0.007467f
C1156 B.n1116 VSUBS 0.007467f
C1157 B.n1117 VSUBS 0.007467f
C1158 B.n1118 VSUBS 0.007467f
C1159 B.n1119 VSUBS 0.007467f
C1160 B.n1120 VSUBS 0.007467f
C1161 B.n1121 VSUBS 0.007467f
C1162 B.n1122 VSUBS 0.007467f
C1163 B.n1123 VSUBS 0.007467f
C1164 B.n1124 VSUBS 0.007467f
C1165 B.n1125 VSUBS 0.007467f
C1166 B.n1126 VSUBS 0.007467f
C1167 B.n1127 VSUBS 0.007467f
C1168 B.n1128 VSUBS 0.007467f
C1169 B.n1129 VSUBS 0.007467f
C1170 B.n1130 VSUBS 0.007467f
C1171 B.n1131 VSUBS 0.007467f
C1172 B.n1132 VSUBS 0.007467f
C1173 B.n1133 VSUBS 0.007467f
C1174 B.n1134 VSUBS 0.007467f
C1175 B.n1135 VSUBS 0.007467f
C1176 B.n1136 VSUBS 0.007467f
C1177 B.n1137 VSUBS 0.007467f
C1178 B.n1138 VSUBS 0.007467f
C1179 B.n1139 VSUBS 0.007467f
C1180 B.n1140 VSUBS 0.007467f
C1181 B.n1141 VSUBS 0.007467f
C1182 B.n1142 VSUBS 0.007467f
C1183 B.n1143 VSUBS 0.007467f
C1184 B.n1144 VSUBS 0.007467f
C1185 B.n1145 VSUBS 0.007467f
C1186 B.n1146 VSUBS 0.007467f
C1187 B.n1147 VSUBS 0.007467f
C1188 B.n1148 VSUBS 0.007467f
C1189 B.n1149 VSUBS 0.007467f
C1190 B.n1150 VSUBS 0.007467f
C1191 B.n1151 VSUBS 0.007467f
C1192 B.n1152 VSUBS 0.007467f
C1193 B.n1153 VSUBS 0.007467f
C1194 B.n1154 VSUBS 0.007467f
C1195 B.n1155 VSUBS 0.007467f
C1196 B.n1156 VSUBS 0.007467f
C1197 B.n1157 VSUBS 0.007467f
C1198 B.n1158 VSUBS 0.007467f
C1199 B.n1159 VSUBS 0.007467f
C1200 B.n1160 VSUBS 0.007467f
C1201 B.n1161 VSUBS 0.007467f
C1202 B.n1162 VSUBS 0.007467f
C1203 B.n1163 VSUBS 0.007467f
C1204 B.n1164 VSUBS 0.007467f
C1205 B.n1165 VSUBS 0.007467f
C1206 B.n1166 VSUBS 0.007467f
C1207 B.n1167 VSUBS 0.007467f
C1208 B.n1168 VSUBS 0.007467f
C1209 B.n1169 VSUBS 0.007467f
C1210 B.n1170 VSUBS 0.007467f
C1211 B.n1171 VSUBS 0.007467f
C1212 B.n1172 VSUBS 0.007467f
C1213 B.n1173 VSUBS 0.007467f
C1214 B.n1174 VSUBS 0.007467f
C1215 B.n1175 VSUBS 0.016907f
C1216 VDD1.t8 VSUBS 4.63734f
C1217 VDD1.t1 VSUBS 0.424509f
C1218 VDD1.t9 VSUBS 0.424509f
C1219 VDD1.n0 VSUBS 3.53814f
C1220 VDD1.n1 VSUBS 1.95277f
C1221 VDD1.t6 VSUBS 4.63732f
C1222 VDD1.t0 VSUBS 0.424509f
C1223 VDD1.t2 VSUBS 0.424509f
C1224 VDD1.n2 VSUBS 3.53814f
C1225 VDD1.n3 VSUBS 1.94305f
C1226 VDD1.t3 VSUBS 0.424509f
C1227 VDD1.t7 VSUBS 0.424509f
C1228 VDD1.n4 VSUBS 3.57942f
C1229 VDD1.n5 VSUBS 5.01218f
C1230 VDD1.t4 VSUBS 0.424509f
C1231 VDD1.t5 VSUBS 0.424509f
C1232 VDD1.n6 VSUBS 3.53813f
C1233 VDD1.n7 VSUBS 5.10394f
C1234 VP.t2 VSUBS 4.1413f
C1235 VP.n0 VSUBS 1.50589f
C1236 VP.n1 VSUBS 0.021876f
C1237 VP.n2 VSUBS 0.042236f
C1238 VP.n3 VSUBS 0.021876f
C1239 VP.n4 VSUBS 0.039564f
C1240 VP.n5 VSUBS 0.021876f
C1241 VP.n6 VSUBS 0.043121f
C1242 VP.n7 VSUBS 0.021876f
C1243 VP.n8 VSUBS 0.040772f
C1244 VP.n9 VSUBS 0.021876f
C1245 VP.t7 VSUBS 4.1413f
C1246 VP.n10 VSUBS 0.043777f
C1247 VP.n11 VSUBS 0.021876f
C1248 VP.n12 VSUBS 0.040772f
C1249 VP.n13 VSUBS 0.021876f
C1250 VP.t9 VSUBS 4.1413f
C1251 VP.n14 VSUBS 0.044149f
C1252 VP.n15 VSUBS 0.021876f
C1253 VP.n16 VSUBS 0.040772f
C1254 VP.t4 VSUBS 4.1413f
C1255 VP.n17 VSUBS 1.50589f
C1256 VP.n18 VSUBS 0.021876f
C1257 VP.n19 VSUBS 0.042236f
C1258 VP.n20 VSUBS 0.021876f
C1259 VP.n21 VSUBS 0.039564f
C1260 VP.n22 VSUBS 0.021876f
C1261 VP.n23 VSUBS 0.043121f
C1262 VP.n24 VSUBS 0.021876f
C1263 VP.n25 VSUBS 0.040772f
C1264 VP.n26 VSUBS 0.021876f
C1265 VP.t0 VSUBS 4.1413f
C1266 VP.n27 VSUBS 0.043777f
C1267 VP.n28 VSUBS 0.021876f
C1268 VP.n29 VSUBS 0.040772f
C1269 VP.t1 VSUBS 4.47307f
C1270 VP.n30 VSUBS 1.43554f
C1271 VP.t8 VSUBS 4.1413f
C1272 VP.n31 VSUBS 1.49541f
C1273 VP.n32 VSUBS 0.02185f
C1274 VP.n33 VSUBS 0.278f
C1275 VP.n34 VSUBS 0.021876f
C1276 VP.n35 VSUBS 0.021876f
C1277 VP.n36 VSUBS 0.040772f
C1278 VP.n37 VSUBS 0.043121f
C1279 VP.n38 VSUBS 0.017749f
C1280 VP.n39 VSUBS 0.021876f
C1281 VP.n40 VSUBS 0.021876f
C1282 VP.n41 VSUBS 0.021876f
C1283 VP.n42 VSUBS 0.040772f
C1284 VP.n43 VSUBS 0.040772f
C1285 VP.n44 VSUBS 1.44641f
C1286 VP.n45 VSUBS 0.021876f
C1287 VP.n46 VSUBS 0.021876f
C1288 VP.n47 VSUBS 0.021876f
C1289 VP.n48 VSUBS 0.040772f
C1290 VP.n49 VSUBS 0.043777f
C1291 VP.n50 VSUBS 0.017749f
C1292 VP.n51 VSUBS 0.021876f
C1293 VP.n52 VSUBS 0.021876f
C1294 VP.n53 VSUBS 0.021876f
C1295 VP.n54 VSUBS 0.040772f
C1296 VP.n55 VSUBS 0.040772f
C1297 VP.t5 VSUBS 4.1413f
C1298 VP.n56 VSUBS 1.42577f
C1299 VP.n57 VSUBS 0.02185f
C1300 VP.n58 VSUBS 0.021876f
C1301 VP.n59 VSUBS 0.021876f
C1302 VP.n60 VSUBS 0.021876f
C1303 VP.n61 VSUBS 0.040772f
C1304 VP.n62 VSUBS 0.044149f
C1305 VP.n63 VSUBS 0.018261f
C1306 VP.n64 VSUBS 0.021876f
C1307 VP.n65 VSUBS 0.021876f
C1308 VP.n66 VSUBS 0.021876f
C1309 VP.n67 VSUBS 0.040772f
C1310 VP.n68 VSUBS 0.040772f
C1311 VP.n69 VSUBS 0.023058f
C1312 VP.n70 VSUBS 0.035308f
C1313 VP.n71 VSUBS 1.76138f
C1314 VP.n72 VSUBS 1.77364f
C1315 VP.t3 VSUBS 4.1413f
C1316 VP.n73 VSUBS 1.50589f
C1317 VP.n74 VSUBS 0.023058f
C1318 VP.n75 VSUBS 0.035308f
C1319 VP.n76 VSUBS 0.021876f
C1320 VP.n77 VSUBS 0.021876f
C1321 VP.n78 VSUBS 0.040772f
C1322 VP.n79 VSUBS 0.042236f
C1323 VP.n80 VSUBS 0.018261f
C1324 VP.n81 VSUBS 0.021876f
C1325 VP.n82 VSUBS 0.021876f
C1326 VP.n83 VSUBS 0.021876f
C1327 VP.n84 VSUBS 0.040772f
C1328 VP.n85 VSUBS 0.039564f
C1329 VP.n86 VSUBS 1.42577f
C1330 VP.n87 VSUBS 0.02185f
C1331 VP.n88 VSUBS 0.021876f
C1332 VP.n89 VSUBS 0.021876f
C1333 VP.n90 VSUBS 0.021876f
C1334 VP.n91 VSUBS 0.040772f
C1335 VP.n92 VSUBS 0.043121f
C1336 VP.n93 VSUBS 0.017749f
C1337 VP.n94 VSUBS 0.021876f
C1338 VP.n95 VSUBS 0.021876f
C1339 VP.n96 VSUBS 0.021876f
C1340 VP.n97 VSUBS 0.040772f
C1341 VP.n98 VSUBS 0.040772f
C1342 VP.n99 VSUBS 1.44641f
C1343 VP.n100 VSUBS 0.021876f
C1344 VP.n101 VSUBS 0.021876f
C1345 VP.n102 VSUBS 0.021876f
C1346 VP.n103 VSUBS 0.040772f
C1347 VP.n104 VSUBS 0.043777f
C1348 VP.n105 VSUBS 0.017749f
C1349 VP.n106 VSUBS 0.021876f
C1350 VP.n107 VSUBS 0.021876f
C1351 VP.n108 VSUBS 0.021876f
C1352 VP.n109 VSUBS 0.040772f
C1353 VP.n110 VSUBS 0.040772f
C1354 VP.t6 VSUBS 4.1413f
C1355 VP.n111 VSUBS 1.42577f
C1356 VP.n112 VSUBS 0.02185f
C1357 VP.n113 VSUBS 0.021876f
C1358 VP.n114 VSUBS 0.021876f
C1359 VP.n115 VSUBS 0.021876f
C1360 VP.n116 VSUBS 0.040772f
C1361 VP.n117 VSUBS 0.044149f
C1362 VP.n118 VSUBS 0.018261f
C1363 VP.n119 VSUBS 0.021876f
C1364 VP.n120 VSUBS 0.021876f
C1365 VP.n121 VSUBS 0.021876f
C1366 VP.n122 VSUBS 0.040772f
C1367 VP.n123 VSUBS 0.040772f
C1368 VP.n124 VSUBS 0.023058f
C1369 VP.n125 VSUBS 0.035308f
C1370 VP.n126 VSUBS 0.065954f
C1371 VTAIL.t8 VSUBS 0.41004f
C1372 VTAIL.t14 VSUBS 0.41004f
C1373 VTAIL.n0 VSUBS 3.24004f
C1374 VTAIL.n1 VSUBS 1.1327f
C1375 VTAIL.t5 VSUBS 4.22906f
C1376 VTAIL.n2 VSUBS 1.33485f
C1377 VTAIL.t4 VSUBS 0.41004f
C1378 VTAIL.t0 VSUBS 0.41004f
C1379 VTAIL.n3 VSUBS 3.24004f
C1380 VTAIL.n4 VSUBS 1.31955f
C1381 VTAIL.t19 VSUBS 0.41004f
C1382 VTAIL.t1 VSUBS 0.41004f
C1383 VTAIL.n5 VSUBS 3.24004f
C1384 VTAIL.n6 VSUBS 3.45252f
C1385 VTAIL.t11 VSUBS 0.41004f
C1386 VTAIL.t16 VSUBS 0.41004f
C1387 VTAIL.n7 VSUBS 3.24005f
C1388 VTAIL.n8 VSUBS 3.45251f
C1389 VTAIL.t10 VSUBS 0.41004f
C1390 VTAIL.t17 VSUBS 0.41004f
C1391 VTAIL.n9 VSUBS 3.24005f
C1392 VTAIL.n10 VSUBS 1.31955f
C1393 VTAIL.t13 VSUBS 4.22909f
C1394 VTAIL.n11 VSUBS 1.33482f
C1395 VTAIL.t6 VSUBS 0.41004f
C1396 VTAIL.t3 VSUBS 0.41004f
C1397 VTAIL.n12 VSUBS 3.24005f
C1398 VTAIL.n13 VSUBS 1.20557f
C1399 VTAIL.t2 VSUBS 0.41004f
C1400 VTAIL.t18 VSUBS 0.41004f
C1401 VTAIL.n14 VSUBS 3.24005f
C1402 VTAIL.n15 VSUBS 1.31955f
C1403 VTAIL.t7 VSUBS 4.22906f
C1404 VTAIL.n16 VSUBS 3.26933f
C1405 VTAIL.t15 VSUBS 4.22906f
C1406 VTAIL.n17 VSUBS 3.26933f
C1407 VTAIL.t12 VSUBS 0.41004f
C1408 VTAIL.t9 VSUBS 0.41004f
C1409 VTAIL.n18 VSUBS 3.24004f
C1410 VTAIL.n19 VSUBS 1.07997f
C1411 VDD2.t6 VSUBS 4.64936f
C1412 VDD2.t4 VSUBS 0.425612f
C1413 VDD2.t2 VSUBS 0.425612f
C1414 VDD2.n0 VSUBS 3.54733f
C1415 VDD2.n1 VSUBS 1.94809f
C1416 VDD2.t7 VSUBS 0.425612f
C1417 VDD2.t5 VSUBS 0.425612f
C1418 VDD2.n2 VSUBS 3.58872f
C1419 VDD2.n3 VSUBS 4.83985f
C1420 VDD2.t1 VSUBS 4.60126f
C1421 VDD2.n4 VSUBS 5.06455f
C1422 VDD2.t8 VSUBS 0.425612f
C1423 VDD2.t0 VSUBS 0.425612f
C1424 VDD2.n5 VSUBS 3.54733f
C1425 VDD2.n6 VSUBS 0.986989f
C1426 VDD2.t9 VSUBS 0.425612f
C1427 VDD2.t3 VSUBS 0.425612f
C1428 VDD2.n7 VSUBS 3.58865f
C1429 VN.t2 VSUBS 3.87245f
C1430 VN.n0 VSUBS 1.40813f
C1431 VN.n1 VSUBS 0.020456f
C1432 VN.n2 VSUBS 0.039494f
C1433 VN.n3 VSUBS 0.020456f
C1434 VN.n4 VSUBS 0.036996f
C1435 VN.n5 VSUBS 0.020456f
C1436 VN.n6 VSUBS 0.040321f
C1437 VN.n7 VSUBS 0.020456f
C1438 VN.n8 VSUBS 0.038125f
C1439 VN.n9 VSUBS 0.020456f
C1440 VN.t5 VSUBS 3.87245f
C1441 VN.n10 VSUBS 0.040935f
C1442 VN.n11 VSUBS 0.020456f
C1443 VN.n12 VSUBS 0.038125f
C1444 VN.t9 VSUBS 4.18269f
C1445 VN.n13 VSUBS 1.34234f
C1446 VN.t3 VSUBS 3.87245f
C1447 VN.n14 VSUBS 1.39833f
C1448 VN.n15 VSUBS 0.020432f
C1449 VN.n16 VSUBS 0.259953f
C1450 VN.n17 VSUBS 0.020456f
C1451 VN.n18 VSUBS 0.020456f
C1452 VN.n19 VSUBS 0.038125f
C1453 VN.n20 VSUBS 0.040321f
C1454 VN.n21 VSUBS 0.016597f
C1455 VN.n22 VSUBS 0.020456f
C1456 VN.n23 VSUBS 0.020456f
C1457 VN.n24 VSUBS 0.020456f
C1458 VN.n25 VSUBS 0.038125f
C1459 VN.n26 VSUBS 0.038125f
C1460 VN.n27 VSUBS 1.35251f
C1461 VN.n28 VSUBS 0.020456f
C1462 VN.n29 VSUBS 0.020456f
C1463 VN.n30 VSUBS 0.020456f
C1464 VN.n31 VSUBS 0.038125f
C1465 VN.n32 VSUBS 0.040935f
C1466 VN.n33 VSUBS 0.016597f
C1467 VN.n34 VSUBS 0.020456f
C1468 VN.n35 VSUBS 0.020456f
C1469 VN.n36 VSUBS 0.020456f
C1470 VN.n37 VSUBS 0.038125f
C1471 VN.n38 VSUBS 0.038125f
C1472 VN.t8 VSUBS 3.87245f
C1473 VN.n39 VSUBS 1.33321f
C1474 VN.n40 VSUBS 0.020432f
C1475 VN.n41 VSUBS 0.020456f
C1476 VN.n42 VSUBS 0.020456f
C1477 VN.n43 VSUBS 0.020456f
C1478 VN.n44 VSUBS 0.038125f
C1479 VN.n45 VSUBS 0.041283f
C1480 VN.n46 VSUBS 0.017076f
C1481 VN.n47 VSUBS 0.020456f
C1482 VN.n48 VSUBS 0.020456f
C1483 VN.n49 VSUBS 0.020456f
C1484 VN.n50 VSUBS 0.038125f
C1485 VN.n51 VSUBS 0.038125f
C1486 VN.n52 VSUBS 0.021561f
C1487 VN.n53 VSUBS 0.033016f
C1488 VN.n54 VSUBS 0.061672f
C1489 VN.t6 VSUBS 3.87245f
C1490 VN.n55 VSUBS 1.40813f
C1491 VN.n56 VSUBS 0.020456f
C1492 VN.n57 VSUBS 0.039494f
C1493 VN.n58 VSUBS 0.020456f
C1494 VN.n59 VSUBS 0.036996f
C1495 VN.n60 VSUBS 0.020456f
C1496 VN.t1 VSUBS 3.87245f
C1497 VN.n61 VSUBS 1.33321f
C1498 VN.n62 VSUBS 0.040321f
C1499 VN.n63 VSUBS 0.020456f
C1500 VN.n64 VSUBS 0.038125f
C1501 VN.n65 VSUBS 0.020456f
C1502 VN.t7 VSUBS 3.87245f
C1503 VN.n66 VSUBS 0.040935f
C1504 VN.n67 VSUBS 0.020456f
C1505 VN.n68 VSUBS 0.038125f
C1506 VN.t4 VSUBS 4.18269f
C1507 VN.n69 VSUBS 1.34234f
C1508 VN.t0 VSUBS 3.87245f
C1509 VN.n70 VSUBS 1.39833f
C1510 VN.n71 VSUBS 0.020432f
C1511 VN.n72 VSUBS 0.259953f
C1512 VN.n73 VSUBS 0.020456f
C1513 VN.n74 VSUBS 0.020456f
C1514 VN.n75 VSUBS 0.038125f
C1515 VN.n76 VSUBS 0.040321f
C1516 VN.n77 VSUBS 0.016597f
C1517 VN.n78 VSUBS 0.020456f
C1518 VN.n79 VSUBS 0.020456f
C1519 VN.n80 VSUBS 0.020456f
C1520 VN.n81 VSUBS 0.038125f
C1521 VN.n82 VSUBS 0.038125f
C1522 VN.n83 VSUBS 1.35251f
C1523 VN.n84 VSUBS 0.020456f
C1524 VN.n85 VSUBS 0.020456f
C1525 VN.n86 VSUBS 0.020456f
C1526 VN.n87 VSUBS 0.038125f
C1527 VN.n88 VSUBS 0.040935f
C1528 VN.n89 VSUBS 0.016597f
C1529 VN.n90 VSUBS 0.020456f
C1530 VN.n91 VSUBS 0.020456f
C1531 VN.n92 VSUBS 0.020456f
C1532 VN.n93 VSUBS 0.038125f
C1533 VN.n94 VSUBS 0.038125f
C1534 VN.n95 VSUBS 0.020432f
C1535 VN.n96 VSUBS 0.020456f
C1536 VN.n97 VSUBS 0.020456f
C1537 VN.n98 VSUBS 0.020456f
C1538 VN.n99 VSUBS 0.038125f
C1539 VN.n100 VSUBS 0.041283f
C1540 VN.n101 VSUBS 0.017076f
C1541 VN.n102 VSUBS 0.020456f
C1542 VN.n103 VSUBS 0.020456f
C1543 VN.n104 VSUBS 0.020456f
C1544 VN.n105 VSUBS 0.038125f
C1545 VN.n106 VSUBS 0.038125f
C1546 VN.n107 VSUBS 0.021561f
C1547 VN.n108 VSUBS 0.033016f
C1548 VN.n109 VSUBS 1.65477f
.ends

