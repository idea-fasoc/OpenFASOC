* NGSPICE file created from diff_pair_sample_0088.ext - technology: sky130A

.subckt diff_pair_sample_0088 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=0.39
X1 VDD1.t3 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=0.39
X2 VTAIL.t4 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=0.39
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=0.39
X4 VTAIL.t6 VN.t2 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=0.39
X5 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=0.39
X6 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=0.39
X7 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=0.39
X8 VDD2.t0 VN.t3 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=0.39
X9 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53605 pd=15.7 as=5.9943 ps=31.52 w=15.37 l=0.39
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=0 ps=0 w=15.37 l=0.39
X11 VTAIL.t1 VP.t3 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=5.9943 pd=31.52 as=2.53605 ps=15.7 w=15.37 l=0.39
R0 VN.n0 VN.t3 1075.23
R1 VN.n0 VN.t1 1075.23
R2 VN.n1 VN.t0 1075.23
R3 VN.n1 VN.t2 1075.23
R4 VN VN.n1 203.863
R5 VN VN.n0 161.351
R6 VTAIL.n682 VTAIL.n602 289.615
R7 VTAIL.n80 VTAIL.n0 289.615
R8 VTAIL.n166 VTAIL.n86 289.615
R9 VTAIL.n252 VTAIL.n172 289.615
R10 VTAIL.n596 VTAIL.n516 289.615
R11 VTAIL.n510 VTAIL.n430 289.615
R12 VTAIL.n424 VTAIL.n344 289.615
R13 VTAIL.n338 VTAIL.n258 289.615
R14 VTAIL.n631 VTAIL.n630 185
R15 VTAIL.n633 VTAIL.n632 185
R16 VTAIL.n626 VTAIL.n625 185
R17 VTAIL.n639 VTAIL.n638 185
R18 VTAIL.n641 VTAIL.n640 185
R19 VTAIL.n622 VTAIL.n621 185
R20 VTAIL.n647 VTAIL.n646 185
R21 VTAIL.n649 VTAIL.n648 185
R22 VTAIL.n618 VTAIL.n617 185
R23 VTAIL.n655 VTAIL.n654 185
R24 VTAIL.n657 VTAIL.n656 185
R25 VTAIL.n614 VTAIL.n613 185
R26 VTAIL.n663 VTAIL.n662 185
R27 VTAIL.n665 VTAIL.n664 185
R28 VTAIL.n610 VTAIL.n609 185
R29 VTAIL.n672 VTAIL.n671 185
R30 VTAIL.n673 VTAIL.n608 185
R31 VTAIL.n675 VTAIL.n674 185
R32 VTAIL.n606 VTAIL.n605 185
R33 VTAIL.n681 VTAIL.n680 185
R34 VTAIL.n683 VTAIL.n682 185
R35 VTAIL.n29 VTAIL.n28 185
R36 VTAIL.n31 VTAIL.n30 185
R37 VTAIL.n24 VTAIL.n23 185
R38 VTAIL.n37 VTAIL.n36 185
R39 VTAIL.n39 VTAIL.n38 185
R40 VTAIL.n20 VTAIL.n19 185
R41 VTAIL.n45 VTAIL.n44 185
R42 VTAIL.n47 VTAIL.n46 185
R43 VTAIL.n16 VTAIL.n15 185
R44 VTAIL.n53 VTAIL.n52 185
R45 VTAIL.n55 VTAIL.n54 185
R46 VTAIL.n12 VTAIL.n11 185
R47 VTAIL.n61 VTAIL.n60 185
R48 VTAIL.n63 VTAIL.n62 185
R49 VTAIL.n8 VTAIL.n7 185
R50 VTAIL.n70 VTAIL.n69 185
R51 VTAIL.n71 VTAIL.n6 185
R52 VTAIL.n73 VTAIL.n72 185
R53 VTAIL.n4 VTAIL.n3 185
R54 VTAIL.n79 VTAIL.n78 185
R55 VTAIL.n81 VTAIL.n80 185
R56 VTAIL.n115 VTAIL.n114 185
R57 VTAIL.n117 VTAIL.n116 185
R58 VTAIL.n110 VTAIL.n109 185
R59 VTAIL.n123 VTAIL.n122 185
R60 VTAIL.n125 VTAIL.n124 185
R61 VTAIL.n106 VTAIL.n105 185
R62 VTAIL.n131 VTAIL.n130 185
R63 VTAIL.n133 VTAIL.n132 185
R64 VTAIL.n102 VTAIL.n101 185
R65 VTAIL.n139 VTAIL.n138 185
R66 VTAIL.n141 VTAIL.n140 185
R67 VTAIL.n98 VTAIL.n97 185
R68 VTAIL.n147 VTAIL.n146 185
R69 VTAIL.n149 VTAIL.n148 185
R70 VTAIL.n94 VTAIL.n93 185
R71 VTAIL.n156 VTAIL.n155 185
R72 VTAIL.n157 VTAIL.n92 185
R73 VTAIL.n159 VTAIL.n158 185
R74 VTAIL.n90 VTAIL.n89 185
R75 VTAIL.n165 VTAIL.n164 185
R76 VTAIL.n167 VTAIL.n166 185
R77 VTAIL.n201 VTAIL.n200 185
R78 VTAIL.n203 VTAIL.n202 185
R79 VTAIL.n196 VTAIL.n195 185
R80 VTAIL.n209 VTAIL.n208 185
R81 VTAIL.n211 VTAIL.n210 185
R82 VTAIL.n192 VTAIL.n191 185
R83 VTAIL.n217 VTAIL.n216 185
R84 VTAIL.n219 VTAIL.n218 185
R85 VTAIL.n188 VTAIL.n187 185
R86 VTAIL.n225 VTAIL.n224 185
R87 VTAIL.n227 VTAIL.n226 185
R88 VTAIL.n184 VTAIL.n183 185
R89 VTAIL.n233 VTAIL.n232 185
R90 VTAIL.n235 VTAIL.n234 185
R91 VTAIL.n180 VTAIL.n179 185
R92 VTAIL.n242 VTAIL.n241 185
R93 VTAIL.n243 VTAIL.n178 185
R94 VTAIL.n245 VTAIL.n244 185
R95 VTAIL.n176 VTAIL.n175 185
R96 VTAIL.n251 VTAIL.n250 185
R97 VTAIL.n253 VTAIL.n252 185
R98 VTAIL.n597 VTAIL.n596 185
R99 VTAIL.n595 VTAIL.n594 185
R100 VTAIL.n520 VTAIL.n519 185
R101 VTAIL.n524 VTAIL.n522 185
R102 VTAIL.n589 VTAIL.n588 185
R103 VTAIL.n587 VTAIL.n586 185
R104 VTAIL.n526 VTAIL.n525 185
R105 VTAIL.n581 VTAIL.n580 185
R106 VTAIL.n579 VTAIL.n578 185
R107 VTAIL.n530 VTAIL.n529 185
R108 VTAIL.n573 VTAIL.n572 185
R109 VTAIL.n571 VTAIL.n570 185
R110 VTAIL.n534 VTAIL.n533 185
R111 VTAIL.n565 VTAIL.n564 185
R112 VTAIL.n563 VTAIL.n562 185
R113 VTAIL.n538 VTAIL.n537 185
R114 VTAIL.n557 VTAIL.n556 185
R115 VTAIL.n555 VTAIL.n554 185
R116 VTAIL.n542 VTAIL.n541 185
R117 VTAIL.n549 VTAIL.n548 185
R118 VTAIL.n547 VTAIL.n546 185
R119 VTAIL.n511 VTAIL.n510 185
R120 VTAIL.n509 VTAIL.n508 185
R121 VTAIL.n434 VTAIL.n433 185
R122 VTAIL.n438 VTAIL.n436 185
R123 VTAIL.n503 VTAIL.n502 185
R124 VTAIL.n501 VTAIL.n500 185
R125 VTAIL.n440 VTAIL.n439 185
R126 VTAIL.n495 VTAIL.n494 185
R127 VTAIL.n493 VTAIL.n492 185
R128 VTAIL.n444 VTAIL.n443 185
R129 VTAIL.n487 VTAIL.n486 185
R130 VTAIL.n485 VTAIL.n484 185
R131 VTAIL.n448 VTAIL.n447 185
R132 VTAIL.n479 VTAIL.n478 185
R133 VTAIL.n477 VTAIL.n476 185
R134 VTAIL.n452 VTAIL.n451 185
R135 VTAIL.n471 VTAIL.n470 185
R136 VTAIL.n469 VTAIL.n468 185
R137 VTAIL.n456 VTAIL.n455 185
R138 VTAIL.n463 VTAIL.n462 185
R139 VTAIL.n461 VTAIL.n460 185
R140 VTAIL.n425 VTAIL.n424 185
R141 VTAIL.n423 VTAIL.n422 185
R142 VTAIL.n348 VTAIL.n347 185
R143 VTAIL.n352 VTAIL.n350 185
R144 VTAIL.n417 VTAIL.n416 185
R145 VTAIL.n415 VTAIL.n414 185
R146 VTAIL.n354 VTAIL.n353 185
R147 VTAIL.n409 VTAIL.n408 185
R148 VTAIL.n407 VTAIL.n406 185
R149 VTAIL.n358 VTAIL.n357 185
R150 VTAIL.n401 VTAIL.n400 185
R151 VTAIL.n399 VTAIL.n398 185
R152 VTAIL.n362 VTAIL.n361 185
R153 VTAIL.n393 VTAIL.n392 185
R154 VTAIL.n391 VTAIL.n390 185
R155 VTAIL.n366 VTAIL.n365 185
R156 VTAIL.n385 VTAIL.n384 185
R157 VTAIL.n383 VTAIL.n382 185
R158 VTAIL.n370 VTAIL.n369 185
R159 VTAIL.n377 VTAIL.n376 185
R160 VTAIL.n375 VTAIL.n374 185
R161 VTAIL.n339 VTAIL.n338 185
R162 VTAIL.n337 VTAIL.n336 185
R163 VTAIL.n262 VTAIL.n261 185
R164 VTAIL.n266 VTAIL.n264 185
R165 VTAIL.n331 VTAIL.n330 185
R166 VTAIL.n329 VTAIL.n328 185
R167 VTAIL.n268 VTAIL.n267 185
R168 VTAIL.n323 VTAIL.n322 185
R169 VTAIL.n321 VTAIL.n320 185
R170 VTAIL.n272 VTAIL.n271 185
R171 VTAIL.n315 VTAIL.n314 185
R172 VTAIL.n313 VTAIL.n312 185
R173 VTAIL.n276 VTAIL.n275 185
R174 VTAIL.n307 VTAIL.n306 185
R175 VTAIL.n305 VTAIL.n304 185
R176 VTAIL.n280 VTAIL.n279 185
R177 VTAIL.n299 VTAIL.n298 185
R178 VTAIL.n297 VTAIL.n296 185
R179 VTAIL.n284 VTAIL.n283 185
R180 VTAIL.n291 VTAIL.n290 185
R181 VTAIL.n289 VTAIL.n288 185
R182 VTAIL.n629 VTAIL.t5 147.659
R183 VTAIL.n27 VTAIL.t4 147.659
R184 VTAIL.n113 VTAIL.t3 147.659
R185 VTAIL.n199 VTAIL.t0 147.659
R186 VTAIL.n545 VTAIL.t2 147.659
R187 VTAIL.n459 VTAIL.t1 147.659
R188 VTAIL.n373 VTAIL.t7 147.659
R189 VTAIL.n287 VTAIL.t6 147.659
R190 VTAIL.n632 VTAIL.n631 104.615
R191 VTAIL.n632 VTAIL.n625 104.615
R192 VTAIL.n639 VTAIL.n625 104.615
R193 VTAIL.n640 VTAIL.n639 104.615
R194 VTAIL.n640 VTAIL.n621 104.615
R195 VTAIL.n647 VTAIL.n621 104.615
R196 VTAIL.n648 VTAIL.n647 104.615
R197 VTAIL.n648 VTAIL.n617 104.615
R198 VTAIL.n655 VTAIL.n617 104.615
R199 VTAIL.n656 VTAIL.n655 104.615
R200 VTAIL.n656 VTAIL.n613 104.615
R201 VTAIL.n663 VTAIL.n613 104.615
R202 VTAIL.n664 VTAIL.n663 104.615
R203 VTAIL.n664 VTAIL.n609 104.615
R204 VTAIL.n672 VTAIL.n609 104.615
R205 VTAIL.n673 VTAIL.n672 104.615
R206 VTAIL.n674 VTAIL.n673 104.615
R207 VTAIL.n674 VTAIL.n605 104.615
R208 VTAIL.n681 VTAIL.n605 104.615
R209 VTAIL.n682 VTAIL.n681 104.615
R210 VTAIL.n30 VTAIL.n29 104.615
R211 VTAIL.n30 VTAIL.n23 104.615
R212 VTAIL.n37 VTAIL.n23 104.615
R213 VTAIL.n38 VTAIL.n37 104.615
R214 VTAIL.n38 VTAIL.n19 104.615
R215 VTAIL.n45 VTAIL.n19 104.615
R216 VTAIL.n46 VTAIL.n45 104.615
R217 VTAIL.n46 VTAIL.n15 104.615
R218 VTAIL.n53 VTAIL.n15 104.615
R219 VTAIL.n54 VTAIL.n53 104.615
R220 VTAIL.n54 VTAIL.n11 104.615
R221 VTAIL.n61 VTAIL.n11 104.615
R222 VTAIL.n62 VTAIL.n61 104.615
R223 VTAIL.n62 VTAIL.n7 104.615
R224 VTAIL.n70 VTAIL.n7 104.615
R225 VTAIL.n71 VTAIL.n70 104.615
R226 VTAIL.n72 VTAIL.n71 104.615
R227 VTAIL.n72 VTAIL.n3 104.615
R228 VTAIL.n79 VTAIL.n3 104.615
R229 VTAIL.n80 VTAIL.n79 104.615
R230 VTAIL.n116 VTAIL.n115 104.615
R231 VTAIL.n116 VTAIL.n109 104.615
R232 VTAIL.n123 VTAIL.n109 104.615
R233 VTAIL.n124 VTAIL.n123 104.615
R234 VTAIL.n124 VTAIL.n105 104.615
R235 VTAIL.n131 VTAIL.n105 104.615
R236 VTAIL.n132 VTAIL.n131 104.615
R237 VTAIL.n132 VTAIL.n101 104.615
R238 VTAIL.n139 VTAIL.n101 104.615
R239 VTAIL.n140 VTAIL.n139 104.615
R240 VTAIL.n140 VTAIL.n97 104.615
R241 VTAIL.n147 VTAIL.n97 104.615
R242 VTAIL.n148 VTAIL.n147 104.615
R243 VTAIL.n148 VTAIL.n93 104.615
R244 VTAIL.n156 VTAIL.n93 104.615
R245 VTAIL.n157 VTAIL.n156 104.615
R246 VTAIL.n158 VTAIL.n157 104.615
R247 VTAIL.n158 VTAIL.n89 104.615
R248 VTAIL.n165 VTAIL.n89 104.615
R249 VTAIL.n166 VTAIL.n165 104.615
R250 VTAIL.n202 VTAIL.n201 104.615
R251 VTAIL.n202 VTAIL.n195 104.615
R252 VTAIL.n209 VTAIL.n195 104.615
R253 VTAIL.n210 VTAIL.n209 104.615
R254 VTAIL.n210 VTAIL.n191 104.615
R255 VTAIL.n217 VTAIL.n191 104.615
R256 VTAIL.n218 VTAIL.n217 104.615
R257 VTAIL.n218 VTAIL.n187 104.615
R258 VTAIL.n225 VTAIL.n187 104.615
R259 VTAIL.n226 VTAIL.n225 104.615
R260 VTAIL.n226 VTAIL.n183 104.615
R261 VTAIL.n233 VTAIL.n183 104.615
R262 VTAIL.n234 VTAIL.n233 104.615
R263 VTAIL.n234 VTAIL.n179 104.615
R264 VTAIL.n242 VTAIL.n179 104.615
R265 VTAIL.n243 VTAIL.n242 104.615
R266 VTAIL.n244 VTAIL.n243 104.615
R267 VTAIL.n244 VTAIL.n175 104.615
R268 VTAIL.n251 VTAIL.n175 104.615
R269 VTAIL.n252 VTAIL.n251 104.615
R270 VTAIL.n596 VTAIL.n595 104.615
R271 VTAIL.n595 VTAIL.n519 104.615
R272 VTAIL.n524 VTAIL.n519 104.615
R273 VTAIL.n588 VTAIL.n524 104.615
R274 VTAIL.n588 VTAIL.n587 104.615
R275 VTAIL.n587 VTAIL.n525 104.615
R276 VTAIL.n580 VTAIL.n525 104.615
R277 VTAIL.n580 VTAIL.n579 104.615
R278 VTAIL.n579 VTAIL.n529 104.615
R279 VTAIL.n572 VTAIL.n529 104.615
R280 VTAIL.n572 VTAIL.n571 104.615
R281 VTAIL.n571 VTAIL.n533 104.615
R282 VTAIL.n564 VTAIL.n533 104.615
R283 VTAIL.n564 VTAIL.n563 104.615
R284 VTAIL.n563 VTAIL.n537 104.615
R285 VTAIL.n556 VTAIL.n537 104.615
R286 VTAIL.n556 VTAIL.n555 104.615
R287 VTAIL.n555 VTAIL.n541 104.615
R288 VTAIL.n548 VTAIL.n541 104.615
R289 VTAIL.n548 VTAIL.n547 104.615
R290 VTAIL.n510 VTAIL.n509 104.615
R291 VTAIL.n509 VTAIL.n433 104.615
R292 VTAIL.n438 VTAIL.n433 104.615
R293 VTAIL.n502 VTAIL.n438 104.615
R294 VTAIL.n502 VTAIL.n501 104.615
R295 VTAIL.n501 VTAIL.n439 104.615
R296 VTAIL.n494 VTAIL.n439 104.615
R297 VTAIL.n494 VTAIL.n493 104.615
R298 VTAIL.n493 VTAIL.n443 104.615
R299 VTAIL.n486 VTAIL.n443 104.615
R300 VTAIL.n486 VTAIL.n485 104.615
R301 VTAIL.n485 VTAIL.n447 104.615
R302 VTAIL.n478 VTAIL.n447 104.615
R303 VTAIL.n478 VTAIL.n477 104.615
R304 VTAIL.n477 VTAIL.n451 104.615
R305 VTAIL.n470 VTAIL.n451 104.615
R306 VTAIL.n470 VTAIL.n469 104.615
R307 VTAIL.n469 VTAIL.n455 104.615
R308 VTAIL.n462 VTAIL.n455 104.615
R309 VTAIL.n462 VTAIL.n461 104.615
R310 VTAIL.n424 VTAIL.n423 104.615
R311 VTAIL.n423 VTAIL.n347 104.615
R312 VTAIL.n352 VTAIL.n347 104.615
R313 VTAIL.n416 VTAIL.n352 104.615
R314 VTAIL.n416 VTAIL.n415 104.615
R315 VTAIL.n415 VTAIL.n353 104.615
R316 VTAIL.n408 VTAIL.n353 104.615
R317 VTAIL.n408 VTAIL.n407 104.615
R318 VTAIL.n407 VTAIL.n357 104.615
R319 VTAIL.n400 VTAIL.n357 104.615
R320 VTAIL.n400 VTAIL.n399 104.615
R321 VTAIL.n399 VTAIL.n361 104.615
R322 VTAIL.n392 VTAIL.n361 104.615
R323 VTAIL.n392 VTAIL.n391 104.615
R324 VTAIL.n391 VTAIL.n365 104.615
R325 VTAIL.n384 VTAIL.n365 104.615
R326 VTAIL.n384 VTAIL.n383 104.615
R327 VTAIL.n383 VTAIL.n369 104.615
R328 VTAIL.n376 VTAIL.n369 104.615
R329 VTAIL.n376 VTAIL.n375 104.615
R330 VTAIL.n338 VTAIL.n337 104.615
R331 VTAIL.n337 VTAIL.n261 104.615
R332 VTAIL.n266 VTAIL.n261 104.615
R333 VTAIL.n330 VTAIL.n266 104.615
R334 VTAIL.n330 VTAIL.n329 104.615
R335 VTAIL.n329 VTAIL.n267 104.615
R336 VTAIL.n322 VTAIL.n267 104.615
R337 VTAIL.n322 VTAIL.n321 104.615
R338 VTAIL.n321 VTAIL.n271 104.615
R339 VTAIL.n314 VTAIL.n271 104.615
R340 VTAIL.n314 VTAIL.n313 104.615
R341 VTAIL.n313 VTAIL.n275 104.615
R342 VTAIL.n306 VTAIL.n275 104.615
R343 VTAIL.n306 VTAIL.n305 104.615
R344 VTAIL.n305 VTAIL.n279 104.615
R345 VTAIL.n298 VTAIL.n279 104.615
R346 VTAIL.n298 VTAIL.n297 104.615
R347 VTAIL.n297 VTAIL.n283 104.615
R348 VTAIL.n290 VTAIL.n283 104.615
R349 VTAIL.n290 VTAIL.n289 104.615
R350 VTAIL.n631 VTAIL.t5 52.3082
R351 VTAIL.n29 VTAIL.t4 52.3082
R352 VTAIL.n115 VTAIL.t3 52.3082
R353 VTAIL.n201 VTAIL.t0 52.3082
R354 VTAIL.n547 VTAIL.t2 52.3082
R355 VTAIL.n461 VTAIL.t1 52.3082
R356 VTAIL.n375 VTAIL.t7 52.3082
R357 VTAIL.n289 VTAIL.t6 52.3082
R358 VTAIL.n687 VTAIL.n686 32.3793
R359 VTAIL.n85 VTAIL.n84 32.3793
R360 VTAIL.n171 VTAIL.n170 32.3793
R361 VTAIL.n257 VTAIL.n256 32.3793
R362 VTAIL.n601 VTAIL.n600 32.3793
R363 VTAIL.n515 VTAIL.n514 32.3793
R364 VTAIL.n429 VTAIL.n428 32.3793
R365 VTAIL.n343 VTAIL.n342 32.3793
R366 VTAIL.n687 VTAIL.n601 26.2548
R367 VTAIL.n343 VTAIL.n257 26.2548
R368 VTAIL.n630 VTAIL.n629 15.6677
R369 VTAIL.n28 VTAIL.n27 15.6677
R370 VTAIL.n114 VTAIL.n113 15.6677
R371 VTAIL.n200 VTAIL.n199 15.6677
R372 VTAIL.n546 VTAIL.n545 15.6677
R373 VTAIL.n460 VTAIL.n459 15.6677
R374 VTAIL.n374 VTAIL.n373 15.6677
R375 VTAIL.n288 VTAIL.n287 15.6677
R376 VTAIL.n675 VTAIL.n606 13.1884
R377 VTAIL.n73 VTAIL.n4 13.1884
R378 VTAIL.n159 VTAIL.n90 13.1884
R379 VTAIL.n245 VTAIL.n176 13.1884
R380 VTAIL.n522 VTAIL.n520 13.1884
R381 VTAIL.n436 VTAIL.n434 13.1884
R382 VTAIL.n350 VTAIL.n348 13.1884
R383 VTAIL.n264 VTAIL.n262 13.1884
R384 VTAIL.n633 VTAIL.n628 12.8005
R385 VTAIL.n676 VTAIL.n608 12.8005
R386 VTAIL.n680 VTAIL.n679 12.8005
R387 VTAIL.n31 VTAIL.n26 12.8005
R388 VTAIL.n74 VTAIL.n6 12.8005
R389 VTAIL.n78 VTAIL.n77 12.8005
R390 VTAIL.n117 VTAIL.n112 12.8005
R391 VTAIL.n160 VTAIL.n92 12.8005
R392 VTAIL.n164 VTAIL.n163 12.8005
R393 VTAIL.n203 VTAIL.n198 12.8005
R394 VTAIL.n246 VTAIL.n178 12.8005
R395 VTAIL.n250 VTAIL.n249 12.8005
R396 VTAIL.n594 VTAIL.n593 12.8005
R397 VTAIL.n590 VTAIL.n589 12.8005
R398 VTAIL.n549 VTAIL.n544 12.8005
R399 VTAIL.n508 VTAIL.n507 12.8005
R400 VTAIL.n504 VTAIL.n503 12.8005
R401 VTAIL.n463 VTAIL.n458 12.8005
R402 VTAIL.n422 VTAIL.n421 12.8005
R403 VTAIL.n418 VTAIL.n417 12.8005
R404 VTAIL.n377 VTAIL.n372 12.8005
R405 VTAIL.n336 VTAIL.n335 12.8005
R406 VTAIL.n332 VTAIL.n331 12.8005
R407 VTAIL.n291 VTAIL.n286 12.8005
R408 VTAIL.n634 VTAIL.n626 12.0247
R409 VTAIL.n671 VTAIL.n670 12.0247
R410 VTAIL.n683 VTAIL.n604 12.0247
R411 VTAIL.n32 VTAIL.n24 12.0247
R412 VTAIL.n69 VTAIL.n68 12.0247
R413 VTAIL.n81 VTAIL.n2 12.0247
R414 VTAIL.n118 VTAIL.n110 12.0247
R415 VTAIL.n155 VTAIL.n154 12.0247
R416 VTAIL.n167 VTAIL.n88 12.0247
R417 VTAIL.n204 VTAIL.n196 12.0247
R418 VTAIL.n241 VTAIL.n240 12.0247
R419 VTAIL.n253 VTAIL.n174 12.0247
R420 VTAIL.n597 VTAIL.n518 12.0247
R421 VTAIL.n586 VTAIL.n523 12.0247
R422 VTAIL.n550 VTAIL.n542 12.0247
R423 VTAIL.n511 VTAIL.n432 12.0247
R424 VTAIL.n500 VTAIL.n437 12.0247
R425 VTAIL.n464 VTAIL.n456 12.0247
R426 VTAIL.n425 VTAIL.n346 12.0247
R427 VTAIL.n414 VTAIL.n351 12.0247
R428 VTAIL.n378 VTAIL.n370 12.0247
R429 VTAIL.n339 VTAIL.n260 12.0247
R430 VTAIL.n328 VTAIL.n265 12.0247
R431 VTAIL.n292 VTAIL.n284 12.0247
R432 VTAIL.n638 VTAIL.n637 11.249
R433 VTAIL.n669 VTAIL.n610 11.249
R434 VTAIL.n684 VTAIL.n602 11.249
R435 VTAIL.n36 VTAIL.n35 11.249
R436 VTAIL.n67 VTAIL.n8 11.249
R437 VTAIL.n82 VTAIL.n0 11.249
R438 VTAIL.n122 VTAIL.n121 11.249
R439 VTAIL.n153 VTAIL.n94 11.249
R440 VTAIL.n168 VTAIL.n86 11.249
R441 VTAIL.n208 VTAIL.n207 11.249
R442 VTAIL.n239 VTAIL.n180 11.249
R443 VTAIL.n254 VTAIL.n172 11.249
R444 VTAIL.n598 VTAIL.n516 11.249
R445 VTAIL.n585 VTAIL.n526 11.249
R446 VTAIL.n554 VTAIL.n553 11.249
R447 VTAIL.n512 VTAIL.n430 11.249
R448 VTAIL.n499 VTAIL.n440 11.249
R449 VTAIL.n468 VTAIL.n467 11.249
R450 VTAIL.n426 VTAIL.n344 11.249
R451 VTAIL.n413 VTAIL.n354 11.249
R452 VTAIL.n382 VTAIL.n381 11.249
R453 VTAIL.n340 VTAIL.n258 11.249
R454 VTAIL.n327 VTAIL.n268 11.249
R455 VTAIL.n296 VTAIL.n295 11.249
R456 VTAIL.n641 VTAIL.n624 10.4732
R457 VTAIL.n666 VTAIL.n665 10.4732
R458 VTAIL.n39 VTAIL.n22 10.4732
R459 VTAIL.n64 VTAIL.n63 10.4732
R460 VTAIL.n125 VTAIL.n108 10.4732
R461 VTAIL.n150 VTAIL.n149 10.4732
R462 VTAIL.n211 VTAIL.n194 10.4732
R463 VTAIL.n236 VTAIL.n235 10.4732
R464 VTAIL.n582 VTAIL.n581 10.4732
R465 VTAIL.n557 VTAIL.n540 10.4732
R466 VTAIL.n496 VTAIL.n495 10.4732
R467 VTAIL.n471 VTAIL.n454 10.4732
R468 VTAIL.n410 VTAIL.n409 10.4732
R469 VTAIL.n385 VTAIL.n368 10.4732
R470 VTAIL.n324 VTAIL.n323 10.4732
R471 VTAIL.n299 VTAIL.n282 10.4732
R472 VTAIL.n642 VTAIL.n622 9.69747
R473 VTAIL.n662 VTAIL.n612 9.69747
R474 VTAIL.n40 VTAIL.n20 9.69747
R475 VTAIL.n60 VTAIL.n10 9.69747
R476 VTAIL.n126 VTAIL.n106 9.69747
R477 VTAIL.n146 VTAIL.n96 9.69747
R478 VTAIL.n212 VTAIL.n192 9.69747
R479 VTAIL.n232 VTAIL.n182 9.69747
R480 VTAIL.n578 VTAIL.n528 9.69747
R481 VTAIL.n558 VTAIL.n538 9.69747
R482 VTAIL.n492 VTAIL.n442 9.69747
R483 VTAIL.n472 VTAIL.n452 9.69747
R484 VTAIL.n406 VTAIL.n356 9.69747
R485 VTAIL.n386 VTAIL.n366 9.69747
R486 VTAIL.n320 VTAIL.n270 9.69747
R487 VTAIL.n300 VTAIL.n280 9.69747
R488 VTAIL.n686 VTAIL.n685 9.45567
R489 VTAIL.n84 VTAIL.n83 9.45567
R490 VTAIL.n170 VTAIL.n169 9.45567
R491 VTAIL.n256 VTAIL.n255 9.45567
R492 VTAIL.n600 VTAIL.n599 9.45567
R493 VTAIL.n514 VTAIL.n513 9.45567
R494 VTAIL.n428 VTAIL.n427 9.45567
R495 VTAIL.n342 VTAIL.n341 9.45567
R496 VTAIL.n685 VTAIL.n684 9.3005
R497 VTAIL.n604 VTAIL.n603 9.3005
R498 VTAIL.n679 VTAIL.n678 9.3005
R499 VTAIL.n651 VTAIL.n650 9.3005
R500 VTAIL.n620 VTAIL.n619 9.3005
R501 VTAIL.n645 VTAIL.n644 9.3005
R502 VTAIL.n643 VTAIL.n642 9.3005
R503 VTAIL.n624 VTAIL.n623 9.3005
R504 VTAIL.n637 VTAIL.n636 9.3005
R505 VTAIL.n635 VTAIL.n634 9.3005
R506 VTAIL.n628 VTAIL.n627 9.3005
R507 VTAIL.n653 VTAIL.n652 9.3005
R508 VTAIL.n616 VTAIL.n615 9.3005
R509 VTAIL.n659 VTAIL.n658 9.3005
R510 VTAIL.n661 VTAIL.n660 9.3005
R511 VTAIL.n612 VTAIL.n611 9.3005
R512 VTAIL.n667 VTAIL.n666 9.3005
R513 VTAIL.n669 VTAIL.n668 9.3005
R514 VTAIL.n670 VTAIL.n607 9.3005
R515 VTAIL.n677 VTAIL.n676 9.3005
R516 VTAIL.n83 VTAIL.n82 9.3005
R517 VTAIL.n2 VTAIL.n1 9.3005
R518 VTAIL.n77 VTAIL.n76 9.3005
R519 VTAIL.n49 VTAIL.n48 9.3005
R520 VTAIL.n18 VTAIL.n17 9.3005
R521 VTAIL.n43 VTAIL.n42 9.3005
R522 VTAIL.n41 VTAIL.n40 9.3005
R523 VTAIL.n22 VTAIL.n21 9.3005
R524 VTAIL.n35 VTAIL.n34 9.3005
R525 VTAIL.n33 VTAIL.n32 9.3005
R526 VTAIL.n26 VTAIL.n25 9.3005
R527 VTAIL.n51 VTAIL.n50 9.3005
R528 VTAIL.n14 VTAIL.n13 9.3005
R529 VTAIL.n57 VTAIL.n56 9.3005
R530 VTAIL.n59 VTAIL.n58 9.3005
R531 VTAIL.n10 VTAIL.n9 9.3005
R532 VTAIL.n65 VTAIL.n64 9.3005
R533 VTAIL.n67 VTAIL.n66 9.3005
R534 VTAIL.n68 VTAIL.n5 9.3005
R535 VTAIL.n75 VTAIL.n74 9.3005
R536 VTAIL.n169 VTAIL.n168 9.3005
R537 VTAIL.n88 VTAIL.n87 9.3005
R538 VTAIL.n163 VTAIL.n162 9.3005
R539 VTAIL.n135 VTAIL.n134 9.3005
R540 VTAIL.n104 VTAIL.n103 9.3005
R541 VTAIL.n129 VTAIL.n128 9.3005
R542 VTAIL.n127 VTAIL.n126 9.3005
R543 VTAIL.n108 VTAIL.n107 9.3005
R544 VTAIL.n121 VTAIL.n120 9.3005
R545 VTAIL.n119 VTAIL.n118 9.3005
R546 VTAIL.n112 VTAIL.n111 9.3005
R547 VTAIL.n137 VTAIL.n136 9.3005
R548 VTAIL.n100 VTAIL.n99 9.3005
R549 VTAIL.n143 VTAIL.n142 9.3005
R550 VTAIL.n145 VTAIL.n144 9.3005
R551 VTAIL.n96 VTAIL.n95 9.3005
R552 VTAIL.n151 VTAIL.n150 9.3005
R553 VTAIL.n153 VTAIL.n152 9.3005
R554 VTAIL.n154 VTAIL.n91 9.3005
R555 VTAIL.n161 VTAIL.n160 9.3005
R556 VTAIL.n255 VTAIL.n254 9.3005
R557 VTAIL.n174 VTAIL.n173 9.3005
R558 VTAIL.n249 VTAIL.n248 9.3005
R559 VTAIL.n221 VTAIL.n220 9.3005
R560 VTAIL.n190 VTAIL.n189 9.3005
R561 VTAIL.n215 VTAIL.n214 9.3005
R562 VTAIL.n213 VTAIL.n212 9.3005
R563 VTAIL.n194 VTAIL.n193 9.3005
R564 VTAIL.n207 VTAIL.n206 9.3005
R565 VTAIL.n205 VTAIL.n204 9.3005
R566 VTAIL.n198 VTAIL.n197 9.3005
R567 VTAIL.n223 VTAIL.n222 9.3005
R568 VTAIL.n186 VTAIL.n185 9.3005
R569 VTAIL.n229 VTAIL.n228 9.3005
R570 VTAIL.n231 VTAIL.n230 9.3005
R571 VTAIL.n182 VTAIL.n181 9.3005
R572 VTAIL.n237 VTAIL.n236 9.3005
R573 VTAIL.n239 VTAIL.n238 9.3005
R574 VTAIL.n240 VTAIL.n177 9.3005
R575 VTAIL.n247 VTAIL.n246 9.3005
R576 VTAIL.n532 VTAIL.n531 9.3005
R577 VTAIL.n575 VTAIL.n574 9.3005
R578 VTAIL.n577 VTAIL.n576 9.3005
R579 VTAIL.n528 VTAIL.n527 9.3005
R580 VTAIL.n583 VTAIL.n582 9.3005
R581 VTAIL.n585 VTAIL.n584 9.3005
R582 VTAIL.n523 VTAIL.n521 9.3005
R583 VTAIL.n591 VTAIL.n590 9.3005
R584 VTAIL.n599 VTAIL.n598 9.3005
R585 VTAIL.n518 VTAIL.n517 9.3005
R586 VTAIL.n593 VTAIL.n592 9.3005
R587 VTAIL.n569 VTAIL.n568 9.3005
R588 VTAIL.n567 VTAIL.n566 9.3005
R589 VTAIL.n536 VTAIL.n535 9.3005
R590 VTAIL.n561 VTAIL.n560 9.3005
R591 VTAIL.n559 VTAIL.n558 9.3005
R592 VTAIL.n540 VTAIL.n539 9.3005
R593 VTAIL.n553 VTAIL.n552 9.3005
R594 VTAIL.n551 VTAIL.n550 9.3005
R595 VTAIL.n544 VTAIL.n543 9.3005
R596 VTAIL.n446 VTAIL.n445 9.3005
R597 VTAIL.n489 VTAIL.n488 9.3005
R598 VTAIL.n491 VTAIL.n490 9.3005
R599 VTAIL.n442 VTAIL.n441 9.3005
R600 VTAIL.n497 VTAIL.n496 9.3005
R601 VTAIL.n499 VTAIL.n498 9.3005
R602 VTAIL.n437 VTAIL.n435 9.3005
R603 VTAIL.n505 VTAIL.n504 9.3005
R604 VTAIL.n513 VTAIL.n512 9.3005
R605 VTAIL.n432 VTAIL.n431 9.3005
R606 VTAIL.n507 VTAIL.n506 9.3005
R607 VTAIL.n483 VTAIL.n482 9.3005
R608 VTAIL.n481 VTAIL.n480 9.3005
R609 VTAIL.n450 VTAIL.n449 9.3005
R610 VTAIL.n475 VTAIL.n474 9.3005
R611 VTAIL.n473 VTAIL.n472 9.3005
R612 VTAIL.n454 VTAIL.n453 9.3005
R613 VTAIL.n467 VTAIL.n466 9.3005
R614 VTAIL.n465 VTAIL.n464 9.3005
R615 VTAIL.n458 VTAIL.n457 9.3005
R616 VTAIL.n360 VTAIL.n359 9.3005
R617 VTAIL.n403 VTAIL.n402 9.3005
R618 VTAIL.n405 VTAIL.n404 9.3005
R619 VTAIL.n356 VTAIL.n355 9.3005
R620 VTAIL.n411 VTAIL.n410 9.3005
R621 VTAIL.n413 VTAIL.n412 9.3005
R622 VTAIL.n351 VTAIL.n349 9.3005
R623 VTAIL.n419 VTAIL.n418 9.3005
R624 VTAIL.n427 VTAIL.n426 9.3005
R625 VTAIL.n346 VTAIL.n345 9.3005
R626 VTAIL.n421 VTAIL.n420 9.3005
R627 VTAIL.n397 VTAIL.n396 9.3005
R628 VTAIL.n395 VTAIL.n394 9.3005
R629 VTAIL.n364 VTAIL.n363 9.3005
R630 VTAIL.n389 VTAIL.n388 9.3005
R631 VTAIL.n387 VTAIL.n386 9.3005
R632 VTAIL.n368 VTAIL.n367 9.3005
R633 VTAIL.n381 VTAIL.n380 9.3005
R634 VTAIL.n379 VTAIL.n378 9.3005
R635 VTAIL.n372 VTAIL.n371 9.3005
R636 VTAIL.n274 VTAIL.n273 9.3005
R637 VTAIL.n317 VTAIL.n316 9.3005
R638 VTAIL.n319 VTAIL.n318 9.3005
R639 VTAIL.n270 VTAIL.n269 9.3005
R640 VTAIL.n325 VTAIL.n324 9.3005
R641 VTAIL.n327 VTAIL.n326 9.3005
R642 VTAIL.n265 VTAIL.n263 9.3005
R643 VTAIL.n333 VTAIL.n332 9.3005
R644 VTAIL.n341 VTAIL.n340 9.3005
R645 VTAIL.n260 VTAIL.n259 9.3005
R646 VTAIL.n335 VTAIL.n334 9.3005
R647 VTAIL.n311 VTAIL.n310 9.3005
R648 VTAIL.n309 VTAIL.n308 9.3005
R649 VTAIL.n278 VTAIL.n277 9.3005
R650 VTAIL.n303 VTAIL.n302 9.3005
R651 VTAIL.n301 VTAIL.n300 9.3005
R652 VTAIL.n282 VTAIL.n281 9.3005
R653 VTAIL.n295 VTAIL.n294 9.3005
R654 VTAIL.n293 VTAIL.n292 9.3005
R655 VTAIL.n286 VTAIL.n285 9.3005
R656 VTAIL.n646 VTAIL.n645 8.92171
R657 VTAIL.n661 VTAIL.n614 8.92171
R658 VTAIL.n44 VTAIL.n43 8.92171
R659 VTAIL.n59 VTAIL.n12 8.92171
R660 VTAIL.n130 VTAIL.n129 8.92171
R661 VTAIL.n145 VTAIL.n98 8.92171
R662 VTAIL.n216 VTAIL.n215 8.92171
R663 VTAIL.n231 VTAIL.n184 8.92171
R664 VTAIL.n577 VTAIL.n530 8.92171
R665 VTAIL.n562 VTAIL.n561 8.92171
R666 VTAIL.n491 VTAIL.n444 8.92171
R667 VTAIL.n476 VTAIL.n475 8.92171
R668 VTAIL.n405 VTAIL.n358 8.92171
R669 VTAIL.n390 VTAIL.n389 8.92171
R670 VTAIL.n319 VTAIL.n272 8.92171
R671 VTAIL.n304 VTAIL.n303 8.92171
R672 VTAIL.n649 VTAIL.n620 8.14595
R673 VTAIL.n658 VTAIL.n657 8.14595
R674 VTAIL.n47 VTAIL.n18 8.14595
R675 VTAIL.n56 VTAIL.n55 8.14595
R676 VTAIL.n133 VTAIL.n104 8.14595
R677 VTAIL.n142 VTAIL.n141 8.14595
R678 VTAIL.n219 VTAIL.n190 8.14595
R679 VTAIL.n228 VTAIL.n227 8.14595
R680 VTAIL.n574 VTAIL.n573 8.14595
R681 VTAIL.n565 VTAIL.n536 8.14595
R682 VTAIL.n488 VTAIL.n487 8.14595
R683 VTAIL.n479 VTAIL.n450 8.14595
R684 VTAIL.n402 VTAIL.n401 8.14595
R685 VTAIL.n393 VTAIL.n364 8.14595
R686 VTAIL.n316 VTAIL.n315 8.14595
R687 VTAIL.n307 VTAIL.n278 8.14595
R688 VTAIL.n650 VTAIL.n618 7.3702
R689 VTAIL.n654 VTAIL.n616 7.3702
R690 VTAIL.n48 VTAIL.n16 7.3702
R691 VTAIL.n52 VTAIL.n14 7.3702
R692 VTAIL.n134 VTAIL.n102 7.3702
R693 VTAIL.n138 VTAIL.n100 7.3702
R694 VTAIL.n220 VTAIL.n188 7.3702
R695 VTAIL.n224 VTAIL.n186 7.3702
R696 VTAIL.n570 VTAIL.n532 7.3702
R697 VTAIL.n566 VTAIL.n534 7.3702
R698 VTAIL.n484 VTAIL.n446 7.3702
R699 VTAIL.n480 VTAIL.n448 7.3702
R700 VTAIL.n398 VTAIL.n360 7.3702
R701 VTAIL.n394 VTAIL.n362 7.3702
R702 VTAIL.n312 VTAIL.n274 7.3702
R703 VTAIL.n308 VTAIL.n276 7.3702
R704 VTAIL.n653 VTAIL.n618 6.59444
R705 VTAIL.n654 VTAIL.n653 6.59444
R706 VTAIL.n51 VTAIL.n16 6.59444
R707 VTAIL.n52 VTAIL.n51 6.59444
R708 VTAIL.n137 VTAIL.n102 6.59444
R709 VTAIL.n138 VTAIL.n137 6.59444
R710 VTAIL.n223 VTAIL.n188 6.59444
R711 VTAIL.n224 VTAIL.n223 6.59444
R712 VTAIL.n570 VTAIL.n569 6.59444
R713 VTAIL.n569 VTAIL.n534 6.59444
R714 VTAIL.n484 VTAIL.n483 6.59444
R715 VTAIL.n483 VTAIL.n448 6.59444
R716 VTAIL.n398 VTAIL.n397 6.59444
R717 VTAIL.n397 VTAIL.n362 6.59444
R718 VTAIL.n312 VTAIL.n311 6.59444
R719 VTAIL.n311 VTAIL.n276 6.59444
R720 VTAIL.n650 VTAIL.n649 5.81868
R721 VTAIL.n657 VTAIL.n616 5.81868
R722 VTAIL.n48 VTAIL.n47 5.81868
R723 VTAIL.n55 VTAIL.n14 5.81868
R724 VTAIL.n134 VTAIL.n133 5.81868
R725 VTAIL.n141 VTAIL.n100 5.81868
R726 VTAIL.n220 VTAIL.n219 5.81868
R727 VTAIL.n227 VTAIL.n186 5.81868
R728 VTAIL.n573 VTAIL.n532 5.81868
R729 VTAIL.n566 VTAIL.n565 5.81868
R730 VTAIL.n487 VTAIL.n446 5.81868
R731 VTAIL.n480 VTAIL.n479 5.81868
R732 VTAIL.n401 VTAIL.n360 5.81868
R733 VTAIL.n394 VTAIL.n393 5.81868
R734 VTAIL.n315 VTAIL.n274 5.81868
R735 VTAIL.n308 VTAIL.n307 5.81868
R736 VTAIL.n646 VTAIL.n620 5.04292
R737 VTAIL.n658 VTAIL.n614 5.04292
R738 VTAIL.n44 VTAIL.n18 5.04292
R739 VTAIL.n56 VTAIL.n12 5.04292
R740 VTAIL.n130 VTAIL.n104 5.04292
R741 VTAIL.n142 VTAIL.n98 5.04292
R742 VTAIL.n216 VTAIL.n190 5.04292
R743 VTAIL.n228 VTAIL.n184 5.04292
R744 VTAIL.n574 VTAIL.n530 5.04292
R745 VTAIL.n562 VTAIL.n536 5.04292
R746 VTAIL.n488 VTAIL.n444 5.04292
R747 VTAIL.n476 VTAIL.n450 5.04292
R748 VTAIL.n402 VTAIL.n358 5.04292
R749 VTAIL.n390 VTAIL.n364 5.04292
R750 VTAIL.n316 VTAIL.n272 5.04292
R751 VTAIL.n304 VTAIL.n278 5.04292
R752 VTAIL.n629 VTAIL.n627 4.38563
R753 VTAIL.n27 VTAIL.n25 4.38563
R754 VTAIL.n113 VTAIL.n111 4.38563
R755 VTAIL.n199 VTAIL.n197 4.38563
R756 VTAIL.n545 VTAIL.n543 4.38563
R757 VTAIL.n459 VTAIL.n457 4.38563
R758 VTAIL.n373 VTAIL.n371 4.38563
R759 VTAIL.n287 VTAIL.n285 4.38563
R760 VTAIL.n645 VTAIL.n622 4.26717
R761 VTAIL.n662 VTAIL.n661 4.26717
R762 VTAIL.n43 VTAIL.n20 4.26717
R763 VTAIL.n60 VTAIL.n59 4.26717
R764 VTAIL.n129 VTAIL.n106 4.26717
R765 VTAIL.n146 VTAIL.n145 4.26717
R766 VTAIL.n215 VTAIL.n192 4.26717
R767 VTAIL.n232 VTAIL.n231 4.26717
R768 VTAIL.n578 VTAIL.n577 4.26717
R769 VTAIL.n561 VTAIL.n538 4.26717
R770 VTAIL.n492 VTAIL.n491 4.26717
R771 VTAIL.n475 VTAIL.n452 4.26717
R772 VTAIL.n406 VTAIL.n405 4.26717
R773 VTAIL.n389 VTAIL.n366 4.26717
R774 VTAIL.n320 VTAIL.n319 4.26717
R775 VTAIL.n303 VTAIL.n280 4.26717
R776 VTAIL.n642 VTAIL.n641 3.49141
R777 VTAIL.n665 VTAIL.n612 3.49141
R778 VTAIL.n40 VTAIL.n39 3.49141
R779 VTAIL.n63 VTAIL.n10 3.49141
R780 VTAIL.n126 VTAIL.n125 3.49141
R781 VTAIL.n149 VTAIL.n96 3.49141
R782 VTAIL.n212 VTAIL.n211 3.49141
R783 VTAIL.n235 VTAIL.n182 3.49141
R784 VTAIL.n581 VTAIL.n528 3.49141
R785 VTAIL.n558 VTAIL.n557 3.49141
R786 VTAIL.n495 VTAIL.n442 3.49141
R787 VTAIL.n472 VTAIL.n471 3.49141
R788 VTAIL.n409 VTAIL.n356 3.49141
R789 VTAIL.n386 VTAIL.n385 3.49141
R790 VTAIL.n323 VTAIL.n270 3.49141
R791 VTAIL.n300 VTAIL.n299 3.49141
R792 VTAIL.n638 VTAIL.n624 2.71565
R793 VTAIL.n666 VTAIL.n610 2.71565
R794 VTAIL.n686 VTAIL.n602 2.71565
R795 VTAIL.n36 VTAIL.n22 2.71565
R796 VTAIL.n64 VTAIL.n8 2.71565
R797 VTAIL.n84 VTAIL.n0 2.71565
R798 VTAIL.n122 VTAIL.n108 2.71565
R799 VTAIL.n150 VTAIL.n94 2.71565
R800 VTAIL.n170 VTAIL.n86 2.71565
R801 VTAIL.n208 VTAIL.n194 2.71565
R802 VTAIL.n236 VTAIL.n180 2.71565
R803 VTAIL.n256 VTAIL.n172 2.71565
R804 VTAIL.n600 VTAIL.n516 2.71565
R805 VTAIL.n582 VTAIL.n526 2.71565
R806 VTAIL.n554 VTAIL.n540 2.71565
R807 VTAIL.n514 VTAIL.n430 2.71565
R808 VTAIL.n496 VTAIL.n440 2.71565
R809 VTAIL.n468 VTAIL.n454 2.71565
R810 VTAIL.n428 VTAIL.n344 2.71565
R811 VTAIL.n410 VTAIL.n354 2.71565
R812 VTAIL.n382 VTAIL.n368 2.71565
R813 VTAIL.n342 VTAIL.n258 2.71565
R814 VTAIL.n324 VTAIL.n268 2.71565
R815 VTAIL.n296 VTAIL.n282 2.71565
R816 VTAIL.n637 VTAIL.n626 1.93989
R817 VTAIL.n671 VTAIL.n669 1.93989
R818 VTAIL.n684 VTAIL.n683 1.93989
R819 VTAIL.n35 VTAIL.n24 1.93989
R820 VTAIL.n69 VTAIL.n67 1.93989
R821 VTAIL.n82 VTAIL.n81 1.93989
R822 VTAIL.n121 VTAIL.n110 1.93989
R823 VTAIL.n155 VTAIL.n153 1.93989
R824 VTAIL.n168 VTAIL.n167 1.93989
R825 VTAIL.n207 VTAIL.n196 1.93989
R826 VTAIL.n241 VTAIL.n239 1.93989
R827 VTAIL.n254 VTAIL.n253 1.93989
R828 VTAIL.n598 VTAIL.n597 1.93989
R829 VTAIL.n586 VTAIL.n585 1.93989
R830 VTAIL.n553 VTAIL.n542 1.93989
R831 VTAIL.n512 VTAIL.n511 1.93989
R832 VTAIL.n500 VTAIL.n499 1.93989
R833 VTAIL.n467 VTAIL.n456 1.93989
R834 VTAIL.n426 VTAIL.n425 1.93989
R835 VTAIL.n414 VTAIL.n413 1.93989
R836 VTAIL.n381 VTAIL.n370 1.93989
R837 VTAIL.n340 VTAIL.n339 1.93989
R838 VTAIL.n328 VTAIL.n327 1.93989
R839 VTAIL.n295 VTAIL.n284 1.93989
R840 VTAIL.n634 VTAIL.n633 1.16414
R841 VTAIL.n670 VTAIL.n608 1.16414
R842 VTAIL.n680 VTAIL.n604 1.16414
R843 VTAIL.n32 VTAIL.n31 1.16414
R844 VTAIL.n68 VTAIL.n6 1.16414
R845 VTAIL.n78 VTAIL.n2 1.16414
R846 VTAIL.n118 VTAIL.n117 1.16414
R847 VTAIL.n154 VTAIL.n92 1.16414
R848 VTAIL.n164 VTAIL.n88 1.16414
R849 VTAIL.n204 VTAIL.n203 1.16414
R850 VTAIL.n240 VTAIL.n178 1.16414
R851 VTAIL.n250 VTAIL.n174 1.16414
R852 VTAIL.n594 VTAIL.n518 1.16414
R853 VTAIL.n589 VTAIL.n523 1.16414
R854 VTAIL.n550 VTAIL.n549 1.16414
R855 VTAIL.n508 VTAIL.n432 1.16414
R856 VTAIL.n503 VTAIL.n437 1.16414
R857 VTAIL.n464 VTAIL.n463 1.16414
R858 VTAIL.n422 VTAIL.n346 1.16414
R859 VTAIL.n417 VTAIL.n351 1.16414
R860 VTAIL.n378 VTAIL.n377 1.16414
R861 VTAIL.n336 VTAIL.n260 1.16414
R862 VTAIL.n331 VTAIL.n265 1.16414
R863 VTAIL.n292 VTAIL.n291 1.16414
R864 VTAIL.n429 VTAIL.n343 0.62119
R865 VTAIL.n601 VTAIL.n515 0.62119
R866 VTAIL.n257 VTAIL.n171 0.62119
R867 VTAIL.n515 VTAIL.n429 0.470328
R868 VTAIL.n171 VTAIL.n85 0.470328
R869 VTAIL.n630 VTAIL.n628 0.388379
R870 VTAIL.n676 VTAIL.n675 0.388379
R871 VTAIL.n679 VTAIL.n606 0.388379
R872 VTAIL.n28 VTAIL.n26 0.388379
R873 VTAIL.n74 VTAIL.n73 0.388379
R874 VTAIL.n77 VTAIL.n4 0.388379
R875 VTAIL.n114 VTAIL.n112 0.388379
R876 VTAIL.n160 VTAIL.n159 0.388379
R877 VTAIL.n163 VTAIL.n90 0.388379
R878 VTAIL.n200 VTAIL.n198 0.388379
R879 VTAIL.n246 VTAIL.n245 0.388379
R880 VTAIL.n249 VTAIL.n176 0.388379
R881 VTAIL.n593 VTAIL.n520 0.388379
R882 VTAIL.n590 VTAIL.n522 0.388379
R883 VTAIL.n546 VTAIL.n544 0.388379
R884 VTAIL.n507 VTAIL.n434 0.388379
R885 VTAIL.n504 VTAIL.n436 0.388379
R886 VTAIL.n460 VTAIL.n458 0.388379
R887 VTAIL.n421 VTAIL.n348 0.388379
R888 VTAIL.n418 VTAIL.n350 0.388379
R889 VTAIL.n374 VTAIL.n372 0.388379
R890 VTAIL.n335 VTAIL.n262 0.388379
R891 VTAIL.n332 VTAIL.n264 0.388379
R892 VTAIL.n288 VTAIL.n286 0.388379
R893 VTAIL VTAIL.n85 0.369034
R894 VTAIL VTAIL.n687 0.252655
R895 VTAIL.n635 VTAIL.n627 0.155672
R896 VTAIL.n636 VTAIL.n635 0.155672
R897 VTAIL.n636 VTAIL.n623 0.155672
R898 VTAIL.n643 VTAIL.n623 0.155672
R899 VTAIL.n644 VTAIL.n643 0.155672
R900 VTAIL.n644 VTAIL.n619 0.155672
R901 VTAIL.n651 VTAIL.n619 0.155672
R902 VTAIL.n652 VTAIL.n651 0.155672
R903 VTAIL.n652 VTAIL.n615 0.155672
R904 VTAIL.n659 VTAIL.n615 0.155672
R905 VTAIL.n660 VTAIL.n659 0.155672
R906 VTAIL.n660 VTAIL.n611 0.155672
R907 VTAIL.n667 VTAIL.n611 0.155672
R908 VTAIL.n668 VTAIL.n667 0.155672
R909 VTAIL.n668 VTAIL.n607 0.155672
R910 VTAIL.n677 VTAIL.n607 0.155672
R911 VTAIL.n678 VTAIL.n677 0.155672
R912 VTAIL.n678 VTAIL.n603 0.155672
R913 VTAIL.n685 VTAIL.n603 0.155672
R914 VTAIL.n33 VTAIL.n25 0.155672
R915 VTAIL.n34 VTAIL.n33 0.155672
R916 VTAIL.n34 VTAIL.n21 0.155672
R917 VTAIL.n41 VTAIL.n21 0.155672
R918 VTAIL.n42 VTAIL.n41 0.155672
R919 VTAIL.n42 VTAIL.n17 0.155672
R920 VTAIL.n49 VTAIL.n17 0.155672
R921 VTAIL.n50 VTAIL.n49 0.155672
R922 VTAIL.n50 VTAIL.n13 0.155672
R923 VTAIL.n57 VTAIL.n13 0.155672
R924 VTAIL.n58 VTAIL.n57 0.155672
R925 VTAIL.n58 VTAIL.n9 0.155672
R926 VTAIL.n65 VTAIL.n9 0.155672
R927 VTAIL.n66 VTAIL.n65 0.155672
R928 VTAIL.n66 VTAIL.n5 0.155672
R929 VTAIL.n75 VTAIL.n5 0.155672
R930 VTAIL.n76 VTAIL.n75 0.155672
R931 VTAIL.n76 VTAIL.n1 0.155672
R932 VTAIL.n83 VTAIL.n1 0.155672
R933 VTAIL.n119 VTAIL.n111 0.155672
R934 VTAIL.n120 VTAIL.n119 0.155672
R935 VTAIL.n120 VTAIL.n107 0.155672
R936 VTAIL.n127 VTAIL.n107 0.155672
R937 VTAIL.n128 VTAIL.n127 0.155672
R938 VTAIL.n128 VTAIL.n103 0.155672
R939 VTAIL.n135 VTAIL.n103 0.155672
R940 VTAIL.n136 VTAIL.n135 0.155672
R941 VTAIL.n136 VTAIL.n99 0.155672
R942 VTAIL.n143 VTAIL.n99 0.155672
R943 VTAIL.n144 VTAIL.n143 0.155672
R944 VTAIL.n144 VTAIL.n95 0.155672
R945 VTAIL.n151 VTAIL.n95 0.155672
R946 VTAIL.n152 VTAIL.n151 0.155672
R947 VTAIL.n152 VTAIL.n91 0.155672
R948 VTAIL.n161 VTAIL.n91 0.155672
R949 VTAIL.n162 VTAIL.n161 0.155672
R950 VTAIL.n162 VTAIL.n87 0.155672
R951 VTAIL.n169 VTAIL.n87 0.155672
R952 VTAIL.n205 VTAIL.n197 0.155672
R953 VTAIL.n206 VTAIL.n205 0.155672
R954 VTAIL.n206 VTAIL.n193 0.155672
R955 VTAIL.n213 VTAIL.n193 0.155672
R956 VTAIL.n214 VTAIL.n213 0.155672
R957 VTAIL.n214 VTAIL.n189 0.155672
R958 VTAIL.n221 VTAIL.n189 0.155672
R959 VTAIL.n222 VTAIL.n221 0.155672
R960 VTAIL.n222 VTAIL.n185 0.155672
R961 VTAIL.n229 VTAIL.n185 0.155672
R962 VTAIL.n230 VTAIL.n229 0.155672
R963 VTAIL.n230 VTAIL.n181 0.155672
R964 VTAIL.n237 VTAIL.n181 0.155672
R965 VTAIL.n238 VTAIL.n237 0.155672
R966 VTAIL.n238 VTAIL.n177 0.155672
R967 VTAIL.n247 VTAIL.n177 0.155672
R968 VTAIL.n248 VTAIL.n247 0.155672
R969 VTAIL.n248 VTAIL.n173 0.155672
R970 VTAIL.n255 VTAIL.n173 0.155672
R971 VTAIL.n599 VTAIL.n517 0.155672
R972 VTAIL.n592 VTAIL.n517 0.155672
R973 VTAIL.n592 VTAIL.n591 0.155672
R974 VTAIL.n591 VTAIL.n521 0.155672
R975 VTAIL.n584 VTAIL.n521 0.155672
R976 VTAIL.n584 VTAIL.n583 0.155672
R977 VTAIL.n583 VTAIL.n527 0.155672
R978 VTAIL.n576 VTAIL.n527 0.155672
R979 VTAIL.n576 VTAIL.n575 0.155672
R980 VTAIL.n575 VTAIL.n531 0.155672
R981 VTAIL.n568 VTAIL.n531 0.155672
R982 VTAIL.n568 VTAIL.n567 0.155672
R983 VTAIL.n567 VTAIL.n535 0.155672
R984 VTAIL.n560 VTAIL.n535 0.155672
R985 VTAIL.n560 VTAIL.n559 0.155672
R986 VTAIL.n559 VTAIL.n539 0.155672
R987 VTAIL.n552 VTAIL.n539 0.155672
R988 VTAIL.n552 VTAIL.n551 0.155672
R989 VTAIL.n551 VTAIL.n543 0.155672
R990 VTAIL.n513 VTAIL.n431 0.155672
R991 VTAIL.n506 VTAIL.n431 0.155672
R992 VTAIL.n506 VTAIL.n505 0.155672
R993 VTAIL.n505 VTAIL.n435 0.155672
R994 VTAIL.n498 VTAIL.n435 0.155672
R995 VTAIL.n498 VTAIL.n497 0.155672
R996 VTAIL.n497 VTAIL.n441 0.155672
R997 VTAIL.n490 VTAIL.n441 0.155672
R998 VTAIL.n490 VTAIL.n489 0.155672
R999 VTAIL.n489 VTAIL.n445 0.155672
R1000 VTAIL.n482 VTAIL.n445 0.155672
R1001 VTAIL.n482 VTAIL.n481 0.155672
R1002 VTAIL.n481 VTAIL.n449 0.155672
R1003 VTAIL.n474 VTAIL.n449 0.155672
R1004 VTAIL.n474 VTAIL.n473 0.155672
R1005 VTAIL.n473 VTAIL.n453 0.155672
R1006 VTAIL.n466 VTAIL.n453 0.155672
R1007 VTAIL.n466 VTAIL.n465 0.155672
R1008 VTAIL.n465 VTAIL.n457 0.155672
R1009 VTAIL.n427 VTAIL.n345 0.155672
R1010 VTAIL.n420 VTAIL.n345 0.155672
R1011 VTAIL.n420 VTAIL.n419 0.155672
R1012 VTAIL.n419 VTAIL.n349 0.155672
R1013 VTAIL.n412 VTAIL.n349 0.155672
R1014 VTAIL.n412 VTAIL.n411 0.155672
R1015 VTAIL.n411 VTAIL.n355 0.155672
R1016 VTAIL.n404 VTAIL.n355 0.155672
R1017 VTAIL.n404 VTAIL.n403 0.155672
R1018 VTAIL.n403 VTAIL.n359 0.155672
R1019 VTAIL.n396 VTAIL.n359 0.155672
R1020 VTAIL.n396 VTAIL.n395 0.155672
R1021 VTAIL.n395 VTAIL.n363 0.155672
R1022 VTAIL.n388 VTAIL.n363 0.155672
R1023 VTAIL.n388 VTAIL.n387 0.155672
R1024 VTAIL.n387 VTAIL.n367 0.155672
R1025 VTAIL.n380 VTAIL.n367 0.155672
R1026 VTAIL.n380 VTAIL.n379 0.155672
R1027 VTAIL.n379 VTAIL.n371 0.155672
R1028 VTAIL.n341 VTAIL.n259 0.155672
R1029 VTAIL.n334 VTAIL.n259 0.155672
R1030 VTAIL.n334 VTAIL.n333 0.155672
R1031 VTAIL.n333 VTAIL.n263 0.155672
R1032 VTAIL.n326 VTAIL.n263 0.155672
R1033 VTAIL.n326 VTAIL.n325 0.155672
R1034 VTAIL.n325 VTAIL.n269 0.155672
R1035 VTAIL.n318 VTAIL.n269 0.155672
R1036 VTAIL.n318 VTAIL.n317 0.155672
R1037 VTAIL.n317 VTAIL.n273 0.155672
R1038 VTAIL.n310 VTAIL.n273 0.155672
R1039 VTAIL.n310 VTAIL.n309 0.155672
R1040 VTAIL.n309 VTAIL.n277 0.155672
R1041 VTAIL.n302 VTAIL.n277 0.155672
R1042 VTAIL.n302 VTAIL.n301 0.155672
R1043 VTAIL.n301 VTAIL.n281 0.155672
R1044 VTAIL.n294 VTAIL.n281 0.155672
R1045 VTAIL.n294 VTAIL.n293 0.155672
R1046 VTAIL.n293 VTAIL.n285 0.155672
R1047 VDD2.n2 VDD2.n0 99.8804
R1048 VDD2.n2 VDD2.n1 61.0363
R1049 VDD2.n1 VDD2.t1 1.28872
R1050 VDD2.n1 VDD2.t3 1.28872
R1051 VDD2.n0 VDD2.t2 1.28872
R1052 VDD2.n0 VDD2.t0 1.28872
R1053 VDD2 VDD2.n2 0.0586897
R1054 B.n58 B.t15 1159.59
R1055 B.n64 B.t4 1159.59
R1056 B.n151 B.t12 1159.59
R1057 B.n145 B.t8 1159.59
R1058 B.n468 B.n91 585
R1059 B.n91 B.n30 585
R1060 B.n470 B.n469 585
R1061 B.n472 B.n90 585
R1062 B.n475 B.n474 585
R1063 B.n476 B.n89 585
R1064 B.n478 B.n477 585
R1065 B.n480 B.n88 585
R1066 B.n483 B.n482 585
R1067 B.n484 B.n87 585
R1068 B.n486 B.n485 585
R1069 B.n488 B.n86 585
R1070 B.n491 B.n490 585
R1071 B.n492 B.n85 585
R1072 B.n494 B.n493 585
R1073 B.n496 B.n84 585
R1074 B.n499 B.n498 585
R1075 B.n500 B.n83 585
R1076 B.n502 B.n501 585
R1077 B.n504 B.n82 585
R1078 B.n507 B.n506 585
R1079 B.n508 B.n81 585
R1080 B.n510 B.n509 585
R1081 B.n512 B.n80 585
R1082 B.n515 B.n514 585
R1083 B.n516 B.n79 585
R1084 B.n518 B.n517 585
R1085 B.n520 B.n78 585
R1086 B.n523 B.n522 585
R1087 B.n524 B.n77 585
R1088 B.n526 B.n525 585
R1089 B.n528 B.n76 585
R1090 B.n531 B.n530 585
R1091 B.n532 B.n75 585
R1092 B.n534 B.n533 585
R1093 B.n536 B.n74 585
R1094 B.n539 B.n538 585
R1095 B.n540 B.n73 585
R1096 B.n542 B.n541 585
R1097 B.n544 B.n72 585
R1098 B.n547 B.n546 585
R1099 B.n548 B.n71 585
R1100 B.n550 B.n549 585
R1101 B.n552 B.n70 585
R1102 B.n555 B.n554 585
R1103 B.n556 B.n69 585
R1104 B.n558 B.n557 585
R1105 B.n560 B.n68 585
R1106 B.n563 B.n562 585
R1107 B.n564 B.n67 585
R1108 B.n566 B.n565 585
R1109 B.n568 B.n66 585
R1110 B.n571 B.n570 585
R1111 B.n573 B.n63 585
R1112 B.n575 B.n574 585
R1113 B.n577 B.n62 585
R1114 B.n580 B.n579 585
R1115 B.n581 B.n61 585
R1116 B.n583 B.n582 585
R1117 B.n585 B.n60 585
R1118 B.n588 B.n587 585
R1119 B.n589 B.n57 585
R1120 B.n592 B.n591 585
R1121 B.n594 B.n56 585
R1122 B.n597 B.n596 585
R1123 B.n598 B.n55 585
R1124 B.n600 B.n599 585
R1125 B.n602 B.n54 585
R1126 B.n605 B.n604 585
R1127 B.n606 B.n53 585
R1128 B.n608 B.n607 585
R1129 B.n610 B.n52 585
R1130 B.n613 B.n612 585
R1131 B.n614 B.n51 585
R1132 B.n616 B.n615 585
R1133 B.n618 B.n50 585
R1134 B.n621 B.n620 585
R1135 B.n622 B.n49 585
R1136 B.n624 B.n623 585
R1137 B.n626 B.n48 585
R1138 B.n629 B.n628 585
R1139 B.n630 B.n47 585
R1140 B.n632 B.n631 585
R1141 B.n634 B.n46 585
R1142 B.n637 B.n636 585
R1143 B.n638 B.n45 585
R1144 B.n640 B.n639 585
R1145 B.n642 B.n44 585
R1146 B.n645 B.n644 585
R1147 B.n646 B.n43 585
R1148 B.n648 B.n647 585
R1149 B.n650 B.n42 585
R1150 B.n653 B.n652 585
R1151 B.n654 B.n41 585
R1152 B.n656 B.n655 585
R1153 B.n658 B.n40 585
R1154 B.n661 B.n660 585
R1155 B.n662 B.n39 585
R1156 B.n664 B.n663 585
R1157 B.n666 B.n38 585
R1158 B.n669 B.n668 585
R1159 B.n670 B.n37 585
R1160 B.n672 B.n671 585
R1161 B.n674 B.n36 585
R1162 B.n677 B.n676 585
R1163 B.n678 B.n35 585
R1164 B.n680 B.n679 585
R1165 B.n682 B.n34 585
R1166 B.n685 B.n684 585
R1167 B.n686 B.n33 585
R1168 B.n688 B.n687 585
R1169 B.n690 B.n32 585
R1170 B.n693 B.n692 585
R1171 B.n694 B.n31 585
R1172 B.n467 B.n29 585
R1173 B.n697 B.n29 585
R1174 B.n466 B.n28 585
R1175 B.n698 B.n28 585
R1176 B.n465 B.n27 585
R1177 B.n699 B.n27 585
R1178 B.n464 B.n463 585
R1179 B.n463 B.n23 585
R1180 B.n462 B.n22 585
R1181 B.n705 B.n22 585
R1182 B.n461 B.n21 585
R1183 B.n706 B.n21 585
R1184 B.n460 B.n20 585
R1185 B.n707 B.n20 585
R1186 B.n459 B.n458 585
R1187 B.n458 B.n16 585
R1188 B.n457 B.n15 585
R1189 B.n713 B.n15 585
R1190 B.n456 B.n14 585
R1191 B.n714 B.n14 585
R1192 B.n455 B.n13 585
R1193 B.n715 B.n13 585
R1194 B.n454 B.n453 585
R1195 B.n453 B.n12 585
R1196 B.n452 B.n451 585
R1197 B.n452 B.n8 585
R1198 B.n450 B.n7 585
R1199 B.n722 B.n7 585
R1200 B.n449 B.n6 585
R1201 B.n723 B.n6 585
R1202 B.n448 B.n5 585
R1203 B.n724 B.n5 585
R1204 B.n447 B.n446 585
R1205 B.n446 B.n4 585
R1206 B.n445 B.n92 585
R1207 B.n445 B.n444 585
R1208 B.n434 B.n93 585
R1209 B.n437 B.n93 585
R1210 B.n436 B.n435 585
R1211 B.n438 B.n436 585
R1212 B.n433 B.n97 585
R1213 B.n101 B.n97 585
R1214 B.n432 B.n431 585
R1215 B.n431 B.n430 585
R1216 B.n99 B.n98 585
R1217 B.n100 B.n99 585
R1218 B.n423 B.n422 585
R1219 B.n424 B.n423 585
R1220 B.n421 B.n106 585
R1221 B.n106 B.n105 585
R1222 B.n420 B.n419 585
R1223 B.n419 B.n418 585
R1224 B.n108 B.n107 585
R1225 B.n109 B.n108 585
R1226 B.n411 B.n410 585
R1227 B.n412 B.n411 585
R1228 B.n409 B.n114 585
R1229 B.n114 B.n113 585
R1230 B.n408 B.n407 585
R1231 B.n407 B.n406 585
R1232 B.n403 B.n118 585
R1233 B.n402 B.n401 585
R1234 B.n399 B.n119 585
R1235 B.n399 B.n117 585
R1236 B.n398 B.n397 585
R1237 B.n396 B.n395 585
R1238 B.n394 B.n121 585
R1239 B.n392 B.n391 585
R1240 B.n390 B.n122 585
R1241 B.n389 B.n388 585
R1242 B.n386 B.n123 585
R1243 B.n384 B.n383 585
R1244 B.n382 B.n124 585
R1245 B.n381 B.n380 585
R1246 B.n378 B.n125 585
R1247 B.n376 B.n375 585
R1248 B.n374 B.n126 585
R1249 B.n373 B.n372 585
R1250 B.n370 B.n127 585
R1251 B.n368 B.n367 585
R1252 B.n366 B.n128 585
R1253 B.n365 B.n364 585
R1254 B.n362 B.n129 585
R1255 B.n360 B.n359 585
R1256 B.n358 B.n130 585
R1257 B.n357 B.n356 585
R1258 B.n354 B.n131 585
R1259 B.n352 B.n351 585
R1260 B.n350 B.n132 585
R1261 B.n349 B.n348 585
R1262 B.n346 B.n133 585
R1263 B.n344 B.n343 585
R1264 B.n342 B.n134 585
R1265 B.n341 B.n340 585
R1266 B.n338 B.n135 585
R1267 B.n336 B.n335 585
R1268 B.n334 B.n136 585
R1269 B.n333 B.n332 585
R1270 B.n330 B.n137 585
R1271 B.n328 B.n327 585
R1272 B.n326 B.n138 585
R1273 B.n325 B.n324 585
R1274 B.n322 B.n139 585
R1275 B.n320 B.n319 585
R1276 B.n318 B.n140 585
R1277 B.n317 B.n316 585
R1278 B.n314 B.n141 585
R1279 B.n312 B.n311 585
R1280 B.n310 B.n142 585
R1281 B.n309 B.n308 585
R1282 B.n306 B.n143 585
R1283 B.n304 B.n303 585
R1284 B.n302 B.n144 585
R1285 B.n300 B.n299 585
R1286 B.n297 B.n147 585
R1287 B.n295 B.n294 585
R1288 B.n293 B.n148 585
R1289 B.n292 B.n291 585
R1290 B.n289 B.n149 585
R1291 B.n287 B.n286 585
R1292 B.n285 B.n150 585
R1293 B.n284 B.n283 585
R1294 B.n281 B.n280 585
R1295 B.n279 B.n278 585
R1296 B.n277 B.n155 585
R1297 B.n275 B.n274 585
R1298 B.n273 B.n156 585
R1299 B.n272 B.n271 585
R1300 B.n269 B.n157 585
R1301 B.n267 B.n266 585
R1302 B.n265 B.n158 585
R1303 B.n264 B.n263 585
R1304 B.n261 B.n159 585
R1305 B.n259 B.n258 585
R1306 B.n257 B.n160 585
R1307 B.n256 B.n255 585
R1308 B.n253 B.n161 585
R1309 B.n251 B.n250 585
R1310 B.n249 B.n162 585
R1311 B.n248 B.n247 585
R1312 B.n245 B.n163 585
R1313 B.n243 B.n242 585
R1314 B.n241 B.n164 585
R1315 B.n240 B.n239 585
R1316 B.n237 B.n165 585
R1317 B.n235 B.n234 585
R1318 B.n233 B.n166 585
R1319 B.n232 B.n231 585
R1320 B.n229 B.n167 585
R1321 B.n227 B.n226 585
R1322 B.n225 B.n168 585
R1323 B.n224 B.n223 585
R1324 B.n221 B.n169 585
R1325 B.n219 B.n218 585
R1326 B.n217 B.n170 585
R1327 B.n216 B.n215 585
R1328 B.n213 B.n171 585
R1329 B.n211 B.n210 585
R1330 B.n209 B.n172 585
R1331 B.n208 B.n207 585
R1332 B.n205 B.n173 585
R1333 B.n203 B.n202 585
R1334 B.n201 B.n174 585
R1335 B.n200 B.n199 585
R1336 B.n197 B.n175 585
R1337 B.n195 B.n194 585
R1338 B.n193 B.n176 585
R1339 B.n192 B.n191 585
R1340 B.n189 B.n177 585
R1341 B.n187 B.n186 585
R1342 B.n185 B.n178 585
R1343 B.n184 B.n183 585
R1344 B.n181 B.n179 585
R1345 B.n116 B.n115 585
R1346 B.n405 B.n404 585
R1347 B.n406 B.n405 585
R1348 B.n112 B.n111 585
R1349 B.n113 B.n112 585
R1350 B.n414 B.n413 585
R1351 B.n413 B.n412 585
R1352 B.n415 B.n110 585
R1353 B.n110 B.n109 585
R1354 B.n417 B.n416 585
R1355 B.n418 B.n417 585
R1356 B.n104 B.n103 585
R1357 B.n105 B.n104 585
R1358 B.n426 B.n425 585
R1359 B.n425 B.n424 585
R1360 B.n427 B.n102 585
R1361 B.n102 B.n100 585
R1362 B.n429 B.n428 585
R1363 B.n430 B.n429 585
R1364 B.n96 B.n95 585
R1365 B.n101 B.n96 585
R1366 B.n440 B.n439 585
R1367 B.n439 B.n438 585
R1368 B.n441 B.n94 585
R1369 B.n437 B.n94 585
R1370 B.n443 B.n442 585
R1371 B.n444 B.n443 585
R1372 B.n3 B.n0 585
R1373 B.n4 B.n3 585
R1374 B.n721 B.n1 585
R1375 B.n722 B.n721 585
R1376 B.n720 B.n719 585
R1377 B.n720 B.n8 585
R1378 B.n718 B.n9 585
R1379 B.n12 B.n9 585
R1380 B.n717 B.n716 585
R1381 B.n716 B.n715 585
R1382 B.n11 B.n10 585
R1383 B.n714 B.n11 585
R1384 B.n712 B.n711 585
R1385 B.n713 B.n712 585
R1386 B.n710 B.n17 585
R1387 B.n17 B.n16 585
R1388 B.n709 B.n708 585
R1389 B.n708 B.n707 585
R1390 B.n19 B.n18 585
R1391 B.n706 B.n19 585
R1392 B.n704 B.n703 585
R1393 B.n705 B.n704 585
R1394 B.n702 B.n24 585
R1395 B.n24 B.n23 585
R1396 B.n701 B.n700 585
R1397 B.n700 B.n699 585
R1398 B.n26 B.n25 585
R1399 B.n698 B.n26 585
R1400 B.n696 B.n695 585
R1401 B.n697 B.n696 585
R1402 B.n725 B.n724 585
R1403 B.n723 B.n2 585
R1404 B.n696 B.n31 473.281
R1405 B.n91 B.n29 473.281
R1406 B.n407 B.n116 473.281
R1407 B.n405 B.n118 473.281
R1408 B.n64 B.t6 353.952
R1409 B.n151 B.t14 353.952
R1410 B.n58 B.t16 353.952
R1411 B.n145 B.t11 353.952
R1412 B.n65 B.t7 339.988
R1413 B.n152 B.t13 339.988
R1414 B.n59 B.t17 339.988
R1415 B.n146 B.t10 339.988
R1416 B.n471 B.n30 256.663
R1417 B.n473 B.n30 256.663
R1418 B.n479 B.n30 256.663
R1419 B.n481 B.n30 256.663
R1420 B.n487 B.n30 256.663
R1421 B.n489 B.n30 256.663
R1422 B.n495 B.n30 256.663
R1423 B.n497 B.n30 256.663
R1424 B.n503 B.n30 256.663
R1425 B.n505 B.n30 256.663
R1426 B.n511 B.n30 256.663
R1427 B.n513 B.n30 256.663
R1428 B.n519 B.n30 256.663
R1429 B.n521 B.n30 256.663
R1430 B.n527 B.n30 256.663
R1431 B.n529 B.n30 256.663
R1432 B.n535 B.n30 256.663
R1433 B.n537 B.n30 256.663
R1434 B.n543 B.n30 256.663
R1435 B.n545 B.n30 256.663
R1436 B.n551 B.n30 256.663
R1437 B.n553 B.n30 256.663
R1438 B.n559 B.n30 256.663
R1439 B.n561 B.n30 256.663
R1440 B.n567 B.n30 256.663
R1441 B.n569 B.n30 256.663
R1442 B.n576 B.n30 256.663
R1443 B.n578 B.n30 256.663
R1444 B.n584 B.n30 256.663
R1445 B.n586 B.n30 256.663
R1446 B.n593 B.n30 256.663
R1447 B.n595 B.n30 256.663
R1448 B.n601 B.n30 256.663
R1449 B.n603 B.n30 256.663
R1450 B.n609 B.n30 256.663
R1451 B.n611 B.n30 256.663
R1452 B.n617 B.n30 256.663
R1453 B.n619 B.n30 256.663
R1454 B.n625 B.n30 256.663
R1455 B.n627 B.n30 256.663
R1456 B.n633 B.n30 256.663
R1457 B.n635 B.n30 256.663
R1458 B.n641 B.n30 256.663
R1459 B.n643 B.n30 256.663
R1460 B.n649 B.n30 256.663
R1461 B.n651 B.n30 256.663
R1462 B.n657 B.n30 256.663
R1463 B.n659 B.n30 256.663
R1464 B.n665 B.n30 256.663
R1465 B.n667 B.n30 256.663
R1466 B.n673 B.n30 256.663
R1467 B.n675 B.n30 256.663
R1468 B.n681 B.n30 256.663
R1469 B.n683 B.n30 256.663
R1470 B.n689 B.n30 256.663
R1471 B.n691 B.n30 256.663
R1472 B.n400 B.n117 256.663
R1473 B.n120 B.n117 256.663
R1474 B.n393 B.n117 256.663
R1475 B.n387 B.n117 256.663
R1476 B.n385 B.n117 256.663
R1477 B.n379 B.n117 256.663
R1478 B.n377 B.n117 256.663
R1479 B.n371 B.n117 256.663
R1480 B.n369 B.n117 256.663
R1481 B.n363 B.n117 256.663
R1482 B.n361 B.n117 256.663
R1483 B.n355 B.n117 256.663
R1484 B.n353 B.n117 256.663
R1485 B.n347 B.n117 256.663
R1486 B.n345 B.n117 256.663
R1487 B.n339 B.n117 256.663
R1488 B.n337 B.n117 256.663
R1489 B.n331 B.n117 256.663
R1490 B.n329 B.n117 256.663
R1491 B.n323 B.n117 256.663
R1492 B.n321 B.n117 256.663
R1493 B.n315 B.n117 256.663
R1494 B.n313 B.n117 256.663
R1495 B.n307 B.n117 256.663
R1496 B.n305 B.n117 256.663
R1497 B.n298 B.n117 256.663
R1498 B.n296 B.n117 256.663
R1499 B.n290 B.n117 256.663
R1500 B.n288 B.n117 256.663
R1501 B.n282 B.n117 256.663
R1502 B.n154 B.n117 256.663
R1503 B.n276 B.n117 256.663
R1504 B.n270 B.n117 256.663
R1505 B.n268 B.n117 256.663
R1506 B.n262 B.n117 256.663
R1507 B.n260 B.n117 256.663
R1508 B.n254 B.n117 256.663
R1509 B.n252 B.n117 256.663
R1510 B.n246 B.n117 256.663
R1511 B.n244 B.n117 256.663
R1512 B.n238 B.n117 256.663
R1513 B.n236 B.n117 256.663
R1514 B.n230 B.n117 256.663
R1515 B.n228 B.n117 256.663
R1516 B.n222 B.n117 256.663
R1517 B.n220 B.n117 256.663
R1518 B.n214 B.n117 256.663
R1519 B.n212 B.n117 256.663
R1520 B.n206 B.n117 256.663
R1521 B.n204 B.n117 256.663
R1522 B.n198 B.n117 256.663
R1523 B.n196 B.n117 256.663
R1524 B.n190 B.n117 256.663
R1525 B.n188 B.n117 256.663
R1526 B.n182 B.n117 256.663
R1527 B.n180 B.n117 256.663
R1528 B.n727 B.n726 256.663
R1529 B.n692 B.n690 163.367
R1530 B.n688 B.n33 163.367
R1531 B.n684 B.n682 163.367
R1532 B.n680 B.n35 163.367
R1533 B.n676 B.n674 163.367
R1534 B.n672 B.n37 163.367
R1535 B.n668 B.n666 163.367
R1536 B.n664 B.n39 163.367
R1537 B.n660 B.n658 163.367
R1538 B.n656 B.n41 163.367
R1539 B.n652 B.n650 163.367
R1540 B.n648 B.n43 163.367
R1541 B.n644 B.n642 163.367
R1542 B.n640 B.n45 163.367
R1543 B.n636 B.n634 163.367
R1544 B.n632 B.n47 163.367
R1545 B.n628 B.n626 163.367
R1546 B.n624 B.n49 163.367
R1547 B.n620 B.n618 163.367
R1548 B.n616 B.n51 163.367
R1549 B.n612 B.n610 163.367
R1550 B.n608 B.n53 163.367
R1551 B.n604 B.n602 163.367
R1552 B.n600 B.n55 163.367
R1553 B.n596 B.n594 163.367
R1554 B.n592 B.n57 163.367
R1555 B.n587 B.n585 163.367
R1556 B.n583 B.n61 163.367
R1557 B.n579 B.n577 163.367
R1558 B.n575 B.n63 163.367
R1559 B.n570 B.n568 163.367
R1560 B.n566 B.n67 163.367
R1561 B.n562 B.n560 163.367
R1562 B.n558 B.n69 163.367
R1563 B.n554 B.n552 163.367
R1564 B.n550 B.n71 163.367
R1565 B.n546 B.n544 163.367
R1566 B.n542 B.n73 163.367
R1567 B.n538 B.n536 163.367
R1568 B.n534 B.n75 163.367
R1569 B.n530 B.n528 163.367
R1570 B.n526 B.n77 163.367
R1571 B.n522 B.n520 163.367
R1572 B.n518 B.n79 163.367
R1573 B.n514 B.n512 163.367
R1574 B.n510 B.n81 163.367
R1575 B.n506 B.n504 163.367
R1576 B.n502 B.n83 163.367
R1577 B.n498 B.n496 163.367
R1578 B.n494 B.n85 163.367
R1579 B.n490 B.n488 163.367
R1580 B.n486 B.n87 163.367
R1581 B.n482 B.n480 163.367
R1582 B.n478 B.n89 163.367
R1583 B.n474 B.n472 163.367
R1584 B.n470 B.n91 163.367
R1585 B.n407 B.n114 163.367
R1586 B.n411 B.n114 163.367
R1587 B.n411 B.n108 163.367
R1588 B.n419 B.n108 163.367
R1589 B.n419 B.n106 163.367
R1590 B.n423 B.n106 163.367
R1591 B.n423 B.n99 163.367
R1592 B.n431 B.n99 163.367
R1593 B.n431 B.n97 163.367
R1594 B.n436 B.n97 163.367
R1595 B.n436 B.n93 163.367
R1596 B.n445 B.n93 163.367
R1597 B.n446 B.n445 163.367
R1598 B.n446 B.n5 163.367
R1599 B.n6 B.n5 163.367
R1600 B.n7 B.n6 163.367
R1601 B.n452 B.n7 163.367
R1602 B.n453 B.n452 163.367
R1603 B.n453 B.n13 163.367
R1604 B.n14 B.n13 163.367
R1605 B.n15 B.n14 163.367
R1606 B.n458 B.n15 163.367
R1607 B.n458 B.n20 163.367
R1608 B.n21 B.n20 163.367
R1609 B.n22 B.n21 163.367
R1610 B.n463 B.n22 163.367
R1611 B.n463 B.n27 163.367
R1612 B.n28 B.n27 163.367
R1613 B.n29 B.n28 163.367
R1614 B.n401 B.n399 163.367
R1615 B.n399 B.n398 163.367
R1616 B.n395 B.n394 163.367
R1617 B.n392 B.n122 163.367
R1618 B.n388 B.n386 163.367
R1619 B.n384 B.n124 163.367
R1620 B.n380 B.n378 163.367
R1621 B.n376 B.n126 163.367
R1622 B.n372 B.n370 163.367
R1623 B.n368 B.n128 163.367
R1624 B.n364 B.n362 163.367
R1625 B.n360 B.n130 163.367
R1626 B.n356 B.n354 163.367
R1627 B.n352 B.n132 163.367
R1628 B.n348 B.n346 163.367
R1629 B.n344 B.n134 163.367
R1630 B.n340 B.n338 163.367
R1631 B.n336 B.n136 163.367
R1632 B.n332 B.n330 163.367
R1633 B.n328 B.n138 163.367
R1634 B.n324 B.n322 163.367
R1635 B.n320 B.n140 163.367
R1636 B.n316 B.n314 163.367
R1637 B.n312 B.n142 163.367
R1638 B.n308 B.n306 163.367
R1639 B.n304 B.n144 163.367
R1640 B.n299 B.n297 163.367
R1641 B.n295 B.n148 163.367
R1642 B.n291 B.n289 163.367
R1643 B.n287 B.n150 163.367
R1644 B.n283 B.n281 163.367
R1645 B.n278 B.n277 163.367
R1646 B.n275 B.n156 163.367
R1647 B.n271 B.n269 163.367
R1648 B.n267 B.n158 163.367
R1649 B.n263 B.n261 163.367
R1650 B.n259 B.n160 163.367
R1651 B.n255 B.n253 163.367
R1652 B.n251 B.n162 163.367
R1653 B.n247 B.n245 163.367
R1654 B.n243 B.n164 163.367
R1655 B.n239 B.n237 163.367
R1656 B.n235 B.n166 163.367
R1657 B.n231 B.n229 163.367
R1658 B.n227 B.n168 163.367
R1659 B.n223 B.n221 163.367
R1660 B.n219 B.n170 163.367
R1661 B.n215 B.n213 163.367
R1662 B.n211 B.n172 163.367
R1663 B.n207 B.n205 163.367
R1664 B.n203 B.n174 163.367
R1665 B.n199 B.n197 163.367
R1666 B.n195 B.n176 163.367
R1667 B.n191 B.n189 163.367
R1668 B.n187 B.n178 163.367
R1669 B.n183 B.n181 163.367
R1670 B.n405 B.n112 163.367
R1671 B.n413 B.n112 163.367
R1672 B.n413 B.n110 163.367
R1673 B.n417 B.n110 163.367
R1674 B.n417 B.n104 163.367
R1675 B.n425 B.n104 163.367
R1676 B.n425 B.n102 163.367
R1677 B.n429 B.n102 163.367
R1678 B.n429 B.n96 163.367
R1679 B.n439 B.n96 163.367
R1680 B.n439 B.n94 163.367
R1681 B.n443 B.n94 163.367
R1682 B.n443 B.n3 163.367
R1683 B.n725 B.n3 163.367
R1684 B.n721 B.n2 163.367
R1685 B.n721 B.n720 163.367
R1686 B.n720 B.n9 163.367
R1687 B.n716 B.n9 163.367
R1688 B.n716 B.n11 163.367
R1689 B.n712 B.n11 163.367
R1690 B.n712 B.n17 163.367
R1691 B.n708 B.n17 163.367
R1692 B.n708 B.n19 163.367
R1693 B.n704 B.n19 163.367
R1694 B.n704 B.n24 163.367
R1695 B.n700 B.n24 163.367
R1696 B.n700 B.n26 163.367
R1697 B.n696 B.n26 163.367
R1698 B.n691 B.n31 71.676
R1699 B.n690 B.n689 71.676
R1700 B.n683 B.n33 71.676
R1701 B.n682 B.n681 71.676
R1702 B.n675 B.n35 71.676
R1703 B.n674 B.n673 71.676
R1704 B.n667 B.n37 71.676
R1705 B.n666 B.n665 71.676
R1706 B.n659 B.n39 71.676
R1707 B.n658 B.n657 71.676
R1708 B.n651 B.n41 71.676
R1709 B.n650 B.n649 71.676
R1710 B.n643 B.n43 71.676
R1711 B.n642 B.n641 71.676
R1712 B.n635 B.n45 71.676
R1713 B.n634 B.n633 71.676
R1714 B.n627 B.n47 71.676
R1715 B.n626 B.n625 71.676
R1716 B.n619 B.n49 71.676
R1717 B.n618 B.n617 71.676
R1718 B.n611 B.n51 71.676
R1719 B.n610 B.n609 71.676
R1720 B.n603 B.n53 71.676
R1721 B.n602 B.n601 71.676
R1722 B.n595 B.n55 71.676
R1723 B.n594 B.n593 71.676
R1724 B.n586 B.n57 71.676
R1725 B.n585 B.n584 71.676
R1726 B.n578 B.n61 71.676
R1727 B.n577 B.n576 71.676
R1728 B.n569 B.n63 71.676
R1729 B.n568 B.n567 71.676
R1730 B.n561 B.n67 71.676
R1731 B.n560 B.n559 71.676
R1732 B.n553 B.n69 71.676
R1733 B.n552 B.n551 71.676
R1734 B.n545 B.n71 71.676
R1735 B.n544 B.n543 71.676
R1736 B.n537 B.n73 71.676
R1737 B.n536 B.n535 71.676
R1738 B.n529 B.n75 71.676
R1739 B.n528 B.n527 71.676
R1740 B.n521 B.n77 71.676
R1741 B.n520 B.n519 71.676
R1742 B.n513 B.n79 71.676
R1743 B.n512 B.n511 71.676
R1744 B.n505 B.n81 71.676
R1745 B.n504 B.n503 71.676
R1746 B.n497 B.n83 71.676
R1747 B.n496 B.n495 71.676
R1748 B.n489 B.n85 71.676
R1749 B.n488 B.n487 71.676
R1750 B.n481 B.n87 71.676
R1751 B.n480 B.n479 71.676
R1752 B.n473 B.n89 71.676
R1753 B.n472 B.n471 71.676
R1754 B.n471 B.n470 71.676
R1755 B.n474 B.n473 71.676
R1756 B.n479 B.n478 71.676
R1757 B.n482 B.n481 71.676
R1758 B.n487 B.n486 71.676
R1759 B.n490 B.n489 71.676
R1760 B.n495 B.n494 71.676
R1761 B.n498 B.n497 71.676
R1762 B.n503 B.n502 71.676
R1763 B.n506 B.n505 71.676
R1764 B.n511 B.n510 71.676
R1765 B.n514 B.n513 71.676
R1766 B.n519 B.n518 71.676
R1767 B.n522 B.n521 71.676
R1768 B.n527 B.n526 71.676
R1769 B.n530 B.n529 71.676
R1770 B.n535 B.n534 71.676
R1771 B.n538 B.n537 71.676
R1772 B.n543 B.n542 71.676
R1773 B.n546 B.n545 71.676
R1774 B.n551 B.n550 71.676
R1775 B.n554 B.n553 71.676
R1776 B.n559 B.n558 71.676
R1777 B.n562 B.n561 71.676
R1778 B.n567 B.n566 71.676
R1779 B.n570 B.n569 71.676
R1780 B.n576 B.n575 71.676
R1781 B.n579 B.n578 71.676
R1782 B.n584 B.n583 71.676
R1783 B.n587 B.n586 71.676
R1784 B.n593 B.n592 71.676
R1785 B.n596 B.n595 71.676
R1786 B.n601 B.n600 71.676
R1787 B.n604 B.n603 71.676
R1788 B.n609 B.n608 71.676
R1789 B.n612 B.n611 71.676
R1790 B.n617 B.n616 71.676
R1791 B.n620 B.n619 71.676
R1792 B.n625 B.n624 71.676
R1793 B.n628 B.n627 71.676
R1794 B.n633 B.n632 71.676
R1795 B.n636 B.n635 71.676
R1796 B.n641 B.n640 71.676
R1797 B.n644 B.n643 71.676
R1798 B.n649 B.n648 71.676
R1799 B.n652 B.n651 71.676
R1800 B.n657 B.n656 71.676
R1801 B.n660 B.n659 71.676
R1802 B.n665 B.n664 71.676
R1803 B.n668 B.n667 71.676
R1804 B.n673 B.n672 71.676
R1805 B.n676 B.n675 71.676
R1806 B.n681 B.n680 71.676
R1807 B.n684 B.n683 71.676
R1808 B.n689 B.n688 71.676
R1809 B.n692 B.n691 71.676
R1810 B.n400 B.n118 71.676
R1811 B.n398 B.n120 71.676
R1812 B.n394 B.n393 71.676
R1813 B.n387 B.n122 71.676
R1814 B.n386 B.n385 71.676
R1815 B.n379 B.n124 71.676
R1816 B.n378 B.n377 71.676
R1817 B.n371 B.n126 71.676
R1818 B.n370 B.n369 71.676
R1819 B.n363 B.n128 71.676
R1820 B.n362 B.n361 71.676
R1821 B.n355 B.n130 71.676
R1822 B.n354 B.n353 71.676
R1823 B.n347 B.n132 71.676
R1824 B.n346 B.n345 71.676
R1825 B.n339 B.n134 71.676
R1826 B.n338 B.n337 71.676
R1827 B.n331 B.n136 71.676
R1828 B.n330 B.n329 71.676
R1829 B.n323 B.n138 71.676
R1830 B.n322 B.n321 71.676
R1831 B.n315 B.n140 71.676
R1832 B.n314 B.n313 71.676
R1833 B.n307 B.n142 71.676
R1834 B.n306 B.n305 71.676
R1835 B.n298 B.n144 71.676
R1836 B.n297 B.n296 71.676
R1837 B.n290 B.n148 71.676
R1838 B.n289 B.n288 71.676
R1839 B.n282 B.n150 71.676
R1840 B.n281 B.n154 71.676
R1841 B.n277 B.n276 71.676
R1842 B.n270 B.n156 71.676
R1843 B.n269 B.n268 71.676
R1844 B.n262 B.n158 71.676
R1845 B.n261 B.n260 71.676
R1846 B.n254 B.n160 71.676
R1847 B.n253 B.n252 71.676
R1848 B.n246 B.n162 71.676
R1849 B.n245 B.n244 71.676
R1850 B.n238 B.n164 71.676
R1851 B.n237 B.n236 71.676
R1852 B.n230 B.n166 71.676
R1853 B.n229 B.n228 71.676
R1854 B.n222 B.n168 71.676
R1855 B.n221 B.n220 71.676
R1856 B.n214 B.n170 71.676
R1857 B.n213 B.n212 71.676
R1858 B.n206 B.n172 71.676
R1859 B.n205 B.n204 71.676
R1860 B.n198 B.n174 71.676
R1861 B.n197 B.n196 71.676
R1862 B.n190 B.n176 71.676
R1863 B.n189 B.n188 71.676
R1864 B.n182 B.n178 71.676
R1865 B.n181 B.n180 71.676
R1866 B.n401 B.n400 71.676
R1867 B.n395 B.n120 71.676
R1868 B.n393 B.n392 71.676
R1869 B.n388 B.n387 71.676
R1870 B.n385 B.n384 71.676
R1871 B.n380 B.n379 71.676
R1872 B.n377 B.n376 71.676
R1873 B.n372 B.n371 71.676
R1874 B.n369 B.n368 71.676
R1875 B.n364 B.n363 71.676
R1876 B.n361 B.n360 71.676
R1877 B.n356 B.n355 71.676
R1878 B.n353 B.n352 71.676
R1879 B.n348 B.n347 71.676
R1880 B.n345 B.n344 71.676
R1881 B.n340 B.n339 71.676
R1882 B.n337 B.n336 71.676
R1883 B.n332 B.n331 71.676
R1884 B.n329 B.n328 71.676
R1885 B.n324 B.n323 71.676
R1886 B.n321 B.n320 71.676
R1887 B.n316 B.n315 71.676
R1888 B.n313 B.n312 71.676
R1889 B.n308 B.n307 71.676
R1890 B.n305 B.n304 71.676
R1891 B.n299 B.n298 71.676
R1892 B.n296 B.n295 71.676
R1893 B.n291 B.n290 71.676
R1894 B.n288 B.n287 71.676
R1895 B.n283 B.n282 71.676
R1896 B.n278 B.n154 71.676
R1897 B.n276 B.n275 71.676
R1898 B.n271 B.n270 71.676
R1899 B.n268 B.n267 71.676
R1900 B.n263 B.n262 71.676
R1901 B.n260 B.n259 71.676
R1902 B.n255 B.n254 71.676
R1903 B.n252 B.n251 71.676
R1904 B.n247 B.n246 71.676
R1905 B.n244 B.n243 71.676
R1906 B.n239 B.n238 71.676
R1907 B.n236 B.n235 71.676
R1908 B.n231 B.n230 71.676
R1909 B.n228 B.n227 71.676
R1910 B.n223 B.n222 71.676
R1911 B.n220 B.n219 71.676
R1912 B.n215 B.n214 71.676
R1913 B.n212 B.n211 71.676
R1914 B.n207 B.n206 71.676
R1915 B.n204 B.n203 71.676
R1916 B.n199 B.n198 71.676
R1917 B.n196 B.n195 71.676
R1918 B.n191 B.n190 71.676
R1919 B.n188 B.n187 71.676
R1920 B.n183 B.n182 71.676
R1921 B.n180 B.n116 71.676
R1922 B.n726 B.n725 71.676
R1923 B.n726 B.n2 71.676
R1924 B.n406 B.n117 64.4089
R1925 B.n697 B.n30 64.4089
R1926 B.n590 B.n59 59.5399
R1927 B.n572 B.n65 59.5399
R1928 B.n153 B.n152 59.5399
R1929 B.n301 B.n146 59.5399
R1930 B.n406 B.n113 36.197
R1931 B.n412 B.n113 36.197
R1932 B.n412 B.n109 36.197
R1933 B.n418 B.n109 36.197
R1934 B.n424 B.n105 36.197
R1935 B.n424 B.n100 36.197
R1936 B.n430 B.n100 36.197
R1937 B.n430 B.n101 36.197
R1938 B.n438 B.n437 36.197
R1939 B.n444 B.n4 36.197
R1940 B.n724 B.n4 36.197
R1941 B.n724 B.n723 36.197
R1942 B.n723 B.n722 36.197
R1943 B.n722 B.n8 36.197
R1944 B.n715 B.n12 36.197
R1945 B.n714 B.n713 36.197
R1946 B.n713 B.n16 36.197
R1947 B.n707 B.n16 36.197
R1948 B.n707 B.n706 36.197
R1949 B.n705 B.n23 36.197
R1950 B.n699 B.n23 36.197
R1951 B.n699 B.n698 36.197
R1952 B.n698 B.n697 36.197
R1953 B.n404 B.n403 30.7517
R1954 B.n408 B.n115 30.7517
R1955 B.n468 B.n467 30.7517
R1956 B.n695 B.n694 30.7517
R1957 B.n437 B.t3 30.3417
R1958 B.n12 B.t1 30.3417
R1959 B.n101 B.t0 26.0832
R1960 B.t2 B.n714 26.0832
R1961 B.t9 B.n105 21.8248
R1962 B.n706 B.t5 21.8248
R1963 B B.n727 18.0485
R1964 B.n418 B.t9 14.3726
R1965 B.t5 B.n705 14.3726
R1966 B.n59 B.n58 13.9641
R1967 B.n65 B.n64 13.9641
R1968 B.n152 B.n151 13.9641
R1969 B.n146 B.n145 13.9641
R1970 B.n404 B.n111 10.6151
R1971 B.n414 B.n111 10.6151
R1972 B.n415 B.n414 10.6151
R1973 B.n416 B.n415 10.6151
R1974 B.n416 B.n103 10.6151
R1975 B.n426 B.n103 10.6151
R1976 B.n427 B.n426 10.6151
R1977 B.n428 B.n427 10.6151
R1978 B.n428 B.n95 10.6151
R1979 B.n440 B.n95 10.6151
R1980 B.n441 B.n440 10.6151
R1981 B.n442 B.n441 10.6151
R1982 B.n442 B.n0 10.6151
R1983 B.n403 B.n402 10.6151
R1984 B.n402 B.n119 10.6151
R1985 B.n397 B.n119 10.6151
R1986 B.n397 B.n396 10.6151
R1987 B.n396 B.n121 10.6151
R1988 B.n391 B.n121 10.6151
R1989 B.n391 B.n390 10.6151
R1990 B.n390 B.n389 10.6151
R1991 B.n389 B.n123 10.6151
R1992 B.n383 B.n123 10.6151
R1993 B.n383 B.n382 10.6151
R1994 B.n382 B.n381 10.6151
R1995 B.n381 B.n125 10.6151
R1996 B.n375 B.n125 10.6151
R1997 B.n375 B.n374 10.6151
R1998 B.n374 B.n373 10.6151
R1999 B.n373 B.n127 10.6151
R2000 B.n367 B.n127 10.6151
R2001 B.n367 B.n366 10.6151
R2002 B.n366 B.n365 10.6151
R2003 B.n365 B.n129 10.6151
R2004 B.n359 B.n129 10.6151
R2005 B.n359 B.n358 10.6151
R2006 B.n358 B.n357 10.6151
R2007 B.n357 B.n131 10.6151
R2008 B.n351 B.n131 10.6151
R2009 B.n351 B.n350 10.6151
R2010 B.n350 B.n349 10.6151
R2011 B.n349 B.n133 10.6151
R2012 B.n343 B.n133 10.6151
R2013 B.n343 B.n342 10.6151
R2014 B.n342 B.n341 10.6151
R2015 B.n341 B.n135 10.6151
R2016 B.n335 B.n135 10.6151
R2017 B.n335 B.n334 10.6151
R2018 B.n334 B.n333 10.6151
R2019 B.n333 B.n137 10.6151
R2020 B.n327 B.n137 10.6151
R2021 B.n327 B.n326 10.6151
R2022 B.n326 B.n325 10.6151
R2023 B.n325 B.n139 10.6151
R2024 B.n319 B.n139 10.6151
R2025 B.n319 B.n318 10.6151
R2026 B.n318 B.n317 10.6151
R2027 B.n317 B.n141 10.6151
R2028 B.n311 B.n141 10.6151
R2029 B.n311 B.n310 10.6151
R2030 B.n310 B.n309 10.6151
R2031 B.n309 B.n143 10.6151
R2032 B.n303 B.n143 10.6151
R2033 B.n303 B.n302 10.6151
R2034 B.n300 B.n147 10.6151
R2035 B.n294 B.n147 10.6151
R2036 B.n294 B.n293 10.6151
R2037 B.n293 B.n292 10.6151
R2038 B.n292 B.n149 10.6151
R2039 B.n286 B.n149 10.6151
R2040 B.n286 B.n285 10.6151
R2041 B.n285 B.n284 10.6151
R2042 B.n280 B.n279 10.6151
R2043 B.n279 B.n155 10.6151
R2044 B.n274 B.n155 10.6151
R2045 B.n274 B.n273 10.6151
R2046 B.n273 B.n272 10.6151
R2047 B.n272 B.n157 10.6151
R2048 B.n266 B.n157 10.6151
R2049 B.n266 B.n265 10.6151
R2050 B.n265 B.n264 10.6151
R2051 B.n264 B.n159 10.6151
R2052 B.n258 B.n159 10.6151
R2053 B.n258 B.n257 10.6151
R2054 B.n257 B.n256 10.6151
R2055 B.n256 B.n161 10.6151
R2056 B.n250 B.n161 10.6151
R2057 B.n250 B.n249 10.6151
R2058 B.n249 B.n248 10.6151
R2059 B.n248 B.n163 10.6151
R2060 B.n242 B.n163 10.6151
R2061 B.n242 B.n241 10.6151
R2062 B.n241 B.n240 10.6151
R2063 B.n240 B.n165 10.6151
R2064 B.n234 B.n165 10.6151
R2065 B.n234 B.n233 10.6151
R2066 B.n233 B.n232 10.6151
R2067 B.n232 B.n167 10.6151
R2068 B.n226 B.n167 10.6151
R2069 B.n226 B.n225 10.6151
R2070 B.n225 B.n224 10.6151
R2071 B.n224 B.n169 10.6151
R2072 B.n218 B.n169 10.6151
R2073 B.n218 B.n217 10.6151
R2074 B.n217 B.n216 10.6151
R2075 B.n216 B.n171 10.6151
R2076 B.n210 B.n171 10.6151
R2077 B.n210 B.n209 10.6151
R2078 B.n209 B.n208 10.6151
R2079 B.n208 B.n173 10.6151
R2080 B.n202 B.n173 10.6151
R2081 B.n202 B.n201 10.6151
R2082 B.n201 B.n200 10.6151
R2083 B.n200 B.n175 10.6151
R2084 B.n194 B.n175 10.6151
R2085 B.n194 B.n193 10.6151
R2086 B.n193 B.n192 10.6151
R2087 B.n192 B.n177 10.6151
R2088 B.n186 B.n177 10.6151
R2089 B.n186 B.n185 10.6151
R2090 B.n185 B.n184 10.6151
R2091 B.n184 B.n179 10.6151
R2092 B.n179 B.n115 10.6151
R2093 B.n409 B.n408 10.6151
R2094 B.n410 B.n409 10.6151
R2095 B.n410 B.n107 10.6151
R2096 B.n420 B.n107 10.6151
R2097 B.n421 B.n420 10.6151
R2098 B.n422 B.n421 10.6151
R2099 B.n422 B.n98 10.6151
R2100 B.n432 B.n98 10.6151
R2101 B.n433 B.n432 10.6151
R2102 B.n435 B.n433 10.6151
R2103 B.n435 B.n434 10.6151
R2104 B.n434 B.n92 10.6151
R2105 B.n447 B.n92 10.6151
R2106 B.n448 B.n447 10.6151
R2107 B.n449 B.n448 10.6151
R2108 B.n450 B.n449 10.6151
R2109 B.n451 B.n450 10.6151
R2110 B.n454 B.n451 10.6151
R2111 B.n455 B.n454 10.6151
R2112 B.n456 B.n455 10.6151
R2113 B.n457 B.n456 10.6151
R2114 B.n459 B.n457 10.6151
R2115 B.n460 B.n459 10.6151
R2116 B.n461 B.n460 10.6151
R2117 B.n462 B.n461 10.6151
R2118 B.n464 B.n462 10.6151
R2119 B.n465 B.n464 10.6151
R2120 B.n466 B.n465 10.6151
R2121 B.n467 B.n466 10.6151
R2122 B.n719 B.n1 10.6151
R2123 B.n719 B.n718 10.6151
R2124 B.n718 B.n717 10.6151
R2125 B.n717 B.n10 10.6151
R2126 B.n711 B.n10 10.6151
R2127 B.n711 B.n710 10.6151
R2128 B.n710 B.n709 10.6151
R2129 B.n709 B.n18 10.6151
R2130 B.n703 B.n18 10.6151
R2131 B.n703 B.n702 10.6151
R2132 B.n702 B.n701 10.6151
R2133 B.n701 B.n25 10.6151
R2134 B.n695 B.n25 10.6151
R2135 B.n694 B.n693 10.6151
R2136 B.n693 B.n32 10.6151
R2137 B.n687 B.n32 10.6151
R2138 B.n687 B.n686 10.6151
R2139 B.n686 B.n685 10.6151
R2140 B.n685 B.n34 10.6151
R2141 B.n679 B.n34 10.6151
R2142 B.n679 B.n678 10.6151
R2143 B.n678 B.n677 10.6151
R2144 B.n677 B.n36 10.6151
R2145 B.n671 B.n36 10.6151
R2146 B.n671 B.n670 10.6151
R2147 B.n670 B.n669 10.6151
R2148 B.n669 B.n38 10.6151
R2149 B.n663 B.n38 10.6151
R2150 B.n663 B.n662 10.6151
R2151 B.n662 B.n661 10.6151
R2152 B.n661 B.n40 10.6151
R2153 B.n655 B.n40 10.6151
R2154 B.n655 B.n654 10.6151
R2155 B.n654 B.n653 10.6151
R2156 B.n653 B.n42 10.6151
R2157 B.n647 B.n42 10.6151
R2158 B.n647 B.n646 10.6151
R2159 B.n646 B.n645 10.6151
R2160 B.n645 B.n44 10.6151
R2161 B.n639 B.n44 10.6151
R2162 B.n639 B.n638 10.6151
R2163 B.n638 B.n637 10.6151
R2164 B.n637 B.n46 10.6151
R2165 B.n631 B.n46 10.6151
R2166 B.n631 B.n630 10.6151
R2167 B.n630 B.n629 10.6151
R2168 B.n629 B.n48 10.6151
R2169 B.n623 B.n48 10.6151
R2170 B.n623 B.n622 10.6151
R2171 B.n622 B.n621 10.6151
R2172 B.n621 B.n50 10.6151
R2173 B.n615 B.n50 10.6151
R2174 B.n615 B.n614 10.6151
R2175 B.n614 B.n613 10.6151
R2176 B.n613 B.n52 10.6151
R2177 B.n607 B.n52 10.6151
R2178 B.n607 B.n606 10.6151
R2179 B.n606 B.n605 10.6151
R2180 B.n605 B.n54 10.6151
R2181 B.n599 B.n54 10.6151
R2182 B.n599 B.n598 10.6151
R2183 B.n598 B.n597 10.6151
R2184 B.n597 B.n56 10.6151
R2185 B.n591 B.n56 10.6151
R2186 B.n589 B.n588 10.6151
R2187 B.n588 B.n60 10.6151
R2188 B.n582 B.n60 10.6151
R2189 B.n582 B.n581 10.6151
R2190 B.n581 B.n580 10.6151
R2191 B.n580 B.n62 10.6151
R2192 B.n574 B.n62 10.6151
R2193 B.n574 B.n573 10.6151
R2194 B.n571 B.n66 10.6151
R2195 B.n565 B.n66 10.6151
R2196 B.n565 B.n564 10.6151
R2197 B.n564 B.n563 10.6151
R2198 B.n563 B.n68 10.6151
R2199 B.n557 B.n68 10.6151
R2200 B.n557 B.n556 10.6151
R2201 B.n556 B.n555 10.6151
R2202 B.n555 B.n70 10.6151
R2203 B.n549 B.n70 10.6151
R2204 B.n549 B.n548 10.6151
R2205 B.n548 B.n547 10.6151
R2206 B.n547 B.n72 10.6151
R2207 B.n541 B.n72 10.6151
R2208 B.n541 B.n540 10.6151
R2209 B.n540 B.n539 10.6151
R2210 B.n539 B.n74 10.6151
R2211 B.n533 B.n74 10.6151
R2212 B.n533 B.n532 10.6151
R2213 B.n532 B.n531 10.6151
R2214 B.n531 B.n76 10.6151
R2215 B.n525 B.n76 10.6151
R2216 B.n525 B.n524 10.6151
R2217 B.n524 B.n523 10.6151
R2218 B.n523 B.n78 10.6151
R2219 B.n517 B.n78 10.6151
R2220 B.n517 B.n516 10.6151
R2221 B.n516 B.n515 10.6151
R2222 B.n515 B.n80 10.6151
R2223 B.n509 B.n80 10.6151
R2224 B.n509 B.n508 10.6151
R2225 B.n508 B.n507 10.6151
R2226 B.n507 B.n82 10.6151
R2227 B.n501 B.n82 10.6151
R2228 B.n501 B.n500 10.6151
R2229 B.n500 B.n499 10.6151
R2230 B.n499 B.n84 10.6151
R2231 B.n493 B.n84 10.6151
R2232 B.n493 B.n492 10.6151
R2233 B.n492 B.n491 10.6151
R2234 B.n491 B.n86 10.6151
R2235 B.n485 B.n86 10.6151
R2236 B.n485 B.n484 10.6151
R2237 B.n484 B.n483 10.6151
R2238 B.n483 B.n88 10.6151
R2239 B.n477 B.n88 10.6151
R2240 B.n477 B.n476 10.6151
R2241 B.n476 B.n475 10.6151
R2242 B.n475 B.n90 10.6151
R2243 B.n469 B.n90 10.6151
R2244 B.n469 B.n468 10.6151
R2245 B.n438 B.t0 10.1142
R2246 B.n715 B.t2 10.1142
R2247 B.n727 B.n0 8.11757
R2248 B.n727 B.n1 8.11757
R2249 B.n301 B.n300 7.18099
R2250 B.n284 B.n153 7.18099
R2251 B.n590 B.n589 7.18099
R2252 B.n573 B.n572 7.18099
R2253 B.n444 B.t3 5.85581
R2254 B.t1 B.n8 5.85581
R2255 B.n302 B.n301 3.43465
R2256 B.n280 B.n153 3.43465
R2257 B.n591 B.n590 3.43465
R2258 B.n572 B.n571 3.43465
R2259 VP.n1 VP.t2 1075.23
R2260 VP.n1 VP.t1 1075.23
R2261 VP.n0 VP.t0 1075.23
R2262 VP.n0 VP.t3 1075.23
R2263 VP.n2 VP.n0 203.482
R2264 VP.n2 VP.n1 161.3
R2265 VP VP.n2 0.0516364
R2266 VDD1 VDD1.n1 100.406
R2267 VDD1 VDD1.n0 61.0945
R2268 VDD1.n0 VDD1.t0 1.28872
R2269 VDD1.n0 VDD1.t3 1.28872
R2270 VDD1.n1 VDD1.t2 1.28872
R2271 VDD1.n1 VDD1.t1 1.28872
C0 VTAIL VN 2.33017f
C1 VN VDD2 2.96876f
C2 VTAIL VDD2 10.566299f
C3 VN VP 5.21377f
C4 VTAIL VP 2.34427f
C5 VP VDD2 0.25482f
C6 VN VDD1 0.148144f
C7 VTAIL VDD1 10.5269f
C8 VDD1 VDD2 0.497497f
C9 VDD1 VP 3.07526f
C10 VDD2 B 2.79073f
C11 VDD1 B 7.21497f
C12 VTAIL B 10.459539f
C13 VN B 9.01823f
C14 VP B 4.47137f
C15 VDD1.t0 B 0.380904f
C16 VDD1.t3 B 0.380904f
C17 VDD1.n0 B 3.44735f
C18 VDD1.t2 B 0.380904f
C19 VDD1.t1 B 0.380904f
C20 VDD1.n1 B 4.27449f
C21 VP.t3 B 1.01448f
C22 VP.t0 B 1.01448f
C23 VP.n0 B 1.28195f
C24 VP.t1 B 1.01448f
C25 VP.t2 B 1.01448f
C26 VP.n1 B 0.768441f
C27 VP.n2 B 4.4562f
C28 VDD2.t2 B 0.384176f
C29 VDD2.t0 B 0.384176f
C30 VDD2.n0 B 4.27957f
C31 VDD2.t1 B 0.384176f
C32 VDD2.t3 B 0.384176f
C33 VDD2.n1 B 3.47664f
C34 VDD2.n2 B 4.23702f
C35 VTAIL.n0 B 0.023049f
C36 VTAIL.n1 B 0.01767f
C37 VTAIL.n2 B 0.009495f
C38 VTAIL.n3 B 0.022443f
C39 VTAIL.n4 B 0.009774f
C40 VTAIL.n5 B 0.01767f
C41 VTAIL.n6 B 0.010054f
C42 VTAIL.n7 B 0.022443f
C43 VTAIL.n8 B 0.010054f
C44 VTAIL.n9 B 0.01767f
C45 VTAIL.n10 B 0.009495f
C46 VTAIL.n11 B 0.022443f
C47 VTAIL.n12 B 0.010054f
C48 VTAIL.n13 B 0.01767f
C49 VTAIL.n14 B 0.009495f
C50 VTAIL.n15 B 0.022443f
C51 VTAIL.n16 B 0.010054f
C52 VTAIL.n17 B 0.01767f
C53 VTAIL.n18 B 0.009495f
C54 VTAIL.n19 B 0.022443f
C55 VTAIL.n20 B 0.010054f
C56 VTAIL.n21 B 0.01767f
C57 VTAIL.n22 B 0.009495f
C58 VTAIL.n23 B 0.022443f
C59 VTAIL.n24 B 0.010054f
C60 VTAIL.n25 B 1.17961f
C61 VTAIL.n26 B 0.009495f
C62 VTAIL.t4 B 0.037028f
C63 VTAIL.n27 B 0.116888f
C64 VTAIL.n28 B 0.013258f
C65 VTAIL.n29 B 0.016832f
C66 VTAIL.n30 B 0.022443f
C67 VTAIL.n31 B 0.010054f
C68 VTAIL.n32 B 0.009495f
C69 VTAIL.n33 B 0.01767f
C70 VTAIL.n34 B 0.01767f
C71 VTAIL.n35 B 0.009495f
C72 VTAIL.n36 B 0.010054f
C73 VTAIL.n37 B 0.022443f
C74 VTAIL.n38 B 0.022443f
C75 VTAIL.n39 B 0.010054f
C76 VTAIL.n40 B 0.009495f
C77 VTAIL.n41 B 0.01767f
C78 VTAIL.n42 B 0.01767f
C79 VTAIL.n43 B 0.009495f
C80 VTAIL.n44 B 0.010054f
C81 VTAIL.n45 B 0.022443f
C82 VTAIL.n46 B 0.022443f
C83 VTAIL.n47 B 0.010054f
C84 VTAIL.n48 B 0.009495f
C85 VTAIL.n49 B 0.01767f
C86 VTAIL.n50 B 0.01767f
C87 VTAIL.n51 B 0.009495f
C88 VTAIL.n52 B 0.010054f
C89 VTAIL.n53 B 0.022443f
C90 VTAIL.n54 B 0.022443f
C91 VTAIL.n55 B 0.010054f
C92 VTAIL.n56 B 0.009495f
C93 VTAIL.n57 B 0.01767f
C94 VTAIL.n58 B 0.01767f
C95 VTAIL.n59 B 0.009495f
C96 VTAIL.n60 B 0.010054f
C97 VTAIL.n61 B 0.022443f
C98 VTAIL.n62 B 0.022443f
C99 VTAIL.n63 B 0.010054f
C100 VTAIL.n64 B 0.009495f
C101 VTAIL.n65 B 0.01767f
C102 VTAIL.n66 B 0.01767f
C103 VTAIL.n67 B 0.009495f
C104 VTAIL.n68 B 0.009495f
C105 VTAIL.n69 B 0.010054f
C106 VTAIL.n70 B 0.022443f
C107 VTAIL.n71 B 0.022443f
C108 VTAIL.n72 B 0.022443f
C109 VTAIL.n73 B 0.009774f
C110 VTAIL.n74 B 0.009495f
C111 VTAIL.n75 B 0.01767f
C112 VTAIL.n76 B 0.01767f
C113 VTAIL.n77 B 0.009495f
C114 VTAIL.n78 B 0.010054f
C115 VTAIL.n79 B 0.022443f
C116 VTAIL.n80 B 0.045423f
C117 VTAIL.n81 B 0.010054f
C118 VTAIL.n82 B 0.009495f
C119 VTAIL.n83 B 0.041085f
C120 VTAIL.n84 B 0.025098f
C121 VTAIL.n85 B 0.062962f
C122 VTAIL.n86 B 0.023049f
C123 VTAIL.n87 B 0.01767f
C124 VTAIL.n88 B 0.009495f
C125 VTAIL.n89 B 0.022443f
C126 VTAIL.n90 B 0.009774f
C127 VTAIL.n91 B 0.01767f
C128 VTAIL.n92 B 0.010054f
C129 VTAIL.n93 B 0.022443f
C130 VTAIL.n94 B 0.010054f
C131 VTAIL.n95 B 0.01767f
C132 VTAIL.n96 B 0.009495f
C133 VTAIL.n97 B 0.022443f
C134 VTAIL.n98 B 0.010054f
C135 VTAIL.n99 B 0.01767f
C136 VTAIL.n100 B 0.009495f
C137 VTAIL.n101 B 0.022443f
C138 VTAIL.n102 B 0.010054f
C139 VTAIL.n103 B 0.01767f
C140 VTAIL.n104 B 0.009495f
C141 VTAIL.n105 B 0.022443f
C142 VTAIL.n106 B 0.010054f
C143 VTAIL.n107 B 0.01767f
C144 VTAIL.n108 B 0.009495f
C145 VTAIL.n109 B 0.022443f
C146 VTAIL.n110 B 0.010054f
C147 VTAIL.n111 B 1.17961f
C148 VTAIL.n112 B 0.009495f
C149 VTAIL.t3 B 0.037028f
C150 VTAIL.n113 B 0.116888f
C151 VTAIL.n114 B 0.013258f
C152 VTAIL.n115 B 0.016832f
C153 VTAIL.n116 B 0.022443f
C154 VTAIL.n117 B 0.010054f
C155 VTAIL.n118 B 0.009495f
C156 VTAIL.n119 B 0.01767f
C157 VTAIL.n120 B 0.01767f
C158 VTAIL.n121 B 0.009495f
C159 VTAIL.n122 B 0.010054f
C160 VTAIL.n123 B 0.022443f
C161 VTAIL.n124 B 0.022443f
C162 VTAIL.n125 B 0.010054f
C163 VTAIL.n126 B 0.009495f
C164 VTAIL.n127 B 0.01767f
C165 VTAIL.n128 B 0.01767f
C166 VTAIL.n129 B 0.009495f
C167 VTAIL.n130 B 0.010054f
C168 VTAIL.n131 B 0.022443f
C169 VTAIL.n132 B 0.022443f
C170 VTAIL.n133 B 0.010054f
C171 VTAIL.n134 B 0.009495f
C172 VTAIL.n135 B 0.01767f
C173 VTAIL.n136 B 0.01767f
C174 VTAIL.n137 B 0.009495f
C175 VTAIL.n138 B 0.010054f
C176 VTAIL.n139 B 0.022443f
C177 VTAIL.n140 B 0.022443f
C178 VTAIL.n141 B 0.010054f
C179 VTAIL.n142 B 0.009495f
C180 VTAIL.n143 B 0.01767f
C181 VTAIL.n144 B 0.01767f
C182 VTAIL.n145 B 0.009495f
C183 VTAIL.n146 B 0.010054f
C184 VTAIL.n147 B 0.022443f
C185 VTAIL.n148 B 0.022443f
C186 VTAIL.n149 B 0.010054f
C187 VTAIL.n150 B 0.009495f
C188 VTAIL.n151 B 0.01767f
C189 VTAIL.n152 B 0.01767f
C190 VTAIL.n153 B 0.009495f
C191 VTAIL.n154 B 0.009495f
C192 VTAIL.n155 B 0.010054f
C193 VTAIL.n156 B 0.022443f
C194 VTAIL.n157 B 0.022443f
C195 VTAIL.n158 B 0.022443f
C196 VTAIL.n159 B 0.009774f
C197 VTAIL.n160 B 0.009495f
C198 VTAIL.n161 B 0.01767f
C199 VTAIL.n162 B 0.01767f
C200 VTAIL.n163 B 0.009495f
C201 VTAIL.n164 B 0.010054f
C202 VTAIL.n165 B 0.022443f
C203 VTAIL.n166 B 0.045423f
C204 VTAIL.n167 B 0.010054f
C205 VTAIL.n168 B 0.009495f
C206 VTAIL.n169 B 0.041085f
C207 VTAIL.n170 B 0.025098f
C208 VTAIL.n171 B 0.077319f
C209 VTAIL.n172 B 0.023049f
C210 VTAIL.n173 B 0.01767f
C211 VTAIL.n174 B 0.009495f
C212 VTAIL.n175 B 0.022443f
C213 VTAIL.n176 B 0.009774f
C214 VTAIL.n177 B 0.01767f
C215 VTAIL.n178 B 0.010054f
C216 VTAIL.n179 B 0.022443f
C217 VTAIL.n180 B 0.010054f
C218 VTAIL.n181 B 0.01767f
C219 VTAIL.n182 B 0.009495f
C220 VTAIL.n183 B 0.022443f
C221 VTAIL.n184 B 0.010054f
C222 VTAIL.n185 B 0.01767f
C223 VTAIL.n186 B 0.009495f
C224 VTAIL.n187 B 0.022443f
C225 VTAIL.n188 B 0.010054f
C226 VTAIL.n189 B 0.01767f
C227 VTAIL.n190 B 0.009495f
C228 VTAIL.n191 B 0.022443f
C229 VTAIL.n192 B 0.010054f
C230 VTAIL.n193 B 0.01767f
C231 VTAIL.n194 B 0.009495f
C232 VTAIL.n195 B 0.022443f
C233 VTAIL.n196 B 0.010054f
C234 VTAIL.n197 B 1.17961f
C235 VTAIL.n198 B 0.009495f
C236 VTAIL.t0 B 0.037028f
C237 VTAIL.n199 B 0.116888f
C238 VTAIL.n200 B 0.013258f
C239 VTAIL.n201 B 0.016832f
C240 VTAIL.n202 B 0.022443f
C241 VTAIL.n203 B 0.010054f
C242 VTAIL.n204 B 0.009495f
C243 VTAIL.n205 B 0.01767f
C244 VTAIL.n206 B 0.01767f
C245 VTAIL.n207 B 0.009495f
C246 VTAIL.n208 B 0.010054f
C247 VTAIL.n209 B 0.022443f
C248 VTAIL.n210 B 0.022443f
C249 VTAIL.n211 B 0.010054f
C250 VTAIL.n212 B 0.009495f
C251 VTAIL.n213 B 0.01767f
C252 VTAIL.n214 B 0.01767f
C253 VTAIL.n215 B 0.009495f
C254 VTAIL.n216 B 0.010054f
C255 VTAIL.n217 B 0.022443f
C256 VTAIL.n218 B 0.022443f
C257 VTAIL.n219 B 0.010054f
C258 VTAIL.n220 B 0.009495f
C259 VTAIL.n221 B 0.01767f
C260 VTAIL.n222 B 0.01767f
C261 VTAIL.n223 B 0.009495f
C262 VTAIL.n224 B 0.010054f
C263 VTAIL.n225 B 0.022443f
C264 VTAIL.n226 B 0.022443f
C265 VTAIL.n227 B 0.010054f
C266 VTAIL.n228 B 0.009495f
C267 VTAIL.n229 B 0.01767f
C268 VTAIL.n230 B 0.01767f
C269 VTAIL.n231 B 0.009495f
C270 VTAIL.n232 B 0.010054f
C271 VTAIL.n233 B 0.022443f
C272 VTAIL.n234 B 0.022443f
C273 VTAIL.n235 B 0.010054f
C274 VTAIL.n236 B 0.009495f
C275 VTAIL.n237 B 0.01767f
C276 VTAIL.n238 B 0.01767f
C277 VTAIL.n239 B 0.009495f
C278 VTAIL.n240 B 0.009495f
C279 VTAIL.n241 B 0.010054f
C280 VTAIL.n242 B 0.022443f
C281 VTAIL.n243 B 0.022443f
C282 VTAIL.n244 B 0.022443f
C283 VTAIL.n245 B 0.009774f
C284 VTAIL.n246 B 0.009495f
C285 VTAIL.n247 B 0.01767f
C286 VTAIL.n248 B 0.01767f
C287 VTAIL.n249 B 0.009495f
C288 VTAIL.n250 B 0.010054f
C289 VTAIL.n251 B 0.022443f
C290 VTAIL.n252 B 0.045423f
C291 VTAIL.n253 B 0.010054f
C292 VTAIL.n254 B 0.009495f
C293 VTAIL.n255 B 0.041085f
C294 VTAIL.n256 B 0.025098f
C295 VTAIL.n257 B 1.08134f
C296 VTAIL.n258 B 0.023049f
C297 VTAIL.n259 B 0.01767f
C298 VTAIL.n260 B 0.009495f
C299 VTAIL.n261 B 0.022443f
C300 VTAIL.n262 B 0.009774f
C301 VTAIL.n263 B 0.01767f
C302 VTAIL.n264 B 0.009774f
C303 VTAIL.n265 B 0.009495f
C304 VTAIL.n266 B 0.022443f
C305 VTAIL.n267 B 0.022443f
C306 VTAIL.n268 B 0.010054f
C307 VTAIL.n269 B 0.01767f
C308 VTAIL.n270 B 0.009495f
C309 VTAIL.n271 B 0.022443f
C310 VTAIL.n272 B 0.010054f
C311 VTAIL.n273 B 0.01767f
C312 VTAIL.n274 B 0.009495f
C313 VTAIL.n275 B 0.022443f
C314 VTAIL.n276 B 0.010054f
C315 VTAIL.n277 B 0.01767f
C316 VTAIL.n278 B 0.009495f
C317 VTAIL.n279 B 0.022443f
C318 VTAIL.n280 B 0.010054f
C319 VTAIL.n281 B 0.01767f
C320 VTAIL.n282 B 0.009495f
C321 VTAIL.n283 B 0.022443f
C322 VTAIL.n284 B 0.010054f
C323 VTAIL.n285 B 1.17961f
C324 VTAIL.n286 B 0.009495f
C325 VTAIL.t6 B 0.037028f
C326 VTAIL.n287 B 0.116888f
C327 VTAIL.n288 B 0.013258f
C328 VTAIL.n289 B 0.016832f
C329 VTAIL.n290 B 0.022443f
C330 VTAIL.n291 B 0.010054f
C331 VTAIL.n292 B 0.009495f
C332 VTAIL.n293 B 0.01767f
C333 VTAIL.n294 B 0.01767f
C334 VTAIL.n295 B 0.009495f
C335 VTAIL.n296 B 0.010054f
C336 VTAIL.n297 B 0.022443f
C337 VTAIL.n298 B 0.022443f
C338 VTAIL.n299 B 0.010054f
C339 VTAIL.n300 B 0.009495f
C340 VTAIL.n301 B 0.01767f
C341 VTAIL.n302 B 0.01767f
C342 VTAIL.n303 B 0.009495f
C343 VTAIL.n304 B 0.010054f
C344 VTAIL.n305 B 0.022443f
C345 VTAIL.n306 B 0.022443f
C346 VTAIL.n307 B 0.010054f
C347 VTAIL.n308 B 0.009495f
C348 VTAIL.n309 B 0.01767f
C349 VTAIL.n310 B 0.01767f
C350 VTAIL.n311 B 0.009495f
C351 VTAIL.n312 B 0.010054f
C352 VTAIL.n313 B 0.022443f
C353 VTAIL.n314 B 0.022443f
C354 VTAIL.n315 B 0.010054f
C355 VTAIL.n316 B 0.009495f
C356 VTAIL.n317 B 0.01767f
C357 VTAIL.n318 B 0.01767f
C358 VTAIL.n319 B 0.009495f
C359 VTAIL.n320 B 0.010054f
C360 VTAIL.n321 B 0.022443f
C361 VTAIL.n322 B 0.022443f
C362 VTAIL.n323 B 0.010054f
C363 VTAIL.n324 B 0.009495f
C364 VTAIL.n325 B 0.01767f
C365 VTAIL.n326 B 0.01767f
C366 VTAIL.n327 B 0.009495f
C367 VTAIL.n328 B 0.010054f
C368 VTAIL.n329 B 0.022443f
C369 VTAIL.n330 B 0.022443f
C370 VTAIL.n331 B 0.010054f
C371 VTAIL.n332 B 0.009495f
C372 VTAIL.n333 B 0.01767f
C373 VTAIL.n334 B 0.01767f
C374 VTAIL.n335 B 0.009495f
C375 VTAIL.n336 B 0.010054f
C376 VTAIL.n337 B 0.022443f
C377 VTAIL.n338 B 0.045423f
C378 VTAIL.n339 B 0.010054f
C379 VTAIL.n340 B 0.009495f
C380 VTAIL.n341 B 0.041085f
C381 VTAIL.n342 B 0.025098f
C382 VTAIL.n343 B 1.08134f
C383 VTAIL.n344 B 0.023049f
C384 VTAIL.n345 B 0.01767f
C385 VTAIL.n346 B 0.009495f
C386 VTAIL.n347 B 0.022443f
C387 VTAIL.n348 B 0.009774f
C388 VTAIL.n349 B 0.01767f
C389 VTAIL.n350 B 0.009774f
C390 VTAIL.n351 B 0.009495f
C391 VTAIL.n352 B 0.022443f
C392 VTAIL.n353 B 0.022443f
C393 VTAIL.n354 B 0.010054f
C394 VTAIL.n355 B 0.01767f
C395 VTAIL.n356 B 0.009495f
C396 VTAIL.n357 B 0.022443f
C397 VTAIL.n358 B 0.010054f
C398 VTAIL.n359 B 0.01767f
C399 VTAIL.n360 B 0.009495f
C400 VTAIL.n361 B 0.022443f
C401 VTAIL.n362 B 0.010054f
C402 VTAIL.n363 B 0.01767f
C403 VTAIL.n364 B 0.009495f
C404 VTAIL.n365 B 0.022443f
C405 VTAIL.n366 B 0.010054f
C406 VTAIL.n367 B 0.01767f
C407 VTAIL.n368 B 0.009495f
C408 VTAIL.n369 B 0.022443f
C409 VTAIL.n370 B 0.010054f
C410 VTAIL.n371 B 1.17961f
C411 VTAIL.n372 B 0.009495f
C412 VTAIL.t7 B 0.037028f
C413 VTAIL.n373 B 0.116888f
C414 VTAIL.n374 B 0.013258f
C415 VTAIL.n375 B 0.016832f
C416 VTAIL.n376 B 0.022443f
C417 VTAIL.n377 B 0.010054f
C418 VTAIL.n378 B 0.009495f
C419 VTAIL.n379 B 0.01767f
C420 VTAIL.n380 B 0.01767f
C421 VTAIL.n381 B 0.009495f
C422 VTAIL.n382 B 0.010054f
C423 VTAIL.n383 B 0.022443f
C424 VTAIL.n384 B 0.022443f
C425 VTAIL.n385 B 0.010054f
C426 VTAIL.n386 B 0.009495f
C427 VTAIL.n387 B 0.01767f
C428 VTAIL.n388 B 0.01767f
C429 VTAIL.n389 B 0.009495f
C430 VTAIL.n390 B 0.010054f
C431 VTAIL.n391 B 0.022443f
C432 VTAIL.n392 B 0.022443f
C433 VTAIL.n393 B 0.010054f
C434 VTAIL.n394 B 0.009495f
C435 VTAIL.n395 B 0.01767f
C436 VTAIL.n396 B 0.01767f
C437 VTAIL.n397 B 0.009495f
C438 VTAIL.n398 B 0.010054f
C439 VTAIL.n399 B 0.022443f
C440 VTAIL.n400 B 0.022443f
C441 VTAIL.n401 B 0.010054f
C442 VTAIL.n402 B 0.009495f
C443 VTAIL.n403 B 0.01767f
C444 VTAIL.n404 B 0.01767f
C445 VTAIL.n405 B 0.009495f
C446 VTAIL.n406 B 0.010054f
C447 VTAIL.n407 B 0.022443f
C448 VTAIL.n408 B 0.022443f
C449 VTAIL.n409 B 0.010054f
C450 VTAIL.n410 B 0.009495f
C451 VTAIL.n411 B 0.01767f
C452 VTAIL.n412 B 0.01767f
C453 VTAIL.n413 B 0.009495f
C454 VTAIL.n414 B 0.010054f
C455 VTAIL.n415 B 0.022443f
C456 VTAIL.n416 B 0.022443f
C457 VTAIL.n417 B 0.010054f
C458 VTAIL.n418 B 0.009495f
C459 VTAIL.n419 B 0.01767f
C460 VTAIL.n420 B 0.01767f
C461 VTAIL.n421 B 0.009495f
C462 VTAIL.n422 B 0.010054f
C463 VTAIL.n423 B 0.022443f
C464 VTAIL.n424 B 0.045423f
C465 VTAIL.n425 B 0.010054f
C466 VTAIL.n426 B 0.009495f
C467 VTAIL.n427 B 0.041085f
C468 VTAIL.n428 B 0.025098f
C469 VTAIL.n429 B 0.077319f
C470 VTAIL.n430 B 0.023049f
C471 VTAIL.n431 B 0.01767f
C472 VTAIL.n432 B 0.009495f
C473 VTAIL.n433 B 0.022443f
C474 VTAIL.n434 B 0.009774f
C475 VTAIL.n435 B 0.01767f
C476 VTAIL.n436 B 0.009774f
C477 VTAIL.n437 B 0.009495f
C478 VTAIL.n438 B 0.022443f
C479 VTAIL.n439 B 0.022443f
C480 VTAIL.n440 B 0.010054f
C481 VTAIL.n441 B 0.01767f
C482 VTAIL.n442 B 0.009495f
C483 VTAIL.n443 B 0.022443f
C484 VTAIL.n444 B 0.010054f
C485 VTAIL.n445 B 0.01767f
C486 VTAIL.n446 B 0.009495f
C487 VTAIL.n447 B 0.022443f
C488 VTAIL.n448 B 0.010054f
C489 VTAIL.n449 B 0.01767f
C490 VTAIL.n450 B 0.009495f
C491 VTAIL.n451 B 0.022443f
C492 VTAIL.n452 B 0.010054f
C493 VTAIL.n453 B 0.01767f
C494 VTAIL.n454 B 0.009495f
C495 VTAIL.n455 B 0.022443f
C496 VTAIL.n456 B 0.010054f
C497 VTAIL.n457 B 1.17961f
C498 VTAIL.n458 B 0.009495f
C499 VTAIL.t1 B 0.037028f
C500 VTAIL.n459 B 0.116888f
C501 VTAIL.n460 B 0.013258f
C502 VTAIL.n461 B 0.016832f
C503 VTAIL.n462 B 0.022443f
C504 VTAIL.n463 B 0.010054f
C505 VTAIL.n464 B 0.009495f
C506 VTAIL.n465 B 0.01767f
C507 VTAIL.n466 B 0.01767f
C508 VTAIL.n467 B 0.009495f
C509 VTAIL.n468 B 0.010054f
C510 VTAIL.n469 B 0.022443f
C511 VTAIL.n470 B 0.022443f
C512 VTAIL.n471 B 0.010054f
C513 VTAIL.n472 B 0.009495f
C514 VTAIL.n473 B 0.01767f
C515 VTAIL.n474 B 0.01767f
C516 VTAIL.n475 B 0.009495f
C517 VTAIL.n476 B 0.010054f
C518 VTAIL.n477 B 0.022443f
C519 VTAIL.n478 B 0.022443f
C520 VTAIL.n479 B 0.010054f
C521 VTAIL.n480 B 0.009495f
C522 VTAIL.n481 B 0.01767f
C523 VTAIL.n482 B 0.01767f
C524 VTAIL.n483 B 0.009495f
C525 VTAIL.n484 B 0.010054f
C526 VTAIL.n485 B 0.022443f
C527 VTAIL.n486 B 0.022443f
C528 VTAIL.n487 B 0.010054f
C529 VTAIL.n488 B 0.009495f
C530 VTAIL.n489 B 0.01767f
C531 VTAIL.n490 B 0.01767f
C532 VTAIL.n491 B 0.009495f
C533 VTAIL.n492 B 0.010054f
C534 VTAIL.n493 B 0.022443f
C535 VTAIL.n494 B 0.022443f
C536 VTAIL.n495 B 0.010054f
C537 VTAIL.n496 B 0.009495f
C538 VTAIL.n497 B 0.01767f
C539 VTAIL.n498 B 0.01767f
C540 VTAIL.n499 B 0.009495f
C541 VTAIL.n500 B 0.010054f
C542 VTAIL.n501 B 0.022443f
C543 VTAIL.n502 B 0.022443f
C544 VTAIL.n503 B 0.010054f
C545 VTAIL.n504 B 0.009495f
C546 VTAIL.n505 B 0.01767f
C547 VTAIL.n506 B 0.01767f
C548 VTAIL.n507 B 0.009495f
C549 VTAIL.n508 B 0.010054f
C550 VTAIL.n509 B 0.022443f
C551 VTAIL.n510 B 0.045423f
C552 VTAIL.n511 B 0.010054f
C553 VTAIL.n512 B 0.009495f
C554 VTAIL.n513 B 0.041085f
C555 VTAIL.n514 B 0.025098f
C556 VTAIL.n515 B 0.077319f
C557 VTAIL.n516 B 0.023049f
C558 VTAIL.n517 B 0.01767f
C559 VTAIL.n518 B 0.009495f
C560 VTAIL.n519 B 0.022443f
C561 VTAIL.n520 B 0.009774f
C562 VTAIL.n521 B 0.01767f
C563 VTAIL.n522 B 0.009774f
C564 VTAIL.n523 B 0.009495f
C565 VTAIL.n524 B 0.022443f
C566 VTAIL.n525 B 0.022443f
C567 VTAIL.n526 B 0.010054f
C568 VTAIL.n527 B 0.01767f
C569 VTAIL.n528 B 0.009495f
C570 VTAIL.n529 B 0.022443f
C571 VTAIL.n530 B 0.010054f
C572 VTAIL.n531 B 0.01767f
C573 VTAIL.n532 B 0.009495f
C574 VTAIL.n533 B 0.022443f
C575 VTAIL.n534 B 0.010054f
C576 VTAIL.n535 B 0.01767f
C577 VTAIL.n536 B 0.009495f
C578 VTAIL.n537 B 0.022443f
C579 VTAIL.n538 B 0.010054f
C580 VTAIL.n539 B 0.01767f
C581 VTAIL.n540 B 0.009495f
C582 VTAIL.n541 B 0.022443f
C583 VTAIL.n542 B 0.010054f
C584 VTAIL.n543 B 1.17961f
C585 VTAIL.n544 B 0.009495f
C586 VTAIL.t2 B 0.037028f
C587 VTAIL.n545 B 0.116888f
C588 VTAIL.n546 B 0.013258f
C589 VTAIL.n547 B 0.016832f
C590 VTAIL.n548 B 0.022443f
C591 VTAIL.n549 B 0.010054f
C592 VTAIL.n550 B 0.009495f
C593 VTAIL.n551 B 0.01767f
C594 VTAIL.n552 B 0.01767f
C595 VTAIL.n553 B 0.009495f
C596 VTAIL.n554 B 0.010054f
C597 VTAIL.n555 B 0.022443f
C598 VTAIL.n556 B 0.022443f
C599 VTAIL.n557 B 0.010054f
C600 VTAIL.n558 B 0.009495f
C601 VTAIL.n559 B 0.01767f
C602 VTAIL.n560 B 0.01767f
C603 VTAIL.n561 B 0.009495f
C604 VTAIL.n562 B 0.010054f
C605 VTAIL.n563 B 0.022443f
C606 VTAIL.n564 B 0.022443f
C607 VTAIL.n565 B 0.010054f
C608 VTAIL.n566 B 0.009495f
C609 VTAIL.n567 B 0.01767f
C610 VTAIL.n568 B 0.01767f
C611 VTAIL.n569 B 0.009495f
C612 VTAIL.n570 B 0.010054f
C613 VTAIL.n571 B 0.022443f
C614 VTAIL.n572 B 0.022443f
C615 VTAIL.n573 B 0.010054f
C616 VTAIL.n574 B 0.009495f
C617 VTAIL.n575 B 0.01767f
C618 VTAIL.n576 B 0.01767f
C619 VTAIL.n577 B 0.009495f
C620 VTAIL.n578 B 0.010054f
C621 VTAIL.n579 B 0.022443f
C622 VTAIL.n580 B 0.022443f
C623 VTAIL.n581 B 0.010054f
C624 VTAIL.n582 B 0.009495f
C625 VTAIL.n583 B 0.01767f
C626 VTAIL.n584 B 0.01767f
C627 VTAIL.n585 B 0.009495f
C628 VTAIL.n586 B 0.010054f
C629 VTAIL.n587 B 0.022443f
C630 VTAIL.n588 B 0.022443f
C631 VTAIL.n589 B 0.010054f
C632 VTAIL.n590 B 0.009495f
C633 VTAIL.n591 B 0.01767f
C634 VTAIL.n592 B 0.01767f
C635 VTAIL.n593 B 0.009495f
C636 VTAIL.n594 B 0.010054f
C637 VTAIL.n595 B 0.022443f
C638 VTAIL.n596 B 0.045423f
C639 VTAIL.n597 B 0.010054f
C640 VTAIL.n598 B 0.009495f
C641 VTAIL.n599 B 0.041085f
C642 VTAIL.n600 B 0.025098f
C643 VTAIL.n601 B 1.08134f
C644 VTAIL.n602 B 0.023049f
C645 VTAIL.n603 B 0.01767f
C646 VTAIL.n604 B 0.009495f
C647 VTAIL.n605 B 0.022443f
C648 VTAIL.n606 B 0.009774f
C649 VTAIL.n607 B 0.01767f
C650 VTAIL.n608 B 0.010054f
C651 VTAIL.n609 B 0.022443f
C652 VTAIL.n610 B 0.010054f
C653 VTAIL.n611 B 0.01767f
C654 VTAIL.n612 B 0.009495f
C655 VTAIL.n613 B 0.022443f
C656 VTAIL.n614 B 0.010054f
C657 VTAIL.n615 B 0.01767f
C658 VTAIL.n616 B 0.009495f
C659 VTAIL.n617 B 0.022443f
C660 VTAIL.n618 B 0.010054f
C661 VTAIL.n619 B 0.01767f
C662 VTAIL.n620 B 0.009495f
C663 VTAIL.n621 B 0.022443f
C664 VTAIL.n622 B 0.010054f
C665 VTAIL.n623 B 0.01767f
C666 VTAIL.n624 B 0.009495f
C667 VTAIL.n625 B 0.022443f
C668 VTAIL.n626 B 0.010054f
C669 VTAIL.n627 B 1.17961f
C670 VTAIL.n628 B 0.009495f
C671 VTAIL.t5 B 0.037028f
C672 VTAIL.n629 B 0.116888f
C673 VTAIL.n630 B 0.013258f
C674 VTAIL.n631 B 0.016832f
C675 VTAIL.n632 B 0.022443f
C676 VTAIL.n633 B 0.010054f
C677 VTAIL.n634 B 0.009495f
C678 VTAIL.n635 B 0.01767f
C679 VTAIL.n636 B 0.01767f
C680 VTAIL.n637 B 0.009495f
C681 VTAIL.n638 B 0.010054f
C682 VTAIL.n639 B 0.022443f
C683 VTAIL.n640 B 0.022443f
C684 VTAIL.n641 B 0.010054f
C685 VTAIL.n642 B 0.009495f
C686 VTAIL.n643 B 0.01767f
C687 VTAIL.n644 B 0.01767f
C688 VTAIL.n645 B 0.009495f
C689 VTAIL.n646 B 0.010054f
C690 VTAIL.n647 B 0.022443f
C691 VTAIL.n648 B 0.022443f
C692 VTAIL.n649 B 0.010054f
C693 VTAIL.n650 B 0.009495f
C694 VTAIL.n651 B 0.01767f
C695 VTAIL.n652 B 0.01767f
C696 VTAIL.n653 B 0.009495f
C697 VTAIL.n654 B 0.010054f
C698 VTAIL.n655 B 0.022443f
C699 VTAIL.n656 B 0.022443f
C700 VTAIL.n657 B 0.010054f
C701 VTAIL.n658 B 0.009495f
C702 VTAIL.n659 B 0.01767f
C703 VTAIL.n660 B 0.01767f
C704 VTAIL.n661 B 0.009495f
C705 VTAIL.n662 B 0.010054f
C706 VTAIL.n663 B 0.022443f
C707 VTAIL.n664 B 0.022443f
C708 VTAIL.n665 B 0.010054f
C709 VTAIL.n666 B 0.009495f
C710 VTAIL.n667 B 0.01767f
C711 VTAIL.n668 B 0.01767f
C712 VTAIL.n669 B 0.009495f
C713 VTAIL.n670 B 0.009495f
C714 VTAIL.n671 B 0.010054f
C715 VTAIL.n672 B 0.022443f
C716 VTAIL.n673 B 0.022443f
C717 VTAIL.n674 B 0.022443f
C718 VTAIL.n675 B 0.009774f
C719 VTAIL.n676 B 0.009495f
C720 VTAIL.n677 B 0.01767f
C721 VTAIL.n678 B 0.01767f
C722 VTAIL.n679 B 0.009495f
C723 VTAIL.n680 B 0.010054f
C724 VTAIL.n681 B 0.022443f
C725 VTAIL.n682 B 0.045423f
C726 VTAIL.n683 B 0.010054f
C727 VTAIL.n684 B 0.009495f
C728 VTAIL.n685 B 0.041085f
C729 VTAIL.n686 B 0.025098f
C730 VTAIL.n687 B 1.06035f
C731 VN.t1 B 0.997097f
C732 VN.t3 B 0.997097f
C733 VN.n0 B 0.755298f
C734 VN.t2 B 0.997097f
C735 VN.t0 B 0.997097f
C736 VN.n1 B 1.27155f
.ends

