* NGSPICE file created from diff_pair_sample_0156.ext - technology: sky130A

.subckt diff_pair_sample_0156 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=4.446 ps=23.58 w=11.4 l=1.43
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=0 ps=0 w=11.4 l=1.43
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=4.446 ps=23.58 w=11.4 l=1.43
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=0 ps=0 w=11.4 l=1.43
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=4.446 ps=23.58 w=11.4 l=1.43
X5 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=4.446 ps=23.58 w=11.4 l=1.43
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=0 ps=0 w=11.4 l=1.43
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.446 pd=23.58 as=0 ps=0 w=11.4 l=1.43
R0 VP.n0 VP.t0 341.637
R1 VP.n0 VP.t1 300.538
R2 VP VP.n0 0.146778
R3 VTAIL.n242 VTAIL.n186 289.615
R4 VTAIL.n56 VTAIL.n0 289.615
R5 VTAIL.n180 VTAIL.n124 289.615
R6 VTAIL.n118 VTAIL.n62 289.615
R7 VTAIL.n207 VTAIL.n206 185
R8 VTAIL.n209 VTAIL.n208 185
R9 VTAIL.n202 VTAIL.n201 185
R10 VTAIL.n215 VTAIL.n214 185
R11 VTAIL.n217 VTAIL.n216 185
R12 VTAIL.n198 VTAIL.n197 185
R13 VTAIL.n224 VTAIL.n223 185
R14 VTAIL.n225 VTAIL.n196 185
R15 VTAIL.n227 VTAIL.n226 185
R16 VTAIL.n194 VTAIL.n193 185
R17 VTAIL.n233 VTAIL.n232 185
R18 VTAIL.n235 VTAIL.n234 185
R19 VTAIL.n190 VTAIL.n189 185
R20 VTAIL.n241 VTAIL.n240 185
R21 VTAIL.n243 VTAIL.n242 185
R22 VTAIL.n21 VTAIL.n20 185
R23 VTAIL.n23 VTAIL.n22 185
R24 VTAIL.n16 VTAIL.n15 185
R25 VTAIL.n29 VTAIL.n28 185
R26 VTAIL.n31 VTAIL.n30 185
R27 VTAIL.n12 VTAIL.n11 185
R28 VTAIL.n38 VTAIL.n37 185
R29 VTAIL.n39 VTAIL.n10 185
R30 VTAIL.n41 VTAIL.n40 185
R31 VTAIL.n8 VTAIL.n7 185
R32 VTAIL.n47 VTAIL.n46 185
R33 VTAIL.n49 VTAIL.n48 185
R34 VTAIL.n4 VTAIL.n3 185
R35 VTAIL.n55 VTAIL.n54 185
R36 VTAIL.n57 VTAIL.n56 185
R37 VTAIL.n181 VTAIL.n180 185
R38 VTAIL.n179 VTAIL.n178 185
R39 VTAIL.n128 VTAIL.n127 185
R40 VTAIL.n173 VTAIL.n172 185
R41 VTAIL.n171 VTAIL.n170 185
R42 VTAIL.n132 VTAIL.n131 185
R43 VTAIL.n136 VTAIL.n134 185
R44 VTAIL.n165 VTAIL.n164 185
R45 VTAIL.n163 VTAIL.n162 185
R46 VTAIL.n138 VTAIL.n137 185
R47 VTAIL.n157 VTAIL.n156 185
R48 VTAIL.n155 VTAIL.n154 185
R49 VTAIL.n142 VTAIL.n141 185
R50 VTAIL.n149 VTAIL.n148 185
R51 VTAIL.n147 VTAIL.n146 185
R52 VTAIL.n119 VTAIL.n118 185
R53 VTAIL.n117 VTAIL.n116 185
R54 VTAIL.n66 VTAIL.n65 185
R55 VTAIL.n111 VTAIL.n110 185
R56 VTAIL.n109 VTAIL.n108 185
R57 VTAIL.n70 VTAIL.n69 185
R58 VTAIL.n74 VTAIL.n72 185
R59 VTAIL.n103 VTAIL.n102 185
R60 VTAIL.n101 VTAIL.n100 185
R61 VTAIL.n76 VTAIL.n75 185
R62 VTAIL.n95 VTAIL.n94 185
R63 VTAIL.n93 VTAIL.n92 185
R64 VTAIL.n80 VTAIL.n79 185
R65 VTAIL.n87 VTAIL.n86 185
R66 VTAIL.n85 VTAIL.n84 185
R67 VTAIL.n205 VTAIL.t0 149.524
R68 VTAIL.n19 VTAIL.t2 149.524
R69 VTAIL.n145 VTAIL.t3 149.524
R70 VTAIL.n83 VTAIL.t1 149.524
R71 VTAIL.n208 VTAIL.n207 104.615
R72 VTAIL.n208 VTAIL.n201 104.615
R73 VTAIL.n215 VTAIL.n201 104.615
R74 VTAIL.n216 VTAIL.n215 104.615
R75 VTAIL.n216 VTAIL.n197 104.615
R76 VTAIL.n224 VTAIL.n197 104.615
R77 VTAIL.n225 VTAIL.n224 104.615
R78 VTAIL.n226 VTAIL.n225 104.615
R79 VTAIL.n226 VTAIL.n193 104.615
R80 VTAIL.n233 VTAIL.n193 104.615
R81 VTAIL.n234 VTAIL.n233 104.615
R82 VTAIL.n234 VTAIL.n189 104.615
R83 VTAIL.n241 VTAIL.n189 104.615
R84 VTAIL.n242 VTAIL.n241 104.615
R85 VTAIL.n22 VTAIL.n21 104.615
R86 VTAIL.n22 VTAIL.n15 104.615
R87 VTAIL.n29 VTAIL.n15 104.615
R88 VTAIL.n30 VTAIL.n29 104.615
R89 VTAIL.n30 VTAIL.n11 104.615
R90 VTAIL.n38 VTAIL.n11 104.615
R91 VTAIL.n39 VTAIL.n38 104.615
R92 VTAIL.n40 VTAIL.n39 104.615
R93 VTAIL.n40 VTAIL.n7 104.615
R94 VTAIL.n47 VTAIL.n7 104.615
R95 VTAIL.n48 VTAIL.n47 104.615
R96 VTAIL.n48 VTAIL.n3 104.615
R97 VTAIL.n55 VTAIL.n3 104.615
R98 VTAIL.n56 VTAIL.n55 104.615
R99 VTAIL.n180 VTAIL.n179 104.615
R100 VTAIL.n179 VTAIL.n127 104.615
R101 VTAIL.n172 VTAIL.n127 104.615
R102 VTAIL.n172 VTAIL.n171 104.615
R103 VTAIL.n171 VTAIL.n131 104.615
R104 VTAIL.n136 VTAIL.n131 104.615
R105 VTAIL.n164 VTAIL.n136 104.615
R106 VTAIL.n164 VTAIL.n163 104.615
R107 VTAIL.n163 VTAIL.n137 104.615
R108 VTAIL.n156 VTAIL.n137 104.615
R109 VTAIL.n156 VTAIL.n155 104.615
R110 VTAIL.n155 VTAIL.n141 104.615
R111 VTAIL.n148 VTAIL.n141 104.615
R112 VTAIL.n148 VTAIL.n147 104.615
R113 VTAIL.n118 VTAIL.n117 104.615
R114 VTAIL.n117 VTAIL.n65 104.615
R115 VTAIL.n110 VTAIL.n65 104.615
R116 VTAIL.n110 VTAIL.n109 104.615
R117 VTAIL.n109 VTAIL.n69 104.615
R118 VTAIL.n74 VTAIL.n69 104.615
R119 VTAIL.n102 VTAIL.n74 104.615
R120 VTAIL.n102 VTAIL.n101 104.615
R121 VTAIL.n101 VTAIL.n75 104.615
R122 VTAIL.n94 VTAIL.n75 104.615
R123 VTAIL.n94 VTAIL.n93 104.615
R124 VTAIL.n93 VTAIL.n79 104.615
R125 VTAIL.n86 VTAIL.n79 104.615
R126 VTAIL.n86 VTAIL.n85 104.615
R127 VTAIL.n207 VTAIL.t0 52.3082
R128 VTAIL.n21 VTAIL.t2 52.3082
R129 VTAIL.n147 VTAIL.t3 52.3082
R130 VTAIL.n85 VTAIL.t1 52.3082
R131 VTAIL.n247 VTAIL.n246 32.1853
R132 VTAIL.n61 VTAIL.n60 32.1853
R133 VTAIL.n185 VTAIL.n184 32.1853
R134 VTAIL.n123 VTAIL.n122 32.1853
R135 VTAIL.n123 VTAIL.n61 25.2289
R136 VTAIL.n247 VTAIL.n185 23.7117
R137 VTAIL.n227 VTAIL.n194 13.1884
R138 VTAIL.n41 VTAIL.n8 13.1884
R139 VTAIL.n134 VTAIL.n132 13.1884
R140 VTAIL.n72 VTAIL.n70 13.1884
R141 VTAIL.n228 VTAIL.n196 12.8005
R142 VTAIL.n232 VTAIL.n231 12.8005
R143 VTAIL.n42 VTAIL.n10 12.8005
R144 VTAIL.n46 VTAIL.n45 12.8005
R145 VTAIL.n170 VTAIL.n169 12.8005
R146 VTAIL.n166 VTAIL.n165 12.8005
R147 VTAIL.n108 VTAIL.n107 12.8005
R148 VTAIL.n104 VTAIL.n103 12.8005
R149 VTAIL.n223 VTAIL.n222 12.0247
R150 VTAIL.n235 VTAIL.n192 12.0247
R151 VTAIL.n37 VTAIL.n36 12.0247
R152 VTAIL.n49 VTAIL.n6 12.0247
R153 VTAIL.n173 VTAIL.n130 12.0247
R154 VTAIL.n162 VTAIL.n135 12.0247
R155 VTAIL.n111 VTAIL.n68 12.0247
R156 VTAIL.n100 VTAIL.n73 12.0247
R157 VTAIL.n221 VTAIL.n198 11.249
R158 VTAIL.n236 VTAIL.n190 11.249
R159 VTAIL.n35 VTAIL.n12 11.249
R160 VTAIL.n50 VTAIL.n4 11.249
R161 VTAIL.n174 VTAIL.n128 11.249
R162 VTAIL.n161 VTAIL.n138 11.249
R163 VTAIL.n112 VTAIL.n66 11.249
R164 VTAIL.n99 VTAIL.n76 11.249
R165 VTAIL.n218 VTAIL.n217 10.4732
R166 VTAIL.n240 VTAIL.n239 10.4732
R167 VTAIL.n32 VTAIL.n31 10.4732
R168 VTAIL.n54 VTAIL.n53 10.4732
R169 VTAIL.n178 VTAIL.n177 10.4732
R170 VTAIL.n158 VTAIL.n157 10.4732
R171 VTAIL.n116 VTAIL.n115 10.4732
R172 VTAIL.n96 VTAIL.n95 10.4732
R173 VTAIL.n206 VTAIL.n205 10.2747
R174 VTAIL.n20 VTAIL.n19 10.2747
R175 VTAIL.n146 VTAIL.n145 10.2747
R176 VTAIL.n84 VTAIL.n83 10.2747
R177 VTAIL.n214 VTAIL.n200 9.69747
R178 VTAIL.n243 VTAIL.n188 9.69747
R179 VTAIL.n28 VTAIL.n14 9.69747
R180 VTAIL.n57 VTAIL.n2 9.69747
R181 VTAIL.n181 VTAIL.n126 9.69747
R182 VTAIL.n154 VTAIL.n140 9.69747
R183 VTAIL.n119 VTAIL.n64 9.69747
R184 VTAIL.n92 VTAIL.n78 9.69747
R185 VTAIL.n246 VTAIL.n245 9.45567
R186 VTAIL.n60 VTAIL.n59 9.45567
R187 VTAIL.n184 VTAIL.n183 9.45567
R188 VTAIL.n122 VTAIL.n121 9.45567
R189 VTAIL.n245 VTAIL.n244 9.3005
R190 VTAIL.n188 VTAIL.n187 9.3005
R191 VTAIL.n239 VTAIL.n238 9.3005
R192 VTAIL.n237 VTAIL.n236 9.3005
R193 VTAIL.n192 VTAIL.n191 9.3005
R194 VTAIL.n231 VTAIL.n230 9.3005
R195 VTAIL.n204 VTAIL.n203 9.3005
R196 VTAIL.n211 VTAIL.n210 9.3005
R197 VTAIL.n213 VTAIL.n212 9.3005
R198 VTAIL.n200 VTAIL.n199 9.3005
R199 VTAIL.n219 VTAIL.n218 9.3005
R200 VTAIL.n221 VTAIL.n220 9.3005
R201 VTAIL.n222 VTAIL.n195 9.3005
R202 VTAIL.n229 VTAIL.n228 9.3005
R203 VTAIL.n59 VTAIL.n58 9.3005
R204 VTAIL.n2 VTAIL.n1 9.3005
R205 VTAIL.n53 VTAIL.n52 9.3005
R206 VTAIL.n51 VTAIL.n50 9.3005
R207 VTAIL.n6 VTAIL.n5 9.3005
R208 VTAIL.n45 VTAIL.n44 9.3005
R209 VTAIL.n18 VTAIL.n17 9.3005
R210 VTAIL.n25 VTAIL.n24 9.3005
R211 VTAIL.n27 VTAIL.n26 9.3005
R212 VTAIL.n14 VTAIL.n13 9.3005
R213 VTAIL.n33 VTAIL.n32 9.3005
R214 VTAIL.n35 VTAIL.n34 9.3005
R215 VTAIL.n36 VTAIL.n9 9.3005
R216 VTAIL.n43 VTAIL.n42 9.3005
R217 VTAIL.n144 VTAIL.n143 9.3005
R218 VTAIL.n151 VTAIL.n150 9.3005
R219 VTAIL.n153 VTAIL.n152 9.3005
R220 VTAIL.n140 VTAIL.n139 9.3005
R221 VTAIL.n159 VTAIL.n158 9.3005
R222 VTAIL.n161 VTAIL.n160 9.3005
R223 VTAIL.n135 VTAIL.n133 9.3005
R224 VTAIL.n167 VTAIL.n166 9.3005
R225 VTAIL.n183 VTAIL.n182 9.3005
R226 VTAIL.n126 VTAIL.n125 9.3005
R227 VTAIL.n177 VTAIL.n176 9.3005
R228 VTAIL.n175 VTAIL.n174 9.3005
R229 VTAIL.n130 VTAIL.n129 9.3005
R230 VTAIL.n169 VTAIL.n168 9.3005
R231 VTAIL.n82 VTAIL.n81 9.3005
R232 VTAIL.n89 VTAIL.n88 9.3005
R233 VTAIL.n91 VTAIL.n90 9.3005
R234 VTAIL.n78 VTAIL.n77 9.3005
R235 VTAIL.n97 VTAIL.n96 9.3005
R236 VTAIL.n99 VTAIL.n98 9.3005
R237 VTAIL.n73 VTAIL.n71 9.3005
R238 VTAIL.n105 VTAIL.n104 9.3005
R239 VTAIL.n121 VTAIL.n120 9.3005
R240 VTAIL.n64 VTAIL.n63 9.3005
R241 VTAIL.n115 VTAIL.n114 9.3005
R242 VTAIL.n113 VTAIL.n112 9.3005
R243 VTAIL.n68 VTAIL.n67 9.3005
R244 VTAIL.n107 VTAIL.n106 9.3005
R245 VTAIL.n213 VTAIL.n202 8.92171
R246 VTAIL.n244 VTAIL.n186 8.92171
R247 VTAIL.n27 VTAIL.n16 8.92171
R248 VTAIL.n58 VTAIL.n0 8.92171
R249 VTAIL.n182 VTAIL.n124 8.92171
R250 VTAIL.n153 VTAIL.n142 8.92171
R251 VTAIL.n120 VTAIL.n62 8.92171
R252 VTAIL.n91 VTAIL.n80 8.92171
R253 VTAIL.n210 VTAIL.n209 8.14595
R254 VTAIL.n24 VTAIL.n23 8.14595
R255 VTAIL.n150 VTAIL.n149 8.14595
R256 VTAIL.n88 VTAIL.n87 8.14595
R257 VTAIL.n206 VTAIL.n204 7.3702
R258 VTAIL.n20 VTAIL.n18 7.3702
R259 VTAIL.n146 VTAIL.n144 7.3702
R260 VTAIL.n84 VTAIL.n82 7.3702
R261 VTAIL.n209 VTAIL.n204 5.81868
R262 VTAIL.n23 VTAIL.n18 5.81868
R263 VTAIL.n149 VTAIL.n144 5.81868
R264 VTAIL.n87 VTAIL.n82 5.81868
R265 VTAIL.n210 VTAIL.n202 5.04292
R266 VTAIL.n246 VTAIL.n186 5.04292
R267 VTAIL.n24 VTAIL.n16 5.04292
R268 VTAIL.n60 VTAIL.n0 5.04292
R269 VTAIL.n184 VTAIL.n124 5.04292
R270 VTAIL.n150 VTAIL.n142 5.04292
R271 VTAIL.n122 VTAIL.n62 5.04292
R272 VTAIL.n88 VTAIL.n80 5.04292
R273 VTAIL.n214 VTAIL.n213 4.26717
R274 VTAIL.n244 VTAIL.n243 4.26717
R275 VTAIL.n28 VTAIL.n27 4.26717
R276 VTAIL.n58 VTAIL.n57 4.26717
R277 VTAIL.n182 VTAIL.n181 4.26717
R278 VTAIL.n154 VTAIL.n153 4.26717
R279 VTAIL.n120 VTAIL.n119 4.26717
R280 VTAIL.n92 VTAIL.n91 4.26717
R281 VTAIL.n217 VTAIL.n200 3.49141
R282 VTAIL.n240 VTAIL.n188 3.49141
R283 VTAIL.n31 VTAIL.n14 3.49141
R284 VTAIL.n54 VTAIL.n2 3.49141
R285 VTAIL.n178 VTAIL.n126 3.49141
R286 VTAIL.n157 VTAIL.n140 3.49141
R287 VTAIL.n116 VTAIL.n64 3.49141
R288 VTAIL.n95 VTAIL.n78 3.49141
R289 VTAIL.n205 VTAIL.n203 2.84303
R290 VTAIL.n19 VTAIL.n17 2.84303
R291 VTAIL.n145 VTAIL.n143 2.84303
R292 VTAIL.n83 VTAIL.n81 2.84303
R293 VTAIL.n218 VTAIL.n198 2.71565
R294 VTAIL.n239 VTAIL.n190 2.71565
R295 VTAIL.n32 VTAIL.n12 2.71565
R296 VTAIL.n53 VTAIL.n4 2.71565
R297 VTAIL.n177 VTAIL.n128 2.71565
R298 VTAIL.n158 VTAIL.n138 2.71565
R299 VTAIL.n115 VTAIL.n66 2.71565
R300 VTAIL.n96 VTAIL.n76 2.71565
R301 VTAIL.n223 VTAIL.n221 1.93989
R302 VTAIL.n236 VTAIL.n235 1.93989
R303 VTAIL.n37 VTAIL.n35 1.93989
R304 VTAIL.n50 VTAIL.n49 1.93989
R305 VTAIL.n174 VTAIL.n173 1.93989
R306 VTAIL.n162 VTAIL.n161 1.93989
R307 VTAIL.n112 VTAIL.n111 1.93989
R308 VTAIL.n100 VTAIL.n99 1.93989
R309 VTAIL.n185 VTAIL.n123 1.22895
R310 VTAIL.n222 VTAIL.n196 1.16414
R311 VTAIL.n232 VTAIL.n192 1.16414
R312 VTAIL.n36 VTAIL.n10 1.16414
R313 VTAIL.n46 VTAIL.n6 1.16414
R314 VTAIL.n170 VTAIL.n130 1.16414
R315 VTAIL.n165 VTAIL.n135 1.16414
R316 VTAIL.n108 VTAIL.n68 1.16414
R317 VTAIL.n103 VTAIL.n73 1.16414
R318 VTAIL VTAIL.n61 0.907828
R319 VTAIL.n228 VTAIL.n227 0.388379
R320 VTAIL.n231 VTAIL.n194 0.388379
R321 VTAIL.n42 VTAIL.n41 0.388379
R322 VTAIL.n45 VTAIL.n8 0.388379
R323 VTAIL.n169 VTAIL.n132 0.388379
R324 VTAIL.n166 VTAIL.n134 0.388379
R325 VTAIL.n107 VTAIL.n70 0.388379
R326 VTAIL.n104 VTAIL.n72 0.388379
R327 VTAIL VTAIL.n247 0.321621
R328 VTAIL.n211 VTAIL.n203 0.155672
R329 VTAIL.n212 VTAIL.n211 0.155672
R330 VTAIL.n212 VTAIL.n199 0.155672
R331 VTAIL.n219 VTAIL.n199 0.155672
R332 VTAIL.n220 VTAIL.n219 0.155672
R333 VTAIL.n220 VTAIL.n195 0.155672
R334 VTAIL.n229 VTAIL.n195 0.155672
R335 VTAIL.n230 VTAIL.n229 0.155672
R336 VTAIL.n230 VTAIL.n191 0.155672
R337 VTAIL.n237 VTAIL.n191 0.155672
R338 VTAIL.n238 VTAIL.n237 0.155672
R339 VTAIL.n238 VTAIL.n187 0.155672
R340 VTAIL.n245 VTAIL.n187 0.155672
R341 VTAIL.n25 VTAIL.n17 0.155672
R342 VTAIL.n26 VTAIL.n25 0.155672
R343 VTAIL.n26 VTAIL.n13 0.155672
R344 VTAIL.n33 VTAIL.n13 0.155672
R345 VTAIL.n34 VTAIL.n33 0.155672
R346 VTAIL.n34 VTAIL.n9 0.155672
R347 VTAIL.n43 VTAIL.n9 0.155672
R348 VTAIL.n44 VTAIL.n43 0.155672
R349 VTAIL.n44 VTAIL.n5 0.155672
R350 VTAIL.n51 VTAIL.n5 0.155672
R351 VTAIL.n52 VTAIL.n51 0.155672
R352 VTAIL.n52 VTAIL.n1 0.155672
R353 VTAIL.n59 VTAIL.n1 0.155672
R354 VTAIL.n183 VTAIL.n125 0.155672
R355 VTAIL.n176 VTAIL.n125 0.155672
R356 VTAIL.n176 VTAIL.n175 0.155672
R357 VTAIL.n175 VTAIL.n129 0.155672
R358 VTAIL.n168 VTAIL.n129 0.155672
R359 VTAIL.n168 VTAIL.n167 0.155672
R360 VTAIL.n167 VTAIL.n133 0.155672
R361 VTAIL.n160 VTAIL.n133 0.155672
R362 VTAIL.n160 VTAIL.n159 0.155672
R363 VTAIL.n159 VTAIL.n139 0.155672
R364 VTAIL.n152 VTAIL.n139 0.155672
R365 VTAIL.n152 VTAIL.n151 0.155672
R366 VTAIL.n151 VTAIL.n143 0.155672
R367 VTAIL.n121 VTAIL.n63 0.155672
R368 VTAIL.n114 VTAIL.n63 0.155672
R369 VTAIL.n114 VTAIL.n113 0.155672
R370 VTAIL.n113 VTAIL.n67 0.155672
R371 VTAIL.n106 VTAIL.n67 0.155672
R372 VTAIL.n106 VTAIL.n105 0.155672
R373 VTAIL.n105 VTAIL.n71 0.155672
R374 VTAIL.n98 VTAIL.n71 0.155672
R375 VTAIL.n98 VTAIL.n97 0.155672
R376 VTAIL.n97 VTAIL.n77 0.155672
R377 VTAIL.n90 VTAIL.n77 0.155672
R378 VTAIL.n90 VTAIL.n89 0.155672
R379 VTAIL.n89 VTAIL.n81 0.155672
R380 VDD1.n56 VDD1.n0 289.615
R381 VDD1.n117 VDD1.n61 289.615
R382 VDD1.n57 VDD1.n56 185
R383 VDD1.n55 VDD1.n54 185
R384 VDD1.n4 VDD1.n3 185
R385 VDD1.n49 VDD1.n48 185
R386 VDD1.n47 VDD1.n46 185
R387 VDD1.n8 VDD1.n7 185
R388 VDD1.n12 VDD1.n10 185
R389 VDD1.n41 VDD1.n40 185
R390 VDD1.n39 VDD1.n38 185
R391 VDD1.n14 VDD1.n13 185
R392 VDD1.n33 VDD1.n32 185
R393 VDD1.n31 VDD1.n30 185
R394 VDD1.n18 VDD1.n17 185
R395 VDD1.n25 VDD1.n24 185
R396 VDD1.n23 VDD1.n22 185
R397 VDD1.n82 VDD1.n81 185
R398 VDD1.n84 VDD1.n83 185
R399 VDD1.n77 VDD1.n76 185
R400 VDD1.n90 VDD1.n89 185
R401 VDD1.n92 VDD1.n91 185
R402 VDD1.n73 VDD1.n72 185
R403 VDD1.n99 VDD1.n98 185
R404 VDD1.n100 VDD1.n71 185
R405 VDD1.n102 VDD1.n101 185
R406 VDD1.n69 VDD1.n68 185
R407 VDD1.n108 VDD1.n107 185
R408 VDD1.n110 VDD1.n109 185
R409 VDD1.n65 VDD1.n64 185
R410 VDD1.n116 VDD1.n115 185
R411 VDD1.n118 VDD1.n117 185
R412 VDD1.n21 VDD1.t1 149.524
R413 VDD1.n80 VDD1.t0 149.524
R414 VDD1.n56 VDD1.n55 104.615
R415 VDD1.n55 VDD1.n3 104.615
R416 VDD1.n48 VDD1.n3 104.615
R417 VDD1.n48 VDD1.n47 104.615
R418 VDD1.n47 VDD1.n7 104.615
R419 VDD1.n12 VDD1.n7 104.615
R420 VDD1.n40 VDD1.n12 104.615
R421 VDD1.n40 VDD1.n39 104.615
R422 VDD1.n39 VDD1.n13 104.615
R423 VDD1.n32 VDD1.n13 104.615
R424 VDD1.n32 VDD1.n31 104.615
R425 VDD1.n31 VDD1.n17 104.615
R426 VDD1.n24 VDD1.n17 104.615
R427 VDD1.n24 VDD1.n23 104.615
R428 VDD1.n83 VDD1.n82 104.615
R429 VDD1.n83 VDD1.n76 104.615
R430 VDD1.n90 VDD1.n76 104.615
R431 VDD1.n91 VDD1.n90 104.615
R432 VDD1.n91 VDD1.n72 104.615
R433 VDD1.n99 VDD1.n72 104.615
R434 VDD1.n100 VDD1.n99 104.615
R435 VDD1.n101 VDD1.n100 104.615
R436 VDD1.n101 VDD1.n68 104.615
R437 VDD1.n108 VDD1.n68 104.615
R438 VDD1.n109 VDD1.n108 104.615
R439 VDD1.n109 VDD1.n64 104.615
R440 VDD1.n116 VDD1.n64 104.615
R441 VDD1.n117 VDD1.n116 104.615
R442 VDD1 VDD1.n121 86.2898
R443 VDD1.n23 VDD1.t1 52.3082
R444 VDD1.n82 VDD1.t0 52.3082
R445 VDD1 VDD1.n60 49.3016
R446 VDD1.n10 VDD1.n8 13.1884
R447 VDD1.n102 VDD1.n69 13.1884
R448 VDD1.n46 VDD1.n45 12.8005
R449 VDD1.n42 VDD1.n41 12.8005
R450 VDD1.n103 VDD1.n71 12.8005
R451 VDD1.n107 VDD1.n106 12.8005
R452 VDD1.n49 VDD1.n6 12.0247
R453 VDD1.n38 VDD1.n11 12.0247
R454 VDD1.n98 VDD1.n97 12.0247
R455 VDD1.n110 VDD1.n67 12.0247
R456 VDD1.n50 VDD1.n4 11.249
R457 VDD1.n37 VDD1.n14 11.249
R458 VDD1.n96 VDD1.n73 11.249
R459 VDD1.n111 VDD1.n65 11.249
R460 VDD1.n54 VDD1.n53 10.4732
R461 VDD1.n34 VDD1.n33 10.4732
R462 VDD1.n93 VDD1.n92 10.4732
R463 VDD1.n115 VDD1.n114 10.4732
R464 VDD1.n22 VDD1.n21 10.2747
R465 VDD1.n81 VDD1.n80 10.2747
R466 VDD1.n57 VDD1.n2 9.69747
R467 VDD1.n30 VDD1.n16 9.69747
R468 VDD1.n89 VDD1.n75 9.69747
R469 VDD1.n118 VDD1.n63 9.69747
R470 VDD1.n60 VDD1.n59 9.45567
R471 VDD1.n121 VDD1.n120 9.45567
R472 VDD1.n20 VDD1.n19 9.3005
R473 VDD1.n27 VDD1.n26 9.3005
R474 VDD1.n29 VDD1.n28 9.3005
R475 VDD1.n16 VDD1.n15 9.3005
R476 VDD1.n35 VDD1.n34 9.3005
R477 VDD1.n37 VDD1.n36 9.3005
R478 VDD1.n11 VDD1.n9 9.3005
R479 VDD1.n43 VDD1.n42 9.3005
R480 VDD1.n59 VDD1.n58 9.3005
R481 VDD1.n2 VDD1.n1 9.3005
R482 VDD1.n53 VDD1.n52 9.3005
R483 VDD1.n51 VDD1.n50 9.3005
R484 VDD1.n6 VDD1.n5 9.3005
R485 VDD1.n45 VDD1.n44 9.3005
R486 VDD1.n120 VDD1.n119 9.3005
R487 VDD1.n63 VDD1.n62 9.3005
R488 VDD1.n114 VDD1.n113 9.3005
R489 VDD1.n112 VDD1.n111 9.3005
R490 VDD1.n67 VDD1.n66 9.3005
R491 VDD1.n106 VDD1.n105 9.3005
R492 VDD1.n79 VDD1.n78 9.3005
R493 VDD1.n86 VDD1.n85 9.3005
R494 VDD1.n88 VDD1.n87 9.3005
R495 VDD1.n75 VDD1.n74 9.3005
R496 VDD1.n94 VDD1.n93 9.3005
R497 VDD1.n96 VDD1.n95 9.3005
R498 VDD1.n97 VDD1.n70 9.3005
R499 VDD1.n104 VDD1.n103 9.3005
R500 VDD1.n58 VDD1.n0 8.92171
R501 VDD1.n29 VDD1.n18 8.92171
R502 VDD1.n88 VDD1.n77 8.92171
R503 VDD1.n119 VDD1.n61 8.92171
R504 VDD1.n26 VDD1.n25 8.14595
R505 VDD1.n85 VDD1.n84 8.14595
R506 VDD1.n22 VDD1.n20 7.3702
R507 VDD1.n81 VDD1.n79 7.3702
R508 VDD1.n25 VDD1.n20 5.81868
R509 VDD1.n84 VDD1.n79 5.81868
R510 VDD1.n60 VDD1.n0 5.04292
R511 VDD1.n26 VDD1.n18 5.04292
R512 VDD1.n85 VDD1.n77 5.04292
R513 VDD1.n121 VDD1.n61 5.04292
R514 VDD1.n58 VDD1.n57 4.26717
R515 VDD1.n30 VDD1.n29 4.26717
R516 VDD1.n89 VDD1.n88 4.26717
R517 VDD1.n119 VDD1.n118 4.26717
R518 VDD1.n54 VDD1.n2 3.49141
R519 VDD1.n33 VDD1.n16 3.49141
R520 VDD1.n92 VDD1.n75 3.49141
R521 VDD1.n115 VDD1.n63 3.49141
R522 VDD1.n21 VDD1.n19 2.84303
R523 VDD1.n80 VDD1.n78 2.84303
R524 VDD1.n53 VDD1.n4 2.71565
R525 VDD1.n34 VDD1.n14 2.71565
R526 VDD1.n93 VDD1.n73 2.71565
R527 VDD1.n114 VDD1.n65 2.71565
R528 VDD1.n50 VDD1.n49 1.93989
R529 VDD1.n38 VDD1.n37 1.93989
R530 VDD1.n98 VDD1.n96 1.93989
R531 VDD1.n111 VDD1.n110 1.93989
R532 VDD1.n46 VDD1.n6 1.16414
R533 VDD1.n41 VDD1.n11 1.16414
R534 VDD1.n97 VDD1.n71 1.16414
R535 VDD1.n107 VDD1.n67 1.16414
R536 VDD1.n45 VDD1.n8 0.388379
R537 VDD1.n42 VDD1.n10 0.388379
R538 VDD1.n103 VDD1.n102 0.388379
R539 VDD1.n106 VDD1.n69 0.388379
R540 VDD1.n59 VDD1.n1 0.155672
R541 VDD1.n52 VDD1.n1 0.155672
R542 VDD1.n52 VDD1.n51 0.155672
R543 VDD1.n51 VDD1.n5 0.155672
R544 VDD1.n44 VDD1.n5 0.155672
R545 VDD1.n44 VDD1.n43 0.155672
R546 VDD1.n43 VDD1.n9 0.155672
R547 VDD1.n36 VDD1.n9 0.155672
R548 VDD1.n36 VDD1.n35 0.155672
R549 VDD1.n35 VDD1.n15 0.155672
R550 VDD1.n28 VDD1.n15 0.155672
R551 VDD1.n28 VDD1.n27 0.155672
R552 VDD1.n27 VDD1.n19 0.155672
R553 VDD1.n86 VDD1.n78 0.155672
R554 VDD1.n87 VDD1.n86 0.155672
R555 VDD1.n87 VDD1.n74 0.155672
R556 VDD1.n94 VDD1.n74 0.155672
R557 VDD1.n95 VDD1.n94 0.155672
R558 VDD1.n95 VDD1.n70 0.155672
R559 VDD1.n104 VDD1.n70 0.155672
R560 VDD1.n105 VDD1.n104 0.155672
R561 VDD1.n105 VDD1.n66 0.155672
R562 VDD1.n112 VDD1.n66 0.155672
R563 VDD1.n113 VDD1.n112 0.155672
R564 VDD1.n113 VDD1.n62 0.155672
R565 VDD1.n120 VDD1.n62 0.155672
R566 B.n428 B.n85 585
R567 B.n85 B.n36 585
R568 B.n430 B.n429 585
R569 B.n432 B.n84 585
R570 B.n435 B.n434 585
R571 B.n436 B.n83 585
R572 B.n438 B.n437 585
R573 B.n440 B.n82 585
R574 B.n443 B.n442 585
R575 B.n444 B.n81 585
R576 B.n446 B.n445 585
R577 B.n448 B.n80 585
R578 B.n451 B.n450 585
R579 B.n452 B.n79 585
R580 B.n454 B.n453 585
R581 B.n456 B.n78 585
R582 B.n459 B.n458 585
R583 B.n460 B.n77 585
R584 B.n462 B.n461 585
R585 B.n464 B.n76 585
R586 B.n467 B.n466 585
R587 B.n468 B.n75 585
R588 B.n470 B.n469 585
R589 B.n472 B.n74 585
R590 B.n475 B.n474 585
R591 B.n476 B.n73 585
R592 B.n478 B.n477 585
R593 B.n480 B.n72 585
R594 B.n483 B.n482 585
R595 B.n484 B.n71 585
R596 B.n486 B.n485 585
R597 B.n488 B.n70 585
R598 B.n491 B.n490 585
R599 B.n492 B.n69 585
R600 B.n494 B.n493 585
R601 B.n496 B.n68 585
R602 B.n499 B.n498 585
R603 B.n500 B.n67 585
R604 B.n502 B.n501 585
R605 B.n504 B.n66 585
R606 B.n507 B.n506 585
R607 B.n509 B.n63 585
R608 B.n511 B.n510 585
R609 B.n513 B.n62 585
R610 B.n516 B.n515 585
R611 B.n517 B.n61 585
R612 B.n519 B.n518 585
R613 B.n521 B.n60 585
R614 B.n524 B.n523 585
R615 B.n525 B.n57 585
R616 B.n528 B.n527 585
R617 B.n530 B.n56 585
R618 B.n533 B.n532 585
R619 B.n534 B.n55 585
R620 B.n536 B.n535 585
R621 B.n538 B.n54 585
R622 B.n541 B.n540 585
R623 B.n542 B.n53 585
R624 B.n544 B.n543 585
R625 B.n546 B.n52 585
R626 B.n549 B.n548 585
R627 B.n550 B.n51 585
R628 B.n552 B.n551 585
R629 B.n554 B.n50 585
R630 B.n557 B.n556 585
R631 B.n558 B.n49 585
R632 B.n560 B.n559 585
R633 B.n562 B.n48 585
R634 B.n565 B.n564 585
R635 B.n566 B.n47 585
R636 B.n568 B.n567 585
R637 B.n570 B.n46 585
R638 B.n573 B.n572 585
R639 B.n574 B.n45 585
R640 B.n576 B.n575 585
R641 B.n578 B.n44 585
R642 B.n581 B.n580 585
R643 B.n582 B.n43 585
R644 B.n584 B.n583 585
R645 B.n586 B.n42 585
R646 B.n589 B.n588 585
R647 B.n590 B.n41 585
R648 B.n592 B.n591 585
R649 B.n594 B.n40 585
R650 B.n597 B.n596 585
R651 B.n598 B.n39 585
R652 B.n600 B.n599 585
R653 B.n602 B.n38 585
R654 B.n605 B.n604 585
R655 B.n606 B.n37 585
R656 B.n427 B.n35 585
R657 B.n609 B.n35 585
R658 B.n426 B.n34 585
R659 B.n610 B.n34 585
R660 B.n425 B.n33 585
R661 B.n611 B.n33 585
R662 B.n424 B.n423 585
R663 B.n423 B.n29 585
R664 B.n422 B.n28 585
R665 B.n617 B.n28 585
R666 B.n421 B.n27 585
R667 B.n618 B.n27 585
R668 B.n420 B.n26 585
R669 B.n619 B.n26 585
R670 B.n419 B.n418 585
R671 B.n418 B.n22 585
R672 B.n417 B.n21 585
R673 B.n625 B.n21 585
R674 B.n416 B.n20 585
R675 B.n626 B.n20 585
R676 B.n415 B.n19 585
R677 B.n627 B.n19 585
R678 B.n414 B.n413 585
R679 B.n413 B.n15 585
R680 B.n412 B.n14 585
R681 B.n633 B.n14 585
R682 B.n411 B.n13 585
R683 B.n634 B.n13 585
R684 B.n410 B.n12 585
R685 B.n635 B.n12 585
R686 B.n409 B.n408 585
R687 B.n408 B.n407 585
R688 B.n406 B.n405 585
R689 B.n406 B.n8 585
R690 B.n404 B.n7 585
R691 B.n642 B.n7 585
R692 B.n403 B.n6 585
R693 B.n643 B.n6 585
R694 B.n402 B.n5 585
R695 B.n644 B.n5 585
R696 B.n401 B.n400 585
R697 B.n400 B.n4 585
R698 B.n399 B.n86 585
R699 B.n399 B.n398 585
R700 B.n389 B.n87 585
R701 B.n88 B.n87 585
R702 B.n391 B.n390 585
R703 B.n392 B.n391 585
R704 B.n388 B.n93 585
R705 B.n93 B.n92 585
R706 B.n387 B.n386 585
R707 B.n386 B.n385 585
R708 B.n95 B.n94 585
R709 B.n96 B.n95 585
R710 B.n378 B.n377 585
R711 B.n379 B.n378 585
R712 B.n376 B.n101 585
R713 B.n101 B.n100 585
R714 B.n375 B.n374 585
R715 B.n374 B.n373 585
R716 B.n103 B.n102 585
R717 B.n104 B.n103 585
R718 B.n366 B.n365 585
R719 B.n367 B.n366 585
R720 B.n364 B.n108 585
R721 B.n112 B.n108 585
R722 B.n363 B.n362 585
R723 B.n362 B.n361 585
R724 B.n110 B.n109 585
R725 B.n111 B.n110 585
R726 B.n354 B.n353 585
R727 B.n355 B.n354 585
R728 B.n352 B.n117 585
R729 B.n117 B.n116 585
R730 B.n351 B.n350 585
R731 B.n350 B.n349 585
R732 B.n346 B.n121 585
R733 B.n345 B.n344 585
R734 B.n342 B.n122 585
R735 B.n342 B.n120 585
R736 B.n341 B.n340 585
R737 B.n339 B.n338 585
R738 B.n337 B.n124 585
R739 B.n335 B.n334 585
R740 B.n333 B.n125 585
R741 B.n332 B.n331 585
R742 B.n329 B.n126 585
R743 B.n327 B.n326 585
R744 B.n325 B.n127 585
R745 B.n324 B.n323 585
R746 B.n321 B.n128 585
R747 B.n319 B.n318 585
R748 B.n317 B.n129 585
R749 B.n316 B.n315 585
R750 B.n313 B.n130 585
R751 B.n311 B.n310 585
R752 B.n309 B.n131 585
R753 B.n308 B.n307 585
R754 B.n305 B.n132 585
R755 B.n303 B.n302 585
R756 B.n301 B.n133 585
R757 B.n300 B.n299 585
R758 B.n297 B.n134 585
R759 B.n295 B.n294 585
R760 B.n293 B.n135 585
R761 B.n292 B.n291 585
R762 B.n289 B.n136 585
R763 B.n287 B.n286 585
R764 B.n285 B.n137 585
R765 B.n284 B.n283 585
R766 B.n281 B.n138 585
R767 B.n279 B.n278 585
R768 B.n277 B.n139 585
R769 B.n276 B.n275 585
R770 B.n273 B.n140 585
R771 B.n271 B.n270 585
R772 B.n269 B.n141 585
R773 B.n267 B.n266 585
R774 B.n264 B.n144 585
R775 B.n262 B.n261 585
R776 B.n260 B.n145 585
R777 B.n259 B.n258 585
R778 B.n256 B.n146 585
R779 B.n254 B.n253 585
R780 B.n252 B.n147 585
R781 B.n251 B.n250 585
R782 B.n248 B.n247 585
R783 B.n246 B.n245 585
R784 B.n244 B.n152 585
R785 B.n242 B.n241 585
R786 B.n240 B.n153 585
R787 B.n239 B.n238 585
R788 B.n236 B.n154 585
R789 B.n234 B.n233 585
R790 B.n232 B.n155 585
R791 B.n231 B.n230 585
R792 B.n228 B.n156 585
R793 B.n226 B.n225 585
R794 B.n224 B.n157 585
R795 B.n223 B.n222 585
R796 B.n220 B.n158 585
R797 B.n218 B.n217 585
R798 B.n216 B.n159 585
R799 B.n215 B.n214 585
R800 B.n212 B.n160 585
R801 B.n210 B.n209 585
R802 B.n208 B.n161 585
R803 B.n207 B.n206 585
R804 B.n204 B.n162 585
R805 B.n202 B.n201 585
R806 B.n200 B.n163 585
R807 B.n199 B.n198 585
R808 B.n196 B.n164 585
R809 B.n194 B.n193 585
R810 B.n192 B.n165 585
R811 B.n191 B.n190 585
R812 B.n188 B.n166 585
R813 B.n186 B.n185 585
R814 B.n184 B.n167 585
R815 B.n183 B.n182 585
R816 B.n180 B.n168 585
R817 B.n178 B.n177 585
R818 B.n176 B.n169 585
R819 B.n175 B.n174 585
R820 B.n172 B.n170 585
R821 B.n119 B.n118 585
R822 B.n348 B.n347 585
R823 B.n349 B.n348 585
R824 B.n115 B.n114 585
R825 B.n116 B.n115 585
R826 B.n357 B.n356 585
R827 B.n356 B.n355 585
R828 B.n358 B.n113 585
R829 B.n113 B.n111 585
R830 B.n360 B.n359 585
R831 B.n361 B.n360 585
R832 B.n107 B.n106 585
R833 B.n112 B.n107 585
R834 B.n369 B.n368 585
R835 B.n368 B.n367 585
R836 B.n370 B.n105 585
R837 B.n105 B.n104 585
R838 B.n372 B.n371 585
R839 B.n373 B.n372 585
R840 B.n99 B.n98 585
R841 B.n100 B.n99 585
R842 B.n381 B.n380 585
R843 B.n380 B.n379 585
R844 B.n382 B.n97 585
R845 B.n97 B.n96 585
R846 B.n384 B.n383 585
R847 B.n385 B.n384 585
R848 B.n91 B.n90 585
R849 B.n92 B.n91 585
R850 B.n394 B.n393 585
R851 B.n393 B.n392 585
R852 B.n395 B.n89 585
R853 B.n89 B.n88 585
R854 B.n397 B.n396 585
R855 B.n398 B.n397 585
R856 B.n3 B.n0 585
R857 B.n4 B.n3 585
R858 B.n641 B.n1 585
R859 B.n642 B.n641 585
R860 B.n640 B.n639 585
R861 B.n640 B.n8 585
R862 B.n638 B.n9 585
R863 B.n407 B.n9 585
R864 B.n637 B.n636 585
R865 B.n636 B.n635 585
R866 B.n11 B.n10 585
R867 B.n634 B.n11 585
R868 B.n632 B.n631 585
R869 B.n633 B.n632 585
R870 B.n630 B.n16 585
R871 B.n16 B.n15 585
R872 B.n629 B.n628 585
R873 B.n628 B.n627 585
R874 B.n18 B.n17 585
R875 B.n626 B.n18 585
R876 B.n624 B.n623 585
R877 B.n625 B.n624 585
R878 B.n622 B.n23 585
R879 B.n23 B.n22 585
R880 B.n621 B.n620 585
R881 B.n620 B.n619 585
R882 B.n25 B.n24 585
R883 B.n618 B.n25 585
R884 B.n616 B.n615 585
R885 B.n617 B.n616 585
R886 B.n614 B.n30 585
R887 B.n30 B.n29 585
R888 B.n613 B.n612 585
R889 B.n612 B.n611 585
R890 B.n32 B.n31 585
R891 B.n610 B.n32 585
R892 B.n608 B.n607 585
R893 B.n609 B.n608 585
R894 B.n645 B.n644 585
R895 B.n643 B.n2 585
R896 B.n608 B.n37 516.524
R897 B.n85 B.n35 516.524
R898 B.n350 B.n119 516.524
R899 B.n348 B.n121 516.524
R900 B.n58 B.t6 397.296
R901 B.n64 B.t13 397.296
R902 B.n148 B.t2 397.296
R903 B.n142 B.t10 397.296
R904 B.n64 B.t14 305.981
R905 B.n148 B.t5 305.981
R906 B.n58 B.t8 305.981
R907 B.n142 B.t12 305.981
R908 B.n65 B.t15 271.848
R909 B.n149 B.t4 271.848
R910 B.n59 B.t9 271.848
R911 B.n143 B.t11 271.848
R912 B.n431 B.n36 256.663
R913 B.n433 B.n36 256.663
R914 B.n439 B.n36 256.663
R915 B.n441 B.n36 256.663
R916 B.n447 B.n36 256.663
R917 B.n449 B.n36 256.663
R918 B.n455 B.n36 256.663
R919 B.n457 B.n36 256.663
R920 B.n463 B.n36 256.663
R921 B.n465 B.n36 256.663
R922 B.n471 B.n36 256.663
R923 B.n473 B.n36 256.663
R924 B.n479 B.n36 256.663
R925 B.n481 B.n36 256.663
R926 B.n487 B.n36 256.663
R927 B.n489 B.n36 256.663
R928 B.n495 B.n36 256.663
R929 B.n497 B.n36 256.663
R930 B.n503 B.n36 256.663
R931 B.n505 B.n36 256.663
R932 B.n512 B.n36 256.663
R933 B.n514 B.n36 256.663
R934 B.n520 B.n36 256.663
R935 B.n522 B.n36 256.663
R936 B.n529 B.n36 256.663
R937 B.n531 B.n36 256.663
R938 B.n537 B.n36 256.663
R939 B.n539 B.n36 256.663
R940 B.n545 B.n36 256.663
R941 B.n547 B.n36 256.663
R942 B.n553 B.n36 256.663
R943 B.n555 B.n36 256.663
R944 B.n561 B.n36 256.663
R945 B.n563 B.n36 256.663
R946 B.n569 B.n36 256.663
R947 B.n571 B.n36 256.663
R948 B.n577 B.n36 256.663
R949 B.n579 B.n36 256.663
R950 B.n585 B.n36 256.663
R951 B.n587 B.n36 256.663
R952 B.n593 B.n36 256.663
R953 B.n595 B.n36 256.663
R954 B.n601 B.n36 256.663
R955 B.n603 B.n36 256.663
R956 B.n343 B.n120 256.663
R957 B.n123 B.n120 256.663
R958 B.n336 B.n120 256.663
R959 B.n330 B.n120 256.663
R960 B.n328 B.n120 256.663
R961 B.n322 B.n120 256.663
R962 B.n320 B.n120 256.663
R963 B.n314 B.n120 256.663
R964 B.n312 B.n120 256.663
R965 B.n306 B.n120 256.663
R966 B.n304 B.n120 256.663
R967 B.n298 B.n120 256.663
R968 B.n296 B.n120 256.663
R969 B.n290 B.n120 256.663
R970 B.n288 B.n120 256.663
R971 B.n282 B.n120 256.663
R972 B.n280 B.n120 256.663
R973 B.n274 B.n120 256.663
R974 B.n272 B.n120 256.663
R975 B.n265 B.n120 256.663
R976 B.n263 B.n120 256.663
R977 B.n257 B.n120 256.663
R978 B.n255 B.n120 256.663
R979 B.n249 B.n120 256.663
R980 B.n151 B.n120 256.663
R981 B.n243 B.n120 256.663
R982 B.n237 B.n120 256.663
R983 B.n235 B.n120 256.663
R984 B.n229 B.n120 256.663
R985 B.n227 B.n120 256.663
R986 B.n221 B.n120 256.663
R987 B.n219 B.n120 256.663
R988 B.n213 B.n120 256.663
R989 B.n211 B.n120 256.663
R990 B.n205 B.n120 256.663
R991 B.n203 B.n120 256.663
R992 B.n197 B.n120 256.663
R993 B.n195 B.n120 256.663
R994 B.n189 B.n120 256.663
R995 B.n187 B.n120 256.663
R996 B.n181 B.n120 256.663
R997 B.n179 B.n120 256.663
R998 B.n173 B.n120 256.663
R999 B.n171 B.n120 256.663
R1000 B.n647 B.n646 256.663
R1001 B.n604 B.n602 163.367
R1002 B.n600 B.n39 163.367
R1003 B.n596 B.n594 163.367
R1004 B.n592 B.n41 163.367
R1005 B.n588 B.n586 163.367
R1006 B.n584 B.n43 163.367
R1007 B.n580 B.n578 163.367
R1008 B.n576 B.n45 163.367
R1009 B.n572 B.n570 163.367
R1010 B.n568 B.n47 163.367
R1011 B.n564 B.n562 163.367
R1012 B.n560 B.n49 163.367
R1013 B.n556 B.n554 163.367
R1014 B.n552 B.n51 163.367
R1015 B.n548 B.n546 163.367
R1016 B.n544 B.n53 163.367
R1017 B.n540 B.n538 163.367
R1018 B.n536 B.n55 163.367
R1019 B.n532 B.n530 163.367
R1020 B.n528 B.n57 163.367
R1021 B.n523 B.n521 163.367
R1022 B.n519 B.n61 163.367
R1023 B.n515 B.n513 163.367
R1024 B.n511 B.n63 163.367
R1025 B.n506 B.n504 163.367
R1026 B.n502 B.n67 163.367
R1027 B.n498 B.n496 163.367
R1028 B.n494 B.n69 163.367
R1029 B.n490 B.n488 163.367
R1030 B.n486 B.n71 163.367
R1031 B.n482 B.n480 163.367
R1032 B.n478 B.n73 163.367
R1033 B.n474 B.n472 163.367
R1034 B.n470 B.n75 163.367
R1035 B.n466 B.n464 163.367
R1036 B.n462 B.n77 163.367
R1037 B.n458 B.n456 163.367
R1038 B.n454 B.n79 163.367
R1039 B.n450 B.n448 163.367
R1040 B.n446 B.n81 163.367
R1041 B.n442 B.n440 163.367
R1042 B.n438 B.n83 163.367
R1043 B.n434 B.n432 163.367
R1044 B.n430 B.n85 163.367
R1045 B.n350 B.n117 163.367
R1046 B.n354 B.n117 163.367
R1047 B.n354 B.n110 163.367
R1048 B.n362 B.n110 163.367
R1049 B.n362 B.n108 163.367
R1050 B.n366 B.n108 163.367
R1051 B.n366 B.n103 163.367
R1052 B.n374 B.n103 163.367
R1053 B.n374 B.n101 163.367
R1054 B.n378 B.n101 163.367
R1055 B.n378 B.n95 163.367
R1056 B.n386 B.n95 163.367
R1057 B.n386 B.n93 163.367
R1058 B.n391 B.n93 163.367
R1059 B.n391 B.n87 163.367
R1060 B.n399 B.n87 163.367
R1061 B.n400 B.n399 163.367
R1062 B.n400 B.n5 163.367
R1063 B.n6 B.n5 163.367
R1064 B.n7 B.n6 163.367
R1065 B.n406 B.n7 163.367
R1066 B.n408 B.n406 163.367
R1067 B.n408 B.n12 163.367
R1068 B.n13 B.n12 163.367
R1069 B.n14 B.n13 163.367
R1070 B.n413 B.n14 163.367
R1071 B.n413 B.n19 163.367
R1072 B.n20 B.n19 163.367
R1073 B.n21 B.n20 163.367
R1074 B.n418 B.n21 163.367
R1075 B.n418 B.n26 163.367
R1076 B.n27 B.n26 163.367
R1077 B.n28 B.n27 163.367
R1078 B.n423 B.n28 163.367
R1079 B.n423 B.n33 163.367
R1080 B.n34 B.n33 163.367
R1081 B.n35 B.n34 163.367
R1082 B.n344 B.n342 163.367
R1083 B.n342 B.n341 163.367
R1084 B.n338 B.n337 163.367
R1085 B.n335 B.n125 163.367
R1086 B.n331 B.n329 163.367
R1087 B.n327 B.n127 163.367
R1088 B.n323 B.n321 163.367
R1089 B.n319 B.n129 163.367
R1090 B.n315 B.n313 163.367
R1091 B.n311 B.n131 163.367
R1092 B.n307 B.n305 163.367
R1093 B.n303 B.n133 163.367
R1094 B.n299 B.n297 163.367
R1095 B.n295 B.n135 163.367
R1096 B.n291 B.n289 163.367
R1097 B.n287 B.n137 163.367
R1098 B.n283 B.n281 163.367
R1099 B.n279 B.n139 163.367
R1100 B.n275 B.n273 163.367
R1101 B.n271 B.n141 163.367
R1102 B.n266 B.n264 163.367
R1103 B.n262 B.n145 163.367
R1104 B.n258 B.n256 163.367
R1105 B.n254 B.n147 163.367
R1106 B.n250 B.n248 163.367
R1107 B.n245 B.n244 163.367
R1108 B.n242 B.n153 163.367
R1109 B.n238 B.n236 163.367
R1110 B.n234 B.n155 163.367
R1111 B.n230 B.n228 163.367
R1112 B.n226 B.n157 163.367
R1113 B.n222 B.n220 163.367
R1114 B.n218 B.n159 163.367
R1115 B.n214 B.n212 163.367
R1116 B.n210 B.n161 163.367
R1117 B.n206 B.n204 163.367
R1118 B.n202 B.n163 163.367
R1119 B.n198 B.n196 163.367
R1120 B.n194 B.n165 163.367
R1121 B.n190 B.n188 163.367
R1122 B.n186 B.n167 163.367
R1123 B.n182 B.n180 163.367
R1124 B.n178 B.n169 163.367
R1125 B.n174 B.n172 163.367
R1126 B.n348 B.n115 163.367
R1127 B.n356 B.n115 163.367
R1128 B.n356 B.n113 163.367
R1129 B.n360 B.n113 163.367
R1130 B.n360 B.n107 163.367
R1131 B.n368 B.n107 163.367
R1132 B.n368 B.n105 163.367
R1133 B.n372 B.n105 163.367
R1134 B.n372 B.n99 163.367
R1135 B.n380 B.n99 163.367
R1136 B.n380 B.n97 163.367
R1137 B.n384 B.n97 163.367
R1138 B.n384 B.n91 163.367
R1139 B.n393 B.n91 163.367
R1140 B.n393 B.n89 163.367
R1141 B.n397 B.n89 163.367
R1142 B.n397 B.n3 163.367
R1143 B.n645 B.n3 163.367
R1144 B.n641 B.n2 163.367
R1145 B.n641 B.n640 163.367
R1146 B.n640 B.n9 163.367
R1147 B.n636 B.n9 163.367
R1148 B.n636 B.n11 163.367
R1149 B.n632 B.n11 163.367
R1150 B.n632 B.n16 163.367
R1151 B.n628 B.n16 163.367
R1152 B.n628 B.n18 163.367
R1153 B.n624 B.n18 163.367
R1154 B.n624 B.n23 163.367
R1155 B.n620 B.n23 163.367
R1156 B.n620 B.n25 163.367
R1157 B.n616 B.n25 163.367
R1158 B.n616 B.n30 163.367
R1159 B.n612 B.n30 163.367
R1160 B.n612 B.n32 163.367
R1161 B.n608 B.n32 163.367
R1162 B.n349 B.n120 79.8206
R1163 B.n609 B.n36 79.8206
R1164 B.n603 B.n37 71.676
R1165 B.n602 B.n601 71.676
R1166 B.n595 B.n39 71.676
R1167 B.n594 B.n593 71.676
R1168 B.n587 B.n41 71.676
R1169 B.n586 B.n585 71.676
R1170 B.n579 B.n43 71.676
R1171 B.n578 B.n577 71.676
R1172 B.n571 B.n45 71.676
R1173 B.n570 B.n569 71.676
R1174 B.n563 B.n47 71.676
R1175 B.n562 B.n561 71.676
R1176 B.n555 B.n49 71.676
R1177 B.n554 B.n553 71.676
R1178 B.n547 B.n51 71.676
R1179 B.n546 B.n545 71.676
R1180 B.n539 B.n53 71.676
R1181 B.n538 B.n537 71.676
R1182 B.n531 B.n55 71.676
R1183 B.n530 B.n529 71.676
R1184 B.n522 B.n57 71.676
R1185 B.n521 B.n520 71.676
R1186 B.n514 B.n61 71.676
R1187 B.n513 B.n512 71.676
R1188 B.n505 B.n63 71.676
R1189 B.n504 B.n503 71.676
R1190 B.n497 B.n67 71.676
R1191 B.n496 B.n495 71.676
R1192 B.n489 B.n69 71.676
R1193 B.n488 B.n487 71.676
R1194 B.n481 B.n71 71.676
R1195 B.n480 B.n479 71.676
R1196 B.n473 B.n73 71.676
R1197 B.n472 B.n471 71.676
R1198 B.n465 B.n75 71.676
R1199 B.n464 B.n463 71.676
R1200 B.n457 B.n77 71.676
R1201 B.n456 B.n455 71.676
R1202 B.n449 B.n79 71.676
R1203 B.n448 B.n447 71.676
R1204 B.n441 B.n81 71.676
R1205 B.n440 B.n439 71.676
R1206 B.n433 B.n83 71.676
R1207 B.n432 B.n431 71.676
R1208 B.n431 B.n430 71.676
R1209 B.n434 B.n433 71.676
R1210 B.n439 B.n438 71.676
R1211 B.n442 B.n441 71.676
R1212 B.n447 B.n446 71.676
R1213 B.n450 B.n449 71.676
R1214 B.n455 B.n454 71.676
R1215 B.n458 B.n457 71.676
R1216 B.n463 B.n462 71.676
R1217 B.n466 B.n465 71.676
R1218 B.n471 B.n470 71.676
R1219 B.n474 B.n473 71.676
R1220 B.n479 B.n478 71.676
R1221 B.n482 B.n481 71.676
R1222 B.n487 B.n486 71.676
R1223 B.n490 B.n489 71.676
R1224 B.n495 B.n494 71.676
R1225 B.n498 B.n497 71.676
R1226 B.n503 B.n502 71.676
R1227 B.n506 B.n505 71.676
R1228 B.n512 B.n511 71.676
R1229 B.n515 B.n514 71.676
R1230 B.n520 B.n519 71.676
R1231 B.n523 B.n522 71.676
R1232 B.n529 B.n528 71.676
R1233 B.n532 B.n531 71.676
R1234 B.n537 B.n536 71.676
R1235 B.n540 B.n539 71.676
R1236 B.n545 B.n544 71.676
R1237 B.n548 B.n547 71.676
R1238 B.n553 B.n552 71.676
R1239 B.n556 B.n555 71.676
R1240 B.n561 B.n560 71.676
R1241 B.n564 B.n563 71.676
R1242 B.n569 B.n568 71.676
R1243 B.n572 B.n571 71.676
R1244 B.n577 B.n576 71.676
R1245 B.n580 B.n579 71.676
R1246 B.n585 B.n584 71.676
R1247 B.n588 B.n587 71.676
R1248 B.n593 B.n592 71.676
R1249 B.n596 B.n595 71.676
R1250 B.n601 B.n600 71.676
R1251 B.n604 B.n603 71.676
R1252 B.n343 B.n121 71.676
R1253 B.n341 B.n123 71.676
R1254 B.n337 B.n336 71.676
R1255 B.n330 B.n125 71.676
R1256 B.n329 B.n328 71.676
R1257 B.n322 B.n127 71.676
R1258 B.n321 B.n320 71.676
R1259 B.n314 B.n129 71.676
R1260 B.n313 B.n312 71.676
R1261 B.n306 B.n131 71.676
R1262 B.n305 B.n304 71.676
R1263 B.n298 B.n133 71.676
R1264 B.n297 B.n296 71.676
R1265 B.n290 B.n135 71.676
R1266 B.n289 B.n288 71.676
R1267 B.n282 B.n137 71.676
R1268 B.n281 B.n280 71.676
R1269 B.n274 B.n139 71.676
R1270 B.n273 B.n272 71.676
R1271 B.n265 B.n141 71.676
R1272 B.n264 B.n263 71.676
R1273 B.n257 B.n145 71.676
R1274 B.n256 B.n255 71.676
R1275 B.n249 B.n147 71.676
R1276 B.n248 B.n151 71.676
R1277 B.n244 B.n243 71.676
R1278 B.n237 B.n153 71.676
R1279 B.n236 B.n235 71.676
R1280 B.n229 B.n155 71.676
R1281 B.n228 B.n227 71.676
R1282 B.n221 B.n157 71.676
R1283 B.n220 B.n219 71.676
R1284 B.n213 B.n159 71.676
R1285 B.n212 B.n211 71.676
R1286 B.n205 B.n161 71.676
R1287 B.n204 B.n203 71.676
R1288 B.n197 B.n163 71.676
R1289 B.n196 B.n195 71.676
R1290 B.n189 B.n165 71.676
R1291 B.n188 B.n187 71.676
R1292 B.n181 B.n167 71.676
R1293 B.n180 B.n179 71.676
R1294 B.n173 B.n169 71.676
R1295 B.n172 B.n171 71.676
R1296 B.n344 B.n343 71.676
R1297 B.n338 B.n123 71.676
R1298 B.n336 B.n335 71.676
R1299 B.n331 B.n330 71.676
R1300 B.n328 B.n327 71.676
R1301 B.n323 B.n322 71.676
R1302 B.n320 B.n319 71.676
R1303 B.n315 B.n314 71.676
R1304 B.n312 B.n311 71.676
R1305 B.n307 B.n306 71.676
R1306 B.n304 B.n303 71.676
R1307 B.n299 B.n298 71.676
R1308 B.n296 B.n295 71.676
R1309 B.n291 B.n290 71.676
R1310 B.n288 B.n287 71.676
R1311 B.n283 B.n282 71.676
R1312 B.n280 B.n279 71.676
R1313 B.n275 B.n274 71.676
R1314 B.n272 B.n271 71.676
R1315 B.n266 B.n265 71.676
R1316 B.n263 B.n262 71.676
R1317 B.n258 B.n257 71.676
R1318 B.n255 B.n254 71.676
R1319 B.n250 B.n249 71.676
R1320 B.n245 B.n151 71.676
R1321 B.n243 B.n242 71.676
R1322 B.n238 B.n237 71.676
R1323 B.n235 B.n234 71.676
R1324 B.n230 B.n229 71.676
R1325 B.n227 B.n226 71.676
R1326 B.n222 B.n221 71.676
R1327 B.n219 B.n218 71.676
R1328 B.n214 B.n213 71.676
R1329 B.n211 B.n210 71.676
R1330 B.n206 B.n205 71.676
R1331 B.n203 B.n202 71.676
R1332 B.n198 B.n197 71.676
R1333 B.n195 B.n194 71.676
R1334 B.n190 B.n189 71.676
R1335 B.n187 B.n186 71.676
R1336 B.n182 B.n181 71.676
R1337 B.n179 B.n178 71.676
R1338 B.n174 B.n173 71.676
R1339 B.n171 B.n119 71.676
R1340 B.n646 B.n645 71.676
R1341 B.n646 B.n2 71.676
R1342 B.n526 B.n59 59.5399
R1343 B.n508 B.n65 59.5399
R1344 B.n150 B.n149 59.5399
R1345 B.n268 B.n143 59.5399
R1346 B.n349 B.n116 44.8581
R1347 B.n355 B.n116 44.8581
R1348 B.n355 B.n111 44.8581
R1349 B.n361 B.n111 44.8581
R1350 B.n361 B.n112 44.8581
R1351 B.n367 B.n104 44.8581
R1352 B.n373 B.n104 44.8581
R1353 B.n373 B.n100 44.8581
R1354 B.n379 B.n100 44.8581
R1355 B.n379 B.n96 44.8581
R1356 B.n385 B.n96 44.8581
R1357 B.n385 B.n92 44.8581
R1358 B.n392 B.n92 44.8581
R1359 B.n398 B.n88 44.8581
R1360 B.n398 B.n4 44.8581
R1361 B.n644 B.n4 44.8581
R1362 B.n644 B.n643 44.8581
R1363 B.n643 B.n642 44.8581
R1364 B.n642 B.n8 44.8581
R1365 B.n407 B.n8 44.8581
R1366 B.n635 B.n634 44.8581
R1367 B.n634 B.n633 44.8581
R1368 B.n633 B.n15 44.8581
R1369 B.n627 B.n15 44.8581
R1370 B.n627 B.n626 44.8581
R1371 B.n626 B.n625 44.8581
R1372 B.n625 B.n22 44.8581
R1373 B.n619 B.n22 44.8581
R1374 B.n618 B.n617 44.8581
R1375 B.n617 B.n29 44.8581
R1376 B.n611 B.n29 44.8581
R1377 B.n611 B.n610 44.8581
R1378 B.n610 B.n609 44.8581
R1379 B.n112 B.t3 41.5597
R1380 B.t7 B.n618 41.5597
R1381 B.n59 B.n58 34.1338
R1382 B.n65 B.n64 34.1338
R1383 B.n149 B.n148 34.1338
R1384 B.n143 B.n142 34.1338
R1385 B.n347 B.n346 33.5615
R1386 B.n351 B.n118 33.5615
R1387 B.n428 B.n427 33.5615
R1388 B.n607 B.n606 33.5615
R1389 B.t1 B.n88 31.005
R1390 B.n407 B.t0 31.005
R1391 B B.n647 18.0485
R1392 B.n392 B.t1 13.8536
R1393 B.n635 B.t0 13.8536
R1394 B.n347 B.n114 10.6151
R1395 B.n357 B.n114 10.6151
R1396 B.n358 B.n357 10.6151
R1397 B.n359 B.n358 10.6151
R1398 B.n359 B.n106 10.6151
R1399 B.n369 B.n106 10.6151
R1400 B.n370 B.n369 10.6151
R1401 B.n371 B.n370 10.6151
R1402 B.n371 B.n98 10.6151
R1403 B.n381 B.n98 10.6151
R1404 B.n382 B.n381 10.6151
R1405 B.n383 B.n382 10.6151
R1406 B.n383 B.n90 10.6151
R1407 B.n394 B.n90 10.6151
R1408 B.n395 B.n394 10.6151
R1409 B.n396 B.n395 10.6151
R1410 B.n396 B.n0 10.6151
R1411 B.n346 B.n345 10.6151
R1412 B.n345 B.n122 10.6151
R1413 B.n340 B.n122 10.6151
R1414 B.n340 B.n339 10.6151
R1415 B.n339 B.n124 10.6151
R1416 B.n334 B.n124 10.6151
R1417 B.n334 B.n333 10.6151
R1418 B.n333 B.n332 10.6151
R1419 B.n332 B.n126 10.6151
R1420 B.n326 B.n126 10.6151
R1421 B.n326 B.n325 10.6151
R1422 B.n325 B.n324 10.6151
R1423 B.n324 B.n128 10.6151
R1424 B.n318 B.n128 10.6151
R1425 B.n318 B.n317 10.6151
R1426 B.n317 B.n316 10.6151
R1427 B.n316 B.n130 10.6151
R1428 B.n310 B.n130 10.6151
R1429 B.n310 B.n309 10.6151
R1430 B.n309 B.n308 10.6151
R1431 B.n308 B.n132 10.6151
R1432 B.n302 B.n132 10.6151
R1433 B.n302 B.n301 10.6151
R1434 B.n301 B.n300 10.6151
R1435 B.n300 B.n134 10.6151
R1436 B.n294 B.n134 10.6151
R1437 B.n294 B.n293 10.6151
R1438 B.n293 B.n292 10.6151
R1439 B.n292 B.n136 10.6151
R1440 B.n286 B.n136 10.6151
R1441 B.n286 B.n285 10.6151
R1442 B.n285 B.n284 10.6151
R1443 B.n284 B.n138 10.6151
R1444 B.n278 B.n138 10.6151
R1445 B.n278 B.n277 10.6151
R1446 B.n277 B.n276 10.6151
R1447 B.n276 B.n140 10.6151
R1448 B.n270 B.n140 10.6151
R1449 B.n270 B.n269 10.6151
R1450 B.n267 B.n144 10.6151
R1451 B.n261 B.n144 10.6151
R1452 B.n261 B.n260 10.6151
R1453 B.n260 B.n259 10.6151
R1454 B.n259 B.n146 10.6151
R1455 B.n253 B.n146 10.6151
R1456 B.n253 B.n252 10.6151
R1457 B.n252 B.n251 10.6151
R1458 B.n247 B.n246 10.6151
R1459 B.n246 B.n152 10.6151
R1460 B.n241 B.n152 10.6151
R1461 B.n241 B.n240 10.6151
R1462 B.n240 B.n239 10.6151
R1463 B.n239 B.n154 10.6151
R1464 B.n233 B.n154 10.6151
R1465 B.n233 B.n232 10.6151
R1466 B.n232 B.n231 10.6151
R1467 B.n231 B.n156 10.6151
R1468 B.n225 B.n156 10.6151
R1469 B.n225 B.n224 10.6151
R1470 B.n224 B.n223 10.6151
R1471 B.n223 B.n158 10.6151
R1472 B.n217 B.n158 10.6151
R1473 B.n217 B.n216 10.6151
R1474 B.n216 B.n215 10.6151
R1475 B.n215 B.n160 10.6151
R1476 B.n209 B.n160 10.6151
R1477 B.n209 B.n208 10.6151
R1478 B.n208 B.n207 10.6151
R1479 B.n207 B.n162 10.6151
R1480 B.n201 B.n162 10.6151
R1481 B.n201 B.n200 10.6151
R1482 B.n200 B.n199 10.6151
R1483 B.n199 B.n164 10.6151
R1484 B.n193 B.n164 10.6151
R1485 B.n193 B.n192 10.6151
R1486 B.n192 B.n191 10.6151
R1487 B.n191 B.n166 10.6151
R1488 B.n185 B.n166 10.6151
R1489 B.n185 B.n184 10.6151
R1490 B.n184 B.n183 10.6151
R1491 B.n183 B.n168 10.6151
R1492 B.n177 B.n168 10.6151
R1493 B.n177 B.n176 10.6151
R1494 B.n176 B.n175 10.6151
R1495 B.n175 B.n170 10.6151
R1496 B.n170 B.n118 10.6151
R1497 B.n352 B.n351 10.6151
R1498 B.n353 B.n352 10.6151
R1499 B.n353 B.n109 10.6151
R1500 B.n363 B.n109 10.6151
R1501 B.n364 B.n363 10.6151
R1502 B.n365 B.n364 10.6151
R1503 B.n365 B.n102 10.6151
R1504 B.n375 B.n102 10.6151
R1505 B.n376 B.n375 10.6151
R1506 B.n377 B.n376 10.6151
R1507 B.n377 B.n94 10.6151
R1508 B.n387 B.n94 10.6151
R1509 B.n388 B.n387 10.6151
R1510 B.n390 B.n388 10.6151
R1511 B.n390 B.n389 10.6151
R1512 B.n389 B.n86 10.6151
R1513 B.n401 B.n86 10.6151
R1514 B.n402 B.n401 10.6151
R1515 B.n403 B.n402 10.6151
R1516 B.n404 B.n403 10.6151
R1517 B.n405 B.n404 10.6151
R1518 B.n409 B.n405 10.6151
R1519 B.n410 B.n409 10.6151
R1520 B.n411 B.n410 10.6151
R1521 B.n412 B.n411 10.6151
R1522 B.n414 B.n412 10.6151
R1523 B.n415 B.n414 10.6151
R1524 B.n416 B.n415 10.6151
R1525 B.n417 B.n416 10.6151
R1526 B.n419 B.n417 10.6151
R1527 B.n420 B.n419 10.6151
R1528 B.n421 B.n420 10.6151
R1529 B.n422 B.n421 10.6151
R1530 B.n424 B.n422 10.6151
R1531 B.n425 B.n424 10.6151
R1532 B.n426 B.n425 10.6151
R1533 B.n427 B.n426 10.6151
R1534 B.n639 B.n1 10.6151
R1535 B.n639 B.n638 10.6151
R1536 B.n638 B.n637 10.6151
R1537 B.n637 B.n10 10.6151
R1538 B.n631 B.n10 10.6151
R1539 B.n631 B.n630 10.6151
R1540 B.n630 B.n629 10.6151
R1541 B.n629 B.n17 10.6151
R1542 B.n623 B.n17 10.6151
R1543 B.n623 B.n622 10.6151
R1544 B.n622 B.n621 10.6151
R1545 B.n621 B.n24 10.6151
R1546 B.n615 B.n24 10.6151
R1547 B.n615 B.n614 10.6151
R1548 B.n614 B.n613 10.6151
R1549 B.n613 B.n31 10.6151
R1550 B.n607 B.n31 10.6151
R1551 B.n606 B.n605 10.6151
R1552 B.n605 B.n38 10.6151
R1553 B.n599 B.n38 10.6151
R1554 B.n599 B.n598 10.6151
R1555 B.n598 B.n597 10.6151
R1556 B.n597 B.n40 10.6151
R1557 B.n591 B.n40 10.6151
R1558 B.n591 B.n590 10.6151
R1559 B.n590 B.n589 10.6151
R1560 B.n589 B.n42 10.6151
R1561 B.n583 B.n42 10.6151
R1562 B.n583 B.n582 10.6151
R1563 B.n582 B.n581 10.6151
R1564 B.n581 B.n44 10.6151
R1565 B.n575 B.n44 10.6151
R1566 B.n575 B.n574 10.6151
R1567 B.n574 B.n573 10.6151
R1568 B.n573 B.n46 10.6151
R1569 B.n567 B.n46 10.6151
R1570 B.n567 B.n566 10.6151
R1571 B.n566 B.n565 10.6151
R1572 B.n565 B.n48 10.6151
R1573 B.n559 B.n48 10.6151
R1574 B.n559 B.n558 10.6151
R1575 B.n558 B.n557 10.6151
R1576 B.n557 B.n50 10.6151
R1577 B.n551 B.n50 10.6151
R1578 B.n551 B.n550 10.6151
R1579 B.n550 B.n549 10.6151
R1580 B.n549 B.n52 10.6151
R1581 B.n543 B.n52 10.6151
R1582 B.n543 B.n542 10.6151
R1583 B.n542 B.n541 10.6151
R1584 B.n541 B.n54 10.6151
R1585 B.n535 B.n54 10.6151
R1586 B.n535 B.n534 10.6151
R1587 B.n534 B.n533 10.6151
R1588 B.n533 B.n56 10.6151
R1589 B.n527 B.n56 10.6151
R1590 B.n525 B.n524 10.6151
R1591 B.n524 B.n60 10.6151
R1592 B.n518 B.n60 10.6151
R1593 B.n518 B.n517 10.6151
R1594 B.n517 B.n516 10.6151
R1595 B.n516 B.n62 10.6151
R1596 B.n510 B.n62 10.6151
R1597 B.n510 B.n509 10.6151
R1598 B.n507 B.n66 10.6151
R1599 B.n501 B.n66 10.6151
R1600 B.n501 B.n500 10.6151
R1601 B.n500 B.n499 10.6151
R1602 B.n499 B.n68 10.6151
R1603 B.n493 B.n68 10.6151
R1604 B.n493 B.n492 10.6151
R1605 B.n492 B.n491 10.6151
R1606 B.n491 B.n70 10.6151
R1607 B.n485 B.n70 10.6151
R1608 B.n485 B.n484 10.6151
R1609 B.n484 B.n483 10.6151
R1610 B.n483 B.n72 10.6151
R1611 B.n477 B.n72 10.6151
R1612 B.n477 B.n476 10.6151
R1613 B.n476 B.n475 10.6151
R1614 B.n475 B.n74 10.6151
R1615 B.n469 B.n74 10.6151
R1616 B.n469 B.n468 10.6151
R1617 B.n468 B.n467 10.6151
R1618 B.n467 B.n76 10.6151
R1619 B.n461 B.n76 10.6151
R1620 B.n461 B.n460 10.6151
R1621 B.n460 B.n459 10.6151
R1622 B.n459 B.n78 10.6151
R1623 B.n453 B.n78 10.6151
R1624 B.n453 B.n452 10.6151
R1625 B.n452 B.n451 10.6151
R1626 B.n451 B.n80 10.6151
R1627 B.n445 B.n80 10.6151
R1628 B.n445 B.n444 10.6151
R1629 B.n444 B.n443 10.6151
R1630 B.n443 B.n82 10.6151
R1631 B.n437 B.n82 10.6151
R1632 B.n437 B.n436 10.6151
R1633 B.n436 B.n435 10.6151
R1634 B.n435 B.n84 10.6151
R1635 B.n429 B.n84 10.6151
R1636 B.n429 B.n428 10.6151
R1637 B.n647 B.n0 8.11757
R1638 B.n647 B.n1 8.11757
R1639 B.n268 B.n267 6.5566
R1640 B.n251 B.n150 6.5566
R1641 B.n526 B.n525 6.5566
R1642 B.n509 B.n508 6.5566
R1643 B.n269 B.n268 4.05904
R1644 B.n247 B.n150 4.05904
R1645 B.n527 B.n526 4.05904
R1646 B.n508 B.n507 4.05904
R1647 B.n367 B.t3 3.29885
R1648 B.n619 B.t7 3.29885
R1649 VN VN.t1 341.923
R1650 VN VN.t0 300.683
R1651 VDD2.n117 VDD2.n61 289.615
R1652 VDD2.n56 VDD2.n0 289.615
R1653 VDD2.n118 VDD2.n117 185
R1654 VDD2.n116 VDD2.n115 185
R1655 VDD2.n65 VDD2.n64 185
R1656 VDD2.n110 VDD2.n109 185
R1657 VDD2.n108 VDD2.n107 185
R1658 VDD2.n69 VDD2.n68 185
R1659 VDD2.n73 VDD2.n71 185
R1660 VDD2.n102 VDD2.n101 185
R1661 VDD2.n100 VDD2.n99 185
R1662 VDD2.n75 VDD2.n74 185
R1663 VDD2.n94 VDD2.n93 185
R1664 VDD2.n92 VDD2.n91 185
R1665 VDD2.n79 VDD2.n78 185
R1666 VDD2.n86 VDD2.n85 185
R1667 VDD2.n84 VDD2.n83 185
R1668 VDD2.n21 VDD2.n20 185
R1669 VDD2.n23 VDD2.n22 185
R1670 VDD2.n16 VDD2.n15 185
R1671 VDD2.n29 VDD2.n28 185
R1672 VDD2.n31 VDD2.n30 185
R1673 VDD2.n12 VDD2.n11 185
R1674 VDD2.n38 VDD2.n37 185
R1675 VDD2.n39 VDD2.n10 185
R1676 VDD2.n41 VDD2.n40 185
R1677 VDD2.n8 VDD2.n7 185
R1678 VDD2.n47 VDD2.n46 185
R1679 VDD2.n49 VDD2.n48 185
R1680 VDD2.n4 VDD2.n3 185
R1681 VDD2.n55 VDD2.n54 185
R1682 VDD2.n57 VDD2.n56 185
R1683 VDD2.n82 VDD2.t0 149.524
R1684 VDD2.n19 VDD2.t1 149.524
R1685 VDD2.n117 VDD2.n116 104.615
R1686 VDD2.n116 VDD2.n64 104.615
R1687 VDD2.n109 VDD2.n64 104.615
R1688 VDD2.n109 VDD2.n108 104.615
R1689 VDD2.n108 VDD2.n68 104.615
R1690 VDD2.n73 VDD2.n68 104.615
R1691 VDD2.n101 VDD2.n73 104.615
R1692 VDD2.n101 VDD2.n100 104.615
R1693 VDD2.n100 VDD2.n74 104.615
R1694 VDD2.n93 VDD2.n74 104.615
R1695 VDD2.n93 VDD2.n92 104.615
R1696 VDD2.n92 VDD2.n78 104.615
R1697 VDD2.n85 VDD2.n78 104.615
R1698 VDD2.n85 VDD2.n84 104.615
R1699 VDD2.n22 VDD2.n21 104.615
R1700 VDD2.n22 VDD2.n15 104.615
R1701 VDD2.n29 VDD2.n15 104.615
R1702 VDD2.n30 VDD2.n29 104.615
R1703 VDD2.n30 VDD2.n11 104.615
R1704 VDD2.n38 VDD2.n11 104.615
R1705 VDD2.n39 VDD2.n38 104.615
R1706 VDD2.n40 VDD2.n39 104.615
R1707 VDD2.n40 VDD2.n7 104.615
R1708 VDD2.n47 VDD2.n7 104.615
R1709 VDD2.n48 VDD2.n47 104.615
R1710 VDD2.n48 VDD2.n3 104.615
R1711 VDD2.n55 VDD2.n3 104.615
R1712 VDD2.n56 VDD2.n55 104.615
R1713 VDD2.n122 VDD2.n60 85.3856
R1714 VDD2.n84 VDD2.t0 52.3082
R1715 VDD2.n21 VDD2.t1 52.3082
R1716 VDD2.n122 VDD2.n121 48.8641
R1717 VDD2.n71 VDD2.n69 13.1884
R1718 VDD2.n41 VDD2.n8 13.1884
R1719 VDD2.n107 VDD2.n106 12.8005
R1720 VDD2.n103 VDD2.n102 12.8005
R1721 VDD2.n42 VDD2.n10 12.8005
R1722 VDD2.n46 VDD2.n45 12.8005
R1723 VDD2.n110 VDD2.n67 12.0247
R1724 VDD2.n99 VDD2.n72 12.0247
R1725 VDD2.n37 VDD2.n36 12.0247
R1726 VDD2.n49 VDD2.n6 12.0247
R1727 VDD2.n111 VDD2.n65 11.249
R1728 VDD2.n98 VDD2.n75 11.249
R1729 VDD2.n35 VDD2.n12 11.249
R1730 VDD2.n50 VDD2.n4 11.249
R1731 VDD2.n115 VDD2.n114 10.4732
R1732 VDD2.n95 VDD2.n94 10.4732
R1733 VDD2.n32 VDD2.n31 10.4732
R1734 VDD2.n54 VDD2.n53 10.4732
R1735 VDD2.n83 VDD2.n82 10.2747
R1736 VDD2.n20 VDD2.n19 10.2747
R1737 VDD2.n118 VDD2.n63 9.69747
R1738 VDD2.n91 VDD2.n77 9.69747
R1739 VDD2.n28 VDD2.n14 9.69747
R1740 VDD2.n57 VDD2.n2 9.69747
R1741 VDD2.n121 VDD2.n120 9.45567
R1742 VDD2.n60 VDD2.n59 9.45567
R1743 VDD2.n81 VDD2.n80 9.3005
R1744 VDD2.n88 VDD2.n87 9.3005
R1745 VDD2.n90 VDD2.n89 9.3005
R1746 VDD2.n77 VDD2.n76 9.3005
R1747 VDD2.n96 VDD2.n95 9.3005
R1748 VDD2.n98 VDD2.n97 9.3005
R1749 VDD2.n72 VDD2.n70 9.3005
R1750 VDD2.n104 VDD2.n103 9.3005
R1751 VDD2.n120 VDD2.n119 9.3005
R1752 VDD2.n63 VDD2.n62 9.3005
R1753 VDD2.n114 VDD2.n113 9.3005
R1754 VDD2.n112 VDD2.n111 9.3005
R1755 VDD2.n67 VDD2.n66 9.3005
R1756 VDD2.n106 VDD2.n105 9.3005
R1757 VDD2.n59 VDD2.n58 9.3005
R1758 VDD2.n2 VDD2.n1 9.3005
R1759 VDD2.n53 VDD2.n52 9.3005
R1760 VDD2.n51 VDD2.n50 9.3005
R1761 VDD2.n6 VDD2.n5 9.3005
R1762 VDD2.n45 VDD2.n44 9.3005
R1763 VDD2.n18 VDD2.n17 9.3005
R1764 VDD2.n25 VDD2.n24 9.3005
R1765 VDD2.n27 VDD2.n26 9.3005
R1766 VDD2.n14 VDD2.n13 9.3005
R1767 VDD2.n33 VDD2.n32 9.3005
R1768 VDD2.n35 VDD2.n34 9.3005
R1769 VDD2.n36 VDD2.n9 9.3005
R1770 VDD2.n43 VDD2.n42 9.3005
R1771 VDD2.n119 VDD2.n61 8.92171
R1772 VDD2.n90 VDD2.n79 8.92171
R1773 VDD2.n27 VDD2.n16 8.92171
R1774 VDD2.n58 VDD2.n0 8.92171
R1775 VDD2.n87 VDD2.n86 8.14595
R1776 VDD2.n24 VDD2.n23 8.14595
R1777 VDD2.n83 VDD2.n81 7.3702
R1778 VDD2.n20 VDD2.n18 7.3702
R1779 VDD2.n86 VDD2.n81 5.81868
R1780 VDD2.n23 VDD2.n18 5.81868
R1781 VDD2.n121 VDD2.n61 5.04292
R1782 VDD2.n87 VDD2.n79 5.04292
R1783 VDD2.n24 VDD2.n16 5.04292
R1784 VDD2.n60 VDD2.n0 5.04292
R1785 VDD2.n119 VDD2.n118 4.26717
R1786 VDD2.n91 VDD2.n90 4.26717
R1787 VDD2.n28 VDD2.n27 4.26717
R1788 VDD2.n58 VDD2.n57 4.26717
R1789 VDD2.n115 VDD2.n63 3.49141
R1790 VDD2.n94 VDD2.n77 3.49141
R1791 VDD2.n31 VDD2.n14 3.49141
R1792 VDD2.n54 VDD2.n2 3.49141
R1793 VDD2.n82 VDD2.n80 2.84303
R1794 VDD2.n19 VDD2.n17 2.84303
R1795 VDD2.n114 VDD2.n65 2.71565
R1796 VDD2.n95 VDD2.n75 2.71565
R1797 VDD2.n32 VDD2.n12 2.71565
R1798 VDD2.n53 VDD2.n4 2.71565
R1799 VDD2.n111 VDD2.n110 1.93989
R1800 VDD2.n99 VDD2.n98 1.93989
R1801 VDD2.n37 VDD2.n35 1.93989
R1802 VDD2.n50 VDD2.n49 1.93989
R1803 VDD2.n107 VDD2.n67 1.16414
R1804 VDD2.n102 VDD2.n72 1.16414
R1805 VDD2.n36 VDD2.n10 1.16414
R1806 VDD2.n46 VDD2.n6 1.16414
R1807 VDD2 VDD2.n122 0.438
R1808 VDD2.n106 VDD2.n69 0.388379
R1809 VDD2.n103 VDD2.n71 0.388379
R1810 VDD2.n42 VDD2.n41 0.388379
R1811 VDD2.n45 VDD2.n8 0.388379
R1812 VDD2.n120 VDD2.n62 0.155672
R1813 VDD2.n113 VDD2.n62 0.155672
R1814 VDD2.n113 VDD2.n112 0.155672
R1815 VDD2.n112 VDD2.n66 0.155672
R1816 VDD2.n105 VDD2.n66 0.155672
R1817 VDD2.n105 VDD2.n104 0.155672
R1818 VDD2.n104 VDD2.n70 0.155672
R1819 VDD2.n97 VDD2.n70 0.155672
R1820 VDD2.n97 VDD2.n96 0.155672
R1821 VDD2.n96 VDD2.n76 0.155672
R1822 VDD2.n89 VDD2.n76 0.155672
R1823 VDD2.n89 VDD2.n88 0.155672
R1824 VDD2.n88 VDD2.n80 0.155672
R1825 VDD2.n25 VDD2.n17 0.155672
R1826 VDD2.n26 VDD2.n25 0.155672
R1827 VDD2.n26 VDD2.n13 0.155672
R1828 VDD2.n33 VDD2.n13 0.155672
R1829 VDD2.n34 VDD2.n33 0.155672
R1830 VDD2.n34 VDD2.n9 0.155672
R1831 VDD2.n43 VDD2.n9 0.155672
R1832 VDD2.n44 VDD2.n43 0.155672
R1833 VDD2.n44 VDD2.n5 0.155672
R1834 VDD2.n51 VDD2.n5 0.155672
R1835 VDD2.n52 VDD2.n51 0.155672
R1836 VDD2.n52 VDD2.n1 0.155672
R1837 VDD2.n59 VDD2.n1 0.155672
C0 VTAIL VDD2 4.94444f
C1 VDD1 VDD2 0.538277f
C2 VN VP 4.79659f
C3 VTAIL VN 1.97262f
C4 VTAIL VP 1.98703f
C5 VDD1 VN 0.147252f
C6 VDD1 VP 2.49115f
C7 VN VDD2 2.35797f
C8 VDD2 VP 0.283663f
C9 VDD1 VTAIL 4.90328f
C10 VDD2 B 3.910869f
C11 VDD1 B 6.35344f
C12 VTAIL B 6.494531f
C13 VN B 8.46161f
C14 VP B 4.883409f
C15 VDD2.n0 B 0.027934f
C16 VDD2.n1 B 0.020263f
C17 VDD2.n2 B 0.010888f
C18 VDD2.n3 B 0.025736f
C19 VDD2.n4 B 0.011529f
C20 VDD2.n5 B 0.020263f
C21 VDD2.n6 B 0.010888f
C22 VDD2.n7 B 0.025736f
C23 VDD2.n8 B 0.011209f
C24 VDD2.n9 B 0.020263f
C25 VDD2.n10 B 0.011529f
C26 VDD2.n11 B 0.025736f
C27 VDD2.n12 B 0.011529f
C28 VDD2.n13 B 0.020263f
C29 VDD2.n14 B 0.010888f
C30 VDD2.n15 B 0.025736f
C31 VDD2.n16 B 0.011529f
C32 VDD2.n17 B 0.968149f
C33 VDD2.n18 B 0.010888f
C34 VDD2.t1 B 0.043401f
C35 VDD2.n19 B 0.141426f
C36 VDD2.n20 B 0.018194f
C37 VDD2.n21 B 0.019302f
C38 VDD2.n22 B 0.025736f
C39 VDD2.n23 B 0.011529f
C40 VDD2.n24 B 0.010888f
C41 VDD2.n25 B 0.020263f
C42 VDD2.n26 B 0.020263f
C43 VDD2.n27 B 0.010888f
C44 VDD2.n28 B 0.011529f
C45 VDD2.n29 B 0.025736f
C46 VDD2.n30 B 0.025736f
C47 VDD2.n31 B 0.011529f
C48 VDD2.n32 B 0.010888f
C49 VDD2.n33 B 0.020263f
C50 VDD2.n34 B 0.020263f
C51 VDD2.n35 B 0.010888f
C52 VDD2.n36 B 0.010888f
C53 VDD2.n37 B 0.011529f
C54 VDD2.n38 B 0.025736f
C55 VDD2.n39 B 0.025736f
C56 VDD2.n40 B 0.025736f
C57 VDD2.n41 B 0.011209f
C58 VDD2.n42 B 0.010888f
C59 VDD2.n43 B 0.020263f
C60 VDD2.n44 B 0.020263f
C61 VDD2.n45 B 0.010888f
C62 VDD2.n46 B 0.011529f
C63 VDD2.n47 B 0.025736f
C64 VDD2.n48 B 0.025736f
C65 VDD2.n49 B 0.011529f
C66 VDD2.n50 B 0.010888f
C67 VDD2.n51 B 0.020263f
C68 VDD2.n52 B 0.020263f
C69 VDD2.n53 B 0.010888f
C70 VDD2.n54 B 0.011529f
C71 VDD2.n55 B 0.025736f
C72 VDD2.n56 B 0.054747f
C73 VDD2.n57 B 0.011529f
C74 VDD2.n58 B 0.010888f
C75 VDD2.n59 B 0.046837f
C76 VDD2.n60 B 0.517395f
C77 VDD2.n61 B 0.027934f
C78 VDD2.n62 B 0.020263f
C79 VDD2.n63 B 0.010888f
C80 VDD2.n64 B 0.025736f
C81 VDD2.n65 B 0.011529f
C82 VDD2.n66 B 0.020263f
C83 VDD2.n67 B 0.010888f
C84 VDD2.n68 B 0.025736f
C85 VDD2.n69 B 0.011209f
C86 VDD2.n70 B 0.020263f
C87 VDD2.n71 B 0.011209f
C88 VDD2.n72 B 0.010888f
C89 VDD2.n73 B 0.025736f
C90 VDD2.n74 B 0.025736f
C91 VDD2.n75 B 0.011529f
C92 VDD2.n76 B 0.020263f
C93 VDD2.n77 B 0.010888f
C94 VDD2.n78 B 0.025736f
C95 VDD2.n79 B 0.011529f
C96 VDD2.n80 B 0.968149f
C97 VDD2.n81 B 0.010888f
C98 VDD2.t0 B 0.043401f
C99 VDD2.n82 B 0.141426f
C100 VDD2.n83 B 0.018194f
C101 VDD2.n84 B 0.019302f
C102 VDD2.n85 B 0.025736f
C103 VDD2.n86 B 0.011529f
C104 VDD2.n87 B 0.010888f
C105 VDD2.n88 B 0.020263f
C106 VDD2.n89 B 0.020263f
C107 VDD2.n90 B 0.010888f
C108 VDD2.n91 B 0.011529f
C109 VDD2.n92 B 0.025736f
C110 VDD2.n93 B 0.025736f
C111 VDD2.n94 B 0.011529f
C112 VDD2.n95 B 0.010888f
C113 VDD2.n96 B 0.020263f
C114 VDD2.n97 B 0.020263f
C115 VDD2.n98 B 0.010888f
C116 VDD2.n99 B 0.011529f
C117 VDD2.n100 B 0.025736f
C118 VDD2.n101 B 0.025736f
C119 VDD2.n102 B 0.011529f
C120 VDD2.n103 B 0.010888f
C121 VDD2.n104 B 0.020263f
C122 VDD2.n105 B 0.020263f
C123 VDD2.n106 B 0.010888f
C124 VDD2.n107 B 0.011529f
C125 VDD2.n108 B 0.025736f
C126 VDD2.n109 B 0.025736f
C127 VDD2.n110 B 0.011529f
C128 VDD2.n111 B 0.010888f
C129 VDD2.n112 B 0.020263f
C130 VDD2.n113 B 0.020263f
C131 VDD2.n114 B 0.010888f
C132 VDD2.n115 B 0.011529f
C133 VDD2.n116 B 0.025736f
C134 VDD2.n117 B 0.054747f
C135 VDD2.n118 B 0.011529f
C136 VDD2.n119 B 0.010888f
C137 VDD2.n120 B 0.046837f
C138 VDD2.n121 B 0.044525f
C139 VDD2.n122 B 2.23759f
C140 VN.t0 B 1.73526f
C141 VN.t1 B 1.9584f
C142 VDD1.n0 B 0.02803f
C143 VDD1.n1 B 0.020332f
C144 VDD1.n2 B 0.010925f
C145 VDD1.n3 B 0.025824f
C146 VDD1.n4 B 0.011568f
C147 VDD1.n5 B 0.020332f
C148 VDD1.n6 B 0.010925f
C149 VDD1.n7 B 0.025824f
C150 VDD1.n8 B 0.011247f
C151 VDD1.n9 B 0.020332f
C152 VDD1.n10 B 0.011247f
C153 VDD1.n11 B 0.010925f
C154 VDD1.n12 B 0.025824f
C155 VDD1.n13 B 0.025824f
C156 VDD1.n14 B 0.011568f
C157 VDD1.n15 B 0.020332f
C158 VDD1.n16 B 0.010925f
C159 VDD1.n17 B 0.025824f
C160 VDD1.n18 B 0.011568f
C161 VDD1.n19 B 0.971452f
C162 VDD1.n20 B 0.010925f
C163 VDD1.t1 B 0.04355f
C164 VDD1.n21 B 0.141908f
C165 VDD1.n22 B 0.018256f
C166 VDD1.n23 B 0.019368f
C167 VDD1.n24 B 0.025824f
C168 VDD1.n25 B 0.011568f
C169 VDD1.n26 B 0.010925f
C170 VDD1.n27 B 0.020332f
C171 VDD1.n28 B 0.020332f
C172 VDD1.n29 B 0.010925f
C173 VDD1.n30 B 0.011568f
C174 VDD1.n31 B 0.025824f
C175 VDD1.n32 B 0.025824f
C176 VDD1.n33 B 0.011568f
C177 VDD1.n34 B 0.010925f
C178 VDD1.n35 B 0.020332f
C179 VDD1.n36 B 0.020332f
C180 VDD1.n37 B 0.010925f
C181 VDD1.n38 B 0.011568f
C182 VDD1.n39 B 0.025824f
C183 VDD1.n40 B 0.025824f
C184 VDD1.n41 B 0.011568f
C185 VDD1.n42 B 0.010925f
C186 VDD1.n43 B 0.020332f
C187 VDD1.n44 B 0.020332f
C188 VDD1.n45 B 0.010925f
C189 VDD1.n46 B 0.011568f
C190 VDD1.n47 B 0.025824f
C191 VDD1.n48 B 0.025824f
C192 VDD1.n49 B 0.011568f
C193 VDD1.n50 B 0.010925f
C194 VDD1.n51 B 0.020332f
C195 VDD1.n52 B 0.020332f
C196 VDD1.n53 B 0.010925f
C197 VDD1.n54 B 0.011568f
C198 VDD1.n55 B 0.025824f
C199 VDD1.n56 B 0.054934f
C200 VDD1.n57 B 0.011568f
C201 VDD1.n58 B 0.010925f
C202 VDD1.n59 B 0.046996f
C203 VDD1.n60 B 0.045279f
C204 VDD1.n61 B 0.02803f
C205 VDD1.n62 B 0.020332f
C206 VDD1.n63 B 0.010925f
C207 VDD1.n64 B 0.025824f
C208 VDD1.n65 B 0.011568f
C209 VDD1.n66 B 0.020332f
C210 VDD1.n67 B 0.010925f
C211 VDD1.n68 B 0.025824f
C212 VDD1.n69 B 0.011247f
C213 VDD1.n70 B 0.020332f
C214 VDD1.n71 B 0.011568f
C215 VDD1.n72 B 0.025824f
C216 VDD1.n73 B 0.011568f
C217 VDD1.n74 B 0.020332f
C218 VDD1.n75 B 0.010925f
C219 VDD1.n76 B 0.025824f
C220 VDD1.n77 B 0.011568f
C221 VDD1.n78 B 0.971452f
C222 VDD1.n79 B 0.010925f
C223 VDD1.t0 B 0.04355f
C224 VDD1.n80 B 0.141908f
C225 VDD1.n81 B 0.018256f
C226 VDD1.n82 B 0.019368f
C227 VDD1.n83 B 0.025824f
C228 VDD1.n84 B 0.011568f
C229 VDD1.n85 B 0.010925f
C230 VDD1.n86 B 0.020332f
C231 VDD1.n87 B 0.020332f
C232 VDD1.n88 B 0.010925f
C233 VDD1.n89 B 0.011568f
C234 VDD1.n90 B 0.025824f
C235 VDD1.n91 B 0.025824f
C236 VDD1.n92 B 0.011568f
C237 VDD1.n93 B 0.010925f
C238 VDD1.n94 B 0.020332f
C239 VDD1.n95 B 0.020332f
C240 VDD1.n96 B 0.010925f
C241 VDD1.n97 B 0.010925f
C242 VDD1.n98 B 0.011568f
C243 VDD1.n99 B 0.025824f
C244 VDD1.n100 B 0.025824f
C245 VDD1.n101 B 0.025824f
C246 VDD1.n102 B 0.011247f
C247 VDD1.n103 B 0.010925f
C248 VDD1.n104 B 0.020332f
C249 VDD1.n105 B 0.020332f
C250 VDD1.n106 B 0.010925f
C251 VDD1.n107 B 0.011568f
C252 VDD1.n108 B 0.025824f
C253 VDD1.n109 B 0.025824f
C254 VDD1.n110 B 0.011568f
C255 VDD1.n111 B 0.010925f
C256 VDD1.n112 B 0.020332f
C257 VDD1.n113 B 0.020332f
C258 VDD1.n114 B 0.010925f
C259 VDD1.n115 B 0.011568f
C260 VDD1.n116 B 0.025824f
C261 VDD1.n117 B 0.054934f
C262 VDD1.n118 B 0.011568f
C263 VDD1.n119 B 0.010925f
C264 VDD1.n120 B 0.046996f
C265 VDD1.n121 B 0.550642f
C266 VTAIL.n0 B 0.020103f
C267 VTAIL.n1 B 0.014582f
C268 VTAIL.n2 B 0.007836f
C269 VTAIL.n3 B 0.018521f
C270 VTAIL.n4 B 0.008297f
C271 VTAIL.n5 B 0.014582f
C272 VTAIL.n6 B 0.007836f
C273 VTAIL.n7 B 0.018521f
C274 VTAIL.n8 B 0.008066f
C275 VTAIL.n9 B 0.014582f
C276 VTAIL.n10 B 0.008297f
C277 VTAIL.n11 B 0.018521f
C278 VTAIL.n12 B 0.008297f
C279 VTAIL.n13 B 0.014582f
C280 VTAIL.n14 B 0.007836f
C281 VTAIL.n15 B 0.018521f
C282 VTAIL.n16 B 0.008297f
C283 VTAIL.n17 B 0.696723f
C284 VTAIL.n18 B 0.007836f
C285 VTAIL.t2 B 0.031234f
C286 VTAIL.n19 B 0.101776f
C287 VTAIL.n20 B 0.013093f
C288 VTAIL.n21 B 0.013891f
C289 VTAIL.n22 B 0.018521f
C290 VTAIL.n23 B 0.008297f
C291 VTAIL.n24 B 0.007836f
C292 VTAIL.n25 B 0.014582f
C293 VTAIL.n26 B 0.014582f
C294 VTAIL.n27 B 0.007836f
C295 VTAIL.n28 B 0.008297f
C296 VTAIL.n29 B 0.018521f
C297 VTAIL.n30 B 0.018521f
C298 VTAIL.n31 B 0.008297f
C299 VTAIL.n32 B 0.007836f
C300 VTAIL.n33 B 0.014582f
C301 VTAIL.n34 B 0.014582f
C302 VTAIL.n35 B 0.007836f
C303 VTAIL.n36 B 0.007836f
C304 VTAIL.n37 B 0.008297f
C305 VTAIL.n38 B 0.018521f
C306 VTAIL.n39 B 0.018521f
C307 VTAIL.n40 B 0.018521f
C308 VTAIL.n41 B 0.008066f
C309 VTAIL.n42 B 0.007836f
C310 VTAIL.n43 B 0.014582f
C311 VTAIL.n44 B 0.014582f
C312 VTAIL.n45 B 0.007836f
C313 VTAIL.n46 B 0.008297f
C314 VTAIL.n47 B 0.018521f
C315 VTAIL.n48 B 0.018521f
C316 VTAIL.n49 B 0.008297f
C317 VTAIL.n50 B 0.007836f
C318 VTAIL.n51 B 0.014582f
C319 VTAIL.n52 B 0.014582f
C320 VTAIL.n53 B 0.007836f
C321 VTAIL.n54 B 0.008297f
C322 VTAIL.n55 B 0.018521f
C323 VTAIL.n56 B 0.039399f
C324 VTAIL.n57 B 0.008297f
C325 VTAIL.n58 B 0.007836f
C326 VTAIL.n59 B 0.033706f
C327 VTAIL.n60 B 0.021974f
C328 VTAIL.n61 B 0.857511f
C329 VTAIL.n62 B 0.020103f
C330 VTAIL.n63 B 0.014582f
C331 VTAIL.n64 B 0.007836f
C332 VTAIL.n65 B 0.018521f
C333 VTAIL.n66 B 0.008297f
C334 VTAIL.n67 B 0.014582f
C335 VTAIL.n68 B 0.007836f
C336 VTAIL.n69 B 0.018521f
C337 VTAIL.n70 B 0.008066f
C338 VTAIL.n71 B 0.014582f
C339 VTAIL.n72 B 0.008066f
C340 VTAIL.n73 B 0.007836f
C341 VTAIL.n74 B 0.018521f
C342 VTAIL.n75 B 0.018521f
C343 VTAIL.n76 B 0.008297f
C344 VTAIL.n77 B 0.014582f
C345 VTAIL.n78 B 0.007836f
C346 VTAIL.n79 B 0.018521f
C347 VTAIL.n80 B 0.008297f
C348 VTAIL.n81 B 0.696723f
C349 VTAIL.n82 B 0.007836f
C350 VTAIL.t1 B 0.031234f
C351 VTAIL.n83 B 0.101776f
C352 VTAIL.n84 B 0.013093f
C353 VTAIL.n85 B 0.013891f
C354 VTAIL.n86 B 0.018521f
C355 VTAIL.n87 B 0.008297f
C356 VTAIL.n88 B 0.007836f
C357 VTAIL.n89 B 0.014582f
C358 VTAIL.n90 B 0.014582f
C359 VTAIL.n91 B 0.007836f
C360 VTAIL.n92 B 0.008297f
C361 VTAIL.n93 B 0.018521f
C362 VTAIL.n94 B 0.018521f
C363 VTAIL.n95 B 0.008297f
C364 VTAIL.n96 B 0.007836f
C365 VTAIL.n97 B 0.014582f
C366 VTAIL.n98 B 0.014582f
C367 VTAIL.n99 B 0.007836f
C368 VTAIL.n100 B 0.008297f
C369 VTAIL.n101 B 0.018521f
C370 VTAIL.n102 B 0.018521f
C371 VTAIL.n103 B 0.008297f
C372 VTAIL.n104 B 0.007836f
C373 VTAIL.n105 B 0.014582f
C374 VTAIL.n106 B 0.014582f
C375 VTAIL.n107 B 0.007836f
C376 VTAIL.n108 B 0.008297f
C377 VTAIL.n109 B 0.018521f
C378 VTAIL.n110 B 0.018521f
C379 VTAIL.n111 B 0.008297f
C380 VTAIL.n112 B 0.007836f
C381 VTAIL.n113 B 0.014582f
C382 VTAIL.n114 B 0.014582f
C383 VTAIL.n115 B 0.007836f
C384 VTAIL.n116 B 0.008297f
C385 VTAIL.n117 B 0.018521f
C386 VTAIL.n118 B 0.039399f
C387 VTAIL.n119 B 0.008297f
C388 VTAIL.n120 B 0.007836f
C389 VTAIL.n121 B 0.033706f
C390 VTAIL.n122 B 0.021974f
C391 VTAIL.n123 B 0.872599f
C392 VTAIL.n124 B 0.020103f
C393 VTAIL.n125 B 0.014582f
C394 VTAIL.n126 B 0.007836f
C395 VTAIL.n127 B 0.018521f
C396 VTAIL.n128 B 0.008297f
C397 VTAIL.n129 B 0.014582f
C398 VTAIL.n130 B 0.007836f
C399 VTAIL.n131 B 0.018521f
C400 VTAIL.n132 B 0.008066f
C401 VTAIL.n133 B 0.014582f
C402 VTAIL.n134 B 0.008066f
C403 VTAIL.n135 B 0.007836f
C404 VTAIL.n136 B 0.018521f
C405 VTAIL.n137 B 0.018521f
C406 VTAIL.n138 B 0.008297f
C407 VTAIL.n139 B 0.014582f
C408 VTAIL.n140 B 0.007836f
C409 VTAIL.n141 B 0.018521f
C410 VTAIL.n142 B 0.008297f
C411 VTAIL.n143 B 0.696723f
C412 VTAIL.n144 B 0.007836f
C413 VTAIL.t3 B 0.031234f
C414 VTAIL.n145 B 0.101776f
C415 VTAIL.n146 B 0.013093f
C416 VTAIL.n147 B 0.013891f
C417 VTAIL.n148 B 0.018521f
C418 VTAIL.n149 B 0.008297f
C419 VTAIL.n150 B 0.007836f
C420 VTAIL.n151 B 0.014582f
C421 VTAIL.n152 B 0.014582f
C422 VTAIL.n153 B 0.007836f
C423 VTAIL.n154 B 0.008297f
C424 VTAIL.n155 B 0.018521f
C425 VTAIL.n156 B 0.018521f
C426 VTAIL.n157 B 0.008297f
C427 VTAIL.n158 B 0.007836f
C428 VTAIL.n159 B 0.014582f
C429 VTAIL.n160 B 0.014582f
C430 VTAIL.n161 B 0.007836f
C431 VTAIL.n162 B 0.008297f
C432 VTAIL.n163 B 0.018521f
C433 VTAIL.n164 B 0.018521f
C434 VTAIL.n165 B 0.008297f
C435 VTAIL.n166 B 0.007836f
C436 VTAIL.n167 B 0.014582f
C437 VTAIL.n168 B 0.014582f
C438 VTAIL.n169 B 0.007836f
C439 VTAIL.n170 B 0.008297f
C440 VTAIL.n171 B 0.018521f
C441 VTAIL.n172 B 0.018521f
C442 VTAIL.n173 B 0.008297f
C443 VTAIL.n174 B 0.007836f
C444 VTAIL.n175 B 0.014582f
C445 VTAIL.n176 B 0.014582f
C446 VTAIL.n177 B 0.007836f
C447 VTAIL.n178 B 0.008297f
C448 VTAIL.n179 B 0.018521f
C449 VTAIL.n180 B 0.039399f
C450 VTAIL.n181 B 0.008297f
C451 VTAIL.n182 B 0.007836f
C452 VTAIL.n183 B 0.033706f
C453 VTAIL.n184 B 0.021974f
C454 VTAIL.n185 B 0.801309f
C455 VTAIL.n186 B 0.020103f
C456 VTAIL.n187 B 0.014582f
C457 VTAIL.n188 B 0.007836f
C458 VTAIL.n189 B 0.018521f
C459 VTAIL.n190 B 0.008297f
C460 VTAIL.n191 B 0.014582f
C461 VTAIL.n192 B 0.007836f
C462 VTAIL.n193 B 0.018521f
C463 VTAIL.n194 B 0.008066f
C464 VTAIL.n195 B 0.014582f
C465 VTAIL.n196 B 0.008297f
C466 VTAIL.n197 B 0.018521f
C467 VTAIL.n198 B 0.008297f
C468 VTAIL.n199 B 0.014582f
C469 VTAIL.n200 B 0.007836f
C470 VTAIL.n201 B 0.018521f
C471 VTAIL.n202 B 0.008297f
C472 VTAIL.n203 B 0.696723f
C473 VTAIL.n204 B 0.007836f
C474 VTAIL.t0 B 0.031234f
C475 VTAIL.n205 B 0.101776f
C476 VTAIL.n206 B 0.013093f
C477 VTAIL.n207 B 0.013891f
C478 VTAIL.n208 B 0.018521f
C479 VTAIL.n209 B 0.008297f
C480 VTAIL.n210 B 0.007836f
C481 VTAIL.n211 B 0.014582f
C482 VTAIL.n212 B 0.014582f
C483 VTAIL.n213 B 0.007836f
C484 VTAIL.n214 B 0.008297f
C485 VTAIL.n215 B 0.018521f
C486 VTAIL.n216 B 0.018521f
C487 VTAIL.n217 B 0.008297f
C488 VTAIL.n218 B 0.007836f
C489 VTAIL.n219 B 0.014582f
C490 VTAIL.n220 B 0.014582f
C491 VTAIL.n221 B 0.007836f
C492 VTAIL.n222 B 0.007836f
C493 VTAIL.n223 B 0.008297f
C494 VTAIL.n224 B 0.018521f
C495 VTAIL.n225 B 0.018521f
C496 VTAIL.n226 B 0.018521f
C497 VTAIL.n227 B 0.008066f
C498 VTAIL.n228 B 0.007836f
C499 VTAIL.n229 B 0.014582f
C500 VTAIL.n230 B 0.014582f
C501 VTAIL.n231 B 0.007836f
C502 VTAIL.n232 B 0.008297f
C503 VTAIL.n233 B 0.018521f
C504 VTAIL.n234 B 0.018521f
C505 VTAIL.n235 B 0.008297f
C506 VTAIL.n236 B 0.007836f
C507 VTAIL.n237 B 0.014582f
C508 VTAIL.n238 B 0.014582f
C509 VTAIL.n239 B 0.007836f
C510 VTAIL.n240 B 0.008297f
C511 VTAIL.n241 B 0.018521f
C512 VTAIL.n242 B 0.039399f
C513 VTAIL.n243 B 0.008297f
C514 VTAIL.n244 B 0.007836f
C515 VTAIL.n245 B 0.033706f
C516 VTAIL.n246 B 0.021974f
C517 VTAIL.n247 B 0.758677f
C518 VP.t0 B 1.99504f
C519 VP.t1 B 1.77076f
C520 VP.n0 B 3.5f
.ends

