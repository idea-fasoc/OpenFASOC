* NGSPICE file created from diff_pair_sample_0499.ext - technology: sky130A

.subckt diff_pair_sample_0499 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=0 ps=0 w=6.24 l=2.27
X1 B.t8 B.t6 B.t7 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=0 ps=0 w=6.24 l=2.27
X2 VDD1.t9 VP.t0 VTAIL.t16 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=1.0296 ps=6.57 w=6.24 l=2.27
X3 B.t5 B.t3 B.t4 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=0 ps=0 w=6.24 l=2.27
X4 VTAIL.t14 VP.t1 VDD1.t8 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X5 VDD2.t9 VN.t0 VTAIL.t9 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=1.0296 ps=6.57 w=6.24 l=2.27
X6 VDD2.t8 VN.t1 VTAIL.t2 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=2.4336 ps=13.26 w=6.24 l=2.27
X7 VTAIL.t3 VN.t2 VDD2.t7 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X8 VDD1.t7 VP.t2 VTAIL.t17 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=2.4336 ps=13.26 w=6.24 l=2.27
X9 VTAIL.t15 VP.t3 VDD1.t6 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X10 VDD2.t6 VN.t3 VTAIL.t1 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=1.0296 ps=6.57 w=6.24 l=2.27
X11 VDD2.t5 VN.t4 VTAIL.t5 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X12 VDD1.t5 VP.t4 VTAIL.t18 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=1.0296 ps=6.57 w=6.24 l=2.27
X13 VDD1.t4 VP.t5 VTAIL.t19 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X14 VTAIL.t10 VP.t6 VDD1.t3 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X15 VTAIL.t4 VN.t5 VDD2.t4 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X16 VTAIL.t0 VN.t6 VDD2.t3 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X17 VTAIL.t8 VN.t7 VDD2.t2 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X18 VDD1.t2 VP.t7 VTAIL.t12 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X19 VDD2.t1 VN.t8 VTAIL.t7 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=2.4336 ps=13.26 w=6.24 l=2.27
X20 VDD2.t0 VN.t9 VTAIL.t6 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X21 VDD1.t1 VP.t8 VTAIL.t11 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=2.4336 ps=13.26 w=6.24 l=2.27
X22 VTAIL.t13 VP.t9 VDD1.t0 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=1.0296 pd=6.57 as=1.0296 ps=6.57 w=6.24 l=2.27
X23 B.t2 B.t0 B.t1 w_n4090_n2216# sky130_fd_pr__pfet_01v8 ad=2.4336 pd=13.26 as=0 ps=0 w=6.24 l=2.27
R0 B.n512 B.n511 585
R1 B.n513 B.n62 585
R2 B.n515 B.n514 585
R3 B.n516 B.n61 585
R4 B.n518 B.n517 585
R5 B.n519 B.n60 585
R6 B.n521 B.n520 585
R7 B.n522 B.n59 585
R8 B.n524 B.n523 585
R9 B.n525 B.n58 585
R10 B.n527 B.n526 585
R11 B.n528 B.n57 585
R12 B.n530 B.n529 585
R13 B.n531 B.n56 585
R14 B.n533 B.n532 585
R15 B.n534 B.n55 585
R16 B.n536 B.n535 585
R17 B.n537 B.n54 585
R18 B.n539 B.n538 585
R19 B.n540 B.n53 585
R20 B.n542 B.n541 585
R21 B.n543 B.n52 585
R22 B.n545 B.n544 585
R23 B.n546 B.n51 585
R24 B.n548 B.n547 585
R25 B.n550 B.n549 585
R26 B.n551 B.n47 585
R27 B.n553 B.n552 585
R28 B.n554 B.n46 585
R29 B.n556 B.n555 585
R30 B.n557 B.n45 585
R31 B.n559 B.n558 585
R32 B.n560 B.n44 585
R33 B.n562 B.n561 585
R34 B.n564 B.n41 585
R35 B.n566 B.n565 585
R36 B.n567 B.n40 585
R37 B.n569 B.n568 585
R38 B.n570 B.n39 585
R39 B.n572 B.n571 585
R40 B.n573 B.n38 585
R41 B.n575 B.n574 585
R42 B.n576 B.n37 585
R43 B.n578 B.n577 585
R44 B.n579 B.n36 585
R45 B.n581 B.n580 585
R46 B.n582 B.n35 585
R47 B.n584 B.n583 585
R48 B.n585 B.n34 585
R49 B.n587 B.n586 585
R50 B.n588 B.n33 585
R51 B.n590 B.n589 585
R52 B.n591 B.n32 585
R53 B.n593 B.n592 585
R54 B.n594 B.n31 585
R55 B.n596 B.n595 585
R56 B.n597 B.n30 585
R57 B.n599 B.n598 585
R58 B.n600 B.n29 585
R59 B.n510 B.n63 585
R60 B.n509 B.n508 585
R61 B.n507 B.n64 585
R62 B.n506 B.n505 585
R63 B.n504 B.n65 585
R64 B.n503 B.n502 585
R65 B.n501 B.n66 585
R66 B.n500 B.n499 585
R67 B.n498 B.n67 585
R68 B.n497 B.n496 585
R69 B.n495 B.n68 585
R70 B.n494 B.n493 585
R71 B.n492 B.n69 585
R72 B.n491 B.n490 585
R73 B.n489 B.n70 585
R74 B.n488 B.n487 585
R75 B.n486 B.n71 585
R76 B.n485 B.n484 585
R77 B.n483 B.n72 585
R78 B.n482 B.n481 585
R79 B.n480 B.n73 585
R80 B.n479 B.n478 585
R81 B.n477 B.n74 585
R82 B.n476 B.n475 585
R83 B.n474 B.n75 585
R84 B.n473 B.n472 585
R85 B.n471 B.n76 585
R86 B.n470 B.n469 585
R87 B.n468 B.n77 585
R88 B.n467 B.n466 585
R89 B.n465 B.n78 585
R90 B.n464 B.n463 585
R91 B.n462 B.n79 585
R92 B.n461 B.n460 585
R93 B.n459 B.n80 585
R94 B.n458 B.n457 585
R95 B.n456 B.n81 585
R96 B.n455 B.n454 585
R97 B.n453 B.n82 585
R98 B.n452 B.n451 585
R99 B.n450 B.n83 585
R100 B.n449 B.n448 585
R101 B.n447 B.n84 585
R102 B.n446 B.n445 585
R103 B.n444 B.n85 585
R104 B.n443 B.n442 585
R105 B.n441 B.n86 585
R106 B.n440 B.n439 585
R107 B.n438 B.n87 585
R108 B.n437 B.n436 585
R109 B.n435 B.n88 585
R110 B.n434 B.n433 585
R111 B.n432 B.n89 585
R112 B.n431 B.n430 585
R113 B.n429 B.n90 585
R114 B.n428 B.n427 585
R115 B.n426 B.n91 585
R116 B.n425 B.n424 585
R117 B.n423 B.n92 585
R118 B.n422 B.n421 585
R119 B.n420 B.n93 585
R120 B.n419 B.n418 585
R121 B.n417 B.n94 585
R122 B.n416 B.n415 585
R123 B.n414 B.n95 585
R124 B.n413 B.n412 585
R125 B.n411 B.n96 585
R126 B.n410 B.n409 585
R127 B.n408 B.n97 585
R128 B.n407 B.n406 585
R129 B.n405 B.n98 585
R130 B.n404 B.n403 585
R131 B.n402 B.n99 585
R132 B.n401 B.n400 585
R133 B.n399 B.n100 585
R134 B.n398 B.n397 585
R135 B.n396 B.n101 585
R136 B.n395 B.n394 585
R137 B.n393 B.n102 585
R138 B.n392 B.n391 585
R139 B.n390 B.n103 585
R140 B.n389 B.n388 585
R141 B.n387 B.n104 585
R142 B.n386 B.n385 585
R143 B.n384 B.n105 585
R144 B.n383 B.n382 585
R145 B.n381 B.n106 585
R146 B.n380 B.n379 585
R147 B.n378 B.n107 585
R148 B.n377 B.n376 585
R149 B.n375 B.n108 585
R150 B.n374 B.n373 585
R151 B.n372 B.n109 585
R152 B.n371 B.n370 585
R153 B.n369 B.n110 585
R154 B.n368 B.n367 585
R155 B.n366 B.n111 585
R156 B.n365 B.n364 585
R157 B.n363 B.n112 585
R158 B.n362 B.n361 585
R159 B.n360 B.n113 585
R160 B.n359 B.n358 585
R161 B.n357 B.n114 585
R162 B.n356 B.n355 585
R163 B.n354 B.n115 585
R164 B.n353 B.n352 585
R165 B.n351 B.n116 585
R166 B.n350 B.n349 585
R167 B.n348 B.n117 585
R168 B.n258 B.n151 585
R169 B.n260 B.n259 585
R170 B.n261 B.n150 585
R171 B.n263 B.n262 585
R172 B.n264 B.n149 585
R173 B.n266 B.n265 585
R174 B.n267 B.n148 585
R175 B.n269 B.n268 585
R176 B.n270 B.n147 585
R177 B.n272 B.n271 585
R178 B.n273 B.n146 585
R179 B.n275 B.n274 585
R180 B.n276 B.n145 585
R181 B.n278 B.n277 585
R182 B.n279 B.n144 585
R183 B.n281 B.n280 585
R184 B.n282 B.n143 585
R185 B.n284 B.n283 585
R186 B.n285 B.n142 585
R187 B.n287 B.n286 585
R188 B.n288 B.n141 585
R189 B.n290 B.n289 585
R190 B.n291 B.n140 585
R191 B.n293 B.n292 585
R192 B.n294 B.n137 585
R193 B.n297 B.n296 585
R194 B.n298 B.n136 585
R195 B.n300 B.n299 585
R196 B.n301 B.n135 585
R197 B.n303 B.n302 585
R198 B.n304 B.n134 585
R199 B.n306 B.n305 585
R200 B.n307 B.n133 585
R201 B.n309 B.n308 585
R202 B.n311 B.n310 585
R203 B.n312 B.n129 585
R204 B.n314 B.n313 585
R205 B.n315 B.n128 585
R206 B.n317 B.n316 585
R207 B.n318 B.n127 585
R208 B.n320 B.n319 585
R209 B.n321 B.n126 585
R210 B.n323 B.n322 585
R211 B.n324 B.n125 585
R212 B.n326 B.n325 585
R213 B.n327 B.n124 585
R214 B.n329 B.n328 585
R215 B.n330 B.n123 585
R216 B.n332 B.n331 585
R217 B.n333 B.n122 585
R218 B.n335 B.n334 585
R219 B.n336 B.n121 585
R220 B.n338 B.n337 585
R221 B.n339 B.n120 585
R222 B.n341 B.n340 585
R223 B.n342 B.n119 585
R224 B.n344 B.n343 585
R225 B.n345 B.n118 585
R226 B.n347 B.n346 585
R227 B.n257 B.n256 585
R228 B.n255 B.n152 585
R229 B.n254 B.n253 585
R230 B.n252 B.n153 585
R231 B.n251 B.n250 585
R232 B.n249 B.n154 585
R233 B.n248 B.n247 585
R234 B.n246 B.n155 585
R235 B.n245 B.n244 585
R236 B.n243 B.n156 585
R237 B.n242 B.n241 585
R238 B.n240 B.n157 585
R239 B.n239 B.n238 585
R240 B.n237 B.n158 585
R241 B.n236 B.n235 585
R242 B.n234 B.n159 585
R243 B.n233 B.n232 585
R244 B.n231 B.n160 585
R245 B.n230 B.n229 585
R246 B.n228 B.n161 585
R247 B.n227 B.n226 585
R248 B.n225 B.n162 585
R249 B.n224 B.n223 585
R250 B.n222 B.n163 585
R251 B.n221 B.n220 585
R252 B.n219 B.n164 585
R253 B.n218 B.n217 585
R254 B.n216 B.n165 585
R255 B.n215 B.n214 585
R256 B.n213 B.n166 585
R257 B.n212 B.n211 585
R258 B.n210 B.n167 585
R259 B.n209 B.n208 585
R260 B.n207 B.n168 585
R261 B.n206 B.n205 585
R262 B.n204 B.n169 585
R263 B.n203 B.n202 585
R264 B.n201 B.n170 585
R265 B.n200 B.n199 585
R266 B.n198 B.n171 585
R267 B.n197 B.n196 585
R268 B.n195 B.n172 585
R269 B.n194 B.n193 585
R270 B.n192 B.n173 585
R271 B.n191 B.n190 585
R272 B.n189 B.n174 585
R273 B.n188 B.n187 585
R274 B.n186 B.n175 585
R275 B.n185 B.n184 585
R276 B.n183 B.n176 585
R277 B.n182 B.n181 585
R278 B.n180 B.n177 585
R279 B.n179 B.n178 585
R280 B.n2 B.n0 585
R281 B.n681 B.n1 585
R282 B.n680 B.n679 585
R283 B.n678 B.n3 585
R284 B.n677 B.n676 585
R285 B.n675 B.n4 585
R286 B.n674 B.n673 585
R287 B.n672 B.n5 585
R288 B.n671 B.n670 585
R289 B.n669 B.n6 585
R290 B.n668 B.n667 585
R291 B.n666 B.n7 585
R292 B.n665 B.n664 585
R293 B.n663 B.n8 585
R294 B.n662 B.n661 585
R295 B.n660 B.n9 585
R296 B.n659 B.n658 585
R297 B.n657 B.n10 585
R298 B.n656 B.n655 585
R299 B.n654 B.n11 585
R300 B.n653 B.n652 585
R301 B.n651 B.n12 585
R302 B.n650 B.n649 585
R303 B.n648 B.n13 585
R304 B.n647 B.n646 585
R305 B.n645 B.n14 585
R306 B.n644 B.n643 585
R307 B.n642 B.n15 585
R308 B.n641 B.n640 585
R309 B.n639 B.n16 585
R310 B.n638 B.n637 585
R311 B.n636 B.n17 585
R312 B.n635 B.n634 585
R313 B.n633 B.n18 585
R314 B.n632 B.n631 585
R315 B.n630 B.n19 585
R316 B.n629 B.n628 585
R317 B.n627 B.n20 585
R318 B.n626 B.n625 585
R319 B.n624 B.n21 585
R320 B.n623 B.n622 585
R321 B.n621 B.n22 585
R322 B.n620 B.n619 585
R323 B.n618 B.n23 585
R324 B.n617 B.n616 585
R325 B.n615 B.n24 585
R326 B.n614 B.n613 585
R327 B.n612 B.n25 585
R328 B.n611 B.n610 585
R329 B.n609 B.n26 585
R330 B.n608 B.n607 585
R331 B.n606 B.n27 585
R332 B.n605 B.n604 585
R333 B.n603 B.n28 585
R334 B.n602 B.n601 585
R335 B.n683 B.n682 585
R336 B.n256 B.n151 492.5
R337 B.n602 B.n29 492.5
R338 B.n346 B.n117 492.5
R339 B.n512 B.n63 492.5
R340 B.n130 B.t3 273.736
R341 B.n138 B.t9 273.736
R342 B.n42 B.t0 273.736
R343 B.n48 B.t6 273.736
R344 B.n130 B.t5 163.423
R345 B.n48 B.t7 163.423
R346 B.n138 B.t11 163.416
R347 B.n42 B.t1 163.416
R348 B.n256 B.n255 163.367
R349 B.n255 B.n254 163.367
R350 B.n254 B.n153 163.367
R351 B.n250 B.n153 163.367
R352 B.n250 B.n249 163.367
R353 B.n249 B.n248 163.367
R354 B.n248 B.n155 163.367
R355 B.n244 B.n155 163.367
R356 B.n244 B.n243 163.367
R357 B.n243 B.n242 163.367
R358 B.n242 B.n157 163.367
R359 B.n238 B.n157 163.367
R360 B.n238 B.n237 163.367
R361 B.n237 B.n236 163.367
R362 B.n236 B.n159 163.367
R363 B.n232 B.n159 163.367
R364 B.n232 B.n231 163.367
R365 B.n231 B.n230 163.367
R366 B.n230 B.n161 163.367
R367 B.n226 B.n161 163.367
R368 B.n226 B.n225 163.367
R369 B.n225 B.n224 163.367
R370 B.n224 B.n163 163.367
R371 B.n220 B.n163 163.367
R372 B.n220 B.n219 163.367
R373 B.n219 B.n218 163.367
R374 B.n218 B.n165 163.367
R375 B.n214 B.n165 163.367
R376 B.n214 B.n213 163.367
R377 B.n213 B.n212 163.367
R378 B.n212 B.n167 163.367
R379 B.n208 B.n167 163.367
R380 B.n208 B.n207 163.367
R381 B.n207 B.n206 163.367
R382 B.n206 B.n169 163.367
R383 B.n202 B.n169 163.367
R384 B.n202 B.n201 163.367
R385 B.n201 B.n200 163.367
R386 B.n200 B.n171 163.367
R387 B.n196 B.n171 163.367
R388 B.n196 B.n195 163.367
R389 B.n195 B.n194 163.367
R390 B.n194 B.n173 163.367
R391 B.n190 B.n173 163.367
R392 B.n190 B.n189 163.367
R393 B.n189 B.n188 163.367
R394 B.n188 B.n175 163.367
R395 B.n184 B.n175 163.367
R396 B.n184 B.n183 163.367
R397 B.n183 B.n182 163.367
R398 B.n182 B.n177 163.367
R399 B.n178 B.n177 163.367
R400 B.n178 B.n2 163.367
R401 B.n682 B.n2 163.367
R402 B.n682 B.n681 163.367
R403 B.n681 B.n680 163.367
R404 B.n680 B.n3 163.367
R405 B.n676 B.n3 163.367
R406 B.n676 B.n675 163.367
R407 B.n675 B.n674 163.367
R408 B.n674 B.n5 163.367
R409 B.n670 B.n5 163.367
R410 B.n670 B.n669 163.367
R411 B.n669 B.n668 163.367
R412 B.n668 B.n7 163.367
R413 B.n664 B.n7 163.367
R414 B.n664 B.n663 163.367
R415 B.n663 B.n662 163.367
R416 B.n662 B.n9 163.367
R417 B.n658 B.n9 163.367
R418 B.n658 B.n657 163.367
R419 B.n657 B.n656 163.367
R420 B.n656 B.n11 163.367
R421 B.n652 B.n11 163.367
R422 B.n652 B.n651 163.367
R423 B.n651 B.n650 163.367
R424 B.n650 B.n13 163.367
R425 B.n646 B.n13 163.367
R426 B.n646 B.n645 163.367
R427 B.n645 B.n644 163.367
R428 B.n644 B.n15 163.367
R429 B.n640 B.n15 163.367
R430 B.n640 B.n639 163.367
R431 B.n639 B.n638 163.367
R432 B.n638 B.n17 163.367
R433 B.n634 B.n17 163.367
R434 B.n634 B.n633 163.367
R435 B.n633 B.n632 163.367
R436 B.n632 B.n19 163.367
R437 B.n628 B.n19 163.367
R438 B.n628 B.n627 163.367
R439 B.n627 B.n626 163.367
R440 B.n626 B.n21 163.367
R441 B.n622 B.n21 163.367
R442 B.n622 B.n621 163.367
R443 B.n621 B.n620 163.367
R444 B.n620 B.n23 163.367
R445 B.n616 B.n23 163.367
R446 B.n616 B.n615 163.367
R447 B.n615 B.n614 163.367
R448 B.n614 B.n25 163.367
R449 B.n610 B.n25 163.367
R450 B.n610 B.n609 163.367
R451 B.n609 B.n608 163.367
R452 B.n608 B.n27 163.367
R453 B.n604 B.n27 163.367
R454 B.n604 B.n603 163.367
R455 B.n603 B.n602 163.367
R456 B.n260 B.n151 163.367
R457 B.n261 B.n260 163.367
R458 B.n262 B.n261 163.367
R459 B.n262 B.n149 163.367
R460 B.n266 B.n149 163.367
R461 B.n267 B.n266 163.367
R462 B.n268 B.n267 163.367
R463 B.n268 B.n147 163.367
R464 B.n272 B.n147 163.367
R465 B.n273 B.n272 163.367
R466 B.n274 B.n273 163.367
R467 B.n274 B.n145 163.367
R468 B.n278 B.n145 163.367
R469 B.n279 B.n278 163.367
R470 B.n280 B.n279 163.367
R471 B.n280 B.n143 163.367
R472 B.n284 B.n143 163.367
R473 B.n285 B.n284 163.367
R474 B.n286 B.n285 163.367
R475 B.n286 B.n141 163.367
R476 B.n290 B.n141 163.367
R477 B.n291 B.n290 163.367
R478 B.n292 B.n291 163.367
R479 B.n292 B.n137 163.367
R480 B.n297 B.n137 163.367
R481 B.n298 B.n297 163.367
R482 B.n299 B.n298 163.367
R483 B.n299 B.n135 163.367
R484 B.n303 B.n135 163.367
R485 B.n304 B.n303 163.367
R486 B.n305 B.n304 163.367
R487 B.n305 B.n133 163.367
R488 B.n309 B.n133 163.367
R489 B.n310 B.n309 163.367
R490 B.n310 B.n129 163.367
R491 B.n314 B.n129 163.367
R492 B.n315 B.n314 163.367
R493 B.n316 B.n315 163.367
R494 B.n316 B.n127 163.367
R495 B.n320 B.n127 163.367
R496 B.n321 B.n320 163.367
R497 B.n322 B.n321 163.367
R498 B.n322 B.n125 163.367
R499 B.n326 B.n125 163.367
R500 B.n327 B.n326 163.367
R501 B.n328 B.n327 163.367
R502 B.n328 B.n123 163.367
R503 B.n332 B.n123 163.367
R504 B.n333 B.n332 163.367
R505 B.n334 B.n333 163.367
R506 B.n334 B.n121 163.367
R507 B.n338 B.n121 163.367
R508 B.n339 B.n338 163.367
R509 B.n340 B.n339 163.367
R510 B.n340 B.n119 163.367
R511 B.n344 B.n119 163.367
R512 B.n345 B.n344 163.367
R513 B.n346 B.n345 163.367
R514 B.n350 B.n117 163.367
R515 B.n351 B.n350 163.367
R516 B.n352 B.n351 163.367
R517 B.n352 B.n115 163.367
R518 B.n356 B.n115 163.367
R519 B.n357 B.n356 163.367
R520 B.n358 B.n357 163.367
R521 B.n358 B.n113 163.367
R522 B.n362 B.n113 163.367
R523 B.n363 B.n362 163.367
R524 B.n364 B.n363 163.367
R525 B.n364 B.n111 163.367
R526 B.n368 B.n111 163.367
R527 B.n369 B.n368 163.367
R528 B.n370 B.n369 163.367
R529 B.n370 B.n109 163.367
R530 B.n374 B.n109 163.367
R531 B.n375 B.n374 163.367
R532 B.n376 B.n375 163.367
R533 B.n376 B.n107 163.367
R534 B.n380 B.n107 163.367
R535 B.n381 B.n380 163.367
R536 B.n382 B.n381 163.367
R537 B.n382 B.n105 163.367
R538 B.n386 B.n105 163.367
R539 B.n387 B.n386 163.367
R540 B.n388 B.n387 163.367
R541 B.n388 B.n103 163.367
R542 B.n392 B.n103 163.367
R543 B.n393 B.n392 163.367
R544 B.n394 B.n393 163.367
R545 B.n394 B.n101 163.367
R546 B.n398 B.n101 163.367
R547 B.n399 B.n398 163.367
R548 B.n400 B.n399 163.367
R549 B.n400 B.n99 163.367
R550 B.n404 B.n99 163.367
R551 B.n405 B.n404 163.367
R552 B.n406 B.n405 163.367
R553 B.n406 B.n97 163.367
R554 B.n410 B.n97 163.367
R555 B.n411 B.n410 163.367
R556 B.n412 B.n411 163.367
R557 B.n412 B.n95 163.367
R558 B.n416 B.n95 163.367
R559 B.n417 B.n416 163.367
R560 B.n418 B.n417 163.367
R561 B.n418 B.n93 163.367
R562 B.n422 B.n93 163.367
R563 B.n423 B.n422 163.367
R564 B.n424 B.n423 163.367
R565 B.n424 B.n91 163.367
R566 B.n428 B.n91 163.367
R567 B.n429 B.n428 163.367
R568 B.n430 B.n429 163.367
R569 B.n430 B.n89 163.367
R570 B.n434 B.n89 163.367
R571 B.n435 B.n434 163.367
R572 B.n436 B.n435 163.367
R573 B.n436 B.n87 163.367
R574 B.n440 B.n87 163.367
R575 B.n441 B.n440 163.367
R576 B.n442 B.n441 163.367
R577 B.n442 B.n85 163.367
R578 B.n446 B.n85 163.367
R579 B.n447 B.n446 163.367
R580 B.n448 B.n447 163.367
R581 B.n448 B.n83 163.367
R582 B.n452 B.n83 163.367
R583 B.n453 B.n452 163.367
R584 B.n454 B.n453 163.367
R585 B.n454 B.n81 163.367
R586 B.n458 B.n81 163.367
R587 B.n459 B.n458 163.367
R588 B.n460 B.n459 163.367
R589 B.n460 B.n79 163.367
R590 B.n464 B.n79 163.367
R591 B.n465 B.n464 163.367
R592 B.n466 B.n465 163.367
R593 B.n466 B.n77 163.367
R594 B.n470 B.n77 163.367
R595 B.n471 B.n470 163.367
R596 B.n472 B.n471 163.367
R597 B.n472 B.n75 163.367
R598 B.n476 B.n75 163.367
R599 B.n477 B.n476 163.367
R600 B.n478 B.n477 163.367
R601 B.n478 B.n73 163.367
R602 B.n482 B.n73 163.367
R603 B.n483 B.n482 163.367
R604 B.n484 B.n483 163.367
R605 B.n484 B.n71 163.367
R606 B.n488 B.n71 163.367
R607 B.n489 B.n488 163.367
R608 B.n490 B.n489 163.367
R609 B.n490 B.n69 163.367
R610 B.n494 B.n69 163.367
R611 B.n495 B.n494 163.367
R612 B.n496 B.n495 163.367
R613 B.n496 B.n67 163.367
R614 B.n500 B.n67 163.367
R615 B.n501 B.n500 163.367
R616 B.n502 B.n501 163.367
R617 B.n502 B.n65 163.367
R618 B.n506 B.n65 163.367
R619 B.n507 B.n506 163.367
R620 B.n508 B.n507 163.367
R621 B.n508 B.n63 163.367
R622 B.n598 B.n29 163.367
R623 B.n598 B.n597 163.367
R624 B.n597 B.n596 163.367
R625 B.n596 B.n31 163.367
R626 B.n592 B.n31 163.367
R627 B.n592 B.n591 163.367
R628 B.n591 B.n590 163.367
R629 B.n590 B.n33 163.367
R630 B.n586 B.n33 163.367
R631 B.n586 B.n585 163.367
R632 B.n585 B.n584 163.367
R633 B.n584 B.n35 163.367
R634 B.n580 B.n35 163.367
R635 B.n580 B.n579 163.367
R636 B.n579 B.n578 163.367
R637 B.n578 B.n37 163.367
R638 B.n574 B.n37 163.367
R639 B.n574 B.n573 163.367
R640 B.n573 B.n572 163.367
R641 B.n572 B.n39 163.367
R642 B.n568 B.n39 163.367
R643 B.n568 B.n567 163.367
R644 B.n567 B.n566 163.367
R645 B.n566 B.n41 163.367
R646 B.n561 B.n41 163.367
R647 B.n561 B.n560 163.367
R648 B.n560 B.n559 163.367
R649 B.n559 B.n45 163.367
R650 B.n555 B.n45 163.367
R651 B.n555 B.n554 163.367
R652 B.n554 B.n553 163.367
R653 B.n553 B.n47 163.367
R654 B.n549 B.n47 163.367
R655 B.n549 B.n548 163.367
R656 B.n548 B.n51 163.367
R657 B.n544 B.n51 163.367
R658 B.n544 B.n543 163.367
R659 B.n543 B.n542 163.367
R660 B.n542 B.n53 163.367
R661 B.n538 B.n53 163.367
R662 B.n538 B.n537 163.367
R663 B.n537 B.n536 163.367
R664 B.n536 B.n55 163.367
R665 B.n532 B.n55 163.367
R666 B.n532 B.n531 163.367
R667 B.n531 B.n530 163.367
R668 B.n530 B.n57 163.367
R669 B.n526 B.n57 163.367
R670 B.n526 B.n525 163.367
R671 B.n525 B.n524 163.367
R672 B.n524 B.n59 163.367
R673 B.n520 B.n59 163.367
R674 B.n520 B.n519 163.367
R675 B.n519 B.n518 163.367
R676 B.n518 B.n61 163.367
R677 B.n514 B.n61 163.367
R678 B.n514 B.n513 163.367
R679 B.n513 B.n512 163.367
R680 B.n131 B.t4 112.999
R681 B.n49 B.t8 112.999
R682 B.n139 B.t10 112.992
R683 B.n43 B.t2 112.992
R684 B.n132 B.n131 59.5399
R685 B.n295 B.n139 59.5399
R686 B.n563 B.n43 59.5399
R687 B.n50 B.n49 59.5399
R688 B.n131 B.n130 50.4247
R689 B.n139 B.n138 50.4247
R690 B.n43 B.n42 50.4247
R691 B.n49 B.n48 50.4247
R692 B.n601 B.n600 32.0005
R693 B.n511 B.n510 32.0005
R694 B.n348 B.n347 32.0005
R695 B.n258 B.n257 32.0005
R696 B B.n683 18.0485
R697 B.n600 B.n599 10.6151
R698 B.n599 B.n30 10.6151
R699 B.n595 B.n30 10.6151
R700 B.n595 B.n594 10.6151
R701 B.n594 B.n593 10.6151
R702 B.n593 B.n32 10.6151
R703 B.n589 B.n32 10.6151
R704 B.n589 B.n588 10.6151
R705 B.n588 B.n587 10.6151
R706 B.n587 B.n34 10.6151
R707 B.n583 B.n34 10.6151
R708 B.n583 B.n582 10.6151
R709 B.n582 B.n581 10.6151
R710 B.n581 B.n36 10.6151
R711 B.n577 B.n36 10.6151
R712 B.n577 B.n576 10.6151
R713 B.n576 B.n575 10.6151
R714 B.n575 B.n38 10.6151
R715 B.n571 B.n38 10.6151
R716 B.n571 B.n570 10.6151
R717 B.n570 B.n569 10.6151
R718 B.n569 B.n40 10.6151
R719 B.n565 B.n40 10.6151
R720 B.n565 B.n564 10.6151
R721 B.n562 B.n44 10.6151
R722 B.n558 B.n44 10.6151
R723 B.n558 B.n557 10.6151
R724 B.n557 B.n556 10.6151
R725 B.n556 B.n46 10.6151
R726 B.n552 B.n46 10.6151
R727 B.n552 B.n551 10.6151
R728 B.n551 B.n550 10.6151
R729 B.n547 B.n546 10.6151
R730 B.n546 B.n545 10.6151
R731 B.n545 B.n52 10.6151
R732 B.n541 B.n52 10.6151
R733 B.n541 B.n540 10.6151
R734 B.n540 B.n539 10.6151
R735 B.n539 B.n54 10.6151
R736 B.n535 B.n54 10.6151
R737 B.n535 B.n534 10.6151
R738 B.n534 B.n533 10.6151
R739 B.n533 B.n56 10.6151
R740 B.n529 B.n56 10.6151
R741 B.n529 B.n528 10.6151
R742 B.n528 B.n527 10.6151
R743 B.n527 B.n58 10.6151
R744 B.n523 B.n58 10.6151
R745 B.n523 B.n522 10.6151
R746 B.n522 B.n521 10.6151
R747 B.n521 B.n60 10.6151
R748 B.n517 B.n60 10.6151
R749 B.n517 B.n516 10.6151
R750 B.n516 B.n515 10.6151
R751 B.n515 B.n62 10.6151
R752 B.n511 B.n62 10.6151
R753 B.n349 B.n348 10.6151
R754 B.n349 B.n116 10.6151
R755 B.n353 B.n116 10.6151
R756 B.n354 B.n353 10.6151
R757 B.n355 B.n354 10.6151
R758 B.n355 B.n114 10.6151
R759 B.n359 B.n114 10.6151
R760 B.n360 B.n359 10.6151
R761 B.n361 B.n360 10.6151
R762 B.n361 B.n112 10.6151
R763 B.n365 B.n112 10.6151
R764 B.n366 B.n365 10.6151
R765 B.n367 B.n366 10.6151
R766 B.n367 B.n110 10.6151
R767 B.n371 B.n110 10.6151
R768 B.n372 B.n371 10.6151
R769 B.n373 B.n372 10.6151
R770 B.n373 B.n108 10.6151
R771 B.n377 B.n108 10.6151
R772 B.n378 B.n377 10.6151
R773 B.n379 B.n378 10.6151
R774 B.n379 B.n106 10.6151
R775 B.n383 B.n106 10.6151
R776 B.n384 B.n383 10.6151
R777 B.n385 B.n384 10.6151
R778 B.n385 B.n104 10.6151
R779 B.n389 B.n104 10.6151
R780 B.n390 B.n389 10.6151
R781 B.n391 B.n390 10.6151
R782 B.n391 B.n102 10.6151
R783 B.n395 B.n102 10.6151
R784 B.n396 B.n395 10.6151
R785 B.n397 B.n396 10.6151
R786 B.n397 B.n100 10.6151
R787 B.n401 B.n100 10.6151
R788 B.n402 B.n401 10.6151
R789 B.n403 B.n402 10.6151
R790 B.n403 B.n98 10.6151
R791 B.n407 B.n98 10.6151
R792 B.n408 B.n407 10.6151
R793 B.n409 B.n408 10.6151
R794 B.n409 B.n96 10.6151
R795 B.n413 B.n96 10.6151
R796 B.n414 B.n413 10.6151
R797 B.n415 B.n414 10.6151
R798 B.n415 B.n94 10.6151
R799 B.n419 B.n94 10.6151
R800 B.n420 B.n419 10.6151
R801 B.n421 B.n420 10.6151
R802 B.n421 B.n92 10.6151
R803 B.n425 B.n92 10.6151
R804 B.n426 B.n425 10.6151
R805 B.n427 B.n426 10.6151
R806 B.n427 B.n90 10.6151
R807 B.n431 B.n90 10.6151
R808 B.n432 B.n431 10.6151
R809 B.n433 B.n432 10.6151
R810 B.n433 B.n88 10.6151
R811 B.n437 B.n88 10.6151
R812 B.n438 B.n437 10.6151
R813 B.n439 B.n438 10.6151
R814 B.n439 B.n86 10.6151
R815 B.n443 B.n86 10.6151
R816 B.n444 B.n443 10.6151
R817 B.n445 B.n444 10.6151
R818 B.n445 B.n84 10.6151
R819 B.n449 B.n84 10.6151
R820 B.n450 B.n449 10.6151
R821 B.n451 B.n450 10.6151
R822 B.n451 B.n82 10.6151
R823 B.n455 B.n82 10.6151
R824 B.n456 B.n455 10.6151
R825 B.n457 B.n456 10.6151
R826 B.n457 B.n80 10.6151
R827 B.n461 B.n80 10.6151
R828 B.n462 B.n461 10.6151
R829 B.n463 B.n462 10.6151
R830 B.n463 B.n78 10.6151
R831 B.n467 B.n78 10.6151
R832 B.n468 B.n467 10.6151
R833 B.n469 B.n468 10.6151
R834 B.n469 B.n76 10.6151
R835 B.n473 B.n76 10.6151
R836 B.n474 B.n473 10.6151
R837 B.n475 B.n474 10.6151
R838 B.n475 B.n74 10.6151
R839 B.n479 B.n74 10.6151
R840 B.n480 B.n479 10.6151
R841 B.n481 B.n480 10.6151
R842 B.n481 B.n72 10.6151
R843 B.n485 B.n72 10.6151
R844 B.n486 B.n485 10.6151
R845 B.n487 B.n486 10.6151
R846 B.n487 B.n70 10.6151
R847 B.n491 B.n70 10.6151
R848 B.n492 B.n491 10.6151
R849 B.n493 B.n492 10.6151
R850 B.n493 B.n68 10.6151
R851 B.n497 B.n68 10.6151
R852 B.n498 B.n497 10.6151
R853 B.n499 B.n498 10.6151
R854 B.n499 B.n66 10.6151
R855 B.n503 B.n66 10.6151
R856 B.n504 B.n503 10.6151
R857 B.n505 B.n504 10.6151
R858 B.n505 B.n64 10.6151
R859 B.n509 B.n64 10.6151
R860 B.n510 B.n509 10.6151
R861 B.n259 B.n258 10.6151
R862 B.n259 B.n150 10.6151
R863 B.n263 B.n150 10.6151
R864 B.n264 B.n263 10.6151
R865 B.n265 B.n264 10.6151
R866 B.n265 B.n148 10.6151
R867 B.n269 B.n148 10.6151
R868 B.n270 B.n269 10.6151
R869 B.n271 B.n270 10.6151
R870 B.n271 B.n146 10.6151
R871 B.n275 B.n146 10.6151
R872 B.n276 B.n275 10.6151
R873 B.n277 B.n276 10.6151
R874 B.n277 B.n144 10.6151
R875 B.n281 B.n144 10.6151
R876 B.n282 B.n281 10.6151
R877 B.n283 B.n282 10.6151
R878 B.n283 B.n142 10.6151
R879 B.n287 B.n142 10.6151
R880 B.n288 B.n287 10.6151
R881 B.n289 B.n288 10.6151
R882 B.n289 B.n140 10.6151
R883 B.n293 B.n140 10.6151
R884 B.n294 B.n293 10.6151
R885 B.n296 B.n136 10.6151
R886 B.n300 B.n136 10.6151
R887 B.n301 B.n300 10.6151
R888 B.n302 B.n301 10.6151
R889 B.n302 B.n134 10.6151
R890 B.n306 B.n134 10.6151
R891 B.n307 B.n306 10.6151
R892 B.n308 B.n307 10.6151
R893 B.n312 B.n311 10.6151
R894 B.n313 B.n312 10.6151
R895 B.n313 B.n128 10.6151
R896 B.n317 B.n128 10.6151
R897 B.n318 B.n317 10.6151
R898 B.n319 B.n318 10.6151
R899 B.n319 B.n126 10.6151
R900 B.n323 B.n126 10.6151
R901 B.n324 B.n323 10.6151
R902 B.n325 B.n324 10.6151
R903 B.n325 B.n124 10.6151
R904 B.n329 B.n124 10.6151
R905 B.n330 B.n329 10.6151
R906 B.n331 B.n330 10.6151
R907 B.n331 B.n122 10.6151
R908 B.n335 B.n122 10.6151
R909 B.n336 B.n335 10.6151
R910 B.n337 B.n336 10.6151
R911 B.n337 B.n120 10.6151
R912 B.n341 B.n120 10.6151
R913 B.n342 B.n341 10.6151
R914 B.n343 B.n342 10.6151
R915 B.n343 B.n118 10.6151
R916 B.n347 B.n118 10.6151
R917 B.n257 B.n152 10.6151
R918 B.n253 B.n152 10.6151
R919 B.n253 B.n252 10.6151
R920 B.n252 B.n251 10.6151
R921 B.n251 B.n154 10.6151
R922 B.n247 B.n154 10.6151
R923 B.n247 B.n246 10.6151
R924 B.n246 B.n245 10.6151
R925 B.n245 B.n156 10.6151
R926 B.n241 B.n156 10.6151
R927 B.n241 B.n240 10.6151
R928 B.n240 B.n239 10.6151
R929 B.n239 B.n158 10.6151
R930 B.n235 B.n158 10.6151
R931 B.n235 B.n234 10.6151
R932 B.n234 B.n233 10.6151
R933 B.n233 B.n160 10.6151
R934 B.n229 B.n160 10.6151
R935 B.n229 B.n228 10.6151
R936 B.n228 B.n227 10.6151
R937 B.n227 B.n162 10.6151
R938 B.n223 B.n162 10.6151
R939 B.n223 B.n222 10.6151
R940 B.n222 B.n221 10.6151
R941 B.n221 B.n164 10.6151
R942 B.n217 B.n164 10.6151
R943 B.n217 B.n216 10.6151
R944 B.n216 B.n215 10.6151
R945 B.n215 B.n166 10.6151
R946 B.n211 B.n166 10.6151
R947 B.n211 B.n210 10.6151
R948 B.n210 B.n209 10.6151
R949 B.n209 B.n168 10.6151
R950 B.n205 B.n168 10.6151
R951 B.n205 B.n204 10.6151
R952 B.n204 B.n203 10.6151
R953 B.n203 B.n170 10.6151
R954 B.n199 B.n170 10.6151
R955 B.n199 B.n198 10.6151
R956 B.n198 B.n197 10.6151
R957 B.n197 B.n172 10.6151
R958 B.n193 B.n172 10.6151
R959 B.n193 B.n192 10.6151
R960 B.n192 B.n191 10.6151
R961 B.n191 B.n174 10.6151
R962 B.n187 B.n174 10.6151
R963 B.n187 B.n186 10.6151
R964 B.n186 B.n185 10.6151
R965 B.n185 B.n176 10.6151
R966 B.n181 B.n176 10.6151
R967 B.n181 B.n180 10.6151
R968 B.n180 B.n179 10.6151
R969 B.n179 B.n0 10.6151
R970 B.n679 B.n1 10.6151
R971 B.n679 B.n678 10.6151
R972 B.n678 B.n677 10.6151
R973 B.n677 B.n4 10.6151
R974 B.n673 B.n4 10.6151
R975 B.n673 B.n672 10.6151
R976 B.n672 B.n671 10.6151
R977 B.n671 B.n6 10.6151
R978 B.n667 B.n6 10.6151
R979 B.n667 B.n666 10.6151
R980 B.n666 B.n665 10.6151
R981 B.n665 B.n8 10.6151
R982 B.n661 B.n8 10.6151
R983 B.n661 B.n660 10.6151
R984 B.n660 B.n659 10.6151
R985 B.n659 B.n10 10.6151
R986 B.n655 B.n10 10.6151
R987 B.n655 B.n654 10.6151
R988 B.n654 B.n653 10.6151
R989 B.n653 B.n12 10.6151
R990 B.n649 B.n12 10.6151
R991 B.n649 B.n648 10.6151
R992 B.n648 B.n647 10.6151
R993 B.n647 B.n14 10.6151
R994 B.n643 B.n14 10.6151
R995 B.n643 B.n642 10.6151
R996 B.n642 B.n641 10.6151
R997 B.n641 B.n16 10.6151
R998 B.n637 B.n16 10.6151
R999 B.n637 B.n636 10.6151
R1000 B.n636 B.n635 10.6151
R1001 B.n635 B.n18 10.6151
R1002 B.n631 B.n18 10.6151
R1003 B.n631 B.n630 10.6151
R1004 B.n630 B.n629 10.6151
R1005 B.n629 B.n20 10.6151
R1006 B.n625 B.n20 10.6151
R1007 B.n625 B.n624 10.6151
R1008 B.n624 B.n623 10.6151
R1009 B.n623 B.n22 10.6151
R1010 B.n619 B.n22 10.6151
R1011 B.n619 B.n618 10.6151
R1012 B.n618 B.n617 10.6151
R1013 B.n617 B.n24 10.6151
R1014 B.n613 B.n24 10.6151
R1015 B.n613 B.n612 10.6151
R1016 B.n612 B.n611 10.6151
R1017 B.n611 B.n26 10.6151
R1018 B.n607 B.n26 10.6151
R1019 B.n607 B.n606 10.6151
R1020 B.n606 B.n605 10.6151
R1021 B.n605 B.n28 10.6151
R1022 B.n601 B.n28 10.6151
R1023 B.n563 B.n562 6.5566
R1024 B.n550 B.n50 6.5566
R1025 B.n296 B.n295 6.5566
R1026 B.n308 B.n132 6.5566
R1027 B.n564 B.n563 4.05904
R1028 B.n547 B.n50 4.05904
R1029 B.n295 B.n294 4.05904
R1030 B.n311 B.n132 4.05904
R1031 B.n683 B.n0 2.81026
R1032 B.n683 B.n1 2.81026
R1033 VP.n22 VP.n21 161.3
R1034 VP.n23 VP.n18 161.3
R1035 VP.n25 VP.n24 161.3
R1036 VP.n26 VP.n17 161.3
R1037 VP.n28 VP.n27 161.3
R1038 VP.n29 VP.n16 161.3
R1039 VP.n31 VP.n30 161.3
R1040 VP.n32 VP.n15 161.3
R1041 VP.n34 VP.n33 161.3
R1042 VP.n35 VP.n14 161.3
R1043 VP.n37 VP.n36 161.3
R1044 VP.n39 VP.n13 161.3
R1045 VP.n41 VP.n40 161.3
R1046 VP.n42 VP.n12 161.3
R1047 VP.n44 VP.n43 161.3
R1048 VP.n45 VP.n11 161.3
R1049 VP.n82 VP.n0 161.3
R1050 VP.n81 VP.n80 161.3
R1051 VP.n79 VP.n1 161.3
R1052 VP.n78 VP.n77 161.3
R1053 VP.n76 VP.n2 161.3
R1054 VP.n74 VP.n73 161.3
R1055 VP.n72 VP.n3 161.3
R1056 VP.n71 VP.n70 161.3
R1057 VP.n69 VP.n4 161.3
R1058 VP.n68 VP.n67 161.3
R1059 VP.n66 VP.n5 161.3
R1060 VP.n65 VP.n64 161.3
R1061 VP.n63 VP.n6 161.3
R1062 VP.n62 VP.n61 161.3
R1063 VP.n60 VP.n7 161.3
R1064 VP.n59 VP.n58 161.3
R1065 VP.n56 VP.n8 161.3
R1066 VP.n55 VP.n54 161.3
R1067 VP.n53 VP.n9 161.3
R1068 VP.n52 VP.n51 161.3
R1069 VP.n50 VP.n10 161.3
R1070 VP.n49 VP.n48 101.072
R1071 VP.n84 VP.n83 101.072
R1072 VP.n47 VP.n46 101.072
R1073 VP.n19 VP.t4 97.2042
R1074 VP.n20 VP.n19 67.3861
R1075 VP.n5 VP.t7 66.249
R1076 VP.n49 VP.t0 66.249
R1077 VP.n57 VP.t1 66.249
R1078 VP.n75 VP.t9 66.249
R1079 VP.n83 VP.t8 66.249
R1080 VP.n16 VP.t5 66.249
R1081 VP.n46 VP.t2 66.249
R1082 VP.n38 VP.t3 66.249
R1083 VP.n20 VP.t6 66.249
R1084 VP.n63 VP.n62 56.5617
R1085 VP.n70 VP.n69 56.5617
R1086 VP.n33 VP.n32 56.5617
R1087 VP.n26 VP.n25 56.5617
R1088 VP.n55 VP.n9 50.2647
R1089 VP.n77 VP.n1 50.2647
R1090 VP.n40 VP.n12 50.2647
R1091 VP.n48 VP.n47 46.8936
R1092 VP.n51 VP.n9 30.8893
R1093 VP.n81 VP.n1 30.8893
R1094 VP.n44 VP.n12 30.8893
R1095 VP.n51 VP.n50 24.5923
R1096 VP.n56 VP.n55 24.5923
R1097 VP.n58 VP.n7 24.5923
R1098 VP.n62 VP.n7 24.5923
R1099 VP.n64 VP.n63 24.5923
R1100 VP.n64 VP.n5 24.5923
R1101 VP.n68 VP.n5 24.5923
R1102 VP.n69 VP.n68 24.5923
R1103 VP.n70 VP.n3 24.5923
R1104 VP.n74 VP.n3 24.5923
R1105 VP.n77 VP.n76 24.5923
R1106 VP.n82 VP.n81 24.5923
R1107 VP.n45 VP.n44 24.5923
R1108 VP.n33 VP.n14 24.5923
R1109 VP.n37 VP.n14 24.5923
R1110 VP.n40 VP.n39 24.5923
R1111 VP.n27 VP.n26 24.5923
R1112 VP.n27 VP.n16 24.5923
R1113 VP.n31 VP.n16 24.5923
R1114 VP.n32 VP.n31 24.5923
R1115 VP.n21 VP.n18 24.5923
R1116 VP.n25 VP.n18 24.5923
R1117 VP.n57 VP.n56 19.674
R1118 VP.n76 VP.n75 19.674
R1119 VP.n39 VP.n38 19.674
R1120 VP.n22 VP.n19 10.0049
R1121 VP.n50 VP.n49 9.83723
R1122 VP.n83 VP.n82 9.83723
R1123 VP.n46 VP.n45 9.83723
R1124 VP.n58 VP.n57 4.91887
R1125 VP.n75 VP.n74 4.91887
R1126 VP.n38 VP.n37 4.91887
R1127 VP.n21 VP.n20 4.91887
R1128 VP.n47 VP.n11 0.278335
R1129 VP.n48 VP.n10 0.278335
R1130 VP.n84 VP.n0 0.278335
R1131 VP.n23 VP.n22 0.189894
R1132 VP.n24 VP.n23 0.189894
R1133 VP.n24 VP.n17 0.189894
R1134 VP.n28 VP.n17 0.189894
R1135 VP.n29 VP.n28 0.189894
R1136 VP.n30 VP.n29 0.189894
R1137 VP.n30 VP.n15 0.189894
R1138 VP.n34 VP.n15 0.189894
R1139 VP.n35 VP.n34 0.189894
R1140 VP.n36 VP.n35 0.189894
R1141 VP.n36 VP.n13 0.189894
R1142 VP.n41 VP.n13 0.189894
R1143 VP.n42 VP.n41 0.189894
R1144 VP.n43 VP.n42 0.189894
R1145 VP.n43 VP.n11 0.189894
R1146 VP.n52 VP.n10 0.189894
R1147 VP.n53 VP.n52 0.189894
R1148 VP.n54 VP.n53 0.189894
R1149 VP.n54 VP.n8 0.189894
R1150 VP.n59 VP.n8 0.189894
R1151 VP.n60 VP.n59 0.189894
R1152 VP.n61 VP.n60 0.189894
R1153 VP.n61 VP.n6 0.189894
R1154 VP.n65 VP.n6 0.189894
R1155 VP.n66 VP.n65 0.189894
R1156 VP.n67 VP.n66 0.189894
R1157 VP.n67 VP.n4 0.189894
R1158 VP.n71 VP.n4 0.189894
R1159 VP.n72 VP.n71 0.189894
R1160 VP.n73 VP.n72 0.189894
R1161 VP.n73 VP.n2 0.189894
R1162 VP.n78 VP.n2 0.189894
R1163 VP.n79 VP.n78 0.189894
R1164 VP.n80 VP.n79 0.189894
R1165 VP.n80 VP.n0 0.189894
R1166 VP VP.n84 0.153485
R1167 VTAIL.n11 VTAIL.t2 76.4315
R1168 VTAIL.n17 VTAIL.t7 76.4314
R1169 VTAIL.n2 VTAIL.t11 76.4314
R1170 VTAIL.n16 VTAIL.t17 76.4313
R1171 VTAIL.n15 VTAIL.n14 71.2224
R1172 VTAIL.n13 VTAIL.n12 71.2224
R1173 VTAIL.n10 VTAIL.n9 71.2224
R1174 VTAIL.n8 VTAIL.n7 71.2224
R1175 VTAIL.n19 VTAIL.n18 71.2222
R1176 VTAIL.n1 VTAIL.n0 71.2222
R1177 VTAIL.n4 VTAIL.n3 71.2222
R1178 VTAIL.n6 VTAIL.n5 71.2222
R1179 VTAIL.n8 VTAIL.n6 22.2289
R1180 VTAIL.n17 VTAIL.n16 19.9876
R1181 VTAIL.n18 VTAIL.t6 5.20963
R1182 VTAIL.n18 VTAIL.t0 5.20963
R1183 VTAIL.n0 VTAIL.t9 5.20963
R1184 VTAIL.n0 VTAIL.t8 5.20963
R1185 VTAIL.n3 VTAIL.t12 5.20963
R1186 VTAIL.n3 VTAIL.t13 5.20963
R1187 VTAIL.n5 VTAIL.t16 5.20963
R1188 VTAIL.n5 VTAIL.t14 5.20963
R1189 VTAIL.n14 VTAIL.t19 5.20963
R1190 VTAIL.n14 VTAIL.t15 5.20963
R1191 VTAIL.n12 VTAIL.t18 5.20963
R1192 VTAIL.n12 VTAIL.t10 5.20963
R1193 VTAIL.n9 VTAIL.t5 5.20963
R1194 VTAIL.n9 VTAIL.t3 5.20963
R1195 VTAIL.n7 VTAIL.t1 5.20963
R1196 VTAIL.n7 VTAIL.t4 5.20963
R1197 VTAIL.n10 VTAIL.n8 2.24188
R1198 VTAIL.n11 VTAIL.n10 2.24188
R1199 VTAIL.n15 VTAIL.n13 2.24188
R1200 VTAIL.n16 VTAIL.n15 2.24188
R1201 VTAIL.n6 VTAIL.n4 2.24188
R1202 VTAIL.n4 VTAIL.n2 2.24188
R1203 VTAIL.n19 VTAIL.n17 2.24188
R1204 VTAIL VTAIL.n1 1.73972
R1205 VTAIL.n13 VTAIL.n11 1.59102
R1206 VTAIL.n2 VTAIL.n1 1.59102
R1207 VTAIL VTAIL.n19 0.502655
R1208 VDD1.n1 VDD1.t5 95.3516
R1209 VDD1.n3 VDD1.t9 95.3515
R1210 VDD1.n5 VDD1.n4 89.5266
R1211 VDD1.n1 VDD1.n0 87.9012
R1212 VDD1.n7 VDD1.n6 87.901
R1213 VDD1.n3 VDD1.n2 87.901
R1214 VDD1.n7 VDD1.n5 41.4449
R1215 VDD1.n6 VDD1.t6 5.20963
R1216 VDD1.n6 VDD1.t7 5.20963
R1217 VDD1.n0 VDD1.t3 5.20963
R1218 VDD1.n0 VDD1.t4 5.20963
R1219 VDD1.n4 VDD1.t0 5.20963
R1220 VDD1.n4 VDD1.t1 5.20963
R1221 VDD1.n2 VDD1.t8 5.20963
R1222 VDD1.n2 VDD1.t2 5.20963
R1223 VDD1 VDD1.n7 1.62334
R1224 VDD1 VDD1.n1 0.619035
R1225 VDD1.n5 VDD1.n3 0.505499
R1226 VN.n71 VN.n37 161.3
R1227 VN.n70 VN.n69 161.3
R1228 VN.n68 VN.n38 161.3
R1229 VN.n67 VN.n66 161.3
R1230 VN.n65 VN.n39 161.3
R1231 VN.n63 VN.n62 161.3
R1232 VN.n61 VN.n40 161.3
R1233 VN.n60 VN.n59 161.3
R1234 VN.n58 VN.n41 161.3
R1235 VN.n57 VN.n56 161.3
R1236 VN.n55 VN.n42 161.3
R1237 VN.n54 VN.n53 161.3
R1238 VN.n52 VN.n43 161.3
R1239 VN.n51 VN.n50 161.3
R1240 VN.n49 VN.n44 161.3
R1241 VN.n48 VN.n47 161.3
R1242 VN.n34 VN.n0 161.3
R1243 VN.n33 VN.n32 161.3
R1244 VN.n31 VN.n1 161.3
R1245 VN.n30 VN.n29 161.3
R1246 VN.n28 VN.n2 161.3
R1247 VN.n26 VN.n25 161.3
R1248 VN.n24 VN.n3 161.3
R1249 VN.n23 VN.n22 161.3
R1250 VN.n21 VN.n4 161.3
R1251 VN.n20 VN.n19 161.3
R1252 VN.n18 VN.n5 161.3
R1253 VN.n17 VN.n16 161.3
R1254 VN.n15 VN.n6 161.3
R1255 VN.n14 VN.n13 161.3
R1256 VN.n12 VN.n7 161.3
R1257 VN.n11 VN.n10 161.3
R1258 VN.n36 VN.n35 101.072
R1259 VN.n73 VN.n72 101.072
R1260 VN.n8 VN.t0 97.2042
R1261 VN.n45 VN.t1 97.2042
R1262 VN.n9 VN.n8 67.3861
R1263 VN.n46 VN.n45 67.3861
R1264 VN.n5 VN.t9 66.249
R1265 VN.n9 VN.t7 66.249
R1266 VN.n27 VN.t6 66.249
R1267 VN.n35 VN.t8 66.249
R1268 VN.n42 VN.t4 66.249
R1269 VN.n46 VN.t2 66.249
R1270 VN.n64 VN.t5 66.249
R1271 VN.n72 VN.t3 66.249
R1272 VN.n15 VN.n14 56.5617
R1273 VN.n22 VN.n21 56.5617
R1274 VN.n52 VN.n51 56.5617
R1275 VN.n59 VN.n58 56.5617
R1276 VN.n29 VN.n1 50.2647
R1277 VN.n66 VN.n38 50.2647
R1278 VN VN.n73 47.1724
R1279 VN.n33 VN.n1 30.8893
R1280 VN.n70 VN.n38 30.8893
R1281 VN.n10 VN.n7 24.5923
R1282 VN.n14 VN.n7 24.5923
R1283 VN.n16 VN.n15 24.5923
R1284 VN.n16 VN.n5 24.5923
R1285 VN.n20 VN.n5 24.5923
R1286 VN.n21 VN.n20 24.5923
R1287 VN.n22 VN.n3 24.5923
R1288 VN.n26 VN.n3 24.5923
R1289 VN.n29 VN.n28 24.5923
R1290 VN.n34 VN.n33 24.5923
R1291 VN.n51 VN.n44 24.5923
R1292 VN.n47 VN.n44 24.5923
R1293 VN.n58 VN.n57 24.5923
R1294 VN.n57 VN.n42 24.5923
R1295 VN.n53 VN.n42 24.5923
R1296 VN.n53 VN.n52 24.5923
R1297 VN.n66 VN.n65 24.5923
R1298 VN.n63 VN.n40 24.5923
R1299 VN.n59 VN.n40 24.5923
R1300 VN.n71 VN.n70 24.5923
R1301 VN.n28 VN.n27 19.674
R1302 VN.n65 VN.n64 19.674
R1303 VN.n48 VN.n45 10.0049
R1304 VN.n11 VN.n8 10.0049
R1305 VN.n35 VN.n34 9.83723
R1306 VN.n72 VN.n71 9.83723
R1307 VN.n10 VN.n9 4.91887
R1308 VN.n27 VN.n26 4.91887
R1309 VN.n47 VN.n46 4.91887
R1310 VN.n64 VN.n63 4.91887
R1311 VN.n73 VN.n37 0.278335
R1312 VN.n36 VN.n0 0.278335
R1313 VN.n69 VN.n37 0.189894
R1314 VN.n69 VN.n68 0.189894
R1315 VN.n68 VN.n67 0.189894
R1316 VN.n67 VN.n39 0.189894
R1317 VN.n62 VN.n39 0.189894
R1318 VN.n62 VN.n61 0.189894
R1319 VN.n61 VN.n60 0.189894
R1320 VN.n60 VN.n41 0.189894
R1321 VN.n56 VN.n41 0.189894
R1322 VN.n56 VN.n55 0.189894
R1323 VN.n55 VN.n54 0.189894
R1324 VN.n54 VN.n43 0.189894
R1325 VN.n50 VN.n43 0.189894
R1326 VN.n50 VN.n49 0.189894
R1327 VN.n49 VN.n48 0.189894
R1328 VN.n12 VN.n11 0.189894
R1329 VN.n13 VN.n12 0.189894
R1330 VN.n13 VN.n6 0.189894
R1331 VN.n17 VN.n6 0.189894
R1332 VN.n18 VN.n17 0.189894
R1333 VN.n19 VN.n18 0.189894
R1334 VN.n19 VN.n4 0.189894
R1335 VN.n23 VN.n4 0.189894
R1336 VN.n24 VN.n23 0.189894
R1337 VN.n25 VN.n24 0.189894
R1338 VN.n25 VN.n2 0.189894
R1339 VN.n30 VN.n2 0.189894
R1340 VN.n31 VN.n30 0.189894
R1341 VN.n32 VN.n31 0.189894
R1342 VN.n32 VN.n0 0.189894
R1343 VN VN.n36 0.153485
R1344 VDD2.n1 VDD2.t9 95.3515
R1345 VDD2.n4 VDD2.t6 93.1102
R1346 VDD2.n3 VDD2.n2 89.5266
R1347 VDD2 VDD2.n7 89.5238
R1348 VDD2.n6 VDD2.n5 87.9012
R1349 VDD2.n1 VDD2.n0 87.901
R1350 VDD2.n4 VDD2.n3 39.7412
R1351 VDD2.n7 VDD2.t7 5.20963
R1352 VDD2.n7 VDD2.t8 5.20963
R1353 VDD2.n5 VDD2.t4 5.20963
R1354 VDD2.n5 VDD2.t5 5.20963
R1355 VDD2.n2 VDD2.t3 5.20963
R1356 VDD2.n2 VDD2.t1 5.20963
R1357 VDD2.n0 VDD2.t2 5.20963
R1358 VDD2.n0 VDD2.t0 5.20963
R1359 VDD2.n6 VDD2.n4 2.24188
R1360 VDD2 VDD2.n6 0.619035
R1361 VDD2.n3 VDD2.n1 0.505499
C0 VN VDD1 0.152968f
C1 VDD2 B 2.00531f
C2 VTAIL VDD2 7.57848f
C3 w_n4090_n2216# VP 9.074201f
C4 VDD2 VDD1 1.95912f
C5 w_n4090_n2216# B 8.3846f
C6 VTAIL w_n4090_n2216# 2.35179f
C7 w_n4090_n2216# VDD1 2.26088f
C8 VDD2 VN 5.63351f
C9 VP B 2.02399f
C10 VTAIL VP 6.57849f
C11 VP VDD1 6.01914f
C12 VTAIL B 2.32337f
C13 w_n4090_n2216# VN 8.54272f
C14 B VDD1 1.90024f
C15 VTAIL VDD1 7.52862f
C16 w_n4090_n2216# VDD2 2.38737f
C17 VN VP 6.84317f
C18 VN B 1.1321f
C19 VTAIL VN 6.56428f
C20 VDD2 VP 0.541351f
C21 VDD2 VSUBS 1.834705f
C22 VDD1 VSUBS 1.627915f
C23 VTAIL VSUBS 0.646557f
C24 VN VSUBS 6.8394f
C25 VP VSUBS 3.408026f
C26 B VSUBS 4.470204f
C27 w_n4090_n2216# VSUBS 0.113031p
C28 VDD2.t9 VSUBS 1.33689f
C29 VDD2.t2 VSUBS 0.147719f
C30 VDD2.t0 VSUBS 0.147719f
C31 VDD2.n0 VSUBS 0.984704f
C32 VDD2.n1 VSUBS 1.53976f
C33 VDD2.t3 VSUBS 0.147719f
C34 VDD2.t1 VSUBS 0.147719f
C35 VDD2.n2 VSUBS 1.00074f
C36 VDD2.n3 VSUBS 3.10593f
C37 VDD2.t6 VSUBS 1.31821f
C38 VDD2.n4 VSUBS 3.29092f
C39 VDD2.t4 VSUBS 0.147719f
C40 VDD2.t5 VSUBS 0.147719f
C41 VDD2.n5 VSUBS 0.984709f
C42 VDD2.n6 VSUBS 0.773149f
C43 VDD2.t7 VSUBS 0.147719f
C44 VDD2.t8 VSUBS 0.147719f
C45 VDD2.n7 VSUBS 1.0007f
C46 VN.n0 VSUBS 0.048733f
C47 VN.t8 VSUBS 1.38903f
C48 VN.n1 VSUBS 0.034853f
C49 VN.n2 VSUBS 0.036966f
C50 VN.t6 VSUBS 1.38903f
C51 VN.n3 VSUBS 0.06855f
C52 VN.n4 VSUBS 0.036966f
C53 VN.t9 VSUBS 1.38903f
C54 VN.n5 VSUBS 0.55769f
C55 VN.n6 VSUBS 0.036966f
C56 VN.n7 VSUBS 0.06855f
C57 VN.t0 VSUBS 1.61816f
C58 VN.n8 VSUBS 0.609819f
C59 VN.t7 VSUBS 1.38903f
C60 VN.n9 VSUBS 0.611098f
C61 VN.n10 VSUBS 0.041477f
C62 VN.n11 VSUBS 0.316634f
C63 VN.n12 VSUBS 0.036966f
C64 VN.n13 VSUBS 0.036966f
C65 VN.n14 VSUBS 0.048622f
C66 VN.n15 VSUBS 0.05885f
C67 VN.n16 VSUBS 0.06855f
C68 VN.n17 VSUBS 0.036966f
C69 VN.n18 VSUBS 0.036966f
C70 VN.n19 VSUBS 0.036966f
C71 VN.n20 VSUBS 0.06855f
C72 VN.n21 VSUBS 0.05885f
C73 VN.n22 VSUBS 0.048622f
C74 VN.n23 VSUBS 0.036966f
C75 VN.n24 VSUBS 0.036966f
C76 VN.n25 VSUBS 0.036966f
C77 VN.n26 VSUBS 0.041477f
C78 VN.n27 VSUBS 0.522981f
C79 VN.n28 VSUBS 0.061782f
C80 VN.n29 VSUBS 0.067513f
C81 VN.n30 VSUBS 0.036966f
C82 VN.n31 VSUBS 0.036966f
C83 VN.n32 VSUBS 0.036966f
C84 VN.n33 VSUBS 0.073655f
C85 VN.n34 VSUBS 0.048245f
C86 VN.n35 VSUBS 0.629288f
C87 VN.n36 VSUBS 0.056487f
C88 VN.n37 VSUBS 0.048733f
C89 VN.t3 VSUBS 1.38903f
C90 VN.n38 VSUBS 0.034853f
C91 VN.n39 VSUBS 0.036966f
C92 VN.t5 VSUBS 1.38903f
C93 VN.n40 VSUBS 0.06855f
C94 VN.n41 VSUBS 0.036966f
C95 VN.t4 VSUBS 1.38903f
C96 VN.n42 VSUBS 0.55769f
C97 VN.n43 VSUBS 0.036966f
C98 VN.n44 VSUBS 0.06855f
C99 VN.t1 VSUBS 1.61816f
C100 VN.n45 VSUBS 0.609819f
C101 VN.t2 VSUBS 1.38903f
C102 VN.n46 VSUBS 0.611098f
C103 VN.n47 VSUBS 0.041477f
C104 VN.n48 VSUBS 0.316634f
C105 VN.n49 VSUBS 0.036966f
C106 VN.n50 VSUBS 0.036966f
C107 VN.n51 VSUBS 0.048622f
C108 VN.n52 VSUBS 0.05885f
C109 VN.n53 VSUBS 0.06855f
C110 VN.n54 VSUBS 0.036966f
C111 VN.n55 VSUBS 0.036966f
C112 VN.n56 VSUBS 0.036966f
C113 VN.n57 VSUBS 0.06855f
C114 VN.n58 VSUBS 0.05885f
C115 VN.n59 VSUBS 0.048622f
C116 VN.n60 VSUBS 0.036966f
C117 VN.n61 VSUBS 0.036966f
C118 VN.n62 VSUBS 0.036966f
C119 VN.n63 VSUBS 0.041477f
C120 VN.n64 VSUBS 0.522981f
C121 VN.n65 VSUBS 0.061782f
C122 VN.n66 VSUBS 0.067513f
C123 VN.n67 VSUBS 0.036966f
C124 VN.n68 VSUBS 0.036966f
C125 VN.n69 VSUBS 0.036966f
C126 VN.n70 VSUBS 0.073655f
C127 VN.n71 VSUBS 0.048245f
C128 VN.n72 VSUBS 0.629288f
C129 VN.n73 VSUBS 1.88368f
C130 VDD1.t5 VSUBS 1.19267f
C131 VDD1.t3 VSUBS 0.131783f
C132 VDD1.t4 VSUBS 0.131783f
C133 VDD1.n0 VSUBS 0.878477f
C134 VDD1.n1 VSUBS 1.38219f
C135 VDD1.t9 VSUBS 1.19267f
C136 VDD1.t8 VSUBS 0.131783f
C137 VDD1.t2 VSUBS 0.131783f
C138 VDD1.n2 VSUBS 0.878473f
C139 VDD1.n3 VSUBS 1.37365f
C140 VDD1.t0 VSUBS 0.131783f
C141 VDD1.t1 VSUBS 0.131783f
C142 VDD1.n4 VSUBS 0.892776f
C143 VDD1.n5 VSUBS 2.89048f
C144 VDD1.t6 VSUBS 0.131783f
C145 VDD1.t7 VSUBS 0.131783f
C146 VDD1.n6 VSUBS 0.878472f
C147 VDD1.n7 VSUBS 2.99285f
C148 VTAIL.t9 VSUBS 0.160635f
C149 VTAIL.t8 VSUBS 0.160635f
C150 VTAIL.n0 VSUBS 0.945667f
C151 VTAIL.n1 VSUBS 0.97093f
C152 VTAIL.t11 VSUBS 1.3004f
C153 VTAIL.n2 VSUBS 1.107f
C154 VTAIL.t12 VSUBS 0.160635f
C155 VTAIL.t13 VSUBS 0.160635f
C156 VTAIL.n3 VSUBS 0.945667f
C157 VTAIL.n4 VSUBS 1.09196f
C158 VTAIL.t16 VSUBS 0.160635f
C159 VTAIL.t14 VSUBS 0.160635f
C160 VTAIL.n5 VSUBS 0.945667f
C161 VTAIL.n6 VSUBS 2.3344f
C162 VTAIL.t1 VSUBS 0.160635f
C163 VTAIL.t4 VSUBS 0.160635f
C164 VTAIL.n7 VSUBS 0.945673f
C165 VTAIL.n8 VSUBS 2.33439f
C166 VTAIL.t5 VSUBS 0.160635f
C167 VTAIL.t3 VSUBS 0.160635f
C168 VTAIL.n9 VSUBS 0.945673f
C169 VTAIL.n10 VSUBS 1.09195f
C170 VTAIL.t2 VSUBS 1.30041f
C171 VTAIL.n11 VSUBS 1.10699f
C172 VTAIL.t18 VSUBS 0.160635f
C173 VTAIL.t10 VSUBS 0.160635f
C174 VTAIL.n12 VSUBS 0.945673f
C175 VTAIL.n13 VSUBS 1.02363f
C176 VTAIL.t19 VSUBS 0.160635f
C177 VTAIL.t15 VSUBS 0.160635f
C178 VTAIL.n14 VSUBS 0.945673f
C179 VTAIL.n15 VSUBS 1.09195f
C180 VTAIL.t17 VSUBS 1.3004f
C181 VTAIL.n16 VSUBS 2.18249f
C182 VTAIL.t7 VSUBS 1.3004f
C183 VTAIL.n17 VSUBS 2.18249f
C184 VTAIL.t6 VSUBS 0.160635f
C185 VTAIL.t0 VSUBS 0.160635f
C186 VTAIL.n18 VSUBS 0.945667f
C187 VTAIL.n19 VSUBS 0.909397f
C188 VP.n0 VSUBS 0.054152f
C189 VP.t8 VSUBS 1.54348f
C190 VP.n1 VSUBS 0.038729f
C191 VP.n2 VSUBS 0.041076f
C192 VP.t9 VSUBS 1.54348f
C193 VP.n3 VSUBS 0.076172f
C194 VP.n4 VSUBS 0.041076f
C195 VP.t7 VSUBS 1.54348f
C196 VP.n5 VSUBS 0.6197f
C197 VP.n6 VSUBS 0.041076f
C198 VP.n7 VSUBS 0.076172f
C199 VP.n8 VSUBS 0.041076f
C200 VP.t1 VSUBS 1.54348f
C201 VP.n9 VSUBS 0.038729f
C202 VP.n10 VSUBS 0.054152f
C203 VP.t0 VSUBS 1.54348f
C204 VP.n11 VSUBS 0.054152f
C205 VP.t2 VSUBS 1.54348f
C206 VP.n12 VSUBS 0.038729f
C207 VP.n13 VSUBS 0.041076f
C208 VP.t3 VSUBS 1.54348f
C209 VP.n14 VSUBS 0.076172f
C210 VP.n15 VSUBS 0.041076f
C211 VP.t5 VSUBS 1.54348f
C212 VP.n16 VSUBS 0.6197f
C213 VP.n17 VSUBS 0.041076f
C214 VP.n18 VSUBS 0.076172f
C215 VP.t4 VSUBS 1.79809f
C216 VP.n19 VSUBS 0.677625f
C217 VP.t6 VSUBS 1.54348f
C218 VP.n20 VSUBS 0.679047f
C219 VP.n21 VSUBS 0.046089f
C220 VP.n22 VSUBS 0.351841f
C221 VP.n23 VSUBS 0.041076f
C222 VP.n24 VSUBS 0.041076f
C223 VP.n25 VSUBS 0.054028f
C224 VP.n26 VSUBS 0.065393f
C225 VP.n27 VSUBS 0.076172f
C226 VP.n28 VSUBS 0.041076f
C227 VP.n29 VSUBS 0.041076f
C228 VP.n30 VSUBS 0.041076f
C229 VP.n31 VSUBS 0.076172f
C230 VP.n32 VSUBS 0.065393f
C231 VP.n33 VSUBS 0.054028f
C232 VP.n34 VSUBS 0.041076f
C233 VP.n35 VSUBS 0.041076f
C234 VP.n36 VSUBS 0.041076f
C235 VP.n37 VSUBS 0.046089f
C236 VP.n38 VSUBS 0.581132f
C237 VP.n39 VSUBS 0.068651f
C238 VP.n40 VSUBS 0.07502f
C239 VP.n41 VSUBS 0.041076f
C240 VP.n42 VSUBS 0.041076f
C241 VP.n43 VSUBS 0.041076f
C242 VP.n44 VSUBS 0.081845f
C243 VP.n45 VSUBS 0.05361f
C244 VP.n46 VSUBS 0.699259f
C245 VP.n47 VSUBS 2.07082f
C246 VP.n48 VSUBS 2.1024f
C247 VP.n49 VSUBS 0.699259f
C248 VP.n50 VSUBS 0.05361f
C249 VP.n51 VSUBS 0.081845f
C250 VP.n52 VSUBS 0.041076f
C251 VP.n53 VSUBS 0.041076f
C252 VP.n54 VSUBS 0.041076f
C253 VP.n55 VSUBS 0.07502f
C254 VP.n56 VSUBS 0.068651f
C255 VP.n57 VSUBS 0.581132f
C256 VP.n58 VSUBS 0.046089f
C257 VP.n59 VSUBS 0.041076f
C258 VP.n60 VSUBS 0.041076f
C259 VP.n61 VSUBS 0.041076f
C260 VP.n62 VSUBS 0.054028f
C261 VP.n63 VSUBS 0.065393f
C262 VP.n64 VSUBS 0.076172f
C263 VP.n65 VSUBS 0.041076f
C264 VP.n66 VSUBS 0.041076f
C265 VP.n67 VSUBS 0.041076f
C266 VP.n68 VSUBS 0.076172f
C267 VP.n69 VSUBS 0.065393f
C268 VP.n70 VSUBS 0.054028f
C269 VP.n71 VSUBS 0.041076f
C270 VP.n72 VSUBS 0.041076f
C271 VP.n73 VSUBS 0.041076f
C272 VP.n74 VSUBS 0.046089f
C273 VP.n75 VSUBS 0.581132f
C274 VP.n76 VSUBS 0.068651f
C275 VP.n77 VSUBS 0.07502f
C276 VP.n78 VSUBS 0.041076f
C277 VP.n79 VSUBS 0.041076f
C278 VP.n80 VSUBS 0.041076f
C279 VP.n81 VSUBS 0.081845f
C280 VP.n82 VSUBS 0.05361f
C281 VP.n83 VSUBS 0.699259f
C282 VP.n84 VSUBS 0.062768f
C283 B.n0 VSUBS 0.006604f
C284 B.n1 VSUBS 0.006604f
C285 B.n2 VSUBS 0.010443f
C286 B.n3 VSUBS 0.010443f
C287 B.n4 VSUBS 0.010443f
C288 B.n5 VSUBS 0.010443f
C289 B.n6 VSUBS 0.010443f
C290 B.n7 VSUBS 0.010443f
C291 B.n8 VSUBS 0.010443f
C292 B.n9 VSUBS 0.010443f
C293 B.n10 VSUBS 0.010443f
C294 B.n11 VSUBS 0.010443f
C295 B.n12 VSUBS 0.010443f
C296 B.n13 VSUBS 0.010443f
C297 B.n14 VSUBS 0.010443f
C298 B.n15 VSUBS 0.010443f
C299 B.n16 VSUBS 0.010443f
C300 B.n17 VSUBS 0.010443f
C301 B.n18 VSUBS 0.010443f
C302 B.n19 VSUBS 0.010443f
C303 B.n20 VSUBS 0.010443f
C304 B.n21 VSUBS 0.010443f
C305 B.n22 VSUBS 0.010443f
C306 B.n23 VSUBS 0.010443f
C307 B.n24 VSUBS 0.010443f
C308 B.n25 VSUBS 0.010443f
C309 B.n26 VSUBS 0.010443f
C310 B.n27 VSUBS 0.010443f
C311 B.n28 VSUBS 0.010443f
C312 B.n29 VSUBS 0.024742f
C313 B.n30 VSUBS 0.010443f
C314 B.n31 VSUBS 0.010443f
C315 B.n32 VSUBS 0.010443f
C316 B.n33 VSUBS 0.010443f
C317 B.n34 VSUBS 0.010443f
C318 B.n35 VSUBS 0.010443f
C319 B.n36 VSUBS 0.010443f
C320 B.n37 VSUBS 0.010443f
C321 B.n38 VSUBS 0.010443f
C322 B.n39 VSUBS 0.010443f
C323 B.n40 VSUBS 0.010443f
C324 B.n41 VSUBS 0.010443f
C325 B.t2 VSUBS 0.27406f
C326 B.t1 VSUBS 0.301477f
C327 B.t0 VSUBS 0.990628f
C328 B.n42 VSUBS 0.172279f
C329 B.n43 VSUBS 0.103748f
C330 B.n44 VSUBS 0.010443f
C331 B.n45 VSUBS 0.010443f
C332 B.n46 VSUBS 0.010443f
C333 B.n47 VSUBS 0.010443f
C334 B.t8 VSUBS 0.274059f
C335 B.t7 VSUBS 0.301475f
C336 B.t6 VSUBS 0.990628f
C337 B.n48 VSUBS 0.172281f
C338 B.n49 VSUBS 0.103749f
C339 B.n50 VSUBS 0.024196f
C340 B.n51 VSUBS 0.010443f
C341 B.n52 VSUBS 0.010443f
C342 B.n53 VSUBS 0.010443f
C343 B.n54 VSUBS 0.010443f
C344 B.n55 VSUBS 0.010443f
C345 B.n56 VSUBS 0.010443f
C346 B.n57 VSUBS 0.010443f
C347 B.n58 VSUBS 0.010443f
C348 B.n59 VSUBS 0.010443f
C349 B.n60 VSUBS 0.010443f
C350 B.n61 VSUBS 0.010443f
C351 B.n62 VSUBS 0.010443f
C352 B.n63 VSUBS 0.023482f
C353 B.n64 VSUBS 0.010443f
C354 B.n65 VSUBS 0.010443f
C355 B.n66 VSUBS 0.010443f
C356 B.n67 VSUBS 0.010443f
C357 B.n68 VSUBS 0.010443f
C358 B.n69 VSUBS 0.010443f
C359 B.n70 VSUBS 0.010443f
C360 B.n71 VSUBS 0.010443f
C361 B.n72 VSUBS 0.010443f
C362 B.n73 VSUBS 0.010443f
C363 B.n74 VSUBS 0.010443f
C364 B.n75 VSUBS 0.010443f
C365 B.n76 VSUBS 0.010443f
C366 B.n77 VSUBS 0.010443f
C367 B.n78 VSUBS 0.010443f
C368 B.n79 VSUBS 0.010443f
C369 B.n80 VSUBS 0.010443f
C370 B.n81 VSUBS 0.010443f
C371 B.n82 VSUBS 0.010443f
C372 B.n83 VSUBS 0.010443f
C373 B.n84 VSUBS 0.010443f
C374 B.n85 VSUBS 0.010443f
C375 B.n86 VSUBS 0.010443f
C376 B.n87 VSUBS 0.010443f
C377 B.n88 VSUBS 0.010443f
C378 B.n89 VSUBS 0.010443f
C379 B.n90 VSUBS 0.010443f
C380 B.n91 VSUBS 0.010443f
C381 B.n92 VSUBS 0.010443f
C382 B.n93 VSUBS 0.010443f
C383 B.n94 VSUBS 0.010443f
C384 B.n95 VSUBS 0.010443f
C385 B.n96 VSUBS 0.010443f
C386 B.n97 VSUBS 0.010443f
C387 B.n98 VSUBS 0.010443f
C388 B.n99 VSUBS 0.010443f
C389 B.n100 VSUBS 0.010443f
C390 B.n101 VSUBS 0.010443f
C391 B.n102 VSUBS 0.010443f
C392 B.n103 VSUBS 0.010443f
C393 B.n104 VSUBS 0.010443f
C394 B.n105 VSUBS 0.010443f
C395 B.n106 VSUBS 0.010443f
C396 B.n107 VSUBS 0.010443f
C397 B.n108 VSUBS 0.010443f
C398 B.n109 VSUBS 0.010443f
C399 B.n110 VSUBS 0.010443f
C400 B.n111 VSUBS 0.010443f
C401 B.n112 VSUBS 0.010443f
C402 B.n113 VSUBS 0.010443f
C403 B.n114 VSUBS 0.010443f
C404 B.n115 VSUBS 0.010443f
C405 B.n116 VSUBS 0.010443f
C406 B.n117 VSUBS 0.023482f
C407 B.n118 VSUBS 0.010443f
C408 B.n119 VSUBS 0.010443f
C409 B.n120 VSUBS 0.010443f
C410 B.n121 VSUBS 0.010443f
C411 B.n122 VSUBS 0.010443f
C412 B.n123 VSUBS 0.010443f
C413 B.n124 VSUBS 0.010443f
C414 B.n125 VSUBS 0.010443f
C415 B.n126 VSUBS 0.010443f
C416 B.n127 VSUBS 0.010443f
C417 B.n128 VSUBS 0.010443f
C418 B.n129 VSUBS 0.010443f
C419 B.t4 VSUBS 0.274059f
C420 B.t5 VSUBS 0.301475f
C421 B.t3 VSUBS 0.990628f
C422 B.n130 VSUBS 0.172281f
C423 B.n131 VSUBS 0.103749f
C424 B.n132 VSUBS 0.024196f
C425 B.n133 VSUBS 0.010443f
C426 B.n134 VSUBS 0.010443f
C427 B.n135 VSUBS 0.010443f
C428 B.n136 VSUBS 0.010443f
C429 B.n137 VSUBS 0.010443f
C430 B.t10 VSUBS 0.27406f
C431 B.t11 VSUBS 0.301477f
C432 B.t9 VSUBS 0.990628f
C433 B.n138 VSUBS 0.172279f
C434 B.n139 VSUBS 0.103748f
C435 B.n140 VSUBS 0.010443f
C436 B.n141 VSUBS 0.010443f
C437 B.n142 VSUBS 0.010443f
C438 B.n143 VSUBS 0.010443f
C439 B.n144 VSUBS 0.010443f
C440 B.n145 VSUBS 0.010443f
C441 B.n146 VSUBS 0.010443f
C442 B.n147 VSUBS 0.010443f
C443 B.n148 VSUBS 0.010443f
C444 B.n149 VSUBS 0.010443f
C445 B.n150 VSUBS 0.010443f
C446 B.n151 VSUBS 0.024742f
C447 B.n152 VSUBS 0.010443f
C448 B.n153 VSUBS 0.010443f
C449 B.n154 VSUBS 0.010443f
C450 B.n155 VSUBS 0.010443f
C451 B.n156 VSUBS 0.010443f
C452 B.n157 VSUBS 0.010443f
C453 B.n158 VSUBS 0.010443f
C454 B.n159 VSUBS 0.010443f
C455 B.n160 VSUBS 0.010443f
C456 B.n161 VSUBS 0.010443f
C457 B.n162 VSUBS 0.010443f
C458 B.n163 VSUBS 0.010443f
C459 B.n164 VSUBS 0.010443f
C460 B.n165 VSUBS 0.010443f
C461 B.n166 VSUBS 0.010443f
C462 B.n167 VSUBS 0.010443f
C463 B.n168 VSUBS 0.010443f
C464 B.n169 VSUBS 0.010443f
C465 B.n170 VSUBS 0.010443f
C466 B.n171 VSUBS 0.010443f
C467 B.n172 VSUBS 0.010443f
C468 B.n173 VSUBS 0.010443f
C469 B.n174 VSUBS 0.010443f
C470 B.n175 VSUBS 0.010443f
C471 B.n176 VSUBS 0.010443f
C472 B.n177 VSUBS 0.010443f
C473 B.n178 VSUBS 0.010443f
C474 B.n179 VSUBS 0.010443f
C475 B.n180 VSUBS 0.010443f
C476 B.n181 VSUBS 0.010443f
C477 B.n182 VSUBS 0.010443f
C478 B.n183 VSUBS 0.010443f
C479 B.n184 VSUBS 0.010443f
C480 B.n185 VSUBS 0.010443f
C481 B.n186 VSUBS 0.010443f
C482 B.n187 VSUBS 0.010443f
C483 B.n188 VSUBS 0.010443f
C484 B.n189 VSUBS 0.010443f
C485 B.n190 VSUBS 0.010443f
C486 B.n191 VSUBS 0.010443f
C487 B.n192 VSUBS 0.010443f
C488 B.n193 VSUBS 0.010443f
C489 B.n194 VSUBS 0.010443f
C490 B.n195 VSUBS 0.010443f
C491 B.n196 VSUBS 0.010443f
C492 B.n197 VSUBS 0.010443f
C493 B.n198 VSUBS 0.010443f
C494 B.n199 VSUBS 0.010443f
C495 B.n200 VSUBS 0.010443f
C496 B.n201 VSUBS 0.010443f
C497 B.n202 VSUBS 0.010443f
C498 B.n203 VSUBS 0.010443f
C499 B.n204 VSUBS 0.010443f
C500 B.n205 VSUBS 0.010443f
C501 B.n206 VSUBS 0.010443f
C502 B.n207 VSUBS 0.010443f
C503 B.n208 VSUBS 0.010443f
C504 B.n209 VSUBS 0.010443f
C505 B.n210 VSUBS 0.010443f
C506 B.n211 VSUBS 0.010443f
C507 B.n212 VSUBS 0.010443f
C508 B.n213 VSUBS 0.010443f
C509 B.n214 VSUBS 0.010443f
C510 B.n215 VSUBS 0.010443f
C511 B.n216 VSUBS 0.010443f
C512 B.n217 VSUBS 0.010443f
C513 B.n218 VSUBS 0.010443f
C514 B.n219 VSUBS 0.010443f
C515 B.n220 VSUBS 0.010443f
C516 B.n221 VSUBS 0.010443f
C517 B.n222 VSUBS 0.010443f
C518 B.n223 VSUBS 0.010443f
C519 B.n224 VSUBS 0.010443f
C520 B.n225 VSUBS 0.010443f
C521 B.n226 VSUBS 0.010443f
C522 B.n227 VSUBS 0.010443f
C523 B.n228 VSUBS 0.010443f
C524 B.n229 VSUBS 0.010443f
C525 B.n230 VSUBS 0.010443f
C526 B.n231 VSUBS 0.010443f
C527 B.n232 VSUBS 0.010443f
C528 B.n233 VSUBS 0.010443f
C529 B.n234 VSUBS 0.010443f
C530 B.n235 VSUBS 0.010443f
C531 B.n236 VSUBS 0.010443f
C532 B.n237 VSUBS 0.010443f
C533 B.n238 VSUBS 0.010443f
C534 B.n239 VSUBS 0.010443f
C535 B.n240 VSUBS 0.010443f
C536 B.n241 VSUBS 0.010443f
C537 B.n242 VSUBS 0.010443f
C538 B.n243 VSUBS 0.010443f
C539 B.n244 VSUBS 0.010443f
C540 B.n245 VSUBS 0.010443f
C541 B.n246 VSUBS 0.010443f
C542 B.n247 VSUBS 0.010443f
C543 B.n248 VSUBS 0.010443f
C544 B.n249 VSUBS 0.010443f
C545 B.n250 VSUBS 0.010443f
C546 B.n251 VSUBS 0.010443f
C547 B.n252 VSUBS 0.010443f
C548 B.n253 VSUBS 0.010443f
C549 B.n254 VSUBS 0.010443f
C550 B.n255 VSUBS 0.010443f
C551 B.n256 VSUBS 0.023482f
C552 B.n257 VSUBS 0.023482f
C553 B.n258 VSUBS 0.024742f
C554 B.n259 VSUBS 0.010443f
C555 B.n260 VSUBS 0.010443f
C556 B.n261 VSUBS 0.010443f
C557 B.n262 VSUBS 0.010443f
C558 B.n263 VSUBS 0.010443f
C559 B.n264 VSUBS 0.010443f
C560 B.n265 VSUBS 0.010443f
C561 B.n266 VSUBS 0.010443f
C562 B.n267 VSUBS 0.010443f
C563 B.n268 VSUBS 0.010443f
C564 B.n269 VSUBS 0.010443f
C565 B.n270 VSUBS 0.010443f
C566 B.n271 VSUBS 0.010443f
C567 B.n272 VSUBS 0.010443f
C568 B.n273 VSUBS 0.010443f
C569 B.n274 VSUBS 0.010443f
C570 B.n275 VSUBS 0.010443f
C571 B.n276 VSUBS 0.010443f
C572 B.n277 VSUBS 0.010443f
C573 B.n278 VSUBS 0.010443f
C574 B.n279 VSUBS 0.010443f
C575 B.n280 VSUBS 0.010443f
C576 B.n281 VSUBS 0.010443f
C577 B.n282 VSUBS 0.010443f
C578 B.n283 VSUBS 0.010443f
C579 B.n284 VSUBS 0.010443f
C580 B.n285 VSUBS 0.010443f
C581 B.n286 VSUBS 0.010443f
C582 B.n287 VSUBS 0.010443f
C583 B.n288 VSUBS 0.010443f
C584 B.n289 VSUBS 0.010443f
C585 B.n290 VSUBS 0.010443f
C586 B.n291 VSUBS 0.010443f
C587 B.n292 VSUBS 0.010443f
C588 B.n293 VSUBS 0.010443f
C589 B.n294 VSUBS 0.007218f
C590 B.n295 VSUBS 0.024196f
C591 B.n296 VSUBS 0.008447f
C592 B.n297 VSUBS 0.010443f
C593 B.n298 VSUBS 0.010443f
C594 B.n299 VSUBS 0.010443f
C595 B.n300 VSUBS 0.010443f
C596 B.n301 VSUBS 0.010443f
C597 B.n302 VSUBS 0.010443f
C598 B.n303 VSUBS 0.010443f
C599 B.n304 VSUBS 0.010443f
C600 B.n305 VSUBS 0.010443f
C601 B.n306 VSUBS 0.010443f
C602 B.n307 VSUBS 0.010443f
C603 B.n308 VSUBS 0.008447f
C604 B.n309 VSUBS 0.010443f
C605 B.n310 VSUBS 0.010443f
C606 B.n311 VSUBS 0.007218f
C607 B.n312 VSUBS 0.010443f
C608 B.n313 VSUBS 0.010443f
C609 B.n314 VSUBS 0.010443f
C610 B.n315 VSUBS 0.010443f
C611 B.n316 VSUBS 0.010443f
C612 B.n317 VSUBS 0.010443f
C613 B.n318 VSUBS 0.010443f
C614 B.n319 VSUBS 0.010443f
C615 B.n320 VSUBS 0.010443f
C616 B.n321 VSUBS 0.010443f
C617 B.n322 VSUBS 0.010443f
C618 B.n323 VSUBS 0.010443f
C619 B.n324 VSUBS 0.010443f
C620 B.n325 VSUBS 0.010443f
C621 B.n326 VSUBS 0.010443f
C622 B.n327 VSUBS 0.010443f
C623 B.n328 VSUBS 0.010443f
C624 B.n329 VSUBS 0.010443f
C625 B.n330 VSUBS 0.010443f
C626 B.n331 VSUBS 0.010443f
C627 B.n332 VSUBS 0.010443f
C628 B.n333 VSUBS 0.010443f
C629 B.n334 VSUBS 0.010443f
C630 B.n335 VSUBS 0.010443f
C631 B.n336 VSUBS 0.010443f
C632 B.n337 VSUBS 0.010443f
C633 B.n338 VSUBS 0.010443f
C634 B.n339 VSUBS 0.010443f
C635 B.n340 VSUBS 0.010443f
C636 B.n341 VSUBS 0.010443f
C637 B.n342 VSUBS 0.010443f
C638 B.n343 VSUBS 0.010443f
C639 B.n344 VSUBS 0.010443f
C640 B.n345 VSUBS 0.010443f
C641 B.n346 VSUBS 0.024742f
C642 B.n347 VSUBS 0.024742f
C643 B.n348 VSUBS 0.023482f
C644 B.n349 VSUBS 0.010443f
C645 B.n350 VSUBS 0.010443f
C646 B.n351 VSUBS 0.010443f
C647 B.n352 VSUBS 0.010443f
C648 B.n353 VSUBS 0.010443f
C649 B.n354 VSUBS 0.010443f
C650 B.n355 VSUBS 0.010443f
C651 B.n356 VSUBS 0.010443f
C652 B.n357 VSUBS 0.010443f
C653 B.n358 VSUBS 0.010443f
C654 B.n359 VSUBS 0.010443f
C655 B.n360 VSUBS 0.010443f
C656 B.n361 VSUBS 0.010443f
C657 B.n362 VSUBS 0.010443f
C658 B.n363 VSUBS 0.010443f
C659 B.n364 VSUBS 0.010443f
C660 B.n365 VSUBS 0.010443f
C661 B.n366 VSUBS 0.010443f
C662 B.n367 VSUBS 0.010443f
C663 B.n368 VSUBS 0.010443f
C664 B.n369 VSUBS 0.010443f
C665 B.n370 VSUBS 0.010443f
C666 B.n371 VSUBS 0.010443f
C667 B.n372 VSUBS 0.010443f
C668 B.n373 VSUBS 0.010443f
C669 B.n374 VSUBS 0.010443f
C670 B.n375 VSUBS 0.010443f
C671 B.n376 VSUBS 0.010443f
C672 B.n377 VSUBS 0.010443f
C673 B.n378 VSUBS 0.010443f
C674 B.n379 VSUBS 0.010443f
C675 B.n380 VSUBS 0.010443f
C676 B.n381 VSUBS 0.010443f
C677 B.n382 VSUBS 0.010443f
C678 B.n383 VSUBS 0.010443f
C679 B.n384 VSUBS 0.010443f
C680 B.n385 VSUBS 0.010443f
C681 B.n386 VSUBS 0.010443f
C682 B.n387 VSUBS 0.010443f
C683 B.n388 VSUBS 0.010443f
C684 B.n389 VSUBS 0.010443f
C685 B.n390 VSUBS 0.010443f
C686 B.n391 VSUBS 0.010443f
C687 B.n392 VSUBS 0.010443f
C688 B.n393 VSUBS 0.010443f
C689 B.n394 VSUBS 0.010443f
C690 B.n395 VSUBS 0.010443f
C691 B.n396 VSUBS 0.010443f
C692 B.n397 VSUBS 0.010443f
C693 B.n398 VSUBS 0.010443f
C694 B.n399 VSUBS 0.010443f
C695 B.n400 VSUBS 0.010443f
C696 B.n401 VSUBS 0.010443f
C697 B.n402 VSUBS 0.010443f
C698 B.n403 VSUBS 0.010443f
C699 B.n404 VSUBS 0.010443f
C700 B.n405 VSUBS 0.010443f
C701 B.n406 VSUBS 0.010443f
C702 B.n407 VSUBS 0.010443f
C703 B.n408 VSUBS 0.010443f
C704 B.n409 VSUBS 0.010443f
C705 B.n410 VSUBS 0.010443f
C706 B.n411 VSUBS 0.010443f
C707 B.n412 VSUBS 0.010443f
C708 B.n413 VSUBS 0.010443f
C709 B.n414 VSUBS 0.010443f
C710 B.n415 VSUBS 0.010443f
C711 B.n416 VSUBS 0.010443f
C712 B.n417 VSUBS 0.010443f
C713 B.n418 VSUBS 0.010443f
C714 B.n419 VSUBS 0.010443f
C715 B.n420 VSUBS 0.010443f
C716 B.n421 VSUBS 0.010443f
C717 B.n422 VSUBS 0.010443f
C718 B.n423 VSUBS 0.010443f
C719 B.n424 VSUBS 0.010443f
C720 B.n425 VSUBS 0.010443f
C721 B.n426 VSUBS 0.010443f
C722 B.n427 VSUBS 0.010443f
C723 B.n428 VSUBS 0.010443f
C724 B.n429 VSUBS 0.010443f
C725 B.n430 VSUBS 0.010443f
C726 B.n431 VSUBS 0.010443f
C727 B.n432 VSUBS 0.010443f
C728 B.n433 VSUBS 0.010443f
C729 B.n434 VSUBS 0.010443f
C730 B.n435 VSUBS 0.010443f
C731 B.n436 VSUBS 0.010443f
C732 B.n437 VSUBS 0.010443f
C733 B.n438 VSUBS 0.010443f
C734 B.n439 VSUBS 0.010443f
C735 B.n440 VSUBS 0.010443f
C736 B.n441 VSUBS 0.010443f
C737 B.n442 VSUBS 0.010443f
C738 B.n443 VSUBS 0.010443f
C739 B.n444 VSUBS 0.010443f
C740 B.n445 VSUBS 0.010443f
C741 B.n446 VSUBS 0.010443f
C742 B.n447 VSUBS 0.010443f
C743 B.n448 VSUBS 0.010443f
C744 B.n449 VSUBS 0.010443f
C745 B.n450 VSUBS 0.010443f
C746 B.n451 VSUBS 0.010443f
C747 B.n452 VSUBS 0.010443f
C748 B.n453 VSUBS 0.010443f
C749 B.n454 VSUBS 0.010443f
C750 B.n455 VSUBS 0.010443f
C751 B.n456 VSUBS 0.010443f
C752 B.n457 VSUBS 0.010443f
C753 B.n458 VSUBS 0.010443f
C754 B.n459 VSUBS 0.010443f
C755 B.n460 VSUBS 0.010443f
C756 B.n461 VSUBS 0.010443f
C757 B.n462 VSUBS 0.010443f
C758 B.n463 VSUBS 0.010443f
C759 B.n464 VSUBS 0.010443f
C760 B.n465 VSUBS 0.010443f
C761 B.n466 VSUBS 0.010443f
C762 B.n467 VSUBS 0.010443f
C763 B.n468 VSUBS 0.010443f
C764 B.n469 VSUBS 0.010443f
C765 B.n470 VSUBS 0.010443f
C766 B.n471 VSUBS 0.010443f
C767 B.n472 VSUBS 0.010443f
C768 B.n473 VSUBS 0.010443f
C769 B.n474 VSUBS 0.010443f
C770 B.n475 VSUBS 0.010443f
C771 B.n476 VSUBS 0.010443f
C772 B.n477 VSUBS 0.010443f
C773 B.n478 VSUBS 0.010443f
C774 B.n479 VSUBS 0.010443f
C775 B.n480 VSUBS 0.010443f
C776 B.n481 VSUBS 0.010443f
C777 B.n482 VSUBS 0.010443f
C778 B.n483 VSUBS 0.010443f
C779 B.n484 VSUBS 0.010443f
C780 B.n485 VSUBS 0.010443f
C781 B.n486 VSUBS 0.010443f
C782 B.n487 VSUBS 0.010443f
C783 B.n488 VSUBS 0.010443f
C784 B.n489 VSUBS 0.010443f
C785 B.n490 VSUBS 0.010443f
C786 B.n491 VSUBS 0.010443f
C787 B.n492 VSUBS 0.010443f
C788 B.n493 VSUBS 0.010443f
C789 B.n494 VSUBS 0.010443f
C790 B.n495 VSUBS 0.010443f
C791 B.n496 VSUBS 0.010443f
C792 B.n497 VSUBS 0.010443f
C793 B.n498 VSUBS 0.010443f
C794 B.n499 VSUBS 0.010443f
C795 B.n500 VSUBS 0.010443f
C796 B.n501 VSUBS 0.010443f
C797 B.n502 VSUBS 0.010443f
C798 B.n503 VSUBS 0.010443f
C799 B.n504 VSUBS 0.010443f
C800 B.n505 VSUBS 0.010443f
C801 B.n506 VSUBS 0.010443f
C802 B.n507 VSUBS 0.010443f
C803 B.n508 VSUBS 0.010443f
C804 B.n509 VSUBS 0.010443f
C805 B.n510 VSUBS 0.024742f
C806 B.n511 VSUBS 0.023482f
C807 B.n512 VSUBS 0.024742f
C808 B.n513 VSUBS 0.010443f
C809 B.n514 VSUBS 0.010443f
C810 B.n515 VSUBS 0.010443f
C811 B.n516 VSUBS 0.010443f
C812 B.n517 VSUBS 0.010443f
C813 B.n518 VSUBS 0.010443f
C814 B.n519 VSUBS 0.010443f
C815 B.n520 VSUBS 0.010443f
C816 B.n521 VSUBS 0.010443f
C817 B.n522 VSUBS 0.010443f
C818 B.n523 VSUBS 0.010443f
C819 B.n524 VSUBS 0.010443f
C820 B.n525 VSUBS 0.010443f
C821 B.n526 VSUBS 0.010443f
C822 B.n527 VSUBS 0.010443f
C823 B.n528 VSUBS 0.010443f
C824 B.n529 VSUBS 0.010443f
C825 B.n530 VSUBS 0.010443f
C826 B.n531 VSUBS 0.010443f
C827 B.n532 VSUBS 0.010443f
C828 B.n533 VSUBS 0.010443f
C829 B.n534 VSUBS 0.010443f
C830 B.n535 VSUBS 0.010443f
C831 B.n536 VSUBS 0.010443f
C832 B.n537 VSUBS 0.010443f
C833 B.n538 VSUBS 0.010443f
C834 B.n539 VSUBS 0.010443f
C835 B.n540 VSUBS 0.010443f
C836 B.n541 VSUBS 0.010443f
C837 B.n542 VSUBS 0.010443f
C838 B.n543 VSUBS 0.010443f
C839 B.n544 VSUBS 0.010443f
C840 B.n545 VSUBS 0.010443f
C841 B.n546 VSUBS 0.010443f
C842 B.n547 VSUBS 0.007218f
C843 B.n548 VSUBS 0.010443f
C844 B.n549 VSUBS 0.010443f
C845 B.n550 VSUBS 0.008447f
C846 B.n551 VSUBS 0.010443f
C847 B.n552 VSUBS 0.010443f
C848 B.n553 VSUBS 0.010443f
C849 B.n554 VSUBS 0.010443f
C850 B.n555 VSUBS 0.010443f
C851 B.n556 VSUBS 0.010443f
C852 B.n557 VSUBS 0.010443f
C853 B.n558 VSUBS 0.010443f
C854 B.n559 VSUBS 0.010443f
C855 B.n560 VSUBS 0.010443f
C856 B.n561 VSUBS 0.010443f
C857 B.n562 VSUBS 0.008447f
C858 B.n563 VSUBS 0.024196f
C859 B.n564 VSUBS 0.007218f
C860 B.n565 VSUBS 0.010443f
C861 B.n566 VSUBS 0.010443f
C862 B.n567 VSUBS 0.010443f
C863 B.n568 VSUBS 0.010443f
C864 B.n569 VSUBS 0.010443f
C865 B.n570 VSUBS 0.010443f
C866 B.n571 VSUBS 0.010443f
C867 B.n572 VSUBS 0.010443f
C868 B.n573 VSUBS 0.010443f
C869 B.n574 VSUBS 0.010443f
C870 B.n575 VSUBS 0.010443f
C871 B.n576 VSUBS 0.010443f
C872 B.n577 VSUBS 0.010443f
C873 B.n578 VSUBS 0.010443f
C874 B.n579 VSUBS 0.010443f
C875 B.n580 VSUBS 0.010443f
C876 B.n581 VSUBS 0.010443f
C877 B.n582 VSUBS 0.010443f
C878 B.n583 VSUBS 0.010443f
C879 B.n584 VSUBS 0.010443f
C880 B.n585 VSUBS 0.010443f
C881 B.n586 VSUBS 0.010443f
C882 B.n587 VSUBS 0.010443f
C883 B.n588 VSUBS 0.010443f
C884 B.n589 VSUBS 0.010443f
C885 B.n590 VSUBS 0.010443f
C886 B.n591 VSUBS 0.010443f
C887 B.n592 VSUBS 0.010443f
C888 B.n593 VSUBS 0.010443f
C889 B.n594 VSUBS 0.010443f
C890 B.n595 VSUBS 0.010443f
C891 B.n596 VSUBS 0.010443f
C892 B.n597 VSUBS 0.010443f
C893 B.n598 VSUBS 0.010443f
C894 B.n599 VSUBS 0.010443f
C895 B.n600 VSUBS 0.024742f
C896 B.n601 VSUBS 0.023482f
C897 B.n602 VSUBS 0.023482f
C898 B.n603 VSUBS 0.010443f
C899 B.n604 VSUBS 0.010443f
C900 B.n605 VSUBS 0.010443f
C901 B.n606 VSUBS 0.010443f
C902 B.n607 VSUBS 0.010443f
C903 B.n608 VSUBS 0.010443f
C904 B.n609 VSUBS 0.010443f
C905 B.n610 VSUBS 0.010443f
C906 B.n611 VSUBS 0.010443f
C907 B.n612 VSUBS 0.010443f
C908 B.n613 VSUBS 0.010443f
C909 B.n614 VSUBS 0.010443f
C910 B.n615 VSUBS 0.010443f
C911 B.n616 VSUBS 0.010443f
C912 B.n617 VSUBS 0.010443f
C913 B.n618 VSUBS 0.010443f
C914 B.n619 VSUBS 0.010443f
C915 B.n620 VSUBS 0.010443f
C916 B.n621 VSUBS 0.010443f
C917 B.n622 VSUBS 0.010443f
C918 B.n623 VSUBS 0.010443f
C919 B.n624 VSUBS 0.010443f
C920 B.n625 VSUBS 0.010443f
C921 B.n626 VSUBS 0.010443f
C922 B.n627 VSUBS 0.010443f
C923 B.n628 VSUBS 0.010443f
C924 B.n629 VSUBS 0.010443f
C925 B.n630 VSUBS 0.010443f
C926 B.n631 VSUBS 0.010443f
C927 B.n632 VSUBS 0.010443f
C928 B.n633 VSUBS 0.010443f
C929 B.n634 VSUBS 0.010443f
C930 B.n635 VSUBS 0.010443f
C931 B.n636 VSUBS 0.010443f
C932 B.n637 VSUBS 0.010443f
C933 B.n638 VSUBS 0.010443f
C934 B.n639 VSUBS 0.010443f
C935 B.n640 VSUBS 0.010443f
C936 B.n641 VSUBS 0.010443f
C937 B.n642 VSUBS 0.010443f
C938 B.n643 VSUBS 0.010443f
C939 B.n644 VSUBS 0.010443f
C940 B.n645 VSUBS 0.010443f
C941 B.n646 VSUBS 0.010443f
C942 B.n647 VSUBS 0.010443f
C943 B.n648 VSUBS 0.010443f
C944 B.n649 VSUBS 0.010443f
C945 B.n650 VSUBS 0.010443f
C946 B.n651 VSUBS 0.010443f
C947 B.n652 VSUBS 0.010443f
C948 B.n653 VSUBS 0.010443f
C949 B.n654 VSUBS 0.010443f
C950 B.n655 VSUBS 0.010443f
C951 B.n656 VSUBS 0.010443f
C952 B.n657 VSUBS 0.010443f
C953 B.n658 VSUBS 0.010443f
C954 B.n659 VSUBS 0.010443f
C955 B.n660 VSUBS 0.010443f
C956 B.n661 VSUBS 0.010443f
C957 B.n662 VSUBS 0.010443f
C958 B.n663 VSUBS 0.010443f
C959 B.n664 VSUBS 0.010443f
C960 B.n665 VSUBS 0.010443f
C961 B.n666 VSUBS 0.010443f
C962 B.n667 VSUBS 0.010443f
C963 B.n668 VSUBS 0.010443f
C964 B.n669 VSUBS 0.010443f
C965 B.n670 VSUBS 0.010443f
C966 B.n671 VSUBS 0.010443f
C967 B.n672 VSUBS 0.010443f
C968 B.n673 VSUBS 0.010443f
C969 B.n674 VSUBS 0.010443f
C970 B.n675 VSUBS 0.010443f
C971 B.n676 VSUBS 0.010443f
C972 B.n677 VSUBS 0.010443f
C973 B.n678 VSUBS 0.010443f
C974 B.n679 VSUBS 0.010443f
C975 B.n680 VSUBS 0.010443f
C976 B.n681 VSUBS 0.010443f
C977 B.n682 VSUBS 0.010443f
C978 B.n683 VSUBS 0.023647f
.ends

