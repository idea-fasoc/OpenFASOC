* NGSPICE file created from diff_pair_sample_1065.ext - technology: sky130A

.subckt diff_pair_sample_1065 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t5 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X1 VDD2.t4 VN.t1 VTAIL.t14 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=6.3999 ps=33.6 w=16.41 l=2.06
X2 VTAIL.t0 VP.t0 VDD1.t7 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=2.70765 ps=16.74 w=16.41 l=2.06
X3 B.t11 B.t9 B.t10 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=2.06
X4 VDD1.t6 VP.t1 VTAIL.t4 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=6.3999 ps=33.6 w=16.41 l=2.06
X5 VDD1.t5 VP.t2 VTAIL.t1 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X6 VTAIL.t13 VN.t2 VDD2.t1 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=2.70765 ps=16.74 w=16.41 l=2.06
X7 B.t8 B.t6 B.t7 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=2.06
X8 VTAIL.t12 VN.t3 VDD2.t0 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=2.70765 ps=16.74 w=16.41 l=2.06
X9 VDD2.t3 VN.t4 VTAIL.t11 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=6.3999 ps=33.6 w=16.41 l=2.06
X10 VTAIL.t5 VP.t3 VDD1.t4 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X11 B.t5 B.t3 B.t4 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=2.06
X12 VDD2.t2 VN.t5 VTAIL.t10 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X13 VTAIL.t9 VN.t6 VDD2.t7 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X14 VDD1.t3 VP.t4 VTAIL.t3 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X15 B.t2 B.t0 B.t1 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=0 ps=0 w=16.41 l=2.06
X16 VTAIL.t2 VP.t5 VDD1.t2 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
X17 VTAIL.t6 VP.t6 VDD1.t1 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=6.3999 pd=33.6 as=2.70765 ps=16.74 w=16.41 l=2.06
X18 VDD1.t0 VP.t7 VTAIL.t7 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=6.3999 ps=33.6 w=16.41 l=2.06
X19 VDD2.t6 VN.t7 VTAIL.t8 w_n3360_n4250# sky130_fd_pr__pfet_01v8 ad=2.70765 pd=16.74 as=2.70765 ps=16.74 w=16.41 l=2.06
R0 VN.n5 VN.t3 225.405
R1 VN.n28 VN.t4 225.405
R2 VN.n6 VN.t7 191.982
R3 VN.n13 VN.t6 191.982
R4 VN.n21 VN.t1 191.982
R5 VN.n29 VN.t0 191.982
R6 VN.n36 VN.t5 191.982
R7 VN.n44 VN.t2 191.982
R8 VN.n43 VN.n23 161.3
R9 VN.n42 VN.n41 161.3
R10 VN.n40 VN.n24 161.3
R11 VN.n39 VN.n38 161.3
R12 VN.n37 VN.n25 161.3
R13 VN.n35 VN.n34 161.3
R14 VN.n33 VN.n26 161.3
R15 VN.n32 VN.n31 161.3
R16 VN.n30 VN.n27 161.3
R17 VN.n20 VN.n0 161.3
R18 VN.n19 VN.n18 161.3
R19 VN.n17 VN.n1 161.3
R20 VN.n16 VN.n15 161.3
R21 VN.n14 VN.n2 161.3
R22 VN.n12 VN.n11 161.3
R23 VN.n10 VN.n3 161.3
R24 VN.n9 VN.n8 161.3
R25 VN.n7 VN.n4 161.3
R26 VN.n22 VN.n21 94.3636
R27 VN.n45 VN.n44 94.3636
R28 VN.n8 VN.n3 56.5193
R29 VN.n31 VN.n26 56.5193
R30 VN.n19 VN.n1 54.0911
R31 VN.n42 VN.n24 54.0911
R32 VN VN.n45 51.9754
R33 VN.n6 VN.n5 48.7053
R34 VN.n29 VN.n28 48.7053
R35 VN.n15 VN.n1 26.8957
R36 VN.n38 VN.n24 26.8957
R37 VN.n8 VN.n7 24.4675
R38 VN.n12 VN.n3 24.4675
R39 VN.n15 VN.n14 24.4675
R40 VN.n20 VN.n19 24.4675
R41 VN.n31 VN.n30 24.4675
R42 VN.n38 VN.n37 24.4675
R43 VN.n35 VN.n26 24.4675
R44 VN.n43 VN.n42 24.4675
R45 VN.n7 VN.n6 21.7761
R46 VN.n13 VN.n12 21.7761
R47 VN.n30 VN.n29 21.7761
R48 VN.n36 VN.n35 21.7761
R49 VN.n21 VN.n20 16.3934
R50 VN.n44 VN.n43 16.3934
R51 VN.n28 VN.n27 9.30567
R52 VN.n5 VN.n4 9.30567
R53 VN.n14 VN.n13 2.69187
R54 VN.n37 VN.n36 2.69187
R55 VN.n45 VN.n23 0.278367
R56 VN.n22 VN.n0 0.278367
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153454
R74 VDD2.n2 VDD2.n1 69.9842
R75 VDD2.n2 VDD2.n0 69.9842
R76 VDD2 VDD2.n5 69.9814
R77 VDD2.n4 VDD2.n3 69.0097
R78 VDD2.n4 VDD2.n2 47.1334
R79 VDD2.n5 VDD2.t5 1.9813
R80 VDD2.n5 VDD2.t3 1.9813
R81 VDD2.n3 VDD2.t1 1.9813
R82 VDD2.n3 VDD2.t2 1.9813
R83 VDD2.n1 VDD2.t7 1.9813
R84 VDD2.n1 VDD2.t4 1.9813
R85 VDD2.n0 VDD2.t0 1.9813
R86 VDD2.n0 VDD2.t6 1.9813
R87 VDD2 VDD2.n4 1.08886
R88 VTAIL.n11 VTAIL.t0 54.3117
R89 VTAIL.n10 VTAIL.t11 54.3117
R90 VTAIL.n7 VTAIL.t13 54.3117
R91 VTAIL.n15 VTAIL.t14 54.3114
R92 VTAIL.n2 VTAIL.t12 54.3114
R93 VTAIL.n3 VTAIL.t4 54.3114
R94 VTAIL.n6 VTAIL.t6 54.3114
R95 VTAIL.n14 VTAIL.t7 54.3114
R96 VTAIL.n13 VTAIL.n12 52.3309
R97 VTAIL.n9 VTAIL.n8 52.3309
R98 VTAIL.n1 VTAIL.n0 52.3306
R99 VTAIL.n5 VTAIL.n4 52.3306
R100 VTAIL.n15 VTAIL.n14 28.5738
R101 VTAIL.n7 VTAIL.n6 28.5738
R102 VTAIL.n9 VTAIL.n7 2.06084
R103 VTAIL.n10 VTAIL.n9 2.06084
R104 VTAIL.n13 VTAIL.n11 2.06084
R105 VTAIL.n14 VTAIL.n13 2.06084
R106 VTAIL.n6 VTAIL.n5 2.06084
R107 VTAIL.n5 VTAIL.n3 2.06084
R108 VTAIL.n2 VTAIL.n1 2.06084
R109 VTAIL VTAIL.n15 2.00266
R110 VTAIL.n0 VTAIL.t8 1.9813
R111 VTAIL.n0 VTAIL.t9 1.9813
R112 VTAIL.n4 VTAIL.t1 1.9813
R113 VTAIL.n4 VTAIL.t2 1.9813
R114 VTAIL.n12 VTAIL.t3 1.9813
R115 VTAIL.n12 VTAIL.t5 1.9813
R116 VTAIL.n8 VTAIL.t10 1.9813
R117 VTAIL.n8 VTAIL.t15 1.9813
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 VP.n13 VP.t0 225.405
R122 VP.n7 VP.t6 191.982
R123 VP.n40 VP.t2 191.982
R124 VP.n47 VP.t5 191.982
R125 VP.n55 VP.t1 191.982
R126 VP.n29 VP.t7 191.982
R127 VP.n21 VP.t3 191.982
R128 VP.n14 VP.t4 191.982
R129 VP.n15 VP.n12 161.3
R130 VP.n17 VP.n16 161.3
R131 VP.n18 VP.n11 161.3
R132 VP.n20 VP.n19 161.3
R133 VP.n22 VP.n10 161.3
R134 VP.n24 VP.n23 161.3
R135 VP.n25 VP.n9 161.3
R136 VP.n27 VP.n26 161.3
R137 VP.n28 VP.n8 161.3
R138 VP.n54 VP.n0 161.3
R139 VP.n53 VP.n52 161.3
R140 VP.n51 VP.n1 161.3
R141 VP.n50 VP.n49 161.3
R142 VP.n48 VP.n2 161.3
R143 VP.n46 VP.n45 161.3
R144 VP.n44 VP.n3 161.3
R145 VP.n43 VP.n42 161.3
R146 VP.n41 VP.n4 161.3
R147 VP.n39 VP.n38 161.3
R148 VP.n37 VP.n5 161.3
R149 VP.n36 VP.n35 161.3
R150 VP.n34 VP.n6 161.3
R151 VP.n33 VP.n32 161.3
R152 VP.n31 VP.n7 94.3636
R153 VP.n56 VP.n55 94.3636
R154 VP.n30 VP.n29 94.3636
R155 VP.n42 VP.n3 56.5193
R156 VP.n16 VP.n11 56.5193
R157 VP.n35 VP.n34 54.0911
R158 VP.n53 VP.n1 54.0911
R159 VP.n27 VP.n9 54.0911
R160 VP.n31 VP.n30 51.6966
R161 VP.n14 VP.n13 48.7053
R162 VP.n35 VP.n5 26.8957
R163 VP.n49 VP.n1 26.8957
R164 VP.n23 VP.n9 26.8957
R165 VP.n34 VP.n33 24.4675
R166 VP.n39 VP.n5 24.4675
R167 VP.n42 VP.n41 24.4675
R168 VP.n46 VP.n3 24.4675
R169 VP.n49 VP.n48 24.4675
R170 VP.n54 VP.n53 24.4675
R171 VP.n28 VP.n27 24.4675
R172 VP.n20 VP.n11 24.4675
R173 VP.n23 VP.n22 24.4675
R174 VP.n16 VP.n15 24.4675
R175 VP.n41 VP.n40 21.7761
R176 VP.n47 VP.n46 21.7761
R177 VP.n21 VP.n20 21.7761
R178 VP.n15 VP.n14 21.7761
R179 VP.n33 VP.n7 16.3934
R180 VP.n55 VP.n54 16.3934
R181 VP.n29 VP.n28 16.3934
R182 VP.n13 VP.n12 9.30567
R183 VP.n40 VP.n39 2.69187
R184 VP.n48 VP.n47 2.69187
R185 VP.n22 VP.n21 2.69187
R186 VP.n30 VP.n8 0.278367
R187 VP.n32 VP.n31 0.278367
R188 VP.n56 VP.n0 0.278367
R189 VP.n17 VP.n12 0.189894
R190 VP.n18 VP.n17 0.189894
R191 VP.n19 VP.n18 0.189894
R192 VP.n19 VP.n10 0.189894
R193 VP.n24 VP.n10 0.189894
R194 VP.n25 VP.n24 0.189894
R195 VP.n26 VP.n25 0.189894
R196 VP.n26 VP.n8 0.189894
R197 VP.n32 VP.n6 0.189894
R198 VP.n36 VP.n6 0.189894
R199 VP.n37 VP.n36 0.189894
R200 VP.n38 VP.n37 0.189894
R201 VP.n38 VP.n4 0.189894
R202 VP.n43 VP.n4 0.189894
R203 VP.n44 VP.n43 0.189894
R204 VP.n45 VP.n44 0.189894
R205 VP.n45 VP.n2 0.189894
R206 VP.n50 VP.n2 0.189894
R207 VP.n51 VP.n50 0.189894
R208 VP.n52 VP.n51 0.189894
R209 VP.n52 VP.n0 0.189894
R210 VP VP.n56 0.153454
R211 VDD1 VDD1.n0 70.098
R212 VDD1.n3 VDD1.n2 69.9842
R213 VDD1.n3 VDD1.n1 69.9842
R214 VDD1.n5 VDD1.n4 69.0095
R215 VDD1.n5 VDD1.n3 47.7164
R216 VDD1.n4 VDD1.t4 1.9813
R217 VDD1.n4 VDD1.t0 1.9813
R218 VDD1.n0 VDD1.t7 1.9813
R219 VDD1.n0 VDD1.t3 1.9813
R220 VDD1.n2 VDD1.t2 1.9813
R221 VDD1.n2 VDD1.t6 1.9813
R222 VDD1.n1 VDD1.t1 1.9813
R223 VDD1.n1 VDD1.t5 1.9813
R224 VDD1 VDD1.n5 0.972483
R225 B.n590 B.n589 585
R226 B.n591 B.n86 585
R227 B.n593 B.n592 585
R228 B.n594 B.n85 585
R229 B.n596 B.n595 585
R230 B.n597 B.n84 585
R231 B.n599 B.n598 585
R232 B.n600 B.n83 585
R233 B.n602 B.n601 585
R234 B.n603 B.n82 585
R235 B.n605 B.n604 585
R236 B.n606 B.n81 585
R237 B.n608 B.n607 585
R238 B.n609 B.n80 585
R239 B.n611 B.n610 585
R240 B.n612 B.n79 585
R241 B.n614 B.n613 585
R242 B.n615 B.n78 585
R243 B.n617 B.n616 585
R244 B.n618 B.n77 585
R245 B.n620 B.n619 585
R246 B.n621 B.n76 585
R247 B.n623 B.n622 585
R248 B.n624 B.n75 585
R249 B.n626 B.n625 585
R250 B.n627 B.n74 585
R251 B.n629 B.n628 585
R252 B.n630 B.n73 585
R253 B.n632 B.n631 585
R254 B.n633 B.n72 585
R255 B.n635 B.n634 585
R256 B.n636 B.n71 585
R257 B.n638 B.n637 585
R258 B.n639 B.n70 585
R259 B.n641 B.n640 585
R260 B.n642 B.n69 585
R261 B.n644 B.n643 585
R262 B.n645 B.n68 585
R263 B.n647 B.n646 585
R264 B.n648 B.n67 585
R265 B.n650 B.n649 585
R266 B.n651 B.n66 585
R267 B.n653 B.n652 585
R268 B.n654 B.n65 585
R269 B.n656 B.n655 585
R270 B.n657 B.n64 585
R271 B.n659 B.n658 585
R272 B.n660 B.n63 585
R273 B.n662 B.n661 585
R274 B.n663 B.n62 585
R275 B.n665 B.n664 585
R276 B.n666 B.n61 585
R277 B.n668 B.n667 585
R278 B.n669 B.n60 585
R279 B.n671 B.n670 585
R280 B.n673 B.n57 585
R281 B.n675 B.n674 585
R282 B.n676 B.n56 585
R283 B.n678 B.n677 585
R284 B.n679 B.n55 585
R285 B.n681 B.n680 585
R286 B.n682 B.n54 585
R287 B.n684 B.n683 585
R288 B.n685 B.n51 585
R289 B.n688 B.n687 585
R290 B.n689 B.n50 585
R291 B.n691 B.n690 585
R292 B.n692 B.n49 585
R293 B.n694 B.n693 585
R294 B.n695 B.n48 585
R295 B.n697 B.n696 585
R296 B.n698 B.n47 585
R297 B.n700 B.n699 585
R298 B.n701 B.n46 585
R299 B.n703 B.n702 585
R300 B.n704 B.n45 585
R301 B.n706 B.n705 585
R302 B.n707 B.n44 585
R303 B.n709 B.n708 585
R304 B.n710 B.n43 585
R305 B.n712 B.n711 585
R306 B.n713 B.n42 585
R307 B.n715 B.n714 585
R308 B.n716 B.n41 585
R309 B.n718 B.n717 585
R310 B.n719 B.n40 585
R311 B.n721 B.n720 585
R312 B.n722 B.n39 585
R313 B.n724 B.n723 585
R314 B.n725 B.n38 585
R315 B.n727 B.n726 585
R316 B.n728 B.n37 585
R317 B.n730 B.n729 585
R318 B.n731 B.n36 585
R319 B.n733 B.n732 585
R320 B.n734 B.n35 585
R321 B.n736 B.n735 585
R322 B.n737 B.n34 585
R323 B.n739 B.n738 585
R324 B.n740 B.n33 585
R325 B.n742 B.n741 585
R326 B.n743 B.n32 585
R327 B.n745 B.n744 585
R328 B.n746 B.n31 585
R329 B.n748 B.n747 585
R330 B.n749 B.n30 585
R331 B.n751 B.n750 585
R332 B.n752 B.n29 585
R333 B.n754 B.n753 585
R334 B.n755 B.n28 585
R335 B.n757 B.n756 585
R336 B.n758 B.n27 585
R337 B.n760 B.n759 585
R338 B.n761 B.n26 585
R339 B.n763 B.n762 585
R340 B.n764 B.n25 585
R341 B.n766 B.n765 585
R342 B.n767 B.n24 585
R343 B.n769 B.n768 585
R344 B.n588 B.n87 585
R345 B.n587 B.n586 585
R346 B.n585 B.n88 585
R347 B.n584 B.n583 585
R348 B.n582 B.n89 585
R349 B.n581 B.n580 585
R350 B.n579 B.n90 585
R351 B.n578 B.n577 585
R352 B.n576 B.n91 585
R353 B.n575 B.n574 585
R354 B.n573 B.n92 585
R355 B.n572 B.n571 585
R356 B.n570 B.n93 585
R357 B.n569 B.n568 585
R358 B.n567 B.n94 585
R359 B.n566 B.n565 585
R360 B.n564 B.n95 585
R361 B.n563 B.n562 585
R362 B.n561 B.n96 585
R363 B.n560 B.n559 585
R364 B.n558 B.n97 585
R365 B.n557 B.n556 585
R366 B.n555 B.n98 585
R367 B.n554 B.n553 585
R368 B.n552 B.n99 585
R369 B.n551 B.n550 585
R370 B.n549 B.n100 585
R371 B.n548 B.n547 585
R372 B.n546 B.n101 585
R373 B.n545 B.n544 585
R374 B.n543 B.n102 585
R375 B.n542 B.n541 585
R376 B.n540 B.n103 585
R377 B.n539 B.n538 585
R378 B.n537 B.n104 585
R379 B.n536 B.n535 585
R380 B.n534 B.n105 585
R381 B.n533 B.n532 585
R382 B.n531 B.n106 585
R383 B.n530 B.n529 585
R384 B.n528 B.n107 585
R385 B.n527 B.n526 585
R386 B.n525 B.n108 585
R387 B.n524 B.n523 585
R388 B.n522 B.n109 585
R389 B.n521 B.n520 585
R390 B.n519 B.n110 585
R391 B.n518 B.n517 585
R392 B.n516 B.n111 585
R393 B.n515 B.n514 585
R394 B.n513 B.n112 585
R395 B.n512 B.n511 585
R396 B.n510 B.n113 585
R397 B.n509 B.n508 585
R398 B.n507 B.n114 585
R399 B.n506 B.n505 585
R400 B.n504 B.n115 585
R401 B.n503 B.n502 585
R402 B.n501 B.n116 585
R403 B.n500 B.n499 585
R404 B.n498 B.n117 585
R405 B.n497 B.n496 585
R406 B.n495 B.n118 585
R407 B.n494 B.n493 585
R408 B.n492 B.n119 585
R409 B.n491 B.n490 585
R410 B.n489 B.n120 585
R411 B.n488 B.n487 585
R412 B.n486 B.n121 585
R413 B.n485 B.n484 585
R414 B.n483 B.n122 585
R415 B.n482 B.n481 585
R416 B.n480 B.n123 585
R417 B.n479 B.n478 585
R418 B.n477 B.n124 585
R419 B.n476 B.n475 585
R420 B.n474 B.n125 585
R421 B.n473 B.n472 585
R422 B.n471 B.n126 585
R423 B.n470 B.n469 585
R424 B.n468 B.n127 585
R425 B.n467 B.n466 585
R426 B.n465 B.n128 585
R427 B.n464 B.n463 585
R428 B.n462 B.n129 585
R429 B.n461 B.n460 585
R430 B.n459 B.n130 585
R431 B.n279 B.n194 585
R432 B.n281 B.n280 585
R433 B.n282 B.n193 585
R434 B.n284 B.n283 585
R435 B.n285 B.n192 585
R436 B.n287 B.n286 585
R437 B.n288 B.n191 585
R438 B.n290 B.n289 585
R439 B.n291 B.n190 585
R440 B.n293 B.n292 585
R441 B.n294 B.n189 585
R442 B.n296 B.n295 585
R443 B.n297 B.n188 585
R444 B.n299 B.n298 585
R445 B.n300 B.n187 585
R446 B.n302 B.n301 585
R447 B.n303 B.n186 585
R448 B.n305 B.n304 585
R449 B.n306 B.n185 585
R450 B.n308 B.n307 585
R451 B.n309 B.n184 585
R452 B.n311 B.n310 585
R453 B.n312 B.n183 585
R454 B.n314 B.n313 585
R455 B.n315 B.n182 585
R456 B.n317 B.n316 585
R457 B.n318 B.n181 585
R458 B.n320 B.n319 585
R459 B.n321 B.n180 585
R460 B.n323 B.n322 585
R461 B.n324 B.n179 585
R462 B.n326 B.n325 585
R463 B.n327 B.n178 585
R464 B.n329 B.n328 585
R465 B.n330 B.n177 585
R466 B.n332 B.n331 585
R467 B.n333 B.n176 585
R468 B.n335 B.n334 585
R469 B.n336 B.n175 585
R470 B.n338 B.n337 585
R471 B.n339 B.n174 585
R472 B.n341 B.n340 585
R473 B.n342 B.n173 585
R474 B.n344 B.n343 585
R475 B.n345 B.n172 585
R476 B.n347 B.n346 585
R477 B.n348 B.n171 585
R478 B.n350 B.n349 585
R479 B.n351 B.n170 585
R480 B.n353 B.n352 585
R481 B.n354 B.n169 585
R482 B.n356 B.n355 585
R483 B.n357 B.n168 585
R484 B.n359 B.n358 585
R485 B.n360 B.n165 585
R486 B.n363 B.n362 585
R487 B.n364 B.n164 585
R488 B.n366 B.n365 585
R489 B.n367 B.n163 585
R490 B.n369 B.n368 585
R491 B.n370 B.n162 585
R492 B.n372 B.n371 585
R493 B.n373 B.n161 585
R494 B.n375 B.n374 585
R495 B.n377 B.n376 585
R496 B.n378 B.n157 585
R497 B.n380 B.n379 585
R498 B.n381 B.n156 585
R499 B.n383 B.n382 585
R500 B.n384 B.n155 585
R501 B.n386 B.n385 585
R502 B.n387 B.n154 585
R503 B.n389 B.n388 585
R504 B.n390 B.n153 585
R505 B.n392 B.n391 585
R506 B.n393 B.n152 585
R507 B.n395 B.n394 585
R508 B.n396 B.n151 585
R509 B.n398 B.n397 585
R510 B.n399 B.n150 585
R511 B.n401 B.n400 585
R512 B.n402 B.n149 585
R513 B.n404 B.n403 585
R514 B.n405 B.n148 585
R515 B.n407 B.n406 585
R516 B.n408 B.n147 585
R517 B.n410 B.n409 585
R518 B.n411 B.n146 585
R519 B.n413 B.n412 585
R520 B.n414 B.n145 585
R521 B.n416 B.n415 585
R522 B.n417 B.n144 585
R523 B.n419 B.n418 585
R524 B.n420 B.n143 585
R525 B.n422 B.n421 585
R526 B.n423 B.n142 585
R527 B.n425 B.n424 585
R528 B.n426 B.n141 585
R529 B.n428 B.n427 585
R530 B.n429 B.n140 585
R531 B.n431 B.n430 585
R532 B.n432 B.n139 585
R533 B.n434 B.n433 585
R534 B.n435 B.n138 585
R535 B.n437 B.n436 585
R536 B.n438 B.n137 585
R537 B.n440 B.n439 585
R538 B.n441 B.n136 585
R539 B.n443 B.n442 585
R540 B.n444 B.n135 585
R541 B.n446 B.n445 585
R542 B.n447 B.n134 585
R543 B.n449 B.n448 585
R544 B.n450 B.n133 585
R545 B.n452 B.n451 585
R546 B.n453 B.n132 585
R547 B.n455 B.n454 585
R548 B.n456 B.n131 585
R549 B.n458 B.n457 585
R550 B.n278 B.n277 585
R551 B.n276 B.n195 585
R552 B.n275 B.n274 585
R553 B.n273 B.n196 585
R554 B.n272 B.n271 585
R555 B.n270 B.n197 585
R556 B.n269 B.n268 585
R557 B.n267 B.n198 585
R558 B.n266 B.n265 585
R559 B.n264 B.n199 585
R560 B.n263 B.n262 585
R561 B.n261 B.n200 585
R562 B.n260 B.n259 585
R563 B.n258 B.n201 585
R564 B.n257 B.n256 585
R565 B.n255 B.n202 585
R566 B.n254 B.n253 585
R567 B.n252 B.n203 585
R568 B.n251 B.n250 585
R569 B.n249 B.n204 585
R570 B.n248 B.n247 585
R571 B.n246 B.n205 585
R572 B.n245 B.n244 585
R573 B.n243 B.n206 585
R574 B.n242 B.n241 585
R575 B.n240 B.n207 585
R576 B.n239 B.n238 585
R577 B.n237 B.n208 585
R578 B.n236 B.n235 585
R579 B.n234 B.n209 585
R580 B.n233 B.n232 585
R581 B.n231 B.n210 585
R582 B.n230 B.n229 585
R583 B.n228 B.n211 585
R584 B.n227 B.n226 585
R585 B.n225 B.n212 585
R586 B.n224 B.n223 585
R587 B.n222 B.n213 585
R588 B.n221 B.n220 585
R589 B.n219 B.n214 585
R590 B.n218 B.n217 585
R591 B.n216 B.n215 585
R592 B.n2 B.n0 585
R593 B.n833 B.n1 585
R594 B.n832 B.n831 585
R595 B.n830 B.n3 585
R596 B.n829 B.n828 585
R597 B.n827 B.n4 585
R598 B.n826 B.n825 585
R599 B.n824 B.n5 585
R600 B.n823 B.n822 585
R601 B.n821 B.n6 585
R602 B.n820 B.n819 585
R603 B.n818 B.n7 585
R604 B.n817 B.n816 585
R605 B.n815 B.n8 585
R606 B.n814 B.n813 585
R607 B.n812 B.n9 585
R608 B.n811 B.n810 585
R609 B.n809 B.n10 585
R610 B.n808 B.n807 585
R611 B.n806 B.n11 585
R612 B.n805 B.n804 585
R613 B.n803 B.n12 585
R614 B.n802 B.n801 585
R615 B.n800 B.n13 585
R616 B.n799 B.n798 585
R617 B.n797 B.n14 585
R618 B.n796 B.n795 585
R619 B.n794 B.n15 585
R620 B.n793 B.n792 585
R621 B.n791 B.n16 585
R622 B.n790 B.n789 585
R623 B.n788 B.n17 585
R624 B.n787 B.n786 585
R625 B.n785 B.n18 585
R626 B.n784 B.n783 585
R627 B.n782 B.n19 585
R628 B.n781 B.n780 585
R629 B.n779 B.n20 585
R630 B.n778 B.n777 585
R631 B.n776 B.n21 585
R632 B.n775 B.n774 585
R633 B.n773 B.n22 585
R634 B.n772 B.n771 585
R635 B.n770 B.n23 585
R636 B.n835 B.n834 585
R637 B.n279 B.n278 521.33
R638 B.n768 B.n23 521.33
R639 B.n459 B.n458 521.33
R640 B.n590 B.n87 521.33
R641 B.n158 B.t6 399.036
R642 B.n166 B.t9 399.036
R643 B.n52 B.t0 399.036
R644 B.n58 B.t3 399.036
R645 B.n278 B.n195 163.367
R646 B.n274 B.n195 163.367
R647 B.n274 B.n273 163.367
R648 B.n273 B.n272 163.367
R649 B.n272 B.n197 163.367
R650 B.n268 B.n197 163.367
R651 B.n268 B.n267 163.367
R652 B.n267 B.n266 163.367
R653 B.n266 B.n199 163.367
R654 B.n262 B.n199 163.367
R655 B.n262 B.n261 163.367
R656 B.n261 B.n260 163.367
R657 B.n260 B.n201 163.367
R658 B.n256 B.n201 163.367
R659 B.n256 B.n255 163.367
R660 B.n255 B.n254 163.367
R661 B.n254 B.n203 163.367
R662 B.n250 B.n203 163.367
R663 B.n250 B.n249 163.367
R664 B.n249 B.n248 163.367
R665 B.n248 B.n205 163.367
R666 B.n244 B.n205 163.367
R667 B.n244 B.n243 163.367
R668 B.n243 B.n242 163.367
R669 B.n242 B.n207 163.367
R670 B.n238 B.n207 163.367
R671 B.n238 B.n237 163.367
R672 B.n237 B.n236 163.367
R673 B.n236 B.n209 163.367
R674 B.n232 B.n209 163.367
R675 B.n232 B.n231 163.367
R676 B.n231 B.n230 163.367
R677 B.n230 B.n211 163.367
R678 B.n226 B.n211 163.367
R679 B.n226 B.n225 163.367
R680 B.n225 B.n224 163.367
R681 B.n224 B.n213 163.367
R682 B.n220 B.n213 163.367
R683 B.n220 B.n219 163.367
R684 B.n219 B.n218 163.367
R685 B.n218 B.n215 163.367
R686 B.n215 B.n2 163.367
R687 B.n834 B.n2 163.367
R688 B.n834 B.n833 163.367
R689 B.n833 B.n832 163.367
R690 B.n832 B.n3 163.367
R691 B.n828 B.n3 163.367
R692 B.n828 B.n827 163.367
R693 B.n827 B.n826 163.367
R694 B.n826 B.n5 163.367
R695 B.n822 B.n5 163.367
R696 B.n822 B.n821 163.367
R697 B.n821 B.n820 163.367
R698 B.n820 B.n7 163.367
R699 B.n816 B.n7 163.367
R700 B.n816 B.n815 163.367
R701 B.n815 B.n814 163.367
R702 B.n814 B.n9 163.367
R703 B.n810 B.n9 163.367
R704 B.n810 B.n809 163.367
R705 B.n809 B.n808 163.367
R706 B.n808 B.n11 163.367
R707 B.n804 B.n11 163.367
R708 B.n804 B.n803 163.367
R709 B.n803 B.n802 163.367
R710 B.n802 B.n13 163.367
R711 B.n798 B.n13 163.367
R712 B.n798 B.n797 163.367
R713 B.n797 B.n796 163.367
R714 B.n796 B.n15 163.367
R715 B.n792 B.n15 163.367
R716 B.n792 B.n791 163.367
R717 B.n791 B.n790 163.367
R718 B.n790 B.n17 163.367
R719 B.n786 B.n17 163.367
R720 B.n786 B.n785 163.367
R721 B.n785 B.n784 163.367
R722 B.n784 B.n19 163.367
R723 B.n780 B.n19 163.367
R724 B.n780 B.n779 163.367
R725 B.n779 B.n778 163.367
R726 B.n778 B.n21 163.367
R727 B.n774 B.n21 163.367
R728 B.n774 B.n773 163.367
R729 B.n773 B.n772 163.367
R730 B.n772 B.n23 163.367
R731 B.n280 B.n279 163.367
R732 B.n280 B.n193 163.367
R733 B.n284 B.n193 163.367
R734 B.n285 B.n284 163.367
R735 B.n286 B.n285 163.367
R736 B.n286 B.n191 163.367
R737 B.n290 B.n191 163.367
R738 B.n291 B.n290 163.367
R739 B.n292 B.n291 163.367
R740 B.n292 B.n189 163.367
R741 B.n296 B.n189 163.367
R742 B.n297 B.n296 163.367
R743 B.n298 B.n297 163.367
R744 B.n298 B.n187 163.367
R745 B.n302 B.n187 163.367
R746 B.n303 B.n302 163.367
R747 B.n304 B.n303 163.367
R748 B.n304 B.n185 163.367
R749 B.n308 B.n185 163.367
R750 B.n309 B.n308 163.367
R751 B.n310 B.n309 163.367
R752 B.n310 B.n183 163.367
R753 B.n314 B.n183 163.367
R754 B.n315 B.n314 163.367
R755 B.n316 B.n315 163.367
R756 B.n316 B.n181 163.367
R757 B.n320 B.n181 163.367
R758 B.n321 B.n320 163.367
R759 B.n322 B.n321 163.367
R760 B.n322 B.n179 163.367
R761 B.n326 B.n179 163.367
R762 B.n327 B.n326 163.367
R763 B.n328 B.n327 163.367
R764 B.n328 B.n177 163.367
R765 B.n332 B.n177 163.367
R766 B.n333 B.n332 163.367
R767 B.n334 B.n333 163.367
R768 B.n334 B.n175 163.367
R769 B.n338 B.n175 163.367
R770 B.n339 B.n338 163.367
R771 B.n340 B.n339 163.367
R772 B.n340 B.n173 163.367
R773 B.n344 B.n173 163.367
R774 B.n345 B.n344 163.367
R775 B.n346 B.n345 163.367
R776 B.n346 B.n171 163.367
R777 B.n350 B.n171 163.367
R778 B.n351 B.n350 163.367
R779 B.n352 B.n351 163.367
R780 B.n352 B.n169 163.367
R781 B.n356 B.n169 163.367
R782 B.n357 B.n356 163.367
R783 B.n358 B.n357 163.367
R784 B.n358 B.n165 163.367
R785 B.n363 B.n165 163.367
R786 B.n364 B.n363 163.367
R787 B.n365 B.n364 163.367
R788 B.n365 B.n163 163.367
R789 B.n369 B.n163 163.367
R790 B.n370 B.n369 163.367
R791 B.n371 B.n370 163.367
R792 B.n371 B.n161 163.367
R793 B.n375 B.n161 163.367
R794 B.n376 B.n375 163.367
R795 B.n376 B.n157 163.367
R796 B.n380 B.n157 163.367
R797 B.n381 B.n380 163.367
R798 B.n382 B.n381 163.367
R799 B.n382 B.n155 163.367
R800 B.n386 B.n155 163.367
R801 B.n387 B.n386 163.367
R802 B.n388 B.n387 163.367
R803 B.n388 B.n153 163.367
R804 B.n392 B.n153 163.367
R805 B.n393 B.n392 163.367
R806 B.n394 B.n393 163.367
R807 B.n394 B.n151 163.367
R808 B.n398 B.n151 163.367
R809 B.n399 B.n398 163.367
R810 B.n400 B.n399 163.367
R811 B.n400 B.n149 163.367
R812 B.n404 B.n149 163.367
R813 B.n405 B.n404 163.367
R814 B.n406 B.n405 163.367
R815 B.n406 B.n147 163.367
R816 B.n410 B.n147 163.367
R817 B.n411 B.n410 163.367
R818 B.n412 B.n411 163.367
R819 B.n412 B.n145 163.367
R820 B.n416 B.n145 163.367
R821 B.n417 B.n416 163.367
R822 B.n418 B.n417 163.367
R823 B.n418 B.n143 163.367
R824 B.n422 B.n143 163.367
R825 B.n423 B.n422 163.367
R826 B.n424 B.n423 163.367
R827 B.n424 B.n141 163.367
R828 B.n428 B.n141 163.367
R829 B.n429 B.n428 163.367
R830 B.n430 B.n429 163.367
R831 B.n430 B.n139 163.367
R832 B.n434 B.n139 163.367
R833 B.n435 B.n434 163.367
R834 B.n436 B.n435 163.367
R835 B.n436 B.n137 163.367
R836 B.n440 B.n137 163.367
R837 B.n441 B.n440 163.367
R838 B.n442 B.n441 163.367
R839 B.n442 B.n135 163.367
R840 B.n446 B.n135 163.367
R841 B.n447 B.n446 163.367
R842 B.n448 B.n447 163.367
R843 B.n448 B.n133 163.367
R844 B.n452 B.n133 163.367
R845 B.n453 B.n452 163.367
R846 B.n454 B.n453 163.367
R847 B.n454 B.n131 163.367
R848 B.n458 B.n131 163.367
R849 B.n460 B.n459 163.367
R850 B.n460 B.n129 163.367
R851 B.n464 B.n129 163.367
R852 B.n465 B.n464 163.367
R853 B.n466 B.n465 163.367
R854 B.n466 B.n127 163.367
R855 B.n470 B.n127 163.367
R856 B.n471 B.n470 163.367
R857 B.n472 B.n471 163.367
R858 B.n472 B.n125 163.367
R859 B.n476 B.n125 163.367
R860 B.n477 B.n476 163.367
R861 B.n478 B.n477 163.367
R862 B.n478 B.n123 163.367
R863 B.n482 B.n123 163.367
R864 B.n483 B.n482 163.367
R865 B.n484 B.n483 163.367
R866 B.n484 B.n121 163.367
R867 B.n488 B.n121 163.367
R868 B.n489 B.n488 163.367
R869 B.n490 B.n489 163.367
R870 B.n490 B.n119 163.367
R871 B.n494 B.n119 163.367
R872 B.n495 B.n494 163.367
R873 B.n496 B.n495 163.367
R874 B.n496 B.n117 163.367
R875 B.n500 B.n117 163.367
R876 B.n501 B.n500 163.367
R877 B.n502 B.n501 163.367
R878 B.n502 B.n115 163.367
R879 B.n506 B.n115 163.367
R880 B.n507 B.n506 163.367
R881 B.n508 B.n507 163.367
R882 B.n508 B.n113 163.367
R883 B.n512 B.n113 163.367
R884 B.n513 B.n512 163.367
R885 B.n514 B.n513 163.367
R886 B.n514 B.n111 163.367
R887 B.n518 B.n111 163.367
R888 B.n519 B.n518 163.367
R889 B.n520 B.n519 163.367
R890 B.n520 B.n109 163.367
R891 B.n524 B.n109 163.367
R892 B.n525 B.n524 163.367
R893 B.n526 B.n525 163.367
R894 B.n526 B.n107 163.367
R895 B.n530 B.n107 163.367
R896 B.n531 B.n530 163.367
R897 B.n532 B.n531 163.367
R898 B.n532 B.n105 163.367
R899 B.n536 B.n105 163.367
R900 B.n537 B.n536 163.367
R901 B.n538 B.n537 163.367
R902 B.n538 B.n103 163.367
R903 B.n542 B.n103 163.367
R904 B.n543 B.n542 163.367
R905 B.n544 B.n543 163.367
R906 B.n544 B.n101 163.367
R907 B.n548 B.n101 163.367
R908 B.n549 B.n548 163.367
R909 B.n550 B.n549 163.367
R910 B.n550 B.n99 163.367
R911 B.n554 B.n99 163.367
R912 B.n555 B.n554 163.367
R913 B.n556 B.n555 163.367
R914 B.n556 B.n97 163.367
R915 B.n560 B.n97 163.367
R916 B.n561 B.n560 163.367
R917 B.n562 B.n561 163.367
R918 B.n562 B.n95 163.367
R919 B.n566 B.n95 163.367
R920 B.n567 B.n566 163.367
R921 B.n568 B.n567 163.367
R922 B.n568 B.n93 163.367
R923 B.n572 B.n93 163.367
R924 B.n573 B.n572 163.367
R925 B.n574 B.n573 163.367
R926 B.n574 B.n91 163.367
R927 B.n578 B.n91 163.367
R928 B.n579 B.n578 163.367
R929 B.n580 B.n579 163.367
R930 B.n580 B.n89 163.367
R931 B.n584 B.n89 163.367
R932 B.n585 B.n584 163.367
R933 B.n586 B.n585 163.367
R934 B.n586 B.n87 163.367
R935 B.n768 B.n767 163.367
R936 B.n767 B.n766 163.367
R937 B.n766 B.n25 163.367
R938 B.n762 B.n25 163.367
R939 B.n762 B.n761 163.367
R940 B.n761 B.n760 163.367
R941 B.n760 B.n27 163.367
R942 B.n756 B.n27 163.367
R943 B.n756 B.n755 163.367
R944 B.n755 B.n754 163.367
R945 B.n754 B.n29 163.367
R946 B.n750 B.n29 163.367
R947 B.n750 B.n749 163.367
R948 B.n749 B.n748 163.367
R949 B.n748 B.n31 163.367
R950 B.n744 B.n31 163.367
R951 B.n744 B.n743 163.367
R952 B.n743 B.n742 163.367
R953 B.n742 B.n33 163.367
R954 B.n738 B.n33 163.367
R955 B.n738 B.n737 163.367
R956 B.n737 B.n736 163.367
R957 B.n736 B.n35 163.367
R958 B.n732 B.n35 163.367
R959 B.n732 B.n731 163.367
R960 B.n731 B.n730 163.367
R961 B.n730 B.n37 163.367
R962 B.n726 B.n37 163.367
R963 B.n726 B.n725 163.367
R964 B.n725 B.n724 163.367
R965 B.n724 B.n39 163.367
R966 B.n720 B.n39 163.367
R967 B.n720 B.n719 163.367
R968 B.n719 B.n718 163.367
R969 B.n718 B.n41 163.367
R970 B.n714 B.n41 163.367
R971 B.n714 B.n713 163.367
R972 B.n713 B.n712 163.367
R973 B.n712 B.n43 163.367
R974 B.n708 B.n43 163.367
R975 B.n708 B.n707 163.367
R976 B.n707 B.n706 163.367
R977 B.n706 B.n45 163.367
R978 B.n702 B.n45 163.367
R979 B.n702 B.n701 163.367
R980 B.n701 B.n700 163.367
R981 B.n700 B.n47 163.367
R982 B.n696 B.n47 163.367
R983 B.n696 B.n695 163.367
R984 B.n695 B.n694 163.367
R985 B.n694 B.n49 163.367
R986 B.n690 B.n49 163.367
R987 B.n690 B.n689 163.367
R988 B.n689 B.n688 163.367
R989 B.n688 B.n51 163.367
R990 B.n683 B.n51 163.367
R991 B.n683 B.n682 163.367
R992 B.n682 B.n681 163.367
R993 B.n681 B.n55 163.367
R994 B.n677 B.n55 163.367
R995 B.n677 B.n676 163.367
R996 B.n676 B.n675 163.367
R997 B.n675 B.n57 163.367
R998 B.n670 B.n57 163.367
R999 B.n670 B.n669 163.367
R1000 B.n669 B.n668 163.367
R1001 B.n668 B.n61 163.367
R1002 B.n664 B.n61 163.367
R1003 B.n664 B.n663 163.367
R1004 B.n663 B.n662 163.367
R1005 B.n662 B.n63 163.367
R1006 B.n658 B.n63 163.367
R1007 B.n658 B.n657 163.367
R1008 B.n657 B.n656 163.367
R1009 B.n656 B.n65 163.367
R1010 B.n652 B.n65 163.367
R1011 B.n652 B.n651 163.367
R1012 B.n651 B.n650 163.367
R1013 B.n650 B.n67 163.367
R1014 B.n646 B.n67 163.367
R1015 B.n646 B.n645 163.367
R1016 B.n645 B.n644 163.367
R1017 B.n644 B.n69 163.367
R1018 B.n640 B.n69 163.367
R1019 B.n640 B.n639 163.367
R1020 B.n639 B.n638 163.367
R1021 B.n638 B.n71 163.367
R1022 B.n634 B.n71 163.367
R1023 B.n634 B.n633 163.367
R1024 B.n633 B.n632 163.367
R1025 B.n632 B.n73 163.367
R1026 B.n628 B.n73 163.367
R1027 B.n628 B.n627 163.367
R1028 B.n627 B.n626 163.367
R1029 B.n626 B.n75 163.367
R1030 B.n622 B.n75 163.367
R1031 B.n622 B.n621 163.367
R1032 B.n621 B.n620 163.367
R1033 B.n620 B.n77 163.367
R1034 B.n616 B.n77 163.367
R1035 B.n616 B.n615 163.367
R1036 B.n615 B.n614 163.367
R1037 B.n614 B.n79 163.367
R1038 B.n610 B.n79 163.367
R1039 B.n610 B.n609 163.367
R1040 B.n609 B.n608 163.367
R1041 B.n608 B.n81 163.367
R1042 B.n604 B.n81 163.367
R1043 B.n604 B.n603 163.367
R1044 B.n603 B.n602 163.367
R1045 B.n602 B.n83 163.367
R1046 B.n598 B.n83 163.367
R1047 B.n598 B.n597 163.367
R1048 B.n597 B.n596 163.367
R1049 B.n596 B.n85 163.367
R1050 B.n592 B.n85 163.367
R1051 B.n592 B.n591 163.367
R1052 B.n591 B.n590 163.367
R1053 B.n158 B.t8 154.474
R1054 B.n58 B.t4 154.474
R1055 B.n166 B.t11 154.452
R1056 B.n52 B.t1 154.452
R1057 B.n159 B.t7 108.123
R1058 B.n59 B.t5 108.123
R1059 B.n167 B.t10 108.102
R1060 B.n53 B.t2 108.102
R1061 B.n160 B.n159 59.5399
R1062 B.n361 B.n167 59.5399
R1063 B.n686 B.n53 59.5399
R1064 B.n672 B.n59 59.5399
R1065 B.n159 B.n158 46.352
R1066 B.n167 B.n166 46.352
R1067 B.n53 B.n52 46.352
R1068 B.n59 B.n58 46.352
R1069 B.n770 B.n769 33.8737
R1070 B.n589 B.n588 33.8737
R1071 B.n457 B.n130 33.8737
R1072 B.n277 B.n194 33.8737
R1073 B B.n835 18.0485
R1074 B.n769 B.n24 10.6151
R1075 B.n765 B.n24 10.6151
R1076 B.n765 B.n764 10.6151
R1077 B.n764 B.n763 10.6151
R1078 B.n763 B.n26 10.6151
R1079 B.n759 B.n26 10.6151
R1080 B.n759 B.n758 10.6151
R1081 B.n758 B.n757 10.6151
R1082 B.n757 B.n28 10.6151
R1083 B.n753 B.n28 10.6151
R1084 B.n753 B.n752 10.6151
R1085 B.n752 B.n751 10.6151
R1086 B.n751 B.n30 10.6151
R1087 B.n747 B.n30 10.6151
R1088 B.n747 B.n746 10.6151
R1089 B.n746 B.n745 10.6151
R1090 B.n745 B.n32 10.6151
R1091 B.n741 B.n32 10.6151
R1092 B.n741 B.n740 10.6151
R1093 B.n740 B.n739 10.6151
R1094 B.n739 B.n34 10.6151
R1095 B.n735 B.n34 10.6151
R1096 B.n735 B.n734 10.6151
R1097 B.n734 B.n733 10.6151
R1098 B.n733 B.n36 10.6151
R1099 B.n729 B.n36 10.6151
R1100 B.n729 B.n728 10.6151
R1101 B.n728 B.n727 10.6151
R1102 B.n727 B.n38 10.6151
R1103 B.n723 B.n38 10.6151
R1104 B.n723 B.n722 10.6151
R1105 B.n722 B.n721 10.6151
R1106 B.n721 B.n40 10.6151
R1107 B.n717 B.n40 10.6151
R1108 B.n717 B.n716 10.6151
R1109 B.n716 B.n715 10.6151
R1110 B.n715 B.n42 10.6151
R1111 B.n711 B.n42 10.6151
R1112 B.n711 B.n710 10.6151
R1113 B.n710 B.n709 10.6151
R1114 B.n709 B.n44 10.6151
R1115 B.n705 B.n44 10.6151
R1116 B.n705 B.n704 10.6151
R1117 B.n704 B.n703 10.6151
R1118 B.n703 B.n46 10.6151
R1119 B.n699 B.n46 10.6151
R1120 B.n699 B.n698 10.6151
R1121 B.n698 B.n697 10.6151
R1122 B.n697 B.n48 10.6151
R1123 B.n693 B.n48 10.6151
R1124 B.n693 B.n692 10.6151
R1125 B.n692 B.n691 10.6151
R1126 B.n691 B.n50 10.6151
R1127 B.n687 B.n50 10.6151
R1128 B.n685 B.n684 10.6151
R1129 B.n684 B.n54 10.6151
R1130 B.n680 B.n54 10.6151
R1131 B.n680 B.n679 10.6151
R1132 B.n679 B.n678 10.6151
R1133 B.n678 B.n56 10.6151
R1134 B.n674 B.n56 10.6151
R1135 B.n674 B.n673 10.6151
R1136 B.n671 B.n60 10.6151
R1137 B.n667 B.n60 10.6151
R1138 B.n667 B.n666 10.6151
R1139 B.n666 B.n665 10.6151
R1140 B.n665 B.n62 10.6151
R1141 B.n661 B.n62 10.6151
R1142 B.n661 B.n660 10.6151
R1143 B.n660 B.n659 10.6151
R1144 B.n659 B.n64 10.6151
R1145 B.n655 B.n64 10.6151
R1146 B.n655 B.n654 10.6151
R1147 B.n654 B.n653 10.6151
R1148 B.n653 B.n66 10.6151
R1149 B.n649 B.n66 10.6151
R1150 B.n649 B.n648 10.6151
R1151 B.n648 B.n647 10.6151
R1152 B.n647 B.n68 10.6151
R1153 B.n643 B.n68 10.6151
R1154 B.n643 B.n642 10.6151
R1155 B.n642 B.n641 10.6151
R1156 B.n641 B.n70 10.6151
R1157 B.n637 B.n70 10.6151
R1158 B.n637 B.n636 10.6151
R1159 B.n636 B.n635 10.6151
R1160 B.n635 B.n72 10.6151
R1161 B.n631 B.n72 10.6151
R1162 B.n631 B.n630 10.6151
R1163 B.n630 B.n629 10.6151
R1164 B.n629 B.n74 10.6151
R1165 B.n625 B.n74 10.6151
R1166 B.n625 B.n624 10.6151
R1167 B.n624 B.n623 10.6151
R1168 B.n623 B.n76 10.6151
R1169 B.n619 B.n76 10.6151
R1170 B.n619 B.n618 10.6151
R1171 B.n618 B.n617 10.6151
R1172 B.n617 B.n78 10.6151
R1173 B.n613 B.n78 10.6151
R1174 B.n613 B.n612 10.6151
R1175 B.n612 B.n611 10.6151
R1176 B.n611 B.n80 10.6151
R1177 B.n607 B.n80 10.6151
R1178 B.n607 B.n606 10.6151
R1179 B.n606 B.n605 10.6151
R1180 B.n605 B.n82 10.6151
R1181 B.n601 B.n82 10.6151
R1182 B.n601 B.n600 10.6151
R1183 B.n600 B.n599 10.6151
R1184 B.n599 B.n84 10.6151
R1185 B.n595 B.n84 10.6151
R1186 B.n595 B.n594 10.6151
R1187 B.n594 B.n593 10.6151
R1188 B.n593 B.n86 10.6151
R1189 B.n589 B.n86 10.6151
R1190 B.n461 B.n130 10.6151
R1191 B.n462 B.n461 10.6151
R1192 B.n463 B.n462 10.6151
R1193 B.n463 B.n128 10.6151
R1194 B.n467 B.n128 10.6151
R1195 B.n468 B.n467 10.6151
R1196 B.n469 B.n468 10.6151
R1197 B.n469 B.n126 10.6151
R1198 B.n473 B.n126 10.6151
R1199 B.n474 B.n473 10.6151
R1200 B.n475 B.n474 10.6151
R1201 B.n475 B.n124 10.6151
R1202 B.n479 B.n124 10.6151
R1203 B.n480 B.n479 10.6151
R1204 B.n481 B.n480 10.6151
R1205 B.n481 B.n122 10.6151
R1206 B.n485 B.n122 10.6151
R1207 B.n486 B.n485 10.6151
R1208 B.n487 B.n486 10.6151
R1209 B.n487 B.n120 10.6151
R1210 B.n491 B.n120 10.6151
R1211 B.n492 B.n491 10.6151
R1212 B.n493 B.n492 10.6151
R1213 B.n493 B.n118 10.6151
R1214 B.n497 B.n118 10.6151
R1215 B.n498 B.n497 10.6151
R1216 B.n499 B.n498 10.6151
R1217 B.n499 B.n116 10.6151
R1218 B.n503 B.n116 10.6151
R1219 B.n504 B.n503 10.6151
R1220 B.n505 B.n504 10.6151
R1221 B.n505 B.n114 10.6151
R1222 B.n509 B.n114 10.6151
R1223 B.n510 B.n509 10.6151
R1224 B.n511 B.n510 10.6151
R1225 B.n511 B.n112 10.6151
R1226 B.n515 B.n112 10.6151
R1227 B.n516 B.n515 10.6151
R1228 B.n517 B.n516 10.6151
R1229 B.n517 B.n110 10.6151
R1230 B.n521 B.n110 10.6151
R1231 B.n522 B.n521 10.6151
R1232 B.n523 B.n522 10.6151
R1233 B.n523 B.n108 10.6151
R1234 B.n527 B.n108 10.6151
R1235 B.n528 B.n527 10.6151
R1236 B.n529 B.n528 10.6151
R1237 B.n529 B.n106 10.6151
R1238 B.n533 B.n106 10.6151
R1239 B.n534 B.n533 10.6151
R1240 B.n535 B.n534 10.6151
R1241 B.n535 B.n104 10.6151
R1242 B.n539 B.n104 10.6151
R1243 B.n540 B.n539 10.6151
R1244 B.n541 B.n540 10.6151
R1245 B.n541 B.n102 10.6151
R1246 B.n545 B.n102 10.6151
R1247 B.n546 B.n545 10.6151
R1248 B.n547 B.n546 10.6151
R1249 B.n547 B.n100 10.6151
R1250 B.n551 B.n100 10.6151
R1251 B.n552 B.n551 10.6151
R1252 B.n553 B.n552 10.6151
R1253 B.n553 B.n98 10.6151
R1254 B.n557 B.n98 10.6151
R1255 B.n558 B.n557 10.6151
R1256 B.n559 B.n558 10.6151
R1257 B.n559 B.n96 10.6151
R1258 B.n563 B.n96 10.6151
R1259 B.n564 B.n563 10.6151
R1260 B.n565 B.n564 10.6151
R1261 B.n565 B.n94 10.6151
R1262 B.n569 B.n94 10.6151
R1263 B.n570 B.n569 10.6151
R1264 B.n571 B.n570 10.6151
R1265 B.n571 B.n92 10.6151
R1266 B.n575 B.n92 10.6151
R1267 B.n576 B.n575 10.6151
R1268 B.n577 B.n576 10.6151
R1269 B.n577 B.n90 10.6151
R1270 B.n581 B.n90 10.6151
R1271 B.n582 B.n581 10.6151
R1272 B.n583 B.n582 10.6151
R1273 B.n583 B.n88 10.6151
R1274 B.n587 B.n88 10.6151
R1275 B.n588 B.n587 10.6151
R1276 B.n281 B.n194 10.6151
R1277 B.n282 B.n281 10.6151
R1278 B.n283 B.n282 10.6151
R1279 B.n283 B.n192 10.6151
R1280 B.n287 B.n192 10.6151
R1281 B.n288 B.n287 10.6151
R1282 B.n289 B.n288 10.6151
R1283 B.n289 B.n190 10.6151
R1284 B.n293 B.n190 10.6151
R1285 B.n294 B.n293 10.6151
R1286 B.n295 B.n294 10.6151
R1287 B.n295 B.n188 10.6151
R1288 B.n299 B.n188 10.6151
R1289 B.n300 B.n299 10.6151
R1290 B.n301 B.n300 10.6151
R1291 B.n301 B.n186 10.6151
R1292 B.n305 B.n186 10.6151
R1293 B.n306 B.n305 10.6151
R1294 B.n307 B.n306 10.6151
R1295 B.n307 B.n184 10.6151
R1296 B.n311 B.n184 10.6151
R1297 B.n312 B.n311 10.6151
R1298 B.n313 B.n312 10.6151
R1299 B.n313 B.n182 10.6151
R1300 B.n317 B.n182 10.6151
R1301 B.n318 B.n317 10.6151
R1302 B.n319 B.n318 10.6151
R1303 B.n319 B.n180 10.6151
R1304 B.n323 B.n180 10.6151
R1305 B.n324 B.n323 10.6151
R1306 B.n325 B.n324 10.6151
R1307 B.n325 B.n178 10.6151
R1308 B.n329 B.n178 10.6151
R1309 B.n330 B.n329 10.6151
R1310 B.n331 B.n330 10.6151
R1311 B.n331 B.n176 10.6151
R1312 B.n335 B.n176 10.6151
R1313 B.n336 B.n335 10.6151
R1314 B.n337 B.n336 10.6151
R1315 B.n337 B.n174 10.6151
R1316 B.n341 B.n174 10.6151
R1317 B.n342 B.n341 10.6151
R1318 B.n343 B.n342 10.6151
R1319 B.n343 B.n172 10.6151
R1320 B.n347 B.n172 10.6151
R1321 B.n348 B.n347 10.6151
R1322 B.n349 B.n348 10.6151
R1323 B.n349 B.n170 10.6151
R1324 B.n353 B.n170 10.6151
R1325 B.n354 B.n353 10.6151
R1326 B.n355 B.n354 10.6151
R1327 B.n355 B.n168 10.6151
R1328 B.n359 B.n168 10.6151
R1329 B.n360 B.n359 10.6151
R1330 B.n362 B.n164 10.6151
R1331 B.n366 B.n164 10.6151
R1332 B.n367 B.n366 10.6151
R1333 B.n368 B.n367 10.6151
R1334 B.n368 B.n162 10.6151
R1335 B.n372 B.n162 10.6151
R1336 B.n373 B.n372 10.6151
R1337 B.n374 B.n373 10.6151
R1338 B.n378 B.n377 10.6151
R1339 B.n379 B.n378 10.6151
R1340 B.n379 B.n156 10.6151
R1341 B.n383 B.n156 10.6151
R1342 B.n384 B.n383 10.6151
R1343 B.n385 B.n384 10.6151
R1344 B.n385 B.n154 10.6151
R1345 B.n389 B.n154 10.6151
R1346 B.n390 B.n389 10.6151
R1347 B.n391 B.n390 10.6151
R1348 B.n391 B.n152 10.6151
R1349 B.n395 B.n152 10.6151
R1350 B.n396 B.n395 10.6151
R1351 B.n397 B.n396 10.6151
R1352 B.n397 B.n150 10.6151
R1353 B.n401 B.n150 10.6151
R1354 B.n402 B.n401 10.6151
R1355 B.n403 B.n402 10.6151
R1356 B.n403 B.n148 10.6151
R1357 B.n407 B.n148 10.6151
R1358 B.n408 B.n407 10.6151
R1359 B.n409 B.n408 10.6151
R1360 B.n409 B.n146 10.6151
R1361 B.n413 B.n146 10.6151
R1362 B.n414 B.n413 10.6151
R1363 B.n415 B.n414 10.6151
R1364 B.n415 B.n144 10.6151
R1365 B.n419 B.n144 10.6151
R1366 B.n420 B.n419 10.6151
R1367 B.n421 B.n420 10.6151
R1368 B.n421 B.n142 10.6151
R1369 B.n425 B.n142 10.6151
R1370 B.n426 B.n425 10.6151
R1371 B.n427 B.n426 10.6151
R1372 B.n427 B.n140 10.6151
R1373 B.n431 B.n140 10.6151
R1374 B.n432 B.n431 10.6151
R1375 B.n433 B.n432 10.6151
R1376 B.n433 B.n138 10.6151
R1377 B.n437 B.n138 10.6151
R1378 B.n438 B.n437 10.6151
R1379 B.n439 B.n438 10.6151
R1380 B.n439 B.n136 10.6151
R1381 B.n443 B.n136 10.6151
R1382 B.n444 B.n443 10.6151
R1383 B.n445 B.n444 10.6151
R1384 B.n445 B.n134 10.6151
R1385 B.n449 B.n134 10.6151
R1386 B.n450 B.n449 10.6151
R1387 B.n451 B.n450 10.6151
R1388 B.n451 B.n132 10.6151
R1389 B.n455 B.n132 10.6151
R1390 B.n456 B.n455 10.6151
R1391 B.n457 B.n456 10.6151
R1392 B.n277 B.n276 10.6151
R1393 B.n276 B.n275 10.6151
R1394 B.n275 B.n196 10.6151
R1395 B.n271 B.n196 10.6151
R1396 B.n271 B.n270 10.6151
R1397 B.n270 B.n269 10.6151
R1398 B.n269 B.n198 10.6151
R1399 B.n265 B.n198 10.6151
R1400 B.n265 B.n264 10.6151
R1401 B.n264 B.n263 10.6151
R1402 B.n263 B.n200 10.6151
R1403 B.n259 B.n200 10.6151
R1404 B.n259 B.n258 10.6151
R1405 B.n258 B.n257 10.6151
R1406 B.n257 B.n202 10.6151
R1407 B.n253 B.n202 10.6151
R1408 B.n253 B.n252 10.6151
R1409 B.n252 B.n251 10.6151
R1410 B.n251 B.n204 10.6151
R1411 B.n247 B.n204 10.6151
R1412 B.n247 B.n246 10.6151
R1413 B.n246 B.n245 10.6151
R1414 B.n245 B.n206 10.6151
R1415 B.n241 B.n206 10.6151
R1416 B.n241 B.n240 10.6151
R1417 B.n240 B.n239 10.6151
R1418 B.n239 B.n208 10.6151
R1419 B.n235 B.n208 10.6151
R1420 B.n235 B.n234 10.6151
R1421 B.n234 B.n233 10.6151
R1422 B.n233 B.n210 10.6151
R1423 B.n229 B.n210 10.6151
R1424 B.n229 B.n228 10.6151
R1425 B.n228 B.n227 10.6151
R1426 B.n227 B.n212 10.6151
R1427 B.n223 B.n212 10.6151
R1428 B.n223 B.n222 10.6151
R1429 B.n222 B.n221 10.6151
R1430 B.n221 B.n214 10.6151
R1431 B.n217 B.n214 10.6151
R1432 B.n217 B.n216 10.6151
R1433 B.n216 B.n0 10.6151
R1434 B.n831 B.n1 10.6151
R1435 B.n831 B.n830 10.6151
R1436 B.n830 B.n829 10.6151
R1437 B.n829 B.n4 10.6151
R1438 B.n825 B.n4 10.6151
R1439 B.n825 B.n824 10.6151
R1440 B.n824 B.n823 10.6151
R1441 B.n823 B.n6 10.6151
R1442 B.n819 B.n6 10.6151
R1443 B.n819 B.n818 10.6151
R1444 B.n818 B.n817 10.6151
R1445 B.n817 B.n8 10.6151
R1446 B.n813 B.n8 10.6151
R1447 B.n813 B.n812 10.6151
R1448 B.n812 B.n811 10.6151
R1449 B.n811 B.n10 10.6151
R1450 B.n807 B.n10 10.6151
R1451 B.n807 B.n806 10.6151
R1452 B.n806 B.n805 10.6151
R1453 B.n805 B.n12 10.6151
R1454 B.n801 B.n12 10.6151
R1455 B.n801 B.n800 10.6151
R1456 B.n800 B.n799 10.6151
R1457 B.n799 B.n14 10.6151
R1458 B.n795 B.n14 10.6151
R1459 B.n795 B.n794 10.6151
R1460 B.n794 B.n793 10.6151
R1461 B.n793 B.n16 10.6151
R1462 B.n789 B.n16 10.6151
R1463 B.n789 B.n788 10.6151
R1464 B.n788 B.n787 10.6151
R1465 B.n787 B.n18 10.6151
R1466 B.n783 B.n18 10.6151
R1467 B.n783 B.n782 10.6151
R1468 B.n782 B.n781 10.6151
R1469 B.n781 B.n20 10.6151
R1470 B.n777 B.n20 10.6151
R1471 B.n777 B.n776 10.6151
R1472 B.n776 B.n775 10.6151
R1473 B.n775 B.n22 10.6151
R1474 B.n771 B.n22 10.6151
R1475 B.n771 B.n770 10.6151
R1476 B.n686 B.n685 6.5566
R1477 B.n673 B.n672 6.5566
R1478 B.n362 B.n361 6.5566
R1479 B.n374 B.n160 6.5566
R1480 B.n687 B.n686 4.05904
R1481 B.n672 B.n671 4.05904
R1482 B.n361 B.n360 4.05904
R1483 B.n377 B.n160 4.05904
R1484 B.n835 B.n0 2.81026
R1485 B.n835 B.n1 2.81026
C0 VP VDD1 11.4479f
C1 VP B 1.87704f
C2 B VDD1 1.60449f
C3 VDD2 VP 0.46219f
C4 VDD2 VDD1 1.49626f
C5 VN VTAIL 11.1724f
C6 w_n3360_n4250# VN 6.77449f
C7 VDD2 B 1.68353f
C8 w_n3360_n4250# VTAIL 5.19131f
C9 VP VN 7.82188f
C10 VN VDD1 0.150733f
C11 VP VTAIL 11.1865f
C12 VTAIL VDD1 9.77569f
C13 VN B 1.15137f
C14 w_n3360_n4250# VP 7.2091f
C15 w_n3360_n4250# VDD1 1.8974f
C16 B VTAIL 6.1157f
C17 VDD2 VN 11.1375f
C18 VDD2 VTAIL 9.82649f
C19 w_n3360_n4250# B 10.525099f
C20 w_n3360_n4250# VDD2 1.98946f
C21 VDD2 VSUBS 1.770167f
C22 VDD1 VSUBS 2.322464f
C23 VTAIL VSUBS 1.449225f
C24 VN VSUBS 6.26391f
C25 VP VSUBS 3.197766f
C26 B VSUBS 4.770194f
C27 w_n3360_n4250# VSUBS 0.174868p
C28 B.n0 VSUBS 0.004128f
C29 B.n1 VSUBS 0.004128f
C30 B.n2 VSUBS 0.006528f
C31 B.n3 VSUBS 0.006528f
C32 B.n4 VSUBS 0.006528f
C33 B.n5 VSUBS 0.006528f
C34 B.n6 VSUBS 0.006528f
C35 B.n7 VSUBS 0.006528f
C36 B.n8 VSUBS 0.006528f
C37 B.n9 VSUBS 0.006528f
C38 B.n10 VSUBS 0.006528f
C39 B.n11 VSUBS 0.006528f
C40 B.n12 VSUBS 0.006528f
C41 B.n13 VSUBS 0.006528f
C42 B.n14 VSUBS 0.006528f
C43 B.n15 VSUBS 0.006528f
C44 B.n16 VSUBS 0.006528f
C45 B.n17 VSUBS 0.006528f
C46 B.n18 VSUBS 0.006528f
C47 B.n19 VSUBS 0.006528f
C48 B.n20 VSUBS 0.006528f
C49 B.n21 VSUBS 0.006528f
C50 B.n22 VSUBS 0.006528f
C51 B.n23 VSUBS 0.015059f
C52 B.n24 VSUBS 0.006528f
C53 B.n25 VSUBS 0.006528f
C54 B.n26 VSUBS 0.006528f
C55 B.n27 VSUBS 0.006528f
C56 B.n28 VSUBS 0.006528f
C57 B.n29 VSUBS 0.006528f
C58 B.n30 VSUBS 0.006528f
C59 B.n31 VSUBS 0.006528f
C60 B.n32 VSUBS 0.006528f
C61 B.n33 VSUBS 0.006528f
C62 B.n34 VSUBS 0.006528f
C63 B.n35 VSUBS 0.006528f
C64 B.n36 VSUBS 0.006528f
C65 B.n37 VSUBS 0.006528f
C66 B.n38 VSUBS 0.006528f
C67 B.n39 VSUBS 0.006528f
C68 B.n40 VSUBS 0.006528f
C69 B.n41 VSUBS 0.006528f
C70 B.n42 VSUBS 0.006528f
C71 B.n43 VSUBS 0.006528f
C72 B.n44 VSUBS 0.006528f
C73 B.n45 VSUBS 0.006528f
C74 B.n46 VSUBS 0.006528f
C75 B.n47 VSUBS 0.006528f
C76 B.n48 VSUBS 0.006528f
C77 B.n49 VSUBS 0.006528f
C78 B.n50 VSUBS 0.006528f
C79 B.n51 VSUBS 0.006528f
C80 B.t2 VSUBS 0.513158f
C81 B.t1 VSUBS 0.529906f
C82 B.t0 VSUBS 1.38281f
C83 B.n52 VSUBS 0.262921f
C84 B.n53 VSUBS 0.065118f
C85 B.n54 VSUBS 0.006528f
C86 B.n55 VSUBS 0.006528f
C87 B.n56 VSUBS 0.006528f
C88 B.n57 VSUBS 0.006528f
C89 B.t5 VSUBS 0.513142f
C90 B.t4 VSUBS 0.529892f
C91 B.t3 VSUBS 1.38281f
C92 B.n58 VSUBS 0.262935f
C93 B.n59 VSUBS 0.065135f
C94 B.n60 VSUBS 0.006528f
C95 B.n61 VSUBS 0.006528f
C96 B.n62 VSUBS 0.006528f
C97 B.n63 VSUBS 0.006528f
C98 B.n64 VSUBS 0.006528f
C99 B.n65 VSUBS 0.006528f
C100 B.n66 VSUBS 0.006528f
C101 B.n67 VSUBS 0.006528f
C102 B.n68 VSUBS 0.006528f
C103 B.n69 VSUBS 0.006528f
C104 B.n70 VSUBS 0.006528f
C105 B.n71 VSUBS 0.006528f
C106 B.n72 VSUBS 0.006528f
C107 B.n73 VSUBS 0.006528f
C108 B.n74 VSUBS 0.006528f
C109 B.n75 VSUBS 0.006528f
C110 B.n76 VSUBS 0.006528f
C111 B.n77 VSUBS 0.006528f
C112 B.n78 VSUBS 0.006528f
C113 B.n79 VSUBS 0.006528f
C114 B.n80 VSUBS 0.006528f
C115 B.n81 VSUBS 0.006528f
C116 B.n82 VSUBS 0.006528f
C117 B.n83 VSUBS 0.006528f
C118 B.n84 VSUBS 0.006528f
C119 B.n85 VSUBS 0.006528f
C120 B.n86 VSUBS 0.006528f
C121 B.n87 VSUBS 0.015059f
C122 B.n88 VSUBS 0.006528f
C123 B.n89 VSUBS 0.006528f
C124 B.n90 VSUBS 0.006528f
C125 B.n91 VSUBS 0.006528f
C126 B.n92 VSUBS 0.006528f
C127 B.n93 VSUBS 0.006528f
C128 B.n94 VSUBS 0.006528f
C129 B.n95 VSUBS 0.006528f
C130 B.n96 VSUBS 0.006528f
C131 B.n97 VSUBS 0.006528f
C132 B.n98 VSUBS 0.006528f
C133 B.n99 VSUBS 0.006528f
C134 B.n100 VSUBS 0.006528f
C135 B.n101 VSUBS 0.006528f
C136 B.n102 VSUBS 0.006528f
C137 B.n103 VSUBS 0.006528f
C138 B.n104 VSUBS 0.006528f
C139 B.n105 VSUBS 0.006528f
C140 B.n106 VSUBS 0.006528f
C141 B.n107 VSUBS 0.006528f
C142 B.n108 VSUBS 0.006528f
C143 B.n109 VSUBS 0.006528f
C144 B.n110 VSUBS 0.006528f
C145 B.n111 VSUBS 0.006528f
C146 B.n112 VSUBS 0.006528f
C147 B.n113 VSUBS 0.006528f
C148 B.n114 VSUBS 0.006528f
C149 B.n115 VSUBS 0.006528f
C150 B.n116 VSUBS 0.006528f
C151 B.n117 VSUBS 0.006528f
C152 B.n118 VSUBS 0.006528f
C153 B.n119 VSUBS 0.006528f
C154 B.n120 VSUBS 0.006528f
C155 B.n121 VSUBS 0.006528f
C156 B.n122 VSUBS 0.006528f
C157 B.n123 VSUBS 0.006528f
C158 B.n124 VSUBS 0.006528f
C159 B.n125 VSUBS 0.006528f
C160 B.n126 VSUBS 0.006528f
C161 B.n127 VSUBS 0.006528f
C162 B.n128 VSUBS 0.006528f
C163 B.n129 VSUBS 0.006528f
C164 B.n130 VSUBS 0.015059f
C165 B.n131 VSUBS 0.006528f
C166 B.n132 VSUBS 0.006528f
C167 B.n133 VSUBS 0.006528f
C168 B.n134 VSUBS 0.006528f
C169 B.n135 VSUBS 0.006528f
C170 B.n136 VSUBS 0.006528f
C171 B.n137 VSUBS 0.006528f
C172 B.n138 VSUBS 0.006528f
C173 B.n139 VSUBS 0.006528f
C174 B.n140 VSUBS 0.006528f
C175 B.n141 VSUBS 0.006528f
C176 B.n142 VSUBS 0.006528f
C177 B.n143 VSUBS 0.006528f
C178 B.n144 VSUBS 0.006528f
C179 B.n145 VSUBS 0.006528f
C180 B.n146 VSUBS 0.006528f
C181 B.n147 VSUBS 0.006528f
C182 B.n148 VSUBS 0.006528f
C183 B.n149 VSUBS 0.006528f
C184 B.n150 VSUBS 0.006528f
C185 B.n151 VSUBS 0.006528f
C186 B.n152 VSUBS 0.006528f
C187 B.n153 VSUBS 0.006528f
C188 B.n154 VSUBS 0.006528f
C189 B.n155 VSUBS 0.006528f
C190 B.n156 VSUBS 0.006528f
C191 B.n157 VSUBS 0.006528f
C192 B.t7 VSUBS 0.513142f
C193 B.t8 VSUBS 0.529892f
C194 B.t6 VSUBS 1.38281f
C195 B.n158 VSUBS 0.262935f
C196 B.n159 VSUBS 0.065135f
C197 B.n160 VSUBS 0.015125f
C198 B.n161 VSUBS 0.006528f
C199 B.n162 VSUBS 0.006528f
C200 B.n163 VSUBS 0.006528f
C201 B.n164 VSUBS 0.006528f
C202 B.n165 VSUBS 0.006528f
C203 B.t10 VSUBS 0.513158f
C204 B.t11 VSUBS 0.529906f
C205 B.t9 VSUBS 1.38281f
C206 B.n166 VSUBS 0.262921f
C207 B.n167 VSUBS 0.065118f
C208 B.n168 VSUBS 0.006528f
C209 B.n169 VSUBS 0.006528f
C210 B.n170 VSUBS 0.006528f
C211 B.n171 VSUBS 0.006528f
C212 B.n172 VSUBS 0.006528f
C213 B.n173 VSUBS 0.006528f
C214 B.n174 VSUBS 0.006528f
C215 B.n175 VSUBS 0.006528f
C216 B.n176 VSUBS 0.006528f
C217 B.n177 VSUBS 0.006528f
C218 B.n178 VSUBS 0.006528f
C219 B.n179 VSUBS 0.006528f
C220 B.n180 VSUBS 0.006528f
C221 B.n181 VSUBS 0.006528f
C222 B.n182 VSUBS 0.006528f
C223 B.n183 VSUBS 0.006528f
C224 B.n184 VSUBS 0.006528f
C225 B.n185 VSUBS 0.006528f
C226 B.n186 VSUBS 0.006528f
C227 B.n187 VSUBS 0.006528f
C228 B.n188 VSUBS 0.006528f
C229 B.n189 VSUBS 0.006528f
C230 B.n190 VSUBS 0.006528f
C231 B.n191 VSUBS 0.006528f
C232 B.n192 VSUBS 0.006528f
C233 B.n193 VSUBS 0.006528f
C234 B.n194 VSUBS 0.016238f
C235 B.n195 VSUBS 0.006528f
C236 B.n196 VSUBS 0.006528f
C237 B.n197 VSUBS 0.006528f
C238 B.n198 VSUBS 0.006528f
C239 B.n199 VSUBS 0.006528f
C240 B.n200 VSUBS 0.006528f
C241 B.n201 VSUBS 0.006528f
C242 B.n202 VSUBS 0.006528f
C243 B.n203 VSUBS 0.006528f
C244 B.n204 VSUBS 0.006528f
C245 B.n205 VSUBS 0.006528f
C246 B.n206 VSUBS 0.006528f
C247 B.n207 VSUBS 0.006528f
C248 B.n208 VSUBS 0.006528f
C249 B.n209 VSUBS 0.006528f
C250 B.n210 VSUBS 0.006528f
C251 B.n211 VSUBS 0.006528f
C252 B.n212 VSUBS 0.006528f
C253 B.n213 VSUBS 0.006528f
C254 B.n214 VSUBS 0.006528f
C255 B.n215 VSUBS 0.006528f
C256 B.n216 VSUBS 0.006528f
C257 B.n217 VSUBS 0.006528f
C258 B.n218 VSUBS 0.006528f
C259 B.n219 VSUBS 0.006528f
C260 B.n220 VSUBS 0.006528f
C261 B.n221 VSUBS 0.006528f
C262 B.n222 VSUBS 0.006528f
C263 B.n223 VSUBS 0.006528f
C264 B.n224 VSUBS 0.006528f
C265 B.n225 VSUBS 0.006528f
C266 B.n226 VSUBS 0.006528f
C267 B.n227 VSUBS 0.006528f
C268 B.n228 VSUBS 0.006528f
C269 B.n229 VSUBS 0.006528f
C270 B.n230 VSUBS 0.006528f
C271 B.n231 VSUBS 0.006528f
C272 B.n232 VSUBS 0.006528f
C273 B.n233 VSUBS 0.006528f
C274 B.n234 VSUBS 0.006528f
C275 B.n235 VSUBS 0.006528f
C276 B.n236 VSUBS 0.006528f
C277 B.n237 VSUBS 0.006528f
C278 B.n238 VSUBS 0.006528f
C279 B.n239 VSUBS 0.006528f
C280 B.n240 VSUBS 0.006528f
C281 B.n241 VSUBS 0.006528f
C282 B.n242 VSUBS 0.006528f
C283 B.n243 VSUBS 0.006528f
C284 B.n244 VSUBS 0.006528f
C285 B.n245 VSUBS 0.006528f
C286 B.n246 VSUBS 0.006528f
C287 B.n247 VSUBS 0.006528f
C288 B.n248 VSUBS 0.006528f
C289 B.n249 VSUBS 0.006528f
C290 B.n250 VSUBS 0.006528f
C291 B.n251 VSUBS 0.006528f
C292 B.n252 VSUBS 0.006528f
C293 B.n253 VSUBS 0.006528f
C294 B.n254 VSUBS 0.006528f
C295 B.n255 VSUBS 0.006528f
C296 B.n256 VSUBS 0.006528f
C297 B.n257 VSUBS 0.006528f
C298 B.n258 VSUBS 0.006528f
C299 B.n259 VSUBS 0.006528f
C300 B.n260 VSUBS 0.006528f
C301 B.n261 VSUBS 0.006528f
C302 B.n262 VSUBS 0.006528f
C303 B.n263 VSUBS 0.006528f
C304 B.n264 VSUBS 0.006528f
C305 B.n265 VSUBS 0.006528f
C306 B.n266 VSUBS 0.006528f
C307 B.n267 VSUBS 0.006528f
C308 B.n268 VSUBS 0.006528f
C309 B.n269 VSUBS 0.006528f
C310 B.n270 VSUBS 0.006528f
C311 B.n271 VSUBS 0.006528f
C312 B.n272 VSUBS 0.006528f
C313 B.n273 VSUBS 0.006528f
C314 B.n274 VSUBS 0.006528f
C315 B.n275 VSUBS 0.006528f
C316 B.n276 VSUBS 0.006528f
C317 B.n277 VSUBS 0.015059f
C318 B.n278 VSUBS 0.015059f
C319 B.n279 VSUBS 0.016238f
C320 B.n280 VSUBS 0.006528f
C321 B.n281 VSUBS 0.006528f
C322 B.n282 VSUBS 0.006528f
C323 B.n283 VSUBS 0.006528f
C324 B.n284 VSUBS 0.006528f
C325 B.n285 VSUBS 0.006528f
C326 B.n286 VSUBS 0.006528f
C327 B.n287 VSUBS 0.006528f
C328 B.n288 VSUBS 0.006528f
C329 B.n289 VSUBS 0.006528f
C330 B.n290 VSUBS 0.006528f
C331 B.n291 VSUBS 0.006528f
C332 B.n292 VSUBS 0.006528f
C333 B.n293 VSUBS 0.006528f
C334 B.n294 VSUBS 0.006528f
C335 B.n295 VSUBS 0.006528f
C336 B.n296 VSUBS 0.006528f
C337 B.n297 VSUBS 0.006528f
C338 B.n298 VSUBS 0.006528f
C339 B.n299 VSUBS 0.006528f
C340 B.n300 VSUBS 0.006528f
C341 B.n301 VSUBS 0.006528f
C342 B.n302 VSUBS 0.006528f
C343 B.n303 VSUBS 0.006528f
C344 B.n304 VSUBS 0.006528f
C345 B.n305 VSUBS 0.006528f
C346 B.n306 VSUBS 0.006528f
C347 B.n307 VSUBS 0.006528f
C348 B.n308 VSUBS 0.006528f
C349 B.n309 VSUBS 0.006528f
C350 B.n310 VSUBS 0.006528f
C351 B.n311 VSUBS 0.006528f
C352 B.n312 VSUBS 0.006528f
C353 B.n313 VSUBS 0.006528f
C354 B.n314 VSUBS 0.006528f
C355 B.n315 VSUBS 0.006528f
C356 B.n316 VSUBS 0.006528f
C357 B.n317 VSUBS 0.006528f
C358 B.n318 VSUBS 0.006528f
C359 B.n319 VSUBS 0.006528f
C360 B.n320 VSUBS 0.006528f
C361 B.n321 VSUBS 0.006528f
C362 B.n322 VSUBS 0.006528f
C363 B.n323 VSUBS 0.006528f
C364 B.n324 VSUBS 0.006528f
C365 B.n325 VSUBS 0.006528f
C366 B.n326 VSUBS 0.006528f
C367 B.n327 VSUBS 0.006528f
C368 B.n328 VSUBS 0.006528f
C369 B.n329 VSUBS 0.006528f
C370 B.n330 VSUBS 0.006528f
C371 B.n331 VSUBS 0.006528f
C372 B.n332 VSUBS 0.006528f
C373 B.n333 VSUBS 0.006528f
C374 B.n334 VSUBS 0.006528f
C375 B.n335 VSUBS 0.006528f
C376 B.n336 VSUBS 0.006528f
C377 B.n337 VSUBS 0.006528f
C378 B.n338 VSUBS 0.006528f
C379 B.n339 VSUBS 0.006528f
C380 B.n340 VSUBS 0.006528f
C381 B.n341 VSUBS 0.006528f
C382 B.n342 VSUBS 0.006528f
C383 B.n343 VSUBS 0.006528f
C384 B.n344 VSUBS 0.006528f
C385 B.n345 VSUBS 0.006528f
C386 B.n346 VSUBS 0.006528f
C387 B.n347 VSUBS 0.006528f
C388 B.n348 VSUBS 0.006528f
C389 B.n349 VSUBS 0.006528f
C390 B.n350 VSUBS 0.006528f
C391 B.n351 VSUBS 0.006528f
C392 B.n352 VSUBS 0.006528f
C393 B.n353 VSUBS 0.006528f
C394 B.n354 VSUBS 0.006528f
C395 B.n355 VSUBS 0.006528f
C396 B.n356 VSUBS 0.006528f
C397 B.n357 VSUBS 0.006528f
C398 B.n358 VSUBS 0.006528f
C399 B.n359 VSUBS 0.006528f
C400 B.n360 VSUBS 0.004512f
C401 B.n361 VSUBS 0.015125f
C402 B.n362 VSUBS 0.00528f
C403 B.n363 VSUBS 0.006528f
C404 B.n364 VSUBS 0.006528f
C405 B.n365 VSUBS 0.006528f
C406 B.n366 VSUBS 0.006528f
C407 B.n367 VSUBS 0.006528f
C408 B.n368 VSUBS 0.006528f
C409 B.n369 VSUBS 0.006528f
C410 B.n370 VSUBS 0.006528f
C411 B.n371 VSUBS 0.006528f
C412 B.n372 VSUBS 0.006528f
C413 B.n373 VSUBS 0.006528f
C414 B.n374 VSUBS 0.00528f
C415 B.n375 VSUBS 0.006528f
C416 B.n376 VSUBS 0.006528f
C417 B.n377 VSUBS 0.004512f
C418 B.n378 VSUBS 0.006528f
C419 B.n379 VSUBS 0.006528f
C420 B.n380 VSUBS 0.006528f
C421 B.n381 VSUBS 0.006528f
C422 B.n382 VSUBS 0.006528f
C423 B.n383 VSUBS 0.006528f
C424 B.n384 VSUBS 0.006528f
C425 B.n385 VSUBS 0.006528f
C426 B.n386 VSUBS 0.006528f
C427 B.n387 VSUBS 0.006528f
C428 B.n388 VSUBS 0.006528f
C429 B.n389 VSUBS 0.006528f
C430 B.n390 VSUBS 0.006528f
C431 B.n391 VSUBS 0.006528f
C432 B.n392 VSUBS 0.006528f
C433 B.n393 VSUBS 0.006528f
C434 B.n394 VSUBS 0.006528f
C435 B.n395 VSUBS 0.006528f
C436 B.n396 VSUBS 0.006528f
C437 B.n397 VSUBS 0.006528f
C438 B.n398 VSUBS 0.006528f
C439 B.n399 VSUBS 0.006528f
C440 B.n400 VSUBS 0.006528f
C441 B.n401 VSUBS 0.006528f
C442 B.n402 VSUBS 0.006528f
C443 B.n403 VSUBS 0.006528f
C444 B.n404 VSUBS 0.006528f
C445 B.n405 VSUBS 0.006528f
C446 B.n406 VSUBS 0.006528f
C447 B.n407 VSUBS 0.006528f
C448 B.n408 VSUBS 0.006528f
C449 B.n409 VSUBS 0.006528f
C450 B.n410 VSUBS 0.006528f
C451 B.n411 VSUBS 0.006528f
C452 B.n412 VSUBS 0.006528f
C453 B.n413 VSUBS 0.006528f
C454 B.n414 VSUBS 0.006528f
C455 B.n415 VSUBS 0.006528f
C456 B.n416 VSUBS 0.006528f
C457 B.n417 VSUBS 0.006528f
C458 B.n418 VSUBS 0.006528f
C459 B.n419 VSUBS 0.006528f
C460 B.n420 VSUBS 0.006528f
C461 B.n421 VSUBS 0.006528f
C462 B.n422 VSUBS 0.006528f
C463 B.n423 VSUBS 0.006528f
C464 B.n424 VSUBS 0.006528f
C465 B.n425 VSUBS 0.006528f
C466 B.n426 VSUBS 0.006528f
C467 B.n427 VSUBS 0.006528f
C468 B.n428 VSUBS 0.006528f
C469 B.n429 VSUBS 0.006528f
C470 B.n430 VSUBS 0.006528f
C471 B.n431 VSUBS 0.006528f
C472 B.n432 VSUBS 0.006528f
C473 B.n433 VSUBS 0.006528f
C474 B.n434 VSUBS 0.006528f
C475 B.n435 VSUBS 0.006528f
C476 B.n436 VSUBS 0.006528f
C477 B.n437 VSUBS 0.006528f
C478 B.n438 VSUBS 0.006528f
C479 B.n439 VSUBS 0.006528f
C480 B.n440 VSUBS 0.006528f
C481 B.n441 VSUBS 0.006528f
C482 B.n442 VSUBS 0.006528f
C483 B.n443 VSUBS 0.006528f
C484 B.n444 VSUBS 0.006528f
C485 B.n445 VSUBS 0.006528f
C486 B.n446 VSUBS 0.006528f
C487 B.n447 VSUBS 0.006528f
C488 B.n448 VSUBS 0.006528f
C489 B.n449 VSUBS 0.006528f
C490 B.n450 VSUBS 0.006528f
C491 B.n451 VSUBS 0.006528f
C492 B.n452 VSUBS 0.006528f
C493 B.n453 VSUBS 0.006528f
C494 B.n454 VSUBS 0.006528f
C495 B.n455 VSUBS 0.006528f
C496 B.n456 VSUBS 0.006528f
C497 B.n457 VSUBS 0.016238f
C498 B.n458 VSUBS 0.016238f
C499 B.n459 VSUBS 0.015059f
C500 B.n460 VSUBS 0.006528f
C501 B.n461 VSUBS 0.006528f
C502 B.n462 VSUBS 0.006528f
C503 B.n463 VSUBS 0.006528f
C504 B.n464 VSUBS 0.006528f
C505 B.n465 VSUBS 0.006528f
C506 B.n466 VSUBS 0.006528f
C507 B.n467 VSUBS 0.006528f
C508 B.n468 VSUBS 0.006528f
C509 B.n469 VSUBS 0.006528f
C510 B.n470 VSUBS 0.006528f
C511 B.n471 VSUBS 0.006528f
C512 B.n472 VSUBS 0.006528f
C513 B.n473 VSUBS 0.006528f
C514 B.n474 VSUBS 0.006528f
C515 B.n475 VSUBS 0.006528f
C516 B.n476 VSUBS 0.006528f
C517 B.n477 VSUBS 0.006528f
C518 B.n478 VSUBS 0.006528f
C519 B.n479 VSUBS 0.006528f
C520 B.n480 VSUBS 0.006528f
C521 B.n481 VSUBS 0.006528f
C522 B.n482 VSUBS 0.006528f
C523 B.n483 VSUBS 0.006528f
C524 B.n484 VSUBS 0.006528f
C525 B.n485 VSUBS 0.006528f
C526 B.n486 VSUBS 0.006528f
C527 B.n487 VSUBS 0.006528f
C528 B.n488 VSUBS 0.006528f
C529 B.n489 VSUBS 0.006528f
C530 B.n490 VSUBS 0.006528f
C531 B.n491 VSUBS 0.006528f
C532 B.n492 VSUBS 0.006528f
C533 B.n493 VSUBS 0.006528f
C534 B.n494 VSUBS 0.006528f
C535 B.n495 VSUBS 0.006528f
C536 B.n496 VSUBS 0.006528f
C537 B.n497 VSUBS 0.006528f
C538 B.n498 VSUBS 0.006528f
C539 B.n499 VSUBS 0.006528f
C540 B.n500 VSUBS 0.006528f
C541 B.n501 VSUBS 0.006528f
C542 B.n502 VSUBS 0.006528f
C543 B.n503 VSUBS 0.006528f
C544 B.n504 VSUBS 0.006528f
C545 B.n505 VSUBS 0.006528f
C546 B.n506 VSUBS 0.006528f
C547 B.n507 VSUBS 0.006528f
C548 B.n508 VSUBS 0.006528f
C549 B.n509 VSUBS 0.006528f
C550 B.n510 VSUBS 0.006528f
C551 B.n511 VSUBS 0.006528f
C552 B.n512 VSUBS 0.006528f
C553 B.n513 VSUBS 0.006528f
C554 B.n514 VSUBS 0.006528f
C555 B.n515 VSUBS 0.006528f
C556 B.n516 VSUBS 0.006528f
C557 B.n517 VSUBS 0.006528f
C558 B.n518 VSUBS 0.006528f
C559 B.n519 VSUBS 0.006528f
C560 B.n520 VSUBS 0.006528f
C561 B.n521 VSUBS 0.006528f
C562 B.n522 VSUBS 0.006528f
C563 B.n523 VSUBS 0.006528f
C564 B.n524 VSUBS 0.006528f
C565 B.n525 VSUBS 0.006528f
C566 B.n526 VSUBS 0.006528f
C567 B.n527 VSUBS 0.006528f
C568 B.n528 VSUBS 0.006528f
C569 B.n529 VSUBS 0.006528f
C570 B.n530 VSUBS 0.006528f
C571 B.n531 VSUBS 0.006528f
C572 B.n532 VSUBS 0.006528f
C573 B.n533 VSUBS 0.006528f
C574 B.n534 VSUBS 0.006528f
C575 B.n535 VSUBS 0.006528f
C576 B.n536 VSUBS 0.006528f
C577 B.n537 VSUBS 0.006528f
C578 B.n538 VSUBS 0.006528f
C579 B.n539 VSUBS 0.006528f
C580 B.n540 VSUBS 0.006528f
C581 B.n541 VSUBS 0.006528f
C582 B.n542 VSUBS 0.006528f
C583 B.n543 VSUBS 0.006528f
C584 B.n544 VSUBS 0.006528f
C585 B.n545 VSUBS 0.006528f
C586 B.n546 VSUBS 0.006528f
C587 B.n547 VSUBS 0.006528f
C588 B.n548 VSUBS 0.006528f
C589 B.n549 VSUBS 0.006528f
C590 B.n550 VSUBS 0.006528f
C591 B.n551 VSUBS 0.006528f
C592 B.n552 VSUBS 0.006528f
C593 B.n553 VSUBS 0.006528f
C594 B.n554 VSUBS 0.006528f
C595 B.n555 VSUBS 0.006528f
C596 B.n556 VSUBS 0.006528f
C597 B.n557 VSUBS 0.006528f
C598 B.n558 VSUBS 0.006528f
C599 B.n559 VSUBS 0.006528f
C600 B.n560 VSUBS 0.006528f
C601 B.n561 VSUBS 0.006528f
C602 B.n562 VSUBS 0.006528f
C603 B.n563 VSUBS 0.006528f
C604 B.n564 VSUBS 0.006528f
C605 B.n565 VSUBS 0.006528f
C606 B.n566 VSUBS 0.006528f
C607 B.n567 VSUBS 0.006528f
C608 B.n568 VSUBS 0.006528f
C609 B.n569 VSUBS 0.006528f
C610 B.n570 VSUBS 0.006528f
C611 B.n571 VSUBS 0.006528f
C612 B.n572 VSUBS 0.006528f
C613 B.n573 VSUBS 0.006528f
C614 B.n574 VSUBS 0.006528f
C615 B.n575 VSUBS 0.006528f
C616 B.n576 VSUBS 0.006528f
C617 B.n577 VSUBS 0.006528f
C618 B.n578 VSUBS 0.006528f
C619 B.n579 VSUBS 0.006528f
C620 B.n580 VSUBS 0.006528f
C621 B.n581 VSUBS 0.006528f
C622 B.n582 VSUBS 0.006528f
C623 B.n583 VSUBS 0.006528f
C624 B.n584 VSUBS 0.006528f
C625 B.n585 VSUBS 0.006528f
C626 B.n586 VSUBS 0.006528f
C627 B.n587 VSUBS 0.006528f
C628 B.n588 VSUBS 0.015803f
C629 B.n589 VSUBS 0.015494f
C630 B.n590 VSUBS 0.016238f
C631 B.n591 VSUBS 0.006528f
C632 B.n592 VSUBS 0.006528f
C633 B.n593 VSUBS 0.006528f
C634 B.n594 VSUBS 0.006528f
C635 B.n595 VSUBS 0.006528f
C636 B.n596 VSUBS 0.006528f
C637 B.n597 VSUBS 0.006528f
C638 B.n598 VSUBS 0.006528f
C639 B.n599 VSUBS 0.006528f
C640 B.n600 VSUBS 0.006528f
C641 B.n601 VSUBS 0.006528f
C642 B.n602 VSUBS 0.006528f
C643 B.n603 VSUBS 0.006528f
C644 B.n604 VSUBS 0.006528f
C645 B.n605 VSUBS 0.006528f
C646 B.n606 VSUBS 0.006528f
C647 B.n607 VSUBS 0.006528f
C648 B.n608 VSUBS 0.006528f
C649 B.n609 VSUBS 0.006528f
C650 B.n610 VSUBS 0.006528f
C651 B.n611 VSUBS 0.006528f
C652 B.n612 VSUBS 0.006528f
C653 B.n613 VSUBS 0.006528f
C654 B.n614 VSUBS 0.006528f
C655 B.n615 VSUBS 0.006528f
C656 B.n616 VSUBS 0.006528f
C657 B.n617 VSUBS 0.006528f
C658 B.n618 VSUBS 0.006528f
C659 B.n619 VSUBS 0.006528f
C660 B.n620 VSUBS 0.006528f
C661 B.n621 VSUBS 0.006528f
C662 B.n622 VSUBS 0.006528f
C663 B.n623 VSUBS 0.006528f
C664 B.n624 VSUBS 0.006528f
C665 B.n625 VSUBS 0.006528f
C666 B.n626 VSUBS 0.006528f
C667 B.n627 VSUBS 0.006528f
C668 B.n628 VSUBS 0.006528f
C669 B.n629 VSUBS 0.006528f
C670 B.n630 VSUBS 0.006528f
C671 B.n631 VSUBS 0.006528f
C672 B.n632 VSUBS 0.006528f
C673 B.n633 VSUBS 0.006528f
C674 B.n634 VSUBS 0.006528f
C675 B.n635 VSUBS 0.006528f
C676 B.n636 VSUBS 0.006528f
C677 B.n637 VSUBS 0.006528f
C678 B.n638 VSUBS 0.006528f
C679 B.n639 VSUBS 0.006528f
C680 B.n640 VSUBS 0.006528f
C681 B.n641 VSUBS 0.006528f
C682 B.n642 VSUBS 0.006528f
C683 B.n643 VSUBS 0.006528f
C684 B.n644 VSUBS 0.006528f
C685 B.n645 VSUBS 0.006528f
C686 B.n646 VSUBS 0.006528f
C687 B.n647 VSUBS 0.006528f
C688 B.n648 VSUBS 0.006528f
C689 B.n649 VSUBS 0.006528f
C690 B.n650 VSUBS 0.006528f
C691 B.n651 VSUBS 0.006528f
C692 B.n652 VSUBS 0.006528f
C693 B.n653 VSUBS 0.006528f
C694 B.n654 VSUBS 0.006528f
C695 B.n655 VSUBS 0.006528f
C696 B.n656 VSUBS 0.006528f
C697 B.n657 VSUBS 0.006528f
C698 B.n658 VSUBS 0.006528f
C699 B.n659 VSUBS 0.006528f
C700 B.n660 VSUBS 0.006528f
C701 B.n661 VSUBS 0.006528f
C702 B.n662 VSUBS 0.006528f
C703 B.n663 VSUBS 0.006528f
C704 B.n664 VSUBS 0.006528f
C705 B.n665 VSUBS 0.006528f
C706 B.n666 VSUBS 0.006528f
C707 B.n667 VSUBS 0.006528f
C708 B.n668 VSUBS 0.006528f
C709 B.n669 VSUBS 0.006528f
C710 B.n670 VSUBS 0.006528f
C711 B.n671 VSUBS 0.004512f
C712 B.n672 VSUBS 0.015125f
C713 B.n673 VSUBS 0.00528f
C714 B.n674 VSUBS 0.006528f
C715 B.n675 VSUBS 0.006528f
C716 B.n676 VSUBS 0.006528f
C717 B.n677 VSUBS 0.006528f
C718 B.n678 VSUBS 0.006528f
C719 B.n679 VSUBS 0.006528f
C720 B.n680 VSUBS 0.006528f
C721 B.n681 VSUBS 0.006528f
C722 B.n682 VSUBS 0.006528f
C723 B.n683 VSUBS 0.006528f
C724 B.n684 VSUBS 0.006528f
C725 B.n685 VSUBS 0.00528f
C726 B.n686 VSUBS 0.015125f
C727 B.n687 VSUBS 0.004512f
C728 B.n688 VSUBS 0.006528f
C729 B.n689 VSUBS 0.006528f
C730 B.n690 VSUBS 0.006528f
C731 B.n691 VSUBS 0.006528f
C732 B.n692 VSUBS 0.006528f
C733 B.n693 VSUBS 0.006528f
C734 B.n694 VSUBS 0.006528f
C735 B.n695 VSUBS 0.006528f
C736 B.n696 VSUBS 0.006528f
C737 B.n697 VSUBS 0.006528f
C738 B.n698 VSUBS 0.006528f
C739 B.n699 VSUBS 0.006528f
C740 B.n700 VSUBS 0.006528f
C741 B.n701 VSUBS 0.006528f
C742 B.n702 VSUBS 0.006528f
C743 B.n703 VSUBS 0.006528f
C744 B.n704 VSUBS 0.006528f
C745 B.n705 VSUBS 0.006528f
C746 B.n706 VSUBS 0.006528f
C747 B.n707 VSUBS 0.006528f
C748 B.n708 VSUBS 0.006528f
C749 B.n709 VSUBS 0.006528f
C750 B.n710 VSUBS 0.006528f
C751 B.n711 VSUBS 0.006528f
C752 B.n712 VSUBS 0.006528f
C753 B.n713 VSUBS 0.006528f
C754 B.n714 VSUBS 0.006528f
C755 B.n715 VSUBS 0.006528f
C756 B.n716 VSUBS 0.006528f
C757 B.n717 VSUBS 0.006528f
C758 B.n718 VSUBS 0.006528f
C759 B.n719 VSUBS 0.006528f
C760 B.n720 VSUBS 0.006528f
C761 B.n721 VSUBS 0.006528f
C762 B.n722 VSUBS 0.006528f
C763 B.n723 VSUBS 0.006528f
C764 B.n724 VSUBS 0.006528f
C765 B.n725 VSUBS 0.006528f
C766 B.n726 VSUBS 0.006528f
C767 B.n727 VSUBS 0.006528f
C768 B.n728 VSUBS 0.006528f
C769 B.n729 VSUBS 0.006528f
C770 B.n730 VSUBS 0.006528f
C771 B.n731 VSUBS 0.006528f
C772 B.n732 VSUBS 0.006528f
C773 B.n733 VSUBS 0.006528f
C774 B.n734 VSUBS 0.006528f
C775 B.n735 VSUBS 0.006528f
C776 B.n736 VSUBS 0.006528f
C777 B.n737 VSUBS 0.006528f
C778 B.n738 VSUBS 0.006528f
C779 B.n739 VSUBS 0.006528f
C780 B.n740 VSUBS 0.006528f
C781 B.n741 VSUBS 0.006528f
C782 B.n742 VSUBS 0.006528f
C783 B.n743 VSUBS 0.006528f
C784 B.n744 VSUBS 0.006528f
C785 B.n745 VSUBS 0.006528f
C786 B.n746 VSUBS 0.006528f
C787 B.n747 VSUBS 0.006528f
C788 B.n748 VSUBS 0.006528f
C789 B.n749 VSUBS 0.006528f
C790 B.n750 VSUBS 0.006528f
C791 B.n751 VSUBS 0.006528f
C792 B.n752 VSUBS 0.006528f
C793 B.n753 VSUBS 0.006528f
C794 B.n754 VSUBS 0.006528f
C795 B.n755 VSUBS 0.006528f
C796 B.n756 VSUBS 0.006528f
C797 B.n757 VSUBS 0.006528f
C798 B.n758 VSUBS 0.006528f
C799 B.n759 VSUBS 0.006528f
C800 B.n760 VSUBS 0.006528f
C801 B.n761 VSUBS 0.006528f
C802 B.n762 VSUBS 0.006528f
C803 B.n763 VSUBS 0.006528f
C804 B.n764 VSUBS 0.006528f
C805 B.n765 VSUBS 0.006528f
C806 B.n766 VSUBS 0.006528f
C807 B.n767 VSUBS 0.006528f
C808 B.n768 VSUBS 0.016238f
C809 B.n769 VSUBS 0.016238f
C810 B.n770 VSUBS 0.015059f
C811 B.n771 VSUBS 0.006528f
C812 B.n772 VSUBS 0.006528f
C813 B.n773 VSUBS 0.006528f
C814 B.n774 VSUBS 0.006528f
C815 B.n775 VSUBS 0.006528f
C816 B.n776 VSUBS 0.006528f
C817 B.n777 VSUBS 0.006528f
C818 B.n778 VSUBS 0.006528f
C819 B.n779 VSUBS 0.006528f
C820 B.n780 VSUBS 0.006528f
C821 B.n781 VSUBS 0.006528f
C822 B.n782 VSUBS 0.006528f
C823 B.n783 VSUBS 0.006528f
C824 B.n784 VSUBS 0.006528f
C825 B.n785 VSUBS 0.006528f
C826 B.n786 VSUBS 0.006528f
C827 B.n787 VSUBS 0.006528f
C828 B.n788 VSUBS 0.006528f
C829 B.n789 VSUBS 0.006528f
C830 B.n790 VSUBS 0.006528f
C831 B.n791 VSUBS 0.006528f
C832 B.n792 VSUBS 0.006528f
C833 B.n793 VSUBS 0.006528f
C834 B.n794 VSUBS 0.006528f
C835 B.n795 VSUBS 0.006528f
C836 B.n796 VSUBS 0.006528f
C837 B.n797 VSUBS 0.006528f
C838 B.n798 VSUBS 0.006528f
C839 B.n799 VSUBS 0.006528f
C840 B.n800 VSUBS 0.006528f
C841 B.n801 VSUBS 0.006528f
C842 B.n802 VSUBS 0.006528f
C843 B.n803 VSUBS 0.006528f
C844 B.n804 VSUBS 0.006528f
C845 B.n805 VSUBS 0.006528f
C846 B.n806 VSUBS 0.006528f
C847 B.n807 VSUBS 0.006528f
C848 B.n808 VSUBS 0.006528f
C849 B.n809 VSUBS 0.006528f
C850 B.n810 VSUBS 0.006528f
C851 B.n811 VSUBS 0.006528f
C852 B.n812 VSUBS 0.006528f
C853 B.n813 VSUBS 0.006528f
C854 B.n814 VSUBS 0.006528f
C855 B.n815 VSUBS 0.006528f
C856 B.n816 VSUBS 0.006528f
C857 B.n817 VSUBS 0.006528f
C858 B.n818 VSUBS 0.006528f
C859 B.n819 VSUBS 0.006528f
C860 B.n820 VSUBS 0.006528f
C861 B.n821 VSUBS 0.006528f
C862 B.n822 VSUBS 0.006528f
C863 B.n823 VSUBS 0.006528f
C864 B.n824 VSUBS 0.006528f
C865 B.n825 VSUBS 0.006528f
C866 B.n826 VSUBS 0.006528f
C867 B.n827 VSUBS 0.006528f
C868 B.n828 VSUBS 0.006528f
C869 B.n829 VSUBS 0.006528f
C870 B.n830 VSUBS 0.006528f
C871 B.n831 VSUBS 0.006528f
C872 B.n832 VSUBS 0.006528f
C873 B.n833 VSUBS 0.006528f
C874 B.n834 VSUBS 0.006528f
C875 B.n835 VSUBS 0.014782f
C876 VDD1.t7 VSUBS 0.320623f
C877 VDD1.t3 VSUBS 0.320623f
C878 VDD1.n0 VSUBS 2.64124f
C879 VDD1.t1 VSUBS 0.320623f
C880 VDD1.t5 VSUBS 0.320623f
C881 VDD1.n1 VSUBS 2.63993f
C882 VDD1.t2 VSUBS 0.320623f
C883 VDD1.t6 VSUBS 0.320623f
C884 VDD1.n2 VSUBS 2.63993f
C885 VDD1.n3 VSUBS 3.81179f
C886 VDD1.t4 VSUBS 0.320623f
C887 VDD1.t0 VSUBS 0.320623f
C888 VDD1.n4 VSUBS 2.62967f
C889 VDD1.n5 VSUBS 3.37504f
C890 VP.n0 VSUBS 0.041048f
C891 VP.t1 VSUBS 2.88966f
C892 VP.n1 VSUBS 0.034003f
C893 VP.n2 VSUBS 0.031135f
C894 VP.t5 VSUBS 2.88966f
C895 VP.n3 VSUBS 0.045451f
C896 VP.n4 VSUBS 0.031135f
C897 VP.t2 VSUBS 2.88966f
C898 VP.n5 VSUBS 0.060353f
C899 VP.n6 VSUBS 0.031135f
C900 VP.t6 VSUBS 2.88966f
C901 VP.n7 VSUBS 1.10388f
C902 VP.n8 VSUBS 0.041048f
C903 VP.t7 VSUBS 2.88966f
C904 VP.n9 VSUBS 0.034003f
C905 VP.n10 VSUBS 0.031135f
C906 VP.t3 VSUBS 2.88966f
C907 VP.n11 VSUBS 0.045451f
C908 VP.n12 VSUBS 0.26096f
C909 VP.t4 VSUBS 2.88966f
C910 VP.t0 VSUBS 3.0637f
C911 VP.n13 VSUBS 1.08199f
C912 VP.n14 VSUBS 1.10024f
C913 VP.n15 VSUBS 0.054874f
C914 VP.n16 VSUBS 0.045451f
C915 VP.n17 VSUBS 0.031135f
C916 VP.n18 VSUBS 0.031135f
C917 VP.n19 VSUBS 0.031135f
C918 VP.n20 VSUBS 0.054874f
C919 VP.n21 VSUBS 1.01184f
C920 VP.n22 VSUBS 0.032529f
C921 VP.n23 VSUBS 0.060353f
C922 VP.n24 VSUBS 0.031135f
C923 VP.n25 VSUBS 0.031135f
C924 VP.n26 VSUBS 0.031135f
C925 VP.n27 VSUBS 0.054573f
C926 VP.n28 VSUBS 0.048572f
C927 VP.n29 VSUBS 1.10388f
C928 VP.n30 VSUBS 1.80792f
C929 VP.n31 VSUBS 1.82957f
C930 VP.n32 VSUBS 0.041048f
C931 VP.n33 VSUBS 0.048572f
C932 VP.n34 VSUBS 0.054573f
C933 VP.n35 VSUBS 0.034003f
C934 VP.n36 VSUBS 0.031135f
C935 VP.n37 VSUBS 0.031135f
C936 VP.n38 VSUBS 0.031135f
C937 VP.n39 VSUBS 0.032529f
C938 VP.n40 VSUBS 1.01184f
C939 VP.n41 VSUBS 0.054874f
C940 VP.n42 VSUBS 0.045451f
C941 VP.n43 VSUBS 0.031135f
C942 VP.n44 VSUBS 0.031135f
C943 VP.n45 VSUBS 0.031135f
C944 VP.n46 VSUBS 0.054874f
C945 VP.n47 VSUBS 1.01184f
C946 VP.n48 VSUBS 0.032529f
C947 VP.n49 VSUBS 0.060353f
C948 VP.n50 VSUBS 0.031135f
C949 VP.n51 VSUBS 0.031135f
C950 VP.n52 VSUBS 0.031135f
C951 VP.n53 VSUBS 0.054573f
C952 VP.n54 VSUBS 0.048572f
C953 VP.n55 VSUBS 1.10388f
C954 VP.n56 VSUBS 0.041036f
C955 VTAIL.t8 VSUBS 0.306227f
C956 VTAIL.t9 VSUBS 0.306227f
C957 VTAIL.n0 VSUBS 2.3657f
C958 VTAIL.n1 VSUBS 0.737296f
C959 VTAIL.t12 VSUBS 3.09529f
C960 VTAIL.n2 VSUBS 0.87419f
C961 VTAIL.t4 VSUBS 3.09529f
C962 VTAIL.n3 VSUBS 0.87419f
C963 VTAIL.t1 VSUBS 0.306227f
C964 VTAIL.t2 VSUBS 0.306227f
C965 VTAIL.n4 VSUBS 2.3657f
C966 VTAIL.n5 VSUBS 0.889643f
C967 VTAIL.t6 VSUBS 3.09529f
C968 VTAIL.n6 VSUBS 2.39243f
C969 VTAIL.t13 VSUBS 3.0953f
C970 VTAIL.n7 VSUBS 2.39242f
C971 VTAIL.t10 VSUBS 0.306227f
C972 VTAIL.t15 VSUBS 0.306227f
C973 VTAIL.n8 VSUBS 2.3657f
C974 VTAIL.n9 VSUBS 0.889638f
C975 VTAIL.t11 VSUBS 3.0953f
C976 VTAIL.n10 VSUBS 0.874184f
C977 VTAIL.t0 VSUBS 3.0953f
C978 VTAIL.n11 VSUBS 0.874184f
C979 VTAIL.t3 VSUBS 0.306227f
C980 VTAIL.t5 VSUBS 0.306227f
C981 VTAIL.n12 VSUBS 2.3657f
C982 VTAIL.n13 VSUBS 0.889638f
C983 VTAIL.t7 VSUBS 3.09529f
C984 VTAIL.n14 VSUBS 2.39243f
C985 VTAIL.t14 VSUBS 3.09529f
C986 VTAIL.n15 VSUBS 2.388f
C987 VDD2.t0 VSUBS 0.317453f
C988 VDD2.t6 VSUBS 0.317453f
C989 VDD2.n0 VSUBS 2.61383f
C990 VDD2.t7 VSUBS 0.317453f
C991 VDD2.t4 VSUBS 0.317453f
C992 VDD2.n1 VSUBS 2.61383f
C993 VDD2.n2 VSUBS 3.723f
C994 VDD2.t1 VSUBS 0.317453f
C995 VDD2.t2 VSUBS 0.317453f
C996 VDD2.n3 VSUBS 2.60368f
C997 VDD2.n4 VSUBS 3.31153f
C998 VDD2.t5 VSUBS 0.317453f
C999 VDD2.t3 VSUBS 0.317453f
C1000 VDD2.n5 VSUBS 2.61379f
C1001 VN.n0 VSUBS 0.040237f
C1002 VN.t1 VSUBS 2.83257f
C1003 VN.n1 VSUBS 0.033331f
C1004 VN.n2 VSUBS 0.030519f
C1005 VN.t6 VSUBS 2.83257f
C1006 VN.n3 VSUBS 0.044553f
C1007 VN.n4 VSUBS 0.255804f
C1008 VN.t7 VSUBS 2.83257f
C1009 VN.t3 VSUBS 3.00317f
C1010 VN.n5 VSUBS 1.06061f
C1011 VN.n6 VSUBS 1.0785f
C1012 VN.n7 VSUBS 0.05379f
C1013 VN.n8 VSUBS 0.044553f
C1014 VN.n9 VSUBS 0.030519f
C1015 VN.n10 VSUBS 0.030519f
C1016 VN.n11 VSUBS 0.030519f
C1017 VN.n12 VSUBS 0.05379f
C1018 VN.n13 VSUBS 0.991845f
C1019 VN.n14 VSUBS 0.031886f
C1020 VN.n15 VSUBS 0.059161f
C1021 VN.n16 VSUBS 0.030519f
C1022 VN.n17 VSUBS 0.030519f
C1023 VN.n18 VSUBS 0.030519f
C1024 VN.n19 VSUBS 0.053494f
C1025 VN.n20 VSUBS 0.047612f
C1026 VN.n21 VSUBS 1.08207f
C1027 VN.n22 VSUBS 0.040225f
C1028 VN.n23 VSUBS 0.040237f
C1029 VN.t2 VSUBS 2.83257f
C1030 VN.n24 VSUBS 0.033331f
C1031 VN.n25 VSUBS 0.030519f
C1032 VN.t5 VSUBS 2.83257f
C1033 VN.n26 VSUBS 0.044553f
C1034 VN.n27 VSUBS 0.255804f
C1035 VN.t0 VSUBS 2.83257f
C1036 VN.t4 VSUBS 3.00317f
C1037 VN.n28 VSUBS 1.06061f
C1038 VN.n29 VSUBS 1.0785f
C1039 VN.n30 VSUBS 0.05379f
C1040 VN.n31 VSUBS 0.044553f
C1041 VN.n32 VSUBS 0.030519f
C1042 VN.n33 VSUBS 0.030519f
C1043 VN.n34 VSUBS 0.030519f
C1044 VN.n35 VSUBS 0.05379f
C1045 VN.n36 VSUBS 0.991845f
C1046 VN.n37 VSUBS 0.031886f
C1047 VN.n38 VSUBS 0.059161f
C1048 VN.n39 VSUBS 0.030519f
C1049 VN.n40 VSUBS 0.030519f
C1050 VN.n41 VSUBS 0.030519f
C1051 VN.n42 VSUBS 0.053494f
C1052 VN.n43 VSUBS 0.047612f
C1053 VN.n44 VSUBS 1.08207f
C1054 VN.n45 VSUBS 1.78852f
.ends

