* NGSPICE file created from diff_pair_sample_1367.ext - technology: sky130A

.subckt diff_pair_sample_1367 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=2.6235 ps=16.23 w=15.9 l=1.69
X1 B.t11 B.t9 B.t10 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=0 ps=0 w=15.9 l=1.69
X2 VTAIL.t6 VP.t1 VDD1.t1 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=2.6235 ps=16.23 w=15.9 l=1.69
X3 VDD2.t3 VN.t0 VTAIL.t3 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=2.6235 pd=16.23 as=6.201 ps=32.58 w=15.9 l=1.69
X4 B.t8 B.t6 B.t7 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=0 ps=0 w=15.9 l=1.69
X5 VDD1.t0 VP.t2 VTAIL.t5 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=2.6235 pd=16.23 as=6.201 ps=32.58 w=15.9 l=1.69
X6 B.t5 B.t3 B.t4 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=0 ps=0 w=15.9 l=1.69
X7 VTAIL.t1 VN.t1 VDD2.t2 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=2.6235 ps=16.23 w=15.9 l=1.69
X8 B.t2 B.t0 B.t1 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=0 ps=0 w=15.9 l=1.69
X9 VDD1.t3 VP.t3 VTAIL.t4 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=2.6235 pd=16.23 as=6.201 ps=32.58 w=15.9 l=1.69
X10 VTAIL.t2 VN.t2 VDD2.t1 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=6.201 pd=32.58 as=2.6235 ps=16.23 w=15.9 l=1.69
X11 VDD2.t0 VN.t3 VTAIL.t0 w_n2182_n4148# sky130_fd_pr__pfet_01v8 ad=2.6235 pd=16.23 as=6.201 ps=32.58 w=15.9 l=1.69
R0 VP.n3 VP.t0 261.692
R1 VP.n3 VP.t2 261.271
R2 VP.n5 VP.t1 226.74
R3 VP.n13 VP.t3 226.74
R4 VP.n5 VP.n4 185.4
R5 VP.n14 VP.n13 185.4
R6 VP.n12 VP.n0 161.3
R7 VP.n11 VP.n10 161.3
R8 VP.n9 VP.n1 161.3
R9 VP.n8 VP.n7 161.3
R10 VP.n6 VP.n2 161.3
R11 VP.n4 VP.n3 55.8727
R12 VP.n7 VP.n1 40.577
R13 VP.n11 VP.n1 40.577
R14 VP.n7 VP.n6 24.5923
R15 VP.n12 VP.n11 24.5923
R16 VP.n6 VP.n5 0.492337
R17 VP.n13 VP.n12 0.492337
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VDD1 VDD1.n1 116.686
R26 VDD1 VDD1.n0 73.5727
R27 VDD1.n0 VDD1.t2 2.04484
R28 VDD1.n0 VDD1.t0 2.04484
R29 VDD1.n1 VDD1.t1 2.04484
R30 VDD1.n1 VDD1.t3 2.04484
R31 VTAIL.n5 VTAIL.t7 58.8802
R32 VTAIL.n4 VTAIL.t3 58.8802
R33 VTAIL.n3 VTAIL.t2 58.8802
R34 VTAIL.n6 VTAIL.t5 58.88
R35 VTAIL.n7 VTAIL.t0 58.88
R36 VTAIL.n0 VTAIL.t1 58.88
R37 VTAIL.n1 VTAIL.t4 58.88
R38 VTAIL.n2 VTAIL.t6 58.88
R39 VTAIL.n7 VTAIL.n6 27.8152
R40 VTAIL.n3 VTAIL.n2 27.8152
R41 VTAIL.n4 VTAIL.n3 1.74188
R42 VTAIL.n6 VTAIL.n5 1.74188
R43 VTAIL.n2 VTAIL.n1 1.74188
R44 VTAIL VTAIL.n0 0.929379
R45 VTAIL VTAIL.n7 0.813
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 B.n473 B.n472 585
R49 B.n474 B.n77 585
R50 B.n476 B.n475 585
R51 B.n477 B.n76 585
R52 B.n479 B.n478 585
R53 B.n480 B.n75 585
R54 B.n482 B.n481 585
R55 B.n483 B.n74 585
R56 B.n485 B.n484 585
R57 B.n486 B.n73 585
R58 B.n488 B.n487 585
R59 B.n489 B.n72 585
R60 B.n491 B.n490 585
R61 B.n492 B.n71 585
R62 B.n494 B.n493 585
R63 B.n495 B.n70 585
R64 B.n497 B.n496 585
R65 B.n498 B.n69 585
R66 B.n500 B.n499 585
R67 B.n501 B.n68 585
R68 B.n503 B.n502 585
R69 B.n504 B.n67 585
R70 B.n506 B.n505 585
R71 B.n507 B.n66 585
R72 B.n509 B.n508 585
R73 B.n510 B.n65 585
R74 B.n512 B.n511 585
R75 B.n513 B.n64 585
R76 B.n515 B.n514 585
R77 B.n516 B.n63 585
R78 B.n518 B.n517 585
R79 B.n519 B.n62 585
R80 B.n521 B.n520 585
R81 B.n522 B.n61 585
R82 B.n524 B.n523 585
R83 B.n525 B.n60 585
R84 B.n527 B.n526 585
R85 B.n528 B.n59 585
R86 B.n530 B.n529 585
R87 B.n531 B.n58 585
R88 B.n533 B.n532 585
R89 B.n534 B.n57 585
R90 B.n536 B.n535 585
R91 B.n537 B.n56 585
R92 B.n539 B.n538 585
R93 B.n540 B.n55 585
R94 B.n542 B.n541 585
R95 B.n543 B.n54 585
R96 B.n545 B.n544 585
R97 B.n546 B.n53 585
R98 B.n548 B.n547 585
R99 B.n549 B.n49 585
R100 B.n551 B.n550 585
R101 B.n552 B.n48 585
R102 B.n554 B.n553 585
R103 B.n555 B.n47 585
R104 B.n557 B.n556 585
R105 B.n558 B.n46 585
R106 B.n560 B.n559 585
R107 B.n561 B.n45 585
R108 B.n563 B.n562 585
R109 B.n564 B.n44 585
R110 B.n566 B.n565 585
R111 B.n568 B.n41 585
R112 B.n570 B.n569 585
R113 B.n571 B.n40 585
R114 B.n573 B.n572 585
R115 B.n574 B.n39 585
R116 B.n576 B.n575 585
R117 B.n577 B.n38 585
R118 B.n579 B.n578 585
R119 B.n580 B.n37 585
R120 B.n582 B.n581 585
R121 B.n583 B.n36 585
R122 B.n585 B.n584 585
R123 B.n586 B.n35 585
R124 B.n588 B.n587 585
R125 B.n589 B.n34 585
R126 B.n591 B.n590 585
R127 B.n592 B.n33 585
R128 B.n594 B.n593 585
R129 B.n595 B.n32 585
R130 B.n597 B.n596 585
R131 B.n598 B.n31 585
R132 B.n600 B.n599 585
R133 B.n601 B.n30 585
R134 B.n603 B.n602 585
R135 B.n604 B.n29 585
R136 B.n606 B.n605 585
R137 B.n607 B.n28 585
R138 B.n609 B.n608 585
R139 B.n610 B.n27 585
R140 B.n612 B.n611 585
R141 B.n613 B.n26 585
R142 B.n615 B.n614 585
R143 B.n616 B.n25 585
R144 B.n618 B.n617 585
R145 B.n619 B.n24 585
R146 B.n621 B.n620 585
R147 B.n622 B.n23 585
R148 B.n624 B.n623 585
R149 B.n625 B.n22 585
R150 B.n627 B.n626 585
R151 B.n628 B.n21 585
R152 B.n630 B.n629 585
R153 B.n631 B.n20 585
R154 B.n633 B.n632 585
R155 B.n634 B.n19 585
R156 B.n636 B.n635 585
R157 B.n637 B.n18 585
R158 B.n639 B.n638 585
R159 B.n640 B.n17 585
R160 B.n642 B.n641 585
R161 B.n643 B.n16 585
R162 B.n645 B.n644 585
R163 B.n646 B.n15 585
R164 B.n471 B.n78 585
R165 B.n470 B.n469 585
R166 B.n468 B.n79 585
R167 B.n467 B.n466 585
R168 B.n465 B.n80 585
R169 B.n464 B.n463 585
R170 B.n462 B.n81 585
R171 B.n461 B.n460 585
R172 B.n459 B.n82 585
R173 B.n458 B.n457 585
R174 B.n456 B.n83 585
R175 B.n455 B.n454 585
R176 B.n453 B.n84 585
R177 B.n452 B.n451 585
R178 B.n450 B.n85 585
R179 B.n449 B.n448 585
R180 B.n447 B.n86 585
R181 B.n446 B.n445 585
R182 B.n444 B.n87 585
R183 B.n443 B.n442 585
R184 B.n441 B.n88 585
R185 B.n440 B.n439 585
R186 B.n438 B.n89 585
R187 B.n437 B.n436 585
R188 B.n435 B.n90 585
R189 B.n434 B.n433 585
R190 B.n432 B.n91 585
R191 B.n431 B.n430 585
R192 B.n429 B.n92 585
R193 B.n428 B.n427 585
R194 B.n426 B.n93 585
R195 B.n425 B.n424 585
R196 B.n423 B.n94 585
R197 B.n422 B.n421 585
R198 B.n420 B.n95 585
R199 B.n419 B.n418 585
R200 B.n417 B.n96 585
R201 B.n416 B.n415 585
R202 B.n414 B.n97 585
R203 B.n413 B.n412 585
R204 B.n411 B.n98 585
R205 B.n410 B.n409 585
R206 B.n408 B.n99 585
R207 B.n407 B.n406 585
R208 B.n405 B.n100 585
R209 B.n404 B.n403 585
R210 B.n402 B.n101 585
R211 B.n401 B.n400 585
R212 B.n399 B.n102 585
R213 B.n398 B.n397 585
R214 B.n396 B.n103 585
R215 B.n395 B.n394 585
R216 B.n393 B.n104 585
R217 B.n218 B.n217 585
R218 B.n219 B.n166 585
R219 B.n221 B.n220 585
R220 B.n222 B.n165 585
R221 B.n224 B.n223 585
R222 B.n225 B.n164 585
R223 B.n227 B.n226 585
R224 B.n228 B.n163 585
R225 B.n230 B.n229 585
R226 B.n231 B.n162 585
R227 B.n233 B.n232 585
R228 B.n234 B.n161 585
R229 B.n236 B.n235 585
R230 B.n237 B.n160 585
R231 B.n239 B.n238 585
R232 B.n240 B.n159 585
R233 B.n242 B.n241 585
R234 B.n243 B.n158 585
R235 B.n245 B.n244 585
R236 B.n246 B.n157 585
R237 B.n248 B.n247 585
R238 B.n249 B.n156 585
R239 B.n251 B.n250 585
R240 B.n252 B.n155 585
R241 B.n254 B.n253 585
R242 B.n255 B.n154 585
R243 B.n257 B.n256 585
R244 B.n258 B.n153 585
R245 B.n260 B.n259 585
R246 B.n261 B.n152 585
R247 B.n263 B.n262 585
R248 B.n264 B.n151 585
R249 B.n266 B.n265 585
R250 B.n267 B.n150 585
R251 B.n269 B.n268 585
R252 B.n270 B.n149 585
R253 B.n272 B.n271 585
R254 B.n273 B.n148 585
R255 B.n275 B.n274 585
R256 B.n276 B.n147 585
R257 B.n278 B.n277 585
R258 B.n279 B.n146 585
R259 B.n281 B.n280 585
R260 B.n282 B.n145 585
R261 B.n284 B.n283 585
R262 B.n285 B.n144 585
R263 B.n287 B.n286 585
R264 B.n288 B.n143 585
R265 B.n290 B.n289 585
R266 B.n291 B.n142 585
R267 B.n293 B.n292 585
R268 B.n294 B.n141 585
R269 B.n296 B.n295 585
R270 B.n298 B.n138 585
R271 B.n300 B.n299 585
R272 B.n301 B.n137 585
R273 B.n303 B.n302 585
R274 B.n304 B.n136 585
R275 B.n306 B.n305 585
R276 B.n307 B.n135 585
R277 B.n309 B.n308 585
R278 B.n310 B.n134 585
R279 B.n312 B.n311 585
R280 B.n314 B.n313 585
R281 B.n315 B.n130 585
R282 B.n317 B.n316 585
R283 B.n318 B.n129 585
R284 B.n320 B.n319 585
R285 B.n321 B.n128 585
R286 B.n323 B.n322 585
R287 B.n324 B.n127 585
R288 B.n326 B.n325 585
R289 B.n327 B.n126 585
R290 B.n329 B.n328 585
R291 B.n330 B.n125 585
R292 B.n332 B.n331 585
R293 B.n333 B.n124 585
R294 B.n335 B.n334 585
R295 B.n336 B.n123 585
R296 B.n338 B.n337 585
R297 B.n339 B.n122 585
R298 B.n341 B.n340 585
R299 B.n342 B.n121 585
R300 B.n344 B.n343 585
R301 B.n345 B.n120 585
R302 B.n347 B.n346 585
R303 B.n348 B.n119 585
R304 B.n350 B.n349 585
R305 B.n351 B.n118 585
R306 B.n353 B.n352 585
R307 B.n354 B.n117 585
R308 B.n356 B.n355 585
R309 B.n357 B.n116 585
R310 B.n359 B.n358 585
R311 B.n360 B.n115 585
R312 B.n362 B.n361 585
R313 B.n363 B.n114 585
R314 B.n365 B.n364 585
R315 B.n366 B.n113 585
R316 B.n368 B.n367 585
R317 B.n369 B.n112 585
R318 B.n371 B.n370 585
R319 B.n372 B.n111 585
R320 B.n374 B.n373 585
R321 B.n375 B.n110 585
R322 B.n377 B.n376 585
R323 B.n378 B.n109 585
R324 B.n380 B.n379 585
R325 B.n381 B.n108 585
R326 B.n383 B.n382 585
R327 B.n384 B.n107 585
R328 B.n386 B.n385 585
R329 B.n387 B.n106 585
R330 B.n389 B.n388 585
R331 B.n390 B.n105 585
R332 B.n392 B.n391 585
R333 B.n216 B.n167 585
R334 B.n215 B.n214 585
R335 B.n213 B.n168 585
R336 B.n212 B.n211 585
R337 B.n210 B.n169 585
R338 B.n209 B.n208 585
R339 B.n207 B.n170 585
R340 B.n206 B.n205 585
R341 B.n204 B.n171 585
R342 B.n203 B.n202 585
R343 B.n201 B.n172 585
R344 B.n200 B.n199 585
R345 B.n198 B.n173 585
R346 B.n197 B.n196 585
R347 B.n195 B.n174 585
R348 B.n194 B.n193 585
R349 B.n192 B.n175 585
R350 B.n191 B.n190 585
R351 B.n189 B.n176 585
R352 B.n188 B.n187 585
R353 B.n186 B.n177 585
R354 B.n185 B.n184 585
R355 B.n183 B.n178 585
R356 B.n182 B.n181 585
R357 B.n180 B.n179 585
R358 B.n2 B.n0 585
R359 B.n685 B.n1 585
R360 B.n684 B.n683 585
R361 B.n682 B.n3 585
R362 B.n681 B.n680 585
R363 B.n679 B.n4 585
R364 B.n678 B.n677 585
R365 B.n676 B.n5 585
R366 B.n675 B.n674 585
R367 B.n673 B.n6 585
R368 B.n672 B.n671 585
R369 B.n670 B.n7 585
R370 B.n669 B.n668 585
R371 B.n667 B.n8 585
R372 B.n666 B.n665 585
R373 B.n664 B.n9 585
R374 B.n663 B.n662 585
R375 B.n661 B.n10 585
R376 B.n660 B.n659 585
R377 B.n658 B.n11 585
R378 B.n657 B.n656 585
R379 B.n655 B.n12 585
R380 B.n654 B.n653 585
R381 B.n652 B.n13 585
R382 B.n651 B.n650 585
R383 B.n649 B.n14 585
R384 B.n648 B.n647 585
R385 B.n687 B.n686 585
R386 B.n217 B.n216 468.476
R387 B.n648 B.n15 468.476
R388 B.n391 B.n104 468.476
R389 B.n473 B.n78 468.476
R390 B.n131 B.t6 432.824
R391 B.n139 B.t9 432.824
R392 B.n42 B.t0 432.824
R393 B.n50 B.t3 432.824
R394 B.n216 B.n215 163.367
R395 B.n215 B.n168 163.367
R396 B.n211 B.n168 163.367
R397 B.n211 B.n210 163.367
R398 B.n210 B.n209 163.367
R399 B.n209 B.n170 163.367
R400 B.n205 B.n170 163.367
R401 B.n205 B.n204 163.367
R402 B.n204 B.n203 163.367
R403 B.n203 B.n172 163.367
R404 B.n199 B.n172 163.367
R405 B.n199 B.n198 163.367
R406 B.n198 B.n197 163.367
R407 B.n197 B.n174 163.367
R408 B.n193 B.n174 163.367
R409 B.n193 B.n192 163.367
R410 B.n192 B.n191 163.367
R411 B.n191 B.n176 163.367
R412 B.n187 B.n176 163.367
R413 B.n187 B.n186 163.367
R414 B.n186 B.n185 163.367
R415 B.n185 B.n178 163.367
R416 B.n181 B.n178 163.367
R417 B.n181 B.n180 163.367
R418 B.n180 B.n2 163.367
R419 B.n686 B.n2 163.367
R420 B.n686 B.n685 163.367
R421 B.n685 B.n684 163.367
R422 B.n684 B.n3 163.367
R423 B.n680 B.n3 163.367
R424 B.n680 B.n679 163.367
R425 B.n679 B.n678 163.367
R426 B.n678 B.n5 163.367
R427 B.n674 B.n5 163.367
R428 B.n674 B.n673 163.367
R429 B.n673 B.n672 163.367
R430 B.n672 B.n7 163.367
R431 B.n668 B.n7 163.367
R432 B.n668 B.n667 163.367
R433 B.n667 B.n666 163.367
R434 B.n666 B.n9 163.367
R435 B.n662 B.n9 163.367
R436 B.n662 B.n661 163.367
R437 B.n661 B.n660 163.367
R438 B.n660 B.n11 163.367
R439 B.n656 B.n11 163.367
R440 B.n656 B.n655 163.367
R441 B.n655 B.n654 163.367
R442 B.n654 B.n13 163.367
R443 B.n650 B.n13 163.367
R444 B.n650 B.n649 163.367
R445 B.n649 B.n648 163.367
R446 B.n217 B.n166 163.367
R447 B.n221 B.n166 163.367
R448 B.n222 B.n221 163.367
R449 B.n223 B.n222 163.367
R450 B.n223 B.n164 163.367
R451 B.n227 B.n164 163.367
R452 B.n228 B.n227 163.367
R453 B.n229 B.n228 163.367
R454 B.n229 B.n162 163.367
R455 B.n233 B.n162 163.367
R456 B.n234 B.n233 163.367
R457 B.n235 B.n234 163.367
R458 B.n235 B.n160 163.367
R459 B.n239 B.n160 163.367
R460 B.n240 B.n239 163.367
R461 B.n241 B.n240 163.367
R462 B.n241 B.n158 163.367
R463 B.n245 B.n158 163.367
R464 B.n246 B.n245 163.367
R465 B.n247 B.n246 163.367
R466 B.n247 B.n156 163.367
R467 B.n251 B.n156 163.367
R468 B.n252 B.n251 163.367
R469 B.n253 B.n252 163.367
R470 B.n253 B.n154 163.367
R471 B.n257 B.n154 163.367
R472 B.n258 B.n257 163.367
R473 B.n259 B.n258 163.367
R474 B.n259 B.n152 163.367
R475 B.n263 B.n152 163.367
R476 B.n264 B.n263 163.367
R477 B.n265 B.n264 163.367
R478 B.n265 B.n150 163.367
R479 B.n269 B.n150 163.367
R480 B.n270 B.n269 163.367
R481 B.n271 B.n270 163.367
R482 B.n271 B.n148 163.367
R483 B.n275 B.n148 163.367
R484 B.n276 B.n275 163.367
R485 B.n277 B.n276 163.367
R486 B.n277 B.n146 163.367
R487 B.n281 B.n146 163.367
R488 B.n282 B.n281 163.367
R489 B.n283 B.n282 163.367
R490 B.n283 B.n144 163.367
R491 B.n287 B.n144 163.367
R492 B.n288 B.n287 163.367
R493 B.n289 B.n288 163.367
R494 B.n289 B.n142 163.367
R495 B.n293 B.n142 163.367
R496 B.n294 B.n293 163.367
R497 B.n295 B.n294 163.367
R498 B.n295 B.n138 163.367
R499 B.n300 B.n138 163.367
R500 B.n301 B.n300 163.367
R501 B.n302 B.n301 163.367
R502 B.n302 B.n136 163.367
R503 B.n306 B.n136 163.367
R504 B.n307 B.n306 163.367
R505 B.n308 B.n307 163.367
R506 B.n308 B.n134 163.367
R507 B.n312 B.n134 163.367
R508 B.n313 B.n312 163.367
R509 B.n313 B.n130 163.367
R510 B.n317 B.n130 163.367
R511 B.n318 B.n317 163.367
R512 B.n319 B.n318 163.367
R513 B.n319 B.n128 163.367
R514 B.n323 B.n128 163.367
R515 B.n324 B.n323 163.367
R516 B.n325 B.n324 163.367
R517 B.n325 B.n126 163.367
R518 B.n329 B.n126 163.367
R519 B.n330 B.n329 163.367
R520 B.n331 B.n330 163.367
R521 B.n331 B.n124 163.367
R522 B.n335 B.n124 163.367
R523 B.n336 B.n335 163.367
R524 B.n337 B.n336 163.367
R525 B.n337 B.n122 163.367
R526 B.n341 B.n122 163.367
R527 B.n342 B.n341 163.367
R528 B.n343 B.n342 163.367
R529 B.n343 B.n120 163.367
R530 B.n347 B.n120 163.367
R531 B.n348 B.n347 163.367
R532 B.n349 B.n348 163.367
R533 B.n349 B.n118 163.367
R534 B.n353 B.n118 163.367
R535 B.n354 B.n353 163.367
R536 B.n355 B.n354 163.367
R537 B.n355 B.n116 163.367
R538 B.n359 B.n116 163.367
R539 B.n360 B.n359 163.367
R540 B.n361 B.n360 163.367
R541 B.n361 B.n114 163.367
R542 B.n365 B.n114 163.367
R543 B.n366 B.n365 163.367
R544 B.n367 B.n366 163.367
R545 B.n367 B.n112 163.367
R546 B.n371 B.n112 163.367
R547 B.n372 B.n371 163.367
R548 B.n373 B.n372 163.367
R549 B.n373 B.n110 163.367
R550 B.n377 B.n110 163.367
R551 B.n378 B.n377 163.367
R552 B.n379 B.n378 163.367
R553 B.n379 B.n108 163.367
R554 B.n383 B.n108 163.367
R555 B.n384 B.n383 163.367
R556 B.n385 B.n384 163.367
R557 B.n385 B.n106 163.367
R558 B.n389 B.n106 163.367
R559 B.n390 B.n389 163.367
R560 B.n391 B.n390 163.367
R561 B.n395 B.n104 163.367
R562 B.n396 B.n395 163.367
R563 B.n397 B.n396 163.367
R564 B.n397 B.n102 163.367
R565 B.n401 B.n102 163.367
R566 B.n402 B.n401 163.367
R567 B.n403 B.n402 163.367
R568 B.n403 B.n100 163.367
R569 B.n407 B.n100 163.367
R570 B.n408 B.n407 163.367
R571 B.n409 B.n408 163.367
R572 B.n409 B.n98 163.367
R573 B.n413 B.n98 163.367
R574 B.n414 B.n413 163.367
R575 B.n415 B.n414 163.367
R576 B.n415 B.n96 163.367
R577 B.n419 B.n96 163.367
R578 B.n420 B.n419 163.367
R579 B.n421 B.n420 163.367
R580 B.n421 B.n94 163.367
R581 B.n425 B.n94 163.367
R582 B.n426 B.n425 163.367
R583 B.n427 B.n426 163.367
R584 B.n427 B.n92 163.367
R585 B.n431 B.n92 163.367
R586 B.n432 B.n431 163.367
R587 B.n433 B.n432 163.367
R588 B.n433 B.n90 163.367
R589 B.n437 B.n90 163.367
R590 B.n438 B.n437 163.367
R591 B.n439 B.n438 163.367
R592 B.n439 B.n88 163.367
R593 B.n443 B.n88 163.367
R594 B.n444 B.n443 163.367
R595 B.n445 B.n444 163.367
R596 B.n445 B.n86 163.367
R597 B.n449 B.n86 163.367
R598 B.n450 B.n449 163.367
R599 B.n451 B.n450 163.367
R600 B.n451 B.n84 163.367
R601 B.n455 B.n84 163.367
R602 B.n456 B.n455 163.367
R603 B.n457 B.n456 163.367
R604 B.n457 B.n82 163.367
R605 B.n461 B.n82 163.367
R606 B.n462 B.n461 163.367
R607 B.n463 B.n462 163.367
R608 B.n463 B.n80 163.367
R609 B.n467 B.n80 163.367
R610 B.n468 B.n467 163.367
R611 B.n469 B.n468 163.367
R612 B.n469 B.n78 163.367
R613 B.n644 B.n15 163.367
R614 B.n644 B.n643 163.367
R615 B.n643 B.n642 163.367
R616 B.n642 B.n17 163.367
R617 B.n638 B.n17 163.367
R618 B.n638 B.n637 163.367
R619 B.n637 B.n636 163.367
R620 B.n636 B.n19 163.367
R621 B.n632 B.n19 163.367
R622 B.n632 B.n631 163.367
R623 B.n631 B.n630 163.367
R624 B.n630 B.n21 163.367
R625 B.n626 B.n21 163.367
R626 B.n626 B.n625 163.367
R627 B.n625 B.n624 163.367
R628 B.n624 B.n23 163.367
R629 B.n620 B.n23 163.367
R630 B.n620 B.n619 163.367
R631 B.n619 B.n618 163.367
R632 B.n618 B.n25 163.367
R633 B.n614 B.n25 163.367
R634 B.n614 B.n613 163.367
R635 B.n613 B.n612 163.367
R636 B.n612 B.n27 163.367
R637 B.n608 B.n27 163.367
R638 B.n608 B.n607 163.367
R639 B.n607 B.n606 163.367
R640 B.n606 B.n29 163.367
R641 B.n602 B.n29 163.367
R642 B.n602 B.n601 163.367
R643 B.n601 B.n600 163.367
R644 B.n600 B.n31 163.367
R645 B.n596 B.n31 163.367
R646 B.n596 B.n595 163.367
R647 B.n595 B.n594 163.367
R648 B.n594 B.n33 163.367
R649 B.n590 B.n33 163.367
R650 B.n590 B.n589 163.367
R651 B.n589 B.n588 163.367
R652 B.n588 B.n35 163.367
R653 B.n584 B.n35 163.367
R654 B.n584 B.n583 163.367
R655 B.n583 B.n582 163.367
R656 B.n582 B.n37 163.367
R657 B.n578 B.n37 163.367
R658 B.n578 B.n577 163.367
R659 B.n577 B.n576 163.367
R660 B.n576 B.n39 163.367
R661 B.n572 B.n39 163.367
R662 B.n572 B.n571 163.367
R663 B.n571 B.n570 163.367
R664 B.n570 B.n41 163.367
R665 B.n565 B.n41 163.367
R666 B.n565 B.n564 163.367
R667 B.n564 B.n563 163.367
R668 B.n563 B.n45 163.367
R669 B.n559 B.n45 163.367
R670 B.n559 B.n558 163.367
R671 B.n558 B.n557 163.367
R672 B.n557 B.n47 163.367
R673 B.n553 B.n47 163.367
R674 B.n553 B.n552 163.367
R675 B.n552 B.n551 163.367
R676 B.n551 B.n49 163.367
R677 B.n547 B.n49 163.367
R678 B.n547 B.n546 163.367
R679 B.n546 B.n545 163.367
R680 B.n545 B.n54 163.367
R681 B.n541 B.n54 163.367
R682 B.n541 B.n540 163.367
R683 B.n540 B.n539 163.367
R684 B.n539 B.n56 163.367
R685 B.n535 B.n56 163.367
R686 B.n535 B.n534 163.367
R687 B.n534 B.n533 163.367
R688 B.n533 B.n58 163.367
R689 B.n529 B.n58 163.367
R690 B.n529 B.n528 163.367
R691 B.n528 B.n527 163.367
R692 B.n527 B.n60 163.367
R693 B.n523 B.n60 163.367
R694 B.n523 B.n522 163.367
R695 B.n522 B.n521 163.367
R696 B.n521 B.n62 163.367
R697 B.n517 B.n62 163.367
R698 B.n517 B.n516 163.367
R699 B.n516 B.n515 163.367
R700 B.n515 B.n64 163.367
R701 B.n511 B.n64 163.367
R702 B.n511 B.n510 163.367
R703 B.n510 B.n509 163.367
R704 B.n509 B.n66 163.367
R705 B.n505 B.n66 163.367
R706 B.n505 B.n504 163.367
R707 B.n504 B.n503 163.367
R708 B.n503 B.n68 163.367
R709 B.n499 B.n68 163.367
R710 B.n499 B.n498 163.367
R711 B.n498 B.n497 163.367
R712 B.n497 B.n70 163.367
R713 B.n493 B.n70 163.367
R714 B.n493 B.n492 163.367
R715 B.n492 B.n491 163.367
R716 B.n491 B.n72 163.367
R717 B.n487 B.n72 163.367
R718 B.n487 B.n486 163.367
R719 B.n486 B.n485 163.367
R720 B.n485 B.n74 163.367
R721 B.n481 B.n74 163.367
R722 B.n481 B.n480 163.367
R723 B.n480 B.n479 163.367
R724 B.n479 B.n76 163.367
R725 B.n475 B.n76 163.367
R726 B.n475 B.n474 163.367
R727 B.n474 B.n473 163.367
R728 B.n131 B.t8 150.657
R729 B.n50 B.t4 150.657
R730 B.n139 B.t11 150.637
R731 B.n42 B.t1 150.637
R732 B.n132 B.t7 111.481
R733 B.n51 B.t5 111.481
R734 B.n140 B.t10 111.462
R735 B.n43 B.t2 111.462
R736 B.n133 B.n132 59.5399
R737 B.n297 B.n140 59.5399
R738 B.n567 B.n43 59.5399
R739 B.n52 B.n51 59.5399
R740 B.n132 B.n131 39.1763
R741 B.n140 B.n139 39.1763
R742 B.n43 B.n42 39.1763
R743 B.n51 B.n50 39.1763
R744 B.n647 B.n646 30.4395
R745 B.n472 B.n471 30.4395
R746 B.n393 B.n392 30.4395
R747 B.n218 B.n167 30.4395
R748 B B.n687 18.0485
R749 B.n646 B.n645 10.6151
R750 B.n645 B.n16 10.6151
R751 B.n641 B.n16 10.6151
R752 B.n641 B.n640 10.6151
R753 B.n640 B.n639 10.6151
R754 B.n639 B.n18 10.6151
R755 B.n635 B.n18 10.6151
R756 B.n635 B.n634 10.6151
R757 B.n634 B.n633 10.6151
R758 B.n633 B.n20 10.6151
R759 B.n629 B.n20 10.6151
R760 B.n629 B.n628 10.6151
R761 B.n628 B.n627 10.6151
R762 B.n627 B.n22 10.6151
R763 B.n623 B.n22 10.6151
R764 B.n623 B.n622 10.6151
R765 B.n622 B.n621 10.6151
R766 B.n621 B.n24 10.6151
R767 B.n617 B.n24 10.6151
R768 B.n617 B.n616 10.6151
R769 B.n616 B.n615 10.6151
R770 B.n615 B.n26 10.6151
R771 B.n611 B.n26 10.6151
R772 B.n611 B.n610 10.6151
R773 B.n610 B.n609 10.6151
R774 B.n609 B.n28 10.6151
R775 B.n605 B.n28 10.6151
R776 B.n605 B.n604 10.6151
R777 B.n604 B.n603 10.6151
R778 B.n603 B.n30 10.6151
R779 B.n599 B.n30 10.6151
R780 B.n599 B.n598 10.6151
R781 B.n598 B.n597 10.6151
R782 B.n597 B.n32 10.6151
R783 B.n593 B.n32 10.6151
R784 B.n593 B.n592 10.6151
R785 B.n592 B.n591 10.6151
R786 B.n591 B.n34 10.6151
R787 B.n587 B.n34 10.6151
R788 B.n587 B.n586 10.6151
R789 B.n586 B.n585 10.6151
R790 B.n585 B.n36 10.6151
R791 B.n581 B.n36 10.6151
R792 B.n581 B.n580 10.6151
R793 B.n580 B.n579 10.6151
R794 B.n579 B.n38 10.6151
R795 B.n575 B.n38 10.6151
R796 B.n575 B.n574 10.6151
R797 B.n574 B.n573 10.6151
R798 B.n573 B.n40 10.6151
R799 B.n569 B.n40 10.6151
R800 B.n569 B.n568 10.6151
R801 B.n566 B.n44 10.6151
R802 B.n562 B.n44 10.6151
R803 B.n562 B.n561 10.6151
R804 B.n561 B.n560 10.6151
R805 B.n560 B.n46 10.6151
R806 B.n556 B.n46 10.6151
R807 B.n556 B.n555 10.6151
R808 B.n555 B.n554 10.6151
R809 B.n554 B.n48 10.6151
R810 B.n550 B.n549 10.6151
R811 B.n549 B.n548 10.6151
R812 B.n548 B.n53 10.6151
R813 B.n544 B.n53 10.6151
R814 B.n544 B.n543 10.6151
R815 B.n543 B.n542 10.6151
R816 B.n542 B.n55 10.6151
R817 B.n538 B.n55 10.6151
R818 B.n538 B.n537 10.6151
R819 B.n537 B.n536 10.6151
R820 B.n536 B.n57 10.6151
R821 B.n532 B.n57 10.6151
R822 B.n532 B.n531 10.6151
R823 B.n531 B.n530 10.6151
R824 B.n530 B.n59 10.6151
R825 B.n526 B.n59 10.6151
R826 B.n526 B.n525 10.6151
R827 B.n525 B.n524 10.6151
R828 B.n524 B.n61 10.6151
R829 B.n520 B.n61 10.6151
R830 B.n520 B.n519 10.6151
R831 B.n519 B.n518 10.6151
R832 B.n518 B.n63 10.6151
R833 B.n514 B.n63 10.6151
R834 B.n514 B.n513 10.6151
R835 B.n513 B.n512 10.6151
R836 B.n512 B.n65 10.6151
R837 B.n508 B.n65 10.6151
R838 B.n508 B.n507 10.6151
R839 B.n507 B.n506 10.6151
R840 B.n506 B.n67 10.6151
R841 B.n502 B.n67 10.6151
R842 B.n502 B.n501 10.6151
R843 B.n501 B.n500 10.6151
R844 B.n500 B.n69 10.6151
R845 B.n496 B.n69 10.6151
R846 B.n496 B.n495 10.6151
R847 B.n495 B.n494 10.6151
R848 B.n494 B.n71 10.6151
R849 B.n490 B.n71 10.6151
R850 B.n490 B.n489 10.6151
R851 B.n489 B.n488 10.6151
R852 B.n488 B.n73 10.6151
R853 B.n484 B.n73 10.6151
R854 B.n484 B.n483 10.6151
R855 B.n483 B.n482 10.6151
R856 B.n482 B.n75 10.6151
R857 B.n478 B.n75 10.6151
R858 B.n478 B.n477 10.6151
R859 B.n477 B.n476 10.6151
R860 B.n476 B.n77 10.6151
R861 B.n472 B.n77 10.6151
R862 B.n394 B.n393 10.6151
R863 B.n394 B.n103 10.6151
R864 B.n398 B.n103 10.6151
R865 B.n399 B.n398 10.6151
R866 B.n400 B.n399 10.6151
R867 B.n400 B.n101 10.6151
R868 B.n404 B.n101 10.6151
R869 B.n405 B.n404 10.6151
R870 B.n406 B.n405 10.6151
R871 B.n406 B.n99 10.6151
R872 B.n410 B.n99 10.6151
R873 B.n411 B.n410 10.6151
R874 B.n412 B.n411 10.6151
R875 B.n412 B.n97 10.6151
R876 B.n416 B.n97 10.6151
R877 B.n417 B.n416 10.6151
R878 B.n418 B.n417 10.6151
R879 B.n418 B.n95 10.6151
R880 B.n422 B.n95 10.6151
R881 B.n423 B.n422 10.6151
R882 B.n424 B.n423 10.6151
R883 B.n424 B.n93 10.6151
R884 B.n428 B.n93 10.6151
R885 B.n429 B.n428 10.6151
R886 B.n430 B.n429 10.6151
R887 B.n430 B.n91 10.6151
R888 B.n434 B.n91 10.6151
R889 B.n435 B.n434 10.6151
R890 B.n436 B.n435 10.6151
R891 B.n436 B.n89 10.6151
R892 B.n440 B.n89 10.6151
R893 B.n441 B.n440 10.6151
R894 B.n442 B.n441 10.6151
R895 B.n442 B.n87 10.6151
R896 B.n446 B.n87 10.6151
R897 B.n447 B.n446 10.6151
R898 B.n448 B.n447 10.6151
R899 B.n448 B.n85 10.6151
R900 B.n452 B.n85 10.6151
R901 B.n453 B.n452 10.6151
R902 B.n454 B.n453 10.6151
R903 B.n454 B.n83 10.6151
R904 B.n458 B.n83 10.6151
R905 B.n459 B.n458 10.6151
R906 B.n460 B.n459 10.6151
R907 B.n460 B.n81 10.6151
R908 B.n464 B.n81 10.6151
R909 B.n465 B.n464 10.6151
R910 B.n466 B.n465 10.6151
R911 B.n466 B.n79 10.6151
R912 B.n470 B.n79 10.6151
R913 B.n471 B.n470 10.6151
R914 B.n219 B.n218 10.6151
R915 B.n220 B.n219 10.6151
R916 B.n220 B.n165 10.6151
R917 B.n224 B.n165 10.6151
R918 B.n225 B.n224 10.6151
R919 B.n226 B.n225 10.6151
R920 B.n226 B.n163 10.6151
R921 B.n230 B.n163 10.6151
R922 B.n231 B.n230 10.6151
R923 B.n232 B.n231 10.6151
R924 B.n232 B.n161 10.6151
R925 B.n236 B.n161 10.6151
R926 B.n237 B.n236 10.6151
R927 B.n238 B.n237 10.6151
R928 B.n238 B.n159 10.6151
R929 B.n242 B.n159 10.6151
R930 B.n243 B.n242 10.6151
R931 B.n244 B.n243 10.6151
R932 B.n244 B.n157 10.6151
R933 B.n248 B.n157 10.6151
R934 B.n249 B.n248 10.6151
R935 B.n250 B.n249 10.6151
R936 B.n250 B.n155 10.6151
R937 B.n254 B.n155 10.6151
R938 B.n255 B.n254 10.6151
R939 B.n256 B.n255 10.6151
R940 B.n256 B.n153 10.6151
R941 B.n260 B.n153 10.6151
R942 B.n261 B.n260 10.6151
R943 B.n262 B.n261 10.6151
R944 B.n262 B.n151 10.6151
R945 B.n266 B.n151 10.6151
R946 B.n267 B.n266 10.6151
R947 B.n268 B.n267 10.6151
R948 B.n268 B.n149 10.6151
R949 B.n272 B.n149 10.6151
R950 B.n273 B.n272 10.6151
R951 B.n274 B.n273 10.6151
R952 B.n274 B.n147 10.6151
R953 B.n278 B.n147 10.6151
R954 B.n279 B.n278 10.6151
R955 B.n280 B.n279 10.6151
R956 B.n280 B.n145 10.6151
R957 B.n284 B.n145 10.6151
R958 B.n285 B.n284 10.6151
R959 B.n286 B.n285 10.6151
R960 B.n286 B.n143 10.6151
R961 B.n290 B.n143 10.6151
R962 B.n291 B.n290 10.6151
R963 B.n292 B.n291 10.6151
R964 B.n292 B.n141 10.6151
R965 B.n296 B.n141 10.6151
R966 B.n299 B.n298 10.6151
R967 B.n299 B.n137 10.6151
R968 B.n303 B.n137 10.6151
R969 B.n304 B.n303 10.6151
R970 B.n305 B.n304 10.6151
R971 B.n305 B.n135 10.6151
R972 B.n309 B.n135 10.6151
R973 B.n310 B.n309 10.6151
R974 B.n311 B.n310 10.6151
R975 B.n315 B.n314 10.6151
R976 B.n316 B.n315 10.6151
R977 B.n316 B.n129 10.6151
R978 B.n320 B.n129 10.6151
R979 B.n321 B.n320 10.6151
R980 B.n322 B.n321 10.6151
R981 B.n322 B.n127 10.6151
R982 B.n326 B.n127 10.6151
R983 B.n327 B.n326 10.6151
R984 B.n328 B.n327 10.6151
R985 B.n328 B.n125 10.6151
R986 B.n332 B.n125 10.6151
R987 B.n333 B.n332 10.6151
R988 B.n334 B.n333 10.6151
R989 B.n334 B.n123 10.6151
R990 B.n338 B.n123 10.6151
R991 B.n339 B.n338 10.6151
R992 B.n340 B.n339 10.6151
R993 B.n340 B.n121 10.6151
R994 B.n344 B.n121 10.6151
R995 B.n345 B.n344 10.6151
R996 B.n346 B.n345 10.6151
R997 B.n346 B.n119 10.6151
R998 B.n350 B.n119 10.6151
R999 B.n351 B.n350 10.6151
R1000 B.n352 B.n351 10.6151
R1001 B.n352 B.n117 10.6151
R1002 B.n356 B.n117 10.6151
R1003 B.n357 B.n356 10.6151
R1004 B.n358 B.n357 10.6151
R1005 B.n358 B.n115 10.6151
R1006 B.n362 B.n115 10.6151
R1007 B.n363 B.n362 10.6151
R1008 B.n364 B.n363 10.6151
R1009 B.n364 B.n113 10.6151
R1010 B.n368 B.n113 10.6151
R1011 B.n369 B.n368 10.6151
R1012 B.n370 B.n369 10.6151
R1013 B.n370 B.n111 10.6151
R1014 B.n374 B.n111 10.6151
R1015 B.n375 B.n374 10.6151
R1016 B.n376 B.n375 10.6151
R1017 B.n376 B.n109 10.6151
R1018 B.n380 B.n109 10.6151
R1019 B.n381 B.n380 10.6151
R1020 B.n382 B.n381 10.6151
R1021 B.n382 B.n107 10.6151
R1022 B.n386 B.n107 10.6151
R1023 B.n387 B.n386 10.6151
R1024 B.n388 B.n387 10.6151
R1025 B.n388 B.n105 10.6151
R1026 B.n392 B.n105 10.6151
R1027 B.n214 B.n167 10.6151
R1028 B.n214 B.n213 10.6151
R1029 B.n213 B.n212 10.6151
R1030 B.n212 B.n169 10.6151
R1031 B.n208 B.n169 10.6151
R1032 B.n208 B.n207 10.6151
R1033 B.n207 B.n206 10.6151
R1034 B.n206 B.n171 10.6151
R1035 B.n202 B.n171 10.6151
R1036 B.n202 B.n201 10.6151
R1037 B.n201 B.n200 10.6151
R1038 B.n200 B.n173 10.6151
R1039 B.n196 B.n173 10.6151
R1040 B.n196 B.n195 10.6151
R1041 B.n195 B.n194 10.6151
R1042 B.n194 B.n175 10.6151
R1043 B.n190 B.n175 10.6151
R1044 B.n190 B.n189 10.6151
R1045 B.n189 B.n188 10.6151
R1046 B.n188 B.n177 10.6151
R1047 B.n184 B.n177 10.6151
R1048 B.n184 B.n183 10.6151
R1049 B.n183 B.n182 10.6151
R1050 B.n182 B.n179 10.6151
R1051 B.n179 B.n0 10.6151
R1052 B.n683 B.n1 10.6151
R1053 B.n683 B.n682 10.6151
R1054 B.n682 B.n681 10.6151
R1055 B.n681 B.n4 10.6151
R1056 B.n677 B.n4 10.6151
R1057 B.n677 B.n676 10.6151
R1058 B.n676 B.n675 10.6151
R1059 B.n675 B.n6 10.6151
R1060 B.n671 B.n6 10.6151
R1061 B.n671 B.n670 10.6151
R1062 B.n670 B.n669 10.6151
R1063 B.n669 B.n8 10.6151
R1064 B.n665 B.n8 10.6151
R1065 B.n665 B.n664 10.6151
R1066 B.n664 B.n663 10.6151
R1067 B.n663 B.n10 10.6151
R1068 B.n659 B.n10 10.6151
R1069 B.n659 B.n658 10.6151
R1070 B.n658 B.n657 10.6151
R1071 B.n657 B.n12 10.6151
R1072 B.n653 B.n12 10.6151
R1073 B.n653 B.n652 10.6151
R1074 B.n652 B.n651 10.6151
R1075 B.n651 B.n14 10.6151
R1076 B.n647 B.n14 10.6151
R1077 B.n568 B.n567 9.36635
R1078 B.n550 B.n52 9.36635
R1079 B.n297 B.n296 9.36635
R1080 B.n314 B.n133 9.36635
R1081 B.n687 B.n0 2.81026
R1082 B.n687 B.n1 2.81026
R1083 B.n567 B.n566 1.24928
R1084 B.n52 B.n48 1.24928
R1085 B.n298 B.n297 1.24928
R1086 B.n311 B.n133 1.24928
R1087 VN.n0 VN.t1 261.692
R1088 VN.n1 VN.t0 261.692
R1089 VN.n0 VN.t3 261.271
R1090 VN.n1 VN.t2 261.271
R1091 VN VN.n1 56.2534
R1092 VN VN.n0 9.56781
R1093 VDD2.n2 VDD2.n0 116.16
R1094 VDD2.n2 VDD2.n1 73.5145
R1095 VDD2.n1 VDD2.t1 2.04484
R1096 VDD2.n1 VDD2.t3 2.04484
R1097 VDD2.n0 VDD2.t2 2.04484
R1098 VDD2.n0 VDD2.t0 2.04484
R1099 VDD2 VDD2.n2 0.0586897
C0 B VN 0.984837f
C1 VTAIL B 5.68208f
C2 B VDD2 1.24418f
C3 VTAIL VN 5.25255f
C4 VP B 1.44227f
C5 w_n2182_n4148# B 9.21935f
C6 VDD2 VN 5.63579f
C7 VP VN 6.25722f
C8 w_n2182_n4148# VN 3.60692f
C9 VTAIL VDD2 6.60793f
C10 VP VTAIL 5.26666f
C11 VDD1 B 1.20689f
C12 w_n2182_n4148# VTAIL 4.89205f
C13 VP VDD2 0.336555f
C14 VDD1 VN 0.148332f
C15 w_n2182_n4148# VDD2 1.41167f
C16 VP w_n2182_n4148# 3.88513f
C17 VDD1 VTAIL 6.55982f
C18 VDD1 VDD2 0.804487f
C19 VDD1 VP 5.82351f
C20 VDD1 w_n2182_n4148# 1.37591f
C21 VDD2 VSUBS 0.899029f
C22 VDD1 VSUBS 5.7682f
C23 VTAIL VSUBS 1.260888f
C24 VN VSUBS 5.34816f
C25 VP VSUBS 1.933729f
C26 B VSUBS 3.817887f
C27 w_n2182_n4148# VSUBS 0.110889p
C28 VDD2.t2 VSUBS 0.332873f
C29 VDD2.t0 VSUBS 0.332873f
C30 VDD2.n0 VSUBS 3.51862f
C31 VDD2.t1 VSUBS 0.332873f
C32 VDD2.t3 VSUBS 0.332873f
C33 VDD2.n1 VSUBS 2.7364f
C34 VDD2.n2 VSUBS 4.45913f
C35 VN.t1 VSUBS 3.03965f
C36 VN.t3 VSUBS 3.0377f
C37 VN.n0 VSUBS 2.13622f
C38 VN.t0 VSUBS 3.03965f
C39 VN.t2 VSUBS 3.0377f
C40 VN.n1 VSUBS 3.93827f
C41 B.n0 VSUBS 0.004345f
C42 B.n1 VSUBS 0.004345f
C43 B.n2 VSUBS 0.006871f
C44 B.n3 VSUBS 0.006871f
C45 B.n4 VSUBS 0.006871f
C46 B.n5 VSUBS 0.006871f
C47 B.n6 VSUBS 0.006871f
C48 B.n7 VSUBS 0.006871f
C49 B.n8 VSUBS 0.006871f
C50 B.n9 VSUBS 0.006871f
C51 B.n10 VSUBS 0.006871f
C52 B.n11 VSUBS 0.006871f
C53 B.n12 VSUBS 0.006871f
C54 B.n13 VSUBS 0.006871f
C55 B.n14 VSUBS 0.006871f
C56 B.n15 VSUBS 0.015814f
C57 B.n16 VSUBS 0.006871f
C58 B.n17 VSUBS 0.006871f
C59 B.n18 VSUBS 0.006871f
C60 B.n19 VSUBS 0.006871f
C61 B.n20 VSUBS 0.006871f
C62 B.n21 VSUBS 0.006871f
C63 B.n22 VSUBS 0.006871f
C64 B.n23 VSUBS 0.006871f
C65 B.n24 VSUBS 0.006871f
C66 B.n25 VSUBS 0.006871f
C67 B.n26 VSUBS 0.006871f
C68 B.n27 VSUBS 0.006871f
C69 B.n28 VSUBS 0.006871f
C70 B.n29 VSUBS 0.006871f
C71 B.n30 VSUBS 0.006871f
C72 B.n31 VSUBS 0.006871f
C73 B.n32 VSUBS 0.006871f
C74 B.n33 VSUBS 0.006871f
C75 B.n34 VSUBS 0.006871f
C76 B.n35 VSUBS 0.006871f
C77 B.n36 VSUBS 0.006871f
C78 B.n37 VSUBS 0.006871f
C79 B.n38 VSUBS 0.006871f
C80 B.n39 VSUBS 0.006871f
C81 B.n40 VSUBS 0.006871f
C82 B.n41 VSUBS 0.006871f
C83 B.t2 VSUBS 0.522021f
C84 B.t1 VSUBS 0.53689f
C85 B.t0 VSUBS 1.14174f
C86 B.n42 VSUBS 0.246736f
C87 B.n43 VSUBS 0.066974f
C88 B.n44 VSUBS 0.006871f
C89 B.n45 VSUBS 0.006871f
C90 B.n46 VSUBS 0.006871f
C91 B.n47 VSUBS 0.006871f
C92 B.n48 VSUBS 0.003839f
C93 B.n49 VSUBS 0.006871f
C94 B.t5 VSUBS 0.522006f
C95 B.t4 VSUBS 0.536877f
C96 B.t3 VSUBS 1.14174f
C97 B.n50 VSUBS 0.24675f
C98 B.n51 VSUBS 0.06699f
C99 B.n52 VSUBS 0.015918f
C100 B.n53 VSUBS 0.006871f
C101 B.n54 VSUBS 0.006871f
C102 B.n55 VSUBS 0.006871f
C103 B.n56 VSUBS 0.006871f
C104 B.n57 VSUBS 0.006871f
C105 B.n58 VSUBS 0.006871f
C106 B.n59 VSUBS 0.006871f
C107 B.n60 VSUBS 0.006871f
C108 B.n61 VSUBS 0.006871f
C109 B.n62 VSUBS 0.006871f
C110 B.n63 VSUBS 0.006871f
C111 B.n64 VSUBS 0.006871f
C112 B.n65 VSUBS 0.006871f
C113 B.n66 VSUBS 0.006871f
C114 B.n67 VSUBS 0.006871f
C115 B.n68 VSUBS 0.006871f
C116 B.n69 VSUBS 0.006871f
C117 B.n70 VSUBS 0.006871f
C118 B.n71 VSUBS 0.006871f
C119 B.n72 VSUBS 0.006871f
C120 B.n73 VSUBS 0.006871f
C121 B.n74 VSUBS 0.006871f
C122 B.n75 VSUBS 0.006871f
C123 B.n76 VSUBS 0.006871f
C124 B.n77 VSUBS 0.006871f
C125 B.n78 VSUBS 0.014901f
C126 B.n79 VSUBS 0.006871f
C127 B.n80 VSUBS 0.006871f
C128 B.n81 VSUBS 0.006871f
C129 B.n82 VSUBS 0.006871f
C130 B.n83 VSUBS 0.006871f
C131 B.n84 VSUBS 0.006871f
C132 B.n85 VSUBS 0.006871f
C133 B.n86 VSUBS 0.006871f
C134 B.n87 VSUBS 0.006871f
C135 B.n88 VSUBS 0.006871f
C136 B.n89 VSUBS 0.006871f
C137 B.n90 VSUBS 0.006871f
C138 B.n91 VSUBS 0.006871f
C139 B.n92 VSUBS 0.006871f
C140 B.n93 VSUBS 0.006871f
C141 B.n94 VSUBS 0.006871f
C142 B.n95 VSUBS 0.006871f
C143 B.n96 VSUBS 0.006871f
C144 B.n97 VSUBS 0.006871f
C145 B.n98 VSUBS 0.006871f
C146 B.n99 VSUBS 0.006871f
C147 B.n100 VSUBS 0.006871f
C148 B.n101 VSUBS 0.006871f
C149 B.n102 VSUBS 0.006871f
C150 B.n103 VSUBS 0.006871f
C151 B.n104 VSUBS 0.014901f
C152 B.n105 VSUBS 0.006871f
C153 B.n106 VSUBS 0.006871f
C154 B.n107 VSUBS 0.006871f
C155 B.n108 VSUBS 0.006871f
C156 B.n109 VSUBS 0.006871f
C157 B.n110 VSUBS 0.006871f
C158 B.n111 VSUBS 0.006871f
C159 B.n112 VSUBS 0.006871f
C160 B.n113 VSUBS 0.006871f
C161 B.n114 VSUBS 0.006871f
C162 B.n115 VSUBS 0.006871f
C163 B.n116 VSUBS 0.006871f
C164 B.n117 VSUBS 0.006871f
C165 B.n118 VSUBS 0.006871f
C166 B.n119 VSUBS 0.006871f
C167 B.n120 VSUBS 0.006871f
C168 B.n121 VSUBS 0.006871f
C169 B.n122 VSUBS 0.006871f
C170 B.n123 VSUBS 0.006871f
C171 B.n124 VSUBS 0.006871f
C172 B.n125 VSUBS 0.006871f
C173 B.n126 VSUBS 0.006871f
C174 B.n127 VSUBS 0.006871f
C175 B.n128 VSUBS 0.006871f
C176 B.n129 VSUBS 0.006871f
C177 B.n130 VSUBS 0.006871f
C178 B.t7 VSUBS 0.522006f
C179 B.t8 VSUBS 0.536877f
C180 B.t6 VSUBS 1.14174f
C181 B.n131 VSUBS 0.24675f
C182 B.n132 VSUBS 0.06699f
C183 B.n133 VSUBS 0.015918f
C184 B.n134 VSUBS 0.006871f
C185 B.n135 VSUBS 0.006871f
C186 B.n136 VSUBS 0.006871f
C187 B.n137 VSUBS 0.006871f
C188 B.n138 VSUBS 0.006871f
C189 B.t10 VSUBS 0.522021f
C190 B.t11 VSUBS 0.53689f
C191 B.t9 VSUBS 1.14174f
C192 B.n139 VSUBS 0.246736f
C193 B.n140 VSUBS 0.066974f
C194 B.n141 VSUBS 0.006871f
C195 B.n142 VSUBS 0.006871f
C196 B.n143 VSUBS 0.006871f
C197 B.n144 VSUBS 0.006871f
C198 B.n145 VSUBS 0.006871f
C199 B.n146 VSUBS 0.006871f
C200 B.n147 VSUBS 0.006871f
C201 B.n148 VSUBS 0.006871f
C202 B.n149 VSUBS 0.006871f
C203 B.n150 VSUBS 0.006871f
C204 B.n151 VSUBS 0.006871f
C205 B.n152 VSUBS 0.006871f
C206 B.n153 VSUBS 0.006871f
C207 B.n154 VSUBS 0.006871f
C208 B.n155 VSUBS 0.006871f
C209 B.n156 VSUBS 0.006871f
C210 B.n157 VSUBS 0.006871f
C211 B.n158 VSUBS 0.006871f
C212 B.n159 VSUBS 0.006871f
C213 B.n160 VSUBS 0.006871f
C214 B.n161 VSUBS 0.006871f
C215 B.n162 VSUBS 0.006871f
C216 B.n163 VSUBS 0.006871f
C217 B.n164 VSUBS 0.006871f
C218 B.n165 VSUBS 0.006871f
C219 B.n166 VSUBS 0.006871f
C220 B.n167 VSUBS 0.014901f
C221 B.n168 VSUBS 0.006871f
C222 B.n169 VSUBS 0.006871f
C223 B.n170 VSUBS 0.006871f
C224 B.n171 VSUBS 0.006871f
C225 B.n172 VSUBS 0.006871f
C226 B.n173 VSUBS 0.006871f
C227 B.n174 VSUBS 0.006871f
C228 B.n175 VSUBS 0.006871f
C229 B.n176 VSUBS 0.006871f
C230 B.n177 VSUBS 0.006871f
C231 B.n178 VSUBS 0.006871f
C232 B.n179 VSUBS 0.006871f
C233 B.n180 VSUBS 0.006871f
C234 B.n181 VSUBS 0.006871f
C235 B.n182 VSUBS 0.006871f
C236 B.n183 VSUBS 0.006871f
C237 B.n184 VSUBS 0.006871f
C238 B.n185 VSUBS 0.006871f
C239 B.n186 VSUBS 0.006871f
C240 B.n187 VSUBS 0.006871f
C241 B.n188 VSUBS 0.006871f
C242 B.n189 VSUBS 0.006871f
C243 B.n190 VSUBS 0.006871f
C244 B.n191 VSUBS 0.006871f
C245 B.n192 VSUBS 0.006871f
C246 B.n193 VSUBS 0.006871f
C247 B.n194 VSUBS 0.006871f
C248 B.n195 VSUBS 0.006871f
C249 B.n196 VSUBS 0.006871f
C250 B.n197 VSUBS 0.006871f
C251 B.n198 VSUBS 0.006871f
C252 B.n199 VSUBS 0.006871f
C253 B.n200 VSUBS 0.006871f
C254 B.n201 VSUBS 0.006871f
C255 B.n202 VSUBS 0.006871f
C256 B.n203 VSUBS 0.006871f
C257 B.n204 VSUBS 0.006871f
C258 B.n205 VSUBS 0.006871f
C259 B.n206 VSUBS 0.006871f
C260 B.n207 VSUBS 0.006871f
C261 B.n208 VSUBS 0.006871f
C262 B.n209 VSUBS 0.006871f
C263 B.n210 VSUBS 0.006871f
C264 B.n211 VSUBS 0.006871f
C265 B.n212 VSUBS 0.006871f
C266 B.n213 VSUBS 0.006871f
C267 B.n214 VSUBS 0.006871f
C268 B.n215 VSUBS 0.006871f
C269 B.n216 VSUBS 0.014901f
C270 B.n217 VSUBS 0.015814f
C271 B.n218 VSUBS 0.015814f
C272 B.n219 VSUBS 0.006871f
C273 B.n220 VSUBS 0.006871f
C274 B.n221 VSUBS 0.006871f
C275 B.n222 VSUBS 0.006871f
C276 B.n223 VSUBS 0.006871f
C277 B.n224 VSUBS 0.006871f
C278 B.n225 VSUBS 0.006871f
C279 B.n226 VSUBS 0.006871f
C280 B.n227 VSUBS 0.006871f
C281 B.n228 VSUBS 0.006871f
C282 B.n229 VSUBS 0.006871f
C283 B.n230 VSUBS 0.006871f
C284 B.n231 VSUBS 0.006871f
C285 B.n232 VSUBS 0.006871f
C286 B.n233 VSUBS 0.006871f
C287 B.n234 VSUBS 0.006871f
C288 B.n235 VSUBS 0.006871f
C289 B.n236 VSUBS 0.006871f
C290 B.n237 VSUBS 0.006871f
C291 B.n238 VSUBS 0.006871f
C292 B.n239 VSUBS 0.006871f
C293 B.n240 VSUBS 0.006871f
C294 B.n241 VSUBS 0.006871f
C295 B.n242 VSUBS 0.006871f
C296 B.n243 VSUBS 0.006871f
C297 B.n244 VSUBS 0.006871f
C298 B.n245 VSUBS 0.006871f
C299 B.n246 VSUBS 0.006871f
C300 B.n247 VSUBS 0.006871f
C301 B.n248 VSUBS 0.006871f
C302 B.n249 VSUBS 0.006871f
C303 B.n250 VSUBS 0.006871f
C304 B.n251 VSUBS 0.006871f
C305 B.n252 VSUBS 0.006871f
C306 B.n253 VSUBS 0.006871f
C307 B.n254 VSUBS 0.006871f
C308 B.n255 VSUBS 0.006871f
C309 B.n256 VSUBS 0.006871f
C310 B.n257 VSUBS 0.006871f
C311 B.n258 VSUBS 0.006871f
C312 B.n259 VSUBS 0.006871f
C313 B.n260 VSUBS 0.006871f
C314 B.n261 VSUBS 0.006871f
C315 B.n262 VSUBS 0.006871f
C316 B.n263 VSUBS 0.006871f
C317 B.n264 VSUBS 0.006871f
C318 B.n265 VSUBS 0.006871f
C319 B.n266 VSUBS 0.006871f
C320 B.n267 VSUBS 0.006871f
C321 B.n268 VSUBS 0.006871f
C322 B.n269 VSUBS 0.006871f
C323 B.n270 VSUBS 0.006871f
C324 B.n271 VSUBS 0.006871f
C325 B.n272 VSUBS 0.006871f
C326 B.n273 VSUBS 0.006871f
C327 B.n274 VSUBS 0.006871f
C328 B.n275 VSUBS 0.006871f
C329 B.n276 VSUBS 0.006871f
C330 B.n277 VSUBS 0.006871f
C331 B.n278 VSUBS 0.006871f
C332 B.n279 VSUBS 0.006871f
C333 B.n280 VSUBS 0.006871f
C334 B.n281 VSUBS 0.006871f
C335 B.n282 VSUBS 0.006871f
C336 B.n283 VSUBS 0.006871f
C337 B.n284 VSUBS 0.006871f
C338 B.n285 VSUBS 0.006871f
C339 B.n286 VSUBS 0.006871f
C340 B.n287 VSUBS 0.006871f
C341 B.n288 VSUBS 0.006871f
C342 B.n289 VSUBS 0.006871f
C343 B.n290 VSUBS 0.006871f
C344 B.n291 VSUBS 0.006871f
C345 B.n292 VSUBS 0.006871f
C346 B.n293 VSUBS 0.006871f
C347 B.n294 VSUBS 0.006871f
C348 B.n295 VSUBS 0.006871f
C349 B.n296 VSUBS 0.006466f
C350 B.n297 VSUBS 0.015918f
C351 B.n298 VSUBS 0.003839f
C352 B.n299 VSUBS 0.006871f
C353 B.n300 VSUBS 0.006871f
C354 B.n301 VSUBS 0.006871f
C355 B.n302 VSUBS 0.006871f
C356 B.n303 VSUBS 0.006871f
C357 B.n304 VSUBS 0.006871f
C358 B.n305 VSUBS 0.006871f
C359 B.n306 VSUBS 0.006871f
C360 B.n307 VSUBS 0.006871f
C361 B.n308 VSUBS 0.006871f
C362 B.n309 VSUBS 0.006871f
C363 B.n310 VSUBS 0.006871f
C364 B.n311 VSUBS 0.003839f
C365 B.n312 VSUBS 0.006871f
C366 B.n313 VSUBS 0.006871f
C367 B.n314 VSUBS 0.006466f
C368 B.n315 VSUBS 0.006871f
C369 B.n316 VSUBS 0.006871f
C370 B.n317 VSUBS 0.006871f
C371 B.n318 VSUBS 0.006871f
C372 B.n319 VSUBS 0.006871f
C373 B.n320 VSUBS 0.006871f
C374 B.n321 VSUBS 0.006871f
C375 B.n322 VSUBS 0.006871f
C376 B.n323 VSUBS 0.006871f
C377 B.n324 VSUBS 0.006871f
C378 B.n325 VSUBS 0.006871f
C379 B.n326 VSUBS 0.006871f
C380 B.n327 VSUBS 0.006871f
C381 B.n328 VSUBS 0.006871f
C382 B.n329 VSUBS 0.006871f
C383 B.n330 VSUBS 0.006871f
C384 B.n331 VSUBS 0.006871f
C385 B.n332 VSUBS 0.006871f
C386 B.n333 VSUBS 0.006871f
C387 B.n334 VSUBS 0.006871f
C388 B.n335 VSUBS 0.006871f
C389 B.n336 VSUBS 0.006871f
C390 B.n337 VSUBS 0.006871f
C391 B.n338 VSUBS 0.006871f
C392 B.n339 VSUBS 0.006871f
C393 B.n340 VSUBS 0.006871f
C394 B.n341 VSUBS 0.006871f
C395 B.n342 VSUBS 0.006871f
C396 B.n343 VSUBS 0.006871f
C397 B.n344 VSUBS 0.006871f
C398 B.n345 VSUBS 0.006871f
C399 B.n346 VSUBS 0.006871f
C400 B.n347 VSUBS 0.006871f
C401 B.n348 VSUBS 0.006871f
C402 B.n349 VSUBS 0.006871f
C403 B.n350 VSUBS 0.006871f
C404 B.n351 VSUBS 0.006871f
C405 B.n352 VSUBS 0.006871f
C406 B.n353 VSUBS 0.006871f
C407 B.n354 VSUBS 0.006871f
C408 B.n355 VSUBS 0.006871f
C409 B.n356 VSUBS 0.006871f
C410 B.n357 VSUBS 0.006871f
C411 B.n358 VSUBS 0.006871f
C412 B.n359 VSUBS 0.006871f
C413 B.n360 VSUBS 0.006871f
C414 B.n361 VSUBS 0.006871f
C415 B.n362 VSUBS 0.006871f
C416 B.n363 VSUBS 0.006871f
C417 B.n364 VSUBS 0.006871f
C418 B.n365 VSUBS 0.006871f
C419 B.n366 VSUBS 0.006871f
C420 B.n367 VSUBS 0.006871f
C421 B.n368 VSUBS 0.006871f
C422 B.n369 VSUBS 0.006871f
C423 B.n370 VSUBS 0.006871f
C424 B.n371 VSUBS 0.006871f
C425 B.n372 VSUBS 0.006871f
C426 B.n373 VSUBS 0.006871f
C427 B.n374 VSUBS 0.006871f
C428 B.n375 VSUBS 0.006871f
C429 B.n376 VSUBS 0.006871f
C430 B.n377 VSUBS 0.006871f
C431 B.n378 VSUBS 0.006871f
C432 B.n379 VSUBS 0.006871f
C433 B.n380 VSUBS 0.006871f
C434 B.n381 VSUBS 0.006871f
C435 B.n382 VSUBS 0.006871f
C436 B.n383 VSUBS 0.006871f
C437 B.n384 VSUBS 0.006871f
C438 B.n385 VSUBS 0.006871f
C439 B.n386 VSUBS 0.006871f
C440 B.n387 VSUBS 0.006871f
C441 B.n388 VSUBS 0.006871f
C442 B.n389 VSUBS 0.006871f
C443 B.n390 VSUBS 0.006871f
C444 B.n391 VSUBS 0.015814f
C445 B.n392 VSUBS 0.015814f
C446 B.n393 VSUBS 0.014901f
C447 B.n394 VSUBS 0.006871f
C448 B.n395 VSUBS 0.006871f
C449 B.n396 VSUBS 0.006871f
C450 B.n397 VSUBS 0.006871f
C451 B.n398 VSUBS 0.006871f
C452 B.n399 VSUBS 0.006871f
C453 B.n400 VSUBS 0.006871f
C454 B.n401 VSUBS 0.006871f
C455 B.n402 VSUBS 0.006871f
C456 B.n403 VSUBS 0.006871f
C457 B.n404 VSUBS 0.006871f
C458 B.n405 VSUBS 0.006871f
C459 B.n406 VSUBS 0.006871f
C460 B.n407 VSUBS 0.006871f
C461 B.n408 VSUBS 0.006871f
C462 B.n409 VSUBS 0.006871f
C463 B.n410 VSUBS 0.006871f
C464 B.n411 VSUBS 0.006871f
C465 B.n412 VSUBS 0.006871f
C466 B.n413 VSUBS 0.006871f
C467 B.n414 VSUBS 0.006871f
C468 B.n415 VSUBS 0.006871f
C469 B.n416 VSUBS 0.006871f
C470 B.n417 VSUBS 0.006871f
C471 B.n418 VSUBS 0.006871f
C472 B.n419 VSUBS 0.006871f
C473 B.n420 VSUBS 0.006871f
C474 B.n421 VSUBS 0.006871f
C475 B.n422 VSUBS 0.006871f
C476 B.n423 VSUBS 0.006871f
C477 B.n424 VSUBS 0.006871f
C478 B.n425 VSUBS 0.006871f
C479 B.n426 VSUBS 0.006871f
C480 B.n427 VSUBS 0.006871f
C481 B.n428 VSUBS 0.006871f
C482 B.n429 VSUBS 0.006871f
C483 B.n430 VSUBS 0.006871f
C484 B.n431 VSUBS 0.006871f
C485 B.n432 VSUBS 0.006871f
C486 B.n433 VSUBS 0.006871f
C487 B.n434 VSUBS 0.006871f
C488 B.n435 VSUBS 0.006871f
C489 B.n436 VSUBS 0.006871f
C490 B.n437 VSUBS 0.006871f
C491 B.n438 VSUBS 0.006871f
C492 B.n439 VSUBS 0.006871f
C493 B.n440 VSUBS 0.006871f
C494 B.n441 VSUBS 0.006871f
C495 B.n442 VSUBS 0.006871f
C496 B.n443 VSUBS 0.006871f
C497 B.n444 VSUBS 0.006871f
C498 B.n445 VSUBS 0.006871f
C499 B.n446 VSUBS 0.006871f
C500 B.n447 VSUBS 0.006871f
C501 B.n448 VSUBS 0.006871f
C502 B.n449 VSUBS 0.006871f
C503 B.n450 VSUBS 0.006871f
C504 B.n451 VSUBS 0.006871f
C505 B.n452 VSUBS 0.006871f
C506 B.n453 VSUBS 0.006871f
C507 B.n454 VSUBS 0.006871f
C508 B.n455 VSUBS 0.006871f
C509 B.n456 VSUBS 0.006871f
C510 B.n457 VSUBS 0.006871f
C511 B.n458 VSUBS 0.006871f
C512 B.n459 VSUBS 0.006871f
C513 B.n460 VSUBS 0.006871f
C514 B.n461 VSUBS 0.006871f
C515 B.n462 VSUBS 0.006871f
C516 B.n463 VSUBS 0.006871f
C517 B.n464 VSUBS 0.006871f
C518 B.n465 VSUBS 0.006871f
C519 B.n466 VSUBS 0.006871f
C520 B.n467 VSUBS 0.006871f
C521 B.n468 VSUBS 0.006871f
C522 B.n469 VSUBS 0.006871f
C523 B.n470 VSUBS 0.006871f
C524 B.n471 VSUBS 0.015772f
C525 B.n472 VSUBS 0.014943f
C526 B.n473 VSUBS 0.015814f
C527 B.n474 VSUBS 0.006871f
C528 B.n475 VSUBS 0.006871f
C529 B.n476 VSUBS 0.006871f
C530 B.n477 VSUBS 0.006871f
C531 B.n478 VSUBS 0.006871f
C532 B.n479 VSUBS 0.006871f
C533 B.n480 VSUBS 0.006871f
C534 B.n481 VSUBS 0.006871f
C535 B.n482 VSUBS 0.006871f
C536 B.n483 VSUBS 0.006871f
C537 B.n484 VSUBS 0.006871f
C538 B.n485 VSUBS 0.006871f
C539 B.n486 VSUBS 0.006871f
C540 B.n487 VSUBS 0.006871f
C541 B.n488 VSUBS 0.006871f
C542 B.n489 VSUBS 0.006871f
C543 B.n490 VSUBS 0.006871f
C544 B.n491 VSUBS 0.006871f
C545 B.n492 VSUBS 0.006871f
C546 B.n493 VSUBS 0.006871f
C547 B.n494 VSUBS 0.006871f
C548 B.n495 VSUBS 0.006871f
C549 B.n496 VSUBS 0.006871f
C550 B.n497 VSUBS 0.006871f
C551 B.n498 VSUBS 0.006871f
C552 B.n499 VSUBS 0.006871f
C553 B.n500 VSUBS 0.006871f
C554 B.n501 VSUBS 0.006871f
C555 B.n502 VSUBS 0.006871f
C556 B.n503 VSUBS 0.006871f
C557 B.n504 VSUBS 0.006871f
C558 B.n505 VSUBS 0.006871f
C559 B.n506 VSUBS 0.006871f
C560 B.n507 VSUBS 0.006871f
C561 B.n508 VSUBS 0.006871f
C562 B.n509 VSUBS 0.006871f
C563 B.n510 VSUBS 0.006871f
C564 B.n511 VSUBS 0.006871f
C565 B.n512 VSUBS 0.006871f
C566 B.n513 VSUBS 0.006871f
C567 B.n514 VSUBS 0.006871f
C568 B.n515 VSUBS 0.006871f
C569 B.n516 VSUBS 0.006871f
C570 B.n517 VSUBS 0.006871f
C571 B.n518 VSUBS 0.006871f
C572 B.n519 VSUBS 0.006871f
C573 B.n520 VSUBS 0.006871f
C574 B.n521 VSUBS 0.006871f
C575 B.n522 VSUBS 0.006871f
C576 B.n523 VSUBS 0.006871f
C577 B.n524 VSUBS 0.006871f
C578 B.n525 VSUBS 0.006871f
C579 B.n526 VSUBS 0.006871f
C580 B.n527 VSUBS 0.006871f
C581 B.n528 VSUBS 0.006871f
C582 B.n529 VSUBS 0.006871f
C583 B.n530 VSUBS 0.006871f
C584 B.n531 VSUBS 0.006871f
C585 B.n532 VSUBS 0.006871f
C586 B.n533 VSUBS 0.006871f
C587 B.n534 VSUBS 0.006871f
C588 B.n535 VSUBS 0.006871f
C589 B.n536 VSUBS 0.006871f
C590 B.n537 VSUBS 0.006871f
C591 B.n538 VSUBS 0.006871f
C592 B.n539 VSUBS 0.006871f
C593 B.n540 VSUBS 0.006871f
C594 B.n541 VSUBS 0.006871f
C595 B.n542 VSUBS 0.006871f
C596 B.n543 VSUBS 0.006871f
C597 B.n544 VSUBS 0.006871f
C598 B.n545 VSUBS 0.006871f
C599 B.n546 VSUBS 0.006871f
C600 B.n547 VSUBS 0.006871f
C601 B.n548 VSUBS 0.006871f
C602 B.n549 VSUBS 0.006871f
C603 B.n550 VSUBS 0.006466f
C604 B.n551 VSUBS 0.006871f
C605 B.n552 VSUBS 0.006871f
C606 B.n553 VSUBS 0.006871f
C607 B.n554 VSUBS 0.006871f
C608 B.n555 VSUBS 0.006871f
C609 B.n556 VSUBS 0.006871f
C610 B.n557 VSUBS 0.006871f
C611 B.n558 VSUBS 0.006871f
C612 B.n559 VSUBS 0.006871f
C613 B.n560 VSUBS 0.006871f
C614 B.n561 VSUBS 0.006871f
C615 B.n562 VSUBS 0.006871f
C616 B.n563 VSUBS 0.006871f
C617 B.n564 VSUBS 0.006871f
C618 B.n565 VSUBS 0.006871f
C619 B.n566 VSUBS 0.003839f
C620 B.n567 VSUBS 0.015918f
C621 B.n568 VSUBS 0.006466f
C622 B.n569 VSUBS 0.006871f
C623 B.n570 VSUBS 0.006871f
C624 B.n571 VSUBS 0.006871f
C625 B.n572 VSUBS 0.006871f
C626 B.n573 VSUBS 0.006871f
C627 B.n574 VSUBS 0.006871f
C628 B.n575 VSUBS 0.006871f
C629 B.n576 VSUBS 0.006871f
C630 B.n577 VSUBS 0.006871f
C631 B.n578 VSUBS 0.006871f
C632 B.n579 VSUBS 0.006871f
C633 B.n580 VSUBS 0.006871f
C634 B.n581 VSUBS 0.006871f
C635 B.n582 VSUBS 0.006871f
C636 B.n583 VSUBS 0.006871f
C637 B.n584 VSUBS 0.006871f
C638 B.n585 VSUBS 0.006871f
C639 B.n586 VSUBS 0.006871f
C640 B.n587 VSUBS 0.006871f
C641 B.n588 VSUBS 0.006871f
C642 B.n589 VSUBS 0.006871f
C643 B.n590 VSUBS 0.006871f
C644 B.n591 VSUBS 0.006871f
C645 B.n592 VSUBS 0.006871f
C646 B.n593 VSUBS 0.006871f
C647 B.n594 VSUBS 0.006871f
C648 B.n595 VSUBS 0.006871f
C649 B.n596 VSUBS 0.006871f
C650 B.n597 VSUBS 0.006871f
C651 B.n598 VSUBS 0.006871f
C652 B.n599 VSUBS 0.006871f
C653 B.n600 VSUBS 0.006871f
C654 B.n601 VSUBS 0.006871f
C655 B.n602 VSUBS 0.006871f
C656 B.n603 VSUBS 0.006871f
C657 B.n604 VSUBS 0.006871f
C658 B.n605 VSUBS 0.006871f
C659 B.n606 VSUBS 0.006871f
C660 B.n607 VSUBS 0.006871f
C661 B.n608 VSUBS 0.006871f
C662 B.n609 VSUBS 0.006871f
C663 B.n610 VSUBS 0.006871f
C664 B.n611 VSUBS 0.006871f
C665 B.n612 VSUBS 0.006871f
C666 B.n613 VSUBS 0.006871f
C667 B.n614 VSUBS 0.006871f
C668 B.n615 VSUBS 0.006871f
C669 B.n616 VSUBS 0.006871f
C670 B.n617 VSUBS 0.006871f
C671 B.n618 VSUBS 0.006871f
C672 B.n619 VSUBS 0.006871f
C673 B.n620 VSUBS 0.006871f
C674 B.n621 VSUBS 0.006871f
C675 B.n622 VSUBS 0.006871f
C676 B.n623 VSUBS 0.006871f
C677 B.n624 VSUBS 0.006871f
C678 B.n625 VSUBS 0.006871f
C679 B.n626 VSUBS 0.006871f
C680 B.n627 VSUBS 0.006871f
C681 B.n628 VSUBS 0.006871f
C682 B.n629 VSUBS 0.006871f
C683 B.n630 VSUBS 0.006871f
C684 B.n631 VSUBS 0.006871f
C685 B.n632 VSUBS 0.006871f
C686 B.n633 VSUBS 0.006871f
C687 B.n634 VSUBS 0.006871f
C688 B.n635 VSUBS 0.006871f
C689 B.n636 VSUBS 0.006871f
C690 B.n637 VSUBS 0.006871f
C691 B.n638 VSUBS 0.006871f
C692 B.n639 VSUBS 0.006871f
C693 B.n640 VSUBS 0.006871f
C694 B.n641 VSUBS 0.006871f
C695 B.n642 VSUBS 0.006871f
C696 B.n643 VSUBS 0.006871f
C697 B.n644 VSUBS 0.006871f
C698 B.n645 VSUBS 0.006871f
C699 B.n646 VSUBS 0.015814f
C700 B.n647 VSUBS 0.014901f
C701 B.n648 VSUBS 0.014901f
C702 B.n649 VSUBS 0.006871f
C703 B.n650 VSUBS 0.006871f
C704 B.n651 VSUBS 0.006871f
C705 B.n652 VSUBS 0.006871f
C706 B.n653 VSUBS 0.006871f
C707 B.n654 VSUBS 0.006871f
C708 B.n655 VSUBS 0.006871f
C709 B.n656 VSUBS 0.006871f
C710 B.n657 VSUBS 0.006871f
C711 B.n658 VSUBS 0.006871f
C712 B.n659 VSUBS 0.006871f
C713 B.n660 VSUBS 0.006871f
C714 B.n661 VSUBS 0.006871f
C715 B.n662 VSUBS 0.006871f
C716 B.n663 VSUBS 0.006871f
C717 B.n664 VSUBS 0.006871f
C718 B.n665 VSUBS 0.006871f
C719 B.n666 VSUBS 0.006871f
C720 B.n667 VSUBS 0.006871f
C721 B.n668 VSUBS 0.006871f
C722 B.n669 VSUBS 0.006871f
C723 B.n670 VSUBS 0.006871f
C724 B.n671 VSUBS 0.006871f
C725 B.n672 VSUBS 0.006871f
C726 B.n673 VSUBS 0.006871f
C727 B.n674 VSUBS 0.006871f
C728 B.n675 VSUBS 0.006871f
C729 B.n676 VSUBS 0.006871f
C730 B.n677 VSUBS 0.006871f
C731 B.n678 VSUBS 0.006871f
C732 B.n679 VSUBS 0.006871f
C733 B.n680 VSUBS 0.006871f
C734 B.n681 VSUBS 0.006871f
C735 B.n682 VSUBS 0.006871f
C736 B.n683 VSUBS 0.006871f
C737 B.n684 VSUBS 0.006871f
C738 B.n685 VSUBS 0.006871f
C739 B.n686 VSUBS 0.006871f
C740 B.n687 VSUBS 0.015557f
C741 VTAIL.t1 VSUBS 2.84968f
C742 VTAIL.n0 VSUBS 0.703232f
C743 VTAIL.t4 VSUBS 2.84968f
C744 VTAIL.n1 VSUBS 0.761545f
C745 VTAIL.t6 VSUBS 2.84968f
C746 VTAIL.n2 VSUBS 2.1391f
C747 VTAIL.t2 VSUBS 2.8497f
C748 VTAIL.n3 VSUBS 2.13908f
C749 VTAIL.t3 VSUBS 2.8497f
C750 VTAIL.n4 VSUBS 0.761524f
C751 VTAIL.t7 VSUBS 2.8497f
C752 VTAIL.n5 VSUBS 0.761524f
C753 VTAIL.t5 VSUBS 2.84968f
C754 VTAIL.n6 VSUBS 2.1391f
C755 VTAIL.t0 VSUBS 2.84968f
C756 VTAIL.n7 VSUBS 2.07243f
C757 VDD1.t2 VSUBS 0.335638f
C758 VDD1.t0 VSUBS 0.335638f
C759 VDD1.n0 VSUBS 2.75965f
C760 VDD1.t1 VSUBS 0.335638f
C761 VDD1.t3 VSUBS 0.335638f
C762 VDD1.n1 VSUBS 3.57364f
C763 VP.n0 VSUBS 0.040109f
C764 VP.t3 VSUBS 2.95705f
C765 VP.n1 VSUBS 0.032394f
C766 VP.n2 VSUBS 0.040109f
C767 VP.t1 VSUBS 2.95705f
C768 VP.t0 VSUBS 3.12096f
C769 VP.t2 VSUBS 3.11895f
C770 VP.n3 VSUBS 4.01933f
C771 VP.n4 VSUBS 2.35947f
C772 VP.n5 VSUBS 1.121f
C773 VP.n6 VSUBS 0.038394f
C774 VP.n7 VSUBS 0.079296f
C775 VP.n8 VSUBS 0.040109f
C776 VP.n9 VSUBS 0.040109f
C777 VP.n10 VSUBS 0.040109f
C778 VP.n11 VSUBS 0.079296f
C779 VP.n12 VSUBS 0.038394f
C780 VP.n13 VSUBS 1.121f
C781 VP.n14 VSUBS 0.04266f
.ends

