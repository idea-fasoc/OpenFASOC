* NGSPICE file created from diff_pair_sample_0506.ext - technology: sky130A

.subckt diff_pair_sample_0506 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=1.7238 ps=9.62 w=4.42 l=0.21
X1 B.t11 B.t9 B.t10 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=0 ps=0 w=4.42 l=0.21
X2 B.t8 B.t6 B.t7 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=0 ps=0 w=4.42 l=0.21
X3 B.t5 B.t3 B.t4 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=0 ps=0 w=4.42 l=0.21
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=1.7238 ps=9.62 w=4.42 l=0.21
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=1.7238 ps=9.62 w=4.42 l=0.21
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=1.7238 ps=9.62 w=4.42 l=0.21
X7 B.t2 B.t0 B.t1 w_n1186_n1856# sky130_fd_pr__pfet_01v8 ad=1.7238 pd=9.62 as=0 ps=0 w=4.42 l=0.21
R0 VP.n0 VP.t0 874.429
R1 VP.n0 VP.t1 841.838
R2 VP VP.n0 0.0516364
R3 VTAIL.n1 VTAIL.t0 103.329
R4 VTAIL.n3 VTAIL.t1 103.329
R5 VTAIL.n0 VTAIL.t2 103.329
R6 VTAIL.n2 VTAIL.t3 103.329
R7 VTAIL.n1 VTAIL.n0 17.1255
R8 VTAIL.n3 VTAIL.n2 16.66
R9 VTAIL.n2 VTAIL.n1 0.703086
R10 VTAIL VTAIL.n0 0.644897
R11 VTAIL VTAIL.n3 0.0586897
R12 VDD1 VDD1.t0 149.066
R13 VDD1 VDD1.t1 120.181
R14 B.n58 B.t9 740.73
R15 B.n64 B.t3 740.73
R16 B.n18 B.t0 740.73
R17 B.n24 B.t6 740.73
R18 B.n205 B.n204 585
R19 B.n206 B.n35 585
R20 B.n208 B.n207 585
R21 B.n209 B.n34 585
R22 B.n211 B.n210 585
R23 B.n212 B.n33 585
R24 B.n214 B.n213 585
R25 B.n215 B.n32 585
R26 B.n217 B.n216 585
R27 B.n218 B.n31 585
R28 B.n220 B.n219 585
R29 B.n221 B.n30 585
R30 B.n223 B.n222 585
R31 B.n224 B.n29 585
R32 B.n226 B.n225 585
R33 B.n227 B.n28 585
R34 B.n229 B.n228 585
R35 B.n230 B.n27 585
R36 B.n232 B.n231 585
R37 B.n234 B.n233 585
R38 B.n235 B.n23 585
R39 B.n237 B.n236 585
R40 B.n238 B.n22 585
R41 B.n240 B.n239 585
R42 B.n241 B.n21 585
R43 B.n243 B.n242 585
R44 B.n244 B.n20 585
R45 B.n246 B.n245 585
R46 B.n247 B.n17 585
R47 B.n250 B.n249 585
R48 B.n251 B.n16 585
R49 B.n253 B.n252 585
R50 B.n254 B.n15 585
R51 B.n256 B.n255 585
R52 B.n257 B.n14 585
R53 B.n259 B.n258 585
R54 B.n260 B.n13 585
R55 B.n262 B.n261 585
R56 B.n263 B.n12 585
R57 B.n265 B.n264 585
R58 B.n266 B.n11 585
R59 B.n268 B.n267 585
R60 B.n269 B.n10 585
R61 B.n271 B.n270 585
R62 B.n272 B.n9 585
R63 B.n274 B.n273 585
R64 B.n275 B.n8 585
R65 B.n277 B.n276 585
R66 B.n203 B.n36 585
R67 B.n202 B.n201 585
R68 B.n200 B.n37 585
R69 B.n199 B.n198 585
R70 B.n197 B.n38 585
R71 B.n196 B.n195 585
R72 B.n194 B.n39 585
R73 B.n193 B.n192 585
R74 B.n191 B.n40 585
R75 B.n190 B.n189 585
R76 B.n188 B.n41 585
R77 B.n187 B.n186 585
R78 B.n185 B.n42 585
R79 B.n184 B.n183 585
R80 B.n182 B.n43 585
R81 B.n181 B.n180 585
R82 B.n179 B.n44 585
R83 B.n178 B.n177 585
R84 B.n176 B.n45 585
R85 B.n175 B.n174 585
R86 B.n173 B.n46 585
R87 B.n172 B.n171 585
R88 B.n170 B.n47 585
R89 B.n97 B.n96 585
R90 B.n98 B.n75 585
R91 B.n100 B.n99 585
R92 B.n101 B.n74 585
R93 B.n103 B.n102 585
R94 B.n104 B.n73 585
R95 B.n106 B.n105 585
R96 B.n107 B.n72 585
R97 B.n109 B.n108 585
R98 B.n110 B.n71 585
R99 B.n112 B.n111 585
R100 B.n113 B.n70 585
R101 B.n115 B.n114 585
R102 B.n116 B.n69 585
R103 B.n118 B.n117 585
R104 B.n119 B.n68 585
R105 B.n121 B.n120 585
R106 B.n122 B.n67 585
R107 B.n124 B.n123 585
R108 B.n126 B.n125 585
R109 B.n127 B.n63 585
R110 B.n129 B.n128 585
R111 B.n130 B.n62 585
R112 B.n132 B.n131 585
R113 B.n133 B.n61 585
R114 B.n135 B.n134 585
R115 B.n136 B.n60 585
R116 B.n138 B.n137 585
R117 B.n139 B.n57 585
R118 B.n142 B.n141 585
R119 B.n143 B.n56 585
R120 B.n145 B.n144 585
R121 B.n146 B.n55 585
R122 B.n148 B.n147 585
R123 B.n149 B.n54 585
R124 B.n151 B.n150 585
R125 B.n152 B.n53 585
R126 B.n154 B.n153 585
R127 B.n155 B.n52 585
R128 B.n157 B.n156 585
R129 B.n158 B.n51 585
R130 B.n160 B.n159 585
R131 B.n161 B.n50 585
R132 B.n163 B.n162 585
R133 B.n164 B.n49 585
R134 B.n166 B.n165 585
R135 B.n167 B.n48 585
R136 B.n169 B.n168 585
R137 B.n95 B.n76 585
R138 B.n94 B.n93 585
R139 B.n92 B.n77 585
R140 B.n91 B.n90 585
R141 B.n89 B.n78 585
R142 B.n88 B.n87 585
R143 B.n86 B.n79 585
R144 B.n85 B.n84 585
R145 B.n83 B.n80 585
R146 B.n82 B.n81 585
R147 B.n2 B.n0 585
R148 B.n293 B.n1 585
R149 B.n292 B.n291 585
R150 B.n290 B.n3 585
R151 B.n289 B.n288 585
R152 B.n287 B.n4 585
R153 B.n286 B.n285 585
R154 B.n284 B.n5 585
R155 B.n283 B.n282 585
R156 B.n281 B.n6 585
R157 B.n280 B.n279 585
R158 B.n278 B.n7 585
R159 B.n295 B.n294 585
R160 B.n96 B.n95 574.183
R161 B.n276 B.n7 574.183
R162 B.n168 B.n47 574.183
R163 B.n204 B.n203 574.183
R164 B.n95 B.n94 163.367
R165 B.n94 B.n77 163.367
R166 B.n90 B.n77 163.367
R167 B.n90 B.n89 163.367
R168 B.n89 B.n88 163.367
R169 B.n88 B.n79 163.367
R170 B.n84 B.n79 163.367
R171 B.n84 B.n83 163.367
R172 B.n83 B.n82 163.367
R173 B.n82 B.n2 163.367
R174 B.n294 B.n2 163.367
R175 B.n294 B.n293 163.367
R176 B.n293 B.n292 163.367
R177 B.n292 B.n3 163.367
R178 B.n288 B.n3 163.367
R179 B.n288 B.n287 163.367
R180 B.n287 B.n286 163.367
R181 B.n286 B.n5 163.367
R182 B.n282 B.n5 163.367
R183 B.n282 B.n281 163.367
R184 B.n281 B.n280 163.367
R185 B.n280 B.n7 163.367
R186 B.n96 B.n75 163.367
R187 B.n100 B.n75 163.367
R188 B.n101 B.n100 163.367
R189 B.n102 B.n101 163.367
R190 B.n102 B.n73 163.367
R191 B.n106 B.n73 163.367
R192 B.n107 B.n106 163.367
R193 B.n108 B.n107 163.367
R194 B.n108 B.n71 163.367
R195 B.n112 B.n71 163.367
R196 B.n113 B.n112 163.367
R197 B.n114 B.n113 163.367
R198 B.n114 B.n69 163.367
R199 B.n118 B.n69 163.367
R200 B.n119 B.n118 163.367
R201 B.n120 B.n119 163.367
R202 B.n120 B.n67 163.367
R203 B.n124 B.n67 163.367
R204 B.n125 B.n124 163.367
R205 B.n125 B.n63 163.367
R206 B.n129 B.n63 163.367
R207 B.n130 B.n129 163.367
R208 B.n131 B.n130 163.367
R209 B.n131 B.n61 163.367
R210 B.n135 B.n61 163.367
R211 B.n136 B.n135 163.367
R212 B.n137 B.n136 163.367
R213 B.n137 B.n57 163.367
R214 B.n142 B.n57 163.367
R215 B.n143 B.n142 163.367
R216 B.n144 B.n143 163.367
R217 B.n144 B.n55 163.367
R218 B.n148 B.n55 163.367
R219 B.n149 B.n148 163.367
R220 B.n150 B.n149 163.367
R221 B.n150 B.n53 163.367
R222 B.n154 B.n53 163.367
R223 B.n155 B.n154 163.367
R224 B.n156 B.n155 163.367
R225 B.n156 B.n51 163.367
R226 B.n160 B.n51 163.367
R227 B.n161 B.n160 163.367
R228 B.n162 B.n161 163.367
R229 B.n162 B.n49 163.367
R230 B.n166 B.n49 163.367
R231 B.n167 B.n166 163.367
R232 B.n168 B.n167 163.367
R233 B.n172 B.n47 163.367
R234 B.n173 B.n172 163.367
R235 B.n174 B.n173 163.367
R236 B.n174 B.n45 163.367
R237 B.n178 B.n45 163.367
R238 B.n179 B.n178 163.367
R239 B.n180 B.n179 163.367
R240 B.n180 B.n43 163.367
R241 B.n184 B.n43 163.367
R242 B.n185 B.n184 163.367
R243 B.n186 B.n185 163.367
R244 B.n186 B.n41 163.367
R245 B.n190 B.n41 163.367
R246 B.n191 B.n190 163.367
R247 B.n192 B.n191 163.367
R248 B.n192 B.n39 163.367
R249 B.n196 B.n39 163.367
R250 B.n197 B.n196 163.367
R251 B.n198 B.n197 163.367
R252 B.n198 B.n37 163.367
R253 B.n202 B.n37 163.367
R254 B.n203 B.n202 163.367
R255 B.n276 B.n275 163.367
R256 B.n275 B.n274 163.367
R257 B.n274 B.n9 163.367
R258 B.n270 B.n9 163.367
R259 B.n270 B.n269 163.367
R260 B.n269 B.n268 163.367
R261 B.n268 B.n11 163.367
R262 B.n264 B.n11 163.367
R263 B.n264 B.n263 163.367
R264 B.n263 B.n262 163.367
R265 B.n262 B.n13 163.367
R266 B.n258 B.n13 163.367
R267 B.n258 B.n257 163.367
R268 B.n257 B.n256 163.367
R269 B.n256 B.n15 163.367
R270 B.n252 B.n15 163.367
R271 B.n252 B.n251 163.367
R272 B.n251 B.n250 163.367
R273 B.n250 B.n17 163.367
R274 B.n245 B.n17 163.367
R275 B.n245 B.n244 163.367
R276 B.n244 B.n243 163.367
R277 B.n243 B.n21 163.367
R278 B.n239 B.n21 163.367
R279 B.n239 B.n238 163.367
R280 B.n238 B.n237 163.367
R281 B.n237 B.n23 163.367
R282 B.n233 B.n23 163.367
R283 B.n233 B.n232 163.367
R284 B.n232 B.n27 163.367
R285 B.n228 B.n27 163.367
R286 B.n228 B.n227 163.367
R287 B.n227 B.n226 163.367
R288 B.n226 B.n29 163.367
R289 B.n222 B.n29 163.367
R290 B.n222 B.n221 163.367
R291 B.n221 B.n220 163.367
R292 B.n220 B.n31 163.367
R293 B.n216 B.n31 163.367
R294 B.n216 B.n215 163.367
R295 B.n215 B.n214 163.367
R296 B.n214 B.n33 163.367
R297 B.n210 B.n33 163.367
R298 B.n210 B.n209 163.367
R299 B.n209 B.n208 163.367
R300 B.n208 B.n35 163.367
R301 B.n204 B.n35 163.367
R302 B.n58 B.t11 135.544
R303 B.n24 B.t7 135.544
R304 B.n64 B.t5 135.542
R305 B.n18 B.t1 135.542
R306 B.n59 B.t10 125.073
R307 B.n25 B.t8 125.073
R308 B.n65 B.t4 125.069
R309 B.n19 B.t2 125.069
R310 B.n140 B.n59 59.5399
R311 B.n66 B.n65 59.5399
R312 B.n248 B.n19 59.5399
R313 B.n26 B.n25 59.5399
R314 B.n278 B.n277 37.3078
R315 B.n205 B.n36 37.3078
R316 B.n170 B.n169 37.3078
R317 B.n97 B.n76 37.3078
R318 B B.n295 18.0485
R319 B.n277 B.n8 10.6151
R320 B.n273 B.n8 10.6151
R321 B.n273 B.n272 10.6151
R322 B.n272 B.n271 10.6151
R323 B.n271 B.n10 10.6151
R324 B.n267 B.n10 10.6151
R325 B.n267 B.n266 10.6151
R326 B.n266 B.n265 10.6151
R327 B.n265 B.n12 10.6151
R328 B.n261 B.n12 10.6151
R329 B.n261 B.n260 10.6151
R330 B.n260 B.n259 10.6151
R331 B.n259 B.n14 10.6151
R332 B.n255 B.n14 10.6151
R333 B.n255 B.n254 10.6151
R334 B.n254 B.n253 10.6151
R335 B.n253 B.n16 10.6151
R336 B.n249 B.n16 10.6151
R337 B.n247 B.n246 10.6151
R338 B.n246 B.n20 10.6151
R339 B.n242 B.n20 10.6151
R340 B.n242 B.n241 10.6151
R341 B.n241 B.n240 10.6151
R342 B.n240 B.n22 10.6151
R343 B.n236 B.n22 10.6151
R344 B.n236 B.n235 10.6151
R345 B.n235 B.n234 10.6151
R346 B.n231 B.n230 10.6151
R347 B.n230 B.n229 10.6151
R348 B.n229 B.n28 10.6151
R349 B.n225 B.n28 10.6151
R350 B.n225 B.n224 10.6151
R351 B.n224 B.n223 10.6151
R352 B.n223 B.n30 10.6151
R353 B.n219 B.n30 10.6151
R354 B.n219 B.n218 10.6151
R355 B.n218 B.n217 10.6151
R356 B.n217 B.n32 10.6151
R357 B.n213 B.n32 10.6151
R358 B.n213 B.n212 10.6151
R359 B.n212 B.n211 10.6151
R360 B.n211 B.n34 10.6151
R361 B.n207 B.n34 10.6151
R362 B.n207 B.n206 10.6151
R363 B.n206 B.n205 10.6151
R364 B.n171 B.n170 10.6151
R365 B.n171 B.n46 10.6151
R366 B.n175 B.n46 10.6151
R367 B.n176 B.n175 10.6151
R368 B.n177 B.n176 10.6151
R369 B.n177 B.n44 10.6151
R370 B.n181 B.n44 10.6151
R371 B.n182 B.n181 10.6151
R372 B.n183 B.n182 10.6151
R373 B.n183 B.n42 10.6151
R374 B.n187 B.n42 10.6151
R375 B.n188 B.n187 10.6151
R376 B.n189 B.n188 10.6151
R377 B.n189 B.n40 10.6151
R378 B.n193 B.n40 10.6151
R379 B.n194 B.n193 10.6151
R380 B.n195 B.n194 10.6151
R381 B.n195 B.n38 10.6151
R382 B.n199 B.n38 10.6151
R383 B.n200 B.n199 10.6151
R384 B.n201 B.n200 10.6151
R385 B.n201 B.n36 10.6151
R386 B.n98 B.n97 10.6151
R387 B.n99 B.n98 10.6151
R388 B.n99 B.n74 10.6151
R389 B.n103 B.n74 10.6151
R390 B.n104 B.n103 10.6151
R391 B.n105 B.n104 10.6151
R392 B.n105 B.n72 10.6151
R393 B.n109 B.n72 10.6151
R394 B.n110 B.n109 10.6151
R395 B.n111 B.n110 10.6151
R396 B.n111 B.n70 10.6151
R397 B.n115 B.n70 10.6151
R398 B.n116 B.n115 10.6151
R399 B.n117 B.n116 10.6151
R400 B.n117 B.n68 10.6151
R401 B.n121 B.n68 10.6151
R402 B.n122 B.n121 10.6151
R403 B.n123 B.n122 10.6151
R404 B.n127 B.n126 10.6151
R405 B.n128 B.n127 10.6151
R406 B.n128 B.n62 10.6151
R407 B.n132 B.n62 10.6151
R408 B.n133 B.n132 10.6151
R409 B.n134 B.n133 10.6151
R410 B.n134 B.n60 10.6151
R411 B.n138 B.n60 10.6151
R412 B.n139 B.n138 10.6151
R413 B.n141 B.n56 10.6151
R414 B.n145 B.n56 10.6151
R415 B.n146 B.n145 10.6151
R416 B.n147 B.n146 10.6151
R417 B.n147 B.n54 10.6151
R418 B.n151 B.n54 10.6151
R419 B.n152 B.n151 10.6151
R420 B.n153 B.n152 10.6151
R421 B.n153 B.n52 10.6151
R422 B.n157 B.n52 10.6151
R423 B.n158 B.n157 10.6151
R424 B.n159 B.n158 10.6151
R425 B.n159 B.n50 10.6151
R426 B.n163 B.n50 10.6151
R427 B.n164 B.n163 10.6151
R428 B.n165 B.n164 10.6151
R429 B.n165 B.n48 10.6151
R430 B.n169 B.n48 10.6151
R431 B.n93 B.n76 10.6151
R432 B.n93 B.n92 10.6151
R433 B.n92 B.n91 10.6151
R434 B.n91 B.n78 10.6151
R435 B.n87 B.n78 10.6151
R436 B.n87 B.n86 10.6151
R437 B.n86 B.n85 10.6151
R438 B.n85 B.n80 10.6151
R439 B.n81 B.n80 10.6151
R440 B.n81 B.n0 10.6151
R441 B.n291 B.n1 10.6151
R442 B.n291 B.n290 10.6151
R443 B.n290 B.n289 10.6151
R444 B.n289 B.n4 10.6151
R445 B.n285 B.n4 10.6151
R446 B.n285 B.n284 10.6151
R447 B.n284 B.n283 10.6151
R448 B.n283 B.n6 10.6151
R449 B.n279 B.n6 10.6151
R450 B.n279 B.n278 10.6151
R451 B.n59 B.n58 10.4732
R452 B.n65 B.n64 10.4732
R453 B.n19 B.n18 10.4732
R454 B.n25 B.n24 10.4732
R455 B.n249 B.n248 8.74196
R456 B.n231 B.n26 8.74196
R457 B.n123 B.n66 8.74196
R458 B.n141 B.n140 8.74196
R459 B.n295 B.n0 2.81026
R460 B.n295 B.n1 2.81026
R461 B.n248 B.n247 1.87367
R462 B.n234 B.n26 1.87367
R463 B.n126 B.n66 1.87367
R464 B.n140 B.n139 1.87367
R465 VN VN.t1 874.811
R466 VN VN.t0 841.889
R467 VDD2.n0 VDD2.t1 148.425
R468 VDD2.n0 VDD2.t0 120.007
R469 VDD2 VDD2.n0 0.175069
C0 VN VP 2.94675f
C1 VN w_n1186_n1856# 1.33291f
C2 VDD2 VN 0.61739f
C3 VP VDD1 0.700389f
C4 w_n1186_n1856# VDD1 0.941443f
C5 VP VTAIL 0.436841f
C6 VDD2 VDD1 0.419458f
C7 w_n1186_n1856# VTAIL 1.66003f
C8 VDD2 VTAIL 3.5297f
C9 B VP 0.783625f
C10 B w_n1186_n1856# 4.14854f
C11 VDD2 B 0.804374f
C12 VN VDD1 0.152705f
C13 VN VTAIL 0.422478f
C14 VTAIL VDD1 3.49578f
C15 VN B 0.55342f
C16 VP w_n1186_n1856# 1.47849f
C17 VDD2 VP 0.237931f
C18 VDD2 w_n1186_n1856# 0.940961f
C19 B VDD1 0.792954f
C20 B VTAIL 1.14825f
C21 VDD2 VSUBS 0.439404f
C22 VDD1 VSUBS 2.682535f
C23 VTAIL VSUBS 0.135393f
C24 VN VSUBS 3.67455f
C25 VP VSUBS 0.626199f
C26 B VSUBS 1.438791f
C27 w_n1186_n1856# VSUBS 27.6528f
C28 VDD2.t1 VSUBS 0.779499f
C29 VDD2.t0 VSUBS 0.592637f
C30 VDD2.n0 VSUBS 2.10048f
C31 VN.t0 VSUBS 0.139078f
C32 VN.t1 VSUBS 0.187442f
C33 B.n0 VSUBS 0.004722f
C34 B.n1 VSUBS 0.004722f
C35 B.n2 VSUBS 0.007467f
C36 B.n3 VSUBS 0.007467f
C37 B.n4 VSUBS 0.007467f
C38 B.n5 VSUBS 0.007467f
C39 B.n6 VSUBS 0.007467f
C40 B.n7 VSUBS 0.018664f
C41 B.n8 VSUBS 0.007467f
C42 B.n9 VSUBS 0.007467f
C43 B.n10 VSUBS 0.007467f
C44 B.n11 VSUBS 0.007467f
C45 B.n12 VSUBS 0.007467f
C46 B.n13 VSUBS 0.007467f
C47 B.n14 VSUBS 0.007467f
C48 B.n15 VSUBS 0.007467f
C49 B.n16 VSUBS 0.007467f
C50 B.n17 VSUBS 0.007467f
C51 B.t2 VSUBS 0.127012f
C52 B.t1 VSUBS 0.131121f
C53 B.t0 VSUBS 0.040418f
C54 B.n18 VSUBS 0.068979f
C55 B.n19 VSUBS 0.06383f
C56 B.n20 VSUBS 0.007467f
C57 B.n21 VSUBS 0.007467f
C58 B.n22 VSUBS 0.007467f
C59 B.n23 VSUBS 0.007467f
C60 B.t8 VSUBS 0.127012f
C61 B.t7 VSUBS 0.131121f
C62 B.t6 VSUBS 0.040418f
C63 B.n24 VSUBS 0.068979f
C64 B.n25 VSUBS 0.06383f
C65 B.n26 VSUBS 0.017301f
C66 B.n27 VSUBS 0.007467f
C67 B.n28 VSUBS 0.007467f
C68 B.n29 VSUBS 0.007467f
C69 B.n30 VSUBS 0.007467f
C70 B.n31 VSUBS 0.007467f
C71 B.n32 VSUBS 0.007467f
C72 B.n33 VSUBS 0.007467f
C73 B.n34 VSUBS 0.007467f
C74 B.n35 VSUBS 0.007467f
C75 B.n36 VSUBS 0.019437f
C76 B.n37 VSUBS 0.007467f
C77 B.n38 VSUBS 0.007467f
C78 B.n39 VSUBS 0.007467f
C79 B.n40 VSUBS 0.007467f
C80 B.n41 VSUBS 0.007467f
C81 B.n42 VSUBS 0.007467f
C82 B.n43 VSUBS 0.007467f
C83 B.n44 VSUBS 0.007467f
C84 B.n45 VSUBS 0.007467f
C85 B.n46 VSUBS 0.007467f
C86 B.n47 VSUBS 0.018664f
C87 B.n48 VSUBS 0.007467f
C88 B.n49 VSUBS 0.007467f
C89 B.n50 VSUBS 0.007467f
C90 B.n51 VSUBS 0.007467f
C91 B.n52 VSUBS 0.007467f
C92 B.n53 VSUBS 0.007467f
C93 B.n54 VSUBS 0.007467f
C94 B.n55 VSUBS 0.007467f
C95 B.n56 VSUBS 0.007467f
C96 B.n57 VSUBS 0.007467f
C97 B.t10 VSUBS 0.127012f
C98 B.t11 VSUBS 0.131121f
C99 B.t9 VSUBS 0.040418f
C100 B.n58 VSUBS 0.068979f
C101 B.n59 VSUBS 0.06383f
C102 B.n60 VSUBS 0.007467f
C103 B.n61 VSUBS 0.007467f
C104 B.n62 VSUBS 0.007467f
C105 B.n63 VSUBS 0.007467f
C106 B.t4 VSUBS 0.127012f
C107 B.t5 VSUBS 0.131121f
C108 B.t3 VSUBS 0.040418f
C109 B.n64 VSUBS 0.068979f
C110 B.n65 VSUBS 0.06383f
C111 B.n66 VSUBS 0.017301f
C112 B.n67 VSUBS 0.007467f
C113 B.n68 VSUBS 0.007467f
C114 B.n69 VSUBS 0.007467f
C115 B.n70 VSUBS 0.007467f
C116 B.n71 VSUBS 0.007467f
C117 B.n72 VSUBS 0.007467f
C118 B.n73 VSUBS 0.007467f
C119 B.n74 VSUBS 0.007467f
C120 B.n75 VSUBS 0.007467f
C121 B.n76 VSUBS 0.018664f
C122 B.n77 VSUBS 0.007467f
C123 B.n78 VSUBS 0.007467f
C124 B.n79 VSUBS 0.007467f
C125 B.n80 VSUBS 0.007467f
C126 B.n81 VSUBS 0.007467f
C127 B.n82 VSUBS 0.007467f
C128 B.n83 VSUBS 0.007467f
C129 B.n84 VSUBS 0.007467f
C130 B.n85 VSUBS 0.007467f
C131 B.n86 VSUBS 0.007467f
C132 B.n87 VSUBS 0.007467f
C133 B.n88 VSUBS 0.007467f
C134 B.n89 VSUBS 0.007467f
C135 B.n90 VSUBS 0.007467f
C136 B.n91 VSUBS 0.007467f
C137 B.n92 VSUBS 0.007467f
C138 B.n93 VSUBS 0.007467f
C139 B.n94 VSUBS 0.007467f
C140 B.n95 VSUBS 0.018664f
C141 B.n96 VSUBS 0.01955f
C142 B.n97 VSUBS 0.01955f
C143 B.n98 VSUBS 0.007467f
C144 B.n99 VSUBS 0.007467f
C145 B.n100 VSUBS 0.007467f
C146 B.n101 VSUBS 0.007467f
C147 B.n102 VSUBS 0.007467f
C148 B.n103 VSUBS 0.007467f
C149 B.n104 VSUBS 0.007467f
C150 B.n105 VSUBS 0.007467f
C151 B.n106 VSUBS 0.007467f
C152 B.n107 VSUBS 0.007467f
C153 B.n108 VSUBS 0.007467f
C154 B.n109 VSUBS 0.007467f
C155 B.n110 VSUBS 0.007467f
C156 B.n111 VSUBS 0.007467f
C157 B.n112 VSUBS 0.007467f
C158 B.n113 VSUBS 0.007467f
C159 B.n114 VSUBS 0.007467f
C160 B.n115 VSUBS 0.007467f
C161 B.n116 VSUBS 0.007467f
C162 B.n117 VSUBS 0.007467f
C163 B.n118 VSUBS 0.007467f
C164 B.n119 VSUBS 0.007467f
C165 B.n120 VSUBS 0.007467f
C166 B.n121 VSUBS 0.007467f
C167 B.n122 VSUBS 0.007467f
C168 B.n123 VSUBS 0.006808f
C169 B.n124 VSUBS 0.007467f
C170 B.n125 VSUBS 0.007467f
C171 B.n126 VSUBS 0.004392f
C172 B.n127 VSUBS 0.007467f
C173 B.n128 VSUBS 0.007467f
C174 B.n129 VSUBS 0.007467f
C175 B.n130 VSUBS 0.007467f
C176 B.n131 VSUBS 0.007467f
C177 B.n132 VSUBS 0.007467f
C178 B.n133 VSUBS 0.007467f
C179 B.n134 VSUBS 0.007467f
C180 B.n135 VSUBS 0.007467f
C181 B.n136 VSUBS 0.007467f
C182 B.n137 VSUBS 0.007467f
C183 B.n138 VSUBS 0.007467f
C184 B.n139 VSUBS 0.004392f
C185 B.n140 VSUBS 0.017301f
C186 B.n141 VSUBS 0.006808f
C187 B.n142 VSUBS 0.007467f
C188 B.n143 VSUBS 0.007467f
C189 B.n144 VSUBS 0.007467f
C190 B.n145 VSUBS 0.007467f
C191 B.n146 VSUBS 0.007467f
C192 B.n147 VSUBS 0.007467f
C193 B.n148 VSUBS 0.007467f
C194 B.n149 VSUBS 0.007467f
C195 B.n150 VSUBS 0.007467f
C196 B.n151 VSUBS 0.007467f
C197 B.n152 VSUBS 0.007467f
C198 B.n153 VSUBS 0.007467f
C199 B.n154 VSUBS 0.007467f
C200 B.n155 VSUBS 0.007467f
C201 B.n156 VSUBS 0.007467f
C202 B.n157 VSUBS 0.007467f
C203 B.n158 VSUBS 0.007467f
C204 B.n159 VSUBS 0.007467f
C205 B.n160 VSUBS 0.007467f
C206 B.n161 VSUBS 0.007467f
C207 B.n162 VSUBS 0.007467f
C208 B.n163 VSUBS 0.007467f
C209 B.n164 VSUBS 0.007467f
C210 B.n165 VSUBS 0.007467f
C211 B.n166 VSUBS 0.007467f
C212 B.n167 VSUBS 0.007467f
C213 B.n168 VSUBS 0.01955f
C214 B.n169 VSUBS 0.01955f
C215 B.n170 VSUBS 0.018664f
C216 B.n171 VSUBS 0.007467f
C217 B.n172 VSUBS 0.007467f
C218 B.n173 VSUBS 0.007467f
C219 B.n174 VSUBS 0.007467f
C220 B.n175 VSUBS 0.007467f
C221 B.n176 VSUBS 0.007467f
C222 B.n177 VSUBS 0.007467f
C223 B.n178 VSUBS 0.007467f
C224 B.n179 VSUBS 0.007467f
C225 B.n180 VSUBS 0.007467f
C226 B.n181 VSUBS 0.007467f
C227 B.n182 VSUBS 0.007467f
C228 B.n183 VSUBS 0.007467f
C229 B.n184 VSUBS 0.007467f
C230 B.n185 VSUBS 0.007467f
C231 B.n186 VSUBS 0.007467f
C232 B.n187 VSUBS 0.007467f
C233 B.n188 VSUBS 0.007467f
C234 B.n189 VSUBS 0.007467f
C235 B.n190 VSUBS 0.007467f
C236 B.n191 VSUBS 0.007467f
C237 B.n192 VSUBS 0.007467f
C238 B.n193 VSUBS 0.007467f
C239 B.n194 VSUBS 0.007467f
C240 B.n195 VSUBS 0.007467f
C241 B.n196 VSUBS 0.007467f
C242 B.n197 VSUBS 0.007467f
C243 B.n198 VSUBS 0.007467f
C244 B.n199 VSUBS 0.007467f
C245 B.n200 VSUBS 0.007467f
C246 B.n201 VSUBS 0.007467f
C247 B.n202 VSUBS 0.007467f
C248 B.n203 VSUBS 0.018664f
C249 B.n204 VSUBS 0.01955f
C250 B.n205 VSUBS 0.018777f
C251 B.n206 VSUBS 0.007467f
C252 B.n207 VSUBS 0.007467f
C253 B.n208 VSUBS 0.007467f
C254 B.n209 VSUBS 0.007467f
C255 B.n210 VSUBS 0.007467f
C256 B.n211 VSUBS 0.007467f
C257 B.n212 VSUBS 0.007467f
C258 B.n213 VSUBS 0.007467f
C259 B.n214 VSUBS 0.007467f
C260 B.n215 VSUBS 0.007467f
C261 B.n216 VSUBS 0.007467f
C262 B.n217 VSUBS 0.007467f
C263 B.n218 VSUBS 0.007467f
C264 B.n219 VSUBS 0.007467f
C265 B.n220 VSUBS 0.007467f
C266 B.n221 VSUBS 0.007467f
C267 B.n222 VSUBS 0.007467f
C268 B.n223 VSUBS 0.007467f
C269 B.n224 VSUBS 0.007467f
C270 B.n225 VSUBS 0.007467f
C271 B.n226 VSUBS 0.007467f
C272 B.n227 VSUBS 0.007467f
C273 B.n228 VSUBS 0.007467f
C274 B.n229 VSUBS 0.007467f
C275 B.n230 VSUBS 0.007467f
C276 B.n231 VSUBS 0.006808f
C277 B.n232 VSUBS 0.007467f
C278 B.n233 VSUBS 0.007467f
C279 B.n234 VSUBS 0.004392f
C280 B.n235 VSUBS 0.007467f
C281 B.n236 VSUBS 0.007467f
C282 B.n237 VSUBS 0.007467f
C283 B.n238 VSUBS 0.007467f
C284 B.n239 VSUBS 0.007467f
C285 B.n240 VSUBS 0.007467f
C286 B.n241 VSUBS 0.007467f
C287 B.n242 VSUBS 0.007467f
C288 B.n243 VSUBS 0.007467f
C289 B.n244 VSUBS 0.007467f
C290 B.n245 VSUBS 0.007467f
C291 B.n246 VSUBS 0.007467f
C292 B.n247 VSUBS 0.004392f
C293 B.n248 VSUBS 0.017301f
C294 B.n249 VSUBS 0.006808f
C295 B.n250 VSUBS 0.007467f
C296 B.n251 VSUBS 0.007467f
C297 B.n252 VSUBS 0.007467f
C298 B.n253 VSUBS 0.007467f
C299 B.n254 VSUBS 0.007467f
C300 B.n255 VSUBS 0.007467f
C301 B.n256 VSUBS 0.007467f
C302 B.n257 VSUBS 0.007467f
C303 B.n258 VSUBS 0.007467f
C304 B.n259 VSUBS 0.007467f
C305 B.n260 VSUBS 0.007467f
C306 B.n261 VSUBS 0.007467f
C307 B.n262 VSUBS 0.007467f
C308 B.n263 VSUBS 0.007467f
C309 B.n264 VSUBS 0.007467f
C310 B.n265 VSUBS 0.007467f
C311 B.n266 VSUBS 0.007467f
C312 B.n267 VSUBS 0.007467f
C313 B.n268 VSUBS 0.007467f
C314 B.n269 VSUBS 0.007467f
C315 B.n270 VSUBS 0.007467f
C316 B.n271 VSUBS 0.007467f
C317 B.n272 VSUBS 0.007467f
C318 B.n273 VSUBS 0.007467f
C319 B.n274 VSUBS 0.007467f
C320 B.n275 VSUBS 0.007467f
C321 B.n276 VSUBS 0.01955f
C322 B.n277 VSUBS 0.01955f
C323 B.n278 VSUBS 0.018664f
C324 B.n279 VSUBS 0.007467f
C325 B.n280 VSUBS 0.007467f
C326 B.n281 VSUBS 0.007467f
C327 B.n282 VSUBS 0.007467f
C328 B.n283 VSUBS 0.007467f
C329 B.n284 VSUBS 0.007467f
C330 B.n285 VSUBS 0.007467f
C331 B.n286 VSUBS 0.007467f
C332 B.n287 VSUBS 0.007467f
C333 B.n288 VSUBS 0.007467f
C334 B.n289 VSUBS 0.007467f
C335 B.n290 VSUBS 0.007467f
C336 B.n291 VSUBS 0.007467f
C337 B.n292 VSUBS 0.007467f
C338 B.n293 VSUBS 0.007467f
C339 B.n294 VSUBS 0.007467f
C340 B.n295 VSUBS 0.016908f
C341 VDD1.t1 VSUBS 0.58063f
C342 VDD1.t0 VSUBS 0.77522f
C343 VTAIL.t2 VSUBS 0.621256f
C344 VTAIL.n0 VSUBS 1.14198f
C345 VTAIL.t0 VSUBS 0.621258f
C346 VTAIL.n1 VSUBS 1.14639f
C347 VTAIL.t3 VSUBS 0.621256f
C348 VTAIL.n2 VSUBS 1.1111f
C349 VTAIL.t1 VSUBS 0.621256f
C350 VTAIL.n3 VSUBS 1.06224f
C351 VP.t0 VSUBS 0.190027f
C352 VP.t1 VSUBS 0.142278f
C353 VP.n0 VSUBS 2.56198f
.ends

