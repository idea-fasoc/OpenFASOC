* NGSPICE file created from diff_pair_sample_1109.ext - technology: sky130A

.subckt diff_pair_sample_1109 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=1.8525 ps=10.28 w=4.75 l=1.34
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=0 ps=0 w=4.75 l=1.34
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=1.8525 ps=10.28 w=4.75 l=1.34
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=0 ps=0 w=4.75 l=1.34
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=0 ps=0 w=4.75 l=1.34
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=1.8525 ps=10.28 w=4.75 l=1.34
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=1.8525 ps=10.28 w=4.75 l=1.34
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8525 pd=10.28 as=0 ps=0 w=4.75 l=1.34
R0 VP.n0 VP.t0 231.351
R1 VP.n0 VP.t1 195.529
R2 VP VP.n0 0.146778
R3 VTAIL.n90 VTAIL.n72 289.615
R4 VTAIL.n18 VTAIL.n0 289.615
R5 VTAIL.n66 VTAIL.n48 289.615
R6 VTAIL.n42 VTAIL.n24 289.615
R7 VTAIL.n81 VTAIL.n80 185
R8 VTAIL.n83 VTAIL.n82 185
R9 VTAIL.n76 VTAIL.n75 185
R10 VTAIL.n89 VTAIL.n88 185
R11 VTAIL.n91 VTAIL.n90 185
R12 VTAIL.n9 VTAIL.n8 185
R13 VTAIL.n11 VTAIL.n10 185
R14 VTAIL.n4 VTAIL.n3 185
R15 VTAIL.n17 VTAIL.n16 185
R16 VTAIL.n19 VTAIL.n18 185
R17 VTAIL.n67 VTAIL.n66 185
R18 VTAIL.n65 VTAIL.n64 185
R19 VTAIL.n52 VTAIL.n51 185
R20 VTAIL.n59 VTAIL.n58 185
R21 VTAIL.n57 VTAIL.n56 185
R22 VTAIL.n43 VTAIL.n42 185
R23 VTAIL.n41 VTAIL.n40 185
R24 VTAIL.n28 VTAIL.n27 185
R25 VTAIL.n35 VTAIL.n34 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n79 VTAIL.t0 147.714
R28 VTAIL.n7 VTAIL.t3 147.714
R29 VTAIL.n55 VTAIL.t2 147.714
R30 VTAIL.n31 VTAIL.t1 147.714
R31 VTAIL.n82 VTAIL.n81 104.615
R32 VTAIL.n82 VTAIL.n75 104.615
R33 VTAIL.n89 VTAIL.n75 104.615
R34 VTAIL.n90 VTAIL.n89 104.615
R35 VTAIL.n10 VTAIL.n9 104.615
R36 VTAIL.n10 VTAIL.n3 104.615
R37 VTAIL.n17 VTAIL.n3 104.615
R38 VTAIL.n18 VTAIL.n17 104.615
R39 VTAIL.n66 VTAIL.n65 104.615
R40 VTAIL.n65 VTAIL.n51 104.615
R41 VTAIL.n58 VTAIL.n51 104.615
R42 VTAIL.n58 VTAIL.n57 104.615
R43 VTAIL.n42 VTAIL.n41 104.615
R44 VTAIL.n41 VTAIL.n27 104.615
R45 VTAIL.n34 VTAIL.n27 104.615
R46 VTAIL.n34 VTAIL.n33 104.615
R47 VTAIL.n81 VTAIL.t0 52.3082
R48 VTAIL.n9 VTAIL.t3 52.3082
R49 VTAIL.n57 VTAIL.t2 52.3082
R50 VTAIL.n33 VTAIL.t1 52.3082
R51 VTAIL.n95 VTAIL.n94 35.8702
R52 VTAIL.n23 VTAIL.n22 35.8702
R53 VTAIL.n71 VTAIL.n70 35.8702
R54 VTAIL.n47 VTAIL.n46 35.8702
R55 VTAIL.n47 VTAIL.n23 19.341
R56 VTAIL.n95 VTAIL.n71 17.9014
R57 VTAIL.n80 VTAIL.n79 15.6631
R58 VTAIL.n8 VTAIL.n7 15.6631
R59 VTAIL.n56 VTAIL.n55 15.6631
R60 VTAIL.n32 VTAIL.n31 15.6631
R61 VTAIL.n83 VTAIL.n78 12.8005
R62 VTAIL.n11 VTAIL.n6 12.8005
R63 VTAIL.n59 VTAIL.n54 12.8005
R64 VTAIL.n35 VTAIL.n30 12.8005
R65 VTAIL.n84 VTAIL.n76 12.0247
R66 VTAIL.n12 VTAIL.n4 12.0247
R67 VTAIL.n60 VTAIL.n52 12.0247
R68 VTAIL.n36 VTAIL.n28 12.0247
R69 VTAIL.n88 VTAIL.n87 11.249
R70 VTAIL.n16 VTAIL.n15 11.249
R71 VTAIL.n64 VTAIL.n63 11.249
R72 VTAIL.n40 VTAIL.n39 11.249
R73 VTAIL.n91 VTAIL.n74 10.4732
R74 VTAIL.n19 VTAIL.n2 10.4732
R75 VTAIL.n67 VTAIL.n50 10.4732
R76 VTAIL.n43 VTAIL.n26 10.4732
R77 VTAIL.n92 VTAIL.n72 9.69747
R78 VTAIL.n20 VTAIL.n0 9.69747
R79 VTAIL.n68 VTAIL.n48 9.69747
R80 VTAIL.n44 VTAIL.n24 9.69747
R81 VTAIL.n94 VTAIL.n93 9.45567
R82 VTAIL.n22 VTAIL.n21 9.45567
R83 VTAIL.n70 VTAIL.n69 9.45567
R84 VTAIL.n46 VTAIL.n45 9.45567
R85 VTAIL.n93 VTAIL.n92 9.3005
R86 VTAIL.n74 VTAIL.n73 9.3005
R87 VTAIL.n87 VTAIL.n86 9.3005
R88 VTAIL.n85 VTAIL.n84 9.3005
R89 VTAIL.n78 VTAIL.n77 9.3005
R90 VTAIL.n21 VTAIL.n20 9.3005
R91 VTAIL.n2 VTAIL.n1 9.3005
R92 VTAIL.n15 VTAIL.n14 9.3005
R93 VTAIL.n13 VTAIL.n12 9.3005
R94 VTAIL.n6 VTAIL.n5 9.3005
R95 VTAIL.n69 VTAIL.n68 9.3005
R96 VTAIL.n50 VTAIL.n49 9.3005
R97 VTAIL.n63 VTAIL.n62 9.3005
R98 VTAIL.n61 VTAIL.n60 9.3005
R99 VTAIL.n54 VTAIL.n53 9.3005
R100 VTAIL.n45 VTAIL.n44 9.3005
R101 VTAIL.n26 VTAIL.n25 9.3005
R102 VTAIL.n39 VTAIL.n38 9.3005
R103 VTAIL.n37 VTAIL.n36 9.3005
R104 VTAIL.n30 VTAIL.n29 9.3005
R105 VTAIL.n79 VTAIL.n77 4.39059
R106 VTAIL.n7 VTAIL.n5 4.39059
R107 VTAIL.n55 VTAIL.n53 4.39059
R108 VTAIL.n31 VTAIL.n29 4.39059
R109 VTAIL.n94 VTAIL.n72 4.26717
R110 VTAIL.n22 VTAIL.n0 4.26717
R111 VTAIL.n70 VTAIL.n48 4.26717
R112 VTAIL.n46 VTAIL.n24 4.26717
R113 VTAIL.n92 VTAIL.n91 3.49141
R114 VTAIL.n20 VTAIL.n19 3.49141
R115 VTAIL.n68 VTAIL.n67 3.49141
R116 VTAIL.n44 VTAIL.n43 3.49141
R117 VTAIL.n88 VTAIL.n74 2.71565
R118 VTAIL.n16 VTAIL.n2 2.71565
R119 VTAIL.n64 VTAIL.n50 2.71565
R120 VTAIL.n40 VTAIL.n26 2.71565
R121 VTAIL.n87 VTAIL.n76 1.93989
R122 VTAIL.n15 VTAIL.n4 1.93989
R123 VTAIL.n63 VTAIL.n52 1.93989
R124 VTAIL.n39 VTAIL.n28 1.93989
R125 VTAIL.n71 VTAIL.n47 1.19016
R126 VTAIL.n84 VTAIL.n83 1.16414
R127 VTAIL.n12 VTAIL.n11 1.16414
R128 VTAIL.n60 VTAIL.n59 1.16414
R129 VTAIL.n36 VTAIL.n35 1.16414
R130 VTAIL VTAIL.n23 0.888431
R131 VTAIL.n80 VTAIL.n78 0.388379
R132 VTAIL.n8 VTAIL.n6 0.388379
R133 VTAIL.n56 VTAIL.n54 0.388379
R134 VTAIL.n32 VTAIL.n30 0.388379
R135 VTAIL VTAIL.n95 0.302224
R136 VTAIL.n85 VTAIL.n77 0.155672
R137 VTAIL.n86 VTAIL.n85 0.155672
R138 VTAIL.n86 VTAIL.n73 0.155672
R139 VTAIL.n93 VTAIL.n73 0.155672
R140 VTAIL.n13 VTAIL.n5 0.155672
R141 VTAIL.n14 VTAIL.n13 0.155672
R142 VTAIL.n14 VTAIL.n1 0.155672
R143 VTAIL.n21 VTAIL.n1 0.155672
R144 VTAIL.n69 VTAIL.n49 0.155672
R145 VTAIL.n62 VTAIL.n49 0.155672
R146 VTAIL.n62 VTAIL.n61 0.155672
R147 VTAIL.n61 VTAIL.n53 0.155672
R148 VTAIL.n45 VTAIL.n25 0.155672
R149 VTAIL.n38 VTAIL.n25 0.155672
R150 VTAIL.n38 VTAIL.n37 0.155672
R151 VTAIL.n37 VTAIL.n29 0.155672
R152 VDD1.n18 VDD1.n0 289.615
R153 VDD1.n41 VDD1.n23 289.615
R154 VDD1.n19 VDD1.n18 185
R155 VDD1.n17 VDD1.n16 185
R156 VDD1.n4 VDD1.n3 185
R157 VDD1.n11 VDD1.n10 185
R158 VDD1.n9 VDD1.n8 185
R159 VDD1.n32 VDD1.n31 185
R160 VDD1.n34 VDD1.n33 185
R161 VDD1.n27 VDD1.n26 185
R162 VDD1.n40 VDD1.n39 185
R163 VDD1.n42 VDD1.n41 185
R164 VDD1.n7 VDD1.t1 147.714
R165 VDD1.n30 VDD1.t0 147.714
R166 VDD1.n18 VDD1.n17 104.615
R167 VDD1.n17 VDD1.n3 104.615
R168 VDD1.n10 VDD1.n3 104.615
R169 VDD1.n10 VDD1.n9 104.615
R170 VDD1.n33 VDD1.n32 104.615
R171 VDD1.n33 VDD1.n26 104.615
R172 VDD1.n40 VDD1.n26 104.615
R173 VDD1.n41 VDD1.n40 104.615
R174 VDD1 VDD1.n45 84.0673
R175 VDD1 VDD1.n22 52.9671
R176 VDD1.n9 VDD1.t1 52.3082
R177 VDD1.n32 VDD1.t0 52.3082
R178 VDD1.n8 VDD1.n7 15.6631
R179 VDD1.n31 VDD1.n30 15.6631
R180 VDD1.n11 VDD1.n6 12.8005
R181 VDD1.n34 VDD1.n29 12.8005
R182 VDD1.n12 VDD1.n4 12.0247
R183 VDD1.n35 VDD1.n27 12.0247
R184 VDD1.n16 VDD1.n15 11.249
R185 VDD1.n39 VDD1.n38 11.249
R186 VDD1.n19 VDD1.n2 10.4732
R187 VDD1.n42 VDD1.n25 10.4732
R188 VDD1.n20 VDD1.n0 9.69747
R189 VDD1.n43 VDD1.n23 9.69747
R190 VDD1.n22 VDD1.n21 9.45567
R191 VDD1.n45 VDD1.n44 9.45567
R192 VDD1.n21 VDD1.n20 9.3005
R193 VDD1.n2 VDD1.n1 9.3005
R194 VDD1.n15 VDD1.n14 9.3005
R195 VDD1.n13 VDD1.n12 9.3005
R196 VDD1.n6 VDD1.n5 9.3005
R197 VDD1.n44 VDD1.n43 9.3005
R198 VDD1.n25 VDD1.n24 9.3005
R199 VDD1.n38 VDD1.n37 9.3005
R200 VDD1.n36 VDD1.n35 9.3005
R201 VDD1.n29 VDD1.n28 9.3005
R202 VDD1.n7 VDD1.n5 4.39059
R203 VDD1.n30 VDD1.n28 4.39059
R204 VDD1.n22 VDD1.n0 4.26717
R205 VDD1.n45 VDD1.n23 4.26717
R206 VDD1.n20 VDD1.n19 3.49141
R207 VDD1.n43 VDD1.n42 3.49141
R208 VDD1.n16 VDD1.n2 2.71565
R209 VDD1.n39 VDD1.n25 2.71565
R210 VDD1.n15 VDD1.n4 1.93989
R211 VDD1.n38 VDD1.n27 1.93989
R212 VDD1.n12 VDD1.n11 1.16414
R213 VDD1.n35 VDD1.n34 1.16414
R214 VDD1.n8 VDD1.n6 0.388379
R215 VDD1.n31 VDD1.n29 0.388379
R216 VDD1.n21 VDD1.n1 0.155672
R217 VDD1.n14 VDD1.n1 0.155672
R218 VDD1.n14 VDD1.n13 0.155672
R219 VDD1.n13 VDD1.n5 0.155672
R220 VDD1.n36 VDD1.n28 0.155672
R221 VDD1.n37 VDD1.n36 0.155672
R222 VDD1.n37 VDD1.n24 0.155672
R223 VDD1.n44 VDD1.n24 0.155672
R224 B.n309 B.n308 585
R225 B.n311 B.n66 585
R226 B.n314 B.n313 585
R227 B.n315 B.n65 585
R228 B.n317 B.n316 585
R229 B.n319 B.n64 585
R230 B.n322 B.n321 585
R231 B.n323 B.n63 585
R232 B.n325 B.n324 585
R233 B.n327 B.n62 585
R234 B.n330 B.n329 585
R235 B.n331 B.n61 585
R236 B.n333 B.n332 585
R237 B.n335 B.n60 585
R238 B.n338 B.n337 585
R239 B.n339 B.n59 585
R240 B.n341 B.n340 585
R241 B.n343 B.n58 585
R242 B.n345 B.n344 585
R243 B.n347 B.n346 585
R244 B.n350 B.n349 585
R245 B.n351 B.n53 585
R246 B.n353 B.n352 585
R247 B.n355 B.n52 585
R248 B.n358 B.n357 585
R249 B.n359 B.n51 585
R250 B.n361 B.n360 585
R251 B.n363 B.n50 585
R252 B.n366 B.n365 585
R253 B.n367 B.n47 585
R254 B.n370 B.n369 585
R255 B.n372 B.n46 585
R256 B.n375 B.n374 585
R257 B.n376 B.n45 585
R258 B.n378 B.n377 585
R259 B.n380 B.n44 585
R260 B.n383 B.n382 585
R261 B.n384 B.n43 585
R262 B.n386 B.n385 585
R263 B.n388 B.n42 585
R264 B.n391 B.n390 585
R265 B.n392 B.n41 585
R266 B.n394 B.n393 585
R267 B.n396 B.n40 585
R268 B.n399 B.n398 585
R269 B.n400 B.n39 585
R270 B.n402 B.n401 585
R271 B.n404 B.n38 585
R272 B.n407 B.n406 585
R273 B.n408 B.n37 585
R274 B.n307 B.n35 585
R275 B.n411 B.n35 585
R276 B.n306 B.n34 585
R277 B.n412 B.n34 585
R278 B.n305 B.n33 585
R279 B.n413 B.n33 585
R280 B.n304 B.n303 585
R281 B.n303 B.n29 585
R282 B.n302 B.n28 585
R283 B.n419 B.n28 585
R284 B.n301 B.n27 585
R285 B.n420 B.n27 585
R286 B.n300 B.n26 585
R287 B.n421 B.n26 585
R288 B.n299 B.n298 585
R289 B.n298 B.n22 585
R290 B.n297 B.n21 585
R291 B.n427 B.n21 585
R292 B.n296 B.n20 585
R293 B.n428 B.n20 585
R294 B.n295 B.n19 585
R295 B.n429 B.n19 585
R296 B.n294 B.n293 585
R297 B.n293 B.n15 585
R298 B.n292 B.n14 585
R299 B.n435 B.n14 585
R300 B.n291 B.n13 585
R301 B.n436 B.n13 585
R302 B.n290 B.n12 585
R303 B.n437 B.n12 585
R304 B.n289 B.n288 585
R305 B.n288 B.n8 585
R306 B.n287 B.n7 585
R307 B.n443 B.n7 585
R308 B.n286 B.n6 585
R309 B.n444 B.n6 585
R310 B.n285 B.n5 585
R311 B.n445 B.n5 585
R312 B.n284 B.n283 585
R313 B.n283 B.n4 585
R314 B.n282 B.n67 585
R315 B.n282 B.n281 585
R316 B.n272 B.n68 585
R317 B.n69 B.n68 585
R318 B.n274 B.n273 585
R319 B.n275 B.n274 585
R320 B.n271 B.n73 585
R321 B.n77 B.n73 585
R322 B.n270 B.n269 585
R323 B.n269 B.n268 585
R324 B.n75 B.n74 585
R325 B.n76 B.n75 585
R326 B.n261 B.n260 585
R327 B.n262 B.n261 585
R328 B.n259 B.n82 585
R329 B.n82 B.n81 585
R330 B.n258 B.n257 585
R331 B.n257 B.n256 585
R332 B.n84 B.n83 585
R333 B.n85 B.n84 585
R334 B.n249 B.n248 585
R335 B.n250 B.n249 585
R336 B.n247 B.n89 585
R337 B.n93 B.n89 585
R338 B.n246 B.n245 585
R339 B.n245 B.n244 585
R340 B.n91 B.n90 585
R341 B.n92 B.n91 585
R342 B.n237 B.n236 585
R343 B.n238 B.n237 585
R344 B.n235 B.n98 585
R345 B.n98 B.n97 585
R346 B.n234 B.n233 585
R347 B.n233 B.n232 585
R348 B.n229 B.n102 585
R349 B.n228 B.n227 585
R350 B.n225 B.n103 585
R351 B.n225 B.n101 585
R352 B.n224 B.n223 585
R353 B.n222 B.n221 585
R354 B.n220 B.n105 585
R355 B.n218 B.n217 585
R356 B.n216 B.n106 585
R357 B.n215 B.n214 585
R358 B.n212 B.n107 585
R359 B.n210 B.n209 585
R360 B.n208 B.n108 585
R361 B.n207 B.n206 585
R362 B.n204 B.n109 585
R363 B.n202 B.n201 585
R364 B.n200 B.n110 585
R365 B.n199 B.n198 585
R366 B.n196 B.n111 585
R367 B.n194 B.n193 585
R368 B.n192 B.n112 585
R369 B.n190 B.n189 585
R370 B.n187 B.n115 585
R371 B.n185 B.n184 585
R372 B.n183 B.n116 585
R373 B.n182 B.n181 585
R374 B.n179 B.n117 585
R375 B.n177 B.n176 585
R376 B.n175 B.n118 585
R377 B.n174 B.n173 585
R378 B.n171 B.n119 585
R379 B.n169 B.n168 585
R380 B.n167 B.n120 585
R381 B.n166 B.n165 585
R382 B.n163 B.n124 585
R383 B.n161 B.n160 585
R384 B.n159 B.n125 585
R385 B.n158 B.n157 585
R386 B.n155 B.n126 585
R387 B.n153 B.n152 585
R388 B.n151 B.n127 585
R389 B.n150 B.n149 585
R390 B.n147 B.n128 585
R391 B.n145 B.n144 585
R392 B.n143 B.n129 585
R393 B.n142 B.n141 585
R394 B.n139 B.n130 585
R395 B.n137 B.n136 585
R396 B.n135 B.n131 585
R397 B.n134 B.n133 585
R398 B.n100 B.n99 585
R399 B.n101 B.n100 585
R400 B.n231 B.n230 585
R401 B.n232 B.n231 585
R402 B.n96 B.n95 585
R403 B.n97 B.n96 585
R404 B.n240 B.n239 585
R405 B.n239 B.n238 585
R406 B.n241 B.n94 585
R407 B.n94 B.n92 585
R408 B.n243 B.n242 585
R409 B.n244 B.n243 585
R410 B.n88 B.n87 585
R411 B.n93 B.n88 585
R412 B.n252 B.n251 585
R413 B.n251 B.n250 585
R414 B.n253 B.n86 585
R415 B.n86 B.n85 585
R416 B.n255 B.n254 585
R417 B.n256 B.n255 585
R418 B.n80 B.n79 585
R419 B.n81 B.n80 585
R420 B.n264 B.n263 585
R421 B.n263 B.n262 585
R422 B.n265 B.n78 585
R423 B.n78 B.n76 585
R424 B.n267 B.n266 585
R425 B.n268 B.n267 585
R426 B.n72 B.n71 585
R427 B.n77 B.n72 585
R428 B.n277 B.n276 585
R429 B.n276 B.n275 585
R430 B.n278 B.n70 585
R431 B.n70 B.n69 585
R432 B.n280 B.n279 585
R433 B.n281 B.n280 585
R434 B.n2 B.n0 585
R435 B.n4 B.n2 585
R436 B.n3 B.n1 585
R437 B.n444 B.n3 585
R438 B.n442 B.n441 585
R439 B.n443 B.n442 585
R440 B.n440 B.n9 585
R441 B.n9 B.n8 585
R442 B.n439 B.n438 585
R443 B.n438 B.n437 585
R444 B.n11 B.n10 585
R445 B.n436 B.n11 585
R446 B.n434 B.n433 585
R447 B.n435 B.n434 585
R448 B.n432 B.n16 585
R449 B.n16 B.n15 585
R450 B.n431 B.n430 585
R451 B.n430 B.n429 585
R452 B.n18 B.n17 585
R453 B.n428 B.n18 585
R454 B.n426 B.n425 585
R455 B.n427 B.n426 585
R456 B.n424 B.n23 585
R457 B.n23 B.n22 585
R458 B.n423 B.n422 585
R459 B.n422 B.n421 585
R460 B.n25 B.n24 585
R461 B.n420 B.n25 585
R462 B.n418 B.n417 585
R463 B.n419 B.n418 585
R464 B.n416 B.n30 585
R465 B.n30 B.n29 585
R466 B.n415 B.n414 585
R467 B.n414 B.n413 585
R468 B.n32 B.n31 585
R469 B.n412 B.n32 585
R470 B.n410 B.n409 585
R471 B.n411 B.n410 585
R472 B.n447 B.n446 585
R473 B.n446 B.n445 585
R474 B.n231 B.n102 502.111
R475 B.n410 B.n37 502.111
R476 B.n233 B.n100 502.111
R477 B.n309 B.n35 502.111
R478 B.n121 B.t9 290.219
R479 B.n113 B.t13 290.219
R480 B.n48 B.t6 290.219
R481 B.n54 B.t2 290.219
R482 B.n310 B.n36 256.663
R483 B.n312 B.n36 256.663
R484 B.n318 B.n36 256.663
R485 B.n320 B.n36 256.663
R486 B.n326 B.n36 256.663
R487 B.n328 B.n36 256.663
R488 B.n334 B.n36 256.663
R489 B.n336 B.n36 256.663
R490 B.n342 B.n36 256.663
R491 B.n57 B.n36 256.663
R492 B.n348 B.n36 256.663
R493 B.n354 B.n36 256.663
R494 B.n356 B.n36 256.663
R495 B.n362 B.n36 256.663
R496 B.n364 B.n36 256.663
R497 B.n371 B.n36 256.663
R498 B.n373 B.n36 256.663
R499 B.n379 B.n36 256.663
R500 B.n381 B.n36 256.663
R501 B.n387 B.n36 256.663
R502 B.n389 B.n36 256.663
R503 B.n395 B.n36 256.663
R504 B.n397 B.n36 256.663
R505 B.n403 B.n36 256.663
R506 B.n405 B.n36 256.663
R507 B.n226 B.n101 256.663
R508 B.n104 B.n101 256.663
R509 B.n219 B.n101 256.663
R510 B.n213 B.n101 256.663
R511 B.n211 B.n101 256.663
R512 B.n205 B.n101 256.663
R513 B.n203 B.n101 256.663
R514 B.n197 B.n101 256.663
R515 B.n195 B.n101 256.663
R516 B.n188 B.n101 256.663
R517 B.n186 B.n101 256.663
R518 B.n180 B.n101 256.663
R519 B.n178 B.n101 256.663
R520 B.n172 B.n101 256.663
R521 B.n170 B.n101 256.663
R522 B.n164 B.n101 256.663
R523 B.n162 B.n101 256.663
R524 B.n156 B.n101 256.663
R525 B.n154 B.n101 256.663
R526 B.n148 B.n101 256.663
R527 B.n146 B.n101 256.663
R528 B.n140 B.n101 256.663
R529 B.n138 B.n101 256.663
R530 B.n132 B.n101 256.663
R531 B.n121 B.t12 190.327
R532 B.n54 B.t4 190.327
R533 B.n113 B.t15 190.327
R534 B.n48 B.t7 190.327
R535 B.n231 B.n96 163.367
R536 B.n239 B.n96 163.367
R537 B.n239 B.n94 163.367
R538 B.n243 B.n94 163.367
R539 B.n243 B.n88 163.367
R540 B.n251 B.n88 163.367
R541 B.n251 B.n86 163.367
R542 B.n255 B.n86 163.367
R543 B.n255 B.n80 163.367
R544 B.n263 B.n80 163.367
R545 B.n263 B.n78 163.367
R546 B.n267 B.n78 163.367
R547 B.n267 B.n72 163.367
R548 B.n276 B.n72 163.367
R549 B.n276 B.n70 163.367
R550 B.n280 B.n70 163.367
R551 B.n280 B.n2 163.367
R552 B.n446 B.n2 163.367
R553 B.n446 B.n3 163.367
R554 B.n442 B.n3 163.367
R555 B.n442 B.n9 163.367
R556 B.n438 B.n9 163.367
R557 B.n438 B.n11 163.367
R558 B.n434 B.n11 163.367
R559 B.n434 B.n16 163.367
R560 B.n430 B.n16 163.367
R561 B.n430 B.n18 163.367
R562 B.n426 B.n18 163.367
R563 B.n426 B.n23 163.367
R564 B.n422 B.n23 163.367
R565 B.n422 B.n25 163.367
R566 B.n418 B.n25 163.367
R567 B.n418 B.n30 163.367
R568 B.n414 B.n30 163.367
R569 B.n414 B.n32 163.367
R570 B.n410 B.n32 163.367
R571 B.n227 B.n225 163.367
R572 B.n225 B.n224 163.367
R573 B.n221 B.n220 163.367
R574 B.n218 B.n106 163.367
R575 B.n214 B.n212 163.367
R576 B.n210 B.n108 163.367
R577 B.n206 B.n204 163.367
R578 B.n202 B.n110 163.367
R579 B.n198 B.n196 163.367
R580 B.n194 B.n112 163.367
R581 B.n189 B.n187 163.367
R582 B.n185 B.n116 163.367
R583 B.n181 B.n179 163.367
R584 B.n177 B.n118 163.367
R585 B.n173 B.n171 163.367
R586 B.n169 B.n120 163.367
R587 B.n165 B.n163 163.367
R588 B.n161 B.n125 163.367
R589 B.n157 B.n155 163.367
R590 B.n153 B.n127 163.367
R591 B.n149 B.n147 163.367
R592 B.n145 B.n129 163.367
R593 B.n141 B.n139 163.367
R594 B.n137 B.n131 163.367
R595 B.n133 B.n100 163.367
R596 B.n233 B.n98 163.367
R597 B.n237 B.n98 163.367
R598 B.n237 B.n91 163.367
R599 B.n245 B.n91 163.367
R600 B.n245 B.n89 163.367
R601 B.n249 B.n89 163.367
R602 B.n249 B.n84 163.367
R603 B.n257 B.n84 163.367
R604 B.n257 B.n82 163.367
R605 B.n261 B.n82 163.367
R606 B.n261 B.n75 163.367
R607 B.n269 B.n75 163.367
R608 B.n269 B.n73 163.367
R609 B.n274 B.n73 163.367
R610 B.n274 B.n68 163.367
R611 B.n282 B.n68 163.367
R612 B.n283 B.n282 163.367
R613 B.n283 B.n5 163.367
R614 B.n6 B.n5 163.367
R615 B.n7 B.n6 163.367
R616 B.n288 B.n7 163.367
R617 B.n288 B.n12 163.367
R618 B.n13 B.n12 163.367
R619 B.n14 B.n13 163.367
R620 B.n293 B.n14 163.367
R621 B.n293 B.n19 163.367
R622 B.n20 B.n19 163.367
R623 B.n21 B.n20 163.367
R624 B.n298 B.n21 163.367
R625 B.n298 B.n26 163.367
R626 B.n27 B.n26 163.367
R627 B.n28 B.n27 163.367
R628 B.n303 B.n28 163.367
R629 B.n303 B.n33 163.367
R630 B.n34 B.n33 163.367
R631 B.n35 B.n34 163.367
R632 B.n406 B.n404 163.367
R633 B.n402 B.n39 163.367
R634 B.n398 B.n396 163.367
R635 B.n394 B.n41 163.367
R636 B.n390 B.n388 163.367
R637 B.n386 B.n43 163.367
R638 B.n382 B.n380 163.367
R639 B.n378 B.n45 163.367
R640 B.n374 B.n372 163.367
R641 B.n370 B.n47 163.367
R642 B.n365 B.n363 163.367
R643 B.n361 B.n51 163.367
R644 B.n357 B.n355 163.367
R645 B.n353 B.n53 163.367
R646 B.n349 B.n347 163.367
R647 B.n344 B.n343 163.367
R648 B.n341 B.n59 163.367
R649 B.n337 B.n335 163.367
R650 B.n333 B.n61 163.367
R651 B.n329 B.n327 163.367
R652 B.n325 B.n63 163.367
R653 B.n321 B.n319 163.367
R654 B.n317 B.n65 163.367
R655 B.n313 B.n311 163.367
R656 B.n122 B.t11 157.94
R657 B.n55 B.t5 157.94
R658 B.n114 B.t14 157.94
R659 B.n49 B.t8 157.94
R660 B.n232 B.n101 130.575
R661 B.n411 B.n36 130.575
R662 B.n232 B.n97 74.614
R663 B.n238 B.n97 74.614
R664 B.n238 B.n92 74.614
R665 B.n244 B.n92 74.614
R666 B.n244 B.n93 74.614
R667 B.n250 B.n85 74.614
R668 B.n256 B.n85 74.614
R669 B.n256 B.n81 74.614
R670 B.n262 B.n81 74.614
R671 B.n262 B.n76 74.614
R672 B.n268 B.n76 74.614
R673 B.n268 B.n77 74.614
R674 B.n275 B.n69 74.614
R675 B.n281 B.n69 74.614
R676 B.n281 B.n4 74.614
R677 B.n445 B.n4 74.614
R678 B.n445 B.n444 74.614
R679 B.n444 B.n443 74.614
R680 B.n443 B.n8 74.614
R681 B.n437 B.n8 74.614
R682 B.n436 B.n435 74.614
R683 B.n435 B.n15 74.614
R684 B.n429 B.n15 74.614
R685 B.n429 B.n428 74.614
R686 B.n428 B.n427 74.614
R687 B.n427 B.n22 74.614
R688 B.n421 B.n22 74.614
R689 B.n420 B.n419 74.614
R690 B.n419 B.n29 74.614
R691 B.n413 B.n29 74.614
R692 B.n413 B.n412 74.614
R693 B.n412 B.n411 74.614
R694 B.n226 B.n102 71.676
R695 B.n224 B.n104 71.676
R696 B.n220 B.n219 71.676
R697 B.n213 B.n106 71.676
R698 B.n212 B.n211 71.676
R699 B.n205 B.n108 71.676
R700 B.n204 B.n203 71.676
R701 B.n197 B.n110 71.676
R702 B.n196 B.n195 71.676
R703 B.n188 B.n112 71.676
R704 B.n187 B.n186 71.676
R705 B.n180 B.n116 71.676
R706 B.n179 B.n178 71.676
R707 B.n172 B.n118 71.676
R708 B.n171 B.n170 71.676
R709 B.n164 B.n120 71.676
R710 B.n163 B.n162 71.676
R711 B.n156 B.n125 71.676
R712 B.n155 B.n154 71.676
R713 B.n148 B.n127 71.676
R714 B.n147 B.n146 71.676
R715 B.n140 B.n129 71.676
R716 B.n139 B.n138 71.676
R717 B.n132 B.n131 71.676
R718 B.n405 B.n37 71.676
R719 B.n404 B.n403 71.676
R720 B.n397 B.n39 71.676
R721 B.n396 B.n395 71.676
R722 B.n389 B.n41 71.676
R723 B.n388 B.n387 71.676
R724 B.n381 B.n43 71.676
R725 B.n380 B.n379 71.676
R726 B.n373 B.n45 71.676
R727 B.n372 B.n371 71.676
R728 B.n364 B.n47 71.676
R729 B.n363 B.n362 71.676
R730 B.n356 B.n51 71.676
R731 B.n355 B.n354 71.676
R732 B.n348 B.n53 71.676
R733 B.n347 B.n57 71.676
R734 B.n343 B.n342 71.676
R735 B.n336 B.n59 71.676
R736 B.n335 B.n334 71.676
R737 B.n328 B.n61 71.676
R738 B.n327 B.n326 71.676
R739 B.n320 B.n63 71.676
R740 B.n319 B.n318 71.676
R741 B.n312 B.n65 71.676
R742 B.n311 B.n310 71.676
R743 B.n310 B.n309 71.676
R744 B.n313 B.n312 71.676
R745 B.n318 B.n317 71.676
R746 B.n321 B.n320 71.676
R747 B.n326 B.n325 71.676
R748 B.n329 B.n328 71.676
R749 B.n334 B.n333 71.676
R750 B.n337 B.n336 71.676
R751 B.n342 B.n341 71.676
R752 B.n344 B.n57 71.676
R753 B.n349 B.n348 71.676
R754 B.n354 B.n353 71.676
R755 B.n357 B.n356 71.676
R756 B.n362 B.n361 71.676
R757 B.n365 B.n364 71.676
R758 B.n371 B.n370 71.676
R759 B.n374 B.n373 71.676
R760 B.n379 B.n378 71.676
R761 B.n382 B.n381 71.676
R762 B.n387 B.n386 71.676
R763 B.n390 B.n389 71.676
R764 B.n395 B.n394 71.676
R765 B.n398 B.n397 71.676
R766 B.n403 B.n402 71.676
R767 B.n406 B.n405 71.676
R768 B.n227 B.n226 71.676
R769 B.n221 B.n104 71.676
R770 B.n219 B.n218 71.676
R771 B.n214 B.n213 71.676
R772 B.n211 B.n210 71.676
R773 B.n206 B.n205 71.676
R774 B.n203 B.n202 71.676
R775 B.n198 B.n197 71.676
R776 B.n195 B.n194 71.676
R777 B.n189 B.n188 71.676
R778 B.n186 B.n185 71.676
R779 B.n181 B.n180 71.676
R780 B.n178 B.n177 71.676
R781 B.n173 B.n172 71.676
R782 B.n170 B.n169 71.676
R783 B.n165 B.n164 71.676
R784 B.n162 B.n161 71.676
R785 B.n157 B.n156 71.676
R786 B.n154 B.n153 71.676
R787 B.n149 B.n148 71.676
R788 B.n146 B.n145 71.676
R789 B.n141 B.n140 71.676
R790 B.n138 B.n137 71.676
R791 B.n133 B.n132 71.676
R792 B.n77 B.t1 70.2249
R793 B.t0 B.n436 70.2249
R794 B.n93 B.t10 61.4469
R795 B.t3 B.n420 61.4469
R796 B.n123 B.n122 59.5399
R797 B.n191 B.n114 59.5399
R798 B.n368 B.n49 59.5399
R799 B.n56 B.n55 59.5399
R800 B.n409 B.n408 32.6249
R801 B.n308 B.n307 32.6249
R802 B.n234 B.n99 32.6249
R803 B.n230 B.n229 32.6249
R804 B.n122 B.n121 32.3884
R805 B.n114 B.n113 32.3884
R806 B.n49 B.n48 32.3884
R807 B.n55 B.n54 32.3884
R808 B B.n447 18.0485
R809 B.n250 B.t10 13.1676
R810 B.n421 B.t3 13.1676
R811 B.n408 B.n407 10.6151
R812 B.n407 B.n38 10.6151
R813 B.n401 B.n38 10.6151
R814 B.n401 B.n400 10.6151
R815 B.n400 B.n399 10.6151
R816 B.n399 B.n40 10.6151
R817 B.n393 B.n40 10.6151
R818 B.n393 B.n392 10.6151
R819 B.n392 B.n391 10.6151
R820 B.n391 B.n42 10.6151
R821 B.n385 B.n42 10.6151
R822 B.n385 B.n384 10.6151
R823 B.n384 B.n383 10.6151
R824 B.n383 B.n44 10.6151
R825 B.n377 B.n44 10.6151
R826 B.n377 B.n376 10.6151
R827 B.n376 B.n375 10.6151
R828 B.n375 B.n46 10.6151
R829 B.n369 B.n46 10.6151
R830 B.n367 B.n366 10.6151
R831 B.n366 B.n50 10.6151
R832 B.n360 B.n50 10.6151
R833 B.n360 B.n359 10.6151
R834 B.n359 B.n358 10.6151
R835 B.n358 B.n52 10.6151
R836 B.n352 B.n52 10.6151
R837 B.n352 B.n351 10.6151
R838 B.n351 B.n350 10.6151
R839 B.n346 B.n345 10.6151
R840 B.n345 B.n58 10.6151
R841 B.n340 B.n58 10.6151
R842 B.n340 B.n339 10.6151
R843 B.n339 B.n338 10.6151
R844 B.n338 B.n60 10.6151
R845 B.n332 B.n60 10.6151
R846 B.n332 B.n331 10.6151
R847 B.n331 B.n330 10.6151
R848 B.n330 B.n62 10.6151
R849 B.n324 B.n62 10.6151
R850 B.n324 B.n323 10.6151
R851 B.n323 B.n322 10.6151
R852 B.n322 B.n64 10.6151
R853 B.n316 B.n64 10.6151
R854 B.n316 B.n315 10.6151
R855 B.n315 B.n314 10.6151
R856 B.n314 B.n66 10.6151
R857 B.n308 B.n66 10.6151
R858 B.n235 B.n234 10.6151
R859 B.n236 B.n235 10.6151
R860 B.n236 B.n90 10.6151
R861 B.n246 B.n90 10.6151
R862 B.n247 B.n246 10.6151
R863 B.n248 B.n247 10.6151
R864 B.n248 B.n83 10.6151
R865 B.n258 B.n83 10.6151
R866 B.n259 B.n258 10.6151
R867 B.n260 B.n259 10.6151
R868 B.n260 B.n74 10.6151
R869 B.n270 B.n74 10.6151
R870 B.n271 B.n270 10.6151
R871 B.n273 B.n271 10.6151
R872 B.n273 B.n272 10.6151
R873 B.n272 B.n67 10.6151
R874 B.n284 B.n67 10.6151
R875 B.n285 B.n284 10.6151
R876 B.n286 B.n285 10.6151
R877 B.n287 B.n286 10.6151
R878 B.n289 B.n287 10.6151
R879 B.n290 B.n289 10.6151
R880 B.n291 B.n290 10.6151
R881 B.n292 B.n291 10.6151
R882 B.n294 B.n292 10.6151
R883 B.n295 B.n294 10.6151
R884 B.n296 B.n295 10.6151
R885 B.n297 B.n296 10.6151
R886 B.n299 B.n297 10.6151
R887 B.n300 B.n299 10.6151
R888 B.n301 B.n300 10.6151
R889 B.n302 B.n301 10.6151
R890 B.n304 B.n302 10.6151
R891 B.n305 B.n304 10.6151
R892 B.n306 B.n305 10.6151
R893 B.n307 B.n306 10.6151
R894 B.n229 B.n228 10.6151
R895 B.n228 B.n103 10.6151
R896 B.n223 B.n103 10.6151
R897 B.n223 B.n222 10.6151
R898 B.n222 B.n105 10.6151
R899 B.n217 B.n105 10.6151
R900 B.n217 B.n216 10.6151
R901 B.n216 B.n215 10.6151
R902 B.n215 B.n107 10.6151
R903 B.n209 B.n107 10.6151
R904 B.n209 B.n208 10.6151
R905 B.n208 B.n207 10.6151
R906 B.n207 B.n109 10.6151
R907 B.n201 B.n109 10.6151
R908 B.n201 B.n200 10.6151
R909 B.n200 B.n199 10.6151
R910 B.n199 B.n111 10.6151
R911 B.n193 B.n111 10.6151
R912 B.n193 B.n192 10.6151
R913 B.n190 B.n115 10.6151
R914 B.n184 B.n115 10.6151
R915 B.n184 B.n183 10.6151
R916 B.n183 B.n182 10.6151
R917 B.n182 B.n117 10.6151
R918 B.n176 B.n117 10.6151
R919 B.n176 B.n175 10.6151
R920 B.n175 B.n174 10.6151
R921 B.n174 B.n119 10.6151
R922 B.n168 B.n167 10.6151
R923 B.n167 B.n166 10.6151
R924 B.n166 B.n124 10.6151
R925 B.n160 B.n124 10.6151
R926 B.n160 B.n159 10.6151
R927 B.n159 B.n158 10.6151
R928 B.n158 B.n126 10.6151
R929 B.n152 B.n126 10.6151
R930 B.n152 B.n151 10.6151
R931 B.n151 B.n150 10.6151
R932 B.n150 B.n128 10.6151
R933 B.n144 B.n128 10.6151
R934 B.n144 B.n143 10.6151
R935 B.n143 B.n142 10.6151
R936 B.n142 B.n130 10.6151
R937 B.n136 B.n130 10.6151
R938 B.n136 B.n135 10.6151
R939 B.n135 B.n134 10.6151
R940 B.n134 B.n99 10.6151
R941 B.n230 B.n95 10.6151
R942 B.n240 B.n95 10.6151
R943 B.n241 B.n240 10.6151
R944 B.n242 B.n241 10.6151
R945 B.n242 B.n87 10.6151
R946 B.n252 B.n87 10.6151
R947 B.n253 B.n252 10.6151
R948 B.n254 B.n253 10.6151
R949 B.n254 B.n79 10.6151
R950 B.n264 B.n79 10.6151
R951 B.n265 B.n264 10.6151
R952 B.n266 B.n265 10.6151
R953 B.n266 B.n71 10.6151
R954 B.n277 B.n71 10.6151
R955 B.n278 B.n277 10.6151
R956 B.n279 B.n278 10.6151
R957 B.n279 B.n0 10.6151
R958 B.n441 B.n1 10.6151
R959 B.n441 B.n440 10.6151
R960 B.n440 B.n439 10.6151
R961 B.n439 B.n10 10.6151
R962 B.n433 B.n10 10.6151
R963 B.n433 B.n432 10.6151
R964 B.n432 B.n431 10.6151
R965 B.n431 B.n17 10.6151
R966 B.n425 B.n17 10.6151
R967 B.n425 B.n424 10.6151
R968 B.n424 B.n423 10.6151
R969 B.n423 B.n24 10.6151
R970 B.n417 B.n24 10.6151
R971 B.n417 B.n416 10.6151
R972 B.n416 B.n415 10.6151
R973 B.n415 B.n31 10.6151
R974 B.n409 B.n31 10.6151
R975 B.n369 B.n368 9.36635
R976 B.n346 B.n56 9.36635
R977 B.n192 B.n191 9.36635
R978 B.n168 B.n123 9.36635
R979 B.n275 B.t1 4.38953
R980 B.n437 B.t0 4.38953
R981 B.n447 B.n0 2.81026
R982 B.n447 B.n1 2.81026
R983 B.n368 B.n367 1.24928
R984 B.n350 B.n56 1.24928
R985 B.n191 B.n190 1.24928
R986 B.n123 B.n119 1.24928
R987 VN VN.t1 231.637
R988 VN VN.t0 195.674
R989 VDD2.n41 VDD2.n23 289.615
R990 VDD2.n18 VDD2.n0 289.615
R991 VDD2.n42 VDD2.n41 185
R992 VDD2.n40 VDD2.n39 185
R993 VDD2.n27 VDD2.n26 185
R994 VDD2.n34 VDD2.n33 185
R995 VDD2.n32 VDD2.n31 185
R996 VDD2.n9 VDD2.n8 185
R997 VDD2.n11 VDD2.n10 185
R998 VDD2.n4 VDD2.n3 185
R999 VDD2.n17 VDD2.n16 185
R1000 VDD2.n19 VDD2.n18 185
R1001 VDD2.n30 VDD2.t0 147.714
R1002 VDD2.n7 VDD2.t1 147.714
R1003 VDD2.n41 VDD2.n40 104.615
R1004 VDD2.n40 VDD2.n26 104.615
R1005 VDD2.n33 VDD2.n26 104.615
R1006 VDD2.n33 VDD2.n32 104.615
R1007 VDD2.n10 VDD2.n9 104.615
R1008 VDD2.n10 VDD2.n3 104.615
R1009 VDD2.n17 VDD2.n3 104.615
R1010 VDD2.n18 VDD2.n17 104.615
R1011 VDD2.n46 VDD2.n22 83.1826
R1012 VDD2.n46 VDD2.n45 52.549
R1013 VDD2.n32 VDD2.t0 52.3082
R1014 VDD2.n9 VDD2.t1 52.3082
R1015 VDD2.n31 VDD2.n30 15.6631
R1016 VDD2.n8 VDD2.n7 15.6631
R1017 VDD2.n34 VDD2.n29 12.8005
R1018 VDD2.n11 VDD2.n6 12.8005
R1019 VDD2.n35 VDD2.n27 12.0247
R1020 VDD2.n12 VDD2.n4 12.0247
R1021 VDD2.n39 VDD2.n38 11.249
R1022 VDD2.n16 VDD2.n15 11.249
R1023 VDD2.n42 VDD2.n25 10.4732
R1024 VDD2.n19 VDD2.n2 10.4732
R1025 VDD2.n43 VDD2.n23 9.69747
R1026 VDD2.n20 VDD2.n0 9.69747
R1027 VDD2.n45 VDD2.n44 9.45567
R1028 VDD2.n22 VDD2.n21 9.45567
R1029 VDD2.n44 VDD2.n43 9.3005
R1030 VDD2.n25 VDD2.n24 9.3005
R1031 VDD2.n38 VDD2.n37 9.3005
R1032 VDD2.n36 VDD2.n35 9.3005
R1033 VDD2.n29 VDD2.n28 9.3005
R1034 VDD2.n21 VDD2.n20 9.3005
R1035 VDD2.n2 VDD2.n1 9.3005
R1036 VDD2.n15 VDD2.n14 9.3005
R1037 VDD2.n13 VDD2.n12 9.3005
R1038 VDD2.n6 VDD2.n5 9.3005
R1039 VDD2.n30 VDD2.n28 4.39059
R1040 VDD2.n7 VDD2.n5 4.39059
R1041 VDD2.n45 VDD2.n23 4.26717
R1042 VDD2.n22 VDD2.n0 4.26717
R1043 VDD2.n43 VDD2.n42 3.49141
R1044 VDD2.n20 VDD2.n19 3.49141
R1045 VDD2.n39 VDD2.n25 2.71565
R1046 VDD2.n16 VDD2.n2 2.71565
R1047 VDD2.n38 VDD2.n27 1.93989
R1048 VDD2.n15 VDD2.n4 1.93989
R1049 VDD2.n35 VDD2.n34 1.16414
R1050 VDD2.n12 VDD2.n11 1.16414
R1051 VDD2 VDD2.n46 0.418603
R1052 VDD2.n31 VDD2.n29 0.388379
R1053 VDD2.n8 VDD2.n6 0.388379
R1054 VDD2.n44 VDD2.n24 0.155672
R1055 VDD2.n37 VDD2.n24 0.155672
R1056 VDD2.n37 VDD2.n36 0.155672
R1057 VDD2.n36 VDD2.n28 0.155672
R1058 VDD2.n13 VDD2.n5 0.155672
R1059 VDD2.n14 VDD2.n13 0.155672
R1060 VDD2.n14 VDD2.n1 0.155672
R1061 VDD2.n21 VDD2.n1 0.155672
C0 VP VDD2 0.283596f
C1 VP VN 3.52183f
C2 VDD1 VDD2 0.527025f
C3 VDD1 VN 0.151408f
C4 VDD2 VTAIL 2.94218f
C5 VTAIL VN 1.06452f
C6 VP VDD1 1.24051f
C7 VDD2 VN 1.11017f
C8 VP VTAIL 1.07876f
C9 VDD1 VTAIL 2.89918f
C10 VDD2 B 2.650861f
C11 VDD1 B 4.04157f
C12 VTAIL B 3.715207f
C13 VN B 6.36095f
C14 VP B 4.237451f
C15 VDD2.n0 B 0.022175f
C16 VDD2.n1 B 0.014985f
C17 VDD2.n2 B 0.008052f
C18 VDD2.n3 B 0.019033f
C19 VDD2.n4 B 0.008526f
C20 VDD2.n5 B 0.269578f
C21 VDD2.n6 B 0.008052f
C22 VDD2.t1 B 0.031349f
C23 VDD2.n7 B 0.060176f
C24 VDD2.n8 B 0.011232f
C25 VDD2.n9 B 0.014275f
C26 VDD2.n10 B 0.019033f
C27 VDD2.n11 B 0.008526f
C28 VDD2.n12 B 0.008052f
C29 VDD2.n13 B 0.014985f
C30 VDD2.n14 B 0.014985f
C31 VDD2.n15 B 0.008052f
C32 VDD2.n16 B 0.008526f
C33 VDD2.n17 B 0.019033f
C34 VDD2.n18 B 0.043169f
C35 VDD2.n19 B 0.008526f
C36 VDD2.n20 B 0.008052f
C37 VDD2.n21 B 0.038526f
C38 VDD2.n22 B 0.248195f
C39 VDD2.n23 B 0.022175f
C40 VDD2.n24 B 0.014985f
C41 VDD2.n25 B 0.008052f
C42 VDD2.n26 B 0.019033f
C43 VDD2.n27 B 0.008526f
C44 VDD2.n28 B 0.269578f
C45 VDD2.n29 B 0.008052f
C46 VDD2.t0 B 0.031349f
C47 VDD2.n30 B 0.060176f
C48 VDD2.n31 B 0.011232f
C49 VDD2.n32 B 0.014275f
C50 VDD2.n33 B 0.019033f
C51 VDD2.n34 B 0.008526f
C52 VDD2.n35 B 0.008052f
C53 VDD2.n36 B 0.014985f
C54 VDD2.n37 B 0.014985f
C55 VDD2.n38 B 0.008052f
C56 VDD2.n39 B 0.008526f
C57 VDD2.n40 B 0.019033f
C58 VDD2.n41 B 0.043169f
C59 VDD2.n42 B 0.008526f
C60 VDD2.n43 B 0.008052f
C61 VDD2.n44 B 0.038526f
C62 VDD2.n45 B 0.034791f
C63 VDD2.n46 B 1.22786f
C64 VN.t0 B 0.642263f
C65 VN.t1 B 0.812008f
C66 VDD1.n0 B 0.02176f
C67 VDD1.n1 B 0.014704f
C68 VDD1.n2 B 0.007901f
C69 VDD1.n3 B 0.018676f
C70 VDD1.n4 B 0.008366f
C71 VDD1.n5 B 0.26453f
C72 VDD1.n6 B 0.007901f
C73 VDD1.t1 B 0.030762f
C74 VDD1.n7 B 0.059049f
C75 VDD1.n8 B 0.011022f
C76 VDD1.n9 B 0.014007f
C77 VDD1.n10 B 0.018676f
C78 VDD1.n11 B 0.008366f
C79 VDD1.n12 B 0.007901f
C80 VDD1.n13 B 0.014704f
C81 VDD1.n14 B 0.014704f
C82 VDD1.n15 B 0.007901f
C83 VDD1.n16 B 0.008366f
C84 VDD1.n17 B 0.018676f
C85 VDD1.n18 B 0.042361f
C86 VDD1.n19 B 0.008366f
C87 VDD1.n20 B 0.007901f
C88 VDD1.n21 B 0.037805f
C89 VDD1.n22 B 0.034536f
C90 VDD1.n23 B 0.02176f
C91 VDD1.n24 B 0.014704f
C92 VDD1.n25 B 0.007901f
C93 VDD1.n26 B 0.018676f
C94 VDD1.n27 B 0.008366f
C95 VDD1.n28 B 0.26453f
C96 VDD1.n29 B 0.007901f
C97 VDD1.t0 B 0.030762f
C98 VDD1.n30 B 0.059049f
C99 VDD1.n31 B 0.011022f
C100 VDD1.n32 B 0.014007f
C101 VDD1.n33 B 0.018676f
C102 VDD1.n34 B 0.008366f
C103 VDD1.n35 B 0.007901f
C104 VDD1.n36 B 0.014704f
C105 VDD1.n37 B 0.014704f
C106 VDD1.n38 B 0.007901f
C107 VDD1.n39 B 0.008366f
C108 VDD1.n40 B 0.018676f
C109 VDD1.n41 B 0.042361f
C110 VDD1.n42 B 0.008366f
C111 VDD1.n43 B 0.007901f
C112 VDD1.n44 B 0.037805f
C113 VDD1.n45 B 0.262176f
C114 VTAIL.n0 B 0.025331f
C115 VTAIL.n1 B 0.017118f
C116 VTAIL.n2 B 0.009198f
C117 VTAIL.n3 B 0.021741f
C118 VTAIL.n4 B 0.009739f
C119 VTAIL.n5 B 0.307943f
C120 VTAIL.n6 B 0.009198f
C121 VTAIL.t3 B 0.03581f
C122 VTAIL.n7 B 0.06874f
C123 VTAIL.n8 B 0.01283f
C124 VTAIL.n9 B 0.016306f
C125 VTAIL.n10 B 0.021741f
C126 VTAIL.n11 B 0.009739f
C127 VTAIL.n12 B 0.009198f
C128 VTAIL.n13 B 0.017118f
C129 VTAIL.n14 B 0.017118f
C130 VTAIL.n15 B 0.009198f
C131 VTAIL.n16 B 0.009739f
C132 VTAIL.n17 B 0.021741f
C133 VTAIL.n18 B 0.049313f
C134 VTAIL.n19 B 0.009739f
C135 VTAIL.n20 B 0.009198f
C136 VTAIL.n21 B 0.044009f
C137 VTAIL.n22 B 0.027953f
C138 VTAIL.n23 B 0.6833f
C139 VTAIL.n24 B 0.025331f
C140 VTAIL.n25 B 0.017118f
C141 VTAIL.n26 B 0.009198f
C142 VTAIL.n27 B 0.021741f
C143 VTAIL.n28 B 0.009739f
C144 VTAIL.n29 B 0.307943f
C145 VTAIL.n30 B 0.009198f
C146 VTAIL.t1 B 0.03581f
C147 VTAIL.n31 B 0.06874f
C148 VTAIL.n32 B 0.01283f
C149 VTAIL.n33 B 0.016306f
C150 VTAIL.n34 B 0.021741f
C151 VTAIL.n35 B 0.009739f
C152 VTAIL.n36 B 0.009198f
C153 VTAIL.n37 B 0.017118f
C154 VTAIL.n38 B 0.017118f
C155 VTAIL.n39 B 0.009198f
C156 VTAIL.n40 B 0.009739f
C157 VTAIL.n41 B 0.021741f
C158 VTAIL.n42 B 0.049313f
C159 VTAIL.n43 B 0.009739f
C160 VTAIL.n44 B 0.009198f
C161 VTAIL.n45 B 0.044009f
C162 VTAIL.n46 B 0.027953f
C163 VTAIL.n47 B 0.699942f
C164 VTAIL.n48 B 0.025331f
C165 VTAIL.n49 B 0.017118f
C166 VTAIL.n50 B 0.009198f
C167 VTAIL.n51 B 0.021741f
C168 VTAIL.n52 B 0.009739f
C169 VTAIL.n53 B 0.307943f
C170 VTAIL.n54 B 0.009198f
C171 VTAIL.t2 B 0.03581f
C172 VTAIL.n55 B 0.06874f
C173 VTAIL.n56 B 0.01283f
C174 VTAIL.n57 B 0.016306f
C175 VTAIL.n58 B 0.021741f
C176 VTAIL.n59 B 0.009739f
C177 VTAIL.n60 B 0.009198f
C178 VTAIL.n61 B 0.017118f
C179 VTAIL.n62 B 0.017118f
C180 VTAIL.n63 B 0.009198f
C181 VTAIL.n64 B 0.009739f
C182 VTAIL.n65 B 0.021741f
C183 VTAIL.n66 B 0.049313f
C184 VTAIL.n67 B 0.009739f
C185 VTAIL.n68 B 0.009198f
C186 VTAIL.n69 B 0.044009f
C187 VTAIL.n70 B 0.027953f
C188 VTAIL.n71 B 0.620536f
C189 VTAIL.n72 B 0.025331f
C190 VTAIL.n73 B 0.017118f
C191 VTAIL.n74 B 0.009198f
C192 VTAIL.n75 B 0.021741f
C193 VTAIL.n76 B 0.009739f
C194 VTAIL.n77 B 0.307943f
C195 VTAIL.n78 B 0.009198f
C196 VTAIL.t0 B 0.03581f
C197 VTAIL.n79 B 0.06874f
C198 VTAIL.n80 B 0.01283f
C199 VTAIL.n81 B 0.016306f
C200 VTAIL.n82 B 0.021741f
C201 VTAIL.n83 B 0.009739f
C202 VTAIL.n84 B 0.009198f
C203 VTAIL.n85 B 0.017118f
C204 VTAIL.n86 B 0.017118f
C205 VTAIL.n87 B 0.009198f
C206 VTAIL.n88 B 0.009739f
C207 VTAIL.n89 B 0.021741f
C208 VTAIL.n90 B 0.049313f
C209 VTAIL.n91 B 0.009739f
C210 VTAIL.n92 B 0.009198f
C211 VTAIL.n93 B 0.044009f
C212 VTAIL.n94 B 0.027953f
C213 VTAIL.n95 B 0.571561f
C214 VP.t0 B 0.817753f
C215 VP.t1 B 0.649633f
C216 VP.n0 B 2.00526f
.ends

