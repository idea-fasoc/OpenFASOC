* NGSPICE file created from diff_pair_sample_0790.ext - technology: sky130A

.subckt diff_pair_sample_0790 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t6 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=5.0544 ps=26.7 w=12.96 l=1.39
X1 B.t11 B.t9 B.t10 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=0 ps=0 w=12.96 l=1.39
X2 VTAIL.t5 VN.t0 VDD2.t5 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=2.1384 ps=13.29 w=12.96 l=1.39
X3 VDD2.t4 VN.t1 VTAIL.t2 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=2.1384 ps=13.29 w=12.96 l=1.39
X4 VDD1.t4 VP.t1 VTAIL.t10 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=2.1384 ps=13.29 w=12.96 l=1.39
X5 VDD1.t3 VP.t2 VTAIL.t8 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=5.0544 ps=26.7 w=12.96 l=1.39
X6 VTAIL.t9 VP.t3 VDD1.t2 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=2.1384 ps=13.29 w=12.96 l=1.39
X7 VDD2.t3 VN.t2 VTAIL.t3 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=2.1384 ps=13.29 w=12.96 l=1.39
X8 VDD2.t2 VN.t3 VTAIL.t4 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=5.0544 ps=26.7 w=12.96 l=1.39
X9 B.t8 B.t6 B.t7 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=0 ps=0 w=12.96 l=1.39
X10 VDD2.t1 VN.t4 VTAIL.t1 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=5.0544 ps=26.7 w=12.96 l=1.39
X11 VDD1.t1 VP.t4 VTAIL.t11 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=2.1384 ps=13.29 w=12.96 l=1.39
X12 VTAIL.t7 VP.t5 VDD1.t0 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=2.1384 ps=13.29 w=12.96 l=1.39
X13 B.t5 B.t3 B.t4 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=0 ps=0 w=12.96 l=1.39
X14 B.t2 B.t0 B.t1 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=5.0544 pd=26.7 as=0 ps=0 w=12.96 l=1.39
X15 VTAIL.t0 VN.t5 VDD2.t0 w_n2346_n3560# sky130_fd_pr__pfet_01v8 ad=2.1384 pd=13.29 as=2.1384 ps=13.29 w=12.96 l=1.39
R0 VP.n7 VP.t4 259.094
R1 VP.n20 VP.t5 224.702
R2 VP.n14 VP.t1 224.702
R3 VP.n26 VP.t0 224.702
R4 VP.n6 VP.t3 224.702
R5 VP.n12 VP.t2 224.702
R6 VP.n15 VP.n14 174.933
R7 VP.n27 VP.n26 174.933
R8 VP.n13 VP.n12 174.933
R9 VP.n8 VP.n5 161.3
R10 VP.n10 VP.n9 161.3
R11 VP.n11 VP.n4 161.3
R12 VP.n25 VP.n0 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n22 VP.n1 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n19 VP.n2 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n3 161.3
R19 VP.n19 VP.n18 54.0429
R20 VP.n24 VP.n1 54.0429
R21 VP.n10 VP.n5 54.0429
R22 VP.n15 VP.n13 44.5687
R23 VP.n7 VP.n6 41.7088
R24 VP.n18 VP.n3 26.7783
R25 VP.n25 VP.n24 26.7783
R26 VP.n11 VP.n10 26.7783
R27 VP.n20 VP.n19 24.3439
R28 VP.n20 VP.n1 24.3439
R29 VP.n6 VP.n5 24.3439
R30 VP.n8 VP.n7 17.7134
R31 VP.n14 VP.n3 10.7116
R32 VP.n26 VP.n25 10.7116
R33 VP.n12 VP.n11 10.7116
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n4 0.189894
R36 VP.n13 VP.n4 0.189894
R37 VP.n16 VP.n15 0.189894
R38 VP.n17 VP.n16 0.189894
R39 VP.n17 VP.n2 0.189894
R40 VP.n21 VP.n2 0.189894
R41 VP.n22 VP.n21 0.189894
R42 VP.n23 VP.n22 0.189894
R43 VP.n23 VP.n0 0.189894
R44 VP.n27 VP.n0 0.189894
R45 VP VP.n27 0.0516364
R46 VTAIL.n7 VTAIL.t4 60.4663
R47 VTAIL.n11 VTAIL.t1 60.4652
R48 VTAIL.n2 VTAIL.t6 60.4652
R49 VTAIL.n10 VTAIL.t8 60.4652
R50 VTAIL.n9 VTAIL.n8 57.9583
R51 VTAIL.n6 VTAIL.n5 57.9583
R52 VTAIL.n1 VTAIL.n0 57.9571
R53 VTAIL.n4 VTAIL.n3 57.9571
R54 VTAIL.n6 VTAIL.n4 26.5048
R55 VTAIL.n11 VTAIL.n10 25.0221
R56 VTAIL.n0 VTAIL.t3 2.5086
R57 VTAIL.n0 VTAIL.t0 2.5086
R58 VTAIL.n3 VTAIL.t10 2.5086
R59 VTAIL.n3 VTAIL.t7 2.5086
R60 VTAIL.n8 VTAIL.t11 2.5086
R61 VTAIL.n8 VTAIL.t9 2.5086
R62 VTAIL.n5 VTAIL.t2 2.5086
R63 VTAIL.n5 VTAIL.t5 2.5086
R64 VTAIL.n7 VTAIL.n6 1.48326
R65 VTAIL.n10 VTAIL.n9 1.48326
R66 VTAIL.n4 VTAIL.n2 1.48326
R67 VTAIL.n9 VTAIL.n7 1.21171
R68 VTAIL.n2 VTAIL.n1 1.21171
R69 VTAIL VTAIL.n11 1.05438
R70 VTAIL VTAIL.n1 0.429379
R71 VDD1 VDD1.t1 78.3154
R72 VDD1.n1 VDD1.t4 78.2007
R73 VDD1.n1 VDD1.n0 74.9512
R74 VDD1.n3 VDD1.n2 74.6359
R75 VDD1.n3 VDD1.n1 41.0311
R76 VDD1.n2 VDD1.t2 2.5086
R77 VDD1.n2 VDD1.t3 2.5086
R78 VDD1.n0 VDD1.t0 2.5086
R79 VDD1.n0 VDD1.t5 2.5086
R80 VDD1 VDD1.n3 0.313
R81 B.n354 B.n353 585
R82 B.n352 B.n99 585
R83 B.n351 B.n350 585
R84 B.n349 B.n100 585
R85 B.n348 B.n347 585
R86 B.n346 B.n101 585
R87 B.n345 B.n344 585
R88 B.n343 B.n102 585
R89 B.n342 B.n341 585
R90 B.n340 B.n103 585
R91 B.n339 B.n338 585
R92 B.n337 B.n104 585
R93 B.n336 B.n335 585
R94 B.n334 B.n105 585
R95 B.n333 B.n332 585
R96 B.n331 B.n106 585
R97 B.n330 B.n329 585
R98 B.n328 B.n107 585
R99 B.n327 B.n326 585
R100 B.n325 B.n108 585
R101 B.n324 B.n323 585
R102 B.n322 B.n109 585
R103 B.n321 B.n320 585
R104 B.n319 B.n110 585
R105 B.n318 B.n317 585
R106 B.n316 B.n111 585
R107 B.n315 B.n314 585
R108 B.n313 B.n112 585
R109 B.n312 B.n311 585
R110 B.n310 B.n113 585
R111 B.n309 B.n308 585
R112 B.n307 B.n114 585
R113 B.n306 B.n305 585
R114 B.n304 B.n115 585
R115 B.n303 B.n302 585
R116 B.n301 B.n116 585
R117 B.n300 B.n299 585
R118 B.n298 B.n117 585
R119 B.n297 B.n296 585
R120 B.n295 B.n118 585
R121 B.n294 B.n293 585
R122 B.n292 B.n119 585
R123 B.n291 B.n290 585
R124 B.n289 B.n120 585
R125 B.n288 B.n287 585
R126 B.n283 B.n121 585
R127 B.n282 B.n281 585
R128 B.n280 B.n122 585
R129 B.n279 B.n278 585
R130 B.n277 B.n123 585
R131 B.n276 B.n275 585
R132 B.n274 B.n124 585
R133 B.n273 B.n272 585
R134 B.n271 B.n125 585
R135 B.n269 B.n268 585
R136 B.n267 B.n128 585
R137 B.n266 B.n265 585
R138 B.n264 B.n129 585
R139 B.n263 B.n262 585
R140 B.n261 B.n130 585
R141 B.n260 B.n259 585
R142 B.n258 B.n131 585
R143 B.n257 B.n256 585
R144 B.n255 B.n132 585
R145 B.n254 B.n253 585
R146 B.n252 B.n133 585
R147 B.n251 B.n250 585
R148 B.n249 B.n134 585
R149 B.n248 B.n247 585
R150 B.n246 B.n135 585
R151 B.n245 B.n244 585
R152 B.n243 B.n136 585
R153 B.n242 B.n241 585
R154 B.n240 B.n137 585
R155 B.n239 B.n238 585
R156 B.n237 B.n138 585
R157 B.n236 B.n235 585
R158 B.n234 B.n139 585
R159 B.n233 B.n232 585
R160 B.n231 B.n140 585
R161 B.n230 B.n229 585
R162 B.n228 B.n141 585
R163 B.n227 B.n226 585
R164 B.n225 B.n142 585
R165 B.n224 B.n223 585
R166 B.n222 B.n143 585
R167 B.n221 B.n220 585
R168 B.n219 B.n144 585
R169 B.n218 B.n217 585
R170 B.n216 B.n145 585
R171 B.n215 B.n214 585
R172 B.n213 B.n146 585
R173 B.n212 B.n211 585
R174 B.n210 B.n147 585
R175 B.n209 B.n208 585
R176 B.n207 B.n148 585
R177 B.n206 B.n205 585
R178 B.n204 B.n149 585
R179 B.n355 B.n98 585
R180 B.n357 B.n356 585
R181 B.n358 B.n97 585
R182 B.n360 B.n359 585
R183 B.n361 B.n96 585
R184 B.n363 B.n362 585
R185 B.n364 B.n95 585
R186 B.n366 B.n365 585
R187 B.n367 B.n94 585
R188 B.n369 B.n368 585
R189 B.n370 B.n93 585
R190 B.n372 B.n371 585
R191 B.n373 B.n92 585
R192 B.n375 B.n374 585
R193 B.n376 B.n91 585
R194 B.n378 B.n377 585
R195 B.n379 B.n90 585
R196 B.n381 B.n380 585
R197 B.n382 B.n89 585
R198 B.n384 B.n383 585
R199 B.n385 B.n88 585
R200 B.n387 B.n386 585
R201 B.n388 B.n87 585
R202 B.n390 B.n389 585
R203 B.n391 B.n86 585
R204 B.n393 B.n392 585
R205 B.n394 B.n85 585
R206 B.n396 B.n395 585
R207 B.n397 B.n84 585
R208 B.n399 B.n398 585
R209 B.n400 B.n83 585
R210 B.n402 B.n401 585
R211 B.n403 B.n82 585
R212 B.n405 B.n404 585
R213 B.n406 B.n81 585
R214 B.n408 B.n407 585
R215 B.n409 B.n80 585
R216 B.n411 B.n410 585
R217 B.n412 B.n79 585
R218 B.n414 B.n413 585
R219 B.n415 B.n78 585
R220 B.n417 B.n416 585
R221 B.n418 B.n77 585
R222 B.n420 B.n419 585
R223 B.n421 B.n76 585
R224 B.n423 B.n422 585
R225 B.n424 B.n75 585
R226 B.n426 B.n425 585
R227 B.n427 B.n74 585
R228 B.n429 B.n428 585
R229 B.n430 B.n73 585
R230 B.n432 B.n431 585
R231 B.n433 B.n72 585
R232 B.n435 B.n434 585
R233 B.n436 B.n71 585
R234 B.n438 B.n437 585
R235 B.n439 B.n70 585
R236 B.n441 B.n440 585
R237 B.n589 B.n16 585
R238 B.n588 B.n587 585
R239 B.n586 B.n17 585
R240 B.n585 B.n584 585
R241 B.n583 B.n18 585
R242 B.n582 B.n581 585
R243 B.n580 B.n19 585
R244 B.n579 B.n578 585
R245 B.n577 B.n20 585
R246 B.n576 B.n575 585
R247 B.n574 B.n21 585
R248 B.n573 B.n572 585
R249 B.n571 B.n22 585
R250 B.n570 B.n569 585
R251 B.n568 B.n23 585
R252 B.n567 B.n566 585
R253 B.n565 B.n24 585
R254 B.n564 B.n563 585
R255 B.n562 B.n25 585
R256 B.n561 B.n560 585
R257 B.n559 B.n26 585
R258 B.n558 B.n557 585
R259 B.n556 B.n27 585
R260 B.n555 B.n554 585
R261 B.n553 B.n28 585
R262 B.n552 B.n551 585
R263 B.n550 B.n29 585
R264 B.n549 B.n548 585
R265 B.n547 B.n30 585
R266 B.n546 B.n545 585
R267 B.n544 B.n31 585
R268 B.n543 B.n542 585
R269 B.n541 B.n32 585
R270 B.n540 B.n539 585
R271 B.n538 B.n33 585
R272 B.n537 B.n536 585
R273 B.n535 B.n34 585
R274 B.n534 B.n533 585
R275 B.n532 B.n35 585
R276 B.n531 B.n530 585
R277 B.n529 B.n36 585
R278 B.n528 B.n527 585
R279 B.n526 B.n37 585
R280 B.n525 B.n524 585
R281 B.n523 B.n522 585
R282 B.n521 B.n41 585
R283 B.n520 B.n519 585
R284 B.n518 B.n42 585
R285 B.n517 B.n516 585
R286 B.n515 B.n43 585
R287 B.n514 B.n513 585
R288 B.n512 B.n44 585
R289 B.n511 B.n510 585
R290 B.n509 B.n45 585
R291 B.n507 B.n506 585
R292 B.n505 B.n48 585
R293 B.n504 B.n503 585
R294 B.n502 B.n49 585
R295 B.n501 B.n500 585
R296 B.n499 B.n50 585
R297 B.n498 B.n497 585
R298 B.n496 B.n51 585
R299 B.n495 B.n494 585
R300 B.n493 B.n52 585
R301 B.n492 B.n491 585
R302 B.n490 B.n53 585
R303 B.n489 B.n488 585
R304 B.n487 B.n54 585
R305 B.n486 B.n485 585
R306 B.n484 B.n55 585
R307 B.n483 B.n482 585
R308 B.n481 B.n56 585
R309 B.n480 B.n479 585
R310 B.n478 B.n57 585
R311 B.n477 B.n476 585
R312 B.n475 B.n58 585
R313 B.n474 B.n473 585
R314 B.n472 B.n59 585
R315 B.n471 B.n470 585
R316 B.n469 B.n60 585
R317 B.n468 B.n467 585
R318 B.n466 B.n61 585
R319 B.n465 B.n464 585
R320 B.n463 B.n62 585
R321 B.n462 B.n461 585
R322 B.n460 B.n63 585
R323 B.n459 B.n458 585
R324 B.n457 B.n64 585
R325 B.n456 B.n455 585
R326 B.n454 B.n65 585
R327 B.n453 B.n452 585
R328 B.n451 B.n66 585
R329 B.n450 B.n449 585
R330 B.n448 B.n67 585
R331 B.n447 B.n446 585
R332 B.n445 B.n68 585
R333 B.n444 B.n443 585
R334 B.n442 B.n69 585
R335 B.n591 B.n590 585
R336 B.n592 B.n15 585
R337 B.n594 B.n593 585
R338 B.n595 B.n14 585
R339 B.n597 B.n596 585
R340 B.n598 B.n13 585
R341 B.n600 B.n599 585
R342 B.n601 B.n12 585
R343 B.n603 B.n602 585
R344 B.n604 B.n11 585
R345 B.n606 B.n605 585
R346 B.n607 B.n10 585
R347 B.n609 B.n608 585
R348 B.n610 B.n9 585
R349 B.n612 B.n611 585
R350 B.n613 B.n8 585
R351 B.n615 B.n614 585
R352 B.n616 B.n7 585
R353 B.n618 B.n617 585
R354 B.n619 B.n6 585
R355 B.n621 B.n620 585
R356 B.n622 B.n5 585
R357 B.n624 B.n623 585
R358 B.n625 B.n4 585
R359 B.n627 B.n626 585
R360 B.n628 B.n3 585
R361 B.n630 B.n629 585
R362 B.n631 B.n0 585
R363 B.n2 B.n1 585
R364 B.n164 B.n163 585
R365 B.n165 B.n162 585
R366 B.n167 B.n166 585
R367 B.n168 B.n161 585
R368 B.n170 B.n169 585
R369 B.n171 B.n160 585
R370 B.n173 B.n172 585
R371 B.n174 B.n159 585
R372 B.n176 B.n175 585
R373 B.n177 B.n158 585
R374 B.n179 B.n178 585
R375 B.n180 B.n157 585
R376 B.n182 B.n181 585
R377 B.n183 B.n156 585
R378 B.n185 B.n184 585
R379 B.n186 B.n155 585
R380 B.n188 B.n187 585
R381 B.n189 B.n154 585
R382 B.n191 B.n190 585
R383 B.n192 B.n153 585
R384 B.n194 B.n193 585
R385 B.n195 B.n152 585
R386 B.n197 B.n196 585
R387 B.n198 B.n151 585
R388 B.n200 B.n199 585
R389 B.n201 B.n150 585
R390 B.n203 B.n202 585
R391 B.n202 B.n149 511.721
R392 B.n355 B.n354 511.721
R393 B.n440 B.n69 511.721
R394 B.n590 B.n589 511.721
R395 B.n126 B.t0 429.707
R396 B.n284 B.t9 429.707
R397 B.n46 B.t6 429.707
R398 B.n38 B.t3 429.707
R399 B.n633 B.n632 256.663
R400 B.n632 B.n631 235.042
R401 B.n632 B.n2 235.042
R402 B.n206 B.n149 163.367
R403 B.n207 B.n206 163.367
R404 B.n208 B.n207 163.367
R405 B.n208 B.n147 163.367
R406 B.n212 B.n147 163.367
R407 B.n213 B.n212 163.367
R408 B.n214 B.n213 163.367
R409 B.n214 B.n145 163.367
R410 B.n218 B.n145 163.367
R411 B.n219 B.n218 163.367
R412 B.n220 B.n219 163.367
R413 B.n220 B.n143 163.367
R414 B.n224 B.n143 163.367
R415 B.n225 B.n224 163.367
R416 B.n226 B.n225 163.367
R417 B.n226 B.n141 163.367
R418 B.n230 B.n141 163.367
R419 B.n231 B.n230 163.367
R420 B.n232 B.n231 163.367
R421 B.n232 B.n139 163.367
R422 B.n236 B.n139 163.367
R423 B.n237 B.n236 163.367
R424 B.n238 B.n237 163.367
R425 B.n238 B.n137 163.367
R426 B.n242 B.n137 163.367
R427 B.n243 B.n242 163.367
R428 B.n244 B.n243 163.367
R429 B.n244 B.n135 163.367
R430 B.n248 B.n135 163.367
R431 B.n249 B.n248 163.367
R432 B.n250 B.n249 163.367
R433 B.n250 B.n133 163.367
R434 B.n254 B.n133 163.367
R435 B.n255 B.n254 163.367
R436 B.n256 B.n255 163.367
R437 B.n256 B.n131 163.367
R438 B.n260 B.n131 163.367
R439 B.n261 B.n260 163.367
R440 B.n262 B.n261 163.367
R441 B.n262 B.n129 163.367
R442 B.n266 B.n129 163.367
R443 B.n267 B.n266 163.367
R444 B.n268 B.n267 163.367
R445 B.n268 B.n125 163.367
R446 B.n273 B.n125 163.367
R447 B.n274 B.n273 163.367
R448 B.n275 B.n274 163.367
R449 B.n275 B.n123 163.367
R450 B.n279 B.n123 163.367
R451 B.n280 B.n279 163.367
R452 B.n281 B.n280 163.367
R453 B.n281 B.n121 163.367
R454 B.n288 B.n121 163.367
R455 B.n289 B.n288 163.367
R456 B.n290 B.n289 163.367
R457 B.n290 B.n119 163.367
R458 B.n294 B.n119 163.367
R459 B.n295 B.n294 163.367
R460 B.n296 B.n295 163.367
R461 B.n296 B.n117 163.367
R462 B.n300 B.n117 163.367
R463 B.n301 B.n300 163.367
R464 B.n302 B.n301 163.367
R465 B.n302 B.n115 163.367
R466 B.n306 B.n115 163.367
R467 B.n307 B.n306 163.367
R468 B.n308 B.n307 163.367
R469 B.n308 B.n113 163.367
R470 B.n312 B.n113 163.367
R471 B.n313 B.n312 163.367
R472 B.n314 B.n313 163.367
R473 B.n314 B.n111 163.367
R474 B.n318 B.n111 163.367
R475 B.n319 B.n318 163.367
R476 B.n320 B.n319 163.367
R477 B.n320 B.n109 163.367
R478 B.n324 B.n109 163.367
R479 B.n325 B.n324 163.367
R480 B.n326 B.n325 163.367
R481 B.n326 B.n107 163.367
R482 B.n330 B.n107 163.367
R483 B.n331 B.n330 163.367
R484 B.n332 B.n331 163.367
R485 B.n332 B.n105 163.367
R486 B.n336 B.n105 163.367
R487 B.n337 B.n336 163.367
R488 B.n338 B.n337 163.367
R489 B.n338 B.n103 163.367
R490 B.n342 B.n103 163.367
R491 B.n343 B.n342 163.367
R492 B.n344 B.n343 163.367
R493 B.n344 B.n101 163.367
R494 B.n348 B.n101 163.367
R495 B.n349 B.n348 163.367
R496 B.n350 B.n349 163.367
R497 B.n350 B.n99 163.367
R498 B.n354 B.n99 163.367
R499 B.n440 B.n439 163.367
R500 B.n439 B.n438 163.367
R501 B.n438 B.n71 163.367
R502 B.n434 B.n71 163.367
R503 B.n434 B.n433 163.367
R504 B.n433 B.n432 163.367
R505 B.n432 B.n73 163.367
R506 B.n428 B.n73 163.367
R507 B.n428 B.n427 163.367
R508 B.n427 B.n426 163.367
R509 B.n426 B.n75 163.367
R510 B.n422 B.n75 163.367
R511 B.n422 B.n421 163.367
R512 B.n421 B.n420 163.367
R513 B.n420 B.n77 163.367
R514 B.n416 B.n77 163.367
R515 B.n416 B.n415 163.367
R516 B.n415 B.n414 163.367
R517 B.n414 B.n79 163.367
R518 B.n410 B.n79 163.367
R519 B.n410 B.n409 163.367
R520 B.n409 B.n408 163.367
R521 B.n408 B.n81 163.367
R522 B.n404 B.n81 163.367
R523 B.n404 B.n403 163.367
R524 B.n403 B.n402 163.367
R525 B.n402 B.n83 163.367
R526 B.n398 B.n83 163.367
R527 B.n398 B.n397 163.367
R528 B.n397 B.n396 163.367
R529 B.n396 B.n85 163.367
R530 B.n392 B.n85 163.367
R531 B.n392 B.n391 163.367
R532 B.n391 B.n390 163.367
R533 B.n390 B.n87 163.367
R534 B.n386 B.n87 163.367
R535 B.n386 B.n385 163.367
R536 B.n385 B.n384 163.367
R537 B.n384 B.n89 163.367
R538 B.n380 B.n89 163.367
R539 B.n380 B.n379 163.367
R540 B.n379 B.n378 163.367
R541 B.n378 B.n91 163.367
R542 B.n374 B.n91 163.367
R543 B.n374 B.n373 163.367
R544 B.n373 B.n372 163.367
R545 B.n372 B.n93 163.367
R546 B.n368 B.n93 163.367
R547 B.n368 B.n367 163.367
R548 B.n367 B.n366 163.367
R549 B.n366 B.n95 163.367
R550 B.n362 B.n95 163.367
R551 B.n362 B.n361 163.367
R552 B.n361 B.n360 163.367
R553 B.n360 B.n97 163.367
R554 B.n356 B.n97 163.367
R555 B.n356 B.n355 163.367
R556 B.n589 B.n588 163.367
R557 B.n588 B.n17 163.367
R558 B.n584 B.n17 163.367
R559 B.n584 B.n583 163.367
R560 B.n583 B.n582 163.367
R561 B.n582 B.n19 163.367
R562 B.n578 B.n19 163.367
R563 B.n578 B.n577 163.367
R564 B.n577 B.n576 163.367
R565 B.n576 B.n21 163.367
R566 B.n572 B.n21 163.367
R567 B.n572 B.n571 163.367
R568 B.n571 B.n570 163.367
R569 B.n570 B.n23 163.367
R570 B.n566 B.n23 163.367
R571 B.n566 B.n565 163.367
R572 B.n565 B.n564 163.367
R573 B.n564 B.n25 163.367
R574 B.n560 B.n25 163.367
R575 B.n560 B.n559 163.367
R576 B.n559 B.n558 163.367
R577 B.n558 B.n27 163.367
R578 B.n554 B.n27 163.367
R579 B.n554 B.n553 163.367
R580 B.n553 B.n552 163.367
R581 B.n552 B.n29 163.367
R582 B.n548 B.n29 163.367
R583 B.n548 B.n547 163.367
R584 B.n547 B.n546 163.367
R585 B.n546 B.n31 163.367
R586 B.n542 B.n31 163.367
R587 B.n542 B.n541 163.367
R588 B.n541 B.n540 163.367
R589 B.n540 B.n33 163.367
R590 B.n536 B.n33 163.367
R591 B.n536 B.n535 163.367
R592 B.n535 B.n534 163.367
R593 B.n534 B.n35 163.367
R594 B.n530 B.n35 163.367
R595 B.n530 B.n529 163.367
R596 B.n529 B.n528 163.367
R597 B.n528 B.n37 163.367
R598 B.n524 B.n37 163.367
R599 B.n524 B.n523 163.367
R600 B.n523 B.n41 163.367
R601 B.n519 B.n41 163.367
R602 B.n519 B.n518 163.367
R603 B.n518 B.n517 163.367
R604 B.n517 B.n43 163.367
R605 B.n513 B.n43 163.367
R606 B.n513 B.n512 163.367
R607 B.n512 B.n511 163.367
R608 B.n511 B.n45 163.367
R609 B.n506 B.n45 163.367
R610 B.n506 B.n505 163.367
R611 B.n505 B.n504 163.367
R612 B.n504 B.n49 163.367
R613 B.n500 B.n49 163.367
R614 B.n500 B.n499 163.367
R615 B.n499 B.n498 163.367
R616 B.n498 B.n51 163.367
R617 B.n494 B.n51 163.367
R618 B.n494 B.n493 163.367
R619 B.n493 B.n492 163.367
R620 B.n492 B.n53 163.367
R621 B.n488 B.n53 163.367
R622 B.n488 B.n487 163.367
R623 B.n487 B.n486 163.367
R624 B.n486 B.n55 163.367
R625 B.n482 B.n55 163.367
R626 B.n482 B.n481 163.367
R627 B.n481 B.n480 163.367
R628 B.n480 B.n57 163.367
R629 B.n476 B.n57 163.367
R630 B.n476 B.n475 163.367
R631 B.n475 B.n474 163.367
R632 B.n474 B.n59 163.367
R633 B.n470 B.n59 163.367
R634 B.n470 B.n469 163.367
R635 B.n469 B.n468 163.367
R636 B.n468 B.n61 163.367
R637 B.n464 B.n61 163.367
R638 B.n464 B.n463 163.367
R639 B.n463 B.n462 163.367
R640 B.n462 B.n63 163.367
R641 B.n458 B.n63 163.367
R642 B.n458 B.n457 163.367
R643 B.n457 B.n456 163.367
R644 B.n456 B.n65 163.367
R645 B.n452 B.n65 163.367
R646 B.n452 B.n451 163.367
R647 B.n451 B.n450 163.367
R648 B.n450 B.n67 163.367
R649 B.n446 B.n67 163.367
R650 B.n446 B.n445 163.367
R651 B.n445 B.n444 163.367
R652 B.n444 B.n69 163.367
R653 B.n590 B.n15 163.367
R654 B.n594 B.n15 163.367
R655 B.n595 B.n594 163.367
R656 B.n596 B.n595 163.367
R657 B.n596 B.n13 163.367
R658 B.n600 B.n13 163.367
R659 B.n601 B.n600 163.367
R660 B.n602 B.n601 163.367
R661 B.n602 B.n11 163.367
R662 B.n606 B.n11 163.367
R663 B.n607 B.n606 163.367
R664 B.n608 B.n607 163.367
R665 B.n608 B.n9 163.367
R666 B.n612 B.n9 163.367
R667 B.n613 B.n612 163.367
R668 B.n614 B.n613 163.367
R669 B.n614 B.n7 163.367
R670 B.n618 B.n7 163.367
R671 B.n619 B.n618 163.367
R672 B.n620 B.n619 163.367
R673 B.n620 B.n5 163.367
R674 B.n624 B.n5 163.367
R675 B.n625 B.n624 163.367
R676 B.n626 B.n625 163.367
R677 B.n626 B.n3 163.367
R678 B.n630 B.n3 163.367
R679 B.n631 B.n630 163.367
R680 B.n164 B.n2 163.367
R681 B.n165 B.n164 163.367
R682 B.n166 B.n165 163.367
R683 B.n166 B.n161 163.367
R684 B.n170 B.n161 163.367
R685 B.n171 B.n170 163.367
R686 B.n172 B.n171 163.367
R687 B.n172 B.n159 163.367
R688 B.n176 B.n159 163.367
R689 B.n177 B.n176 163.367
R690 B.n178 B.n177 163.367
R691 B.n178 B.n157 163.367
R692 B.n182 B.n157 163.367
R693 B.n183 B.n182 163.367
R694 B.n184 B.n183 163.367
R695 B.n184 B.n155 163.367
R696 B.n188 B.n155 163.367
R697 B.n189 B.n188 163.367
R698 B.n190 B.n189 163.367
R699 B.n190 B.n153 163.367
R700 B.n194 B.n153 163.367
R701 B.n195 B.n194 163.367
R702 B.n196 B.n195 163.367
R703 B.n196 B.n151 163.367
R704 B.n200 B.n151 163.367
R705 B.n201 B.n200 163.367
R706 B.n202 B.n201 163.367
R707 B.n284 B.t10 141.036
R708 B.n46 B.t8 141.036
R709 B.n126 B.t1 141.019
R710 B.n38 B.t5 141.019
R711 B.n285 B.t11 107.677
R712 B.n47 B.t7 107.677
R713 B.n127 B.t2 107.662
R714 B.n39 B.t4 107.662
R715 B.n270 B.n127 59.5399
R716 B.n286 B.n285 59.5399
R717 B.n508 B.n47 59.5399
R718 B.n40 B.n39 59.5399
R719 B.n127 B.n126 33.3581
R720 B.n285 B.n284 33.3581
R721 B.n47 B.n46 33.3581
R722 B.n39 B.n38 33.3581
R723 B.n591 B.n16 33.2493
R724 B.n442 B.n441 33.2493
R725 B.n353 B.n98 33.2493
R726 B.n204 B.n203 33.2493
R727 B B.n633 18.0485
R728 B.n592 B.n591 10.6151
R729 B.n593 B.n592 10.6151
R730 B.n593 B.n14 10.6151
R731 B.n597 B.n14 10.6151
R732 B.n598 B.n597 10.6151
R733 B.n599 B.n598 10.6151
R734 B.n599 B.n12 10.6151
R735 B.n603 B.n12 10.6151
R736 B.n604 B.n603 10.6151
R737 B.n605 B.n604 10.6151
R738 B.n605 B.n10 10.6151
R739 B.n609 B.n10 10.6151
R740 B.n610 B.n609 10.6151
R741 B.n611 B.n610 10.6151
R742 B.n611 B.n8 10.6151
R743 B.n615 B.n8 10.6151
R744 B.n616 B.n615 10.6151
R745 B.n617 B.n616 10.6151
R746 B.n617 B.n6 10.6151
R747 B.n621 B.n6 10.6151
R748 B.n622 B.n621 10.6151
R749 B.n623 B.n622 10.6151
R750 B.n623 B.n4 10.6151
R751 B.n627 B.n4 10.6151
R752 B.n628 B.n627 10.6151
R753 B.n629 B.n628 10.6151
R754 B.n629 B.n0 10.6151
R755 B.n587 B.n16 10.6151
R756 B.n587 B.n586 10.6151
R757 B.n586 B.n585 10.6151
R758 B.n585 B.n18 10.6151
R759 B.n581 B.n18 10.6151
R760 B.n581 B.n580 10.6151
R761 B.n580 B.n579 10.6151
R762 B.n579 B.n20 10.6151
R763 B.n575 B.n20 10.6151
R764 B.n575 B.n574 10.6151
R765 B.n574 B.n573 10.6151
R766 B.n573 B.n22 10.6151
R767 B.n569 B.n22 10.6151
R768 B.n569 B.n568 10.6151
R769 B.n568 B.n567 10.6151
R770 B.n567 B.n24 10.6151
R771 B.n563 B.n24 10.6151
R772 B.n563 B.n562 10.6151
R773 B.n562 B.n561 10.6151
R774 B.n561 B.n26 10.6151
R775 B.n557 B.n26 10.6151
R776 B.n557 B.n556 10.6151
R777 B.n556 B.n555 10.6151
R778 B.n555 B.n28 10.6151
R779 B.n551 B.n28 10.6151
R780 B.n551 B.n550 10.6151
R781 B.n550 B.n549 10.6151
R782 B.n549 B.n30 10.6151
R783 B.n545 B.n30 10.6151
R784 B.n545 B.n544 10.6151
R785 B.n544 B.n543 10.6151
R786 B.n543 B.n32 10.6151
R787 B.n539 B.n32 10.6151
R788 B.n539 B.n538 10.6151
R789 B.n538 B.n537 10.6151
R790 B.n537 B.n34 10.6151
R791 B.n533 B.n34 10.6151
R792 B.n533 B.n532 10.6151
R793 B.n532 B.n531 10.6151
R794 B.n531 B.n36 10.6151
R795 B.n527 B.n36 10.6151
R796 B.n527 B.n526 10.6151
R797 B.n526 B.n525 10.6151
R798 B.n522 B.n521 10.6151
R799 B.n521 B.n520 10.6151
R800 B.n520 B.n42 10.6151
R801 B.n516 B.n42 10.6151
R802 B.n516 B.n515 10.6151
R803 B.n515 B.n514 10.6151
R804 B.n514 B.n44 10.6151
R805 B.n510 B.n44 10.6151
R806 B.n510 B.n509 10.6151
R807 B.n507 B.n48 10.6151
R808 B.n503 B.n48 10.6151
R809 B.n503 B.n502 10.6151
R810 B.n502 B.n501 10.6151
R811 B.n501 B.n50 10.6151
R812 B.n497 B.n50 10.6151
R813 B.n497 B.n496 10.6151
R814 B.n496 B.n495 10.6151
R815 B.n495 B.n52 10.6151
R816 B.n491 B.n52 10.6151
R817 B.n491 B.n490 10.6151
R818 B.n490 B.n489 10.6151
R819 B.n489 B.n54 10.6151
R820 B.n485 B.n54 10.6151
R821 B.n485 B.n484 10.6151
R822 B.n484 B.n483 10.6151
R823 B.n483 B.n56 10.6151
R824 B.n479 B.n56 10.6151
R825 B.n479 B.n478 10.6151
R826 B.n478 B.n477 10.6151
R827 B.n477 B.n58 10.6151
R828 B.n473 B.n58 10.6151
R829 B.n473 B.n472 10.6151
R830 B.n472 B.n471 10.6151
R831 B.n471 B.n60 10.6151
R832 B.n467 B.n60 10.6151
R833 B.n467 B.n466 10.6151
R834 B.n466 B.n465 10.6151
R835 B.n465 B.n62 10.6151
R836 B.n461 B.n62 10.6151
R837 B.n461 B.n460 10.6151
R838 B.n460 B.n459 10.6151
R839 B.n459 B.n64 10.6151
R840 B.n455 B.n64 10.6151
R841 B.n455 B.n454 10.6151
R842 B.n454 B.n453 10.6151
R843 B.n453 B.n66 10.6151
R844 B.n449 B.n66 10.6151
R845 B.n449 B.n448 10.6151
R846 B.n448 B.n447 10.6151
R847 B.n447 B.n68 10.6151
R848 B.n443 B.n68 10.6151
R849 B.n443 B.n442 10.6151
R850 B.n441 B.n70 10.6151
R851 B.n437 B.n70 10.6151
R852 B.n437 B.n436 10.6151
R853 B.n436 B.n435 10.6151
R854 B.n435 B.n72 10.6151
R855 B.n431 B.n72 10.6151
R856 B.n431 B.n430 10.6151
R857 B.n430 B.n429 10.6151
R858 B.n429 B.n74 10.6151
R859 B.n425 B.n74 10.6151
R860 B.n425 B.n424 10.6151
R861 B.n424 B.n423 10.6151
R862 B.n423 B.n76 10.6151
R863 B.n419 B.n76 10.6151
R864 B.n419 B.n418 10.6151
R865 B.n418 B.n417 10.6151
R866 B.n417 B.n78 10.6151
R867 B.n413 B.n78 10.6151
R868 B.n413 B.n412 10.6151
R869 B.n412 B.n411 10.6151
R870 B.n411 B.n80 10.6151
R871 B.n407 B.n80 10.6151
R872 B.n407 B.n406 10.6151
R873 B.n406 B.n405 10.6151
R874 B.n405 B.n82 10.6151
R875 B.n401 B.n82 10.6151
R876 B.n401 B.n400 10.6151
R877 B.n400 B.n399 10.6151
R878 B.n399 B.n84 10.6151
R879 B.n395 B.n84 10.6151
R880 B.n395 B.n394 10.6151
R881 B.n394 B.n393 10.6151
R882 B.n393 B.n86 10.6151
R883 B.n389 B.n86 10.6151
R884 B.n389 B.n388 10.6151
R885 B.n388 B.n387 10.6151
R886 B.n387 B.n88 10.6151
R887 B.n383 B.n88 10.6151
R888 B.n383 B.n382 10.6151
R889 B.n382 B.n381 10.6151
R890 B.n381 B.n90 10.6151
R891 B.n377 B.n90 10.6151
R892 B.n377 B.n376 10.6151
R893 B.n376 B.n375 10.6151
R894 B.n375 B.n92 10.6151
R895 B.n371 B.n92 10.6151
R896 B.n371 B.n370 10.6151
R897 B.n370 B.n369 10.6151
R898 B.n369 B.n94 10.6151
R899 B.n365 B.n94 10.6151
R900 B.n365 B.n364 10.6151
R901 B.n364 B.n363 10.6151
R902 B.n363 B.n96 10.6151
R903 B.n359 B.n96 10.6151
R904 B.n359 B.n358 10.6151
R905 B.n358 B.n357 10.6151
R906 B.n357 B.n98 10.6151
R907 B.n163 B.n1 10.6151
R908 B.n163 B.n162 10.6151
R909 B.n167 B.n162 10.6151
R910 B.n168 B.n167 10.6151
R911 B.n169 B.n168 10.6151
R912 B.n169 B.n160 10.6151
R913 B.n173 B.n160 10.6151
R914 B.n174 B.n173 10.6151
R915 B.n175 B.n174 10.6151
R916 B.n175 B.n158 10.6151
R917 B.n179 B.n158 10.6151
R918 B.n180 B.n179 10.6151
R919 B.n181 B.n180 10.6151
R920 B.n181 B.n156 10.6151
R921 B.n185 B.n156 10.6151
R922 B.n186 B.n185 10.6151
R923 B.n187 B.n186 10.6151
R924 B.n187 B.n154 10.6151
R925 B.n191 B.n154 10.6151
R926 B.n192 B.n191 10.6151
R927 B.n193 B.n192 10.6151
R928 B.n193 B.n152 10.6151
R929 B.n197 B.n152 10.6151
R930 B.n198 B.n197 10.6151
R931 B.n199 B.n198 10.6151
R932 B.n199 B.n150 10.6151
R933 B.n203 B.n150 10.6151
R934 B.n205 B.n204 10.6151
R935 B.n205 B.n148 10.6151
R936 B.n209 B.n148 10.6151
R937 B.n210 B.n209 10.6151
R938 B.n211 B.n210 10.6151
R939 B.n211 B.n146 10.6151
R940 B.n215 B.n146 10.6151
R941 B.n216 B.n215 10.6151
R942 B.n217 B.n216 10.6151
R943 B.n217 B.n144 10.6151
R944 B.n221 B.n144 10.6151
R945 B.n222 B.n221 10.6151
R946 B.n223 B.n222 10.6151
R947 B.n223 B.n142 10.6151
R948 B.n227 B.n142 10.6151
R949 B.n228 B.n227 10.6151
R950 B.n229 B.n228 10.6151
R951 B.n229 B.n140 10.6151
R952 B.n233 B.n140 10.6151
R953 B.n234 B.n233 10.6151
R954 B.n235 B.n234 10.6151
R955 B.n235 B.n138 10.6151
R956 B.n239 B.n138 10.6151
R957 B.n240 B.n239 10.6151
R958 B.n241 B.n240 10.6151
R959 B.n241 B.n136 10.6151
R960 B.n245 B.n136 10.6151
R961 B.n246 B.n245 10.6151
R962 B.n247 B.n246 10.6151
R963 B.n247 B.n134 10.6151
R964 B.n251 B.n134 10.6151
R965 B.n252 B.n251 10.6151
R966 B.n253 B.n252 10.6151
R967 B.n253 B.n132 10.6151
R968 B.n257 B.n132 10.6151
R969 B.n258 B.n257 10.6151
R970 B.n259 B.n258 10.6151
R971 B.n259 B.n130 10.6151
R972 B.n263 B.n130 10.6151
R973 B.n264 B.n263 10.6151
R974 B.n265 B.n264 10.6151
R975 B.n265 B.n128 10.6151
R976 B.n269 B.n128 10.6151
R977 B.n272 B.n271 10.6151
R978 B.n272 B.n124 10.6151
R979 B.n276 B.n124 10.6151
R980 B.n277 B.n276 10.6151
R981 B.n278 B.n277 10.6151
R982 B.n278 B.n122 10.6151
R983 B.n282 B.n122 10.6151
R984 B.n283 B.n282 10.6151
R985 B.n287 B.n283 10.6151
R986 B.n291 B.n120 10.6151
R987 B.n292 B.n291 10.6151
R988 B.n293 B.n292 10.6151
R989 B.n293 B.n118 10.6151
R990 B.n297 B.n118 10.6151
R991 B.n298 B.n297 10.6151
R992 B.n299 B.n298 10.6151
R993 B.n299 B.n116 10.6151
R994 B.n303 B.n116 10.6151
R995 B.n304 B.n303 10.6151
R996 B.n305 B.n304 10.6151
R997 B.n305 B.n114 10.6151
R998 B.n309 B.n114 10.6151
R999 B.n310 B.n309 10.6151
R1000 B.n311 B.n310 10.6151
R1001 B.n311 B.n112 10.6151
R1002 B.n315 B.n112 10.6151
R1003 B.n316 B.n315 10.6151
R1004 B.n317 B.n316 10.6151
R1005 B.n317 B.n110 10.6151
R1006 B.n321 B.n110 10.6151
R1007 B.n322 B.n321 10.6151
R1008 B.n323 B.n322 10.6151
R1009 B.n323 B.n108 10.6151
R1010 B.n327 B.n108 10.6151
R1011 B.n328 B.n327 10.6151
R1012 B.n329 B.n328 10.6151
R1013 B.n329 B.n106 10.6151
R1014 B.n333 B.n106 10.6151
R1015 B.n334 B.n333 10.6151
R1016 B.n335 B.n334 10.6151
R1017 B.n335 B.n104 10.6151
R1018 B.n339 B.n104 10.6151
R1019 B.n340 B.n339 10.6151
R1020 B.n341 B.n340 10.6151
R1021 B.n341 B.n102 10.6151
R1022 B.n345 B.n102 10.6151
R1023 B.n346 B.n345 10.6151
R1024 B.n347 B.n346 10.6151
R1025 B.n347 B.n100 10.6151
R1026 B.n351 B.n100 10.6151
R1027 B.n352 B.n351 10.6151
R1028 B.n353 B.n352 10.6151
R1029 B.n525 B.n40 9.36635
R1030 B.n508 B.n507 9.36635
R1031 B.n270 B.n269 9.36635
R1032 B.n286 B.n120 9.36635
R1033 B.n633 B.n0 8.11757
R1034 B.n633 B.n1 8.11757
R1035 B.n522 B.n40 1.24928
R1036 B.n509 B.n508 1.24928
R1037 B.n271 B.n270 1.24928
R1038 B.n287 B.n286 1.24928
R1039 VN.n3 VN.t2 259.094
R1040 VN.n13 VN.t3 259.094
R1041 VN.n2 VN.t5 224.702
R1042 VN.n8 VN.t4 224.702
R1043 VN.n12 VN.t0 224.702
R1044 VN.n18 VN.t1 224.702
R1045 VN.n9 VN.n8 174.933
R1046 VN.n19 VN.n18 174.933
R1047 VN.n17 VN.n10 161.3
R1048 VN.n16 VN.n15 161.3
R1049 VN.n14 VN.n11 161.3
R1050 VN.n7 VN.n0 161.3
R1051 VN.n6 VN.n5 161.3
R1052 VN.n4 VN.n1 161.3
R1053 VN.n6 VN.n1 54.0429
R1054 VN.n16 VN.n11 54.0429
R1055 VN VN.n19 44.9494
R1056 VN.n3 VN.n2 41.7088
R1057 VN.n13 VN.n12 41.7088
R1058 VN.n7 VN.n6 26.7783
R1059 VN.n17 VN.n16 26.7783
R1060 VN.n2 VN.n1 24.3439
R1061 VN.n12 VN.n11 24.3439
R1062 VN.n14 VN.n13 17.7134
R1063 VN.n4 VN.n3 17.7134
R1064 VN.n8 VN.n7 10.7116
R1065 VN.n18 VN.n17 10.7116
R1066 VN.n19 VN.n10 0.189894
R1067 VN.n15 VN.n10 0.189894
R1068 VN.n15 VN.n14 0.189894
R1069 VN.n5 VN.n4 0.189894
R1070 VN.n5 VN.n0 0.189894
R1071 VN.n9 VN.n0 0.189894
R1072 VN VN.n9 0.0516364
R1073 VDD2.n1 VDD2.t3 78.2007
R1074 VDD2.n2 VDD2.t4 77.1451
R1075 VDD2.n1 VDD2.n0 74.9512
R1076 VDD2 VDD2.n3 74.9484
R1077 VDD2.n2 VDD2.n1 39.7067
R1078 VDD2.n3 VDD2.t5 2.5086
R1079 VDD2.n3 VDD2.t2 2.5086
R1080 VDD2.n0 VDD2.t0 2.5086
R1081 VDD2.n0 VDD2.t1 2.5086
R1082 VDD2 VDD2.n2 1.17076
C0 w_n2346_n3560# VN 4.17557f
C1 VP VDD2 0.355675f
C2 VDD1 VDD2 0.96602f
C3 VTAIL w_n2346_n3560# 3.04505f
C4 VDD1 VP 6.37086f
C5 B w_n2346_n3560# 8.274281f
C6 VTAIL VN 6.00933f
C7 B VN 0.919674f
C8 VTAIL B 3.31734f
C9 w_n2346_n3560# VDD2 2.10777f
C10 w_n2346_n3560# VP 4.47551f
C11 VN VDD2 6.16799f
C12 VDD1 w_n2346_n3560# 2.0617f
C13 VN VP 5.93322f
C14 VDD1 VN 0.148764f
C15 VTAIL VDD2 8.602849f
C16 B VDD2 1.88169f
C17 VTAIL VP 6.02379f
C18 VDD1 VTAIL 8.56243f
C19 B VP 1.41435f
C20 VDD1 B 1.83646f
C21 VDD2 VSUBS 1.522718f
C22 VDD1 VSUBS 1.895537f
C23 VTAIL VSUBS 0.982548f
C24 VN VSUBS 4.84387f
C25 VP VSUBS 2.024248f
C26 B VSUBS 3.522257f
C27 w_n2346_n3560# VSUBS 0.10267p
C28 VDD2.t3 VSUBS 2.66215f
C29 VDD2.t0 VSUBS 0.255505f
C30 VDD2.t1 VSUBS 0.255505f
C31 VDD2.n0 VSUBS 2.03993f
C32 VDD2.n1 VSUBS 2.95287f
C33 VDD2.t4 VSUBS 2.65361f
C34 VDD2.n2 VSUBS 2.80121f
C35 VDD2.t5 VSUBS 0.255505f
C36 VDD2.t2 VSUBS 0.255505f
C37 VDD2.n3 VSUBS 2.0399f
C38 VN.n0 VSUBS 0.041406f
C39 VN.t4 VSUBS 2.03659f
C40 VN.n1 VSUBS 0.072927f
C41 VN.t2 VSUBS 2.15434f
C42 VN.t5 VSUBS 2.03659f
C43 VN.n2 VSUBS 0.829177f
C44 VN.n3 VSUBS 0.823724f
C45 VN.n4 VSUBS 0.259139f
C46 VN.n5 VSUBS 0.041406f
C47 VN.n6 VSUBS 0.045356f
C48 VN.n7 VSUBS 0.059246f
C49 VN.n8 VSUBS 0.814359f
C50 VN.n9 VSUBS 0.038788f
C51 VN.n10 VSUBS 0.041406f
C52 VN.t1 VSUBS 2.03659f
C53 VN.n11 VSUBS 0.072927f
C54 VN.t3 VSUBS 2.15434f
C55 VN.t0 VSUBS 2.03659f
C56 VN.n12 VSUBS 0.829177f
C57 VN.n13 VSUBS 0.823724f
C58 VN.n14 VSUBS 0.259139f
C59 VN.n15 VSUBS 0.041406f
C60 VN.n16 VSUBS 0.045356f
C61 VN.n17 VSUBS 0.059246f
C62 VN.n18 VSUBS 0.814359f
C63 VN.n19 VSUBS 1.91707f
C64 B.n0 VSUBS 0.005881f
C65 B.n1 VSUBS 0.005881f
C66 B.n2 VSUBS 0.008698f
C67 B.n3 VSUBS 0.006665f
C68 B.n4 VSUBS 0.006665f
C69 B.n5 VSUBS 0.006665f
C70 B.n6 VSUBS 0.006665f
C71 B.n7 VSUBS 0.006665f
C72 B.n8 VSUBS 0.006665f
C73 B.n9 VSUBS 0.006665f
C74 B.n10 VSUBS 0.006665f
C75 B.n11 VSUBS 0.006665f
C76 B.n12 VSUBS 0.006665f
C77 B.n13 VSUBS 0.006665f
C78 B.n14 VSUBS 0.006665f
C79 B.n15 VSUBS 0.006665f
C80 B.n16 VSUBS 0.015904f
C81 B.n17 VSUBS 0.006665f
C82 B.n18 VSUBS 0.006665f
C83 B.n19 VSUBS 0.006665f
C84 B.n20 VSUBS 0.006665f
C85 B.n21 VSUBS 0.006665f
C86 B.n22 VSUBS 0.006665f
C87 B.n23 VSUBS 0.006665f
C88 B.n24 VSUBS 0.006665f
C89 B.n25 VSUBS 0.006665f
C90 B.n26 VSUBS 0.006665f
C91 B.n27 VSUBS 0.006665f
C92 B.n28 VSUBS 0.006665f
C93 B.n29 VSUBS 0.006665f
C94 B.n30 VSUBS 0.006665f
C95 B.n31 VSUBS 0.006665f
C96 B.n32 VSUBS 0.006665f
C97 B.n33 VSUBS 0.006665f
C98 B.n34 VSUBS 0.006665f
C99 B.n35 VSUBS 0.006665f
C100 B.n36 VSUBS 0.006665f
C101 B.n37 VSUBS 0.006665f
C102 B.t4 VSUBS 0.405335f
C103 B.t5 VSUBS 0.418148f
C104 B.t3 VSUBS 0.741781f
C105 B.n38 VSUBS 0.179702f
C106 B.n39 VSUBS 0.063673f
C107 B.n40 VSUBS 0.015443f
C108 B.n41 VSUBS 0.006665f
C109 B.n42 VSUBS 0.006665f
C110 B.n43 VSUBS 0.006665f
C111 B.n44 VSUBS 0.006665f
C112 B.n45 VSUBS 0.006665f
C113 B.t7 VSUBS 0.405326f
C114 B.t8 VSUBS 0.41814f
C115 B.t6 VSUBS 0.741781f
C116 B.n46 VSUBS 0.179711f
C117 B.n47 VSUBS 0.063682f
C118 B.n48 VSUBS 0.006665f
C119 B.n49 VSUBS 0.006665f
C120 B.n50 VSUBS 0.006665f
C121 B.n51 VSUBS 0.006665f
C122 B.n52 VSUBS 0.006665f
C123 B.n53 VSUBS 0.006665f
C124 B.n54 VSUBS 0.006665f
C125 B.n55 VSUBS 0.006665f
C126 B.n56 VSUBS 0.006665f
C127 B.n57 VSUBS 0.006665f
C128 B.n58 VSUBS 0.006665f
C129 B.n59 VSUBS 0.006665f
C130 B.n60 VSUBS 0.006665f
C131 B.n61 VSUBS 0.006665f
C132 B.n62 VSUBS 0.006665f
C133 B.n63 VSUBS 0.006665f
C134 B.n64 VSUBS 0.006665f
C135 B.n65 VSUBS 0.006665f
C136 B.n66 VSUBS 0.006665f
C137 B.n67 VSUBS 0.006665f
C138 B.n68 VSUBS 0.006665f
C139 B.n69 VSUBS 0.015904f
C140 B.n70 VSUBS 0.006665f
C141 B.n71 VSUBS 0.006665f
C142 B.n72 VSUBS 0.006665f
C143 B.n73 VSUBS 0.006665f
C144 B.n74 VSUBS 0.006665f
C145 B.n75 VSUBS 0.006665f
C146 B.n76 VSUBS 0.006665f
C147 B.n77 VSUBS 0.006665f
C148 B.n78 VSUBS 0.006665f
C149 B.n79 VSUBS 0.006665f
C150 B.n80 VSUBS 0.006665f
C151 B.n81 VSUBS 0.006665f
C152 B.n82 VSUBS 0.006665f
C153 B.n83 VSUBS 0.006665f
C154 B.n84 VSUBS 0.006665f
C155 B.n85 VSUBS 0.006665f
C156 B.n86 VSUBS 0.006665f
C157 B.n87 VSUBS 0.006665f
C158 B.n88 VSUBS 0.006665f
C159 B.n89 VSUBS 0.006665f
C160 B.n90 VSUBS 0.006665f
C161 B.n91 VSUBS 0.006665f
C162 B.n92 VSUBS 0.006665f
C163 B.n93 VSUBS 0.006665f
C164 B.n94 VSUBS 0.006665f
C165 B.n95 VSUBS 0.006665f
C166 B.n96 VSUBS 0.006665f
C167 B.n97 VSUBS 0.006665f
C168 B.n98 VSUBS 0.016432f
C169 B.n99 VSUBS 0.006665f
C170 B.n100 VSUBS 0.006665f
C171 B.n101 VSUBS 0.006665f
C172 B.n102 VSUBS 0.006665f
C173 B.n103 VSUBS 0.006665f
C174 B.n104 VSUBS 0.006665f
C175 B.n105 VSUBS 0.006665f
C176 B.n106 VSUBS 0.006665f
C177 B.n107 VSUBS 0.006665f
C178 B.n108 VSUBS 0.006665f
C179 B.n109 VSUBS 0.006665f
C180 B.n110 VSUBS 0.006665f
C181 B.n111 VSUBS 0.006665f
C182 B.n112 VSUBS 0.006665f
C183 B.n113 VSUBS 0.006665f
C184 B.n114 VSUBS 0.006665f
C185 B.n115 VSUBS 0.006665f
C186 B.n116 VSUBS 0.006665f
C187 B.n117 VSUBS 0.006665f
C188 B.n118 VSUBS 0.006665f
C189 B.n119 VSUBS 0.006665f
C190 B.n120 VSUBS 0.006273f
C191 B.n121 VSUBS 0.006665f
C192 B.n122 VSUBS 0.006665f
C193 B.n123 VSUBS 0.006665f
C194 B.n124 VSUBS 0.006665f
C195 B.n125 VSUBS 0.006665f
C196 B.t2 VSUBS 0.405335f
C197 B.t1 VSUBS 0.418148f
C198 B.t0 VSUBS 0.741781f
C199 B.n126 VSUBS 0.179702f
C200 B.n127 VSUBS 0.063673f
C201 B.n128 VSUBS 0.006665f
C202 B.n129 VSUBS 0.006665f
C203 B.n130 VSUBS 0.006665f
C204 B.n131 VSUBS 0.006665f
C205 B.n132 VSUBS 0.006665f
C206 B.n133 VSUBS 0.006665f
C207 B.n134 VSUBS 0.006665f
C208 B.n135 VSUBS 0.006665f
C209 B.n136 VSUBS 0.006665f
C210 B.n137 VSUBS 0.006665f
C211 B.n138 VSUBS 0.006665f
C212 B.n139 VSUBS 0.006665f
C213 B.n140 VSUBS 0.006665f
C214 B.n141 VSUBS 0.006665f
C215 B.n142 VSUBS 0.006665f
C216 B.n143 VSUBS 0.006665f
C217 B.n144 VSUBS 0.006665f
C218 B.n145 VSUBS 0.006665f
C219 B.n146 VSUBS 0.006665f
C220 B.n147 VSUBS 0.006665f
C221 B.n148 VSUBS 0.006665f
C222 B.n149 VSUBS 0.015904f
C223 B.n150 VSUBS 0.006665f
C224 B.n151 VSUBS 0.006665f
C225 B.n152 VSUBS 0.006665f
C226 B.n153 VSUBS 0.006665f
C227 B.n154 VSUBS 0.006665f
C228 B.n155 VSUBS 0.006665f
C229 B.n156 VSUBS 0.006665f
C230 B.n157 VSUBS 0.006665f
C231 B.n158 VSUBS 0.006665f
C232 B.n159 VSUBS 0.006665f
C233 B.n160 VSUBS 0.006665f
C234 B.n161 VSUBS 0.006665f
C235 B.n162 VSUBS 0.006665f
C236 B.n163 VSUBS 0.006665f
C237 B.n164 VSUBS 0.006665f
C238 B.n165 VSUBS 0.006665f
C239 B.n166 VSUBS 0.006665f
C240 B.n167 VSUBS 0.006665f
C241 B.n168 VSUBS 0.006665f
C242 B.n169 VSUBS 0.006665f
C243 B.n170 VSUBS 0.006665f
C244 B.n171 VSUBS 0.006665f
C245 B.n172 VSUBS 0.006665f
C246 B.n173 VSUBS 0.006665f
C247 B.n174 VSUBS 0.006665f
C248 B.n175 VSUBS 0.006665f
C249 B.n176 VSUBS 0.006665f
C250 B.n177 VSUBS 0.006665f
C251 B.n178 VSUBS 0.006665f
C252 B.n179 VSUBS 0.006665f
C253 B.n180 VSUBS 0.006665f
C254 B.n181 VSUBS 0.006665f
C255 B.n182 VSUBS 0.006665f
C256 B.n183 VSUBS 0.006665f
C257 B.n184 VSUBS 0.006665f
C258 B.n185 VSUBS 0.006665f
C259 B.n186 VSUBS 0.006665f
C260 B.n187 VSUBS 0.006665f
C261 B.n188 VSUBS 0.006665f
C262 B.n189 VSUBS 0.006665f
C263 B.n190 VSUBS 0.006665f
C264 B.n191 VSUBS 0.006665f
C265 B.n192 VSUBS 0.006665f
C266 B.n193 VSUBS 0.006665f
C267 B.n194 VSUBS 0.006665f
C268 B.n195 VSUBS 0.006665f
C269 B.n196 VSUBS 0.006665f
C270 B.n197 VSUBS 0.006665f
C271 B.n198 VSUBS 0.006665f
C272 B.n199 VSUBS 0.006665f
C273 B.n200 VSUBS 0.006665f
C274 B.n201 VSUBS 0.006665f
C275 B.n202 VSUBS 0.015659f
C276 B.n203 VSUBS 0.015659f
C277 B.n204 VSUBS 0.015904f
C278 B.n205 VSUBS 0.006665f
C279 B.n206 VSUBS 0.006665f
C280 B.n207 VSUBS 0.006665f
C281 B.n208 VSUBS 0.006665f
C282 B.n209 VSUBS 0.006665f
C283 B.n210 VSUBS 0.006665f
C284 B.n211 VSUBS 0.006665f
C285 B.n212 VSUBS 0.006665f
C286 B.n213 VSUBS 0.006665f
C287 B.n214 VSUBS 0.006665f
C288 B.n215 VSUBS 0.006665f
C289 B.n216 VSUBS 0.006665f
C290 B.n217 VSUBS 0.006665f
C291 B.n218 VSUBS 0.006665f
C292 B.n219 VSUBS 0.006665f
C293 B.n220 VSUBS 0.006665f
C294 B.n221 VSUBS 0.006665f
C295 B.n222 VSUBS 0.006665f
C296 B.n223 VSUBS 0.006665f
C297 B.n224 VSUBS 0.006665f
C298 B.n225 VSUBS 0.006665f
C299 B.n226 VSUBS 0.006665f
C300 B.n227 VSUBS 0.006665f
C301 B.n228 VSUBS 0.006665f
C302 B.n229 VSUBS 0.006665f
C303 B.n230 VSUBS 0.006665f
C304 B.n231 VSUBS 0.006665f
C305 B.n232 VSUBS 0.006665f
C306 B.n233 VSUBS 0.006665f
C307 B.n234 VSUBS 0.006665f
C308 B.n235 VSUBS 0.006665f
C309 B.n236 VSUBS 0.006665f
C310 B.n237 VSUBS 0.006665f
C311 B.n238 VSUBS 0.006665f
C312 B.n239 VSUBS 0.006665f
C313 B.n240 VSUBS 0.006665f
C314 B.n241 VSUBS 0.006665f
C315 B.n242 VSUBS 0.006665f
C316 B.n243 VSUBS 0.006665f
C317 B.n244 VSUBS 0.006665f
C318 B.n245 VSUBS 0.006665f
C319 B.n246 VSUBS 0.006665f
C320 B.n247 VSUBS 0.006665f
C321 B.n248 VSUBS 0.006665f
C322 B.n249 VSUBS 0.006665f
C323 B.n250 VSUBS 0.006665f
C324 B.n251 VSUBS 0.006665f
C325 B.n252 VSUBS 0.006665f
C326 B.n253 VSUBS 0.006665f
C327 B.n254 VSUBS 0.006665f
C328 B.n255 VSUBS 0.006665f
C329 B.n256 VSUBS 0.006665f
C330 B.n257 VSUBS 0.006665f
C331 B.n258 VSUBS 0.006665f
C332 B.n259 VSUBS 0.006665f
C333 B.n260 VSUBS 0.006665f
C334 B.n261 VSUBS 0.006665f
C335 B.n262 VSUBS 0.006665f
C336 B.n263 VSUBS 0.006665f
C337 B.n264 VSUBS 0.006665f
C338 B.n265 VSUBS 0.006665f
C339 B.n266 VSUBS 0.006665f
C340 B.n267 VSUBS 0.006665f
C341 B.n268 VSUBS 0.006665f
C342 B.n269 VSUBS 0.006273f
C343 B.n270 VSUBS 0.015443f
C344 B.n271 VSUBS 0.003725f
C345 B.n272 VSUBS 0.006665f
C346 B.n273 VSUBS 0.006665f
C347 B.n274 VSUBS 0.006665f
C348 B.n275 VSUBS 0.006665f
C349 B.n276 VSUBS 0.006665f
C350 B.n277 VSUBS 0.006665f
C351 B.n278 VSUBS 0.006665f
C352 B.n279 VSUBS 0.006665f
C353 B.n280 VSUBS 0.006665f
C354 B.n281 VSUBS 0.006665f
C355 B.n282 VSUBS 0.006665f
C356 B.n283 VSUBS 0.006665f
C357 B.t11 VSUBS 0.405326f
C358 B.t10 VSUBS 0.41814f
C359 B.t9 VSUBS 0.741781f
C360 B.n284 VSUBS 0.179711f
C361 B.n285 VSUBS 0.063682f
C362 B.n286 VSUBS 0.015443f
C363 B.n287 VSUBS 0.003725f
C364 B.n288 VSUBS 0.006665f
C365 B.n289 VSUBS 0.006665f
C366 B.n290 VSUBS 0.006665f
C367 B.n291 VSUBS 0.006665f
C368 B.n292 VSUBS 0.006665f
C369 B.n293 VSUBS 0.006665f
C370 B.n294 VSUBS 0.006665f
C371 B.n295 VSUBS 0.006665f
C372 B.n296 VSUBS 0.006665f
C373 B.n297 VSUBS 0.006665f
C374 B.n298 VSUBS 0.006665f
C375 B.n299 VSUBS 0.006665f
C376 B.n300 VSUBS 0.006665f
C377 B.n301 VSUBS 0.006665f
C378 B.n302 VSUBS 0.006665f
C379 B.n303 VSUBS 0.006665f
C380 B.n304 VSUBS 0.006665f
C381 B.n305 VSUBS 0.006665f
C382 B.n306 VSUBS 0.006665f
C383 B.n307 VSUBS 0.006665f
C384 B.n308 VSUBS 0.006665f
C385 B.n309 VSUBS 0.006665f
C386 B.n310 VSUBS 0.006665f
C387 B.n311 VSUBS 0.006665f
C388 B.n312 VSUBS 0.006665f
C389 B.n313 VSUBS 0.006665f
C390 B.n314 VSUBS 0.006665f
C391 B.n315 VSUBS 0.006665f
C392 B.n316 VSUBS 0.006665f
C393 B.n317 VSUBS 0.006665f
C394 B.n318 VSUBS 0.006665f
C395 B.n319 VSUBS 0.006665f
C396 B.n320 VSUBS 0.006665f
C397 B.n321 VSUBS 0.006665f
C398 B.n322 VSUBS 0.006665f
C399 B.n323 VSUBS 0.006665f
C400 B.n324 VSUBS 0.006665f
C401 B.n325 VSUBS 0.006665f
C402 B.n326 VSUBS 0.006665f
C403 B.n327 VSUBS 0.006665f
C404 B.n328 VSUBS 0.006665f
C405 B.n329 VSUBS 0.006665f
C406 B.n330 VSUBS 0.006665f
C407 B.n331 VSUBS 0.006665f
C408 B.n332 VSUBS 0.006665f
C409 B.n333 VSUBS 0.006665f
C410 B.n334 VSUBS 0.006665f
C411 B.n335 VSUBS 0.006665f
C412 B.n336 VSUBS 0.006665f
C413 B.n337 VSUBS 0.006665f
C414 B.n338 VSUBS 0.006665f
C415 B.n339 VSUBS 0.006665f
C416 B.n340 VSUBS 0.006665f
C417 B.n341 VSUBS 0.006665f
C418 B.n342 VSUBS 0.006665f
C419 B.n343 VSUBS 0.006665f
C420 B.n344 VSUBS 0.006665f
C421 B.n345 VSUBS 0.006665f
C422 B.n346 VSUBS 0.006665f
C423 B.n347 VSUBS 0.006665f
C424 B.n348 VSUBS 0.006665f
C425 B.n349 VSUBS 0.006665f
C426 B.n350 VSUBS 0.006665f
C427 B.n351 VSUBS 0.006665f
C428 B.n352 VSUBS 0.006665f
C429 B.n353 VSUBS 0.01513f
C430 B.n354 VSUBS 0.015904f
C431 B.n355 VSUBS 0.015659f
C432 B.n356 VSUBS 0.006665f
C433 B.n357 VSUBS 0.006665f
C434 B.n358 VSUBS 0.006665f
C435 B.n359 VSUBS 0.006665f
C436 B.n360 VSUBS 0.006665f
C437 B.n361 VSUBS 0.006665f
C438 B.n362 VSUBS 0.006665f
C439 B.n363 VSUBS 0.006665f
C440 B.n364 VSUBS 0.006665f
C441 B.n365 VSUBS 0.006665f
C442 B.n366 VSUBS 0.006665f
C443 B.n367 VSUBS 0.006665f
C444 B.n368 VSUBS 0.006665f
C445 B.n369 VSUBS 0.006665f
C446 B.n370 VSUBS 0.006665f
C447 B.n371 VSUBS 0.006665f
C448 B.n372 VSUBS 0.006665f
C449 B.n373 VSUBS 0.006665f
C450 B.n374 VSUBS 0.006665f
C451 B.n375 VSUBS 0.006665f
C452 B.n376 VSUBS 0.006665f
C453 B.n377 VSUBS 0.006665f
C454 B.n378 VSUBS 0.006665f
C455 B.n379 VSUBS 0.006665f
C456 B.n380 VSUBS 0.006665f
C457 B.n381 VSUBS 0.006665f
C458 B.n382 VSUBS 0.006665f
C459 B.n383 VSUBS 0.006665f
C460 B.n384 VSUBS 0.006665f
C461 B.n385 VSUBS 0.006665f
C462 B.n386 VSUBS 0.006665f
C463 B.n387 VSUBS 0.006665f
C464 B.n388 VSUBS 0.006665f
C465 B.n389 VSUBS 0.006665f
C466 B.n390 VSUBS 0.006665f
C467 B.n391 VSUBS 0.006665f
C468 B.n392 VSUBS 0.006665f
C469 B.n393 VSUBS 0.006665f
C470 B.n394 VSUBS 0.006665f
C471 B.n395 VSUBS 0.006665f
C472 B.n396 VSUBS 0.006665f
C473 B.n397 VSUBS 0.006665f
C474 B.n398 VSUBS 0.006665f
C475 B.n399 VSUBS 0.006665f
C476 B.n400 VSUBS 0.006665f
C477 B.n401 VSUBS 0.006665f
C478 B.n402 VSUBS 0.006665f
C479 B.n403 VSUBS 0.006665f
C480 B.n404 VSUBS 0.006665f
C481 B.n405 VSUBS 0.006665f
C482 B.n406 VSUBS 0.006665f
C483 B.n407 VSUBS 0.006665f
C484 B.n408 VSUBS 0.006665f
C485 B.n409 VSUBS 0.006665f
C486 B.n410 VSUBS 0.006665f
C487 B.n411 VSUBS 0.006665f
C488 B.n412 VSUBS 0.006665f
C489 B.n413 VSUBS 0.006665f
C490 B.n414 VSUBS 0.006665f
C491 B.n415 VSUBS 0.006665f
C492 B.n416 VSUBS 0.006665f
C493 B.n417 VSUBS 0.006665f
C494 B.n418 VSUBS 0.006665f
C495 B.n419 VSUBS 0.006665f
C496 B.n420 VSUBS 0.006665f
C497 B.n421 VSUBS 0.006665f
C498 B.n422 VSUBS 0.006665f
C499 B.n423 VSUBS 0.006665f
C500 B.n424 VSUBS 0.006665f
C501 B.n425 VSUBS 0.006665f
C502 B.n426 VSUBS 0.006665f
C503 B.n427 VSUBS 0.006665f
C504 B.n428 VSUBS 0.006665f
C505 B.n429 VSUBS 0.006665f
C506 B.n430 VSUBS 0.006665f
C507 B.n431 VSUBS 0.006665f
C508 B.n432 VSUBS 0.006665f
C509 B.n433 VSUBS 0.006665f
C510 B.n434 VSUBS 0.006665f
C511 B.n435 VSUBS 0.006665f
C512 B.n436 VSUBS 0.006665f
C513 B.n437 VSUBS 0.006665f
C514 B.n438 VSUBS 0.006665f
C515 B.n439 VSUBS 0.006665f
C516 B.n440 VSUBS 0.015659f
C517 B.n441 VSUBS 0.015659f
C518 B.n442 VSUBS 0.015904f
C519 B.n443 VSUBS 0.006665f
C520 B.n444 VSUBS 0.006665f
C521 B.n445 VSUBS 0.006665f
C522 B.n446 VSUBS 0.006665f
C523 B.n447 VSUBS 0.006665f
C524 B.n448 VSUBS 0.006665f
C525 B.n449 VSUBS 0.006665f
C526 B.n450 VSUBS 0.006665f
C527 B.n451 VSUBS 0.006665f
C528 B.n452 VSUBS 0.006665f
C529 B.n453 VSUBS 0.006665f
C530 B.n454 VSUBS 0.006665f
C531 B.n455 VSUBS 0.006665f
C532 B.n456 VSUBS 0.006665f
C533 B.n457 VSUBS 0.006665f
C534 B.n458 VSUBS 0.006665f
C535 B.n459 VSUBS 0.006665f
C536 B.n460 VSUBS 0.006665f
C537 B.n461 VSUBS 0.006665f
C538 B.n462 VSUBS 0.006665f
C539 B.n463 VSUBS 0.006665f
C540 B.n464 VSUBS 0.006665f
C541 B.n465 VSUBS 0.006665f
C542 B.n466 VSUBS 0.006665f
C543 B.n467 VSUBS 0.006665f
C544 B.n468 VSUBS 0.006665f
C545 B.n469 VSUBS 0.006665f
C546 B.n470 VSUBS 0.006665f
C547 B.n471 VSUBS 0.006665f
C548 B.n472 VSUBS 0.006665f
C549 B.n473 VSUBS 0.006665f
C550 B.n474 VSUBS 0.006665f
C551 B.n475 VSUBS 0.006665f
C552 B.n476 VSUBS 0.006665f
C553 B.n477 VSUBS 0.006665f
C554 B.n478 VSUBS 0.006665f
C555 B.n479 VSUBS 0.006665f
C556 B.n480 VSUBS 0.006665f
C557 B.n481 VSUBS 0.006665f
C558 B.n482 VSUBS 0.006665f
C559 B.n483 VSUBS 0.006665f
C560 B.n484 VSUBS 0.006665f
C561 B.n485 VSUBS 0.006665f
C562 B.n486 VSUBS 0.006665f
C563 B.n487 VSUBS 0.006665f
C564 B.n488 VSUBS 0.006665f
C565 B.n489 VSUBS 0.006665f
C566 B.n490 VSUBS 0.006665f
C567 B.n491 VSUBS 0.006665f
C568 B.n492 VSUBS 0.006665f
C569 B.n493 VSUBS 0.006665f
C570 B.n494 VSUBS 0.006665f
C571 B.n495 VSUBS 0.006665f
C572 B.n496 VSUBS 0.006665f
C573 B.n497 VSUBS 0.006665f
C574 B.n498 VSUBS 0.006665f
C575 B.n499 VSUBS 0.006665f
C576 B.n500 VSUBS 0.006665f
C577 B.n501 VSUBS 0.006665f
C578 B.n502 VSUBS 0.006665f
C579 B.n503 VSUBS 0.006665f
C580 B.n504 VSUBS 0.006665f
C581 B.n505 VSUBS 0.006665f
C582 B.n506 VSUBS 0.006665f
C583 B.n507 VSUBS 0.006273f
C584 B.n508 VSUBS 0.015443f
C585 B.n509 VSUBS 0.003725f
C586 B.n510 VSUBS 0.006665f
C587 B.n511 VSUBS 0.006665f
C588 B.n512 VSUBS 0.006665f
C589 B.n513 VSUBS 0.006665f
C590 B.n514 VSUBS 0.006665f
C591 B.n515 VSUBS 0.006665f
C592 B.n516 VSUBS 0.006665f
C593 B.n517 VSUBS 0.006665f
C594 B.n518 VSUBS 0.006665f
C595 B.n519 VSUBS 0.006665f
C596 B.n520 VSUBS 0.006665f
C597 B.n521 VSUBS 0.006665f
C598 B.n522 VSUBS 0.003725f
C599 B.n523 VSUBS 0.006665f
C600 B.n524 VSUBS 0.006665f
C601 B.n525 VSUBS 0.006273f
C602 B.n526 VSUBS 0.006665f
C603 B.n527 VSUBS 0.006665f
C604 B.n528 VSUBS 0.006665f
C605 B.n529 VSUBS 0.006665f
C606 B.n530 VSUBS 0.006665f
C607 B.n531 VSUBS 0.006665f
C608 B.n532 VSUBS 0.006665f
C609 B.n533 VSUBS 0.006665f
C610 B.n534 VSUBS 0.006665f
C611 B.n535 VSUBS 0.006665f
C612 B.n536 VSUBS 0.006665f
C613 B.n537 VSUBS 0.006665f
C614 B.n538 VSUBS 0.006665f
C615 B.n539 VSUBS 0.006665f
C616 B.n540 VSUBS 0.006665f
C617 B.n541 VSUBS 0.006665f
C618 B.n542 VSUBS 0.006665f
C619 B.n543 VSUBS 0.006665f
C620 B.n544 VSUBS 0.006665f
C621 B.n545 VSUBS 0.006665f
C622 B.n546 VSUBS 0.006665f
C623 B.n547 VSUBS 0.006665f
C624 B.n548 VSUBS 0.006665f
C625 B.n549 VSUBS 0.006665f
C626 B.n550 VSUBS 0.006665f
C627 B.n551 VSUBS 0.006665f
C628 B.n552 VSUBS 0.006665f
C629 B.n553 VSUBS 0.006665f
C630 B.n554 VSUBS 0.006665f
C631 B.n555 VSUBS 0.006665f
C632 B.n556 VSUBS 0.006665f
C633 B.n557 VSUBS 0.006665f
C634 B.n558 VSUBS 0.006665f
C635 B.n559 VSUBS 0.006665f
C636 B.n560 VSUBS 0.006665f
C637 B.n561 VSUBS 0.006665f
C638 B.n562 VSUBS 0.006665f
C639 B.n563 VSUBS 0.006665f
C640 B.n564 VSUBS 0.006665f
C641 B.n565 VSUBS 0.006665f
C642 B.n566 VSUBS 0.006665f
C643 B.n567 VSUBS 0.006665f
C644 B.n568 VSUBS 0.006665f
C645 B.n569 VSUBS 0.006665f
C646 B.n570 VSUBS 0.006665f
C647 B.n571 VSUBS 0.006665f
C648 B.n572 VSUBS 0.006665f
C649 B.n573 VSUBS 0.006665f
C650 B.n574 VSUBS 0.006665f
C651 B.n575 VSUBS 0.006665f
C652 B.n576 VSUBS 0.006665f
C653 B.n577 VSUBS 0.006665f
C654 B.n578 VSUBS 0.006665f
C655 B.n579 VSUBS 0.006665f
C656 B.n580 VSUBS 0.006665f
C657 B.n581 VSUBS 0.006665f
C658 B.n582 VSUBS 0.006665f
C659 B.n583 VSUBS 0.006665f
C660 B.n584 VSUBS 0.006665f
C661 B.n585 VSUBS 0.006665f
C662 B.n586 VSUBS 0.006665f
C663 B.n587 VSUBS 0.006665f
C664 B.n588 VSUBS 0.006665f
C665 B.n589 VSUBS 0.015904f
C666 B.n590 VSUBS 0.015659f
C667 B.n591 VSUBS 0.015659f
C668 B.n592 VSUBS 0.006665f
C669 B.n593 VSUBS 0.006665f
C670 B.n594 VSUBS 0.006665f
C671 B.n595 VSUBS 0.006665f
C672 B.n596 VSUBS 0.006665f
C673 B.n597 VSUBS 0.006665f
C674 B.n598 VSUBS 0.006665f
C675 B.n599 VSUBS 0.006665f
C676 B.n600 VSUBS 0.006665f
C677 B.n601 VSUBS 0.006665f
C678 B.n602 VSUBS 0.006665f
C679 B.n603 VSUBS 0.006665f
C680 B.n604 VSUBS 0.006665f
C681 B.n605 VSUBS 0.006665f
C682 B.n606 VSUBS 0.006665f
C683 B.n607 VSUBS 0.006665f
C684 B.n608 VSUBS 0.006665f
C685 B.n609 VSUBS 0.006665f
C686 B.n610 VSUBS 0.006665f
C687 B.n611 VSUBS 0.006665f
C688 B.n612 VSUBS 0.006665f
C689 B.n613 VSUBS 0.006665f
C690 B.n614 VSUBS 0.006665f
C691 B.n615 VSUBS 0.006665f
C692 B.n616 VSUBS 0.006665f
C693 B.n617 VSUBS 0.006665f
C694 B.n618 VSUBS 0.006665f
C695 B.n619 VSUBS 0.006665f
C696 B.n620 VSUBS 0.006665f
C697 B.n621 VSUBS 0.006665f
C698 B.n622 VSUBS 0.006665f
C699 B.n623 VSUBS 0.006665f
C700 B.n624 VSUBS 0.006665f
C701 B.n625 VSUBS 0.006665f
C702 B.n626 VSUBS 0.006665f
C703 B.n627 VSUBS 0.006665f
C704 B.n628 VSUBS 0.006665f
C705 B.n629 VSUBS 0.006665f
C706 B.n630 VSUBS 0.006665f
C707 B.n631 VSUBS 0.008698f
C708 B.n632 VSUBS 0.009266f
C709 B.n633 VSUBS 0.018425f
C710 VDD1.t1 VSUBS 2.6801f
C711 VDD1.t4 VSUBS 2.67905f
C712 VDD1.t0 VSUBS 0.257127f
C713 VDD1.t5 VSUBS 0.257127f
C714 VDD1.n0 VSUBS 2.05288f
C715 VDD1.n1 VSUBS 3.06605f
C716 VDD1.t2 VSUBS 0.257127f
C717 VDD1.t3 VSUBS 0.257127f
C718 VDD1.n2 VSUBS 2.05028f
C719 VDD1.n3 VSUBS 2.78675f
C720 VTAIL.t3 VSUBS 0.287734f
C721 VTAIL.t0 VSUBS 0.287734f
C722 VTAIL.n0 VSUBS 2.14767f
C723 VTAIL.n1 VSUBS 0.77194f
C724 VTAIL.t6 VSUBS 2.8227f
C725 VTAIL.n2 VSUBS 0.977051f
C726 VTAIL.t10 VSUBS 0.287734f
C727 VTAIL.t7 VSUBS 0.287734f
C728 VTAIL.n3 VSUBS 2.14767f
C729 VTAIL.n4 VSUBS 2.41923f
C730 VTAIL.t2 VSUBS 0.287734f
C731 VTAIL.t5 VSUBS 0.287734f
C732 VTAIL.n5 VSUBS 2.14769f
C733 VTAIL.n6 VSUBS 2.41921f
C734 VTAIL.t4 VSUBS 2.82272f
C735 VTAIL.n7 VSUBS 0.977026f
C736 VTAIL.t11 VSUBS 0.287734f
C737 VTAIL.t9 VSUBS 0.287734f
C738 VTAIL.n8 VSUBS 2.14769f
C739 VTAIL.n9 VSUBS 0.867328f
C740 VTAIL.t8 VSUBS 2.8227f
C741 VTAIL.n10 VSUBS 2.3947f
C742 VTAIL.t1 VSUBS 2.8227f
C743 VTAIL.n11 VSUBS 2.35588f
C744 VP.n0 VSUBS 0.042445f
C745 VP.t0 VSUBS 2.0877f
C746 VP.n1 VSUBS 0.074757f
C747 VP.n2 VSUBS 0.042445f
C748 VP.t5 VSUBS 2.0877f
C749 VP.n3 VSUBS 0.060733f
C750 VP.n4 VSUBS 0.042445f
C751 VP.t2 VSUBS 2.0877f
C752 VP.n5 VSUBS 0.074757f
C753 VP.t4 VSUBS 2.20841f
C754 VP.t3 VSUBS 2.0877f
C755 VP.n6 VSUBS 0.849986f
C756 VP.n7 VSUBS 0.844397f
C757 VP.n8 VSUBS 0.265643f
C758 VP.n9 VSUBS 0.042445f
C759 VP.n10 VSUBS 0.046494f
C760 VP.n11 VSUBS 0.060733f
C761 VP.n12 VSUBS 0.834797f
C762 VP.n13 VSUBS 1.93742f
C763 VP.t1 VSUBS 2.0877f
C764 VP.n14 VSUBS 0.834797f
C765 VP.n15 VSUBS 1.97155f
C766 VP.n16 VSUBS 0.042445f
C767 VP.n17 VSUBS 0.042445f
C768 VP.n18 VSUBS 0.046494f
C769 VP.n19 VSUBS 0.074757f
C770 VP.n20 VSUBS 0.793776f
C771 VP.n21 VSUBS 0.042445f
C772 VP.n22 VSUBS 0.042445f
C773 VP.n23 VSUBS 0.042445f
C774 VP.n24 VSUBS 0.046494f
C775 VP.n25 VSUBS 0.060733f
C776 VP.n26 VSUBS 0.834797f
C777 VP.n27 VSUBS 0.039762f
.ends

