* NGSPICE file created from diff_pair_sample_0766.ext - technology: sky130A

.subckt diff_pair_sample_0766 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X1 VTAIL.t9 VP.t0 VDD1.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X2 VDD1.t8 VP.t1 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=2.12
X3 VDD2.t8 VN.t1 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X4 VDD1.t7 VP.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=2.12
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=2.12
X6 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X7 VDD1.t5 VP.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X8 VTAIL.t15 VN.t2 VDD2.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X9 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=2.12
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=2.12
X11 VTAIL.t10 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X12 VTAIL.t4 VP.t5 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X13 VTAIL.t3 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X14 VDD1.t2 VP.t7 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=2.12
X15 VDD2.t5 VN.t4 VTAIL.t18 B.t1 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=2.12
X16 VDD2.t4 VN.t5 VTAIL.t16 B.t7 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=2.12
X17 VDD2.t3 VN.t6 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.585 ps=3.78 w=1.5 l=2.12
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0 ps=0 w=1.5 l=2.12
X19 VDD2.t2 VN.t7 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=2.12
X20 VDD1.t1 VP.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.585 pd=3.78 as=0.2475 ps=1.83 w=1.5 l=2.12
X21 VDD1.t0 VP.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X22 VTAIL.t13 VN.t8 VDD2.t1 B.t9 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
X23 VTAIL.t14 VN.t9 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2475 pd=1.83 as=0.2475 ps=1.83 w=1.5 l=2.12
R0 VN.n63 VN.n33 161.3
R1 VN.n62 VN.n61 161.3
R2 VN.n60 VN.n34 161.3
R3 VN.n59 VN.n58 161.3
R4 VN.n57 VN.n35 161.3
R5 VN.n55 VN.n54 161.3
R6 VN.n53 VN.n36 161.3
R7 VN.n52 VN.n51 161.3
R8 VN.n50 VN.n37 161.3
R9 VN.n49 VN.n48 161.3
R10 VN.n47 VN.n38 161.3
R11 VN.n46 VN.n45 161.3
R12 VN.n44 VN.n39 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n30 VN.n0 161.3
R15 VN.n29 VN.n28 161.3
R16 VN.n27 VN.n1 161.3
R17 VN.n26 VN.n25 161.3
R18 VN.n24 VN.n2 161.3
R19 VN.n22 VN.n21 161.3
R20 VN.n20 VN.n3 161.3
R21 VN.n19 VN.n18 161.3
R22 VN.n17 VN.n4 161.3
R23 VN.n16 VN.n15 161.3
R24 VN.n14 VN.n5 161.3
R25 VN.n13 VN.n12 161.3
R26 VN.n11 VN.n6 161.3
R27 VN.n10 VN.n9 161.3
R28 VN.n32 VN.n31 91.2348
R29 VN.n65 VN.n64 91.2348
R30 VN.n12 VN.n11 56.5617
R31 VN.n18 VN.n3 56.5617
R32 VN.n29 VN.n1 56.5617
R33 VN.n45 VN.n44 56.5617
R34 VN.n51 VN.n36 56.5617
R35 VN.n62 VN.n34 56.5617
R36 VN.n8 VN.t7 51.2161
R37 VN.n41 VN.t6 51.2161
R38 VN.n8 VN.n7 48.5947
R39 VN.n41 VN.n40 48.5947
R40 VN VN.n65 42.8808
R41 VN.n11 VN.n10 24.5923
R42 VN.n12 VN.n5 24.5923
R43 VN.n16 VN.n5 24.5923
R44 VN.n17 VN.n16 24.5923
R45 VN.n18 VN.n17 24.5923
R46 VN.n22 VN.n3 24.5923
R47 VN.n25 VN.n24 24.5923
R48 VN.n25 VN.n1 24.5923
R49 VN.n30 VN.n29 24.5923
R50 VN.n44 VN.n43 24.5923
R51 VN.n51 VN.n50 24.5923
R52 VN.n50 VN.n49 24.5923
R53 VN.n49 VN.n38 24.5923
R54 VN.n45 VN.n38 24.5923
R55 VN.n58 VN.n34 24.5923
R56 VN.n58 VN.n57 24.5923
R57 VN.n55 VN.n36 24.5923
R58 VN.n63 VN.n62 24.5923
R59 VN.n10 VN.n7 22.1332
R60 VN.n23 VN.n22 22.1332
R61 VN.n43 VN.n40 22.1332
R62 VN.n56 VN.n55 22.1332
R63 VN.n31 VN.n30 19.674
R64 VN.n64 VN.n63 19.674
R65 VN.n16 VN.t0 17.0524
R66 VN.n7 VN.t8 17.0524
R67 VN.n23 VN.t3 17.0524
R68 VN.n31 VN.t5 17.0524
R69 VN.n49 VN.t1 17.0524
R70 VN.n40 VN.t2 17.0524
R71 VN.n56 VN.t9 17.0524
R72 VN.n64 VN.t4 17.0524
R73 VN.n42 VN.n41 8.9882
R74 VN.n9 VN.n8 8.9882
R75 VN.n24 VN.n23 2.45968
R76 VN.n57 VN.n56 2.45968
R77 VN.n65 VN.n33 0.278335
R78 VN.n32 VN.n0 0.278335
R79 VN.n61 VN.n33 0.189894
R80 VN.n61 VN.n60 0.189894
R81 VN.n60 VN.n59 0.189894
R82 VN.n59 VN.n35 0.189894
R83 VN.n54 VN.n35 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n52 0.189894
R86 VN.n52 VN.n37 0.189894
R87 VN.n48 VN.n37 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n46 0.189894
R90 VN.n46 VN.n39 0.189894
R91 VN.n42 VN.n39 0.189894
R92 VN.n9 VN.n6 0.189894
R93 VN.n13 VN.n6 0.189894
R94 VN.n14 VN.n13 0.189894
R95 VN.n15 VN.n14 0.189894
R96 VN.n15 VN.n4 0.189894
R97 VN.n19 VN.n4 0.189894
R98 VN.n20 VN.n19 0.189894
R99 VN.n21 VN.n20 0.189894
R100 VN.n21 VN.n2 0.189894
R101 VN.n26 VN.n2 0.189894
R102 VN.n27 VN.n26 0.189894
R103 VN.n28 VN.n27 0.189894
R104 VN.n28 VN.n0 0.189894
R105 VN VN.n32 0.153485
R106 VTAIL.n11 VTAIL.t17 114.085
R107 VTAIL.n17 VTAIL.t16 114.085
R108 VTAIL.n2 VTAIL.t6 114.085
R109 VTAIL.n16 VTAIL.t7 114.085
R110 VTAIL.n15 VTAIL.n14 100.885
R111 VTAIL.n13 VTAIL.n12 100.885
R112 VTAIL.n10 VTAIL.n9 100.885
R113 VTAIL.n8 VTAIL.n7 100.885
R114 VTAIL.n19 VTAIL.n18 100.885
R115 VTAIL.n1 VTAIL.n0 100.885
R116 VTAIL.n4 VTAIL.n3 100.885
R117 VTAIL.n6 VTAIL.n5 100.885
R118 VTAIL.n8 VTAIL.n6 17.8841
R119 VTAIL.n17 VTAIL.n16 15.7721
R120 VTAIL.n18 VTAIL.t11 13.2005
R121 VTAIL.n18 VTAIL.t10 13.2005
R122 VTAIL.n0 VTAIL.t19 13.2005
R123 VTAIL.n0 VTAIL.t13 13.2005
R124 VTAIL.n3 VTAIL.t2 13.2005
R125 VTAIL.n3 VTAIL.t5 13.2005
R126 VTAIL.n5 VTAIL.t1 13.2005
R127 VTAIL.n5 VTAIL.t4 13.2005
R128 VTAIL.n14 VTAIL.t0 13.2005
R129 VTAIL.n14 VTAIL.t3 13.2005
R130 VTAIL.n12 VTAIL.t8 13.2005
R131 VTAIL.n12 VTAIL.t9 13.2005
R132 VTAIL.n9 VTAIL.t12 13.2005
R133 VTAIL.n9 VTAIL.t15 13.2005
R134 VTAIL.n7 VTAIL.t18 13.2005
R135 VTAIL.n7 VTAIL.t14 13.2005
R136 VTAIL.n10 VTAIL.n8 2.11257
R137 VTAIL.n11 VTAIL.n10 2.11257
R138 VTAIL.n15 VTAIL.n13 2.11257
R139 VTAIL.n16 VTAIL.n15 2.11257
R140 VTAIL.n6 VTAIL.n4 2.11257
R141 VTAIL.n4 VTAIL.n2 2.11257
R142 VTAIL.n19 VTAIL.n17 2.11257
R143 VTAIL VTAIL.n1 1.64274
R144 VTAIL.n13 VTAIL.n11 1.52636
R145 VTAIL.n2 VTAIL.n1 1.52636
R146 VTAIL VTAIL.n19 0.470328
R147 VDD2.n1 VDD2.t2 132.876
R148 VDD2.n4 VDD2.t5 130.764
R149 VDD2.n3 VDD2.n2 119.093
R150 VDD2 VDD2.n7 119.09
R151 VDD2.n6 VDD2.n5 117.564
R152 VDD2.n1 VDD2.n0 117.564
R153 VDD2.n4 VDD2.n3 35.0407
R154 VDD2.n7 VDD2.t7 13.2005
R155 VDD2.n7 VDD2.t3 13.2005
R156 VDD2.n5 VDD2.t0 13.2005
R157 VDD2.n5 VDD2.t8 13.2005
R158 VDD2.n2 VDD2.t6 13.2005
R159 VDD2.n2 VDD2.t4 13.2005
R160 VDD2.n0 VDD2.t1 13.2005
R161 VDD2.n0 VDD2.t9 13.2005
R162 VDD2.n6 VDD2.n4 2.11257
R163 VDD2 VDD2.n6 0.586707
R164 VDD2.n3 VDD2.n1 0.473171
R165 B.n577 B.n576 585
R166 B.n578 B.n577 585
R167 B.n173 B.n111 585
R168 B.n172 B.n171 585
R169 B.n170 B.n169 585
R170 B.n168 B.n167 585
R171 B.n166 B.n165 585
R172 B.n164 B.n163 585
R173 B.n162 B.n161 585
R174 B.n160 B.n159 585
R175 B.n158 B.n157 585
R176 B.n156 B.n155 585
R177 B.n154 B.n153 585
R178 B.n152 B.n151 585
R179 B.n150 B.n149 585
R180 B.n148 B.n147 585
R181 B.n146 B.n145 585
R182 B.n144 B.n143 585
R183 B.n142 B.n141 585
R184 B.n140 B.n139 585
R185 B.n138 B.n137 585
R186 B.n135 B.n134 585
R187 B.n133 B.n132 585
R188 B.n131 B.n130 585
R189 B.n129 B.n128 585
R190 B.n127 B.n126 585
R191 B.n125 B.n124 585
R192 B.n123 B.n122 585
R193 B.n121 B.n120 585
R194 B.n119 B.n118 585
R195 B.n96 B.n95 585
R196 B.n581 B.n580 585
R197 B.n575 B.n112 585
R198 B.n112 B.n93 585
R199 B.n574 B.n92 585
R200 B.n585 B.n92 585
R201 B.n573 B.n91 585
R202 B.n586 B.n91 585
R203 B.n572 B.n90 585
R204 B.n587 B.n90 585
R205 B.n571 B.n570 585
R206 B.n570 B.n86 585
R207 B.n569 B.n85 585
R208 B.n593 B.n85 585
R209 B.n568 B.n84 585
R210 B.n594 B.n84 585
R211 B.n567 B.n83 585
R212 B.n595 B.n83 585
R213 B.n566 B.n565 585
R214 B.n565 B.n79 585
R215 B.n564 B.n78 585
R216 B.n601 B.n78 585
R217 B.n563 B.n77 585
R218 B.n602 B.n77 585
R219 B.n562 B.n76 585
R220 B.n603 B.n76 585
R221 B.n561 B.n560 585
R222 B.n560 B.n72 585
R223 B.n559 B.n71 585
R224 B.n609 B.n71 585
R225 B.n558 B.n70 585
R226 B.n610 B.n70 585
R227 B.n557 B.n69 585
R228 B.n611 B.n69 585
R229 B.n556 B.n555 585
R230 B.n555 B.n65 585
R231 B.n554 B.n64 585
R232 B.n617 B.n64 585
R233 B.n553 B.n63 585
R234 B.n618 B.n63 585
R235 B.n552 B.n62 585
R236 B.n619 B.n62 585
R237 B.n551 B.n550 585
R238 B.n550 B.n58 585
R239 B.n549 B.n57 585
R240 B.n625 B.n57 585
R241 B.n548 B.n56 585
R242 B.n626 B.n56 585
R243 B.n547 B.n55 585
R244 B.n627 B.n55 585
R245 B.n546 B.n545 585
R246 B.n545 B.n54 585
R247 B.n544 B.n50 585
R248 B.n633 B.n50 585
R249 B.n543 B.n49 585
R250 B.n634 B.n49 585
R251 B.n542 B.n48 585
R252 B.n635 B.n48 585
R253 B.n541 B.n540 585
R254 B.n540 B.n44 585
R255 B.n539 B.n43 585
R256 B.n641 B.n43 585
R257 B.n538 B.n42 585
R258 B.n642 B.n42 585
R259 B.n537 B.n41 585
R260 B.n643 B.n41 585
R261 B.n536 B.n535 585
R262 B.n535 B.n37 585
R263 B.n534 B.n36 585
R264 B.n649 B.n36 585
R265 B.n533 B.n35 585
R266 B.n650 B.n35 585
R267 B.n532 B.n34 585
R268 B.n651 B.n34 585
R269 B.n531 B.n530 585
R270 B.n530 B.n30 585
R271 B.n529 B.n29 585
R272 B.n657 B.n29 585
R273 B.n528 B.n28 585
R274 B.n658 B.n28 585
R275 B.n527 B.n27 585
R276 B.n659 B.n27 585
R277 B.n526 B.n525 585
R278 B.n525 B.n23 585
R279 B.n524 B.n22 585
R280 B.n665 B.n22 585
R281 B.n523 B.n21 585
R282 B.n666 B.n21 585
R283 B.n522 B.n20 585
R284 B.n667 B.n20 585
R285 B.n521 B.n520 585
R286 B.n520 B.n16 585
R287 B.n519 B.n15 585
R288 B.n673 B.n15 585
R289 B.n518 B.n14 585
R290 B.n674 B.n14 585
R291 B.n517 B.n13 585
R292 B.n675 B.n13 585
R293 B.n516 B.n515 585
R294 B.n515 B.n12 585
R295 B.n514 B.n513 585
R296 B.n514 B.n8 585
R297 B.n512 B.n7 585
R298 B.n682 B.n7 585
R299 B.n511 B.n6 585
R300 B.n683 B.n6 585
R301 B.n510 B.n5 585
R302 B.n684 B.n5 585
R303 B.n509 B.n508 585
R304 B.n508 B.n4 585
R305 B.n507 B.n174 585
R306 B.n507 B.n506 585
R307 B.n497 B.n175 585
R308 B.n176 B.n175 585
R309 B.n499 B.n498 585
R310 B.n500 B.n499 585
R311 B.n496 B.n180 585
R312 B.n184 B.n180 585
R313 B.n495 B.n494 585
R314 B.n494 B.n493 585
R315 B.n182 B.n181 585
R316 B.n183 B.n182 585
R317 B.n486 B.n485 585
R318 B.n487 B.n486 585
R319 B.n484 B.n189 585
R320 B.n189 B.n188 585
R321 B.n483 B.n482 585
R322 B.n482 B.n481 585
R323 B.n191 B.n190 585
R324 B.n192 B.n191 585
R325 B.n474 B.n473 585
R326 B.n475 B.n474 585
R327 B.n472 B.n197 585
R328 B.n197 B.n196 585
R329 B.n471 B.n470 585
R330 B.n470 B.n469 585
R331 B.n199 B.n198 585
R332 B.n200 B.n199 585
R333 B.n462 B.n461 585
R334 B.n463 B.n462 585
R335 B.n460 B.n205 585
R336 B.n205 B.n204 585
R337 B.n459 B.n458 585
R338 B.n458 B.n457 585
R339 B.n207 B.n206 585
R340 B.n208 B.n207 585
R341 B.n450 B.n449 585
R342 B.n451 B.n450 585
R343 B.n448 B.n213 585
R344 B.n213 B.n212 585
R345 B.n447 B.n446 585
R346 B.n446 B.n445 585
R347 B.n215 B.n214 585
R348 B.n216 B.n215 585
R349 B.n438 B.n437 585
R350 B.n439 B.n438 585
R351 B.n436 B.n221 585
R352 B.n221 B.n220 585
R353 B.n435 B.n434 585
R354 B.n434 B.n433 585
R355 B.n223 B.n222 585
R356 B.n426 B.n223 585
R357 B.n425 B.n424 585
R358 B.n427 B.n425 585
R359 B.n423 B.n228 585
R360 B.n228 B.n227 585
R361 B.n422 B.n421 585
R362 B.n421 B.n420 585
R363 B.n230 B.n229 585
R364 B.n231 B.n230 585
R365 B.n413 B.n412 585
R366 B.n414 B.n413 585
R367 B.n411 B.n236 585
R368 B.n236 B.n235 585
R369 B.n410 B.n409 585
R370 B.n409 B.n408 585
R371 B.n238 B.n237 585
R372 B.n239 B.n238 585
R373 B.n401 B.n400 585
R374 B.n402 B.n401 585
R375 B.n399 B.n244 585
R376 B.n244 B.n243 585
R377 B.n398 B.n397 585
R378 B.n397 B.n396 585
R379 B.n246 B.n245 585
R380 B.n247 B.n246 585
R381 B.n389 B.n388 585
R382 B.n390 B.n389 585
R383 B.n387 B.n252 585
R384 B.n252 B.n251 585
R385 B.n386 B.n385 585
R386 B.n385 B.n384 585
R387 B.n254 B.n253 585
R388 B.n255 B.n254 585
R389 B.n377 B.n376 585
R390 B.n378 B.n377 585
R391 B.n375 B.n260 585
R392 B.n260 B.n259 585
R393 B.n374 B.n373 585
R394 B.n373 B.n372 585
R395 B.n262 B.n261 585
R396 B.n263 B.n262 585
R397 B.n365 B.n364 585
R398 B.n366 B.n365 585
R399 B.n363 B.n268 585
R400 B.n268 B.n267 585
R401 B.n362 B.n361 585
R402 B.n361 B.n360 585
R403 B.n270 B.n269 585
R404 B.n271 B.n270 585
R405 B.n356 B.n355 585
R406 B.n274 B.n273 585
R407 B.n352 B.n351 585
R408 B.n353 B.n352 585
R409 B.n350 B.n289 585
R410 B.n349 B.n348 585
R411 B.n347 B.n346 585
R412 B.n345 B.n344 585
R413 B.n343 B.n342 585
R414 B.n341 B.n340 585
R415 B.n339 B.n338 585
R416 B.n337 B.n336 585
R417 B.n335 B.n334 585
R418 B.n333 B.n332 585
R419 B.n331 B.n330 585
R420 B.n329 B.n328 585
R421 B.n327 B.n326 585
R422 B.n325 B.n324 585
R423 B.n323 B.n322 585
R424 B.n321 B.n320 585
R425 B.n319 B.n318 585
R426 B.n316 B.n315 585
R427 B.n314 B.n313 585
R428 B.n312 B.n311 585
R429 B.n310 B.n309 585
R430 B.n308 B.n307 585
R431 B.n306 B.n305 585
R432 B.n304 B.n303 585
R433 B.n302 B.n301 585
R434 B.n300 B.n299 585
R435 B.n298 B.n297 585
R436 B.n296 B.n295 585
R437 B.n357 B.n272 585
R438 B.n272 B.n271 585
R439 B.n359 B.n358 585
R440 B.n360 B.n359 585
R441 B.n266 B.n265 585
R442 B.n267 B.n266 585
R443 B.n368 B.n367 585
R444 B.n367 B.n366 585
R445 B.n369 B.n264 585
R446 B.n264 B.n263 585
R447 B.n371 B.n370 585
R448 B.n372 B.n371 585
R449 B.n258 B.n257 585
R450 B.n259 B.n258 585
R451 B.n380 B.n379 585
R452 B.n379 B.n378 585
R453 B.n381 B.n256 585
R454 B.n256 B.n255 585
R455 B.n383 B.n382 585
R456 B.n384 B.n383 585
R457 B.n250 B.n249 585
R458 B.n251 B.n250 585
R459 B.n392 B.n391 585
R460 B.n391 B.n390 585
R461 B.n393 B.n248 585
R462 B.n248 B.n247 585
R463 B.n395 B.n394 585
R464 B.n396 B.n395 585
R465 B.n242 B.n241 585
R466 B.n243 B.n242 585
R467 B.n404 B.n403 585
R468 B.n403 B.n402 585
R469 B.n405 B.n240 585
R470 B.n240 B.n239 585
R471 B.n407 B.n406 585
R472 B.n408 B.n407 585
R473 B.n234 B.n233 585
R474 B.n235 B.n234 585
R475 B.n416 B.n415 585
R476 B.n415 B.n414 585
R477 B.n417 B.n232 585
R478 B.n232 B.n231 585
R479 B.n419 B.n418 585
R480 B.n420 B.n419 585
R481 B.n226 B.n225 585
R482 B.n227 B.n226 585
R483 B.n429 B.n428 585
R484 B.n428 B.n427 585
R485 B.n430 B.n224 585
R486 B.n426 B.n224 585
R487 B.n432 B.n431 585
R488 B.n433 B.n432 585
R489 B.n219 B.n218 585
R490 B.n220 B.n219 585
R491 B.n441 B.n440 585
R492 B.n440 B.n439 585
R493 B.n442 B.n217 585
R494 B.n217 B.n216 585
R495 B.n444 B.n443 585
R496 B.n445 B.n444 585
R497 B.n211 B.n210 585
R498 B.n212 B.n211 585
R499 B.n453 B.n452 585
R500 B.n452 B.n451 585
R501 B.n454 B.n209 585
R502 B.n209 B.n208 585
R503 B.n456 B.n455 585
R504 B.n457 B.n456 585
R505 B.n203 B.n202 585
R506 B.n204 B.n203 585
R507 B.n465 B.n464 585
R508 B.n464 B.n463 585
R509 B.n466 B.n201 585
R510 B.n201 B.n200 585
R511 B.n468 B.n467 585
R512 B.n469 B.n468 585
R513 B.n195 B.n194 585
R514 B.n196 B.n195 585
R515 B.n477 B.n476 585
R516 B.n476 B.n475 585
R517 B.n478 B.n193 585
R518 B.n193 B.n192 585
R519 B.n480 B.n479 585
R520 B.n481 B.n480 585
R521 B.n187 B.n186 585
R522 B.n188 B.n187 585
R523 B.n489 B.n488 585
R524 B.n488 B.n487 585
R525 B.n490 B.n185 585
R526 B.n185 B.n183 585
R527 B.n492 B.n491 585
R528 B.n493 B.n492 585
R529 B.n179 B.n178 585
R530 B.n184 B.n179 585
R531 B.n502 B.n501 585
R532 B.n501 B.n500 585
R533 B.n503 B.n177 585
R534 B.n177 B.n176 585
R535 B.n505 B.n504 585
R536 B.n506 B.n505 585
R537 B.n3 B.n0 585
R538 B.n4 B.n3 585
R539 B.n681 B.n1 585
R540 B.n682 B.n681 585
R541 B.n680 B.n679 585
R542 B.n680 B.n8 585
R543 B.n678 B.n9 585
R544 B.n12 B.n9 585
R545 B.n677 B.n676 585
R546 B.n676 B.n675 585
R547 B.n11 B.n10 585
R548 B.n674 B.n11 585
R549 B.n672 B.n671 585
R550 B.n673 B.n672 585
R551 B.n670 B.n17 585
R552 B.n17 B.n16 585
R553 B.n669 B.n668 585
R554 B.n668 B.n667 585
R555 B.n19 B.n18 585
R556 B.n666 B.n19 585
R557 B.n664 B.n663 585
R558 B.n665 B.n664 585
R559 B.n662 B.n24 585
R560 B.n24 B.n23 585
R561 B.n661 B.n660 585
R562 B.n660 B.n659 585
R563 B.n26 B.n25 585
R564 B.n658 B.n26 585
R565 B.n656 B.n655 585
R566 B.n657 B.n656 585
R567 B.n654 B.n31 585
R568 B.n31 B.n30 585
R569 B.n653 B.n652 585
R570 B.n652 B.n651 585
R571 B.n33 B.n32 585
R572 B.n650 B.n33 585
R573 B.n648 B.n647 585
R574 B.n649 B.n648 585
R575 B.n646 B.n38 585
R576 B.n38 B.n37 585
R577 B.n645 B.n644 585
R578 B.n644 B.n643 585
R579 B.n40 B.n39 585
R580 B.n642 B.n40 585
R581 B.n640 B.n639 585
R582 B.n641 B.n640 585
R583 B.n638 B.n45 585
R584 B.n45 B.n44 585
R585 B.n637 B.n636 585
R586 B.n636 B.n635 585
R587 B.n47 B.n46 585
R588 B.n634 B.n47 585
R589 B.n632 B.n631 585
R590 B.n633 B.n632 585
R591 B.n630 B.n51 585
R592 B.n54 B.n51 585
R593 B.n629 B.n628 585
R594 B.n628 B.n627 585
R595 B.n53 B.n52 585
R596 B.n626 B.n53 585
R597 B.n624 B.n623 585
R598 B.n625 B.n624 585
R599 B.n622 B.n59 585
R600 B.n59 B.n58 585
R601 B.n621 B.n620 585
R602 B.n620 B.n619 585
R603 B.n61 B.n60 585
R604 B.n618 B.n61 585
R605 B.n616 B.n615 585
R606 B.n617 B.n616 585
R607 B.n614 B.n66 585
R608 B.n66 B.n65 585
R609 B.n613 B.n612 585
R610 B.n612 B.n611 585
R611 B.n68 B.n67 585
R612 B.n610 B.n68 585
R613 B.n608 B.n607 585
R614 B.n609 B.n608 585
R615 B.n606 B.n73 585
R616 B.n73 B.n72 585
R617 B.n605 B.n604 585
R618 B.n604 B.n603 585
R619 B.n75 B.n74 585
R620 B.n602 B.n75 585
R621 B.n600 B.n599 585
R622 B.n601 B.n600 585
R623 B.n598 B.n80 585
R624 B.n80 B.n79 585
R625 B.n597 B.n596 585
R626 B.n596 B.n595 585
R627 B.n82 B.n81 585
R628 B.n594 B.n82 585
R629 B.n592 B.n591 585
R630 B.n593 B.n592 585
R631 B.n590 B.n87 585
R632 B.n87 B.n86 585
R633 B.n589 B.n588 585
R634 B.n588 B.n587 585
R635 B.n89 B.n88 585
R636 B.n586 B.n89 585
R637 B.n584 B.n583 585
R638 B.n585 B.n584 585
R639 B.n582 B.n94 585
R640 B.n94 B.n93 585
R641 B.n685 B.n684 585
R642 B.n683 B.n2 585
R643 B.n580 B.n94 478.086
R644 B.n577 B.n112 478.086
R645 B.n295 B.n270 478.086
R646 B.n355 B.n272 478.086
R647 B.n578 B.n110 256.663
R648 B.n578 B.n109 256.663
R649 B.n578 B.n108 256.663
R650 B.n578 B.n107 256.663
R651 B.n578 B.n106 256.663
R652 B.n578 B.n105 256.663
R653 B.n578 B.n104 256.663
R654 B.n578 B.n103 256.663
R655 B.n578 B.n102 256.663
R656 B.n578 B.n101 256.663
R657 B.n578 B.n100 256.663
R658 B.n578 B.n99 256.663
R659 B.n578 B.n98 256.663
R660 B.n578 B.n97 256.663
R661 B.n579 B.n578 256.663
R662 B.n354 B.n353 256.663
R663 B.n353 B.n275 256.663
R664 B.n353 B.n276 256.663
R665 B.n353 B.n277 256.663
R666 B.n353 B.n278 256.663
R667 B.n353 B.n279 256.663
R668 B.n353 B.n280 256.663
R669 B.n353 B.n281 256.663
R670 B.n353 B.n282 256.663
R671 B.n353 B.n283 256.663
R672 B.n353 B.n284 256.663
R673 B.n353 B.n285 256.663
R674 B.n353 B.n286 256.663
R675 B.n353 B.n287 256.663
R676 B.n353 B.n288 256.663
R677 B.n687 B.n686 256.663
R678 B.n116 B.t21 224.238
R679 B.n113 B.t17 224.238
R680 B.n293 B.t14 224.238
R681 B.n290 B.t10 224.238
R682 B.n353 B.n271 183.47
R683 B.n578 B.n93 183.47
R684 B.n118 B.n96 163.367
R685 B.n122 B.n121 163.367
R686 B.n126 B.n125 163.367
R687 B.n130 B.n129 163.367
R688 B.n134 B.n133 163.367
R689 B.n139 B.n138 163.367
R690 B.n143 B.n142 163.367
R691 B.n147 B.n146 163.367
R692 B.n151 B.n150 163.367
R693 B.n155 B.n154 163.367
R694 B.n159 B.n158 163.367
R695 B.n163 B.n162 163.367
R696 B.n167 B.n166 163.367
R697 B.n171 B.n170 163.367
R698 B.n577 B.n111 163.367
R699 B.n361 B.n270 163.367
R700 B.n361 B.n268 163.367
R701 B.n365 B.n268 163.367
R702 B.n365 B.n262 163.367
R703 B.n373 B.n262 163.367
R704 B.n373 B.n260 163.367
R705 B.n377 B.n260 163.367
R706 B.n377 B.n254 163.367
R707 B.n385 B.n254 163.367
R708 B.n385 B.n252 163.367
R709 B.n389 B.n252 163.367
R710 B.n389 B.n246 163.367
R711 B.n397 B.n246 163.367
R712 B.n397 B.n244 163.367
R713 B.n401 B.n244 163.367
R714 B.n401 B.n238 163.367
R715 B.n409 B.n238 163.367
R716 B.n409 B.n236 163.367
R717 B.n413 B.n236 163.367
R718 B.n413 B.n230 163.367
R719 B.n421 B.n230 163.367
R720 B.n421 B.n228 163.367
R721 B.n425 B.n228 163.367
R722 B.n425 B.n223 163.367
R723 B.n434 B.n223 163.367
R724 B.n434 B.n221 163.367
R725 B.n438 B.n221 163.367
R726 B.n438 B.n215 163.367
R727 B.n446 B.n215 163.367
R728 B.n446 B.n213 163.367
R729 B.n450 B.n213 163.367
R730 B.n450 B.n207 163.367
R731 B.n458 B.n207 163.367
R732 B.n458 B.n205 163.367
R733 B.n462 B.n205 163.367
R734 B.n462 B.n199 163.367
R735 B.n470 B.n199 163.367
R736 B.n470 B.n197 163.367
R737 B.n474 B.n197 163.367
R738 B.n474 B.n191 163.367
R739 B.n482 B.n191 163.367
R740 B.n482 B.n189 163.367
R741 B.n486 B.n189 163.367
R742 B.n486 B.n182 163.367
R743 B.n494 B.n182 163.367
R744 B.n494 B.n180 163.367
R745 B.n499 B.n180 163.367
R746 B.n499 B.n175 163.367
R747 B.n507 B.n175 163.367
R748 B.n508 B.n507 163.367
R749 B.n508 B.n5 163.367
R750 B.n6 B.n5 163.367
R751 B.n7 B.n6 163.367
R752 B.n514 B.n7 163.367
R753 B.n515 B.n514 163.367
R754 B.n515 B.n13 163.367
R755 B.n14 B.n13 163.367
R756 B.n15 B.n14 163.367
R757 B.n520 B.n15 163.367
R758 B.n520 B.n20 163.367
R759 B.n21 B.n20 163.367
R760 B.n22 B.n21 163.367
R761 B.n525 B.n22 163.367
R762 B.n525 B.n27 163.367
R763 B.n28 B.n27 163.367
R764 B.n29 B.n28 163.367
R765 B.n530 B.n29 163.367
R766 B.n530 B.n34 163.367
R767 B.n35 B.n34 163.367
R768 B.n36 B.n35 163.367
R769 B.n535 B.n36 163.367
R770 B.n535 B.n41 163.367
R771 B.n42 B.n41 163.367
R772 B.n43 B.n42 163.367
R773 B.n540 B.n43 163.367
R774 B.n540 B.n48 163.367
R775 B.n49 B.n48 163.367
R776 B.n50 B.n49 163.367
R777 B.n545 B.n50 163.367
R778 B.n545 B.n55 163.367
R779 B.n56 B.n55 163.367
R780 B.n57 B.n56 163.367
R781 B.n550 B.n57 163.367
R782 B.n550 B.n62 163.367
R783 B.n63 B.n62 163.367
R784 B.n64 B.n63 163.367
R785 B.n555 B.n64 163.367
R786 B.n555 B.n69 163.367
R787 B.n70 B.n69 163.367
R788 B.n71 B.n70 163.367
R789 B.n560 B.n71 163.367
R790 B.n560 B.n76 163.367
R791 B.n77 B.n76 163.367
R792 B.n78 B.n77 163.367
R793 B.n565 B.n78 163.367
R794 B.n565 B.n83 163.367
R795 B.n84 B.n83 163.367
R796 B.n85 B.n84 163.367
R797 B.n570 B.n85 163.367
R798 B.n570 B.n90 163.367
R799 B.n91 B.n90 163.367
R800 B.n92 B.n91 163.367
R801 B.n112 B.n92 163.367
R802 B.n352 B.n274 163.367
R803 B.n352 B.n289 163.367
R804 B.n348 B.n347 163.367
R805 B.n344 B.n343 163.367
R806 B.n340 B.n339 163.367
R807 B.n336 B.n335 163.367
R808 B.n332 B.n331 163.367
R809 B.n328 B.n327 163.367
R810 B.n324 B.n323 163.367
R811 B.n320 B.n319 163.367
R812 B.n315 B.n314 163.367
R813 B.n311 B.n310 163.367
R814 B.n307 B.n306 163.367
R815 B.n303 B.n302 163.367
R816 B.n299 B.n298 163.367
R817 B.n359 B.n272 163.367
R818 B.n359 B.n266 163.367
R819 B.n367 B.n266 163.367
R820 B.n367 B.n264 163.367
R821 B.n371 B.n264 163.367
R822 B.n371 B.n258 163.367
R823 B.n379 B.n258 163.367
R824 B.n379 B.n256 163.367
R825 B.n383 B.n256 163.367
R826 B.n383 B.n250 163.367
R827 B.n391 B.n250 163.367
R828 B.n391 B.n248 163.367
R829 B.n395 B.n248 163.367
R830 B.n395 B.n242 163.367
R831 B.n403 B.n242 163.367
R832 B.n403 B.n240 163.367
R833 B.n407 B.n240 163.367
R834 B.n407 B.n234 163.367
R835 B.n415 B.n234 163.367
R836 B.n415 B.n232 163.367
R837 B.n419 B.n232 163.367
R838 B.n419 B.n226 163.367
R839 B.n428 B.n226 163.367
R840 B.n428 B.n224 163.367
R841 B.n432 B.n224 163.367
R842 B.n432 B.n219 163.367
R843 B.n440 B.n219 163.367
R844 B.n440 B.n217 163.367
R845 B.n444 B.n217 163.367
R846 B.n444 B.n211 163.367
R847 B.n452 B.n211 163.367
R848 B.n452 B.n209 163.367
R849 B.n456 B.n209 163.367
R850 B.n456 B.n203 163.367
R851 B.n464 B.n203 163.367
R852 B.n464 B.n201 163.367
R853 B.n468 B.n201 163.367
R854 B.n468 B.n195 163.367
R855 B.n476 B.n195 163.367
R856 B.n476 B.n193 163.367
R857 B.n480 B.n193 163.367
R858 B.n480 B.n187 163.367
R859 B.n488 B.n187 163.367
R860 B.n488 B.n185 163.367
R861 B.n492 B.n185 163.367
R862 B.n492 B.n179 163.367
R863 B.n501 B.n179 163.367
R864 B.n501 B.n177 163.367
R865 B.n505 B.n177 163.367
R866 B.n505 B.n3 163.367
R867 B.n685 B.n3 163.367
R868 B.n681 B.n2 163.367
R869 B.n681 B.n680 163.367
R870 B.n680 B.n9 163.367
R871 B.n676 B.n9 163.367
R872 B.n676 B.n11 163.367
R873 B.n672 B.n11 163.367
R874 B.n672 B.n17 163.367
R875 B.n668 B.n17 163.367
R876 B.n668 B.n19 163.367
R877 B.n664 B.n19 163.367
R878 B.n664 B.n24 163.367
R879 B.n660 B.n24 163.367
R880 B.n660 B.n26 163.367
R881 B.n656 B.n26 163.367
R882 B.n656 B.n31 163.367
R883 B.n652 B.n31 163.367
R884 B.n652 B.n33 163.367
R885 B.n648 B.n33 163.367
R886 B.n648 B.n38 163.367
R887 B.n644 B.n38 163.367
R888 B.n644 B.n40 163.367
R889 B.n640 B.n40 163.367
R890 B.n640 B.n45 163.367
R891 B.n636 B.n45 163.367
R892 B.n636 B.n47 163.367
R893 B.n632 B.n47 163.367
R894 B.n632 B.n51 163.367
R895 B.n628 B.n51 163.367
R896 B.n628 B.n53 163.367
R897 B.n624 B.n53 163.367
R898 B.n624 B.n59 163.367
R899 B.n620 B.n59 163.367
R900 B.n620 B.n61 163.367
R901 B.n616 B.n61 163.367
R902 B.n616 B.n66 163.367
R903 B.n612 B.n66 163.367
R904 B.n612 B.n68 163.367
R905 B.n608 B.n68 163.367
R906 B.n608 B.n73 163.367
R907 B.n604 B.n73 163.367
R908 B.n604 B.n75 163.367
R909 B.n600 B.n75 163.367
R910 B.n600 B.n80 163.367
R911 B.n596 B.n80 163.367
R912 B.n596 B.n82 163.367
R913 B.n592 B.n82 163.367
R914 B.n592 B.n87 163.367
R915 B.n588 B.n87 163.367
R916 B.n588 B.n89 163.367
R917 B.n584 B.n89 163.367
R918 B.n584 B.n94 163.367
R919 B.n113 B.t19 154.855
R920 B.n293 B.t16 154.855
R921 B.n116 B.t22 154.855
R922 B.n290 B.t13 154.855
R923 B.n360 B.n271 110.406
R924 B.n360 B.n267 110.406
R925 B.n366 B.n267 110.406
R926 B.n366 B.n263 110.406
R927 B.n372 B.n263 110.406
R928 B.n372 B.n259 110.406
R929 B.n378 B.n259 110.406
R930 B.n384 B.n255 110.406
R931 B.n384 B.n251 110.406
R932 B.n390 B.n251 110.406
R933 B.n390 B.n247 110.406
R934 B.n396 B.n247 110.406
R935 B.n396 B.n243 110.406
R936 B.n402 B.n243 110.406
R937 B.n402 B.n239 110.406
R938 B.n408 B.n239 110.406
R939 B.n414 B.n235 110.406
R940 B.n414 B.n231 110.406
R941 B.n420 B.n231 110.406
R942 B.n420 B.n227 110.406
R943 B.n427 B.n227 110.406
R944 B.n427 B.n426 110.406
R945 B.n433 B.n220 110.406
R946 B.n439 B.n220 110.406
R947 B.n439 B.n216 110.406
R948 B.n445 B.n216 110.406
R949 B.n445 B.n212 110.406
R950 B.n451 B.n212 110.406
R951 B.n457 B.n208 110.406
R952 B.n457 B.n204 110.406
R953 B.n463 B.n204 110.406
R954 B.n463 B.n200 110.406
R955 B.n469 B.n200 110.406
R956 B.n469 B.n196 110.406
R957 B.n475 B.n196 110.406
R958 B.n481 B.n192 110.406
R959 B.n481 B.n188 110.406
R960 B.n487 B.n188 110.406
R961 B.n487 B.n183 110.406
R962 B.n493 B.n183 110.406
R963 B.n493 B.n184 110.406
R964 B.n500 B.n176 110.406
R965 B.n506 B.n176 110.406
R966 B.n506 B.n4 110.406
R967 B.n684 B.n4 110.406
R968 B.n684 B.n683 110.406
R969 B.n683 B.n682 110.406
R970 B.n682 B.n8 110.406
R971 B.n12 B.n8 110.406
R972 B.n675 B.n12 110.406
R973 B.n674 B.n673 110.406
R974 B.n673 B.n16 110.406
R975 B.n667 B.n16 110.406
R976 B.n667 B.n666 110.406
R977 B.n666 B.n665 110.406
R978 B.n665 B.n23 110.406
R979 B.n659 B.n658 110.406
R980 B.n658 B.n657 110.406
R981 B.n657 B.n30 110.406
R982 B.n651 B.n30 110.406
R983 B.n651 B.n650 110.406
R984 B.n650 B.n649 110.406
R985 B.n649 B.n37 110.406
R986 B.n643 B.n642 110.406
R987 B.n642 B.n641 110.406
R988 B.n641 B.n44 110.406
R989 B.n635 B.n44 110.406
R990 B.n635 B.n634 110.406
R991 B.n634 B.n633 110.406
R992 B.n627 B.n54 110.406
R993 B.n627 B.n626 110.406
R994 B.n626 B.n625 110.406
R995 B.n625 B.n58 110.406
R996 B.n619 B.n58 110.406
R997 B.n619 B.n618 110.406
R998 B.n617 B.n65 110.406
R999 B.n611 B.n65 110.406
R1000 B.n611 B.n610 110.406
R1001 B.n610 B.n609 110.406
R1002 B.n609 B.n72 110.406
R1003 B.n603 B.n72 110.406
R1004 B.n603 B.n602 110.406
R1005 B.n602 B.n601 110.406
R1006 B.n601 B.n79 110.406
R1007 B.n595 B.n594 110.406
R1008 B.n594 B.n593 110.406
R1009 B.n593 B.n86 110.406
R1010 B.n587 B.n86 110.406
R1011 B.n587 B.n586 110.406
R1012 B.n586 B.n585 110.406
R1013 B.n585 B.n93 110.406
R1014 B.n114 B.t20 107.34
R1015 B.n294 B.t15 107.34
R1016 B.n117 B.t23 107.338
R1017 B.n291 B.t12 107.338
R1018 B.t11 B.n255 103.912
R1019 B.t18 B.n79 103.912
R1020 B.t5 B.n192 100.665
R1021 B.t9 B.n23 100.665
R1022 B.n451 B.t2 97.4175
R1023 B.n643 B.t0 97.4175
R1024 B.n500 B.t6 77.9341
R1025 B.n675 B.t8 77.9341
R1026 B.n426 B.t4 74.6868
R1027 B.n54 B.t3 74.6868
R1028 B.n580 B.n579 71.676
R1029 B.n118 B.n97 71.676
R1030 B.n122 B.n98 71.676
R1031 B.n126 B.n99 71.676
R1032 B.n130 B.n100 71.676
R1033 B.n134 B.n101 71.676
R1034 B.n139 B.n102 71.676
R1035 B.n143 B.n103 71.676
R1036 B.n147 B.n104 71.676
R1037 B.n151 B.n105 71.676
R1038 B.n155 B.n106 71.676
R1039 B.n159 B.n107 71.676
R1040 B.n163 B.n108 71.676
R1041 B.n167 B.n109 71.676
R1042 B.n171 B.n110 71.676
R1043 B.n111 B.n110 71.676
R1044 B.n170 B.n109 71.676
R1045 B.n166 B.n108 71.676
R1046 B.n162 B.n107 71.676
R1047 B.n158 B.n106 71.676
R1048 B.n154 B.n105 71.676
R1049 B.n150 B.n104 71.676
R1050 B.n146 B.n103 71.676
R1051 B.n142 B.n102 71.676
R1052 B.n138 B.n101 71.676
R1053 B.n133 B.n100 71.676
R1054 B.n129 B.n99 71.676
R1055 B.n125 B.n98 71.676
R1056 B.n121 B.n97 71.676
R1057 B.n579 B.n96 71.676
R1058 B.n355 B.n354 71.676
R1059 B.n289 B.n275 71.676
R1060 B.n347 B.n276 71.676
R1061 B.n343 B.n277 71.676
R1062 B.n339 B.n278 71.676
R1063 B.n335 B.n279 71.676
R1064 B.n331 B.n280 71.676
R1065 B.n327 B.n281 71.676
R1066 B.n323 B.n282 71.676
R1067 B.n319 B.n283 71.676
R1068 B.n314 B.n284 71.676
R1069 B.n310 B.n285 71.676
R1070 B.n306 B.n286 71.676
R1071 B.n302 B.n287 71.676
R1072 B.n298 B.n288 71.676
R1073 B.n354 B.n274 71.676
R1074 B.n348 B.n275 71.676
R1075 B.n344 B.n276 71.676
R1076 B.n340 B.n277 71.676
R1077 B.n336 B.n278 71.676
R1078 B.n332 B.n279 71.676
R1079 B.n328 B.n280 71.676
R1080 B.n324 B.n281 71.676
R1081 B.n320 B.n282 71.676
R1082 B.n315 B.n283 71.676
R1083 B.n311 B.n284 71.676
R1084 B.n307 B.n285 71.676
R1085 B.n303 B.n286 71.676
R1086 B.n299 B.n287 71.676
R1087 B.n295 B.n288 71.676
R1088 B.n686 B.n685 71.676
R1089 B.n686 B.n2 71.676
R1090 B.n136 B.n117 59.5399
R1091 B.n115 B.n114 59.5399
R1092 B.n317 B.n294 59.5399
R1093 B.n292 B.n291 59.5399
R1094 B.t1 B.n235 58.4507
R1095 B.n618 B.t7 58.4507
R1096 B.n408 B.t1 51.9562
R1097 B.t7 B.n617 51.9562
R1098 B.n117 B.n116 47.5157
R1099 B.n114 B.n113 47.5157
R1100 B.n294 B.n293 47.5157
R1101 B.n291 B.n290 47.5157
R1102 B.n433 B.t4 35.7201
R1103 B.n633 B.t3 35.7201
R1104 B.n184 B.t6 32.4728
R1105 B.t8 B.n674 32.4728
R1106 B.n357 B.n356 31.0639
R1107 B.n296 B.n269 31.0639
R1108 B.n576 B.n575 31.0639
R1109 B.n582 B.n581 31.0639
R1110 B B.n687 18.0485
R1111 B.t2 B.n208 12.9894
R1112 B.t0 B.n37 12.9894
R1113 B.n358 B.n357 10.6151
R1114 B.n358 B.n265 10.6151
R1115 B.n368 B.n265 10.6151
R1116 B.n369 B.n368 10.6151
R1117 B.n370 B.n369 10.6151
R1118 B.n370 B.n257 10.6151
R1119 B.n380 B.n257 10.6151
R1120 B.n381 B.n380 10.6151
R1121 B.n382 B.n381 10.6151
R1122 B.n382 B.n249 10.6151
R1123 B.n392 B.n249 10.6151
R1124 B.n393 B.n392 10.6151
R1125 B.n394 B.n393 10.6151
R1126 B.n394 B.n241 10.6151
R1127 B.n404 B.n241 10.6151
R1128 B.n405 B.n404 10.6151
R1129 B.n406 B.n405 10.6151
R1130 B.n406 B.n233 10.6151
R1131 B.n416 B.n233 10.6151
R1132 B.n417 B.n416 10.6151
R1133 B.n418 B.n417 10.6151
R1134 B.n418 B.n225 10.6151
R1135 B.n429 B.n225 10.6151
R1136 B.n430 B.n429 10.6151
R1137 B.n431 B.n430 10.6151
R1138 B.n431 B.n218 10.6151
R1139 B.n441 B.n218 10.6151
R1140 B.n442 B.n441 10.6151
R1141 B.n443 B.n442 10.6151
R1142 B.n443 B.n210 10.6151
R1143 B.n453 B.n210 10.6151
R1144 B.n454 B.n453 10.6151
R1145 B.n455 B.n454 10.6151
R1146 B.n455 B.n202 10.6151
R1147 B.n465 B.n202 10.6151
R1148 B.n466 B.n465 10.6151
R1149 B.n467 B.n466 10.6151
R1150 B.n467 B.n194 10.6151
R1151 B.n477 B.n194 10.6151
R1152 B.n478 B.n477 10.6151
R1153 B.n479 B.n478 10.6151
R1154 B.n479 B.n186 10.6151
R1155 B.n489 B.n186 10.6151
R1156 B.n490 B.n489 10.6151
R1157 B.n491 B.n490 10.6151
R1158 B.n491 B.n178 10.6151
R1159 B.n502 B.n178 10.6151
R1160 B.n503 B.n502 10.6151
R1161 B.n504 B.n503 10.6151
R1162 B.n504 B.n0 10.6151
R1163 B.n356 B.n273 10.6151
R1164 B.n351 B.n273 10.6151
R1165 B.n351 B.n350 10.6151
R1166 B.n350 B.n349 10.6151
R1167 B.n349 B.n346 10.6151
R1168 B.n346 B.n345 10.6151
R1169 B.n345 B.n342 10.6151
R1170 B.n342 B.n341 10.6151
R1171 B.n341 B.n338 10.6151
R1172 B.n338 B.n337 10.6151
R1173 B.n334 B.n333 10.6151
R1174 B.n333 B.n330 10.6151
R1175 B.n330 B.n329 10.6151
R1176 B.n329 B.n326 10.6151
R1177 B.n326 B.n325 10.6151
R1178 B.n325 B.n322 10.6151
R1179 B.n322 B.n321 10.6151
R1180 B.n321 B.n318 10.6151
R1181 B.n316 B.n313 10.6151
R1182 B.n313 B.n312 10.6151
R1183 B.n312 B.n309 10.6151
R1184 B.n309 B.n308 10.6151
R1185 B.n308 B.n305 10.6151
R1186 B.n305 B.n304 10.6151
R1187 B.n304 B.n301 10.6151
R1188 B.n301 B.n300 10.6151
R1189 B.n300 B.n297 10.6151
R1190 B.n297 B.n296 10.6151
R1191 B.n362 B.n269 10.6151
R1192 B.n363 B.n362 10.6151
R1193 B.n364 B.n363 10.6151
R1194 B.n364 B.n261 10.6151
R1195 B.n374 B.n261 10.6151
R1196 B.n375 B.n374 10.6151
R1197 B.n376 B.n375 10.6151
R1198 B.n376 B.n253 10.6151
R1199 B.n386 B.n253 10.6151
R1200 B.n387 B.n386 10.6151
R1201 B.n388 B.n387 10.6151
R1202 B.n388 B.n245 10.6151
R1203 B.n398 B.n245 10.6151
R1204 B.n399 B.n398 10.6151
R1205 B.n400 B.n399 10.6151
R1206 B.n400 B.n237 10.6151
R1207 B.n410 B.n237 10.6151
R1208 B.n411 B.n410 10.6151
R1209 B.n412 B.n411 10.6151
R1210 B.n412 B.n229 10.6151
R1211 B.n422 B.n229 10.6151
R1212 B.n423 B.n422 10.6151
R1213 B.n424 B.n423 10.6151
R1214 B.n424 B.n222 10.6151
R1215 B.n435 B.n222 10.6151
R1216 B.n436 B.n435 10.6151
R1217 B.n437 B.n436 10.6151
R1218 B.n437 B.n214 10.6151
R1219 B.n447 B.n214 10.6151
R1220 B.n448 B.n447 10.6151
R1221 B.n449 B.n448 10.6151
R1222 B.n449 B.n206 10.6151
R1223 B.n459 B.n206 10.6151
R1224 B.n460 B.n459 10.6151
R1225 B.n461 B.n460 10.6151
R1226 B.n461 B.n198 10.6151
R1227 B.n471 B.n198 10.6151
R1228 B.n472 B.n471 10.6151
R1229 B.n473 B.n472 10.6151
R1230 B.n473 B.n190 10.6151
R1231 B.n483 B.n190 10.6151
R1232 B.n484 B.n483 10.6151
R1233 B.n485 B.n484 10.6151
R1234 B.n485 B.n181 10.6151
R1235 B.n495 B.n181 10.6151
R1236 B.n496 B.n495 10.6151
R1237 B.n498 B.n496 10.6151
R1238 B.n498 B.n497 10.6151
R1239 B.n497 B.n174 10.6151
R1240 B.n509 B.n174 10.6151
R1241 B.n510 B.n509 10.6151
R1242 B.n511 B.n510 10.6151
R1243 B.n512 B.n511 10.6151
R1244 B.n513 B.n512 10.6151
R1245 B.n516 B.n513 10.6151
R1246 B.n517 B.n516 10.6151
R1247 B.n518 B.n517 10.6151
R1248 B.n519 B.n518 10.6151
R1249 B.n521 B.n519 10.6151
R1250 B.n522 B.n521 10.6151
R1251 B.n523 B.n522 10.6151
R1252 B.n524 B.n523 10.6151
R1253 B.n526 B.n524 10.6151
R1254 B.n527 B.n526 10.6151
R1255 B.n528 B.n527 10.6151
R1256 B.n529 B.n528 10.6151
R1257 B.n531 B.n529 10.6151
R1258 B.n532 B.n531 10.6151
R1259 B.n533 B.n532 10.6151
R1260 B.n534 B.n533 10.6151
R1261 B.n536 B.n534 10.6151
R1262 B.n537 B.n536 10.6151
R1263 B.n538 B.n537 10.6151
R1264 B.n539 B.n538 10.6151
R1265 B.n541 B.n539 10.6151
R1266 B.n542 B.n541 10.6151
R1267 B.n543 B.n542 10.6151
R1268 B.n544 B.n543 10.6151
R1269 B.n546 B.n544 10.6151
R1270 B.n547 B.n546 10.6151
R1271 B.n548 B.n547 10.6151
R1272 B.n549 B.n548 10.6151
R1273 B.n551 B.n549 10.6151
R1274 B.n552 B.n551 10.6151
R1275 B.n553 B.n552 10.6151
R1276 B.n554 B.n553 10.6151
R1277 B.n556 B.n554 10.6151
R1278 B.n557 B.n556 10.6151
R1279 B.n558 B.n557 10.6151
R1280 B.n559 B.n558 10.6151
R1281 B.n561 B.n559 10.6151
R1282 B.n562 B.n561 10.6151
R1283 B.n563 B.n562 10.6151
R1284 B.n564 B.n563 10.6151
R1285 B.n566 B.n564 10.6151
R1286 B.n567 B.n566 10.6151
R1287 B.n568 B.n567 10.6151
R1288 B.n569 B.n568 10.6151
R1289 B.n571 B.n569 10.6151
R1290 B.n572 B.n571 10.6151
R1291 B.n573 B.n572 10.6151
R1292 B.n574 B.n573 10.6151
R1293 B.n575 B.n574 10.6151
R1294 B.n679 B.n1 10.6151
R1295 B.n679 B.n678 10.6151
R1296 B.n678 B.n677 10.6151
R1297 B.n677 B.n10 10.6151
R1298 B.n671 B.n10 10.6151
R1299 B.n671 B.n670 10.6151
R1300 B.n670 B.n669 10.6151
R1301 B.n669 B.n18 10.6151
R1302 B.n663 B.n18 10.6151
R1303 B.n663 B.n662 10.6151
R1304 B.n662 B.n661 10.6151
R1305 B.n661 B.n25 10.6151
R1306 B.n655 B.n25 10.6151
R1307 B.n655 B.n654 10.6151
R1308 B.n654 B.n653 10.6151
R1309 B.n653 B.n32 10.6151
R1310 B.n647 B.n32 10.6151
R1311 B.n647 B.n646 10.6151
R1312 B.n646 B.n645 10.6151
R1313 B.n645 B.n39 10.6151
R1314 B.n639 B.n39 10.6151
R1315 B.n639 B.n638 10.6151
R1316 B.n638 B.n637 10.6151
R1317 B.n637 B.n46 10.6151
R1318 B.n631 B.n46 10.6151
R1319 B.n631 B.n630 10.6151
R1320 B.n630 B.n629 10.6151
R1321 B.n629 B.n52 10.6151
R1322 B.n623 B.n52 10.6151
R1323 B.n623 B.n622 10.6151
R1324 B.n622 B.n621 10.6151
R1325 B.n621 B.n60 10.6151
R1326 B.n615 B.n60 10.6151
R1327 B.n615 B.n614 10.6151
R1328 B.n614 B.n613 10.6151
R1329 B.n613 B.n67 10.6151
R1330 B.n607 B.n67 10.6151
R1331 B.n607 B.n606 10.6151
R1332 B.n606 B.n605 10.6151
R1333 B.n605 B.n74 10.6151
R1334 B.n599 B.n74 10.6151
R1335 B.n599 B.n598 10.6151
R1336 B.n598 B.n597 10.6151
R1337 B.n597 B.n81 10.6151
R1338 B.n591 B.n81 10.6151
R1339 B.n591 B.n590 10.6151
R1340 B.n590 B.n589 10.6151
R1341 B.n589 B.n88 10.6151
R1342 B.n583 B.n88 10.6151
R1343 B.n583 B.n582 10.6151
R1344 B.n581 B.n95 10.6151
R1345 B.n119 B.n95 10.6151
R1346 B.n120 B.n119 10.6151
R1347 B.n123 B.n120 10.6151
R1348 B.n124 B.n123 10.6151
R1349 B.n127 B.n124 10.6151
R1350 B.n128 B.n127 10.6151
R1351 B.n131 B.n128 10.6151
R1352 B.n132 B.n131 10.6151
R1353 B.n135 B.n132 10.6151
R1354 B.n140 B.n137 10.6151
R1355 B.n141 B.n140 10.6151
R1356 B.n144 B.n141 10.6151
R1357 B.n145 B.n144 10.6151
R1358 B.n148 B.n145 10.6151
R1359 B.n149 B.n148 10.6151
R1360 B.n152 B.n149 10.6151
R1361 B.n153 B.n152 10.6151
R1362 B.n157 B.n156 10.6151
R1363 B.n160 B.n157 10.6151
R1364 B.n161 B.n160 10.6151
R1365 B.n164 B.n161 10.6151
R1366 B.n165 B.n164 10.6151
R1367 B.n168 B.n165 10.6151
R1368 B.n169 B.n168 10.6151
R1369 B.n172 B.n169 10.6151
R1370 B.n173 B.n172 10.6151
R1371 B.n576 B.n173 10.6151
R1372 B.n475 B.t5 9.7422
R1373 B.n659 B.t9 9.7422
R1374 B.n687 B.n0 8.11757
R1375 B.n687 B.n1 8.11757
R1376 B.n334 B.n292 6.5566
R1377 B.n318 B.n317 6.5566
R1378 B.n137 B.n136 6.5566
R1379 B.n153 B.n115 6.5566
R1380 B.n378 B.t11 6.49496
R1381 B.n595 B.t18 6.49496
R1382 B.n337 B.n292 4.05904
R1383 B.n317 B.n316 4.05904
R1384 B.n136 B.n135 4.05904
R1385 B.n156 B.n115 4.05904
R1386 VP.n20 VP.n19 161.3
R1387 VP.n21 VP.n16 161.3
R1388 VP.n23 VP.n22 161.3
R1389 VP.n24 VP.n15 161.3
R1390 VP.n26 VP.n25 161.3
R1391 VP.n27 VP.n14 161.3
R1392 VP.n29 VP.n28 161.3
R1393 VP.n30 VP.n13 161.3
R1394 VP.n32 VP.n31 161.3
R1395 VP.n34 VP.n12 161.3
R1396 VP.n36 VP.n35 161.3
R1397 VP.n37 VP.n11 161.3
R1398 VP.n39 VP.n38 161.3
R1399 VP.n40 VP.n10 161.3
R1400 VP.n74 VP.n0 161.3
R1401 VP.n73 VP.n72 161.3
R1402 VP.n71 VP.n1 161.3
R1403 VP.n70 VP.n69 161.3
R1404 VP.n68 VP.n2 161.3
R1405 VP.n66 VP.n65 161.3
R1406 VP.n64 VP.n3 161.3
R1407 VP.n63 VP.n62 161.3
R1408 VP.n61 VP.n4 161.3
R1409 VP.n60 VP.n59 161.3
R1410 VP.n58 VP.n5 161.3
R1411 VP.n57 VP.n56 161.3
R1412 VP.n55 VP.n6 161.3
R1413 VP.n54 VP.n53 161.3
R1414 VP.n52 VP.n51 161.3
R1415 VP.n50 VP.n8 161.3
R1416 VP.n49 VP.n48 161.3
R1417 VP.n47 VP.n9 161.3
R1418 VP.n46 VP.n45 161.3
R1419 VP.n44 VP.n43 91.2348
R1420 VP.n76 VP.n75 91.2348
R1421 VP.n42 VP.n41 91.2348
R1422 VP.n49 VP.n9 56.5617
R1423 VP.n56 VP.n55 56.5617
R1424 VP.n62 VP.n3 56.5617
R1425 VP.n73 VP.n1 56.5617
R1426 VP.n39 VP.n11 56.5617
R1427 VP.n28 VP.n13 56.5617
R1428 VP.n22 VP.n21 56.5617
R1429 VP.n18 VP.t7 51.2161
R1430 VP.n18 VP.n17 48.5947
R1431 VP.n43 VP.n42 42.6019
R1432 VP.n45 VP.n9 24.5923
R1433 VP.n50 VP.n49 24.5923
R1434 VP.n51 VP.n50 24.5923
R1435 VP.n55 VP.n54 24.5923
R1436 VP.n56 VP.n5 24.5923
R1437 VP.n60 VP.n5 24.5923
R1438 VP.n61 VP.n60 24.5923
R1439 VP.n62 VP.n61 24.5923
R1440 VP.n66 VP.n3 24.5923
R1441 VP.n69 VP.n68 24.5923
R1442 VP.n69 VP.n1 24.5923
R1443 VP.n74 VP.n73 24.5923
R1444 VP.n40 VP.n39 24.5923
R1445 VP.n32 VP.n13 24.5923
R1446 VP.n35 VP.n34 24.5923
R1447 VP.n35 VP.n11 24.5923
R1448 VP.n22 VP.n15 24.5923
R1449 VP.n26 VP.n15 24.5923
R1450 VP.n27 VP.n26 24.5923
R1451 VP.n28 VP.n27 24.5923
R1452 VP.n21 VP.n20 24.5923
R1453 VP.n54 VP.n7 22.1332
R1454 VP.n67 VP.n66 22.1332
R1455 VP.n33 VP.n32 22.1332
R1456 VP.n20 VP.n17 22.1332
R1457 VP.n45 VP.n44 19.674
R1458 VP.n75 VP.n74 19.674
R1459 VP.n41 VP.n40 19.674
R1460 VP.n60 VP.t4 17.0524
R1461 VP.n44 VP.t8 17.0524
R1462 VP.n7 VP.t5 17.0524
R1463 VP.n67 VP.t3 17.0524
R1464 VP.n75 VP.t2 17.0524
R1465 VP.n26 VP.t9 17.0524
R1466 VP.n41 VP.t1 17.0524
R1467 VP.n33 VP.t6 17.0524
R1468 VP.n17 VP.t0 17.0524
R1469 VP.n19 VP.n18 8.9882
R1470 VP.n51 VP.n7 2.45968
R1471 VP.n68 VP.n67 2.45968
R1472 VP.n34 VP.n33 2.45968
R1473 VP.n42 VP.n10 0.278335
R1474 VP.n46 VP.n43 0.278335
R1475 VP.n76 VP.n0 0.278335
R1476 VP.n19 VP.n16 0.189894
R1477 VP.n23 VP.n16 0.189894
R1478 VP.n24 VP.n23 0.189894
R1479 VP.n25 VP.n24 0.189894
R1480 VP.n25 VP.n14 0.189894
R1481 VP.n29 VP.n14 0.189894
R1482 VP.n30 VP.n29 0.189894
R1483 VP.n31 VP.n30 0.189894
R1484 VP.n31 VP.n12 0.189894
R1485 VP.n36 VP.n12 0.189894
R1486 VP.n37 VP.n36 0.189894
R1487 VP.n38 VP.n37 0.189894
R1488 VP.n38 VP.n10 0.189894
R1489 VP.n47 VP.n46 0.189894
R1490 VP.n48 VP.n47 0.189894
R1491 VP.n48 VP.n8 0.189894
R1492 VP.n52 VP.n8 0.189894
R1493 VP.n53 VP.n52 0.189894
R1494 VP.n53 VP.n6 0.189894
R1495 VP.n57 VP.n6 0.189894
R1496 VP.n58 VP.n57 0.189894
R1497 VP.n59 VP.n58 0.189894
R1498 VP.n59 VP.n4 0.189894
R1499 VP.n63 VP.n4 0.189894
R1500 VP.n64 VP.n63 0.189894
R1501 VP.n65 VP.n64 0.189894
R1502 VP.n65 VP.n2 0.189894
R1503 VP.n70 VP.n2 0.189894
R1504 VP.n71 VP.n70 0.189894
R1505 VP.n72 VP.n71 0.189894
R1506 VP.n72 VP.n0 0.189894
R1507 VP VP.n76 0.153485
R1508 VDD1.n1 VDD1.t2 132.876
R1509 VDD1.n3 VDD1.t1 132.876
R1510 VDD1.n5 VDD1.n4 119.093
R1511 VDD1.n1 VDD1.n0 117.564
R1512 VDD1.n7 VDD1.n6 117.564
R1513 VDD1.n3 VDD1.n2 117.564
R1514 VDD1.n7 VDD1.n5 36.6798
R1515 VDD1.n6 VDD1.t3 13.2005
R1516 VDD1.n6 VDD1.t8 13.2005
R1517 VDD1.n0 VDD1.t9 13.2005
R1518 VDD1.n0 VDD1.t0 13.2005
R1519 VDD1.n4 VDD1.t6 13.2005
R1520 VDD1.n4 VDD1.t7 13.2005
R1521 VDD1.n2 VDD1.t4 13.2005
R1522 VDD1.n2 VDD1.t5 13.2005
R1523 VDD1 VDD1.n7 1.52636
R1524 VDD1 VDD1.n1 0.586707
R1525 VDD1.n5 VDD1.n3 0.473171
C0 VTAIL VN 2.92279f
C1 VDD2 VP 0.530655f
C2 VN VDD1 0.159996f
C3 VTAIL VDD2 5.07393f
C4 VDD2 VDD1 1.86169f
C5 VDD2 VN 1.71436f
C6 VTAIL VP 2.93693f
C7 VP VDD1 2.0814f
C8 VTAIL VDD1 5.02386f
C9 VN VP 5.74874f
C10 VDD2 B 4.595554f
C11 VDD1 B 4.742323f
C12 VTAIL B 3.236315f
C13 VN B 14.740919f
C14 VP B 13.383558f
C15 VDD1.t2 B 0.231487f
C16 VDD1.t9 B 0.028772f
C17 VDD1.t0 B 0.028772f
C18 VDD1.n0 B 0.169355f
C19 VDD1.n1 B 0.734714f
C20 VDD1.t1 B 0.231486f
C21 VDD1.t4 B 0.028772f
C22 VDD1.t5 B 0.028772f
C23 VDD1.n2 B 0.169355f
C24 VDD1.n3 B 0.727025f
C25 VDD1.t6 B 0.028772f
C26 VDD1.t7 B 0.028772f
C27 VDD1.n4 B 0.175274f
C28 VDD1.n5 B 2.04185f
C29 VDD1.t3 B 0.028772f
C30 VDD1.t8 B 0.028772f
C31 VDD1.n6 B 0.169355f
C32 VDD1.n7 B 2.05473f
C33 VP.n0 B 0.045472f
C34 VP.t2 B 0.239083f
C35 VP.n1 B 0.042983f
C36 VP.n2 B 0.034493f
C37 VP.t3 B 0.239083f
C38 VP.n3 B 0.052526f
C39 VP.n4 B 0.034493f
C40 VP.t4 B 0.239083f
C41 VP.n5 B 0.063963f
C42 VP.n6 B 0.034493f
C43 VP.t5 B 0.239083f
C44 VP.n7 B 0.134041f
C45 VP.n8 B 0.034493f
C46 VP.n9 B 0.057298f
C47 VP.n10 B 0.045472f
C48 VP.t1 B 0.239083f
C49 VP.n11 B 0.042983f
C50 VP.n12 B 0.034493f
C51 VP.t6 B 0.239083f
C52 VP.n13 B 0.052526f
C53 VP.n14 B 0.034493f
C54 VP.t9 B 0.239083f
C55 VP.n15 B 0.063963f
C56 VP.n16 B 0.034493f
C57 VP.t0 B 0.239083f
C58 VP.n17 B 0.23338f
C59 VP.t7 B 0.452597f
C60 VP.n18 B 0.201743f
C61 VP.n19 B 0.290946f
C62 VP.n20 B 0.060806f
C63 VP.n21 B 0.052526f
C64 VP.n22 B 0.047755f
C65 VP.n23 B 0.034493f
C66 VP.n24 B 0.034493f
C67 VP.n25 B 0.034493f
C68 VP.n26 B 0.166428f
C69 VP.n27 B 0.063963f
C70 VP.n28 B 0.047755f
C71 VP.n29 B 0.034493f
C72 VP.n30 B 0.034493f
C73 VP.n31 B 0.034493f
C74 VP.n32 B 0.060806f
C75 VP.n33 B 0.134041f
C76 VP.n34 B 0.035544f
C77 VP.n35 B 0.063963f
C78 VP.n36 B 0.034493f
C79 VP.n37 B 0.034493f
C80 VP.n38 B 0.034493f
C81 VP.n39 B 0.057298f
C82 VP.n40 B 0.057648f
C83 VP.n41 B 0.244941f
C84 VP.n42 B 1.48808f
C85 VP.n43 B 1.51726f
C86 VP.t8 B 0.239083f
C87 VP.n44 B 0.244941f
C88 VP.n45 B 0.057648f
C89 VP.n46 B 0.045472f
C90 VP.n47 B 0.034493f
C91 VP.n48 B 0.034493f
C92 VP.n49 B 0.042983f
C93 VP.n50 B 0.063963f
C94 VP.n51 B 0.035544f
C95 VP.n52 B 0.034493f
C96 VP.n53 B 0.034493f
C97 VP.n54 B 0.060806f
C98 VP.n55 B 0.052526f
C99 VP.n56 B 0.047755f
C100 VP.n57 B 0.034493f
C101 VP.n58 B 0.034493f
C102 VP.n59 B 0.034493f
C103 VP.n60 B 0.166428f
C104 VP.n61 B 0.063963f
C105 VP.n62 B 0.047755f
C106 VP.n63 B 0.034493f
C107 VP.n64 B 0.034493f
C108 VP.n65 B 0.034493f
C109 VP.n66 B 0.060806f
C110 VP.n67 B 0.134041f
C111 VP.n68 B 0.035544f
C112 VP.n69 B 0.063963f
C113 VP.n70 B 0.034493f
C114 VP.n71 B 0.034493f
C115 VP.n72 B 0.034493f
C116 VP.n73 B 0.057298f
C117 VP.n74 B 0.057648f
C118 VP.n75 B 0.244941f
C119 VP.n76 B 0.042768f
C120 VDD2.t2 B 0.168405f
C121 VDD2.t1 B 0.020932f
C122 VDD2.t9 B 0.020932f
C123 VDD2.n0 B 0.123205f
C124 VDD2.n1 B 0.528908f
C125 VDD2.t6 B 0.020932f
C126 VDD2.t4 B 0.020932f
C127 VDD2.n2 B 0.127511f
C128 VDD2.n3 B 1.4125f
C129 VDD2.t5 B 0.164205f
C130 VDD2.n4 B 1.43178f
C131 VDD2.t0 B 0.020932f
C132 VDD2.t8 B 0.020932f
C133 VDD2.n5 B 0.123205f
C134 VDD2.n6 B 0.274429f
C135 VDD2.t7 B 0.020932f
C136 VDD2.t3 B 0.020932f
C137 VDD2.n7 B 0.127497f
C138 VTAIL.t19 B 0.044676f
C139 VTAIL.t13 B 0.044676f
C140 VTAIL.n0 B 0.221493f
C141 VTAIL.n1 B 0.633043f
C142 VTAIL.t6 B 0.308782f
C143 VTAIL.n2 B 0.724658f
C144 VTAIL.t2 B 0.044676f
C145 VTAIL.t5 B 0.044676f
C146 VTAIL.n3 B 0.221493f
C147 VTAIL.n4 B 0.761295f
C148 VTAIL.t1 B 0.044676f
C149 VTAIL.t4 B 0.044676f
C150 VTAIL.n5 B 0.221493f
C151 VTAIL.n6 B 1.68683f
C152 VTAIL.t18 B 0.044676f
C153 VTAIL.t14 B 0.044676f
C154 VTAIL.n7 B 0.221494f
C155 VTAIL.n8 B 1.68683f
C156 VTAIL.t12 B 0.044676f
C157 VTAIL.t15 B 0.044676f
C158 VTAIL.n9 B 0.221494f
C159 VTAIL.n10 B 0.761295f
C160 VTAIL.t17 B 0.308782f
C161 VTAIL.n11 B 0.724658f
C162 VTAIL.t8 B 0.044676f
C163 VTAIL.t9 B 0.044676f
C164 VTAIL.n12 B 0.221494f
C165 VTAIL.n13 B 0.690101f
C166 VTAIL.t0 B 0.044676f
C167 VTAIL.t3 B 0.044676f
C168 VTAIL.n14 B 0.221494f
C169 VTAIL.n15 B 0.761295f
C170 VTAIL.t7 B 0.308782f
C171 VTAIL.n16 B 1.46488f
C172 VTAIL.t16 B 0.308782f
C173 VTAIL.n17 B 1.46488f
C174 VTAIL.t11 B 0.044676f
C175 VTAIL.t10 B 0.044676f
C176 VTAIL.n18 B 0.221493f
C177 VTAIL.n19 B 0.561849f
C178 VN.n0 B 0.036383f
C179 VN.t5 B 0.191294f
C180 VN.n1 B 0.034391f
C181 VN.n2 B 0.027598f
C182 VN.t3 B 0.191294f
C183 VN.n3 B 0.042027f
C184 VN.n4 B 0.027598f
C185 VN.t0 B 0.191294f
C186 VN.n5 B 0.051178f
C187 VN.n6 B 0.027598f
C188 VN.t8 B 0.191294f
C189 VN.n7 B 0.18673f
C190 VN.t7 B 0.362128f
C191 VN.n8 B 0.161417f
C192 VN.n9 B 0.232789f
C193 VN.n10 B 0.048651f
C194 VN.n11 B 0.042027f
C195 VN.n12 B 0.038209f
C196 VN.n13 B 0.027598f
C197 VN.n14 B 0.027598f
C198 VN.n15 B 0.027598f
C199 VN.n16 B 0.133161f
C200 VN.n17 B 0.051178f
C201 VN.n18 B 0.038209f
C202 VN.n19 B 0.027598f
C203 VN.n20 B 0.027598f
C204 VN.n21 B 0.027598f
C205 VN.n22 B 0.048651f
C206 VN.n23 B 0.107248f
C207 VN.n24 B 0.028439f
C208 VN.n25 B 0.051178f
C209 VN.n26 B 0.027598f
C210 VN.n27 B 0.027598f
C211 VN.n28 B 0.027598f
C212 VN.n29 B 0.045845f
C213 VN.n30 B 0.046125f
C214 VN.n31 B 0.195981f
C215 VN.n32 B 0.034219f
C216 VN.n33 B 0.036383f
C217 VN.t4 B 0.191294f
C218 VN.n34 B 0.034391f
C219 VN.n35 B 0.027598f
C220 VN.t9 B 0.191294f
C221 VN.n36 B 0.042027f
C222 VN.n37 B 0.027598f
C223 VN.t1 B 0.191294f
C224 VN.n38 B 0.051178f
C225 VN.n39 B 0.027598f
C226 VN.t2 B 0.191294f
C227 VN.n40 B 0.18673f
C228 VN.t6 B 0.362128f
C229 VN.n41 B 0.161417f
C230 VN.n42 B 0.232789f
C231 VN.n43 B 0.048651f
C232 VN.n44 B 0.042027f
C233 VN.n45 B 0.038209f
C234 VN.n46 B 0.027598f
C235 VN.n47 B 0.027598f
C236 VN.n48 B 0.027598f
C237 VN.n49 B 0.133161f
C238 VN.n50 B 0.051178f
C239 VN.n51 B 0.038209f
C240 VN.n52 B 0.027598f
C241 VN.n53 B 0.027598f
C242 VN.n54 B 0.027598f
C243 VN.n55 B 0.048651f
C244 VN.n56 B 0.107248f
C245 VN.n57 B 0.028439f
C246 VN.n58 B 0.051178f
C247 VN.n59 B 0.027598f
C248 VN.n60 B 0.027598f
C249 VN.n61 B 0.027598f
C250 VN.n62 B 0.045845f
C251 VN.n63 B 0.046125f
C252 VN.n64 B 0.195981f
C253 VN.n65 B 1.20586f
.ends

