* NGSPICE file created from diff_pair_sample_0102.ext - technology: sky130A

.subckt diff_pair_sample_0102 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=6.9186 ps=36.26 w=17.74 l=3.41
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=0 ps=0 w=17.74 l=3.41
X2 VDD1.t4 VP.t1 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=2.9271 ps=18.07 w=17.74 l=3.41
X3 VTAIL.t5 VN.t0 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=2.9271 ps=18.07 w=17.74 l=3.41
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=0 ps=0 w=17.74 l=3.41
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=0 ps=0 w=17.74 l=3.41
X6 VTAIL.t10 VP.t2 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=2.9271 ps=18.07 w=17.74 l=3.41
X7 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=2.9271 ps=18.07 w=17.74 l=3.41
X8 VDD2.t3 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=6.9186 ps=36.26 w=17.74 l=3.41
X9 VDD2.t2 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=2.9271 ps=18.07 w=17.74 l=3.41
X10 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=6.9186 ps=36.26 w=17.74 l=3.41
X11 VDD1.t2 VP.t3 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=6.9186 ps=36.26 w=17.74 l=3.41
X12 VTAIL.t9 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=2.9271 ps=18.07 w=17.74 l=3.41
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=0 ps=0 w=17.74 l=3.41
X14 VTAIL.t4 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9271 pd=18.07 as=2.9271 ps=18.07 w=17.74 l=3.41
X15 VDD1.t0 VP.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=6.9186 pd=36.26 as=2.9271 ps=18.07 w=17.74 l=3.41
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n50 VP.n49 161.3
R8 VP.n48 VP.n1 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n2 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n42 VP.n3 161.3
R13 VP.n41 VP.n40 161.3
R14 VP.n39 VP.n4 161.3
R15 VP.n38 VP.n37 161.3
R16 VP.n36 VP.n5 161.3
R17 VP.n35 VP.n34 161.3
R18 VP.n33 VP.n6 161.3
R19 VP.n32 VP.n31 161.3
R20 VP.n30 VP.n7 161.3
R21 VP.n29 VP.n28 161.3
R22 VP.n14 VP.t1 159.168
R23 VP.n4 VP.t4 125.377
R24 VP.n8 VP.t5 125.377
R25 VP.n0 VP.t0 125.377
R26 VP.n13 VP.t2 125.377
R27 VP.n9 VP.t3 125.377
R28 VP.n27 VP.n8 78.4415
R29 VP.n51 VP.n0 78.4415
R30 VP.n26 VP.n9 78.4415
R31 VP.n27 VP.n26 56.295
R32 VP.n35 VP.n6 53.171
R33 VP.n43 VP.n2 53.171
R34 VP.n18 VP.n11 53.171
R35 VP.n14 VP.n13 50.2542
R36 VP.n31 VP.n6 27.983
R37 VP.n47 VP.n2 27.983
R38 VP.n22 VP.n11 27.983
R39 VP.n30 VP.n29 24.5923
R40 VP.n31 VP.n30 24.5923
R41 VP.n36 VP.n35 24.5923
R42 VP.n37 VP.n36 24.5923
R43 VP.n37 VP.n4 24.5923
R44 VP.n41 VP.n4 24.5923
R45 VP.n42 VP.n41 24.5923
R46 VP.n43 VP.n42 24.5923
R47 VP.n48 VP.n47 24.5923
R48 VP.n49 VP.n48 24.5923
R49 VP.n23 VP.n22 24.5923
R50 VP.n24 VP.n23 24.5923
R51 VP.n16 VP.n13 24.5923
R52 VP.n17 VP.n16 24.5923
R53 VP.n18 VP.n17 24.5923
R54 VP.n29 VP.n8 11.8046
R55 VP.n49 VP.n0 11.8046
R56 VP.n24 VP.n9 11.8046
R57 VP.n15 VP.n14 3.08084
R58 VP.n26 VP.n25 0.354861
R59 VP.n28 VP.n27 0.354861
R60 VP.n51 VP.n50 0.354861
R61 VP VP.n51 0.267071
R62 VP.n15 VP.n12 0.189894
R63 VP.n19 VP.n12 0.189894
R64 VP.n20 VP.n19 0.189894
R65 VP.n21 VP.n20 0.189894
R66 VP.n21 VP.n10 0.189894
R67 VP.n25 VP.n10 0.189894
R68 VP.n28 VP.n7 0.189894
R69 VP.n32 VP.n7 0.189894
R70 VP.n33 VP.n32 0.189894
R71 VP.n34 VP.n33 0.189894
R72 VP.n34 VP.n5 0.189894
R73 VP.n38 VP.n5 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n40 VP.n39 0.189894
R76 VP.n40 VP.n3 0.189894
R77 VP.n44 VP.n3 0.189894
R78 VP.n45 VP.n44 0.189894
R79 VP.n46 VP.n45 0.189894
R80 VP.n46 VP.n1 0.189894
R81 VP.n50 VP.n1 0.189894
R82 VTAIL.n7 VTAIL.t0 48.7801
R83 VTAIL.n11 VTAIL.t1 48.7791
R84 VTAIL.n2 VTAIL.t8 48.7791
R85 VTAIL.n10 VTAIL.t7 48.7791
R86 VTAIL.n9 VTAIL.n8 47.664
R87 VTAIL.n6 VTAIL.n5 47.664
R88 VTAIL.n1 VTAIL.n0 47.663
R89 VTAIL.n4 VTAIL.n3 47.663
R90 VTAIL.n6 VTAIL.n4 34.1083
R91 VTAIL.n11 VTAIL.n10 30.8841
R92 VTAIL.n7 VTAIL.n6 3.22464
R93 VTAIL.n10 VTAIL.n9 3.22464
R94 VTAIL.n4 VTAIL.n2 3.22464
R95 VTAIL VTAIL.n11 2.36041
R96 VTAIL.n9 VTAIL.n7 2.0824
R97 VTAIL.n2 VTAIL.n1 2.0824
R98 VTAIL.n0 VTAIL.t3 1.11662
R99 VTAIL.n0 VTAIL.t5 1.11662
R100 VTAIL.n3 VTAIL.t6 1.11662
R101 VTAIL.n3 VTAIL.t9 1.11662
R102 VTAIL.n8 VTAIL.t11 1.11662
R103 VTAIL.n8 VTAIL.t10 1.11662
R104 VTAIL.n5 VTAIL.t2 1.11662
R105 VTAIL.n5 VTAIL.t4 1.11662
R106 VTAIL VTAIL.n1 0.864724
R107 VDD1 VDD1.t4 67.9352
R108 VDD1.n1 VDD1.t0 67.8207
R109 VDD1.n1 VDD1.n0 65.0924
R110 VDD1.n3 VDD1.n2 64.3418
R111 VDD1.n3 VDD1.n1 51.6819
R112 VDD1.n2 VDD1.t3 1.11662
R113 VDD1.n2 VDD1.t2 1.11662
R114 VDD1.n0 VDD1.t1 1.11662
R115 VDD1.n0 VDD1.t5 1.11662
R116 VDD1 VDD1.n3 0.748345
R117 B.n1064 B.n1063 585
R118 B.n1065 B.n1064 585
R119 B.n415 B.n160 585
R120 B.n414 B.n413 585
R121 B.n412 B.n411 585
R122 B.n410 B.n409 585
R123 B.n408 B.n407 585
R124 B.n406 B.n405 585
R125 B.n404 B.n403 585
R126 B.n402 B.n401 585
R127 B.n400 B.n399 585
R128 B.n398 B.n397 585
R129 B.n396 B.n395 585
R130 B.n394 B.n393 585
R131 B.n392 B.n391 585
R132 B.n390 B.n389 585
R133 B.n388 B.n387 585
R134 B.n386 B.n385 585
R135 B.n384 B.n383 585
R136 B.n382 B.n381 585
R137 B.n380 B.n379 585
R138 B.n378 B.n377 585
R139 B.n376 B.n375 585
R140 B.n374 B.n373 585
R141 B.n372 B.n371 585
R142 B.n370 B.n369 585
R143 B.n368 B.n367 585
R144 B.n366 B.n365 585
R145 B.n364 B.n363 585
R146 B.n362 B.n361 585
R147 B.n360 B.n359 585
R148 B.n358 B.n357 585
R149 B.n356 B.n355 585
R150 B.n354 B.n353 585
R151 B.n352 B.n351 585
R152 B.n350 B.n349 585
R153 B.n348 B.n347 585
R154 B.n346 B.n345 585
R155 B.n344 B.n343 585
R156 B.n342 B.n341 585
R157 B.n340 B.n339 585
R158 B.n338 B.n337 585
R159 B.n336 B.n335 585
R160 B.n334 B.n333 585
R161 B.n332 B.n331 585
R162 B.n330 B.n329 585
R163 B.n328 B.n327 585
R164 B.n326 B.n325 585
R165 B.n324 B.n323 585
R166 B.n322 B.n321 585
R167 B.n320 B.n319 585
R168 B.n318 B.n317 585
R169 B.n316 B.n315 585
R170 B.n314 B.n313 585
R171 B.n312 B.n311 585
R172 B.n310 B.n309 585
R173 B.n308 B.n307 585
R174 B.n306 B.n305 585
R175 B.n304 B.n303 585
R176 B.n302 B.n301 585
R177 B.n300 B.n299 585
R178 B.n298 B.n297 585
R179 B.n296 B.n295 585
R180 B.n294 B.n293 585
R181 B.n292 B.n291 585
R182 B.n290 B.n289 585
R183 B.n288 B.n287 585
R184 B.n286 B.n285 585
R185 B.n284 B.n283 585
R186 B.n281 B.n280 585
R187 B.n279 B.n278 585
R188 B.n277 B.n276 585
R189 B.n275 B.n274 585
R190 B.n273 B.n272 585
R191 B.n271 B.n270 585
R192 B.n269 B.n268 585
R193 B.n267 B.n266 585
R194 B.n265 B.n264 585
R195 B.n263 B.n262 585
R196 B.n261 B.n260 585
R197 B.n259 B.n258 585
R198 B.n257 B.n256 585
R199 B.n255 B.n254 585
R200 B.n253 B.n252 585
R201 B.n251 B.n250 585
R202 B.n249 B.n248 585
R203 B.n247 B.n246 585
R204 B.n245 B.n244 585
R205 B.n243 B.n242 585
R206 B.n241 B.n240 585
R207 B.n239 B.n238 585
R208 B.n237 B.n236 585
R209 B.n235 B.n234 585
R210 B.n233 B.n232 585
R211 B.n231 B.n230 585
R212 B.n229 B.n228 585
R213 B.n227 B.n226 585
R214 B.n225 B.n224 585
R215 B.n223 B.n222 585
R216 B.n221 B.n220 585
R217 B.n219 B.n218 585
R218 B.n217 B.n216 585
R219 B.n215 B.n214 585
R220 B.n213 B.n212 585
R221 B.n211 B.n210 585
R222 B.n209 B.n208 585
R223 B.n207 B.n206 585
R224 B.n205 B.n204 585
R225 B.n203 B.n202 585
R226 B.n201 B.n200 585
R227 B.n199 B.n198 585
R228 B.n197 B.n196 585
R229 B.n195 B.n194 585
R230 B.n193 B.n192 585
R231 B.n191 B.n190 585
R232 B.n189 B.n188 585
R233 B.n187 B.n186 585
R234 B.n185 B.n184 585
R235 B.n183 B.n182 585
R236 B.n181 B.n180 585
R237 B.n179 B.n178 585
R238 B.n177 B.n176 585
R239 B.n175 B.n174 585
R240 B.n173 B.n172 585
R241 B.n171 B.n170 585
R242 B.n169 B.n168 585
R243 B.n167 B.n166 585
R244 B.n95 B.n94 585
R245 B.n1062 B.n96 585
R246 B.n1066 B.n96 585
R247 B.n1061 B.n1060 585
R248 B.n1060 B.n92 585
R249 B.n1059 B.n91 585
R250 B.n1072 B.n91 585
R251 B.n1058 B.n90 585
R252 B.n1073 B.n90 585
R253 B.n1057 B.n89 585
R254 B.n1074 B.n89 585
R255 B.n1056 B.n1055 585
R256 B.n1055 B.n85 585
R257 B.n1054 B.n84 585
R258 B.n1080 B.n84 585
R259 B.n1053 B.n83 585
R260 B.n1081 B.n83 585
R261 B.n1052 B.n82 585
R262 B.n1082 B.n82 585
R263 B.n1051 B.n1050 585
R264 B.n1050 B.n78 585
R265 B.n1049 B.n77 585
R266 B.n1088 B.n77 585
R267 B.n1048 B.n76 585
R268 B.n1089 B.n76 585
R269 B.n1047 B.n75 585
R270 B.n1090 B.n75 585
R271 B.n1046 B.n1045 585
R272 B.n1045 B.n71 585
R273 B.n1044 B.n70 585
R274 B.n1096 B.n70 585
R275 B.n1043 B.n69 585
R276 B.n1097 B.n69 585
R277 B.n1042 B.n68 585
R278 B.n1098 B.n68 585
R279 B.n1041 B.n1040 585
R280 B.n1040 B.n64 585
R281 B.n1039 B.n63 585
R282 B.n1104 B.n63 585
R283 B.n1038 B.n62 585
R284 B.n1105 B.n62 585
R285 B.n1037 B.n61 585
R286 B.n1106 B.n61 585
R287 B.n1036 B.n1035 585
R288 B.n1035 B.n57 585
R289 B.n1034 B.n56 585
R290 B.n1112 B.n56 585
R291 B.n1033 B.n55 585
R292 B.n1113 B.n55 585
R293 B.n1032 B.n54 585
R294 B.n1114 B.n54 585
R295 B.n1031 B.n1030 585
R296 B.n1030 B.n50 585
R297 B.n1029 B.n49 585
R298 B.n1120 B.n49 585
R299 B.n1028 B.n48 585
R300 B.n1121 B.n48 585
R301 B.n1027 B.n47 585
R302 B.n1122 B.n47 585
R303 B.n1026 B.n1025 585
R304 B.n1025 B.n43 585
R305 B.n1024 B.n42 585
R306 B.n1128 B.n42 585
R307 B.n1023 B.n41 585
R308 B.n1129 B.n41 585
R309 B.n1022 B.n40 585
R310 B.n1130 B.n40 585
R311 B.n1021 B.n1020 585
R312 B.n1020 B.n39 585
R313 B.n1019 B.n35 585
R314 B.n1136 B.n35 585
R315 B.n1018 B.n34 585
R316 B.n1137 B.n34 585
R317 B.n1017 B.n33 585
R318 B.n1138 B.n33 585
R319 B.n1016 B.n1015 585
R320 B.n1015 B.n29 585
R321 B.n1014 B.n28 585
R322 B.n1144 B.n28 585
R323 B.n1013 B.n27 585
R324 B.n1145 B.n27 585
R325 B.n1012 B.n26 585
R326 B.n1146 B.n26 585
R327 B.n1011 B.n1010 585
R328 B.n1010 B.n22 585
R329 B.n1009 B.n21 585
R330 B.n1152 B.n21 585
R331 B.n1008 B.n20 585
R332 B.n1153 B.n20 585
R333 B.n1007 B.n19 585
R334 B.n1154 B.n19 585
R335 B.n1006 B.n1005 585
R336 B.n1005 B.n15 585
R337 B.n1004 B.n14 585
R338 B.n1160 B.n14 585
R339 B.n1003 B.n13 585
R340 B.n1161 B.n13 585
R341 B.n1002 B.n12 585
R342 B.n1162 B.n12 585
R343 B.n1001 B.n1000 585
R344 B.n1000 B.n8 585
R345 B.n999 B.n7 585
R346 B.n1168 B.n7 585
R347 B.n998 B.n6 585
R348 B.n1169 B.n6 585
R349 B.n997 B.n5 585
R350 B.n1170 B.n5 585
R351 B.n996 B.n995 585
R352 B.n995 B.n4 585
R353 B.n994 B.n416 585
R354 B.n994 B.n993 585
R355 B.n984 B.n417 585
R356 B.n418 B.n417 585
R357 B.n986 B.n985 585
R358 B.n987 B.n986 585
R359 B.n983 B.n423 585
R360 B.n423 B.n422 585
R361 B.n982 B.n981 585
R362 B.n981 B.n980 585
R363 B.n425 B.n424 585
R364 B.n426 B.n425 585
R365 B.n973 B.n972 585
R366 B.n974 B.n973 585
R367 B.n971 B.n431 585
R368 B.n431 B.n430 585
R369 B.n970 B.n969 585
R370 B.n969 B.n968 585
R371 B.n433 B.n432 585
R372 B.n434 B.n433 585
R373 B.n961 B.n960 585
R374 B.n962 B.n961 585
R375 B.n959 B.n439 585
R376 B.n439 B.n438 585
R377 B.n958 B.n957 585
R378 B.n957 B.n956 585
R379 B.n441 B.n440 585
R380 B.n442 B.n441 585
R381 B.n949 B.n948 585
R382 B.n950 B.n949 585
R383 B.n947 B.n447 585
R384 B.n447 B.n446 585
R385 B.n946 B.n945 585
R386 B.n945 B.n944 585
R387 B.n449 B.n448 585
R388 B.n937 B.n449 585
R389 B.n936 B.n935 585
R390 B.n938 B.n936 585
R391 B.n934 B.n454 585
R392 B.n454 B.n453 585
R393 B.n933 B.n932 585
R394 B.n932 B.n931 585
R395 B.n456 B.n455 585
R396 B.n457 B.n456 585
R397 B.n924 B.n923 585
R398 B.n925 B.n924 585
R399 B.n922 B.n462 585
R400 B.n462 B.n461 585
R401 B.n921 B.n920 585
R402 B.n920 B.n919 585
R403 B.n464 B.n463 585
R404 B.n465 B.n464 585
R405 B.n912 B.n911 585
R406 B.n913 B.n912 585
R407 B.n910 B.n470 585
R408 B.n470 B.n469 585
R409 B.n909 B.n908 585
R410 B.n908 B.n907 585
R411 B.n472 B.n471 585
R412 B.n473 B.n472 585
R413 B.n900 B.n899 585
R414 B.n901 B.n900 585
R415 B.n898 B.n478 585
R416 B.n478 B.n477 585
R417 B.n897 B.n896 585
R418 B.n896 B.n895 585
R419 B.n480 B.n479 585
R420 B.n481 B.n480 585
R421 B.n888 B.n887 585
R422 B.n889 B.n888 585
R423 B.n886 B.n486 585
R424 B.n486 B.n485 585
R425 B.n885 B.n884 585
R426 B.n884 B.n883 585
R427 B.n488 B.n487 585
R428 B.n489 B.n488 585
R429 B.n876 B.n875 585
R430 B.n877 B.n876 585
R431 B.n874 B.n494 585
R432 B.n494 B.n493 585
R433 B.n873 B.n872 585
R434 B.n872 B.n871 585
R435 B.n496 B.n495 585
R436 B.n497 B.n496 585
R437 B.n864 B.n863 585
R438 B.n865 B.n864 585
R439 B.n862 B.n502 585
R440 B.n502 B.n501 585
R441 B.n861 B.n860 585
R442 B.n860 B.n859 585
R443 B.n504 B.n503 585
R444 B.n505 B.n504 585
R445 B.n852 B.n851 585
R446 B.n853 B.n852 585
R447 B.n850 B.n510 585
R448 B.n510 B.n509 585
R449 B.n849 B.n848 585
R450 B.n848 B.n847 585
R451 B.n512 B.n511 585
R452 B.n513 B.n512 585
R453 B.n840 B.n839 585
R454 B.n841 B.n840 585
R455 B.n516 B.n515 585
R456 B.n585 B.n584 585
R457 B.n586 B.n582 585
R458 B.n582 B.n517 585
R459 B.n588 B.n587 585
R460 B.n590 B.n581 585
R461 B.n593 B.n592 585
R462 B.n594 B.n580 585
R463 B.n596 B.n595 585
R464 B.n598 B.n579 585
R465 B.n601 B.n600 585
R466 B.n602 B.n578 585
R467 B.n604 B.n603 585
R468 B.n606 B.n577 585
R469 B.n609 B.n608 585
R470 B.n610 B.n576 585
R471 B.n612 B.n611 585
R472 B.n614 B.n575 585
R473 B.n617 B.n616 585
R474 B.n618 B.n574 585
R475 B.n620 B.n619 585
R476 B.n622 B.n573 585
R477 B.n625 B.n624 585
R478 B.n626 B.n572 585
R479 B.n628 B.n627 585
R480 B.n630 B.n571 585
R481 B.n633 B.n632 585
R482 B.n634 B.n570 585
R483 B.n636 B.n635 585
R484 B.n638 B.n569 585
R485 B.n641 B.n640 585
R486 B.n642 B.n568 585
R487 B.n644 B.n643 585
R488 B.n646 B.n567 585
R489 B.n649 B.n648 585
R490 B.n650 B.n566 585
R491 B.n652 B.n651 585
R492 B.n654 B.n565 585
R493 B.n657 B.n656 585
R494 B.n658 B.n564 585
R495 B.n660 B.n659 585
R496 B.n662 B.n563 585
R497 B.n665 B.n664 585
R498 B.n666 B.n562 585
R499 B.n668 B.n667 585
R500 B.n670 B.n561 585
R501 B.n673 B.n672 585
R502 B.n674 B.n560 585
R503 B.n676 B.n675 585
R504 B.n678 B.n559 585
R505 B.n681 B.n680 585
R506 B.n682 B.n558 585
R507 B.n684 B.n683 585
R508 B.n686 B.n557 585
R509 B.n689 B.n688 585
R510 B.n690 B.n556 585
R511 B.n692 B.n691 585
R512 B.n694 B.n555 585
R513 B.n697 B.n696 585
R514 B.n698 B.n552 585
R515 B.n701 B.n700 585
R516 B.n703 B.n551 585
R517 B.n706 B.n705 585
R518 B.n707 B.n550 585
R519 B.n709 B.n708 585
R520 B.n711 B.n549 585
R521 B.n714 B.n713 585
R522 B.n715 B.n548 585
R523 B.n720 B.n719 585
R524 B.n722 B.n547 585
R525 B.n725 B.n724 585
R526 B.n726 B.n546 585
R527 B.n728 B.n727 585
R528 B.n730 B.n545 585
R529 B.n733 B.n732 585
R530 B.n734 B.n544 585
R531 B.n736 B.n735 585
R532 B.n738 B.n543 585
R533 B.n741 B.n740 585
R534 B.n742 B.n542 585
R535 B.n744 B.n743 585
R536 B.n746 B.n541 585
R537 B.n749 B.n748 585
R538 B.n750 B.n540 585
R539 B.n752 B.n751 585
R540 B.n754 B.n539 585
R541 B.n757 B.n756 585
R542 B.n758 B.n538 585
R543 B.n760 B.n759 585
R544 B.n762 B.n537 585
R545 B.n765 B.n764 585
R546 B.n766 B.n536 585
R547 B.n768 B.n767 585
R548 B.n770 B.n535 585
R549 B.n773 B.n772 585
R550 B.n774 B.n534 585
R551 B.n776 B.n775 585
R552 B.n778 B.n533 585
R553 B.n781 B.n780 585
R554 B.n782 B.n532 585
R555 B.n784 B.n783 585
R556 B.n786 B.n531 585
R557 B.n789 B.n788 585
R558 B.n790 B.n530 585
R559 B.n792 B.n791 585
R560 B.n794 B.n529 585
R561 B.n797 B.n796 585
R562 B.n798 B.n528 585
R563 B.n800 B.n799 585
R564 B.n802 B.n527 585
R565 B.n805 B.n804 585
R566 B.n806 B.n526 585
R567 B.n808 B.n807 585
R568 B.n810 B.n525 585
R569 B.n813 B.n812 585
R570 B.n814 B.n524 585
R571 B.n816 B.n815 585
R572 B.n818 B.n523 585
R573 B.n821 B.n820 585
R574 B.n822 B.n522 585
R575 B.n824 B.n823 585
R576 B.n826 B.n521 585
R577 B.n829 B.n828 585
R578 B.n830 B.n520 585
R579 B.n832 B.n831 585
R580 B.n834 B.n519 585
R581 B.n837 B.n836 585
R582 B.n838 B.n518 585
R583 B.n843 B.n842 585
R584 B.n842 B.n841 585
R585 B.n844 B.n514 585
R586 B.n514 B.n513 585
R587 B.n846 B.n845 585
R588 B.n847 B.n846 585
R589 B.n508 B.n507 585
R590 B.n509 B.n508 585
R591 B.n855 B.n854 585
R592 B.n854 B.n853 585
R593 B.n856 B.n506 585
R594 B.n506 B.n505 585
R595 B.n858 B.n857 585
R596 B.n859 B.n858 585
R597 B.n500 B.n499 585
R598 B.n501 B.n500 585
R599 B.n867 B.n866 585
R600 B.n866 B.n865 585
R601 B.n868 B.n498 585
R602 B.n498 B.n497 585
R603 B.n870 B.n869 585
R604 B.n871 B.n870 585
R605 B.n492 B.n491 585
R606 B.n493 B.n492 585
R607 B.n879 B.n878 585
R608 B.n878 B.n877 585
R609 B.n880 B.n490 585
R610 B.n490 B.n489 585
R611 B.n882 B.n881 585
R612 B.n883 B.n882 585
R613 B.n484 B.n483 585
R614 B.n485 B.n484 585
R615 B.n891 B.n890 585
R616 B.n890 B.n889 585
R617 B.n892 B.n482 585
R618 B.n482 B.n481 585
R619 B.n894 B.n893 585
R620 B.n895 B.n894 585
R621 B.n476 B.n475 585
R622 B.n477 B.n476 585
R623 B.n903 B.n902 585
R624 B.n902 B.n901 585
R625 B.n904 B.n474 585
R626 B.n474 B.n473 585
R627 B.n906 B.n905 585
R628 B.n907 B.n906 585
R629 B.n468 B.n467 585
R630 B.n469 B.n468 585
R631 B.n915 B.n914 585
R632 B.n914 B.n913 585
R633 B.n916 B.n466 585
R634 B.n466 B.n465 585
R635 B.n918 B.n917 585
R636 B.n919 B.n918 585
R637 B.n460 B.n459 585
R638 B.n461 B.n460 585
R639 B.n927 B.n926 585
R640 B.n926 B.n925 585
R641 B.n928 B.n458 585
R642 B.n458 B.n457 585
R643 B.n930 B.n929 585
R644 B.n931 B.n930 585
R645 B.n452 B.n451 585
R646 B.n453 B.n452 585
R647 B.n940 B.n939 585
R648 B.n939 B.n938 585
R649 B.n941 B.n450 585
R650 B.n937 B.n450 585
R651 B.n943 B.n942 585
R652 B.n944 B.n943 585
R653 B.n445 B.n444 585
R654 B.n446 B.n445 585
R655 B.n952 B.n951 585
R656 B.n951 B.n950 585
R657 B.n953 B.n443 585
R658 B.n443 B.n442 585
R659 B.n955 B.n954 585
R660 B.n956 B.n955 585
R661 B.n437 B.n436 585
R662 B.n438 B.n437 585
R663 B.n964 B.n963 585
R664 B.n963 B.n962 585
R665 B.n965 B.n435 585
R666 B.n435 B.n434 585
R667 B.n967 B.n966 585
R668 B.n968 B.n967 585
R669 B.n429 B.n428 585
R670 B.n430 B.n429 585
R671 B.n976 B.n975 585
R672 B.n975 B.n974 585
R673 B.n977 B.n427 585
R674 B.n427 B.n426 585
R675 B.n979 B.n978 585
R676 B.n980 B.n979 585
R677 B.n421 B.n420 585
R678 B.n422 B.n421 585
R679 B.n989 B.n988 585
R680 B.n988 B.n987 585
R681 B.n990 B.n419 585
R682 B.n419 B.n418 585
R683 B.n992 B.n991 585
R684 B.n993 B.n992 585
R685 B.n2 B.n0 585
R686 B.n4 B.n2 585
R687 B.n3 B.n1 585
R688 B.n1169 B.n3 585
R689 B.n1167 B.n1166 585
R690 B.n1168 B.n1167 585
R691 B.n1165 B.n9 585
R692 B.n9 B.n8 585
R693 B.n1164 B.n1163 585
R694 B.n1163 B.n1162 585
R695 B.n11 B.n10 585
R696 B.n1161 B.n11 585
R697 B.n1159 B.n1158 585
R698 B.n1160 B.n1159 585
R699 B.n1157 B.n16 585
R700 B.n16 B.n15 585
R701 B.n1156 B.n1155 585
R702 B.n1155 B.n1154 585
R703 B.n18 B.n17 585
R704 B.n1153 B.n18 585
R705 B.n1151 B.n1150 585
R706 B.n1152 B.n1151 585
R707 B.n1149 B.n23 585
R708 B.n23 B.n22 585
R709 B.n1148 B.n1147 585
R710 B.n1147 B.n1146 585
R711 B.n25 B.n24 585
R712 B.n1145 B.n25 585
R713 B.n1143 B.n1142 585
R714 B.n1144 B.n1143 585
R715 B.n1141 B.n30 585
R716 B.n30 B.n29 585
R717 B.n1140 B.n1139 585
R718 B.n1139 B.n1138 585
R719 B.n32 B.n31 585
R720 B.n1137 B.n32 585
R721 B.n1135 B.n1134 585
R722 B.n1136 B.n1135 585
R723 B.n1133 B.n36 585
R724 B.n39 B.n36 585
R725 B.n1132 B.n1131 585
R726 B.n1131 B.n1130 585
R727 B.n38 B.n37 585
R728 B.n1129 B.n38 585
R729 B.n1127 B.n1126 585
R730 B.n1128 B.n1127 585
R731 B.n1125 B.n44 585
R732 B.n44 B.n43 585
R733 B.n1124 B.n1123 585
R734 B.n1123 B.n1122 585
R735 B.n46 B.n45 585
R736 B.n1121 B.n46 585
R737 B.n1119 B.n1118 585
R738 B.n1120 B.n1119 585
R739 B.n1117 B.n51 585
R740 B.n51 B.n50 585
R741 B.n1116 B.n1115 585
R742 B.n1115 B.n1114 585
R743 B.n53 B.n52 585
R744 B.n1113 B.n53 585
R745 B.n1111 B.n1110 585
R746 B.n1112 B.n1111 585
R747 B.n1109 B.n58 585
R748 B.n58 B.n57 585
R749 B.n1108 B.n1107 585
R750 B.n1107 B.n1106 585
R751 B.n60 B.n59 585
R752 B.n1105 B.n60 585
R753 B.n1103 B.n1102 585
R754 B.n1104 B.n1103 585
R755 B.n1101 B.n65 585
R756 B.n65 B.n64 585
R757 B.n1100 B.n1099 585
R758 B.n1099 B.n1098 585
R759 B.n67 B.n66 585
R760 B.n1097 B.n67 585
R761 B.n1095 B.n1094 585
R762 B.n1096 B.n1095 585
R763 B.n1093 B.n72 585
R764 B.n72 B.n71 585
R765 B.n1092 B.n1091 585
R766 B.n1091 B.n1090 585
R767 B.n74 B.n73 585
R768 B.n1089 B.n74 585
R769 B.n1087 B.n1086 585
R770 B.n1088 B.n1087 585
R771 B.n1085 B.n79 585
R772 B.n79 B.n78 585
R773 B.n1084 B.n1083 585
R774 B.n1083 B.n1082 585
R775 B.n81 B.n80 585
R776 B.n1081 B.n81 585
R777 B.n1079 B.n1078 585
R778 B.n1080 B.n1079 585
R779 B.n1077 B.n86 585
R780 B.n86 B.n85 585
R781 B.n1076 B.n1075 585
R782 B.n1075 B.n1074 585
R783 B.n88 B.n87 585
R784 B.n1073 B.n88 585
R785 B.n1071 B.n1070 585
R786 B.n1072 B.n1071 585
R787 B.n1069 B.n93 585
R788 B.n93 B.n92 585
R789 B.n1068 B.n1067 585
R790 B.n1067 B.n1066 585
R791 B.n1172 B.n1171 585
R792 B.n1171 B.n1170 585
R793 B.n842 B.n516 482.89
R794 B.n1067 B.n95 482.89
R795 B.n840 B.n518 482.89
R796 B.n1064 B.n96 482.89
R797 B.n716 B.t6 334.387
R798 B.n553 B.t10 334.387
R799 B.n164 B.t13 334.387
R800 B.n161 B.t17 334.387
R801 B.n1065 B.n159 256.663
R802 B.n1065 B.n158 256.663
R803 B.n1065 B.n157 256.663
R804 B.n1065 B.n156 256.663
R805 B.n1065 B.n155 256.663
R806 B.n1065 B.n154 256.663
R807 B.n1065 B.n153 256.663
R808 B.n1065 B.n152 256.663
R809 B.n1065 B.n151 256.663
R810 B.n1065 B.n150 256.663
R811 B.n1065 B.n149 256.663
R812 B.n1065 B.n148 256.663
R813 B.n1065 B.n147 256.663
R814 B.n1065 B.n146 256.663
R815 B.n1065 B.n145 256.663
R816 B.n1065 B.n144 256.663
R817 B.n1065 B.n143 256.663
R818 B.n1065 B.n142 256.663
R819 B.n1065 B.n141 256.663
R820 B.n1065 B.n140 256.663
R821 B.n1065 B.n139 256.663
R822 B.n1065 B.n138 256.663
R823 B.n1065 B.n137 256.663
R824 B.n1065 B.n136 256.663
R825 B.n1065 B.n135 256.663
R826 B.n1065 B.n134 256.663
R827 B.n1065 B.n133 256.663
R828 B.n1065 B.n132 256.663
R829 B.n1065 B.n131 256.663
R830 B.n1065 B.n130 256.663
R831 B.n1065 B.n129 256.663
R832 B.n1065 B.n128 256.663
R833 B.n1065 B.n127 256.663
R834 B.n1065 B.n126 256.663
R835 B.n1065 B.n125 256.663
R836 B.n1065 B.n124 256.663
R837 B.n1065 B.n123 256.663
R838 B.n1065 B.n122 256.663
R839 B.n1065 B.n121 256.663
R840 B.n1065 B.n120 256.663
R841 B.n1065 B.n119 256.663
R842 B.n1065 B.n118 256.663
R843 B.n1065 B.n117 256.663
R844 B.n1065 B.n116 256.663
R845 B.n1065 B.n115 256.663
R846 B.n1065 B.n114 256.663
R847 B.n1065 B.n113 256.663
R848 B.n1065 B.n112 256.663
R849 B.n1065 B.n111 256.663
R850 B.n1065 B.n110 256.663
R851 B.n1065 B.n109 256.663
R852 B.n1065 B.n108 256.663
R853 B.n1065 B.n107 256.663
R854 B.n1065 B.n106 256.663
R855 B.n1065 B.n105 256.663
R856 B.n1065 B.n104 256.663
R857 B.n1065 B.n103 256.663
R858 B.n1065 B.n102 256.663
R859 B.n1065 B.n101 256.663
R860 B.n1065 B.n100 256.663
R861 B.n1065 B.n99 256.663
R862 B.n1065 B.n98 256.663
R863 B.n1065 B.n97 256.663
R864 B.n583 B.n517 256.663
R865 B.n589 B.n517 256.663
R866 B.n591 B.n517 256.663
R867 B.n597 B.n517 256.663
R868 B.n599 B.n517 256.663
R869 B.n605 B.n517 256.663
R870 B.n607 B.n517 256.663
R871 B.n613 B.n517 256.663
R872 B.n615 B.n517 256.663
R873 B.n621 B.n517 256.663
R874 B.n623 B.n517 256.663
R875 B.n629 B.n517 256.663
R876 B.n631 B.n517 256.663
R877 B.n637 B.n517 256.663
R878 B.n639 B.n517 256.663
R879 B.n645 B.n517 256.663
R880 B.n647 B.n517 256.663
R881 B.n653 B.n517 256.663
R882 B.n655 B.n517 256.663
R883 B.n661 B.n517 256.663
R884 B.n663 B.n517 256.663
R885 B.n669 B.n517 256.663
R886 B.n671 B.n517 256.663
R887 B.n677 B.n517 256.663
R888 B.n679 B.n517 256.663
R889 B.n685 B.n517 256.663
R890 B.n687 B.n517 256.663
R891 B.n693 B.n517 256.663
R892 B.n695 B.n517 256.663
R893 B.n702 B.n517 256.663
R894 B.n704 B.n517 256.663
R895 B.n710 B.n517 256.663
R896 B.n712 B.n517 256.663
R897 B.n721 B.n517 256.663
R898 B.n723 B.n517 256.663
R899 B.n729 B.n517 256.663
R900 B.n731 B.n517 256.663
R901 B.n737 B.n517 256.663
R902 B.n739 B.n517 256.663
R903 B.n745 B.n517 256.663
R904 B.n747 B.n517 256.663
R905 B.n753 B.n517 256.663
R906 B.n755 B.n517 256.663
R907 B.n761 B.n517 256.663
R908 B.n763 B.n517 256.663
R909 B.n769 B.n517 256.663
R910 B.n771 B.n517 256.663
R911 B.n777 B.n517 256.663
R912 B.n779 B.n517 256.663
R913 B.n785 B.n517 256.663
R914 B.n787 B.n517 256.663
R915 B.n793 B.n517 256.663
R916 B.n795 B.n517 256.663
R917 B.n801 B.n517 256.663
R918 B.n803 B.n517 256.663
R919 B.n809 B.n517 256.663
R920 B.n811 B.n517 256.663
R921 B.n817 B.n517 256.663
R922 B.n819 B.n517 256.663
R923 B.n825 B.n517 256.663
R924 B.n827 B.n517 256.663
R925 B.n833 B.n517 256.663
R926 B.n835 B.n517 256.663
R927 B.n842 B.n514 163.367
R928 B.n846 B.n514 163.367
R929 B.n846 B.n508 163.367
R930 B.n854 B.n508 163.367
R931 B.n854 B.n506 163.367
R932 B.n858 B.n506 163.367
R933 B.n858 B.n500 163.367
R934 B.n866 B.n500 163.367
R935 B.n866 B.n498 163.367
R936 B.n870 B.n498 163.367
R937 B.n870 B.n492 163.367
R938 B.n878 B.n492 163.367
R939 B.n878 B.n490 163.367
R940 B.n882 B.n490 163.367
R941 B.n882 B.n484 163.367
R942 B.n890 B.n484 163.367
R943 B.n890 B.n482 163.367
R944 B.n894 B.n482 163.367
R945 B.n894 B.n476 163.367
R946 B.n902 B.n476 163.367
R947 B.n902 B.n474 163.367
R948 B.n906 B.n474 163.367
R949 B.n906 B.n468 163.367
R950 B.n914 B.n468 163.367
R951 B.n914 B.n466 163.367
R952 B.n918 B.n466 163.367
R953 B.n918 B.n460 163.367
R954 B.n926 B.n460 163.367
R955 B.n926 B.n458 163.367
R956 B.n930 B.n458 163.367
R957 B.n930 B.n452 163.367
R958 B.n939 B.n452 163.367
R959 B.n939 B.n450 163.367
R960 B.n943 B.n450 163.367
R961 B.n943 B.n445 163.367
R962 B.n951 B.n445 163.367
R963 B.n951 B.n443 163.367
R964 B.n955 B.n443 163.367
R965 B.n955 B.n437 163.367
R966 B.n963 B.n437 163.367
R967 B.n963 B.n435 163.367
R968 B.n967 B.n435 163.367
R969 B.n967 B.n429 163.367
R970 B.n975 B.n429 163.367
R971 B.n975 B.n427 163.367
R972 B.n979 B.n427 163.367
R973 B.n979 B.n421 163.367
R974 B.n988 B.n421 163.367
R975 B.n988 B.n419 163.367
R976 B.n992 B.n419 163.367
R977 B.n992 B.n2 163.367
R978 B.n1171 B.n2 163.367
R979 B.n1171 B.n3 163.367
R980 B.n1167 B.n3 163.367
R981 B.n1167 B.n9 163.367
R982 B.n1163 B.n9 163.367
R983 B.n1163 B.n11 163.367
R984 B.n1159 B.n11 163.367
R985 B.n1159 B.n16 163.367
R986 B.n1155 B.n16 163.367
R987 B.n1155 B.n18 163.367
R988 B.n1151 B.n18 163.367
R989 B.n1151 B.n23 163.367
R990 B.n1147 B.n23 163.367
R991 B.n1147 B.n25 163.367
R992 B.n1143 B.n25 163.367
R993 B.n1143 B.n30 163.367
R994 B.n1139 B.n30 163.367
R995 B.n1139 B.n32 163.367
R996 B.n1135 B.n32 163.367
R997 B.n1135 B.n36 163.367
R998 B.n1131 B.n36 163.367
R999 B.n1131 B.n38 163.367
R1000 B.n1127 B.n38 163.367
R1001 B.n1127 B.n44 163.367
R1002 B.n1123 B.n44 163.367
R1003 B.n1123 B.n46 163.367
R1004 B.n1119 B.n46 163.367
R1005 B.n1119 B.n51 163.367
R1006 B.n1115 B.n51 163.367
R1007 B.n1115 B.n53 163.367
R1008 B.n1111 B.n53 163.367
R1009 B.n1111 B.n58 163.367
R1010 B.n1107 B.n58 163.367
R1011 B.n1107 B.n60 163.367
R1012 B.n1103 B.n60 163.367
R1013 B.n1103 B.n65 163.367
R1014 B.n1099 B.n65 163.367
R1015 B.n1099 B.n67 163.367
R1016 B.n1095 B.n67 163.367
R1017 B.n1095 B.n72 163.367
R1018 B.n1091 B.n72 163.367
R1019 B.n1091 B.n74 163.367
R1020 B.n1087 B.n74 163.367
R1021 B.n1087 B.n79 163.367
R1022 B.n1083 B.n79 163.367
R1023 B.n1083 B.n81 163.367
R1024 B.n1079 B.n81 163.367
R1025 B.n1079 B.n86 163.367
R1026 B.n1075 B.n86 163.367
R1027 B.n1075 B.n88 163.367
R1028 B.n1071 B.n88 163.367
R1029 B.n1071 B.n93 163.367
R1030 B.n1067 B.n93 163.367
R1031 B.n584 B.n582 163.367
R1032 B.n588 B.n582 163.367
R1033 B.n592 B.n590 163.367
R1034 B.n596 B.n580 163.367
R1035 B.n600 B.n598 163.367
R1036 B.n604 B.n578 163.367
R1037 B.n608 B.n606 163.367
R1038 B.n612 B.n576 163.367
R1039 B.n616 B.n614 163.367
R1040 B.n620 B.n574 163.367
R1041 B.n624 B.n622 163.367
R1042 B.n628 B.n572 163.367
R1043 B.n632 B.n630 163.367
R1044 B.n636 B.n570 163.367
R1045 B.n640 B.n638 163.367
R1046 B.n644 B.n568 163.367
R1047 B.n648 B.n646 163.367
R1048 B.n652 B.n566 163.367
R1049 B.n656 B.n654 163.367
R1050 B.n660 B.n564 163.367
R1051 B.n664 B.n662 163.367
R1052 B.n668 B.n562 163.367
R1053 B.n672 B.n670 163.367
R1054 B.n676 B.n560 163.367
R1055 B.n680 B.n678 163.367
R1056 B.n684 B.n558 163.367
R1057 B.n688 B.n686 163.367
R1058 B.n692 B.n556 163.367
R1059 B.n696 B.n694 163.367
R1060 B.n701 B.n552 163.367
R1061 B.n705 B.n703 163.367
R1062 B.n709 B.n550 163.367
R1063 B.n713 B.n711 163.367
R1064 B.n720 B.n548 163.367
R1065 B.n724 B.n722 163.367
R1066 B.n728 B.n546 163.367
R1067 B.n732 B.n730 163.367
R1068 B.n736 B.n544 163.367
R1069 B.n740 B.n738 163.367
R1070 B.n744 B.n542 163.367
R1071 B.n748 B.n746 163.367
R1072 B.n752 B.n540 163.367
R1073 B.n756 B.n754 163.367
R1074 B.n760 B.n538 163.367
R1075 B.n764 B.n762 163.367
R1076 B.n768 B.n536 163.367
R1077 B.n772 B.n770 163.367
R1078 B.n776 B.n534 163.367
R1079 B.n780 B.n778 163.367
R1080 B.n784 B.n532 163.367
R1081 B.n788 B.n786 163.367
R1082 B.n792 B.n530 163.367
R1083 B.n796 B.n794 163.367
R1084 B.n800 B.n528 163.367
R1085 B.n804 B.n802 163.367
R1086 B.n808 B.n526 163.367
R1087 B.n812 B.n810 163.367
R1088 B.n816 B.n524 163.367
R1089 B.n820 B.n818 163.367
R1090 B.n824 B.n522 163.367
R1091 B.n828 B.n826 163.367
R1092 B.n832 B.n520 163.367
R1093 B.n836 B.n834 163.367
R1094 B.n840 B.n512 163.367
R1095 B.n848 B.n512 163.367
R1096 B.n848 B.n510 163.367
R1097 B.n852 B.n510 163.367
R1098 B.n852 B.n504 163.367
R1099 B.n860 B.n504 163.367
R1100 B.n860 B.n502 163.367
R1101 B.n864 B.n502 163.367
R1102 B.n864 B.n496 163.367
R1103 B.n872 B.n496 163.367
R1104 B.n872 B.n494 163.367
R1105 B.n876 B.n494 163.367
R1106 B.n876 B.n488 163.367
R1107 B.n884 B.n488 163.367
R1108 B.n884 B.n486 163.367
R1109 B.n888 B.n486 163.367
R1110 B.n888 B.n480 163.367
R1111 B.n896 B.n480 163.367
R1112 B.n896 B.n478 163.367
R1113 B.n900 B.n478 163.367
R1114 B.n900 B.n472 163.367
R1115 B.n908 B.n472 163.367
R1116 B.n908 B.n470 163.367
R1117 B.n912 B.n470 163.367
R1118 B.n912 B.n464 163.367
R1119 B.n920 B.n464 163.367
R1120 B.n920 B.n462 163.367
R1121 B.n924 B.n462 163.367
R1122 B.n924 B.n456 163.367
R1123 B.n932 B.n456 163.367
R1124 B.n932 B.n454 163.367
R1125 B.n936 B.n454 163.367
R1126 B.n936 B.n449 163.367
R1127 B.n945 B.n449 163.367
R1128 B.n945 B.n447 163.367
R1129 B.n949 B.n447 163.367
R1130 B.n949 B.n441 163.367
R1131 B.n957 B.n441 163.367
R1132 B.n957 B.n439 163.367
R1133 B.n961 B.n439 163.367
R1134 B.n961 B.n433 163.367
R1135 B.n969 B.n433 163.367
R1136 B.n969 B.n431 163.367
R1137 B.n973 B.n431 163.367
R1138 B.n973 B.n425 163.367
R1139 B.n981 B.n425 163.367
R1140 B.n981 B.n423 163.367
R1141 B.n986 B.n423 163.367
R1142 B.n986 B.n417 163.367
R1143 B.n994 B.n417 163.367
R1144 B.n995 B.n994 163.367
R1145 B.n995 B.n5 163.367
R1146 B.n6 B.n5 163.367
R1147 B.n7 B.n6 163.367
R1148 B.n1000 B.n7 163.367
R1149 B.n1000 B.n12 163.367
R1150 B.n13 B.n12 163.367
R1151 B.n14 B.n13 163.367
R1152 B.n1005 B.n14 163.367
R1153 B.n1005 B.n19 163.367
R1154 B.n20 B.n19 163.367
R1155 B.n21 B.n20 163.367
R1156 B.n1010 B.n21 163.367
R1157 B.n1010 B.n26 163.367
R1158 B.n27 B.n26 163.367
R1159 B.n28 B.n27 163.367
R1160 B.n1015 B.n28 163.367
R1161 B.n1015 B.n33 163.367
R1162 B.n34 B.n33 163.367
R1163 B.n35 B.n34 163.367
R1164 B.n1020 B.n35 163.367
R1165 B.n1020 B.n40 163.367
R1166 B.n41 B.n40 163.367
R1167 B.n42 B.n41 163.367
R1168 B.n1025 B.n42 163.367
R1169 B.n1025 B.n47 163.367
R1170 B.n48 B.n47 163.367
R1171 B.n49 B.n48 163.367
R1172 B.n1030 B.n49 163.367
R1173 B.n1030 B.n54 163.367
R1174 B.n55 B.n54 163.367
R1175 B.n56 B.n55 163.367
R1176 B.n1035 B.n56 163.367
R1177 B.n1035 B.n61 163.367
R1178 B.n62 B.n61 163.367
R1179 B.n63 B.n62 163.367
R1180 B.n1040 B.n63 163.367
R1181 B.n1040 B.n68 163.367
R1182 B.n69 B.n68 163.367
R1183 B.n70 B.n69 163.367
R1184 B.n1045 B.n70 163.367
R1185 B.n1045 B.n75 163.367
R1186 B.n76 B.n75 163.367
R1187 B.n77 B.n76 163.367
R1188 B.n1050 B.n77 163.367
R1189 B.n1050 B.n82 163.367
R1190 B.n83 B.n82 163.367
R1191 B.n84 B.n83 163.367
R1192 B.n1055 B.n84 163.367
R1193 B.n1055 B.n89 163.367
R1194 B.n90 B.n89 163.367
R1195 B.n91 B.n90 163.367
R1196 B.n1060 B.n91 163.367
R1197 B.n1060 B.n96 163.367
R1198 B.n168 B.n167 163.367
R1199 B.n172 B.n171 163.367
R1200 B.n176 B.n175 163.367
R1201 B.n180 B.n179 163.367
R1202 B.n184 B.n183 163.367
R1203 B.n188 B.n187 163.367
R1204 B.n192 B.n191 163.367
R1205 B.n196 B.n195 163.367
R1206 B.n200 B.n199 163.367
R1207 B.n204 B.n203 163.367
R1208 B.n208 B.n207 163.367
R1209 B.n212 B.n211 163.367
R1210 B.n216 B.n215 163.367
R1211 B.n220 B.n219 163.367
R1212 B.n224 B.n223 163.367
R1213 B.n228 B.n227 163.367
R1214 B.n232 B.n231 163.367
R1215 B.n236 B.n235 163.367
R1216 B.n240 B.n239 163.367
R1217 B.n244 B.n243 163.367
R1218 B.n248 B.n247 163.367
R1219 B.n252 B.n251 163.367
R1220 B.n256 B.n255 163.367
R1221 B.n260 B.n259 163.367
R1222 B.n264 B.n263 163.367
R1223 B.n268 B.n267 163.367
R1224 B.n272 B.n271 163.367
R1225 B.n276 B.n275 163.367
R1226 B.n280 B.n279 163.367
R1227 B.n285 B.n284 163.367
R1228 B.n289 B.n288 163.367
R1229 B.n293 B.n292 163.367
R1230 B.n297 B.n296 163.367
R1231 B.n301 B.n300 163.367
R1232 B.n305 B.n304 163.367
R1233 B.n309 B.n308 163.367
R1234 B.n313 B.n312 163.367
R1235 B.n317 B.n316 163.367
R1236 B.n321 B.n320 163.367
R1237 B.n325 B.n324 163.367
R1238 B.n329 B.n328 163.367
R1239 B.n333 B.n332 163.367
R1240 B.n337 B.n336 163.367
R1241 B.n341 B.n340 163.367
R1242 B.n345 B.n344 163.367
R1243 B.n349 B.n348 163.367
R1244 B.n353 B.n352 163.367
R1245 B.n357 B.n356 163.367
R1246 B.n361 B.n360 163.367
R1247 B.n365 B.n364 163.367
R1248 B.n369 B.n368 163.367
R1249 B.n373 B.n372 163.367
R1250 B.n377 B.n376 163.367
R1251 B.n381 B.n380 163.367
R1252 B.n385 B.n384 163.367
R1253 B.n389 B.n388 163.367
R1254 B.n393 B.n392 163.367
R1255 B.n397 B.n396 163.367
R1256 B.n401 B.n400 163.367
R1257 B.n405 B.n404 163.367
R1258 B.n409 B.n408 163.367
R1259 B.n413 B.n412 163.367
R1260 B.n1064 B.n160 163.367
R1261 B.n716 B.t9 140.962
R1262 B.n161 B.t18 140.962
R1263 B.n553 B.t12 140.938
R1264 B.n164 B.t15 140.938
R1265 B.n717 B.n716 72.5338
R1266 B.n554 B.n553 72.5338
R1267 B.n165 B.n164 72.5338
R1268 B.n162 B.n161 72.5338
R1269 B.n583 B.n516 71.676
R1270 B.n589 B.n588 71.676
R1271 B.n592 B.n591 71.676
R1272 B.n597 B.n596 71.676
R1273 B.n600 B.n599 71.676
R1274 B.n605 B.n604 71.676
R1275 B.n608 B.n607 71.676
R1276 B.n613 B.n612 71.676
R1277 B.n616 B.n615 71.676
R1278 B.n621 B.n620 71.676
R1279 B.n624 B.n623 71.676
R1280 B.n629 B.n628 71.676
R1281 B.n632 B.n631 71.676
R1282 B.n637 B.n636 71.676
R1283 B.n640 B.n639 71.676
R1284 B.n645 B.n644 71.676
R1285 B.n648 B.n647 71.676
R1286 B.n653 B.n652 71.676
R1287 B.n656 B.n655 71.676
R1288 B.n661 B.n660 71.676
R1289 B.n664 B.n663 71.676
R1290 B.n669 B.n668 71.676
R1291 B.n672 B.n671 71.676
R1292 B.n677 B.n676 71.676
R1293 B.n680 B.n679 71.676
R1294 B.n685 B.n684 71.676
R1295 B.n688 B.n687 71.676
R1296 B.n693 B.n692 71.676
R1297 B.n696 B.n695 71.676
R1298 B.n702 B.n701 71.676
R1299 B.n705 B.n704 71.676
R1300 B.n710 B.n709 71.676
R1301 B.n713 B.n712 71.676
R1302 B.n721 B.n720 71.676
R1303 B.n724 B.n723 71.676
R1304 B.n729 B.n728 71.676
R1305 B.n732 B.n731 71.676
R1306 B.n737 B.n736 71.676
R1307 B.n740 B.n739 71.676
R1308 B.n745 B.n744 71.676
R1309 B.n748 B.n747 71.676
R1310 B.n753 B.n752 71.676
R1311 B.n756 B.n755 71.676
R1312 B.n761 B.n760 71.676
R1313 B.n764 B.n763 71.676
R1314 B.n769 B.n768 71.676
R1315 B.n772 B.n771 71.676
R1316 B.n777 B.n776 71.676
R1317 B.n780 B.n779 71.676
R1318 B.n785 B.n784 71.676
R1319 B.n788 B.n787 71.676
R1320 B.n793 B.n792 71.676
R1321 B.n796 B.n795 71.676
R1322 B.n801 B.n800 71.676
R1323 B.n804 B.n803 71.676
R1324 B.n809 B.n808 71.676
R1325 B.n812 B.n811 71.676
R1326 B.n817 B.n816 71.676
R1327 B.n820 B.n819 71.676
R1328 B.n825 B.n824 71.676
R1329 B.n828 B.n827 71.676
R1330 B.n833 B.n832 71.676
R1331 B.n836 B.n835 71.676
R1332 B.n97 B.n95 71.676
R1333 B.n168 B.n98 71.676
R1334 B.n172 B.n99 71.676
R1335 B.n176 B.n100 71.676
R1336 B.n180 B.n101 71.676
R1337 B.n184 B.n102 71.676
R1338 B.n188 B.n103 71.676
R1339 B.n192 B.n104 71.676
R1340 B.n196 B.n105 71.676
R1341 B.n200 B.n106 71.676
R1342 B.n204 B.n107 71.676
R1343 B.n208 B.n108 71.676
R1344 B.n212 B.n109 71.676
R1345 B.n216 B.n110 71.676
R1346 B.n220 B.n111 71.676
R1347 B.n224 B.n112 71.676
R1348 B.n228 B.n113 71.676
R1349 B.n232 B.n114 71.676
R1350 B.n236 B.n115 71.676
R1351 B.n240 B.n116 71.676
R1352 B.n244 B.n117 71.676
R1353 B.n248 B.n118 71.676
R1354 B.n252 B.n119 71.676
R1355 B.n256 B.n120 71.676
R1356 B.n260 B.n121 71.676
R1357 B.n264 B.n122 71.676
R1358 B.n268 B.n123 71.676
R1359 B.n272 B.n124 71.676
R1360 B.n276 B.n125 71.676
R1361 B.n280 B.n126 71.676
R1362 B.n285 B.n127 71.676
R1363 B.n289 B.n128 71.676
R1364 B.n293 B.n129 71.676
R1365 B.n297 B.n130 71.676
R1366 B.n301 B.n131 71.676
R1367 B.n305 B.n132 71.676
R1368 B.n309 B.n133 71.676
R1369 B.n313 B.n134 71.676
R1370 B.n317 B.n135 71.676
R1371 B.n321 B.n136 71.676
R1372 B.n325 B.n137 71.676
R1373 B.n329 B.n138 71.676
R1374 B.n333 B.n139 71.676
R1375 B.n337 B.n140 71.676
R1376 B.n341 B.n141 71.676
R1377 B.n345 B.n142 71.676
R1378 B.n349 B.n143 71.676
R1379 B.n353 B.n144 71.676
R1380 B.n357 B.n145 71.676
R1381 B.n361 B.n146 71.676
R1382 B.n365 B.n147 71.676
R1383 B.n369 B.n148 71.676
R1384 B.n373 B.n149 71.676
R1385 B.n377 B.n150 71.676
R1386 B.n381 B.n151 71.676
R1387 B.n385 B.n152 71.676
R1388 B.n389 B.n153 71.676
R1389 B.n393 B.n154 71.676
R1390 B.n397 B.n155 71.676
R1391 B.n401 B.n156 71.676
R1392 B.n405 B.n157 71.676
R1393 B.n409 B.n158 71.676
R1394 B.n413 B.n159 71.676
R1395 B.n160 B.n159 71.676
R1396 B.n412 B.n158 71.676
R1397 B.n408 B.n157 71.676
R1398 B.n404 B.n156 71.676
R1399 B.n400 B.n155 71.676
R1400 B.n396 B.n154 71.676
R1401 B.n392 B.n153 71.676
R1402 B.n388 B.n152 71.676
R1403 B.n384 B.n151 71.676
R1404 B.n380 B.n150 71.676
R1405 B.n376 B.n149 71.676
R1406 B.n372 B.n148 71.676
R1407 B.n368 B.n147 71.676
R1408 B.n364 B.n146 71.676
R1409 B.n360 B.n145 71.676
R1410 B.n356 B.n144 71.676
R1411 B.n352 B.n143 71.676
R1412 B.n348 B.n142 71.676
R1413 B.n344 B.n141 71.676
R1414 B.n340 B.n140 71.676
R1415 B.n336 B.n139 71.676
R1416 B.n332 B.n138 71.676
R1417 B.n328 B.n137 71.676
R1418 B.n324 B.n136 71.676
R1419 B.n320 B.n135 71.676
R1420 B.n316 B.n134 71.676
R1421 B.n312 B.n133 71.676
R1422 B.n308 B.n132 71.676
R1423 B.n304 B.n131 71.676
R1424 B.n300 B.n130 71.676
R1425 B.n296 B.n129 71.676
R1426 B.n292 B.n128 71.676
R1427 B.n288 B.n127 71.676
R1428 B.n284 B.n126 71.676
R1429 B.n279 B.n125 71.676
R1430 B.n275 B.n124 71.676
R1431 B.n271 B.n123 71.676
R1432 B.n267 B.n122 71.676
R1433 B.n263 B.n121 71.676
R1434 B.n259 B.n120 71.676
R1435 B.n255 B.n119 71.676
R1436 B.n251 B.n118 71.676
R1437 B.n247 B.n117 71.676
R1438 B.n243 B.n116 71.676
R1439 B.n239 B.n115 71.676
R1440 B.n235 B.n114 71.676
R1441 B.n231 B.n113 71.676
R1442 B.n227 B.n112 71.676
R1443 B.n223 B.n111 71.676
R1444 B.n219 B.n110 71.676
R1445 B.n215 B.n109 71.676
R1446 B.n211 B.n108 71.676
R1447 B.n207 B.n107 71.676
R1448 B.n203 B.n106 71.676
R1449 B.n199 B.n105 71.676
R1450 B.n195 B.n104 71.676
R1451 B.n191 B.n103 71.676
R1452 B.n187 B.n102 71.676
R1453 B.n183 B.n101 71.676
R1454 B.n179 B.n100 71.676
R1455 B.n175 B.n99 71.676
R1456 B.n171 B.n98 71.676
R1457 B.n167 B.n97 71.676
R1458 B.n584 B.n583 71.676
R1459 B.n590 B.n589 71.676
R1460 B.n591 B.n580 71.676
R1461 B.n598 B.n597 71.676
R1462 B.n599 B.n578 71.676
R1463 B.n606 B.n605 71.676
R1464 B.n607 B.n576 71.676
R1465 B.n614 B.n613 71.676
R1466 B.n615 B.n574 71.676
R1467 B.n622 B.n621 71.676
R1468 B.n623 B.n572 71.676
R1469 B.n630 B.n629 71.676
R1470 B.n631 B.n570 71.676
R1471 B.n638 B.n637 71.676
R1472 B.n639 B.n568 71.676
R1473 B.n646 B.n645 71.676
R1474 B.n647 B.n566 71.676
R1475 B.n654 B.n653 71.676
R1476 B.n655 B.n564 71.676
R1477 B.n662 B.n661 71.676
R1478 B.n663 B.n562 71.676
R1479 B.n670 B.n669 71.676
R1480 B.n671 B.n560 71.676
R1481 B.n678 B.n677 71.676
R1482 B.n679 B.n558 71.676
R1483 B.n686 B.n685 71.676
R1484 B.n687 B.n556 71.676
R1485 B.n694 B.n693 71.676
R1486 B.n695 B.n552 71.676
R1487 B.n703 B.n702 71.676
R1488 B.n704 B.n550 71.676
R1489 B.n711 B.n710 71.676
R1490 B.n712 B.n548 71.676
R1491 B.n722 B.n721 71.676
R1492 B.n723 B.n546 71.676
R1493 B.n730 B.n729 71.676
R1494 B.n731 B.n544 71.676
R1495 B.n738 B.n737 71.676
R1496 B.n739 B.n542 71.676
R1497 B.n746 B.n745 71.676
R1498 B.n747 B.n540 71.676
R1499 B.n754 B.n753 71.676
R1500 B.n755 B.n538 71.676
R1501 B.n762 B.n761 71.676
R1502 B.n763 B.n536 71.676
R1503 B.n770 B.n769 71.676
R1504 B.n771 B.n534 71.676
R1505 B.n778 B.n777 71.676
R1506 B.n779 B.n532 71.676
R1507 B.n786 B.n785 71.676
R1508 B.n787 B.n530 71.676
R1509 B.n794 B.n793 71.676
R1510 B.n795 B.n528 71.676
R1511 B.n802 B.n801 71.676
R1512 B.n803 B.n526 71.676
R1513 B.n810 B.n809 71.676
R1514 B.n811 B.n524 71.676
R1515 B.n818 B.n817 71.676
R1516 B.n819 B.n522 71.676
R1517 B.n826 B.n825 71.676
R1518 B.n827 B.n520 71.676
R1519 B.n834 B.n833 71.676
R1520 B.n835 B.n518 71.676
R1521 B.n717 B.t8 68.4282
R1522 B.n162 B.t19 68.4282
R1523 B.n554 B.t11 68.4044
R1524 B.n165 B.t16 68.4044
R1525 B.n841 B.n517 62.6118
R1526 B.n1066 B.n1065 62.6118
R1527 B.n718 B.n717 59.5399
R1528 B.n699 B.n554 59.5399
R1529 B.n282 B.n165 59.5399
R1530 B.n163 B.n162 59.5399
R1531 B.n841 B.n513 32.501
R1532 B.n847 B.n513 32.501
R1533 B.n847 B.n509 32.501
R1534 B.n853 B.n509 32.501
R1535 B.n853 B.n505 32.501
R1536 B.n859 B.n505 32.501
R1537 B.n859 B.n501 32.501
R1538 B.n865 B.n501 32.501
R1539 B.n871 B.n497 32.501
R1540 B.n871 B.n493 32.501
R1541 B.n877 B.n493 32.501
R1542 B.n877 B.n489 32.501
R1543 B.n883 B.n489 32.501
R1544 B.n883 B.n485 32.501
R1545 B.n889 B.n485 32.501
R1546 B.n889 B.n481 32.501
R1547 B.n895 B.n481 32.501
R1548 B.n895 B.n477 32.501
R1549 B.n901 B.n477 32.501
R1550 B.n901 B.n473 32.501
R1551 B.n907 B.n473 32.501
R1552 B.n913 B.n469 32.501
R1553 B.n913 B.n465 32.501
R1554 B.n919 B.n465 32.501
R1555 B.n919 B.n461 32.501
R1556 B.n925 B.n461 32.501
R1557 B.n925 B.n457 32.501
R1558 B.n931 B.n457 32.501
R1559 B.n931 B.n453 32.501
R1560 B.n938 B.n453 32.501
R1561 B.n938 B.n937 32.501
R1562 B.n944 B.n446 32.501
R1563 B.n950 B.n446 32.501
R1564 B.n950 B.n442 32.501
R1565 B.n956 B.n442 32.501
R1566 B.n956 B.n438 32.501
R1567 B.n962 B.n438 32.501
R1568 B.n962 B.n434 32.501
R1569 B.n968 B.n434 32.501
R1570 B.n968 B.n430 32.501
R1571 B.n974 B.n430 32.501
R1572 B.n980 B.n426 32.501
R1573 B.n980 B.n422 32.501
R1574 B.n987 B.n422 32.501
R1575 B.n987 B.n418 32.501
R1576 B.n993 B.n418 32.501
R1577 B.n993 B.n4 32.501
R1578 B.n1170 B.n4 32.501
R1579 B.n1170 B.n1169 32.501
R1580 B.n1169 B.n1168 32.501
R1581 B.n1168 B.n8 32.501
R1582 B.n1162 B.n8 32.501
R1583 B.n1162 B.n1161 32.501
R1584 B.n1161 B.n1160 32.501
R1585 B.n1160 B.n15 32.501
R1586 B.n1154 B.n1153 32.501
R1587 B.n1153 B.n1152 32.501
R1588 B.n1152 B.n22 32.501
R1589 B.n1146 B.n22 32.501
R1590 B.n1146 B.n1145 32.501
R1591 B.n1145 B.n1144 32.501
R1592 B.n1144 B.n29 32.501
R1593 B.n1138 B.n29 32.501
R1594 B.n1138 B.n1137 32.501
R1595 B.n1137 B.n1136 32.501
R1596 B.n1130 B.n39 32.501
R1597 B.n1130 B.n1129 32.501
R1598 B.n1129 B.n1128 32.501
R1599 B.n1128 B.n43 32.501
R1600 B.n1122 B.n43 32.501
R1601 B.n1122 B.n1121 32.501
R1602 B.n1121 B.n1120 32.501
R1603 B.n1120 B.n50 32.501
R1604 B.n1114 B.n50 32.501
R1605 B.n1114 B.n1113 32.501
R1606 B.n1112 B.n57 32.501
R1607 B.n1106 B.n57 32.501
R1608 B.n1106 B.n1105 32.501
R1609 B.n1105 B.n1104 32.501
R1610 B.n1104 B.n64 32.501
R1611 B.n1098 B.n64 32.501
R1612 B.n1098 B.n1097 32.501
R1613 B.n1097 B.n1096 32.501
R1614 B.n1096 B.n71 32.501
R1615 B.n1090 B.n71 32.501
R1616 B.n1090 B.n1089 32.501
R1617 B.n1089 B.n1088 32.501
R1618 B.n1088 B.n78 32.501
R1619 B.n1082 B.n1081 32.501
R1620 B.n1081 B.n1080 32.501
R1621 B.n1080 B.n85 32.501
R1622 B.n1074 B.n85 32.501
R1623 B.n1074 B.n1073 32.501
R1624 B.n1073 B.n1072 32.501
R1625 B.n1072 B.n92 32.501
R1626 B.n1066 B.n92 32.501
R1627 B.n1068 B.n94 31.3761
R1628 B.n1063 B.n1062 31.3761
R1629 B.n839 B.n838 31.3761
R1630 B.n843 B.n515 31.3761
R1631 B.n907 B.t2 29.1554
R1632 B.n937 B.t4 29.1554
R1633 B.n974 B.t0 29.1554
R1634 B.n1154 B.t3 29.1554
R1635 B.n39 B.t5 29.1554
R1636 B.t1 B.n1112 29.1554
R1637 B.n865 B.t7 22.4641
R1638 B.n1082 B.t14 22.4641
R1639 B B.n1172 18.0485
R1640 B.n166 B.n94 10.6151
R1641 B.n169 B.n166 10.6151
R1642 B.n170 B.n169 10.6151
R1643 B.n173 B.n170 10.6151
R1644 B.n174 B.n173 10.6151
R1645 B.n177 B.n174 10.6151
R1646 B.n178 B.n177 10.6151
R1647 B.n181 B.n178 10.6151
R1648 B.n182 B.n181 10.6151
R1649 B.n185 B.n182 10.6151
R1650 B.n186 B.n185 10.6151
R1651 B.n189 B.n186 10.6151
R1652 B.n190 B.n189 10.6151
R1653 B.n193 B.n190 10.6151
R1654 B.n194 B.n193 10.6151
R1655 B.n197 B.n194 10.6151
R1656 B.n198 B.n197 10.6151
R1657 B.n201 B.n198 10.6151
R1658 B.n202 B.n201 10.6151
R1659 B.n205 B.n202 10.6151
R1660 B.n206 B.n205 10.6151
R1661 B.n209 B.n206 10.6151
R1662 B.n210 B.n209 10.6151
R1663 B.n213 B.n210 10.6151
R1664 B.n214 B.n213 10.6151
R1665 B.n217 B.n214 10.6151
R1666 B.n218 B.n217 10.6151
R1667 B.n221 B.n218 10.6151
R1668 B.n222 B.n221 10.6151
R1669 B.n225 B.n222 10.6151
R1670 B.n226 B.n225 10.6151
R1671 B.n229 B.n226 10.6151
R1672 B.n230 B.n229 10.6151
R1673 B.n233 B.n230 10.6151
R1674 B.n234 B.n233 10.6151
R1675 B.n237 B.n234 10.6151
R1676 B.n238 B.n237 10.6151
R1677 B.n241 B.n238 10.6151
R1678 B.n242 B.n241 10.6151
R1679 B.n245 B.n242 10.6151
R1680 B.n246 B.n245 10.6151
R1681 B.n249 B.n246 10.6151
R1682 B.n250 B.n249 10.6151
R1683 B.n253 B.n250 10.6151
R1684 B.n254 B.n253 10.6151
R1685 B.n257 B.n254 10.6151
R1686 B.n258 B.n257 10.6151
R1687 B.n261 B.n258 10.6151
R1688 B.n262 B.n261 10.6151
R1689 B.n265 B.n262 10.6151
R1690 B.n266 B.n265 10.6151
R1691 B.n269 B.n266 10.6151
R1692 B.n270 B.n269 10.6151
R1693 B.n273 B.n270 10.6151
R1694 B.n274 B.n273 10.6151
R1695 B.n277 B.n274 10.6151
R1696 B.n278 B.n277 10.6151
R1697 B.n281 B.n278 10.6151
R1698 B.n286 B.n283 10.6151
R1699 B.n287 B.n286 10.6151
R1700 B.n290 B.n287 10.6151
R1701 B.n291 B.n290 10.6151
R1702 B.n294 B.n291 10.6151
R1703 B.n295 B.n294 10.6151
R1704 B.n298 B.n295 10.6151
R1705 B.n299 B.n298 10.6151
R1706 B.n303 B.n302 10.6151
R1707 B.n306 B.n303 10.6151
R1708 B.n307 B.n306 10.6151
R1709 B.n310 B.n307 10.6151
R1710 B.n311 B.n310 10.6151
R1711 B.n314 B.n311 10.6151
R1712 B.n315 B.n314 10.6151
R1713 B.n318 B.n315 10.6151
R1714 B.n319 B.n318 10.6151
R1715 B.n322 B.n319 10.6151
R1716 B.n323 B.n322 10.6151
R1717 B.n326 B.n323 10.6151
R1718 B.n327 B.n326 10.6151
R1719 B.n330 B.n327 10.6151
R1720 B.n331 B.n330 10.6151
R1721 B.n334 B.n331 10.6151
R1722 B.n335 B.n334 10.6151
R1723 B.n338 B.n335 10.6151
R1724 B.n339 B.n338 10.6151
R1725 B.n342 B.n339 10.6151
R1726 B.n343 B.n342 10.6151
R1727 B.n346 B.n343 10.6151
R1728 B.n347 B.n346 10.6151
R1729 B.n350 B.n347 10.6151
R1730 B.n351 B.n350 10.6151
R1731 B.n354 B.n351 10.6151
R1732 B.n355 B.n354 10.6151
R1733 B.n358 B.n355 10.6151
R1734 B.n359 B.n358 10.6151
R1735 B.n362 B.n359 10.6151
R1736 B.n363 B.n362 10.6151
R1737 B.n366 B.n363 10.6151
R1738 B.n367 B.n366 10.6151
R1739 B.n370 B.n367 10.6151
R1740 B.n371 B.n370 10.6151
R1741 B.n374 B.n371 10.6151
R1742 B.n375 B.n374 10.6151
R1743 B.n378 B.n375 10.6151
R1744 B.n379 B.n378 10.6151
R1745 B.n382 B.n379 10.6151
R1746 B.n383 B.n382 10.6151
R1747 B.n386 B.n383 10.6151
R1748 B.n387 B.n386 10.6151
R1749 B.n390 B.n387 10.6151
R1750 B.n391 B.n390 10.6151
R1751 B.n394 B.n391 10.6151
R1752 B.n395 B.n394 10.6151
R1753 B.n398 B.n395 10.6151
R1754 B.n399 B.n398 10.6151
R1755 B.n402 B.n399 10.6151
R1756 B.n403 B.n402 10.6151
R1757 B.n406 B.n403 10.6151
R1758 B.n407 B.n406 10.6151
R1759 B.n410 B.n407 10.6151
R1760 B.n411 B.n410 10.6151
R1761 B.n414 B.n411 10.6151
R1762 B.n415 B.n414 10.6151
R1763 B.n1063 B.n415 10.6151
R1764 B.n839 B.n511 10.6151
R1765 B.n849 B.n511 10.6151
R1766 B.n850 B.n849 10.6151
R1767 B.n851 B.n850 10.6151
R1768 B.n851 B.n503 10.6151
R1769 B.n861 B.n503 10.6151
R1770 B.n862 B.n861 10.6151
R1771 B.n863 B.n862 10.6151
R1772 B.n863 B.n495 10.6151
R1773 B.n873 B.n495 10.6151
R1774 B.n874 B.n873 10.6151
R1775 B.n875 B.n874 10.6151
R1776 B.n875 B.n487 10.6151
R1777 B.n885 B.n487 10.6151
R1778 B.n886 B.n885 10.6151
R1779 B.n887 B.n886 10.6151
R1780 B.n887 B.n479 10.6151
R1781 B.n897 B.n479 10.6151
R1782 B.n898 B.n897 10.6151
R1783 B.n899 B.n898 10.6151
R1784 B.n899 B.n471 10.6151
R1785 B.n909 B.n471 10.6151
R1786 B.n910 B.n909 10.6151
R1787 B.n911 B.n910 10.6151
R1788 B.n911 B.n463 10.6151
R1789 B.n921 B.n463 10.6151
R1790 B.n922 B.n921 10.6151
R1791 B.n923 B.n922 10.6151
R1792 B.n923 B.n455 10.6151
R1793 B.n933 B.n455 10.6151
R1794 B.n934 B.n933 10.6151
R1795 B.n935 B.n934 10.6151
R1796 B.n935 B.n448 10.6151
R1797 B.n946 B.n448 10.6151
R1798 B.n947 B.n946 10.6151
R1799 B.n948 B.n947 10.6151
R1800 B.n948 B.n440 10.6151
R1801 B.n958 B.n440 10.6151
R1802 B.n959 B.n958 10.6151
R1803 B.n960 B.n959 10.6151
R1804 B.n960 B.n432 10.6151
R1805 B.n970 B.n432 10.6151
R1806 B.n971 B.n970 10.6151
R1807 B.n972 B.n971 10.6151
R1808 B.n972 B.n424 10.6151
R1809 B.n982 B.n424 10.6151
R1810 B.n983 B.n982 10.6151
R1811 B.n985 B.n983 10.6151
R1812 B.n985 B.n984 10.6151
R1813 B.n984 B.n416 10.6151
R1814 B.n996 B.n416 10.6151
R1815 B.n997 B.n996 10.6151
R1816 B.n998 B.n997 10.6151
R1817 B.n999 B.n998 10.6151
R1818 B.n1001 B.n999 10.6151
R1819 B.n1002 B.n1001 10.6151
R1820 B.n1003 B.n1002 10.6151
R1821 B.n1004 B.n1003 10.6151
R1822 B.n1006 B.n1004 10.6151
R1823 B.n1007 B.n1006 10.6151
R1824 B.n1008 B.n1007 10.6151
R1825 B.n1009 B.n1008 10.6151
R1826 B.n1011 B.n1009 10.6151
R1827 B.n1012 B.n1011 10.6151
R1828 B.n1013 B.n1012 10.6151
R1829 B.n1014 B.n1013 10.6151
R1830 B.n1016 B.n1014 10.6151
R1831 B.n1017 B.n1016 10.6151
R1832 B.n1018 B.n1017 10.6151
R1833 B.n1019 B.n1018 10.6151
R1834 B.n1021 B.n1019 10.6151
R1835 B.n1022 B.n1021 10.6151
R1836 B.n1023 B.n1022 10.6151
R1837 B.n1024 B.n1023 10.6151
R1838 B.n1026 B.n1024 10.6151
R1839 B.n1027 B.n1026 10.6151
R1840 B.n1028 B.n1027 10.6151
R1841 B.n1029 B.n1028 10.6151
R1842 B.n1031 B.n1029 10.6151
R1843 B.n1032 B.n1031 10.6151
R1844 B.n1033 B.n1032 10.6151
R1845 B.n1034 B.n1033 10.6151
R1846 B.n1036 B.n1034 10.6151
R1847 B.n1037 B.n1036 10.6151
R1848 B.n1038 B.n1037 10.6151
R1849 B.n1039 B.n1038 10.6151
R1850 B.n1041 B.n1039 10.6151
R1851 B.n1042 B.n1041 10.6151
R1852 B.n1043 B.n1042 10.6151
R1853 B.n1044 B.n1043 10.6151
R1854 B.n1046 B.n1044 10.6151
R1855 B.n1047 B.n1046 10.6151
R1856 B.n1048 B.n1047 10.6151
R1857 B.n1049 B.n1048 10.6151
R1858 B.n1051 B.n1049 10.6151
R1859 B.n1052 B.n1051 10.6151
R1860 B.n1053 B.n1052 10.6151
R1861 B.n1054 B.n1053 10.6151
R1862 B.n1056 B.n1054 10.6151
R1863 B.n1057 B.n1056 10.6151
R1864 B.n1058 B.n1057 10.6151
R1865 B.n1059 B.n1058 10.6151
R1866 B.n1061 B.n1059 10.6151
R1867 B.n1062 B.n1061 10.6151
R1868 B.n585 B.n515 10.6151
R1869 B.n586 B.n585 10.6151
R1870 B.n587 B.n586 10.6151
R1871 B.n587 B.n581 10.6151
R1872 B.n593 B.n581 10.6151
R1873 B.n594 B.n593 10.6151
R1874 B.n595 B.n594 10.6151
R1875 B.n595 B.n579 10.6151
R1876 B.n601 B.n579 10.6151
R1877 B.n602 B.n601 10.6151
R1878 B.n603 B.n602 10.6151
R1879 B.n603 B.n577 10.6151
R1880 B.n609 B.n577 10.6151
R1881 B.n610 B.n609 10.6151
R1882 B.n611 B.n610 10.6151
R1883 B.n611 B.n575 10.6151
R1884 B.n617 B.n575 10.6151
R1885 B.n618 B.n617 10.6151
R1886 B.n619 B.n618 10.6151
R1887 B.n619 B.n573 10.6151
R1888 B.n625 B.n573 10.6151
R1889 B.n626 B.n625 10.6151
R1890 B.n627 B.n626 10.6151
R1891 B.n627 B.n571 10.6151
R1892 B.n633 B.n571 10.6151
R1893 B.n634 B.n633 10.6151
R1894 B.n635 B.n634 10.6151
R1895 B.n635 B.n569 10.6151
R1896 B.n641 B.n569 10.6151
R1897 B.n642 B.n641 10.6151
R1898 B.n643 B.n642 10.6151
R1899 B.n643 B.n567 10.6151
R1900 B.n649 B.n567 10.6151
R1901 B.n650 B.n649 10.6151
R1902 B.n651 B.n650 10.6151
R1903 B.n651 B.n565 10.6151
R1904 B.n657 B.n565 10.6151
R1905 B.n658 B.n657 10.6151
R1906 B.n659 B.n658 10.6151
R1907 B.n659 B.n563 10.6151
R1908 B.n665 B.n563 10.6151
R1909 B.n666 B.n665 10.6151
R1910 B.n667 B.n666 10.6151
R1911 B.n667 B.n561 10.6151
R1912 B.n673 B.n561 10.6151
R1913 B.n674 B.n673 10.6151
R1914 B.n675 B.n674 10.6151
R1915 B.n675 B.n559 10.6151
R1916 B.n681 B.n559 10.6151
R1917 B.n682 B.n681 10.6151
R1918 B.n683 B.n682 10.6151
R1919 B.n683 B.n557 10.6151
R1920 B.n689 B.n557 10.6151
R1921 B.n690 B.n689 10.6151
R1922 B.n691 B.n690 10.6151
R1923 B.n691 B.n555 10.6151
R1924 B.n697 B.n555 10.6151
R1925 B.n698 B.n697 10.6151
R1926 B.n700 B.n551 10.6151
R1927 B.n706 B.n551 10.6151
R1928 B.n707 B.n706 10.6151
R1929 B.n708 B.n707 10.6151
R1930 B.n708 B.n549 10.6151
R1931 B.n714 B.n549 10.6151
R1932 B.n715 B.n714 10.6151
R1933 B.n719 B.n715 10.6151
R1934 B.n725 B.n547 10.6151
R1935 B.n726 B.n725 10.6151
R1936 B.n727 B.n726 10.6151
R1937 B.n727 B.n545 10.6151
R1938 B.n733 B.n545 10.6151
R1939 B.n734 B.n733 10.6151
R1940 B.n735 B.n734 10.6151
R1941 B.n735 B.n543 10.6151
R1942 B.n741 B.n543 10.6151
R1943 B.n742 B.n741 10.6151
R1944 B.n743 B.n742 10.6151
R1945 B.n743 B.n541 10.6151
R1946 B.n749 B.n541 10.6151
R1947 B.n750 B.n749 10.6151
R1948 B.n751 B.n750 10.6151
R1949 B.n751 B.n539 10.6151
R1950 B.n757 B.n539 10.6151
R1951 B.n758 B.n757 10.6151
R1952 B.n759 B.n758 10.6151
R1953 B.n759 B.n537 10.6151
R1954 B.n765 B.n537 10.6151
R1955 B.n766 B.n765 10.6151
R1956 B.n767 B.n766 10.6151
R1957 B.n767 B.n535 10.6151
R1958 B.n773 B.n535 10.6151
R1959 B.n774 B.n773 10.6151
R1960 B.n775 B.n774 10.6151
R1961 B.n775 B.n533 10.6151
R1962 B.n781 B.n533 10.6151
R1963 B.n782 B.n781 10.6151
R1964 B.n783 B.n782 10.6151
R1965 B.n783 B.n531 10.6151
R1966 B.n789 B.n531 10.6151
R1967 B.n790 B.n789 10.6151
R1968 B.n791 B.n790 10.6151
R1969 B.n791 B.n529 10.6151
R1970 B.n797 B.n529 10.6151
R1971 B.n798 B.n797 10.6151
R1972 B.n799 B.n798 10.6151
R1973 B.n799 B.n527 10.6151
R1974 B.n805 B.n527 10.6151
R1975 B.n806 B.n805 10.6151
R1976 B.n807 B.n806 10.6151
R1977 B.n807 B.n525 10.6151
R1978 B.n813 B.n525 10.6151
R1979 B.n814 B.n813 10.6151
R1980 B.n815 B.n814 10.6151
R1981 B.n815 B.n523 10.6151
R1982 B.n821 B.n523 10.6151
R1983 B.n822 B.n821 10.6151
R1984 B.n823 B.n822 10.6151
R1985 B.n823 B.n521 10.6151
R1986 B.n829 B.n521 10.6151
R1987 B.n830 B.n829 10.6151
R1988 B.n831 B.n830 10.6151
R1989 B.n831 B.n519 10.6151
R1990 B.n837 B.n519 10.6151
R1991 B.n838 B.n837 10.6151
R1992 B.n844 B.n843 10.6151
R1993 B.n845 B.n844 10.6151
R1994 B.n845 B.n507 10.6151
R1995 B.n855 B.n507 10.6151
R1996 B.n856 B.n855 10.6151
R1997 B.n857 B.n856 10.6151
R1998 B.n857 B.n499 10.6151
R1999 B.n867 B.n499 10.6151
R2000 B.n868 B.n867 10.6151
R2001 B.n869 B.n868 10.6151
R2002 B.n869 B.n491 10.6151
R2003 B.n879 B.n491 10.6151
R2004 B.n880 B.n879 10.6151
R2005 B.n881 B.n880 10.6151
R2006 B.n881 B.n483 10.6151
R2007 B.n891 B.n483 10.6151
R2008 B.n892 B.n891 10.6151
R2009 B.n893 B.n892 10.6151
R2010 B.n893 B.n475 10.6151
R2011 B.n903 B.n475 10.6151
R2012 B.n904 B.n903 10.6151
R2013 B.n905 B.n904 10.6151
R2014 B.n905 B.n467 10.6151
R2015 B.n915 B.n467 10.6151
R2016 B.n916 B.n915 10.6151
R2017 B.n917 B.n916 10.6151
R2018 B.n917 B.n459 10.6151
R2019 B.n927 B.n459 10.6151
R2020 B.n928 B.n927 10.6151
R2021 B.n929 B.n928 10.6151
R2022 B.n929 B.n451 10.6151
R2023 B.n940 B.n451 10.6151
R2024 B.n941 B.n940 10.6151
R2025 B.n942 B.n941 10.6151
R2026 B.n942 B.n444 10.6151
R2027 B.n952 B.n444 10.6151
R2028 B.n953 B.n952 10.6151
R2029 B.n954 B.n953 10.6151
R2030 B.n954 B.n436 10.6151
R2031 B.n964 B.n436 10.6151
R2032 B.n965 B.n964 10.6151
R2033 B.n966 B.n965 10.6151
R2034 B.n966 B.n428 10.6151
R2035 B.n976 B.n428 10.6151
R2036 B.n977 B.n976 10.6151
R2037 B.n978 B.n977 10.6151
R2038 B.n978 B.n420 10.6151
R2039 B.n989 B.n420 10.6151
R2040 B.n990 B.n989 10.6151
R2041 B.n991 B.n990 10.6151
R2042 B.n991 B.n0 10.6151
R2043 B.n1166 B.n1 10.6151
R2044 B.n1166 B.n1165 10.6151
R2045 B.n1165 B.n1164 10.6151
R2046 B.n1164 B.n10 10.6151
R2047 B.n1158 B.n10 10.6151
R2048 B.n1158 B.n1157 10.6151
R2049 B.n1157 B.n1156 10.6151
R2050 B.n1156 B.n17 10.6151
R2051 B.n1150 B.n17 10.6151
R2052 B.n1150 B.n1149 10.6151
R2053 B.n1149 B.n1148 10.6151
R2054 B.n1148 B.n24 10.6151
R2055 B.n1142 B.n24 10.6151
R2056 B.n1142 B.n1141 10.6151
R2057 B.n1141 B.n1140 10.6151
R2058 B.n1140 B.n31 10.6151
R2059 B.n1134 B.n31 10.6151
R2060 B.n1134 B.n1133 10.6151
R2061 B.n1133 B.n1132 10.6151
R2062 B.n1132 B.n37 10.6151
R2063 B.n1126 B.n37 10.6151
R2064 B.n1126 B.n1125 10.6151
R2065 B.n1125 B.n1124 10.6151
R2066 B.n1124 B.n45 10.6151
R2067 B.n1118 B.n45 10.6151
R2068 B.n1118 B.n1117 10.6151
R2069 B.n1117 B.n1116 10.6151
R2070 B.n1116 B.n52 10.6151
R2071 B.n1110 B.n52 10.6151
R2072 B.n1110 B.n1109 10.6151
R2073 B.n1109 B.n1108 10.6151
R2074 B.n1108 B.n59 10.6151
R2075 B.n1102 B.n59 10.6151
R2076 B.n1102 B.n1101 10.6151
R2077 B.n1101 B.n1100 10.6151
R2078 B.n1100 B.n66 10.6151
R2079 B.n1094 B.n66 10.6151
R2080 B.n1094 B.n1093 10.6151
R2081 B.n1093 B.n1092 10.6151
R2082 B.n1092 B.n73 10.6151
R2083 B.n1086 B.n73 10.6151
R2084 B.n1086 B.n1085 10.6151
R2085 B.n1085 B.n1084 10.6151
R2086 B.n1084 B.n80 10.6151
R2087 B.n1078 B.n80 10.6151
R2088 B.n1078 B.n1077 10.6151
R2089 B.n1077 B.n1076 10.6151
R2090 B.n1076 B.n87 10.6151
R2091 B.n1070 B.n87 10.6151
R2092 B.n1070 B.n1069 10.6151
R2093 B.n1069 B.n1068 10.6151
R2094 B.t7 B.n497 10.0374
R2095 B.t14 B.n78 10.0374
R2096 B.n283 B.n282 6.5566
R2097 B.n299 B.n163 6.5566
R2098 B.n700 B.n699 6.5566
R2099 B.n719 B.n718 6.5566
R2100 B.n282 B.n281 4.05904
R2101 B.n302 B.n163 4.05904
R2102 B.n699 B.n698 4.05904
R2103 B.n718 B.n547 4.05904
R2104 B.t2 B.n469 3.34614
R2105 B.n944 B.t4 3.34614
R2106 B.t0 B.n426 3.34614
R2107 B.t3 B.n15 3.34614
R2108 B.n1136 B.t5 3.34614
R2109 B.n1113 B.t1 3.34614
R2110 B.n1172 B.n0 2.81026
R2111 B.n1172 B.n1 2.81026
R2112 VN.n34 VN.n33 161.3
R2113 VN.n32 VN.n19 161.3
R2114 VN.n31 VN.n30 161.3
R2115 VN.n29 VN.n20 161.3
R2116 VN.n28 VN.n27 161.3
R2117 VN.n26 VN.n21 161.3
R2118 VN.n25 VN.n24 161.3
R2119 VN.n16 VN.n15 161.3
R2120 VN.n14 VN.n1 161.3
R2121 VN.n13 VN.n12 161.3
R2122 VN.n11 VN.n2 161.3
R2123 VN.n10 VN.n9 161.3
R2124 VN.n8 VN.n3 161.3
R2125 VN.n7 VN.n6 161.3
R2126 VN.n23 VN.t4 159.168
R2127 VN.n5 VN.t3 159.168
R2128 VN.n4 VN.t0 125.377
R2129 VN.n0 VN.t2 125.377
R2130 VN.n22 VN.t5 125.377
R2131 VN.n18 VN.t1 125.377
R2132 VN.n17 VN.n0 78.4415
R2133 VN.n35 VN.n18 78.4415
R2134 VN VN.n35 56.4603
R2135 VN.n9 VN.n2 53.171
R2136 VN.n27 VN.n20 53.171
R2137 VN.n5 VN.n4 50.2542
R2138 VN.n23 VN.n22 50.2542
R2139 VN.n13 VN.n2 27.983
R2140 VN.n31 VN.n20 27.983
R2141 VN.n7 VN.n4 24.5923
R2142 VN.n8 VN.n7 24.5923
R2143 VN.n9 VN.n8 24.5923
R2144 VN.n14 VN.n13 24.5923
R2145 VN.n15 VN.n14 24.5923
R2146 VN.n27 VN.n26 24.5923
R2147 VN.n26 VN.n25 24.5923
R2148 VN.n25 VN.n22 24.5923
R2149 VN.n33 VN.n32 24.5923
R2150 VN.n32 VN.n31 24.5923
R2151 VN.n15 VN.n0 11.8046
R2152 VN.n33 VN.n18 11.8046
R2153 VN.n24 VN.n23 3.08085
R2154 VN.n6 VN.n5 3.08085
R2155 VN.n35 VN.n34 0.354861
R2156 VN.n17 VN.n16 0.354861
R2157 VN VN.n17 0.267071
R2158 VN.n34 VN.n19 0.189894
R2159 VN.n30 VN.n19 0.189894
R2160 VN.n30 VN.n29 0.189894
R2161 VN.n29 VN.n28 0.189894
R2162 VN.n28 VN.n21 0.189894
R2163 VN.n24 VN.n21 0.189894
R2164 VN.n6 VN.n3 0.189894
R2165 VN.n10 VN.n3 0.189894
R2166 VN.n11 VN.n10 0.189894
R2167 VN.n12 VN.n11 0.189894
R2168 VN.n12 VN.n1 0.189894
R2169 VN.n16 VN.n1 0.189894
R2170 VDD2.n1 VDD2.t2 67.8207
R2171 VDD2.n2 VDD2.t4 65.4589
R2172 VDD2.n1 VDD2.n0 65.0924
R2173 VDD2 VDD2.n3 65.0896
R2174 VDD2.n2 VDD2.n1 49.4868
R2175 VDD2 VDD2.n2 2.47679
R2176 VDD2.n3 VDD2.t0 1.11662
R2177 VDD2.n3 VDD2.t1 1.11662
R2178 VDD2.n0 VDD2.t5 1.11662
R2179 VDD2.n0 VDD2.t3 1.11662
C0 VN VDD1 0.152202f
C1 VDD1 VTAIL 9.87287f
C2 VN VDD2 10.2157f
C3 VDD2 VTAIL 9.92884f
C4 VDD1 VP 10.587299f
C5 VN VTAIL 10.301f
C6 VDD2 VP 0.527729f
C7 VN VP 8.772191f
C8 VDD2 VDD1 1.72363f
C9 VTAIL VP 10.3153f
C10 VDD2 B 7.610508f
C11 VDD1 B 7.975062f
C12 VTAIL B 10.674242f
C13 VN B 15.71879f
C14 VP B 14.350806f
C15 VDD2.t2 B 3.46404f
C16 VDD2.t5 B 0.295494f
C17 VDD2.t3 B 0.295494f
C18 VDD2.n0 B 2.70443f
C19 VDD2.n1 B 3.03303f
C20 VDD2.t4 B 3.45045f
C21 VDD2.n2 B 2.90351f
C22 VDD2.t0 B 0.295494f
C23 VDD2.t1 B 0.295494f
C24 VDD2.n3 B 2.70439f
C25 VN.t2 B 3.07484f
C26 VN.n0 B 1.13255f
C27 VN.n1 B 0.018485f
C28 VN.n2 B 0.019336f
C29 VN.n3 B 0.018485f
C30 VN.t0 B 3.07484f
C31 VN.n4 B 1.13412f
C32 VN.t3 B 3.32919f
C33 VN.n5 B 1.0768f
C34 VN.n6 B 0.22558f
C35 VN.n7 B 0.034278f
C36 VN.n8 B 0.034278f
C37 VN.n9 B 0.032641f
C38 VN.n10 B 0.018485f
C39 VN.n11 B 0.018485f
C40 VN.n12 B 0.018485f
C41 VN.n13 B 0.036042f
C42 VN.n14 B 0.034278f
C43 VN.n15 B 0.025478f
C44 VN.n16 B 0.029829f
C45 VN.n17 B 0.047653f
C46 VN.t1 B 3.07484f
C47 VN.n18 B 1.13255f
C48 VN.n19 B 0.018485f
C49 VN.n20 B 0.019336f
C50 VN.n21 B 0.018485f
C51 VN.t5 B 3.07484f
C52 VN.n22 B 1.13412f
C53 VN.t4 B 3.32919f
C54 VN.n23 B 1.0768f
C55 VN.n24 B 0.22558f
C56 VN.n25 B 0.034278f
C57 VN.n26 B 0.034278f
C58 VN.n27 B 0.032641f
C59 VN.n28 B 0.018485f
C60 VN.n29 B 0.018485f
C61 VN.n30 B 0.018485f
C62 VN.n31 B 0.036042f
C63 VN.n32 B 0.034278f
C64 VN.n33 B 0.025478f
C65 VN.n34 B 0.029829f
C66 VN.n35 B 1.25186f
C67 VDD1.t4 B 3.52026f
C68 VDD1.t0 B 3.51935f
C69 VDD1.t1 B 0.300212f
C70 VDD1.t5 B 0.300212f
C71 VDD1.n0 B 2.74761f
C72 VDD1.n1 B 3.21001f
C73 VDD1.t3 B 0.300212f
C74 VDD1.t2 B 0.300212f
C75 VDD1.n2 B 2.74238f
C76 VDD1.n3 B 2.94802f
C77 VTAIL.t3 B 0.320807f
C78 VTAIL.t5 B 0.320807f
C79 VTAIL.n0 B 2.86898f
C80 VTAIL.n1 B 0.427914f
C81 VTAIL.t8 B 3.66558f
C82 VTAIL.n2 B 0.68026f
C83 VTAIL.t6 B 0.320807f
C84 VTAIL.t9 B 0.320807f
C85 VTAIL.n3 B 2.86898f
C86 VTAIL.n4 B 2.36244f
C87 VTAIL.t2 B 0.320807f
C88 VTAIL.t4 B 0.320807f
C89 VTAIL.n5 B 2.86897f
C90 VTAIL.n6 B 2.36245f
C91 VTAIL.t0 B 3.66558f
C92 VTAIL.n7 B 0.680262f
C93 VTAIL.t11 B 0.320807f
C94 VTAIL.t10 B 0.320807f
C95 VTAIL.n8 B 2.86897f
C96 VTAIL.n9 B 0.601943f
C97 VTAIL.t7 B 3.66556f
C98 VTAIL.n10 B 2.20304f
C99 VTAIL.t1 B 3.66558f
C100 VTAIL.n11 B 2.1393f
C101 VP.t0 B 3.11958f
C102 VP.n0 B 1.14903f
C103 VP.n1 B 0.018754f
C104 VP.n2 B 0.019618f
C105 VP.n3 B 0.018754f
C106 VP.t4 B 3.11958f
C107 VP.n4 B 1.09455f
C108 VP.n5 B 0.018754f
C109 VP.n6 B 0.019618f
C110 VP.n7 B 0.018754f
C111 VP.t5 B 3.11958f
C112 VP.n8 B 1.14903f
C113 VP.t3 B 3.11958f
C114 VP.n9 B 1.14903f
C115 VP.n10 B 0.018754f
C116 VP.n11 B 0.019618f
C117 VP.n12 B 0.018754f
C118 VP.t2 B 3.11958f
C119 VP.n13 B 1.15062f
C120 VP.t1 B 3.37763f
C121 VP.n14 B 1.09247f
C122 VP.n15 B 0.228863f
C123 VP.n16 B 0.034777f
C124 VP.n17 B 0.034777f
C125 VP.n18 B 0.033116f
C126 VP.n19 B 0.018754f
C127 VP.n20 B 0.018754f
C128 VP.n21 B 0.018754f
C129 VP.n22 B 0.036566f
C130 VP.n23 B 0.034777f
C131 VP.n24 B 0.025849f
C132 VP.n25 B 0.030263f
C133 VP.n26 B 1.2627f
C134 VP.n27 B 1.27471f
C135 VP.n28 B 0.030263f
C136 VP.n29 B 0.025849f
C137 VP.n30 B 0.034777f
C138 VP.n31 B 0.036566f
C139 VP.n32 B 0.018754f
C140 VP.n33 B 0.018754f
C141 VP.n34 B 0.018754f
C142 VP.n35 B 0.033116f
C143 VP.n36 B 0.034777f
C144 VP.n37 B 0.034777f
C145 VP.n38 B 0.018754f
C146 VP.n39 B 0.018754f
C147 VP.n40 B 0.018754f
C148 VP.n41 B 0.034777f
C149 VP.n42 B 0.034777f
C150 VP.n43 B 0.033116f
C151 VP.n44 B 0.018754f
C152 VP.n45 B 0.018754f
C153 VP.n46 B 0.018754f
C154 VP.n47 B 0.036566f
C155 VP.n48 B 0.034777f
C156 VP.n49 B 0.025849f
C157 VP.n50 B 0.030263f
C158 VP.n51 B 0.048346f
.ends

