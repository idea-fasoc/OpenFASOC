* NGSPICE file created from diff_pair_sample_0970.ext - technology: sky130A

.subckt diff_pair_sample_0970 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=0 ps=0 w=17.95 l=1.58
X1 VDD2.t5 VN.t0 VTAIL.t11 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=7.0005 ps=36.68 w=17.95 l=1.58
X2 VTAIL.t8 VN.t1 VDD2.t4 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=2.96175 ps=18.28 w=17.95 l=1.58
X3 VDD1.t5 VP.t0 VTAIL.t4 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=2.96175 ps=18.28 w=17.95 l=1.58
X4 VDD2.t3 VN.t2 VTAIL.t6 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=2.96175 ps=18.28 w=17.95 l=1.58
X5 VDD1.t4 VP.t1 VTAIL.t5 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=7.0005 ps=36.68 w=17.95 l=1.58
X6 VDD1.t3 VP.t2 VTAIL.t0 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=2.96175 ps=18.28 w=17.95 l=1.58
X7 VDD2.t2 VN.t3 VTAIL.t9 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=7.0005 ps=36.68 w=17.95 l=1.58
X8 VDD1.t2 VP.t3 VTAIL.t2 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=7.0005 ps=36.68 w=17.95 l=1.58
X9 B.t8 B.t6 B.t7 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=0 ps=0 w=17.95 l=1.58
X10 B.t5 B.t3 B.t4 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=0 ps=0 w=17.95 l=1.58
X11 B.t2 B.t0 B.t1 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=0 ps=0 w=17.95 l=1.58
X12 VDD2.t1 VN.t4 VTAIL.t10 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=7.0005 pd=36.68 as=2.96175 ps=18.28 w=17.95 l=1.58
X13 VTAIL.t7 VN.t5 VDD2.t0 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=2.96175 ps=18.28 w=17.95 l=1.58
X14 VTAIL.t3 VP.t4 VDD1.t1 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=2.96175 ps=18.28 w=17.95 l=1.58
X15 VTAIL.t1 VP.t5 VDD1.t0 w_n2498_n4558# sky130_fd_pr__pfet_01v8 ad=2.96175 pd=18.28 as=2.96175 ps=18.28 w=17.95 l=1.58
R0 B.n436 B.n117 585
R1 B.n435 B.n434 585
R2 B.n433 B.n118 585
R3 B.n432 B.n431 585
R4 B.n430 B.n119 585
R5 B.n429 B.n428 585
R6 B.n427 B.n120 585
R7 B.n426 B.n425 585
R8 B.n424 B.n121 585
R9 B.n423 B.n422 585
R10 B.n421 B.n122 585
R11 B.n420 B.n419 585
R12 B.n418 B.n123 585
R13 B.n417 B.n416 585
R14 B.n415 B.n124 585
R15 B.n414 B.n413 585
R16 B.n412 B.n125 585
R17 B.n411 B.n410 585
R18 B.n409 B.n126 585
R19 B.n408 B.n407 585
R20 B.n406 B.n127 585
R21 B.n405 B.n404 585
R22 B.n403 B.n128 585
R23 B.n402 B.n401 585
R24 B.n400 B.n129 585
R25 B.n399 B.n398 585
R26 B.n397 B.n130 585
R27 B.n396 B.n395 585
R28 B.n394 B.n131 585
R29 B.n393 B.n392 585
R30 B.n391 B.n132 585
R31 B.n390 B.n389 585
R32 B.n388 B.n133 585
R33 B.n387 B.n386 585
R34 B.n385 B.n134 585
R35 B.n384 B.n383 585
R36 B.n382 B.n135 585
R37 B.n381 B.n380 585
R38 B.n379 B.n136 585
R39 B.n378 B.n377 585
R40 B.n376 B.n137 585
R41 B.n375 B.n374 585
R42 B.n373 B.n138 585
R43 B.n372 B.n371 585
R44 B.n370 B.n139 585
R45 B.n369 B.n368 585
R46 B.n367 B.n140 585
R47 B.n366 B.n365 585
R48 B.n364 B.n141 585
R49 B.n363 B.n362 585
R50 B.n361 B.n142 585
R51 B.n360 B.n359 585
R52 B.n358 B.n143 585
R53 B.n357 B.n356 585
R54 B.n355 B.n144 585
R55 B.n354 B.n353 585
R56 B.n352 B.n145 585
R57 B.n351 B.n350 585
R58 B.n349 B.n146 585
R59 B.n347 B.n346 585
R60 B.n345 B.n149 585
R61 B.n344 B.n343 585
R62 B.n342 B.n150 585
R63 B.n341 B.n340 585
R64 B.n339 B.n151 585
R65 B.n338 B.n337 585
R66 B.n336 B.n152 585
R67 B.n335 B.n334 585
R68 B.n333 B.n153 585
R69 B.n332 B.n331 585
R70 B.n327 B.n154 585
R71 B.n326 B.n325 585
R72 B.n324 B.n155 585
R73 B.n323 B.n322 585
R74 B.n321 B.n156 585
R75 B.n320 B.n319 585
R76 B.n318 B.n157 585
R77 B.n317 B.n316 585
R78 B.n315 B.n158 585
R79 B.n314 B.n313 585
R80 B.n312 B.n159 585
R81 B.n311 B.n310 585
R82 B.n309 B.n160 585
R83 B.n308 B.n307 585
R84 B.n306 B.n161 585
R85 B.n305 B.n304 585
R86 B.n303 B.n162 585
R87 B.n302 B.n301 585
R88 B.n300 B.n163 585
R89 B.n299 B.n298 585
R90 B.n297 B.n164 585
R91 B.n296 B.n295 585
R92 B.n294 B.n165 585
R93 B.n293 B.n292 585
R94 B.n291 B.n166 585
R95 B.n290 B.n289 585
R96 B.n288 B.n167 585
R97 B.n287 B.n286 585
R98 B.n285 B.n168 585
R99 B.n284 B.n283 585
R100 B.n282 B.n169 585
R101 B.n281 B.n280 585
R102 B.n279 B.n170 585
R103 B.n278 B.n277 585
R104 B.n276 B.n171 585
R105 B.n275 B.n274 585
R106 B.n273 B.n172 585
R107 B.n272 B.n271 585
R108 B.n270 B.n173 585
R109 B.n269 B.n268 585
R110 B.n267 B.n174 585
R111 B.n266 B.n265 585
R112 B.n264 B.n175 585
R113 B.n263 B.n262 585
R114 B.n261 B.n176 585
R115 B.n260 B.n259 585
R116 B.n258 B.n177 585
R117 B.n257 B.n256 585
R118 B.n255 B.n178 585
R119 B.n254 B.n253 585
R120 B.n252 B.n179 585
R121 B.n251 B.n250 585
R122 B.n249 B.n180 585
R123 B.n248 B.n247 585
R124 B.n246 B.n181 585
R125 B.n245 B.n244 585
R126 B.n243 B.n182 585
R127 B.n242 B.n241 585
R128 B.n438 B.n437 585
R129 B.n439 B.n116 585
R130 B.n441 B.n440 585
R131 B.n442 B.n115 585
R132 B.n444 B.n443 585
R133 B.n445 B.n114 585
R134 B.n447 B.n446 585
R135 B.n448 B.n113 585
R136 B.n450 B.n449 585
R137 B.n451 B.n112 585
R138 B.n453 B.n452 585
R139 B.n454 B.n111 585
R140 B.n456 B.n455 585
R141 B.n457 B.n110 585
R142 B.n459 B.n458 585
R143 B.n460 B.n109 585
R144 B.n462 B.n461 585
R145 B.n463 B.n108 585
R146 B.n465 B.n464 585
R147 B.n466 B.n107 585
R148 B.n468 B.n467 585
R149 B.n469 B.n106 585
R150 B.n471 B.n470 585
R151 B.n472 B.n105 585
R152 B.n474 B.n473 585
R153 B.n475 B.n104 585
R154 B.n477 B.n476 585
R155 B.n478 B.n103 585
R156 B.n480 B.n479 585
R157 B.n481 B.n102 585
R158 B.n483 B.n482 585
R159 B.n484 B.n101 585
R160 B.n486 B.n485 585
R161 B.n487 B.n100 585
R162 B.n489 B.n488 585
R163 B.n490 B.n99 585
R164 B.n492 B.n491 585
R165 B.n493 B.n98 585
R166 B.n495 B.n494 585
R167 B.n496 B.n97 585
R168 B.n498 B.n497 585
R169 B.n499 B.n96 585
R170 B.n501 B.n500 585
R171 B.n502 B.n95 585
R172 B.n504 B.n503 585
R173 B.n505 B.n94 585
R174 B.n507 B.n506 585
R175 B.n508 B.n93 585
R176 B.n510 B.n509 585
R177 B.n511 B.n92 585
R178 B.n513 B.n512 585
R179 B.n514 B.n91 585
R180 B.n516 B.n515 585
R181 B.n517 B.n90 585
R182 B.n519 B.n518 585
R183 B.n520 B.n89 585
R184 B.n522 B.n521 585
R185 B.n523 B.n88 585
R186 B.n525 B.n524 585
R187 B.n526 B.n87 585
R188 B.n528 B.n527 585
R189 B.n529 B.n86 585
R190 B.n722 B.n17 585
R191 B.n721 B.n720 585
R192 B.n719 B.n18 585
R193 B.n718 B.n717 585
R194 B.n716 B.n19 585
R195 B.n715 B.n714 585
R196 B.n713 B.n20 585
R197 B.n712 B.n711 585
R198 B.n710 B.n21 585
R199 B.n709 B.n708 585
R200 B.n707 B.n22 585
R201 B.n706 B.n705 585
R202 B.n704 B.n23 585
R203 B.n703 B.n702 585
R204 B.n701 B.n24 585
R205 B.n700 B.n699 585
R206 B.n698 B.n25 585
R207 B.n697 B.n696 585
R208 B.n695 B.n26 585
R209 B.n694 B.n693 585
R210 B.n692 B.n27 585
R211 B.n691 B.n690 585
R212 B.n689 B.n28 585
R213 B.n688 B.n687 585
R214 B.n686 B.n29 585
R215 B.n685 B.n684 585
R216 B.n683 B.n30 585
R217 B.n682 B.n681 585
R218 B.n680 B.n31 585
R219 B.n679 B.n678 585
R220 B.n677 B.n32 585
R221 B.n676 B.n675 585
R222 B.n674 B.n33 585
R223 B.n673 B.n672 585
R224 B.n671 B.n34 585
R225 B.n670 B.n669 585
R226 B.n668 B.n35 585
R227 B.n667 B.n666 585
R228 B.n665 B.n36 585
R229 B.n664 B.n663 585
R230 B.n662 B.n37 585
R231 B.n661 B.n660 585
R232 B.n659 B.n38 585
R233 B.n658 B.n657 585
R234 B.n656 B.n39 585
R235 B.n655 B.n654 585
R236 B.n653 B.n40 585
R237 B.n652 B.n651 585
R238 B.n650 B.n41 585
R239 B.n649 B.n648 585
R240 B.n647 B.n42 585
R241 B.n646 B.n645 585
R242 B.n644 B.n43 585
R243 B.n643 B.n642 585
R244 B.n641 B.n44 585
R245 B.n640 B.n639 585
R246 B.n638 B.n45 585
R247 B.n637 B.n636 585
R248 B.n635 B.n46 585
R249 B.n634 B.n633 585
R250 B.n632 B.n47 585
R251 B.n631 B.n630 585
R252 B.n629 B.n51 585
R253 B.n628 B.n627 585
R254 B.n626 B.n52 585
R255 B.n625 B.n624 585
R256 B.n623 B.n53 585
R257 B.n622 B.n621 585
R258 B.n620 B.n54 585
R259 B.n618 B.n617 585
R260 B.n616 B.n57 585
R261 B.n615 B.n614 585
R262 B.n613 B.n58 585
R263 B.n612 B.n611 585
R264 B.n610 B.n59 585
R265 B.n609 B.n608 585
R266 B.n607 B.n60 585
R267 B.n606 B.n605 585
R268 B.n604 B.n61 585
R269 B.n603 B.n602 585
R270 B.n601 B.n62 585
R271 B.n600 B.n599 585
R272 B.n598 B.n63 585
R273 B.n597 B.n596 585
R274 B.n595 B.n64 585
R275 B.n594 B.n593 585
R276 B.n592 B.n65 585
R277 B.n591 B.n590 585
R278 B.n589 B.n66 585
R279 B.n588 B.n587 585
R280 B.n586 B.n67 585
R281 B.n585 B.n584 585
R282 B.n583 B.n68 585
R283 B.n582 B.n581 585
R284 B.n580 B.n69 585
R285 B.n579 B.n578 585
R286 B.n577 B.n70 585
R287 B.n576 B.n575 585
R288 B.n574 B.n71 585
R289 B.n573 B.n572 585
R290 B.n571 B.n72 585
R291 B.n570 B.n569 585
R292 B.n568 B.n73 585
R293 B.n567 B.n566 585
R294 B.n565 B.n74 585
R295 B.n564 B.n563 585
R296 B.n562 B.n75 585
R297 B.n561 B.n560 585
R298 B.n559 B.n76 585
R299 B.n558 B.n557 585
R300 B.n556 B.n77 585
R301 B.n555 B.n554 585
R302 B.n553 B.n78 585
R303 B.n552 B.n551 585
R304 B.n550 B.n79 585
R305 B.n549 B.n548 585
R306 B.n547 B.n80 585
R307 B.n546 B.n545 585
R308 B.n544 B.n81 585
R309 B.n543 B.n542 585
R310 B.n541 B.n82 585
R311 B.n540 B.n539 585
R312 B.n538 B.n83 585
R313 B.n537 B.n536 585
R314 B.n535 B.n84 585
R315 B.n534 B.n533 585
R316 B.n532 B.n85 585
R317 B.n531 B.n530 585
R318 B.n724 B.n723 585
R319 B.n725 B.n16 585
R320 B.n727 B.n726 585
R321 B.n728 B.n15 585
R322 B.n730 B.n729 585
R323 B.n731 B.n14 585
R324 B.n733 B.n732 585
R325 B.n734 B.n13 585
R326 B.n736 B.n735 585
R327 B.n737 B.n12 585
R328 B.n739 B.n738 585
R329 B.n740 B.n11 585
R330 B.n742 B.n741 585
R331 B.n743 B.n10 585
R332 B.n745 B.n744 585
R333 B.n746 B.n9 585
R334 B.n748 B.n747 585
R335 B.n749 B.n8 585
R336 B.n751 B.n750 585
R337 B.n752 B.n7 585
R338 B.n754 B.n753 585
R339 B.n755 B.n6 585
R340 B.n757 B.n756 585
R341 B.n758 B.n5 585
R342 B.n760 B.n759 585
R343 B.n761 B.n4 585
R344 B.n763 B.n762 585
R345 B.n764 B.n3 585
R346 B.n766 B.n765 585
R347 B.n767 B.n0 585
R348 B.n2 B.n1 585
R349 B.n198 B.n197 585
R350 B.n200 B.n199 585
R351 B.n201 B.n196 585
R352 B.n203 B.n202 585
R353 B.n204 B.n195 585
R354 B.n206 B.n205 585
R355 B.n207 B.n194 585
R356 B.n209 B.n208 585
R357 B.n210 B.n193 585
R358 B.n212 B.n211 585
R359 B.n213 B.n192 585
R360 B.n215 B.n214 585
R361 B.n216 B.n191 585
R362 B.n218 B.n217 585
R363 B.n219 B.n190 585
R364 B.n221 B.n220 585
R365 B.n222 B.n189 585
R366 B.n224 B.n223 585
R367 B.n225 B.n188 585
R368 B.n227 B.n226 585
R369 B.n228 B.n187 585
R370 B.n230 B.n229 585
R371 B.n231 B.n186 585
R372 B.n233 B.n232 585
R373 B.n234 B.n185 585
R374 B.n236 B.n235 585
R375 B.n237 B.n184 585
R376 B.n239 B.n238 585
R377 B.n240 B.n183 585
R378 B.n241 B.n240 497.305
R379 B.n437 B.n436 497.305
R380 B.n531 B.n86 497.305
R381 B.n724 B.n17 497.305
R382 B.n328 B.t0 479.521
R383 B.n147 B.t6 479.521
R384 B.n55 B.t3 479.521
R385 B.n48 B.t9 479.521
R386 B.n769 B.n768 256.663
R387 B.n768 B.n767 235.042
R388 B.n768 B.n2 235.042
R389 B.n241 B.n182 163.367
R390 B.n245 B.n182 163.367
R391 B.n246 B.n245 163.367
R392 B.n247 B.n246 163.367
R393 B.n247 B.n180 163.367
R394 B.n251 B.n180 163.367
R395 B.n252 B.n251 163.367
R396 B.n253 B.n252 163.367
R397 B.n253 B.n178 163.367
R398 B.n257 B.n178 163.367
R399 B.n258 B.n257 163.367
R400 B.n259 B.n258 163.367
R401 B.n259 B.n176 163.367
R402 B.n263 B.n176 163.367
R403 B.n264 B.n263 163.367
R404 B.n265 B.n264 163.367
R405 B.n265 B.n174 163.367
R406 B.n269 B.n174 163.367
R407 B.n270 B.n269 163.367
R408 B.n271 B.n270 163.367
R409 B.n271 B.n172 163.367
R410 B.n275 B.n172 163.367
R411 B.n276 B.n275 163.367
R412 B.n277 B.n276 163.367
R413 B.n277 B.n170 163.367
R414 B.n281 B.n170 163.367
R415 B.n282 B.n281 163.367
R416 B.n283 B.n282 163.367
R417 B.n283 B.n168 163.367
R418 B.n287 B.n168 163.367
R419 B.n288 B.n287 163.367
R420 B.n289 B.n288 163.367
R421 B.n289 B.n166 163.367
R422 B.n293 B.n166 163.367
R423 B.n294 B.n293 163.367
R424 B.n295 B.n294 163.367
R425 B.n295 B.n164 163.367
R426 B.n299 B.n164 163.367
R427 B.n300 B.n299 163.367
R428 B.n301 B.n300 163.367
R429 B.n301 B.n162 163.367
R430 B.n305 B.n162 163.367
R431 B.n306 B.n305 163.367
R432 B.n307 B.n306 163.367
R433 B.n307 B.n160 163.367
R434 B.n311 B.n160 163.367
R435 B.n312 B.n311 163.367
R436 B.n313 B.n312 163.367
R437 B.n313 B.n158 163.367
R438 B.n317 B.n158 163.367
R439 B.n318 B.n317 163.367
R440 B.n319 B.n318 163.367
R441 B.n319 B.n156 163.367
R442 B.n323 B.n156 163.367
R443 B.n324 B.n323 163.367
R444 B.n325 B.n324 163.367
R445 B.n325 B.n154 163.367
R446 B.n332 B.n154 163.367
R447 B.n333 B.n332 163.367
R448 B.n334 B.n333 163.367
R449 B.n334 B.n152 163.367
R450 B.n338 B.n152 163.367
R451 B.n339 B.n338 163.367
R452 B.n340 B.n339 163.367
R453 B.n340 B.n150 163.367
R454 B.n344 B.n150 163.367
R455 B.n345 B.n344 163.367
R456 B.n346 B.n345 163.367
R457 B.n346 B.n146 163.367
R458 B.n351 B.n146 163.367
R459 B.n352 B.n351 163.367
R460 B.n353 B.n352 163.367
R461 B.n353 B.n144 163.367
R462 B.n357 B.n144 163.367
R463 B.n358 B.n357 163.367
R464 B.n359 B.n358 163.367
R465 B.n359 B.n142 163.367
R466 B.n363 B.n142 163.367
R467 B.n364 B.n363 163.367
R468 B.n365 B.n364 163.367
R469 B.n365 B.n140 163.367
R470 B.n369 B.n140 163.367
R471 B.n370 B.n369 163.367
R472 B.n371 B.n370 163.367
R473 B.n371 B.n138 163.367
R474 B.n375 B.n138 163.367
R475 B.n376 B.n375 163.367
R476 B.n377 B.n376 163.367
R477 B.n377 B.n136 163.367
R478 B.n381 B.n136 163.367
R479 B.n382 B.n381 163.367
R480 B.n383 B.n382 163.367
R481 B.n383 B.n134 163.367
R482 B.n387 B.n134 163.367
R483 B.n388 B.n387 163.367
R484 B.n389 B.n388 163.367
R485 B.n389 B.n132 163.367
R486 B.n393 B.n132 163.367
R487 B.n394 B.n393 163.367
R488 B.n395 B.n394 163.367
R489 B.n395 B.n130 163.367
R490 B.n399 B.n130 163.367
R491 B.n400 B.n399 163.367
R492 B.n401 B.n400 163.367
R493 B.n401 B.n128 163.367
R494 B.n405 B.n128 163.367
R495 B.n406 B.n405 163.367
R496 B.n407 B.n406 163.367
R497 B.n407 B.n126 163.367
R498 B.n411 B.n126 163.367
R499 B.n412 B.n411 163.367
R500 B.n413 B.n412 163.367
R501 B.n413 B.n124 163.367
R502 B.n417 B.n124 163.367
R503 B.n418 B.n417 163.367
R504 B.n419 B.n418 163.367
R505 B.n419 B.n122 163.367
R506 B.n423 B.n122 163.367
R507 B.n424 B.n423 163.367
R508 B.n425 B.n424 163.367
R509 B.n425 B.n120 163.367
R510 B.n429 B.n120 163.367
R511 B.n430 B.n429 163.367
R512 B.n431 B.n430 163.367
R513 B.n431 B.n118 163.367
R514 B.n435 B.n118 163.367
R515 B.n436 B.n435 163.367
R516 B.n527 B.n86 163.367
R517 B.n527 B.n526 163.367
R518 B.n526 B.n525 163.367
R519 B.n525 B.n88 163.367
R520 B.n521 B.n88 163.367
R521 B.n521 B.n520 163.367
R522 B.n520 B.n519 163.367
R523 B.n519 B.n90 163.367
R524 B.n515 B.n90 163.367
R525 B.n515 B.n514 163.367
R526 B.n514 B.n513 163.367
R527 B.n513 B.n92 163.367
R528 B.n509 B.n92 163.367
R529 B.n509 B.n508 163.367
R530 B.n508 B.n507 163.367
R531 B.n507 B.n94 163.367
R532 B.n503 B.n94 163.367
R533 B.n503 B.n502 163.367
R534 B.n502 B.n501 163.367
R535 B.n501 B.n96 163.367
R536 B.n497 B.n96 163.367
R537 B.n497 B.n496 163.367
R538 B.n496 B.n495 163.367
R539 B.n495 B.n98 163.367
R540 B.n491 B.n98 163.367
R541 B.n491 B.n490 163.367
R542 B.n490 B.n489 163.367
R543 B.n489 B.n100 163.367
R544 B.n485 B.n100 163.367
R545 B.n485 B.n484 163.367
R546 B.n484 B.n483 163.367
R547 B.n483 B.n102 163.367
R548 B.n479 B.n102 163.367
R549 B.n479 B.n478 163.367
R550 B.n478 B.n477 163.367
R551 B.n477 B.n104 163.367
R552 B.n473 B.n104 163.367
R553 B.n473 B.n472 163.367
R554 B.n472 B.n471 163.367
R555 B.n471 B.n106 163.367
R556 B.n467 B.n106 163.367
R557 B.n467 B.n466 163.367
R558 B.n466 B.n465 163.367
R559 B.n465 B.n108 163.367
R560 B.n461 B.n108 163.367
R561 B.n461 B.n460 163.367
R562 B.n460 B.n459 163.367
R563 B.n459 B.n110 163.367
R564 B.n455 B.n110 163.367
R565 B.n455 B.n454 163.367
R566 B.n454 B.n453 163.367
R567 B.n453 B.n112 163.367
R568 B.n449 B.n112 163.367
R569 B.n449 B.n448 163.367
R570 B.n448 B.n447 163.367
R571 B.n447 B.n114 163.367
R572 B.n443 B.n114 163.367
R573 B.n443 B.n442 163.367
R574 B.n442 B.n441 163.367
R575 B.n441 B.n116 163.367
R576 B.n437 B.n116 163.367
R577 B.n720 B.n17 163.367
R578 B.n720 B.n719 163.367
R579 B.n719 B.n718 163.367
R580 B.n718 B.n19 163.367
R581 B.n714 B.n19 163.367
R582 B.n714 B.n713 163.367
R583 B.n713 B.n712 163.367
R584 B.n712 B.n21 163.367
R585 B.n708 B.n21 163.367
R586 B.n708 B.n707 163.367
R587 B.n707 B.n706 163.367
R588 B.n706 B.n23 163.367
R589 B.n702 B.n23 163.367
R590 B.n702 B.n701 163.367
R591 B.n701 B.n700 163.367
R592 B.n700 B.n25 163.367
R593 B.n696 B.n25 163.367
R594 B.n696 B.n695 163.367
R595 B.n695 B.n694 163.367
R596 B.n694 B.n27 163.367
R597 B.n690 B.n27 163.367
R598 B.n690 B.n689 163.367
R599 B.n689 B.n688 163.367
R600 B.n688 B.n29 163.367
R601 B.n684 B.n29 163.367
R602 B.n684 B.n683 163.367
R603 B.n683 B.n682 163.367
R604 B.n682 B.n31 163.367
R605 B.n678 B.n31 163.367
R606 B.n678 B.n677 163.367
R607 B.n677 B.n676 163.367
R608 B.n676 B.n33 163.367
R609 B.n672 B.n33 163.367
R610 B.n672 B.n671 163.367
R611 B.n671 B.n670 163.367
R612 B.n670 B.n35 163.367
R613 B.n666 B.n35 163.367
R614 B.n666 B.n665 163.367
R615 B.n665 B.n664 163.367
R616 B.n664 B.n37 163.367
R617 B.n660 B.n37 163.367
R618 B.n660 B.n659 163.367
R619 B.n659 B.n658 163.367
R620 B.n658 B.n39 163.367
R621 B.n654 B.n39 163.367
R622 B.n654 B.n653 163.367
R623 B.n653 B.n652 163.367
R624 B.n652 B.n41 163.367
R625 B.n648 B.n41 163.367
R626 B.n648 B.n647 163.367
R627 B.n647 B.n646 163.367
R628 B.n646 B.n43 163.367
R629 B.n642 B.n43 163.367
R630 B.n642 B.n641 163.367
R631 B.n641 B.n640 163.367
R632 B.n640 B.n45 163.367
R633 B.n636 B.n45 163.367
R634 B.n636 B.n635 163.367
R635 B.n635 B.n634 163.367
R636 B.n634 B.n47 163.367
R637 B.n630 B.n47 163.367
R638 B.n630 B.n629 163.367
R639 B.n629 B.n628 163.367
R640 B.n628 B.n52 163.367
R641 B.n624 B.n52 163.367
R642 B.n624 B.n623 163.367
R643 B.n623 B.n622 163.367
R644 B.n622 B.n54 163.367
R645 B.n617 B.n54 163.367
R646 B.n617 B.n616 163.367
R647 B.n616 B.n615 163.367
R648 B.n615 B.n58 163.367
R649 B.n611 B.n58 163.367
R650 B.n611 B.n610 163.367
R651 B.n610 B.n609 163.367
R652 B.n609 B.n60 163.367
R653 B.n605 B.n60 163.367
R654 B.n605 B.n604 163.367
R655 B.n604 B.n603 163.367
R656 B.n603 B.n62 163.367
R657 B.n599 B.n62 163.367
R658 B.n599 B.n598 163.367
R659 B.n598 B.n597 163.367
R660 B.n597 B.n64 163.367
R661 B.n593 B.n64 163.367
R662 B.n593 B.n592 163.367
R663 B.n592 B.n591 163.367
R664 B.n591 B.n66 163.367
R665 B.n587 B.n66 163.367
R666 B.n587 B.n586 163.367
R667 B.n586 B.n585 163.367
R668 B.n585 B.n68 163.367
R669 B.n581 B.n68 163.367
R670 B.n581 B.n580 163.367
R671 B.n580 B.n579 163.367
R672 B.n579 B.n70 163.367
R673 B.n575 B.n70 163.367
R674 B.n575 B.n574 163.367
R675 B.n574 B.n573 163.367
R676 B.n573 B.n72 163.367
R677 B.n569 B.n72 163.367
R678 B.n569 B.n568 163.367
R679 B.n568 B.n567 163.367
R680 B.n567 B.n74 163.367
R681 B.n563 B.n74 163.367
R682 B.n563 B.n562 163.367
R683 B.n562 B.n561 163.367
R684 B.n561 B.n76 163.367
R685 B.n557 B.n76 163.367
R686 B.n557 B.n556 163.367
R687 B.n556 B.n555 163.367
R688 B.n555 B.n78 163.367
R689 B.n551 B.n78 163.367
R690 B.n551 B.n550 163.367
R691 B.n550 B.n549 163.367
R692 B.n549 B.n80 163.367
R693 B.n545 B.n80 163.367
R694 B.n545 B.n544 163.367
R695 B.n544 B.n543 163.367
R696 B.n543 B.n82 163.367
R697 B.n539 B.n82 163.367
R698 B.n539 B.n538 163.367
R699 B.n538 B.n537 163.367
R700 B.n537 B.n84 163.367
R701 B.n533 B.n84 163.367
R702 B.n533 B.n532 163.367
R703 B.n532 B.n531 163.367
R704 B.n725 B.n724 163.367
R705 B.n726 B.n725 163.367
R706 B.n726 B.n15 163.367
R707 B.n730 B.n15 163.367
R708 B.n731 B.n730 163.367
R709 B.n732 B.n731 163.367
R710 B.n732 B.n13 163.367
R711 B.n736 B.n13 163.367
R712 B.n737 B.n736 163.367
R713 B.n738 B.n737 163.367
R714 B.n738 B.n11 163.367
R715 B.n742 B.n11 163.367
R716 B.n743 B.n742 163.367
R717 B.n744 B.n743 163.367
R718 B.n744 B.n9 163.367
R719 B.n748 B.n9 163.367
R720 B.n749 B.n748 163.367
R721 B.n750 B.n749 163.367
R722 B.n750 B.n7 163.367
R723 B.n754 B.n7 163.367
R724 B.n755 B.n754 163.367
R725 B.n756 B.n755 163.367
R726 B.n756 B.n5 163.367
R727 B.n760 B.n5 163.367
R728 B.n761 B.n760 163.367
R729 B.n762 B.n761 163.367
R730 B.n762 B.n3 163.367
R731 B.n766 B.n3 163.367
R732 B.n767 B.n766 163.367
R733 B.n198 B.n2 163.367
R734 B.n199 B.n198 163.367
R735 B.n199 B.n196 163.367
R736 B.n203 B.n196 163.367
R737 B.n204 B.n203 163.367
R738 B.n205 B.n204 163.367
R739 B.n205 B.n194 163.367
R740 B.n209 B.n194 163.367
R741 B.n210 B.n209 163.367
R742 B.n211 B.n210 163.367
R743 B.n211 B.n192 163.367
R744 B.n215 B.n192 163.367
R745 B.n216 B.n215 163.367
R746 B.n217 B.n216 163.367
R747 B.n217 B.n190 163.367
R748 B.n221 B.n190 163.367
R749 B.n222 B.n221 163.367
R750 B.n223 B.n222 163.367
R751 B.n223 B.n188 163.367
R752 B.n227 B.n188 163.367
R753 B.n228 B.n227 163.367
R754 B.n229 B.n228 163.367
R755 B.n229 B.n186 163.367
R756 B.n233 B.n186 163.367
R757 B.n234 B.n233 163.367
R758 B.n235 B.n234 163.367
R759 B.n235 B.n184 163.367
R760 B.n239 B.n184 163.367
R761 B.n240 B.n239 163.367
R762 B.n147 B.t7 148.488
R763 B.n55 B.t5 148.488
R764 B.n328 B.t1 148.464
R765 B.n48 B.t11 148.464
R766 B.n148 B.t8 111.445
R767 B.n56 B.t4 111.445
R768 B.n329 B.t2 111.422
R769 B.n49 B.t10 111.422
R770 B.n330 B.n329 59.5399
R771 B.n348 B.n148 59.5399
R772 B.n619 B.n56 59.5399
R773 B.n50 B.n49 59.5399
R774 B.n329 B.n328 37.0429
R775 B.n148 B.n147 37.0429
R776 B.n56 B.n55 37.0429
R777 B.n49 B.n48 37.0429
R778 B.n723 B.n722 32.3127
R779 B.n530 B.n529 32.3127
R780 B.n438 B.n117 32.3127
R781 B.n242 B.n183 32.3127
R782 B B.n769 18.0485
R783 B.n723 B.n16 10.6151
R784 B.n727 B.n16 10.6151
R785 B.n728 B.n727 10.6151
R786 B.n729 B.n728 10.6151
R787 B.n729 B.n14 10.6151
R788 B.n733 B.n14 10.6151
R789 B.n734 B.n733 10.6151
R790 B.n735 B.n734 10.6151
R791 B.n735 B.n12 10.6151
R792 B.n739 B.n12 10.6151
R793 B.n740 B.n739 10.6151
R794 B.n741 B.n740 10.6151
R795 B.n741 B.n10 10.6151
R796 B.n745 B.n10 10.6151
R797 B.n746 B.n745 10.6151
R798 B.n747 B.n746 10.6151
R799 B.n747 B.n8 10.6151
R800 B.n751 B.n8 10.6151
R801 B.n752 B.n751 10.6151
R802 B.n753 B.n752 10.6151
R803 B.n753 B.n6 10.6151
R804 B.n757 B.n6 10.6151
R805 B.n758 B.n757 10.6151
R806 B.n759 B.n758 10.6151
R807 B.n759 B.n4 10.6151
R808 B.n763 B.n4 10.6151
R809 B.n764 B.n763 10.6151
R810 B.n765 B.n764 10.6151
R811 B.n765 B.n0 10.6151
R812 B.n722 B.n721 10.6151
R813 B.n721 B.n18 10.6151
R814 B.n717 B.n18 10.6151
R815 B.n717 B.n716 10.6151
R816 B.n716 B.n715 10.6151
R817 B.n715 B.n20 10.6151
R818 B.n711 B.n20 10.6151
R819 B.n711 B.n710 10.6151
R820 B.n710 B.n709 10.6151
R821 B.n709 B.n22 10.6151
R822 B.n705 B.n22 10.6151
R823 B.n705 B.n704 10.6151
R824 B.n704 B.n703 10.6151
R825 B.n703 B.n24 10.6151
R826 B.n699 B.n24 10.6151
R827 B.n699 B.n698 10.6151
R828 B.n698 B.n697 10.6151
R829 B.n697 B.n26 10.6151
R830 B.n693 B.n26 10.6151
R831 B.n693 B.n692 10.6151
R832 B.n692 B.n691 10.6151
R833 B.n691 B.n28 10.6151
R834 B.n687 B.n28 10.6151
R835 B.n687 B.n686 10.6151
R836 B.n686 B.n685 10.6151
R837 B.n685 B.n30 10.6151
R838 B.n681 B.n30 10.6151
R839 B.n681 B.n680 10.6151
R840 B.n680 B.n679 10.6151
R841 B.n679 B.n32 10.6151
R842 B.n675 B.n32 10.6151
R843 B.n675 B.n674 10.6151
R844 B.n674 B.n673 10.6151
R845 B.n673 B.n34 10.6151
R846 B.n669 B.n34 10.6151
R847 B.n669 B.n668 10.6151
R848 B.n668 B.n667 10.6151
R849 B.n667 B.n36 10.6151
R850 B.n663 B.n36 10.6151
R851 B.n663 B.n662 10.6151
R852 B.n662 B.n661 10.6151
R853 B.n661 B.n38 10.6151
R854 B.n657 B.n38 10.6151
R855 B.n657 B.n656 10.6151
R856 B.n656 B.n655 10.6151
R857 B.n655 B.n40 10.6151
R858 B.n651 B.n40 10.6151
R859 B.n651 B.n650 10.6151
R860 B.n650 B.n649 10.6151
R861 B.n649 B.n42 10.6151
R862 B.n645 B.n42 10.6151
R863 B.n645 B.n644 10.6151
R864 B.n644 B.n643 10.6151
R865 B.n643 B.n44 10.6151
R866 B.n639 B.n44 10.6151
R867 B.n639 B.n638 10.6151
R868 B.n638 B.n637 10.6151
R869 B.n637 B.n46 10.6151
R870 B.n633 B.n632 10.6151
R871 B.n632 B.n631 10.6151
R872 B.n631 B.n51 10.6151
R873 B.n627 B.n51 10.6151
R874 B.n627 B.n626 10.6151
R875 B.n626 B.n625 10.6151
R876 B.n625 B.n53 10.6151
R877 B.n621 B.n53 10.6151
R878 B.n621 B.n620 10.6151
R879 B.n618 B.n57 10.6151
R880 B.n614 B.n57 10.6151
R881 B.n614 B.n613 10.6151
R882 B.n613 B.n612 10.6151
R883 B.n612 B.n59 10.6151
R884 B.n608 B.n59 10.6151
R885 B.n608 B.n607 10.6151
R886 B.n607 B.n606 10.6151
R887 B.n606 B.n61 10.6151
R888 B.n602 B.n61 10.6151
R889 B.n602 B.n601 10.6151
R890 B.n601 B.n600 10.6151
R891 B.n600 B.n63 10.6151
R892 B.n596 B.n63 10.6151
R893 B.n596 B.n595 10.6151
R894 B.n595 B.n594 10.6151
R895 B.n594 B.n65 10.6151
R896 B.n590 B.n65 10.6151
R897 B.n590 B.n589 10.6151
R898 B.n589 B.n588 10.6151
R899 B.n588 B.n67 10.6151
R900 B.n584 B.n67 10.6151
R901 B.n584 B.n583 10.6151
R902 B.n583 B.n582 10.6151
R903 B.n582 B.n69 10.6151
R904 B.n578 B.n69 10.6151
R905 B.n578 B.n577 10.6151
R906 B.n577 B.n576 10.6151
R907 B.n576 B.n71 10.6151
R908 B.n572 B.n71 10.6151
R909 B.n572 B.n571 10.6151
R910 B.n571 B.n570 10.6151
R911 B.n570 B.n73 10.6151
R912 B.n566 B.n73 10.6151
R913 B.n566 B.n565 10.6151
R914 B.n565 B.n564 10.6151
R915 B.n564 B.n75 10.6151
R916 B.n560 B.n75 10.6151
R917 B.n560 B.n559 10.6151
R918 B.n559 B.n558 10.6151
R919 B.n558 B.n77 10.6151
R920 B.n554 B.n77 10.6151
R921 B.n554 B.n553 10.6151
R922 B.n553 B.n552 10.6151
R923 B.n552 B.n79 10.6151
R924 B.n548 B.n79 10.6151
R925 B.n548 B.n547 10.6151
R926 B.n547 B.n546 10.6151
R927 B.n546 B.n81 10.6151
R928 B.n542 B.n81 10.6151
R929 B.n542 B.n541 10.6151
R930 B.n541 B.n540 10.6151
R931 B.n540 B.n83 10.6151
R932 B.n536 B.n83 10.6151
R933 B.n536 B.n535 10.6151
R934 B.n535 B.n534 10.6151
R935 B.n534 B.n85 10.6151
R936 B.n530 B.n85 10.6151
R937 B.n529 B.n528 10.6151
R938 B.n528 B.n87 10.6151
R939 B.n524 B.n87 10.6151
R940 B.n524 B.n523 10.6151
R941 B.n523 B.n522 10.6151
R942 B.n522 B.n89 10.6151
R943 B.n518 B.n89 10.6151
R944 B.n518 B.n517 10.6151
R945 B.n517 B.n516 10.6151
R946 B.n516 B.n91 10.6151
R947 B.n512 B.n91 10.6151
R948 B.n512 B.n511 10.6151
R949 B.n511 B.n510 10.6151
R950 B.n510 B.n93 10.6151
R951 B.n506 B.n93 10.6151
R952 B.n506 B.n505 10.6151
R953 B.n505 B.n504 10.6151
R954 B.n504 B.n95 10.6151
R955 B.n500 B.n95 10.6151
R956 B.n500 B.n499 10.6151
R957 B.n499 B.n498 10.6151
R958 B.n498 B.n97 10.6151
R959 B.n494 B.n97 10.6151
R960 B.n494 B.n493 10.6151
R961 B.n493 B.n492 10.6151
R962 B.n492 B.n99 10.6151
R963 B.n488 B.n99 10.6151
R964 B.n488 B.n487 10.6151
R965 B.n487 B.n486 10.6151
R966 B.n486 B.n101 10.6151
R967 B.n482 B.n101 10.6151
R968 B.n482 B.n481 10.6151
R969 B.n481 B.n480 10.6151
R970 B.n480 B.n103 10.6151
R971 B.n476 B.n103 10.6151
R972 B.n476 B.n475 10.6151
R973 B.n475 B.n474 10.6151
R974 B.n474 B.n105 10.6151
R975 B.n470 B.n105 10.6151
R976 B.n470 B.n469 10.6151
R977 B.n469 B.n468 10.6151
R978 B.n468 B.n107 10.6151
R979 B.n464 B.n107 10.6151
R980 B.n464 B.n463 10.6151
R981 B.n463 B.n462 10.6151
R982 B.n462 B.n109 10.6151
R983 B.n458 B.n109 10.6151
R984 B.n458 B.n457 10.6151
R985 B.n457 B.n456 10.6151
R986 B.n456 B.n111 10.6151
R987 B.n452 B.n111 10.6151
R988 B.n452 B.n451 10.6151
R989 B.n451 B.n450 10.6151
R990 B.n450 B.n113 10.6151
R991 B.n446 B.n113 10.6151
R992 B.n446 B.n445 10.6151
R993 B.n445 B.n444 10.6151
R994 B.n444 B.n115 10.6151
R995 B.n440 B.n115 10.6151
R996 B.n440 B.n439 10.6151
R997 B.n439 B.n438 10.6151
R998 B.n197 B.n1 10.6151
R999 B.n200 B.n197 10.6151
R1000 B.n201 B.n200 10.6151
R1001 B.n202 B.n201 10.6151
R1002 B.n202 B.n195 10.6151
R1003 B.n206 B.n195 10.6151
R1004 B.n207 B.n206 10.6151
R1005 B.n208 B.n207 10.6151
R1006 B.n208 B.n193 10.6151
R1007 B.n212 B.n193 10.6151
R1008 B.n213 B.n212 10.6151
R1009 B.n214 B.n213 10.6151
R1010 B.n214 B.n191 10.6151
R1011 B.n218 B.n191 10.6151
R1012 B.n219 B.n218 10.6151
R1013 B.n220 B.n219 10.6151
R1014 B.n220 B.n189 10.6151
R1015 B.n224 B.n189 10.6151
R1016 B.n225 B.n224 10.6151
R1017 B.n226 B.n225 10.6151
R1018 B.n226 B.n187 10.6151
R1019 B.n230 B.n187 10.6151
R1020 B.n231 B.n230 10.6151
R1021 B.n232 B.n231 10.6151
R1022 B.n232 B.n185 10.6151
R1023 B.n236 B.n185 10.6151
R1024 B.n237 B.n236 10.6151
R1025 B.n238 B.n237 10.6151
R1026 B.n238 B.n183 10.6151
R1027 B.n243 B.n242 10.6151
R1028 B.n244 B.n243 10.6151
R1029 B.n244 B.n181 10.6151
R1030 B.n248 B.n181 10.6151
R1031 B.n249 B.n248 10.6151
R1032 B.n250 B.n249 10.6151
R1033 B.n250 B.n179 10.6151
R1034 B.n254 B.n179 10.6151
R1035 B.n255 B.n254 10.6151
R1036 B.n256 B.n255 10.6151
R1037 B.n256 B.n177 10.6151
R1038 B.n260 B.n177 10.6151
R1039 B.n261 B.n260 10.6151
R1040 B.n262 B.n261 10.6151
R1041 B.n262 B.n175 10.6151
R1042 B.n266 B.n175 10.6151
R1043 B.n267 B.n266 10.6151
R1044 B.n268 B.n267 10.6151
R1045 B.n268 B.n173 10.6151
R1046 B.n272 B.n173 10.6151
R1047 B.n273 B.n272 10.6151
R1048 B.n274 B.n273 10.6151
R1049 B.n274 B.n171 10.6151
R1050 B.n278 B.n171 10.6151
R1051 B.n279 B.n278 10.6151
R1052 B.n280 B.n279 10.6151
R1053 B.n280 B.n169 10.6151
R1054 B.n284 B.n169 10.6151
R1055 B.n285 B.n284 10.6151
R1056 B.n286 B.n285 10.6151
R1057 B.n286 B.n167 10.6151
R1058 B.n290 B.n167 10.6151
R1059 B.n291 B.n290 10.6151
R1060 B.n292 B.n291 10.6151
R1061 B.n292 B.n165 10.6151
R1062 B.n296 B.n165 10.6151
R1063 B.n297 B.n296 10.6151
R1064 B.n298 B.n297 10.6151
R1065 B.n298 B.n163 10.6151
R1066 B.n302 B.n163 10.6151
R1067 B.n303 B.n302 10.6151
R1068 B.n304 B.n303 10.6151
R1069 B.n304 B.n161 10.6151
R1070 B.n308 B.n161 10.6151
R1071 B.n309 B.n308 10.6151
R1072 B.n310 B.n309 10.6151
R1073 B.n310 B.n159 10.6151
R1074 B.n314 B.n159 10.6151
R1075 B.n315 B.n314 10.6151
R1076 B.n316 B.n315 10.6151
R1077 B.n316 B.n157 10.6151
R1078 B.n320 B.n157 10.6151
R1079 B.n321 B.n320 10.6151
R1080 B.n322 B.n321 10.6151
R1081 B.n322 B.n155 10.6151
R1082 B.n326 B.n155 10.6151
R1083 B.n327 B.n326 10.6151
R1084 B.n331 B.n327 10.6151
R1085 B.n335 B.n153 10.6151
R1086 B.n336 B.n335 10.6151
R1087 B.n337 B.n336 10.6151
R1088 B.n337 B.n151 10.6151
R1089 B.n341 B.n151 10.6151
R1090 B.n342 B.n341 10.6151
R1091 B.n343 B.n342 10.6151
R1092 B.n343 B.n149 10.6151
R1093 B.n347 B.n149 10.6151
R1094 B.n350 B.n349 10.6151
R1095 B.n350 B.n145 10.6151
R1096 B.n354 B.n145 10.6151
R1097 B.n355 B.n354 10.6151
R1098 B.n356 B.n355 10.6151
R1099 B.n356 B.n143 10.6151
R1100 B.n360 B.n143 10.6151
R1101 B.n361 B.n360 10.6151
R1102 B.n362 B.n361 10.6151
R1103 B.n362 B.n141 10.6151
R1104 B.n366 B.n141 10.6151
R1105 B.n367 B.n366 10.6151
R1106 B.n368 B.n367 10.6151
R1107 B.n368 B.n139 10.6151
R1108 B.n372 B.n139 10.6151
R1109 B.n373 B.n372 10.6151
R1110 B.n374 B.n373 10.6151
R1111 B.n374 B.n137 10.6151
R1112 B.n378 B.n137 10.6151
R1113 B.n379 B.n378 10.6151
R1114 B.n380 B.n379 10.6151
R1115 B.n380 B.n135 10.6151
R1116 B.n384 B.n135 10.6151
R1117 B.n385 B.n384 10.6151
R1118 B.n386 B.n385 10.6151
R1119 B.n386 B.n133 10.6151
R1120 B.n390 B.n133 10.6151
R1121 B.n391 B.n390 10.6151
R1122 B.n392 B.n391 10.6151
R1123 B.n392 B.n131 10.6151
R1124 B.n396 B.n131 10.6151
R1125 B.n397 B.n396 10.6151
R1126 B.n398 B.n397 10.6151
R1127 B.n398 B.n129 10.6151
R1128 B.n402 B.n129 10.6151
R1129 B.n403 B.n402 10.6151
R1130 B.n404 B.n403 10.6151
R1131 B.n404 B.n127 10.6151
R1132 B.n408 B.n127 10.6151
R1133 B.n409 B.n408 10.6151
R1134 B.n410 B.n409 10.6151
R1135 B.n410 B.n125 10.6151
R1136 B.n414 B.n125 10.6151
R1137 B.n415 B.n414 10.6151
R1138 B.n416 B.n415 10.6151
R1139 B.n416 B.n123 10.6151
R1140 B.n420 B.n123 10.6151
R1141 B.n421 B.n420 10.6151
R1142 B.n422 B.n421 10.6151
R1143 B.n422 B.n121 10.6151
R1144 B.n426 B.n121 10.6151
R1145 B.n427 B.n426 10.6151
R1146 B.n428 B.n427 10.6151
R1147 B.n428 B.n119 10.6151
R1148 B.n432 B.n119 10.6151
R1149 B.n433 B.n432 10.6151
R1150 B.n434 B.n433 10.6151
R1151 B.n434 B.n117 10.6151
R1152 B.n50 B.n46 9.36635
R1153 B.n619 B.n618 9.36635
R1154 B.n331 B.n330 9.36635
R1155 B.n349 B.n348 9.36635
R1156 B.n769 B.n0 8.11757
R1157 B.n769 B.n1 8.11757
R1158 B.n633 B.n50 1.24928
R1159 B.n620 B.n619 1.24928
R1160 B.n330 B.n153 1.24928
R1161 B.n348 B.n347 1.24928
R1162 VN.n2 VN.t2 306.377
R1163 VN.n14 VN.t3 306.377
R1164 VN.n3 VN.t5 273.795
R1165 VN.n10 VN.t0 273.795
R1166 VN.n15 VN.t1 273.795
R1167 VN.n22 VN.t4 273.795
R1168 VN.n11 VN.n10 177.939
R1169 VN.n23 VN.n22 177.939
R1170 VN.n21 VN.n12 161.3
R1171 VN.n20 VN.n19 161.3
R1172 VN.n18 VN.n13 161.3
R1173 VN.n17 VN.n16 161.3
R1174 VN.n9 VN.n0 161.3
R1175 VN.n8 VN.n7 161.3
R1176 VN.n6 VN.n1 161.3
R1177 VN.n5 VN.n4 161.3
R1178 VN.n8 VN.n1 56.5193
R1179 VN.n20 VN.n13 56.5193
R1180 VN.n3 VN.n2 53.9242
R1181 VN.n15 VN.n14 53.9242
R1182 VN VN.n23 49.4759
R1183 VN.n4 VN.n1 24.4675
R1184 VN.n9 VN.n8 24.4675
R1185 VN.n16 VN.n13 24.4675
R1186 VN.n21 VN.n20 24.4675
R1187 VN.n17 VN.n14 17.9992
R1188 VN.n5 VN.n2 17.9992
R1189 VN.n4 VN.n3 12.234
R1190 VN.n16 VN.n15 12.234
R1191 VN.n10 VN.n9 7.82994
R1192 VN.n22 VN.n21 7.82994
R1193 VN.n23 VN.n12 0.189894
R1194 VN.n19 VN.n12 0.189894
R1195 VN.n19 VN.n18 0.189894
R1196 VN.n18 VN.n17 0.189894
R1197 VN.n6 VN.n5 0.189894
R1198 VN.n7 VN.n6 0.189894
R1199 VN.n7 VN.n0 0.189894
R1200 VN.n11 VN.n0 0.189894
R1201 VN VN.n11 0.0516364
R1202 VTAIL.n7 VTAIL.t9 55.3403
R1203 VTAIL.n11 VTAIL.t11 55.3401
R1204 VTAIL.n2 VTAIL.t5 55.3401
R1205 VTAIL.n10 VTAIL.t2 55.3401
R1206 VTAIL.n9 VTAIL.n8 53.5295
R1207 VTAIL.n6 VTAIL.n5 53.5295
R1208 VTAIL.n1 VTAIL.n0 53.5292
R1209 VTAIL.n4 VTAIL.n3 53.5292
R1210 VTAIL.n6 VTAIL.n4 31.1341
R1211 VTAIL.n11 VTAIL.n10 29.4876
R1212 VTAIL.n0 VTAIL.t6 1.81136
R1213 VTAIL.n0 VTAIL.t7 1.81136
R1214 VTAIL.n3 VTAIL.t0 1.81136
R1215 VTAIL.n3 VTAIL.t3 1.81136
R1216 VTAIL.n8 VTAIL.t4 1.81136
R1217 VTAIL.n8 VTAIL.t1 1.81136
R1218 VTAIL.n5 VTAIL.t10 1.81136
R1219 VTAIL.n5 VTAIL.t8 1.81136
R1220 VTAIL.n7 VTAIL.n6 1.64705
R1221 VTAIL.n10 VTAIL.n9 1.64705
R1222 VTAIL.n4 VTAIL.n2 1.64705
R1223 VTAIL.n9 VTAIL.n7 1.2936
R1224 VTAIL.n2 VTAIL.n1 1.2936
R1225 VTAIL VTAIL.n11 1.17722
R1226 VTAIL VTAIL.n1 0.470328
R1227 VDD2.n1 VDD2.t3 73.1984
R1228 VDD2.n2 VDD2.t1 72.0191
R1229 VDD2.n1 VDD2.n0 70.5643
R1230 VDD2 VDD2.n3 70.5615
R1231 VDD2.n2 VDD2.n1 44.5407
R1232 VDD2.n3 VDD2.t4 1.81136
R1233 VDD2.n3 VDD2.t2 1.81136
R1234 VDD2.n0 VDD2.t0 1.81136
R1235 VDD2.n0 VDD2.t5 1.81136
R1236 VDD2 VDD2.n2 1.2936
R1237 VP.n6 VP.t0 306.377
R1238 VP.n17 VP.t2 273.795
R1239 VP.n24 VP.t4 273.795
R1240 VP.n31 VP.t1 273.795
R1241 VP.n14 VP.t3 273.795
R1242 VP.n7 VP.t5 273.795
R1243 VP.n17 VP.n16 177.939
R1244 VP.n32 VP.n31 177.939
R1245 VP.n15 VP.n14 177.939
R1246 VP.n9 VP.n8 161.3
R1247 VP.n10 VP.n5 161.3
R1248 VP.n12 VP.n11 161.3
R1249 VP.n13 VP.n4 161.3
R1250 VP.n30 VP.n0 161.3
R1251 VP.n29 VP.n28 161.3
R1252 VP.n27 VP.n1 161.3
R1253 VP.n26 VP.n25 161.3
R1254 VP.n23 VP.n2 161.3
R1255 VP.n22 VP.n21 161.3
R1256 VP.n20 VP.n3 161.3
R1257 VP.n19 VP.n18 161.3
R1258 VP.n22 VP.n3 56.5193
R1259 VP.n29 VP.n1 56.5193
R1260 VP.n12 VP.n5 56.5193
R1261 VP.n7 VP.n6 53.9242
R1262 VP.n16 VP.n15 49.0952
R1263 VP.n18 VP.n3 24.4675
R1264 VP.n23 VP.n22 24.4675
R1265 VP.n25 VP.n1 24.4675
R1266 VP.n30 VP.n29 24.4675
R1267 VP.n13 VP.n12 24.4675
R1268 VP.n8 VP.n5 24.4675
R1269 VP.n9 VP.n6 17.9991
R1270 VP.n24 VP.n23 12.234
R1271 VP.n25 VP.n24 12.234
R1272 VP.n8 VP.n7 12.234
R1273 VP.n18 VP.n17 7.82994
R1274 VP.n31 VP.n30 7.82994
R1275 VP.n14 VP.n13 7.82994
R1276 VP.n10 VP.n9 0.189894
R1277 VP.n11 VP.n10 0.189894
R1278 VP.n11 VP.n4 0.189894
R1279 VP.n15 VP.n4 0.189894
R1280 VP.n19 VP.n16 0.189894
R1281 VP.n20 VP.n19 0.189894
R1282 VP.n21 VP.n20 0.189894
R1283 VP.n21 VP.n2 0.189894
R1284 VP.n26 VP.n2 0.189894
R1285 VP.n27 VP.n26 0.189894
R1286 VP.n28 VP.n27 0.189894
R1287 VP.n28 VP.n0 0.189894
R1288 VP.n32 VP.n0 0.189894
R1289 VP VP.n32 0.0516364
R1290 VDD1 VDD1.t5 73.3122
R1291 VDD1.n1 VDD1.t3 73.1984
R1292 VDD1.n1 VDD1.n0 70.5643
R1293 VDD1.n3 VDD1.n2 70.2081
R1294 VDD1.n3 VDD1.n1 45.947
R1295 VDD1.n2 VDD1.t0 1.81136
R1296 VDD1.n2 VDD1.t2 1.81136
R1297 VDD1.n0 VDD1.t1 1.81136
R1298 VDD1.n0 VDD1.t4 1.81136
R1299 VDD1 VDD1.n3 0.353948
C0 w_n2498_n4558# VDD2 2.51785f
C1 VDD1 B 2.27251f
C2 B VP 1.55058f
C3 w_n2498_n4558# B 9.93584f
C4 VDD1 VP 8.96701f
C5 VN VDD2 8.74885f
C6 w_n2498_n4558# VDD1 2.46553f
C7 VTAIL VDD2 10.6275f
C8 w_n2498_n4558# VP 4.91402f
C9 VN B 1.02125f
C10 VTAIL B 4.44217f
C11 VN VDD1 0.149412f
C12 VN VP 7.03729f
C13 VTAIL VDD1 10.587099f
C14 VTAIL VP 8.44177f
C15 VN w_n2498_n4558# 4.59391f
C16 VTAIL w_n2498_n4558# 3.78127f
C17 VDD2 B 2.32224f
C18 VDD2 VDD1 1.03885f
C19 VDD2 VP 0.372671f
C20 VTAIL VN 8.42721f
C21 VDD2 VSUBS 1.807258f
C22 VDD1 VSUBS 2.210118f
C23 VTAIL VSUBS 1.199512f
C24 VN VSUBS 5.26563f
C25 VP VSUBS 2.355026f
C26 B VSUBS 4.133428f
C27 w_n2498_n4558# VSUBS 0.139239p
C28 VDD1.t5 VSUBS 4.15143f
C29 VDD1.t3 VSUBS 4.15013f
C30 VDD1.t1 VSUBS 0.383378f
C31 VDD1.t4 VSUBS 0.383378f
C32 VDD1.n0 VSUBS 3.19312f
C33 VDD1.n1 VSUBS 3.80428f
C34 VDD1.t0 VSUBS 0.383378f
C35 VDD1.t2 VSUBS 0.383378f
C36 VDD1.n2 VSUBS 3.1895f
C37 VDD1.n3 VSUBS 3.5003f
C38 VP.n0 VSUBS 0.037137f
C39 VP.t1 VSUBS 2.89683f
C40 VP.n1 VSUBS 0.04956f
C41 VP.n2 VSUBS 0.037137f
C42 VP.t4 VSUBS 2.89683f
C43 VP.n3 VSUBS 0.058873f
C44 VP.n4 VSUBS 0.037137f
C45 VP.t3 VSUBS 2.89683f
C46 VP.n5 VSUBS 0.04956f
C47 VP.t0 VSUBS 3.02101f
C48 VP.n6 VSUBS 1.1104f
C49 VP.t5 VSUBS 2.89683f
C50 VP.n7 VSUBS 1.08966f
C51 VP.n8 VSUBS 0.052128f
C52 VP.n9 VSUBS 0.236002f
C53 VP.n10 VSUBS 0.037137f
C54 VP.n11 VSUBS 0.037137f
C55 VP.n12 VSUBS 0.058873f
C56 VP.n13 VSUBS 0.045977f
C57 VP.n14 VSUBS 1.09566f
C58 VP.n15 VSUBS 1.97206f
C59 VP.n16 VSUBS 1.99925f
C60 VP.t2 VSUBS 2.89683f
C61 VP.n17 VSUBS 1.09566f
C62 VP.n18 VSUBS 0.045977f
C63 VP.n19 VSUBS 0.037137f
C64 VP.n20 VSUBS 0.037137f
C65 VP.n21 VSUBS 0.037137f
C66 VP.n22 VSUBS 0.04956f
C67 VP.n23 VSUBS 0.052128f
C68 VP.n24 VSUBS 1.01805f
C69 VP.n25 VSUBS 0.052128f
C70 VP.n26 VSUBS 0.037137f
C71 VP.n27 VSUBS 0.037137f
C72 VP.n28 VSUBS 0.037137f
C73 VP.n29 VSUBS 0.058873f
C74 VP.n30 VSUBS 0.045977f
C75 VP.n31 VSUBS 1.09566f
C76 VP.n32 VSUBS 0.036785f
C77 VDD2.t3 VSUBS 4.115951f
C78 VDD2.t0 VSUBS 0.38022f
C79 VDD2.t5 VSUBS 0.38022f
C80 VDD2.n0 VSUBS 3.16682f
C81 VDD2.n1 VSUBS 3.66459f
C82 VDD2.t1 VSUBS 4.10415f
C83 VDD2.n2 VSUBS 3.5158f
C84 VDD2.t4 VSUBS 0.38022f
C85 VDD2.t2 VSUBS 0.38022f
C86 VDD2.n3 VSUBS 3.16677f
C87 VTAIL.t6 VSUBS 0.384995f
C88 VTAIL.t7 VSUBS 0.384995f
C89 VTAIL.n0 VSUBS 3.03963f
C90 VTAIL.n1 VSUBS 0.810011f
C91 VTAIL.t5 VSUBS 3.96839f
C92 VTAIL.n2 VSUBS 1.03415f
C93 VTAIL.t0 VSUBS 0.384995f
C94 VTAIL.t3 VSUBS 0.384995f
C95 VTAIL.n3 VSUBS 3.03963f
C96 VTAIL.n4 VSUBS 2.80984f
C97 VTAIL.t10 VSUBS 0.384995f
C98 VTAIL.t8 VSUBS 0.384995f
C99 VTAIL.n5 VSUBS 3.03963f
C100 VTAIL.n6 VSUBS 2.80983f
C101 VTAIL.t9 VSUBS 3.9684f
C102 VTAIL.n7 VSUBS 1.03414f
C103 VTAIL.t4 VSUBS 0.384995f
C104 VTAIL.t1 VSUBS 0.384995f
C105 VTAIL.n8 VSUBS 3.03963f
C106 VTAIL.n9 VSUBS 0.912917f
C107 VTAIL.t2 VSUBS 3.96839f
C108 VTAIL.n10 VSUBS 2.78706f
C109 VTAIL.t11 VSUBS 3.96839f
C110 VTAIL.n11 VSUBS 2.74598f
C111 VN.n0 VSUBS 0.036311f
C112 VN.t0 VSUBS 2.83246f
C113 VN.n1 VSUBS 0.048458f
C114 VN.t2 VSUBS 2.95388f
C115 VN.n2 VSUBS 1.08573f
C116 VN.t5 VSUBS 2.83246f
C117 VN.n3 VSUBS 1.06544f
C118 VN.n4 VSUBS 0.05097f
C119 VN.n5 VSUBS 0.230758f
C120 VN.n6 VSUBS 0.036311f
C121 VN.n7 VSUBS 0.036311f
C122 VN.n8 VSUBS 0.057565f
C123 VN.n9 VSUBS 0.044955f
C124 VN.n10 VSUBS 1.07132f
C125 VN.n11 VSUBS 0.035967f
C126 VN.n12 VSUBS 0.036311f
C127 VN.t4 VSUBS 2.83246f
C128 VN.n13 VSUBS 0.048458f
C129 VN.t3 VSUBS 2.95388f
C130 VN.n14 VSUBS 1.08573f
C131 VN.t1 VSUBS 2.83246f
C132 VN.n15 VSUBS 1.06544f
C133 VN.n16 VSUBS 0.05097f
C134 VN.n17 VSUBS 0.230758f
C135 VN.n18 VSUBS 0.036311f
C136 VN.n19 VSUBS 0.036311f
C137 VN.n20 VSUBS 0.057565f
C138 VN.n21 VSUBS 0.044955f
C139 VN.n22 VSUBS 1.07132f
C140 VN.n23 VSUBS 1.95187f
C141 B.n0 VSUBS 0.007005f
C142 B.n1 VSUBS 0.007005f
C143 B.n2 VSUBS 0.010361f
C144 B.n3 VSUBS 0.007939f
C145 B.n4 VSUBS 0.007939f
C146 B.n5 VSUBS 0.007939f
C147 B.n6 VSUBS 0.007939f
C148 B.n7 VSUBS 0.007939f
C149 B.n8 VSUBS 0.007939f
C150 B.n9 VSUBS 0.007939f
C151 B.n10 VSUBS 0.007939f
C152 B.n11 VSUBS 0.007939f
C153 B.n12 VSUBS 0.007939f
C154 B.n13 VSUBS 0.007939f
C155 B.n14 VSUBS 0.007939f
C156 B.n15 VSUBS 0.007939f
C157 B.n16 VSUBS 0.007939f
C158 B.n17 VSUBS 0.019037f
C159 B.n18 VSUBS 0.007939f
C160 B.n19 VSUBS 0.007939f
C161 B.n20 VSUBS 0.007939f
C162 B.n21 VSUBS 0.007939f
C163 B.n22 VSUBS 0.007939f
C164 B.n23 VSUBS 0.007939f
C165 B.n24 VSUBS 0.007939f
C166 B.n25 VSUBS 0.007939f
C167 B.n26 VSUBS 0.007939f
C168 B.n27 VSUBS 0.007939f
C169 B.n28 VSUBS 0.007939f
C170 B.n29 VSUBS 0.007939f
C171 B.n30 VSUBS 0.007939f
C172 B.n31 VSUBS 0.007939f
C173 B.n32 VSUBS 0.007939f
C174 B.n33 VSUBS 0.007939f
C175 B.n34 VSUBS 0.007939f
C176 B.n35 VSUBS 0.007939f
C177 B.n36 VSUBS 0.007939f
C178 B.n37 VSUBS 0.007939f
C179 B.n38 VSUBS 0.007939f
C180 B.n39 VSUBS 0.007939f
C181 B.n40 VSUBS 0.007939f
C182 B.n41 VSUBS 0.007939f
C183 B.n42 VSUBS 0.007939f
C184 B.n43 VSUBS 0.007939f
C185 B.n44 VSUBS 0.007939f
C186 B.n45 VSUBS 0.007939f
C187 B.n46 VSUBS 0.007472f
C188 B.n47 VSUBS 0.007939f
C189 B.t10 VSUBS 0.687208f
C190 B.t11 VSUBS 0.703588f
C191 B.t9 VSUBS 1.37368f
C192 B.n48 VSUBS 0.315029f
C193 B.n49 VSUBS 0.076973f
C194 B.n50 VSUBS 0.018395f
C195 B.n51 VSUBS 0.007939f
C196 B.n52 VSUBS 0.007939f
C197 B.n53 VSUBS 0.007939f
C198 B.n54 VSUBS 0.007939f
C199 B.t4 VSUBS 0.687183f
C200 B.t5 VSUBS 0.703567f
C201 B.t3 VSUBS 1.37368f
C202 B.n55 VSUBS 0.31505f
C203 B.n56 VSUBS 0.076997f
C204 B.n57 VSUBS 0.007939f
C205 B.n58 VSUBS 0.007939f
C206 B.n59 VSUBS 0.007939f
C207 B.n60 VSUBS 0.007939f
C208 B.n61 VSUBS 0.007939f
C209 B.n62 VSUBS 0.007939f
C210 B.n63 VSUBS 0.007939f
C211 B.n64 VSUBS 0.007939f
C212 B.n65 VSUBS 0.007939f
C213 B.n66 VSUBS 0.007939f
C214 B.n67 VSUBS 0.007939f
C215 B.n68 VSUBS 0.007939f
C216 B.n69 VSUBS 0.007939f
C217 B.n70 VSUBS 0.007939f
C218 B.n71 VSUBS 0.007939f
C219 B.n72 VSUBS 0.007939f
C220 B.n73 VSUBS 0.007939f
C221 B.n74 VSUBS 0.007939f
C222 B.n75 VSUBS 0.007939f
C223 B.n76 VSUBS 0.007939f
C224 B.n77 VSUBS 0.007939f
C225 B.n78 VSUBS 0.007939f
C226 B.n79 VSUBS 0.007939f
C227 B.n80 VSUBS 0.007939f
C228 B.n81 VSUBS 0.007939f
C229 B.n82 VSUBS 0.007939f
C230 B.n83 VSUBS 0.007939f
C231 B.n84 VSUBS 0.007939f
C232 B.n85 VSUBS 0.007939f
C233 B.n86 VSUBS 0.017858f
C234 B.n87 VSUBS 0.007939f
C235 B.n88 VSUBS 0.007939f
C236 B.n89 VSUBS 0.007939f
C237 B.n90 VSUBS 0.007939f
C238 B.n91 VSUBS 0.007939f
C239 B.n92 VSUBS 0.007939f
C240 B.n93 VSUBS 0.007939f
C241 B.n94 VSUBS 0.007939f
C242 B.n95 VSUBS 0.007939f
C243 B.n96 VSUBS 0.007939f
C244 B.n97 VSUBS 0.007939f
C245 B.n98 VSUBS 0.007939f
C246 B.n99 VSUBS 0.007939f
C247 B.n100 VSUBS 0.007939f
C248 B.n101 VSUBS 0.007939f
C249 B.n102 VSUBS 0.007939f
C250 B.n103 VSUBS 0.007939f
C251 B.n104 VSUBS 0.007939f
C252 B.n105 VSUBS 0.007939f
C253 B.n106 VSUBS 0.007939f
C254 B.n107 VSUBS 0.007939f
C255 B.n108 VSUBS 0.007939f
C256 B.n109 VSUBS 0.007939f
C257 B.n110 VSUBS 0.007939f
C258 B.n111 VSUBS 0.007939f
C259 B.n112 VSUBS 0.007939f
C260 B.n113 VSUBS 0.007939f
C261 B.n114 VSUBS 0.007939f
C262 B.n115 VSUBS 0.007939f
C263 B.n116 VSUBS 0.007939f
C264 B.n117 VSUBS 0.018089f
C265 B.n118 VSUBS 0.007939f
C266 B.n119 VSUBS 0.007939f
C267 B.n120 VSUBS 0.007939f
C268 B.n121 VSUBS 0.007939f
C269 B.n122 VSUBS 0.007939f
C270 B.n123 VSUBS 0.007939f
C271 B.n124 VSUBS 0.007939f
C272 B.n125 VSUBS 0.007939f
C273 B.n126 VSUBS 0.007939f
C274 B.n127 VSUBS 0.007939f
C275 B.n128 VSUBS 0.007939f
C276 B.n129 VSUBS 0.007939f
C277 B.n130 VSUBS 0.007939f
C278 B.n131 VSUBS 0.007939f
C279 B.n132 VSUBS 0.007939f
C280 B.n133 VSUBS 0.007939f
C281 B.n134 VSUBS 0.007939f
C282 B.n135 VSUBS 0.007939f
C283 B.n136 VSUBS 0.007939f
C284 B.n137 VSUBS 0.007939f
C285 B.n138 VSUBS 0.007939f
C286 B.n139 VSUBS 0.007939f
C287 B.n140 VSUBS 0.007939f
C288 B.n141 VSUBS 0.007939f
C289 B.n142 VSUBS 0.007939f
C290 B.n143 VSUBS 0.007939f
C291 B.n144 VSUBS 0.007939f
C292 B.n145 VSUBS 0.007939f
C293 B.n146 VSUBS 0.007939f
C294 B.t8 VSUBS 0.687183f
C295 B.t7 VSUBS 0.703567f
C296 B.t6 VSUBS 1.37368f
C297 B.n147 VSUBS 0.31505f
C298 B.n148 VSUBS 0.076997f
C299 B.n149 VSUBS 0.007939f
C300 B.n150 VSUBS 0.007939f
C301 B.n151 VSUBS 0.007939f
C302 B.n152 VSUBS 0.007939f
C303 B.n153 VSUBS 0.004437f
C304 B.n154 VSUBS 0.007939f
C305 B.n155 VSUBS 0.007939f
C306 B.n156 VSUBS 0.007939f
C307 B.n157 VSUBS 0.007939f
C308 B.n158 VSUBS 0.007939f
C309 B.n159 VSUBS 0.007939f
C310 B.n160 VSUBS 0.007939f
C311 B.n161 VSUBS 0.007939f
C312 B.n162 VSUBS 0.007939f
C313 B.n163 VSUBS 0.007939f
C314 B.n164 VSUBS 0.007939f
C315 B.n165 VSUBS 0.007939f
C316 B.n166 VSUBS 0.007939f
C317 B.n167 VSUBS 0.007939f
C318 B.n168 VSUBS 0.007939f
C319 B.n169 VSUBS 0.007939f
C320 B.n170 VSUBS 0.007939f
C321 B.n171 VSUBS 0.007939f
C322 B.n172 VSUBS 0.007939f
C323 B.n173 VSUBS 0.007939f
C324 B.n174 VSUBS 0.007939f
C325 B.n175 VSUBS 0.007939f
C326 B.n176 VSUBS 0.007939f
C327 B.n177 VSUBS 0.007939f
C328 B.n178 VSUBS 0.007939f
C329 B.n179 VSUBS 0.007939f
C330 B.n180 VSUBS 0.007939f
C331 B.n181 VSUBS 0.007939f
C332 B.n182 VSUBS 0.007939f
C333 B.n183 VSUBS 0.017858f
C334 B.n184 VSUBS 0.007939f
C335 B.n185 VSUBS 0.007939f
C336 B.n186 VSUBS 0.007939f
C337 B.n187 VSUBS 0.007939f
C338 B.n188 VSUBS 0.007939f
C339 B.n189 VSUBS 0.007939f
C340 B.n190 VSUBS 0.007939f
C341 B.n191 VSUBS 0.007939f
C342 B.n192 VSUBS 0.007939f
C343 B.n193 VSUBS 0.007939f
C344 B.n194 VSUBS 0.007939f
C345 B.n195 VSUBS 0.007939f
C346 B.n196 VSUBS 0.007939f
C347 B.n197 VSUBS 0.007939f
C348 B.n198 VSUBS 0.007939f
C349 B.n199 VSUBS 0.007939f
C350 B.n200 VSUBS 0.007939f
C351 B.n201 VSUBS 0.007939f
C352 B.n202 VSUBS 0.007939f
C353 B.n203 VSUBS 0.007939f
C354 B.n204 VSUBS 0.007939f
C355 B.n205 VSUBS 0.007939f
C356 B.n206 VSUBS 0.007939f
C357 B.n207 VSUBS 0.007939f
C358 B.n208 VSUBS 0.007939f
C359 B.n209 VSUBS 0.007939f
C360 B.n210 VSUBS 0.007939f
C361 B.n211 VSUBS 0.007939f
C362 B.n212 VSUBS 0.007939f
C363 B.n213 VSUBS 0.007939f
C364 B.n214 VSUBS 0.007939f
C365 B.n215 VSUBS 0.007939f
C366 B.n216 VSUBS 0.007939f
C367 B.n217 VSUBS 0.007939f
C368 B.n218 VSUBS 0.007939f
C369 B.n219 VSUBS 0.007939f
C370 B.n220 VSUBS 0.007939f
C371 B.n221 VSUBS 0.007939f
C372 B.n222 VSUBS 0.007939f
C373 B.n223 VSUBS 0.007939f
C374 B.n224 VSUBS 0.007939f
C375 B.n225 VSUBS 0.007939f
C376 B.n226 VSUBS 0.007939f
C377 B.n227 VSUBS 0.007939f
C378 B.n228 VSUBS 0.007939f
C379 B.n229 VSUBS 0.007939f
C380 B.n230 VSUBS 0.007939f
C381 B.n231 VSUBS 0.007939f
C382 B.n232 VSUBS 0.007939f
C383 B.n233 VSUBS 0.007939f
C384 B.n234 VSUBS 0.007939f
C385 B.n235 VSUBS 0.007939f
C386 B.n236 VSUBS 0.007939f
C387 B.n237 VSUBS 0.007939f
C388 B.n238 VSUBS 0.007939f
C389 B.n239 VSUBS 0.007939f
C390 B.n240 VSUBS 0.017858f
C391 B.n241 VSUBS 0.019037f
C392 B.n242 VSUBS 0.019037f
C393 B.n243 VSUBS 0.007939f
C394 B.n244 VSUBS 0.007939f
C395 B.n245 VSUBS 0.007939f
C396 B.n246 VSUBS 0.007939f
C397 B.n247 VSUBS 0.007939f
C398 B.n248 VSUBS 0.007939f
C399 B.n249 VSUBS 0.007939f
C400 B.n250 VSUBS 0.007939f
C401 B.n251 VSUBS 0.007939f
C402 B.n252 VSUBS 0.007939f
C403 B.n253 VSUBS 0.007939f
C404 B.n254 VSUBS 0.007939f
C405 B.n255 VSUBS 0.007939f
C406 B.n256 VSUBS 0.007939f
C407 B.n257 VSUBS 0.007939f
C408 B.n258 VSUBS 0.007939f
C409 B.n259 VSUBS 0.007939f
C410 B.n260 VSUBS 0.007939f
C411 B.n261 VSUBS 0.007939f
C412 B.n262 VSUBS 0.007939f
C413 B.n263 VSUBS 0.007939f
C414 B.n264 VSUBS 0.007939f
C415 B.n265 VSUBS 0.007939f
C416 B.n266 VSUBS 0.007939f
C417 B.n267 VSUBS 0.007939f
C418 B.n268 VSUBS 0.007939f
C419 B.n269 VSUBS 0.007939f
C420 B.n270 VSUBS 0.007939f
C421 B.n271 VSUBS 0.007939f
C422 B.n272 VSUBS 0.007939f
C423 B.n273 VSUBS 0.007939f
C424 B.n274 VSUBS 0.007939f
C425 B.n275 VSUBS 0.007939f
C426 B.n276 VSUBS 0.007939f
C427 B.n277 VSUBS 0.007939f
C428 B.n278 VSUBS 0.007939f
C429 B.n279 VSUBS 0.007939f
C430 B.n280 VSUBS 0.007939f
C431 B.n281 VSUBS 0.007939f
C432 B.n282 VSUBS 0.007939f
C433 B.n283 VSUBS 0.007939f
C434 B.n284 VSUBS 0.007939f
C435 B.n285 VSUBS 0.007939f
C436 B.n286 VSUBS 0.007939f
C437 B.n287 VSUBS 0.007939f
C438 B.n288 VSUBS 0.007939f
C439 B.n289 VSUBS 0.007939f
C440 B.n290 VSUBS 0.007939f
C441 B.n291 VSUBS 0.007939f
C442 B.n292 VSUBS 0.007939f
C443 B.n293 VSUBS 0.007939f
C444 B.n294 VSUBS 0.007939f
C445 B.n295 VSUBS 0.007939f
C446 B.n296 VSUBS 0.007939f
C447 B.n297 VSUBS 0.007939f
C448 B.n298 VSUBS 0.007939f
C449 B.n299 VSUBS 0.007939f
C450 B.n300 VSUBS 0.007939f
C451 B.n301 VSUBS 0.007939f
C452 B.n302 VSUBS 0.007939f
C453 B.n303 VSUBS 0.007939f
C454 B.n304 VSUBS 0.007939f
C455 B.n305 VSUBS 0.007939f
C456 B.n306 VSUBS 0.007939f
C457 B.n307 VSUBS 0.007939f
C458 B.n308 VSUBS 0.007939f
C459 B.n309 VSUBS 0.007939f
C460 B.n310 VSUBS 0.007939f
C461 B.n311 VSUBS 0.007939f
C462 B.n312 VSUBS 0.007939f
C463 B.n313 VSUBS 0.007939f
C464 B.n314 VSUBS 0.007939f
C465 B.n315 VSUBS 0.007939f
C466 B.n316 VSUBS 0.007939f
C467 B.n317 VSUBS 0.007939f
C468 B.n318 VSUBS 0.007939f
C469 B.n319 VSUBS 0.007939f
C470 B.n320 VSUBS 0.007939f
C471 B.n321 VSUBS 0.007939f
C472 B.n322 VSUBS 0.007939f
C473 B.n323 VSUBS 0.007939f
C474 B.n324 VSUBS 0.007939f
C475 B.n325 VSUBS 0.007939f
C476 B.n326 VSUBS 0.007939f
C477 B.n327 VSUBS 0.007939f
C478 B.t2 VSUBS 0.687208f
C479 B.t1 VSUBS 0.703588f
C480 B.t0 VSUBS 1.37368f
C481 B.n328 VSUBS 0.315029f
C482 B.n329 VSUBS 0.076973f
C483 B.n330 VSUBS 0.018395f
C484 B.n331 VSUBS 0.007472f
C485 B.n332 VSUBS 0.007939f
C486 B.n333 VSUBS 0.007939f
C487 B.n334 VSUBS 0.007939f
C488 B.n335 VSUBS 0.007939f
C489 B.n336 VSUBS 0.007939f
C490 B.n337 VSUBS 0.007939f
C491 B.n338 VSUBS 0.007939f
C492 B.n339 VSUBS 0.007939f
C493 B.n340 VSUBS 0.007939f
C494 B.n341 VSUBS 0.007939f
C495 B.n342 VSUBS 0.007939f
C496 B.n343 VSUBS 0.007939f
C497 B.n344 VSUBS 0.007939f
C498 B.n345 VSUBS 0.007939f
C499 B.n346 VSUBS 0.007939f
C500 B.n347 VSUBS 0.004437f
C501 B.n348 VSUBS 0.018395f
C502 B.n349 VSUBS 0.007472f
C503 B.n350 VSUBS 0.007939f
C504 B.n351 VSUBS 0.007939f
C505 B.n352 VSUBS 0.007939f
C506 B.n353 VSUBS 0.007939f
C507 B.n354 VSUBS 0.007939f
C508 B.n355 VSUBS 0.007939f
C509 B.n356 VSUBS 0.007939f
C510 B.n357 VSUBS 0.007939f
C511 B.n358 VSUBS 0.007939f
C512 B.n359 VSUBS 0.007939f
C513 B.n360 VSUBS 0.007939f
C514 B.n361 VSUBS 0.007939f
C515 B.n362 VSUBS 0.007939f
C516 B.n363 VSUBS 0.007939f
C517 B.n364 VSUBS 0.007939f
C518 B.n365 VSUBS 0.007939f
C519 B.n366 VSUBS 0.007939f
C520 B.n367 VSUBS 0.007939f
C521 B.n368 VSUBS 0.007939f
C522 B.n369 VSUBS 0.007939f
C523 B.n370 VSUBS 0.007939f
C524 B.n371 VSUBS 0.007939f
C525 B.n372 VSUBS 0.007939f
C526 B.n373 VSUBS 0.007939f
C527 B.n374 VSUBS 0.007939f
C528 B.n375 VSUBS 0.007939f
C529 B.n376 VSUBS 0.007939f
C530 B.n377 VSUBS 0.007939f
C531 B.n378 VSUBS 0.007939f
C532 B.n379 VSUBS 0.007939f
C533 B.n380 VSUBS 0.007939f
C534 B.n381 VSUBS 0.007939f
C535 B.n382 VSUBS 0.007939f
C536 B.n383 VSUBS 0.007939f
C537 B.n384 VSUBS 0.007939f
C538 B.n385 VSUBS 0.007939f
C539 B.n386 VSUBS 0.007939f
C540 B.n387 VSUBS 0.007939f
C541 B.n388 VSUBS 0.007939f
C542 B.n389 VSUBS 0.007939f
C543 B.n390 VSUBS 0.007939f
C544 B.n391 VSUBS 0.007939f
C545 B.n392 VSUBS 0.007939f
C546 B.n393 VSUBS 0.007939f
C547 B.n394 VSUBS 0.007939f
C548 B.n395 VSUBS 0.007939f
C549 B.n396 VSUBS 0.007939f
C550 B.n397 VSUBS 0.007939f
C551 B.n398 VSUBS 0.007939f
C552 B.n399 VSUBS 0.007939f
C553 B.n400 VSUBS 0.007939f
C554 B.n401 VSUBS 0.007939f
C555 B.n402 VSUBS 0.007939f
C556 B.n403 VSUBS 0.007939f
C557 B.n404 VSUBS 0.007939f
C558 B.n405 VSUBS 0.007939f
C559 B.n406 VSUBS 0.007939f
C560 B.n407 VSUBS 0.007939f
C561 B.n408 VSUBS 0.007939f
C562 B.n409 VSUBS 0.007939f
C563 B.n410 VSUBS 0.007939f
C564 B.n411 VSUBS 0.007939f
C565 B.n412 VSUBS 0.007939f
C566 B.n413 VSUBS 0.007939f
C567 B.n414 VSUBS 0.007939f
C568 B.n415 VSUBS 0.007939f
C569 B.n416 VSUBS 0.007939f
C570 B.n417 VSUBS 0.007939f
C571 B.n418 VSUBS 0.007939f
C572 B.n419 VSUBS 0.007939f
C573 B.n420 VSUBS 0.007939f
C574 B.n421 VSUBS 0.007939f
C575 B.n422 VSUBS 0.007939f
C576 B.n423 VSUBS 0.007939f
C577 B.n424 VSUBS 0.007939f
C578 B.n425 VSUBS 0.007939f
C579 B.n426 VSUBS 0.007939f
C580 B.n427 VSUBS 0.007939f
C581 B.n428 VSUBS 0.007939f
C582 B.n429 VSUBS 0.007939f
C583 B.n430 VSUBS 0.007939f
C584 B.n431 VSUBS 0.007939f
C585 B.n432 VSUBS 0.007939f
C586 B.n433 VSUBS 0.007939f
C587 B.n434 VSUBS 0.007939f
C588 B.n435 VSUBS 0.007939f
C589 B.n436 VSUBS 0.019037f
C590 B.n437 VSUBS 0.017858f
C591 B.n438 VSUBS 0.018806f
C592 B.n439 VSUBS 0.007939f
C593 B.n440 VSUBS 0.007939f
C594 B.n441 VSUBS 0.007939f
C595 B.n442 VSUBS 0.007939f
C596 B.n443 VSUBS 0.007939f
C597 B.n444 VSUBS 0.007939f
C598 B.n445 VSUBS 0.007939f
C599 B.n446 VSUBS 0.007939f
C600 B.n447 VSUBS 0.007939f
C601 B.n448 VSUBS 0.007939f
C602 B.n449 VSUBS 0.007939f
C603 B.n450 VSUBS 0.007939f
C604 B.n451 VSUBS 0.007939f
C605 B.n452 VSUBS 0.007939f
C606 B.n453 VSUBS 0.007939f
C607 B.n454 VSUBS 0.007939f
C608 B.n455 VSUBS 0.007939f
C609 B.n456 VSUBS 0.007939f
C610 B.n457 VSUBS 0.007939f
C611 B.n458 VSUBS 0.007939f
C612 B.n459 VSUBS 0.007939f
C613 B.n460 VSUBS 0.007939f
C614 B.n461 VSUBS 0.007939f
C615 B.n462 VSUBS 0.007939f
C616 B.n463 VSUBS 0.007939f
C617 B.n464 VSUBS 0.007939f
C618 B.n465 VSUBS 0.007939f
C619 B.n466 VSUBS 0.007939f
C620 B.n467 VSUBS 0.007939f
C621 B.n468 VSUBS 0.007939f
C622 B.n469 VSUBS 0.007939f
C623 B.n470 VSUBS 0.007939f
C624 B.n471 VSUBS 0.007939f
C625 B.n472 VSUBS 0.007939f
C626 B.n473 VSUBS 0.007939f
C627 B.n474 VSUBS 0.007939f
C628 B.n475 VSUBS 0.007939f
C629 B.n476 VSUBS 0.007939f
C630 B.n477 VSUBS 0.007939f
C631 B.n478 VSUBS 0.007939f
C632 B.n479 VSUBS 0.007939f
C633 B.n480 VSUBS 0.007939f
C634 B.n481 VSUBS 0.007939f
C635 B.n482 VSUBS 0.007939f
C636 B.n483 VSUBS 0.007939f
C637 B.n484 VSUBS 0.007939f
C638 B.n485 VSUBS 0.007939f
C639 B.n486 VSUBS 0.007939f
C640 B.n487 VSUBS 0.007939f
C641 B.n488 VSUBS 0.007939f
C642 B.n489 VSUBS 0.007939f
C643 B.n490 VSUBS 0.007939f
C644 B.n491 VSUBS 0.007939f
C645 B.n492 VSUBS 0.007939f
C646 B.n493 VSUBS 0.007939f
C647 B.n494 VSUBS 0.007939f
C648 B.n495 VSUBS 0.007939f
C649 B.n496 VSUBS 0.007939f
C650 B.n497 VSUBS 0.007939f
C651 B.n498 VSUBS 0.007939f
C652 B.n499 VSUBS 0.007939f
C653 B.n500 VSUBS 0.007939f
C654 B.n501 VSUBS 0.007939f
C655 B.n502 VSUBS 0.007939f
C656 B.n503 VSUBS 0.007939f
C657 B.n504 VSUBS 0.007939f
C658 B.n505 VSUBS 0.007939f
C659 B.n506 VSUBS 0.007939f
C660 B.n507 VSUBS 0.007939f
C661 B.n508 VSUBS 0.007939f
C662 B.n509 VSUBS 0.007939f
C663 B.n510 VSUBS 0.007939f
C664 B.n511 VSUBS 0.007939f
C665 B.n512 VSUBS 0.007939f
C666 B.n513 VSUBS 0.007939f
C667 B.n514 VSUBS 0.007939f
C668 B.n515 VSUBS 0.007939f
C669 B.n516 VSUBS 0.007939f
C670 B.n517 VSUBS 0.007939f
C671 B.n518 VSUBS 0.007939f
C672 B.n519 VSUBS 0.007939f
C673 B.n520 VSUBS 0.007939f
C674 B.n521 VSUBS 0.007939f
C675 B.n522 VSUBS 0.007939f
C676 B.n523 VSUBS 0.007939f
C677 B.n524 VSUBS 0.007939f
C678 B.n525 VSUBS 0.007939f
C679 B.n526 VSUBS 0.007939f
C680 B.n527 VSUBS 0.007939f
C681 B.n528 VSUBS 0.007939f
C682 B.n529 VSUBS 0.017858f
C683 B.n530 VSUBS 0.019037f
C684 B.n531 VSUBS 0.019037f
C685 B.n532 VSUBS 0.007939f
C686 B.n533 VSUBS 0.007939f
C687 B.n534 VSUBS 0.007939f
C688 B.n535 VSUBS 0.007939f
C689 B.n536 VSUBS 0.007939f
C690 B.n537 VSUBS 0.007939f
C691 B.n538 VSUBS 0.007939f
C692 B.n539 VSUBS 0.007939f
C693 B.n540 VSUBS 0.007939f
C694 B.n541 VSUBS 0.007939f
C695 B.n542 VSUBS 0.007939f
C696 B.n543 VSUBS 0.007939f
C697 B.n544 VSUBS 0.007939f
C698 B.n545 VSUBS 0.007939f
C699 B.n546 VSUBS 0.007939f
C700 B.n547 VSUBS 0.007939f
C701 B.n548 VSUBS 0.007939f
C702 B.n549 VSUBS 0.007939f
C703 B.n550 VSUBS 0.007939f
C704 B.n551 VSUBS 0.007939f
C705 B.n552 VSUBS 0.007939f
C706 B.n553 VSUBS 0.007939f
C707 B.n554 VSUBS 0.007939f
C708 B.n555 VSUBS 0.007939f
C709 B.n556 VSUBS 0.007939f
C710 B.n557 VSUBS 0.007939f
C711 B.n558 VSUBS 0.007939f
C712 B.n559 VSUBS 0.007939f
C713 B.n560 VSUBS 0.007939f
C714 B.n561 VSUBS 0.007939f
C715 B.n562 VSUBS 0.007939f
C716 B.n563 VSUBS 0.007939f
C717 B.n564 VSUBS 0.007939f
C718 B.n565 VSUBS 0.007939f
C719 B.n566 VSUBS 0.007939f
C720 B.n567 VSUBS 0.007939f
C721 B.n568 VSUBS 0.007939f
C722 B.n569 VSUBS 0.007939f
C723 B.n570 VSUBS 0.007939f
C724 B.n571 VSUBS 0.007939f
C725 B.n572 VSUBS 0.007939f
C726 B.n573 VSUBS 0.007939f
C727 B.n574 VSUBS 0.007939f
C728 B.n575 VSUBS 0.007939f
C729 B.n576 VSUBS 0.007939f
C730 B.n577 VSUBS 0.007939f
C731 B.n578 VSUBS 0.007939f
C732 B.n579 VSUBS 0.007939f
C733 B.n580 VSUBS 0.007939f
C734 B.n581 VSUBS 0.007939f
C735 B.n582 VSUBS 0.007939f
C736 B.n583 VSUBS 0.007939f
C737 B.n584 VSUBS 0.007939f
C738 B.n585 VSUBS 0.007939f
C739 B.n586 VSUBS 0.007939f
C740 B.n587 VSUBS 0.007939f
C741 B.n588 VSUBS 0.007939f
C742 B.n589 VSUBS 0.007939f
C743 B.n590 VSUBS 0.007939f
C744 B.n591 VSUBS 0.007939f
C745 B.n592 VSUBS 0.007939f
C746 B.n593 VSUBS 0.007939f
C747 B.n594 VSUBS 0.007939f
C748 B.n595 VSUBS 0.007939f
C749 B.n596 VSUBS 0.007939f
C750 B.n597 VSUBS 0.007939f
C751 B.n598 VSUBS 0.007939f
C752 B.n599 VSUBS 0.007939f
C753 B.n600 VSUBS 0.007939f
C754 B.n601 VSUBS 0.007939f
C755 B.n602 VSUBS 0.007939f
C756 B.n603 VSUBS 0.007939f
C757 B.n604 VSUBS 0.007939f
C758 B.n605 VSUBS 0.007939f
C759 B.n606 VSUBS 0.007939f
C760 B.n607 VSUBS 0.007939f
C761 B.n608 VSUBS 0.007939f
C762 B.n609 VSUBS 0.007939f
C763 B.n610 VSUBS 0.007939f
C764 B.n611 VSUBS 0.007939f
C765 B.n612 VSUBS 0.007939f
C766 B.n613 VSUBS 0.007939f
C767 B.n614 VSUBS 0.007939f
C768 B.n615 VSUBS 0.007939f
C769 B.n616 VSUBS 0.007939f
C770 B.n617 VSUBS 0.007939f
C771 B.n618 VSUBS 0.007472f
C772 B.n619 VSUBS 0.018395f
C773 B.n620 VSUBS 0.004437f
C774 B.n621 VSUBS 0.007939f
C775 B.n622 VSUBS 0.007939f
C776 B.n623 VSUBS 0.007939f
C777 B.n624 VSUBS 0.007939f
C778 B.n625 VSUBS 0.007939f
C779 B.n626 VSUBS 0.007939f
C780 B.n627 VSUBS 0.007939f
C781 B.n628 VSUBS 0.007939f
C782 B.n629 VSUBS 0.007939f
C783 B.n630 VSUBS 0.007939f
C784 B.n631 VSUBS 0.007939f
C785 B.n632 VSUBS 0.007939f
C786 B.n633 VSUBS 0.004437f
C787 B.n634 VSUBS 0.007939f
C788 B.n635 VSUBS 0.007939f
C789 B.n636 VSUBS 0.007939f
C790 B.n637 VSUBS 0.007939f
C791 B.n638 VSUBS 0.007939f
C792 B.n639 VSUBS 0.007939f
C793 B.n640 VSUBS 0.007939f
C794 B.n641 VSUBS 0.007939f
C795 B.n642 VSUBS 0.007939f
C796 B.n643 VSUBS 0.007939f
C797 B.n644 VSUBS 0.007939f
C798 B.n645 VSUBS 0.007939f
C799 B.n646 VSUBS 0.007939f
C800 B.n647 VSUBS 0.007939f
C801 B.n648 VSUBS 0.007939f
C802 B.n649 VSUBS 0.007939f
C803 B.n650 VSUBS 0.007939f
C804 B.n651 VSUBS 0.007939f
C805 B.n652 VSUBS 0.007939f
C806 B.n653 VSUBS 0.007939f
C807 B.n654 VSUBS 0.007939f
C808 B.n655 VSUBS 0.007939f
C809 B.n656 VSUBS 0.007939f
C810 B.n657 VSUBS 0.007939f
C811 B.n658 VSUBS 0.007939f
C812 B.n659 VSUBS 0.007939f
C813 B.n660 VSUBS 0.007939f
C814 B.n661 VSUBS 0.007939f
C815 B.n662 VSUBS 0.007939f
C816 B.n663 VSUBS 0.007939f
C817 B.n664 VSUBS 0.007939f
C818 B.n665 VSUBS 0.007939f
C819 B.n666 VSUBS 0.007939f
C820 B.n667 VSUBS 0.007939f
C821 B.n668 VSUBS 0.007939f
C822 B.n669 VSUBS 0.007939f
C823 B.n670 VSUBS 0.007939f
C824 B.n671 VSUBS 0.007939f
C825 B.n672 VSUBS 0.007939f
C826 B.n673 VSUBS 0.007939f
C827 B.n674 VSUBS 0.007939f
C828 B.n675 VSUBS 0.007939f
C829 B.n676 VSUBS 0.007939f
C830 B.n677 VSUBS 0.007939f
C831 B.n678 VSUBS 0.007939f
C832 B.n679 VSUBS 0.007939f
C833 B.n680 VSUBS 0.007939f
C834 B.n681 VSUBS 0.007939f
C835 B.n682 VSUBS 0.007939f
C836 B.n683 VSUBS 0.007939f
C837 B.n684 VSUBS 0.007939f
C838 B.n685 VSUBS 0.007939f
C839 B.n686 VSUBS 0.007939f
C840 B.n687 VSUBS 0.007939f
C841 B.n688 VSUBS 0.007939f
C842 B.n689 VSUBS 0.007939f
C843 B.n690 VSUBS 0.007939f
C844 B.n691 VSUBS 0.007939f
C845 B.n692 VSUBS 0.007939f
C846 B.n693 VSUBS 0.007939f
C847 B.n694 VSUBS 0.007939f
C848 B.n695 VSUBS 0.007939f
C849 B.n696 VSUBS 0.007939f
C850 B.n697 VSUBS 0.007939f
C851 B.n698 VSUBS 0.007939f
C852 B.n699 VSUBS 0.007939f
C853 B.n700 VSUBS 0.007939f
C854 B.n701 VSUBS 0.007939f
C855 B.n702 VSUBS 0.007939f
C856 B.n703 VSUBS 0.007939f
C857 B.n704 VSUBS 0.007939f
C858 B.n705 VSUBS 0.007939f
C859 B.n706 VSUBS 0.007939f
C860 B.n707 VSUBS 0.007939f
C861 B.n708 VSUBS 0.007939f
C862 B.n709 VSUBS 0.007939f
C863 B.n710 VSUBS 0.007939f
C864 B.n711 VSUBS 0.007939f
C865 B.n712 VSUBS 0.007939f
C866 B.n713 VSUBS 0.007939f
C867 B.n714 VSUBS 0.007939f
C868 B.n715 VSUBS 0.007939f
C869 B.n716 VSUBS 0.007939f
C870 B.n717 VSUBS 0.007939f
C871 B.n718 VSUBS 0.007939f
C872 B.n719 VSUBS 0.007939f
C873 B.n720 VSUBS 0.007939f
C874 B.n721 VSUBS 0.007939f
C875 B.n722 VSUBS 0.019037f
C876 B.n723 VSUBS 0.017858f
C877 B.n724 VSUBS 0.017858f
C878 B.n725 VSUBS 0.007939f
C879 B.n726 VSUBS 0.007939f
C880 B.n727 VSUBS 0.007939f
C881 B.n728 VSUBS 0.007939f
C882 B.n729 VSUBS 0.007939f
C883 B.n730 VSUBS 0.007939f
C884 B.n731 VSUBS 0.007939f
C885 B.n732 VSUBS 0.007939f
C886 B.n733 VSUBS 0.007939f
C887 B.n734 VSUBS 0.007939f
C888 B.n735 VSUBS 0.007939f
C889 B.n736 VSUBS 0.007939f
C890 B.n737 VSUBS 0.007939f
C891 B.n738 VSUBS 0.007939f
C892 B.n739 VSUBS 0.007939f
C893 B.n740 VSUBS 0.007939f
C894 B.n741 VSUBS 0.007939f
C895 B.n742 VSUBS 0.007939f
C896 B.n743 VSUBS 0.007939f
C897 B.n744 VSUBS 0.007939f
C898 B.n745 VSUBS 0.007939f
C899 B.n746 VSUBS 0.007939f
C900 B.n747 VSUBS 0.007939f
C901 B.n748 VSUBS 0.007939f
C902 B.n749 VSUBS 0.007939f
C903 B.n750 VSUBS 0.007939f
C904 B.n751 VSUBS 0.007939f
C905 B.n752 VSUBS 0.007939f
C906 B.n753 VSUBS 0.007939f
C907 B.n754 VSUBS 0.007939f
C908 B.n755 VSUBS 0.007939f
C909 B.n756 VSUBS 0.007939f
C910 B.n757 VSUBS 0.007939f
C911 B.n758 VSUBS 0.007939f
C912 B.n759 VSUBS 0.007939f
C913 B.n760 VSUBS 0.007939f
C914 B.n761 VSUBS 0.007939f
C915 B.n762 VSUBS 0.007939f
C916 B.n763 VSUBS 0.007939f
C917 B.n764 VSUBS 0.007939f
C918 B.n765 VSUBS 0.007939f
C919 B.n766 VSUBS 0.007939f
C920 B.n767 VSUBS 0.010361f
C921 B.n768 VSUBS 0.011037f
C922 B.n769 VSUBS 0.021948f
.ends

