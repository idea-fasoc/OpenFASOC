* NGSPICE file created from diff_pair_sample_0778.ext - technology: sky130A

.subckt diff_pair_sample_0778 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=0.45
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=0.45
X2 VTAIL.t11 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=0.45
X3 VDD1.t4 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=0.45
X4 VDD1.t3 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=0.45
X5 VDD1.t2 VP.t3 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=0.45
X6 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=0.45
X7 VDD2.t3 VN.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=0.45
X8 VDD1.t1 VP.t4 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=0.45
X9 VDD2.t5 VN.t2 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=1.1817 ps=6.84 w=3.03 l=0.45
X10 VTAIL.t4 VN.t3 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=0.45
X11 VDD2.t2 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=0.45
X12 VDD2.t1 VN.t5 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0.49995 ps=3.36 w=3.03 l=0.45
X13 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=0.45
X14 VTAIL.t1 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.49995 pd=3.36 as=0.49995 ps=3.36 w=3.03 l=0.45
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1817 pd=6.84 as=0 ps=0 w=3.03 l=0.45
R0 VN.n0 VN.t5 276.01
R1 VN.n4 VN.t1 276.01
R2 VN.n2 VN.t2 258.139
R3 VN.n6 VN.t4 258.139
R4 VN.n1 VN.t3 250.105
R5 VN.n5 VN.t0 250.105
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 71.9573
R9 VN.n3 VN.n0 71.9573
R10 VN.n2 VN.n1 40.1672
R11 VN.n6 VN.n5 40.1672
R12 VN VN.n7 33.9342
R13 VN.n5 VN.n4 17.8513
R14 VN.n1 VN.n0 17.8513
R15 VN VN.n3 0.0516364
R16 VDD2.n1 VDD2.t1 87.3384
R17 VDD2.n2 VDD2.t2 86.8896
R18 VDD2.n1 VDD2.n0 80.4676
R19 VDD2 VDD2.n3 80.4648
R20 VDD2.n2 VDD2.n1 28.5127
R21 VDD2.n3 VDD2.t4 6.53515
R22 VDD2.n3 VDD2.t3 6.53515
R23 VDD2.n0 VDD2.t0 6.53515
R24 VDD2.n0 VDD2.t5 6.53515
R25 VDD2 VDD2.n2 0.563
R26 VTAIL.n7 VTAIL.t6 70.2108
R27 VTAIL.n10 VTAIL.t8 70.2108
R28 VTAIL.n11 VTAIL.t5 70.2107
R29 VTAIL.n2 VTAIL.t0 70.2107
R30 VTAIL.n9 VTAIL.n8 63.6761
R31 VTAIL.n6 VTAIL.n5 63.6761
R32 VTAIL.n1 VTAIL.n0 63.676
R33 VTAIL.n4 VTAIL.n3 63.676
R34 VTAIL.n6 VTAIL.n4 16.3238
R35 VTAIL.n11 VTAIL.n10 15.6514
R36 VTAIL.n0 VTAIL.t2 6.53515
R37 VTAIL.n0 VTAIL.t4 6.53515
R38 VTAIL.n3 VTAIL.t10 6.53515
R39 VTAIL.n3 VTAIL.t11 6.53515
R40 VTAIL.n8 VTAIL.t9 6.53515
R41 VTAIL.n8 VTAIL.t1 6.53515
R42 VTAIL.n5 VTAIL.t3 6.53515
R43 VTAIL.n5 VTAIL.t7 6.53515
R44 VTAIL.n9 VTAIL.n7 0.806535
R45 VTAIL.n2 VTAIL.n1 0.806535
R46 VTAIL.n7 VTAIL.n6 0.672914
R47 VTAIL.n10 VTAIL.n9 0.672914
R48 VTAIL.n4 VTAIL.n2 0.672914
R49 VTAIL VTAIL.n11 0.446621
R50 VTAIL VTAIL.n1 0.226793
R51 B.n352 B.n351 585
R52 B.n138 B.n55 585
R53 B.n137 B.n136 585
R54 B.n135 B.n134 585
R55 B.n133 B.n132 585
R56 B.n131 B.n130 585
R57 B.n129 B.n128 585
R58 B.n127 B.n126 585
R59 B.n125 B.n124 585
R60 B.n123 B.n122 585
R61 B.n121 B.n120 585
R62 B.n119 B.n118 585
R63 B.n117 B.n116 585
R64 B.n115 B.n114 585
R65 B.n113 B.n112 585
R66 B.n110 B.n109 585
R67 B.n108 B.n107 585
R68 B.n106 B.n105 585
R69 B.n104 B.n103 585
R70 B.n102 B.n101 585
R71 B.n100 B.n99 585
R72 B.n98 B.n97 585
R73 B.n96 B.n95 585
R74 B.n94 B.n93 585
R75 B.n92 B.n91 585
R76 B.n89 B.n88 585
R77 B.n87 B.n86 585
R78 B.n85 B.n84 585
R79 B.n83 B.n82 585
R80 B.n81 B.n80 585
R81 B.n79 B.n78 585
R82 B.n77 B.n76 585
R83 B.n75 B.n74 585
R84 B.n73 B.n72 585
R85 B.n71 B.n70 585
R86 B.n69 B.n68 585
R87 B.n67 B.n66 585
R88 B.n65 B.n64 585
R89 B.n63 B.n62 585
R90 B.n61 B.n60 585
R91 B.n350 B.n35 585
R92 B.n355 B.n35 585
R93 B.n349 B.n34 585
R94 B.n356 B.n34 585
R95 B.n348 B.n347 585
R96 B.n347 B.n30 585
R97 B.n346 B.n29 585
R98 B.n362 B.n29 585
R99 B.n345 B.n28 585
R100 B.n363 B.n28 585
R101 B.n344 B.n27 585
R102 B.n364 B.n27 585
R103 B.n343 B.n342 585
R104 B.n342 B.n23 585
R105 B.n341 B.n22 585
R106 B.n370 B.n22 585
R107 B.n340 B.n21 585
R108 B.n371 B.n21 585
R109 B.n339 B.n20 585
R110 B.n372 B.n20 585
R111 B.n338 B.n337 585
R112 B.n337 B.n19 585
R113 B.n336 B.n15 585
R114 B.n378 B.n15 585
R115 B.n335 B.n14 585
R116 B.n379 B.n14 585
R117 B.n334 B.n13 585
R118 B.n380 B.n13 585
R119 B.n333 B.n332 585
R120 B.n332 B.n12 585
R121 B.n331 B.n330 585
R122 B.n331 B.n8 585
R123 B.n329 B.n7 585
R124 B.n387 B.n7 585
R125 B.n328 B.n6 585
R126 B.n388 B.n6 585
R127 B.n327 B.n5 585
R128 B.n389 B.n5 585
R129 B.n326 B.n325 585
R130 B.n325 B.n4 585
R131 B.n324 B.n139 585
R132 B.n324 B.n323 585
R133 B.n313 B.n140 585
R134 B.n316 B.n140 585
R135 B.n315 B.n314 585
R136 B.n317 B.n315 585
R137 B.n312 B.n144 585
R138 B.n147 B.n144 585
R139 B.n311 B.n310 585
R140 B.n310 B.n309 585
R141 B.n146 B.n145 585
R142 B.n302 B.n146 585
R143 B.n301 B.n300 585
R144 B.n303 B.n301 585
R145 B.n299 B.n152 585
R146 B.n152 B.n151 585
R147 B.n298 B.n297 585
R148 B.n297 B.n296 585
R149 B.n154 B.n153 585
R150 B.n155 B.n154 585
R151 B.n289 B.n288 585
R152 B.n290 B.n289 585
R153 B.n287 B.n159 585
R154 B.n163 B.n159 585
R155 B.n286 B.n285 585
R156 B.n285 B.n284 585
R157 B.n161 B.n160 585
R158 B.n162 B.n161 585
R159 B.n277 B.n276 585
R160 B.n278 B.n277 585
R161 B.n275 B.n168 585
R162 B.n168 B.n167 585
R163 B.n270 B.n269 585
R164 B.n268 B.n190 585
R165 B.n267 B.n189 585
R166 B.n272 B.n189 585
R167 B.n266 B.n265 585
R168 B.n264 B.n263 585
R169 B.n262 B.n261 585
R170 B.n260 B.n259 585
R171 B.n258 B.n257 585
R172 B.n256 B.n255 585
R173 B.n254 B.n253 585
R174 B.n252 B.n251 585
R175 B.n250 B.n249 585
R176 B.n248 B.n247 585
R177 B.n246 B.n245 585
R178 B.n244 B.n243 585
R179 B.n242 B.n241 585
R180 B.n240 B.n239 585
R181 B.n238 B.n237 585
R182 B.n236 B.n235 585
R183 B.n234 B.n233 585
R184 B.n232 B.n231 585
R185 B.n230 B.n229 585
R186 B.n228 B.n227 585
R187 B.n226 B.n225 585
R188 B.n224 B.n223 585
R189 B.n222 B.n221 585
R190 B.n220 B.n219 585
R191 B.n218 B.n217 585
R192 B.n216 B.n215 585
R193 B.n214 B.n213 585
R194 B.n212 B.n211 585
R195 B.n210 B.n209 585
R196 B.n208 B.n207 585
R197 B.n206 B.n205 585
R198 B.n204 B.n203 585
R199 B.n202 B.n201 585
R200 B.n200 B.n199 585
R201 B.n198 B.n197 585
R202 B.n170 B.n169 585
R203 B.n274 B.n273 585
R204 B.n273 B.n272 585
R205 B.n166 B.n165 585
R206 B.n167 B.n166 585
R207 B.n280 B.n279 585
R208 B.n279 B.n278 585
R209 B.n281 B.n164 585
R210 B.n164 B.n162 585
R211 B.n283 B.n282 585
R212 B.n284 B.n283 585
R213 B.n158 B.n157 585
R214 B.n163 B.n158 585
R215 B.n292 B.n291 585
R216 B.n291 B.n290 585
R217 B.n293 B.n156 585
R218 B.n156 B.n155 585
R219 B.n295 B.n294 585
R220 B.n296 B.n295 585
R221 B.n150 B.n149 585
R222 B.n151 B.n150 585
R223 B.n305 B.n304 585
R224 B.n304 B.n303 585
R225 B.n306 B.n148 585
R226 B.n302 B.n148 585
R227 B.n308 B.n307 585
R228 B.n309 B.n308 585
R229 B.n143 B.n142 585
R230 B.n147 B.n143 585
R231 B.n319 B.n318 585
R232 B.n318 B.n317 585
R233 B.n320 B.n141 585
R234 B.n316 B.n141 585
R235 B.n322 B.n321 585
R236 B.n323 B.n322 585
R237 B.n3 B.n0 585
R238 B.n4 B.n3 585
R239 B.n386 B.n1 585
R240 B.n387 B.n386 585
R241 B.n385 B.n384 585
R242 B.n385 B.n8 585
R243 B.n383 B.n9 585
R244 B.n12 B.n9 585
R245 B.n382 B.n381 585
R246 B.n381 B.n380 585
R247 B.n11 B.n10 585
R248 B.n379 B.n11 585
R249 B.n377 B.n376 585
R250 B.n378 B.n377 585
R251 B.n375 B.n16 585
R252 B.n19 B.n16 585
R253 B.n374 B.n373 585
R254 B.n373 B.n372 585
R255 B.n18 B.n17 585
R256 B.n371 B.n18 585
R257 B.n369 B.n368 585
R258 B.n370 B.n369 585
R259 B.n367 B.n24 585
R260 B.n24 B.n23 585
R261 B.n366 B.n365 585
R262 B.n365 B.n364 585
R263 B.n26 B.n25 585
R264 B.n363 B.n26 585
R265 B.n361 B.n360 585
R266 B.n362 B.n361 585
R267 B.n359 B.n31 585
R268 B.n31 B.n30 585
R269 B.n358 B.n357 585
R270 B.n357 B.n356 585
R271 B.n33 B.n32 585
R272 B.n355 B.n33 585
R273 B.n390 B.n389 585
R274 B.n388 B.n2 585
R275 B.n60 B.n33 468.476
R276 B.n352 B.n35 468.476
R277 B.n273 B.n168 468.476
R278 B.n270 B.n166 468.476
R279 B.n58 B.t10 370.021
R280 B.n56 B.t6 370.021
R281 B.n194 B.t13 370.021
R282 B.n191 B.t17 370.021
R283 B.n354 B.n353 256.663
R284 B.n354 B.n54 256.663
R285 B.n354 B.n53 256.663
R286 B.n354 B.n52 256.663
R287 B.n354 B.n51 256.663
R288 B.n354 B.n50 256.663
R289 B.n354 B.n49 256.663
R290 B.n354 B.n48 256.663
R291 B.n354 B.n47 256.663
R292 B.n354 B.n46 256.663
R293 B.n354 B.n45 256.663
R294 B.n354 B.n44 256.663
R295 B.n354 B.n43 256.663
R296 B.n354 B.n42 256.663
R297 B.n354 B.n41 256.663
R298 B.n354 B.n40 256.663
R299 B.n354 B.n39 256.663
R300 B.n354 B.n38 256.663
R301 B.n354 B.n37 256.663
R302 B.n354 B.n36 256.663
R303 B.n272 B.n271 256.663
R304 B.n272 B.n171 256.663
R305 B.n272 B.n172 256.663
R306 B.n272 B.n173 256.663
R307 B.n272 B.n174 256.663
R308 B.n272 B.n175 256.663
R309 B.n272 B.n176 256.663
R310 B.n272 B.n177 256.663
R311 B.n272 B.n178 256.663
R312 B.n272 B.n179 256.663
R313 B.n272 B.n180 256.663
R314 B.n272 B.n181 256.663
R315 B.n272 B.n182 256.663
R316 B.n272 B.n183 256.663
R317 B.n272 B.n184 256.663
R318 B.n272 B.n185 256.663
R319 B.n272 B.n186 256.663
R320 B.n272 B.n187 256.663
R321 B.n272 B.n188 256.663
R322 B.n392 B.n391 256.663
R323 B.n64 B.n63 163.367
R324 B.n68 B.n67 163.367
R325 B.n72 B.n71 163.367
R326 B.n76 B.n75 163.367
R327 B.n80 B.n79 163.367
R328 B.n84 B.n83 163.367
R329 B.n88 B.n87 163.367
R330 B.n93 B.n92 163.367
R331 B.n97 B.n96 163.367
R332 B.n101 B.n100 163.367
R333 B.n105 B.n104 163.367
R334 B.n109 B.n108 163.367
R335 B.n114 B.n113 163.367
R336 B.n118 B.n117 163.367
R337 B.n122 B.n121 163.367
R338 B.n126 B.n125 163.367
R339 B.n130 B.n129 163.367
R340 B.n134 B.n133 163.367
R341 B.n136 B.n55 163.367
R342 B.n277 B.n168 163.367
R343 B.n277 B.n161 163.367
R344 B.n285 B.n161 163.367
R345 B.n285 B.n159 163.367
R346 B.n289 B.n159 163.367
R347 B.n289 B.n154 163.367
R348 B.n297 B.n154 163.367
R349 B.n297 B.n152 163.367
R350 B.n301 B.n152 163.367
R351 B.n301 B.n146 163.367
R352 B.n310 B.n146 163.367
R353 B.n310 B.n144 163.367
R354 B.n315 B.n144 163.367
R355 B.n315 B.n140 163.367
R356 B.n324 B.n140 163.367
R357 B.n325 B.n324 163.367
R358 B.n325 B.n5 163.367
R359 B.n6 B.n5 163.367
R360 B.n7 B.n6 163.367
R361 B.n331 B.n7 163.367
R362 B.n332 B.n331 163.367
R363 B.n332 B.n13 163.367
R364 B.n14 B.n13 163.367
R365 B.n15 B.n14 163.367
R366 B.n337 B.n15 163.367
R367 B.n337 B.n20 163.367
R368 B.n21 B.n20 163.367
R369 B.n22 B.n21 163.367
R370 B.n342 B.n22 163.367
R371 B.n342 B.n27 163.367
R372 B.n28 B.n27 163.367
R373 B.n29 B.n28 163.367
R374 B.n347 B.n29 163.367
R375 B.n347 B.n34 163.367
R376 B.n35 B.n34 163.367
R377 B.n190 B.n189 163.367
R378 B.n265 B.n189 163.367
R379 B.n263 B.n262 163.367
R380 B.n259 B.n258 163.367
R381 B.n255 B.n254 163.367
R382 B.n251 B.n250 163.367
R383 B.n247 B.n246 163.367
R384 B.n243 B.n242 163.367
R385 B.n239 B.n238 163.367
R386 B.n235 B.n234 163.367
R387 B.n231 B.n230 163.367
R388 B.n227 B.n226 163.367
R389 B.n223 B.n222 163.367
R390 B.n219 B.n218 163.367
R391 B.n215 B.n214 163.367
R392 B.n211 B.n210 163.367
R393 B.n207 B.n206 163.367
R394 B.n203 B.n202 163.367
R395 B.n199 B.n198 163.367
R396 B.n273 B.n170 163.367
R397 B.n279 B.n166 163.367
R398 B.n279 B.n164 163.367
R399 B.n283 B.n164 163.367
R400 B.n283 B.n158 163.367
R401 B.n291 B.n158 163.367
R402 B.n291 B.n156 163.367
R403 B.n295 B.n156 163.367
R404 B.n295 B.n150 163.367
R405 B.n304 B.n150 163.367
R406 B.n304 B.n148 163.367
R407 B.n308 B.n148 163.367
R408 B.n308 B.n143 163.367
R409 B.n318 B.n143 163.367
R410 B.n318 B.n141 163.367
R411 B.n322 B.n141 163.367
R412 B.n322 B.n3 163.367
R413 B.n390 B.n3 163.367
R414 B.n386 B.n2 163.367
R415 B.n386 B.n385 163.367
R416 B.n385 B.n9 163.367
R417 B.n381 B.n9 163.367
R418 B.n381 B.n11 163.367
R419 B.n377 B.n11 163.367
R420 B.n377 B.n16 163.367
R421 B.n373 B.n16 163.367
R422 B.n373 B.n18 163.367
R423 B.n369 B.n18 163.367
R424 B.n369 B.n24 163.367
R425 B.n365 B.n24 163.367
R426 B.n365 B.n26 163.367
R427 B.n361 B.n26 163.367
R428 B.n361 B.n31 163.367
R429 B.n357 B.n31 163.367
R430 B.n357 B.n33 163.367
R431 B.n272 B.n167 144.371
R432 B.n355 B.n354 144.371
R433 B.n56 B.t8 96.2585
R434 B.n194 B.t16 96.2585
R435 B.n58 B.t11 96.2567
R436 B.n191 B.t19 96.2567
R437 B.n278 B.n167 90.0667
R438 B.n278 B.n162 90.0667
R439 B.n284 B.n162 90.0667
R440 B.n284 B.n163 90.0667
R441 B.n290 B.n155 90.0667
R442 B.n296 B.n155 90.0667
R443 B.n296 B.n151 90.0667
R444 B.n303 B.n151 90.0667
R445 B.n303 B.n302 90.0667
R446 B.n309 B.n147 90.0667
R447 B.n317 B.n316 90.0667
R448 B.n323 B.n4 90.0667
R449 B.n389 B.n4 90.0667
R450 B.n389 B.n388 90.0667
R451 B.n388 B.n387 90.0667
R452 B.n387 B.n8 90.0667
R453 B.n380 B.n12 90.0667
R454 B.n379 B.n378 90.0667
R455 B.n372 B.n19 90.0667
R456 B.n372 B.n371 90.0667
R457 B.n371 B.n370 90.0667
R458 B.n370 B.n23 90.0667
R459 B.n364 B.n23 90.0667
R460 B.n363 B.n362 90.0667
R461 B.n362 B.n30 90.0667
R462 B.n356 B.n30 90.0667
R463 B.n356 B.n355 90.0667
R464 B.n57 B.t9 81.1313
R465 B.n195 B.t15 81.1313
R466 B.n59 B.t12 81.1295
R467 B.n192 B.t18 81.1295
R468 B.n309 B.t3 75.4972
R469 B.n378 B.t4 75.4972
R470 B.n60 B.n36 71.676
R471 B.n64 B.n37 71.676
R472 B.n68 B.n38 71.676
R473 B.n72 B.n39 71.676
R474 B.n76 B.n40 71.676
R475 B.n80 B.n41 71.676
R476 B.n84 B.n42 71.676
R477 B.n88 B.n43 71.676
R478 B.n93 B.n44 71.676
R479 B.n97 B.n45 71.676
R480 B.n101 B.n46 71.676
R481 B.n105 B.n47 71.676
R482 B.n109 B.n48 71.676
R483 B.n114 B.n49 71.676
R484 B.n118 B.n50 71.676
R485 B.n122 B.n51 71.676
R486 B.n126 B.n52 71.676
R487 B.n130 B.n53 71.676
R488 B.n134 B.n54 71.676
R489 B.n353 B.n55 71.676
R490 B.n353 B.n352 71.676
R491 B.n136 B.n54 71.676
R492 B.n133 B.n53 71.676
R493 B.n129 B.n52 71.676
R494 B.n125 B.n51 71.676
R495 B.n121 B.n50 71.676
R496 B.n117 B.n49 71.676
R497 B.n113 B.n48 71.676
R498 B.n108 B.n47 71.676
R499 B.n104 B.n46 71.676
R500 B.n100 B.n45 71.676
R501 B.n96 B.n44 71.676
R502 B.n92 B.n43 71.676
R503 B.n87 B.n42 71.676
R504 B.n83 B.n41 71.676
R505 B.n79 B.n40 71.676
R506 B.n75 B.n39 71.676
R507 B.n71 B.n38 71.676
R508 B.n67 B.n37 71.676
R509 B.n63 B.n36 71.676
R510 B.n271 B.n270 71.676
R511 B.n265 B.n171 71.676
R512 B.n262 B.n172 71.676
R513 B.n258 B.n173 71.676
R514 B.n254 B.n174 71.676
R515 B.n250 B.n175 71.676
R516 B.n246 B.n176 71.676
R517 B.n242 B.n177 71.676
R518 B.n238 B.n178 71.676
R519 B.n234 B.n179 71.676
R520 B.n230 B.n180 71.676
R521 B.n226 B.n181 71.676
R522 B.n222 B.n182 71.676
R523 B.n218 B.n183 71.676
R524 B.n214 B.n184 71.676
R525 B.n210 B.n185 71.676
R526 B.n206 B.n186 71.676
R527 B.n202 B.n187 71.676
R528 B.n198 B.n188 71.676
R529 B.n271 B.n190 71.676
R530 B.n263 B.n171 71.676
R531 B.n259 B.n172 71.676
R532 B.n255 B.n173 71.676
R533 B.n251 B.n174 71.676
R534 B.n247 B.n175 71.676
R535 B.n243 B.n176 71.676
R536 B.n239 B.n177 71.676
R537 B.n235 B.n178 71.676
R538 B.n231 B.n179 71.676
R539 B.n227 B.n180 71.676
R540 B.n223 B.n181 71.676
R541 B.n219 B.n182 71.676
R542 B.n215 B.n183 71.676
R543 B.n211 B.n184 71.676
R544 B.n207 B.n185 71.676
R545 B.n203 B.n186 71.676
R546 B.n199 B.n187 71.676
R547 B.n188 B.n170 71.676
R548 B.n391 B.n390 71.676
R549 B.n391 B.n2 71.676
R550 B.n316 B.t0 67.5502
R551 B.n12 B.t2 67.5502
R552 B.n163 B.t14 59.6031
R553 B.t7 B.n363 59.6031
R554 B.n90 B.n59 59.5399
R555 B.n111 B.n57 59.5399
R556 B.n196 B.n195 59.5399
R557 B.n193 B.n192 59.5399
R558 B.n317 B.t5 49.0071
R559 B.n380 B.t1 49.0071
R560 B.n147 B.t5 41.0601
R561 B.t1 B.n379 41.0601
R562 B.n290 B.t14 30.4641
R563 B.n364 B.t7 30.4641
R564 B.n269 B.n165 30.4395
R565 B.n275 B.n274 30.4395
R566 B.n61 B.n32 30.4395
R567 B.n351 B.n350 30.4395
R568 B.n323 B.t0 22.5171
R569 B.t2 B.n8 22.5171
R570 B B.n392 18.0485
R571 B.n59 B.n58 15.1278
R572 B.n57 B.n56 15.1278
R573 B.n195 B.n194 15.1278
R574 B.n192 B.n191 15.1278
R575 B.n302 B.t3 14.57
R576 B.n19 B.t4 14.57
R577 B.n280 B.n165 10.6151
R578 B.n281 B.n280 10.6151
R579 B.n282 B.n281 10.6151
R580 B.n282 B.n157 10.6151
R581 B.n292 B.n157 10.6151
R582 B.n293 B.n292 10.6151
R583 B.n294 B.n293 10.6151
R584 B.n294 B.n149 10.6151
R585 B.n305 B.n149 10.6151
R586 B.n306 B.n305 10.6151
R587 B.n307 B.n306 10.6151
R588 B.n307 B.n142 10.6151
R589 B.n319 B.n142 10.6151
R590 B.n320 B.n319 10.6151
R591 B.n321 B.n320 10.6151
R592 B.n321 B.n0 10.6151
R593 B.n269 B.n268 10.6151
R594 B.n268 B.n267 10.6151
R595 B.n267 B.n266 10.6151
R596 B.n266 B.n264 10.6151
R597 B.n264 B.n261 10.6151
R598 B.n261 B.n260 10.6151
R599 B.n260 B.n257 10.6151
R600 B.n257 B.n256 10.6151
R601 B.n256 B.n253 10.6151
R602 B.n253 B.n252 10.6151
R603 B.n252 B.n249 10.6151
R604 B.n249 B.n248 10.6151
R605 B.n248 B.n245 10.6151
R606 B.n245 B.n244 10.6151
R607 B.n241 B.n240 10.6151
R608 B.n240 B.n237 10.6151
R609 B.n237 B.n236 10.6151
R610 B.n236 B.n233 10.6151
R611 B.n233 B.n232 10.6151
R612 B.n232 B.n229 10.6151
R613 B.n229 B.n228 10.6151
R614 B.n228 B.n225 10.6151
R615 B.n225 B.n224 10.6151
R616 B.n221 B.n220 10.6151
R617 B.n220 B.n217 10.6151
R618 B.n217 B.n216 10.6151
R619 B.n216 B.n213 10.6151
R620 B.n213 B.n212 10.6151
R621 B.n212 B.n209 10.6151
R622 B.n209 B.n208 10.6151
R623 B.n208 B.n205 10.6151
R624 B.n205 B.n204 10.6151
R625 B.n204 B.n201 10.6151
R626 B.n201 B.n200 10.6151
R627 B.n200 B.n197 10.6151
R628 B.n197 B.n169 10.6151
R629 B.n274 B.n169 10.6151
R630 B.n276 B.n275 10.6151
R631 B.n276 B.n160 10.6151
R632 B.n286 B.n160 10.6151
R633 B.n287 B.n286 10.6151
R634 B.n288 B.n287 10.6151
R635 B.n288 B.n153 10.6151
R636 B.n298 B.n153 10.6151
R637 B.n299 B.n298 10.6151
R638 B.n300 B.n299 10.6151
R639 B.n300 B.n145 10.6151
R640 B.n311 B.n145 10.6151
R641 B.n312 B.n311 10.6151
R642 B.n314 B.n312 10.6151
R643 B.n314 B.n313 10.6151
R644 B.n313 B.n139 10.6151
R645 B.n326 B.n139 10.6151
R646 B.n327 B.n326 10.6151
R647 B.n328 B.n327 10.6151
R648 B.n329 B.n328 10.6151
R649 B.n330 B.n329 10.6151
R650 B.n333 B.n330 10.6151
R651 B.n334 B.n333 10.6151
R652 B.n335 B.n334 10.6151
R653 B.n336 B.n335 10.6151
R654 B.n338 B.n336 10.6151
R655 B.n339 B.n338 10.6151
R656 B.n340 B.n339 10.6151
R657 B.n341 B.n340 10.6151
R658 B.n343 B.n341 10.6151
R659 B.n344 B.n343 10.6151
R660 B.n345 B.n344 10.6151
R661 B.n346 B.n345 10.6151
R662 B.n348 B.n346 10.6151
R663 B.n349 B.n348 10.6151
R664 B.n350 B.n349 10.6151
R665 B.n384 B.n1 10.6151
R666 B.n384 B.n383 10.6151
R667 B.n383 B.n382 10.6151
R668 B.n382 B.n10 10.6151
R669 B.n376 B.n10 10.6151
R670 B.n376 B.n375 10.6151
R671 B.n375 B.n374 10.6151
R672 B.n374 B.n17 10.6151
R673 B.n368 B.n17 10.6151
R674 B.n368 B.n367 10.6151
R675 B.n367 B.n366 10.6151
R676 B.n366 B.n25 10.6151
R677 B.n360 B.n25 10.6151
R678 B.n360 B.n359 10.6151
R679 B.n359 B.n358 10.6151
R680 B.n358 B.n32 10.6151
R681 B.n62 B.n61 10.6151
R682 B.n65 B.n62 10.6151
R683 B.n66 B.n65 10.6151
R684 B.n69 B.n66 10.6151
R685 B.n70 B.n69 10.6151
R686 B.n73 B.n70 10.6151
R687 B.n74 B.n73 10.6151
R688 B.n77 B.n74 10.6151
R689 B.n78 B.n77 10.6151
R690 B.n81 B.n78 10.6151
R691 B.n82 B.n81 10.6151
R692 B.n85 B.n82 10.6151
R693 B.n86 B.n85 10.6151
R694 B.n89 B.n86 10.6151
R695 B.n94 B.n91 10.6151
R696 B.n95 B.n94 10.6151
R697 B.n98 B.n95 10.6151
R698 B.n99 B.n98 10.6151
R699 B.n102 B.n99 10.6151
R700 B.n103 B.n102 10.6151
R701 B.n106 B.n103 10.6151
R702 B.n107 B.n106 10.6151
R703 B.n110 B.n107 10.6151
R704 B.n115 B.n112 10.6151
R705 B.n116 B.n115 10.6151
R706 B.n119 B.n116 10.6151
R707 B.n120 B.n119 10.6151
R708 B.n123 B.n120 10.6151
R709 B.n124 B.n123 10.6151
R710 B.n127 B.n124 10.6151
R711 B.n128 B.n127 10.6151
R712 B.n131 B.n128 10.6151
R713 B.n132 B.n131 10.6151
R714 B.n135 B.n132 10.6151
R715 B.n137 B.n135 10.6151
R716 B.n138 B.n137 10.6151
R717 B.n351 B.n138 10.6151
R718 B.n244 B.n193 9.36635
R719 B.n221 B.n196 9.36635
R720 B.n90 B.n89 9.36635
R721 B.n112 B.n111 9.36635
R722 B.n392 B.n0 8.11757
R723 B.n392 B.n1 8.11757
R724 B.n241 B.n193 1.24928
R725 B.n224 B.n196 1.24928
R726 B.n91 B.n90 1.24928
R727 B.n111 B.n110 1.24928
R728 VP.n1 VP.t3 276.01
R729 VP.n8 VP.t2 258.139
R730 VP.n6 VP.t1 258.139
R731 VP.n3 VP.t4 258.139
R732 VP.n7 VP.t0 250.105
R733 VP.n2 VP.t5 250.105
R734 VP.n9 VP.n8 161.3
R735 VP.n4 VP.n3 161.3
R736 VP.n7 VP.n0 161.3
R737 VP.n6 VP.n5 161.3
R738 VP.n4 VP.n1 71.9573
R739 VP.n7 VP.n6 40.1672
R740 VP.n8 VP.n7 40.1672
R741 VP.n3 VP.n2 40.1672
R742 VP.n5 VP.n4 33.5535
R743 VP.n2 VP.n1 17.8513
R744 VP.n5 VP.n0 0.189894
R745 VP.n9 VP.n0 0.189894
R746 VP VP.n9 0.0516364
R747 VDD1 VDD1.t2 87.4521
R748 VDD1.n1 VDD1.t4 87.3384
R749 VDD1.n1 VDD1.n0 80.4676
R750 VDD1.n3 VDD1.n2 80.3549
R751 VDD1.n3 VDD1.n1 29.4319
R752 VDD1.n2 VDD1.t0 6.53515
R753 VDD1.n2 VDD1.t1 6.53515
R754 VDD1.n0 VDD1.t5 6.53515
R755 VDD1.n0 VDD1.t3 6.53515
R756 VDD1 VDD1.n3 0.110414
C0 VDD1 VP 1.23207f
C1 VDD2 VDD1 0.618824f
C2 VP VN 3.18008f
C3 VP VTAIL 1.16273f
C4 VDD2 VN 1.10626f
C5 VDD2 VTAIL 4.28681f
C6 VDD1 VN 0.152862f
C7 VDD1 VTAIL 4.24972f
C8 VN VTAIL 1.14848f
C9 VDD2 VP 0.280574f
C10 VDD2 B 2.610269f
C11 VDD1 B 2.780495f
C12 VTAIL B 2.776284f
C13 VN B 5.273161f
C14 VP B 4.276602f
C15 VDD1.t2 B 0.42465f
C16 VDD1.t4 B 0.424326f
C17 VDD1.t5 B 0.04562f
C18 VDD1.t3 B 0.04562f
C19 VDD1.n0 B 0.329779f
C20 VDD1.n1 B 1.13251f
C21 VDD1.t0 B 0.04562f
C22 VDD1.t1 B 0.04562f
C23 VDD1.n2 B 0.329483f
C24 VDD1.n3 B 1.11094f
C25 VP.n0 B 0.031906f
C26 VP.t1 B 0.132759f
C27 VP.t3 B 0.137784f
C28 VP.n1 B 0.07277f
C29 VP.t5 B 0.130501f
C30 VP.n2 B 0.083055f
C31 VP.t4 B 0.132759f
C32 VP.n3 B 0.077551f
C33 VP.n4 B 0.94849f
C34 VP.n5 B 0.909071f
C35 VP.n6 B 0.077551f
C36 VP.t0 B 0.130501f
C37 VP.n7 B 0.083055f
C38 VP.t2 B 0.132759f
C39 VP.n8 B 0.077551f
C40 VP.n9 B 0.024726f
C41 VTAIL.t2 B 0.055646f
C42 VTAIL.t4 B 0.055646f
C43 VTAIL.n0 B 0.354137f
C44 VTAIL.n1 B 0.280197f
C45 VTAIL.t0 B 0.463992f
C46 VTAIL.n2 B 0.355511f
C47 VTAIL.t10 B 0.055646f
C48 VTAIL.t11 B 0.055646f
C49 VTAIL.n3 B 0.354137f
C50 VTAIL.n4 B 0.865245f
C51 VTAIL.t3 B 0.055646f
C52 VTAIL.t7 B 0.055646f
C53 VTAIL.n5 B 0.354139f
C54 VTAIL.n6 B 0.865243f
C55 VTAIL.t6 B 0.463995f
C56 VTAIL.n7 B 0.355508f
C57 VTAIL.t9 B 0.055646f
C58 VTAIL.t1 B 0.055646f
C59 VTAIL.n8 B 0.354139f
C60 VTAIL.n9 B 0.313602f
C61 VTAIL.t8 B 0.463995f
C62 VTAIL.n10 B 0.856796f
C63 VTAIL.t5 B 0.463992f
C64 VTAIL.n11 B 0.839852f
C65 VDD2.t1 B 0.441832f
C66 VDD2.t0 B 0.047503f
C67 VDD2.t5 B 0.047503f
C68 VDD2.n0 B 0.343385f
C69 VDD2.n1 B 1.12531f
C70 VDD2.t2 B 0.440656f
C71 VDD2.n2 B 1.15535f
C72 VDD2.t4 B 0.047503f
C73 VDD2.t3 B 0.047503f
C74 VDD2.n3 B 0.343373f
C75 VN.t5 B 0.135879f
C76 VN.n0 B 0.071764f
C77 VN.t3 B 0.128697f
C78 VN.n1 B 0.081907f
C79 VN.t2 B 0.130924f
C80 VN.n2 B 0.076479f
C81 VN.n3 B 0.096967f
C82 VN.t1 B 0.135879f
C83 VN.n4 B 0.071764f
C84 VN.t4 B 0.130924f
C85 VN.t0 B 0.128697f
C86 VN.n5 B 0.081907f
C87 VN.n6 B 0.076479f
C88 VN.n7 B 0.956362f
.ends

